* NGSPICE file created from tg_sample_0001.ext - technology: sky130A

.subckt tg_sample_0001 VIN VGN VGP VSS VCC VOUT
X0 VOUT.t0 VGN.t0 VIN.t0 VSS.t8 sky130_fd_pr__nfet_01v8 ad=4.9959 pd=26.4 as=4.9959 ps=26.4 w=12.81 l=3.16
X1 VSS.t7 VSS.t4 VSS.t6 VSS.t5 sky130_fd_pr__nfet_01v8 ad=4.9959 pd=26.4 as=0 ps=0 w=12.81 l=3.16
X2 VCC.t7 VCC.t4 VCC.t6 VCC.t5 sky130_fd_pr__pfet_01v8 ad=1.3221 pd=7.56 as=0 ps=0 w=3.39 l=1.3
X3 VCC.t3 VCC.t0 VCC.t2 VCC.t1 sky130_fd_pr__pfet_01v8 ad=1.3221 pd=7.56 as=0 ps=0 w=3.39 l=1.3
X4 VOUT.t1 VGP.t0 VIN.t1 VCC.t8 sky130_fd_pr__pfet_01v8 ad=1.3221 pd=7.56 as=1.3221 ps=7.56 w=3.39 l=1.3
X5 VSS.t3 VSS.t0 VSS.t2 VSS.t1 sky130_fd_pr__nfet_01v8 ad=4.9959 pd=26.4 as=0 ps=0 w=12.81 l=3.16
R0 VGN VGN.t0 137.034
R1 VIN.n10 VIN.n0 756.745
R2 VIN.n4 VIN.n3 585
R3 VIN.n9 VIN.n8 585
R4 VIN.n11 VIN.n10 585
R5 VIN.n5 VIN.t1 338.558
R6 VIN.n79 VIN.n15 289.615
R7 VIN.n80 VIN.n79 185
R8 VIN.n78 VIN.n77 185
R9 VIN.n19 VIN.n18 185
R10 VIN.n72 VIN.n71 185
R11 VIN.n70 VIN.n69 185
R12 VIN.n23 VIN.n22 185
R13 VIN.n64 VIN.n63 185
R14 VIN.n62 VIN.n61 185
R15 VIN.n60 VIN.n26 185
R16 VIN.n30 VIN.n27 185
R17 VIN.n55 VIN.n54 185
R18 VIN.n53 VIN.n52 185
R19 VIN.n32 VIN.n31 185
R20 VIN.n47 VIN.n46 185
R21 VIN.n45 VIN.n44 185
R22 VIN.n36 VIN.n35 185
R23 VIN.n39 VIN.n38 185
R24 VIN.n9 VIN.n3 171.744
R25 VIN.n10 VIN.n9 171.744
R26 VIN.t0 VIN.n37 149.524
R27 VIN.n79 VIN.n78 104.615
R28 VIN.n78 VIN.n18 104.615
R29 VIN.n71 VIN.n18 104.615
R30 VIN.n71 VIN.n70 104.615
R31 VIN.n70 VIN.n22 104.615
R32 VIN.n63 VIN.n22 104.615
R33 VIN.n63 VIN.n62 104.615
R34 VIN.n62 VIN.n26 104.615
R35 VIN.n30 VIN.n26 104.615
R36 VIN.n54 VIN.n30 104.615
R37 VIN.n54 VIN.n53 104.615
R38 VIN.n53 VIN.n31 104.615
R39 VIN.n46 VIN.n31 104.615
R40 VIN.n46 VIN.n45 104.615
R41 VIN.n45 VIN.n35 104.615
R42 VIN.n38 VIN.n35 104.615
R43 VIN.t1 VIN.n3 85.8723
R44 VIN.n38 VIN.t0 52.3082
R45 VIN VIN.n14 42.9097
R46 VIN VIN.n83 33.1122
R47 VIN.n61 VIN.n60 13.1884
R48 VIN.n64 VIN.n25 12.8005
R49 VIN.n59 VIN.n27 12.8005
R50 VIN.n65 VIN.n23 12.0247
R51 VIN.n56 VIN.n55 12.0247
R52 VIN.n69 VIN.n68 11.249
R53 VIN.n52 VIN.n29 11.249
R54 VIN.n5 VIN.n4 10.6058
R55 VIN.n72 VIN.n21 10.4732
R56 VIN.n51 VIN.n32 10.4732
R57 VIN.n39 VIN.n37 10.2747
R58 VIN.n73 VIN.n19 9.69747
R59 VIN.n48 VIN.n47 9.69747
R60 VIN.n14 VIN.n0 9.69747
R61 VIN.n83 VIN.n82 9.45567
R62 VIN.n14 VIN.n13 9.45567
R63 VIN.n41 VIN.n40 9.3005
R64 VIN.n43 VIN.n42 9.3005
R65 VIN.n34 VIN.n33 9.3005
R66 VIN.n49 VIN.n48 9.3005
R67 VIN.n51 VIN.n50 9.3005
R68 VIN.n29 VIN.n28 9.3005
R69 VIN.n57 VIN.n56 9.3005
R70 VIN.n59 VIN.n58 9.3005
R71 VIN.n82 VIN.n81 9.3005
R72 VIN.n17 VIN.n16 9.3005
R73 VIN.n76 VIN.n75 9.3005
R74 VIN.n74 VIN.n73 9.3005
R75 VIN.n21 VIN.n20 9.3005
R76 VIN.n68 VIN.n67 9.3005
R77 VIN.n66 VIN.n65 9.3005
R78 VIN.n25 VIN.n24 9.3005
R79 VIN.n7 VIN.n6 9.3005
R80 VIN.n2 VIN.n1 9.3005
R81 VIN.n13 VIN.n12 9.3005
R82 VIN.n77 VIN.n76 8.92171
R83 VIN.n44 VIN.n34 8.92171
R84 VIN.n12 VIN.n11 8.92171
R85 VIN.n80 VIN.n17 8.14595
R86 VIN.n43 VIN.n36 8.14595
R87 VIN.n8 VIN.n2 8.14595
R88 VIN.n81 VIN.n15 7.3702
R89 VIN.n40 VIN.n39 7.3702
R90 VIN.n7 VIN.n4 7.3702
R91 VIN.n83 VIN.n15 6.59444
R92 VIN.n81 VIN.n80 5.81868
R93 VIN.n40 VIN.n36 5.81868
R94 VIN.n8 VIN.n7 5.81868
R95 VIN.n77 VIN.n17 5.04292
R96 VIN.n44 VIN.n43 5.04292
R97 VIN.n11 VIN.n2 5.04292
R98 VIN.n76 VIN.n19 4.26717
R99 VIN.n47 VIN.n34 4.26717
R100 VIN.n12 VIN.n0 4.26717
R101 VIN.n73 VIN.n72 3.49141
R102 VIN.n48 VIN.n32 3.49141
R103 VIN.n41 VIN.n37 2.84303
R104 VIN.n69 VIN.n21 2.71565
R105 VIN.n52 VIN.n51 2.71565
R106 VIN.n6 VIN.n5 2.5326
R107 VIN.n68 VIN.n23 1.93989
R108 VIN.n55 VIN.n29 1.93989
R109 VIN.n65 VIN.n64 1.16414
R110 VIN.n56 VIN.n27 1.16414
R111 VIN.n61 VIN.n25 0.388379
R112 VIN.n60 VIN.n59 0.388379
R113 VIN.n82 VIN.n16 0.155672
R114 VIN.n75 VIN.n16 0.155672
R115 VIN.n75 VIN.n74 0.155672
R116 VIN.n74 VIN.n20 0.155672
R117 VIN.n67 VIN.n20 0.155672
R118 VIN.n67 VIN.n66 0.155672
R119 VIN.n66 VIN.n24 0.155672
R120 VIN.n58 VIN.n24 0.155672
R121 VIN.n58 VIN.n57 0.155672
R122 VIN.n57 VIN.n28 0.155672
R123 VIN.n50 VIN.n28 0.155672
R124 VIN.n50 VIN.n49 0.155672
R125 VIN.n49 VIN.n33 0.155672
R126 VIN.n42 VIN.n33 0.155672
R127 VIN.n42 VIN.n41 0.155672
R128 VIN.n6 VIN.n1 0.155672
R129 VIN.n13 VIN.n1 0.155672
R130 VOUT.n10 VOUT.n0 756.745
R131 VOUT.n4 VOUT.n3 585
R132 VOUT.n9 VOUT.n8 585
R133 VOUT.n11 VOUT.n10 585
R134 VOUT.n5 VOUT.t1 338.558
R135 VOUT.n79 VOUT.n15 289.615
R136 VOUT.n80 VOUT.n79 185
R137 VOUT.n78 VOUT.n77 185
R138 VOUT.n19 VOUT.n18 185
R139 VOUT.n72 VOUT.n71 185
R140 VOUT.n70 VOUT.n69 185
R141 VOUT.n23 VOUT.n22 185
R142 VOUT.n64 VOUT.n63 185
R143 VOUT.n62 VOUT.n61 185
R144 VOUT.n60 VOUT.n26 185
R145 VOUT.n30 VOUT.n27 185
R146 VOUT.n55 VOUT.n54 185
R147 VOUT.n53 VOUT.n52 185
R148 VOUT.n32 VOUT.n31 185
R149 VOUT.n47 VOUT.n46 185
R150 VOUT.n45 VOUT.n44 185
R151 VOUT.n36 VOUT.n35 185
R152 VOUT.n39 VOUT.n38 185
R153 VOUT.n9 VOUT.n3 171.744
R154 VOUT.n10 VOUT.n9 171.744
R155 VOUT.t0 VOUT.n37 149.524
R156 VOUT.n79 VOUT.n78 104.615
R157 VOUT.n78 VOUT.n18 104.615
R158 VOUT.n71 VOUT.n18 104.615
R159 VOUT.n71 VOUT.n70 104.615
R160 VOUT.n70 VOUT.n22 104.615
R161 VOUT.n63 VOUT.n22 104.615
R162 VOUT.n63 VOUT.n62 104.615
R163 VOUT.n62 VOUT.n26 104.615
R164 VOUT.n30 VOUT.n26 104.615
R165 VOUT.n54 VOUT.n30 104.615
R166 VOUT.n54 VOUT.n53 104.615
R167 VOUT.n53 VOUT.n31 104.615
R168 VOUT.n46 VOUT.n31 104.615
R169 VOUT.n46 VOUT.n45 104.615
R170 VOUT.n45 VOUT.n35 104.615
R171 VOUT.n38 VOUT.n35 104.615
R172 VOUT.t1 VOUT.n3 85.8723
R173 VOUT VOUT.n83 60.9461
R174 VOUT.n38 VOUT.t0 52.3082
R175 VOUT VOUT.n14 47.942
R176 VOUT.n61 VOUT.n60 13.1884
R177 VOUT.n64 VOUT.n25 12.8005
R178 VOUT.n59 VOUT.n27 12.8005
R179 VOUT.n65 VOUT.n23 12.0247
R180 VOUT.n56 VOUT.n55 12.0247
R181 VOUT.n69 VOUT.n68 11.249
R182 VOUT.n52 VOUT.n29 11.249
R183 VOUT.n5 VOUT.n4 10.6058
R184 VOUT.n72 VOUT.n21 10.4732
R185 VOUT.n51 VOUT.n32 10.4732
R186 VOUT.n39 VOUT.n37 10.2747
R187 VOUT.n14 VOUT.n0 9.69747
R188 VOUT.n73 VOUT.n19 9.69747
R189 VOUT.n48 VOUT.n47 9.69747
R190 VOUT.n14 VOUT.n13 9.45567
R191 VOUT.n83 VOUT.n82 9.45567
R192 VOUT.n7 VOUT.n6 9.3005
R193 VOUT.n2 VOUT.n1 9.3005
R194 VOUT.n13 VOUT.n12 9.3005
R195 VOUT.n41 VOUT.n40 9.3005
R196 VOUT.n43 VOUT.n42 9.3005
R197 VOUT.n34 VOUT.n33 9.3005
R198 VOUT.n49 VOUT.n48 9.3005
R199 VOUT.n51 VOUT.n50 9.3005
R200 VOUT.n29 VOUT.n28 9.3005
R201 VOUT.n57 VOUT.n56 9.3005
R202 VOUT.n59 VOUT.n58 9.3005
R203 VOUT.n82 VOUT.n81 9.3005
R204 VOUT.n17 VOUT.n16 9.3005
R205 VOUT.n76 VOUT.n75 9.3005
R206 VOUT.n74 VOUT.n73 9.3005
R207 VOUT.n21 VOUT.n20 9.3005
R208 VOUT.n68 VOUT.n67 9.3005
R209 VOUT.n66 VOUT.n65 9.3005
R210 VOUT.n25 VOUT.n24 9.3005
R211 VOUT.n12 VOUT.n11 8.92171
R212 VOUT.n77 VOUT.n76 8.92171
R213 VOUT.n44 VOUT.n34 8.92171
R214 VOUT.n8 VOUT.n2 8.14595
R215 VOUT.n80 VOUT.n17 8.14595
R216 VOUT.n43 VOUT.n36 8.14595
R217 VOUT.n7 VOUT.n4 7.3702
R218 VOUT.n81 VOUT.n15 7.3702
R219 VOUT.n40 VOUT.n39 7.3702
R220 VOUT.n83 VOUT.n15 6.59444
R221 VOUT.n8 VOUT.n7 5.81868
R222 VOUT.n81 VOUT.n80 5.81868
R223 VOUT.n40 VOUT.n36 5.81868
R224 VOUT.n11 VOUT.n2 5.04292
R225 VOUT.n77 VOUT.n17 5.04292
R226 VOUT.n44 VOUT.n43 5.04292
R227 VOUT.n12 VOUT.n0 4.26717
R228 VOUT.n76 VOUT.n19 4.26717
R229 VOUT.n47 VOUT.n34 4.26717
R230 VOUT.n73 VOUT.n72 3.49141
R231 VOUT.n48 VOUT.n32 3.49141
R232 VOUT.n41 VOUT.n37 2.84303
R233 VOUT.n69 VOUT.n21 2.71565
R234 VOUT.n52 VOUT.n51 2.71565
R235 VOUT.n6 VOUT.n5 2.5326
R236 VOUT.n68 VOUT.n23 1.93989
R237 VOUT.n55 VOUT.n29 1.93989
R238 VOUT.n65 VOUT.n64 1.16414
R239 VOUT.n56 VOUT.n27 1.16414
R240 VOUT.n61 VOUT.n25 0.388379
R241 VOUT.n60 VOUT.n59 0.388379
R242 VOUT.n6 VOUT.n1 0.155672
R243 VOUT.n13 VOUT.n1 0.155672
R244 VOUT.n82 VOUT.n16 0.155672
R245 VOUT.n75 VOUT.n16 0.155672
R246 VOUT.n75 VOUT.n74 0.155672
R247 VOUT.n74 VOUT.n20 0.155672
R248 VOUT.n67 VOUT.n20 0.155672
R249 VOUT.n67 VOUT.n66 0.155672
R250 VOUT.n66 VOUT.n24 0.155672
R251 VOUT.n58 VOUT.n24 0.155672
R252 VOUT.n58 VOUT.n57 0.155672
R253 VOUT.n57 VOUT.n28 0.155672
R254 VOUT.n50 VOUT.n28 0.155672
R255 VOUT.n50 VOUT.n49 0.155672
R256 VOUT.n49 VOUT.n33 0.155672
R257 VOUT.n42 VOUT.n33 0.155672
R258 VOUT.n42 VOUT.n41 0.155672
R259 VSS.n195 VSS.n79 627.038
R260 VSS.n107 VSS.n77 627.038
R261 VSS.n396 VSS.n23 627.038
R262 VSS.n398 VSS.n19 627.038
R263 VSS.n80 VSS.n79 585
R264 VSS.n79 VSS.n78 585
R265 VSS.n200 VSS.n199 585
R266 VSS.n201 VSS.n200 585
R267 VSS.n71 VSS.n70 585
R268 VSS.n72 VSS.n71 585
R269 VSS.n211 VSS.n210 585
R270 VSS.n210 VSS.n209 585
R271 VSS.n68 VSS.n67 585
R272 VSS.n67 VSS.n66 585
R273 VSS.n216 VSS.n215 585
R274 VSS.n217 VSS.n216 585
R275 VSS.n59 VSS.n58 585
R276 VSS.n60 VSS.n59 585
R277 VSS.n227 VSS.n226 585
R278 VSS.n226 VSS.n225 585
R279 VSS.n55 VSS.n53 585
R280 VSS.n53 VSS.n51 585
R281 VSS.n233 VSS.n232 585
R282 VSS.n234 VSS.n233 585
R283 VSS.n56 VSS.n54 585
R284 VSS.n54 VSS.n52 585
R285 VSS.n44 VSS.n43 585
R286 VSS.n45 VSS.n44 585
R287 VSS.n245 VSS.n244 585
R288 VSS.n244 VSS.n243 585
R289 VSS.n41 VSS.n40 585
R290 VSS.n40 VSS.t8 585
R291 VSS.n250 VSS.n249 585
R292 VSS.n251 VSS.n250 585
R293 VSS.n39 VSS.n38 585
R294 VSS.n252 VSS.n39 585
R295 VSS.n256 VSS.n255 585
R296 VSS.n255 VSS.n254 585
R297 VSS.n36 VSS.n35 585
R298 VSS.n35 VSS.n34 585
R299 VSS.n261 VSS.n260 585
R300 VSS.n262 VSS.n261 585
R301 VSS.n33 VSS.n32 585
R302 VSS.n263 VSS.n33 585
R303 VSS.n267 VSS.n266 585
R304 VSS.n266 VSS.n265 585
R305 VSS.n30 VSS.n29 585
R306 VSS.n29 VSS.n28 585
R307 VSS.n272 VSS.n271 585
R308 VSS.n273 VSS.n272 585
R309 VSS.n27 VSS.n26 585
R310 VSS.n274 VSS.n27 585
R311 VSS.n278 VSS.n277 585
R312 VSS.n277 VSS.n276 585
R313 VSS.n24 VSS.n22 585
R314 VSS.n22 VSS.n20 585
R315 VSS.n396 VSS.n395 585
R316 VSS.n397 VSS.n396 585
R317 VSS.n399 VSS.n398 585
R318 VSS.n398 VSS.n397 585
R319 VSS.n400 VSS.n18 585
R320 VSS.n20 VSS.n18 585
R321 VSS.n275 VSS.n16 585
R322 VSS.n276 VSS.n275 585
R323 VSS.n404 VSS.n15 585
R324 VSS.n274 VSS.n15 585
R325 VSS.n405 VSS.n14 585
R326 VSS.n273 VSS.n14 585
R327 VSS.n406 VSS.n13 585
R328 VSS.n28 VSS.n13 585
R329 VSS.n264 VSS.n11 585
R330 VSS.n265 VSS.n264 585
R331 VSS.n410 VSS.n10 585
R332 VSS.n263 VSS.n10 585
R333 VSS.n411 VSS.n9 585
R334 VSS.n262 VSS.n9 585
R335 VSS.n412 VSS.n8 585
R336 VSS.n34 VSS.n8 585
R337 VSS.n253 VSS.n6 585
R338 VSS.n254 VSS.n253 585
R339 VSS.n416 VSS.n5 585
R340 VSS.n252 VSS.n5 585
R341 VSS.n417 VSS.n4 585
R342 VSS.n251 VSS.n4 585
R343 VSS.n418 VSS.n3 585
R344 VSS.t8 VSS.n3 585
R345 VSS.n242 VSS.n2 585
R346 VSS.n243 VSS.n242 585
R347 VSS.n241 VSS.n240 585
R348 VSS.n241 VSS.n45 585
R349 VSS.n47 VSS.n46 585
R350 VSS.n52 VSS.n46 585
R351 VSS.n236 VSS.n235 585
R352 VSS.n235 VSS.n234 585
R353 VSS.n50 VSS.n49 585
R354 VSS.n51 VSS.n50 585
R355 VSS.n224 VSS.n223 585
R356 VSS.n225 VSS.n224 585
R357 VSS.n62 VSS.n61 585
R358 VSS.n61 VSS.n60 585
R359 VSS.n219 VSS.n218 585
R360 VSS.n218 VSS.n217 585
R361 VSS.n65 VSS.n64 585
R362 VSS.n66 VSS.n65 585
R363 VSS.n208 VSS.n207 585
R364 VSS.n209 VSS.n208 585
R365 VSS.n74 VSS.n73 585
R366 VSS.n73 VSS.n72 585
R367 VSS.n203 VSS.n202 585
R368 VSS.n202 VSS.n201 585
R369 VSS.n77 VSS.n76 585
R370 VSS.n78 VSS.n77 585
R371 VSS.n313 VSS.n19 585
R372 VSS.n317 VSS.n314 585
R373 VSS.n319 VSS.n318 585
R374 VSS.n321 VSS.n310 585
R375 VSS.n323 VSS.n322 585
R376 VSS.n325 VSS.n308 585
R377 VSS.n327 VSS.n326 585
R378 VSS.n328 VSS.n307 585
R379 VSS.n330 VSS.n329 585
R380 VSS.n332 VSS.n305 585
R381 VSS.n334 VSS.n333 585
R382 VSS.n335 VSS.n304 585
R383 VSS.n337 VSS.n336 585
R384 VSS.n339 VSS.n302 585
R385 VSS.n341 VSS.n340 585
R386 VSS.n342 VSS.n301 585
R387 VSS.n344 VSS.n343 585
R388 VSS.n346 VSS.n299 585
R389 VSS.n348 VSS.n347 585
R390 VSS.n349 VSS.n298 585
R391 VSS.n351 VSS.n350 585
R392 VSS.n353 VSS.n296 585
R393 VSS.n355 VSS.n354 585
R394 VSS.n356 VSS.n295 585
R395 VSS.n358 VSS.n357 585
R396 VSS.n360 VSS.n293 585
R397 VSS.n362 VSS.n361 585
R398 VSS.n363 VSS.n292 585
R399 VSS.n365 VSS.n364 585
R400 VSS.n367 VSS.n290 585
R401 VSS.n369 VSS.n368 585
R402 VSS.n370 VSS.n289 585
R403 VSS.n372 VSS.n371 585
R404 VSS.n374 VSS.n287 585
R405 VSS.n376 VSS.n375 585
R406 VSS.n377 VSS.n286 585
R407 VSS.n379 VSS.n378 585
R408 VSS.n381 VSS.n284 585
R409 VSS.n383 VSS.n382 585
R410 VSS.n384 VSS.n283 585
R411 VSS.n386 VSS.n385 585
R412 VSS.n388 VSS.n282 585
R413 VSS.n389 VSS.n281 585
R414 VSS.n392 VSS.n391 585
R415 VSS.n393 VSS.n23 585
R416 VSS.n23 VSS.n21 585
R417 VSS.n196 VSS.n195 585
R418 VSS.n82 VSS.n81 585
R419 VSS.n192 VSS.n191 585
R420 VSS.n193 VSS.n192 585
R421 VSS.n190 VSS.n104 585
R422 VSS.n189 VSS.n188 585
R423 VSS.n187 VSS.n186 585
R424 VSS.n185 VSS.n184 585
R425 VSS.n183 VSS.n182 585
R426 VSS.n181 VSS.n180 585
R427 VSS.n179 VSS.n178 585
R428 VSS.n177 VSS.n176 585
R429 VSS.n175 VSS.n174 585
R430 VSS.n173 VSS.n172 585
R431 VSS.n171 VSS.n170 585
R432 VSS.n169 VSS.n168 585
R433 VSS.n167 VSS.n166 585
R434 VSS.n165 VSS.n164 585
R435 VSS.n163 VSS.n162 585
R436 VSS.n161 VSS.n160 585
R437 VSS.n159 VSS.n158 585
R438 VSS.n157 VSS.n156 585
R439 VSS.n155 VSS.n154 585
R440 VSS.n153 VSS.n152 585
R441 VSS.n151 VSS.n150 585
R442 VSS.n149 VSS.n148 585
R443 VSS.n147 VSS.n146 585
R444 VSS.n145 VSS.n144 585
R445 VSS.n143 VSS.n142 585
R446 VSS.n141 VSS.n140 585
R447 VSS.n139 VSS.n138 585
R448 VSS.n137 VSS.n136 585
R449 VSS.n135 VSS.n134 585
R450 VSS.n133 VSS.n132 585
R451 VSS.n131 VSS.n130 585
R452 VSS.n129 VSS.n128 585
R453 VSS.n127 VSS.n126 585
R454 VSS.n125 VSS.n124 585
R455 VSS.n123 VSS.n122 585
R456 VSS.n121 VSS.n120 585
R457 VSS.n119 VSS.n118 585
R458 VSS.n117 VSS.n116 585
R459 VSS.n115 VSS.n114 585
R460 VSS.n112 VSS.n111 585
R461 VSS.n110 VSS.n109 585
R462 VSS.n108 VSS.n107 585
R463 VSS.n311 VSS.t2 363.926
R464 VSS.n105 VSS.t7 363.926
R465 VSS.n311 VSS.t0 306.457
R466 VSS.n105 VSS.t4 306.457
R467 VSS.n312 VSS.t3 296.241
R468 VSS.n106 VSS.t6 296.241
R469 VSS.n316 VSS.n21 256.663
R470 VSS.n315 VSS.n21 256.663
R471 VSS.n324 VSS.n21 256.663
R472 VSS.n309 VSS.n21 256.663
R473 VSS.n331 VSS.n21 256.663
R474 VSS.n306 VSS.n21 256.663
R475 VSS.n338 VSS.n21 256.663
R476 VSS.n303 VSS.n21 256.663
R477 VSS.n345 VSS.n21 256.663
R478 VSS.n300 VSS.n21 256.663
R479 VSS.n352 VSS.n21 256.663
R480 VSS.n297 VSS.n21 256.663
R481 VSS.n359 VSS.n21 256.663
R482 VSS.n294 VSS.n21 256.663
R483 VSS.n366 VSS.n21 256.663
R484 VSS.n291 VSS.n21 256.663
R485 VSS.n373 VSS.n21 256.663
R486 VSS.n288 VSS.n21 256.663
R487 VSS.n380 VSS.n21 256.663
R488 VSS.n285 VSS.n21 256.663
R489 VSS.n387 VSS.n21 256.663
R490 VSS.n390 VSS.n21 256.663
R491 VSS.n194 VSS.n193 256.663
R492 VSS.n193 VSS.n83 256.663
R493 VSS.n193 VSS.n84 256.663
R494 VSS.n193 VSS.n85 256.663
R495 VSS.n193 VSS.n86 256.663
R496 VSS.n193 VSS.n87 256.663
R497 VSS.n193 VSS.n88 256.663
R498 VSS.n193 VSS.n89 256.663
R499 VSS.n193 VSS.n90 256.663
R500 VSS.n193 VSS.n91 256.663
R501 VSS.n193 VSS.n92 256.663
R502 VSS.n193 VSS.n93 256.663
R503 VSS.n193 VSS.n94 256.663
R504 VSS.n193 VSS.n95 256.663
R505 VSS.n193 VSS.n96 256.663
R506 VSS.n193 VSS.n97 256.663
R507 VSS.n193 VSS.n98 256.663
R508 VSS.n193 VSS.n99 256.663
R509 VSS.n193 VSS.n100 256.663
R510 VSS.n193 VSS.n101 256.663
R511 VSS.n193 VSS.n102 256.663
R512 VSS.n193 VSS.n103 256.663
R513 VSS.n200 VSS.n79 240.244
R514 VSS.n200 VSS.n71 240.244
R515 VSS.n210 VSS.n71 240.244
R516 VSS.n210 VSS.n67 240.244
R517 VSS.n216 VSS.n67 240.244
R518 VSS.n216 VSS.n59 240.244
R519 VSS.n226 VSS.n59 240.244
R520 VSS.n226 VSS.n53 240.244
R521 VSS.n233 VSS.n53 240.244
R522 VSS.n233 VSS.n54 240.244
R523 VSS.n54 VSS.n44 240.244
R524 VSS.n244 VSS.n44 240.244
R525 VSS.n244 VSS.n40 240.244
R526 VSS.n250 VSS.n40 240.244
R527 VSS.n250 VSS.n39 240.244
R528 VSS.n255 VSS.n39 240.244
R529 VSS.n255 VSS.n35 240.244
R530 VSS.n261 VSS.n35 240.244
R531 VSS.n261 VSS.n33 240.244
R532 VSS.n266 VSS.n33 240.244
R533 VSS.n266 VSS.n29 240.244
R534 VSS.n272 VSS.n29 240.244
R535 VSS.n272 VSS.n27 240.244
R536 VSS.n277 VSS.n27 240.244
R537 VSS.n277 VSS.n22 240.244
R538 VSS.n396 VSS.n22 240.244
R539 VSS.n202 VSS.n77 240.244
R540 VSS.n202 VSS.n73 240.244
R541 VSS.n208 VSS.n73 240.244
R542 VSS.n208 VSS.n65 240.244
R543 VSS.n218 VSS.n65 240.244
R544 VSS.n218 VSS.n61 240.244
R545 VSS.n224 VSS.n61 240.244
R546 VSS.n224 VSS.n50 240.244
R547 VSS.n235 VSS.n50 240.244
R548 VSS.n235 VSS.n46 240.244
R549 VSS.n241 VSS.n46 240.244
R550 VSS.n242 VSS.n241 240.244
R551 VSS.n242 VSS.n3 240.244
R552 VSS.n4 VSS.n3 240.244
R553 VSS.n5 VSS.n4 240.244
R554 VSS.n253 VSS.n5 240.244
R555 VSS.n253 VSS.n8 240.244
R556 VSS.n9 VSS.n8 240.244
R557 VSS.n10 VSS.n9 240.244
R558 VSS.n264 VSS.n10 240.244
R559 VSS.n264 VSS.n13 240.244
R560 VSS.n14 VSS.n13 240.244
R561 VSS.n15 VSS.n14 240.244
R562 VSS.n275 VSS.n15 240.244
R563 VSS.n275 VSS.n18 240.244
R564 VSS.n398 VSS.n18 240.244
R565 VSS.n193 VSS.n78 231.38
R566 VSS.n397 VSS.n21 231.38
R567 VSS.n192 VSS.n82 163.367
R568 VSS.n192 VSS.n104 163.367
R569 VSS.n188 VSS.n187 163.367
R570 VSS.n184 VSS.n183 163.367
R571 VSS.n180 VSS.n179 163.367
R572 VSS.n176 VSS.n175 163.367
R573 VSS.n172 VSS.n171 163.367
R574 VSS.n168 VSS.n167 163.367
R575 VSS.n164 VSS.n163 163.367
R576 VSS.n160 VSS.n159 163.367
R577 VSS.n156 VSS.n155 163.367
R578 VSS.n152 VSS.n151 163.367
R579 VSS.n148 VSS.n147 163.367
R580 VSS.n144 VSS.n143 163.367
R581 VSS.n140 VSS.n139 163.367
R582 VSS.n136 VSS.n135 163.367
R583 VSS.n132 VSS.n131 163.367
R584 VSS.n128 VSS.n127 163.367
R585 VSS.n124 VSS.n123 163.367
R586 VSS.n120 VSS.n119 163.367
R587 VSS.n116 VSS.n115 163.367
R588 VSS.n111 VSS.n110 163.367
R589 VSS.n391 VSS.n23 163.367
R590 VSS.n389 VSS.n388 163.367
R591 VSS.n386 VSS.n283 163.367
R592 VSS.n382 VSS.n381 163.367
R593 VSS.n379 VSS.n286 163.367
R594 VSS.n375 VSS.n374 163.367
R595 VSS.n372 VSS.n289 163.367
R596 VSS.n368 VSS.n367 163.367
R597 VSS.n365 VSS.n292 163.367
R598 VSS.n361 VSS.n360 163.367
R599 VSS.n358 VSS.n295 163.367
R600 VSS.n354 VSS.n353 163.367
R601 VSS.n351 VSS.n298 163.367
R602 VSS.n347 VSS.n346 163.367
R603 VSS.n344 VSS.n301 163.367
R604 VSS.n340 VSS.n339 163.367
R605 VSS.n337 VSS.n304 163.367
R606 VSS.n333 VSS.n332 163.367
R607 VSS.n330 VSS.n307 163.367
R608 VSS.n326 VSS.n325 163.367
R609 VSS.n323 VSS.n310 163.367
R610 VSS.n318 VSS.n317 163.367
R611 VSS.n201 VSS.n78 126.438
R612 VSS.n201 VSS.n72 126.438
R613 VSS.n209 VSS.n72 126.438
R614 VSS.n217 VSS.n66 126.438
R615 VSS.n217 VSS.n60 126.438
R616 VSS.n225 VSS.n60 126.438
R617 VSS.n225 VSS.n51 126.438
R618 VSS.n234 VSS.n51 126.438
R619 VSS.n234 VSS.n52 126.438
R620 VSS.n52 VSS.n45 126.438
R621 VSS.n243 VSS.n45 126.438
R622 VSS.n243 VSS.t8 126.438
R623 VSS.n251 VSS.t8 126.438
R624 VSS.n252 VSS.n251 126.438
R625 VSS.n254 VSS.n252 126.438
R626 VSS.n254 VSS.n34 126.438
R627 VSS.n262 VSS.n34 126.438
R628 VSS.n263 VSS.n262 126.438
R629 VSS.n265 VSS.n263 126.438
R630 VSS.n265 VSS.n28 126.438
R631 VSS.n273 VSS.n28 126.438
R632 VSS.n276 VSS.n274 126.438
R633 VSS.n276 VSS.n20 126.438
R634 VSS.n397 VSS.n20 126.438
R635 VSS.n209 VSS.t5 106.207
R636 VSS.n274 VSS.t1 106.207
R637 VSS.n195 VSS.n194 71.676
R638 VSS.n104 VSS.n83 71.676
R639 VSS.n187 VSS.n84 71.676
R640 VSS.n183 VSS.n85 71.676
R641 VSS.n179 VSS.n86 71.676
R642 VSS.n175 VSS.n87 71.676
R643 VSS.n171 VSS.n88 71.676
R644 VSS.n167 VSS.n89 71.676
R645 VSS.n163 VSS.n90 71.676
R646 VSS.n159 VSS.n91 71.676
R647 VSS.n155 VSS.n92 71.676
R648 VSS.n151 VSS.n93 71.676
R649 VSS.n147 VSS.n94 71.676
R650 VSS.n143 VSS.n95 71.676
R651 VSS.n139 VSS.n96 71.676
R652 VSS.n135 VSS.n97 71.676
R653 VSS.n131 VSS.n98 71.676
R654 VSS.n127 VSS.n99 71.676
R655 VSS.n123 VSS.n100 71.676
R656 VSS.n119 VSS.n101 71.676
R657 VSS.n115 VSS.n102 71.676
R658 VSS.n110 VSS.n103 71.676
R659 VSS.n390 VSS.n389 71.676
R660 VSS.n387 VSS.n386 71.676
R661 VSS.n382 VSS.n285 71.676
R662 VSS.n380 VSS.n379 71.676
R663 VSS.n375 VSS.n288 71.676
R664 VSS.n373 VSS.n372 71.676
R665 VSS.n368 VSS.n291 71.676
R666 VSS.n366 VSS.n365 71.676
R667 VSS.n361 VSS.n294 71.676
R668 VSS.n359 VSS.n358 71.676
R669 VSS.n354 VSS.n297 71.676
R670 VSS.n352 VSS.n351 71.676
R671 VSS.n347 VSS.n300 71.676
R672 VSS.n345 VSS.n344 71.676
R673 VSS.n340 VSS.n303 71.676
R674 VSS.n338 VSS.n337 71.676
R675 VSS.n333 VSS.n306 71.676
R676 VSS.n331 VSS.n330 71.676
R677 VSS.n326 VSS.n309 71.676
R678 VSS.n324 VSS.n323 71.676
R679 VSS.n318 VSS.n315 71.676
R680 VSS.n316 VSS.n19 71.676
R681 VSS.n317 VSS.n316 71.676
R682 VSS.n315 VSS.n310 71.676
R683 VSS.n325 VSS.n324 71.676
R684 VSS.n309 VSS.n307 71.676
R685 VSS.n332 VSS.n331 71.676
R686 VSS.n306 VSS.n304 71.676
R687 VSS.n339 VSS.n338 71.676
R688 VSS.n303 VSS.n301 71.676
R689 VSS.n346 VSS.n345 71.676
R690 VSS.n300 VSS.n298 71.676
R691 VSS.n353 VSS.n352 71.676
R692 VSS.n297 VSS.n295 71.676
R693 VSS.n360 VSS.n359 71.676
R694 VSS.n294 VSS.n292 71.676
R695 VSS.n367 VSS.n366 71.676
R696 VSS.n291 VSS.n289 71.676
R697 VSS.n374 VSS.n373 71.676
R698 VSS.n288 VSS.n286 71.676
R699 VSS.n381 VSS.n380 71.676
R700 VSS.n285 VSS.n283 71.676
R701 VSS.n388 VSS.n387 71.676
R702 VSS.n391 VSS.n390 71.676
R703 VSS.n194 VSS.n82 71.676
R704 VSS.n188 VSS.n83 71.676
R705 VSS.n184 VSS.n84 71.676
R706 VSS.n180 VSS.n85 71.676
R707 VSS.n176 VSS.n86 71.676
R708 VSS.n172 VSS.n87 71.676
R709 VSS.n168 VSS.n88 71.676
R710 VSS.n164 VSS.n89 71.676
R711 VSS.n160 VSS.n90 71.676
R712 VSS.n156 VSS.n91 71.676
R713 VSS.n152 VSS.n92 71.676
R714 VSS.n148 VSS.n93 71.676
R715 VSS.n144 VSS.n94 71.676
R716 VSS.n140 VSS.n95 71.676
R717 VSS.n136 VSS.n96 71.676
R718 VSS.n132 VSS.n97 71.676
R719 VSS.n128 VSS.n98 71.676
R720 VSS.n124 VSS.n99 71.676
R721 VSS.n120 VSS.n100 71.676
R722 VSS.n116 VSS.n101 71.676
R723 VSS.n111 VSS.n102 71.676
R724 VSS.n107 VSS.n103 71.676
R725 VSS.n312 VSS.n311 67.6854
R726 VSS.n106 VSS.n105 67.6854
R727 VSS.n320 VSS.n312 34.3278
R728 VSS.n113 VSS.n106 34.3278
R729 VSS.n394 VSS.n393 28.1551
R730 VSS.n313 VSS.n17 28.1551
R731 VSS.n197 VSS.n196 28.1551
R732 VSS.n108 VSS.n75 28.1551
R733 VSS.t5 VSS.n66 20.2304
R734 VSS.t1 VSS.n273 20.2304
R735 VSS.n199 VSS.n80 19.3944
R736 VSS.n199 VSS.n70 19.3944
R737 VSS.n211 VSS.n70 19.3944
R738 VSS.n211 VSS.n68 19.3944
R739 VSS.n215 VSS.n68 19.3944
R740 VSS.n215 VSS.n58 19.3944
R741 VSS.n227 VSS.n58 19.3944
R742 VSS.n227 VSS.n55 19.3944
R743 VSS.n232 VSS.n55 19.3944
R744 VSS.n232 VSS.n56 19.3944
R745 VSS.n56 VSS.n43 19.3944
R746 VSS.n245 VSS.n43 19.3944
R747 VSS.n245 VSS.n41 19.3944
R748 VSS.n249 VSS.n41 19.3944
R749 VSS.n249 VSS.n38 19.3944
R750 VSS.n256 VSS.n38 19.3944
R751 VSS.n256 VSS.n36 19.3944
R752 VSS.n260 VSS.n36 19.3944
R753 VSS.n260 VSS.n32 19.3944
R754 VSS.n267 VSS.n32 19.3944
R755 VSS.n267 VSS.n30 19.3944
R756 VSS.n271 VSS.n30 19.3944
R757 VSS.n271 VSS.n26 19.3944
R758 VSS.n278 VSS.n26 19.3944
R759 VSS.n278 VSS.n24 19.3944
R760 VSS.n395 VSS.n24 19.3944
R761 VSS.n203 VSS.n76 19.3944
R762 VSS.n203 VSS.n74 19.3944
R763 VSS.n207 VSS.n74 19.3944
R764 VSS.n207 VSS.n64 19.3944
R765 VSS.n219 VSS.n64 19.3944
R766 VSS.n219 VSS.n62 19.3944
R767 VSS.n223 VSS.n62 19.3944
R768 VSS.n223 VSS.n49 19.3944
R769 VSS.n236 VSS.n49 19.3944
R770 VSS.n236 VSS.n47 19.3944
R771 VSS.n240 VSS.n47 19.3944
R772 VSS.n240 VSS.n2 19.3944
R773 VSS.n418 VSS.n2 19.3944
R774 VSS.n418 VSS.n417 19.3944
R775 VSS.n417 VSS.n416 19.3944
R776 VSS.n416 VSS.n6 19.3944
R777 VSS.n412 VSS.n6 19.3944
R778 VSS.n412 VSS.n411 19.3944
R779 VSS.n411 VSS.n410 19.3944
R780 VSS.n410 VSS.n11 19.3944
R781 VSS.n406 VSS.n11 19.3944
R782 VSS.n406 VSS.n405 19.3944
R783 VSS.n405 VSS.n404 19.3944
R784 VSS.n404 VSS.n16 19.3944
R785 VSS.n400 VSS.n16 19.3944
R786 VSS.n400 VSS.n399 19.3944
R787 VSS.n393 VSS.n392 10.6151
R788 VSS.n392 VSS.n281 10.6151
R789 VSS.n282 VSS.n281 10.6151
R790 VSS.n385 VSS.n282 10.6151
R791 VSS.n385 VSS.n384 10.6151
R792 VSS.n384 VSS.n383 10.6151
R793 VSS.n383 VSS.n284 10.6151
R794 VSS.n378 VSS.n284 10.6151
R795 VSS.n378 VSS.n377 10.6151
R796 VSS.n377 VSS.n376 10.6151
R797 VSS.n376 VSS.n287 10.6151
R798 VSS.n371 VSS.n287 10.6151
R799 VSS.n371 VSS.n370 10.6151
R800 VSS.n370 VSS.n369 10.6151
R801 VSS.n369 VSS.n290 10.6151
R802 VSS.n364 VSS.n290 10.6151
R803 VSS.n364 VSS.n363 10.6151
R804 VSS.n363 VSS.n362 10.6151
R805 VSS.n362 VSS.n293 10.6151
R806 VSS.n357 VSS.n293 10.6151
R807 VSS.n357 VSS.n356 10.6151
R808 VSS.n356 VSS.n355 10.6151
R809 VSS.n355 VSS.n296 10.6151
R810 VSS.n350 VSS.n296 10.6151
R811 VSS.n350 VSS.n349 10.6151
R812 VSS.n349 VSS.n348 10.6151
R813 VSS.n348 VSS.n299 10.6151
R814 VSS.n343 VSS.n299 10.6151
R815 VSS.n343 VSS.n342 10.6151
R816 VSS.n342 VSS.n341 10.6151
R817 VSS.n341 VSS.n302 10.6151
R818 VSS.n336 VSS.n302 10.6151
R819 VSS.n336 VSS.n335 10.6151
R820 VSS.n335 VSS.n334 10.6151
R821 VSS.n334 VSS.n305 10.6151
R822 VSS.n329 VSS.n305 10.6151
R823 VSS.n329 VSS.n328 10.6151
R824 VSS.n328 VSS.n327 10.6151
R825 VSS.n327 VSS.n308 10.6151
R826 VSS.n322 VSS.n308 10.6151
R827 VSS.n322 VSS.n321 10.6151
R828 VSS.n319 VSS.n314 10.6151
R829 VSS.n314 VSS.n313 10.6151
R830 VSS.n196 VSS.n81 10.6151
R831 VSS.n191 VSS.n81 10.6151
R832 VSS.n191 VSS.n190 10.6151
R833 VSS.n190 VSS.n189 10.6151
R834 VSS.n189 VSS.n186 10.6151
R835 VSS.n186 VSS.n185 10.6151
R836 VSS.n185 VSS.n182 10.6151
R837 VSS.n182 VSS.n181 10.6151
R838 VSS.n181 VSS.n178 10.6151
R839 VSS.n178 VSS.n177 10.6151
R840 VSS.n177 VSS.n174 10.6151
R841 VSS.n174 VSS.n173 10.6151
R842 VSS.n173 VSS.n170 10.6151
R843 VSS.n170 VSS.n169 10.6151
R844 VSS.n169 VSS.n166 10.6151
R845 VSS.n166 VSS.n165 10.6151
R846 VSS.n165 VSS.n162 10.6151
R847 VSS.n162 VSS.n161 10.6151
R848 VSS.n161 VSS.n158 10.6151
R849 VSS.n158 VSS.n157 10.6151
R850 VSS.n157 VSS.n154 10.6151
R851 VSS.n154 VSS.n153 10.6151
R852 VSS.n153 VSS.n150 10.6151
R853 VSS.n150 VSS.n149 10.6151
R854 VSS.n149 VSS.n146 10.6151
R855 VSS.n146 VSS.n145 10.6151
R856 VSS.n145 VSS.n142 10.6151
R857 VSS.n142 VSS.n141 10.6151
R858 VSS.n141 VSS.n138 10.6151
R859 VSS.n138 VSS.n137 10.6151
R860 VSS.n137 VSS.n134 10.6151
R861 VSS.n134 VSS.n133 10.6151
R862 VSS.n133 VSS.n130 10.6151
R863 VSS.n130 VSS.n129 10.6151
R864 VSS.n129 VSS.n126 10.6151
R865 VSS.n126 VSS.n125 10.6151
R866 VSS.n125 VSS.n122 10.6151
R867 VSS.n122 VSS.n121 10.6151
R868 VSS.n121 VSS.n118 10.6151
R869 VSS.n118 VSS.n117 10.6151
R870 VSS.n117 VSS.n114 10.6151
R871 VSS.n112 VSS.n109 10.6151
R872 VSS.n109 VSS.n108 10.6151
R873 VSS.n417 VSS.n0 9.3005
R874 VSS.n416 VSS.n415 9.3005
R875 VSS.n414 VSS.n6 9.3005
R876 VSS.n413 VSS.n412 9.3005
R877 VSS.n411 VSS.n7 9.3005
R878 VSS.n410 VSS.n409 9.3005
R879 VSS.n408 VSS.n11 9.3005
R880 VSS.n407 VSS.n406 9.3005
R881 VSS.n405 VSS.n12 9.3005
R882 VSS.n404 VSS.n403 9.3005
R883 VSS.n402 VSS.n16 9.3005
R884 VSS.n401 VSS.n400 9.3005
R885 VSS.n399 VSS.n17 9.3005
R886 VSS.n197 VSS.n80 9.3005
R887 VSS.n199 VSS.n198 9.3005
R888 VSS.n70 VSS.n69 9.3005
R889 VSS.n212 VSS.n211 9.3005
R890 VSS.n213 VSS.n68 9.3005
R891 VSS.n215 VSS.n214 9.3005
R892 VSS.n58 VSS.n57 9.3005
R893 VSS.n228 VSS.n227 9.3005
R894 VSS.n229 VSS.n55 9.3005
R895 VSS.n232 VSS.n231 9.3005
R896 VSS.n230 VSS.n56 9.3005
R897 VSS.n43 VSS.n42 9.3005
R898 VSS.n246 VSS.n245 9.3005
R899 VSS.n247 VSS.n41 9.3005
R900 VSS.n249 VSS.n248 9.3005
R901 VSS.n38 VSS.n37 9.3005
R902 VSS.n257 VSS.n256 9.3005
R903 VSS.n258 VSS.n36 9.3005
R904 VSS.n260 VSS.n259 9.3005
R905 VSS.n32 VSS.n31 9.3005
R906 VSS.n268 VSS.n267 9.3005
R907 VSS.n269 VSS.n30 9.3005
R908 VSS.n271 VSS.n270 9.3005
R909 VSS.n26 VSS.n25 9.3005
R910 VSS.n279 VSS.n278 9.3005
R911 VSS.n280 VSS.n24 9.3005
R912 VSS.n395 VSS.n394 9.3005
R913 VSS.n204 VSS.n203 9.3005
R914 VSS.n205 VSS.n74 9.3005
R915 VSS.n207 VSS.n206 9.3005
R916 VSS.n64 VSS.n63 9.3005
R917 VSS.n220 VSS.n219 9.3005
R918 VSS.n221 VSS.n62 9.3005
R919 VSS.n223 VSS.n222 9.3005
R920 VSS.n49 VSS.n48 9.3005
R921 VSS.n237 VSS.n236 9.3005
R922 VSS.n238 VSS.n47 9.3005
R923 VSS.n240 VSS.n239 9.3005
R924 VSS.n2 VSS.n1 9.3005
R925 VSS.n76 VSS.n75 9.3005
R926 VSS.n419 VSS.n418 9.3005
R927 VSS.n321 VSS.n320 9.05416
R928 VSS.n114 VSS.n113 9.05416
R929 VSS.n320 VSS.n319 1.56148
R930 VSS.n113 VSS.n112 1.56148
R931 VSS.n415 VSS.n0 0.152939
R932 VSS.n415 VSS.n414 0.152939
R933 VSS.n414 VSS.n413 0.152939
R934 VSS.n413 VSS.n7 0.152939
R935 VSS.n409 VSS.n7 0.152939
R936 VSS.n409 VSS.n408 0.152939
R937 VSS.n408 VSS.n407 0.152939
R938 VSS.n407 VSS.n12 0.152939
R939 VSS.n403 VSS.n12 0.152939
R940 VSS.n403 VSS.n402 0.152939
R941 VSS.n402 VSS.n401 0.152939
R942 VSS.n401 VSS.n17 0.152939
R943 VSS.n198 VSS.n197 0.152939
R944 VSS.n198 VSS.n69 0.152939
R945 VSS.n212 VSS.n69 0.152939
R946 VSS.n213 VSS.n212 0.152939
R947 VSS.n214 VSS.n213 0.152939
R948 VSS.n214 VSS.n57 0.152939
R949 VSS.n228 VSS.n57 0.152939
R950 VSS.n229 VSS.n228 0.152939
R951 VSS.n231 VSS.n229 0.152939
R952 VSS.n231 VSS.n230 0.152939
R953 VSS.n230 VSS.n42 0.152939
R954 VSS.n246 VSS.n42 0.152939
R955 VSS.n247 VSS.n246 0.152939
R956 VSS.n248 VSS.n247 0.152939
R957 VSS.n248 VSS.n37 0.152939
R958 VSS.n257 VSS.n37 0.152939
R959 VSS.n258 VSS.n257 0.152939
R960 VSS.n259 VSS.n258 0.152939
R961 VSS.n259 VSS.n31 0.152939
R962 VSS.n268 VSS.n31 0.152939
R963 VSS.n269 VSS.n268 0.152939
R964 VSS.n270 VSS.n269 0.152939
R965 VSS.n270 VSS.n25 0.152939
R966 VSS.n279 VSS.n25 0.152939
R967 VSS.n280 VSS.n279 0.152939
R968 VSS.n394 VSS.n280 0.152939
R969 VSS.n204 VSS.n75 0.152939
R970 VSS.n205 VSS.n204 0.152939
R971 VSS.n206 VSS.n205 0.152939
R972 VSS.n206 VSS.n63 0.152939
R973 VSS.n220 VSS.n63 0.152939
R974 VSS.n221 VSS.n220 0.152939
R975 VSS.n222 VSS.n221 0.152939
R976 VSS.n222 VSS.n48 0.152939
R977 VSS.n237 VSS.n48 0.152939
R978 VSS.n238 VSS.n237 0.152939
R979 VSS.n239 VSS.n238 0.152939
R980 VSS.n239 VSS.n1 0.152939
R981 VSS.n419 VSS.n1 0.13922
R982 VSS VSS.n0 0.0767195
R983 VSS VSS.n419 0.063
R984 VCC.n177 VCC.n13 431.707
R985 VCC.n151 VCC.n28 431.707
R986 VCC.n69 VCC.n57 431.707
R987 VCC.n102 VCC.n59 431.707
R988 VCC.n15 VCC.t4 267.454
R989 VCC.n71 VCC.t0 267.454
R990 VCC.n15 VCC.t6 260.858
R991 VCC.n71 VCC.t3 260.858
R992 VCC.n16 VCC.t7 229.245
R993 VCC.n72 VCC.t2 229.245
R994 VCC.n148 VCC.n28 185
R995 VCC.n144 VCC.n28 185
R996 VCC.n147 VCC.n146 185
R997 VCC.n146 VCC.n145 185
R998 VCC.n31 VCC.n30 185
R999 VCC.n143 VCC.n31 185
R1000 VCC.n141 VCC.n140 185
R1001 VCC.n142 VCC.n141 185
R1002 VCC.n35 VCC.n34 185
R1003 VCC.n34 VCC.n33 185
R1004 VCC.n135 VCC.n134 185
R1005 VCC.n134 VCC.n133 185
R1006 VCC.n38 VCC.n37 185
R1007 VCC.n132 VCC.n38 185
R1008 VCC.n131 VCC.n130 185
R1009 VCC.t8 VCC.n131 185
R1010 VCC.n41 VCC.n40 185
R1011 VCC.n40 VCC.n39 185
R1012 VCC.n126 VCC.n125 185
R1013 VCC.n125 VCC.n124 185
R1014 VCC.n44 VCC.n43 185
R1015 VCC.n45 VCC.n44 185
R1016 VCC.n115 VCC.n114 185
R1017 VCC.n116 VCC.n115 185
R1018 VCC.n54 VCC.n53 185
R1019 VCC.n53 VCC.n52 185
R1020 VCC.n110 VCC.n109 185
R1021 VCC.n109 VCC.n108 185
R1022 VCC.n57 VCC.n56 185
R1023 VCC.n58 VCC.n57 185
R1024 VCC.n60 VCC.n59 185
R1025 VCC.n59 VCC.n58 185
R1026 VCC.n107 VCC.n106 185
R1027 VCC.n108 VCC.n107 185
R1028 VCC.n51 VCC.n50 185
R1029 VCC.n52 VCC.n51 185
R1030 VCC.n118 VCC.n117 185
R1031 VCC.n117 VCC.n116 185
R1032 VCC.n48 VCC.n46 185
R1033 VCC.n46 VCC.n45 185
R1034 VCC.n123 VCC.n122 185
R1035 VCC.n124 VCC.n123 185
R1036 VCC.n47 VCC.n2 185
R1037 VCC.n47 VCC.n39 185
R1038 VCC.n189 VCC.n3 185
R1039 VCC.t8 VCC.n3 185
R1040 VCC.n188 VCC.n4 185
R1041 VCC.n132 VCC.n4 185
R1042 VCC.n187 VCC.n5 185
R1043 VCC.n133 VCC.n5 185
R1044 VCC.n32 VCC.n6 185
R1045 VCC.n33 VCC.n32 185
R1046 VCC.n183 VCC.n8 185
R1047 VCC.n142 VCC.n8 185
R1048 VCC.n182 VCC.n9 185
R1049 VCC.n143 VCC.n9 185
R1050 VCC.n181 VCC.n10 185
R1051 VCC.n145 VCC.n10 185
R1052 VCC.n13 VCC.n11 185
R1053 VCC.n144 VCC.n13 185
R1054 VCC.n151 VCC.n150 185
R1055 VCC.n153 VCC.n26 185
R1056 VCC.n155 VCC.n154 185
R1057 VCC.n156 VCC.n25 185
R1058 VCC.n158 VCC.n157 185
R1059 VCC.n160 VCC.n23 185
R1060 VCC.n162 VCC.n161 185
R1061 VCC.n163 VCC.n22 185
R1062 VCC.n165 VCC.n164 185
R1063 VCC.n167 VCC.n20 185
R1064 VCC.n169 VCC.n168 185
R1065 VCC.n170 VCC.n19 185
R1066 VCC.n172 VCC.n171 185
R1067 VCC.n174 VCC.n18 185
R1068 VCC.n175 VCC.n12 185
R1069 VCC.n178 VCC.n177 185
R1070 VCC.n103 VCC.n102 185
R1071 VCC.n62 VCC.n61 185
R1072 VCC.n99 VCC.n98 185
R1073 VCC.n100 VCC.n99 185
R1074 VCC.n97 VCC.n70 185
R1075 VCC.n96 VCC.n95 185
R1076 VCC.n94 VCC.n93 185
R1077 VCC.n92 VCC.n91 185
R1078 VCC.n90 VCC.n89 185
R1079 VCC.n88 VCC.n87 185
R1080 VCC.n86 VCC.n85 185
R1081 VCC.n84 VCC.n83 185
R1082 VCC.n82 VCC.n81 185
R1083 VCC.n80 VCC.n79 185
R1084 VCC.n78 VCC.n77 185
R1085 VCC.n76 VCC.n75 185
R1086 VCC.n74 VCC.n69 185
R1087 VCC.n100 VCC.n69 185
R1088 VCC.n109 VCC.n57 146.341
R1089 VCC.n109 VCC.n53 146.341
R1090 VCC.n115 VCC.n53 146.341
R1091 VCC.n115 VCC.n44 146.341
R1092 VCC.n125 VCC.n44 146.341
R1093 VCC.n125 VCC.n40 146.341
R1094 VCC.n131 VCC.n40 146.341
R1095 VCC.n131 VCC.n38 146.341
R1096 VCC.n134 VCC.n38 146.341
R1097 VCC.n134 VCC.n34 146.341
R1098 VCC.n141 VCC.n34 146.341
R1099 VCC.n141 VCC.n31 146.341
R1100 VCC.n146 VCC.n31 146.341
R1101 VCC.n146 VCC.n28 146.341
R1102 VCC.n107 VCC.n59 146.341
R1103 VCC.n107 VCC.n51 146.341
R1104 VCC.n117 VCC.n51 146.341
R1105 VCC.n117 VCC.n46 146.341
R1106 VCC.n123 VCC.n46 146.341
R1107 VCC.n123 VCC.n47 146.341
R1108 VCC.n47 VCC.n3 146.341
R1109 VCC.n4 VCC.n3 146.341
R1110 VCC.n5 VCC.n4 146.341
R1111 VCC.n32 VCC.n5 146.341
R1112 VCC.n32 VCC.n8 146.341
R1113 VCC.n9 VCC.n8 146.341
R1114 VCC.n10 VCC.n9 146.341
R1115 VCC.n13 VCC.n10 146.341
R1116 VCC.n100 VCC.n58 126.034
R1117 VCC.n144 VCC.n14 126.034
R1118 VCC.n175 VCC.n174 99.5127
R1119 VCC.n172 VCC.n19 99.5127
R1120 VCC.n168 VCC.n167 99.5127
R1121 VCC.n165 VCC.n22 99.5127
R1122 VCC.n161 VCC.n160 99.5127
R1123 VCC.n158 VCC.n25 99.5127
R1124 VCC.n154 VCC.n153 99.5127
R1125 VCC.n99 VCC.n62 99.5127
R1126 VCC.n99 VCC.n70 99.5127
R1127 VCC.n95 VCC.n94 99.5127
R1128 VCC.n91 VCC.n90 99.5127
R1129 VCC.n87 VCC.n86 99.5127
R1130 VCC.n83 VCC.n82 99.5127
R1131 VCC.n79 VCC.n78 99.5127
R1132 VCC.n75 VCC.n69 99.5127
R1133 VCC.n152 VCC.n14 72.8958
R1134 VCC.n27 VCC.n14 72.8958
R1135 VCC.n159 VCC.n14 72.8958
R1136 VCC.n24 VCC.n14 72.8958
R1137 VCC.n166 VCC.n14 72.8958
R1138 VCC.n21 VCC.n14 72.8958
R1139 VCC.n173 VCC.n14 72.8958
R1140 VCC.n176 VCC.n14 72.8958
R1141 VCC.n101 VCC.n100 72.8958
R1142 VCC.n100 VCC.n63 72.8958
R1143 VCC.n100 VCC.n64 72.8958
R1144 VCC.n100 VCC.n65 72.8958
R1145 VCC.n100 VCC.n66 72.8958
R1146 VCC.n100 VCC.n67 72.8958
R1147 VCC.n100 VCC.n68 72.8958
R1148 VCC.n108 VCC.n58 63.3338
R1149 VCC.n116 VCC.n52 63.3338
R1150 VCC.n116 VCC.n45 63.3338
R1151 VCC.n124 VCC.n45 63.3338
R1152 VCC.n124 VCC.n39 63.3338
R1153 VCC.t8 VCC.n39 63.3338
R1154 VCC.n132 VCC.t8 63.3338
R1155 VCC.n133 VCC.n132 63.3338
R1156 VCC.n133 VCC.n33 63.3338
R1157 VCC.n142 VCC.n33 63.3338
R1158 VCC.n143 VCC.n142 63.3338
R1159 VCC.n145 VCC.n144 63.3338
R1160 VCC.n176 VCC.n175 39.2114
R1161 VCC.n173 VCC.n172 39.2114
R1162 VCC.n168 VCC.n21 39.2114
R1163 VCC.n166 VCC.n165 39.2114
R1164 VCC.n161 VCC.n24 39.2114
R1165 VCC.n159 VCC.n158 39.2114
R1166 VCC.n154 VCC.n27 39.2114
R1167 VCC.n152 VCC.n151 39.2114
R1168 VCC.n102 VCC.n101 39.2114
R1169 VCC.n70 VCC.n63 39.2114
R1170 VCC.n94 VCC.n64 39.2114
R1171 VCC.n90 VCC.n65 39.2114
R1172 VCC.n86 VCC.n66 39.2114
R1173 VCC.n82 VCC.n67 39.2114
R1174 VCC.n78 VCC.n68 39.2114
R1175 VCC.n153 VCC.n152 39.2114
R1176 VCC.n27 VCC.n25 39.2114
R1177 VCC.n160 VCC.n159 39.2114
R1178 VCC.n24 VCC.n22 39.2114
R1179 VCC.n167 VCC.n166 39.2114
R1180 VCC.n21 VCC.n19 39.2114
R1181 VCC.n174 VCC.n173 39.2114
R1182 VCC.n177 VCC.n176 39.2114
R1183 VCC.n101 VCC.n62 39.2114
R1184 VCC.n95 VCC.n63 39.2114
R1185 VCC.n91 VCC.n64 39.2114
R1186 VCC.n87 VCC.n65 39.2114
R1187 VCC.n83 VCC.n66 39.2114
R1188 VCC.n79 VCC.n67 39.2114
R1189 VCC.n75 VCC.n68 39.2114
R1190 VCC.n108 VCC.t1 35.4672
R1191 VCC.n145 VCC.t5 35.4672
R1192 VCC.n16 VCC.n15 31.6126
R1193 VCC.n72 VCC.n71 31.6126
R1194 VCC.n179 VCC.n178 30.9892
R1195 VCC.n150 VCC.n149 30.9892
R1196 VCC.n104 VCC.n103 30.9892
R1197 VCC.n74 VCC.n55 30.9892
R1198 VCC.n17 VCC.n16 29.2853
R1199 VCC.n73 VCC.n72 29.2853
R1200 VCC.t1 VCC.n52 27.8672
R1201 VCC.t5 VCC.n143 27.8672
R1202 VCC.n110 VCC.n56 19.3944
R1203 VCC.n110 VCC.n54 19.3944
R1204 VCC.n114 VCC.n54 19.3944
R1205 VCC.n114 VCC.n43 19.3944
R1206 VCC.n126 VCC.n43 19.3944
R1207 VCC.n126 VCC.n41 19.3944
R1208 VCC.n130 VCC.n41 19.3944
R1209 VCC.n130 VCC.n37 19.3944
R1210 VCC.n135 VCC.n37 19.3944
R1211 VCC.n135 VCC.n35 19.3944
R1212 VCC.n140 VCC.n35 19.3944
R1213 VCC.n140 VCC.n30 19.3944
R1214 VCC.n147 VCC.n30 19.3944
R1215 VCC.n148 VCC.n147 19.3944
R1216 VCC.n106 VCC.n60 19.3944
R1217 VCC.n106 VCC.n50 19.3944
R1218 VCC.n118 VCC.n50 19.3944
R1219 VCC.n118 VCC.n48 19.3944
R1220 VCC.n122 VCC.n48 19.3944
R1221 VCC.n122 VCC.n2 19.3944
R1222 VCC.n189 VCC.n2 19.3944
R1223 VCC.n189 VCC.n188 19.3944
R1224 VCC.n188 VCC.n187 19.3944
R1225 VCC.n187 VCC.n6 19.3944
R1226 VCC.n183 VCC.n6 19.3944
R1227 VCC.n183 VCC.n182 19.3944
R1228 VCC.n182 VCC.n181 19.3944
R1229 VCC.n181 VCC.n11 19.3944
R1230 VCC.n178 VCC.n12 10.6151
R1231 VCC.n171 VCC.n18 10.6151
R1232 VCC.n171 VCC.n170 10.6151
R1233 VCC.n170 VCC.n169 10.6151
R1234 VCC.n169 VCC.n20 10.6151
R1235 VCC.n164 VCC.n20 10.6151
R1236 VCC.n164 VCC.n163 10.6151
R1237 VCC.n163 VCC.n162 10.6151
R1238 VCC.n162 VCC.n23 10.6151
R1239 VCC.n157 VCC.n23 10.6151
R1240 VCC.n157 VCC.n156 10.6151
R1241 VCC.n156 VCC.n155 10.6151
R1242 VCC.n155 VCC.n26 10.6151
R1243 VCC.n150 VCC.n26 10.6151
R1244 VCC.n103 VCC.n61 10.6151
R1245 VCC.n98 VCC.n97 10.6151
R1246 VCC.n97 VCC.n96 10.6151
R1247 VCC.n96 VCC.n93 10.6151
R1248 VCC.n93 VCC.n92 10.6151
R1249 VCC.n92 VCC.n89 10.6151
R1250 VCC.n89 VCC.n88 10.6151
R1251 VCC.n88 VCC.n85 10.6151
R1252 VCC.n85 VCC.n84 10.6151
R1253 VCC.n84 VCC.n81 10.6151
R1254 VCC.n81 VCC.n80 10.6151
R1255 VCC.n80 VCC.n77 10.6151
R1256 VCC.n77 VCC.n76 10.6151
R1257 VCC.n76 VCC.n74 10.6151
R1258 VCC.n188 VCC.n0 9.3005
R1259 VCC.n187 VCC.n186 9.3005
R1260 VCC.n185 VCC.n6 9.3005
R1261 VCC.n184 VCC.n183 9.3005
R1262 VCC.n182 VCC.n7 9.3005
R1263 VCC.n181 VCC.n180 9.3005
R1264 VCC.n179 VCC.n11 9.3005
R1265 VCC.n111 VCC.n110 9.3005
R1266 VCC.n112 VCC.n54 9.3005
R1267 VCC.n114 VCC.n113 9.3005
R1268 VCC.n43 VCC.n42 9.3005
R1269 VCC.n127 VCC.n126 9.3005
R1270 VCC.n128 VCC.n41 9.3005
R1271 VCC.n130 VCC.n129 9.3005
R1272 VCC.n37 VCC.n36 9.3005
R1273 VCC.n136 VCC.n135 9.3005
R1274 VCC.n137 VCC.n35 9.3005
R1275 VCC.n140 VCC.n139 9.3005
R1276 VCC.n138 VCC.n30 9.3005
R1277 VCC.n147 VCC.n29 9.3005
R1278 VCC.n149 VCC.n148 9.3005
R1279 VCC.n56 VCC.n55 9.3005
R1280 VCC.n104 VCC.n60 9.3005
R1281 VCC.n106 VCC.n105 9.3005
R1282 VCC.n50 VCC.n49 9.3005
R1283 VCC.n119 VCC.n118 9.3005
R1284 VCC.n120 VCC.n48 9.3005
R1285 VCC.n122 VCC.n121 9.3005
R1286 VCC.n2 VCC.n1 9.3005
R1287 VCC.n190 VCC.n189 9.3005
R1288 VCC.n17 VCC.n12 5.30782
R1289 VCC.n18 VCC.n17 5.30782
R1290 VCC.n73 VCC.n61 5.30782
R1291 VCC.n98 VCC.n73 5.30782
R1292 VCC.n186 VCC.n0 0.152939
R1293 VCC.n186 VCC.n185 0.152939
R1294 VCC.n185 VCC.n184 0.152939
R1295 VCC.n184 VCC.n7 0.152939
R1296 VCC.n180 VCC.n7 0.152939
R1297 VCC.n180 VCC.n179 0.152939
R1298 VCC.n111 VCC.n55 0.152939
R1299 VCC.n112 VCC.n111 0.152939
R1300 VCC.n113 VCC.n112 0.152939
R1301 VCC.n113 VCC.n42 0.152939
R1302 VCC.n127 VCC.n42 0.152939
R1303 VCC.n128 VCC.n127 0.152939
R1304 VCC.n129 VCC.n128 0.152939
R1305 VCC.n129 VCC.n36 0.152939
R1306 VCC.n136 VCC.n36 0.152939
R1307 VCC.n137 VCC.n136 0.152939
R1308 VCC.n139 VCC.n137 0.152939
R1309 VCC.n139 VCC.n138 0.152939
R1310 VCC.n138 VCC.n29 0.152939
R1311 VCC.n149 VCC.n29 0.152939
R1312 VCC.n105 VCC.n104 0.152939
R1313 VCC.n105 VCC.n49 0.152939
R1314 VCC.n119 VCC.n49 0.152939
R1315 VCC.n120 VCC.n119 0.152939
R1316 VCC.n121 VCC.n120 0.152939
R1317 VCC.n121 VCC.n1 0.152939
R1318 VCC.n190 VCC.n1 0.13922
R1319 VCC VCC.n0 0.0767195
R1320 VCC VCC.n190 0.063
R1321 VGP VGP.t0 174.048
C0 VCC VIN 0.718344f
C1 VCC VGN 0.015036f
C2 VIN VOUT 1.27059f
C3 VGP VIN 0.305185f
C4 VGN VOUT 1.08508f
C5 VGP VGN 0.0052f
C6 VGN VIN 1.23266f
C7 VCC VOUT 0.918948f
C8 VGP VCC 0.664026f
C9 VGP VOUT 0.240022f
C10 VGN VSS 1.71021f
C11 VOUT VSS 1.87415f
C12 VIN VSS 1.64173f
C13 VGP VSS 0.179333f
C14 VCC VSS 10.5468f
.ends

