* NGSPICE file created from diff_pair_sample_1466.ext - technology: sky130A

.subckt diff_pair_sample_1466 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2230_n2590# sky130_fd_pr__pfet_01v8 ad=3.1629 pd=17 as=0 ps=0 w=8.11 l=2.82
X1 B.t8 B.t6 B.t7 w_n2230_n2590# sky130_fd_pr__pfet_01v8 ad=3.1629 pd=17 as=0 ps=0 w=8.11 l=2.82
X2 VDD1.t1 VP.t0 VTAIL.t3 w_n2230_n2590# sky130_fd_pr__pfet_01v8 ad=3.1629 pd=17 as=3.1629 ps=17 w=8.11 l=2.82
X3 VDD2.t1 VN.t0 VTAIL.t1 w_n2230_n2590# sky130_fd_pr__pfet_01v8 ad=3.1629 pd=17 as=3.1629 ps=17 w=8.11 l=2.82
X4 B.t5 B.t3 B.t4 w_n2230_n2590# sky130_fd_pr__pfet_01v8 ad=3.1629 pd=17 as=0 ps=0 w=8.11 l=2.82
X5 VDD2.t0 VN.t1 VTAIL.t0 w_n2230_n2590# sky130_fd_pr__pfet_01v8 ad=3.1629 pd=17 as=3.1629 ps=17 w=8.11 l=2.82
X6 B.t2 B.t0 B.t1 w_n2230_n2590# sky130_fd_pr__pfet_01v8 ad=3.1629 pd=17 as=0 ps=0 w=8.11 l=2.82
X7 VDD1.t0 VP.t1 VTAIL.t2 w_n2230_n2590# sky130_fd_pr__pfet_01v8 ad=3.1629 pd=17 as=3.1629 ps=17 w=8.11 l=2.82
R0 B.n277 B.n276 585
R1 B.n275 B.n82 585
R2 B.n274 B.n273 585
R3 B.n272 B.n83 585
R4 B.n271 B.n270 585
R5 B.n269 B.n84 585
R6 B.n268 B.n267 585
R7 B.n266 B.n85 585
R8 B.n265 B.n264 585
R9 B.n263 B.n86 585
R10 B.n262 B.n261 585
R11 B.n260 B.n87 585
R12 B.n259 B.n258 585
R13 B.n257 B.n88 585
R14 B.n256 B.n255 585
R15 B.n254 B.n89 585
R16 B.n253 B.n252 585
R17 B.n251 B.n90 585
R18 B.n250 B.n249 585
R19 B.n248 B.n91 585
R20 B.n247 B.n246 585
R21 B.n245 B.n92 585
R22 B.n244 B.n243 585
R23 B.n242 B.n93 585
R24 B.n241 B.n240 585
R25 B.n239 B.n94 585
R26 B.n238 B.n237 585
R27 B.n236 B.n95 585
R28 B.n235 B.n234 585
R29 B.n233 B.n96 585
R30 B.n232 B.n231 585
R31 B.n227 B.n97 585
R32 B.n226 B.n225 585
R33 B.n224 B.n98 585
R34 B.n223 B.n222 585
R35 B.n221 B.n99 585
R36 B.n220 B.n219 585
R37 B.n218 B.n100 585
R38 B.n217 B.n216 585
R39 B.n215 B.n101 585
R40 B.n213 B.n212 585
R41 B.n211 B.n104 585
R42 B.n210 B.n209 585
R43 B.n208 B.n105 585
R44 B.n207 B.n206 585
R45 B.n205 B.n106 585
R46 B.n204 B.n203 585
R47 B.n202 B.n107 585
R48 B.n201 B.n200 585
R49 B.n199 B.n108 585
R50 B.n198 B.n197 585
R51 B.n196 B.n109 585
R52 B.n195 B.n194 585
R53 B.n193 B.n110 585
R54 B.n192 B.n191 585
R55 B.n190 B.n111 585
R56 B.n189 B.n188 585
R57 B.n187 B.n112 585
R58 B.n186 B.n185 585
R59 B.n184 B.n113 585
R60 B.n183 B.n182 585
R61 B.n181 B.n114 585
R62 B.n180 B.n179 585
R63 B.n178 B.n115 585
R64 B.n177 B.n176 585
R65 B.n175 B.n116 585
R66 B.n174 B.n173 585
R67 B.n172 B.n117 585
R68 B.n171 B.n170 585
R69 B.n169 B.n118 585
R70 B.n278 B.n81 585
R71 B.n280 B.n279 585
R72 B.n281 B.n80 585
R73 B.n283 B.n282 585
R74 B.n284 B.n79 585
R75 B.n286 B.n285 585
R76 B.n287 B.n78 585
R77 B.n289 B.n288 585
R78 B.n290 B.n77 585
R79 B.n292 B.n291 585
R80 B.n293 B.n76 585
R81 B.n295 B.n294 585
R82 B.n296 B.n75 585
R83 B.n298 B.n297 585
R84 B.n299 B.n74 585
R85 B.n301 B.n300 585
R86 B.n302 B.n73 585
R87 B.n304 B.n303 585
R88 B.n305 B.n72 585
R89 B.n307 B.n306 585
R90 B.n308 B.n71 585
R91 B.n310 B.n309 585
R92 B.n311 B.n70 585
R93 B.n313 B.n312 585
R94 B.n314 B.n69 585
R95 B.n316 B.n315 585
R96 B.n317 B.n68 585
R97 B.n319 B.n318 585
R98 B.n320 B.n67 585
R99 B.n322 B.n321 585
R100 B.n323 B.n66 585
R101 B.n325 B.n324 585
R102 B.n326 B.n65 585
R103 B.n328 B.n327 585
R104 B.n329 B.n64 585
R105 B.n331 B.n330 585
R106 B.n332 B.n63 585
R107 B.n334 B.n333 585
R108 B.n335 B.n62 585
R109 B.n337 B.n336 585
R110 B.n338 B.n61 585
R111 B.n340 B.n339 585
R112 B.n341 B.n60 585
R113 B.n343 B.n342 585
R114 B.n344 B.n59 585
R115 B.n346 B.n345 585
R116 B.n347 B.n58 585
R117 B.n349 B.n348 585
R118 B.n350 B.n57 585
R119 B.n352 B.n351 585
R120 B.n353 B.n56 585
R121 B.n355 B.n354 585
R122 B.n356 B.n55 585
R123 B.n358 B.n357 585
R124 B.n464 B.n15 585
R125 B.n463 B.n462 585
R126 B.n461 B.n16 585
R127 B.n460 B.n459 585
R128 B.n458 B.n17 585
R129 B.n457 B.n456 585
R130 B.n455 B.n18 585
R131 B.n454 B.n453 585
R132 B.n452 B.n19 585
R133 B.n451 B.n450 585
R134 B.n449 B.n20 585
R135 B.n448 B.n447 585
R136 B.n446 B.n21 585
R137 B.n445 B.n444 585
R138 B.n443 B.n22 585
R139 B.n442 B.n441 585
R140 B.n440 B.n23 585
R141 B.n439 B.n438 585
R142 B.n437 B.n24 585
R143 B.n436 B.n435 585
R144 B.n434 B.n25 585
R145 B.n433 B.n432 585
R146 B.n431 B.n26 585
R147 B.n430 B.n429 585
R148 B.n428 B.n27 585
R149 B.n427 B.n426 585
R150 B.n425 B.n28 585
R151 B.n424 B.n423 585
R152 B.n422 B.n29 585
R153 B.n421 B.n420 585
R154 B.n419 B.n418 585
R155 B.n417 B.n33 585
R156 B.n416 B.n415 585
R157 B.n414 B.n34 585
R158 B.n413 B.n412 585
R159 B.n411 B.n35 585
R160 B.n410 B.n409 585
R161 B.n408 B.n36 585
R162 B.n407 B.n406 585
R163 B.n405 B.n37 585
R164 B.n403 B.n402 585
R165 B.n401 B.n40 585
R166 B.n400 B.n399 585
R167 B.n398 B.n41 585
R168 B.n397 B.n396 585
R169 B.n395 B.n42 585
R170 B.n394 B.n393 585
R171 B.n392 B.n43 585
R172 B.n391 B.n390 585
R173 B.n389 B.n44 585
R174 B.n388 B.n387 585
R175 B.n386 B.n45 585
R176 B.n385 B.n384 585
R177 B.n383 B.n46 585
R178 B.n382 B.n381 585
R179 B.n380 B.n47 585
R180 B.n379 B.n378 585
R181 B.n377 B.n48 585
R182 B.n376 B.n375 585
R183 B.n374 B.n49 585
R184 B.n373 B.n372 585
R185 B.n371 B.n50 585
R186 B.n370 B.n369 585
R187 B.n368 B.n51 585
R188 B.n367 B.n366 585
R189 B.n365 B.n52 585
R190 B.n364 B.n363 585
R191 B.n362 B.n53 585
R192 B.n361 B.n360 585
R193 B.n359 B.n54 585
R194 B.n466 B.n465 585
R195 B.n467 B.n14 585
R196 B.n469 B.n468 585
R197 B.n470 B.n13 585
R198 B.n472 B.n471 585
R199 B.n473 B.n12 585
R200 B.n475 B.n474 585
R201 B.n476 B.n11 585
R202 B.n478 B.n477 585
R203 B.n479 B.n10 585
R204 B.n481 B.n480 585
R205 B.n482 B.n9 585
R206 B.n484 B.n483 585
R207 B.n485 B.n8 585
R208 B.n487 B.n486 585
R209 B.n488 B.n7 585
R210 B.n490 B.n489 585
R211 B.n491 B.n6 585
R212 B.n493 B.n492 585
R213 B.n494 B.n5 585
R214 B.n496 B.n495 585
R215 B.n497 B.n4 585
R216 B.n499 B.n498 585
R217 B.n500 B.n3 585
R218 B.n502 B.n501 585
R219 B.n503 B.n0 585
R220 B.n2 B.n1 585
R221 B.n132 B.n131 585
R222 B.n133 B.n130 585
R223 B.n135 B.n134 585
R224 B.n136 B.n129 585
R225 B.n138 B.n137 585
R226 B.n139 B.n128 585
R227 B.n141 B.n140 585
R228 B.n142 B.n127 585
R229 B.n144 B.n143 585
R230 B.n145 B.n126 585
R231 B.n147 B.n146 585
R232 B.n148 B.n125 585
R233 B.n150 B.n149 585
R234 B.n151 B.n124 585
R235 B.n153 B.n152 585
R236 B.n154 B.n123 585
R237 B.n156 B.n155 585
R238 B.n157 B.n122 585
R239 B.n159 B.n158 585
R240 B.n160 B.n121 585
R241 B.n162 B.n161 585
R242 B.n163 B.n120 585
R243 B.n165 B.n164 585
R244 B.n166 B.n119 585
R245 B.n168 B.n167 585
R246 B.n169 B.n168 516.524
R247 B.n276 B.n81 516.524
R248 B.n359 B.n358 516.524
R249 B.n466 B.n15 516.524
R250 B.n228 B.t10 366.914
R251 B.n38 B.t2 366.914
R252 B.n102 B.t7 366.914
R253 B.n30 B.t5 366.914
R254 B.n229 B.t11 305.824
R255 B.n39 B.t1 305.824
R256 B.n103 B.t8 305.824
R257 B.n31 B.t4 305.824
R258 B.n102 B.t6 277.666
R259 B.n228 B.t9 277.666
R260 B.n38 B.t0 277.666
R261 B.n30 B.t3 277.666
R262 B.n505 B.n504 256.663
R263 B.n504 B.n503 235.042
R264 B.n504 B.n2 235.042
R265 B.n170 B.n169 163.367
R266 B.n170 B.n117 163.367
R267 B.n174 B.n117 163.367
R268 B.n175 B.n174 163.367
R269 B.n176 B.n175 163.367
R270 B.n176 B.n115 163.367
R271 B.n180 B.n115 163.367
R272 B.n181 B.n180 163.367
R273 B.n182 B.n181 163.367
R274 B.n182 B.n113 163.367
R275 B.n186 B.n113 163.367
R276 B.n187 B.n186 163.367
R277 B.n188 B.n187 163.367
R278 B.n188 B.n111 163.367
R279 B.n192 B.n111 163.367
R280 B.n193 B.n192 163.367
R281 B.n194 B.n193 163.367
R282 B.n194 B.n109 163.367
R283 B.n198 B.n109 163.367
R284 B.n199 B.n198 163.367
R285 B.n200 B.n199 163.367
R286 B.n200 B.n107 163.367
R287 B.n204 B.n107 163.367
R288 B.n205 B.n204 163.367
R289 B.n206 B.n205 163.367
R290 B.n206 B.n105 163.367
R291 B.n210 B.n105 163.367
R292 B.n211 B.n210 163.367
R293 B.n212 B.n211 163.367
R294 B.n212 B.n101 163.367
R295 B.n217 B.n101 163.367
R296 B.n218 B.n217 163.367
R297 B.n219 B.n218 163.367
R298 B.n219 B.n99 163.367
R299 B.n223 B.n99 163.367
R300 B.n224 B.n223 163.367
R301 B.n225 B.n224 163.367
R302 B.n225 B.n97 163.367
R303 B.n232 B.n97 163.367
R304 B.n233 B.n232 163.367
R305 B.n234 B.n233 163.367
R306 B.n234 B.n95 163.367
R307 B.n238 B.n95 163.367
R308 B.n239 B.n238 163.367
R309 B.n240 B.n239 163.367
R310 B.n240 B.n93 163.367
R311 B.n244 B.n93 163.367
R312 B.n245 B.n244 163.367
R313 B.n246 B.n245 163.367
R314 B.n246 B.n91 163.367
R315 B.n250 B.n91 163.367
R316 B.n251 B.n250 163.367
R317 B.n252 B.n251 163.367
R318 B.n252 B.n89 163.367
R319 B.n256 B.n89 163.367
R320 B.n257 B.n256 163.367
R321 B.n258 B.n257 163.367
R322 B.n258 B.n87 163.367
R323 B.n262 B.n87 163.367
R324 B.n263 B.n262 163.367
R325 B.n264 B.n263 163.367
R326 B.n264 B.n85 163.367
R327 B.n268 B.n85 163.367
R328 B.n269 B.n268 163.367
R329 B.n270 B.n269 163.367
R330 B.n270 B.n83 163.367
R331 B.n274 B.n83 163.367
R332 B.n275 B.n274 163.367
R333 B.n276 B.n275 163.367
R334 B.n358 B.n55 163.367
R335 B.n354 B.n55 163.367
R336 B.n354 B.n353 163.367
R337 B.n353 B.n352 163.367
R338 B.n352 B.n57 163.367
R339 B.n348 B.n57 163.367
R340 B.n348 B.n347 163.367
R341 B.n347 B.n346 163.367
R342 B.n346 B.n59 163.367
R343 B.n342 B.n59 163.367
R344 B.n342 B.n341 163.367
R345 B.n341 B.n340 163.367
R346 B.n340 B.n61 163.367
R347 B.n336 B.n61 163.367
R348 B.n336 B.n335 163.367
R349 B.n335 B.n334 163.367
R350 B.n334 B.n63 163.367
R351 B.n330 B.n63 163.367
R352 B.n330 B.n329 163.367
R353 B.n329 B.n328 163.367
R354 B.n328 B.n65 163.367
R355 B.n324 B.n65 163.367
R356 B.n324 B.n323 163.367
R357 B.n323 B.n322 163.367
R358 B.n322 B.n67 163.367
R359 B.n318 B.n67 163.367
R360 B.n318 B.n317 163.367
R361 B.n317 B.n316 163.367
R362 B.n316 B.n69 163.367
R363 B.n312 B.n69 163.367
R364 B.n312 B.n311 163.367
R365 B.n311 B.n310 163.367
R366 B.n310 B.n71 163.367
R367 B.n306 B.n71 163.367
R368 B.n306 B.n305 163.367
R369 B.n305 B.n304 163.367
R370 B.n304 B.n73 163.367
R371 B.n300 B.n73 163.367
R372 B.n300 B.n299 163.367
R373 B.n299 B.n298 163.367
R374 B.n298 B.n75 163.367
R375 B.n294 B.n75 163.367
R376 B.n294 B.n293 163.367
R377 B.n293 B.n292 163.367
R378 B.n292 B.n77 163.367
R379 B.n288 B.n77 163.367
R380 B.n288 B.n287 163.367
R381 B.n287 B.n286 163.367
R382 B.n286 B.n79 163.367
R383 B.n282 B.n79 163.367
R384 B.n282 B.n281 163.367
R385 B.n281 B.n280 163.367
R386 B.n280 B.n81 163.367
R387 B.n462 B.n15 163.367
R388 B.n462 B.n461 163.367
R389 B.n461 B.n460 163.367
R390 B.n460 B.n17 163.367
R391 B.n456 B.n17 163.367
R392 B.n456 B.n455 163.367
R393 B.n455 B.n454 163.367
R394 B.n454 B.n19 163.367
R395 B.n450 B.n19 163.367
R396 B.n450 B.n449 163.367
R397 B.n449 B.n448 163.367
R398 B.n448 B.n21 163.367
R399 B.n444 B.n21 163.367
R400 B.n444 B.n443 163.367
R401 B.n443 B.n442 163.367
R402 B.n442 B.n23 163.367
R403 B.n438 B.n23 163.367
R404 B.n438 B.n437 163.367
R405 B.n437 B.n436 163.367
R406 B.n436 B.n25 163.367
R407 B.n432 B.n25 163.367
R408 B.n432 B.n431 163.367
R409 B.n431 B.n430 163.367
R410 B.n430 B.n27 163.367
R411 B.n426 B.n27 163.367
R412 B.n426 B.n425 163.367
R413 B.n425 B.n424 163.367
R414 B.n424 B.n29 163.367
R415 B.n420 B.n29 163.367
R416 B.n420 B.n419 163.367
R417 B.n419 B.n33 163.367
R418 B.n415 B.n33 163.367
R419 B.n415 B.n414 163.367
R420 B.n414 B.n413 163.367
R421 B.n413 B.n35 163.367
R422 B.n409 B.n35 163.367
R423 B.n409 B.n408 163.367
R424 B.n408 B.n407 163.367
R425 B.n407 B.n37 163.367
R426 B.n402 B.n37 163.367
R427 B.n402 B.n401 163.367
R428 B.n401 B.n400 163.367
R429 B.n400 B.n41 163.367
R430 B.n396 B.n41 163.367
R431 B.n396 B.n395 163.367
R432 B.n395 B.n394 163.367
R433 B.n394 B.n43 163.367
R434 B.n390 B.n43 163.367
R435 B.n390 B.n389 163.367
R436 B.n389 B.n388 163.367
R437 B.n388 B.n45 163.367
R438 B.n384 B.n45 163.367
R439 B.n384 B.n383 163.367
R440 B.n383 B.n382 163.367
R441 B.n382 B.n47 163.367
R442 B.n378 B.n47 163.367
R443 B.n378 B.n377 163.367
R444 B.n377 B.n376 163.367
R445 B.n376 B.n49 163.367
R446 B.n372 B.n49 163.367
R447 B.n372 B.n371 163.367
R448 B.n371 B.n370 163.367
R449 B.n370 B.n51 163.367
R450 B.n366 B.n51 163.367
R451 B.n366 B.n365 163.367
R452 B.n365 B.n364 163.367
R453 B.n364 B.n53 163.367
R454 B.n360 B.n53 163.367
R455 B.n360 B.n359 163.367
R456 B.n467 B.n466 163.367
R457 B.n468 B.n467 163.367
R458 B.n468 B.n13 163.367
R459 B.n472 B.n13 163.367
R460 B.n473 B.n472 163.367
R461 B.n474 B.n473 163.367
R462 B.n474 B.n11 163.367
R463 B.n478 B.n11 163.367
R464 B.n479 B.n478 163.367
R465 B.n480 B.n479 163.367
R466 B.n480 B.n9 163.367
R467 B.n484 B.n9 163.367
R468 B.n485 B.n484 163.367
R469 B.n486 B.n485 163.367
R470 B.n486 B.n7 163.367
R471 B.n490 B.n7 163.367
R472 B.n491 B.n490 163.367
R473 B.n492 B.n491 163.367
R474 B.n492 B.n5 163.367
R475 B.n496 B.n5 163.367
R476 B.n497 B.n496 163.367
R477 B.n498 B.n497 163.367
R478 B.n498 B.n3 163.367
R479 B.n502 B.n3 163.367
R480 B.n503 B.n502 163.367
R481 B.n132 B.n2 163.367
R482 B.n133 B.n132 163.367
R483 B.n134 B.n133 163.367
R484 B.n134 B.n129 163.367
R485 B.n138 B.n129 163.367
R486 B.n139 B.n138 163.367
R487 B.n140 B.n139 163.367
R488 B.n140 B.n127 163.367
R489 B.n144 B.n127 163.367
R490 B.n145 B.n144 163.367
R491 B.n146 B.n145 163.367
R492 B.n146 B.n125 163.367
R493 B.n150 B.n125 163.367
R494 B.n151 B.n150 163.367
R495 B.n152 B.n151 163.367
R496 B.n152 B.n123 163.367
R497 B.n156 B.n123 163.367
R498 B.n157 B.n156 163.367
R499 B.n158 B.n157 163.367
R500 B.n158 B.n121 163.367
R501 B.n162 B.n121 163.367
R502 B.n163 B.n162 163.367
R503 B.n164 B.n163 163.367
R504 B.n164 B.n119 163.367
R505 B.n168 B.n119 163.367
R506 B.n103 B.n102 61.0914
R507 B.n229 B.n228 61.0914
R508 B.n39 B.n38 61.0914
R509 B.n31 B.n30 61.0914
R510 B.n214 B.n103 59.5399
R511 B.n230 B.n229 59.5399
R512 B.n404 B.n39 59.5399
R513 B.n32 B.n31 59.5399
R514 B.n465 B.n464 33.5615
R515 B.n357 B.n54 33.5615
R516 B.n278 B.n277 33.5615
R517 B.n167 B.n118 33.5615
R518 B B.n505 18.0485
R519 B.n465 B.n14 10.6151
R520 B.n469 B.n14 10.6151
R521 B.n470 B.n469 10.6151
R522 B.n471 B.n470 10.6151
R523 B.n471 B.n12 10.6151
R524 B.n475 B.n12 10.6151
R525 B.n476 B.n475 10.6151
R526 B.n477 B.n476 10.6151
R527 B.n477 B.n10 10.6151
R528 B.n481 B.n10 10.6151
R529 B.n482 B.n481 10.6151
R530 B.n483 B.n482 10.6151
R531 B.n483 B.n8 10.6151
R532 B.n487 B.n8 10.6151
R533 B.n488 B.n487 10.6151
R534 B.n489 B.n488 10.6151
R535 B.n489 B.n6 10.6151
R536 B.n493 B.n6 10.6151
R537 B.n494 B.n493 10.6151
R538 B.n495 B.n494 10.6151
R539 B.n495 B.n4 10.6151
R540 B.n499 B.n4 10.6151
R541 B.n500 B.n499 10.6151
R542 B.n501 B.n500 10.6151
R543 B.n501 B.n0 10.6151
R544 B.n464 B.n463 10.6151
R545 B.n463 B.n16 10.6151
R546 B.n459 B.n16 10.6151
R547 B.n459 B.n458 10.6151
R548 B.n458 B.n457 10.6151
R549 B.n457 B.n18 10.6151
R550 B.n453 B.n18 10.6151
R551 B.n453 B.n452 10.6151
R552 B.n452 B.n451 10.6151
R553 B.n451 B.n20 10.6151
R554 B.n447 B.n20 10.6151
R555 B.n447 B.n446 10.6151
R556 B.n446 B.n445 10.6151
R557 B.n445 B.n22 10.6151
R558 B.n441 B.n22 10.6151
R559 B.n441 B.n440 10.6151
R560 B.n440 B.n439 10.6151
R561 B.n439 B.n24 10.6151
R562 B.n435 B.n24 10.6151
R563 B.n435 B.n434 10.6151
R564 B.n434 B.n433 10.6151
R565 B.n433 B.n26 10.6151
R566 B.n429 B.n26 10.6151
R567 B.n429 B.n428 10.6151
R568 B.n428 B.n427 10.6151
R569 B.n427 B.n28 10.6151
R570 B.n423 B.n28 10.6151
R571 B.n423 B.n422 10.6151
R572 B.n422 B.n421 10.6151
R573 B.n418 B.n417 10.6151
R574 B.n417 B.n416 10.6151
R575 B.n416 B.n34 10.6151
R576 B.n412 B.n34 10.6151
R577 B.n412 B.n411 10.6151
R578 B.n411 B.n410 10.6151
R579 B.n410 B.n36 10.6151
R580 B.n406 B.n36 10.6151
R581 B.n406 B.n405 10.6151
R582 B.n403 B.n40 10.6151
R583 B.n399 B.n40 10.6151
R584 B.n399 B.n398 10.6151
R585 B.n398 B.n397 10.6151
R586 B.n397 B.n42 10.6151
R587 B.n393 B.n42 10.6151
R588 B.n393 B.n392 10.6151
R589 B.n392 B.n391 10.6151
R590 B.n391 B.n44 10.6151
R591 B.n387 B.n44 10.6151
R592 B.n387 B.n386 10.6151
R593 B.n386 B.n385 10.6151
R594 B.n385 B.n46 10.6151
R595 B.n381 B.n46 10.6151
R596 B.n381 B.n380 10.6151
R597 B.n380 B.n379 10.6151
R598 B.n379 B.n48 10.6151
R599 B.n375 B.n48 10.6151
R600 B.n375 B.n374 10.6151
R601 B.n374 B.n373 10.6151
R602 B.n373 B.n50 10.6151
R603 B.n369 B.n50 10.6151
R604 B.n369 B.n368 10.6151
R605 B.n368 B.n367 10.6151
R606 B.n367 B.n52 10.6151
R607 B.n363 B.n52 10.6151
R608 B.n363 B.n362 10.6151
R609 B.n362 B.n361 10.6151
R610 B.n361 B.n54 10.6151
R611 B.n357 B.n356 10.6151
R612 B.n356 B.n355 10.6151
R613 B.n355 B.n56 10.6151
R614 B.n351 B.n56 10.6151
R615 B.n351 B.n350 10.6151
R616 B.n350 B.n349 10.6151
R617 B.n349 B.n58 10.6151
R618 B.n345 B.n58 10.6151
R619 B.n345 B.n344 10.6151
R620 B.n344 B.n343 10.6151
R621 B.n343 B.n60 10.6151
R622 B.n339 B.n60 10.6151
R623 B.n339 B.n338 10.6151
R624 B.n338 B.n337 10.6151
R625 B.n337 B.n62 10.6151
R626 B.n333 B.n62 10.6151
R627 B.n333 B.n332 10.6151
R628 B.n332 B.n331 10.6151
R629 B.n331 B.n64 10.6151
R630 B.n327 B.n64 10.6151
R631 B.n327 B.n326 10.6151
R632 B.n326 B.n325 10.6151
R633 B.n325 B.n66 10.6151
R634 B.n321 B.n66 10.6151
R635 B.n321 B.n320 10.6151
R636 B.n320 B.n319 10.6151
R637 B.n319 B.n68 10.6151
R638 B.n315 B.n68 10.6151
R639 B.n315 B.n314 10.6151
R640 B.n314 B.n313 10.6151
R641 B.n313 B.n70 10.6151
R642 B.n309 B.n70 10.6151
R643 B.n309 B.n308 10.6151
R644 B.n308 B.n307 10.6151
R645 B.n307 B.n72 10.6151
R646 B.n303 B.n72 10.6151
R647 B.n303 B.n302 10.6151
R648 B.n302 B.n301 10.6151
R649 B.n301 B.n74 10.6151
R650 B.n297 B.n74 10.6151
R651 B.n297 B.n296 10.6151
R652 B.n296 B.n295 10.6151
R653 B.n295 B.n76 10.6151
R654 B.n291 B.n76 10.6151
R655 B.n291 B.n290 10.6151
R656 B.n290 B.n289 10.6151
R657 B.n289 B.n78 10.6151
R658 B.n285 B.n78 10.6151
R659 B.n285 B.n284 10.6151
R660 B.n284 B.n283 10.6151
R661 B.n283 B.n80 10.6151
R662 B.n279 B.n80 10.6151
R663 B.n279 B.n278 10.6151
R664 B.n131 B.n1 10.6151
R665 B.n131 B.n130 10.6151
R666 B.n135 B.n130 10.6151
R667 B.n136 B.n135 10.6151
R668 B.n137 B.n136 10.6151
R669 B.n137 B.n128 10.6151
R670 B.n141 B.n128 10.6151
R671 B.n142 B.n141 10.6151
R672 B.n143 B.n142 10.6151
R673 B.n143 B.n126 10.6151
R674 B.n147 B.n126 10.6151
R675 B.n148 B.n147 10.6151
R676 B.n149 B.n148 10.6151
R677 B.n149 B.n124 10.6151
R678 B.n153 B.n124 10.6151
R679 B.n154 B.n153 10.6151
R680 B.n155 B.n154 10.6151
R681 B.n155 B.n122 10.6151
R682 B.n159 B.n122 10.6151
R683 B.n160 B.n159 10.6151
R684 B.n161 B.n160 10.6151
R685 B.n161 B.n120 10.6151
R686 B.n165 B.n120 10.6151
R687 B.n166 B.n165 10.6151
R688 B.n167 B.n166 10.6151
R689 B.n171 B.n118 10.6151
R690 B.n172 B.n171 10.6151
R691 B.n173 B.n172 10.6151
R692 B.n173 B.n116 10.6151
R693 B.n177 B.n116 10.6151
R694 B.n178 B.n177 10.6151
R695 B.n179 B.n178 10.6151
R696 B.n179 B.n114 10.6151
R697 B.n183 B.n114 10.6151
R698 B.n184 B.n183 10.6151
R699 B.n185 B.n184 10.6151
R700 B.n185 B.n112 10.6151
R701 B.n189 B.n112 10.6151
R702 B.n190 B.n189 10.6151
R703 B.n191 B.n190 10.6151
R704 B.n191 B.n110 10.6151
R705 B.n195 B.n110 10.6151
R706 B.n196 B.n195 10.6151
R707 B.n197 B.n196 10.6151
R708 B.n197 B.n108 10.6151
R709 B.n201 B.n108 10.6151
R710 B.n202 B.n201 10.6151
R711 B.n203 B.n202 10.6151
R712 B.n203 B.n106 10.6151
R713 B.n207 B.n106 10.6151
R714 B.n208 B.n207 10.6151
R715 B.n209 B.n208 10.6151
R716 B.n209 B.n104 10.6151
R717 B.n213 B.n104 10.6151
R718 B.n216 B.n215 10.6151
R719 B.n216 B.n100 10.6151
R720 B.n220 B.n100 10.6151
R721 B.n221 B.n220 10.6151
R722 B.n222 B.n221 10.6151
R723 B.n222 B.n98 10.6151
R724 B.n226 B.n98 10.6151
R725 B.n227 B.n226 10.6151
R726 B.n231 B.n227 10.6151
R727 B.n235 B.n96 10.6151
R728 B.n236 B.n235 10.6151
R729 B.n237 B.n236 10.6151
R730 B.n237 B.n94 10.6151
R731 B.n241 B.n94 10.6151
R732 B.n242 B.n241 10.6151
R733 B.n243 B.n242 10.6151
R734 B.n243 B.n92 10.6151
R735 B.n247 B.n92 10.6151
R736 B.n248 B.n247 10.6151
R737 B.n249 B.n248 10.6151
R738 B.n249 B.n90 10.6151
R739 B.n253 B.n90 10.6151
R740 B.n254 B.n253 10.6151
R741 B.n255 B.n254 10.6151
R742 B.n255 B.n88 10.6151
R743 B.n259 B.n88 10.6151
R744 B.n260 B.n259 10.6151
R745 B.n261 B.n260 10.6151
R746 B.n261 B.n86 10.6151
R747 B.n265 B.n86 10.6151
R748 B.n266 B.n265 10.6151
R749 B.n267 B.n266 10.6151
R750 B.n267 B.n84 10.6151
R751 B.n271 B.n84 10.6151
R752 B.n272 B.n271 10.6151
R753 B.n273 B.n272 10.6151
R754 B.n273 B.n82 10.6151
R755 B.n277 B.n82 10.6151
R756 B.n421 B.n32 9.36635
R757 B.n404 B.n403 9.36635
R758 B.n214 B.n213 9.36635
R759 B.n230 B.n96 9.36635
R760 B.n505 B.n0 8.11757
R761 B.n505 B.n1 8.11757
R762 B.n418 B.n32 1.24928
R763 B.n405 B.n404 1.24928
R764 B.n215 B.n214 1.24928
R765 B.n231 B.n230 1.24928
R766 VP.n0 VP.t0 152.698
R767 VP.n0 VP.t1 110.406
R768 VP VP.n0 0.431811
R769 VTAIL.n170 VTAIL.n132 756.745
R770 VTAIL.n38 VTAIL.n0 756.745
R771 VTAIL.n126 VTAIL.n88 756.745
R772 VTAIL.n82 VTAIL.n44 756.745
R773 VTAIL.n147 VTAIL.n146 585
R774 VTAIL.n144 VTAIL.n143 585
R775 VTAIL.n153 VTAIL.n152 585
R776 VTAIL.n155 VTAIL.n154 585
R777 VTAIL.n140 VTAIL.n139 585
R778 VTAIL.n161 VTAIL.n160 585
R779 VTAIL.n163 VTAIL.n162 585
R780 VTAIL.n136 VTAIL.n135 585
R781 VTAIL.n169 VTAIL.n168 585
R782 VTAIL.n171 VTAIL.n170 585
R783 VTAIL.n15 VTAIL.n14 585
R784 VTAIL.n12 VTAIL.n11 585
R785 VTAIL.n21 VTAIL.n20 585
R786 VTAIL.n23 VTAIL.n22 585
R787 VTAIL.n8 VTAIL.n7 585
R788 VTAIL.n29 VTAIL.n28 585
R789 VTAIL.n31 VTAIL.n30 585
R790 VTAIL.n4 VTAIL.n3 585
R791 VTAIL.n37 VTAIL.n36 585
R792 VTAIL.n39 VTAIL.n38 585
R793 VTAIL.n127 VTAIL.n126 585
R794 VTAIL.n125 VTAIL.n124 585
R795 VTAIL.n92 VTAIL.n91 585
R796 VTAIL.n119 VTAIL.n118 585
R797 VTAIL.n117 VTAIL.n116 585
R798 VTAIL.n96 VTAIL.n95 585
R799 VTAIL.n111 VTAIL.n110 585
R800 VTAIL.n109 VTAIL.n108 585
R801 VTAIL.n100 VTAIL.n99 585
R802 VTAIL.n103 VTAIL.n102 585
R803 VTAIL.n83 VTAIL.n82 585
R804 VTAIL.n81 VTAIL.n80 585
R805 VTAIL.n48 VTAIL.n47 585
R806 VTAIL.n75 VTAIL.n74 585
R807 VTAIL.n73 VTAIL.n72 585
R808 VTAIL.n52 VTAIL.n51 585
R809 VTAIL.n67 VTAIL.n66 585
R810 VTAIL.n65 VTAIL.n64 585
R811 VTAIL.n56 VTAIL.n55 585
R812 VTAIL.n59 VTAIL.n58 585
R813 VTAIL.t0 VTAIL.n145 327.473
R814 VTAIL.t2 VTAIL.n13 327.473
R815 VTAIL.t3 VTAIL.n101 327.473
R816 VTAIL.t1 VTAIL.n57 327.473
R817 VTAIL.n146 VTAIL.n143 171.744
R818 VTAIL.n153 VTAIL.n143 171.744
R819 VTAIL.n154 VTAIL.n153 171.744
R820 VTAIL.n154 VTAIL.n139 171.744
R821 VTAIL.n161 VTAIL.n139 171.744
R822 VTAIL.n162 VTAIL.n161 171.744
R823 VTAIL.n162 VTAIL.n135 171.744
R824 VTAIL.n169 VTAIL.n135 171.744
R825 VTAIL.n170 VTAIL.n169 171.744
R826 VTAIL.n14 VTAIL.n11 171.744
R827 VTAIL.n21 VTAIL.n11 171.744
R828 VTAIL.n22 VTAIL.n21 171.744
R829 VTAIL.n22 VTAIL.n7 171.744
R830 VTAIL.n29 VTAIL.n7 171.744
R831 VTAIL.n30 VTAIL.n29 171.744
R832 VTAIL.n30 VTAIL.n3 171.744
R833 VTAIL.n37 VTAIL.n3 171.744
R834 VTAIL.n38 VTAIL.n37 171.744
R835 VTAIL.n126 VTAIL.n125 171.744
R836 VTAIL.n125 VTAIL.n91 171.744
R837 VTAIL.n118 VTAIL.n91 171.744
R838 VTAIL.n118 VTAIL.n117 171.744
R839 VTAIL.n117 VTAIL.n95 171.744
R840 VTAIL.n110 VTAIL.n95 171.744
R841 VTAIL.n110 VTAIL.n109 171.744
R842 VTAIL.n109 VTAIL.n99 171.744
R843 VTAIL.n102 VTAIL.n99 171.744
R844 VTAIL.n82 VTAIL.n81 171.744
R845 VTAIL.n81 VTAIL.n47 171.744
R846 VTAIL.n74 VTAIL.n47 171.744
R847 VTAIL.n74 VTAIL.n73 171.744
R848 VTAIL.n73 VTAIL.n51 171.744
R849 VTAIL.n66 VTAIL.n51 171.744
R850 VTAIL.n66 VTAIL.n65 171.744
R851 VTAIL.n65 VTAIL.n55 171.744
R852 VTAIL.n58 VTAIL.n55 171.744
R853 VTAIL.n146 VTAIL.t0 85.8723
R854 VTAIL.n14 VTAIL.t2 85.8723
R855 VTAIL.n102 VTAIL.t3 85.8723
R856 VTAIL.n58 VTAIL.t1 85.8723
R857 VTAIL.n175 VTAIL.n174 31.2157
R858 VTAIL.n43 VTAIL.n42 31.2157
R859 VTAIL.n131 VTAIL.n130 31.2157
R860 VTAIL.n87 VTAIL.n86 31.2157
R861 VTAIL.n87 VTAIL.n43 24.7893
R862 VTAIL.n175 VTAIL.n131 22.0738
R863 VTAIL.n147 VTAIL.n145 16.3894
R864 VTAIL.n15 VTAIL.n13 16.3894
R865 VTAIL.n103 VTAIL.n101 16.3894
R866 VTAIL.n59 VTAIL.n57 16.3894
R867 VTAIL.n148 VTAIL.n144 12.8005
R868 VTAIL.n16 VTAIL.n12 12.8005
R869 VTAIL.n104 VTAIL.n100 12.8005
R870 VTAIL.n60 VTAIL.n56 12.8005
R871 VTAIL.n152 VTAIL.n151 12.0247
R872 VTAIL.n20 VTAIL.n19 12.0247
R873 VTAIL.n108 VTAIL.n107 12.0247
R874 VTAIL.n64 VTAIL.n63 12.0247
R875 VTAIL.n155 VTAIL.n142 11.249
R876 VTAIL.n23 VTAIL.n10 11.249
R877 VTAIL.n111 VTAIL.n98 11.249
R878 VTAIL.n67 VTAIL.n54 11.249
R879 VTAIL.n156 VTAIL.n140 10.4732
R880 VTAIL.n24 VTAIL.n8 10.4732
R881 VTAIL.n112 VTAIL.n96 10.4732
R882 VTAIL.n68 VTAIL.n52 10.4732
R883 VTAIL.n160 VTAIL.n159 9.69747
R884 VTAIL.n28 VTAIL.n27 9.69747
R885 VTAIL.n116 VTAIL.n115 9.69747
R886 VTAIL.n72 VTAIL.n71 9.69747
R887 VTAIL.n174 VTAIL.n173 9.45567
R888 VTAIL.n42 VTAIL.n41 9.45567
R889 VTAIL.n130 VTAIL.n129 9.45567
R890 VTAIL.n86 VTAIL.n85 9.45567
R891 VTAIL.n134 VTAIL.n133 9.3005
R892 VTAIL.n173 VTAIL.n172 9.3005
R893 VTAIL.n165 VTAIL.n164 9.3005
R894 VTAIL.n138 VTAIL.n137 9.3005
R895 VTAIL.n159 VTAIL.n158 9.3005
R896 VTAIL.n157 VTAIL.n156 9.3005
R897 VTAIL.n142 VTAIL.n141 9.3005
R898 VTAIL.n151 VTAIL.n150 9.3005
R899 VTAIL.n149 VTAIL.n148 9.3005
R900 VTAIL.n167 VTAIL.n166 9.3005
R901 VTAIL.n2 VTAIL.n1 9.3005
R902 VTAIL.n41 VTAIL.n40 9.3005
R903 VTAIL.n33 VTAIL.n32 9.3005
R904 VTAIL.n6 VTAIL.n5 9.3005
R905 VTAIL.n27 VTAIL.n26 9.3005
R906 VTAIL.n25 VTAIL.n24 9.3005
R907 VTAIL.n10 VTAIL.n9 9.3005
R908 VTAIL.n19 VTAIL.n18 9.3005
R909 VTAIL.n17 VTAIL.n16 9.3005
R910 VTAIL.n35 VTAIL.n34 9.3005
R911 VTAIL.n90 VTAIL.n89 9.3005
R912 VTAIL.n123 VTAIL.n122 9.3005
R913 VTAIL.n121 VTAIL.n120 9.3005
R914 VTAIL.n94 VTAIL.n93 9.3005
R915 VTAIL.n115 VTAIL.n114 9.3005
R916 VTAIL.n113 VTAIL.n112 9.3005
R917 VTAIL.n98 VTAIL.n97 9.3005
R918 VTAIL.n107 VTAIL.n106 9.3005
R919 VTAIL.n105 VTAIL.n104 9.3005
R920 VTAIL.n129 VTAIL.n128 9.3005
R921 VTAIL.n85 VTAIL.n84 9.3005
R922 VTAIL.n46 VTAIL.n45 9.3005
R923 VTAIL.n79 VTAIL.n78 9.3005
R924 VTAIL.n77 VTAIL.n76 9.3005
R925 VTAIL.n50 VTAIL.n49 9.3005
R926 VTAIL.n71 VTAIL.n70 9.3005
R927 VTAIL.n69 VTAIL.n68 9.3005
R928 VTAIL.n54 VTAIL.n53 9.3005
R929 VTAIL.n63 VTAIL.n62 9.3005
R930 VTAIL.n61 VTAIL.n60 9.3005
R931 VTAIL.n163 VTAIL.n138 8.92171
R932 VTAIL.n31 VTAIL.n6 8.92171
R933 VTAIL.n119 VTAIL.n94 8.92171
R934 VTAIL.n75 VTAIL.n50 8.92171
R935 VTAIL.n164 VTAIL.n136 8.14595
R936 VTAIL.n174 VTAIL.n132 8.14595
R937 VTAIL.n32 VTAIL.n4 8.14595
R938 VTAIL.n42 VTAIL.n0 8.14595
R939 VTAIL.n130 VTAIL.n88 8.14595
R940 VTAIL.n120 VTAIL.n92 8.14595
R941 VTAIL.n86 VTAIL.n44 8.14595
R942 VTAIL.n76 VTAIL.n48 8.14595
R943 VTAIL.n168 VTAIL.n167 7.3702
R944 VTAIL.n172 VTAIL.n171 7.3702
R945 VTAIL.n36 VTAIL.n35 7.3702
R946 VTAIL.n40 VTAIL.n39 7.3702
R947 VTAIL.n128 VTAIL.n127 7.3702
R948 VTAIL.n124 VTAIL.n123 7.3702
R949 VTAIL.n84 VTAIL.n83 7.3702
R950 VTAIL.n80 VTAIL.n79 7.3702
R951 VTAIL.n168 VTAIL.n134 6.59444
R952 VTAIL.n171 VTAIL.n134 6.59444
R953 VTAIL.n36 VTAIL.n2 6.59444
R954 VTAIL.n39 VTAIL.n2 6.59444
R955 VTAIL.n127 VTAIL.n90 6.59444
R956 VTAIL.n124 VTAIL.n90 6.59444
R957 VTAIL.n83 VTAIL.n46 6.59444
R958 VTAIL.n80 VTAIL.n46 6.59444
R959 VTAIL.n167 VTAIL.n136 5.81868
R960 VTAIL.n172 VTAIL.n132 5.81868
R961 VTAIL.n35 VTAIL.n4 5.81868
R962 VTAIL.n40 VTAIL.n0 5.81868
R963 VTAIL.n128 VTAIL.n88 5.81868
R964 VTAIL.n123 VTAIL.n92 5.81868
R965 VTAIL.n84 VTAIL.n44 5.81868
R966 VTAIL.n79 VTAIL.n48 5.81868
R967 VTAIL.n164 VTAIL.n163 5.04292
R968 VTAIL.n32 VTAIL.n31 5.04292
R969 VTAIL.n120 VTAIL.n119 5.04292
R970 VTAIL.n76 VTAIL.n75 5.04292
R971 VTAIL.n160 VTAIL.n138 4.26717
R972 VTAIL.n28 VTAIL.n6 4.26717
R973 VTAIL.n116 VTAIL.n94 4.26717
R974 VTAIL.n72 VTAIL.n50 4.26717
R975 VTAIL.n149 VTAIL.n145 3.70995
R976 VTAIL.n17 VTAIL.n13 3.70995
R977 VTAIL.n61 VTAIL.n57 3.70995
R978 VTAIL.n105 VTAIL.n101 3.70995
R979 VTAIL.n159 VTAIL.n140 3.49141
R980 VTAIL.n27 VTAIL.n8 3.49141
R981 VTAIL.n115 VTAIL.n96 3.49141
R982 VTAIL.n71 VTAIL.n52 3.49141
R983 VTAIL.n156 VTAIL.n155 2.71565
R984 VTAIL.n24 VTAIL.n23 2.71565
R985 VTAIL.n112 VTAIL.n111 2.71565
R986 VTAIL.n68 VTAIL.n67 2.71565
R987 VTAIL.n152 VTAIL.n142 1.93989
R988 VTAIL.n20 VTAIL.n10 1.93989
R989 VTAIL.n108 VTAIL.n98 1.93989
R990 VTAIL.n64 VTAIL.n54 1.93989
R991 VTAIL.n131 VTAIL.n87 1.82809
R992 VTAIL VTAIL.n43 1.2074
R993 VTAIL.n151 VTAIL.n144 1.16414
R994 VTAIL.n19 VTAIL.n12 1.16414
R995 VTAIL.n107 VTAIL.n100 1.16414
R996 VTAIL.n63 VTAIL.n56 1.16414
R997 VTAIL VTAIL.n175 0.62119
R998 VTAIL.n148 VTAIL.n147 0.388379
R999 VTAIL.n16 VTAIL.n15 0.388379
R1000 VTAIL.n104 VTAIL.n103 0.388379
R1001 VTAIL.n60 VTAIL.n59 0.388379
R1002 VTAIL.n150 VTAIL.n149 0.155672
R1003 VTAIL.n150 VTAIL.n141 0.155672
R1004 VTAIL.n157 VTAIL.n141 0.155672
R1005 VTAIL.n158 VTAIL.n157 0.155672
R1006 VTAIL.n158 VTAIL.n137 0.155672
R1007 VTAIL.n165 VTAIL.n137 0.155672
R1008 VTAIL.n166 VTAIL.n165 0.155672
R1009 VTAIL.n166 VTAIL.n133 0.155672
R1010 VTAIL.n173 VTAIL.n133 0.155672
R1011 VTAIL.n18 VTAIL.n17 0.155672
R1012 VTAIL.n18 VTAIL.n9 0.155672
R1013 VTAIL.n25 VTAIL.n9 0.155672
R1014 VTAIL.n26 VTAIL.n25 0.155672
R1015 VTAIL.n26 VTAIL.n5 0.155672
R1016 VTAIL.n33 VTAIL.n5 0.155672
R1017 VTAIL.n34 VTAIL.n33 0.155672
R1018 VTAIL.n34 VTAIL.n1 0.155672
R1019 VTAIL.n41 VTAIL.n1 0.155672
R1020 VTAIL.n129 VTAIL.n89 0.155672
R1021 VTAIL.n122 VTAIL.n89 0.155672
R1022 VTAIL.n122 VTAIL.n121 0.155672
R1023 VTAIL.n121 VTAIL.n93 0.155672
R1024 VTAIL.n114 VTAIL.n93 0.155672
R1025 VTAIL.n114 VTAIL.n113 0.155672
R1026 VTAIL.n113 VTAIL.n97 0.155672
R1027 VTAIL.n106 VTAIL.n97 0.155672
R1028 VTAIL.n106 VTAIL.n105 0.155672
R1029 VTAIL.n85 VTAIL.n45 0.155672
R1030 VTAIL.n78 VTAIL.n45 0.155672
R1031 VTAIL.n78 VTAIL.n77 0.155672
R1032 VTAIL.n77 VTAIL.n49 0.155672
R1033 VTAIL.n70 VTAIL.n49 0.155672
R1034 VTAIL.n70 VTAIL.n69 0.155672
R1035 VTAIL.n69 VTAIL.n53 0.155672
R1036 VTAIL.n62 VTAIL.n53 0.155672
R1037 VTAIL.n62 VTAIL.n61 0.155672
R1038 VDD1.n38 VDD1.n0 756.745
R1039 VDD1.n81 VDD1.n43 756.745
R1040 VDD1.n39 VDD1.n38 585
R1041 VDD1.n37 VDD1.n36 585
R1042 VDD1.n4 VDD1.n3 585
R1043 VDD1.n31 VDD1.n30 585
R1044 VDD1.n29 VDD1.n28 585
R1045 VDD1.n8 VDD1.n7 585
R1046 VDD1.n23 VDD1.n22 585
R1047 VDD1.n21 VDD1.n20 585
R1048 VDD1.n12 VDD1.n11 585
R1049 VDD1.n15 VDD1.n14 585
R1050 VDD1.n58 VDD1.n57 585
R1051 VDD1.n55 VDD1.n54 585
R1052 VDD1.n64 VDD1.n63 585
R1053 VDD1.n66 VDD1.n65 585
R1054 VDD1.n51 VDD1.n50 585
R1055 VDD1.n72 VDD1.n71 585
R1056 VDD1.n74 VDD1.n73 585
R1057 VDD1.n47 VDD1.n46 585
R1058 VDD1.n80 VDD1.n79 585
R1059 VDD1.n82 VDD1.n81 585
R1060 VDD1.t1 VDD1.n13 327.473
R1061 VDD1.t0 VDD1.n56 327.473
R1062 VDD1.n38 VDD1.n37 171.744
R1063 VDD1.n37 VDD1.n3 171.744
R1064 VDD1.n30 VDD1.n3 171.744
R1065 VDD1.n30 VDD1.n29 171.744
R1066 VDD1.n29 VDD1.n7 171.744
R1067 VDD1.n22 VDD1.n7 171.744
R1068 VDD1.n22 VDD1.n21 171.744
R1069 VDD1.n21 VDD1.n11 171.744
R1070 VDD1.n14 VDD1.n11 171.744
R1071 VDD1.n57 VDD1.n54 171.744
R1072 VDD1.n64 VDD1.n54 171.744
R1073 VDD1.n65 VDD1.n64 171.744
R1074 VDD1.n65 VDD1.n50 171.744
R1075 VDD1.n72 VDD1.n50 171.744
R1076 VDD1.n73 VDD1.n72 171.744
R1077 VDD1.n73 VDD1.n46 171.744
R1078 VDD1.n80 VDD1.n46 171.744
R1079 VDD1.n81 VDD1.n80 171.744
R1080 VDD1.n14 VDD1.t1 85.8723
R1081 VDD1.n57 VDD1.t0 85.8723
R1082 VDD1 VDD1.n85 85.18
R1083 VDD1 VDD1.n42 48.6315
R1084 VDD1.n15 VDD1.n13 16.3894
R1085 VDD1.n58 VDD1.n56 16.3894
R1086 VDD1.n16 VDD1.n12 12.8005
R1087 VDD1.n59 VDD1.n55 12.8005
R1088 VDD1.n20 VDD1.n19 12.0247
R1089 VDD1.n63 VDD1.n62 12.0247
R1090 VDD1.n23 VDD1.n10 11.249
R1091 VDD1.n66 VDD1.n53 11.249
R1092 VDD1.n24 VDD1.n8 10.4732
R1093 VDD1.n67 VDD1.n51 10.4732
R1094 VDD1.n28 VDD1.n27 9.69747
R1095 VDD1.n71 VDD1.n70 9.69747
R1096 VDD1.n42 VDD1.n41 9.45567
R1097 VDD1.n85 VDD1.n84 9.45567
R1098 VDD1.n2 VDD1.n1 9.3005
R1099 VDD1.n35 VDD1.n34 9.3005
R1100 VDD1.n33 VDD1.n32 9.3005
R1101 VDD1.n6 VDD1.n5 9.3005
R1102 VDD1.n27 VDD1.n26 9.3005
R1103 VDD1.n25 VDD1.n24 9.3005
R1104 VDD1.n10 VDD1.n9 9.3005
R1105 VDD1.n19 VDD1.n18 9.3005
R1106 VDD1.n17 VDD1.n16 9.3005
R1107 VDD1.n41 VDD1.n40 9.3005
R1108 VDD1.n45 VDD1.n44 9.3005
R1109 VDD1.n84 VDD1.n83 9.3005
R1110 VDD1.n76 VDD1.n75 9.3005
R1111 VDD1.n49 VDD1.n48 9.3005
R1112 VDD1.n70 VDD1.n69 9.3005
R1113 VDD1.n68 VDD1.n67 9.3005
R1114 VDD1.n53 VDD1.n52 9.3005
R1115 VDD1.n62 VDD1.n61 9.3005
R1116 VDD1.n60 VDD1.n59 9.3005
R1117 VDD1.n78 VDD1.n77 9.3005
R1118 VDD1.n31 VDD1.n6 8.92171
R1119 VDD1.n74 VDD1.n49 8.92171
R1120 VDD1.n42 VDD1.n0 8.14595
R1121 VDD1.n32 VDD1.n4 8.14595
R1122 VDD1.n75 VDD1.n47 8.14595
R1123 VDD1.n85 VDD1.n43 8.14595
R1124 VDD1.n40 VDD1.n39 7.3702
R1125 VDD1.n36 VDD1.n35 7.3702
R1126 VDD1.n79 VDD1.n78 7.3702
R1127 VDD1.n83 VDD1.n82 7.3702
R1128 VDD1.n39 VDD1.n2 6.59444
R1129 VDD1.n36 VDD1.n2 6.59444
R1130 VDD1.n79 VDD1.n45 6.59444
R1131 VDD1.n82 VDD1.n45 6.59444
R1132 VDD1.n40 VDD1.n0 5.81868
R1133 VDD1.n35 VDD1.n4 5.81868
R1134 VDD1.n78 VDD1.n47 5.81868
R1135 VDD1.n83 VDD1.n43 5.81868
R1136 VDD1.n32 VDD1.n31 5.04292
R1137 VDD1.n75 VDD1.n74 5.04292
R1138 VDD1.n28 VDD1.n6 4.26717
R1139 VDD1.n71 VDD1.n49 4.26717
R1140 VDD1.n60 VDD1.n56 3.70995
R1141 VDD1.n17 VDD1.n13 3.70995
R1142 VDD1.n27 VDD1.n8 3.49141
R1143 VDD1.n70 VDD1.n51 3.49141
R1144 VDD1.n24 VDD1.n23 2.71565
R1145 VDD1.n67 VDD1.n66 2.71565
R1146 VDD1.n20 VDD1.n10 1.93989
R1147 VDD1.n63 VDD1.n53 1.93989
R1148 VDD1.n19 VDD1.n12 1.16414
R1149 VDD1.n62 VDD1.n55 1.16414
R1150 VDD1.n16 VDD1.n15 0.388379
R1151 VDD1.n59 VDD1.n58 0.388379
R1152 VDD1.n41 VDD1.n1 0.155672
R1153 VDD1.n34 VDD1.n1 0.155672
R1154 VDD1.n34 VDD1.n33 0.155672
R1155 VDD1.n33 VDD1.n5 0.155672
R1156 VDD1.n26 VDD1.n5 0.155672
R1157 VDD1.n26 VDD1.n25 0.155672
R1158 VDD1.n25 VDD1.n9 0.155672
R1159 VDD1.n18 VDD1.n9 0.155672
R1160 VDD1.n18 VDD1.n17 0.155672
R1161 VDD1.n61 VDD1.n60 0.155672
R1162 VDD1.n61 VDD1.n52 0.155672
R1163 VDD1.n68 VDD1.n52 0.155672
R1164 VDD1.n69 VDD1.n68 0.155672
R1165 VDD1.n69 VDD1.n48 0.155672
R1166 VDD1.n76 VDD1.n48 0.155672
R1167 VDD1.n77 VDD1.n76 0.155672
R1168 VDD1.n77 VDD1.n44 0.155672
R1169 VDD1.n84 VDD1.n44 0.155672
R1170 VN VN.t0 152.7
R1171 VN VN.t1 110.837
R1172 VDD2.n81 VDD2.n43 756.745
R1173 VDD2.n38 VDD2.n0 756.745
R1174 VDD2.n82 VDD2.n81 585
R1175 VDD2.n80 VDD2.n79 585
R1176 VDD2.n47 VDD2.n46 585
R1177 VDD2.n74 VDD2.n73 585
R1178 VDD2.n72 VDD2.n71 585
R1179 VDD2.n51 VDD2.n50 585
R1180 VDD2.n66 VDD2.n65 585
R1181 VDD2.n64 VDD2.n63 585
R1182 VDD2.n55 VDD2.n54 585
R1183 VDD2.n58 VDD2.n57 585
R1184 VDD2.n15 VDD2.n14 585
R1185 VDD2.n12 VDD2.n11 585
R1186 VDD2.n21 VDD2.n20 585
R1187 VDD2.n23 VDD2.n22 585
R1188 VDD2.n8 VDD2.n7 585
R1189 VDD2.n29 VDD2.n28 585
R1190 VDD2.n31 VDD2.n30 585
R1191 VDD2.n4 VDD2.n3 585
R1192 VDD2.n37 VDD2.n36 585
R1193 VDD2.n39 VDD2.n38 585
R1194 VDD2.t1 VDD2.n56 327.473
R1195 VDD2.t0 VDD2.n13 327.473
R1196 VDD2.n81 VDD2.n80 171.744
R1197 VDD2.n80 VDD2.n46 171.744
R1198 VDD2.n73 VDD2.n46 171.744
R1199 VDD2.n73 VDD2.n72 171.744
R1200 VDD2.n72 VDD2.n50 171.744
R1201 VDD2.n65 VDD2.n50 171.744
R1202 VDD2.n65 VDD2.n64 171.744
R1203 VDD2.n64 VDD2.n54 171.744
R1204 VDD2.n57 VDD2.n54 171.744
R1205 VDD2.n14 VDD2.n11 171.744
R1206 VDD2.n21 VDD2.n11 171.744
R1207 VDD2.n22 VDD2.n21 171.744
R1208 VDD2.n22 VDD2.n7 171.744
R1209 VDD2.n29 VDD2.n7 171.744
R1210 VDD2.n30 VDD2.n29 171.744
R1211 VDD2.n30 VDD2.n3 171.744
R1212 VDD2.n37 VDD2.n3 171.744
R1213 VDD2.n38 VDD2.n37 171.744
R1214 VDD2.n57 VDD2.t1 85.8723
R1215 VDD2.n14 VDD2.t0 85.8723
R1216 VDD2.n86 VDD2.n42 83.9763
R1217 VDD2.n86 VDD2.n85 47.8944
R1218 VDD2.n58 VDD2.n56 16.3894
R1219 VDD2.n15 VDD2.n13 16.3894
R1220 VDD2.n59 VDD2.n55 12.8005
R1221 VDD2.n16 VDD2.n12 12.8005
R1222 VDD2.n63 VDD2.n62 12.0247
R1223 VDD2.n20 VDD2.n19 12.0247
R1224 VDD2.n66 VDD2.n53 11.249
R1225 VDD2.n23 VDD2.n10 11.249
R1226 VDD2.n67 VDD2.n51 10.4732
R1227 VDD2.n24 VDD2.n8 10.4732
R1228 VDD2.n71 VDD2.n70 9.69747
R1229 VDD2.n28 VDD2.n27 9.69747
R1230 VDD2.n85 VDD2.n84 9.45567
R1231 VDD2.n42 VDD2.n41 9.45567
R1232 VDD2.n45 VDD2.n44 9.3005
R1233 VDD2.n78 VDD2.n77 9.3005
R1234 VDD2.n76 VDD2.n75 9.3005
R1235 VDD2.n49 VDD2.n48 9.3005
R1236 VDD2.n70 VDD2.n69 9.3005
R1237 VDD2.n68 VDD2.n67 9.3005
R1238 VDD2.n53 VDD2.n52 9.3005
R1239 VDD2.n62 VDD2.n61 9.3005
R1240 VDD2.n60 VDD2.n59 9.3005
R1241 VDD2.n84 VDD2.n83 9.3005
R1242 VDD2.n2 VDD2.n1 9.3005
R1243 VDD2.n41 VDD2.n40 9.3005
R1244 VDD2.n33 VDD2.n32 9.3005
R1245 VDD2.n6 VDD2.n5 9.3005
R1246 VDD2.n27 VDD2.n26 9.3005
R1247 VDD2.n25 VDD2.n24 9.3005
R1248 VDD2.n10 VDD2.n9 9.3005
R1249 VDD2.n19 VDD2.n18 9.3005
R1250 VDD2.n17 VDD2.n16 9.3005
R1251 VDD2.n35 VDD2.n34 9.3005
R1252 VDD2.n74 VDD2.n49 8.92171
R1253 VDD2.n31 VDD2.n6 8.92171
R1254 VDD2.n85 VDD2.n43 8.14595
R1255 VDD2.n75 VDD2.n47 8.14595
R1256 VDD2.n32 VDD2.n4 8.14595
R1257 VDD2.n42 VDD2.n0 8.14595
R1258 VDD2.n83 VDD2.n82 7.3702
R1259 VDD2.n79 VDD2.n78 7.3702
R1260 VDD2.n36 VDD2.n35 7.3702
R1261 VDD2.n40 VDD2.n39 7.3702
R1262 VDD2.n82 VDD2.n45 6.59444
R1263 VDD2.n79 VDD2.n45 6.59444
R1264 VDD2.n36 VDD2.n2 6.59444
R1265 VDD2.n39 VDD2.n2 6.59444
R1266 VDD2.n83 VDD2.n43 5.81868
R1267 VDD2.n78 VDD2.n47 5.81868
R1268 VDD2.n35 VDD2.n4 5.81868
R1269 VDD2.n40 VDD2.n0 5.81868
R1270 VDD2.n75 VDD2.n74 5.04292
R1271 VDD2.n32 VDD2.n31 5.04292
R1272 VDD2.n71 VDD2.n49 4.26717
R1273 VDD2.n28 VDD2.n6 4.26717
R1274 VDD2.n17 VDD2.n13 3.70995
R1275 VDD2.n60 VDD2.n56 3.70995
R1276 VDD2.n70 VDD2.n51 3.49141
R1277 VDD2.n27 VDD2.n8 3.49141
R1278 VDD2.n67 VDD2.n66 2.71565
R1279 VDD2.n24 VDD2.n23 2.71565
R1280 VDD2.n63 VDD2.n53 1.93989
R1281 VDD2.n20 VDD2.n10 1.93989
R1282 VDD2.n62 VDD2.n55 1.16414
R1283 VDD2.n19 VDD2.n12 1.16414
R1284 VDD2 VDD2.n86 0.737569
R1285 VDD2.n59 VDD2.n58 0.388379
R1286 VDD2.n16 VDD2.n15 0.388379
R1287 VDD2.n84 VDD2.n44 0.155672
R1288 VDD2.n77 VDD2.n44 0.155672
R1289 VDD2.n77 VDD2.n76 0.155672
R1290 VDD2.n76 VDD2.n48 0.155672
R1291 VDD2.n69 VDD2.n48 0.155672
R1292 VDD2.n69 VDD2.n68 0.155672
R1293 VDD2.n68 VDD2.n52 0.155672
R1294 VDD2.n61 VDD2.n52 0.155672
R1295 VDD2.n61 VDD2.n60 0.155672
R1296 VDD2.n18 VDD2.n17 0.155672
R1297 VDD2.n18 VDD2.n9 0.155672
R1298 VDD2.n25 VDD2.n9 0.155672
R1299 VDD2.n26 VDD2.n25 0.155672
R1300 VDD2.n26 VDD2.n5 0.155672
R1301 VDD2.n33 VDD2.n5 0.155672
R1302 VDD2.n34 VDD2.n33 0.155672
R1303 VDD2.n34 VDD2.n1 0.155672
R1304 VDD2.n41 VDD2.n1 0.155672
C0 VDD1 w_n2230_n2590# 1.53674f
C1 VN VDD2 1.98227f
C2 VTAIL VDD1 4.08726f
C3 VP VDD2 0.342011f
C4 w_n2230_n2590# B 7.95576f
C5 VN VP 4.83987f
C6 VTAIL B 2.85969f
C7 w_n2230_n2590# VDD2 1.56534f
C8 VDD1 B 1.42638f
C9 VN w_n2230_n2590# 3.03486f
C10 VTAIL VDD2 4.14041f
C11 VTAIL VN 1.84337f
C12 w_n2230_n2590# VP 3.31939f
C13 VTAIL VP 1.85758f
C14 VDD1 VDD2 0.700799f
C15 VDD1 VN 0.148223f
C16 VDD1 VP 2.17427f
C17 VDD2 B 1.45841f
C18 VN B 1.04128f
C19 VTAIL w_n2230_n2590# 2.20591f
C20 VP B 1.50995f
C21 VDD2 VSUBS 0.741508f
C22 VDD1 VSUBS 3.352813f
C23 VTAIL VSUBS 0.840954f
C24 VN VSUBS 5.604179f
C25 VP VSUBS 1.604308f
C26 B VSUBS 3.742006f
C27 w_n2230_n2590# VSUBS 71.6365f
C28 VDD2.n0 VSUBS 0.015588f
C29 VDD2.n1 VSUBS 0.013865f
C30 VDD2.n2 VSUBS 0.007451f
C31 VDD2.n3 VSUBS 0.01761f
C32 VDD2.n4 VSUBS 0.007889f
C33 VDD2.n5 VSUBS 0.013865f
C34 VDD2.n6 VSUBS 0.007451f
C35 VDD2.n7 VSUBS 0.01761f
C36 VDD2.n8 VSUBS 0.007889f
C37 VDD2.n9 VSUBS 0.013865f
C38 VDD2.n10 VSUBS 0.007451f
C39 VDD2.n11 VSUBS 0.01761f
C40 VDD2.n12 VSUBS 0.007889f
C41 VDD2.n13 VSUBS 0.069652f
C42 VDD2.t0 VSUBS 0.037556f
C43 VDD2.n14 VSUBS 0.013208f
C44 VDD2.n15 VSUBS 0.011203f
C45 VDD2.n16 VSUBS 0.007451f
C46 VDD2.n17 VSUBS 0.451448f
C47 VDD2.n18 VSUBS 0.013865f
C48 VDD2.n19 VSUBS 0.007451f
C49 VDD2.n20 VSUBS 0.007889f
C50 VDD2.n21 VSUBS 0.01761f
C51 VDD2.n22 VSUBS 0.01761f
C52 VDD2.n23 VSUBS 0.007889f
C53 VDD2.n24 VSUBS 0.007451f
C54 VDD2.n25 VSUBS 0.013865f
C55 VDD2.n26 VSUBS 0.013865f
C56 VDD2.n27 VSUBS 0.007451f
C57 VDD2.n28 VSUBS 0.007889f
C58 VDD2.n29 VSUBS 0.01761f
C59 VDD2.n30 VSUBS 0.01761f
C60 VDD2.n31 VSUBS 0.007889f
C61 VDD2.n32 VSUBS 0.007451f
C62 VDD2.n33 VSUBS 0.013865f
C63 VDD2.n34 VSUBS 0.013865f
C64 VDD2.n35 VSUBS 0.007451f
C65 VDD2.n36 VSUBS 0.007889f
C66 VDD2.n37 VSUBS 0.01761f
C67 VDD2.n38 VSUBS 0.043837f
C68 VDD2.n39 VSUBS 0.007889f
C69 VDD2.n40 VSUBS 0.007451f
C70 VDD2.n41 VSUBS 0.031102f
C71 VDD2.n42 VSUBS 0.345676f
C72 VDD2.n43 VSUBS 0.015588f
C73 VDD2.n44 VSUBS 0.013865f
C74 VDD2.n45 VSUBS 0.007451f
C75 VDD2.n46 VSUBS 0.01761f
C76 VDD2.n47 VSUBS 0.007889f
C77 VDD2.n48 VSUBS 0.013865f
C78 VDD2.n49 VSUBS 0.007451f
C79 VDD2.n50 VSUBS 0.01761f
C80 VDD2.n51 VSUBS 0.007889f
C81 VDD2.n52 VSUBS 0.013865f
C82 VDD2.n53 VSUBS 0.007451f
C83 VDD2.n54 VSUBS 0.01761f
C84 VDD2.n55 VSUBS 0.007889f
C85 VDD2.n56 VSUBS 0.069652f
C86 VDD2.t1 VSUBS 0.037556f
C87 VDD2.n57 VSUBS 0.013208f
C88 VDD2.n58 VSUBS 0.011203f
C89 VDD2.n59 VSUBS 0.007451f
C90 VDD2.n60 VSUBS 0.451447f
C91 VDD2.n61 VSUBS 0.013865f
C92 VDD2.n62 VSUBS 0.007451f
C93 VDD2.n63 VSUBS 0.007889f
C94 VDD2.n64 VSUBS 0.01761f
C95 VDD2.n65 VSUBS 0.01761f
C96 VDD2.n66 VSUBS 0.007889f
C97 VDD2.n67 VSUBS 0.007451f
C98 VDD2.n68 VSUBS 0.013865f
C99 VDD2.n69 VSUBS 0.013865f
C100 VDD2.n70 VSUBS 0.007451f
C101 VDD2.n71 VSUBS 0.007889f
C102 VDD2.n72 VSUBS 0.01761f
C103 VDD2.n73 VSUBS 0.01761f
C104 VDD2.n74 VSUBS 0.007889f
C105 VDD2.n75 VSUBS 0.007451f
C106 VDD2.n76 VSUBS 0.013865f
C107 VDD2.n77 VSUBS 0.013865f
C108 VDD2.n78 VSUBS 0.007451f
C109 VDD2.n79 VSUBS 0.007889f
C110 VDD2.n80 VSUBS 0.01761f
C111 VDD2.n81 VSUBS 0.043837f
C112 VDD2.n82 VSUBS 0.007889f
C113 VDD2.n83 VSUBS 0.007451f
C114 VDD2.n84 VSUBS 0.031102f
C115 VDD2.n85 VSUBS 0.03165f
C116 VDD2.n86 VSUBS 1.4869f
C117 VN.t1 VSUBS 2.03208f
C118 VN.t0 VSUBS 2.54088f
C119 VDD1.n0 VSUBS 0.023657f
C120 VDD1.n1 VSUBS 0.021042f
C121 VDD1.n2 VSUBS 0.011307f
C122 VDD1.n3 VSUBS 0.026726f
C123 VDD1.n4 VSUBS 0.011972f
C124 VDD1.n5 VSUBS 0.021042f
C125 VDD1.n6 VSUBS 0.011307f
C126 VDD1.n7 VSUBS 0.026726f
C127 VDD1.n8 VSUBS 0.011972f
C128 VDD1.n9 VSUBS 0.021042f
C129 VDD1.n10 VSUBS 0.011307f
C130 VDD1.n11 VSUBS 0.026726f
C131 VDD1.n12 VSUBS 0.011972f
C132 VDD1.n13 VSUBS 0.105707f
C133 VDD1.t1 VSUBS 0.056997f
C134 VDD1.n14 VSUBS 0.020045f
C135 VDD1.n15 VSUBS 0.017001f
C136 VDD1.n16 VSUBS 0.011307f
C137 VDD1.n17 VSUBS 0.68513f
C138 VDD1.n18 VSUBS 0.021042f
C139 VDD1.n19 VSUBS 0.011307f
C140 VDD1.n20 VSUBS 0.011972f
C141 VDD1.n21 VSUBS 0.026726f
C142 VDD1.n22 VSUBS 0.026726f
C143 VDD1.n23 VSUBS 0.011972f
C144 VDD1.n24 VSUBS 0.011307f
C145 VDD1.n25 VSUBS 0.021042f
C146 VDD1.n26 VSUBS 0.021042f
C147 VDD1.n27 VSUBS 0.011307f
C148 VDD1.n28 VSUBS 0.011972f
C149 VDD1.n29 VSUBS 0.026726f
C150 VDD1.n30 VSUBS 0.026726f
C151 VDD1.n31 VSUBS 0.011972f
C152 VDD1.n32 VSUBS 0.011307f
C153 VDD1.n33 VSUBS 0.021042f
C154 VDD1.n34 VSUBS 0.021042f
C155 VDD1.n35 VSUBS 0.011307f
C156 VDD1.n36 VSUBS 0.011972f
C157 VDD1.n37 VSUBS 0.026726f
C158 VDD1.n38 VSUBS 0.066528f
C159 VDD1.n39 VSUBS 0.011972f
C160 VDD1.n40 VSUBS 0.011307f
C161 VDD1.n41 VSUBS 0.047201f
C162 VDD1.n42 VSUBS 0.049393f
C163 VDD1.n43 VSUBS 0.023657f
C164 VDD1.n44 VSUBS 0.021042f
C165 VDD1.n45 VSUBS 0.011307f
C166 VDD1.n46 VSUBS 0.026726f
C167 VDD1.n47 VSUBS 0.011972f
C168 VDD1.n48 VSUBS 0.021042f
C169 VDD1.n49 VSUBS 0.011307f
C170 VDD1.n50 VSUBS 0.026726f
C171 VDD1.n51 VSUBS 0.011972f
C172 VDD1.n52 VSUBS 0.021042f
C173 VDD1.n53 VSUBS 0.011307f
C174 VDD1.n54 VSUBS 0.026726f
C175 VDD1.n55 VSUBS 0.011972f
C176 VDD1.n56 VSUBS 0.105707f
C177 VDD1.t0 VSUBS 0.056997f
C178 VDD1.n57 VSUBS 0.020045f
C179 VDD1.n58 VSUBS 0.017001f
C180 VDD1.n59 VSUBS 0.011307f
C181 VDD1.n60 VSUBS 0.68513f
C182 VDD1.n61 VSUBS 0.021042f
C183 VDD1.n62 VSUBS 0.011307f
C184 VDD1.n63 VSUBS 0.011972f
C185 VDD1.n64 VSUBS 0.026726f
C186 VDD1.n65 VSUBS 0.026726f
C187 VDD1.n66 VSUBS 0.011972f
C188 VDD1.n67 VSUBS 0.011307f
C189 VDD1.n68 VSUBS 0.021042f
C190 VDD1.n69 VSUBS 0.021042f
C191 VDD1.n70 VSUBS 0.011307f
C192 VDD1.n71 VSUBS 0.011972f
C193 VDD1.n72 VSUBS 0.026726f
C194 VDD1.n73 VSUBS 0.026726f
C195 VDD1.n74 VSUBS 0.011972f
C196 VDD1.n75 VSUBS 0.011307f
C197 VDD1.n76 VSUBS 0.021042f
C198 VDD1.n77 VSUBS 0.021042f
C199 VDD1.n78 VSUBS 0.011307f
C200 VDD1.n79 VSUBS 0.011972f
C201 VDD1.n80 VSUBS 0.026726f
C202 VDD1.n81 VSUBS 0.066528f
C203 VDD1.n82 VSUBS 0.011972f
C204 VDD1.n83 VSUBS 0.011307f
C205 VDD1.n84 VSUBS 0.047201f
C206 VDD1.n85 VSUBS 0.564856f
C207 VTAIL.n0 VSUBS 0.027738f
C208 VTAIL.n1 VSUBS 0.024672f
C209 VTAIL.n2 VSUBS 0.013257f
C210 VTAIL.n3 VSUBS 0.031336f
C211 VTAIL.n4 VSUBS 0.014037f
C212 VTAIL.n5 VSUBS 0.024672f
C213 VTAIL.n6 VSUBS 0.013257f
C214 VTAIL.n7 VSUBS 0.031336f
C215 VTAIL.n8 VSUBS 0.014037f
C216 VTAIL.n9 VSUBS 0.024672f
C217 VTAIL.n10 VSUBS 0.013257f
C218 VTAIL.n11 VSUBS 0.031336f
C219 VTAIL.n12 VSUBS 0.014037f
C220 VTAIL.n13 VSUBS 0.12394f
C221 VTAIL.t2 VSUBS 0.066828f
C222 VTAIL.n14 VSUBS 0.023502f
C223 VTAIL.n15 VSUBS 0.019934f
C224 VTAIL.n16 VSUBS 0.013257f
C225 VTAIL.n17 VSUBS 0.803309f
C226 VTAIL.n18 VSUBS 0.024672f
C227 VTAIL.n19 VSUBS 0.013257f
C228 VTAIL.n20 VSUBS 0.014037f
C229 VTAIL.n21 VSUBS 0.031336f
C230 VTAIL.n22 VSUBS 0.031336f
C231 VTAIL.n23 VSUBS 0.014037f
C232 VTAIL.n24 VSUBS 0.013257f
C233 VTAIL.n25 VSUBS 0.024672f
C234 VTAIL.n26 VSUBS 0.024672f
C235 VTAIL.n27 VSUBS 0.013257f
C236 VTAIL.n28 VSUBS 0.014037f
C237 VTAIL.n29 VSUBS 0.031336f
C238 VTAIL.n30 VSUBS 0.031336f
C239 VTAIL.n31 VSUBS 0.014037f
C240 VTAIL.n32 VSUBS 0.013257f
C241 VTAIL.n33 VSUBS 0.024672f
C242 VTAIL.n34 VSUBS 0.024672f
C243 VTAIL.n35 VSUBS 0.013257f
C244 VTAIL.n36 VSUBS 0.014037f
C245 VTAIL.n37 VSUBS 0.031336f
C246 VTAIL.n38 VSUBS 0.078003f
C247 VTAIL.n39 VSUBS 0.014037f
C248 VTAIL.n40 VSUBS 0.013257f
C249 VTAIL.n41 VSUBS 0.055342f
C250 VTAIL.n42 VSUBS 0.03927f
C251 VTAIL.n43 VSUBS 1.43876f
C252 VTAIL.n44 VSUBS 0.027738f
C253 VTAIL.n45 VSUBS 0.024672f
C254 VTAIL.n46 VSUBS 0.013257f
C255 VTAIL.n47 VSUBS 0.031336f
C256 VTAIL.n48 VSUBS 0.014037f
C257 VTAIL.n49 VSUBS 0.024672f
C258 VTAIL.n50 VSUBS 0.013257f
C259 VTAIL.n51 VSUBS 0.031336f
C260 VTAIL.n52 VSUBS 0.014037f
C261 VTAIL.n53 VSUBS 0.024672f
C262 VTAIL.n54 VSUBS 0.013257f
C263 VTAIL.n55 VSUBS 0.031336f
C264 VTAIL.n56 VSUBS 0.014037f
C265 VTAIL.n57 VSUBS 0.12394f
C266 VTAIL.t1 VSUBS 0.066828f
C267 VTAIL.n58 VSUBS 0.023502f
C268 VTAIL.n59 VSUBS 0.019934f
C269 VTAIL.n60 VSUBS 0.013257f
C270 VTAIL.n61 VSUBS 0.803309f
C271 VTAIL.n62 VSUBS 0.024672f
C272 VTAIL.n63 VSUBS 0.013257f
C273 VTAIL.n64 VSUBS 0.014037f
C274 VTAIL.n65 VSUBS 0.031336f
C275 VTAIL.n66 VSUBS 0.031336f
C276 VTAIL.n67 VSUBS 0.014037f
C277 VTAIL.n68 VSUBS 0.013257f
C278 VTAIL.n69 VSUBS 0.024672f
C279 VTAIL.n70 VSUBS 0.024672f
C280 VTAIL.n71 VSUBS 0.013257f
C281 VTAIL.n72 VSUBS 0.014037f
C282 VTAIL.n73 VSUBS 0.031336f
C283 VTAIL.n74 VSUBS 0.031336f
C284 VTAIL.n75 VSUBS 0.014037f
C285 VTAIL.n76 VSUBS 0.013257f
C286 VTAIL.n77 VSUBS 0.024672f
C287 VTAIL.n78 VSUBS 0.024672f
C288 VTAIL.n79 VSUBS 0.013257f
C289 VTAIL.n80 VSUBS 0.014037f
C290 VTAIL.n81 VSUBS 0.031336f
C291 VTAIL.n82 VSUBS 0.078003f
C292 VTAIL.n83 VSUBS 0.014037f
C293 VTAIL.n84 VSUBS 0.013257f
C294 VTAIL.n85 VSUBS 0.055342f
C295 VTAIL.n86 VSUBS 0.03927f
C296 VTAIL.n87 VSUBS 1.4881f
C297 VTAIL.n88 VSUBS 0.027738f
C298 VTAIL.n89 VSUBS 0.024672f
C299 VTAIL.n90 VSUBS 0.013257f
C300 VTAIL.n91 VSUBS 0.031336f
C301 VTAIL.n92 VSUBS 0.014037f
C302 VTAIL.n93 VSUBS 0.024672f
C303 VTAIL.n94 VSUBS 0.013257f
C304 VTAIL.n95 VSUBS 0.031336f
C305 VTAIL.n96 VSUBS 0.014037f
C306 VTAIL.n97 VSUBS 0.024672f
C307 VTAIL.n98 VSUBS 0.013257f
C308 VTAIL.n99 VSUBS 0.031336f
C309 VTAIL.n100 VSUBS 0.014037f
C310 VTAIL.n101 VSUBS 0.12394f
C311 VTAIL.t3 VSUBS 0.066828f
C312 VTAIL.n102 VSUBS 0.023502f
C313 VTAIL.n103 VSUBS 0.019934f
C314 VTAIL.n104 VSUBS 0.013257f
C315 VTAIL.n105 VSUBS 0.803308f
C316 VTAIL.n106 VSUBS 0.024672f
C317 VTAIL.n107 VSUBS 0.013257f
C318 VTAIL.n108 VSUBS 0.014037f
C319 VTAIL.n109 VSUBS 0.031336f
C320 VTAIL.n110 VSUBS 0.031336f
C321 VTAIL.n111 VSUBS 0.014037f
C322 VTAIL.n112 VSUBS 0.013257f
C323 VTAIL.n113 VSUBS 0.024672f
C324 VTAIL.n114 VSUBS 0.024672f
C325 VTAIL.n115 VSUBS 0.013257f
C326 VTAIL.n116 VSUBS 0.014037f
C327 VTAIL.n117 VSUBS 0.031336f
C328 VTAIL.n118 VSUBS 0.031336f
C329 VTAIL.n119 VSUBS 0.014037f
C330 VTAIL.n120 VSUBS 0.013257f
C331 VTAIL.n121 VSUBS 0.024672f
C332 VTAIL.n122 VSUBS 0.024672f
C333 VTAIL.n123 VSUBS 0.013257f
C334 VTAIL.n124 VSUBS 0.014037f
C335 VTAIL.n125 VSUBS 0.031336f
C336 VTAIL.n126 VSUBS 0.078003f
C337 VTAIL.n127 VSUBS 0.014037f
C338 VTAIL.n128 VSUBS 0.013257f
C339 VTAIL.n129 VSUBS 0.055342f
C340 VTAIL.n130 VSUBS 0.03927f
C341 VTAIL.n131 VSUBS 1.27222f
C342 VTAIL.n132 VSUBS 0.027738f
C343 VTAIL.n133 VSUBS 0.024672f
C344 VTAIL.n134 VSUBS 0.013257f
C345 VTAIL.n135 VSUBS 0.031336f
C346 VTAIL.n136 VSUBS 0.014037f
C347 VTAIL.n137 VSUBS 0.024672f
C348 VTAIL.n138 VSUBS 0.013257f
C349 VTAIL.n139 VSUBS 0.031336f
C350 VTAIL.n140 VSUBS 0.014037f
C351 VTAIL.n141 VSUBS 0.024672f
C352 VTAIL.n142 VSUBS 0.013257f
C353 VTAIL.n143 VSUBS 0.031336f
C354 VTAIL.n144 VSUBS 0.014037f
C355 VTAIL.n145 VSUBS 0.12394f
C356 VTAIL.t0 VSUBS 0.066828f
C357 VTAIL.n146 VSUBS 0.023502f
C358 VTAIL.n147 VSUBS 0.019934f
C359 VTAIL.n148 VSUBS 0.013257f
C360 VTAIL.n149 VSUBS 0.803309f
C361 VTAIL.n150 VSUBS 0.024672f
C362 VTAIL.n151 VSUBS 0.013257f
C363 VTAIL.n152 VSUBS 0.014037f
C364 VTAIL.n153 VSUBS 0.031336f
C365 VTAIL.n154 VSUBS 0.031336f
C366 VTAIL.n155 VSUBS 0.014037f
C367 VTAIL.n156 VSUBS 0.013257f
C368 VTAIL.n157 VSUBS 0.024672f
C369 VTAIL.n158 VSUBS 0.024672f
C370 VTAIL.n159 VSUBS 0.013257f
C371 VTAIL.n160 VSUBS 0.014037f
C372 VTAIL.n161 VSUBS 0.031336f
C373 VTAIL.n162 VSUBS 0.031336f
C374 VTAIL.n163 VSUBS 0.014037f
C375 VTAIL.n164 VSUBS 0.013257f
C376 VTAIL.n165 VSUBS 0.024672f
C377 VTAIL.n166 VSUBS 0.024672f
C378 VTAIL.n167 VSUBS 0.013257f
C379 VTAIL.n168 VSUBS 0.014037f
C380 VTAIL.n169 VSUBS 0.031336f
C381 VTAIL.n170 VSUBS 0.078003f
C382 VTAIL.n171 VSUBS 0.014037f
C383 VTAIL.n172 VSUBS 0.013257f
C384 VTAIL.n173 VSUBS 0.055342f
C385 VTAIL.n174 VSUBS 0.03927f
C386 VTAIL.n175 VSUBS 1.17628f
C387 VP.t1 VSUBS 2.69361f
C388 VP.t0 VSUBS 3.36959f
C389 VP.n0 VSUBS 4.13296f
C390 B.n0 VSUBS 0.006145f
C391 B.n1 VSUBS 0.006145f
C392 B.n2 VSUBS 0.009088f
C393 B.n3 VSUBS 0.006965f
C394 B.n4 VSUBS 0.006965f
C395 B.n5 VSUBS 0.006965f
C396 B.n6 VSUBS 0.006965f
C397 B.n7 VSUBS 0.006965f
C398 B.n8 VSUBS 0.006965f
C399 B.n9 VSUBS 0.006965f
C400 B.n10 VSUBS 0.006965f
C401 B.n11 VSUBS 0.006965f
C402 B.n12 VSUBS 0.006965f
C403 B.n13 VSUBS 0.006965f
C404 B.n14 VSUBS 0.006965f
C405 B.n15 VSUBS 0.01709f
C406 B.n16 VSUBS 0.006965f
C407 B.n17 VSUBS 0.006965f
C408 B.n18 VSUBS 0.006965f
C409 B.n19 VSUBS 0.006965f
C410 B.n20 VSUBS 0.006965f
C411 B.n21 VSUBS 0.006965f
C412 B.n22 VSUBS 0.006965f
C413 B.n23 VSUBS 0.006965f
C414 B.n24 VSUBS 0.006965f
C415 B.n25 VSUBS 0.006965f
C416 B.n26 VSUBS 0.006965f
C417 B.n27 VSUBS 0.006965f
C418 B.n28 VSUBS 0.006965f
C419 B.n29 VSUBS 0.006965f
C420 B.t4 VSUBS 0.128357f
C421 B.t5 VSUBS 0.15886f
C422 B.t3 VSUBS 1.06502f
C423 B.n30 VSUBS 0.261725f
C424 B.n31 VSUBS 0.193138f
C425 B.n32 VSUBS 0.016136f
C426 B.n33 VSUBS 0.006965f
C427 B.n34 VSUBS 0.006965f
C428 B.n35 VSUBS 0.006965f
C429 B.n36 VSUBS 0.006965f
C430 B.n37 VSUBS 0.006965f
C431 B.t1 VSUBS 0.128359f
C432 B.t2 VSUBS 0.158862f
C433 B.t0 VSUBS 1.06502f
C434 B.n38 VSUBS 0.261723f
C435 B.n39 VSUBS 0.193136f
C436 B.n40 VSUBS 0.006965f
C437 B.n41 VSUBS 0.006965f
C438 B.n42 VSUBS 0.006965f
C439 B.n43 VSUBS 0.006965f
C440 B.n44 VSUBS 0.006965f
C441 B.n45 VSUBS 0.006965f
C442 B.n46 VSUBS 0.006965f
C443 B.n47 VSUBS 0.006965f
C444 B.n48 VSUBS 0.006965f
C445 B.n49 VSUBS 0.006965f
C446 B.n50 VSUBS 0.006965f
C447 B.n51 VSUBS 0.006965f
C448 B.n52 VSUBS 0.006965f
C449 B.n53 VSUBS 0.006965f
C450 B.n54 VSUBS 0.01709f
C451 B.n55 VSUBS 0.006965f
C452 B.n56 VSUBS 0.006965f
C453 B.n57 VSUBS 0.006965f
C454 B.n58 VSUBS 0.006965f
C455 B.n59 VSUBS 0.006965f
C456 B.n60 VSUBS 0.006965f
C457 B.n61 VSUBS 0.006965f
C458 B.n62 VSUBS 0.006965f
C459 B.n63 VSUBS 0.006965f
C460 B.n64 VSUBS 0.006965f
C461 B.n65 VSUBS 0.006965f
C462 B.n66 VSUBS 0.006965f
C463 B.n67 VSUBS 0.006965f
C464 B.n68 VSUBS 0.006965f
C465 B.n69 VSUBS 0.006965f
C466 B.n70 VSUBS 0.006965f
C467 B.n71 VSUBS 0.006965f
C468 B.n72 VSUBS 0.006965f
C469 B.n73 VSUBS 0.006965f
C470 B.n74 VSUBS 0.006965f
C471 B.n75 VSUBS 0.006965f
C472 B.n76 VSUBS 0.006965f
C473 B.n77 VSUBS 0.006965f
C474 B.n78 VSUBS 0.006965f
C475 B.n79 VSUBS 0.006965f
C476 B.n80 VSUBS 0.006965f
C477 B.n81 VSUBS 0.016094f
C478 B.n82 VSUBS 0.006965f
C479 B.n83 VSUBS 0.006965f
C480 B.n84 VSUBS 0.006965f
C481 B.n85 VSUBS 0.006965f
C482 B.n86 VSUBS 0.006965f
C483 B.n87 VSUBS 0.006965f
C484 B.n88 VSUBS 0.006965f
C485 B.n89 VSUBS 0.006965f
C486 B.n90 VSUBS 0.006965f
C487 B.n91 VSUBS 0.006965f
C488 B.n92 VSUBS 0.006965f
C489 B.n93 VSUBS 0.006965f
C490 B.n94 VSUBS 0.006965f
C491 B.n95 VSUBS 0.006965f
C492 B.n96 VSUBS 0.006555f
C493 B.n97 VSUBS 0.006965f
C494 B.n98 VSUBS 0.006965f
C495 B.n99 VSUBS 0.006965f
C496 B.n100 VSUBS 0.006965f
C497 B.n101 VSUBS 0.006965f
C498 B.t8 VSUBS 0.128357f
C499 B.t7 VSUBS 0.15886f
C500 B.t6 VSUBS 1.06502f
C501 B.n102 VSUBS 0.261725f
C502 B.n103 VSUBS 0.193138f
C503 B.n104 VSUBS 0.006965f
C504 B.n105 VSUBS 0.006965f
C505 B.n106 VSUBS 0.006965f
C506 B.n107 VSUBS 0.006965f
C507 B.n108 VSUBS 0.006965f
C508 B.n109 VSUBS 0.006965f
C509 B.n110 VSUBS 0.006965f
C510 B.n111 VSUBS 0.006965f
C511 B.n112 VSUBS 0.006965f
C512 B.n113 VSUBS 0.006965f
C513 B.n114 VSUBS 0.006965f
C514 B.n115 VSUBS 0.006965f
C515 B.n116 VSUBS 0.006965f
C516 B.n117 VSUBS 0.006965f
C517 B.n118 VSUBS 0.01709f
C518 B.n119 VSUBS 0.006965f
C519 B.n120 VSUBS 0.006965f
C520 B.n121 VSUBS 0.006965f
C521 B.n122 VSUBS 0.006965f
C522 B.n123 VSUBS 0.006965f
C523 B.n124 VSUBS 0.006965f
C524 B.n125 VSUBS 0.006965f
C525 B.n126 VSUBS 0.006965f
C526 B.n127 VSUBS 0.006965f
C527 B.n128 VSUBS 0.006965f
C528 B.n129 VSUBS 0.006965f
C529 B.n130 VSUBS 0.006965f
C530 B.n131 VSUBS 0.006965f
C531 B.n132 VSUBS 0.006965f
C532 B.n133 VSUBS 0.006965f
C533 B.n134 VSUBS 0.006965f
C534 B.n135 VSUBS 0.006965f
C535 B.n136 VSUBS 0.006965f
C536 B.n137 VSUBS 0.006965f
C537 B.n138 VSUBS 0.006965f
C538 B.n139 VSUBS 0.006965f
C539 B.n140 VSUBS 0.006965f
C540 B.n141 VSUBS 0.006965f
C541 B.n142 VSUBS 0.006965f
C542 B.n143 VSUBS 0.006965f
C543 B.n144 VSUBS 0.006965f
C544 B.n145 VSUBS 0.006965f
C545 B.n146 VSUBS 0.006965f
C546 B.n147 VSUBS 0.006965f
C547 B.n148 VSUBS 0.006965f
C548 B.n149 VSUBS 0.006965f
C549 B.n150 VSUBS 0.006965f
C550 B.n151 VSUBS 0.006965f
C551 B.n152 VSUBS 0.006965f
C552 B.n153 VSUBS 0.006965f
C553 B.n154 VSUBS 0.006965f
C554 B.n155 VSUBS 0.006965f
C555 B.n156 VSUBS 0.006965f
C556 B.n157 VSUBS 0.006965f
C557 B.n158 VSUBS 0.006965f
C558 B.n159 VSUBS 0.006965f
C559 B.n160 VSUBS 0.006965f
C560 B.n161 VSUBS 0.006965f
C561 B.n162 VSUBS 0.006965f
C562 B.n163 VSUBS 0.006965f
C563 B.n164 VSUBS 0.006965f
C564 B.n165 VSUBS 0.006965f
C565 B.n166 VSUBS 0.006965f
C566 B.n167 VSUBS 0.016094f
C567 B.n168 VSUBS 0.016094f
C568 B.n169 VSUBS 0.01709f
C569 B.n170 VSUBS 0.006965f
C570 B.n171 VSUBS 0.006965f
C571 B.n172 VSUBS 0.006965f
C572 B.n173 VSUBS 0.006965f
C573 B.n174 VSUBS 0.006965f
C574 B.n175 VSUBS 0.006965f
C575 B.n176 VSUBS 0.006965f
C576 B.n177 VSUBS 0.006965f
C577 B.n178 VSUBS 0.006965f
C578 B.n179 VSUBS 0.006965f
C579 B.n180 VSUBS 0.006965f
C580 B.n181 VSUBS 0.006965f
C581 B.n182 VSUBS 0.006965f
C582 B.n183 VSUBS 0.006965f
C583 B.n184 VSUBS 0.006965f
C584 B.n185 VSUBS 0.006965f
C585 B.n186 VSUBS 0.006965f
C586 B.n187 VSUBS 0.006965f
C587 B.n188 VSUBS 0.006965f
C588 B.n189 VSUBS 0.006965f
C589 B.n190 VSUBS 0.006965f
C590 B.n191 VSUBS 0.006965f
C591 B.n192 VSUBS 0.006965f
C592 B.n193 VSUBS 0.006965f
C593 B.n194 VSUBS 0.006965f
C594 B.n195 VSUBS 0.006965f
C595 B.n196 VSUBS 0.006965f
C596 B.n197 VSUBS 0.006965f
C597 B.n198 VSUBS 0.006965f
C598 B.n199 VSUBS 0.006965f
C599 B.n200 VSUBS 0.006965f
C600 B.n201 VSUBS 0.006965f
C601 B.n202 VSUBS 0.006965f
C602 B.n203 VSUBS 0.006965f
C603 B.n204 VSUBS 0.006965f
C604 B.n205 VSUBS 0.006965f
C605 B.n206 VSUBS 0.006965f
C606 B.n207 VSUBS 0.006965f
C607 B.n208 VSUBS 0.006965f
C608 B.n209 VSUBS 0.006965f
C609 B.n210 VSUBS 0.006965f
C610 B.n211 VSUBS 0.006965f
C611 B.n212 VSUBS 0.006965f
C612 B.n213 VSUBS 0.006555f
C613 B.n214 VSUBS 0.016136f
C614 B.n215 VSUBS 0.003892f
C615 B.n216 VSUBS 0.006965f
C616 B.n217 VSUBS 0.006965f
C617 B.n218 VSUBS 0.006965f
C618 B.n219 VSUBS 0.006965f
C619 B.n220 VSUBS 0.006965f
C620 B.n221 VSUBS 0.006965f
C621 B.n222 VSUBS 0.006965f
C622 B.n223 VSUBS 0.006965f
C623 B.n224 VSUBS 0.006965f
C624 B.n225 VSUBS 0.006965f
C625 B.n226 VSUBS 0.006965f
C626 B.n227 VSUBS 0.006965f
C627 B.t11 VSUBS 0.128359f
C628 B.t10 VSUBS 0.158862f
C629 B.t9 VSUBS 1.06502f
C630 B.n228 VSUBS 0.261723f
C631 B.n229 VSUBS 0.193136f
C632 B.n230 VSUBS 0.016136f
C633 B.n231 VSUBS 0.003892f
C634 B.n232 VSUBS 0.006965f
C635 B.n233 VSUBS 0.006965f
C636 B.n234 VSUBS 0.006965f
C637 B.n235 VSUBS 0.006965f
C638 B.n236 VSUBS 0.006965f
C639 B.n237 VSUBS 0.006965f
C640 B.n238 VSUBS 0.006965f
C641 B.n239 VSUBS 0.006965f
C642 B.n240 VSUBS 0.006965f
C643 B.n241 VSUBS 0.006965f
C644 B.n242 VSUBS 0.006965f
C645 B.n243 VSUBS 0.006965f
C646 B.n244 VSUBS 0.006965f
C647 B.n245 VSUBS 0.006965f
C648 B.n246 VSUBS 0.006965f
C649 B.n247 VSUBS 0.006965f
C650 B.n248 VSUBS 0.006965f
C651 B.n249 VSUBS 0.006965f
C652 B.n250 VSUBS 0.006965f
C653 B.n251 VSUBS 0.006965f
C654 B.n252 VSUBS 0.006965f
C655 B.n253 VSUBS 0.006965f
C656 B.n254 VSUBS 0.006965f
C657 B.n255 VSUBS 0.006965f
C658 B.n256 VSUBS 0.006965f
C659 B.n257 VSUBS 0.006965f
C660 B.n258 VSUBS 0.006965f
C661 B.n259 VSUBS 0.006965f
C662 B.n260 VSUBS 0.006965f
C663 B.n261 VSUBS 0.006965f
C664 B.n262 VSUBS 0.006965f
C665 B.n263 VSUBS 0.006965f
C666 B.n264 VSUBS 0.006965f
C667 B.n265 VSUBS 0.006965f
C668 B.n266 VSUBS 0.006965f
C669 B.n267 VSUBS 0.006965f
C670 B.n268 VSUBS 0.006965f
C671 B.n269 VSUBS 0.006965f
C672 B.n270 VSUBS 0.006965f
C673 B.n271 VSUBS 0.006965f
C674 B.n272 VSUBS 0.006965f
C675 B.n273 VSUBS 0.006965f
C676 B.n274 VSUBS 0.006965f
C677 B.n275 VSUBS 0.006965f
C678 B.n276 VSUBS 0.01709f
C679 B.n277 VSUBS 0.016289f
C680 B.n278 VSUBS 0.016895f
C681 B.n279 VSUBS 0.006965f
C682 B.n280 VSUBS 0.006965f
C683 B.n281 VSUBS 0.006965f
C684 B.n282 VSUBS 0.006965f
C685 B.n283 VSUBS 0.006965f
C686 B.n284 VSUBS 0.006965f
C687 B.n285 VSUBS 0.006965f
C688 B.n286 VSUBS 0.006965f
C689 B.n287 VSUBS 0.006965f
C690 B.n288 VSUBS 0.006965f
C691 B.n289 VSUBS 0.006965f
C692 B.n290 VSUBS 0.006965f
C693 B.n291 VSUBS 0.006965f
C694 B.n292 VSUBS 0.006965f
C695 B.n293 VSUBS 0.006965f
C696 B.n294 VSUBS 0.006965f
C697 B.n295 VSUBS 0.006965f
C698 B.n296 VSUBS 0.006965f
C699 B.n297 VSUBS 0.006965f
C700 B.n298 VSUBS 0.006965f
C701 B.n299 VSUBS 0.006965f
C702 B.n300 VSUBS 0.006965f
C703 B.n301 VSUBS 0.006965f
C704 B.n302 VSUBS 0.006965f
C705 B.n303 VSUBS 0.006965f
C706 B.n304 VSUBS 0.006965f
C707 B.n305 VSUBS 0.006965f
C708 B.n306 VSUBS 0.006965f
C709 B.n307 VSUBS 0.006965f
C710 B.n308 VSUBS 0.006965f
C711 B.n309 VSUBS 0.006965f
C712 B.n310 VSUBS 0.006965f
C713 B.n311 VSUBS 0.006965f
C714 B.n312 VSUBS 0.006965f
C715 B.n313 VSUBS 0.006965f
C716 B.n314 VSUBS 0.006965f
C717 B.n315 VSUBS 0.006965f
C718 B.n316 VSUBS 0.006965f
C719 B.n317 VSUBS 0.006965f
C720 B.n318 VSUBS 0.006965f
C721 B.n319 VSUBS 0.006965f
C722 B.n320 VSUBS 0.006965f
C723 B.n321 VSUBS 0.006965f
C724 B.n322 VSUBS 0.006965f
C725 B.n323 VSUBS 0.006965f
C726 B.n324 VSUBS 0.006965f
C727 B.n325 VSUBS 0.006965f
C728 B.n326 VSUBS 0.006965f
C729 B.n327 VSUBS 0.006965f
C730 B.n328 VSUBS 0.006965f
C731 B.n329 VSUBS 0.006965f
C732 B.n330 VSUBS 0.006965f
C733 B.n331 VSUBS 0.006965f
C734 B.n332 VSUBS 0.006965f
C735 B.n333 VSUBS 0.006965f
C736 B.n334 VSUBS 0.006965f
C737 B.n335 VSUBS 0.006965f
C738 B.n336 VSUBS 0.006965f
C739 B.n337 VSUBS 0.006965f
C740 B.n338 VSUBS 0.006965f
C741 B.n339 VSUBS 0.006965f
C742 B.n340 VSUBS 0.006965f
C743 B.n341 VSUBS 0.006965f
C744 B.n342 VSUBS 0.006965f
C745 B.n343 VSUBS 0.006965f
C746 B.n344 VSUBS 0.006965f
C747 B.n345 VSUBS 0.006965f
C748 B.n346 VSUBS 0.006965f
C749 B.n347 VSUBS 0.006965f
C750 B.n348 VSUBS 0.006965f
C751 B.n349 VSUBS 0.006965f
C752 B.n350 VSUBS 0.006965f
C753 B.n351 VSUBS 0.006965f
C754 B.n352 VSUBS 0.006965f
C755 B.n353 VSUBS 0.006965f
C756 B.n354 VSUBS 0.006965f
C757 B.n355 VSUBS 0.006965f
C758 B.n356 VSUBS 0.006965f
C759 B.n357 VSUBS 0.016094f
C760 B.n358 VSUBS 0.016094f
C761 B.n359 VSUBS 0.01709f
C762 B.n360 VSUBS 0.006965f
C763 B.n361 VSUBS 0.006965f
C764 B.n362 VSUBS 0.006965f
C765 B.n363 VSUBS 0.006965f
C766 B.n364 VSUBS 0.006965f
C767 B.n365 VSUBS 0.006965f
C768 B.n366 VSUBS 0.006965f
C769 B.n367 VSUBS 0.006965f
C770 B.n368 VSUBS 0.006965f
C771 B.n369 VSUBS 0.006965f
C772 B.n370 VSUBS 0.006965f
C773 B.n371 VSUBS 0.006965f
C774 B.n372 VSUBS 0.006965f
C775 B.n373 VSUBS 0.006965f
C776 B.n374 VSUBS 0.006965f
C777 B.n375 VSUBS 0.006965f
C778 B.n376 VSUBS 0.006965f
C779 B.n377 VSUBS 0.006965f
C780 B.n378 VSUBS 0.006965f
C781 B.n379 VSUBS 0.006965f
C782 B.n380 VSUBS 0.006965f
C783 B.n381 VSUBS 0.006965f
C784 B.n382 VSUBS 0.006965f
C785 B.n383 VSUBS 0.006965f
C786 B.n384 VSUBS 0.006965f
C787 B.n385 VSUBS 0.006965f
C788 B.n386 VSUBS 0.006965f
C789 B.n387 VSUBS 0.006965f
C790 B.n388 VSUBS 0.006965f
C791 B.n389 VSUBS 0.006965f
C792 B.n390 VSUBS 0.006965f
C793 B.n391 VSUBS 0.006965f
C794 B.n392 VSUBS 0.006965f
C795 B.n393 VSUBS 0.006965f
C796 B.n394 VSUBS 0.006965f
C797 B.n395 VSUBS 0.006965f
C798 B.n396 VSUBS 0.006965f
C799 B.n397 VSUBS 0.006965f
C800 B.n398 VSUBS 0.006965f
C801 B.n399 VSUBS 0.006965f
C802 B.n400 VSUBS 0.006965f
C803 B.n401 VSUBS 0.006965f
C804 B.n402 VSUBS 0.006965f
C805 B.n403 VSUBS 0.006555f
C806 B.n404 VSUBS 0.016136f
C807 B.n405 VSUBS 0.003892f
C808 B.n406 VSUBS 0.006965f
C809 B.n407 VSUBS 0.006965f
C810 B.n408 VSUBS 0.006965f
C811 B.n409 VSUBS 0.006965f
C812 B.n410 VSUBS 0.006965f
C813 B.n411 VSUBS 0.006965f
C814 B.n412 VSUBS 0.006965f
C815 B.n413 VSUBS 0.006965f
C816 B.n414 VSUBS 0.006965f
C817 B.n415 VSUBS 0.006965f
C818 B.n416 VSUBS 0.006965f
C819 B.n417 VSUBS 0.006965f
C820 B.n418 VSUBS 0.003892f
C821 B.n419 VSUBS 0.006965f
C822 B.n420 VSUBS 0.006965f
C823 B.n421 VSUBS 0.006555f
C824 B.n422 VSUBS 0.006965f
C825 B.n423 VSUBS 0.006965f
C826 B.n424 VSUBS 0.006965f
C827 B.n425 VSUBS 0.006965f
C828 B.n426 VSUBS 0.006965f
C829 B.n427 VSUBS 0.006965f
C830 B.n428 VSUBS 0.006965f
C831 B.n429 VSUBS 0.006965f
C832 B.n430 VSUBS 0.006965f
C833 B.n431 VSUBS 0.006965f
C834 B.n432 VSUBS 0.006965f
C835 B.n433 VSUBS 0.006965f
C836 B.n434 VSUBS 0.006965f
C837 B.n435 VSUBS 0.006965f
C838 B.n436 VSUBS 0.006965f
C839 B.n437 VSUBS 0.006965f
C840 B.n438 VSUBS 0.006965f
C841 B.n439 VSUBS 0.006965f
C842 B.n440 VSUBS 0.006965f
C843 B.n441 VSUBS 0.006965f
C844 B.n442 VSUBS 0.006965f
C845 B.n443 VSUBS 0.006965f
C846 B.n444 VSUBS 0.006965f
C847 B.n445 VSUBS 0.006965f
C848 B.n446 VSUBS 0.006965f
C849 B.n447 VSUBS 0.006965f
C850 B.n448 VSUBS 0.006965f
C851 B.n449 VSUBS 0.006965f
C852 B.n450 VSUBS 0.006965f
C853 B.n451 VSUBS 0.006965f
C854 B.n452 VSUBS 0.006965f
C855 B.n453 VSUBS 0.006965f
C856 B.n454 VSUBS 0.006965f
C857 B.n455 VSUBS 0.006965f
C858 B.n456 VSUBS 0.006965f
C859 B.n457 VSUBS 0.006965f
C860 B.n458 VSUBS 0.006965f
C861 B.n459 VSUBS 0.006965f
C862 B.n460 VSUBS 0.006965f
C863 B.n461 VSUBS 0.006965f
C864 B.n462 VSUBS 0.006965f
C865 B.n463 VSUBS 0.006965f
C866 B.n464 VSUBS 0.01709f
C867 B.n465 VSUBS 0.016094f
C868 B.n466 VSUBS 0.016094f
C869 B.n467 VSUBS 0.006965f
C870 B.n468 VSUBS 0.006965f
C871 B.n469 VSUBS 0.006965f
C872 B.n470 VSUBS 0.006965f
C873 B.n471 VSUBS 0.006965f
C874 B.n472 VSUBS 0.006965f
C875 B.n473 VSUBS 0.006965f
C876 B.n474 VSUBS 0.006965f
C877 B.n475 VSUBS 0.006965f
C878 B.n476 VSUBS 0.006965f
C879 B.n477 VSUBS 0.006965f
C880 B.n478 VSUBS 0.006965f
C881 B.n479 VSUBS 0.006965f
C882 B.n480 VSUBS 0.006965f
C883 B.n481 VSUBS 0.006965f
C884 B.n482 VSUBS 0.006965f
C885 B.n483 VSUBS 0.006965f
C886 B.n484 VSUBS 0.006965f
C887 B.n485 VSUBS 0.006965f
C888 B.n486 VSUBS 0.006965f
C889 B.n487 VSUBS 0.006965f
C890 B.n488 VSUBS 0.006965f
C891 B.n489 VSUBS 0.006965f
C892 B.n490 VSUBS 0.006965f
C893 B.n491 VSUBS 0.006965f
C894 B.n492 VSUBS 0.006965f
C895 B.n493 VSUBS 0.006965f
C896 B.n494 VSUBS 0.006965f
C897 B.n495 VSUBS 0.006965f
C898 B.n496 VSUBS 0.006965f
C899 B.n497 VSUBS 0.006965f
C900 B.n498 VSUBS 0.006965f
C901 B.n499 VSUBS 0.006965f
C902 B.n500 VSUBS 0.006965f
C903 B.n501 VSUBS 0.006965f
C904 B.n502 VSUBS 0.006965f
C905 B.n503 VSUBS 0.009088f
C906 B.n504 VSUBS 0.009682f
C907 B.n505 VSUBS 0.019253f
.ends

