* NGSPICE file created from diff_pair_sample_0376.ext - technology: sky130A

.subckt diff_pair_sample_0376 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t10 VN.t0 VDD2.t1 w_n3810_n3168# sky130_fd_pr__pfet_01v8 ad=1.815 pd=11.33 as=1.815 ps=11.33 w=11 l=3.22
X1 VDD1.t5 VP.t0 VTAIL.t2 w_n3810_n3168# sky130_fd_pr__pfet_01v8 ad=4.29 pd=22.78 as=1.815 ps=11.33 w=11 l=3.22
X2 B.t11 B.t9 B.t10 w_n3810_n3168# sky130_fd_pr__pfet_01v8 ad=4.29 pd=22.78 as=0 ps=0 w=11 l=3.22
X3 B.t8 B.t6 B.t7 w_n3810_n3168# sky130_fd_pr__pfet_01v8 ad=4.29 pd=22.78 as=0 ps=0 w=11 l=3.22
X4 VDD2.t4 VN.t1 VTAIL.t9 w_n3810_n3168# sky130_fd_pr__pfet_01v8 ad=1.815 pd=11.33 as=4.29 ps=22.78 w=11 l=3.22
X5 VDD1.t4 VP.t1 VTAIL.t3 w_n3810_n3168# sky130_fd_pr__pfet_01v8 ad=1.815 pd=11.33 as=4.29 ps=22.78 w=11 l=3.22
X6 VDD1.t3 VP.t2 VTAIL.t1 w_n3810_n3168# sky130_fd_pr__pfet_01v8 ad=4.29 pd=22.78 as=1.815 ps=11.33 w=11 l=3.22
X7 B.t5 B.t3 B.t4 w_n3810_n3168# sky130_fd_pr__pfet_01v8 ad=4.29 pd=22.78 as=0 ps=0 w=11 l=3.22
X8 VDD2.t0 VN.t2 VTAIL.t8 w_n3810_n3168# sky130_fd_pr__pfet_01v8 ad=1.815 pd=11.33 as=4.29 ps=22.78 w=11 l=3.22
X9 VTAIL.t4 VP.t3 VDD1.t2 w_n3810_n3168# sky130_fd_pr__pfet_01v8 ad=1.815 pd=11.33 as=1.815 ps=11.33 w=11 l=3.22
X10 VDD1.t1 VP.t4 VTAIL.t11 w_n3810_n3168# sky130_fd_pr__pfet_01v8 ad=1.815 pd=11.33 as=4.29 ps=22.78 w=11 l=3.22
X11 B.t2 B.t0 B.t1 w_n3810_n3168# sky130_fd_pr__pfet_01v8 ad=4.29 pd=22.78 as=0 ps=0 w=11 l=3.22
X12 VTAIL.t0 VP.t5 VDD1.t0 w_n3810_n3168# sky130_fd_pr__pfet_01v8 ad=1.815 pd=11.33 as=1.815 ps=11.33 w=11 l=3.22
X13 VDD2.t2 VN.t3 VTAIL.t7 w_n3810_n3168# sky130_fd_pr__pfet_01v8 ad=4.29 pd=22.78 as=1.815 ps=11.33 w=11 l=3.22
X14 VDD2.t5 VN.t4 VTAIL.t6 w_n3810_n3168# sky130_fd_pr__pfet_01v8 ad=4.29 pd=22.78 as=1.815 ps=11.33 w=11 l=3.22
X15 VTAIL.t5 VN.t5 VDD2.t3 w_n3810_n3168# sky130_fd_pr__pfet_01v8 ad=1.815 pd=11.33 as=1.815 ps=11.33 w=11 l=3.22
R0 VN.n34 VN.n33 161.3
R1 VN.n32 VN.n19 161.3
R2 VN.n31 VN.n30 161.3
R3 VN.n29 VN.n20 161.3
R4 VN.n28 VN.n27 161.3
R5 VN.n26 VN.n21 161.3
R6 VN.n25 VN.n24 161.3
R7 VN.n16 VN.n15 161.3
R8 VN.n14 VN.n1 161.3
R9 VN.n13 VN.n12 161.3
R10 VN.n11 VN.n2 161.3
R11 VN.n10 VN.n9 161.3
R12 VN.n8 VN.n3 161.3
R13 VN.n7 VN.n6 161.3
R14 VN.n5 VN.t4 115.365
R15 VN.n23 VN.t2 115.365
R16 VN.n4 VN.t5 82.3297
R17 VN.n0 VN.t1 82.3297
R18 VN.n22 VN.t0 82.3297
R19 VN.n18 VN.t3 82.3297
R20 VN.n17 VN.n0 75.4905
R21 VN.n35 VN.n18 75.4905
R22 VN.n23 VN.n22 62.2128
R23 VN.n5 VN.n4 62.2128
R24 VN VN.n35 50.608
R25 VN.n13 VN.n2 42.999
R26 VN.n31 VN.n20 42.999
R27 VN.n9 VN.n2 38.1551
R28 VN.n27 VN.n20 38.1551
R29 VN.n8 VN.n7 24.5923
R30 VN.n9 VN.n8 24.5923
R31 VN.n14 VN.n13 24.5923
R32 VN.n15 VN.n14 24.5923
R33 VN.n27 VN.n26 24.5923
R34 VN.n26 VN.n25 24.5923
R35 VN.n33 VN.n32 24.5923
R36 VN.n32 VN.n31 24.5923
R37 VN.n15 VN.n0 14.7556
R38 VN.n33 VN.n18 14.7556
R39 VN.n7 VN.n4 12.2964
R40 VN.n25 VN.n22 12.2964
R41 VN.n6 VN.n5 4.14385
R42 VN.n24 VN.n23 4.14385
R43 VN.n35 VN.n34 0.354861
R44 VN.n17 VN.n16 0.354861
R45 VN VN.n17 0.267071
R46 VN.n34 VN.n19 0.189894
R47 VN.n30 VN.n19 0.189894
R48 VN.n30 VN.n29 0.189894
R49 VN.n29 VN.n28 0.189894
R50 VN.n28 VN.n21 0.189894
R51 VN.n24 VN.n21 0.189894
R52 VN.n6 VN.n3 0.189894
R53 VN.n10 VN.n3 0.189894
R54 VN.n11 VN.n10 0.189894
R55 VN.n12 VN.n11 0.189894
R56 VN.n12 VN.n1 0.189894
R57 VN.n16 VN.n1 0.189894
R58 VDD2.n1 VDD2.t5 79.724
R59 VDD2.n2 VDD2.t2 77.4842
R60 VDD2.n1 VDD2.n0 75.2388
R61 VDD2 VDD2.n3 75.236
R62 VDD2.n2 VDD2.n1 43.1442
R63 VDD2.n3 VDD2.t1 2.9555
R64 VDD2.n3 VDD2.t0 2.9555
R65 VDD2.n0 VDD2.t3 2.9555
R66 VDD2.n0 VDD2.t4 2.9555
R67 VDD2 VDD2.n2 2.35395
R68 VTAIL.n7 VTAIL.t8 60.8054
R69 VTAIL.n11 VTAIL.t9 60.8053
R70 VTAIL.n2 VTAIL.t3 60.8053
R71 VTAIL.n10 VTAIL.t11 60.8053
R72 VTAIL.n9 VTAIL.n8 57.8505
R73 VTAIL.n6 VTAIL.n5 57.8505
R74 VTAIL.n1 VTAIL.n0 57.8503
R75 VTAIL.n4 VTAIL.n3 57.8503
R76 VTAIL.n6 VTAIL.n4 27.9703
R77 VTAIL.n11 VTAIL.n10 24.91
R78 VTAIL.n7 VTAIL.n6 3.06084
R79 VTAIL.n10 VTAIL.n9 3.06084
R80 VTAIL.n4 VTAIL.n2 3.06084
R81 VTAIL.n0 VTAIL.t6 2.9555
R82 VTAIL.n0 VTAIL.t5 2.9555
R83 VTAIL.n3 VTAIL.t1 2.9555
R84 VTAIL.n3 VTAIL.t4 2.9555
R85 VTAIL.n8 VTAIL.t2 2.9555
R86 VTAIL.n8 VTAIL.t0 2.9555
R87 VTAIL.n5 VTAIL.t7 2.9555
R88 VTAIL.n5 VTAIL.t10 2.9555
R89 VTAIL VTAIL.n11 2.23757
R90 VTAIL.n9 VTAIL.n7 2.0005
R91 VTAIL.n2 VTAIL.n1 2.0005
R92 VTAIL VTAIL.n1 0.823776
R93 VP.n16 VP.n15 161.3
R94 VP.n17 VP.n12 161.3
R95 VP.n19 VP.n18 161.3
R96 VP.n20 VP.n11 161.3
R97 VP.n22 VP.n21 161.3
R98 VP.n23 VP.n10 161.3
R99 VP.n25 VP.n24 161.3
R100 VP.n49 VP.n48 161.3
R101 VP.n47 VP.n1 161.3
R102 VP.n46 VP.n45 161.3
R103 VP.n44 VP.n2 161.3
R104 VP.n43 VP.n42 161.3
R105 VP.n41 VP.n3 161.3
R106 VP.n40 VP.n39 161.3
R107 VP.n38 VP.n37 161.3
R108 VP.n36 VP.n5 161.3
R109 VP.n35 VP.n34 161.3
R110 VP.n33 VP.n6 161.3
R111 VP.n32 VP.n31 161.3
R112 VP.n30 VP.n7 161.3
R113 VP.n29 VP.n28 161.3
R114 VP.n14 VP.t0 115.365
R115 VP.n8 VP.t2 82.3297
R116 VP.n4 VP.t3 82.3297
R117 VP.n0 VP.t1 82.3297
R118 VP.n9 VP.t4 82.3297
R119 VP.n13 VP.t5 82.3297
R120 VP.n27 VP.n8 75.4905
R121 VP.n50 VP.n0 75.4905
R122 VP.n26 VP.n9 75.4905
R123 VP.n14 VP.n13 62.2128
R124 VP.n27 VP.n26 50.4427
R125 VP.n31 VP.n6 42.999
R126 VP.n46 VP.n2 42.999
R127 VP.n22 VP.n11 42.999
R128 VP.n35 VP.n6 38.1551
R129 VP.n42 VP.n2 38.1551
R130 VP.n18 VP.n11 38.1551
R131 VP.n30 VP.n29 24.5923
R132 VP.n31 VP.n30 24.5923
R133 VP.n36 VP.n35 24.5923
R134 VP.n37 VP.n36 24.5923
R135 VP.n41 VP.n40 24.5923
R136 VP.n42 VP.n41 24.5923
R137 VP.n47 VP.n46 24.5923
R138 VP.n48 VP.n47 24.5923
R139 VP.n23 VP.n22 24.5923
R140 VP.n24 VP.n23 24.5923
R141 VP.n17 VP.n16 24.5923
R142 VP.n18 VP.n17 24.5923
R143 VP.n29 VP.n8 14.7556
R144 VP.n48 VP.n0 14.7556
R145 VP.n24 VP.n9 14.7556
R146 VP.n37 VP.n4 12.2964
R147 VP.n40 VP.n4 12.2964
R148 VP.n16 VP.n13 12.2964
R149 VP.n15 VP.n14 4.14382
R150 VP.n26 VP.n25 0.354861
R151 VP.n28 VP.n27 0.354861
R152 VP.n50 VP.n49 0.354861
R153 VP VP.n50 0.267071
R154 VP.n15 VP.n12 0.189894
R155 VP.n19 VP.n12 0.189894
R156 VP.n20 VP.n19 0.189894
R157 VP.n21 VP.n20 0.189894
R158 VP.n21 VP.n10 0.189894
R159 VP.n25 VP.n10 0.189894
R160 VP.n28 VP.n7 0.189894
R161 VP.n32 VP.n7 0.189894
R162 VP.n33 VP.n32 0.189894
R163 VP.n34 VP.n33 0.189894
R164 VP.n34 VP.n5 0.189894
R165 VP.n38 VP.n5 0.189894
R166 VP.n39 VP.n38 0.189894
R167 VP.n39 VP.n3 0.189894
R168 VP.n43 VP.n3 0.189894
R169 VP.n44 VP.n43 0.189894
R170 VP.n45 VP.n44 0.189894
R171 VP.n45 VP.n1 0.189894
R172 VP.n49 VP.n1 0.189894
R173 VDD1 VDD1.t5 79.8377
R174 VDD1.n1 VDD1.t3 79.724
R175 VDD1.n1 VDD1.n0 75.2388
R176 VDD1.n3 VDD1.n2 74.5291
R177 VDD1.n3 VDD1.n1 45.2574
R178 VDD1.n2 VDD1.t0 2.9555
R179 VDD1.n2 VDD1.t1 2.9555
R180 VDD1.n0 VDD1.t2 2.9555
R181 VDD1.n0 VDD1.t4 2.9555
R182 VDD1 VDD1.n3 0.707397
R183 B.n556 B.n75 585
R184 B.n558 B.n557 585
R185 B.n559 B.n74 585
R186 B.n561 B.n560 585
R187 B.n562 B.n73 585
R188 B.n564 B.n563 585
R189 B.n565 B.n72 585
R190 B.n567 B.n566 585
R191 B.n568 B.n71 585
R192 B.n570 B.n569 585
R193 B.n571 B.n70 585
R194 B.n573 B.n572 585
R195 B.n574 B.n69 585
R196 B.n576 B.n575 585
R197 B.n577 B.n68 585
R198 B.n579 B.n578 585
R199 B.n580 B.n67 585
R200 B.n582 B.n581 585
R201 B.n583 B.n66 585
R202 B.n585 B.n584 585
R203 B.n586 B.n65 585
R204 B.n588 B.n587 585
R205 B.n589 B.n64 585
R206 B.n591 B.n590 585
R207 B.n592 B.n63 585
R208 B.n594 B.n593 585
R209 B.n595 B.n62 585
R210 B.n597 B.n596 585
R211 B.n598 B.n61 585
R212 B.n600 B.n599 585
R213 B.n601 B.n60 585
R214 B.n603 B.n602 585
R215 B.n604 B.n59 585
R216 B.n606 B.n605 585
R217 B.n607 B.n58 585
R218 B.n609 B.n608 585
R219 B.n610 B.n57 585
R220 B.n612 B.n611 585
R221 B.n613 B.n54 585
R222 B.n616 B.n615 585
R223 B.n617 B.n53 585
R224 B.n619 B.n618 585
R225 B.n620 B.n52 585
R226 B.n622 B.n621 585
R227 B.n623 B.n51 585
R228 B.n625 B.n624 585
R229 B.n626 B.n47 585
R230 B.n628 B.n627 585
R231 B.n629 B.n46 585
R232 B.n631 B.n630 585
R233 B.n632 B.n45 585
R234 B.n634 B.n633 585
R235 B.n635 B.n44 585
R236 B.n637 B.n636 585
R237 B.n638 B.n43 585
R238 B.n640 B.n639 585
R239 B.n641 B.n42 585
R240 B.n643 B.n642 585
R241 B.n644 B.n41 585
R242 B.n646 B.n645 585
R243 B.n647 B.n40 585
R244 B.n649 B.n648 585
R245 B.n650 B.n39 585
R246 B.n652 B.n651 585
R247 B.n653 B.n38 585
R248 B.n655 B.n654 585
R249 B.n656 B.n37 585
R250 B.n658 B.n657 585
R251 B.n659 B.n36 585
R252 B.n661 B.n660 585
R253 B.n662 B.n35 585
R254 B.n664 B.n663 585
R255 B.n665 B.n34 585
R256 B.n667 B.n666 585
R257 B.n668 B.n33 585
R258 B.n670 B.n669 585
R259 B.n671 B.n32 585
R260 B.n673 B.n672 585
R261 B.n674 B.n31 585
R262 B.n676 B.n675 585
R263 B.n677 B.n30 585
R264 B.n679 B.n678 585
R265 B.n680 B.n29 585
R266 B.n682 B.n681 585
R267 B.n683 B.n28 585
R268 B.n685 B.n684 585
R269 B.n686 B.n27 585
R270 B.n555 B.n554 585
R271 B.n553 B.n76 585
R272 B.n552 B.n551 585
R273 B.n550 B.n77 585
R274 B.n549 B.n548 585
R275 B.n547 B.n78 585
R276 B.n546 B.n545 585
R277 B.n544 B.n79 585
R278 B.n543 B.n542 585
R279 B.n541 B.n80 585
R280 B.n540 B.n539 585
R281 B.n538 B.n81 585
R282 B.n537 B.n536 585
R283 B.n535 B.n82 585
R284 B.n534 B.n533 585
R285 B.n532 B.n83 585
R286 B.n531 B.n530 585
R287 B.n529 B.n84 585
R288 B.n528 B.n527 585
R289 B.n526 B.n85 585
R290 B.n525 B.n524 585
R291 B.n523 B.n86 585
R292 B.n522 B.n521 585
R293 B.n520 B.n87 585
R294 B.n519 B.n518 585
R295 B.n517 B.n88 585
R296 B.n516 B.n515 585
R297 B.n514 B.n89 585
R298 B.n513 B.n512 585
R299 B.n511 B.n90 585
R300 B.n510 B.n509 585
R301 B.n508 B.n91 585
R302 B.n507 B.n506 585
R303 B.n505 B.n92 585
R304 B.n504 B.n503 585
R305 B.n502 B.n93 585
R306 B.n501 B.n500 585
R307 B.n499 B.n94 585
R308 B.n498 B.n497 585
R309 B.n496 B.n95 585
R310 B.n495 B.n494 585
R311 B.n493 B.n96 585
R312 B.n492 B.n491 585
R313 B.n490 B.n97 585
R314 B.n489 B.n488 585
R315 B.n487 B.n98 585
R316 B.n486 B.n485 585
R317 B.n484 B.n99 585
R318 B.n483 B.n482 585
R319 B.n481 B.n100 585
R320 B.n480 B.n479 585
R321 B.n478 B.n101 585
R322 B.n477 B.n476 585
R323 B.n475 B.n102 585
R324 B.n474 B.n473 585
R325 B.n472 B.n103 585
R326 B.n471 B.n470 585
R327 B.n469 B.n104 585
R328 B.n468 B.n467 585
R329 B.n466 B.n105 585
R330 B.n465 B.n464 585
R331 B.n463 B.n106 585
R332 B.n462 B.n461 585
R333 B.n460 B.n107 585
R334 B.n459 B.n458 585
R335 B.n457 B.n108 585
R336 B.n456 B.n455 585
R337 B.n454 B.n109 585
R338 B.n453 B.n452 585
R339 B.n451 B.n110 585
R340 B.n450 B.n449 585
R341 B.n448 B.n111 585
R342 B.n447 B.n446 585
R343 B.n445 B.n112 585
R344 B.n444 B.n443 585
R345 B.n442 B.n113 585
R346 B.n441 B.n440 585
R347 B.n439 B.n114 585
R348 B.n438 B.n437 585
R349 B.n436 B.n115 585
R350 B.n435 B.n434 585
R351 B.n433 B.n116 585
R352 B.n432 B.n431 585
R353 B.n430 B.n117 585
R354 B.n429 B.n428 585
R355 B.n427 B.n118 585
R356 B.n426 B.n425 585
R357 B.n424 B.n119 585
R358 B.n423 B.n422 585
R359 B.n421 B.n120 585
R360 B.n420 B.n419 585
R361 B.n418 B.n121 585
R362 B.n417 B.n416 585
R363 B.n415 B.n122 585
R364 B.n414 B.n413 585
R365 B.n412 B.n123 585
R366 B.n411 B.n410 585
R367 B.n409 B.n124 585
R368 B.n408 B.n407 585
R369 B.n406 B.n125 585
R370 B.n405 B.n404 585
R371 B.n270 B.n171 585
R372 B.n272 B.n271 585
R373 B.n273 B.n170 585
R374 B.n275 B.n274 585
R375 B.n276 B.n169 585
R376 B.n278 B.n277 585
R377 B.n279 B.n168 585
R378 B.n281 B.n280 585
R379 B.n282 B.n167 585
R380 B.n284 B.n283 585
R381 B.n285 B.n166 585
R382 B.n287 B.n286 585
R383 B.n288 B.n165 585
R384 B.n290 B.n289 585
R385 B.n291 B.n164 585
R386 B.n293 B.n292 585
R387 B.n294 B.n163 585
R388 B.n296 B.n295 585
R389 B.n297 B.n162 585
R390 B.n299 B.n298 585
R391 B.n300 B.n161 585
R392 B.n302 B.n301 585
R393 B.n303 B.n160 585
R394 B.n305 B.n304 585
R395 B.n306 B.n159 585
R396 B.n308 B.n307 585
R397 B.n309 B.n158 585
R398 B.n311 B.n310 585
R399 B.n312 B.n157 585
R400 B.n314 B.n313 585
R401 B.n315 B.n156 585
R402 B.n317 B.n316 585
R403 B.n318 B.n155 585
R404 B.n320 B.n319 585
R405 B.n321 B.n154 585
R406 B.n323 B.n322 585
R407 B.n324 B.n153 585
R408 B.n326 B.n325 585
R409 B.n327 B.n150 585
R410 B.n330 B.n329 585
R411 B.n331 B.n149 585
R412 B.n333 B.n332 585
R413 B.n334 B.n148 585
R414 B.n336 B.n335 585
R415 B.n337 B.n147 585
R416 B.n339 B.n338 585
R417 B.n340 B.n146 585
R418 B.n345 B.n344 585
R419 B.n346 B.n145 585
R420 B.n348 B.n347 585
R421 B.n349 B.n144 585
R422 B.n351 B.n350 585
R423 B.n352 B.n143 585
R424 B.n354 B.n353 585
R425 B.n355 B.n142 585
R426 B.n357 B.n356 585
R427 B.n358 B.n141 585
R428 B.n360 B.n359 585
R429 B.n361 B.n140 585
R430 B.n363 B.n362 585
R431 B.n364 B.n139 585
R432 B.n366 B.n365 585
R433 B.n367 B.n138 585
R434 B.n369 B.n368 585
R435 B.n370 B.n137 585
R436 B.n372 B.n371 585
R437 B.n373 B.n136 585
R438 B.n375 B.n374 585
R439 B.n376 B.n135 585
R440 B.n378 B.n377 585
R441 B.n379 B.n134 585
R442 B.n381 B.n380 585
R443 B.n382 B.n133 585
R444 B.n384 B.n383 585
R445 B.n385 B.n132 585
R446 B.n387 B.n386 585
R447 B.n388 B.n131 585
R448 B.n390 B.n389 585
R449 B.n391 B.n130 585
R450 B.n393 B.n392 585
R451 B.n394 B.n129 585
R452 B.n396 B.n395 585
R453 B.n397 B.n128 585
R454 B.n399 B.n398 585
R455 B.n400 B.n127 585
R456 B.n402 B.n401 585
R457 B.n403 B.n126 585
R458 B.n269 B.n268 585
R459 B.n267 B.n172 585
R460 B.n266 B.n265 585
R461 B.n264 B.n173 585
R462 B.n263 B.n262 585
R463 B.n261 B.n174 585
R464 B.n260 B.n259 585
R465 B.n258 B.n175 585
R466 B.n257 B.n256 585
R467 B.n255 B.n176 585
R468 B.n254 B.n253 585
R469 B.n252 B.n177 585
R470 B.n251 B.n250 585
R471 B.n249 B.n178 585
R472 B.n248 B.n247 585
R473 B.n246 B.n179 585
R474 B.n245 B.n244 585
R475 B.n243 B.n180 585
R476 B.n242 B.n241 585
R477 B.n240 B.n181 585
R478 B.n239 B.n238 585
R479 B.n237 B.n182 585
R480 B.n236 B.n235 585
R481 B.n234 B.n183 585
R482 B.n233 B.n232 585
R483 B.n231 B.n184 585
R484 B.n230 B.n229 585
R485 B.n228 B.n185 585
R486 B.n227 B.n226 585
R487 B.n225 B.n186 585
R488 B.n224 B.n223 585
R489 B.n222 B.n187 585
R490 B.n221 B.n220 585
R491 B.n219 B.n188 585
R492 B.n218 B.n217 585
R493 B.n216 B.n189 585
R494 B.n215 B.n214 585
R495 B.n213 B.n190 585
R496 B.n212 B.n211 585
R497 B.n210 B.n191 585
R498 B.n209 B.n208 585
R499 B.n207 B.n192 585
R500 B.n206 B.n205 585
R501 B.n204 B.n193 585
R502 B.n203 B.n202 585
R503 B.n201 B.n194 585
R504 B.n200 B.n199 585
R505 B.n198 B.n195 585
R506 B.n197 B.n196 585
R507 B.n2 B.n0 585
R508 B.n761 B.n1 585
R509 B.n760 B.n759 585
R510 B.n758 B.n3 585
R511 B.n757 B.n756 585
R512 B.n755 B.n4 585
R513 B.n754 B.n753 585
R514 B.n752 B.n5 585
R515 B.n751 B.n750 585
R516 B.n749 B.n6 585
R517 B.n748 B.n747 585
R518 B.n746 B.n7 585
R519 B.n745 B.n744 585
R520 B.n743 B.n8 585
R521 B.n742 B.n741 585
R522 B.n740 B.n9 585
R523 B.n739 B.n738 585
R524 B.n737 B.n10 585
R525 B.n736 B.n735 585
R526 B.n734 B.n11 585
R527 B.n733 B.n732 585
R528 B.n731 B.n12 585
R529 B.n730 B.n729 585
R530 B.n728 B.n13 585
R531 B.n727 B.n726 585
R532 B.n725 B.n14 585
R533 B.n724 B.n723 585
R534 B.n722 B.n15 585
R535 B.n721 B.n720 585
R536 B.n719 B.n16 585
R537 B.n718 B.n717 585
R538 B.n716 B.n17 585
R539 B.n715 B.n714 585
R540 B.n713 B.n18 585
R541 B.n712 B.n711 585
R542 B.n710 B.n19 585
R543 B.n709 B.n708 585
R544 B.n707 B.n20 585
R545 B.n706 B.n705 585
R546 B.n704 B.n21 585
R547 B.n703 B.n702 585
R548 B.n701 B.n22 585
R549 B.n700 B.n699 585
R550 B.n698 B.n23 585
R551 B.n697 B.n696 585
R552 B.n695 B.n24 585
R553 B.n694 B.n693 585
R554 B.n692 B.n25 585
R555 B.n691 B.n690 585
R556 B.n689 B.n26 585
R557 B.n688 B.n687 585
R558 B.n763 B.n762 585
R559 B.n270 B.n269 473.281
R560 B.n688 B.n27 473.281
R561 B.n405 B.n126 473.281
R562 B.n556 B.n555 473.281
R563 B.n341 B.t6 291.152
R564 B.n151 B.t0 291.152
R565 B.n48 B.t3 291.152
R566 B.n55 B.t9 291.152
R567 B.n341 B.t8 178.535
R568 B.n55 B.t10 178.535
R569 B.n151 B.t2 178.522
R570 B.n48 B.t4 178.522
R571 B.n269 B.n172 163.367
R572 B.n265 B.n172 163.367
R573 B.n265 B.n264 163.367
R574 B.n264 B.n263 163.367
R575 B.n263 B.n174 163.367
R576 B.n259 B.n174 163.367
R577 B.n259 B.n258 163.367
R578 B.n258 B.n257 163.367
R579 B.n257 B.n176 163.367
R580 B.n253 B.n176 163.367
R581 B.n253 B.n252 163.367
R582 B.n252 B.n251 163.367
R583 B.n251 B.n178 163.367
R584 B.n247 B.n178 163.367
R585 B.n247 B.n246 163.367
R586 B.n246 B.n245 163.367
R587 B.n245 B.n180 163.367
R588 B.n241 B.n180 163.367
R589 B.n241 B.n240 163.367
R590 B.n240 B.n239 163.367
R591 B.n239 B.n182 163.367
R592 B.n235 B.n182 163.367
R593 B.n235 B.n234 163.367
R594 B.n234 B.n233 163.367
R595 B.n233 B.n184 163.367
R596 B.n229 B.n184 163.367
R597 B.n229 B.n228 163.367
R598 B.n228 B.n227 163.367
R599 B.n227 B.n186 163.367
R600 B.n223 B.n186 163.367
R601 B.n223 B.n222 163.367
R602 B.n222 B.n221 163.367
R603 B.n221 B.n188 163.367
R604 B.n217 B.n188 163.367
R605 B.n217 B.n216 163.367
R606 B.n216 B.n215 163.367
R607 B.n215 B.n190 163.367
R608 B.n211 B.n190 163.367
R609 B.n211 B.n210 163.367
R610 B.n210 B.n209 163.367
R611 B.n209 B.n192 163.367
R612 B.n205 B.n192 163.367
R613 B.n205 B.n204 163.367
R614 B.n204 B.n203 163.367
R615 B.n203 B.n194 163.367
R616 B.n199 B.n194 163.367
R617 B.n199 B.n198 163.367
R618 B.n198 B.n197 163.367
R619 B.n197 B.n2 163.367
R620 B.n762 B.n2 163.367
R621 B.n762 B.n761 163.367
R622 B.n761 B.n760 163.367
R623 B.n760 B.n3 163.367
R624 B.n756 B.n3 163.367
R625 B.n756 B.n755 163.367
R626 B.n755 B.n754 163.367
R627 B.n754 B.n5 163.367
R628 B.n750 B.n5 163.367
R629 B.n750 B.n749 163.367
R630 B.n749 B.n748 163.367
R631 B.n748 B.n7 163.367
R632 B.n744 B.n7 163.367
R633 B.n744 B.n743 163.367
R634 B.n743 B.n742 163.367
R635 B.n742 B.n9 163.367
R636 B.n738 B.n9 163.367
R637 B.n738 B.n737 163.367
R638 B.n737 B.n736 163.367
R639 B.n736 B.n11 163.367
R640 B.n732 B.n11 163.367
R641 B.n732 B.n731 163.367
R642 B.n731 B.n730 163.367
R643 B.n730 B.n13 163.367
R644 B.n726 B.n13 163.367
R645 B.n726 B.n725 163.367
R646 B.n725 B.n724 163.367
R647 B.n724 B.n15 163.367
R648 B.n720 B.n15 163.367
R649 B.n720 B.n719 163.367
R650 B.n719 B.n718 163.367
R651 B.n718 B.n17 163.367
R652 B.n714 B.n17 163.367
R653 B.n714 B.n713 163.367
R654 B.n713 B.n712 163.367
R655 B.n712 B.n19 163.367
R656 B.n708 B.n19 163.367
R657 B.n708 B.n707 163.367
R658 B.n707 B.n706 163.367
R659 B.n706 B.n21 163.367
R660 B.n702 B.n21 163.367
R661 B.n702 B.n701 163.367
R662 B.n701 B.n700 163.367
R663 B.n700 B.n23 163.367
R664 B.n696 B.n23 163.367
R665 B.n696 B.n695 163.367
R666 B.n695 B.n694 163.367
R667 B.n694 B.n25 163.367
R668 B.n690 B.n25 163.367
R669 B.n690 B.n689 163.367
R670 B.n689 B.n688 163.367
R671 B.n271 B.n270 163.367
R672 B.n271 B.n170 163.367
R673 B.n275 B.n170 163.367
R674 B.n276 B.n275 163.367
R675 B.n277 B.n276 163.367
R676 B.n277 B.n168 163.367
R677 B.n281 B.n168 163.367
R678 B.n282 B.n281 163.367
R679 B.n283 B.n282 163.367
R680 B.n283 B.n166 163.367
R681 B.n287 B.n166 163.367
R682 B.n288 B.n287 163.367
R683 B.n289 B.n288 163.367
R684 B.n289 B.n164 163.367
R685 B.n293 B.n164 163.367
R686 B.n294 B.n293 163.367
R687 B.n295 B.n294 163.367
R688 B.n295 B.n162 163.367
R689 B.n299 B.n162 163.367
R690 B.n300 B.n299 163.367
R691 B.n301 B.n300 163.367
R692 B.n301 B.n160 163.367
R693 B.n305 B.n160 163.367
R694 B.n306 B.n305 163.367
R695 B.n307 B.n306 163.367
R696 B.n307 B.n158 163.367
R697 B.n311 B.n158 163.367
R698 B.n312 B.n311 163.367
R699 B.n313 B.n312 163.367
R700 B.n313 B.n156 163.367
R701 B.n317 B.n156 163.367
R702 B.n318 B.n317 163.367
R703 B.n319 B.n318 163.367
R704 B.n319 B.n154 163.367
R705 B.n323 B.n154 163.367
R706 B.n324 B.n323 163.367
R707 B.n325 B.n324 163.367
R708 B.n325 B.n150 163.367
R709 B.n330 B.n150 163.367
R710 B.n331 B.n330 163.367
R711 B.n332 B.n331 163.367
R712 B.n332 B.n148 163.367
R713 B.n336 B.n148 163.367
R714 B.n337 B.n336 163.367
R715 B.n338 B.n337 163.367
R716 B.n338 B.n146 163.367
R717 B.n345 B.n146 163.367
R718 B.n346 B.n345 163.367
R719 B.n347 B.n346 163.367
R720 B.n347 B.n144 163.367
R721 B.n351 B.n144 163.367
R722 B.n352 B.n351 163.367
R723 B.n353 B.n352 163.367
R724 B.n353 B.n142 163.367
R725 B.n357 B.n142 163.367
R726 B.n358 B.n357 163.367
R727 B.n359 B.n358 163.367
R728 B.n359 B.n140 163.367
R729 B.n363 B.n140 163.367
R730 B.n364 B.n363 163.367
R731 B.n365 B.n364 163.367
R732 B.n365 B.n138 163.367
R733 B.n369 B.n138 163.367
R734 B.n370 B.n369 163.367
R735 B.n371 B.n370 163.367
R736 B.n371 B.n136 163.367
R737 B.n375 B.n136 163.367
R738 B.n376 B.n375 163.367
R739 B.n377 B.n376 163.367
R740 B.n377 B.n134 163.367
R741 B.n381 B.n134 163.367
R742 B.n382 B.n381 163.367
R743 B.n383 B.n382 163.367
R744 B.n383 B.n132 163.367
R745 B.n387 B.n132 163.367
R746 B.n388 B.n387 163.367
R747 B.n389 B.n388 163.367
R748 B.n389 B.n130 163.367
R749 B.n393 B.n130 163.367
R750 B.n394 B.n393 163.367
R751 B.n395 B.n394 163.367
R752 B.n395 B.n128 163.367
R753 B.n399 B.n128 163.367
R754 B.n400 B.n399 163.367
R755 B.n401 B.n400 163.367
R756 B.n401 B.n126 163.367
R757 B.n406 B.n405 163.367
R758 B.n407 B.n406 163.367
R759 B.n407 B.n124 163.367
R760 B.n411 B.n124 163.367
R761 B.n412 B.n411 163.367
R762 B.n413 B.n412 163.367
R763 B.n413 B.n122 163.367
R764 B.n417 B.n122 163.367
R765 B.n418 B.n417 163.367
R766 B.n419 B.n418 163.367
R767 B.n419 B.n120 163.367
R768 B.n423 B.n120 163.367
R769 B.n424 B.n423 163.367
R770 B.n425 B.n424 163.367
R771 B.n425 B.n118 163.367
R772 B.n429 B.n118 163.367
R773 B.n430 B.n429 163.367
R774 B.n431 B.n430 163.367
R775 B.n431 B.n116 163.367
R776 B.n435 B.n116 163.367
R777 B.n436 B.n435 163.367
R778 B.n437 B.n436 163.367
R779 B.n437 B.n114 163.367
R780 B.n441 B.n114 163.367
R781 B.n442 B.n441 163.367
R782 B.n443 B.n442 163.367
R783 B.n443 B.n112 163.367
R784 B.n447 B.n112 163.367
R785 B.n448 B.n447 163.367
R786 B.n449 B.n448 163.367
R787 B.n449 B.n110 163.367
R788 B.n453 B.n110 163.367
R789 B.n454 B.n453 163.367
R790 B.n455 B.n454 163.367
R791 B.n455 B.n108 163.367
R792 B.n459 B.n108 163.367
R793 B.n460 B.n459 163.367
R794 B.n461 B.n460 163.367
R795 B.n461 B.n106 163.367
R796 B.n465 B.n106 163.367
R797 B.n466 B.n465 163.367
R798 B.n467 B.n466 163.367
R799 B.n467 B.n104 163.367
R800 B.n471 B.n104 163.367
R801 B.n472 B.n471 163.367
R802 B.n473 B.n472 163.367
R803 B.n473 B.n102 163.367
R804 B.n477 B.n102 163.367
R805 B.n478 B.n477 163.367
R806 B.n479 B.n478 163.367
R807 B.n479 B.n100 163.367
R808 B.n483 B.n100 163.367
R809 B.n484 B.n483 163.367
R810 B.n485 B.n484 163.367
R811 B.n485 B.n98 163.367
R812 B.n489 B.n98 163.367
R813 B.n490 B.n489 163.367
R814 B.n491 B.n490 163.367
R815 B.n491 B.n96 163.367
R816 B.n495 B.n96 163.367
R817 B.n496 B.n495 163.367
R818 B.n497 B.n496 163.367
R819 B.n497 B.n94 163.367
R820 B.n501 B.n94 163.367
R821 B.n502 B.n501 163.367
R822 B.n503 B.n502 163.367
R823 B.n503 B.n92 163.367
R824 B.n507 B.n92 163.367
R825 B.n508 B.n507 163.367
R826 B.n509 B.n508 163.367
R827 B.n509 B.n90 163.367
R828 B.n513 B.n90 163.367
R829 B.n514 B.n513 163.367
R830 B.n515 B.n514 163.367
R831 B.n515 B.n88 163.367
R832 B.n519 B.n88 163.367
R833 B.n520 B.n519 163.367
R834 B.n521 B.n520 163.367
R835 B.n521 B.n86 163.367
R836 B.n525 B.n86 163.367
R837 B.n526 B.n525 163.367
R838 B.n527 B.n526 163.367
R839 B.n527 B.n84 163.367
R840 B.n531 B.n84 163.367
R841 B.n532 B.n531 163.367
R842 B.n533 B.n532 163.367
R843 B.n533 B.n82 163.367
R844 B.n537 B.n82 163.367
R845 B.n538 B.n537 163.367
R846 B.n539 B.n538 163.367
R847 B.n539 B.n80 163.367
R848 B.n543 B.n80 163.367
R849 B.n544 B.n543 163.367
R850 B.n545 B.n544 163.367
R851 B.n545 B.n78 163.367
R852 B.n549 B.n78 163.367
R853 B.n550 B.n549 163.367
R854 B.n551 B.n550 163.367
R855 B.n551 B.n76 163.367
R856 B.n555 B.n76 163.367
R857 B.n684 B.n27 163.367
R858 B.n684 B.n683 163.367
R859 B.n683 B.n682 163.367
R860 B.n682 B.n29 163.367
R861 B.n678 B.n29 163.367
R862 B.n678 B.n677 163.367
R863 B.n677 B.n676 163.367
R864 B.n676 B.n31 163.367
R865 B.n672 B.n31 163.367
R866 B.n672 B.n671 163.367
R867 B.n671 B.n670 163.367
R868 B.n670 B.n33 163.367
R869 B.n666 B.n33 163.367
R870 B.n666 B.n665 163.367
R871 B.n665 B.n664 163.367
R872 B.n664 B.n35 163.367
R873 B.n660 B.n35 163.367
R874 B.n660 B.n659 163.367
R875 B.n659 B.n658 163.367
R876 B.n658 B.n37 163.367
R877 B.n654 B.n37 163.367
R878 B.n654 B.n653 163.367
R879 B.n653 B.n652 163.367
R880 B.n652 B.n39 163.367
R881 B.n648 B.n39 163.367
R882 B.n648 B.n647 163.367
R883 B.n647 B.n646 163.367
R884 B.n646 B.n41 163.367
R885 B.n642 B.n41 163.367
R886 B.n642 B.n641 163.367
R887 B.n641 B.n640 163.367
R888 B.n640 B.n43 163.367
R889 B.n636 B.n43 163.367
R890 B.n636 B.n635 163.367
R891 B.n635 B.n634 163.367
R892 B.n634 B.n45 163.367
R893 B.n630 B.n45 163.367
R894 B.n630 B.n629 163.367
R895 B.n629 B.n628 163.367
R896 B.n628 B.n47 163.367
R897 B.n624 B.n47 163.367
R898 B.n624 B.n623 163.367
R899 B.n623 B.n622 163.367
R900 B.n622 B.n52 163.367
R901 B.n618 B.n52 163.367
R902 B.n618 B.n617 163.367
R903 B.n617 B.n616 163.367
R904 B.n616 B.n54 163.367
R905 B.n611 B.n54 163.367
R906 B.n611 B.n610 163.367
R907 B.n610 B.n609 163.367
R908 B.n609 B.n58 163.367
R909 B.n605 B.n58 163.367
R910 B.n605 B.n604 163.367
R911 B.n604 B.n603 163.367
R912 B.n603 B.n60 163.367
R913 B.n599 B.n60 163.367
R914 B.n599 B.n598 163.367
R915 B.n598 B.n597 163.367
R916 B.n597 B.n62 163.367
R917 B.n593 B.n62 163.367
R918 B.n593 B.n592 163.367
R919 B.n592 B.n591 163.367
R920 B.n591 B.n64 163.367
R921 B.n587 B.n64 163.367
R922 B.n587 B.n586 163.367
R923 B.n586 B.n585 163.367
R924 B.n585 B.n66 163.367
R925 B.n581 B.n66 163.367
R926 B.n581 B.n580 163.367
R927 B.n580 B.n579 163.367
R928 B.n579 B.n68 163.367
R929 B.n575 B.n68 163.367
R930 B.n575 B.n574 163.367
R931 B.n574 B.n573 163.367
R932 B.n573 B.n70 163.367
R933 B.n569 B.n70 163.367
R934 B.n569 B.n568 163.367
R935 B.n568 B.n567 163.367
R936 B.n567 B.n72 163.367
R937 B.n563 B.n72 163.367
R938 B.n563 B.n562 163.367
R939 B.n562 B.n561 163.367
R940 B.n561 B.n74 163.367
R941 B.n557 B.n74 163.367
R942 B.n557 B.n556 163.367
R943 B.n342 B.t7 109.686
R944 B.n56 B.t11 109.686
R945 B.n152 B.t1 109.674
R946 B.n49 B.t5 109.674
R947 B.n342 B.n341 68.849
R948 B.n152 B.n151 68.849
R949 B.n49 B.n48 68.849
R950 B.n56 B.n55 68.849
R951 B.n343 B.n342 59.5399
R952 B.n328 B.n152 59.5399
R953 B.n50 B.n49 59.5399
R954 B.n614 B.n56 59.5399
R955 B.n687 B.n686 30.7517
R956 B.n554 B.n75 30.7517
R957 B.n404 B.n403 30.7517
R958 B.n268 B.n171 30.7517
R959 B B.n763 18.0485
R960 B.n686 B.n685 10.6151
R961 B.n685 B.n28 10.6151
R962 B.n681 B.n28 10.6151
R963 B.n681 B.n680 10.6151
R964 B.n680 B.n679 10.6151
R965 B.n679 B.n30 10.6151
R966 B.n675 B.n30 10.6151
R967 B.n675 B.n674 10.6151
R968 B.n674 B.n673 10.6151
R969 B.n673 B.n32 10.6151
R970 B.n669 B.n32 10.6151
R971 B.n669 B.n668 10.6151
R972 B.n668 B.n667 10.6151
R973 B.n667 B.n34 10.6151
R974 B.n663 B.n34 10.6151
R975 B.n663 B.n662 10.6151
R976 B.n662 B.n661 10.6151
R977 B.n661 B.n36 10.6151
R978 B.n657 B.n36 10.6151
R979 B.n657 B.n656 10.6151
R980 B.n656 B.n655 10.6151
R981 B.n655 B.n38 10.6151
R982 B.n651 B.n38 10.6151
R983 B.n651 B.n650 10.6151
R984 B.n650 B.n649 10.6151
R985 B.n649 B.n40 10.6151
R986 B.n645 B.n40 10.6151
R987 B.n645 B.n644 10.6151
R988 B.n644 B.n643 10.6151
R989 B.n643 B.n42 10.6151
R990 B.n639 B.n42 10.6151
R991 B.n639 B.n638 10.6151
R992 B.n638 B.n637 10.6151
R993 B.n637 B.n44 10.6151
R994 B.n633 B.n44 10.6151
R995 B.n633 B.n632 10.6151
R996 B.n632 B.n631 10.6151
R997 B.n631 B.n46 10.6151
R998 B.n627 B.n626 10.6151
R999 B.n626 B.n625 10.6151
R1000 B.n625 B.n51 10.6151
R1001 B.n621 B.n51 10.6151
R1002 B.n621 B.n620 10.6151
R1003 B.n620 B.n619 10.6151
R1004 B.n619 B.n53 10.6151
R1005 B.n615 B.n53 10.6151
R1006 B.n613 B.n612 10.6151
R1007 B.n612 B.n57 10.6151
R1008 B.n608 B.n57 10.6151
R1009 B.n608 B.n607 10.6151
R1010 B.n607 B.n606 10.6151
R1011 B.n606 B.n59 10.6151
R1012 B.n602 B.n59 10.6151
R1013 B.n602 B.n601 10.6151
R1014 B.n601 B.n600 10.6151
R1015 B.n600 B.n61 10.6151
R1016 B.n596 B.n61 10.6151
R1017 B.n596 B.n595 10.6151
R1018 B.n595 B.n594 10.6151
R1019 B.n594 B.n63 10.6151
R1020 B.n590 B.n63 10.6151
R1021 B.n590 B.n589 10.6151
R1022 B.n589 B.n588 10.6151
R1023 B.n588 B.n65 10.6151
R1024 B.n584 B.n65 10.6151
R1025 B.n584 B.n583 10.6151
R1026 B.n583 B.n582 10.6151
R1027 B.n582 B.n67 10.6151
R1028 B.n578 B.n67 10.6151
R1029 B.n578 B.n577 10.6151
R1030 B.n577 B.n576 10.6151
R1031 B.n576 B.n69 10.6151
R1032 B.n572 B.n69 10.6151
R1033 B.n572 B.n571 10.6151
R1034 B.n571 B.n570 10.6151
R1035 B.n570 B.n71 10.6151
R1036 B.n566 B.n71 10.6151
R1037 B.n566 B.n565 10.6151
R1038 B.n565 B.n564 10.6151
R1039 B.n564 B.n73 10.6151
R1040 B.n560 B.n73 10.6151
R1041 B.n560 B.n559 10.6151
R1042 B.n559 B.n558 10.6151
R1043 B.n558 B.n75 10.6151
R1044 B.n404 B.n125 10.6151
R1045 B.n408 B.n125 10.6151
R1046 B.n409 B.n408 10.6151
R1047 B.n410 B.n409 10.6151
R1048 B.n410 B.n123 10.6151
R1049 B.n414 B.n123 10.6151
R1050 B.n415 B.n414 10.6151
R1051 B.n416 B.n415 10.6151
R1052 B.n416 B.n121 10.6151
R1053 B.n420 B.n121 10.6151
R1054 B.n421 B.n420 10.6151
R1055 B.n422 B.n421 10.6151
R1056 B.n422 B.n119 10.6151
R1057 B.n426 B.n119 10.6151
R1058 B.n427 B.n426 10.6151
R1059 B.n428 B.n427 10.6151
R1060 B.n428 B.n117 10.6151
R1061 B.n432 B.n117 10.6151
R1062 B.n433 B.n432 10.6151
R1063 B.n434 B.n433 10.6151
R1064 B.n434 B.n115 10.6151
R1065 B.n438 B.n115 10.6151
R1066 B.n439 B.n438 10.6151
R1067 B.n440 B.n439 10.6151
R1068 B.n440 B.n113 10.6151
R1069 B.n444 B.n113 10.6151
R1070 B.n445 B.n444 10.6151
R1071 B.n446 B.n445 10.6151
R1072 B.n446 B.n111 10.6151
R1073 B.n450 B.n111 10.6151
R1074 B.n451 B.n450 10.6151
R1075 B.n452 B.n451 10.6151
R1076 B.n452 B.n109 10.6151
R1077 B.n456 B.n109 10.6151
R1078 B.n457 B.n456 10.6151
R1079 B.n458 B.n457 10.6151
R1080 B.n458 B.n107 10.6151
R1081 B.n462 B.n107 10.6151
R1082 B.n463 B.n462 10.6151
R1083 B.n464 B.n463 10.6151
R1084 B.n464 B.n105 10.6151
R1085 B.n468 B.n105 10.6151
R1086 B.n469 B.n468 10.6151
R1087 B.n470 B.n469 10.6151
R1088 B.n470 B.n103 10.6151
R1089 B.n474 B.n103 10.6151
R1090 B.n475 B.n474 10.6151
R1091 B.n476 B.n475 10.6151
R1092 B.n476 B.n101 10.6151
R1093 B.n480 B.n101 10.6151
R1094 B.n481 B.n480 10.6151
R1095 B.n482 B.n481 10.6151
R1096 B.n482 B.n99 10.6151
R1097 B.n486 B.n99 10.6151
R1098 B.n487 B.n486 10.6151
R1099 B.n488 B.n487 10.6151
R1100 B.n488 B.n97 10.6151
R1101 B.n492 B.n97 10.6151
R1102 B.n493 B.n492 10.6151
R1103 B.n494 B.n493 10.6151
R1104 B.n494 B.n95 10.6151
R1105 B.n498 B.n95 10.6151
R1106 B.n499 B.n498 10.6151
R1107 B.n500 B.n499 10.6151
R1108 B.n500 B.n93 10.6151
R1109 B.n504 B.n93 10.6151
R1110 B.n505 B.n504 10.6151
R1111 B.n506 B.n505 10.6151
R1112 B.n506 B.n91 10.6151
R1113 B.n510 B.n91 10.6151
R1114 B.n511 B.n510 10.6151
R1115 B.n512 B.n511 10.6151
R1116 B.n512 B.n89 10.6151
R1117 B.n516 B.n89 10.6151
R1118 B.n517 B.n516 10.6151
R1119 B.n518 B.n517 10.6151
R1120 B.n518 B.n87 10.6151
R1121 B.n522 B.n87 10.6151
R1122 B.n523 B.n522 10.6151
R1123 B.n524 B.n523 10.6151
R1124 B.n524 B.n85 10.6151
R1125 B.n528 B.n85 10.6151
R1126 B.n529 B.n528 10.6151
R1127 B.n530 B.n529 10.6151
R1128 B.n530 B.n83 10.6151
R1129 B.n534 B.n83 10.6151
R1130 B.n535 B.n534 10.6151
R1131 B.n536 B.n535 10.6151
R1132 B.n536 B.n81 10.6151
R1133 B.n540 B.n81 10.6151
R1134 B.n541 B.n540 10.6151
R1135 B.n542 B.n541 10.6151
R1136 B.n542 B.n79 10.6151
R1137 B.n546 B.n79 10.6151
R1138 B.n547 B.n546 10.6151
R1139 B.n548 B.n547 10.6151
R1140 B.n548 B.n77 10.6151
R1141 B.n552 B.n77 10.6151
R1142 B.n553 B.n552 10.6151
R1143 B.n554 B.n553 10.6151
R1144 B.n272 B.n171 10.6151
R1145 B.n273 B.n272 10.6151
R1146 B.n274 B.n273 10.6151
R1147 B.n274 B.n169 10.6151
R1148 B.n278 B.n169 10.6151
R1149 B.n279 B.n278 10.6151
R1150 B.n280 B.n279 10.6151
R1151 B.n280 B.n167 10.6151
R1152 B.n284 B.n167 10.6151
R1153 B.n285 B.n284 10.6151
R1154 B.n286 B.n285 10.6151
R1155 B.n286 B.n165 10.6151
R1156 B.n290 B.n165 10.6151
R1157 B.n291 B.n290 10.6151
R1158 B.n292 B.n291 10.6151
R1159 B.n292 B.n163 10.6151
R1160 B.n296 B.n163 10.6151
R1161 B.n297 B.n296 10.6151
R1162 B.n298 B.n297 10.6151
R1163 B.n298 B.n161 10.6151
R1164 B.n302 B.n161 10.6151
R1165 B.n303 B.n302 10.6151
R1166 B.n304 B.n303 10.6151
R1167 B.n304 B.n159 10.6151
R1168 B.n308 B.n159 10.6151
R1169 B.n309 B.n308 10.6151
R1170 B.n310 B.n309 10.6151
R1171 B.n310 B.n157 10.6151
R1172 B.n314 B.n157 10.6151
R1173 B.n315 B.n314 10.6151
R1174 B.n316 B.n315 10.6151
R1175 B.n316 B.n155 10.6151
R1176 B.n320 B.n155 10.6151
R1177 B.n321 B.n320 10.6151
R1178 B.n322 B.n321 10.6151
R1179 B.n322 B.n153 10.6151
R1180 B.n326 B.n153 10.6151
R1181 B.n327 B.n326 10.6151
R1182 B.n329 B.n149 10.6151
R1183 B.n333 B.n149 10.6151
R1184 B.n334 B.n333 10.6151
R1185 B.n335 B.n334 10.6151
R1186 B.n335 B.n147 10.6151
R1187 B.n339 B.n147 10.6151
R1188 B.n340 B.n339 10.6151
R1189 B.n344 B.n340 10.6151
R1190 B.n348 B.n145 10.6151
R1191 B.n349 B.n348 10.6151
R1192 B.n350 B.n349 10.6151
R1193 B.n350 B.n143 10.6151
R1194 B.n354 B.n143 10.6151
R1195 B.n355 B.n354 10.6151
R1196 B.n356 B.n355 10.6151
R1197 B.n356 B.n141 10.6151
R1198 B.n360 B.n141 10.6151
R1199 B.n361 B.n360 10.6151
R1200 B.n362 B.n361 10.6151
R1201 B.n362 B.n139 10.6151
R1202 B.n366 B.n139 10.6151
R1203 B.n367 B.n366 10.6151
R1204 B.n368 B.n367 10.6151
R1205 B.n368 B.n137 10.6151
R1206 B.n372 B.n137 10.6151
R1207 B.n373 B.n372 10.6151
R1208 B.n374 B.n373 10.6151
R1209 B.n374 B.n135 10.6151
R1210 B.n378 B.n135 10.6151
R1211 B.n379 B.n378 10.6151
R1212 B.n380 B.n379 10.6151
R1213 B.n380 B.n133 10.6151
R1214 B.n384 B.n133 10.6151
R1215 B.n385 B.n384 10.6151
R1216 B.n386 B.n385 10.6151
R1217 B.n386 B.n131 10.6151
R1218 B.n390 B.n131 10.6151
R1219 B.n391 B.n390 10.6151
R1220 B.n392 B.n391 10.6151
R1221 B.n392 B.n129 10.6151
R1222 B.n396 B.n129 10.6151
R1223 B.n397 B.n396 10.6151
R1224 B.n398 B.n397 10.6151
R1225 B.n398 B.n127 10.6151
R1226 B.n402 B.n127 10.6151
R1227 B.n403 B.n402 10.6151
R1228 B.n268 B.n267 10.6151
R1229 B.n267 B.n266 10.6151
R1230 B.n266 B.n173 10.6151
R1231 B.n262 B.n173 10.6151
R1232 B.n262 B.n261 10.6151
R1233 B.n261 B.n260 10.6151
R1234 B.n260 B.n175 10.6151
R1235 B.n256 B.n175 10.6151
R1236 B.n256 B.n255 10.6151
R1237 B.n255 B.n254 10.6151
R1238 B.n254 B.n177 10.6151
R1239 B.n250 B.n177 10.6151
R1240 B.n250 B.n249 10.6151
R1241 B.n249 B.n248 10.6151
R1242 B.n248 B.n179 10.6151
R1243 B.n244 B.n179 10.6151
R1244 B.n244 B.n243 10.6151
R1245 B.n243 B.n242 10.6151
R1246 B.n242 B.n181 10.6151
R1247 B.n238 B.n181 10.6151
R1248 B.n238 B.n237 10.6151
R1249 B.n237 B.n236 10.6151
R1250 B.n236 B.n183 10.6151
R1251 B.n232 B.n183 10.6151
R1252 B.n232 B.n231 10.6151
R1253 B.n231 B.n230 10.6151
R1254 B.n230 B.n185 10.6151
R1255 B.n226 B.n185 10.6151
R1256 B.n226 B.n225 10.6151
R1257 B.n225 B.n224 10.6151
R1258 B.n224 B.n187 10.6151
R1259 B.n220 B.n187 10.6151
R1260 B.n220 B.n219 10.6151
R1261 B.n219 B.n218 10.6151
R1262 B.n218 B.n189 10.6151
R1263 B.n214 B.n189 10.6151
R1264 B.n214 B.n213 10.6151
R1265 B.n213 B.n212 10.6151
R1266 B.n212 B.n191 10.6151
R1267 B.n208 B.n191 10.6151
R1268 B.n208 B.n207 10.6151
R1269 B.n207 B.n206 10.6151
R1270 B.n206 B.n193 10.6151
R1271 B.n202 B.n193 10.6151
R1272 B.n202 B.n201 10.6151
R1273 B.n201 B.n200 10.6151
R1274 B.n200 B.n195 10.6151
R1275 B.n196 B.n195 10.6151
R1276 B.n196 B.n0 10.6151
R1277 B.n759 B.n1 10.6151
R1278 B.n759 B.n758 10.6151
R1279 B.n758 B.n757 10.6151
R1280 B.n757 B.n4 10.6151
R1281 B.n753 B.n4 10.6151
R1282 B.n753 B.n752 10.6151
R1283 B.n752 B.n751 10.6151
R1284 B.n751 B.n6 10.6151
R1285 B.n747 B.n6 10.6151
R1286 B.n747 B.n746 10.6151
R1287 B.n746 B.n745 10.6151
R1288 B.n745 B.n8 10.6151
R1289 B.n741 B.n8 10.6151
R1290 B.n741 B.n740 10.6151
R1291 B.n740 B.n739 10.6151
R1292 B.n739 B.n10 10.6151
R1293 B.n735 B.n10 10.6151
R1294 B.n735 B.n734 10.6151
R1295 B.n734 B.n733 10.6151
R1296 B.n733 B.n12 10.6151
R1297 B.n729 B.n12 10.6151
R1298 B.n729 B.n728 10.6151
R1299 B.n728 B.n727 10.6151
R1300 B.n727 B.n14 10.6151
R1301 B.n723 B.n14 10.6151
R1302 B.n723 B.n722 10.6151
R1303 B.n722 B.n721 10.6151
R1304 B.n721 B.n16 10.6151
R1305 B.n717 B.n16 10.6151
R1306 B.n717 B.n716 10.6151
R1307 B.n716 B.n715 10.6151
R1308 B.n715 B.n18 10.6151
R1309 B.n711 B.n18 10.6151
R1310 B.n711 B.n710 10.6151
R1311 B.n710 B.n709 10.6151
R1312 B.n709 B.n20 10.6151
R1313 B.n705 B.n20 10.6151
R1314 B.n705 B.n704 10.6151
R1315 B.n704 B.n703 10.6151
R1316 B.n703 B.n22 10.6151
R1317 B.n699 B.n22 10.6151
R1318 B.n699 B.n698 10.6151
R1319 B.n698 B.n697 10.6151
R1320 B.n697 B.n24 10.6151
R1321 B.n693 B.n24 10.6151
R1322 B.n693 B.n692 10.6151
R1323 B.n692 B.n691 10.6151
R1324 B.n691 B.n26 10.6151
R1325 B.n687 B.n26 10.6151
R1326 B.n627 B.n50 6.5566
R1327 B.n615 B.n614 6.5566
R1328 B.n329 B.n328 6.5566
R1329 B.n344 B.n343 6.5566
R1330 B.n50 B.n46 4.05904
R1331 B.n614 B.n613 4.05904
R1332 B.n328 B.n327 4.05904
R1333 B.n343 B.n145 4.05904
R1334 B.n763 B.n0 2.81026
R1335 B.n763 B.n1 2.81026
C0 B w_n3810_n3168# 10.2521f
C1 VN VTAIL 6.78729f
C2 VTAIL VDD1 7.57008f
C3 VTAIL VDD2 7.62583f
C4 VN w_n3810_n3168# 7.34893f
C5 w_n3810_n3168# VDD1 2.3702f
C6 VDD2 w_n3810_n3168# 2.47508f
C7 B VN 1.29056f
C8 VTAIL VP 6.80153f
C9 B VDD1 2.17506f
C10 B VDD2 2.26402f
C11 w_n3810_n3168# VP 7.84323f
C12 VN VDD2 6.43238f
C13 VN VDD1 0.151755f
C14 VDD2 VDD1 1.64755f
C15 B VP 2.11898f
C16 VTAIL w_n3810_n3168# 2.88527f
C17 VN VP 7.340681f
C18 VDD1 VP 6.78868f
C19 VDD2 VP 0.51099f
C20 B VTAIL 3.70091f
C21 VDD2 VSUBS 2.053486f
C22 VDD1 VSUBS 2.59128f
C23 VTAIL VSUBS 1.277671f
C24 VN VSUBS 6.4065f
C25 VP VSUBS 3.387505f
C26 B VSUBS 5.166743f
C27 w_n3810_n3168# VSUBS 0.148819p
C28 B.n0 VSUBS 0.005658f
C29 B.n1 VSUBS 0.005658f
C30 B.n2 VSUBS 0.008948f
C31 B.n3 VSUBS 0.008948f
C32 B.n4 VSUBS 0.008948f
C33 B.n5 VSUBS 0.008948f
C34 B.n6 VSUBS 0.008948f
C35 B.n7 VSUBS 0.008948f
C36 B.n8 VSUBS 0.008948f
C37 B.n9 VSUBS 0.008948f
C38 B.n10 VSUBS 0.008948f
C39 B.n11 VSUBS 0.008948f
C40 B.n12 VSUBS 0.008948f
C41 B.n13 VSUBS 0.008948f
C42 B.n14 VSUBS 0.008948f
C43 B.n15 VSUBS 0.008948f
C44 B.n16 VSUBS 0.008948f
C45 B.n17 VSUBS 0.008948f
C46 B.n18 VSUBS 0.008948f
C47 B.n19 VSUBS 0.008948f
C48 B.n20 VSUBS 0.008948f
C49 B.n21 VSUBS 0.008948f
C50 B.n22 VSUBS 0.008948f
C51 B.n23 VSUBS 0.008948f
C52 B.n24 VSUBS 0.008948f
C53 B.n25 VSUBS 0.008948f
C54 B.n26 VSUBS 0.008948f
C55 B.n27 VSUBS 0.020584f
C56 B.n28 VSUBS 0.008948f
C57 B.n29 VSUBS 0.008948f
C58 B.n30 VSUBS 0.008948f
C59 B.n31 VSUBS 0.008948f
C60 B.n32 VSUBS 0.008948f
C61 B.n33 VSUBS 0.008948f
C62 B.n34 VSUBS 0.008948f
C63 B.n35 VSUBS 0.008948f
C64 B.n36 VSUBS 0.008948f
C65 B.n37 VSUBS 0.008948f
C66 B.n38 VSUBS 0.008948f
C67 B.n39 VSUBS 0.008948f
C68 B.n40 VSUBS 0.008948f
C69 B.n41 VSUBS 0.008948f
C70 B.n42 VSUBS 0.008948f
C71 B.n43 VSUBS 0.008948f
C72 B.n44 VSUBS 0.008948f
C73 B.n45 VSUBS 0.008948f
C74 B.n46 VSUBS 0.006185f
C75 B.n47 VSUBS 0.008948f
C76 B.t5 VSUBS 0.453765f
C77 B.t4 VSUBS 0.485464f
C78 B.t3 VSUBS 2.10114f
C79 B.n48 VSUBS 0.267479f
C80 B.n49 VSUBS 0.094956f
C81 B.n50 VSUBS 0.020731f
C82 B.n51 VSUBS 0.008948f
C83 B.n52 VSUBS 0.008948f
C84 B.n53 VSUBS 0.008948f
C85 B.n54 VSUBS 0.008948f
C86 B.t11 VSUBS 0.453757f
C87 B.t10 VSUBS 0.485457f
C88 B.t9 VSUBS 2.10114f
C89 B.n55 VSUBS 0.267486f
C90 B.n56 VSUBS 0.094963f
C91 B.n57 VSUBS 0.008948f
C92 B.n58 VSUBS 0.008948f
C93 B.n59 VSUBS 0.008948f
C94 B.n60 VSUBS 0.008948f
C95 B.n61 VSUBS 0.008948f
C96 B.n62 VSUBS 0.008948f
C97 B.n63 VSUBS 0.008948f
C98 B.n64 VSUBS 0.008948f
C99 B.n65 VSUBS 0.008948f
C100 B.n66 VSUBS 0.008948f
C101 B.n67 VSUBS 0.008948f
C102 B.n68 VSUBS 0.008948f
C103 B.n69 VSUBS 0.008948f
C104 B.n70 VSUBS 0.008948f
C105 B.n71 VSUBS 0.008948f
C106 B.n72 VSUBS 0.008948f
C107 B.n73 VSUBS 0.008948f
C108 B.n74 VSUBS 0.008948f
C109 B.n75 VSUBS 0.019462f
C110 B.n76 VSUBS 0.008948f
C111 B.n77 VSUBS 0.008948f
C112 B.n78 VSUBS 0.008948f
C113 B.n79 VSUBS 0.008948f
C114 B.n80 VSUBS 0.008948f
C115 B.n81 VSUBS 0.008948f
C116 B.n82 VSUBS 0.008948f
C117 B.n83 VSUBS 0.008948f
C118 B.n84 VSUBS 0.008948f
C119 B.n85 VSUBS 0.008948f
C120 B.n86 VSUBS 0.008948f
C121 B.n87 VSUBS 0.008948f
C122 B.n88 VSUBS 0.008948f
C123 B.n89 VSUBS 0.008948f
C124 B.n90 VSUBS 0.008948f
C125 B.n91 VSUBS 0.008948f
C126 B.n92 VSUBS 0.008948f
C127 B.n93 VSUBS 0.008948f
C128 B.n94 VSUBS 0.008948f
C129 B.n95 VSUBS 0.008948f
C130 B.n96 VSUBS 0.008948f
C131 B.n97 VSUBS 0.008948f
C132 B.n98 VSUBS 0.008948f
C133 B.n99 VSUBS 0.008948f
C134 B.n100 VSUBS 0.008948f
C135 B.n101 VSUBS 0.008948f
C136 B.n102 VSUBS 0.008948f
C137 B.n103 VSUBS 0.008948f
C138 B.n104 VSUBS 0.008948f
C139 B.n105 VSUBS 0.008948f
C140 B.n106 VSUBS 0.008948f
C141 B.n107 VSUBS 0.008948f
C142 B.n108 VSUBS 0.008948f
C143 B.n109 VSUBS 0.008948f
C144 B.n110 VSUBS 0.008948f
C145 B.n111 VSUBS 0.008948f
C146 B.n112 VSUBS 0.008948f
C147 B.n113 VSUBS 0.008948f
C148 B.n114 VSUBS 0.008948f
C149 B.n115 VSUBS 0.008948f
C150 B.n116 VSUBS 0.008948f
C151 B.n117 VSUBS 0.008948f
C152 B.n118 VSUBS 0.008948f
C153 B.n119 VSUBS 0.008948f
C154 B.n120 VSUBS 0.008948f
C155 B.n121 VSUBS 0.008948f
C156 B.n122 VSUBS 0.008948f
C157 B.n123 VSUBS 0.008948f
C158 B.n124 VSUBS 0.008948f
C159 B.n125 VSUBS 0.008948f
C160 B.n126 VSUBS 0.020584f
C161 B.n127 VSUBS 0.008948f
C162 B.n128 VSUBS 0.008948f
C163 B.n129 VSUBS 0.008948f
C164 B.n130 VSUBS 0.008948f
C165 B.n131 VSUBS 0.008948f
C166 B.n132 VSUBS 0.008948f
C167 B.n133 VSUBS 0.008948f
C168 B.n134 VSUBS 0.008948f
C169 B.n135 VSUBS 0.008948f
C170 B.n136 VSUBS 0.008948f
C171 B.n137 VSUBS 0.008948f
C172 B.n138 VSUBS 0.008948f
C173 B.n139 VSUBS 0.008948f
C174 B.n140 VSUBS 0.008948f
C175 B.n141 VSUBS 0.008948f
C176 B.n142 VSUBS 0.008948f
C177 B.n143 VSUBS 0.008948f
C178 B.n144 VSUBS 0.008948f
C179 B.n145 VSUBS 0.006185f
C180 B.n146 VSUBS 0.008948f
C181 B.n147 VSUBS 0.008948f
C182 B.n148 VSUBS 0.008948f
C183 B.n149 VSUBS 0.008948f
C184 B.n150 VSUBS 0.008948f
C185 B.t1 VSUBS 0.453765f
C186 B.t2 VSUBS 0.485464f
C187 B.t0 VSUBS 2.10114f
C188 B.n151 VSUBS 0.267479f
C189 B.n152 VSUBS 0.094956f
C190 B.n153 VSUBS 0.008948f
C191 B.n154 VSUBS 0.008948f
C192 B.n155 VSUBS 0.008948f
C193 B.n156 VSUBS 0.008948f
C194 B.n157 VSUBS 0.008948f
C195 B.n158 VSUBS 0.008948f
C196 B.n159 VSUBS 0.008948f
C197 B.n160 VSUBS 0.008948f
C198 B.n161 VSUBS 0.008948f
C199 B.n162 VSUBS 0.008948f
C200 B.n163 VSUBS 0.008948f
C201 B.n164 VSUBS 0.008948f
C202 B.n165 VSUBS 0.008948f
C203 B.n166 VSUBS 0.008948f
C204 B.n167 VSUBS 0.008948f
C205 B.n168 VSUBS 0.008948f
C206 B.n169 VSUBS 0.008948f
C207 B.n170 VSUBS 0.008948f
C208 B.n171 VSUBS 0.020584f
C209 B.n172 VSUBS 0.008948f
C210 B.n173 VSUBS 0.008948f
C211 B.n174 VSUBS 0.008948f
C212 B.n175 VSUBS 0.008948f
C213 B.n176 VSUBS 0.008948f
C214 B.n177 VSUBS 0.008948f
C215 B.n178 VSUBS 0.008948f
C216 B.n179 VSUBS 0.008948f
C217 B.n180 VSUBS 0.008948f
C218 B.n181 VSUBS 0.008948f
C219 B.n182 VSUBS 0.008948f
C220 B.n183 VSUBS 0.008948f
C221 B.n184 VSUBS 0.008948f
C222 B.n185 VSUBS 0.008948f
C223 B.n186 VSUBS 0.008948f
C224 B.n187 VSUBS 0.008948f
C225 B.n188 VSUBS 0.008948f
C226 B.n189 VSUBS 0.008948f
C227 B.n190 VSUBS 0.008948f
C228 B.n191 VSUBS 0.008948f
C229 B.n192 VSUBS 0.008948f
C230 B.n193 VSUBS 0.008948f
C231 B.n194 VSUBS 0.008948f
C232 B.n195 VSUBS 0.008948f
C233 B.n196 VSUBS 0.008948f
C234 B.n197 VSUBS 0.008948f
C235 B.n198 VSUBS 0.008948f
C236 B.n199 VSUBS 0.008948f
C237 B.n200 VSUBS 0.008948f
C238 B.n201 VSUBS 0.008948f
C239 B.n202 VSUBS 0.008948f
C240 B.n203 VSUBS 0.008948f
C241 B.n204 VSUBS 0.008948f
C242 B.n205 VSUBS 0.008948f
C243 B.n206 VSUBS 0.008948f
C244 B.n207 VSUBS 0.008948f
C245 B.n208 VSUBS 0.008948f
C246 B.n209 VSUBS 0.008948f
C247 B.n210 VSUBS 0.008948f
C248 B.n211 VSUBS 0.008948f
C249 B.n212 VSUBS 0.008948f
C250 B.n213 VSUBS 0.008948f
C251 B.n214 VSUBS 0.008948f
C252 B.n215 VSUBS 0.008948f
C253 B.n216 VSUBS 0.008948f
C254 B.n217 VSUBS 0.008948f
C255 B.n218 VSUBS 0.008948f
C256 B.n219 VSUBS 0.008948f
C257 B.n220 VSUBS 0.008948f
C258 B.n221 VSUBS 0.008948f
C259 B.n222 VSUBS 0.008948f
C260 B.n223 VSUBS 0.008948f
C261 B.n224 VSUBS 0.008948f
C262 B.n225 VSUBS 0.008948f
C263 B.n226 VSUBS 0.008948f
C264 B.n227 VSUBS 0.008948f
C265 B.n228 VSUBS 0.008948f
C266 B.n229 VSUBS 0.008948f
C267 B.n230 VSUBS 0.008948f
C268 B.n231 VSUBS 0.008948f
C269 B.n232 VSUBS 0.008948f
C270 B.n233 VSUBS 0.008948f
C271 B.n234 VSUBS 0.008948f
C272 B.n235 VSUBS 0.008948f
C273 B.n236 VSUBS 0.008948f
C274 B.n237 VSUBS 0.008948f
C275 B.n238 VSUBS 0.008948f
C276 B.n239 VSUBS 0.008948f
C277 B.n240 VSUBS 0.008948f
C278 B.n241 VSUBS 0.008948f
C279 B.n242 VSUBS 0.008948f
C280 B.n243 VSUBS 0.008948f
C281 B.n244 VSUBS 0.008948f
C282 B.n245 VSUBS 0.008948f
C283 B.n246 VSUBS 0.008948f
C284 B.n247 VSUBS 0.008948f
C285 B.n248 VSUBS 0.008948f
C286 B.n249 VSUBS 0.008948f
C287 B.n250 VSUBS 0.008948f
C288 B.n251 VSUBS 0.008948f
C289 B.n252 VSUBS 0.008948f
C290 B.n253 VSUBS 0.008948f
C291 B.n254 VSUBS 0.008948f
C292 B.n255 VSUBS 0.008948f
C293 B.n256 VSUBS 0.008948f
C294 B.n257 VSUBS 0.008948f
C295 B.n258 VSUBS 0.008948f
C296 B.n259 VSUBS 0.008948f
C297 B.n260 VSUBS 0.008948f
C298 B.n261 VSUBS 0.008948f
C299 B.n262 VSUBS 0.008948f
C300 B.n263 VSUBS 0.008948f
C301 B.n264 VSUBS 0.008948f
C302 B.n265 VSUBS 0.008948f
C303 B.n266 VSUBS 0.008948f
C304 B.n267 VSUBS 0.008948f
C305 B.n268 VSUBS 0.019681f
C306 B.n269 VSUBS 0.019681f
C307 B.n270 VSUBS 0.020584f
C308 B.n271 VSUBS 0.008948f
C309 B.n272 VSUBS 0.008948f
C310 B.n273 VSUBS 0.008948f
C311 B.n274 VSUBS 0.008948f
C312 B.n275 VSUBS 0.008948f
C313 B.n276 VSUBS 0.008948f
C314 B.n277 VSUBS 0.008948f
C315 B.n278 VSUBS 0.008948f
C316 B.n279 VSUBS 0.008948f
C317 B.n280 VSUBS 0.008948f
C318 B.n281 VSUBS 0.008948f
C319 B.n282 VSUBS 0.008948f
C320 B.n283 VSUBS 0.008948f
C321 B.n284 VSUBS 0.008948f
C322 B.n285 VSUBS 0.008948f
C323 B.n286 VSUBS 0.008948f
C324 B.n287 VSUBS 0.008948f
C325 B.n288 VSUBS 0.008948f
C326 B.n289 VSUBS 0.008948f
C327 B.n290 VSUBS 0.008948f
C328 B.n291 VSUBS 0.008948f
C329 B.n292 VSUBS 0.008948f
C330 B.n293 VSUBS 0.008948f
C331 B.n294 VSUBS 0.008948f
C332 B.n295 VSUBS 0.008948f
C333 B.n296 VSUBS 0.008948f
C334 B.n297 VSUBS 0.008948f
C335 B.n298 VSUBS 0.008948f
C336 B.n299 VSUBS 0.008948f
C337 B.n300 VSUBS 0.008948f
C338 B.n301 VSUBS 0.008948f
C339 B.n302 VSUBS 0.008948f
C340 B.n303 VSUBS 0.008948f
C341 B.n304 VSUBS 0.008948f
C342 B.n305 VSUBS 0.008948f
C343 B.n306 VSUBS 0.008948f
C344 B.n307 VSUBS 0.008948f
C345 B.n308 VSUBS 0.008948f
C346 B.n309 VSUBS 0.008948f
C347 B.n310 VSUBS 0.008948f
C348 B.n311 VSUBS 0.008948f
C349 B.n312 VSUBS 0.008948f
C350 B.n313 VSUBS 0.008948f
C351 B.n314 VSUBS 0.008948f
C352 B.n315 VSUBS 0.008948f
C353 B.n316 VSUBS 0.008948f
C354 B.n317 VSUBS 0.008948f
C355 B.n318 VSUBS 0.008948f
C356 B.n319 VSUBS 0.008948f
C357 B.n320 VSUBS 0.008948f
C358 B.n321 VSUBS 0.008948f
C359 B.n322 VSUBS 0.008948f
C360 B.n323 VSUBS 0.008948f
C361 B.n324 VSUBS 0.008948f
C362 B.n325 VSUBS 0.008948f
C363 B.n326 VSUBS 0.008948f
C364 B.n327 VSUBS 0.006185f
C365 B.n328 VSUBS 0.020731f
C366 B.n329 VSUBS 0.007237f
C367 B.n330 VSUBS 0.008948f
C368 B.n331 VSUBS 0.008948f
C369 B.n332 VSUBS 0.008948f
C370 B.n333 VSUBS 0.008948f
C371 B.n334 VSUBS 0.008948f
C372 B.n335 VSUBS 0.008948f
C373 B.n336 VSUBS 0.008948f
C374 B.n337 VSUBS 0.008948f
C375 B.n338 VSUBS 0.008948f
C376 B.n339 VSUBS 0.008948f
C377 B.n340 VSUBS 0.008948f
C378 B.t7 VSUBS 0.453757f
C379 B.t8 VSUBS 0.485457f
C380 B.t6 VSUBS 2.10114f
C381 B.n341 VSUBS 0.267486f
C382 B.n342 VSUBS 0.094963f
C383 B.n343 VSUBS 0.020731f
C384 B.n344 VSUBS 0.007237f
C385 B.n345 VSUBS 0.008948f
C386 B.n346 VSUBS 0.008948f
C387 B.n347 VSUBS 0.008948f
C388 B.n348 VSUBS 0.008948f
C389 B.n349 VSUBS 0.008948f
C390 B.n350 VSUBS 0.008948f
C391 B.n351 VSUBS 0.008948f
C392 B.n352 VSUBS 0.008948f
C393 B.n353 VSUBS 0.008948f
C394 B.n354 VSUBS 0.008948f
C395 B.n355 VSUBS 0.008948f
C396 B.n356 VSUBS 0.008948f
C397 B.n357 VSUBS 0.008948f
C398 B.n358 VSUBS 0.008948f
C399 B.n359 VSUBS 0.008948f
C400 B.n360 VSUBS 0.008948f
C401 B.n361 VSUBS 0.008948f
C402 B.n362 VSUBS 0.008948f
C403 B.n363 VSUBS 0.008948f
C404 B.n364 VSUBS 0.008948f
C405 B.n365 VSUBS 0.008948f
C406 B.n366 VSUBS 0.008948f
C407 B.n367 VSUBS 0.008948f
C408 B.n368 VSUBS 0.008948f
C409 B.n369 VSUBS 0.008948f
C410 B.n370 VSUBS 0.008948f
C411 B.n371 VSUBS 0.008948f
C412 B.n372 VSUBS 0.008948f
C413 B.n373 VSUBS 0.008948f
C414 B.n374 VSUBS 0.008948f
C415 B.n375 VSUBS 0.008948f
C416 B.n376 VSUBS 0.008948f
C417 B.n377 VSUBS 0.008948f
C418 B.n378 VSUBS 0.008948f
C419 B.n379 VSUBS 0.008948f
C420 B.n380 VSUBS 0.008948f
C421 B.n381 VSUBS 0.008948f
C422 B.n382 VSUBS 0.008948f
C423 B.n383 VSUBS 0.008948f
C424 B.n384 VSUBS 0.008948f
C425 B.n385 VSUBS 0.008948f
C426 B.n386 VSUBS 0.008948f
C427 B.n387 VSUBS 0.008948f
C428 B.n388 VSUBS 0.008948f
C429 B.n389 VSUBS 0.008948f
C430 B.n390 VSUBS 0.008948f
C431 B.n391 VSUBS 0.008948f
C432 B.n392 VSUBS 0.008948f
C433 B.n393 VSUBS 0.008948f
C434 B.n394 VSUBS 0.008948f
C435 B.n395 VSUBS 0.008948f
C436 B.n396 VSUBS 0.008948f
C437 B.n397 VSUBS 0.008948f
C438 B.n398 VSUBS 0.008948f
C439 B.n399 VSUBS 0.008948f
C440 B.n400 VSUBS 0.008948f
C441 B.n401 VSUBS 0.008948f
C442 B.n402 VSUBS 0.008948f
C443 B.n403 VSUBS 0.020584f
C444 B.n404 VSUBS 0.019681f
C445 B.n405 VSUBS 0.019681f
C446 B.n406 VSUBS 0.008948f
C447 B.n407 VSUBS 0.008948f
C448 B.n408 VSUBS 0.008948f
C449 B.n409 VSUBS 0.008948f
C450 B.n410 VSUBS 0.008948f
C451 B.n411 VSUBS 0.008948f
C452 B.n412 VSUBS 0.008948f
C453 B.n413 VSUBS 0.008948f
C454 B.n414 VSUBS 0.008948f
C455 B.n415 VSUBS 0.008948f
C456 B.n416 VSUBS 0.008948f
C457 B.n417 VSUBS 0.008948f
C458 B.n418 VSUBS 0.008948f
C459 B.n419 VSUBS 0.008948f
C460 B.n420 VSUBS 0.008948f
C461 B.n421 VSUBS 0.008948f
C462 B.n422 VSUBS 0.008948f
C463 B.n423 VSUBS 0.008948f
C464 B.n424 VSUBS 0.008948f
C465 B.n425 VSUBS 0.008948f
C466 B.n426 VSUBS 0.008948f
C467 B.n427 VSUBS 0.008948f
C468 B.n428 VSUBS 0.008948f
C469 B.n429 VSUBS 0.008948f
C470 B.n430 VSUBS 0.008948f
C471 B.n431 VSUBS 0.008948f
C472 B.n432 VSUBS 0.008948f
C473 B.n433 VSUBS 0.008948f
C474 B.n434 VSUBS 0.008948f
C475 B.n435 VSUBS 0.008948f
C476 B.n436 VSUBS 0.008948f
C477 B.n437 VSUBS 0.008948f
C478 B.n438 VSUBS 0.008948f
C479 B.n439 VSUBS 0.008948f
C480 B.n440 VSUBS 0.008948f
C481 B.n441 VSUBS 0.008948f
C482 B.n442 VSUBS 0.008948f
C483 B.n443 VSUBS 0.008948f
C484 B.n444 VSUBS 0.008948f
C485 B.n445 VSUBS 0.008948f
C486 B.n446 VSUBS 0.008948f
C487 B.n447 VSUBS 0.008948f
C488 B.n448 VSUBS 0.008948f
C489 B.n449 VSUBS 0.008948f
C490 B.n450 VSUBS 0.008948f
C491 B.n451 VSUBS 0.008948f
C492 B.n452 VSUBS 0.008948f
C493 B.n453 VSUBS 0.008948f
C494 B.n454 VSUBS 0.008948f
C495 B.n455 VSUBS 0.008948f
C496 B.n456 VSUBS 0.008948f
C497 B.n457 VSUBS 0.008948f
C498 B.n458 VSUBS 0.008948f
C499 B.n459 VSUBS 0.008948f
C500 B.n460 VSUBS 0.008948f
C501 B.n461 VSUBS 0.008948f
C502 B.n462 VSUBS 0.008948f
C503 B.n463 VSUBS 0.008948f
C504 B.n464 VSUBS 0.008948f
C505 B.n465 VSUBS 0.008948f
C506 B.n466 VSUBS 0.008948f
C507 B.n467 VSUBS 0.008948f
C508 B.n468 VSUBS 0.008948f
C509 B.n469 VSUBS 0.008948f
C510 B.n470 VSUBS 0.008948f
C511 B.n471 VSUBS 0.008948f
C512 B.n472 VSUBS 0.008948f
C513 B.n473 VSUBS 0.008948f
C514 B.n474 VSUBS 0.008948f
C515 B.n475 VSUBS 0.008948f
C516 B.n476 VSUBS 0.008948f
C517 B.n477 VSUBS 0.008948f
C518 B.n478 VSUBS 0.008948f
C519 B.n479 VSUBS 0.008948f
C520 B.n480 VSUBS 0.008948f
C521 B.n481 VSUBS 0.008948f
C522 B.n482 VSUBS 0.008948f
C523 B.n483 VSUBS 0.008948f
C524 B.n484 VSUBS 0.008948f
C525 B.n485 VSUBS 0.008948f
C526 B.n486 VSUBS 0.008948f
C527 B.n487 VSUBS 0.008948f
C528 B.n488 VSUBS 0.008948f
C529 B.n489 VSUBS 0.008948f
C530 B.n490 VSUBS 0.008948f
C531 B.n491 VSUBS 0.008948f
C532 B.n492 VSUBS 0.008948f
C533 B.n493 VSUBS 0.008948f
C534 B.n494 VSUBS 0.008948f
C535 B.n495 VSUBS 0.008948f
C536 B.n496 VSUBS 0.008948f
C537 B.n497 VSUBS 0.008948f
C538 B.n498 VSUBS 0.008948f
C539 B.n499 VSUBS 0.008948f
C540 B.n500 VSUBS 0.008948f
C541 B.n501 VSUBS 0.008948f
C542 B.n502 VSUBS 0.008948f
C543 B.n503 VSUBS 0.008948f
C544 B.n504 VSUBS 0.008948f
C545 B.n505 VSUBS 0.008948f
C546 B.n506 VSUBS 0.008948f
C547 B.n507 VSUBS 0.008948f
C548 B.n508 VSUBS 0.008948f
C549 B.n509 VSUBS 0.008948f
C550 B.n510 VSUBS 0.008948f
C551 B.n511 VSUBS 0.008948f
C552 B.n512 VSUBS 0.008948f
C553 B.n513 VSUBS 0.008948f
C554 B.n514 VSUBS 0.008948f
C555 B.n515 VSUBS 0.008948f
C556 B.n516 VSUBS 0.008948f
C557 B.n517 VSUBS 0.008948f
C558 B.n518 VSUBS 0.008948f
C559 B.n519 VSUBS 0.008948f
C560 B.n520 VSUBS 0.008948f
C561 B.n521 VSUBS 0.008948f
C562 B.n522 VSUBS 0.008948f
C563 B.n523 VSUBS 0.008948f
C564 B.n524 VSUBS 0.008948f
C565 B.n525 VSUBS 0.008948f
C566 B.n526 VSUBS 0.008948f
C567 B.n527 VSUBS 0.008948f
C568 B.n528 VSUBS 0.008948f
C569 B.n529 VSUBS 0.008948f
C570 B.n530 VSUBS 0.008948f
C571 B.n531 VSUBS 0.008948f
C572 B.n532 VSUBS 0.008948f
C573 B.n533 VSUBS 0.008948f
C574 B.n534 VSUBS 0.008948f
C575 B.n535 VSUBS 0.008948f
C576 B.n536 VSUBS 0.008948f
C577 B.n537 VSUBS 0.008948f
C578 B.n538 VSUBS 0.008948f
C579 B.n539 VSUBS 0.008948f
C580 B.n540 VSUBS 0.008948f
C581 B.n541 VSUBS 0.008948f
C582 B.n542 VSUBS 0.008948f
C583 B.n543 VSUBS 0.008948f
C584 B.n544 VSUBS 0.008948f
C585 B.n545 VSUBS 0.008948f
C586 B.n546 VSUBS 0.008948f
C587 B.n547 VSUBS 0.008948f
C588 B.n548 VSUBS 0.008948f
C589 B.n549 VSUBS 0.008948f
C590 B.n550 VSUBS 0.008948f
C591 B.n551 VSUBS 0.008948f
C592 B.n552 VSUBS 0.008948f
C593 B.n553 VSUBS 0.008948f
C594 B.n554 VSUBS 0.020803f
C595 B.n555 VSUBS 0.019681f
C596 B.n556 VSUBS 0.020584f
C597 B.n557 VSUBS 0.008948f
C598 B.n558 VSUBS 0.008948f
C599 B.n559 VSUBS 0.008948f
C600 B.n560 VSUBS 0.008948f
C601 B.n561 VSUBS 0.008948f
C602 B.n562 VSUBS 0.008948f
C603 B.n563 VSUBS 0.008948f
C604 B.n564 VSUBS 0.008948f
C605 B.n565 VSUBS 0.008948f
C606 B.n566 VSUBS 0.008948f
C607 B.n567 VSUBS 0.008948f
C608 B.n568 VSUBS 0.008948f
C609 B.n569 VSUBS 0.008948f
C610 B.n570 VSUBS 0.008948f
C611 B.n571 VSUBS 0.008948f
C612 B.n572 VSUBS 0.008948f
C613 B.n573 VSUBS 0.008948f
C614 B.n574 VSUBS 0.008948f
C615 B.n575 VSUBS 0.008948f
C616 B.n576 VSUBS 0.008948f
C617 B.n577 VSUBS 0.008948f
C618 B.n578 VSUBS 0.008948f
C619 B.n579 VSUBS 0.008948f
C620 B.n580 VSUBS 0.008948f
C621 B.n581 VSUBS 0.008948f
C622 B.n582 VSUBS 0.008948f
C623 B.n583 VSUBS 0.008948f
C624 B.n584 VSUBS 0.008948f
C625 B.n585 VSUBS 0.008948f
C626 B.n586 VSUBS 0.008948f
C627 B.n587 VSUBS 0.008948f
C628 B.n588 VSUBS 0.008948f
C629 B.n589 VSUBS 0.008948f
C630 B.n590 VSUBS 0.008948f
C631 B.n591 VSUBS 0.008948f
C632 B.n592 VSUBS 0.008948f
C633 B.n593 VSUBS 0.008948f
C634 B.n594 VSUBS 0.008948f
C635 B.n595 VSUBS 0.008948f
C636 B.n596 VSUBS 0.008948f
C637 B.n597 VSUBS 0.008948f
C638 B.n598 VSUBS 0.008948f
C639 B.n599 VSUBS 0.008948f
C640 B.n600 VSUBS 0.008948f
C641 B.n601 VSUBS 0.008948f
C642 B.n602 VSUBS 0.008948f
C643 B.n603 VSUBS 0.008948f
C644 B.n604 VSUBS 0.008948f
C645 B.n605 VSUBS 0.008948f
C646 B.n606 VSUBS 0.008948f
C647 B.n607 VSUBS 0.008948f
C648 B.n608 VSUBS 0.008948f
C649 B.n609 VSUBS 0.008948f
C650 B.n610 VSUBS 0.008948f
C651 B.n611 VSUBS 0.008948f
C652 B.n612 VSUBS 0.008948f
C653 B.n613 VSUBS 0.006185f
C654 B.n614 VSUBS 0.020731f
C655 B.n615 VSUBS 0.007237f
C656 B.n616 VSUBS 0.008948f
C657 B.n617 VSUBS 0.008948f
C658 B.n618 VSUBS 0.008948f
C659 B.n619 VSUBS 0.008948f
C660 B.n620 VSUBS 0.008948f
C661 B.n621 VSUBS 0.008948f
C662 B.n622 VSUBS 0.008948f
C663 B.n623 VSUBS 0.008948f
C664 B.n624 VSUBS 0.008948f
C665 B.n625 VSUBS 0.008948f
C666 B.n626 VSUBS 0.008948f
C667 B.n627 VSUBS 0.007237f
C668 B.n628 VSUBS 0.008948f
C669 B.n629 VSUBS 0.008948f
C670 B.n630 VSUBS 0.008948f
C671 B.n631 VSUBS 0.008948f
C672 B.n632 VSUBS 0.008948f
C673 B.n633 VSUBS 0.008948f
C674 B.n634 VSUBS 0.008948f
C675 B.n635 VSUBS 0.008948f
C676 B.n636 VSUBS 0.008948f
C677 B.n637 VSUBS 0.008948f
C678 B.n638 VSUBS 0.008948f
C679 B.n639 VSUBS 0.008948f
C680 B.n640 VSUBS 0.008948f
C681 B.n641 VSUBS 0.008948f
C682 B.n642 VSUBS 0.008948f
C683 B.n643 VSUBS 0.008948f
C684 B.n644 VSUBS 0.008948f
C685 B.n645 VSUBS 0.008948f
C686 B.n646 VSUBS 0.008948f
C687 B.n647 VSUBS 0.008948f
C688 B.n648 VSUBS 0.008948f
C689 B.n649 VSUBS 0.008948f
C690 B.n650 VSUBS 0.008948f
C691 B.n651 VSUBS 0.008948f
C692 B.n652 VSUBS 0.008948f
C693 B.n653 VSUBS 0.008948f
C694 B.n654 VSUBS 0.008948f
C695 B.n655 VSUBS 0.008948f
C696 B.n656 VSUBS 0.008948f
C697 B.n657 VSUBS 0.008948f
C698 B.n658 VSUBS 0.008948f
C699 B.n659 VSUBS 0.008948f
C700 B.n660 VSUBS 0.008948f
C701 B.n661 VSUBS 0.008948f
C702 B.n662 VSUBS 0.008948f
C703 B.n663 VSUBS 0.008948f
C704 B.n664 VSUBS 0.008948f
C705 B.n665 VSUBS 0.008948f
C706 B.n666 VSUBS 0.008948f
C707 B.n667 VSUBS 0.008948f
C708 B.n668 VSUBS 0.008948f
C709 B.n669 VSUBS 0.008948f
C710 B.n670 VSUBS 0.008948f
C711 B.n671 VSUBS 0.008948f
C712 B.n672 VSUBS 0.008948f
C713 B.n673 VSUBS 0.008948f
C714 B.n674 VSUBS 0.008948f
C715 B.n675 VSUBS 0.008948f
C716 B.n676 VSUBS 0.008948f
C717 B.n677 VSUBS 0.008948f
C718 B.n678 VSUBS 0.008948f
C719 B.n679 VSUBS 0.008948f
C720 B.n680 VSUBS 0.008948f
C721 B.n681 VSUBS 0.008948f
C722 B.n682 VSUBS 0.008948f
C723 B.n683 VSUBS 0.008948f
C724 B.n684 VSUBS 0.008948f
C725 B.n685 VSUBS 0.008948f
C726 B.n686 VSUBS 0.020584f
C727 B.n687 VSUBS 0.019681f
C728 B.n688 VSUBS 0.019681f
C729 B.n689 VSUBS 0.008948f
C730 B.n690 VSUBS 0.008948f
C731 B.n691 VSUBS 0.008948f
C732 B.n692 VSUBS 0.008948f
C733 B.n693 VSUBS 0.008948f
C734 B.n694 VSUBS 0.008948f
C735 B.n695 VSUBS 0.008948f
C736 B.n696 VSUBS 0.008948f
C737 B.n697 VSUBS 0.008948f
C738 B.n698 VSUBS 0.008948f
C739 B.n699 VSUBS 0.008948f
C740 B.n700 VSUBS 0.008948f
C741 B.n701 VSUBS 0.008948f
C742 B.n702 VSUBS 0.008948f
C743 B.n703 VSUBS 0.008948f
C744 B.n704 VSUBS 0.008948f
C745 B.n705 VSUBS 0.008948f
C746 B.n706 VSUBS 0.008948f
C747 B.n707 VSUBS 0.008948f
C748 B.n708 VSUBS 0.008948f
C749 B.n709 VSUBS 0.008948f
C750 B.n710 VSUBS 0.008948f
C751 B.n711 VSUBS 0.008948f
C752 B.n712 VSUBS 0.008948f
C753 B.n713 VSUBS 0.008948f
C754 B.n714 VSUBS 0.008948f
C755 B.n715 VSUBS 0.008948f
C756 B.n716 VSUBS 0.008948f
C757 B.n717 VSUBS 0.008948f
C758 B.n718 VSUBS 0.008948f
C759 B.n719 VSUBS 0.008948f
C760 B.n720 VSUBS 0.008948f
C761 B.n721 VSUBS 0.008948f
C762 B.n722 VSUBS 0.008948f
C763 B.n723 VSUBS 0.008948f
C764 B.n724 VSUBS 0.008948f
C765 B.n725 VSUBS 0.008948f
C766 B.n726 VSUBS 0.008948f
C767 B.n727 VSUBS 0.008948f
C768 B.n728 VSUBS 0.008948f
C769 B.n729 VSUBS 0.008948f
C770 B.n730 VSUBS 0.008948f
C771 B.n731 VSUBS 0.008948f
C772 B.n732 VSUBS 0.008948f
C773 B.n733 VSUBS 0.008948f
C774 B.n734 VSUBS 0.008948f
C775 B.n735 VSUBS 0.008948f
C776 B.n736 VSUBS 0.008948f
C777 B.n737 VSUBS 0.008948f
C778 B.n738 VSUBS 0.008948f
C779 B.n739 VSUBS 0.008948f
C780 B.n740 VSUBS 0.008948f
C781 B.n741 VSUBS 0.008948f
C782 B.n742 VSUBS 0.008948f
C783 B.n743 VSUBS 0.008948f
C784 B.n744 VSUBS 0.008948f
C785 B.n745 VSUBS 0.008948f
C786 B.n746 VSUBS 0.008948f
C787 B.n747 VSUBS 0.008948f
C788 B.n748 VSUBS 0.008948f
C789 B.n749 VSUBS 0.008948f
C790 B.n750 VSUBS 0.008948f
C791 B.n751 VSUBS 0.008948f
C792 B.n752 VSUBS 0.008948f
C793 B.n753 VSUBS 0.008948f
C794 B.n754 VSUBS 0.008948f
C795 B.n755 VSUBS 0.008948f
C796 B.n756 VSUBS 0.008948f
C797 B.n757 VSUBS 0.008948f
C798 B.n758 VSUBS 0.008948f
C799 B.n759 VSUBS 0.008948f
C800 B.n760 VSUBS 0.008948f
C801 B.n761 VSUBS 0.008948f
C802 B.n762 VSUBS 0.008948f
C803 B.n763 VSUBS 0.020261f
C804 VDD1.t5 VSUBS 2.53722f
C805 VDD1.t3 VSUBS 2.53574f
C806 VDD1.t2 VSUBS 0.250182f
C807 VDD1.t4 VSUBS 0.250182f
C808 VDD1.n0 VSUBS 1.92787f
C809 VDD1.n1 VSUBS 4.34433f
C810 VDD1.t0 VSUBS 0.250182f
C811 VDD1.t1 VSUBS 0.250182f
C812 VDD1.n2 VSUBS 1.91941f
C813 VDD1.n3 VSUBS 3.6222f
C814 VP.t1 VSUBS 2.97282f
C815 VP.n0 VSUBS 1.16827f
C816 VP.n1 VSUBS 0.030885f
C817 VP.n2 VSUBS 0.025191f
C818 VP.n3 VSUBS 0.030885f
C819 VP.t3 VSUBS 2.97282f
C820 VP.n4 VSUBS 1.05018f
C821 VP.n5 VSUBS 0.030885f
C822 VP.n6 VSUBS 0.025191f
C823 VP.n7 VSUBS 0.030885f
C824 VP.t2 VSUBS 2.97282f
C825 VP.n8 VSUBS 1.16827f
C826 VP.t4 VSUBS 2.97282f
C827 VP.n9 VSUBS 1.16827f
C828 VP.n10 VSUBS 0.030885f
C829 VP.n11 VSUBS 0.025191f
C830 VP.n12 VSUBS 0.030885f
C831 VP.t5 VSUBS 2.97282f
C832 VP.n13 VSUBS 1.15143f
C833 VP.t0 VSUBS 3.3355f
C834 VP.n14 VSUBS 1.09599f
C835 VP.n15 VSUBS 0.35974f
C836 VP.n16 VSUBS 0.043136f
C837 VP.n17 VSUBS 0.057273f
C838 VP.n18 VSUBS 0.061695f
C839 VP.n19 VSUBS 0.030885f
C840 VP.n20 VSUBS 0.030885f
C841 VP.n21 VSUBS 0.030885f
C842 VP.n22 VSUBS 0.060178f
C843 VP.n23 VSUBS 0.057273f
C844 VP.n24 VSUBS 0.045963f
C845 VP.n25 VSUBS 0.049839f
C846 VP.n26 VSUBS 1.77744f
C847 VP.n27 VSUBS 1.79951f
C848 VP.n28 VSUBS 0.049839f
C849 VP.n29 VSUBS 0.045963f
C850 VP.n30 VSUBS 0.057273f
C851 VP.n31 VSUBS 0.060178f
C852 VP.n32 VSUBS 0.030885f
C853 VP.n33 VSUBS 0.030885f
C854 VP.n34 VSUBS 0.030885f
C855 VP.n35 VSUBS 0.061695f
C856 VP.n36 VSUBS 0.057273f
C857 VP.n37 VSUBS 0.043136f
C858 VP.n38 VSUBS 0.030885f
C859 VP.n39 VSUBS 0.030885f
C860 VP.n40 VSUBS 0.043136f
C861 VP.n41 VSUBS 0.057273f
C862 VP.n42 VSUBS 0.061695f
C863 VP.n43 VSUBS 0.030885f
C864 VP.n44 VSUBS 0.030885f
C865 VP.n45 VSUBS 0.030885f
C866 VP.n46 VSUBS 0.060178f
C867 VP.n47 VSUBS 0.057273f
C868 VP.n48 VSUBS 0.045963f
C869 VP.n49 VSUBS 0.049839f
C870 VP.n50 VSUBS 0.073651f
C871 VTAIL.t6 VSUBS 0.261679f
C872 VTAIL.t5 VSUBS 0.261679f
C873 VTAIL.n0 VSUBS 1.84814f
C874 VTAIL.n1 VSUBS 0.951325f
C875 VTAIL.t3 VSUBS 2.45002f
C876 VTAIL.n2 VSUBS 1.28011f
C877 VTAIL.t1 VSUBS 0.261679f
C878 VTAIL.t4 VSUBS 0.261679f
C879 VTAIL.n3 VSUBS 1.84814f
C880 VTAIL.n4 VSUBS 2.8968f
C881 VTAIL.t7 VSUBS 0.261679f
C882 VTAIL.t10 VSUBS 0.261679f
C883 VTAIL.n5 VSUBS 1.84814f
C884 VTAIL.n6 VSUBS 2.8968f
C885 VTAIL.t8 VSUBS 2.45004f
C886 VTAIL.n7 VSUBS 1.28009f
C887 VTAIL.t2 VSUBS 0.261679f
C888 VTAIL.t0 VSUBS 0.261679f
C889 VTAIL.n8 VSUBS 1.84814f
C890 VTAIL.n9 VSUBS 1.16832f
C891 VTAIL.t11 VSUBS 2.45002f
C892 VTAIL.n10 VSUBS 2.71173f
C893 VTAIL.t9 VSUBS 2.45002f
C894 VTAIL.n11 VSUBS 2.63187f
C895 VDD2.t5 VSUBS 2.52317f
C896 VDD2.t3 VSUBS 0.248941f
C897 VDD2.t4 VSUBS 0.248941f
C898 VDD2.n0 VSUBS 1.91831f
C899 VDD2.n1 VSUBS 4.16286f
C900 VDD2.t2 VSUBS 2.49959f
C901 VDD2.n2 VSUBS 3.61714f
C902 VDD2.t1 VSUBS 0.248941f
C903 VDD2.t0 VSUBS 0.248941f
C904 VDD2.n3 VSUBS 1.91826f
C905 VN.t1 VSUBS 2.67948f
C906 VN.n0 VSUBS 1.05299f
C907 VN.n1 VSUBS 0.027837f
C908 VN.n2 VSUBS 0.022706f
C909 VN.n3 VSUBS 0.027837f
C910 VN.t5 VSUBS 2.67948f
C911 VN.n4 VSUBS 1.03781f
C912 VN.t4 VSUBS 3.00638f
C913 VN.n5 VSUBS 0.987843f
C914 VN.n6 VSUBS 0.324243f
C915 VN.n7 VSUBS 0.038879f
C916 VN.n8 VSUBS 0.051621f
C917 VN.n9 VSUBS 0.055607f
C918 VN.n10 VSUBS 0.027837f
C919 VN.n11 VSUBS 0.027837f
C920 VN.n12 VSUBS 0.027837f
C921 VN.n13 VSUBS 0.05424f
C922 VN.n14 VSUBS 0.051621f
C923 VN.n15 VSUBS 0.041428f
C924 VN.n16 VSUBS 0.044922f
C925 VN.n17 VSUBS 0.066383f
C926 VN.t3 VSUBS 2.67948f
C927 VN.n18 VSUBS 1.05299f
C928 VN.n19 VSUBS 0.027837f
C929 VN.n20 VSUBS 0.022706f
C930 VN.n21 VSUBS 0.027837f
C931 VN.t0 VSUBS 2.67948f
C932 VN.n22 VSUBS 1.03781f
C933 VN.t2 VSUBS 3.00638f
C934 VN.n23 VSUBS 0.987843f
C935 VN.n24 VSUBS 0.324243f
C936 VN.n25 VSUBS 0.038879f
C937 VN.n26 VSUBS 0.051621f
C938 VN.n27 VSUBS 0.055607f
C939 VN.n28 VSUBS 0.027837f
C940 VN.n29 VSUBS 0.027837f
C941 VN.n30 VSUBS 0.027837f
C942 VN.n31 VSUBS 0.05424f
C943 VN.n32 VSUBS 0.051621f
C944 VN.n33 VSUBS 0.041428f
C945 VN.n34 VSUBS 0.044922f
C946 VN.n35 VSUBS 1.61341f
.ends

