* NGSPICE file created from diff_pair_sample_1066.ext - technology: sky130A

.subckt diff_pair_sample_1066 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t11 VN.t0 VDD2.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=0.7425 pd=4.83 as=0.7425 ps=4.83 w=4.5 l=2.34
X1 VTAIL.t2 VP.t0 VDD1.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=0.7425 pd=4.83 as=0.7425 ps=4.83 w=4.5 l=2.34
X2 B.t19 B.t17 B.t18 B.t7 sky130_fd_pr__nfet_01v8 ad=1.755 pd=9.78 as=0 ps=0 w=4.5 l=2.34
X3 VTAIL.t10 VN.t1 VDD2.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.7425 pd=4.83 as=0.7425 ps=4.83 w=4.5 l=2.34
X4 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=1.755 pd=9.78 as=0 ps=0 w=4.5 l=2.34
X5 VDD1.t4 VP.t1 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=0.7425 pd=4.83 as=1.755 ps=9.78 w=4.5 l=2.34
X6 VDD1.t3 VP.t2 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.7425 pd=4.83 as=1.755 ps=9.78 w=4.5 l=2.34
X7 VDD1.t2 VP.t3 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.755 pd=9.78 as=0.7425 ps=4.83 w=4.5 l=2.34
X8 VDD1.t1 VP.t4 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.755 pd=9.78 as=0.7425 ps=4.83 w=4.5 l=2.34
X9 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=1.755 pd=9.78 as=0 ps=0 w=4.5 l=2.34
X10 VDD2.t0 VN.t2 VTAIL.t9 B.t0 sky130_fd_pr__nfet_01v8 ad=0.7425 pd=4.83 as=1.755 ps=9.78 w=4.5 l=2.34
X11 VTAIL.t3 VP.t5 VDD1.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=0.7425 pd=4.83 as=0.7425 ps=4.83 w=4.5 l=2.34
X12 VDD2.t4 VN.t3 VTAIL.t8 B.t4 sky130_fd_pr__nfet_01v8 ad=1.755 pd=9.78 as=0.7425 ps=4.83 w=4.5 l=2.34
X13 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=1.755 pd=9.78 as=0 ps=0 w=4.5 l=2.34
X14 VDD2.t2 VN.t4 VTAIL.t7 B.t5 sky130_fd_pr__nfet_01v8 ad=0.7425 pd=4.83 as=1.755 ps=9.78 w=4.5 l=2.34
X15 VDD2.t5 VN.t5 VTAIL.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=1.755 pd=9.78 as=0.7425 ps=4.83 w=4.5 l=2.34
R0 VN.n25 VN.n14 161.3
R1 VN.n24 VN.n23 161.3
R2 VN.n22 VN.n15 161.3
R3 VN.n21 VN.n20 161.3
R4 VN.n19 VN.n16 161.3
R5 VN.n11 VN.n0 161.3
R6 VN.n10 VN.n9 161.3
R7 VN.n8 VN.n1 161.3
R8 VN.n7 VN.n6 161.3
R9 VN.n5 VN.n2 161.3
R10 VN.n13 VN.n12 102.547
R11 VN.n27 VN.n26 102.547
R12 VN.n3 VN.t5 79.5466
R13 VN.n17 VN.t2 79.5466
R14 VN.n6 VN.n1 56.5617
R15 VN.n20 VN.n15 56.5617
R16 VN.n18 VN.n17 47.9848
R17 VN.n4 VN.n3 47.9848
R18 VN.n4 VN.t1 46.3467
R19 VN.n12 VN.t4 46.3467
R20 VN.n18 VN.t0 46.3467
R21 VN.n26 VN.t3 46.3467
R22 VN VN.n27 42.1838
R23 VN.n5 VN.n4 24.5923
R24 VN.n6 VN.n5 24.5923
R25 VN.n10 VN.n1 24.5923
R26 VN.n11 VN.n10 24.5923
R27 VN.n20 VN.n19 24.5923
R28 VN.n19 VN.n18 24.5923
R29 VN.n25 VN.n24 24.5923
R30 VN.n24 VN.n15 24.5923
R31 VN.n12 VN.n11 8.36172
R32 VN.n26 VN.n25 8.36172
R33 VN.n17 VN.n16 6.93618
R34 VN.n3 VN.n2 6.93618
R35 VN.n27 VN.n14 0.278335
R36 VN.n13 VN.n0 0.278335
R37 VN.n23 VN.n14 0.189894
R38 VN.n23 VN.n22 0.189894
R39 VN.n22 VN.n21 0.189894
R40 VN.n21 VN.n16 0.189894
R41 VN.n7 VN.n2 0.189894
R42 VN.n8 VN.n7 0.189894
R43 VN.n9 VN.n8 0.189894
R44 VN.n9 VN.n0 0.189894
R45 VN VN.n13 0.153485
R46 VDD2.n43 VDD2.n25 289.615
R47 VDD2.n18 VDD2.n0 289.615
R48 VDD2.n44 VDD2.n43 185
R49 VDD2.n42 VDD2.n41 185
R50 VDD2.n29 VDD2.n28 185
R51 VDD2.n36 VDD2.n35 185
R52 VDD2.n34 VDD2.n33 185
R53 VDD2.n9 VDD2.n8 185
R54 VDD2.n11 VDD2.n10 185
R55 VDD2.n4 VDD2.n3 185
R56 VDD2.n17 VDD2.n16 185
R57 VDD2.n19 VDD2.n18 185
R58 VDD2.n32 VDD2.t4 147.714
R59 VDD2.n7 VDD2.t5 147.714
R60 VDD2.n43 VDD2.n42 104.615
R61 VDD2.n42 VDD2.n28 104.615
R62 VDD2.n35 VDD2.n28 104.615
R63 VDD2.n35 VDD2.n34 104.615
R64 VDD2.n10 VDD2.n9 104.615
R65 VDD2.n10 VDD2.n3 104.615
R66 VDD2.n17 VDD2.n3 104.615
R67 VDD2.n18 VDD2.n17 104.615
R68 VDD2.n24 VDD2.n23 69.9981
R69 VDD2 VDD2.n49 69.9953
R70 VDD2.n34 VDD2.t4 52.3082
R71 VDD2.n9 VDD2.t5 52.3082
R72 VDD2.n24 VDD2.n22 49.3714
R73 VDD2.n48 VDD2.n47 47.7005
R74 VDD2.n48 VDD2.n24 35.0752
R75 VDD2.n33 VDD2.n32 15.6631
R76 VDD2.n8 VDD2.n7 15.6631
R77 VDD2.n36 VDD2.n31 12.8005
R78 VDD2.n11 VDD2.n6 12.8005
R79 VDD2.n37 VDD2.n29 12.0247
R80 VDD2.n12 VDD2.n4 12.0247
R81 VDD2.n41 VDD2.n40 11.249
R82 VDD2.n16 VDD2.n15 11.249
R83 VDD2.n44 VDD2.n27 10.4732
R84 VDD2.n19 VDD2.n2 10.4732
R85 VDD2.n45 VDD2.n25 9.69747
R86 VDD2.n20 VDD2.n0 9.69747
R87 VDD2.n47 VDD2.n46 9.45567
R88 VDD2.n22 VDD2.n21 9.45567
R89 VDD2.n46 VDD2.n45 9.3005
R90 VDD2.n27 VDD2.n26 9.3005
R91 VDD2.n40 VDD2.n39 9.3005
R92 VDD2.n38 VDD2.n37 9.3005
R93 VDD2.n31 VDD2.n30 9.3005
R94 VDD2.n21 VDD2.n20 9.3005
R95 VDD2.n2 VDD2.n1 9.3005
R96 VDD2.n15 VDD2.n14 9.3005
R97 VDD2.n13 VDD2.n12 9.3005
R98 VDD2.n6 VDD2.n5 9.3005
R99 VDD2.n49 VDD2.t1 4.4005
R100 VDD2.n49 VDD2.t0 4.4005
R101 VDD2.n23 VDD2.t3 4.4005
R102 VDD2.n23 VDD2.t2 4.4005
R103 VDD2.n32 VDD2.n30 4.39059
R104 VDD2.n7 VDD2.n5 4.39059
R105 VDD2.n47 VDD2.n25 4.26717
R106 VDD2.n22 VDD2.n0 4.26717
R107 VDD2.n45 VDD2.n44 3.49141
R108 VDD2.n20 VDD2.n19 3.49141
R109 VDD2.n41 VDD2.n27 2.71565
R110 VDD2.n16 VDD2.n2 2.71565
R111 VDD2.n40 VDD2.n29 1.93989
R112 VDD2.n15 VDD2.n4 1.93989
R113 VDD2 VDD2.n48 1.78498
R114 VDD2.n37 VDD2.n36 1.16414
R115 VDD2.n12 VDD2.n11 1.16414
R116 VDD2.n33 VDD2.n31 0.388379
R117 VDD2.n8 VDD2.n6 0.388379
R118 VDD2.n46 VDD2.n26 0.155672
R119 VDD2.n39 VDD2.n26 0.155672
R120 VDD2.n39 VDD2.n38 0.155672
R121 VDD2.n38 VDD2.n30 0.155672
R122 VDD2.n13 VDD2.n5 0.155672
R123 VDD2.n14 VDD2.n13 0.155672
R124 VDD2.n14 VDD2.n1 0.155672
R125 VDD2.n21 VDD2.n1 0.155672
R126 VTAIL.n98 VTAIL.n80 289.615
R127 VTAIL.n20 VTAIL.n2 289.615
R128 VTAIL.n74 VTAIL.n56 289.615
R129 VTAIL.n48 VTAIL.n30 289.615
R130 VTAIL.n89 VTAIL.n88 185
R131 VTAIL.n91 VTAIL.n90 185
R132 VTAIL.n84 VTAIL.n83 185
R133 VTAIL.n97 VTAIL.n96 185
R134 VTAIL.n99 VTAIL.n98 185
R135 VTAIL.n11 VTAIL.n10 185
R136 VTAIL.n13 VTAIL.n12 185
R137 VTAIL.n6 VTAIL.n5 185
R138 VTAIL.n19 VTAIL.n18 185
R139 VTAIL.n21 VTAIL.n20 185
R140 VTAIL.n75 VTAIL.n74 185
R141 VTAIL.n73 VTAIL.n72 185
R142 VTAIL.n60 VTAIL.n59 185
R143 VTAIL.n67 VTAIL.n66 185
R144 VTAIL.n65 VTAIL.n64 185
R145 VTAIL.n49 VTAIL.n48 185
R146 VTAIL.n47 VTAIL.n46 185
R147 VTAIL.n34 VTAIL.n33 185
R148 VTAIL.n41 VTAIL.n40 185
R149 VTAIL.n39 VTAIL.n38 185
R150 VTAIL.n87 VTAIL.t7 147.714
R151 VTAIL.n9 VTAIL.t0 147.714
R152 VTAIL.n63 VTAIL.t5 147.714
R153 VTAIL.n37 VTAIL.t9 147.714
R154 VTAIL.n90 VTAIL.n89 104.615
R155 VTAIL.n90 VTAIL.n83 104.615
R156 VTAIL.n97 VTAIL.n83 104.615
R157 VTAIL.n98 VTAIL.n97 104.615
R158 VTAIL.n12 VTAIL.n11 104.615
R159 VTAIL.n12 VTAIL.n5 104.615
R160 VTAIL.n19 VTAIL.n5 104.615
R161 VTAIL.n20 VTAIL.n19 104.615
R162 VTAIL.n74 VTAIL.n73 104.615
R163 VTAIL.n73 VTAIL.n59 104.615
R164 VTAIL.n66 VTAIL.n59 104.615
R165 VTAIL.n66 VTAIL.n65 104.615
R166 VTAIL.n48 VTAIL.n47 104.615
R167 VTAIL.n47 VTAIL.n33 104.615
R168 VTAIL.n40 VTAIL.n33 104.615
R169 VTAIL.n40 VTAIL.n39 104.615
R170 VTAIL.n55 VTAIL.n54 52.7994
R171 VTAIL.n29 VTAIL.n28 52.7994
R172 VTAIL.n1 VTAIL.n0 52.7992
R173 VTAIL.n27 VTAIL.n26 52.7992
R174 VTAIL.n89 VTAIL.t7 52.3082
R175 VTAIL.n11 VTAIL.t0 52.3082
R176 VTAIL.n65 VTAIL.t5 52.3082
R177 VTAIL.n39 VTAIL.t9 52.3082
R178 VTAIL.n103 VTAIL.n102 31.0217
R179 VTAIL.n25 VTAIL.n24 31.0217
R180 VTAIL.n79 VTAIL.n78 31.0217
R181 VTAIL.n53 VTAIL.n52 31.0217
R182 VTAIL.n29 VTAIL.n27 20.8496
R183 VTAIL.n103 VTAIL.n79 18.5479
R184 VTAIL.n88 VTAIL.n87 15.6631
R185 VTAIL.n10 VTAIL.n9 15.6631
R186 VTAIL.n64 VTAIL.n63 15.6631
R187 VTAIL.n38 VTAIL.n37 15.6631
R188 VTAIL.n91 VTAIL.n86 12.8005
R189 VTAIL.n13 VTAIL.n8 12.8005
R190 VTAIL.n67 VTAIL.n62 12.8005
R191 VTAIL.n41 VTAIL.n36 12.8005
R192 VTAIL.n92 VTAIL.n84 12.0247
R193 VTAIL.n14 VTAIL.n6 12.0247
R194 VTAIL.n68 VTAIL.n60 12.0247
R195 VTAIL.n42 VTAIL.n34 12.0247
R196 VTAIL.n96 VTAIL.n95 11.249
R197 VTAIL.n18 VTAIL.n17 11.249
R198 VTAIL.n72 VTAIL.n71 11.249
R199 VTAIL.n46 VTAIL.n45 11.249
R200 VTAIL.n99 VTAIL.n82 10.4732
R201 VTAIL.n21 VTAIL.n4 10.4732
R202 VTAIL.n75 VTAIL.n58 10.4732
R203 VTAIL.n49 VTAIL.n32 10.4732
R204 VTAIL.n100 VTAIL.n80 9.69747
R205 VTAIL.n22 VTAIL.n2 9.69747
R206 VTAIL.n76 VTAIL.n56 9.69747
R207 VTAIL.n50 VTAIL.n30 9.69747
R208 VTAIL.n102 VTAIL.n101 9.45567
R209 VTAIL.n24 VTAIL.n23 9.45567
R210 VTAIL.n78 VTAIL.n77 9.45567
R211 VTAIL.n52 VTAIL.n51 9.45567
R212 VTAIL.n101 VTAIL.n100 9.3005
R213 VTAIL.n82 VTAIL.n81 9.3005
R214 VTAIL.n95 VTAIL.n94 9.3005
R215 VTAIL.n93 VTAIL.n92 9.3005
R216 VTAIL.n86 VTAIL.n85 9.3005
R217 VTAIL.n23 VTAIL.n22 9.3005
R218 VTAIL.n4 VTAIL.n3 9.3005
R219 VTAIL.n17 VTAIL.n16 9.3005
R220 VTAIL.n15 VTAIL.n14 9.3005
R221 VTAIL.n8 VTAIL.n7 9.3005
R222 VTAIL.n77 VTAIL.n76 9.3005
R223 VTAIL.n58 VTAIL.n57 9.3005
R224 VTAIL.n71 VTAIL.n70 9.3005
R225 VTAIL.n69 VTAIL.n68 9.3005
R226 VTAIL.n62 VTAIL.n61 9.3005
R227 VTAIL.n51 VTAIL.n50 9.3005
R228 VTAIL.n32 VTAIL.n31 9.3005
R229 VTAIL.n45 VTAIL.n44 9.3005
R230 VTAIL.n43 VTAIL.n42 9.3005
R231 VTAIL.n36 VTAIL.n35 9.3005
R232 VTAIL.n0 VTAIL.t6 4.4005
R233 VTAIL.n0 VTAIL.t10 4.4005
R234 VTAIL.n26 VTAIL.t4 4.4005
R235 VTAIL.n26 VTAIL.t2 4.4005
R236 VTAIL.n54 VTAIL.t1 4.4005
R237 VTAIL.n54 VTAIL.t3 4.4005
R238 VTAIL.n28 VTAIL.t8 4.4005
R239 VTAIL.n28 VTAIL.t11 4.4005
R240 VTAIL.n87 VTAIL.n85 4.39059
R241 VTAIL.n9 VTAIL.n7 4.39059
R242 VTAIL.n63 VTAIL.n61 4.39059
R243 VTAIL.n37 VTAIL.n35 4.39059
R244 VTAIL.n102 VTAIL.n80 4.26717
R245 VTAIL.n24 VTAIL.n2 4.26717
R246 VTAIL.n78 VTAIL.n56 4.26717
R247 VTAIL.n52 VTAIL.n30 4.26717
R248 VTAIL.n100 VTAIL.n99 3.49141
R249 VTAIL.n22 VTAIL.n21 3.49141
R250 VTAIL.n76 VTAIL.n75 3.49141
R251 VTAIL.n50 VTAIL.n49 3.49141
R252 VTAIL.n96 VTAIL.n82 2.71565
R253 VTAIL.n18 VTAIL.n4 2.71565
R254 VTAIL.n72 VTAIL.n58 2.71565
R255 VTAIL.n46 VTAIL.n32 2.71565
R256 VTAIL.n53 VTAIL.n29 2.30222
R257 VTAIL.n79 VTAIL.n55 2.30222
R258 VTAIL.n27 VTAIL.n25 2.30222
R259 VTAIL.n95 VTAIL.n84 1.93989
R260 VTAIL.n17 VTAIL.n6 1.93989
R261 VTAIL.n71 VTAIL.n60 1.93989
R262 VTAIL.n45 VTAIL.n34 1.93989
R263 VTAIL VTAIL.n103 1.6686
R264 VTAIL.n55 VTAIL.n53 1.62119
R265 VTAIL.n25 VTAIL.n1 1.62119
R266 VTAIL.n92 VTAIL.n91 1.16414
R267 VTAIL.n14 VTAIL.n13 1.16414
R268 VTAIL.n68 VTAIL.n67 1.16414
R269 VTAIL.n42 VTAIL.n41 1.16414
R270 VTAIL VTAIL.n1 0.634121
R271 VTAIL.n88 VTAIL.n86 0.388379
R272 VTAIL.n10 VTAIL.n8 0.388379
R273 VTAIL.n64 VTAIL.n62 0.388379
R274 VTAIL.n38 VTAIL.n36 0.388379
R275 VTAIL.n93 VTAIL.n85 0.155672
R276 VTAIL.n94 VTAIL.n93 0.155672
R277 VTAIL.n94 VTAIL.n81 0.155672
R278 VTAIL.n101 VTAIL.n81 0.155672
R279 VTAIL.n15 VTAIL.n7 0.155672
R280 VTAIL.n16 VTAIL.n15 0.155672
R281 VTAIL.n16 VTAIL.n3 0.155672
R282 VTAIL.n23 VTAIL.n3 0.155672
R283 VTAIL.n77 VTAIL.n57 0.155672
R284 VTAIL.n70 VTAIL.n57 0.155672
R285 VTAIL.n70 VTAIL.n69 0.155672
R286 VTAIL.n69 VTAIL.n61 0.155672
R287 VTAIL.n51 VTAIL.n31 0.155672
R288 VTAIL.n44 VTAIL.n31 0.155672
R289 VTAIL.n44 VTAIL.n43 0.155672
R290 VTAIL.n43 VTAIL.n35 0.155672
R291 B.n571 B.n570 585
R292 B.n572 B.n571 585
R293 B.n197 B.n99 585
R294 B.n196 B.n195 585
R295 B.n194 B.n193 585
R296 B.n192 B.n191 585
R297 B.n190 B.n189 585
R298 B.n188 B.n187 585
R299 B.n186 B.n185 585
R300 B.n184 B.n183 585
R301 B.n182 B.n181 585
R302 B.n180 B.n179 585
R303 B.n178 B.n177 585
R304 B.n176 B.n175 585
R305 B.n174 B.n173 585
R306 B.n172 B.n171 585
R307 B.n170 B.n169 585
R308 B.n168 B.n167 585
R309 B.n166 B.n165 585
R310 B.n164 B.n163 585
R311 B.n162 B.n161 585
R312 B.n159 B.n158 585
R313 B.n157 B.n156 585
R314 B.n155 B.n154 585
R315 B.n153 B.n152 585
R316 B.n151 B.n150 585
R317 B.n149 B.n148 585
R318 B.n147 B.n146 585
R319 B.n145 B.n144 585
R320 B.n143 B.n142 585
R321 B.n141 B.n140 585
R322 B.n139 B.n138 585
R323 B.n137 B.n136 585
R324 B.n135 B.n134 585
R325 B.n133 B.n132 585
R326 B.n131 B.n130 585
R327 B.n129 B.n128 585
R328 B.n127 B.n126 585
R329 B.n125 B.n124 585
R330 B.n123 B.n122 585
R331 B.n121 B.n120 585
R332 B.n119 B.n118 585
R333 B.n117 B.n116 585
R334 B.n115 B.n114 585
R335 B.n113 B.n112 585
R336 B.n111 B.n110 585
R337 B.n109 B.n108 585
R338 B.n107 B.n106 585
R339 B.n75 B.n74 585
R340 B.n575 B.n574 585
R341 B.n569 B.n100 585
R342 B.n100 B.n72 585
R343 B.n568 B.n71 585
R344 B.n579 B.n71 585
R345 B.n567 B.n70 585
R346 B.n580 B.n70 585
R347 B.n566 B.n69 585
R348 B.n581 B.n69 585
R349 B.n565 B.n564 585
R350 B.n564 B.n65 585
R351 B.n563 B.n64 585
R352 B.n587 B.n64 585
R353 B.n562 B.n63 585
R354 B.n588 B.n63 585
R355 B.n561 B.n62 585
R356 B.n589 B.n62 585
R357 B.n560 B.n559 585
R358 B.n559 B.n58 585
R359 B.n558 B.n57 585
R360 B.n595 B.n57 585
R361 B.n557 B.n56 585
R362 B.n596 B.n56 585
R363 B.n556 B.n55 585
R364 B.n597 B.n55 585
R365 B.n555 B.n554 585
R366 B.n554 B.n51 585
R367 B.n553 B.n50 585
R368 B.n603 B.n50 585
R369 B.n552 B.n49 585
R370 B.n604 B.n49 585
R371 B.n551 B.n48 585
R372 B.n605 B.n48 585
R373 B.n550 B.n549 585
R374 B.n549 B.n44 585
R375 B.n548 B.n43 585
R376 B.n611 B.n43 585
R377 B.n547 B.n42 585
R378 B.n612 B.n42 585
R379 B.n546 B.n41 585
R380 B.n613 B.n41 585
R381 B.n545 B.n544 585
R382 B.n544 B.n37 585
R383 B.n543 B.n36 585
R384 B.n619 B.n36 585
R385 B.n542 B.n35 585
R386 B.n620 B.n35 585
R387 B.n541 B.n34 585
R388 B.n621 B.n34 585
R389 B.n540 B.n539 585
R390 B.n539 B.n30 585
R391 B.n538 B.n29 585
R392 B.n627 B.n29 585
R393 B.n537 B.n28 585
R394 B.n628 B.n28 585
R395 B.n536 B.n27 585
R396 B.n629 B.n27 585
R397 B.n535 B.n534 585
R398 B.n534 B.n23 585
R399 B.n533 B.n22 585
R400 B.n635 B.n22 585
R401 B.n532 B.n21 585
R402 B.n636 B.n21 585
R403 B.n531 B.n20 585
R404 B.n637 B.n20 585
R405 B.n530 B.n529 585
R406 B.n529 B.n16 585
R407 B.n528 B.n15 585
R408 B.n643 B.n15 585
R409 B.n527 B.n14 585
R410 B.n644 B.n14 585
R411 B.n526 B.n13 585
R412 B.n645 B.n13 585
R413 B.n525 B.n524 585
R414 B.n524 B.n12 585
R415 B.n523 B.n522 585
R416 B.n523 B.n8 585
R417 B.n521 B.n7 585
R418 B.n652 B.n7 585
R419 B.n520 B.n6 585
R420 B.n653 B.n6 585
R421 B.n519 B.n5 585
R422 B.n654 B.n5 585
R423 B.n518 B.n517 585
R424 B.n517 B.n4 585
R425 B.n516 B.n198 585
R426 B.n516 B.n515 585
R427 B.n506 B.n199 585
R428 B.n200 B.n199 585
R429 B.n508 B.n507 585
R430 B.n509 B.n508 585
R431 B.n505 B.n205 585
R432 B.n205 B.n204 585
R433 B.n504 B.n503 585
R434 B.n503 B.n502 585
R435 B.n207 B.n206 585
R436 B.n208 B.n207 585
R437 B.n495 B.n494 585
R438 B.n496 B.n495 585
R439 B.n493 B.n213 585
R440 B.n213 B.n212 585
R441 B.n492 B.n491 585
R442 B.n491 B.n490 585
R443 B.n215 B.n214 585
R444 B.n216 B.n215 585
R445 B.n483 B.n482 585
R446 B.n484 B.n483 585
R447 B.n481 B.n220 585
R448 B.n224 B.n220 585
R449 B.n480 B.n479 585
R450 B.n479 B.n478 585
R451 B.n222 B.n221 585
R452 B.n223 B.n222 585
R453 B.n471 B.n470 585
R454 B.n472 B.n471 585
R455 B.n469 B.n229 585
R456 B.n229 B.n228 585
R457 B.n468 B.n467 585
R458 B.n467 B.n466 585
R459 B.n231 B.n230 585
R460 B.n232 B.n231 585
R461 B.n459 B.n458 585
R462 B.n460 B.n459 585
R463 B.n457 B.n236 585
R464 B.n240 B.n236 585
R465 B.n456 B.n455 585
R466 B.n455 B.n454 585
R467 B.n238 B.n237 585
R468 B.n239 B.n238 585
R469 B.n447 B.n446 585
R470 B.n448 B.n447 585
R471 B.n445 B.n245 585
R472 B.n245 B.n244 585
R473 B.n444 B.n443 585
R474 B.n443 B.n442 585
R475 B.n247 B.n246 585
R476 B.n248 B.n247 585
R477 B.n435 B.n434 585
R478 B.n436 B.n435 585
R479 B.n433 B.n253 585
R480 B.n253 B.n252 585
R481 B.n432 B.n431 585
R482 B.n431 B.n430 585
R483 B.n255 B.n254 585
R484 B.n256 B.n255 585
R485 B.n423 B.n422 585
R486 B.n424 B.n423 585
R487 B.n421 B.n261 585
R488 B.n261 B.n260 585
R489 B.n420 B.n419 585
R490 B.n419 B.n418 585
R491 B.n263 B.n262 585
R492 B.n264 B.n263 585
R493 B.n411 B.n410 585
R494 B.n412 B.n411 585
R495 B.n409 B.n269 585
R496 B.n269 B.n268 585
R497 B.n408 B.n407 585
R498 B.n407 B.n406 585
R499 B.n271 B.n270 585
R500 B.n272 B.n271 585
R501 B.n402 B.n401 585
R502 B.n275 B.n274 585
R503 B.n398 B.n397 585
R504 B.n399 B.n398 585
R505 B.n396 B.n299 585
R506 B.n395 B.n394 585
R507 B.n393 B.n392 585
R508 B.n391 B.n390 585
R509 B.n389 B.n388 585
R510 B.n387 B.n386 585
R511 B.n385 B.n384 585
R512 B.n383 B.n382 585
R513 B.n381 B.n380 585
R514 B.n379 B.n378 585
R515 B.n377 B.n376 585
R516 B.n375 B.n374 585
R517 B.n373 B.n372 585
R518 B.n371 B.n370 585
R519 B.n369 B.n368 585
R520 B.n367 B.n366 585
R521 B.n365 B.n364 585
R522 B.n362 B.n361 585
R523 B.n360 B.n359 585
R524 B.n358 B.n357 585
R525 B.n356 B.n355 585
R526 B.n354 B.n353 585
R527 B.n352 B.n351 585
R528 B.n350 B.n349 585
R529 B.n348 B.n347 585
R530 B.n346 B.n345 585
R531 B.n344 B.n343 585
R532 B.n342 B.n341 585
R533 B.n340 B.n339 585
R534 B.n338 B.n337 585
R535 B.n336 B.n335 585
R536 B.n334 B.n333 585
R537 B.n332 B.n331 585
R538 B.n330 B.n329 585
R539 B.n328 B.n327 585
R540 B.n326 B.n325 585
R541 B.n324 B.n323 585
R542 B.n322 B.n321 585
R543 B.n320 B.n319 585
R544 B.n318 B.n317 585
R545 B.n316 B.n315 585
R546 B.n314 B.n313 585
R547 B.n312 B.n311 585
R548 B.n310 B.n309 585
R549 B.n308 B.n307 585
R550 B.n306 B.n305 585
R551 B.n403 B.n273 585
R552 B.n273 B.n272 585
R553 B.n405 B.n404 585
R554 B.n406 B.n405 585
R555 B.n267 B.n266 585
R556 B.n268 B.n267 585
R557 B.n414 B.n413 585
R558 B.n413 B.n412 585
R559 B.n415 B.n265 585
R560 B.n265 B.n264 585
R561 B.n417 B.n416 585
R562 B.n418 B.n417 585
R563 B.n259 B.n258 585
R564 B.n260 B.n259 585
R565 B.n426 B.n425 585
R566 B.n425 B.n424 585
R567 B.n427 B.n257 585
R568 B.n257 B.n256 585
R569 B.n429 B.n428 585
R570 B.n430 B.n429 585
R571 B.n251 B.n250 585
R572 B.n252 B.n251 585
R573 B.n438 B.n437 585
R574 B.n437 B.n436 585
R575 B.n439 B.n249 585
R576 B.n249 B.n248 585
R577 B.n441 B.n440 585
R578 B.n442 B.n441 585
R579 B.n243 B.n242 585
R580 B.n244 B.n243 585
R581 B.n450 B.n449 585
R582 B.n449 B.n448 585
R583 B.n451 B.n241 585
R584 B.n241 B.n239 585
R585 B.n453 B.n452 585
R586 B.n454 B.n453 585
R587 B.n235 B.n234 585
R588 B.n240 B.n235 585
R589 B.n462 B.n461 585
R590 B.n461 B.n460 585
R591 B.n463 B.n233 585
R592 B.n233 B.n232 585
R593 B.n465 B.n464 585
R594 B.n466 B.n465 585
R595 B.n227 B.n226 585
R596 B.n228 B.n227 585
R597 B.n474 B.n473 585
R598 B.n473 B.n472 585
R599 B.n475 B.n225 585
R600 B.n225 B.n223 585
R601 B.n477 B.n476 585
R602 B.n478 B.n477 585
R603 B.n219 B.n218 585
R604 B.n224 B.n219 585
R605 B.n486 B.n485 585
R606 B.n485 B.n484 585
R607 B.n487 B.n217 585
R608 B.n217 B.n216 585
R609 B.n489 B.n488 585
R610 B.n490 B.n489 585
R611 B.n211 B.n210 585
R612 B.n212 B.n211 585
R613 B.n498 B.n497 585
R614 B.n497 B.n496 585
R615 B.n499 B.n209 585
R616 B.n209 B.n208 585
R617 B.n501 B.n500 585
R618 B.n502 B.n501 585
R619 B.n203 B.n202 585
R620 B.n204 B.n203 585
R621 B.n511 B.n510 585
R622 B.n510 B.n509 585
R623 B.n512 B.n201 585
R624 B.n201 B.n200 585
R625 B.n514 B.n513 585
R626 B.n515 B.n514 585
R627 B.n3 B.n0 585
R628 B.n4 B.n3 585
R629 B.n651 B.n1 585
R630 B.n652 B.n651 585
R631 B.n650 B.n649 585
R632 B.n650 B.n8 585
R633 B.n648 B.n9 585
R634 B.n12 B.n9 585
R635 B.n647 B.n646 585
R636 B.n646 B.n645 585
R637 B.n11 B.n10 585
R638 B.n644 B.n11 585
R639 B.n642 B.n641 585
R640 B.n643 B.n642 585
R641 B.n640 B.n17 585
R642 B.n17 B.n16 585
R643 B.n639 B.n638 585
R644 B.n638 B.n637 585
R645 B.n19 B.n18 585
R646 B.n636 B.n19 585
R647 B.n634 B.n633 585
R648 B.n635 B.n634 585
R649 B.n632 B.n24 585
R650 B.n24 B.n23 585
R651 B.n631 B.n630 585
R652 B.n630 B.n629 585
R653 B.n26 B.n25 585
R654 B.n628 B.n26 585
R655 B.n626 B.n625 585
R656 B.n627 B.n626 585
R657 B.n624 B.n31 585
R658 B.n31 B.n30 585
R659 B.n623 B.n622 585
R660 B.n622 B.n621 585
R661 B.n33 B.n32 585
R662 B.n620 B.n33 585
R663 B.n618 B.n617 585
R664 B.n619 B.n618 585
R665 B.n616 B.n38 585
R666 B.n38 B.n37 585
R667 B.n615 B.n614 585
R668 B.n614 B.n613 585
R669 B.n40 B.n39 585
R670 B.n612 B.n40 585
R671 B.n610 B.n609 585
R672 B.n611 B.n610 585
R673 B.n608 B.n45 585
R674 B.n45 B.n44 585
R675 B.n607 B.n606 585
R676 B.n606 B.n605 585
R677 B.n47 B.n46 585
R678 B.n604 B.n47 585
R679 B.n602 B.n601 585
R680 B.n603 B.n602 585
R681 B.n600 B.n52 585
R682 B.n52 B.n51 585
R683 B.n599 B.n598 585
R684 B.n598 B.n597 585
R685 B.n54 B.n53 585
R686 B.n596 B.n54 585
R687 B.n594 B.n593 585
R688 B.n595 B.n594 585
R689 B.n592 B.n59 585
R690 B.n59 B.n58 585
R691 B.n591 B.n590 585
R692 B.n590 B.n589 585
R693 B.n61 B.n60 585
R694 B.n588 B.n61 585
R695 B.n586 B.n585 585
R696 B.n587 B.n586 585
R697 B.n584 B.n66 585
R698 B.n66 B.n65 585
R699 B.n583 B.n582 585
R700 B.n582 B.n581 585
R701 B.n68 B.n67 585
R702 B.n580 B.n68 585
R703 B.n578 B.n577 585
R704 B.n579 B.n578 585
R705 B.n576 B.n73 585
R706 B.n73 B.n72 585
R707 B.n655 B.n654 585
R708 B.n653 B.n2 585
R709 B.n574 B.n73 478.086
R710 B.n571 B.n100 478.086
R711 B.n305 B.n271 478.086
R712 B.n401 B.n273 478.086
R713 B.n572 B.n98 256.663
R714 B.n572 B.n97 256.663
R715 B.n572 B.n96 256.663
R716 B.n572 B.n95 256.663
R717 B.n572 B.n94 256.663
R718 B.n572 B.n93 256.663
R719 B.n572 B.n92 256.663
R720 B.n572 B.n91 256.663
R721 B.n572 B.n90 256.663
R722 B.n572 B.n89 256.663
R723 B.n572 B.n88 256.663
R724 B.n572 B.n87 256.663
R725 B.n572 B.n86 256.663
R726 B.n572 B.n85 256.663
R727 B.n572 B.n84 256.663
R728 B.n572 B.n83 256.663
R729 B.n572 B.n82 256.663
R730 B.n572 B.n81 256.663
R731 B.n572 B.n80 256.663
R732 B.n572 B.n79 256.663
R733 B.n572 B.n78 256.663
R734 B.n572 B.n77 256.663
R735 B.n572 B.n76 256.663
R736 B.n573 B.n572 256.663
R737 B.n400 B.n399 256.663
R738 B.n399 B.n276 256.663
R739 B.n399 B.n277 256.663
R740 B.n399 B.n278 256.663
R741 B.n399 B.n279 256.663
R742 B.n399 B.n280 256.663
R743 B.n399 B.n281 256.663
R744 B.n399 B.n282 256.663
R745 B.n399 B.n283 256.663
R746 B.n399 B.n284 256.663
R747 B.n399 B.n285 256.663
R748 B.n399 B.n286 256.663
R749 B.n399 B.n287 256.663
R750 B.n399 B.n288 256.663
R751 B.n399 B.n289 256.663
R752 B.n399 B.n290 256.663
R753 B.n399 B.n291 256.663
R754 B.n399 B.n292 256.663
R755 B.n399 B.n293 256.663
R756 B.n399 B.n294 256.663
R757 B.n399 B.n295 256.663
R758 B.n399 B.n296 256.663
R759 B.n399 B.n297 256.663
R760 B.n399 B.n298 256.663
R761 B.n657 B.n656 256.663
R762 B.n103 B.t14 253.964
R763 B.n101 B.t10 253.964
R764 B.n302 B.t17 253.964
R765 B.n300 B.t6 253.964
R766 B.n101 B.t12 204.873
R767 B.n302 B.t19 204.873
R768 B.n103 B.t15 204.873
R769 B.n300 B.t9 204.873
R770 B.n106 B.n75 163.367
R771 B.n110 B.n109 163.367
R772 B.n114 B.n113 163.367
R773 B.n118 B.n117 163.367
R774 B.n122 B.n121 163.367
R775 B.n126 B.n125 163.367
R776 B.n130 B.n129 163.367
R777 B.n134 B.n133 163.367
R778 B.n138 B.n137 163.367
R779 B.n142 B.n141 163.367
R780 B.n146 B.n145 163.367
R781 B.n150 B.n149 163.367
R782 B.n154 B.n153 163.367
R783 B.n158 B.n157 163.367
R784 B.n163 B.n162 163.367
R785 B.n167 B.n166 163.367
R786 B.n171 B.n170 163.367
R787 B.n175 B.n174 163.367
R788 B.n179 B.n178 163.367
R789 B.n183 B.n182 163.367
R790 B.n187 B.n186 163.367
R791 B.n191 B.n190 163.367
R792 B.n195 B.n194 163.367
R793 B.n571 B.n99 163.367
R794 B.n407 B.n271 163.367
R795 B.n407 B.n269 163.367
R796 B.n411 B.n269 163.367
R797 B.n411 B.n263 163.367
R798 B.n419 B.n263 163.367
R799 B.n419 B.n261 163.367
R800 B.n423 B.n261 163.367
R801 B.n423 B.n255 163.367
R802 B.n431 B.n255 163.367
R803 B.n431 B.n253 163.367
R804 B.n435 B.n253 163.367
R805 B.n435 B.n247 163.367
R806 B.n443 B.n247 163.367
R807 B.n443 B.n245 163.367
R808 B.n447 B.n245 163.367
R809 B.n447 B.n238 163.367
R810 B.n455 B.n238 163.367
R811 B.n455 B.n236 163.367
R812 B.n459 B.n236 163.367
R813 B.n459 B.n231 163.367
R814 B.n467 B.n231 163.367
R815 B.n467 B.n229 163.367
R816 B.n471 B.n229 163.367
R817 B.n471 B.n222 163.367
R818 B.n479 B.n222 163.367
R819 B.n479 B.n220 163.367
R820 B.n483 B.n220 163.367
R821 B.n483 B.n215 163.367
R822 B.n491 B.n215 163.367
R823 B.n491 B.n213 163.367
R824 B.n495 B.n213 163.367
R825 B.n495 B.n207 163.367
R826 B.n503 B.n207 163.367
R827 B.n503 B.n205 163.367
R828 B.n508 B.n205 163.367
R829 B.n508 B.n199 163.367
R830 B.n516 B.n199 163.367
R831 B.n517 B.n516 163.367
R832 B.n517 B.n5 163.367
R833 B.n6 B.n5 163.367
R834 B.n7 B.n6 163.367
R835 B.n523 B.n7 163.367
R836 B.n524 B.n523 163.367
R837 B.n524 B.n13 163.367
R838 B.n14 B.n13 163.367
R839 B.n15 B.n14 163.367
R840 B.n529 B.n15 163.367
R841 B.n529 B.n20 163.367
R842 B.n21 B.n20 163.367
R843 B.n22 B.n21 163.367
R844 B.n534 B.n22 163.367
R845 B.n534 B.n27 163.367
R846 B.n28 B.n27 163.367
R847 B.n29 B.n28 163.367
R848 B.n539 B.n29 163.367
R849 B.n539 B.n34 163.367
R850 B.n35 B.n34 163.367
R851 B.n36 B.n35 163.367
R852 B.n544 B.n36 163.367
R853 B.n544 B.n41 163.367
R854 B.n42 B.n41 163.367
R855 B.n43 B.n42 163.367
R856 B.n549 B.n43 163.367
R857 B.n549 B.n48 163.367
R858 B.n49 B.n48 163.367
R859 B.n50 B.n49 163.367
R860 B.n554 B.n50 163.367
R861 B.n554 B.n55 163.367
R862 B.n56 B.n55 163.367
R863 B.n57 B.n56 163.367
R864 B.n559 B.n57 163.367
R865 B.n559 B.n62 163.367
R866 B.n63 B.n62 163.367
R867 B.n64 B.n63 163.367
R868 B.n564 B.n64 163.367
R869 B.n564 B.n69 163.367
R870 B.n70 B.n69 163.367
R871 B.n71 B.n70 163.367
R872 B.n100 B.n71 163.367
R873 B.n398 B.n275 163.367
R874 B.n398 B.n299 163.367
R875 B.n394 B.n393 163.367
R876 B.n390 B.n389 163.367
R877 B.n386 B.n385 163.367
R878 B.n382 B.n381 163.367
R879 B.n378 B.n377 163.367
R880 B.n374 B.n373 163.367
R881 B.n370 B.n369 163.367
R882 B.n366 B.n365 163.367
R883 B.n361 B.n360 163.367
R884 B.n357 B.n356 163.367
R885 B.n353 B.n352 163.367
R886 B.n349 B.n348 163.367
R887 B.n345 B.n344 163.367
R888 B.n341 B.n340 163.367
R889 B.n337 B.n336 163.367
R890 B.n333 B.n332 163.367
R891 B.n329 B.n328 163.367
R892 B.n325 B.n324 163.367
R893 B.n321 B.n320 163.367
R894 B.n317 B.n316 163.367
R895 B.n313 B.n312 163.367
R896 B.n309 B.n308 163.367
R897 B.n405 B.n273 163.367
R898 B.n405 B.n267 163.367
R899 B.n413 B.n267 163.367
R900 B.n413 B.n265 163.367
R901 B.n417 B.n265 163.367
R902 B.n417 B.n259 163.367
R903 B.n425 B.n259 163.367
R904 B.n425 B.n257 163.367
R905 B.n429 B.n257 163.367
R906 B.n429 B.n251 163.367
R907 B.n437 B.n251 163.367
R908 B.n437 B.n249 163.367
R909 B.n441 B.n249 163.367
R910 B.n441 B.n243 163.367
R911 B.n449 B.n243 163.367
R912 B.n449 B.n241 163.367
R913 B.n453 B.n241 163.367
R914 B.n453 B.n235 163.367
R915 B.n461 B.n235 163.367
R916 B.n461 B.n233 163.367
R917 B.n465 B.n233 163.367
R918 B.n465 B.n227 163.367
R919 B.n473 B.n227 163.367
R920 B.n473 B.n225 163.367
R921 B.n477 B.n225 163.367
R922 B.n477 B.n219 163.367
R923 B.n485 B.n219 163.367
R924 B.n485 B.n217 163.367
R925 B.n489 B.n217 163.367
R926 B.n489 B.n211 163.367
R927 B.n497 B.n211 163.367
R928 B.n497 B.n209 163.367
R929 B.n501 B.n209 163.367
R930 B.n501 B.n203 163.367
R931 B.n510 B.n203 163.367
R932 B.n510 B.n201 163.367
R933 B.n514 B.n201 163.367
R934 B.n514 B.n3 163.367
R935 B.n655 B.n3 163.367
R936 B.n651 B.n2 163.367
R937 B.n651 B.n650 163.367
R938 B.n650 B.n9 163.367
R939 B.n646 B.n9 163.367
R940 B.n646 B.n11 163.367
R941 B.n642 B.n11 163.367
R942 B.n642 B.n17 163.367
R943 B.n638 B.n17 163.367
R944 B.n638 B.n19 163.367
R945 B.n634 B.n19 163.367
R946 B.n634 B.n24 163.367
R947 B.n630 B.n24 163.367
R948 B.n630 B.n26 163.367
R949 B.n626 B.n26 163.367
R950 B.n626 B.n31 163.367
R951 B.n622 B.n31 163.367
R952 B.n622 B.n33 163.367
R953 B.n618 B.n33 163.367
R954 B.n618 B.n38 163.367
R955 B.n614 B.n38 163.367
R956 B.n614 B.n40 163.367
R957 B.n610 B.n40 163.367
R958 B.n610 B.n45 163.367
R959 B.n606 B.n45 163.367
R960 B.n606 B.n47 163.367
R961 B.n602 B.n47 163.367
R962 B.n602 B.n52 163.367
R963 B.n598 B.n52 163.367
R964 B.n598 B.n54 163.367
R965 B.n594 B.n54 163.367
R966 B.n594 B.n59 163.367
R967 B.n590 B.n59 163.367
R968 B.n590 B.n61 163.367
R969 B.n586 B.n61 163.367
R970 B.n586 B.n66 163.367
R971 B.n582 B.n66 163.367
R972 B.n582 B.n68 163.367
R973 B.n578 B.n68 163.367
R974 B.n578 B.n73 163.367
R975 B.n102 B.t13 153.091
R976 B.n303 B.t18 153.091
R977 B.n104 B.t16 153.091
R978 B.n301 B.t8 153.091
R979 B.n399 B.n272 140.666
R980 B.n572 B.n72 140.666
R981 B.n406 B.n272 76.5222
R982 B.n406 B.n268 76.5222
R983 B.n412 B.n268 76.5222
R984 B.n412 B.n264 76.5222
R985 B.n418 B.n264 76.5222
R986 B.n418 B.n260 76.5222
R987 B.n424 B.n260 76.5222
R988 B.n430 B.n256 76.5222
R989 B.n430 B.n252 76.5222
R990 B.n436 B.n252 76.5222
R991 B.n436 B.n248 76.5222
R992 B.n442 B.n248 76.5222
R993 B.n442 B.n244 76.5222
R994 B.n448 B.n244 76.5222
R995 B.n448 B.n239 76.5222
R996 B.n454 B.n239 76.5222
R997 B.n454 B.n240 76.5222
R998 B.n460 B.n232 76.5222
R999 B.n466 B.n232 76.5222
R1000 B.n466 B.n228 76.5222
R1001 B.n472 B.n228 76.5222
R1002 B.n472 B.n223 76.5222
R1003 B.n478 B.n223 76.5222
R1004 B.n478 B.n224 76.5222
R1005 B.n484 B.n216 76.5222
R1006 B.n490 B.n216 76.5222
R1007 B.n490 B.n212 76.5222
R1008 B.n496 B.n212 76.5222
R1009 B.n496 B.n208 76.5222
R1010 B.n502 B.n208 76.5222
R1011 B.n509 B.n204 76.5222
R1012 B.n509 B.n200 76.5222
R1013 B.n515 B.n200 76.5222
R1014 B.n515 B.n4 76.5222
R1015 B.n654 B.n4 76.5222
R1016 B.n654 B.n653 76.5222
R1017 B.n653 B.n652 76.5222
R1018 B.n652 B.n8 76.5222
R1019 B.n12 B.n8 76.5222
R1020 B.n645 B.n12 76.5222
R1021 B.n645 B.n644 76.5222
R1022 B.n643 B.n16 76.5222
R1023 B.n637 B.n16 76.5222
R1024 B.n637 B.n636 76.5222
R1025 B.n636 B.n635 76.5222
R1026 B.n635 B.n23 76.5222
R1027 B.n629 B.n23 76.5222
R1028 B.n628 B.n627 76.5222
R1029 B.n627 B.n30 76.5222
R1030 B.n621 B.n30 76.5222
R1031 B.n621 B.n620 76.5222
R1032 B.n620 B.n619 76.5222
R1033 B.n619 B.n37 76.5222
R1034 B.n613 B.n37 76.5222
R1035 B.n612 B.n611 76.5222
R1036 B.n611 B.n44 76.5222
R1037 B.n605 B.n44 76.5222
R1038 B.n605 B.n604 76.5222
R1039 B.n604 B.n603 76.5222
R1040 B.n603 B.n51 76.5222
R1041 B.n597 B.n51 76.5222
R1042 B.n597 B.n596 76.5222
R1043 B.n596 B.n595 76.5222
R1044 B.n595 B.n58 76.5222
R1045 B.n589 B.n588 76.5222
R1046 B.n588 B.n587 76.5222
R1047 B.n587 B.n65 76.5222
R1048 B.n581 B.n65 76.5222
R1049 B.n581 B.n580 76.5222
R1050 B.n580 B.n579 76.5222
R1051 B.n579 B.n72 76.5222
R1052 B.n502 B.t0 74.2716
R1053 B.t1 B.n643 74.2716
R1054 B.n574 B.n573 71.676
R1055 B.n106 B.n76 71.676
R1056 B.n110 B.n77 71.676
R1057 B.n114 B.n78 71.676
R1058 B.n118 B.n79 71.676
R1059 B.n122 B.n80 71.676
R1060 B.n126 B.n81 71.676
R1061 B.n130 B.n82 71.676
R1062 B.n134 B.n83 71.676
R1063 B.n138 B.n84 71.676
R1064 B.n142 B.n85 71.676
R1065 B.n146 B.n86 71.676
R1066 B.n150 B.n87 71.676
R1067 B.n154 B.n88 71.676
R1068 B.n158 B.n89 71.676
R1069 B.n163 B.n90 71.676
R1070 B.n167 B.n91 71.676
R1071 B.n171 B.n92 71.676
R1072 B.n175 B.n93 71.676
R1073 B.n179 B.n94 71.676
R1074 B.n183 B.n95 71.676
R1075 B.n187 B.n96 71.676
R1076 B.n191 B.n97 71.676
R1077 B.n195 B.n98 71.676
R1078 B.n99 B.n98 71.676
R1079 B.n194 B.n97 71.676
R1080 B.n190 B.n96 71.676
R1081 B.n186 B.n95 71.676
R1082 B.n182 B.n94 71.676
R1083 B.n178 B.n93 71.676
R1084 B.n174 B.n92 71.676
R1085 B.n170 B.n91 71.676
R1086 B.n166 B.n90 71.676
R1087 B.n162 B.n89 71.676
R1088 B.n157 B.n88 71.676
R1089 B.n153 B.n87 71.676
R1090 B.n149 B.n86 71.676
R1091 B.n145 B.n85 71.676
R1092 B.n141 B.n84 71.676
R1093 B.n137 B.n83 71.676
R1094 B.n133 B.n82 71.676
R1095 B.n129 B.n81 71.676
R1096 B.n125 B.n80 71.676
R1097 B.n121 B.n79 71.676
R1098 B.n117 B.n78 71.676
R1099 B.n113 B.n77 71.676
R1100 B.n109 B.n76 71.676
R1101 B.n573 B.n75 71.676
R1102 B.n401 B.n400 71.676
R1103 B.n299 B.n276 71.676
R1104 B.n393 B.n277 71.676
R1105 B.n389 B.n278 71.676
R1106 B.n385 B.n279 71.676
R1107 B.n381 B.n280 71.676
R1108 B.n377 B.n281 71.676
R1109 B.n373 B.n282 71.676
R1110 B.n369 B.n283 71.676
R1111 B.n365 B.n284 71.676
R1112 B.n360 B.n285 71.676
R1113 B.n356 B.n286 71.676
R1114 B.n352 B.n287 71.676
R1115 B.n348 B.n288 71.676
R1116 B.n344 B.n289 71.676
R1117 B.n340 B.n290 71.676
R1118 B.n336 B.n291 71.676
R1119 B.n332 B.n292 71.676
R1120 B.n328 B.n293 71.676
R1121 B.n324 B.n294 71.676
R1122 B.n320 B.n295 71.676
R1123 B.n316 B.n296 71.676
R1124 B.n312 B.n297 71.676
R1125 B.n308 B.n298 71.676
R1126 B.n400 B.n275 71.676
R1127 B.n394 B.n276 71.676
R1128 B.n390 B.n277 71.676
R1129 B.n386 B.n278 71.676
R1130 B.n382 B.n279 71.676
R1131 B.n378 B.n280 71.676
R1132 B.n374 B.n281 71.676
R1133 B.n370 B.n282 71.676
R1134 B.n366 B.n283 71.676
R1135 B.n361 B.n284 71.676
R1136 B.n357 B.n285 71.676
R1137 B.n353 B.n286 71.676
R1138 B.n349 B.n287 71.676
R1139 B.n345 B.n288 71.676
R1140 B.n341 B.n289 71.676
R1141 B.n337 B.n290 71.676
R1142 B.n333 B.n291 71.676
R1143 B.n329 B.n292 71.676
R1144 B.n325 B.n293 71.676
R1145 B.n321 B.n294 71.676
R1146 B.n317 B.n295 71.676
R1147 B.n313 B.n296 71.676
R1148 B.n309 B.n297 71.676
R1149 B.n305 B.n298 71.676
R1150 B.n656 B.n655 71.676
R1151 B.n656 B.n2 71.676
R1152 B.n484 B.t2 67.5197
R1153 B.n629 B.t3 67.5197
R1154 B.t7 B.n256 60.7678
R1155 B.t11 B.n58 60.7678
R1156 B.n105 B.n104 59.5399
R1157 B.n160 B.n102 59.5399
R1158 B.n304 B.n303 59.5399
R1159 B.n363 B.n301 59.5399
R1160 B.n460 B.t4 56.2665
R1161 B.n613 B.t5 56.2665
R1162 B.n104 B.n103 51.7823
R1163 B.n102 B.n101 51.7823
R1164 B.n303 B.n302 51.7823
R1165 B.n301 B.n300 51.7823
R1166 B.n403 B.n402 31.0639
R1167 B.n306 B.n270 31.0639
R1168 B.n570 B.n569 31.0639
R1169 B.n576 B.n575 31.0639
R1170 B.n240 B.t4 20.2563
R1171 B.t5 B.n612 20.2563
R1172 B B.n657 18.0485
R1173 B.n424 B.t7 15.755
R1174 B.n589 B.t11 15.755
R1175 B.n404 B.n403 10.6151
R1176 B.n404 B.n266 10.6151
R1177 B.n414 B.n266 10.6151
R1178 B.n415 B.n414 10.6151
R1179 B.n416 B.n415 10.6151
R1180 B.n416 B.n258 10.6151
R1181 B.n426 B.n258 10.6151
R1182 B.n427 B.n426 10.6151
R1183 B.n428 B.n427 10.6151
R1184 B.n428 B.n250 10.6151
R1185 B.n438 B.n250 10.6151
R1186 B.n439 B.n438 10.6151
R1187 B.n440 B.n439 10.6151
R1188 B.n440 B.n242 10.6151
R1189 B.n450 B.n242 10.6151
R1190 B.n451 B.n450 10.6151
R1191 B.n452 B.n451 10.6151
R1192 B.n452 B.n234 10.6151
R1193 B.n462 B.n234 10.6151
R1194 B.n463 B.n462 10.6151
R1195 B.n464 B.n463 10.6151
R1196 B.n464 B.n226 10.6151
R1197 B.n474 B.n226 10.6151
R1198 B.n475 B.n474 10.6151
R1199 B.n476 B.n475 10.6151
R1200 B.n476 B.n218 10.6151
R1201 B.n486 B.n218 10.6151
R1202 B.n487 B.n486 10.6151
R1203 B.n488 B.n487 10.6151
R1204 B.n488 B.n210 10.6151
R1205 B.n498 B.n210 10.6151
R1206 B.n499 B.n498 10.6151
R1207 B.n500 B.n499 10.6151
R1208 B.n500 B.n202 10.6151
R1209 B.n511 B.n202 10.6151
R1210 B.n512 B.n511 10.6151
R1211 B.n513 B.n512 10.6151
R1212 B.n513 B.n0 10.6151
R1213 B.n402 B.n274 10.6151
R1214 B.n397 B.n274 10.6151
R1215 B.n397 B.n396 10.6151
R1216 B.n396 B.n395 10.6151
R1217 B.n395 B.n392 10.6151
R1218 B.n392 B.n391 10.6151
R1219 B.n391 B.n388 10.6151
R1220 B.n388 B.n387 10.6151
R1221 B.n387 B.n384 10.6151
R1222 B.n384 B.n383 10.6151
R1223 B.n383 B.n380 10.6151
R1224 B.n380 B.n379 10.6151
R1225 B.n379 B.n376 10.6151
R1226 B.n376 B.n375 10.6151
R1227 B.n375 B.n372 10.6151
R1228 B.n372 B.n371 10.6151
R1229 B.n371 B.n368 10.6151
R1230 B.n368 B.n367 10.6151
R1231 B.n367 B.n364 10.6151
R1232 B.n362 B.n359 10.6151
R1233 B.n359 B.n358 10.6151
R1234 B.n358 B.n355 10.6151
R1235 B.n355 B.n354 10.6151
R1236 B.n354 B.n351 10.6151
R1237 B.n351 B.n350 10.6151
R1238 B.n350 B.n347 10.6151
R1239 B.n347 B.n346 10.6151
R1240 B.n343 B.n342 10.6151
R1241 B.n342 B.n339 10.6151
R1242 B.n339 B.n338 10.6151
R1243 B.n338 B.n335 10.6151
R1244 B.n335 B.n334 10.6151
R1245 B.n334 B.n331 10.6151
R1246 B.n331 B.n330 10.6151
R1247 B.n330 B.n327 10.6151
R1248 B.n327 B.n326 10.6151
R1249 B.n326 B.n323 10.6151
R1250 B.n323 B.n322 10.6151
R1251 B.n322 B.n319 10.6151
R1252 B.n319 B.n318 10.6151
R1253 B.n318 B.n315 10.6151
R1254 B.n315 B.n314 10.6151
R1255 B.n314 B.n311 10.6151
R1256 B.n311 B.n310 10.6151
R1257 B.n310 B.n307 10.6151
R1258 B.n307 B.n306 10.6151
R1259 B.n408 B.n270 10.6151
R1260 B.n409 B.n408 10.6151
R1261 B.n410 B.n409 10.6151
R1262 B.n410 B.n262 10.6151
R1263 B.n420 B.n262 10.6151
R1264 B.n421 B.n420 10.6151
R1265 B.n422 B.n421 10.6151
R1266 B.n422 B.n254 10.6151
R1267 B.n432 B.n254 10.6151
R1268 B.n433 B.n432 10.6151
R1269 B.n434 B.n433 10.6151
R1270 B.n434 B.n246 10.6151
R1271 B.n444 B.n246 10.6151
R1272 B.n445 B.n444 10.6151
R1273 B.n446 B.n445 10.6151
R1274 B.n446 B.n237 10.6151
R1275 B.n456 B.n237 10.6151
R1276 B.n457 B.n456 10.6151
R1277 B.n458 B.n457 10.6151
R1278 B.n458 B.n230 10.6151
R1279 B.n468 B.n230 10.6151
R1280 B.n469 B.n468 10.6151
R1281 B.n470 B.n469 10.6151
R1282 B.n470 B.n221 10.6151
R1283 B.n480 B.n221 10.6151
R1284 B.n481 B.n480 10.6151
R1285 B.n482 B.n481 10.6151
R1286 B.n482 B.n214 10.6151
R1287 B.n492 B.n214 10.6151
R1288 B.n493 B.n492 10.6151
R1289 B.n494 B.n493 10.6151
R1290 B.n494 B.n206 10.6151
R1291 B.n504 B.n206 10.6151
R1292 B.n505 B.n504 10.6151
R1293 B.n507 B.n505 10.6151
R1294 B.n507 B.n506 10.6151
R1295 B.n506 B.n198 10.6151
R1296 B.n518 B.n198 10.6151
R1297 B.n519 B.n518 10.6151
R1298 B.n520 B.n519 10.6151
R1299 B.n521 B.n520 10.6151
R1300 B.n522 B.n521 10.6151
R1301 B.n525 B.n522 10.6151
R1302 B.n526 B.n525 10.6151
R1303 B.n527 B.n526 10.6151
R1304 B.n528 B.n527 10.6151
R1305 B.n530 B.n528 10.6151
R1306 B.n531 B.n530 10.6151
R1307 B.n532 B.n531 10.6151
R1308 B.n533 B.n532 10.6151
R1309 B.n535 B.n533 10.6151
R1310 B.n536 B.n535 10.6151
R1311 B.n537 B.n536 10.6151
R1312 B.n538 B.n537 10.6151
R1313 B.n540 B.n538 10.6151
R1314 B.n541 B.n540 10.6151
R1315 B.n542 B.n541 10.6151
R1316 B.n543 B.n542 10.6151
R1317 B.n545 B.n543 10.6151
R1318 B.n546 B.n545 10.6151
R1319 B.n547 B.n546 10.6151
R1320 B.n548 B.n547 10.6151
R1321 B.n550 B.n548 10.6151
R1322 B.n551 B.n550 10.6151
R1323 B.n552 B.n551 10.6151
R1324 B.n553 B.n552 10.6151
R1325 B.n555 B.n553 10.6151
R1326 B.n556 B.n555 10.6151
R1327 B.n557 B.n556 10.6151
R1328 B.n558 B.n557 10.6151
R1329 B.n560 B.n558 10.6151
R1330 B.n561 B.n560 10.6151
R1331 B.n562 B.n561 10.6151
R1332 B.n563 B.n562 10.6151
R1333 B.n565 B.n563 10.6151
R1334 B.n566 B.n565 10.6151
R1335 B.n567 B.n566 10.6151
R1336 B.n568 B.n567 10.6151
R1337 B.n569 B.n568 10.6151
R1338 B.n649 B.n1 10.6151
R1339 B.n649 B.n648 10.6151
R1340 B.n648 B.n647 10.6151
R1341 B.n647 B.n10 10.6151
R1342 B.n641 B.n10 10.6151
R1343 B.n641 B.n640 10.6151
R1344 B.n640 B.n639 10.6151
R1345 B.n639 B.n18 10.6151
R1346 B.n633 B.n18 10.6151
R1347 B.n633 B.n632 10.6151
R1348 B.n632 B.n631 10.6151
R1349 B.n631 B.n25 10.6151
R1350 B.n625 B.n25 10.6151
R1351 B.n625 B.n624 10.6151
R1352 B.n624 B.n623 10.6151
R1353 B.n623 B.n32 10.6151
R1354 B.n617 B.n32 10.6151
R1355 B.n617 B.n616 10.6151
R1356 B.n616 B.n615 10.6151
R1357 B.n615 B.n39 10.6151
R1358 B.n609 B.n39 10.6151
R1359 B.n609 B.n608 10.6151
R1360 B.n608 B.n607 10.6151
R1361 B.n607 B.n46 10.6151
R1362 B.n601 B.n46 10.6151
R1363 B.n601 B.n600 10.6151
R1364 B.n600 B.n599 10.6151
R1365 B.n599 B.n53 10.6151
R1366 B.n593 B.n53 10.6151
R1367 B.n593 B.n592 10.6151
R1368 B.n592 B.n591 10.6151
R1369 B.n591 B.n60 10.6151
R1370 B.n585 B.n60 10.6151
R1371 B.n585 B.n584 10.6151
R1372 B.n584 B.n583 10.6151
R1373 B.n583 B.n67 10.6151
R1374 B.n577 B.n67 10.6151
R1375 B.n577 B.n576 10.6151
R1376 B.n575 B.n74 10.6151
R1377 B.n107 B.n74 10.6151
R1378 B.n108 B.n107 10.6151
R1379 B.n111 B.n108 10.6151
R1380 B.n112 B.n111 10.6151
R1381 B.n115 B.n112 10.6151
R1382 B.n116 B.n115 10.6151
R1383 B.n119 B.n116 10.6151
R1384 B.n120 B.n119 10.6151
R1385 B.n123 B.n120 10.6151
R1386 B.n124 B.n123 10.6151
R1387 B.n127 B.n124 10.6151
R1388 B.n128 B.n127 10.6151
R1389 B.n131 B.n128 10.6151
R1390 B.n132 B.n131 10.6151
R1391 B.n135 B.n132 10.6151
R1392 B.n136 B.n135 10.6151
R1393 B.n139 B.n136 10.6151
R1394 B.n140 B.n139 10.6151
R1395 B.n144 B.n143 10.6151
R1396 B.n147 B.n144 10.6151
R1397 B.n148 B.n147 10.6151
R1398 B.n151 B.n148 10.6151
R1399 B.n152 B.n151 10.6151
R1400 B.n155 B.n152 10.6151
R1401 B.n156 B.n155 10.6151
R1402 B.n159 B.n156 10.6151
R1403 B.n164 B.n161 10.6151
R1404 B.n165 B.n164 10.6151
R1405 B.n168 B.n165 10.6151
R1406 B.n169 B.n168 10.6151
R1407 B.n172 B.n169 10.6151
R1408 B.n173 B.n172 10.6151
R1409 B.n176 B.n173 10.6151
R1410 B.n177 B.n176 10.6151
R1411 B.n180 B.n177 10.6151
R1412 B.n181 B.n180 10.6151
R1413 B.n184 B.n181 10.6151
R1414 B.n185 B.n184 10.6151
R1415 B.n188 B.n185 10.6151
R1416 B.n189 B.n188 10.6151
R1417 B.n192 B.n189 10.6151
R1418 B.n193 B.n192 10.6151
R1419 B.n196 B.n193 10.6151
R1420 B.n197 B.n196 10.6151
R1421 B.n570 B.n197 10.6151
R1422 B.n224 B.t2 9.00306
R1423 B.t3 B.n628 9.00306
R1424 B.n657 B.n0 8.11757
R1425 B.n657 B.n1 8.11757
R1426 B.n363 B.n362 6.5566
R1427 B.n346 B.n304 6.5566
R1428 B.n143 B.n105 6.5566
R1429 B.n160 B.n159 6.5566
R1430 B.n364 B.n363 4.05904
R1431 B.n343 B.n304 4.05904
R1432 B.n140 B.n105 4.05904
R1433 B.n161 B.n160 4.05904
R1434 B.t0 B.n204 2.25114
R1435 B.n644 B.t1 2.25114
R1436 VP.n11 VP.n8 161.3
R1437 VP.n13 VP.n12 161.3
R1438 VP.n14 VP.n7 161.3
R1439 VP.n16 VP.n15 161.3
R1440 VP.n17 VP.n6 161.3
R1441 VP.n37 VP.n0 161.3
R1442 VP.n36 VP.n35 161.3
R1443 VP.n34 VP.n1 161.3
R1444 VP.n33 VP.n32 161.3
R1445 VP.n31 VP.n2 161.3
R1446 VP.n30 VP.n29 161.3
R1447 VP.n28 VP.n3 161.3
R1448 VP.n27 VP.n26 161.3
R1449 VP.n25 VP.n4 161.3
R1450 VP.n24 VP.n23 161.3
R1451 VP.n22 VP.n5 161.3
R1452 VP.n21 VP.n20 102.547
R1453 VP.n39 VP.n38 102.547
R1454 VP.n19 VP.n18 102.547
R1455 VP.n9 VP.t3 79.5466
R1456 VP.n26 VP.n25 56.5617
R1457 VP.n32 VP.n1 56.5617
R1458 VP.n12 VP.n7 56.5617
R1459 VP.n10 VP.n9 47.9848
R1460 VP.n30 VP.t0 46.3467
R1461 VP.n20 VP.t4 46.3467
R1462 VP.n38 VP.t2 46.3467
R1463 VP.n10 VP.t5 46.3467
R1464 VP.n18 VP.t1 46.3467
R1465 VP.n21 VP.n19 41.905
R1466 VP.n24 VP.n5 24.5923
R1467 VP.n25 VP.n24 24.5923
R1468 VP.n26 VP.n3 24.5923
R1469 VP.n30 VP.n3 24.5923
R1470 VP.n31 VP.n30 24.5923
R1471 VP.n32 VP.n31 24.5923
R1472 VP.n36 VP.n1 24.5923
R1473 VP.n37 VP.n36 24.5923
R1474 VP.n16 VP.n7 24.5923
R1475 VP.n17 VP.n16 24.5923
R1476 VP.n11 VP.n10 24.5923
R1477 VP.n12 VP.n11 24.5923
R1478 VP.n20 VP.n5 8.36172
R1479 VP.n38 VP.n37 8.36172
R1480 VP.n18 VP.n17 8.36172
R1481 VP.n9 VP.n8 6.93618
R1482 VP.n19 VP.n6 0.278335
R1483 VP.n22 VP.n21 0.278335
R1484 VP.n39 VP.n0 0.278335
R1485 VP.n13 VP.n8 0.189894
R1486 VP.n14 VP.n13 0.189894
R1487 VP.n15 VP.n14 0.189894
R1488 VP.n15 VP.n6 0.189894
R1489 VP.n23 VP.n22 0.189894
R1490 VP.n23 VP.n4 0.189894
R1491 VP.n27 VP.n4 0.189894
R1492 VP.n28 VP.n27 0.189894
R1493 VP.n29 VP.n28 0.189894
R1494 VP.n29 VP.n2 0.189894
R1495 VP.n33 VP.n2 0.189894
R1496 VP.n34 VP.n33 0.189894
R1497 VP.n35 VP.n34 0.189894
R1498 VP.n35 VP.n0 0.189894
R1499 VP VP.n39 0.153485
R1500 VDD1.n18 VDD1.n0 289.615
R1501 VDD1.n41 VDD1.n23 289.615
R1502 VDD1.n19 VDD1.n18 185
R1503 VDD1.n17 VDD1.n16 185
R1504 VDD1.n4 VDD1.n3 185
R1505 VDD1.n11 VDD1.n10 185
R1506 VDD1.n9 VDD1.n8 185
R1507 VDD1.n32 VDD1.n31 185
R1508 VDD1.n34 VDD1.n33 185
R1509 VDD1.n27 VDD1.n26 185
R1510 VDD1.n40 VDD1.n39 185
R1511 VDD1.n42 VDD1.n41 185
R1512 VDD1.n7 VDD1.t2 147.714
R1513 VDD1.n30 VDD1.t1 147.714
R1514 VDD1.n18 VDD1.n17 104.615
R1515 VDD1.n17 VDD1.n3 104.615
R1516 VDD1.n10 VDD1.n3 104.615
R1517 VDD1.n10 VDD1.n9 104.615
R1518 VDD1.n33 VDD1.n32 104.615
R1519 VDD1.n33 VDD1.n26 104.615
R1520 VDD1.n40 VDD1.n26 104.615
R1521 VDD1.n41 VDD1.n40 104.615
R1522 VDD1.n47 VDD1.n46 69.9981
R1523 VDD1.n49 VDD1.n48 69.478
R1524 VDD1.n9 VDD1.t2 52.3082
R1525 VDD1.n32 VDD1.t1 52.3082
R1526 VDD1 VDD1.n22 49.485
R1527 VDD1.n47 VDD1.n45 49.3714
R1528 VDD1.n49 VDD1.n47 36.8091
R1529 VDD1.n8 VDD1.n7 15.6631
R1530 VDD1.n31 VDD1.n30 15.6631
R1531 VDD1.n11 VDD1.n6 12.8005
R1532 VDD1.n34 VDD1.n29 12.8005
R1533 VDD1.n12 VDD1.n4 12.0247
R1534 VDD1.n35 VDD1.n27 12.0247
R1535 VDD1.n16 VDD1.n15 11.249
R1536 VDD1.n39 VDD1.n38 11.249
R1537 VDD1.n19 VDD1.n2 10.4732
R1538 VDD1.n42 VDD1.n25 10.4732
R1539 VDD1.n20 VDD1.n0 9.69747
R1540 VDD1.n43 VDD1.n23 9.69747
R1541 VDD1.n22 VDD1.n21 9.45567
R1542 VDD1.n45 VDD1.n44 9.45567
R1543 VDD1.n21 VDD1.n20 9.3005
R1544 VDD1.n2 VDD1.n1 9.3005
R1545 VDD1.n15 VDD1.n14 9.3005
R1546 VDD1.n13 VDD1.n12 9.3005
R1547 VDD1.n6 VDD1.n5 9.3005
R1548 VDD1.n44 VDD1.n43 9.3005
R1549 VDD1.n25 VDD1.n24 9.3005
R1550 VDD1.n38 VDD1.n37 9.3005
R1551 VDD1.n36 VDD1.n35 9.3005
R1552 VDD1.n29 VDD1.n28 9.3005
R1553 VDD1.n48 VDD1.t0 4.4005
R1554 VDD1.n48 VDD1.t4 4.4005
R1555 VDD1.n46 VDD1.t5 4.4005
R1556 VDD1.n46 VDD1.t3 4.4005
R1557 VDD1.n7 VDD1.n5 4.39059
R1558 VDD1.n30 VDD1.n28 4.39059
R1559 VDD1.n22 VDD1.n0 4.26717
R1560 VDD1.n45 VDD1.n23 4.26717
R1561 VDD1.n20 VDD1.n19 3.49141
R1562 VDD1.n43 VDD1.n42 3.49141
R1563 VDD1.n16 VDD1.n2 2.71565
R1564 VDD1.n39 VDD1.n25 2.71565
R1565 VDD1.n15 VDD1.n4 1.93989
R1566 VDD1.n38 VDD1.n27 1.93989
R1567 VDD1.n12 VDD1.n11 1.16414
R1568 VDD1.n35 VDD1.n34 1.16414
R1569 VDD1 VDD1.n49 0.517741
R1570 VDD1.n8 VDD1.n6 0.388379
R1571 VDD1.n31 VDD1.n29 0.388379
R1572 VDD1.n21 VDD1.n1 0.155672
R1573 VDD1.n14 VDD1.n1 0.155672
R1574 VDD1.n14 VDD1.n13 0.155672
R1575 VDD1.n13 VDD1.n5 0.155672
R1576 VDD1.n36 VDD1.n28 0.155672
R1577 VDD1.n37 VDD1.n36 0.155672
R1578 VDD1.n37 VDD1.n24 0.155672
R1579 VDD1.n44 VDD1.n24 0.155672
C0 VDD1 VTAIL 4.86838f
C1 VDD1 VN 0.1548f
C2 VP VDD1 2.98974f
C3 VDD2 VDD1 1.30527f
C4 VN VTAIL 3.28251f
C5 VP VTAIL 3.2967f
C6 VP VN 5.28978f
C7 VDD2 VTAIL 4.9191f
C8 VDD2 VN 2.7064f
C9 VP VDD2 0.440503f
C10 VDD2 B 4.446501f
C11 VDD1 B 4.566324f
C12 VTAIL B 4.359386f
C13 VN B 11.40347f
C14 VP B 10.035871f
C15 VDD1.n0 B 0.029643f
C16 VDD1.n1 B 0.022609f
C17 VDD1.n2 B 0.012149f
C18 VDD1.n3 B 0.028715f
C19 VDD1.n4 B 0.012864f
C20 VDD1.n5 B 0.381723f
C21 VDD1.n6 B 0.012149f
C22 VDD1.t2 B 0.046984f
C23 VDD1.n7 B 0.088767f
C24 VDD1.n8 B 0.016946f
C25 VDD1.n9 B 0.021537f
C26 VDD1.n10 B 0.028715f
C27 VDD1.n11 B 0.012864f
C28 VDD1.n12 B 0.012149f
C29 VDD1.n13 B 0.022609f
C30 VDD1.n14 B 0.022609f
C31 VDD1.n15 B 0.012149f
C32 VDD1.n16 B 0.012864f
C33 VDD1.n17 B 0.028715f
C34 VDD1.n18 B 0.058388f
C35 VDD1.n19 B 0.012864f
C36 VDD1.n20 B 0.012149f
C37 VDD1.n21 B 0.050405f
C38 VDD1.n22 B 0.05407f
C39 VDD1.n23 B 0.029643f
C40 VDD1.n24 B 0.022609f
C41 VDD1.n25 B 0.012149f
C42 VDD1.n26 B 0.028715f
C43 VDD1.n27 B 0.012864f
C44 VDD1.n28 B 0.381723f
C45 VDD1.n29 B 0.012149f
C46 VDD1.t1 B 0.046984f
C47 VDD1.n30 B 0.088767f
C48 VDD1.n31 B 0.016946f
C49 VDD1.n32 B 0.021537f
C50 VDD1.n33 B 0.028715f
C51 VDD1.n34 B 0.012864f
C52 VDD1.n35 B 0.012149f
C53 VDD1.n36 B 0.022609f
C54 VDD1.n37 B 0.022609f
C55 VDD1.n38 B 0.012149f
C56 VDD1.n39 B 0.012864f
C57 VDD1.n40 B 0.028715f
C58 VDD1.n41 B 0.058388f
C59 VDD1.n42 B 0.012864f
C60 VDD1.n43 B 0.012149f
C61 VDD1.n44 B 0.050405f
C62 VDD1.n45 B 0.053418f
C63 VDD1.t5 B 0.080397f
C64 VDD1.t3 B 0.080397f
C65 VDD1.n46 B 0.647496f
C66 VDD1.n47 B 2.00362f
C67 VDD1.t0 B 0.080397f
C68 VDD1.t4 B 0.080397f
C69 VDD1.n48 B 0.644571f
C70 VDD1.n49 B 1.92018f
C71 VP.n0 B 0.039478f
C72 VP.t2 B 0.818238f
C73 VP.n1 B 0.036488f
C74 VP.n2 B 0.029946f
C75 VP.t0 B 0.818238f
C76 VP.n3 B 0.055531f
C77 VP.n4 B 0.029946f
C78 VP.n5 B 0.037438f
C79 VP.n6 B 0.039478f
C80 VP.t1 B 0.818238f
C81 VP.n7 B 0.036488f
C82 VP.n8 B 0.281352f
C83 VP.t5 B 0.818238f
C84 VP.t3 B 1.02372f
C85 VP.n9 B 0.386449f
C86 VP.n10 B 0.418807f
C87 VP.n11 B 0.055531f
C88 VP.n12 B 0.050573f
C89 VP.n13 B 0.029946f
C90 VP.n14 B 0.029946f
C91 VP.n15 B 0.029946f
C92 VP.n16 B 0.055531f
C93 VP.n17 B 0.037438f
C94 VP.n18 B 0.408643f
C95 VP.n19 B 1.2668f
C96 VP.t4 B 0.818238f
C97 VP.n20 B 0.408643f
C98 VP.n21 B 1.29256f
C99 VP.n22 B 0.039478f
C100 VP.n23 B 0.029946f
C101 VP.n24 B 0.055531f
C102 VP.n25 B 0.036488f
C103 VP.n26 B 0.050573f
C104 VP.n27 B 0.029946f
C105 VP.n28 B 0.029946f
C106 VP.n29 B 0.029946f
C107 VP.n30 B 0.350097f
C108 VP.n31 B 0.055531f
C109 VP.n32 B 0.050573f
C110 VP.n33 B 0.029946f
C111 VP.n34 B 0.029946f
C112 VP.n35 B 0.029946f
C113 VP.n36 B 0.055531f
C114 VP.n37 B 0.037438f
C115 VP.n38 B 0.408643f
C116 VP.n39 B 0.047358f
C117 VTAIL.t6 B 0.101165f
C118 VTAIL.t10 B 0.101165f
C119 VTAIL.n0 B 0.742058f
C120 VTAIL.n1 B 0.460918f
C121 VTAIL.n2 B 0.0373f
C122 VTAIL.n3 B 0.028449f
C123 VTAIL.n4 B 0.015287f
C124 VTAIL.n5 B 0.036133f
C125 VTAIL.n6 B 0.016186f
C126 VTAIL.n7 B 0.480331f
C127 VTAIL.n8 B 0.015287f
C128 VTAIL.t0 B 0.059121f
C129 VTAIL.n9 B 0.111698f
C130 VTAIL.n10 B 0.021324f
C131 VTAIL.n11 B 0.0271f
C132 VTAIL.n12 B 0.036133f
C133 VTAIL.n13 B 0.016186f
C134 VTAIL.n14 B 0.015287f
C135 VTAIL.n15 B 0.028449f
C136 VTAIL.n16 B 0.028449f
C137 VTAIL.n17 B 0.015287f
C138 VTAIL.n18 B 0.016186f
C139 VTAIL.n19 B 0.036133f
C140 VTAIL.n20 B 0.073471f
C141 VTAIL.n21 B 0.016186f
C142 VTAIL.n22 B 0.015287f
C143 VTAIL.n23 B 0.063426f
C144 VTAIL.n24 B 0.040548f
C145 VTAIL.n25 B 0.382546f
C146 VTAIL.t4 B 0.101165f
C147 VTAIL.t2 B 0.101165f
C148 VTAIL.n26 B 0.742058f
C149 VTAIL.n27 B 1.62931f
C150 VTAIL.t8 B 0.101165f
C151 VTAIL.t11 B 0.101165f
C152 VTAIL.n28 B 0.742063f
C153 VTAIL.n29 B 1.62931f
C154 VTAIL.n30 B 0.0373f
C155 VTAIL.n31 B 0.028449f
C156 VTAIL.n32 B 0.015287f
C157 VTAIL.n33 B 0.036133f
C158 VTAIL.n34 B 0.016186f
C159 VTAIL.n35 B 0.480331f
C160 VTAIL.n36 B 0.015287f
C161 VTAIL.t9 B 0.059121f
C162 VTAIL.n37 B 0.111698f
C163 VTAIL.n38 B 0.021324f
C164 VTAIL.n39 B 0.0271f
C165 VTAIL.n40 B 0.036133f
C166 VTAIL.n41 B 0.016186f
C167 VTAIL.n42 B 0.015287f
C168 VTAIL.n43 B 0.028449f
C169 VTAIL.n44 B 0.028449f
C170 VTAIL.n45 B 0.015287f
C171 VTAIL.n46 B 0.016186f
C172 VTAIL.n47 B 0.036133f
C173 VTAIL.n48 B 0.073471f
C174 VTAIL.n49 B 0.016186f
C175 VTAIL.n50 B 0.015287f
C176 VTAIL.n51 B 0.063426f
C177 VTAIL.n52 B 0.040548f
C178 VTAIL.n53 B 0.382546f
C179 VTAIL.t1 B 0.101165f
C180 VTAIL.t3 B 0.101165f
C181 VTAIL.n54 B 0.742063f
C182 VTAIL.n55 B 0.613826f
C183 VTAIL.n56 B 0.0373f
C184 VTAIL.n57 B 0.028449f
C185 VTAIL.n58 B 0.015287f
C186 VTAIL.n59 B 0.036133f
C187 VTAIL.n60 B 0.016186f
C188 VTAIL.n61 B 0.480331f
C189 VTAIL.n62 B 0.015287f
C190 VTAIL.t5 B 0.059121f
C191 VTAIL.n63 B 0.111698f
C192 VTAIL.n64 B 0.021324f
C193 VTAIL.n65 B 0.0271f
C194 VTAIL.n66 B 0.036133f
C195 VTAIL.n67 B 0.016186f
C196 VTAIL.n68 B 0.015287f
C197 VTAIL.n69 B 0.028449f
C198 VTAIL.n70 B 0.028449f
C199 VTAIL.n71 B 0.015287f
C200 VTAIL.n72 B 0.016186f
C201 VTAIL.n73 B 0.036133f
C202 VTAIL.n74 B 0.073471f
C203 VTAIL.n75 B 0.016186f
C204 VTAIL.n76 B 0.015287f
C205 VTAIL.n77 B 0.063426f
C206 VTAIL.n78 B 0.040548f
C207 VTAIL.n79 B 1.18703f
C208 VTAIL.n80 B 0.0373f
C209 VTAIL.n81 B 0.028449f
C210 VTAIL.n82 B 0.015287f
C211 VTAIL.n83 B 0.036133f
C212 VTAIL.n84 B 0.016186f
C213 VTAIL.n85 B 0.480331f
C214 VTAIL.n86 B 0.015287f
C215 VTAIL.t7 B 0.059121f
C216 VTAIL.n87 B 0.111698f
C217 VTAIL.n88 B 0.021324f
C218 VTAIL.n89 B 0.0271f
C219 VTAIL.n90 B 0.036133f
C220 VTAIL.n91 B 0.016186f
C221 VTAIL.n92 B 0.015287f
C222 VTAIL.n93 B 0.028449f
C223 VTAIL.n94 B 0.028449f
C224 VTAIL.n95 B 0.015287f
C225 VTAIL.n96 B 0.016186f
C226 VTAIL.n97 B 0.036133f
C227 VTAIL.n98 B 0.073471f
C228 VTAIL.n99 B 0.016186f
C229 VTAIL.n100 B 0.015287f
C230 VTAIL.n101 B 0.063426f
C231 VTAIL.n102 B 0.040548f
C232 VTAIL.n103 B 1.12895f
C233 VDD2.n0 B 0.028822f
C234 VDD2.n1 B 0.021982f
C235 VDD2.n2 B 0.011812f
C236 VDD2.n3 B 0.02792f
C237 VDD2.n4 B 0.012507f
C238 VDD2.n5 B 0.37115f
C239 VDD2.n6 B 0.011812f
C240 VDD2.t5 B 0.045682f
C241 VDD2.n7 B 0.086309f
C242 VDD2.n8 B 0.016477f
C243 VDD2.n9 B 0.02094f
C244 VDD2.n10 B 0.02792f
C245 VDD2.n11 B 0.012507f
C246 VDD2.n12 B 0.011812f
C247 VDD2.n13 B 0.021982f
C248 VDD2.n14 B 0.021982f
C249 VDD2.n15 B 0.011812f
C250 VDD2.n16 B 0.012507f
C251 VDD2.n17 B 0.02792f
C252 VDD2.n18 B 0.056771f
C253 VDD2.n19 B 0.012507f
C254 VDD2.n20 B 0.011812f
C255 VDD2.n21 B 0.049009f
C256 VDD2.n22 B 0.051939f
C257 VDD2.t3 B 0.07817f
C258 VDD2.t2 B 0.07817f
C259 VDD2.n23 B 0.629562f
C260 VDD2.n24 B 1.85101f
C261 VDD2.n25 B 0.028822f
C262 VDD2.n26 B 0.021982f
C263 VDD2.n27 B 0.011812f
C264 VDD2.n28 B 0.02792f
C265 VDD2.n29 B 0.012507f
C266 VDD2.n30 B 0.37115f
C267 VDD2.n31 B 0.011812f
C268 VDD2.t4 B 0.045682f
C269 VDD2.n32 B 0.086309f
C270 VDD2.n33 B 0.016477f
C271 VDD2.n34 B 0.02094f
C272 VDD2.n35 B 0.02792f
C273 VDD2.n36 B 0.012507f
C274 VDD2.n37 B 0.011812f
C275 VDD2.n38 B 0.021982f
C276 VDD2.n39 B 0.021982f
C277 VDD2.n40 B 0.011812f
C278 VDD2.n41 B 0.012507f
C279 VDD2.n42 B 0.02792f
C280 VDD2.n43 B 0.056771f
C281 VDD2.n44 B 0.012507f
C282 VDD2.n45 B 0.011812f
C283 VDD2.n46 B 0.049009f
C284 VDD2.n47 B 0.046525f
C285 VDD2.n48 B 1.66907f
C286 VDD2.t1 B 0.07817f
C287 VDD2.t0 B 0.07817f
C288 VDD2.n49 B 0.629538f
C289 VN.n0 B 0.038318f
C290 VN.t4 B 0.794194f
C291 VN.n1 B 0.035416f
C292 VN.n2 B 0.273084f
C293 VN.t1 B 0.794194f
C294 VN.t5 B 0.993634f
C295 VN.n3 B 0.375093f
C296 VN.n4 B 0.406501f
C297 VN.n5 B 0.0539f
C298 VN.n6 B 0.049087f
C299 VN.n7 B 0.029066f
C300 VN.n8 B 0.029066f
C301 VN.n9 B 0.029066f
C302 VN.n10 B 0.0539f
C303 VN.n11 B 0.036338f
C304 VN.n12 B 0.396636f
C305 VN.n13 B 0.045967f
C306 VN.n14 B 0.038318f
C307 VN.t3 B 0.794194f
C308 VN.n15 B 0.035416f
C309 VN.n16 B 0.273084f
C310 VN.t0 B 0.794194f
C311 VN.t2 B 0.993634f
C312 VN.n17 B 0.375093f
C313 VN.n18 B 0.406501f
C314 VN.n19 B 0.0539f
C315 VN.n20 B 0.049087f
C316 VN.n21 B 0.029066f
C317 VN.n22 B 0.029066f
C318 VN.n23 B 0.029066f
C319 VN.n24 B 0.0539f
C320 VN.n25 B 0.036338f
C321 VN.n26 B 0.396636f
C322 VN.n27 B 1.24568f
.ends

