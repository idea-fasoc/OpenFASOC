* NGSPICE file created from diff_pair_sample_1639.ext - technology: sky130A

.subckt diff_pair_sample_1639 VTAIL VN VP B VDD2 VDD1
X0 B.t17 B.t15 B.t16 B.t5 sky130_fd_pr__nfet_01v8 ad=3.7908 pd=20.22 as=0 ps=0 w=9.72 l=2.71
X1 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=3.7908 pd=20.22 as=0 ps=0 w=9.72 l=2.71
X2 VTAIL.t7 VN.t0 VDD2.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=3.7908 pd=20.22 as=1.6038 ps=10.05 w=9.72 l=2.71
X3 VTAIL.t0 VP.t0 VDD1.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=3.7908 pd=20.22 as=1.6038 ps=10.05 w=9.72 l=2.71
X4 VTAIL.t2 VP.t1 VDD1.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=3.7908 pd=20.22 as=1.6038 ps=10.05 w=9.72 l=2.71
X5 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=3.7908 pd=20.22 as=0 ps=0 w=9.72 l=2.71
X6 VDD1.t1 VP.t2 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.6038 pd=10.05 as=3.7908 ps=20.22 w=9.72 l=2.71
X7 VDD2.t0 VN.t1 VTAIL.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=1.6038 pd=10.05 as=3.7908 ps=20.22 w=9.72 l=2.71
X8 VDD2.t3 VN.t2 VTAIL.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=1.6038 pd=10.05 as=3.7908 ps=20.22 w=9.72 l=2.71
X9 VDD1.t0 VP.t3 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.6038 pd=10.05 as=3.7908 ps=20.22 w=9.72 l=2.71
X10 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=3.7908 pd=20.22 as=0 ps=0 w=9.72 l=2.71
X11 VTAIL.t4 VN.t3 VDD2.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=3.7908 pd=20.22 as=1.6038 ps=10.05 w=9.72 l=2.71
R0 B.n686 B.n685 585
R1 B.n687 B.n686 585
R2 B.n264 B.n106 585
R3 B.n263 B.n262 585
R4 B.n261 B.n260 585
R5 B.n259 B.n258 585
R6 B.n257 B.n256 585
R7 B.n255 B.n254 585
R8 B.n253 B.n252 585
R9 B.n251 B.n250 585
R10 B.n249 B.n248 585
R11 B.n247 B.n246 585
R12 B.n245 B.n244 585
R13 B.n243 B.n242 585
R14 B.n241 B.n240 585
R15 B.n239 B.n238 585
R16 B.n237 B.n236 585
R17 B.n235 B.n234 585
R18 B.n233 B.n232 585
R19 B.n231 B.n230 585
R20 B.n229 B.n228 585
R21 B.n227 B.n226 585
R22 B.n225 B.n224 585
R23 B.n223 B.n222 585
R24 B.n221 B.n220 585
R25 B.n219 B.n218 585
R26 B.n217 B.n216 585
R27 B.n215 B.n214 585
R28 B.n213 B.n212 585
R29 B.n211 B.n210 585
R30 B.n209 B.n208 585
R31 B.n207 B.n206 585
R32 B.n205 B.n204 585
R33 B.n203 B.n202 585
R34 B.n201 B.n200 585
R35 B.n199 B.n198 585
R36 B.n197 B.n196 585
R37 B.n195 B.n194 585
R38 B.n193 B.n192 585
R39 B.n191 B.n190 585
R40 B.n189 B.n188 585
R41 B.n187 B.n186 585
R42 B.n185 B.n184 585
R43 B.n183 B.n182 585
R44 B.n181 B.n180 585
R45 B.n178 B.n177 585
R46 B.n176 B.n175 585
R47 B.n174 B.n173 585
R48 B.n172 B.n171 585
R49 B.n170 B.n169 585
R50 B.n168 B.n167 585
R51 B.n166 B.n165 585
R52 B.n164 B.n163 585
R53 B.n162 B.n161 585
R54 B.n160 B.n159 585
R55 B.n158 B.n157 585
R56 B.n156 B.n155 585
R57 B.n154 B.n153 585
R58 B.n152 B.n151 585
R59 B.n150 B.n149 585
R60 B.n148 B.n147 585
R61 B.n146 B.n145 585
R62 B.n144 B.n143 585
R63 B.n142 B.n141 585
R64 B.n140 B.n139 585
R65 B.n138 B.n137 585
R66 B.n136 B.n135 585
R67 B.n134 B.n133 585
R68 B.n132 B.n131 585
R69 B.n130 B.n129 585
R70 B.n128 B.n127 585
R71 B.n126 B.n125 585
R72 B.n124 B.n123 585
R73 B.n122 B.n121 585
R74 B.n120 B.n119 585
R75 B.n118 B.n117 585
R76 B.n116 B.n115 585
R77 B.n114 B.n113 585
R78 B.n67 B.n66 585
R79 B.n690 B.n689 585
R80 B.n684 B.n107 585
R81 B.n107 B.n64 585
R82 B.n683 B.n63 585
R83 B.n694 B.n63 585
R84 B.n682 B.n62 585
R85 B.n695 B.n62 585
R86 B.n681 B.n61 585
R87 B.n696 B.n61 585
R88 B.n680 B.n679 585
R89 B.n679 B.n57 585
R90 B.n678 B.n56 585
R91 B.n702 B.n56 585
R92 B.n677 B.n55 585
R93 B.n703 B.n55 585
R94 B.n676 B.n54 585
R95 B.n704 B.n54 585
R96 B.n675 B.n674 585
R97 B.n674 B.n50 585
R98 B.n673 B.n49 585
R99 B.n710 B.n49 585
R100 B.n672 B.n48 585
R101 B.n711 B.n48 585
R102 B.n671 B.n47 585
R103 B.n712 B.n47 585
R104 B.n670 B.n669 585
R105 B.n669 B.n43 585
R106 B.n668 B.n42 585
R107 B.n718 B.n42 585
R108 B.n667 B.n41 585
R109 B.n719 B.n41 585
R110 B.n666 B.n40 585
R111 B.n720 B.n40 585
R112 B.n665 B.n664 585
R113 B.n664 B.n36 585
R114 B.n663 B.n35 585
R115 B.n726 B.n35 585
R116 B.n662 B.n34 585
R117 B.n727 B.n34 585
R118 B.n661 B.n33 585
R119 B.n728 B.n33 585
R120 B.n660 B.n659 585
R121 B.n659 B.n29 585
R122 B.n658 B.n28 585
R123 B.n734 B.n28 585
R124 B.n657 B.n27 585
R125 B.n735 B.n27 585
R126 B.n656 B.n26 585
R127 B.n736 B.n26 585
R128 B.n655 B.n654 585
R129 B.n654 B.n22 585
R130 B.n653 B.n21 585
R131 B.n742 B.n21 585
R132 B.n652 B.n20 585
R133 B.n743 B.n20 585
R134 B.n651 B.n19 585
R135 B.n744 B.n19 585
R136 B.n650 B.n649 585
R137 B.n649 B.n18 585
R138 B.n648 B.n14 585
R139 B.n750 B.n14 585
R140 B.n647 B.n13 585
R141 B.n751 B.n13 585
R142 B.n646 B.n12 585
R143 B.n752 B.n12 585
R144 B.n645 B.n644 585
R145 B.n644 B.n8 585
R146 B.n643 B.n7 585
R147 B.n758 B.n7 585
R148 B.n642 B.n6 585
R149 B.n759 B.n6 585
R150 B.n641 B.n5 585
R151 B.n760 B.n5 585
R152 B.n640 B.n639 585
R153 B.n639 B.n4 585
R154 B.n638 B.n265 585
R155 B.n638 B.n637 585
R156 B.n628 B.n266 585
R157 B.n267 B.n266 585
R158 B.n630 B.n629 585
R159 B.n631 B.n630 585
R160 B.n627 B.n272 585
R161 B.n272 B.n271 585
R162 B.n626 B.n625 585
R163 B.n625 B.n624 585
R164 B.n274 B.n273 585
R165 B.n617 B.n274 585
R166 B.n616 B.n615 585
R167 B.n618 B.n616 585
R168 B.n614 B.n279 585
R169 B.n279 B.n278 585
R170 B.n613 B.n612 585
R171 B.n612 B.n611 585
R172 B.n281 B.n280 585
R173 B.n282 B.n281 585
R174 B.n604 B.n603 585
R175 B.n605 B.n604 585
R176 B.n602 B.n287 585
R177 B.n287 B.n286 585
R178 B.n601 B.n600 585
R179 B.n600 B.n599 585
R180 B.n289 B.n288 585
R181 B.n290 B.n289 585
R182 B.n592 B.n591 585
R183 B.n593 B.n592 585
R184 B.n590 B.n295 585
R185 B.n295 B.n294 585
R186 B.n589 B.n588 585
R187 B.n588 B.n587 585
R188 B.n297 B.n296 585
R189 B.n298 B.n297 585
R190 B.n580 B.n579 585
R191 B.n581 B.n580 585
R192 B.n578 B.n303 585
R193 B.n303 B.n302 585
R194 B.n577 B.n576 585
R195 B.n576 B.n575 585
R196 B.n305 B.n304 585
R197 B.n306 B.n305 585
R198 B.n568 B.n567 585
R199 B.n569 B.n568 585
R200 B.n566 B.n311 585
R201 B.n311 B.n310 585
R202 B.n565 B.n564 585
R203 B.n564 B.n563 585
R204 B.n313 B.n312 585
R205 B.n314 B.n313 585
R206 B.n556 B.n555 585
R207 B.n557 B.n556 585
R208 B.n554 B.n319 585
R209 B.n319 B.n318 585
R210 B.n553 B.n552 585
R211 B.n552 B.n551 585
R212 B.n321 B.n320 585
R213 B.n322 B.n321 585
R214 B.n544 B.n543 585
R215 B.n545 B.n544 585
R216 B.n542 B.n327 585
R217 B.n327 B.n326 585
R218 B.n541 B.n540 585
R219 B.n540 B.n539 585
R220 B.n329 B.n328 585
R221 B.n330 B.n329 585
R222 B.n535 B.n534 585
R223 B.n333 B.n332 585
R224 B.n531 B.n530 585
R225 B.n532 B.n531 585
R226 B.n529 B.n372 585
R227 B.n528 B.n527 585
R228 B.n526 B.n525 585
R229 B.n524 B.n523 585
R230 B.n522 B.n521 585
R231 B.n520 B.n519 585
R232 B.n518 B.n517 585
R233 B.n516 B.n515 585
R234 B.n514 B.n513 585
R235 B.n512 B.n511 585
R236 B.n510 B.n509 585
R237 B.n508 B.n507 585
R238 B.n506 B.n505 585
R239 B.n504 B.n503 585
R240 B.n502 B.n501 585
R241 B.n500 B.n499 585
R242 B.n498 B.n497 585
R243 B.n496 B.n495 585
R244 B.n494 B.n493 585
R245 B.n492 B.n491 585
R246 B.n490 B.n489 585
R247 B.n488 B.n487 585
R248 B.n486 B.n485 585
R249 B.n484 B.n483 585
R250 B.n482 B.n481 585
R251 B.n480 B.n479 585
R252 B.n478 B.n477 585
R253 B.n476 B.n475 585
R254 B.n474 B.n473 585
R255 B.n472 B.n471 585
R256 B.n470 B.n469 585
R257 B.n468 B.n467 585
R258 B.n466 B.n465 585
R259 B.n464 B.n463 585
R260 B.n462 B.n461 585
R261 B.n460 B.n459 585
R262 B.n458 B.n457 585
R263 B.n456 B.n455 585
R264 B.n454 B.n453 585
R265 B.n452 B.n451 585
R266 B.n450 B.n449 585
R267 B.n447 B.n446 585
R268 B.n445 B.n444 585
R269 B.n443 B.n442 585
R270 B.n441 B.n440 585
R271 B.n439 B.n438 585
R272 B.n437 B.n436 585
R273 B.n435 B.n434 585
R274 B.n433 B.n432 585
R275 B.n431 B.n430 585
R276 B.n429 B.n428 585
R277 B.n427 B.n426 585
R278 B.n425 B.n424 585
R279 B.n423 B.n422 585
R280 B.n421 B.n420 585
R281 B.n419 B.n418 585
R282 B.n417 B.n416 585
R283 B.n415 B.n414 585
R284 B.n413 B.n412 585
R285 B.n411 B.n410 585
R286 B.n409 B.n408 585
R287 B.n407 B.n406 585
R288 B.n405 B.n404 585
R289 B.n403 B.n402 585
R290 B.n401 B.n400 585
R291 B.n399 B.n398 585
R292 B.n397 B.n396 585
R293 B.n395 B.n394 585
R294 B.n393 B.n392 585
R295 B.n391 B.n390 585
R296 B.n389 B.n388 585
R297 B.n387 B.n386 585
R298 B.n385 B.n384 585
R299 B.n383 B.n382 585
R300 B.n381 B.n380 585
R301 B.n379 B.n378 585
R302 B.n536 B.n331 585
R303 B.n331 B.n330 585
R304 B.n538 B.n537 585
R305 B.n539 B.n538 585
R306 B.n325 B.n324 585
R307 B.n326 B.n325 585
R308 B.n547 B.n546 585
R309 B.n546 B.n545 585
R310 B.n548 B.n323 585
R311 B.n323 B.n322 585
R312 B.n550 B.n549 585
R313 B.n551 B.n550 585
R314 B.n317 B.n316 585
R315 B.n318 B.n317 585
R316 B.n559 B.n558 585
R317 B.n558 B.n557 585
R318 B.n560 B.n315 585
R319 B.n315 B.n314 585
R320 B.n562 B.n561 585
R321 B.n563 B.n562 585
R322 B.n309 B.n308 585
R323 B.n310 B.n309 585
R324 B.n571 B.n570 585
R325 B.n570 B.n569 585
R326 B.n572 B.n307 585
R327 B.n307 B.n306 585
R328 B.n574 B.n573 585
R329 B.n575 B.n574 585
R330 B.n301 B.n300 585
R331 B.n302 B.n301 585
R332 B.n583 B.n582 585
R333 B.n582 B.n581 585
R334 B.n584 B.n299 585
R335 B.n299 B.n298 585
R336 B.n586 B.n585 585
R337 B.n587 B.n586 585
R338 B.n293 B.n292 585
R339 B.n294 B.n293 585
R340 B.n595 B.n594 585
R341 B.n594 B.n593 585
R342 B.n596 B.n291 585
R343 B.n291 B.n290 585
R344 B.n598 B.n597 585
R345 B.n599 B.n598 585
R346 B.n285 B.n284 585
R347 B.n286 B.n285 585
R348 B.n607 B.n606 585
R349 B.n606 B.n605 585
R350 B.n608 B.n283 585
R351 B.n283 B.n282 585
R352 B.n610 B.n609 585
R353 B.n611 B.n610 585
R354 B.n277 B.n276 585
R355 B.n278 B.n277 585
R356 B.n620 B.n619 585
R357 B.n619 B.n618 585
R358 B.n621 B.n275 585
R359 B.n617 B.n275 585
R360 B.n623 B.n622 585
R361 B.n624 B.n623 585
R362 B.n270 B.n269 585
R363 B.n271 B.n270 585
R364 B.n633 B.n632 585
R365 B.n632 B.n631 585
R366 B.n634 B.n268 585
R367 B.n268 B.n267 585
R368 B.n636 B.n635 585
R369 B.n637 B.n636 585
R370 B.n2 B.n0 585
R371 B.n4 B.n2 585
R372 B.n3 B.n1 585
R373 B.n759 B.n3 585
R374 B.n757 B.n756 585
R375 B.n758 B.n757 585
R376 B.n755 B.n9 585
R377 B.n9 B.n8 585
R378 B.n754 B.n753 585
R379 B.n753 B.n752 585
R380 B.n11 B.n10 585
R381 B.n751 B.n11 585
R382 B.n749 B.n748 585
R383 B.n750 B.n749 585
R384 B.n747 B.n15 585
R385 B.n18 B.n15 585
R386 B.n746 B.n745 585
R387 B.n745 B.n744 585
R388 B.n17 B.n16 585
R389 B.n743 B.n17 585
R390 B.n741 B.n740 585
R391 B.n742 B.n741 585
R392 B.n739 B.n23 585
R393 B.n23 B.n22 585
R394 B.n738 B.n737 585
R395 B.n737 B.n736 585
R396 B.n25 B.n24 585
R397 B.n735 B.n25 585
R398 B.n733 B.n732 585
R399 B.n734 B.n733 585
R400 B.n731 B.n30 585
R401 B.n30 B.n29 585
R402 B.n730 B.n729 585
R403 B.n729 B.n728 585
R404 B.n32 B.n31 585
R405 B.n727 B.n32 585
R406 B.n725 B.n724 585
R407 B.n726 B.n725 585
R408 B.n723 B.n37 585
R409 B.n37 B.n36 585
R410 B.n722 B.n721 585
R411 B.n721 B.n720 585
R412 B.n39 B.n38 585
R413 B.n719 B.n39 585
R414 B.n717 B.n716 585
R415 B.n718 B.n717 585
R416 B.n715 B.n44 585
R417 B.n44 B.n43 585
R418 B.n714 B.n713 585
R419 B.n713 B.n712 585
R420 B.n46 B.n45 585
R421 B.n711 B.n46 585
R422 B.n709 B.n708 585
R423 B.n710 B.n709 585
R424 B.n707 B.n51 585
R425 B.n51 B.n50 585
R426 B.n706 B.n705 585
R427 B.n705 B.n704 585
R428 B.n53 B.n52 585
R429 B.n703 B.n53 585
R430 B.n701 B.n700 585
R431 B.n702 B.n701 585
R432 B.n699 B.n58 585
R433 B.n58 B.n57 585
R434 B.n698 B.n697 585
R435 B.n697 B.n696 585
R436 B.n60 B.n59 585
R437 B.n695 B.n60 585
R438 B.n693 B.n692 585
R439 B.n694 B.n693 585
R440 B.n691 B.n65 585
R441 B.n65 B.n64 585
R442 B.n762 B.n761 585
R443 B.n761 B.n760 585
R444 B.n534 B.n331 521.33
R445 B.n689 B.n65 521.33
R446 B.n378 B.n329 521.33
R447 B.n686 B.n107 521.33
R448 B.n376 B.t12 294.647
R449 B.n373 B.t8 294.647
R450 B.n111 B.t15 294.647
R451 B.n108 B.t4 294.647
R452 B.n687 B.n105 256.663
R453 B.n687 B.n104 256.663
R454 B.n687 B.n103 256.663
R455 B.n687 B.n102 256.663
R456 B.n687 B.n101 256.663
R457 B.n687 B.n100 256.663
R458 B.n687 B.n99 256.663
R459 B.n687 B.n98 256.663
R460 B.n687 B.n97 256.663
R461 B.n687 B.n96 256.663
R462 B.n687 B.n95 256.663
R463 B.n687 B.n94 256.663
R464 B.n687 B.n93 256.663
R465 B.n687 B.n92 256.663
R466 B.n687 B.n91 256.663
R467 B.n687 B.n90 256.663
R468 B.n687 B.n89 256.663
R469 B.n687 B.n88 256.663
R470 B.n687 B.n87 256.663
R471 B.n687 B.n86 256.663
R472 B.n687 B.n85 256.663
R473 B.n687 B.n84 256.663
R474 B.n687 B.n83 256.663
R475 B.n687 B.n82 256.663
R476 B.n687 B.n81 256.663
R477 B.n687 B.n80 256.663
R478 B.n687 B.n79 256.663
R479 B.n687 B.n78 256.663
R480 B.n687 B.n77 256.663
R481 B.n687 B.n76 256.663
R482 B.n687 B.n75 256.663
R483 B.n687 B.n74 256.663
R484 B.n687 B.n73 256.663
R485 B.n687 B.n72 256.663
R486 B.n687 B.n71 256.663
R487 B.n687 B.n70 256.663
R488 B.n687 B.n69 256.663
R489 B.n687 B.n68 256.663
R490 B.n688 B.n687 256.663
R491 B.n533 B.n532 256.663
R492 B.n532 B.n334 256.663
R493 B.n532 B.n335 256.663
R494 B.n532 B.n336 256.663
R495 B.n532 B.n337 256.663
R496 B.n532 B.n338 256.663
R497 B.n532 B.n339 256.663
R498 B.n532 B.n340 256.663
R499 B.n532 B.n341 256.663
R500 B.n532 B.n342 256.663
R501 B.n532 B.n343 256.663
R502 B.n532 B.n344 256.663
R503 B.n532 B.n345 256.663
R504 B.n532 B.n346 256.663
R505 B.n532 B.n347 256.663
R506 B.n532 B.n348 256.663
R507 B.n532 B.n349 256.663
R508 B.n532 B.n350 256.663
R509 B.n532 B.n351 256.663
R510 B.n532 B.n352 256.663
R511 B.n532 B.n353 256.663
R512 B.n532 B.n354 256.663
R513 B.n532 B.n355 256.663
R514 B.n532 B.n356 256.663
R515 B.n532 B.n357 256.663
R516 B.n532 B.n358 256.663
R517 B.n532 B.n359 256.663
R518 B.n532 B.n360 256.663
R519 B.n532 B.n361 256.663
R520 B.n532 B.n362 256.663
R521 B.n532 B.n363 256.663
R522 B.n532 B.n364 256.663
R523 B.n532 B.n365 256.663
R524 B.n532 B.n366 256.663
R525 B.n532 B.n367 256.663
R526 B.n532 B.n368 256.663
R527 B.n532 B.n369 256.663
R528 B.n532 B.n370 256.663
R529 B.n532 B.n371 256.663
R530 B.n538 B.n331 163.367
R531 B.n538 B.n325 163.367
R532 B.n546 B.n325 163.367
R533 B.n546 B.n323 163.367
R534 B.n550 B.n323 163.367
R535 B.n550 B.n317 163.367
R536 B.n558 B.n317 163.367
R537 B.n558 B.n315 163.367
R538 B.n562 B.n315 163.367
R539 B.n562 B.n309 163.367
R540 B.n570 B.n309 163.367
R541 B.n570 B.n307 163.367
R542 B.n574 B.n307 163.367
R543 B.n574 B.n301 163.367
R544 B.n582 B.n301 163.367
R545 B.n582 B.n299 163.367
R546 B.n586 B.n299 163.367
R547 B.n586 B.n293 163.367
R548 B.n594 B.n293 163.367
R549 B.n594 B.n291 163.367
R550 B.n598 B.n291 163.367
R551 B.n598 B.n285 163.367
R552 B.n606 B.n285 163.367
R553 B.n606 B.n283 163.367
R554 B.n610 B.n283 163.367
R555 B.n610 B.n277 163.367
R556 B.n619 B.n277 163.367
R557 B.n619 B.n275 163.367
R558 B.n623 B.n275 163.367
R559 B.n623 B.n270 163.367
R560 B.n632 B.n270 163.367
R561 B.n632 B.n268 163.367
R562 B.n636 B.n268 163.367
R563 B.n636 B.n2 163.367
R564 B.n761 B.n2 163.367
R565 B.n761 B.n3 163.367
R566 B.n757 B.n3 163.367
R567 B.n757 B.n9 163.367
R568 B.n753 B.n9 163.367
R569 B.n753 B.n11 163.367
R570 B.n749 B.n11 163.367
R571 B.n749 B.n15 163.367
R572 B.n745 B.n15 163.367
R573 B.n745 B.n17 163.367
R574 B.n741 B.n17 163.367
R575 B.n741 B.n23 163.367
R576 B.n737 B.n23 163.367
R577 B.n737 B.n25 163.367
R578 B.n733 B.n25 163.367
R579 B.n733 B.n30 163.367
R580 B.n729 B.n30 163.367
R581 B.n729 B.n32 163.367
R582 B.n725 B.n32 163.367
R583 B.n725 B.n37 163.367
R584 B.n721 B.n37 163.367
R585 B.n721 B.n39 163.367
R586 B.n717 B.n39 163.367
R587 B.n717 B.n44 163.367
R588 B.n713 B.n44 163.367
R589 B.n713 B.n46 163.367
R590 B.n709 B.n46 163.367
R591 B.n709 B.n51 163.367
R592 B.n705 B.n51 163.367
R593 B.n705 B.n53 163.367
R594 B.n701 B.n53 163.367
R595 B.n701 B.n58 163.367
R596 B.n697 B.n58 163.367
R597 B.n697 B.n60 163.367
R598 B.n693 B.n60 163.367
R599 B.n693 B.n65 163.367
R600 B.n531 B.n333 163.367
R601 B.n531 B.n372 163.367
R602 B.n527 B.n526 163.367
R603 B.n523 B.n522 163.367
R604 B.n519 B.n518 163.367
R605 B.n515 B.n514 163.367
R606 B.n511 B.n510 163.367
R607 B.n507 B.n506 163.367
R608 B.n503 B.n502 163.367
R609 B.n499 B.n498 163.367
R610 B.n495 B.n494 163.367
R611 B.n491 B.n490 163.367
R612 B.n487 B.n486 163.367
R613 B.n483 B.n482 163.367
R614 B.n479 B.n478 163.367
R615 B.n475 B.n474 163.367
R616 B.n471 B.n470 163.367
R617 B.n467 B.n466 163.367
R618 B.n463 B.n462 163.367
R619 B.n459 B.n458 163.367
R620 B.n455 B.n454 163.367
R621 B.n451 B.n450 163.367
R622 B.n446 B.n445 163.367
R623 B.n442 B.n441 163.367
R624 B.n438 B.n437 163.367
R625 B.n434 B.n433 163.367
R626 B.n430 B.n429 163.367
R627 B.n426 B.n425 163.367
R628 B.n422 B.n421 163.367
R629 B.n418 B.n417 163.367
R630 B.n414 B.n413 163.367
R631 B.n410 B.n409 163.367
R632 B.n406 B.n405 163.367
R633 B.n402 B.n401 163.367
R634 B.n398 B.n397 163.367
R635 B.n394 B.n393 163.367
R636 B.n390 B.n389 163.367
R637 B.n386 B.n385 163.367
R638 B.n382 B.n381 163.367
R639 B.n540 B.n329 163.367
R640 B.n540 B.n327 163.367
R641 B.n544 B.n327 163.367
R642 B.n544 B.n321 163.367
R643 B.n552 B.n321 163.367
R644 B.n552 B.n319 163.367
R645 B.n556 B.n319 163.367
R646 B.n556 B.n313 163.367
R647 B.n564 B.n313 163.367
R648 B.n564 B.n311 163.367
R649 B.n568 B.n311 163.367
R650 B.n568 B.n305 163.367
R651 B.n576 B.n305 163.367
R652 B.n576 B.n303 163.367
R653 B.n580 B.n303 163.367
R654 B.n580 B.n297 163.367
R655 B.n588 B.n297 163.367
R656 B.n588 B.n295 163.367
R657 B.n592 B.n295 163.367
R658 B.n592 B.n289 163.367
R659 B.n600 B.n289 163.367
R660 B.n600 B.n287 163.367
R661 B.n604 B.n287 163.367
R662 B.n604 B.n281 163.367
R663 B.n612 B.n281 163.367
R664 B.n612 B.n279 163.367
R665 B.n616 B.n279 163.367
R666 B.n616 B.n274 163.367
R667 B.n625 B.n274 163.367
R668 B.n625 B.n272 163.367
R669 B.n630 B.n272 163.367
R670 B.n630 B.n266 163.367
R671 B.n638 B.n266 163.367
R672 B.n639 B.n638 163.367
R673 B.n639 B.n5 163.367
R674 B.n6 B.n5 163.367
R675 B.n7 B.n6 163.367
R676 B.n644 B.n7 163.367
R677 B.n644 B.n12 163.367
R678 B.n13 B.n12 163.367
R679 B.n14 B.n13 163.367
R680 B.n649 B.n14 163.367
R681 B.n649 B.n19 163.367
R682 B.n20 B.n19 163.367
R683 B.n21 B.n20 163.367
R684 B.n654 B.n21 163.367
R685 B.n654 B.n26 163.367
R686 B.n27 B.n26 163.367
R687 B.n28 B.n27 163.367
R688 B.n659 B.n28 163.367
R689 B.n659 B.n33 163.367
R690 B.n34 B.n33 163.367
R691 B.n35 B.n34 163.367
R692 B.n664 B.n35 163.367
R693 B.n664 B.n40 163.367
R694 B.n41 B.n40 163.367
R695 B.n42 B.n41 163.367
R696 B.n669 B.n42 163.367
R697 B.n669 B.n47 163.367
R698 B.n48 B.n47 163.367
R699 B.n49 B.n48 163.367
R700 B.n674 B.n49 163.367
R701 B.n674 B.n54 163.367
R702 B.n55 B.n54 163.367
R703 B.n56 B.n55 163.367
R704 B.n679 B.n56 163.367
R705 B.n679 B.n61 163.367
R706 B.n62 B.n61 163.367
R707 B.n63 B.n62 163.367
R708 B.n107 B.n63 163.367
R709 B.n113 B.n67 163.367
R710 B.n117 B.n116 163.367
R711 B.n121 B.n120 163.367
R712 B.n125 B.n124 163.367
R713 B.n129 B.n128 163.367
R714 B.n133 B.n132 163.367
R715 B.n137 B.n136 163.367
R716 B.n141 B.n140 163.367
R717 B.n145 B.n144 163.367
R718 B.n149 B.n148 163.367
R719 B.n153 B.n152 163.367
R720 B.n157 B.n156 163.367
R721 B.n161 B.n160 163.367
R722 B.n165 B.n164 163.367
R723 B.n169 B.n168 163.367
R724 B.n173 B.n172 163.367
R725 B.n177 B.n176 163.367
R726 B.n182 B.n181 163.367
R727 B.n186 B.n185 163.367
R728 B.n190 B.n189 163.367
R729 B.n194 B.n193 163.367
R730 B.n198 B.n197 163.367
R731 B.n202 B.n201 163.367
R732 B.n206 B.n205 163.367
R733 B.n210 B.n209 163.367
R734 B.n214 B.n213 163.367
R735 B.n218 B.n217 163.367
R736 B.n222 B.n221 163.367
R737 B.n226 B.n225 163.367
R738 B.n230 B.n229 163.367
R739 B.n234 B.n233 163.367
R740 B.n238 B.n237 163.367
R741 B.n242 B.n241 163.367
R742 B.n246 B.n245 163.367
R743 B.n250 B.n249 163.367
R744 B.n254 B.n253 163.367
R745 B.n258 B.n257 163.367
R746 B.n262 B.n261 163.367
R747 B.n686 B.n106 163.367
R748 B.n376 B.t14 131.01
R749 B.n108 B.t6 131.01
R750 B.n373 B.t11 130.999
R751 B.n111 B.t16 130.999
R752 B.n532 B.n330 87.2963
R753 B.n687 B.n64 87.2963
R754 B.n377 B.t13 72.0523
R755 B.n109 B.t7 72.0523
R756 B.n374 B.t10 72.0405
R757 B.n112 B.t17 72.0405
R758 B.n534 B.n533 71.676
R759 B.n372 B.n334 71.676
R760 B.n526 B.n335 71.676
R761 B.n522 B.n336 71.676
R762 B.n518 B.n337 71.676
R763 B.n514 B.n338 71.676
R764 B.n510 B.n339 71.676
R765 B.n506 B.n340 71.676
R766 B.n502 B.n341 71.676
R767 B.n498 B.n342 71.676
R768 B.n494 B.n343 71.676
R769 B.n490 B.n344 71.676
R770 B.n486 B.n345 71.676
R771 B.n482 B.n346 71.676
R772 B.n478 B.n347 71.676
R773 B.n474 B.n348 71.676
R774 B.n470 B.n349 71.676
R775 B.n466 B.n350 71.676
R776 B.n462 B.n351 71.676
R777 B.n458 B.n352 71.676
R778 B.n454 B.n353 71.676
R779 B.n450 B.n354 71.676
R780 B.n445 B.n355 71.676
R781 B.n441 B.n356 71.676
R782 B.n437 B.n357 71.676
R783 B.n433 B.n358 71.676
R784 B.n429 B.n359 71.676
R785 B.n425 B.n360 71.676
R786 B.n421 B.n361 71.676
R787 B.n417 B.n362 71.676
R788 B.n413 B.n363 71.676
R789 B.n409 B.n364 71.676
R790 B.n405 B.n365 71.676
R791 B.n401 B.n366 71.676
R792 B.n397 B.n367 71.676
R793 B.n393 B.n368 71.676
R794 B.n389 B.n369 71.676
R795 B.n385 B.n370 71.676
R796 B.n381 B.n371 71.676
R797 B.n689 B.n688 71.676
R798 B.n113 B.n68 71.676
R799 B.n117 B.n69 71.676
R800 B.n121 B.n70 71.676
R801 B.n125 B.n71 71.676
R802 B.n129 B.n72 71.676
R803 B.n133 B.n73 71.676
R804 B.n137 B.n74 71.676
R805 B.n141 B.n75 71.676
R806 B.n145 B.n76 71.676
R807 B.n149 B.n77 71.676
R808 B.n153 B.n78 71.676
R809 B.n157 B.n79 71.676
R810 B.n161 B.n80 71.676
R811 B.n165 B.n81 71.676
R812 B.n169 B.n82 71.676
R813 B.n173 B.n83 71.676
R814 B.n177 B.n84 71.676
R815 B.n182 B.n85 71.676
R816 B.n186 B.n86 71.676
R817 B.n190 B.n87 71.676
R818 B.n194 B.n88 71.676
R819 B.n198 B.n89 71.676
R820 B.n202 B.n90 71.676
R821 B.n206 B.n91 71.676
R822 B.n210 B.n92 71.676
R823 B.n214 B.n93 71.676
R824 B.n218 B.n94 71.676
R825 B.n222 B.n95 71.676
R826 B.n226 B.n96 71.676
R827 B.n230 B.n97 71.676
R828 B.n234 B.n98 71.676
R829 B.n238 B.n99 71.676
R830 B.n242 B.n100 71.676
R831 B.n246 B.n101 71.676
R832 B.n250 B.n102 71.676
R833 B.n254 B.n103 71.676
R834 B.n258 B.n104 71.676
R835 B.n262 B.n105 71.676
R836 B.n106 B.n105 71.676
R837 B.n261 B.n104 71.676
R838 B.n257 B.n103 71.676
R839 B.n253 B.n102 71.676
R840 B.n249 B.n101 71.676
R841 B.n245 B.n100 71.676
R842 B.n241 B.n99 71.676
R843 B.n237 B.n98 71.676
R844 B.n233 B.n97 71.676
R845 B.n229 B.n96 71.676
R846 B.n225 B.n95 71.676
R847 B.n221 B.n94 71.676
R848 B.n217 B.n93 71.676
R849 B.n213 B.n92 71.676
R850 B.n209 B.n91 71.676
R851 B.n205 B.n90 71.676
R852 B.n201 B.n89 71.676
R853 B.n197 B.n88 71.676
R854 B.n193 B.n87 71.676
R855 B.n189 B.n86 71.676
R856 B.n185 B.n85 71.676
R857 B.n181 B.n84 71.676
R858 B.n176 B.n83 71.676
R859 B.n172 B.n82 71.676
R860 B.n168 B.n81 71.676
R861 B.n164 B.n80 71.676
R862 B.n160 B.n79 71.676
R863 B.n156 B.n78 71.676
R864 B.n152 B.n77 71.676
R865 B.n148 B.n76 71.676
R866 B.n144 B.n75 71.676
R867 B.n140 B.n74 71.676
R868 B.n136 B.n73 71.676
R869 B.n132 B.n72 71.676
R870 B.n128 B.n71 71.676
R871 B.n124 B.n70 71.676
R872 B.n120 B.n69 71.676
R873 B.n116 B.n68 71.676
R874 B.n688 B.n67 71.676
R875 B.n533 B.n333 71.676
R876 B.n527 B.n334 71.676
R877 B.n523 B.n335 71.676
R878 B.n519 B.n336 71.676
R879 B.n515 B.n337 71.676
R880 B.n511 B.n338 71.676
R881 B.n507 B.n339 71.676
R882 B.n503 B.n340 71.676
R883 B.n499 B.n341 71.676
R884 B.n495 B.n342 71.676
R885 B.n491 B.n343 71.676
R886 B.n487 B.n344 71.676
R887 B.n483 B.n345 71.676
R888 B.n479 B.n346 71.676
R889 B.n475 B.n347 71.676
R890 B.n471 B.n348 71.676
R891 B.n467 B.n349 71.676
R892 B.n463 B.n350 71.676
R893 B.n459 B.n351 71.676
R894 B.n455 B.n352 71.676
R895 B.n451 B.n353 71.676
R896 B.n446 B.n354 71.676
R897 B.n442 B.n355 71.676
R898 B.n438 B.n356 71.676
R899 B.n434 B.n357 71.676
R900 B.n430 B.n358 71.676
R901 B.n426 B.n359 71.676
R902 B.n422 B.n360 71.676
R903 B.n418 B.n361 71.676
R904 B.n414 B.n362 71.676
R905 B.n410 B.n363 71.676
R906 B.n406 B.n364 71.676
R907 B.n402 B.n365 71.676
R908 B.n398 B.n366 71.676
R909 B.n394 B.n367 71.676
R910 B.n390 B.n368 71.676
R911 B.n386 B.n369 71.676
R912 B.n382 B.n370 71.676
R913 B.n378 B.n371 71.676
R914 B.n448 B.n377 59.5399
R915 B.n375 B.n374 59.5399
R916 B.n179 B.n112 59.5399
R917 B.n110 B.n109 59.5399
R918 B.n377 B.n376 58.9581
R919 B.n374 B.n373 58.9581
R920 B.n112 B.n111 58.9581
R921 B.n109 B.n108 58.9581
R922 B.n539 B.n330 49.8838
R923 B.n539 B.n326 49.8838
R924 B.n545 B.n326 49.8838
R925 B.n545 B.n322 49.8838
R926 B.n551 B.n322 49.8838
R927 B.n551 B.n318 49.8838
R928 B.n557 B.n318 49.8838
R929 B.n563 B.n314 49.8838
R930 B.n563 B.n310 49.8838
R931 B.n569 B.n310 49.8838
R932 B.n569 B.n306 49.8838
R933 B.n575 B.n306 49.8838
R934 B.n575 B.n302 49.8838
R935 B.n581 B.n302 49.8838
R936 B.n581 B.n298 49.8838
R937 B.n587 B.n298 49.8838
R938 B.n587 B.n294 49.8838
R939 B.n593 B.n294 49.8838
R940 B.n599 B.n290 49.8838
R941 B.n599 B.n286 49.8838
R942 B.n605 B.n286 49.8838
R943 B.n605 B.n282 49.8838
R944 B.n611 B.n282 49.8838
R945 B.n611 B.n278 49.8838
R946 B.n618 B.n278 49.8838
R947 B.n618 B.n617 49.8838
R948 B.n624 B.n271 49.8838
R949 B.n631 B.n271 49.8838
R950 B.n631 B.n267 49.8838
R951 B.n637 B.n267 49.8838
R952 B.n637 B.n4 49.8838
R953 B.n760 B.n4 49.8838
R954 B.n760 B.n759 49.8838
R955 B.n759 B.n758 49.8838
R956 B.n758 B.n8 49.8838
R957 B.n752 B.n8 49.8838
R958 B.n752 B.n751 49.8838
R959 B.n751 B.n750 49.8838
R960 B.n744 B.n18 49.8838
R961 B.n744 B.n743 49.8838
R962 B.n743 B.n742 49.8838
R963 B.n742 B.n22 49.8838
R964 B.n736 B.n22 49.8838
R965 B.n736 B.n735 49.8838
R966 B.n735 B.n734 49.8838
R967 B.n734 B.n29 49.8838
R968 B.n728 B.n727 49.8838
R969 B.n727 B.n726 49.8838
R970 B.n726 B.n36 49.8838
R971 B.n720 B.n36 49.8838
R972 B.n720 B.n719 49.8838
R973 B.n719 B.n718 49.8838
R974 B.n718 B.n43 49.8838
R975 B.n712 B.n43 49.8838
R976 B.n712 B.n711 49.8838
R977 B.n711 B.n710 49.8838
R978 B.n710 B.n50 49.8838
R979 B.n704 B.n703 49.8838
R980 B.n703 B.n702 49.8838
R981 B.n702 B.n57 49.8838
R982 B.n696 B.n57 49.8838
R983 B.n696 B.n695 49.8838
R984 B.n695 B.n694 49.8838
R985 B.n694 B.n64 49.8838
R986 B.n593 B.t2 49.1502
R987 B.n728 B.t3 49.1502
R988 B.n617 B.t1 46.2159
R989 B.n18 B.t0 46.2159
R990 B.n557 B.t9 41.8144
R991 B.n704 B.t5 41.8144
R992 B.n691 B.n690 33.8737
R993 B.n685 B.n684 33.8737
R994 B.n379 B.n328 33.8737
R995 B.n536 B.n535 33.8737
R996 B B.n762 18.0485
R997 B.n690 B.n66 10.6151
R998 B.n114 B.n66 10.6151
R999 B.n115 B.n114 10.6151
R1000 B.n118 B.n115 10.6151
R1001 B.n119 B.n118 10.6151
R1002 B.n122 B.n119 10.6151
R1003 B.n123 B.n122 10.6151
R1004 B.n126 B.n123 10.6151
R1005 B.n127 B.n126 10.6151
R1006 B.n130 B.n127 10.6151
R1007 B.n131 B.n130 10.6151
R1008 B.n134 B.n131 10.6151
R1009 B.n135 B.n134 10.6151
R1010 B.n138 B.n135 10.6151
R1011 B.n139 B.n138 10.6151
R1012 B.n142 B.n139 10.6151
R1013 B.n143 B.n142 10.6151
R1014 B.n146 B.n143 10.6151
R1015 B.n147 B.n146 10.6151
R1016 B.n150 B.n147 10.6151
R1017 B.n151 B.n150 10.6151
R1018 B.n154 B.n151 10.6151
R1019 B.n155 B.n154 10.6151
R1020 B.n158 B.n155 10.6151
R1021 B.n159 B.n158 10.6151
R1022 B.n162 B.n159 10.6151
R1023 B.n163 B.n162 10.6151
R1024 B.n166 B.n163 10.6151
R1025 B.n167 B.n166 10.6151
R1026 B.n170 B.n167 10.6151
R1027 B.n171 B.n170 10.6151
R1028 B.n174 B.n171 10.6151
R1029 B.n175 B.n174 10.6151
R1030 B.n178 B.n175 10.6151
R1031 B.n183 B.n180 10.6151
R1032 B.n184 B.n183 10.6151
R1033 B.n187 B.n184 10.6151
R1034 B.n188 B.n187 10.6151
R1035 B.n191 B.n188 10.6151
R1036 B.n192 B.n191 10.6151
R1037 B.n195 B.n192 10.6151
R1038 B.n196 B.n195 10.6151
R1039 B.n200 B.n199 10.6151
R1040 B.n203 B.n200 10.6151
R1041 B.n204 B.n203 10.6151
R1042 B.n207 B.n204 10.6151
R1043 B.n208 B.n207 10.6151
R1044 B.n211 B.n208 10.6151
R1045 B.n212 B.n211 10.6151
R1046 B.n215 B.n212 10.6151
R1047 B.n216 B.n215 10.6151
R1048 B.n219 B.n216 10.6151
R1049 B.n220 B.n219 10.6151
R1050 B.n223 B.n220 10.6151
R1051 B.n224 B.n223 10.6151
R1052 B.n227 B.n224 10.6151
R1053 B.n228 B.n227 10.6151
R1054 B.n231 B.n228 10.6151
R1055 B.n232 B.n231 10.6151
R1056 B.n235 B.n232 10.6151
R1057 B.n236 B.n235 10.6151
R1058 B.n239 B.n236 10.6151
R1059 B.n240 B.n239 10.6151
R1060 B.n243 B.n240 10.6151
R1061 B.n244 B.n243 10.6151
R1062 B.n247 B.n244 10.6151
R1063 B.n248 B.n247 10.6151
R1064 B.n251 B.n248 10.6151
R1065 B.n252 B.n251 10.6151
R1066 B.n255 B.n252 10.6151
R1067 B.n256 B.n255 10.6151
R1068 B.n259 B.n256 10.6151
R1069 B.n260 B.n259 10.6151
R1070 B.n263 B.n260 10.6151
R1071 B.n264 B.n263 10.6151
R1072 B.n685 B.n264 10.6151
R1073 B.n541 B.n328 10.6151
R1074 B.n542 B.n541 10.6151
R1075 B.n543 B.n542 10.6151
R1076 B.n543 B.n320 10.6151
R1077 B.n553 B.n320 10.6151
R1078 B.n554 B.n553 10.6151
R1079 B.n555 B.n554 10.6151
R1080 B.n555 B.n312 10.6151
R1081 B.n565 B.n312 10.6151
R1082 B.n566 B.n565 10.6151
R1083 B.n567 B.n566 10.6151
R1084 B.n567 B.n304 10.6151
R1085 B.n577 B.n304 10.6151
R1086 B.n578 B.n577 10.6151
R1087 B.n579 B.n578 10.6151
R1088 B.n579 B.n296 10.6151
R1089 B.n589 B.n296 10.6151
R1090 B.n590 B.n589 10.6151
R1091 B.n591 B.n590 10.6151
R1092 B.n591 B.n288 10.6151
R1093 B.n601 B.n288 10.6151
R1094 B.n602 B.n601 10.6151
R1095 B.n603 B.n602 10.6151
R1096 B.n603 B.n280 10.6151
R1097 B.n613 B.n280 10.6151
R1098 B.n614 B.n613 10.6151
R1099 B.n615 B.n614 10.6151
R1100 B.n615 B.n273 10.6151
R1101 B.n626 B.n273 10.6151
R1102 B.n627 B.n626 10.6151
R1103 B.n629 B.n627 10.6151
R1104 B.n629 B.n628 10.6151
R1105 B.n628 B.n265 10.6151
R1106 B.n640 B.n265 10.6151
R1107 B.n641 B.n640 10.6151
R1108 B.n642 B.n641 10.6151
R1109 B.n643 B.n642 10.6151
R1110 B.n645 B.n643 10.6151
R1111 B.n646 B.n645 10.6151
R1112 B.n647 B.n646 10.6151
R1113 B.n648 B.n647 10.6151
R1114 B.n650 B.n648 10.6151
R1115 B.n651 B.n650 10.6151
R1116 B.n652 B.n651 10.6151
R1117 B.n653 B.n652 10.6151
R1118 B.n655 B.n653 10.6151
R1119 B.n656 B.n655 10.6151
R1120 B.n657 B.n656 10.6151
R1121 B.n658 B.n657 10.6151
R1122 B.n660 B.n658 10.6151
R1123 B.n661 B.n660 10.6151
R1124 B.n662 B.n661 10.6151
R1125 B.n663 B.n662 10.6151
R1126 B.n665 B.n663 10.6151
R1127 B.n666 B.n665 10.6151
R1128 B.n667 B.n666 10.6151
R1129 B.n668 B.n667 10.6151
R1130 B.n670 B.n668 10.6151
R1131 B.n671 B.n670 10.6151
R1132 B.n672 B.n671 10.6151
R1133 B.n673 B.n672 10.6151
R1134 B.n675 B.n673 10.6151
R1135 B.n676 B.n675 10.6151
R1136 B.n677 B.n676 10.6151
R1137 B.n678 B.n677 10.6151
R1138 B.n680 B.n678 10.6151
R1139 B.n681 B.n680 10.6151
R1140 B.n682 B.n681 10.6151
R1141 B.n683 B.n682 10.6151
R1142 B.n684 B.n683 10.6151
R1143 B.n535 B.n332 10.6151
R1144 B.n530 B.n332 10.6151
R1145 B.n530 B.n529 10.6151
R1146 B.n529 B.n528 10.6151
R1147 B.n528 B.n525 10.6151
R1148 B.n525 B.n524 10.6151
R1149 B.n524 B.n521 10.6151
R1150 B.n521 B.n520 10.6151
R1151 B.n520 B.n517 10.6151
R1152 B.n517 B.n516 10.6151
R1153 B.n516 B.n513 10.6151
R1154 B.n513 B.n512 10.6151
R1155 B.n512 B.n509 10.6151
R1156 B.n509 B.n508 10.6151
R1157 B.n508 B.n505 10.6151
R1158 B.n505 B.n504 10.6151
R1159 B.n504 B.n501 10.6151
R1160 B.n501 B.n500 10.6151
R1161 B.n500 B.n497 10.6151
R1162 B.n497 B.n496 10.6151
R1163 B.n496 B.n493 10.6151
R1164 B.n493 B.n492 10.6151
R1165 B.n492 B.n489 10.6151
R1166 B.n489 B.n488 10.6151
R1167 B.n488 B.n485 10.6151
R1168 B.n485 B.n484 10.6151
R1169 B.n484 B.n481 10.6151
R1170 B.n481 B.n480 10.6151
R1171 B.n480 B.n477 10.6151
R1172 B.n477 B.n476 10.6151
R1173 B.n476 B.n473 10.6151
R1174 B.n473 B.n472 10.6151
R1175 B.n472 B.n469 10.6151
R1176 B.n469 B.n468 10.6151
R1177 B.n465 B.n464 10.6151
R1178 B.n464 B.n461 10.6151
R1179 B.n461 B.n460 10.6151
R1180 B.n460 B.n457 10.6151
R1181 B.n457 B.n456 10.6151
R1182 B.n456 B.n453 10.6151
R1183 B.n453 B.n452 10.6151
R1184 B.n452 B.n449 10.6151
R1185 B.n447 B.n444 10.6151
R1186 B.n444 B.n443 10.6151
R1187 B.n443 B.n440 10.6151
R1188 B.n440 B.n439 10.6151
R1189 B.n439 B.n436 10.6151
R1190 B.n436 B.n435 10.6151
R1191 B.n435 B.n432 10.6151
R1192 B.n432 B.n431 10.6151
R1193 B.n431 B.n428 10.6151
R1194 B.n428 B.n427 10.6151
R1195 B.n427 B.n424 10.6151
R1196 B.n424 B.n423 10.6151
R1197 B.n423 B.n420 10.6151
R1198 B.n420 B.n419 10.6151
R1199 B.n419 B.n416 10.6151
R1200 B.n416 B.n415 10.6151
R1201 B.n415 B.n412 10.6151
R1202 B.n412 B.n411 10.6151
R1203 B.n411 B.n408 10.6151
R1204 B.n408 B.n407 10.6151
R1205 B.n407 B.n404 10.6151
R1206 B.n404 B.n403 10.6151
R1207 B.n403 B.n400 10.6151
R1208 B.n400 B.n399 10.6151
R1209 B.n399 B.n396 10.6151
R1210 B.n396 B.n395 10.6151
R1211 B.n395 B.n392 10.6151
R1212 B.n392 B.n391 10.6151
R1213 B.n391 B.n388 10.6151
R1214 B.n388 B.n387 10.6151
R1215 B.n387 B.n384 10.6151
R1216 B.n384 B.n383 10.6151
R1217 B.n383 B.n380 10.6151
R1218 B.n380 B.n379 10.6151
R1219 B.n537 B.n536 10.6151
R1220 B.n537 B.n324 10.6151
R1221 B.n547 B.n324 10.6151
R1222 B.n548 B.n547 10.6151
R1223 B.n549 B.n548 10.6151
R1224 B.n549 B.n316 10.6151
R1225 B.n559 B.n316 10.6151
R1226 B.n560 B.n559 10.6151
R1227 B.n561 B.n560 10.6151
R1228 B.n561 B.n308 10.6151
R1229 B.n571 B.n308 10.6151
R1230 B.n572 B.n571 10.6151
R1231 B.n573 B.n572 10.6151
R1232 B.n573 B.n300 10.6151
R1233 B.n583 B.n300 10.6151
R1234 B.n584 B.n583 10.6151
R1235 B.n585 B.n584 10.6151
R1236 B.n585 B.n292 10.6151
R1237 B.n595 B.n292 10.6151
R1238 B.n596 B.n595 10.6151
R1239 B.n597 B.n596 10.6151
R1240 B.n597 B.n284 10.6151
R1241 B.n607 B.n284 10.6151
R1242 B.n608 B.n607 10.6151
R1243 B.n609 B.n608 10.6151
R1244 B.n609 B.n276 10.6151
R1245 B.n620 B.n276 10.6151
R1246 B.n621 B.n620 10.6151
R1247 B.n622 B.n621 10.6151
R1248 B.n622 B.n269 10.6151
R1249 B.n633 B.n269 10.6151
R1250 B.n634 B.n633 10.6151
R1251 B.n635 B.n634 10.6151
R1252 B.n635 B.n0 10.6151
R1253 B.n756 B.n1 10.6151
R1254 B.n756 B.n755 10.6151
R1255 B.n755 B.n754 10.6151
R1256 B.n754 B.n10 10.6151
R1257 B.n748 B.n10 10.6151
R1258 B.n748 B.n747 10.6151
R1259 B.n747 B.n746 10.6151
R1260 B.n746 B.n16 10.6151
R1261 B.n740 B.n16 10.6151
R1262 B.n740 B.n739 10.6151
R1263 B.n739 B.n738 10.6151
R1264 B.n738 B.n24 10.6151
R1265 B.n732 B.n24 10.6151
R1266 B.n732 B.n731 10.6151
R1267 B.n731 B.n730 10.6151
R1268 B.n730 B.n31 10.6151
R1269 B.n724 B.n31 10.6151
R1270 B.n724 B.n723 10.6151
R1271 B.n723 B.n722 10.6151
R1272 B.n722 B.n38 10.6151
R1273 B.n716 B.n38 10.6151
R1274 B.n716 B.n715 10.6151
R1275 B.n715 B.n714 10.6151
R1276 B.n714 B.n45 10.6151
R1277 B.n708 B.n45 10.6151
R1278 B.n708 B.n707 10.6151
R1279 B.n707 B.n706 10.6151
R1280 B.n706 B.n52 10.6151
R1281 B.n700 B.n52 10.6151
R1282 B.n700 B.n699 10.6151
R1283 B.n699 B.n698 10.6151
R1284 B.n698 B.n59 10.6151
R1285 B.n692 B.n59 10.6151
R1286 B.n692 B.n691 10.6151
R1287 B.t9 B.n314 8.06986
R1288 B.t5 B.n50 8.06986
R1289 B.n180 B.n179 6.5566
R1290 B.n196 B.n110 6.5566
R1291 B.n465 B.n375 6.5566
R1292 B.n449 B.n448 6.5566
R1293 B.n179 B.n178 4.05904
R1294 B.n199 B.n110 4.05904
R1295 B.n468 B.n375 4.05904
R1296 B.n448 B.n447 4.05904
R1297 B.n624 B.t1 3.66839
R1298 B.n750 B.t0 3.66839
R1299 B.n762 B.n0 2.81026
R1300 B.n762 B.n1 2.81026
R1301 B.t2 B.n290 0.734078
R1302 B.t3 B.n29 0.734078
R1303 VN.n0 VN.t3 120.481
R1304 VN.n1 VN.t1 120.481
R1305 VN.n0 VN.t2 119.611
R1306 VN.n1 VN.t0 119.611
R1307 VN VN.n1 48.7598
R1308 VN VN.n0 3.64997
R1309 VDD2.n2 VDD2.n0 105.096
R1310 VDD2.n2 VDD2.n1 65.1392
R1311 VDD2.n1 VDD2.t2 2.03754
R1312 VDD2.n1 VDD2.t0 2.03754
R1313 VDD2.n0 VDD2.t1 2.03754
R1314 VDD2.n0 VDD2.t3 2.03754
R1315 VDD2 VDD2.n2 0.0586897
R1316 VTAIL.n5 VTAIL.t0 50.4976
R1317 VTAIL.n4 VTAIL.t6 50.4976
R1318 VTAIL.n3 VTAIL.t7 50.4976
R1319 VTAIL.n7 VTAIL.t5 50.4975
R1320 VTAIL.n0 VTAIL.t4 50.4975
R1321 VTAIL.n1 VTAIL.t1 50.4975
R1322 VTAIL.n2 VTAIL.t2 50.4975
R1323 VTAIL.n6 VTAIL.t3 50.4975
R1324 VTAIL.n7 VTAIL.n6 23.3669
R1325 VTAIL.n3 VTAIL.n2 23.3669
R1326 VTAIL.n4 VTAIL.n3 2.62119
R1327 VTAIL.n6 VTAIL.n5 2.62119
R1328 VTAIL.n2 VTAIL.n1 2.62119
R1329 VTAIL VTAIL.n0 1.36903
R1330 VTAIL VTAIL.n7 1.25266
R1331 VTAIL.n5 VTAIL.n4 0.470328
R1332 VTAIL.n1 VTAIL.n0 0.470328
R1333 VP.n16 VP.n0 161.3
R1334 VP.n15 VP.n14 161.3
R1335 VP.n13 VP.n1 161.3
R1336 VP.n12 VP.n11 161.3
R1337 VP.n10 VP.n2 161.3
R1338 VP.n9 VP.n8 161.3
R1339 VP.n7 VP.n3 161.3
R1340 VP.n4 VP.t0 120.481
R1341 VP.n4 VP.t3 119.611
R1342 VP.n6 VP.n5 109.632
R1343 VP.n18 VP.n17 109.632
R1344 VP.n5 VP.t1 86.4403
R1345 VP.n17 VP.t2 86.4403
R1346 VP.n6 VP.n4 48.4809
R1347 VP.n11 VP.n10 40.4106
R1348 VP.n11 VP.n1 40.4106
R1349 VP.n9 VP.n3 24.3439
R1350 VP.n10 VP.n9 24.3439
R1351 VP.n15 VP.n1 24.3439
R1352 VP.n16 VP.n15 24.3439
R1353 VP.n5 VP.n3 0.974237
R1354 VP.n17 VP.n16 0.974237
R1355 VP.n7 VP.n6 0.278398
R1356 VP.n18 VP.n0 0.278398
R1357 VP.n8 VP.n7 0.189894
R1358 VP.n8 VP.n2 0.189894
R1359 VP.n12 VP.n2 0.189894
R1360 VP.n13 VP.n12 0.189894
R1361 VP.n14 VP.n13 0.189894
R1362 VP.n14 VP.n0 0.189894
R1363 VP VP.n18 0.153422
R1364 VDD1 VDD1.n1 105.621
R1365 VDD1 VDD1.n0 65.1974
R1366 VDD1.n0 VDD1.t3 2.03754
R1367 VDD1.n0 VDD1.t0 2.03754
R1368 VDD1.n1 VDD1.t2 2.03754
R1369 VDD1.n1 VDD1.t1 2.03754
C0 VDD1 VTAIL 4.89272f
C1 VDD1 VN 0.148601f
C2 VDD1 VDD2 1.04657f
C3 VTAIL VP 3.97602f
C4 VP VN 5.85514f
C5 VDD2 VP 0.400807f
C6 VTAIL VN 3.96191f
C7 VDD2 VTAIL 4.94767f
C8 VDD2 VN 3.93985f
C9 VDD1 VP 4.19129f
C10 VDD2 B 3.65667f
C11 VDD1 B 7.63375f
C12 VTAIL B 8.769053f
C13 VN B 10.731991f
C14 VP B 9.019561f
C15 VDD1.t3 B 0.210815f
C16 VDD1.t0 B 0.210815f
C17 VDD1.n0 B 1.85497f
C18 VDD1.t2 B 0.210815f
C19 VDD1.t1 B 0.210815f
C20 VDD1.n1 B 2.47278f
C21 VP.n0 B 0.034569f
C22 VP.t2 B 1.8691f
C23 VP.n1 B 0.052388f
C24 VP.n2 B 0.026219f
C25 VP.n3 B 0.025833f
C26 VP.t3 B 2.10237f
C27 VP.t0 B 2.10838f
C28 VP.n4 B 2.72066f
C29 VP.t1 B 1.8691f
C30 VP.n5 B 0.749148f
C31 VP.n6 B 1.37821f
C32 VP.n7 B 0.034569f
C33 VP.n8 B 0.026219f
C34 VP.n9 B 0.04911f
C35 VP.n10 B 0.052388f
C36 VP.n11 B 0.021217f
C37 VP.n12 B 0.026219f
C38 VP.n13 B 0.026219f
C39 VP.n14 B 0.026219f
C40 VP.n15 B 0.04911f
C41 VP.n16 B 0.025833f
C42 VP.n17 B 0.749148f
C43 VP.n18 B 0.048951f
C44 VTAIL.t4 B 1.42641f
C45 VTAIL.n0 B 0.318993f
C46 VTAIL.t1 B 1.42641f
C47 VTAIL.n1 B 0.388619f
C48 VTAIL.t2 B 1.42641f
C49 VTAIL.n2 B 1.20856f
C50 VTAIL.t7 B 1.42642f
C51 VTAIL.n3 B 1.20855f
C52 VTAIL.t6 B 1.42642f
C53 VTAIL.n4 B 0.388609f
C54 VTAIL.t0 B 1.42642f
C55 VTAIL.n5 B 0.388609f
C56 VTAIL.t3 B 1.42641f
C57 VTAIL.n6 B 1.20856f
C58 VTAIL.t5 B 1.42641f
C59 VTAIL.n7 B 1.13246f
C60 VDD2.t1 B 0.206161f
C61 VDD2.t3 B 0.206161f
C62 VDD2.n0 B 2.39297f
C63 VDD2.t2 B 0.206161f
C64 VDD2.t0 B 0.206161f
C65 VDD2.n1 B 1.81361f
C66 VDD2.n2 B 3.53635f
C67 VN.t3 B 2.05814f
C68 VN.t2 B 2.05228f
C69 VN.n0 B 1.31f
C70 VN.t1 B 2.05814f
C71 VN.t0 B 2.05228f
C72 VN.n1 B 2.66943f
.ends

