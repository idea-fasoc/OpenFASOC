* NGSPICE file created from diff_pair_sample_1073.ext - technology: sky130A

.subckt diff_pair_sample_1073 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=4.056 pd=21.58 as=0 ps=0 w=10.4 l=3.37
X1 B.t12 B.t10 B.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=4.056 pd=21.58 as=0 ps=0 w=10.4 l=3.37
X2 VDD1.t1 VP.t0 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=4.056 pd=21.58 as=4.056 ps=21.58 w=10.4 l=3.37
X3 VDD2.t1 VN.t0 VTAIL.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=4.056 pd=21.58 as=4.056 ps=21.58 w=10.4 l=3.37
X4 VDD2.t0 VN.t1 VTAIL.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=4.056 pd=21.58 as=4.056 ps=21.58 w=10.4 l=3.37
X5 VDD1.t0 VP.t1 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=4.056 pd=21.58 as=4.056 ps=21.58 w=10.4 l=3.37
X6 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=4.056 pd=21.58 as=0 ps=0 w=10.4 l=3.37
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=4.056 pd=21.58 as=0 ps=0 w=10.4 l=3.37
R0 B.n504 B.n104 585
R1 B.n104 B.n57 585
R2 B.n506 B.n505 585
R3 B.n508 B.n103 585
R4 B.n511 B.n510 585
R5 B.n512 B.n102 585
R6 B.n514 B.n513 585
R7 B.n516 B.n101 585
R8 B.n519 B.n518 585
R9 B.n520 B.n100 585
R10 B.n522 B.n521 585
R11 B.n524 B.n99 585
R12 B.n527 B.n526 585
R13 B.n528 B.n98 585
R14 B.n530 B.n529 585
R15 B.n532 B.n97 585
R16 B.n535 B.n534 585
R17 B.n536 B.n96 585
R18 B.n538 B.n537 585
R19 B.n540 B.n95 585
R20 B.n543 B.n542 585
R21 B.n544 B.n94 585
R22 B.n546 B.n545 585
R23 B.n548 B.n93 585
R24 B.n551 B.n550 585
R25 B.n552 B.n92 585
R26 B.n554 B.n553 585
R27 B.n556 B.n91 585
R28 B.n559 B.n558 585
R29 B.n560 B.n90 585
R30 B.n562 B.n561 585
R31 B.n564 B.n89 585
R32 B.n567 B.n566 585
R33 B.n568 B.n88 585
R34 B.n570 B.n569 585
R35 B.n572 B.n87 585
R36 B.n574 B.n573 585
R37 B.n576 B.n575 585
R38 B.n579 B.n578 585
R39 B.n580 B.n82 585
R40 B.n582 B.n581 585
R41 B.n584 B.n81 585
R42 B.n587 B.n586 585
R43 B.n588 B.n80 585
R44 B.n590 B.n589 585
R45 B.n592 B.n79 585
R46 B.n595 B.n594 585
R47 B.n597 B.n76 585
R48 B.n599 B.n598 585
R49 B.n601 B.n75 585
R50 B.n604 B.n603 585
R51 B.n605 B.n74 585
R52 B.n607 B.n606 585
R53 B.n609 B.n73 585
R54 B.n612 B.n611 585
R55 B.n613 B.n72 585
R56 B.n615 B.n614 585
R57 B.n617 B.n71 585
R58 B.n620 B.n619 585
R59 B.n621 B.n70 585
R60 B.n623 B.n622 585
R61 B.n625 B.n69 585
R62 B.n628 B.n627 585
R63 B.n629 B.n68 585
R64 B.n631 B.n630 585
R65 B.n633 B.n67 585
R66 B.n636 B.n635 585
R67 B.n637 B.n66 585
R68 B.n639 B.n638 585
R69 B.n641 B.n65 585
R70 B.n644 B.n643 585
R71 B.n645 B.n64 585
R72 B.n647 B.n646 585
R73 B.n649 B.n63 585
R74 B.n652 B.n651 585
R75 B.n653 B.n62 585
R76 B.n655 B.n654 585
R77 B.n657 B.n61 585
R78 B.n660 B.n659 585
R79 B.n661 B.n60 585
R80 B.n663 B.n662 585
R81 B.n665 B.n59 585
R82 B.n668 B.n667 585
R83 B.n669 B.n58 585
R84 B.n503 B.n56 585
R85 B.n672 B.n56 585
R86 B.n502 B.n55 585
R87 B.n673 B.n55 585
R88 B.n501 B.n54 585
R89 B.n674 B.n54 585
R90 B.n500 B.n499 585
R91 B.n499 B.n50 585
R92 B.n498 B.n49 585
R93 B.n680 B.n49 585
R94 B.n497 B.n48 585
R95 B.n681 B.n48 585
R96 B.n496 B.n47 585
R97 B.n682 B.n47 585
R98 B.n495 B.n494 585
R99 B.n494 B.n43 585
R100 B.n493 B.n42 585
R101 B.n688 B.n42 585
R102 B.n492 B.n41 585
R103 B.n689 B.n41 585
R104 B.n491 B.n40 585
R105 B.n690 B.n40 585
R106 B.n490 B.n489 585
R107 B.n489 B.n36 585
R108 B.n488 B.n35 585
R109 B.n696 B.n35 585
R110 B.n487 B.n34 585
R111 B.n697 B.n34 585
R112 B.n486 B.n33 585
R113 B.n698 B.n33 585
R114 B.n485 B.n484 585
R115 B.n484 B.n29 585
R116 B.n483 B.n28 585
R117 B.n704 B.n28 585
R118 B.n482 B.n27 585
R119 B.n705 B.n27 585
R120 B.n481 B.n26 585
R121 B.n706 B.n26 585
R122 B.n480 B.n479 585
R123 B.n479 B.n22 585
R124 B.n478 B.n21 585
R125 B.n712 B.n21 585
R126 B.n477 B.n20 585
R127 B.n713 B.n20 585
R128 B.n476 B.n19 585
R129 B.n714 B.n19 585
R130 B.n475 B.n474 585
R131 B.n474 B.n15 585
R132 B.n473 B.n14 585
R133 B.n720 B.n14 585
R134 B.n472 B.n13 585
R135 B.n721 B.n13 585
R136 B.n471 B.n12 585
R137 B.n722 B.n12 585
R138 B.n470 B.n469 585
R139 B.n469 B.n8 585
R140 B.n468 B.n7 585
R141 B.n728 B.n7 585
R142 B.n467 B.n6 585
R143 B.n729 B.n6 585
R144 B.n466 B.n5 585
R145 B.n730 B.n5 585
R146 B.n465 B.n464 585
R147 B.n464 B.n4 585
R148 B.n463 B.n105 585
R149 B.n463 B.n462 585
R150 B.n453 B.n106 585
R151 B.n107 B.n106 585
R152 B.n455 B.n454 585
R153 B.n456 B.n455 585
R154 B.n452 B.n112 585
R155 B.n112 B.n111 585
R156 B.n451 B.n450 585
R157 B.n450 B.n449 585
R158 B.n114 B.n113 585
R159 B.n115 B.n114 585
R160 B.n442 B.n441 585
R161 B.n443 B.n442 585
R162 B.n440 B.n120 585
R163 B.n120 B.n119 585
R164 B.n439 B.n438 585
R165 B.n438 B.n437 585
R166 B.n122 B.n121 585
R167 B.n123 B.n122 585
R168 B.n430 B.n429 585
R169 B.n431 B.n430 585
R170 B.n428 B.n128 585
R171 B.n128 B.n127 585
R172 B.n427 B.n426 585
R173 B.n426 B.n425 585
R174 B.n130 B.n129 585
R175 B.n131 B.n130 585
R176 B.n418 B.n417 585
R177 B.n419 B.n418 585
R178 B.n416 B.n136 585
R179 B.n136 B.n135 585
R180 B.n415 B.n414 585
R181 B.n414 B.n413 585
R182 B.n138 B.n137 585
R183 B.n139 B.n138 585
R184 B.n406 B.n405 585
R185 B.n407 B.n406 585
R186 B.n404 B.n144 585
R187 B.n144 B.n143 585
R188 B.n403 B.n402 585
R189 B.n402 B.n401 585
R190 B.n146 B.n145 585
R191 B.n147 B.n146 585
R192 B.n394 B.n393 585
R193 B.n395 B.n394 585
R194 B.n392 B.n152 585
R195 B.n152 B.n151 585
R196 B.n391 B.n390 585
R197 B.n390 B.n389 585
R198 B.n154 B.n153 585
R199 B.n155 B.n154 585
R200 B.n382 B.n381 585
R201 B.n383 B.n382 585
R202 B.n380 B.n160 585
R203 B.n160 B.n159 585
R204 B.n379 B.n378 585
R205 B.n378 B.n377 585
R206 B.n374 B.n164 585
R207 B.n373 B.n372 585
R208 B.n370 B.n165 585
R209 B.n370 B.n163 585
R210 B.n369 B.n368 585
R211 B.n367 B.n366 585
R212 B.n365 B.n167 585
R213 B.n363 B.n362 585
R214 B.n361 B.n168 585
R215 B.n360 B.n359 585
R216 B.n357 B.n169 585
R217 B.n355 B.n354 585
R218 B.n353 B.n170 585
R219 B.n352 B.n351 585
R220 B.n349 B.n171 585
R221 B.n347 B.n346 585
R222 B.n345 B.n172 585
R223 B.n344 B.n343 585
R224 B.n341 B.n173 585
R225 B.n339 B.n338 585
R226 B.n337 B.n174 585
R227 B.n336 B.n335 585
R228 B.n333 B.n175 585
R229 B.n331 B.n330 585
R230 B.n329 B.n176 585
R231 B.n328 B.n327 585
R232 B.n325 B.n177 585
R233 B.n323 B.n322 585
R234 B.n321 B.n178 585
R235 B.n320 B.n319 585
R236 B.n317 B.n179 585
R237 B.n315 B.n314 585
R238 B.n313 B.n180 585
R239 B.n312 B.n311 585
R240 B.n309 B.n181 585
R241 B.n307 B.n306 585
R242 B.n305 B.n182 585
R243 B.n304 B.n303 585
R244 B.n301 B.n300 585
R245 B.n299 B.n298 585
R246 B.n297 B.n187 585
R247 B.n295 B.n294 585
R248 B.n293 B.n188 585
R249 B.n292 B.n291 585
R250 B.n289 B.n189 585
R251 B.n287 B.n286 585
R252 B.n285 B.n190 585
R253 B.n283 B.n282 585
R254 B.n280 B.n193 585
R255 B.n278 B.n277 585
R256 B.n276 B.n194 585
R257 B.n275 B.n274 585
R258 B.n272 B.n195 585
R259 B.n270 B.n269 585
R260 B.n268 B.n196 585
R261 B.n267 B.n266 585
R262 B.n264 B.n197 585
R263 B.n262 B.n261 585
R264 B.n260 B.n198 585
R265 B.n259 B.n258 585
R266 B.n256 B.n199 585
R267 B.n254 B.n253 585
R268 B.n252 B.n200 585
R269 B.n251 B.n250 585
R270 B.n248 B.n201 585
R271 B.n246 B.n245 585
R272 B.n244 B.n202 585
R273 B.n243 B.n242 585
R274 B.n240 B.n203 585
R275 B.n238 B.n237 585
R276 B.n236 B.n204 585
R277 B.n235 B.n234 585
R278 B.n232 B.n205 585
R279 B.n230 B.n229 585
R280 B.n228 B.n206 585
R281 B.n227 B.n226 585
R282 B.n224 B.n207 585
R283 B.n222 B.n221 585
R284 B.n220 B.n208 585
R285 B.n219 B.n218 585
R286 B.n216 B.n209 585
R287 B.n214 B.n213 585
R288 B.n212 B.n211 585
R289 B.n162 B.n161 585
R290 B.n376 B.n375 585
R291 B.n377 B.n376 585
R292 B.n158 B.n157 585
R293 B.n159 B.n158 585
R294 B.n385 B.n384 585
R295 B.n384 B.n383 585
R296 B.n386 B.n156 585
R297 B.n156 B.n155 585
R298 B.n388 B.n387 585
R299 B.n389 B.n388 585
R300 B.n150 B.n149 585
R301 B.n151 B.n150 585
R302 B.n397 B.n396 585
R303 B.n396 B.n395 585
R304 B.n398 B.n148 585
R305 B.n148 B.n147 585
R306 B.n400 B.n399 585
R307 B.n401 B.n400 585
R308 B.n142 B.n141 585
R309 B.n143 B.n142 585
R310 B.n409 B.n408 585
R311 B.n408 B.n407 585
R312 B.n410 B.n140 585
R313 B.n140 B.n139 585
R314 B.n412 B.n411 585
R315 B.n413 B.n412 585
R316 B.n134 B.n133 585
R317 B.n135 B.n134 585
R318 B.n421 B.n420 585
R319 B.n420 B.n419 585
R320 B.n422 B.n132 585
R321 B.n132 B.n131 585
R322 B.n424 B.n423 585
R323 B.n425 B.n424 585
R324 B.n126 B.n125 585
R325 B.n127 B.n126 585
R326 B.n433 B.n432 585
R327 B.n432 B.n431 585
R328 B.n434 B.n124 585
R329 B.n124 B.n123 585
R330 B.n436 B.n435 585
R331 B.n437 B.n436 585
R332 B.n118 B.n117 585
R333 B.n119 B.n118 585
R334 B.n445 B.n444 585
R335 B.n444 B.n443 585
R336 B.n446 B.n116 585
R337 B.n116 B.n115 585
R338 B.n448 B.n447 585
R339 B.n449 B.n448 585
R340 B.n110 B.n109 585
R341 B.n111 B.n110 585
R342 B.n458 B.n457 585
R343 B.n457 B.n456 585
R344 B.n459 B.n108 585
R345 B.n108 B.n107 585
R346 B.n461 B.n460 585
R347 B.n462 B.n461 585
R348 B.n2 B.n0 585
R349 B.n4 B.n2 585
R350 B.n3 B.n1 585
R351 B.n729 B.n3 585
R352 B.n727 B.n726 585
R353 B.n728 B.n727 585
R354 B.n725 B.n9 585
R355 B.n9 B.n8 585
R356 B.n724 B.n723 585
R357 B.n723 B.n722 585
R358 B.n11 B.n10 585
R359 B.n721 B.n11 585
R360 B.n719 B.n718 585
R361 B.n720 B.n719 585
R362 B.n717 B.n16 585
R363 B.n16 B.n15 585
R364 B.n716 B.n715 585
R365 B.n715 B.n714 585
R366 B.n18 B.n17 585
R367 B.n713 B.n18 585
R368 B.n711 B.n710 585
R369 B.n712 B.n711 585
R370 B.n709 B.n23 585
R371 B.n23 B.n22 585
R372 B.n708 B.n707 585
R373 B.n707 B.n706 585
R374 B.n25 B.n24 585
R375 B.n705 B.n25 585
R376 B.n703 B.n702 585
R377 B.n704 B.n703 585
R378 B.n701 B.n30 585
R379 B.n30 B.n29 585
R380 B.n700 B.n699 585
R381 B.n699 B.n698 585
R382 B.n32 B.n31 585
R383 B.n697 B.n32 585
R384 B.n695 B.n694 585
R385 B.n696 B.n695 585
R386 B.n693 B.n37 585
R387 B.n37 B.n36 585
R388 B.n692 B.n691 585
R389 B.n691 B.n690 585
R390 B.n39 B.n38 585
R391 B.n689 B.n39 585
R392 B.n687 B.n686 585
R393 B.n688 B.n687 585
R394 B.n685 B.n44 585
R395 B.n44 B.n43 585
R396 B.n684 B.n683 585
R397 B.n683 B.n682 585
R398 B.n46 B.n45 585
R399 B.n681 B.n46 585
R400 B.n679 B.n678 585
R401 B.n680 B.n679 585
R402 B.n677 B.n51 585
R403 B.n51 B.n50 585
R404 B.n676 B.n675 585
R405 B.n675 B.n674 585
R406 B.n53 B.n52 585
R407 B.n673 B.n53 585
R408 B.n671 B.n670 585
R409 B.n672 B.n671 585
R410 B.n732 B.n731 585
R411 B.n731 B.n730 585
R412 B.n376 B.n164 511.721
R413 B.n671 B.n58 511.721
R414 B.n378 B.n162 511.721
R415 B.n104 B.n56 511.721
R416 B.n191 B.t2 283.348
R417 B.n183 B.t10 283.348
R418 B.n77 B.t13 283.348
R419 B.n83 B.t6 283.348
R420 B.n507 B.n57 256.663
R421 B.n509 B.n57 256.663
R422 B.n515 B.n57 256.663
R423 B.n517 B.n57 256.663
R424 B.n523 B.n57 256.663
R425 B.n525 B.n57 256.663
R426 B.n531 B.n57 256.663
R427 B.n533 B.n57 256.663
R428 B.n539 B.n57 256.663
R429 B.n541 B.n57 256.663
R430 B.n547 B.n57 256.663
R431 B.n549 B.n57 256.663
R432 B.n555 B.n57 256.663
R433 B.n557 B.n57 256.663
R434 B.n563 B.n57 256.663
R435 B.n565 B.n57 256.663
R436 B.n571 B.n57 256.663
R437 B.n86 B.n57 256.663
R438 B.n577 B.n57 256.663
R439 B.n583 B.n57 256.663
R440 B.n585 B.n57 256.663
R441 B.n591 B.n57 256.663
R442 B.n593 B.n57 256.663
R443 B.n600 B.n57 256.663
R444 B.n602 B.n57 256.663
R445 B.n608 B.n57 256.663
R446 B.n610 B.n57 256.663
R447 B.n616 B.n57 256.663
R448 B.n618 B.n57 256.663
R449 B.n624 B.n57 256.663
R450 B.n626 B.n57 256.663
R451 B.n632 B.n57 256.663
R452 B.n634 B.n57 256.663
R453 B.n640 B.n57 256.663
R454 B.n642 B.n57 256.663
R455 B.n648 B.n57 256.663
R456 B.n650 B.n57 256.663
R457 B.n656 B.n57 256.663
R458 B.n658 B.n57 256.663
R459 B.n664 B.n57 256.663
R460 B.n666 B.n57 256.663
R461 B.n371 B.n163 256.663
R462 B.n166 B.n163 256.663
R463 B.n364 B.n163 256.663
R464 B.n358 B.n163 256.663
R465 B.n356 B.n163 256.663
R466 B.n350 B.n163 256.663
R467 B.n348 B.n163 256.663
R468 B.n342 B.n163 256.663
R469 B.n340 B.n163 256.663
R470 B.n334 B.n163 256.663
R471 B.n332 B.n163 256.663
R472 B.n326 B.n163 256.663
R473 B.n324 B.n163 256.663
R474 B.n318 B.n163 256.663
R475 B.n316 B.n163 256.663
R476 B.n310 B.n163 256.663
R477 B.n308 B.n163 256.663
R478 B.n302 B.n163 256.663
R479 B.n186 B.n163 256.663
R480 B.n296 B.n163 256.663
R481 B.n290 B.n163 256.663
R482 B.n288 B.n163 256.663
R483 B.n281 B.n163 256.663
R484 B.n279 B.n163 256.663
R485 B.n273 B.n163 256.663
R486 B.n271 B.n163 256.663
R487 B.n265 B.n163 256.663
R488 B.n263 B.n163 256.663
R489 B.n257 B.n163 256.663
R490 B.n255 B.n163 256.663
R491 B.n249 B.n163 256.663
R492 B.n247 B.n163 256.663
R493 B.n241 B.n163 256.663
R494 B.n239 B.n163 256.663
R495 B.n233 B.n163 256.663
R496 B.n231 B.n163 256.663
R497 B.n225 B.n163 256.663
R498 B.n223 B.n163 256.663
R499 B.n217 B.n163 256.663
R500 B.n215 B.n163 256.663
R501 B.n210 B.n163 256.663
R502 B.n376 B.n158 163.367
R503 B.n384 B.n158 163.367
R504 B.n384 B.n156 163.367
R505 B.n388 B.n156 163.367
R506 B.n388 B.n150 163.367
R507 B.n396 B.n150 163.367
R508 B.n396 B.n148 163.367
R509 B.n400 B.n148 163.367
R510 B.n400 B.n142 163.367
R511 B.n408 B.n142 163.367
R512 B.n408 B.n140 163.367
R513 B.n412 B.n140 163.367
R514 B.n412 B.n134 163.367
R515 B.n420 B.n134 163.367
R516 B.n420 B.n132 163.367
R517 B.n424 B.n132 163.367
R518 B.n424 B.n126 163.367
R519 B.n432 B.n126 163.367
R520 B.n432 B.n124 163.367
R521 B.n436 B.n124 163.367
R522 B.n436 B.n118 163.367
R523 B.n444 B.n118 163.367
R524 B.n444 B.n116 163.367
R525 B.n448 B.n116 163.367
R526 B.n448 B.n110 163.367
R527 B.n457 B.n110 163.367
R528 B.n457 B.n108 163.367
R529 B.n461 B.n108 163.367
R530 B.n461 B.n2 163.367
R531 B.n731 B.n2 163.367
R532 B.n731 B.n3 163.367
R533 B.n727 B.n3 163.367
R534 B.n727 B.n9 163.367
R535 B.n723 B.n9 163.367
R536 B.n723 B.n11 163.367
R537 B.n719 B.n11 163.367
R538 B.n719 B.n16 163.367
R539 B.n715 B.n16 163.367
R540 B.n715 B.n18 163.367
R541 B.n711 B.n18 163.367
R542 B.n711 B.n23 163.367
R543 B.n707 B.n23 163.367
R544 B.n707 B.n25 163.367
R545 B.n703 B.n25 163.367
R546 B.n703 B.n30 163.367
R547 B.n699 B.n30 163.367
R548 B.n699 B.n32 163.367
R549 B.n695 B.n32 163.367
R550 B.n695 B.n37 163.367
R551 B.n691 B.n37 163.367
R552 B.n691 B.n39 163.367
R553 B.n687 B.n39 163.367
R554 B.n687 B.n44 163.367
R555 B.n683 B.n44 163.367
R556 B.n683 B.n46 163.367
R557 B.n679 B.n46 163.367
R558 B.n679 B.n51 163.367
R559 B.n675 B.n51 163.367
R560 B.n675 B.n53 163.367
R561 B.n671 B.n53 163.367
R562 B.n372 B.n370 163.367
R563 B.n370 B.n369 163.367
R564 B.n366 B.n365 163.367
R565 B.n363 B.n168 163.367
R566 B.n359 B.n357 163.367
R567 B.n355 B.n170 163.367
R568 B.n351 B.n349 163.367
R569 B.n347 B.n172 163.367
R570 B.n343 B.n341 163.367
R571 B.n339 B.n174 163.367
R572 B.n335 B.n333 163.367
R573 B.n331 B.n176 163.367
R574 B.n327 B.n325 163.367
R575 B.n323 B.n178 163.367
R576 B.n319 B.n317 163.367
R577 B.n315 B.n180 163.367
R578 B.n311 B.n309 163.367
R579 B.n307 B.n182 163.367
R580 B.n303 B.n301 163.367
R581 B.n298 B.n297 163.367
R582 B.n295 B.n188 163.367
R583 B.n291 B.n289 163.367
R584 B.n287 B.n190 163.367
R585 B.n282 B.n280 163.367
R586 B.n278 B.n194 163.367
R587 B.n274 B.n272 163.367
R588 B.n270 B.n196 163.367
R589 B.n266 B.n264 163.367
R590 B.n262 B.n198 163.367
R591 B.n258 B.n256 163.367
R592 B.n254 B.n200 163.367
R593 B.n250 B.n248 163.367
R594 B.n246 B.n202 163.367
R595 B.n242 B.n240 163.367
R596 B.n238 B.n204 163.367
R597 B.n234 B.n232 163.367
R598 B.n230 B.n206 163.367
R599 B.n226 B.n224 163.367
R600 B.n222 B.n208 163.367
R601 B.n218 B.n216 163.367
R602 B.n214 B.n211 163.367
R603 B.n378 B.n160 163.367
R604 B.n382 B.n160 163.367
R605 B.n382 B.n154 163.367
R606 B.n390 B.n154 163.367
R607 B.n390 B.n152 163.367
R608 B.n394 B.n152 163.367
R609 B.n394 B.n146 163.367
R610 B.n402 B.n146 163.367
R611 B.n402 B.n144 163.367
R612 B.n406 B.n144 163.367
R613 B.n406 B.n138 163.367
R614 B.n414 B.n138 163.367
R615 B.n414 B.n136 163.367
R616 B.n418 B.n136 163.367
R617 B.n418 B.n130 163.367
R618 B.n426 B.n130 163.367
R619 B.n426 B.n128 163.367
R620 B.n430 B.n128 163.367
R621 B.n430 B.n122 163.367
R622 B.n438 B.n122 163.367
R623 B.n438 B.n120 163.367
R624 B.n442 B.n120 163.367
R625 B.n442 B.n114 163.367
R626 B.n450 B.n114 163.367
R627 B.n450 B.n112 163.367
R628 B.n455 B.n112 163.367
R629 B.n455 B.n106 163.367
R630 B.n463 B.n106 163.367
R631 B.n464 B.n463 163.367
R632 B.n464 B.n5 163.367
R633 B.n6 B.n5 163.367
R634 B.n7 B.n6 163.367
R635 B.n469 B.n7 163.367
R636 B.n469 B.n12 163.367
R637 B.n13 B.n12 163.367
R638 B.n14 B.n13 163.367
R639 B.n474 B.n14 163.367
R640 B.n474 B.n19 163.367
R641 B.n20 B.n19 163.367
R642 B.n21 B.n20 163.367
R643 B.n479 B.n21 163.367
R644 B.n479 B.n26 163.367
R645 B.n27 B.n26 163.367
R646 B.n28 B.n27 163.367
R647 B.n484 B.n28 163.367
R648 B.n484 B.n33 163.367
R649 B.n34 B.n33 163.367
R650 B.n35 B.n34 163.367
R651 B.n489 B.n35 163.367
R652 B.n489 B.n40 163.367
R653 B.n41 B.n40 163.367
R654 B.n42 B.n41 163.367
R655 B.n494 B.n42 163.367
R656 B.n494 B.n47 163.367
R657 B.n48 B.n47 163.367
R658 B.n49 B.n48 163.367
R659 B.n499 B.n49 163.367
R660 B.n499 B.n54 163.367
R661 B.n55 B.n54 163.367
R662 B.n56 B.n55 163.367
R663 B.n667 B.n665 163.367
R664 B.n663 B.n60 163.367
R665 B.n659 B.n657 163.367
R666 B.n655 B.n62 163.367
R667 B.n651 B.n649 163.367
R668 B.n647 B.n64 163.367
R669 B.n643 B.n641 163.367
R670 B.n639 B.n66 163.367
R671 B.n635 B.n633 163.367
R672 B.n631 B.n68 163.367
R673 B.n627 B.n625 163.367
R674 B.n623 B.n70 163.367
R675 B.n619 B.n617 163.367
R676 B.n615 B.n72 163.367
R677 B.n611 B.n609 163.367
R678 B.n607 B.n74 163.367
R679 B.n603 B.n601 163.367
R680 B.n599 B.n76 163.367
R681 B.n594 B.n592 163.367
R682 B.n590 B.n80 163.367
R683 B.n586 B.n584 163.367
R684 B.n582 B.n82 163.367
R685 B.n578 B.n576 163.367
R686 B.n573 B.n572 163.367
R687 B.n570 B.n88 163.367
R688 B.n566 B.n564 163.367
R689 B.n562 B.n90 163.367
R690 B.n558 B.n556 163.367
R691 B.n554 B.n92 163.367
R692 B.n550 B.n548 163.367
R693 B.n546 B.n94 163.367
R694 B.n542 B.n540 163.367
R695 B.n538 B.n96 163.367
R696 B.n534 B.n532 163.367
R697 B.n530 B.n98 163.367
R698 B.n526 B.n524 163.367
R699 B.n522 B.n100 163.367
R700 B.n518 B.n516 163.367
R701 B.n514 B.n102 163.367
R702 B.n510 B.n508 163.367
R703 B.n506 B.n104 163.367
R704 B.n191 B.t5 143.678
R705 B.n83 B.t8 143.678
R706 B.n183 B.t12 143.665
R707 B.n77 B.t14 143.665
R708 B.n377 B.n163 80.7023
R709 B.n672 B.n57 80.7023
R710 B.n192 B.t4 71.92
R711 B.n84 B.t9 71.92
R712 B.n184 B.t11 71.9073
R713 B.n78 B.t15 71.9073
R714 B.n192 B.n191 71.7581
R715 B.n184 B.n183 71.7581
R716 B.n78 B.n77 71.7581
R717 B.n84 B.n83 71.7581
R718 B.n371 B.n164 71.676
R719 B.n369 B.n166 71.676
R720 B.n365 B.n364 71.676
R721 B.n358 B.n168 71.676
R722 B.n357 B.n356 71.676
R723 B.n350 B.n170 71.676
R724 B.n349 B.n348 71.676
R725 B.n342 B.n172 71.676
R726 B.n341 B.n340 71.676
R727 B.n334 B.n174 71.676
R728 B.n333 B.n332 71.676
R729 B.n326 B.n176 71.676
R730 B.n325 B.n324 71.676
R731 B.n318 B.n178 71.676
R732 B.n317 B.n316 71.676
R733 B.n310 B.n180 71.676
R734 B.n309 B.n308 71.676
R735 B.n302 B.n182 71.676
R736 B.n301 B.n186 71.676
R737 B.n297 B.n296 71.676
R738 B.n290 B.n188 71.676
R739 B.n289 B.n288 71.676
R740 B.n281 B.n190 71.676
R741 B.n280 B.n279 71.676
R742 B.n273 B.n194 71.676
R743 B.n272 B.n271 71.676
R744 B.n265 B.n196 71.676
R745 B.n264 B.n263 71.676
R746 B.n257 B.n198 71.676
R747 B.n256 B.n255 71.676
R748 B.n249 B.n200 71.676
R749 B.n248 B.n247 71.676
R750 B.n241 B.n202 71.676
R751 B.n240 B.n239 71.676
R752 B.n233 B.n204 71.676
R753 B.n232 B.n231 71.676
R754 B.n225 B.n206 71.676
R755 B.n224 B.n223 71.676
R756 B.n217 B.n208 71.676
R757 B.n216 B.n215 71.676
R758 B.n211 B.n210 71.676
R759 B.n666 B.n58 71.676
R760 B.n665 B.n664 71.676
R761 B.n658 B.n60 71.676
R762 B.n657 B.n656 71.676
R763 B.n650 B.n62 71.676
R764 B.n649 B.n648 71.676
R765 B.n642 B.n64 71.676
R766 B.n641 B.n640 71.676
R767 B.n634 B.n66 71.676
R768 B.n633 B.n632 71.676
R769 B.n626 B.n68 71.676
R770 B.n625 B.n624 71.676
R771 B.n618 B.n70 71.676
R772 B.n617 B.n616 71.676
R773 B.n610 B.n72 71.676
R774 B.n609 B.n608 71.676
R775 B.n602 B.n74 71.676
R776 B.n601 B.n600 71.676
R777 B.n593 B.n76 71.676
R778 B.n592 B.n591 71.676
R779 B.n585 B.n80 71.676
R780 B.n584 B.n583 71.676
R781 B.n577 B.n82 71.676
R782 B.n576 B.n86 71.676
R783 B.n572 B.n571 71.676
R784 B.n565 B.n88 71.676
R785 B.n564 B.n563 71.676
R786 B.n557 B.n90 71.676
R787 B.n556 B.n555 71.676
R788 B.n549 B.n92 71.676
R789 B.n548 B.n547 71.676
R790 B.n541 B.n94 71.676
R791 B.n540 B.n539 71.676
R792 B.n533 B.n96 71.676
R793 B.n532 B.n531 71.676
R794 B.n525 B.n98 71.676
R795 B.n524 B.n523 71.676
R796 B.n517 B.n100 71.676
R797 B.n516 B.n515 71.676
R798 B.n509 B.n102 71.676
R799 B.n508 B.n507 71.676
R800 B.n507 B.n506 71.676
R801 B.n510 B.n509 71.676
R802 B.n515 B.n514 71.676
R803 B.n518 B.n517 71.676
R804 B.n523 B.n522 71.676
R805 B.n526 B.n525 71.676
R806 B.n531 B.n530 71.676
R807 B.n534 B.n533 71.676
R808 B.n539 B.n538 71.676
R809 B.n542 B.n541 71.676
R810 B.n547 B.n546 71.676
R811 B.n550 B.n549 71.676
R812 B.n555 B.n554 71.676
R813 B.n558 B.n557 71.676
R814 B.n563 B.n562 71.676
R815 B.n566 B.n565 71.676
R816 B.n571 B.n570 71.676
R817 B.n573 B.n86 71.676
R818 B.n578 B.n577 71.676
R819 B.n583 B.n582 71.676
R820 B.n586 B.n585 71.676
R821 B.n591 B.n590 71.676
R822 B.n594 B.n593 71.676
R823 B.n600 B.n599 71.676
R824 B.n603 B.n602 71.676
R825 B.n608 B.n607 71.676
R826 B.n611 B.n610 71.676
R827 B.n616 B.n615 71.676
R828 B.n619 B.n618 71.676
R829 B.n624 B.n623 71.676
R830 B.n627 B.n626 71.676
R831 B.n632 B.n631 71.676
R832 B.n635 B.n634 71.676
R833 B.n640 B.n639 71.676
R834 B.n643 B.n642 71.676
R835 B.n648 B.n647 71.676
R836 B.n651 B.n650 71.676
R837 B.n656 B.n655 71.676
R838 B.n659 B.n658 71.676
R839 B.n664 B.n663 71.676
R840 B.n667 B.n666 71.676
R841 B.n372 B.n371 71.676
R842 B.n366 B.n166 71.676
R843 B.n364 B.n363 71.676
R844 B.n359 B.n358 71.676
R845 B.n356 B.n355 71.676
R846 B.n351 B.n350 71.676
R847 B.n348 B.n347 71.676
R848 B.n343 B.n342 71.676
R849 B.n340 B.n339 71.676
R850 B.n335 B.n334 71.676
R851 B.n332 B.n331 71.676
R852 B.n327 B.n326 71.676
R853 B.n324 B.n323 71.676
R854 B.n319 B.n318 71.676
R855 B.n316 B.n315 71.676
R856 B.n311 B.n310 71.676
R857 B.n308 B.n307 71.676
R858 B.n303 B.n302 71.676
R859 B.n298 B.n186 71.676
R860 B.n296 B.n295 71.676
R861 B.n291 B.n290 71.676
R862 B.n288 B.n287 71.676
R863 B.n282 B.n281 71.676
R864 B.n279 B.n278 71.676
R865 B.n274 B.n273 71.676
R866 B.n271 B.n270 71.676
R867 B.n266 B.n265 71.676
R868 B.n263 B.n262 71.676
R869 B.n258 B.n257 71.676
R870 B.n255 B.n254 71.676
R871 B.n250 B.n249 71.676
R872 B.n247 B.n246 71.676
R873 B.n242 B.n241 71.676
R874 B.n239 B.n238 71.676
R875 B.n234 B.n233 71.676
R876 B.n231 B.n230 71.676
R877 B.n226 B.n225 71.676
R878 B.n223 B.n222 71.676
R879 B.n218 B.n217 71.676
R880 B.n215 B.n214 71.676
R881 B.n210 B.n162 71.676
R882 B.n284 B.n192 59.5399
R883 B.n185 B.n184 59.5399
R884 B.n596 B.n78 59.5399
R885 B.n85 B.n84 59.5399
R886 B.n377 B.n159 47.7198
R887 B.n383 B.n159 47.7198
R888 B.n383 B.n155 47.7198
R889 B.n389 B.n155 47.7198
R890 B.n389 B.n151 47.7198
R891 B.n395 B.n151 47.7198
R892 B.n395 B.n147 47.7198
R893 B.n401 B.n147 47.7198
R894 B.n407 B.n143 47.7198
R895 B.n407 B.n139 47.7198
R896 B.n413 B.n139 47.7198
R897 B.n413 B.n135 47.7198
R898 B.n419 B.n135 47.7198
R899 B.n419 B.n131 47.7198
R900 B.n425 B.n131 47.7198
R901 B.n425 B.n127 47.7198
R902 B.n431 B.n127 47.7198
R903 B.n431 B.n123 47.7198
R904 B.n437 B.n123 47.7198
R905 B.n437 B.n119 47.7198
R906 B.n443 B.n119 47.7198
R907 B.n449 B.n115 47.7198
R908 B.n449 B.n111 47.7198
R909 B.n456 B.n111 47.7198
R910 B.n456 B.n107 47.7198
R911 B.n462 B.n107 47.7198
R912 B.n462 B.n4 47.7198
R913 B.n730 B.n4 47.7198
R914 B.n730 B.n729 47.7198
R915 B.n729 B.n728 47.7198
R916 B.n728 B.n8 47.7198
R917 B.n722 B.n8 47.7198
R918 B.n722 B.n721 47.7198
R919 B.n721 B.n720 47.7198
R920 B.n720 B.n15 47.7198
R921 B.n714 B.n713 47.7198
R922 B.n713 B.n712 47.7198
R923 B.n712 B.n22 47.7198
R924 B.n706 B.n22 47.7198
R925 B.n706 B.n705 47.7198
R926 B.n705 B.n704 47.7198
R927 B.n704 B.n29 47.7198
R928 B.n698 B.n29 47.7198
R929 B.n698 B.n697 47.7198
R930 B.n697 B.n696 47.7198
R931 B.n696 B.n36 47.7198
R932 B.n690 B.n36 47.7198
R933 B.n690 B.n689 47.7198
R934 B.n688 B.n43 47.7198
R935 B.n682 B.n43 47.7198
R936 B.n682 B.n681 47.7198
R937 B.n681 B.n680 47.7198
R938 B.n680 B.n50 47.7198
R939 B.n674 B.n50 47.7198
R940 B.n674 B.n673 47.7198
R941 B.n673 B.n672 47.7198
R942 B.n443 B.t0 45.6145
R943 B.n714 B.t1 45.6145
R944 B.n401 B.t3 41.404
R945 B.t7 B.n688 41.404
R946 B.n670 B.n669 33.2493
R947 B.n504 B.n503 33.2493
R948 B.n379 B.n161 33.2493
R949 B.n375 B.n374 33.2493
R950 B B.n732 18.0485
R951 B.n669 B.n668 10.6151
R952 B.n668 B.n59 10.6151
R953 B.n662 B.n59 10.6151
R954 B.n662 B.n661 10.6151
R955 B.n661 B.n660 10.6151
R956 B.n660 B.n61 10.6151
R957 B.n654 B.n61 10.6151
R958 B.n654 B.n653 10.6151
R959 B.n653 B.n652 10.6151
R960 B.n652 B.n63 10.6151
R961 B.n646 B.n63 10.6151
R962 B.n646 B.n645 10.6151
R963 B.n645 B.n644 10.6151
R964 B.n644 B.n65 10.6151
R965 B.n638 B.n65 10.6151
R966 B.n638 B.n637 10.6151
R967 B.n637 B.n636 10.6151
R968 B.n636 B.n67 10.6151
R969 B.n630 B.n67 10.6151
R970 B.n630 B.n629 10.6151
R971 B.n629 B.n628 10.6151
R972 B.n628 B.n69 10.6151
R973 B.n622 B.n69 10.6151
R974 B.n622 B.n621 10.6151
R975 B.n621 B.n620 10.6151
R976 B.n620 B.n71 10.6151
R977 B.n614 B.n71 10.6151
R978 B.n614 B.n613 10.6151
R979 B.n613 B.n612 10.6151
R980 B.n612 B.n73 10.6151
R981 B.n606 B.n73 10.6151
R982 B.n606 B.n605 10.6151
R983 B.n605 B.n604 10.6151
R984 B.n604 B.n75 10.6151
R985 B.n598 B.n75 10.6151
R986 B.n598 B.n597 10.6151
R987 B.n595 B.n79 10.6151
R988 B.n589 B.n79 10.6151
R989 B.n589 B.n588 10.6151
R990 B.n588 B.n587 10.6151
R991 B.n587 B.n81 10.6151
R992 B.n581 B.n81 10.6151
R993 B.n581 B.n580 10.6151
R994 B.n580 B.n579 10.6151
R995 B.n575 B.n574 10.6151
R996 B.n574 B.n87 10.6151
R997 B.n569 B.n87 10.6151
R998 B.n569 B.n568 10.6151
R999 B.n568 B.n567 10.6151
R1000 B.n567 B.n89 10.6151
R1001 B.n561 B.n89 10.6151
R1002 B.n561 B.n560 10.6151
R1003 B.n560 B.n559 10.6151
R1004 B.n559 B.n91 10.6151
R1005 B.n553 B.n91 10.6151
R1006 B.n553 B.n552 10.6151
R1007 B.n552 B.n551 10.6151
R1008 B.n551 B.n93 10.6151
R1009 B.n545 B.n93 10.6151
R1010 B.n545 B.n544 10.6151
R1011 B.n544 B.n543 10.6151
R1012 B.n543 B.n95 10.6151
R1013 B.n537 B.n95 10.6151
R1014 B.n537 B.n536 10.6151
R1015 B.n536 B.n535 10.6151
R1016 B.n535 B.n97 10.6151
R1017 B.n529 B.n97 10.6151
R1018 B.n529 B.n528 10.6151
R1019 B.n528 B.n527 10.6151
R1020 B.n527 B.n99 10.6151
R1021 B.n521 B.n99 10.6151
R1022 B.n521 B.n520 10.6151
R1023 B.n520 B.n519 10.6151
R1024 B.n519 B.n101 10.6151
R1025 B.n513 B.n101 10.6151
R1026 B.n513 B.n512 10.6151
R1027 B.n512 B.n511 10.6151
R1028 B.n511 B.n103 10.6151
R1029 B.n505 B.n103 10.6151
R1030 B.n505 B.n504 10.6151
R1031 B.n380 B.n379 10.6151
R1032 B.n381 B.n380 10.6151
R1033 B.n381 B.n153 10.6151
R1034 B.n391 B.n153 10.6151
R1035 B.n392 B.n391 10.6151
R1036 B.n393 B.n392 10.6151
R1037 B.n393 B.n145 10.6151
R1038 B.n403 B.n145 10.6151
R1039 B.n404 B.n403 10.6151
R1040 B.n405 B.n404 10.6151
R1041 B.n405 B.n137 10.6151
R1042 B.n415 B.n137 10.6151
R1043 B.n416 B.n415 10.6151
R1044 B.n417 B.n416 10.6151
R1045 B.n417 B.n129 10.6151
R1046 B.n427 B.n129 10.6151
R1047 B.n428 B.n427 10.6151
R1048 B.n429 B.n428 10.6151
R1049 B.n429 B.n121 10.6151
R1050 B.n439 B.n121 10.6151
R1051 B.n440 B.n439 10.6151
R1052 B.n441 B.n440 10.6151
R1053 B.n441 B.n113 10.6151
R1054 B.n451 B.n113 10.6151
R1055 B.n452 B.n451 10.6151
R1056 B.n454 B.n452 10.6151
R1057 B.n454 B.n453 10.6151
R1058 B.n453 B.n105 10.6151
R1059 B.n465 B.n105 10.6151
R1060 B.n466 B.n465 10.6151
R1061 B.n467 B.n466 10.6151
R1062 B.n468 B.n467 10.6151
R1063 B.n470 B.n468 10.6151
R1064 B.n471 B.n470 10.6151
R1065 B.n472 B.n471 10.6151
R1066 B.n473 B.n472 10.6151
R1067 B.n475 B.n473 10.6151
R1068 B.n476 B.n475 10.6151
R1069 B.n477 B.n476 10.6151
R1070 B.n478 B.n477 10.6151
R1071 B.n480 B.n478 10.6151
R1072 B.n481 B.n480 10.6151
R1073 B.n482 B.n481 10.6151
R1074 B.n483 B.n482 10.6151
R1075 B.n485 B.n483 10.6151
R1076 B.n486 B.n485 10.6151
R1077 B.n487 B.n486 10.6151
R1078 B.n488 B.n487 10.6151
R1079 B.n490 B.n488 10.6151
R1080 B.n491 B.n490 10.6151
R1081 B.n492 B.n491 10.6151
R1082 B.n493 B.n492 10.6151
R1083 B.n495 B.n493 10.6151
R1084 B.n496 B.n495 10.6151
R1085 B.n497 B.n496 10.6151
R1086 B.n498 B.n497 10.6151
R1087 B.n500 B.n498 10.6151
R1088 B.n501 B.n500 10.6151
R1089 B.n502 B.n501 10.6151
R1090 B.n503 B.n502 10.6151
R1091 B.n374 B.n373 10.6151
R1092 B.n373 B.n165 10.6151
R1093 B.n368 B.n165 10.6151
R1094 B.n368 B.n367 10.6151
R1095 B.n367 B.n167 10.6151
R1096 B.n362 B.n167 10.6151
R1097 B.n362 B.n361 10.6151
R1098 B.n361 B.n360 10.6151
R1099 B.n360 B.n169 10.6151
R1100 B.n354 B.n169 10.6151
R1101 B.n354 B.n353 10.6151
R1102 B.n353 B.n352 10.6151
R1103 B.n352 B.n171 10.6151
R1104 B.n346 B.n171 10.6151
R1105 B.n346 B.n345 10.6151
R1106 B.n345 B.n344 10.6151
R1107 B.n344 B.n173 10.6151
R1108 B.n338 B.n173 10.6151
R1109 B.n338 B.n337 10.6151
R1110 B.n337 B.n336 10.6151
R1111 B.n336 B.n175 10.6151
R1112 B.n330 B.n175 10.6151
R1113 B.n330 B.n329 10.6151
R1114 B.n329 B.n328 10.6151
R1115 B.n328 B.n177 10.6151
R1116 B.n322 B.n177 10.6151
R1117 B.n322 B.n321 10.6151
R1118 B.n321 B.n320 10.6151
R1119 B.n320 B.n179 10.6151
R1120 B.n314 B.n179 10.6151
R1121 B.n314 B.n313 10.6151
R1122 B.n313 B.n312 10.6151
R1123 B.n312 B.n181 10.6151
R1124 B.n306 B.n181 10.6151
R1125 B.n306 B.n305 10.6151
R1126 B.n305 B.n304 10.6151
R1127 B.n300 B.n299 10.6151
R1128 B.n299 B.n187 10.6151
R1129 B.n294 B.n187 10.6151
R1130 B.n294 B.n293 10.6151
R1131 B.n293 B.n292 10.6151
R1132 B.n292 B.n189 10.6151
R1133 B.n286 B.n189 10.6151
R1134 B.n286 B.n285 10.6151
R1135 B.n283 B.n193 10.6151
R1136 B.n277 B.n193 10.6151
R1137 B.n277 B.n276 10.6151
R1138 B.n276 B.n275 10.6151
R1139 B.n275 B.n195 10.6151
R1140 B.n269 B.n195 10.6151
R1141 B.n269 B.n268 10.6151
R1142 B.n268 B.n267 10.6151
R1143 B.n267 B.n197 10.6151
R1144 B.n261 B.n197 10.6151
R1145 B.n261 B.n260 10.6151
R1146 B.n260 B.n259 10.6151
R1147 B.n259 B.n199 10.6151
R1148 B.n253 B.n199 10.6151
R1149 B.n253 B.n252 10.6151
R1150 B.n252 B.n251 10.6151
R1151 B.n251 B.n201 10.6151
R1152 B.n245 B.n201 10.6151
R1153 B.n245 B.n244 10.6151
R1154 B.n244 B.n243 10.6151
R1155 B.n243 B.n203 10.6151
R1156 B.n237 B.n203 10.6151
R1157 B.n237 B.n236 10.6151
R1158 B.n236 B.n235 10.6151
R1159 B.n235 B.n205 10.6151
R1160 B.n229 B.n205 10.6151
R1161 B.n229 B.n228 10.6151
R1162 B.n228 B.n227 10.6151
R1163 B.n227 B.n207 10.6151
R1164 B.n221 B.n207 10.6151
R1165 B.n221 B.n220 10.6151
R1166 B.n220 B.n219 10.6151
R1167 B.n219 B.n209 10.6151
R1168 B.n213 B.n209 10.6151
R1169 B.n213 B.n212 10.6151
R1170 B.n212 B.n161 10.6151
R1171 B.n375 B.n157 10.6151
R1172 B.n385 B.n157 10.6151
R1173 B.n386 B.n385 10.6151
R1174 B.n387 B.n386 10.6151
R1175 B.n387 B.n149 10.6151
R1176 B.n397 B.n149 10.6151
R1177 B.n398 B.n397 10.6151
R1178 B.n399 B.n398 10.6151
R1179 B.n399 B.n141 10.6151
R1180 B.n409 B.n141 10.6151
R1181 B.n410 B.n409 10.6151
R1182 B.n411 B.n410 10.6151
R1183 B.n411 B.n133 10.6151
R1184 B.n421 B.n133 10.6151
R1185 B.n422 B.n421 10.6151
R1186 B.n423 B.n422 10.6151
R1187 B.n423 B.n125 10.6151
R1188 B.n433 B.n125 10.6151
R1189 B.n434 B.n433 10.6151
R1190 B.n435 B.n434 10.6151
R1191 B.n435 B.n117 10.6151
R1192 B.n445 B.n117 10.6151
R1193 B.n446 B.n445 10.6151
R1194 B.n447 B.n446 10.6151
R1195 B.n447 B.n109 10.6151
R1196 B.n458 B.n109 10.6151
R1197 B.n459 B.n458 10.6151
R1198 B.n460 B.n459 10.6151
R1199 B.n460 B.n0 10.6151
R1200 B.n726 B.n1 10.6151
R1201 B.n726 B.n725 10.6151
R1202 B.n725 B.n724 10.6151
R1203 B.n724 B.n10 10.6151
R1204 B.n718 B.n10 10.6151
R1205 B.n718 B.n717 10.6151
R1206 B.n717 B.n716 10.6151
R1207 B.n716 B.n17 10.6151
R1208 B.n710 B.n17 10.6151
R1209 B.n710 B.n709 10.6151
R1210 B.n709 B.n708 10.6151
R1211 B.n708 B.n24 10.6151
R1212 B.n702 B.n24 10.6151
R1213 B.n702 B.n701 10.6151
R1214 B.n701 B.n700 10.6151
R1215 B.n700 B.n31 10.6151
R1216 B.n694 B.n31 10.6151
R1217 B.n694 B.n693 10.6151
R1218 B.n693 B.n692 10.6151
R1219 B.n692 B.n38 10.6151
R1220 B.n686 B.n38 10.6151
R1221 B.n686 B.n685 10.6151
R1222 B.n685 B.n684 10.6151
R1223 B.n684 B.n45 10.6151
R1224 B.n678 B.n45 10.6151
R1225 B.n678 B.n677 10.6151
R1226 B.n677 B.n676 10.6151
R1227 B.n676 B.n52 10.6151
R1228 B.n670 B.n52 10.6151
R1229 B.n596 B.n595 6.5566
R1230 B.n579 B.n85 6.5566
R1231 B.n300 B.n185 6.5566
R1232 B.n285 B.n284 6.5566
R1233 B.t3 B.n143 6.31629
R1234 B.n689 B.t7 6.31629
R1235 B.n597 B.n596 4.05904
R1236 B.n575 B.n85 4.05904
R1237 B.n304 B.n185 4.05904
R1238 B.n284 B.n283 4.05904
R1239 B.n732 B.n0 2.81026
R1240 B.n732 B.n1 2.81026
R1241 B.t0 B.n115 2.10576
R1242 B.t1 B.n15 2.10576
R1243 VP.n0 VP.t1 158.59
R1244 VP.n0 VP.t0 113.105
R1245 VP VP.n0 0.526368
R1246 VTAIL.n1 VTAIL.t1 49.2596
R1247 VTAIL.n2 VTAIL.t2 49.2593
R1248 VTAIL.n3 VTAIL.t0 49.2593
R1249 VTAIL.n0 VTAIL.t3 49.2593
R1250 VTAIL.n1 VTAIL.n0 27.7117
R1251 VTAIL.n3 VTAIL.n2 24.5221
R1252 VTAIL.n2 VTAIL.n1 2.06516
R1253 VTAIL VTAIL.n0 1.32593
R1254 VTAIL VTAIL.n3 0.739724
R1255 VDD1 VDD1.t1 106.264
R1256 VDD1 VDD1.t0 66.7937
R1257 VN VN.t1 158.499
R1258 VN VN.t0 113.63
R1259 VDD2.n0 VDD2.t1 104.942
R1260 VDD2.n0 VDD2.t0 65.9381
R1261 VDD2 VDD2.n0 0.856103
C0 VN VTAIL 2.32121f
C1 VP VDD1 2.74505f
C2 VDD2 VTAIL 4.86194f
C3 VN VDD1 0.148141f
C4 VDD2 VDD1 0.768418f
C5 VP VN 5.52503f
C6 VTAIL VDD1 4.8052f
C7 VP VDD2 0.364978f
C8 VN VDD2 2.53021f
C9 VP VTAIL 2.33543f
C10 VDD2 B 4.41336f
C11 VDD1 B 7.5758f
C12 VTAIL B 7.076122f
C13 VN B 11.09327f
C14 VP B 7.2501f
C15 VDD2.t1 B 2.43752f
C16 VDD2.t0 B 1.9039f
C17 VDD2.n0 B 2.89553f
C18 VN.t0 B 2.93204f
C19 VN.t1 B 3.55687f
C20 VDD1.t0 B 1.91366f
C21 VDD1.t1 B 2.48567f
C22 VTAIL.t3 B 1.91249f
C23 VTAIL.n0 B 1.72177f
C24 VTAIL.t1 B 1.91249f
C25 VTAIL.n1 B 1.77295f
C26 VTAIL.t2 B 1.91249f
C27 VTAIL.n2 B 1.55207f
C28 VTAIL.t0 B 1.91249f
C29 VTAIL.n3 B 1.46028f
C30 VP.t1 B 3.63912f
C31 VP.t0 B 2.99562f
C32 VP.n0 B 3.76697f
.ends

