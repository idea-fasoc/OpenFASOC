* NGSPICE file created from diff_pair_sample_1697.ext - technology: sky130A

.subckt diff_pair_sample_1697 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t16 w_n6022_n4064# sky130_fd_pr__pfet_01v8 ad=6.0372 pd=31.74 as=2.5542 ps=15.81 w=15.48 l=3.88
X1 VDD2.t9 VN.t0 VTAIL.t1 w_n6022_n4064# sky130_fd_pr__pfet_01v8 ad=2.5542 pd=15.81 as=2.5542 ps=15.81 w=15.48 l=3.88
X2 B.t11 B.t9 B.t10 w_n6022_n4064# sky130_fd_pr__pfet_01v8 ad=6.0372 pd=31.74 as=0 ps=0 w=15.48 l=3.88
X3 VDD1.t8 VP.t1 VTAIL.t8 w_n6022_n4064# sky130_fd_pr__pfet_01v8 ad=2.5542 pd=15.81 as=6.0372 ps=31.74 w=15.48 l=3.88
X4 VTAIL.t9 VP.t2 VDD1.t7 w_n6022_n4064# sky130_fd_pr__pfet_01v8 ad=2.5542 pd=15.81 as=2.5542 ps=15.81 w=15.48 l=3.88
X5 VDD2.t8 VN.t1 VTAIL.t0 w_n6022_n4064# sky130_fd_pr__pfet_01v8 ad=2.5542 pd=15.81 as=6.0372 ps=31.74 w=15.48 l=3.88
X6 VDD2.t7 VN.t2 VTAIL.t7 w_n6022_n4064# sky130_fd_pr__pfet_01v8 ad=6.0372 pd=31.74 as=2.5542 ps=15.81 w=15.48 l=3.88
X7 VTAIL.t6 VN.t3 VDD2.t6 w_n6022_n4064# sky130_fd_pr__pfet_01v8 ad=2.5542 pd=15.81 as=2.5542 ps=15.81 w=15.48 l=3.88
X8 VTAIL.t10 VP.t3 VDD1.t6 w_n6022_n4064# sky130_fd_pr__pfet_01v8 ad=2.5542 pd=15.81 as=2.5542 ps=15.81 w=15.48 l=3.88
X9 B.t8 B.t6 B.t7 w_n6022_n4064# sky130_fd_pr__pfet_01v8 ad=6.0372 pd=31.74 as=0 ps=0 w=15.48 l=3.88
X10 VTAIL.t5 VN.t4 VDD2.t5 w_n6022_n4064# sky130_fd_pr__pfet_01v8 ad=2.5542 pd=15.81 as=2.5542 ps=15.81 w=15.48 l=3.88
X11 VTAIL.t18 VN.t5 VDD2.t4 w_n6022_n4064# sky130_fd_pr__pfet_01v8 ad=2.5542 pd=15.81 as=2.5542 ps=15.81 w=15.48 l=3.88
X12 VDD2.t3 VN.t6 VTAIL.t19 w_n6022_n4064# sky130_fd_pr__pfet_01v8 ad=2.5542 pd=15.81 as=6.0372 ps=31.74 w=15.48 l=3.88
X13 B.t5 B.t3 B.t4 w_n6022_n4064# sky130_fd_pr__pfet_01v8 ad=6.0372 pd=31.74 as=0 ps=0 w=15.48 l=3.88
X14 VDD1.t5 VP.t4 VTAIL.t14 w_n6022_n4064# sky130_fd_pr__pfet_01v8 ad=2.5542 pd=15.81 as=2.5542 ps=15.81 w=15.48 l=3.88
X15 B.t2 B.t0 B.t1 w_n6022_n4064# sky130_fd_pr__pfet_01v8 ad=6.0372 pd=31.74 as=0 ps=0 w=15.48 l=3.88
X16 VTAIL.t11 VP.t5 VDD1.t4 w_n6022_n4064# sky130_fd_pr__pfet_01v8 ad=2.5542 pd=15.81 as=2.5542 ps=15.81 w=15.48 l=3.88
X17 VTAIL.t4 VN.t7 VDD2.t2 w_n6022_n4064# sky130_fd_pr__pfet_01v8 ad=2.5542 pd=15.81 as=2.5542 ps=15.81 w=15.48 l=3.88
X18 VDD2.t1 VN.t8 VTAIL.t3 w_n6022_n4064# sky130_fd_pr__pfet_01v8 ad=2.5542 pd=15.81 as=2.5542 ps=15.81 w=15.48 l=3.88
X19 VDD2.t0 VN.t9 VTAIL.t2 w_n6022_n4064# sky130_fd_pr__pfet_01v8 ad=6.0372 pd=31.74 as=2.5542 ps=15.81 w=15.48 l=3.88
X20 VDD1.t3 VP.t6 VTAIL.t15 w_n6022_n4064# sky130_fd_pr__pfet_01v8 ad=6.0372 pd=31.74 as=2.5542 ps=15.81 w=15.48 l=3.88
X21 VDD1.t2 VP.t7 VTAIL.t17 w_n6022_n4064# sky130_fd_pr__pfet_01v8 ad=2.5542 pd=15.81 as=2.5542 ps=15.81 w=15.48 l=3.88
X22 VTAIL.t13 VP.t8 VDD1.t1 w_n6022_n4064# sky130_fd_pr__pfet_01v8 ad=2.5542 pd=15.81 as=2.5542 ps=15.81 w=15.48 l=3.88
X23 VDD1.t0 VP.t9 VTAIL.t12 w_n6022_n4064# sky130_fd_pr__pfet_01v8 ad=2.5542 pd=15.81 as=6.0372 ps=31.74 w=15.48 l=3.88
R0 VP.n32 VP.n29 161.3
R1 VP.n34 VP.n33 161.3
R2 VP.n35 VP.n28 161.3
R3 VP.n37 VP.n36 161.3
R4 VP.n38 VP.n27 161.3
R5 VP.n40 VP.n39 161.3
R6 VP.n41 VP.n26 161.3
R7 VP.n43 VP.n42 161.3
R8 VP.n44 VP.n25 161.3
R9 VP.n46 VP.n45 161.3
R10 VP.n47 VP.n24 161.3
R11 VP.n49 VP.n48 161.3
R12 VP.n50 VP.n23 161.3
R13 VP.n52 VP.n51 161.3
R14 VP.n53 VP.n22 161.3
R15 VP.n55 VP.n54 161.3
R16 VP.n56 VP.n21 161.3
R17 VP.n59 VP.n58 161.3
R18 VP.n60 VP.n20 161.3
R19 VP.n62 VP.n61 161.3
R20 VP.n63 VP.n19 161.3
R21 VP.n65 VP.n64 161.3
R22 VP.n66 VP.n18 161.3
R23 VP.n68 VP.n67 161.3
R24 VP.n69 VP.n17 161.3
R25 VP.n124 VP.n0 161.3
R26 VP.n123 VP.n122 161.3
R27 VP.n121 VP.n1 161.3
R28 VP.n120 VP.n119 161.3
R29 VP.n118 VP.n2 161.3
R30 VP.n117 VP.n116 161.3
R31 VP.n115 VP.n3 161.3
R32 VP.n114 VP.n113 161.3
R33 VP.n111 VP.n4 161.3
R34 VP.n110 VP.n109 161.3
R35 VP.n108 VP.n5 161.3
R36 VP.n107 VP.n106 161.3
R37 VP.n105 VP.n6 161.3
R38 VP.n104 VP.n103 161.3
R39 VP.n102 VP.n7 161.3
R40 VP.n101 VP.n100 161.3
R41 VP.n99 VP.n8 161.3
R42 VP.n98 VP.n97 161.3
R43 VP.n96 VP.n9 161.3
R44 VP.n95 VP.n94 161.3
R45 VP.n93 VP.n10 161.3
R46 VP.n92 VP.n91 161.3
R47 VP.n90 VP.n11 161.3
R48 VP.n89 VP.n88 161.3
R49 VP.n87 VP.n12 161.3
R50 VP.n85 VP.n84 161.3
R51 VP.n83 VP.n13 161.3
R52 VP.n82 VP.n81 161.3
R53 VP.n80 VP.n14 161.3
R54 VP.n79 VP.n78 161.3
R55 VP.n77 VP.n15 161.3
R56 VP.n76 VP.n75 161.3
R57 VP.n74 VP.n16 161.3
R58 VP.n30 VP.t6 128.481
R59 VP.n99 VP.t7 96.1521
R60 VP.n73 VP.t0 96.1521
R61 VP.n86 VP.t3 96.1521
R62 VP.n112 VP.t8 96.1521
R63 VP.n125 VP.t1 96.1521
R64 VP.n44 VP.t4 96.1521
R65 VP.n70 VP.t9 96.1521
R66 VP.n57 VP.t2 96.1521
R67 VP.n31 VP.t5 96.1521
R68 VP.n31 VP.n30 64.9805
R69 VP.n72 VP.n71 62.9325
R70 VP.n73 VP.n72 61.7228
R71 VP.n126 VP.n125 61.7228
R72 VP.n71 VP.n70 61.7228
R73 VP.n80 VP.n79 56.5617
R74 VP.n119 VP.n118 56.5617
R75 VP.n64 VP.n63 56.5617
R76 VP.n93 VP.n92 50.7491
R77 VP.n106 VP.n105 50.7491
R78 VP.n51 VP.n50 50.7491
R79 VP.n38 VP.n37 50.7491
R80 VP.n94 VP.n93 30.405
R81 VP.n105 VP.n104 30.405
R82 VP.n50 VP.n49 30.405
R83 VP.n39 VP.n38 30.405
R84 VP.n75 VP.n74 24.5923
R85 VP.n75 VP.n15 24.5923
R86 VP.n79 VP.n15 24.5923
R87 VP.n81 VP.n80 24.5923
R88 VP.n81 VP.n13 24.5923
R89 VP.n85 VP.n13 24.5923
R90 VP.n88 VP.n87 24.5923
R91 VP.n88 VP.n11 24.5923
R92 VP.n92 VP.n11 24.5923
R93 VP.n94 VP.n9 24.5923
R94 VP.n98 VP.n9 24.5923
R95 VP.n99 VP.n98 24.5923
R96 VP.n100 VP.n99 24.5923
R97 VP.n100 VP.n7 24.5923
R98 VP.n104 VP.n7 24.5923
R99 VP.n106 VP.n5 24.5923
R100 VP.n110 VP.n5 24.5923
R101 VP.n111 VP.n110 24.5923
R102 VP.n113 VP.n3 24.5923
R103 VP.n117 VP.n3 24.5923
R104 VP.n118 VP.n117 24.5923
R105 VP.n119 VP.n1 24.5923
R106 VP.n123 VP.n1 24.5923
R107 VP.n124 VP.n123 24.5923
R108 VP.n64 VP.n18 24.5923
R109 VP.n68 VP.n18 24.5923
R110 VP.n69 VP.n68 24.5923
R111 VP.n51 VP.n22 24.5923
R112 VP.n55 VP.n22 24.5923
R113 VP.n56 VP.n55 24.5923
R114 VP.n58 VP.n20 24.5923
R115 VP.n62 VP.n20 24.5923
R116 VP.n63 VP.n62 24.5923
R117 VP.n39 VP.n26 24.5923
R118 VP.n43 VP.n26 24.5923
R119 VP.n44 VP.n43 24.5923
R120 VP.n45 VP.n44 24.5923
R121 VP.n45 VP.n24 24.5923
R122 VP.n49 VP.n24 24.5923
R123 VP.n33 VP.n32 24.5923
R124 VP.n33 VP.n28 24.5923
R125 VP.n37 VP.n28 24.5923
R126 VP.n74 VP.n73 20.6576
R127 VP.n125 VP.n124 20.6576
R128 VP.n70 VP.n69 20.6576
R129 VP.n86 VP.n85 14.2638
R130 VP.n113 VP.n112 14.2638
R131 VP.n58 VP.n57 14.2638
R132 VP.n87 VP.n86 10.3291
R133 VP.n112 VP.n111 10.3291
R134 VP.n57 VP.n56 10.3291
R135 VP.n32 VP.n31 10.3291
R136 VP.n30 VP.n29 2.66362
R137 VP.n71 VP.n17 0.417304
R138 VP.n72 VP.n16 0.417304
R139 VP.n126 VP.n0 0.417304
R140 VP VP.n126 0.394524
R141 VP.n34 VP.n29 0.189894
R142 VP.n35 VP.n34 0.189894
R143 VP.n36 VP.n35 0.189894
R144 VP.n36 VP.n27 0.189894
R145 VP.n40 VP.n27 0.189894
R146 VP.n41 VP.n40 0.189894
R147 VP.n42 VP.n41 0.189894
R148 VP.n42 VP.n25 0.189894
R149 VP.n46 VP.n25 0.189894
R150 VP.n47 VP.n46 0.189894
R151 VP.n48 VP.n47 0.189894
R152 VP.n48 VP.n23 0.189894
R153 VP.n52 VP.n23 0.189894
R154 VP.n53 VP.n52 0.189894
R155 VP.n54 VP.n53 0.189894
R156 VP.n54 VP.n21 0.189894
R157 VP.n59 VP.n21 0.189894
R158 VP.n60 VP.n59 0.189894
R159 VP.n61 VP.n60 0.189894
R160 VP.n61 VP.n19 0.189894
R161 VP.n65 VP.n19 0.189894
R162 VP.n66 VP.n65 0.189894
R163 VP.n67 VP.n66 0.189894
R164 VP.n67 VP.n17 0.189894
R165 VP.n76 VP.n16 0.189894
R166 VP.n77 VP.n76 0.189894
R167 VP.n78 VP.n77 0.189894
R168 VP.n78 VP.n14 0.189894
R169 VP.n82 VP.n14 0.189894
R170 VP.n83 VP.n82 0.189894
R171 VP.n84 VP.n83 0.189894
R172 VP.n84 VP.n12 0.189894
R173 VP.n89 VP.n12 0.189894
R174 VP.n90 VP.n89 0.189894
R175 VP.n91 VP.n90 0.189894
R176 VP.n91 VP.n10 0.189894
R177 VP.n95 VP.n10 0.189894
R178 VP.n96 VP.n95 0.189894
R179 VP.n97 VP.n96 0.189894
R180 VP.n97 VP.n8 0.189894
R181 VP.n101 VP.n8 0.189894
R182 VP.n102 VP.n101 0.189894
R183 VP.n103 VP.n102 0.189894
R184 VP.n103 VP.n6 0.189894
R185 VP.n107 VP.n6 0.189894
R186 VP.n108 VP.n107 0.189894
R187 VP.n109 VP.n108 0.189894
R188 VP.n109 VP.n4 0.189894
R189 VP.n114 VP.n4 0.189894
R190 VP.n115 VP.n114 0.189894
R191 VP.n116 VP.n115 0.189894
R192 VP.n116 VP.n2 0.189894
R193 VP.n120 VP.n2 0.189894
R194 VP.n121 VP.n120 0.189894
R195 VP.n122 VP.n121 0.189894
R196 VP.n122 VP.n0 0.189894
R197 VTAIL.n352 VTAIL.n272 756.745
R198 VTAIL.n82 VTAIL.n2 756.745
R199 VTAIL.n266 VTAIL.n186 756.745
R200 VTAIL.n176 VTAIL.n96 756.745
R201 VTAIL.n301 VTAIL.n300 585
R202 VTAIL.n303 VTAIL.n302 585
R203 VTAIL.n296 VTAIL.n295 585
R204 VTAIL.n309 VTAIL.n308 585
R205 VTAIL.n311 VTAIL.n310 585
R206 VTAIL.n292 VTAIL.n291 585
R207 VTAIL.n317 VTAIL.n316 585
R208 VTAIL.n319 VTAIL.n318 585
R209 VTAIL.n288 VTAIL.n287 585
R210 VTAIL.n325 VTAIL.n324 585
R211 VTAIL.n327 VTAIL.n326 585
R212 VTAIL.n284 VTAIL.n283 585
R213 VTAIL.n333 VTAIL.n332 585
R214 VTAIL.n335 VTAIL.n334 585
R215 VTAIL.n280 VTAIL.n279 585
R216 VTAIL.n342 VTAIL.n341 585
R217 VTAIL.n343 VTAIL.n278 585
R218 VTAIL.n345 VTAIL.n344 585
R219 VTAIL.n276 VTAIL.n275 585
R220 VTAIL.n351 VTAIL.n350 585
R221 VTAIL.n353 VTAIL.n352 585
R222 VTAIL.n31 VTAIL.n30 585
R223 VTAIL.n33 VTAIL.n32 585
R224 VTAIL.n26 VTAIL.n25 585
R225 VTAIL.n39 VTAIL.n38 585
R226 VTAIL.n41 VTAIL.n40 585
R227 VTAIL.n22 VTAIL.n21 585
R228 VTAIL.n47 VTAIL.n46 585
R229 VTAIL.n49 VTAIL.n48 585
R230 VTAIL.n18 VTAIL.n17 585
R231 VTAIL.n55 VTAIL.n54 585
R232 VTAIL.n57 VTAIL.n56 585
R233 VTAIL.n14 VTAIL.n13 585
R234 VTAIL.n63 VTAIL.n62 585
R235 VTAIL.n65 VTAIL.n64 585
R236 VTAIL.n10 VTAIL.n9 585
R237 VTAIL.n72 VTAIL.n71 585
R238 VTAIL.n73 VTAIL.n8 585
R239 VTAIL.n75 VTAIL.n74 585
R240 VTAIL.n6 VTAIL.n5 585
R241 VTAIL.n81 VTAIL.n80 585
R242 VTAIL.n83 VTAIL.n82 585
R243 VTAIL.n267 VTAIL.n266 585
R244 VTAIL.n265 VTAIL.n264 585
R245 VTAIL.n190 VTAIL.n189 585
R246 VTAIL.n194 VTAIL.n192 585
R247 VTAIL.n259 VTAIL.n258 585
R248 VTAIL.n257 VTAIL.n256 585
R249 VTAIL.n196 VTAIL.n195 585
R250 VTAIL.n251 VTAIL.n250 585
R251 VTAIL.n249 VTAIL.n248 585
R252 VTAIL.n200 VTAIL.n199 585
R253 VTAIL.n243 VTAIL.n242 585
R254 VTAIL.n241 VTAIL.n240 585
R255 VTAIL.n204 VTAIL.n203 585
R256 VTAIL.n235 VTAIL.n234 585
R257 VTAIL.n233 VTAIL.n232 585
R258 VTAIL.n208 VTAIL.n207 585
R259 VTAIL.n227 VTAIL.n226 585
R260 VTAIL.n225 VTAIL.n224 585
R261 VTAIL.n212 VTAIL.n211 585
R262 VTAIL.n219 VTAIL.n218 585
R263 VTAIL.n217 VTAIL.n216 585
R264 VTAIL.n177 VTAIL.n176 585
R265 VTAIL.n175 VTAIL.n174 585
R266 VTAIL.n100 VTAIL.n99 585
R267 VTAIL.n104 VTAIL.n102 585
R268 VTAIL.n169 VTAIL.n168 585
R269 VTAIL.n167 VTAIL.n166 585
R270 VTAIL.n106 VTAIL.n105 585
R271 VTAIL.n161 VTAIL.n160 585
R272 VTAIL.n159 VTAIL.n158 585
R273 VTAIL.n110 VTAIL.n109 585
R274 VTAIL.n153 VTAIL.n152 585
R275 VTAIL.n151 VTAIL.n150 585
R276 VTAIL.n114 VTAIL.n113 585
R277 VTAIL.n145 VTAIL.n144 585
R278 VTAIL.n143 VTAIL.n142 585
R279 VTAIL.n118 VTAIL.n117 585
R280 VTAIL.n137 VTAIL.n136 585
R281 VTAIL.n135 VTAIL.n134 585
R282 VTAIL.n122 VTAIL.n121 585
R283 VTAIL.n129 VTAIL.n128 585
R284 VTAIL.n127 VTAIL.n126 585
R285 VTAIL.n299 VTAIL.t0 327.466
R286 VTAIL.n29 VTAIL.t8 327.466
R287 VTAIL.n215 VTAIL.t12 327.466
R288 VTAIL.n125 VTAIL.t19 327.466
R289 VTAIL.n302 VTAIL.n301 171.744
R290 VTAIL.n302 VTAIL.n295 171.744
R291 VTAIL.n309 VTAIL.n295 171.744
R292 VTAIL.n310 VTAIL.n309 171.744
R293 VTAIL.n310 VTAIL.n291 171.744
R294 VTAIL.n317 VTAIL.n291 171.744
R295 VTAIL.n318 VTAIL.n317 171.744
R296 VTAIL.n318 VTAIL.n287 171.744
R297 VTAIL.n325 VTAIL.n287 171.744
R298 VTAIL.n326 VTAIL.n325 171.744
R299 VTAIL.n326 VTAIL.n283 171.744
R300 VTAIL.n333 VTAIL.n283 171.744
R301 VTAIL.n334 VTAIL.n333 171.744
R302 VTAIL.n334 VTAIL.n279 171.744
R303 VTAIL.n342 VTAIL.n279 171.744
R304 VTAIL.n343 VTAIL.n342 171.744
R305 VTAIL.n344 VTAIL.n343 171.744
R306 VTAIL.n344 VTAIL.n275 171.744
R307 VTAIL.n351 VTAIL.n275 171.744
R308 VTAIL.n352 VTAIL.n351 171.744
R309 VTAIL.n32 VTAIL.n31 171.744
R310 VTAIL.n32 VTAIL.n25 171.744
R311 VTAIL.n39 VTAIL.n25 171.744
R312 VTAIL.n40 VTAIL.n39 171.744
R313 VTAIL.n40 VTAIL.n21 171.744
R314 VTAIL.n47 VTAIL.n21 171.744
R315 VTAIL.n48 VTAIL.n47 171.744
R316 VTAIL.n48 VTAIL.n17 171.744
R317 VTAIL.n55 VTAIL.n17 171.744
R318 VTAIL.n56 VTAIL.n55 171.744
R319 VTAIL.n56 VTAIL.n13 171.744
R320 VTAIL.n63 VTAIL.n13 171.744
R321 VTAIL.n64 VTAIL.n63 171.744
R322 VTAIL.n64 VTAIL.n9 171.744
R323 VTAIL.n72 VTAIL.n9 171.744
R324 VTAIL.n73 VTAIL.n72 171.744
R325 VTAIL.n74 VTAIL.n73 171.744
R326 VTAIL.n74 VTAIL.n5 171.744
R327 VTAIL.n81 VTAIL.n5 171.744
R328 VTAIL.n82 VTAIL.n81 171.744
R329 VTAIL.n266 VTAIL.n265 171.744
R330 VTAIL.n265 VTAIL.n189 171.744
R331 VTAIL.n194 VTAIL.n189 171.744
R332 VTAIL.n258 VTAIL.n194 171.744
R333 VTAIL.n258 VTAIL.n257 171.744
R334 VTAIL.n257 VTAIL.n195 171.744
R335 VTAIL.n250 VTAIL.n195 171.744
R336 VTAIL.n250 VTAIL.n249 171.744
R337 VTAIL.n249 VTAIL.n199 171.744
R338 VTAIL.n242 VTAIL.n199 171.744
R339 VTAIL.n242 VTAIL.n241 171.744
R340 VTAIL.n241 VTAIL.n203 171.744
R341 VTAIL.n234 VTAIL.n203 171.744
R342 VTAIL.n234 VTAIL.n233 171.744
R343 VTAIL.n233 VTAIL.n207 171.744
R344 VTAIL.n226 VTAIL.n207 171.744
R345 VTAIL.n226 VTAIL.n225 171.744
R346 VTAIL.n225 VTAIL.n211 171.744
R347 VTAIL.n218 VTAIL.n211 171.744
R348 VTAIL.n218 VTAIL.n217 171.744
R349 VTAIL.n176 VTAIL.n175 171.744
R350 VTAIL.n175 VTAIL.n99 171.744
R351 VTAIL.n104 VTAIL.n99 171.744
R352 VTAIL.n168 VTAIL.n104 171.744
R353 VTAIL.n168 VTAIL.n167 171.744
R354 VTAIL.n167 VTAIL.n105 171.744
R355 VTAIL.n160 VTAIL.n105 171.744
R356 VTAIL.n160 VTAIL.n159 171.744
R357 VTAIL.n159 VTAIL.n109 171.744
R358 VTAIL.n152 VTAIL.n109 171.744
R359 VTAIL.n152 VTAIL.n151 171.744
R360 VTAIL.n151 VTAIL.n113 171.744
R361 VTAIL.n144 VTAIL.n113 171.744
R362 VTAIL.n144 VTAIL.n143 171.744
R363 VTAIL.n143 VTAIL.n117 171.744
R364 VTAIL.n136 VTAIL.n117 171.744
R365 VTAIL.n136 VTAIL.n135 171.744
R366 VTAIL.n135 VTAIL.n121 171.744
R367 VTAIL.n128 VTAIL.n121 171.744
R368 VTAIL.n128 VTAIL.n127 171.744
R369 VTAIL.n301 VTAIL.t0 85.8723
R370 VTAIL.n31 VTAIL.t8 85.8723
R371 VTAIL.n217 VTAIL.t12 85.8723
R372 VTAIL.n127 VTAIL.t19 85.8723
R373 VTAIL.n185 VTAIL.n184 55.9066
R374 VTAIL.n183 VTAIL.n182 55.9066
R375 VTAIL.n95 VTAIL.n94 55.9066
R376 VTAIL.n93 VTAIL.n92 55.9066
R377 VTAIL.n359 VTAIL.n358 55.9065
R378 VTAIL.n1 VTAIL.n0 55.9065
R379 VTAIL.n89 VTAIL.n88 55.9065
R380 VTAIL.n91 VTAIL.n90 55.9065
R381 VTAIL.n357 VTAIL.n356 34.5126
R382 VTAIL.n87 VTAIL.n86 34.5126
R383 VTAIL.n271 VTAIL.n270 34.5126
R384 VTAIL.n181 VTAIL.n180 34.5126
R385 VTAIL.n93 VTAIL.n91 32.9703
R386 VTAIL.n357 VTAIL.n271 29.341
R387 VTAIL.n300 VTAIL.n299 16.3895
R388 VTAIL.n30 VTAIL.n29 16.3895
R389 VTAIL.n216 VTAIL.n215 16.3895
R390 VTAIL.n126 VTAIL.n125 16.3895
R391 VTAIL.n345 VTAIL.n276 13.1884
R392 VTAIL.n75 VTAIL.n6 13.1884
R393 VTAIL.n192 VTAIL.n190 13.1884
R394 VTAIL.n102 VTAIL.n100 13.1884
R395 VTAIL.n303 VTAIL.n298 12.8005
R396 VTAIL.n346 VTAIL.n278 12.8005
R397 VTAIL.n350 VTAIL.n349 12.8005
R398 VTAIL.n33 VTAIL.n28 12.8005
R399 VTAIL.n76 VTAIL.n8 12.8005
R400 VTAIL.n80 VTAIL.n79 12.8005
R401 VTAIL.n264 VTAIL.n263 12.8005
R402 VTAIL.n260 VTAIL.n259 12.8005
R403 VTAIL.n219 VTAIL.n214 12.8005
R404 VTAIL.n174 VTAIL.n173 12.8005
R405 VTAIL.n170 VTAIL.n169 12.8005
R406 VTAIL.n129 VTAIL.n124 12.8005
R407 VTAIL.n304 VTAIL.n296 12.0247
R408 VTAIL.n341 VTAIL.n340 12.0247
R409 VTAIL.n353 VTAIL.n274 12.0247
R410 VTAIL.n34 VTAIL.n26 12.0247
R411 VTAIL.n71 VTAIL.n70 12.0247
R412 VTAIL.n83 VTAIL.n4 12.0247
R413 VTAIL.n267 VTAIL.n188 12.0247
R414 VTAIL.n256 VTAIL.n193 12.0247
R415 VTAIL.n220 VTAIL.n212 12.0247
R416 VTAIL.n177 VTAIL.n98 12.0247
R417 VTAIL.n166 VTAIL.n103 12.0247
R418 VTAIL.n130 VTAIL.n122 12.0247
R419 VTAIL.n308 VTAIL.n307 11.249
R420 VTAIL.n339 VTAIL.n280 11.249
R421 VTAIL.n354 VTAIL.n272 11.249
R422 VTAIL.n38 VTAIL.n37 11.249
R423 VTAIL.n69 VTAIL.n10 11.249
R424 VTAIL.n84 VTAIL.n2 11.249
R425 VTAIL.n268 VTAIL.n186 11.249
R426 VTAIL.n255 VTAIL.n196 11.249
R427 VTAIL.n224 VTAIL.n223 11.249
R428 VTAIL.n178 VTAIL.n96 11.249
R429 VTAIL.n165 VTAIL.n106 11.249
R430 VTAIL.n134 VTAIL.n133 11.249
R431 VTAIL.n311 VTAIL.n294 10.4732
R432 VTAIL.n336 VTAIL.n335 10.4732
R433 VTAIL.n41 VTAIL.n24 10.4732
R434 VTAIL.n66 VTAIL.n65 10.4732
R435 VTAIL.n252 VTAIL.n251 10.4732
R436 VTAIL.n227 VTAIL.n210 10.4732
R437 VTAIL.n162 VTAIL.n161 10.4732
R438 VTAIL.n137 VTAIL.n120 10.4732
R439 VTAIL.n312 VTAIL.n292 9.69747
R440 VTAIL.n332 VTAIL.n282 9.69747
R441 VTAIL.n42 VTAIL.n22 9.69747
R442 VTAIL.n62 VTAIL.n12 9.69747
R443 VTAIL.n248 VTAIL.n198 9.69747
R444 VTAIL.n228 VTAIL.n208 9.69747
R445 VTAIL.n158 VTAIL.n108 9.69747
R446 VTAIL.n138 VTAIL.n118 9.69747
R447 VTAIL.n356 VTAIL.n355 9.45567
R448 VTAIL.n86 VTAIL.n85 9.45567
R449 VTAIL.n270 VTAIL.n269 9.45567
R450 VTAIL.n180 VTAIL.n179 9.45567
R451 VTAIL.n355 VTAIL.n354 9.3005
R452 VTAIL.n274 VTAIL.n273 9.3005
R453 VTAIL.n349 VTAIL.n348 9.3005
R454 VTAIL.n321 VTAIL.n320 9.3005
R455 VTAIL.n290 VTAIL.n289 9.3005
R456 VTAIL.n315 VTAIL.n314 9.3005
R457 VTAIL.n313 VTAIL.n312 9.3005
R458 VTAIL.n294 VTAIL.n293 9.3005
R459 VTAIL.n307 VTAIL.n306 9.3005
R460 VTAIL.n305 VTAIL.n304 9.3005
R461 VTAIL.n298 VTAIL.n297 9.3005
R462 VTAIL.n323 VTAIL.n322 9.3005
R463 VTAIL.n286 VTAIL.n285 9.3005
R464 VTAIL.n329 VTAIL.n328 9.3005
R465 VTAIL.n331 VTAIL.n330 9.3005
R466 VTAIL.n282 VTAIL.n281 9.3005
R467 VTAIL.n337 VTAIL.n336 9.3005
R468 VTAIL.n339 VTAIL.n338 9.3005
R469 VTAIL.n340 VTAIL.n277 9.3005
R470 VTAIL.n347 VTAIL.n346 9.3005
R471 VTAIL.n85 VTAIL.n84 9.3005
R472 VTAIL.n4 VTAIL.n3 9.3005
R473 VTAIL.n79 VTAIL.n78 9.3005
R474 VTAIL.n51 VTAIL.n50 9.3005
R475 VTAIL.n20 VTAIL.n19 9.3005
R476 VTAIL.n45 VTAIL.n44 9.3005
R477 VTAIL.n43 VTAIL.n42 9.3005
R478 VTAIL.n24 VTAIL.n23 9.3005
R479 VTAIL.n37 VTAIL.n36 9.3005
R480 VTAIL.n35 VTAIL.n34 9.3005
R481 VTAIL.n28 VTAIL.n27 9.3005
R482 VTAIL.n53 VTAIL.n52 9.3005
R483 VTAIL.n16 VTAIL.n15 9.3005
R484 VTAIL.n59 VTAIL.n58 9.3005
R485 VTAIL.n61 VTAIL.n60 9.3005
R486 VTAIL.n12 VTAIL.n11 9.3005
R487 VTAIL.n67 VTAIL.n66 9.3005
R488 VTAIL.n69 VTAIL.n68 9.3005
R489 VTAIL.n70 VTAIL.n7 9.3005
R490 VTAIL.n77 VTAIL.n76 9.3005
R491 VTAIL.n202 VTAIL.n201 9.3005
R492 VTAIL.n245 VTAIL.n244 9.3005
R493 VTAIL.n247 VTAIL.n246 9.3005
R494 VTAIL.n198 VTAIL.n197 9.3005
R495 VTAIL.n253 VTAIL.n252 9.3005
R496 VTAIL.n255 VTAIL.n254 9.3005
R497 VTAIL.n193 VTAIL.n191 9.3005
R498 VTAIL.n261 VTAIL.n260 9.3005
R499 VTAIL.n269 VTAIL.n268 9.3005
R500 VTAIL.n188 VTAIL.n187 9.3005
R501 VTAIL.n263 VTAIL.n262 9.3005
R502 VTAIL.n239 VTAIL.n238 9.3005
R503 VTAIL.n237 VTAIL.n236 9.3005
R504 VTAIL.n206 VTAIL.n205 9.3005
R505 VTAIL.n231 VTAIL.n230 9.3005
R506 VTAIL.n229 VTAIL.n228 9.3005
R507 VTAIL.n210 VTAIL.n209 9.3005
R508 VTAIL.n223 VTAIL.n222 9.3005
R509 VTAIL.n221 VTAIL.n220 9.3005
R510 VTAIL.n214 VTAIL.n213 9.3005
R511 VTAIL.n112 VTAIL.n111 9.3005
R512 VTAIL.n155 VTAIL.n154 9.3005
R513 VTAIL.n157 VTAIL.n156 9.3005
R514 VTAIL.n108 VTAIL.n107 9.3005
R515 VTAIL.n163 VTAIL.n162 9.3005
R516 VTAIL.n165 VTAIL.n164 9.3005
R517 VTAIL.n103 VTAIL.n101 9.3005
R518 VTAIL.n171 VTAIL.n170 9.3005
R519 VTAIL.n179 VTAIL.n178 9.3005
R520 VTAIL.n98 VTAIL.n97 9.3005
R521 VTAIL.n173 VTAIL.n172 9.3005
R522 VTAIL.n149 VTAIL.n148 9.3005
R523 VTAIL.n147 VTAIL.n146 9.3005
R524 VTAIL.n116 VTAIL.n115 9.3005
R525 VTAIL.n141 VTAIL.n140 9.3005
R526 VTAIL.n139 VTAIL.n138 9.3005
R527 VTAIL.n120 VTAIL.n119 9.3005
R528 VTAIL.n133 VTAIL.n132 9.3005
R529 VTAIL.n131 VTAIL.n130 9.3005
R530 VTAIL.n124 VTAIL.n123 9.3005
R531 VTAIL.n316 VTAIL.n315 8.92171
R532 VTAIL.n331 VTAIL.n284 8.92171
R533 VTAIL.n46 VTAIL.n45 8.92171
R534 VTAIL.n61 VTAIL.n14 8.92171
R535 VTAIL.n247 VTAIL.n200 8.92171
R536 VTAIL.n232 VTAIL.n231 8.92171
R537 VTAIL.n157 VTAIL.n110 8.92171
R538 VTAIL.n142 VTAIL.n141 8.92171
R539 VTAIL.n319 VTAIL.n290 8.14595
R540 VTAIL.n328 VTAIL.n327 8.14595
R541 VTAIL.n49 VTAIL.n20 8.14595
R542 VTAIL.n58 VTAIL.n57 8.14595
R543 VTAIL.n244 VTAIL.n243 8.14595
R544 VTAIL.n235 VTAIL.n206 8.14595
R545 VTAIL.n154 VTAIL.n153 8.14595
R546 VTAIL.n145 VTAIL.n116 8.14595
R547 VTAIL.n320 VTAIL.n288 7.3702
R548 VTAIL.n324 VTAIL.n286 7.3702
R549 VTAIL.n50 VTAIL.n18 7.3702
R550 VTAIL.n54 VTAIL.n16 7.3702
R551 VTAIL.n240 VTAIL.n202 7.3702
R552 VTAIL.n236 VTAIL.n204 7.3702
R553 VTAIL.n150 VTAIL.n112 7.3702
R554 VTAIL.n146 VTAIL.n114 7.3702
R555 VTAIL.n323 VTAIL.n288 6.59444
R556 VTAIL.n324 VTAIL.n323 6.59444
R557 VTAIL.n53 VTAIL.n18 6.59444
R558 VTAIL.n54 VTAIL.n53 6.59444
R559 VTAIL.n240 VTAIL.n239 6.59444
R560 VTAIL.n239 VTAIL.n204 6.59444
R561 VTAIL.n150 VTAIL.n149 6.59444
R562 VTAIL.n149 VTAIL.n114 6.59444
R563 VTAIL.n320 VTAIL.n319 5.81868
R564 VTAIL.n327 VTAIL.n286 5.81868
R565 VTAIL.n50 VTAIL.n49 5.81868
R566 VTAIL.n57 VTAIL.n16 5.81868
R567 VTAIL.n243 VTAIL.n202 5.81868
R568 VTAIL.n236 VTAIL.n235 5.81868
R569 VTAIL.n153 VTAIL.n112 5.81868
R570 VTAIL.n146 VTAIL.n145 5.81868
R571 VTAIL.n316 VTAIL.n290 5.04292
R572 VTAIL.n328 VTAIL.n284 5.04292
R573 VTAIL.n46 VTAIL.n20 5.04292
R574 VTAIL.n58 VTAIL.n14 5.04292
R575 VTAIL.n244 VTAIL.n200 5.04292
R576 VTAIL.n232 VTAIL.n206 5.04292
R577 VTAIL.n154 VTAIL.n110 5.04292
R578 VTAIL.n142 VTAIL.n116 5.04292
R579 VTAIL.n315 VTAIL.n292 4.26717
R580 VTAIL.n332 VTAIL.n331 4.26717
R581 VTAIL.n45 VTAIL.n22 4.26717
R582 VTAIL.n62 VTAIL.n61 4.26717
R583 VTAIL.n248 VTAIL.n247 4.26717
R584 VTAIL.n231 VTAIL.n208 4.26717
R585 VTAIL.n158 VTAIL.n157 4.26717
R586 VTAIL.n141 VTAIL.n118 4.26717
R587 VTAIL.n299 VTAIL.n297 3.70982
R588 VTAIL.n29 VTAIL.n27 3.70982
R589 VTAIL.n215 VTAIL.n213 3.70982
R590 VTAIL.n125 VTAIL.n123 3.70982
R591 VTAIL.n95 VTAIL.n93 3.62981
R592 VTAIL.n181 VTAIL.n95 3.62981
R593 VTAIL.n185 VTAIL.n183 3.62981
R594 VTAIL.n271 VTAIL.n185 3.62981
R595 VTAIL.n91 VTAIL.n89 3.62981
R596 VTAIL.n89 VTAIL.n87 3.62981
R597 VTAIL.n359 VTAIL.n357 3.62981
R598 VTAIL.n312 VTAIL.n311 3.49141
R599 VTAIL.n335 VTAIL.n282 3.49141
R600 VTAIL.n42 VTAIL.n41 3.49141
R601 VTAIL.n65 VTAIL.n12 3.49141
R602 VTAIL.n251 VTAIL.n198 3.49141
R603 VTAIL.n228 VTAIL.n227 3.49141
R604 VTAIL.n161 VTAIL.n108 3.49141
R605 VTAIL.n138 VTAIL.n137 3.49141
R606 VTAIL VTAIL.n1 2.78067
R607 VTAIL.n308 VTAIL.n294 2.71565
R608 VTAIL.n336 VTAIL.n280 2.71565
R609 VTAIL.n356 VTAIL.n272 2.71565
R610 VTAIL.n38 VTAIL.n24 2.71565
R611 VTAIL.n66 VTAIL.n10 2.71565
R612 VTAIL.n86 VTAIL.n2 2.71565
R613 VTAIL.n270 VTAIL.n186 2.71565
R614 VTAIL.n252 VTAIL.n196 2.71565
R615 VTAIL.n224 VTAIL.n210 2.71565
R616 VTAIL.n180 VTAIL.n96 2.71565
R617 VTAIL.n162 VTAIL.n106 2.71565
R618 VTAIL.n134 VTAIL.n120 2.71565
R619 VTAIL.n183 VTAIL.n181 2.28498
R620 VTAIL.n87 VTAIL.n1 2.28498
R621 VTAIL.n358 VTAIL.t1 2.10031
R622 VTAIL.n358 VTAIL.t4 2.10031
R623 VTAIL.n0 VTAIL.t2 2.10031
R624 VTAIL.n0 VTAIL.t18 2.10031
R625 VTAIL.n88 VTAIL.t17 2.10031
R626 VTAIL.n88 VTAIL.t13 2.10031
R627 VTAIL.n90 VTAIL.t16 2.10031
R628 VTAIL.n90 VTAIL.t10 2.10031
R629 VTAIL.n184 VTAIL.t14 2.10031
R630 VTAIL.n184 VTAIL.t9 2.10031
R631 VTAIL.n182 VTAIL.t15 2.10031
R632 VTAIL.n182 VTAIL.t11 2.10031
R633 VTAIL.n94 VTAIL.t3 2.10031
R634 VTAIL.n94 VTAIL.t5 2.10031
R635 VTAIL.n92 VTAIL.t7 2.10031
R636 VTAIL.n92 VTAIL.t6 2.10031
R637 VTAIL.n307 VTAIL.n296 1.93989
R638 VTAIL.n341 VTAIL.n339 1.93989
R639 VTAIL.n354 VTAIL.n353 1.93989
R640 VTAIL.n37 VTAIL.n26 1.93989
R641 VTAIL.n71 VTAIL.n69 1.93989
R642 VTAIL.n84 VTAIL.n83 1.93989
R643 VTAIL.n268 VTAIL.n267 1.93989
R644 VTAIL.n256 VTAIL.n255 1.93989
R645 VTAIL.n223 VTAIL.n212 1.93989
R646 VTAIL.n178 VTAIL.n177 1.93989
R647 VTAIL.n166 VTAIL.n165 1.93989
R648 VTAIL.n133 VTAIL.n122 1.93989
R649 VTAIL.n304 VTAIL.n303 1.16414
R650 VTAIL.n340 VTAIL.n278 1.16414
R651 VTAIL.n350 VTAIL.n274 1.16414
R652 VTAIL.n34 VTAIL.n33 1.16414
R653 VTAIL.n70 VTAIL.n8 1.16414
R654 VTAIL.n80 VTAIL.n4 1.16414
R655 VTAIL.n264 VTAIL.n188 1.16414
R656 VTAIL.n259 VTAIL.n193 1.16414
R657 VTAIL.n220 VTAIL.n219 1.16414
R658 VTAIL.n174 VTAIL.n98 1.16414
R659 VTAIL.n169 VTAIL.n103 1.16414
R660 VTAIL.n130 VTAIL.n129 1.16414
R661 VTAIL VTAIL.n359 0.849638
R662 VTAIL.n300 VTAIL.n298 0.388379
R663 VTAIL.n346 VTAIL.n345 0.388379
R664 VTAIL.n349 VTAIL.n276 0.388379
R665 VTAIL.n30 VTAIL.n28 0.388379
R666 VTAIL.n76 VTAIL.n75 0.388379
R667 VTAIL.n79 VTAIL.n6 0.388379
R668 VTAIL.n263 VTAIL.n190 0.388379
R669 VTAIL.n260 VTAIL.n192 0.388379
R670 VTAIL.n216 VTAIL.n214 0.388379
R671 VTAIL.n173 VTAIL.n100 0.388379
R672 VTAIL.n170 VTAIL.n102 0.388379
R673 VTAIL.n126 VTAIL.n124 0.388379
R674 VTAIL.n305 VTAIL.n297 0.155672
R675 VTAIL.n306 VTAIL.n305 0.155672
R676 VTAIL.n306 VTAIL.n293 0.155672
R677 VTAIL.n313 VTAIL.n293 0.155672
R678 VTAIL.n314 VTAIL.n313 0.155672
R679 VTAIL.n314 VTAIL.n289 0.155672
R680 VTAIL.n321 VTAIL.n289 0.155672
R681 VTAIL.n322 VTAIL.n321 0.155672
R682 VTAIL.n322 VTAIL.n285 0.155672
R683 VTAIL.n329 VTAIL.n285 0.155672
R684 VTAIL.n330 VTAIL.n329 0.155672
R685 VTAIL.n330 VTAIL.n281 0.155672
R686 VTAIL.n337 VTAIL.n281 0.155672
R687 VTAIL.n338 VTAIL.n337 0.155672
R688 VTAIL.n338 VTAIL.n277 0.155672
R689 VTAIL.n347 VTAIL.n277 0.155672
R690 VTAIL.n348 VTAIL.n347 0.155672
R691 VTAIL.n348 VTAIL.n273 0.155672
R692 VTAIL.n355 VTAIL.n273 0.155672
R693 VTAIL.n35 VTAIL.n27 0.155672
R694 VTAIL.n36 VTAIL.n35 0.155672
R695 VTAIL.n36 VTAIL.n23 0.155672
R696 VTAIL.n43 VTAIL.n23 0.155672
R697 VTAIL.n44 VTAIL.n43 0.155672
R698 VTAIL.n44 VTAIL.n19 0.155672
R699 VTAIL.n51 VTAIL.n19 0.155672
R700 VTAIL.n52 VTAIL.n51 0.155672
R701 VTAIL.n52 VTAIL.n15 0.155672
R702 VTAIL.n59 VTAIL.n15 0.155672
R703 VTAIL.n60 VTAIL.n59 0.155672
R704 VTAIL.n60 VTAIL.n11 0.155672
R705 VTAIL.n67 VTAIL.n11 0.155672
R706 VTAIL.n68 VTAIL.n67 0.155672
R707 VTAIL.n68 VTAIL.n7 0.155672
R708 VTAIL.n77 VTAIL.n7 0.155672
R709 VTAIL.n78 VTAIL.n77 0.155672
R710 VTAIL.n78 VTAIL.n3 0.155672
R711 VTAIL.n85 VTAIL.n3 0.155672
R712 VTAIL.n269 VTAIL.n187 0.155672
R713 VTAIL.n262 VTAIL.n187 0.155672
R714 VTAIL.n262 VTAIL.n261 0.155672
R715 VTAIL.n261 VTAIL.n191 0.155672
R716 VTAIL.n254 VTAIL.n191 0.155672
R717 VTAIL.n254 VTAIL.n253 0.155672
R718 VTAIL.n253 VTAIL.n197 0.155672
R719 VTAIL.n246 VTAIL.n197 0.155672
R720 VTAIL.n246 VTAIL.n245 0.155672
R721 VTAIL.n245 VTAIL.n201 0.155672
R722 VTAIL.n238 VTAIL.n201 0.155672
R723 VTAIL.n238 VTAIL.n237 0.155672
R724 VTAIL.n237 VTAIL.n205 0.155672
R725 VTAIL.n230 VTAIL.n205 0.155672
R726 VTAIL.n230 VTAIL.n229 0.155672
R727 VTAIL.n229 VTAIL.n209 0.155672
R728 VTAIL.n222 VTAIL.n209 0.155672
R729 VTAIL.n222 VTAIL.n221 0.155672
R730 VTAIL.n221 VTAIL.n213 0.155672
R731 VTAIL.n179 VTAIL.n97 0.155672
R732 VTAIL.n172 VTAIL.n97 0.155672
R733 VTAIL.n172 VTAIL.n171 0.155672
R734 VTAIL.n171 VTAIL.n101 0.155672
R735 VTAIL.n164 VTAIL.n101 0.155672
R736 VTAIL.n164 VTAIL.n163 0.155672
R737 VTAIL.n163 VTAIL.n107 0.155672
R738 VTAIL.n156 VTAIL.n107 0.155672
R739 VTAIL.n156 VTAIL.n155 0.155672
R740 VTAIL.n155 VTAIL.n111 0.155672
R741 VTAIL.n148 VTAIL.n111 0.155672
R742 VTAIL.n148 VTAIL.n147 0.155672
R743 VTAIL.n147 VTAIL.n115 0.155672
R744 VTAIL.n140 VTAIL.n115 0.155672
R745 VTAIL.n140 VTAIL.n139 0.155672
R746 VTAIL.n139 VTAIL.n119 0.155672
R747 VTAIL.n132 VTAIL.n119 0.155672
R748 VTAIL.n132 VTAIL.n131 0.155672
R749 VTAIL.n131 VTAIL.n123 0.155672
R750 VDD1.n80 VDD1.n0 756.745
R751 VDD1.n167 VDD1.n87 756.745
R752 VDD1.n81 VDD1.n80 585
R753 VDD1.n79 VDD1.n78 585
R754 VDD1.n4 VDD1.n3 585
R755 VDD1.n8 VDD1.n6 585
R756 VDD1.n73 VDD1.n72 585
R757 VDD1.n71 VDD1.n70 585
R758 VDD1.n10 VDD1.n9 585
R759 VDD1.n65 VDD1.n64 585
R760 VDD1.n63 VDD1.n62 585
R761 VDD1.n14 VDD1.n13 585
R762 VDD1.n57 VDD1.n56 585
R763 VDD1.n55 VDD1.n54 585
R764 VDD1.n18 VDD1.n17 585
R765 VDD1.n49 VDD1.n48 585
R766 VDD1.n47 VDD1.n46 585
R767 VDD1.n22 VDD1.n21 585
R768 VDD1.n41 VDD1.n40 585
R769 VDD1.n39 VDD1.n38 585
R770 VDD1.n26 VDD1.n25 585
R771 VDD1.n33 VDD1.n32 585
R772 VDD1.n31 VDD1.n30 585
R773 VDD1.n116 VDD1.n115 585
R774 VDD1.n118 VDD1.n117 585
R775 VDD1.n111 VDD1.n110 585
R776 VDD1.n124 VDD1.n123 585
R777 VDD1.n126 VDD1.n125 585
R778 VDD1.n107 VDD1.n106 585
R779 VDD1.n132 VDD1.n131 585
R780 VDD1.n134 VDD1.n133 585
R781 VDD1.n103 VDD1.n102 585
R782 VDD1.n140 VDD1.n139 585
R783 VDD1.n142 VDD1.n141 585
R784 VDD1.n99 VDD1.n98 585
R785 VDD1.n148 VDD1.n147 585
R786 VDD1.n150 VDD1.n149 585
R787 VDD1.n95 VDD1.n94 585
R788 VDD1.n157 VDD1.n156 585
R789 VDD1.n158 VDD1.n93 585
R790 VDD1.n160 VDD1.n159 585
R791 VDD1.n91 VDD1.n90 585
R792 VDD1.n166 VDD1.n165 585
R793 VDD1.n168 VDD1.n167 585
R794 VDD1.n29 VDD1.t3 327.466
R795 VDD1.n114 VDD1.t9 327.466
R796 VDD1.n80 VDD1.n79 171.744
R797 VDD1.n79 VDD1.n3 171.744
R798 VDD1.n8 VDD1.n3 171.744
R799 VDD1.n72 VDD1.n8 171.744
R800 VDD1.n72 VDD1.n71 171.744
R801 VDD1.n71 VDD1.n9 171.744
R802 VDD1.n64 VDD1.n9 171.744
R803 VDD1.n64 VDD1.n63 171.744
R804 VDD1.n63 VDD1.n13 171.744
R805 VDD1.n56 VDD1.n13 171.744
R806 VDD1.n56 VDD1.n55 171.744
R807 VDD1.n55 VDD1.n17 171.744
R808 VDD1.n48 VDD1.n17 171.744
R809 VDD1.n48 VDD1.n47 171.744
R810 VDD1.n47 VDD1.n21 171.744
R811 VDD1.n40 VDD1.n21 171.744
R812 VDD1.n40 VDD1.n39 171.744
R813 VDD1.n39 VDD1.n25 171.744
R814 VDD1.n32 VDD1.n25 171.744
R815 VDD1.n32 VDD1.n31 171.744
R816 VDD1.n117 VDD1.n116 171.744
R817 VDD1.n117 VDD1.n110 171.744
R818 VDD1.n124 VDD1.n110 171.744
R819 VDD1.n125 VDD1.n124 171.744
R820 VDD1.n125 VDD1.n106 171.744
R821 VDD1.n132 VDD1.n106 171.744
R822 VDD1.n133 VDD1.n132 171.744
R823 VDD1.n133 VDD1.n102 171.744
R824 VDD1.n140 VDD1.n102 171.744
R825 VDD1.n141 VDD1.n140 171.744
R826 VDD1.n141 VDD1.n98 171.744
R827 VDD1.n148 VDD1.n98 171.744
R828 VDD1.n149 VDD1.n148 171.744
R829 VDD1.n149 VDD1.n94 171.744
R830 VDD1.n157 VDD1.n94 171.744
R831 VDD1.n158 VDD1.n157 171.744
R832 VDD1.n159 VDD1.n158 171.744
R833 VDD1.n159 VDD1.n90 171.744
R834 VDD1.n166 VDD1.n90 171.744
R835 VDD1.n167 VDD1.n166 171.744
R836 VDD1.n31 VDD1.t3 85.8723
R837 VDD1.n116 VDD1.t9 85.8723
R838 VDD1.n175 VDD1.n174 75.2519
R839 VDD1.n86 VDD1.n85 72.5854
R840 VDD1.n173 VDD1.n172 72.5852
R841 VDD1.n177 VDD1.n176 72.5852
R842 VDD1.n177 VDD1.n175 56.697
R843 VDD1.n86 VDD1.n84 54.8207
R844 VDD1.n173 VDD1.n171 54.8207
R845 VDD1.n30 VDD1.n29 16.3895
R846 VDD1.n115 VDD1.n114 16.3895
R847 VDD1.n6 VDD1.n4 13.1884
R848 VDD1.n160 VDD1.n91 13.1884
R849 VDD1.n78 VDD1.n77 12.8005
R850 VDD1.n74 VDD1.n73 12.8005
R851 VDD1.n33 VDD1.n28 12.8005
R852 VDD1.n118 VDD1.n113 12.8005
R853 VDD1.n161 VDD1.n93 12.8005
R854 VDD1.n165 VDD1.n164 12.8005
R855 VDD1.n81 VDD1.n2 12.0247
R856 VDD1.n70 VDD1.n7 12.0247
R857 VDD1.n34 VDD1.n26 12.0247
R858 VDD1.n119 VDD1.n111 12.0247
R859 VDD1.n156 VDD1.n155 12.0247
R860 VDD1.n168 VDD1.n89 12.0247
R861 VDD1.n82 VDD1.n0 11.249
R862 VDD1.n69 VDD1.n10 11.249
R863 VDD1.n38 VDD1.n37 11.249
R864 VDD1.n123 VDD1.n122 11.249
R865 VDD1.n154 VDD1.n95 11.249
R866 VDD1.n169 VDD1.n87 11.249
R867 VDD1.n66 VDD1.n65 10.4732
R868 VDD1.n41 VDD1.n24 10.4732
R869 VDD1.n126 VDD1.n109 10.4732
R870 VDD1.n151 VDD1.n150 10.4732
R871 VDD1.n62 VDD1.n12 9.69747
R872 VDD1.n42 VDD1.n22 9.69747
R873 VDD1.n127 VDD1.n107 9.69747
R874 VDD1.n147 VDD1.n97 9.69747
R875 VDD1.n84 VDD1.n83 9.45567
R876 VDD1.n171 VDD1.n170 9.45567
R877 VDD1.n16 VDD1.n15 9.3005
R878 VDD1.n59 VDD1.n58 9.3005
R879 VDD1.n61 VDD1.n60 9.3005
R880 VDD1.n12 VDD1.n11 9.3005
R881 VDD1.n67 VDD1.n66 9.3005
R882 VDD1.n69 VDD1.n68 9.3005
R883 VDD1.n7 VDD1.n5 9.3005
R884 VDD1.n75 VDD1.n74 9.3005
R885 VDD1.n83 VDD1.n82 9.3005
R886 VDD1.n2 VDD1.n1 9.3005
R887 VDD1.n77 VDD1.n76 9.3005
R888 VDD1.n53 VDD1.n52 9.3005
R889 VDD1.n51 VDD1.n50 9.3005
R890 VDD1.n20 VDD1.n19 9.3005
R891 VDD1.n45 VDD1.n44 9.3005
R892 VDD1.n43 VDD1.n42 9.3005
R893 VDD1.n24 VDD1.n23 9.3005
R894 VDD1.n37 VDD1.n36 9.3005
R895 VDD1.n35 VDD1.n34 9.3005
R896 VDD1.n28 VDD1.n27 9.3005
R897 VDD1.n170 VDD1.n169 9.3005
R898 VDD1.n89 VDD1.n88 9.3005
R899 VDD1.n164 VDD1.n163 9.3005
R900 VDD1.n136 VDD1.n135 9.3005
R901 VDD1.n105 VDD1.n104 9.3005
R902 VDD1.n130 VDD1.n129 9.3005
R903 VDD1.n128 VDD1.n127 9.3005
R904 VDD1.n109 VDD1.n108 9.3005
R905 VDD1.n122 VDD1.n121 9.3005
R906 VDD1.n120 VDD1.n119 9.3005
R907 VDD1.n113 VDD1.n112 9.3005
R908 VDD1.n138 VDD1.n137 9.3005
R909 VDD1.n101 VDD1.n100 9.3005
R910 VDD1.n144 VDD1.n143 9.3005
R911 VDD1.n146 VDD1.n145 9.3005
R912 VDD1.n97 VDD1.n96 9.3005
R913 VDD1.n152 VDD1.n151 9.3005
R914 VDD1.n154 VDD1.n153 9.3005
R915 VDD1.n155 VDD1.n92 9.3005
R916 VDD1.n162 VDD1.n161 9.3005
R917 VDD1.n61 VDD1.n14 8.92171
R918 VDD1.n46 VDD1.n45 8.92171
R919 VDD1.n131 VDD1.n130 8.92171
R920 VDD1.n146 VDD1.n99 8.92171
R921 VDD1.n58 VDD1.n57 8.14595
R922 VDD1.n49 VDD1.n20 8.14595
R923 VDD1.n134 VDD1.n105 8.14595
R924 VDD1.n143 VDD1.n142 8.14595
R925 VDD1.n54 VDD1.n16 7.3702
R926 VDD1.n50 VDD1.n18 7.3702
R927 VDD1.n135 VDD1.n103 7.3702
R928 VDD1.n139 VDD1.n101 7.3702
R929 VDD1.n54 VDD1.n53 6.59444
R930 VDD1.n53 VDD1.n18 6.59444
R931 VDD1.n138 VDD1.n103 6.59444
R932 VDD1.n139 VDD1.n138 6.59444
R933 VDD1.n57 VDD1.n16 5.81868
R934 VDD1.n50 VDD1.n49 5.81868
R935 VDD1.n135 VDD1.n134 5.81868
R936 VDD1.n142 VDD1.n101 5.81868
R937 VDD1.n58 VDD1.n14 5.04292
R938 VDD1.n46 VDD1.n20 5.04292
R939 VDD1.n131 VDD1.n105 5.04292
R940 VDD1.n143 VDD1.n99 5.04292
R941 VDD1.n62 VDD1.n61 4.26717
R942 VDD1.n45 VDD1.n22 4.26717
R943 VDD1.n130 VDD1.n107 4.26717
R944 VDD1.n147 VDD1.n146 4.26717
R945 VDD1.n29 VDD1.n27 3.70982
R946 VDD1.n114 VDD1.n112 3.70982
R947 VDD1.n65 VDD1.n12 3.49141
R948 VDD1.n42 VDD1.n41 3.49141
R949 VDD1.n127 VDD1.n126 3.49141
R950 VDD1.n150 VDD1.n97 3.49141
R951 VDD1.n84 VDD1.n0 2.71565
R952 VDD1.n66 VDD1.n10 2.71565
R953 VDD1.n38 VDD1.n24 2.71565
R954 VDD1.n123 VDD1.n109 2.71565
R955 VDD1.n151 VDD1.n95 2.71565
R956 VDD1.n171 VDD1.n87 2.71565
R957 VDD1 VDD1.n177 2.66429
R958 VDD1.n176 VDD1.t7 2.10031
R959 VDD1.n176 VDD1.t0 2.10031
R960 VDD1.n85 VDD1.t4 2.10031
R961 VDD1.n85 VDD1.t5 2.10031
R962 VDD1.n174 VDD1.t1 2.10031
R963 VDD1.n174 VDD1.t8 2.10031
R964 VDD1.n172 VDD1.t6 2.10031
R965 VDD1.n172 VDD1.t2 2.10031
R966 VDD1.n82 VDD1.n81 1.93989
R967 VDD1.n70 VDD1.n69 1.93989
R968 VDD1.n37 VDD1.n26 1.93989
R969 VDD1.n122 VDD1.n111 1.93989
R970 VDD1.n156 VDD1.n154 1.93989
R971 VDD1.n169 VDD1.n168 1.93989
R972 VDD1.n78 VDD1.n2 1.16414
R973 VDD1.n73 VDD1.n7 1.16414
R974 VDD1.n34 VDD1.n33 1.16414
R975 VDD1.n119 VDD1.n118 1.16414
R976 VDD1.n155 VDD1.n93 1.16414
R977 VDD1.n165 VDD1.n89 1.16414
R978 VDD1 VDD1.n86 0.966017
R979 VDD1.n175 VDD1.n173 0.852482
R980 VDD1.n77 VDD1.n4 0.388379
R981 VDD1.n74 VDD1.n6 0.388379
R982 VDD1.n30 VDD1.n28 0.388379
R983 VDD1.n115 VDD1.n113 0.388379
R984 VDD1.n161 VDD1.n160 0.388379
R985 VDD1.n164 VDD1.n91 0.388379
R986 VDD1.n83 VDD1.n1 0.155672
R987 VDD1.n76 VDD1.n1 0.155672
R988 VDD1.n76 VDD1.n75 0.155672
R989 VDD1.n75 VDD1.n5 0.155672
R990 VDD1.n68 VDD1.n5 0.155672
R991 VDD1.n68 VDD1.n67 0.155672
R992 VDD1.n67 VDD1.n11 0.155672
R993 VDD1.n60 VDD1.n11 0.155672
R994 VDD1.n60 VDD1.n59 0.155672
R995 VDD1.n59 VDD1.n15 0.155672
R996 VDD1.n52 VDD1.n15 0.155672
R997 VDD1.n52 VDD1.n51 0.155672
R998 VDD1.n51 VDD1.n19 0.155672
R999 VDD1.n44 VDD1.n19 0.155672
R1000 VDD1.n44 VDD1.n43 0.155672
R1001 VDD1.n43 VDD1.n23 0.155672
R1002 VDD1.n36 VDD1.n23 0.155672
R1003 VDD1.n36 VDD1.n35 0.155672
R1004 VDD1.n35 VDD1.n27 0.155672
R1005 VDD1.n120 VDD1.n112 0.155672
R1006 VDD1.n121 VDD1.n120 0.155672
R1007 VDD1.n121 VDD1.n108 0.155672
R1008 VDD1.n128 VDD1.n108 0.155672
R1009 VDD1.n129 VDD1.n128 0.155672
R1010 VDD1.n129 VDD1.n104 0.155672
R1011 VDD1.n136 VDD1.n104 0.155672
R1012 VDD1.n137 VDD1.n136 0.155672
R1013 VDD1.n137 VDD1.n100 0.155672
R1014 VDD1.n144 VDD1.n100 0.155672
R1015 VDD1.n145 VDD1.n144 0.155672
R1016 VDD1.n145 VDD1.n96 0.155672
R1017 VDD1.n152 VDD1.n96 0.155672
R1018 VDD1.n153 VDD1.n152 0.155672
R1019 VDD1.n153 VDD1.n92 0.155672
R1020 VDD1.n162 VDD1.n92 0.155672
R1021 VDD1.n163 VDD1.n162 0.155672
R1022 VDD1.n163 VDD1.n88 0.155672
R1023 VDD1.n170 VDD1.n88 0.155672
R1024 VN.n107 VN.n55 161.3
R1025 VN.n106 VN.n105 161.3
R1026 VN.n104 VN.n56 161.3
R1027 VN.n103 VN.n102 161.3
R1028 VN.n101 VN.n57 161.3
R1029 VN.n100 VN.n99 161.3
R1030 VN.n98 VN.n58 161.3
R1031 VN.n97 VN.n96 161.3
R1032 VN.n94 VN.n59 161.3
R1033 VN.n93 VN.n92 161.3
R1034 VN.n91 VN.n60 161.3
R1035 VN.n90 VN.n89 161.3
R1036 VN.n88 VN.n61 161.3
R1037 VN.n87 VN.n86 161.3
R1038 VN.n85 VN.n62 161.3
R1039 VN.n84 VN.n83 161.3
R1040 VN.n82 VN.n63 161.3
R1041 VN.n81 VN.n80 161.3
R1042 VN.n79 VN.n64 161.3
R1043 VN.n78 VN.n77 161.3
R1044 VN.n76 VN.n65 161.3
R1045 VN.n75 VN.n74 161.3
R1046 VN.n73 VN.n66 161.3
R1047 VN.n72 VN.n71 161.3
R1048 VN.n70 VN.n67 161.3
R1049 VN.n52 VN.n0 161.3
R1050 VN.n51 VN.n50 161.3
R1051 VN.n49 VN.n1 161.3
R1052 VN.n48 VN.n47 161.3
R1053 VN.n46 VN.n2 161.3
R1054 VN.n45 VN.n44 161.3
R1055 VN.n43 VN.n3 161.3
R1056 VN.n42 VN.n41 161.3
R1057 VN.n39 VN.n4 161.3
R1058 VN.n38 VN.n37 161.3
R1059 VN.n36 VN.n5 161.3
R1060 VN.n35 VN.n34 161.3
R1061 VN.n33 VN.n6 161.3
R1062 VN.n32 VN.n31 161.3
R1063 VN.n30 VN.n7 161.3
R1064 VN.n29 VN.n28 161.3
R1065 VN.n27 VN.n8 161.3
R1066 VN.n26 VN.n25 161.3
R1067 VN.n24 VN.n9 161.3
R1068 VN.n23 VN.n22 161.3
R1069 VN.n21 VN.n10 161.3
R1070 VN.n20 VN.n19 161.3
R1071 VN.n18 VN.n11 161.3
R1072 VN.n17 VN.n16 161.3
R1073 VN.n15 VN.n12 161.3
R1074 VN.n13 VN.t9 128.482
R1075 VN.n68 VN.t6 128.482
R1076 VN.n27 VN.t0 96.1521
R1077 VN.n14 VN.t5 96.1521
R1078 VN.n40 VN.t7 96.1521
R1079 VN.n53 VN.t1 96.1521
R1080 VN.n82 VN.t8 96.1521
R1081 VN.n69 VN.t4 96.1521
R1082 VN.n95 VN.t3 96.1521
R1083 VN.n108 VN.t2 96.1521
R1084 VN.n14 VN.n13 64.9805
R1085 VN.n69 VN.n68 64.9805
R1086 VN VN.n109 62.9703
R1087 VN.n54 VN.n53 61.7228
R1088 VN.n109 VN.n108 61.7228
R1089 VN.n47 VN.n46 56.5617
R1090 VN.n102 VN.n101 56.5617
R1091 VN.n21 VN.n20 50.7491
R1092 VN.n34 VN.n33 50.7491
R1093 VN.n76 VN.n75 50.7491
R1094 VN.n89 VN.n88 50.7491
R1095 VN.n22 VN.n21 30.405
R1096 VN.n33 VN.n32 30.405
R1097 VN.n77 VN.n76 30.405
R1098 VN.n88 VN.n87 30.405
R1099 VN.n16 VN.n15 24.5923
R1100 VN.n16 VN.n11 24.5923
R1101 VN.n20 VN.n11 24.5923
R1102 VN.n22 VN.n9 24.5923
R1103 VN.n26 VN.n9 24.5923
R1104 VN.n27 VN.n26 24.5923
R1105 VN.n28 VN.n27 24.5923
R1106 VN.n28 VN.n7 24.5923
R1107 VN.n32 VN.n7 24.5923
R1108 VN.n34 VN.n5 24.5923
R1109 VN.n38 VN.n5 24.5923
R1110 VN.n39 VN.n38 24.5923
R1111 VN.n41 VN.n3 24.5923
R1112 VN.n45 VN.n3 24.5923
R1113 VN.n46 VN.n45 24.5923
R1114 VN.n47 VN.n1 24.5923
R1115 VN.n51 VN.n1 24.5923
R1116 VN.n52 VN.n51 24.5923
R1117 VN.n75 VN.n66 24.5923
R1118 VN.n71 VN.n66 24.5923
R1119 VN.n71 VN.n70 24.5923
R1120 VN.n87 VN.n62 24.5923
R1121 VN.n83 VN.n62 24.5923
R1122 VN.n83 VN.n82 24.5923
R1123 VN.n82 VN.n81 24.5923
R1124 VN.n81 VN.n64 24.5923
R1125 VN.n77 VN.n64 24.5923
R1126 VN.n101 VN.n100 24.5923
R1127 VN.n100 VN.n58 24.5923
R1128 VN.n96 VN.n58 24.5923
R1129 VN.n94 VN.n93 24.5923
R1130 VN.n93 VN.n60 24.5923
R1131 VN.n89 VN.n60 24.5923
R1132 VN.n107 VN.n106 24.5923
R1133 VN.n106 VN.n56 24.5923
R1134 VN.n102 VN.n56 24.5923
R1135 VN.n53 VN.n52 20.6576
R1136 VN.n108 VN.n107 20.6576
R1137 VN.n41 VN.n40 14.2638
R1138 VN.n96 VN.n95 14.2638
R1139 VN.n15 VN.n14 10.3291
R1140 VN.n40 VN.n39 10.3291
R1141 VN.n70 VN.n69 10.3291
R1142 VN.n95 VN.n94 10.3291
R1143 VN.n68 VN.n67 2.66364
R1144 VN.n13 VN.n12 2.66364
R1145 VN.n109 VN.n55 0.417304
R1146 VN.n54 VN.n0 0.417304
R1147 VN VN.n54 0.394524
R1148 VN.n105 VN.n55 0.189894
R1149 VN.n105 VN.n104 0.189894
R1150 VN.n104 VN.n103 0.189894
R1151 VN.n103 VN.n57 0.189894
R1152 VN.n99 VN.n57 0.189894
R1153 VN.n99 VN.n98 0.189894
R1154 VN.n98 VN.n97 0.189894
R1155 VN.n97 VN.n59 0.189894
R1156 VN.n92 VN.n59 0.189894
R1157 VN.n92 VN.n91 0.189894
R1158 VN.n91 VN.n90 0.189894
R1159 VN.n90 VN.n61 0.189894
R1160 VN.n86 VN.n61 0.189894
R1161 VN.n86 VN.n85 0.189894
R1162 VN.n85 VN.n84 0.189894
R1163 VN.n84 VN.n63 0.189894
R1164 VN.n80 VN.n63 0.189894
R1165 VN.n80 VN.n79 0.189894
R1166 VN.n79 VN.n78 0.189894
R1167 VN.n78 VN.n65 0.189894
R1168 VN.n74 VN.n65 0.189894
R1169 VN.n74 VN.n73 0.189894
R1170 VN.n73 VN.n72 0.189894
R1171 VN.n72 VN.n67 0.189894
R1172 VN.n17 VN.n12 0.189894
R1173 VN.n18 VN.n17 0.189894
R1174 VN.n19 VN.n18 0.189894
R1175 VN.n19 VN.n10 0.189894
R1176 VN.n23 VN.n10 0.189894
R1177 VN.n24 VN.n23 0.189894
R1178 VN.n25 VN.n24 0.189894
R1179 VN.n25 VN.n8 0.189894
R1180 VN.n29 VN.n8 0.189894
R1181 VN.n30 VN.n29 0.189894
R1182 VN.n31 VN.n30 0.189894
R1183 VN.n31 VN.n6 0.189894
R1184 VN.n35 VN.n6 0.189894
R1185 VN.n36 VN.n35 0.189894
R1186 VN.n37 VN.n36 0.189894
R1187 VN.n37 VN.n4 0.189894
R1188 VN.n42 VN.n4 0.189894
R1189 VN.n43 VN.n42 0.189894
R1190 VN.n44 VN.n43 0.189894
R1191 VN.n44 VN.n2 0.189894
R1192 VN.n48 VN.n2 0.189894
R1193 VN.n49 VN.n48 0.189894
R1194 VN.n50 VN.n49 0.189894
R1195 VN.n50 VN.n0 0.189894
R1196 VDD2.n169 VDD2.n89 756.745
R1197 VDD2.n80 VDD2.n0 756.745
R1198 VDD2.n170 VDD2.n169 585
R1199 VDD2.n168 VDD2.n167 585
R1200 VDD2.n93 VDD2.n92 585
R1201 VDD2.n97 VDD2.n95 585
R1202 VDD2.n162 VDD2.n161 585
R1203 VDD2.n160 VDD2.n159 585
R1204 VDD2.n99 VDD2.n98 585
R1205 VDD2.n154 VDD2.n153 585
R1206 VDD2.n152 VDD2.n151 585
R1207 VDD2.n103 VDD2.n102 585
R1208 VDD2.n146 VDD2.n145 585
R1209 VDD2.n144 VDD2.n143 585
R1210 VDD2.n107 VDD2.n106 585
R1211 VDD2.n138 VDD2.n137 585
R1212 VDD2.n136 VDD2.n135 585
R1213 VDD2.n111 VDD2.n110 585
R1214 VDD2.n130 VDD2.n129 585
R1215 VDD2.n128 VDD2.n127 585
R1216 VDD2.n115 VDD2.n114 585
R1217 VDD2.n122 VDD2.n121 585
R1218 VDD2.n120 VDD2.n119 585
R1219 VDD2.n29 VDD2.n28 585
R1220 VDD2.n31 VDD2.n30 585
R1221 VDD2.n24 VDD2.n23 585
R1222 VDD2.n37 VDD2.n36 585
R1223 VDD2.n39 VDD2.n38 585
R1224 VDD2.n20 VDD2.n19 585
R1225 VDD2.n45 VDD2.n44 585
R1226 VDD2.n47 VDD2.n46 585
R1227 VDD2.n16 VDD2.n15 585
R1228 VDD2.n53 VDD2.n52 585
R1229 VDD2.n55 VDD2.n54 585
R1230 VDD2.n12 VDD2.n11 585
R1231 VDD2.n61 VDD2.n60 585
R1232 VDD2.n63 VDD2.n62 585
R1233 VDD2.n8 VDD2.n7 585
R1234 VDD2.n70 VDD2.n69 585
R1235 VDD2.n71 VDD2.n6 585
R1236 VDD2.n73 VDD2.n72 585
R1237 VDD2.n4 VDD2.n3 585
R1238 VDD2.n79 VDD2.n78 585
R1239 VDD2.n81 VDD2.n80 585
R1240 VDD2.n118 VDD2.t7 327.466
R1241 VDD2.n27 VDD2.t0 327.466
R1242 VDD2.n169 VDD2.n168 171.744
R1243 VDD2.n168 VDD2.n92 171.744
R1244 VDD2.n97 VDD2.n92 171.744
R1245 VDD2.n161 VDD2.n97 171.744
R1246 VDD2.n161 VDD2.n160 171.744
R1247 VDD2.n160 VDD2.n98 171.744
R1248 VDD2.n153 VDD2.n98 171.744
R1249 VDD2.n153 VDD2.n152 171.744
R1250 VDD2.n152 VDD2.n102 171.744
R1251 VDD2.n145 VDD2.n102 171.744
R1252 VDD2.n145 VDD2.n144 171.744
R1253 VDD2.n144 VDD2.n106 171.744
R1254 VDD2.n137 VDD2.n106 171.744
R1255 VDD2.n137 VDD2.n136 171.744
R1256 VDD2.n136 VDD2.n110 171.744
R1257 VDD2.n129 VDD2.n110 171.744
R1258 VDD2.n129 VDD2.n128 171.744
R1259 VDD2.n128 VDD2.n114 171.744
R1260 VDD2.n121 VDD2.n114 171.744
R1261 VDD2.n121 VDD2.n120 171.744
R1262 VDD2.n30 VDD2.n29 171.744
R1263 VDD2.n30 VDD2.n23 171.744
R1264 VDD2.n37 VDD2.n23 171.744
R1265 VDD2.n38 VDD2.n37 171.744
R1266 VDD2.n38 VDD2.n19 171.744
R1267 VDD2.n45 VDD2.n19 171.744
R1268 VDD2.n46 VDD2.n45 171.744
R1269 VDD2.n46 VDD2.n15 171.744
R1270 VDD2.n53 VDD2.n15 171.744
R1271 VDD2.n54 VDD2.n53 171.744
R1272 VDD2.n54 VDD2.n11 171.744
R1273 VDD2.n61 VDD2.n11 171.744
R1274 VDD2.n62 VDD2.n61 171.744
R1275 VDD2.n62 VDD2.n7 171.744
R1276 VDD2.n70 VDD2.n7 171.744
R1277 VDD2.n71 VDD2.n70 171.744
R1278 VDD2.n72 VDD2.n71 171.744
R1279 VDD2.n72 VDD2.n3 171.744
R1280 VDD2.n79 VDD2.n3 171.744
R1281 VDD2.n80 VDD2.n79 171.744
R1282 VDD2.n120 VDD2.t7 85.8723
R1283 VDD2.n29 VDD2.t0 85.8723
R1284 VDD2.n88 VDD2.n87 75.2519
R1285 VDD2 VDD2.n177 75.249
R1286 VDD2.n176 VDD2.n175 72.5854
R1287 VDD2.n86 VDD2.n85 72.5852
R1288 VDD2.n86 VDD2.n84 54.8207
R1289 VDD2.n174 VDD2.n88 54.2993
R1290 VDD2.n174 VDD2.n173 51.1914
R1291 VDD2.n119 VDD2.n118 16.3895
R1292 VDD2.n28 VDD2.n27 16.3895
R1293 VDD2.n95 VDD2.n93 13.1884
R1294 VDD2.n73 VDD2.n4 13.1884
R1295 VDD2.n167 VDD2.n166 12.8005
R1296 VDD2.n163 VDD2.n162 12.8005
R1297 VDD2.n122 VDD2.n117 12.8005
R1298 VDD2.n31 VDD2.n26 12.8005
R1299 VDD2.n74 VDD2.n6 12.8005
R1300 VDD2.n78 VDD2.n77 12.8005
R1301 VDD2.n170 VDD2.n91 12.0247
R1302 VDD2.n159 VDD2.n96 12.0247
R1303 VDD2.n123 VDD2.n115 12.0247
R1304 VDD2.n32 VDD2.n24 12.0247
R1305 VDD2.n69 VDD2.n68 12.0247
R1306 VDD2.n81 VDD2.n2 12.0247
R1307 VDD2.n171 VDD2.n89 11.249
R1308 VDD2.n158 VDD2.n99 11.249
R1309 VDD2.n127 VDD2.n126 11.249
R1310 VDD2.n36 VDD2.n35 11.249
R1311 VDD2.n67 VDD2.n8 11.249
R1312 VDD2.n82 VDD2.n0 11.249
R1313 VDD2.n155 VDD2.n154 10.4732
R1314 VDD2.n130 VDD2.n113 10.4732
R1315 VDD2.n39 VDD2.n22 10.4732
R1316 VDD2.n64 VDD2.n63 10.4732
R1317 VDD2.n151 VDD2.n101 9.69747
R1318 VDD2.n131 VDD2.n111 9.69747
R1319 VDD2.n40 VDD2.n20 9.69747
R1320 VDD2.n60 VDD2.n10 9.69747
R1321 VDD2.n173 VDD2.n172 9.45567
R1322 VDD2.n84 VDD2.n83 9.45567
R1323 VDD2.n105 VDD2.n104 9.3005
R1324 VDD2.n148 VDD2.n147 9.3005
R1325 VDD2.n150 VDD2.n149 9.3005
R1326 VDD2.n101 VDD2.n100 9.3005
R1327 VDD2.n156 VDD2.n155 9.3005
R1328 VDD2.n158 VDD2.n157 9.3005
R1329 VDD2.n96 VDD2.n94 9.3005
R1330 VDD2.n164 VDD2.n163 9.3005
R1331 VDD2.n172 VDD2.n171 9.3005
R1332 VDD2.n91 VDD2.n90 9.3005
R1333 VDD2.n166 VDD2.n165 9.3005
R1334 VDD2.n142 VDD2.n141 9.3005
R1335 VDD2.n140 VDD2.n139 9.3005
R1336 VDD2.n109 VDD2.n108 9.3005
R1337 VDD2.n134 VDD2.n133 9.3005
R1338 VDD2.n132 VDD2.n131 9.3005
R1339 VDD2.n113 VDD2.n112 9.3005
R1340 VDD2.n126 VDD2.n125 9.3005
R1341 VDD2.n124 VDD2.n123 9.3005
R1342 VDD2.n117 VDD2.n116 9.3005
R1343 VDD2.n83 VDD2.n82 9.3005
R1344 VDD2.n2 VDD2.n1 9.3005
R1345 VDD2.n77 VDD2.n76 9.3005
R1346 VDD2.n49 VDD2.n48 9.3005
R1347 VDD2.n18 VDD2.n17 9.3005
R1348 VDD2.n43 VDD2.n42 9.3005
R1349 VDD2.n41 VDD2.n40 9.3005
R1350 VDD2.n22 VDD2.n21 9.3005
R1351 VDD2.n35 VDD2.n34 9.3005
R1352 VDD2.n33 VDD2.n32 9.3005
R1353 VDD2.n26 VDD2.n25 9.3005
R1354 VDD2.n51 VDD2.n50 9.3005
R1355 VDD2.n14 VDD2.n13 9.3005
R1356 VDD2.n57 VDD2.n56 9.3005
R1357 VDD2.n59 VDD2.n58 9.3005
R1358 VDD2.n10 VDD2.n9 9.3005
R1359 VDD2.n65 VDD2.n64 9.3005
R1360 VDD2.n67 VDD2.n66 9.3005
R1361 VDD2.n68 VDD2.n5 9.3005
R1362 VDD2.n75 VDD2.n74 9.3005
R1363 VDD2.n150 VDD2.n103 8.92171
R1364 VDD2.n135 VDD2.n134 8.92171
R1365 VDD2.n44 VDD2.n43 8.92171
R1366 VDD2.n59 VDD2.n12 8.92171
R1367 VDD2.n147 VDD2.n146 8.14595
R1368 VDD2.n138 VDD2.n109 8.14595
R1369 VDD2.n47 VDD2.n18 8.14595
R1370 VDD2.n56 VDD2.n55 8.14595
R1371 VDD2.n143 VDD2.n105 7.3702
R1372 VDD2.n139 VDD2.n107 7.3702
R1373 VDD2.n48 VDD2.n16 7.3702
R1374 VDD2.n52 VDD2.n14 7.3702
R1375 VDD2.n143 VDD2.n142 6.59444
R1376 VDD2.n142 VDD2.n107 6.59444
R1377 VDD2.n51 VDD2.n16 6.59444
R1378 VDD2.n52 VDD2.n51 6.59444
R1379 VDD2.n146 VDD2.n105 5.81868
R1380 VDD2.n139 VDD2.n138 5.81868
R1381 VDD2.n48 VDD2.n47 5.81868
R1382 VDD2.n55 VDD2.n14 5.81868
R1383 VDD2.n147 VDD2.n103 5.04292
R1384 VDD2.n135 VDD2.n109 5.04292
R1385 VDD2.n44 VDD2.n18 5.04292
R1386 VDD2.n56 VDD2.n12 5.04292
R1387 VDD2.n151 VDD2.n150 4.26717
R1388 VDD2.n134 VDD2.n111 4.26717
R1389 VDD2.n43 VDD2.n20 4.26717
R1390 VDD2.n60 VDD2.n59 4.26717
R1391 VDD2.n118 VDD2.n116 3.70982
R1392 VDD2.n27 VDD2.n25 3.70982
R1393 VDD2.n176 VDD2.n174 3.62981
R1394 VDD2.n154 VDD2.n101 3.49141
R1395 VDD2.n131 VDD2.n130 3.49141
R1396 VDD2.n40 VDD2.n39 3.49141
R1397 VDD2.n63 VDD2.n10 3.49141
R1398 VDD2.n173 VDD2.n89 2.71565
R1399 VDD2.n155 VDD2.n99 2.71565
R1400 VDD2.n127 VDD2.n113 2.71565
R1401 VDD2.n36 VDD2.n22 2.71565
R1402 VDD2.n64 VDD2.n8 2.71565
R1403 VDD2.n84 VDD2.n0 2.71565
R1404 VDD2.n177 VDD2.t5 2.10031
R1405 VDD2.n177 VDD2.t3 2.10031
R1406 VDD2.n175 VDD2.t6 2.10031
R1407 VDD2.n175 VDD2.t1 2.10031
R1408 VDD2.n87 VDD2.t2 2.10031
R1409 VDD2.n87 VDD2.t8 2.10031
R1410 VDD2.n85 VDD2.t4 2.10031
R1411 VDD2.n85 VDD2.t9 2.10031
R1412 VDD2.n171 VDD2.n170 1.93989
R1413 VDD2.n159 VDD2.n158 1.93989
R1414 VDD2.n126 VDD2.n115 1.93989
R1415 VDD2.n35 VDD2.n24 1.93989
R1416 VDD2.n69 VDD2.n67 1.93989
R1417 VDD2.n82 VDD2.n81 1.93989
R1418 VDD2.n167 VDD2.n91 1.16414
R1419 VDD2.n162 VDD2.n96 1.16414
R1420 VDD2.n123 VDD2.n122 1.16414
R1421 VDD2.n32 VDD2.n31 1.16414
R1422 VDD2.n68 VDD2.n6 1.16414
R1423 VDD2.n78 VDD2.n2 1.16414
R1424 VDD2 VDD2.n176 0.966017
R1425 VDD2.n88 VDD2.n86 0.852482
R1426 VDD2.n166 VDD2.n93 0.388379
R1427 VDD2.n163 VDD2.n95 0.388379
R1428 VDD2.n119 VDD2.n117 0.388379
R1429 VDD2.n28 VDD2.n26 0.388379
R1430 VDD2.n74 VDD2.n73 0.388379
R1431 VDD2.n77 VDD2.n4 0.388379
R1432 VDD2.n172 VDD2.n90 0.155672
R1433 VDD2.n165 VDD2.n90 0.155672
R1434 VDD2.n165 VDD2.n164 0.155672
R1435 VDD2.n164 VDD2.n94 0.155672
R1436 VDD2.n157 VDD2.n94 0.155672
R1437 VDD2.n157 VDD2.n156 0.155672
R1438 VDD2.n156 VDD2.n100 0.155672
R1439 VDD2.n149 VDD2.n100 0.155672
R1440 VDD2.n149 VDD2.n148 0.155672
R1441 VDD2.n148 VDD2.n104 0.155672
R1442 VDD2.n141 VDD2.n104 0.155672
R1443 VDD2.n141 VDD2.n140 0.155672
R1444 VDD2.n140 VDD2.n108 0.155672
R1445 VDD2.n133 VDD2.n108 0.155672
R1446 VDD2.n133 VDD2.n132 0.155672
R1447 VDD2.n132 VDD2.n112 0.155672
R1448 VDD2.n125 VDD2.n112 0.155672
R1449 VDD2.n125 VDD2.n124 0.155672
R1450 VDD2.n124 VDD2.n116 0.155672
R1451 VDD2.n33 VDD2.n25 0.155672
R1452 VDD2.n34 VDD2.n33 0.155672
R1453 VDD2.n34 VDD2.n21 0.155672
R1454 VDD2.n41 VDD2.n21 0.155672
R1455 VDD2.n42 VDD2.n41 0.155672
R1456 VDD2.n42 VDD2.n17 0.155672
R1457 VDD2.n49 VDD2.n17 0.155672
R1458 VDD2.n50 VDD2.n49 0.155672
R1459 VDD2.n50 VDD2.n13 0.155672
R1460 VDD2.n57 VDD2.n13 0.155672
R1461 VDD2.n58 VDD2.n57 0.155672
R1462 VDD2.n58 VDD2.n9 0.155672
R1463 VDD2.n65 VDD2.n9 0.155672
R1464 VDD2.n66 VDD2.n65 0.155672
R1465 VDD2.n66 VDD2.n5 0.155672
R1466 VDD2.n75 VDD2.n5 0.155672
R1467 VDD2.n76 VDD2.n75 0.155672
R1468 VDD2.n76 VDD2.n1 0.155672
R1469 VDD2.n83 VDD2.n1 0.155672
R1470 B.n580 B.n579 585
R1471 B.n578 B.n187 585
R1472 B.n577 B.n576 585
R1473 B.n575 B.n188 585
R1474 B.n574 B.n573 585
R1475 B.n572 B.n189 585
R1476 B.n571 B.n570 585
R1477 B.n569 B.n190 585
R1478 B.n568 B.n567 585
R1479 B.n566 B.n191 585
R1480 B.n565 B.n564 585
R1481 B.n563 B.n192 585
R1482 B.n562 B.n561 585
R1483 B.n560 B.n193 585
R1484 B.n559 B.n558 585
R1485 B.n557 B.n194 585
R1486 B.n556 B.n555 585
R1487 B.n554 B.n195 585
R1488 B.n553 B.n552 585
R1489 B.n551 B.n196 585
R1490 B.n550 B.n549 585
R1491 B.n548 B.n197 585
R1492 B.n547 B.n546 585
R1493 B.n545 B.n198 585
R1494 B.n544 B.n543 585
R1495 B.n542 B.n199 585
R1496 B.n541 B.n540 585
R1497 B.n539 B.n200 585
R1498 B.n538 B.n537 585
R1499 B.n536 B.n201 585
R1500 B.n535 B.n534 585
R1501 B.n533 B.n202 585
R1502 B.n532 B.n531 585
R1503 B.n530 B.n203 585
R1504 B.n529 B.n528 585
R1505 B.n527 B.n204 585
R1506 B.n526 B.n525 585
R1507 B.n524 B.n205 585
R1508 B.n523 B.n522 585
R1509 B.n521 B.n206 585
R1510 B.n520 B.n519 585
R1511 B.n518 B.n207 585
R1512 B.n517 B.n516 585
R1513 B.n515 B.n208 585
R1514 B.n514 B.n513 585
R1515 B.n512 B.n209 585
R1516 B.n511 B.n510 585
R1517 B.n509 B.n210 585
R1518 B.n508 B.n507 585
R1519 B.n506 B.n211 585
R1520 B.n505 B.n504 585
R1521 B.n503 B.n212 585
R1522 B.n502 B.n501 585
R1523 B.n497 B.n213 585
R1524 B.n496 B.n495 585
R1525 B.n494 B.n214 585
R1526 B.n493 B.n492 585
R1527 B.n491 B.n215 585
R1528 B.n490 B.n489 585
R1529 B.n488 B.n216 585
R1530 B.n487 B.n486 585
R1531 B.n484 B.n217 585
R1532 B.n483 B.n482 585
R1533 B.n481 B.n220 585
R1534 B.n480 B.n479 585
R1535 B.n478 B.n221 585
R1536 B.n477 B.n476 585
R1537 B.n475 B.n222 585
R1538 B.n474 B.n473 585
R1539 B.n472 B.n223 585
R1540 B.n471 B.n470 585
R1541 B.n469 B.n224 585
R1542 B.n468 B.n467 585
R1543 B.n466 B.n225 585
R1544 B.n465 B.n464 585
R1545 B.n463 B.n226 585
R1546 B.n462 B.n461 585
R1547 B.n460 B.n227 585
R1548 B.n459 B.n458 585
R1549 B.n457 B.n228 585
R1550 B.n456 B.n455 585
R1551 B.n454 B.n229 585
R1552 B.n453 B.n452 585
R1553 B.n451 B.n230 585
R1554 B.n450 B.n449 585
R1555 B.n448 B.n231 585
R1556 B.n447 B.n446 585
R1557 B.n445 B.n232 585
R1558 B.n444 B.n443 585
R1559 B.n442 B.n233 585
R1560 B.n441 B.n440 585
R1561 B.n439 B.n234 585
R1562 B.n438 B.n437 585
R1563 B.n436 B.n235 585
R1564 B.n435 B.n434 585
R1565 B.n433 B.n236 585
R1566 B.n432 B.n431 585
R1567 B.n430 B.n237 585
R1568 B.n429 B.n428 585
R1569 B.n427 B.n238 585
R1570 B.n426 B.n425 585
R1571 B.n424 B.n239 585
R1572 B.n423 B.n422 585
R1573 B.n421 B.n240 585
R1574 B.n420 B.n419 585
R1575 B.n418 B.n241 585
R1576 B.n417 B.n416 585
R1577 B.n415 B.n242 585
R1578 B.n414 B.n413 585
R1579 B.n412 B.n243 585
R1580 B.n411 B.n410 585
R1581 B.n409 B.n244 585
R1582 B.n408 B.n407 585
R1583 B.n581 B.n186 585
R1584 B.n583 B.n582 585
R1585 B.n584 B.n185 585
R1586 B.n586 B.n585 585
R1587 B.n587 B.n184 585
R1588 B.n589 B.n588 585
R1589 B.n590 B.n183 585
R1590 B.n592 B.n591 585
R1591 B.n593 B.n182 585
R1592 B.n595 B.n594 585
R1593 B.n596 B.n181 585
R1594 B.n598 B.n597 585
R1595 B.n599 B.n180 585
R1596 B.n601 B.n600 585
R1597 B.n602 B.n179 585
R1598 B.n604 B.n603 585
R1599 B.n605 B.n178 585
R1600 B.n607 B.n606 585
R1601 B.n608 B.n177 585
R1602 B.n610 B.n609 585
R1603 B.n611 B.n176 585
R1604 B.n613 B.n612 585
R1605 B.n614 B.n175 585
R1606 B.n616 B.n615 585
R1607 B.n617 B.n174 585
R1608 B.n619 B.n618 585
R1609 B.n620 B.n173 585
R1610 B.n622 B.n621 585
R1611 B.n623 B.n172 585
R1612 B.n625 B.n624 585
R1613 B.n626 B.n171 585
R1614 B.n628 B.n627 585
R1615 B.n629 B.n170 585
R1616 B.n631 B.n630 585
R1617 B.n632 B.n169 585
R1618 B.n634 B.n633 585
R1619 B.n635 B.n168 585
R1620 B.n637 B.n636 585
R1621 B.n638 B.n167 585
R1622 B.n640 B.n639 585
R1623 B.n641 B.n166 585
R1624 B.n643 B.n642 585
R1625 B.n644 B.n165 585
R1626 B.n646 B.n645 585
R1627 B.n647 B.n164 585
R1628 B.n649 B.n648 585
R1629 B.n650 B.n163 585
R1630 B.n652 B.n651 585
R1631 B.n653 B.n162 585
R1632 B.n655 B.n654 585
R1633 B.n656 B.n161 585
R1634 B.n658 B.n657 585
R1635 B.n659 B.n160 585
R1636 B.n661 B.n660 585
R1637 B.n662 B.n159 585
R1638 B.n664 B.n663 585
R1639 B.n665 B.n158 585
R1640 B.n667 B.n666 585
R1641 B.n668 B.n157 585
R1642 B.n670 B.n669 585
R1643 B.n671 B.n156 585
R1644 B.n673 B.n672 585
R1645 B.n674 B.n155 585
R1646 B.n676 B.n675 585
R1647 B.n677 B.n154 585
R1648 B.n679 B.n678 585
R1649 B.n680 B.n153 585
R1650 B.n682 B.n681 585
R1651 B.n683 B.n152 585
R1652 B.n685 B.n684 585
R1653 B.n686 B.n151 585
R1654 B.n688 B.n687 585
R1655 B.n689 B.n150 585
R1656 B.n691 B.n690 585
R1657 B.n692 B.n149 585
R1658 B.n694 B.n693 585
R1659 B.n695 B.n148 585
R1660 B.n697 B.n696 585
R1661 B.n698 B.n147 585
R1662 B.n700 B.n699 585
R1663 B.n701 B.n146 585
R1664 B.n703 B.n702 585
R1665 B.n704 B.n145 585
R1666 B.n706 B.n705 585
R1667 B.n707 B.n144 585
R1668 B.n709 B.n708 585
R1669 B.n710 B.n143 585
R1670 B.n712 B.n711 585
R1671 B.n713 B.n142 585
R1672 B.n715 B.n714 585
R1673 B.n716 B.n141 585
R1674 B.n718 B.n717 585
R1675 B.n719 B.n140 585
R1676 B.n721 B.n720 585
R1677 B.n722 B.n139 585
R1678 B.n724 B.n723 585
R1679 B.n725 B.n138 585
R1680 B.n727 B.n726 585
R1681 B.n728 B.n137 585
R1682 B.n730 B.n729 585
R1683 B.n731 B.n136 585
R1684 B.n733 B.n732 585
R1685 B.n734 B.n135 585
R1686 B.n736 B.n735 585
R1687 B.n737 B.n134 585
R1688 B.n739 B.n738 585
R1689 B.n740 B.n133 585
R1690 B.n742 B.n741 585
R1691 B.n743 B.n132 585
R1692 B.n745 B.n744 585
R1693 B.n746 B.n131 585
R1694 B.n748 B.n747 585
R1695 B.n749 B.n130 585
R1696 B.n751 B.n750 585
R1697 B.n752 B.n129 585
R1698 B.n754 B.n753 585
R1699 B.n755 B.n128 585
R1700 B.n757 B.n756 585
R1701 B.n758 B.n127 585
R1702 B.n760 B.n759 585
R1703 B.n761 B.n126 585
R1704 B.n763 B.n762 585
R1705 B.n764 B.n125 585
R1706 B.n766 B.n765 585
R1707 B.n767 B.n124 585
R1708 B.n769 B.n768 585
R1709 B.n770 B.n123 585
R1710 B.n772 B.n771 585
R1711 B.n773 B.n122 585
R1712 B.n775 B.n774 585
R1713 B.n776 B.n121 585
R1714 B.n778 B.n777 585
R1715 B.n779 B.n120 585
R1716 B.n781 B.n780 585
R1717 B.n782 B.n119 585
R1718 B.n784 B.n783 585
R1719 B.n785 B.n118 585
R1720 B.n787 B.n786 585
R1721 B.n788 B.n117 585
R1722 B.n790 B.n789 585
R1723 B.n791 B.n116 585
R1724 B.n793 B.n792 585
R1725 B.n794 B.n115 585
R1726 B.n796 B.n795 585
R1727 B.n797 B.n114 585
R1728 B.n799 B.n798 585
R1729 B.n800 B.n113 585
R1730 B.n802 B.n801 585
R1731 B.n803 B.n112 585
R1732 B.n805 B.n804 585
R1733 B.n806 B.n111 585
R1734 B.n808 B.n807 585
R1735 B.n809 B.n110 585
R1736 B.n811 B.n810 585
R1737 B.n812 B.n109 585
R1738 B.n814 B.n813 585
R1739 B.n815 B.n108 585
R1740 B.n817 B.n816 585
R1741 B.n818 B.n107 585
R1742 B.n820 B.n819 585
R1743 B.n821 B.n106 585
R1744 B.n823 B.n822 585
R1745 B.n824 B.n105 585
R1746 B.n826 B.n825 585
R1747 B.n827 B.n104 585
R1748 B.n829 B.n828 585
R1749 B.n1000 B.n43 585
R1750 B.n999 B.n998 585
R1751 B.n997 B.n44 585
R1752 B.n996 B.n995 585
R1753 B.n994 B.n45 585
R1754 B.n993 B.n992 585
R1755 B.n991 B.n46 585
R1756 B.n990 B.n989 585
R1757 B.n988 B.n47 585
R1758 B.n987 B.n986 585
R1759 B.n985 B.n48 585
R1760 B.n984 B.n983 585
R1761 B.n982 B.n49 585
R1762 B.n981 B.n980 585
R1763 B.n979 B.n50 585
R1764 B.n978 B.n977 585
R1765 B.n976 B.n51 585
R1766 B.n975 B.n974 585
R1767 B.n973 B.n52 585
R1768 B.n972 B.n971 585
R1769 B.n970 B.n53 585
R1770 B.n969 B.n968 585
R1771 B.n967 B.n54 585
R1772 B.n966 B.n965 585
R1773 B.n964 B.n55 585
R1774 B.n963 B.n962 585
R1775 B.n961 B.n56 585
R1776 B.n960 B.n959 585
R1777 B.n958 B.n57 585
R1778 B.n957 B.n956 585
R1779 B.n955 B.n58 585
R1780 B.n954 B.n953 585
R1781 B.n952 B.n59 585
R1782 B.n951 B.n950 585
R1783 B.n949 B.n60 585
R1784 B.n948 B.n947 585
R1785 B.n946 B.n61 585
R1786 B.n945 B.n944 585
R1787 B.n943 B.n62 585
R1788 B.n942 B.n941 585
R1789 B.n940 B.n63 585
R1790 B.n939 B.n938 585
R1791 B.n937 B.n64 585
R1792 B.n936 B.n935 585
R1793 B.n934 B.n65 585
R1794 B.n933 B.n932 585
R1795 B.n931 B.n66 585
R1796 B.n930 B.n929 585
R1797 B.n928 B.n67 585
R1798 B.n927 B.n926 585
R1799 B.n925 B.n68 585
R1800 B.n924 B.n923 585
R1801 B.n921 B.n69 585
R1802 B.n920 B.n919 585
R1803 B.n918 B.n72 585
R1804 B.n917 B.n916 585
R1805 B.n915 B.n73 585
R1806 B.n914 B.n913 585
R1807 B.n912 B.n74 585
R1808 B.n911 B.n910 585
R1809 B.n909 B.n75 585
R1810 B.n907 B.n906 585
R1811 B.n905 B.n78 585
R1812 B.n904 B.n903 585
R1813 B.n902 B.n79 585
R1814 B.n901 B.n900 585
R1815 B.n899 B.n80 585
R1816 B.n898 B.n897 585
R1817 B.n896 B.n81 585
R1818 B.n895 B.n894 585
R1819 B.n893 B.n82 585
R1820 B.n892 B.n891 585
R1821 B.n890 B.n83 585
R1822 B.n889 B.n888 585
R1823 B.n887 B.n84 585
R1824 B.n886 B.n885 585
R1825 B.n884 B.n85 585
R1826 B.n883 B.n882 585
R1827 B.n881 B.n86 585
R1828 B.n880 B.n879 585
R1829 B.n878 B.n87 585
R1830 B.n877 B.n876 585
R1831 B.n875 B.n88 585
R1832 B.n874 B.n873 585
R1833 B.n872 B.n89 585
R1834 B.n871 B.n870 585
R1835 B.n869 B.n90 585
R1836 B.n868 B.n867 585
R1837 B.n866 B.n91 585
R1838 B.n865 B.n864 585
R1839 B.n863 B.n92 585
R1840 B.n862 B.n861 585
R1841 B.n860 B.n93 585
R1842 B.n859 B.n858 585
R1843 B.n857 B.n94 585
R1844 B.n856 B.n855 585
R1845 B.n854 B.n95 585
R1846 B.n853 B.n852 585
R1847 B.n851 B.n96 585
R1848 B.n850 B.n849 585
R1849 B.n848 B.n97 585
R1850 B.n847 B.n846 585
R1851 B.n845 B.n98 585
R1852 B.n844 B.n843 585
R1853 B.n842 B.n99 585
R1854 B.n841 B.n840 585
R1855 B.n839 B.n100 585
R1856 B.n838 B.n837 585
R1857 B.n836 B.n101 585
R1858 B.n835 B.n834 585
R1859 B.n833 B.n102 585
R1860 B.n832 B.n831 585
R1861 B.n830 B.n103 585
R1862 B.n1002 B.n1001 585
R1863 B.n1003 B.n42 585
R1864 B.n1005 B.n1004 585
R1865 B.n1006 B.n41 585
R1866 B.n1008 B.n1007 585
R1867 B.n1009 B.n40 585
R1868 B.n1011 B.n1010 585
R1869 B.n1012 B.n39 585
R1870 B.n1014 B.n1013 585
R1871 B.n1015 B.n38 585
R1872 B.n1017 B.n1016 585
R1873 B.n1018 B.n37 585
R1874 B.n1020 B.n1019 585
R1875 B.n1021 B.n36 585
R1876 B.n1023 B.n1022 585
R1877 B.n1024 B.n35 585
R1878 B.n1026 B.n1025 585
R1879 B.n1027 B.n34 585
R1880 B.n1029 B.n1028 585
R1881 B.n1030 B.n33 585
R1882 B.n1032 B.n1031 585
R1883 B.n1033 B.n32 585
R1884 B.n1035 B.n1034 585
R1885 B.n1036 B.n31 585
R1886 B.n1038 B.n1037 585
R1887 B.n1039 B.n30 585
R1888 B.n1041 B.n1040 585
R1889 B.n1042 B.n29 585
R1890 B.n1044 B.n1043 585
R1891 B.n1045 B.n28 585
R1892 B.n1047 B.n1046 585
R1893 B.n1048 B.n27 585
R1894 B.n1050 B.n1049 585
R1895 B.n1051 B.n26 585
R1896 B.n1053 B.n1052 585
R1897 B.n1054 B.n25 585
R1898 B.n1056 B.n1055 585
R1899 B.n1057 B.n24 585
R1900 B.n1059 B.n1058 585
R1901 B.n1060 B.n23 585
R1902 B.n1062 B.n1061 585
R1903 B.n1063 B.n22 585
R1904 B.n1065 B.n1064 585
R1905 B.n1066 B.n21 585
R1906 B.n1068 B.n1067 585
R1907 B.n1069 B.n20 585
R1908 B.n1071 B.n1070 585
R1909 B.n1072 B.n19 585
R1910 B.n1074 B.n1073 585
R1911 B.n1075 B.n18 585
R1912 B.n1077 B.n1076 585
R1913 B.n1078 B.n17 585
R1914 B.n1080 B.n1079 585
R1915 B.n1081 B.n16 585
R1916 B.n1083 B.n1082 585
R1917 B.n1084 B.n15 585
R1918 B.n1086 B.n1085 585
R1919 B.n1087 B.n14 585
R1920 B.n1089 B.n1088 585
R1921 B.n1090 B.n13 585
R1922 B.n1092 B.n1091 585
R1923 B.n1093 B.n12 585
R1924 B.n1095 B.n1094 585
R1925 B.n1096 B.n11 585
R1926 B.n1098 B.n1097 585
R1927 B.n1099 B.n10 585
R1928 B.n1101 B.n1100 585
R1929 B.n1102 B.n9 585
R1930 B.n1104 B.n1103 585
R1931 B.n1105 B.n8 585
R1932 B.n1107 B.n1106 585
R1933 B.n1108 B.n7 585
R1934 B.n1110 B.n1109 585
R1935 B.n1111 B.n6 585
R1936 B.n1113 B.n1112 585
R1937 B.n1114 B.n5 585
R1938 B.n1116 B.n1115 585
R1939 B.n1117 B.n4 585
R1940 B.n1119 B.n1118 585
R1941 B.n1120 B.n3 585
R1942 B.n1122 B.n1121 585
R1943 B.n1123 B.n0 585
R1944 B.n2 B.n1 585
R1945 B.n286 B.n285 585
R1946 B.n288 B.n287 585
R1947 B.n289 B.n284 585
R1948 B.n291 B.n290 585
R1949 B.n292 B.n283 585
R1950 B.n294 B.n293 585
R1951 B.n295 B.n282 585
R1952 B.n297 B.n296 585
R1953 B.n298 B.n281 585
R1954 B.n300 B.n299 585
R1955 B.n301 B.n280 585
R1956 B.n303 B.n302 585
R1957 B.n304 B.n279 585
R1958 B.n306 B.n305 585
R1959 B.n307 B.n278 585
R1960 B.n309 B.n308 585
R1961 B.n310 B.n277 585
R1962 B.n312 B.n311 585
R1963 B.n313 B.n276 585
R1964 B.n315 B.n314 585
R1965 B.n316 B.n275 585
R1966 B.n318 B.n317 585
R1967 B.n319 B.n274 585
R1968 B.n321 B.n320 585
R1969 B.n322 B.n273 585
R1970 B.n324 B.n323 585
R1971 B.n325 B.n272 585
R1972 B.n327 B.n326 585
R1973 B.n328 B.n271 585
R1974 B.n330 B.n329 585
R1975 B.n331 B.n270 585
R1976 B.n333 B.n332 585
R1977 B.n334 B.n269 585
R1978 B.n336 B.n335 585
R1979 B.n337 B.n268 585
R1980 B.n339 B.n338 585
R1981 B.n340 B.n267 585
R1982 B.n342 B.n341 585
R1983 B.n343 B.n266 585
R1984 B.n345 B.n344 585
R1985 B.n346 B.n265 585
R1986 B.n348 B.n347 585
R1987 B.n349 B.n264 585
R1988 B.n351 B.n350 585
R1989 B.n352 B.n263 585
R1990 B.n354 B.n353 585
R1991 B.n355 B.n262 585
R1992 B.n357 B.n356 585
R1993 B.n358 B.n261 585
R1994 B.n360 B.n359 585
R1995 B.n361 B.n260 585
R1996 B.n363 B.n362 585
R1997 B.n364 B.n259 585
R1998 B.n366 B.n365 585
R1999 B.n367 B.n258 585
R2000 B.n369 B.n368 585
R2001 B.n370 B.n257 585
R2002 B.n372 B.n371 585
R2003 B.n373 B.n256 585
R2004 B.n375 B.n374 585
R2005 B.n376 B.n255 585
R2006 B.n378 B.n377 585
R2007 B.n379 B.n254 585
R2008 B.n381 B.n380 585
R2009 B.n382 B.n253 585
R2010 B.n384 B.n383 585
R2011 B.n385 B.n252 585
R2012 B.n387 B.n386 585
R2013 B.n388 B.n251 585
R2014 B.n390 B.n389 585
R2015 B.n391 B.n250 585
R2016 B.n393 B.n392 585
R2017 B.n394 B.n249 585
R2018 B.n396 B.n395 585
R2019 B.n397 B.n248 585
R2020 B.n399 B.n398 585
R2021 B.n400 B.n247 585
R2022 B.n402 B.n401 585
R2023 B.n403 B.n246 585
R2024 B.n405 B.n404 585
R2025 B.n406 B.n245 585
R2026 B.n498 B.t10 519.968
R2027 B.n76 B.t2 519.968
R2028 B.n218 B.t7 519.968
R2029 B.n70 B.t5 519.968
R2030 B.n408 B.n245 506.916
R2031 B.n581 B.n580 506.916
R2032 B.n828 B.n103 506.916
R2033 B.n1002 B.n43 506.916
R2034 B.n499 B.t11 438.32
R2035 B.n77 B.t1 438.32
R2036 B.n219 B.t8 438.32
R2037 B.n71 B.t4 438.32
R2038 B.n218 B.t6 305.557
R2039 B.n498 B.t9 305.557
R2040 B.n76 B.t0 305.557
R2041 B.n70 B.t3 305.557
R2042 B.n1125 B.n1124 256.663
R2043 B.n1124 B.n1123 235.042
R2044 B.n1124 B.n2 235.042
R2045 B.n409 B.n408 163.367
R2046 B.n410 B.n409 163.367
R2047 B.n410 B.n243 163.367
R2048 B.n414 B.n243 163.367
R2049 B.n415 B.n414 163.367
R2050 B.n416 B.n415 163.367
R2051 B.n416 B.n241 163.367
R2052 B.n420 B.n241 163.367
R2053 B.n421 B.n420 163.367
R2054 B.n422 B.n421 163.367
R2055 B.n422 B.n239 163.367
R2056 B.n426 B.n239 163.367
R2057 B.n427 B.n426 163.367
R2058 B.n428 B.n427 163.367
R2059 B.n428 B.n237 163.367
R2060 B.n432 B.n237 163.367
R2061 B.n433 B.n432 163.367
R2062 B.n434 B.n433 163.367
R2063 B.n434 B.n235 163.367
R2064 B.n438 B.n235 163.367
R2065 B.n439 B.n438 163.367
R2066 B.n440 B.n439 163.367
R2067 B.n440 B.n233 163.367
R2068 B.n444 B.n233 163.367
R2069 B.n445 B.n444 163.367
R2070 B.n446 B.n445 163.367
R2071 B.n446 B.n231 163.367
R2072 B.n450 B.n231 163.367
R2073 B.n451 B.n450 163.367
R2074 B.n452 B.n451 163.367
R2075 B.n452 B.n229 163.367
R2076 B.n456 B.n229 163.367
R2077 B.n457 B.n456 163.367
R2078 B.n458 B.n457 163.367
R2079 B.n458 B.n227 163.367
R2080 B.n462 B.n227 163.367
R2081 B.n463 B.n462 163.367
R2082 B.n464 B.n463 163.367
R2083 B.n464 B.n225 163.367
R2084 B.n468 B.n225 163.367
R2085 B.n469 B.n468 163.367
R2086 B.n470 B.n469 163.367
R2087 B.n470 B.n223 163.367
R2088 B.n474 B.n223 163.367
R2089 B.n475 B.n474 163.367
R2090 B.n476 B.n475 163.367
R2091 B.n476 B.n221 163.367
R2092 B.n480 B.n221 163.367
R2093 B.n481 B.n480 163.367
R2094 B.n482 B.n481 163.367
R2095 B.n482 B.n217 163.367
R2096 B.n487 B.n217 163.367
R2097 B.n488 B.n487 163.367
R2098 B.n489 B.n488 163.367
R2099 B.n489 B.n215 163.367
R2100 B.n493 B.n215 163.367
R2101 B.n494 B.n493 163.367
R2102 B.n495 B.n494 163.367
R2103 B.n495 B.n213 163.367
R2104 B.n502 B.n213 163.367
R2105 B.n503 B.n502 163.367
R2106 B.n504 B.n503 163.367
R2107 B.n504 B.n211 163.367
R2108 B.n508 B.n211 163.367
R2109 B.n509 B.n508 163.367
R2110 B.n510 B.n509 163.367
R2111 B.n510 B.n209 163.367
R2112 B.n514 B.n209 163.367
R2113 B.n515 B.n514 163.367
R2114 B.n516 B.n515 163.367
R2115 B.n516 B.n207 163.367
R2116 B.n520 B.n207 163.367
R2117 B.n521 B.n520 163.367
R2118 B.n522 B.n521 163.367
R2119 B.n522 B.n205 163.367
R2120 B.n526 B.n205 163.367
R2121 B.n527 B.n526 163.367
R2122 B.n528 B.n527 163.367
R2123 B.n528 B.n203 163.367
R2124 B.n532 B.n203 163.367
R2125 B.n533 B.n532 163.367
R2126 B.n534 B.n533 163.367
R2127 B.n534 B.n201 163.367
R2128 B.n538 B.n201 163.367
R2129 B.n539 B.n538 163.367
R2130 B.n540 B.n539 163.367
R2131 B.n540 B.n199 163.367
R2132 B.n544 B.n199 163.367
R2133 B.n545 B.n544 163.367
R2134 B.n546 B.n545 163.367
R2135 B.n546 B.n197 163.367
R2136 B.n550 B.n197 163.367
R2137 B.n551 B.n550 163.367
R2138 B.n552 B.n551 163.367
R2139 B.n552 B.n195 163.367
R2140 B.n556 B.n195 163.367
R2141 B.n557 B.n556 163.367
R2142 B.n558 B.n557 163.367
R2143 B.n558 B.n193 163.367
R2144 B.n562 B.n193 163.367
R2145 B.n563 B.n562 163.367
R2146 B.n564 B.n563 163.367
R2147 B.n564 B.n191 163.367
R2148 B.n568 B.n191 163.367
R2149 B.n569 B.n568 163.367
R2150 B.n570 B.n569 163.367
R2151 B.n570 B.n189 163.367
R2152 B.n574 B.n189 163.367
R2153 B.n575 B.n574 163.367
R2154 B.n576 B.n575 163.367
R2155 B.n576 B.n187 163.367
R2156 B.n580 B.n187 163.367
R2157 B.n828 B.n827 163.367
R2158 B.n827 B.n826 163.367
R2159 B.n826 B.n105 163.367
R2160 B.n822 B.n105 163.367
R2161 B.n822 B.n821 163.367
R2162 B.n821 B.n820 163.367
R2163 B.n820 B.n107 163.367
R2164 B.n816 B.n107 163.367
R2165 B.n816 B.n815 163.367
R2166 B.n815 B.n814 163.367
R2167 B.n814 B.n109 163.367
R2168 B.n810 B.n109 163.367
R2169 B.n810 B.n809 163.367
R2170 B.n809 B.n808 163.367
R2171 B.n808 B.n111 163.367
R2172 B.n804 B.n111 163.367
R2173 B.n804 B.n803 163.367
R2174 B.n803 B.n802 163.367
R2175 B.n802 B.n113 163.367
R2176 B.n798 B.n113 163.367
R2177 B.n798 B.n797 163.367
R2178 B.n797 B.n796 163.367
R2179 B.n796 B.n115 163.367
R2180 B.n792 B.n115 163.367
R2181 B.n792 B.n791 163.367
R2182 B.n791 B.n790 163.367
R2183 B.n790 B.n117 163.367
R2184 B.n786 B.n117 163.367
R2185 B.n786 B.n785 163.367
R2186 B.n785 B.n784 163.367
R2187 B.n784 B.n119 163.367
R2188 B.n780 B.n119 163.367
R2189 B.n780 B.n779 163.367
R2190 B.n779 B.n778 163.367
R2191 B.n778 B.n121 163.367
R2192 B.n774 B.n121 163.367
R2193 B.n774 B.n773 163.367
R2194 B.n773 B.n772 163.367
R2195 B.n772 B.n123 163.367
R2196 B.n768 B.n123 163.367
R2197 B.n768 B.n767 163.367
R2198 B.n767 B.n766 163.367
R2199 B.n766 B.n125 163.367
R2200 B.n762 B.n125 163.367
R2201 B.n762 B.n761 163.367
R2202 B.n761 B.n760 163.367
R2203 B.n760 B.n127 163.367
R2204 B.n756 B.n127 163.367
R2205 B.n756 B.n755 163.367
R2206 B.n755 B.n754 163.367
R2207 B.n754 B.n129 163.367
R2208 B.n750 B.n129 163.367
R2209 B.n750 B.n749 163.367
R2210 B.n749 B.n748 163.367
R2211 B.n748 B.n131 163.367
R2212 B.n744 B.n131 163.367
R2213 B.n744 B.n743 163.367
R2214 B.n743 B.n742 163.367
R2215 B.n742 B.n133 163.367
R2216 B.n738 B.n133 163.367
R2217 B.n738 B.n737 163.367
R2218 B.n737 B.n736 163.367
R2219 B.n736 B.n135 163.367
R2220 B.n732 B.n135 163.367
R2221 B.n732 B.n731 163.367
R2222 B.n731 B.n730 163.367
R2223 B.n730 B.n137 163.367
R2224 B.n726 B.n137 163.367
R2225 B.n726 B.n725 163.367
R2226 B.n725 B.n724 163.367
R2227 B.n724 B.n139 163.367
R2228 B.n720 B.n139 163.367
R2229 B.n720 B.n719 163.367
R2230 B.n719 B.n718 163.367
R2231 B.n718 B.n141 163.367
R2232 B.n714 B.n141 163.367
R2233 B.n714 B.n713 163.367
R2234 B.n713 B.n712 163.367
R2235 B.n712 B.n143 163.367
R2236 B.n708 B.n143 163.367
R2237 B.n708 B.n707 163.367
R2238 B.n707 B.n706 163.367
R2239 B.n706 B.n145 163.367
R2240 B.n702 B.n145 163.367
R2241 B.n702 B.n701 163.367
R2242 B.n701 B.n700 163.367
R2243 B.n700 B.n147 163.367
R2244 B.n696 B.n147 163.367
R2245 B.n696 B.n695 163.367
R2246 B.n695 B.n694 163.367
R2247 B.n694 B.n149 163.367
R2248 B.n690 B.n149 163.367
R2249 B.n690 B.n689 163.367
R2250 B.n689 B.n688 163.367
R2251 B.n688 B.n151 163.367
R2252 B.n684 B.n151 163.367
R2253 B.n684 B.n683 163.367
R2254 B.n683 B.n682 163.367
R2255 B.n682 B.n153 163.367
R2256 B.n678 B.n153 163.367
R2257 B.n678 B.n677 163.367
R2258 B.n677 B.n676 163.367
R2259 B.n676 B.n155 163.367
R2260 B.n672 B.n155 163.367
R2261 B.n672 B.n671 163.367
R2262 B.n671 B.n670 163.367
R2263 B.n670 B.n157 163.367
R2264 B.n666 B.n157 163.367
R2265 B.n666 B.n665 163.367
R2266 B.n665 B.n664 163.367
R2267 B.n664 B.n159 163.367
R2268 B.n660 B.n159 163.367
R2269 B.n660 B.n659 163.367
R2270 B.n659 B.n658 163.367
R2271 B.n658 B.n161 163.367
R2272 B.n654 B.n161 163.367
R2273 B.n654 B.n653 163.367
R2274 B.n653 B.n652 163.367
R2275 B.n652 B.n163 163.367
R2276 B.n648 B.n163 163.367
R2277 B.n648 B.n647 163.367
R2278 B.n647 B.n646 163.367
R2279 B.n646 B.n165 163.367
R2280 B.n642 B.n165 163.367
R2281 B.n642 B.n641 163.367
R2282 B.n641 B.n640 163.367
R2283 B.n640 B.n167 163.367
R2284 B.n636 B.n167 163.367
R2285 B.n636 B.n635 163.367
R2286 B.n635 B.n634 163.367
R2287 B.n634 B.n169 163.367
R2288 B.n630 B.n169 163.367
R2289 B.n630 B.n629 163.367
R2290 B.n629 B.n628 163.367
R2291 B.n628 B.n171 163.367
R2292 B.n624 B.n171 163.367
R2293 B.n624 B.n623 163.367
R2294 B.n623 B.n622 163.367
R2295 B.n622 B.n173 163.367
R2296 B.n618 B.n173 163.367
R2297 B.n618 B.n617 163.367
R2298 B.n617 B.n616 163.367
R2299 B.n616 B.n175 163.367
R2300 B.n612 B.n175 163.367
R2301 B.n612 B.n611 163.367
R2302 B.n611 B.n610 163.367
R2303 B.n610 B.n177 163.367
R2304 B.n606 B.n177 163.367
R2305 B.n606 B.n605 163.367
R2306 B.n605 B.n604 163.367
R2307 B.n604 B.n179 163.367
R2308 B.n600 B.n179 163.367
R2309 B.n600 B.n599 163.367
R2310 B.n599 B.n598 163.367
R2311 B.n598 B.n181 163.367
R2312 B.n594 B.n181 163.367
R2313 B.n594 B.n593 163.367
R2314 B.n593 B.n592 163.367
R2315 B.n592 B.n183 163.367
R2316 B.n588 B.n183 163.367
R2317 B.n588 B.n587 163.367
R2318 B.n587 B.n586 163.367
R2319 B.n586 B.n185 163.367
R2320 B.n582 B.n185 163.367
R2321 B.n582 B.n581 163.367
R2322 B.n998 B.n43 163.367
R2323 B.n998 B.n997 163.367
R2324 B.n997 B.n996 163.367
R2325 B.n996 B.n45 163.367
R2326 B.n992 B.n45 163.367
R2327 B.n992 B.n991 163.367
R2328 B.n991 B.n990 163.367
R2329 B.n990 B.n47 163.367
R2330 B.n986 B.n47 163.367
R2331 B.n986 B.n985 163.367
R2332 B.n985 B.n984 163.367
R2333 B.n984 B.n49 163.367
R2334 B.n980 B.n49 163.367
R2335 B.n980 B.n979 163.367
R2336 B.n979 B.n978 163.367
R2337 B.n978 B.n51 163.367
R2338 B.n974 B.n51 163.367
R2339 B.n974 B.n973 163.367
R2340 B.n973 B.n972 163.367
R2341 B.n972 B.n53 163.367
R2342 B.n968 B.n53 163.367
R2343 B.n968 B.n967 163.367
R2344 B.n967 B.n966 163.367
R2345 B.n966 B.n55 163.367
R2346 B.n962 B.n55 163.367
R2347 B.n962 B.n961 163.367
R2348 B.n961 B.n960 163.367
R2349 B.n960 B.n57 163.367
R2350 B.n956 B.n57 163.367
R2351 B.n956 B.n955 163.367
R2352 B.n955 B.n954 163.367
R2353 B.n954 B.n59 163.367
R2354 B.n950 B.n59 163.367
R2355 B.n950 B.n949 163.367
R2356 B.n949 B.n948 163.367
R2357 B.n948 B.n61 163.367
R2358 B.n944 B.n61 163.367
R2359 B.n944 B.n943 163.367
R2360 B.n943 B.n942 163.367
R2361 B.n942 B.n63 163.367
R2362 B.n938 B.n63 163.367
R2363 B.n938 B.n937 163.367
R2364 B.n937 B.n936 163.367
R2365 B.n936 B.n65 163.367
R2366 B.n932 B.n65 163.367
R2367 B.n932 B.n931 163.367
R2368 B.n931 B.n930 163.367
R2369 B.n930 B.n67 163.367
R2370 B.n926 B.n67 163.367
R2371 B.n926 B.n925 163.367
R2372 B.n925 B.n924 163.367
R2373 B.n924 B.n69 163.367
R2374 B.n919 B.n69 163.367
R2375 B.n919 B.n918 163.367
R2376 B.n918 B.n917 163.367
R2377 B.n917 B.n73 163.367
R2378 B.n913 B.n73 163.367
R2379 B.n913 B.n912 163.367
R2380 B.n912 B.n911 163.367
R2381 B.n911 B.n75 163.367
R2382 B.n906 B.n75 163.367
R2383 B.n906 B.n905 163.367
R2384 B.n905 B.n904 163.367
R2385 B.n904 B.n79 163.367
R2386 B.n900 B.n79 163.367
R2387 B.n900 B.n899 163.367
R2388 B.n899 B.n898 163.367
R2389 B.n898 B.n81 163.367
R2390 B.n894 B.n81 163.367
R2391 B.n894 B.n893 163.367
R2392 B.n893 B.n892 163.367
R2393 B.n892 B.n83 163.367
R2394 B.n888 B.n83 163.367
R2395 B.n888 B.n887 163.367
R2396 B.n887 B.n886 163.367
R2397 B.n886 B.n85 163.367
R2398 B.n882 B.n85 163.367
R2399 B.n882 B.n881 163.367
R2400 B.n881 B.n880 163.367
R2401 B.n880 B.n87 163.367
R2402 B.n876 B.n87 163.367
R2403 B.n876 B.n875 163.367
R2404 B.n875 B.n874 163.367
R2405 B.n874 B.n89 163.367
R2406 B.n870 B.n89 163.367
R2407 B.n870 B.n869 163.367
R2408 B.n869 B.n868 163.367
R2409 B.n868 B.n91 163.367
R2410 B.n864 B.n91 163.367
R2411 B.n864 B.n863 163.367
R2412 B.n863 B.n862 163.367
R2413 B.n862 B.n93 163.367
R2414 B.n858 B.n93 163.367
R2415 B.n858 B.n857 163.367
R2416 B.n857 B.n856 163.367
R2417 B.n856 B.n95 163.367
R2418 B.n852 B.n95 163.367
R2419 B.n852 B.n851 163.367
R2420 B.n851 B.n850 163.367
R2421 B.n850 B.n97 163.367
R2422 B.n846 B.n97 163.367
R2423 B.n846 B.n845 163.367
R2424 B.n845 B.n844 163.367
R2425 B.n844 B.n99 163.367
R2426 B.n840 B.n99 163.367
R2427 B.n840 B.n839 163.367
R2428 B.n839 B.n838 163.367
R2429 B.n838 B.n101 163.367
R2430 B.n834 B.n101 163.367
R2431 B.n834 B.n833 163.367
R2432 B.n833 B.n832 163.367
R2433 B.n832 B.n103 163.367
R2434 B.n1003 B.n1002 163.367
R2435 B.n1004 B.n1003 163.367
R2436 B.n1004 B.n41 163.367
R2437 B.n1008 B.n41 163.367
R2438 B.n1009 B.n1008 163.367
R2439 B.n1010 B.n1009 163.367
R2440 B.n1010 B.n39 163.367
R2441 B.n1014 B.n39 163.367
R2442 B.n1015 B.n1014 163.367
R2443 B.n1016 B.n1015 163.367
R2444 B.n1016 B.n37 163.367
R2445 B.n1020 B.n37 163.367
R2446 B.n1021 B.n1020 163.367
R2447 B.n1022 B.n1021 163.367
R2448 B.n1022 B.n35 163.367
R2449 B.n1026 B.n35 163.367
R2450 B.n1027 B.n1026 163.367
R2451 B.n1028 B.n1027 163.367
R2452 B.n1028 B.n33 163.367
R2453 B.n1032 B.n33 163.367
R2454 B.n1033 B.n1032 163.367
R2455 B.n1034 B.n1033 163.367
R2456 B.n1034 B.n31 163.367
R2457 B.n1038 B.n31 163.367
R2458 B.n1039 B.n1038 163.367
R2459 B.n1040 B.n1039 163.367
R2460 B.n1040 B.n29 163.367
R2461 B.n1044 B.n29 163.367
R2462 B.n1045 B.n1044 163.367
R2463 B.n1046 B.n1045 163.367
R2464 B.n1046 B.n27 163.367
R2465 B.n1050 B.n27 163.367
R2466 B.n1051 B.n1050 163.367
R2467 B.n1052 B.n1051 163.367
R2468 B.n1052 B.n25 163.367
R2469 B.n1056 B.n25 163.367
R2470 B.n1057 B.n1056 163.367
R2471 B.n1058 B.n1057 163.367
R2472 B.n1058 B.n23 163.367
R2473 B.n1062 B.n23 163.367
R2474 B.n1063 B.n1062 163.367
R2475 B.n1064 B.n1063 163.367
R2476 B.n1064 B.n21 163.367
R2477 B.n1068 B.n21 163.367
R2478 B.n1069 B.n1068 163.367
R2479 B.n1070 B.n1069 163.367
R2480 B.n1070 B.n19 163.367
R2481 B.n1074 B.n19 163.367
R2482 B.n1075 B.n1074 163.367
R2483 B.n1076 B.n1075 163.367
R2484 B.n1076 B.n17 163.367
R2485 B.n1080 B.n17 163.367
R2486 B.n1081 B.n1080 163.367
R2487 B.n1082 B.n1081 163.367
R2488 B.n1082 B.n15 163.367
R2489 B.n1086 B.n15 163.367
R2490 B.n1087 B.n1086 163.367
R2491 B.n1088 B.n1087 163.367
R2492 B.n1088 B.n13 163.367
R2493 B.n1092 B.n13 163.367
R2494 B.n1093 B.n1092 163.367
R2495 B.n1094 B.n1093 163.367
R2496 B.n1094 B.n11 163.367
R2497 B.n1098 B.n11 163.367
R2498 B.n1099 B.n1098 163.367
R2499 B.n1100 B.n1099 163.367
R2500 B.n1100 B.n9 163.367
R2501 B.n1104 B.n9 163.367
R2502 B.n1105 B.n1104 163.367
R2503 B.n1106 B.n1105 163.367
R2504 B.n1106 B.n7 163.367
R2505 B.n1110 B.n7 163.367
R2506 B.n1111 B.n1110 163.367
R2507 B.n1112 B.n1111 163.367
R2508 B.n1112 B.n5 163.367
R2509 B.n1116 B.n5 163.367
R2510 B.n1117 B.n1116 163.367
R2511 B.n1118 B.n1117 163.367
R2512 B.n1118 B.n3 163.367
R2513 B.n1122 B.n3 163.367
R2514 B.n1123 B.n1122 163.367
R2515 B.n285 B.n2 163.367
R2516 B.n288 B.n285 163.367
R2517 B.n289 B.n288 163.367
R2518 B.n290 B.n289 163.367
R2519 B.n290 B.n283 163.367
R2520 B.n294 B.n283 163.367
R2521 B.n295 B.n294 163.367
R2522 B.n296 B.n295 163.367
R2523 B.n296 B.n281 163.367
R2524 B.n300 B.n281 163.367
R2525 B.n301 B.n300 163.367
R2526 B.n302 B.n301 163.367
R2527 B.n302 B.n279 163.367
R2528 B.n306 B.n279 163.367
R2529 B.n307 B.n306 163.367
R2530 B.n308 B.n307 163.367
R2531 B.n308 B.n277 163.367
R2532 B.n312 B.n277 163.367
R2533 B.n313 B.n312 163.367
R2534 B.n314 B.n313 163.367
R2535 B.n314 B.n275 163.367
R2536 B.n318 B.n275 163.367
R2537 B.n319 B.n318 163.367
R2538 B.n320 B.n319 163.367
R2539 B.n320 B.n273 163.367
R2540 B.n324 B.n273 163.367
R2541 B.n325 B.n324 163.367
R2542 B.n326 B.n325 163.367
R2543 B.n326 B.n271 163.367
R2544 B.n330 B.n271 163.367
R2545 B.n331 B.n330 163.367
R2546 B.n332 B.n331 163.367
R2547 B.n332 B.n269 163.367
R2548 B.n336 B.n269 163.367
R2549 B.n337 B.n336 163.367
R2550 B.n338 B.n337 163.367
R2551 B.n338 B.n267 163.367
R2552 B.n342 B.n267 163.367
R2553 B.n343 B.n342 163.367
R2554 B.n344 B.n343 163.367
R2555 B.n344 B.n265 163.367
R2556 B.n348 B.n265 163.367
R2557 B.n349 B.n348 163.367
R2558 B.n350 B.n349 163.367
R2559 B.n350 B.n263 163.367
R2560 B.n354 B.n263 163.367
R2561 B.n355 B.n354 163.367
R2562 B.n356 B.n355 163.367
R2563 B.n356 B.n261 163.367
R2564 B.n360 B.n261 163.367
R2565 B.n361 B.n360 163.367
R2566 B.n362 B.n361 163.367
R2567 B.n362 B.n259 163.367
R2568 B.n366 B.n259 163.367
R2569 B.n367 B.n366 163.367
R2570 B.n368 B.n367 163.367
R2571 B.n368 B.n257 163.367
R2572 B.n372 B.n257 163.367
R2573 B.n373 B.n372 163.367
R2574 B.n374 B.n373 163.367
R2575 B.n374 B.n255 163.367
R2576 B.n378 B.n255 163.367
R2577 B.n379 B.n378 163.367
R2578 B.n380 B.n379 163.367
R2579 B.n380 B.n253 163.367
R2580 B.n384 B.n253 163.367
R2581 B.n385 B.n384 163.367
R2582 B.n386 B.n385 163.367
R2583 B.n386 B.n251 163.367
R2584 B.n390 B.n251 163.367
R2585 B.n391 B.n390 163.367
R2586 B.n392 B.n391 163.367
R2587 B.n392 B.n249 163.367
R2588 B.n396 B.n249 163.367
R2589 B.n397 B.n396 163.367
R2590 B.n398 B.n397 163.367
R2591 B.n398 B.n247 163.367
R2592 B.n402 B.n247 163.367
R2593 B.n403 B.n402 163.367
R2594 B.n404 B.n403 163.367
R2595 B.n404 B.n245 163.367
R2596 B.n219 B.n218 81.649
R2597 B.n499 B.n498 81.649
R2598 B.n77 B.n76 81.649
R2599 B.n71 B.n70 81.649
R2600 B.n485 B.n219 59.5399
R2601 B.n500 B.n499 59.5399
R2602 B.n908 B.n77 59.5399
R2603 B.n922 B.n71 59.5399
R2604 B.n1001 B.n1000 32.9371
R2605 B.n830 B.n829 32.9371
R2606 B.n579 B.n186 32.9371
R2607 B.n407 B.n406 32.9371
R2608 B B.n1125 18.0485
R2609 B.n1001 B.n42 10.6151
R2610 B.n1005 B.n42 10.6151
R2611 B.n1006 B.n1005 10.6151
R2612 B.n1007 B.n1006 10.6151
R2613 B.n1007 B.n40 10.6151
R2614 B.n1011 B.n40 10.6151
R2615 B.n1012 B.n1011 10.6151
R2616 B.n1013 B.n1012 10.6151
R2617 B.n1013 B.n38 10.6151
R2618 B.n1017 B.n38 10.6151
R2619 B.n1018 B.n1017 10.6151
R2620 B.n1019 B.n1018 10.6151
R2621 B.n1019 B.n36 10.6151
R2622 B.n1023 B.n36 10.6151
R2623 B.n1024 B.n1023 10.6151
R2624 B.n1025 B.n1024 10.6151
R2625 B.n1025 B.n34 10.6151
R2626 B.n1029 B.n34 10.6151
R2627 B.n1030 B.n1029 10.6151
R2628 B.n1031 B.n1030 10.6151
R2629 B.n1031 B.n32 10.6151
R2630 B.n1035 B.n32 10.6151
R2631 B.n1036 B.n1035 10.6151
R2632 B.n1037 B.n1036 10.6151
R2633 B.n1037 B.n30 10.6151
R2634 B.n1041 B.n30 10.6151
R2635 B.n1042 B.n1041 10.6151
R2636 B.n1043 B.n1042 10.6151
R2637 B.n1043 B.n28 10.6151
R2638 B.n1047 B.n28 10.6151
R2639 B.n1048 B.n1047 10.6151
R2640 B.n1049 B.n1048 10.6151
R2641 B.n1049 B.n26 10.6151
R2642 B.n1053 B.n26 10.6151
R2643 B.n1054 B.n1053 10.6151
R2644 B.n1055 B.n1054 10.6151
R2645 B.n1055 B.n24 10.6151
R2646 B.n1059 B.n24 10.6151
R2647 B.n1060 B.n1059 10.6151
R2648 B.n1061 B.n1060 10.6151
R2649 B.n1061 B.n22 10.6151
R2650 B.n1065 B.n22 10.6151
R2651 B.n1066 B.n1065 10.6151
R2652 B.n1067 B.n1066 10.6151
R2653 B.n1067 B.n20 10.6151
R2654 B.n1071 B.n20 10.6151
R2655 B.n1072 B.n1071 10.6151
R2656 B.n1073 B.n1072 10.6151
R2657 B.n1073 B.n18 10.6151
R2658 B.n1077 B.n18 10.6151
R2659 B.n1078 B.n1077 10.6151
R2660 B.n1079 B.n1078 10.6151
R2661 B.n1079 B.n16 10.6151
R2662 B.n1083 B.n16 10.6151
R2663 B.n1084 B.n1083 10.6151
R2664 B.n1085 B.n1084 10.6151
R2665 B.n1085 B.n14 10.6151
R2666 B.n1089 B.n14 10.6151
R2667 B.n1090 B.n1089 10.6151
R2668 B.n1091 B.n1090 10.6151
R2669 B.n1091 B.n12 10.6151
R2670 B.n1095 B.n12 10.6151
R2671 B.n1096 B.n1095 10.6151
R2672 B.n1097 B.n1096 10.6151
R2673 B.n1097 B.n10 10.6151
R2674 B.n1101 B.n10 10.6151
R2675 B.n1102 B.n1101 10.6151
R2676 B.n1103 B.n1102 10.6151
R2677 B.n1103 B.n8 10.6151
R2678 B.n1107 B.n8 10.6151
R2679 B.n1108 B.n1107 10.6151
R2680 B.n1109 B.n1108 10.6151
R2681 B.n1109 B.n6 10.6151
R2682 B.n1113 B.n6 10.6151
R2683 B.n1114 B.n1113 10.6151
R2684 B.n1115 B.n1114 10.6151
R2685 B.n1115 B.n4 10.6151
R2686 B.n1119 B.n4 10.6151
R2687 B.n1120 B.n1119 10.6151
R2688 B.n1121 B.n1120 10.6151
R2689 B.n1121 B.n0 10.6151
R2690 B.n1000 B.n999 10.6151
R2691 B.n999 B.n44 10.6151
R2692 B.n995 B.n44 10.6151
R2693 B.n995 B.n994 10.6151
R2694 B.n994 B.n993 10.6151
R2695 B.n993 B.n46 10.6151
R2696 B.n989 B.n46 10.6151
R2697 B.n989 B.n988 10.6151
R2698 B.n988 B.n987 10.6151
R2699 B.n987 B.n48 10.6151
R2700 B.n983 B.n48 10.6151
R2701 B.n983 B.n982 10.6151
R2702 B.n982 B.n981 10.6151
R2703 B.n981 B.n50 10.6151
R2704 B.n977 B.n50 10.6151
R2705 B.n977 B.n976 10.6151
R2706 B.n976 B.n975 10.6151
R2707 B.n975 B.n52 10.6151
R2708 B.n971 B.n52 10.6151
R2709 B.n971 B.n970 10.6151
R2710 B.n970 B.n969 10.6151
R2711 B.n969 B.n54 10.6151
R2712 B.n965 B.n54 10.6151
R2713 B.n965 B.n964 10.6151
R2714 B.n964 B.n963 10.6151
R2715 B.n963 B.n56 10.6151
R2716 B.n959 B.n56 10.6151
R2717 B.n959 B.n958 10.6151
R2718 B.n958 B.n957 10.6151
R2719 B.n957 B.n58 10.6151
R2720 B.n953 B.n58 10.6151
R2721 B.n953 B.n952 10.6151
R2722 B.n952 B.n951 10.6151
R2723 B.n951 B.n60 10.6151
R2724 B.n947 B.n60 10.6151
R2725 B.n947 B.n946 10.6151
R2726 B.n946 B.n945 10.6151
R2727 B.n945 B.n62 10.6151
R2728 B.n941 B.n62 10.6151
R2729 B.n941 B.n940 10.6151
R2730 B.n940 B.n939 10.6151
R2731 B.n939 B.n64 10.6151
R2732 B.n935 B.n64 10.6151
R2733 B.n935 B.n934 10.6151
R2734 B.n934 B.n933 10.6151
R2735 B.n933 B.n66 10.6151
R2736 B.n929 B.n66 10.6151
R2737 B.n929 B.n928 10.6151
R2738 B.n928 B.n927 10.6151
R2739 B.n927 B.n68 10.6151
R2740 B.n923 B.n68 10.6151
R2741 B.n921 B.n920 10.6151
R2742 B.n920 B.n72 10.6151
R2743 B.n916 B.n72 10.6151
R2744 B.n916 B.n915 10.6151
R2745 B.n915 B.n914 10.6151
R2746 B.n914 B.n74 10.6151
R2747 B.n910 B.n74 10.6151
R2748 B.n910 B.n909 10.6151
R2749 B.n907 B.n78 10.6151
R2750 B.n903 B.n78 10.6151
R2751 B.n903 B.n902 10.6151
R2752 B.n902 B.n901 10.6151
R2753 B.n901 B.n80 10.6151
R2754 B.n897 B.n80 10.6151
R2755 B.n897 B.n896 10.6151
R2756 B.n896 B.n895 10.6151
R2757 B.n895 B.n82 10.6151
R2758 B.n891 B.n82 10.6151
R2759 B.n891 B.n890 10.6151
R2760 B.n890 B.n889 10.6151
R2761 B.n889 B.n84 10.6151
R2762 B.n885 B.n84 10.6151
R2763 B.n885 B.n884 10.6151
R2764 B.n884 B.n883 10.6151
R2765 B.n883 B.n86 10.6151
R2766 B.n879 B.n86 10.6151
R2767 B.n879 B.n878 10.6151
R2768 B.n878 B.n877 10.6151
R2769 B.n877 B.n88 10.6151
R2770 B.n873 B.n88 10.6151
R2771 B.n873 B.n872 10.6151
R2772 B.n872 B.n871 10.6151
R2773 B.n871 B.n90 10.6151
R2774 B.n867 B.n90 10.6151
R2775 B.n867 B.n866 10.6151
R2776 B.n866 B.n865 10.6151
R2777 B.n865 B.n92 10.6151
R2778 B.n861 B.n92 10.6151
R2779 B.n861 B.n860 10.6151
R2780 B.n860 B.n859 10.6151
R2781 B.n859 B.n94 10.6151
R2782 B.n855 B.n94 10.6151
R2783 B.n855 B.n854 10.6151
R2784 B.n854 B.n853 10.6151
R2785 B.n853 B.n96 10.6151
R2786 B.n849 B.n96 10.6151
R2787 B.n849 B.n848 10.6151
R2788 B.n848 B.n847 10.6151
R2789 B.n847 B.n98 10.6151
R2790 B.n843 B.n98 10.6151
R2791 B.n843 B.n842 10.6151
R2792 B.n842 B.n841 10.6151
R2793 B.n841 B.n100 10.6151
R2794 B.n837 B.n100 10.6151
R2795 B.n837 B.n836 10.6151
R2796 B.n836 B.n835 10.6151
R2797 B.n835 B.n102 10.6151
R2798 B.n831 B.n102 10.6151
R2799 B.n831 B.n830 10.6151
R2800 B.n829 B.n104 10.6151
R2801 B.n825 B.n104 10.6151
R2802 B.n825 B.n824 10.6151
R2803 B.n824 B.n823 10.6151
R2804 B.n823 B.n106 10.6151
R2805 B.n819 B.n106 10.6151
R2806 B.n819 B.n818 10.6151
R2807 B.n818 B.n817 10.6151
R2808 B.n817 B.n108 10.6151
R2809 B.n813 B.n108 10.6151
R2810 B.n813 B.n812 10.6151
R2811 B.n812 B.n811 10.6151
R2812 B.n811 B.n110 10.6151
R2813 B.n807 B.n110 10.6151
R2814 B.n807 B.n806 10.6151
R2815 B.n806 B.n805 10.6151
R2816 B.n805 B.n112 10.6151
R2817 B.n801 B.n112 10.6151
R2818 B.n801 B.n800 10.6151
R2819 B.n800 B.n799 10.6151
R2820 B.n799 B.n114 10.6151
R2821 B.n795 B.n114 10.6151
R2822 B.n795 B.n794 10.6151
R2823 B.n794 B.n793 10.6151
R2824 B.n793 B.n116 10.6151
R2825 B.n789 B.n116 10.6151
R2826 B.n789 B.n788 10.6151
R2827 B.n788 B.n787 10.6151
R2828 B.n787 B.n118 10.6151
R2829 B.n783 B.n118 10.6151
R2830 B.n783 B.n782 10.6151
R2831 B.n782 B.n781 10.6151
R2832 B.n781 B.n120 10.6151
R2833 B.n777 B.n120 10.6151
R2834 B.n777 B.n776 10.6151
R2835 B.n776 B.n775 10.6151
R2836 B.n775 B.n122 10.6151
R2837 B.n771 B.n122 10.6151
R2838 B.n771 B.n770 10.6151
R2839 B.n770 B.n769 10.6151
R2840 B.n769 B.n124 10.6151
R2841 B.n765 B.n124 10.6151
R2842 B.n765 B.n764 10.6151
R2843 B.n764 B.n763 10.6151
R2844 B.n763 B.n126 10.6151
R2845 B.n759 B.n126 10.6151
R2846 B.n759 B.n758 10.6151
R2847 B.n758 B.n757 10.6151
R2848 B.n757 B.n128 10.6151
R2849 B.n753 B.n128 10.6151
R2850 B.n753 B.n752 10.6151
R2851 B.n752 B.n751 10.6151
R2852 B.n751 B.n130 10.6151
R2853 B.n747 B.n130 10.6151
R2854 B.n747 B.n746 10.6151
R2855 B.n746 B.n745 10.6151
R2856 B.n745 B.n132 10.6151
R2857 B.n741 B.n132 10.6151
R2858 B.n741 B.n740 10.6151
R2859 B.n740 B.n739 10.6151
R2860 B.n739 B.n134 10.6151
R2861 B.n735 B.n134 10.6151
R2862 B.n735 B.n734 10.6151
R2863 B.n734 B.n733 10.6151
R2864 B.n733 B.n136 10.6151
R2865 B.n729 B.n136 10.6151
R2866 B.n729 B.n728 10.6151
R2867 B.n728 B.n727 10.6151
R2868 B.n727 B.n138 10.6151
R2869 B.n723 B.n138 10.6151
R2870 B.n723 B.n722 10.6151
R2871 B.n722 B.n721 10.6151
R2872 B.n721 B.n140 10.6151
R2873 B.n717 B.n140 10.6151
R2874 B.n717 B.n716 10.6151
R2875 B.n716 B.n715 10.6151
R2876 B.n715 B.n142 10.6151
R2877 B.n711 B.n142 10.6151
R2878 B.n711 B.n710 10.6151
R2879 B.n710 B.n709 10.6151
R2880 B.n709 B.n144 10.6151
R2881 B.n705 B.n144 10.6151
R2882 B.n705 B.n704 10.6151
R2883 B.n704 B.n703 10.6151
R2884 B.n703 B.n146 10.6151
R2885 B.n699 B.n146 10.6151
R2886 B.n699 B.n698 10.6151
R2887 B.n698 B.n697 10.6151
R2888 B.n697 B.n148 10.6151
R2889 B.n693 B.n148 10.6151
R2890 B.n693 B.n692 10.6151
R2891 B.n692 B.n691 10.6151
R2892 B.n691 B.n150 10.6151
R2893 B.n687 B.n150 10.6151
R2894 B.n687 B.n686 10.6151
R2895 B.n686 B.n685 10.6151
R2896 B.n685 B.n152 10.6151
R2897 B.n681 B.n152 10.6151
R2898 B.n681 B.n680 10.6151
R2899 B.n680 B.n679 10.6151
R2900 B.n679 B.n154 10.6151
R2901 B.n675 B.n154 10.6151
R2902 B.n675 B.n674 10.6151
R2903 B.n674 B.n673 10.6151
R2904 B.n673 B.n156 10.6151
R2905 B.n669 B.n156 10.6151
R2906 B.n669 B.n668 10.6151
R2907 B.n668 B.n667 10.6151
R2908 B.n667 B.n158 10.6151
R2909 B.n663 B.n158 10.6151
R2910 B.n663 B.n662 10.6151
R2911 B.n662 B.n661 10.6151
R2912 B.n661 B.n160 10.6151
R2913 B.n657 B.n160 10.6151
R2914 B.n657 B.n656 10.6151
R2915 B.n656 B.n655 10.6151
R2916 B.n655 B.n162 10.6151
R2917 B.n651 B.n162 10.6151
R2918 B.n651 B.n650 10.6151
R2919 B.n650 B.n649 10.6151
R2920 B.n649 B.n164 10.6151
R2921 B.n645 B.n164 10.6151
R2922 B.n645 B.n644 10.6151
R2923 B.n644 B.n643 10.6151
R2924 B.n643 B.n166 10.6151
R2925 B.n639 B.n166 10.6151
R2926 B.n639 B.n638 10.6151
R2927 B.n638 B.n637 10.6151
R2928 B.n637 B.n168 10.6151
R2929 B.n633 B.n168 10.6151
R2930 B.n633 B.n632 10.6151
R2931 B.n632 B.n631 10.6151
R2932 B.n631 B.n170 10.6151
R2933 B.n627 B.n170 10.6151
R2934 B.n627 B.n626 10.6151
R2935 B.n626 B.n625 10.6151
R2936 B.n625 B.n172 10.6151
R2937 B.n621 B.n172 10.6151
R2938 B.n621 B.n620 10.6151
R2939 B.n620 B.n619 10.6151
R2940 B.n619 B.n174 10.6151
R2941 B.n615 B.n174 10.6151
R2942 B.n615 B.n614 10.6151
R2943 B.n614 B.n613 10.6151
R2944 B.n613 B.n176 10.6151
R2945 B.n609 B.n176 10.6151
R2946 B.n609 B.n608 10.6151
R2947 B.n608 B.n607 10.6151
R2948 B.n607 B.n178 10.6151
R2949 B.n603 B.n178 10.6151
R2950 B.n603 B.n602 10.6151
R2951 B.n602 B.n601 10.6151
R2952 B.n601 B.n180 10.6151
R2953 B.n597 B.n180 10.6151
R2954 B.n597 B.n596 10.6151
R2955 B.n596 B.n595 10.6151
R2956 B.n595 B.n182 10.6151
R2957 B.n591 B.n182 10.6151
R2958 B.n591 B.n590 10.6151
R2959 B.n590 B.n589 10.6151
R2960 B.n589 B.n184 10.6151
R2961 B.n585 B.n184 10.6151
R2962 B.n585 B.n584 10.6151
R2963 B.n584 B.n583 10.6151
R2964 B.n583 B.n186 10.6151
R2965 B.n286 B.n1 10.6151
R2966 B.n287 B.n286 10.6151
R2967 B.n287 B.n284 10.6151
R2968 B.n291 B.n284 10.6151
R2969 B.n292 B.n291 10.6151
R2970 B.n293 B.n292 10.6151
R2971 B.n293 B.n282 10.6151
R2972 B.n297 B.n282 10.6151
R2973 B.n298 B.n297 10.6151
R2974 B.n299 B.n298 10.6151
R2975 B.n299 B.n280 10.6151
R2976 B.n303 B.n280 10.6151
R2977 B.n304 B.n303 10.6151
R2978 B.n305 B.n304 10.6151
R2979 B.n305 B.n278 10.6151
R2980 B.n309 B.n278 10.6151
R2981 B.n310 B.n309 10.6151
R2982 B.n311 B.n310 10.6151
R2983 B.n311 B.n276 10.6151
R2984 B.n315 B.n276 10.6151
R2985 B.n316 B.n315 10.6151
R2986 B.n317 B.n316 10.6151
R2987 B.n317 B.n274 10.6151
R2988 B.n321 B.n274 10.6151
R2989 B.n322 B.n321 10.6151
R2990 B.n323 B.n322 10.6151
R2991 B.n323 B.n272 10.6151
R2992 B.n327 B.n272 10.6151
R2993 B.n328 B.n327 10.6151
R2994 B.n329 B.n328 10.6151
R2995 B.n329 B.n270 10.6151
R2996 B.n333 B.n270 10.6151
R2997 B.n334 B.n333 10.6151
R2998 B.n335 B.n334 10.6151
R2999 B.n335 B.n268 10.6151
R3000 B.n339 B.n268 10.6151
R3001 B.n340 B.n339 10.6151
R3002 B.n341 B.n340 10.6151
R3003 B.n341 B.n266 10.6151
R3004 B.n345 B.n266 10.6151
R3005 B.n346 B.n345 10.6151
R3006 B.n347 B.n346 10.6151
R3007 B.n347 B.n264 10.6151
R3008 B.n351 B.n264 10.6151
R3009 B.n352 B.n351 10.6151
R3010 B.n353 B.n352 10.6151
R3011 B.n353 B.n262 10.6151
R3012 B.n357 B.n262 10.6151
R3013 B.n358 B.n357 10.6151
R3014 B.n359 B.n358 10.6151
R3015 B.n359 B.n260 10.6151
R3016 B.n363 B.n260 10.6151
R3017 B.n364 B.n363 10.6151
R3018 B.n365 B.n364 10.6151
R3019 B.n365 B.n258 10.6151
R3020 B.n369 B.n258 10.6151
R3021 B.n370 B.n369 10.6151
R3022 B.n371 B.n370 10.6151
R3023 B.n371 B.n256 10.6151
R3024 B.n375 B.n256 10.6151
R3025 B.n376 B.n375 10.6151
R3026 B.n377 B.n376 10.6151
R3027 B.n377 B.n254 10.6151
R3028 B.n381 B.n254 10.6151
R3029 B.n382 B.n381 10.6151
R3030 B.n383 B.n382 10.6151
R3031 B.n383 B.n252 10.6151
R3032 B.n387 B.n252 10.6151
R3033 B.n388 B.n387 10.6151
R3034 B.n389 B.n388 10.6151
R3035 B.n389 B.n250 10.6151
R3036 B.n393 B.n250 10.6151
R3037 B.n394 B.n393 10.6151
R3038 B.n395 B.n394 10.6151
R3039 B.n395 B.n248 10.6151
R3040 B.n399 B.n248 10.6151
R3041 B.n400 B.n399 10.6151
R3042 B.n401 B.n400 10.6151
R3043 B.n401 B.n246 10.6151
R3044 B.n405 B.n246 10.6151
R3045 B.n406 B.n405 10.6151
R3046 B.n407 B.n244 10.6151
R3047 B.n411 B.n244 10.6151
R3048 B.n412 B.n411 10.6151
R3049 B.n413 B.n412 10.6151
R3050 B.n413 B.n242 10.6151
R3051 B.n417 B.n242 10.6151
R3052 B.n418 B.n417 10.6151
R3053 B.n419 B.n418 10.6151
R3054 B.n419 B.n240 10.6151
R3055 B.n423 B.n240 10.6151
R3056 B.n424 B.n423 10.6151
R3057 B.n425 B.n424 10.6151
R3058 B.n425 B.n238 10.6151
R3059 B.n429 B.n238 10.6151
R3060 B.n430 B.n429 10.6151
R3061 B.n431 B.n430 10.6151
R3062 B.n431 B.n236 10.6151
R3063 B.n435 B.n236 10.6151
R3064 B.n436 B.n435 10.6151
R3065 B.n437 B.n436 10.6151
R3066 B.n437 B.n234 10.6151
R3067 B.n441 B.n234 10.6151
R3068 B.n442 B.n441 10.6151
R3069 B.n443 B.n442 10.6151
R3070 B.n443 B.n232 10.6151
R3071 B.n447 B.n232 10.6151
R3072 B.n448 B.n447 10.6151
R3073 B.n449 B.n448 10.6151
R3074 B.n449 B.n230 10.6151
R3075 B.n453 B.n230 10.6151
R3076 B.n454 B.n453 10.6151
R3077 B.n455 B.n454 10.6151
R3078 B.n455 B.n228 10.6151
R3079 B.n459 B.n228 10.6151
R3080 B.n460 B.n459 10.6151
R3081 B.n461 B.n460 10.6151
R3082 B.n461 B.n226 10.6151
R3083 B.n465 B.n226 10.6151
R3084 B.n466 B.n465 10.6151
R3085 B.n467 B.n466 10.6151
R3086 B.n467 B.n224 10.6151
R3087 B.n471 B.n224 10.6151
R3088 B.n472 B.n471 10.6151
R3089 B.n473 B.n472 10.6151
R3090 B.n473 B.n222 10.6151
R3091 B.n477 B.n222 10.6151
R3092 B.n478 B.n477 10.6151
R3093 B.n479 B.n478 10.6151
R3094 B.n479 B.n220 10.6151
R3095 B.n483 B.n220 10.6151
R3096 B.n484 B.n483 10.6151
R3097 B.n486 B.n216 10.6151
R3098 B.n490 B.n216 10.6151
R3099 B.n491 B.n490 10.6151
R3100 B.n492 B.n491 10.6151
R3101 B.n492 B.n214 10.6151
R3102 B.n496 B.n214 10.6151
R3103 B.n497 B.n496 10.6151
R3104 B.n501 B.n497 10.6151
R3105 B.n505 B.n212 10.6151
R3106 B.n506 B.n505 10.6151
R3107 B.n507 B.n506 10.6151
R3108 B.n507 B.n210 10.6151
R3109 B.n511 B.n210 10.6151
R3110 B.n512 B.n511 10.6151
R3111 B.n513 B.n512 10.6151
R3112 B.n513 B.n208 10.6151
R3113 B.n517 B.n208 10.6151
R3114 B.n518 B.n517 10.6151
R3115 B.n519 B.n518 10.6151
R3116 B.n519 B.n206 10.6151
R3117 B.n523 B.n206 10.6151
R3118 B.n524 B.n523 10.6151
R3119 B.n525 B.n524 10.6151
R3120 B.n525 B.n204 10.6151
R3121 B.n529 B.n204 10.6151
R3122 B.n530 B.n529 10.6151
R3123 B.n531 B.n530 10.6151
R3124 B.n531 B.n202 10.6151
R3125 B.n535 B.n202 10.6151
R3126 B.n536 B.n535 10.6151
R3127 B.n537 B.n536 10.6151
R3128 B.n537 B.n200 10.6151
R3129 B.n541 B.n200 10.6151
R3130 B.n542 B.n541 10.6151
R3131 B.n543 B.n542 10.6151
R3132 B.n543 B.n198 10.6151
R3133 B.n547 B.n198 10.6151
R3134 B.n548 B.n547 10.6151
R3135 B.n549 B.n548 10.6151
R3136 B.n549 B.n196 10.6151
R3137 B.n553 B.n196 10.6151
R3138 B.n554 B.n553 10.6151
R3139 B.n555 B.n554 10.6151
R3140 B.n555 B.n194 10.6151
R3141 B.n559 B.n194 10.6151
R3142 B.n560 B.n559 10.6151
R3143 B.n561 B.n560 10.6151
R3144 B.n561 B.n192 10.6151
R3145 B.n565 B.n192 10.6151
R3146 B.n566 B.n565 10.6151
R3147 B.n567 B.n566 10.6151
R3148 B.n567 B.n190 10.6151
R3149 B.n571 B.n190 10.6151
R3150 B.n572 B.n571 10.6151
R3151 B.n573 B.n572 10.6151
R3152 B.n573 B.n188 10.6151
R3153 B.n577 B.n188 10.6151
R3154 B.n578 B.n577 10.6151
R3155 B.n579 B.n578 10.6151
R3156 B.n1125 B.n0 8.11757
R3157 B.n1125 B.n1 8.11757
R3158 B.n922 B.n921 6.5566
R3159 B.n909 B.n908 6.5566
R3160 B.n486 B.n485 6.5566
R3161 B.n501 B.n500 6.5566
R3162 B.n923 B.n922 4.05904
R3163 B.n908 B.n907 4.05904
R3164 B.n485 B.n484 4.05904
R3165 B.n500 B.n212 4.05904
C0 VDD1 VDD2 3.00913f
C1 B VP 2.98679f
C2 B VN 1.65469f
C3 VTAIL B 5.04322f
C4 w_n6022_n4064# B 13.6743f
C5 VDD1 B 3.25824f
C6 B VDD2 3.426f
C7 VP VN 10.9252f
C8 VTAIL VP 15.5913f
C9 w_n6022_n4064# VP 14.1122f
C10 VTAIL VN 15.5762f
C11 VDD1 VP 15.139401f
C12 w_n6022_n4064# VN 13.3242f
C13 VTAIL w_n6022_n4064# 3.86239f
C14 VDD1 VN 0.156686f
C15 VTAIL VDD1 12.407201f
C16 VP VDD2 0.746667f
C17 VDD1 w_n6022_n4064# 3.50847f
C18 VN VDD2 14.553f
C19 VTAIL VDD2 12.4672f
C20 w_n6022_n4064# VDD2 3.71855f
C21 VDD2 VSUBS 2.70118f
C22 VDD1 VSUBS 2.591437f
C23 VTAIL VSUBS 1.724658f
C24 VN VSUBS 9.94759f
C25 VP VSUBS 6.010328f
C26 B VSUBS 7.246088f
C27 w_n6022_n4064# VSUBS 0.299968p
C28 B.n0 VSUBS 0.007026f
C29 B.n1 VSUBS 0.007026f
C30 B.n2 VSUBS 0.010392f
C31 B.n3 VSUBS 0.007963f
C32 B.n4 VSUBS 0.007963f
C33 B.n5 VSUBS 0.007963f
C34 B.n6 VSUBS 0.007963f
C35 B.n7 VSUBS 0.007963f
C36 B.n8 VSUBS 0.007963f
C37 B.n9 VSUBS 0.007963f
C38 B.n10 VSUBS 0.007963f
C39 B.n11 VSUBS 0.007963f
C40 B.n12 VSUBS 0.007963f
C41 B.n13 VSUBS 0.007963f
C42 B.n14 VSUBS 0.007963f
C43 B.n15 VSUBS 0.007963f
C44 B.n16 VSUBS 0.007963f
C45 B.n17 VSUBS 0.007963f
C46 B.n18 VSUBS 0.007963f
C47 B.n19 VSUBS 0.007963f
C48 B.n20 VSUBS 0.007963f
C49 B.n21 VSUBS 0.007963f
C50 B.n22 VSUBS 0.007963f
C51 B.n23 VSUBS 0.007963f
C52 B.n24 VSUBS 0.007963f
C53 B.n25 VSUBS 0.007963f
C54 B.n26 VSUBS 0.007963f
C55 B.n27 VSUBS 0.007963f
C56 B.n28 VSUBS 0.007963f
C57 B.n29 VSUBS 0.007963f
C58 B.n30 VSUBS 0.007963f
C59 B.n31 VSUBS 0.007963f
C60 B.n32 VSUBS 0.007963f
C61 B.n33 VSUBS 0.007963f
C62 B.n34 VSUBS 0.007963f
C63 B.n35 VSUBS 0.007963f
C64 B.n36 VSUBS 0.007963f
C65 B.n37 VSUBS 0.007963f
C66 B.n38 VSUBS 0.007963f
C67 B.n39 VSUBS 0.007963f
C68 B.n40 VSUBS 0.007963f
C69 B.n41 VSUBS 0.007963f
C70 B.n42 VSUBS 0.007963f
C71 B.n43 VSUBS 0.018999f
C72 B.n44 VSUBS 0.007963f
C73 B.n45 VSUBS 0.007963f
C74 B.n46 VSUBS 0.007963f
C75 B.n47 VSUBS 0.007963f
C76 B.n48 VSUBS 0.007963f
C77 B.n49 VSUBS 0.007963f
C78 B.n50 VSUBS 0.007963f
C79 B.n51 VSUBS 0.007963f
C80 B.n52 VSUBS 0.007963f
C81 B.n53 VSUBS 0.007963f
C82 B.n54 VSUBS 0.007963f
C83 B.n55 VSUBS 0.007963f
C84 B.n56 VSUBS 0.007963f
C85 B.n57 VSUBS 0.007963f
C86 B.n58 VSUBS 0.007963f
C87 B.n59 VSUBS 0.007963f
C88 B.n60 VSUBS 0.007963f
C89 B.n61 VSUBS 0.007963f
C90 B.n62 VSUBS 0.007963f
C91 B.n63 VSUBS 0.007963f
C92 B.n64 VSUBS 0.007963f
C93 B.n65 VSUBS 0.007963f
C94 B.n66 VSUBS 0.007963f
C95 B.n67 VSUBS 0.007963f
C96 B.n68 VSUBS 0.007963f
C97 B.n69 VSUBS 0.007963f
C98 B.t4 VSUBS 0.330935f
C99 B.t5 VSUBS 0.383292f
C100 B.t3 VSUBS 3.1461f
C101 B.n70 VSUBS 0.611987f
C102 B.n71 VSUBS 0.344788f
C103 B.n72 VSUBS 0.007963f
C104 B.n73 VSUBS 0.007963f
C105 B.n74 VSUBS 0.007963f
C106 B.n75 VSUBS 0.007963f
C107 B.t1 VSUBS 0.330939f
C108 B.t2 VSUBS 0.383296f
C109 B.t0 VSUBS 3.1461f
C110 B.n76 VSUBS 0.611984f
C111 B.n77 VSUBS 0.344784f
C112 B.n78 VSUBS 0.007963f
C113 B.n79 VSUBS 0.007963f
C114 B.n80 VSUBS 0.007963f
C115 B.n81 VSUBS 0.007963f
C116 B.n82 VSUBS 0.007963f
C117 B.n83 VSUBS 0.007963f
C118 B.n84 VSUBS 0.007963f
C119 B.n85 VSUBS 0.007963f
C120 B.n86 VSUBS 0.007963f
C121 B.n87 VSUBS 0.007963f
C122 B.n88 VSUBS 0.007963f
C123 B.n89 VSUBS 0.007963f
C124 B.n90 VSUBS 0.007963f
C125 B.n91 VSUBS 0.007963f
C126 B.n92 VSUBS 0.007963f
C127 B.n93 VSUBS 0.007963f
C128 B.n94 VSUBS 0.007963f
C129 B.n95 VSUBS 0.007963f
C130 B.n96 VSUBS 0.007963f
C131 B.n97 VSUBS 0.007963f
C132 B.n98 VSUBS 0.007963f
C133 B.n99 VSUBS 0.007963f
C134 B.n100 VSUBS 0.007963f
C135 B.n101 VSUBS 0.007963f
C136 B.n102 VSUBS 0.007963f
C137 B.n103 VSUBS 0.018999f
C138 B.n104 VSUBS 0.007963f
C139 B.n105 VSUBS 0.007963f
C140 B.n106 VSUBS 0.007963f
C141 B.n107 VSUBS 0.007963f
C142 B.n108 VSUBS 0.007963f
C143 B.n109 VSUBS 0.007963f
C144 B.n110 VSUBS 0.007963f
C145 B.n111 VSUBS 0.007963f
C146 B.n112 VSUBS 0.007963f
C147 B.n113 VSUBS 0.007963f
C148 B.n114 VSUBS 0.007963f
C149 B.n115 VSUBS 0.007963f
C150 B.n116 VSUBS 0.007963f
C151 B.n117 VSUBS 0.007963f
C152 B.n118 VSUBS 0.007963f
C153 B.n119 VSUBS 0.007963f
C154 B.n120 VSUBS 0.007963f
C155 B.n121 VSUBS 0.007963f
C156 B.n122 VSUBS 0.007963f
C157 B.n123 VSUBS 0.007963f
C158 B.n124 VSUBS 0.007963f
C159 B.n125 VSUBS 0.007963f
C160 B.n126 VSUBS 0.007963f
C161 B.n127 VSUBS 0.007963f
C162 B.n128 VSUBS 0.007963f
C163 B.n129 VSUBS 0.007963f
C164 B.n130 VSUBS 0.007963f
C165 B.n131 VSUBS 0.007963f
C166 B.n132 VSUBS 0.007963f
C167 B.n133 VSUBS 0.007963f
C168 B.n134 VSUBS 0.007963f
C169 B.n135 VSUBS 0.007963f
C170 B.n136 VSUBS 0.007963f
C171 B.n137 VSUBS 0.007963f
C172 B.n138 VSUBS 0.007963f
C173 B.n139 VSUBS 0.007963f
C174 B.n140 VSUBS 0.007963f
C175 B.n141 VSUBS 0.007963f
C176 B.n142 VSUBS 0.007963f
C177 B.n143 VSUBS 0.007963f
C178 B.n144 VSUBS 0.007963f
C179 B.n145 VSUBS 0.007963f
C180 B.n146 VSUBS 0.007963f
C181 B.n147 VSUBS 0.007963f
C182 B.n148 VSUBS 0.007963f
C183 B.n149 VSUBS 0.007963f
C184 B.n150 VSUBS 0.007963f
C185 B.n151 VSUBS 0.007963f
C186 B.n152 VSUBS 0.007963f
C187 B.n153 VSUBS 0.007963f
C188 B.n154 VSUBS 0.007963f
C189 B.n155 VSUBS 0.007963f
C190 B.n156 VSUBS 0.007963f
C191 B.n157 VSUBS 0.007963f
C192 B.n158 VSUBS 0.007963f
C193 B.n159 VSUBS 0.007963f
C194 B.n160 VSUBS 0.007963f
C195 B.n161 VSUBS 0.007963f
C196 B.n162 VSUBS 0.007963f
C197 B.n163 VSUBS 0.007963f
C198 B.n164 VSUBS 0.007963f
C199 B.n165 VSUBS 0.007963f
C200 B.n166 VSUBS 0.007963f
C201 B.n167 VSUBS 0.007963f
C202 B.n168 VSUBS 0.007963f
C203 B.n169 VSUBS 0.007963f
C204 B.n170 VSUBS 0.007963f
C205 B.n171 VSUBS 0.007963f
C206 B.n172 VSUBS 0.007963f
C207 B.n173 VSUBS 0.007963f
C208 B.n174 VSUBS 0.007963f
C209 B.n175 VSUBS 0.007963f
C210 B.n176 VSUBS 0.007963f
C211 B.n177 VSUBS 0.007963f
C212 B.n178 VSUBS 0.007963f
C213 B.n179 VSUBS 0.007963f
C214 B.n180 VSUBS 0.007963f
C215 B.n181 VSUBS 0.007963f
C216 B.n182 VSUBS 0.007963f
C217 B.n183 VSUBS 0.007963f
C218 B.n184 VSUBS 0.007963f
C219 B.n185 VSUBS 0.007963f
C220 B.n186 VSUBS 0.019409f
C221 B.n187 VSUBS 0.007963f
C222 B.n188 VSUBS 0.007963f
C223 B.n189 VSUBS 0.007963f
C224 B.n190 VSUBS 0.007963f
C225 B.n191 VSUBS 0.007963f
C226 B.n192 VSUBS 0.007963f
C227 B.n193 VSUBS 0.007963f
C228 B.n194 VSUBS 0.007963f
C229 B.n195 VSUBS 0.007963f
C230 B.n196 VSUBS 0.007963f
C231 B.n197 VSUBS 0.007963f
C232 B.n198 VSUBS 0.007963f
C233 B.n199 VSUBS 0.007963f
C234 B.n200 VSUBS 0.007963f
C235 B.n201 VSUBS 0.007963f
C236 B.n202 VSUBS 0.007963f
C237 B.n203 VSUBS 0.007963f
C238 B.n204 VSUBS 0.007963f
C239 B.n205 VSUBS 0.007963f
C240 B.n206 VSUBS 0.007963f
C241 B.n207 VSUBS 0.007963f
C242 B.n208 VSUBS 0.007963f
C243 B.n209 VSUBS 0.007963f
C244 B.n210 VSUBS 0.007963f
C245 B.n211 VSUBS 0.007963f
C246 B.n212 VSUBS 0.005504f
C247 B.n213 VSUBS 0.007963f
C248 B.n214 VSUBS 0.007963f
C249 B.n215 VSUBS 0.007963f
C250 B.n216 VSUBS 0.007963f
C251 B.n217 VSUBS 0.007963f
C252 B.t8 VSUBS 0.330935f
C253 B.t7 VSUBS 0.383292f
C254 B.t6 VSUBS 3.1461f
C255 B.n218 VSUBS 0.611987f
C256 B.n219 VSUBS 0.344788f
C257 B.n220 VSUBS 0.007963f
C258 B.n221 VSUBS 0.007963f
C259 B.n222 VSUBS 0.007963f
C260 B.n223 VSUBS 0.007963f
C261 B.n224 VSUBS 0.007963f
C262 B.n225 VSUBS 0.007963f
C263 B.n226 VSUBS 0.007963f
C264 B.n227 VSUBS 0.007963f
C265 B.n228 VSUBS 0.007963f
C266 B.n229 VSUBS 0.007963f
C267 B.n230 VSUBS 0.007963f
C268 B.n231 VSUBS 0.007963f
C269 B.n232 VSUBS 0.007963f
C270 B.n233 VSUBS 0.007963f
C271 B.n234 VSUBS 0.007963f
C272 B.n235 VSUBS 0.007963f
C273 B.n236 VSUBS 0.007963f
C274 B.n237 VSUBS 0.007963f
C275 B.n238 VSUBS 0.007963f
C276 B.n239 VSUBS 0.007963f
C277 B.n240 VSUBS 0.007963f
C278 B.n241 VSUBS 0.007963f
C279 B.n242 VSUBS 0.007963f
C280 B.n243 VSUBS 0.007963f
C281 B.n244 VSUBS 0.007963f
C282 B.n245 VSUBS 0.018476f
C283 B.n246 VSUBS 0.007963f
C284 B.n247 VSUBS 0.007963f
C285 B.n248 VSUBS 0.007963f
C286 B.n249 VSUBS 0.007963f
C287 B.n250 VSUBS 0.007963f
C288 B.n251 VSUBS 0.007963f
C289 B.n252 VSUBS 0.007963f
C290 B.n253 VSUBS 0.007963f
C291 B.n254 VSUBS 0.007963f
C292 B.n255 VSUBS 0.007963f
C293 B.n256 VSUBS 0.007963f
C294 B.n257 VSUBS 0.007963f
C295 B.n258 VSUBS 0.007963f
C296 B.n259 VSUBS 0.007963f
C297 B.n260 VSUBS 0.007963f
C298 B.n261 VSUBS 0.007963f
C299 B.n262 VSUBS 0.007963f
C300 B.n263 VSUBS 0.007963f
C301 B.n264 VSUBS 0.007963f
C302 B.n265 VSUBS 0.007963f
C303 B.n266 VSUBS 0.007963f
C304 B.n267 VSUBS 0.007963f
C305 B.n268 VSUBS 0.007963f
C306 B.n269 VSUBS 0.007963f
C307 B.n270 VSUBS 0.007963f
C308 B.n271 VSUBS 0.007963f
C309 B.n272 VSUBS 0.007963f
C310 B.n273 VSUBS 0.007963f
C311 B.n274 VSUBS 0.007963f
C312 B.n275 VSUBS 0.007963f
C313 B.n276 VSUBS 0.007963f
C314 B.n277 VSUBS 0.007963f
C315 B.n278 VSUBS 0.007963f
C316 B.n279 VSUBS 0.007963f
C317 B.n280 VSUBS 0.007963f
C318 B.n281 VSUBS 0.007963f
C319 B.n282 VSUBS 0.007963f
C320 B.n283 VSUBS 0.007963f
C321 B.n284 VSUBS 0.007963f
C322 B.n285 VSUBS 0.007963f
C323 B.n286 VSUBS 0.007963f
C324 B.n287 VSUBS 0.007963f
C325 B.n288 VSUBS 0.007963f
C326 B.n289 VSUBS 0.007963f
C327 B.n290 VSUBS 0.007963f
C328 B.n291 VSUBS 0.007963f
C329 B.n292 VSUBS 0.007963f
C330 B.n293 VSUBS 0.007963f
C331 B.n294 VSUBS 0.007963f
C332 B.n295 VSUBS 0.007963f
C333 B.n296 VSUBS 0.007963f
C334 B.n297 VSUBS 0.007963f
C335 B.n298 VSUBS 0.007963f
C336 B.n299 VSUBS 0.007963f
C337 B.n300 VSUBS 0.007963f
C338 B.n301 VSUBS 0.007963f
C339 B.n302 VSUBS 0.007963f
C340 B.n303 VSUBS 0.007963f
C341 B.n304 VSUBS 0.007963f
C342 B.n305 VSUBS 0.007963f
C343 B.n306 VSUBS 0.007963f
C344 B.n307 VSUBS 0.007963f
C345 B.n308 VSUBS 0.007963f
C346 B.n309 VSUBS 0.007963f
C347 B.n310 VSUBS 0.007963f
C348 B.n311 VSUBS 0.007963f
C349 B.n312 VSUBS 0.007963f
C350 B.n313 VSUBS 0.007963f
C351 B.n314 VSUBS 0.007963f
C352 B.n315 VSUBS 0.007963f
C353 B.n316 VSUBS 0.007963f
C354 B.n317 VSUBS 0.007963f
C355 B.n318 VSUBS 0.007963f
C356 B.n319 VSUBS 0.007963f
C357 B.n320 VSUBS 0.007963f
C358 B.n321 VSUBS 0.007963f
C359 B.n322 VSUBS 0.007963f
C360 B.n323 VSUBS 0.007963f
C361 B.n324 VSUBS 0.007963f
C362 B.n325 VSUBS 0.007963f
C363 B.n326 VSUBS 0.007963f
C364 B.n327 VSUBS 0.007963f
C365 B.n328 VSUBS 0.007963f
C366 B.n329 VSUBS 0.007963f
C367 B.n330 VSUBS 0.007963f
C368 B.n331 VSUBS 0.007963f
C369 B.n332 VSUBS 0.007963f
C370 B.n333 VSUBS 0.007963f
C371 B.n334 VSUBS 0.007963f
C372 B.n335 VSUBS 0.007963f
C373 B.n336 VSUBS 0.007963f
C374 B.n337 VSUBS 0.007963f
C375 B.n338 VSUBS 0.007963f
C376 B.n339 VSUBS 0.007963f
C377 B.n340 VSUBS 0.007963f
C378 B.n341 VSUBS 0.007963f
C379 B.n342 VSUBS 0.007963f
C380 B.n343 VSUBS 0.007963f
C381 B.n344 VSUBS 0.007963f
C382 B.n345 VSUBS 0.007963f
C383 B.n346 VSUBS 0.007963f
C384 B.n347 VSUBS 0.007963f
C385 B.n348 VSUBS 0.007963f
C386 B.n349 VSUBS 0.007963f
C387 B.n350 VSUBS 0.007963f
C388 B.n351 VSUBS 0.007963f
C389 B.n352 VSUBS 0.007963f
C390 B.n353 VSUBS 0.007963f
C391 B.n354 VSUBS 0.007963f
C392 B.n355 VSUBS 0.007963f
C393 B.n356 VSUBS 0.007963f
C394 B.n357 VSUBS 0.007963f
C395 B.n358 VSUBS 0.007963f
C396 B.n359 VSUBS 0.007963f
C397 B.n360 VSUBS 0.007963f
C398 B.n361 VSUBS 0.007963f
C399 B.n362 VSUBS 0.007963f
C400 B.n363 VSUBS 0.007963f
C401 B.n364 VSUBS 0.007963f
C402 B.n365 VSUBS 0.007963f
C403 B.n366 VSUBS 0.007963f
C404 B.n367 VSUBS 0.007963f
C405 B.n368 VSUBS 0.007963f
C406 B.n369 VSUBS 0.007963f
C407 B.n370 VSUBS 0.007963f
C408 B.n371 VSUBS 0.007963f
C409 B.n372 VSUBS 0.007963f
C410 B.n373 VSUBS 0.007963f
C411 B.n374 VSUBS 0.007963f
C412 B.n375 VSUBS 0.007963f
C413 B.n376 VSUBS 0.007963f
C414 B.n377 VSUBS 0.007963f
C415 B.n378 VSUBS 0.007963f
C416 B.n379 VSUBS 0.007963f
C417 B.n380 VSUBS 0.007963f
C418 B.n381 VSUBS 0.007963f
C419 B.n382 VSUBS 0.007963f
C420 B.n383 VSUBS 0.007963f
C421 B.n384 VSUBS 0.007963f
C422 B.n385 VSUBS 0.007963f
C423 B.n386 VSUBS 0.007963f
C424 B.n387 VSUBS 0.007963f
C425 B.n388 VSUBS 0.007963f
C426 B.n389 VSUBS 0.007963f
C427 B.n390 VSUBS 0.007963f
C428 B.n391 VSUBS 0.007963f
C429 B.n392 VSUBS 0.007963f
C430 B.n393 VSUBS 0.007963f
C431 B.n394 VSUBS 0.007963f
C432 B.n395 VSUBS 0.007963f
C433 B.n396 VSUBS 0.007963f
C434 B.n397 VSUBS 0.007963f
C435 B.n398 VSUBS 0.007963f
C436 B.n399 VSUBS 0.007963f
C437 B.n400 VSUBS 0.007963f
C438 B.n401 VSUBS 0.007963f
C439 B.n402 VSUBS 0.007963f
C440 B.n403 VSUBS 0.007963f
C441 B.n404 VSUBS 0.007963f
C442 B.n405 VSUBS 0.007963f
C443 B.n406 VSUBS 0.018476f
C444 B.n407 VSUBS 0.018999f
C445 B.n408 VSUBS 0.018999f
C446 B.n409 VSUBS 0.007963f
C447 B.n410 VSUBS 0.007963f
C448 B.n411 VSUBS 0.007963f
C449 B.n412 VSUBS 0.007963f
C450 B.n413 VSUBS 0.007963f
C451 B.n414 VSUBS 0.007963f
C452 B.n415 VSUBS 0.007963f
C453 B.n416 VSUBS 0.007963f
C454 B.n417 VSUBS 0.007963f
C455 B.n418 VSUBS 0.007963f
C456 B.n419 VSUBS 0.007963f
C457 B.n420 VSUBS 0.007963f
C458 B.n421 VSUBS 0.007963f
C459 B.n422 VSUBS 0.007963f
C460 B.n423 VSUBS 0.007963f
C461 B.n424 VSUBS 0.007963f
C462 B.n425 VSUBS 0.007963f
C463 B.n426 VSUBS 0.007963f
C464 B.n427 VSUBS 0.007963f
C465 B.n428 VSUBS 0.007963f
C466 B.n429 VSUBS 0.007963f
C467 B.n430 VSUBS 0.007963f
C468 B.n431 VSUBS 0.007963f
C469 B.n432 VSUBS 0.007963f
C470 B.n433 VSUBS 0.007963f
C471 B.n434 VSUBS 0.007963f
C472 B.n435 VSUBS 0.007963f
C473 B.n436 VSUBS 0.007963f
C474 B.n437 VSUBS 0.007963f
C475 B.n438 VSUBS 0.007963f
C476 B.n439 VSUBS 0.007963f
C477 B.n440 VSUBS 0.007963f
C478 B.n441 VSUBS 0.007963f
C479 B.n442 VSUBS 0.007963f
C480 B.n443 VSUBS 0.007963f
C481 B.n444 VSUBS 0.007963f
C482 B.n445 VSUBS 0.007963f
C483 B.n446 VSUBS 0.007963f
C484 B.n447 VSUBS 0.007963f
C485 B.n448 VSUBS 0.007963f
C486 B.n449 VSUBS 0.007963f
C487 B.n450 VSUBS 0.007963f
C488 B.n451 VSUBS 0.007963f
C489 B.n452 VSUBS 0.007963f
C490 B.n453 VSUBS 0.007963f
C491 B.n454 VSUBS 0.007963f
C492 B.n455 VSUBS 0.007963f
C493 B.n456 VSUBS 0.007963f
C494 B.n457 VSUBS 0.007963f
C495 B.n458 VSUBS 0.007963f
C496 B.n459 VSUBS 0.007963f
C497 B.n460 VSUBS 0.007963f
C498 B.n461 VSUBS 0.007963f
C499 B.n462 VSUBS 0.007963f
C500 B.n463 VSUBS 0.007963f
C501 B.n464 VSUBS 0.007963f
C502 B.n465 VSUBS 0.007963f
C503 B.n466 VSUBS 0.007963f
C504 B.n467 VSUBS 0.007963f
C505 B.n468 VSUBS 0.007963f
C506 B.n469 VSUBS 0.007963f
C507 B.n470 VSUBS 0.007963f
C508 B.n471 VSUBS 0.007963f
C509 B.n472 VSUBS 0.007963f
C510 B.n473 VSUBS 0.007963f
C511 B.n474 VSUBS 0.007963f
C512 B.n475 VSUBS 0.007963f
C513 B.n476 VSUBS 0.007963f
C514 B.n477 VSUBS 0.007963f
C515 B.n478 VSUBS 0.007963f
C516 B.n479 VSUBS 0.007963f
C517 B.n480 VSUBS 0.007963f
C518 B.n481 VSUBS 0.007963f
C519 B.n482 VSUBS 0.007963f
C520 B.n483 VSUBS 0.007963f
C521 B.n484 VSUBS 0.005504f
C522 B.n485 VSUBS 0.01845f
C523 B.n486 VSUBS 0.006441f
C524 B.n487 VSUBS 0.007963f
C525 B.n488 VSUBS 0.007963f
C526 B.n489 VSUBS 0.007963f
C527 B.n490 VSUBS 0.007963f
C528 B.n491 VSUBS 0.007963f
C529 B.n492 VSUBS 0.007963f
C530 B.n493 VSUBS 0.007963f
C531 B.n494 VSUBS 0.007963f
C532 B.n495 VSUBS 0.007963f
C533 B.n496 VSUBS 0.007963f
C534 B.n497 VSUBS 0.007963f
C535 B.t11 VSUBS 0.330939f
C536 B.t10 VSUBS 0.383296f
C537 B.t9 VSUBS 3.1461f
C538 B.n498 VSUBS 0.611984f
C539 B.n499 VSUBS 0.344784f
C540 B.n500 VSUBS 0.01845f
C541 B.n501 VSUBS 0.006441f
C542 B.n502 VSUBS 0.007963f
C543 B.n503 VSUBS 0.007963f
C544 B.n504 VSUBS 0.007963f
C545 B.n505 VSUBS 0.007963f
C546 B.n506 VSUBS 0.007963f
C547 B.n507 VSUBS 0.007963f
C548 B.n508 VSUBS 0.007963f
C549 B.n509 VSUBS 0.007963f
C550 B.n510 VSUBS 0.007963f
C551 B.n511 VSUBS 0.007963f
C552 B.n512 VSUBS 0.007963f
C553 B.n513 VSUBS 0.007963f
C554 B.n514 VSUBS 0.007963f
C555 B.n515 VSUBS 0.007963f
C556 B.n516 VSUBS 0.007963f
C557 B.n517 VSUBS 0.007963f
C558 B.n518 VSUBS 0.007963f
C559 B.n519 VSUBS 0.007963f
C560 B.n520 VSUBS 0.007963f
C561 B.n521 VSUBS 0.007963f
C562 B.n522 VSUBS 0.007963f
C563 B.n523 VSUBS 0.007963f
C564 B.n524 VSUBS 0.007963f
C565 B.n525 VSUBS 0.007963f
C566 B.n526 VSUBS 0.007963f
C567 B.n527 VSUBS 0.007963f
C568 B.n528 VSUBS 0.007963f
C569 B.n529 VSUBS 0.007963f
C570 B.n530 VSUBS 0.007963f
C571 B.n531 VSUBS 0.007963f
C572 B.n532 VSUBS 0.007963f
C573 B.n533 VSUBS 0.007963f
C574 B.n534 VSUBS 0.007963f
C575 B.n535 VSUBS 0.007963f
C576 B.n536 VSUBS 0.007963f
C577 B.n537 VSUBS 0.007963f
C578 B.n538 VSUBS 0.007963f
C579 B.n539 VSUBS 0.007963f
C580 B.n540 VSUBS 0.007963f
C581 B.n541 VSUBS 0.007963f
C582 B.n542 VSUBS 0.007963f
C583 B.n543 VSUBS 0.007963f
C584 B.n544 VSUBS 0.007963f
C585 B.n545 VSUBS 0.007963f
C586 B.n546 VSUBS 0.007963f
C587 B.n547 VSUBS 0.007963f
C588 B.n548 VSUBS 0.007963f
C589 B.n549 VSUBS 0.007963f
C590 B.n550 VSUBS 0.007963f
C591 B.n551 VSUBS 0.007963f
C592 B.n552 VSUBS 0.007963f
C593 B.n553 VSUBS 0.007963f
C594 B.n554 VSUBS 0.007963f
C595 B.n555 VSUBS 0.007963f
C596 B.n556 VSUBS 0.007963f
C597 B.n557 VSUBS 0.007963f
C598 B.n558 VSUBS 0.007963f
C599 B.n559 VSUBS 0.007963f
C600 B.n560 VSUBS 0.007963f
C601 B.n561 VSUBS 0.007963f
C602 B.n562 VSUBS 0.007963f
C603 B.n563 VSUBS 0.007963f
C604 B.n564 VSUBS 0.007963f
C605 B.n565 VSUBS 0.007963f
C606 B.n566 VSUBS 0.007963f
C607 B.n567 VSUBS 0.007963f
C608 B.n568 VSUBS 0.007963f
C609 B.n569 VSUBS 0.007963f
C610 B.n570 VSUBS 0.007963f
C611 B.n571 VSUBS 0.007963f
C612 B.n572 VSUBS 0.007963f
C613 B.n573 VSUBS 0.007963f
C614 B.n574 VSUBS 0.007963f
C615 B.n575 VSUBS 0.007963f
C616 B.n576 VSUBS 0.007963f
C617 B.n577 VSUBS 0.007963f
C618 B.n578 VSUBS 0.007963f
C619 B.n579 VSUBS 0.018066f
C620 B.n580 VSUBS 0.018999f
C621 B.n581 VSUBS 0.018476f
C622 B.n582 VSUBS 0.007963f
C623 B.n583 VSUBS 0.007963f
C624 B.n584 VSUBS 0.007963f
C625 B.n585 VSUBS 0.007963f
C626 B.n586 VSUBS 0.007963f
C627 B.n587 VSUBS 0.007963f
C628 B.n588 VSUBS 0.007963f
C629 B.n589 VSUBS 0.007963f
C630 B.n590 VSUBS 0.007963f
C631 B.n591 VSUBS 0.007963f
C632 B.n592 VSUBS 0.007963f
C633 B.n593 VSUBS 0.007963f
C634 B.n594 VSUBS 0.007963f
C635 B.n595 VSUBS 0.007963f
C636 B.n596 VSUBS 0.007963f
C637 B.n597 VSUBS 0.007963f
C638 B.n598 VSUBS 0.007963f
C639 B.n599 VSUBS 0.007963f
C640 B.n600 VSUBS 0.007963f
C641 B.n601 VSUBS 0.007963f
C642 B.n602 VSUBS 0.007963f
C643 B.n603 VSUBS 0.007963f
C644 B.n604 VSUBS 0.007963f
C645 B.n605 VSUBS 0.007963f
C646 B.n606 VSUBS 0.007963f
C647 B.n607 VSUBS 0.007963f
C648 B.n608 VSUBS 0.007963f
C649 B.n609 VSUBS 0.007963f
C650 B.n610 VSUBS 0.007963f
C651 B.n611 VSUBS 0.007963f
C652 B.n612 VSUBS 0.007963f
C653 B.n613 VSUBS 0.007963f
C654 B.n614 VSUBS 0.007963f
C655 B.n615 VSUBS 0.007963f
C656 B.n616 VSUBS 0.007963f
C657 B.n617 VSUBS 0.007963f
C658 B.n618 VSUBS 0.007963f
C659 B.n619 VSUBS 0.007963f
C660 B.n620 VSUBS 0.007963f
C661 B.n621 VSUBS 0.007963f
C662 B.n622 VSUBS 0.007963f
C663 B.n623 VSUBS 0.007963f
C664 B.n624 VSUBS 0.007963f
C665 B.n625 VSUBS 0.007963f
C666 B.n626 VSUBS 0.007963f
C667 B.n627 VSUBS 0.007963f
C668 B.n628 VSUBS 0.007963f
C669 B.n629 VSUBS 0.007963f
C670 B.n630 VSUBS 0.007963f
C671 B.n631 VSUBS 0.007963f
C672 B.n632 VSUBS 0.007963f
C673 B.n633 VSUBS 0.007963f
C674 B.n634 VSUBS 0.007963f
C675 B.n635 VSUBS 0.007963f
C676 B.n636 VSUBS 0.007963f
C677 B.n637 VSUBS 0.007963f
C678 B.n638 VSUBS 0.007963f
C679 B.n639 VSUBS 0.007963f
C680 B.n640 VSUBS 0.007963f
C681 B.n641 VSUBS 0.007963f
C682 B.n642 VSUBS 0.007963f
C683 B.n643 VSUBS 0.007963f
C684 B.n644 VSUBS 0.007963f
C685 B.n645 VSUBS 0.007963f
C686 B.n646 VSUBS 0.007963f
C687 B.n647 VSUBS 0.007963f
C688 B.n648 VSUBS 0.007963f
C689 B.n649 VSUBS 0.007963f
C690 B.n650 VSUBS 0.007963f
C691 B.n651 VSUBS 0.007963f
C692 B.n652 VSUBS 0.007963f
C693 B.n653 VSUBS 0.007963f
C694 B.n654 VSUBS 0.007963f
C695 B.n655 VSUBS 0.007963f
C696 B.n656 VSUBS 0.007963f
C697 B.n657 VSUBS 0.007963f
C698 B.n658 VSUBS 0.007963f
C699 B.n659 VSUBS 0.007963f
C700 B.n660 VSUBS 0.007963f
C701 B.n661 VSUBS 0.007963f
C702 B.n662 VSUBS 0.007963f
C703 B.n663 VSUBS 0.007963f
C704 B.n664 VSUBS 0.007963f
C705 B.n665 VSUBS 0.007963f
C706 B.n666 VSUBS 0.007963f
C707 B.n667 VSUBS 0.007963f
C708 B.n668 VSUBS 0.007963f
C709 B.n669 VSUBS 0.007963f
C710 B.n670 VSUBS 0.007963f
C711 B.n671 VSUBS 0.007963f
C712 B.n672 VSUBS 0.007963f
C713 B.n673 VSUBS 0.007963f
C714 B.n674 VSUBS 0.007963f
C715 B.n675 VSUBS 0.007963f
C716 B.n676 VSUBS 0.007963f
C717 B.n677 VSUBS 0.007963f
C718 B.n678 VSUBS 0.007963f
C719 B.n679 VSUBS 0.007963f
C720 B.n680 VSUBS 0.007963f
C721 B.n681 VSUBS 0.007963f
C722 B.n682 VSUBS 0.007963f
C723 B.n683 VSUBS 0.007963f
C724 B.n684 VSUBS 0.007963f
C725 B.n685 VSUBS 0.007963f
C726 B.n686 VSUBS 0.007963f
C727 B.n687 VSUBS 0.007963f
C728 B.n688 VSUBS 0.007963f
C729 B.n689 VSUBS 0.007963f
C730 B.n690 VSUBS 0.007963f
C731 B.n691 VSUBS 0.007963f
C732 B.n692 VSUBS 0.007963f
C733 B.n693 VSUBS 0.007963f
C734 B.n694 VSUBS 0.007963f
C735 B.n695 VSUBS 0.007963f
C736 B.n696 VSUBS 0.007963f
C737 B.n697 VSUBS 0.007963f
C738 B.n698 VSUBS 0.007963f
C739 B.n699 VSUBS 0.007963f
C740 B.n700 VSUBS 0.007963f
C741 B.n701 VSUBS 0.007963f
C742 B.n702 VSUBS 0.007963f
C743 B.n703 VSUBS 0.007963f
C744 B.n704 VSUBS 0.007963f
C745 B.n705 VSUBS 0.007963f
C746 B.n706 VSUBS 0.007963f
C747 B.n707 VSUBS 0.007963f
C748 B.n708 VSUBS 0.007963f
C749 B.n709 VSUBS 0.007963f
C750 B.n710 VSUBS 0.007963f
C751 B.n711 VSUBS 0.007963f
C752 B.n712 VSUBS 0.007963f
C753 B.n713 VSUBS 0.007963f
C754 B.n714 VSUBS 0.007963f
C755 B.n715 VSUBS 0.007963f
C756 B.n716 VSUBS 0.007963f
C757 B.n717 VSUBS 0.007963f
C758 B.n718 VSUBS 0.007963f
C759 B.n719 VSUBS 0.007963f
C760 B.n720 VSUBS 0.007963f
C761 B.n721 VSUBS 0.007963f
C762 B.n722 VSUBS 0.007963f
C763 B.n723 VSUBS 0.007963f
C764 B.n724 VSUBS 0.007963f
C765 B.n725 VSUBS 0.007963f
C766 B.n726 VSUBS 0.007963f
C767 B.n727 VSUBS 0.007963f
C768 B.n728 VSUBS 0.007963f
C769 B.n729 VSUBS 0.007963f
C770 B.n730 VSUBS 0.007963f
C771 B.n731 VSUBS 0.007963f
C772 B.n732 VSUBS 0.007963f
C773 B.n733 VSUBS 0.007963f
C774 B.n734 VSUBS 0.007963f
C775 B.n735 VSUBS 0.007963f
C776 B.n736 VSUBS 0.007963f
C777 B.n737 VSUBS 0.007963f
C778 B.n738 VSUBS 0.007963f
C779 B.n739 VSUBS 0.007963f
C780 B.n740 VSUBS 0.007963f
C781 B.n741 VSUBS 0.007963f
C782 B.n742 VSUBS 0.007963f
C783 B.n743 VSUBS 0.007963f
C784 B.n744 VSUBS 0.007963f
C785 B.n745 VSUBS 0.007963f
C786 B.n746 VSUBS 0.007963f
C787 B.n747 VSUBS 0.007963f
C788 B.n748 VSUBS 0.007963f
C789 B.n749 VSUBS 0.007963f
C790 B.n750 VSUBS 0.007963f
C791 B.n751 VSUBS 0.007963f
C792 B.n752 VSUBS 0.007963f
C793 B.n753 VSUBS 0.007963f
C794 B.n754 VSUBS 0.007963f
C795 B.n755 VSUBS 0.007963f
C796 B.n756 VSUBS 0.007963f
C797 B.n757 VSUBS 0.007963f
C798 B.n758 VSUBS 0.007963f
C799 B.n759 VSUBS 0.007963f
C800 B.n760 VSUBS 0.007963f
C801 B.n761 VSUBS 0.007963f
C802 B.n762 VSUBS 0.007963f
C803 B.n763 VSUBS 0.007963f
C804 B.n764 VSUBS 0.007963f
C805 B.n765 VSUBS 0.007963f
C806 B.n766 VSUBS 0.007963f
C807 B.n767 VSUBS 0.007963f
C808 B.n768 VSUBS 0.007963f
C809 B.n769 VSUBS 0.007963f
C810 B.n770 VSUBS 0.007963f
C811 B.n771 VSUBS 0.007963f
C812 B.n772 VSUBS 0.007963f
C813 B.n773 VSUBS 0.007963f
C814 B.n774 VSUBS 0.007963f
C815 B.n775 VSUBS 0.007963f
C816 B.n776 VSUBS 0.007963f
C817 B.n777 VSUBS 0.007963f
C818 B.n778 VSUBS 0.007963f
C819 B.n779 VSUBS 0.007963f
C820 B.n780 VSUBS 0.007963f
C821 B.n781 VSUBS 0.007963f
C822 B.n782 VSUBS 0.007963f
C823 B.n783 VSUBS 0.007963f
C824 B.n784 VSUBS 0.007963f
C825 B.n785 VSUBS 0.007963f
C826 B.n786 VSUBS 0.007963f
C827 B.n787 VSUBS 0.007963f
C828 B.n788 VSUBS 0.007963f
C829 B.n789 VSUBS 0.007963f
C830 B.n790 VSUBS 0.007963f
C831 B.n791 VSUBS 0.007963f
C832 B.n792 VSUBS 0.007963f
C833 B.n793 VSUBS 0.007963f
C834 B.n794 VSUBS 0.007963f
C835 B.n795 VSUBS 0.007963f
C836 B.n796 VSUBS 0.007963f
C837 B.n797 VSUBS 0.007963f
C838 B.n798 VSUBS 0.007963f
C839 B.n799 VSUBS 0.007963f
C840 B.n800 VSUBS 0.007963f
C841 B.n801 VSUBS 0.007963f
C842 B.n802 VSUBS 0.007963f
C843 B.n803 VSUBS 0.007963f
C844 B.n804 VSUBS 0.007963f
C845 B.n805 VSUBS 0.007963f
C846 B.n806 VSUBS 0.007963f
C847 B.n807 VSUBS 0.007963f
C848 B.n808 VSUBS 0.007963f
C849 B.n809 VSUBS 0.007963f
C850 B.n810 VSUBS 0.007963f
C851 B.n811 VSUBS 0.007963f
C852 B.n812 VSUBS 0.007963f
C853 B.n813 VSUBS 0.007963f
C854 B.n814 VSUBS 0.007963f
C855 B.n815 VSUBS 0.007963f
C856 B.n816 VSUBS 0.007963f
C857 B.n817 VSUBS 0.007963f
C858 B.n818 VSUBS 0.007963f
C859 B.n819 VSUBS 0.007963f
C860 B.n820 VSUBS 0.007963f
C861 B.n821 VSUBS 0.007963f
C862 B.n822 VSUBS 0.007963f
C863 B.n823 VSUBS 0.007963f
C864 B.n824 VSUBS 0.007963f
C865 B.n825 VSUBS 0.007963f
C866 B.n826 VSUBS 0.007963f
C867 B.n827 VSUBS 0.007963f
C868 B.n828 VSUBS 0.018476f
C869 B.n829 VSUBS 0.018476f
C870 B.n830 VSUBS 0.018999f
C871 B.n831 VSUBS 0.007963f
C872 B.n832 VSUBS 0.007963f
C873 B.n833 VSUBS 0.007963f
C874 B.n834 VSUBS 0.007963f
C875 B.n835 VSUBS 0.007963f
C876 B.n836 VSUBS 0.007963f
C877 B.n837 VSUBS 0.007963f
C878 B.n838 VSUBS 0.007963f
C879 B.n839 VSUBS 0.007963f
C880 B.n840 VSUBS 0.007963f
C881 B.n841 VSUBS 0.007963f
C882 B.n842 VSUBS 0.007963f
C883 B.n843 VSUBS 0.007963f
C884 B.n844 VSUBS 0.007963f
C885 B.n845 VSUBS 0.007963f
C886 B.n846 VSUBS 0.007963f
C887 B.n847 VSUBS 0.007963f
C888 B.n848 VSUBS 0.007963f
C889 B.n849 VSUBS 0.007963f
C890 B.n850 VSUBS 0.007963f
C891 B.n851 VSUBS 0.007963f
C892 B.n852 VSUBS 0.007963f
C893 B.n853 VSUBS 0.007963f
C894 B.n854 VSUBS 0.007963f
C895 B.n855 VSUBS 0.007963f
C896 B.n856 VSUBS 0.007963f
C897 B.n857 VSUBS 0.007963f
C898 B.n858 VSUBS 0.007963f
C899 B.n859 VSUBS 0.007963f
C900 B.n860 VSUBS 0.007963f
C901 B.n861 VSUBS 0.007963f
C902 B.n862 VSUBS 0.007963f
C903 B.n863 VSUBS 0.007963f
C904 B.n864 VSUBS 0.007963f
C905 B.n865 VSUBS 0.007963f
C906 B.n866 VSUBS 0.007963f
C907 B.n867 VSUBS 0.007963f
C908 B.n868 VSUBS 0.007963f
C909 B.n869 VSUBS 0.007963f
C910 B.n870 VSUBS 0.007963f
C911 B.n871 VSUBS 0.007963f
C912 B.n872 VSUBS 0.007963f
C913 B.n873 VSUBS 0.007963f
C914 B.n874 VSUBS 0.007963f
C915 B.n875 VSUBS 0.007963f
C916 B.n876 VSUBS 0.007963f
C917 B.n877 VSUBS 0.007963f
C918 B.n878 VSUBS 0.007963f
C919 B.n879 VSUBS 0.007963f
C920 B.n880 VSUBS 0.007963f
C921 B.n881 VSUBS 0.007963f
C922 B.n882 VSUBS 0.007963f
C923 B.n883 VSUBS 0.007963f
C924 B.n884 VSUBS 0.007963f
C925 B.n885 VSUBS 0.007963f
C926 B.n886 VSUBS 0.007963f
C927 B.n887 VSUBS 0.007963f
C928 B.n888 VSUBS 0.007963f
C929 B.n889 VSUBS 0.007963f
C930 B.n890 VSUBS 0.007963f
C931 B.n891 VSUBS 0.007963f
C932 B.n892 VSUBS 0.007963f
C933 B.n893 VSUBS 0.007963f
C934 B.n894 VSUBS 0.007963f
C935 B.n895 VSUBS 0.007963f
C936 B.n896 VSUBS 0.007963f
C937 B.n897 VSUBS 0.007963f
C938 B.n898 VSUBS 0.007963f
C939 B.n899 VSUBS 0.007963f
C940 B.n900 VSUBS 0.007963f
C941 B.n901 VSUBS 0.007963f
C942 B.n902 VSUBS 0.007963f
C943 B.n903 VSUBS 0.007963f
C944 B.n904 VSUBS 0.007963f
C945 B.n905 VSUBS 0.007963f
C946 B.n906 VSUBS 0.007963f
C947 B.n907 VSUBS 0.005504f
C948 B.n908 VSUBS 0.01845f
C949 B.n909 VSUBS 0.006441f
C950 B.n910 VSUBS 0.007963f
C951 B.n911 VSUBS 0.007963f
C952 B.n912 VSUBS 0.007963f
C953 B.n913 VSUBS 0.007963f
C954 B.n914 VSUBS 0.007963f
C955 B.n915 VSUBS 0.007963f
C956 B.n916 VSUBS 0.007963f
C957 B.n917 VSUBS 0.007963f
C958 B.n918 VSUBS 0.007963f
C959 B.n919 VSUBS 0.007963f
C960 B.n920 VSUBS 0.007963f
C961 B.n921 VSUBS 0.006441f
C962 B.n922 VSUBS 0.01845f
C963 B.n923 VSUBS 0.005504f
C964 B.n924 VSUBS 0.007963f
C965 B.n925 VSUBS 0.007963f
C966 B.n926 VSUBS 0.007963f
C967 B.n927 VSUBS 0.007963f
C968 B.n928 VSUBS 0.007963f
C969 B.n929 VSUBS 0.007963f
C970 B.n930 VSUBS 0.007963f
C971 B.n931 VSUBS 0.007963f
C972 B.n932 VSUBS 0.007963f
C973 B.n933 VSUBS 0.007963f
C974 B.n934 VSUBS 0.007963f
C975 B.n935 VSUBS 0.007963f
C976 B.n936 VSUBS 0.007963f
C977 B.n937 VSUBS 0.007963f
C978 B.n938 VSUBS 0.007963f
C979 B.n939 VSUBS 0.007963f
C980 B.n940 VSUBS 0.007963f
C981 B.n941 VSUBS 0.007963f
C982 B.n942 VSUBS 0.007963f
C983 B.n943 VSUBS 0.007963f
C984 B.n944 VSUBS 0.007963f
C985 B.n945 VSUBS 0.007963f
C986 B.n946 VSUBS 0.007963f
C987 B.n947 VSUBS 0.007963f
C988 B.n948 VSUBS 0.007963f
C989 B.n949 VSUBS 0.007963f
C990 B.n950 VSUBS 0.007963f
C991 B.n951 VSUBS 0.007963f
C992 B.n952 VSUBS 0.007963f
C993 B.n953 VSUBS 0.007963f
C994 B.n954 VSUBS 0.007963f
C995 B.n955 VSUBS 0.007963f
C996 B.n956 VSUBS 0.007963f
C997 B.n957 VSUBS 0.007963f
C998 B.n958 VSUBS 0.007963f
C999 B.n959 VSUBS 0.007963f
C1000 B.n960 VSUBS 0.007963f
C1001 B.n961 VSUBS 0.007963f
C1002 B.n962 VSUBS 0.007963f
C1003 B.n963 VSUBS 0.007963f
C1004 B.n964 VSUBS 0.007963f
C1005 B.n965 VSUBS 0.007963f
C1006 B.n966 VSUBS 0.007963f
C1007 B.n967 VSUBS 0.007963f
C1008 B.n968 VSUBS 0.007963f
C1009 B.n969 VSUBS 0.007963f
C1010 B.n970 VSUBS 0.007963f
C1011 B.n971 VSUBS 0.007963f
C1012 B.n972 VSUBS 0.007963f
C1013 B.n973 VSUBS 0.007963f
C1014 B.n974 VSUBS 0.007963f
C1015 B.n975 VSUBS 0.007963f
C1016 B.n976 VSUBS 0.007963f
C1017 B.n977 VSUBS 0.007963f
C1018 B.n978 VSUBS 0.007963f
C1019 B.n979 VSUBS 0.007963f
C1020 B.n980 VSUBS 0.007963f
C1021 B.n981 VSUBS 0.007963f
C1022 B.n982 VSUBS 0.007963f
C1023 B.n983 VSUBS 0.007963f
C1024 B.n984 VSUBS 0.007963f
C1025 B.n985 VSUBS 0.007963f
C1026 B.n986 VSUBS 0.007963f
C1027 B.n987 VSUBS 0.007963f
C1028 B.n988 VSUBS 0.007963f
C1029 B.n989 VSUBS 0.007963f
C1030 B.n990 VSUBS 0.007963f
C1031 B.n991 VSUBS 0.007963f
C1032 B.n992 VSUBS 0.007963f
C1033 B.n993 VSUBS 0.007963f
C1034 B.n994 VSUBS 0.007963f
C1035 B.n995 VSUBS 0.007963f
C1036 B.n996 VSUBS 0.007963f
C1037 B.n997 VSUBS 0.007963f
C1038 B.n998 VSUBS 0.007963f
C1039 B.n999 VSUBS 0.007963f
C1040 B.n1000 VSUBS 0.018999f
C1041 B.n1001 VSUBS 0.018476f
C1042 B.n1002 VSUBS 0.018476f
C1043 B.n1003 VSUBS 0.007963f
C1044 B.n1004 VSUBS 0.007963f
C1045 B.n1005 VSUBS 0.007963f
C1046 B.n1006 VSUBS 0.007963f
C1047 B.n1007 VSUBS 0.007963f
C1048 B.n1008 VSUBS 0.007963f
C1049 B.n1009 VSUBS 0.007963f
C1050 B.n1010 VSUBS 0.007963f
C1051 B.n1011 VSUBS 0.007963f
C1052 B.n1012 VSUBS 0.007963f
C1053 B.n1013 VSUBS 0.007963f
C1054 B.n1014 VSUBS 0.007963f
C1055 B.n1015 VSUBS 0.007963f
C1056 B.n1016 VSUBS 0.007963f
C1057 B.n1017 VSUBS 0.007963f
C1058 B.n1018 VSUBS 0.007963f
C1059 B.n1019 VSUBS 0.007963f
C1060 B.n1020 VSUBS 0.007963f
C1061 B.n1021 VSUBS 0.007963f
C1062 B.n1022 VSUBS 0.007963f
C1063 B.n1023 VSUBS 0.007963f
C1064 B.n1024 VSUBS 0.007963f
C1065 B.n1025 VSUBS 0.007963f
C1066 B.n1026 VSUBS 0.007963f
C1067 B.n1027 VSUBS 0.007963f
C1068 B.n1028 VSUBS 0.007963f
C1069 B.n1029 VSUBS 0.007963f
C1070 B.n1030 VSUBS 0.007963f
C1071 B.n1031 VSUBS 0.007963f
C1072 B.n1032 VSUBS 0.007963f
C1073 B.n1033 VSUBS 0.007963f
C1074 B.n1034 VSUBS 0.007963f
C1075 B.n1035 VSUBS 0.007963f
C1076 B.n1036 VSUBS 0.007963f
C1077 B.n1037 VSUBS 0.007963f
C1078 B.n1038 VSUBS 0.007963f
C1079 B.n1039 VSUBS 0.007963f
C1080 B.n1040 VSUBS 0.007963f
C1081 B.n1041 VSUBS 0.007963f
C1082 B.n1042 VSUBS 0.007963f
C1083 B.n1043 VSUBS 0.007963f
C1084 B.n1044 VSUBS 0.007963f
C1085 B.n1045 VSUBS 0.007963f
C1086 B.n1046 VSUBS 0.007963f
C1087 B.n1047 VSUBS 0.007963f
C1088 B.n1048 VSUBS 0.007963f
C1089 B.n1049 VSUBS 0.007963f
C1090 B.n1050 VSUBS 0.007963f
C1091 B.n1051 VSUBS 0.007963f
C1092 B.n1052 VSUBS 0.007963f
C1093 B.n1053 VSUBS 0.007963f
C1094 B.n1054 VSUBS 0.007963f
C1095 B.n1055 VSUBS 0.007963f
C1096 B.n1056 VSUBS 0.007963f
C1097 B.n1057 VSUBS 0.007963f
C1098 B.n1058 VSUBS 0.007963f
C1099 B.n1059 VSUBS 0.007963f
C1100 B.n1060 VSUBS 0.007963f
C1101 B.n1061 VSUBS 0.007963f
C1102 B.n1062 VSUBS 0.007963f
C1103 B.n1063 VSUBS 0.007963f
C1104 B.n1064 VSUBS 0.007963f
C1105 B.n1065 VSUBS 0.007963f
C1106 B.n1066 VSUBS 0.007963f
C1107 B.n1067 VSUBS 0.007963f
C1108 B.n1068 VSUBS 0.007963f
C1109 B.n1069 VSUBS 0.007963f
C1110 B.n1070 VSUBS 0.007963f
C1111 B.n1071 VSUBS 0.007963f
C1112 B.n1072 VSUBS 0.007963f
C1113 B.n1073 VSUBS 0.007963f
C1114 B.n1074 VSUBS 0.007963f
C1115 B.n1075 VSUBS 0.007963f
C1116 B.n1076 VSUBS 0.007963f
C1117 B.n1077 VSUBS 0.007963f
C1118 B.n1078 VSUBS 0.007963f
C1119 B.n1079 VSUBS 0.007963f
C1120 B.n1080 VSUBS 0.007963f
C1121 B.n1081 VSUBS 0.007963f
C1122 B.n1082 VSUBS 0.007963f
C1123 B.n1083 VSUBS 0.007963f
C1124 B.n1084 VSUBS 0.007963f
C1125 B.n1085 VSUBS 0.007963f
C1126 B.n1086 VSUBS 0.007963f
C1127 B.n1087 VSUBS 0.007963f
C1128 B.n1088 VSUBS 0.007963f
C1129 B.n1089 VSUBS 0.007963f
C1130 B.n1090 VSUBS 0.007963f
C1131 B.n1091 VSUBS 0.007963f
C1132 B.n1092 VSUBS 0.007963f
C1133 B.n1093 VSUBS 0.007963f
C1134 B.n1094 VSUBS 0.007963f
C1135 B.n1095 VSUBS 0.007963f
C1136 B.n1096 VSUBS 0.007963f
C1137 B.n1097 VSUBS 0.007963f
C1138 B.n1098 VSUBS 0.007963f
C1139 B.n1099 VSUBS 0.007963f
C1140 B.n1100 VSUBS 0.007963f
C1141 B.n1101 VSUBS 0.007963f
C1142 B.n1102 VSUBS 0.007963f
C1143 B.n1103 VSUBS 0.007963f
C1144 B.n1104 VSUBS 0.007963f
C1145 B.n1105 VSUBS 0.007963f
C1146 B.n1106 VSUBS 0.007963f
C1147 B.n1107 VSUBS 0.007963f
C1148 B.n1108 VSUBS 0.007963f
C1149 B.n1109 VSUBS 0.007963f
C1150 B.n1110 VSUBS 0.007963f
C1151 B.n1111 VSUBS 0.007963f
C1152 B.n1112 VSUBS 0.007963f
C1153 B.n1113 VSUBS 0.007963f
C1154 B.n1114 VSUBS 0.007963f
C1155 B.n1115 VSUBS 0.007963f
C1156 B.n1116 VSUBS 0.007963f
C1157 B.n1117 VSUBS 0.007963f
C1158 B.n1118 VSUBS 0.007963f
C1159 B.n1119 VSUBS 0.007963f
C1160 B.n1120 VSUBS 0.007963f
C1161 B.n1121 VSUBS 0.007963f
C1162 B.n1122 VSUBS 0.007963f
C1163 B.n1123 VSUBS 0.010392f
C1164 B.n1124 VSUBS 0.01107f
C1165 B.n1125 VSUBS 0.022013f
C1166 VDD2.n0 VSUBS 0.032299f
C1167 VDD2.n1 VSUBS 0.029972f
C1168 VDD2.n2 VSUBS 0.016106f
C1169 VDD2.n3 VSUBS 0.038068f
C1170 VDD2.n4 VSUBS 0.016579f
C1171 VDD2.n5 VSUBS 0.029972f
C1172 VDD2.n6 VSUBS 0.017053f
C1173 VDD2.n7 VSUBS 0.038068f
C1174 VDD2.n8 VSUBS 0.017053f
C1175 VDD2.n9 VSUBS 0.029972f
C1176 VDD2.n10 VSUBS 0.016106f
C1177 VDD2.n11 VSUBS 0.038068f
C1178 VDD2.n12 VSUBS 0.017053f
C1179 VDD2.n13 VSUBS 0.029972f
C1180 VDD2.n14 VSUBS 0.016106f
C1181 VDD2.n15 VSUBS 0.038068f
C1182 VDD2.n16 VSUBS 0.017053f
C1183 VDD2.n17 VSUBS 0.029972f
C1184 VDD2.n18 VSUBS 0.016106f
C1185 VDD2.n19 VSUBS 0.038068f
C1186 VDD2.n20 VSUBS 0.017053f
C1187 VDD2.n21 VSUBS 0.029972f
C1188 VDD2.n22 VSUBS 0.016106f
C1189 VDD2.n23 VSUBS 0.038068f
C1190 VDD2.n24 VSUBS 0.017053f
C1191 VDD2.n25 VSUBS 1.97909f
C1192 VDD2.n26 VSUBS 0.016106f
C1193 VDD2.t0 VSUBS 0.081532f
C1194 VDD2.n27 VSUBS 0.215521f
C1195 VDD2.n28 VSUBS 0.024217f
C1196 VDD2.n29 VSUBS 0.028551f
C1197 VDD2.n30 VSUBS 0.038068f
C1198 VDD2.n31 VSUBS 0.017053f
C1199 VDD2.n32 VSUBS 0.016106f
C1200 VDD2.n33 VSUBS 0.029972f
C1201 VDD2.n34 VSUBS 0.029972f
C1202 VDD2.n35 VSUBS 0.016106f
C1203 VDD2.n36 VSUBS 0.017053f
C1204 VDD2.n37 VSUBS 0.038068f
C1205 VDD2.n38 VSUBS 0.038068f
C1206 VDD2.n39 VSUBS 0.017053f
C1207 VDD2.n40 VSUBS 0.016106f
C1208 VDD2.n41 VSUBS 0.029972f
C1209 VDD2.n42 VSUBS 0.029972f
C1210 VDD2.n43 VSUBS 0.016106f
C1211 VDD2.n44 VSUBS 0.017053f
C1212 VDD2.n45 VSUBS 0.038068f
C1213 VDD2.n46 VSUBS 0.038068f
C1214 VDD2.n47 VSUBS 0.017053f
C1215 VDD2.n48 VSUBS 0.016106f
C1216 VDD2.n49 VSUBS 0.029972f
C1217 VDD2.n50 VSUBS 0.029972f
C1218 VDD2.n51 VSUBS 0.016106f
C1219 VDD2.n52 VSUBS 0.017053f
C1220 VDD2.n53 VSUBS 0.038068f
C1221 VDD2.n54 VSUBS 0.038068f
C1222 VDD2.n55 VSUBS 0.017053f
C1223 VDD2.n56 VSUBS 0.016106f
C1224 VDD2.n57 VSUBS 0.029972f
C1225 VDD2.n58 VSUBS 0.029972f
C1226 VDD2.n59 VSUBS 0.016106f
C1227 VDD2.n60 VSUBS 0.017053f
C1228 VDD2.n61 VSUBS 0.038068f
C1229 VDD2.n62 VSUBS 0.038068f
C1230 VDD2.n63 VSUBS 0.017053f
C1231 VDD2.n64 VSUBS 0.016106f
C1232 VDD2.n65 VSUBS 0.029972f
C1233 VDD2.n66 VSUBS 0.029972f
C1234 VDD2.n67 VSUBS 0.016106f
C1235 VDD2.n68 VSUBS 0.016106f
C1236 VDD2.n69 VSUBS 0.017053f
C1237 VDD2.n70 VSUBS 0.038068f
C1238 VDD2.n71 VSUBS 0.038068f
C1239 VDD2.n72 VSUBS 0.038068f
C1240 VDD2.n73 VSUBS 0.016579f
C1241 VDD2.n74 VSUBS 0.016106f
C1242 VDD2.n75 VSUBS 0.029972f
C1243 VDD2.n76 VSUBS 0.029972f
C1244 VDD2.n77 VSUBS 0.016106f
C1245 VDD2.n78 VSUBS 0.017053f
C1246 VDD2.n79 VSUBS 0.038068f
C1247 VDD2.n80 VSUBS 0.090001f
C1248 VDD2.n81 VSUBS 0.017053f
C1249 VDD2.n82 VSUBS 0.016106f
C1250 VDD2.n83 VSUBS 0.074192f
C1251 VDD2.n84 VSUBS 0.093182f
C1252 VDD2.t4 VSUBS 0.366642f
C1253 VDD2.t9 VSUBS 0.366642f
C1254 VDD2.n85 VSUBS 2.99817f
C1255 VDD2.n86 VSUBS 1.38417f
C1256 VDD2.t2 VSUBS 0.366642f
C1257 VDD2.t8 VSUBS 0.366642f
C1258 VDD2.n87 VSUBS 3.04024f
C1259 VDD2.n88 VSUBS 4.85631f
C1260 VDD2.n89 VSUBS 0.032299f
C1261 VDD2.n90 VSUBS 0.029972f
C1262 VDD2.n91 VSUBS 0.016106f
C1263 VDD2.n92 VSUBS 0.038068f
C1264 VDD2.n93 VSUBS 0.016579f
C1265 VDD2.n94 VSUBS 0.029972f
C1266 VDD2.n95 VSUBS 0.016579f
C1267 VDD2.n96 VSUBS 0.016106f
C1268 VDD2.n97 VSUBS 0.038068f
C1269 VDD2.n98 VSUBS 0.038068f
C1270 VDD2.n99 VSUBS 0.017053f
C1271 VDD2.n100 VSUBS 0.029972f
C1272 VDD2.n101 VSUBS 0.016106f
C1273 VDD2.n102 VSUBS 0.038068f
C1274 VDD2.n103 VSUBS 0.017053f
C1275 VDD2.n104 VSUBS 0.029972f
C1276 VDD2.n105 VSUBS 0.016106f
C1277 VDD2.n106 VSUBS 0.038068f
C1278 VDD2.n107 VSUBS 0.017053f
C1279 VDD2.n108 VSUBS 0.029972f
C1280 VDD2.n109 VSUBS 0.016106f
C1281 VDD2.n110 VSUBS 0.038068f
C1282 VDD2.n111 VSUBS 0.017053f
C1283 VDD2.n112 VSUBS 0.029972f
C1284 VDD2.n113 VSUBS 0.016106f
C1285 VDD2.n114 VSUBS 0.038068f
C1286 VDD2.n115 VSUBS 0.017053f
C1287 VDD2.n116 VSUBS 1.97909f
C1288 VDD2.n117 VSUBS 0.016106f
C1289 VDD2.t7 VSUBS 0.081532f
C1290 VDD2.n118 VSUBS 0.215521f
C1291 VDD2.n119 VSUBS 0.024217f
C1292 VDD2.n120 VSUBS 0.028551f
C1293 VDD2.n121 VSUBS 0.038068f
C1294 VDD2.n122 VSUBS 0.017053f
C1295 VDD2.n123 VSUBS 0.016106f
C1296 VDD2.n124 VSUBS 0.029972f
C1297 VDD2.n125 VSUBS 0.029972f
C1298 VDD2.n126 VSUBS 0.016106f
C1299 VDD2.n127 VSUBS 0.017053f
C1300 VDD2.n128 VSUBS 0.038068f
C1301 VDD2.n129 VSUBS 0.038068f
C1302 VDD2.n130 VSUBS 0.017053f
C1303 VDD2.n131 VSUBS 0.016106f
C1304 VDD2.n132 VSUBS 0.029972f
C1305 VDD2.n133 VSUBS 0.029972f
C1306 VDD2.n134 VSUBS 0.016106f
C1307 VDD2.n135 VSUBS 0.017053f
C1308 VDD2.n136 VSUBS 0.038068f
C1309 VDD2.n137 VSUBS 0.038068f
C1310 VDD2.n138 VSUBS 0.017053f
C1311 VDD2.n139 VSUBS 0.016106f
C1312 VDD2.n140 VSUBS 0.029972f
C1313 VDD2.n141 VSUBS 0.029972f
C1314 VDD2.n142 VSUBS 0.016106f
C1315 VDD2.n143 VSUBS 0.017053f
C1316 VDD2.n144 VSUBS 0.038068f
C1317 VDD2.n145 VSUBS 0.038068f
C1318 VDD2.n146 VSUBS 0.017053f
C1319 VDD2.n147 VSUBS 0.016106f
C1320 VDD2.n148 VSUBS 0.029972f
C1321 VDD2.n149 VSUBS 0.029972f
C1322 VDD2.n150 VSUBS 0.016106f
C1323 VDD2.n151 VSUBS 0.017053f
C1324 VDD2.n152 VSUBS 0.038068f
C1325 VDD2.n153 VSUBS 0.038068f
C1326 VDD2.n154 VSUBS 0.017053f
C1327 VDD2.n155 VSUBS 0.016106f
C1328 VDD2.n156 VSUBS 0.029972f
C1329 VDD2.n157 VSUBS 0.029972f
C1330 VDD2.n158 VSUBS 0.016106f
C1331 VDD2.n159 VSUBS 0.017053f
C1332 VDD2.n160 VSUBS 0.038068f
C1333 VDD2.n161 VSUBS 0.038068f
C1334 VDD2.n162 VSUBS 0.017053f
C1335 VDD2.n163 VSUBS 0.016106f
C1336 VDD2.n164 VSUBS 0.029972f
C1337 VDD2.n165 VSUBS 0.029972f
C1338 VDD2.n166 VSUBS 0.016106f
C1339 VDD2.n167 VSUBS 0.017053f
C1340 VDD2.n168 VSUBS 0.038068f
C1341 VDD2.n169 VSUBS 0.090001f
C1342 VDD2.n170 VSUBS 0.017053f
C1343 VDD2.n171 VSUBS 0.016106f
C1344 VDD2.n172 VSUBS 0.074192f
C1345 VDD2.n173 VSUBS 0.06597f
C1346 VDD2.n174 VSUBS 4.38405f
C1347 VDD2.t6 VSUBS 0.366642f
C1348 VDD2.t1 VSUBS 0.366642f
C1349 VDD2.n175 VSUBS 2.99818f
C1350 VDD2.n176 VSUBS 1.01049f
C1351 VDD2.t5 VSUBS 0.366642f
C1352 VDD2.t3 VSUBS 0.366642f
C1353 VDD2.n177 VSUBS 3.04018f
C1354 VN.n0 VSUBS 0.039553f
C1355 VN.t1 VSUBS 3.46423f
C1356 VN.n1 VSUBS 0.039005f
C1357 VN.n2 VSUBS 0.021034f
C1358 VN.n3 VSUBS 0.039005f
C1359 VN.n4 VSUBS 0.021034f
C1360 VN.t7 VSUBS 3.46423f
C1361 VN.n5 VSUBS 0.039005f
C1362 VN.n6 VSUBS 0.021034f
C1363 VN.n7 VSUBS 0.039005f
C1364 VN.n8 VSUBS 0.021034f
C1365 VN.t0 VSUBS 3.46423f
C1366 VN.n9 VSUBS 0.039005f
C1367 VN.n10 VSUBS 0.021034f
C1368 VN.n11 VSUBS 0.039005f
C1369 VN.n12 VSUBS 0.277554f
C1370 VN.t5 VSUBS 3.46423f
C1371 VN.t9 VSUBS 3.8071f
C1372 VN.n13 VSUBS 1.21361f
C1373 VN.n14 VSUBS 1.27341f
C1374 VN.n15 VSUBS 0.027837f
C1375 VN.n16 VSUBS 0.039005f
C1376 VN.n17 VSUBS 0.021034f
C1377 VN.n18 VSUBS 0.021034f
C1378 VN.n19 VSUBS 0.021034f
C1379 VN.n20 VSUBS 0.038211f
C1380 VN.n21 VSUBS 0.020143f
C1381 VN.n22 VSUBS 0.041803f
C1382 VN.n23 VSUBS 0.021034f
C1383 VN.n24 VSUBS 0.021034f
C1384 VN.n25 VSUBS 0.021034f
C1385 VN.n26 VSUBS 0.039005f
C1386 VN.n27 VSUBS 1.21916f
C1387 VN.n28 VSUBS 0.039005f
C1388 VN.n29 VSUBS 0.021034f
C1389 VN.n30 VSUBS 0.021034f
C1390 VN.n31 VSUBS 0.021034f
C1391 VN.n32 VSUBS 0.041803f
C1392 VN.n33 VSUBS 0.020143f
C1393 VN.n34 VSUBS 0.038211f
C1394 VN.n35 VSUBS 0.021034f
C1395 VN.n36 VSUBS 0.021034f
C1396 VN.n37 VSUBS 0.021034f
C1397 VN.n38 VSUBS 0.039005f
C1398 VN.n39 VSUBS 0.027837f
C1399 VN.n40 VSUBS 1.19941f
C1400 VN.n41 VSUBS 0.030918f
C1401 VN.n42 VSUBS 0.021034f
C1402 VN.n43 VSUBS 0.021034f
C1403 VN.n44 VSUBS 0.021034f
C1404 VN.n45 VSUBS 0.039005f
C1405 VN.n46 VSUBS 0.034359f
C1406 VN.n47 VSUBS 0.026793f
C1407 VN.n48 VSUBS 0.021034f
C1408 VN.n49 VSUBS 0.021034f
C1409 VN.n50 VSUBS 0.021034f
C1410 VN.n51 VSUBS 0.039005f
C1411 VN.n52 VSUBS 0.035924f
C1412 VN.n53 VSUBS 1.28987f
C1413 VN.n54 VSUBS 0.065709f
C1414 VN.n55 VSUBS 0.039553f
C1415 VN.t2 VSUBS 3.46423f
C1416 VN.n56 VSUBS 0.039005f
C1417 VN.n57 VSUBS 0.021034f
C1418 VN.n58 VSUBS 0.039005f
C1419 VN.n59 VSUBS 0.021034f
C1420 VN.t3 VSUBS 3.46423f
C1421 VN.n60 VSUBS 0.039005f
C1422 VN.n61 VSUBS 0.021034f
C1423 VN.n62 VSUBS 0.039005f
C1424 VN.n63 VSUBS 0.021034f
C1425 VN.t8 VSUBS 3.46423f
C1426 VN.n64 VSUBS 0.039005f
C1427 VN.n65 VSUBS 0.021034f
C1428 VN.n66 VSUBS 0.039005f
C1429 VN.n67 VSUBS 0.277554f
C1430 VN.t4 VSUBS 3.46423f
C1431 VN.t6 VSUBS 3.8071f
C1432 VN.n68 VSUBS 1.21361f
C1433 VN.n69 VSUBS 1.27341f
C1434 VN.n70 VSUBS 0.027837f
C1435 VN.n71 VSUBS 0.039005f
C1436 VN.n72 VSUBS 0.021034f
C1437 VN.n73 VSUBS 0.021034f
C1438 VN.n74 VSUBS 0.021034f
C1439 VN.n75 VSUBS 0.038211f
C1440 VN.n76 VSUBS 0.020143f
C1441 VN.n77 VSUBS 0.041803f
C1442 VN.n78 VSUBS 0.021034f
C1443 VN.n79 VSUBS 0.021034f
C1444 VN.n80 VSUBS 0.021034f
C1445 VN.n81 VSUBS 0.039005f
C1446 VN.n82 VSUBS 1.21916f
C1447 VN.n83 VSUBS 0.039005f
C1448 VN.n84 VSUBS 0.021034f
C1449 VN.n85 VSUBS 0.021034f
C1450 VN.n86 VSUBS 0.021034f
C1451 VN.n87 VSUBS 0.041803f
C1452 VN.n88 VSUBS 0.020143f
C1453 VN.n89 VSUBS 0.038211f
C1454 VN.n90 VSUBS 0.021034f
C1455 VN.n91 VSUBS 0.021034f
C1456 VN.n92 VSUBS 0.021034f
C1457 VN.n93 VSUBS 0.039005f
C1458 VN.n94 VSUBS 0.027837f
C1459 VN.n95 VSUBS 1.19941f
C1460 VN.n96 VSUBS 0.030918f
C1461 VN.n97 VSUBS 0.021034f
C1462 VN.n98 VSUBS 0.021034f
C1463 VN.n99 VSUBS 0.021034f
C1464 VN.n100 VSUBS 0.039005f
C1465 VN.n101 VSUBS 0.034359f
C1466 VN.n102 VSUBS 0.026793f
C1467 VN.n103 VSUBS 0.021034f
C1468 VN.n104 VSUBS 0.021034f
C1469 VN.n105 VSUBS 0.021034f
C1470 VN.n106 VSUBS 0.039005f
C1471 VN.n107 VSUBS 0.035924f
C1472 VN.n108 VSUBS 1.28987f
C1473 VN.n109 VSUBS 1.67144f
C1474 VDD1.n0 VSUBS 0.03229f
C1475 VDD1.n1 VSUBS 0.029963f
C1476 VDD1.n2 VSUBS 0.016101f
C1477 VDD1.n3 VSUBS 0.038057f
C1478 VDD1.n4 VSUBS 0.016575f
C1479 VDD1.n5 VSUBS 0.029963f
C1480 VDD1.n6 VSUBS 0.016575f
C1481 VDD1.n7 VSUBS 0.016101f
C1482 VDD1.n8 VSUBS 0.038057f
C1483 VDD1.n9 VSUBS 0.038057f
C1484 VDD1.n10 VSUBS 0.017048f
C1485 VDD1.n11 VSUBS 0.029963f
C1486 VDD1.n12 VSUBS 0.016101f
C1487 VDD1.n13 VSUBS 0.038057f
C1488 VDD1.n14 VSUBS 0.017048f
C1489 VDD1.n15 VSUBS 0.029963f
C1490 VDD1.n16 VSUBS 0.016101f
C1491 VDD1.n17 VSUBS 0.038057f
C1492 VDD1.n18 VSUBS 0.017048f
C1493 VDD1.n19 VSUBS 0.029963f
C1494 VDD1.n20 VSUBS 0.016101f
C1495 VDD1.n21 VSUBS 0.038057f
C1496 VDD1.n22 VSUBS 0.017048f
C1497 VDD1.n23 VSUBS 0.029963f
C1498 VDD1.n24 VSUBS 0.016101f
C1499 VDD1.n25 VSUBS 0.038057f
C1500 VDD1.n26 VSUBS 0.017048f
C1501 VDD1.n27 VSUBS 1.97852f
C1502 VDD1.n28 VSUBS 0.016101f
C1503 VDD1.t3 VSUBS 0.081508f
C1504 VDD1.n29 VSUBS 0.215459f
C1505 VDD1.n30 VSUBS 0.02421f
C1506 VDD1.n31 VSUBS 0.028543f
C1507 VDD1.n32 VSUBS 0.038057f
C1508 VDD1.n33 VSUBS 0.017048f
C1509 VDD1.n34 VSUBS 0.016101f
C1510 VDD1.n35 VSUBS 0.029963f
C1511 VDD1.n36 VSUBS 0.029963f
C1512 VDD1.n37 VSUBS 0.016101f
C1513 VDD1.n38 VSUBS 0.017048f
C1514 VDD1.n39 VSUBS 0.038057f
C1515 VDD1.n40 VSUBS 0.038057f
C1516 VDD1.n41 VSUBS 0.017048f
C1517 VDD1.n42 VSUBS 0.016101f
C1518 VDD1.n43 VSUBS 0.029963f
C1519 VDD1.n44 VSUBS 0.029963f
C1520 VDD1.n45 VSUBS 0.016101f
C1521 VDD1.n46 VSUBS 0.017048f
C1522 VDD1.n47 VSUBS 0.038057f
C1523 VDD1.n48 VSUBS 0.038057f
C1524 VDD1.n49 VSUBS 0.017048f
C1525 VDD1.n50 VSUBS 0.016101f
C1526 VDD1.n51 VSUBS 0.029963f
C1527 VDD1.n52 VSUBS 0.029963f
C1528 VDD1.n53 VSUBS 0.016101f
C1529 VDD1.n54 VSUBS 0.017048f
C1530 VDD1.n55 VSUBS 0.038057f
C1531 VDD1.n56 VSUBS 0.038057f
C1532 VDD1.n57 VSUBS 0.017048f
C1533 VDD1.n58 VSUBS 0.016101f
C1534 VDD1.n59 VSUBS 0.029963f
C1535 VDD1.n60 VSUBS 0.029963f
C1536 VDD1.n61 VSUBS 0.016101f
C1537 VDD1.n62 VSUBS 0.017048f
C1538 VDD1.n63 VSUBS 0.038057f
C1539 VDD1.n64 VSUBS 0.038057f
C1540 VDD1.n65 VSUBS 0.017048f
C1541 VDD1.n66 VSUBS 0.016101f
C1542 VDD1.n67 VSUBS 0.029963f
C1543 VDD1.n68 VSUBS 0.029963f
C1544 VDD1.n69 VSUBS 0.016101f
C1545 VDD1.n70 VSUBS 0.017048f
C1546 VDD1.n71 VSUBS 0.038057f
C1547 VDD1.n72 VSUBS 0.038057f
C1548 VDD1.n73 VSUBS 0.017048f
C1549 VDD1.n74 VSUBS 0.016101f
C1550 VDD1.n75 VSUBS 0.029963f
C1551 VDD1.n76 VSUBS 0.029963f
C1552 VDD1.n77 VSUBS 0.016101f
C1553 VDD1.n78 VSUBS 0.017048f
C1554 VDD1.n79 VSUBS 0.038057f
C1555 VDD1.n80 VSUBS 0.089975f
C1556 VDD1.n81 VSUBS 0.017048f
C1557 VDD1.n82 VSUBS 0.016101f
C1558 VDD1.n83 VSUBS 0.074171f
C1559 VDD1.n84 VSUBS 0.093156f
C1560 VDD1.t4 VSUBS 0.366536f
C1561 VDD1.t5 VSUBS 0.366536f
C1562 VDD1.n85 VSUBS 2.99732f
C1563 VDD1.n86 VSUBS 1.39391f
C1564 VDD1.n87 VSUBS 0.03229f
C1565 VDD1.n88 VSUBS 0.029963f
C1566 VDD1.n89 VSUBS 0.016101f
C1567 VDD1.n90 VSUBS 0.038057f
C1568 VDD1.n91 VSUBS 0.016575f
C1569 VDD1.n92 VSUBS 0.029963f
C1570 VDD1.n93 VSUBS 0.017048f
C1571 VDD1.n94 VSUBS 0.038057f
C1572 VDD1.n95 VSUBS 0.017048f
C1573 VDD1.n96 VSUBS 0.029963f
C1574 VDD1.n97 VSUBS 0.016101f
C1575 VDD1.n98 VSUBS 0.038057f
C1576 VDD1.n99 VSUBS 0.017048f
C1577 VDD1.n100 VSUBS 0.029963f
C1578 VDD1.n101 VSUBS 0.016101f
C1579 VDD1.n102 VSUBS 0.038057f
C1580 VDD1.n103 VSUBS 0.017048f
C1581 VDD1.n104 VSUBS 0.029963f
C1582 VDD1.n105 VSUBS 0.016101f
C1583 VDD1.n106 VSUBS 0.038057f
C1584 VDD1.n107 VSUBS 0.017048f
C1585 VDD1.n108 VSUBS 0.029963f
C1586 VDD1.n109 VSUBS 0.016101f
C1587 VDD1.n110 VSUBS 0.038057f
C1588 VDD1.n111 VSUBS 0.017048f
C1589 VDD1.n112 VSUBS 1.97852f
C1590 VDD1.n113 VSUBS 0.016101f
C1591 VDD1.t9 VSUBS 0.081508f
C1592 VDD1.n114 VSUBS 0.215459f
C1593 VDD1.n115 VSUBS 0.02421f
C1594 VDD1.n116 VSUBS 0.028543f
C1595 VDD1.n117 VSUBS 0.038057f
C1596 VDD1.n118 VSUBS 0.017048f
C1597 VDD1.n119 VSUBS 0.016101f
C1598 VDD1.n120 VSUBS 0.029963f
C1599 VDD1.n121 VSUBS 0.029963f
C1600 VDD1.n122 VSUBS 0.016101f
C1601 VDD1.n123 VSUBS 0.017048f
C1602 VDD1.n124 VSUBS 0.038057f
C1603 VDD1.n125 VSUBS 0.038057f
C1604 VDD1.n126 VSUBS 0.017048f
C1605 VDD1.n127 VSUBS 0.016101f
C1606 VDD1.n128 VSUBS 0.029963f
C1607 VDD1.n129 VSUBS 0.029963f
C1608 VDD1.n130 VSUBS 0.016101f
C1609 VDD1.n131 VSUBS 0.017048f
C1610 VDD1.n132 VSUBS 0.038057f
C1611 VDD1.n133 VSUBS 0.038057f
C1612 VDD1.n134 VSUBS 0.017048f
C1613 VDD1.n135 VSUBS 0.016101f
C1614 VDD1.n136 VSUBS 0.029963f
C1615 VDD1.n137 VSUBS 0.029963f
C1616 VDD1.n138 VSUBS 0.016101f
C1617 VDD1.n139 VSUBS 0.017048f
C1618 VDD1.n140 VSUBS 0.038057f
C1619 VDD1.n141 VSUBS 0.038057f
C1620 VDD1.n142 VSUBS 0.017048f
C1621 VDD1.n143 VSUBS 0.016101f
C1622 VDD1.n144 VSUBS 0.029963f
C1623 VDD1.n145 VSUBS 0.029963f
C1624 VDD1.n146 VSUBS 0.016101f
C1625 VDD1.n147 VSUBS 0.017048f
C1626 VDD1.n148 VSUBS 0.038057f
C1627 VDD1.n149 VSUBS 0.038057f
C1628 VDD1.n150 VSUBS 0.017048f
C1629 VDD1.n151 VSUBS 0.016101f
C1630 VDD1.n152 VSUBS 0.029963f
C1631 VDD1.n153 VSUBS 0.029963f
C1632 VDD1.n154 VSUBS 0.016101f
C1633 VDD1.n155 VSUBS 0.016101f
C1634 VDD1.n156 VSUBS 0.017048f
C1635 VDD1.n157 VSUBS 0.038057f
C1636 VDD1.n158 VSUBS 0.038057f
C1637 VDD1.n159 VSUBS 0.038057f
C1638 VDD1.n160 VSUBS 0.016575f
C1639 VDD1.n161 VSUBS 0.016101f
C1640 VDD1.n162 VSUBS 0.029963f
C1641 VDD1.n163 VSUBS 0.029963f
C1642 VDD1.n164 VSUBS 0.016101f
C1643 VDD1.n165 VSUBS 0.017048f
C1644 VDD1.n166 VSUBS 0.038057f
C1645 VDD1.n167 VSUBS 0.089975f
C1646 VDD1.n168 VSUBS 0.017048f
C1647 VDD1.n169 VSUBS 0.016101f
C1648 VDD1.n170 VSUBS 0.074171f
C1649 VDD1.n171 VSUBS 0.093156f
C1650 VDD1.t6 VSUBS 0.366536f
C1651 VDD1.t2 VSUBS 0.366536f
C1652 VDD1.n172 VSUBS 2.99731f
C1653 VDD1.n173 VSUBS 1.38377f
C1654 VDD1.t1 VSUBS 0.366536f
C1655 VDD1.t8 VSUBS 0.366536f
C1656 VDD1.n174 VSUBS 3.03937f
C1657 VDD1.n175 VSUBS 5.05038f
C1658 VDD1.t7 VSUBS 0.366536f
C1659 VDD1.t0 VSUBS 0.366536f
C1660 VDD1.n176 VSUBS 2.99731f
C1661 VDD1.n177 VSUBS 5.07332f
C1662 VTAIL.t2 VSUBS 0.352887f
C1663 VTAIL.t18 VSUBS 0.352887f
C1664 VTAIL.n0 VSUBS 2.72459f
C1665 VTAIL.n1 VSUBS 1.13815f
C1666 VTAIL.n2 VSUBS 0.031088f
C1667 VTAIL.n3 VSUBS 0.028848f
C1668 VTAIL.n4 VSUBS 0.015502f
C1669 VTAIL.n5 VSUBS 0.03664f
C1670 VTAIL.n6 VSUBS 0.015957f
C1671 VTAIL.n7 VSUBS 0.028848f
C1672 VTAIL.n8 VSUBS 0.016413f
C1673 VTAIL.n9 VSUBS 0.03664f
C1674 VTAIL.n10 VSUBS 0.016413f
C1675 VTAIL.n11 VSUBS 0.028848f
C1676 VTAIL.n12 VSUBS 0.015502f
C1677 VTAIL.n13 VSUBS 0.03664f
C1678 VTAIL.n14 VSUBS 0.016413f
C1679 VTAIL.n15 VSUBS 0.028848f
C1680 VTAIL.n16 VSUBS 0.015502f
C1681 VTAIL.n17 VSUBS 0.03664f
C1682 VTAIL.n18 VSUBS 0.016413f
C1683 VTAIL.n19 VSUBS 0.028848f
C1684 VTAIL.n20 VSUBS 0.015502f
C1685 VTAIL.n21 VSUBS 0.03664f
C1686 VTAIL.n22 VSUBS 0.016413f
C1687 VTAIL.n23 VSUBS 0.028848f
C1688 VTAIL.n24 VSUBS 0.015502f
C1689 VTAIL.n25 VSUBS 0.03664f
C1690 VTAIL.n26 VSUBS 0.016413f
C1691 VTAIL.n27 VSUBS 1.90484f
C1692 VTAIL.n28 VSUBS 0.015502f
C1693 VTAIL.t8 VSUBS 0.078473f
C1694 VTAIL.n29 VSUBS 0.207435f
C1695 VTAIL.n30 VSUBS 0.023309f
C1696 VTAIL.n31 VSUBS 0.02748f
C1697 VTAIL.n32 VSUBS 0.03664f
C1698 VTAIL.n33 VSUBS 0.016413f
C1699 VTAIL.n34 VSUBS 0.015502f
C1700 VTAIL.n35 VSUBS 0.028848f
C1701 VTAIL.n36 VSUBS 0.028848f
C1702 VTAIL.n37 VSUBS 0.015502f
C1703 VTAIL.n38 VSUBS 0.016413f
C1704 VTAIL.n39 VSUBS 0.03664f
C1705 VTAIL.n40 VSUBS 0.03664f
C1706 VTAIL.n41 VSUBS 0.016413f
C1707 VTAIL.n42 VSUBS 0.015502f
C1708 VTAIL.n43 VSUBS 0.028848f
C1709 VTAIL.n44 VSUBS 0.028848f
C1710 VTAIL.n45 VSUBS 0.015502f
C1711 VTAIL.n46 VSUBS 0.016413f
C1712 VTAIL.n47 VSUBS 0.03664f
C1713 VTAIL.n48 VSUBS 0.03664f
C1714 VTAIL.n49 VSUBS 0.016413f
C1715 VTAIL.n50 VSUBS 0.015502f
C1716 VTAIL.n51 VSUBS 0.028848f
C1717 VTAIL.n52 VSUBS 0.028848f
C1718 VTAIL.n53 VSUBS 0.015502f
C1719 VTAIL.n54 VSUBS 0.016413f
C1720 VTAIL.n55 VSUBS 0.03664f
C1721 VTAIL.n56 VSUBS 0.03664f
C1722 VTAIL.n57 VSUBS 0.016413f
C1723 VTAIL.n58 VSUBS 0.015502f
C1724 VTAIL.n59 VSUBS 0.028848f
C1725 VTAIL.n60 VSUBS 0.028848f
C1726 VTAIL.n61 VSUBS 0.015502f
C1727 VTAIL.n62 VSUBS 0.016413f
C1728 VTAIL.n63 VSUBS 0.03664f
C1729 VTAIL.n64 VSUBS 0.03664f
C1730 VTAIL.n65 VSUBS 0.016413f
C1731 VTAIL.n66 VSUBS 0.015502f
C1732 VTAIL.n67 VSUBS 0.028848f
C1733 VTAIL.n68 VSUBS 0.028848f
C1734 VTAIL.n69 VSUBS 0.015502f
C1735 VTAIL.n70 VSUBS 0.015502f
C1736 VTAIL.n71 VSUBS 0.016413f
C1737 VTAIL.n72 VSUBS 0.03664f
C1738 VTAIL.n73 VSUBS 0.03664f
C1739 VTAIL.n74 VSUBS 0.03664f
C1740 VTAIL.n75 VSUBS 0.015957f
C1741 VTAIL.n76 VSUBS 0.015502f
C1742 VTAIL.n77 VSUBS 0.028848f
C1743 VTAIL.n78 VSUBS 0.028848f
C1744 VTAIL.n79 VSUBS 0.015502f
C1745 VTAIL.n80 VSUBS 0.016413f
C1746 VTAIL.n81 VSUBS 0.03664f
C1747 VTAIL.n82 VSUBS 0.086624f
C1748 VTAIL.n83 VSUBS 0.016413f
C1749 VTAIL.n84 VSUBS 0.015502f
C1750 VTAIL.n85 VSUBS 0.071409f
C1751 VTAIL.n86 VSUBS 0.043611f
C1752 VTAIL.n87 VSUBS 0.57702f
C1753 VTAIL.t17 VSUBS 0.352887f
C1754 VTAIL.t13 VSUBS 0.352887f
C1755 VTAIL.n88 VSUBS 2.72459f
C1756 VTAIL.n89 VSUBS 1.34209f
C1757 VTAIL.t16 VSUBS 0.352887f
C1758 VTAIL.t10 VSUBS 0.352887f
C1759 VTAIL.n90 VSUBS 2.72459f
C1760 VTAIL.n91 VSUBS 3.31176f
C1761 VTAIL.t7 VSUBS 0.352887f
C1762 VTAIL.t6 VSUBS 0.352887f
C1763 VTAIL.n92 VSUBS 2.72461f
C1764 VTAIL.n93 VSUBS 3.31174f
C1765 VTAIL.t3 VSUBS 0.352887f
C1766 VTAIL.t5 VSUBS 0.352887f
C1767 VTAIL.n94 VSUBS 2.72461f
C1768 VTAIL.n95 VSUBS 1.34207f
C1769 VTAIL.n96 VSUBS 0.031088f
C1770 VTAIL.n97 VSUBS 0.028848f
C1771 VTAIL.n98 VSUBS 0.015502f
C1772 VTAIL.n99 VSUBS 0.03664f
C1773 VTAIL.n100 VSUBS 0.015957f
C1774 VTAIL.n101 VSUBS 0.028848f
C1775 VTAIL.n102 VSUBS 0.015957f
C1776 VTAIL.n103 VSUBS 0.015502f
C1777 VTAIL.n104 VSUBS 0.03664f
C1778 VTAIL.n105 VSUBS 0.03664f
C1779 VTAIL.n106 VSUBS 0.016413f
C1780 VTAIL.n107 VSUBS 0.028848f
C1781 VTAIL.n108 VSUBS 0.015502f
C1782 VTAIL.n109 VSUBS 0.03664f
C1783 VTAIL.n110 VSUBS 0.016413f
C1784 VTAIL.n111 VSUBS 0.028848f
C1785 VTAIL.n112 VSUBS 0.015502f
C1786 VTAIL.n113 VSUBS 0.03664f
C1787 VTAIL.n114 VSUBS 0.016413f
C1788 VTAIL.n115 VSUBS 0.028848f
C1789 VTAIL.n116 VSUBS 0.015502f
C1790 VTAIL.n117 VSUBS 0.03664f
C1791 VTAIL.n118 VSUBS 0.016413f
C1792 VTAIL.n119 VSUBS 0.028848f
C1793 VTAIL.n120 VSUBS 0.015502f
C1794 VTAIL.n121 VSUBS 0.03664f
C1795 VTAIL.n122 VSUBS 0.016413f
C1796 VTAIL.n123 VSUBS 1.90484f
C1797 VTAIL.n124 VSUBS 0.015502f
C1798 VTAIL.t19 VSUBS 0.078473f
C1799 VTAIL.n125 VSUBS 0.207435f
C1800 VTAIL.n126 VSUBS 0.023309f
C1801 VTAIL.n127 VSUBS 0.02748f
C1802 VTAIL.n128 VSUBS 0.03664f
C1803 VTAIL.n129 VSUBS 0.016413f
C1804 VTAIL.n130 VSUBS 0.015502f
C1805 VTAIL.n131 VSUBS 0.028848f
C1806 VTAIL.n132 VSUBS 0.028848f
C1807 VTAIL.n133 VSUBS 0.015502f
C1808 VTAIL.n134 VSUBS 0.016413f
C1809 VTAIL.n135 VSUBS 0.03664f
C1810 VTAIL.n136 VSUBS 0.03664f
C1811 VTAIL.n137 VSUBS 0.016413f
C1812 VTAIL.n138 VSUBS 0.015502f
C1813 VTAIL.n139 VSUBS 0.028848f
C1814 VTAIL.n140 VSUBS 0.028848f
C1815 VTAIL.n141 VSUBS 0.015502f
C1816 VTAIL.n142 VSUBS 0.016413f
C1817 VTAIL.n143 VSUBS 0.03664f
C1818 VTAIL.n144 VSUBS 0.03664f
C1819 VTAIL.n145 VSUBS 0.016413f
C1820 VTAIL.n146 VSUBS 0.015502f
C1821 VTAIL.n147 VSUBS 0.028848f
C1822 VTAIL.n148 VSUBS 0.028848f
C1823 VTAIL.n149 VSUBS 0.015502f
C1824 VTAIL.n150 VSUBS 0.016413f
C1825 VTAIL.n151 VSUBS 0.03664f
C1826 VTAIL.n152 VSUBS 0.03664f
C1827 VTAIL.n153 VSUBS 0.016413f
C1828 VTAIL.n154 VSUBS 0.015502f
C1829 VTAIL.n155 VSUBS 0.028848f
C1830 VTAIL.n156 VSUBS 0.028848f
C1831 VTAIL.n157 VSUBS 0.015502f
C1832 VTAIL.n158 VSUBS 0.016413f
C1833 VTAIL.n159 VSUBS 0.03664f
C1834 VTAIL.n160 VSUBS 0.03664f
C1835 VTAIL.n161 VSUBS 0.016413f
C1836 VTAIL.n162 VSUBS 0.015502f
C1837 VTAIL.n163 VSUBS 0.028848f
C1838 VTAIL.n164 VSUBS 0.028848f
C1839 VTAIL.n165 VSUBS 0.015502f
C1840 VTAIL.n166 VSUBS 0.016413f
C1841 VTAIL.n167 VSUBS 0.03664f
C1842 VTAIL.n168 VSUBS 0.03664f
C1843 VTAIL.n169 VSUBS 0.016413f
C1844 VTAIL.n170 VSUBS 0.015502f
C1845 VTAIL.n171 VSUBS 0.028848f
C1846 VTAIL.n172 VSUBS 0.028848f
C1847 VTAIL.n173 VSUBS 0.015502f
C1848 VTAIL.n174 VSUBS 0.016413f
C1849 VTAIL.n175 VSUBS 0.03664f
C1850 VTAIL.n176 VSUBS 0.086624f
C1851 VTAIL.n177 VSUBS 0.016413f
C1852 VTAIL.n178 VSUBS 0.015502f
C1853 VTAIL.n179 VSUBS 0.071409f
C1854 VTAIL.n180 VSUBS 0.043611f
C1855 VTAIL.n181 VSUBS 0.57702f
C1856 VTAIL.t15 VSUBS 0.352887f
C1857 VTAIL.t11 VSUBS 0.352887f
C1858 VTAIL.n182 VSUBS 2.72461f
C1859 VTAIL.n183 VSUBS 1.21706f
C1860 VTAIL.t14 VSUBS 0.352887f
C1861 VTAIL.t9 VSUBS 0.352887f
C1862 VTAIL.n184 VSUBS 2.72461f
C1863 VTAIL.n185 VSUBS 1.34207f
C1864 VTAIL.n186 VSUBS 0.031088f
C1865 VTAIL.n187 VSUBS 0.028848f
C1866 VTAIL.n188 VSUBS 0.015502f
C1867 VTAIL.n189 VSUBS 0.03664f
C1868 VTAIL.n190 VSUBS 0.015957f
C1869 VTAIL.n191 VSUBS 0.028848f
C1870 VTAIL.n192 VSUBS 0.015957f
C1871 VTAIL.n193 VSUBS 0.015502f
C1872 VTAIL.n194 VSUBS 0.03664f
C1873 VTAIL.n195 VSUBS 0.03664f
C1874 VTAIL.n196 VSUBS 0.016413f
C1875 VTAIL.n197 VSUBS 0.028848f
C1876 VTAIL.n198 VSUBS 0.015502f
C1877 VTAIL.n199 VSUBS 0.03664f
C1878 VTAIL.n200 VSUBS 0.016413f
C1879 VTAIL.n201 VSUBS 0.028848f
C1880 VTAIL.n202 VSUBS 0.015502f
C1881 VTAIL.n203 VSUBS 0.03664f
C1882 VTAIL.n204 VSUBS 0.016413f
C1883 VTAIL.n205 VSUBS 0.028848f
C1884 VTAIL.n206 VSUBS 0.015502f
C1885 VTAIL.n207 VSUBS 0.03664f
C1886 VTAIL.n208 VSUBS 0.016413f
C1887 VTAIL.n209 VSUBS 0.028848f
C1888 VTAIL.n210 VSUBS 0.015502f
C1889 VTAIL.n211 VSUBS 0.03664f
C1890 VTAIL.n212 VSUBS 0.016413f
C1891 VTAIL.n213 VSUBS 1.90484f
C1892 VTAIL.n214 VSUBS 0.015502f
C1893 VTAIL.t12 VSUBS 0.078473f
C1894 VTAIL.n215 VSUBS 0.207435f
C1895 VTAIL.n216 VSUBS 0.023309f
C1896 VTAIL.n217 VSUBS 0.02748f
C1897 VTAIL.n218 VSUBS 0.03664f
C1898 VTAIL.n219 VSUBS 0.016413f
C1899 VTAIL.n220 VSUBS 0.015502f
C1900 VTAIL.n221 VSUBS 0.028848f
C1901 VTAIL.n222 VSUBS 0.028848f
C1902 VTAIL.n223 VSUBS 0.015502f
C1903 VTAIL.n224 VSUBS 0.016413f
C1904 VTAIL.n225 VSUBS 0.03664f
C1905 VTAIL.n226 VSUBS 0.03664f
C1906 VTAIL.n227 VSUBS 0.016413f
C1907 VTAIL.n228 VSUBS 0.015502f
C1908 VTAIL.n229 VSUBS 0.028848f
C1909 VTAIL.n230 VSUBS 0.028848f
C1910 VTAIL.n231 VSUBS 0.015502f
C1911 VTAIL.n232 VSUBS 0.016413f
C1912 VTAIL.n233 VSUBS 0.03664f
C1913 VTAIL.n234 VSUBS 0.03664f
C1914 VTAIL.n235 VSUBS 0.016413f
C1915 VTAIL.n236 VSUBS 0.015502f
C1916 VTAIL.n237 VSUBS 0.028848f
C1917 VTAIL.n238 VSUBS 0.028848f
C1918 VTAIL.n239 VSUBS 0.015502f
C1919 VTAIL.n240 VSUBS 0.016413f
C1920 VTAIL.n241 VSUBS 0.03664f
C1921 VTAIL.n242 VSUBS 0.03664f
C1922 VTAIL.n243 VSUBS 0.016413f
C1923 VTAIL.n244 VSUBS 0.015502f
C1924 VTAIL.n245 VSUBS 0.028848f
C1925 VTAIL.n246 VSUBS 0.028848f
C1926 VTAIL.n247 VSUBS 0.015502f
C1927 VTAIL.n248 VSUBS 0.016413f
C1928 VTAIL.n249 VSUBS 0.03664f
C1929 VTAIL.n250 VSUBS 0.03664f
C1930 VTAIL.n251 VSUBS 0.016413f
C1931 VTAIL.n252 VSUBS 0.015502f
C1932 VTAIL.n253 VSUBS 0.028848f
C1933 VTAIL.n254 VSUBS 0.028848f
C1934 VTAIL.n255 VSUBS 0.015502f
C1935 VTAIL.n256 VSUBS 0.016413f
C1936 VTAIL.n257 VSUBS 0.03664f
C1937 VTAIL.n258 VSUBS 0.03664f
C1938 VTAIL.n259 VSUBS 0.016413f
C1939 VTAIL.n260 VSUBS 0.015502f
C1940 VTAIL.n261 VSUBS 0.028848f
C1941 VTAIL.n262 VSUBS 0.028848f
C1942 VTAIL.n263 VSUBS 0.015502f
C1943 VTAIL.n264 VSUBS 0.016413f
C1944 VTAIL.n265 VSUBS 0.03664f
C1945 VTAIL.n266 VSUBS 0.086624f
C1946 VTAIL.n267 VSUBS 0.016413f
C1947 VTAIL.n268 VSUBS 0.015502f
C1948 VTAIL.n269 VSUBS 0.071409f
C1949 VTAIL.n270 VSUBS 0.043611f
C1950 VTAIL.n271 VSUBS 2.33434f
C1951 VTAIL.n272 VSUBS 0.031088f
C1952 VTAIL.n273 VSUBS 0.028848f
C1953 VTAIL.n274 VSUBS 0.015502f
C1954 VTAIL.n275 VSUBS 0.03664f
C1955 VTAIL.n276 VSUBS 0.015957f
C1956 VTAIL.n277 VSUBS 0.028848f
C1957 VTAIL.n278 VSUBS 0.016413f
C1958 VTAIL.n279 VSUBS 0.03664f
C1959 VTAIL.n280 VSUBS 0.016413f
C1960 VTAIL.n281 VSUBS 0.028848f
C1961 VTAIL.n282 VSUBS 0.015502f
C1962 VTAIL.n283 VSUBS 0.03664f
C1963 VTAIL.n284 VSUBS 0.016413f
C1964 VTAIL.n285 VSUBS 0.028848f
C1965 VTAIL.n286 VSUBS 0.015502f
C1966 VTAIL.n287 VSUBS 0.03664f
C1967 VTAIL.n288 VSUBS 0.016413f
C1968 VTAIL.n289 VSUBS 0.028848f
C1969 VTAIL.n290 VSUBS 0.015502f
C1970 VTAIL.n291 VSUBS 0.03664f
C1971 VTAIL.n292 VSUBS 0.016413f
C1972 VTAIL.n293 VSUBS 0.028848f
C1973 VTAIL.n294 VSUBS 0.015502f
C1974 VTAIL.n295 VSUBS 0.03664f
C1975 VTAIL.n296 VSUBS 0.016413f
C1976 VTAIL.n297 VSUBS 1.90484f
C1977 VTAIL.n298 VSUBS 0.015502f
C1978 VTAIL.t0 VSUBS 0.078473f
C1979 VTAIL.n299 VSUBS 0.207435f
C1980 VTAIL.n300 VSUBS 0.023309f
C1981 VTAIL.n301 VSUBS 0.02748f
C1982 VTAIL.n302 VSUBS 0.03664f
C1983 VTAIL.n303 VSUBS 0.016413f
C1984 VTAIL.n304 VSUBS 0.015502f
C1985 VTAIL.n305 VSUBS 0.028848f
C1986 VTAIL.n306 VSUBS 0.028848f
C1987 VTAIL.n307 VSUBS 0.015502f
C1988 VTAIL.n308 VSUBS 0.016413f
C1989 VTAIL.n309 VSUBS 0.03664f
C1990 VTAIL.n310 VSUBS 0.03664f
C1991 VTAIL.n311 VSUBS 0.016413f
C1992 VTAIL.n312 VSUBS 0.015502f
C1993 VTAIL.n313 VSUBS 0.028848f
C1994 VTAIL.n314 VSUBS 0.028848f
C1995 VTAIL.n315 VSUBS 0.015502f
C1996 VTAIL.n316 VSUBS 0.016413f
C1997 VTAIL.n317 VSUBS 0.03664f
C1998 VTAIL.n318 VSUBS 0.03664f
C1999 VTAIL.n319 VSUBS 0.016413f
C2000 VTAIL.n320 VSUBS 0.015502f
C2001 VTAIL.n321 VSUBS 0.028848f
C2002 VTAIL.n322 VSUBS 0.028848f
C2003 VTAIL.n323 VSUBS 0.015502f
C2004 VTAIL.n324 VSUBS 0.016413f
C2005 VTAIL.n325 VSUBS 0.03664f
C2006 VTAIL.n326 VSUBS 0.03664f
C2007 VTAIL.n327 VSUBS 0.016413f
C2008 VTAIL.n328 VSUBS 0.015502f
C2009 VTAIL.n329 VSUBS 0.028848f
C2010 VTAIL.n330 VSUBS 0.028848f
C2011 VTAIL.n331 VSUBS 0.015502f
C2012 VTAIL.n332 VSUBS 0.016413f
C2013 VTAIL.n333 VSUBS 0.03664f
C2014 VTAIL.n334 VSUBS 0.03664f
C2015 VTAIL.n335 VSUBS 0.016413f
C2016 VTAIL.n336 VSUBS 0.015502f
C2017 VTAIL.n337 VSUBS 0.028848f
C2018 VTAIL.n338 VSUBS 0.028848f
C2019 VTAIL.n339 VSUBS 0.015502f
C2020 VTAIL.n340 VSUBS 0.015502f
C2021 VTAIL.n341 VSUBS 0.016413f
C2022 VTAIL.n342 VSUBS 0.03664f
C2023 VTAIL.n343 VSUBS 0.03664f
C2024 VTAIL.n344 VSUBS 0.03664f
C2025 VTAIL.n345 VSUBS 0.015957f
C2026 VTAIL.n346 VSUBS 0.015502f
C2027 VTAIL.n347 VSUBS 0.028848f
C2028 VTAIL.n348 VSUBS 0.028848f
C2029 VTAIL.n349 VSUBS 0.015502f
C2030 VTAIL.n350 VSUBS 0.016413f
C2031 VTAIL.n351 VSUBS 0.03664f
C2032 VTAIL.n352 VSUBS 0.086624f
C2033 VTAIL.n353 VSUBS 0.016413f
C2034 VTAIL.n354 VSUBS 0.015502f
C2035 VTAIL.n355 VSUBS 0.071409f
C2036 VTAIL.n356 VSUBS 0.043611f
C2037 VTAIL.n357 VSUBS 2.33434f
C2038 VTAIL.t1 VSUBS 0.352887f
C2039 VTAIL.t4 VSUBS 0.352887f
C2040 VTAIL.n358 VSUBS 2.72459f
C2041 VTAIL.n359 VSUBS 1.08366f
C2042 VP.n0 VSUBS 0.042703f
C2043 VP.t1 VSUBS 3.74008f
C2044 VP.n1 VSUBS 0.042111f
C2045 VP.n2 VSUBS 0.022709f
C2046 VP.n3 VSUBS 0.042111f
C2047 VP.n4 VSUBS 0.022709f
C2048 VP.t8 VSUBS 3.74008f
C2049 VP.n5 VSUBS 0.042111f
C2050 VP.n6 VSUBS 0.022709f
C2051 VP.n7 VSUBS 0.042111f
C2052 VP.n8 VSUBS 0.022709f
C2053 VP.t7 VSUBS 3.74008f
C2054 VP.n9 VSUBS 0.042111f
C2055 VP.n10 VSUBS 0.022709f
C2056 VP.n11 VSUBS 0.042111f
C2057 VP.n12 VSUBS 0.022709f
C2058 VP.t3 VSUBS 3.74008f
C2059 VP.n13 VSUBS 0.042111f
C2060 VP.n14 VSUBS 0.022709f
C2061 VP.n15 VSUBS 0.042111f
C2062 VP.n16 VSUBS 0.042703f
C2063 VP.t0 VSUBS 3.74008f
C2064 VP.n17 VSUBS 0.042703f
C2065 VP.t9 VSUBS 3.74008f
C2066 VP.n18 VSUBS 0.042111f
C2067 VP.n19 VSUBS 0.022709f
C2068 VP.n20 VSUBS 0.042111f
C2069 VP.n21 VSUBS 0.022709f
C2070 VP.t2 VSUBS 3.74008f
C2071 VP.n22 VSUBS 0.042111f
C2072 VP.n23 VSUBS 0.022709f
C2073 VP.n24 VSUBS 0.042111f
C2074 VP.n25 VSUBS 0.022709f
C2075 VP.t4 VSUBS 3.74008f
C2076 VP.n26 VSUBS 0.042111f
C2077 VP.n27 VSUBS 0.022709f
C2078 VP.n28 VSUBS 0.042111f
C2079 VP.n29 VSUBS 0.299657f
C2080 VP.t5 VSUBS 3.74008f
C2081 VP.t6 VSUBS 4.11025f
C2082 VP.n30 VSUBS 1.31026f
C2083 VP.n31 VSUBS 1.37481f
C2084 VP.n32 VSUBS 0.030053f
C2085 VP.n33 VSUBS 0.042111f
C2086 VP.n34 VSUBS 0.022709f
C2087 VP.n35 VSUBS 0.022709f
C2088 VP.n36 VSUBS 0.022709f
C2089 VP.n37 VSUBS 0.041254f
C2090 VP.n38 VSUBS 0.021747f
C2091 VP.n39 VSUBS 0.045132f
C2092 VP.n40 VSUBS 0.022709f
C2093 VP.n41 VSUBS 0.022709f
C2094 VP.n42 VSUBS 0.022709f
C2095 VP.n43 VSUBS 0.042111f
C2096 VP.n44 VSUBS 1.31624f
C2097 VP.n45 VSUBS 0.042111f
C2098 VP.n46 VSUBS 0.022709f
C2099 VP.n47 VSUBS 0.022709f
C2100 VP.n48 VSUBS 0.022709f
C2101 VP.n49 VSUBS 0.045132f
C2102 VP.n50 VSUBS 0.021747f
C2103 VP.n51 VSUBS 0.041254f
C2104 VP.n52 VSUBS 0.022709f
C2105 VP.n53 VSUBS 0.022709f
C2106 VP.n54 VSUBS 0.022709f
C2107 VP.n55 VSUBS 0.042111f
C2108 VP.n56 VSUBS 0.030053f
C2109 VP.n57 VSUBS 1.29492f
C2110 VP.n58 VSUBS 0.03338f
C2111 VP.n59 VSUBS 0.022709f
C2112 VP.n60 VSUBS 0.022709f
C2113 VP.n61 VSUBS 0.022709f
C2114 VP.n62 VSUBS 0.042111f
C2115 VP.n63 VSUBS 0.037094f
C2116 VP.n64 VSUBS 0.028927f
C2117 VP.n65 VSUBS 0.022709f
C2118 VP.n66 VSUBS 0.022709f
C2119 VP.n67 VSUBS 0.022709f
C2120 VP.n68 VSUBS 0.042111f
C2121 VP.n69 VSUBS 0.038785f
C2122 VP.n70 VSUBS 1.39258f
C2123 VP.n71 VSUBS 1.79952f
C2124 VP.n72 VSUBS 1.81253f
C2125 VP.n73 VSUBS 1.39258f
C2126 VP.n74 VSUBS 0.038785f
C2127 VP.n75 VSUBS 0.042111f
C2128 VP.n76 VSUBS 0.022709f
C2129 VP.n77 VSUBS 0.022709f
C2130 VP.n78 VSUBS 0.022709f
C2131 VP.n79 VSUBS 0.028927f
C2132 VP.n80 VSUBS 0.037094f
C2133 VP.n81 VSUBS 0.042111f
C2134 VP.n82 VSUBS 0.022709f
C2135 VP.n83 VSUBS 0.022709f
C2136 VP.n84 VSUBS 0.022709f
C2137 VP.n85 VSUBS 0.03338f
C2138 VP.n86 VSUBS 1.29492f
C2139 VP.n87 VSUBS 0.030053f
C2140 VP.n88 VSUBS 0.042111f
C2141 VP.n89 VSUBS 0.022709f
C2142 VP.n90 VSUBS 0.022709f
C2143 VP.n91 VSUBS 0.022709f
C2144 VP.n92 VSUBS 0.041254f
C2145 VP.n93 VSUBS 0.021747f
C2146 VP.n94 VSUBS 0.045132f
C2147 VP.n95 VSUBS 0.022709f
C2148 VP.n96 VSUBS 0.022709f
C2149 VP.n97 VSUBS 0.022709f
C2150 VP.n98 VSUBS 0.042111f
C2151 VP.n99 VSUBS 1.31624f
C2152 VP.n100 VSUBS 0.042111f
C2153 VP.n101 VSUBS 0.022709f
C2154 VP.n102 VSUBS 0.022709f
C2155 VP.n103 VSUBS 0.022709f
C2156 VP.n104 VSUBS 0.045132f
C2157 VP.n105 VSUBS 0.021747f
C2158 VP.n106 VSUBS 0.041254f
C2159 VP.n107 VSUBS 0.022709f
C2160 VP.n108 VSUBS 0.022709f
C2161 VP.n109 VSUBS 0.022709f
C2162 VP.n110 VSUBS 0.042111f
C2163 VP.n111 VSUBS 0.030053f
C2164 VP.n112 VSUBS 1.29492f
C2165 VP.n113 VSUBS 0.03338f
C2166 VP.n114 VSUBS 0.022709f
C2167 VP.n115 VSUBS 0.022709f
C2168 VP.n116 VSUBS 0.022709f
C2169 VP.n117 VSUBS 0.042111f
C2170 VP.n118 VSUBS 0.037094f
C2171 VP.n119 VSUBS 0.028927f
C2172 VP.n120 VSUBS 0.022709f
C2173 VP.n121 VSUBS 0.022709f
C2174 VP.n122 VSUBS 0.022709f
C2175 VP.n123 VSUBS 0.042111f
C2176 VP.n124 VSUBS 0.038785f
C2177 VP.n125 VSUBS 1.39258f
C2178 VP.n126 VSUBS 0.070942f
.ends

