* NGSPICE file created from diff_pair_sample_1273.ext - technology: sky130A

.subckt diff_pair_sample_1273 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t9 VN.t0 VTAIL.t10 B.t0 sky130_fd_pr__nfet_01v8 ad=4.1847 pd=22.24 as=1.77045 ps=11.06 w=10.73 l=1.9
X1 VDD1.t9 VP.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=4.1847 pd=22.24 as=1.77045 ps=11.06 w=10.73 l=1.9
X2 VDD1.t8 VP.t1 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.77045 pd=11.06 as=1.77045 ps=11.06 w=10.73 l=1.9
X3 VDD1.t7 VP.t2 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=1.77045 pd=11.06 as=4.1847 ps=22.24 w=10.73 l=1.9
X4 B.t23 B.t21 B.t22 B.t11 sky130_fd_pr__nfet_01v8 ad=4.1847 pd=22.24 as=0 ps=0 w=10.73 l=1.9
X5 VTAIL.t13 VN.t1 VDD2.t8 B.t2 sky130_fd_pr__nfet_01v8 ad=1.77045 pd=11.06 as=1.77045 ps=11.06 w=10.73 l=1.9
X6 VTAIL.t14 VN.t2 VDD2.t7 B.t9 sky130_fd_pr__nfet_01v8 ad=1.77045 pd=11.06 as=1.77045 ps=11.06 w=10.73 l=1.9
X7 VTAIL.t4 VP.t3 VDD1.t6 B.t4 sky130_fd_pr__nfet_01v8 ad=1.77045 pd=11.06 as=1.77045 ps=11.06 w=10.73 l=1.9
X8 VTAIL.t19 VP.t4 VDD1.t5 B.t9 sky130_fd_pr__nfet_01v8 ad=1.77045 pd=11.06 as=1.77045 ps=11.06 w=10.73 l=1.9
X9 VDD2.t6 VN.t3 VTAIL.t17 B.t1 sky130_fd_pr__nfet_01v8 ad=4.1847 pd=22.24 as=1.77045 ps=11.06 w=10.73 l=1.9
X10 B.t20 B.t18 B.t19 B.t15 sky130_fd_pr__nfet_01v8 ad=4.1847 pd=22.24 as=0 ps=0 w=10.73 l=1.9
X11 VDD2.t5 VN.t4 VTAIL.t16 B.t6 sky130_fd_pr__nfet_01v8 ad=1.77045 pd=11.06 as=4.1847 ps=22.24 w=10.73 l=1.9
X12 VDD2.t4 VN.t5 VTAIL.t12 B.t7 sky130_fd_pr__nfet_01v8 ad=1.77045 pd=11.06 as=4.1847 ps=22.24 w=10.73 l=1.9
X13 VDD2.t3 VN.t6 VTAIL.t18 B.t5 sky130_fd_pr__nfet_01v8 ad=1.77045 pd=11.06 as=1.77045 ps=11.06 w=10.73 l=1.9
X14 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=4.1847 pd=22.24 as=0 ps=0 w=10.73 l=1.9
X15 VDD1.t4 VP.t5 VTAIL.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=1.77045 pd=11.06 as=1.77045 ps=11.06 w=10.73 l=1.9
X16 VTAIL.t3 VP.t6 VDD1.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.77045 pd=11.06 as=1.77045 ps=11.06 w=10.73 l=1.9
X17 VDD1.t2 VP.t7 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=1.77045 pd=11.06 as=4.1847 ps=22.24 w=10.73 l=1.9
X18 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=4.1847 pd=22.24 as=0 ps=0 w=10.73 l=1.9
X19 VTAIL.t9 VN.t7 VDD2.t2 B.t4 sky130_fd_pr__nfet_01v8 ad=1.77045 pd=11.06 as=1.77045 ps=11.06 w=10.73 l=1.9
X20 VDD1.t1 VP.t8 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=4.1847 pd=22.24 as=1.77045 ps=11.06 w=10.73 l=1.9
X21 VDD2.t1 VN.t8 VTAIL.t15 B.t8 sky130_fd_pr__nfet_01v8 ad=1.77045 pd=11.06 as=1.77045 ps=11.06 w=10.73 l=1.9
X22 VTAIL.t2 VP.t9 VDD1.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=1.77045 pd=11.06 as=1.77045 ps=11.06 w=10.73 l=1.9
X23 VTAIL.t11 VN.t9 VDD2.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=1.77045 pd=11.06 as=1.77045 ps=11.06 w=10.73 l=1.9
R0 VN.n7 VN.t0 166.995
R1 VN.n38 VN.t5 166.995
R2 VN.n59 VN.n31 161.3
R3 VN.n58 VN.n57 161.3
R4 VN.n56 VN.n32 161.3
R5 VN.n55 VN.n54 161.3
R6 VN.n52 VN.n33 161.3
R7 VN.n51 VN.n50 161.3
R8 VN.n49 VN.n34 161.3
R9 VN.n48 VN.n47 161.3
R10 VN.n46 VN.n35 161.3
R11 VN.n45 VN.n44 161.3
R12 VN.n43 VN.n36 161.3
R13 VN.n42 VN.n41 161.3
R14 VN.n40 VN.n37 161.3
R15 VN.n28 VN.n0 161.3
R16 VN.n27 VN.n26 161.3
R17 VN.n25 VN.n1 161.3
R18 VN.n24 VN.n23 161.3
R19 VN.n21 VN.n2 161.3
R20 VN.n20 VN.n19 161.3
R21 VN.n18 VN.n3 161.3
R22 VN.n17 VN.n16 161.3
R23 VN.n15 VN.n4 161.3
R24 VN.n14 VN.n13 161.3
R25 VN.n12 VN.n5 161.3
R26 VN.n11 VN.n10 161.3
R27 VN.n9 VN.n6 161.3
R28 VN.n15 VN.t8 136.102
R29 VN.n8 VN.t9 136.102
R30 VN.n22 VN.t7 136.102
R31 VN.n29 VN.t4 136.102
R32 VN.n46 VN.t6 136.102
R33 VN.n39 VN.t2 136.102
R34 VN.n53 VN.t1 136.102
R35 VN.n60 VN.t3 136.102
R36 VN.n30 VN.n29 88.2468
R37 VN.n61 VN.n60 88.2468
R38 VN.n8 VN.n7 58.8387
R39 VN.n39 VN.n38 58.8387
R40 VN.n27 VN.n1 55.548
R41 VN.n58 VN.n32 55.548
R42 VN.n10 VN.n5 51.663
R43 VN.n20 VN.n3 51.663
R44 VN.n41 VN.n36 51.663
R45 VN.n51 VN.n34 51.663
R46 VN VN.n61 48.6686
R47 VN.n14 VN.n5 29.3238
R48 VN.n16 VN.n3 29.3238
R49 VN.n45 VN.n36 29.3238
R50 VN.n47 VN.n34 29.3238
R51 VN.n28 VN.n27 25.4388
R52 VN.n59 VN.n58 25.4388
R53 VN.n10 VN.n9 24.4675
R54 VN.n15 VN.n14 24.4675
R55 VN.n16 VN.n15 24.4675
R56 VN.n21 VN.n20 24.4675
R57 VN.n23 VN.n1 24.4675
R58 VN.n41 VN.n40 24.4675
R59 VN.n47 VN.n46 24.4675
R60 VN.n46 VN.n45 24.4675
R61 VN.n54 VN.n32 24.4675
R62 VN.n52 VN.n51 24.4675
R63 VN.n29 VN.n28 22.5101
R64 VN.n60 VN.n59 22.5101
R65 VN.n23 VN.n22 13.2127
R66 VN.n54 VN.n53 13.2127
R67 VN.n38 VN.n37 12.9374
R68 VN.n7 VN.n6 12.9374
R69 VN.n9 VN.n8 11.2553
R70 VN.n22 VN.n21 11.2553
R71 VN.n40 VN.n39 11.2553
R72 VN.n53 VN.n52 11.2553
R73 VN.n61 VN.n31 0.278367
R74 VN.n30 VN.n0 0.278367
R75 VN.n57 VN.n31 0.189894
R76 VN.n57 VN.n56 0.189894
R77 VN.n56 VN.n55 0.189894
R78 VN.n55 VN.n33 0.189894
R79 VN.n50 VN.n33 0.189894
R80 VN.n50 VN.n49 0.189894
R81 VN.n49 VN.n48 0.189894
R82 VN.n48 VN.n35 0.189894
R83 VN.n44 VN.n35 0.189894
R84 VN.n44 VN.n43 0.189894
R85 VN.n43 VN.n42 0.189894
R86 VN.n42 VN.n37 0.189894
R87 VN.n11 VN.n6 0.189894
R88 VN.n12 VN.n11 0.189894
R89 VN.n13 VN.n12 0.189894
R90 VN.n13 VN.n4 0.189894
R91 VN.n17 VN.n4 0.189894
R92 VN.n18 VN.n17 0.189894
R93 VN.n19 VN.n18 0.189894
R94 VN.n19 VN.n2 0.189894
R95 VN.n24 VN.n2 0.189894
R96 VN.n25 VN.n24 0.189894
R97 VN.n26 VN.n25 0.189894
R98 VN.n26 VN.n0 0.189894
R99 VN VN.n30 0.153454
R100 VTAIL.n240 VTAIL.n188 289.615
R101 VTAIL.n54 VTAIL.n2 289.615
R102 VTAIL.n182 VTAIL.n130 289.615
R103 VTAIL.n120 VTAIL.n68 289.615
R104 VTAIL.n207 VTAIL.n206 185
R105 VTAIL.n204 VTAIL.n203 185
R106 VTAIL.n213 VTAIL.n212 185
R107 VTAIL.n215 VTAIL.n214 185
R108 VTAIL.n200 VTAIL.n199 185
R109 VTAIL.n221 VTAIL.n220 185
R110 VTAIL.n224 VTAIL.n223 185
R111 VTAIL.n222 VTAIL.n196 185
R112 VTAIL.n229 VTAIL.n195 185
R113 VTAIL.n231 VTAIL.n230 185
R114 VTAIL.n233 VTAIL.n232 185
R115 VTAIL.n192 VTAIL.n191 185
R116 VTAIL.n239 VTAIL.n238 185
R117 VTAIL.n241 VTAIL.n240 185
R118 VTAIL.n21 VTAIL.n20 185
R119 VTAIL.n18 VTAIL.n17 185
R120 VTAIL.n27 VTAIL.n26 185
R121 VTAIL.n29 VTAIL.n28 185
R122 VTAIL.n14 VTAIL.n13 185
R123 VTAIL.n35 VTAIL.n34 185
R124 VTAIL.n38 VTAIL.n37 185
R125 VTAIL.n36 VTAIL.n10 185
R126 VTAIL.n43 VTAIL.n9 185
R127 VTAIL.n45 VTAIL.n44 185
R128 VTAIL.n47 VTAIL.n46 185
R129 VTAIL.n6 VTAIL.n5 185
R130 VTAIL.n53 VTAIL.n52 185
R131 VTAIL.n55 VTAIL.n54 185
R132 VTAIL.n183 VTAIL.n182 185
R133 VTAIL.n181 VTAIL.n180 185
R134 VTAIL.n134 VTAIL.n133 185
R135 VTAIL.n175 VTAIL.n174 185
R136 VTAIL.n173 VTAIL.n172 185
R137 VTAIL.n171 VTAIL.n137 185
R138 VTAIL.n141 VTAIL.n138 185
R139 VTAIL.n166 VTAIL.n165 185
R140 VTAIL.n164 VTAIL.n163 185
R141 VTAIL.n143 VTAIL.n142 185
R142 VTAIL.n158 VTAIL.n157 185
R143 VTAIL.n156 VTAIL.n155 185
R144 VTAIL.n147 VTAIL.n146 185
R145 VTAIL.n150 VTAIL.n149 185
R146 VTAIL.n121 VTAIL.n120 185
R147 VTAIL.n119 VTAIL.n118 185
R148 VTAIL.n72 VTAIL.n71 185
R149 VTAIL.n113 VTAIL.n112 185
R150 VTAIL.n111 VTAIL.n110 185
R151 VTAIL.n109 VTAIL.n75 185
R152 VTAIL.n79 VTAIL.n76 185
R153 VTAIL.n104 VTAIL.n103 185
R154 VTAIL.n102 VTAIL.n101 185
R155 VTAIL.n81 VTAIL.n80 185
R156 VTAIL.n96 VTAIL.n95 185
R157 VTAIL.n94 VTAIL.n93 185
R158 VTAIL.n85 VTAIL.n84 185
R159 VTAIL.n88 VTAIL.n87 185
R160 VTAIL.t16 VTAIL.n205 149.524
R161 VTAIL.t7 VTAIL.n19 149.524
R162 VTAIL.t6 VTAIL.n148 149.524
R163 VTAIL.t12 VTAIL.n86 149.524
R164 VTAIL.n206 VTAIL.n203 104.615
R165 VTAIL.n213 VTAIL.n203 104.615
R166 VTAIL.n214 VTAIL.n213 104.615
R167 VTAIL.n214 VTAIL.n199 104.615
R168 VTAIL.n221 VTAIL.n199 104.615
R169 VTAIL.n223 VTAIL.n221 104.615
R170 VTAIL.n223 VTAIL.n222 104.615
R171 VTAIL.n222 VTAIL.n195 104.615
R172 VTAIL.n231 VTAIL.n195 104.615
R173 VTAIL.n232 VTAIL.n231 104.615
R174 VTAIL.n232 VTAIL.n191 104.615
R175 VTAIL.n239 VTAIL.n191 104.615
R176 VTAIL.n240 VTAIL.n239 104.615
R177 VTAIL.n20 VTAIL.n17 104.615
R178 VTAIL.n27 VTAIL.n17 104.615
R179 VTAIL.n28 VTAIL.n27 104.615
R180 VTAIL.n28 VTAIL.n13 104.615
R181 VTAIL.n35 VTAIL.n13 104.615
R182 VTAIL.n37 VTAIL.n35 104.615
R183 VTAIL.n37 VTAIL.n36 104.615
R184 VTAIL.n36 VTAIL.n9 104.615
R185 VTAIL.n45 VTAIL.n9 104.615
R186 VTAIL.n46 VTAIL.n45 104.615
R187 VTAIL.n46 VTAIL.n5 104.615
R188 VTAIL.n53 VTAIL.n5 104.615
R189 VTAIL.n54 VTAIL.n53 104.615
R190 VTAIL.n182 VTAIL.n181 104.615
R191 VTAIL.n181 VTAIL.n133 104.615
R192 VTAIL.n174 VTAIL.n133 104.615
R193 VTAIL.n174 VTAIL.n173 104.615
R194 VTAIL.n173 VTAIL.n137 104.615
R195 VTAIL.n141 VTAIL.n137 104.615
R196 VTAIL.n165 VTAIL.n141 104.615
R197 VTAIL.n165 VTAIL.n164 104.615
R198 VTAIL.n164 VTAIL.n142 104.615
R199 VTAIL.n157 VTAIL.n142 104.615
R200 VTAIL.n157 VTAIL.n156 104.615
R201 VTAIL.n156 VTAIL.n146 104.615
R202 VTAIL.n149 VTAIL.n146 104.615
R203 VTAIL.n120 VTAIL.n119 104.615
R204 VTAIL.n119 VTAIL.n71 104.615
R205 VTAIL.n112 VTAIL.n71 104.615
R206 VTAIL.n112 VTAIL.n111 104.615
R207 VTAIL.n111 VTAIL.n75 104.615
R208 VTAIL.n79 VTAIL.n75 104.615
R209 VTAIL.n103 VTAIL.n79 104.615
R210 VTAIL.n103 VTAIL.n102 104.615
R211 VTAIL.n102 VTAIL.n80 104.615
R212 VTAIL.n95 VTAIL.n80 104.615
R213 VTAIL.n95 VTAIL.n94 104.615
R214 VTAIL.n94 VTAIL.n84 104.615
R215 VTAIL.n87 VTAIL.n84 104.615
R216 VTAIL.n206 VTAIL.t16 52.3082
R217 VTAIL.n20 VTAIL.t7 52.3082
R218 VTAIL.n149 VTAIL.t6 52.3082
R219 VTAIL.n87 VTAIL.t12 52.3082
R220 VTAIL.n129 VTAIL.n128 46.6312
R221 VTAIL.n127 VTAIL.n126 46.6312
R222 VTAIL.n67 VTAIL.n66 46.6312
R223 VTAIL.n65 VTAIL.n64 46.6312
R224 VTAIL.n247 VTAIL.n246 46.631
R225 VTAIL.n1 VTAIL.n0 46.631
R226 VTAIL.n61 VTAIL.n60 46.631
R227 VTAIL.n63 VTAIL.n62 46.631
R228 VTAIL.n245 VTAIL.n244 33.155
R229 VTAIL.n59 VTAIL.n58 33.155
R230 VTAIL.n187 VTAIL.n186 33.155
R231 VTAIL.n125 VTAIL.n124 33.155
R232 VTAIL.n65 VTAIL.n63 25.4617
R233 VTAIL.n245 VTAIL.n187 23.5393
R234 VTAIL.n230 VTAIL.n229 13.1884
R235 VTAIL.n44 VTAIL.n43 13.1884
R236 VTAIL.n172 VTAIL.n171 13.1884
R237 VTAIL.n110 VTAIL.n109 13.1884
R238 VTAIL.n228 VTAIL.n196 12.8005
R239 VTAIL.n233 VTAIL.n194 12.8005
R240 VTAIL.n42 VTAIL.n10 12.8005
R241 VTAIL.n47 VTAIL.n8 12.8005
R242 VTAIL.n175 VTAIL.n136 12.8005
R243 VTAIL.n170 VTAIL.n138 12.8005
R244 VTAIL.n113 VTAIL.n74 12.8005
R245 VTAIL.n108 VTAIL.n76 12.8005
R246 VTAIL.n225 VTAIL.n224 12.0247
R247 VTAIL.n234 VTAIL.n192 12.0247
R248 VTAIL.n39 VTAIL.n38 12.0247
R249 VTAIL.n48 VTAIL.n6 12.0247
R250 VTAIL.n176 VTAIL.n134 12.0247
R251 VTAIL.n167 VTAIL.n166 12.0247
R252 VTAIL.n114 VTAIL.n72 12.0247
R253 VTAIL.n105 VTAIL.n104 12.0247
R254 VTAIL.n220 VTAIL.n198 11.249
R255 VTAIL.n238 VTAIL.n237 11.249
R256 VTAIL.n34 VTAIL.n12 11.249
R257 VTAIL.n52 VTAIL.n51 11.249
R258 VTAIL.n180 VTAIL.n179 11.249
R259 VTAIL.n163 VTAIL.n140 11.249
R260 VTAIL.n118 VTAIL.n117 11.249
R261 VTAIL.n101 VTAIL.n78 11.249
R262 VTAIL.n219 VTAIL.n200 10.4732
R263 VTAIL.n241 VTAIL.n190 10.4732
R264 VTAIL.n33 VTAIL.n14 10.4732
R265 VTAIL.n55 VTAIL.n4 10.4732
R266 VTAIL.n183 VTAIL.n132 10.4732
R267 VTAIL.n162 VTAIL.n143 10.4732
R268 VTAIL.n121 VTAIL.n70 10.4732
R269 VTAIL.n100 VTAIL.n81 10.4732
R270 VTAIL.n207 VTAIL.n205 10.2747
R271 VTAIL.n21 VTAIL.n19 10.2747
R272 VTAIL.n150 VTAIL.n148 10.2747
R273 VTAIL.n88 VTAIL.n86 10.2747
R274 VTAIL.n216 VTAIL.n215 9.69747
R275 VTAIL.n242 VTAIL.n188 9.69747
R276 VTAIL.n30 VTAIL.n29 9.69747
R277 VTAIL.n56 VTAIL.n2 9.69747
R278 VTAIL.n184 VTAIL.n130 9.69747
R279 VTAIL.n159 VTAIL.n158 9.69747
R280 VTAIL.n122 VTAIL.n68 9.69747
R281 VTAIL.n97 VTAIL.n96 9.69747
R282 VTAIL.n244 VTAIL.n243 9.45567
R283 VTAIL.n58 VTAIL.n57 9.45567
R284 VTAIL.n186 VTAIL.n185 9.45567
R285 VTAIL.n124 VTAIL.n123 9.45567
R286 VTAIL.n243 VTAIL.n242 9.3005
R287 VTAIL.n190 VTAIL.n189 9.3005
R288 VTAIL.n237 VTAIL.n236 9.3005
R289 VTAIL.n235 VTAIL.n234 9.3005
R290 VTAIL.n194 VTAIL.n193 9.3005
R291 VTAIL.n209 VTAIL.n208 9.3005
R292 VTAIL.n211 VTAIL.n210 9.3005
R293 VTAIL.n202 VTAIL.n201 9.3005
R294 VTAIL.n217 VTAIL.n216 9.3005
R295 VTAIL.n219 VTAIL.n218 9.3005
R296 VTAIL.n198 VTAIL.n197 9.3005
R297 VTAIL.n226 VTAIL.n225 9.3005
R298 VTAIL.n228 VTAIL.n227 9.3005
R299 VTAIL.n57 VTAIL.n56 9.3005
R300 VTAIL.n4 VTAIL.n3 9.3005
R301 VTAIL.n51 VTAIL.n50 9.3005
R302 VTAIL.n49 VTAIL.n48 9.3005
R303 VTAIL.n8 VTAIL.n7 9.3005
R304 VTAIL.n23 VTAIL.n22 9.3005
R305 VTAIL.n25 VTAIL.n24 9.3005
R306 VTAIL.n16 VTAIL.n15 9.3005
R307 VTAIL.n31 VTAIL.n30 9.3005
R308 VTAIL.n33 VTAIL.n32 9.3005
R309 VTAIL.n12 VTAIL.n11 9.3005
R310 VTAIL.n40 VTAIL.n39 9.3005
R311 VTAIL.n42 VTAIL.n41 9.3005
R312 VTAIL.n152 VTAIL.n151 9.3005
R313 VTAIL.n154 VTAIL.n153 9.3005
R314 VTAIL.n145 VTAIL.n144 9.3005
R315 VTAIL.n160 VTAIL.n159 9.3005
R316 VTAIL.n162 VTAIL.n161 9.3005
R317 VTAIL.n140 VTAIL.n139 9.3005
R318 VTAIL.n168 VTAIL.n167 9.3005
R319 VTAIL.n170 VTAIL.n169 9.3005
R320 VTAIL.n185 VTAIL.n184 9.3005
R321 VTAIL.n132 VTAIL.n131 9.3005
R322 VTAIL.n179 VTAIL.n178 9.3005
R323 VTAIL.n177 VTAIL.n176 9.3005
R324 VTAIL.n136 VTAIL.n135 9.3005
R325 VTAIL.n90 VTAIL.n89 9.3005
R326 VTAIL.n92 VTAIL.n91 9.3005
R327 VTAIL.n83 VTAIL.n82 9.3005
R328 VTAIL.n98 VTAIL.n97 9.3005
R329 VTAIL.n100 VTAIL.n99 9.3005
R330 VTAIL.n78 VTAIL.n77 9.3005
R331 VTAIL.n106 VTAIL.n105 9.3005
R332 VTAIL.n108 VTAIL.n107 9.3005
R333 VTAIL.n123 VTAIL.n122 9.3005
R334 VTAIL.n70 VTAIL.n69 9.3005
R335 VTAIL.n117 VTAIL.n116 9.3005
R336 VTAIL.n115 VTAIL.n114 9.3005
R337 VTAIL.n74 VTAIL.n73 9.3005
R338 VTAIL.n212 VTAIL.n202 8.92171
R339 VTAIL.n26 VTAIL.n16 8.92171
R340 VTAIL.n155 VTAIL.n145 8.92171
R341 VTAIL.n93 VTAIL.n83 8.92171
R342 VTAIL.n211 VTAIL.n204 8.14595
R343 VTAIL.n25 VTAIL.n18 8.14595
R344 VTAIL.n154 VTAIL.n147 8.14595
R345 VTAIL.n92 VTAIL.n85 8.14595
R346 VTAIL.n208 VTAIL.n207 7.3702
R347 VTAIL.n22 VTAIL.n21 7.3702
R348 VTAIL.n151 VTAIL.n150 7.3702
R349 VTAIL.n89 VTAIL.n88 7.3702
R350 VTAIL.n208 VTAIL.n204 5.81868
R351 VTAIL.n22 VTAIL.n18 5.81868
R352 VTAIL.n151 VTAIL.n147 5.81868
R353 VTAIL.n89 VTAIL.n85 5.81868
R354 VTAIL.n212 VTAIL.n211 5.04292
R355 VTAIL.n26 VTAIL.n25 5.04292
R356 VTAIL.n155 VTAIL.n154 5.04292
R357 VTAIL.n93 VTAIL.n92 5.04292
R358 VTAIL.n215 VTAIL.n202 4.26717
R359 VTAIL.n244 VTAIL.n188 4.26717
R360 VTAIL.n29 VTAIL.n16 4.26717
R361 VTAIL.n58 VTAIL.n2 4.26717
R362 VTAIL.n186 VTAIL.n130 4.26717
R363 VTAIL.n158 VTAIL.n145 4.26717
R364 VTAIL.n124 VTAIL.n68 4.26717
R365 VTAIL.n96 VTAIL.n83 4.26717
R366 VTAIL.n216 VTAIL.n200 3.49141
R367 VTAIL.n242 VTAIL.n241 3.49141
R368 VTAIL.n30 VTAIL.n14 3.49141
R369 VTAIL.n56 VTAIL.n55 3.49141
R370 VTAIL.n184 VTAIL.n183 3.49141
R371 VTAIL.n159 VTAIL.n143 3.49141
R372 VTAIL.n122 VTAIL.n121 3.49141
R373 VTAIL.n97 VTAIL.n81 3.49141
R374 VTAIL.n209 VTAIL.n205 2.84303
R375 VTAIL.n23 VTAIL.n19 2.84303
R376 VTAIL.n152 VTAIL.n148 2.84303
R377 VTAIL.n90 VTAIL.n86 2.84303
R378 VTAIL.n220 VTAIL.n219 2.71565
R379 VTAIL.n238 VTAIL.n190 2.71565
R380 VTAIL.n34 VTAIL.n33 2.71565
R381 VTAIL.n52 VTAIL.n4 2.71565
R382 VTAIL.n180 VTAIL.n132 2.71565
R383 VTAIL.n163 VTAIL.n162 2.71565
R384 VTAIL.n118 VTAIL.n70 2.71565
R385 VTAIL.n101 VTAIL.n100 2.71565
R386 VTAIL.n224 VTAIL.n198 1.93989
R387 VTAIL.n237 VTAIL.n192 1.93989
R388 VTAIL.n38 VTAIL.n12 1.93989
R389 VTAIL.n51 VTAIL.n6 1.93989
R390 VTAIL.n179 VTAIL.n134 1.93989
R391 VTAIL.n166 VTAIL.n140 1.93989
R392 VTAIL.n117 VTAIL.n72 1.93989
R393 VTAIL.n104 VTAIL.n78 1.93989
R394 VTAIL.n67 VTAIL.n65 1.92291
R395 VTAIL.n125 VTAIL.n67 1.92291
R396 VTAIL.n129 VTAIL.n127 1.92291
R397 VTAIL.n187 VTAIL.n129 1.92291
R398 VTAIL.n63 VTAIL.n61 1.92291
R399 VTAIL.n61 VTAIL.n59 1.92291
R400 VTAIL.n247 VTAIL.n245 1.92291
R401 VTAIL.n246 VTAIL.t15 1.84579
R402 VTAIL.n246 VTAIL.t9 1.84579
R403 VTAIL.n0 VTAIL.t10 1.84579
R404 VTAIL.n0 VTAIL.t11 1.84579
R405 VTAIL.n60 VTAIL.t5 1.84579
R406 VTAIL.n60 VTAIL.t19 1.84579
R407 VTAIL.n62 VTAIL.t1 1.84579
R408 VTAIL.n62 VTAIL.t2 1.84579
R409 VTAIL.n128 VTAIL.t8 1.84579
R410 VTAIL.n128 VTAIL.t4 1.84579
R411 VTAIL.n126 VTAIL.t0 1.84579
R412 VTAIL.n126 VTAIL.t3 1.84579
R413 VTAIL.n66 VTAIL.t18 1.84579
R414 VTAIL.n66 VTAIL.t14 1.84579
R415 VTAIL.n64 VTAIL.t17 1.84579
R416 VTAIL.n64 VTAIL.t13 1.84579
R417 VTAIL VTAIL.n1 1.5005
R418 VTAIL.n127 VTAIL.n125 1.43153
R419 VTAIL.n59 VTAIL.n1 1.43153
R420 VTAIL.n225 VTAIL.n196 1.16414
R421 VTAIL.n234 VTAIL.n233 1.16414
R422 VTAIL.n39 VTAIL.n10 1.16414
R423 VTAIL.n48 VTAIL.n47 1.16414
R424 VTAIL.n176 VTAIL.n175 1.16414
R425 VTAIL.n167 VTAIL.n138 1.16414
R426 VTAIL.n114 VTAIL.n113 1.16414
R427 VTAIL.n105 VTAIL.n76 1.16414
R428 VTAIL VTAIL.n247 0.422914
R429 VTAIL.n229 VTAIL.n228 0.388379
R430 VTAIL.n230 VTAIL.n194 0.388379
R431 VTAIL.n43 VTAIL.n42 0.388379
R432 VTAIL.n44 VTAIL.n8 0.388379
R433 VTAIL.n172 VTAIL.n136 0.388379
R434 VTAIL.n171 VTAIL.n170 0.388379
R435 VTAIL.n110 VTAIL.n74 0.388379
R436 VTAIL.n109 VTAIL.n108 0.388379
R437 VTAIL.n210 VTAIL.n209 0.155672
R438 VTAIL.n210 VTAIL.n201 0.155672
R439 VTAIL.n217 VTAIL.n201 0.155672
R440 VTAIL.n218 VTAIL.n217 0.155672
R441 VTAIL.n218 VTAIL.n197 0.155672
R442 VTAIL.n226 VTAIL.n197 0.155672
R443 VTAIL.n227 VTAIL.n226 0.155672
R444 VTAIL.n227 VTAIL.n193 0.155672
R445 VTAIL.n235 VTAIL.n193 0.155672
R446 VTAIL.n236 VTAIL.n235 0.155672
R447 VTAIL.n236 VTAIL.n189 0.155672
R448 VTAIL.n243 VTAIL.n189 0.155672
R449 VTAIL.n24 VTAIL.n23 0.155672
R450 VTAIL.n24 VTAIL.n15 0.155672
R451 VTAIL.n31 VTAIL.n15 0.155672
R452 VTAIL.n32 VTAIL.n31 0.155672
R453 VTAIL.n32 VTAIL.n11 0.155672
R454 VTAIL.n40 VTAIL.n11 0.155672
R455 VTAIL.n41 VTAIL.n40 0.155672
R456 VTAIL.n41 VTAIL.n7 0.155672
R457 VTAIL.n49 VTAIL.n7 0.155672
R458 VTAIL.n50 VTAIL.n49 0.155672
R459 VTAIL.n50 VTAIL.n3 0.155672
R460 VTAIL.n57 VTAIL.n3 0.155672
R461 VTAIL.n185 VTAIL.n131 0.155672
R462 VTAIL.n178 VTAIL.n131 0.155672
R463 VTAIL.n178 VTAIL.n177 0.155672
R464 VTAIL.n177 VTAIL.n135 0.155672
R465 VTAIL.n169 VTAIL.n135 0.155672
R466 VTAIL.n169 VTAIL.n168 0.155672
R467 VTAIL.n168 VTAIL.n139 0.155672
R468 VTAIL.n161 VTAIL.n139 0.155672
R469 VTAIL.n161 VTAIL.n160 0.155672
R470 VTAIL.n160 VTAIL.n144 0.155672
R471 VTAIL.n153 VTAIL.n144 0.155672
R472 VTAIL.n153 VTAIL.n152 0.155672
R473 VTAIL.n123 VTAIL.n69 0.155672
R474 VTAIL.n116 VTAIL.n69 0.155672
R475 VTAIL.n116 VTAIL.n115 0.155672
R476 VTAIL.n115 VTAIL.n73 0.155672
R477 VTAIL.n107 VTAIL.n73 0.155672
R478 VTAIL.n107 VTAIL.n106 0.155672
R479 VTAIL.n106 VTAIL.n77 0.155672
R480 VTAIL.n99 VTAIL.n77 0.155672
R481 VTAIL.n99 VTAIL.n98 0.155672
R482 VTAIL.n98 VTAIL.n82 0.155672
R483 VTAIL.n91 VTAIL.n82 0.155672
R484 VTAIL.n91 VTAIL.n90 0.155672
R485 VDD2.n113 VDD2.n61 289.615
R486 VDD2.n52 VDD2.n0 289.615
R487 VDD2.n114 VDD2.n113 185
R488 VDD2.n112 VDD2.n111 185
R489 VDD2.n65 VDD2.n64 185
R490 VDD2.n106 VDD2.n105 185
R491 VDD2.n104 VDD2.n103 185
R492 VDD2.n102 VDD2.n68 185
R493 VDD2.n72 VDD2.n69 185
R494 VDD2.n97 VDD2.n96 185
R495 VDD2.n95 VDD2.n94 185
R496 VDD2.n74 VDD2.n73 185
R497 VDD2.n89 VDD2.n88 185
R498 VDD2.n87 VDD2.n86 185
R499 VDD2.n78 VDD2.n77 185
R500 VDD2.n81 VDD2.n80 185
R501 VDD2.n19 VDD2.n18 185
R502 VDD2.n16 VDD2.n15 185
R503 VDD2.n25 VDD2.n24 185
R504 VDD2.n27 VDD2.n26 185
R505 VDD2.n12 VDD2.n11 185
R506 VDD2.n33 VDD2.n32 185
R507 VDD2.n36 VDD2.n35 185
R508 VDD2.n34 VDD2.n8 185
R509 VDD2.n41 VDD2.n7 185
R510 VDD2.n43 VDD2.n42 185
R511 VDD2.n45 VDD2.n44 185
R512 VDD2.n4 VDD2.n3 185
R513 VDD2.n51 VDD2.n50 185
R514 VDD2.n53 VDD2.n52 185
R515 VDD2.t6 VDD2.n79 149.524
R516 VDD2.t9 VDD2.n17 149.524
R517 VDD2.n113 VDD2.n112 104.615
R518 VDD2.n112 VDD2.n64 104.615
R519 VDD2.n105 VDD2.n64 104.615
R520 VDD2.n105 VDD2.n104 104.615
R521 VDD2.n104 VDD2.n68 104.615
R522 VDD2.n72 VDD2.n68 104.615
R523 VDD2.n96 VDD2.n72 104.615
R524 VDD2.n96 VDD2.n95 104.615
R525 VDD2.n95 VDD2.n73 104.615
R526 VDD2.n88 VDD2.n73 104.615
R527 VDD2.n88 VDD2.n87 104.615
R528 VDD2.n87 VDD2.n77 104.615
R529 VDD2.n80 VDD2.n77 104.615
R530 VDD2.n18 VDD2.n15 104.615
R531 VDD2.n25 VDD2.n15 104.615
R532 VDD2.n26 VDD2.n25 104.615
R533 VDD2.n26 VDD2.n11 104.615
R534 VDD2.n33 VDD2.n11 104.615
R535 VDD2.n35 VDD2.n33 104.615
R536 VDD2.n35 VDD2.n34 104.615
R537 VDD2.n34 VDD2.n7 104.615
R538 VDD2.n43 VDD2.n7 104.615
R539 VDD2.n44 VDD2.n43 104.615
R540 VDD2.n44 VDD2.n3 104.615
R541 VDD2.n51 VDD2.n3 104.615
R542 VDD2.n52 VDD2.n51 104.615
R543 VDD2.n60 VDD2.n59 64.6963
R544 VDD2 VDD2.n121 64.6934
R545 VDD2.n120 VDD2.n119 63.31
R546 VDD2.n58 VDD2.n57 63.3098
R547 VDD2.n80 VDD2.t6 52.3082
R548 VDD2.n18 VDD2.t9 52.3082
R549 VDD2.n58 VDD2.n56 51.7562
R550 VDD2.n118 VDD2.n117 49.8338
R551 VDD2.n118 VDD2.n60 42.0968
R552 VDD2.n103 VDD2.n102 13.1884
R553 VDD2.n42 VDD2.n41 13.1884
R554 VDD2.n106 VDD2.n67 12.8005
R555 VDD2.n101 VDD2.n69 12.8005
R556 VDD2.n40 VDD2.n8 12.8005
R557 VDD2.n45 VDD2.n6 12.8005
R558 VDD2.n107 VDD2.n65 12.0247
R559 VDD2.n98 VDD2.n97 12.0247
R560 VDD2.n37 VDD2.n36 12.0247
R561 VDD2.n46 VDD2.n4 12.0247
R562 VDD2.n111 VDD2.n110 11.249
R563 VDD2.n94 VDD2.n71 11.249
R564 VDD2.n32 VDD2.n10 11.249
R565 VDD2.n50 VDD2.n49 11.249
R566 VDD2.n114 VDD2.n63 10.4732
R567 VDD2.n93 VDD2.n74 10.4732
R568 VDD2.n31 VDD2.n12 10.4732
R569 VDD2.n53 VDD2.n2 10.4732
R570 VDD2.n81 VDD2.n79 10.2747
R571 VDD2.n19 VDD2.n17 10.2747
R572 VDD2.n115 VDD2.n61 9.69747
R573 VDD2.n90 VDD2.n89 9.69747
R574 VDD2.n28 VDD2.n27 9.69747
R575 VDD2.n54 VDD2.n0 9.69747
R576 VDD2.n117 VDD2.n116 9.45567
R577 VDD2.n56 VDD2.n55 9.45567
R578 VDD2.n83 VDD2.n82 9.3005
R579 VDD2.n85 VDD2.n84 9.3005
R580 VDD2.n76 VDD2.n75 9.3005
R581 VDD2.n91 VDD2.n90 9.3005
R582 VDD2.n93 VDD2.n92 9.3005
R583 VDD2.n71 VDD2.n70 9.3005
R584 VDD2.n99 VDD2.n98 9.3005
R585 VDD2.n101 VDD2.n100 9.3005
R586 VDD2.n116 VDD2.n115 9.3005
R587 VDD2.n63 VDD2.n62 9.3005
R588 VDD2.n110 VDD2.n109 9.3005
R589 VDD2.n108 VDD2.n107 9.3005
R590 VDD2.n67 VDD2.n66 9.3005
R591 VDD2.n55 VDD2.n54 9.3005
R592 VDD2.n2 VDD2.n1 9.3005
R593 VDD2.n49 VDD2.n48 9.3005
R594 VDD2.n47 VDD2.n46 9.3005
R595 VDD2.n6 VDD2.n5 9.3005
R596 VDD2.n21 VDD2.n20 9.3005
R597 VDD2.n23 VDD2.n22 9.3005
R598 VDD2.n14 VDD2.n13 9.3005
R599 VDD2.n29 VDD2.n28 9.3005
R600 VDD2.n31 VDD2.n30 9.3005
R601 VDD2.n10 VDD2.n9 9.3005
R602 VDD2.n38 VDD2.n37 9.3005
R603 VDD2.n40 VDD2.n39 9.3005
R604 VDD2.n86 VDD2.n76 8.92171
R605 VDD2.n24 VDD2.n14 8.92171
R606 VDD2.n85 VDD2.n78 8.14595
R607 VDD2.n23 VDD2.n16 8.14595
R608 VDD2.n82 VDD2.n81 7.3702
R609 VDD2.n20 VDD2.n19 7.3702
R610 VDD2.n82 VDD2.n78 5.81868
R611 VDD2.n20 VDD2.n16 5.81868
R612 VDD2.n86 VDD2.n85 5.04292
R613 VDD2.n24 VDD2.n23 5.04292
R614 VDD2.n117 VDD2.n61 4.26717
R615 VDD2.n89 VDD2.n76 4.26717
R616 VDD2.n27 VDD2.n14 4.26717
R617 VDD2.n56 VDD2.n0 4.26717
R618 VDD2.n115 VDD2.n114 3.49141
R619 VDD2.n90 VDD2.n74 3.49141
R620 VDD2.n28 VDD2.n12 3.49141
R621 VDD2.n54 VDD2.n53 3.49141
R622 VDD2.n83 VDD2.n79 2.84303
R623 VDD2.n21 VDD2.n17 2.84303
R624 VDD2.n111 VDD2.n63 2.71565
R625 VDD2.n94 VDD2.n93 2.71565
R626 VDD2.n32 VDD2.n31 2.71565
R627 VDD2.n50 VDD2.n2 2.71565
R628 VDD2.n110 VDD2.n65 1.93989
R629 VDD2.n97 VDD2.n71 1.93989
R630 VDD2.n36 VDD2.n10 1.93989
R631 VDD2.n49 VDD2.n4 1.93989
R632 VDD2.n120 VDD2.n118 1.92291
R633 VDD2.n121 VDD2.t7 1.84579
R634 VDD2.n121 VDD2.t4 1.84579
R635 VDD2.n119 VDD2.t8 1.84579
R636 VDD2.n119 VDD2.t3 1.84579
R637 VDD2.n59 VDD2.t2 1.84579
R638 VDD2.n59 VDD2.t5 1.84579
R639 VDD2.n57 VDD2.t0 1.84579
R640 VDD2.n57 VDD2.t1 1.84579
R641 VDD2.n107 VDD2.n106 1.16414
R642 VDD2.n98 VDD2.n69 1.16414
R643 VDD2.n37 VDD2.n8 1.16414
R644 VDD2.n46 VDD2.n45 1.16414
R645 VDD2 VDD2.n120 0.539293
R646 VDD2.n60 VDD2.n58 0.425757
R647 VDD2.n103 VDD2.n67 0.388379
R648 VDD2.n102 VDD2.n101 0.388379
R649 VDD2.n41 VDD2.n40 0.388379
R650 VDD2.n42 VDD2.n6 0.388379
R651 VDD2.n116 VDD2.n62 0.155672
R652 VDD2.n109 VDD2.n62 0.155672
R653 VDD2.n109 VDD2.n108 0.155672
R654 VDD2.n108 VDD2.n66 0.155672
R655 VDD2.n100 VDD2.n66 0.155672
R656 VDD2.n100 VDD2.n99 0.155672
R657 VDD2.n99 VDD2.n70 0.155672
R658 VDD2.n92 VDD2.n70 0.155672
R659 VDD2.n92 VDD2.n91 0.155672
R660 VDD2.n91 VDD2.n75 0.155672
R661 VDD2.n84 VDD2.n75 0.155672
R662 VDD2.n84 VDD2.n83 0.155672
R663 VDD2.n22 VDD2.n21 0.155672
R664 VDD2.n22 VDD2.n13 0.155672
R665 VDD2.n29 VDD2.n13 0.155672
R666 VDD2.n30 VDD2.n29 0.155672
R667 VDD2.n30 VDD2.n9 0.155672
R668 VDD2.n38 VDD2.n9 0.155672
R669 VDD2.n39 VDD2.n38 0.155672
R670 VDD2.n39 VDD2.n5 0.155672
R671 VDD2.n47 VDD2.n5 0.155672
R672 VDD2.n48 VDD2.n47 0.155672
R673 VDD2.n48 VDD2.n1 0.155672
R674 VDD2.n55 VDD2.n1 0.155672
R675 B.n815 B.n814 585
R676 B.n816 B.n815 585
R677 B.n301 B.n131 585
R678 B.n300 B.n299 585
R679 B.n298 B.n297 585
R680 B.n296 B.n295 585
R681 B.n294 B.n293 585
R682 B.n292 B.n291 585
R683 B.n290 B.n289 585
R684 B.n288 B.n287 585
R685 B.n286 B.n285 585
R686 B.n284 B.n283 585
R687 B.n282 B.n281 585
R688 B.n280 B.n279 585
R689 B.n278 B.n277 585
R690 B.n276 B.n275 585
R691 B.n274 B.n273 585
R692 B.n272 B.n271 585
R693 B.n270 B.n269 585
R694 B.n268 B.n267 585
R695 B.n266 B.n265 585
R696 B.n264 B.n263 585
R697 B.n262 B.n261 585
R698 B.n260 B.n259 585
R699 B.n258 B.n257 585
R700 B.n256 B.n255 585
R701 B.n254 B.n253 585
R702 B.n252 B.n251 585
R703 B.n250 B.n249 585
R704 B.n248 B.n247 585
R705 B.n246 B.n245 585
R706 B.n244 B.n243 585
R707 B.n242 B.n241 585
R708 B.n240 B.n239 585
R709 B.n238 B.n237 585
R710 B.n236 B.n235 585
R711 B.n234 B.n233 585
R712 B.n232 B.n231 585
R713 B.n230 B.n229 585
R714 B.n227 B.n226 585
R715 B.n225 B.n224 585
R716 B.n223 B.n222 585
R717 B.n221 B.n220 585
R718 B.n219 B.n218 585
R719 B.n217 B.n216 585
R720 B.n215 B.n214 585
R721 B.n213 B.n212 585
R722 B.n211 B.n210 585
R723 B.n209 B.n208 585
R724 B.n207 B.n206 585
R725 B.n205 B.n204 585
R726 B.n203 B.n202 585
R727 B.n201 B.n200 585
R728 B.n199 B.n198 585
R729 B.n197 B.n196 585
R730 B.n195 B.n194 585
R731 B.n193 B.n192 585
R732 B.n191 B.n190 585
R733 B.n189 B.n188 585
R734 B.n187 B.n186 585
R735 B.n185 B.n184 585
R736 B.n183 B.n182 585
R737 B.n181 B.n180 585
R738 B.n179 B.n178 585
R739 B.n177 B.n176 585
R740 B.n175 B.n174 585
R741 B.n173 B.n172 585
R742 B.n171 B.n170 585
R743 B.n169 B.n168 585
R744 B.n167 B.n166 585
R745 B.n165 B.n164 585
R746 B.n163 B.n162 585
R747 B.n161 B.n160 585
R748 B.n159 B.n158 585
R749 B.n157 B.n156 585
R750 B.n155 B.n154 585
R751 B.n153 B.n152 585
R752 B.n151 B.n150 585
R753 B.n149 B.n148 585
R754 B.n147 B.n146 585
R755 B.n145 B.n144 585
R756 B.n143 B.n142 585
R757 B.n141 B.n140 585
R758 B.n139 B.n138 585
R759 B.n89 B.n88 585
R760 B.n819 B.n818 585
R761 B.n813 B.n132 585
R762 B.n132 B.n86 585
R763 B.n812 B.n85 585
R764 B.n823 B.n85 585
R765 B.n811 B.n84 585
R766 B.n824 B.n84 585
R767 B.n810 B.n83 585
R768 B.n825 B.n83 585
R769 B.n809 B.n808 585
R770 B.n808 B.n79 585
R771 B.n807 B.n78 585
R772 B.n831 B.n78 585
R773 B.n806 B.n77 585
R774 B.n832 B.n77 585
R775 B.n805 B.n76 585
R776 B.n833 B.n76 585
R777 B.n804 B.n803 585
R778 B.n803 B.n72 585
R779 B.n802 B.n71 585
R780 B.n839 B.n71 585
R781 B.n801 B.n70 585
R782 B.n840 B.n70 585
R783 B.n800 B.n69 585
R784 B.n841 B.n69 585
R785 B.n799 B.n798 585
R786 B.n798 B.n65 585
R787 B.n797 B.n64 585
R788 B.n847 B.n64 585
R789 B.n796 B.n63 585
R790 B.n848 B.n63 585
R791 B.n795 B.n62 585
R792 B.n849 B.n62 585
R793 B.n794 B.n793 585
R794 B.n793 B.n61 585
R795 B.n792 B.n57 585
R796 B.n855 B.n57 585
R797 B.n791 B.n56 585
R798 B.n856 B.n56 585
R799 B.n790 B.n55 585
R800 B.n857 B.n55 585
R801 B.n789 B.n788 585
R802 B.n788 B.n51 585
R803 B.n787 B.n50 585
R804 B.n863 B.n50 585
R805 B.n786 B.n49 585
R806 B.n864 B.n49 585
R807 B.n785 B.n48 585
R808 B.n865 B.n48 585
R809 B.n784 B.n783 585
R810 B.n783 B.n44 585
R811 B.n782 B.n43 585
R812 B.n871 B.n43 585
R813 B.n781 B.n42 585
R814 B.n872 B.n42 585
R815 B.n780 B.n41 585
R816 B.n873 B.n41 585
R817 B.n779 B.n778 585
R818 B.n778 B.n37 585
R819 B.n777 B.n36 585
R820 B.n879 B.n36 585
R821 B.n776 B.n35 585
R822 B.n880 B.n35 585
R823 B.n775 B.n34 585
R824 B.n881 B.n34 585
R825 B.n774 B.n773 585
R826 B.n773 B.n30 585
R827 B.n772 B.n29 585
R828 B.n887 B.n29 585
R829 B.n771 B.n28 585
R830 B.n888 B.n28 585
R831 B.n770 B.n27 585
R832 B.n889 B.n27 585
R833 B.n769 B.n768 585
R834 B.n768 B.n26 585
R835 B.n767 B.n22 585
R836 B.n895 B.n22 585
R837 B.n766 B.n21 585
R838 B.n896 B.n21 585
R839 B.n765 B.n20 585
R840 B.n897 B.n20 585
R841 B.n764 B.n763 585
R842 B.n763 B.n16 585
R843 B.n762 B.n15 585
R844 B.n903 B.n15 585
R845 B.n761 B.n14 585
R846 B.n904 B.n14 585
R847 B.n760 B.n13 585
R848 B.n905 B.n13 585
R849 B.n759 B.n758 585
R850 B.n758 B.n12 585
R851 B.n757 B.n756 585
R852 B.n757 B.n8 585
R853 B.n755 B.n7 585
R854 B.n912 B.n7 585
R855 B.n754 B.n6 585
R856 B.n913 B.n6 585
R857 B.n753 B.n5 585
R858 B.n914 B.n5 585
R859 B.n752 B.n751 585
R860 B.n751 B.n4 585
R861 B.n750 B.n302 585
R862 B.n750 B.n749 585
R863 B.n740 B.n303 585
R864 B.n304 B.n303 585
R865 B.n742 B.n741 585
R866 B.n743 B.n742 585
R867 B.n739 B.n308 585
R868 B.n312 B.n308 585
R869 B.n738 B.n737 585
R870 B.n737 B.n736 585
R871 B.n310 B.n309 585
R872 B.n311 B.n310 585
R873 B.n729 B.n728 585
R874 B.n730 B.n729 585
R875 B.n727 B.n317 585
R876 B.n317 B.n316 585
R877 B.n726 B.n725 585
R878 B.n725 B.n724 585
R879 B.n319 B.n318 585
R880 B.n717 B.n319 585
R881 B.n716 B.n715 585
R882 B.n718 B.n716 585
R883 B.n714 B.n324 585
R884 B.n324 B.n323 585
R885 B.n713 B.n712 585
R886 B.n712 B.n711 585
R887 B.n326 B.n325 585
R888 B.n327 B.n326 585
R889 B.n704 B.n703 585
R890 B.n705 B.n704 585
R891 B.n702 B.n332 585
R892 B.n332 B.n331 585
R893 B.n701 B.n700 585
R894 B.n700 B.n699 585
R895 B.n334 B.n333 585
R896 B.n335 B.n334 585
R897 B.n692 B.n691 585
R898 B.n693 B.n692 585
R899 B.n690 B.n340 585
R900 B.n340 B.n339 585
R901 B.n689 B.n688 585
R902 B.n688 B.n687 585
R903 B.n342 B.n341 585
R904 B.n343 B.n342 585
R905 B.n680 B.n679 585
R906 B.n681 B.n680 585
R907 B.n678 B.n347 585
R908 B.n351 B.n347 585
R909 B.n677 B.n676 585
R910 B.n676 B.n675 585
R911 B.n349 B.n348 585
R912 B.n350 B.n349 585
R913 B.n668 B.n667 585
R914 B.n669 B.n668 585
R915 B.n666 B.n356 585
R916 B.n356 B.n355 585
R917 B.n665 B.n664 585
R918 B.n664 B.n663 585
R919 B.n358 B.n357 585
R920 B.n656 B.n358 585
R921 B.n655 B.n654 585
R922 B.n657 B.n655 585
R923 B.n653 B.n363 585
R924 B.n363 B.n362 585
R925 B.n652 B.n651 585
R926 B.n651 B.n650 585
R927 B.n365 B.n364 585
R928 B.n366 B.n365 585
R929 B.n643 B.n642 585
R930 B.n644 B.n643 585
R931 B.n641 B.n371 585
R932 B.n371 B.n370 585
R933 B.n640 B.n639 585
R934 B.n639 B.n638 585
R935 B.n373 B.n372 585
R936 B.n374 B.n373 585
R937 B.n631 B.n630 585
R938 B.n632 B.n631 585
R939 B.n629 B.n378 585
R940 B.n382 B.n378 585
R941 B.n628 B.n627 585
R942 B.n627 B.n626 585
R943 B.n380 B.n379 585
R944 B.n381 B.n380 585
R945 B.n619 B.n618 585
R946 B.n620 B.n619 585
R947 B.n617 B.n387 585
R948 B.n387 B.n386 585
R949 B.n616 B.n615 585
R950 B.n615 B.n614 585
R951 B.n389 B.n388 585
R952 B.n390 B.n389 585
R953 B.n610 B.n609 585
R954 B.n393 B.n392 585
R955 B.n606 B.n605 585
R956 B.n607 B.n606 585
R957 B.n604 B.n435 585
R958 B.n603 B.n602 585
R959 B.n601 B.n600 585
R960 B.n599 B.n598 585
R961 B.n597 B.n596 585
R962 B.n595 B.n594 585
R963 B.n593 B.n592 585
R964 B.n591 B.n590 585
R965 B.n589 B.n588 585
R966 B.n587 B.n586 585
R967 B.n585 B.n584 585
R968 B.n583 B.n582 585
R969 B.n581 B.n580 585
R970 B.n579 B.n578 585
R971 B.n577 B.n576 585
R972 B.n575 B.n574 585
R973 B.n573 B.n572 585
R974 B.n571 B.n570 585
R975 B.n569 B.n568 585
R976 B.n567 B.n566 585
R977 B.n565 B.n564 585
R978 B.n563 B.n562 585
R979 B.n561 B.n560 585
R980 B.n559 B.n558 585
R981 B.n557 B.n556 585
R982 B.n555 B.n554 585
R983 B.n553 B.n552 585
R984 B.n551 B.n550 585
R985 B.n549 B.n548 585
R986 B.n547 B.n546 585
R987 B.n545 B.n544 585
R988 B.n543 B.n542 585
R989 B.n541 B.n540 585
R990 B.n539 B.n538 585
R991 B.n537 B.n536 585
R992 B.n534 B.n533 585
R993 B.n532 B.n531 585
R994 B.n530 B.n529 585
R995 B.n528 B.n527 585
R996 B.n526 B.n525 585
R997 B.n524 B.n523 585
R998 B.n522 B.n521 585
R999 B.n520 B.n519 585
R1000 B.n518 B.n517 585
R1001 B.n516 B.n515 585
R1002 B.n514 B.n513 585
R1003 B.n512 B.n511 585
R1004 B.n510 B.n509 585
R1005 B.n508 B.n507 585
R1006 B.n506 B.n505 585
R1007 B.n504 B.n503 585
R1008 B.n502 B.n501 585
R1009 B.n500 B.n499 585
R1010 B.n498 B.n497 585
R1011 B.n496 B.n495 585
R1012 B.n494 B.n493 585
R1013 B.n492 B.n491 585
R1014 B.n490 B.n489 585
R1015 B.n488 B.n487 585
R1016 B.n486 B.n485 585
R1017 B.n484 B.n483 585
R1018 B.n482 B.n481 585
R1019 B.n480 B.n479 585
R1020 B.n478 B.n477 585
R1021 B.n476 B.n475 585
R1022 B.n474 B.n473 585
R1023 B.n472 B.n471 585
R1024 B.n470 B.n469 585
R1025 B.n468 B.n467 585
R1026 B.n466 B.n465 585
R1027 B.n464 B.n463 585
R1028 B.n462 B.n461 585
R1029 B.n460 B.n459 585
R1030 B.n458 B.n457 585
R1031 B.n456 B.n455 585
R1032 B.n454 B.n453 585
R1033 B.n452 B.n451 585
R1034 B.n450 B.n449 585
R1035 B.n448 B.n447 585
R1036 B.n446 B.n445 585
R1037 B.n444 B.n443 585
R1038 B.n442 B.n441 585
R1039 B.n611 B.n391 585
R1040 B.n391 B.n390 585
R1041 B.n613 B.n612 585
R1042 B.n614 B.n613 585
R1043 B.n385 B.n384 585
R1044 B.n386 B.n385 585
R1045 B.n622 B.n621 585
R1046 B.n621 B.n620 585
R1047 B.n623 B.n383 585
R1048 B.n383 B.n381 585
R1049 B.n625 B.n624 585
R1050 B.n626 B.n625 585
R1051 B.n377 B.n376 585
R1052 B.n382 B.n377 585
R1053 B.n634 B.n633 585
R1054 B.n633 B.n632 585
R1055 B.n635 B.n375 585
R1056 B.n375 B.n374 585
R1057 B.n637 B.n636 585
R1058 B.n638 B.n637 585
R1059 B.n369 B.n368 585
R1060 B.n370 B.n369 585
R1061 B.n646 B.n645 585
R1062 B.n645 B.n644 585
R1063 B.n647 B.n367 585
R1064 B.n367 B.n366 585
R1065 B.n649 B.n648 585
R1066 B.n650 B.n649 585
R1067 B.n361 B.n360 585
R1068 B.n362 B.n361 585
R1069 B.n659 B.n658 585
R1070 B.n658 B.n657 585
R1071 B.n660 B.n359 585
R1072 B.n656 B.n359 585
R1073 B.n662 B.n661 585
R1074 B.n663 B.n662 585
R1075 B.n354 B.n353 585
R1076 B.n355 B.n354 585
R1077 B.n671 B.n670 585
R1078 B.n670 B.n669 585
R1079 B.n672 B.n352 585
R1080 B.n352 B.n350 585
R1081 B.n674 B.n673 585
R1082 B.n675 B.n674 585
R1083 B.n346 B.n345 585
R1084 B.n351 B.n346 585
R1085 B.n683 B.n682 585
R1086 B.n682 B.n681 585
R1087 B.n684 B.n344 585
R1088 B.n344 B.n343 585
R1089 B.n686 B.n685 585
R1090 B.n687 B.n686 585
R1091 B.n338 B.n337 585
R1092 B.n339 B.n338 585
R1093 B.n695 B.n694 585
R1094 B.n694 B.n693 585
R1095 B.n696 B.n336 585
R1096 B.n336 B.n335 585
R1097 B.n698 B.n697 585
R1098 B.n699 B.n698 585
R1099 B.n330 B.n329 585
R1100 B.n331 B.n330 585
R1101 B.n707 B.n706 585
R1102 B.n706 B.n705 585
R1103 B.n708 B.n328 585
R1104 B.n328 B.n327 585
R1105 B.n710 B.n709 585
R1106 B.n711 B.n710 585
R1107 B.n322 B.n321 585
R1108 B.n323 B.n322 585
R1109 B.n720 B.n719 585
R1110 B.n719 B.n718 585
R1111 B.n721 B.n320 585
R1112 B.n717 B.n320 585
R1113 B.n723 B.n722 585
R1114 B.n724 B.n723 585
R1115 B.n315 B.n314 585
R1116 B.n316 B.n315 585
R1117 B.n732 B.n731 585
R1118 B.n731 B.n730 585
R1119 B.n733 B.n313 585
R1120 B.n313 B.n311 585
R1121 B.n735 B.n734 585
R1122 B.n736 B.n735 585
R1123 B.n307 B.n306 585
R1124 B.n312 B.n307 585
R1125 B.n745 B.n744 585
R1126 B.n744 B.n743 585
R1127 B.n746 B.n305 585
R1128 B.n305 B.n304 585
R1129 B.n748 B.n747 585
R1130 B.n749 B.n748 585
R1131 B.n3 B.n0 585
R1132 B.n4 B.n3 585
R1133 B.n911 B.n1 585
R1134 B.n912 B.n911 585
R1135 B.n910 B.n909 585
R1136 B.n910 B.n8 585
R1137 B.n908 B.n9 585
R1138 B.n12 B.n9 585
R1139 B.n907 B.n906 585
R1140 B.n906 B.n905 585
R1141 B.n11 B.n10 585
R1142 B.n904 B.n11 585
R1143 B.n902 B.n901 585
R1144 B.n903 B.n902 585
R1145 B.n900 B.n17 585
R1146 B.n17 B.n16 585
R1147 B.n899 B.n898 585
R1148 B.n898 B.n897 585
R1149 B.n19 B.n18 585
R1150 B.n896 B.n19 585
R1151 B.n894 B.n893 585
R1152 B.n895 B.n894 585
R1153 B.n892 B.n23 585
R1154 B.n26 B.n23 585
R1155 B.n891 B.n890 585
R1156 B.n890 B.n889 585
R1157 B.n25 B.n24 585
R1158 B.n888 B.n25 585
R1159 B.n886 B.n885 585
R1160 B.n887 B.n886 585
R1161 B.n884 B.n31 585
R1162 B.n31 B.n30 585
R1163 B.n883 B.n882 585
R1164 B.n882 B.n881 585
R1165 B.n33 B.n32 585
R1166 B.n880 B.n33 585
R1167 B.n878 B.n877 585
R1168 B.n879 B.n878 585
R1169 B.n876 B.n38 585
R1170 B.n38 B.n37 585
R1171 B.n875 B.n874 585
R1172 B.n874 B.n873 585
R1173 B.n40 B.n39 585
R1174 B.n872 B.n40 585
R1175 B.n870 B.n869 585
R1176 B.n871 B.n870 585
R1177 B.n868 B.n45 585
R1178 B.n45 B.n44 585
R1179 B.n867 B.n866 585
R1180 B.n866 B.n865 585
R1181 B.n47 B.n46 585
R1182 B.n864 B.n47 585
R1183 B.n862 B.n861 585
R1184 B.n863 B.n862 585
R1185 B.n860 B.n52 585
R1186 B.n52 B.n51 585
R1187 B.n859 B.n858 585
R1188 B.n858 B.n857 585
R1189 B.n54 B.n53 585
R1190 B.n856 B.n54 585
R1191 B.n854 B.n853 585
R1192 B.n855 B.n854 585
R1193 B.n852 B.n58 585
R1194 B.n61 B.n58 585
R1195 B.n851 B.n850 585
R1196 B.n850 B.n849 585
R1197 B.n60 B.n59 585
R1198 B.n848 B.n60 585
R1199 B.n846 B.n845 585
R1200 B.n847 B.n846 585
R1201 B.n844 B.n66 585
R1202 B.n66 B.n65 585
R1203 B.n843 B.n842 585
R1204 B.n842 B.n841 585
R1205 B.n68 B.n67 585
R1206 B.n840 B.n68 585
R1207 B.n838 B.n837 585
R1208 B.n839 B.n838 585
R1209 B.n836 B.n73 585
R1210 B.n73 B.n72 585
R1211 B.n835 B.n834 585
R1212 B.n834 B.n833 585
R1213 B.n75 B.n74 585
R1214 B.n832 B.n75 585
R1215 B.n830 B.n829 585
R1216 B.n831 B.n830 585
R1217 B.n828 B.n80 585
R1218 B.n80 B.n79 585
R1219 B.n827 B.n826 585
R1220 B.n826 B.n825 585
R1221 B.n82 B.n81 585
R1222 B.n824 B.n82 585
R1223 B.n822 B.n821 585
R1224 B.n823 B.n822 585
R1225 B.n820 B.n87 585
R1226 B.n87 B.n86 585
R1227 B.n915 B.n914 585
R1228 B.n913 B.n2 585
R1229 B.n818 B.n87 521.33
R1230 B.n815 B.n132 521.33
R1231 B.n441 B.n389 521.33
R1232 B.n609 B.n391 521.33
R1233 B.n135 B.t10 342.774
R1234 B.n133 B.t21 342.774
R1235 B.n438 B.t18 342.774
R1236 B.n436 B.t14 342.774
R1237 B.n133 B.t22 303.577
R1238 B.n438 B.t20 303.577
R1239 B.n135 B.t12 303.577
R1240 B.n436 B.t17 303.577
R1241 B.n134 B.t23 260.329
R1242 B.n439 B.t19 260.329
R1243 B.n136 B.t13 260.329
R1244 B.n437 B.t16 260.329
R1245 B.n816 B.n130 256.663
R1246 B.n816 B.n129 256.663
R1247 B.n816 B.n128 256.663
R1248 B.n816 B.n127 256.663
R1249 B.n816 B.n126 256.663
R1250 B.n816 B.n125 256.663
R1251 B.n816 B.n124 256.663
R1252 B.n816 B.n123 256.663
R1253 B.n816 B.n122 256.663
R1254 B.n816 B.n121 256.663
R1255 B.n816 B.n120 256.663
R1256 B.n816 B.n119 256.663
R1257 B.n816 B.n118 256.663
R1258 B.n816 B.n117 256.663
R1259 B.n816 B.n116 256.663
R1260 B.n816 B.n115 256.663
R1261 B.n816 B.n114 256.663
R1262 B.n816 B.n113 256.663
R1263 B.n816 B.n112 256.663
R1264 B.n816 B.n111 256.663
R1265 B.n816 B.n110 256.663
R1266 B.n816 B.n109 256.663
R1267 B.n816 B.n108 256.663
R1268 B.n816 B.n107 256.663
R1269 B.n816 B.n106 256.663
R1270 B.n816 B.n105 256.663
R1271 B.n816 B.n104 256.663
R1272 B.n816 B.n103 256.663
R1273 B.n816 B.n102 256.663
R1274 B.n816 B.n101 256.663
R1275 B.n816 B.n100 256.663
R1276 B.n816 B.n99 256.663
R1277 B.n816 B.n98 256.663
R1278 B.n816 B.n97 256.663
R1279 B.n816 B.n96 256.663
R1280 B.n816 B.n95 256.663
R1281 B.n816 B.n94 256.663
R1282 B.n816 B.n93 256.663
R1283 B.n816 B.n92 256.663
R1284 B.n816 B.n91 256.663
R1285 B.n816 B.n90 256.663
R1286 B.n817 B.n816 256.663
R1287 B.n608 B.n607 256.663
R1288 B.n607 B.n394 256.663
R1289 B.n607 B.n395 256.663
R1290 B.n607 B.n396 256.663
R1291 B.n607 B.n397 256.663
R1292 B.n607 B.n398 256.663
R1293 B.n607 B.n399 256.663
R1294 B.n607 B.n400 256.663
R1295 B.n607 B.n401 256.663
R1296 B.n607 B.n402 256.663
R1297 B.n607 B.n403 256.663
R1298 B.n607 B.n404 256.663
R1299 B.n607 B.n405 256.663
R1300 B.n607 B.n406 256.663
R1301 B.n607 B.n407 256.663
R1302 B.n607 B.n408 256.663
R1303 B.n607 B.n409 256.663
R1304 B.n607 B.n410 256.663
R1305 B.n607 B.n411 256.663
R1306 B.n607 B.n412 256.663
R1307 B.n607 B.n413 256.663
R1308 B.n607 B.n414 256.663
R1309 B.n607 B.n415 256.663
R1310 B.n607 B.n416 256.663
R1311 B.n607 B.n417 256.663
R1312 B.n607 B.n418 256.663
R1313 B.n607 B.n419 256.663
R1314 B.n607 B.n420 256.663
R1315 B.n607 B.n421 256.663
R1316 B.n607 B.n422 256.663
R1317 B.n607 B.n423 256.663
R1318 B.n607 B.n424 256.663
R1319 B.n607 B.n425 256.663
R1320 B.n607 B.n426 256.663
R1321 B.n607 B.n427 256.663
R1322 B.n607 B.n428 256.663
R1323 B.n607 B.n429 256.663
R1324 B.n607 B.n430 256.663
R1325 B.n607 B.n431 256.663
R1326 B.n607 B.n432 256.663
R1327 B.n607 B.n433 256.663
R1328 B.n607 B.n434 256.663
R1329 B.n917 B.n916 256.663
R1330 B.n138 B.n89 163.367
R1331 B.n142 B.n141 163.367
R1332 B.n146 B.n145 163.367
R1333 B.n150 B.n149 163.367
R1334 B.n154 B.n153 163.367
R1335 B.n158 B.n157 163.367
R1336 B.n162 B.n161 163.367
R1337 B.n166 B.n165 163.367
R1338 B.n170 B.n169 163.367
R1339 B.n174 B.n173 163.367
R1340 B.n178 B.n177 163.367
R1341 B.n182 B.n181 163.367
R1342 B.n186 B.n185 163.367
R1343 B.n190 B.n189 163.367
R1344 B.n194 B.n193 163.367
R1345 B.n198 B.n197 163.367
R1346 B.n202 B.n201 163.367
R1347 B.n206 B.n205 163.367
R1348 B.n210 B.n209 163.367
R1349 B.n214 B.n213 163.367
R1350 B.n218 B.n217 163.367
R1351 B.n222 B.n221 163.367
R1352 B.n226 B.n225 163.367
R1353 B.n231 B.n230 163.367
R1354 B.n235 B.n234 163.367
R1355 B.n239 B.n238 163.367
R1356 B.n243 B.n242 163.367
R1357 B.n247 B.n246 163.367
R1358 B.n251 B.n250 163.367
R1359 B.n255 B.n254 163.367
R1360 B.n259 B.n258 163.367
R1361 B.n263 B.n262 163.367
R1362 B.n267 B.n266 163.367
R1363 B.n271 B.n270 163.367
R1364 B.n275 B.n274 163.367
R1365 B.n279 B.n278 163.367
R1366 B.n283 B.n282 163.367
R1367 B.n287 B.n286 163.367
R1368 B.n291 B.n290 163.367
R1369 B.n295 B.n294 163.367
R1370 B.n299 B.n298 163.367
R1371 B.n815 B.n131 163.367
R1372 B.n615 B.n389 163.367
R1373 B.n615 B.n387 163.367
R1374 B.n619 B.n387 163.367
R1375 B.n619 B.n380 163.367
R1376 B.n627 B.n380 163.367
R1377 B.n627 B.n378 163.367
R1378 B.n631 B.n378 163.367
R1379 B.n631 B.n373 163.367
R1380 B.n639 B.n373 163.367
R1381 B.n639 B.n371 163.367
R1382 B.n643 B.n371 163.367
R1383 B.n643 B.n365 163.367
R1384 B.n651 B.n365 163.367
R1385 B.n651 B.n363 163.367
R1386 B.n655 B.n363 163.367
R1387 B.n655 B.n358 163.367
R1388 B.n664 B.n358 163.367
R1389 B.n664 B.n356 163.367
R1390 B.n668 B.n356 163.367
R1391 B.n668 B.n349 163.367
R1392 B.n676 B.n349 163.367
R1393 B.n676 B.n347 163.367
R1394 B.n680 B.n347 163.367
R1395 B.n680 B.n342 163.367
R1396 B.n688 B.n342 163.367
R1397 B.n688 B.n340 163.367
R1398 B.n692 B.n340 163.367
R1399 B.n692 B.n334 163.367
R1400 B.n700 B.n334 163.367
R1401 B.n700 B.n332 163.367
R1402 B.n704 B.n332 163.367
R1403 B.n704 B.n326 163.367
R1404 B.n712 B.n326 163.367
R1405 B.n712 B.n324 163.367
R1406 B.n716 B.n324 163.367
R1407 B.n716 B.n319 163.367
R1408 B.n725 B.n319 163.367
R1409 B.n725 B.n317 163.367
R1410 B.n729 B.n317 163.367
R1411 B.n729 B.n310 163.367
R1412 B.n737 B.n310 163.367
R1413 B.n737 B.n308 163.367
R1414 B.n742 B.n308 163.367
R1415 B.n742 B.n303 163.367
R1416 B.n750 B.n303 163.367
R1417 B.n751 B.n750 163.367
R1418 B.n751 B.n5 163.367
R1419 B.n6 B.n5 163.367
R1420 B.n7 B.n6 163.367
R1421 B.n757 B.n7 163.367
R1422 B.n758 B.n757 163.367
R1423 B.n758 B.n13 163.367
R1424 B.n14 B.n13 163.367
R1425 B.n15 B.n14 163.367
R1426 B.n763 B.n15 163.367
R1427 B.n763 B.n20 163.367
R1428 B.n21 B.n20 163.367
R1429 B.n22 B.n21 163.367
R1430 B.n768 B.n22 163.367
R1431 B.n768 B.n27 163.367
R1432 B.n28 B.n27 163.367
R1433 B.n29 B.n28 163.367
R1434 B.n773 B.n29 163.367
R1435 B.n773 B.n34 163.367
R1436 B.n35 B.n34 163.367
R1437 B.n36 B.n35 163.367
R1438 B.n778 B.n36 163.367
R1439 B.n778 B.n41 163.367
R1440 B.n42 B.n41 163.367
R1441 B.n43 B.n42 163.367
R1442 B.n783 B.n43 163.367
R1443 B.n783 B.n48 163.367
R1444 B.n49 B.n48 163.367
R1445 B.n50 B.n49 163.367
R1446 B.n788 B.n50 163.367
R1447 B.n788 B.n55 163.367
R1448 B.n56 B.n55 163.367
R1449 B.n57 B.n56 163.367
R1450 B.n793 B.n57 163.367
R1451 B.n793 B.n62 163.367
R1452 B.n63 B.n62 163.367
R1453 B.n64 B.n63 163.367
R1454 B.n798 B.n64 163.367
R1455 B.n798 B.n69 163.367
R1456 B.n70 B.n69 163.367
R1457 B.n71 B.n70 163.367
R1458 B.n803 B.n71 163.367
R1459 B.n803 B.n76 163.367
R1460 B.n77 B.n76 163.367
R1461 B.n78 B.n77 163.367
R1462 B.n808 B.n78 163.367
R1463 B.n808 B.n83 163.367
R1464 B.n84 B.n83 163.367
R1465 B.n85 B.n84 163.367
R1466 B.n132 B.n85 163.367
R1467 B.n606 B.n393 163.367
R1468 B.n606 B.n435 163.367
R1469 B.n602 B.n601 163.367
R1470 B.n598 B.n597 163.367
R1471 B.n594 B.n593 163.367
R1472 B.n590 B.n589 163.367
R1473 B.n586 B.n585 163.367
R1474 B.n582 B.n581 163.367
R1475 B.n578 B.n577 163.367
R1476 B.n574 B.n573 163.367
R1477 B.n570 B.n569 163.367
R1478 B.n566 B.n565 163.367
R1479 B.n562 B.n561 163.367
R1480 B.n558 B.n557 163.367
R1481 B.n554 B.n553 163.367
R1482 B.n550 B.n549 163.367
R1483 B.n546 B.n545 163.367
R1484 B.n542 B.n541 163.367
R1485 B.n538 B.n537 163.367
R1486 B.n533 B.n532 163.367
R1487 B.n529 B.n528 163.367
R1488 B.n525 B.n524 163.367
R1489 B.n521 B.n520 163.367
R1490 B.n517 B.n516 163.367
R1491 B.n513 B.n512 163.367
R1492 B.n509 B.n508 163.367
R1493 B.n505 B.n504 163.367
R1494 B.n501 B.n500 163.367
R1495 B.n497 B.n496 163.367
R1496 B.n493 B.n492 163.367
R1497 B.n489 B.n488 163.367
R1498 B.n485 B.n484 163.367
R1499 B.n481 B.n480 163.367
R1500 B.n477 B.n476 163.367
R1501 B.n473 B.n472 163.367
R1502 B.n469 B.n468 163.367
R1503 B.n465 B.n464 163.367
R1504 B.n461 B.n460 163.367
R1505 B.n457 B.n456 163.367
R1506 B.n453 B.n452 163.367
R1507 B.n449 B.n448 163.367
R1508 B.n445 B.n444 163.367
R1509 B.n613 B.n391 163.367
R1510 B.n613 B.n385 163.367
R1511 B.n621 B.n385 163.367
R1512 B.n621 B.n383 163.367
R1513 B.n625 B.n383 163.367
R1514 B.n625 B.n377 163.367
R1515 B.n633 B.n377 163.367
R1516 B.n633 B.n375 163.367
R1517 B.n637 B.n375 163.367
R1518 B.n637 B.n369 163.367
R1519 B.n645 B.n369 163.367
R1520 B.n645 B.n367 163.367
R1521 B.n649 B.n367 163.367
R1522 B.n649 B.n361 163.367
R1523 B.n658 B.n361 163.367
R1524 B.n658 B.n359 163.367
R1525 B.n662 B.n359 163.367
R1526 B.n662 B.n354 163.367
R1527 B.n670 B.n354 163.367
R1528 B.n670 B.n352 163.367
R1529 B.n674 B.n352 163.367
R1530 B.n674 B.n346 163.367
R1531 B.n682 B.n346 163.367
R1532 B.n682 B.n344 163.367
R1533 B.n686 B.n344 163.367
R1534 B.n686 B.n338 163.367
R1535 B.n694 B.n338 163.367
R1536 B.n694 B.n336 163.367
R1537 B.n698 B.n336 163.367
R1538 B.n698 B.n330 163.367
R1539 B.n706 B.n330 163.367
R1540 B.n706 B.n328 163.367
R1541 B.n710 B.n328 163.367
R1542 B.n710 B.n322 163.367
R1543 B.n719 B.n322 163.367
R1544 B.n719 B.n320 163.367
R1545 B.n723 B.n320 163.367
R1546 B.n723 B.n315 163.367
R1547 B.n731 B.n315 163.367
R1548 B.n731 B.n313 163.367
R1549 B.n735 B.n313 163.367
R1550 B.n735 B.n307 163.367
R1551 B.n744 B.n307 163.367
R1552 B.n744 B.n305 163.367
R1553 B.n748 B.n305 163.367
R1554 B.n748 B.n3 163.367
R1555 B.n915 B.n3 163.367
R1556 B.n911 B.n2 163.367
R1557 B.n911 B.n910 163.367
R1558 B.n910 B.n9 163.367
R1559 B.n906 B.n9 163.367
R1560 B.n906 B.n11 163.367
R1561 B.n902 B.n11 163.367
R1562 B.n902 B.n17 163.367
R1563 B.n898 B.n17 163.367
R1564 B.n898 B.n19 163.367
R1565 B.n894 B.n19 163.367
R1566 B.n894 B.n23 163.367
R1567 B.n890 B.n23 163.367
R1568 B.n890 B.n25 163.367
R1569 B.n886 B.n25 163.367
R1570 B.n886 B.n31 163.367
R1571 B.n882 B.n31 163.367
R1572 B.n882 B.n33 163.367
R1573 B.n878 B.n33 163.367
R1574 B.n878 B.n38 163.367
R1575 B.n874 B.n38 163.367
R1576 B.n874 B.n40 163.367
R1577 B.n870 B.n40 163.367
R1578 B.n870 B.n45 163.367
R1579 B.n866 B.n45 163.367
R1580 B.n866 B.n47 163.367
R1581 B.n862 B.n47 163.367
R1582 B.n862 B.n52 163.367
R1583 B.n858 B.n52 163.367
R1584 B.n858 B.n54 163.367
R1585 B.n854 B.n54 163.367
R1586 B.n854 B.n58 163.367
R1587 B.n850 B.n58 163.367
R1588 B.n850 B.n60 163.367
R1589 B.n846 B.n60 163.367
R1590 B.n846 B.n66 163.367
R1591 B.n842 B.n66 163.367
R1592 B.n842 B.n68 163.367
R1593 B.n838 B.n68 163.367
R1594 B.n838 B.n73 163.367
R1595 B.n834 B.n73 163.367
R1596 B.n834 B.n75 163.367
R1597 B.n830 B.n75 163.367
R1598 B.n830 B.n80 163.367
R1599 B.n826 B.n80 163.367
R1600 B.n826 B.n82 163.367
R1601 B.n822 B.n82 163.367
R1602 B.n822 B.n87 163.367
R1603 B.n607 B.n390 83.162
R1604 B.n816 B.n86 83.162
R1605 B.n818 B.n817 71.676
R1606 B.n138 B.n90 71.676
R1607 B.n142 B.n91 71.676
R1608 B.n146 B.n92 71.676
R1609 B.n150 B.n93 71.676
R1610 B.n154 B.n94 71.676
R1611 B.n158 B.n95 71.676
R1612 B.n162 B.n96 71.676
R1613 B.n166 B.n97 71.676
R1614 B.n170 B.n98 71.676
R1615 B.n174 B.n99 71.676
R1616 B.n178 B.n100 71.676
R1617 B.n182 B.n101 71.676
R1618 B.n186 B.n102 71.676
R1619 B.n190 B.n103 71.676
R1620 B.n194 B.n104 71.676
R1621 B.n198 B.n105 71.676
R1622 B.n202 B.n106 71.676
R1623 B.n206 B.n107 71.676
R1624 B.n210 B.n108 71.676
R1625 B.n214 B.n109 71.676
R1626 B.n218 B.n110 71.676
R1627 B.n222 B.n111 71.676
R1628 B.n226 B.n112 71.676
R1629 B.n231 B.n113 71.676
R1630 B.n235 B.n114 71.676
R1631 B.n239 B.n115 71.676
R1632 B.n243 B.n116 71.676
R1633 B.n247 B.n117 71.676
R1634 B.n251 B.n118 71.676
R1635 B.n255 B.n119 71.676
R1636 B.n259 B.n120 71.676
R1637 B.n263 B.n121 71.676
R1638 B.n267 B.n122 71.676
R1639 B.n271 B.n123 71.676
R1640 B.n275 B.n124 71.676
R1641 B.n279 B.n125 71.676
R1642 B.n283 B.n126 71.676
R1643 B.n287 B.n127 71.676
R1644 B.n291 B.n128 71.676
R1645 B.n295 B.n129 71.676
R1646 B.n299 B.n130 71.676
R1647 B.n131 B.n130 71.676
R1648 B.n298 B.n129 71.676
R1649 B.n294 B.n128 71.676
R1650 B.n290 B.n127 71.676
R1651 B.n286 B.n126 71.676
R1652 B.n282 B.n125 71.676
R1653 B.n278 B.n124 71.676
R1654 B.n274 B.n123 71.676
R1655 B.n270 B.n122 71.676
R1656 B.n266 B.n121 71.676
R1657 B.n262 B.n120 71.676
R1658 B.n258 B.n119 71.676
R1659 B.n254 B.n118 71.676
R1660 B.n250 B.n117 71.676
R1661 B.n246 B.n116 71.676
R1662 B.n242 B.n115 71.676
R1663 B.n238 B.n114 71.676
R1664 B.n234 B.n113 71.676
R1665 B.n230 B.n112 71.676
R1666 B.n225 B.n111 71.676
R1667 B.n221 B.n110 71.676
R1668 B.n217 B.n109 71.676
R1669 B.n213 B.n108 71.676
R1670 B.n209 B.n107 71.676
R1671 B.n205 B.n106 71.676
R1672 B.n201 B.n105 71.676
R1673 B.n197 B.n104 71.676
R1674 B.n193 B.n103 71.676
R1675 B.n189 B.n102 71.676
R1676 B.n185 B.n101 71.676
R1677 B.n181 B.n100 71.676
R1678 B.n177 B.n99 71.676
R1679 B.n173 B.n98 71.676
R1680 B.n169 B.n97 71.676
R1681 B.n165 B.n96 71.676
R1682 B.n161 B.n95 71.676
R1683 B.n157 B.n94 71.676
R1684 B.n153 B.n93 71.676
R1685 B.n149 B.n92 71.676
R1686 B.n145 B.n91 71.676
R1687 B.n141 B.n90 71.676
R1688 B.n817 B.n89 71.676
R1689 B.n609 B.n608 71.676
R1690 B.n435 B.n394 71.676
R1691 B.n601 B.n395 71.676
R1692 B.n597 B.n396 71.676
R1693 B.n593 B.n397 71.676
R1694 B.n589 B.n398 71.676
R1695 B.n585 B.n399 71.676
R1696 B.n581 B.n400 71.676
R1697 B.n577 B.n401 71.676
R1698 B.n573 B.n402 71.676
R1699 B.n569 B.n403 71.676
R1700 B.n565 B.n404 71.676
R1701 B.n561 B.n405 71.676
R1702 B.n557 B.n406 71.676
R1703 B.n553 B.n407 71.676
R1704 B.n549 B.n408 71.676
R1705 B.n545 B.n409 71.676
R1706 B.n541 B.n410 71.676
R1707 B.n537 B.n411 71.676
R1708 B.n532 B.n412 71.676
R1709 B.n528 B.n413 71.676
R1710 B.n524 B.n414 71.676
R1711 B.n520 B.n415 71.676
R1712 B.n516 B.n416 71.676
R1713 B.n512 B.n417 71.676
R1714 B.n508 B.n418 71.676
R1715 B.n504 B.n419 71.676
R1716 B.n500 B.n420 71.676
R1717 B.n496 B.n421 71.676
R1718 B.n492 B.n422 71.676
R1719 B.n488 B.n423 71.676
R1720 B.n484 B.n424 71.676
R1721 B.n480 B.n425 71.676
R1722 B.n476 B.n426 71.676
R1723 B.n472 B.n427 71.676
R1724 B.n468 B.n428 71.676
R1725 B.n464 B.n429 71.676
R1726 B.n460 B.n430 71.676
R1727 B.n456 B.n431 71.676
R1728 B.n452 B.n432 71.676
R1729 B.n448 B.n433 71.676
R1730 B.n444 B.n434 71.676
R1731 B.n608 B.n393 71.676
R1732 B.n602 B.n394 71.676
R1733 B.n598 B.n395 71.676
R1734 B.n594 B.n396 71.676
R1735 B.n590 B.n397 71.676
R1736 B.n586 B.n398 71.676
R1737 B.n582 B.n399 71.676
R1738 B.n578 B.n400 71.676
R1739 B.n574 B.n401 71.676
R1740 B.n570 B.n402 71.676
R1741 B.n566 B.n403 71.676
R1742 B.n562 B.n404 71.676
R1743 B.n558 B.n405 71.676
R1744 B.n554 B.n406 71.676
R1745 B.n550 B.n407 71.676
R1746 B.n546 B.n408 71.676
R1747 B.n542 B.n409 71.676
R1748 B.n538 B.n410 71.676
R1749 B.n533 B.n411 71.676
R1750 B.n529 B.n412 71.676
R1751 B.n525 B.n413 71.676
R1752 B.n521 B.n414 71.676
R1753 B.n517 B.n415 71.676
R1754 B.n513 B.n416 71.676
R1755 B.n509 B.n417 71.676
R1756 B.n505 B.n418 71.676
R1757 B.n501 B.n419 71.676
R1758 B.n497 B.n420 71.676
R1759 B.n493 B.n421 71.676
R1760 B.n489 B.n422 71.676
R1761 B.n485 B.n423 71.676
R1762 B.n481 B.n424 71.676
R1763 B.n477 B.n425 71.676
R1764 B.n473 B.n426 71.676
R1765 B.n469 B.n427 71.676
R1766 B.n465 B.n428 71.676
R1767 B.n461 B.n429 71.676
R1768 B.n457 B.n430 71.676
R1769 B.n453 B.n431 71.676
R1770 B.n449 B.n432 71.676
R1771 B.n445 B.n433 71.676
R1772 B.n441 B.n434 71.676
R1773 B.n916 B.n915 71.676
R1774 B.n916 B.n2 71.676
R1775 B.n137 B.n136 59.5399
R1776 B.n228 B.n134 59.5399
R1777 B.n440 B.n439 59.5399
R1778 B.n535 B.n437 59.5399
R1779 B.n614 B.n390 46.7359
R1780 B.n614 B.n386 46.7359
R1781 B.n620 B.n386 46.7359
R1782 B.n620 B.n381 46.7359
R1783 B.n626 B.n381 46.7359
R1784 B.n626 B.n382 46.7359
R1785 B.n632 B.n374 46.7359
R1786 B.n638 B.n374 46.7359
R1787 B.n638 B.n370 46.7359
R1788 B.n644 B.n370 46.7359
R1789 B.n644 B.n366 46.7359
R1790 B.n650 B.n366 46.7359
R1791 B.n650 B.n362 46.7359
R1792 B.n657 B.n362 46.7359
R1793 B.n657 B.n656 46.7359
R1794 B.n663 B.n355 46.7359
R1795 B.n669 B.n355 46.7359
R1796 B.n669 B.n350 46.7359
R1797 B.n675 B.n350 46.7359
R1798 B.n675 B.n351 46.7359
R1799 B.n681 B.n343 46.7359
R1800 B.n687 B.n343 46.7359
R1801 B.n687 B.n339 46.7359
R1802 B.n693 B.n339 46.7359
R1803 B.n693 B.n335 46.7359
R1804 B.n699 B.n335 46.7359
R1805 B.n705 B.n331 46.7359
R1806 B.n705 B.n327 46.7359
R1807 B.n711 B.n327 46.7359
R1808 B.n711 B.n323 46.7359
R1809 B.n718 B.n323 46.7359
R1810 B.n718 B.n717 46.7359
R1811 B.n724 B.n316 46.7359
R1812 B.n730 B.n316 46.7359
R1813 B.n730 B.n311 46.7359
R1814 B.n736 B.n311 46.7359
R1815 B.n736 B.n312 46.7359
R1816 B.n743 B.n304 46.7359
R1817 B.n749 B.n304 46.7359
R1818 B.n749 B.n4 46.7359
R1819 B.n914 B.n4 46.7359
R1820 B.n914 B.n913 46.7359
R1821 B.n913 B.n912 46.7359
R1822 B.n912 B.n8 46.7359
R1823 B.n12 B.n8 46.7359
R1824 B.n905 B.n12 46.7359
R1825 B.n904 B.n903 46.7359
R1826 B.n903 B.n16 46.7359
R1827 B.n897 B.n16 46.7359
R1828 B.n897 B.n896 46.7359
R1829 B.n896 B.n895 46.7359
R1830 B.n889 B.n26 46.7359
R1831 B.n889 B.n888 46.7359
R1832 B.n888 B.n887 46.7359
R1833 B.n887 B.n30 46.7359
R1834 B.n881 B.n30 46.7359
R1835 B.n881 B.n880 46.7359
R1836 B.n879 B.n37 46.7359
R1837 B.n873 B.n37 46.7359
R1838 B.n873 B.n872 46.7359
R1839 B.n872 B.n871 46.7359
R1840 B.n871 B.n44 46.7359
R1841 B.n865 B.n44 46.7359
R1842 B.n864 B.n863 46.7359
R1843 B.n863 B.n51 46.7359
R1844 B.n857 B.n51 46.7359
R1845 B.n857 B.n856 46.7359
R1846 B.n856 B.n855 46.7359
R1847 B.n849 B.n61 46.7359
R1848 B.n849 B.n848 46.7359
R1849 B.n848 B.n847 46.7359
R1850 B.n847 B.n65 46.7359
R1851 B.n841 B.n65 46.7359
R1852 B.n841 B.n840 46.7359
R1853 B.n840 B.n839 46.7359
R1854 B.n839 B.n72 46.7359
R1855 B.n833 B.n72 46.7359
R1856 B.n832 B.n831 46.7359
R1857 B.n831 B.n79 46.7359
R1858 B.n825 B.n79 46.7359
R1859 B.n825 B.n824 46.7359
R1860 B.n824 B.n823 46.7359
R1861 B.n823 B.n86 46.7359
R1862 B.n351 B.t2 43.9868
R1863 B.n724 B.t9 43.9868
R1864 B.n895 B.t3 43.9868
R1865 B.t4 B.n864 43.9868
R1866 B.n136 B.n135 43.249
R1867 B.n134 B.n133 43.249
R1868 B.n439 B.n438 43.249
R1869 B.n437 B.n436 43.249
R1870 B.n611 B.n610 33.8737
R1871 B.n442 B.n388 33.8737
R1872 B.n814 B.n813 33.8737
R1873 B.n820 B.n819 33.8737
R1874 B.n382 B.t15 28.8665
R1875 B.n663 B.t1 28.8665
R1876 B.n312 B.t7 28.8665
R1877 B.t0 B.n904 28.8665
R1878 B.n855 B.t6 28.8665
R1879 B.t11 B.n832 28.8665
R1880 B.n699 B.t5 23.3682
R1881 B.t5 B.n331 23.3682
R1882 B.n880 B.t8 23.3682
R1883 B.t8 B.n879 23.3682
R1884 B B.n917 18.0485
R1885 B.n632 B.t15 17.8699
R1886 B.n656 B.t1 17.8699
R1887 B.n743 B.t7 17.8699
R1888 B.n905 B.t0 17.8699
R1889 B.n61 B.t6 17.8699
R1890 B.n833 B.t11 17.8699
R1891 B.n612 B.n611 10.6151
R1892 B.n612 B.n384 10.6151
R1893 B.n622 B.n384 10.6151
R1894 B.n623 B.n622 10.6151
R1895 B.n624 B.n623 10.6151
R1896 B.n624 B.n376 10.6151
R1897 B.n634 B.n376 10.6151
R1898 B.n635 B.n634 10.6151
R1899 B.n636 B.n635 10.6151
R1900 B.n636 B.n368 10.6151
R1901 B.n646 B.n368 10.6151
R1902 B.n647 B.n646 10.6151
R1903 B.n648 B.n647 10.6151
R1904 B.n648 B.n360 10.6151
R1905 B.n659 B.n360 10.6151
R1906 B.n660 B.n659 10.6151
R1907 B.n661 B.n660 10.6151
R1908 B.n661 B.n353 10.6151
R1909 B.n671 B.n353 10.6151
R1910 B.n672 B.n671 10.6151
R1911 B.n673 B.n672 10.6151
R1912 B.n673 B.n345 10.6151
R1913 B.n683 B.n345 10.6151
R1914 B.n684 B.n683 10.6151
R1915 B.n685 B.n684 10.6151
R1916 B.n685 B.n337 10.6151
R1917 B.n695 B.n337 10.6151
R1918 B.n696 B.n695 10.6151
R1919 B.n697 B.n696 10.6151
R1920 B.n697 B.n329 10.6151
R1921 B.n707 B.n329 10.6151
R1922 B.n708 B.n707 10.6151
R1923 B.n709 B.n708 10.6151
R1924 B.n709 B.n321 10.6151
R1925 B.n720 B.n321 10.6151
R1926 B.n721 B.n720 10.6151
R1927 B.n722 B.n721 10.6151
R1928 B.n722 B.n314 10.6151
R1929 B.n732 B.n314 10.6151
R1930 B.n733 B.n732 10.6151
R1931 B.n734 B.n733 10.6151
R1932 B.n734 B.n306 10.6151
R1933 B.n745 B.n306 10.6151
R1934 B.n746 B.n745 10.6151
R1935 B.n747 B.n746 10.6151
R1936 B.n747 B.n0 10.6151
R1937 B.n610 B.n392 10.6151
R1938 B.n605 B.n392 10.6151
R1939 B.n605 B.n604 10.6151
R1940 B.n604 B.n603 10.6151
R1941 B.n603 B.n600 10.6151
R1942 B.n600 B.n599 10.6151
R1943 B.n599 B.n596 10.6151
R1944 B.n596 B.n595 10.6151
R1945 B.n595 B.n592 10.6151
R1946 B.n592 B.n591 10.6151
R1947 B.n591 B.n588 10.6151
R1948 B.n588 B.n587 10.6151
R1949 B.n587 B.n584 10.6151
R1950 B.n584 B.n583 10.6151
R1951 B.n583 B.n580 10.6151
R1952 B.n580 B.n579 10.6151
R1953 B.n579 B.n576 10.6151
R1954 B.n576 B.n575 10.6151
R1955 B.n575 B.n572 10.6151
R1956 B.n572 B.n571 10.6151
R1957 B.n571 B.n568 10.6151
R1958 B.n568 B.n567 10.6151
R1959 B.n567 B.n564 10.6151
R1960 B.n564 B.n563 10.6151
R1961 B.n563 B.n560 10.6151
R1962 B.n560 B.n559 10.6151
R1963 B.n559 B.n556 10.6151
R1964 B.n556 B.n555 10.6151
R1965 B.n555 B.n552 10.6151
R1966 B.n552 B.n551 10.6151
R1967 B.n551 B.n548 10.6151
R1968 B.n548 B.n547 10.6151
R1969 B.n547 B.n544 10.6151
R1970 B.n544 B.n543 10.6151
R1971 B.n543 B.n540 10.6151
R1972 B.n540 B.n539 10.6151
R1973 B.n539 B.n536 10.6151
R1974 B.n534 B.n531 10.6151
R1975 B.n531 B.n530 10.6151
R1976 B.n530 B.n527 10.6151
R1977 B.n527 B.n526 10.6151
R1978 B.n526 B.n523 10.6151
R1979 B.n523 B.n522 10.6151
R1980 B.n522 B.n519 10.6151
R1981 B.n519 B.n518 10.6151
R1982 B.n515 B.n514 10.6151
R1983 B.n514 B.n511 10.6151
R1984 B.n511 B.n510 10.6151
R1985 B.n510 B.n507 10.6151
R1986 B.n507 B.n506 10.6151
R1987 B.n506 B.n503 10.6151
R1988 B.n503 B.n502 10.6151
R1989 B.n502 B.n499 10.6151
R1990 B.n499 B.n498 10.6151
R1991 B.n498 B.n495 10.6151
R1992 B.n495 B.n494 10.6151
R1993 B.n494 B.n491 10.6151
R1994 B.n491 B.n490 10.6151
R1995 B.n490 B.n487 10.6151
R1996 B.n487 B.n486 10.6151
R1997 B.n486 B.n483 10.6151
R1998 B.n483 B.n482 10.6151
R1999 B.n482 B.n479 10.6151
R2000 B.n479 B.n478 10.6151
R2001 B.n478 B.n475 10.6151
R2002 B.n475 B.n474 10.6151
R2003 B.n474 B.n471 10.6151
R2004 B.n471 B.n470 10.6151
R2005 B.n470 B.n467 10.6151
R2006 B.n467 B.n466 10.6151
R2007 B.n466 B.n463 10.6151
R2008 B.n463 B.n462 10.6151
R2009 B.n462 B.n459 10.6151
R2010 B.n459 B.n458 10.6151
R2011 B.n458 B.n455 10.6151
R2012 B.n455 B.n454 10.6151
R2013 B.n454 B.n451 10.6151
R2014 B.n451 B.n450 10.6151
R2015 B.n450 B.n447 10.6151
R2016 B.n447 B.n446 10.6151
R2017 B.n446 B.n443 10.6151
R2018 B.n443 B.n442 10.6151
R2019 B.n616 B.n388 10.6151
R2020 B.n617 B.n616 10.6151
R2021 B.n618 B.n617 10.6151
R2022 B.n618 B.n379 10.6151
R2023 B.n628 B.n379 10.6151
R2024 B.n629 B.n628 10.6151
R2025 B.n630 B.n629 10.6151
R2026 B.n630 B.n372 10.6151
R2027 B.n640 B.n372 10.6151
R2028 B.n641 B.n640 10.6151
R2029 B.n642 B.n641 10.6151
R2030 B.n642 B.n364 10.6151
R2031 B.n652 B.n364 10.6151
R2032 B.n653 B.n652 10.6151
R2033 B.n654 B.n653 10.6151
R2034 B.n654 B.n357 10.6151
R2035 B.n665 B.n357 10.6151
R2036 B.n666 B.n665 10.6151
R2037 B.n667 B.n666 10.6151
R2038 B.n667 B.n348 10.6151
R2039 B.n677 B.n348 10.6151
R2040 B.n678 B.n677 10.6151
R2041 B.n679 B.n678 10.6151
R2042 B.n679 B.n341 10.6151
R2043 B.n689 B.n341 10.6151
R2044 B.n690 B.n689 10.6151
R2045 B.n691 B.n690 10.6151
R2046 B.n691 B.n333 10.6151
R2047 B.n701 B.n333 10.6151
R2048 B.n702 B.n701 10.6151
R2049 B.n703 B.n702 10.6151
R2050 B.n703 B.n325 10.6151
R2051 B.n713 B.n325 10.6151
R2052 B.n714 B.n713 10.6151
R2053 B.n715 B.n714 10.6151
R2054 B.n715 B.n318 10.6151
R2055 B.n726 B.n318 10.6151
R2056 B.n727 B.n726 10.6151
R2057 B.n728 B.n727 10.6151
R2058 B.n728 B.n309 10.6151
R2059 B.n738 B.n309 10.6151
R2060 B.n739 B.n738 10.6151
R2061 B.n741 B.n739 10.6151
R2062 B.n741 B.n740 10.6151
R2063 B.n740 B.n302 10.6151
R2064 B.n752 B.n302 10.6151
R2065 B.n753 B.n752 10.6151
R2066 B.n754 B.n753 10.6151
R2067 B.n755 B.n754 10.6151
R2068 B.n756 B.n755 10.6151
R2069 B.n759 B.n756 10.6151
R2070 B.n760 B.n759 10.6151
R2071 B.n761 B.n760 10.6151
R2072 B.n762 B.n761 10.6151
R2073 B.n764 B.n762 10.6151
R2074 B.n765 B.n764 10.6151
R2075 B.n766 B.n765 10.6151
R2076 B.n767 B.n766 10.6151
R2077 B.n769 B.n767 10.6151
R2078 B.n770 B.n769 10.6151
R2079 B.n771 B.n770 10.6151
R2080 B.n772 B.n771 10.6151
R2081 B.n774 B.n772 10.6151
R2082 B.n775 B.n774 10.6151
R2083 B.n776 B.n775 10.6151
R2084 B.n777 B.n776 10.6151
R2085 B.n779 B.n777 10.6151
R2086 B.n780 B.n779 10.6151
R2087 B.n781 B.n780 10.6151
R2088 B.n782 B.n781 10.6151
R2089 B.n784 B.n782 10.6151
R2090 B.n785 B.n784 10.6151
R2091 B.n786 B.n785 10.6151
R2092 B.n787 B.n786 10.6151
R2093 B.n789 B.n787 10.6151
R2094 B.n790 B.n789 10.6151
R2095 B.n791 B.n790 10.6151
R2096 B.n792 B.n791 10.6151
R2097 B.n794 B.n792 10.6151
R2098 B.n795 B.n794 10.6151
R2099 B.n796 B.n795 10.6151
R2100 B.n797 B.n796 10.6151
R2101 B.n799 B.n797 10.6151
R2102 B.n800 B.n799 10.6151
R2103 B.n801 B.n800 10.6151
R2104 B.n802 B.n801 10.6151
R2105 B.n804 B.n802 10.6151
R2106 B.n805 B.n804 10.6151
R2107 B.n806 B.n805 10.6151
R2108 B.n807 B.n806 10.6151
R2109 B.n809 B.n807 10.6151
R2110 B.n810 B.n809 10.6151
R2111 B.n811 B.n810 10.6151
R2112 B.n812 B.n811 10.6151
R2113 B.n813 B.n812 10.6151
R2114 B.n909 B.n1 10.6151
R2115 B.n909 B.n908 10.6151
R2116 B.n908 B.n907 10.6151
R2117 B.n907 B.n10 10.6151
R2118 B.n901 B.n10 10.6151
R2119 B.n901 B.n900 10.6151
R2120 B.n900 B.n899 10.6151
R2121 B.n899 B.n18 10.6151
R2122 B.n893 B.n18 10.6151
R2123 B.n893 B.n892 10.6151
R2124 B.n892 B.n891 10.6151
R2125 B.n891 B.n24 10.6151
R2126 B.n885 B.n24 10.6151
R2127 B.n885 B.n884 10.6151
R2128 B.n884 B.n883 10.6151
R2129 B.n883 B.n32 10.6151
R2130 B.n877 B.n32 10.6151
R2131 B.n877 B.n876 10.6151
R2132 B.n876 B.n875 10.6151
R2133 B.n875 B.n39 10.6151
R2134 B.n869 B.n39 10.6151
R2135 B.n869 B.n868 10.6151
R2136 B.n868 B.n867 10.6151
R2137 B.n867 B.n46 10.6151
R2138 B.n861 B.n46 10.6151
R2139 B.n861 B.n860 10.6151
R2140 B.n860 B.n859 10.6151
R2141 B.n859 B.n53 10.6151
R2142 B.n853 B.n53 10.6151
R2143 B.n853 B.n852 10.6151
R2144 B.n852 B.n851 10.6151
R2145 B.n851 B.n59 10.6151
R2146 B.n845 B.n59 10.6151
R2147 B.n845 B.n844 10.6151
R2148 B.n844 B.n843 10.6151
R2149 B.n843 B.n67 10.6151
R2150 B.n837 B.n67 10.6151
R2151 B.n837 B.n836 10.6151
R2152 B.n836 B.n835 10.6151
R2153 B.n835 B.n74 10.6151
R2154 B.n829 B.n74 10.6151
R2155 B.n829 B.n828 10.6151
R2156 B.n828 B.n827 10.6151
R2157 B.n827 B.n81 10.6151
R2158 B.n821 B.n81 10.6151
R2159 B.n821 B.n820 10.6151
R2160 B.n819 B.n88 10.6151
R2161 B.n139 B.n88 10.6151
R2162 B.n140 B.n139 10.6151
R2163 B.n143 B.n140 10.6151
R2164 B.n144 B.n143 10.6151
R2165 B.n147 B.n144 10.6151
R2166 B.n148 B.n147 10.6151
R2167 B.n151 B.n148 10.6151
R2168 B.n152 B.n151 10.6151
R2169 B.n155 B.n152 10.6151
R2170 B.n156 B.n155 10.6151
R2171 B.n159 B.n156 10.6151
R2172 B.n160 B.n159 10.6151
R2173 B.n163 B.n160 10.6151
R2174 B.n164 B.n163 10.6151
R2175 B.n167 B.n164 10.6151
R2176 B.n168 B.n167 10.6151
R2177 B.n171 B.n168 10.6151
R2178 B.n172 B.n171 10.6151
R2179 B.n175 B.n172 10.6151
R2180 B.n176 B.n175 10.6151
R2181 B.n179 B.n176 10.6151
R2182 B.n180 B.n179 10.6151
R2183 B.n183 B.n180 10.6151
R2184 B.n184 B.n183 10.6151
R2185 B.n187 B.n184 10.6151
R2186 B.n188 B.n187 10.6151
R2187 B.n191 B.n188 10.6151
R2188 B.n192 B.n191 10.6151
R2189 B.n195 B.n192 10.6151
R2190 B.n196 B.n195 10.6151
R2191 B.n199 B.n196 10.6151
R2192 B.n200 B.n199 10.6151
R2193 B.n203 B.n200 10.6151
R2194 B.n204 B.n203 10.6151
R2195 B.n207 B.n204 10.6151
R2196 B.n208 B.n207 10.6151
R2197 B.n212 B.n211 10.6151
R2198 B.n215 B.n212 10.6151
R2199 B.n216 B.n215 10.6151
R2200 B.n219 B.n216 10.6151
R2201 B.n220 B.n219 10.6151
R2202 B.n223 B.n220 10.6151
R2203 B.n224 B.n223 10.6151
R2204 B.n227 B.n224 10.6151
R2205 B.n232 B.n229 10.6151
R2206 B.n233 B.n232 10.6151
R2207 B.n236 B.n233 10.6151
R2208 B.n237 B.n236 10.6151
R2209 B.n240 B.n237 10.6151
R2210 B.n241 B.n240 10.6151
R2211 B.n244 B.n241 10.6151
R2212 B.n245 B.n244 10.6151
R2213 B.n248 B.n245 10.6151
R2214 B.n249 B.n248 10.6151
R2215 B.n252 B.n249 10.6151
R2216 B.n253 B.n252 10.6151
R2217 B.n256 B.n253 10.6151
R2218 B.n257 B.n256 10.6151
R2219 B.n260 B.n257 10.6151
R2220 B.n261 B.n260 10.6151
R2221 B.n264 B.n261 10.6151
R2222 B.n265 B.n264 10.6151
R2223 B.n268 B.n265 10.6151
R2224 B.n269 B.n268 10.6151
R2225 B.n272 B.n269 10.6151
R2226 B.n273 B.n272 10.6151
R2227 B.n276 B.n273 10.6151
R2228 B.n277 B.n276 10.6151
R2229 B.n280 B.n277 10.6151
R2230 B.n281 B.n280 10.6151
R2231 B.n284 B.n281 10.6151
R2232 B.n285 B.n284 10.6151
R2233 B.n288 B.n285 10.6151
R2234 B.n289 B.n288 10.6151
R2235 B.n292 B.n289 10.6151
R2236 B.n293 B.n292 10.6151
R2237 B.n296 B.n293 10.6151
R2238 B.n297 B.n296 10.6151
R2239 B.n300 B.n297 10.6151
R2240 B.n301 B.n300 10.6151
R2241 B.n814 B.n301 10.6151
R2242 B.n917 B.n0 8.11757
R2243 B.n917 B.n1 8.11757
R2244 B.n535 B.n534 6.5566
R2245 B.n518 B.n440 6.5566
R2246 B.n211 B.n137 6.5566
R2247 B.n228 B.n227 6.5566
R2248 B.n536 B.n535 4.05904
R2249 B.n515 B.n440 4.05904
R2250 B.n208 B.n137 4.05904
R2251 B.n229 B.n228 4.05904
R2252 B.n681 B.t2 2.74964
R2253 B.n717 B.t9 2.74964
R2254 B.n26 B.t3 2.74964
R2255 B.n865 B.t4 2.74964
R2256 VP.n16 VP.t8 166.995
R2257 VP.n18 VP.n15 161.3
R2258 VP.n20 VP.n19 161.3
R2259 VP.n21 VP.n14 161.3
R2260 VP.n23 VP.n22 161.3
R2261 VP.n24 VP.n13 161.3
R2262 VP.n26 VP.n25 161.3
R2263 VP.n27 VP.n12 161.3
R2264 VP.n29 VP.n28 161.3
R2265 VP.n30 VP.n11 161.3
R2266 VP.n33 VP.n32 161.3
R2267 VP.n34 VP.n10 161.3
R2268 VP.n36 VP.n35 161.3
R2269 VP.n37 VP.n9 161.3
R2270 VP.n68 VP.n0 161.3
R2271 VP.n67 VP.n66 161.3
R2272 VP.n65 VP.n1 161.3
R2273 VP.n64 VP.n63 161.3
R2274 VP.n61 VP.n2 161.3
R2275 VP.n60 VP.n59 161.3
R2276 VP.n58 VP.n3 161.3
R2277 VP.n57 VP.n56 161.3
R2278 VP.n55 VP.n4 161.3
R2279 VP.n54 VP.n53 161.3
R2280 VP.n52 VP.n5 161.3
R2281 VP.n51 VP.n50 161.3
R2282 VP.n49 VP.n6 161.3
R2283 VP.n47 VP.n46 161.3
R2284 VP.n45 VP.n7 161.3
R2285 VP.n44 VP.n43 161.3
R2286 VP.n42 VP.n8 161.3
R2287 VP.n55 VP.t1 136.102
R2288 VP.n41 VP.t0 136.102
R2289 VP.n48 VP.t9 136.102
R2290 VP.n62 VP.t4 136.102
R2291 VP.n69 VP.t7 136.102
R2292 VP.n24 VP.t5 136.102
R2293 VP.n38 VP.t2 136.102
R2294 VP.n31 VP.t3 136.102
R2295 VP.n17 VP.t6 136.102
R2296 VP.n41 VP.n40 88.2468
R2297 VP.n70 VP.n69 88.2468
R2298 VP.n39 VP.n38 88.2468
R2299 VP.n17 VP.n16 58.8387
R2300 VP.n43 VP.n7 55.548
R2301 VP.n67 VP.n1 55.548
R2302 VP.n36 VP.n10 55.548
R2303 VP.n50 VP.n5 51.663
R2304 VP.n60 VP.n3 51.663
R2305 VP.n29 VP.n12 51.663
R2306 VP.n19 VP.n14 51.663
R2307 VP.n40 VP.n39 48.3897
R2308 VP.n54 VP.n5 29.3238
R2309 VP.n56 VP.n3 29.3238
R2310 VP.n25 VP.n12 29.3238
R2311 VP.n23 VP.n14 29.3238
R2312 VP.n43 VP.n42 25.4388
R2313 VP.n68 VP.n67 25.4388
R2314 VP.n37 VP.n36 25.4388
R2315 VP.n47 VP.n7 24.4675
R2316 VP.n50 VP.n49 24.4675
R2317 VP.n55 VP.n54 24.4675
R2318 VP.n56 VP.n55 24.4675
R2319 VP.n61 VP.n60 24.4675
R2320 VP.n63 VP.n1 24.4675
R2321 VP.n30 VP.n29 24.4675
R2322 VP.n32 VP.n10 24.4675
R2323 VP.n24 VP.n23 24.4675
R2324 VP.n25 VP.n24 24.4675
R2325 VP.n19 VP.n18 24.4675
R2326 VP.n42 VP.n41 22.5101
R2327 VP.n69 VP.n68 22.5101
R2328 VP.n38 VP.n37 22.5101
R2329 VP.n48 VP.n47 13.2127
R2330 VP.n63 VP.n62 13.2127
R2331 VP.n32 VP.n31 13.2127
R2332 VP.n16 VP.n15 12.9374
R2333 VP.n49 VP.n48 11.2553
R2334 VP.n62 VP.n61 11.2553
R2335 VP.n31 VP.n30 11.2553
R2336 VP.n18 VP.n17 11.2553
R2337 VP.n39 VP.n9 0.278367
R2338 VP.n40 VP.n8 0.278367
R2339 VP.n70 VP.n0 0.278367
R2340 VP.n20 VP.n15 0.189894
R2341 VP.n21 VP.n20 0.189894
R2342 VP.n22 VP.n21 0.189894
R2343 VP.n22 VP.n13 0.189894
R2344 VP.n26 VP.n13 0.189894
R2345 VP.n27 VP.n26 0.189894
R2346 VP.n28 VP.n27 0.189894
R2347 VP.n28 VP.n11 0.189894
R2348 VP.n33 VP.n11 0.189894
R2349 VP.n34 VP.n33 0.189894
R2350 VP.n35 VP.n34 0.189894
R2351 VP.n35 VP.n9 0.189894
R2352 VP.n44 VP.n8 0.189894
R2353 VP.n45 VP.n44 0.189894
R2354 VP.n46 VP.n45 0.189894
R2355 VP.n46 VP.n6 0.189894
R2356 VP.n51 VP.n6 0.189894
R2357 VP.n52 VP.n51 0.189894
R2358 VP.n53 VP.n52 0.189894
R2359 VP.n53 VP.n4 0.189894
R2360 VP.n57 VP.n4 0.189894
R2361 VP.n58 VP.n57 0.189894
R2362 VP.n59 VP.n58 0.189894
R2363 VP.n59 VP.n2 0.189894
R2364 VP.n64 VP.n2 0.189894
R2365 VP.n65 VP.n64 0.189894
R2366 VP.n66 VP.n65 0.189894
R2367 VP.n66 VP.n0 0.189894
R2368 VP VP.n70 0.153454
R2369 VDD1.n52 VDD1.n0 289.615
R2370 VDD1.n111 VDD1.n59 289.615
R2371 VDD1.n53 VDD1.n52 185
R2372 VDD1.n51 VDD1.n50 185
R2373 VDD1.n4 VDD1.n3 185
R2374 VDD1.n45 VDD1.n44 185
R2375 VDD1.n43 VDD1.n42 185
R2376 VDD1.n41 VDD1.n7 185
R2377 VDD1.n11 VDD1.n8 185
R2378 VDD1.n36 VDD1.n35 185
R2379 VDD1.n34 VDD1.n33 185
R2380 VDD1.n13 VDD1.n12 185
R2381 VDD1.n28 VDD1.n27 185
R2382 VDD1.n26 VDD1.n25 185
R2383 VDD1.n17 VDD1.n16 185
R2384 VDD1.n20 VDD1.n19 185
R2385 VDD1.n78 VDD1.n77 185
R2386 VDD1.n75 VDD1.n74 185
R2387 VDD1.n84 VDD1.n83 185
R2388 VDD1.n86 VDD1.n85 185
R2389 VDD1.n71 VDD1.n70 185
R2390 VDD1.n92 VDD1.n91 185
R2391 VDD1.n95 VDD1.n94 185
R2392 VDD1.n93 VDD1.n67 185
R2393 VDD1.n100 VDD1.n66 185
R2394 VDD1.n102 VDD1.n101 185
R2395 VDD1.n104 VDD1.n103 185
R2396 VDD1.n63 VDD1.n62 185
R2397 VDD1.n110 VDD1.n109 185
R2398 VDD1.n112 VDD1.n111 185
R2399 VDD1.t1 VDD1.n18 149.524
R2400 VDD1.t9 VDD1.n76 149.524
R2401 VDD1.n52 VDD1.n51 104.615
R2402 VDD1.n51 VDD1.n3 104.615
R2403 VDD1.n44 VDD1.n3 104.615
R2404 VDD1.n44 VDD1.n43 104.615
R2405 VDD1.n43 VDD1.n7 104.615
R2406 VDD1.n11 VDD1.n7 104.615
R2407 VDD1.n35 VDD1.n11 104.615
R2408 VDD1.n35 VDD1.n34 104.615
R2409 VDD1.n34 VDD1.n12 104.615
R2410 VDD1.n27 VDD1.n12 104.615
R2411 VDD1.n27 VDD1.n26 104.615
R2412 VDD1.n26 VDD1.n16 104.615
R2413 VDD1.n19 VDD1.n16 104.615
R2414 VDD1.n77 VDD1.n74 104.615
R2415 VDD1.n84 VDD1.n74 104.615
R2416 VDD1.n85 VDD1.n84 104.615
R2417 VDD1.n85 VDD1.n70 104.615
R2418 VDD1.n92 VDD1.n70 104.615
R2419 VDD1.n94 VDD1.n92 104.615
R2420 VDD1.n94 VDD1.n93 104.615
R2421 VDD1.n93 VDD1.n66 104.615
R2422 VDD1.n102 VDD1.n66 104.615
R2423 VDD1.n103 VDD1.n102 104.615
R2424 VDD1.n103 VDD1.n62 104.615
R2425 VDD1.n110 VDD1.n62 104.615
R2426 VDD1.n111 VDD1.n110 104.615
R2427 VDD1.n119 VDD1.n118 64.6963
R2428 VDD1.n58 VDD1.n57 63.31
R2429 VDD1.n121 VDD1.n120 63.3098
R2430 VDD1.n117 VDD1.n116 63.3098
R2431 VDD1.n19 VDD1.t1 52.3082
R2432 VDD1.n77 VDD1.t9 52.3082
R2433 VDD1.n58 VDD1.n56 51.7562
R2434 VDD1.n117 VDD1.n115 51.7562
R2435 VDD1.n121 VDD1.n119 43.641
R2436 VDD1.n42 VDD1.n41 13.1884
R2437 VDD1.n101 VDD1.n100 13.1884
R2438 VDD1.n45 VDD1.n6 12.8005
R2439 VDD1.n40 VDD1.n8 12.8005
R2440 VDD1.n99 VDD1.n67 12.8005
R2441 VDD1.n104 VDD1.n65 12.8005
R2442 VDD1.n46 VDD1.n4 12.0247
R2443 VDD1.n37 VDD1.n36 12.0247
R2444 VDD1.n96 VDD1.n95 12.0247
R2445 VDD1.n105 VDD1.n63 12.0247
R2446 VDD1.n50 VDD1.n49 11.249
R2447 VDD1.n33 VDD1.n10 11.249
R2448 VDD1.n91 VDD1.n69 11.249
R2449 VDD1.n109 VDD1.n108 11.249
R2450 VDD1.n53 VDD1.n2 10.4732
R2451 VDD1.n32 VDD1.n13 10.4732
R2452 VDD1.n90 VDD1.n71 10.4732
R2453 VDD1.n112 VDD1.n61 10.4732
R2454 VDD1.n20 VDD1.n18 10.2747
R2455 VDD1.n78 VDD1.n76 10.2747
R2456 VDD1.n54 VDD1.n0 9.69747
R2457 VDD1.n29 VDD1.n28 9.69747
R2458 VDD1.n87 VDD1.n86 9.69747
R2459 VDD1.n113 VDD1.n59 9.69747
R2460 VDD1.n56 VDD1.n55 9.45567
R2461 VDD1.n115 VDD1.n114 9.45567
R2462 VDD1.n22 VDD1.n21 9.3005
R2463 VDD1.n24 VDD1.n23 9.3005
R2464 VDD1.n15 VDD1.n14 9.3005
R2465 VDD1.n30 VDD1.n29 9.3005
R2466 VDD1.n32 VDD1.n31 9.3005
R2467 VDD1.n10 VDD1.n9 9.3005
R2468 VDD1.n38 VDD1.n37 9.3005
R2469 VDD1.n40 VDD1.n39 9.3005
R2470 VDD1.n55 VDD1.n54 9.3005
R2471 VDD1.n2 VDD1.n1 9.3005
R2472 VDD1.n49 VDD1.n48 9.3005
R2473 VDD1.n47 VDD1.n46 9.3005
R2474 VDD1.n6 VDD1.n5 9.3005
R2475 VDD1.n114 VDD1.n113 9.3005
R2476 VDD1.n61 VDD1.n60 9.3005
R2477 VDD1.n108 VDD1.n107 9.3005
R2478 VDD1.n106 VDD1.n105 9.3005
R2479 VDD1.n65 VDD1.n64 9.3005
R2480 VDD1.n80 VDD1.n79 9.3005
R2481 VDD1.n82 VDD1.n81 9.3005
R2482 VDD1.n73 VDD1.n72 9.3005
R2483 VDD1.n88 VDD1.n87 9.3005
R2484 VDD1.n90 VDD1.n89 9.3005
R2485 VDD1.n69 VDD1.n68 9.3005
R2486 VDD1.n97 VDD1.n96 9.3005
R2487 VDD1.n99 VDD1.n98 9.3005
R2488 VDD1.n25 VDD1.n15 8.92171
R2489 VDD1.n83 VDD1.n73 8.92171
R2490 VDD1.n24 VDD1.n17 8.14595
R2491 VDD1.n82 VDD1.n75 8.14595
R2492 VDD1.n21 VDD1.n20 7.3702
R2493 VDD1.n79 VDD1.n78 7.3702
R2494 VDD1.n21 VDD1.n17 5.81868
R2495 VDD1.n79 VDD1.n75 5.81868
R2496 VDD1.n25 VDD1.n24 5.04292
R2497 VDD1.n83 VDD1.n82 5.04292
R2498 VDD1.n56 VDD1.n0 4.26717
R2499 VDD1.n28 VDD1.n15 4.26717
R2500 VDD1.n86 VDD1.n73 4.26717
R2501 VDD1.n115 VDD1.n59 4.26717
R2502 VDD1.n54 VDD1.n53 3.49141
R2503 VDD1.n29 VDD1.n13 3.49141
R2504 VDD1.n87 VDD1.n71 3.49141
R2505 VDD1.n113 VDD1.n112 3.49141
R2506 VDD1.n22 VDD1.n18 2.84303
R2507 VDD1.n80 VDD1.n76 2.84303
R2508 VDD1.n50 VDD1.n2 2.71565
R2509 VDD1.n33 VDD1.n32 2.71565
R2510 VDD1.n91 VDD1.n90 2.71565
R2511 VDD1.n109 VDD1.n61 2.71565
R2512 VDD1.n49 VDD1.n4 1.93989
R2513 VDD1.n36 VDD1.n10 1.93989
R2514 VDD1.n95 VDD1.n69 1.93989
R2515 VDD1.n108 VDD1.n63 1.93989
R2516 VDD1.n120 VDD1.t6 1.84579
R2517 VDD1.n120 VDD1.t7 1.84579
R2518 VDD1.n57 VDD1.t3 1.84579
R2519 VDD1.n57 VDD1.t4 1.84579
R2520 VDD1.n118 VDD1.t5 1.84579
R2521 VDD1.n118 VDD1.t2 1.84579
R2522 VDD1.n116 VDD1.t0 1.84579
R2523 VDD1.n116 VDD1.t8 1.84579
R2524 VDD1 VDD1.n121 1.38412
R2525 VDD1.n46 VDD1.n45 1.16414
R2526 VDD1.n37 VDD1.n8 1.16414
R2527 VDD1.n96 VDD1.n67 1.16414
R2528 VDD1.n105 VDD1.n104 1.16414
R2529 VDD1 VDD1.n58 0.539293
R2530 VDD1.n119 VDD1.n117 0.425757
R2531 VDD1.n42 VDD1.n6 0.388379
R2532 VDD1.n41 VDD1.n40 0.388379
R2533 VDD1.n100 VDD1.n99 0.388379
R2534 VDD1.n101 VDD1.n65 0.388379
R2535 VDD1.n55 VDD1.n1 0.155672
R2536 VDD1.n48 VDD1.n1 0.155672
R2537 VDD1.n48 VDD1.n47 0.155672
R2538 VDD1.n47 VDD1.n5 0.155672
R2539 VDD1.n39 VDD1.n5 0.155672
R2540 VDD1.n39 VDD1.n38 0.155672
R2541 VDD1.n38 VDD1.n9 0.155672
R2542 VDD1.n31 VDD1.n9 0.155672
R2543 VDD1.n31 VDD1.n30 0.155672
R2544 VDD1.n30 VDD1.n14 0.155672
R2545 VDD1.n23 VDD1.n14 0.155672
R2546 VDD1.n23 VDD1.n22 0.155672
R2547 VDD1.n81 VDD1.n80 0.155672
R2548 VDD1.n81 VDD1.n72 0.155672
R2549 VDD1.n88 VDD1.n72 0.155672
R2550 VDD1.n89 VDD1.n88 0.155672
R2551 VDD1.n89 VDD1.n68 0.155672
R2552 VDD1.n97 VDD1.n68 0.155672
R2553 VDD1.n98 VDD1.n97 0.155672
R2554 VDD1.n98 VDD1.n64 0.155672
R2555 VDD1.n106 VDD1.n64 0.155672
R2556 VDD1.n107 VDD1.n106 0.155672
R2557 VDD1.n107 VDD1.n60 0.155672
R2558 VDD1.n114 VDD1.n60 0.155672
C0 VTAIL VDD2 9.85583f
C1 VN VDD1 0.151783f
C2 VTAIL VDD1 9.810121f
C3 VN VTAIL 9.32655f
C4 VP VDD2 0.494228f
C5 VP VDD1 9.26017f
C6 VP VN 7.13278f
C7 VP VTAIL 9.34089f
C8 VDD1 VDD2 1.71903f
C9 VN VDD2 8.92139f
C10 VDD2 B 6.146704f
C11 VDD1 B 6.132433f
C12 VTAIL B 7.158423f
C13 VN B 14.74304f
C14 VP B 13.214104f
C15 VDD1.n0 B 0.031262f
C16 VDD1.n1 B 0.022566f
C17 VDD1.n2 B 0.012126f
C18 VDD1.n3 B 0.028661f
C19 VDD1.n4 B 0.012839f
C20 VDD1.n5 B 0.022566f
C21 VDD1.n6 B 0.012126f
C22 VDD1.n7 B 0.028661f
C23 VDD1.n8 B 0.012839f
C24 VDD1.n9 B 0.022566f
C25 VDD1.n10 B 0.012126f
C26 VDD1.n11 B 0.028661f
C27 VDD1.n12 B 0.028661f
C28 VDD1.n13 B 0.012839f
C29 VDD1.n14 B 0.022566f
C30 VDD1.n15 B 0.012126f
C31 VDD1.n16 B 0.028661f
C32 VDD1.n17 B 0.012839f
C33 VDD1.n18 B 0.151696f
C34 VDD1.t1 B 0.048254f
C35 VDD1.n19 B 0.021496f
C36 VDD1.n20 B 0.020261f
C37 VDD1.n21 B 0.012126f
C38 VDD1.n22 B 1.01094f
C39 VDD1.n23 B 0.022566f
C40 VDD1.n24 B 0.012126f
C41 VDD1.n25 B 0.012839f
C42 VDD1.n26 B 0.028661f
C43 VDD1.n27 B 0.028661f
C44 VDD1.n28 B 0.012839f
C45 VDD1.n29 B 0.012126f
C46 VDD1.n30 B 0.022566f
C47 VDD1.n31 B 0.022566f
C48 VDD1.n32 B 0.012126f
C49 VDD1.n33 B 0.012839f
C50 VDD1.n34 B 0.028661f
C51 VDD1.n35 B 0.028661f
C52 VDD1.n36 B 0.012839f
C53 VDD1.n37 B 0.012126f
C54 VDD1.n38 B 0.022566f
C55 VDD1.n39 B 0.022566f
C56 VDD1.n40 B 0.012126f
C57 VDD1.n41 B 0.012483f
C58 VDD1.n42 B 0.012483f
C59 VDD1.n43 B 0.028661f
C60 VDD1.n44 B 0.028661f
C61 VDD1.n45 B 0.012839f
C62 VDD1.n46 B 0.012126f
C63 VDD1.n47 B 0.022566f
C64 VDD1.n48 B 0.022566f
C65 VDD1.n49 B 0.012126f
C66 VDD1.n50 B 0.012839f
C67 VDD1.n51 B 0.028661f
C68 VDD1.n52 B 0.061239f
C69 VDD1.n53 B 0.012839f
C70 VDD1.n54 B 0.012126f
C71 VDD1.n55 B 0.053701f
C72 VDD1.n56 B 0.056638f
C73 VDD1.t3 B 0.19134f
C74 VDD1.t4 B 0.19134f
C75 VDD1.n57 B 1.69369f
C76 VDD1.n58 B 0.540603f
C77 VDD1.n59 B 0.031262f
C78 VDD1.n60 B 0.022566f
C79 VDD1.n61 B 0.012126f
C80 VDD1.n62 B 0.028661f
C81 VDD1.n63 B 0.012839f
C82 VDD1.n64 B 0.022566f
C83 VDD1.n65 B 0.012126f
C84 VDD1.n66 B 0.028661f
C85 VDD1.n67 B 0.012839f
C86 VDD1.n68 B 0.022566f
C87 VDD1.n69 B 0.012126f
C88 VDD1.n70 B 0.028661f
C89 VDD1.n71 B 0.012839f
C90 VDD1.n72 B 0.022566f
C91 VDD1.n73 B 0.012126f
C92 VDD1.n74 B 0.028661f
C93 VDD1.n75 B 0.012839f
C94 VDD1.n76 B 0.151696f
C95 VDD1.t9 B 0.048254f
C96 VDD1.n77 B 0.021496f
C97 VDD1.n78 B 0.020261f
C98 VDD1.n79 B 0.012126f
C99 VDD1.n80 B 1.01094f
C100 VDD1.n81 B 0.022566f
C101 VDD1.n82 B 0.012126f
C102 VDD1.n83 B 0.012839f
C103 VDD1.n84 B 0.028661f
C104 VDD1.n85 B 0.028661f
C105 VDD1.n86 B 0.012839f
C106 VDD1.n87 B 0.012126f
C107 VDD1.n88 B 0.022566f
C108 VDD1.n89 B 0.022566f
C109 VDD1.n90 B 0.012126f
C110 VDD1.n91 B 0.012839f
C111 VDD1.n92 B 0.028661f
C112 VDD1.n93 B 0.028661f
C113 VDD1.n94 B 0.028661f
C114 VDD1.n95 B 0.012839f
C115 VDD1.n96 B 0.012126f
C116 VDD1.n97 B 0.022566f
C117 VDD1.n98 B 0.022566f
C118 VDD1.n99 B 0.012126f
C119 VDD1.n100 B 0.012483f
C120 VDD1.n101 B 0.012483f
C121 VDD1.n102 B 0.028661f
C122 VDD1.n103 B 0.028661f
C123 VDD1.n104 B 0.012839f
C124 VDD1.n105 B 0.012126f
C125 VDD1.n106 B 0.022566f
C126 VDD1.n107 B 0.022566f
C127 VDD1.n108 B 0.012126f
C128 VDD1.n109 B 0.012839f
C129 VDD1.n110 B 0.028661f
C130 VDD1.n111 B 0.061239f
C131 VDD1.n112 B 0.012839f
C132 VDD1.n113 B 0.012126f
C133 VDD1.n114 B 0.053701f
C134 VDD1.n115 B 0.056638f
C135 VDD1.t0 B 0.19134f
C136 VDD1.t8 B 0.19134f
C137 VDD1.n116 B 1.69368f
C138 VDD1.n117 B 0.533585f
C139 VDD1.t5 B 0.19134f
C140 VDD1.t2 B 0.19134f
C141 VDD1.n118 B 1.70299f
C142 VDD1.n119 B 2.31552f
C143 VDD1.t6 B 0.19134f
C144 VDD1.t7 B 0.19134f
C145 VDD1.n120 B 1.69368f
C146 VDD1.n121 B 2.5128f
C147 VP.n0 B 0.035216f
C148 VP.t7 B 1.47869f
C149 VP.n1 B 0.045932f
C150 VP.n2 B 0.026711f
C151 VP.t4 B 1.47869f
C152 VP.n3 B 0.026505f
C153 VP.n4 B 0.026711f
C154 VP.t1 B 1.47869f
C155 VP.n5 B 0.026505f
C156 VP.n6 B 0.026711f
C157 VP.t9 B 1.47869f
C158 VP.n7 B 0.045932f
C159 VP.n8 B 0.035216f
C160 VP.t0 B 1.47869f
C161 VP.n9 B 0.035216f
C162 VP.t2 B 1.47869f
C163 VP.n10 B 0.045932f
C164 VP.n11 B 0.026711f
C165 VP.t3 B 1.47869f
C166 VP.n12 B 0.026505f
C167 VP.n13 B 0.026711f
C168 VP.t5 B 1.47869f
C169 VP.n14 B 0.026505f
C170 VP.n15 B 0.197578f
C171 VP.t6 B 1.47869f
C172 VP.t8 B 1.60104f
C173 VP.n16 B 0.601772f
C174 VP.n17 B 0.594078f
C175 VP.n18 B 0.036511f
C176 VP.n19 B 0.04823f
C177 VP.n20 B 0.026711f
C178 VP.n21 B 0.026711f
C179 VP.n22 B 0.026711f
C180 VP.n23 B 0.053039f
C181 VP.n24 B 0.558484f
C182 VP.n25 B 0.053039f
C183 VP.n26 B 0.026711f
C184 VP.n27 B 0.026711f
C185 VP.n28 B 0.026711f
C186 VP.n29 B 0.04823f
C187 VP.n30 B 0.036511f
C188 VP.n31 B 0.533279f
C189 VP.n32 B 0.038477f
C190 VP.n33 B 0.026711f
C191 VP.n34 B 0.026711f
C192 VP.n35 B 0.026711f
C193 VP.n36 B 0.031159f
C194 VP.n37 B 0.048717f
C195 VP.n38 B 0.61547f
C196 VP.n39 B 1.40171f
C197 VP.n40 B 1.42155f
C198 VP.n41 B 0.61547f
C199 VP.n42 B 0.048717f
C200 VP.n43 B 0.031159f
C201 VP.n44 B 0.026711f
C202 VP.n45 B 0.026711f
C203 VP.n46 B 0.026711f
C204 VP.n47 B 0.038477f
C205 VP.n48 B 0.533279f
C206 VP.n49 B 0.036511f
C207 VP.n50 B 0.04823f
C208 VP.n51 B 0.026711f
C209 VP.n52 B 0.026711f
C210 VP.n53 B 0.026711f
C211 VP.n54 B 0.053039f
C212 VP.n55 B 0.558484f
C213 VP.n56 B 0.053039f
C214 VP.n57 B 0.026711f
C215 VP.n58 B 0.026711f
C216 VP.n59 B 0.026711f
C217 VP.n60 B 0.04823f
C218 VP.n61 B 0.036511f
C219 VP.n62 B 0.533279f
C220 VP.n63 B 0.038477f
C221 VP.n64 B 0.026711f
C222 VP.n65 B 0.026711f
C223 VP.n66 B 0.026711f
C224 VP.n67 B 0.031159f
C225 VP.n68 B 0.048717f
C226 VP.n69 B 0.61547f
C227 VP.n70 B 0.029876f
C228 VDD2.n0 B 0.030906f
C229 VDD2.n1 B 0.022309f
C230 VDD2.n2 B 0.011988f
C231 VDD2.n3 B 0.028335f
C232 VDD2.n4 B 0.012693f
C233 VDD2.n5 B 0.022309f
C234 VDD2.n6 B 0.011988f
C235 VDD2.n7 B 0.028335f
C236 VDD2.n8 B 0.012693f
C237 VDD2.n9 B 0.022309f
C238 VDD2.n10 B 0.011988f
C239 VDD2.n11 B 0.028335f
C240 VDD2.n12 B 0.012693f
C241 VDD2.n13 B 0.022309f
C242 VDD2.n14 B 0.011988f
C243 VDD2.n15 B 0.028335f
C244 VDD2.n16 B 0.012693f
C245 VDD2.n17 B 0.149968f
C246 VDD2.t9 B 0.047704f
C247 VDD2.n18 B 0.021251f
C248 VDD2.n19 B 0.020031f
C249 VDD2.n20 B 0.011988f
C250 VDD2.n21 B 0.999421f
C251 VDD2.n22 B 0.022309f
C252 VDD2.n23 B 0.011988f
C253 VDD2.n24 B 0.012693f
C254 VDD2.n25 B 0.028335f
C255 VDD2.n26 B 0.028335f
C256 VDD2.n27 B 0.012693f
C257 VDD2.n28 B 0.011988f
C258 VDD2.n29 B 0.022309f
C259 VDD2.n30 B 0.022309f
C260 VDD2.n31 B 0.011988f
C261 VDD2.n32 B 0.012693f
C262 VDD2.n33 B 0.028335f
C263 VDD2.n34 B 0.028335f
C264 VDD2.n35 B 0.028335f
C265 VDD2.n36 B 0.012693f
C266 VDD2.n37 B 0.011988f
C267 VDD2.n38 B 0.022309f
C268 VDD2.n39 B 0.022309f
C269 VDD2.n40 B 0.011988f
C270 VDD2.n41 B 0.01234f
C271 VDD2.n42 B 0.01234f
C272 VDD2.n43 B 0.028335f
C273 VDD2.n44 B 0.028335f
C274 VDD2.n45 B 0.012693f
C275 VDD2.n46 B 0.011988f
C276 VDD2.n47 B 0.022309f
C277 VDD2.n48 B 0.022309f
C278 VDD2.n49 B 0.011988f
C279 VDD2.n50 B 0.012693f
C280 VDD2.n51 B 0.028335f
C281 VDD2.n52 B 0.060541f
C282 VDD2.n53 B 0.012693f
C283 VDD2.n54 B 0.011988f
C284 VDD2.n55 B 0.05309f
C285 VDD2.n56 B 0.055992f
C286 VDD2.t0 B 0.18916f
C287 VDD2.t1 B 0.18916f
C288 VDD2.n57 B 1.67438f
C289 VDD2.n58 B 0.527506f
C290 VDD2.t2 B 0.18916f
C291 VDD2.t5 B 0.18916f
C292 VDD2.n59 B 1.68359f
C293 VDD2.n60 B 2.19468f
C294 VDD2.n61 B 0.030906f
C295 VDD2.n62 B 0.022309f
C296 VDD2.n63 B 0.011988f
C297 VDD2.n64 B 0.028335f
C298 VDD2.n65 B 0.012693f
C299 VDD2.n66 B 0.022309f
C300 VDD2.n67 B 0.011988f
C301 VDD2.n68 B 0.028335f
C302 VDD2.n69 B 0.012693f
C303 VDD2.n70 B 0.022309f
C304 VDD2.n71 B 0.011988f
C305 VDD2.n72 B 0.028335f
C306 VDD2.n73 B 0.028335f
C307 VDD2.n74 B 0.012693f
C308 VDD2.n75 B 0.022309f
C309 VDD2.n76 B 0.011988f
C310 VDD2.n77 B 0.028335f
C311 VDD2.n78 B 0.012693f
C312 VDD2.n79 B 0.149968f
C313 VDD2.t6 B 0.047704f
C314 VDD2.n80 B 0.021251f
C315 VDD2.n81 B 0.020031f
C316 VDD2.n82 B 0.011988f
C317 VDD2.n83 B 0.999421f
C318 VDD2.n84 B 0.022309f
C319 VDD2.n85 B 0.011988f
C320 VDD2.n86 B 0.012693f
C321 VDD2.n87 B 0.028335f
C322 VDD2.n88 B 0.028335f
C323 VDD2.n89 B 0.012693f
C324 VDD2.n90 B 0.011988f
C325 VDD2.n91 B 0.022309f
C326 VDD2.n92 B 0.022309f
C327 VDD2.n93 B 0.011988f
C328 VDD2.n94 B 0.012693f
C329 VDD2.n95 B 0.028335f
C330 VDD2.n96 B 0.028335f
C331 VDD2.n97 B 0.012693f
C332 VDD2.n98 B 0.011988f
C333 VDD2.n99 B 0.022309f
C334 VDD2.n100 B 0.022309f
C335 VDD2.n101 B 0.011988f
C336 VDD2.n102 B 0.01234f
C337 VDD2.n103 B 0.01234f
C338 VDD2.n104 B 0.028335f
C339 VDD2.n105 B 0.028335f
C340 VDD2.n106 B 0.012693f
C341 VDD2.n107 B 0.011988f
C342 VDD2.n108 B 0.022309f
C343 VDD2.n109 B 0.022309f
C344 VDD2.n110 B 0.011988f
C345 VDD2.n111 B 0.012693f
C346 VDD2.n112 B 0.028335f
C347 VDD2.n113 B 0.060541f
C348 VDD2.n114 B 0.012693f
C349 VDD2.n115 B 0.011988f
C350 VDD2.n116 B 0.05309f
C351 VDD2.n117 B 0.049231f
C352 VDD2.n118 B 2.24934f
C353 VDD2.t8 B 0.18916f
C354 VDD2.t3 B 0.18916f
C355 VDD2.n119 B 1.67439f
C356 VDD2.n120 B 0.359185f
C357 VDD2.t7 B 0.18916f
C358 VDD2.t4 B 0.18916f
C359 VDD2.n121 B 1.68356f
C360 VTAIL.t10 B 0.211037f
C361 VTAIL.t11 B 0.211037f
C362 VTAIL.n0 B 1.79699f
C363 VTAIL.n1 B 0.475623f
C364 VTAIL.n2 B 0.03448f
C365 VTAIL.n3 B 0.024889f
C366 VTAIL.n4 B 0.013374f
C367 VTAIL.n5 B 0.031612f
C368 VTAIL.n6 B 0.014161f
C369 VTAIL.n7 B 0.024889f
C370 VTAIL.n8 B 0.013374f
C371 VTAIL.n9 B 0.031612f
C372 VTAIL.n10 B 0.014161f
C373 VTAIL.n11 B 0.024889f
C374 VTAIL.n12 B 0.013374f
C375 VTAIL.n13 B 0.031612f
C376 VTAIL.n14 B 0.014161f
C377 VTAIL.n15 B 0.024889f
C378 VTAIL.n16 B 0.013374f
C379 VTAIL.n17 B 0.031612f
C380 VTAIL.n18 B 0.014161f
C381 VTAIL.n19 B 0.167313f
C382 VTAIL.t7 B 0.053221f
C383 VTAIL.n20 B 0.023709f
C384 VTAIL.n21 B 0.022347f
C385 VTAIL.n22 B 0.013374f
C386 VTAIL.n23 B 1.11501f
C387 VTAIL.n24 B 0.024889f
C388 VTAIL.n25 B 0.013374f
C389 VTAIL.n26 B 0.014161f
C390 VTAIL.n27 B 0.031612f
C391 VTAIL.n28 B 0.031612f
C392 VTAIL.n29 B 0.014161f
C393 VTAIL.n30 B 0.013374f
C394 VTAIL.n31 B 0.024889f
C395 VTAIL.n32 B 0.024889f
C396 VTAIL.n33 B 0.013374f
C397 VTAIL.n34 B 0.014161f
C398 VTAIL.n35 B 0.031612f
C399 VTAIL.n36 B 0.031612f
C400 VTAIL.n37 B 0.031612f
C401 VTAIL.n38 B 0.014161f
C402 VTAIL.n39 B 0.013374f
C403 VTAIL.n40 B 0.024889f
C404 VTAIL.n41 B 0.024889f
C405 VTAIL.n42 B 0.013374f
C406 VTAIL.n43 B 0.013768f
C407 VTAIL.n44 B 0.013768f
C408 VTAIL.n45 B 0.031612f
C409 VTAIL.n46 B 0.031612f
C410 VTAIL.n47 B 0.014161f
C411 VTAIL.n48 B 0.013374f
C412 VTAIL.n49 B 0.024889f
C413 VTAIL.n50 B 0.024889f
C414 VTAIL.n51 B 0.013374f
C415 VTAIL.n52 B 0.014161f
C416 VTAIL.n53 B 0.031612f
C417 VTAIL.n54 B 0.067543f
C418 VTAIL.n55 B 0.014161f
C419 VTAIL.n56 B 0.013374f
C420 VTAIL.n57 B 0.05923f
C421 VTAIL.n58 B 0.037753f
C422 VTAIL.n59 B 0.291156f
C423 VTAIL.t5 B 0.211037f
C424 VTAIL.t19 B 0.211037f
C425 VTAIL.n60 B 1.79699f
C426 VTAIL.n61 B 0.548907f
C427 VTAIL.t1 B 0.211037f
C428 VTAIL.t2 B 0.211037f
C429 VTAIL.n62 B 1.79699f
C430 VTAIL.n63 B 1.78299f
C431 VTAIL.t17 B 0.211037f
C432 VTAIL.t13 B 0.211037f
C433 VTAIL.n64 B 1.797f
C434 VTAIL.n65 B 1.78298f
C435 VTAIL.t18 B 0.211037f
C436 VTAIL.t14 B 0.211037f
C437 VTAIL.n66 B 1.797f
C438 VTAIL.n67 B 0.548897f
C439 VTAIL.n68 B 0.03448f
C440 VTAIL.n69 B 0.024889f
C441 VTAIL.n70 B 0.013374f
C442 VTAIL.n71 B 0.031612f
C443 VTAIL.n72 B 0.014161f
C444 VTAIL.n73 B 0.024889f
C445 VTAIL.n74 B 0.013374f
C446 VTAIL.n75 B 0.031612f
C447 VTAIL.n76 B 0.014161f
C448 VTAIL.n77 B 0.024889f
C449 VTAIL.n78 B 0.013374f
C450 VTAIL.n79 B 0.031612f
C451 VTAIL.n80 B 0.031612f
C452 VTAIL.n81 B 0.014161f
C453 VTAIL.n82 B 0.024889f
C454 VTAIL.n83 B 0.013374f
C455 VTAIL.n84 B 0.031612f
C456 VTAIL.n85 B 0.014161f
C457 VTAIL.n86 B 0.167313f
C458 VTAIL.t12 B 0.053221f
C459 VTAIL.n87 B 0.023709f
C460 VTAIL.n88 B 0.022347f
C461 VTAIL.n89 B 0.013374f
C462 VTAIL.n90 B 1.11501f
C463 VTAIL.n91 B 0.024889f
C464 VTAIL.n92 B 0.013374f
C465 VTAIL.n93 B 0.014161f
C466 VTAIL.n94 B 0.031612f
C467 VTAIL.n95 B 0.031612f
C468 VTAIL.n96 B 0.014161f
C469 VTAIL.n97 B 0.013374f
C470 VTAIL.n98 B 0.024889f
C471 VTAIL.n99 B 0.024889f
C472 VTAIL.n100 B 0.013374f
C473 VTAIL.n101 B 0.014161f
C474 VTAIL.n102 B 0.031612f
C475 VTAIL.n103 B 0.031612f
C476 VTAIL.n104 B 0.014161f
C477 VTAIL.n105 B 0.013374f
C478 VTAIL.n106 B 0.024889f
C479 VTAIL.n107 B 0.024889f
C480 VTAIL.n108 B 0.013374f
C481 VTAIL.n109 B 0.013768f
C482 VTAIL.n110 B 0.013768f
C483 VTAIL.n111 B 0.031612f
C484 VTAIL.n112 B 0.031612f
C485 VTAIL.n113 B 0.014161f
C486 VTAIL.n114 B 0.013374f
C487 VTAIL.n115 B 0.024889f
C488 VTAIL.n116 B 0.024889f
C489 VTAIL.n117 B 0.013374f
C490 VTAIL.n118 B 0.014161f
C491 VTAIL.n119 B 0.031612f
C492 VTAIL.n120 B 0.067543f
C493 VTAIL.n121 B 0.014161f
C494 VTAIL.n122 B 0.013374f
C495 VTAIL.n123 B 0.05923f
C496 VTAIL.n124 B 0.037753f
C497 VTAIL.n125 B 0.291156f
C498 VTAIL.t0 B 0.211037f
C499 VTAIL.t3 B 0.211037f
C500 VTAIL.n126 B 1.797f
C501 VTAIL.n127 B 0.509489f
C502 VTAIL.t8 B 0.211037f
C503 VTAIL.t4 B 0.211037f
C504 VTAIL.n128 B 1.797f
C505 VTAIL.n129 B 0.548897f
C506 VTAIL.n130 B 0.03448f
C507 VTAIL.n131 B 0.024889f
C508 VTAIL.n132 B 0.013374f
C509 VTAIL.n133 B 0.031612f
C510 VTAIL.n134 B 0.014161f
C511 VTAIL.n135 B 0.024889f
C512 VTAIL.n136 B 0.013374f
C513 VTAIL.n137 B 0.031612f
C514 VTAIL.n138 B 0.014161f
C515 VTAIL.n139 B 0.024889f
C516 VTAIL.n140 B 0.013374f
C517 VTAIL.n141 B 0.031612f
C518 VTAIL.n142 B 0.031612f
C519 VTAIL.n143 B 0.014161f
C520 VTAIL.n144 B 0.024889f
C521 VTAIL.n145 B 0.013374f
C522 VTAIL.n146 B 0.031612f
C523 VTAIL.n147 B 0.014161f
C524 VTAIL.n148 B 0.167313f
C525 VTAIL.t6 B 0.053221f
C526 VTAIL.n149 B 0.023709f
C527 VTAIL.n150 B 0.022347f
C528 VTAIL.n151 B 0.013374f
C529 VTAIL.n152 B 1.11501f
C530 VTAIL.n153 B 0.024889f
C531 VTAIL.n154 B 0.013374f
C532 VTAIL.n155 B 0.014161f
C533 VTAIL.n156 B 0.031612f
C534 VTAIL.n157 B 0.031612f
C535 VTAIL.n158 B 0.014161f
C536 VTAIL.n159 B 0.013374f
C537 VTAIL.n160 B 0.024889f
C538 VTAIL.n161 B 0.024889f
C539 VTAIL.n162 B 0.013374f
C540 VTAIL.n163 B 0.014161f
C541 VTAIL.n164 B 0.031612f
C542 VTAIL.n165 B 0.031612f
C543 VTAIL.n166 B 0.014161f
C544 VTAIL.n167 B 0.013374f
C545 VTAIL.n168 B 0.024889f
C546 VTAIL.n169 B 0.024889f
C547 VTAIL.n170 B 0.013374f
C548 VTAIL.n171 B 0.013768f
C549 VTAIL.n172 B 0.013768f
C550 VTAIL.n173 B 0.031612f
C551 VTAIL.n174 B 0.031612f
C552 VTAIL.n175 B 0.014161f
C553 VTAIL.n176 B 0.013374f
C554 VTAIL.n177 B 0.024889f
C555 VTAIL.n178 B 0.024889f
C556 VTAIL.n179 B 0.013374f
C557 VTAIL.n180 B 0.014161f
C558 VTAIL.n181 B 0.031612f
C559 VTAIL.n182 B 0.067543f
C560 VTAIL.n183 B 0.014161f
C561 VTAIL.n184 B 0.013374f
C562 VTAIL.n185 B 0.05923f
C563 VTAIL.n186 B 0.037753f
C564 VTAIL.n187 B 1.41048f
C565 VTAIL.n188 B 0.03448f
C566 VTAIL.n189 B 0.024889f
C567 VTAIL.n190 B 0.013374f
C568 VTAIL.n191 B 0.031612f
C569 VTAIL.n192 B 0.014161f
C570 VTAIL.n193 B 0.024889f
C571 VTAIL.n194 B 0.013374f
C572 VTAIL.n195 B 0.031612f
C573 VTAIL.n196 B 0.014161f
C574 VTAIL.n197 B 0.024889f
C575 VTAIL.n198 B 0.013374f
C576 VTAIL.n199 B 0.031612f
C577 VTAIL.n200 B 0.014161f
C578 VTAIL.n201 B 0.024889f
C579 VTAIL.n202 B 0.013374f
C580 VTAIL.n203 B 0.031612f
C581 VTAIL.n204 B 0.014161f
C582 VTAIL.n205 B 0.167313f
C583 VTAIL.t16 B 0.053221f
C584 VTAIL.n206 B 0.023709f
C585 VTAIL.n207 B 0.022347f
C586 VTAIL.n208 B 0.013374f
C587 VTAIL.n209 B 1.11501f
C588 VTAIL.n210 B 0.024889f
C589 VTAIL.n211 B 0.013374f
C590 VTAIL.n212 B 0.014161f
C591 VTAIL.n213 B 0.031612f
C592 VTAIL.n214 B 0.031612f
C593 VTAIL.n215 B 0.014161f
C594 VTAIL.n216 B 0.013374f
C595 VTAIL.n217 B 0.024889f
C596 VTAIL.n218 B 0.024889f
C597 VTAIL.n219 B 0.013374f
C598 VTAIL.n220 B 0.014161f
C599 VTAIL.n221 B 0.031612f
C600 VTAIL.n222 B 0.031612f
C601 VTAIL.n223 B 0.031612f
C602 VTAIL.n224 B 0.014161f
C603 VTAIL.n225 B 0.013374f
C604 VTAIL.n226 B 0.024889f
C605 VTAIL.n227 B 0.024889f
C606 VTAIL.n228 B 0.013374f
C607 VTAIL.n229 B 0.013768f
C608 VTAIL.n230 B 0.013768f
C609 VTAIL.n231 B 0.031612f
C610 VTAIL.n232 B 0.031612f
C611 VTAIL.n233 B 0.014161f
C612 VTAIL.n234 B 0.013374f
C613 VTAIL.n235 B 0.024889f
C614 VTAIL.n236 B 0.024889f
C615 VTAIL.n237 B 0.013374f
C616 VTAIL.n238 B 0.014161f
C617 VTAIL.n239 B 0.031612f
C618 VTAIL.n240 B 0.067543f
C619 VTAIL.n241 B 0.014161f
C620 VTAIL.n242 B 0.013374f
C621 VTAIL.n243 B 0.05923f
C622 VTAIL.n244 B 0.037753f
C623 VTAIL.n245 B 1.41048f
C624 VTAIL.t15 B 0.211037f
C625 VTAIL.t9 B 0.211037f
C626 VTAIL.n246 B 1.79699f
C627 VTAIL.n247 B 0.428611f
C628 VN.n0 B 0.034617f
C629 VN.t4 B 1.45356f
C630 VN.n1 B 0.045151f
C631 VN.n2 B 0.026257f
C632 VN.t7 B 1.45356f
C633 VN.n3 B 0.026054f
C634 VN.n4 B 0.026257f
C635 VN.t8 B 1.45356f
C636 VN.n5 B 0.026054f
C637 VN.n6 B 0.194219f
C638 VN.t9 B 1.45356f
C639 VN.t0 B 1.57382f
C640 VN.n7 B 0.591542f
C641 VN.n8 B 0.583979f
C642 VN.n9 B 0.03589f
C643 VN.n10 B 0.04741f
C644 VN.n11 B 0.026257f
C645 VN.n12 B 0.026257f
C646 VN.n13 B 0.026257f
C647 VN.n14 B 0.052137f
C648 VN.n15 B 0.548989f
C649 VN.n16 B 0.052137f
C650 VN.n17 B 0.026257f
C651 VN.n18 B 0.026257f
C652 VN.n19 B 0.026257f
C653 VN.n20 B 0.04741f
C654 VN.n21 B 0.03589f
C655 VN.n22 B 0.524213f
C656 VN.n23 B 0.037823f
C657 VN.n24 B 0.026257f
C658 VN.n25 B 0.026257f
C659 VN.n26 B 0.026257f
C660 VN.n27 B 0.030629f
C661 VN.n28 B 0.047889f
C662 VN.n29 B 0.605006f
C663 VN.n30 B 0.029368f
C664 VN.n31 B 0.034617f
C665 VN.t3 B 1.45356f
C666 VN.n32 B 0.045151f
C667 VN.n33 B 0.026257f
C668 VN.t1 B 1.45356f
C669 VN.n34 B 0.026054f
C670 VN.n35 B 0.026257f
C671 VN.t6 B 1.45356f
C672 VN.n36 B 0.026054f
C673 VN.n37 B 0.194219f
C674 VN.t2 B 1.45356f
C675 VN.t5 B 1.57382f
C676 VN.n38 B 0.591542f
C677 VN.n39 B 0.583979f
C678 VN.n40 B 0.03589f
C679 VN.n41 B 0.04741f
C680 VN.n42 B 0.026257f
C681 VN.n43 B 0.026257f
C682 VN.n44 B 0.026257f
C683 VN.n45 B 0.052137f
C684 VN.n46 B 0.548989f
C685 VN.n47 B 0.052137f
C686 VN.n48 B 0.026257f
C687 VN.n49 B 0.026257f
C688 VN.n50 B 0.026257f
C689 VN.n51 B 0.04741f
C690 VN.n52 B 0.03589f
C691 VN.n53 B 0.524213f
C692 VN.n54 B 0.037823f
C693 VN.n55 B 0.026257f
C694 VN.n56 B 0.026257f
C695 VN.n57 B 0.026257f
C696 VN.n58 B 0.030629f
C697 VN.n59 B 0.047889f
C698 VN.n60 B 0.605006f
C699 VN.n61 B 1.39206f
.ends

