* NGSPICE file created from diff_pair_sample_0952.ext - technology: sky130A

.subckt diff_pair_sample_0952 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t9 w_n3794_n2936# sky130_fd_pr__pfet_01v8 ad=1.6236 pd=10.17 as=3.8376 ps=20.46 w=9.84 l=3.2
X1 VDD1.t4 VP.t1 VTAIL.t11 w_n3794_n2936# sky130_fd_pr__pfet_01v8 ad=1.6236 pd=10.17 as=3.8376 ps=20.46 w=9.84 l=3.2
X2 B.t11 B.t9 B.t10 w_n3794_n2936# sky130_fd_pr__pfet_01v8 ad=3.8376 pd=20.46 as=0 ps=0 w=9.84 l=3.2
X3 B.t8 B.t6 B.t7 w_n3794_n2936# sky130_fd_pr__pfet_01v8 ad=3.8376 pd=20.46 as=0 ps=0 w=9.84 l=3.2
X4 VTAIL.t7 VP.t2 VDD1.t3 w_n3794_n2936# sky130_fd_pr__pfet_01v8 ad=1.6236 pd=10.17 as=1.6236 ps=10.17 w=9.84 l=3.2
X5 VDD2.t5 VN.t0 VTAIL.t5 w_n3794_n2936# sky130_fd_pr__pfet_01v8 ad=1.6236 pd=10.17 as=3.8376 ps=20.46 w=9.84 l=3.2
X6 VTAIL.t4 VN.t1 VDD2.t4 w_n3794_n2936# sky130_fd_pr__pfet_01v8 ad=1.6236 pd=10.17 as=1.6236 ps=10.17 w=9.84 l=3.2
X7 VDD2.t3 VN.t2 VTAIL.t2 w_n3794_n2936# sky130_fd_pr__pfet_01v8 ad=3.8376 pd=20.46 as=1.6236 ps=10.17 w=9.84 l=3.2
X8 VTAIL.t0 VN.t3 VDD2.t2 w_n3794_n2936# sky130_fd_pr__pfet_01v8 ad=1.6236 pd=10.17 as=1.6236 ps=10.17 w=9.84 l=3.2
X9 VDD1.t2 VP.t3 VTAIL.t8 w_n3794_n2936# sky130_fd_pr__pfet_01v8 ad=3.8376 pd=20.46 as=1.6236 ps=10.17 w=9.84 l=3.2
X10 B.t5 B.t3 B.t4 w_n3794_n2936# sky130_fd_pr__pfet_01v8 ad=3.8376 pd=20.46 as=0 ps=0 w=9.84 l=3.2
X11 VDD2.t1 VN.t4 VTAIL.t1 w_n3794_n2936# sky130_fd_pr__pfet_01v8 ad=1.6236 pd=10.17 as=3.8376 ps=20.46 w=9.84 l=3.2
X12 B.t2 B.t0 B.t1 w_n3794_n2936# sky130_fd_pr__pfet_01v8 ad=3.8376 pd=20.46 as=0 ps=0 w=9.84 l=3.2
X13 VTAIL.t6 VP.t4 VDD1.t1 w_n3794_n2936# sky130_fd_pr__pfet_01v8 ad=1.6236 pd=10.17 as=1.6236 ps=10.17 w=9.84 l=3.2
X14 VDD1.t0 VP.t5 VTAIL.t10 w_n3794_n2936# sky130_fd_pr__pfet_01v8 ad=3.8376 pd=20.46 as=1.6236 ps=10.17 w=9.84 l=3.2
X15 VDD2.t0 VN.t5 VTAIL.t3 w_n3794_n2936# sky130_fd_pr__pfet_01v8 ad=3.8376 pd=20.46 as=1.6236 ps=10.17 w=9.84 l=3.2
R0 VP.n16 VP.n15 161.3
R1 VP.n17 VP.n12 161.3
R2 VP.n19 VP.n18 161.3
R3 VP.n20 VP.n11 161.3
R4 VP.n22 VP.n21 161.3
R5 VP.n23 VP.n10 161.3
R6 VP.n25 VP.n24 161.3
R7 VP.n49 VP.n48 161.3
R8 VP.n47 VP.n1 161.3
R9 VP.n46 VP.n45 161.3
R10 VP.n44 VP.n2 161.3
R11 VP.n43 VP.n42 161.3
R12 VP.n41 VP.n3 161.3
R13 VP.n40 VP.n39 161.3
R14 VP.n38 VP.n37 161.3
R15 VP.n36 VP.n5 161.3
R16 VP.n35 VP.n34 161.3
R17 VP.n33 VP.n6 161.3
R18 VP.n32 VP.n31 161.3
R19 VP.n30 VP.n7 161.3
R20 VP.n29 VP.n28 161.3
R21 VP.n14 VP.t3 107.028
R22 VP.n27 VP.n8 76.4741
R23 VP.n50 VP.n0 76.4741
R24 VP.n26 VP.n9 76.4741
R25 VP.n8 VP.t5 74.108
R26 VP.n4 VP.t4 74.108
R27 VP.n0 VP.t1 74.108
R28 VP.n9 VP.t0 74.108
R29 VP.n13 VP.t2 74.108
R30 VP.n14 VP.n13 62.2079
R31 VP.n27 VP.n26 49.4655
R32 VP.n31 VP.n6 42.0302
R33 VP.n46 VP.n2 42.0302
R34 VP.n22 VP.n11 42.0302
R35 VP.n35 VP.n6 39.1239
R36 VP.n42 VP.n2 39.1239
R37 VP.n18 VP.n11 39.1239
R38 VP.n30 VP.n29 24.5923
R39 VP.n31 VP.n30 24.5923
R40 VP.n36 VP.n35 24.5923
R41 VP.n37 VP.n36 24.5923
R42 VP.n41 VP.n40 24.5923
R43 VP.n42 VP.n41 24.5923
R44 VP.n47 VP.n46 24.5923
R45 VP.n48 VP.n47 24.5923
R46 VP.n23 VP.n22 24.5923
R47 VP.n24 VP.n23 24.5923
R48 VP.n17 VP.n16 24.5923
R49 VP.n18 VP.n17 24.5923
R50 VP.n29 VP.n8 13.7719
R51 VP.n48 VP.n0 13.7719
R52 VP.n24 VP.n9 13.7719
R53 VP.n37 VP.n4 12.2964
R54 VP.n40 VP.n4 12.2964
R55 VP.n16 VP.n13 12.2964
R56 VP.n15 VP.n14 4.19125
R57 VP.n26 VP.n25 0.354861
R58 VP.n28 VP.n27 0.354861
R59 VP.n50 VP.n49 0.354861
R60 VP VP.n50 0.267071
R61 VP.n15 VP.n12 0.189894
R62 VP.n19 VP.n12 0.189894
R63 VP.n20 VP.n19 0.189894
R64 VP.n21 VP.n20 0.189894
R65 VP.n21 VP.n10 0.189894
R66 VP.n25 VP.n10 0.189894
R67 VP.n28 VP.n7 0.189894
R68 VP.n32 VP.n7 0.189894
R69 VP.n33 VP.n32 0.189894
R70 VP.n34 VP.n33 0.189894
R71 VP.n34 VP.n5 0.189894
R72 VP.n38 VP.n5 0.189894
R73 VP.n39 VP.n38 0.189894
R74 VP.n39 VP.n3 0.189894
R75 VP.n43 VP.n3 0.189894
R76 VP.n44 VP.n43 0.189894
R77 VP.n45 VP.n44 0.189894
R78 VP.n45 VP.n1 0.189894
R79 VP.n49 VP.n1 0.189894
R80 VTAIL.n7 VTAIL.t5 62.4885
R81 VTAIL.n10 VTAIL.t9 62.4885
R82 VTAIL.n11 VTAIL.t1 62.4883
R83 VTAIL.n2 VTAIL.t11 62.4883
R84 VTAIL.n9 VTAIL.n8 59.1851
R85 VTAIL.n6 VTAIL.n5 59.1851
R86 VTAIL.n1 VTAIL.n0 59.1849
R87 VTAIL.n4 VTAIL.n3 59.1849
R88 VTAIL.n6 VTAIL.n4 26.9358
R89 VTAIL.n11 VTAIL.n10 23.8927
R90 VTAIL.n0 VTAIL.t3 3.30385
R91 VTAIL.n0 VTAIL.t0 3.30385
R92 VTAIL.n3 VTAIL.t10 3.30385
R93 VTAIL.n3 VTAIL.t6 3.30385
R94 VTAIL.n8 VTAIL.t8 3.30385
R95 VTAIL.n8 VTAIL.t7 3.30385
R96 VTAIL.n5 VTAIL.t2 3.30385
R97 VTAIL.n5 VTAIL.t4 3.30385
R98 VTAIL.n7 VTAIL.n6 3.0436
R99 VTAIL.n10 VTAIL.n9 3.0436
R100 VTAIL.n4 VTAIL.n2 3.0436
R101 VTAIL VTAIL.n11 2.22464
R102 VTAIL.n9 VTAIL.n7 1.99188
R103 VTAIL.n2 VTAIL.n1 1.99188
R104 VTAIL VTAIL.n1 0.819465
R105 VDD1 VDD1.t2 81.5078
R106 VDD1.n1 VDD1.t0 81.394
R107 VDD1.n1 VDD1.n0 76.5691
R108 VDD1.n3 VDD1.n2 75.8639
R109 VDD1.n3 VDD1.n1 44.1927
R110 VDD1.n2 VDD1.t3 3.30385
R111 VDD1.n2 VDD1.t5 3.30385
R112 VDD1.n0 VDD1.t1 3.30385
R113 VDD1.n0 VDD1.t4 3.30385
R114 VDD1 VDD1.n3 0.703086
R115 B.n382 B.n121 585
R116 B.n381 B.n380 585
R117 B.n379 B.n122 585
R118 B.n378 B.n377 585
R119 B.n376 B.n123 585
R120 B.n375 B.n374 585
R121 B.n373 B.n124 585
R122 B.n372 B.n371 585
R123 B.n370 B.n125 585
R124 B.n369 B.n368 585
R125 B.n367 B.n126 585
R126 B.n366 B.n365 585
R127 B.n364 B.n127 585
R128 B.n363 B.n362 585
R129 B.n361 B.n128 585
R130 B.n360 B.n359 585
R131 B.n358 B.n129 585
R132 B.n357 B.n356 585
R133 B.n355 B.n130 585
R134 B.n354 B.n353 585
R135 B.n352 B.n131 585
R136 B.n351 B.n350 585
R137 B.n349 B.n132 585
R138 B.n348 B.n347 585
R139 B.n346 B.n133 585
R140 B.n345 B.n344 585
R141 B.n343 B.n134 585
R142 B.n342 B.n341 585
R143 B.n340 B.n135 585
R144 B.n339 B.n338 585
R145 B.n337 B.n136 585
R146 B.n336 B.n335 585
R147 B.n334 B.n137 585
R148 B.n333 B.n332 585
R149 B.n331 B.n138 585
R150 B.n330 B.n329 585
R151 B.n325 B.n139 585
R152 B.n324 B.n323 585
R153 B.n322 B.n140 585
R154 B.n321 B.n320 585
R155 B.n319 B.n141 585
R156 B.n318 B.n317 585
R157 B.n316 B.n142 585
R158 B.n315 B.n314 585
R159 B.n313 B.n143 585
R160 B.n311 B.n310 585
R161 B.n309 B.n146 585
R162 B.n308 B.n307 585
R163 B.n306 B.n147 585
R164 B.n305 B.n304 585
R165 B.n303 B.n148 585
R166 B.n302 B.n301 585
R167 B.n300 B.n149 585
R168 B.n299 B.n298 585
R169 B.n297 B.n150 585
R170 B.n296 B.n295 585
R171 B.n294 B.n151 585
R172 B.n293 B.n292 585
R173 B.n291 B.n152 585
R174 B.n290 B.n289 585
R175 B.n288 B.n153 585
R176 B.n287 B.n286 585
R177 B.n285 B.n154 585
R178 B.n284 B.n283 585
R179 B.n282 B.n155 585
R180 B.n281 B.n280 585
R181 B.n279 B.n156 585
R182 B.n278 B.n277 585
R183 B.n276 B.n157 585
R184 B.n275 B.n274 585
R185 B.n273 B.n158 585
R186 B.n272 B.n271 585
R187 B.n270 B.n159 585
R188 B.n269 B.n268 585
R189 B.n267 B.n160 585
R190 B.n266 B.n265 585
R191 B.n264 B.n161 585
R192 B.n263 B.n262 585
R193 B.n261 B.n162 585
R194 B.n260 B.n259 585
R195 B.n384 B.n383 585
R196 B.n385 B.n120 585
R197 B.n387 B.n386 585
R198 B.n388 B.n119 585
R199 B.n390 B.n389 585
R200 B.n391 B.n118 585
R201 B.n393 B.n392 585
R202 B.n394 B.n117 585
R203 B.n396 B.n395 585
R204 B.n397 B.n116 585
R205 B.n399 B.n398 585
R206 B.n400 B.n115 585
R207 B.n402 B.n401 585
R208 B.n403 B.n114 585
R209 B.n405 B.n404 585
R210 B.n406 B.n113 585
R211 B.n408 B.n407 585
R212 B.n409 B.n112 585
R213 B.n411 B.n410 585
R214 B.n412 B.n111 585
R215 B.n414 B.n413 585
R216 B.n415 B.n110 585
R217 B.n417 B.n416 585
R218 B.n418 B.n109 585
R219 B.n420 B.n419 585
R220 B.n421 B.n108 585
R221 B.n423 B.n422 585
R222 B.n424 B.n107 585
R223 B.n426 B.n425 585
R224 B.n427 B.n106 585
R225 B.n429 B.n428 585
R226 B.n430 B.n105 585
R227 B.n432 B.n431 585
R228 B.n433 B.n104 585
R229 B.n435 B.n434 585
R230 B.n436 B.n103 585
R231 B.n438 B.n437 585
R232 B.n439 B.n102 585
R233 B.n441 B.n440 585
R234 B.n442 B.n101 585
R235 B.n444 B.n443 585
R236 B.n445 B.n100 585
R237 B.n447 B.n446 585
R238 B.n448 B.n99 585
R239 B.n450 B.n449 585
R240 B.n451 B.n98 585
R241 B.n453 B.n452 585
R242 B.n454 B.n97 585
R243 B.n456 B.n455 585
R244 B.n457 B.n96 585
R245 B.n459 B.n458 585
R246 B.n460 B.n95 585
R247 B.n462 B.n461 585
R248 B.n463 B.n94 585
R249 B.n465 B.n464 585
R250 B.n466 B.n93 585
R251 B.n468 B.n467 585
R252 B.n469 B.n92 585
R253 B.n471 B.n470 585
R254 B.n472 B.n91 585
R255 B.n474 B.n473 585
R256 B.n475 B.n90 585
R257 B.n477 B.n476 585
R258 B.n478 B.n89 585
R259 B.n480 B.n479 585
R260 B.n481 B.n88 585
R261 B.n483 B.n482 585
R262 B.n484 B.n87 585
R263 B.n486 B.n485 585
R264 B.n487 B.n86 585
R265 B.n489 B.n488 585
R266 B.n490 B.n85 585
R267 B.n492 B.n491 585
R268 B.n493 B.n84 585
R269 B.n495 B.n494 585
R270 B.n496 B.n83 585
R271 B.n498 B.n497 585
R272 B.n499 B.n82 585
R273 B.n501 B.n500 585
R274 B.n502 B.n81 585
R275 B.n504 B.n503 585
R276 B.n505 B.n80 585
R277 B.n507 B.n506 585
R278 B.n508 B.n79 585
R279 B.n510 B.n509 585
R280 B.n511 B.n78 585
R281 B.n513 B.n512 585
R282 B.n514 B.n77 585
R283 B.n516 B.n515 585
R284 B.n517 B.n76 585
R285 B.n519 B.n518 585
R286 B.n520 B.n75 585
R287 B.n522 B.n521 585
R288 B.n523 B.n74 585
R289 B.n525 B.n524 585
R290 B.n526 B.n73 585
R291 B.n528 B.n527 585
R292 B.n529 B.n72 585
R293 B.n531 B.n530 585
R294 B.n532 B.n71 585
R295 B.n654 B.n653 585
R296 B.n652 B.n27 585
R297 B.n651 B.n650 585
R298 B.n649 B.n28 585
R299 B.n648 B.n647 585
R300 B.n646 B.n29 585
R301 B.n645 B.n644 585
R302 B.n643 B.n30 585
R303 B.n642 B.n641 585
R304 B.n640 B.n31 585
R305 B.n639 B.n638 585
R306 B.n637 B.n32 585
R307 B.n636 B.n635 585
R308 B.n634 B.n33 585
R309 B.n633 B.n632 585
R310 B.n631 B.n34 585
R311 B.n630 B.n629 585
R312 B.n628 B.n35 585
R313 B.n627 B.n626 585
R314 B.n625 B.n36 585
R315 B.n624 B.n623 585
R316 B.n622 B.n37 585
R317 B.n621 B.n620 585
R318 B.n619 B.n38 585
R319 B.n618 B.n617 585
R320 B.n616 B.n39 585
R321 B.n615 B.n614 585
R322 B.n613 B.n40 585
R323 B.n612 B.n611 585
R324 B.n610 B.n41 585
R325 B.n609 B.n608 585
R326 B.n607 B.n42 585
R327 B.n606 B.n605 585
R328 B.n604 B.n43 585
R329 B.n603 B.n602 585
R330 B.n601 B.n600 585
R331 B.n599 B.n47 585
R332 B.n598 B.n597 585
R333 B.n596 B.n48 585
R334 B.n595 B.n594 585
R335 B.n593 B.n49 585
R336 B.n592 B.n591 585
R337 B.n590 B.n50 585
R338 B.n589 B.n588 585
R339 B.n587 B.n51 585
R340 B.n585 B.n584 585
R341 B.n583 B.n54 585
R342 B.n582 B.n581 585
R343 B.n580 B.n55 585
R344 B.n579 B.n578 585
R345 B.n577 B.n56 585
R346 B.n576 B.n575 585
R347 B.n574 B.n57 585
R348 B.n573 B.n572 585
R349 B.n571 B.n58 585
R350 B.n570 B.n569 585
R351 B.n568 B.n59 585
R352 B.n567 B.n566 585
R353 B.n565 B.n60 585
R354 B.n564 B.n563 585
R355 B.n562 B.n61 585
R356 B.n561 B.n560 585
R357 B.n559 B.n62 585
R358 B.n558 B.n557 585
R359 B.n556 B.n63 585
R360 B.n555 B.n554 585
R361 B.n553 B.n64 585
R362 B.n552 B.n551 585
R363 B.n550 B.n65 585
R364 B.n549 B.n548 585
R365 B.n547 B.n66 585
R366 B.n546 B.n545 585
R367 B.n544 B.n67 585
R368 B.n543 B.n542 585
R369 B.n541 B.n68 585
R370 B.n540 B.n539 585
R371 B.n538 B.n69 585
R372 B.n537 B.n536 585
R373 B.n535 B.n70 585
R374 B.n534 B.n533 585
R375 B.n655 B.n26 585
R376 B.n657 B.n656 585
R377 B.n658 B.n25 585
R378 B.n660 B.n659 585
R379 B.n661 B.n24 585
R380 B.n663 B.n662 585
R381 B.n664 B.n23 585
R382 B.n666 B.n665 585
R383 B.n667 B.n22 585
R384 B.n669 B.n668 585
R385 B.n670 B.n21 585
R386 B.n672 B.n671 585
R387 B.n673 B.n20 585
R388 B.n675 B.n674 585
R389 B.n676 B.n19 585
R390 B.n678 B.n677 585
R391 B.n679 B.n18 585
R392 B.n681 B.n680 585
R393 B.n682 B.n17 585
R394 B.n684 B.n683 585
R395 B.n685 B.n16 585
R396 B.n687 B.n686 585
R397 B.n688 B.n15 585
R398 B.n690 B.n689 585
R399 B.n691 B.n14 585
R400 B.n693 B.n692 585
R401 B.n694 B.n13 585
R402 B.n696 B.n695 585
R403 B.n697 B.n12 585
R404 B.n699 B.n698 585
R405 B.n700 B.n11 585
R406 B.n702 B.n701 585
R407 B.n703 B.n10 585
R408 B.n705 B.n704 585
R409 B.n706 B.n9 585
R410 B.n708 B.n707 585
R411 B.n709 B.n8 585
R412 B.n711 B.n710 585
R413 B.n712 B.n7 585
R414 B.n714 B.n713 585
R415 B.n715 B.n6 585
R416 B.n717 B.n716 585
R417 B.n718 B.n5 585
R418 B.n720 B.n719 585
R419 B.n721 B.n4 585
R420 B.n723 B.n722 585
R421 B.n724 B.n3 585
R422 B.n726 B.n725 585
R423 B.n727 B.n0 585
R424 B.n2 B.n1 585
R425 B.n188 B.n187 585
R426 B.n189 B.n186 585
R427 B.n191 B.n190 585
R428 B.n192 B.n185 585
R429 B.n194 B.n193 585
R430 B.n195 B.n184 585
R431 B.n197 B.n196 585
R432 B.n198 B.n183 585
R433 B.n200 B.n199 585
R434 B.n201 B.n182 585
R435 B.n203 B.n202 585
R436 B.n204 B.n181 585
R437 B.n206 B.n205 585
R438 B.n207 B.n180 585
R439 B.n209 B.n208 585
R440 B.n210 B.n179 585
R441 B.n212 B.n211 585
R442 B.n213 B.n178 585
R443 B.n215 B.n214 585
R444 B.n216 B.n177 585
R445 B.n218 B.n217 585
R446 B.n219 B.n176 585
R447 B.n221 B.n220 585
R448 B.n222 B.n175 585
R449 B.n224 B.n223 585
R450 B.n225 B.n174 585
R451 B.n227 B.n226 585
R452 B.n228 B.n173 585
R453 B.n230 B.n229 585
R454 B.n231 B.n172 585
R455 B.n233 B.n232 585
R456 B.n234 B.n171 585
R457 B.n236 B.n235 585
R458 B.n237 B.n170 585
R459 B.n239 B.n238 585
R460 B.n240 B.n169 585
R461 B.n242 B.n241 585
R462 B.n243 B.n168 585
R463 B.n245 B.n244 585
R464 B.n246 B.n167 585
R465 B.n248 B.n247 585
R466 B.n249 B.n166 585
R467 B.n251 B.n250 585
R468 B.n252 B.n165 585
R469 B.n254 B.n253 585
R470 B.n255 B.n164 585
R471 B.n257 B.n256 585
R472 B.n258 B.n163 585
R473 B.n260 B.n163 530.939
R474 B.n384 B.n121 530.939
R475 B.n534 B.n71 530.939
R476 B.n655 B.n654 530.939
R477 B.n144 B.t3 282.911
R478 B.n326 B.t6 282.911
R479 B.n52 B.t9 282.911
R480 B.n44 B.t0 282.911
R481 B.n729 B.n728 256.663
R482 B.n728 B.n727 235.042
R483 B.n728 B.n2 235.042
R484 B.n326 B.t7 182.41
R485 B.n52 B.t11 182.41
R486 B.n144 B.t4 182.399
R487 B.n44 B.t2 182.399
R488 B.n261 B.n260 163.367
R489 B.n262 B.n261 163.367
R490 B.n262 B.n161 163.367
R491 B.n266 B.n161 163.367
R492 B.n267 B.n266 163.367
R493 B.n268 B.n267 163.367
R494 B.n268 B.n159 163.367
R495 B.n272 B.n159 163.367
R496 B.n273 B.n272 163.367
R497 B.n274 B.n273 163.367
R498 B.n274 B.n157 163.367
R499 B.n278 B.n157 163.367
R500 B.n279 B.n278 163.367
R501 B.n280 B.n279 163.367
R502 B.n280 B.n155 163.367
R503 B.n284 B.n155 163.367
R504 B.n285 B.n284 163.367
R505 B.n286 B.n285 163.367
R506 B.n286 B.n153 163.367
R507 B.n290 B.n153 163.367
R508 B.n291 B.n290 163.367
R509 B.n292 B.n291 163.367
R510 B.n292 B.n151 163.367
R511 B.n296 B.n151 163.367
R512 B.n297 B.n296 163.367
R513 B.n298 B.n297 163.367
R514 B.n298 B.n149 163.367
R515 B.n302 B.n149 163.367
R516 B.n303 B.n302 163.367
R517 B.n304 B.n303 163.367
R518 B.n304 B.n147 163.367
R519 B.n308 B.n147 163.367
R520 B.n309 B.n308 163.367
R521 B.n310 B.n309 163.367
R522 B.n310 B.n143 163.367
R523 B.n315 B.n143 163.367
R524 B.n316 B.n315 163.367
R525 B.n317 B.n316 163.367
R526 B.n317 B.n141 163.367
R527 B.n321 B.n141 163.367
R528 B.n322 B.n321 163.367
R529 B.n323 B.n322 163.367
R530 B.n323 B.n139 163.367
R531 B.n330 B.n139 163.367
R532 B.n331 B.n330 163.367
R533 B.n332 B.n331 163.367
R534 B.n332 B.n137 163.367
R535 B.n336 B.n137 163.367
R536 B.n337 B.n336 163.367
R537 B.n338 B.n337 163.367
R538 B.n338 B.n135 163.367
R539 B.n342 B.n135 163.367
R540 B.n343 B.n342 163.367
R541 B.n344 B.n343 163.367
R542 B.n344 B.n133 163.367
R543 B.n348 B.n133 163.367
R544 B.n349 B.n348 163.367
R545 B.n350 B.n349 163.367
R546 B.n350 B.n131 163.367
R547 B.n354 B.n131 163.367
R548 B.n355 B.n354 163.367
R549 B.n356 B.n355 163.367
R550 B.n356 B.n129 163.367
R551 B.n360 B.n129 163.367
R552 B.n361 B.n360 163.367
R553 B.n362 B.n361 163.367
R554 B.n362 B.n127 163.367
R555 B.n366 B.n127 163.367
R556 B.n367 B.n366 163.367
R557 B.n368 B.n367 163.367
R558 B.n368 B.n125 163.367
R559 B.n372 B.n125 163.367
R560 B.n373 B.n372 163.367
R561 B.n374 B.n373 163.367
R562 B.n374 B.n123 163.367
R563 B.n378 B.n123 163.367
R564 B.n379 B.n378 163.367
R565 B.n380 B.n379 163.367
R566 B.n380 B.n121 163.367
R567 B.n530 B.n71 163.367
R568 B.n530 B.n529 163.367
R569 B.n529 B.n528 163.367
R570 B.n528 B.n73 163.367
R571 B.n524 B.n73 163.367
R572 B.n524 B.n523 163.367
R573 B.n523 B.n522 163.367
R574 B.n522 B.n75 163.367
R575 B.n518 B.n75 163.367
R576 B.n518 B.n517 163.367
R577 B.n517 B.n516 163.367
R578 B.n516 B.n77 163.367
R579 B.n512 B.n77 163.367
R580 B.n512 B.n511 163.367
R581 B.n511 B.n510 163.367
R582 B.n510 B.n79 163.367
R583 B.n506 B.n79 163.367
R584 B.n506 B.n505 163.367
R585 B.n505 B.n504 163.367
R586 B.n504 B.n81 163.367
R587 B.n500 B.n81 163.367
R588 B.n500 B.n499 163.367
R589 B.n499 B.n498 163.367
R590 B.n498 B.n83 163.367
R591 B.n494 B.n83 163.367
R592 B.n494 B.n493 163.367
R593 B.n493 B.n492 163.367
R594 B.n492 B.n85 163.367
R595 B.n488 B.n85 163.367
R596 B.n488 B.n487 163.367
R597 B.n487 B.n486 163.367
R598 B.n486 B.n87 163.367
R599 B.n482 B.n87 163.367
R600 B.n482 B.n481 163.367
R601 B.n481 B.n480 163.367
R602 B.n480 B.n89 163.367
R603 B.n476 B.n89 163.367
R604 B.n476 B.n475 163.367
R605 B.n475 B.n474 163.367
R606 B.n474 B.n91 163.367
R607 B.n470 B.n91 163.367
R608 B.n470 B.n469 163.367
R609 B.n469 B.n468 163.367
R610 B.n468 B.n93 163.367
R611 B.n464 B.n93 163.367
R612 B.n464 B.n463 163.367
R613 B.n463 B.n462 163.367
R614 B.n462 B.n95 163.367
R615 B.n458 B.n95 163.367
R616 B.n458 B.n457 163.367
R617 B.n457 B.n456 163.367
R618 B.n456 B.n97 163.367
R619 B.n452 B.n97 163.367
R620 B.n452 B.n451 163.367
R621 B.n451 B.n450 163.367
R622 B.n450 B.n99 163.367
R623 B.n446 B.n99 163.367
R624 B.n446 B.n445 163.367
R625 B.n445 B.n444 163.367
R626 B.n444 B.n101 163.367
R627 B.n440 B.n101 163.367
R628 B.n440 B.n439 163.367
R629 B.n439 B.n438 163.367
R630 B.n438 B.n103 163.367
R631 B.n434 B.n103 163.367
R632 B.n434 B.n433 163.367
R633 B.n433 B.n432 163.367
R634 B.n432 B.n105 163.367
R635 B.n428 B.n105 163.367
R636 B.n428 B.n427 163.367
R637 B.n427 B.n426 163.367
R638 B.n426 B.n107 163.367
R639 B.n422 B.n107 163.367
R640 B.n422 B.n421 163.367
R641 B.n421 B.n420 163.367
R642 B.n420 B.n109 163.367
R643 B.n416 B.n109 163.367
R644 B.n416 B.n415 163.367
R645 B.n415 B.n414 163.367
R646 B.n414 B.n111 163.367
R647 B.n410 B.n111 163.367
R648 B.n410 B.n409 163.367
R649 B.n409 B.n408 163.367
R650 B.n408 B.n113 163.367
R651 B.n404 B.n113 163.367
R652 B.n404 B.n403 163.367
R653 B.n403 B.n402 163.367
R654 B.n402 B.n115 163.367
R655 B.n398 B.n115 163.367
R656 B.n398 B.n397 163.367
R657 B.n397 B.n396 163.367
R658 B.n396 B.n117 163.367
R659 B.n392 B.n117 163.367
R660 B.n392 B.n391 163.367
R661 B.n391 B.n390 163.367
R662 B.n390 B.n119 163.367
R663 B.n386 B.n119 163.367
R664 B.n386 B.n385 163.367
R665 B.n385 B.n384 163.367
R666 B.n654 B.n27 163.367
R667 B.n650 B.n27 163.367
R668 B.n650 B.n649 163.367
R669 B.n649 B.n648 163.367
R670 B.n648 B.n29 163.367
R671 B.n644 B.n29 163.367
R672 B.n644 B.n643 163.367
R673 B.n643 B.n642 163.367
R674 B.n642 B.n31 163.367
R675 B.n638 B.n31 163.367
R676 B.n638 B.n637 163.367
R677 B.n637 B.n636 163.367
R678 B.n636 B.n33 163.367
R679 B.n632 B.n33 163.367
R680 B.n632 B.n631 163.367
R681 B.n631 B.n630 163.367
R682 B.n630 B.n35 163.367
R683 B.n626 B.n35 163.367
R684 B.n626 B.n625 163.367
R685 B.n625 B.n624 163.367
R686 B.n624 B.n37 163.367
R687 B.n620 B.n37 163.367
R688 B.n620 B.n619 163.367
R689 B.n619 B.n618 163.367
R690 B.n618 B.n39 163.367
R691 B.n614 B.n39 163.367
R692 B.n614 B.n613 163.367
R693 B.n613 B.n612 163.367
R694 B.n612 B.n41 163.367
R695 B.n608 B.n41 163.367
R696 B.n608 B.n607 163.367
R697 B.n607 B.n606 163.367
R698 B.n606 B.n43 163.367
R699 B.n602 B.n43 163.367
R700 B.n602 B.n601 163.367
R701 B.n601 B.n47 163.367
R702 B.n597 B.n47 163.367
R703 B.n597 B.n596 163.367
R704 B.n596 B.n595 163.367
R705 B.n595 B.n49 163.367
R706 B.n591 B.n49 163.367
R707 B.n591 B.n590 163.367
R708 B.n590 B.n589 163.367
R709 B.n589 B.n51 163.367
R710 B.n584 B.n51 163.367
R711 B.n584 B.n583 163.367
R712 B.n583 B.n582 163.367
R713 B.n582 B.n55 163.367
R714 B.n578 B.n55 163.367
R715 B.n578 B.n577 163.367
R716 B.n577 B.n576 163.367
R717 B.n576 B.n57 163.367
R718 B.n572 B.n57 163.367
R719 B.n572 B.n571 163.367
R720 B.n571 B.n570 163.367
R721 B.n570 B.n59 163.367
R722 B.n566 B.n59 163.367
R723 B.n566 B.n565 163.367
R724 B.n565 B.n564 163.367
R725 B.n564 B.n61 163.367
R726 B.n560 B.n61 163.367
R727 B.n560 B.n559 163.367
R728 B.n559 B.n558 163.367
R729 B.n558 B.n63 163.367
R730 B.n554 B.n63 163.367
R731 B.n554 B.n553 163.367
R732 B.n553 B.n552 163.367
R733 B.n552 B.n65 163.367
R734 B.n548 B.n65 163.367
R735 B.n548 B.n547 163.367
R736 B.n547 B.n546 163.367
R737 B.n546 B.n67 163.367
R738 B.n542 B.n67 163.367
R739 B.n542 B.n541 163.367
R740 B.n541 B.n540 163.367
R741 B.n540 B.n69 163.367
R742 B.n536 B.n69 163.367
R743 B.n536 B.n535 163.367
R744 B.n535 B.n534 163.367
R745 B.n656 B.n655 163.367
R746 B.n656 B.n25 163.367
R747 B.n660 B.n25 163.367
R748 B.n661 B.n660 163.367
R749 B.n662 B.n661 163.367
R750 B.n662 B.n23 163.367
R751 B.n666 B.n23 163.367
R752 B.n667 B.n666 163.367
R753 B.n668 B.n667 163.367
R754 B.n668 B.n21 163.367
R755 B.n672 B.n21 163.367
R756 B.n673 B.n672 163.367
R757 B.n674 B.n673 163.367
R758 B.n674 B.n19 163.367
R759 B.n678 B.n19 163.367
R760 B.n679 B.n678 163.367
R761 B.n680 B.n679 163.367
R762 B.n680 B.n17 163.367
R763 B.n684 B.n17 163.367
R764 B.n685 B.n684 163.367
R765 B.n686 B.n685 163.367
R766 B.n686 B.n15 163.367
R767 B.n690 B.n15 163.367
R768 B.n691 B.n690 163.367
R769 B.n692 B.n691 163.367
R770 B.n692 B.n13 163.367
R771 B.n696 B.n13 163.367
R772 B.n697 B.n696 163.367
R773 B.n698 B.n697 163.367
R774 B.n698 B.n11 163.367
R775 B.n702 B.n11 163.367
R776 B.n703 B.n702 163.367
R777 B.n704 B.n703 163.367
R778 B.n704 B.n9 163.367
R779 B.n708 B.n9 163.367
R780 B.n709 B.n708 163.367
R781 B.n710 B.n709 163.367
R782 B.n710 B.n7 163.367
R783 B.n714 B.n7 163.367
R784 B.n715 B.n714 163.367
R785 B.n716 B.n715 163.367
R786 B.n716 B.n5 163.367
R787 B.n720 B.n5 163.367
R788 B.n721 B.n720 163.367
R789 B.n722 B.n721 163.367
R790 B.n722 B.n3 163.367
R791 B.n726 B.n3 163.367
R792 B.n727 B.n726 163.367
R793 B.n188 B.n2 163.367
R794 B.n189 B.n188 163.367
R795 B.n190 B.n189 163.367
R796 B.n190 B.n185 163.367
R797 B.n194 B.n185 163.367
R798 B.n195 B.n194 163.367
R799 B.n196 B.n195 163.367
R800 B.n196 B.n183 163.367
R801 B.n200 B.n183 163.367
R802 B.n201 B.n200 163.367
R803 B.n202 B.n201 163.367
R804 B.n202 B.n181 163.367
R805 B.n206 B.n181 163.367
R806 B.n207 B.n206 163.367
R807 B.n208 B.n207 163.367
R808 B.n208 B.n179 163.367
R809 B.n212 B.n179 163.367
R810 B.n213 B.n212 163.367
R811 B.n214 B.n213 163.367
R812 B.n214 B.n177 163.367
R813 B.n218 B.n177 163.367
R814 B.n219 B.n218 163.367
R815 B.n220 B.n219 163.367
R816 B.n220 B.n175 163.367
R817 B.n224 B.n175 163.367
R818 B.n225 B.n224 163.367
R819 B.n226 B.n225 163.367
R820 B.n226 B.n173 163.367
R821 B.n230 B.n173 163.367
R822 B.n231 B.n230 163.367
R823 B.n232 B.n231 163.367
R824 B.n232 B.n171 163.367
R825 B.n236 B.n171 163.367
R826 B.n237 B.n236 163.367
R827 B.n238 B.n237 163.367
R828 B.n238 B.n169 163.367
R829 B.n242 B.n169 163.367
R830 B.n243 B.n242 163.367
R831 B.n244 B.n243 163.367
R832 B.n244 B.n167 163.367
R833 B.n248 B.n167 163.367
R834 B.n249 B.n248 163.367
R835 B.n250 B.n249 163.367
R836 B.n250 B.n165 163.367
R837 B.n254 B.n165 163.367
R838 B.n255 B.n254 163.367
R839 B.n256 B.n255 163.367
R840 B.n256 B.n163 163.367
R841 B.n327 B.t8 113.948
R842 B.n53 B.t10 113.948
R843 B.n145 B.t5 113.938
R844 B.n45 B.t1 113.938
R845 B.n145 B.n144 68.4611
R846 B.n327 B.n326 68.4611
R847 B.n53 B.n52 68.4611
R848 B.n45 B.n44 68.4611
R849 B.n312 B.n145 59.5399
R850 B.n328 B.n327 59.5399
R851 B.n586 B.n53 59.5399
R852 B.n46 B.n45 59.5399
R853 B.n653 B.n26 34.4981
R854 B.n533 B.n532 34.4981
R855 B.n383 B.n382 34.4981
R856 B.n259 B.n258 34.4981
R857 B B.n729 18.0485
R858 B.n657 B.n26 10.6151
R859 B.n658 B.n657 10.6151
R860 B.n659 B.n658 10.6151
R861 B.n659 B.n24 10.6151
R862 B.n663 B.n24 10.6151
R863 B.n664 B.n663 10.6151
R864 B.n665 B.n664 10.6151
R865 B.n665 B.n22 10.6151
R866 B.n669 B.n22 10.6151
R867 B.n670 B.n669 10.6151
R868 B.n671 B.n670 10.6151
R869 B.n671 B.n20 10.6151
R870 B.n675 B.n20 10.6151
R871 B.n676 B.n675 10.6151
R872 B.n677 B.n676 10.6151
R873 B.n677 B.n18 10.6151
R874 B.n681 B.n18 10.6151
R875 B.n682 B.n681 10.6151
R876 B.n683 B.n682 10.6151
R877 B.n683 B.n16 10.6151
R878 B.n687 B.n16 10.6151
R879 B.n688 B.n687 10.6151
R880 B.n689 B.n688 10.6151
R881 B.n689 B.n14 10.6151
R882 B.n693 B.n14 10.6151
R883 B.n694 B.n693 10.6151
R884 B.n695 B.n694 10.6151
R885 B.n695 B.n12 10.6151
R886 B.n699 B.n12 10.6151
R887 B.n700 B.n699 10.6151
R888 B.n701 B.n700 10.6151
R889 B.n701 B.n10 10.6151
R890 B.n705 B.n10 10.6151
R891 B.n706 B.n705 10.6151
R892 B.n707 B.n706 10.6151
R893 B.n707 B.n8 10.6151
R894 B.n711 B.n8 10.6151
R895 B.n712 B.n711 10.6151
R896 B.n713 B.n712 10.6151
R897 B.n713 B.n6 10.6151
R898 B.n717 B.n6 10.6151
R899 B.n718 B.n717 10.6151
R900 B.n719 B.n718 10.6151
R901 B.n719 B.n4 10.6151
R902 B.n723 B.n4 10.6151
R903 B.n724 B.n723 10.6151
R904 B.n725 B.n724 10.6151
R905 B.n725 B.n0 10.6151
R906 B.n653 B.n652 10.6151
R907 B.n652 B.n651 10.6151
R908 B.n651 B.n28 10.6151
R909 B.n647 B.n28 10.6151
R910 B.n647 B.n646 10.6151
R911 B.n646 B.n645 10.6151
R912 B.n645 B.n30 10.6151
R913 B.n641 B.n30 10.6151
R914 B.n641 B.n640 10.6151
R915 B.n640 B.n639 10.6151
R916 B.n639 B.n32 10.6151
R917 B.n635 B.n32 10.6151
R918 B.n635 B.n634 10.6151
R919 B.n634 B.n633 10.6151
R920 B.n633 B.n34 10.6151
R921 B.n629 B.n34 10.6151
R922 B.n629 B.n628 10.6151
R923 B.n628 B.n627 10.6151
R924 B.n627 B.n36 10.6151
R925 B.n623 B.n36 10.6151
R926 B.n623 B.n622 10.6151
R927 B.n622 B.n621 10.6151
R928 B.n621 B.n38 10.6151
R929 B.n617 B.n38 10.6151
R930 B.n617 B.n616 10.6151
R931 B.n616 B.n615 10.6151
R932 B.n615 B.n40 10.6151
R933 B.n611 B.n40 10.6151
R934 B.n611 B.n610 10.6151
R935 B.n610 B.n609 10.6151
R936 B.n609 B.n42 10.6151
R937 B.n605 B.n42 10.6151
R938 B.n605 B.n604 10.6151
R939 B.n604 B.n603 10.6151
R940 B.n600 B.n599 10.6151
R941 B.n599 B.n598 10.6151
R942 B.n598 B.n48 10.6151
R943 B.n594 B.n48 10.6151
R944 B.n594 B.n593 10.6151
R945 B.n593 B.n592 10.6151
R946 B.n592 B.n50 10.6151
R947 B.n588 B.n50 10.6151
R948 B.n588 B.n587 10.6151
R949 B.n585 B.n54 10.6151
R950 B.n581 B.n54 10.6151
R951 B.n581 B.n580 10.6151
R952 B.n580 B.n579 10.6151
R953 B.n579 B.n56 10.6151
R954 B.n575 B.n56 10.6151
R955 B.n575 B.n574 10.6151
R956 B.n574 B.n573 10.6151
R957 B.n573 B.n58 10.6151
R958 B.n569 B.n58 10.6151
R959 B.n569 B.n568 10.6151
R960 B.n568 B.n567 10.6151
R961 B.n567 B.n60 10.6151
R962 B.n563 B.n60 10.6151
R963 B.n563 B.n562 10.6151
R964 B.n562 B.n561 10.6151
R965 B.n561 B.n62 10.6151
R966 B.n557 B.n62 10.6151
R967 B.n557 B.n556 10.6151
R968 B.n556 B.n555 10.6151
R969 B.n555 B.n64 10.6151
R970 B.n551 B.n64 10.6151
R971 B.n551 B.n550 10.6151
R972 B.n550 B.n549 10.6151
R973 B.n549 B.n66 10.6151
R974 B.n545 B.n66 10.6151
R975 B.n545 B.n544 10.6151
R976 B.n544 B.n543 10.6151
R977 B.n543 B.n68 10.6151
R978 B.n539 B.n68 10.6151
R979 B.n539 B.n538 10.6151
R980 B.n538 B.n537 10.6151
R981 B.n537 B.n70 10.6151
R982 B.n533 B.n70 10.6151
R983 B.n532 B.n531 10.6151
R984 B.n531 B.n72 10.6151
R985 B.n527 B.n72 10.6151
R986 B.n527 B.n526 10.6151
R987 B.n526 B.n525 10.6151
R988 B.n525 B.n74 10.6151
R989 B.n521 B.n74 10.6151
R990 B.n521 B.n520 10.6151
R991 B.n520 B.n519 10.6151
R992 B.n519 B.n76 10.6151
R993 B.n515 B.n76 10.6151
R994 B.n515 B.n514 10.6151
R995 B.n514 B.n513 10.6151
R996 B.n513 B.n78 10.6151
R997 B.n509 B.n78 10.6151
R998 B.n509 B.n508 10.6151
R999 B.n508 B.n507 10.6151
R1000 B.n507 B.n80 10.6151
R1001 B.n503 B.n80 10.6151
R1002 B.n503 B.n502 10.6151
R1003 B.n502 B.n501 10.6151
R1004 B.n501 B.n82 10.6151
R1005 B.n497 B.n82 10.6151
R1006 B.n497 B.n496 10.6151
R1007 B.n496 B.n495 10.6151
R1008 B.n495 B.n84 10.6151
R1009 B.n491 B.n84 10.6151
R1010 B.n491 B.n490 10.6151
R1011 B.n490 B.n489 10.6151
R1012 B.n489 B.n86 10.6151
R1013 B.n485 B.n86 10.6151
R1014 B.n485 B.n484 10.6151
R1015 B.n484 B.n483 10.6151
R1016 B.n483 B.n88 10.6151
R1017 B.n479 B.n88 10.6151
R1018 B.n479 B.n478 10.6151
R1019 B.n478 B.n477 10.6151
R1020 B.n477 B.n90 10.6151
R1021 B.n473 B.n90 10.6151
R1022 B.n473 B.n472 10.6151
R1023 B.n472 B.n471 10.6151
R1024 B.n471 B.n92 10.6151
R1025 B.n467 B.n92 10.6151
R1026 B.n467 B.n466 10.6151
R1027 B.n466 B.n465 10.6151
R1028 B.n465 B.n94 10.6151
R1029 B.n461 B.n94 10.6151
R1030 B.n461 B.n460 10.6151
R1031 B.n460 B.n459 10.6151
R1032 B.n459 B.n96 10.6151
R1033 B.n455 B.n96 10.6151
R1034 B.n455 B.n454 10.6151
R1035 B.n454 B.n453 10.6151
R1036 B.n453 B.n98 10.6151
R1037 B.n449 B.n98 10.6151
R1038 B.n449 B.n448 10.6151
R1039 B.n448 B.n447 10.6151
R1040 B.n447 B.n100 10.6151
R1041 B.n443 B.n100 10.6151
R1042 B.n443 B.n442 10.6151
R1043 B.n442 B.n441 10.6151
R1044 B.n441 B.n102 10.6151
R1045 B.n437 B.n102 10.6151
R1046 B.n437 B.n436 10.6151
R1047 B.n436 B.n435 10.6151
R1048 B.n435 B.n104 10.6151
R1049 B.n431 B.n104 10.6151
R1050 B.n431 B.n430 10.6151
R1051 B.n430 B.n429 10.6151
R1052 B.n429 B.n106 10.6151
R1053 B.n425 B.n106 10.6151
R1054 B.n425 B.n424 10.6151
R1055 B.n424 B.n423 10.6151
R1056 B.n423 B.n108 10.6151
R1057 B.n419 B.n108 10.6151
R1058 B.n419 B.n418 10.6151
R1059 B.n418 B.n417 10.6151
R1060 B.n417 B.n110 10.6151
R1061 B.n413 B.n110 10.6151
R1062 B.n413 B.n412 10.6151
R1063 B.n412 B.n411 10.6151
R1064 B.n411 B.n112 10.6151
R1065 B.n407 B.n112 10.6151
R1066 B.n407 B.n406 10.6151
R1067 B.n406 B.n405 10.6151
R1068 B.n405 B.n114 10.6151
R1069 B.n401 B.n114 10.6151
R1070 B.n401 B.n400 10.6151
R1071 B.n400 B.n399 10.6151
R1072 B.n399 B.n116 10.6151
R1073 B.n395 B.n116 10.6151
R1074 B.n395 B.n394 10.6151
R1075 B.n394 B.n393 10.6151
R1076 B.n393 B.n118 10.6151
R1077 B.n389 B.n118 10.6151
R1078 B.n389 B.n388 10.6151
R1079 B.n388 B.n387 10.6151
R1080 B.n387 B.n120 10.6151
R1081 B.n383 B.n120 10.6151
R1082 B.n187 B.n1 10.6151
R1083 B.n187 B.n186 10.6151
R1084 B.n191 B.n186 10.6151
R1085 B.n192 B.n191 10.6151
R1086 B.n193 B.n192 10.6151
R1087 B.n193 B.n184 10.6151
R1088 B.n197 B.n184 10.6151
R1089 B.n198 B.n197 10.6151
R1090 B.n199 B.n198 10.6151
R1091 B.n199 B.n182 10.6151
R1092 B.n203 B.n182 10.6151
R1093 B.n204 B.n203 10.6151
R1094 B.n205 B.n204 10.6151
R1095 B.n205 B.n180 10.6151
R1096 B.n209 B.n180 10.6151
R1097 B.n210 B.n209 10.6151
R1098 B.n211 B.n210 10.6151
R1099 B.n211 B.n178 10.6151
R1100 B.n215 B.n178 10.6151
R1101 B.n216 B.n215 10.6151
R1102 B.n217 B.n216 10.6151
R1103 B.n217 B.n176 10.6151
R1104 B.n221 B.n176 10.6151
R1105 B.n222 B.n221 10.6151
R1106 B.n223 B.n222 10.6151
R1107 B.n223 B.n174 10.6151
R1108 B.n227 B.n174 10.6151
R1109 B.n228 B.n227 10.6151
R1110 B.n229 B.n228 10.6151
R1111 B.n229 B.n172 10.6151
R1112 B.n233 B.n172 10.6151
R1113 B.n234 B.n233 10.6151
R1114 B.n235 B.n234 10.6151
R1115 B.n235 B.n170 10.6151
R1116 B.n239 B.n170 10.6151
R1117 B.n240 B.n239 10.6151
R1118 B.n241 B.n240 10.6151
R1119 B.n241 B.n168 10.6151
R1120 B.n245 B.n168 10.6151
R1121 B.n246 B.n245 10.6151
R1122 B.n247 B.n246 10.6151
R1123 B.n247 B.n166 10.6151
R1124 B.n251 B.n166 10.6151
R1125 B.n252 B.n251 10.6151
R1126 B.n253 B.n252 10.6151
R1127 B.n253 B.n164 10.6151
R1128 B.n257 B.n164 10.6151
R1129 B.n258 B.n257 10.6151
R1130 B.n259 B.n162 10.6151
R1131 B.n263 B.n162 10.6151
R1132 B.n264 B.n263 10.6151
R1133 B.n265 B.n264 10.6151
R1134 B.n265 B.n160 10.6151
R1135 B.n269 B.n160 10.6151
R1136 B.n270 B.n269 10.6151
R1137 B.n271 B.n270 10.6151
R1138 B.n271 B.n158 10.6151
R1139 B.n275 B.n158 10.6151
R1140 B.n276 B.n275 10.6151
R1141 B.n277 B.n276 10.6151
R1142 B.n277 B.n156 10.6151
R1143 B.n281 B.n156 10.6151
R1144 B.n282 B.n281 10.6151
R1145 B.n283 B.n282 10.6151
R1146 B.n283 B.n154 10.6151
R1147 B.n287 B.n154 10.6151
R1148 B.n288 B.n287 10.6151
R1149 B.n289 B.n288 10.6151
R1150 B.n289 B.n152 10.6151
R1151 B.n293 B.n152 10.6151
R1152 B.n294 B.n293 10.6151
R1153 B.n295 B.n294 10.6151
R1154 B.n295 B.n150 10.6151
R1155 B.n299 B.n150 10.6151
R1156 B.n300 B.n299 10.6151
R1157 B.n301 B.n300 10.6151
R1158 B.n301 B.n148 10.6151
R1159 B.n305 B.n148 10.6151
R1160 B.n306 B.n305 10.6151
R1161 B.n307 B.n306 10.6151
R1162 B.n307 B.n146 10.6151
R1163 B.n311 B.n146 10.6151
R1164 B.n314 B.n313 10.6151
R1165 B.n314 B.n142 10.6151
R1166 B.n318 B.n142 10.6151
R1167 B.n319 B.n318 10.6151
R1168 B.n320 B.n319 10.6151
R1169 B.n320 B.n140 10.6151
R1170 B.n324 B.n140 10.6151
R1171 B.n325 B.n324 10.6151
R1172 B.n329 B.n325 10.6151
R1173 B.n333 B.n138 10.6151
R1174 B.n334 B.n333 10.6151
R1175 B.n335 B.n334 10.6151
R1176 B.n335 B.n136 10.6151
R1177 B.n339 B.n136 10.6151
R1178 B.n340 B.n339 10.6151
R1179 B.n341 B.n340 10.6151
R1180 B.n341 B.n134 10.6151
R1181 B.n345 B.n134 10.6151
R1182 B.n346 B.n345 10.6151
R1183 B.n347 B.n346 10.6151
R1184 B.n347 B.n132 10.6151
R1185 B.n351 B.n132 10.6151
R1186 B.n352 B.n351 10.6151
R1187 B.n353 B.n352 10.6151
R1188 B.n353 B.n130 10.6151
R1189 B.n357 B.n130 10.6151
R1190 B.n358 B.n357 10.6151
R1191 B.n359 B.n358 10.6151
R1192 B.n359 B.n128 10.6151
R1193 B.n363 B.n128 10.6151
R1194 B.n364 B.n363 10.6151
R1195 B.n365 B.n364 10.6151
R1196 B.n365 B.n126 10.6151
R1197 B.n369 B.n126 10.6151
R1198 B.n370 B.n369 10.6151
R1199 B.n371 B.n370 10.6151
R1200 B.n371 B.n124 10.6151
R1201 B.n375 B.n124 10.6151
R1202 B.n376 B.n375 10.6151
R1203 B.n377 B.n376 10.6151
R1204 B.n377 B.n122 10.6151
R1205 B.n381 B.n122 10.6151
R1206 B.n382 B.n381 10.6151
R1207 B.n603 B.n46 9.36635
R1208 B.n586 B.n585 9.36635
R1209 B.n312 B.n311 9.36635
R1210 B.n328 B.n138 9.36635
R1211 B.n729 B.n0 8.11757
R1212 B.n729 B.n1 8.11757
R1213 B.n600 B.n46 1.24928
R1214 B.n587 B.n586 1.24928
R1215 B.n313 B.n312 1.24928
R1216 B.n329 B.n328 1.24928
R1217 VN.n34 VN.n33 161.3
R1218 VN.n32 VN.n19 161.3
R1219 VN.n31 VN.n30 161.3
R1220 VN.n29 VN.n20 161.3
R1221 VN.n28 VN.n27 161.3
R1222 VN.n26 VN.n21 161.3
R1223 VN.n25 VN.n24 161.3
R1224 VN.n16 VN.n15 161.3
R1225 VN.n14 VN.n1 161.3
R1226 VN.n13 VN.n12 161.3
R1227 VN.n11 VN.n2 161.3
R1228 VN.n10 VN.n9 161.3
R1229 VN.n8 VN.n3 161.3
R1230 VN.n7 VN.n6 161.3
R1231 VN.n23 VN.t0 107.028
R1232 VN.n5 VN.t5 107.028
R1233 VN.n17 VN.n0 76.4741
R1234 VN.n35 VN.n18 76.4741
R1235 VN.n4 VN.t3 74.108
R1236 VN.n0 VN.t4 74.108
R1237 VN.n22 VN.t1 74.108
R1238 VN.n18 VN.t2 74.108
R1239 VN.n5 VN.n4 62.2079
R1240 VN.n23 VN.n22 62.2079
R1241 VN VN.n35 49.6307
R1242 VN.n13 VN.n2 42.0302
R1243 VN.n31 VN.n20 42.0302
R1244 VN.n9 VN.n2 39.1239
R1245 VN.n27 VN.n20 39.1239
R1246 VN.n8 VN.n7 24.5923
R1247 VN.n9 VN.n8 24.5923
R1248 VN.n14 VN.n13 24.5923
R1249 VN.n15 VN.n14 24.5923
R1250 VN.n27 VN.n26 24.5923
R1251 VN.n26 VN.n25 24.5923
R1252 VN.n33 VN.n32 24.5923
R1253 VN.n32 VN.n31 24.5923
R1254 VN.n15 VN.n0 13.7719
R1255 VN.n33 VN.n18 13.7719
R1256 VN.n7 VN.n4 12.2964
R1257 VN.n25 VN.n22 12.2964
R1258 VN.n24 VN.n23 4.19127
R1259 VN.n6 VN.n5 4.19127
R1260 VN.n35 VN.n34 0.354861
R1261 VN.n17 VN.n16 0.354861
R1262 VN VN.n17 0.267071
R1263 VN.n34 VN.n19 0.189894
R1264 VN.n30 VN.n19 0.189894
R1265 VN.n30 VN.n29 0.189894
R1266 VN.n29 VN.n28 0.189894
R1267 VN.n28 VN.n21 0.189894
R1268 VN.n24 VN.n21 0.189894
R1269 VN.n6 VN.n3 0.189894
R1270 VN.n10 VN.n3 0.189894
R1271 VN.n11 VN.n10 0.189894
R1272 VN.n12 VN.n11 0.189894
R1273 VN.n12 VN.n1 0.189894
R1274 VN.n16 VN.n1 0.189894
R1275 VDD2.n1 VDD2.t0 81.394
R1276 VDD2.n2 VDD2.t3 79.1673
R1277 VDD2.n1 VDD2.n0 76.5691
R1278 VDD2 VDD2.n3 76.5665
R1279 VDD2.n2 VDD2.n1 42.0881
R1280 VDD2.n3 VDD2.t4 3.30385
R1281 VDD2.n3 VDD2.t5 3.30385
R1282 VDD2.n0 VDD2.t2 3.30385
R1283 VDD2.n0 VDD2.t1 3.30385
R1284 VDD2 VDD2.n2 2.34102
C0 B VTAIL 3.42433f
C1 w_n3794_n2936# VDD1 2.28527f
C2 VP VDD2 0.509197f
C3 VDD1 VTAIL 7.17153f
C4 VP VN 7.107419f
C5 VP B 2.09746f
C6 w_n3794_n2936# VTAIL 2.72407f
C7 VP VDD1 6.14527f
C8 VN VDD2 5.79055f
C9 B VDD2 2.16556f
C10 VP w_n3794_n2936# 7.78738f
C11 B VN 1.27268f
C12 VP VTAIL 6.20844f
C13 VDD2 VDD1 1.63951f
C14 VN VDD1 0.151709f
C15 w_n3794_n2936# VDD2 2.38951f
C16 B VDD1 2.07708f
C17 w_n3794_n2936# VN 7.29519f
C18 B w_n3794_n2936# 9.89934f
C19 VDD2 VTAIL 7.22734f
C20 VN VTAIL 6.19422f
C21 VDD2 VSUBS 2.037315f
C22 VDD1 VSUBS 2.56265f
C23 VTAIL VSUBS 1.233783f
C24 VN VSUBS 6.36739f
C25 VP VSUBS 3.330145f
C26 B VSUBS 5.049342f
C27 w_n3794_n2936# VSUBS 0.137631p
C28 VDD2.t0 VSUBS 2.23115f
C29 VDD2.t2 VSUBS 0.225921f
C30 VDD2.t1 VSUBS 0.225921f
C31 VDD2.n0 VSUBS 1.68636f
C32 VDD2.n1 VSUBS 4.1393f
C33 VDD2.t3 VSUBS 2.20784f
C34 VDD2.n2 VSUBS 3.5608f
C35 VDD2.t4 VSUBS 0.225921f
C36 VDD2.t5 VSUBS 0.225921f
C37 VDD2.n3 VSUBS 1.68632f
C38 VN.t4 VSUBS 2.48171f
C39 VN.n0 VSUBS 0.991817f
C40 VN.n1 VSUBS 0.029109f
C41 VN.n2 VSUBS 0.023594f
C42 VN.n3 VSUBS 0.029109f
C43 VN.t3 VSUBS 2.48171f
C44 VN.n4 VSUBS 0.978054f
C45 VN.t5 VSUBS 2.81545f
C46 VN.n5 VSUBS 0.930415f
C47 VN.n6 VSUBS 0.338787f
C48 VN.n7 VSUBS 0.040656f
C49 VN.n8 VSUBS 0.05398f
C50 VN.n9 VSUBS 0.05794f
C51 VN.n10 VSUBS 0.029109f
C52 VN.n11 VSUBS 0.029109f
C53 VN.n12 VSUBS 0.029109f
C54 VN.n13 VSUBS 0.057076f
C55 VN.n14 VSUBS 0.05398f
C56 VN.n15 VSUBS 0.042255f
C57 VN.n16 VSUBS 0.046974f
C58 VN.n17 VSUBS 0.070259f
C59 VN.t2 VSUBS 2.48171f
C60 VN.n18 VSUBS 0.991817f
C61 VN.n19 VSUBS 0.029109f
C62 VN.n20 VSUBS 0.023594f
C63 VN.n21 VSUBS 0.029109f
C64 VN.t1 VSUBS 2.48171f
C65 VN.n22 VSUBS 0.978054f
C66 VN.t0 VSUBS 2.81545f
C67 VN.n23 VSUBS 0.930415f
C68 VN.n24 VSUBS 0.338787f
C69 VN.n25 VSUBS 0.040656f
C70 VN.n26 VSUBS 0.05398f
C71 VN.n27 VSUBS 0.05794f
C72 VN.n28 VSUBS 0.029109f
C73 VN.n29 VSUBS 0.029109f
C74 VN.n30 VSUBS 0.029109f
C75 VN.n31 VSUBS 0.057076f
C76 VN.n32 VSUBS 0.05398f
C77 VN.n33 VSUBS 0.042255f
C78 VN.n34 VSUBS 0.046974f
C79 VN.n35 VSUBS 1.64095f
C80 B.n0 VSUBS 0.00823f
C81 B.n1 VSUBS 0.00823f
C82 B.n2 VSUBS 0.012171f
C83 B.n3 VSUBS 0.009327f
C84 B.n4 VSUBS 0.009327f
C85 B.n5 VSUBS 0.009327f
C86 B.n6 VSUBS 0.009327f
C87 B.n7 VSUBS 0.009327f
C88 B.n8 VSUBS 0.009327f
C89 B.n9 VSUBS 0.009327f
C90 B.n10 VSUBS 0.009327f
C91 B.n11 VSUBS 0.009327f
C92 B.n12 VSUBS 0.009327f
C93 B.n13 VSUBS 0.009327f
C94 B.n14 VSUBS 0.009327f
C95 B.n15 VSUBS 0.009327f
C96 B.n16 VSUBS 0.009327f
C97 B.n17 VSUBS 0.009327f
C98 B.n18 VSUBS 0.009327f
C99 B.n19 VSUBS 0.009327f
C100 B.n20 VSUBS 0.009327f
C101 B.n21 VSUBS 0.009327f
C102 B.n22 VSUBS 0.009327f
C103 B.n23 VSUBS 0.009327f
C104 B.n24 VSUBS 0.009327f
C105 B.n25 VSUBS 0.009327f
C106 B.n26 VSUBS 0.022059f
C107 B.n27 VSUBS 0.009327f
C108 B.n28 VSUBS 0.009327f
C109 B.n29 VSUBS 0.009327f
C110 B.n30 VSUBS 0.009327f
C111 B.n31 VSUBS 0.009327f
C112 B.n32 VSUBS 0.009327f
C113 B.n33 VSUBS 0.009327f
C114 B.n34 VSUBS 0.009327f
C115 B.n35 VSUBS 0.009327f
C116 B.n36 VSUBS 0.009327f
C117 B.n37 VSUBS 0.009327f
C118 B.n38 VSUBS 0.009327f
C119 B.n39 VSUBS 0.009327f
C120 B.n40 VSUBS 0.009327f
C121 B.n41 VSUBS 0.009327f
C122 B.n42 VSUBS 0.009327f
C123 B.n43 VSUBS 0.009327f
C124 B.t1 VSUBS 0.417208f
C125 B.t2 VSUBS 0.449291f
C126 B.t0 VSUBS 1.958f
C127 B.n44 VSUBS 0.248488f
C128 B.n45 VSUBS 0.098782f
C129 B.n46 VSUBS 0.02161f
C130 B.n47 VSUBS 0.009327f
C131 B.n48 VSUBS 0.009327f
C132 B.n49 VSUBS 0.009327f
C133 B.n50 VSUBS 0.009327f
C134 B.n51 VSUBS 0.009327f
C135 B.t10 VSUBS 0.417203f
C136 B.t11 VSUBS 0.449286f
C137 B.t9 VSUBS 1.958f
C138 B.n52 VSUBS 0.248493f
C139 B.n53 VSUBS 0.098787f
C140 B.n54 VSUBS 0.009327f
C141 B.n55 VSUBS 0.009327f
C142 B.n56 VSUBS 0.009327f
C143 B.n57 VSUBS 0.009327f
C144 B.n58 VSUBS 0.009327f
C145 B.n59 VSUBS 0.009327f
C146 B.n60 VSUBS 0.009327f
C147 B.n61 VSUBS 0.009327f
C148 B.n62 VSUBS 0.009327f
C149 B.n63 VSUBS 0.009327f
C150 B.n64 VSUBS 0.009327f
C151 B.n65 VSUBS 0.009327f
C152 B.n66 VSUBS 0.009327f
C153 B.n67 VSUBS 0.009327f
C154 B.n68 VSUBS 0.009327f
C155 B.n69 VSUBS 0.009327f
C156 B.n70 VSUBS 0.009327f
C157 B.n71 VSUBS 0.022059f
C158 B.n72 VSUBS 0.009327f
C159 B.n73 VSUBS 0.009327f
C160 B.n74 VSUBS 0.009327f
C161 B.n75 VSUBS 0.009327f
C162 B.n76 VSUBS 0.009327f
C163 B.n77 VSUBS 0.009327f
C164 B.n78 VSUBS 0.009327f
C165 B.n79 VSUBS 0.009327f
C166 B.n80 VSUBS 0.009327f
C167 B.n81 VSUBS 0.009327f
C168 B.n82 VSUBS 0.009327f
C169 B.n83 VSUBS 0.009327f
C170 B.n84 VSUBS 0.009327f
C171 B.n85 VSUBS 0.009327f
C172 B.n86 VSUBS 0.009327f
C173 B.n87 VSUBS 0.009327f
C174 B.n88 VSUBS 0.009327f
C175 B.n89 VSUBS 0.009327f
C176 B.n90 VSUBS 0.009327f
C177 B.n91 VSUBS 0.009327f
C178 B.n92 VSUBS 0.009327f
C179 B.n93 VSUBS 0.009327f
C180 B.n94 VSUBS 0.009327f
C181 B.n95 VSUBS 0.009327f
C182 B.n96 VSUBS 0.009327f
C183 B.n97 VSUBS 0.009327f
C184 B.n98 VSUBS 0.009327f
C185 B.n99 VSUBS 0.009327f
C186 B.n100 VSUBS 0.009327f
C187 B.n101 VSUBS 0.009327f
C188 B.n102 VSUBS 0.009327f
C189 B.n103 VSUBS 0.009327f
C190 B.n104 VSUBS 0.009327f
C191 B.n105 VSUBS 0.009327f
C192 B.n106 VSUBS 0.009327f
C193 B.n107 VSUBS 0.009327f
C194 B.n108 VSUBS 0.009327f
C195 B.n109 VSUBS 0.009327f
C196 B.n110 VSUBS 0.009327f
C197 B.n111 VSUBS 0.009327f
C198 B.n112 VSUBS 0.009327f
C199 B.n113 VSUBS 0.009327f
C200 B.n114 VSUBS 0.009327f
C201 B.n115 VSUBS 0.009327f
C202 B.n116 VSUBS 0.009327f
C203 B.n117 VSUBS 0.009327f
C204 B.n118 VSUBS 0.009327f
C205 B.n119 VSUBS 0.009327f
C206 B.n120 VSUBS 0.009327f
C207 B.n121 VSUBS 0.023205f
C208 B.n122 VSUBS 0.009327f
C209 B.n123 VSUBS 0.009327f
C210 B.n124 VSUBS 0.009327f
C211 B.n125 VSUBS 0.009327f
C212 B.n126 VSUBS 0.009327f
C213 B.n127 VSUBS 0.009327f
C214 B.n128 VSUBS 0.009327f
C215 B.n129 VSUBS 0.009327f
C216 B.n130 VSUBS 0.009327f
C217 B.n131 VSUBS 0.009327f
C218 B.n132 VSUBS 0.009327f
C219 B.n133 VSUBS 0.009327f
C220 B.n134 VSUBS 0.009327f
C221 B.n135 VSUBS 0.009327f
C222 B.n136 VSUBS 0.009327f
C223 B.n137 VSUBS 0.009327f
C224 B.n138 VSUBS 0.008778f
C225 B.n139 VSUBS 0.009327f
C226 B.n140 VSUBS 0.009327f
C227 B.n141 VSUBS 0.009327f
C228 B.n142 VSUBS 0.009327f
C229 B.n143 VSUBS 0.009327f
C230 B.t5 VSUBS 0.417208f
C231 B.t4 VSUBS 0.449291f
C232 B.t3 VSUBS 1.958f
C233 B.n144 VSUBS 0.248488f
C234 B.n145 VSUBS 0.098782f
C235 B.n146 VSUBS 0.009327f
C236 B.n147 VSUBS 0.009327f
C237 B.n148 VSUBS 0.009327f
C238 B.n149 VSUBS 0.009327f
C239 B.n150 VSUBS 0.009327f
C240 B.n151 VSUBS 0.009327f
C241 B.n152 VSUBS 0.009327f
C242 B.n153 VSUBS 0.009327f
C243 B.n154 VSUBS 0.009327f
C244 B.n155 VSUBS 0.009327f
C245 B.n156 VSUBS 0.009327f
C246 B.n157 VSUBS 0.009327f
C247 B.n158 VSUBS 0.009327f
C248 B.n159 VSUBS 0.009327f
C249 B.n160 VSUBS 0.009327f
C250 B.n161 VSUBS 0.009327f
C251 B.n162 VSUBS 0.009327f
C252 B.n163 VSUBS 0.022059f
C253 B.n164 VSUBS 0.009327f
C254 B.n165 VSUBS 0.009327f
C255 B.n166 VSUBS 0.009327f
C256 B.n167 VSUBS 0.009327f
C257 B.n168 VSUBS 0.009327f
C258 B.n169 VSUBS 0.009327f
C259 B.n170 VSUBS 0.009327f
C260 B.n171 VSUBS 0.009327f
C261 B.n172 VSUBS 0.009327f
C262 B.n173 VSUBS 0.009327f
C263 B.n174 VSUBS 0.009327f
C264 B.n175 VSUBS 0.009327f
C265 B.n176 VSUBS 0.009327f
C266 B.n177 VSUBS 0.009327f
C267 B.n178 VSUBS 0.009327f
C268 B.n179 VSUBS 0.009327f
C269 B.n180 VSUBS 0.009327f
C270 B.n181 VSUBS 0.009327f
C271 B.n182 VSUBS 0.009327f
C272 B.n183 VSUBS 0.009327f
C273 B.n184 VSUBS 0.009327f
C274 B.n185 VSUBS 0.009327f
C275 B.n186 VSUBS 0.009327f
C276 B.n187 VSUBS 0.009327f
C277 B.n188 VSUBS 0.009327f
C278 B.n189 VSUBS 0.009327f
C279 B.n190 VSUBS 0.009327f
C280 B.n191 VSUBS 0.009327f
C281 B.n192 VSUBS 0.009327f
C282 B.n193 VSUBS 0.009327f
C283 B.n194 VSUBS 0.009327f
C284 B.n195 VSUBS 0.009327f
C285 B.n196 VSUBS 0.009327f
C286 B.n197 VSUBS 0.009327f
C287 B.n198 VSUBS 0.009327f
C288 B.n199 VSUBS 0.009327f
C289 B.n200 VSUBS 0.009327f
C290 B.n201 VSUBS 0.009327f
C291 B.n202 VSUBS 0.009327f
C292 B.n203 VSUBS 0.009327f
C293 B.n204 VSUBS 0.009327f
C294 B.n205 VSUBS 0.009327f
C295 B.n206 VSUBS 0.009327f
C296 B.n207 VSUBS 0.009327f
C297 B.n208 VSUBS 0.009327f
C298 B.n209 VSUBS 0.009327f
C299 B.n210 VSUBS 0.009327f
C300 B.n211 VSUBS 0.009327f
C301 B.n212 VSUBS 0.009327f
C302 B.n213 VSUBS 0.009327f
C303 B.n214 VSUBS 0.009327f
C304 B.n215 VSUBS 0.009327f
C305 B.n216 VSUBS 0.009327f
C306 B.n217 VSUBS 0.009327f
C307 B.n218 VSUBS 0.009327f
C308 B.n219 VSUBS 0.009327f
C309 B.n220 VSUBS 0.009327f
C310 B.n221 VSUBS 0.009327f
C311 B.n222 VSUBS 0.009327f
C312 B.n223 VSUBS 0.009327f
C313 B.n224 VSUBS 0.009327f
C314 B.n225 VSUBS 0.009327f
C315 B.n226 VSUBS 0.009327f
C316 B.n227 VSUBS 0.009327f
C317 B.n228 VSUBS 0.009327f
C318 B.n229 VSUBS 0.009327f
C319 B.n230 VSUBS 0.009327f
C320 B.n231 VSUBS 0.009327f
C321 B.n232 VSUBS 0.009327f
C322 B.n233 VSUBS 0.009327f
C323 B.n234 VSUBS 0.009327f
C324 B.n235 VSUBS 0.009327f
C325 B.n236 VSUBS 0.009327f
C326 B.n237 VSUBS 0.009327f
C327 B.n238 VSUBS 0.009327f
C328 B.n239 VSUBS 0.009327f
C329 B.n240 VSUBS 0.009327f
C330 B.n241 VSUBS 0.009327f
C331 B.n242 VSUBS 0.009327f
C332 B.n243 VSUBS 0.009327f
C333 B.n244 VSUBS 0.009327f
C334 B.n245 VSUBS 0.009327f
C335 B.n246 VSUBS 0.009327f
C336 B.n247 VSUBS 0.009327f
C337 B.n248 VSUBS 0.009327f
C338 B.n249 VSUBS 0.009327f
C339 B.n250 VSUBS 0.009327f
C340 B.n251 VSUBS 0.009327f
C341 B.n252 VSUBS 0.009327f
C342 B.n253 VSUBS 0.009327f
C343 B.n254 VSUBS 0.009327f
C344 B.n255 VSUBS 0.009327f
C345 B.n256 VSUBS 0.009327f
C346 B.n257 VSUBS 0.009327f
C347 B.n258 VSUBS 0.022059f
C348 B.n259 VSUBS 0.023205f
C349 B.n260 VSUBS 0.023205f
C350 B.n261 VSUBS 0.009327f
C351 B.n262 VSUBS 0.009327f
C352 B.n263 VSUBS 0.009327f
C353 B.n264 VSUBS 0.009327f
C354 B.n265 VSUBS 0.009327f
C355 B.n266 VSUBS 0.009327f
C356 B.n267 VSUBS 0.009327f
C357 B.n268 VSUBS 0.009327f
C358 B.n269 VSUBS 0.009327f
C359 B.n270 VSUBS 0.009327f
C360 B.n271 VSUBS 0.009327f
C361 B.n272 VSUBS 0.009327f
C362 B.n273 VSUBS 0.009327f
C363 B.n274 VSUBS 0.009327f
C364 B.n275 VSUBS 0.009327f
C365 B.n276 VSUBS 0.009327f
C366 B.n277 VSUBS 0.009327f
C367 B.n278 VSUBS 0.009327f
C368 B.n279 VSUBS 0.009327f
C369 B.n280 VSUBS 0.009327f
C370 B.n281 VSUBS 0.009327f
C371 B.n282 VSUBS 0.009327f
C372 B.n283 VSUBS 0.009327f
C373 B.n284 VSUBS 0.009327f
C374 B.n285 VSUBS 0.009327f
C375 B.n286 VSUBS 0.009327f
C376 B.n287 VSUBS 0.009327f
C377 B.n288 VSUBS 0.009327f
C378 B.n289 VSUBS 0.009327f
C379 B.n290 VSUBS 0.009327f
C380 B.n291 VSUBS 0.009327f
C381 B.n292 VSUBS 0.009327f
C382 B.n293 VSUBS 0.009327f
C383 B.n294 VSUBS 0.009327f
C384 B.n295 VSUBS 0.009327f
C385 B.n296 VSUBS 0.009327f
C386 B.n297 VSUBS 0.009327f
C387 B.n298 VSUBS 0.009327f
C388 B.n299 VSUBS 0.009327f
C389 B.n300 VSUBS 0.009327f
C390 B.n301 VSUBS 0.009327f
C391 B.n302 VSUBS 0.009327f
C392 B.n303 VSUBS 0.009327f
C393 B.n304 VSUBS 0.009327f
C394 B.n305 VSUBS 0.009327f
C395 B.n306 VSUBS 0.009327f
C396 B.n307 VSUBS 0.009327f
C397 B.n308 VSUBS 0.009327f
C398 B.n309 VSUBS 0.009327f
C399 B.n310 VSUBS 0.009327f
C400 B.n311 VSUBS 0.008778f
C401 B.n312 VSUBS 0.02161f
C402 B.n313 VSUBS 0.005212f
C403 B.n314 VSUBS 0.009327f
C404 B.n315 VSUBS 0.009327f
C405 B.n316 VSUBS 0.009327f
C406 B.n317 VSUBS 0.009327f
C407 B.n318 VSUBS 0.009327f
C408 B.n319 VSUBS 0.009327f
C409 B.n320 VSUBS 0.009327f
C410 B.n321 VSUBS 0.009327f
C411 B.n322 VSUBS 0.009327f
C412 B.n323 VSUBS 0.009327f
C413 B.n324 VSUBS 0.009327f
C414 B.n325 VSUBS 0.009327f
C415 B.t8 VSUBS 0.417203f
C416 B.t7 VSUBS 0.449286f
C417 B.t6 VSUBS 1.958f
C418 B.n326 VSUBS 0.248493f
C419 B.n327 VSUBS 0.098787f
C420 B.n328 VSUBS 0.02161f
C421 B.n329 VSUBS 0.005212f
C422 B.n330 VSUBS 0.009327f
C423 B.n331 VSUBS 0.009327f
C424 B.n332 VSUBS 0.009327f
C425 B.n333 VSUBS 0.009327f
C426 B.n334 VSUBS 0.009327f
C427 B.n335 VSUBS 0.009327f
C428 B.n336 VSUBS 0.009327f
C429 B.n337 VSUBS 0.009327f
C430 B.n338 VSUBS 0.009327f
C431 B.n339 VSUBS 0.009327f
C432 B.n340 VSUBS 0.009327f
C433 B.n341 VSUBS 0.009327f
C434 B.n342 VSUBS 0.009327f
C435 B.n343 VSUBS 0.009327f
C436 B.n344 VSUBS 0.009327f
C437 B.n345 VSUBS 0.009327f
C438 B.n346 VSUBS 0.009327f
C439 B.n347 VSUBS 0.009327f
C440 B.n348 VSUBS 0.009327f
C441 B.n349 VSUBS 0.009327f
C442 B.n350 VSUBS 0.009327f
C443 B.n351 VSUBS 0.009327f
C444 B.n352 VSUBS 0.009327f
C445 B.n353 VSUBS 0.009327f
C446 B.n354 VSUBS 0.009327f
C447 B.n355 VSUBS 0.009327f
C448 B.n356 VSUBS 0.009327f
C449 B.n357 VSUBS 0.009327f
C450 B.n358 VSUBS 0.009327f
C451 B.n359 VSUBS 0.009327f
C452 B.n360 VSUBS 0.009327f
C453 B.n361 VSUBS 0.009327f
C454 B.n362 VSUBS 0.009327f
C455 B.n363 VSUBS 0.009327f
C456 B.n364 VSUBS 0.009327f
C457 B.n365 VSUBS 0.009327f
C458 B.n366 VSUBS 0.009327f
C459 B.n367 VSUBS 0.009327f
C460 B.n368 VSUBS 0.009327f
C461 B.n369 VSUBS 0.009327f
C462 B.n370 VSUBS 0.009327f
C463 B.n371 VSUBS 0.009327f
C464 B.n372 VSUBS 0.009327f
C465 B.n373 VSUBS 0.009327f
C466 B.n374 VSUBS 0.009327f
C467 B.n375 VSUBS 0.009327f
C468 B.n376 VSUBS 0.009327f
C469 B.n377 VSUBS 0.009327f
C470 B.n378 VSUBS 0.009327f
C471 B.n379 VSUBS 0.009327f
C472 B.n380 VSUBS 0.009327f
C473 B.n381 VSUBS 0.009327f
C474 B.n382 VSUBS 0.022161f
C475 B.n383 VSUBS 0.023103f
C476 B.n384 VSUBS 0.022059f
C477 B.n385 VSUBS 0.009327f
C478 B.n386 VSUBS 0.009327f
C479 B.n387 VSUBS 0.009327f
C480 B.n388 VSUBS 0.009327f
C481 B.n389 VSUBS 0.009327f
C482 B.n390 VSUBS 0.009327f
C483 B.n391 VSUBS 0.009327f
C484 B.n392 VSUBS 0.009327f
C485 B.n393 VSUBS 0.009327f
C486 B.n394 VSUBS 0.009327f
C487 B.n395 VSUBS 0.009327f
C488 B.n396 VSUBS 0.009327f
C489 B.n397 VSUBS 0.009327f
C490 B.n398 VSUBS 0.009327f
C491 B.n399 VSUBS 0.009327f
C492 B.n400 VSUBS 0.009327f
C493 B.n401 VSUBS 0.009327f
C494 B.n402 VSUBS 0.009327f
C495 B.n403 VSUBS 0.009327f
C496 B.n404 VSUBS 0.009327f
C497 B.n405 VSUBS 0.009327f
C498 B.n406 VSUBS 0.009327f
C499 B.n407 VSUBS 0.009327f
C500 B.n408 VSUBS 0.009327f
C501 B.n409 VSUBS 0.009327f
C502 B.n410 VSUBS 0.009327f
C503 B.n411 VSUBS 0.009327f
C504 B.n412 VSUBS 0.009327f
C505 B.n413 VSUBS 0.009327f
C506 B.n414 VSUBS 0.009327f
C507 B.n415 VSUBS 0.009327f
C508 B.n416 VSUBS 0.009327f
C509 B.n417 VSUBS 0.009327f
C510 B.n418 VSUBS 0.009327f
C511 B.n419 VSUBS 0.009327f
C512 B.n420 VSUBS 0.009327f
C513 B.n421 VSUBS 0.009327f
C514 B.n422 VSUBS 0.009327f
C515 B.n423 VSUBS 0.009327f
C516 B.n424 VSUBS 0.009327f
C517 B.n425 VSUBS 0.009327f
C518 B.n426 VSUBS 0.009327f
C519 B.n427 VSUBS 0.009327f
C520 B.n428 VSUBS 0.009327f
C521 B.n429 VSUBS 0.009327f
C522 B.n430 VSUBS 0.009327f
C523 B.n431 VSUBS 0.009327f
C524 B.n432 VSUBS 0.009327f
C525 B.n433 VSUBS 0.009327f
C526 B.n434 VSUBS 0.009327f
C527 B.n435 VSUBS 0.009327f
C528 B.n436 VSUBS 0.009327f
C529 B.n437 VSUBS 0.009327f
C530 B.n438 VSUBS 0.009327f
C531 B.n439 VSUBS 0.009327f
C532 B.n440 VSUBS 0.009327f
C533 B.n441 VSUBS 0.009327f
C534 B.n442 VSUBS 0.009327f
C535 B.n443 VSUBS 0.009327f
C536 B.n444 VSUBS 0.009327f
C537 B.n445 VSUBS 0.009327f
C538 B.n446 VSUBS 0.009327f
C539 B.n447 VSUBS 0.009327f
C540 B.n448 VSUBS 0.009327f
C541 B.n449 VSUBS 0.009327f
C542 B.n450 VSUBS 0.009327f
C543 B.n451 VSUBS 0.009327f
C544 B.n452 VSUBS 0.009327f
C545 B.n453 VSUBS 0.009327f
C546 B.n454 VSUBS 0.009327f
C547 B.n455 VSUBS 0.009327f
C548 B.n456 VSUBS 0.009327f
C549 B.n457 VSUBS 0.009327f
C550 B.n458 VSUBS 0.009327f
C551 B.n459 VSUBS 0.009327f
C552 B.n460 VSUBS 0.009327f
C553 B.n461 VSUBS 0.009327f
C554 B.n462 VSUBS 0.009327f
C555 B.n463 VSUBS 0.009327f
C556 B.n464 VSUBS 0.009327f
C557 B.n465 VSUBS 0.009327f
C558 B.n466 VSUBS 0.009327f
C559 B.n467 VSUBS 0.009327f
C560 B.n468 VSUBS 0.009327f
C561 B.n469 VSUBS 0.009327f
C562 B.n470 VSUBS 0.009327f
C563 B.n471 VSUBS 0.009327f
C564 B.n472 VSUBS 0.009327f
C565 B.n473 VSUBS 0.009327f
C566 B.n474 VSUBS 0.009327f
C567 B.n475 VSUBS 0.009327f
C568 B.n476 VSUBS 0.009327f
C569 B.n477 VSUBS 0.009327f
C570 B.n478 VSUBS 0.009327f
C571 B.n479 VSUBS 0.009327f
C572 B.n480 VSUBS 0.009327f
C573 B.n481 VSUBS 0.009327f
C574 B.n482 VSUBS 0.009327f
C575 B.n483 VSUBS 0.009327f
C576 B.n484 VSUBS 0.009327f
C577 B.n485 VSUBS 0.009327f
C578 B.n486 VSUBS 0.009327f
C579 B.n487 VSUBS 0.009327f
C580 B.n488 VSUBS 0.009327f
C581 B.n489 VSUBS 0.009327f
C582 B.n490 VSUBS 0.009327f
C583 B.n491 VSUBS 0.009327f
C584 B.n492 VSUBS 0.009327f
C585 B.n493 VSUBS 0.009327f
C586 B.n494 VSUBS 0.009327f
C587 B.n495 VSUBS 0.009327f
C588 B.n496 VSUBS 0.009327f
C589 B.n497 VSUBS 0.009327f
C590 B.n498 VSUBS 0.009327f
C591 B.n499 VSUBS 0.009327f
C592 B.n500 VSUBS 0.009327f
C593 B.n501 VSUBS 0.009327f
C594 B.n502 VSUBS 0.009327f
C595 B.n503 VSUBS 0.009327f
C596 B.n504 VSUBS 0.009327f
C597 B.n505 VSUBS 0.009327f
C598 B.n506 VSUBS 0.009327f
C599 B.n507 VSUBS 0.009327f
C600 B.n508 VSUBS 0.009327f
C601 B.n509 VSUBS 0.009327f
C602 B.n510 VSUBS 0.009327f
C603 B.n511 VSUBS 0.009327f
C604 B.n512 VSUBS 0.009327f
C605 B.n513 VSUBS 0.009327f
C606 B.n514 VSUBS 0.009327f
C607 B.n515 VSUBS 0.009327f
C608 B.n516 VSUBS 0.009327f
C609 B.n517 VSUBS 0.009327f
C610 B.n518 VSUBS 0.009327f
C611 B.n519 VSUBS 0.009327f
C612 B.n520 VSUBS 0.009327f
C613 B.n521 VSUBS 0.009327f
C614 B.n522 VSUBS 0.009327f
C615 B.n523 VSUBS 0.009327f
C616 B.n524 VSUBS 0.009327f
C617 B.n525 VSUBS 0.009327f
C618 B.n526 VSUBS 0.009327f
C619 B.n527 VSUBS 0.009327f
C620 B.n528 VSUBS 0.009327f
C621 B.n529 VSUBS 0.009327f
C622 B.n530 VSUBS 0.009327f
C623 B.n531 VSUBS 0.009327f
C624 B.n532 VSUBS 0.022059f
C625 B.n533 VSUBS 0.023205f
C626 B.n534 VSUBS 0.023205f
C627 B.n535 VSUBS 0.009327f
C628 B.n536 VSUBS 0.009327f
C629 B.n537 VSUBS 0.009327f
C630 B.n538 VSUBS 0.009327f
C631 B.n539 VSUBS 0.009327f
C632 B.n540 VSUBS 0.009327f
C633 B.n541 VSUBS 0.009327f
C634 B.n542 VSUBS 0.009327f
C635 B.n543 VSUBS 0.009327f
C636 B.n544 VSUBS 0.009327f
C637 B.n545 VSUBS 0.009327f
C638 B.n546 VSUBS 0.009327f
C639 B.n547 VSUBS 0.009327f
C640 B.n548 VSUBS 0.009327f
C641 B.n549 VSUBS 0.009327f
C642 B.n550 VSUBS 0.009327f
C643 B.n551 VSUBS 0.009327f
C644 B.n552 VSUBS 0.009327f
C645 B.n553 VSUBS 0.009327f
C646 B.n554 VSUBS 0.009327f
C647 B.n555 VSUBS 0.009327f
C648 B.n556 VSUBS 0.009327f
C649 B.n557 VSUBS 0.009327f
C650 B.n558 VSUBS 0.009327f
C651 B.n559 VSUBS 0.009327f
C652 B.n560 VSUBS 0.009327f
C653 B.n561 VSUBS 0.009327f
C654 B.n562 VSUBS 0.009327f
C655 B.n563 VSUBS 0.009327f
C656 B.n564 VSUBS 0.009327f
C657 B.n565 VSUBS 0.009327f
C658 B.n566 VSUBS 0.009327f
C659 B.n567 VSUBS 0.009327f
C660 B.n568 VSUBS 0.009327f
C661 B.n569 VSUBS 0.009327f
C662 B.n570 VSUBS 0.009327f
C663 B.n571 VSUBS 0.009327f
C664 B.n572 VSUBS 0.009327f
C665 B.n573 VSUBS 0.009327f
C666 B.n574 VSUBS 0.009327f
C667 B.n575 VSUBS 0.009327f
C668 B.n576 VSUBS 0.009327f
C669 B.n577 VSUBS 0.009327f
C670 B.n578 VSUBS 0.009327f
C671 B.n579 VSUBS 0.009327f
C672 B.n580 VSUBS 0.009327f
C673 B.n581 VSUBS 0.009327f
C674 B.n582 VSUBS 0.009327f
C675 B.n583 VSUBS 0.009327f
C676 B.n584 VSUBS 0.009327f
C677 B.n585 VSUBS 0.008778f
C678 B.n586 VSUBS 0.02161f
C679 B.n587 VSUBS 0.005212f
C680 B.n588 VSUBS 0.009327f
C681 B.n589 VSUBS 0.009327f
C682 B.n590 VSUBS 0.009327f
C683 B.n591 VSUBS 0.009327f
C684 B.n592 VSUBS 0.009327f
C685 B.n593 VSUBS 0.009327f
C686 B.n594 VSUBS 0.009327f
C687 B.n595 VSUBS 0.009327f
C688 B.n596 VSUBS 0.009327f
C689 B.n597 VSUBS 0.009327f
C690 B.n598 VSUBS 0.009327f
C691 B.n599 VSUBS 0.009327f
C692 B.n600 VSUBS 0.005212f
C693 B.n601 VSUBS 0.009327f
C694 B.n602 VSUBS 0.009327f
C695 B.n603 VSUBS 0.008778f
C696 B.n604 VSUBS 0.009327f
C697 B.n605 VSUBS 0.009327f
C698 B.n606 VSUBS 0.009327f
C699 B.n607 VSUBS 0.009327f
C700 B.n608 VSUBS 0.009327f
C701 B.n609 VSUBS 0.009327f
C702 B.n610 VSUBS 0.009327f
C703 B.n611 VSUBS 0.009327f
C704 B.n612 VSUBS 0.009327f
C705 B.n613 VSUBS 0.009327f
C706 B.n614 VSUBS 0.009327f
C707 B.n615 VSUBS 0.009327f
C708 B.n616 VSUBS 0.009327f
C709 B.n617 VSUBS 0.009327f
C710 B.n618 VSUBS 0.009327f
C711 B.n619 VSUBS 0.009327f
C712 B.n620 VSUBS 0.009327f
C713 B.n621 VSUBS 0.009327f
C714 B.n622 VSUBS 0.009327f
C715 B.n623 VSUBS 0.009327f
C716 B.n624 VSUBS 0.009327f
C717 B.n625 VSUBS 0.009327f
C718 B.n626 VSUBS 0.009327f
C719 B.n627 VSUBS 0.009327f
C720 B.n628 VSUBS 0.009327f
C721 B.n629 VSUBS 0.009327f
C722 B.n630 VSUBS 0.009327f
C723 B.n631 VSUBS 0.009327f
C724 B.n632 VSUBS 0.009327f
C725 B.n633 VSUBS 0.009327f
C726 B.n634 VSUBS 0.009327f
C727 B.n635 VSUBS 0.009327f
C728 B.n636 VSUBS 0.009327f
C729 B.n637 VSUBS 0.009327f
C730 B.n638 VSUBS 0.009327f
C731 B.n639 VSUBS 0.009327f
C732 B.n640 VSUBS 0.009327f
C733 B.n641 VSUBS 0.009327f
C734 B.n642 VSUBS 0.009327f
C735 B.n643 VSUBS 0.009327f
C736 B.n644 VSUBS 0.009327f
C737 B.n645 VSUBS 0.009327f
C738 B.n646 VSUBS 0.009327f
C739 B.n647 VSUBS 0.009327f
C740 B.n648 VSUBS 0.009327f
C741 B.n649 VSUBS 0.009327f
C742 B.n650 VSUBS 0.009327f
C743 B.n651 VSUBS 0.009327f
C744 B.n652 VSUBS 0.009327f
C745 B.n653 VSUBS 0.023205f
C746 B.n654 VSUBS 0.023205f
C747 B.n655 VSUBS 0.022059f
C748 B.n656 VSUBS 0.009327f
C749 B.n657 VSUBS 0.009327f
C750 B.n658 VSUBS 0.009327f
C751 B.n659 VSUBS 0.009327f
C752 B.n660 VSUBS 0.009327f
C753 B.n661 VSUBS 0.009327f
C754 B.n662 VSUBS 0.009327f
C755 B.n663 VSUBS 0.009327f
C756 B.n664 VSUBS 0.009327f
C757 B.n665 VSUBS 0.009327f
C758 B.n666 VSUBS 0.009327f
C759 B.n667 VSUBS 0.009327f
C760 B.n668 VSUBS 0.009327f
C761 B.n669 VSUBS 0.009327f
C762 B.n670 VSUBS 0.009327f
C763 B.n671 VSUBS 0.009327f
C764 B.n672 VSUBS 0.009327f
C765 B.n673 VSUBS 0.009327f
C766 B.n674 VSUBS 0.009327f
C767 B.n675 VSUBS 0.009327f
C768 B.n676 VSUBS 0.009327f
C769 B.n677 VSUBS 0.009327f
C770 B.n678 VSUBS 0.009327f
C771 B.n679 VSUBS 0.009327f
C772 B.n680 VSUBS 0.009327f
C773 B.n681 VSUBS 0.009327f
C774 B.n682 VSUBS 0.009327f
C775 B.n683 VSUBS 0.009327f
C776 B.n684 VSUBS 0.009327f
C777 B.n685 VSUBS 0.009327f
C778 B.n686 VSUBS 0.009327f
C779 B.n687 VSUBS 0.009327f
C780 B.n688 VSUBS 0.009327f
C781 B.n689 VSUBS 0.009327f
C782 B.n690 VSUBS 0.009327f
C783 B.n691 VSUBS 0.009327f
C784 B.n692 VSUBS 0.009327f
C785 B.n693 VSUBS 0.009327f
C786 B.n694 VSUBS 0.009327f
C787 B.n695 VSUBS 0.009327f
C788 B.n696 VSUBS 0.009327f
C789 B.n697 VSUBS 0.009327f
C790 B.n698 VSUBS 0.009327f
C791 B.n699 VSUBS 0.009327f
C792 B.n700 VSUBS 0.009327f
C793 B.n701 VSUBS 0.009327f
C794 B.n702 VSUBS 0.009327f
C795 B.n703 VSUBS 0.009327f
C796 B.n704 VSUBS 0.009327f
C797 B.n705 VSUBS 0.009327f
C798 B.n706 VSUBS 0.009327f
C799 B.n707 VSUBS 0.009327f
C800 B.n708 VSUBS 0.009327f
C801 B.n709 VSUBS 0.009327f
C802 B.n710 VSUBS 0.009327f
C803 B.n711 VSUBS 0.009327f
C804 B.n712 VSUBS 0.009327f
C805 B.n713 VSUBS 0.009327f
C806 B.n714 VSUBS 0.009327f
C807 B.n715 VSUBS 0.009327f
C808 B.n716 VSUBS 0.009327f
C809 B.n717 VSUBS 0.009327f
C810 B.n718 VSUBS 0.009327f
C811 B.n719 VSUBS 0.009327f
C812 B.n720 VSUBS 0.009327f
C813 B.n721 VSUBS 0.009327f
C814 B.n722 VSUBS 0.009327f
C815 B.n723 VSUBS 0.009327f
C816 B.n724 VSUBS 0.009327f
C817 B.n725 VSUBS 0.009327f
C818 B.n726 VSUBS 0.009327f
C819 B.n727 VSUBS 0.012171f
C820 B.n728 VSUBS 0.012966f
C821 B.n729 VSUBS 0.025783f
C822 VDD1.t2 VSUBS 2.23169f
C823 VDD1.t0 VSUBS 2.23023f
C824 VDD1.t1 VSUBS 0.225828f
C825 VDD1.t4 VSUBS 0.225828f
C826 VDD1.n0 VSUBS 1.68566f
C827 VDD1.n1 VSUBS 4.29787f
C828 VDD1.t3 VSUBS 0.225828f
C829 VDD1.t5 VSUBS 0.225828f
C830 VDD1.n2 VSUBS 1.67729f
C831 VDD1.n3 VSUBS 3.55155f
C832 VTAIL.t3 VSUBS 0.237969f
C833 VTAIL.t0 VSUBS 0.237969f
C834 VTAIL.n0 VSUBS 1.60714f
C835 VTAIL.n1 VSUBS 0.970578f
C836 VTAIL.t11 VSUBS 2.14946f
C837 VTAIL.n2 VSUBS 1.29659f
C838 VTAIL.t10 VSUBS 0.237969f
C839 VTAIL.t6 VSUBS 0.237969f
C840 VTAIL.n3 VSUBS 1.60714f
C841 VTAIL.n4 VSUBS 2.84591f
C842 VTAIL.t2 VSUBS 0.237969f
C843 VTAIL.t4 VSUBS 0.237969f
C844 VTAIL.n5 VSUBS 1.60715f
C845 VTAIL.n6 VSUBS 2.8459f
C846 VTAIL.t5 VSUBS 2.14947f
C847 VTAIL.n7 VSUBS 1.29658f
C848 VTAIL.t8 VSUBS 0.237969f
C849 VTAIL.t7 VSUBS 0.237969f
C850 VTAIL.n8 VSUBS 1.60715f
C851 VTAIL.n9 VSUBS 1.18989f
C852 VTAIL.t9 VSUBS 2.14947f
C853 VTAIL.n10 VSUBS 2.6525f
C854 VTAIL.t1 VSUBS 2.14946f
C855 VTAIL.n11 VSUBS 2.57176f
C856 VP.t1 VSUBS 2.75859f
C857 VP.n0 VSUBS 1.10248f
C858 VP.n1 VSUBS 0.032357f
C859 VP.n2 VSUBS 0.026227f
C860 VP.n3 VSUBS 0.032357f
C861 VP.t4 VSUBS 2.75859f
C862 VP.n4 VSUBS 0.981394f
C863 VP.n5 VSUBS 0.032357f
C864 VP.n6 VSUBS 0.026227f
C865 VP.n7 VSUBS 0.032357f
C866 VP.t5 VSUBS 2.75859f
C867 VP.n8 VSUBS 1.10248f
C868 VP.t0 VSUBS 2.75859f
C869 VP.n9 VSUBS 1.10248f
C870 VP.n10 VSUBS 0.032357f
C871 VP.n11 VSUBS 0.026227f
C872 VP.n12 VSUBS 0.032357f
C873 VP.t2 VSUBS 2.75859f
C874 VP.n13 VSUBS 1.08718f
C875 VP.t3 VSUBS 3.12957f
C876 VP.n14 VSUBS 1.03422f
C877 VP.n15 VSUBS 0.376587f
C878 VP.n16 VSUBS 0.045192f
C879 VP.n17 VSUBS 0.060003f
C880 VP.n18 VSUBS 0.064404f
C881 VP.n19 VSUBS 0.032357f
C882 VP.n20 VSUBS 0.032357f
C883 VP.n21 VSUBS 0.032357f
C884 VP.n22 VSUBS 0.063444f
C885 VP.n23 VSUBS 0.060003f
C886 VP.n24 VSUBS 0.046969f
C887 VP.n25 VSUBS 0.052215f
C888 VP.n26 VSUBS 1.81074f
C889 VP.n27 VSUBS 1.83432f
C890 VP.n28 VSUBS 0.052215f
C891 VP.n29 VSUBS 0.046969f
C892 VP.n30 VSUBS 0.060003f
C893 VP.n31 VSUBS 0.063444f
C894 VP.n32 VSUBS 0.032357f
C895 VP.n33 VSUBS 0.032357f
C896 VP.n34 VSUBS 0.032357f
C897 VP.n35 VSUBS 0.064404f
C898 VP.n36 VSUBS 0.060003f
C899 VP.n37 VSUBS 0.045192f
C900 VP.n38 VSUBS 0.032357f
C901 VP.n39 VSUBS 0.032357f
C902 VP.n40 VSUBS 0.045192f
C903 VP.n41 VSUBS 0.060003f
C904 VP.n42 VSUBS 0.064404f
C905 VP.n43 VSUBS 0.032357f
C906 VP.n44 VSUBS 0.032357f
C907 VP.n45 VSUBS 0.032357f
C908 VP.n46 VSUBS 0.063444f
C909 VP.n47 VSUBS 0.060003f
C910 VP.n48 VSUBS 0.046969f
C911 VP.n49 VSUBS 0.052215f
C912 VP.n50 VSUBS 0.078099f
.ends

