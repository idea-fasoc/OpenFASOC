* NGSPICE file created from diff_pair_sample_0967.ext - technology: sky130A

.subckt diff_pair_sample_0967 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t3 w_n2662_n1372# sky130_fd_pr__pfet_01v8 ad=0.7878 pd=4.82 as=0.7878 ps=4.82 w=2.02 l=3.9
X1 VDD2.t1 VN.t0 VTAIL.t1 w_n2662_n1372# sky130_fd_pr__pfet_01v8 ad=0.7878 pd=4.82 as=0.7878 ps=4.82 w=2.02 l=3.9
X2 VDD1.t0 VP.t1 VTAIL.t2 w_n2662_n1372# sky130_fd_pr__pfet_01v8 ad=0.7878 pd=4.82 as=0.7878 ps=4.82 w=2.02 l=3.9
X3 B.t11 B.t9 B.t10 w_n2662_n1372# sky130_fd_pr__pfet_01v8 ad=0.7878 pd=4.82 as=0 ps=0 w=2.02 l=3.9
X4 B.t8 B.t6 B.t7 w_n2662_n1372# sky130_fd_pr__pfet_01v8 ad=0.7878 pd=4.82 as=0 ps=0 w=2.02 l=3.9
X5 B.t5 B.t3 B.t4 w_n2662_n1372# sky130_fd_pr__pfet_01v8 ad=0.7878 pd=4.82 as=0 ps=0 w=2.02 l=3.9
X6 B.t2 B.t0 B.t1 w_n2662_n1372# sky130_fd_pr__pfet_01v8 ad=0.7878 pd=4.82 as=0 ps=0 w=2.02 l=3.9
X7 VDD2.t0 VN.t1 VTAIL.t0 w_n2662_n1372# sky130_fd_pr__pfet_01v8 ad=0.7878 pd=4.82 as=0.7878 ps=4.82 w=2.02 l=3.9
R0 VP.n0 VP.t1 88.0094
R1 VP.n0 VP.t0 47.4662
R2 VP VP.n0 0.621233
R3 VTAIL.n26 VTAIL.n24 756.745
R4 VTAIL.n2 VTAIL.n0 756.745
R5 VTAIL.n18 VTAIL.n16 756.745
R6 VTAIL.n10 VTAIL.n8 756.745
R7 VTAIL.n27 VTAIL.n26 585
R8 VTAIL.n3 VTAIL.n2 585
R9 VTAIL.n19 VTAIL.n18 585
R10 VTAIL.n11 VTAIL.n10 585
R11 VTAIL.t0 VTAIL.n25 417.779
R12 VTAIL.t3 VTAIL.n1 417.779
R13 VTAIL.t2 VTAIL.n17 417.779
R14 VTAIL.t1 VTAIL.n9 417.779
R15 VTAIL.n26 VTAIL.t0 85.8723
R16 VTAIL.n2 VTAIL.t3 85.8723
R17 VTAIL.n18 VTAIL.t2 85.8723
R18 VTAIL.n10 VTAIL.t1 85.8723
R19 VTAIL.n31 VTAIL.n30 31.7975
R20 VTAIL.n7 VTAIL.n6 31.7975
R21 VTAIL.n23 VTAIL.n22 31.7975
R22 VTAIL.n15 VTAIL.n14 31.7975
R23 VTAIL.n15 VTAIL.n7 21.4014
R24 VTAIL.n31 VTAIL.n23 17.7548
R25 VTAIL.n27 VTAIL.n25 9.84608
R26 VTAIL.n3 VTAIL.n1 9.84608
R27 VTAIL.n19 VTAIL.n17 9.84608
R28 VTAIL.n11 VTAIL.n9 9.84608
R29 VTAIL.n30 VTAIL.n29 9.45567
R30 VTAIL.n6 VTAIL.n5 9.45567
R31 VTAIL.n22 VTAIL.n21 9.45567
R32 VTAIL.n14 VTAIL.n13 9.45567
R33 VTAIL.n29 VTAIL.n28 9.3005
R34 VTAIL.n5 VTAIL.n4 9.3005
R35 VTAIL.n21 VTAIL.n20 9.3005
R36 VTAIL.n13 VTAIL.n12 9.3005
R37 VTAIL.n30 VTAIL.n24 8.14595
R38 VTAIL.n6 VTAIL.n0 8.14595
R39 VTAIL.n22 VTAIL.n16 8.14595
R40 VTAIL.n14 VTAIL.n8 8.14595
R41 VTAIL.n28 VTAIL.n27 7.3702
R42 VTAIL.n4 VTAIL.n3 7.3702
R43 VTAIL.n20 VTAIL.n19 7.3702
R44 VTAIL.n12 VTAIL.n11 7.3702
R45 VTAIL.n28 VTAIL.n24 5.81868
R46 VTAIL.n4 VTAIL.n0 5.81868
R47 VTAIL.n20 VTAIL.n16 5.81868
R48 VTAIL.n12 VTAIL.n8 5.81868
R49 VTAIL.n13 VTAIL.n9 3.32369
R50 VTAIL.n29 VTAIL.n25 3.32369
R51 VTAIL.n5 VTAIL.n1 3.32369
R52 VTAIL.n21 VTAIL.n17 3.32369
R53 VTAIL.n23 VTAIL.n15 2.2936
R54 VTAIL VTAIL.n7 1.44016
R55 VTAIL VTAIL.n31 0.853948
R56 VDD1.n2 VDD1.n0 756.745
R57 VDD1.n9 VDD1.n7 756.745
R58 VDD1.n3 VDD1.n2 585
R59 VDD1.n10 VDD1.n9 585
R60 VDD1.t1 VDD1.n8 417.779
R61 VDD1.t0 VDD1.n1 417.779
R62 VDD1.n2 VDD1.t0 85.8723
R63 VDD1.n9 VDD1.t1 85.8723
R64 VDD1 VDD1.n13 82.6066
R65 VDD1 VDD1.n6 49.4461
R66 VDD1.n3 VDD1.n1 9.84608
R67 VDD1.n10 VDD1.n8 9.84608
R68 VDD1.n6 VDD1.n5 9.45567
R69 VDD1.n13 VDD1.n12 9.45567
R70 VDD1.n5 VDD1.n4 9.3005
R71 VDD1.n12 VDD1.n11 9.3005
R72 VDD1.n6 VDD1.n0 8.14595
R73 VDD1.n13 VDD1.n7 8.14595
R74 VDD1.n4 VDD1.n3 7.3702
R75 VDD1.n11 VDD1.n10 7.3702
R76 VDD1.n4 VDD1.n0 5.81868
R77 VDD1.n11 VDD1.n7 5.81868
R78 VDD1.n5 VDD1.n1 3.32369
R79 VDD1.n12 VDD1.n8 3.32369
R80 VN VN.t0 87.8217
R81 VN VN.t1 48.0869
R82 VDD2.n9 VDD2.n7 756.745
R83 VDD2.n2 VDD2.n0 756.745
R84 VDD2.n10 VDD2.n9 585
R85 VDD2.n3 VDD2.n2 585
R86 VDD2.t0 VDD2.n1 417.779
R87 VDD2.t1 VDD2.n8 417.779
R88 VDD2.n9 VDD2.t1 85.8723
R89 VDD2.n2 VDD2.t0 85.8723
R90 VDD2.n14 VDD2.n6 81.1702
R91 VDD2.n14 VDD2.n13 48.4763
R92 VDD2.n10 VDD2.n8 9.84608
R93 VDD2.n3 VDD2.n1 9.84608
R94 VDD2.n13 VDD2.n12 9.45567
R95 VDD2.n6 VDD2.n5 9.45567
R96 VDD2.n12 VDD2.n11 9.3005
R97 VDD2.n5 VDD2.n4 9.3005
R98 VDD2.n13 VDD2.n7 8.14595
R99 VDD2.n6 VDD2.n0 8.14595
R100 VDD2.n11 VDD2.n10 7.3702
R101 VDD2.n4 VDD2.n3 7.3702
R102 VDD2.n11 VDD2.n7 5.81868
R103 VDD2.n4 VDD2.n0 5.81868
R104 VDD2.n12 VDD2.n8 3.32369
R105 VDD2.n5 VDD2.n1 3.32369
R106 VDD2 VDD2.n14 0.970328
R107 B.n313 B.n40 585
R108 B.n315 B.n314 585
R109 B.n316 B.n39 585
R110 B.n318 B.n317 585
R111 B.n319 B.n38 585
R112 B.n321 B.n320 585
R113 B.n322 B.n37 585
R114 B.n324 B.n323 585
R115 B.n325 B.n36 585
R116 B.n327 B.n326 585
R117 B.n328 B.n35 585
R118 B.n330 B.n329 585
R119 B.n332 B.n32 585
R120 B.n334 B.n333 585
R121 B.n335 B.n31 585
R122 B.n337 B.n336 585
R123 B.n338 B.n30 585
R124 B.n340 B.n339 585
R125 B.n341 B.n29 585
R126 B.n343 B.n342 585
R127 B.n344 B.n25 585
R128 B.n346 B.n345 585
R129 B.n347 B.n24 585
R130 B.n349 B.n348 585
R131 B.n350 B.n23 585
R132 B.n352 B.n351 585
R133 B.n353 B.n22 585
R134 B.n355 B.n354 585
R135 B.n356 B.n21 585
R136 B.n358 B.n357 585
R137 B.n359 B.n20 585
R138 B.n361 B.n360 585
R139 B.n362 B.n19 585
R140 B.n364 B.n363 585
R141 B.n312 B.n311 585
R142 B.n310 B.n41 585
R143 B.n309 B.n308 585
R144 B.n307 B.n42 585
R145 B.n306 B.n305 585
R146 B.n304 B.n43 585
R147 B.n303 B.n302 585
R148 B.n301 B.n44 585
R149 B.n300 B.n299 585
R150 B.n298 B.n45 585
R151 B.n297 B.n296 585
R152 B.n295 B.n46 585
R153 B.n294 B.n293 585
R154 B.n292 B.n47 585
R155 B.n291 B.n290 585
R156 B.n289 B.n48 585
R157 B.n288 B.n287 585
R158 B.n286 B.n49 585
R159 B.n285 B.n284 585
R160 B.n283 B.n50 585
R161 B.n282 B.n281 585
R162 B.n280 B.n51 585
R163 B.n279 B.n278 585
R164 B.n277 B.n52 585
R165 B.n276 B.n275 585
R166 B.n274 B.n53 585
R167 B.n273 B.n272 585
R168 B.n271 B.n54 585
R169 B.n270 B.n269 585
R170 B.n268 B.n55 585
R171 B.n267 B.n266 585
R172 B.n265 B.n56 585
R173 B.n264 B.n263 585
R174 B.n262 B.n57 585
R175 B.n261 B.n260 585
R176 B.n259 B.n58 585
R177 B.n258 B.n257 585
R178 B.n256 B.n59 585
R179 B.n255 B.n254 585
R180 B.n253 B.n60 585
R181 B.n252 B.n251 585
R182 B.n250 B.n61 585
R183 B.n249 B.n248 585
R184 B.n247 B.n62 585
R185 B.n246 B.n245 585
R186 B.n244 B.n63 585
R187 B.n243 B.n242 585
R188 B.n241 B.n64 585
R189 B.n240 B.n239 585
R190 B.n238 B.n65 585
R191 B.n237 B.n236 585
R192 B.n235 B.n66 585
R193 B.n234 B.n233 585
R194 B.n232 B.n67 585
R195 B.n231 B.n230 585
R196 B.n229 B.n68 585
R197 B.n228 B.n227 585
R198 B.n226 B.n69 585
R199 B.n225 B.n224 585
R200 B.n223 B.n70 585
R201 B.n222 B.n221 585
R202 B.n220 B.n71 585
R203 B.n219 B.n218 585
R204 B.n217 B.n72 585
R205 B.n216 B.n215 585
R206 B.n214 B.n73 585
R207 B.n213 B.n212 585
R208 B.n160 B.n95 585
R209 B.n162 B.n161 585
R210 B.n163 B.n94 585
R211 B.n165 B.n164 585
R212 B.n166 B.n93 585
R213 B.n168 B.n167 585
R214 B.n169 B.n92 585
R215 B.n171 B.n170 585
R216 B.n172 B.n91 585
R217 B.n174 B.n173 585
R218 B.n175 B.n90 585
R219 B.n177 B.n176 585
R220 B.n179 B.n178 585
R221 B.n180 B.n86 585
R222 B.n182 B.n181 585
R223 B.n183 B.n85 585
R224 B.n185 B.n184 585
R225 B.n186 B.n84 585
R226 B.n188 B.n187 585
R227 B.n189 B.n83 585
R228 B.n191 B.n190 585
R229 B.n192 B.n80 585
R230 B.n195 B.n194 585
R231 B.n196 B.n79 585
R232 B.n198 B.n197 585
R233 B.n199 B.n78 585
R234 B.n201 B.n200 585
R235 B.n202 B.n77 585
R236 B.n204 B.n203 585
R237 B.n205 B.n76 585
R238 B.n207 B.n206 585
R239 B.n208 B.n75 585
R240 B.n210 B.n209 585
R241 B.n211 B.n74 585
R242 B.n159 B.n158 585
R243 B.n157 B.n96 585
R244 B.n156 B.n155 585
R245 B.n154 B.n97 585
R246 B.n153 B.n152 585
R247 B.n151 B.n98 585
R248 B.n150 B.n149 585
R249 B.n148 B.n99 585
R250 B.n147 B.n146 585
R251 B.n145 B.n100 585
R252 B.n144 B.n143 585
R253 B.n142 B.n101 585
R254 B.n141 B.n140 585
R255 B.n139 B.n102 585
R256 B.n138 B.n137 585
R257 B.n136 B.n103 585
R258 B.n135 B.n134 585
R259 B.n133 B.n104 585
R260 B.n132 B.n131 585
R261 B.n130 B.n105 585
R262 B.n129 B.n128 585
R263 B.n127 B.n106 585
R264 B.n126 B.n125 585
R265 B.n124 B.n107 585
R266 B.n123 B.n122 585
R267 B.n121 B.n108 585
R268 B.n120 B.n119 585
R269 B.n118 B.n109 585
R270 B.n117 B.n116 585
R271 B.n115 B.n110 585
R272 B.n114 B.n113 585
R273 B.n112 B.n111 585
R274 B.n2 B.n0 585
R275 B.n413 B.n1 585
R276 B.n412 B.n411 585
R277 B.n410 B.n3 585
R278 B.n409 B.n408 585
R279 B.n407 B.n4 585
R280 B.n406 B.n405 585
R281 B.n404 B.n5 585
R282 B.n403 B.n402 585
R283 B.n401 B.n6 585
R284 B.n400 B.n399 585
R285 B.n398 B.n7 585
R286 B.n397 B.n396 585
R287 B.n395 B.n8 585
R288 B.n394 B.n393 585
R289 B.n392 B.n9 585
R290 B.n391 B.n390 585
R291 B.n389 B.n10 585
R292 B.n388 B.n387 585
R293 B.n386 B.n11 585
R294 B.n385 B.n384 585
R295 B.n383 B.n12 585
R296 B.n382 B.n381 585
R297 B.n380 B.n13 585
R298 B.n379 B.n378 585
R299 B.n377 B.n14 585
R300 B.n376 B.n375 585
R301 B.n374 B.n15 585
R302 B.n373 B.n372 585
R303 B.n371 B.n16 585
R304 B.n370 B.n369 585
R305 B.n368 B.n17 585
R306 B.n367 B.n366 585
R307 B.n365 B.n18 585
R308 B.n415 B.n414 585
R309 B.n160 B.n159 506.916
R310 B.n365 B.n364 506.916
R311 B.n213 B.n74 506.916
R312 B.n311 B.n40 506.916
R313 B.n81 B.t8 330.762
R314 B.n33 B.t4 330.762
R315 B.n87 B.t2 330.762
R316 B.n26 B.t10 330.762
R317 B.n82 B.t7 248.726
R318 B.n34 B.t5 248.726
R319 B.n88 B.t1 248.726
R320 B.n27 B.t11 248.726
R321 B.n81 B.t6 209.764
R322 B.n87 B.t0 209.764
R323 B.n26 B.t9 209.764
R324 B.n33 B.t3 209.764
R325 B.n159 B.n96 163.367
R326 B.n155 B.n96 163.367
R327 B.n155 B.n154 163.367
R328 B.n154 B.n153 163.367
R329 B.n153 B.n98 163.367
R330 B.n149 B.n98 163.367
R331 B.n149 B.n148 163.367
R332 B.n148 B.n147 163.367
R333 B.n147 B.n100 163.367
R334 B.n143 B.n100 163.367
R335 B.n143 B.n142 163.367
R336 B.n142 B.n141 163.367
R337 B.n141 B.n102 163.367
R338 B.n137 B.n102 163.367
R339 B.n137 B.n136 163.367
R340 B.n136 B.n135 163.367
R341 B.n135 B.n104 163.367
R342 B.n131 B.n104 163.367
R343 B.n131 B.n130 163.367
R344 B.n130 B.n129 163.367
R345 B.n129 B.n106 163.367
R346 B.n125 B.n106 163.367
R347 B.n125 B.n124 163.367
R348 B.n124 B.n123 163.367
R349 B.n123 B.n108 163.367
R350 B.n119 B.n108 163.367
R351 B.n119 B.n118 163.367
R352 B.n118 B.n117 163.367
R353 B.n117 B.n110 163.367
R354 B.n113 B.n110 163.367
R355 B.n113 B.n112 163.367
R356 B.n112 B.n2 163.367
R357 B.n414 B.n2 163.367
R358 B.n414 B.n413 163.367
R359 B.n413 B.n412 163.367
R360 B.n412 B.n3 163.367
R361 B.n408 B.n3 163.367
R362 B.n408 B.n407 163.367
R363 B.n407 B.n406 163.367
R364 B.n406 B.n5 163.367
R365 B.n402 B.n5 163.367
R366 B.n402 B.n401 163.367
R367 B.n401 B.n400 163.367
R368 B.n400 B.n7 163.367
R369 B.n396 B.n7 163.367
R370 B.n396 B.n395 163.367
R371 B.n395 B.n394 163.367
R372 B.n394 B.n9 163.367
R373 B.n390 B.n9 163.367
R374 B.n390 B.n389 163.367
R375 B.n389 B.n388 163.367
R376 B.n388 B.n11 163.367
R377 B.n384 B.n11 163.367
R378 B.n384 B.n383 163.367
R379 B.n383 B.n382 163.367
R380 B.n382 B.n13 163.367
R381 B.n378 B.n13 163.367
R382 B.n378 B.n377 163.367
R383 B.n377 B.n376 163.367
R384 B.n376 B.n15 163.367
R385 B.n372 B.n15 163.367
R386 B.n372 B.n371 163.367
R387 B.n371 B.n370 163.367
R388 B.n370 B.n17 163.367
R389 B.n366 B.n17 163.367
R390 B.n366 B.n365 163.367
R391 B.n161 B.n160 163.367
R392 B.n161 B.n94 163.367
R393 B.n165 B.n94 163.367
R394 B.n166 B.n165 163.367
R395 B.n167 B.n166 163.367
R396 B.n167 B.n92 163.367
R397 B.n171 B.n92 163.367
R398 B.n172 B.n171 163.367
R399 B.n173 B.n172 163.367
R400 B.n173 B.n90 163.367
R401 B.n177 B.n90 163.367
R402 B.n178 B.n177 163.367
R403 B.n178 B.n86 163.367
R404 B.n182 B.n86 163.367
R405 B.n183 B.n182 163.367
R406 B.n184 B.n183 163.367
R407 B.n184 B.n84 163.367
R408 B.n188 B.n84 163.367
R409 B.n189 B.n188 163.367
R410 B.n190 B.n189 163.367
R411 B.n190 B.n80 163.367
R412 B.n195 B.n80 163.367
R413 B.n196 B.n195 163.367
R414 B.n197 B.n196 163.367
R415 B.n197 B.n78 163.367
R416 B.n201 B.n78 163.367
R417 B.n202 B.n201 163.367
R418 B.n203 B.n202 163.367
R419 B.n203 B.n76 163.367
R420 B.n207 B.n76 163.367
R421 B.n208 B.n207 163.367
R422 B.n209 B.n208 163.367
R423 B.n209 B.n74 163.367
R424 B.n214 B.n213 163.367
R425 B.n215 B.n214 163.367
R426 B.n215 B.n72 163.367
R427 B.n219 B.n72 163.367
R428 B.n220 B.n219 163.367
R429 B.n221 B.n220 163.367
R430 B.n221 B.n70 163.367
R431 B.n225 B.n70 163.367
R432 B.n226 B.n225 163.367
R433 B.n227 B.n226 163.367
R434 B.n227 B.n68 163.367
R435 B.n231 B.n68 163.367
R436 B.n232 B.n231 163.367
R437 B.n233 B.n232 163.367
R438 B.n233 B.n66 163.367
R439 B.n237 B.n66 163.367
R440 B.n238 B.n237 163.367
R441 B.n239 B.n238 163.367
R442 B.n239 B.n64 163.367
R443 B.n243 B.n64 163.367
R444 B.n244 B.n243 163.367
R445 B.n245 B.n244 163.367
R446 B.n245 B.n62 163.367
R447 B.n249 B.n62 163.367
R448 B.n250 B.n249 163.367
R449 B.n251 B.n250 163.367
R450 B.n251 B.n60 163.367
R451 B.n255 B.n60 163.367
R452 B.n256 B.n255 163.367
R453 B.n257 B.n256 163.367
R454 B.n257 B.n58 163.367
R455 B.n261 B.n58 163.367
R456 B.n262 B.n261 163.367
R457 B.n263 B.n262 163.367
R458 B.n263 B.n56 163.367
R459 B.n267 B.n56 163.367
R460 B.n268 B.n267 163.367
R461 B.n269 B.n268 163.367
R462 B.n269 B.n54 163.367
R463 B.n273 B.n54 163.367
R464 B.n274 B.n273 163.367
R465 B.n275 B.n274 163.367
R466 B.n275 B.n52 163.367
R467 B.n279 B.n52 163.367
R468 B.n280 B.n279 163.367
R469 B.n281 B.n280 163.367
R470 B.n281 B.n50 163.367
R471 B.n285 B.n50 163.367
R472 B.n286 B.n285 163.367
R473 B.n287 B.n286 163.367
R474 B.n287 B.n48 163.367
R475 B.n291 B.n48 163.367
R476 B.n292 B.n291 163.367
R477 B.n293 B.n292 163.367
R478 B.n293 B.n46 163.367
R479 B.n297 B.n46 163.367
R480 B.n298 B.n297 163.367
R481 B.n299 B.n298 163.367
R482 B.n299 B.n44 163.367
R483 B.n303 B.n44 163.367
R484 B.n304 B.n303 163.367
R485 B.n305 B.n304 163.367
R486 B.n305 B.n42 163.367
R487 B.n309 B.n42 163.367
R488 B.n310 B.n309 163.367
R489 B.n311 B.n310 163.367
R490 B.n364 B.n19 163.367
R491 B.n360 B.n19 163.367
R492 B.n360 B.n359 163.367
R493 B.n359 B.n358 163.367
R494 B.n358 B.n21 163.367
R495 B.n354 B.n21 163.367
R496 B.n354 B.n353 163.367
R497 B.n353 B.n352 163.367
R498 B.n352 B.n23 163.367
R499 B.n348 B.n23 163.367
R500 B.n348 B.n347 163.367
R501 B.n347 B.n346 163.367
R502 B.n346 B.n25 163.367
R503 B.n342 B.n25 163.367
R504 B.n342 B.n341 163.367
R505 B.n341 B.n340 163.367
R506 B.n340 B.n30 163.367
R507 B.n336 B.n30 163.367
R508 B.n336 B.n335 163.367
R509 B.n335 B.n334 163.367
R510 B.n334 B.n32 163.367
R511 B.n329 B.n32 163.367
R512 B.n329 B.n328 163.367
R513 B.n328 B.n327 163.367
R514 B.n327 B.n36 163.367
R515 B.n323 B.n36 163.367
R516 B.n323 B.n322 163.367
R517 B.n322 B.n321 163.367
R518 B.n321 B.n38 163.367
R519 B.n317 B.n38 163.367
R520 B.n317 B.n316 163.367
R521 B.n316 B.n315 163.367
R522 B.n315 B.n40 163.367
R523 B.n82 B.n81 82.0369
R524 B.n88 B.n87 82.0369
R525 B.n27 B.n26 82.0369
R526 B.n34 B.n33 82.0369
R527 B.n193 B.n82 59.5399
R528 B.n89 B.n88 59.5399
R529 B.n28 B.n27 59.5399
R530 B.n331 B.n34 59.5399
R531 B.n363 B.n18 32.9371
R532 B.n313 B.n312 32.9371
R533 B.n212 B.n211 32.9371
R534 B.n158 B.n95 32.9371
R535 B B.n415 18.0485
R536 B.n363 B.n362 10.6151
R537 B.n362 B.n361 10.6151
R538 B.n361 B.n20 10.6151
R539 B.n357 B.n20 10.6151
R540 B.n357 B.n356 10.6151
R541 B.n356 B.n355 10.6151
R542 B.n355 B.n22 10.6151
R543 B.n351 B.n22 10.6151
R544 B.n351 B.n350 10.6151
R545 B.n350 B.n349 10.6151
R546 B.n349 B.n24 10.6151
R547 B.n345 B.n344 10.6151
R548 B.n344 B.n343 10.6151
R549 B.n343 B.n29 10.6151
R550 B.n339 B.n29 10.6151
R551 B.n339 B.n338 10.6151
R552 B.n338 B.n337 10.6151
R553 B.n337 B.n31 10.6151
R554 B.n333 B.n31 10.6151
R555 B.n333 B.n332 10.6151
R556 B.n330 B.n35 10.6151
R557 B.n326 B.n35 10.6151
R558 B.n326 B.n325 10.6151
R559 B.n325 B.n324 10.6151
R560 B.n324 B.n37 10.6151
R561 B.n320 B.n37 10.6151
R562 B.n320 B.n319 10.6151
R563 B.n319 B.n318 10.6151
R564 B.n318 B.n39 10.6151
R565 B.n314 B.n39 10.6151
R566 B.n314 B.n313 10.6151
R567 B.n212 B.n73 10.6151
R568 B.n216 B.n73 10.6151
R569 B.n217 B.n216 10.6151
R570 B.n218 B.n217 10.6151
R571 B.n218 B.n71 10.6151
R572 B.n222 B.n71 10.6151
R573 B.n223 B.n222 10.6151
R574 B.n224 B.n223 10.6151
R575 B.n224 B.n69 10.6151
R576 B.n228 B.n69 10.6151
R577 B.n229 B.n228 10.6151
R578 B.n230 B.n229 10.6151
R579 B.n230 B.n67 10.6151
R580 B.n234 B.n67 10.6151
R581 B.n235 B.n234 10.6151
R582 B.n236 B.n235 10.6151
R583 B.n236 B.n65 10.6151
R584 B.n240 B.n65 10.6151
R585 B.n241 B.n240 10.6151
R586 B.n242 B.n241 10.6151
R587 B.n242 B.n63 10.6151
R588 B.n246 B.n63 10.6151
R589 B.n247 B.n246 10.6151
R590 B.n248 B.n247 10.6151
R591 B.n248 B.n61 10.6151
R592 B.n252 B.n61 10.6151
R593 B.n253 B.n252 10.6151
R594 B.n254 B.n253 10.6151
R595 B.n254 B.n59 10.6151
R596 B.n258 B.n59 10.6151
R597 B.n259 B.n258 10.6151
R598 B.n260 B.n259 10.6151
R599 B.n260 B.n57 10.6151
R600 B.n264 B.n57 10.6151
R601 B.n265 B.n264 10.6151
R602 B.n266 B.n265 10.6151
R603 B.n266 B.n55 10.6151
R604 B.n270 B.n55 10.6151
R605 B.n271 B.n270 10.6151
R606 B.n272 B.n271 10.6151
R607 B.n272 B.n53 10.6151
R608 B.n276 B.n53 10.6151
R609 B.n277 B.n276 10.6151
R610 B.n278 B.n277 10.6151
R611 B.n278 B.n51 10.6151
R612 B.n282 B.n51 10.6151
R613 B.n283 B.n282 10.6151
R614 B.n284 B.n283 10.6151
R615 B.n284 B.n49 10.6151
R616 B.n288 B.n49 10.6151
R617 B.n289 B.n288 10.6151
R618 B.n290 B.n289 10.6151
R619 B.n290 B.n47 10.6151
R620 B.n294 B.n47 10.6151
R621 B.n295 B.n294 10.6151
R622 B.n296 B.n295 10.6151
R623 B.n296 B.n45 10.6151
R624 B.n300 B.n45 10.6151
R625 B.n301 B.n300 10.6151
R626 B.n302 B.n301 10.6151
R627 B.n302 B.n43 10.6151
R628 B.n306 B.n43 10.6151
R629 B.n307 B.n306 10.6151
R630 B.n308 B.n307 10.6151
R631 B.n308 B.n41 10.6151
R632 B.n312 B.n41 10.6151
R633 B.n162 B.n95 10.6151
R634 B.n163 B.n162 10.6151
R635 B.n164 B.n163 10.6151
R636 B.n164 B.n93 10.6151
R637 B.n168 B.n93 10.6151
R638 B.n169 B.n168 10.6151
R639 B.n170 B.n169 10.6151
R640 B.n170 B.n91 10.6151
R641 B.n174 B.n91 10.6151
R642 B.n175 B.n174 10.6151
R643 B.n176 B.n175 10.6151
R644 B.n180 B.n179 10.6151
R645 B.n181 B.n180 10.6151
R646 B.n181 B.n85 10.6151
R647 B.n185 B.n85 10.6151
R648 B.n186 B.n185 10.6151
R649 B.n187 B.n186 10.6151
R650 B.n187 B.n83 10.6151
R651 B.n191 B.n83 10.6151
R652 B.n192 B.n191 10.6151
R653 B.n194 B.n79 10.6151
R654 B.n198 B.n79 10.6151
R655 B.n199 B.n198 10.6151
R656 B.n200 B.n199 10.6151
R657 B.n200 B.n77 10.6151
R658 B.n204 B.n77 10.6151
R659 B.n205 B.n204 10.6151
R660 B.n206 B.n205 10.6151
R661 B.n206 B.n75 10.6151
R662 B.n210 B.n75 10.6151
R663 B.n211 B.n210 10.6151
R664 B.n158 B.n157 10.6151
R665 B.n157 B.n156 10.6151
R666 B.n156 B.n97 10.6151
R667 B.n152 B.n97 10.6151
R668 B.n152 B.n151 10.6151
R669 B.n151 B.n150 10.6151
R670 B.n150 B.n99 10.6151
R671 B.n146 B.n99 10.6151
R672 B.n146 B.n145 10.6151
R673 B.n145 B.n144 10.6151
R674 B.n144 B.n101 10.6151
R675 B.n140 B.n101 10.6151
R676 B.n140 B.n139 10.6151
R677 B.n139 B.n138 10.6151
R678 B.n138 B.n103 10.6151
R679 B.n134 B.n103 10.6151
R680 B.n134 B.n133 10.6151
R681 B.n133 B.n132 10.6151
R682 B.n132 B.n105 10.6151
R683 B.n128 B.n105 10.6151
R684 B.n128 B.n127 10.6151
R685 B.n127 B.n126 10.6151
R686 B.n126 B.n107 10.6151
R687 B.n122 B.n107 10.6151
R688 B.n122 B.n121 10.6151
R689 B.n121 B.n120 10.6151
R690 B.n120 B.n109 10.6151
R691 B.n116 B.n109 10.6151
R692 B.n116 B.n115 10.6151
R693 B.n115 B.n114 10.6151
R694 B.n114 B.n111 10.6151
R695 B.n111 B.n0 10.6151
R696 B.n411 B.n1 10.6151
R697 B.n411 B.n410 10.6151
R698 B.n410 B.n409 10.6151
R699 B.n409 B.n4 10.6151
R700 B.n405 B.n4 10.6151
R701 B.n405 B.n404 10.6151
R702 B.n404 B.n403 10.6151
R703 B.n403 B.n6 10.6151
R704 B.n399 B.n6 10.6151
R705 B.n399 B.n398 10.6151
R706 B.n398 B.n397 10.6151
R707 B.n397 B.n8 10.6151
R708 B.n393 B.n8 10.6151
R709 B.n393 B.n392 10.6151
R710 B.n392 B.n391 10.6151
R711 B.n391 B.n10 10.6151
R712 B.n387 B.n10 10.6151
R713 B.n387 B.n386 10.6151
R714 B.n386 B.n385 10.6151
R715 B.n385 B.n12 10.6151
R716 B.n381 B.n12 10.6151
R717 B.n381 B.n380 10.6151
R718 B.n380 B.n379 10.6151
R719 B.n379 B.n14 10.6151
R720 B.n375 B.n14 10.6151
R721 B.n375 B.n374 10.6151
R722 B.n374 B.n373 10.6151
R723 B.n373 B.n16 10.6151
R724 B.n369 B.n16 10.6151
R725 B.n369 B.n368 10.6151
R726 B.n368 B.n367 10.6151
R727 B.n367 B.n18 10.6151
R728 B.n28 B.n24 9.36635
R729 B.n331 B.n330 9.36635
R730 B.n176 B.n89 9.36635
R731 B.n194 B.n193 9.36635
R732 B.n415 B.n0 2.81026
R733 B.n415 B.n1 2.81026
R734 B.n345 B.n28 1.24928
R735 B.n332 B.n331 1.24928
R736 B.n179 B.n89 1.24928
R737 B.n193 B.n192 1.24928
C0 VN VDD1 0.154652f
C1 VDD2 VDD1 0.819908f
C2 VN B 1.09767f
C3 VDD2 B 1.10987f
C4 VN w_n2662_n1372# 3.59656f
C5 VDD2 w_n2662_n1372# 1.28188f
C6 VTAIL VP 1.18021f
C7 VTAIL VDD1 2.86017f
C8 VTAIL B 1.59378f
C9 VP VDD1 0.950138f
C10 VP B 1.66423f
C11 VTAIL w_n2662_n1372# 1.39609f
C12 VP w_n2662_n1372# 3.93395f
C13 VN VDD2 0.712636f
C14 B VDD1 1.06761f
C15 w_n2662_n1372# VDD1 1.24073f
C16 w_n2662_n1372# B 7.4709f
C17 VTAIL VN 1.16597f
C18 VTAIL VDD2 2.92202f
C19 VN VP 4.22932f
C20 VDD2 VP 0.393783f
C21 VDD2 VSUBS 0.685639f
C22 VDD1 VSUBS 2.652063f
C23 VTAIL VSUBS 0.419733f
C24 VN VSUBS 6.29425f
C25 VP VSUBS 1.591953f
C26 B VSUBS 3.798789f
C27 w_n2662_n1372# VSUBS 46.6063f
C28 B.n0 VSUBS 0.005921f
C29 B.n1 VSUBS 0.005921f
C30 B.n2 VSUBS 0.009364f
C31 B.n3 VSUBS 0.009364f
C32 B.n4 VSUBS 0.009364f
C33 B.n5 VSUBS 0.009364f
C34 B.n6 VSUBS 0.009364f
C35 B.n7 VSUBS 0.009364f
C36 B.n8 VSUBS 0.009364f
C37 B.n9 VSUBS 0.009364f
C38 B.n10 VSUBS 0.009364f
C39 B.n11 VSUBS 0.009364f
C40 B.n12 VSUBS 0.009364f
C41 B.n13 VSUBS 0.009364f
C42 B.n14 VSUBS 0.009364f
C43 B.n15 VSUBS 0.009364f
C44 B.n16 VSUBS 0.009364f
C45 B.n17 VSUBS 0.009364f
C46 B.n18 VSUBS 0.021564f
C47 B.n19 VSUBS 0.009364f
C48 B.n20 VSUBS 0.009364f
C49 B.n21 VSUBS 0.009364f
C50 B.n22 VSUBS 0.009364f
C51 B.n23 VSUBS 0.009364f
C52 B.n24 VSUBS 0.008813f
C53 B.n25 VSUBS 0.009364f
C54 B.t11 VSUBS 0.046074f
C55 B.t10 VSUBS 0.066972f
C56 B.t9 VSUBS 0.529111f
C57 B.n26 VSUBS 0.117619f
C58 B.n27 VSUBS 0.097615f
C59 B.n28 VSUBS 0.021694f
C60 B.n29 VSUBS 0.009364f
C61 B.n30 VSUBS 0.009364f
C62 B.n31 VSUBS 0.009364f
C63 B.n32 VSUBS 0.009364f
C64 B.t5 VSUBS 0.046074f
C65 B.t4 VSUBS 0.066972f
C66 B.t3 VSUBS 0.529111f
C67 B.n33 VSUBS 0.117619f
C68 B.n34 VSUBS 0.097615f
C69 B.n35 VSUBS 0.009364f
C70 B.n36 VSUBS 0.009364f
C71 B.n37 VSUBS 0.009364f
C72 B.n38 VSUBS 0.009364f
C73 B.n39 VSUBS 0.009364f
C74 B.n40 VSUBS 0.0225f
C75 B.n41 VSUBS 0.009364f
C76 B.n42 VSUBS 0.009364f
C77 B.n43 VSUBS 0.009364f
C78 B.n44 VSUBS 0.009364f
C79 B.n45 VSUBS 0.009364f
C80 B.n46 VSUBS 0.009364f
C81 B.n47 VSUBS 0.009364f
C82 B.n48 VSUBS 0.009364f
C83 B.n49 VSUBS 0.009364f
C84 B.n50 VSUBS 0.009364f
C85 B.n51 VSUBS 0.009364f
C86 B.n52 VSUBS 0.009364f
C87 B.n53 VSUBS 0.009364f
C88 B.n54 VSUBS 0.009364f
C89 B.n55 VSUBS 0.009364f
C90 B.n56 VSUBS 0.009364f
C91 B.n57 VSUBS 0.009364f
C92 B.n58 VSUBS 0.009364f
C93 B.n59 VSUBS 0.009364f
C94 B.n60 VSUBS 0.009364f
C95 B.n61 VSUBS 0.009364f
C96 B.n62 VSUBS 0.009364f
C97 B.n63 VSUBS 0.009364f
C98 B.n64 VSUBS 0.009364f
C99 B.n65 VSUBS 0.009364f
C100 B.n66 VSUBS 0.009364f
C101 B.n67 VSUBS 0.009364f
C102 B.n68 VSUBS 0.009364f
C103 B.n69 VSUBS 0.009364f
C104 B.n70 VSUBS 0.009364f
C105 B.n71 VSUBS 0.009364f
C106 B.n72 VSUBS 0.009364f
C107 B.n73 VSUBS 0.009364f
C108 B.n74 VSUBS 0.0225f
C109 B.n75 VSUBS 0.009364f
C110 B.n76 VSUBS 0.009364f
C111 B.n77 VSUBS 0.009364f
C112 B.n78 VSUBS 0.009364f
C113 B.n79 VSUBS 0.009364f
C114 B.n80 VSUBS 0.009364f
C115 B.t7 VSUBS 0.046074f
C116 B.t8 VSUBS 0.066972f
C117 B.t6 VSUBS 0.529111f
C118 B.n81 VSUBS 0.117619f
C119 B.n82 VSUBS 0.097615f
C120 B.n83 VSUBS 0.009364f
C121 B.n84 VSUBS 0.009364f
C122 B.n85 VSUBS 0.009364f
C123 B.n86 VSUBS 0.009364f
C124 B.t1 VSUBS 0.046074f
C125 B.t2 VSUBS 0.066972f
C126 B.t0 VSUBS 0.529111f
C127 B.n87 VSUBS 0.117619f
C128 B.n88 VSUBS 0.097615f
C129 B.n89 VSUBS 0.021694f
C130 B.n90 VSUBS 0.009364f
C131 B.n91 VSUBS 0.009364f
C132 B.n92 VSUBS 0.009364f
C133 B.n93 VSUBS 0.009364f
C134 B.n94 VSUBS 0.009364f
C135 B.n95 VSUBS 0.0225f
C136 B.n96 VSUBS 0.009364f
C137 B.n97 VSUBS 0.009364f
C138 B.n98 VSUBS 0.009364f
C139 B.n99 VSUBS 0.009364f
C140 B.n100 VSUBS 0.009364f
C141 B.n101 VSUBS 0.009364f
C142 B.n102 VSUBS 0.009364f
C143 B.n103 VSUBS 0.009364f
C144 B.n104 VSUBS 0.009364f
C145 B.n105 VSUBS 0.009364f
C146 B.n106 VSUBS 0.009364f
C147 B.n107 VSUBS 0.009364f
C148 B.n108 VSUBS 0.009364f
C149 B.n109 VSUBS 0.009364f
C150 B.n110 VSUBS 0.009364f
C151 B.n111 VSUBS 0.009364f
C152 B.n112 VSUBS 0.009364f
C153 B.n113 VSUBS 0.009364f
C154 B.n114 VSUBS 0.009364f
C155 B.n115 VSUBS 0.009364f
C156 B.n116 VSUBS 0.009364f
C157 B.n117 VSUBS 0.009364f
C158 B.n118 VSUBS 0.009364f
C159 B.n119 VSUBS 0.009364f
C160 B.n120 VSUBS 0.009364f
C161 B.n121 VSUBS 0.009364f
C162 B.n122 VSUBS 0.009364f
C163 B.n123 VSUBS 0.009364f
C164 B.n124 VSUBS 0.009364f
C165 B.n125 VSUBS 0.009364f
C166 B.n126 VSUBS 0.009364f
C167 B.n127 VSUBS 0.009364f
C168 B.n128 VSUBS 0.009364f
C169 B.n129 VSUBS 0.009364f
C170 B.n130 VSUBS 0.009364f
C171 B.n131 VSUBS 0.009364f
C172 B.n132 VSUBS 0.009364f
C173 B.n133 VSUBS 0.009364f
C174 B.n134 VSUBS 0.009364f
C175 B.n135 VSUBS 0.009364f
C176 B.n136 VSUBS 0.009364f
C177 B.n137 VSUBS 0.009364f
C178 B.n138 VSUBS 0.009364f
C179 B.n139 VSUBS 0.009364f
C180 B.n140 VSUBS 0.009364f
C181 B.n141 VSUBS 0.009364f
C182 B.n142 VSUBS 0.009364f
C183 B.n143 VSUBS 0.009364f
C184 B.n144 VSUBS 0.009364f
C185 B.n145 VSUBS 0.009364f
C186 B.n146 VSUBS 0.009364f
C187 B.n147 VSUBS 0.009364f
C188 B.n148 VSUBS 0.009364f
C189 B.n149 VSUBS 0.009364f
C190 B.n150 VSUBS 0.009364f
C191 B.n151 VSUBS 0.009364f
C192 B.n152 VSUBS 0.009364f
C193 B.n153 VSUBS 0.009364f
C194 B.n154 VSUBS 0.009364f
C195 B.n155 VSUBS 0.009364f
C196 B.n156 VSUBS 0.009364f
C197 B.n157 VSUBS 0.009364f
C198 B.n158 VSUBS 0.021564f
C199 B.n159 VSUBS 0.021564f
C200 B.n160 VSUBS 0.0225f
C201 B.n161 VSUBS 0.009364f
C202 B.n162 VSUBS 0.009364f
C203 B.n163 VSUBS 0.009364f
C204 B.n164 VSUBS 0.009364f
C205 B.n165 VSUBS 0.009364f
C206 B.n166 VSUBS 0.009364f
C207 B.n167 VSUBS 0.009364f
C208 B.n168 VSUBS 0.009364f
C209 B.n169 VSUBS 0.009364f
C210 B.n170 VSUBS 0.009364f
C211 B.n171 VSUBS 0.009364f
C212 B.n172 VSUBS 0.009364f
C213 B.n173 VSUBS 0.009364f
C214 B.n174 VSUBS 0.009364f
C215 B.n175 VSUBS 0.009364f
C216 B.n176 VSUBS 0.008813f
C217 B.n177 VSUBS 0.009364f
C218 B.n178 VSUBS 0.009364f
C219 B.n179 VSUBS 0.005233f
C220 B.n180 VSUBS 0.009364f
C221 B.n181 VSUBS 0.009364f
C222 B.n182 VSUBS 0.009364f
C223 B.n183 VSUBS 0.009364f
C224 B.n184 VSUBS 0.009364f
C225 B.n185 VSUBS 0.009364f
C226 B.n186 VSUBS 0.009364f
C227 B.n187 VSUBS 0.009364f
C228 B.n188 VSUBS 0.009364f
C229 B.n189 VSUBS 0.009364f
C230 B.n190 VSUBS 0.009364f
C231 B.n191 VSUBS 0.009364f
C232 B.n192 VSUBS 0.005233f
C233 B.n193 VSUBS 0.021694f
C234 B.n194 VSUBS 0.008813f
C235 B.n195 VSUBS 0.009364f
C236 B.n196 VSUBS 0.009364f
C237 B.n197 VSUBS 0.009364f
C238 B.n198 VSUBS 0.009364f
C239 B.n199 VSUBS 0.009364f
C240 B.n200 VSUBS 0.009364f
C241 B.n201 VSUBS 0.009364f
C242 B.n202 VSUBS 0.009364f
C243 B.n203 VSUBS 0.009364f
C244 B.n204 VSUBS 0.009364f
C245 B.n205 VSUBS 0.009364f
C246 B.n206 VSUBS 0.009364f
C247 B.n207 VSUBS 0.009364f
C248 B.n208 VSUBS 0.009364f
C249 B.n209 VSUBS 0.009364f
C250 B.n210 VSUBS 0.009364f
C251 B.n211 VSUBS 0.0225f
C252 B.n212 VSUBS 0.021564f
C253 B.n213 VSUBS 0.021564f
C254 B.n214 VSUBS 0.009364f
C255 B.n215 VSUBS 0.009364f
C256 B.n216 VSUBS 0.009364f
C257 B.n217 VSUBS 0.009364f
C258 B.n218 VSUBS 0.009364f
C259 B.n219 VSUBS 0.009364f
C260 B.n220 VSUBS 0.009364f
C261 B.n221 VSUBS 0.009364f
C262 B.n222 VSUBS 0.009364f
C263 B.n223 VSUBS 0.009364f
C264 B.n224 VSUBS 0.009364f
C265 B.n225 VSUBS 0.009364f
C266 B.n226 VSUBS 0.009364f
C267 B.n227 VSUBS 0.009364f
C268 B.n228 VSUBS 0.009364f
C269 B.n229 VSUBS 0.009364f
C270 B.n230 VSUBS 0.009364f
C271 B.n231 VSUBS 0.009364f
C272 B.n232 VSUBS 0.009364f
C273 B.n233 VSUBS 0.009364f
C274 B.n234 VSUBS 0.009364f
C275 B.n235 VSUBS 0.009364f
C276 B.n236 VSUBS 0.009364f
C277 B.n237 VSUBS 0.009364f
C278 B.n238 VSUBS 0.009364f
C279 B.n239 VSUBS 0.009364f
C280 B.n240 VSUBS 0.009364f
C281 B.n241 VSUBS 0.009364f
C282 B.n242 VSUBS 0.009364f
C283 B.n243 VSUBS 0.009364f
C284 B.n244 VSUBS 0.009364f
C285 B.n245 VSUBS 0.009364f
C286 B.n246 VSUBS 0.009364f
C287 B.n247 VSUBS 0.009364f
C288 B.n248 VSUBS 0.009364f
C289 B.n249 VSUBS 0.009364f
C290 B.n250 VSUBS 0.009364f
C291 B.n251 VSUBS 0.009364f
C292 B.n252 VSUBS 0.009364f
C293 B.n253 VSUBS 0.009364f
C294 B.n254 VSUBS 0.009364f
C295 B.n255 VSUBS 0.009364f
C296 B.n256 VSUBS 0.009364f
C297 B.n257 VSUBS 0.009364f
C298 B.n258 VSUBS 0.009364f
C299 B.n259 VSUBS 0.009364f
C300 B.n260 VSUBS 0.009364f
C301 B.n261 VSUBS 0.009364f
C302 B.n262 VSUBS 0.009364f
C303 B.n263 VSUBS 0.009364f
C304 B.n264 VSUBS 0.009364f
C305 B.n265 VSUBS 0.009364f
C306 B.n266 VSUBS 0.009364f
C307 B.n267 VSUBS 0.009364f
C308 B.n268 VSUBS 0.009364f
C309 B.n269 VSUBS 0.009364f
C310 B.n270 VSUBS 0.009364f
C311 B.n271 VSUBS 0.009364f
C312 B.n272 VSUBS 0.009364f
C313 B.n273 VSUBS 0.009364f
C314 B.n274 VSUBS 0.009364f
C315 B.n275 VSUBS 0.009364f
C316 B.n276 VSUBS 0.009364f
C317 B.n277 VSUBS 0.009364f
C318 B.n278 VSUBS 0.009364f
C319 B.n279 VSUBS 0.009364f
C320 B.n280 VSUBS 0.009364f
C321 B.n281 VSUBS 0.009364f
C322 B.n282 VSUBS 0.009364f
C323 B.n283 VSUBS 0.009364f
C324 B.n284 VSUBS 0.009364f
C325 B.n285 VSUBS 0.009364f
C326 B.n286 VSUBS 0.009364f
C327 B.n287 VSUBS 0.009364f
C328 B.n288 VSUBS 0.009364f
C329 B.n289 VSUBS 0.009364f
C330 B.n290 VSUBS 0.009364f
C331 B.n291 VSUBS 0.009364f
C332 B.n292 VSUBS 0.009364f
C333 B.n293 VSUBS 0.009364f
C334 B.n294 VSUBS 0.009364f
C335 B.n295 VSUBS 0.009364f
C336 B.n296 VSUBS 0.009364f
C337 B.n297 VSUBS 0.009364f
C338 B.n298 VSUBS 0.009364f
C339 B.n299 VSUBS 0.009364f
C340 B.n300 VSUBS 0.009364f
C341 B.n301 VSUBS 0.009364f
C342 B.n302 VSUBS 0.009364f
C343 B.n303 VSUBS 0.009364f
C344 B.n304 VSUBS 0.009364f
C345 B.n305 VSUBS 0.009364f
C346 B.n306 VSUBS 0.009364f
C347 B.n307 VSUBS 0.009364f
C348 B.n308 VSUBS 0.009364f
C349 B.n309 VSUBS 0.009364f
C350 B.n310 VSUBS 0.009364f
C351 B.n311 VSUBS 0.021564f
C352 B.n312 VSUBS 0.022661f
C353 B.n313 VSUBS 0.021403f
C354 B.n314 VSUBS 0.009364f
C355 B.n315 VSUBS 0.009364f
C356 B.n316 VSUBS 0.009364f
C357 B.n317 VSUBS 0.009364f
C358 B.n318 VSUBS 0.009364f
C359 B.n319 VSUBS 0.009364f
C360 B.n320 VSUBS 0.009364f
C361 B.n321 VSUBS 0.009364f
C362 B.n322 VSUBS 0.009364f
C363 B.n323 VSUBS 0.009364f
C364 B.n324 VSUBS 0.009364f
C365 B.n325 VSUBS 0.009364f
C366 B.n326 VSUBS 0.009364f
C367 B.n327 VSUBS 0.009364f
C368 B.n328 VSUBS 0.009364f
C369 B.n329 VSUBS 0.009364f
C370 B.n330 VSUBS 0.008813f
C371 B.n331 VSUBS 0.021694f
C372 B.n332 VSUBS 0.005233f
C373 B.n333 VSUBS 0.009364f
C374 B.n334 VSUBS 0.009364f
C375 B.n335 VSUBS 0.009364f
C376 B.n336 VSUBS 0.009364f
C377 B.n337 VSUBS 0.009364f
C378 B.n338 VSUBS 0.009364f
C379 B.n339 VSUBS 0.009364f
C380 B.n340 VSUBS 0.009364f
C381 B.n341 VSUBS 0.009364f
C382 B.n342 VSUBS 0.009364f
C383 B.n343 VSUBS 0.009364f
C384 B.n344 VSUBS 0.009364f
C385 B.n345 VSUBS 0.005233f
C386 B.n346 VSUBS 0.009364f
C387 B.n347 VSUBS 0.009364f
C388 B.n348 VSUBS 0.009364f
C389 B.n349 VSUBS 0.009364f
C390 B.n350 VSUBS 0.009364f
C391 B.n351 VSUBS 0.009364f
C392 B.n352 VSUBS 0.009364f
C393 B.n353 VSUBS 0.009364f
C394 B.n354 VSUBS 0.009364f
C395 B.n355 VSUBS 0.009364f
C396 B.n356 VSUBS 0.009364f
C397 B.n357 VSUBS 0.009364f
C398 B.n358 VSUBS 0.009364f
C399 B.n359 VSUBS 0.009364f
C400 B.n360 VSUBS 0.009364f
C401 B.n361 VSUBS 0.009364f
C402 B.n362 VSUBS 0.009364f
C403 B.n363 VSUBS 0.0225f
C404 B.n364 VSUBS 0.0225f
C405 B.n365 VSUBS 0.021564f
C406 B.n366 VSUBS 0.009364f
C407 B.n367 VSUBS 0.009364f
C408 B.n368 VSUBS 0.009364f
C409 B.n369 VSUBS 0.009364f
C410 B.n370 VSUBS 0.009364f
C411 B.n371 VSUBS 0.009364f
C412 B.n372 VSUBS 0.009364f
C413 B.n373 VSUBS 0.009364f
C414 B.n374 VSUBS 0.009364f
C415 B.n375 VSUBS 0.009364f
C416 B.n376 VSUBS 0.009364f
C417 B.n377 VSUBS 0.009364f
C418 B.n378 VSUBS 0.009364f
C419 B.n379 VSUBS 0.009364f
C420 B.n380 VSUBS 0.009364f
C421 B.n381 VSUBS 0.009364f
C422 B.n382 VSUBS 0.009364f
C423 B.n383 VSUBS 0.009364f
C424 B.n384 VSUBS 0.009364f
C425 B.n385 VSUBS 0.009364f
C426 B.n386 VSUBS 0.009364f
C427 B.n387 VSUBS 0.009364f
C428 B.n388 VSUBS 0.009364f
C429 B.n389 VSUBS 0.009364f
C430 B.n390 VSUBS 0.009364f
C431 B.n391 VSUBS 0.009364f
C432 B.n392 VSUBS 0.009364f
C433 B.n393 VSUBS 0.009364f
C434 B.n394 VSUBS 0.009364f
C435 B.n395 VSUBS 0.009364f
C436 B.n396 VSUBS 0.009364f
C437 B.n397 VSUBS 0.009364f
C438 B.n398 VSUBS 0.009364f
C439 B.n399 VSUBS 0.009364f
C440 B.n400 VSUBS 0.009364f
C441 B.n401 VSUBS 0.009364f
C442 B.n402 VSUBS 0.009364f
C443 B.n403 VSUBS 0.009364f
C444 B.n404 VSUBS 0.009364f
C445 B.n405 VSUBS 0.009364f
C446 B.n406 VSUBS 0.009364f
C447 B.n407 VSUBS 0.009364f
C448 B.n408 VSUBS 0.009364f
C449 B.n409 VSUBS 0.009364f
C450 B.n410 VSUBS 0.009364f
C451 B.n411 VSUBS 0.009364f
C452 B.n412 VSUBS 0.009364f
C453 B.n413 VSUBS 0.009364f
C454 B.n414 VSUBS 0.009364f
C455 B.n415 VSUBS 0.021202f
C456 VDD2.n0 VSUBS 0.02093f
C457 VDD2.n1 VSUBS 0.054061f
C458 VDD2.t0 VSUBS 0.054279f
C459 VDD2.n2 VSUBS 0.053152f
C460 VDD2.n3 VSUBS 0.015249f
C461 VDD2.n4 VSUBS 0.009892f
C462 VDD2.n5 VSUBS 0.128795f
C463 VDD2.n6 VSUBS 0.363019f
C464 VDD2.n7 VSUBS 0.02093f
C465 VDD2.n8 VSUBS 0.054061f
C466 VDD2.t1 VSUBS 0.054279f
C467 VDD2.n9 VSUBS 0.053152f
C468 VDD2.n10 VSUBS 0.015249f
C469 VDD2.n11 VSUBS 0.009892f
C470 VDD2.n12 VSUBS 0.128795f
C471 VDD2.n13 VSUBS 0.042475f
C472 VDD2.n14 VSUBS 1.65561f
C473 VN.t1 VSUBS 1.42039f
C474 VN.t0 VSUBS 2.53291f
C475 VDD1.n0 VSUBS 0.020451f
C476 VDD1.n1 VSUBS 0.052822f
C477 VDD1.t0 VSUBS 0.053035f
C478 VDD1.n2 VSUBS 0.051935f
C479 VDD1.n3 VSUBS 0.014899f
C480 VDD1.n4 VSUBS 0.009665f
C481 VDD1.n5 VSUBS 0.125845f
C482 VDD1.n6 VSUBS 0.043278f
C483 VDD1.n7 VSUBS 0.020451f
C484 VDD1.n8 VSUBS 0.052822f
C485 VDD1.t1 VSUBS 0.053035f
C486 VDD1.n9 VSUBS 0.051935f
C487 VDD1.n10 VSUBS 0.014899f
C488 VDD1.n11 VSUBS 0.009665f
C489 VDD1.n12 VSUBS 0.125845f
C490 VDD1.n13 VSUBS 0.390242f
C491 VTAIL.n0 VSUBS 0.025389f
C492 VTAIL.n1 VSUBS 0.065577f
C493 VTAIL.t3 VSUBS 0.065842f
C494 VTAIL.n2 VSUBS 0.064475f
C495 VTAIL.n3 VSUBS 0.018497f
C496 VTAIL.n4 VSUBS 0.011999f
C497 VTAIL.n5 VSUBS 0.156232f
C498 VTAIL.n6 VSUBS 0.0361f
C499 VTAIL.n7 VSUBS 1.07567f
C500 VTAIL.n8 VSUBS 0.025389f
C501 VTAIL.n9 VSUBS 0.065577f
C502 VTAIL.t1 VSUBS 0.065841f
C503 VTAIL.n10 VSUBS 0.064475f
C504 VTAIL.n11 VSUBS 0.018497f
C505 VTAIL.n12 VSUBS 0.011999f
C506 VTAIL.n13 VSUBS 0.156232f
C507 VTAIL.n14 VSUBS 0.0361f
C508 VTAIL.n15 VSUBS 1.13708f
C509 VTAIL.n16 VSUBS 0.025389f
C510 VTAIL.n17 VSUBS 0.065577f
C511 VTAIL.t2 VSUBS 0.065842f
C512 VTAIL.n18 VSUBS 0.064475f
C513 VTAIL.n19 VSUBS 0.018497f
C514 VTAIL.n20 VSUBS 0.011999f
C515 VTAIL.n21 VSUBS 0.156232f
C516 VTAIL.n22 VSUBS 0.0361f
C517 VTAIL.n23 VSUBS 0.874705f
C518 VTAIL.n24 VSUBS 0.025389f
C519 VTAIL.n25 VSUBS 0.065577f
C520 VTAIL.t0 VSUBS 0.065842f
C521 VTAIL.n26 VSUBS 0.064475f
C522 VTAIL.n27 VSUBS 0.018497f
C523 VTAIL.n28 VSUBS 0.011999f
C524 VTAIL.n29 VSUBS 0.156232f
C525 VTAIL.n30 VSUBS 0.0361f
C526 VTAIL.n31 VSUBS 0.77112f
C527 VP.t1 VSUBS 2.65381f
C528 VP.t0 VSUBS 1.47941f
C529 VP.n0 VSUBS 3.75561f
.ends

