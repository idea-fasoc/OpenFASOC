* NGSPICE file created from diff_pair_sample_1771.ext - technology: sky130A

.subckt diff_pair_sample_1771 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1978_n4762# sky130_fd_pr__pfet_01v8 ad=7.3983 pd=38.72 as=0 ps=0 w=18.97 l=1.35
X1 VTAIL.t7 VN.t0 VDD2.t3 w_n1978_n4762# sky130_fd_pr__pfet_01v8 ad=7.3983 pd=38.72 as=3.13005 ps=19.3 w=18.97 l=1.35
X2 VTAIL.t0 VP.t0 VDD1.t3 w_n1978_n4762# sky130_fd_pr__pfet_01v8 ad=7.3983 pd=38.72 as=3.13005 ps=19.3 w=18.97 l=1.35
X3 VDD2.t2 VN.t1 VTAIL.t6 w_n1978_n4762# sky130_fd_pr__pfet_01v8 ad=3.13005 pd=19.3 as=7.3983 ps=38.72 w=18.97 l=1.35
X4 VDD2.t0 VN.t2 VTAIL.t5 w_n1978_n4762# sky130_fd_pr__pfet_01v8 ad=3.13005 pd=19.3 as=7.3983 ps=38.72 w=18.97 l=1.35
X5 VDD1.t2 VP.t1 VTAIL.t2 w_n1978_n4762# sky130_fd_pr__pfet_01v8 ad=3.13005 pd=19.3 as=7.3983 ps=38.72 w=18.97 l=1.35
X6 B.t8 B.t6 B.t7 w_n1978_n4762# sky130_fd_pr__pfet_01v8 ad=7.3983 pd=38.72 as=0 ps=0 w=18.97 l=1.35
X7 VDD1.t1 VP.t2 VTAIL.t3 w_n1978_n4762# sky130_fd_pr__pfet_01v8 ad=3.13005 pd=19.3 as=7.3983 ps=38.72 w=18.97 l=1.35
X8 VTAIL.t1 VP.t3 VDD1.t0 w_n1978_n4762# sky130_fd_pr__pfet_01v8 ad=7.3983 pd=38.72 as=3.13005 ps=19.3 w=18.97 l=1.35
X9 B.t5 B.t3 B.t4 w_n1978_n4762# sky130_fd_pr__pfet_01v8 ad=7.3983 pd=38.72 as=0 ps=0 w=18.97 l=1.35
X10 B.t2 B.t0 B.t1 w_n1978_n4762# sky130_fd_pr__pfet_01v8 ad=7.3983 pd=38.72 as=0 ps=0 w=18.97 l=1.35
X11 VTAIL.t4 VN.t3 VDD2.t1 w_n1978_n4762# sky130_fd_pr__pfet_01v8 ad=7.3983 pd=38.72 as=3.13005 ps=19.3 w=18.97 l=1.35
R0 B.n498 B.n85 585
R1 B.n500 B.n499 585
R2 B.n501 B.n84 585
R3 B.n503 B.n502 585
R4 B.n504 B.n83 585
R5 B.n506 B.n505 585
R6 B.n507 B.n82 585
R7 B.n509 B.n508 585
R8 B.n510 B.n81 585
R9 B.n512 B.n511 585
R10 B.n513 B.n80 585
R11 B.n515 B.n514 585
R12 B.n516 B.n79 585
R13 B.n518 B.n517 585
R14 B.n519 B.n78 585
R15 B.n521 B.n520 585
R16 B.n522 B.n77 585
R17 B.n524 B.n523 585
R18 B.n525 B.n76 585
R19 B.n527 B.n526 585
R20 B.n528 B.n75 585
R21 B.n530 B.n529 585
R22 B.n531 B.n74 585
R23 B.n533 B.n532 585
R24 B.n534 B.n73 585
R25 B.n536 B.n535 585
R26 B.n537 B.n72 585
R27 B.n539 B.n538 585
R28 B.n540 B.n71 585
R29 B.n542 B.n541 585
R30 B.n543 B.n70 585
R31 B.n545 B.n544 585
R32 B.n546 B.n69 585
R33 B.n548 B.n547 585
R34 B.n549 B.n68 585
R35 B.n551 B.n550 585
R36 B.n552 B.n67 585
R37 B.n554 B.n553 585
R38 B.n555 B.n66 585
R39 B.n557 B.n556 585
R40 B.n558 B.n65 585
R41 B.n560 B.n559 585
R42 B.n561 B.n64 585
R43 B.n563 B.n562 585
R44 B.n564 B.n63 585
R45 B.n566 B.n565 585
R46 B.n567 B.n62 585
R47 B.n569 B.n568 585
R48 B.n570 B.n61 585
R49 B.n572 B.n571 585
R50 B.n573 B.n60 585
R51 B.n575 B.n574 585
R52 B.n576 B.n59 585
R53 B.n578 B.n577 585
R54 B.n579 B.n58 585
R55 B.n581 B.n580 585
R56 B.n582 B.n57 585
R57 B.n584 B.n583 585
R58 B.n585 B.n56 585
R59 B.n587 B.n586 585
R60 B.n588 B.n55 585
R61 B.n590 B.n589 585
R62 B.n592 B.n52 585
R63 B.n594 B.n593 585
R64 B.n595 B.n51 585
R65 B.n597 B.n596 585
R66 B.n598 B.n50 585
R67 B.n600 B.n599 585
R68 B.n601 B.n49 585
R69 B.n603 B.n602 585
R70 B.n604 B.n45 585
R71 B.n606 B.n605 585
R72 B.n607 B.n44 585
R73 B.n609 B.n608 585
R74 B.n610 B.n43 585
R75 B.n612 B.n611 585
R76 B.n613 B.n42 585
R77 B.n615 B.n614 585
R78 B.n616 B.n41 585
R79 B.n618 B.n617 585
R80 B.n619 B.n40 585
R81 B.n621 B.n620 585
R82 B.n622 B.n39 585
R83 B.n624 B.n623 585
R84 B.n625 B.n38 585
R85 B.n627 B.n626 585
R86 B.n628 B.n37 585
R87 B.n630 B.n629 585
R88 B.n631 B.n36 585
R89 B.n633 B.n632 585
R90 B.n634 B.n35 585
R91 B.n636 B.n635 585
R92 B.n637 B.n34 585
R93 B.n639 B.n638 585
R94 B.n640 B.n33 585
R95 B.n642 B.n641 585
R96 B.n643 B.n32 585
R97 B.n645 B.n644 585
R98 B.n646 B.n31 585
R99 B.n648 B.n647 585
R100 B.n649 B.n30 585
R101 B.n651 B.n650 585
R102 B.n652 B.n29 585
R103 B.n654 B.n653 585
R104 B.n655 B.n28 585
R105 B.n657 B.n656 585
R106 B.n658 B.n27 585
R107 B.n660 B.n659 585
R108 B.n661 B.n26 585
R109 B.n663 B.n662 585
R110 B.n664 B.n25 585
R111 B.n666 B.n665 585
R112 B.n667 B.n24 585
R113 B.n669 B.n668 585
R114 B.n670 B.n23 585
R115 B.n672 B.n671 585
R116 B.n673 B.n22 585
R117 B.n675 B.n674 585
R118 B.n676 B.n21 585
R119 B.n678 B.n677 585
R120 B.n679 B.n20 585
R121 B.n681 B.n680 585
R122 B.n682 B.n19 585
R123 B.n684 B.n683 585
R124 B.n685 B.n18 585
R125 B.n687 B.n686 585
R126 B.n688 B.n17 585
R127 B.n690 B.n689 585
R128 B.n691 B.n16 585
R129 B.n693 B.n692 585
R130 B.n694 B.n15 585
R131 B.n696 B.n695 585
R132 B.n697 B.n14 585
R133 B.n699 B.n698 585
R134 B.n497 B.n496 585
R135 B.n495 B.n86 585
R136 B.n494 B.n493 585
R137 B.n492 B.n87 585
R138 B.n491 B.n490 585
R139 B.n489 B.n88 585
R140 B.n488 B.n487 585
R141 B.n486 B.n89 585
R142 B.n485 B.n484 585
R143 B.n483 B.n90 585
R144 B.n482 B.n481 585
R145 B.n480 B.n91 585
R146 B.n479 B.n478 585
R147 B.n477 B.n92 585
R148 B.n476 B.n475 585
R149 B.n474 B.n93 585
R150 B.n473 B.n472 585
R151 B.n471 B.n94 585
R152 B.n470 B.n469 585
R153 B.n468 B.n95 585
R154 B.n467 B.n466 585
R155 B.n465 B.n96 585
R156 B.n464 B.n463 585
R157 B.n462 B.n97 585
R158 B.n461 B.n460 585
R159 B.n459 B.n98 585
R160 B.n458 B.n457 585
R161 B.n456 B.n99 585
R162 B.n455 B.n454 585
R163 B.n453 B.n100 585
R164 B.n452 B.n451 585
R165 B.n450 B.n101 585
R166 B.n449 B.n448 585
R167 B.n447 B.n102 585
R168 B.n446 B.n445 585
R169 B.n444 B.n103 585
R170 B.n443 B.n442 585
R171 B.n441 B.n104 585
R172 B.n440 B.n439 585
R173 B.n438 B.n105 585
R174 B.n437 B.n436 585
R175 B.n435 B.n106 585
R176 B.n434 B.n433 585
R177 B.n432 B.n107 585
R178 B.n431 B.n430 585
R179 B.n429 B.n108 585
R180 B.n428 B.n427 585
R181 B.n225 B.n180 585
R182 B.n227 B.n226 585
R183 B.n228 B.n179 585
R184 B.n230 B.n229 585
R185 B.n231 B.n178 585
R186 B.n233 B.n232 585
R187 B.n234 B.n177 585
R188 B.n236 B.n235 585
R189 B.n237 B.n176 585
R190 B.n239 B.n238 585
R191 B.n240 B.n175 585
R192 B.n242 B.n241 585
R193 B.n243 B.n174 585
R194 B.n245 B.n244 585
R195 B.n246 B.n173 585
R196 B.n248 B.n247 585
R197 B.n249 B.n172 585
R198 B.n251 B.n250 585
R199 B.n252 B.n171 585
R200 B.n254 B.n253 585
R201 B.n255 B.n170 585
R202 B.n257 B.n256 585
R203 B.n258 B.n169 585
R204 B.n260 B.n259 585
R205 B.n261 B.n168 585
R206 B.n263 B.n262 585
R207 B.n264 B.n167 585
R208 B.n266 B.n265 585
R209 B.n267 B.n166 585
R210 B.n269 B.n268 585
R211 B.n270 B.n165 585
R212 B.n272 B.n271 585
R213 B.n273 B.n164 585
R214 B.n275 B.n274 585
R215 B.n276 B.n163 585
R216 B.n278 B.n277 585
R217 B.n279 B.n162 585
R218 B.n281 B.n280 585
R219 B.n282 B.n161 585
R220 B.n284 B.n283 585
R221 B.n285 B.n160 585
R222 B.n287 B.n286 585
R223 B.n288 B.n159 585
R224 B.n290 B.n289 585
R225 B.n291 B.n158 585
R226 B.n293 B.n292 585
R227 B.n294 B.n157 585
R228 B.n296 B.n295 585
R229 B.n297 B.n156 585
R230 B.n299 B.n298 585
R231 B.n300 B.n155 585
R232 B.n302 B.n301 585
R233 B.n303 B.n154 585
R234 B.n305 B.n304 585
R235 B.n306 B.n153 585
R236 B.n308 B.n307 585
R237 B.n309 B.n152 585
R238 B.n311 B.n310 585
R239 B.n312 B.n151 585
R240 B.n314 B.n313 585
R241 B.n315 B.n150 585
R242 B.n317 B.n316 585
R243 B.n319 B.n318 585
R244 B.n320 B.n146 585
R245 B.n322 B.n321 585
R246 B.n323 B.n145 585
R247 B.n325 B.n324 585
R248 B.n326 B.n144 585
R249 B.n328 B.n327 585
R250 B.n329 B.n143 585
R251 B.n331 B.n330 585
R252 B.n332 B.n140 585
R253 B.n335 B.n334 585
R254 B.n336 B.n139 585
R255 B.n338 B.n337 585
R256 B.n339 B.n138 585
R257 B.n341 B.n340 585
R258 B.n342 B.n137 585
R259 B.n344 B.n343 585
R260 B.n345 B.n136 585
R261 B.n347 B.n346 585
R262 B.n348 B.n135 585
R263 B.n350 B.n349 585
R264 B.n351 B.n134 585
R265 B.n353 B.n352 585
R266 B.n354 B.n133 585
R267 B.n356 B.n355 585
R268 B.n357 B.n132 585
R269 B.n359 B.n358 585
R270 B.n360 B.n131 585
R271 B.n362 B.n361 585
R272 B.n363 B.n130 585
R273 B.n365 B.n364 585
R274 B.n366 B.n129 585
R275 B.n368 B.n367 585
R276 B.n369 B.n128 585
R277 B.n371 B.n370 585
R278 B.n372 B.n127 585
R279 B.n374 B.n373 585
R280 B.n375 B.n126 585
R281 B.n377 B.n376 585
R282 B.n378 B.n125 585
R283 B.n380 B.n379 585
R284 B.n381 B.n124 585
R285 B.n383 B.n382 585
R286 B.n384 B.n123 585
R287 B.n386 B.n385 585
R288 B.n387 B.n122 585
R289 B.n389 B.n388 585
R290 B.n390 B.n121 585
R291 B.n392 B.n391 585
R292 B.n393 B.n120 585
R293 B.n395 B.n394 585
R294 B.n396 B.n119 585
R295 B.n398 B.n397 585
R296 B.n399 B.n118 585
R297 B.n401 B.n400 585
R298 B.n402 B.n117 585
R299 B.n404 B.n403 585
R300 B.n405 B.n116 585
R301 B.n407 B.n406 585
R302 B.n408 B.n115 585
R303 B.n410 B.n409 585
R304 B.n411 B.n114 585
R305 B.n413 B.n412 585
R306 B.n414 B.n113 585
R307 B.n416 B.n415 585
R308 B.n417 B.n112 585
R309 B.n419 B.n418 585
R310 B.n420 B.n111 585
R311 B.n422 B.n421 585
R312 B.n423 B.n110 585
R313 B.n425 B.n424 585
R314 B.n426 B.n109 585
R315 B.n224 B.n223 585
R316 B.n222 B.n181 585
R317 B.n221 B.n220 585
R318 B.n219 B.n182 585
R319 B.n218 B.n217 585
R320 B.n216 B.n183 585
R321 B.n215 B.n214 585
R322 B.n213 B.n184 585
R323 B.n212 B.n211 585
R324 B.n210 B.n185 585
R325 B.n209 B.n208 585
R326 B.n207 B.n186 585
R327 B.n206 B.n205 585
R328 B.n204 B.n187 585
R329 B.n203 B.n202 585
R330 B.n201 B.n188 585
R331 B.n200 B.n199 585
R332 B.n198 B.n189 585
R333 B.n197 B.n196 585
R334 B.n195 B.n190 585
R335 B.n194 B.n193 585
R336 B.n192 B.n191 585
R337 B.n2 B.n0 585
R338 B.n733 B.n1 585
R339 B.n732 B.n731 585
R340 B.n730 B.n3 585
R341 B.n729 B.n728 585
R342 B.n727 B.n4 585
R343 B.n726 B.n725 585
R344 B.n724 B.n5 585
R345 B.n723 B.n722 585
R346 B.n721 B.n6 585
R347 B.n720 B.n719 585
R348 B.n718 B.n7 585
R349 B.n717 B.n716 585
R350 B.n715 B.n8 585
R351 B.n714 B.n713 585
R352 B.n712 B.n9 585
R353 B.n711 B.n710 585
R354 B.n709 B.n10 585
R355 B.n708 B.n707 585
R356 B.n706 B.n11 585
R357 B.n705 B.n704 585
R358 B.n703 B.n12 585
R359 B.n702 B.n701 585
R360 B.n700 B.n13 585
R361 B.n735 B.n734 585
R362 B.n141 B.t3 543.485
R363 B.n147 B.t9 543.485
R364 B.n46 B.t0 543.485
R365 B.n53 B.t6 543.485
R366 B.n141 B.t5 533.889
R367 B.n53 B.t7 533.889
R368 B.n147 B.t11 533.889
R369 B.n46 B.t1 533.889
R370 B.n142 B.t4 501.307
R371 B.n54 B.t8 501.307
R372 B.n148 B.t10 501.307
R373 B.n47 B.t2 501.307
R374 B.n223 B.n180 473.281
R375 B.n698 B.n13 473.281
R376 B.n427 B.n426 473.281
R377 B.n498 B.n497 473.281
R378 B.n223 B.n222 163.367
R379 B.n222 B.n221 163.367
R380 B.n221 B.n182 163.367
R381 B.n217 B.n182 163.367
R382 B.n217 B.n216 163.367
R383 B.n216 B.n215 163.367
R384 B.n215 B.n184 163.367
R385 B.n211 B.n184 163.367
R386 B.n211 B.n210 163.367
R387 B.n210 B.n209 163.367
R388 B.n209 B.n186 163.367
R389 B.n205 B.n186 163.367
R390 B.n205 B.n204 163.367
R391 B.n204 B.n203 163.367
R392 B.n203 B.n188 163.367
R393 B.n199 B.n188 163.367
R394 B.n199 B.n198 163.367
R395 B.n198 B.n197 163.367
R396 B.n197 B.n190 163.367
R397 B.n193 B.n190 163.367
R398 B.n193 B.n192 163.367
R399 B.n192 B.n2 163.367
R400 B.n734 B.n2 163.367
R401 B.n734 B.n733 163.367
R402 B.n733 B.n732 163.367
R403 B.n732 B.n3 163.367
R404 B.n728 B.n3 163.367
R405 B.n728 B.n727 163.367
R406 B.n727 B.n726 163.367
R407 B.n726 B.n5 163.367
R408 B.n722 B.n5 163.367
R409 B.n722 B.n721 163.367
R410 B.n721 B.n720 163.367
R411 B.n720 B.n7 163.367
R412 B.n716 B.n7 163.367
R413 B.n716 B.n715 163.367
R414 B.n715 B.n714 163.367
R415 B.n714 B.n9 163.367
R416 B.n710 B.n9 163.367
R417 B.n710 B.n709 163.367
R418 B.n709 B.n708 163.367
R419 B.n708 B.n11 163.367
R420 B.n704 B.n11 163.367
R421 B.n704 B.n703 163.367
R422 B.n703 B.n702 163.367
R423 B.n702 B.n13 163.367
R424 B.n227 B.n180 163.367
R425 B.n228 B.n227 163.367
R426 B.n229 B.n228 163.367
R427 B.n229 B.n178 163.367
R428 B.n233 B.n178 163.367
R429 B.n234 B.n233 163.367
R430 B.n235 B.n234 163.367
R431 B.n235 B.n176 163.367
R432 B.n239 B.n176 163.367
R433 B.n240 B.n239 163.367
R434 B.n241 B.n240 163.367
R435 B.n241 B.n174 163.367
R436 B.n245 B.n174 163.367
R437 B.n246 B.n245 163.367
R438 B.n247 B.n246 163.367
R439 B.n247 B.n172 163.367
R440 B.n251 B.n172 163.367
R441 B.n252 B.n251 163.367
R442 B.n253 B.n252 163.367
R443 B.n253 B.n170 163.367
R444 B.n257 B.n170 163.367
R445 B.n258 B.n257 163.367
R446 B.n259 B.n258 163.367
R447 B.n259 B.n168 163.367
R448 B.n263 B.n168 163.367
R449 B.n264 B.n263 163.367
R450 B.n265 B.n264 163.367
R451 B.n265 B.n166 163.367
R452 B.n269 B.n166 163.367
R453 B.n270 B.n269 163.367
R454 B.n271 B.n270 163.367
R455 B.n271 B.n164 163.367
R456 B.n275 B.n164 163.367
R457 B.n276 B.n275 163.367
R458 B.n277 B.n276 163.367
R459 B.n277 B.n162 163.367
R460 B.n281 B.n162 163.367
R461 B.n282 B.n281 163.367
R462 B.n283 B.n282 163.367
R463 B.n283 B.n160 163.367
R464 B.n287 B.n160 163.367
R465 B.n288 B.n287 163.367
R466 B.n289 B.n288 163.367
R467 B.n289 B.n158 163.367
R468 B.n293 B.n158 163.367
R469 B.n294 B.n293 163.367
R470 B.n295 B.n294 163.367
R471 B.n295 B.n156 163.367
R472 B.n299 B.n156 163.367
R473 B.n300 B.n299 163.367
R474 B.n301 B.n300 163.367
R475 B.n301 B.n154 163.367
R476 B.n305 B.n154 163.367
R477 B.n306 B.n305 163.367
R478 B.n307 B.n306 163.367
R479 B.n307 B.n152 163.367
R480 B.n311 B.n152 163.367
R481 B.n312 B.n311 163.367
R482 B.n313 B.n312 163.367
R483 B.n313 B.n150 163.367
R484 B.n317 B.n150 163.367
R485 B.n318 B.n317 163.367
R486 B.n318 B.n146 163.367
R487 B.n322 B.n146 163.367
R488 B.n323 B.n322 163.367
R489 B.n324 B.n323 163.367
R490 B.n324 B.n144 163.367
R491 B.n328 B.n144 163.367
R492 B.n329 B.n328 163.367
R493 B.n330 B.n329 163.367
R494 B.n330 B.n140 163.367
R495 B.n335 B.n140 163.367
R496 B.n336 B.n335 163.367
R497 B.n337 B.n336 163.367
R498 B.n337 B.n138 163.367
R499 B.n341 B.n138 163.367
R500 B.n342 B.n341 163.367
R501 B.n343 B.n342 163.367
R502 B.n343 B.n136 163.367
R503 B.n347 B.n136 163.367
R504 B.n348 B.n347 163.367
R505 B.n349 B.n348 163.367
R506 B.n349 B.n134 163.367
R507 B.n353 B.n134 163.367
R508 B.n354 B.n353 163.367
R509 B.n355 B.n354 163.367
R510 B.n355 B.n132 163.367
R511 B.n359 B.n132 163.367
R512 B.n360 B.n359 163.367
R513 B.n361 B.n360 163.367
R514 B.n361 B.n130 163.367
R515 B.n365 B.n130 163.367
R516 B.n366 B.n365 163.367
R517 B.n367 B.n366 163.367
R518 B.n367 B.n128 163.367
R519 B.n371 B.n128 163.367
R520 B.n372 B.n371 163.367
R521 B.n373 B.n372 163.367
R522 B.n373 B.n126 163.367
R523 B.n377 B.n126 163.367
R524 B.n378 B.n377 163.367
R525 B.n379 B.n378 163.367
R526 B.n379 B.n124 163.367
R527 B.n383 B.n124 163.367
R528 B.n384 B.n383 163.367
R529 B.n385 B.n384 163.367
R530 B.n385 B.n122 163.367
R531 B.n389 B.n122 163.367
R532 B.n390 B.n389 163.367
R533 B.n391 B.n390 163.367
R534 B.n391 B.n120 163.367
R535 B.n395 B.n120 163.367
R536 B.n396 B.n395 163.367
R537 B.n397 B.n396 163.367
R538 B.n397 B.n118 163.367
R539 B.n401 B.n118 163.367
R540 B.n402 B.n401 163.367
R541 B.n403 B.n402 163.367
R542 B.n403 B.n116 163.367
R543 B.n407 B.n116 163.367
R544 B.n408 B.n407 163.367
R545 B.n409 B.n408 163.367
R546 B.n409 B.n114 163.367
R547 B.n413 B.n114 163.367
R548 B.n414 B.n413 163.367
R549 B.n415 B.n414 163.367
R550 B.n415 B.n112 163.367
R551 B.n419 B.n112 163.367
R552 B.n420 B.n419 163.367
R553 B.n421 B.n420 163.367
R554 B.n421 B.n110 163.367
R555 B.n425 B.n110 163.367
R556 B.n426 B.n425 163.367
R557 B.n427 B.n108 163.367
R558 B.n431 B.n108 163.367
R559 B.n432 B.n431 163.367
R560 B.n433 B.n432 163.367
R561 B.n433 B.n106 163.367
R562 B.n437 B.n106 163.367
R563 B.n438 B.n437 163.367
R564 B.n439 B.n438 163.367
R565 B.n439 B.n104 163.367
R566 B.n443 B.n104 163.367
R567 B.n444 B.n443 163.367
R568 B.n445 B.n444 163.367
R569 B.n445 B.n102 163.367
R570 B.n449 B.n102 163.367
R571 B.n450 B.n449 163.367
R572 B.n451 B.n450 163.367
R573 B.n451 B.n100 163.367
R574 B.n455 B.n100 163.367
R575 B.n456 B.n455 163.367
R576 B.n457 B.n456 163.367
R577 B.n457 B.n98 163.367
R578 B.n461 B.n98 163.367
R579 B.n462 B.n461 163.367
R580 B.n463 B.n462 163.367
R581 B.n463 B.n96 163.367
R582 B.n467 B.n96 163.367
R583 B.n468 B.n467 163.367
R584 B.n469 B.n468 163.367
R585 B.n469 B.n94 163.367
R586 B.n473 B.n94 163.367
R587 B.n474 B.n473 163.367
R588 B.n475 B.n474 163.367
R589 B.n475 B.n92 163.367
R590 B.n479 B.n92 163.367
R591 B.n480 B.n479 163.367
R592 B.n481 B.n480 163.367
R593 B.n481 B.n90 163.367
R594 B.n485 B.n90 163.367
R595 B.n486 B.n485 163.367
R596 B.n487 B.n486 163.367
R597 B.n487 B.n88 163.367
R598 B.n491 B.n88 163.367
R599 B.n492 B.n491 163.367
R600 B.n493 B.n492 163.367
R601 B.n493 B.n86 163.367
R602 B.n497 B.n86 163.367
R603 B.n698 B.n697 163.367
R604 B.n697 B.n696 163.367
R605 B.n696 B.n15 163.367
R606 B.n692 B.n15 163.367
R607 B.n692 B.n691 163.367
R608 B.n691 B.n690 163.367
R609 B.n690 B.n17 163.367
R610 B.n686 B.n17 163.367
R611 B.n686 B.n685 163.367
R612 B.n685 B.n684 163.367
R613 B.n684 B.n19 163.367
R614 B.n680 B.n19 163.367
R615 B.n680 B.n679 163.367
R616 B.n679 B.n678 163.367
R617 B.n678 B.n21 163.367
R618 B.n674 B.n21 163.367
R619 B.n674 B.n673 163.367
R620 B.n673 B.n672 163.367
R621 B.n672 B.n23 163.367
R622 B.n668 B.n23 163.367
R623 B.n668 B.n667 163.367
R624 B.n667 B.n666 163.367
R625 B.n666 B.n25 163.367
R626 B.n662 B.n25 163.367
R627 B.n662 B.n661 163.367
R628 B.n661 B.n660 163.367
R629 B.n660 B.n27 163.367
R630 B.n656 B.n27 163.367
R631 B.n656 B.n655 163.367
R632 B.n655 B.n654 163.367
R633 B.n654 B.n29 163.367
R634 B.n650 B.n29 163.367
R635 B.n650 B.n649 163.367
R636 B.n649 B.n648 163.367
R637 B.n648 B.n31 163.367
R638 B.n644 B.n31 163.367
R639 B.n644 B.n643 163.367
R640 B.n643 B.n642 163.367
R641 B.n642 B.n33 163.367
R642 B.n638 B.n33 163.367
R643 B.n638 B.n637 163.367
R644 B.n637 B.n636 163.367
R645 B.n636 B.n35 163.367
R646 B.n632 B.n35 163.367
R647 B.n632 B.n631 163.367
R648 B.n631 B.n630 163.367
R649 B.n630 B.n37 163.367
R650 B.n626 B.n37 163.367
R651 B.n626 B.n625 163.367
R652 B.n625 B.n624 163.367
R653 B.n624 B.n39 163.367
R654 B.n620 B.n39 163.367
R655 B.n620 B.n619 163.367
R656 B.n619 B.n618 163.367
R657 B.n618 B.n41 163.367
R658 B.n614 B.n41 163.367
R659 B.n614 B.n613 163.367
R660 B.n613 B.n612 163.367
R661 B.n612 B.n43 163.367
R662 B.n608 B.n43 163.367
R663 B.n608 B.n607 163.367
R664 B.n607 B.n606 163.367
R665 B.n606 B.n45 163.367
R666 B.n602 B.n45 163.367
R667 B.n602 B.n601 163.367
R668 B.n601 B.n600 163.367
R669 B.n600 B.n50 163.367
R670 B.n596 B.n50 163.367
R671 B.n596 B.n595 163.367
R672 B.n595 B.n594 163.367
R673 B.n594 B.n52 163.367
R674 B.n589 B.n52 163.367
R675 B.n589 B.n588 163.367
R676 B.n588 B.n587 163.367
R677 B.n587 B.n56 163.367
R678 B.n583 B.n56 163.367
R679 B.n583 B.n582 163.367
R680 B.n582 B.n581 163.367
R681 B.n581 B.n58 163.367
R682 B.n577 B.n58 163.367
R683 B.n577 B.n576 163.367
R684 B.n576 B.n575 163.367
R685 B.n575 B.n60 163.367
R686 B.n571 B.n60 163.367
R687 B.n571 B.n570 163.367
R688 B.n570 B.n569 163.367
R689 B.n569 B.n62 163.367
R690 B.n565 B.n62 163.367
R691 B.n565 B.n564 163.367
R692 B.n564 B.n563 163.367
R693 B.n563 B.n64 163.367
R694 B.n559 B.n64 163.367
R695 B.n559 B.n558 163.367
R696 B.n558 B.n557 163.367
R697 B.n557 B.n66 163.367
R698 B.n553 B.n66 163.367
R699 B.n553 B.n552 163.367
R700 B.n552 B.n551 163.367
R701 B.n551 B.n68 163.367
R702 B.n547 B.n68 163.367
R703 B.n547 B.n546 163.367
R704 B.n546 B.n545 163.367
R705 B.n545 B.n70 163.367
R706 B.n541 B.n70 163.367
R707 B.n541 B.n540 163.367
R708 B.n540 B.n539 163.367
R709 B.n539 B.n72 163.367
R710 B.n535 B.n72 163.367
R711 B.n535 B.n534 163.367
R712 B.n534 B.n533 163.367
R713 B.n533 B.n74 163.367
R714 B.n529 B.n74 163.367
R715 B.n529 B.n528 163.367
R716 B.n528 B.n527 163.367
R717 B.n527 B.n76 163.367
R718 B.n523 B.n76 163.367
R719 B.n523 B.n522 163.367
R720 B.n522 B.n521 163.367
R721 B.n521 B.n78 163.367
R722 B.n517 B.n78 163.367
R723 B.n517 B.n516 163.367
R724 B.n516 B.n515 163.367
R725 B.n515 B.n80 163.367
R726 B.n511 B.n80 163.367
R727 B.n511 B.n510 163.367
R728 B.n510 B.n509 163.367
R729 B.n509 B.n82 163.367
R730 B.n505 B.n82 163.367
R731 B.n505 B.n504 163.367
R732 B.n504 B.n503 163.367
R733 B.n503 B.n84 163.367
R734 B.n499 B.n84 163.367
R735 B.n499 B.n498 163.367
R736 B.n333 B.n142 59.5399
R737 B.n149 B.n148 59.5399
R738 B.n48 B.n47 59.5399
R739 B.n591 B.n54 59.5399
R740 B.n142 B.n141 32.5823
R741 B.n148 B.n147 32.5823
R742 B.n47 B.n46 32.5823
R743 B.n54 B.n53 32.5823
R744 B.n700 B.n699 30.7517
R745 B.n496 B.n85 30.7517
R746 B.n428 B.n109 30.7517
R747 B.n225 B.n224 30.7517
R748 B B.n735 18.0485
R749 B.n699 B.n14 10.6151
R750 B.n695 B.n14 10.6151
R751 B.n695 B.n694 10.6151
R752 B.n694 B.n693 10.6151
R753 B.n693 B.n16 10.6151
R754 B.n689 B.n16 10.6151
R755 B.n689 B.n688 10.6151
R756 B.n688 B.n687 10.6151
R757 B.n687 B.n18 10.6151
R758 B.n683 B.n18 10.6151
R759 B.n683 B.n682 10.6151
R760 B.n682 B.n681 10.6151
R761 B.n681 B.n20 10.6151
R762 B.n677 B.n20 10.6151
R763 B.n677 B.n676 10.6151
R764 B.n676 B.n675 10.6151
R765 B.n675 B.n22 10.6151
R766 B.n671 B.n22 10.6151
R767 B.n671 B.n670 10.6151
R768 B.n670 B.n669 10.6151
R769 B.n669 B.n24 10.6151
R770 B.n665 B.n24 10.6151
R771 B.n665 B.n664 10.6151
R772 B.n664 B.n663 10.6151
R773 B.n663 B.n26 10.6151
R774 B.n659 B.n26 10.6151
R775 B.n659 B.n658 10.6151
R776 B.n658 B.n657 10.6151
R777 B.n657 B.n28 10.6151
R778 B.n653 B.n28 10.6151
R779 B.n653 B.n652 10.6151
R780 B.n652 B.n651 10.6151
R781 B.n651 B.n30 10.6151
R782 B.n647 B.n30 10.6151
R783 B.n647 B.n646 10.6151
R784 B.n646 B.n645 10.6151
R785 B.n645 B.n32 10.6151
R786 B.n641 B.n32 10.6151
R787 B.n641 B.n640 10.6151
R788 B.n640 B.n639 10.6151
R789 B.n639 B.n34 10.6151
R790 B.n635 B.n34 10.6151
R791 B.n635 B.n634 10.6151
R792 B.n634 B.n633 10.6151
R793 B.n633 B.n36 10.6151
R794 B.n629 B.n36 10.6151
R795 B.n629 B.n628 10.6151
R796 B.n628 B.n627 10.6151
R797 B.n627 B.n38 10.6151
R798 B.n623 B.n38 10.6151
R799 B.n623 B.n622 10.6151
R800 B.n622 B.n621 10.6151
R801 B.n621 B.n40 10.6151
R802 B.n617 B.n40 10.6151
R803 B.n617 B.n616 10.6151
R804 B.n616 B.n615 10.6151
R805 B.n615 B.n42 10.6151
R806 B.n611 B.n42 10.6151
R807 B.n611 B.n610 10.6151
R808 B.n610 B.n609 10.6151
R809 B.n609 B.n44 10.6151
R810 B.n605 B.n604 10.6151
R811 B.n604 B.n603 10.6151
R812 B.n603 B.n49 10.6151
R813 B.n599 B.n49 10.6151
R814 B.n599 B.n598 10.6151
R815 B.n598 B.n597 10.6151
R816 B.n597 B.n51 10.6151
R817 B.n593 B.n51 10.6151
R818 B.n593 B.n592 10.6151
R819 B.n590 B.n55 10.6151
R820 B.n586 B.n55 10.6151
R821 B.n586 B.n585 10.6151
R822 B.n585 B.n584 10.6151
R823 B.n584 B.n57 10.6151
R824 B.n580 B.n57 10.6151
R825 B.n580 B.n579 10.6151
R826 B.n579 B.n578 10.6151
R827 B.n578 B.n59 10.6151
R828 B.n574 B.n59 10.6151
R829 B.n574 B.n573 10.6151
R830 B.n573 B.n572 10.6151
R831 B.n572 B.n61 10.6151
R832 B.n568 B.n61 10.6151
R833 B.n568 B.n567 10.6151
R834 B.n567 B.n566 10.6151
R835 B.n566 B.n63 10.6151
R836 B.n562 B.n63 10.6151
R837 B.n562 B.n561 10.6151
R838 B.n561 B.n560 10.6151
R839 B.n560 B.n65 10.6151
R840 B.n556 B.n65 10.6151
R841 B.n556 B.n555 10.6151
R842 B.n555 B.n554 10.6151
R843 B.n554 B.n67 10.6151
R844 B.n550 B.n67 10.6151
R845 B.n550 B.n549 10.6151
R846 B.n549 B.n548 10.6151
R847 B.n548 B.n69 10.6151
R848 B.n544 B.n69 10.6151
R849 B.n544 B.n543 10.6151
R850 B.n543 B.n542 10.6151
R851 B.n542 B.n71 10.6151
R852 B.n538 B.n71 10.6151
R853 B.n538 B.n537 10.6151
R854 B.n537 B.n536 10.6151
R855 B.n536 B.n73 10.6151
R856 B.n532 B.n73 10.6151
R857 B.n532 B.n531 10.6151
R858 B.n531 B.n530 10.6151
R859 B.n530 B.n75 10.6151
R860 B.n526 B.n75 10.6151
R861 B.n526 B.n525 10.6151
R862 B.n525 B.n524 10.6151
R863 B.n524 B.n77 10.6151
R864 B.n520 B.n77 10.6151
R865 B.n520 B.n519 10.6151
R866 B.n519 B.n518 10.6151
R867 B.n518 B.n79 10.6151
R868 B.n514 B.n79 10.6151
R869 B.n514 B.n513 10.6151
R870 B.n513 B.n512 10.6151
R871 B.n512 B.n81 10.6151
R872 B.n508 B.n81 10.6151
R873 B.n508 B.n507 10.6151
R874 B.n507 B.n506 10.6151
R875 B.n506 B.n83 10.6151
R876 B.n502 B.n83 10.6151
R877 B.n502 B.n501 10.6151
R878 B.n501 B.n500 10.6151
R879 B.n500 B.n85 10.6151
R880 B.n429 B.n428 10.6151
R881 B.n430 B.n429 10.6151
R882 B.n430 B.n107 10.6151
R883 B.n434 B.n107 10.6151
R884 B.n435 B.n434 10.6151
R885 B.n436 B.n435 10.6151
R886 B.n436 B.n105 10.6151
R887 B.n440 B.n105 10.6151
R888 B.n441 B.n440 10.6151
R889 B.n442 B.n441 10.6151
R890 B.n442 B.n103 10.6151
R891 B.n446 B.n103 10.6151
R892 B.n447 B.n446 10.6151
R893 B.n448 B.n447 10.6151
R894 B.n448 B.n101 10.6151
R895 B.n452 B.n101 10.6151
R896 B.n453 B.n452 10.6151
R897 B.n454 B.n453 10.6151
R898 B.n454 B.n99 10.6151
R899 B.n458 B.n99 10.6151
R900 B.n459 B.n458 10.6151
R901 B.n460 B.n459 10.6151
R902 B.n460 B.n97 10.6151
R903 B.n464 B.n97 10.6151
R904 B.n465 B.n464 10.6151
R905 B.n466 B.n465 10.6151
R906 B.n466 B.n95 10.6151
R907 B.n470 B.n95 10.6151
R908 B.n471 B.n470 10.6151
R909 B.n472 B.n471 10.6151
R910 B.n472 B.n93 10.6151
R911 B.n476 B.n93 10.6151
R912 B.n477 B.n476 10.6151
R913 B.n478 B.n477 10.6151
R914 B.n478 B.n91 10.6151
R915 B.n482 B.n91 10.6151
R916 B.n483 B.n482 10.6151
R917 B.n484 B.n483 10.6151
R918 B.n484 B.n89 10.6151
R919 B.n488 B.n89 10.6151
R920 B.n489 B.n488 10.6151
R921 B.n490 B.n489 10.6151
R922 B.n490 B.n87 10.6151
R923 B.n494 B.n87 10.6151
R924 B.n495 B.n494 10.6151
R925 B.n496 B.n495 10.6151
R926 B.n226 B.n225 10.6151
R927 B.n226 B.n179 10.6151
R928 B.n230 B.n179 10.6151
R929 B.n231 B.n230 10.6151
R930 B.n232 B.n231 10.6151
R931 B.n232 B.n177 10.6151
R932 B.n236 B.n177 10.6151
R933 B.n237 B.n236 10.6151
R934 B.n238 B.n237 10.6151
R935 B.n238 B.n175 10.6151
R936 B.n242 B.n175 10.6151
R937 B.n243 B.n242 10.6151
R938 B.n244 B.n243 10.6151
R939 B.n244 B.n173 10.6151
R940 B.n248 B.n173 10.6151
R941 B.n249 B.n248 10.6151
R942 B.n250 B.n249 10.6151
R943 B.n250 B.n171 10.6151
R944 B.n254 B.n171 10.6151
R945 B.n255 B.n254 10.6151
R946 B.n256 B.n255 10.6151
R947 B.n256 B.n169 10.6151
R948 B.n260 B.n169 10.6151
R949 B.n261 B.n260 10.6151
R950 B.n262 B.n261 10.6151
R951 B.n262 B.n167 10.6151
R952 B.n266 B.n167 10.6151
R953 B.n267 B.n266 10.6151
R954 B.n268 B.n267 10.6151
R955 B.n268 B.n165 10.6151
R956 B.n272 B.n165 10.6151
R957 B.n273 B.n272 10.6151
R958 B.n274 B.n273 10.6151
R959 B.n274 B.n163 10.6151
R960 B.n278 B.n163 10.6151
R961 B.n279 B.n278 10.6151
R962 B.n280 B.n279 10.6151
R963 B.n280 B.n161 10.6151
R964 B.n284 B.n161 10.6151
R965 B.n285 B.n284 10.6151
R966 B.n286 B.n285 10.6151
R967 B.n286 B.n159 10.6151
R968 B.n290 B.n159 10.6151
R969 B.n291 B.n290 10.6151
R970 B.n292 B.n291 10.6151
R971 B.n292 B.n157 10.6151
R972 B.n296 B.n157 10.6151
R973 B.n297 B.n296 10.6151
R974 B.n298 B.n297 10.6151
R975 B.n298 B.n155 10.6151
R976 B.n302 B.n155 10.6151
R977 B.n303 B.n302 10.6151
R978 B.n304 B.n303 10.6151
R979 B.n304 B.n153 10.6151
R980 B.n308 B.n153 10.6151
R981 B.n309 B.n308 10.6151
R982 B.n310 B.n309 10.6151
R983 B.n310 B.n151 10.6151
R984 B.n314 B.n151 10.6151
R985 B.n315 B.n314 10.6151
R986 B.n316 B.n315 10.6151
R987 B.n320 B.n319 10.6151
R988 B.n321 B.n320 10.6151
R989 B.n321 B.n145 10.6151
R990 B.n325 B.n145 10.6151
R991 B.n326 B.n325 10.6151
R992 B.n327 B.n326 10.6151
R993 B.n327 B.n143 10.6151
R994 B.n331 B.n143 10.6151
R995 B.n332 B.n331 10.6151
R996 B.n334 B.n139 10.6151
R997 B.n338 B.n139 10.6151
R998 B.n339 B.n338 10.6151
R999 B.n340 B.n339 10.6151
R1000 B.n340 B.n137 10.6151
R1001 B.n344 B.n137 10.6151
R1002 B.n345 B.n344 10.6151
R1003 B.n346 B.n345 10.6151
R1004 B.n346 B.n135 10.6151
R1005 B.n350 B.n135 10.6151
R1006 B.n351 B.n350 10.6151
R1007 B.n352 B.n351 10.6151
R1008 B.n352 B.n133 10.6151
R1009 B.n356 B.n133 10.6151
R1010 B.n357 B.n356 10.6151
R1011 B.n358 B.n357 10.6151
R1012 B.n358 B.n131 10.6151
R1013 B.n362 B.n131 10.6151
R1014 B.n363 B.n362 10.6151
R1015 B.n364 B.n363 10.6151
R1016 B.n364 B.n129 10.6151
R1017 B.n368 B.n129 10.6151
R1018 B.n369 B.n368 10.6151
R1019 B.n370 B.n369 10.6151
R1020 B.n370 B.n127 10.6151
R1021 B.n374 B.n127 10.6151
R1022 B.n375 B.n374 10.6151
R1023 B.n376 B.n375 10.6151
R1024 B.n376 B.n125 10.6151
R1025 B.n380 B.n125 10.6151
R1026 B.n381 B.n380 10.6151
R1027 B.n382 B.n381 10.6151
R1028 B.n382 B.n123 10.6151
R1029 B.n386 B.n123 10.6151
R1030 B.n387 B.n386 10.6151
R1031 B.n388 B.n387 10.6151
R1032 B.n388 B.n121 10.6151
R1033 B.n392 B.n121 10.6151
R1034 B.n393 B.n392 10.6151
R1035 B.n394 B.n393 10.6151
R1036 B.n394 B.n119 10.6151
R1037 B.n398 B.n119 10.6151
R1038 B.n399 B.n398 10.6151
R1039 B.n400 B.n399 10.6151
R1040 B.n400 B.n117 10.6151
R1041 B.n404 B.n117 10.6151
R1042 B.n405 B.n404 10.6151
R1043 B.n406 B.n405 10.6151
R1044 B.n406 B.n115 10.6151
R1045 B.n410 B.n115 10.6151
R1046 B.n411 B.n410 10.6151
R1047 B.n412 B.n411 10.6151
R1048 B.n412 B.n113 10.6151
R1049 B.n416 B.n113 10.6151
R1050 B.n417 B.n416 10.6151
R1051 B.n418 B.n417 10.6151
R1052 B.n418 B.n111 10.6151
R1053 B.n422 B.n111 10.6151
R1054 B.n423 B.n422 10.6151
R1055 B.n424 B.n423 10.6151
R1056 B.n424 B.n109 10.6151
R1057 B.n224 B.n181 10.6151
R1058 B.n220 B.n181 10.6151
R1059 B.n220 B.n219 10.6151
R1060 B.n219 B.n218 10.6151
R1061 B.n218 B.n183 10.6151
R1062 B.n214 B.n183 10.6151
R1063 B.n214 B.n213 10.6151
R1064 B.n213 B.n212 10.6151
R1065 B.n212 B.n185 10.6151
R1066 B.n208 B.n185 10.6151
R1067 B.n208 B.n207 10.6151
R1068 B.n207 B.n206 10.6151
R1069 B.n206 B.n187 10.6151
R1070 B.n202 B.n187 10.6151
R1071 B.n202 B.n201 10.6151
R1072 B.n201 B.n200 10.6151
R1073 B.n200 B.n189 10.6151
R1074 B.n196 B.n189 10.6151
R1075 B.n196 B.n195 10.6151
R1076 B.n195 B.n194 10.6151
R1077 B.n194 B.n191 10.6151
R1078 B.n191 B.n0 10.6151
R1079 B.n731 B.n1 10.6151
R1080 B.n731 B.n730 10.6151
R1081 B.n730 B.n729 10.6151
R1082 B.n729 B.n4 10.6151
R1083 B.n725 B.n4 10.6151
R1084 B.n725 B.n724 10.6151
R1085 B.n724 B.n723 10.6151
R1086 B.n723 B.n6 10.6151
R1087 B.n719 B.n6 10.6151
R1088 B.n719 B.n718 10.6151
R1089 B.n718 B.n717 10.6151
R1090 B.n717 B.n8 10.6151
R1091 B.n713 B.n8 10.6151
R1092 B.n713 B.n712 10.6151
R1093 B.n712 B.n711 10.6151
R1094 B.n711 B.n10 10.6151
R1095 B.n707 B.n10 10.6151
R1096 B.n707 B.n706 10.6151
R1097 B.n706 B.n705 10.6151
R1098 B.n705 B.n12 10.6151
R1099 B.n701 B.n12 10.6151
R1100 B.n701 B.n700 10.6151
R1101 B.n48 B.n44 9.36635
R1102 B.n591 B.n590 9.36635
R1103 B.n316 B.n149 9.36635
R1104 B.n334 B.n333 9.36635
R1105 B.n735 B.n0 2.81026
R1106 B.n735 B.n1 2.81026
R1107 B.n605 B.n48 1.24928
R1108 B.n592 B.n591 1.24928
R1109 B.n319 B.n149 1.24928
R1110 B.n333 B.n332 1.24928
R1111 VN.n0 VN.t0 376.8
R1112 VN.n1 VN.t2 376.8
R1113 VN.n0 VN.t1 376.57
R1114 VN.n1 VN.t3 376.57
R1115 VN VN.n1 65.8428
R1116 VN VN.n0 17.7405
R1117 VDD2.n2 VDD2.n0 112.992
R1118 VDD2.n2 VDD2.n1 68.5787
R1119 VDD2.n1 VDD2.t1 1.714
R1120 VDD2.n1 VDD2.t0 1.714
R1121 VDD2.n0 VDD2.t3 1.714
R1122 VDD2.n0 VDD2.t2 1.714
R1123 VDD2 VDD2.n2 0.0586897
R1124 VTAIL.n842 VTAIL.n742 756.745
R1125 VTAIL.n100 VTAIL.n0 756.745
R1126 VTAIL.n206 VTAIL.n106 756.745
R1127 VTAIL.n312 VTAIL.n212 756.745
R1128 VTAIL.n736 VTAIL.n636 756.745
R1129 VTAIL.n630 VTAIL.n530 756.745
R1130 VTAIL.n524 VTAIL.n424 756.745
R1131 VTAIL.n418 VTAIL.n318 756.745
R1132 VTAIL.n777 VTAIL.n776 585
R1133 VTAIL.n774 VTAIL.n773 585
R1134 VTAIL.n783 VTAIL.n782 585
R1135 VTAIL.n785 VTAIL.n784 585
R1136 VTAIL.n770 VTAIL.n769 585
R1137 VTAIL.n791 VTAIL.n790 585
R1138 VTAIL.n793 VTAIL.n792 585
R1139 VTAIL.n766 VTAIL.n765 585
R1140 VTAIL.n799 VTAIL.n798 585
R1141 VTAIL.n801 VTAIL.n800 585
R1142 VTAIL.n762 VTAIL.n761 585
R1143 VTAIL.n807 VTAIL.n806 585
R1144 VTAIL.n809 VTAIL.n808 585
R1145 VTAIL.n758 VTAIL.n757 585
R1146 VTAIL.n815 VTAIL.n814 585
R1147 VTAIL.n818 VTAIL.n817 585
R1148 VTAIL.n816 VTAIL.n754 585
R1149 VTAIL.n823 VTAIL.n753 585
R1150 VTAIL.n825 VTAIL.n824 585
R1151 VTAIL.n827 VTAIL.n826 585
R1152 VTAIL.n750 VTAIL.n749 585
R1153 VTAIL.n833 VTAIL.n832 585
R1154 VTAIL.n835 VTAIL.n834 585
R1155 VTAIL.n746 VTAIL.n745 585
R1156 VTAIL.n841 VTAIL.n840 585
R1157 VTAIL.n843 VTAIL.n842 585
R1158 VTAIL.n35 VTAIL.n34 585
R1159 VTAIL.n32 VTAIL.n31 585
R1160 VTAIL.n41 VTAIL.n40 585
R1161 VTAIL.n43 VTAIL.n42 585
R1162 VTAIL.n28 VTAIL.n27 585
R1163 VTAIL.n49 VTAIL.n48 585
R1164 VTAIL.n51 VTAIL.n50 585
R1165 VTAIL.n24 VTAIL.n23 585
R1166 VTAIL.n57 VTAIL.n56 585
R1167 VTAIL.n59 VTAIL.n58 585
R1168 VTAIL.n20 VTAIL.n19 585
R1169 VTAIL.n65 VTAIL.n64 585
R1170 VTAIL.n67 VTAIL.n66 585
R1171 VTAIL.n16 VTAIL.n15 585
R1172 VTAIL.n73 VTAIL.n72 585
R1173 VTAIL.n76 VTAIL.n75 585
R1174 VTAIL.n74 VTAIL.n12 585
R1175 VTAIL.n81 VTAIL.n11 585
R1176 VTAIL.n83 VTAIL.n82 585
R1177 VTAIL.n85 VTAIL.n84 585
R1178 VTAIL.n8 VTAIL.n7 585
R1179 VTAIL.n91 VTAIL.n90 585
R1180 VTAIL.n93 VTAIL.n92 585
R1181 VTAIL.n4 VTAIL.n3 585
R1182 VTAIL.n99 VTAIL.n98 585
R1183 VTAIL.n101 VTAIL.n100 585
R1184 VTAIL.n141 VTAIL.n140 585
R1185 VTAIL.n138 VTAIL.n137 585
R1186 VTAIL.n147 VTAIL.n146 585
R1187 VTAIL.n149 VTAIL.n148 585
R1188 VTAIL.n134 VTAIL.n133 585
R1189 VTAIL.n155 VTAIL.n154 585
R1190 VTAIL.n157 VTAIL.n156 585
R1191 VTAIL.n130 VTAIL.n129 585
R1192 VTAIL.n163 VTAIL.n162 585
R1193 VTAIL.n165 VTAIL.n164 585
R1194 VTAIL.n126 VTAIL.n125 585
R1195 VTAIL.n171 VTAIL.n170 585
R1196 VTAIL.n173 VTAIL.n172 585
R1197 VTAIL.n122 VTAIL.n121 585
R1198 VTAIL.n179 VTAIL.n178 585
R1199 VTAIL.n182 VTAIL.n181 585
R1200 VTAIL.n180 VTAIL.n118 585
R1201 VTAIL.n187 VTAIL.n117 585
R1202 VTAIL.n189 VTAIL.n188 585
R1203 VTAIL.n191 VTAIL.n190 585
R1204 VTAIL.n114 VTAIL.n113 585
R1205 VTAIL.n197 VTAIL.n196 585
R1206 VTAIL.n199 VTAIL.n198 585
R1207 VTAIL.n110 VTAIL.n109 585
R1208 VTAIL.n205 VTAIL.n204 585
R1209 VTAIL.n207 VTAIL.n206 585
R1210 VTAIL.n247 VTAIL.n246 585
R1211 VTAIL.n244 VTAIL.n243 585
R1212 VTAIL.n253 VTAIL.n252 585
R1213 VTAIL.n255 VTAIL.n254 585
R1214 VTAIL.n240 VTAIL.n239 585
R1215 VTAIL.n261 VTAIL.n260 585
R1216 VTAIL.n263 VTAIL.n262 585
R1217 VTAIL.n236 VTAIL.n235 585
R1218 VTAIL.n269 VTAIL.n268 585
R1219 VTAIL.n271 VTAIL.n270 585
R1220 VTAIL.n232 VTAIL.n231 585
R1221 VTAIL.n277 VTAIL.n276 585
R1222 VTAIL.n279 VTAIL.n278 585
R1223 VTAIL.n228 VTAIL.n227 585
R1224 VTAIL.n285 VTAIL.n284 585
R1225 VTAIL.n288 VTAIL.n287 585
R1226 VTAIL.n286 VTAIL.n224 585
R1227 VTAIL.n293 VTAIL.n223 585
R1228 VTAIL.n295 VTAIL.n294 585
R1229 VTAIL.n297 VTAIL.n296 585
R1230 VTAIL.n220 VTAIL.n219 585
R1231 VTAIL.n303 VTAIL.n302 585
R1232 VTAIL.n305 VTAIL.n304 585
R1233 VTAIL.n216 VTAIL.n215 585
R1234 VTAIL.n311 VTAIL.n310 585
R1235 VTAIL.n313 VTAIL.n312 585
R1236 VTAIL.n737 VTAIL.n736 585
R1237 VTAIL.n735 VTAIL.n734 585
R1238 VTAIL.n640 VTAIL.n639 585
R1239 VTAIL.n729 VTAIL.n728 585
R1240 VTAIL.n727 VTAIL.n726 585
R1241 VTAIL.n644 VTAIL.n643 585
R1242 VTAIL.n721 VTAIL.n720 585
R1243 VTAIL.n719 VTAIL.n718 585
R1244 VTAIL.n717 VTAIL.n647 585
R1245 VTAIL.n651 VTAIL.n648 585
R1246 VTAIL.n712 VTAIL.n711 585
R1247 VTAIL.n710 VTAIL.n709 585
R1248 VTAIL.n653 VTAIL.n652 585
R1249 VTAIL.n704 VTAIL.n703 585
R1250 VTAIL.n702 VTAIL.n701 585
R1251 VTAIL.n657 VTAIL.n656 585
R1252 VTAIL.n696 VTAIL.n695 585
R1253 VTAIL.n694 VTAIL.n693 585
R1254 VTAIL.n661 VTAIL.n660 585
R1255 VTAIL.n688 VTAIL.n687 585
R1256 VTAIL.n686 VTAIL.n685 585
R1257 VTAIL.n665 VTAIL.n664 585
R1258 VTAIL.n680 VTAIL.n679 585
R1259 VTAIL.n678 VTAIL.n677 585
R1260 VTAIL.n669 VTAIL.n668 585
R1261 VTAIL.n672 VTAIL.n671 585
R1262 VTAIL.n631 VTAIL.n630 585
R1263 VTAIL.n629 VTAIL.n628 585
R1264 VTAIL.n534 VTAIL.n533 585
R1265 VTAIL.n623 VTAIL.n622 585
R1266 VTAIL.n621 VTAIL.n620 585
R1267 VTAIL.n538 VTAIL.n537 585
R1268 VTAIL.n615 VTAIL.n614 585
R1269 VTAIL.n613 VTAIL.n612 585
R1270 VTAIL.n611 VTAIL.n541 585
R1271 VTAIL.n545 VTAIL.n542 585
R1272 VTAIL.n606 VTAIL.n605 585
R1273 VTAIL.n604 VTAIL.n603 585
R1274 VTAIL.n547 VTAIL.n546 585
R1275 VTAIL.n598 VTAIL.n597 585
R1276 VTAIL.n596 VTAIL.n595 585
R1277 VTAIL.n551 VTAIL.n550 585
R1278 VTAIL.n590 VTAIL.n589 585
R1279 VTAIL.n588 VTAIL.n587 585
R1280 VTAIL.n555 VTAIL.n554 585
R1281 VTAIL.n582 VTAIL.n581 585
R1282 VTAIL.n580 VTAIL.n579 585
R1283 VTAIL.n559 VTAIL.n558 585
R1284 VTAIL.n574 VTAIL.n573 585
R1285 VTAIL.n572 VTAIL.n571 585
R1286 VTAIL.n563 VTAIL.n562 585
R1287 VTAIL.n566 VTAIL.n565 585
R1288 VTAIL.n525 VTAIL.n524 585
R1289 VTAIL.n523 VTAIL.n522 585
R1290 VTAIL.n428 VTAIL.n427 585
R1291 VTAIL.n517 VTAIL.n516 585
R1292 VTAIL.n515 VTAIL.n514 585
R1293 VTAIL.n432 VTAIL.n431 585
R1294 VTAIL.n509 VTAIL.n508 585
R1295 VTAIL.n507 VTAIL.n506 585
R1296 VTAIL.n505 VTAIL.n435 585
R1297 VTAIL.n439 VTAIL.n436 585
R1298 VTAIL.n500 VTAIL.n499 585
R1299 VTAIL.n498 VTAIL.n497 585
R1300 VTAIL.n441 VTAIL.n440 585
R1301 VTAIL.n492 VTAIL.n491 585
R1302 VTAIL.n490 VTAIL.n489 585
R1303 VTAIL.n445 VTAIL.n444 585
R1304 VTAIL.n484 VTAIL.n483 585
R1305 VTAIL.n482 VTAIL.n481 585
R1306 VTAIL.n449 VTAIL.n448 585
R1307 VTAIL.n476 VTAIL.n475 585
R1308 VTAIL.n474 VTAIL.n473 585
R1309 VTAIL.n453 VTAIL.n452 585
R1310 VTAIL.n468 VTAIL.n467 585
R1311 VTAIL.n466 VTAIL.n465 585
R1312 VTAIL.n457 VTAIL.n456 585
R1313 VTAIL.n460 VTAIL.n459 585
R1314 VTAIL.n419 VTAIL.n418 585
R1315 VTAIL.n417 VTAIL.n416 585
R1316 VTAIL.n322 VTAIL.n321 585
R1317 VTAIL.n411 VTAIL.n410 585
R1318 VTAIL.n409 VTAIL.n408 585
R1319 VTAIL.n326 VTAIL.n325 585
R1320 VTAIL.n403 VTAIL.n402 585
R1321 VTAIL.n401 VTAIL.n400 585
R1322 VTAIL.n399 VTAIL.n329 585
R1323 VTAIL.n333 VTAIL.n330 585
R1324 VTAIL.n394 VTAIL.n393 585
R1325 VTAIL.n392 VTAIL.n391 585
R1326 VTAIL.n335 VTAIL.n334 585
R1327 VTAIL.n386 VTAIL.n385 585
R1328 VTAIL.n384 VTAIL.n383 585
R1329 VTAIL.n339 VTAIL.n338 585
R1330 VTAIL.n378 VTAIL.n377 585
R1331 VTAIL.n376 VTAIL.n375 585
R1332 VTAIL.n343 VTAIL.n342 585
R1333 VTAIL.n370 VTAIL.n369 585
R1334 VTAIL.n368 VTAIL.n367 585
R1335 VTAIL.n347 VTAIL.n346 585
R1336 VTAIL.n362 VTAIL.n361 585
R1337 VTAIL.n360 VTAIL.n359 585
R1338 VTAIL.n351 VTAIL.n350 585
R1339 VTAIL.n354 VTAIL.n353 585
R1340 VTAIL.t3 VTAIL.n670 327.466
R1341 VTAIL.t0 VTAIL.n564 327.466
R1342 VTAIL.t5 VTAIL.n458 327.466
R1343 VTAIL.t4 VTAIL.n352 327.466
R1344 VTAIL.t6 VTAIL.n775 327.466
R1345 VTAIL.t7 VTAIL.n33 327.466
R1346 VTAIL.t2 VTAIL.n139 327.466
R1347 VTAIL.t1 VTAIL.n245 327.466
R1348 VTAIL.n776 VTAIL.n773 171.744
R1349 VTAIL.n783 VTAIL.n773 171.744
R1350 VTAIL.n784 VTAIL.n783 171.744
R1351 VTAIL.n784 VTAIL.n769 171.744
R1352 VTAIL.n791 VTAIL.n769 171.744
R1353 VTAIL.n792 VTAIL.n791 171.744
R1354 VTAIL.n792 VTAIL.n765 171.744
R1355 VTAIL.n799 VTAIL.n765 171.744
R1356 VTAIL.n800 VTAIL.n799 171.744
R1357 VTAIL.n800 VTAIL.n761 171.744
R1358 VTAIL.n807 VTAIL.n761 171.744
R1359 VTAIL.n808 VTAIL.n807 171.744
R1360 VTAIL.n808 VTAIL.n757 171.744
R1361 VTAIL.n815 VTAIL.n757 171.744
R1362 VTAIL.n817 VTAIL.n815 171.744
R1363 VTAIL.n817 VTAIL.n816 171.744
R1364 VTAIL.n816 VTAIL.n753 171.744
R1365 VTAIL.n825 VTAIL.n753 171.744
R1366 VTAIL.n826 VTAIL.n825 171.744
R1367 VTAIL.n826 VTAIL.n749 171.744
R1368 VTAIL.n833 VTAIL.n749 171.744
R1369 VTAIL.n834 VTAIL.n833 171.744
R1370 VTAIL.n834 VTAIL.n745 171.744
R1371 VTAIL.n841 VTAIL.n745 171.744
R1372 VTAIL.n842 VTAIL.n841 171.744
R1373 VTAIL.n34 VTAIL.n31 171.744
R1374 VTAIL.n41 VTAIL.n31 171.744
R1375 VTAIL.n42 VTAIL.n41 171.744
R1376 VTAIL.n42 VTAIL.n27 171.744
R1377 VTAIL.n49 VTAIL.n27 171.744
R1378 VTAIL.n50 VTAIL.n49 171.744
R1379 VTAIL.n50 VTAIL.n23 171.744
R1380 VTAIL.n57 VTAIL.n23 171.744
R1381 VTAIL.n58 VTAIL.n57 171.744
R1382 VTAIL.n58 VTAIL.n19 171.744
R1383 VTAIL.n65 VTAIL.n19 171.744
R1384 VTAIL.n66 VTAIL.n65 171.744
R1385 VTAIL.n66 VTAIL.n15 171.744
R1386 VTAIL.n73 VTAIL.n15 171.744
R1387 VTAIL.n75 VTAIL.n73 171.744
R1388 VTAIL.n75 VTAIL.n74 171.744
R1389 VTAIL.n74 VTAIL.n11 171.744
R1390 VTAIL.n83 VTAIL.n11 171.744
R1391 VTAIL.n84 VTAIL.n83 171.744
R1392 VTAIL.n84 VTAIL.n7 171.744
R1393 VTAIL.n91 VTAIL.n7 171.744
R1394 VTAIL.n92 VTAIL.n91 171.744
R1395 VTAIL.n92 VTAIL.n3 171.744
R1396 VTAIL.n99 VTAIL.n3 171.744
R1397 VTAIL.n100 VTAIL.n99 171.744
R1398 VTAIL.n140 VTAIL.n137 171.744
R1399 VTAIL.n147 VTAIL.n137 171.744
R1400 VTAIL.n148 VTAIL.n147 171.744
R1401 VTAIL.n148 VTAIL.n133 171.744
R1402 VTAIL.n155 VTAIL.n133 171.744
R1403 VTAIL.n156 VTAIL.n155 171.744
R1404 VTAIL.n156 VTAIL.n129 171.744
R1405 VTAIL.n163 VTAIL.n129 171.744
R1406 VTAIL.n164 VTAIL.n163 171.744
R1407 VTAIL.n164 VTAIL.n125 171.744
R1408 VTAIL.n171 VTAIL.n125 171.744
R1409 VTAIL.n172 VTAIL.n171 171.744
R1410 VTAIL.n172 VTAIL.n121 171.744
R1411 VTAIL.n179 VTAIL.n121 171.744
R1412 VTAIL.n181 VTAIL.n179 171.744
R1413 VTAIL.n181 VTAIL.n180 171.744
R1414 VTAIL.n180 VTAIL.n117 171.744
R1415 VTAIL.n189 VTAIL.n117 171.744
R1416 VTAIL.n190 VTAIL.n189 171.744
R1417 VTAIL.n190 VTAIL.n113 171.744
R1418 VTAIL.n197 VTAIL.n113 171.744
R1419 VTAIL.n198 VTAIL.n197 171.744
R1420 VTAIL.n198 VTAIL.n109 171.744
R1421 VTAIL.n205 VTAIL.n109 171.744
R1422 VTAIL.n206 VTAIL.n205 171.744
R1423 VTAIL.n246 VTAIL.n243 171.744
R1424 VTAIL.n253 VTAIL.n243 171.744
R1425 VTAIL.n254 VTAIL.n253 171.744
R1426 VTAIL.n254 VTAIL.n239 171.744
R1427 VTAIL.n261 VTAIL.n239 171.744
R1428 VTAIL.n262 VTAIL.n261 171.744
R1429 VTAIL.n262 VTAIL.n235 171.744
R1430 VTAIL.n269 VTAIL.n235 171.744
R1431 VTAIL.n270 VTAIL.n269 171.744
R1432 VTAIL.n270 VTAIL.n231 171.744
R1433 VTAIL.n277 VTAIL.n231 171.744
R1434 VTAIL.n278 VTAIL.n277 171.744
R1435 VTAIL.n278 VTAIL.n227 171.744
R1436 VTAIL.n285 VTAIL.n227 171.744
R1437 VTAIL.n287 VTAIL.n285 171.744
R1438 VTAIL.n287 VTAIL.n286 171.744
R1439 VTAIL.n286 VTAIL.n223 171.744
R1440 VTAIL.n295 VTAIL.n223 171.744
R1441 VTAIL.n296 VTAIL.n295 171.744
R1442 VTAIL.n296 VTAIL.n219 171.744
R1443 VTAIL.n303 VTAIL.n219 171.744
R1444 VTAIL.n304 VTAIL.n303 171.744
R1445 VTAIL.n304 VTAIL.n215 171.744
R1446 VTAIL.n311 VTAIL.n215 171.744
R1447 VTAIL.n312 VTAIL.n311 171.744
R1448 VTAIL.n736 VTAIL.n735 171.744
R1449 VTAIL.n735 VTAIL.n639 171.744
R1450 VTAIL.n728 VTAIL.n639 171.744
R1451 VTAIL.n728 VTAIL.n727 171.744
R1452 VTAIL.n727 VTAIL.n643 171.744
R1453 VTAIL.n720 VTAIL.n643 171.744
R1454 VTAIL.n720 VTAIL.n719 171.744
R1455 VTAIL.n719 VTAIL.n647 171.744
R1456 VTAIL.n651 VTAIL.n647 171.744
R1457 VTAIL.n711 VTAIL.n651 171.744
R1458 VTAIL.n711 VTAIL.n710 171.744
R1459 VTAIL.n710 VTAIL.n652 171.744
R1460 VTAIL.n703 VTAIL.n652 171.744
R1461 VTAIL.n703 VTAIL.n702 171.744
R1462 VTAIL.n702 VTAIL.n656 171.744
R1463 VTAIL.n695 VTAIL.n656 171.744
R1464 VTAIL.n695 VTAIL.n694 171.744
R1465 VTAIL.n694 VTAIL.n660 171.744
R1466 VTAIL.n687 VTAIL.n660 171.744
R1467 VTAIL.n687 VTAIL.n686 171.744
R1468 VTAIL.n686 VTAIL.n664 171.744
R1469 VTAIL.n679 VTAIL.n664 171.744
R1470 VTAIL.n679 VTAIL.n678 171.744
R1471 VTAIL.n678 VTAIL.n668 171.744
R1472 VTAIL.n671 VTAIL.n668 171.744
R1473 VTAIL.n630 VTAIL.n629 171.744
R1474 VTAIL.n629 VTAIL.n533 171.744
R1475 VTAIL.n622 VTAIL.n533 171.744
R1476 VTAIL.n622 VTAIL.n621 171.744
R1477 VTAIL.n621 VTAIL.n537 171.744
R1478 VTAIL.n614 VTAIL.n537 171.744
R1479 VTAIL.n614 VTAIL.n613 171.744
R1480 VTAIL.n613 VTAIL.n541 171.744
R1481 VTAIL.n545 VTAIL.n541 171.744
R1482 VTAIL.n605 VTAIL.n545 171.744
R1483 VTAIL.n605 VTAIL.n604 171.744
R1484 VTAIL.n604 VTAIL.n546 171.744
R1485 VTAIL.n597 VTAIL.n546 171.744
R1486 VTAIL.n597 VTAIL.n596 171.744
R1487 VTAIL.n596 VTAIL.n550 171.744
R1488 VTAIL.n589 VTAIL.n550 171.744
R1489 VTAIL.n589 VTAIL.n588 171.744
R1490 VTAIL.n588 VTAIL.n554 171.744
R1491 VTAIL.n581 VTAIL.n554 171.744
R1492 VTAIL.n581 VTAIL.n580 171.744
R1493 VTAIL.n580 VTAIL.n558 171.744
R1494 VTAIL.n573 VTAIL.n558 171.744
R1495 VTAIL.n573 VTAIL.n572 171.744
R1496 VTAIL.n572 VTAIL.n562 171.744
R1497 VTAIL.n565 VTAIL.n562 171.744
R1498 VTAIL.n524 VTAIL.n523 171.744
R1499 VTAIL.n523 VTAIL.n427 171.744
R1500 VTAIL.n516 VTAIL.n427 171.744
R1501 VTAIL.n516 VTAIL.n515 171.744
R1502 VTAIL.n515 VTAIL.n431 171.744
R1503 VTAIL.n508 VTAIL.n431 171.744
R1504 VTAIL.n508 VTAIL.n507 171.744
R1505 VTAIL.n507 VTAIL.n435 171.744
R1506 VTAIL.n439 VTAIL.n435 171.744
R1507 VTAIL.n499 VTAIL.n439 171.744
R1508 VTAIL.n499 VTAIL.n498 171.744
R1509 VTAIL.n498 VTAIL.n440 171.744
R1510 VTAIL.n491 VTAIL.n440 171.744
R1511 VTAIL.n491 VTAIL.n490 171.744
R1512 VTAIL.n490 VTAIL.n444 171.744
R1513 VTAIL.n483 VTAIL.n444 171.744
R1514 VTAIL.n483 VTAIL.n482 171.744
R1515 VTAIL.n482 VTAIL.n448 171.744
R1516 VTAIL.n475 VTAIL.n448 171.744
R1517 VTAIL.n475 VTAIL.n474 171.744
R1518 VTAIL.n474 VTAIL.n452 171.744
R1519 VTAIL.n467 VTAIL.n452 171.744
R1520 VTAIL.n467 VTAIL.n466 171.744
R1521 VTAIL.n466 VTAIL.n456 171.744
R1522 VTAIL.n459 VTAIL.n456 171.744
R1523 VTAIL.n418 VTAIL.n417 171.744
R1524 VTAIL.n417 VTAIL.n321 171.744
R1525 VTAIL.n410 VTAIL.n321 171.744
R1526 VTAIL.n410 VTAIL.n409 171.744
R1527 VTAIL.n409 VTAIL.n325 171.744
R1528 VTAIL.n402 VTAIL.n325 171.744
R1529 VTAIL.n402 VTAIL.n401 171.744
R1530 VTAIL.n401 VTAIL.n329 171.744
R1531 VTAIL.n333 VTAIL.n329 171.744
R1532 VTAIL.n393 VTAIL.n333 171.744
R1533 VTAIL.n393 VTAIL.n392 171.744
R1534 VTAIL.n392 VTAIL.n334 171.744
R1535 VTAIL.n385 VTAIL.n334 171.744
R1536 VTAIL.n385 VTAIL.n384 171.744
R1537 VTAIL.n384 VTAIL.n338 171.744
R1538 VTAIL.n377 VTAIL.n338 171.744
R1539 VTAIL.n377 VTAIL.n376 171.744
R1540 VTAIL.n376 VTAIL.n342 171.744
R1541 VTAIL.n369 VTAIL.n342 171.744
R1542 VTAIL.n369 VTAIL.n368 171.744
R1543 VTAIL.n368 VTAIL.n346 171.744
R1544 VTAIL.n361 VTAIL.n346 171.744
R1545 VTAIL.n361 VTAIL.n360 171.744
R1546 VTAIL.n360 VTAIL.n350 171.744
R1547 VTAIL.n353 VTAIL.n350 171.744
R1548 VTAIL.n776 VTAIL.t6 85.8723
R1549 VTAIL.n34 VTAIL.t7 85.8723
R1550 VTAIL.n140 VTAIL.t2 85.8723
R1551 VTAIL.n246 VTAIL.t1 85.8723
R1552 VTAIL.n671 VTAIL.t3 85.8723
R1553 VTAIL.n565 VTAIL.t0 85.8723
R1554 VTAIL.n459 VTAIL.t5 85.8723
R1555 VTAIL.n353 VTAIL.t4 85.8723
R1556 VTAIL.n847 VTAIL.n846 32.3793
R1557 VTAIL.n105 VTAIL.n104 32.3793
R1558 VTAIL.n211 VTAIL.n210 32.3793
R1559 VTAIL.n317 VTAIL.n316 32.3793
R1560 VTAIL.n741 VTAIL.n740 32.3793
R1561 VTAIL.n635 VTAIL.n634 32.3793
R1562 VTAIL.n529 VTAIL.n528 32.3793
R1563 VTAIL.n423 VTAIL.n422 32.3793
R1564 VTAIL.n847 VTAIL.n741 30.1686
R1565 VTAIL.n423 VTAIL.n317 30.1686
R1566 VTAIL.n777 VTAIL.n775 16.3895
R1567 VTAIL.n35 VTAIL.n33 16.3895
R1568 VTAIL.n141 VTAIL.n139 16.3895
R1569 VTAIL.n247 VTAIL.n245 16.3895
R1570 VTAIL.n672 VTAIL.n670 16.3895
R1571 VTAIL.n566 VTAIL.n564 16.3895
R1572 VTAIL.n460 VTAIL.n458 16.3895
R1573 VTAIL.n354 VTAIL.n352 16.3895
R1574 VTAIL.n824 VTAIL.n823 13.1884
R1575 VTAIL.n82 VTAIL.n81 13.1884
R1576 VTAIL.n188 VTAIL.n187 13.1884
R1577 VTAIL.n294 VTAIL.n293 13.1884
R1578 VTAIL.n718 VTAIL.n717 13.1884
R1579 VTAIL.n612 VTAIL.n611 13.1884
R1580 VTAIL.n506 VTAIL.n505 13.1884
R1581 VTAIL.n400 VTAIL.n399 13.1884
R1582 VTAIL.n778 VTAIL.n774 12.8005
R1583 VTAIL.n822 VTAIL.n754 12.8005
R1584 VTAIL.n827 VTAIL.n752 12.8005
R1585 VTAIL.n36 VTAIL.n32 12.8005
R1586 VTAIL.n80 VTAIL.n12 12.8005
R1587 VTAIL.n85 VTAIL.n10 12.8005
R1588 VTAIL.n142 VTAIL.n138 12.8005
R1589 VTAIL.n186 VTAIL.n118 12.8005
R1590 VTAIL.n191 VTAIL.n116 12.8005
R1591 VTAIL.n248 VTAIL.n244 12.8005
R1592 VTAIL.n292 VTAIL.n224 12.8005
R1593 VTAIL.n297 VTAIL.n222 12.8005
R1594 VTAIL.n721 VTAIL.n646 12.8005
R1595 VTAIL.n716 VTAIL.n648 12.8005
R1596 VTAIL.n673 VTAIL.n669 12.8005
R1597 VTAIL.n615 VTAIL.n540 12.8005
R1598 VTAIL.n610 VTAIL.n542 12.8005
R1599 VTAIL.n567 VTAIL.n563 12.8005
R1600 VTAIL.n509 VTAIL.n434 12.8005
R1601 VTAIL.n504 VTAIL.n436 12.8005
R1602 VTAIL.n461 VTAIL.n457 12.8005
R1603 VTAIL.n403 VTAIL.n328 12.8005
R1604 VTAIL.n398 VTAIL.n330 12.8005
R1605 VTAIL.n355 VTAIL.n351 12.8005
R1606 VTAIL.n782 VTAIL.n781 12.0247
R1607 VTAIL.n819 VTAIL.n818 12.0247
R1608 VTAIL.n828 VTAIL.n750 12.0247
R1609 VTAIL.n40 VTAIL.n39 12.0247
R1610 VTAIL.n77 VTAIL.n76 12.0247
R1611 VTAIL.n86 VTAIL.n8 12.0247
R1612 VTAIL.n146 VTAIL.n145 12.0247
R1613 VTAIL.n183 VTAIL.n182 12.0247
R1614 VTAIL.n192 VTAIL.n114 12.0247
R1615 VTAIL.n252 VTAIL.n251 12.0247
R1616 VTAIL.n289 VTAIL.n288 12.0247
R1617 VTAIL.n298 VTAIL.n220 12.0247
R1618 VTAIL.n722 VTAIL.n644 12.0247
R1619 VTAIL.n713 VTAIL.n712 12.0247
R1620 VTAIL.n677 VTAIL.n676 12.0247
R1621 VTAIL.n616 VTAIL.n538 12.0247
R1622 VTAIL.n607 VTAIL.n606 12.0247
R1623 VTAIL.n571 VTAIL.n570 12.0247
R1624 VTAIL.n510 VTAIL.n432 12.0247
R1625 VTAIL.n501 VTAIL.n500 12.0247
R1626 VTAIL.n465 VTAIL.n464 12.0247
R1627 VTAIL.n404 VTAIL.n326 12.0247
R1628 VTAIL.n395 VTAIL.n394 12.0247
R1629 VTAIL.n359 VTAIL.n358 12.0247
R1630 VTAIL.n785 VTAIL.n772 11.249
R1631 VTAIL.n814 VTAIL.n756 11.249
R1632 VTAIL.n832 VTAIL.n831 11.249
R1633 VTAIL.n43 VTAIL.n30 11.249
R1634 VTAIL.n72 VTAIL.n14 11.249
R1635 VTAIL.n90 VTAIL.n89 11.249
R1636 VTAIL.n149 VTAIL.n136 11.249
R1637 VTAIL.n178 VTAIL.n120 11.249
R1638 VTAIL.n196 VTAIL.n195 11.249
R1639 VTAIL.n255 VTAIL.n242 11.249
R1640 VTAIL.n284 VTAIL.n226 11.249
R1641 VTAIL.n302 VTAIL.n301 11.249
R1642 VTAIL.n726 VTAIL.n725 11.249
R1643 VTAIL.n709 VTAIL.n650 11.249
R1644 VTAIL.n680 VTAIL.n667 11.249
R1645 VTAIL.n620 VTAIL.n619 11.249
R1646 VTAIL.n603 VTAIL.n544 11.249
R1647 VTAIL.n574 VTAIL.n561 11.249
R1648 VTAIL.n514 VTAIL.n513 11.249
R1649 VTAIL.n497 VTAIL.n438 11.249
R1650 VTAIL.n468 VTAIL.n455 11.249
R1651 VTAIL.n408 VTAIL.n407 11.249
R1652 VTAIL.n391 VTAIL.n332 11.249
R1653 VTAIL.n362 VTAIL.n349 11.249
R1654 VTAIL.n786 VTAIL.n770 10.4732
R1655 VTAIL.n813 VTAIL.n758 10.4732
R1656 VTAIL.n835 VTAIL.n748 10.4732
R1657 VTAIL.n44 VTAIL.n28 10.4732
R1658 VTAIL.n71 VTAIL.n16 10.4732
R1659 VTAIL.n93 VTAIL.n6 10.4732
R1660 VTAIL.n150 VTAIL.n134 10.4732
R1661 VTAIL.n177 VTAIL.n122 10.4732
R1662 VTAIL.n199 VTAIL.n112 10.4732
R1663 VTAIL.n256 VTAIL.n240 10.4732
R1664 VTAIL.n283 VTAIL.n228 10.4732
R1665 VTAIL.n305 VTAIL.n218 10.4732
R1666 VTAIL.n729 VTAIL.n642 10.4732
R1667 VTAIL.n708 VTAIL.n653 10.4732
R1668 VTAIL.n681 VTAIL.n665 10.4732
R1669 VTAIL.n623 VTAIL.n536 10.4732
R1670 VTAIL.n602 VTAIL.n547 10.4732
R1671 VTAIL.n575 VTAIL.n559 10.4732
R1672 VTAIL.n517 VTAIL.n430 10.4732
R1673 VTAIL.n496 VTAIL.n441 10.4732
R1674 VTAIL.n469 VTAIL.n453 10.4732
R1675 VTAIL.n411 VTAIL.n324 10.4732
R1676 VTAIL.n390 VTAIL.n335 10.4732
R1677 VTAIL.n363 VTAIL.n347 10.4732
R1678 VTAIL.n790 VTAIL.n789 9.69747
R1679 VTAIL.n810 VTAIL.n809 9.69747
R1680 VTAIL.n836 VTAIL.n746 9.69747
R1681 VTAIL.n48 VTAIL.n47 9.69747
R1682 VTAIL.n68 VTAIL.n67 9.69747
R1683 VTAIL.n94 VTAIL.n4 9.69747
R1684 VTAIL.n154 VTAIL.n153 9.69747
R1685 VTAIL.n174 VTAIL.n173 9.69747
R1686 VTAIL.n200 VTAIL.n110 9.69747
R1687 VTAIL.n260 VTAIL.n259 9.69747
R1688 VTAIL.n280 VTAIL.n279 9.69747
R1689 VTAIL.n306 VTAIL.n216 9.69747
R1690 VTAIL.n730 VTAIL.n640 9.69747
R1691 VTAIL.n705 VTAIL.n704 9.69747
R1692 VTAIL.n685 VTAIL.n684 9.69747
R1693 VTAIL.n624 VTAIL.n534 9.69747
R1694 VTAIL.n599 VTAIL.n598 9.69747
R1695 VTAIL.n579 VTAIL.n578 9.69747
R1696 VTAIL.n518 VTAIL.n428 9.69747
R1697 VTAIL.n493 VTAIL.n492 9.69747
R1698 VTAIL.n473 VTAIL.n472 9.69747
R1699 VTAIL.n412 VTAIL.n322 9.69747
R1700 VTAIL.n387 VTAIL.n386 9.69747
R1701 VTAIL.n367 VTAIL.n366 9.69747
R1702 VTAIL.n846 VTAIL.n845 9.45567
R1703 VTAIL.n104 VTAIL.n103 9.45567
R1704 VTAIL.n210 VTAIL.n209 9.45567
R1705 VTAIL.n316 VTAIL.n315 9.45567
R1706 VTAIL.n740 VTAIL.n739 9.45567
R1707 VTAIL.n634 VTAIL.n633 9.45567
R1708 VTAIL.n528 VTAIL.n527 9.45567
R1709 VTAIL.n422 VTAIL.n421 9.45567
R1710 VTAIL.n744 VTAIL.n743 9.3005
R1711 VTAIL.n839 VTAIL.n838 9.3005
R1712 VTAIL.n837 VTAIL.n836 9.3005
R1713 VTAIL.n748 VTAIL.n747 9.3005
R1714 VTAIL.n831 VTAIL.n830 9.3005
R1715 VTAIL.n829 VTAIL.n828 9.3005
R1716 VTAIL.n752 VTAIL.n751 9.3005
R1717 VTAIL.n797 VTAIL.n796 9.3005
R1718 VTAIL.n795 VTAIL.n794 9.3005
R1719 VTAIL.n768 VTAIL.n767 9.3005
R1720 VTAIL.n789 VTAIL.n788 9.3005
R1721 VTAIL.n787 VTAIL.n786 9.3005
R1722 VTAIL.n772 VTAIL.n771 9.3005
R1723 VTAIL.n781 VTAIL.n780 9.3005
R1724 VTAIL.n779 VTAIL.n778 9.3005
R1725 VTAIL.n764 VTAIL.n763 9.3005
R1726 VTAIL.n803 VTAIL.n802 9.3005
R1727 VTAIL.n805 VTAIL.n804 9.3005
R1728 VTAIL.n760 VTAIL.n759 9.3005
R1729 VTAIL.n811 VTAIL.n810 9.3005
R1730 VTAIL.n813 VTAIL.n812 9.3005
R1731 VTAIL.n756 VTAIL.n755 9.3005
R1732 VTAIL.n820 VTAIL.n819 9.3005
R1733 VTAIL.n822 VTAIL.n821 9.3005
R1734 VTAIL.n845 VTAIL.n844 9.3005
R1735 VTAIL.n2 VTAIL.n1 9.3005
R1736 VTAIL.n97 VTAIL.n96 9.3005
R1737 VTAIL.n95 VTAIL.n94 9.3005
R1738 VTAIL.n6 VTAIL.n5 9.3005
R1739 VTAIL.n89 VTAIL.n88 9.3005
R1740 VTAIL.n87 VTAIL.n86 9.3005
R1741 VTAIL.n10 VTAIL.n9 9.3005
R1742 VTAIL.n55 VTAIL.n54 9.3005
R1743 VTAIL.n53 VTAIL.n52 9.3005
R1744 VTAIL.n26 VTAIL.n25 9.3005
R1745 VTAIL.n47 VTAIL.n46 9.3005
R1746 VTAIL.n45 VTAIL.n44 9.3005
R1747 VTAIL.n30 VTAIL.n29 9.3005
R1748 VTAIL.n39 VTAIL.n38 9.3005
R1749 VTAIL.n37 VTAIL.n36 9.3005
R1750 VTAIL.n22 VTAIL.n21 9.3005
R1751 VTAIL.n61 VTAIL.n60 9.3005
R1752 VTAIL.n63 VTAIL.n62 9.3005
R1753 VTAIL.n18 VTAIL.n17 9.3005
R1754 VTAIL.n69 VTAIL.n68 9.3005
R1755 VTAIL.n71 VTAIL.n70 9.3005
R1756 VTAIL.n14 VTAIL.n13 9.3005
R1757 VTAIL.n78 VTAIL.n77 9.3005
R1758 VTAIL.n80 VTAIL.n79 9.3005
R1759 VTAIL.n103 VTAIL.n102 9.3005
R1760 VTAIL.n108 VTAIL.n107 9.3005
R1761 VTAIL.n203 VTAIL.n202 9.3005
R1762 VTAIL.n201 VTAIL.n200 9.3005
R1763 VTAIL.n112 VTAIL.n111 9.3005
R1764 VTAIL.n195 VTAIL.n194 9.3005
R1765 VTAIL.n193 VTAIL.n192 9.3005
R1766 VTAIL.n116 VTAIL.n115 9.3005
R1767 VTAIL.n161 VTAIL.n160 9.3005
R1768 VTAIL.n159 VTAIL.n158 9.3005
R1769 VTAIL.n132 VTAIL.n131 9.3005
R1770 VTAIL.n153 VTAIL.n152 9.3005
R1771 VTAIL.n151 VTAIL.n150 9.3005
R1772 VTAIL.n136 VTAIL.n135 9.3005
R1773 VTAIL.n145 VTAIL.n144 9.3005
R1774 VTAIL.n143 VTAIL.n142 9.3005
R1775 VTAIL.n128 VTAIL.n127 9.3005
R1776 VTAIL.n167 VTAIL.n166 9.3005
R1777 VTAIL.n169 VTAIL.n168 9.3005
R1778 VTAIL.n124 VTAIL.n123 9.3005
R1779 VTAIL.n175 VTAIL.n174 9.3005
R1780 VTAIL.n177 VTAIL.n176 9.3005
R1781 VTAIL.n120 VTAIL.n119 9.3005
R1782 VTAIL.n184 VTAIL.n183 9.3005
R1783 VTAIL.n186 VTAIL.n185 9.3005
R1784 VTAIL.n209 VTAIL.n208 9.3005
R1785 VTAIL.n214 VTAIL.n213 9.3005
R1786 VTAIL.n309 VTAIL.n308 9.3005
R1787 VTAIL.n307 VTAIL.n306 9.3005
R1788 VTAIL.n218 VTAIL.n217 9.3005
R1789 VTAIL.n301 VTAIL.n300 9.3005
R1790 VTAIL.n299 VTAIL.n298 9.3005
R1791 VTAIL.n222 VTAIL.n221 9.3005
R1792 VTAIL.n267 VTAIL.n266 9.3005
R1793 VTAIL.n265 VTAIL.n264 9.3005
R1794 VTAIL.n238 VTAIL.n237 9.3005
R1795 VTAIL.n259 VTAIL.n258 9.3005
R1796 VTAIL.n257 VTAIL.n256 9.3005
R1797 VTAIL.n242 VTAIL.n241 9.3005
R1798 VTAIL.n251 VTAIL.n250 9.3005
R1799 VTAIL.n249 VTAIL.n248 9.3005
R1800 VTAIL.n234 VTAIL.n233 9.3005
R1801 VTAIL.n273 VTAIL.n272 9.3005
R1802 VTAIL.n275 VTAIL.n274 9.3005
R1803 VTAIL.n230 VTAIL.n229 9.3005
R1804 VTAIL.n281 VTAIL.n280 9.3005
R1805 VTAIL.n283 VTAIL.n282 9.3005
R1806 VTAIL.n226 VTAIL.n225 9.3005
R1807 VTAIL.n290 VTAIL.n289 9.3005
R1808 VTAIL.n292 VTAIL.n291 9.3005
R1809 VTAIL.n315 VTAIL.n314 9.3005
R1810 VTAIL.n698 VTAIL.n697 9.3005
R1811 VTAIL.n700 VTAIL.n699 9.3005
R1812 VTAIL.n655 VTAIL.n654 9.3005
R1813 VTAIL.n706 VTAIL.n705 9.3005
R1814 VTAIL.n708 VTAIL.n707 9.3005
R1815 VTAIL.n650 VTAIL.n649 9.3005
R1816 VTAIL.n714 VTAIL.n713 9.3005
R1817 VTAIL.n716 VTAIL.n715 9.3005
R1818 VTAIL.n739 VTAIL.n738 9.3005
R1819 VTAIL.n638 VTAIL.n637 9.3005
R1820 VTAIL.n733 VTAIL.n732 9.3005
R1821 VTAIL.n731 VTAIL.n730 9.3005
R1822 VTAIL.n642 VTAIL.n641 9.3005
R1823 VTAIL.n725 VTAIL.n724 9.3005
R1824 VTAIL.n723 VTAIL.n722 9.3005
R1825 VTAIL.n646 VTAIL.n645 9.3005
R1826 VTAIL.n659 VTAIL.n658 9.3005
R1827 VTAIL.n692 VTAIL.n691 9.3005
R1828 VTAIL.n690 VTAIL.n689 9.3005
R1829 VTAIL.n663 VTAIL.n662 9.3005
R1830 VTAIL.n684 VTAIL.n683 9.3005
R1831 VTAIL.n682 VTAIL.n681 9.3005
R1832 VTAIL.n667 VTAIL.n666 9.3005
R1833 VTAIL.n676 VTAIL.n675 9.3005
R1834 VTAIL.n674 VTAIL.n673 9.3005
R1835 VTAIL.n592 VTAIL.n591 9.3005
R1836 VTAIL.n594 VTAIL.n593 9.3005
R1837 VTAIL.n549 VTAIL.n548 9.3005
R1838 VTAIL.n600 VTAIL.n599 9.3005
R1839 VTAIL.n602 VTAIL.n601 9.3005
R1840 VTAIL.n544 VTAIL.n543 9.3005
R1841 VTAIL.n608 VTAIL.n607 9.3005
R1842 VTAIL.n610 VTAIL.n609 9.3005
R1843 VTAIL.n633 VTAIL.n632 9.3005
R1844 VTAIL.n532 VTAIL.n531 9.3005
R1845 VTAIL.n627 VTAIL.n626 9.3005
R1846 VTAIL.n625 VTAIL.n624 9.3005
R1847 VTAIL.n536 VTAIL.n535 9.3005
R1848 VTAIL.n619 VTAIL.n618 9.3005
R1849 VTAIL.n617 VTAIL.n616 9.3005
R1850 VTAIL.n540 VTAIL.n539 9.3005
R1851 VTAIL.n553 VTAIL.n552 9.3005
R1852 VTAIL.n586 VTAIL.n585 9.3005
R1853 VTAIL.n584 VTAIL.n583 9.3005
R1854 VTAIL.n557 VTAIL.n556 9.3005
R1855 VTAIL.n578 VTAIL.n577 9.3005
R1856 VTAIL.n576 VTAIL.n575 9.3005
R1857 VTAIL.n561 VTAIL.n560 9.3005
R1858 VTAIL.n570 VTAIL.n569 9.3005
R1859 VTAIL.n568 VTAIL.n567 9.3005
R1860 VTAIL.n486 VTAIL.n485 9.3005
R1861 VTAIL.n488 VTAIL.n487 9.3005
R1862 VTAIL.n443 VTAIL.n442 9.3005
R1863 VTAIL.n494 VTAIL.n493 9.3005
R1864 VTAIL.n496 VTAIL.n495 9.3005
R1865 VTAIL.n438 VTAIL.n437 9.3005
R1866 VTAIL.n502 VTAIL.n501 9.3005
R1867 VTAIL.n504 VTAIL.n503 9.3005
R1868 VTAIL.n527 VTAIL.n526 9.3005
R1869 VTAIL.n426 VTAIL.n425 9.3005
R1870 VTAIL.n521 VTAIL.n520 9.3005
R1871 VTAIL.n519 VTAIL.n518 9.3005
R1872 VTAIL.n430 VTAIL.n429 9.3005
R1873 VTAIL.n513 VTAIL.n512 9.3005
R1874 VTAIL.n511 VTAIL.n510 9.3005
R1875 VTAIL.n434 VTAIL.n433 9.3005
R1876 VTAIL.n447 VTAIL.n446 9.3005
R1877 VTAIL.n480 VTAIL.n479 9.3005
R1878 VTAIL.n478 VTAIL.n477 9.3005
R1879 VTAIL.n451 VTAIL.n450 9.3005
R1880 VTAIL.n472 VTAIL.n471 9.3005
R1881 VTAIL.n470 VTAIL.n469 9.3005
R1882 VTAIL.n455 VTAIL.n454 9.3005
R1883 VTAIL.n464 VTAIL.n463 9.3005
R1884 VTAIL.n462 VTAIL.n461 9.3005
R1885 VTAIL.n380 VTAIL.n379 9.3005
R1886 VTAIL.n382 VTAIL.n381 9.3005
R1887 VTAIL.n337 VTAIL.n336 9.3005
R1888 VTAIL.n388 VTAIL.n387 9.3005
R1889 VTAIL.n390 VTAIL.n389 9.3005
R1890 VTAIL.n332 VTAIL.n331 9.3005
R1891 VTAIL.n396 VTAIL.n395 9.3005
R1892 VTAIL.n398 VTAIL.n397 9.3005
R1893 VTAIL.n421 VTAIL.n420 9.3005
R1894 VTAIL.n320 VTAIL.n319 9.3005
R1895 VTAIL.n415 VTAIL.n414 9.3005
R1896 VTAIL.n413 VTAIL.n412 9.3005
R1897 VTAIL.n324 VTAIL.n323 9.3005
R1898 VTAIL.n407 VTAIL.n406 9.3005
R1899 VTAIL.n405 VTAIL.n404 9.3005
R1900 VTAIL.n328 VTAIL.n327 9.3005
R1901 VTAIL.n341 VTAIL.n340 9.3005
R1902 VTAIL.n374 VTAIL.n373 9.3005
R1903 VTAIL.n372 VTAIL.n371 9.3005
R1904 VTAIL.n345 VTAIL.n344 9.3005
R1905 VTAIL.n366 VTAIL.n365 9.3005
R1906 VTAIL.n364 VTAIL.n363 9.3005
R1907 VTAIL.n349 VTAIL.n348 9.3005
R1908 VTAIL.n358 VTAIL.n357 9.3005
R1909 VTAIL.n356 VTAIL.n355 9.3005
R1910 VTAIL.n793 VTAIL.n768 8.92171
R1911 VTAIL.n806 VTAIL.n760 8.92171
R1912 VTAIL.n840 VTAIL.n839 8.92171
R1913 VTAIL.n51 VTAIL.n26 8.92171
R1914 VTAIL.n64 VTAIL.n18 8.92171
R1915 VTAIL.n98 VTAIL.n97 8.92171
R1916 VTAIL.n157 VTAIL.n132 8.92171
R1917 VTAIL.n170 VTAIL.n124 8.92171
R1918 VTAIL.n204 VTAIL.n203 8.92171
R1919 VTAIL.n263 VTAIL.n238 8.92171
R1920 VTAIL.n276 VTAIL.n230 8.92171
R1921 VTAIL.n310 VTAIL.n309 8.92171
R1922 VTAIL.n734 VTAIL.n733 8.92171
R1923 VTAIL.n701 VTAIL.n655 8.92171
R1924 VTAIL.n688 VTAIL.n663 8.92171
R1925 VTAIL.n628 VTAIL.n627 8.92171
R1926 VTAIL.n595 VTAIL.n549 8.92171
R1927 VTAIL.n582 VTAIL.n557 8.92171
R1928 VTAIL.n522 VTAIL.n521 8.92171
R1929 VTAIL.n489 VTAIL.n443 8.92171
R1930 VTAIL.n476 VTAIL.n451 8.92171
R1931 VTAIL.n416 VTAIL.n415 8.92171
R1932 VTAIL.n383 VTAIL.n337 8.92171
R1933 VTAIL.n370 VTAIL.n345 8.92171
R1934 VTAIL.n794 VTAIL.n766 8.14595
R1935 VTAIL.n805 VTAIL.n762 8.14595
R1936 VTAIL.n843 VTAIL.n744 8.14595
R1937 VTAIL.n52 VTAIL.n24 8.14595
R1938 VTAIL.n63 VTAIL.n20 8.14595
R1939 VTAIL.n101 VTAIL.n2 8.14595
R1940 VTAIL.n158 VTAIL.n130 8.14595
R1941 VTAIL.n169 VTAIL.n126 8.14595
R1942 VTAIL.n207 VTAIL.n108 8.14595
R1943 VTAIL.n264 VTAIL.n236 8.14595
R1944 VTAIL.n275 VTAIL.n232 8.14595
R1945 VTAIL.n313 VTAIL.n214 8.14595
R1946 VTAIL.n737 VTAIL.n638 8.14595
R1947 VTAIL.n700 VTAIL.n657 8.14595
R1948 VTAIL.n689 VTAIL.n661 8.14595
R1949 VTAIL.n631 VTAIL.n532 8.14595
R1950 VTAIL.n594 VTAIL.n551 8.14595
R1951 VTAIL.n583 VTAIL.n555 8.14595
R1952 VTAIL.n525 VTAIL.n426 8.14595
R1953 VTAIL.n488 VTAIL.n445 8.14595
R1954 VTAIL.n477 VTAIL.n449 8.14595
R1955 VTAIL.n419 VTAIL.n320 8.14595
R1956 VTAIL.n382 VTAIL.n339 8.14595
R1957 VTAIL.n371 VTAIL.n343 8.14595
R1958 VTAIL.n798 VTAIL.n797 7.3702
R1959 VTAIL.n802 VTAIL.n801 7.3702
R1960 VTAIL.n844 VTAIL.n742 7.3702
R1961 VTAIL.n56 VTAIL.n55 7.3702
R1962 VTAIL.n60 VTAIL.n59 7.3702
R1963 VTAIL.n102 VTAIL.n0 7.3702
R1964 VTAIL.n162 VTAIL.n161 7.3702
R1965 VTAIL.n166 VTAIL.n165 7.3702
R1966 VTAIL.n208 VTAIL.n106 7.3702
R1967 VTAIL.n268 VTAIL.n267 7.3702
R1968 VTAIL.n272 VTAIL.n271 7.3702
R1969 VTAIL.n314 VTAIL.n212 7.3702
R1970 VTAIL.n738 VTAIL.n636 7.3702
R1971 VTAIL.n697 VTAIL.n696 7.3702
R1972 VTAIL.n693 VTAIL.n692 7.3702
R1973 VTAIL.n632 VTAIL.n530 7.3702
R1974 VTAIL.n591 VTAIL.n590 7.3702
R1975 VTAIL.n587 VTAIL.n586 7.3702
R1976 VTAIL.n526 VTAIL.n424 7.3702
R1977 VTAIL.n485 VTAIL.n484 7.3702
R1978 VTAIL.n481 VTAIL.n480 7.3702
R1979 VTAIL.n420 VTAIL.n318 7.3702
R1980 VTAIL.n379 VTAIL.n378 7.3702
R1981 VTAIL.n375 VTAIL.n374 7.3702
R1982 VTAIL.n798 VTAIL.n764 6.59444
R1983 VTAIL.n801 VTAIL.n764 6.59444
R1984 VTAIL.n846 VTAIL.n742 6.59444
R1985 VTAIL.n56 VTAIL.n22 6.59444
R1986 VTAIL.n59 VTAIL.n22 6.59444
R1987 VTAIL.n104 VTAIL.n0 6.59444
R1988 VTAIL.n162 VTAIL.n128 6.59444
R1989 VTAIL.n165 VTAIL.n128 6.59444
R1990 VTAIL.n210 VTAIL.n106 6.59444
R1991 VTAIL.n268 VTAIL.n234 6.59444
R1992 VTAIL.n271 VTAIL.n234 6.59444
R1993 VTAIL.n316 VTAIL.n212 6.59444
R1994 VTAIL.n740 VTAIL.n636 6.59444
R1995 VTAIL.n696 VTAIL.n659 6.59444
R1996 VTAIL.n693 VTAIL.n659 6.59444
R1997 VTAIL.n634 VTAIL.n530 6.59444
R1998 VTAIL.n590 VTAIL.n553 6.59444
R1999 VTAIL.n587 VTAIL.n553 6.59444
R2000 VTAIL.n528 VTAIL.n424 6.59444
R2001 VTAIL.n484 VTAIL.n447 6.59444
R2002 VTAIL.n481 VTAIL.n447 6.59444
R2003 VTAIL.n422 VTAIL.n318 6.59444
R2004 VTAIL.n378 VTAIL.n341 6.59444
R2005 VTAIL.n375 VTAIL.n341 6.59444
R2006 VTAIL.n797 VTAIL.n766 5.81868
R2007 VTAIL.n802 VTAIL.n762 5.81868
R2008 VTAIL.n844 VTAIL.n843 5.81868
R2009 VTAIL.n55 VTAIL.n24 5.81868
R2010 VTAIL.n60 VTAIL.n20 5.81868
R2011 VTAIL.n102 VTAIL.n101 5.81868
R2012 VTAIL.n161 VTAIL.n130 5.81868
R2013 VTAIL.n166 VTAIL.n126 5.81868
R2014 VTAIL.n208 VTAIL.n207 5.81868
R2015 VTAIL.n267 VTAIL.n236 5.81868
R2016 VTAIL.n272 VTAIL.n232 5.81868
R2017 VTAIL.n314 VTAIL.n313 5.81868
R2018 VTAIL.n738 VTAIL.n737 5.81868
R2019 VTAIL.n697 VTAIL.n657 5.81868
R2020 VTAIL.n692 VTAIL.n661 5.81868
R2021 VTAIL.n632 VTAIL.n631 5.81868
R2022 VTAIL.n591 VTAIL.n551 5.81868
R2023 VTAIL.n586 VTAIL.n555 5.81868
R2024 VTAIL.n526 VTAIL.n525 5.81868
R2025 VTAIL.n485 VTAIL.n445 5.81868
R2026 VTAIL.n480 VTAIL.n449 5.81868
R2027 VTAIL.n420 VTAIL.n419 5.81868
R2028 VTAIL.n379 VTAIL.n339 5.81868
R2029 VTAIL.n374 VTAIL.n343 5.81868
R2030 VTAIL.n794 VTAIL.n793 5.04292
R2031 VTAIL.n806 VTAIL.n805 5.04292
R2032 VTAIL.n840 VTAIL.n744 5.04292
R2033 VTAIL.n52 VTAIL.n51 5.04292
R2034 VTAIL.n64 VTAIL.n63 5.04292
R2035 VTAIL.n98 VTAIL.n2 5.04292
R2036 VTAIL.n158 VTAIL.n157 5.04292
R2037 VTAIL.n170 VTAIL.n169 5.04292
R2038 VTAIL.n204 VTAIL.n108 5.04292
R2039 VTAIL.n264 VTAIL.n263 5.04292
R2040 VTAIL.n276 VTAIL.n275 5.04292
R2041 VTAIL.n310 VTAIL.n214 5.04292
R2042 VTAIL.n734 VTAIL.n638 5.04292
R2043 VTAIL.n701 VTAIL.n700 5.04292
R2044 VTAIL.n689 VTAIL.n688 5.04292
R2045 VTAIL.n628 VTAIL.n532 5.04292
R2046 VTAIL.n595 VTAIL.n594 5.04292
R2047 VTAIL.n583 VTAIL.n582 5.04292
R2048 VTAIL.n522 VTAIL.n426 5.04292
R2049 VTAIL.n489 VTAIL.n488 5.04292
R2050 VTAIL.n477 VTAIL.n476 5.04292
R2051 VTAIL.n416 VTAIL.n320 5.04292
R2052 VTAIL.n383 VTAIL.n382 5.04292
R2053 VTAIL.n371 VTAIL.n370 5.04292
R2054 VTAIL.n790 VTAIL.n768 4.26717
R2055 VTAIL.n809 VTAIL.n760 4.26717
R2056 VTAIL.n839 VTAIL.n746 4.26717
R2057 VTAIL.n48 VTAIL.n26 4.26717
R2058 VTAIL.n67 VTAIL.n18 4.26717
R2059 VTAIL.n97 VTAIL.n4 4.26717
R2060 VTAIL.n154 VTAIL.n132 4.26717
R2061 VTAIL.n173 VTAIL.n124 4.26717
R2062 VTAIL.n203 VTAIL.n110 4.26717
R2063 VTAIL.n260 VTAIL.n238 4.26717
R2064 VTAIL.n279 VTAIL.n230 4.26717
R2065 VTAIL.n309 VTAIL.n216 4.26717
R2066 VTAIL.n733 VTAIL.n640 4.26717
R2067 VTAIL.n704 VTAIL.n655 4.26717
R2068 VTAIL.n685 VTAIL.n663 4.26717
R2069 VTAIL.n627 VTAIL.n534 4.26717
R2070 VTAIL.n598 VTAIL.n549 4.26717
R2071 VTAIL.n579 VTAIL.n557 4.26717
R2072 VTAIL.n521 VTAIL.n428 4.26717
R2073 VTAIL.n492 VTAIL.n443 4.26717
R2074 VTAIL.n473 VTAIL.n451 4.26717
R2075 VTAIL.n415 VTAIL.n322 4.26717
R2076 VTAIL.n386 VTAIL.n337 4.26717
R2077 VTAIL.n367 VTAIL.n345 4.26717
R2078 VTAIL.n779 VTAIL.n775 3.70982
R2079 VTAIL.n37 VTAIL.n33 3.70982
R2080 VTAIL.n143 VTAIL.n139 3.70982
R2081 VTAIL.n249 VTAIL.n245 3.70982
R2082 VTAIL.n674 VTAIL.n670 3.70982
R2083 VTAIL.n568 VTAIL.n564 3.70982
R2084 VTAIL.n462 VTAIL.n458 3.70982
R2085 VTAIL.n356 VTAIL.n352 3.70982
R2086 VTAIL.n789 VTAIL.n770 3.49141
R2087 VTAIL.n810 VTAIL.n758 3.49141
R2088 VTAIL.n836 VTAIL.n835 3.49141
R2089 VTAIL.n47 VTAIL.n28 3.49141
R2090 VTAIL.n68 VTAIL.n16 3.49141
R2091 VTAIL.n94 VTAIL.n93 3.49141
R2092 VTAIL.n153 VTAIL.n134 3.49141
R2093 VTAIL.n174 VTAIL.n122 3.49141
R2094 VTAIL.n200 VTAIL.n199 3.49141
R2095 VTAIL.n259 VTAIL.n240 3.49141
R2096 VTAIL.n280 VTAIL.n228 3.49141
R2097 VTAIL.n306 VTAIL.n305 3.49141
R2098 VTAIL.n730 VTAIL.n729 3.49141
R2099 VTAIL.n705 VTAIL.n653 3.49141
R2100 VTAIL.n684 VTAIL.n665 3.49141
R2101 VTAIL.n624 VTAIL.n623 3.49141
R2102 VTAIL.n599 VTAIL.n547 3.49141
R2103 VTAIL.n578 VTAIL.n559 3.49141
R2104 VTAIL.n518 VTAIL.n517 3.49141
R2105 VTAIL.n493 VTAIL.n441 3.49141
R2106 VTAIL.n472 VTAIL.n453 3.49141
R2107 VTAIL.n412 VTAIL.n411 3.49141
R2108 VTAIL.n387 VTAIL.n335 3.49141
R2109 VTAIL.n366 VTAIL.n347 3.49141
R2110 VTAIL.n786 VTAIL.n785 2.71565
R2111 VTAIL.n814 VTAIL.n813 2.71565
R2112 VTAIL.n832 VTAIL.n748 2.71565
R2113 VTAIL.n44 VTAIL.n43 2.71565
R2114 VTAIL.n72 VTAIL.n71 2.71565
R2115 VTAIL.n90 VTAIL.n6 2.71565
R2116 VTAIL.n150 VTAIL.n149 2.71565
R2117 VTAIL.n178 VTAIL.n177 2.71565
R2118 VTAIL.n196 VTAIL.n112 2.71565
R2119 VTAIL.n256 VTAIL.n255 2.71565
R2120 VTAIL.n284 VTAIL.n283 2.71565
R2121 VTAIL.n302 VTAIL.n218 2.71565
R2122 VTAIL.n726 VTAIL.n642 2.71565
R2123 VTAIL.n709 VTAIL.n708 2.71565
R2124 VTAIL.n681 VTAIL.n680 2.71565
R2125 VTAIL.n620 VTAIL.n536 2.71565
R2126 VTAIL.n603 VTAIL.n602 2.71565
R2127 VTAIL.n575 VTAIL.n574 2.71565
R2128 VTAIL.n514 VTAIL.n430 2.71565
R2129 VTAIL.n497 VTAIL.n496 2.71565
R2130 VTAIL.n469 VTAIL.n468 2.71565
R2131 VTAIL.n408 VTAIL.n324 2.71565
R2132 VTAIL.n391 VTAIL.n390 2.71565
R2133 VTAIL.n363 VTAIL.n362 2.71565
R2134 VTAIL.n782 VTAIL.n772 1.93989
R2135 VTAIL.n818 VTAIL.n756 1.93989
R2136 VTAIL.n831 VTAIL.n750 1.93989
R2137 VTAIL.n40 VTAIL.n30 1.93989
R2138 VTAIL.n76 VTAIL.n14 1.93989
R2139 VTAIL.n89 VTAIL.n8 1.93989
R2140 VTAIL.n146 VTAIL.n136 1.93989
R2141 VTAIL.n182 VTAIL.n120 1.93989
R2142 VTAIL.n195 VTAIL.n114 1.93989
R2143 VTAIL.n252 VTAIL.n242 1.93989
R2144 VTAIL.n288 VTAIL.n226 1.93989
R2145 VTAIL.n301 VTAIL.n220 1.93989
R2146 VTAIL.n725 VTAIL.n644 1.93989
R2147 VTAIL.n712 VTAIL.n650 1.93989
R2148 VTAIL.n677 VTAIL.n667 1.93989
R2149 VTAIL.n619 VTAIL.n538 1.93989
R2150 VTAIL.n606 VTAIL.n544 1.93989
R2151 VTAIL.n571 VTAIL.n561 1.93989
R2152 VTAIL.n513 VTAIL.n432 1.93989
R2153 VTAIL.n500 VTAIL.n438 1.93989
R2154 VTAIL.n465 VTAIL.n455 1.93989
R2155 VTAIL.n407 VTAIL.n326 1.93989
R2156 VTAIL.n394 VTAIL.n332 1.93989
R2157 VTAIL.n359 VTAIL.n349 1.93989
R2158 VTAIL.n529 VTAIL.n423 1.44878
R2159 VTAIL.n741 VTAIL.n635 1.44878
R2160 VTAIL.n317 VTAIL.n211 1.44878
R2161 VTAIL.n781 VTAIL.n774 1.16414
R2162 VTAIL.n819 VTAIL.n754 1.16414
R2163 VTAIL.n828 VTAIL.n827 1.16414
R2164 VTAIL.n39 VTAIL.n32 1.16414
R2165 VTAIL.n77 VTAIL.n12 1.16414
R2166 VTAIL.n86 VTAIL.n85 1.16414
R2167 VTAIL.n145 VTAIL.n138 1.16414
R2168 VTAIL.n183 VTAIL.n118 1.16414
R2169 VTAIL.n192 VTAIL.n191 1.16414
R2170 VTAIL.n251 VTAIL.n244 1.16414
R2171 VTAIL.n289 VTAIL.n224 1.16414
R2172 VTAIL.n298 VTAIL.n297 1.16414
R2173 VTAIL.n722 VTAIL.n721 1.16414
R2174 VTAIL.n713 VTAIL.n648 1.16414
R2175 VTAIL.n676 VTAIL.n669 1.16414
R2176 VTAIL.n616 VTAIL.n615 1.16414
R2177 VTAIL.n607 VTAIL.n542 1.16414
R2178 VTAIL.n570 VTAIL.n563 1.16414
R2179 VTAIL.n510 VTAIL.n509 1.16414
R2180 VTAIL.n501 VTAIL.n436 1.16414
R2181 VTAIL.n464 VTAIL.n457 1.16414
R2182 VTAIL.n404 VTAIL.n403 1.16414
R2183 VTAIL.n395 VTAIL.n330 1.16414
R2184 VTAIL.n358 VTAIL.n351 1.16414
R2185 VTAIL VTAIL.n105 0.782828
R2186 VTAIL VTAIL.n847 0.666448
R2187 VTAIL.n635 VTAIL.n529 0.470328
R2188 VTAIL.n211 VTAIL.n105 0.470328
R2189 VTAIL.n778 VTAIL.n777 0.388379
R2190 VTAIL.n823 VTAIL.n822 0.388379
R2191 VTAIL.n824 VTAIL.n752 0.388379
R2192 VTAIL.n36 VTAIL.n35 0.388379
R2193 VTAIL.n81 VTAIL.n80 0.388379
R2194 VTAIL.n82 VTAIL.n10 0.388379
R2195 VTAIL.n142 VTAIL.n141 0.388379
R2196 VTAIL.n187 VTAIL.n186 0.388379
R2197 VTAIL.n188 VTAIL.n116 0.388379
R2198 VTAIL.n248 VTAIL.n247 0.388379
R2199 VTAIL.n293 VTAIL.n292 0.388379
R2200 VTAIL.n294 VTAIL.n222 0.388379
R2201 VTAIL.n718 VTAIL.n646 0.388379
R2202 VTAIL.n717 VTAIL.n716 0.388379
R2203 VTAIL.n673 VTAIL.n672 0.388379
R2204 VTAIL.n612 VTAIL.n540 0.388379
R2205 VTAIL.n611 VTAIL.n610 0.388379
R2206 VTAIL.n567 VTAIL.n566 0.388379
R2207 VTAIL.n506 VTAIL.n434 0.388379
R2208 VTAIL.n505 VTAIL.n504 0.388379
R2209 VTAIL.n461 VTAIL.n460 0.388379
R2210 VTAIL.n400 VTAIL.n328 0.388379
R2211 VTAIL.n399 VTAIL.n398 0.388379
R2212 VTAIL.n355 VTAIL.n354 0.388379
R2213 VTAIL.n780 VTAIL.n779 0.155672
R2214 VTAIL.n780 VTAIL.n771 0.155672
R2215 VTAIL.n787 VTAIL.n771 0.155672
R2216 VTAIL.n788 VTAIL.n787 0.155672
R2217 VTAIL.n788 VTAIL.n767 0.155672
R2218 VTAIL.n795 VTAIL.n767 0.155672
R2219 VTAIL.n796 VTAIL.n795 0.155672
R2220 VTAIL.n796 VTAIL.n763 0.155672
R2221 VTAIL.n803 VTAIL.n763 0.155672
R2222 VTAIL.n804 VTAIL.n803 0.155672
R2223 VTAIL.n804 VTAIL.n759 0.155672
R2224 VTAIL.n811 VTAIL.n759 0.155672
R2225 VTAIL.n812 VTAIL.n811 0.155672
R2226 VTAIL.n812 VTAIL.n755 0.155672
R2227 VTAIL.n820 VTAIL.n755 0.155672
R2228 VTAIL.n821 VTAIL.n820 0.155672
R2229 VTAIL.n821 VTAIL.n751 0.155672
R2230 VTAIL.n829 VTAIL.n751 0.155672
R2231 VTAIL.n830 VTAIL.n829 0.155672
R2232 VTAIL.n830 VTAIL.n747 0.155672
R2233 VTAIL.n837 VTAIL.n747 0.155672
R2234 VTAIL.n838 VTAIL.n837 0.155672
R2235 VTAIL.n838 VTAIL.n743 0.155672
R2236 VTAIL.n845 VTAIL.n743 0.155672
R2237 VTAIL.n38 VTAIL.n37 0.155672
R2238 VTAIL.n38 VTAIL.n29 0.155672
R2239 VTAIL.n45 VTAIL.n29 0.155672
R2240 VTAIL.n46 VTAIL.n45 0.155672
R2241 VTAIL.n46 VTAIL.n25 0.155672
R2242 VTAIL.n53 VTAIL.n25 0.155672
R2243 VTAIL.n54 VTAIL.n53 0.155672
R2244 VTAIL.n54 VTAIL.n21 0.155672
R2245 VTAIL.n61 VTAIL.n21 0.155672
R2246 VTAIL.n62 VTAIL.n61 0.155672
R2247 VTAIL.n62 VTAIL.n17 0.155672
R2248 VTAIL.n69 VTAIL.n17 0.155672
R2249 VTAIL.n70 VTAIL.n69 0.155672
R2250 VTAIL.n70 VTAIL.n13 0.155672
R2251 VTAIL.n78 VTAIL.n13 0.155672
R2252 VTAIL.n79 VTAIL.n78 0.155672
R2253 VTAIL.n79 VTAIL.n9 0.155672
R2254 VTAIL.n87 VTAIL.n9 0.155672
R2255 VTAIL.n88 VTAIL.n87 0.155672
R2256 VTAIL.n88 VTAIL.n5 0.155672
R2257 VTAIL.n95 VTAIL.n5 0.155672
R2258 VTAIL.n96 VTAIL.n95 0.155672
R2259 VTAIL.n96 VTAIL.n1 0.155672
R2260 VTAIL.n103 VTAIL.n1 0.155672
R2261 VTAIL.n144 VTAIL.n143 0.155672
R2262 VTAIL.n144 VTAIL.n135 0.155672
R2263 VTAIL.n151 VTAIL.n135 0.155672
R2264 VTAIL.n152 VTAIL.n151 0.155672
R2265 VTAIL.n152 VTAIL.n131 0.155672
R2266 VTAIL.n159 VTAIL.n131 0.155672
R2267 VTAIL.n160 VTAIL.n159 0.155672
R2268 VTAIL.n160 VTAIL.n127 0.155672
R2269 VTAIL.n167 VTAIL.n127 0.155672
R2270 VTAIL.n168 VTAIL.n167 0.155672
R2271 VTAIL.n168 VTAIL.n123 0.155672
R2272 VTAIL.n175 VTAIL.n123 0.155672
R2273 VTAIL.n176 VTAIL.n175 0.155672
R2274 VTAIL.n176 VTAIL.n119 0.155672
R2275 VTAIL.n184 VTAIL.n119 0.155672
R2276 VTAIL.n185 VTAIL.n184 0.155672
R2277 VTAIL.n185 VTAIL.n115 0.155672
R2278 VTAIL.n193 VTAIL.n115 0.155672
R2279 VTAIL.n194 VTAIL.n193 0.155672
R2280 VTAIL.n194 VTAIL.n111 0.155672
R2281 VTAIL.n201 VTAIL.n111 0.155672
R2282 VTAIL.n202 VTAIL.n201 0.155672
R2283 VTAIL.n202 VTAIL.n107 0.155672
R2284 VTAIL.n209 VTAIL.n107 0.155672
R2285 VTAIL.n250 VTAIL.n249 0.155672
R2286 VTAIL.n250 VTAIL.n241 0.155672
R2287 VTAIL.n257 VTAIL.n241 0.155672
R2288 VTAIL.n258 VTAIL.n257 0.155672
R2289 VTAIL.n258 VTAIL.n237 0.155672
R2290 VTAIL.n265 VTAIL.n237 0.155672
R2291 VTAIL.n266 VTAIL.n265 0.155672
R2292 VTAIL.n266 VTAIL.n233 0.155672
R2293 VTAIL.n273 VTAIL.n233 0.155672
R2294 VTAIL.n274 VTAIL.n273 0.155672
R2295 VTAIL.n274 VTAIL.n229 0.155672
R2296 VTAIL.n281 VTAIL.n229 0.155672
R2297 VTAIL.n282 VTAIL.n281 0.155672
R2298 VTAIL.n282 VTAIL.n225 0.155672
R2299 VTAIL.n290 VTAIL.n225 0.155672
R2300 VTAIL.n291 VTAIL.n290 0.155672
R2301 VTAIL.n291 VTAIL.n221 0.155672
R2302 VTAIL.n299 VTAIL.n221 0.155672
R2303 VTAIL.n300 VTAIL.n299 0.155672
R2304 VTAIL.n300 VTAIL.n217 0.155672
R2305 VTAIL.n307 VTAIL.n217 0.155672
R2306 VTAIL.n308 VTAIL.n307 0.155672
R2307 VTAIL.n308 VTAIL.n213 0.155672
R2308 VTAIL.n315 VTAIL.n213 0.155672
R2309 VTAIL.n739 VTAIL.n637 0.155672
R2310 VTAIL.n732 VTAIL.n637 0.155672
R2311 VTAIL.n732 VTAIL.n731 0.155672
R2312 VTAIL.n731 VTAIL.n641 0.155672
R2313 VTAIL.n724 VTAIL.n641 0.155672
R2314 VTAIL.n724 VTAIL.n723 0.155672
R2315 VTAIL.n723 VTAIL.n645 0.155672
R2316 VTAIL.n715 VTAIL.n645 0.155672
R2317 VTAIL.n715 VTAIL.n714 0.155672
R2318 VTAIL.n714 VTAIL.n649 0.155672
R2319 VTAIL.n707 VTAIL.n649 0.155672
R2320 VTAIL.n707 VTAIL.n706 0.155672
R2321 VTAIL.n706 VTAIL.n654 0.155672
R2322 VTAIL.n699 VTAIL.n654 0.155672
R2323 VTAIL.n699 VTAIL.n698 0.155672
R2324 VTAIL.n698 VTAIL.n658 0.155672
R2325 VTAIL.n691 VTAIL.n658 0.155672
R2326 VTAIL.n691 VTAIL.n690 0.155672
R2327 VTAIL.n690 VTAIL.n662 0.155672
R2328 VTAIL.n683 VTAIL.n662 0.155672
R2329 VTAIL.n683 VTAIL.n682 0.155672
R2330 VTAIL.n682 VTAIL.n666 0.155672
R2331 VTAIL.n675 VTAIL.n666 0.155672
R2332 VTAIL.n675 VTAIL.n674 0.155672
R2333 VTAIL.n633 VTAIL.n531 0.155672
R2334 VTAIL.n626 VTAIL.n531 0.155672
R2335 VTAIL.n626 VTAIL.n625 0.155672
R2336 VTAIL.n625 VTAIL.n535 0.155672
R2337 VTAIL.n618 VTAIL.n535 0.155672
R2338 VTAIL.n618 VTAIL.n617 0.155672
R2339 VTAIL.n617 VTAIL.n539 0.155672
R2340 VTAIL.n609 VTAIL.n539 0.155672
R2341 VTAIL.n609 VTAIL.n608 0.155672
R2342 VTAIL.n608 VTAIL.n543 0.155672
R2343 VTAIL.n601 VTAIL.n543 0.155672
R2344 VTAIL.n601 VTAIL.n600 0.155672
R2345 VTAIL.n600 VTAIL.n548 0.155672
R2346 VTAIL.n593 VTAIL.n548 0.155672
R2347 VTAIL.n593 VTAIL.n592 0.155672
R2348 VTAIL.n592 VTAIL.n552 0.155672
R2349 VTAIL.n585 VTAIL.n552 0.155672
R2350 VTAIL.n585 VTAIL.n584 0.155672
R2351 VTAIL.n584 VTAIL.n556 0.155672
R2352 VTAIL.n577 VTAIL.n556 0.155672
R2353 VTAIL.n577 VTAIL.n576 0.155672
R2354 VTAIL.n576 VTAIL.n560 0.155672
R2355 VTAIL.n569 VTAIL.n560 0.155672
R2356 VTAIL.n569 VTAIL.n568 0.155672
R2357 VTAIL.n527 VTAIL.n425 0.155672
R2358 VTAIL.n520 VTAIL.n425 0.155672
R2359 VTAIL.n520 VTAIL.n519 0.155672
R2360 VTAIL.n519 VTAIL.n429 0.155672
R2361 VTAIL.n512 VTAIL.n429 0.155672
R2362 VTAIL.n512 VTAIL.n511 0.155672
R2363 VTAIL.n511 VTAIL.n433 0.155672
R2364 VTAIL.n503 VTAIL.n433 0.155672
R2365 VTAIL.n503 VTAIL.n502 0.155672
R2366 VTAIL.n502 VTAIL.n437 0.155672
R2367 VTAIL.n495 VTAIL.n437 0.155672
R2368 VTAIL.n495 VTAIL.n494 0.155672
R2369 VTAIL.n494 VTAIL.n442 0.155672
R2370 VTAIL.n487 VTAIL.n442 0.155672
R2371 VTAIL.n487 VTAIL.n486 0.155672
R2372 VTAIL.n486 VTAIL.n446 0.155672
R2373 VTAIL.n479 VTAIL.n446 0.155672
R2374 VTAIL.n479 VTAIL.n478 0.155672
R2375 VTAIL.n478 VTAIL.n450 0.155672
R2376 VTAIL.n471 VTAIL.n450 0.155672
R2377 VTAIL.n471 VTAIL.n470 0.155672
R2378 VTAIL.n470 VTAIL.n454 0.155672
R2379 VTAIL.n463 VTAIL.n454 0.155672
R2380 VTAIL.n463 VTAIL.n462 0.155672
R2381 VTAIL.n421 VTAIL.n319 0.155672
R2382 VTAIL.n414 VTAIL.n319 0.155672
R2383 VTAIL.n414 VTAIL.n413 0.155672
R2384 VTAIL.n413 VTAIL.n323 0.155672
R2385 VTAIL.n406 VTAIL.n323 0.155672
R2386 VTAIL.n406 VTAIL.n405 0.155672
R2387 VTAIL.n405 VTAIL.n327 0.155672
R2388 VTAIL.n397 VTAIL.n327 0.155672
R2389 VTAIL.n397 VTAIL.n396 0.155672
R2390 VTAIL.n396 VTAIL.n331 0.155672
R2391 VTAIL.n389 VTAIL.n331 0.155672
R2392 VTAIL.n389 VTAIL.n388 0.155672
R2393 VTAIL.n388 VTAIL.n336 0.155672
R2394 VTAIL.n381 VTAIL.n336 0.155672
R2395 VTAIL.n381 VTAIL.n380 0.155672
R2396 VTAIL.n380 VTAIL.n340 0.155672
R2397 VTAIL.n373 VTAIL.n340 0.155672
R2398 VTAIL.n373 VTAIL.n372 0.155672
R2399 VTAIL.n372 VTAIL.n344 0.155672
R2400 VTAIL.n365 VTAIL.n344 0.155672
R2401 VTAIL.n365 VTAIL.n364 0.155672
R2402 VTAIL.n364 VTAIL.n348 0.155672
R2403 VTAIL.n357 VTAIL.n348 0.155672
R2404 VTAIL.n357 VTAIL.n356 0.155672
R2405 VP.n2 VP.t0 376.8
R2406 VP.n2 VP.t2 376.57
R2407 VP.n3 VP.t3 338.651
R2408 VP.n9 VP.t1 338.651
R2409 VP.n4 VP.n3 169.13
R2410 VP.n10 VP.n9 169.13
R2411 VP.n8 VP.n0 161.3
R2412 VP.n7 VP.n6 161.3
R2413 VP.n5 VP.n1 161.3
R2414 VP.n4 VP.n2 65.4621
R2415 VP.n7 VP.n1 40.4934
R2416 VP.n8 VP.n7 40.4934
R2417 VP.n3 VP.n1 16.6381
R2418 VP.n9 VP.n8 16.6381
R2419 VP.n5 VP.n4 0.189894
R2420 VP.n6 VP.n5 0.189894
R2421 VP.n6 VP.n0 0.189894
R2422 VP.n10 VP.n0 0.189894
R2423 VP VP.n10 0.0516364
R2424 VDD1 VDD1.n1 113.516
R2425 VDD1 VDD1.n0 68.6369
R2426 VDD1.n0 VDD1.t3 1.714
R2427 VDD1.n0 VDD1.t1 1.714
R2428 VDD1.n1 VDD1.t0 1.714
R2429 VDD1.n1 VDD1.t2 1.714
C0 VDD2 VN 6.24534f
C1 VN VTAIL 5.66859f
C2 w_n1978_n4762# B 9.66164f
C3 B VP 1.36408f
C4 w_n1978_n4762# VP 3.49669f
C5 VDD1 B 1.22923f
C6 VDD1 w_n1978_n4762# 1.38854f
C7 VDD2 B 1.261f
C8 VDD1 VP 6.41182f
C9 VTAIL B 6.3436f
C10 VDD2 w_n1978_n4762# 1.41686f
C11 VDD2 VP 0.314581f
C12 w_n1978_n4762# VTAIL 5.71231f
C13 VTAIL VP 5.6827f
C14 VN B 0.953175f
C15 w_n1978_n4762# VN 3.24557f
C16 VN VP 6.57852f
C17 VDD1 VDD2 0.720845f
C18 VDD1 VTAIL 7.84203f
C19 VDD2 VTAIL 7.88785f
C20 VDD1 VN 0.147685f
C21 VDD2 VSUBS 0.928891f
C22 VDD1 VSUBS 6.02849f
C23 VTAIL VSUBS 1.316429f
C24 VN VSUBS 5.68113f
C25 VP VSUBS 1.882033f
C26 B VSUBS 3.776929f
C27 w_n1978_n4762# VSUBS 0.115096p
C28 VDD1.t3 VSUBS 0.399825f
C29 VDD1.t1 VSUBS 0.399825f
C30 VDD1.n0 VSUBS 3.34281f
C31 VDD1.t0 VSUBS 0.399825f
C32 VDD1.t2 VSUBS 0.399825f
C33 VDD1.n1 VSUBS 4.29645f
C34 VP.n0 VSUBS 0.043571f
C35 VP.t1 VSUBS 3.07217f
C36 VP.n1 VSUBS 0.073768f
C37 VP.t0 VSUBS 3.19778f
C38 VP.t2 VSUBS 3.197f
C39 VP.n2 VSUBS 4.03887f
C40 VP.t3 VSUBS 3.07217f
C41 VP.n3 VSUBS 1.17444f
C42 VP.n4 VSUBS 2.89739f
C43 VP.n5 VSUBS 0.043571f
C44 VP.n6 VSUBS 0.043571f
C45 VP.n7 VSUBS 0.035223f
C46 VP.n8 VSUBS 0.073768f
C47 VP.n9 VSUBS 1.17444f
C48 VP.n10 VSUBS 0.038231f
C49 VTAIL.n0 VSUBS 0.024173f
C50 VTAIL.n1 VSUBS 0.021664f
C51 VTAIL.n2 VSUBS 0.011641f
C52 VTAIL.n3 VSUBS 0.027516f
C53 VTAIL.n4 VSUBS 0.012326f
C54 VTAIL.n5 VSUBS 0.021664f
C55 VTAIL.n6 VSUBS 0.011641f
C56 VTAIL.n7 VSUBS 0.027516f
C57 VTAIL.n8 VSUBS 0.012326f
C58 VTAIL.n9 VSUBS 0.021664f
C59 VTAIL.n10 VSUBS 0.011641f
C60 VTAIL.n11 VSUBS 0.027516f
C61 VTAIL.n12 VSUBS 0.012326f
C62 VTAIL.n13 VSUBS 0.021664f
C63 VTAIL.n14 VSUBS 0.011641f
C64 VTAIL.n15 VSUBS 0.027516f
C65 VTAIL.n16 VSUBS 0.012326f
C66 VTAIL.n17 VSUBS 0.021664f
C67 VTAIL.n18 VSUBS 0.011641f
C68 VTAIL.n19 VSUBS 0.027516f
C69 VTAIL.n20 VSUBS 0.012326f
C70 VTAIL.n21 VSUBS 0.021664f
C71 VTAIL.n22 VSUBS 0.011641f
C72 VTAIL.n23 VSUBS 0.027516f
C73 VTAIL.n24 VSUBS 0.012326f
C74 VTAIL.n25 VSUBS 0.021664f
C75 VTAIL.n26 VSUBS 0.011641f
C76 VTAIL.n27 VSUBS 0.027516f
C77 VTAIL.n28 VSUBS 0.012326f
C78 VTAIL.n29 VSUBS 0.021664f
C79 VTAIL.n30 VSUBS 0.011641f
C80 VTAIL.n31 VSUBS 0.027516f
C81 VTAIL.n32 VSUBS 0.012326f
C82 VTAIL.n33 VSUBS 0.178082f
C83 VTAIL.t7 VSUBS 0.05912f
C84 VTAIL.n34 VSUBS 0.020637f
C85 VTAIL.n35 VSUBS 0.017504f
C86 VTAIL.n36 VSUBS 0.011641f
C87 VTAIL.n37 VSUBS 1.77374f
C88 VTAIL.n38 VSUBS 0.021664f
C89 VTAIL.n39 VSUBS 0.011641f
C90 VTAIL.n40 VSUBS 0.012326f
C91 VTAIL.n41 VSUBS 0.027516f
C92 VTAIL.n42 VSUBS 0.027516f
C93 VTAIL.n43 VSUBS 0.012326f
C94 VTAIL.n44 VSUBS 0.011641f
C95 VTAIL.n45 VSUBS 0.021664f
C96 VTAIL.n46 VSUBS 0.021664f
C97 VTAIL.n47 VSUBS 0.011641f
C98 VTAIL.n48 VSUBS 0.012326f
C99 VTAIL.n49 VSUBS 0.027516f
C100 VTAIL.n50 VSUBS 0.027516f
C101 VTAIL.n51 VSUBS 0.012326f
C102 VTAIL.n52 VSUBS 0.011641f
C103 VTAIL.n53 VSUBS 0.021664f
C104 VTAIL.n54 VSUBS 0.021664f
C105 VTAIL.n55 VSUBS 0.011641f
C106 VTAIL.n56 VSUBS 0.012326f
C107 VTAIL.n57 VSUBS 0.027516f
C108 VTAIL.n58 VSUBS 0.027516f
C109 VTAIL.n59 VSUBS 0.012326f
C110 VTAIL.n60 VSUBS 0.011641f
C111 VTAIL.n61 VSUBS 0.021664f
C112 VTAIL.n62 VSUBS 0.021664f
C113 VTAIL.n63 VSUBS 0.011641f
C114 VTAIL.n64 VSUBS 0.012326f
C115 VTAIL.n65 VSUBS 0.027516f
C116 VTAIL.n66 VSUBS 0.027516f
C117 VTAIL.n67 VSUBS 0.012326f
C118 VTAIL.n68 VSUBS 0.011641f
C119 VTAIL.n69 VSUBS 0.021664f
C120 VTAIL.n70 VSUBS 0.021664f
C121 VTAIL.n71 VSUBS 0.011641f
C122 VTAIL.n72 VSUBS 0.012326f
C123 VTAIL.n73 VSUBS 0.027516f
C124 VTAIL.n74 VSUBS 0.027516f
C125 VTAIL.n75 VSUBS 0.027516f
C126 VTAIL.n76 VSUBS 0.012326f
C127 VTAIL.n77 VSUBS 0.011641f
C128 VTAIL.n78 VSUBS 0.021664f
C129 VTAIL.n79 VSUBS 0.021664f
C130 VTAIL.n80 VSUBS 0.011641f
C131 VTAIL.n81 VSUBS 0.011984f
C132 VTAIL.n82 VSUBS 0.011984f
C133 VTAIL.n83 VSUBS 0.027516f
C134 VTAIL.n84 VSUBS 0.027516f
C135 VTAIL.n85 VSUBS 0.012326f
C136 VTAIL.n86 VSUBS 0.011641f
C137 VTAIL.n87 VSUBS 0.021664f
C138 VTAIL.n88 VSUBS 0.021664f
C139 VTAIL.n89 VSUBS 0.011641f
C140 VTAIL.n90 VSUBS 0.012326f
C141 VTAIL.n91 VSUBS 0.027516f
C142 VTAIL.n92 VSUBS 0.027516f
C143 VTAIL.n93 VSUBS 0.012326f
C144 VTAIL.n94 VSUBS 0.011641f
C145 VTAIL.n95 VSUBS 0.021664f
C146 VTAIL.n96 VSUBS 0.021664f
C147 VTAIL.n97 VSUBS 0.011641f
C148 VTAIL.n98 VSUBS 0.012326f
C149 VTAIL.n99 VSUBS 0.027516f
C150 VTAIL.n100 VSUBS 0.067869f
C151 VTAIL.n101 VSUBS 0.012326f
C152 VTAIL.n102 VSUBS 0.011641f
C153 VTAIL.n103 VSUBS 0.050371f
C154 VTAIL.n104 VSUBS 0.034195f
C155 VTAIL.n105 VSUBS 0.106078f
C156 VTAIL.n106 VSUBS 0.024173f
C157 VTAIL.n107 VSUBS 0.021664f
C158 VTAIL.n108 VSUBS 0.011641f
C159 VTAIL.n109 VSUBS 0.027516f
C160 VTAIL.n110 VSUBS 0.012326f
C161 VTAIL.n111 VSUBS 0.021664f
C162 VTAIL.n112 VSUBS 0.011641f
C163 VTAIL.n113 VSUBS 0.027516f
C164 VTAIL.n114 VSUBS 0.012326f
C165 VTAIL.n115 VSUBS 0.021664f
C166 VTAIL.n116 VSUBS 0.011641f
C167 VTAIL.n117 VSUBS 0.027516f
C168 VTAIL.n118 VSUBS 0.012326f
C169 VTAIL.n119 VSUBS 0.021664f
C170 VTAIL.n120 VSUBS 0.011641f
C171 VTAIL.n121 VSUBS 0.027516f
C172 VTAIL.n122 VSUBS 0.012326f
C173 VTAIL.n123 VSUBS 0.021664f
C174 VTAIL.n124 VSUBS 0.011641f
C175 VTAIL.n125 VSUBS 0.027516f
C176 VTAIL.n126 VSUBS 0.012326f
C177 VTAIL.n127 VSUBS 0.021664f
C178 VTAIL.n128 VSUBS 0.011641f
C179 VTAIL.n129 VSUBS 0.027516f
C180 VTAIL.n130 VSUBS 0.012326f
C181 VTAIL.n131 VSUBS 0.021664f
C182 VTAIL.n132 VSUBS 0.011641f
C183 VTAIL.n133 VSUBS 0.027516f
C184 VTAIL.n134 VSUBS 0.012326f
C185 VTAIL.n135 VSUBS 0.021664f
C186 VTAIL.n136 VSUBS 0.011641f
C187 VTAIL.n137 VSUBS 0.027516f
C188 VTAIL.n138 VSUBS 0.012326f
C189 VTAIL.n139 VSUBS 0.178082f
C190 VTAIL.t2 VSUBS 0.05912f
C191 VTAIL.n140 VSUBS 0.020637f
C192 VTAIL.n141 VSUBS 0.017504f
C193 VTAIL.n142 VSUBS 0.011641f
C194 VTAIL.n143 VSUBS 1.77374f
C195 VTAIL.n144 VSUBS 0.021664f
C196 VTAIL.n145 VSUBS 0.011641f
C197 VTAIL.n146 VSUBS 0.012326f
C198 VTAIL.n147 VSUBS 0.027516f
C199 VTAIL.n148 VSUBS 0.027516f
C200 VTAIL.n149 VSUBS 0.012326f
C201 VTAIL.n150 VSUBS 0.011641f
C202 VTAIL.n151 VSUBS 0.021664f
C203 VTAIL.n152 VSUBS 0.021664f
C204 VTAIL.n153 VSUBS 0.011641f
C205 VTAIL.n154 VSUBS 0.012326f
C206 VTAIL.n155 VSUBS 0.027516f
C207 VTAIL.n156 VSUBS 0.027516f
C208 VTAIL.n157 VSUBS 0.012326f
C209 VTAIL.n158 VSUBS 0.011641f
C210 VTAIL.n159 VSUBS 0.021664f
C211 VTAIL.n160 VSUBS 0.021664f
C212 VTAIL.n161 VSUBS 0.011641f
C213 VTAIL.n162 VSUBS 0.012326f
C214 VTAIL.n163 VSUBS 0.027516f
C215 VTAIL.n164 VSUBS 0.027516f
C216 VTAIL.n165 VSUBS 0.012326f
C217 VTAIL.n166 VSUBS 0.011641f
C218 VTAIL.n167 VSUBS 0.021664f
C219 VTAIL.n168 VSUBS 0.021664f
C220 VTAIL.n169 VSUBS 0.011641f
C221 VTAIL.n170 VSUBS 0.012326f
C222 VTAIL.n171 VSUBS 0.027516f
C223 VTAIL.n172 VSUBS 0.027516f
C224 VTAIL.n173 VSUBS 0.012326f
C225 VTAIL.n174 VSUBS 0.011641f
C226 VTAIL.n175 VSUBS 0.021664f
C227 VTAIL.n176 VSUBS 0.021664f
C228 VTAIL.n177 VSUBS 0.011641f
C229 VTAIL.n178 VSUBS 0.012326f
C230 VTAIL.n179 VSUBS 0.027516f
C231 VTAIL.n180 VSUBS 0.027516f
C232 VTAIL.n181 VSUBS 0.027516f
C233 VTAIL.n182 VSUBS 0.012326f
C234 VTAIL.n183 VSUBS 0.011641f
C235 VTAIL.n184 VSUBS 0.021664f
C236 VTAIL.n185 VSUBS 0.021664f
C237 VTAIL.n186 VSUBS 0.011641f
C238 VTAIL.n187 VSUBS 0.011984f
C239 VTAIL.n188 VSUBS 0.011984f
C240 VTAIL.n189 VSUBS 0.027516f
C241 VTAIL.n190 VSUBS 0.027516f
C242 VTAIL.n191 VSUBS 0.012326f
C243 VTAIL.n192 VSUBS 0.011641f
C244 VTAIL.n193 VSUBS 0.021664f
C245 VTAIL.n194 VSUBS 0.021664f
C246 VTAIL.n195 VSUBS 0.011641f
C247 VTAIL.n196 VSUBS 0.012326f
C248 VTAIL.n197 VSUBS 0.027516f
C249 VTAIL.n198 VSUBS 0.027516f
C250 VTAIL.n199 VSUBS 0.012326f
C251 VTAIL.n200 VSUBS 0.011641f
C252 VTAIL.n201 VSUBS 0.021664f
C253 VTAIL.n202 VSUBS 0.021664f
C254 VTAIL.n203 VSUBS 0.011641f
C255 VTAIL.n204 VSUBS 0.012326f
C256 VTAIL.n205 VSUBS 0.027516f
C257 VTAIL.n206 VSUBS 0.067869f
C258 VTAIL.n207 VSUBS 0.012326f
C259 VTAIL.n208 VSUBS 0.011641f
C260 VTAIL.n209 VSUBS 0.050371f
C261 VTAIL.n210 VSUBS 0.034195f
C262 VTAIL.n211 VSUBS 0.152566f
C263 VTAIL.n212 VSUBS 0.024173f
C264 VTAIL.n213 VSUBS 0.021664f
C265 VTAIL.n214 VSUBS 0.011641f
C266 VTAIL.n215 VSUBS 0.027516f
C267 VTAIL.n216 VSUBS 0.012326f
C268 VTAIL.n217 VSUBS 0.021664f
C269 VTAIL.n218 VSUBS 0.011641f
C270 VTAIL.n219 VSUBS 0.027516f
C271 VTAIL.n220 VSUBS 0.012326f
C272 VTAIL.n221 VSUBS 0.021664f
C273 VTAIL.n222 VSUBS 0.011641f
C274 VTAIL.n223 VSUBS 0.027516f
C275 VTAIL.n224 VSUBS 0.012326f
C276 VTAIL.n225 VSUBS 0.021664f
C277 VTAIL.n226 VSUBS 0.011641f
C278 VTAIL.n227 VSUBS 0.027516f
C279 VTAIL.n228 VSUBS 0.012326f
C280 VTAIL.n229 VSUBS 0.021664f
C281 VTAIL.n230 VSUBS 0.011641f
C282 VTAIL.n231 VSUBS 0.027516f
C283 VTAIL.n232 VSUBS 0.012326f
C284 VTAIL.n233 VSUBS 0.021664f
C285 VTAIL.n234 VSUBS 0.011641f
C286 VTAIL.n235 VSUBS 0.027516f
C287 VTAIL.n236 VSUBS 0.012326f
C288 VTAIL.n237 VSUBS 0.021664f
C289 VTAIL.n238 VSUBS 0.011641f
C290 VTAIL.n239 VSUBS 0.027516f
C291 VTAIL.n240 VSUBS 0.012326f
C292 VTAIL.n241 VSUBS 0.021664f
C293 VTAIL.n242 VSUBS 0.011641f
C294 VTAIL.n243 VSUBS 0.027516f
C295 VTAIL.n244 VSUBS 0.012326f
C296 VTAIL.n245 VSUBS 0.178082f
C297 VTAIL.t1 VSUBS 0.05912f
C298 VTAIL.n246 VSUBS 0.020637f
C299 VTAIL.n247 VSUBS 0.017504f
C300 VTAIL.n248 VSUBS 0.011641f
C301 VTAIL.n249 VSUBS 1.77374f
C302 VTAIL.n250 VSUBS 0.021664f
C303 VTAIL.n251 VSUBS 0.011641f
C304 VTAIL.n252 VSUBS 0.012326f
C305 VTAIL.n253 VSUBS 0.027516f
C306 VTAIL.n254 VSUBS 0.027516f
C307 VTAIL.n255 VSUBS 0.012326f
C308 VTAIL.n256 VSUBS 0.011641f
C309 VTAIL.n257 VSUBS 0.021664f
C310 VTAIL.n258 VSUBS 0.021664f
C311 VTAIL.n259 VSUBS 0.011641f
C312 VTAIL.n260 VSUBS 0.012326f
C313 VTAIL.n261 VSUBS 0.027516f
C314 VTAIL.n262 VSUBS 0.027516f
C315 VTAIL.n263 VSUBS 0.012326f
C316 VTAIL.n264 VSUBS 0.011641f
C317 VTAIL.n265 VSUBS 0.021664f
C318 VTAIL.n266 VSUBS 0.021664f
C319 VTAIL.n267 VSUBS 0.011641f
C320 VTAIL.n268 VSUBS 0.012326f
C321 VTAIL.n269 VSUBS 0.027516f
C322 VTAIL.n270 VSUBS 0.027516f
C323 VTAIL.n271 VSUBS 0.012326f
C324 VTAIL.n272 VSUBS 0.011641f
C325 VTAIL.n273 VSUBS 0.021664f
C326 VTAIL.n274 VSUBS 0.021664f
C327 VTAIL.n275 VSUBS 0.011641f
C328 VTAIL.n276 VSUBS 0.012326f
C329 VTAIL.n277 VSUBS 0.027516f
C330 VTAIL.n278 VSUBS 0.027516f
C331 VTAIL.n279 VSUBS 0.012326f
C332 VTAIL.n280 VSUBS 0.011641f
C333 VTAIL.n281 VSUBS 0.021664f
C334 VTAIL.n282 VSUBS 0.021664f
C335 VTAIL.n283 VSUBS 0.011641f
C336 VTAIL.n284 VSUBS 0.012326f
C337 VTAIL.n285 VSUBS 0.027516f
C338 VTAIL.n286 VSUBS 0.027516f
C339 VTAIL.n287 VSUBS 0.027516f
C340 VTAIL.n288 VSUBS 0.012326f
C341 VTAIL.n289 VSUBS 0.011641f
C342 VTAIL.n290 VSUBS 0.021664f
C343 VTAIL.n291 VSUBS 0.021664f
C344 VTAIL.n292 VSUBS 0.011641f
C345 VTAIL.n293 VSUBS 0.011984f
C346 VTAIL.n294 VSUBS 0.011984f
C347 VTAIL.n295 VSUBS 0.027516f
C348 VTAIL.n296 VSUBS 0.027516f
C349 VTAIL.n297 VSUBS 0.012326f
C350 VTAIL.n298 VSUBS 0.011641f
C351 VTAIL.n299 VSUBS 0.021664f
C352 VTAIL.n300 VSUBS 0.021664f
C353 VTAIL.n301 VSUBS 0.011641f
C354 VTAIL.n302 VSUBS 0.012326f
C355 VTAIL.n303 VSUBS 0.027516f
C356 VTAIL.n304 VSUBS 0.027516f
C357 VTAIL.n305 VSUBS 0.012326f
C358 VTAIL.n306 VSUBS 0.011641f
C359 VTAIL.n307 VSUBS 0.021664f
C360 VTAIL.n308 VSUBS 0.021664f
C361 VTAIL.n309 VSUBS 0.011641f
C362 VTAIL.n310 VSUBS 0.012326f
C363 VTAIL.n311 VSUBS 0.027516f
C364 VTAIL.n312 VSUBS 0.067869f
C365 VTAIL.n313 VSUBS 0.012326f
C366 VTAIL.n314 VSUBS 0.011641f
C367 VTAIL.n315 VSUBS 0.050371f
C368 VTAIL.n316 VSUBS 0.034195f
C369 VTAIL.n317 VSUBS 1.65673f
C370 VTAIL.n318 VSUBS 0.024173f
C371 VTAIL.n319 VSUBS 0.021664f
C372 VTAIL.n320 VSUBS 0.011641f
C373 VTAIL.n321 VSUBS 0.027516f
C374 VTAIL.n322 VSUBS 0.012326f
C375 VTAIL.n323 VSUBS 0.021664f
C376 VTAIL.n324 VSUBS 0.011641f
C377 VTAIL.n325 VSUBS 0.027516f
C378 VTAIL.n326 VSUBS 0.012326f
C379 VTAIL.n327 VSUBS 0.021664f
C380 VTAIL.n328 VSUBS 0.011641f
C381 VTAIL.n329 VSUBS 0.027516f
C382 VTAIL.n330 VSUBS 0.012326f
C383 VTAIL.n331 VSUBS 0.021664f
C384 VTAIL.n332 VSUBS 0.011641f
C385 VTAIL.n333 VSUBS 0.027516f
C386 VTAIL.n334 VSUBS 0.027516f
C387 VTAIL.n335 VSUBS 0.012326f
C388 VTAIL.n336 VSUBS 0.021664f
C389 VTAIL.n337 VSUBS 0.011641f
C390 VTAIL.n338 VSUBS 0.027516f
C391 VTAIL.n339 VSUBS 0.012326f
C392 VTAIL.n340 VSUBS 0.021664f
C393 VTAIL.n341 VSUBS 0.011641f
C394 VTAIL.n342 VSUBS 0.027516f
C395 VTAIL.n343 VSUBS 0.012326f
C396 VTAIL.n344 VSUBS 0.021664f
C397 VTAIL.n345 VSUBS 0.011641f
C398 VTAIL.n346 VSUBS 0.027516f
C399 VTAIL.n347 VSUBS 0.012326f
C400 VTAIL.n348 VSUBS 0.021664f
C401 VTAIL.n349 VSUBS 0.011641f
C402 VTAIL.n350 VSUBS 0.027516f
C403 VTAIL.n351 VSUBS 0.012326f
C404 VTAIL.n352 VSUBS 0.178082f
C405 VTAIL.t4 VSUBS 0.05912f
C406 VTAIL.n353 VSUBS 0.020637f
C407 VTAIL.n354 VSUBS 0.017504f
C408 VTAIL.n355 VSUBS 0.011641f
C409 VTAIL.n356 VSUBS 1.77374f
C410 VTAIL.n357 VSUBS 0.021664f
C411 VTAIL.n358 VSUBS 0.011641f
C412 VTAIL.n359 VSUBS 0.012326f
C413 VTAIL.n360 VSUBS 0.027516f
C414 VTAIL.n361 VSUBS 0.027516f
C415 VTAIL.n362 VSUBS 0.012326f
C416 VTAIL.n363 VSUBS 0.011641f
C417 VTAIL.n364 VSUBS 0.021664f
C418 VTAIL.n365 VSUBS 0.021664f
C419 VTAIL.n366 VSUBS 0.011641f
C420 VTAIL.n367 VSUBS 0.012326f
C421 VTAIL.n368 VSUBS 0.027516f
C422 VTAIL.n369 VSUBS 0.027516f
C423 VTAIL.n370 VSUBS 0.012326f
C424 VTAIL.n371 VSUBS 0.011641f
C425 VTAIL.n372 VSUBS 0.021664f
C426 VTAIL.n373 VSUBS 0.021664f
C427 VTAIL.n374 VSUBS 0.011641f
C428 VTAIL.n375 VSUBS 0.012326f
C429 VTAIL.n376 VSUBS 0.027516f
C430 VTAIL.n377 VSUBS 0.027516f
C431 VTAIL.n378 VSUBS 0.012326f
C432 VTAIL.n379 VSUBS 0.011641f
C433 VTAIL.n380 VSUBS 0.021664f
C434 VTAIL.n381 VSUBS 0.021664f
C435 VTAIL.n382 VSUBS 0.011641f
C436 VTAIL.n383 VSUBS 0.012326f
C437 VTAIL.n384 VSUBS 0.027516f
C438 VTAIL.n385 VSUBS 0.027516f
C439 VTAIL.n386 VSUBS 0.012326f
C440 VTAIL.n387 VSUBS 0.011641f
C441 VTAIL.n388 VSUBS 0.021664f
C442 VTAIL.n389 VSUBS 0.021664f
C443 VTAIL.n390 VSUBS 0.011641f
C444 VTAIL.n391 VSUBS 0.012326f
C445 VTAIL.n392 VSUBS 0.027516f
C446 VTAIL.n393 VSUBS 0.027516f
C447 VTAIL.n394 VSUBS 0.012326f
C448 VTAIL.n395 VSUBS 0.011641f
C449 VTAIL.n396 VSUBS 0.021664f
C450 VTAIL.n397 VSUBS 0.021664f
C451 VTAIL.n398 VSUBS 0.011641f
C452 VTAIL.n399 VSUBS 0.011984f
C453 VTAIL.n400 VSUBS 0.011984f
C454 VTAIL.n401 VSUBS 0.027516f
C455 VTAIL.n402 VSUBS 0.027516f
C456 VTAIL.n403 VSUBS 0.012326f
C457 VTAIL.n404 VSUBS 0.011641f
C458 VTAIL.n405 VSUBS 0.021664f
C459 VTAIL.n406 VSUBS 0.021664f
C460 VTAIL.n407 VSUBS 0.011641f
C461 VTAIL.n408 VSUBS 0.012326f
C462 VTAIL.n409 VSUBS 0.027516f
C463 VTAIL.n410 VSUBS 0.027516f
C464 VTAIL.n411 VSUBS 0.012326f
C465 VTAIL.n412 VSUBS 0.011641f
C466 VTAIL.n413 VSUBS 0.021664f
C467 VTAIL.n414 VSUBS 0.021664f
C468 VTAIL.n415 VSUBS 0.011641f
C469 VTAIL.n416 VSUBS 0.012326f
C470 VTAIL.n417 VSUBS 0.027516f
C471 VTAIL.n418 VSUBS 0.067869f
C472 VTAIL.n419 VSUBS 0.012326f
C473 VTAIL.n420 VSUBS 0.011641f
C474 VTAIL.n421 VSUBS 0.050371f
C475 VTAIL.n422 VSUBS 0.034195f
C476 VTAIL.n423 VSUBS 1.65673f
C477 VTAIL.n424 VSUBS 0.024173f
C478 VTAIL.n425 VSUBS 0.021664f
C479 VTAIL.n426 VSUBS 0.011641f
C480 VTAIL.n427 VSUBS 0.027516f
C481 VTAIL.n428 VSUBS 0.012326f
C482 VTAIL.n429 VSUBS 0.021664f
C483 VTAIL.n430 VSUBS 0.011641f
C484 VTAIL.n431 VSUBS 0.027516f
C485 VTAIL.n432 VSUBS 0.012326f
C486 VTAIL.n433 VSUBS 0.021664f
C487 VTAIL.n434 VSUBS 0.011641f
C488 VTAIL.n435 VSUBS 0.027516f
C489 VTAIL.n436 VSUBS 0.012326f
C490 VTAIL.n437 VSUBS 0.021664f
C491 VTAIL.n438 VSUBS 0.011641f
C492 VTAIL.n439 VSUBS 0.027516f
C493 VTAIL.n440 VSUBS 0.027516f
C494 VTAIL.n441 VSUBS 0.012326f
C495 VTAIL.n442 VSUBS 0.021664f
C496 VTAIL.n443 VSUBS 0.011641f
C497 VTAIL.n444 VSUBS 0.027516f
C498 VTAIL.n445 VSUBS 0.012326f
C499 VTAIL.n446 VSUBS 0.021664f
C500 VTAIL.n447 VSUBS 0.011641f
C501 VTAIL.n448 VSUBS 0.027516f
C502 VTAIL.n449 VSUBS 0.012326f
C503 VTAIL.n450 VSUBS 0.021664f
C504 VTAIL.n451 VSUBS 0.011641f
C505 VTAIL.n452 VSUBS 0.027516f
C506 VTAIL.n453 VSUBS 0.012326f
C507 VTAIL.n454 VSUBS 0.021664f
C508 VTAIL.n455 VSUBS 0.011641f
C509 VTAIL.n456 VSUBS 0.027516f
C510 VTAIL.n457 VSUBS 0.012326f
C511 VTAIL.n458 VSUBS 0.178082f
C512 VTAIL.t5 VSUBS 0.05912f
C513 VTAIL.n459 VSUBS 0.020637f
C514 VTAIL.n460 VSUBS 0.017504f
C515 VTAIL.n461 VSUBS 0.011641f
C516 VTAIL.n462 VSUBS 1.77374f
C517 VTAIL.n463 VSUBS 0.021664f
C518 VTAIL.n464 VSUBS 0.011641f
C519 VTAIL.n465 VSUBS 0.012326f
C520 VTAIL.n466 VSUBS 0.027516f
C521 VTAIL.n467 VSUBS 0.027516f
C522 VTAIL.n468 VSUBS 0.012326f
C523 VTAIL.n469 VSUBS 0.011641f
C524 VTAIL.n470 VSUBS 0.021664f
C525 VTAIL.n471 VSUBS 0.021664f
C526 VTAIL.n472 VSUBS 0.011641f
C527 VTAIL.n473 VSUBS 0.012326f
C528 VTAIL.n474 VSUBS 0.027516f
C529 VTAIL.n475 VSUBS 0.027516f
C530 VTAIL.n476 VSUBS 0.012326f
C531 VTAIL.n477 VSUBS 0.011641f
C532 VTAIL.n478 VSUBS 0.021664f
C533 VTAIL.n479 VSUBS 0.021664f
C534 VTAIL.n480 VSUBS 0.011641f
C535 VTAIL.n481 VSUBS 0.012326f
C536 VTAIL.n482 VSUBS 0.027516f
C537 VTAIL.n483 VSUBS 0.027516f
C538 VTAIL.n484 VSUBS 0.012326f
C539 VTAIL.n485 VSUBS 0.011641f
C540 VTAIL.n486 VSUBS 0.021664f
C541 VTAIL.n487 VSUBS 0.021664f
C542 VTAIL.n488 VSUBS 0.011641f
C543 VTAIL.n489 VSUBS 0.012326f
C544 VTAIL.n490 VSUBS 0.027516f
C545 VTAIL.n491 VSUBS 0.027516f
C546 VTAIL.n492 VSUBS 0.012326f
C547 VTAIL.n493 VSUBS 0.011641f
C548 VTAIL.n494 VSUBS 0.021664f
C549 VTAIL.n495 VSUBS 0.021664f
C550 VTAIL.n496 VSUBS 0.011641f
C551 VTAIL.n497 VSUBS 0.012326f
C552 VTAIL.n498 VSUBS 0.027516f
C553 VTAIL.n499 VSUBS 0.027516f
C554 VTAIL.n500 VSUBS 0.012326f
C555 VTAIL.n501 VSUBS 0.011641f
C556 VTAIL.n502 VSUBS 0.021664f
C557 VTAIL.n503 VSUBS 0.021664f
C558 VTAIL.n504 VSUBS 0.011641f
C559 VTAIL.n505 VSUBS 0.011984f
C560 VTAIL.n506 VSUBS 0.011984f
C561 VTAIL.n507 VSUBS 0.027516f
C562 VTAIL.n508 VSUBS 0.027516f
C563 VTAIL.n509 VSUBS 0.012326f
C564 VTAIL.n510 VSUBS 0.011641f
C565 VTAIL.n511 VSUBS 0.021664f
C566 VTAIL.n512 VSUBS 0.021664f
C567 VTAIL.n513 VSUBS 0.011641f
C568 VTAIL.n514 VSUBS 0.012326f
C569 VTAIL.n515 VSUBS 0.027516f
C570 VTAIL.n516 VSUBS 0.027516f
C571 VTAIL.n517 VSUBS 0.012326f
C572 VTAIL.n518 VSUBS 0.011641f
C573 VTAIL.n519 VSUBS 0.021664f
C574 VTAIL.n520 VSUBS 0.021664f
C575 VTAIL.n521 VSUBS 0.011641f
C576 VTAIL.n522 VSUBS 0.012326f
C577 VTAIL.n523 VSUBS 0.027516f
C578 VTAIL.n524 VSUBS 0.067869f
C579 VTAIL.n525 VSUBS 0.012326f
C580 VTAIL.n526 VSUBS 0.011641f
C581 VTAIL.n527 VSUBS 0.050371f
C582 VTAIL.n528 VSUBS 0.034195f
C583 VTAIL.n529 VSUBS 0.152566f
C584 VTAIL.n530 VSUBS 0.024173f
C585 VTAIL.n531 VSUBS 0.021664f
C586 VTAIL.n532 VSUBS 0.011641f
C587 VTAIL.n533 VSUBS 0.027516f
C588 VTAIL.n534 VSUBS 0.012326f
C589 VTAIL.n535 VSUBS 0.021664f
C590 VTAIL.n536 VSUBS 0.011641f
C591 VTAIL.n537 VSUBS 0.027516f
C592 VTAIL.n538 VSUBS 0.012326f
C593 VTAIL.n539 VSUBS 0.021664f
C594 VTAIL.n540 VSUBS 0.011641f
C595 VTAIL.n541 VSUBS 0.027516f
C596 VTAIL.n542 VSUBS 0.012326f
C597 VTAIL.n543 VSUBS 0.021664f
C598 VTAIL.n544 VSUBS 0.011641f
C599 VTAIL.n545 VSUBS 0.027516f
C600 VTAIL.n546 VSUBS 0.027516f
C601 VTAIL.n547 VSUBS 0.012326f
C602 VTAIL.n548 VSUBS 0.021664f
C603 VTAIL.n549 VSUBS 0.011641f
C604 VTAIL.n550 VSUBS 0.027516f
C605 VTAIL.n551 VSUBS 0.012326f
C606 VTAIL.n552 VSUBS 0.021664f
C607 VTAIL.n553 VSUBS 0.011641f
C608 VTAIL.n554 VSUBS 0.027516f
C609 VTAIL.n555 VSUBS 0.012326f
C610 VTAIL.n556 VSUBS 0.021664f
C611 VTAIL.n557 VSUBS 0.011641f
C612 VTAIL.n558 VSUBS 0.027516f
C613 VTAIL.n559 VSUBS 0.012326f
C614 VTAIL.n560 VSUBS 0.021664f
C615 VTAIL.n561 VSUBS 0.011641f
C616 VTAIL.n562 VSUBS 0.027516f
C617 VTAIL.n563 VSUBS 0.012326f
C618 VTAIL.n564 VSUBS 0.178082f
C619 VTAIL.t0 VSUBS 0.05912f
C620 VTAIL.n565 VSUBS 0.020637f
C621 VTAIL.n566 VSUBS 0.017504f
C622 VTAIL.n567 VSUBS 0.011641f
C623 VTAIL.n568 VSUBS 1.77374f
C624 VTAIL.n569 VSUBS 0.021664f
C625 VTAIL.n570 VSUBS 0.011641f
C626 VTAIL.n571 VSUBS 0.012326f
C627 VTAIL.n572 VSUBS 0.027516f
C628 VTAIL.n573 VSUBS 0.027516f
C629 VTAIL.n574 VSUBS 0.012326f
C630 VTAIL.n575 VSUBS 0.011641f
C631 VTAIL.n576 VSUBS 0.021664f
C632 VTAIL.n577 VSUBS 0.021664f
C633 VTAIL.n578 VSUBS 0.011641f
C634 VTAIL.n579 VSUBS 0.012326f
C635 VTAIL.n580 VSUBS 0.027516f
C636 VTAIL.n581 VSUBS 0.027516f
C637 VTAIL.n582 VSUBS 0.012326f
C638 VTAIL.n583 VSUBS 0.011641f
C639 VTAIL.n584 VSUBS 0.021664f
C640 VTAIL.n585 VSUBS 0.021664f
C641 VTAIL.n586 VSUBS 0.011641f
C642 VTAIL.n587 VSUBS 0.012326f
C643 VTAIL.n588 VSUBS 0.027516f
C644 VTAIL.n589 VSUBS 0.027516f
C645 VTAIL.n590 VSUBS 0.012326f
C646 VTAIL.n591 VSUBS 0.011641f
C647 VTAIL.n592 VSUBS 0.021664f
C648 VTAIL.n593 VSUBS 0.021664f
C649 VTAIL.n594 VSUBS 0.011641f
C650 VTAIL.n595 VSUBS 0.012326f
C651 VTAIL.n596 VSUBS 0.027516f
C652 VTAIL.n597 VSUBS 0.027516f
C653 VTAIL.n598 VSUBS 0.012326f
C654 VTAIL.n599 VSUBS 0.011641f
C655 VTAIL.n600 VSUBS 0.021664f
C656 VTAIL.n601 VSUBS 0.021664f
C657 VTAIL.n602 VSUBS 0.011641f
C658 VTAIL.n603 VSUBS 0.012326f
C659 VTAIL.n604 VSUBS 0.027516f
C660 VTAIL.n605 VSUBS 0.027516f
C661 VTAIL.n606 VSUBS 0.012326f
C662 VTAIL.n607 VSUBS 0.011641f
C663 VTAIL.n608 VSUBS 0.021664f
C664 VTAIL.n609 VSUBS 0.021664f
C665 VTAIL.n610 VSUBS 0.011641f
C666 VTAIL.n611 VSUBS 0.011984f
C667 VTAIL.n612 VSUBS 0.011984f
C668 VTAIL.n613 VSUBS 0.027516f
C669 VTAIL.n614 VSUBS 0.027516f
C670 VTAIL.n615 VSUBS 0.012326f
C671 VTAIL.n616 VSUBS 0.011641f
C672 VTAIL.n617 VSUBS 0.021664f
C673 VTAIL.n618 VSUBS 0.021664f
C674 VTAIL.n619 VSUBS 0.011641f
C675 VTAIL.n620 VSUBS 0.012326f
C676 VTAIL.n621 VSUBS 0.027516f
C677 VTAIL.n622 VSUBS 0.027516f
C678 VTAIL.n623 VSUBS 0.012326f
C679 VTAIL.n624 VSUBS 0.011641f
C680 VTAIL.n625 VSUBS 0.021664f
C681 VTAIL.n626 VSUBS 0.021664f
C682 VTAIL.n627 VSUBS 0.011641f
C683 VTAIL.n628 VSUBS 0.012326f
C684 VTAIL.n629 VSUBS 0.027516f
C685 VTAIL.n630 VSUBS 0.067869f
C686 VTAIL.n631 VSUBS 0.012326f
C687 VTAIL.n632 VSUBS 0.011641f
C688 VTAIL.n633 VSUBS 0.050371f
C689 VTAIL.n634 VSUBS 0.034195f
C690 VTAIL.n635 VSUBS 0.152566f
C691 VTAIL.n636 VSUBS 0.024173f
C692 VTAIL.n637 VSUBS 0.021664f
C693 VTAIL.n638 VSUBS 0.011641f
C694 VTAIL.n639 VSUBS 0.027516f
C695 VTAIL.n640 VSUBS 0.012326f
C696 VTAIL.n641 VSUBS 0.021664f
C697 VTAIL.n642 VSUBS 0.011641f
C698 VTAIL.n643 VSUBS 0.027516f
C699 VTAIL.n644 VSUBS 0.012326f
C700 VTAIL.n645 VSUBS 0.021664f
C701 VTAIL.n646 VSUBS 0.011641f
C702 VTAIL.n647 VSUBS 0.027516f
C703 VTAIL.n648 VSUBS 0.012326f
C704 VTAIL.n649 VSUBS 0.021664f
C705 VTAIL.n650 VSUBS 0.011641f
C706 VTAIL.n651 VSUBS 0.027516f
C707 VTAIL.n652 VSUBS 0.027516f
C708 VTAIL.n653 VSUBS 0.012326f
C709 VTAIL.n654 VSUBS 0.021664f
C710 VTAIL.n655 VSUBS 0.011641f
C711 VTAIL.n656 VSUBS 0.027516f
C712 VTAIL.n657 VSUBS 0.012326f
C713 VTAIL.n658 VSUBS 0.021664f
C714 VTAIL.n659 VSUBS 0.011641f
C715 VTAIL.n660 VSUBS 0.027516f
C716 VTAIL.n661 VSUBS 0.012326f
C717 VTAIL.n662 VSUBS 0.021664f
C718 VTAIL.n663 VSUBS 0.011641f
C719 VTAIL.n664 VSUBS 0.027516f
C720 VTAIL.n665 VSUBS 0.012326f
C721 VTAIL.n666 VSUBS 0.021664f
C722 VTAIL.n667 VSUBS 0.011641f
C723 VTAIL.n668 VSUBS 0.027516f
C724 VTAIL.n669 VSUBS 0.012326f
C725 VTAIL.n670 VSUBS 0.178082f
C726 VTAIL.t3 VSUBS 0.05912f
C727 VTAIL.n671 VSUBS 0.020637f
C728 VTAIL.n672 VSUBS 0.017504f
C729 VTAIL.n673 VSUBS 0.011641f
C730 VTAIL.n674 VSUBS 1.77374f
C731 VTAIL.n675 VSUBS 0.021664f
C732 VTAIL.n676 VSUBS 0.011641f
C733 VTAIL.n677 VSUBS 0.012326f
C734 VTAIL.n678 VSUBS 0.027516f
C735 VTAIL.n679 VSUBS 0.027516f
C736 VTAIL.n680 VSUBS 0.012326f
C737 VTAIL.n681 VSUBS 0.011641f
C738 VTAIL.n682 VSUBS 0.021664f
C739 VTAIL.n683 VSUBS 0.021664f
C740 VTAIL.n684 VSUBS 0.011641f
C741 VTAIL.n685 VSUBS 0.012326f
C742 VTAIL.n686 VSUBS 0.027516f
C743 VTAIL.n687 VSUBS 0.027516f
C744 VTAIL.n688 VSUBS 0.012326f
C745 VTAIL.n689 VSUBS 0.011641f
C746 VTAIL.n690 VSUBS 0.021664f
C747 VTAIL.n691 VSUBS 0.021664f
C748 VTAIL.n692 VSUBS 0.011641f
C749 VTAIL.n693 VSUBS 0.012326f
C750 VTAIL.n694 VSUBS 0.027516f
C751 VTAIL.n695 VSUBS 0.027516f
C752 VTAIL.n696 VSUBS 0.012326f
C753 VTAIL.n697 VSUBS 0.011641f
C754 VTAIL.n698 VSUBS 0.021664f
C755 VTAIL.n699 VSUBS 0.021664f
C756 VTAIL.n700 VSUBS 0.011641f
C757 VTAIL.n701 VSUBS 0.012326f
C758 VTAIL.n702 VSUBS 0.027516f
C759 VTAIL.n703 VSUBS 0.027516f
C760 VTAIL.n704 VSUBS 0.012326f
C761 VTAIL.n705 VSUBS 0.011641f
C762 VTAIL.n706 VSUBS 0.021664f
C763 VTAIL.n707 VSUBS 0.021664f
C764 VTAIL.n708 VSUBS 0.011641f
C765 VTAIL.n709 VSUBS 0.012326f
C766 VTAIL.n710 VSUBS 0.027516f
C767 VTAIL.n711 VSUBS 0.027516f
C768 VTAIL.n712 VSUBS 0.012326f
C769 VTAIL.n713 VSUBS 0.011641f
C770 VTAIL.n714 VSUBS 0.021664f
C771 VTAIL.n715 VSUBS 0.021664f
C772 VTAIL.n716 VSUBS 0.011641f
C773 VTAIL.n717 VSUBS 0.011984f
C774 VTAIL.n718 VSUBS 0.011984f
C775 VTAIL.n719 VSUBS 0.027516f
C776 VTAIL.n720 VSUBS 0.027516f
C777 VTAIL.n721 VSUBS 0.012326f
C778 VTAIL.n722 VSUBS 0.011641f
C779 VTAIL.n723 VSUBS 0.021664f
C780 VTAIL.n724 VSUBS 0.021664f
C781 VTAIL.n725 VSUBS 0.011641f
C782 VTAIL.n726 VSUBS 0.012326f
C783 VTAIL.n727 VSUBS 0.027516f
C784 VTAIL.n728 VSUBS 0.027516f
C785 VTAIL.n729 VSUBS 0.012326f
C786 VTAIL.n730 VSUBS 0.011641f
C787 VTAIL.n731 VSUBS 0.021664f
C788 VTAIL.n732 VSUBS 0.021664f
C789 VTAIL.n733 VSUBS 0.011641f
C790 VTAIL.n734 VSUBS 0.012326f
C791 VTAIL.n735 VSUBS 0.027516f
C792 VTAIL.n736 VSUBS 0.067869f
C793 VTAIL.n737 VSUBS 0.012326f
C794 VTAIL.n738 VSUBS 0.011641f
C795 VTAIL.n739 VSUBS 0.050371f
C796 VTAIL.n740 VSUBS 0.034195f
C797 VTAIL.n741 VSUBS 1.65673f
C798 VTAIL.n742 VSUBS 0.024173f
C799 VTAIL.n743 VSUBS 0.021664f
C800 VTAIL.n744 VSUBS 0.011641f
C801 VTAIL.n745 VSUBS 0.027516f
C802 VTAIL.n746 VSUBS 0.012326f
C803 VTAIL.n747 VSUBS 0.021664f
C804 VTAIL.n748 VSUBS 0.011641f
C805 VTAIL.n749 VSUBS 0.027516f
C806 VTAIL.n750 VSUBS 0.012326f
C807 VTAIL.n751 VSUBS 0.021664f
C808 VTAIL.n752 VSUBS 0.011641f
C809 VTAIL.n753 VSUBS 0.027516f
C810 VTAIL.n754 VSUBS 0.012326f
C811 VTAIL.n755 VSUBS 0.021664f
C812 VTAIL.n756 VSUBS 0.011641f
C813 VTAIL.n757 VSUBS 0.027516f
C814 VTAIL.n758 VSUBS 0.012326f
C815 VTAIL.n759 VSUBS 0.021664f
C816 VTAIL.n760 VSUBS 0.011641f
C817 VTAIL.n761 VSUBS 0.027516f
C818 VTAIL.n762 VSUBS 0.012326f
C819 VTAIL.n763 VSUBS 0.021664f
C820 VTAIL.n764 VSUBS 0.011641f
C821 VTAIL.n765 VSUBS 0.027516f
C822 VTAIL.n766 VSUBS 0.012326f
C823 VTAIL.n767 VSUBS 0.021664f
C824 VTAIL.n768 VSUBS 0.011641f
C825 VTAIL.n769 VSUBS 0.027516f
C826 VTAIL.n770 VSUBS 0.012326f
C827 VTAIL.n771 VSUBS 0.021664f
C828 VTAIL.n772 VSUBS 0.011641f
C829 VTAIL.n773 VSUBS 0.027516f
C830 VTAIL.n774 VSUBS 0.012326f
C831 VTAIL.n775 VSUBS 0.178082f
C832 VTAIL.t6 VSUBS 0.05912f
C833 VTAIL.n776 VSUBS 0.020637f
C834 VTAIL.n777 VSUBS 0.017504f
C835 VTAIL.n778 VSUBS 0.011641f
C836 VTAIL.n779 VSUBS 1.77374f
C837 VTAIL.n780 VSUBS 0.021664f
C838 VTAIL.n781 VSUBS 0.011641f
C839 VTAIL.n782 VSUBS 0.012326f
C840 VTAIL.n783 VSUBS 0.027516f
C841 VTAIL.n784 VSUBS 0.027516f
C842 VTAIL.n785 VSUBS 0.012326f
C843 VTAIL.n786 VSUBS 0.011641f
C844 VTAIL.n787 VSUBS 0.021664f
C845 VTAIL.n788 VSUBS 0.021664f
C846 VTAIL.n789 VSUBS 0.011641f
C847 VTAIL.n790 VSUBS 0.012326f
C848 VTAIL.n791 VSUBS 0.027516f
C849 VTAIL.n792 VSUBS 0.027516f
C850 VTAIL.n793 VSUBS 0.012326f
C851 VTAIL.n794 VSUBS 0.011641f
C852 VTAIL.n795 VSUBS 0.021664f
C853 VTAIL.n796 VSUBS 0.021664f
C854 VTAIL.n797 VSUBS 0.011641f
C855 VTAIL.n798 VSUBS 0.012326f
C856 VTAIL.n799 VSUBS 0.027516f
C857 VTAIL.n800 VSUBS 0.027516f
C858 VTAIL.n801 VSUBS 0.012326f
C859 VTAIL.n802 VSUBS 0.011641f
C860 VTAIL.n803 VSUBS 0.021664f
C861 VTAIL.n804 VSUBS 0.021664f
C862 VTAIL.n805 VSUBS 0.011641f
C863 VTAIL.n806 VSUBS 0.012326f
C864 VTAIL.n807 VSUBS 0.027516f
C865 VTAIL.n808 VSUBS 0.027516f
C866 VTAIL.n809 VSUBS 0.012326f
C867 VTAIL.n810 VSUBS 0.011641f
C868 VTAIL.n811 VSUBS 0.021664f
C869 VTAIL.n812 VSUBS 0.021664f
C870 VTAIL.n813 VSUBS 0.011641f
C871 VTAIL.n814 VSUBS 0.012326f
C872 VTAIL.n815 VSUBS 0.027516f
C873 VTAIL.n816 VSUBS 0.027516f
C874 VTAIL.n817 VSUBS 0.027516f
C875 VTAIL.n818 VSUBS 0.012326f
C876 VTAIL.n819 VSUBS 0.011641f
C877 VTAIL.n820 VSUBS 0.021664f
C878 VTAIL.n821 VSUBS 0.021664f
C879 VTAIL.n822 VSUBS 0.011641f
C880 VTAIL.n823 VSUBS 0.011984f
C881 VTAIL.n824 VSUBS 0.011984f
C882 VTAIL.n825 VSUBS 0.027516f
C883 VTAIL.n826 VSUBS 0.027516f
C884 VTAIL.n827 VSUBS 0.012326f
C885 VTAIL.n828 VSUBS 0.011641f
C886 VTAIL.n829 VSUBS 0.021664f
C887 VTAIL.n830 VSUBS 0.021664f
C888 VTAIL.n831 VSUBS 0.011641f
C889 VTAIL.n832 VSUBS 0.012326f
C890 VTAIL.n833 VSUBS 0.027516f
C891 VTAIL.n834 VSUBS 0.027516f
C892 VTAIL.n835 VSUBS 0.012326f
C893 VTAIL.n836 VSUBS 0.011641f
C894 VTAIL.n837 VSUBS 0.021664f
C895 VTAIL.n838 VSUBS 0.021664f
C896 VTAIL.n839 VSUBS 0.011641f
C897 VTAIL.n840 VSUBS 0.012326f
C898 VTAIL.n841 VSUBS 0.027516f
C899 VTAIL.n842 VSUBS 0.067869f
C900 VTAIL.n843 VSUBS 0.012326f
C901 VTAIL.n844 VSUBS 0.011641f
C902 VTAIL.n845 VSUBS 0.050371f
C903 VTAIL.n846 VSUBS 0.034195f
C904 VTAIL.n847 VSUBS 1.60212f
C905 VDD2.t3 VSUBS 0.399783f
C906 VDD2.t2 VSUBS 0.399783f
C907 VDD2.n0 VSUBS 4.26843f
C908 VDD2.t1 VSUBS 0.399783f
C909 VDD2.t0 VSUBS 0.399783f
C910 VDD2.n1 VSUBS 3.34189f
C911 VDD2.n2 VSUBS 4.76035f
C912 VN.t0 VSUBS 3.11716f
C913 VN.t1 VSUBS 3.1164f
C914 VN.n0 VSUBS 2.2266f
C915 VN.t2 VSUBS 3.11716f
C916 VN.t3 VSUBS 3.1164f
C917 VN.n1 VSUBS 3.96095f
C918 B.n0 VSUBS 0.004391f
C919 B.n1 VSUBS 0.004391f
C920 B.n2 VSUBS 0.006943f
C921 B.n3 VSUBS 0.006943f
C922 B.n4 VSUBS 0.006943f
C923 B.n5 VSUBS 0.006943f
C924 B.n6 VSUBS 0.006943f
C925 B.n7 VSUBS 0.006943f
C926 B.n8 VSUBS 0.006943f
C927 B.n9 VSUBS 0.006943f
C928 B.n10 VSUBS 0.006943f
C929 B.n11 VSUBS 0.006943f
C930 B.n12 VSUBS 0.006943f
C931 B.n13 VSUBS 0.015187f
C932 B.n14 VSUBS 0.006943f
C933 B.n15 VSUBS 0.006943f
C934 B.n16 VSUBS 0.006943f
C935 B.n17 VSUBS 0.006943f
C936 B.n18 VSUBS 0.006943f
C937 B.n19 VSUBS 0.006943f
C938 B.n20 VSUBS 0.006943f
C939 B.n21 VSUBS 0.006943f
C940 B.n22 VSUBS 0.006943f
C941 B.n23 VSUBS 0.006943f
C942 B.n24 VSUBS 0.006943f
C943 B.n25 VSUBS 0.006943f
C944 B.n26 VSUBS 0.006943f
C945 B.n27 VSUBS 0.006943f
C946 B.n28 VSUBS 0.006943f
C947 B.n29 VSUBS 0.006943f
C948 B.n30 VSUBS 0.006943f
C949 B.n31 VSUBS 0.006943f
C950 B.n32 VSUBS 0.006943f
C951 B.n33 VSUBS 0.006943f
C952 B.n34 VSUBS 0.006943f
C953 B.n35 VSUBS 0.006943f
C954 B.n36 VSUBS 0.006943f
C955 B.n37 VSUBS 0.006943f
C956 B.n38 VSUBS 0.006943f
C957 B.n39 VSUBS 0.006943f
C958 B.n40 VSUBS 0.006943f
C959 B.n41 VSUBS 0.006943f
C960 B.n42 VSUBS 0.006943f
C961 B.n43 VSUBS 0.006943f
C962 B.n44 VSUBS 0.006535f
C963 B.n45 VSUBS 0.006943f
C964 B.t2 VSUBS 0.371744f
C965 B.t1 VSUBS 0.391413f
C966 B.t0 VSUBS 1.06783f
C967 B.n46 VSUBS 0.529617f
C968 B.n47 VSUBS 0.332198f
C969 B.n48 VSUBS 0.016087f
C970 B.n49 VSUBS 0.006943f
C971 B.n50 VSUBS 0.006943f
C972 B.n51 VSUBS 0.006943f
C973 B.n52 VSUBS 0.006943f
C974 B.t8 VSUBS 0.371748f
C975 B.t7 VSUBS 0.391416f
C976 B.t6 VSUBS 1.06783f
C977 B.n53 VSUBS 0.529614f
C978 B.n54 VSUBS 0.332194f
C979 B.n55 VSUBS 0.006943f
C980 B.n56 VSUBS 0.006943f
C981 B.n57 VSUBS 0.006943f
C982 B.n58 VSUBS 0.006943f
C983 B.n59 VSUBS 0.006943f
C984 B.n60 VSUBS 0.006943f
C985 B.n61 VSUBS 0.006943f
C986 B.n62 VSUBS 0.006943f
C987 B.n63 VSUBS 0.006943f
C988 B.n64 VSUBS 0.006943f
C989 B.n65 VSUBS 0.006943f
C990 B.n66 VSUBS 0.006943f
C991 B.n67 VSUBS 0.006943f
C992 B.n68 VSUBS 0.006943f
C993 B.n69 VSUBS 0.006943f
C994 B.n70 VSUBS 0.006943f
C995 B.n71 VSUBS 0.006943f
C996 B.n72 VSUBS 0.006943f
C997 B.n73 VSUBS 0.006943f
C998 B.n74 VSUBS 0.006943f
C999 B.n75 VSUBS 0.006943f
C1000 B.n76 VSUBS 0.006943f
C1001 B.n77 VSUBS 0.006943f
C1002 B.n78 VSUBS 0.006943f
C1003 B.n79 VSUBS 0.006943f
C1004 B.n80 VSUBS 0.006943f
C1005 B.n81 VSUBS 0.006943f
C1006 B.n82 VSUBS 0.006943f
C1007 B.n83 VSUBS 0.006943f
C1008 B.n84 VSUBS 0.006943f
C1009 B.n85 VSUBS 0.015187f
C1010 B.n86 VSUBS 0.006943f
C1011 B.n87 VSUBS 0.006943f
C1012 B.n88 VSUBS 0.006943f
C1013 B.n89 VSUBS 0.006943f
C1014 B.n90 VSUBS 0.006943f
C1015 B.n91 VSUBS 0.006943f
C1016 B.n92 VSUBS 0.006943f
C1017 B.n93 VSUBS 0.006943f
C1018 B.n94 VSUBS 0.006943f
C1019 B.n95 VSUBS 0.006943f
C1020 B.n96 VSUBS 0.006943f
C1021 B.n97 VSUBS 0.006943f
C1022 B.n98 VSUBS 0.006943f
C1023 B.n99 VSUBS 0.006943f
C1024 B.n100 VSUBS 0.006943f
C1025 B.n101 VSUBS 0.006943f
C1026 B.n102 VSUBS 0.006943f
C1027 B.n103 VSUBS 0.006943f
C1028 B.n104 VSUBS 0.006943f
C1029 B.n105 VSUBS 0.006943f
C1030 B.n106 VSUBS 0.006943f
C1031 B.n107 VSUBS 0.006943f
C1032 B.n108 VSUBS 0.006943f
C1033 B.n109 VSUBS 0.016058f
C1034 B.n110 VSUBS 0.006943f
C1035 B.n111 VSUBS 0.006943f
C1036 B.n112 VSUBS 0.006943f
C1037 B.n113 VSUBS 0.006943f
C1038 B.n114 VSUBS 0.006943f
C1039 B.n115 VSUBS 0.006943f
C1040 B.n116 VSUBS 0.006943f
C1041 B.n117 VSUBS 0.006943f
C1042 B.n118 VSUBS 0.006943f
C1043 B.n119 VSUBS 0.006943f
C1044 B.n120 VSUBS 0.006943f
C1045 B.n121 VSUBS 0.006943f
C1046 B.n122 VSUBS 0.006943f
C1047 B.n123 VSUBS 0.006943f
C1048 B.n124 VSUBS 0.006943f
C1049 B.n125 VSUBS 0.006943f
C1050 B.n126 VSUBS 0.006943f
C1051 B.n127 VSUBS 0.006943f
C1052 B.n128 VSUBS 0.006943f
C1053 B.n129 VSUBS 0.006943f
C1054 B.n130 VSUBS 0.006943f
C1055 B.n131 VSUBS 0.006943f
C1056 B.n132 VSUBS 0.006943f
C1057 B.n133 VSUBS 0.006943f
C1058 B.n134 VSUBS 0.006943f
C1059 B.n135 VSUBS 0.006943f
C1060 B.n136 VSUBS 0.006943f
C1061 B.n137 VSUBS 0.006943f
C1062 B.n138 VSUBS 0.006943f
C1063 B.n139 VSUBS 0.006943f
C1064 B.n140 VSUBS 0.006943f
C1065 B.t4 VSUBS 0.371748f
C1066 B.t5 VSUBS 0.391416f
C1067 B.t3 VSUBS 1.06783f
C1068 B.n141 VSUBS 0.529614f
C1069 B.n142 VSUBS 0.332194f
C1070 B.n143 VSUBS 0.006943f
C1071 B.n144 VSUBS 0.006943f
C1072 B.n145 VSUBS 0.006943f
C1073 B.n146 VSUBS 0.006943f
C1074 B.t10 VSUBS 0.371744f
C1075 B.t11 VSUBS 0.391413f
C1076 B.t9 VSUBS 1.06783f
C1077 B.n147 VSUBS 0.529617f
C1078 B.n148 VSUBS 0.332198f
C1079 B.n149 VSUBS 0.016087f
C1080 B.n150 VSUBS 0.006943f
C1081 B.n151 VSUBS 0.006943f
C1082 B.n152 VSUBS 0.006943f
C1083 B.n153 VSUBS 0.006943f
C1084 B.n154 VSUBS 0.006943f
C1085 B.n155 VSUBS 0.006943f
C1086 B.n156 VSUBS 0.006943f
C1087 B.n157 VSUBS 0.006943f
C1088 B.n158 VSUBS 0.006943f
C1089 B.n159 VSUBS 0.006943f
C1090 B.n160 VSUBS 0.006943f
C1091 B.n161 VSUBS 0.006943f
C1092 B.n162 VSUBS 0.006943f
C1093 B.n163 VSUBS 0.006943f
C1094 B.n164 VSUBS 0.006943f
C1095 B.n165 VSUBS 0.006943f
C1096 B.n166 VSUBS 0.006943f
C1097 B.n167 VSUBS 0.006943f
C1098 B.n168 VSUBS 0.006943f
C1099 B.n169 VSUBS 0.006943f
C1100 B.n170 VSUBS 0.006943f
C1101 B.n171 VSUBS 0.006943f
C1102 B.n172 VSUBS 0.006943f
C1103 B.n173 VSUBS 0.006943f
C1104 B.n174 VSUBS 0.006943f
C1105 B.n175 VSUBS 0.006943f
C1106 B.n176 VSUBS 0.006943f
C1107 B.n177 VSUBS 0.006943f
C1108 B.n178 VSUBS 0.006943f
C1109 B.n179 VSUBS 0.006943f
C1110 B.n180 VSUBS 0.016058f
C1111 B.n181 VSUBS 0.006943f
C1112 B.n182 VSUBS 0.006943f
C1113 B.n183 VSUBS 0.006943f
C1114 B.n184 VSUBS 0.006943f
C1115 B.n185 VSUBS 0.006943f
C1116 B.n186 VSUBS 0.006943f
C1117 B.n187 VSUBS 0.006943f
C1118 B.n188 VSUBS 0.006943f
C1119 B.n189 VSUBS 0.006943f
C1120 B.n190 VSUBS 0.006943f
C1121 B.n191 VSUBS 0.006943f
C1122 B.n192 VSUBS 0.006943f
C1123 B.n193 VSUBS 0.006943f
C1124 B.n194 VSUBS 0.006943f
C1125 B.n195 VSUBS 0.006943f
C1126 B.n196 VSUBS 0.006943f
C1127 B.n197 VSUBS 0.006943f
C1128 B.n198 VSUBS 0.006943f
C1129 B.n199 VSUBS 0.006943f
C1130 B.n200 VSUBS 0.006943f
C1131 B.n201 VSUBS 0.006943f
C1132 B.n202 VSUBS 0.006943f
C1133 B.n203 VSUBS 0.006943f
C1134 B.n204 VSUBS 0.006943f
C1135 B.n205 VSUBS 0.006943f
C1136 B.n206 VSUBS 0.006943f
C1137 B.n207 VSUBS 0.006943f
C1138 B.n208 VSUBS 0.006943f
C1139 B.n209 VSUBS 0.006943f
C1140 B.n210 VSUBS 0.006943f
C1141 B.n211 VSUBS 0.006943f
C1142 B.n212 VSUBS 0.006943f
C1143 B.n213 VSUBS 0.006943f
C1144 B.n214 VSUBS 0.006943f
C1145 B.n215 VSUBS 0.006943f
C1146 B.n216 VSUBS 0.006943f
C1147 B.n217 VSUBS 0.006943f
C1148 B.n218 VSUBS 0.006943f
C1149 B.n219 VSUBS 0.006943f
C1150 B.n220 VSUBS 0.006943f
C1151 B.n221 VSUBS 0.006943f
C1152 B.n222 VSUBS 0.006943f
C1153 B.n223 VSUBS 0.015187f
C1154 B.n224 VSUBS 0.015187f
C1155 B.n225 VSUBS 0.016058f
C1156 B.n226 VSUBS 0.006943f
C1157 B.n227 VSUBS 0.006943f
C1158 B.n228 VSUBS 0.006943f
C1159 B.n229 VSUBS 0.006943f
C1160 B.n230 VSUBS 0.006943f
C1161 B.n231 VSUBS 0.006943f
C1162 B.n232 VSUBS 0.006943f
C1163 B.n233 VSUBS 0.006943f
C1164 B.n234 VSUBS 0.006943f
C1165 B.n235 VSUBS 0.006943f
C1166 B.n236 VSUBS 0.006943f
C1167 B.n237 VSUBS 0.006943f
C1168 B.n238 VSUBS 0.006943f
C1169 B.n239 VSUBS 0.006943f
C1170 B.n240 VSUBS 0.006943f
C1171 B.n241 VSUBS 0.006943f
C1172 B.n242 VSUBS 0.006943f
C1173 B.n243 VSUBS 0.006943f
C1174 B.n244 VSUBS 0.006943f
C1175 B.n245 VSUBS 0.006943f
C1176 B.n246 VSUBS 0.006943f
C1177 B.n247 VSUBS 0.006943f
C1178 B.n248 VSUBS 0.006943f
C1179 B.n249 VSUBS 0.006943f
C1180 B.n250 VSUBS 0.006943f
C1181 B.n251 VSUBS 0.006943f
C1182 B.n252 VSUBS 0.006943f
C1183 B.n253 VSUBS 0.006943f
C1184 B.n254 VSUBS 0.006943f
C1185 B.n255 VSUBS 0.006943f
C1186 B.n256 VSUBS 0.006943f
C1187 B.n257 VSUBS 0.006943f
C1188 B.n258 VSUBS 0.006943f
C1189 B.n259 VSUBS 0.006943f
C1190 B.n260 VSUBS 0.006943f
C1191 B.n261 VSUBS 0.006943f
C1192 B.n262 VSUBS 0.006943f
C1193 B.n263 VSUBS 0.006943f
C1194 B.n264 VSUBS 0.006943f
C1195 B.n265 VSUBS 0.006943f
C1196 B.n266 VSUBS 0.006943f
C1197 B.n267 VSUBS 0.006943f
C1198 B.n268 VSUBS 0.006943f
C1199 B.n269 VSUBS 0.006943f
C1200 B.n270 VSUBS 0.006943f
C1201 B.n271 VSUBS 0.006943f
C1202 B.n272 VSUBS 0.006943f
C1203 B.n273 VSUBS 0.006943f
C1204 B.n274 VSUBS 0.006943f
C1205 B.n275 VSUBS 0.006943f
C1206 B.n276 VSUBS 0.006943f
C1207 B.n277 VSUBS 0.006943f
C1208 B.n278 VSUBS 0.006943f
C1209 B.n279 VSUBS 0.006943f
C1210 B.n280 VSUBS 0.006943f
C1211 B.n281 VSUBS 0.006943f
C1212 B.n282 VSUBS 0.006943f
C1213 B.n283 VSUBS 0.006943f
C1214 B.n284 VSUBS 0.006943f
C1215 B.n285 VSUBS 0.006943f
C1216 B.n286 VSUBS 0.006943f
C1217 B.n287 VSUBS 0.006943f
C1218 B.n288 VSUBS 0.006943f
C1219 B.n289 VSUBS 0.006943f
C1220 B.n290 VSUBS 0.006943f
C1221 B.n291 VSUBS 0.006943f
C1222 B.n292 VSUBS 0.006943f
C1223 B.n293 VSUBS 0.006943f
C1224 B.n294 VSUBS 0.006943f
C1225 B.n295 VSUBS 0.006943f
C1226 B.n296 VSUBS 0.006943f
C1227 B.n297 VSUBS 0.006943f
C1228 B.n298 VSUBS 0.006943f
C1229 B.n299 VSUBS 0.006943f
C1230 B.n300 VSUBS 0.006943f
C1231 B.n301 VSUBS 0.006943f
C1232 B.n302 VSUBS 0.006943f
C1233 B.n303 VSUBS 0.006943f
C1234 B.n304 VSUBS 0.006943f
C1235 B.n305 VSUBS 0.006943f
C1236 B.n306 VSUBS 0.006943f
C1237 B.n307 VSUBS 0.006943f
C1238 B.n308 VSUBS 0.006943f
C1239 B.n309 VSUBS 0.006943f
C1240 B.n310 VSUBS 0.006943f
C1241 B.n311 VSUBS 0.006943f
C1242 B.n312 VSUBS 0.006943f
C1243 B.n313 VSUBS 0.006943f
C1244 B.n314 VSUBS 0.006943f
C1245 B.n315 VSUBS 0.006943f
C1246 B.n316 VSUBS 0.006535f
C1247 B.n317 VSUBS 0.006943f
C1248 B.n318 VSUBS 0.006943f
C1249 B.n319 VSUBS 0.00388f
C1250 B.n320 VSUBS 0.006943f
C1251 B.n321 VSUBS 0.006943f
C1252 B.n322 VSUBS 0.006943f
C1253 B.n323 VSUBS 0.006943f
C1254 B.n324 VSUBS 0.006943f
C1255 B.n325 VSUBS 0.006943f
C1256 B.n326 VSUBS 0.006943f
C1257 B.n327 VSUBS 0.006943f
C1258 B.n328 VSUBS 0.006943f
C1259 B.n329 VSUBS 0.006943f
C1260 B.n330 VSUBS 0.006943f
C1261 B.n331 VSUBS 0.006943f
C1262 B.n332 VSUBS 0.00388f
C1263 B.n333 VSUBS 0.016087f
C1264 B.n334 VSUBS 0.006535f
C1265 B.n335 VSUBS 0.006943f
C1266 B.n336 VSUBS 0.006943f
C1267 B.n337 VSUBS 0.006943f
C1268 B.n338 VSUBS 0.006943f
C1269 B.n339 VSUBS 0.006943f
C1270 B.n340 VSUBS 0.006943f
C1271 B.n341 VSUBS 0.006943f
C1272 B.n342 VSUBS 0.006943f
C1273 B.n343 VSUBS 0.006943f
C1274 B.n344 VSUBS 0.006943f
C1275 B.n345 VSUBS 0.006943f
C1276 B.n346 VSUBS 0.006943f
C1277 B.n347 VSUBS 0.006943f
C1278 B.n348 VSUBS 0.006943f
C1279 B.n349 VSUBS 0.006943f
C1280 B.n350 VSUBS 0.006943f
C1281 B.n351 VSUBS 0.006943f
C1282 B.n352 VSUBS 0.006943f
C1283 B.n353 VSUBS 0.006943f
C1284 B.n354 VSUBS 0.006943f
C1285 B.n355 VSUBS 0.006943f
C1286 B.n356 VSUBS 0.006943f
C1287 B.n357 VSUBS 0.006943f
C1288 B.n358 VSUBS 0.006943f
C1289 B.n359 VSUBS 0.006943f
C1290 B.n360 VSUBS 0.006943f
C1291 B.n361 VSUBS 0.006943f
C1292 B.n362 VSUBS 0.006943f
C1293 B.n363 VSUBS 0.006943f
C1294 B.n364 VSUBS 0.006943f
C1295 B.n365 VSUBS 0.006943f
C1296 B.n366 VSUBS 0.006943f
C1297 B.n367 VSUBS 0.006943f
C1298 B.n368 VSUBS 0.006943f
C1299 B.n369 VSUBS 0.006943f
C1300 B.n370 VSUBS 0.006943f
C1301 B.n371 VSUBS 0.006943f
C1302 B.n372 VSUBS 0.006943f
C1303 B.n373 VSUBS 0.006943f
C1304 B.n374 VSUBS 0.006943f
C1305 B.n375 VSUBS 0.006943f
C1306 B.n376 VSUBS 0.006943f
C1307 B.n377 VSUBS 0.006943f
C1308 B.n378 VSUBS 0.006943f
C1309 B.n379 VSUBS 0.006943f
C1310 B.n380 VSUBS 0.006943f
C1311 B.n381 VSUBS 0.006943f
C1312 B.n382 VSUBS 0.006943f
C1313 B.n383 VSUBS 0.006943f
C1314 B.n384 VSUBS 0.006943f
C1315 B.n385 VSUBS 0.006943f
C1316 B.n386 VSUBS 0.006943f
C1317 B.n387 VSUBS 0.006943f
C1318 B.n388 VSUBS 0.006943f
C1319 B.n389 VSUBS 0.006943f
C1320 B.n390 VSUBS 0.006943f
C1321 B.n391 VSUBS 0.006943f
C1322 B.n392 VSUBS 0.006943f
C1323 B.n393 VSUBS 0.006943f
C1324 B.n394 VSUBS 0.006943f
C1325 B.n395 VSUBS 0.006943f
C1326 B.n396 VSUBS 0.006943f
C1327 B.n397 VSUBS 0.006943f
C1328 B.n398 VSUBS 0.006943f
C1329 B.n399 VSUBS 0.006943f
C1330 B.n400 VSUBS 0.006943f
C1331 B.n401 VSUBS 0.006943f
C1332 B.n402 VSUBS 0.006943f
C1333 B.n403 VSUBS 0.006943f
C1334 B.n404 VSUBS 0.006943f
C1335 B.n405 VSUBS 0.006943f
C1336 B.n406 VSUBS 0.006943f
C1337 B.n407 VSUBS 0.006943f
C1338 B.n408 VSUBS 0.006943f
C1339 B.n409 VSUBS 0.006943f
C1340 B.n410 VSUBS 0.006943f
C1341 B.n411 VSUBS 0.006943f
C1342 B.n412 VSUBS 0.006943f
C1343 B.n413 VSUBS 0.006943f
C1344 B.n414 VSUBS 0.006943f
C1345 B.n415 VSUBS 0.006943f
C1346 B.n416 VSUBS 0.006943f
C1347 B.n417 VSUBS 0.006943f
C1348 B.n418 VSUBS 0.006943f
C1349 B.n419 VSUBS 0.006943f
C1350 B.n420 VSUBS 0.006943f
C1351 B.n421 VSUBS 0.006943f
C1352 B.n422 VSUBS 0.006943f
C1353 B.n423 VSUBS 0.006943f
C1354 B.n424 VSUBS 0.006943f
C1355 B.n425 VSUBS 0.006943f
C1356 B.n426 VSUBS 0.016058f
C1357 B.n427 VSUBS 0.015187f
C1358 B.n428 VSUBS 0.015187f
C1359 B.n429 VSUBS 0.006943f
C1360 B.n430 VSUBS 0.006943f
C1361 B.n431 VSUBS 0.006943f
C1362 B.n432 VSUBS 0.006943f
C1363 B.n433 VSUBS 0.006943f
C1364 B.n434 VSUBS 0.006943f
C1365 B.n435 VSUBS 0.006943f
C1366 B.n436 VSUBS 0.006943f
C1367 B.n437 VSUBS 0.006943f
C1368 B.n438 VSUBS 0.006943f
C1369 B.n439 VSUBS 0.006943f
C1370 B.n440 VSUBS 0.006943f
C1371 B.n441 VSUBS 0.006943f
C1372 B.n442 VSUBS 0.006943f
C1373 B.n443 VSUBS 0.006943f
C1374 B.n444 VSUBS 0.006943f
C1375 B.n445 VSUBS 0.006943f
C1376 B.n446 VSUBS 0.006943f
C1377 B.n447 VSUBS 0.006943f
C1378 B.n448 VSUBS 0.006943f
C1379 B.n449 VSUBS 0.006943f
C1380 B.n450 VSUBS 0.006943f
C1381 B.n451 VSUBS 0.006943f
C1382 B.n452 VSUBS 0.006943f
C1383 B.n453 VSUBS 0.006943f
C1384 B.n454 VSUBS 0.006943f
C1385 B.n455 VSUBS 0.006943f
C1386 B.n456 VSUBS 0.006943f
C1387 B.n457 VSUBS 0.006943f
C1388 B.n458 VSUBS 0.006943f
C1389 B.n459 VSUBS 0.006943f
C1390 B.n460 VSUBS 0.006943f
C1391 B.n461 VSUBS 0.006943f
C1392 B.n462 VSUBS 0.006943f
C1393 B.n463 VSUBS 0.006943f
C1394 B.n464 VSUBS 0.006943f
C1395 B.n465 VSUBS 0.006943f
C1396 B.n466 VSUBS 0.006943f
C1397 B.n467 VSUBS 0.006943f
C1398 B.n468 VSUBS 0.006943f
C1399 B.n469 VSUBS 0.006943f
C1400 B.n470 VSUBS 0.006943f
C1401 B.n471 VSUBS 0.006943f
C1402 B.n472 VSUBS 0.006943f
C1403 B.n473 VSUBS 0.006943f
C1404 B.n474 VSUBS 0.006943f
C1405 B.n475 VSUBS 0.006943f
C1406 B.n476 VSUBS 0.006943f
C1407 B.n477 VSUBS 0.006943f
C1408 B.n478 VSUBS 0.006943f
C1409 B.n479 VSUBS 0.006943f
C1410 B.n480 VSUBS 0.006943f
C1411 B.n481 VSUBS 0.006943f
C1412 B.n482 VSUBS 0.006943f
C1413 B.n483 VSUBS 0.006943f
C1414 B.n484 VSUBS 0.006943f
C1415 B.n485 VSUBS 0.006943f
C1416 B.n486 VSUBS 0.006943f
C1417 B.n487 VSUBS 0.006943f
C1418 B.n488 VSUBS 0.006943f
C1419 B.n489 VSUBS 0.006943f
C1420 B.n490 VSUBS 0.006943f
C1421 B.n491 VSUBS 0.006943f
C1422 B.n492 VSUBS 0.006943f
C1423 B.n493 VSUBS 0.006943f
C1424 B.n494 VSUBS 0.006943f
C1425 B.n495 VSUBS 0.006943f
C1426 B.n496 VSUBS 0.016058f
C1427 B.n497 VSUBS 0.015187f
C1428 B.n498 VSUBS 0.016058f
C1429 B.n499 VSUBS 0.006943f
C1430 B.n500 VSUBS 0.006943f
C1431 B.n501 VSUBS 0.006943f
C1432 B.n502 VSUBS 0.006943f
C1433 B.n503 VSUBS 0.006943f
C1434 B.n504 VSUBS 0.006943f
C1435 B.n505 VSUBS 0.006943f
C1436 B.n506 VSUBS 0.006943f
C1437 B.n507 VSUBS 0.006943f
C1438 B.n508 VSUBS 0.006943f
C1439 B.n509 VSUBS 0.006943f
C1440 B.n510 VSUBS 0.006943f
C1441 B.n511 VSUBS 0.006943f
C1442 B.n512 VSUBS 0.006943f
C1443 B.n513 VSUBS 0.006943f
C1444 B.n514 VSUBS 0.006943f
C1445 B.n515 VSUBS 0.006943f
C1446 B.n516 VSUBS 0.006943f
C1447 B.n517 VSUBS 0.006943f
C1448 B.n518 VSUBS 0.006943f
C1449 B.n519 VSUBS 0.006943f
C1450 B.n520 VSUBS 0.006943f
C1451 B.n521 VSUBS 0.006943f
C1452 B.n522 VSUBS 0.006943f
C1453 B.n523 VSUBS 0.006943f
C1454 B.n524 VSUBS 0.006943f
C1455 B.n525 VSUBS 0.006943f
C1456 B.n526 VSUBS 0.006943f
C1457 B.n527 VSUBS 0.006943f
C1458 B.n528 VSUBS 0.006943f
C1459 B.n529 VSUBS 0.006943f
C1460 B.n530 VSUBS 0.006943f
C1461 B.n531 VSUBS 0.006943f
C1462 B.n532 VSUBS 0.006943f
C1463 B.n533 VSUBS 0.006943f
C1464 B.n534 VSUBS 0.006943f
C1465 B.n535 VSUBS 0.006943f
C1466 B.n536 VSUBS 0.006943f
C1467 B.n537 VSUBS 0.006943f
C1468 B.n538 VSUBS 0.006943f
C1469 B.n539 VSUBS 0.006943f
C1470 B.n540 VSUBS 0.006943f
C1471 B.n541 VSUBS 0.006943f
C1472 B.n542 VSUBS 0.006943f
C1473 B.n543 VSUBS 0.006943f
C1474 B.n544 VSUBS 0.006943f
C1475 B.n545 VSUBS 0.006943f
C1476 B.n546 VSUBS 0.006943f
C1477 B.n547 VSUBS 0.006943f
C1478 B.n548 VSUBS 0.006943f
C1479 B.n549 VSUBS 0.006943f
C1480 B.n550 VSUBS 0.006943f
C1481 B.n551 VSUBS 0.006943f
C1482 B.n552 VSUBS 0.006943f
C1483 B.n553 VSUBS 0.006943f
C1484 B.n554 VSUBS 0.006943f
C1485 B.n555 VSUBS 0.006943f
C1486 B.n556 VSUBS 0.006943f
C1487 B.n557 VSUBS 0.006943f
C1488 B.n558 VSUBS 0.006943f
C1489 B.n559 VSUBS 0.006943f
C1490 B.n560 VSUBS 0.006943f
C1491 B.n561 VSUBS 0.006943f
C1492 B.n562 VSUBS 0.006943f
C1493 B.n563 VSUBS 0.006943f
C1494 B.n564 VSUBS 0.006943f
C1495 B.n565 VSUBS 0.006943f
C1496 B.n566 VSUBS 0.006943f
C1497 B.n567 VSUBS 0.006943f
C1498 B.n568 VSUBS 0.006943f
C1499 B.n569 VSUBS 0.006943f
C1500 B.n570 VSUBS 0.006943f
C1501 B.n571 VSUBS 0.006943f
C1502 B.n572 VSUBS 0.006943f
C1503 B.n573 VSUBS 0.006943f
C1504 B.n574 VSUBS 0.006943f
C1505 B.n575 VSUBS 0.006943f
C1506 B.n576 VSUBS 0.006943f
C1507 B.n577 VSUBS 0.006943f
C1508 B.n578 VSUBS 0.006943f
C1509 B.n579 VSUBS 0.006943f
C1510 B.n580 VSUBS 0.006943f
C1511 B.n581 VSUBS 0.006943f
C1512 B.n582 VSUBS 0.006943f
C1513 B.n583 VSUBS 0.006943f
C1514 B.n584 VSUBS 0.006943f
C1515 B.n585 VSUBS 0.006943f
C1516 B.n586 VSUBS 0.006943f
C1517 B.n587 VSUBS 0.006943f
C1518 B.n588 VSUBS 0.006943f
C1519 B.n589 VSUBS 0.006943f
C1520 B.n590 VSUBS 0.006535f
C1521 B.n591 VSUBS 0.016087f
C1522 B.n592 VSUBS 0.00388f
C1523 B.n593 VSUBS 0.006943f
C1524 B.n594 VSUBS 0.006943f
C1525 B.n595 VSUBS 0.006943f
C1526 B.n596 VSUBS 0.006943f
C1527 B.n597 VSUBS 0.006943f
C1528 B.n598 VSUBS 0.006943f
C1529 B.n599 VSUBS 0.006943f
C1530 B.n600 VSUBS 0.006943f
C1531 B.n601 VSUBS 0.006943f
C1532 B.n602 VSUBS 0.006943f
C1533 B.n603 VSUBS 0.006943f
C1534 B.n604 VSUBS 0.006943f
C1535 B.n605 VSUBS 0.00388f
C1536 B.n606 VSUBS 0.006943f
C1537 B.n607 VSUBS 0.006943f
C1538 B.n608 VSUBS 0.006943f
C1539 B.n609 VSUBS 0.006943f
C1540 B.n610 VSUBS 0.006943f
C1541 B.n611 VSUBS 0.006943f
C1542 B.n612 VSUBS 0.006943f
C1543 B.n613 VSUBS 0.006943f
C1544 B.n614 VSUBS 0.006943f
C1545 B.n615 VSUBS 0.006943f
C1546 B.n616 VSUBS 0.006943f
C1547 B.n617 VSUBS 0.006943f
C1548 B.n618 VSUBS 0.006943f
C1549 B.n619 VSUBS 0.006943f
C1550 B.n620 VSUBS 0.006943f
C1551 B.n621 VSUBS 0.006943f
C1552 B.n622 VSUBS 0.006943f
C1553 B.n623 VSUBS 0.006943f
C1554 B.n624 VSUBS 0.006943f
C1555 B.n625 VSUBS 0.006943f
C1556 B.n626 VSUBS 0.006943f
C1557 B.n627 VSUBS 0.006943f
C1558 B.n628 VSUBS 0.006943f
C1559 B.n629 VSUBS 0.006943f
C1560 B.n630 VSUBS 0.006943f
C1561 B.n631 VSUBS 0.006943f
C1562 B.n632 VSUBS 0.006943f
C1563 B.n633 VSUBS 0.006943f
C1564 B.n634 VSUBS 0.006943f
C1565 B.n635 VSUBS 0.006943f
C1566 B.n636 VSUBS 0.006943f
C1567 B.n637 VSUBS 0.006943f
C1568 B.n638 VSUBS 0.006943f
C1569 B.n639 VSUBS 0.006943f
C1570 B.n640 VSUBS 0.006943f
C1571 B.n641 VSUBS 0.006943f
C1572 B.n642 VSUBS 0.006943f
C1573 B.n643 VSUBS 0.006943f
C1574 B.n644 VSUBS 0.006943f
C1575 B.n645 VSUBS 0.006943f
C1576 B.n646 VSUBS 0.006943f
C1577 B.n647 VSUBS 0.006943f
C1578 B.n648 VSUBS 0.006943f
C1579 B.n649 VSUBS 0.006943f
C1580 B.n650 VSUBS 0.006943f
C1581 B.n651 VSUBS 0.006943f
C1582 B.n652 VSUBS 0.006943f
C1583 B.n653 VSUBS 0.006943f
C1584 B.n654 VSUBS 0.006943f
C1585 B.n655 VSUBS 0.006943f
C1586 B.n656 VSUBS 0.006943f
C1587 B.n657 VSUBS 0.006943f
C1588 B.n658 VSUBS 0.006943f
C1589 B.n659 VSUBS 0.006943f
C1590 B.n660 VSUBS 0.006943f
C1591 B.n661 VSUBS 0.006943f
C1592 B.n662 VSUBS 0.006943f
C1593 B.n663 VSUBS 0.006943f
C1594 B.n664 VSUBS 0.006943f
C1595 B.n665 VSUBS 0.006943f
C1596 B.n666 VSUBS 0.006943f
C1597 B.n667 VSUBS 0.006943f
C1598 B.n668 VSUBS 0.006943f
C1599 B.n669 VSUBS 0.006943f
C1600 B.n670 VSUBS 0.006943f
C1601 B.n671 VSUBS 0.006943f
C1602 B.n672 VSUBS 0.006943f
C1603 B.n673 VSUBS 0.006943f
C1604 B.n674 VSUBS 0.006943f
C1605 B.n675 VSUBS 0.006943f
C1606 B.n676 VSUBS 0.006943f
C1607 B.n677 VSUBS 0.006943f
C1608 B.n678 VSUBS 0.006943f
C1609 B.n679 VSUBS 0.006943f
C1610 B.n680 VSUBS 0.006943f
C1611 B.n681 VSUBS 0.006943f
C1612 B.n682 VSUBS 0.006943f
C1613 B.n683 VSUBS 0.006943f
C1614 B.n684 VSUBS 0.006943f
C1615 B.n685 VSUBS 0.006943f
C1616 B.n686 VSUBS 0.006943f
C1617 B.n687 VSUBS 0.006943f
C1618 B.n688 VSUBS 0.006943f
C1619 B.n689 VSUBS 0.006943f
C1620 B.n690 VSUBS 0.006943f
C1621 B.n691 VSUBS 0.006943f
C1622 B.n692 VSUBS 0.006943f
C1623 B.n693 VSUBS 0.006943f
C1624 B.n694 VSUBS 0.006943f
C1625 B.n695 VSUBS 0.006943f
C1626 B.n696 VSUBS 0.006943f
C1627 B.n697 VSUBS 0.006943f
C1628 B.n698 VSUBS 0.016058f
C1629 B.n699 VSUBS 0.016058f
C1630 B.n700 VSUBS 0.015187f
C1631 B.n701 VSUBS 0.006943f
C1632 B.n702 VSUBS 0.006943f
C1633 B.n703 VSUBS 0.006943f
C1634 B.n704 VSUBS 0.006943f
C1635 B.n705 VSUBS 0.006943f
C1636 B.n706 VSUBS 0.006943f
C1637 B.n707 VSUBS 0.006943f
C1638 B.n708 VSUBS 0.006943f
C1639 B.n709 VSUBS 0.006943f
C1640 B.n710 VSUBS 0.006943f
C1641 B.n711 VSUBS 0.006943f
C1642 B.n712 VSUBS 0.006943f
C1643 B.n713 VSUBS 0.006943f
C1644 B.n714 VSUBS 0.006943f
C1645 B.n715 VSUBS 0.006943f
C1646 B.n716 VSUBS 0.006943f
C1647 B.n717 VSUBS 0.006943f
C1648 B.n718 VSUBS 0.006943f
C1649 B.n719 VSUBS 0.006943f
C1650 B.n720 VSUBS 0.006943f
C1651 B.n721 VSUBS 0.006943f
C1652 B.n722 VSUBS 0.006943f
C1653 B.n723 VSUBS 0.006943f
C1654 B.n724 VSUBS 0.006943f
C1655 B.n725 VSUBS 0.006943f
C1656 B.n726 VSUBS 0.006943f
C1657 B.n727 VSUBS 0.006943f
C1658 B.n728 VSUBS 0.006943f
C1659 B.n729 VSUBS 0.006943f
C1660 B.n730 VSUBS 0.006943f
C1661 B.n731 VSUBS 0.006943f
C1662 B.n732 VSUBS 0.006943f
C1663 B.n733 VSUBS 0.006943f
C1664 B.n734 VSUBS 0.006943f
C1665 B.n735 VSUBS 0.015722f
.ends

