* NGSPICE file created from diff_pair_sample_0621.ext - technology: sky130A

.subckt diff_pair_sample_0621 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t18 VN.t0 VDD2.t8 B.t2 sky130_fd_pr__nfet_01v8 ad=1.51965 pd=9.54 as=1.51965 ps=9.54 w=9.21 l=3.35
X1 VDD1.t9 VP.t0 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=3.5919 pd=19.2 as=1.51965 ps=9.54 w=9.21 l=3.35
X2 VDD1.t8 VP.t1 VTAIL.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=1.51965 pd=9.54 as=1.51965 ps=9.54 w=9.21 l=3.35
X3 VDD2.t3 VN.t1 VTAIL.t17 B.t6 sky130_fd_pr__nfet_01v8 ad=3.5919 pd=19.2 as=1.51965 ps=9.54 w=9.21 l=3.35
X4 VTAIL.t16 VN.t2 VDD2.t4 B.t9 sky130_fd_pr__nfet_01v8 ad=1.51965 pd=9.54 as=1.51965 ps=9.54 w=9.21 l=3.35
X5 B.t23 B.t21 B.t22 B.t18 sky130_fd_pr__nfet_01v8 ad=3.5919 pd=19.2 as=0 ps=0 w=9.21 l=3.35
X6 VDD2.t0 VN.t3 VTAIL.t15 B.t0 sky130_fd_pr__nfet_01v8 ad=1.51965 pd=9.54 as=3.5919 ps=19.2 w=9.21 l=3.35
X7 VDD2.t2 VN.t4 VTAIL.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=3.5919 pd=19.2 as=1.51965 ps=9.54 w=9.21 l=3.35
X8 VTAIL.t2 VP.t2 VDD1.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=1.51965 pd=9.54 as=1.51965 ps=9.54 w=9.21 l=3.35
X9 VDD2.t1 VN.t5 VTAIL.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=1.51965 pd=9.54 as=1.51965 ps=9.54 w=9.21 l=3.35
X10 B.t20 B.t17 B.t19 B.t18 sky130_fd_pr__nfet_01v8 ad=3.5919 pd=19.2 as=0 ps=0 w=9.21 l=3.35
X11 VTAIL.t1 VP.t3 VDD1.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=1.51965 pd=9.54 as=1.51965 ps=9.54 w=9.21 l=3.35
X12 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=3.5919 pd=19.2 as=0 ps=0 w=9.21 l=3.35
X13 VDD1.t5 VP.t4 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.51965 pd=9.54 as=1.51965 ps=9.54 w=9.21 l=3.35
X14 VDD2.t6 VN.t6 VTAIL.t12 B.t8 sky130_fd_pr__nfet_01v8 ad=1.51965 pd=9.54 as=1.51965 ps=9.54 w=9.21 l=3.35
X15 VDD1.t4 VP.t5 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.51965 pd=9.54 as=3.5919 ps=19.2 w=9.21 l=3.35
X16 VDD2.t7 VN.t7 VTAIL.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=1.51965 pd=9.54 as=3.5919 ps=19.2 w=9.21 l=3.35
X17 VTAIL.t10 VN.t8 VDD2.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=1.51965 pd=9.54 as=1.51965 ps=9.54 w=9.21 l=3.35
X18 VDD1.t3 VP.t6 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=3.5919 pd=19.2 as=1.51965 ps=9.54 w=9.21 l=3.35
X19 VTAIL.t4 VP.t7 VDD1.t2 B.t4 sky130_fd_pr__nfet_01v8 ad=1.51965 pd=9.54 as=1.51965 ps=9.54 w=9.21 l=3.35
X20 VTAIL.t9 VN.t9 VDD2.t9 B.t4 sky130_fd_pr__nfet_01v8 ad=1.51965 pd=9.54 as=1.51965 ps=9.54 w=9.21 l=3.35
X21 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=3.5919 pd=19.2 as=0 ps=0 w=9.21 l=3.35
X22 VDD1.t1 VP.t8 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.51965 pd=9.54 as=3.5919 ps=19.2 w=9.21 l=3.35
X23 VTAIL.t19 VP.t9 VDD1.t0 B.t9 sky130_fd_pr__nfet_01v8 ad=1.51965 pd=9.54 as=1.51965 ps=9.54 w=9.21 l=3.35
R0 VN.n96 VN.n95 161.3
R1 VN.n94 VN.n50 161.3
R2 VN.n93 VN.n92 161.3
R3 VN.n91 VN.n51 161.3
R4 VN.n90 VN.n89 161.3
R5 VN.n88 VN.n52 161.3
R6 VN.n87 VN.n86 161.3
R7 VN.n85 VN.n84 161.3
R8 VN.n83 VN.n54 161.3
R9 VN.n82 VN.n81 161.3
R10 VN.n80 VN.n55 161.3
R11 VN.n79 VN.n78 161.3
R12 VN.n77 VN.n56 161.3
R13 VN.n76 VN.n75 161.3
R14 VN.n74 VN.n57 161.3
R15 VN.n73 VN.n72 161.3
R16 VN.n71 VN.n58 161.3
R17 VN.n70 VN.n69 161.3
R18 VN.n68 VN.n59 161.3
R19 VN.n67 VN.n66 161.3
R20 VN.n65 VN.n60 161.3
R21 VN.n64 VN.n63 161.3
R22 VN.n47 VN.n46 161.3
R23 VN.n45 VN.n1 161.3
R24 VN.n44 VN.n43 161.3
R25 VN.n42 VN.n2 161.3
R26 VN.n41 VN.n40 161.3
R27 VN.n39 VN.n3 161.3
R28 VN.n38 VN.n37 161.3
R29 VN.n36 VN.n35 161.3
R30 VN.n34 VN.n5 161.3
R31 VN.n33 VN.n32 161.3
R32 VN.n31 VN.n6 161.3
R33 VN.n30 VN.n29 161.3
R34 VN.n28 VN.n7 161.3
R35 VN.n27 VN.n26 161.3
R36 VN.n25 VN.n8 161.3
R37 VN.n24 VN.n23 161.3
R38 VN.n22 VN.n9 161.3
R39 VN.n21 VN.n20 161.3
R40 VN.n19 VN.n10 161.3
R41 VN.n18 VN.n17 161.3
R42 VN.n16 VN.n11 161.3
R43 VN.n15 VN.n14 161.3
R44 VN.n13 VN.t4 99.435
R45 VN.n62 VN.t7 99.435
R46 VN.n48 VN.n0 72.4512
R47 VN.n97 VN.n49 72.4512
R48 VN.n8 VN.t6 66.2575
R49 VN.n12 VN.t0 66.2575
R50 VN.n4 VN.t8 66.2575
R51 VN.n0 VN.t3 66.2575
R52 VN.n57 VN.t5 66.2575
R53 VN.n61 VN.t9 66.2575
R54 VN.n53 VN.t2 66.2575
R55 VN.n49 VN.t1 66.2575
R56 VN.n62 VN.n61 65.6329
R57 VN.n13 VN.n12 65.6329
R58 VN.n21 VN.n10 56.0336
R59 VN.n29 VN.n6 56.0336
R60 VN.n70 VN.n59 56.0336
R61 VN.n78 VN.n55 56.0336
R62 VN VN.n97 55.4147
R63 VN.n44 VN.n2 42.4359
R64 VN.n93 VN.n51 42.4359
R65 VN.n40 VN.n2 38.5509
R66 VN.n89 VN.n51 38.5509
R67 VN.n17 VN.n10 24.9531
R68 VN.n33 VN.n6 24.9531
R69 VN.n66 VN.n59 24.9531
R70 VN.n82 VN.n55 24.9531
R71 VN.n16 VN.n15 24.4675
R72 VN.n17 VN.n16 24.4675
R73 VN.n22 VN.n21 24.4675
R74 VN.n23 VN.n22 24.4675
R75 VN.n23 VN.n8 24.4675
R76 VN.n27 VN.n8 24.4675
R77 VN.n28 VN.n27 24.4675
R78 VN.n29 VN.n28 24.4675
R79 VN.n34 VN.n33 24.4675
R80 VN.n35 VN.n34 24.4675
R81 VN.n39 VN.n38 24.4675
R82 VN.n40 VN.n39 24.4675
R83 VN.n45 VN.n44 24.4675
R84 VN.n46 VN.n45 24.4675
R85 VN.n66 VN.n65 24.4675
R86 VN.n65 VN.n64 24.4675
R87 VN.n78 VN.n77 24.4675
R88 VN.n77 VN.n76 24.4675
R89 VN.n76 VN.n57 24.4675
R90 VN.n72 VN.n57 24.4675
R91 VN.n72 VN.n71 24.4675
R92 VN.n71 VN.n70 24.4675
R93 VN.n89 VN.n88 24.4675
R94 VN.n88 VN.n87 24.4675
R95 VN.n84 VN.n83 24.4675
R96 VN.n83 VN.n82 24.4675
R97 VN.n95 VN.n94 24.4675
R98 VN.n94 VN.n93 24.4675
R99 VN.n46 VN.n0 17.6167
R100 VN.n95 VN.n49 17.6167
R101 VN.n38 VN.n4 15.6594
R102 VN.n87 VN.n53 15.6594
R103 VN.n15 VN.n12 8.80862
R104 VN.n35 VN.n4 8.80862
R105 VN.n64 VN.n61 8.80862
R106 VN.n84 VN.n53 8.80862
R107 VN.n63 VN.n62 4.01768
R108 VN.n14 VN.n13 4.01768
R109 VN.n97 VN.n96 0.354971
R110 VN.n48 VN.n47 0.354971
R111 VN VN.n48 0.26696
R112 VN.n96 VN.n50 0.189894
R113 VN.n92 VN.n50 0.189894
R114 VN.n92 VN.n91 0.189894
R115 VN.n91 VN.n90 0.189894
R116 VN.n90 VN.n52 0.189894
R117 VN.n86 VN.n52 0.189894
R118 VN.n86 VN.n85 0.189894
R119 VN.n85 VN.n54 0.189894
R120 VN.n81 VN.n54 0.189894
R121 VN.n81 VN.n80 0.189894
R122 VN.n80 VN.n79 0.189894
R123 VN.n79 VN.n56 0.189894
R124 VN.n75 VN.n56 0.189894
R125 VN.n75 VN.n74 0.189894
R126 VN.n74 VN.n73 0.189894
R127 VN.n73 VN.n58 0.189894
R128 VN.n69 VN.n58 0.189894
R129 VN.n69 VN.n68 0.189894
R130 VN.n68 VN.n67 0.189894
R131 VN.n67 VN.n60 0.189894
R132 VN.n63 VN.n60 0.189894
R133 VN.n14 VN.n11 0.189894
R134 VN.n18 VN.n11 0.189894
R135 VN.n19 VN.n18 0.189894
R136 VN.n20 VN.n19 0.189894
R137 VN.n20 VN.n9 0.189894
R138 VN.n24 VN.n9 0.189894
R139 VN.n25 VN.n24 0.189894
R140 VN.n26 VN.n25 0.189894
R141 VN.n26 VN.n7 0.189894
R142 VN.n30 VN.n7 0.189894
R143 VN.n31 VN.n30 0.189894
R144 VN.n32 VN.n31 0.189894
R145 VN.n32 VN.n5 0.189894
R146 VN.n36 VN.n5 0.189894
R147 VN.n37 VN.n36 0.189894
R148 VN.n37 VN.n3 0.189894
R149 VN.n41 VN.n3 0.189894
R150 VN.n42 VN.n41 0.189894
R151 VN.n43 VN.n42 0.189894
R152 VN.n43 VN.n1 0.189894
R153 VN.n47 VN.n1 0.189894
R154 VDD2.n97 VDD2.n53 289.615
R155 VDD2.n44 VDD2.n0 289.615
R156 VDD2.n98 VDD2.n97 185
R157 VDD2.n96 VDD2.n95 185
R158 VDD2.n57 VDD2.n56 185
R159 VDD2.n61 VDD2.n59 185
R160 VDD2.n90 VDD2.n89 185
R161 VDD2.n88 VDD2.n87 185
R162 VDD2.n63 VDD2.n62 185
R163 VDD2.n82 VDD2.n81 185
R164 VDD2.n80 VDD2.n79 185
R165 VDD2.n67 VDD2.n66 185
R166 VDD2.n74 VDD2.n73 185
R167 VDD2.n72 VDD2.n71 185
R168 VDD2.n17 VDD2.n16 185
R169 VDD2.n19 VDD2.n18 185
R170 VDD2.n12 VDD2.n11 185
R171 VDD2.n25 VDD2.n24 185
R172 VDD2.n27 VDD2.n26 185
R173 VDD2.n8 VDD2.n7 185
R174 VDD2.n34 VDD2.n33 185
R175 VDD2.n35 VDD2.n6 185
R176 VDD2.n37 VDD2.n36 185
R177 VDD2.n4 VDD2.n3 185
R178 VDD2.n43 VDD2.n42 185
R179 VDD2.n45 VDD2.n44 185
R180 VDD2.n70 VDD2.t3 149.524
R181 VDD2.n15 VDD2.t2 149.524
R182 VDD2.n97 VDD2.n96 104.615
R183 VDD2.n96 VDD2.n56 104.615
R184 VDD2.n61 VDD2.n56 104.615
R185 VDD2.n89 VDD2.n61 104.615
R186 VDD2.n89 VDD2.n88 104.615
R187 VDD2.n88 VDD2.n62 104.615
R188 VDD2.n81 VDD2.n62 104.615
R189 VDD2.n81 VDD2.n80 104.615
R190 VDD2.n80 VDD2.n66 104.615
R191 VDD2.n73 VDD2.n66 104.615
R192 VDD2.n73 VDD2.n72 104.615
R193 VDD2.n18 VDD2.n17 104.615
R194 VDD2.n18 VDD2.n11 104.615
R195 VDD2.n25 VDD2.n11 104.615
R196 VDD2.n26 VDD2.n25 104.615
R197 VDD2.n26 VDD2.n7 104.615
R198 VDD2.n34 VDD2.n7 104.615
R199 VDD2.n35 VDD2.n34 104.615
R200 VDD2.n36 VDD2.n35 104.615
R201 VDD2.n36 VDD2.n3 104.615
R202 VDD2.n43 VDD2.n3 104.615
R203 VDD2.n44 VDD2.n43 104.615
R204 VDD2.n52 VDD2.n51 64.744
R205 VDD2 VDD2.n105 64.7412
R206 VDD2.n104 VDD2.n103 62.4202
R207 VDD2.n50 VDD2.n49 62.4201
R208 VDD2.n72 VDD2.t3 52.3082
R209 VDD2.n17 VDD2.t2 52.3082
R210 VDD2.n50 VDD2.n48 51.4547
R211 VDD2.n102 VDD2.n101 48.2823
R212 VDD2.n102 VDD2.n52 46.7239
R213 VDD2.n59 VDD2.n57 13.1884
R214 VDD2.n37 VDD2.n4 13.1884
R215 VDD2.n95 VDD2.n94 12.8005
R216 VDD2.n91 VDD2.n90 12.8005
R217 VDD2.n38 VDD2.n6 12.8005
R218 VDD2.n42 VDD2.n41 12.8005
R219 VDD2.n98 VDD2.n55 12.0247
R220 VDD2.n87 VDD2.n60 12.0247
R221 VDD2.n33 VDD2.n32 12.0247
R222 VDD2.n45 VDD2.n2 12.0247
R223 VDD2.n99 VDD2.n53 11.249
R224 VDD2.n86 VDD2.n63 11.249
R225 VDD2.n31 VDD2.n8 11.249
R226 VDD2.n46 VDD2.n0 11.249
R227 VDD2.n83 VDD2.n82 10.4732
R228 VDD2.n28 VDD2.n27 10.4732
R229 VDD2.n71 VDD2.n70 10.2747
R230 VDD2.n16 VDD2.n15 10.2747
R231 VDD2.n79 VDD2.n65 9.69747
R232 VDD2.n24 VDD2.n10 9.69747
R233 VDD2.n101 VDD2.n100 9.45567
R234 VDD2.n48 VDD2.n47 9.45567
R235 VDD2.n69 VDD2.n68 9.3005
R236 VDD2.n76 VDD2.n75 9.3005
R237 VDD2.n78 VDD2.n77 9.3005
R238 VDD2.n65 VDD2.n64 9.3005
R239 VDD2.n84 VDD2.n83 9.3005
R240 VDD2.n86 VDD2.n85 9.3005
R241 VDD2.n60 VDD2.n58 9.3005
R242 VDD2.n92 VDD2.n91 9.3005
R243 VDD2.n100 VDD2.n99 9.3005
R244 VDD2.n55 VDD2.n54 9.3005
R245 VDD2.n94 VDD2.n93 9.3005
R246 VDD2.n47 VDD2.n46 9.3005
R247 VDD2.n2 VDD2.n1 9.3005
R248 VDD2.n41 VDD2.n40 9.3005
R249 VDD2.n14 VDD2.n13 9.3005
R250 VDD2.n21 VDD2.n20 9.3005
R251 VDD2.n23 VDD2.n22 9.3005
R252 VDD2.n10 VDD2.n9 9.3005
R253 VDD2.n29 VDD2.n28 9.3005
R254 VDD2.n31 VDD2.n30 9.3005
R255 VDD2.n32 VDD2.n5 9.3005
R256 VDD2.n39 VDD2.n38 9.3005
R257 VDD2.n78 VDD2.n67 8.92171
R258 VDD2.n23 VDD2.n12 8.92171
R259 VDD2.n75 VDD2.n74 8.14595
R260 VDD2.n20 VDD2.n19 8.14595
R261 VDD2.n71 VDD2.n69 7.3702
R262 VDD2.n16 VDD2.n14 7.3702
R263 VDD2.n74 VDD2.n69 5.81868
R264 VDD2.n19 VDD2.n14 5.81868
R265 VDD2.n75 VDD2.n67 5.04292
R266 VDD2.n20 VDD2.n12 5.04292
R267 VDD2.n79 VDD2.n78 4.26717
R268 VDD2.n24 VDD2.n23 4.26717
R269 VDD2.n82 VDD2.n65 3.49141
R270 VDD2.n27 VDD2.n10 3.49141
R271 VDD2.n104 VDD2.n102 3.17291
R272 VDD2.n70 VDD2.n68 2.84303
R273 VDD2.n15 VDD2.n13 2.84303
R274 VDD2.n101 VDD2.n53 2.71565
R275 VDD2.n83 VDD2.n63 2.71565
R276 VDD2.n28 VDD2.n8 2.71565
R277 VDD2.n48 VDD2.n0 2.71565
R278 VDD2.n105 VDD2.t9 2.15034
R279 VDD2.n105 VDD2.t7 2.15034
R280 VDD2.n103 VDD2.t4 2.15034
R281 VDD2.n103 VDD2.t1 2.15034
R282 VDD2.n51 VDD2.t5 2.15034
R283 VDD2.n51 VDD2.t0 2.15034
R284 VDD2.n49 VDD2.t8 2.15034
R285 VDD2.n49 VDD2.t6 2.15034
R286 VDD2.n99 VDD2.n98 1.93989
R287 VDD2.n87 VDD2.n86 1.93989
R288 VDD2.n33 VDD2.n31 1.93989
R289 VDD2.n46 VDD2.n45 1.93989
R290 VDD2.n95 VDD2.n55 1.16414
R291 VDD2.n90 VDD2.n60 1.16414
R292 VDD2.n32 VDD2.n6 1.16414
R293 VDD2.n42 VDD2.n2 1.16414
R294 VDD2 VDD2.n104 0.851793
R295 VDD2.n52 VDD2.n50 0.738257
R296 VDD2.n94 VDD2.n57 0.388379
R297 VDD2.n91 VDD2.n59 0.388379
R298 VDD2.n38 VDD2.n37 0.388379
R299 VDD2.n41 VDD2.n4 0.388379
R300 VDD2.n100 VDD2.n54 0.155672
R301 VDD2.n93 VDD2.n54 0.155672
R302 VDD2.n93 VDD2.n92 0.155672
R303 VDD2.n92 VDD2.n58 0.155672
R304 VDD2.n85 VDD2.n58 0.155672
R305 VDD2.n85 VDD2.n84 0.155672
R306 VDD2.n84 VDD2.n64 0.155672
R307 VDD2.n77 VDD2.n64 0.155672
R308 VDD2.n77 VDD2.n76 0.155672
R309 VDD2.n76 VDD2.n68 0.155672
R310 VDD2.n21 VDD2.n13 0.155672
R311 VDD2.n22 VDD2.n21 0.155672
R312 VDD2.n22 VDD2.n9 0.155672
R313 VDD2.n29 VDD2.n9 0.155672
R314 VDD2.n30 VDD2.n29 0.155672
R315 VDD2.n30 VDD2.n5 0.155672
R316 VDD2.n39 VDD2.n5 0.155672
R317 VDD2.n40 VDD2.n39 0.155672
R318 VDD2.n40 VDD2.n1 0.155672
R319 VDD2.n47 VDD2.n1 0.155672
R320 VTAIL.n208 VTAIL.n164 289.615
R321 VTAIL.n46 VTAIL.n2 289.615
R322 VTAIL.n158 VTAIL.n114 289.615
R323 VTAIL.n104 VTAIL.n60 289.615
R324 VTAIL.n181 VTAIL.n180 185
R325 VTAIL.n183 VTAIL.n182 185
R326 VTAIL.n176 VTAIL.n175 185
R327 VTAIL.n189 VTAIL.n188 185
R328 VTAIL.n191 VTAIL.n190 185
R329 VTAIL.n172 VTAIL.n171 185
R330 VTAIL.n198 VTAIL.n197 185
R331 VTAIL.n199 VTAIL.n170 185
R332 VTAIL.n201 VTAIL.n200 185
R333 VTAIL.n168 VTAIL.n167 185
R334 VTAIL.n207 VTAIL.n206 185
R335 VTAIL.n209 VTAIL.n208 185
R336 VTAIL.n19 VTAIL.n18 185
R337 VTAIL.n21 VTAIL.n20 185
R338 VTAIL.n14 VTAIL.n13 185
R339 VTAIL.n27 VTAIL.n26 185
R340 VTAIL.n29 VTAIL.n28 185
R341 VTAIL.n10 VTAIL.n9 185
R342 VTAIL.n36 VTAIL.n35 185
R343 VTAIL.n37 VTAIL.n8 185
R344 VTAIL.n39 VTAIL.n38 185
R345 VTAIL.n6 VTAIL.n5 185
R346 VTAIL.n45 VTAIL.n44 185
R347 VTAIL.n47 VTAIL.n46 185
R348 VTAIL.n159 VTAIL.n158 185
R349 VTAIL.n157 VTAIL.n156 185
R350 VTAIL.n118 VTAIL.n117 185
R351 VTAIL.n122 VTAIL.n120 185
R352 VTAIL.n151 VTAIL.n150 185
R353 VTAIL.n149 VTAIL.n148 185
R354 VTAIL.n124 VTAIL.n123 185
R355 VTAIL.n143 VTAIL.n142 185
R356 VTAIL.n141 VTAIL.n140 185
R357 VTAIL.n128 VTAIL.n127 185
R358 VTAIL.n135 VTAIL.n134 185
R359 VTAIL.n133 VTAIL.n132 185
R360 VTAIL.n105 VTAIL.n104 185
R361 VTAIL.n103 VTAIL.n102 185
R362 VTAIL.n64 VTAIL.n63 185
R363 VTAIL.n68 VTAIL.n66 185
R364 VTAIL.n97 VTAIL.n96 185
R365 VTAIL.n95 VTAIL.n94 185
R366 VTAIL.n70 VTAIL.n69 185
R367 VTAIL.n89 VTAIL.n88 185
R368 VTAIL.n87 VTAIL.n86 185
R369 VTAIL.n74 VTAIL.n73 185
R370 VTAIL.n81 VTAIL.n80 185
R371 VTAIL.n79 VTAIL.n78 185
R372 VTAIL.n179 VTAIL.t15 149.524
R373 VTAIL.n17 VTAIL.t3 149.524
R374 VTAIL.n131 VTAIL.t0 149.524
R375 VTAIL.n77 VTAIL.t11 149.524
R376 VTAIL.n182 VTAIL.n181 104.615
R377 VTAIL.n182 VTAIL.n175 104.615
R378 VTAIL.n189 VTAIL.n175 104.615
R379 VTAIL.n190 VTAIL.n189 104.615
R380 VTAIL.n190 VTAIL.n171 104.615
R381 VTAIL.n198 VTAIL.n171 104.615
R382 VTAIL.n199 VTAIL.n198 104.615
R383 VTAIL.n200 VTAIL.n199 104.615
R384 VTAIL.n200 VTAIL.n167 104.615
R385 VTAIL.n207 VTAIL.n167 104.615
R386 VTAIL.n208 VTAIL.n207 104.615
R387 VTAIL.n20 VTAIL.n19 104.615
R388 VTAIL.n20 VTAIL.n13 104.615
R389 VTAIL.n27 VTAIL.n13 104.615
R390 VTAIL.n28 VTAIL.n27 104.615
R391 VTAIL.n28 VTAIL.n9 104.615
R392 VTAIL.n36 VTAIL.n9 104.615
R393 VTAIL.n37 VTAIL.n36 104.615
R394 VTAIL.n38 VTAIL.n37 104.615
R395 VTAIL.n38 VTAIL.n5 104.615
R396 VTAIL.n45 VTAIL.n5 104.615
R397 VTAIL.n46 VTAIL.n45 104.615
R398 VTAIL.n158 VTAIL.n157 104.615
R399 VTAIL.n157 VTAIL.n117 104.615
R400 VTAIL.n122 VTAIL.n117 104.615
R401 VTAIL.n150 VTAIL.n122 104.615
R402 VTAIL.n150 VTAIL.n149 104.615
R403 VTAIL.n149 VTAIL.n123 104.615
R404 VTAIL.n142 VTAIL.n123 104.615
R405 VTAIL.n142 VTAIL.n141 104.615
R406 VTAIL.n141 VTAIL.n127 104.615
R407 VTAIL.n134 VTAIL.n127 104.615
R408 VTAIL.n134 VTAIL.n133 104.615
R409 VTAIL.n104 VTAIL.n103 104.615
R410 VTAIL.n103 VTAIL.n63 104.615
R411 VTAIL.n68 VTAIL.n63 104.615
R412 VTAIL.n96 VTAIL.n68 104.615
R413 VTAIL.n96 VTAIL.n95 104.615
R414 VTAIL.n95 VTAIL.n69 104.615
R415 VTAIL.n88 VTAIL.n69 104.615
R416 VTAIL.n88 VTAIL.n87 104.615
R417 VTAIL.n87 VTAIL.n73 104.615
R418 VTAIL.n80 VTAIL.n73 104.615
R419 VTAIL.n80 VTAIL.n79 104.615
R420 VTAIL.n181 VTAIL.t15 52.3082
R421 VTAIL.n19 VTAIL.t3 52.3082
R422 VTAIL.n133 VTAIL.t0 52.3082
R423 VTAIL.n79 VTAIL.t11 52.3082
R424 VTAIL.n113 VTAIL.n112 45.7414
R425 VTAIL.n111 VTAIL.n110 45.7414
R426 VTAIL.n59 VTAIL.n58 45.7414
R427 VTAIL.n57 VTAIL.n56 45.7414
R428 VTAIL.n215 VTAIL.n214 45.7413
R429 VTAIL.n1 VTAIL.n0 45.7413
R430 VTAIL.n53 VTAIL.n52 45.7413
R431 VTAIL.n55 VTAIL.n54 45.7413
R432 VTAIL.n213 VTAIL.n212 31.6035
R433 VTAIL.n51 VTAIL.n50 31.6035
R434 VTAIL.n163 VTAIL.n162 31.6035
R435 VTAIL.n109 VTAIL.n108 31.6035
R436 VTAIL.n57 VTAIL.n55 26.6514
R437 VTAIL.n213 VTAIL.n163 23.4789
R438 VTAIL.n201 VTAIL.n168 13.1884
R439 VTAIL.n39 VTAIL.n6 13.1884
R440 VTAIL.n120 VTAIL.n118 13.1884
R441 VTAIL.n66 VTAIL.n64 13.1884
R442 VTAIL.n202 VTAIL.n170 12.8005
R443 VTAIL.n206 VTAIL.n205 12.8005
R444 VTAIL.n40 VTAIL.n8 12.8005
R445 VTAIL.n44 VTAIL.n43 12.8005
R446 VTAIL.n156 VTAIL.n155 12.8005
R447 VTAIL.n152 VTAIL.n151 12.8005
R448 VTAIL.n102 VTAIL.n101 12.8005
R449 VTAIL.n98 VTAIL.n97 12.8005
R450 VTAIL.n197 VTAIL.n196 12.0247
R451 VTAIL.n209 VTAIL.n166 12.0247
R452 VTAIL.n35 VTAIL.n34 12.0247
R453 VTAIL.n47 VTAIL.n4 12.0247
R454 VTAIL.n159 VTAIL.n116 12.0247
R455 VTAIL.n148 VTAIL.n121 12.0247
R456 VTAIL.n105 VTAIL.n62 12.0247
R457 VTAIL.n94 VTAIL.n67 12.0247
R458 VTAIL.n195 VTAIL.n172 11.249
R459 VTAIL.n210 VTAIL.n164 11.249
R460 VTAIL.n33 VTAIL.n10 11.249
R461 VTAIL.n48 VTAIL.n2 11.249
R462 VTAIL.n160 VTAIL.n114 11.249
R463 VTAIL.n147 VTAIL.n124 11.249
R464 VTAIL.n106 VTAIL.n60 11.249
R465 VTAIL.n93 VTAIL.n70 11.249
R466 VTAIL.n192 VTAIL.n191 10.4732
R467 VTAIL.n30 VTAIL.n29 10.4732
R468 VTAIL.n144 VTAIL.n143 10.4732
R469 VTAIL.n90 VTAIL.n89 10.4732
R470 VTAIL.n180 VTAIL.n179 10.2747
R471 VTAIL.n18 VTAIL.n17 10.2747
R472 VTAIL.n132 VTAIL.n131 10.2747
R473 VTAIL.n78 VTAIL.n77 10.2747
R474 VTAIL.n188 VTAIL.n174 9.69747
R475 VTAIL.n26 VTAIL.n12 9.69747
R476 VTAIL.n140 VTAIL.n126 9.69747
R477 VTAIL.n86 VTAIL.n72 9.69747
R478 VTAIL.n212 VTAIL.n211 9.45567
R479 VTAIL.n50 VTAIL.n49 9.45567
R480 VTAIL.n162 VTAIL.n161 9.45567
R481 VTAIL.n108 VTAIL.n107 9.45567
R482 VTAIL.n211 VTAIL.n210 9.3005
R483 VTAIL.n166 VTAIL.n165 9.3005
R484 VTAIL.n205 VTAIL.n204 9.3005
R485 VTAIL.n178 VTAIL.n177 9.3005
R486 VTAIL.n185 VTAIL.n184 9.3005
R487 VTAIL.n187 VTAIL.n186 9.3005
R488 VTAIL.n174 VTAIL.n173 9.3005
R489 VTAIL.n193 VTAIL.n192 9.3005
R490 VTAIL.n195 VTAIL.n194 9.3005
R491 VTAIL.n196 VTAIL.n169 9.3005
R492 VTAIL.n203 VTAIL.n202 9.3005
R493 VTAIL.n49 VTAIL.n48 9.3005
R494 VTAIL.n4 VTAIL.n3 9.3005
R495 VTAIL.n43 VTAIL.n42 9.3005
R496 VTAIL.n16 VTAIL.n15 9.3005
R497 VTAIL.n23 VTAIL.n22 9.3005
R498 VTAIL.n25 VTAIL.n24 9.3005
R499 VTAIL.n12 VTAIL.n11 9.3005
R500 VTAIL.n31 VTAIL.n30 9.3005
R501 VTAIL.n33 VTAIL.n32 9.3005
R502 VTAIL.n34 VTAIL.n7 9.3005
R503 VTAIL.n41 VTAIL.n40 9.3005
R504 VTAIL.n130 VTAIL.n129 9.3005
R505 VTAIL.n137 VTAIL.n136 9.3005
R506 VTAIL.n139 VTAIL.n138 9.3005
R507 VTAIL.n126 VTAIL.n125 9.3005
R508 VTAIL.n145 VTAIL.n144 9.3005
R509 VTAIL.n147 VTAIL.n146 9.3005
R510 VTAIL.n121 VTAIL.n119 9.3005
R511 VTAIL.n153 VTAIL.n152 9.3005
R512 VTAIL.n161 VTAIL.n160 9.3005
R513 VTAIL.n116 VTAIL.n115 9.3005
R514 VTAIL.n155 VTAIL.n154 9.3005
R515 VTAIL.n76 VTAIL.n75 9.3005
R516 VTAIL.n83 VTAIL.n82 9.3005
R517 VTAIL.n85 VTAIL.n84 9.3005
R518 VTAIL.n72 VTAIL.n71 9.3005
R519 VTAIL.n91 VTAIL.n90 9.3005
R520 VTAIL.n93 VTAIL.n92 9.3005
R521 VTAIL.n67 VTAIL.n65 9.3005
R522 VTAIL.n99 VTAIL.n98 9.3005
R523 VTAIL.n107 VTAIL.n106 9.3005
R524 VTAIL.n62 VTAIL.n61 9.3005
R525 VTAIL.n101 VTAIL.n100 9.3005
R526 VTAIL.n187 VTAIL.n176 8.92171
R527 VTAIL.n25 VTAIL.n14 8.92171
R528 VTAIL.n139 VTAIL.n128 8.92171
R529 VTAIL.n85 VTAIL.n74 8.92171
R530 VTAIL.n184 VTAIL.n183 8.14595
R531 VTAIL.n22 VTAIL.n21 8.14595
R532 VTAIL.n136 VTAIL.n135 8.14595
R533 VTAIL.n82 VTAIL.n81 8.14595
R534 VTAIL.n180 VTAIL.n178 7.3702
R535 VTAIL.n18 VTAIL.n16 7.3702
R536 VTAIL.n132 VTAIL.n130 7.3702
R537 VTAIL.n78 VTAIL.n76 7.3702
R538 VTAIL.n183 VTAIL.n178 5.81868
R539 VTAIL.n21 VTAIL.n16 5.81868
R540 VTAIL.n135 VTAIL.n130 5.81868
R541 VTAIL.n81 VTAIL.n76 5.81868
R542 VTAIL.n184 VTAIL.n176 5.04292
R543 VTAIL.n22 VTAIL.n14 5.04292
R544 VTAIL.n136 VTAIL.n128 5.04292
R545 VTAIL.n82 VTAIL.n74 5.04292
R546 VTAIL.n188 VTAIL.n187 4.26717
R547 VTAIL.n26 VTAIL.n25 4.26717
R548 VTAIL.n140 VTAIL.n139 4.26717
R549 VTAIL.n86 VTAIL.n85 4.26717
R550 VTAIL.n191 VTAIL.n174 3.49141
R551 VTAIL.n29 VTAIL.n12 3.49141
R552 VTAIL.n143 VTAIL.n126 3.49141
R553 VTAIL.n89 VTAIL.n72 3.49141
R554 VTAIL.n59 VTAIL.n57 3.17291
R555 VTAIL.n109 VTAIL.n59 3.17291
R556 VTAIL.n113 VTAIL.n111 3.17291
R557 VTAIL.n163 VTAIL.n113 3.17291
R558 VTAIL.n55 VTAIL.n53 3.17291
R559 VTAIL.n53 VTAIL.n51 3.17291
R560 VTAIL.n215 VTAIL.n213 3.17291
R561 VTAIL.n179 VTAIL.n177 2.84303
R562 VTAIL.n17 VTAIL.n15 2.84303
R563 VTAIL.n131 VTAIL.n129 2.84303
R564 VTAIL.n77 VTAIL.n75 2.84303
R565 VTAIL.n192 VTAIL.n172 2.71565
R566 VTAIL.n212 VTAIL.n164 2.71565
R567 VTAIL.n30 VTAIL.n10 2.71565
R568 VTAIL.n50 VTAIL.n2 2.71565
R569 VTAIL.n162 VTAIL.n114 2.71565
R570 VTAIL.n144 VTAIL.n124 2.71565
R571 VTAIL.n108 VTAIL.n60 2.71565
R572 VTAIL.n90 VTAIL.n70 2.71565
R573 VTAIL VTAIL.n1 2.438
R574 VTAIL.n214 VTAIL.t12 2.15034
R575 VTAIL.n214 VTAIL.t10 2.15034
R576 VTAIL.n0 VTAIL.t14 2.15034
R577 VTAIL.n0 VTAIL.t18 2.15034
R578 VTAIL.n52 VTAIL.t5 2.15034
R579 VTAIL.n52 VTAIL.t4 2.15034
R580 VTAIL.n54 VTAIL.t6 2.15034
R581 VTAIL.n54 VTAIL.t19 2.15034
R582 VTAIL.n112 VTAIL.t8 2.15034
R583 VTAIL.n112 VTAIL.t1 2.15034
R584 VTAIL.n110 VTAIL.t7 2.15034
R585 VTAIL.n110 VTAIL.t2 2.15034
R586 VTAIL.n58 VTAIL.t13 2.15034
R587 VTAIL.n58 VTAIL.t9 2.15034
R588 VTAIL.n56 VTAIL.t17 2.15034
R589 VTAIL.n56 VTAIL.t16 2.15034
R590 VTAIL.n111 VTAIL.n109 2.05653
R591 VTAIL.n51 VTAIL.n1 2.05653
R592 VTAIL.n197 VTAIL.n195 1.93989
R593 VTAIL.n210 VTAIL.n209 1.93989
R594 VTAIL.n35 VTAIL.n33 1.93989
R595 VTAIL.n48 VTAIL.n47 1.93989
R596 VTAIL.n160 VTAIL.n159 1.93989
R597 VTAIL.n148 VTAIL.n147 1.93989
R598 VTAIL.n106 VTAIL.n105 1.93989
R599 VTAIL.n94 VTAIL.n93 1.93989
R600 VTAIL.n196 VTAIL.n170 1.16414
R601 VTAIL.n206 VTAIL.n166 1.16414
R602 VTAIL.n34 VTAIL.n8 1.16414
R603 VTAIL.n44 VTAIL.n4 1.16414
R604 VTAIL.n156 VTAIL.n116 1.16414
R605 VTAIL.n151 VTAIL.n121 1.16414
R606 VTAIL.n102 VTAIL.n62 1.16414
R607 VTAIL.n97 VTAIL.n67 1.16414
R608 VTAIL VTAIL.n215 0.735414
R609 VTAIL.n202 VTAIL.n201 0.388379
R610 VTAIL.n205 VTAIL.n168 0.388379
R611 VTAIL.n40 VTAIL.n39 0.388379
R612 VTAIL.n43 VTAIL.n6 0.388379
R613 VTAIL.n155 VTAIL.n118 0.388379
R614 VTAIL.n152 VTAIL.n120 0.388379
R615 VTAIL.n101 VTAIL.n64 0.388379
R616 VTAIL.n98 VTAIL.n66 0.388379
R617 VTAIL.n185 VTAIL.n177 0.155672
R618 VTAIL.n186 VTAIL.n185 0.155672
R619 VTAIL.n186 VTAIL.n173 0.155672
R620 VTAIL.n193 VTAIL.n173 0.155672
R621 VTAIL.n194 VTAIL.n193 0.155672
R622 VTAIL.n194 VTAIL.n169 0.155672
R623 VTAIL.n203 VTAIL.n169 0.155672
R624 VTAIL.n204 VTAIL.n203 0.155672
R625 VTAIL.n204 VTAIL.n165 0.155672
R626 VTAIL.n211 VTAIL.n165 0.155672
R627 VTAIL.n23 VTAIL.n15 0.155672
R628 VTAIL.n24 VTAIL.n23 0.155672
R629 VTAIL.n24 VTAIL.n11 0.155672
R630 VTAIL.n31 VTAIL.n11 0.155672
R631 VTAIL.n32 VTAIL.n31 0.155672
R632 VTAIL.n32 VTAIL.n7 0.155672
R633 VTAIL.n41 VTAIL.n7 0.155672
R634 VTAIL.n42 VTAIL.n41 0.155672
R635 VTAIL.n42 VTAIL.n3 0.155672
R636 VTAIL.n49 VTAIL.n3 0.155672
R637 VTAIL.n161 VTAIL.n115 0.155672
R638 VTAIL.n154 VTAIL.n115 0.155672
R639 VTAIL.n154 VTAIL.n153 0.155672
R640 VTAIL.n153 VTAIL.n119 0.155672
R641 VTAIL.n146 VTAIL.n119 0.155672
R642 VTAIL.n146 VTAIL.n145 0.155672
R643 VTAIL.n145 VTAIL.n125 0.155672
R644 VTAIL.n138 VTAIL.n125 0.155672
R645 VTAIL.n138 VTAIL.n137 0.155672
R646 VTAIL.n137 VTAIL.n129 0.155672
R647 VTAIL.n107 VTAIL.n61 0.155672
R648 VTAIL.n100 VTAIL.n61 0.155672
R649 VTAIL.n100 VTAIL.n99 0.155672
R650 VTAIL.n99 VTAIL.n65 0.155672
R651 VTAIL.n92 VTAIL.n65 0.155672
R652 VTAIL.n92 VTAIL.n91 0.155672
R653 VTAIL.n91 VTAIL.n71 0.155672
R654 VTAIL.n84 VTAIL.n71 0.155672
R655 VTAIL.n84 VTAIL.n83 0.155672
R656 VTAIL.n83 VTAIL.n75 0.155672
R657 B.n977 B.n976 585
R658 B.n325 B.n170 585
R659 B.n324 B.n323 585
R660 B.n322 B.n321 585
R661 B.n320 B.n319 585
R662 B.n318 B.n317 585
R663 B.n316 B.n315 585
R664 B.n314 B.n313 585
R665 B.n312 B.n311 585
R666 B.n310 B.n309 585
R667 B.n308 B.n307 585
R668 B.n306 B.n305 585
R669 B.n304 B.n303 585
R670 B.n302 B.n301 585
R671 B.n300 B.n299 585
R672 B.n298 B.n297 585
R673 B.n296 B.n295 585
R674 B.n294 B.n293 585
R675 B.n292 B.n291 585
R676 B.n290 B.n289 585
R677 B.n288 B.n287 585
R678 B.n286 B.n285 585
R679 B.n284 B.n283 585
R680 B.n282 B.n281 585
R681 B.n280 B.n279 585
R682 B.n278 B.n277 585
R683 B.n276 B.n275 585
R684 B.n274 B.n273 585
R685 B.n272 B.n271 585
R686 B.n270 B.n269 585
R687 B.n268 B.n267 585
R688 B.n266 B.n265 585
R689 B.n264 B.n263 585
R690 B.n261 B.n260 585
R691 B.n259 B.n258 585
R692 B.n257 B.n256 585
R693 B.n255 B.n254 585
R694 B.n253 B.n252 585
R695 B.n251 B.n250 585
R696 B.n249 B.n248 585
R697 B.n247 B.n246 585
R698 B.n245 B.n244 585
R699 B.n243 B.n242 585
R700 B.n240 B.n239 585
R701 B.n238 B.n237 585
R702 B.n236 B.n235 585
R703 B.n234 B.n233 585
R704 B.n232 B.n231 585
R705 B.n230 B.n229 585
R706 B.n228 B.n227 585
R707 B.n226 B.n225 585
R708 B.n224 B.n223 585
R709 B.n222 B.n221 585
R710 B.n220 B.n219 585
R711 B.n218 B.n217 585
R712 B.n216 B.n215 585
R713 B.n214 B.n213 585
R714 B.n212 B.n211 585
R715 B.n210 B.n209 585
R716 B.n208 B.n207 585
R717 B.n206 B.n205 585
R718 B.n204 B.n203 585
R719 B.n202 B.n201 585
R720 B.n200 B.n199 585
R721 B.n198 B.n197 585
R722 B.n196 B.n195 585
R723 B.n194 B.n193 585
R724 B.n192 B.n191 585
R725 B.n190 B.n189 585
R726 B.n188 B.n187 585
R727 B.n186 B.n185 585
R728 B.n184 B.n183 585
R729 B.n182 B.n181 585
R730 B.n180 B.n179 585
R731 B.n178 B.n177 585
R732 B.n176 B.n175 585
R733 B.n975 B.n132 585
R734 B.n980 B.n132 585
R735 B.n974 B.n131 585
R736 B.n981 B.n131 585
R737 B.n973 B.n972 585
R738 B.n972 B.n127 585
R739 B.n971 B.n126 585
R740 B.n987 B.n126 585
R741 B.n970 B.n125 585
R742 B.n988 B.n125 585
R743 B.n969 B.n124 585
R744 B.n989 B.n124 585
R745 B.n968 B.n967 585
R746 B.n967 B.n120 585
R747 B.n966 B.n119 585
R748 B.n995 B.n119 585
R749 B.n965 B.n118 585
R750 B.n996 B.n118 585
R751 B.n964 B.n117 585
R752 B.n997 B.n117 585
R753 B.n963 B.n962 585
R754 B.n962 B.n113 585
R755 B.n961 B.n112 585
R756 B.n1003 B.n112 585
R757 B.n960 B.n111 585
R758 B.n1004 B.n111 585
R759 B.n959 B.n110 585
R760 B.n1005 B.n110 585
R761 B.n958 B.n957 585
R762 B.n957 B.n106 585
R763 B.n956 B.n105 585
R764 B.n1011 B.n105 585
R765 B.n955 B.n104 585
R766 B.n1012 B.n104 585
R767 B.n954 B.n103 585
R768 B.n1013 B.n103 585
R769 B.n953 B.n952 585
R770 B.n952 B.n99 585
R771 B.n951 B.n98 585
R772 B.n1019 B.n98 585
R773 B.n950 B.n97 585
R774 B.n1020 B.n97 585
R775 B.n949 B.n96 585
R776 B.n1021 B.n96 585
R777 B.n948 B.n947 585
R778 B.n947 B.n95 585
R779 B.n946 B.n91 585
R780 B.n1027 B.n91 585
R781 B.n945 B.n90 585
R782 B.n1028 B.n90 585
R783 B.n944 B.n89 585
R784 B.n1029 B.n89 585
R785 B.n943 B.n942 585
R786 B.n942 B.n85 585
R787 B.n941 B.n84 585
R788 B.n1035 B.n84 585
R789 B.n940 B.n83 585
R790 B.n1036 B.n83 585
R791 B.n939 B.n82 585
R792 B.n1037 B.n82 585
R793 B.n938 B.n937 585
R794 B.n937 B.n78 585
R795 B.n936 B.n77 585
R796 B.n1043 B.n77 585
R797 B.n935 B.n76 585
R798 B.n1044 B.n76 585
R799 B.n934 B.n75 585
R800 B.n1045 B.n75 585
R801 B.n933 B.n932 585
R802 B.n932 B.n71 585
R803 B.n931 B.n70 585
R804 B.n1051 B.n70 585
R805 B.n930 B.n69 585
R806 B.n1052 B.n69 585
R807 B.n929 B.n68 585
R808 B.n1053 B.n68 585
R809 B.n928 B.n927 585
R810 B.n927 B.n64 585
R811 B.n926 B.n63 585
R812 B.n1059 B.n63 585
R813 B.n925 B.n62 585
R814 B.n1060 B.n62 585
R815 B.n924 B.n61 585
R816 B.n1061 B.n61 585
R817 B.n923 B.n922 585
R818 B.n922 B.n57 585
R819 B.n921 B.n56 585
R820 B.n1067 B.n56 585
R821 B.n920 B.n55 585
R822 B.n1068 B.n55 585
R823 B.n919 B.n54 585
R824 B.n1069 B.n54 585
R825 B.n918 B.n917 585
R826 B.n917 B.n50 585
R827 B.n916 B.n49 585
R828 B.n1075 B.n49 585
R829 B.n915 B.n48 585
R830 B.n1076 B.n48 585
R831 B.n914 B.n47 585
R832 B.n1077 B.n47 585
R833 B.n913 B.n912 585
R834 B.n912 B.n43 585
R835 B.n911 B.n42 585
R836 B.n1083 B.n42 585
R837 B.n910 B.n41 585
R838 B.n1084 B.n41 585
R839 B.n909 B.n40 585
R840 B.n1085 B.n40 585
R841 B.n908 B.n907 585
R842 B.n907 B.n36 585
R843 B.n906 B.n35 585
R844 B.n1091 B.n35 585
R845 B.n905 B.n34 585
R846 B.n1092 B.n34 585
R847 B.n904 B.n33 585
R848 B.n1093 B.n33 585
R849 B.n903 B.n902 585
R850 B.n902 B.n29 585
R851 B.n901 B.n28 585
R852 B.n1099 B.n28 585
R853 B.n900 B.n27 585
R854 B.n1100 B.n27 585
R855 B.n899 B.n26 585
R856 B.n1101 B.n26 585
R857 B.n898 B.n897 585
R858 B.n897 B.n22 585
R859 B.n896 B.n21 585
R860 B.n1107 B.n21 585
R861 B.n895 B.n20 585
R862 B.n1108 B.n20 585
R863 B.n894 B.n19 585
R864 B.n1109 B.n19 585
R865 B.n893 B.n892 585
R866 B.n892 B.n15 585
R867 B.n891 B.n14 585
R868 B.n1115 B.n14 585
R869 B.n890 B.n13 585
R870 B.n1116 B.n13 585
R871 B.n889 B.n12 585
R872 B.n1117 B.n12 585
R873 B.n888 B.n887 585
R874 B.n887 B.n8 585
R875 B.n886 B.n7 585
R876 B.n1123 B.n7 585
R877 B.n885 B.n6 585
R878 B.n1124 B.n6 585
R879 B.n884 B.n5 585
R880 B.n1125 B.n5 585
R881 B.n883 B.n882 585
R882 B.n882 B.n4 585
R883 B.n881 B.n326 585
R884 B.n881 B.n880 585
R885 B.n871 B.n327 585
R886 B.n328 B.n327 585
R887 B.n873 B.n872 585
R888 B.n874 B.n873 585
R889 B.n870 B.n333 585
R890 B.n333 B.n332 585
R891 B.n869 B.n868 585
R892 B.n868 B.n867 585
R893 B.n335 B.n334 585
R894 B.n336 B.n335 585
R895 B.n860 B.n859 585
R896 B.n861 B.n860 585
R897 B.n858 B.n341 585
R898 B.n341 B.n340 585
R899 B.n857 B.n856 585
R900 B.n856 B.n855 585
R901 B.n343 B.n342 585
R902 B.n344 B.n343 585
R903 B.n848 B.n847 585
R904 B.n849 B.n848 585
R905 B.n846 B.n349 585
R906 B.n349 B.n348 585
R907 B.n845 B.n844 585
R908 B.n844 B.n843 585
R909 B.n351 B.n350 585
R910 B.n352 B.n351 585
R911 B.n836 B.n835 585
R912 B.n837 B.n836 585
R913 B.n834 B.n357 585
R914 B.n357 B.n356 585
R915 B.n833 B.n832 585
R916 B.n832 B.n831 585
R917 B.n359 B.n358 585
R918 B.n360 B.n359 585
R919 B.n824 B.n823 585
R920 B.n825 B.n824 585
R921 B.n822 B.n365 585
R922 B.n365 B.n364 585
R923 B.n821 B.n820 585
R924 B.n820 B.n819 585
R925 B.n367 B.n366 585
R926 B.n368 B.n367 585
R927 B.n812 B.n811 585
R928 B.n813 B.n812 585
R929 B.n810 B.n373 585
R930 B.n373 B.n372 585
R931 B.n809 B.n808 585
R932 B.n808 B.n807 585
R933 B.n375 B.n374 585
R934 B.n376 B.n375 585
R935 B.n800 B.n799 585
R936 B.n801 B.n800 585
R937 B.n798 B.n380 585
R938 B.n384 B.n380 585
R939 B.n797 B.n796 585
R940 B.n796 B.n795 585
R941 B.n382 B.n381 585
R942 B.n383 B.n382 585
R943 B.n788 B.n787 585
R944 B.n789 B.n788 585
R945 B.n786 B.n389 585
R946 B.n389 B.n388 585
R947 B.n785 B.n784 585
R948 B.n784 B.n783 585
R949 B.n391 B.n390 585
R950 B.n392 B.n391 585
R951 B.n776 B.n775 585
R952 B.n777 B.n776 585
R953 B.n774 B.n397 585
R954 B.n397 B.n396 585
R955 B.n773 B.n772 585
R956 B.n772 B.n771 585
R957 B.n399 B.n398 585
R958 B.n400 B.n399 585
R959 B.n764 B.n763 585
R960 B.n765 B.n764 585
R961 B.n762 B.n405 585
R962 B.n405 B.n404 585
R963 B.n761 B.n760 585
R964 B.n760 B.n759 585
R965 B.n407 B.n406 585
R966 B.n408 B.n407 585
R967 B.n752 B.n751 585
R968 B.n753 B.n752 585
R969 B.n750 B.n413 585
R970 B.n413 B.n412 585
R971 B.n749 B.n748 585
R972 B.n748 B.n747 585
R973 B.n415 B.n414 585
R974 B.n416 B.n415 585
R975 B.n740 B.n739 585
R976 B.n741 B.n740 585
R977 B.n738 B.n421 585
R978 B.n421 B.n420 585
R979 B.n737 B.n736 585
R980 B.n736 B.n735 585
R981 B.n423 B.n422 585
R982 B.n728 B.n423 585
R983 B.n727 B.n726 585
R984 B.n729 B.n727 585
R985 B.n725 B.n428 585
R986 B.n428 B.n427 585
R987 B.n724 B.n723 585
R988 B.n723 B.n722 585
R989 B.n430 B.n429 585
R990 B.n431 B.n430 585
R991 B.n715 B.n714 585
R992 B.n716 B.n715 585
R993 B.n713 B.n436 585
R994 B.n436 B.n435 585
R995 B.n712 B.n711 585
R996 B.n711 B.n710 585
R997 B.n438 B.n437 585
R998 B.n439 B.n438 585
R999 B.n703 B.n702 585
R1000 B.n704 B.n703 585
R1001 B.n701 B.n444 585
R1002 B.n444 B.n443 585
R1003 B.n700 B.n699 585
R1004 B.n699 B.n698 585
R1005 B.n446 B.n445 585
R1006 B.n447 B.n446 585
R1007 B.n691 B.n690 585
R1008 B.n692 B.n691 585
R1009 B.n689 B.n451 585
R1010 B.n455 B.n451 585
R1011 B.n688 B.n687 585
R1012 B.n687 B.n686 585
R1013 B.n453 B.n452 585
R1014 B.n454 B.n453 585
R1015 B.n679 B.n678 585
R1016 B.n680 B.n679 585
R1017 B.n677 B.n460 585
R1018 B.n460 B.n459 585
R1019 B.n676 B.n675 585
R1020 B.n675 B.n674 585
R1021 B.n462 B.n461 585
R1022 B.n463 B.n462 585
R1023 B.n667 B.n666 585
R1024 B.n668 B.n667 585
R1025 B.n665 B.n468 585
R1026 B.n468 B.n467 585
R1027 B.n660 B.n659 585
R1028 B.n658 B.n508 585
R1029 B.n657 B.n507 585
R1030 B.n662 B.n507 585
R1031 B.n656 B.n655 585
R1032 B.n654 B.n653 585
R1033 B.n652 B.n651 585
R1034 B.n650 B.n649 585
R1035 B.n648 B.n647 585
R1036 B.n646 B.n645 585
R1037 B.n644 B.n643 585
R1038 B.n642 B.n641 585
R1039 B.n640 B.n639 585
R1040 B.n638 B.n637 585
R1041 B.n636 B.n635 585
R1042 B.n634 B.n633 585
R1043 B.n632 B.n631 585
R1044 B.n630 B.n629 585
R1045 B.n628 B.n627 585
R1046 B.n626 B.n625 585
R1047 B.n624 B.n623 585
R1048 B.n622 B.n621 585
R1049 B.n620 B.n619 585
R1050 B.n618 B.n617 585
R1051 B.n616 B.n615 585
R1052 B.n614 B.n613 585
R1053 B.n612 B.n611 585
R1054 B.n610 B.n609 585
R1055 B.n608 B.n607 585
R1056 B.n606 B.n605 585
R1057 B.n604 B.n603 585
R1058 B.n602 B.n601 585
R1059 B.n600 B.n599 585
R1060 B.n598 B.n597 585
R1061 B.n596 B.n595 585
R1062 B.n594 B.n593 585
R1063 B.n592 B.n591 585
R1064 B.n590 B.n589 585
R1065 B.n588 B.n587 585
R1066 B.n586 B.n585 585
R1067 B.n584 B.n583 585
R1068 B.n582 B.n581 585
R1069 B.n580 B.n579 585
R1070 B.n578 B.n577 585
R1071 B.n576 B.n575 585
R1072 B.n574 B.n573 585
R1073 B.n572 B.n571 585
R1074 B.n570 B.n569 585
R1075 B.n568 B.n567 585
R1076 B.n566 B.n565 585
R1077 B.n564 B.n563 585
R1078 B.n562 B.n561 585
R1079 B.n560 B.n559 585
R1080 B.n558 B.n557 585
R1081 B.n556 B.n555 585
R1082 B.n554 B.n553 585
R1083 B.n552 B.n551 585
R1084 B.n550 B.n549 585
R1085 B.n548 B.n547 585
R1086 B.n546 B.n545 585
R1087 B.n544 B.n543 585
R1088 B.n542 B.n541 585
R1089 B.n540 B.n539 585
R1090 B.n538 B.n537 585
R1091 B.n536 B.n535 585
R1092 B.n534 B.n533 585
R1093 B.n532 B.n531 585
R1094 B.n530 B.n529 585
R1095 B.n528 B.n527 585
R1096 B.n526 B.n525 585
R1097 B.n524 B.n523 585
R1098 B.n522 B.n521 585
R1099 B.n520 B.n519 585
R1100 B.n518 B.n517 585
R1101 B.n516 B.n515 585
R1102 B.n470 B.n469 585
R1103 B.n664 B.n663 585
R1104 B.n663 B.n662 585
R1105 B.n466 B.n465 585
R1106 B.n467 B.n466 585
R1107 B.n670 B.n669 585
R1108 B.n669 B.n668 585
R1109 B.n671 B.n464 585
R1110 B.n464 B.n463 585
R1111 B.n673 B.n672 585
R1112 B.n674 B.n673 585
R1113 B.n458 B.n457 585
R1114 B.n459 B.n458 585
R1115 B.n682 B.n681 585
R1116 B.n681 B.n680 585
R1117 B.n683 B.n456 585
R1118 B.n456 B.n454 585
R1119 B.n685 B.n684 585
R1120 B.n686 B.n685 585
R1121 B.n450 B.n449 585
R1122 B.n455 B.n450 585
R1123 B.n694 B.n693 585
R1124 B.n693 B.n692 585
R1125 B.n695 B.n448 585
R1126 B.n448 B.n447 585
R1127 B.n697 B.n696 585
R1128 B.n698 B.n697 585
R1129 B.n442 B.n441 585
R1130 B.n443 B.n442 585
R1131 B.n706 B.n705 585
R1132 B.n705 B.n704 585
R1133 B.n707 B.n440 585
R1134 B.n440 B.n439 585
R1135 B.n709 B.n708 585
R1136 B.n710 B.n709 585
R1137 B.n434 B.n433 585
R1138 B.n435 B.n434 585
R1139 B.n718 B.n717 585
R1140 B.n717 B.n716 585
R1141 B.n719 B.n432 585
R1142 B.n432 B.n431 585
R1143 B.n721 B.n720 585
R1144 B.n722 B.n721 585
R1145 B.n426 B.n425 585
R1146 B.n427 B.n426 585
R1147 B.n731 B.n730 585
R1148 B.n730 B.n729 585
R1149 B.n732 B.n424 585
R1150 B.n728 B.n424 585
R1151 B.n734 B.n733 585
R1152 B.n735 B.n734 585
R1153 B.n419 B.n418 585
R1154 B.n420 B.n419 585
R1155 B.n743 B.n742 585
R1156 B.n742 B.n741 585
R1157 B.n744 B.n417 585
R1158 B.n417 B.n416 585
R1159 B.n746 B.n745 585
R1160 B.n747 B.n746 585
R1161 B.n411 B.n410 585
R1162 B.n412 B.n411 585
R1163 B.n755 B.n754 585
R1164 B.n754 B.n753 585
R1165 B.n756 B.n409 585
R1166 B.n409 B.n408 585
R1167 B.n758 B.n757 585
R1168 B.n759 B.n758 585
R1169 B.n403 B.n402 585
R1170 B.n404 B.n403 585
R1171 B.n767 B.n766 585
R1172 B.n766 B.n765 585
R1173 B.n768 B.n401 585
R1174 B.n401 B.n400 585
R1175 B.n770 B.n769 585
R1176 B.n771 B.n770 585
R1177 B.n395 B.n394 585
R1178 B.n396 B.n395 585
R1179 B.n779 B.n778 585
R1180 B.n778 B.n777 585
R1181 B.n780 B.n393 585
R1182 B.n393 B.n392 585
R1183 B.n782 B.n781 585
R1184 B.n783 B.n782 585
R1185 B.n387 B.n386 585
R1186 B.n388 B.n387 585
R1187 B.n791 B.n790 585
R1188 B.n790 B.n789 585
R1189 B.n792 B.n385 585
R1190 B.n385 B.n383 585
R1191 B.n794 B.n793 585
R1192 B.n795 B.n794 585
R1193 B.n379 B.n378 585
R1194 B.n384 B.n379 585
R1195 B.n803 B.n802 585
R1196 B.n802 B.n801 585
R1197 B.n804 B.n377 585
R1198 B.n377 B.n376 585
R1199 B.n806 B.n805 585
R1200 B.n807 B.n806 585
R1201 B.n371 B.n370 585
R1202 B.n372 B.n371 585
R1203 B.n815 B.n814 585
R1204 B.n814 B.n813 585
R1205 B.n816 B.n369 585
R1206 B.n369 B.n368 585
R1207 B.n818 B.n817 585
R1208 B.n819 B.n818 585
R1209 B.n363 B.n362 585
R1210 B.n364 B.n363 585
R1211 B.n827 B.n826 585
R1212 B.n826 B.n825 585
R1213 B.n828 B.n361 585
R1214 B.n361 B.n360 585
R1215 B.n830 B.n829 585
R1216 B.n831 B.n830 585
R1217 B.n355 B.n354 585
R1218 B.n356 B.n355 585
R1219 B.n839 B.n838 585
R1220 B.n838 B.n837 585
R1221 B.n840 B.n353 585
R1222 B.n353 B.n352 585
R1223 B.n842 B.n841 585
R1224 B.n843 B.n842 585
R1225 B.n347 B.n346 585
R1226 B.n348 B.n347 585
R1227 B.n851 B.n850 585
R1228 B.n850 B.n849 585
R1229 B.n852 B.n345 585
R1230 B.n345 B.n344 585
R1231 B.n854 B.n853 585
R1232 B.n855 B.n854 585
R1233 B.n339 B.n338 585
R1234 B.n340 B.n339 585
R1235 B.n863 B.n862 585
R1236 B.n862 B.n861 585
R1237 B.n864 B.n337 585
R1238 B.n337 B.n336 585
R1239 B.n866 B.n865 585
R1240 B.n867 B.n866 585
R1241 B.n331 B.n330 585
R1242 B.n332 B.n331 585
R1243 B.n876 B.n875 585
R1244 B.n875 B.n874 585
R1245 B.n877 B.n329 585
R1246 B.n329 B.n328 585
R1247 B.n879 B.n878 585
R1248 B.n880 B.n879 585
R1249 B.n2 B.n0 585
R1250 B.n4 B.n2 585
R1251 B.n3 B.n1 585
R1252 B.n1124 B.n3 585
R1253 B.n1122 B.n1121 585
R1254 B.n1123 B.n1122 585
R1255 B.n1120 B.n9 585
R1256 B.n9 B.n8 585
R1257 B.n1119 B.n1118 585
R1258 B.n1118 B.n1117 585
R1259 B.n11 B.n10 585
R1260 B.n1116 B.n11 585
R1261 B.n1114 B.n1113 585
R1262 B.n1115 B.n1114 585
R1263 B.n1112 B.n16 585
R1264 B.n16 B.n15 585
R1265 B.n1111 B.n1110 585
R1266 B.n1110 B.n1109 585
R1267 B.n18 B.n17 585
R1268 B.n1108 B.n18 585
R1269 B.n1106 B.n1105 585
R1270 B.n1107 B.n1106 585
R1271 B.n1104 B.n23 585
R1272 B.n23 B.n22 585
R1273 B.n1103 B.n1102 585
R1274 B.n1102 B.n1101 585
R1275 B.n25 B.n24 585
R1276 B.n1100 B.n25 585
R1277 B.n1098 B.n1097 585
R1278 B.n1099 B.n1098 585
R1279 B.n1096 B.n30 585
R1280 B.n30 B.n29 585
R1281 B.n1095 B.n1094 585
R1282 B.n1094 B.n1093 585
R1283 B.n32 B.n31 585
R1284 B.n1092 B.n32 585
R1285 B.n1090 B.n1089 585
R1286 B.n1091 B.n1090 585
R1287 B.n1088 B.n37 585
R1288 B.n37 B.n36 585
R1289 B.n1087 B.n1086 585
R1290 B.n1086 B.n1085 585
R1291 B.n39 B.n38 585
R1292 B.n1084 B.n39 585
R1293 B.n1082 B.n1081 585
R1294 B.n1083 B.n1082 585
R1295 B.n1080 B.n44 585
R1296 B.n44 B.n43 585
R1297 B.n1079 B.n1078 585
R1298 B.n1078 B.n1077 585
R1299 B.n46 B.n45 585
R1300 B.n1076 B.n46 585
R1301 B.n1074 B.n1073 585
R1302 B.n1075 B.n1074 585
R1303 B.n1072 B.n51 585
R1304 B.n51 B.n50 585
R1305 B.n1071 B.n1070 585
R1306 B.n1070 B.n1069 585
R1307 B.n53 B.n52 585
R1308 B.n1068 B.n53 585
R1309 B.n1066 B.n1065 585
R1310 B.n1067 B.n1066 585
R1311 B.n1064 B.n58 585
R1312 B.n58 B.n57 585
R1313 B.n1063 B.n1062 585
R1314 B.n1062 B.n1061 585
R1315 B.n60 B.n59 585
R1316 B.n1060 B.n60 585
R1317 B.n1058 B.n1057 585
R1318 B.n1059 B.n1058 585
R1319 B.n1056 B.n65 585
R1320 B.n65 B.n64 585
R1321 B.n1055 B.n1054 585
R1322 B.n1054 B.n1053 585
R1323 B.n67 B.n66 585
R1324 B.n1052 B.n67 585
R1325 B.n1050 B.n1049 585
R1326 B.n1051 B.n1050 585
R1327 B.n1048 B.n72 585
R1328 B.n72 B.n71 585
R1329 B.n1047 B.n1046 585
R1330 B.n1046 B.n1045 585
R1331 B.n74 B.n73 585
R1332 B.n1044 B.n74 585
R1333 B.n1042 B.n1041 585
R1334 B.n1043 B.n1042 585
R1335 B.n1040 B.n79 585
R1336 B.n79 B.n78 585
R1337 B.n1039 B.n1038 585
R1338 B.n1038 B.n1037 585
R1339 B.n81 B.n80 585
R1340 B.n1036 B.n81 585
R1341 B.n1034 B.n1033 585
R1342 B.n1035 B.n1034 585
R1343 B.n1032 B.n86 585
R1344 B.n86 B.n85 585
R1345 B.n1031 B.n1030 585
R1346 B.n1030 B.n1029 585
R1347 B.n88 B.n87 585
R1348 B.n1028 B.n88 585
R1349 B.n1026 B.n1025 585
R1350 B.n1027 B.n1026 585
R1351 B.n1024 B.n92 585
R1352 B.n95 B.n92 585
R1353 B.n1023 B.n1022 585
R1354 B.n1022 B.n1021 585
R1355 B.n94 B.n93 585
R1356 B.n1020 B.n94 585
R1357 B.n1018 B.n1017 585
R1358 B.n1019 B.n1018 585
R1359 B.n1016 B.n100 585
R1360 B.n100 B.n99 585
R1361 B.n1015 B.n1014 585
R1362 B.n1014 B.n1013 585
R1363 B.n102 B.n101 585
R1364 B.n1012 B.n102 585
R1365 B.n1010 B.n1009 585
R1366 B.n1011 B.n1010 585
R1367 B.n1008 B.n107 585
R1368 B.n107 B.n106 585
R1369 B.n1007 B.n1006 585
R1370 B.n1006 B.n1005 585
R1371 B.n109 B.n108 585
R1372 B.n1004 B.n109 585
R1373 B.n1002 B.n1001 585
R1374 B.n1003 B.n1002 585
R1375 B.n1000 B.n114 585
R1376 B.n114 B.n113 585
R1377 B.n999 B.n998 585
R1378 B.n998 B.n997 585
R1379 B.n116 B.n115 585
R1380 B.n996 B.n116 585
R1381 B.n994 B.n993 585
R1382 B.n995 B.n994 585
R1383 B.n992 B.n121 585
R1384 B.n121 B.n120 585
R1385 B.n991 B.n990 585
R1386 B.n990 B.n989 585
R1387 B.n123 B.n122 585
R1388 B.n988 B.n123 585
R1389 B.n986 B.n985 585
R1390 B.n987 B.n986 585
R1391 B.n984 B.n128 585
R1392 B.n128 B.n127 585
R1393 B.n983 B.n982 585
R1394 B.n982 B.n981 585
R1395 B.n130 B.n129 585
R1396 B.n980 B.n130 585
R1397 B.n1127 B.n1126 585
R1398 B.n1126 B.n1125 585
R1399 B.n660 B.n466 540.549
R1400 B.n175 B.n130 540.549
R1401 B.n663 B.n468 540.549
R1402 B.n977 B.n132 540.549
R1403 B.n512 B.t16 305.171
R1404 B.n171 B.t22 305.171
R1405 B.n509 B.t13 305.171
R1406 B.n173 B.t19 305.171
R1407 B.n512 B.t14 275.212
R1408 B.n509 B.t10 275.212
R1409 B.n173 B.t17 275.212
R1410 B.n171 B.t21 275.212
R1411 B.n979 B.n978 256.663
R1412 B.n979 B.n169 256.663
R1413 B.n979 B.n168 256.663
R1414 B.n979 B.n167 256.663
R1415 B.n979 B.n166 256.663
R1416 B.n979 B.n165 256.663
R1417 B.n979 B.n164 256.663
R1418 B.n979 B.n163 256.663
R1419 B.n979 B.n162 256.663
R1420 B.n979 B.n161 256.663
R1421 B.n979 B.n160 256.663
R1422 B.n979 B.n159 256.663
R1423 B.n979 B.n158 256.663
R1424 B.n979 B.n157 256.663
R1425 B.n979 B.n156 256.663
R1426 B.n979 B.n155 256.663
R1427 B.n979 B.n154 256.663
R1428 B.n979 B.n153 256.663
R1429 B.n979 B.n152 256.663
R1430 B.n979 B.n151 256.663
R1431 B.n979 B.n150 256.663
R1432 B.n979 B.n149 256.663
R1433 B.n979 B.n148 256.663
R1434 B.n979 B.n147 256.663
R1435 B.n979 B.n146 256.663
R1436 B.n979 B.n145 256.663
R1437 B.n979 B.n144 256.663
R1438 B.n979 B.n143 256.663
R1439 B.n979 B.n142 256.663
R1440 B.n979 B.n141 256.663
R1441 B.n979 B.n140 256.663
R1442 B.n979 B.n139 256.663
R1443 B.n979 B.n138 256.663
R1444 B.n979 B.n137 256.663
R1445 B.n979 B.n136 256.663
R1446 B.n979 B.n135 256.663
R1447 B.n979 B.n134 256.663
R1448 B.n979 B.n133 256.663
R1449 B.n662 B.n661 256.663
R1450 B.n662 B.n471 256.663
R1451 B.n662 B.n472 256.663
R1452 B.n662 B.n473 256.663
R1453 B.n662 B.n474 256.663
R1454 B.n662 B.n475 256.663
R1455 B.n662 B.n476 256.663
R1456 B.n662 B.n477 256.663
R1457 B.n662 B.n478 256.663
R1458 B.n662 B.n479 256.663
R1459 B.n662 B.n480 256.663
R1460 B.n662 B.n481 256.663
R1461 B.n662 B.n482 256.663
R1462 B.n662 B.n483 256.663
R1463 B.n662 B.n484 256.663
R1464 B.n662 B.n485 256.663
R1465 B.n662 B.n486 256.663
R1466 B.n662 B.n487 256.663
R1467 B.n662 B.n488 256.663
R1468 B.n662 B.n489 256.663
R1469 B.n662 B.n490 256.663
R1470 B.n662 B.n491 256.663
R1471 B.n662 B.n492 256.663
R1472 B.n662 B.n493 256.663
R1473 B.n662 B.n494 256.663
R1474 B.n662 B.n495 256.663
R1475 B.n662 B.n496 256.663
R1476 B.n662 B.n497 256.663
R1477 B.n662 B.n498 256.663
R1478 B.n662 B.n499 256.663
R1479 B.n662 B.n500 256.663
R1480 B.n662 B.n501 256.663
R1481 B.n662 B.n502 256.663
R1482 B.n662 B.n503 256.663
R1483 B.n662 B.n504 256.663
R1484 B.n662 B.n505 256.663
R1485 B.n662 B.n506 256.663
R1486 B.n513 B.t15 233.803
R1487 B.n172 B.t23 233.803
R1488 B.n510 B.t12 233.803
R1489 B.n174 B.t20 233.803
R1490 B.n669 B.n466 163.367
R1491 B.n669 B.n464 163.367
R1492 B.n673 B.n464 163.367
R1493 B.n673 B.n458 163.367
R1494 B.n681 B.n458 163.367
R1495 B.n681 B.n456 163.367
R1496 B.n685 B.n456 163.367
R1497 B.n685 B.n450 163.367
R1498 B.n693 B.n450 163.367
R1499 B.n693 B.n448 163.367
R1500 B.n697 B.n448 163.367
R1501 B.n697 B.n442 163.367
R1502 B.n705 B.n442 163.367
R1503 B.n705 B.n440 163.367
R1504 B.n709 B.n440 163.367
R1505 B.n709 B.n434 163.367
R1506 B.n717 B.n434 163.367
R1507 B.n717 B.n432 163.367
R1508 B.n721 B.n432 163.367
R1509 B.n721 B.n426 163.367
R1510 B.n730 B.n426 163.367
R1511 B.n730 B.n424 163.367
R1512 B.n734 B.n424 163.367
R1513 B.n734 B.n419 163.367
R1514 B.n742 B.n419 163.367
R1515 B.n742 B.n417 163.367
R1516 B.n746 B.n417 163.367
R1517 B.n746 B.n411 163.367
R1518 B.n754 B.n411 163.367
R1519 B.n754 B.n409 163.367
R1520 B.n758 B.n409 163.367
R1521 B.n758 B.n403 163.367
R1522 B.n766 B.n403 163.367
R1523 B.n766 B.n401 163.367
R1524 B.n770 B.n401 163.367
R1525 B.n770 B.n395 163.367
R1526 B.n778 B.n395 163.367
R1527 B.n778 B.n393 163.367
R1528 B.n782 B.n393 163.367
R1529 B.n782 B.n387 163.367
R1530 B.n790 B.n387 163.367
R1531 B.n790 B.n385 163.367
R1532 B.n794 B.n385 163.367
R1533 B.n794 B.n379 163.367
R1534 B.n802 B.n379 163.367
R1535 B.n802 B.n377 163.367
R1536 B.n806 B.n377 163.367
R1537 B.n806 B.n371 163.367
R1538 B.n814 B.n371 163.367
R1539 B.n814 B.n369 163.367
R1540 B.n818 B.n369 163.367
R1541 B.n818 B.n363 163.367
R1542 B.n826 B.n363 163.367
R1543 B.n826 B.n361 163.367
R1544 B.n830 B.n361 163.367
R1545 B.n830 B.n355 163.367
R1546 B.n838 B.n355 163.367
R1547 B.n838 B.n353 163.367
R1548 B.n842 B.n353 163.367
R1549 B.n842 B.n347 163.367
R1550 B.n850 B.n347 163.367
R1551 B.n850 B.n345 163.367
R1552 B.n854 B.n345 163.367
R1553 B.n854 B.n339 163.367
R1554 B.n862 B.n339 163.367
R1555 B.n862 B.n337 163.367
R1556 B.n866 B.n337 163.367
R1557 B.n866 B.n331 163.367
R1558 B.n875 B.n331 163.367
R1559 B.n875 B.n329 163.367
R1560 B.n879 B.n329 163.367
R1561 B.n879 B.n2 163.367
R1562 B.n1126 B.n2 163.367
R1563 B.n1126 B.n3 163.367
R1564 B.n1122 B.n3 163.367
R1565 B.n1122 B.n9 163.367
R1566 B.n1118 B.n9 163.367
R1567 B.n1118 B.n11 163.367
R1568 B.n1114 B.n11 163.367
R1569 B.n1114 B.n16 163.367
R1570 B.n1110 B.n16 163.367
R1571 B.n1110 B.n18 163.367
R1572 B.n1106 B.n18 163.367
R1573 B.n1106 B.n23 163.367
R1574 B.n1102 B.n23 163.367
R1575 B.n1102 B.n25 163.367
R1576 B.n1098 B.n25 163.367
R1577 B.n1098 B.n30 163.367
R1578 B.n1094 B.n30 163.367
R1579 B.n1094 B.n32 163.367
R1580 B.n1090 B.n32 163.367
R1581 B.n1090 B.n37 163.367
R1582 B.n1086 B.n37 163.367
R1583 B.n1086 B.n39 163.367
R1584 B.n1082 B.n39 163.367
R1585 B.n1082 B.n44 163.367
R1586 B.n1078 B.n44 163.367
R1587 B.n1078 B.n46 163.367
R1588 B.n1074 B.n46 163.367
R1589 B.n1074 B.n51 163.367
R1590 B.n1070 B.n51 163.367
R1591 B.n1070 B.n53 163.367
R1592 B.n1066 B.n53 163.367
R1593 B.n1066 B.n58 163.367
R1594 B.n1062 B.n58 163.367
R1595 B.n1062 B.n60 163.367
R1596 B.n1058 B.n60 163.367
R1597 B.n1058 B.n65 163.367
R1598 B.n1054 B.n65 163.367
R1599 B.n1054 B.n67 163.367
R1600 B.n1050 B.n67 163.367
R1601 B.n1050 B.n72 163.367
R1602 B.n1046 B.n72 163.367
R1603 B.n1046 B.n74 163.367
R1604 B.n1042 B.n74 163.367
R1605 B.n1042 B.n79 163.367
R1606 B.n1038 B.n79 163.367
R1607 B.n1038 B.n81 163.367
R1608 B.n1034 B.n81 163.367
R1609 B.n1034 B.n86 163.367
R1610 B.n1030 B.n86 163.367
R1611 B.n1030 B.n88 163.367
R1612 B.n1026 B.n88 163.367
R1613 B.n1026 B.n92 163.367
R1614 B.n1022 B.n92 163.367
R1615 B.n1022 B.n94 163.367
R1616 B.n1018 B.n94 163.367
R1617 B.n1018 B.n100 163.367
R1618 B.n1014 B.n100 163.367
R1619 B.n1014 B.n102 163.367
R1620 B.n1010 B.n102 163.367
R1621 B.n1010 B.n107 163.367
R1622 B.n1006 B.n107 163.367
R1623 B.n1006 B.n109 163.367
R1624 B.n1002 B.n109 163.367
R1625 B.n1002 B.n114 163.367
R1626 B.n998 B.n114 163.367
R1627 B.n998 B.n116 163.367
R1628 B.n994 B.n116 163.367
R1629 B.n994 B.n121 163.367
R1630 B.n990 B.n121 163.367
R1631 B.n990 B.n123 163.367
R1632 B.n986 B.n123 163.367
R1633 B.n986 B.n128 163.367
R1634 B.n982 B.n128 163.367
R1635 B.n982 B.n130 163.367
R1636 B.n508 B.n507 163.367
R1637 B.n655 B.n507 163.367
R1638 B.n653 B.n652 163.367
R1639 B.n649 B.n648 163.367
R1640 B.n645 B.n644 163.367
R1641 B.n641 B.n640 163.367
R1642 B.n637 B.n636 163.367
R1643 B.n633 B.n632 163.367
R1644 B.n629 B.n628 163.367
R1645 B.n625 B.n624 163.367
R1646 B.n621 B.n620 163.367
R1647 B.n617 B.n616 163.367
R1648 B.n613 B.n612 163.367
R1649 B.n609 B.n608 163.367
R1650 B.n605 B.n604 163.367
R1651 B.n601 B.n600 163.367
R1652 B.n597 B.n596 163.367
R1653 B.n593 B.n592 163.367
R1654 B.n589 B.n588 163.367
R1655 B.n585 B.n584 163.367
R1656 B.n581 B.n580 163.367
R1657 B.n577 B.n576 163.367
R1658 B.n573 B.n572 163.367
R1659 B.n569 B.n568 163.367
R1660 B.n565 B.n564 163.367
R1661 B.n561 B.n560 163.367
R1662 B.n557 B.n556 163.367
R1663 B.n553 B.n552 163.367
R1664 B.n549 B.n548 163.367
R1665 B.n545 B.n544 163.367
R1666 B.n541 B.n540 163.367
R1667 B.n537 B.n536 163.367
R1668 B.n533 B.n532 163.367
R1669 B.n529 B.n528 163.367
R1670 B.n525 B.n524 163.367
R1671 B.n521 B.n520 163.367
R1672 B.n517 B.n516 163.367
R1673 B.n663 B.n470 163.367
R1674 B.n667 B.n468 163.367
R1675 B.n667 B.n462 163.367
R1676 B.n675 B.n462 163.367
R1677 B.n675 B.n460 163.367
R1678 B.n679 B.n460 163.367
R1679 B.n679 B.n453 163.367
R1680 B.n687 B.n453 163.367
R1681 B.n687 B.n451 163.367
R1682 B.n691 B.n451 163.367
R1683 B.n691 B.n446 163.367
R1684 B.n699 B.n446 163.367
R1685 B.n699 B.n444 163.367
R1686 B.n703 B.n444 163.367
R1687 B.n703 B.n438 163.367
R1688 B.n711 B.n438 163.367
R1689 B.n711 B.n436 163.367
R1690 B.n715 B.n436 163.367
R1691 B.n715 B.n430 163.367
R1692 B.n723 B.n430 163.367
R1693 B.n723 B.n428 163.367
R1694 B.n727 B.n428 163.367
R1695 B.n727 B.n423 163.367
R1696 B.n736 B.n423 163.367
R1697 B.n736 B.n421 163.367
R1698 B.n740 B.n421 163.367
R1699 B.n740 B.n415 163.367
R1700 B.n748 B.n415 163.367
R1701 B.n748 B.n413 163.367
R1702 B.n752 B.n413 163.367
R1703 B.n752 B.n407 163.367
R1704 B.n760 B.n407 163.367
R1705 B.n760 B.n405 163.367
R1706 B.n764 B.n405 163.367
R1707 B.n764 B.n399 163.367
R1708 B.n772 B.n399 163.367
R1709 B.n772 B.n397 163.367
R1710 B.n776 B.n397 163.367
R1711 B.n776 B.n391 163.367
R1712 B.n784 B.n391 163.367
R1713 B.n784 B.n389 163.367
R1714 B.n788 B.n389 163.367
R1715 B.n788 B.n382 163.367
R1716 B.n796 B.n382 163.367
R1717 B.n796 B.n380 163.367
R1718 B.n800 B.n380 163.367
R1719 B.n800 B.n375 163.367
R1720 B.n808 B.n375 163.367
R1721 B.n808 B.n373 163.367
R1722 B.n812 B.n373 163.367
R1723 B.n812 B.n367 163.367
R1724 B.n820 B.n367 163.367
R1725 B.n820 B.n365 163.367
R1726 B.n824 B.n365 163.367
R1727 B.n824 B.n359 163.367
R1728 B.n832 B.n359 163.367
R1729 B.n832 B.n357 163.367
R1730 B.n836 B.n357 163.367
R1731 B.n836 B.n351 163.367
R1732 B.n844 B.n351 163.367
R1733 B.n844 B.n349 163.367
R1734 B.n848 B.n349 163.367
R1735 B.n848 B.n343 163.367
R1736 B.n856 B.n343 163.367
R1737 B.n856 B.n341 163.367
R1738 B.n860 B.n341 163.367
R1739 B.n860 B.n335 163.367
R1740 B.n868 B.n335 163.367
R1741 B.n868 B.n333 163.367
R1742 B.n873 B.n333 163.367
R1743 B.n873 B.n327 163.367
R1744 B.n881 B.n327 163.367
R1745 B.n882 B.n881 163.367
R1746 B.n882 B.n5 163.367
R1747 B.n6 B.n5 163.367
R1748 B.n7 B.n6 163.367
R1749 B.n887 B.n7 163.367
R1750 B.n887 B.n12 163.367
R1751 B.n13 B.n12 163.367
R1752 B.n14 B.n13 163.367
R1753 B.n892 B.n14 163.367
R1754 B.n892 B.n19 163.367
R1755 B.n20 B.n19 163.367
R1756 B.n21 B.n20 163.367
R1757 B.n897 B.n21 163.367
R1758 B.n897 B.n26 163.367
R1759 B.n27 B.n26 163.367
R1760 B.n28 B.n27 163.367
R1761 B.n902 B.n28 163.367
R1762 B.n902 B.n33 163.367
R1763 B.n34 B.n33 163.367
R1764 B.n35 B.n34 163.367
R1765 B.n907 B.n35 163.367
R1766 B.n907 B.n40 163.367
R1767 B.n41 B.n40 163.367
R1768 B.n42 B.n41 163.367
R1769 B.n912 B.n42 163.367
R1770 B.n912 B.n47 163.367
R1771 B.n48 B.n47 163.367
R1772 B.n49 B.n48 163.367
R1773 B.n917 B.n49 163.367
R1774 B.n917 B.n54 163.367
R1775 B.n55 B.n54 163.367
R1776 B.n56 B.n55 163.367
R1777 B.n922 B.n56 163.367
R1778 B.n922 B.n61 163.367
R1779 B.n62 B.n61 163.367
R1780 B.n63 B.n62 163.367
R1781 B.n927 B.n63 163.367
R1782 B.n927 B.n68 163.367
R1783 B.n69 B.n68 163.367
R1784 B.n70 B.n69 163.367
R1785 B.n932 B.n70 163.367
R1786 B.n932 B.n75 163.367
R1787 B.n76 B.n75 163.367
R1788 B.n77 B.n76 163.367
R1789 B.n937 B.n77 163.367
R1790 B.n937 B.n82 163.367
R1791 B.n83 B.n82 163.367
R1792 B.n84 B.n83 163.367
R1793 B.n942 B.n84 163.367
R1794 B.n942 B.n89 163.367
R1795 B.n90 B.n89 163.367
R1796 B.n91 B.n90 163.367
R1797 B.n947 B.n91 163.367
R1798 B.n947 B.n96 163.367
R1799 B.n97 B.n96 163.367
R1800 B.n98 B.n97 163.367
R1801 B.n952 B.n98 163.367
R1802 B.n952 B.n103 163.367
R1803 B.n104 B.n103 163.367
R1804 B.n105 B.n104 163.367
R1805 B.n957 B.n105 163.367
R1806 B.n957 B.n110 163.367
R1807 B.n111 B.n110 163.367
R1808 B.n112 B.n111 163.367
R1809 B.n962 B.n112 163.367
R1810 B.n962 B.n117 163.367
R1811 B.n118 B.n117 163.367
R1812 B.n119 B.n118 163.367
R1813 B.n967 B.n119 163.367
R1814 B.n967 B.n124 163.367
R1815 B.n125 B.n124 163.367
R1816 B.n126 B.n125 163.367
R1817 B.n972 B.n126 163.367
R1818 B.n972 B.n131 163.367
R1819 B.n132 B.n131 163.367
R1820 B.n179 B.n178 163.367
R1821 B.n183 B.n182 163.367
R1822 B.n187 B.n186 163.367
R1823 B.n191 B.n190 163.367
R1824 B.n195 B.n194 163.367
R1825 B.n199 B.n198 163.367
R1826 B.n203 B.n202 163.367
R1827 B.n207 B.n206 163.367
R1828 B.n211 B.n210 163.367
R1829 B.n215 B.n214 163.367
R1830 B.n219 B.n218 163.367
R1831 B.n223 B.n222 163.367
R1832 B.n227 B.n226 163.367
R1833 B.n231 B.n230 163.367
R1834 B.n235 B.n234 163.367
R1835 B.n239 B.n238 163.367
R1836 B.n244 B.n243 163.367
R1837 B.n248 B.n247 163.367
R1838 B.n252 B.n251 163.367
R1839 B.n256 B.n255 163.367
R1840 B.n260 B.n259 163.367
R1841 B.n265 B.n264 163.367
R1842 B.n269 B.n268 163.367
R1843 B.n273 B.n272 163.367
R1844 B.n277 B.n276 163.367
R1845 B.n281 B.n280 163.367
R1846 B.n285 B.n284 163.367
R1847 B.n289 B.n288 163.367
R1848 B.n293 B.n292 163.367
R1849 B.n297 B.n296 163.367
R1850 B.n301 B.n300 163.367
R1851 B.n305 B.n304 163.367
R1852 B.n309 B.n308 163.367
R1853 B.n313 B.n312 163.367
R1854 B.n317 B.n316 163.367
R1855 B.n321 B.n320 163.367
R1856 B.n323 B.n170 163.367
R1857 B.n662 B.n467 96.4451
R1858 B.n980 B.n979 96.4451
R1859 B.n661 B.n660 71.676
R1860 B.n655 B.n471 71.676
R1861 B.n652 B.n472 71.676
R1862 B.n648 B.n473 71.676
R1863 B.n644 B.n474 71.676
R1864 B.n640 B.n475 71.676
R1865 B.n636 B.n476 71.676
R1866 B.n632 B.n477 71.676
R1867 B.n628 B.n478 71.676
R1868 B.n624 B.n479 71.676
R1869 B.n620 B.n480 71.676
R1870 B.n616 B.n481 71.676
R1871 B.n612 B.n482 71.676
R1872 B.n608 B.n483 71.676
R1873 B.n604 B.n484 71.676
R1874 B.n600 B.n485 71.676
R1875 B.n596 B.n486 71.676
R1876 B.n592 B.n487 71.676
R1877 B.n588 B.n488 71.676
R1878 B.n584 B.n489 71.676
R1879 B.n580 B.n490 71.676
R1880 B.n576 B.n491 71.676
R1881 B.n572 B.n492 71.676
R1882 B.n568 B.n493 71.676
R1883 B.n564 B.n494 71.676
R1884 B.n560 B.n495 71.676
R1885 B.n556 B.n496 71.676
R1886 B.n552 B.n497 71.676
R1887 B.n548 B.n498 71.676
R1888 B.n544 B.n499 71.676
R1889 B.n540 B.n500 71.676
R1890 B.n536 B.n501 71.676
R1891 B.n532 B.n502 71.676
R1892 B.n528 B.n503 71.676
R1893 B.n524 B.n504 71.676
R1894 B.n520 B.n505 71.676
R1895 B.n516 B.n506 71.676
R1896 B.n175 B.n133 71.676
R1897 B.n179 B.n134 71.676
R1898 B.n183 B.n135 71.676
R1899 B.n187 B.n136 71.676
R1900 B.n191 B.n137 71.676
R1901 B.n195 B.n138 71.676
R1902 B.n199 B.n139 71.676
R1903 B.n203 B.n140 71.676
R1904 B.n207 B.n141 71.676
R1905 B.n211 B.n142 71.676
R1906 B.n215 B.n143 71.676
R1907 B.n219 B.n144 71.676
R1908 B.n223 B.n145 71.676
R1909 B.n227 B.n146 71.676
R1910 B.n231 B.n147 71.676
R1911 B.n235 B.n148 71.676
R1912 B.n239 B.n149 71.676
R1913 B.n244 B.n150 71.676
R1914 B.n248 B.n151 71.676
R1915 B.n252 B.n152 71.676
R1916 B.n256 B.n153 71.676
R1917 B.n260 B.n154 71.676
R1918 B.n265 B.n155 71.676
R1919 B.n269 B.n156 71.676
R1920 B.n273 B.n157 71.676
R1921 B.n277 B.n158 71.676
R1922 B.n281 B.n159 71.676
R1923 B.n285 B.n160 71.676
R1924 B.n289 B.n161 71.676
R1925 B.n293 B.n162 71.676
R1926 B.n297 B.n163 71.676
R1927 B.n301 B.n164 71.676
R1928 B.n305 B.n165 71.676
R1929 B.n309 B.n166 71.676
R1930 B.n313 B.n167 71.676
R1931 B.n317 B.n168 71.676
R1932 B.n321 B.n169 71.676
R1933 B.n978 B.n170 71.676
R1934 B.n978 B.n977 71.676
R1935 B.n323 B.n169 71.676
R1936 B.n320 B.n168 71.676
R1937 B.n316 B.n167 71.676
R1938 B.n312 B.n166 71.676
R1939 B.n308 B.n165 71.676
R1940 B.n304 B.n164 71.676
R1941 B.n300 B.n163 71.676
R1942 B.n296 B.n162 71.676
R1943 B.n292 B.n161 71.676
R1944 B.n288 B.n160 71.676
R1945 B.n284 B.n159 71.676
R1946 B.n280 B.n158 71.676
R1947 B.n276 B.n157 71.676
R1948 B.n272 B.n156 71.676
R1949 B.n268 B.n155 71.676
R1950 B.n264 B.n154 71.676
R1951 B.n259 B.n153 71.676
R1952 B.n255 B.n152 71.676
R1953 B.n251 B.n151 71.676
R1954 B.n247 B.n150 71.676
R1955 B.n243 B.n149 71.676
R1956 B.n238 B.n148 71.676
R1957 B.n234 B.n147 71.676
R1958 B.n230 B.n146 71.676
R1959 B.n226 B.n145 71.676
R1960 B.n222 B.n144 71.676
R1961 B.n218 B.n143 71.676
R1962 B.n214 B.n142 71.676
R1963 B.n210 B.n141 71.676
R1964 B.n206 B.n140 71.676
R1965 B.n202 B.n139 71.676
R1966 B.n198 B.n138 71.676
R1967 B.n194 B.n137 71.676
R1968 B.n190 B.n136 71.676
R1969 B.n186 B.n135 71.676
R1970 B.n182 B.n134 71.676
R1971 B.n178 B.n133 71.676
R1972 B.n661 B.n508 71.676
R1973 B.n653 B.n471 71.676
R1974 B.n649 B.n472 71.676
R1975 B.n645 B.n473 71.676
R1976 B.n641 B.n474 71.676
R1977 B.n637 B.n475 71.676
R1978 B.n633 B.n476 71.676
R1979 B.n629 B.n477 71.676
R1980 B.n625 B.n478 71.676
R1981 B.n621 B.n479 71.676
R1982 B.n617 B.n480 71.676
R1983 B.n613 B.n481 71.676
R1984 B.n609 B.n482 71.676
R1985 B.n605 B.n483 71.676
R1986 B.n601 B.n484 71.676
R1987 B.n597 B.n485 71.676
R1988 B.n593 B.n486 71.676
R1989 B.n589 B.n487 71.676
R1990 B.n585 B.n488 71.676
R1991 B.n581 B.n489 71.676
R1992 B.n577 B.n490 71.676
R1993 B.n573 B.n491 71.676
R1994 B.n569 B.n492 71.676
R1995 B.n565 B.n493 71.676
R1996 B.n561 B.n494 71.676
R1997 B.n557 B.n495 71.676
R1998 B.n553 B.n496 71.676
R1999 B.n549 B.n497 71.676
R2000 B.n545 B.n498 71.676
R2001 B.n541 B.n499 71.676
R2002 B.n537 B.n500 71.676
R2003 B.n533 B.n501 71.676
R2004 B.n529 B.n502 71.676
R2005 B.n525 B.n503 71.676
R2006 B.n521 B.n504 71.676
R2007 B.n517 B.n505 71.676
R2008 B.n506 B.n470 71.676
R2009 B.n513 B.n512 71.3702
R2010 B.n510 B.n509 71.3702
R2011 B.n174 B.n173 71.3702
R2012 B.n172 B.n171 71.3702
R2013 B.n514 B.n513 59.5399
R2014 B.n511 B.n510 59.5399
R2015 B.n241 B.n174 59.5399
R2016 B.n262 B.n172 59.5399
R2017 B.n668 B.n467 51.6401
R2018 B.n668 B.n463 51.6401
R2019 B.n674 B.n463 51.6401
R2020 B.n674 B.n459 51.6401
R2021 B.n680 B.n459 51.6401
R2022 B.n680 B.n454 51.6401
R2023 B.n686 B.n454 51.6401
R2024 B.n686 B.n455 51.6401
R2025 B.n692 B.n447 51.6401
R2026 B.n698 B.n447 51.6401
R2027 B.n698 B.n443 51.6401
R2028 B.n704 B.n443 51.6401
R2029 B.n704 B.n439 51.6401
R2030 B.n710 B.n439 51.6401
R2031 B.n710 B.n435 51.6401
R2032 B.n716 B.n435 51.6401
R2033 B.n716 B.n431 51.6401
R2034 B.n722 B.n431 51.6401
R2035 B.n722 B.n427 51.6401
R2036 B.n729 B.n427 51.6401
R2037 B.n729 B.n728 51.6401
R2038 B.n735 B.n420 51.6401
R2039 B.n741 B.n420 51.6401
R2040 B.n741 B.n416 51.6401
R2041 B.n747 B.n416 51.6401
R2042 B.n747 B.n412 51.6401
R2043 B.n753 B.n412 51.6401
R2044 B.n753 B.n408 51.6401
R2045 B.n759 B.n408 51.6401
R2046 B.n759 B.n404 51.6401
R2047 B.n765 B.n404 51.6401
R2048 B.n771 B.n400 51.6401
R2049 B.n771 B.n396 51.6401
R2050 B.n777 B.n396 51.6401
R2051 B.n777 B.n392 51.6401
R2052 B.n783 B.n392 51.6401
R2053 B.n783 B.n388 51.6401
R2054 B.n789 B.n388 51.6401
R2055 B.n789 B.n383 51.6401
R2056 B.n795 B.n383 51.6401
R2057 B.n795 B.n384 51.6401
R2058 B.n801 B.n376 51.6401
R2059 B.n807 B.n376 51.6401
R2060 B.n807 B.n372 51.6401
R2061 B.n813 B.n372 51.6401
R2062 B.n813 B.n368 51.6401
R2063 B.n819 B.n368 51.6401
R2064 B.n819 B.n364 51.6401
R2065 B.n825 B.n364 51.6401
R2066 B.n825 B.n360 51.6401
R2067 B.n831 B.n360 51.6401
R2068 B.n837 B.n356 51.6401
R2069 B.n837 B.n352 51.6401
R2070 B.n843 B.n352 51.6401
R2071 B.n843 B.n348 51.6401
R2072 B.n849 B.n348 51.6401
R2073 B.n849 B.n344 51.6401
R2074 B.n855 B.n344 51.6401
R2075 B.n855 B.n340 51.6401
R2076 B.n861 B.n340 51.6401
R2077 B.n867 B.n336 51.6401
R2078 B.n867 B.n332 51.6401
R2079 B.n874 B.n332 51.6401
R2080 B.n874 B.n328 51.6401
R2081 B.n880 B.n328 51.6401
R2082 B.n880 B.n4 51.6401
R2083 B.n1125 B.n4 51.6401
R2084 B.n1125 B.n1124 51.6401
R2085 B.n1124 B.n1123 51.6401
R2086 B.n1123 B.n8 51.6401
R2087 B.n1117 B.n8 51.6401
R2088 B.n1117 B.n1116 51.6401
R2089 B.n1116 B.n1115 51.6401
R2090 B.n1115 B.n15 51.6401
R2091 B.n1109 B.n1108 51.6401
R2092 B.n1108 B.n1107 51.6401
R2093 B.n1107 B.n22 51.6401
R2094 B.n1101 B.n22 51.6401
R2095 B.n1101 B.n1100 51.6401
R2096 B.n1100 B.n1099 51.6401
R2097 B.n1099 B.n29 51.6401
R2098 B.n1093 B.n29 51.6401
R2099 B.n1093 B.n1092 51.6401
R2100 B.n1091 B.n36 51.6401
R2101 B.n1085 B.n36 51.6401
R2102 B.n1085 B.n1084 51.6401
R2103 B.n1084 B.n1083 51.6401
R2104 B.n1083 B.n43 51.6401
R2105 B.n1077 B.n43 51.6401
R2106 B.n1077 B.n1076 51.6401
R2107 B.n1076 B.n1075 51.6401
R2108 B.n1075 B.n50 51.6401
R2109 B.n1069 B.n50 51.6401
R2110 B.n1068 B.n1067 51.6401
R2111 B.n1067 B.n57 51.6401
R2112 B.n1061 B.n57 51.6401
R2113 B.n1061 B.n1060 51.6401
R2114 B.n1060 B.n1059 51.6401
R2115 B.n1059 B.n64 51.6401
R2116 B.n1053 B.n64 51.6401
R2117 B.n1053 B.n1052 51.6401
R2118 B.n1052 B.n1051 51.6401
R2119 B.n1051 B.n71 51.6401
R2120 B.n1045 B.n1044 51.6401
R2121 B.n1044 B.n1043 51.6401
R2122 B.n1043 B.n78 51.6401
R2123 B.n1037 B.n78 51.6401
R2124 B.n1037 B.n1036 51.6401
R2125 B.n1036 B.n1035 51.6401
R2126 B.n1035 B.n85 51.6401
R2127 B.n1029 B.n85 51.6401
R2128 B.n1029 B.n1028 51.6401
R2129 B.n1028 B.n1027 51.6401
R2130 B.n1021 B.n95 51.6401
R2131 B.n1021 B.n1020 51.6401
R2132 B.n1020 B.n1019 51.6401
R2133 B.n1019 B.n99 51.6401
R2134 B.n1013 B.n99 51.6401
R2135 B.n1013 B.n1012 51.6401
R2136 B.n1012 B.n1011 51.6401
R2137 B.n1011 B.n106 51.6401
R2138 B.n1005 B.n106 51.6401
R2139 B.n1005 B.n1004 51.6401
R2140 B.n1004 B.n1003 51.6401
R2141 B.n1003 B.n113 51.6401
R2142 B.n997 B.n113 51.6401
R2143 B.n996 B.n995 51.6401
R2144 B.n995 B.n120 51.6401
R2145 B.n989 B.n120 51.6401
R2146 B.n989 B.n988 51.6401
R2147 B.n988 B.n987 51.6401
R2148 B.n987 B.n127 51.6401
R2149 B.n981 B.n127 51.6401
R2150 B.n981 B.n980 51.6401
R2151 B.n861 B.t3 50.8807
R2152 B.n1109 B.t7 50.8807
R2153 B.t4 B.n356 43.2867
R2154 B.n1092 B.t2 43.2867
R2155 B.n728 B.t6 35.6926
R2156 B.n95 B.t0 35.6926
R2157 B.n176 B.n129 35.1225
R2158 B.n976 B.n975 35.1225
R2159 B.n665 B.n664 35.1225
R2160 B.n659 B.n465 35.1225
R2161 B.n455 B.t11 34.1738
R2162 B.n801 B.t5 34.1738
R2163 B.n1069 B.t8 34.1738
R2164 B.t18 B.n996 34.1738
R2165 B.n765 B.t9 26.5797
R2166 B.n1045 B.t1 26.5797
R2167 B.t9 B.n400 25.0609
R2168 B.t1 B.n71 25.0609
R2169 B B.n1127 18.0485
R2170 B.n692 B.t11 17.4668
R2171 B.n384 B.t5 17.4668
R2172 B.t8 B.n1068 17.4668
R2173 B.n997 B.t18 17.4668
R2174 B.n735 B.t6 15.948
R2175 B.n1027 B.t0 15.948
R2176 B.n177 B.n176 10.6151
R2177 B.n180 B.n177 10.6151
R2178 B.n181 B.n180 10.6151
R2179 B.n184 B.n181 10.6151
R2180 B.n185 B.n184 10.6151
R2181 B.n188 B.n185 10.6151
R2182 B.n189 B.n188 10.6151
R2183 B.n192 B.n189 10.6151
R2184 B.n193 B.n192 10.6151
R2185 B.n196 B.n193 10.6151
R2186 B.n197 B.n196 10.6151
R2187 B.n200 B.n197 10.6151
R2188 B.n201 B.n200 10.6151
R2189 B.n204 B.n201 10.6151
R2190 B.n205 B.n204 10.6151
R2191 B.n208 B.n205 10.6151
R2192 B.n209 B.n208 10.6151
R2193 B.n212 B.n209 10.6151
R2194 B.n213 B.n212 10.6151
R2195 B.n216 B.n213 10.6151
R2196 B.n217 B.n216 10.6151
R2197 B.n220 B.n217 10.6151
R2198 B.n221 B.n220 10.6151
R2199 B.n224 B.n221 10.6151
R2200 B.n225 B.n224 10.6151
R2201 B.n228 B.n225 10.6151
R2202 B.n229 B.n228 10.6151
R2203 B.n232 B.n229 10.6151
R2204 B.n233 B.n232 10.6151
R2205 B.n236 B.n233 10.6151
R2206 B.n237 B.n236 10.6151
R2207 B.n240 B.n237 10.6151
R2208 B.n245 B.n242 10.6151
R2209 B.n246 B.n245 10.6151
R2210 B.n249 B.n246 10.6151
R2211 B.n250 B.n249 10.6151
R2212 B.n253 B.n250 10.6151
R2213 B.n254 B.n253 10.6151
R2214 B.n257 B.n254 10.6151
R2215 B.n258 B.n257 10.6151
R2216 B.n261 B.n258 10.6151
R2217 B.n266 B.n263 10.6151
R2218 B.n267 B.n266 10.6151
R2219 B.n270 B.n267 10.6151
R2220 B.n271 B.n270 10.6151
R2221 B.n274 B.n271 10.6151
R2222 B.n275 B.n274 10.6151
R2223 B.n278 B.n275 10.6151
R2224 B.n279 B.n278 10.6151
R2225 B.n282 B.n279 10.6151
R2226 B.n283 B.n282 10.6151
R2227 B.n286 B.n283 10.6151
R2228 B.n287 B.n286 10.6151
R2229 B.n290 B.n287 10.6151
R2230 B.n291 B.n290 10.6151
R2231 B.n294 B.n291 10.6151
R2232 B.n295 B.n294 10.6151
R2233 B.n298 B.n295 10.6151
R2234 B.n299 B.n298 10.6151
R2235 B.n302 B.n299 10.6151
R2236 B.n303 B.n302 10.6151
R2237 B.n306 B.n303 10.6151
R2238 B.n307 B.n306 10.6151
R2239 B.n310 B.n307 10.6151
R2240 B.n311 B.n310 10.6151
R2241 B.n314 B.n311 10.6151
R2242 B.n315 B.n314 10.6151
R2243 B.n318 B.n315 10.6151
R2244 B.n319 B.n318 10.6151
R2245 B.n322 B.n319 10.6151
R2246 B.n324 B.n322 10.6151
R2247 B.n325 B.n324 10.6151
R2248 B.n976 B.n325 10.6151
R2249 B.n666 B.n665 10.6151
R2250 B.n666 B.n461 10.6151
R2251 B.n676 B.n461 10.6151
R2252 B.n677 B.n676 10.6151
R2253 B.n678 B.n677 10.6151
R2254 B.n678 B.n452 10.6151
R2255 B.n688 B.n452 10.6151
R2256 B.n689 B.n688 10.6151
R2257 B.n690 B.n689 10.6151
R2258 B.n690 B.n445 10.6151
R2259 B.n700 B.n445 10.6151
R2260 B.n701 B.n700 10.6151
R2261 B.n702 B.n701 10.6151
R2262 B.n702 B.n437 10.6151
R2263 B.n712 B.n437 10.6151
R2264 B.n713 B.n712 10.6151
R2265 B.n714 B.n713 10.6151
R2266 B.n714 B.n429 10.6151
R2267 B.n724 B.n429 10.6151
R2268 B.n725 B.n724 10.6151
R2269 B.n726 B.n725 10.6151
R2270 B.n726 B.n422 10.6151
R2271 B.n737 B.n422 10.6151
R2272 B.n738 B.n737 10.6151
R2273 B.n739 B.n738 10.6151
R2274 B.n739 B.n414 10.6151
R2275 B.n749 B.n414 10.6151
R2276 B.n750 B.n749 10.6151
R2277 B.n751 B.n750 10.6151
R2278 B.n751 B.n406 10.6151
R2279 B.n761 B.n406 10.6151
R2280 B.n762 B.n761 10.6151
R2281 B.n763 B.n762 10.6151
R2282 B.n763 B.n398 10.6151
R2283 B.n773 B.n398 10.6151
R2284 B.n774 B.n773 10.6151
R2285 B.n775 B.n774 10.6151
R2286 B.n775 B.n390 10.6151
R2287 B.n785 B.n390 10.6151
R2288 B.n786 B.n785 10.6151
R2289 B.n787 B.n786 10.6151
R2290 B.n787 B.n381 10.6151
R2291 B.n797 B.n381 10.6151
R2292 B.n798 B.n797 10.6151
R2293 B.n799 B.n798 10.6151
R2294 B.n799 B.n374 10.6151
R2295 B.n809 B.n374 10.6151
R2296 B.n810 B.n809 10.6151
R2297 B.n811 B.n810 10.6151
R2298 B.n811 B.n366 10.6151
R2299 B.n821 B.n366 10.6151
R2300 B.n822 B.n821 10.6151
R2301 B.n823 B.n822 10.6151
R2302 B.n823 B.n358 10.6151
R2303 B.n833 B.n358 10.6151
R2304 B.n834 B.n833 10.6151
R2305 B.n835 B.n834 10.6151
R2306 B.n835 B.n350 10.6151
R2307 B.n845 B.n350 10.6151
R2308 B.n846 B.n845 10.6151
R2309 B.n847 B.n846 10.6151
R2310 B.n847 B.n342 10.6151
R2311 B.n857 B.n342 10.6151
R2312 B.n858 B.n857 10.6151
R2313 B.n859 B.n858 10.6151
R2314 B.n859 B.n334 10.6151
R2315 B.n869 B.n334 10.6151
R2316 B.n870 B.n869 10.6151
R2317 B.n872 B.n870 10.6151
R2318 B.n872 B.n871 10.6151
R2319 B.n871 B.n326 10.6151
R2320 B.n883 B.n326 10.6151
R2321 B.n884 B.n883 10.6151
R2322 B.n885 B.n884 10.6151
R2323 B.n886 B.n885 10.6151
R2324 B.n888 B.n886 10.6151
R2325 B.n889 B.n888 10.6151
R2326 B.n890 B.n889 10.6151
R2327 B.n891 B.n890 10.6151
R2328 B.n893 B.n891 10.6151
R2329 B.n894 B.n893 10.6151
R2330 B.n895 B.n894 10.6151
R2331 B.n896 B.n895 10.6151
R2332 B.n898 B.n896 10.6151
R2333 B.n899 B.n898 10.6151
R2334 B.n900 B.n899 10.6151
R2335 B.n901 B.n900 10.6151
R2336 B.n903 B.n901 10.6151
R2337 B.n904 B.n903 10.6151
R2338 B.n905 B.n904 10.6151
R2339 B.n906 B.n905 10.6151
R2340 B.n908 B.n906 10.6151
R2341 B.n909 B.n908 10.6151
R2342 B.n910 B.n909 10.6151
R2343 B.n911 B.n910 10.6151
R2344 B.n913 B.n911 10.6151
R2345 B.n914 B.n913 10.6151
R2346 B.n915 B.n914 10.6151
R2347 B.n916 B.n915 10.6151
R2348 B.n918 B.n916 10.6151
R2349 B.n919 B.n918 10.6151
R2350 B.n920 B.n919 10.6151
R2351 B.n921 B.n920 10.6151
R2352 B.n923 B.n921 10.6151
R2353 B.n924 B.n923 10.6151
R2354 B.n925 B.n924 10.6151
R2355 B.n926 B.n925 10.6151
R2356 B.n928 B.n926 10.6151
R2357 B.n929 B.n928 10.6151
R2358 B.n930 B.n929 10.6151
R2359 B.n931 B.n930 10.6151
R2360 B.n933 B.n931 10.6151
R2361 B.n934 B.n933 10.6151
R2362 B.n935 B.n934 10.6151
R2363 B.n936 B.n935 10.6151
R2364 B.n938 B.n936 10.6151
R2365 B.n939 B.n938 10.6151
R2366 B.n940 B.n939 10.6151
R2367 B.n941 B.n940 10.6151
R2368 B.n943 B.n941 10.6151
R2369 B.n944 B.n943 10.6151
R2370 B.n945 B.n944 10.6151
R2371 B.n946 B.n945 10.6151
R2372 B.n948 B.n946 10.6151
R2373 B.n949 B.n948 10.6151
R2374 B.n950 B.n949 10.6151
R2375 B.n951 B.n950 10.6151
R2376 B.n953 B.n951 10.6151
R2377 B.n954 B.n953 10.6151
R2378 B.n955 B.n954 10.6151
R2379 B.n956 B.n955 10.6151
R2380 B.n958 B.n956 10.6151
R2381 B.n959 B.n958 10.6151
R2382 B.n960 B.n959 10.6151
R2383 B.n961 B.n960 10.6151
R2384 B.n963 B.n961 10.6151
R2385 B.n964 B.n963 10.6151
R2386 B.n965 B.n964 10.6151
R2387 B.n966 B.n965 10.6151
R2388 B.n968 B.n966 10.6151
R2389 B.n969 B.n968 10.6151
R2390 B.n970 B.n969 10.6151
R2391 B.n971 B.n970 10.6151
R2392 B.n973 B.n971 10.6151
R2393 B.n974 B.n973 10.6151
R2394 B.n975 B.n974 10.6151
R2395 B.n659 B.n658 10.6151
R2396 B.n658 B.n657 10.6151
R2397 B.n657 B.n656 10.6151
R2398 B.n656 B.n654 10.6151
R2399 B.n654 B.n651 10.6151
R2400 B.n651 B.n650 10.6151
R2401 B.n650 B.n647 10.6151
R2402 B.n647 B.n646 10.6151
R2403 B.n646 B.n643 10.6151
R2404 B.n643 B.n642 10.6151
R2405 B.n642 B.n639 10.6151
R2406 B.n639 B.n638 10.6151
R2407 B.n638 B.n635 10.6151
R2408 B.n635 B.n634 10.6151
R2409 B.n634 B.n631 10.6151
R2410 B.n631 B.n630 10.6151
R2411 B.n630 B.n627 10.6151
R2412 B.n627 B.n626 10.6151
R2413 B.n626 B.n623 10.6151
R2414 B.n623 B.n622 10.6151
R2415 B.n622 B.n619 10.6151
R2416 B.n619 B.n618 10.6151
R2417 B.n618 B.n615 10.6151
R2418 B.n615 B.n614 10.6151
R2419 B.n614 B.n611 10.6151
R2420 B.n611 B.n610 10.6151
R2421 B.n610 B.n607 10.6151
R2422 B.n607 B.n606 10.6151
R2423 B.n606 B.n603 10.6151
R2424 B.n603 B.n602 10.6151
R2425 B.n602 B.n599 10.6151
R2426 B.n599 B.n598 10.6151
R2427 B.n595 B.n594 10.6151
R2428 B.n594 B.n591 10.6151
R2429 B.n591 B.n590 10.6151
R2430 B.n590 B.n587 10.6151
R2431 B.n587 B.n586 10.6151
R2432 B.n586 B.n583 10.6151
R2433 B.n583 B.n582 10.6151
R2434 B.n582 B.n579 10.6151
R2435 B.n579 B.n578 10.6151
R2436 B.n575 B.n574 10.6151
R2437 B.n574 B.n571 10.6151
R2438 B.n571 B.n570 10.6151
R2439 B.n570 B.n567 10.6151
R2440 B.n567 B.n566 10.6151
R2441 B.n566 B.n563 10.6151
R2442 B.n563 B.n562 10.6151
R2443 B.n562 B.n559 10.6151
R2444 B.n559 B.n558 10.6151
R2445 B.n558 B.n555 10.6151
R2446 B.n555 B.n554 10.6151
R2447 B.n554 B.n551 10.6151
R2448 B.n551 B.n550 10.6151
R2449 B.n550 B.n547 10.6151
R2450 B.n547 B.n546 10.6151
R2451 B.n546 B.n543 10.6151
R2452 B.n543 B.n542 10.6151
R2453 B.n542 B.n539 10.6151
R2454 B.n539 B.n538 10.6151
R2455 B.n538 B.n535 10.6151
R2456 B.n535 B.n534 10.6151
R2457 B.n534 B.n531 10.6151
R2458 B.n531 B.n530 10.6151
R2459 B.n530 B.n527 10.6151
R2460 B.n527 B.n526 10.6151
R2461 B.n526 B.n523 10.6151
R2462 B.n523 B.n522 10.6151
R2463 B.n522 B.n519 10.6151
R2464 B.n519 B.n518 10.6151
R2465 B.n518 B.n515 10.6151
R2466 B.n515 B.n469 10.6151
R2467 B.n664 B.n469 10.6151
R2468 B.n670 B.n465 10.6151
R2469 B.n671 B.n670 10.6151
R2470 B.n672 B.n671 10.6151
R2471 B.n672 B.n457 10.6151
R2472 B.n682 B.n457 10.6151
R2473 B.n683 B.n682 10.6151
R2474 B.n684 B.n683 10.6151
R2475 B.n684 B.n449 10.6151
R2476 B.n694 B.n449 10.6151
R2477 B.n695 B.n694 10.6151
R2478 B.n696 B.n695 10.6151
R2479 B.n696 B.n441 10.6151
R2480 B.n706 B.n441 10.6151
R2481 B.n707 B.n706 10.6151
R2482 B.n708 B.n707 10.6151
R2483 B.n708 B.n433 10.6151
R2484 B.n718 B.n433 10.6151
R2485 B.n719 B.n718 10.6151
R2486 B.n720 B.n719 10.6151
R2487 B.n720 B.n425 10.6151
R2488 B.n731 B.n425 10.6151
R2489 B.n732 B.n731 10.6151
R2490 B.n733 B.n732 10.6151
R2491 B.n733 B.n418 10.6151
R2492 B.n743 B.n418 10.6151
R2493 B.n744 B.n743 10.6151
R2494 B.n745 B.n744 10.6151
R2495 B.n745 B.n410 10.6151
R2496 B.n755 B.n410 10.6151
R2497 B.n756 B.n755 10.6151
R2498 B.n757 B.n756 10.6151
R2499 B.n757 B.n402 10.6151
R2500 B.n767 B.n402 10.6151
R2501 B.n768 B.n767 10.6151
R2502 B.n769 B.n768 10.6151
R2503 B.n769 B.n394 10.6151
R2504 B.n779 B.n394 10.6151
R2505 B.n780 B.n779 10.6151
R2506 B.n781 B.n780 10.6151
R2507 B.n781 B.n386 10.6151
R2508 B.n791 B.n386 10.6151
R2509 B.n792 B.n791 10.6151
R2510 B.n793 B.n792 10.6151
R2511 B.n793 B.n378 10.6151
R2512 B.n803 B.n378 10.6151
R2513 B.n804 B.n803 10.6151
R2514 B.n805 B.n804 10.6151
R2515 B.n805 B.n370 10.6151
R2516 B.n815 B.n370 10.6151
R2517 B.n816 B.n815 10.6151
R2518 B.n817 B.n816 10.6151
R2519 B.n817 B.n362 10.6151
R2520 B.n827 B.n362 10.6151
R2521 B.n828 B.n827 10.6151
R2522 B.n829 B.n828 10.6151
R2523 B.n829 B.n354 10.6151
R2524 B.n839 B.n354 10.6151
R2525 B.n840 B.n839 10.6151
R2526 B.n841 B.n840 10.6151
R2527 B.n841 B.n346 10.6151
R2528 B.n851 B.n346 10.6151
R2529 B.n852 B.n851 10.6151
R2530 B.n853 B.n852 10.6151
R2531 B.n853 B.n338 10.6151
R2532 B.n863 B.n338 10.6151
R2533 B.n864 B.n863 10.6151
R2534 B.n865 B.n864 10.6151
R2535 B.n865 B.n330 10.6151
R2536 B.n876 B.n330 10.6151
R2537 B.n877 B.n876 10.6151
R2538 B.n878 B.n877 10.6151
R2539 B.n878 B.n0 10.6151
R2540 B.n1121 B.n1 10.6151
R2541 B.n1121 B.n1120 10.6151
R2542 B.n1120 B.n1119 10.6151
R2543 B.n1119 B.n10 10.6151
R2544 B.n1113 B.n10 10.6151
R2545 B.n1113 B.n1112 10.6151
R2546 B.n1112 B.n1111 10.6151
R2547 B.n1111 B.n17 10.6151
R2548 B.n1105 B.n17 10.6151
R2549 B.n1105 B.n1104 10.6151
R2550 B.n1104 B.n1103 10.6151
R2551 B.n1103 B.n24 10.6151
R2552 B.n1097 B.n24 10.6151
R2553 B.n1097 B.n1096 10.6151
R2554 B.n1096 B.n1095 10.6151
R2555 B.n1095 B.n31 10.6151
R2556 B.n1089 B.n31 10.6151
R2557 B.n1089 B.n1088 10.6151
R2558 B.n1088 B.n1087 10.6151
R2559 B.n1087 B.n38 10.6151
R2560 B.n1081 B.n38 10.6151
R2561 B.n1081 B.n1080 10.6151
R2562 B.n1080 B.n1079 10.6151
R2563 B.n1079 B.n45 10.6151
R2564 B.n1073 B.n45 10.6151
R2565 B.n1073 B.n1072 10.6151
R2566 B.n1072 B.n1071 10.6151
R2567 B.n1071 B.n52 10.6151
R2568 B.n1065 B.n52 10.6151
R2569 B.n1065 B.n1064 10.6151
R2570 B.n1064 B.n1063 10.6151
R2571 B.n1063 B.n59 10.6151
R2572 B.n1057 B.n59 10.6151
R2573 B.n1057 B.n1056 10.6151
R2574 B.n1056 B.n1055 10.6151
R2575 B.n1055 B.n66 10.6151
R2576 B.n1049 B.n66 10.6151
R2577 B.n1049 B.n1048 10.6151
R2578 B.n1048 B.n1047 10.6151
R2579 B.n1047 B.n73 10.6151
R2580 B.n1041 B.n73 10.6151
R2581 B.n1041 B.n1040 10.6151
R2582 B.n1040 B.n1039 10.6151
R2583 B.n1039 B.n80 10.6151
R2584 B.n1033 B.n80 10.6151
R2585 B.n1033 B.n1032 10.6151
R2586 B.n1032 B.n1031 10.6151
R2587 B.n1031 B.n87 10.6151
R2588 B.n1025 B.n87 10.6151
R2589 B.n1025 B.n1024 10.6151
R2590 B.n1024 B.n1023 10.6151
R2591 B.n1023 B.n93 10.6151
R2592 B.n1017 B.n93 10.6151
R2593 B.n1017 B.n1016 10.6151
R2594 B.n1016 B.n1015 10.6151
R2595 B.n1015 B.n101 10.6151
R2596 B.n1009 B.n101 10.6151
R2597 B.n1009 B.n1008 10.6151
R2598 B.n1008 B.n1007 10.6151
R2599 B.n1007 B.n108 10.6151
R2600 B.n1001 B.n108 10.6151
R2601 B.n1001 B.n1000 10.6151
R2602 B.n1000 B.n999 10.6151
R2603 B.n999 B.n115 10.6151
R2604 B.n993 B.n115 10.6151
R2605 B.n993 B.n992 10.6151
R2606 B.n992 B.n991 10.6151
R2607 B.n991 B.n122 10.6151
R2608 B.n985 B.n122 10.6151
R2609 B.n985 B.n984 10.6151
R2610 B.n984 B.n983 10.6151
R2611 B.n983 B.n129 10.6151
R2612 B.n241 B.n240 9.36635
R2613 B.n263 B.n262 9.36635
R2614 B.n598 B.n511 9.36635
R2615 B.n575 B.n514 9.36635
R2616 B.n831 B.t4 8.35397
R2617 B.t2 B.n1091 8.35397
R2618 B.n1127 B.n0 2.81026
R2619 B.n1127 B.n1 2.81026
R2620 B.n242 B.n241 1.24928
R2621 B.n262 B.n261 1.24928
R2622 B.n595 B.n511 1.24928
R2623 B.n578 B.n514 1.24928
R2624 B.t3 B.n336 0.759906
R2625 B.t7 B.n15 0.759906
R2626 VP.n32 VP.n31 161.3
R2627 VP.n33 VP.n28 161.3
R2628 VP.n35 VP.n34 161.3
R2629 VP.n36 VP.n27 161.3
R2630 VP.n38 VP.n37 161.3
R2631 VP.n39 VP.n26 161.3
R2632 VP.n41 VP.n40 161.3
R2633 VP.n42 VP.n25 161.3
R2634 VP.n44 VP.n43 161.3
R2635 VP.n45 VP.n24 161.3
R2636 VP.n47 VP.n46 161.3
R2637 VP.n48 VP.n23 161.3
R2638 VP.n50 VP.n49 161.3
R2639 VP.n51 VP.n22 161.3
R2640 VP.n53 VP.n52 161.3
R2641 VP.n55 VP.n54 161.3
R2642 VP.n56 VP.n20 161.3
R2643 VP.n58 VP.n57 161.3
R2644 VP.n59 VP.n19 161.3
R2645 VP.n61 VP.n60 161.3
R2646 VP.n62 VP.n18 161.3
R2647 VP.n64 VP.n63 161.3
R2648 VP.n111 VP.n110 161.3
R2649 VP.n109 VP.n1 161.3
R2650 VP.n108 VP.n107 161.3
R2651 VP.n106 VP.n2 161.3
R2652 VP.n105 VP.n104 161.3
R2653 VP.n103 VP.n3 161.3
R2654 VP.n102 VP.n101 161.3
R2655 VP.n100 VP.n99 161.3
R2656 VP.n98 VP.n5 161.3
R2657 VP.n97 VP.n96 161.3
R2658 VP.n95 VP.n6 161.3
R2659 VP.n94 VP.n93 161.3
R2660 VP.n92 VP.n7 161.3
R2661 VP.n91 VP.n90 161.3
R2662 VP.n89 VP.n8 161.3
R2663 VP.n88 VP.n87 161.3
R2664 VP.n86 VP.n9 161.3
R2665 VP.n85 VP.n84 161.3
R2666 VP.n83 VP.n10 161.3
R2667 VP.n82 VP.n81 161.3
R2668 VP.n80 VP.n11 161.3
R2669 VP.n79 VP.n78 161.3
R2670 VP.n77 VP.n76 161.3
R2671 VP.n75 VP.n13 161.3
R2672 VP.n74 VP.n73 161.3
R2673 VP.n72 VP.n14 161.3
R2674 VP.n71 VP.n70 161.3
R2675 VP.n69 VP.n15 161.3
R2676 VP.n68 VP.n67 161.3
R2677 VP.n30 VP.t0 99.4348
R2678 VP.n66 VP.n16 72.4512
R2679 VP.n112 VP.n0 72.4512
R2680 VP.n65 VP.n17 72.4512
R2681 VP.n8 VP.t4 66.2575
R2682 VP.n16 VP.t6 66.2575
R2683 VP.n12 VP.t9 66.2575
R2684 VP.n4 VP.t7 66.2575
R2685 VP.n0 VP.t8 66.2575
R2686 VP.n25 VP.t1 66.2575
R2687 VP.n17 VP.t5 66.2575
R2688 VP.n21 VP.t3 66.2575
R2689 VP.n29 VP.t2 66.2575
R2690 VP.n30 VP.n29 65.6329
R2691 VP.n85 VP.n10 56.0336
R2692 VP.n93 VP.n6 56.0336
R2693 VP.n46 VP.n23 56.0336
R2694 VP.n38 VP.n27 56.0336
R2695 VP.n66 VP.n65 55.2493
R2696 VP.n70 VP.n14 42.4359
R2697 VP.n108 VP.n2 42.4359
R2698 VP.n61 VP.n19 42.4359
R2699 VP.n74 VP.n14 38.5509
R2700 VP.n104 VP.n2 38.5509
R2701 VP.n57 VP.n19 38.5509
R2702 VP.n81 VP.n10 24.9531
R2703 VP.n97 VP.n6 24.9531
R2704 VP.n50 VP.n23 24.9531
R2705 VP.n34 VP.n27 24.9531
R2706 VP.n69 VP.n68 24.4675
R2707 VP.n70 VP.n69 24.4675
R2708 VP.n75 VP.n74 24.4675
R2709 VP.n76 VP.n75 24.4675
R2710 VP.n80 VP.n79 24.4675
R2711 VP.n81 VP.n80 24.4675
R2712 VP.n86 VP.n85 24.4675
R2713 VP.n87 VP.n86 24.4675
R2714 VP.n87 VP.n8 24.4675
R2715 VP.n91 VP.n8 24.4675
R2716 VP.n92 VP.n91 24.4675
R2717 VP.n93 VP.n92 24.4675
R2718 VP.n98 VP.n97 24.4675
R2719 VP.n99 VP.n98 24.4675
R2720 VP.n103 VP.n102 24.4675
R2721 VP.n104 VP.n103 24.4675
R2722 VP.n109 VP.n108 24.4675
R2723 VP.n110 VP.n109 24.4675
R2724 VP.n62 VP.n61 24.4675
R2725 VP.n63 VP.n62 24.4675
R2726 VP.n51 VP.n50 24.4675
R2727 VP.n52 VP.n51 24.4675
R2728 VP.n56 VP.n55 24.4675
R2729 VP.n57 VP.n56 24.4675
R2730 VP.n39 VP.n38 24.4675
R2731 VP.n40 VP.n39 24.4675
R2732 VP.n40 VP.n25 24.4675
R2733 VP.n44 VP.n25 24.4675
R2734 VP.n45 VP.n44 24.4675
R2735 VP.n46 VP.n45 24.4675
R2736 VP.n33 VP.n32 24.4675
R2737 VP.n34 VP.n33 24.4675
R2738 VP.n68 VP.n16 17.6167
R2739 VP.n110 VP.n0 17.6167
R2740 VP.n63 VP.n17 17.6167
R2741 VP.n76 VP.n12 15.6594
R2742 VP.n102 VP.n4 15.6594
R2743 VP.n55 VP.n21 15.6594
R2744 VP.n79 VP.n12 8.80862
R2745 VP.n99 VP.n4 8.80862
R2746 VP.n52 VP.n21 8.80862
R2747 VP.n32 VP.n29 8.80862
R2748 VP.n31 VP.n30 4.01766
R2749 VP.n65 VP.n64 0.354971
R2750 VP.n67 VP.n66 0.354971
R2751 VP.n112 VP.n111 0.354971
R2752 VP VP.n112 0.26696
R2753 VP.n31 VP.n28 0.189894
R2754 VP.n35 VP.n28 0.189894
R2755 VP.n36 VP.n35 0.189894
R2756 VP.n37 VP.n36 0.189894
R2757 VP.n37 VP.n26 0.189894
R2758 VP.n41 VP.n26 0.189894
R2759 VP.n42 VP.n41 0.189894
R2760 VP.n43 VP.n42 0.189894
R2761 VP.n43 VP.n24 0.189894
R2762 VP.n47 VP.n24 0.189894
R2763 VP.n48 VP.n47 0.189894
R2764 VP.n49 VP.n48 0.189894
R2765 VP.n49 VP.n22 0.189894
R2766 VP.n53 VP.n22 0.189894
R2767 VP.n54 VP.n53 0.189894
R2768 VP.n54 VP.n20 0.189894
R2769 VP.n58 VP.n20 0.189894
R2770 VP.n59 VP.n58 0.189894
R2771 VP.n60 VP.n59 0.189894
R2772 VP.n60 VP.n18 0.189894
R2773 VP.n64 VP.n18 0.189894
R2774 VP.n67 VP.n15 0.189894
R2775 VP.n71 VP.n15 0.189894
R2776 VP.n72 VP.n71 0.189894
R2777 VP.n73 VP.n72 0.189894
R2778 VP.n73 VP.n13 0.189894
R2779 VP.n77 VP.n13 0.189894
R2780 VP.n78 VP.n77 0.189894
R2781 VP.n78 VP.n11 0.189894
R2782 VP.n82 VP.n11 0.189894
R2783 VP.n83 VP.n82 0.189894
R2784 VP.n84 VP.n83 0.189894
R2785 VP.n84 VP.n9 0.189894
R2786 VP.n88 VP.n9 0.189894
R2787 VP.n89 VP.n88 0.189894
R2788 VP.n90 VP.n89 0.189894
R2789 VP.n90 VP.n7 0.189894
R2790 VP.n94 VP.n7 0.189894
R2791 VP.n95 VP.n94 0.189894
R2792 VP.n96 VP.n95 0.189894
R2793 VP.n96 VP.n5 0.189894
R2794 VP.n100 VP.n5 0.189894
R2795 VP.n101 VP.n100 0.189894
R2796 VP.n101 VP.n3 0.189894
R2797 VP.n105 VP.n3 0.189894
R2798 VP.n106 VP.n105 0.189894
R2799 VP.n107 VP.n106 0.189894
R2800 VP.n107 VP.n1 0.189894
R2801 VP.n111 VP.n1 0.189894
R2802 VDD1.n44 VDD1.n0 289.615
R2803 VDD1.n95 VDD1.n51 289.615
R2804 VDD1.n45 VDD1.n44 185
R2805 VDD1.n43 VDD1.n42 185
R2806 VDD1.n4 VDD1.n3 185
R2807 VDD1.n8 VDD1.n6 185
R2808 VDD1.n37 VDD1.n36 185
R2809 VDD1.n35 VDD1.n34 185
R2810 VDD1.n10 VDD1.n9 185
R2811 VDD1.n29 VDD1.n28 185
R2812 VDD1.n27 VDD1.n26 185
R2813 VDD1.n14 VDD1.n13 185
R2814 VDD1.n21 VDD1.n20 185
R2815 VDD1.n19 VDD1.n18 185
R2816 VDD1.n68 VDD1.n67 185
R2817 VDD1.n70 VDD1.n69 185
R2818 VDD1.n63 VDD1.n62 185
R2819 VDD1.n76 VDD1.n75 185
R2820 VDD1.n78 VDD1.n77 185
R2821 VDD1.n59 VDD1.n58 185
R2822 VDD1.n85 VDD1.n84 185
R2823 VDD1.n86 VDD1.n57 185
R2824 VDD1.n88 VDD1.n87 185
R2825 VDD1.n55 VDD1.n54 185
R2826 VDD1.n94 VDD1.n93 185
R2827 VDD1.n96 VDD1.n95 185
R2828 VDD1.n17 VDD1.t9 149.524
R2829 VDD1.n66 VDD1.t3 149.524
R2830 VDD1.n44 VDD1.n43 104.615
R2831 VDD1.n43 VDD1.n3 104.615
R2832 VDD1.n8 VDD1.n3 104.615
R2833 VDD1.n36 VDD1.n8 104.615
R2834 VDD1.n36 VDD1.n35 104.615
R2835 VDD1.n35 VDD1.n9 104.615
R2836 VDD1.n28 VDD1.n9 104.615
R2837 VDD1.n28 VDD1.n27 104.615
R2838 VDD1.n27 VDD1.n13 104.615
R2839 VDD1.n20 VDD1.n13 104.615
R2840 VDD1.n20 VDD1.n19 104.615
R2841 VDD1.n69 VDD1.n68 104.615
R2842 VDD1.n69 VDD1.n62 104.615
R2843 VDD1.n76 VDD1.n62 104.615
R2844 VDD1.n77 VDD1.n76 104.615
R2845 VDD1.n77 VDD1.n58 104.615
R2846 VDD1.n85 VDD1.n58 104.615
R2847 VDD1.n86 VDD1.n85 104.615
R2848 VDD1.n87 VDD1.n86 104.615
R2849 VDD1.n87 VDD1.n54 104.615
R2850 VDD1.n94 VDD1.n54 104.615
R2851 VDD1.n95 VDD1.n94 104.615
R2852 VDD1.n103 VDD1.n102 64.744
R2853 VDD1.n50 VDD1.n49 62.4202
R2854 VDD1.n105 VDD1.n104 62.4201
R2855 VDD1.n101 VDD1.n100 62.4201
R2856 VDD1.n19 VDD1.t9 52.3082
R2857 VDD1.n68 VDD1.t3 52.3082
R2858 VDD1.n50 VDD1.n48 51.4547
R2859 VDD1.n101 VDD1.n99 51.4547
R2860 VDD1.n105 VDD1.n103 48.8931
R2861 VDD1.n6 VDD1.n4 13.1884
R2862 VDD1.n88 VDD1.n55 13.1884
R2863 VDD1.n42 VDD1.n41 12.8005
R2864 VDD1.n38 VDD1.n37 12.8005
R2865 VDD1.n89 VDD1.n57 12.8005
R2866 VDD1.n93 VDD1.n92 12.8005
R2867 VDD1.n45 VDD1.n2 12.0247
R2868 VDD1.n34 VDD1.n7 12.0247
R2869 VDD1.n84 VDD1.n83 12.0247
R2870 VDD1.n96 VDD1.n53 12.0247
R2871 VDD1.n46 VDD1.n0 11.249
R2872 VDD1.n33 VDD1.n10 11.249
R2873 VDD1.n82 VDD1.n59 11.249
R2874 VDD1.n97 VDD1.n51 11.249
R2875 VDD1.n30 VDD1.n29 10.4732
R2876 VDD1.n79 VDD1.n78 10.4732
R2877 VDD1.n18 VDD1.n17 10.2747
R2878 VDD1.n67 VDD1.n66 10.2747
R2879 VDD1.n26 VDD1.n12 9.69747
R2880 VDD1.n75 VDD1.n61 9.69747
R2881 VDD1.n48 VDD1.n47 9.45567
R2882 VDD1.n99 VDD1.n98 9.45567
R2883 VDD1.n16 VDD1.n15 9.3005
R2884 VDD1.n23 VDD1.n22 9.3005
R2885 VDD1.n25 VDD1.n24 9.3005
R2886 VDD1.n12 VDD1.n11 9.3005
R2887 VDD1.n31 VDD1.n30 9.3005
R2888 VDD1.n33 VDD1.n32 9.3005
R2889 VDD1.n7 VDD1.n5 9.3005
R2890 VDD1.n39 VDD1.n38 9.3005
R2891 VDD1.n47 VDD1.n46 9.3005
R2892 VDD1.n2 VDD1.n1 9.3005
R2893 VDD1.n41 VDD1.n40 9.3005
R2894 VDD1.n98 VDD1.n97 9.3005
R2895 VDD1.n53 VDD1.n52 9.3005
R2896 VDD1.n92 VDD1.n91 9.3005
R2897 VDD1.n65 VDD1.n64 9.3005
R2898 VDD1.n72 VDD1.n71 9.3005
R2899 VDD1.n74 VDD1.n73 9.3005
R2900 VDD1.n61 VDD1.n60 9.3005
R2901 VDD1.n80 VDD1.n79 9.3005
R2902 VDD1.n82 VDD1.n81 9.3005
R2903 VDD1.n83 VDD1.n56 9.3005
R2904 VDD1.n90 VDD1.n89 9.3005
R2905 VDD1.n25 VDD1.n14 8.92171
R2906 VDD1.n74 VDD1.n63 8.92171
R2907 VDD1.n22 VDD1.n21 8.14595
R2908 VDD1.n71 VDD1.n70 8.14595
R2909 VDD1.n18 VDD1.n16 7.3702
R2910 VDD1.n67 VDD1.n65 7.3702
R2911 VDD1.n21 VDD1.n16 5.81868
R2912 VDD1.n70 VDD1.n65 5.81868
R2913 VDD1.n22 VDD1.n14 5.04292
R2914 VDD1.n71 VDD1.n63 5.04292
R2915 VDD1.n26 VDD1.n25 4.26717
R2916 VDD1.n75 VDD1.n74 4.26717
R2917 VDD1.n29 VDD1.n12 3.49141
R2918 VDD1.n78 VDD1.n61 3.49141
R2919 VDD1.n17 VDD1.n15 2.84303
R2920 VDD1.n66 VDD1.n64 2.84303
R2921 VDD1.n48 VDD1.n0 2.71565
R2922 VDD1.n30 VDD1.n10 2.71565
R2923 VDD1.n79 VDD1.n59 2.71565
R2924 VDD1.n99 VDD1.n51 2.71565
R2925 VDD1 VDD1.n105 2.32162
R2926 VDD1.n104 VDD1.t6 2.15034
R2927 VDD1.n104 VDD1.t4 2.15034
R2928 VDD1.n49 VDD1.t7 2.15034
R2929 VDD1.n49 VDD1.t8 2.15034
R2930 VDD1.n102 VDD1.t2 2.15034
R2931 VDD1.n102 VDD1.t1 2.15034
R2932 VDD1.n100 VDD1.t0 2.15034
R2933 VDD1.n100 VDD1.t5 2.15034
R2934 VDD1.n46 VDD1.n45 1.93989
R2935 VDD1.n34 VDD1.n33 1.93989
R2936 VDD1.n84 VDD1.n82 1.93989
R2937 VDD1.n97 VDD1.n96 1.93989
R2938 VDD1.n42 VDD1.n2 1.16414
R2939 VDD1.n37 VDD1.n7 1.16414
R2940 VDD1.n83 VDD1.n57 1.16414
R2941 VDD1.n93 VDD1.n53 1.16414
R2942 VDD1 VDD1.n50 0.851793
R2943 VDD1.n103 VDD1.n101 0.738257
R2944 VDD1.n41 VDD1.n4 0.388379
R2945 VDD1.n38 VDD1.n6 0.388379
R2946 VDD1.n89 VDD1.n88 0.388379
R2947 VDD1.n92 VDD1.n55 0.388379
R2948 VDD1.n47 VDD1.n1 0.155672
R2949 VDD1.n40 VDD1.n1 0.155672
R2950 VDD1.n40 VDD1.n39 0.155672
R2951 VDD1.n39 VDD1.n5 0.155672
R2952 VDD1.n32 VDD1.n5 0.155672
R2953 VDD1.n32 VDD1.n31 0.155672
R2954 VDD1.n31 VDD1.n11 0.155672
R2955 VDD1.n24 VDD1.n11 0.155672
R2956 VDD1.n24 VDD1.n23 0.155672
R2957 VDD1.n23 VDD1.n15 0.155672
R2958 VDD1.n72 VDD1.n64 0.155672
R2959 VDD1.n73 VDD1.n72 0.155672
R2960 VDD1.n73 VDD1.n60 0.155672
R2961 VDD1.n80 VDD1.n60 0.155672
R2962 VDD1.n81 VDD1.n80 0.155672
R2963 VDD1.n81 VDD1.n56 0.155672
R2964 VDD1.n90 VDD1.n56 0.155672
R2965 VDD1.n91 VDD1.n90 0.155672
R2966 VDD1.n91 VDD1.n52 0.155672
R2967 VDD1.n98 VDD1.n52 0.155672
C0 VP VN 8.985769f
C1 VDD1 VDD2 2.66191f
C2 VP VTAIL 9.800691f
C3 VDD2 VP 0.678979f
C4 VDD1 VP 9.212951f
C5 VN VTAIL 9.786481f
C6 VDD2 VN 8.69246f
C7 VDD2 VTAIL 9.62444f
C8 VDD1 VN 0.154964f
C9 VDD1 VTAIL 9.5673f
C10 VDD2 B 7.615208f
C11 VDD1 B 7.568449f
C12 VTAIL B 7.654774f
C13 VN B 21.51902f
C14 VP B 20.104988f
C15 VDD1.n0 B 0.033019f
C16 VDD1.n1 B 0.025848f
C17 VDD1.n2 B 0.01389f
C18 VDD1.n3 B 0.03283f
C19 VDD1.n4 B 0.014298f
C20 VDD1.n5 B 0.025848f
C21 VDD1.n6 B 0.014298f
C22 VDD1.n7 B 0.01389f
C23 VDD1.n8 B 0.03283f
C24 VDD1.n9 B 0.03283f
C25 VDD1.n10 B 0.014707f
C26 VDD1.n11 B 0.025848f
C27 VDD1.n12 B 0.01389f
C28 VDD1.n13 B 0.03283f
C29 VDD1.n14 B 0.014707f
C30 VDD1.n15 B 0.983234f
C31 VDD1.n16 B 0.01389f
C32 VDD1.t9 B 0.055063f
C33 VDD1.n17 B 0.158683f
C34 VDD1.n18 B 0.023209f
C35 VDD1.n19 B 0.024623f
C36 VDD1.n20 B 0.03283f
C37 VDD1.n21 B 0.014707f
C38 VDD1.n22 B 0.01389f
C39 VDD1.n23 B 0.025848f
C40 VDD1.n24 B 0.025848f
C41 VDD1.n25 B 0.01389f
C42 VDD1.n26 B 0.014707f
C43 VDD1.n27 B 0.03283f
C44 VDD1.n28 B 0.03283f
C45 VDD1.n29 B 0.014707f
C46 VDD1.n30 B 0.01389f
C47 VDD1.n31 B 0.025848f
C48 VDD1.n32 B 0.025848f
C49 VDD1.n33 B 0.01389f
C50 VDD1.n34 B 0.014707f
C51 VDD1.n35 B 0.03283f
C52 VDD1.n36 B 0.03283f
C53 VDD1.n37 B 0.014707f
C54 VDD1.n38 B 0.01389f
C55 VDD1.n39 B 0.025848f
C56 VDD1.n40 B 0.025848f
C57 VDD1.n41 B 0.01389f
C58 VDD1.n42 B 0.014707f
C59 VDD1.n43 B 0.03283f
C60 VDD1.n44 B 0.065213f
C61 VDD1.n45 B 0.014707f
C62 VDD1.n46 B 0.01389f
C63 VDD1.n47 B 0.058688f
C64 VDD1.n48 B 0.073033f
C65 VDD1.t7 B 0.188126f
C66 VDD1.t8 B 0.188126f
C67 VDD1.n49 B 1.64602f
C68 VDD1.n50 B 0.838997f
C69 VDD1.n51 B 0.033019f
C70 VDD1.n52 B 0.025848f
C71 VDD1.n53 B 0.01389f
C72 VDD1.n54 B 0.03283f
C73 VDD1.n55 B 0.014298f
C74 VDD1.n56 B 0.025848f
C75 VDD1.n57 B 0.014707f
C76 VDD1.n58 B 0.03283f
C77 VDD1.n59 B 0.014707f
C78 VDD1.n60 B 0.025848f
C79 VDD1.n61 B 0.01389f
C80 VDD1.n62 B 0.03283f
C81 VDD1.n63 B 0.014707f
C82 VDD1.n64 B 0.983234f
C83 VDD1.n65 B 0.01389f
C84 VDD1.t3 B 0.055063f
C85 VDD1.n66 B 0.158683f
C86 VDD1.n67 B 0.023209f
C87 VDD1.n68 B 0.024623f
C88 VDD1.n69 B 0.03283f
C89 VDD1.n70 B 0.014707f
C90 VDD1.n71 B 0.01389f
C91 VDD1.n72 B 0.025848f
C92 VDD1.n73 B 0.025848f
C93 VDD1.n74 B 0.01389f
C94 VDD1.n75 B 0.014707f
C95 VDD1.n76 B 0.03283f
C96 VDD1.n77 B 0.03283f
C97 VDD1.n78 B 0.014707f
C98 VDD1.n79 B 0.01389f
C99 VDD1.n80 B 0.025848f
C100 VDD1.n81 B 0.025848f
C101 VDD1.n82 B 0.01389f
C102 VDD1.n83 B 0.01389f
C103 VDD1.n84 B 0.014707f
C104 VDD1.n85 B 0.03283f
C105 VDD1.n86 B 0.03283f
C106 VDD1.n87 B 0.03283f
C107 VDD1.n88 B 0.014298f
C108 VDD1.n89 B 0.01389f
C109 VDD1.n90 B 0.025848f
C110 VDD1.n91 B 0.025848f
C111 VDD1.n92 B 0.01389f
C112 VDD1.n93 B 0.014707f
C113 VDD1.n94 B 0.03283f
C114 VDD1.n95 B 0.065213f
C115 VDD1.n96 B 0.014707f
C116 VDD1.n97 B 0.01389f
C117 VDD1.n98 B 0.058688f
C118 VDD1.n99 B 0.073033f
C119 VDD1.t0 B 0.188126f
C120 VDD1.t5 B 0.188126f
C121 VDD1.n100 B 1.64602f
C122 VDD1.n101 B 0.83036f
C123 VDD1.t2 B 0.188126f
C124 VDD1.t1 B 0.188126f
C125 VDD1.n102 B 1.67036f
C126 VDD1.n103 B 3.37463f
C127 VDD1.t6 B 0.188126f
C128 VDD1.t4 B 0.188126f
C129 VDD1.n104 B 1.64602f
C130 VDD1.n105 B 3.37946f
C131 VP.t8 B 1.61637f
C132 VP.n0 B 0.658067f
C133 VP.n1 B 0.019396f
C134 VP.n2 B 0.015779f
C135 VP.n3 B 0.019396f
C136 VP.t7 B 1.61637f
C137 VP.n4 B 0.576868f
C138 VP.n5 B 0.019396f
C139 VP.n6 B 0.023158f
C140 VP.n7 B 0.019396f
C141 VP.t4 B 1.61637f
C142 VP.n8 B 0.59517f
C143 VP.n9 B 0.019396f
C144 VP.n10 B 0.023158f
C145 VP.n11 B 0.019396f
C146 VP.t9 B 1.61637f
C147 VP.n12 B 0.576868f
C148 VP.n13 B 0.019396f
C149 VP.n14 B 0.015779f
C150 VP.n15 B 0.019396f
C151 VP.t6 B 1.61637f
C152 VP.n16 B 0.658067f
C153 VP.t5 B 1.61637f
C154 VP.n17 B 0.658067f
C155 VP.n18 B 0.019396f
C156 VP.n19 B 0.015779f
C157 VP.n20 B 0.019396f
C158 VP.t3 B 1.61637f
C159 VP.n21 B 0.576868f
C160 VP.n22 B 0.019396f
C161 VP.n23 B 0.023158f
C162 VP.n24 B 0.019396f
C163 VP.t1 B 1.61637f
C164 VP.n25 B 0.59517f
C165 VP.n26 B 0.019396f
C166 VP.n27 B 0.023158f
C167 VP.n28 B 0.019396f
C168 VP.t2 B 1.61637f
C169 VP.n29 B 0.639773f
C170 VP.t0 B 1.85636f
C171 VP.n30 B 0.608094f
C172 VP.n31 B 0.227933f
C173 VP.n32 B 0.024727f
C174 VP.n33 B 0.036149f
C175 VP.n34 B 0.036488f
C176 VP.n35 B 0.019396f
C177 VP.n36 B 0.019396f
C178 VP.n37 B 0.019396f
C179 VP.n38 B 0.033131f
C180 VP.n39 B 0.036149f
C181 VP.n40 B 0.036149f
C182 VP.n41 B 0.019396f
C183 VP.n42 B 0.019396f
C184 VP.n43 B 0.019396f
C185 VP.n44 B 0.036149f
C186 VP.n45 B 0.036149f
C187 VP.n46 B 0.033131f
C188 VP.n47 B 0.019396f
C189 VP.n48 B 0.019396f
C190 VP.n49 B 0.019396f
C191 VP.n50 B 0.036488f
C192 VP.n51 B 0.036149f
C193 VP.n52 B 0.024727f
C194 VP.n53 B 0.019396f
C195 VP.n54 B 0.019396f
C196 VP.n55 B 0.029724f
C197 VP.n56 B 0.036149f
C198 VP.n57 B 0.038886f
C199 VP.n58 B 0.019396f
C200 VP.n59 B 0.019396f
C201 VP.n60 B 0.019396f
C202 VP.n61 B 0.038112f
C203 VP.n62 B 0.036149f
C204 VP.n63 B 0.031151f
C205 VP.n64 B 0.031304f
C206 VP.n65 B 1.26889f
C207 VP.n66 B 1.28151f
C208 VP.n67 B 0.031304f
C209 VP.n68 B 0.031151f
C210 VP.n69 B 0.036149f
C211 VP.n70 B 0.038112f
C212 VP.n71 B 0.019396f
C213 VP.n72 B 0.019396f
C214 VP.n73 B 0.019396f
C215 VP.n74 B 0.038886f
C216 VP.n75 B 0.036149f
C217 VP.n76 B 0.029724f
C218 VP.n77 B 0.019396f
C219 VP.n78 B 0.019396f
C220 VP.n79 B 0.024727f
C221 VP.n80 B 0.036149f
C222 VP.n81 B 0.036488f
C223 VP.n82 B 0.019396f
C224 VP.n83 B 0.019396f
C225 VP.n84 B 0.019396f
C226 VP.n85 B 0.033131f
C227 VP.n86 B 0.036149f
C228 VP.n87 B 0.036149f
C229 VP.n88 B 0.019396f
C230 VP.n89 B 0.019396f
C231 VP.n90 B 0.019396f
C232 VP.n91 B 0.036149f
C233 VP.n92 B 0.036149f
C234 VP.n93 B 0.033131f
C235 VP.n94 B 0.019396f
C236 VP.n95 B 0.019396f
C237 VP.n96 B 0.019396f
C238 VP.n97 B 0.036488f
C239 VP.n98 B 0.036149f
C240 VP.n99 B 0.024727f
C241 VP.n100 B 0.019396f
C242 VP.n101 B 0.019396f
C243 VP.n102 B 0.029724f
C244 VP.n103 B 0.036149f
C245 VP.n104 B 0.038886f
C246 VP.n105 B 0.019396f
C247 VP.n106 B 0.019396f
C248 VP.n107 B 0.019396f
C249 VP.n108 B 0.038112f
C250 VP.n109 B 0.036149f
C251 VP.n110 B 0.031151f
C252 VP.n111 B 0.031304f
C253 VP.n112 B 0.044848f
C254 VTAIL.t14 B 0.194865f
C255 VTAIL.t18 B 0.194865f
C256 VTAIL.n0 B 1.6276f
C257 VTAIL.n1 B 0.645975f
C258 VTAIL.n2 B 0.034202f
C259 VTAIL.n3 B 0.026774f
C260 VTAIL.n4 B 0.014387f
C261 VTAIL.n5 B 0.034007f
C262 VTAIL.n6 B 0.014811f
C263 VTAIL.n7 B 0.026774f
C264 VTAIL.n8 B 0.015234f
C265 VTAIL.n9 B 0.034007f
C266 VTAIL.n10 B 0.015234f
C267 VTAIL.n11 B 0.026774f
C268 VTAIL.n12 B 0.014387f
C269 VTAIL.n13 B 0.034007f
C270 VTAIL.n14 B 0.015234f
C271 VTAIL.n15 B 1.01846f
C272 VTAIL.n16 B 0.014387f
C273 VTAIL.t3 B 0.057036f
C274 VTAIL.n17 B 0.164367f
C275 VTAIL.n18 B 0.02404f
C276 VTAIL.n19 B 0.025505f
C277 VTAIL.n20 B 0.034007f
C278 VTAIL.n21 B 0.015234f
C279 VTAIL.n22 B 0.014387f
C280 VTAIL.n23 B 0.026774f
C281 VTAIL.n24 B 0.026774f
C282 VTAIL.n25 B 0.014387f
C283 VTAIL.n26 B 0.015234f
C284 VTAIL.n27 B 0.034007f
C285 VTAIL.n28 B 0.034007f
C286 VTAIL.n29 B 0.015234f
C287 VTAIL.n30 B 0.014387f
C288 VTAIL.n31 B 0.026774f
C289 VTAIL.n32 B 0.026774f
C290 VTAIL.n33 B 0.014387f
C291 VTAIL.n34 B 0.014387f
C292 VTAIL.n35 B 0.015234f
C293 VTAIL.n36 B 0.034007f
C294 VTAIL.n37 B 0.034007f
C295 VTAIL.n38 B 0.034007f
C296 VTAIL.n39 B 0.014811f
C297 VTAIL.n40 B 0.014387f
C298 VTAIL.n41 B 0.026774f
C299 VTAIL.n42 B 0.026774f
C300 VTAIL.n43 B 0.014387f
C301 VTAIL.n44 B 0.015234f
C302 VTAIL.n45 B 0.034007f
C303 VTAIL.n46 B 0.067549f
C304 VTAIL.n47 B 0.015234f
C305 VTAIL.n48 B 0.014387f
C306 VTAIL.n49 B 0.060791f
C307 VTAIL.n50 B 0.037138f
C308 VTAIL.n51 B 0.473323f
C309 VTAIL.t5 B 0.194865f
C310 VTAIL.t4 B 0.194865f
C311 VTAIL.n52 B 1.6276f
C312 VTAIL.n53 B 0.805692f
C313 VTAIL.t6 B 0.194865f
C314 VTAIL.t19 B 0.194865f
C315 VTAIL.n54 B 1.6276f
C316 VTAIL.n55 B 2.12806f
C317 VTAIL.t17 B 0.194865f
C318 VTAIL.t16 B 0.194865f
C319 VTAIL.n56 B 1.62761f
C320 VTAIL.n57 B 2.12805f
C321 VTAIL.t13 B 0.194865f
C322 VTAIL.t9 B 0.194865f
C323 VTAIL.n58 B 1.62761f
C324 VTAIL.n59 B 0.805682f
C325 VTAIL.n60 B 0.034202f
C326 VTAIL.n61 B 0.026774f
C327 VTAIL.n62 B 0.014387f
C328 VTAIL.n63 B 0.034007f
C329 VTAIL.n64 B 0.014811f
C330 VTAIL.n65 B 0.026774f
C331 VTAIL.n66 B 0.014811f
C332 VTAIL.n67 B 0.014387f
C333 VTAIL.n68 B 0.034007f
C334 VTAIL.n69 B 0.034007f
C335 VTAIL.n70 B 0.015234f
C336 VTAIL.n71 B 0.026774f
C337 VTAIL.n72 B 0.014387f
C338 VTAIL.n73 B 0.034007f
C339 VTAIL.n74 B 0.015234f
C340 VTAIL.n75 B 1.01846f
C341 VTAIL.n76 B 0.014387f
C342 VTAIL.t11 B 0.057036f
C343 VTAIL.n77 B 0.164367f
C344 VTAIL.n78 B 0.02404f
C345 VTAIL.n79 B 0.025505f
C346 VTAIL.n80 B 0.034007f
C347 VTAIL.n81 B 0.015234f
C348 VTAIL.n82 B 0.014387f
C349 VTAIL.n83 B 0.026774f
C350 VTAIL.n84 B 0.026774f
C351 VTAIL.n85 B 0.014387f
C352 VTAIL.n86 B 0.015234f
C353 VTAIL.n87 B 0.034007f
C354 VTAIL.n88 B 0.034007f
C355 VTAIL.n89 B 0.015234f
C356 VTAIL.n90 B 0.014387f
C357 VTAIL.n91 B 0.026774f
C358 VTAIL.n92 B 0.026774f
C359 VTAIL.n93 B 0.014387f
C360 VTAIL.n94 B 0.015234f
C361 VTAIL.n95 B 0.034007f
C362 VTAIL.n96 B 0.034007f
C363 VTAIL.n97 B 0.015234f
C364 VTAIL.n98 B 0.014387f
C365 VTAIL.n99 B 0.026774f
C366 VTAIL.n100 B 0.026774f
C367 VTAIL.n101 B 0.014387f
C368 VTAIL.n102 B 0.015234f
C369 VTAIL.n103 B 0.034007f
C370 VTAIL.n104 B 0.067549f
C371 VTAIL.n105 B 0.015234f
C372 VTAIL.n106 B 0.014387f
C373 VTAIL.n107 B 0.060791f
C374 VTAIL.n108 B 0.037138f
C375 VTAIL.n109 B 0.473323f
C376 VTAIL.t7 B 0.194865f
C377 VTAIL.t2 B 0.194865f
C378 VTAIL.n110 B 1.62761f
C379 VTAIL.n111 B 0.709368f
C380 VTAIL.t8 B 0.194865f
C381 VTAIL.t1 B 0.194865f
C382 VTAIL.n112 B 1.62761f
C383 VTAIL.n113 B 0.805682f
C384 VTAIL.n114 B 0.034202f
C385 VTAIL.n115 B 0.026774f
C386 VTAIL.n116 B 0.014387f
C387 VTAIL.n117 B 0.034007f
C388 VTAIL.n118 B 0.014811f
C389 VTAIL.n119 B 0.026774f
C390 VTAIL.n120 B 0.014811f
C391 VTAIL.n121 B 0.014387f
C392 VTAIL.n122 B 0.034007f
C393 VTAIL.n123 B 0.034007f
C394 VTAIL.n124 B 0.015234f
C395 VTAIL.n125 B 0.026774f
C396 VTAIL.n126 B 0.014387f
C397 VTAIL.n127 B 0.034007f
C398 VTAIL.n128 B 0.015234f
C399 VTAIL.n129 B 1.01846f
C400 VTAIL.n130 B 0.014387f
C401 VTAIL.t0 B 0.057036f
C402 VTAIL.n131 B 0.164367f
C403 VTAIL.n132 B 0.02404f
C404 VTAIL.n133 B 0.025505f
C405 VTAIL.n134 B 0.034007f
C406 VTAIL.n135 B 0.015234f
C407 VTAIL.n136 B 0.014387f
C408 VTAIL.n137 B 0.026774f
C409 VTAIL.n138 B 0.026774f
C410 VTAIL.n139 B 0.014387f
C411 VTAIL.n140 B 0.015234f
C412 VTAIL.n141 B 0.034007f
C413 VTAIL.n142 B 0.034007f
C414 VTAIL.n143 B 0.015234f
C415 VTAIL.n144 B 0.014387f
C416 VTAIL.n145 B 0.026774f
C417 VTAIL.n146 B 0.026774f
C418 VTAIL.n147 B 0.014387f
C419 VTAIL.n148 B 0.015234f
C420 VTAIL.n149 B 0.034007f
C421 VTAIL.n150 B 0.034007f
C422 VTAIL.n151 B 0.015234f
C423 VTAIL.n152 B 0.014387f
C424 VTAIL.n153 B 0.026774f
C425 VTAIL.n154 B 0.026774f
C426 VTAIL.n155 B 0.014387f
C427 VTAIL.n156 B 0.015234f
C428 VTAIL.n157 B 0.034007f
C429 VTAIL.n158 B 0.067549f
C430 VTAIL.n159 B 0.015234f
C431 VTAIL.n160 B 0.014387f
C432 VTAIL.n161 B 0.060791f
C433 VTAIL.n162 B 0.037138f
C434 VTAIL.n163 B 1.61831f
C435 VTAIL.n164 B 0.034202f
C436 VTAIL.n165 B 0.026774f
C437 VTAIL.n166 B 0.014387f
C438 VTAIL.n167 B 0.034007f
C439 VTAIL.n168 B 0.014811f
C440 VTAIL.n169 B 0.026774f
C441 VTAIL.n170 B 0.015234f
C442 VTAIL.n171 B 0.034007f
C443 VTAIL.n172 B 0.015234f
C444 VTAIL.n173 B 0.026774f
C445 VTAIL.n174 B 0.014387f
C446 VTAIL.n175 B 0.034007f
C447 VTAIL.n176 B 0.015234f
C448 VTAIL.n177 B 1.01846f
C449 VTAIL.n178 B 0.014387f
C450 VTAIL.t15 B 0.057036f
C451 VTAIL.n179 B 0.164367f
C452 VTAIL.n180 B 0.02404f
C453 VTAIL.n181 B 0.025505f
C454 VTAIL.n182 B 0.034007f
C455 VTAIL.n183 B 0.015234f
C456 VTAIL.n184 B 0.014387f
C457 VTAIL.n185 B 0.026774f
C458 VTAIL.n186 B 0.026774f
C459 VTAIL.n187 B 0.014387f
C460 VTAIL.n188 B 0.015234f
C461 VTAIL.n189 B 0.034007f
C462 VTAIL.n190 B 0.034007f
C463 VTAIL.n191 B 0.015234f
C464 VTAIL.n192 B 0.014387f
C465 VTAIL.n193 B 0.026774f
C466 VTAIL.n194 B 0.026774f
C467 VTAIL.n195 B 0.014387f
C468 VTAIL.n196 B 0.014387f
C469 VTAIL.n197 B 0.015234f
C470 VTAIL.n198 B 0.034007f
C471 VTAIL.n199 B 0.034007f
C472 VTAIL.n200 B 0.034007f
C473 VTAIL.n201 B 0.014811f
C474 VTAIL.n202 B 0.014387f
C475 VTAIL.n203 B 0.026774f
C476 VTAIL.n204 B 0.026774f
C477 VTAIL.n205 B 0.014387f
C478 VTAIL.n206 B 0.015234f
C479 VTAIL.n207 B 0.034007f
C480 VTAIL.n208 B 0.067549f
C481 VTAIL.n209 B 0.015234f
C482 VTAIL.n210 B 0.014387f
C483 VTAIL.n211 B 0.060791f
C484 VTAIL.n212 B 0.037138f
C485 VTAIL.n213 B 1.61831f
C486 VTAIL.t12 B 0.194865f
C487 VTAIL.t10 B 0.194865f
C488 VTAIL.n214 B 1.6276f
C489 VTAIL.n215 B 0.595402f
C490 VDD2.n0 B 0.032395f
C491 VDD2.n1 B 0.02536f
C492 VDD2.n2 B 0.013627f
C493 VDD2.n3 B 0.03221f
C494 VDD2.n4 B 0.014028f
C495 VDD2.n5 B 0.02536f
C496 VDD2.n6 B 0.014429f
C497 VDD2.n7 B 0.03221f
C498 VDD2.n8 B 0.014429f
C499 VDD2.n9 B 0.02536f
C500 VDD2.n10 B 0.013627f
C501 VDD2.n11 B 0.03221f
C502 VDD2.n12 B 0.014429f
C503 VDD2.n13 B 0.964651f
C504 VDD2.n14 B 0.013627f
C505 VDD2.t2 B 0.054023f
C506 VDD2.n15 B 0.155684f
C507 VDD2.n16 B 0.02277f
C508 VDD2.n17 B 0.024157f
C509 VDD2.n18 B 0.03221f
C510 VDD2.n19 B 0.014429f
C511 VDD2.n20 B 0.013627f
C512 VDD2.n21 B 0.02536f
C513 VDD2.n22 B 0.02536f
C514 VDD2.n23 B 0.013627f
C515 VDD2.n24 B 0.014429f
C516 VDD2.n25 B 0.03221f
C517 VDD2.n26 B 0.03221f
C518 VDD2.n27 B 0.014429f
C519 VDD2.n28 B 0.013627f
C520 VDD2.n29 B 0.02536f
C521 VDD2.n30 B 0.02536f
C522 VDD2.n31 B 0.013627f
C523 VDD2.n32 B 0.013627f
C524 VDD2.n33 B 0.014429f
C525 VDD2.n34 B 0.03221f
C526 VDD2.n35 B 0.03221f
C527 VDD2.n36 B 0.03221f
C528 VDD2.n37 B 0.014028f
C529 VDD2.n38 B 0.013627f
C530 VDD2.n39 B 0.02536f
C531 VDD2.n40 B 0.02536f
C532 VDD2.n41 B 0.013627f
C533 VDD2.n42 B 0.014429f
C534 VDD2.n43 B 0.03221f
C535 VDD2.n44 B 0.06398f
C536 VDD2.n45 B 0.014429f
C537 VDD2.n46 B 0.013627f
C538 VDD2.n47 B 0.057579f
C539 VDD2.n48 B 0.071652f
C540 VDD2.t8 B 0.18457f
C541 VDD2.t6 B 0.18457f
C542 VDD2.n49 B 1.61491f
C543 VDD2.n50 B 0.814666f
C544 VDD2.t5 B 0.18457f
C545 VDD2.t0 B 0.18457f
C546 VDD2.n51 B 1.63879f
C547 VDD2.n52 B 3.1655f
C548 VDD2.n53 B 0.032395f
C549 VDD2.n54 B 0.02536f
C550 VDD2.n55 B 0.013627f
C551 VDD2.n56 B 0.03221f
C552 VDD2.n57 B 0.014028f
C553 VDD2.n58 B 0.02536f
C554 VDD2.n59 B 0.014028f
C555 VDD2.n60 B 0.013627f
C556 VDD2.n61 B 0.03221f
C557 VDD2.n62 B 0.03221f
C558 VDD2.n63 B 0.014429f
C559 VDD2.n64 B 0.02536f
C560 VDD2.n65 B 0.013627f
C561 VDD2.n66 B 0.03221f
C562 VDD2.n67 B 0.014429f
C563 VDD2.n68 B 0.964651f
C564 VDD2.n69 B 0.013627f
C565 VDD2.t3 B 0.054023f
C566 VDD2.n70 B 0.155684f
C567 VDD2.n71 B 0.02277f
C568 VDD2.n72 B 0.024157f
C569 VDD2.n73 B 0.03221f
C570 VDD2.n74 B 0.014429f
C571 VDD2.n75 B 0.013627f
C572 VDD2.n76 B 0.02536f
C573 VDD2.n77 B 0.02536f
C574 VDD2.n78 B 0.013627f
C575 VDD2.n79 B 0.014429f
C576 VDD2.n80 B 0.03221f
C577 VDD2.n81 B 0.03221f
C578 VDD2.n82 B 0.014429f
C579 VDD2.n83 B 0.013627f
C580 VDD2.n84 B 0.02536f
C581 VDD2.n85 B 0.02536f
C582 VDD2.n86 B 0.013627f
C583 VDD2.n87 B 0.014429f
C584 VDD2.n88 B 0.03221f
C585 VDD2.n89 B 0.03221f
C586 VDD2.n90 B 0.014429f
C587 VDD2.n91 B 0.013627f
C588 VDD2.n92 B 0.02536f
C589 VDD2.n93 B 0.02536f
C590 VDD2.n94 B 0.013627f
C591 VDD2.n95 B 0.014429f
C592 VDD2.n96 B 0.03221f
C593 VDD2.n97 B 0.06398f
C594 VDD2.n98 B 0.014429f
C595 VDD2.n99 B 0.013627f
C596 VDD2.n100 B 0.057579f
C597 VDD2.n101 B 0.052695f
C598 VDD2.n102 B 3.00979f
C599 VDD2.t4 B 0.18457f
C600 VDD2.t1 B 0.18457f
C601 VDD2.n103 B 1.61492f
C602 VDD2.n104 B 0.534625f
C603 VDD2.t9 B 0.18457f
C604 VDD2.t7 B 0.18457f
C605 VDD2.n105 B 1.63875f
C606 VN.t3 B 1.58596f
C607 VN.n0 B 0.645687f
C608 VN.n1 B 0.019031f
C609 VN.n2 B 0.015483f
C610 VN.n3 B 0.019031f
C611 VN.t8 B 1.58596f
C612 VN.n4 B 0.566016f
C613 VN.n5 B 0.019031f
C614 VN.n6 B 0.022722f
C615 VN.n7 B 0.019031f
C616 VN.t6 B 1.58596f
C617 VN.n8 B 0.583973f
C618 VN.n9 B 0.019031f
C619 VN.n10 B 0.022722f
C620 VN.n11 B 0.019031f
C621 VN.t0 B 1.58596f
C622 VN.n12 B 0.627737f
C623 VN.t4 B 1.82144f
C624 VN.n13 B 0.596653f
C625 VN.n14 B 0.223645f
C626 VN.n15 B 0.024262f
C627 VN.n16 B 0.035469f
C628 VN.n17 B 0.035802f
C629 VN.n18 B 0.019031f
C630 VN.n19 B 0.019031f
C631 VN.n20 B 0.019031f
C632 VN.n21 B 0.032508f
C633 VN.n22 B 0.035469f
C634 VN.n23 B 0.035469f
C635 VN.n24 B 0.019031f
C636 VN.n25 B 0.019031f
C637 VN.n26 B 0.019031f
C638 VN.n27 B 0.035469f
C639 VN.n28 B 0.035469f
C640 VN.n29 B 0.032508f
C641 VN.n30 B 0.019031f
C642 VN.n31 B 0.019031f
C643 VN.n32 B 0.019031f
C644 VN.n33 B 0.035802f
C645 VN.n34 B 0.035469f
C646 VN.n35 B 0.024262f
C647 VN.n36 B 0.019031f
C648 VN.n37 B 0.019031f
C649 VN.n38 B 0.029165f
C650 VN.n39 B 0.035469f
C651 VN.n40 B 0.038154f
C652 VN.n41 B 0.019031f
C653 VN.n42 B 0.019031f
C654 VN.n43 B 0.019031f
C655 VN.n44 B 0.037395f
C656 VN.n45 B 0.035469f
C657 VN.n46 B 0.030566f
C658 VN.n47 B 0.030715f
C659 VN.n48 B 0.044004f
C660 VN.t1 B 1.58596f
C661 VN.n49 B 0.645687f
C662 VN.n50 B 0.019031f
C663 VN.n51 B 0.015483f
C664 VN.n52 B 0.019031f
C665 VN.t2 B 1.58596f
C666 VN.n53 B 0.566016f
C667 VN.n54 B 0.019031f
C668 VN.n55 B 0.022722f
C669 VN.n56 B 0.019031f
C670 VN.t5 B 1.58596f
C671 VN.n57 B 0.583973f
C672 VN.n58 B 0.019031f
C673 VN.n59 B 0.022722f
C674 VN.n60 B 0.019031f
C675 VN.t9 B 1.58596f
C676 VN.n61 B 0.627737f
C677 VN.t7 B 1.82144f
C678 VN.n62 B 0.596653f
C679 VN.n63 B 0.223645f
C680 VN.n64 B 0.024262f
C681 VN.n65 B 0.035469f
C682 VN.n66 B 0.035802f
C683 VN.n67 B 0.019031f
C684 VN.n68 B 0.019031f
C685 VN.n69 B 0.019031f
C686 VN.n70 B 0.032508f
C687 VN.n71 B 0.035469f
C688 VN.n72 B 0.035469f
C689 VN.n73 B 0.019031f
C690 VN.n74 B 0.019031f
C691 VN.n75 B 0.019031f
C692 VN.n76 B 0.035469f
C693 VN.n77 B 0.035469f
C694 VN.n78 B 0.032508f
C695 VN.n79 B 0.019031f
C696 VN.n80 B 0.019031f
C697 VN.n81 B 0.019031f
C698 VN.n82 B 0.035802f
C699 VN.n83 B 0.035469f
C700 VN.n84 B 0.024262f
C701 VN.n85 B 0.019031f
C702 VN.n86 B 0.019031f
C703 VN.n87 B 0.029165f
C704 VN.n88 B 0.035469f
C705 VN.n89 B 0.038154f
C706 VN.n90 B 0.019031f
C707 VN.n91 B 0.019031f
C708 VN.n92 B 0.019031f
C709 VN.n93 B 0.037395f
C710 VN.n94 B 0.035469f
C711 VN.n95 B 0.030566f
C712 VN.n96 B 0.030715f
C713 VN.n97 B 1.25255f
.ends

