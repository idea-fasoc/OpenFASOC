* NGSPICE file created from diff_pair_sample_0693.ext - technology: sky130A

.subckt diff_pair_sample_0693 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=6.4662 pd=33.94 as=6.4662 ps=33.94 w=16.58 l=3.24
X1 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=6.4662 pd=33.94 as=0 ps=0 w=16.58 l=3.24
X2 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=6.4662 pd=33.94 as=0 ps=0 w=16.58 l=3.24
X3 VDD2.t1 VN.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=6.4662 pd=33.94 as=6.4662 ps=33.94 w=16.58 l=3.24
X4 B.t8 B.t6 B.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=6.4662 pd=33.94 as=0 ps=0 w=16.58 l=3.24
X5 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=6.4662 pd=33.94 as=0 ps=0 w=16.58 l=3.24
X6 VDD2.t0 VN.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=6.4662 pd=33.94 as=6.4662 ps=33.94 w=16.58 l=3.24
X7 VDD1.t0 VP.t1 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=6.4662 pd=33.94 as=6.4662 ps=33.94 w=16.58 l=3.24
R0 VP.n0 VP.t0 211.995
R1 VP.n0 VP.t1 162.173
R2 VP VP.n0 0.526373
R3 VTAIL.n1 VTAIL.t1 47.9802
R4 VTAIL.n2 VTAIL.t3 47.98
R5 VTAIL.n3 VTAIL.t0 47.98
R6 VTAIL.n0 VTAIL.t2 47.98
R7 VTAIL.n1 VTAIL.n0 32.8152
R8 VTAIL.n3 VTAIL.n2 29.7376
R9 VTAIL.n2 VTAIL.n1 2.00912
R10 VTAIL VTAIL.n0 1.29791
R11 VTAIL VTAIL.n3 0.711707
R12 VDD1 VDD1.t0 110.061
R13 VDD1 VDD1.t1 65.4864
R14 B.n845 B.n844 585
R15 B.n358 B.n115 585
R16 B.n357 B.n356 585
R17 B.n355 B.n354 585
R18 B.n353 B.n352 585
R19 B.n351 B.n350 585
R20 B.n349 B.n348 585
R21 B.n347 B.n346 585
R22 B.n345 B.n344 585
R23 B.n343 B.n342 585
R24 B.n341 B.n340 585
R25 B.n339 B.n338 585
R26 B.n337 B.n336 585
R27 B.n335 B.n334 585
R28 B.n333 B.n332 585
R29 B.n331 B.n330 585
R30 B.n329 B.n328 585
R31 B.n327 B.n326 585
R32 B.n325 B.n324 585
R33 B.n323 B.n322 585
R34 B.n321 B.n320 585
R35 B.n319 B.n318 585
R36 B.n317 B.n316 585
R37 B.n315 B.n314 585
R38 B.n313 B.n312 585
R39 B.n311 B.n310 585
R40 B.n309 B.n308 585
R41 B.n307 B.n306 585
R42 B.n305 B.n304 585
R43 B.n303 B.n302 585
R44 B.n301 B.n300 585
R45 B.n299 B.n298 585
R46 B.n297 B.n296 585
R47 B.n295 B.n294 585
R48 B.n293 B.n292 585
R49 B.n291 B.n290 585
R50 B.n289 B.n288 585
R51 B.n287 B.n286 585
R52 B.n285 B.n284 585
R53 B.n283 B.n282 585
R54 B.n281 B.n280 585
R55 B.n279 B.n278 585
R56 B.n277 B.n276 585
R57 B.n275 B.n274 585
R58 B.n273 B.n272 585
R59 B.n271 B.n270 585
R60 B.n269 B.n268 585
R61 B.n267 B.n266 585
R62 B.n265 B.n264 585
R63 B.n263 B.n262 585
R64 B.n261 B.n260 585
R65 B.n259 B.n258 585
R66 B.n257 B.n256 585
R67 B.n255 B.n254 585
R68 B.n253 B.n252 585
R69 B.n250 B.n249 585
R70 B.n248 B.n247 585
R71 B.n246 B.n245 585
R72 B.n244 B.n243 585
R73 B.n242 B.n241 585
R74 B.n240 B.n239 585
R75 B.n238 B.n237 585
R76 B.n236 B.n235 585
R77 B.n234 B.n233 585
R78 B.n232 B.n231 585
R79 B.n229 B.n228 585
R80 B.n227 B.n226 585
R81 B.n225 B.n224 585
R82 B.n223 B.n222 585
R83 B.n221 B.n220 585
R84 B.n219 B.n218 585
R85 B.n217 B.n216 585
R86 B.n215 B.n214 585
R87 B.n213 B.n212 585
R88 B.n211 B.n210 585
R89 B.n209 B.n208 585
R90 B.n207 B.n206 585
R91 B.n205 B.n204 585
R92 B.n203 B.n202 585
R93 B.n201 B.n200 585
R94 B.n199 B.n198 585
R95 B.n197 B.n196 585
R96 B.n195 B.n194 585
R97 B.n193 B.n192 585
R98 B.n191 B.n190 585
R99 B.n189 B.n188 585
R100 B.n187 B.n186 585
R101 B.n185 B.n184 585
R102 B.n183 B.n182 585
R103 B.n181 B.n180 585
R104 B.n179 B.n178 585
R105 B.n177 B.n176 585
R106 B.n175 B.n174 585
R107 B.n173 B.n172 585
R108 B.n171 B.n170 585
R109 B.n169 B.n168 585
R110 B.n167 B.n166 585
R111 B.n165 B.n164 585
R112 B.n163 B.n162 585
R113 B.n161 B.n160 585
R114 B.n159 B.n158 585
R115 B.n157 B.n156 585
R116 B.n155 B.n154 585
R117 B.n153 B.n152 585
R118 B.n151 B.n150 585
R119 B.n149 B.n148 585
R120 B.n147 B.n146 585
R121 B.n145 B.n144 585
R122 B.n143 B.n142 585
R123 B.n141 B.n140 585
R124 B.n139 B.n138 585
R125 B.n137 B.n136 585
R126 B.n135 B.n134 585
R127 B.n133 B.n132 585
R128 B.n131 B.n130 585
R129 B.n129 B.n128 585
R130 B.n127 B.n126 585
R131 B.n125 B.n124 585
R132 B.n123 B.n122 585
R133 B.n121 B.n120 585
R134 B.n843 B.n55 585
R135 B.n848 B.n55 585
R136 B.n842 B.n54 585
R137 B.n849 B.n54 585
R138 B.n841 B.n840 585
R139 B.n840 B.n50 585
R140 B.n839 B.n49 585
R141 B.n855 B.n49 585
R142 B.n838 B.n48 585
R143 B.n856 B.n48 585
R144 B.n837 B.n47 585
R145 B.n857 B.n47 585
R146 B.n836 B.n835 585
R147 B.n835 B.n43 585
R148 B.n834 B.n42 585
R149 B.n863 B.n42 585
R150 B.n833 B.n41 585
R151 B.n864 B.n41 585
R152 B.n832 B.n40 585
R153 B.n865 B.n40 585
R154 B.n831 B.n830 585
R155 B.n830 B.n36 585
R156 B.n829 B.n35 585
R157 B.n871 B.n35 585
R158 B.n828 B.n34 585
R159 B.n872 B.n34 585
R160 B.n827 B.n33 585
R161 B.n873 B.n33 585
R162 B.n826 B.n825 585
R163 B.n825 B.n29 585
R164 B.n824 B.n28 585
R165 B.n879 B.n28 585
R166 B.n823 B.n27 585
R167 B.n880 B.n27 585
R168 B.n822 B.n26 585
R169 B.n881 B.n26 585
R170 B.n821 B.n820 585
R171 B.n820 B.n22 585
R172 B.n819 B.n21 585
R173 B.n887 B.n21 585
R174 B.n818 B.n20 585
R175 B.n888 B.n20 585
R176 B.n817 B.n19 585
R177 B.n889 B.n19 585
R178 B.n816 B.n815 585
R179 B.n815 B.n18 585
R180 B.n814 B.n14 585
R181 B.n895 B.n14 585
R182 B.n813 B.n13 585
R183 B.n896 B.n13 585
R184 B.n812 B.n12 585
R185 B.n897 B.n12 585
R186 B.n811 B.n810 585
R187 B.n810 B.n8 585
R188 B.n809 B.n7 585
R189 B.n903 B.n7 585
R190 B.n808 B.n6 585
R191 B.n904 B.n6 585
R192 B.n807 B.n5 585
R193 B.n905 B.n5 585
R194 B.n806 B.n805 585
R195 B.n805 B.n4 585
R196 B.n804 B.n359 585
R197 B.n804 B.n803 585
R198 B.n794 B.n360 585
R199 B.n361 B.n360 585
R200 B.n796 B.n795 585
R201 B.n797 B.n796 585
R202 B.n793 B.n366 585
R203 B.n366 B.n365 585
R204 B.n792 B.n791 585
R205 B.n791 B.n790 585
R206 B.n368 B.n367 585
R207 B.n783 B.n368 585
R208 B.n782 B.n781 585
R209 B.n784 B.n782 585
R210 B.n780 B.n373 585
R211 B.n373 B.n372 585
R212 B.n779 B.n778 585
R213 B.n778 B.n777 585
R214 B.n375 B.n374 585
R215 B.n376 B.n375 585
R216 B.n770 B.n769 585
R217 B.n771 B.n770 585
R218 B.n768 B.n381 585
R219 B.n381 B.n380 585
R220 B.n767 B.n766 585
R221 B.n766 B.n765 585
R222 B.n383 B.n382 585
R223 B.n384 B.n383 585
R224 B.n758 B.n757 585
R225 B.n759 B.n758 585
R226 B.n756 B.n389 585
R227 B.n389 B.n388 585
R228 B.n755 B.n754 585
R229 B.n754 B.n753 585
R230 B.n391 B.n390 585
R231 B.n392 B.n391 585
R232 B.n746 B.n745 585
R233 B.n747 B.n746 585
R234 B.n744 B.n396 585
R235 B.n400 B.n396 585
R236 B.n743 B.n742 585
R237 B.n742 B.n741 585
R238 B.n398 B.n397 585
R239 B.n399 B.n398 585
R240 B.n734 B.n733 585
R241 B.n735 B.n734 585
R242 B.n732 B.n405 585
R243 B.n405 B.n404 585
R244 B.n731 B.n730 585
R245 B.n730 B.n729 585
R246 B.n407 B.n406 585
R247 B.n408 B.n407 585
R248 B.n722 B.n721 585
R249 B.n723 B.n722 585
R250 B.n720 B.n413 585
R251 B.n413 B.n412 585
R252 B.n715 B.n714 585
R253 B.n713 B.n475 585
R254 B.n712 B.n474 585
R255 B.n717 B.n474 585
R256 B.n711 B.n710 585
R257 B.n709 B.n708 585
R258 B.n707 B.n706 585
R259 B.n705 B.n704 585
R260 B.n703 B.n702 585
R261 B.n701 B.n700 585
R262 B.n699 B.n698 585
R263 B.n697 B.n696 585
R264 B.n695 B.n694 585
R265 B.n693 B.n692 585
R266 B.n691 B.n690 585
R267 B.n689 B.n688 585
R268 B.n687 B.n686 585
R269 B.n685 B.n684 585
R270 B.n683 B.n682 585
R271 B.n681 B.n680 585
R272 B.n679 B.n678 585
R273 B.n677 B.n676 585
R274 B.n675 B.n674 585
R275 B.n673 B.n672 585
R276 B.n671 B.n670 585
R277 B.n669 B.n668 585
R278 B.n667 B.n666 585
R279 B.n665 B.n664 585
R280 B.n663 B.n662 585
R281 B.n661 B.n660 585
R282 B.n659 B.n658 585
R283 B.n657 B.n656 585
R284 B.n655 B.n654 585
R285 B.n653 B.n652 585
R286 B.n651 B.n650 585
R287 B.n649 B.n648 585
R288 B.n647 B.n646 585
R289 B.n645 B.n644 585
R290 B.n643 B.n642 585
R291 B.n641 B.n640 585
R292 B.n639 B.n638 585
R293 B.n637 B.n636 585
R294 B.n635 B.n634 585
R295 B.n633 B.n632 585
R296 B.n631 B.n630 585
R297 B.n629 B.n628 585
R298 B.n627 B.n626 585
R299 B.n625 B.n624 585
R300 B.n623 B.n622 585
R301 B.n621 B.n620 585
R302 B.n619 B.n618 585
R303 B.n617 B.n616 585
R304 B.n615 B.n614 585
R305 B.n613 B.n612 585
R306 B.n611 B.n610 585
R307 B.n609 B.n608 585
R308 B.n607 B.n606 585
R309 B.n605 B.n604 585
R310 B.n603 B.n602 585
R311 B.n601 B.n600 585
R312 B.n599 B.n598 585
R313 B.n597 B.n596 585
R314 B.n595 B.n594 585
R315 B.n593 B.n592 585
R316 B.n591 B.n590 585
R317 B.n589 B.n588 585
R318 B.n587 B.n586 585
R319 B.n585 B.n584 585
R320 B.n583 B.n582 585
R321 B.n581 B.n580 585
R322 B.n579 B.n578 585
R323 B.n577 B.n576 585
R324 B.n575 B.n574 585
R325 B.n573 B.n572 585
R326 B.n571 B.n570 585
R327 B.n569 B.n568 585
R328 B.n567 B.n566 585
R329 B.n565 B.n564 585
R330 B.n563 B.n562 585
R331 B.n561 B.n560 585
R332 B.n559 B.n558 585
R333 B.n557 B.n556 585
R334 B.n555 B.n554 585
R335 B.n553 B.n552 585
R336 B.n551 B.n550 585
R337 B.n549 B.n548 585
R338 B.n547 B.n546 585
R339 B.n545 B.n544 585
R340 B.n543 B.n542 585
R341 B.n541 B.n540 585
R342 B.n539 B.n538 585
R343 B.n537 B.n536 585
R344 B.n535 B.n534 585
R345 B.n533 B.n532 585
R346 B.n531 B.n530 585
R347 B.n529 B.n528 585
R348 B.n527 B.n526 585
R349 B.n525 B.n524 585
R350 B.n523 B.n522 585
R351 B.n521 B.n520 585
R352 B.n519 B.n518 585
R353 B.n517 B.n516 585
R354 B.n515 B.n514 585
R355 B.n513 B.n512 585
R356 B.n511 B.n510 585
R357 B.n509 B.n508 585
R358 B.n507 B.n506 585
R359 B.n505 B.n504 585
R360 B.n503 B.n502 585
R361 B.n501 B.n500 585
R362 B.n499 B.n498 585
R363 B.n497 B.n496 585
R364 B.n495 B.n494 585
R365 B.n493 B.n492 585
R366 B.n491 B.n490 585
R367 B.n489 B.n488 585
R368 B.n487 B.n486 585
R369 B.n485 B.n484 585
R370 B.n483 B.n482 585
R371 B.n415 B.n414 585
R372 B.n719 B.n718 585
R373 B.n718 B.n717 585
R374 B.n411 B.n410 585
R375 B.n412 B.n411 585
R376 B.n725 B.n724 585
R377 B.n724 B.n723 585
R378 B.n726 B.n409 585
R379 B.n409 B.n408 585
R380 B.n728 B.n727 585
R381 B.n729 B.n728 585
R382 B.n403 B.n402 585
R383 B.n404 B.n403 585
R384 B.n737 B.n736 585
R385 B.n736 B.n735 585
R386 B.n738 B.n401 585
R387 B.n401 B.n399 585
R388 B.n740 B.n739 585
R389 B.n741 B.n740 585
R390 B.n395 B.n394 585
R391 B.n400 B.n395 585
R392 B.n749 B.n748 585
R393 B.n748 B.n747 585
R394 B.n750 B.n393 585
R395 B.n393 B.n392 585
R396 B.n752 B.n751 585
R397 B.n753 B.n752 585
R398 B.n387 B.n386 585
R399 B.n388 B.n387 585
R400 B.n761 B.n760 585
R401 B.n760 B.n759 585
R402 B.n762 B.n385 585
R403 B.n385 B.n384 585
R404 B.n764 B.n763 585
R405 B.n765 B.n764 585
R406 B.n379 B.n378 585
R407 B.n380 B.n379 585
R408 B.n773 B.n772 585
R409 B.n772 B.n771 585
R410 B.n774 B.n377 585
R411 B.n377 B.n376 585
R412 B.n776 B.n775 585
R413 B.n777 B.n776 585
R414 B.n371 B.n370 585
R415 B.n372 B.n371 585
R416 B.n786 B.n785 585
R417 B.n785 B.n784 585
R418 B.n787 B.n369 585
R419 B.n783 B.n369 585
R420 B.n789 B.n788 585
R421 B.n790 B.n789 585
R422 B.n364 B.n363 585
R423 B.n365 B.n364 585
R424 B.n799 B.n798 585
R425 B.n798 B.n797 585
R426 B.n800 B.n362 585
R427 B.n362 B.n361 585
R428 B.n802 B.n801 585
R429 B.n803 B.n802 585
R430 B.n2 B.n0 585
R431 B.n4 B.n2 585
R432 B.n3 B.n1 585
R433 B.n904 B.n3 585
R434 B.n902 B.n901 585
R435 B.n903 B.n902 585
R436 B.n900 B.n9 585
R437 B.n9 B.n8 585
R438 B.n899 B.n898 585
R439 B.n898 B.n897 585
R440 B.n11 B.n10 585
R441 B.n896 B.n11 585
R442 B.n894 B.n893 585
R443 B.n895 B.n894 585
R444 B.n892 B.n15 585
R445 B.n18 B.n15 585
R446 B.n891 B.n890 585
R447 B.n890 B.n889 585
R448 B.n17 B.n16 585
R449 B.n888 B.n17 585
R450 B.n886 B.n885 585
R451 B.n887 B.n886 585
R452 B.n884 B.n23 585
R453 B.n23 B.n22 585
R454 B.n883 B.n882 585
R455 B.n882 B.n881 585
R456 B.n25 B.n24 585
R457 B.n880 B.n25 585
R458 B.n878 B.n877 585
R459 B.n879 B.n878 585
R460 B.n876 B.n30 585
R461 B.n30 B.n29 585
R462 B.n875 B.n874 585
R463 B.n874 B.n873 585
R464 B.n32 B.n31 585
R465 B.n872 B.n32 585
R466 B.n870 B.n869 585
R467 B.n871 B.n870 585
R468 B.n868 B.n37 585
R469 B.n37 B.n36 585
R470 B.n867 B.n866 585
R471 B.n866 B.n865 585
R472 B.n39 B.n38 585
R473 B.n864 B.n39 585
R474 B.n862 B.n861 585
R475 B.n863 B.n862 585
R476 B.n860 B.n44 585
R477 B.n44 B.n43 585
R478 B.n859 B.n858 585
R479 B.n858 B.n857 585
R480 B.n46 B.n45 585
R481 B.n856 B.n46 585
R482 B.n854 B.n853 585
R483 B.n855 B.n854 585
R484 B.n852 B.n51 585
R485 B.n51 B.n50 585
R486 B.n851 B.n850 585
R487 B.n850 B.n849 585
R488 B.n53 B.n52 585
R489 B.n848 B.n53 585
R490 B.n907 B.n906 585
R491 B.n906 B.n905 585
R492 B.n715 B.n411 497.305
R493 B.n120 B.n53 497.305
R494 B.n718 B.n413 497.305
R495 B.n845 B.n55 497.305
R496 B.n479 B.t6 332.171
R497 B.n476 B.t2 332.171
R498 B.n118 B.t13 332.171
R499 B.n116 B.t9 332.171
R500 B.n847 B.n846 256.663
R501 B.n847 B.n114 256.663
R502 B.n847 B.n113 256.663
R503 B.n847 B.n112 256.663
R504 B.n847 B.n111 256.663
R505 B.n847 B.n110 256.663
R506 B.n847 B.n109 256.663
R507 B.n847 B.n108 256.663
R508 B.n847 B.n107 256.663
R509 B.n847 B.n106 256.663
R510 B.n847 B.n105 256.663
R511 B.n847 B.n104 256.663
R512 B.n847 B.n103 256.663
R513 B.n847 B.n102 256.663
R514 B.n847 B.n101 256.663
R515 B.n847 B.n100 256.663
R516 B.n847 B.n99 256.663
R517 B.n847 B.n98 256.663
R518 B.n847 B.n97 256.663
R519 B.n847 B.n96 256.663
R520 B.n847 B.n95 256.663
R521 B.n847 B.n94 256.663
R522 B.n847 B.n93 256.663
R523 B.n847 B.n92 256.663
R524 B.n847 B.n91 256.663
R525 B.n847 B.n90 256.663
R526 B.n847 B.n89 256.663
R527 B.n847 B.n88 256.663
R528 B.n847 B.n87 256.663
R529 B.n847 B.n86 256.663
R530 B.n847 B.n85 256.663
R531 B.n847 B.n84 256.663
R532 B.n847 B.n83 256.663
R533 B.n847 B.n82 256.663
R534 B.n847 B.n81 256.663
R535 B.n847 B.n80 256.663
R536 B.n847 B.n79 256.663
R537 B.n847 B.n78 256.663
R538 B.n847 B.n77 256.663
R539 B.n847 B.n76 256.663
R540 B.n847 B.n75 256.663
R541 B.n847 B.n74 256.663
R542 B.n847 B.n73 256.663
R543 B.n847 B.n72 256.663
R544 B.n847 B.n71 256.663
R545 B.n847 B.n70 256.663
R546 B.n847 B.n69 256.663
R547 B.n847 B.n68 256.663
R548 B.n847 B.n67 256.663
R549 B.n847 B.n66 256.663
R550 B.n847 B.n65 256.663
R551 B.n847 B.n64 256.663
R552 B.n847 B.n63 256.663
R553 B.n847 B.n62 256.663
R554 B.n847 B.n61 256.663
R555 B.n847 B.n60 256.663
R556 B.n847 B.n59 256.663
R557 B.n847 B.n58 256.663
R558 B.n847 B.n57 256.663
R559 B.n847 B.n56 256.663
R560 B.n717 B.n716 256.663
R561 B.n717 B.n416 256.663
R562 B.n717 B.n417 256.663
R563 B.n717 B.n418 256.663
R564 B.n717 B.n419 256.663
R565 B.n717 B.n420 256.663
R566 B.n717 B.n421 256.663
R567 B.n717 B.n422 256.663
R568 B.n717 B.n423 256.663
R569 B.n717 B.n424 256.663
R570 B.n717 B.n425 256.663
R571 B.n717 B.n426 256.663
R572 B.n717 B.n427 256.663
R573 B.n717 B.n428 256.663
R574 B.n717 B.n429 256.663
R575 B.n717 B.n430 256.663
R576 B.n717 B.n431 256.663
R577 B.n717 B.n432 256.663
R578 B.n717 B.n433 256.663
R579 B.n717 B.n434 256.663
R580 B.n717 B.n435 256.663
R581 B.n717 B.n436 256.663
R582 B.n717 B.n437 256.663
R583 B.n717 B.n438 256.663
R584 B.n717 B.n439 256.663
R585 B.n717 B.n440 256.663
R586 B.n717 B.n441 256.663
R587 B.n717 B.n442 256.663
R588 B.n717 B.n443 256.663
R589 B.n717 B.n444 256.663
R590 B.n717 B.n445 256.663
R591 B.n717 B.n446 256.663
R592 B.n717 B.n447 256.663
R593 B.n717 B.n448 256.663
R594 B.n717 B.n449 256.663
R595 B.n717 B.n450 256.663
R596 B.n717 B.n451 256.663
R597 B.n717 B.n452 256.663
R598 B.n717 B.n453 256.663
R599 B.n717 B.n454 256.663
R600 B.n717 B.n455 256.663
R601 B.n717 B.n456 256.663
R602 B.n717 B.n457 256.663
R603 B.n717 B.n458 256.663
R604 B.n717 B.n459 256.663
R605 B.n717 B.n460 256.663
R606 B.n717 B.n461 256.663
R607 B.n717 B.n462 256.663
R608 B.n717 B.n463 256.663
R609 B.n717 B.n464 256.663
R610 B.n717 B.n465 256.663
R611 B.n717 B.n466 256.663
R612 B.n717 B.n467 256.663
R613 B.n717 B.n468 256.663
R614 B.n717 B.n469 256.663
R615 B.n717 B.n470 256.663
R616 B.n717 B.n471 256.663
R617 B.n717 B.n472 256.663
R618 B.n717 B.n473 256.663
R619 B.n724 B.n411 163.367
R620 B.n724 B.n409 163.367
R621 B.n728 B.n409 163.367
R622 B.n728 B.n403 163.367
R623 B.n736 B.n403 163.367
R624 B.n736 B.n401 163.367
R625 B.n740 B.n401 163.367
R626 B.n740 B.n395 163.367
R627 B.n748 B.n395 163.367
R628 B.n748 B.n393 163.367
R629 B.n752 B.n393 163.367
R630 B.n752 B.n387 163.367
R631 B.n760 B.n387 163.367
R632 B.n760 B.n385 163.367
R633 B.n764 B.n385 163.367
R634 B.n764 B.n379 163.367
R635 B.n772 B.n379 163.367
R636 B.n772 B.n377 163.367
R637 B.n776 B.n377 163.367
R638 B.n776 B.n371 163.367
R639 B.n785 B.n371 163.367
R640 B.n785 B.n369 163.367
R641 B.n789 B.n369 163.367
R642 B.n789 B.n364 163.367
R643 B.n798 B.n364 163.367
R644 B.n798 B.n362 163.367
R645 B.n802 B.n362 163.367
R646 B.n802 B.n2 163.367
R647 B.n906 B.n2 163.367
R648 B.n906 B.n3 163.367
R649 B.n902 B.n3 163.367
R650 B.n902 B.n9 163.367
R651 B.n898 B.n9 163.367
R652 B.n898 B.n11 163.367
R653 B.n894 B.n11 163.367
R654 B.n894 B.n15 163.367
R655 B.n890 B.n15 163.367
R656 B.n890 B.n17 163.367
R657 B.n886 B.n17 163.367
R658 B.n886 B.n23 163.367
R659 B.n882 B.n23 163.367
R660 B.n882 B.n25 163.367
R661 B.n878 B.n25 163.367
R662 B.n878 B.n30 163.367
R663 B.n874 B.n30 163.367
R664 B.n874 B.n32 163.367
R665 B.n870 B.n32 163.367
R666 B.n870 B.n37 163.367
R667 B.n866 B.n37 163.367
R668 B.n866 B.n39 163.367
R669 B.n862 B.n39 163.367
R670 B.n862 B.n44 163.367
R671 B.n858 B.n44 163.367
R672 B.n858 B.n46 163.367
R673 B.n854 B.n46 163.367
R674 B.n854 B.n51 163.367
R675 B.n850 B.n51 163.367
R676 B.n850 B.n53 163.367
R677 B.n475 B.n474 163.367
R678 B.n710 B.n474 163.367
R679 B.n708 B.n707 163.367
R680 B.n704 B.n703 163.367
R681 B.n700 B.n699 163.367
R682 B.n696 B.n695 163.367
R683 B.n692 B.n691 163.367
R684 B.n688 B.n687 163.367
R685 B.n684 B.n683 163.367
R686 B.n680 B.n679 163.367
R687 B.n676 B.n675 163.367
R688 B.n672 B.n671 163.367
R689 B.n668 B.n667 163.367
R690 B.n664 B.n663 163.367
R691 B.n660 B.n659 163.367
R692 B.n656 B.n655 163.367
R693 B.n652 B.n651 163.367
R694 B.n648 B.n647 163.367
R695 B.n644 B.n643 163.367
R696 B.n640 B.n639 163.367
R697 B.n636 B.n635 163.367
R698 B.n632 B.n631 163.367
R699 B.n628 B.n627 163.367
R700 B.n624 B.n623 163.367
R701 B.n620 B.n619 163.367
R702 B.n616 B.n615 163.367
R703 B.n612 B.n611 163.367
R704 B.n608 B.n607 163.367
R705 B.n604 B.n603 163.367
R706 B.n600 B.n599 163.367
R707 B.n596 B.n595 163.367
R708 B.n592 B.n591 163.367
R709 B.n588 B.n587 163.367
R710 B.n584 B.n583 163.367
R711 B.n580 B.n579 163.367
R712 B.n576 B.n575 163.367
R713 B.n572 B.n571 163.367
R714 B.n568 B.n567 163.367
R715 B.n564 B.n563 163.367
R716 B.n560 B.n559 163.367
R717 B.n556 B.n555 163.367
R718 B.n552 B.n551 163.367
R719 B.n548 B.n547 163.367
R720 B.n544 B.n543 163.367
R721 B.n540 B.n539 163.367
R722 B.n536 B.n535 163.367
R723 B.n532 B.n531 163.367
R724 B.n528 B.n527 163.367
R725 B.n524 B.n523 163.367
R726 B.n520 B.n519 163.367
R727 B.n516 B.n515 163.367
R728 B.n512 B.n511 163.367
R729 B.n508 B.n507 163.367
R730 B.n504 B.n503 163.367
R731 B.n500 B.n499 163.367
R732 B.n496 B.n495 163.367
R733 B.n492 B.n491 163.367
R734 B.n488 B.n487 163.367
R735 B.n484 B.n483 163.367
R736 B.n718 B.n415 163.367
R737 B.n722 B.n413 163.367
R738 B.n722 B.n407 163.367
R739 B.n730 B.n407 163.367
R740 B.n730 B.n405 163.367
R741 B.n734 B.n405 163.367
R742 B.n734 B.n398 163.367
R743 B.n742 B.n398 163.367
R744 B.n742 B.n396 163.367
R745 B.n746 B.n396 163.367
R746 B.n746 B.n391 163.367
R747 B.n754 B.n391 163.367
R748 B.n754 B.n389 163.367
R749 B.n758 B.n389 163.367
R750 B.n758 B.n383 163.367
R751 B.n766 B.n383 163.367
R752 B.n766 B.n381 163.367
R753 B.n770 B.n381 163.367
R754 B.n770 B.n375 163.367
R755 B.n778 B.n375 163.367
R756 B.n778 B.n373 163.367
R757 B.n782 B.n373 163.367
R758 B.n782 B.n368 163.367
R759 B.n791 B.n368 163.367
R760 B.n791 B.n366 163.367
R761 B.n796 B.n366 163.367
R762 B.n796 B.n360 163.367
R763 B.n804 B.n360 163.367
R764 B.n805 B.n804 163.367
R765 B.n805 B.n5 163.367
R766 B.n6 B.n5 163.367
R767 B.n7 B.n6 163.367
R768 B.n810 B.n7 163.367
R769 B.n810 B.n12 163.367
R770 B.n13 B.n12 163.367
R771 B.n14 B.n13 163.367
R772 B.n815 B.n14 163.367
R773 B.n815 B.n19 163.367
R774 B.n20 B.n19 163.367
R775 B.n21 B.n20 163.367
R776 B.n820 B.n21 163.367
R777 B.n820 B.n26 163.367
R778 B.n27 B.n26 163.367
R779 B.n28 B.n27 163.367
R780 B.n825 B.n28 163.367
R781 B.n825 B.n33 163.367
R782 B.n34 B.n33 163.367
R783 B.n35 B.n34 163.367
R784 B.n830 B.n35 163.367
R785 B.n830 B.n40 163.367
R786 B.n41 B.n40 163.367
R787 B.n42 B.n41 163.367
R788 B.n835 B.n42 163.367
R789 B.n835 B.n47 163.367
R790 B.n48 B.n47 163.367
R791 B.n49 B.n48 163.367
R792 B.n840 B.n49 163.367
R793 B.n840 B.n54 163.367
R794 B.n55 B.n54 163.367
R795 B.n124 B.n123 163.367
R796 B.n128 B.n127 163.367
R797 B.n132 B.n131 163.367
R798 B.n136 B.n135 163.367
R799 B.n140 B.n139 163.367
R800 B.n144 B.n143 163.367
R801 B.n148 B.n147 163.367
R802 B.n152 B.n151 163.367
R803 B.n156 B.n155 163.367
R804 B.n160 B.n159 163.367
R805 B.n164 B.n163 163.367
R806 B.n168 B.n167 163.367
R807 B.n172 B.n171 163.367
R808 B.n176 B.n175 163.367
R809 B.n180 B.n179 163.367
R810 B.n184 B.n183 163.367
R811 B.n188 B.n187 163.367
R812 B.n192 B.n191 163.367
R813 B.n196 B.n195 163.367
R814 B.n200 B.n199 163.367
R815 B.n204 B.n203 163.367
R816 B.n208 B.n207 163.367
R817 B.n212 B.n211 163.367
R818 B.n216 B.n215 163.367
R819 B.n220 B.n219 163.367
R820 B.n224 B.n223 163.367
R821 B.n228 B.n227 163.367
R822 B.n233 B.n232 163.367
R823 B.n237 B.n236 163.367
R824 B.n241 B.n240 163.367
R825 B.n245 B.n244 163.367
R826 B.n249 B.n248 163.367
R827 B.n254 B.n253 163.367
R828 B.n258 B.n257 163.367
R829 B.n262 B.n261 163.367
R830 B.n266 B.n265 163.367
R831 B.n270 B.n269 163.367
R832 B.n274 B.n273 163.367
R833 B.n278 B.n277 163.367
R834 B.n282 B.n281 163.367
R835 B.n286 B.n285 163.367
R836 B.n290 B.n289 163.367
R837 B.n294 B.n293 163.367
R838 B.n298 B.n297 163.367
R839 B.n302 B.n301 163.367
R840 B.n306 B.n305 163.367
R841 B.n310 B.n309 163.367
R842 B.n314 B.n313 163.367
R843 B.n318 B.n317 163.367
R844 B.n322 B.n321 163.367
R845 B.n326 B.n325 163.367
R846 B.n330 B.n329 163.367
R847 B.n334 B.n333 163.367
R848 B.n338 B.n337 163.367
R849 B.n342 B.n341 163.367
R850 B.n346 B.n345 163.367
R851 B.n350 B.n349 163.367
R852 B.n354 B.n353 163.367
R853 B.n356 B.n115 163.367
R854 B.n479 B.t8 141.619
R855 B.n116 B.t11 141.619
R856 B.n476 B.t5 141.597
R857 B.n118 B.t14 141.597
R858 B.n480 B.t7 72.383
R859 B.n117 B.t12 72.383
R860 B.n477 B.t4 72.3613
R861 B.n119 B.t15 72.3613
R862 B.n716 B.n715 71.676
R863 B.n710 B.n416 71.676
R864 B.n707 B.n417 71.676
R865 B.n703 B.n418 71.676
R866 B.n699 B.n419 71.676
R867 B.n695 B.n420 71.676
R868 B.n691 B.n421 71.676
R869 B.n687 B.n422 71.676
R870 B.n683 B.n423 71.676
R871 B.n679 B.n424 71.676
R872 B.n675 B.n425 71.676
R873 B.n671 B.n426 71.676
R874 B.n667 B.n427 71.676
R875 B.n663 B.n428 71.676
R876 B.n659 B.n429 71.676
R877 B.n655 B.n430 71.676
R878 B.n651 B.n431 71.676
R879 B.n647 B.n432 71.676
R880 B.n643 B.n433 71.676
R881 B.n639 B.n434 71.676
R882 B.n635 B.n435 71.676
R883 B.n631 B.n436 71.676
R884 B.n627 B.n437 71.676
R885 B.n623 B.n438 71.676
R886 B.n619 B.n439 71.676
R887 B.n615 B.n440 71.676
R888 B.n611 B.n441 71.676
R889 B.n607 B.n442 71.676
R890 B.n603 B.n443 71.676
R891 B.n599 B.n444 71.676
R892 B.n595 B.n445 71.676
R893 B.n591 B.n446 71.676
R894 B.n587 B.n447 71.676
R895 B.n583 B.n448 71.676
R896 B.n579 B.n449 71.676
R897 B.n575 B.n450 71.676
R898 B.n571 B.n451 71.676
R899 B.n567 B.n452 71.676
R900 B.n563 B.n453 71.676
R901 B.n559 B.n454 71.676
R902 B.n555 B.n455 71.676
R903 B.n551 B.n456 71.676
R904 B.n547 B.n457 71.676
R905 B.n543 B.n458 71.676
R906 B.n539 B.n459 71.676
R907 B.n535 B.n460 71.676
R908 B.n531 B.n461 71.676
R909 B.n527 B.n462 71.676
R910 B.n523 B.n463 71.676
R911 B.n519 B.n464 71.676
R912 B.n515 B.n465 71.676
R913 B.n511 B.n466 71.676
R914 B.n507 B.n467 71.676
R915 B.n503 B.n468 71.676
R916 B.n499 B.n469 71.676
R917 B.n495 B.n470 71.676
R918 B.n491 B.n471 71.676
R919 B.n487 B.n472 71.676
R920 B.n483 B.n473 71.676
R921 B.n120 B.n56 71.676
R922 B.n124 B.n57 71.676
R923 B.n128 B.n58 71.676
R924 B.n132 B.n59 71.676
R925 B.n136 B.n60 71.676
R926 B.n140 B.n61 71.676
R927 B.n144 B.n62 71.676
R928 B.n148 B.n63 71.676
R929 B.n152 B.n64 71.676
R930 B.n156 B.n65 71.676
R931 B.n160 B.n66 71.676
R932 B.n164 B.n67 71.676
R933 B.n168 B.n68 71.676
R934 B.n172 B.n69 71.676
R935 B.n176 B.n70 71.676
R936 B.n180 B.n71 71.676
R937 B.n184 B.n72 71.676
R938 B.n188 B.n73 71.676
R939 B.n192 B.n74 71.676
R940 B.n196 B.n75 71.676
R941 B.n200 B.n76 71.676
R942 B.n204 B.n77 71.676
R943 B.n208 B.n78 71.676
R944 B.n212 B.n79 71.676
R945 B.n216 B.n80 71.676
R946 B.n220 B.n81 71.676
R947 B.n224 B.n82 71.676
R948 B.n228 B.n83 71.676
R949 B.n233 B.n84 71.676
R950 B.n237 B.n85 71.676
R951 B.n241 B.n86 71.676
R952 B.n245 B.n87 71.676
R953 B.n249 B.n88 71.676
R954 B.n254 B.n89 71.676
R955 B.n258 B.n90 71.676
R956 B.n262 B.n91 71.676
R957 B.n266 B.n92 71.676
R958 B.n270 B.n93 71.676
R959 B.n274 B.n94 71.676
R960 B.n278 B.n95 71.676
R961 B.n282 B.n96 71.676
R962 B.n286 B.n97 71.676
R963 B.n290 B.n98 71.676
R964 B.n294 B.n99 71.676
R965 B.n298 B.n100 71.676
R966 B.n302 B.n101 71.676
R967 B.n306 B.n102 71.676
R968 B.n310 B.n103 71.676
R969 B.n314 B.n104 71.676
R970 B.n318 B.n105 71.676
R971 B.n322 B.n106 71.676
R972 B.n326 B.n107 71.676
R973 B.n330 B.n108 71.676
R974 B.n334 B.n109 71.676
R975 B.n338 B.n110 71.676
R976 B.n342 B.n111 71.676
R977 B.n346 B.n112 71.676
R978 B.n350 B.n113 71.676
R979 B.n354 B.n114 71.676
R980 B.n846 B.n115 71.676
R981 B.n846 B.n845 71.676
R982 B.n356 B.n114 71.676
R983 B.n353 B.n113 71.676
R984 B.n349 B.n112 71.676
R985 B.n345 B.n111 71.676
R986 B.n341 B.n110 71.676
R987 B.n337 B.n109 71.676
R988 B.n333 B.n108 71.676
R989 B.n329 B.n107 71.676
R990 B.n325 B.n106 71.676
R991 B.n321 B.n105 71.676
R992 B.n317 B.n104 71.676
R993 B.n313 B.n103 71.676
R994 B.n309 B.n102 71.676
R995 B.n305 B.n101 71.676
R996 B.n301 B.n100 71.676
R997 B.n297 B.n99 71.676
R998 B.n293 B.n98 71.676
R999 B.n289 B.n97 71.676
R1000 B.n285 B.n96 71.676
R1001 B.n281 B.n95 71.676
R1002 B.n277 B.n94 71.676
R1003 B.n273 B.n93 71.676
R1004 B.n269 B.n92 71.676
R1005 B.n265 B.n91 71.676
R1006 B.n261 B.n90 71.676
R1007 B.n257 B.n89 71.676
R1008 B.n253 B.n88 71.676
R1009 B.n248 B.n87 71.676
R1010 B.n244 B.n86 71.676
R1011 B.n240 B.n85 71.676
R1012 B.n236 B.n84 71.676
R1013 B.n232 B.n83 71.676
R1014 B.n227 B.n82 71.676
R1015 B.n223 B.n81 71.676
R1016 B.n219 B.n80 71.676
R1017 B.n215 B.n79 71.676
R1018 B.n211 B.n78 71.676
R1019 B.n207 B.n77 71.676
R1020 B.n203 B.n76 71.676
R1021 B.n199 B.n75 71.676
R1022 B.n195 B.n74 71.676
R1023 B.n191 B.n73 71.676
R1024 B.n187 B.n72 71.676
R1025 B.n183 B.n71 71.676
R1026 B.n179 B.n70 71.676
R1027 B.n175 B.n69 71.676
R1028 B.n171 B.n68 71.676
R1029 B.n167 B.n67 71.676
R1030 B.n163 B.n66 71.676
R1031 B.n159 B.n65 71.676
R1032 B.n155 B.n64 71.676
R1033 B.n151 B.n63 71.676
R1034 B.n147 B.n62 71.676
R1035 B.n143 B.n61 71.676
R1036 B.n139 B.n60 71.676
R1037 B.n135 B.n59 71.676
R1038 B.n131 B.n58 71.676
R1039 B.n127 B.n57 71.676
R1040 B.n123 B.n56 71.676
R1041 B.n716 B.n475 71.676
R1042 B.n708 B.n416 71.676
R1043 B.n704 B.n417 71.676
R1044 B.n700 B.n418 71.676
R1045 B.n696 B.n419 71.676
R1046 B.n692 B.n420 71.676
R1047 B.n688 B.n421 71.676
R1048 B.n684 B.n422 71.676
R1049 B.n680 B.n423 71.676
R1050 B.n676 B.n424 71.676
R1051 B.n672 B.n425 71.676
R1052 B.n668 B.n426 71.676
R1053 B.n664 B.n427 71.676
R1054 B.n660 B.n428 71.676
R1055 B.n656 B.n429 71.676
R1056 B.n652 B.n430 71.676
R1057 B.n648 B.n431 71.676
R1058 B.n644 B.n432 71.676
R1059 B.n640 B.n433 71.676
R1060 B.n636 B.n434 71.676
R1061 B.n632 B.n435 71.676
R1062 B.n628 B.n436 71.676
R1063 B.n624 B.n437 71.676
R1064 B.n620 B.n438 71.676
R1065 B.n616 B.n439 71.676
R1066 B.n612 B.n440 71.676
R1067 B.n608 B.n441 71.676
R1068 B.n604 B.n442 71.676
R1069 B.n600 B.n443 71.676
R1070 B.n596 B.n444 71.676
R1071 B.n592 B.n445 71.676
R1072 B.n588 B.n446 71.676
R1073 B.n584 B.n447 71.676
R1074 B.n580 B.n448 71.676
R1075 B.n576 B.n449 71.676
R1076 B.n572 B.n450 71.676
R1077 B.n568 B.n451 71.676
R1078 B.n564 B.n452 71.676
R1079 B.n560 B.n453 71.676
R1080 B.n556 B.n454 71.676
R1081 B.n552 B.n455 71.676
R1082 B.n548 B.n456 71.676
R1083 B.n544 B.n457 71.676
R1084 B.n540 B.n458 71.676
R1085 B.n536 B.n459 71.676
R1086 B.n532 B.n460 71.676
R1087 B.n528 B.n461 71.676
R1088 B.n524 B.n462 71.676
R1089 B.n520 B.n463 71.676
R1090 B.n516 B.n464 71.676
R1091 B.n512 B.n465 71.676
R1092 B.n508 B.n466 71.676
R1093 B.n504 B.n467 71.676
R1094 B.n500 B.n468 71.676
R1095 B.n496 B.n469 71.676
R1096 B.n492 B.n470 71.676
R1097 B.n488 B.n471 71.676
R1098 B.n484 B.n472 71.676
R1099 B.n473 B.n415 71.676
R1100 B.n480 B.n479 69.2369
R1101 B.n477 B.n476 69.2369
R1102 B.n119 B.n118 69.2369
R1103 B.n117 B.n116 69.2369
R1104 B.n717 B.n412 65.9351
R1105 B.n848 B.n847 65.9351
R1106 B.n481 B.n480 59.5399
R1107 B.n478 B.n477 59.5399
R1108 B.n230 B.n119 59.5399
R1109 B.n251 B.n117 59.5399
R1110 B.n723 B.n412 34.2261
R1111 B.n723 B.n408 34.2261
R1112 B.n729 B.n408 34.2261
R1113 B.n729 B.n404 34.2261
R1114 B.n735 B.n404 34.2261
R1115 B.n735 B.n399 34.2261
R1116 B.n741 B.n399 34.2261
R1117 B.n741 B.n400 34.2261
R1118 B.n747 B.n392 34.2261
R1119 B.n753 B.n392 34.2261
R1120 B.n753 B.n388 34.2261
R1121 B.n759 B.n388 34.2261
R1122 B.n759 B.n384 34.2261
R1123 B.n765 B.n384 34.2261
R1124 B.n765 B.n380 34.2261
R1125 B.n771 B.n380 34.2261
R1126 B.n771 B.n376 34.2261
R1127 B.n777 B.n376 34.2261
R1128 B.n777 B.n372 34.2261
R1129 B.n784 B.n372 34.2261
R1130 B.n784 B.n783 34.2261
R1131 B.n790 B.n365 34.2261
R1132 B.n797 B.n365 34.2261
R1133 B.n797 B.n361 34.2261
R1134 B.n803 B.n361 34.2261
R1135 B.n803 B.n4 34.2261
R1136 B.n905 B.n4 34.2261
R1137 B.n905 B.n904 34.2261
R1138 B.n904 B.n903 34.2261
R1139 B.n903 B.n8 34.2261
R1140 B.n897 B.n8 34.2261
R1141 B.n897 B.n896 34.2261
R1142 B.n896 B.n895 34.2261
R1143 B.n889 B.n18 34.2261
R1144 B.n889 B.n888 34.2261
R1145 B.n888 B.n887 34.2261
R1146 B.n887 B.n22 34.2261
R1147 B.n881 B.n22 34.2261
R1148 B.n881 B.n880 34.2261
R1149 B.n880 B.n879 34.2261
R1150 B.n879 B.n29 34.2261
R1151 B.n873 B.n29 34.2261
R1152 B.n873 B.n872 34.2261
R1153 B.n872 B.n871 34.2261
R1154 B.n871 B.n36 34.2261
R1155 B.n865 B.n36 34.2261
R1156 B.n864 B.n863 34.2261
R1157 B.n863 B.n43 34.2261
R1158 B.n857 B.n43 34.2261
R1159 B.n857 B.n856 34.2261
R1160 B.n856 B.n855 34.2261
R1161 B.n855 B.n50 34.2261
R1162 B.n849 B.n50 34.2261
R1163 B.n849 B.n848 34.2261
R1164 B.n121 B.n52 32.3127
R1165 B.n844 B.n843 32.3127
R1166 B.n720 B.n719 32.3127
R1167 B.n714 B.n410 32.3127
R1168 B.n790 B.t1 29.1929
R1169 B.n895 B.t0 29.1929
R1170 B.n747 B.t3 19.1266
R1171 B.n865 B.t10 19.1266
R1172 B B.n907 18.0485
R1173 B.n400 B.t3 15.1
R1174 B.t10 B.n864 15.1
R1175 B.n122 B.n121 10.6151
R1176 B.n125 B.n122 10.6151
R1177 B.n126 B.n125 10.6151
R1178 B.n129 B.n126 10.6151
R1179 B.n130 B.n129 10.6151
R1180 B.n133 B.n130 10.6151
R1181 B.n134 B.n133 10.6151
R1182 B.n137 B.n134 10.6151
R1183 B.n138 B.n137 10.6151
R1184 B.n141 B.n138 10.6151
R1185 B.n142 B.n141 10.6151
R1186 B.n145 B.n142 10.6151
R1187 B.n146 B.n145 10.6151
R1188 B.n149 B.n146 10.6151
R1189 B.n150 B.n149 10.6151
R1190 B.n153 B.n150 10.6151
R1191 B.n154 B.n153 10.6151
R1192 B.n157 B.n154 10.6151
R1193 B.n158 B.n157 10.6151
R1194 B.n161 B.n158 10.6151
R1195 B.n162 B.n161 10.6151
R1196 B.n165 B.n162 10.6151
R1197 B.n166 B.n165 10.6151
R1198 B.n169 B.n166 10.6151
R1199 B.n170 B.n169 10.6151
R1200 B.n173 B.n170 10.6151
R1201 B.n174 B.n173 10.6151
R1202 B.n177 B.n174 10.6151
R1203 B.n178 B.n177 10.6151
R1204 B.n181 B.n178 10.6151
R1205 B.n182 B.n181 10.6151
R1206 B.n185 B.n182 10.6151
R1207 B.n186 B.n185 10.6151
R1208 B.n189 B.n186 10.6151
R1209 B.n190 B.n189 10.6151
R1210 B.n193 B.n190 10.6151
R1211 B.n194 B.n193 10.6151
R1212 B.n197 B.n194 10.6151
R1213 B.n198 B.n197 10.6151
R1214 B.n201 B.n198 10.6151
R1215 B.n202 B.n201 10.6151
R1216 B.n205 B.n202 10.6151
R1217 B.n206 B.n205 10.6151
R1218 B.n209 B.n206 10.6151
R1219 B.n210 B.n209 10.6151
R1220 B.n213 B.n210 10.6151
R1221 B.n214 B.n213 10.6151
R1222 B.n217 B.n214 10.6151
R1223 B.n218 B.n217 10.6151
R1224 B.n221 B.n218 10.6151
R1225 B.n222 B.n221 10.6151
R1226 B.n225 B.n222 10.6151
R1227 B.n226 B.n225 10.6151
R1228 B.n229 B.n226 10.6151
R1229 B.n234 B.n231 10.6151
R1230 B.n235 B.n234 10.6151
R1231 B.n238 B.n235 10.6151
R1232 B.n239 B.n238 10.6151
R1233 B.n242 B.n239 10.6151
R1234 B.n243 B.n242 10.6151
R1235 B.n246 B.n243 10.6151
R1236 B.n247 B.n246 10.6151
R1237 B.n250 B.n247 10.6151
R1238 B.n255 B.n252 10.6151
R1239 B.n256 B.n255 10.6151
R1240 B.n259 B.n256 10.6151
R1241 B.n260 B.n259 10.6151
R1242 B.n263 B.n260 10.6151
R1243 B.n264 B.n263 10.6151
R1244 B.n267 B.n264 10.6151
R1245 B.n268 B.n267 10.6151
R1246 B.n271 B.n268 10.6151
R1247 B.n272 B.n271 10.6151
R1248 B.n275 B.n272 10.6151
R1249 B.n276 B.n275 10.6151
R1250 B.n279 B.n276 10.6151
R1251 B.n280 B.n279 10.6151
R1252 B.n283 B.n280 10.6151
R1253 B.n284 B.n283 10.6151
R1254 B.n287 B.n284 10.6151
R1255 B.n288 B.n287 10.6151
R1256 B.n291 B.n288 10.6151
R1257 B.n292 B.n291 10.6151
R1258 B.n295 B.n292 10.6151
R1259 B.n296 B.n295 10.6151
R1260 B.n299 B.n296 10.6151
R1261 B.n300 B.n299 10.6151
R1262 B.n303 B.n300 10.6151
R1263 B.n304 B.n303 10.6151
R1264 B.n307 B.n304 10.6151
R1265 B.n308 B.n307 10.6151
R1266 B.n311 B.n308 10.6151
R1267 B.n312 B.n311 10.6151
R1268 B.n315 B.n312 10.6151
R1269 B.n316 B.n315 10.6151
R1270 B.n319 B.n316 10.6151
R1271 B.n320 B.n319 10.6151
R1272 B.n323 B.n320 10.6151
R1273 B.n324 B.n323 10.6151
R1274 B.n327 B.n324 10.6151
R1275 B.n328 B.n327 10.6151
R1276 B.n331 B.n328 10.6151
R1277 B.n332 B.n331 10.6151
R1278 B.n335 B.n332 10.6151
R1279 B.n336 B.n335 10.6151
R1280 B.n339 B.n336 10.6151
R1281 B.n340 B.n339 10.6151
R1282 B.n343 B.n340 10.6151
R1283 B.n344 B.n343 10.6151
R1284 B.n347 B.n344 10.6151
R1285 B.n348 B.n347 10.6151
R1286 B.n351 B.n348 10.6151
R1287 B.n352 B.n351 10.6151
R1288 B.n355 B.n352 10.6151
R1289 B.n357 B.n355 10.6151
R1290 B.n358 B.n357 10.6151
R1291 B.n844 B.n358 10.6151
R1292 B.n721 B.n720 10.6151
R1293 B.n721 B.n406 10.6151
R1294 B.n731 B.n406 10.6151
R1295 B.n732 B.n731 10.6151
R1296 B.n733 B.n732 10.6151
R1297 B.n733 B.n397 10.6151
R1298 B.n743 B.n397 10.6151
R1299 B.n744 B.n743 10.6151
R1300 B.n745 B.n744 10.6151
R1301 B.n745 B.n390 10.6151
R1302 B.n755 B.n390 10.6151
R1303 B.n756 B.n755 10.6151
R1304 B.n757 B.n756 10.6151
R1305 B.n757 B.n382 10.6151
R1306 B.n767 B.n382 10.6151
R1307 B.n768 B.n767 10.6151
R1308 B.n769 B.n768 10.6151
R1309 B.n769 B.n374 10.6151
R1310 B.n779 B.n374 10.6151
R1311 B.n780 B.n779 10.6151
R1312 B.n781 B.n780 10.6151
R1313 B.n781 B.n367 10.6151
R1314 B.n792 B.n367 10.6151
R1315 B.n793 B.n792 10.6151
R1316 B.n795 B.n793 10.6151
R1317 B.n795 B.n794 10.6151
R1318 B.n794 B.n359 10.6151
R1319 B.n806 B.n359 10.6151
R1320 B.n807 B.n806 10.6151
R1321 B.n808 B.n807 10.6151
R1322 B.n809 B.n808 10.6151
R1323 B.n811 B.n809 10.6151
R1324 B.n812 B.n811 10.6151
R1325 B.n813 B.n812 10.6151
R1326 B.n814 B.n813 10.6151
R1327 B.n816 B.n814 10.6151
R1328 B.n817 B.n816 10.6151
R1329 B.n818 B.n817 10.6151
R1330 B.n819 B.n818 10.6151
R1331 B.n821 B.n819 10.6151
R1332 B.n822 B.n821 10.6151
R1333 B.n823 B.n822 10.6151
R1334 B.n824 B.n823 10.6151
R1335 B.n826 B.n824 10.6151
R1336 B.n827 B.n826 10.6151
R1337 B.n828 B.n827 10.6151
R1338 B.n829 B.n828 10.6151
R1339 B.n831 B.n829 10.6151
R1340 B.n832 B.n831 10.6151
R1341 B.n833 B.n832 10.6151
R1342 B.n834 B.n833 10.6151
R1343 B.n836 B.n834 10.6151
R1344 B.n837 B.n836 10.6151
R1345 B.n838 B.n837 10.6151
R1346 B.n839 B.n838 10.6151
R1347 B.n841 B.n839 10.6151
R1348 B.n842 B.n841 10.6151
R1349 B.n843 B.n842 10.6151
R1350 B.n714 B.n713 10.6151
R1351 B.n713 B.n712 10.6151
R1352 B.n712 B.n711 10.6151
R1353 B.n711 B.n709 10.6151
R1354 B.n709 B.n706 10.6151
R1355 B.n706 B.n705 10.6151
R1356 B.n705 B.n702 10.6151
R1357 B.n702 B.n701 10.6151
R1358 B.n701 B.n698 10.6151
R1359 B.n698 B.n697 10.6151
R1360 B.n697 B.n694 10.6151
R1361 B.n694 B.n693 10.6151
R1362 B.n693 B.n690 10.6151
R1363 B.n690 B.n689 10.6151
R1364 B.n689 B.n686 10.6151
R1365 B.n686 B.n685 10.6151
R1366 B.n685 B.n682 10.6151
R1367 B.n682 B.n681 10.6151
R1368 B.n681 B.n678 10.6151
R1369 B.n678 B.n677 10.6151
R1370 B.n677 B.n674 10.6151
R1371 B.n674 B.n673 10.6151
R1372 B.n673 B.n670 10.6151
R1373 B.n670 B.n669 10.6151
R1374 B.n669 B.n666 10.6151
R1375 B.n666 B.n665 10.6151
R1376 B.n665 B.n662 10.6151
R1377 B.n662 B.n661 10.6151
R1378 B.n661 B.n658 10.6151
R1379 B.n658 B.n657 10.6151
R1380 B.n657 B.n654 10.6151
R1381 B.n654 B.n653 10.6151
R1382 B.n653 B.n650 10.6151
R1383 B.n650 B.n649 10.6151
R1384 B.n649 B.n646 10.6151
R1385 B.n646 B.n645 10.6151
R1386 B.n645 B.n642 10.6151
R1387 B.n642 B.n641 10.6151
R1388 B.n641 B.n638 10.6151
R1389 B.n638 B.n637 10.6151
R1390 B.n637 B.n634 10.6151
R1391 B.n634 B.n633 10.6151
R1392 B.n633 B.n630 10.6151
R1393 B.n630 B.n629 10.6151
R1394 B.n629 B.n626 10.6151
R1395 B.n626 B.n625 10.6151
R1396 B.n625 B.n622 10.6151
R1397 B.n622 B.n621 10.6151
R1398 B.n621 B.n618 10.6151
R1399 B.n618 B.n617 10.6151
R1400 B.n617 B.n614 10.6151
R1401 B.n614 B.n613 10.6151
R1402 B.n613 B.n610 10.6151
R1403 B.n610 B.n609 10.6151
R1404 B.n606 B.n605 10.6151
R1405 B.n605 B.n602 10.6151
R1406 B.n602 B.n601 10.6151
R1407 B.n601 B.n598 10.6151
R1408 B.n598 B.n597 10.6151
R1409 B.n597 B.n594 10.6151
R1410 B.n594 B.n593 10.6151
R1411 B.n593 B.n590 10.6151
R1412 B.n590 B.n589 10.6151
R1413 B.n586 B.n585 10.6151
R1414 B.n585 B.n582 10.6151
R1415 B.n582 B.n581 10.6151
R1416 B.n581 B.n578 10.6151
R1417 B.n578 B.n577 10.6151
R1418 B.n577 B.n574 10.6151
R1419 B.n574 B.n573 10.6151
R1420 B.n573 B.n570 10.6151
R1421 B.n570 B.n569 10.6151
R1422 B.n569 B.n566 10.6151
R1423 B.n566 B.n565 10.6151
R1424 B.n565 B.n562 10.6151
R1425 B.n562 B.n561 10.6151
R1426 B.n561 B.n558 10.6151
R1427 B.n558 B.n557 10.6151
R1428 B.n557 B.n554 10.6151
R1429 B.n554 B.n553 10.6151
R1430 B.n553 B.n550 10.6151
R1431 B.n550 B.n549 10.6151
R1432 B.n549 B.n546 10.6151
R1433 B.n546 B.n545 10.6151
R1434 B.n545 B.n542 10.6151
R1435 B.n542 B.n541 10.6151
R1436 B.n541 B.n538 10.6151
R1437 B.n538 B.n537 10.6151
R1438 B.n537 B.n534 10.6151
R1439 B.n534 B.n533 10.6151
R1440 B.n533 B.n530 10.6151
R1441 B.n530 B.n529 10.6151
R1442 B.n529 B.n526 10.6151
R1443 B.n526 B.n525 10.6151
R1444 B.n525 B.n522 10.6151
R1445 B.n522 B.n521 10.6151
R1446 B.n521 B.n518 10.6151
R1447 B.n518 B.n517 10.6151
R1448 B.n517 B.n514 10.6151
R1449 B.n514 B.n513 10.6151
R1450 B.n513 B.n510 10.6151
R1451 B.n510 B.n509 10.6151
R1452 B.n509 B.n506 10.6151
R1453 B.n506 B.n505 10.6151
R1454 B.n505 B.n502 10.6151
R1455 B.n502 B.n501 10.6151
R1456 B.n501 B.n498 10.6151
R1457 B.n498 B.n497 10.6151
R1458 B.n497 B.n494 10.6151
R1459 B.n494 B.n493 10.6151
R1460 B.n493 B.n490 10.6151
R1461 B.n490 B.n489 10.6151
R1462 B.n489 B.n486 10.6151
R1463 B.n486 B.n485 10.6151
R1464 B.n485 B.n482 10.6151
R1465 B.n482 B.n414 10.6151
R1466 B.n719 B.n414 10.6151
R1467 B.n725 B.n410 10.6151
R1468 B.n726 B.n725 10.6151
R1469 B.n727 B.n726 10.6151
R1470 B.n727 B.n402 10.6151
R1471 B.n737 B.n402 10.6151
R1472 B.n738 B.n737 10.6151
R1473 B.n739 B.n738 10.6151
R1474 B.n739 B.n394 10.6151
R1475 B.n749 B.n394 10.6151
R1476 B.n750 B.n749 10.6151
R1477 B.n751 B.n750 10.6151
R1478 B.n751 B.n386 10.6151
R1479 B.n761 B.n386 10.6151
R1480 B.n762 B.n761 10.6151
R1481 B.n763 B.n762 10.6151
R1482 B.n763 B.n378 10.6151
R1483 B.n773 B.n378 10.6151
R1484 B.n774 B.n773 10.6151
R1485 B.n775 B.n774 10.6151
R1486 B.n775 B.n370 10.6151
R1487 B.n786 B.n370 10.6151
R1488 B.n787 B.n786 10.6151
R1489 B.n788 B.n787 10.6151
R1490 B.n788 B.n363 10.6151
R1491 B.n799 B.n363 10.6151
R1492 B.n800 B.n799 10.6151
R1493 B.n801 B.n800 10.6151
R1494 B.n801 B.n0 10.6151
R1495 B.n901 B.n1 10.6151
R1496 B.n901 B.n900 10.6151
R1497 B.n900 B.n899 10.6151
R1498 B.n899 B.n10 10.6151
R1499 B.n893 B.n10 10.6151
R1500 B.n893 B.n892 10.6151
R1501 B.n892 B.n891 10.6151
R1502 B.n891 B.n16 10.6151
R1503 B.n885 B.n16 10.6151
R1504 B.n885 B.n884 10.6151
R1505 B.n884 B.n883 10.6151
R1506 B.n883 B.n24 10.6151
R1507 B.n877 B.n24 10.6151
R1508 B.n877 B.n876 10.6151
R1509 B.n876 B.n875 10.6151
R1510 B.n875 B.n31 10.6151
R1511 B.n869 B.n31 10.6151
R1512 B.n869 B.n868 10.6151
R1513 B.n868 B.n867 10.6151
R1514 B.n867 B.n38 10.6151
R1515 B.n861 B.n38 10.6151
R1516 B.n861 B.n860 10.6151
R1517 B.n860 B.n859 10.6151
R1518 B.n859 B.n45 10.6151
R1519 B.n853 B.n45 10.6151
R1520 B.n853 B.n852 10.6151
R1521 B.n852 B.n851 10.6151
R1522 B.n851 B.n52 10.6151
R1523 B.n230 B.n229 9.36635
R1524 B.n252 B.n251 9.36635
R1525 B.n609 B.n478 9.36635
R1526 B.n586 B.n481 9.36635
R1527 B.n783 B.t1 5.03367
R1528 B.n18 B.t0 5.03367
R1529 B.n907 B.n0 2.81026
R1530 B.n907 B.n1 2.81026
R1531 B.n231 B.n230 1.24928
R1532 B.n251 B.n250 1.24928
R1533 B.n606 B.n478 1.24928
R1534 B.n589 B.n481 1.24928
R1535 VN VN.t1 211.904
R1536 VN VN.t0 162.698
R1537 VDD2.n0 VDD2.t1 108.766
R1538 VDD2.n0 VDD2.t0 64.6588
R1539 VDD2 VDD2.n0 0.828086
C0 VTAIL VP 3.3761f
C1 VDD1 VP 4.07313f
C2 VP VN 6.60369f
C3 VDD2 VP 0.36059f
C4 VDD1 VTAIL 6.34855f
C5 VTAIL VN 3.3618f
C6 VDD2 VTAIL 6.40319f
C7 VDD1 VN 0.14875f
C8 VDD2 VDD1 0.752984f
C9 VDD2 VN 3.86421f
C10 VDD2 B 5.473763f
C11 VDD1 B 9.062779f
C12 VTAIL B 9.546313f
C13 VN B 12.437881f
C14 VP B 7.511174f
C15 VDD2.t1 B 3.75232f
C16 VDD2.t0 B 3.0623f
C17 VDD2.n0 B 3.3314f
C18 VN.t0 B 4.18613f
C19 VN.t1 B 4.82571f
C20 VDD1.t1 B 3.0734f
C21 VDD1.t0 B 3.80479f
C22 VTAIL.t2 B 2.98481f
C23 VTAIL.n0 B 1.94378f
C24 VTAIL.t1 B 2.98482f
C25 VTAIL.n1 B 1.98983f
C26 VTAIL.t3 B 2.98481f
C27 VTAIL.n2 B 1.79054f
C28 VTAIL.t0 B 2.98481f
C29 VTAIL.n3 B 1.70652f
C30 VP.t0 B 4.90824f
C31 VP.t1 B 4.25316f
C32 VP.n0 B 4.84839f
.ends

