* NGSPICE file created from diff_pair_sample_1687.ext - technology: sky130A

.subckt diff_pair_sample_1687 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t3 VN.t0 VDD2.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=3.9273 pd=20.92 as=1.66155 ps=10.4 w=10.07 l=3.76
X1 B.t17 B.t15 B.t16 B.t12 sky130_fd_pr__nfet_01v8 ad=3.9273 pd=20.92 as=0 ps=0 w=10.07 l=3.76
X2 VDD1.t3 VP.t0 VTAIL.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=1.66155 pd=10.4 as=3.9273 ps=20.92 w=10.07 l=3.76
X3 VTAIL.t2 VN.t1 VDD2.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=3.9273 pd=20.92 as=1.66155 ps=10.4 w=10.07 l=3.76
X4 VDD1.t2 VP.t1 VTAIL.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=1.66155 pd=10.4 as=3.9273 ps=20.92 w=10.07 l=3.76
X5 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=3.9273 pd=20.92 as=0 ps=0 w=10.07 l=3.76
X6 VTAIL.t4 VP.t2 VDD1.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=3.9273 pd=20.92 as=1.66155 ps=10.4 w=10.07 l=3.76
X7 VTAIL.t5 VP.t3 VDD1.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=3.9273 pd=20.92 as=1.66155 ps=10.4 w=10.07 l=3.76
X8 VDD2.t3 VN.t2 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.66155 pd=10.4 as=3.9273 ps=20.92 w=10.07 l=3.76
X9 B.t10 B.t8 B.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=3.9273 pd=20.92 as=0 ps=0 w=10.07 l=3.76
X10 VDD2.t2 VN.t3 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.66155 pd=10.4 as=3.9273 ps=20.92 w=10.07 l=3.76
X11 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=3.9273 pd=20.92 as=0 ps=0 w=10.07 l=3.76
R0 VN.n0 VN.t0 98.2304
R1 VN.n1 VN.t2 98.2304
R2 VN.n0 VN.t3 96.8902
R3 VN.n1 VN.t1 96.8902
R4 VN VN.n1 50.4833
R5 VN VN.n0 1.88864
R6 VDD2.n2 VDD2.n0 107.746
R7 VDD2.n2 VDD2.n1 64.7735
R8 VDD2.n1 VDD2.t1 1.96674
R9 VDD2.n1 VDD2.t3 1.96674
R10 VDD2.n0 VDD2.t0 1.96674
R11 VDD2.n0 VDD2.t2 1.96674
R12 VDD2 VDD2.n2 0.0586897
R13 VTAIL.n426 VTAIL.n378 289.615
R14 VTAIL.n48 VTAIL.n0 289.615
R15 VTAIL.n102 VTAIL.n54 289.615
R16 VTAIL.n156 VTAIL.n108 289.615
R17 VTAIL.n372 VTAIL.n324 289.615
R18 VTAIL.n318 VTAIL.n270 289.615
R19 VTAIL.n264 VTAIL.n216 289.615
R20 VTAIL.n210 VTAIL.n162 289.615
R21 VTAIL.n394 VTAIL.n393 185
R22 VTAIL.n399 VTAIL.n398 185
R23 VTAIL.n401 VTAIL.n400 185
R24 VTAIL.n390 VTAIL.n389 185
R25 VTAIL.n407 VTAIL.n406 185
R26 VTAIL.n409 VTAIL.n408 185
R27 VTAIL.n386 VTAIL.n385 185
R28 VTAIL.n416 VTAIL.n415 185
R29 VTAIL.n417 VTAIL.n384 185
R30 VTAIL.n419 VTAIL.n418 185
R31 VTAIL.n382 VTAIL.n381 185
R32 VTAIL.n425 VTAIL.n424 185
R33 VTAIL.n427 VTAIL.n426 185
R34 VTAIL.n16 VTAIL.n15 185
R35 VTAIL.n21 VTAIL.n20 185
R36 VTAIL.n23 VTAIL.n22 185
R37 VTAIL.n12 VTAIL.n11 185
R38 VTAIL.n29 VTAIL.n28 185
R39 VTAIL.n31 VTAIL.n30 185
R40 VTAIL.n8 VTAIL.n7 185
R41 VTAIL.n38 VTAIL.n37 185
R42 VTAIL.n39 VTAIL.n6 185
R43 VTAIL.n41 VTAIL.n40 185
R44 VTAIL.n4 VTAIL.n3 185
R45 VTAIL.n47 VTAIL.n46 185
R46 VTAIL.n49 VTAIL.n48 185
R47 VTAIL.n70 VTAIL.n69 185
R48 VTAIL.n75 VTAIL.n74 185
R49 VTAIL.n77 VTAIL.n76 185
R50 VTAIL.n66 VTAIL.n65 185
R51 VTAIL.n83 VTAIL.n82 185
R52 VTAIL.n85 VTAIL.n84 185
R53 VTAIL.n62 VTAIL.n61 185
R54 VTAIL.n92 VTAIL.n91 185
R55 VTAIL.n93 VTAIL.n60 185
R56 VTAIL.n95 VTAIL.n94 185
R57 VTAIL.n58 VTAIL.n57 185
R58 VTAIL.n101 VTAIL.n100 185
R59 VTAIL.n103 VTAIL.n102 185
R60 VTAIL.n124 VTAIL.n123 185
R61 VTAIL.n129 VTAIL.n128 185
R62 VTAIL.n131 VTAIL.n130 185
R63 VTAIL.n120 VTAIL.n119 185
R64 VTAIL.n137 VTAIL.n136 185
R65 VTAIL.n139 VTAIL.n138 185
R66 VTAIL.n116 VTAIL.n115 185
R67 VTAIL.n146 VTAIL.n145 185
R68 VTAIL.n147 VTAIL.n114 185
R69 VTAIL.n149 VTAIL.n148 185
R70 VTAIL.n112 VTAIL.n111 185
R71 VTAIL.n155 VTAIL.n154 185
R72 VTAIL.n157 VTAIL.n156 185
R73 VTAIL.n373 VTAIL.n372 185
R74 VTAIL.n371 VTAIL.n370 185
R75 VTAIL.n328 VTAIL.n327 185
R76 VTAIL.n365 VTAIL.n364 185
R77 VTAIL.n363 VTAIL.n330 185
R78 VTAIL.n362 VTAIL.n361 185
R79 VTAIL.n333 VTAIL.n331 185
R80 VTAIL.n356 VTAIL.n355 185
R81 VTAIL.n354 VTAIL.n353 185
R82 VTAIL.n337 VTAIL.n336 185
R83 VTAIL.n348 VTAIL.n347 185
R84 VTAIL.n346 VTAIL.n345 185
R85 VTAIL.n341 VTAIL.n340 185
R86 VTAIL.n319 VTAIL.n318 185
R87 VTAIL.n317 VTAIL.n316 185
R88 VTAIL.n274 VTAIL.n273 185
R89 VTAIL.n311 VTAIL.n310 185
R90 VTAIL.n309 VTAIL.n276 185
R91 VTAIL.n308 VTAIL.n307 185
R92 VTAIL.n279 VTAIL.n277 185
R93 VTAIL.n302 VTAIL.n301 185
R94 VTAIL.n300 VTAIL.n299 185
R95 VTAIL.n283 VTAIL.n282 185
R96 VTAIL.n294 VTAIL.n293 185
R97 VTAIL.n292 VTAIL.n291 185
R98 VTAIL.n287 VTAIL.n286 185
R99 VTAIL.n265 VTAIL.n264 185
R100 VTAIL.n263 VTAIL.n262 185
R101 VTAIL.n220 VTAIL.n219 185
R102 VTAIL.n257 VTAIL.n256 185
R103 VTAIL.n255 VTAIL.n222 185
R104 VTAIL.n254 VTAIL.n253 185
R105 VTAIL.n225 VTAIL.n223 185
R106 VTAIL.n248 VTAIL.n247 185
R107 VTAIL.n246 VTAIL.n245 185
R108 VTAIL.n229 VTAIL.n228 185
R109 VTAIL.n240 VTAIL.n239 185
R110 VTAIL.n238 VTAIL.n237 185
R111 VTAIL.n233 VTAIL.n232 185
R112 VTAIL.n211 VTAIL.n210 185
R113 VTAIL.n209 VTAIL.n208 185
R114 VTAIL.n166 VTAIL.n165 185
R115 VTAIL.n203 VTAIL.n202 185
R116 VTAIL.n201 VTAIL.n168 185
R117 VTAIL.n200 VTAIL.n199 185
R118 VTAIL.n171 VTAIL.n169 185
R119 VTAIL.n194 VTAIL.n193 185
R120 VTAIL.n192 VTAIL.n191 185
R121 VTAIL.n175 VTAIL.n174 185
R122 VTAIL.n186 VTAIL.n185 185
R123 VTAIL.n184 VTAIL.n183 185
R124 VTAIL.n179 VTAIL.n178 185
R125 VTAIL.n395 VTAIL.t0 149.524
R126 VTAIL.n17 VTAIL.t3 149.524
R127 VTAIL.n71 VTAIL.t7 149.524
R128 VTAIL.n125 VTAIL.t5 149.524
R129 VTAIL.n342 VTAIL.t6 149.524
R130 VTAIL.n288 VTAIL.t4 149.524
R131 VTAIL.n234 VTAIL.t1 149.524
R132 VTAIL.n180 VTAIL.t2 149.524
R133 VTAIL.n399 VTAIL.n393 104.615
R134 VTAIL.n400 VTAIL.n399 104.615
R135 VTAIL.n400 VTAIL.n389 104.615
R136 VTAIL.n407 VTAIL.n389 104.615
R137 VTAIL.n408 VTAIL.n407 104.615
R138 VTAIL.n408 VTAIL.n385 104.615
R139 VTAIL.n416 VTAIL.n385 104.615
R140 VTAIL.n417 VTAIL.n416 104.615
R141 VTAIL.n418 VTAIL.n417 104.615
R142 VTAIL.n418 VTAIL.n381 104.615
R143 VTAIL.n425 VTAIL.n381 104.615
R144 VTAIL.n426 VTAIL.n425 104.615
R145 VTAIL.n21 VTAIL.n15 104.615
R146 VTAIL.n22 VTAIL.n21 104.615
R147 VTAIL.n22 VTAIL.n11 104.615
R148 VTAIL.n29 VTAIL.n11 104.615
R149 VTAIL.n30 VTAIL.n29 104.615
R150 VTAIL.n30 VTAIL.n7 104.615
R151 VTAIL.n38 VTAIL.n7 104.615
R152 VTAIL.n39 VTAIL.n38 104.615
R153 VTAIL.n40 VTAIL.n39 104.615
R154 VTAIL.n40 VTAIL.n3 104.615
R155 VTAIL.n47 VTAIL.n3 104.615
R156 VTAIL.n48 VTAIL.n47 104.615
R157 VTAIL.n75 VTAIL.n69 104.615
R158 VTAIL.n76 VTAIL.n75 104.615
R159 VTAIL.n76 VTAIL.n65 104.615
R160 VTAIL.n83 VTAIL.n65 104.615
R161 VTAIL.n84 VTAIL.n83 104.615
R162 VTAIL.n84 VTAIL.n61 104.615
R163 VTAIL.n92 VTAIL.n61 104.615
R164 VTAIL.n93 VTAIL.n92 104.615
R165 VTAIL.n94 VTAIL.n93 104.615
R166 VTAIL.n94 VTAIL.n57 104.615
R167 VTAIL.n101 VTAIL.n57 104.615
R168 VTAIL.n102 VTAIL.n101 104.615
R169 VTAIL.n129 VTAIL.n123 104.615
R170 VTAIL.n130 VTAIL.n129 104.615
R171 VTAIL.n130 VTAIL.n119 104.615
R172 VTAIL.n137 VTAIL.n119 104.615
R173 VTAIL.n138 VTAIL.n137 104.615
R174 VTAIL.n138 VTAIL.n115 104.615
R175 VTAIL.n146 VTAIL.n115 104.615
R176 VTAIL.n147 VTAIL.n146 104.615
R177 VTAIL.n148 VTAIL.n147 104.615
R178 VTAIL.n148 VTAIL.n111 104.615
R179 VTAIL.n155 VTAIL.n111 104.615
R180 VTAIL.n156 VTAIL.n155 104.615
R181 VTAIL.n372 VTAIL.n371 104.615
R182 VTAIL.n371 VTAIL.n327 104.615
R183 VTAIL.n364 VTAIL.n327 104.615
R184 VTAIL.n364 VTAIL.n363 104.615
R185 VTAIL.n363 VTAIL.n362 104.615
R186 VTAIL.n362 VTAIL.n331 104.615
R187 VTAIL.n355 VTAIL.n331 104.615
R188 VTAIL.n355 VTAIL.n354 104.615
R189 VTAIL.n354 VTAIL.n336 104.615
R190 VTAIL.n347 VTAIL.n336 104.615
R191 VTAIL.n347 VTAIL.n346 104.615
R192 VTAIL.n346 VTAIL.n340 104.615
R193 VTAIL.n318 VTAIL.n317 104.615
R194 VTAIL.n317 VTAIL.n273 104.615
R195 VTAIL.n310 VTAIL.n273 104.615
R196 VTAIL.n310 VTAIL.n309 104.615
R197 VTAIL.n309 VTAIL.n308 104.615
R198 VTAIL.n308 VTAIL.n277 104.615
R199 VTAIL.n301 VTAIL.n277 104.615
R200 VTAIL.n301 VTAIL.n300 104.615
R201 VTAIL.n300 VTAIL.n282 104.615
R202 VTAIL.n293 VTAIL.n282 104.615
R203 VTAIL.n293 VTAIL.n292 104.615
R204 VTAIL.n292 VTAIL.n286 104.615
R205 VTAIL.n264 VTAIL.n263 104.615
R206 VTAIL.n263 VTAIL.n219 104.615
R207 VTAIL.n256 VTAIL.n219 104.615
R208 VTAIL.n256 VTAIL.n255 104.615
R209 VTAIL.n255 VTAIL.n254 104.615
R210 VTAIL.n254 VTAIL.n223 104.615
R211 VTAIL.n247 VTAIL.n223 104.615
R212 VTAIL.n247 VTAIL.n246 104.615
R213 VTAIL.n246 VTAIL.n228 104.615
R214 VTAIL.n239 VTAIL.n228 104.615
R215 VTAIL.n239 VTAIL.n238 104.615
R216 VTAIL.n238 VTAIL.n232 104.615
R217 VTAIL.n210 VTAIL.n209 104.615
R218 VTAIL.n209 VTAIL.n165 104.615
R219 VTAIL.n202 VTAIL.n165 104.615
R220 VTAIL.n202 VTAIL.n201 104.615
R221 VTAIL.n201 VTAIL.n200 104.615
R222 VTAIL.n200 VTAIL.n169 104.615
R223 VTAIL.n193 VTAIL.n169 104.615
R224 VTAIL.n193 VTAIL.n192 104.615
R225 VTAIL.n192 VTAIL.n174 104.615
R226 VTAIL.n185 VTAIL.n174 104.615
R227 VTAIL.n185 VTAIL.n184 104.615
R228 VTAIL.n184 VTAIL.n178 104.615
R229 VTAIL.t0 VTAIL.n393 52.3082
R230 VTAIL.t3 VTAIL.n15 52.3082
R231 VTAIL.t7 VTAIL.n69 52.3082
R232 VTAIL.t5 VTAIL.n123 52.3082
R233 VTAIL.t6 VTAIL.n340 52.3082
R234 VTAIL.t4 VTAIL.n286 52.3082
R235 VTAIL.t1 VTAIL.n232 52.3082
R236 VTAIL.t2 VTAIL.n178 52.3082
R237 VTAIL.n431 VTAIL.n430 34.3187
R238 VTAIL.n53 VTAIL.n52 34.3187
R239 VTAIL.n107 VTAIL.n106 34.3187
R240 VTAIL.n161 VTAIL.n160 34.3187
R241 VTAIL.n377 VTAIL.n376 34.3187
R242 VTAIL.n323 VTAIL.n322 34.3187
R243 VTAIL.n269 VTAIL.n268 34.3187
R244 VTAIL.n215 VTAIL.n214 34.3187
R245 VTAIL.n431 VTAIL.n377 24.5738
R246 VTAIL.n215 VTAIL.n161 24.5738
R247 VTAIL.n419 VTAIL.n384 13.1884
R248 VTAIL.n41 VTAIL.n6 13.1884
R249 VTAIL.n95 VTAIL.n60 13.1884
R250 VTAIL.n149 VTAIL.n114 13.1884
R251 VTAIL.n365 VTAIL.n330 13.1884
R252 VTAIL.n311 VTAIL.n276 13.1884
R253 VTAIL.n257 VTAIL.n222 13.1884
R254 VTAIL.n203 VTAIL.n168 13.1884
R255 VTAIL.n415 VTAIL.n414 12.8005
R256 VTAIL.n420 VTAIL.n382 12.8005
R257 VTAIL.n37 VTAIL.n36 12.8005
R258 VTAIL.n42 VTAIL.n4 12.8005
R259 VTAIL.n91 VTAIL.n90 12.8005
R260 VTAIL.n96 VTAIL.n58 12.8005
R261 VTAIL.n145 VTAIL.n144 12.8005
R262 VTAIL.n150 VTAIL.n112 12.8005
R263 VTAIL.n366 VTAIL.n328 12.8005
R264 VTAIL.n361 VTAIL.n332 12.8005
R265 VTAIL.n312 VTAIL.n274 12.8005
R266 VTAIL.n307 VTAIL.n278 12.8005
R267 VTAIL.n258 VTAIL.n220 12.8005
R268 VTAIL.n253 VTAIL.n224 12.8005
R269 VTAIL.n204 VTAIL.n166 12.8005
R270 VTAIL.n199 VTAIL.n170 12.8005
R271 VTAIL.n413 VTAIL.n386 12.0247
R272 VTAIL.n424 VTAIL.n423 12.0247
R273 VTAIL.n35 VTAIL.n8 12.0247
R274 VTAIL.n46 VTAIL.n45 12.0247
R275 VTAIL.n89 VTAIL.n62 12.0247
R276 VTAIL.n100 VTAIL.n99 12.0247
R277 VTAIL.n143 VTAIL.n116 12.0247
R278 VTAIL.n154 VTAIL.n153 12.0247
R279 VTAIL.n370 VTAIL.n369 12.0247
R280 VTAIL.n360 VTAIL.n333 12.0247
R281 VTAIL.n316 VTAIL.n315 12.0247
R282 VTAIL.n306 VTAIL.n279 12.0247
R283 VTAIL.n262 VTAIL.n261 12.0247
R284 VTAIL.n252 VTAIL.n225 12.0247
R285 VTAIL.n208 VTAIL.n207 12.0247
R286 VTAIL.n198 VTAIL.n171 12.0247
R287 VTAIL.n410 VTAIL.n409 11.249
R288 VTAIL.n427 VTAIL.n380 11.249
R289 VTAIL.n32 VTAIL.n31 11.249
R290 VTAIL.n49 VTAIL.n2 11.249
R291 VTAIL.n86 VTAIL.n85 11.249
R292 VTAIL.n103 VTAIL.n56 11.249
R293 VTAIL.n140 VTAIL.n139 11.249
R294 VTAIL.n157 VTAIL.n110 11.249
R295 VTAIL.n373 VTAIL.n326 11.249
R296 VTAIL.n357 VTAIL.n356 11.249
R297 VTAIL.n319 VTAIL.n272 11.249
R298 VTAIL.n303 VTAIL.n302 11.249
R299 VTAIL.n265 VTAIL.n218 11.249
R300 VTAIL.n249 VTAIL.n248 11.249
R301 VTAIL.n211 VTAIL.n164 11.249
R302 VTAIL.n195 VTAIL.n194 11.249
R303 VTAIL.n406 VTAIL.n388 10.4732
R304 VTAIL.n428 VTAIL.n378 10.4732
R305 VTAIL.n28 VTAIL.n10 10.4732
R306 VTAIL.n50 VTAIL.n0 10.4732
R307 VTAIL.n82 VTAIL.n64 10.4732
R308 VTAIL.n104 VTAIL.n54 10.4732
R309 VTAIL.n136 VTAIL.n118 10.4732
R310 VTAIL.n158 VTAIL.n108 10.4732
R311 VTAIL.n374 VTAIL.n324 10.4732
R312 VTAIL.n353 VTAIL.n335 10.4732
R313 VTAIL.n320 VTAIL.n270 10.4732
R314 VTAIL.n299 VTAIL.n281 10.4732
R315 VTAIL.n266 VTAIL.n216 10.4732
R316 VTAIL.n245 VTAIL.n227 10.4732
R317 VTAIL.n212 VTAIL.n162 10.4732
R318 VTAIL.n191 VTAIL.n173 10.4732
R319 VTAIL.n395 VTAIL.n394 10.2747
R320 VTAIL.n17 VTAIL.n16 10.2747
R321 VTAIL.n71 VTAIL.n70 10.2747
R322 VTAIL.n125 VTAIL.n124 10.2747
R323 VTAIL.n342 VTAIL.n341 10.2747
R324 VTAIL.n288 VTAIL.n287 10.2747
R325 VTAIL.n234 VTAIL.n233 10.2747
R326 VTAIL.n180 VTAIL.n179 10.2747
R327 VTAIL.n405 VTAIL.n390 9.69747
R328 VTAIL.n27 VTAIL.n12 9.69747
R329 VTAIL.n81 VTAIL.n66 9.69747
R330 VTAIL.n135 VTAIL.n120 9.69747
R331 VTAIL.n352 VTAIL.n337 9.69747
R332 VTAIL.n298 VTAIL.n283 9.69747
R333 VTAIL.n244 VTAIL.n229 9.69747
R334 VTAIL.n190 VTAIL.n175 9.69747
R335 VTAIL.n430 VTAIL.n429 9.45567
R336 VTAIL.n52 VTAIL.n51 9.45567
R337 VTAIL.n106 VTAIL.n105 9.45567
R338 VTAIL.n160 VTAIL.n159 9.45567
R339 VTAIL.n376 VTAIL.n375 9.45567
R340 VTAIL.n322 VTAIL.n321 9.45567
R341 VTAIL.n268 VTAIL.n267 9.45567
R342 VTAIL.n214 VTAIL.n213 9.45567
R343 VTAIL.n429 VTAIL.n428 9.3005
R344 VTAIL.n380 VTAIL.n379 9.3005
R345 VTAIL.n423 VTAIL.n422 9.3005
R346 VTAIL.n421 VTAIL.n420 9.3005
R347 VTAIL.n397 VTAIL.n396 9.3005
R348 VTAIL.n392 VTAIL.n391 9.3005
R349 VTAIL.n403 VTAIL.n402 9.3005
R350 VTAIL.n405 VTAIL.n404 9.3005
R351 VTAIL.n388 VTAIL.n387 9.3005
R352 VTAIL.n411 VTAIL.n410 9.3005
R353 VTAIL.n413 VTAIL.n412 9.3005
R354 VTAIL.n414 VTAIL.n383 9.3005
R355 VTAIL.n51 VTAIL.n50 9.3005
R356 VTAIL.n2 VTAIL.n1 9.3005
R357 VTAIL.n45 VTAIL.n44 9.3005
R358 VTAIL.n43 VTAIL.n42 9.3005
R359 VTAIL.n19 VTAIL.n18 9.3005
R360 VTAIL.n14 VTAIL.n13 9.3005
R361 VTAIL.n25 VTAIL.n24 9.3005
R362 VTAIL.n27 VTAIL.n26 9.3005
R363 VTAIL.n10 VTAIL.n9 9.3005
R364 VTAIL.n33 VTAIL.n32 9.3005
R365 VTAIL.n35 VTAIL.n34 9.3005
R366 VTAIL.n36 VTAIL.n5 9.3005
R367 VTAIL.n105 VTAIL.n104 9.3005
R368 VTAIL.n56 VTAIL.n55 9.3005
R369 VTAIL.n99 VTAIL.n98 9.3005
R370 VTAIL.n97 VTAIL.n96 9.3005
R371 VTAIL.n73 VTAIL.n72 9.3005
R372 VTAIL.n68 VTAIL.n67 9.3005
R373 VTAIL.n79 VTAIL.n78 9.3005
R374 VTAIL.n81 VTAIL.n80 9.3005
R375 VTAIL.n64 VTAIL.n63 9.3005
R376 VTAIL.n87 VTAIL.n86 9.3005
R377 VTAIL.n89 VTAIL.n88 9.3005
R378 VTAIL.n90 VTAIL.n59 9.3005
R379 VTAIL.n159 VTAIL.n158 9.3005
R380 VTAIL.n110 VTAIL.n109 9.3005
R381 VTAIL.n153 VTAIL.n152 9.3005
R382 VTAIL.n151 VTAIL.n150 9.3005
R383 VTAIL.n127 VTAIL.n126 9.3005
R384 VTAIL.n122 VTAIL.n121 9.3005
R385 VTAIL.n133 VTAIL.n132 9.3005
R386 VTAIL.n135 VTAIL.n134 9.3005
R387 VTAIL.n118 VTAIL.n117 9.3005
R388 VTAIL.n141 VTAIL.n140 9.3005
R389 VTAIL.n143 VTAIL.n142 9.3005
R390 VTAIL.n144 VTAIL.n113 9.3005
R391 VTAIL.n344 VTAIL.n343 9.3005
R392 VTAIL.n339 VTAIL.n338 9.3005
R393 VTAIL.n350 VTAIL.n349 9.3005
R394 VTAIL.n352 VTAIL.n351 9.3005
R395 VTAIL.n335 VTAIL.n334 9.3005
R396 VTAIL.n358 VTAIL.n357 9.3005
R397 VTAIL.n360 VTAIL.n359 9.3005
R398 VTAIL.n332 VTAIL.n329 9.3005
R399 VTAIL.n375 VTAIL.n374 9.3005
R400 VTAIL.n326 VTAIL.n325 9.3005
R401 VTAIL.n369 VTAIL.n368 9.3005
R402 VTAIL.n367 VTAIL.n366 9.3005
R403 VTAIL.n290 VTAIL.n289 9.3005
R404 VTAIL.n285 VTAIL.n284 9.3005
R405 VTAIL.n296 VTAIL.n295 9.3005
R406 VTAIL.n298 VTAIL.n297 9.3005
R407 VTAIL.n281 VTAIL.n280 9.3005
R408 VTAIL.n304 VTAIL.n303 9.3005
R409 VTAIL.n306 VTAIL.n305 9.3005
R410 VTAIL.n278 VTAIL.n275 9.3005
R411 VTAIL.n321 VTAIL.n320 9.3005
R412 VTAIL.n272 VTAIL.n271 9.3005
R413 VTAIL.n315 VTAIL.n314 9.3005
R414 VTAIL.n313 VTAIL.n312 9.3005
R415 VTAIL.n236 VTAIL.n235 9.3005
R416 VTAIL.n231 VTAIL.n230 9.3005
R417 VTAIL.n242 VTAIL.n241 9.3005
R418 VTAIL.n244 VTAIL.n243 9.3005
R419 VTAIL.n227 VTAIL.n226 9.3005
R420 VTAIL.n250 VTAIL.n249 9.3005
R421 VTAIL.n252 VTAIL.n251 9.3005
R422 VTAIL.n224 VTAIL.n221 9.3005
R423 VTAIL.n267 VTAIL.n266 9.3005
R424 VTAIL.n218 VTAIL.n217 9.3005
R425 VTAIL.n261 VTAIL.n260 9.3005
R426 VTAIL.n259 VTAIL.n258 9.3005
R427 VTAIL.n182 VTAIL.n181 9.3005
R428 VTAIL.n177 VTAIL.n176 9.3005
R429 VTAIL.n188 VTAIL.n187 9.3005
R430 VTAIL.n190 VTAIL.n189 9.3005
R431 VTAIL.n173 VTAIL.n172 9.3005
R432 VTAIL.n196 VTAIL.n195 9.3005
R433 VTAIL.n198 VTAIL.n197 9.3005
R434 VTAIL.n170 VTAIL.n167 9.3005
R435 VTAIL.n213 VTAIL.n212 9.3005
R436 VTAIL.n164 VTAIL.n163 9.3005
R437 VTAIL.n207 VTAIL.n206 9.3005
R438 VTAIL.n205 VTAIL.n204 9.3005
R439 VTAIL.n402 VTAIL.n401 8.92171
R440 VTAIL.n24 VTAIL.n23 8.92171
R441 VTAIL.n78 VTAIL.n77 8.92171
R442 VTAIL.n132 VTAIL.n131 8.92171
R443 VTAIL.n349 VTAIL.n348 8.92171
R444 VTAIL.n295 VTAIL.n294 8.92171
R445 VTAIL.n241 VTAIL.n240 8.92171
R446 VTAIL.n187 VTAIL.n186 8.92171
R447 VTAIL.n398 VTAIL.n392 8.14595
R448 VTAIL.n20 VTAIL.n14 8.14595
R449 VTAIL.n74 VTAIL.n68 8.14595
R450 VTAIL.n128 VTAIL.n122 8.14595
R451 VTAIL.n345 VTAIL.n339 8.14595
R452 VTAIL.n291 VTAIL.n285 8.14595
R453 VTAIL.n237 VTAIL.n231 8.14595
R454 VTAIL.n183 VTAIL.n177 8.14595
R455 VTAIL.n397 VTAIL.n394 7.3702
R456 VTAIL.n19 VTAIL.n16 7.3702
R457 VTAIL.n73 VTAIL.n70 7.3702
R458 VTAIL.n127 VTAIL.n124 7.3702
R459 VTAIL.n344 VTAIL.n341 7.3702
R460 VTAIL.n290 VTAIL.n287 7.3702
R461 VTAIL.n236 VTAIL.n233 7.3702
R462 VTAIL.n182 VTAIL.n179 7.3702
R463 VTAIL.n398 VTAIL.n397 5.81868
R464 VTAIL.n20 VTAIL.n19 5.81868
R465 VTAIL.n74 VTAIL.n73 5.81868
R466 VTAIL.n128 VTAIL.n127 5.81868
R467 VTAIL.n345 VTAIL.n344 5.81868
R468 VTAIL.n291 VTAIL.n290 5.81868
R469 VTAIL.n237 VTAIL.n236 5.81868
R470 VTAIL.n183 VTAIL.n182 5.81868
R471 VTAIL.n401 VTAIL.n392 5.04292
R472 VTAIL.n23 VTAIL.n14 5.04292
R473 VTAIL.n77 VTAIL.n68 5.04292
R474 VTAIL.n131 VTAIL.n122 5.04292
R475 VTAIL.n348 VTAIL.n339 5.04292
R476 VTAIL.n294 VTAIL.n285 5.04292
R477 VTAIL.n240 VTAIL.n231 5.04292
R478 VTAIL.n186 VTAIL.n177 5.04292
R479 VTAIL.n402 VTAIL.n390 4.26717
R480 VTAIL.n24 VTAIL.n12 4.26717
R481 VTAIL.n78 VTAIL.n66 4.26717
R482 VTAIL.n132 VTAIL.n120 4.26717
R483 VTAIL.n349 VTAIL.n337 4.26717
R484 VTAIL.n295 VTAIL.n283 4.26717
R485 VTAIL.n241 VTAIL.n229 4.26717
R486 VTAIL.n187 VTAIL.n175 4.26717
R487 VTAIL.n269 VTAIL.n215 3.52636
R488 VTAIL.n377 VTAIL.n323 3.52636
R489 VTAIL.n161 VTAIL.n107 3.52636
R490 VTAIL.n406 VTAIL.n405 3.49141
R491 VTAIL.n430 VTAIL.n378 3.49141
R492 VTAIL.n28 VTAIL.n27 3.49141
R493 VTAIL.n52 VTAIL.n0 3.49141
R494 VTAIL.n82 VTAIL.n81 3.49141
R495 VTAIL.n106 VTAIL.n54 3.49141
R496 VTAIL.n136 VTAIL.n135 3.49141
R497 VTAIL.n160 VTAIL.n108 3.49141
R498 VTAIL.n376 VTAIL.n324 3.49141
R499 VTAIL.n353 VTAIL.n352 3.49141
R500 VTAIL.n322 VTAIL.n270 3.49141
R501 VTAIL.n299 VTAIL.n298 3.49141
R502 VTAIL.n268 VTAIL.n216 3.49141
R503 VTAIL.n245 VTAIL.n244 3.49141
R504 VTAIL.n214 VTAIL.n162 3.49141
R505 VTAIL.n191 VTAIL.n190 3.49141
R506 VTAIL.n396 VTAIL.n395 2.84303
R507 VTAIL.n18 VTAIL.n17 2.84303
R508 VTAIL.n72 VTAIL.n71 2.84303
R509 VTAIL.n126 VTAIL.n125 2.84303
R510 VTAIL.n343 VTAIL.n342 2.84303
R511 VTAIL.n289 VTAIL.n288 2.84303
R512 VTAIL.n235 VTAIL.n234 2.84303
R513 VTAIL.n181 VTAIL.n180 2.84303
R514 VTAIL.n409 VTAIL.n388 2.71565
R515 VTAIL.n428 VTAIL.n427 2.71565
R516 VTAIL.n31 VTAIL.n10 2.71565
R517 VTAIL.n50 VTAIL.n49 2.71565
R518 VTAIL.n85 VTAIL.n64 2.71565
R519 VTAIL.n104 VTAIL.n103 2.71565
R520 VTAIL.n139 VTAIL.n118 2.71565
R521 VTAIL.n158 VTAIL.n157 2.71565
R522 VTAIL.n374 VTAIL.n373 2.71565
R523 VTAIL.n356 VTAIL.n335 2.71565
R524 VTAIL.n320 VTAIL.n319 2.71565
R525 VTAIL.n302 VTAIL.n281 2.71565
R526 VTAIL.n266 VTAIL.n265 2.71565
R527 VTAIL.n248 VTAIL.n227 2.71565
R528 VTAIL.n212 VTAIL.n211 2.71565
R529 VTAIL.n194 VTAIL.n173 2.71565
R530 VTAIL.n410 VTAIL.n386 1.93989
R531 VTAIL.n424 VTAIL.n380 1.93989
R532 VTAIL.n32 VTAIL.n8 1.93989
R533 VTAIL.n46 VTAIL.n2 1.93989
R534 VTAIL.n86 VTAIL.n62 1.93989
R535 VTAIL.n100 VTAIL.n56 1.93989
R536 VTAIL.n140 VTAIL.n116 1.93989
R537 VTAIL.n154 VTAIL.n110 1.93989
R538 VTAIL.n370 VTAIL.n326 1.93989
R539 VTAIL.n357 VTAIL.n333 1.93989
R540 VTAIL.n316 VTAIL.n272 1.93989
R541 VTAIL.n303 VTAIL.n279 1.93989
R542 VTAIL.n262 VTAIL.n218 1.93989
R543 VTAIL.n249 VTAIL.n225 1.93989
R544 VTAIL.n208 VTAIL.n164 1.93989
R545 VTAIL.n195 VTAIL.n171 1.93989
R546 VTAIL VTAIL.n53 1.82162
R547 VTAIL VTAIL.n431 1.70524
R548 VTAIL.n415 VTAIL.n413 1.16414
R549 VTAIL.n423 VTAIL.n382 1.16414
R550 VTAIL.n37 VTAIL.n35 1.16414
R551 VTAIL.n45 VTAIL.n4 1.16414
R552 VTAIL.n91 VTAIL.n89 1.16414
R553 VTAIL.n99 VTAIL.n58 1.16414
R554 VTAIL.n145 VTAIL.n143 1.16414
R555 VTAIL.n153 VTAIL.n112 1.16414
R556 VTAIL.n369 VTAIL.n328 1.16414
R557 VTAIL.n361 VTAIL.n360 1.16414
R558 VTAIL.n315 VTAIL.n274 1.16414
R559 VTAIL.n307 VTAIL.n306 1.16414
R560 VTAIL.n261 VTAIL.n220 1.16414
R561 VTAIL.n253 VTAIL.n252 1.16414
R562 VTAIL.n207 VTAIL.n166 1.16414
R563 VTAIL.n199 VTAIL.n198 1.16414
R564 VTAIL.n323 VTAIL.n269 0.470328
R565 VTAIL.n107 VTAIL.n53 0.470328
R566 VTAIL.n414 VTAIL.n384 0.388379
R567 VTAIL.n420 VTAIL.n419 0.388379
R568 VTAIL.n36 VTAIL.n6 0.388379
R569 VTAIL.n42 VTAIL.n41 0.388379
R570 VTAIL.n90 VTAIL.n60 0.388379
R571 VTAIL.n96 VTAIL.n95 0.388379
R572 VTAIL.n144 VTAIL.n114 0.388379
R573 VTAIL.n150 VTAIL.n149 0.388379
R574 VTAIL.n366 VTAIL.n365 0.388379
R575 VTAIL.n332 VTAIL.n330 0.388379
R576 VTAIL.n312 VTAIL.n311 0.388379
R577 VTAIL.n278 VTAIL.n276 0.388379
R578 VTAIL.n258 VTAIL.n257 0.388379
R579 VTAIL.n224 VTAIL.n222 0.388379
R580 VTAIL.n204 VTAIL.n203 0.388379
R581 VTAIL.n170 VTAIL.n168 0.388379
R582 VTAIL.n396 VTAIL.n391 0.155672
R583 VTAIL.n403 VTAIL.n391 0.155672
R584 VTAIL.n404 VTAIL.n403 0.155672
R585 VTAIL.n404 VTAIL.n387 0.155672
R586 VTAIL.n411 VTAIL.n387 0.155672
R587 VTAIL.n412 VTAIL.n411 0.155672
R588 VTAIL.n412 VTAIL.n383 0.155672
R589 VTAIL.n421 VTAIL.n383 0.155672
R590 VTAIL.n422 VTAIL.n421 0.155672
R591 VTAIL.n422 VTAIL.n379 0.155672
R592 VTAIL.n429 VTAIL.n379 0.155672
R593 VTAIL.n18 VTAIL.n13 0.155672
R594 VTAIL.n25 VTAIL.n13 0.155672
R595 VTAIL.n26 VTAIL.n25 0.155672
R596 VTAIL.n26 VTAIL.n9 0.155672
R597 VTAIL.n33 VTAIL.n9 0.155672
R598 VTAIL.n34 VTAIL.n33 0.155672
R599 VTAIL.n34 VTAIL.n5 0.155672
R600 VTAIL.n43 VTAIL.n5 0.155672
R601 VTAIL.n44 VTAIL.n43 0.155672
R602 VTAIL.n44 VTAIL.n1 0.155672
R603 VTAIL.n51 VTAIL.n1 0.155672
R604 VTAIL.n72 VTAIL.n67 0.155672
R605 VTAIL.n79 VTAIL.n67 0.155672
R606 VTAIL.n80 VTAIL.n79 0.155672
R607 VTAIL.n80 VTAIL.n63 0.155672
R608 VTAIL.n87 VTAIL.n63 0.155672
R609 VTAIL.n88 VTAIL.n87 0.155672
R610 VTAIL.n88 VTAIL.n59 0.155672
R611 VTAIL.n97 VTAIL.n59 0.155672
R612 VTAIL.n98 VTAIL.n97 0.155672
R613 VTAIL.n98 VTAIL.n55 0.155672
R614 VTAIL.n105 VTAIL.n55 0.155672
R615 VTAIL.n126 VTAIL.n121 0.155672
R616 VTAIL.n133 VTAIL.n121 0.155672
R617 VTAIL.n134 VTAIL.n133 0.155672
R618 VTAIL.n134 VTAIL.n117 0.155672
R619 VTAIL.n141 VTAIL.n117 0.155672
R620 VTAIL.n142 VTAIL.n141 0.155672
R621 VTAIL.n142 VTAIL.n113 0.155672
R622 VTAIL.n151 VTAIL.n113 0.155672
R623 VTAIL.n152 VTAIL.n151 0.155672
R624 VTAIL.n152 VTAIL.n109 0.155672
R625 VTAIL.n159 VTAIL.n109 0.155672
R626 VTAIL.n375 VTAIL.n325 0.155672
R627 VTAIL.n368 VTAIL.n325 0.155672
R628 VTAIL.n368 VTAIL.n367 0.155672
R629 VTAIL.n367 VTAIL.n329 0.155672
R630 VTAIL.n359 VTAIL.n329 0.155672
R631 VTAIL.n359 VTAIL.n358 0.155672
R632 VTAIL.n358 VTAIL.n334 0.155672
R633 VTAIL.n351 VTAIL.n334 0.155672
R634 VTAIL.n351 VTAIL.n350 0.155672
R635 VTAIL.n350 VTAIL.n338 0.155672
R636 VTAIL.n343 VTAIL.n338 0.155672
R637 VTAIL.n321 VTAIL.n271 0.155672
R638 VTAIL.n314 VTAIL.n271 0.155672
R639 VTAIL.n314 VTAIL.n313 0.155672
R640 VTAIL.n313 VTAIL.n275 0.155672
R641 VTAIL.n305 VTAIL.n275 0.155672
R642 VTAIL.n305 VTAIL.n304 0.155672
R643 VTAIL.n304 VTAIL.n280 0.155672
R644 VTAIL.n297 VTAIL.n280 0.155672
R645 VTAIL.n297 VTAIL.n296 0.155672
R646 VTAIL.n296 VTAIL.n284 0.155672
R647 VTAIL.n289 VTAIL.n284 0.155672
R648 VTAIL.n267 VTAIL.n217 0.155672
R649 VTAIL.n260 VTAIL.n217 0.155672
R650 VTAIL.n260 VTAIL.n259 0.155672
R651 VTAIL.n259 VTAIL.n221 0.155672
R652 VTAIL.n251 VTAIL.n221 0.155672
R653 VTAIL.n251 VTAIL.n250 0.155672
R654 VTAIL.n250 VTAIL.n226 0.155672
R655 VTAIL.n243 VTAIL.n226 0.155672
R656 VTAIL.n243 VTAIL.n242 0.155672
R657 VTAIL.n242 VTAIL.n230 0.155672
R658 VTAIL.n235 VTAIL.n230 0.155672
R659 VTAIL.n213 VTAIL.n163 0.155672
R660 VTAIL.n206 VTAIL.n163 0.155672
R661 VTAIL.n206 VTAIL.n205 0.155672
R662 VTAIL.n205 VTAIL.n167 0.155672
R663 VTAIL.n197 VTAIL.n167 0.155672
R664 VTAIL.n197 VTAIL.n196 0.155672
R665 VTAIL.n196 VTAIL.n172 0.155672
R666 VTAIL.n189 VTAIL.n172 0.155672
R667 VTAIL.n189 VTAIL.n188 0.155672
R668 VTAIL.n188 VTAIL.n176 0.155672
R669 VTAIL.n181 VTAIL.n176 0.155672
R670 B.n770 B.n769 585
R671 B.n771 B.n770 585
R672 B.n286 B.n123 585
R673 B.n285 B.n284 585
R674 B.n283 B.n282 585
R675 B.n281 B.n280 585
R676 B.n279 B.n278 585
R677 B.n277 B.n276 585
R678 B.n275 B.n274 585
R679 B.n273 B.n272 585
R680 B.n271 B.n270 585
R681 B.n269 B.n268 585
R682 B.n267 B.n266 585
R683 B.n265 B.n264 585
R684 B.n263 B.n262 585
R685 B.n261 B.n260 585
R686 B.n259 B.n258 585
R687 B.n257 B.n256 585
R688 B.n255 B.n254 585
R689 B.n253 B.n252 585
R690 B.n251 B.n250 585
R691 B.n249 B.n248 585
R692 B.n247 B.n246 585
R693 B.n245 B.n244 585
R694 B.n243 B.n242 585
R695 B.n241 B.n240 585
R696 B.n239 B.n238 585
R697 B.n237 B.n236 585
R698 B.n235 B.n234 585
R699 B.n233 B.n232 585
R700 B.n231 B.n230 585
R701 B.n229 B.n228 585
R702 B.n227 B.n226 585
R703 B.n225 B.n224 585
R704 B.n223 B.n222 585
R705 B.n221 B.n220 585
R706 B.n219 B.n218 585
R707 B.n216 B.n215 585
R708 B.n214 B.n213 585
R709 B.n212 B.n211 585
R710 B.n210 B.n209 585
R711 B.n208 B.n207 585
R712 B.n206 B.n205 585
R713 B.n204 B.n203 585
R714 B.n202 B.n201 585
R715 B.n200 B.n199 585
R716 B.n198 B.n197 585
R717 B.n196 B.n195 585
R718 B.n194 B.n193 585
R719 B.n192 B.n191 585
R720 B.n190 B.n189 585
R721 B.n188 B.n187 585
R722 B.n186 B.n185 585
R723 B.n184 B.n183 585
R724 B.n182 B.n181 585
R725 B.n180 B.n179 585
R726 B.n178 B.n177 585
R727 B.n176 B.n175 585
R728 B.n174 B.n173 585
R729 B.n172 B.n171 585
R730 B.n170 B.n169 585
R731 B.n168 B.n167 585
R732 B.n166 B.n165 585
R733 B.n164 B.n163 585
R734 B.n162 B.n161 585
R735 B.n160 B.n159 585
R736 B.n158 B.n157 585
R737 B.n156 B.n155 585
R738 B.n154 B.n153 585
R739 B.n152 B.n151 585
R740 B.n150 B.n149 585
R741 B.n148 B.n147 585
R742 B.n146 B.n145 585
R743 B.n144 B.n143 585
R744 B.n142 B.n141 585
R745 B.n140 B.n139 585
R746 B.n138 B.n137 585
R747 B.n136 B.n135 585
R748 B.n134 B.n133 585
R749 B.n132 B.n131 585
R750 B.n130 B.n129 585
R751 B.n81 B.n80 585
R752 B.n768 B.n82 585
R753 B.n772 B.n82 585
R754 B.n767 B.n766 585
R755 B.n766 B.n78 585
R756 B.n765 B.n77 585
R757 B.n778 B.n77 585
R758 B.n764 B.n76 585
R759 B.n779 B.n76 585
R760 B.n763 B.n75 585
R761 B.n780 B.n75 585
R762 B.n762 B.n761 585
R763 B.n761 B.n71 585
R764 B.n760 B.n70 585
R765 B.n786 B.n70 585
R766 B.n759 B.n69 585
R767 B.n787 B.n69 585
R768 B.n758 B.n68 585
R769 B.n788 B.n68 585
R770 B.n757 B.n756 585
R771 B.n756 B.n67 585
R772 B.n755 B.n63 585
R773 B.n794 B.n63 585
R774 B.n754 B.n62 585
R775 B.n795 B.n62 585
R776 B.n753 B.n61 585
R777 B.n796 B.n61 585
R778 B.n752 B.n751 585
R779 B.n751 B.n57 585
R780 B.n750 B.n56 585
R781 B.n802 B.n56 585
R782 B.n749 B.n55 585
R783 B.n803 B.n55 585
R784 B.n748 B.n54 585
R785 B.n804 B.n54 585
R786 B.n747 B.n746 585
R787 B.n746 B.n50 585
R788 B.n745 B.n49 585
R789 B.n810 B.n49 585
R790 B.n744 B.n48 585
R791 B.n811 B.n48 585
R792 B.n743 B.n47 585
R793 B.n812 B.n47 585
R794 B.n742 B.n741 585
R795 B.n741 B.n43 585
R796 B.n740 B.n42 585
R797 B.n818 B.n42 585
R798 B.n739 B.n41 585
R799 B.n819 B.n41 585
R800 B.n738 B.n40 585
R801 B.n820 B.n40 585
R802 B.n737 B.n736 585
R803 B.n736 B.n36 585
R804 B.n735 B.n35 585
R805 B.n826 B.n35 585
R806 B.n734 B.n34 585
R807 B.n827 B.n34 585
R808 B.n733 B.n33 585
R809 B.n828 B.n33 585
R810 B.n732 B.n731 585
R811 B.n731 B.n29 585
R812 B.n730 B.n28 585
R813 B.n834 B.n28 585
R814 B.n729 B.n27 585
R815 B.n835 B.n27 585
R816 B.n728 B.n26 585
R817 B.n836 B.n26 585
R818 B.n727 B.n726 585
R819 B.n726 B.n22 585
R820 B.n725 B.n21 585
R821 B.n842 B.n21 585
R822 B.n724 B.n20 585
R823 B.n843 B.n20 585
R824 B.n723 B.n19 585
R825 B.n844 B.n19 585
R826 B.n722 B.n721 585
R827 B.n721 B.n15 585
R828 B.n720 B.n14 585
R829 B.n850 B.n14 585
R830 B.n719 B.n13 585
R831 B.n851 B.n13 585
R832 B.n718 B.n12 585
R833 B.n852 B.n12 585
R834 B.n717 B.n716 585
R835 B.n716 B.n8 585
R836 B.n715 B.n7 585
R837 B.n858 B.n7 585
R838 B.n714 B.n6 585
R839 B.n859 B.n6 585
R840 B.n713 B.n5 585
R841 B.n860 B.n5 585
R842 B.n712 B.n711 585
R843 B.n711 B.n4 585
R844 B.n710 B.n287 585
R845 B.n710 B.n709 585
R846 B.n700 B.n288 585
R847 B.n289 B.n288 585
R848 B.n702 B.n701 585
R849 B.n703 B.n702 585
R850 B.n699 B.n294 585
R851 B.n294 B.n293 585
R852 B.n698 B.n697 585
R853 B.n697 B.n696 585
R854 B.n296 B.n295 585
R855 B.n297 B.n296 585
R856 B.n689 B.n688 585
R857 B.n690 B.n689 585
R858 B.n687 B.n302 585
R859 B.n302 B.n301 585
R860 B.n686 B.n685 585
R861 B.n685 B.n684 585
R862 B.n304 B.n303 585
R863 B.n305 B.n304 585
R864 B.n677 B.n676 585
R865 B.n678 B.n677 585
R866 B.n675 B.n310 585
R867 B.n310 B.n309 585
R868 B.n674 B.n673 585
R869 B.n673 B.n672 585
R870 B.n312 B.n311 585
R871 B.n313 B.n312 585
R872 B.n665 B.n664 585
R873 B.n666 B.n665 585
R874 B.n663 B.n318 585
R875 B.n318 B.n317 585
R876 B.n662 B.n661 585
R877 B.n661 B.n660 585
R878 B.n320 B.n319 585
R879 B.n321 B.n320 585
R880 B.n653 B.n652 585
R881 B.n654 B.n653 585
R882 B.n651 B.n326 585
R883 B.n326 B.n325 585
R884 B.n650 B.n649 585
R885 B.n649 B.n648 585
R886 B.n328 B.n327 585
R887 B.n329 B.n328 585
R888 B.n641 B.n640 585
R889 B.n642 B.n641 585
R890 B.n639 B.n334 585
R891 B.n334 B.n333 585
R892 B.n638 B.n637 585
R893 B.n637 B.n636 585
R894 B.n336 B.n335 585
R895 B.n337 B.n336 585
R896 B.n629 B.n628 585
R897 B.n630 B.n629 585
R898 B.n627 B.n342 585
R899 B.n342 B.n341 585
R900 B.n626 B.n625 585
R901 B.n625 B.n624 585
R902 B.n344 B.n343 585
R903 B.n345 B.n344 585
R904 B.n617 B.n616 585
R905 B.n618 B.n617 585
R906 B.n615 B.n350 585
R907 B.n350 B.n349 585
R908 B.n614 B.n613 585
R909 B.n613 B.n612 585
R910 B.n352 B.n351 585
R911 B.n605 B.n352 585
R912 B.n604 B.n603 585
R913 B.n606 B.n604 585
R914 B.n602 B.n357 585
R915 B.n357 B.n356 585
R916 B.n601 B.n600 585
R917 B.n600 B.n599 585
R918 B.n359 B.n358 585
R919 B.n360 B.n359 585
R920 B.n592 B.n591 585
R921 B.n593 B.n592 585
R922 B.n590 B.n365 585
R923 B.n365 B.n364 585
R924 B.n589 B.n588 585
R925 B.n588 B.n587 585
R926 B.n367 B.n366 585
R927 B.n368 B.n367 585
R928 B.n580 B.n579 585
R929 B.n581 B.n580 585
R930 B.n371 B.n370 585
R931 B.n419 B.n417 585
R932 B.n420 B.n416 585
R933 B.n420 B.n372 585
R934 B.n423 B.n422 585
R935 B.n424 B.n415 585
R936 B.n426 B.n425 585
R937 B.n428 B.n414 585
R938 B.n431 B.n430 585
R939 B.n432 B.n413 585
R940 B.n434 B.n433 585
R941 B.n436 B.n412 585
R942 B.n439 B.n438 585
R943 B.n440 B.n411 585
R944 B.n442 B.n441 585
R945 B.n444 B.n410 585
R946 B.n447 B.n446 585
R947 B.n448 B.n409 585
R948 B.n450 B.n449 585
R949 B.n452 B.n408 585
R950 B.n455 B.n454 585
R951 B.n456 B.n407 585
R952 B.n458 B.n457 585
R953 B.n460 B.n406 585
R954 B.n463 B.n462 585
R955 B.n464 B.n405 585
R956 B.n466 B.n465 585
R957 B.n468 B.n404 585
R958 B.n471 B.n470 585
R959 B.n472 B.n403 585
R960 B.n474 B.n473 585
R961 B.n476 B.n402 585
R962 B.n479 B.n478 585
R963 B.n480 B.n401 585
R964 B.n482 B.n481 585
R965 B.n484 B.n400 585
R966 B.n487 B.n486 585
R967 B.n489 B.n397 585
R968 B.n491 B.n490 585
R969 B.n493 B.n396 585
R970 B.n496 B.n495 585
R971 B.n497 B.n395 585
R972 B.n499 B.n498 585
R973 B.n501 B.n394 585
R974 B.n504 B.n503 585
R975 B.n505 B.n391 585
R976 B.n508 B.n507 585
R977 B.n510 B.n390 585
R978 B.n513 B.n512 585
R979 B.n514 B.n389 585
R980 B.n516 B.n515 585
R981 B.n518 B.n388 585
R982 B.n521 B.n520 585
R983 B.n522 B.n387 585
R984 B.n524 B.n523 585
R985 B.n526 B.n386 585
R986 B.n529 B.n528 585
R987 B.n530 B.n385 585
R988 B.n532 B.n531 585
R989 B.n534 B.n384 585
R990 B.n537 B.n536 585
R991 B.n538 B.n383 585
R992 B.n540 B.n539 585
R993 B.n542 B.n382 585
R994 B.n545 B.n544 585
R995 B.n546 B.n381 585
R996 B.n548 B.n547 585
R997 B.n550 B.n380 585
R998 B.n553 B.n552 585
R999 B.n554 B.n379 585
R1000 B.n556 B.n555 585
R1001 B.n558 B.n378 585
R1002 B.n561 B.n560 585
R1003 B.n562 B.n377 585
R1004 B.n564 B.n563 585
R1005 B.n566 B.n376 585
R1006 B.n569 B.n568 585
R1007 B.n570 B.n375 585
R1008 B.n572 B.n571 585
R1009 B.n574 B.n374 585
R1010 B.n577 B.n576 585
R1011 B.n578 B.n373 585
R1012 B.n583 B.n582 585
R1013 B.n582 B.n581 585
R1014 B.n584 B.n369 585
R1015 B.n369 B.n368 585
R1016 B.n586 B.n585 585
R1017 B.n587 B.n586 585
R1018 B.n363 B.n362 585
R1019 B.n364 B.n363 585
R1020 B.n595 B.n594 585
R1021 B.n594 B.n593 585
R1022 B.n596 B.n361 585
R1023 B.n361 B.n360 585
R1024 B.n598 B.n597 585
R1025 B.n599 B.n598 585
R1026 B.n355 B.n354 585
R1027 B.n356 B.n355 585
R1028 B.n608 B.n607 585
R1029 B.n607 B.n606 585
R1030 B.n609 B.n353 585
R1031 B.n605 B.n353 585
R1032 B.n611 B.n610 585
R1033 B.n612 B.n611 585
R1034 B.n348 B.n347 585
R1035 B.n349 B.n348 585
R1036 B.n620 B.n619 585
R1037 B.n619 B.n618 585
R1038 B.n621 B.n346 585
R1039 B.n346 B.n345 585
R1040 B.n623 B.n622 585
R1041 B.n624 B.n623 585
R1042 B.n340 B.n339 585
R1043 B.n341 B.n340 585
R1044 B.n632 B.n631 585
R1045 B.n631 B.n630 585
R1046 B.n633 B.n338 585
R1047 B.n338 B.n337 585
R1048 B.n635 B.n634 585
R1049 B.n636 B.n635 585
R1050 B.n332 B.n331 585
R1051 B.n333 B.n332 585
R1052 B.n644 B.n643 585
R1053 B.n643 B.n642 585
R1054 B.n645 B.n330 585
R1055 B.n330 B.n329 585
R1056 B.n647 B.n646 585
R1057 B.n648 B.n647 585
R1058 B.n324 B.n323 585
R1059 B.n325 B.n324 585
R1060 B.n656 B.n655 585
R1061 B.n655 B.n654 585
R1062 B.n657 B.n322 585
R1063 B.n322 B.n321 585
R1064 B.n659 B.n658 585
R1065 B.n660 B.n659 585
R1066 B.n316 B.n315 585
R1067 B.n317 B.n316 585
R1068 B.n668 B.n667 585
R1069 B.n667 B.n666 585
R1070 B.n669 B.n314 585
R1071 B.n314 B.n313 585
R1072 B.n671 B.n670 585
R1073 B.n672 B.n671 585
R1074 B.n308 B.n307 585
R1075 B.n309 B.n308 585
R1076 B.n680 B.n679 585
R1077 B.n679 B.n678 585
R1078 B.n681 B.n306 585
R1079 B.n306 B.n305 585
R1080 B.n683 B.n682 585
R1081 B.n684 B.n683 585
R1082 B.n300 B.n299 585
R1083 B.n301 B.n300 585
R1084 B.n692 B.n691 585
R1085 B.n691 B.n690 585
R1086 B.n693 B.n298 585
R1087 B.n298 B.n297 585
R1088 B.n695 B.n694 585
R1089 B.n696 B.n695 585
R1090 B.n292 B.n291 585
R1091 B.n293 B.n292 585
R1092 B.n705 B.n704 585
R1093 B.n704 B.n703 585
R1094 B.n706 B.n290 585
R1095 B.n290 B.n289 585
R1096 B.n708 B.n707 585
R1097 B.n709 B.n708 585
R1098 B.n2 B.n0 585
R1099 B.n4 B.n2 585
R1100 B.n3 B.n1 585
R1101 B.n859 B.n3 585
R1102 B.n857 B.n856 585
R1103 B.n858 B.n857 585
R1104 B.n855 B.n9 585
R1105 B.n9 B.n8 585
R1106 B.n854 B.n853 585
R1107 B.n853 B.n852 585
R1108 B.n11 B.n10 585
R1109 B.n851 B.n11 585
R1110 B.n849 B.n848 585
R1111 B.n850 B.n849 585
R1112 B.n847 B.n16 585
R1113 B.n16 B.n15 585
R1114 B.n846 B.n845 585
R1115 B.n845 B.n844 585
R1116 B.n18 B.n17 585
R1117 B.n843 B.n18 585
R1118 B.n841 B.n840 585
R1119 B.n842 B.n841 585
R1120 B.n839 B.n23 585
R1121 B.n23 B.n22 585
R1122 B.n838 B.n837 585
R1123 B.n837 B.n836 585
R1124 B.n25 B.n24 585
R1125 B.n835 B.n25 585
R1126 B.n833 B.n832 585
R1127 B.n834 B.n833 585
R1128 B.n831 B.n30 585
R1129 B.n30 B.n29 585
R1130 B.n830 B.n829 585
R1131 B.n829 B.n828 585
R1132 B.n32 B.n31 585
R1133 B.n827 B.n32 585
R1134 B.n825 B.n824 585
R1135 B.n826 B.n825 585
R1136 B.n823 B.n37 585
R1137 B.n37 B.n36 585
R1138 B.n822 B.n821 585
R1139 B.n821 B.n820 585
R1140 B.n39 B.n38 585
R1141 B.n819 B.n39 585
R1142 B.n817 B.n816 585
R1143 B.n818 B.n817 585
R1144 B.n815 B.n44 585
R1145 B.n44 B.n43 585
R1146 B.n814 B.n813 585
R1147 B.n813 B.n812 585
R1148 B.n46 B.n45 585
R1149 B.n811 B.n46 585
R1150 B.n809 B.n808 585
R1151 B.n810 B.n809 585
R1152 B.n807 B.n51 585
R1153 B.n51 B.n50 585
R1154 B.n806 B.n805 585
R1155 B.n805 B.n804 585
R1156 B.n53 B.n52 585
R1157 B.n803 B.n53 585
R1158 B.n801 B.n800 585
R1159 B.n802 B.n801 585
R1160 B.n799 B.n58 585
R1161 B.n58 B.n57 585
R1162 B.n798 B.n797 585
R1163 B.n797 B.n796 585
R1164 B.n60 B.n59 585
R1165 B.n795 B.n60 585
R1166 B.n793 B.n792 585
R1167 B.n794 B.n793 585
R1168 B.n791 B.n64 585
R1169 B.n67 B.n64 585
R1170 B.n790 B.n789 585
R1171 B.n789 B.n788 585
R1172 B.n66 B.n65 585
R1173 B.n787 B.n66 585
R1174 B.n785 B.n784 585
R1175 B.n786 B.n785 585
R1176 B.n783 B.n72 585
R1177 B.n72 B.n71 585
R1178 B.n782 B.n781 585
R1179 B.n781 B.n780 585
R1180 B.n74 B.n73 585
R1181 B.n779 B.n74 585
R1182 B.n777 B.n776 585
R1183 B.n778 B.n777 585
R1184 B.n775 B.n79 585
R1185 B.n79 B.n78 585
R1186 B.n774 B.n773 585
R1187 B.n773 B.n772 585
R1188 B.n862 B.n861 585
R1189 B.n861 B.n860 585
R1190 B.n582 B.n371 569.379
R1191 B.n773 B.n81 569.379
R1192 B.n580 B.n373 569.379
R1193 B.n770 B.n82 569.379
R1194 B.n392 B.t7 328.325
R1195 B.n124 B.t16 328.325
R1196 B.n398 B.t10 328.325
R1197 B.n126 B.t13 328.325
R1198 B.n392 B.t4 273.858
R1199 B.n398 B.t8 273.858
R1200 B.n126 B.t11 273.858
R1201 B.n124 B.t15 273.858
R1202 B.n771 B.n122 256.663
R1203 B.n771 B.n121 256.663
R1204 B.n771 B.n120 256.663
R1205 B.n771 B.n119 256.663
R1206 B.n771 B.n118 256.663
R1207 B.n771 B.n117 256.663
R1208 B.n771 B.n116 256.663
R1209 B.n771 B.n115 256.663
R1210 B.n771 B.n114 256.663
R1211 B.n771 B.n113 256.663
R1212 B.n771 B.n112 256.663
R1213 B.n771 B.n111 256.663
R1214 B.n771 B.n110 256.663
R1215 B.n771 B.n109 256.663
R1216 B.n771 B.n108 256.663
R1217 B.n771 B.n107 256.663
R1218 B.n771 B.n106 256.663
R1219 B.n771 B.n105 256.663
R1220 B.n771 B.n104 256.663
R1221 B.n771 B.n103 256.663
R1222 B.n771 B.n102 256.663
R1223 B.n771 B.n101 256.663
R1224 B.n771 B.n100 256.663
R1225 B.n771 B.n99 256.663
R1226 B.n771 B.n98 256.663
R1227 B.n771 B.n97 256.663
R1228 B.n771 B.n96 256.663
R1229 B.n771 B.n95 256.663
R1230 B.n771 B.n94 256.663
R1231 B.n771 B.n93 256.663
R1232 B.n771 B.n92 256.663
R1233 B.n771 B.n91 256.663
R1234 B.n771 B.n90 256.663
R1235 B.n771 B.n89 256.663
R1236 B.n771 B.n88 256.663
R1237 B.n771 B.n87 256.663
R1238 B.n771 B.n86 256.663
R1239 B.n771 B.n85 256.663
R1240 B.n771 B.n84 256.663
R1241 B.n771 B.n83 256.663
R1242 B.n418 B.n372 256.663
R1243 B.n421 B.n372 256.663
R1244 B.n427 B.n372 256.663
R1245 B.n429 B.n372 256.663
R1246 B.n435 B.n372 256.663
R1247 B.n437 B.n372 256.663
R1248 B.n443 B.n372 256.663
R1249 B.n445 B.n372 256.663
R1250 B.n451 B.n372 256.663
R1251 B.n453 B.n372 256.663
R1252 B.n459 B.n372 256.663
R1253 B.n461 B.n372 256.663
R1254 B.n467 B.n372 256.663
R1255 B.n469 B.n372 256.663
R1256 B.n475 B.n372 256.663
R1257 B.n477 B.n372 256.663
R1258 B.n483 B.n372 256.663
R1259 B.n485 B.n372 256.663
R1260 B.n492 B.n372 256.663
R1261 B.n494 B.n372 256.663
R1262 B.n500 B.n372 256.663
R1263 B.n502 B.n372 256.663
R1264 B.n509 B.n372 256.663
R1265 B.n511 B.n372 256.663
R1266 B.n517 B.n372 256.663
R1267 B.n519 B.n372 256.663
R1268 B.n525 B.n372 256.663
R1269 B.n527 B.n372 256.663
R1270 B.n533 B.n372 256.663
R1271 B.n535 B.n372 256.663
R1272 B.n541 B.n372 256.663
R1273 B.n543 B.n372 256.663
R1274 B.n549 B.n372 256.663
R1275 B.n551 B.n372 256.663
R1276 B.n557 B.n372 256.663
R1277 B.n559 B.n372 256.663
R1278 B.n565 B.n372 256.663
R1279 B.n567 B.n372 256.663
R1280 B.n573 B.n372 256.663
R1281 B.n575 B.n372 256.663
R1282 B.n393 B.t6 249.005
R1283 B.n125 B.t17 249.005
R1284 B.n399 B.t9 249.005
R1285 B.n127 B.t14 249.005
R1286 B.n582 B.n369 163.367
R1287 B.n586 B.n369 163.367
R1288 B.n586 B.n363 163.367
R1289 B.n594 B.n363 163.367
R1290 B.n594 B.n361 163.367
R1291 B.n598 B.n361 163.367
R1292 B.n598 B.n355 163.367
R1293 B.n607 B.n355 163.367
R1294 B.n607 B.n353 163.367
R1295 B.n611 B.n353 163.367
R1296 B.n611 B.n348 163.367
R1297 B.n619 B.n348 163.367
R1298 B.n619 B.n346 163.367
R1299 B.n623 B.n346 163.367
R1300 B.n623 B.n340 163.367
R1301 B.n631 B.n340 163.367
R1302 B.n631 B.n338 163.367
R1303 B.n635 B.n338 163.367
R1304 B.n635 B.n332 163.367
R1305 B.n643 B.n332 163.367
R1306 B.n643 B.n330 163.367
R1307 B.n647 B.n330 163.367
R1308 B.n647 B.n324 163.367
R1309 B.n655 B.n324 163.367
R1310 B.n655 B.n322 163.367
R1311 B.n659 B.n322 163.367
R1312 B.n659 B.n316 163.367
R1313 B.n667 B.n316 163.367
R1314 B.n667 B.n314 163.367
R1315 B.n671 B.n314 163.367
R1316 B.n671 B.n308 163.367
R1317 B.n679 B.n308 163.367
R1318 B.n679 B.n306 163.367
R1319 B.n683 B.n306 163.367
R1320 B.n683 B.n300 163.367
R1321 B.n691 B.n300 163.367
R1322 B.n691 B.n298 163.367
R1323 B.n695 B.n298 163.367
R1324 B.n695 B.n292 163.367
R1325 B.n704 B.n292 163.367
R1326 B.n704 B.n290 163.367
R1327 B.n708 B.n290 163.367
R1328 B.n708 B.n2 163.367
R1329 B.n861 B.n2 163.367
R1330 B.n861 B.n3 163.367
R1331 B.n857 B.n3 163.367
R1332 B.n857 B.n9 163.367
R1333 B.n853 B.n9 163.367
R1334 B.n853 B.n11 163.367
R1335 B.n849 B.n11 163.367
R1336 B.n849 B.n16 163.367
R1337 B.n845 B.n16 163.367
R1338 B.n845 B.n18 163.367
R1339 B.n841 B.n18 163.367
R1340 B.n841 B.n23 163.367
R1341 B.n837 B.n23 163.367
R1342 B.n837 B.n25 163.367
R1343 B.n833 B.n25 163.367
R1344 B.n833 B.n30 163.367
R1345 B.n829 B.n30 163.367
R1346 B.n829 B.n32 163.367
R1347 B.n825 B.n32 163.367
R1348 B.n825 B.n37 163.367
R1349 B.n821 B.n37 163.367
R1350 B.n821 B.n39 163.367
R1351 B.n817 B.n39 163.367
R1352 B.n817 B.n44 163.367
R1353 B.n813 B.n44 163.367
R1354 B.n813 B.n46 163.367
R1355 B.n809 B.n46 163.367
R1356 B.n809 B.n51 163.367
R1357 B.n805 B.n51 163.367
R1358 B.n805 B.n53 163.367
R1359 B.n801 B.n53 163.367
R1360 B.n801 B.n58 163.367
R1361 B.n797 B.n58 163.367
R1362 B.n797 B.n60 163.367
R1363 B.n793 B.n60 163.367
R1364 B.n793 B.n64 163.367
R1365 B.n789 B.n64 163.367
R1366 B.n789 B.n66 163.367
R1367 B.n785 B.n66 163.367
R1368 B.n785 B.n72 163.367
R1369 B.n781 B.n72 163.367
R1370 B.n781 B.n74 163.367
R1371 B.n777 B.n74 163.367
R1372 B.n777 B.n79 163.367
R1373 B.n773 B.n79 163.367
R1374 B.n420 B.n419 163.367
R1375 B.n422 B.n420 163.367
R1376 B.n426 B.n415 163.367
R1377 B.n430 B.n428 163.367
R1378 B.n434 B.n413 163.367
R1379 B.n438 B.n436 163.367
R1380 B.n442 B.n411 163.367
R1381 B.n446 B.n444 163.367
R1382 B.n450 B.n409 163.367
R1383 B.n454 B.n452 163.367
R1384 B.n458 B.n407 163.367
R1385 B.n462 B.n460 163.367
R1386 B.n466 B.n405 163.367
R1387 B.n470 B.n468 163.367
R1388 B.n474 B.n403 163.367
R1389 B.n478 B.n476 163.367
R1390 B.n482 B.n401 163.367
R1391 B.n486 B.n484 163.367
R1392 B.n491 B.n397 163.367
R1393 B.n495 B.n493 163.367
R1394 B.n499 B.n395 163.367
R1395 B.n503 B.n501 163.367
R1396 B.n508 B.n391 163.367
R1397 B.n512 B.n510 163.367
R1398 B.n516 B.n389 163.367
R1399 B.n520 B.n518 163.367
R1400 B.n524 B.n387 163.367
R1401 B.n528 B.n526 163.367
R1402 B.n532 B.n385 163.367
R1403 B.n536 B.n534 163.367
R1404 B.n540 B.n383 163.367
R1405 B.n544 B.n542 163.367
R1406 B.n548 B.n381 163.367
R1407 B.n552 B.n550 163.367
R1408 B.n556 B.n379 163.367
R1409 B.n560 B.n558 163.367
R1410 B.n564 B.n377 163.367
R1411 B.n568 B.n566 163.367
R1412 B.n572 B.n375 163.367
R1413 B.n576 B.n574 163.367
R1414 B.n580 B.n367 163.367
R1415 B.n588 B.n367 163.367
R1416 B.n588 B.n365 163.367
R1417 B.n592 B.n365 163.367
R1418 B.n592 B.n359 163.367
R1419 B.n600 B.n359 163.367
R1420 B.n600 B.n357 163.367
R1421 B.n604 B.n357 163.367
R1422 B.n604 B.n352 163.367
R1423 B.n613 B.n352 163.367
R1424 B.n613 B.n350 163.367
R1425 B.n617 B.n350 163.367
R1426 B.n617 B.n344 163.367
R1427 B.n625 B.n344 163.367
R1428 B.n625 B.n342 163.367
R1429 B.n629 B.n342 163.367
R1430 B.n629 B.n336 163.367
R1431 B.n637 B.n336 163.367
R1432 B.n637 B.n334 163.367
R1433 B.n641 B.n334 163.367
R1434 B.n641 B.n328 163.367
R1435 B.n649 B.n328 163.367
R1436 B.n649 B.n326 163.367
R1437 B.n653 B.n326 163.367
R1438 B.n653 B.n320 163.367
R1439 B.n661 B.n320 163.367
R1440 B.n661 B.n318 163.367
R1441 B.n665 B.n318 163.367
R1442 B.n665 B.n312 163.367
R1443 B.n673 B.n312 163.367
R1444 B.n673 B.n310 163.367
R1445 B.n677 B.n310 163.367
R1446 B.n677 B.n304 163.367
R1447 B.n685 B.n304 163.367
R1448 B.n685 B.n302 163.367
R1449 B.n689 B.n302 163.367
R1450 B.n689 B.n296 163.367
R1451 B.n697 B.n296 163.367
R1452 B.n697 B.n294 163.367
R1453 B.n702 B.n294 163.367
R1454 B.n702 B.n288 163.367
R1455 B.n710 B.n288 163.367
R1456 B.n711 B.n710 163.367
R1457 B.n711 B.n5 163.367
R1458 B.n6 B.n5 163.367
R1459 B.n7 B.n6 163.367
R1460 B.n716 B.n7 163.367
R1461 B.n716 B.n12 163.367
R1462 B.n13 B.n12 163.367
R1463 B.n14 B.n13 163.367
R1464 B.n721 B.n14 163.367
R1465 B.n721 B.n19 163.367
R1466 B.n20 B.n19 163.367
R1467 B.n21 B.n20 163.367
R1468 B.n726 B.n21 163.367
R1469 B.n726 B.n26 163.367
R1470 B.n27 B.n26 163.367
R1471 B.n28 B.n27 163.367
R1472 B.n731 B.n28 163.367
R1473 B.n731 B.n33 163.367
R1474 B.n34 B.n33 163.367
R1475 B.n35 B.n34 163.367
R1476 B.n736 B.n35 163.367
R1477 B.n736 B.n40 163.367
R1478 B.n41 B.n40 163.367
R1479 B.n42 B.n41 163.367
R1480 B.n741 B.n42 163.367
R1481 B.n741 B.n47 163.367
R1482 B.n48 B.n47 163.367
R1483 B.n49 B.n48 163.367
R1484 B.n746 B.n49 163.367
R1485 B.n746 B.n54 163.367
R1486 B.n55 B.n54 163.367
R1487 B.n56 B.n55 163.367
R1488 B.n751 B.n56 163.367
R1489 B.n751 B.n61 163.367
R1490 B.n62 B.n61 163.367
R1491 B.n63 B.n62 163.367
R1492 B.n756 B.n63 163.367
R1493 B.n756 B.n68 163.367
R1494 B.n69 B.n68 163.367
R1495 B.n70 B.n69 163.367
R1496 B.n761 B.n70 163.367
R1497 B.n761 B.n75 163.367
R1498 B.n76 B.n75 163.367
R1499 B.n77 B.n76 163.367
R1500 B.n766 B.n77 163.367
R1501 B.n766 B.n82 163.367
R1502 B.n131 B.n130 163.367
R1503 B.n135 B.n134 163.367
R1504 B.n139 B.n138 163.367
R1505 B.n143 B.n142 163.367
R1506 B.n147 B.n146 163.367
R1507 B.n151 B.n150 163.367
R1508 B.n155 B.n154 163.367
R1509 B.n159 B.n158 163.367
R1510 B.n163 B.n162 163.367
R1511 B.n167 B.n166 163.367
R1512 B.n171 B.n170 163.367
R1513 B.n175 B.n174 163.367
R1514 B.n179 B.n178 163.367
R1515 B.n183 B.n182 163.367
R1516 B.n187 B.n186 163.367
R1517 B.n191 B.n190 163.367
R1518 B.n195 B.n194 163.367
R1519 B.n199 B.n198 163.367
R1520 B.n203 B.n202 163.367
R1521 B.n207 B.n206 163.367
R1522 B.n211 B.n210 163.367
R1523 B.n215 B.n214 163.367
R1524 B.n220 B.n219 163.367
R1525 B.n224 B.n223 163.367
R1526 B.n228 B.n227 163.367
R1527 B.n232 B.n231 163.367
R1528 B.n236 B.n235 163.367
R1529 B.n240 B.n239 163.367
R1530 B.n244 B.n243 163.367
R1531 B.n248 B.n247 163.367
R1532 B.n252 B.n251 163.367
R1533 B.n256 B.n255 163.367
R1534 B.n260 B.n259 163.367
R1535 B.n264 B.n263 163.367
R1536 B.n268 B.n267 163.367
R1537 B.n272 B.n271 163.367
R1538 B.n276 B.n275 163.367
R1539 B.n280 B.n279 163.367
R1540 B.n284 B.n283 163.367
R1541 B.n770 B.n123 163.367
R1542 B.n581 B.n372 98.2084
R1543 B.n772 B.n771 98.2084
R1544 B.n393 B.n392 79.3217
R1545 B.n399 B.n398 79.3217
R1546 B.n127 B.n126 79.3217
R1547 B.n125 B.n124 79.3217
R1548 B.n418 B.n371 71.676
R1549 B.n422 B.n421 71.676
R1550 B.n427 B.n426 71.676
R1551 B.n430 B.n429 71.676
R1552 B.n435 B.n434 71.676
R1553 B.n438 B.n437 71.676
R1554 B.n443 B.n442 71.676
R1555 B.n446 B.n445 71.676
R1556 B.n451 B.n450 71.676
R1557 B.n454 B.n453 71.676
R1558 B.n459 B.n458 71.676
R1559 B.n462 B.n461 71.676
R1560 B.n467 B.n466 71.676
R1561 B.n470 B.n469 71.676
R1562 B.n475 B.n474 71.676
R1563 B.n478 B.n477 71.676
R1564 B.n483 B.n482 71.676
R1565 B.n486 B.n485 71.676
R1566 B.n492 B.n491 71.676
R1567 B.n495 B.n494 71.676
R1568 B.n500 B.n499 71.676
R1569 B.n503 B.n502 71.676
R1570 B.n509 B.n508 71.676
R1571 B.n512 B.n511 71.676
R1572 B.n517 B.n516 71.676
R1573 B.n520 B.n519 71.676
R1574 B.n525 B.n524 71.676
R1575 B.n528 B.n527 71.676
R1576 B.n533 B.n532 71.676
R1577 B.n536 B.n535 71.676
R1578 B.n541 B.n540 71.676
R1579 B.n544 B.n543 71.676
R1580 B.n549 B.n548 71.676
R1581 B.n552 B.n551 71.676
R1582 B.n557 B.n556 71.676
R1583 B.n560 B.n559 71.676
R1584 B.n565 B.n564 71.676
R1585 B.n568 B.n567 71.676
R1586 B.n573 B.n572 71.676
R1587 B.n576 B.n575 71.676
R1588 B.n83 B.n81 71.676
R1589 B.n131 B.n84 71.676
R1590 B.n135 B.n85 71.676
R1591 B.n139 B.n86 71.676
R1592 B.n143 B.n87 71.676
R1593 B.n147 B.n88 71.676
R1594 B.n151 B.n89 71.676
R1595 B.n155 B.n90 71.676
R1596 B.n159 B.n91 71.676
R1597 B.n163 B.n92 71.676
R1598 B.n167 B.n93 71.676
R1599 B.n171 B.n94 71.676
R1600 B.n175 B.n95 71.676
R1601 B.n179 B.n96 71.676
R1602 B.n183 B.n97 71.676
R1603 B.n187 B.n98 71.676
R1604 B.n191 B.n99 71.676
R1605 B.n195 B.n100 71.676
R1606 B.n199 B.n101 71.676
R1607 B.n203 B.n102 71.676
R1608 B.n207 B.n103 71.676
R1609 B.n211 B.n104 71.676
R1610 B.n215 B.n105 71.676
R1611 B.n220 B.n106 71.676
R1612 B.n224 B.n107 71.676
R1613 B.n228 B.n108 71.676
R1614 B.n232 B.n109 71.676
R1615 B.n236 B.n110 71.676
R1616 B.n240 B.n111 71.676
R1617 B.n244 B.n112 71.676
R1618 B.n248 B.n113 71.676
R1619 B.n252 B.n114 71.676
R1620 B.n256 B.n115 71.676
R1621 B.n260 B.n116 71.676
R1622 B.n264 B.n117 71.676
R1623 B.n268 B.n118 71.676
R1624 B.n272 B.n119 71.676
R1625 B.n276 B.n120 71.676
R1626 B.n280 B.n121 71.676
R1627 B.n284 B.n122 71.676
R1628 B.n123 B.n122 71.676
R1629 B.n283 B.n121 71.676
R1630 B.n279 B.n120 71.676
R1631 B.n275 B.n119 71.676
R1632 B.n271 B.n118 71.676
R1633 B.n267 B.n117 71.676
R1634 B.n263 B.n116 71.676
R1635 B.n259 B.n115 71.676
R1636 B.n255 B.n114 71.676
R1637 B.n251 B.n113 71.676
R1638 B.n247 B.n112 71.676
R1639 B.n243 B.n111 71.676
R1640 B.n239 B.n110 71.676
R1641 B.n235 B.n109 71.676
R1642 B.n231 B.n108 71.676
R1643 B.n227 B.n107 71.676
R1644 B.n223 B.n106 71.676
R1645 B.n219 B.n105 71.676
R1646 B.n214 B.n104 71.676
R1647 B.n210 B.n103 71.676
R1648 B.n206 B.n102 71.676
R1649 B.n202 B.n101 71.676
R1650 B.n198 B.n100 71.676
R1651 B.n194 B.n99 71.676
R1652 B.n190 B.n98 71.676
R1653 B.n186 B.n97 71.676
R1654 B.n182 B.n96 71.676
R1655 B.n178 B.n95 71.676
R1656 B.n174 B.n94 71.676
R1657 B.n170 B.n93 71.676
R1658 B.n166 B.n92 71.676
R1659 B.n162 B.n91 71.676
R1660 B.n158 B.n90 71.676
R1661 B.n154 B.n89 71.676
R1662 B.n150 B.n88 71.676
R1663 B.n146 B.n87 71.676
R1664 B.n142 B.n86 71.676
R1665 B.n138 B.n85 71.676
R1666 B.n134 B.n84 71.676
R1667 B.n130 B.n83 71.676
R1668 B.n419 B.n418 71.676
R1669 B.n421 B.n415 71.676
R1670 B.n428 B.n427 71.676
R1671 B.n429 B.n413 71.676
R1672 B.n436 B.n435 71.676
R1673 B.n437 B.n411 71.676
R1674 B.n444 B.n443 71.676
R1675 B.n445 B.n409 71.676
R1676 B.n452 B.n451 71.676
R1677 B.n453 B.n407 71.676
R1678 B.n460 B.n459 71.676
R1679 B.n461 B.n405 71.676
R1680 B.n468 B.n467 71.676
R1681 B.n469 B.n403 71.676
R1682 B.n476 B.n475 71.676
R1683 B.n477 B.n401 71.676
R1684 B.n484 B.n483 71.676
R1685 B.n485 B.n397 71.676
R1686 B.n493 B.n492 71.676
R1687 B.n494 B.n395 71.676
R1688 B.n501 B.n500 71.676
R1689 B.n502 B.n391 71.676
R1690 B.n510 B.n509 71.676
R1691 B.n511 B.n389 71.676
R1692 B.n518 B.n517 71.676
R1693 B.n519 B.n387 71.676
R1694 B.n526 B.n525 71.676
R1695 B.n527 B.n385 71.676
R1696 B.n534 B.n533 71.676
R1697 B.n535 B.n383 71.676
R1698 B.n542 B.n541 71.676
R1699 B.n543 B.n381 71.676
R1700 B.n550 B.n549 71.676
R1701 B.n551 B.n379 71.676
R1702 B.n558 B.n557 71.676
R1703 B.n559 B.n377 71.676
R1704 B.n566 B.n565 71.676
R1705 B.n567 B.n375 71.676
R1706 B.n574 B.n573 71.676
R1707 B.n575 B.n373 71.676
R1708 B.n506 B.n393 59.5399
R1709 B.n488 B.n399 59.5399
R1710 B.n128 B.n127 59.5399
R1711 B.n217 B.n125 59.5399
R1712 B.n581 B.n368 48.746
R1713 B.n587 B.n368 48.746
R1714 B.n587 B.n364 48.746
R1715 B.n593 B.n364 48.746
R1716 B.n593 B.n360 48.746
R1717 B.n599 B.n360 48.746
R1718 B.n599 B.n356 48.746
R1719 B.n606 B.n356 48.746
R1720 B.n606 B.n605 48.746
R1721 B.n612 B.n349 48.746
R1722 B.n618 B.n349 48.746
R1723 B.n618 B.n345 48.746
R1724 B.n624 B.n345 48.746
R1725 B.n624 B.n341 48.746
R1726 B.n630 B.n341 48.746
R1727 B.n630 B.n337 48.746
R1728 B.n636 B.n337 48.746
R1729 B.n636 B.n333 48.746
R1730 B.n642 B.n333 48.746
R1731 B.n642 B.n329 48.746
R1732 B.n648 B.n329 48.746
R1733 B.n648 B.n325 48.746
R1734 B.n654 B.n325 48.746
R1735 B.n660 B.n321 48.746
R1736 B.n660 B.n317 48.746
R1737 B.n666 B.n317 48.746
R1738 B.n666 B.n313 48.746
R1739 B.n672 B.n313 48.746
R1740 B.n672 B.n309 48.746
R1741 B.n678 B.n309 48.746
R1742 B.n678 B.n305 48.746
R1743 B.n684 B.n305 48.746
R1744 B.n684 B.n301 48.746
R1745 B.n690 B.n301 48.746
R1746 B.n696 B.n297 48.746
R1747 B.n696 B.n293 48.746
R1748 B.n703 B.n293 48.746
R1749 B.n703 B.n289 48.746
R1750 B.n709 B.n289 48.746
R1751 B.n709 B.n4 48.746
R1752 B.n860 B.n4 48.746
R1753 B.n860 B.n859 48.746
R1754 B.n859 B.n858 48.746
R1755 B.n858 B.n8 48.746
R1756 B.n852 B.n8 48.746
R1757 B.n852 B.n851 48.746
R1758 B.n851 B.n850 48.746
R1759 B.n850 B.n15 48.746
R1760 B.n844 B.n843 48.746
R1761 B.n843 B.n842 48.746
R1762 B.n842 B.n22 48.746
R1763 B.n836 B.n22 48.746
R1764 B.n836 B.n835 48.746
R1765 B.n835 B.n834 48.746
R1766 B.n834 B.n29 48.746
R1767 B.n828 B.n29 48.746
R1768 B.n828 B.n827 48.746
R1769 B.n827 B.n826 48.746
R1770 B.n826 B.n36 48.746
R1771 B.n820 B.n819 48.746
R1772 B.n819 B.n818 48.746
R1773 B.n818 B.n43 48.746
R1774 B.n812 B.n43 48.746
R1775 B.n812 B.n811 48.746
R1776 B.n811 B.n810 48.746
R1777 B.n810 B.n50 48.746
R1778 B.n804 B.n50 48.746
R1779 B.n804 B.n803 48.746
R1780 B.n803 B.n802 48.746
R1781 B.n802 B.n57 48.746
R1782 B.n796 B.n57 48.746
R1783 B.n796 B.n795 48.746
R1784 B.n795 B.n794 48.746
R1785 B.n788 B.n67 48.746
R1786 B.n788 B.n787 48.746
R1787 B.n787 B.n786 48.746
R1788 B.n786 B.n71 48.746
R1789 B.n780 B.n71 48.746
R1790 B.n780 B.n779 48.746
R1791 B.n779 B.n778 48.746
R1792 B.n778 B.n78 48.746
R1793 B.n772 B.n78 48.746
R1794 B.n612 B.t5 43.0113
R1795 B.n794 B.t12 43.0113
R1796 B.n774 B.n80 36.9956
R1797 B.n769 B.n768 36.9956
R1798 B.n579 B.n578 36.9956
R1799 B.n583 B.n370 36.9956
R1800 B.t2 B.n321 31.5417
R1801 B.t0 B.n36 31.5417
R1802 B.t1 B.n297 30.108
R1803 B.t3 B.n15 30.108
R1804 B.n690 B.t1 18.6385
R1805 B.n844 B.t3 18.6385
R1806 B B.n862 18.0485
R1807 B.n654 B.t2 17.2048
R1808 B.n820 B.t0 17.2048
R1809 B.n129 B.n80 10.6151
R1810 B.n132 B.n129 10.6151
R1811 B.n133 B.n132 10.6151
R1812 B.n136 B.n133 10.6151
R1813 B.n137 B.n136 10.6151
R1814 B.n140 B.n137 10.6151
R1815 B.n141 B.n140 10.6151
R1816 B.n144 B.n141 10.6151
R1817 B.n145 B.n144 10.6151
R1818 B.n148 B.n145 10.6151
R1819 B.n149 B.n148 10.6151
R1820 B.n152 B.n149 10.6151
R1821 B.n153 B.n152 10.6151
R1822 B.n156 B.n153 10.6151
R1823 B.n157 B.n156 10.6151
R1824 B.n160 B.n157 10.6151
R1825 B.n161 B.n160 10.6151
R1826 B.n164 B.n161 10.6151
R1827 B.n165 B.n164 10.6151
R1828 B.n168 B.n165 10.6151
R1829 B.n169 B.n168 10.6151
R1830 B.n172 B.n169 10.6151
R1831 B.n173 B.n172 10.6151
R1832 B.n176 B.n173 10.6151
R1833 B.n177 B.n176 10.6151
R1834 B.n180 B.n177 10.6151
R1835 B.n181 B.n180 10.6151
R1836 B.n184 B.n181 10.6151
R1837 B.n185 B.n184 10.6151
R1838 B.n188 B.n185 10.6151
R1839 B.n189 B.n188 10.6151
R1840 B.n192 B.n189 10.6151
R1841 B.n193 B.n192 10.6151
R1842 B.n196 B.n193 10.6151
R1843 B.n197 B.n196 10.6151
R1844 B.n201 B.n200 10.6151
R1845 B.n204 B.n201 10.6151
R1846 B.n205 B.n204 10.6151
R1847 B.n208 B.n205 10.6151
R1848 B.n209 B.n208 10.6151
R1849 B.n212 B.n209 10.6151
R1850 B.n213 B.n212 10.6151
R1851 B.n216 B.n213 10.6151
R1852 B.n221 B.n218 10.6151
R1853 B.n222 B.n221 10.6151
R1854 B.n225 B.n222 10.6151
R1855 B.n226 B.n225 10.6151
R1856 B.n229 B.n226 10.6151
R1857 B.n230 B.n229 10.6151
R1858 B.n233 B.n230 10.6151
R1859 B.n234 B.n233 10.6151
R1860 B.n237 B.n234 10.6151
R1861 B.n238 B.n237 10.6151
R1862 B.n241 B.n238 10.6151
R1863 B.n242 B.n241 10.6151
R1864 B.n245 B.n242 10.6151
R1865 B.n246 B.n245 10.6151
R1866 B.n249 B.n246 10.6151
R1867 B.n250 B.n249 10.6151
R1868 B.n253 B.n250 10.6151
R1869 B.n254 B.n253 10.6151
R1870 B.n257 B.n254 10.6151
R1871 B.n258 B.n257 10.6151
R1872 B.n261 B.n258 10.6151
R1873 B.n262 B.n261 10.6151
R1874 B.n265 B.n262 10.6151
R1875 B.n266 B.n265 10.6151
R1876 B.n269 B.n266 10.6151
R1877 B.n270 B.n269 10.6151
R1878 B.n273 B.n270 10.6151
R1879 B.n274 B.n273 10.6151
R1880 B.n277 B.n274 10.6151
R1881 B.n278 B.n277 10.6151
R1882 B.n281 B.n278 10.6151
R1883 B.n282 B.n281 10.6151
R1884 B.n285 B.n282 10.6151
R1885 B.n286 B.n285 10.6151
R1886 B.n769 B.n286 10.6151
R1887 B.n579 B.n366 10.6151
R1888 B.n589 B.n366 10.6151
R1889 B.n590 B.n589 10.6151
R1890 B.n591 B.n590 10.6151
R1891 B.n591 B.n358 10.6151
R1892 B.n601 B.n358 10.6151
R1893 B.n602 B.n601 10.6151
R1894 B.n603 B.n602 10.6151
R1895 B.n603 B.n351 10.6151
R1896 B.n614 B.n351 10.6151
R1897 B.n615 B.n614 10.6151
R1898 B.n616 B.n615 10.6151
R1899 B.n616 B.n343 10.6151
R1900 B.n626 B.n343 10.6151
R1901 B.n627 B.n626 10.6151
R1902 B.n628 B.n627 10.6151
R1903 B.n628 B.n335 10.6151
R1904 B.n638 B.n335 10.6151
R1905 B.n639 B.n638 10.6151
R1906 B.n640 B.n639 10.6151
R1907 B.n640 B.n327 10.6151
R1908 B.n650 B.n327 10.6151
R1909 B.n651 B.n650 10.6151
R1910 B.n652 B.n651 10.6151
R1911 B.n652 B.n319 10.6151
R1912 B.n662 B.n319 10.6151
R1913 B.n663 B.n662 10.6151
R1914 B.n664 B.n663 10.6151
R1915 B.n664 B.n311 10.6151
R1916 B.n674 B.n311 10.6151
R1917 B.n675 B.n674 10.6151
R1918 B.n676 B.n675 10.6151
R1919 B.n676 B.n303 10.6151
R1920 B.n686 B.n303 10.6151
R1921 B.n687 B.n686 10.6151
R1922 B.n688 B.n687 10.6151
R1923 B.n688 B.n295 10.6151
R1924 B.n698 B.n295 10.6151
R1925 B.n699 B.n698 10.6151
R1926 B.n701 B.n699 10.6151
R1927 B.n701 B.n700 10.6151
R1928 B.n700 B.n287 10.6151
R1929 B.n712 B.n287 10.6151
R1930 B.n713 B.n712 10.6151
R1931 B.n714 B.n713 10.6151
R1932 B.n715 B.n714 10.6151
R1933 B.n717 B.n715 10.6151
R1934 B.n718 B.n717 10.6151
R1935 B.n719 B.n718 10.6151
R1936 B.n720 B.n719 10.6151
R1937 B.n722 B.n720 10.6151
R1938 B.n723 B.n722 10.6151
R1939 B.n724 B.n723 10.6151
R1940 B.n725 B.n724 10.6151
R1941 B.n727 B.n725 10.6151
R1942 B.n728 B.n727 10.6151
R1943 B.n729 B.n728 10.6151
R1944 B.n730 B.n729 10.6151
R1945 B.n732 B.n730 10.6151
R1946 B.n733 B.n732 10.6151
R1947 B.n734 B.n733 10.6151
R1948 B.n735 B.n734 10.6151
R1949 B.n737 B.n735 10.6151
R1950 B.n738 B.n737 10.6151
R1951 B.n739 B.n738 10.6151
R1952 B.n740 B.n739 10.6151
R1953 B.n742 B.n740 10.6151
R1954 B.n743 B.n742 10.6151
R1955 B.n744 B.n743 10.6151
R1956 B.n745 B.n744 10.6151
R1957 B.n747 B.n745 10.6151
R1958 B.n748 B.n747 10.6151
R1959 B.n749 B.n748 10.6151
R1960 B.n750 B.n749 10.6151
R1961 B.n752 B.n750 10.6151
R1962 B.n753 B.n752 10.6151
R1963 B.n754 B.n753 10.6151
R1964 B.n755 B.n754 10.6151
R1965 B.n757 B.n755 10.6151
R1966 B.n758 B.n757 10.6151
R1967 B.n759 B.n758 10.6151
R1968 B.n760 B.n759 10.6151
R1969 B.n762 B.n760 10.6151
R1970 B.n763 B.n762 10.6151
R1971 B.n764 B.n763 10.6151
R1972 B.n765 B.n764 10.6151
R1973 B.n767 B.n765 10.6151
R1974 B.n768 B.n767 10.6151
R1975 B.n417 B.n370 10.6151
R1976 B.n417 B.n416 10.6151
R1977 B.n423 B.n416 10.6151
R1978 B.n424 B.n423 10.6151
R1979 B.n425 B.n424 10.6151
R1980 B.n425 B.n414 10.6151
R1981 B.n431 B.n414 10.6151
R1982 B.n432 B.n431 10.6151
R1983 B.n433 B.n432 10.6151
R1984 B.n433 B.n412 10.6151
R1985 B.n439 B.n412 10.6151
R1986 B.n440 B.n439 10.6151
R1987 B.n441 B.n440 10.6151
R1988 B.n441 B.n410 10.6151
R1989 B.n447 B.n410 10.6151
R1990 B.n448 B.n447 10.6151
R1991 B.n449 B.n448 10.6151
R1992 B.n449 B.n408 10.6151
R1993 B.n455 B.n408 10.6151
R1994 B.n456 B.n455 10.6151
R1995 B.n457 B.n456 10.6151
R1996 B.n457 B.n406 10.6151
R1997 B.n463 B.n406 10.6151
R1998 B.n464 B.n463 10.6151
R1999 B.n465 B.n464 10.6151
R2000 B.n465 B.n404 10.6151
R2001 B.n471 B.n404 10.6151
R2002 B.n472 B.n471 10.6151
R2003 B.n473 B.n472 10.6151
R2004 B.n473 B.n402 10.6151
R2005 B.n479 B.n402 10.6151
R2006 B.n480 B.n479 10.6151
R2007 B.n481 B.n480 10.6151
R2008 B.n481 B.n400 10.6151
R2009 B.n487 B.n400 10.6151
R2010 B.n490 B.n489 10.6151
R2011 B.n490 B.n396 10.6151
R2012 B.n496 B.n396 10.6151
R2013 B.n497 B.n496 10.6151
R2014 B.n498 B.n497 10.6151
R2015 B.n498 B.n394 10.6151
R2016 B.n504 B.n394 10.6151
R2017 B.n505 B.n504 10.6151
R2018 B.n507 B.n390 10.6151
R2019 B.n513 B.n390 10.6151
R2020 B.n514 B.n513 10.6151
R2021 B.n515 B.n514 10.6151
R2022 B.n515 B.n388 10.6151
R2023 B.n521 B.n388 10.6151
R2024 B.n522 B.n521 10.6151
R2025 B.n523 B.n522 10.6151
R2026 B.n523 B.n386 10.6151
R2027 B.n529 B.n386 10.6151
R2028 B.n530 B.n529 10.6151
R2029 B.n531 B.n530 10.6151
R2030 B.n531 B.n384 10.6151
R2031 B.n537 B.n384 10.6151
R2032 B.n538 B.n537 10.6151
R2033 B.n539 B.n538 10.6151
R2034 B.n539 B.n382 10.6151
R2035 B.n545 B.n382 10.6151
R2036 B.n546 B.n545 10.6151
R2037 B.n547 B.n546 10.6151
R2038 B.n547 B.n380 10.6151
R2039 B.n553 B.n380 10.6151
R2040 B.n554 B.n553 10.6151
R2041 B.n555 B.n554 10.6151
R2042 B.n555 B.n378 10.6151
R2043 B.n561 B.n378 10.6151
R2044 B.n562 B.n561 10.6151
R2045 B.n563 B.n562 10.6151
R2046 B.n563 B.n376 10.6151
R2047 B.n569 B.n376 10.6151
R2048 B.n570 B.n569 10.6151
R2049 B.n571 B.n570 10.6151
R2050 B.n571 B.n374 10.6151
R2051 B.n577 B.n374 10.6151
R2052 B.n578 B.n577 10.6151
R2053 B.n584 B.n583 10.6151
R2054 B.n585 B.n584 10.6151
R2055 B.n585 B.n362 10.6151
R2056 B.n595 B.n362 10.6151
R2057 B.n596 B.n595 10.6151
R2058 B.n597 B.n596 10.6151
R2059 B.n597 B.n354 10.6151
R2060 B.n608 B.n354 10.6151
R2061 B.n609 B.n608 10.6151
R2062 B.n610 B.n609 10.6151
R2063 B.n610 B.n347 10.6151
R2064 B.n620 B.n347 10.6151
R2065 B.n621 B.n620 10.6151
R2066 B.n622 B.n621 10.6151
R2067 B.n622 B.n339 10.6151
R2068 B.n632 B.n339 10.6151
R2069 B.n633 B.n632 10.6151
R2070 B.n634 B.n633 10.6151
R2071 B.n634 B.n331 10.6151
R2072 B.n644 B.n331 10.6151
R2073 B.n645 B.n644 10.6151
R2074 B.n646 B.n645 10.6151
R2075 B.n646 B.n323 10.6151
R2076 B.n656 B.n323 10.6151
R2077 B.n657 B.n656 10.6151
R2078 B.n658 B.n657 10.6151
R2079 B.n658 B.n315 10.6151
R2080 B.n668 B.n315 10.6151
R2081 B.n669 B.n668 10.6151
R2082 B.n670 B.n669 10.6151
R2083 B.n670 B.n307 10.6151
R2084 B.n680 B.n307 10.6151
R2085 B.n681 B.n680 10.6151
R2086 B.n682 B.n681 10.6151
R2087 B.n682 B.n299 10.6151
R2088 B.n692 B.n299 10.6151
R2089 B.n693 B.n692 10.6151
R2090 B.n694 B.n693 10.6151
R2091 B.n694 B.n291 10.6151
R2092 B.n705 B.n291 10.6151
R2093 B.n706 B.n705 10.6151
R2094 B.n707 B.n706 10.6151
R2095 B.n707 B.n0 10.6151
R2096 B.n856 B.n1 10.6151
R2097 B.n856 B.n855 10.6151
R2098 B.n855 B.n854 10.6151
R2099 B.n854 B.n10 10.6151
R2100 B.n848 B.n10 10.6151
R2101 B.n848 B.n847 10.6151
R2102 B.n847 B.n846 10.6151
R2103 B.n846 B.n17 10.6151
R2104 B.n840 B.n17 10.6151
R2105 B.n840 B.n839 10.6151
R2106 B.n839 B.n838 10.6151
R2107 B.n838 B.n24 10.6151
R2108 B.n832 B.n24 10.6151
R2109 B.n832 B.n831 10.6151
R2110 B.n831 B.n830 10.6151
R2111 B.n830 B.n31 10.6151
R2112 B.n824 B.n31 10.6151
R2113 B.n824 B.n823 10.6151
R2114 B.n823 B.n822 10.6151
R2115 B.n822 B.n38 10.6151
R2116 B.n816 B.n38 10.6151
R2117 B.n816 B.n815 10.6151
R2118 B.n815 B.n814 10.6151
R2119 B.n814 B.n45 10.6151
R2120 B.n808 B.n45 10.6151
R2121 B.n808 B.n807 10.6151
R2122 B.n807 B.n806 10.6151
R2123 B.n806 B.n52 10.6151
R2124 B.n800 B.n52 10.6151
R2125 B.n800 B.n799 10.6151
R2126 B.n799 B.n798 10.6151
R2127 B.n798 B.n59 10.6151
R2128 B.n792 B.n59 10.6151
R2129 B.n792 B.n791 10.6151
R2130 B.n791 B.n790 10.6151
R2131 B.n790 B.n65 10.6151
R2132 B.n784 B.n65 10.6151
R2133 B.n784 B.n783 10.6151
R2134 B.n783 B.n782 10.6151
R2135 B.n782 B.n73 10.6151
R2136 B.n776 B.n73 10.6151
R2137 B.n776 B.n775 10.6151
R2138 B.n775 B.n774 10.6151
R2139 B.n200 B.n128 6.5566
R2140 B.n217 B.n216 6.5566
R2141 B.n489 B.n488 6.5566
R2142 B.n506 B.n505 6.5566
R2143 B.n605 B.t5 5.73527
R2144 B.n67 B.t12 5.73527
R2145 B.n197 B.n128 4.05904
R2146 B.n218 B.n217 4.05904
R2147 B.n488 B.n487 4.05904
R2148 B.n507 B.n506 4.05904
R2149 B.n862 B.n0 2.81026
R2150 B.n862 B.n1 2.81026
R2151 VP.n21 VP.n20 161.3
R2152 VP.n19 VP.n1 161.3
R2153 VP.n18 VP.n17 161.3
R2154 VP.n16 VP.n2 161.3
R2155 VP.n15 VP.n14 161.3
R2156 VP.n13 VP.n3 161.3
R2157 VP.n12 VP.n11 161.3
R2158 VP.n10 VP.n4 161.3
R2159 VP.n9 VP.n8 161.3
R2160 VP.n5 VP.t2 98.2303
R2161 VP.n5 VP.t1 96.8902
R2162 VP.n7 VP.n6 87.8654
R2163 VP.n22 VP.n0 87.8654
R2164 VP.n7 VP.t3 64.5449
R2165 VP.n0 VP.t0 64.5449
R2166 VP.n6 VP.n5 50.318
R2167 VP.n14 VP.n13 40.4934
R2168 VP.n14 VP.n2 40.4934
R2169 VP.n8 VP.n4 24.4675
R2170 VP.n12 VP.n4 24.4675
R2171 VP.n13 VP.n12 24.4675
R2172 VP.n18 VP.n2 24.4675
R2173 VP.n19 VP.n18 24.4675
R2174 VP.n20 VP.n19 24.4675
R2175 VP.n8 VP.n7 2.20253
R2176 VP.n20 VP.n0 2.20253
R2177 VP.n9 VP.n6 0.354971
R2178 VP.n22 VP.n21 0.354971
R2179 VP VP.n22 0.26696
R2180 VP.n10 VP.n9 0.189894
R2181 VP.n11 VP.n10 0.189894
R2182 VP.n11 VP.n3 0.189894
R2183 VP.n15 VP.n3 0.189894
R2184 VP.n16 VP.n15 0.189894
R2185 VP.n17 VP.n16 0.189894
R2186 VP.n17 VP.n1 0.189894
R2187 VP.n21 VP.n1 0.189894
R2188 VDD1 VDD1.n1 108.272
R2189 VDD1 VDD1.n0 64.8317
R2190 VDD1.n0 VDD1.t1 1.96674
R2191 VDD1.n0 VDD1.t2 1.96674
R2192 VDD1.n1 VDD1.t0 1.96674
R2193 VDD1.n1 VDD1.t3 1.96674
C0 VTAIL VN 4.44444f
C1 VP VDD2 0.467972f
C2 VDD2 VN 4.27415f
C3 VTAIL VDD2 5.39223f
C4 VP VDD1 4.59119f
C5 VDD1 VN 0.149902f
C6 VTAIL VDD1 5.33025f
C7 VDD1 VDD2 1.30724f
C8 VP VN 6.67137f
C9 VP VTAIL 4.45855f
C10 VDD2 B 4.275334f
C11 VDD1 B 8.68393f
C12 VTAIL B 9.537073f
C13 VN B 12.82328f
C14 VP B 11.276844f
C15 VDD1.t1 B 0.222257f
C16 VDD1.t2 B 0.222257f
C17 VDD1.n0 B 1.96045f
C18 VDD1.t0 B 0.222257f
C19 VDD1.t3 B 0.222257f
C20 VDD1.n1 B 2.6582f
C21 VP.t0 B 2.1877f
C22 VP.n0 B 0.852292f
C23 VP.n1 B 0.021323f
C24 VP.n2 B 0.042379f
C25 VP.n3 B 0.021323f
C26 VP.n4 B 0.039741f
C27 VP.t2 B 2.51308f
C28 VP.t1 B 2.5007f
C29 VP.n5 B 2.83231f
C30 VP.n6 B 1.24292f
C31 VP.t3 B 2.1877f
C32 VP.n7 B 0.852292f
C33 VP.n8 B 0.021885f
C34 VP.n9 B 0.034415f
C35 VP.n10 B 0.021323f
C36 VP.n11 B 0.021323f
C37 VP.n12 B 0.039741f
C38 VP.n13 B 0.042379f
C39 VP.n14 B 0.017238f
C40 VP.n15 B 0.021323f
C41 VP.n16 B 0.021323f
C42 VP.n17 B 0.021323f
C43 VP.n18 B 0.039741f
C44 VP.n19 B 0.039741f
C45 VP.n20 B 0.021885f
C46 VP.n21 B 0.034415f
C47 VP.n22 B 0.065448f
C48 VTAIL.n0 B 0.024983f
C49 VTAIL.n1 B 0.017859f
C50 VTAIL.n2 B 0.009597f
C51 VTAIL.n3 B 0.022684f
C52 VTAIL.n4 B 0.010161f
C53 VTAIL.n5 B 0.017859f
C54 VTAIL.n6 B 0.009879f
C55 VTAIL.n7 B 0.022684f
C56 VTAIL.n8 B 0.010161f
C57 VTAIL.n9 B 0.017859f
C58 VTAIL.n10 B 0.009597f
C59 VTAIL.n11 B 0.022684f
C60 VTAIL.n12 B 0.010161f
C61 VTAIL.n13 B 0.017859f
C62 VTAIL.n14 B 0.009597f
C63 VTAIL.n15 B 0.017013f
C64 VTAIL.n16 B 0.016036f
C65 VTAIL.t3 B 0.038127f
C66 VTAIL.n17 B 0.115534f
C67 VTAIL.n18 B 0.747661f
C68 VTAIL.n19 B 0.009597f
C69 VTAIL.n20 B 0.010161f
C70 VTAIL.n21 B 0.022684f
C71 VTAIL.n22 B 0.022684f
C72 VTAIL.n23 B 0.010161f
C73 VTAIL.n24 B 0.009597f
C74 VTAIL.n25 B 0.017859f
C75 VTAIL.n26 B 0.017859f
C76 VTAIL.n27 B 0.009597f
C77 VTAIL.n28 B 0.010161f
C78 VTAIL.n29 B 0.022684f
C79 VTAIL.n30 B 0.022684f
C80 VTAIL.n31 B 0.010161f
C81 VTAIL.n32 B 0.009597f
C82 VTAIL.n33 B 0.017859f
C83 VTAIL.n34 B 0.017859f
C84 VTAIL.n35 B 0.009597f
C85 VTAIL.n36 B 0.009597f
C86 VTAIL.n37 B 0.010161f
C87 VTAIL.n38 B 0.022684f
C88 VTAIL.n39 B 0.022684f
C89 VTAIL.n40 B 0.022684f
C90 VTAIL.n41 B 0.009879f
C91 VTAIL.n42 B 0.009597f
C92 VTAIL.n43 B 0.017859f
C93 VTAIL.n44 B 0.017859f
C94 VTAIL.n45 B 0.009597f
C95 VTAIL.n46 B 0.010161f
C96 VTAIL.n47 B 0.022684f
C97 VTAIL.n48 B 0.048893f
C98 VTAIL.n49 B 0.010161f
C99 VTAIL.n50 B 0.009597f
C100 VTAIL.n51 B 0.043965f
C101 VTAIL.n52 B 0.027416f
C102 VTAIL.n53 B 0.148608f
C103 VTAIL.n54 B 0.024983f
C104 VTAIL.n55 B 0.017859f
C105 VTAIL.n56 B 0.009597f
C106 VTAIL.n57 B 0.022684f
C107 VTAIL.n58 B 0.010161f
C108 VTAIL.n59 B 0.017859f
C109 VTAIL.n60 B 0.009879f
C110 VTAIL.n61 B 0.022684f
C111 VTAIL.n62 B 0.010161f
C112 VTAIL.n63 B 0.017859f
C113 VTAIL.n64 B 0.009597f
C114 VTAIL.n65 B 0.022684f
C115 VTAIL.n66 B 0.010161f
C116 VTAIL.n67 B 0.017859f
C117 VTAIL.n68 B 0.009597f
C118 VTAIL.n69 B 0.017013f
C119 VTAIL.n70 B 0.016036f
C120 VTAIL.t7 B 0.038127f
C121 VTAIL.n71 B 0.115534f
C122 VTAIL.n72 B 0.747661f
C123 VTAIL.n73 B 0.009597f
C124 VTAIL.n74 B 0.010161f
C125 VTAIL.n75 B 0.022684f
C126 VTAIL.n76 B 0.022684f
C127 VTAIL.n77 B 0.010161f
C128 VTAIL.n78 B 0.009597f
C129 VTAIL.n79 B 0.017859f
C130 VTAIL.n80 B 0.017859f
C131 VTAIL.n81 B 0.009597f
C132 VTAIL.n82 B 0.010161f
C133 VTAIL.n83 B 0.022684f
C134 VTAIL.n84 B 0.022684f
C135 VTAIL.n85 B 0.010161f
C136 VTAIL.n86 B 0.009597f
C137 VTAIL.n87 B 0.017859f
C138 VTAIL.n88 B 0.017859f
C139 VTAIL.n89 B 0.009597f
C140 VTAIL.n90 B 0.009597f
C141 VTAIL.n91 B 0.010161f
C142 VTAIL.n92 B 0.022684f
C143 VTAIL.n93 B 0.022684f
C144 VTAIL.n94 B 0.022684f
C145 VTAIL.n95 B 0.009879f
C146 VTAIL.n96 B 0.009597f
C147 VTAIL.n97 B 0.017859f
C148 VTAIL.n98 B 0.017859f
C149 VTAIL.n99 B 0.009597f
C150 VTAIL.n100 B 0.010161f
C151 VTAIL.n101 B 0.022684f
C152 VTAIL.n102 B 0.048893f
C153 VTAIL.n103 B 0.010161f
C154 VTAIL.n104 B 0.009597f
C155 VTAIL.n105 B 0.043965f
C156 VTAIL.n106 B 0.027416f
C157 VTAIL.n107 B 0.24671f
C158 VTAIL.n108 B 0.024983f
C159 VTAIL.n109 B 0.017859f
C160 VTAIL.n110 B 0.009597f
C161 VTAIL.n111 B 0.022684f
C162 VTAIL.n112 B 0.010161f
C163 VTAIL.n113 B 0.017859f
C164 VTAIL.n114 B 0.009879f
C165 VTAIL.n115 B 0.022684f
C166 VTAIL.n116 B 0.010161f
C167 VTAIL.n117 B 0.017859f
C168 VTAIL.n118 B 0.009597f
C169 VTAIL.n119 B 0.022684f
C170 VTAIL.n120 B 0.010161f
C171 VTAIL.n121 B 0.017859f
C172 VTAIL.n122 B 0.009597f
C173 VTAIL.n123 B 0.017013f
C174 VTAIL.n124 B 0.016036f
C175 VTAIL.t5 B 0.038127f
C176 VTAIL.n125 B 0.115534f
C177 VTAIL.n126 B 0.747661f
C178 VTAIL.n127 B 0.009597f
C179 VTAIL.n128 B 0.010161f
C180 VTAIL.n129 B 0.022684f
C181 VTAIL.n130 B 0.022684f
C182 VTAIL.n131 B 0.010161f
C183 VTAIL.n132 B 0.009597f
C184 VTAIL.n133 B 0.017859f
C185 VTAIL.n134 B 0.017859f
C186 VTAIL.n135 B 0.009597f
C187 VTAIL.n136 B 0.010161f
C188 VTAIL.n137 B 0.022684f
C189 VTAIL.n138 B 0.022684f
C190 VTAIL.n139 B 0.010161f
C191 VTAIL.n140 B 0.009597f
C192 VTAIL.n141 B 0.017859f
C193 VTAIL.n142 B 0.017859f
C194 VTAIL.n143 B 0.009597f
C195 VTAIL.n144 B 0.009597f
C196 VTAIL.n145 B 0.010161f
C197 VTAIL.n146 B 0.022684f
C198 VTAIL.n147 B 0.022684f
C199 VTAIL.n148 B 0.022684f
C200 VTAIL.n149 B 0.009879f
C201 VTAIL.n150 B 0.009597f
C202 VTAIL.n151 B 0.017859f
C203 VTAIL.n152 B 0.017859f
C204 VTAIL.n153 B 0.009597f
C205 VTAIL.n154 B 0.010161f
C206 VTAIL.n155 B 0.022684f
C207 VTAIL.n156 B 0.048893f
C208 VTAIL.n157 B 0.010161f
C209 VTAIL.n158 B 0.009597f
C210 VTAIL.n159 B 0.043965f
C211 VTAIL.n160 B 0.027416f
C212 VTAIL.n161 B 1.16474f
C213 VTAIL.n162 B 0.024983f
C214 VTAIL.n163 B 0.017859f
C215 VTAIL.n164 B 0.009597f
C216 VTAIL.n165 B 0.022684f
C217 VTAIL.n166 B 0.010161f
C218 VTAIL.n167 B 0.017859f
C219 VTAIL.n168 B 0.009879f
C220 VTAIL.n169 B 0.022684f
C221 VTAIL.n170 B 0.009597f
C222 VTAIL.n171 B 0.010161f
C223 VTAIL.n172 B 0.017859f
C224 VTAIL.n173 B 0.009597f
C225 VTAIL.n174 B 0.022684f
C226 VTAIL.n175 B 0.010161f
C227 VTAIL.n176 B 0.017859f
C228 VTAIL.n177 B 0.009597f
C229 VTAIL.n178 B 0.017013f
C230 VTAIL.n179 B 0.016036f
C231 VTAIL.t2 B 0.038127f
C232 VTAIL.n180 B 0.115534f
C233 VTAIL.n181 B 0.747661f
C234 VTAIL.n182 B 0.009597f
C235 VTAIL.n183 B 0.010161f
C236 VTAIL.n184 B 0.022684f
C237 VTAIL.n185 B 0.022684f
C238 VTAIL.n186 B 0.010161f
C239 VTAIL.n187 B 0.009597f
C240 VTAIL.n188 B 0.017859f
C241 VTAIL.n189 B 0.017859f
C242 VTAIL.n190 B 0.009597f
C243 VTAIL.n191 B 0.010161f
C244 VTAIL.n192 B 0.022684f
C245 VTAIL.n193 B 0.022684f
C246 VTAIL.n194 B 0.010161f
C247 VTAIL.n195 B 0.009597f
C248 VTAIL.n196 B 0.017859f
C249 VTAIL.n197 B 0.017859f
C250 VTAIL.n198 B 0.009597f
C251 VTAIL.n199 B 0.010161f
C252 VTAIL.n200 B 0.022684f
C253 VTAIL.n201 B 0.022684f
C254 VTAIL.n202 B 0.022684f
C255 VTAIL.n203 B 0.009879f
C256 VTAIL.n204 B 0.009597f
C257 VTAIL.n205 B 0.017859f
C258 VTAIL.n206 B 0.017859f
C259 VTAIL.n207 B 0.009597f
C260 VTAIL.n208 B 0.010161f
C261 VTAIL.n209 B 0.022684f
C262 VTAIL.n210 B 0.048893f
C263 VTAIL.n211 B 0.010161f
C264 VTAIL.n212 B 0.009597f
C265 VTAIL.n213 B 0.043965f
C266 VTAIL.n214 B 0.027416f
C267 VTAIL.n215 B 1.16474f
C268 VTAIL.n216 B 0.024983f
C269 VTAIL.n217 B 0.017859f
C270 VTAIL.n218 B 0.009597f
C271 VTAIL.n219 B 0.022684f
C272 VTAIL.n220 B 0.010161f
C273 VTAIL.n221 B 0.017859f
C274 VTAIL.n222 B 0.009879f
C275 VTAIL.n223 B 0.022684f
C276 VTAIL.n224 B 0.009597f
C277 VTAIL.n225 B 0.010161f
C278 VTAIL.n226 B 0.017859f
C279 VTAIL.n227 B 0.009597f
C280 VTAIL.n228 B 0.022684f
C281 VTAIL.n229 B 0.010161f
C282 VTAIL.n230 B 0.017859f
C283 VTAIL.n231 B 0.009597f
C284 VTAIL.n232 B 0.017013f
C285 VTAIL.n233 B 0.016036f
C286 VTAIL.t1 B 0.038127f
C287 VTAIL.n234 B 0.115534f
C288 VTAIL.n235 B 0.747661f
C289 VTAIL.n236 B 0.009597f
C290 VTAIL.n237 B 0.010161f
C291 VTAIL.n238 B 0.022684f
C292 VTAIL.n239 B 0.022684f
C293 VTAIL.n240 B 0.010161f
C294 VTAIL.n241 B 0.009597f
C295 VTAIL.n242 B 0.017859f
C296 VTAIL.n243 B 0.017859f
C297 VTAIL.n244 B 0.009597f
C298 VTAIL.n245 B 0.010161f
C299 VTAIL.n246 B 0.022684f
C300 VTAIL.n247 B 0.022684f
C301 VTAIL.n248 B 0.010161f
C302 VTAIL.n249 B 0.009597f
C303 VTAIL.n250 B 0.017859f
C304 VTAIL.n251 B 0.017859f
C305 VTAIL.n252 B 0.009597f
C306 VTAIL.n253 B 0.010161f
C307 VTAIL.n254 B 0.022684f
C308 VTAIL.n255 B 0.022684f
C309 VTAIL.n256 B 0.022684f
C310 VTAIL.n257 B 0.009879f
C311 VTAIL.n258 B 0.009597f
C312 VTAIL.n259 B 0.017859f
C313 VTAIL.n260 B 0.017859f
C314 VTAIL.n261 B 0.009597f
C315 VTAIL.n262 B 0.010161f
C316 VTAIL.n263 B 0.022684f
C317 VTAIL.n264 B 0.048893f
C318 VTAIL.n265 B 0.010161f
C319 VTAIL.n266 B 0.009597f
C320 VTAIL.n267 B 0.043965f
C321 VTAIL.n268 B 0.027416f
C322 VTAIL.n269 B 0.24671f
C323 VTAIL.n270 B 0.024983f
C324 VTAIL.n271 B 0.017859f
C325 VTAIL.n272 B 0.009597f
C326 VTAIL.n273 B 0.022684f
C327 VTAIL.n274 B 0.010161f
C328 VTAIL.n275 B 0.017859f
C329 VTAIL.n276 B 0.009879f
C330 VTAIL.n277 B 0.022684f
C331 VTAIL.n278 B 0.009597f
C332 VTAIL.n279 B 0.010161f
C333 VTAIL.n280 B 0.017859f
C334 VTAIL.n281 B 0.009597f
C335 VTAIL.n282 B 0.022684f
C336 VTAIL.n283 B 0.010161f
C337 VTAIL.n284 B 0.017859f
C338 VTAIL.n285 B 0.009597f
C339 VTAIL.n286 B 0.017013f
C340 VTAIL.n287 B 0.016036f
C341 VTAIL.t4 B 0.038127f
C342 VTAIL.n288 B 0.115534f
C343 VTAIL.n289 B 0.747661f
C344 VTAIL.n290 B 0.009597f
C345 VTAIL.n291 B 0.010161f
C346 VTAIL.n292 B 0.022684f
C347 VTAIL.n293 B 0.022684f
C348 VTAIL.n294 B 0.010161f
C349 VTAIL.n295 B 0.009597f
C350 VTAIL.n296 B 0.017859f
C351 VTAIL.n297 B 0.017859f
C352 VTAIL.n298 B 0.009597f
C353 VTAIL.n299 B 0.010161f
C354 VTAIL.n300 B 0.022684f
C355 VTAIL.n301 B 0.022684f
C356 VTAIL.n302 B 0.010161f
C357 VTAIL.n303 B 0.009597f
C358 VTAIL.n304 B 0.017859f
C359 VTAIL.n305 B 0.017859f
C360 VTAIL.n306 B 0.009597f
C361 VTAIL.n307 B 0.010161f
C362 VTAIL.n308 B 0.022684f
C363 VTAIL.n309 B 0.022684f
C364 VTAIL.n310 B 0.022684f
C365 VTAIL.n311 B 0.009879f
C366 VTAIL.n312 B 0.009597f
C367 VTAIL.n313 B 0.017859f
C368 VTAIL.n314 B 0.017859f
C369 VTAIL.n315 B 0.009597f
C370 VTAIL.n316 B 0.010161f
C371 VTAIL.n317 B 0.022684f
C372 VTAIL.n318 B 0.048893f
C373 VTAIL.n319 B 0.010161f
C374 VTAIL.n320 B 0.009597f
C375 VTAIL.n321 B 0.043965f
C376 VTAIL.n322 B 0.027416f
C377 VTAIL.n323 B 0.24671f
C378 VTAIL.n324 B 0.024983f
C379 VTAIL.n325 B 0.017859f
C380 VTAIL.n326 B 0.009597f
C381 VTAIL.n327 B 0.022684f
C382 VTAIL.n328 B 0.010161f
C383 VTAIL.n329 B 0.017859f
C384 VTAIL.n330 B 0.009879f
C385 VTAIL.n331 B 0.022684f
C386 VTAIL.n332 B 0.009597f
C387 VTAIL.n333 B 0.010161f
C388 VTAIL.n334 B 0.017859f
C389 VTAIL.n335 B 0.009597f
C390 VTAIL.n336 B 0.022684f
C391 VTAIL.n337 B 0.010161f
C392 VTAIL.n338 B 0.017859f
C393 VTAIL.n339 B 0.009597f
C394 VTAIL.n340 B 0.017013f
C395 VTAIL.n341 B 0.016036f
C396 VTAIL.t6 B 0.038127f
C397 VTAIL.n342 B 0.115534f
C398 VTAIL.n343 B 0.747661f
C399 VTAIL.n344 B 0.009597f
C400 VTAIL.n345 B 0.010161f
C401 VTAIL.n346 B 0.022684f
C402 VTAIL.n347 B 0.022684f
C403 VTAIL.n348 B 0.010161f
C404 VTAIL.n349 B 0.009597f
C405 VTAIL.n350 B 0.017859f
C406 VTAIL.n351 B 0.017859f
C407 VTAIL.n352 B 0.009597f
C408 VTAIL.n353 B 0.010161f
C409 VTAIL.n354 B 0.022684f
C410 VTAIL.n355 B 0.022684f
C411 VTAIL.n356 B 0.010161f
C412 VTAIL.n357 B 0.009597f
C413 VTAIL.n358 B 0.017859f
C414 VTAIL.n359 B 0.017859f
C415 VTAIL.n360 B 0.009597f
C416 VTAIL.n361 B 0.010161f
C417 VTAIL.n362 B 0.022684f
C418 VTAIL.n363 B 0.022684f
C419 VTAIL.n364 B 0.022684f
C420 VTAIL.n365 B 0.009879f
C421 VTAIL.n366 B 0.009597f
C422 VTAIL.n367 B 0.017859f
C423 VTAIL.n368 B 0.017859f
C424 VTAIL.n369 B 0.009597f
C425 VTAIL.n370 B 0.010161f
C426 VTAIL.n371 B 0.022684f
C427 VTAIL.n372 B 0.048893f
C428 VTAIL.n373 B 0.010161f
C429 VTAIL.n374 B 0.009597f
C430 VTAIL.n375 B 0.043965f
C431 VTAIL.n376 B 0.027416f
C432 VTAIL.n377 B 1.16474f
C433 VTAIL.n378 B 0.024983f
C434 VTAIL.n379 B 0.017859f
C435 VTAIL.n380 B 0.009597f
C436 VTAIL.n381 B 0.022684f
C437 VTAIL.n382 B 0.010161f
C438 VTAIL.n383 B 0.017859f
C439 VTAIL.n384 B 0.009879f
C440 VTAIL.n385 B 0.022684f
C441 VTAIL.n386 B 0.010161f
C442 VTAIL.n387 B 0.017859f
C443 VTAIL.n388 B 0.009597f
C444 VTAIL.n389 B 0.022684f
C445 VTAIL.n390 B 0.010161f
C446 VTAIL.n391 B 0.017859f
C447 VTAIL.n392 B 0.009597f
C448 VTAIL.n393 B 0.017013f
C449 VTAIL.n394 B 0.016036f
C450 VTAIL.t0 B 0.038127f
C451 VTAIL.n395 B 0.115534f
C452 VTAIL.n396 B 0.747661f
C453 VTAIL.n397 B 0.009597f
C454 VTAIL.n398 B 0.010161f
C455 VTAIL.n399 B 0.022684f
C456 VTAIL.n400 B 0.022684f
C457 VTAIL.n401 B 0.010161f
C458 VTAIL.n402 B 0.009597f
C459 VTAIL.n403 B 0.017859f
C460 VTAIL.n404 B 0.017859f
C461 VTAIL.n405 B 0.009597f
C462 VTAIL.n406 B 0.010161f
C463 VTAIL.n407 B 0.022684f
C464 VTAIL.n408 B 0.022684f
C465 VTAIL.n409 B 0.010161f
C466 VTAIL.n410 B 0.009597f
C467 VTAIL.n411 B 0.017859f
C468 VTAIL.n412 B 0.017859f
C469 VTAIL.n413 B 0.009597f
C470 VTAIL.n414 B 0.009597f
C471 VTAIL.n415 B 0.010161f
C472 VTAIL.n416 B 0.022684f
C473 VTAIL.n417 B 0.022684f
C474 VTAIL.n418 B 0.022684f
C475 VTAIL.n419 B 0.009879f
C476 VTAIL.n420 B 0.009597f
C477 VTAIL.n421 B 0.017859f
C478 VTAIL.n422 B 0.017859f
C479 VTAIL.n423 B 0.009597f
C480 VTAIL.n424 B 0.010161f
C481 VTAIL.n425 B 0.022684f
C482 VTAIL.n426 B 0.048893f
C483 VTAIL.n427 B 0.010161f
C484 VTAIL.n428 B 0.009597f
C485 VTAIL.n429 B 0.043965f
C486 VTAIL.n430 B 0.027416f
C487 VTAIL.n431 B 1.05994f
C488 VDD2.t0 B 0.22006f
C489 VDD2.t2 B 0.22006f
C490 VDD2.n0 B 2.60511f
C491 VDD2.t1 B 0.22006f
C492 VDD2.t3 B 0.22006f
C493 VDD2.n1 B 1.94057f
C494 VDD2.n2 B 3.95394f
C495 VN.t3 B 2.43277f
C496 VN.t0 B 2.44482f
C497 VN.n0 B 1.45322f
C498 VN.t1 B 2.43277f
C499 VN.t2 B 2.44482f
C500 VN.n1 B 2.76381f
.ends

