* NGSPICE file created from diff_pair_sample_0934.ext - technology: sky130A

.subckt diff_pair_sample_0934 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t2 w_n1290_n3148# sky130_fd_pr__pfet_01v8 ad=4.2432 pd=22.54 as=4.2432 ps=22.54 w=10.88 l=0.47
X1 B.t11 B.t9 B.t10 w_n1290_n3148# sky130_fd_pr__pfet_01v8 ad=4.2432 pd=22.54 as=0 ps=0 w=10.88 l=0.47
X2 VDD1.t1 VP.t0 VTAIL.t1 w_n1290_n3148# sky130_fd_pr__pfet_01v8 ad=4.2432 pd=22.54 as=4.2432 ps=22.54 w=10.88 l=0.47
X3 B.t8 B.t6 B.t7 w_n1290_n3148# sky130_fd_pr__pfet_01v8 ad=4.2432 pd=22.54 as=0 ps=0 w=10.88 l=0.47
X4 B.t5 B.t3 B.t4 w_n1290_n3148# sky130_fd_pr__pfet_01v8 ad=4.2432 pd=22.54 as=0 ps=0 w=10.88 l=0.47
X5 VDD2.t0 VN.t1 VTAIL.t3 w_n1290_n3148# sky130_fd_pr__pfet_01v8 ad=4.2432 pd=22.54 as=4.2432 ps=22.54 w=10.88 l=0.47
X6 B.t2 B.t0 B.t1 w_n1290_n3148# sky130_fd_pr__pfet_01v8 ad=4.2432 pd=22.54 as=0 ps=0 w=10.88 l=0.47
X7 VDD1.t0 VP.t1 VTAIL.t0 w_n1290_n3148# sky130_fd_pr__pfet_01v8 ad=4.2432 pd=22.54 as=4.2432 ps=22.54 w=10.88 l=0.47
R0 VN VN.t1 842.351
R1 VN VN.t0 803.847
R2 VTAIL.n1 VTAIL.t3 64.953
R3 VTAIL.n3 VTAIL.t2 64.952
R4 VTAIL.n0 VTAIL.t0 64.952
R5 VTAIL.n2 VTAIL.t1 64.9518
R6 VTAIL.n1 VTAIL.n0 23.1427
R7 VTAIL.n3 VTAIL.n2 22.4531
R8 VTAIL.n2 VTAIL.n1 0.815155
R9 VTAIL VTAIL.n0 0.700931
R10 VTAIL VTAIL.n3 0.114724
R11 VDD2.n0 VDD2.t1 116.067
R12 VDD2.n0 VDD2.t0 81.6306
R13 VDD2 VDD2.n0 0.231103
R14 B.n89 B.t6 765.067
R15 B.n97 B.t3 765.067
R16 B.n28 B.t9 765.067
R17 B.n36 B.t0 765.067
R18 B.n313 B.n56 585
R19 B.n315 B.n314 585
R20 B.n316 B.n55 585
R21 B.n318 B.n317 585
R22 B.n319 B.n54 585
R23 B.n321 B.n320 585
R24 B.n322 B.n53 585
R25 B.n324 B.n323 585
R26 B.n325 B.n52 585
R27 B.n327 B.n326 585
R28 B.n328 B.n51 585
R29 B.n330 B.n329 585
R30 B.n331 B.n50 585
R31 B.n333 B.n332 585
R32 B.n334 B.n49 585
R33 B.n336 B.n335 585
R34 B.n337 B.n48 585
R35 B.n339 B.n338 585
R36 B.n340 B.n47 585
R37 B.n342 B.n341 585
R38 B.n343 B.n46 585
R39 B.n345 B.n344 585
R40 B.n346 B.n45 585
R41 B.n348 B.n347 585
R42 B.n349 B.n44 585
R43 B.n351 B.n350 585
R44 B.n352 B.n43 585
R45 B.n354 B.n353 585
R46 B.n355 B.n42 585
R47 B.n357 B.n356 585
R48 B.n358 B.n41 585
R49 B.n360 B.n359 585
R50 B.n361 B.n40 585
R51 B.n363 B.n362 585
R52 B.n364 B.n39 585
R53 B.n366 B.n365 585
R54 B.n367 B.n35 585
R55 B.n369 B.n368 585
R56 B.n370 B.n34 585
R57 B.n372 B.n371 585
R58 B.n373 B.n33 585
R59 B.n375 B.n374 585
R60 B.n376 B.n32 585
R61 B.n378 B.n377 585
R62 B.n379 B.n31 585
R63 B.n381 B.n380 585
R64 B.n382 B.n30 585
R65 B.n384 B.n383 585
R66 B.n386 B.n27 585
R67 B.n388 B.n387 585
R68 B.n389 B.n26 585
R69 B.n391 B.n390 585
R70 B.n392 B.n25 585
R71 B.n394 B.n393 585
R72 B.n395 B.n24 585
R73 B.n397 B.n396 585
R74 B.n398 B.n23 585
R75 B.n400 B.n399 585
R76 B.n401 B.n22 585
R77 B.n403 B.n402 585
R78 B.n404 B.n21 585
R79 B.n406 B.n405 585
R80 B.n407 B.n20 585
R81 B.n409 B.n408 585
R82 B.n410 B.n19 585
R83 B.n412 B.n411 585
R84 B.n413 B.n18 585
R85 B.n415 B.n414 585
R86 B.n416 B.n17 585
R87 B.n418 B.n417 585
R88 B.n419 B.n16 585
R89 B.n421 B.n420 585
R90 B.n422 B.n15 585
R91 B.n424 B.n423 585
R92 B.n425 B.n14 585
R93 B.n427 B.n426 585
R94 B.n428 B.n13 585
R95 B.n430 B.n429 585
R96 B.n431 B.n12 585
R97 B.n433 B.n432 585
R98 B.n434 B.n11 585
R99 B.n436 B.n435 585
R100 B.n437 B.n10 585
R101 B.n439 B.n438 585
R102 B.n440 B.n9 585
R103 B.n442 B.n441 585
R104 B.n312 B.n311 585
R105 B.n310 B.n57 585
R106 B.n309 B.n308 585
R107 B.n307 B.n58 585
R108 B.n306 B.n305 585
R109 B.n304 B.n59 585
R110 B.n303 B.n302 585
R111 B.n301 B.n60 585
R112 B.n300 B.n299 585
R113 B.n298 B.n61 585
R114 B.n297 B.n296 585
R115 B.n295 B.n62 585
R116 B.n294 B.n293 585
R117 B.n292 B.n63 585
R118 B.n291 B.n290 585
R119 B.n289 B.n64 585
R120 B.n288 B.n287 585
R121 B.n286 B.n65 585
R122 B.n285 B.n284 585
R123 B.n283 B.n66 585
R124 B.n282 B.n281 585
R125 B.n280 B.n67 585
R126 B.n279 B.n278 585
R127 B.n277 B.n68 585
R128 B.n276 B.n275 585
R129 B.n274 B.n69 585
R130 B.n273 B.n272 585
R131 B.n142 B.n117 585
R132 B.n144 B.n143 585
R133 B.n145 B.n116 585
R134 B.n147 B.n146 585
R135 B.n148 B.n115 585
R136 B.n150 B.n149 585
R137 B.n151 B.n114 585
R138 B.n153 B.n152 585
R139 B.n154 B.n113 585
R140 B.n156 B.n155 585
R141 B.n157 B.n112 585
R142 B.n159 B.n158 585
R143 B.n160 B.n111 585
R144 B.n162 B.n161 585
R145 B.n163 B.n110 585
R146 B.n165 B.n164 585
R147 B.n166 B.n109 585
R148 B.n168 B.n167 585
R149 B.n169 B.n108 585
R150 B.n171 B.n170 585
R151 B.n172 B.n107 585
R152 B.n174 B.n173 585
R153 B.n175 B.n106 585
R154 B.n177 B.n176 585
R155 B.n178 B.n105 585
R156 B.n180 B.n179 585
R157 B.n181 B.n104 585
R158 B.n183 B.n182 585
R159 B.n184 B.n103 585
R160 B.n186 B.n185 585
R161 B.n187 B.n102 585
R162 B.n189 B.n188 585
R163 B.n190 B.n101 585
R164 B.n192 B.n191 585
R165 B.n193 B.n100 585
R166 B.n195 B.n194 585
R167 B.n196 B.n99 585
R168 B.n198 B.n197 585
R169 B.n200 B.n96 585
R170 B.n202 B.n201 585
R171 B.n203 B.n95 585
R172 B.n205 B.n204 585
R173 B.n206 B.n94 585
R174 B.n208 B.n207 585
R175 B.n209 B.n93 585
R176 B.n211 B.n210 585
R177 B.n212 B.n92 585
R178 B.n214 B.n213 585
R179 B.n216 B.n215 585
R180 B.n217 B.n88 585
R181 B.n219 B.n218 585
R182 B.n220 B.n87 585
R183 B.n222 B.n221 585
R184 B.n223 B.n86 585
R185 B.n225 B.n224 585
R186 B.n226 B.n85 585
R187 B.n228 B.n227 585
R188 B.n229 B.n84 585
R189 B.n231 B.n230 585
R190 B.n232 B.n83 585
R191 B.n234 B.n233 585
R192 B.n235 B.n82 585
R193 B.n237 B.n236 585
R194 B.n238 B.n81 585
R195 B.n240 B.n239 585
R196 B.n241 B.n80 585
R197 B.n243 B.n242 585
R198 B.n244 B.n79 585
R199 B.n246 B.n245 585
R200 B.n247 B.n78 585
R201 B.n249 B.n248 585
R202 B.n250 B.n77 585
R203 B.n252 B.n251 585
R204 B.n253 B.n76 585
R205 B.n255 B.n254 585
R206 B.n256 B.n75 585
R207 B.n258 B.n257 585
R208 B.n259 B.n74 585
R209 B.n261 B.n260 585
R210 B.n262 B.n73 585
R211 B.n264 B.n263 585
R212 B.n265 B.n72 585
R213 B.n267 B.n266 585
R214 B.n268 B.n71 585
R215 B.n270 B.n269 585
R216 B.n271 B.n70 585
R217 B.n141 B.n140 585
R218 B.n139 B.n118 585
R219 B.n138 B.n137 585
R220 B.n136 B.n119 585
R221 B.n135 B.n134 585
R222 B.n133 B.n120 585
R223 B.n132 B.n131 585
R224 B.n130 B.n121 585
R225 B.n129 B.n128 585
R226 B.n127 B.n122 585
R227 B.n126 B.n125 585
R228 B.n124 B.n123 585
R229 B.n2 B.n0 585
R230 B.n461 B.n1 585
R231 B.n460 B.n459 585
R232 B.n458 B.n3 585
R233 B.n457 B.n456 585
R234 B.n455 B.n4 585
R235 B.n454 B.n453 585
R236 B.n452 B.n5 585
R237 B.n451 B.n450 585
R238 B.n449 B.n6 585
R239 B.n448 B.n447 585
R240 B.n446 B.n7 585
R241 B.n445 B.n444 585
R242 B.n443 B.n8 585
R243 B.n463 B.n462 585
R244 B.n142 B.n141 497.305
R245 B.n443 B.n442 497.305
R246 B.n273 B.n70 497.305
R247 B.n311 B.n56 497.305
R248 B.n141 B.n118 163.367
R249 B.n137 B.n118 163.367
R250 B.n137 B.n136 163.367
R251 B.n136 B.n135 163.367
R252 B.n135 B.n120 163.367
R253 B.n131 B.n120 163.367
R254 B.n131 B.n130 163.367
R255 B.n130 B.n129 163.367
R256 B.n129 B.n122 163.367
R257 B.n125 B.n122 163.367
R258 B.n125 B.n124 163.367
R259 B.n124 B.n2 163.367
R260 B.n462 B.n2 163.367
R261 B.n462 B.n461 163.367
R262 B.n461 B.n460 163.367
R263 B.n460 B.n3 163.367
R264 B.n456 B.n3 163.367
R265 B.n456 B.n455 163.367
R266 B.n455 B.n454 163.367
R267 B.n454 B.n5 163.367
R268 B.n450 B.n5 163.367
R269 B.n450 B.n449 163.367
R270 B.n449 B.n448 163.367
R271 B.n448 B.n7 163.367
R272 B.n444 B.n7 163.367
R273 B.n444 B.n443 163.367
R274 B.n143 B.n142 163.367
R275 B.n143 B.n116 163.367
R276 B.n147 B.n116 163.367
R277 B.n148 B.n147 163.367
R278 B.n149 B.n148 163.367
R279 B.n149 B.n114 163.367
R280 B.n153 B.n114 163.367
R281 B.n154 B.n153 163.367
R282 B.n155 B.n154 163.367
R283 B.n155 B.n112 163.367
R284 B.n159 B.n112 163.367
R285 B.n160 B.n159 163.367
R286 B.n161 B.n160 163.367
R287 B.n161 B.n110 163.367
R288 B.n165 B.n110 163.367
R289 B.n166 B.n165 163.367
R290 B.n167 B.n166 163.367
R291 B.n167 B.n108 163.367
R292 B.n171 B.n108 163.367
R293 B.n172 B.n171 163.367
R294 B.n173 B.n172 163.367
R295 B.n173 B.n106 163.367
R296 B.n177 B.n106 163.367
R297 B.n178 B.n177 163.367
R298 B.n179 B.n178 163.367
R299 B.n179 B.n104 163.367
R300 B.n183 B.n104 163.367
R301 B.n184 B.n183 163.367
R302 B.n185 B.n184 163.367
R303 B.n185 B.n102 163.367
R304 B.n189 B.n102 163.367
R305 B.n190 B.n189 163.367
R306 B.n191 B.n190 163.367
R307 B.n191 B.n100 163.367
R308 B.n195 B.n100 163.367
R309 B.n196 B.n195 163.367
R310 B.n197 B.n196 163.367
R311 B.n197 B.n96 163.367
R312 B.n202 B.n96 163.367
R313 B.n203 B.n202 163.367
R314 B.n204 B.n203 163.367
R315 B.n204 B.n94 163.367
R316 B.n208 B.n94 163.367
R317 B.n209 B.n208 163.367
R318 B.n210 B.n209 163.367
R319 B.n210 B.n92 163.367
R320 B.n214 B.n92 163.367
R321 B.n215 B.n214 163.367
R322 B.n215 B.n88 163.367
R323 B.n219 B.n88 163.367
R324 B.n220 B.n219 163.367
R325 B.n221 B.n220 163.367
R326 B.n221 B.n86 163.367
R327 B.n225 B.n86 163.367
R328 B.n226 B.n225 163.367
R329 B.n227 B.n226 163.367
R330 B.n227 B.n84 163.367
R331 B.n231 B.n84 163.367
R332 B.n232 B.n231 163.367
R333 B.n233 B.n232 163.367
R334 B.n233 B.n82 163.367
R335 B.n237 B.n82 163.367
R336 B.n238 B.n237 163.367
R337 B.n239 B.n238 163.367
R338 B.n239 B.n80 163.367
R339 B.n243 B.n80 163.367
R340 B.n244 B.n243 163.367
R341 B.n245 B.n244 163.367
R342 B.n245 B.n78 163.367
R343 B.n249 B.n78 163.367
R344 B.n250 B.n249 163.367
R345 B.n251 B.n250 163.367
R346 B.n251 B.n76 163.367
R347 B.n255 B.n76 163.367
R348 B.n256 B.n255 163.367
R349 B.n257 B.n256 163.367
R350 B.n257 B.n74 163.367
R351 B.n261 B.n74 163.367
R352 B.n262 B.n261 163.367
R353 B.n263 B.n262 163.367
R354 B.n263 B.n72 163.367
R355 B.n267 B.n72 163.367
R356 B.n268 B.n267 163.367
R357 B.n269 B.n268 163.367
R358 B.n269 B.n70 163.367
R359 B.n274 B.n273 163.367
R360 B.n275 B.n274 163.367
R361 B.n275 B.n68 163.367
R362 B.n279 B.n68 163.367
R363 B.n280 B.n279 163.367
R364 B.n281 B.n280 163.367
R365 B.n281 B.n66 163.367
R366 B.n285 B.n66 163.367
R367 B.n286 B.n285 163.367
R368 B.n287 B.n286 163.367
R369 B.n287 B.n64 163.367
R370 B.n291 B.n64 163.367
R371 B.n292 B.n291 163.367
R372 B.n293 B.n292 163.367
R373 B.n293 B.n62 163.367
R374 B.n297 B.n62 163.367
R375 B.n298 B.n297 163.367
R376 B.n299 B.n298 163.367
R377 B.n299 B.n60 163.367
R378 B.n303 B.n60 163.367
R379 B.n304 B.n303 163.367
R380 B.n305 B.n304 163.367
R381 B.n305 B.n58 163.367
R382 B.n309 B.n58 163.367
R383 B.n310 B.n309 163.367
R384 B.n311 B.n310 163.367
R385 B.n442 B.n9 163.367
R386 B.n438 B.n9 163.367
R387 B.n438 B.n437 163.367
R388 B.n437 B.n436 163.367
R389 B.n436 B.n11 163.367
R390 B.n432 B.n11 163.367
R391 B.n432 B.n431 163.367
R392 B.n431 B.n430 163.367
R393 B.n430 B.n13 163.367
R394 B.n426 B.n13 163.367
R395 B.n426 B.n425 163.367
R396 B.n425 B.n424 163.367
R397 B.n424 B.n15 163.367
R398 B.n420 B.n15 163.367
R399 B.n420 B.n419 163.367
R400 B.n419 B.n418 163.367
R401 B.n418 B.n17 163.367
R402 B.n414 B.n17 163.367
R403 B.n414 B.n413 163.367
R404 B.n413 B.n412 163.367
R405 B.n412 B.n19 163.367
R406 B.n408 B.n19 163.367
R407 B.n408 B.n407 163.367
R408 B.n407 B.n406 163.367
R409 B.n406 B.n21 163.367
R410 B.n402 B.n21 163.367
R411 B.n402 B.n401 163.367
R412 B.n401 B.n400 163.367
R413 B.n400 B.n23 163.367
R414 B.n396 B.n23 163.367
R415 B.n396 B.n395 163.367
R416 B.n395 B.n394 163.367
R417 B.n394 B.n25 163.367
R418 B.n390 B.n25 163.367
R419 B.n390 B.n389 163.367
R420 B.n389 B.n388 163.367
R421 B.n388 B.n27 163.367
R422 B.n383 B.n27 163.367
R423 B.n383 B.n382 163.367
R424 B.n382 B.n381 163.367
R425 B.n381 B.n31 163.367
R426 B.n377 B.n31 163.367
R427 B.n377 B.n376 163.367
R428 B.n376 B.n375 163.367
R429 B.n375 B.n33 163.367
R430 B.n371 B.n33 163.367
R431 B.n371 B.n370 163.367
R432 B.n370 B.n369 163.367
R433 B.n369 B.n35 163.367
R434 B.n365 B.n35 163.367
R435 B.n365 B.n364 163.367
R436 B.n364 B.n363 163.367
R437 B.n363 B.n40 163.367
R438 B.n359 B.n40 163.367
R439 B.n359 B.n358 163.367
R440 B.n358 B.n357 163.367
R441 B.n357 B.n42 163.367
R442 B.n353 B.n42 163.367
R443 B.n353 B.n352 163.367
R444 B.n352 B.n351 163.367
R445 B.n351 B.n44 163.367
R446 B.n347 B.n44 163.367
R447 B.n347 B.n346 163.367
R448 B.n346 B.n345 163.367
R449 B.n345 B.n46 163.367
R450 B.n341 B.n46 163.367
R451 B.n341 B.n340 163.367
R452 B.n340 B.n339 163.367
R453 B.n339 B.n48 163.367
R454 B.n335 B.n48 163.367
R455 B.n335 B.n334 163.367
R456 B.n334 B.n333 163.367
R457 B.n333 B.n50 163.367
R458 B.n329 B.n50 163.367
R459 B.n329 B.n328 163.367
R460 B.n328 B.n327 163.367
R461 B.n327 B.n52 163.367
R462 B.n323 B.n52 163.367
R463 B.n323 B.n322 163.367
R464 B.n322 B.n321 163.367
R465 B.n321 B.n54 163.367
R466 B.n317 B.n54 163.367
R467 B.n317 B.n316 163.367
R468 B.n316 B.n315 163.367
R469 B.n315 B.n56 163.367
R470 B.n89 B.t8 122.906
R471 B.n36 B.t1 122.906
R472 B.n97 B.t5 122.894
R473 B.n28 B.t10 122.894
R474 B.n90 B.t7 107.391
R475 B.n37 B.t2 107.391
R476 B.n98 B.t4 107.379
R477 B.n29 B.t11 107.379
R478 B.n91 B.n90 59.5399
R479 B.n199 B.n98 59.5399
R480 B.n385 B.n29 59.5399
R481 B.n38 B.n37 59.5399
R482 B.n441 B.n8 32.3127
R483 B.n313 B.n312 32.3127
R484 B.n272 B.n271 32.3127
R485 B.n140 B.n117 32.3127
R486 B B.n463 18.0485
R487 B.n90 B.n89 15.5157
R488 B.n98 B.n97 15.5157
R489 B.n29 B.n28 15.5157
R490 B.n37 B.n36 15.5157
R491 B.n441 B.n440 10.6151
R492 B.n440 B.n439 10.6151
R493 B.n439 B.n10 10.6151
R494 B.n435 B.n10 10.6151
R495 B.n435 B.n434 10.6151
R496 B.n434 B.n433 10.6151
R497 B.n433 B.n12 10.6151
R498 B.n429 B.n12 10.6151
R499 B.n429 B.n428 10.6151
R500 B.n428 B.n427 10.6151
R501 B.n427 B.n14 10.6151
R502 B.n423 B.n14 10.6151
R503 B.n423 B.n422 10.6151
R504 B.n422 B.n421 10.6151
R505 B.n421 B.n16 10.6151
R506 B.n417 B.n16 10.6151
R507 B.n417 B.n416 10.6151
R508 B.n416 B.n415 10.6151
R509 B.n415 B.n18 10.6151
R510 B.n411 B.n18 10.6151
R511 B.n411 B.n410 10.6151
R512 B.n410 B.n409 10.6151
R513 B.n409 B.n20 10.6151
R514 B.n405 B.n20 10.6151
R515 B.n405 B.n404 10.6151
R516 B.n404 B.n403 10.6151
R517 B.n403 B.n22 10.6151
R518 B.n399 B.n22 10.6151
R519 B.n399 B.n398 10.6151
R520 B.n398 B.n397 10.6151
R521 B.n397 B.n24 10.6151
R522 B.n393 B.n24 10.6151
R523 B.n393 B.n392 10.6151
R524 B.n392 B.n391 10.6151
R525 B.n391 B.n26 10.6151
R526 B.n387 B.n26 10.6151
R527 B.n387 B.n386 10.6151
R528 B.n384 B.n30 10.6151
R529 B.n380 B.n30 10.6151
R530 B.n380 B.n379 10.6151
R531 B.n379 B.n378 10.6151
R532 B.n378 B.n32 10.6151
R533 B.n374 B.n32 10.6151
R534 B.n374 B.n373 10.6151
R535 B.n373 B.n372 10.6151
R536 B.n372 B.n34 10.6151
R537 B.n368 B.n367 10.6151
R538 B.n367 B.n366 10.6151
R539 B.n366 B.n39 10.6151
R540 B.n362 B.n39 10.6151
R541 B.n362 B.n361 10.6151
R542 B.n361 B.n360 10.6151
R543 B.n360 B.n41 10.6151
R544 B.n356 B.n41 10.6151
R545 B.n356 B.n355 10.6151
R546 B.n355 B.n354 10.6151
R547 B.n354 B.n43 10.6151
R548 B.n350 B.n43 10.6151
R549 B.n350 B.n349 10.6151
R550 B.n349 B.n348 10.6151
R551 B.n348 B.n45 10.6151
R552 B.n344 B.n45 10.6151
R553 B.n344 B.n343 10.6151
R554 B.n343 B.n342 10.6151
R555 B.n342 B.n47 10.6151
R556 B.n338 B.n47 10.6151
R557 B.n338 B.n337 10.6151
R558 B.n337 B.n336 10.6151
R559 B.n336 B.n49 10.6151
R560 B.n332 B.n49 10.6151
R561 B.n332 B.n331 10.6151
R562 B.n331 B.n330 10.6151
R563 B.n330 B.n51 10.6151
R564 B.n326 B.n51 10.6151
R565 B.n326 B.n325 10.6151
R566 B.n325 B.n324 10.6151
R567 B.n324 B.n53 10.6151
R568 B.n320 B.n53 10.6151
R569 B.n320 B.n319 10.6151
R570 B.n319 B.n318 10.6151
R571 B.n318 B.n55 10.6151
R572 B.n314 B.n55 10.6151
R573 B.n314 B.n313 10.6151
R574 B.n272 B.n69 10.6151
R575 B.n276 B.n69 10.6151
R576 B.n277 B.n276 10.6151
R577 B.n278 B.n277 10.6151
R578 B.n278 B.n67 10.6151
R579 B.n282 B.n67 10.6151
R580 B.n283 B.n282 10.6151
R581 B.n284 B.n283 10.6151
R582 B.n284 B.n65 10.6151
R583 B.n288 B.n65 10.6151
R584 B.n289 B.n288 10.6151
R585 B.n290 B.n289 10.6151
R586 B.n290 B.n63 10.6151
R587 B.n294 B.n63 10.6151
R588 B.n295 B.n294 10.6151
R589 B.n296 B.n295 10.6151
R590 B.n296 B.n61 10.6151
R591 B.n300 B.n61 10.6151
R592 B.n301 B.n300 10.6151
R593 B.n302 B.n301 10.6151
R594 B.n302 B.n59 10.6151
R595 B.n306 B.n59 10.6151
R596 B.n307 B.n306 10.6151
R597 B.n308 B.n307 10.6151
R598 B.n308 B.n57 10.6151
R599 B.n312 B.n57 10.6151
R600 B.n144 B.n117 10.6151
R601 B.n145 B.n144 10.6151
R602 B.n146 B.n145 10.6151
R603 B.n146 B.n115 10.6151
R604 B.n150 B.n115 10.6151
R605 B.n151 B.n150 10.6151
R606 B.n152 B.n151 10.6151
R607 B.n152 B.n113 10.6151
R608 B.n156 B.n113 10.6151
R609 B.n157 B.n156 10.6151
R610 B.n158 B.n157 10.6151
R611 B.n158 B.n111 10.6151
R612 B.n162 B.n111 10.6151
R613 B.n163 B.n162 10.6151
R614 B.n164 B.n163 10.6151
R615 B.n164 B.n109 10.6151
R616 B.n168 B.n109 10.6151
R617 B.n169 B.n168 10.6151
R618 B.n170 B.n169 10.6151
R619 B.n170 B.n107 10.6151
R620 B.n174 B.n107 10.6151
R621 B.n175 B.n174 10.6151
R622 B.n176 B.n175 10.6151
R623 B.n176 B.n105 10.6151
R624 B.n180 B.n105 10.6151
R625 B.n181 B.n180 10.6151
R626 B.n182 B.n181 10.6151
R627 B.n182 B.n103 10.6151
R628 B.n186 B.n103 10.6151
R629 B.n187 B.n186 10.6151
R630 B.n188 B.n187 10.6151
R631 B.n188 B.n101 10.6151
R632 B.n192 B.n101 10.6151
R633 B.n193 B.n192 10.6151
R634 B.n194 B.n193 10.6151
R635 B.n194 B.n99 10.6151
R636 B.n198 B.n99 10.6151
R637 B.n201 B.n200 10.6151
R638 B.n201 B.n95 10.6151
R639 B.n205 B.n95 10.6151
R640 B.n206 B.n205 10.6151
R641 B.n207 B.n206 10.6151
R642 B.n207 B.n93 10.6151
R643 B.n211 B.n93 10.6151
R644 B.n212 B.n211 10.6151
R645 B.n213 B.n212 10.6151
R646 B.n217 B.n216 10.6151
R647 B.n218 B.n217 10.6151
R648 B.n218 B.n87 10.6151
R649 B.n222 B.n87 10.6151
R650 B.n223 B.n222 10.6151
R651 B.n224 B.n223 10.6151
R652 B.n224 B.n85 10.6151
R653 B.n228 B.n85 10.6151
R654 B.n229 B.n228 10.6151
R655 B.n230 B.n229 10.6151
R656 B.n230 B.n83 10.6151
R657 B.n234 B.n83 10.6151
R658 B.n235 B.n234 10.6151
R659 B.n236 B.n235 10.6151
R660 B.n236 B.n81 10.6151
R661 B.n240 B.n81 10.6151
R662 B.n241 B.n240 10.6151
R663 B.n242 B.n241 10.6151
R664 B.n242 B.n79 10.6151
R665 B.n246 B.n79 10.6151
R666 B.n247 B.n246 10.6151
R667 B.n248 B.n247 10.6151
R668 B.n248 B.n77 10.6151
R669 B.n252 B.n77 10.6151
R670 B.n253 B.n252 10.6151
R671 B.n254 B.n253 10.6151
R672 B.n254 B.n75 10.6151
R673 B.n258 B.n75 10.6151
R674 B.n259 B.n258 10.6151
R675 B.n260 B.n259 10.6151
R676 B.n260 B.n73 10.6151
R677 B.n264 B.n73 10.6151
R678 B.n265 B.n264 10.6151
R679 B.n266 B.n265 10.6151
R680 B.n266 B.n71 10.6151
R681 B.n270 B.n71 10.6151
R682 B.n271 B.n270 10.6151
R683 B.n140 B.n139 10.6151
R684 B.n139 B.n138 10.6151
R685 B.n138 B.n119 10.6151
R686 B.n134 B.n119 10.6151
R687 B.n134 B.n133 10.6151
R688 B.n133 B.n132 10.6151
R689 B.n132 B.n121 10.6151
R690 B.n128 B.n121 10.6151
R691 B.n128 B.n127 10.6151
R692 B.n127 B.n126 10.6151
R693 B.n126 B.n123 10.6151
R694 B.n123 B.n0 10.6151
R695 B.n459 B.n1 10.6151
R696 B.n459 B.n458 10.6151
R697 B.n458 B.n457 10.6151
R698 B.n457 B.n4 10.6151
R699 B.n453 B.n4 10.6151
R700 B.n453 B.n452 10.6151
R701 B.n452 B.n451 10.6151
R702 B.n451 B.n6 10.6151
R703 B.n447 B.n6 10.6151
R704 B.n447 B.n446 10.6151
R705 B.n446 B.n445 10.6151
R706 B.n445 B.n8 10.6151
R707 B.n386 B.n385 8.74196
R708 B.n368 B.n38 8.74196
R709 B.n199 B.n198 8.74196
R710 B.n216 B.n91 8.74196
R711 B.n463 B.n0 2.81026
R712 B.n463 B.n1 2.81026
R713 B.n385 B.n384 1.87367
R714 B.n38 B.n34 1.87367
R715 B.n200 B.n199 1.87367
R716 B.n213 B.n91 1.87367
R717 VP.n0 VP.t0 841.971
R718 VP.n0 VP.t1 803.797
R719 VP VP.n0 0.0516364
R720 VDD1 VDD1.t0 116.763
R721 VDD1 VDD1.t1 81.8612
C0 VTAIL VDD1 5.72824f
C1 B w_n1290_n3148# 6.19685f
C2 w_n1290_n3148# VN 1.58815f
C3 VP VDD2 0.244942f
C4 B VN 0.67236f
C5 VP VDD1 1.66501f
C6 w_n1290_n3148# VTAIL 2.78066f
C7 B VTAIL 2.39352f
C8 VTAIL VN 1.07592f
C9 VDD1 VDD2 0.440684f
C10 VP w_n1290_n3148# 1.74788f
C11 B VP 0.926416f
C12 VP VN 4.25229f
C13 w_n1290_n3148# VDD2 1.46663f
C14 w_n1290_n3148# VDD1 1.46428f
C15 B VDD2 1.30556f
C16 VP VTAIL 1.09055f
C17 VN VDD2 1.57255f
C18 B VDD1 1.29259f
C19 VN VDD1 0.148151f
C20 VTAIL VDD2 5.76025f
C21 VDD2 VSUBS 0.688848f
C22 VDD1 VSUBS 3.202831f
C23 VTAIL VSUBS 0.246296f
C24 VN VSUBS 4.52988f
C25 VP VSUBS 0.999273f
C26 B VSUBS 2.23395f
C27 w_n1290_n3148# VSUBS 50.0778f
C28 VDD1.t1 VSUBS 1.46857f
C29 VDD1.t0 VSUBS 1.82403f
C30 VP.t0 VSUBS 0.67626f
C31 VP.t1 VSUBS 0.607136f
C32 VP.n0 VSUBS 3.00866f
C33 B.n0 VSUBS 0.004931f
C34 B.n1 VSUBS 0.004931f
C35 B.n2 VSUBS 0.007798f
C36 B.n3 VSUBS 0.007798f
C37 B.n4 VSUBS 0.007798f
C38 B.n5 VSUBS 0.007798f
C39 B.n6 VSUBS 0.007798f
C40 B.n7 VSUBS 0.007798f
C41 B.n8 VSUBS 0.017949f
C42 B.n9 VSUBS 0.007798f
C43 B.n10 VSUBS 0.007798f
C44 B.n11 VSUBS 0.007798f
C45 B.n12 VSUBS 0.007798f
C46 B.n13 VSUBS 0.007798f
C47 B.n14 VSUBS 0.007798f
C48 B.n15 VSUBS 0.007798f
C49 B.n16 VSUBS 0.007798f
C50 B.n17 VSUBS 0.007798f
C51 B.n18 VSUBS 0.007798f
C52 B.n19 VSUBS 0.007798f
C53 B.n20 VSUBS 0.007798f
C54 B.n21 VSUBS 0.007798f
C55 B.n22 VSUBS 0.007798f
C56 B.n23 VSUBS 0.007798f
C57 B.n24 VSUBS 0.007798f
C58 B.n25 VSUBS 0.007798f
C59 B.n26 VSUBS 0.007798f
C60 B.n27 VSUBS 0.007798f
C61 B.t11 VSUBS 0.39063f
C62 B.t10 VSUBS 0.398073f
C63 B.t9 VSUBS 0.230272f
C64 B.n28 VSUBS 0.120783f
C65 B.n29 VSUBS 0.070076f
C66 B.n30 VSUBS 0.007798f
C67 B.n31 VSUBS 0.007798f
C68 B.n32 VSUBS 0.007798f
C69 B.n33 VSUBS 0.007798f
C70 B.n34 VSUBS 0.004587f
C71 B.n35 VSUBS 0.007798f
C72 B.t2 VSUBS 0.390623f
C73 B.t1 VSUBS 0.398066f
C74 B.t0 VSUBS 0.230272f
C75 B.n36 VSUBS 0.120789f
C76 B.n37 VSUBS 0.070083f
C77 B.n38 VSUBS 0.018068f
C78 B.n39 VSUBS 0.007798f
C79 B.n40 VSUBS 0.007798f
C80 B.n41 VSUBS 0.007798f
C81 B.n42 VSUBS 0.007798f
C82 B.n43 VSUBS 0.007798f
C83 B.n44 VSUBS 0.007798f
C84 B.n45 VSUBS 0.007798f
C85 B.n46 VSUBS 0.007798f
C86 B.n47 VSUBS 0.007798f
C87 B.n48 VSUBS 0.007798f
C88 B.n49 VSUBS 0.007798f
C89 B.n50 VSUBS 0.007798f
C90 B.n51 VSUBS 0.007798f
C91 B.n52 VSUBS 0.007798f
C92 B.n53 VSUBS 0.007798f
C93 B.n54 VSUBS 0.007798f
C94 B.n55 VSUBS 0.007798f
C95 B.n56 VSUBS 0.01829f
C96 B.n57 VSUBS 0.007798f
C97 B.n58 VSUBS 0.007798f
C98 B.n59 VSUBS 0.007798f
C99 B.n60 VSUBS 0.007798f
C100 B.n61 VSUBS 0.007798f
C101 B.n62 VSUBS 0.007798f
C102 B.n63 VSUBS 0.007798f
C103 B.n64 VSUBS 0.007798f
C104 B.n65 VSUBS 0.007798f
C105 B.n66 VSUBS 0.007798f
C106 B.n67 VSUBS 0.007798f
C107 B.n68 VSUBS 0.007798f
C108 B.n69 VSUBS 0.007798f
C109 B.n70 VSUBS 0.01829f
C110 B.n71 VSUBS 0.007798f
C111 B.n72 VSUBS 0.007798f
C112 B.n73 VSUBS 0.007798f
C113 B.n74 VSUBS 0.007798f
C114 B.n75 VSUBS 0.007798f
C115 B.n76 VSUBS 0.007798f
C116 B.n77 VSUBS 0.007798f
C117 B.n78 VSUBS 0.007798f
C118 B.n79 VSUBS 0.007798f
C119 B.n80 VSUBS 0.007798f
C120 B.n81 VSUBS 0.007798f
C121 B.n82 VSUBS 0.007798f
C122 B.n83 VSUBS 0.007798f
C123 B.n84 VSUBS 0.007798f
C124 B.n85 VSUBS 0.007798f
C125 B.n86 VSUBS 0.007798f
C126 B.n87 VSUBS 0.007798f
C127 B.n88 VSUBS 0.007798f
C128 B.t7 VSUBS 0.390623f
C129 B.t8 VSUBS 0.398066f
C130 B.t6 VSUBS 0.230272f
C131 B.n89 VSUBS 0.120789f
C132 B.n90 VSUBS 0.070083f
C133 B.n91 VSUBS 0.018068f
C134 B.n92 VSUBS 0.007798f
C135 B.n93 VSUBS 0.007798f
C136 B.n94 VSUBS 0.007798f
C137 B.n95 VSUBS 0.007798f
C138 B.n96 VSUBS 0.007798f
C139 B.t4 VSUBS 0.39063f
C140 B.t5 VSUBS 0.398073f
C141 B.t3 VSUBS 0.230272f
C142 B.n97 VSUBS 0.120783f
C143 B.n98 VSUBS 0.070076f
C144 B.n99 VSUBS 0.007798f
C145 B.n100 VSUBS 0.007798f
C146 B.n101 VSUBS 0.007798f
C147 B.n102 VSUBS 0.007798f
C148 B.n103 VSUBS 0.007798f
C149 B.n104 VSUBS 0.007798f
C150 B.n105 VSUBS 0.007798f
C151 B.n106 VSUBS 0.007798f
C152 B.n107 VSUBS 0.007798f
C153 B.n108 VSUBS 0.007798f
C154 B.n109 VSUBS 0.007798f
C155 B.n110 VSUBS 0.007798f
C156 B.n111 VSUBS 0.007798f
C157 B.n112 VSUBS 0.007798f
C158 B.n113 VSUBS 0.007798f
C159 B.n114 VSUBS 0.007798f
C160 B.n115 VSUBS 0.007798f
C161 B.n116 VSUBS 0.007798f
C162 B.n117 VSUBS 0.01829f
C163 B.n118 VSUBS 0.007798f
C164 B.n119 VSUBS 0.007798f
C165 B.n120 VSUBS 0.007798f
C166 B.n121 VSUBS 0.007798f
C167 B.n122 VSUBS 0.007798f
C168 B.n123 VSUBS 0.007798f
C169 B.n124 VSUBS 0.007798f
C170 B.n125 VSUBS 0.007798f
C171 B.n126 VSUBS 0.007798f
C172 B.n127 VSUBS 0.007798f
C173 B.n128 VSUBS 0.007798f
C174 B.n129 VSUBS 0.007798f
C175 B.n130 VSUBS 0.007798f
C176 B.n131 VSUBS 0.007798f
C177 B.n132 VSUBS 0.007798f
C178 B.n133 VSUBS 0.007798f
C179 B.n134 VSUBS 0.007798f
C180 B.n135 VSUBS 0.007798f
C181 B.n136 VSUBS 0.007798f
C182 B.n137 VSUBS 0.007798f
C183 B.n138 VSUBS 0.007798f
C184 B.n139 VSUBS 0.007798f
C185 B.n140 VSUBS 0.017949f
C186 B.n141 VSUBS 0.017949f
C187 B.n142 VSUBS 0.01829f
C188 B.n143 VSUBS 0.007798f
C189 B.n144 VSUBS 0.007798f
C190 B.n145 VSUBS 0.007798f
C191 B.n146 VSUBS 0.007798f
C192 B.n147 VSUBS 0.007798f
C193 B.n148 VSUBS 0.007798f
C194 B.n149 VSUBS 0.007798f
C195 B.n150 VSUBS 0.007798f
C196 B.n151 VSUBS 0.007798f
C197 B.n152 VSUBS 0.007798f
C198 B.n153 VSUBS 0.007798f
C199 B.n154 VSUBS 0.007798f
C200 B.n155 VSUBS 0.007798f
C201 B.n156 VSUBS 0.007798f
C202 B.n157 VSUBS 0.007798f
C203 B.n158 VSUBS 0.007798f
C204 B.n159 VSUBS 0.007798f
C205 B.n160 VSUBS 0.007798f
C206 B.n161 VSUBS 0.007798f
C207 B.n162 VSUBS 0.007798f
C208 B.n163 VSUBS 0.007798f
C209 B.n164 VSUBS 0.007798f
C210 B.n165 VSUBS 0.007798f
C211 B.n166 VSUBS 0.007798f
C212 B.n167 VSUBS 0.007798f
C213 B.n168 VSUBS 0.007798f
C214 B.n169 VSUBS 0.007798f
C215 B.n170 VSUBS 0.007798f
C216 B.n171 VSUBS 0.007798f
C217 B.n172 VSUBS 0.007798f
C218 B.n173 VSUBS 0.007798f
C219 B.n174 VSUBS 0.007798f
C220 B.n175 VSUBS 0.007798f
C221 B.n176 VSUBS 0.007798f
C222 B.n177 VSUBS 0.007798f
C223 B.n178 VSUBS 0.007798f
C224 B.n179 VSUBS 0.007798f
C225 B.n180 VSUBS 0.007798f
C226 B.n181 VSUBS 0.007798f
C227 B.n182 VSUBS 0.007798f
C228 B.n183 VSUBS 0.007798f
C229 B.n184 VSUBS 0.007798f
C230 B.n185 VSUBS 0.007798f
C231 B.n186 VSUBS 0.007798f
C232 B.n187 VSUBS 0.007798f
C233 B.n188 VSUBS 0.007798f
C234 B.n189 VSUBS 0.007798f
C235 B.n190 VSUBS 0.007798f
C236 B.n191 VSUBS 0.007798f
C237 B.n192 VSUBS 0.007798f
C238 B.n193 VSUBS 0.007798f
C239 B.n194 VSUBS 0.007798f
C240 B.n195 VSUBS 0.007798f
C241 B.n196 VSUBS 0.007798f
C242 B.n197 VSUBS 0.007798f
C243 B.n198 VSUBS 0.00711f
C244 B.n199 VSUBS 0.018068f
C245 B.n200 VSUBS 0.004587f
C246 B.n201 VSUBS 0.007798f
C247 B.n202 VSUBS 0.007798f
C248 B.n203 VSUBS 0.007798f
C249 B.n204 VSUBS 0.007798f
C250 B.n205 VSUBS 0.007798f
C251 B.n206 VSUBS 0.007798f
C252 B.n207 VSUBS 0.007798f
C253 B.n208 VSUBS 0.007798f
C254 B.n209 VSUBS 0.007798f
C255 B.n210 VSUBS 0.007798f
C256 B.n211 VSUBS 0.007798f
C257 B.n212 VSUBS 0.007798f
C258 B.n213 VSUBS 0.004587f
C259 B.n214 VSUBS 0.007798f
C260 B.n215 VSUBS 0.007798f
C261 B.n216 VSUBS 0.00711f
C262 B.n217 VSUBS 0.007798f
C263 B.n218 VSUBS 0.007798f
C264 B.n219 VSUBS 0.007798f
C265 B.n220 VSUBS 0.007798f
C266 B.n221 VSUBS 0.007798f
C267 B.n222 VSUBS 0.007798f
C268 B.n223 VSUBS 0.007798f
C269 B.n224 VSUBS 0.007798f
C270 B.n225 VSUBS 0.007798f
C271 B.n226 VSUBS 0.007798f
C272 B.n227 VSUBS 0.007798f
C273 B.n228 VSUBS 0.007798f
C274 B.n229 VSUBS 0.007798f
C275 B.n230 VSUBS 0.007798f
C276 B.n231 VSUBS 0.007798f
C277 B.n232 VSUBS 0.007798f
C278 B.n233 VSUBS 0.007798f
C279 B.n234 VSUBS 0.007798f
C280 B.n235 VSUBS 0.007798f
C281 B.n236 VSUBS 0.007798f
C282 B.n237 VSUBS 0.007798f
C283 B.n238 VSUBS 0.007798f
C284 B.n239 VSUBS 0.007798f
C285 B.n240 VSUBS 0.007798f
C286 B.n241 VSUBS 0.007798f
C287 B.n242 VSUBS 0.007798f
C288 B.n243 VSUBS 0.007798f
C289 B.n244 VSUBS 0.007798f
C290 B.n245 VSUBS 0.007798f
C291 B.n246 VSUBS 0.007798f
C292 B.n247 VSUBS 0.007798f
C293 B.n248 VSUBS 0.007798f
C294 B.n249 VSUBS 0.007798f
C295 B.n250 VSUBS 0.007798f
C296 B.n251 VSUBS 0.007798f
C297 B.n252 VSUBS 0.007798f
C298 B.n253 VSUBS 0.007798f
C299 B.n254 VSUBS 0.007798f
C300 B.n255 VSUBS 0.007798f
C301 B.n256 VSUBS 0.007798f
C302 B.n257 VSUBS 0.007798f
C303 B.n258 VSUBS 0.007798f
C304 B.n259 VSUBS 0.007798f
C305 B.n260 VSUBS 0.007798f
C306 B.n261 VSUBS 0.007798f
C307 B.n262 VSUBS 0.007798f
C308 B.n263 VSUBS 0.007798f
C309 B.n264 VSUBS 0.007798f
C310 B.n265 VSUBS 0.007798f
C311 B.n266 VSUBS 0.007798f
C312 B.n267 VSUBS 0.007798f
C313 B.n268 VSUBS 0.007798f
C314 B.n269 VSUBS 0.007798f
C315 B.n270 VSUBS 0.007798f
C316 B.n271 VSUBS 0.01829f
C317 B.n272 VSUBS 0.017949f
C318 B.n273 VSUBS 0.017949f
C319 B.n274 VSUBS 0.007798f
C320 B.n275 VSUBS 0.007798f
C321 B.n276 VSUBS 0.007798f
C322 B.n277 VSUBS 0.007798f
C323 B.n278 VSUBS 0.007798f
C324 B.n279 VSUBS 0.007798f
C325 B.n280 VSUBS 0.007798f
C326 B.n281 VSUBS 0.007798f
C327 B.n282 VSUBS 0.007798f
C328 B.n283 VSUBS 0.007798f
C329 B.n284 VSUBS 0.007798f
C330 B.n285 VSUBS 0.007798f
C331 B.n286 VSUBS 0.007798f
C332 B.n287 VSUBS 0.007798f
C333 B.n288 VSUBS 0.007798f
C334 B.n289 VSUBS 0.007798f
C335 B.n290 VSUBS 0.007798f
C336 B.n291 VSUBS 0.007798f
C337 B.n292 VSUBS 0.007798f
C338 B.n293 VSUBS 0.007798f
C339 B.n294 VSUBS 0.007798f
C340 B.n295 VSUBS 0.007798f
C341 B.n296 VSUBS 0.007798f
C342 B.n297 VSUBS 0.007798f
C343 B.n298 VSUBS 0.007798f
C344 B.n299 VSUBS 0.007798f
C345 B.n300 VSUBS 0.007798f
C346 B.n301 VSUBS 0.007798f
C347 B.n302 VSUBS 0.007798f
C348 B.n303 VSUBS 0.007798f
C349 B.n304 VSUBS 0.007798f
C350 B.n305 VSUBS 0.007798f
C351 B.n306 VSUBS 0.007798f
C352 B.n307 VSUBS 0.007798f
C353 B.n308 VSUBS 0.007798f
C354 B.n309 VSUBS 0.007798f
C355 B.n310 VSUBS 0.007798f
C356 B.n311 VSUBS 0.017949f
C357 B.n312 VSUBS 0.018881f
C358 B.n313 VSUBS 0.017359f
C359 B.n314 VSUBS 0.007798f
C360 B.n315 VSUBS 0.007798f
C361 B.n316 VSUBS 0.007798f
C362 B.n317 VSUBS 0.007798f
C363 B.n318 VSUBS 0.007798f
C364 B.n319 VSUBS 0.007798f
C365 B.n320 VSUBS 0.007798f
C366 B.n321 VSUBS 0.007798f
C367 B.n322 VSUBS 0.007798f
C368 B.n323 VSUBS 0.007798f
C369 B.n324 VSUBS 0.007798f
C370 B.n325 VSUBS 0.007798f
C371 B.n326 VSUBS 0.007798f
C372 B.n327 VSUBS 0.007798f
C373 B.n328 VSUBS 0.007798f
C374 B.n329 VSUBS 0.007798f
C375 B.n330 VSUBS 0.007798f
C376 B.n331 VSUBS 0.007798f
C377 B.n332 VSUBS 0.007798f
C378 B.n333 VSUBS 0.007798f
C379 B.n334 VSUBS 0.007798f
C380 B.n335 VSUBS 0.007798f
C381 B.n336 VSUBS 0.007798f
C382 B.n337 VSUBS 0.007798f
C383 B.n338 VSUBS 0.007798f
C384 B.n339 VSUBS 0.007798f
C385 B.n340 VSUBS 0.007798f
C386 B.n341 VSUBS 0.007798f
C387 B.n342 VSUBS 0.007798f
C388 B.n343 VSUBS 0.007798f
C389 B.n344 VSUBS 0.007798f
C390 B.n345 VSUBS 0.007798f
C391 B.n346 VSUBS 0.007798f
C392 B.n347 VSUBS 0.007798f
C393 B.n348 VSUBS 0.007798f
C394 B.n349 VSUBS 0.007798f
C395 B.n350 VSUBS 0.007798f
C396 B.n351 VSUBS 0.007798f
C397 B.n352 VSUBS 0.007798f
C398 B.n353 VSUBS 0.007798f
C399 B.n354 VSUBS 0.007798f
C400 B.n355 VSUBS 0.007798f
C401 B.n356 VSUBS 0.007798f
C402 B.n357 VSUBS 0.007798f
C403 B.n358 VSUBS 0.007798f
C404 B.n359 VSUBS 0.007798f
C405 B.n360 VSUBS 0.007798f
C406 B.n361 VSUBS 0.007798f
C407 B.n362 VSUBS 0.007798f
C408 B.n363 VSUBS 0.007798f
C409 B.n364 VSUBS 0.007798f
C410 B.n365 VSUBS 0.007798f
C411 B.n366 VSUBS 0.007798f
C412 B.n367 VSUBS 0.007798f
C413 B.n368 VSUBS 0.00711f
C414 B.n369 VSUBS 0.007798f
C415 B.n370 VSUBS 0.007798f
C416 B.n371 VSUBS 0.007798f
C417 B.n372 VSUBS 0.007798f
C418 B.n373 VSUBS 0.007798f
C419 B.n374 VSUBS 0.007798f
C420 B.n375 VSUBS 0.007798f
C421 B.n376 VSUBS 0.007798f
C422 B.n377 VSUBS 0.007798f
C423 B.n378 VSUBS 0.007798f
C424 B.n379 VSUBS 0.007798f
C425 B.n380 VSUBS 0.007798f
C426 B.n381 VSUBS 0.007798f
C427 B.n382 VSUBS 0.007798f
C428 B.n383 VSUBS 0.007798f
C429 B.n384 VSUBS 0.004587f
C430 B.n385 VSUBS 0.018068f
C431 B.n386 VSUBS 0.00711f
C432 B.n387 VSUBS 0.007798f
C433 B.n388 VSUBS 0.007798f
C434 B.n389 VSUBS 0.007798f
C435 B.n390 VSUBS 0.007798f
C436 B.n391 VSUBS 0.007798f
C437 B.n392 VSUBS 0.007798f
C438 B.n393 VSUBS 0.007798f
C439 B.n394 VSUBS 0.007798f
C440 B.n395 VSUBS 0.007798f
C441 B.n396 VSUBS 0.007798f
C442 B.n397 VSUBS 0.007798f
C443 B.n398 VSUBS 0.007798f
C444 B.n399 VSUBS 0.007798f
C445 B.n400 VSUBS 0.007798f
C446 B.n401 VSUBS 0.007798f
C447 B.n402 VSUBS 0.007798f
C448 B.n403 VSUBS 0.007798f
C449 B.n404 VSUBS 0.007798f
C450 B.n405 VSUBS 0.007798f
C451 B.n406 VSUBS 0.007798f
C452 B.n407 VSUBS 0.007798f
C453 B.n408 VSUBS 0.007798f
C454 B.n409 VSUBS 0.007798f
C455 B.n410 VSUBS 0.007798f
C456 B.n411 VSUBS 0.007798f
C457 B.n412 VSUBS 0.007798f
C458 B.n413 VSUBS 0.007798f
C459 B.n414 VSUBS 0.007798f
C460 B.n415 VSUBS 0.007798f
C461 B.n416 VSUBS 0.007798f
C462 B.n417 VSUBS 0.007798f
C463 B.n418 VSUBS 0.007798f
C464 B.n419 VSUBS 0.007798f
C465 B.n420 VSUBS 0.007798f
C466 B.n421 VSUBS 0.007798f
C467 B.n422 VSUBS 0.007798f
C468 B.n423 VSUBS 0.007798f
C469 B.n424 VSUBS 0.007798f
C470 B.n425 VSUBS 0.007798f
C471 B.n426 VSUBS 0.007798f
C472 B.n427 VSUBS 0.007798f
C473 B.n428 VSUBS 0.007798f
C474 B.n429 VSUBS 0.007798f
C475 B.n430 VSUBS 0.007798f
C476 B.n431 VSUBS 0.007798f
C477 B.n432 VSUBS 0.007798f
C478 B.n433 VSUBS 0.007798f
C479 B.n434 VSUBS 0.007798f
C480 B.n435 VSUBS 0.007798f
C481 B.n436 VSUBS 0.007798f
C482 B.n437 VSUBS 0.007798f
C483 B.n438 VSUBS 0.007798f
C484 B.n439 VSUBS 0.007798f
C485 B.n440 VSUBS 0.007798f
C486 B.n441 VSUBS 0.01829f
C487 B.n442 VSUBS 0.01829f
C488 B.n443 VSUBS 0.017949f
C489 B.n444 VSUBS 0.007798f
C490 B.n445 VSUBS 0.007798f
C491 B.n446 VSUBS 0.007798f
C492 B.n447 VSUBS 0.007798f
C493 B.n448 VSUBS 0.007798f
C494 B.n449 VSUBS 0.007798f
C495 B.n450 VSUBS 0.007798f
C496 B.n451 VSUBS 0.007798f
C497 B.n452 VSUBS 0.007798f
C498 B.n453 VSUBS 0.007798f
C499 B.n454 VSUBS 0.007798f
C500 B.n455 VSUBS 0.007798f
C501 B.n456 VSUBS 0.007798f
C502 B.n457 VSUBS 0.007798f
C503 B.n458 VSUBS 0.007798f
C504 B.n459 VSUBS 0.007798f
C505 B.n460 VSUBS 0.007798f
C506 B.n461 VSUBS 0.007798f
C507 B.n462 VSUBS 0.007798f
C508 B.n463 VSUBS 0.017658f
C509 VDD2.t1 VSUBS 1.85908f
C510 VDD2.t0 VSUBS 1.50973f
C511 VDD2.n0 VSUBS 2.39864f
C512 VTAIL.t0 VSUBS 2.19351f
C513 VTAIL.n0 VSUBS 2.00134f
C514 VTAIL.t3 VSUBS 2.19351f
C515 VTAIL.n1 VSUBS 2.01117f
C516 VTAIL.t1 VSUBS 2.1935f
C517 VTAIL.n2 VSUBS 1.95181f
C518 VTAIL.t2 VSUBS 2.19351f
C519 VTAIL.n3 VSUBS 1.8915f
C520 VN.t0 VSUBS 0.599608f
C521 VN.t1 VSUBS 0.669659f
.ends

