* NGSPICE file created from diff_pair_sample_1185.ext - technology: sky130A

.subckt diff_pair_sample_1185 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t4 VN.t0 VDD2.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.5031 pd=3.36 as=0.21285 ps=1.62 w=1.29 l=0.87
X1 VTAIL.t7 VP.t0 VDD1.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.5031 pd=3.36 as=0.21285 ps=1.62 w=1.29 l=0.87
X2 B.t17 B.t15 B.t16 B.t9 sky130_fd_pr__nfet_01v8 ad=0.5031 pd=3.36 as=0 ps=0 w=1.29 l=0.87
X3 B.t14 B.t12 B.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=0.5031 pd=3.36 as=0 ps=0 w=1.29 l=0.87
X4 VTAIL.t3 VN.t1 VDD2.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=0.5031 pd=3.36 as=0.21285 ps=1.62 w=1.29 l=0.87
X5 VTAIL.t6 VP.t1 VDD1.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.5031 pd=3.36 as=0.21285 ps=1.62 w=1.29 l=0.87
X6 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=0.5031 pd=3.36 as=0 ps=0 w=1.29 l=0.87
X7 VDD2.t2 VN.t2 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=0.21285 pd=1.62 as=0.5031 ps=3.36 w=1.29 l=0.87
X8 VDD2.t0 VN.t3 VTAIL.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=0.21285 pd=1.62 as=0.5031 ps=3.36 w=1.29 l=0.87
X9 VDD1.t1 VP.t2 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.21285 pd=1.62 as=0.5031 ps=3.36 w=1.29 l=0.87
X10 VDD1.t0 VP.t3 VTAIL.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=0.21285 pd=1.62 as=0.5031 ps=3.36 w=1.29 l=0.87
X11 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=0.5031 pd=3.36 as=0 ps=0 w=1.29 l=0.87
R0 VN.n0 VN.t1 102.162
R1 VN.n1 VN.t2 102.162
R2 VN.n0 VN.t3 102.112
R3 VN.n1 VN.t0 102.112
R4 VN VN.n1 77.9822
R5 VN VN.n0 44.7132
R6 VDD2.n2 VDD2.n0 174.554
R7 VDD2.n2 VDD2.n1 146.623
R8 VDD2.n1 VDD2.t3 15.3493
R9 VDD2.n1 VDD2.t2 15.3493
R10 VDD2.n0 VDD2.t1 15.3493
R11 VDD2.n0 VDD2.t0 15.3493
R12 VDD2 VDD2.n2 0.0586897
R13 VTAIL.n7 VTAIL.t1 156.102
R14 VTAIL.n0 VTAIL.t3 156.102
R15 VTAIL.n1 VTAIL.t5 156.102
R16 VTAIL.n2 VTAIL.t7 156.102
R17 VTAIL.n6 VTAIL.t0 156.102
R18 VTAIL.n5 VTAIL.t6 156.102
R19 VTAIL.n4 VTAIL.t2 156.102
R20 VTAIL.n3 VTAIL.t4 156.102
R21 VTAIL.n7 VTAIL.n6 14.5134
R22 VTAIL.n3 VTAIL.n2 14.5134
R23 VTAIL.n4 VTAIL.n3 1.03498
R24 VTAIL.n6 VTAIL.n5 1.03498
R25 VTAIL.n2 VTAIL.n1 1.03498
R26 VTAIL VTAIL.n0 0.575931
R27 VTAIL.n5 VTAIL.n4 0.470328
R28 VTAIL.n1 VTAIL.n0 0.470328
R29 VTAIL VTAIL.n7 0.459552
R30 B.n254 B.n253 585
R31 B.n255 B.n58 585
R32 B.n257 B.n256 585
R33 B.n259 B.n57 585
R34 B.n262 B.n261 585
R35 B.n263 B.n56 585
R36 B.n265 B.n264 585
R37 B.n267 B.n55 585
R38 B.n269 B.n268 585
R39 B.n271 B.n270 585
R40 B.n274 B.n273 585
R41 B.n275 B.n50 585
R42 B.n277 B.n276 585
R43 B.n279 B.n49 585
R44 B.n282 B.n281 585
R45 B.n283 B.n48 585
R46 B.n285 B.n284 585
R47 B.n287 B.n47 585
R48 B.n289 B.n288 585
R49 B.n291 B.n290 585
R50 B.n294 B.n293 585
R51 B.n295 B.n42 585
R52 B.n297 B.n296 585
R53 B.n299 B.n41 585
R54 B.n302 B.n301 585
R55 B.n303 B.n40 585
R56 B.n305 B.n304 585
R57 B.n307 B.n39 585
R58 B.n310 B.n309 585
R59 B.n311 B.n38 585
R60 B.n251 B.n36 585
R61 B.n314 B.n36 585
R62 B.n250 B.n35 585
R63 B.n315 B.n35 585
R64 B.n249 B.n34 585
R65 B.n316 B.n34 585
R66 B.n248 B.n247 585
R67 B.n247 B.n30 585
R68 B.n246 B.n29 585
R69 B.n322 B.n29 585
R70 B.n245 B.n28 585
R71 B.n323 B.n28 585
R72 B.n244 B.n27 585
R73 B.n324 B.n27 585
R74 B.n243 B.n242 585
R75 B.n242 B.n23 585
R76 B.n241 B.n22 585
R77 B.n330 B.n22 585
R78 B.n240 B.n21 585
R79 B.n331 B.n21 585
R80 B.n239 B.n20 585
R81 B.n332 B.n20 585
R82 B.n238 B.n237 585
R83 B.n237 B.n19 585
R84 B.n236 B.n15 585
R85 B.n338 B.n15 585
R86 B.n235 B.n14 585
R87 B.n339 B.n14 585
R88 B.n234 B.n13 585
R89 B.n340 B.n13 585
R90 B.n233 B.n232 585
R91 B.n232 B.n12 585
R92 B.n231 B.n230 585
R93 B.n231 B.n8 585
R94 B.n229 B.n7 585
R95 B.n347 B.n7 585
R96 B.n228 B.n6 585
R97 B.n348 B.n6 585
R98 B.n227 B.n5 585
R99 B.n349 B.n5 585
R100 B.n226 B.n225 585
R101 B.n225 B.n4 585
R102 B.n224 B.n59 585
R103 B.n224 B.n223 585
R104 B.n213 B.n60 585
R105 B.n216 B.n60 585
R106 B.n215 B.n214 585
R107 B.n217 B.n215 585
R108 B.n212 B.n65 585
R109 B.n65 B.n64 585
R110 B.n211 B.n210 585
R111 B.n210 B.n209 585
R112 B.n67 B.n66 585
R113 B.n202 B.n67 585
R114 B.n201 B.n200 585
R115 B.n203 B.n201 585
R116 B.n199 B.n72 585
R117 B.n72 B.n71 585
R118 B.n198 B.n197 585
R119 B.n197 B.n196 585
R120 B.n74 B.n73 585
R121 B.n75 B.n74 585
R122 B.n189 B.n188 585
R123 B.n190 B.n189 585
R124 B.n187 B.n80 585
R125 B.n80 B.n79 585
R126 B.n186 B.n185 585
R127 B.n185 B.n184 585
R128 B.n82 B.n81 585
R129 B.n83 B.n82 585
R130 B.n177 B.n176 585
R131 B.n178 B.n177 585
R132 B.n175 B.n88 585
R133 B.n88 B.n87 585
R134 B.n174 B.n173 585
R135 B.n173 B.n172 585
R136 B.n169 B.n92 585
R137 B.n168 B.n167 585
R138 B.n165 B.n93 585
R139 B.n165 B.n91 585
R140 B.n164 B.n163 585
R141 B.n162 B.n161 585
R142 B.n160 B.n95 585
R143 B.n158 B.n157 585
R144 B.n156 B.n96 585
R145 B.n155 B.n154 585
R146 B.n152 B.n97 585
R147 B.n150 B.n149 585
R148 B.n148 B.n98 585
R149 B.n147 B.n146 585
R150 B.n144 B.n102 585
R151 B.n142 B.n141 585
R152 B.n140 B.n103 585
R153 B.n139 B.n138 585
R154 B.n136 B.n104 585
R155 B.n134 B.n133 585
R156 B.n132 B.n105 585
R157 B.n130 B.n129 585
R158 B.n127 B.n108 585
R159 B.n125 B.n124 585
R160 B.n123 B.n109 585
R161 B.n122 B.n121 585
R162 B.n119 B.n110 585
R163 B.n117 B.n116 585
R164 B.n115 B.n111 585
R165 B.n114 B.n113 585
R166 B.n90 B.n89 585
R167 B.n91 B.n90 585
R168 B.n171 B.n170 585
R169 B.n172 B.n171 585
R170 B.n86 B.n85 585
R171 B.n87 B.n86 585
R172 B.n180 B.n179 585
R173 B.n179 B.n178 585
R174 B.n181 B.n84 585
R175 B.n84 B.n83 585
R176 B.n183 B.n182 585
R177 B.n184 B.n183 585
R178 B.n78 B.n77 585
R179 B.n79 B.n78 585
R180 B.n192 B.n191 585
R181 B.n191 B.n190 585
R182 B.n193 B.n76 585
R183 B.n76 B.n75 585
R184 B.n195 B.n194 585
R185 B.n196 B.n195 585
R186 B.n70 B.n69 585
R187 B.n71 B.n70 585
R188 B.n205 B.n204 585
R189 B.n204 B.n203 585
R190 B.n206 B.n68 585
R191 B.n202 B.n68 585
R192 B.n208 B.n207 585
R193 B.n209 B.n208 585
R194 B.n63 B.n62 585
R195 B.n64 B.n63 585
R196 B.n219 B.n218 585
R197 B.n218 B.n217 585
R198 B.n220 B.n61 585
R199 B.n216 B.n61 585
R200 B.n222 B.n221 585
R201 B.n223 B.n222 585
R202 B.n3 B.n0 585
R203 B.n4 B.n3 585
R204 B.n346 B.n1 585
R205 B.n347 B.n346 585
R206 B.n345 B.n344 585
R207 B.n345 B.n8 585
R208 B.n343 B.n9 585
R209 B.n12 B.n9 585
R210 B.n342 B.n341 585
R211 B.n341 B.n340 585
R212 B.n11 B.n10 585
R213 B.n339 B.n11 585
R214 B.n337 B.n336 585
R215 B.n338 B.n337 585
R216 B.n335 B.n16 585
R217 B.n19 B.n16 585
R218 B.n334 B.n333 585
R219 B.n333 B.n332 585
R220 B.n18 B.n17 585
R221 B.n331 B.n18 585
R222 B.n329 B.n328 585
R223 B.n330 B.n329 585
R224 B.n327 B.n24 585
R225 B.n24 B.n23 585
R226 B.n326 B.n325 585
R227 B.n325 B.n324 585
R228 B.n26 B.n25 585
R229 B.n323 B.n26 585
R230 B.n321 B.n320 585
R231 B.n322 B.n321 585
R232 B.n319 B.n31 585
R233 B.n31 B.n30 585
R234 B.n318 B.n317 585
R235 B.n317 B.n316 585
R236 B.n33 B.n32 585
R237 B.n315 B.n33 585
R238 B.n313 B.n312 585
R239 B.n314 B.n313 585
R240 B.n350 B.n349 585
R241 B.n348 B.n2 585
R242 B.n313 B.n38 516.524
R243 B.n253 B.n36 516.524
R244 B.n173 B.n90 516.524
R245 B.n171 B.n92 516.524
R246 B.n252 B.n37 256.663
R247 B.n258 B.n37 256.663
R248 B.n260 B.n37 256.663
R249 B.n266 B.n37 256.663
R250 B.n54 B.n37 256.663
R251 B.n272 B.n37 256.663
R252 B.n278 B.n37 256.663
R253 B.n280 B.n37 256.663
R254 B.n286 B.n37 256.663
R255 B.n46 B.n37 256.663
R256 B.n292 B.n37 256.663
R257 B.n298 B.n37 256.663
R258 B.n300 B.n37 256.663
R259 B.n306 B.n37 256.663
R260 B.n308 B.n37 256.663
R261 B.n166 B.n91 256.663
R262 B.n94 B.n91 256.663
R263 B.n159 B.n91 256.663
R264 B.n153 B.n91 256.663
R265 B.n151 B.n91 256.663
R266 B.n145 B.n91 256.663
R267 B.n143 B.n91 256.663
R268 B.n137 B.n91 256.663
R269 B.n135 B.n91 256.663
R270 B.n128 B.n91 256.663
R271 B.n126 B.n91 256.663
R272 B.n120 B.n91 256.663
R273 B.n118 B.n91 256.663
R274 B.n112 B.n91 256.663
R275 B.n352 B.n351 256.663
R276 B.n43 B.t4 237.69
R277 B.n51 B.t12 237.69
R278 B.n106 B.t8 237.69
R279 B.n99 B.t15 237.69
R280 B.n172 B.n91 229.552
R281 B.n314 B.n37 229.552
R282 B.n43 B.t6 173.257
R283 B.n51 B.t13 173.257
R284 B.n106 B.t11 173.257
R285 B.n99 B.t17 173.257
R286 B.n309 B.n307 163.367
R287 B.n305 B.n40 163.367
R288 B.n301 B.n299 163.367
R289 B.n297 B.n42 163.367
R290 B.n293 B.n291 163.367
R291 B.n288 B.n287 163.367
R292 B.n285 B.n48 163.367
R293 B.n281 B.n279 163.367
R294 B.n277 B.n50 163.367
R295 B.n273 B.n271 163.367
R296 B.n268 B.n267 163.367
R297 B.n265 B.n56 163.367
R298 B.n261 B.n259 163.367
R299 B.n257 B.n58 163.367
R300 B.n173 B.n88 163.367
R301 B.n177 B.n88 163.367
R302 B.n177 B.n82 163.367
R303 B.n185 B.n82 163.367
R304 B.n185 B.n80 163.367
R305 B.n189 B.n80 163.367
R306 B.n189 B.n74 163.367
R307 B.n197 B.n74 163.367
R308 B.n197 B.n72 163.367
R309 B.n201 B.n72 163.367
R310 B.n201 B.n67 163.367
R311 B.n210 B.n67 163.367
R312 B.n210 B.n65 163.367
R313 B.n215 B.n65 163.367
R314 B.n215 B.n60 163.367
R315 B.n224 B.n60 163.367
R316 B.n225 B.n224 163.367
R317 B.n225 B.n5 163.367
R318 B.n6 B.n5 163.367
R319 B.n7 B.n6 163.367
R320 B.n231 B.n7 163.367
R321 B.n232 B.n231 163.367
R322 B.n232 B.n13 163.367
R323 B.n14 B.n13 163.367
R324 B.n15 B.n14 163.367
R325 B.n237 B.n15 163.367
R326 B.n237 B.n20 163.367
R327 B.n21 B.n20 163.367
R328 B.n22 B.n21 163.367
R329 B.n242 B.n22 163.367
R330 B.n242 B.n27 163.367
R331 B.n28 B.n27 163.367
R332 B.n29 B.n28 163.367
R333 B.n247 B.n29 163.367
R334 B.n247 B.n34 163.367
R335 B.n35 B.n34 163.367
R336 B.n36 B.n35 163.367
R337 B.n167 B.n165 163.367
R338 B.n165 B.n164 163.367
R339 B.n161 B.n160 163.367
R340 B.n158 B.n96 163.367
R341 B.n154 B.n152 163.367
R342 B.n150 B.n98 163.367
R343 B.n146 B.n144 163.367
R344 B.n142 B.n103 163.367
R345 B.n138 B.n136 163.367
R346 B.n134 B.n105 163.367
R347 B.n129 B.n127 163.367
R348 B.n125 B.n109 163.367
R349 B.n121 B.n119 163.367
R350 B.n117 B.n111 163.367
R351 B.n113 B.n90 163.367
R352 B.n171 B.n86 163.367
R353 B.n179 B.n86 163.367
R354 B.n179 B.n84 163.367
R355 B.n183 B.n84 163.367
R356 B.n183 B.n78 163.367
R357 B.n191 B.n78 163.367
R358 B.n191 B.n76 163.367
R359 B.n195 B.n76 163.367
R360 B.n195 B.n70 163.367
R361 B.n204 B.n70 163.367
R362 B.n204 B.n68 163.367
R363 B.n208 B.n68 163.367
R364 B.n208 B.n63 163.367
R365 B.n218 B.n63 163.367
R366 B.n218 B.n61 163.367
R367 B.n222 B.n61 163.367
R368 B.n222 B.n3 163.367
R369 B.n350 B.n3 163.367
R370 B.n346 B.n2 163.367
R371 B.n346 B.n345 163.367
R372 B.n345 B.n9 163.367
R373 B.n341 B.n9 163.367
R374 B.n341 B.n11 163.367
R375 B.n337 B.n11 163.367
R376 B.n337 B.n16 163.367
R377 B.n333 B.n16 163.367
R378 B.n333 B.n18 163.367
R379 B.n329 B.n18 163.367
R380 B.n329 B.n24 163.367
R381 B.n325 B.n24 163.367
R382 B.n325 B.n26 163.367
R383 B.n321 B.n26 163.367
R384 B.n321 B.n31 163.367
R385 B.n317 B.n31 163.367
R386 B.n317 B.n33 163.367
R387 B.n313 B.n33 163.367
R388 B.n44 B.t7 149.984
R389 B.n52 B.t14 149.984
R390 B.n107 B.t10 149.984
R391 B.n100 B.t16 149.984
R392 B.n172 B.n87 113.939
R393 B.n178 B.n87 113.939
R394 B.n178 B.n83 113.939
R395 B.n184 B.n83 113.939
R396 B.n190 B.n79 113.939
R397 B.n190 B.n75 113.939
R398 B.n196 B.n75 113.939
R399 B.n196 B.n71 113.939
R400 B.n203 B.n71 113.939
R401 B.n203 B.n202 113.939
R402 B.n209 B.n64 113.939
R403 B.n217 B.n64 113.939
R404 B.n217 B.n216 113.939
R405 B.n223 B.n4 113.939
R406 B.n349 B.n4 113.939
R407 B.n349 B.n348 113.939
R408 B.n348 B.n347 113.939
R409 B.n347 B.n8 113.939
R410 B.n340 B.n12 113.939
R411 B.n340 B.n339 113.939
R412 B.n339 B.n338 113.939
R413 B.n332 B.n19 113.939
R414 B.n332 B.n331 113.939
R415 B.n331 B.n330 113.939
R416 B.n330 B.n23 113.939
R417 B.n324 B.n23 113.939
R418 B.n324 B.n323 113.939
R419 B.n322 B.n30 113.939
R420 B.n316 B.n30 113.939
R421 B.n316 B.n315 113.939
R422 B.n315 B.n314 113.939
R423 B.n184 B.t9 98.8581
R424 B.n223 B.t1 98.8581
R425 B.t2 B.n8 98.8581
R426 B.t5 B.n322 98.8581
R427 B.n308 B.n38 71.676
R428 B.n307 B.n306 71.676
R429 B.n300 B.n40 71.676
R430 B.n299 B.n298 71.676
R431 B.n292 B.n42 71.676
R432 B.n291 B.n46 71.676
R433 B.n287 B.n286 71.676
R434 B.n280 B.n48 71.676
R435 B.n279 B.n278 71.676
R436 B.n272 B.n50 71.676
R437 B.n271 B.n54 71.676
R438 B.n267 B.n266 71.676
R439 B.n260 B.n56 71.676
R440 B.n259 B.n258 71.676
R441 B.n252 B.n58 71.676
R442 B.n253 B.n252 71.676
R443 B.n258 B.n257 71.676
R444 B.n261 B.n260 71.676
R445 B.n266 B.n265 71.676
R446 B.n268 B.n54 71.676
R447 B.n273 B.n272 71.676
R448 B.n278 B.n277 71.676
R449 B.n281 B.n280 71.676
R450 B.n286 B.n285 71.676
R451 B.n288 B.n46 71.676
R452 B.n293 B.n292 71.676
R453 B.n298 B.n297 71.676
R454 B.n301 B.n300 71.676
R455 B.n306 B.n305 71.676
R456 B.n309 B.n308 71.676
R457 B.n166 B.n92 71.676
R458 B.n164 B.n94 71.676
R459 B.n160 B.n159 71.676
R460 B.n153 B.n96 71.676
R461 B.n152 B.n151 71.676
R462 B.n145 B.n98 71.676
R463 B.n144 B.n143 71.676
R464 B.n137 B.n103 71.676
R465 B.n136 B.n135 71.676
R466 B.n128 B.n105 71.676
R467 B.n127 B.n126 71.676
R468 B.n120 B.n109 71.676
R469 B.n119 B.n118 71.676
R470 B.n112 B.n111 71.676
R471 B.n167 B.n166 71.676
R472 B.n161 B.n94 71.676
R473 B.n159 B.n158 71.676
R474 B.n154 B.n153 71.676
R475 B.n151 B.n150 71.676
R476 B.n146 B.n145 71.676
R477 B.n143 B.n142 71.676
R478 B.n138 B.n137 71.676
R479 B.n135 B.n134 71.676
R480 B.n129 B.n128 71.676
R481 B.n126 B.n125 71.676
R482 B.n121 B.n120 71.676
R483 B.n118 B.n117 71.676
R484 B.n113 B.n112 71.676
R485 B.n351 B.n350 71.676
R486 B.n351 B.n2 71.676
R487 B.n202 B.t3 68.6981
R488 B.n19 B.t0 68.6981
R489 B.n45 B.n44 59.5399
R490 B.n53 B.n52 59.5399
R491 B.n131 B.n107 59.5399
R492 B.n101 B.n100 59.5399
R493 B.n209 B.t3 45.2404
R494 B.n338 B.t0 45.2404
R495 B.n170 B.n169 33.5615
R496 B.n174 B.n89 33.5615
R497 B.n254 B.n251 33.5615
R498 B.n312 B.n311 33.5615
R499 B.n44 B.n43 23.2732
R500 B.n52 B.n51 23.2732
R501 B.n107 B.n106 23.2732
R502 B.n100 B.n99 23.2732
R503 B B.n352 18.0485
R504 B.t9 B.n79 15.0805
R505 B.n216 B.t1 15.0805
R506 B.n12 B.t2 15.0805
R507 B.n323 B.t5 15.0805
R508 B.n170 B.n85 10.6151
R509 B.n180 B.n85 10.6151
R510 B.n181 B.n180 10.6151
R511 B.n182 B.n181 10.6151
R512 B.n182 B.n77 10.6151
R513 B.n192 B.n77 10.6151
R514 B.n193 B.n192 10.6151
R515 B.n194 B.n193 10.6151
R516 B.n194 B.n69 10.6151
R517 B.n205 B.n69 10.6151
R518 B.n206 B.n205 10.6151
R519 B.n207 B.n206 10.6151
R520 B.n207 B.n62 10.6151
R521 B.n219 B.n62 10.6151
R522 B.n220 B.n219 10.6151
R523 B.n221 B.n220 10.6151
R524 B.n221 B.n0 10.6151
R525 B.n169 B.n168 10.6151
R526 B.n168 B.n93 10.6151
R527 B.n163 B.n93 10.6151
R528 B.n163 B.n162 10.6151
R529 B.n162 B.n95 10.6151
R530 B.n157 B.n95 10.6151
R531 B.n157 B.n156 10.6151
R532 B.n156 B.n155 10.6151
R533 B.n155 B.n97 10.6151
R534 B.n149 B.n148 10.6151
R535 B.n148 B.n147 10.6151
R536 B.n147 B.n102 10.6151
R537 B.n141 B.n102 10.6151
R538 B.n141 B.n140 10.6151
R539 B.n140 B.n139 10.6151
R540 B.n139 B.n104 10.6151
R541 B.n133 B.n104 10.6151
R542 B.n133 B.n132 10.6151
R543 B.n130 B.n108 10.6151
R544 B.n124 B.n108 10.6151
R545 B.n124 B.n123 10.6151
R546 B.n123 B.n122 10.6151
R547 B.n122 B.n110 10.6151
R548 B.n116 B.n110 10.6151
R549 B.n116 B.n115 10.6151
R550 B.n115 B.n114 10.6151
R551 B.n114 B.n89 10.6151
R552 B.n175 B.n174 10.6151
R553 B.n176 B.n175 10.6151
R554 B.n176 B.n81 10.6151
R555 B.n186 B.n81 10.6151
R556 B.n187 B.n186 10.6151
R557 B.n188 B.n187 10.6151
R558 B.n188 B.n73 10.6151
R559 B.n198 B.n73 10.6151
R560 B.n199 B.n198 10.6151
R561 B.n200 B.n199 10.6151
R562 B.n200 B.n66 10.6151
R563 B.n211 B.n66 10.6151
R564 B.n212 B.n211 10.6151
R565 B.n214 B.n212 10.6151
R566 B.n214 B.n213 10.6151
R567 B.n213 B.n59 10.6151
R568 B.n226 B.n59 10.6151
R569 B.n227 B.n226 10.6151
R570 B.n228 B.n227 10.6151
R571 B.n229 B.n228 10.6151
R572 B.n230 B.n229 10.6151
R573 B.n233 B.n230 10.6151
R574 B.n234 B.n233 10.6151
R575 B.n235 B.n234 10.6151
R576 B.n236 B.n235 10.6151
R577 B.n238 B.n236 10.6151
R578 B.n239 B.n238 10.6151
R579 B.n240 B.n239 10.6151
R580 B.n241 B.n240 10.6151
R581 B.n243 B.n241 10.6151
R582 B.n244 B.n243 10.6151
R583 B.n245 B.n244 10.6151
R584 B.n246 B.n245 10.6151
R585 B.n248 B.n246 10.6151
R586 B.n249 B.n248 10.6151
R587 B.n250 B.n249 10.6151
R588 B.n251 B.n250 10.6151
R589 B.n344 B.n1 10.6151
R590 B.n344 B.n343 10.6151
R591 B.n343 B.n342 10.6151
R592 B.n342 B.n10 10.6151
R593 B.n336 B.n10 10.6151
R594 B.n336 B.n335 10.6151
R595 B.n335 B.n334 10.6151
R596 B.n334 B.n17 10.6151
R597 B.n328 B.n17 10.6151
R598 B.n328 B.n327 10.6151
R599 B.n327 B.n326 10.6151
R600 B.n326 B.n25 10.6151
R601 B.n320 B.n25 10.6151
R602 B.n320 B.n319 10.6151
R603 B.n319 B.n318 10.6151
R604 B.n318 B.n32 10.6151
R605 B.n312 B.n32 10.6151
R606 B.n311 B.n310 10.6151
R607 B.n310 B.n39 10.6151
R608 B.n304 B.n39 10.6151
R609 B.n304 B.n303 10.6151
R610 B.n303 B.n302 10.6151
R611 B.n302 B.n41 10.6151
R612 B.n296 B.n41 10.6151
R613 B.n296 B.n295 10.6151
R614 B.n295 B.n294 10.6151
R615 B.n290 B.n289 10.6151
R616 B.n289 B.n47 10.6151
R617 B.n284 B.n47 10.6151
R618 B.n284 B.n283 10.6151
R619 B.n283 B.n282 10.6151
R620 B.n282 B.n49 10.6151
R621 B.n276 B.n49 10.6151
R622 B.n276 B.n275 10.6151
R623 B.n275 B.n274 10.6151
R624 B.n270 B.n269 10.6151
R625 B.n269 B.n55 10.6151
R626 B.n264 B.n55 10.6151
R627 B.n264 B.n263 10.6151
R628 B.n263 B.n262 10.6151
R629 B.n262 B.n57 10.6151
R630 B.n256 B.n57 10.6151
R631 B.n256 B.n255 10.6151
R632 B.n255 B.n254 10.6151
R633 B.n101 B.n97 9.36635
R634 B.n131 B.n130 9.36635
R635 B.n294 B.n45 9.36635
R636 B.n270 B.n53 9.36635
R637 B.n352 B.n0 8.11757
R638 B.n352 B.n1 8.11757
R639 B.n149 B.n101 1.24928
R640 B.n132 B.n131 1.24928
R641 B.n290 B.n45 1.24928
R642 B.n274 B.n53 1.24928
R643 VP.n6 VP.n5 161.3
R644 VP.n4 VP.n0 161.3
R645 VP.n3 VP.n2 161.3
R646 VP.n1 VP.t1 102.162
R647 VP.n1 VP.t2 102.112
R648 VP.n3 VP.t0 81.1649
R649 VP.n5 VP.t3 81.1649
R650 VP.n2 VP.n1 77.6015
R651 VP.n4 VP.n3 24.1005
R652 VP.n5 VP.n4 24.1005
R653 VP.n2 VP.n0 0.189894
R654 VP.n6 VP.n0 0.189894
R655 VP VP.n6 0.0516364
R656 VDD1 VDD1.n1 175.078
R657 VDD1 VDD1.n0 146.681
R658 VDD1.n0 VDD1.t2 15.3493
R659 VDD1.n0 VDD1.t1 15.3493
R660 VDD1.n1 VDD1.t3 15.3493
R661 VDD1.n1 VDD1.t0 15.3493
C0 VDD2 VDD1 0.606243f
C1 VDD2 VP 0.291548f
C2 VDD2 VN 0.641046f
C3 VDD2 VTAIL 2.11369f
C4 VDD1 VP 0.777514f
C5 VDD1 VN 0.153835f
C6 VP VN 2.96607f
C7 VDD1 VTAIL 2.07108f
C8 VTAIL VP 0.858212f
C9 VTAIL VN 0.844105f
C10 VDD2 B 1.923289f
C11 VDD1 B 3.74022f
C12 VTAIL B 2.544327f
C13 VN B 6.07742f
C14 VP B 4.341271f
C15 VDD1.t2 B 0.020243f
C16 VDD1.t1 B 0.020243f
C17 VDD1.n0 B 0.101456f
C18 VDD1.t3 B 0.020243f
C19 VDD1.t0 B 0.020243f
C20 VDD1.n1 B 0.211108f
C21 VP.n0 B 0.034922f
C22 VP.t2 B 0.150316f
C23 VP.t1 B 0.15039f
C24 VP.n1 B 0.602276f
C25 VP.n2 B 1.53845f
C26 VP.t0 B 0.128002f
C27 VP.n3 B 0.106263f
C28 VP.n4 B 0.007925f
C29 VP.t3 B 0.128002f
C30 VP.n5 B 0.106263f
C31 VP.n6 B 0.027063f
C32 VTAIL.t3 B 0.111123f
C33 VTAIL.n0 B 0.208186f
C34 VTAIL.t5 B 0.111123f
C35 VTAIL.n1 B 0.235915f
C36 VTAIL.t7 B 0.111123f
C37 VTAIL.n2 B 0.59184f
C38 VTAIL.t4 B 0.111123f
C39 VTAIL.n3 B 0.59184f
C40 VTAIL.t2 B 0.111123f
C41 VTAIL.n4 B 0.235915f
C42 VTAIL.t6 B 0.111123f
C43 VTAIL.n5 B 0.235915f
C44 VTAIL.t0 B 0.111123f
C45 VTAIL.n6 B 0.59184f
C46 VTAIL.t1 B 0.111123f
C47 VTAIL.n7 B 0.557082f
C48 VDD2.t1 B 0.020976f
C49 VDD2.t0 B 0.020976f
C50 VDD2.n0 B 0.210181f
C51 VDD2.t3 B 0.020976f
C52 VDD2.t2 B 0.020976f
C53 VDD2.n1 B 0.105037f
C54 VDD2.n2 B 1.62786f
C55 VN.t1 B 0.147969f
C56 VN.t3 B 0.147896f
C57 VN.n0 B 0.173298f
C58 VN.t2 B 0.147969f
C59 VN.t0 B 0.147896f
C60 VN.n1 B 0.60516f
.ends

