* NGSPICE file created from diff_pair_sample_0462.ext - technology: sky130A

.subckt diff_pair_sample_0462 VTAIL VN VP B VDD2 VDD1
X0 B.t23 B.t21 B.t22 B.t15 sky130_fd_pr__nfet_01v8 ad=3.1122 pd=16.74 as=0 ps=0 w=7.98 l=1.04
X1 VTAIL.t18 VN.t0 VDD2.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=1.3167 pd=8.31 as=1.3167 ps=8.31 w=7.98 l=1.04
X2 VTAIL.t0 VP.t0 VDD1.t9 B.t2 sky130_fd_pr__nfet_01v8 ad=1.3167 pd=8.31 as=1.3167 ps=8.31 w=7.98 l=1.04
X3 B.t20 B.t18 B.t19 B.t11 sky130_fd_pr__nfet_01v8 ad=3.1122 pd=16.74 as=0 ps=0 w=7.98 l=1.04
X4 VTAIL.t6 VP.t1 VDD1.t8 B.t0 sky130_fd_pr__nfet_01v8 ad=1.3167 pd=8.31 as=1.3167 ps=8.31 w=7.98 l=1.04
X5 VDD1.t7 VP.t2 VTAIL.t5 B.t7 sky130_fd_pr__nfet_01v8 ad=3.1122 pd=16.74 as=1.3167 ps=8.31 w=7.98 l=1.04
X6 VDD1.t6 VP.t3 VTAIL.t19 B.t1 sky130_fd_pr__nfet_01v8 ad=1.3167 pd=8.31 as=1.3167 ps=8.31 w=7.98 l=1.04
X7 VTAIL.t17 VN.t1 VDD2.t7 B.t0 sky130_fd_pr__nfet_01v8 ad=1.3167 pd=8.31 as=1.3167 ps=8.31 w=7.98 l=1.04
X8 VDD1.t5 VP.t4 VTAIL.t7 B.t9 sky130_fd_pr__nfet_01v8 ad=1.3167 pd=8.31 as=3.1122 ps=16.74 w=7.98 l=1.04
X9 VDD1.t4 VP.t5 VTAIL.t8 B.t5 sky130_fd_pr__nfet_01v8 ad=3.1122 pd=16.74 as=1.3167 ps=8.31 w=7.98 l=1.04
X10 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=3.1122 pd=16.74 as=0 ps=0 w=7.98 l=1.04
X11 VDD2.t4 VN.t2 VTAIL.t16 B.t6 sky130_fd_pr__nfet_01v8 ad=1.3167 pd=8.31 as=1.3167 ps=8.31 w=7.98 l=1.04
X12 VTAIL.t15 VN.t3 VDD2.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=1.3167 pd=8.31 as=1.3167 ps=8.31 w=7.98 l=1.04
X13 VDD2.t8 VN.t4 VTAIL.t14 B.t1 sky130_fd_pr__nfet_01v8 ad=1.3167 pd=8.31 as=1.3167 ps=8.31 w=7.98 l=1.04
X14 VDD2.t1 VN.t5 VTAIL.t13 B.t3 sky130_fd_pr__nfet_01v8 ad=1.3167 pd=8.31 as=3.1122 ps=16.74 w=7.98 l=1.04
X15 VTAIL.t12 VN.t6 VDD2.t9 B.t8 sky130_fd_pr__nfet_01v8 ad=1.3167 pd=8.31 as=1.3167 ps=8.31 w=7.98 l=1.04
X16 VDD2.t3 VN.t7 VTAIL.t11 B.t5 sky130_fd_pr__nfet_01v8 ad=3.1122 pd=16.74 as=1.3167 ps=8.31 w=7.98 l=1.04
X17 VTAIL.t4 VP.t6 VDD1.t3 B.t4 sky130_fd_pr__nfet_01v8 ad=1.3167 pd=8.31 as=1.3167 ps=8.31 w=7.98 l=1.04
X18 VDD2.t2 VN.t8 VTAIL.t10 B.t7 sky130_fd_pr__nfet_01v8 ad=3.1122 pd=16.74 as=1.3167 ps=8.31 w=7.98 l=1.04
X19 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=3.1122 pd=16.74 as=0 ps=0 w=7.98 l=1.04
X20 VDD2.t0 VN.t9 VTAIL.t9 B.t9 sky130_fd_pr__nfet_01v8 ad=1.3167 pd=8.31 as=3.1122 ps=16.74 w=7.98 l=1.04
X21 VDD1.t2 VP.t7 VTAIL.t2 B.t6 sky130_fd_pr__nfet_01v8 ad=1.3167 pd=8.31 as=1.3167 ps=8.31 w=7.98 l=1.04
X22 VTAIL.t3 VP.t8 VDD1.t1 B.t8 sky130_fd_pr__nfet_01v8 ad=1.3167 pd=8.31 as=1.3167 ps=8.31 w=7.98 l=1.04
X23 VDD1.t0 VP.t9 VTAIL.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=1.3167 pd=8.31 as=3.1122 ps=16.74 w=7.98 l=1.04
R0 B.n617 B.n616 585
R1 B.n618 B.n617 585
R2 B.n235 B.n96 585
R3 B.n234 B.n233 585
R4 B.n232 B.n231 585
R5 B.n230 B.n229 585
R6 B.n228 B.n227 585
R7 B.n226 B.n225 585
R8 B.n224 B.n223 585
R9 B.n222 B.n221 585
R10 B.n220 B.n219 585
R11 B.n218 B.n217 585
R12 B.n216 B.n215 585
R13 B.n214 B.n213 585
R14 B.n212 B.n211 585
R15 B.n210 B.n209 585
R16 B.n208 B.n207 585
R17 B.n206 B.n205 585
R18 B.n204 B.n203 585
R19 B.n202 B.n201 585
R20 B.n200 B.n199 585
R21 B.n198 B.n197 585
R22 B.n196 B.n195 585
R23 B.n194 B.n193 585
R24 B.n192 B.n191 585
R25 B.n190 B.n189 585
R26 B.n188 B.n187 585
R27 B.n186 B.n185 585
R28 B.n184 B.n183 585
R29 B.n182 B.n181 585
R30 B.n180 B.n179 585
R31 B.n177 B.n176 585
R32 B.n175 B.n174 585
R33 B.n173 B.n172 585
R34 B.n171 B.n170 585
R35 B.n169 B.n168 585
R36 B.n167 B.n166 585
R37 B.n165 B.n164 585
R38 B.n163 B.n162 585
R39 B.n161 B.n160 585
R40 B.n159 B.n158 585
R41 B.n157 B.n156 585
R42 B.n155 B.n154 585
R43 B.n153 B.n152 585
R44 B.n151 B.n150 585
R45 B.n149 B.n148 585
R46 B.n147 B.n146 585
R47 B.n145 B.n144 585
R48 B.n143 B.n142 585
R49 B.n141 B.n140 585
R50 B.n139 B.n138 585
R51 B.n137 B.n136 585
R52 B.n135 B.n134 585
R53 B.n133 B.n132 585
R54 B.n131 B.n130 585
R55 B.n129 B.n128 585
R56 B.n127 B.n126 585
R57 B.n125 B.n124 585
R58 B.n123 B.n122 585
R59 B.n121 B.n120 585
R60 B.n119 B.n118 585
R61 B.n117 B.n116 585
R62 B.n115 B.n114 585
R63 B.n113 B.n112 585
R64 B.n111 B.n110 585
R65 B.n109 B.n108 585
R66 B.n107 B.n106 585
R67 B.n105 B.n104 585
R68 B.n103 B.n102 585
R69 B.n60 B.n59 585
R70 B.n615 B.n61 585
R71 B.n619 B.n61 585
R72 B.n614 B.n613 585
R73 B.n613 B.n57 585
R74 B.n612 B.n56 585
R75 B.n625 B.n56 585
R76 B.n611 B.n55 585
R77 B.n626 B.n55 585
R78 B.n610 B.n54 585
R79 B.n627 B.n54 585
R80 B.n609 B.n608 585
R81 B.n608 B.n53 585
R82 B.n607 B.n49 585
R83 B.n633 B.n49 585
R84 B.n606 B.n48 585
R85 B.n634 B.n48 585
R86 B.n605 B.n47 585
R87 B.n635 B.n47 585
R88 B.n604 B.n603 585
R89 B.n603 B.n43 585
R90 B.n602 B.n42 585
R91 B.n641 B.n42 585
R92 B.n601 B.n41 585
R93 B.n642 B.n41 585
R94 B.n600 B.n40 585
R95 B.n643 B.n40 585
R96 B.n599 B.n598 585
R97 B.n598 B.n36 585
R98 B.n597 B.n35 585
R99 B.n649 B.n35 585
R100 B.n596 B.n34 585
R101 B.n650 B.n34 585
R102 B.n595 B.n33 585
R103 B.n651 B.n33 585
R104 B.n594 B.n593 585
R105 B.n593 B.n29 585
R106 B.n592 B.n28 585
R107 B.n657 B.n28 585
R108 B.n591 B.n27 585
R109 B.n658 B.n27 585
R110 B.n590 B.n26 585
R111 B.n659 B.n26 585
R112 B.n589 B.n588 585
R113 B.n588 B.n22 585
R114 B.n587 B.n21 585
R115 B.n665 B.n21 585
R116 B.n586 B.n20 585
R117 B.n666 B.n20 585
R118 B.n585 B.n19 585
R119 B.n667 B.n19 585
R120 B.n584 B.n583 585
R121 B.n583 B.n15 585
R122 B.n582 B.n14 585
R123 B.n673 B.n14 585
R124 B.n581 B.n13 585
R125 B.n674 B.n13 585
R126 B.n580 B.n12 585
R127 B.n675 B.n12 585
R128 B.n579 B.n578 585
R129 B.n578 B.n577 585
R130 B.n576 B.n575 585
R131 B.n576 B.n8 585
R132 B.n574 B.n7 585
R133 B.n682 B.n7 585
R134 B.n573 B.n6 585
R135 B.n683 B.n6 585
R136 B.n572 B.n5 585
R137 B.n684 B.n5 585
R138 B.n571 B.n570 585
R139 B.n570 B.n4 585
R140 B.n569 B.n236 585
R141 B.n569 B.n568 585
R142 B.n559 B.n237 585
R143 B.n238 B.n237 585
R144 B.n561 B.n560 585
R145 B.n562 B.n561 585
R146 B.n558 B.n243 585
R147 B.n243 B.n242 585
R148 B.n557 B.n556 585
R149 B.n556 B.n555 585
R150 B.n245 B.n244 585
R151 B.n246 B.n245 585
R152 B.n548 B.n547 585
R153 B.n549 B.n548 585
R154 B.n546 B.n251 585
R155 B.n251 B.n250 585
R156 B.n545 B.n544 585
R157 B.n544 B.n543 585
R158 B.n253 B.n252 585
R159 B.n254 B.n253 585
R160 B.n536 B.n535 585
R161 B.n537 B.n536 585
R162 B.n534 B.n259 585
R163 B.n259 B.n258 585
R164 B.n533 B.n532 585
R165 B.n532 B.n531 585
R166 B.n261 B.n260 585
R167 B.n262 B.n261 585
R168 B.n524 B.n523 585
R169 B.n525 B.n524 585
R170 B.n522 B.n267 585
R171 B.n267 B.n266 585
R172 B.n521 B.n520 585
R173 B.n520 B.n519 585
R174 B.n269 B.n268 585
R175 B.n270 B.n269 585
R176 B.n512 B.n511 585
R177 B.n513 B.n512 585
R178 B.n510 B.n275 585
R179 B.n275 B.n274 585
R180 B.n509 B.n508 585
R181 B.n508 B.n507 585
R182 B.n277 B.n276 585
R183 B.n278 B.n277 585
R184 B.n500 B.n499 585
R185 B.n501 B.n500 585
R186 B.n498 B.n283 585
R187 B.n283 B.n282 585
R188 B.n497 B.n496 585
R189 B.n496 B.n495 585
R190 B.n285 B.n284 585
R191 B.n488 B.n285 585
R192 B.n487 B.n486 585
R193 B.n489 B.n487 585
R194 B.n485 B.n290 585
R195 B.n290 B.n289 585
R196 B.n484 B.n483 585
R197 B.n483 B.n482 585
R198 B.n292 B.n291 585
R199 B.n293 B.n292 585
R200 B.n475 B.n474 585
R201 B.n476 B.n475 585
R202 B.n296 B.n295 585
R203 B.n337 B.n335 585
R204 B.n338 B.n334 585
R205 B.n338 B.n297 585
R206 B.n341 B.n340 585
R207 B.n342 B.n333 585
R208 B.n344 B.n343 585
R209 B.n346 B.n332 585
R210 B.n349 B.n348 585
R211 B.n350 B.n331 585
R212 B.n352 B.n351 585
R213 B.n354 B.n330 585
R214 B.n357 B.n356 585
R215 B.n358 B.n329 585
R216 B.n360 B.n359 585
R217 B.n362 B.n328 585
R218 B.n365 B.n364 585
R219 B.n366 B.n327 585
R220 B.n368 B.n367 585
R221 B.n370 B.n326 585
R222 B.n373 B.n372 585
R223 B.n374 B.n325 585
R224 B.n376 B.n375 585
R225 B.n378 B.n324 585
R226 B.n381 B.n380 585
R227 B.n382 B.n323 585
R228 B.n384 B.n383 585
R229 B.n386 B.n322 585
R230 B.n389 B.n388 585
R231 B.n390 B.n321 585
R232 B.n395 B.n394 585
R233 B.n397 B.n320 585
R234 B.n400 B.n399 585
R235 B.n401 B.n319 585
R236 B.n403 B.n402 585
R237 B.n405 B.n318 585
R238 B.n408 B.n407 585
R239 B.n409 B.n317 585
R240 B.n411 B.n410 585
R241 B.n413 B.n316 585
R242 B.n416 B.n415 585
R243 B.n417 B.n312 585
R244 B.n419 B.n418 585
R245 B.n421 B.n311 585
R246 B.n424 B.n423 585
R247 B.n425 B.n310 585
R248 B.n427 B.n426 585
R249 B.n429 B.n309 585
R250 B.n432 B.n431 585
R251 B.n433 B.n308 585
R252 B.n435 B.n434 585
R253 B.n437 B.n307 585
R254 B.n440 B.n439 585
R255 B.n441 B.n306 585
R256 B.n443 B.n442 585
R257 B.n445 B.n305 585
R258 B.n448 B.n447 585
R259 B.n449 B.n304 585
R260 B.n451 B.n450 585
R261 B.n453 B.n303 585
R262 B.n456 B.n455 585
R263 B.n457 B.n302 585
R264 B.n459 B.n458 585
R265 B.n461 B.n301 585
R266 B.n464 B.n463 585
R267 B.n465 B.n300 585
R268 B.n467 B.n466 585
R269 B.n469 B.n299 585
R270 B.n472 B.n471 585
R271 B.n473 B.n298 585
R272 B.n478 B.n477 585
R273 B.n477 B.n476 585
R274 B.n479 B.n294 585
R275 B.n294 B.n293 585
R276 B.n481 B.n480 585
R277 B.n482 B.n481 585
R278 B.n288 B.n287 585
R279 B.n289 B.n288 585
R280 B.n491 B.n490 585
R281 B.n490 B.n489 585
R282 B.n492 B.n286 585
R283 B.n488 B.n286 585
R284 B.n494 B.n493 585
R285 B.n495 B.n494 585
R286 B.n281 B.n280 585
R287 B.n282 B.n281 585
R288 B.n503 B.n502 585
R289 B.n502 B.n501 585
R290 B.n504 B.n279 585
R291 B.n279 B.n278 585
R292 B.n506 B.n505 585
R293 B.n507 B.n506 585
R294 B.n273 B.n272 585
R295 B.n274 B.n273 585
R296 B.n515 B.n514 585
R297 B.n514 B.n513 585
R298 B.n516 B.n271 585
R299 B.n271 B.n270 585
R300 B.n518 B.n517 585
R301 B.n519 B.n518 585
R302 B.n265 B.n264 585
R303 B.n266 B.n265 585
R304 B.n527 B.n526 585
R305 B.n526 B.n525 585
R306 B.n528 B.n263 585
R307 B.n263 B.n262 585
R308 B.n530 B.n529 585
R309 B.n531 B.n530 585
R310 B.n257 B.n256 585
R311 B.n258 B.n257 585
R312 B.n539 B.n538 585
R313 B.n538 B.n537 585
R314 B.n540 B.n255 585
R315 B.n255 B.n254 585
R316 B.n542 B.n541 585
R317 B.n543 B.n542 585
R318 B.n249 B.n248 585
R319 B.n250 B.n249 585
R320 B.n551 B.n550 585
R321 B.n550 B.n549 585
R322 B.n552 B.n247 585
R323 B.n247 B.n246 585
R324 B.n554 B.n553 585
R325 B.n555 B.n554 585
R326 B.n241 B.n240 585
R327 B.n242 B.n241 585
R328 B.n564 B.n563 585
R329 B.n563 B.n562 585
R330 B.n565 B.n239 585
R331 B.n239 B.n238 585
R332 B.n567 B.n566 585
R333 B.n568 B.n567 585
R334 B.n3 B.n0 585
R335 B.n4 B.n3 585
R336 B.n681 B.n1 585
R337 B.n682 B.n681 585
R338 B.n680 B.n679 585
R339 B.n680 B.n8 585
R340 B.n678 B.n9 585
R341 B.n577 B.n9 585
R342 B.n677 B.n676 585
R343 B.n676 B.n675 585
R344 B.n11 B.n10 585
R345 B.n674 B.n11 585
R346 B.n672 B.n671 585
R347 B.n673 B.n672 585
R348 B.n670 B.n16 585
R349 B.n16 B.n15 585
R350 B.n669 B.n668 585
R351 B.n668 B.n667 585
R352 B.n18 B.n17 585
R353 B.n666 B.n18 585
R354 B.n664 B.n663 585
R355 B.n665 B.n664 585
R356 B.n662 B.n23 585
R357 B.n23 B.n22 585
R358 B.n661 B.n660 585
R359 B.n660 B.n659 585
R360 B.n25 B.n24 585
R361 B.n658 B.n25 585
R362 B.n656 B.n655 585
R363 B.n657 B.n656 585
R364 B.n654 B.n30 585
R365 B.n30 B.n29 585
R366 B.n653 B.n652 585
R367 B.n652 B.n651 585
R368 B.n32 B.n31 585
R369 B.n650 B.n32 585
R370 B.n648 B.n647 585
R371 B.n649 B.n648 585
R372 B.n646 B.n37 585
R373 B.n37 B.n36 585
R374 B.n645 B.n644 585
R375 B.n644 B.n643 585
R376 B.n39 B.n38 585
R377 B.n642 B.n39 585
R378 B.n640 B.n639 585
R379 B.n641 B.n640 585
R380 B.n638 B.n44 585
R381 B.n44 B.n43 585
R382 B.n637 B.n636 585
R383 B.n636 B.n635 585
R384 B.n46 B.n45 585
R385 B.n634 B.n46 585
R386 B.n632 B.n631 585
R387 B.n633 B.n632 585
R388 B.n630 B.n50 585
R389 B.n53 B.n50 585
R390 B.n629 B.n628 585
R391 B.n628 B.n627 585
R392 B.n52 B.n51 585
R393 B.n626 B.n52 585
R394 B.n624 B.n623 585
R395 B.n625 B.n624 585
R396 B.n622 B.n58 585
R397 B.n58 B.n57 585
R398 B.n621 B.n620 585
R399 B.n620 B.n619 585
R400 B.n685 B.n684 585
R401 B.n683 B.n2 585
R402 B.n620 B.n60 478.086
R403 B.n617 B.n61 478.086
R404 B.n475 B.n298 478.086
R405 B.n477 B.n296 478.086
R406 B.n99 B.t14 388.111
R407 B.n97 B.t21 388.111
R408 B.n313 B.t18 388.111
R409 B.n391 B.t10 388.111
R410 B.n618 B.n95 256.663
R411 B.n618 B.n94 256.663
R412 B.n618 B.n93 256.663
R413 B.n618 B.n92 256.663
R414 B.n618 B.n91 256.663
R415 B.n618 B.n90 256.663
R416 B.n618 B.n89 256.663
R417 B.n618 B.n88 256.663
R418 B.n618 B.n87 256.663
R419 B.n618 B.n86 256.663
R420 B.n618 B.n85 256.663
R421 B.n618 B.n84 256.663
R422 B.n618 B.n83 256.663
R423 B.n618 B.n82 256.663
R424 B.n618 B.n81 256.663
R425 B.n618 B.n80 256.663
R426 B.n618 B.n79 256.663
R427 B.n618 B.n78 256.663
R428 B.n618 B.n77 256.663
R429 B.n618 B.n76 256.663
R430 B.n618 B.n75 256.663
R431 B.n618 B.n74 256.663
R432 B.n618 B.n73 256.663
R433 B.n618 B.n72 256.663
R434 B.n618 B.n71 256.663
R435 B.n618 B.n70 256.663
R436 B.n618 B.n69 256.663
R437 B.n618 B.n68 256.663
R438 B.n618 B.n67 256.663
R439 B.n618 B.n66 256.663
R440 B.n618 B.n65 256.663
R441 B.n618 B.n64 256.663
R442 B.n618 B.n63 256.663
R443 B.n618 B.n62 256.663
R444 B.n336 B.n297 256.663
R445 B.n339 B.n297 256.663
R446 B.n345 B.n297 256.663
R447 B.n347 B.n297 256.663
R448 B.n353 B.n297 256.663
R449 B.n355 B.n297 256.663
R450 B.n361 B.n297 256.663
R451 B.n363 B.n297 256.663
R452 B.n369 B.n297 256.663
R453 B.n371 B.n297 256.663
R454 B.n377 B.n297 256.663
R455 B.n379 B.n297 256.663
R456 B.n385 B.n297 256.663
R457 B.n387 B.n297 256.663
R458 B.n396 B.n297 256.663
R459 B.n398 B.n297 256.663
R460 B.n404 B.n297 256.663
R461 B.n406 B.n297 256.663
R462 B.n412 B.n297 256.663
R463 B.n414 B.n297 256.663
R464 B.n420 B.n297 256.663
R465 B.n422 B.n297 256.663
R466 B.n428 B.n297 256.663
R467 B.n430 B.n297 256.663
R468 B.n436 B.n297 256.663
R469 B.n438 B.n297 256.663
R470 B.n444 B.n297 256.663
R471 B.n446 B.n297 256.663
R472 B.n452 B.n297 256.663
R473 B.n454 B.n297 256.663
R474 B.n460 B.n297 256.663
R475 B.n462 B.n297 256.663
R476 B.n468 B.n297 256.663
R477 B.n470 B.n297 256.663
R478 B.n687 B.n686 256.663
R479 B.n97 B.t22 239.472
R480 B.n313 B.t20 239.472
R481 B.n99 B.t16 239.472
R482 B.n391 B.t13 239.472
R483 B.n98 B.t23 212.904
R484 B.n314 B.t19 212.904
R485 B.n100 B.t17 212.904
R486 B.n392 B.t12 212.904
R487 B.n104 B.n103 163.367
R488 B.n108 B.n107 163.367
R489 B.n112 B.n111 163.367
R490 B.n116 B.n115 163.367
R491 B.n120 B.n119 163.367
R492 B.n124 B.n123 163.367
R493 B.n128 B.n127 163.367
R494 B.n132 B.n131 163.367
R495 B.n136 B.n135 163.367
R496 B.n140 B.n139 163.367
R497 B.n144 B.n143 163.367
R498 B.n148 B.n147 163.367
R499 B.n152 B.n151 163.367
R500 B.n156 B.n155 163.367
R501 B.n160 B.n159 163.367
R502 B.n164 B.n163 163.367
R503 B.n168 B.n167 163.367
R504 B.n172 B.n171 163.367
R505 B.n176 B.n175 163.367
R506 B.n181 B.n180 163.367
R507 B.n185 B.n184 163.367
R508 B.n189 B.n188 163.367
R509 B.n193 B.n192 163.367
R510 B.n197 B.n196 163.367
R511 B.n201 B.n200 163.367
R512 B.n205 B.n204 163.367
R513 B.n209 B.n208 163.367
R514 B.n213 B.n212 163.367
R515 B.n217 B.n216 163.367
R516 B.n221 B.n220 163.367
R517 B.n225 B.n224 163.367
R518 B.n229 B.n228 163.367
R519 B.n233 B.n232 163.367
R520 B.n617 B.n96 163.367
R521 B.n475 B.n292 163.367
R522 B.n483 B.n292 163.367
R523 B.n483 B.n290 163.367
R524 B.n487 B.n290 163.367
R525 B.n487 B.n285 163.367
R526 B.n496 B.n285 163.367
R527 B.n496 B.n283 163.367
R528 B.n500 B.n283 163.367
R529 B.n500 B.n277 163.367
R530 B.n508 B.n277 163.367
R531 B.n508 B.n275 163.367
R532 B.n512 B.n275 163.367
R533 B.n512 B.n269 163.367
R534 B.n520 B.n269 163.367
R535 B.n520 B.n267 163.367
R536 B.n524 B.n267 163.367
R537 B.n524 B.n261 163.367
R538 B.n532 B.n261 163.367
R539 B.n532 B.n259 163.367
R540 B.n536 B.n259 163.367
R541 B.n536 B.n253 163.367
R542 B.n544 B.n253 163.367
R543 B.n544 B.n251 163.367
R544 B.n548 B.n251 163.367
R545 B.n548 B.n245 163.367
R546 B.n556 B.n245 163.367
R547 B.n556 B.n243 163.367
R548 B.n561 B.n243 163.367
R549 B.n561 B.n237 163.367
R550 B.n569 B.n237 163.367
R551 B.n570 B.n569 163.367
R552 B.n570 B.n5 163.367
R553 B.n6 B.n5 163.367
R554 B.n7 B.n6 163.367
R555 B.n576 B.n7 163.367
R556 B.n578 B.n576 163.367
R557 B.n578 B.n12 163.367
R558 B.n13 B.n12 163.367
R559 B.n14 B.n13 163.367
R560 B.n583 B.n14 163.367
R561 B.n583 B.n19 163.367
R562 B.n20 B.n19 163.367
R563 B.n21 B.n20 163.367
R564 B.n588 B.n21 163.367
R565 B.n588 B.n26 163.367
R566 B.n27 B.n26 163.367
R567 B.n28 B.n27 163.367
R568 B.n593 B.n28 163.367
R569 B.n593 B.n33 163.367
R570 B.n34 B.n33 163.367
R571 B.n35 B.n34 163.367
R572 B.n598 B.n35 163.367
R573 B.n598 B.n40 163.367
R574 B.n41 B.n40 163.367
R575 B.n42 B.n41 163.367
R576 B.n603 B.n42 163.367
R577 B.n603 B.n47 163.367
R578 B.n48 B.n47 163.367
R579 B.n49 B.n48 163.367
R580 B.n608 B.n49 163.367
R581 B.n608 B.n54 163.367
R582 B.n55 B.n54 163.367
R583 B.n56 B.n55 163.367
R584 B.n613 B.n56 163.367
R585 B.n613 B.n61 163.367
R586 B.n338 B.n337 163.367
R587 B.n340 B.n338 163.367
R588 B.n344 B.n333 163.367
R589 B.n348 B.n346 163.367
R590 B.n352 B.n331 163.367
R591 B.n356 B.n354 163.367
R592 B.n360 B.n329 163.367
R593 B.n364 B.n362 163.367
R594 B.n368 B.n327 163.367
R595 B.n372 B.n370 163.367
R596 B.n376 B.n325 163.367
R597 B.n380 B.n378 163.367
R598 B.n384 B.n323 163.367
R599 B.n388 B.n386 163.367
R600 B.n395 B.n321 163.367
R601 B.n399 B.n397 163.367
R602 B.n403 B.n319 163.367
R603 B.n407 B.n405 163.367
R604 B.n411 B.n317 163.367
R605 B.n415 B.n413 163.367
R606 B.n419 B.n312 163.367
R607 B.n423 B.n421 163.367
R608 B.n427 B.n310 163.367
R609 B.n431 B.n429 163.367
R610 B.n435 B.n308 163.367
R611 B.n439 B.n437 163.367
R612 B.n443 B.n306 163.367
R613 B.n447 B.n445 163.367
R614 B.n451 B.n304 163.367
R615 B.n455 B.n453 163.367
R616 B.n459 B.n302 163.367
R617 B.n463 B.n461 163.367
R618 B.n467 B.n300 163.367
R619 B.n471 B.n469 163.367
R620 B.n477 B.n294 163.367
R621 B.n481 B.n294 163.367
R622 B.n481 B.n288 163.367
R623 B.n490 B.n288 163.367
R624 B.n490 B.n286 163.367
R625 B.n494 B.n286 163.367
R626 B.n494 B.n281 163.367
R627 B.n502 B.n281 163.367
R628 B.n502 B.n279 163.367
R629 B.n506 B.n279 163.367
R630 B.n506 B.n273 163.367
R631 B.n514 B.n273 163.367
R632 B.n514 B.n271 163.367
R633 B.n518 B.n271 163.367
R634 B.n518 B.n265 163.367
R635 B.n526 B.n265 163.367
R636 B.n526 B.n263 163.367
R637 B.n530 B.n263 163.367
R638 B.n530 B.n257 163.367
R639 B.n538 B.n257 163.367
R640 B.n538 B.n255 163.367
R641 B.n542 B.n255 163.367
R642 B.n542 B.n249 163.367
R643 B.n550 B.n249 163.367
R644 B.n550 B.n247 163.367
R645 B.n554 B.n247 163.367
R646 B.n554 B.n241 163.367
R647 B.n563 B.n241 163.367
R648 B.n563 B.n239 163.367
R649 B.n567 B.n239 163.367
R650 B.n567 B.n3 163.367
R651 B.n685 B.n3 163.367
R652 B.n681 B.n2 163.367
R653 B.n681 B.n680 163.367
R654 B.n680 B.n9 163.367
R655 B.n676 B.n9 163.367
R656 B.n676 B.n11 163.367
R657 B.n672 B.n11 163.367
R658 B.n672 B.n16 163.367
R659 B.n668 B.n16 163.367
R660 B.n668 B.n18 163.367
R661 B.n664 B.n18 163.367
R662 B.n664 B.n23 163.367
R663 B.n660 B.n23 163.367
R664 B.n660 B.n25 163.367
R665 B.n656 B.n25 163.367
R666 B.n656 B.n30 163.367
R667 B.n652 B.n30 163.367
R668 B.n652 B.n32 163.367
R669 B.n648 B.n32 163.367
R670 B.n648 B.n37 163.367
R671 B.n644 B.n37 163.367
R672 B.n644 B.n39 163.367
R673 B.n640 B.n39 163.367
R674 B.n640 B.n44 163.367
R675 B.n636 B.n44 163.367
R676 B.n636 B.n46 163.367
R677 B.n632 B.n46 163.367
R678 B.n632 B.n50 163.367
R679 B.n628 B.n50 163.367
R680 B.n628 B.n52 163.367
R681 B.n624 B.n52 163.367
R682 B.n624 B.n58 163.367
R683 B.n620 B.n58 163.367
R684 B.n476 B.n297 90.4569
R685 B.n619 B.n618 90.4569
R686 B.n62 B.n60 71.676
R687 B.n104 B.n63 71.676
R688 B.n108 B.n64 71.676
R689 B.n112 B.n65 71.676
R690 B.n116 B.n66 71.676
R691 B.n120 B.n67 71.676
R692 B.n124 B.n68 71.676
R693 B.n128 B.n69 71.676
R694 B.n132 B.n70 71.676
R695 B.n136 B.n71 71.676
R696 B.n140 B.n72 71.676
R697 B.n144 B.n73 71.676
R698 B.n148 B.n74 71.676
R699 B.n152 B.n75 71.676
R700 B.n156 B.n76 71.676
R701 B.n160 B.n77 71.676
R702 B.n164 B.n78 71.676
R703 B.n168 B.n79 71.676
R704 B.n172 B.n80 71.676
R705 B.n176 B.n81 71.676
R706 B.n181 B.n82 71.676
R707 B.n185 B.n83 71.676
R708 B.n189 B.n84 71.676
R709 B.n193 B.n85 71.676
R710 B.n197 B.n86 71.676
R711 B.n201 B.n87 71.676
R712 B.n205 B.n88 71.676
R713 B.n209 B.n89 71.676
R714 B.n213 B.n90 71.676
R715 B.n217 B.n91 71.676
R716 B.n221 B.n92 71.676
R717 B.n225 B.n93 71.676
R718 B.n229 B.n94 71.676
R719 B.n233 B.n95 71.676
R720 B.n96 B.n95 71.676
R721 B.n232 B.n94 71.676
R722 B.n228 B.n93 71.676
R723 B.n224 B.n92 71.676
R724 B.n220 B.n91 71.676
R725 B.n216 B.n90 71.676
R726 B.n212 B.n89 71.676
R727 B.n208 B.n88 71.676
R728 B.n204 B.n87 71.676
R729 B.n200 B.n86 71.676
R730 B.n196 B.n85 71.676
R731 B.n192 B.n84 71.676
R732 B.n188 B.n83 71.676
R733 B.n184 B.n82 71.676
R734 B.n180 B.n81 71.676
R735 B.n175 B.n80 71.676
R736 B.n171 B.n79 71.676
R737 B.n167 B.n78 71.676
R738 B.n163 B.n77 71.676
R739 B.n159 B.n76 71.676
R740 B.n155 B.n75 71.676
R741 B.n151 B.n74 71.676
R742 B.n147 B.n73 71.676
R743 B.n143 B.n72 71.676
R744 B.n139 B.n71 71.676
R745 B.n135 B.n70 71.676
R746 B.n131 B.n69 71.676
R747 B.n127 B.n68 71.676
R748 B.n123 B.n67 71.676
R749 B.n119 B.n66 71.676
R750 B.n115 B.n65 71.676
R751 B.n111 B.n64 71.676
R752 B.n107 B.n63 71.676
R753 B.n103 B.n62 71.676
R754 B.n336 B.n296 71.676
R755 B.n340 B.n339 71.676
R756 B.n345 B.n344 71.676
R757 B.n348 B.n347 71.676
R758 B.n353 B.n352 71.676
R759 B.n356 B.n355 71.676
R760 B.n361 B.n360 71.676
R761 B.n364 B.n363 71.676
R762 B.n369 B.n368 71.676
R763 B.n372 B.n371 71.676
R764 B.n377 B.n376 71.676
R765 B.n380 B.n379 71.676
R766 B.n385 B.n384 71.676
R767 B.n388 B.n387 71.676
R768 B.n396 B.n395 71.676
R769 B.n399 B.n398 71.676
R770 B.n404 B.n403 71.676
R771 B.n407 B.n406 71.676
R772 B.n412 B.n411 71.676
R773 B.n415 B.n414 71.676
R774 B.n420 B.n419 71.676
R775 B.n423 B.n422 71.676
R776 B.n428 B.n427 71.676
R777 B.n431 B.n430 71.676
R778 B.n436 B.n435 71.676
R779 B.n439 B.n438 71.676
R780 B.n444 B.n443 71.676
R781 B.n447 B.n446 71.676
R782 B.n452 B.n451 71.676
R783 B.n455 B.n454 71.676
R784 B.n460 B.n459 71.676
R785 B.n463 B.n462 71.676
R786 B.n468 B.n467 71.676
R787 B.n471 B.n470 71.676
R788 B.n337 B.n336 71.676
R789 B.n339 B.n333 71.676
R790 B.n346 B.n345 71.676
R791 B.n347 B.n331 71.676
R792 B.n354 B.n353 71.676
R793 B.n355 B.n329 71.676
R794 B.n362 B.n361 71.676
R795 B.n363 B.n327 71.676
R796 B.n370 B.n369 71.676
R797 B.n371 B.n325 71.676
R798 B.n378 B.n377 71.676
R799 B.n379 B.n323 71.676
R800 B.n386 B.n385 71.676
R801 B.n387 B.n321 71.676
R802 B.n397 B.n396 71.676
R803 B.n398 B.n319 71.676
R804 B.n405 B.n404 71.676
R805 B.n406 B.n317 71.676
R806 B.n413 B.n412 71.676
R807 B.n414 B.n312 71.676
R808 B.n421 B.n420 71.676
R809 B.n422 B.n310 71.676
R810 B.n429 B.n428 71.676
R811 B.n430 B.n308 71.676
R812 B.n437 B.n436 71.676
R813 B.n438 B.n306 71.676
R814 B.n445 B.n444 71.676
R815 B.n446 B.n304 71.676
R816 B.n453 B.n452 71.676
R817 B.n454 B.n302 71.676
R818 B.n461 B.n460 71.676
R819 B.n462 B.n300 71.676
R820 B.n469 B.n468 71.676
R821 B.n470 B.n298 71.676
R822 B.n686 B.n685 71.676
R823 B.n686 B.n2 71.676
R824 B.n101 B.n100 59.5399
R825 B.n178 B.n98 59.5399
R826 B.n315 B.n314 59.5399
R827 B.n393 B.n392 59.5399
R828 B.n476 B.n293 56.432
R829 B.n482 B.n293 56.432
R830 B.n482 B.n289 56.432
R831 B.n489 B.n289 56.432
R832 B.n489 B.n488 56.432
R833 B.n495 B.n282 56.432
R834 B.n501 B.n282 56.432
R835 B.n501 B.n278 56.432
R836 B.n507 B.n278 56.432
R837 B.n507 B.n274 56.432
R838 B.n513 B.n274 56.432
R839 B.n519 B.n270 56.432
R840 B.n519 B.n266 56.432
R841 B.n525 B.n266 56.432
R842 B.n531 B.n262 56.432
R843 B.n531 B.n258 56.432
R844 B.n537 B.n258 56.432
R845 B.n543 B.n254 56.432
R846 B.n543 B.n250 56.432
R847 B.n549 B.n250 56.432
R848 B.n555 B.n246 56.432
R849 B.n555 B.n242 56.432
R850 B.n562 B.n242 56.432
R851 B.n568 B.n238 56.432
R852 B.n568 B.n4 56.432
R853 B.n684 B.n4 56.432
R854 B.n684 B.n683 56.432
R855 B.n683 B.n682 56.432
R856 B.n682 B.n8 56.432
R857 B.n577 B.n8 56.432
R858 B.n675 B.n674 56.432
R859 B.n674 B.n673 56.432
R860 B.n673 B.n15 56.432
R861 B.n667 B.n666 56.432
R862 B.n666 B.n665 56.432
R863 B.n665 B.n22 56.432
R864 B.n659 B.n658 56.432
R865 B.n658 B.n657 56.432
R866 B.n657 B.n29 56.432
R867 B.n651 B.n650 56.432
R868 B.n650 B.n649 56.432
R869 B.n649 B.n36 56.432
R870 B.n643 B.n642 56.432
R871 B.n642 B.n641 56.432
R872 B.n641 B.n43 56.432
R873 B.n635 B.n43 56.432
R874 B.n635 B.n634 56.432
R875 B.n634 B.n633 56.432
R876 B.n627 B.n53 56.432
R877 B.n627 B.n626 56.432
R878 B.n626 B.n625 56.432
R879 B.n625 B.n57 56.432
R880 B.n619 B.n57 56.432
R881 B.n562 B.t3 49.793
R882 B.n675 B.t5 49.793
R883 B.n549 B.t0 48.1333
R884 B.n667 B.t8 48.1333
R885 B.n537 B.t6 46.4735
R886 B.n659 B.t1 46.4735
R887 B.n525 B.t2 44.8138
R888 B.n651 B.t4 44.8138
R889 B.n513 B.t7 43.154
R890 B.n643 B.t9 43.154
R891 B.n478 B.n295 31.0639
R892 B.n474 B.n473 31.0639
R893 B.n616 B.n615 31.0639
R894 B.n621 B.n59 31.0639
R895 B.n488 B.t11 29.876
R896 B.n53 B.t15 29.876
R897 B.n100 B.n99 26.5702
R898 B.n98 B.n97 26.5702
R899 B.n314 B.n313 26.5702
R900 B.n392 B.n391 26.5702
R901 B.n495 B.t11 26.5565
R902 B.n633 B.t15 26.5565
R903 B B.n687 18.0485
R904 B.t7 B.n270 13.2785
R905 B.t9 B.n36 13.2785
R906 B.t2 B.n262 11.6188
R907 B.t4 B.n29 11.6188
R908 B.n479 B.n478 10.6151
R909 B.n480 B.n479 10.6151
R910 B.n480 B.n287 10.6151
R911 B.n491 B.n287 10.6151
R912 B.n492 B.n491 10.6151
R913 B.n493 B.n492 10.6151
R914 B.n493 B.n280 10.6151
R915 B.n503 B.n280 10.6151
R916 B.n504 B.n503 10.6151
R917 B.n505 B.n504 10.6151
R918 B.n505 B.n272 10.6151
R919 B.n515 B.n272 10.6151
R920 B.n516 B.n515 10.6151
R921 B.n517 B.n516 10.6151
R922 B.n517 B.n264 10.6151
R923 B.n527 B.n264 10.6151
R924 B.n528 B.n527 10.6151
R925 B.n529 B.n528 10.6151
R926 B.n529 B.n256 10.6151
R927 B.n539 B.n256 10.6151
R928 B.n540 B.n539 10.6151
R929 B.n541 B.n540 10.6151
R930 B.n541 B.n248 10.6151
R931 B.n551 B.n248 10.6151
R932 B.n552 B.n551 10.6151
R933 B.n553 B.n552 10.6151
R934 B.n553 B.n240 10.6151
R935 B.n564 B.n240 10.6151
R936 B.n565 B.n564 10.6151
R937 B.n566 B.n565 10.6151
R938 B.n566 B.n0 10.6151
R939 B.n335 B.n295 10.6151
R940 B.n335 B.n334 10.6151
R941 B.n341 B.n334 10.6151
R942 B.n342 B.n341 10.6151
R943 B.n343 B.n342 10.6151
R944 B.n343 B.n332 10.6151
R945 B.n349 B.n332 10.6151
R946 B.n350 B.n349 10.6151
R947 B.n351 B.n350 10.6151
R948 B.n351 B.n330 10.6151
R949 B.n357 B.n330 10.6151
R950 B.n358 B.n357 10.6151
R951 B.n359 B.n358 10.6151
R952 B.n359 B.n328 10.6151
R953 B.n365 B.n328 10.6151
R954 B.n366 B.n365 10.6151
R955 B.n367 B.n366 10.6151
R956 B.n367 B.n326 10.6151
R957 B.n373 B.n326 10.6151
R958 B.n374 B.n373 10.6151
R959 B.n375 B.n374 10.6151
R960 B.n375 B.n324 10.6151
R961 B.n381 B.n324 10.6151
R962 B.n382 B.n381 10.6151
R963 B.n383 B.n382 10.6151
R964 B.n383 B.n322 10.6151
R965 B.n389 B.n322 10.6151
R966 B.n390 B.n389 10.6151
R967 B.n394 B.n390 10.6151
R968 B.n400 B.n320 10.6151
R969 B.n401 B.n400 10.6151
R970 B.n402 B.n401 10.6151
R971 B.n402 B.n318 10.6151
R972 B.n408 B.n318 10.6151
R973 B.n409 B.n408 10.6151
R974 B.n410 B.n409 10.6151
R975 B.n410 B.n316 10.6151
R976 B.n417 B.n416 10.6151
R977 B.n418 B.n417 10.6151
R978 B.n418 B.n311 10.6151
R979 B.n424 B.n311 10.6151
R980 B.n425 B.n424 10.6151
R981 B.n426 B.n425 10.6151
R982 B.n426 B.n309 10.6151
R983 B.n432 B.n309 10.6151
R984 B.n433 B.n432 10.6151
R985 B.n434 B.n433 10.6151
R986 B.n434 B.n307 10.6151
R987 B.n440 B.n307 10.6151
R988 B.n441 B.n440 10.6151
R989 B.n442 B.n441 10.6151
R990 B.n442 B.n305 10.6151
R991 B.n448 B.n305 10.6151
R992 B.n449 B.n448 10.6151
R993 B.n450 B.n449 10.6151
R994 B.n450 B.n303 10.6151
R995 B.n456 B.n303 10.6151
R996 B.n457 B.n456 10.6151
R997 B.n458 B.n457 10.6151
R998 B.n458 B.n301 10.6151
R999 B.n464 B.n301 10.6151
R1000 B.n465 B.n464 10.6151
R1001 B.n466 B.n465 10.6151
R1002 B.n466 B.n299 10.6151
R1003 B.n472 B.n299 10.6151
R1004 B.n473 B.n472 10.6151
R1005 B.n474 B.n291 10.6151
R1006 B.n484 B.n291 10.6151
R1007 B.n485 B.n484 10.6151
R1008 B.n486 B.n485 10.6151
R1009 B.n486 B.n284 10.6151
R1010 B.n497 B.n284 10.6151
R1011 B.n498 B.n497 10.6151
R1012 B.n499 B.n498 10.6151
R1013 B.n499 B.n276 10.6151
R1014 B.n509 B.n276 10.6151
R1015 B.n510 B.n509 10.6151
R1016 B.n511 B.n510 10.6151
R1017 B.n511 B.n268 10.6151
R1018 B.n521 B.n268 10.6151
R1019 B.n522 B.n521 10.6151
R1020 B.n523 B.n522 10.6151
R1021 B.n523 B.n260 10.6151
R1022 B.n533 B.n260 10.6151
R1023 B.n534 B.n533 10.6151
R1024 B.n535 B.n534 10.6151
R1025 B.n535 B.n252 10.6151
R1026 B.n545 B.n252 10.6151
R1027 B.n546 B.n545 10.6151
R1028 B.n547 B.n546 10.6151
R1029 B.n547 B.n244 10.6151
R1030 B.n557 B.n244 10.6151
R1031 B.n558 B.n557 10.6151
R1032 B.n560 B.n558 10.6151
R1033 B.n560 B.n559 10.6151
R1034 B.n559 B.n236 10.6151
R1035 B.n571 B.n236 10.6151
R1036 B.n572 B.n571 10.6151
R1037 B.n573 B.n572 10.6151
R1038 B.n574 B.n573 10.6151
R1039 B.n575 B.n574 10.6151
R1040 B.n579 B.n575 10.6151
R1041 B.n580 B.n579 10.6151
R1042 B.n581 B.n580 10.6151
R1043 B.n582 B.n581 10.6151
R1044 B.n584 B.n582 10.6151
R1045 B.n585 B.n584 10.6151
R1046 B.n586 B.n585 10.6151
R1047 B.n587 B.n586 10.6151
R1048 B.n589 B.n587 10.6151
R1049 B.n590 B.n589 10.6151
R1050 B.n591 B.n590 10.6151
R1051 B.n592 B.n591 10.6151
R1052 B.n594 B.n592 10.6151
R1053 B.n595 B.n594 10.6151
R1054 B.n596 B.n595 10.6151
R1055 B.n597 B.n596 10.6151
R1056 B.n599 B.n597 10.6151
R1057 B.n600 B.n599 10.6151
R1058 B.n601 B.n600 10.6151
R1059 B.n602 B.n601 10.6151
R1060 B.n604 B.n602 10.6151
R1061 B.n605 B.n604 10.6151
R1062 B.n606 B.n605 10.6151
R1063 B.n607 B.n606 10.6151
R1064 B.n609 B.n607 10.6151
R1065 B.n610 B.n609 10.6151
R1066 B.n611 B.n610 10.6151
R1067 B.n612 B.n611 10.6151
R1068 B.n614 B.n612 10.6151
R1069 B.n615 B.n614 10.6151
R1070 B.n679 B.n1 10.6151
R1071 B.n679 B.n678 10.6151
R1072 B.n678 B.n677 10.6151
R1073 B.n677 B.n10 10.6151
R1074 B.n671 B.n10 10.6151
R1075 B.n671 B.n670 10.6151
R1076 B.n670 B.n669 10.6151
R1077 B.n669 B.n17 10.6151
R1078 B.n663 B.n17 10.6151
R1079 B.n663 B.n662 10.6151
R1080 B.n662 B.n661 10.6151
R1081 B.n661 B.n24 10.6151
R1082 B.n655 B.n24 10.6151
R1083 B.n655 B.n654 10.6151
R1084 B.n654 B.n653 10.6151
R1085 B.n653 B.n31 10.6151
R1086 B.n647 B.n31 10.6151
R1087 B.n647 B.n646 10.6151
R1088 B.n646 B.n645 10.6151
R1089 B.n645 B.n38 10.6151
R1090 B.n639 B.n38 10.6151
R1091 B.n639 B.n638 10.6151
R1092 B.n638 B.n637 10.6151
R1093 B.n637 B.n45 10.6151
R1094 B.n631 B.n45 10.6151
R1095 B.n631 B.n630 10.6151
R1096 B.n630 B.n629 10.6151
R1097 B.n629 B.n51 10.6151
R1098 B.n623 B.n51 10.6151
R1099 B.n623 B.n622 10.6151
R1100 B.n622 B.n621 10.6151
R1101 B.n102 B.n59 10.6151
R1102 B.n105 B.n102 10.6151
R1103 B.n106 B.n105 10.6151
R1104 B.n109 B.n106 10.6151
R1105 B.n110 B.n109 10.6151
R1106 B.n113 B.n110 10.6151
R1107 B.n114 B.n113 10.6151
R1108 B.n117 B.n114 10.6151
R1109 B.n118 B.n117 10.6151
R1110 B.n121 B.n118 10.6151
R1111 B.n122 B.n121 10.6151
R1112 B.n125 B.n122 10.6151
R1113 B.n126 B.n125 10.6151
R1114 B.n129 B.n126 10.6151
R1115 B.n130 B.n129 10.6151
R1116 B.n133 B.n130 10.6151
R1117 B.n134 B.n133 10.6151
R1118 B.n137 B.n134 10.6151
R1119 B.n138 B.n137 10.6151
R1120 B.n141 B.n138 10.6151
R1121 B.n142 B.n141 10.6151
R1122 B.n145 B.n142 10.6151
R1123 B.n146 B.n145 10.6151
R1124 B.n149 B.n146 10.6151
R1125 B.n150 B.n149 10.6151
R1126 B.n153 B.n150 10.6151
R1127 B.n154 B.n153 10.6151
R1128 B.n157 B.n154 10.6151
R1129 B.n158 B.n157 10.6151
R1130 B.n162 B.n161 10.6151
R1131 B.n165 B.n162 10.6151
R1132 B.n166 B.n165 10.6151
R1133 B.n169 B.n166 10.6151
R1134 B.n170 B.n169 10.6151
R1135 B.n173 B.n170 10.6151
R1136 B.n174 B.n173 10.6151
R1137 B.n177 B.n174 10.6151
R1138 B.n182 B.n179 10.6151
R1139 B.n183 B.n182 10.6151
R1140 B.n186 B.n183 10.6151
R1141 B.n187 B.n186 10.6151
R1142 B.n190 B.n187 10.6151
R1143 B.n191 B.n190 10.6151
R1144 B.n194 B.n191 10.6151
R1145 B.n195 B.n194 10.6151
R1146 B.n198 B.n195 10.6151
R1147 B.n199 B.n198 10.6151
R1148 B.n202 B.n199 10.6151
R1149 B.n203 B.n202 10.6151
R1150 B.n206 B.n203 10.6151
R1151 B.n207 B.n206 10.6151
R1152 B.n210 B.n207 10.6151
R1153 B.n211 B.n210 10.6151
R1154 B.n214 B.n211 10.6151
R1155 B.n215 B.n214 10.6151
R1156 B.n218 B.n215 10.6151
R1157 B.n219 B.n218 10.6151
R1158 B.n222 B.n219 10.6151
R1159 B.n223 B.n222 10.6151
R1160 B.n226 B.n223 10.6151
R1161 B.n227 B.n226 10.6151
R1162 B.n230 B.n227 10.6151
R1163 B.n231 B.n230 10.6151
R1164 B.n234 B.n231 10.6151
R1165 B.n235 B.n234 10.6151
R1166 B.n616 B.n235 10.6151
R1167 B.t6 B.n254 9.95901
R1168 B.t1 B.n22 9.95901
R1169 B.t0 B.n246 8.29925
R1170 B.t8 B.n15 8.29925
R1171 B.n687 B.n0 8.11757
R1172 B.n687 B.n1 8.11757
R1173 B.t3 B.n238 6.6395
R1174 B.n577 B.t5 6.6395
R1175 B.n393 B.n320 6.5566
R1176 B.n316 B.n315 6.5566
R1177 B.n161 B.n101 6.5566
R1178 B.n178 B.n177 6.5566
R1179 B.n394 B.n393 4.05904
R1180 B.n416 B.n315 4.05904
R1181 B.n158 B.n101 4.05904
R1182 B.n179 B.n178 4.05904
R1183 VN.n5 VN.t7 238.131
R1184 VN.n25 VN.t5 238.131
R1185 VN.n18 VN.t9 223.157
R1186 VN.n38 VN.t8 223.157
R1187 VN.n4 VN.t6 184.922
R1188 VN.n10 VN.t4 184.922
R1189 VN.n16 VN.t3 184.922
R1190 VN.n24 VN.t1 184.922
R1191 VN.n30 VN.t2 184.922
R1192 VN.n36 VN.t0 184.922
R1193 VN.n37 VN.n20 161.3
R1194 VN.n35 VN.n34 161.3
R1195 VN.n33 VN.n21 161.3
R1196 VN.n32 VN.n31 161.3
R1197 VN.n29 VN.n22 161.3
R1198 VN.n28 VN.n27 161.3
R1199 VN.n26 VN.n23 161.3
R1200 VN.n17 VN.n0 161.3
R1201 VN.n15 VN.n14 161.3
R1202 VN.n13 VN.n1 161.3
R1203 VN.n12 VN.n11 161.3
R1204 VN.n9 VN.n2 161.3
R1205 VN.n8 VN.n7 161.3
R1206 VN.n6 VN.n3 161.3
R1207 VN.n39 VN.n38 80.6037
R1208 VN.n19 VN.n18 80.6037
R1209 VN.n18 VN.n17 55.0167
R1210 VN.n38 VN.n37 55.0167
R1211 VN.n5 VN.n4 48.3607
R1212 VN.n25 VN.n24 48.3607
R1213 VN.n9 VN.n8 46.7399
R1214 VN.n11 VN.n1 46.7399
R1215 VN.n29 VN.n28 46.7399
R1216 VN.n31 VN.n21 46.7399
R1217 VN.n26 VN.n25 44.0902
R1218 VN.n6 VN.n5 44.0902
R1219 VN VN.n39 42.0938
R1220 VN.n8 VN.n3 34.0813
R1221 VN.n15 VN.n1 34.0813
R1222 VN.n28 VN.n23 34.0813
R1223 VN.n35 VN.n21 34.0813
R1224 VN.n17 VN.n16 18.5015
R1225 VN.n37 VN.n36 18.5015
R1226 VN.n10 VN.n9 12.1722
R1227 VN.n11 VN.n10 12.1722
R1228 VN.n31 VN.n30 12.1722
R1229 VN.n30 VN.n29 12.1722
R1230 VN.n4 VN.n3 5.84292
R1231 VN.n16 VN.n15 5.84292
R1232 VN.n24 VN.n23 5.84292
R1233 VN.n36 VN.n35 5.84292
R1234 VN.n39 VN.n20 0.285035
R1235 VN.n19 VN.n0 0.285035
R1236 VN.n34 VN.n20 0.189894
R1237 VN.n34 VN.n33 0.189894
R1238 VN.n33 VN.n32 0.189894
R1239 VN.n32 VN.n22 0.189894
R1240 VN.n27 VN.n22 0.189894
R1241 VN.n27 VN.n26 0.189894
R1242 VN.n7 VN.n6 0.189894
R1243 VN.n7 VN.n2 0.189894
R1244 VN.n12 VN.n2 0.189894
R1245 VN.n13 VN.n12 0.189894
R1246 VN.n14 VN.n13 0.189894
R1247 VN.n14 VN.n0 0.189894
R1248 VN VN.n19 0.146778
R1249 VDD2.n81 VDD2.n45 289.615
R1250 VDD2.n36 VDD2.n0 289.615
R1251 VDD2.n82 VDD2.n81 185
R1252 VDD2.n80 VDD2.n47 185
R1253 VDD2.n79 VDD2.n78 185
R1254 VDD2.n50 VDD2.n48 185
R1255 VDD2.n73 VDD2.n72 185
R1256 VDD2.n71 VDD2.n70 185
R1257 VDD2.n54 VDD2.n53 185
R1258 VDD2.n65 VDD2.n64 185
R1259 VDD2.n63 VDD2.n62 185
R1260 VDD2.n58 VDD2.n57 185
R1261 VDD2.n12 VDD2.n11 185
R1262 VDD2.n17 VDD2.n16 185
R1263 VDD2.n19 VDD2.n18 185
R1264 VDD2.n8 VDD2.n7 185
R1265 VDD2.n25 VDD2.n24 185
R1266 VDD2.n27 VDD2.n26 185
R1267 VDD2.n4 VDD2.n3 185
R1268 VDD2.n34 VDD2.n33 185
R1269 VDD2.n35 VDD2.n2 185
R1270 VDD2.n37 VDD2.n36 185
R1271 VDD2.n59 VDD2.t2 149.524
R1272 VDD2.n13 VDD2.t3 149.524
R1273 VDD2.n81 VDD2.n80 104.615
R1274 VDD2.n80 VDD2.n79 104.615
R1275 VDD2.n79 VDD2.n48 104.615
R1276 VDD2.n72 VDD2.n48 104.615
R1277 VDD2.n72 VDD2.n71 104.615
R1278 VDD2.n71 VDD2.n53 104.615
R1279 VDD2.n64 VDD2.n53 104.615
R1280 VDD2.n64 VDD2.n63 104.615
R1281 VDD2.n63 VDD2.n57 104.615
R1282 VDD2.n17 VDD2.n11 104.615
R1283 VDD2.n18 VDD2.n17 104.615
R1284 VDD2.n18 VDD2.n7 104.615
R1285 VDD2.n25 VDD2.n7 104.615
R1286 VDD2.n26 VDD2.n25 104.615
R1287 VDD2.n26 VDD2.n3 104.615
R1288 VDD2.n34 VDD2.n3 104.615
R1289 VDD2.n35 VDD2.n34 104.615
R1290 VDD2.n36 VDD2.n35 104.615
R1291 VDD2.n44 VDD2.n43 68.2991
R1292 VDD2 VDD2.n89 68.2963
R1293 VDD2.n88 VDD2.n87 67.4689
R1294 VDD2.n42 VDD2.n41 67.4687
R1295 VDD2.n42 VDD2.n40 53.5361
R1296 VDD2.n86 VDD2.n85 52.355
R1297 VDD2.t2 VDD2.n57 52.3082
R1298 VDD2.t3 VDD2.n11 52.3082
R1299 VDD2.n86 VDD2.n44 36.2045
R1300 VDD2.n82 VDD2.n47 13.1884
R1301 VDD2.n37 VDD2.n2 13.1884
R1302 VDD2.n83 VDD2.n45 12.8005
R1303 VDD2.n78 VDD2.n49 12.8005
R1304 VDD2.n33 VDD2.n32 12.8005
R1305 VDD2.n38 VDD2.n0 12.8005
R1306 VDD2.n77 VDD2.n50 12.0247
R1307 VDD2.n31 VDD2.n4 12.0247
R1308 VDD2.n74 VDD2.n73 11.249
R1309 VDD2.n28 VDD2.n27 11.249
R1310 VDD2.n70 VDD2.n52 10.4732
R1311 VDD2.n24 VDD2.n6 10.4732
R1312 VDD2.n59 VDD2.n58 10.2747
R1313 VDD2.n13 VDD2.n12 10.2747
R1314 VDD2.n69 VDD2.n54 9.69747
R1315 VDD2.n23 VDD2.n8 9.69747
R1316 VDD2.n85 VDD2.n84 9.45567
R1317 VDD2.n40 VDD2.n39 9.45567
R1318 VDD2.n61 VDD2.n60 9.3005
R1319 VDD2.n56 VDD2.n55 9.3005
R1320 VDD2.n67 VDD2.n66 9.3005
R1321 VDD2.n69 VDD2.n68 9.3005
R1322 VDD2.n52 VDD2.n51 9.3005
R1323 VDD2.n75 VDD2.n74 9.3005
R1324 VDD2.n77 VDD2.n76 9.3005
R1325 VDD2.n49 VDD2.n46 9.3005
R1326 VDD2.n84 VDD2.n83 9.3005
R1327 VDD2.n39 VDD2.n38 9.3005
R1328 VDD2.n15 VDD2.n14 9.3005
R1329 VDD2.n10 VDD2.n9 9.3005
R1330 VDD2.n21 VDD2.n20 9.3005
R1331 VDD2.n23 VDD2.n22 9.3005
R1332 VDD2.n6 VDD2.n5 9.3005
R1333 VDD2.n29 VDD2.n28 9.3005
R1334 VDD2.n31 VDD2.n30 9.3005
R1335 VDD2.n32 VDD2.n1 9.3005
R1336 VDD2.n66 VDD2.n65 8.92171
R1337 VDD2.n20 VDD2.n19 8.92171
R1338 VDD2.n62 VDD2.n56 8.14595
R1339 VDD2.n16 VDD2.n10 8.14595
R1340 VDD2.n61 VDD2.n58 7.3702
R1341 VDD2.n15 VDD2.n12 7.3702
R1342 VDD2.n62 VDD2.n61 5.81868
R1343 VDD2.n16 VDD2.n15 5.81868
R1344 VDD2.n65 VDD2.n56 5.04292
R1345 VDD2.n19 VDD2.n10 5.04292
R1346 VDD2.n66 VDD2.n54 4.26717
R1347 VDD2.n20 VDD2.n8 4.26717
R1348 VDD2.n70 VDD2.n69 3.49141
R1349 VDD2.n24 VDD2.n23 3.49141
R1350 VDD2.n60 VDD2.n59 2.84304
R1351 VDD2.n14 VDD2.n13 2.84304
R1352 VDD2.n73 VDD2.n52 2.71565
R1353 VDD2.n27 VDD2.n6 2.71565
R1354 VDD2.n89 VDD2.t7 2.4817
R1355 VDD2.n89 VDD2.t1 2.4817
R1356 VDD2.n87 VDD2.t6 2.4817
R1357 VDD2.n87 VDD2.t4 2.4817
R1358 VDD2.n43 VDD2.t5 2.4817
R1359 VDD2.n43 VDD2.t0 2.4817
R1360 VDD2.n41 VDD2.t9 2.4817
R1361 VDD2.n41 VDD2.t8 2.4817
R1362 VDD2.n74 VDD2.n50 1.93989
R1363 VDD2.n28 VDD2.n4 1.93989
R1364 VDD2.n88 VDD2.n86 1.18153
R1365 VDD2.n85 VDD2.n45 1.16414
R1366 VDD2.n78 VDD2.n77 1.16414
R1367 VDD2.n33 VDD2.n31 1.16414
R1368 VDD2.n40 VDD2.n0 1.16414
R1369 VDD2.n83 VDD2.n82 0.388379
R1370 VDD2.n49 VDD2.n47 0.388379
R1371 VDD2.n32 VDD2.n2 0.388379
R1372 VDD2.n38 VDD2.n37 0.388379
R1373 VDD2 VDD2.n88 0.353948
R1374 VDD2.n44 VDD2.n42 0.240413
R1375 VDD2.n84 VDD2.n46 0.155672
R1376 VDD2.n76 VDD2.n46 0.155672
R1377 VDD2.n76 VDD2.n75 0.155672
R1378 VDD2.n75 VDD2.n51 0.155672
R1379 VDD2.n68 VDD2.n51 0.155672
R1380 VDD2.n68 VDD2.n67 0.155672
R1381 VDD2.n67 VDD2.n55 0.155672
R1382 VDD2.n60 VDD2.n55 0.155672
R1383 VDD2.n14 VDD2.n9 0.155672
R1384 VDD2.n21 VDD2.n9 0.155672
R1385 VDD2.n22 VDD2.n21 0.155672
R1386 VDD2.n22 VDD2.n5 0.155672
R1387 VDD2.n29 VDD2.n5 0.155672
R1388 VDD2.n30 VDD2.n29 0.155672
R1389 VDD2.n30 VDD2.n1 0.155672
R1390 VDD2.n39 VDD2.n1 0.155672
R1391 VTAIL.n176 VTAIL.n140 289.615
R1392 VTAIL.n38 VTAIL.n2 289.615
R1393 VTAIL.n134 VTAIL.n98 289.615
R1394 VTAIL.n88 VTAIL.n52 289.615
R1395 VTAIL.n152 VTAIL.n151 185
R1396 VTAIL.n157 VTAIL.n156 185
R1397 VTAIL.n159 VTAIL.n158 185
R1398 VTAIL.n148 VTAIL.n147 185
R1399 VTAIL.n165 VTAIL.n164 185
R1400 VTAIL.n167 VTAIL.n166 185
R1401 VTAIL.n144 VTAIL.n143 185
R1402 VTAIL.n174 VTAIL.n173 185
R1403 VTAIL.n175 VTAIL.n142 185
R1404 VTAIL.n177 VTAIL.n176 185
R1405 VTAIL.n14 VTAIL.n13 185
R1406 VTAIL.n19 VTAIL.n18 185
R1407 VTAIL.n21 VTAIL.n20 185
R1408 VTAIL.n10 VTAIL.n9 185
R1409 VTAIL.n27 VTAIL.n26 185
R1410 VTAIL.n29 VTAIL.n28 185
R1411 VTAIL.n6 VTAIL.n5 185
R1412 VTAIL.n36 VTAIL.n35 185
R1413 VTAIL.n37 VTAIL.n4 185
R1414 VTAIL.n39 VTAIL.n38 185
R1415 VTAIL.n135 VTAIL.n134 185
R1416 VTAIL.n133 VTAIL.n100 185
R1417 VTAIL.n132 VTAIL.n131 185
R1418 VTAIL.n103 VTAIL.n101 185
R1419 VTAIL.n126 VTAIL.n125 185
R1420 VTAIL.n124 VTAIL.n123 185
R1421 VTAIL.n107 VTAIL.n106 185
R1422 VTAIL.n118 VTAIL.n117 185
R1423 VTAIL.n116 VTAIL.n115 185
R1424 VTAIL.n111 VTAIL.n110 185
R1425 VTAIL.n89 VTAIL.n88 185
R1426 VTAIL.n87 VTAIL.n54 185
R1427 VTAIL.n86 VTAIL.n85 185
R1428 VTAIL.n57 VTAIL.n55 185
R1429 VTAIL.n80 VTAIL.n79 185
R1430 VTAIL.n78 VTAIL.n77 185
R1431 VTAIL.n61 VTAIL.n60 185
R1432 VTAIL.n72 VTAIL.n71 185
R1433 VTAIL.n70 VTAIL.n69 185
R1434 VTAIL.n65 VTAIL.n64 185
R1435 VTAIL.n153 VTAIL.t9 149.524
R1436 VTAIL.n15 VTAIL.t1 149.524
R1437 VTAIL.n112 VTAIL.t7 149.524
R1438 VTAIL.n66 VTAIL.t13 149.524
R1439 VTAIL.n157 VTAIL.n151 104.615
R1440 VTAIL.n158 VTAIL.n157 104.615
R1441 VTAIL.n158 VTAIL.n147 104.615
R1442 VTAIL.n165 VTAIL.n147 104.615
R1443 VTAIL.n166 VTAIL.n165 104.615
R1444 VTAIL.n166 VTAIL.n143 104.615
R1445 VTAIL.n174 VTAIL.n143 104.615
R1446 VTAIL.n175 VTAIL.n174 104.615
R1447 VTAIL.n176 VTAIL.n175 104.615
R1448 VTAIL.n19 VTAIL.n13 104.615
R1449 VTAIL.n20 VTAIL.n19 104.615
R1450 VTAIL.n20 VTAIL.n9 104.615
R1451 VTAIL.n27 VTAIL.n9 104.615
R1452 VTAIL.n28 VTAIL.n27 104.615
R1453 VTAIL.n28 VTAIL.n5 104.615
R1454 VTAIL.n36 VTAIL.n5 104.615
R1455 VTAIL.n37 VTAIL.n36 104.615
R1456 VTAIL.n38 VTAIL.n37 104.615
R1457 VTAIL.n134 VTAIL.n133 104.615
R1458 VTAIL.n133 VTAIL.n132 104.615
R1459 VTAIL.n132 VTAIL.n101 104.615
R1460 VTAIL.n125 VTAIL.n101 104.615
R1461 VTAIL.n125 VTAIL.n124 104.615
R1462 VTAIL.n124 VTAIL.n106 104.615
R1463 VTAIL.n117 VTAIL.n106 104.615
R1464 VTAIL.n117 VTAIL.n116 104.615
R1465 VTAIL.n116 VTAIL.n110 104.615
R1466 VTAIL.n88 VTAIL.n87 104.615
R1467 VTAIL.n87 VTAIL.n86 104.615
R1468 VTAIL.n86 VTAIL.n55 104.615
R1469 VTAIL.n79 VTAIL.n55 104.615
R1470 VTAIL.n79 VTAIL.n78 104.615
R1471 VTAIL.n78 VTAIL.n60 104.615
R1472 VTAIL.n71 VTAIL.n60 104.615
R1473 VTAIL.n71 VTAIL.n70 104.615
R1474 VTAIL.n70 VTAIL.n64 104.615
R1475 VTAIL.t9 VTAIL.n151 52.3082
R1476 VTAIL.t1 VTAIL.n13 52.3082
R1477 VTAIL.t7 VTAIL.n110 52.3082
R1478 VTAIL.t13 VTAIL.n64 52.3082
R1479 VTAIL.n97 VTAIL.n96 50.7901
R1480 VTAIL.n95 VTAIL.n94 50.7901
R1481 VTAIL.n51 VTAIL.n50 50.7901
R1482 VTAIL.n49 VTAIL.n48 50.7901
R1483 VTAIL.n183 VTAIL.n182 50.7899
R1484 VTAIL.n1 VTAIL.n0 50.7899
R1485 VTAIL.n45 VTAIL.n44 50.7899
R1486 VTAIL.n47 VTAIL.n46 50.7899
R1487 VTAIL.n181 VTAIL.n180 35.6763
R1488 VTAIL.n43 VTAIL.n42 35.6763
R1489 VTAIL.n139 VTAIL.n138 35.6763
R1490 VTAIL.n93 VTAIL.n92 35.6763
R1491 VTAIL.n49 VTAIL.n47 21.6083
R1492 VTAIL.n181 VTAIL.n139 20.4272
R1493 VTAIL.n177 VTAIL.n142 13.1884
R1494 VTAIL.n39 VTAIL.n4 13.1884
R1495 VTAIL.n135 VTAIL.n100 13.1884
R1496 VTAIL.n89 VTAIL.n54 13.1884
R1497 VTAIL.n173 VTAIL.n172 12.8005
R1498 VTAIL.n178 VTAIL.n140 12.8005
R1499 VTAIL.n35 VTAIL.n34 12.8005
R1500 VTAIL.n40 VTAIL.n2 12.8005
R1501 VTAIL.n136 VTAIL.n98 12.8005
R1502 VTAIL.n131 VTAIL.n102 12.8005
R1503 VTAIL.n90 VTAIL.n52 12.8005
R1504 VTAIL.n85 VTAIL.n56 12.8005
R1505 VTAIL.n171 VTAIL.n144 12.0247
R1506 VTAIL.n33 VTAIL.n6 12.0247
R1507 VTAIL.n130 VTAIL.n103 12.0247
R1508 VTAIL.n84 VTAIL.n57 12.0247
R1509 VTAIL.n168 VTAIL.n167 11.249
R1510 VTAIL.n30 VTAIL.n29 11.249
R1511 VTAIL.n127 VTAIL.n126 11.249
R1512 VTAIL.n81 VTAIL.n80 11.249
R1513 VTAIL.n164 VTAIL.n146 10.4732
R1514 VTAIL.n26 VTAIL.n8 10.4732
R1515 VTAIL.n123 VTAIL.n105 10.4732
R1516 VTAIL.n77 VTAIL.n59 10.4732
R1517 VTAIL.n153 VTAIL.n152 10.2747
R1518 VTAIL.n15 VTAIL.n14 10.2747
R1519 VTAIL.n112 VTAIL.n111 10.2747
R1520 VTAIL.n66 VTAIL.n65 10.2747
R1521 VTAIL.n163 VTAIL.n148 9.69747
R1522 VTAIL.n25 VTAIL.n10 9.69747
R1523 VTAIL.n122 VTAIL.n107 9.69747
R1524 VTAIL.n76 VTAIL.n61 9.69747
R1525 VTAIL.n180 VTAIL.n179 9.45567
R1526 VTAIL.n42 VTAIL.n41 9.45567
R1527 VTAIL.n138 VTAIL.n137 9.45567
R1528 VTAIL.n92 VTAIL.n91 9.45567
R1529 VTAIL.n179 VTAIL.n178 9.3005
R1530 VTAIL.n155 VTAIL.n154 9.3005
R1531 VTAIL.n150 VTAIL.n149 9.3005
R1532 VTAIL.n161 VTAIL.n160 9.3005
R1533 VTAIL.n163 VTAIL.n162 9.3005
R1534 VTAIL.n146 VTAIL.n145 9.3005
R1535 VTAIL.n169 VTAIL.n168 9.3005
R1536 VTAIL.n171 VTAIL.n170 9.3005
R1537 VTAIL.n172 VTAIL.n141 9.3005
R1538 VTAIL.n41 VTAIL.n40 9.3005
R1539 VTAIL.n17 VTAIL.n16 9.3005
R1540 VTAIL.n12 VTAIL.n11 9.3005
R1541 VTAIL.n23 VTAIL.n22 9.3005
R1542 VTAIL.n25 VTAIL.n24 9.3005
R1543 VTAIL.n8 VTAIL.n7 9.3005
R1544 VTAIL.n31 VTAIL.n30 9.3005
R1545 VTAIL.n33 VTAIL.n32 9.3005
R1546 VTAIL.n34 VTAIL.n3 9.3005
R1547 VTAIL.n114 VTAIL.n113 9.3005
R1548 VTAIL.n109 VTAIL.n108 9.3005
R1549 VTAIL.n120 VTAIL.n119 9.3005
R1550 VTAIL.n122 VTAIL.n121 9.3005
R1551 VTAIL.n105 VTAIL.n104 9.3005
R1552 VTAIL.n128 VTAIL.n127 9.3005
R1553 VTAIL.n130 VTAIL.n129 9.3005
R1554 VTAIL.n102 VTAIL.n99 9.3005
R1555 VTAIL.n137 VTAIL.n136 9.3005
R1556 VTAIL.n68 VTAIL.n67 9.3005
R1557 VTAIL.n63 VTAIL.n62 9.3005
R1558 VTAIL.n74 VTAIL.n73 9.3005
R1559 VTAIL.n76 VTAIL.n75 9.3005
R1560 VTAIL.n59 VTAIL.n58 9.3005
R1561 VTAIL.n82 VTAIL.n81 9.3005
R1562 VTAIL.n84 VTAIL.n83 9.3005
R1563 VTAIL.n56 VTAIL.n53 9.3005
R1564 VTAIL.n91 VTAIL.n90 9.3005
R1565 VTAIL.n160 VTAIL.n159 8.92171
R1566 VTAIL.n22 VTAIL.n21 8.92171
R1567 VTAIL.n119 VTAIL.n118 8.92171
R1568 VTAIL.n73 VTAIL.n72 8.92171
R1569 VTAIL.n156 VTAIL.n150 8.14595
R1570 VTAIL.n18 VTAIL.n12 8.14595
R1571 VTAIL.n115 VTAIL.n109 8.14595
R1572 VTAIL.n69 VTAIL.n63 8.14595
R1573 VTAIL.n155 VTAIL.n152 7.3702
R1574 VTAIL.n17 VTAIL.n14 7.3702
R1575 VTAIL.n114 VTAIL.n111 7.3702
R1576 VTAIL.n68 VTAIL.n65 7.3702
R1577 VTAIL.n156 VTAIL.n155 5.81868
R1578 VTAIL.n18 VTAIL.n17 5.81868
R1579 VTAIL.n115 VTAIL.n114 5.81868
R1580 VTAIL.n69 VTAIL.n68 5.81868
R1581 VTAIL.n159 VTAIL.n150 5.04292
R1582 VTAIL.n21 VTAIL.n12 5.04292
R1583 VTAIL.n118 VTAIL.n109 5.04292
R1584 VTAIL.n72 VTAIL.n63 5.04292
R1585 VTAIL.n160 VTAIL.n148 4.26717
R1586 VTAIL.n22 VTAIL.n10 4.26717
R1587 VTAIL.n119 VTAIL.n107 4.26717
R1588 VTAIL.n73 VTAIL.n61 4.26717
R1589 VTAIL.n164 VTAIL.n163 3.49141
R1590 VTAIL.n26 VTAIL.n25 3.49141
R1591 VTAIL.n123 VTAIL.n122 3.49141
R1592 VTAIL.n77 VTAIL.n76 3.49141
R1593 VTAIL.n154 VTAIL.n153 2.84304
R1594 VTAIL.n16 VTAIL.n15 2.84304
R1595 VTAIL.n113 VTAIL.n112 2.84304
R1596 VTAIL.n67 VTAIL.n66 2.84304
R1597 VTAIL.n167 VTAIL.n146 2.71565
R1598 VTAIL.n29 VTAIL.n8 2.71565
R1599 VTAIL.n126 VTAIL.n105 2.71565
R1600 VTAIL.n80 VTAIL.n59 2.71565
R1601 VTAIL.n182 VTAIL.t14 2.4817
R1602 VTAIL.n182 VTAIL.t15 2.4817
R1603 VTAIL.n0 VTAIL.t11 2.4817
R1604 VTAIL.n0 VTAIL.t12 2.4817
R1605 VTAIL.n44 VTAIL.t2 2.4817
R1606 VTAIL.n44 VTAIL.t6 2.4817
R1607 VTAIL.n46 VTAIL.t5 2.4817
R1608 VTAIL.n46 VTAIL.t0 2.4817
R1609 VTAIL.n96 VTAIL.t19 2.4817
R1610 VTAIL.n96 VTAIL.t4 2.4817
R1611 VTAIL.n94 VTAIL.t8 2.4817
R1612 VTAIL.n94 VTAIL.t3 2.4817
R1613 VTAIL.n50 VTAIL.t16 2.4817
R1614 VTAIL.n50 VTAIL.t17 2.4817
R1615 VTAIL.n48 VTAIL.t10 2.4817
R1616 VTAIL.n48 VTAIL.t18 2.4817
R1617 VTAIL.n168 VTAIL.n144 1.93989
R1618 VTAIL.n30 VTAIL.n6 1.93989
R1619 VTAIL.n127 VTAIL.n103 1.93989
R1620 VTAIL.n81 VTAIL.n57 1.93989
R1621 VTAIL.n51 VTAIL.n49 1.18153
R1622 VTAIL.n93 VTAIL.n51 1.18153
R1623 VTAIL.n97 VTAIL.n95 1.18153
R1624 VTAIL.n139 VTAIL.n97 1.18153
R1625 VTAIL.n47 VTAIL.n45 1.18153
R1626 VTAIL.n45 VTAIL.n43 1.18153
R1627 VTAIL.n183 VTAIL.n181 1.18153
R1628 VTAIL.n173 VTAIL.n171 1.16414
R1629 VTAIL.n180 VTAIL.n140 1.16414
R1630 VTAIL.n35 VTAIL.n33 1.16414
R1631 VTAIL.n42 VTAIL.n2 1.16414
R1632 VTAIL.n138 VTAIL.n98 1.16414
R1633 VTAIL.n131 VTAIL.n130 1.16414
R1634 VTAIL.n92 VTAIL.n52 1.16414
R1635 VTAIL.n85 VTAIL.n84 1.16414
R1636 VTAIL.n95 VTAIL.n93 1.06084
R1637 VTAIL.n43 VTAIL.n1 1.06084
R1638 VTAIL VTAIL.n1 0.944465
R1639 VTAIL.n172 VTAIL.n142 0.388379
R1640 VTAIL.n178 VTAIL.n177 0.388379
R1641 VTAIL.n34 VTAIL.n4 0.388379
R1642 VTAIL.n40 VTAIL.n39 0.388379
R1643 VTAIL.n136 VTAIL.n135 0.388379
R1644 VTAIL.n102 VTAIL.n100 0.388379
R1645 VTAIL.n90 VTAIL.n89 0.388379
R1646 VTAIL.n56 VTAIL.n54 0.388379
R1647 VTAIL VTAIL.n183 0.237569
R1648 VTAIL.n154 VTAIL.n149 0.155672
R1649 VTAIL.n161 VTAIL.n149 0.155672
R1650 VTAIL.n162 VTAIL.n161 0.155672
R1651 VTAIL.n162 VTAIL.n145 0.155672
R1652 VTAIL.n169 VTAIL.n145 0.155672
R1653 VTAIL.n170 VTAIL.n169 0.155672
R1654 VTAIL.n170 VTAIL.n141 0.155672
R1655 VTAIL.n179 VTAIL.n141 0.155672
R1656 VTAIL.n16 VTAIL.n11 0.155672
R1657 VTAIL.n23 VTAIL.n11 0.155672
R1658 VTAIL.n24 VTAIL.n23 0.155672
R1659 VTAIL.n24 VTAIL.n7 0.155672
R1660 VTAIL.n31 VTAIL.n7 0.155672
R1661 VTAIL.n32 VTAIL.n31 0.155672
R1662 VTAIL.n32 VTAIL.n3 0.155672
R1663 VTAIL.n41 VTAIL.n3 0.155672
R1664 VTAIL.n137 VTAIL.n99 0.155672
R1665 VTAIL.n129 VTAIL.n99 0.155672
R1666 VTAIL.n129 VTAIL.n128 0.155672
R1667 VTAIL.n128 VTAIL.n104 0.155672
R1668 VTAIL.n121 VTAIL.n104 0.155672
R1669 VTAIL.n121 VTAIL.n120 0.155672
R1670 VTAIL.n120 VTAIL.n108 0.155672
R1671 VTAIL.n113 VTAIL.n108 0.155672
R1672 VTAIL.n91 VTAIL.n53 0.155672
R1673 VTAIL.n83 VTAIL.n53 0.155672
R1674 VTAIL.n83 VTAIL.n82 0.155672
R1675 VTAIL.n82 VTAIL.n58 0.155672
R1676 VTAIL.n75 VTAIL.n58 0.155672
R1677 VTAIL.n75 VTAIL.n74 0.155672
R1678 VTAIL.n74 VTAIL.n62 0.155672
R1679 VTAIL.n67 VTAIL.n62 0.155672
R1680 VP.n9 VP.t5 238.131
R1681 VP.n25 VP.t2 223.157
R1682 VP.n41 VP.t9 223.157
R1683 VP.n22 VP.t4 223.157
R1684 VP.n26 VP.t0 184.922
R1685 VP.n33 VP.t7 184.922
R1686 VP.n39 VP.t1 184.922
R1687 VP.n20 VP.t6 184.922
R1688 VP.n14 VP.t3 184.922
R1689 VP.n8 VP.t8 184.922
R1690 VP.n10 VP.n7 161.3
R1691 VP.n12 VP.n11 161.3
R1692 VP.n13 VP.n6 161.3
R1693 VP.n16 VP.n15 161.3
R1694 VP.n17 VP.n5 161.3
R1695 VP.n19 VP.n18 161.3
R1696 VP.n21 VP.n4 161.3
R1697 VP.n40 VP.n0 161.3
R1698 VP.n38 VP.n37 161.3
R1699 VP.n36 VP.n1 161.3
R1700 VP.n35 VP.n34 161.3
R1701 VP.n32 VP.n2 161.3
R1702 VP.n31 VP.n30 161.3
R1703 VP.n29 VP.n3 161.3
R1704 VP.n28 VP.n27 161.3
R1705 VP.n23 VP.n22 80.6037
R1706 VP.n42 VP.n41 80.6037
R1707 VP.n25 VP.n24 80.6037
R1708 VP.n27 VP.n25 55.0167
R1709 VP.n41 VP.n40 55.0167
R1710 VP.n22 VP.n21 55.0167
R1711 VP.n9 VP.n8 48.3607
R1712 VP.n32 VP.n31 46.7399
R1713 VP.n34 VP.n1 46.7399
R1714 VP.n15 VP.n5 46.7399
R1715 VP.n13 VP.n12 46.7399
R1716 VP.n10 VP.n9 44.0902
R1717 VP.n24 VP.n23 41.8082
R1718 VP.n31 VP.n3 34.0813
R1719 VP.n38 VP.n1 34.0813
R1720 VP.n19 VP.n5 34.0813
R1721 VP.n12 VP.n7 34.0813
R1722 VP.n27 VP.n26 18.5015
R1723 VP.n40 VP.n39 18.5015
R1724 VP.n21 VP.n20 18.5015
R1725 VP.n33 VP.n32 12.1722
R1726 VP.n34 VP.n33 12.1722
R1727 VP.n14 VP.n13 12.1722
R1728 VP.n15 VP.n14 12.1722
R1729 VP.n26 VP.n3 5.84292
R1730 VP.n39 VP.n38 5.84292
R1731 VP.n20 VP.n19 5.84292
R1732 VP.n8 VP.n7 5.84292
R1733 VP.n23 VP.n4 0.285035
R1734 VP.n28 VP.n24 0.285035
R1735 VP.n42 VP.n0 0.285035
R1736 VP.n11 VP.n10 0.189894
R1737 VP.n11 VP.n6 0.189894
R1738 VP.n16 VP.n6 0.189894
R1739 VP.n17 VP.n16 0.189894
R1740 VP.n18 VP.n17 0.189894
R1741 VP.n18 VP.n4 0.189894
R1742 VP.n29 VP.n28 0.189894
R1743 VP.n30 VP.n29 0.189894
R1744 VP.n30 VP.n2 0.189894
R1745 VP.n35 VP.n2 0.189894
R1746 VP.n36 VP.n35 0.189894
R1747 VP.n37 VP.n36 0.189894
R1748 VP.n37 VP.n0 0.189894
R1749 VP VP.n42 0.146778
R1750 VDD1.n36 VDD1.n0 289.615
R1751 VDD1.n79 VDD1.n43 289.615
R1752 VDD1.n37 VDD1.n36 185
R1753 VDD1.n35 VDD1.n2 185
R1754 VDD1.n34 VDD1.n33 185
R1755 VDD1.n5 VDD1.n3 185
R1756 VDD1.n28 VDD1.n27 185
R1757 VDD1.n26 VDD1.n25 185
R1758 VDD1.n9 VDD1.n8 185
R1759 VDD1.n20 VDD1.n19 185
R1760 VDD1.n18 VDD1.n17 185
R1761 VDD1.n13 VDD1.n12 185
R1762 VDD1.n55 VDD1.n54 185
R1763 VDD1.n60 VDD1.n59 185
R1764 VDD1.n62 VDD1.n61 185
R1765 VDD1.n51 VDD1.n50 185
R1766 VDD1.n68 VDD1.n67 185
R1767 VDD1.n70 VDD1.n69 185
R1768 VDD1.n47 VDD1.n46 185
R1769 VDD1.n77 VDD1.n76 185
R1770 VDD1.n78 VDD1.n45 185
R1771 VDD1.n80 VDD1.n79 185
R1772 VDD1.n14 VDD1.t4 149.524
R1773 VDD1.n56 VDD1.t7 149.524
R1774 VDD1.n36 VDD1.n35 104.615
R1775 VDD1.n35 VDD1.n34 104.615
R1776 VDD1.n34 VDD1.n3 104.615
R1777 VDD1.n27 VDD1.n3 104.615
R1778 VDD1.n27 VDD1.n26 104.615
R1779 VDD1.n26 VDD1.n8 104.615
R1780 VDD1.n19 VDD1.n8 104.615
R1781 VDD1.n19 VDD1.n18 104.615
R1782 VDD1.n18 VDD1.n12 104.615
R1783 VDD1.n60 VDD1.n54 104.615
R1784 VDD1.n61 VDD1.n60 104.615
R1785 VDD1.n61 VDD1.n50 104.615
R1786 VDD1.n68 VDD1.n50 104.615
R1787 VDD1.n69 VDD1.n68 104.615
R1788 VDD1.n69 VDD1.n46 104.615
R1789 VDD1.n77 VDD1.n46 104.615
R1790 VDD1.n78 VDD1.n77 104.615
R1791 VDD1.n79 VDD1.n78 104.615
R1792 VDD1.n87 VDD1.n86 68.2991
R1793 VDD1.n42 VDD1.n41 67.4689
R1794 VDD1.n89 VDD1.n88 67.4687
R1795 VDD1.n85 VDD1.n84 67.4687
R1796 VDD1.n42 VDD1.n40 53.5361
R1797 VDD1.n85 VDD1.n83 53.5361
R1798 VDD1.t4 VDD1.n12 52.3082
R1799 VDD1.t7 VDD1.n54 52.3082
R1800 VDD1.n89 VDD1.n87 37.378
R1801 VDD1.n37 VDD1.n2 13.1884
R1802 VDD1.n80 VDD1.n45 13.1884
R1803 VDD1.n38 VDD1.n0 12.8005
R1804 VDD1.n33 VDD1.n4 12.8005
R1805 VDD1.n76 VDD1.n75 12.8005
R1806 VDD1.n81 VDD1.n43 12.8005
R1807 VDD1.n32 VDD1.n5 12.0247
R1808 VDD1.n74 VDD1.n47 12.0247
R1809 VDD1.n29 VDD1.n28 11.249
R1810 VDD1.n71 VDD1.n70 11.249
R1811 VDD1.n25 VDD1.n7 10.4732
R1812 VDD1.n67 VDD1.n49 10.4732
R1813 VDD1.n14 VDD1.n13 10.2747
R1814 VDD1.n56 VDD1.n55 10.2747
R1815 VDD1.n24 VDD1.n9 9.69747
R1816 VDD1.n66 VDD1.n51 9.69747
R1817 VDD1.n40 VDD1.n39 9.45567
R1818 VDD1.n83 VDD1.n82 9.45567
R1819 VDD1.n16 VDD1.n15 9.3005
R1820 VDD1.n11 VDD1.n10 9.3005
R1821 VDD1.n22 VDD1.n21 9.3005
R1822 VDD1.n24 VDD1.n23 9.3005
R1823 VDD1.n7 VDD1.n6 9.3005
R1824 VDD1.n30 VDD1.n29 9.3005
R1825 VDD1.n32 VDD1.n31 9.3005
R1826 VDD1.n4 VDD1.n1 9.3005
R1827 VDD1.n39 VDD1.n38 9.3005
R1828 VDD1.n82 VDD1.n81 9.3005
R1829 VDD1.n58 VDD1.n57 9.3005
R1830 VDD1.n53 VDD1.n52 9.3005
R1831 VDD1.n64 VDD1.n63 9.3005
R1832 VDD1.n66 VDD1.n65 9.3005
R1833 VDD1.n49 VDD1.n48 9.3005
R1834 VDD1.n72 VDD1.n71 9.3005
R1835 VDD1.n74 VDD1.n73 9.3005
R1836 VDD1.n75 VDD1.n44 9.3005
R1837 VDD1.n21 VDD1.n20 8.92171
R1838 VDD1.n63 VDD1.n62 8.92171
R1839 VDD1.n17 VDD1.n11 8.14595
R1840 VDD1.n59 VDD1.n53 8.14595
R1841 VDD1.n16 VDD1.n13 7.3702
R1842 VDD1.n58 VDD1.n55 7.3702
R1843 VDD1.n17 VDD1.n16 5.81868
R1844 VDD1.n59 VDD1.n58 5.81868
R1845 VDD1.n20 VDD1.n11 5.04292
R1846 VDD1.n62 VDD1.n53 5.04292
R1847 VDD1.n21 VDD1.n9 4.26717
R1848 VDD1.n63 VDD1.n51 4.26717
R1849 VDD1.n25 VDD1.n24 3.49141
R1850 VDD1.n67 VDD1.n66 3.49141
R1851 VDD1.n15 VDD1.n14 2.84304
R1852 VDD1.n57 VDD1.n56 2.84304
R1853 VDD1.n28 VDD1.n7 2.71565
R1854 VDD1.n70 VDD1.n49 2.71565
R1855 VDD1.n88 VDD1.t3 2.4817
R1856 VDD1.n88 VDD1.t5 2.4817
R1857 VDD1.n41 VDD1.t1 2.4817
R1858 VDD1.n41 VDD1.t6 2.4817
R1859 VDD1.n86 VDD1.t8 2.4817
R1860 VDD1.n86 VDD1.t0 2.4817
R1861 VDD1.n84 VDD1.t9 2.4817
R1862 VDD1.n84 VDD1.t2 2.4817
R1863 VDD1.n29 VDD1.n5 1.93989
R1864 VDD1.n71 VDD1.n47 1.93989
R1865 VDD1.n40 VDD1.n0 1.16414
R1866 VDD1.n33 VDD1.n32 1.16414
R1867 VDD1.n76 VDD1.n74 1.16414
R1868 VDD1.n83 VDD1.n43 1.16414
R1869 VDD1 VDD1.n89 0.828086
R1870 VDD1.n38 VDD1.n37 0.388379
R1871 VDD1.n4 VDD1.n2 0.388379
R1872 VDD1.n75 VDD1.n45 0.388379
R1873 VDD1.n81 VDD1.n80 0.388379
R1874 VDD1 VDD1.n42 0.353948
R1875 VDD1.n87 VDD1.n85 0.240413
R1876 VDD1.n39 VDD1.n1 0.155672
R1877 VDD1.n31 VDD1.n1 0.155672
R1878 VDD1.n31 VDD1.n30 0.155672
R1879 VDD1.n30 VDD1.n6 0.155672
R1880 VDD1.n23 VDD1.n6 0.155672
R1881 VDD1.n23 VDD1.n22 0.155672
R1882 VDD1.n22 VDD1.n10 0.155672
R1883 VDD1.n15 VDD1.n10 0.155672
R1884 VDD1.n57 VDD1.n52 0.155672
R1885 VDD1.n64 VDD1.n52 0.155672
R1886 VDD1.n65 VDD1.n64 0.155672
R1887 VDD1.n65 VDD1.n48 0.155672
R1888 VDD1.n72 VDD1.n48 0.155672
R1889 VDD1.n73 VDD1.n72 0.155672
R1890 VDD1.n73 VDD1.n44 0.155672
R1891 VDD1.n82 VDD1.n44 0.155672
C0 VP VTAIL 5.68331f
C1 VP VDD1 5.75376f
C2 VP VN 5.35585f
C3 VDD2 VTAIL 9.09546f
C4 VDD1 VDD2 1.18538f
C5 VDD1 VTAIL 9.05596f
C6 VDD2 VN 5.52244f
C7 VN VTAIL 5.66893f
C8 VDD1 VN 0.149409f
C9 VP VDD2 0.383892f
C10 VDD2 B 4.644681f
C11 VDD1 B 4.600157f
C12 VTAIL B 5.372356f
C13 VN B 10.537011f
C14 VP B 8.884112f
C15 VDD1.n0 B 0.032222f
C16 VDD1.n1 B 0.023604f
C17 VDD1.n2 B 0.013057f
C18 VDD1.n3 B 0.02998f
C19 VDD1.n4 B 0.012684f
C20 VDD1.n5 B 0.01343f
C21 VDD1.n6 B 0.023604f
C22 VDD1.n7 B 0.012684f
C23 VDD1.n8 B 0.02998f
C24 VDD1.n9 B 0.01343f
C25 VDD1.n10 B 0.023604f
C26 VDD1.n11 B 0.012684f
C27 VDD1.n12 B 0.022485f
C28 VDD1.n13 B 0.021194f
C29 VDD1.t4 B 0.050141f
C30 VDD1.n14 B 0.133786f
C31 VDD1.n15 B 0.768688f
C32 VDD1.n16 B 0.012684f
C33 VDD1.n17 B 0.01343f
C34 VDD1.n18 B 0.02998f
C35 VDD1.n19 B 0.02998f
C36 VDD1.n20 B 0.01343f
C37 VDD1.n21 B 0.012684f
C38 VDD1.n22 B 0.023604f
C39 VDD1.n23 B 0.023604f
C40 VDD1.n24 B 0.012684f
C41 VDD1.n25 B 0.01343f
C42 VDD1.n26 B 0.02998f
C43 VDD1.n27 B 0.02998f
C44 VDD1.n28 B 0.01343f
C45 VDD1.n29 B 0.012684f
C46 VDD1.n30 B 0.023604f
C47 VDD1.n31 B 0.023604f
C48 VDD1.n32 B 0.012684f
C49 VDD1.n33 B 0.01343f
C50 VDD1.n34 B 0.02998f
C51 VDD1.n35 B 0.02998f
C52 VDD1.n36 B 0.063212f
C53 VDD1.n37 B 0.013057f
C54 VDD1.n38 B 0.012684f
C55 VDD1.n39 B 0.060364f
C56 VDD1.n40 B 0.054681f
C57 VDD1.t1 B 0.148849f
C58 VDD1.t6 B 0.148849f
C59 VDD1.n41 B 1.2898f
C60 VDD1.n42 B 0.438834f
C61 VDD1.n43 B 0.032222f
C62 VDD1.n44 B 0.023604f
C63 VDD1.n45 B 0.013057f
C64 VDD1.n46 B 0.02998f
C65 VDD1.n47 B 0.01343f
C66 VDD1.n48 B 0.023604f
C67 VDD1.n49 B 0.012684f
C68 VDD1.n50 B 0.02998f
C69 VDD1.n51 B 0.01343f
C70 VDD1.n52 B 0.023604f
C71 VDD1.n53 B 0.012684f
C72 VDD1.n54 B 0.022485f
C73 VDD1.n55 B 0.021194f
C74 VDD1.t7 B 0.050141f
C75 VDD1.n56 B 0.133786f
C76 VDD1.n57 B 0.768688f
C77 VDD1.n58 B 0.012684f
C78 VDD1.n59 B 0.01343f
C79 VDD1.n60 B 0.02998f
C80 VDD1.n61 B 0.02998f
C81 VDD1.n62 B 0.01343f
C82 VDD1.n63 B 0.012684f
C83 VDD1.n64 B 0.023604f
C84 VDD1.n65 B 0.023604f
C85 VDD1.n66 B 0.012684f
C86 VDD1.n67 B 0.01343f
C87 VDD1.n68 B 0.02998f
C88 VDD1.n69 B 0.02998f
C89 VDD1.n70 B 0.01343f
C90 VDD1.n71 B 0.012684f
C91 VDD1.n72 B 0.023604f
C92 VDD1.n73 B 0.023604f
C93 VDD1.n74 B 0.012684f
C94 VDD1.n75 B 0.012684f
C95 VDD1.n76 B 0.01343f
C96 VDD1.n77 B 0.02998f
C97 VDD1.n78 B 0.02998f
C98 VDD1.n79 B 0.063212f
C99 VDD1.n80 B 0.013057f
C100 VDD1.n81 B 0.012684f
C101 VDD1.n82 B 0.060364f
C102 VDD1.n83 B 0.054681f
C103 VDD1.t9 B 0.148849f
C104 VDD1.t2 B 0.148849f
C105 VDD1.n84 B 1.2898f
C106 VDD1.n85 B 0.432486f
C107 VDD1.t8 B 0.148849f
C108 VDD1.t0 B 0.148849f
C109 VDD1.n86 B 1.29405f
C110 VDD1.n87 B 1.81073f
C111 VDD1.t3 B 0.148849f
C112 VDD1.t5 B 0.148849f
C113 VDD1.n88 B 1.2898f
C114 VDD1.n89 B 2.08165f
C115 VP.n0 B 0.050394f
C116 VP.t1 B 0.84168f
C117 VP.n1 B 0.032678f
C118 VP.n2 B 0.037766f
C119 VP.t7 B 0.84168f
C120 VP.n3 B 0.050182f
C121 VP.n4 B 0.050394f
C122 VP.t4 B 0.90222f
C123 VP.t6 B 0.84168f
C124 VP.n5 B 0.032678f
C125 VP.n6 B 0.037766f
C126 VP.t3 B 0.84168f
C127 VP.n7 B 0.050182f
C128 VP.t8 B 0.84168f
C129 VP.n8 B 0.360138f
C130 VP.t5 B 0.926707f
C131 VP.n9 B 0.385567f
C132 VP.n10 B 0.162371f
C133 VP.n11 B 0.037766f
C134 VP.n12 B 0.032678f
C135 VP.n13 B 0.054615f
C136 VP.n14 B 0.327717f
C137 VP.n15 B 0.054615f
C138 VP.n16 B 0.037766f
C139 VP.n17 B 0.037766f
C140 VP.n18 B 0.037766f
C141 VP.n19 B 0.050182f
C142 VP.n20 B 0.327717f
C143 VP.n21 B 0.052509f
C144 VP.n22 B 0.389165f
C145 VP.n23 B 1.56049f
C146 VP.n24 B 1.59287f
C147 VP.t2 B 0.90222f
C148 VP.n25 B 0.389165f
C149 VP.t0 B 0.84168f
C150 VP.n26 B 0.327717f
C151 VP.n27 B 0.052509f
C152 VP.n28 B 0.050394f
C153 VP.n29 B 0.037766f
C154 VP.n30 B 0.037766f
C155 VP.n31 B 0.032678f
C156 VP.n32 B 0.054615f
C157 VP.n33 B 0.327717f
C158 VP.n34 B 0.054615f
C159 VP.n35 B 0.037766f
C160 VP.n36 B 0.037766f
C161 VP.n37 B 0.037766f
C162 VP.n38 B 0.050182f
C163 VP.n39 B 0.327717f
C164 VP.n40 B 0.052509f
C165 VP.t9 B 0.90222f
C166 VP.n41 B 0.389165f
C167 VP.n42 B 0.035369f
C168 VTAIL.t11 B 0.163115f
C169 VTAIL.t12 B 0.163115f
C170 VTAIL.n0 B 1.34789f
C171 VTAIL.n1 B 0.401892f
C172 VTAIL.n2 B 0.03531f
C173 VTAIL.n3 B 0.025867f
C174 VTAIL.n4 B 0.014308f
C175 VTAIL.n5 B 0.032853f
C176 VTAIL.n6 B 0.014717f
C177 VTAIL.n7 B 0.025867f
C178 VTAIL.n8 B 0.013899f
C179 VTAIL.n9 B 0.032853f
C180 VTAIL.n10 B 0.014717f
C181 VTAIL.n11 B 0.025867f
C182 VTAIL.n12 B 0.013899f
C183 VTAIL.n13 B 0.02464f
C184 VTAIL.n14 B 0.023225f
C185 VTAIL.t1 B 0.054947f
C186 VTAIL.n15 B 0.146608f
C187 VTAIL.n16 B 0.842361f
C188 VTAIL.n17 B 0.013899f
C189 VTAIL.n18 B 0.014717f
C190 VTAIL.n19 B 0.032853f
C191 VTAIL.n20 B 0.032853f
C192 VTAIL.n21 B 0.014717f
C193 VTAIL.n22 B 0.013899f
C194 VTAIL.n23 B 0.025867f
C195 VTAIL.n24 B 0.025867f
C196 VTAIL.n25 B 0.013899f
C197 VTAIL.n26 B 0.014717f
C198 VTAIL.n27 B 0.032853f
C199 VTAIL.n28 B 0.032853f
C200 VTAIL.n29 B 0.014717f
C201 VTAIL.n30 B 0.013899f
C202 VTAIL.n31 B 0.025867f
C203 VTAIL.n32 B 0.025867f
C204 VTAIL.n33 B 0.013899f
C205 VTAIL.n34 B 0.013899f
C206 VTAIL.n35 B 0.014717f
C207 VTAIL.n36 B 0.032853f
C208 VTAIL.n37 B 0.032853f
C209 VTAIL.n38 B 0.06927f
C210 VTAIL.n39 B 0.014308f
C211 VTAIL.n40 B 0.013899f
C212 VTAIL.n41 B 0.06615f
C213 VTAIL.n42 B 0.038756f
C214 VTAIL.n43 B 0.212504f
C215 VTAIL.t2 B 0.163115f
C216 VTAIL.t6 B 0.163115f
C217 VTAIL.n44 B 1.34789f
C218 VTAIL.n45 B 0.43171f
C219 VTAIL.t5 B 0.163115f
C220 VTAIL.t0 B 0.163115f
C221 VTAIL.n46 B 1.34789f
C222 VTAIL.n47 B 1.45489f
C223 VTAIL.t10 B 0.163115f
C224 VTAIL.t18 B 0.163115f
C225 VTAIL.n48 B 1.34789f
C226 VTAIL.n49 B 1.45488f
C227 VTAIL.t16 B 0.163115f
C228 VTAIL.t17 B 0.163115f
C229 VTAIL.n50 B 1.34789f
C230 VTAIL.n51 B 0.431702f
C231 VTAIL.n52 B 0.03531f
C232 VTAIL.n53 B 0.025867f
C233 VTAIL.n54 B 0.014308f
C234 VTAIL.n55 B 0.032853f
C235 VTAIL.n56 B 0.013899f
C236 VTAIL.n57 B 0.014717f
C237 VTAIL.n58 B 0.025867f
C238 VTAIL.n59 B 0.013899f
C239 VTAIL.n60 B 0.032853f
C240 VTAIL.n61 B 0.014717f
C241 VTAIL.n62 B 0.025867f
C242 VTAIL.n63 B 0.013899f
C243 VTAIL.n64 B 0.02464f
C244 VTAIL.n65 B 0.023225f
C245 VTAIL.t13 B 0.054947f
C246 VTAIL.n66 B 0.146608f
C247 VTAIL.n67 B 0.842361f
C248 VTAIL.n68 B 0.013899f
C249 VTAIL.n69 B 0.014717f
C250 VTAIL.n70 B 0.032853f
C251 VTAIL.n71 B 0.032853f
C252 VTAIL.n72 B 0.014717f
C253 VTAIL.n73 B 0.013899f
C254 VTAIL.n74 B 0.025867f
C255 VTAIL.n75 B 0.025867f
C256 VTAIL.n76 B 0.013899f
C257 VTAIL.n77 B 0.014717f
C258 VTAIL.n78 B 0.032853f
C259 VTAIL.n79 B 0.032853f
C260 VTAIL.n80 B 0.014717f
C261 VTAIL.n81 B 0.013899f
C262 VTAIL.n82 B 0.025867f
C263 VTAIL.n83 B 0.025867f
C264 VTAIL.n84 B 0.013899f
C265 VTAIL.n85 B 0.014717f
C266 VTAIL.n86 B 0.032853f
C267 VTAIL.n87 B 0.032853f
C268 VTAIL.n88 B 0.06927f
C269 VTAIL.n89 B 0.014308f
C270 VTAIL.n90 B 0.013899f
C271 VTAIL.n91 B 0.06615f
C272 VTAIL.n92 B 0.038756f
C273 VTAIL.n93 B 0.212504f
C274 VTAIL.t8 B 0.163115f
C275 VTAIL.t3 B 0.163115f
C276 VTAIL.n94 B 1.34789f
C277 VTAIL.n95 B 0.421643f
C278 VTAIL.t19 B 0.163115f
C279 VTAIL.t4 B 0.163115f
C280 VTAIL.n96 B 1.34789f
C281 VTAIL.n97 B 0.431702f
C282 VTAIL.n98 B 0.03531f
C283 VTAIL.n99 B 0.025867f
C284 VTAIL.n100 B 0.014308f
C285 VTAIL.n101 B 0.032853f
C286 VTAIL.n102 B 0.013899f
C287 VTAIL.n103 B 0.014717f
C288 VTAIL.n104 B 0.025867f
C289 VTAIL.n105 B 0.013899f
C290 VTAIL.n106 B 0.032853f
C291 VTAIL.n107 B 0.014717f
C292 VTAIL.n108 B 0.025867f
C293 VTAIL.n109 B 0.013899f
C294 VTAIL.n110 B 0.02464f
C295 VTAIL.n111 B 0.023225f
C296 VTAIL.t7 B 0.054947f
C297 VTAIL.n112 B 0.146608f
C298 VTAIL.n113 B 0.842361f
C299 VTAIL.n114 B 0.013899f
C300 VTAIL.n115 B 0.014717f
C301 VTAIL.n116 B 0.032853f
C302 VTAIL.n117 B 0.032853f
C303 VTAIL.n118 B 0.014717f
C304 VTAIL.n119 B 0.013899f
C305 VTAIL.n120 B 0.025867f
C306 VTAIL.n121 B 0.025867f
C307 VTAIL.n122 B 0.013899f
C308 VTAIL.n123 B 0.014717f
C309 VTAIL.n124 B 0.032853f
C310 VTAIL.n125 B 0.032853f
C311 VTAIL.n126 B 0.014717f
C312 VTAIL.n127 B 0.013899f
C313 VTAIL.n128 B 0.025867f
C314 VTAIL.n129 B 0.025867f
C315 VTAIL.n130 B 0.013899f
C316 VTAIL.n131 B 0.014717f
C317 VTAIL.n132 B 0.032853f
C318 VTAIL.n133 B 0.032853f
C319 VTAIL.n134 B 0.06927f
C320 VTAIL.n135 B 0.014308f
C321 VTAIL.n136 B 0.013899f
C322 VTAIL.n137 B 0.06615f
C323 VTAIL.n138 B 0.038756f
C324 VTAIL.n139 B 1.1473f
C325 VTAIL.n140 B 0.03531f
C326 VTAIL.n141 B 0.025867f
C327 VTAIL.n142 B 0.014308f
C328 VTAIL.n143 B 0.032853f
C329 VTAIL.n144 B 0.014717f
C330 VTAIL.n145 B 0.025867f
C331 VTAIL.n146 B 0.013899f
C332 VTAIL.n147 B 0.032853f
C333 VTAIL.n148 B 0.014717f
C334 VTAIL.n149 B 0.025867f
C335 VTAIL.n150 B 0.013899f
C336 VTAIL.n151 B 0.02464f
C337 VTAIL.n152 B 0.023225f
C338 VTAIL.t9 B 0.054947f
C339 VTAIL.n153 B 0.146608f
C340 VTAIL.n154 B 0.842361f
C341 VTAIL.n155 B 0.013899f
C342 VTAIL.n156 B 0.014717f
C343 VTAIL.n157 B 0.032853f
C344 VTAIL.n158 B 0.032853f
C345 VTAIL.n159 B 0.014717f
C346 VTAIL.n160 B 0.013899f
C347 VTAIL.n161 B 0.025867f
C348 VTAIL.n162 B 0.025867f
C349 VTAIL.n163 B 0.013899f
C350 VTAIL.n164 B 0.014717f
C351 VTAIL.n165 B 0.032853f
C352 VTAIL.n166 B 0.032853f
C353 VTAIL.n167 B 0.014717f
C354 VTAIL.n168 B 0.013899f
C355 VTAIL.n169 B 0.025867f
C356 VTAIL.n170 B 0.025867f
C357 VTAIL.n171 B 0.013899f
C358 VTAIL.n172 B 0.013899f
C359 VTAIL.n173 B 0.014717f
C360 VTAIL.n174 B 0.032853f
C361 VTAIL.n175 B 0.032853f
C362 VTAIL.n176 B 0.06927f
C363 VTAIL.n177 B 0.014308f
C364 VTAIL.n178 B 0.013899f
C365 VTAIL.n179 B 0.06615f
C366 VTAIL.n180 B 0.038756f
C367 VTAIL.n181 B 1.1473f
C368 VTAIL.t14 B 0.163115f
C369 VTAIL.t15 B 0.163115f
C370 VTAIL.n182 B 1.34789f
C371 VTAIL.n183 B 0.353033f
C372 VDD2.n0 B 0.031759f
C373 VDD2.n1 B 0.023265f
C374 VDD2.n2 B 0.012869f
C375 VDD2.n3 B 0.029549f
C376 VDD2.n4 B 0.013237f
C377 VDD2.n5 B 0.023265f
C378 VDD2.n6 B 0.012502f
C379 VDD2.n7 B 0.029549f
C380 VDD2.n8 B 0.013237f
C381 VDD2.n9 B 0.023265f
C382 VDD2.n10 B 0.012502f
C383 VDD2.n11 B 0.022162f
C384 VDD2.n12 B 0.020889f
C385 VDD2.t3 B 0.049421f
C386 VDD2.n13 B 0.131863f
C387 VDD2.n14 B 0.757644f
C388 VDD2.n15 B 0.012502f
C389 VDD2.n16 B 0.013237f
C390 VDD2.n17 B 0.029549f
C391 VDD2.n18 B 0.029549f
C392 VDD2.n19 B 0.013237f
C393 VDD2.n20 B 0.012502f
C394 VDD2.n21 B 0.023265f
C395 VDD2.n22 B 0.023265f
C396 VDD2.n23 B 0.012502f
C397 VDD2.n24 B 0.013237f
C398 VDD2.n25 B 0.029549f
C399 VDD2.n26 B 0.029549f
C400 VDD2.n27 B 0.013237f
C401 VDD2.n28 B 0.012502f
C402 VDD2.n29 B 0.023265f
C403 VDD2.n30 B 0.023265f
C404 VDD2.n31 B 0.012502f
C405 VDD2.n32 B 0.012502f
C406 VDD2.n33 B 0.013237f
C407 VDD2.n34 B 0.029549f
C408 VDD2.n35 B 0.029549f
C409 VDD2.n36 B 0.062304f
C410 VDD2.n37 B 0.012869f
C411 VDD2.n38 B 0.012502f
C412 VDD2.n39 B 0.059497f
C413 VDD2.n40 B 0.053896f
C414 VDD2.t9 B 0.14671f
C415 VDD2.t8 B 0.14671f
C416 VDD2.n41 B 1.27127f
C417 VDD2.n42 B 0.426272f
C418 VDD2.t5 B 0.14671f
C419 VDD2.t0 B 0.14671f
C420 VDD2.n43 B 1.27546f
C421 VDD2.n44 B 1.70728f
C422 VDD2.n45 B 0.031759f
C423 VDD2.n46 B 0.023265f
C424 VDD2.n47 B 0.012869f
C425 VDD2.n48 B 0.029549f
C426 VDD2.n49 B 0.012502f
C427 VDD2.n50 B 0.013237f
C428 VDD2.n51 B 0.023265f
C429 VDD2.n52 B 0.012502f
C430 VDD2.n53 B 0.029549f
C431 VDD2.n54 B 0.013237f
C432 VDD2.n55 B 0.023265f
C433 VDD2.n56 B 0.012502f
C434 VDD2.n57 B 0.022162f
C435 VDD2.n58 B 0.020889f
C436 VDD2.t2 B 0.049421f
C437 VDD2.n59 B 0.131863f
C438 VDD2.n60 B 0.757644f
C439 VDD2.n61 B 0.012502f
C440 VDD2.n62 B 0.013237f
C441 VDD2.n63 B 0.029549f
C442 VDD2.n64 B 0.029549f
C443 VDD2.n65 B 0.013237f
C444 VDD2.n66 B 0.012502f
C445 VDD2.n67 B 0.023265f
C446 VDD2.n68 B 0.023265f
C447 VDD2.n69 B 0.012502f
C448 VDD2.n70 B 0.013237f
C449 VDD2.n71 B 0.029549f
C450 VDD2.n72 B 0.029549f
C451 VDD2.n73 B 0.013237f
C452 VDD2.n74 B 0.012502f
C453 VDD2.n75 B 0.023265f
C454 VDD2.n76 B 0.023265f
C455 VDD2.n77 B 0.012502f
C456 VDD2.n78 B 0.013237f
C457 VDD2.n79 B 0.029549f
C458 VDD2.n80 B 0.029549f
C459 VDD2.n81 B 0.062304f
C460 VDD2.n82 B 0.012869f
C461 VDD2.n83 B 0.012502f
C462 VDD2.n84 B 0.059497f
C463 VDD2.n85 B 0.050882f
C464 VDD2.n86 B 1.836f
C465 VDD2.t6 B 0.14671f
C466 VDD2.t4 B 0.14671f
C467 VDD2.n87 B 1.27127f
C468 VDD2.n88 B 0.298932f
C469 VDD2.t7 B 0.14671f
C470 VDD2.t1 B 0.14671f
C471 VDD2.n89 B 1.27543f
C472 VN.n0 B 0.049344f
C473 VN.t3 B 0.82415f
C474 VN.n1 B 0.031997f
C475 VN.n2 B 0.036979f
C476 VN.t4 B 0.82415f
C477 VN.n3 B 0.049137f
C478 VN.t7 B 0.907406f
C479 VN.t6 B 0.82415f
C480 VN.n4 B 0.352637f
C481 VN.n5 B 0.377537f
C482 VN.n6 B 0.158989f
C483 VN.n7 B 0.036979f
C484 VN.n8 B 0.031997f
C485 VN.n9 B 0.053477f
C486 VN.n10 B 0.320891f
C487 VN.n11 B 0.053477f
C488 VN.n12 B 0.036979f
C489 VN.n13 B 0.036979f
C490 VN.n14 B 0.036979f
C491 VN.n15 B 0.049137f
C492 VN.n16 B 0.320891f
C493 VN.n17 B 0.051416f
C494 VN.t9 B 0.883429f
C495 VN.n18 B 0.38106f
C496 VN.n19 B 0.034633f
C497 VN.n20 B 0.049344f
C498 VN.t0 B 0.82415f
C499 VN.n21 B 0.031997f
C500 VN.n22 B 0.036979f
C501 VN.t2 B 0.82415f
C502 VN.n23 B 0.049137f
C503 VN.t5 B 0.907406f
C504 VN.t1 B 0.82415f
C505 VN.n24 B 0.352637f
C506 VN.n25 B 0.377537f
C507 VN.n26 B 0.158989f
C508 VN.n27 B 0.036979f
C509 VN.n28 B 0.031997f
C510 VN.n29 B 0.053477f
C511 VN.n30 B 0.320891f
C512 VN.n31 B 0.053477f
C513 VN.n32 B 0.036979f
C514 VN.n33 B 0.036979f
C515 VN.n34 B 0.036979f
C516 VN.n35 B 0.049137f
C517 VN.n36 B 0.320891f
C518 VN.n37 B 0.051416f
C519 VN.t8 B 0.883429f
C520 VN.n38 B 0.38106f
C521 VN.n39 B 1.54875f
.ends

