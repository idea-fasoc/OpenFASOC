* NGSPICE file created from diff_pair_sample_0634.ext - technology: sky130A

.subckt diff_pair_sample_0634 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2102_n1302# sky130_fd_pr__pfet_01v8 ad=0.6513 pd=4.12 as=0 ps=0 w=1.67 l=2.5
X1 B.t8 B.t6 B.t7 w_n2102_n1302# sky130_fd_pr__pfet_01v8 ad=0.6513 pd=4.12 as=0 ps=0 w=1.67 l=2.5
X2 B.t5 B.t3 B.t4 w_n2102_n1302# sky130_fd_pr__pfet_01v8 ad=0.6513 pd=4.12 as=0 ps=0 w=1.67 l=2.5
X3 VDD2.t1 VN.t0 VTAIL.t3 w_n2102_n1302# sky130_fd_pr__pfet_01v8 ad=0.6513 pd=4.12 as=0.6513 ps=4.12 w=1.67 l=2.5
X4 VDD2.t0 VN.t1 VTAIL.t2 w_n2102_n1302# sky130_fd_pr__pfet_01v8 ad=0.6513 pd=4.12 as=0.6513 ps=4.12 w=1.67 l=2.5
X5 VDD1.t1 VP.t0 VTAIL.t0 w_n2102_n1302# sky130_fd_pr__pfet_01v8 ad=0.6513 pd=4.12 as=0.6513 ps=4.12 w=1.67 l=2.5
X6 B.t2 B.t0 B.t1 w_n2102_n1302# sky130_fd_pr__pfet_01v8 ad=0.6513 pd=4.12 as=0 ps=0 w=1.67 l=2.5
X7 VDD1.t0 VP.t1 VTAIL.t1 w_n2102_n1302# sky130_fd_pr__pfet_01v8 ad=0.6513 pd=4.12 as=0.6513 ps=4.12 w=1.67 l=2.5
R0 B.n175 B.n60 585
R1 B.n174 B.n173 585
R2 B.n172 B.n61 585
R3 B.n171 B.n170 585
R4 B.n169 B.n62 585
R5 B.n168 B.n167 585
R6 B.n166 B.n63 585
R7 B.n165 B.n164 585
R8 B.n163 B.n64 585
R9 B.n162 B.n161 585
R10 B.n160 B.n65 585
R11 B.n159 B.n158 585
R12 B.n154 B.n66 585
R13 B.n153 B.n152 585
R14 B.n151 B.n67 585
R15 B.n150 B.n149 585
R16 B.n148 B.n68 585
R17 B.n147 B.n146 585
R18 B.n145 B.n69 585
R19 B.n144 B.n143 585
R20 B.n142 B.n70 585
R21 B.n140 B.n139 585
R22 B.n138 B.n73 585
R23 B.n137 B.n136 585
R24 B.n135 B.n74 585
R25 B.n134 B.n133 585
R26 B.n132 B.n75 585
R27 B.n131 B.n130 585
R28 B.n129 B.n76 585
R29 B.n128 B.n127 585
R30 B.n126 B.n77 585
R31 B.n125 B.n124 585
R32 B.n177 B.n176 585
R33 B.n178 B.n59 585
R34 B.n180 B.n179 585
R35 B.n181 B.n58 585
R36 B.n183 B.n182 585
R37 B.n184 B.n57 585
R38 B.n186 B.n185 585
R39 B.n187 B.n56 585
R40 B.n189 B.n188 585
R41 B.n190 B.n55 585
R42 B.n192 B.n191 585
R43 B.n193 B.n54 585
R44 B.n195 B.n194 585
R45 B.n196 B.n53 585
R46 B.n198 B.n197 585
R47 B.n199 B.n52 585
R48 B.n201 B.n200 585
R49 B.n202 B.n51 585
R50 B.n204 B.n203 585
R51 B.n205 B.n50 585
R52 B.n207 B.n206 585
R53 B.n208 B.n49 585
R54 B.n210 B.n209 585
R55 B.n211 B.n48 585
R56 B.n213 B.n212 585
R57 B.n214 B.n47 585
R58 B.n216 B.n215 585
R59 B.n217 B.n46 585
R60 B.n219 B.n218 585
R61 B.n220 B.n45 585
R62 B.n222 B.n221 585
R63 B.n223 B.n44 585
R64 B.n225 B.n224 585
R65 B.n226 B.n43 585
R66 B.n228 B.n227 585
R67 B.n229 B.n42 585
R68 B.n231 B.n230 585
R69 B.n232 B.n41 585
R70 B.n234 B.n233 585
R71 B.n235 B.n40 585
R72 B.n237 B.n236 585
R73 B.n238 B.n39 585
R74 B.n240 B.n239 585
R75 B.n241 B.n38 585
R76 B.n243 B.n242 585
R77 B.n244 B.n37 585
R78 B.n246 B.n245 585
R79 B.n247 B.n36 585
R80 B.n249 B.n248 585
R81 B.n250 B.n35 585
R82 B.n299 B.n14 585
R83 B.n298 B.n297 585
R84 B.n296 B.n15 585
R85 B.n295 B.n294 585
R86 B.n293 B.n16 585
R87 B.n292 B.n291 585
R88 B.n290 B.n17 585
R89 B.n289 B.n288 585
R90 B.n287 B.n18 585
R91 B.n286 B.n285 585
R92 B.n284 B.n19 585
R93 B.n282 B.n281 585
R94 B.n280 B.n22 585
R95 B.n279 B.n278 585
R96 B.n277 B.n23 585
R97 B.n276 B.n275 585
R98 B.n274 B.n24 585
R99 B.n273 B.n272 585
R100 B.n271 B.n25 585
R101 B.n270 B.n269 585
R102 B.n268 B.n26 585
R103 B.n267 B.n266 585
R104 B.n265 B.n27 585
R105 B.n264 B.n263 585
R106 B.n262 B.n31 585
R107 B.n261 B.n260 585
R108 B.n259 B.n32 585
R109 B.n258 B.n257 585
R110 B.n256 B.n33 585
R111 B.n255 B.n254 585
R112 B.n253 B.n34 585
R113 B.n252 B.n251 585
R114 B.n301 B.n300 585
R115 B.n302 B.n13 585
R116 B.n304 B.n303 585
R117 B.n305 B.n12 585
R118 B.n307 B.n306 585
R119 B.n308 B.n11 585
R120 B.n310 B.n309 585
R121 B.n311 B.n10 585
R122 B.n313 B.n312 585
R123 B.n314 B.n9 585
R124 B.n316 B.n315 585
R125 B.n317 B.n8 585
R126 B.n319 B.n318 585
R127 B.n320 B.n7 585
R128 B.n322 B.n321 585
R129 B.n323 B.n6 585
R130 B.n325 B.n324 585
R131 B.n326 B.n5 585
R132 B.n328 B.n327 585
R133 B.n329 B.n4 585
R134 B.n331 B.n330 585
R135 B.n332 B.n3 585
R136 B.n334 B.n333 585
R137 B.n335 B.n0 585
R138 B.n2 B.n1 585
R139 B.n90 B.n89 585
R140 B.n92 B.n91 585
R141 B.n93 B.n88 585
R142 B.n95 B.n94 585
R143 B.n96 B.n87 585
R144 B.n98 B.n97 585
R145 B.n99 B.n86 585
R146 B.n101 B.n100 585
R147 B.n102 B.n85 585
R148 B.n104 B.n103 585
R149 B.n105 B.n84 585
R150 B.n107 B.n106 585
R151 B.n108 B.n83 585
R152 B.n110 B.n109 585
R153 B.n111 B.n82 585
R154 B.n113 B.n112 585
R155 B.n114 B.n81 585
R156 B.n116 B.n115 585
R157 B.n117 B.n80 585
R158 B.n119 B.n118 585
R159 B.n120 B.n79 585
R160 B.n122 B.n121 585
R161 B.n123 B.n78 585
R162 B.n125 B.n78 545.355
R163 B.n177 B.n60 545.355
R164 B.n251 B.n250 545.355
R165 B.n300 B.n299 545.355
R166 B.n155 B.t10 305.423
R167 B.n28 B.t8 305.423
R168 B.n71 B.t1 305.423
R169 B.n20 B.t5 305.423
R170 B.n337 B.n336 256.663
R171 B.n156 B.t11 250.538
R172 B.n29 B.t7 250.538
R173 B.n72 B.t2 250.538
R174 B.n21 B.t4 250.538
R175 B.n336 B.n335 235.042
R176 B.n336 B.n2 235.042
R177 B.n71 B.t0 223.989
R178 B.n155 B.t9 223.989
R179 B.n28 B.t6 223.989
R180 B.n20 B.t3 223.989
R181 B.n126 B.n125 163.367
R182 B.n127 B.n126 163.367
R183 B.n127 B.n76 163.367
R184 B.n131 B.n76 163.367
R185 B.n132 B.n131 163.367
R186 B.n133 B.n132 163.367
R187 B.n133 B.n74 163.367
R188 B.n137 B.n74 163.367
R189 B.n138 B.n137 163.367
R190 B.n139 B.n138 163.367
R191 B.n139 B.n70 163.367
R192 B.n144 B.n70 163.367
R193 B.n145 B.n144 163.367
R194 B.n146 B.n145 163.367
R195 B.n146 B.n68 163.367
R196 B.n150 B.n68 163.367
R197 B.n151 B.n150 163.367
R198 B.n152 B.n151 163.367
R199 B.n152 B.n66 163.367
R200 B.n159 B.n66 163.367
R201 B.n160 B.n159 163.367
R202 B.n161 B.n160 163.367
R203 B.n161 B.n64 163.367
R204 B.n165 B.n64 163.367
R205 B.n166 B.n165 163.367
R206 B.n167 B.n166 163.367
R207 B.n167 B.n62 163.367
R208 B.n171 B.n62 163.367
R209 B.n172 B.n171 163.367
R210 B.n173 B.n172 163.367
R211 B.n173 B.n60 163.367
R212 B.n250 B.n249 163.367
R213 B.n249 B.n36 163.367
R214 B.n245 B.n36 163.367
R215 B.n245 B.n244 163.367
R216 B.n244 B.n243 163.367
R217 B.n243 B.n38 163.367
R218 B.n239 B.n38 163.367
R219 B.n239 B.n238 163.367
R220 B.n238 B.n237 163.367
R221 B.n237 B.n40 163.367
R222 B.n233 B.n40 163.367
R223 B.n233 B.n232 163.367
R224 B.n232 B.n231 163.367
R225 B.n231 B.n42 163.367
R226 B.n227 B.n42 163.367
R227 B.n227 B.n226 163.367
R228 B.n226 B.n225 163.367
R229 B.n225 B.n44 163.367
R230 B.n221 B.n44 163.367
R231 B.n221 B.n220 163.367
R232 B.n220 B.n219 163.367
R233 B.n219 B.n46 163.367
R234 B.n215 B.n46 163.367
R235 B.n215 B.n214 163.367
R236 B.n214 B.n213 163.367
R237 B.n213 B.n48 163.367
R238 B.n209 B.n48 163.367
R239 B.n209 B.n208 163.367
R240 B.n208 B.n207 163.367
R241 B.n207 B.n50 163.367
R242 B.n203 B.n50 163.367
R243 B.n203 B.n202 163.367
R244 B.n202 B.n201 163.367
R245 B.n201 B.n52 163.367
R246 B.n197 B.n52 163.367
R247 B.n197 B.n196 163.367
R248 B.n196 B.n195 163.367
R249 B.n195 B.n54 163.367
R250 B.n191 B.n54 163.367
R251 B.n191 B.n190 163.367
R252 B.n190 B.n189 163.367
R253 B.n189 B.n56 163.367
R254 B.n185 B.n56 163.367
R255 B.n185 B.n184 163.367
R256 B.n184 B.n183 163.367
R257 B.n183 B.n58 163.367
R258 B.n179 B.n58 163.367
R259 B.n179 B.n178 163.367
R260 B.n178 B.n177 163.367
R261 B.n299 B.n298 163.367
R262 B.n298 B.n15 163.367
R263 B.n294 B.n15 163.367
R264 B.n294 B.n293 163.367
R265 B.n293 B.n292 163.367
R266 B.n292 B.n17 163.367
R267 B.n288 B.n17 163.367
R268 B.n288 B.n287 163.367
R269 B.n287 B.n286 163.367
R270 B.n286 B.n19 163.367
R271 B.n281 B.n19 163.367
R272 B.n281 B.n280 163.367
R273 B.n280 B.n279 163.367
R274 B.n279 B.n23 163.367
R275 B.n275 B.n23 163.367
R276 B.n275 B.n274 163.367
R277 B.n274 B.n273 163.367
R278 B.n273 B.n25 163.367
R279 B.n269 B.n25 163.367
R280 B.n269 B.n268 163.367
R281 B.n268 B.n267 163.367
R282 B.n267 B.n27 163.367
R283 B.n263 B.n27 163.367
R284 B.n263 B.n262 163.367
R285 B.n262 B.n261 163.367
R286 B.n261 B.n32 163.367
R287 B.n257 B.n32 163.367
R288 B.n257 B.n256 163.367
R289 B.n256 B.n255 163.367
R290 B.n255 B.n34 163.367
R291 B.n251 B.n34 163.367
R292 B.n300 B.n13 163.367
R293 B.n304 B.n13 163.367
R294 B.n305 B.n304 163.367
R295 B.n306 B.n305 163.367
R296 B.n306 B.n11 163.367
R297 B.n310 B.n11 163.367
R298 B.n311 B.n310 163.367
R299 B.n312 B.n311 163.367
R300 B.n312 B.n9 163.367
R301 B.n316 B.n9 163.367
R302 B.n317 B.n316 163.367
R303 B.n318 B.n317 163.367
R304 B.n318 B.n7 163.367
R305 B.n322 B.n7 163.367
R306 B.n323 B.n322 163.367
R307 B.n324 B.n323 163.367
R308 B.n324 B.n5 163.367
R309 B.n328 B.n5 163.367
R310 B.n329 B.n328 163.367
R311 B.n330 B.n329 163.367
R312 B.n330 B.n3 163.367
R313 B.n334 B.n3 163.367
R314 B.n335 B.n334 163.367
R315 B.n90 B.n2 163.367
R316 B.n91 B.n90 163.367
R317 B.n91 B.n88 163.367
R318 B.n95 B.n88 163.367
R319 B.n96 B.n95 163.367
R320 B.n97 B.n96 163.367
R321 B.n97 B.n86 163.367
R322 B.n101 B.n86 163.367
R323 B.n102 B.n101 163.367
R324 B.n103 B.n102 163.367
R325 B.n103 B.n84 163.367
R326 B.n107 B.n84 163.367
R327 B.n108 B.n107 163.367
R328 B.n109 B.n108 163.367
R329 B.n109 B.n82 163.367
R330 B.n113 B.n82 163.367
R331 B.n114 B.n113 163.367
R332 B.n115 B.n114 163.367
R333 B.n115 B.n80 163.367
R334 B.n119 B.n80 163.367
R335 B.n120 B.n119 163.367
R336 B.n121 B.n120 163.367
R337 B.n121 B.n78 163.367
R338 B.n141 B.n72 59.5399
R339 B.n157 B.n156 59.5399
R340 B.n30 B.n29 59.5399
R341 B.n283 B.n21 59.5399
R342 B.n72 B.n71 54.8853
R343 B.n156 B.n155 54.8853
R344 B.n29 B.n28 54.8853
R345 B.n21 B.n20 54.8853
R346 B.n301 B.n14 35.4346
R347 B.n252 B.n35 35.4346
R348 B.n176 B.n175 35.4346
R349 B.n124 B.n123 35.4346
R350 B B.n337 18.0485
R351 B.n302 B.n301 10.6151
R352 B.n303 B.n302 10.6151
R353 B.n303 B.n12 10.6151
R354 B.n307 B.n12 10.6151
R355 B.n308 B.n307 10.6151
R356 B.n309 B.n308 10.6151
R357 B.n309 B.n10 10.6151
R358 B.n313 B.n10 10.6151
R359 B.n314 B.n313 10.6151
R360 B.n315 B.n314 10.6151
R361 B.n315 B.n8 10.6151
R362 B.n319 B.n8 10.6151
R363 B.n320 B.n319 10.6151
R364 B.n321 B.n320 10.6151
R365 B.n321 B.n6 10.6151
R366 B.n325 B.n6 10.6151
R367 B.n326 B.n325 10.6151
R368 B.n327 B.n326 10.6151
R369 B.n327 B.n4 10.6151
R370 B.n331 B.n4 10.6151
R371 B.n332 B.n331 10.6151
R372 B.n333 B.n332 10.6151
R373 B.n333 B.n0 10.6151
R374 B.n297 B.n14 10.6151
R375 B.n297 B.n296 10.6151
R376 B.n296 B.n295 10.6151
R377 B.n295 B.n16 10.6151
R378 B.n291 B.n16 10.6151
R379 B.n291 B.n290 10.6151
R380 B.n290 B.n289 10.6151
R381 B.n289 B.n18 10.6151
R382 B.n285 B.n18 10.6151
R383 B.n285 B.n284 10.6151
R384 B.n282 B.n22 10.6151
R385 B.n278 B.n22 10.6151
R386 B.n278 B.n277 10.6151
R387 B.n277 B.n276 10.6151
R388 B.n276 B.n24 10.6151
R389 B.n272 B.n24 10.6151
R390 B.n272 B.n271 10.6151
R391 B.n271 B.n270 10.6151
R392 B.n270 B.n26 10.6151
R393 B.n266 B.n265 10.6151
R394 B.n265 B.n264 10.6151
R395 B.n264 B.n31 10.6151
R396 B.n260 B.n31 10.6151
R397 B.n260 B.n259 10.6151
R398 B.n259 B.n258 10.6151
R399 B.n258 B.n33 10.6151
R400 B.n254 B.n33 10.6151
R401 B.n254 B.n253 10.6151
R402 B.n253 B.n252 10.6151
R403 B.n248 B.n35 10.6151
R404 B.n248 B.n247 10.6151
R405 B.n247 B.n246 10.6151
R406 B.n246 B.n37 10.6151
R407 B.n242 B.n37 10.6151
R408 B.n242 B.n241 10.6151
R409 B.n241 B.n240 10.6151
R410 B.n240 B.n39 10.6151
R411 B.n236 B.n39 10.6151
R412 B.n236 B.n235 10.6151
R413 B.n235 B.n234 10.6151
R414 B.n234 B.n41 10.6151
R415 B.n230 B.n41 10.6151
R416 B.n230 B.n229 10.6151
R417 B.n229 B.n228 10.6151
R418 B.n228 B.n43 10.6151
R419 B.n224 B.n43 10.6151
R420 B.n224 B.n223 10.6151
R421 B.n223 B.n222 10.6151
R422 B.n222 B.n45 10.6151
R423 B.n218 B.n45 10.6151
R424 B.n218 B.n217 10.6151
R425 B.n217 B.n216 10.6151
R426 B.n216 B.n47 10.6151
R427 B.n212 B.n47 10.6151
R428 B.n212 B.n211 10.6151
R429 B.n211 B.n210 10.6151
R430 B.n210 B.n49 10.6151
R431 B.n206 B.n49 10.6151
R432 B.n206 B.n205 10.6151
R433 B.n205 B.n204 10.6151
R434 B.n204 B.n51 10.6151
R435 B.n200 B.n51 10.6151
R436 B.n200 B.n199 10.6151
R437 B.n199 B.n198 10.6151
R438 B.n198 B.n53 10.6151
R439 B.n194 B.n53 10.6151
R440 B.n194 B.n193 10.6151
R441 B.n193 B.n192 10.6151
R442 B.n192 B.n55 10.6151
R443 B.n188 B.n55 10.6151
R444 B.n188 B.n187 10.6151
R445 B.n187 B.n186 10.6151
R446 B.n186 B.n57 10.6151
R447 B.n182 B.n57 10.6151
R448 B.n182 B.n181 10.6151
R449 B.n181 B.n180 10.6151
R450 B.n180 B.n59 10.6151
R451 B.n176 B.n59 10.6151
R452 B.n89 B.n1 10.6151
R453 B.n92 B.n89 10.6151
R454 B.n93 B.n92 10.6151
R455 B.n94 B.n93 10.6151
R456 B.n94 B.n87 10.6151
R457 B.n98 B.n87 10.6151
R458 B.n99 B.n98 10.6151
R459 B.n100 B.n99 10.6151
R460 B.n100 B.n85 10.6151
R461 B.n104 B.n85 10.6151
R462 B.n105 B.n104 10.6151
R463 B.n106 B.n105 10.6151
R464 B.n106 B.n83 10.6151
R465 B.n110 B.n83 10.6151
R466 B.n111 B.n110 10.6151
R467 B.n112 B.n111 10.6151
R468 B.n112 B.n81 10.6151
R469 B.n116 B.n81 10.6151
R470 B.n117 B.n116 10.6151
R471 B.n118 B.n117 10.6151
R472 B.n118 B.n79 10.6151
R473 B.n122 B.n79 10.6151
R474 B.n123 B.n122 10.6151
R475 B.n124 B.n77 10.6151
R476 B.n128 B.n77 10.6151
R477 B.n129 B.n128 10.6151
R478 B.n130 B.n129 10.6151
R479 B.n130 B.n75 10.6151
R480 B.n134 B.n75 10.6151
R481 B.n135 B.n134 10.6151
R482 B.n136 B.n135 10.6151
R483 B.n136 B.n73 10.6151
R484 B.n140 B.n73 10.6151
R485 B.n143 B.n142 10.6151
R486 B.n143 B.n69 10.6151
R487 B.n147 B.n69 10.6151
R488 B.n148 B.n147 10.6151
R489 B.n149 B.n148 10.6151
R490 B.n149 B.n67 10.6151
R491 B.n153 B.n67 10.6151
R492 B.n154 B.n153 10.6151
R493 B.n158 B.n154 10.6151
R494 B.n162 B.n65 10.6151
R495 B.n163 B.n162 10.6151
R496 B.n164 B.n163 10.6151
R497 B.n164 B.n63 10.6151
R498 B.n168 B.n63 10.6151
R499 B.n169 B.n168 10.6151
R500 B.n170 B.n169 10.6151
R501 B.n170 B.n61 10.6151
R502 B.n174 B.n61 10.6151
R503 B.n175 B.n174 10.6151
R504 B.n284 B.n283 9.36635
R505 B.n266 B.n30 9.36635
R506 B.n141 B.n140 9.36635
R507 B.n157 B.n65 9.36635
R508 B.n337 B.n0 8.11757
R509 B.n337 B.n1 8.11757
R510 B.n283 B.n282 1.24928
R511 B.n30 B.n26 1.24928
R512 B.n142 B.n141 1.24928
R513 B.n158 B.n157 1.24928
R514 VN VN.t0 101.931
R515 VN VN.t1 65.6059
R516 VTAIL.n3 VTAIL.t2 252.702
R517 VTAIL.n0 VTAIL.t0 252.702
R518 VTAIL.n2 VTAIL.t1 252.702
R519 VTAIL.n1 VTAIL.t3 252.702
R520 VTAIL.n1 VTAIL.n0 18.6858
R521 VTAIL.n3 VTAIL.n2 16.2462
R522 VTAIL.n2 VTAIL.n1 1.69016
R523 VTAIL VTAIL.n0 1.13843
R524 VTAIL VTAIL.n3 0.552224
R525 VDD2.n0 VDD2.t0 299.361
R526 VDD2.n0 VDD2.t1 269.382
R527 VDD2 VDD2.n0 0.668603
R528 VP.n0 VP.t1 101.835
R529 VP.n0 VP.t0 65.2696
R530 VP VP.n0 0.336784
R531 VDD1 VDD1.t1 300.495
R532 VDD1 VDD1.t0 270.05
C0 B w_n2102_n1302# 5.83557f
C1 VDD1 VN 0.15487f
C2 w_n2102_n1302# VP 2.92848f
C3 VTAIL B 1.20676f
C4 VDD2 B 0.905731f
C5 VDD2 VP 0.335664f
C6 VTAIL VP 0.925625f
C7 VN w_n2102_n1302# 2.66663f
C8 VDD1 w_n2102_n1302# 1.04368f
C9 VTAIL VN 0.911492f
C10 VDD2 VN 0.604384f
C11 VDD1 VTAIL 2.30319f
C12 VDD2 VDD1 0.661364f
C13 B VP 1.30583f
C14 VTAIL w_n2102_n1302# 1.23864f
C15 VDD2 w_n2102_n1302# 1.06754f
C16 VDD2 VTAIL 2.35552f
C17 VN B 0.867275f
C18 VDD1 B 0.87613f
C19 VN VP 3.50171f
C20 VDD1 VP 0.783526f
C21 VDD2 VSUBS 0.535909f
C22 VDD1 VSUBS 2.618156f
C23 VTAIL VSUBS 0.345479f
C24 VN VSUBS 5.4133f
C25 VP VSUBS 1.171986f
C26 B VSUBS 2.808639f
C27 w_n2102_n1302# VSUBS 35.036102f
C28 VDD1.t0 VSUBS 0.137362f
C29 VDD1.t1 VSUBS 0.222831f
C30 VP.t1 VSUBS 1.77932f
C31 VP.t0 VSUBS 0.998627f
C32 VP.n0 VSUBS 3.49444f
C33 VDD2.t0 VSUBS 0.230394f
C34 VDD2.t1 VSUBS 0.146768f
C35 VDD2.n0 VSUBS 1.91115f
C36 VTAIL.t0 VSUBS 0.163322f
C37 VTAIL.n0 VSUBS 1.05958f
C38 VTAIL.t3 VSUBS 0.163323f
C39 VTAIL.n1 VSUBS 1.09915f
C40 VTAIL.t1 VSUBS 0.163323f
C41 VTAIL.n2 VSUBS 0.924208f
C42 VTAIL.t2 VSUBS 0.163322f
C43 VTAIL.n3 VSUBS 0.842612f
C44 VN.t1 VSUBS 0.957654f
C45 VN.t0 VSUBS 1.71179f
C46 B.n0 VSUBS 0.008632f
C47 B.n1 VSUBS 0.008632f
C48 B.n2 VSUBS 0.012766f
C49 B.n3 VSUBS 0.009783f
C50 B.n4 VSUBS 0.009783f
C51 B.n5 VSUBS 0.009783f
C52 B.n6 VSUBS 0.009783f
C53 B.n7 VSUBS 0.009783f
C54 B.n8 VSUBS 0.009783f
C55 B.n9 VSUBS 0.009783f
C56 B.n10 VSUBS 0.009783f
C57 B.n11 VSUBS 0.009783f
C58 B.n12 VSUBS 0.009783f
C59 B.n13 VSUBS 0.009783f
C60 B.n14 VSUBS 0.024884f
C61 B.n15 VSUBS 0.009783f
C62 B.n16 VSUBS 0.009783f
C63 B.n17 VSUBS 0.009783f
C64 B.n18 VSUBS 0.009783f
C65 B.n19 VSUBS 0.009783f
C66 B.t4 VSUBS 0.048104f
C67 B.t5 VSUBS 0.059295f
C68 B.t3 VSUBS 0.28901f
C69 B.n20 VSUBS 0.095474f
C70 B.n21 VSUBS 0.076226f
C71 B.n22 VSUBS 0.009783f
C72 B.n23 VSUBS 0.009783f
C73 B.n24 VSUBS 0.009783f
C74 B.n25 VSUBS 0.009783f
C75 B.n26 VSUBS 0.005467f
C76 B.n27 VSUBS 0.009783f
C77 B.t7 VSUBS 0.048104f
C78 B.t8 VSUBS 0.059295f
C79 B.t6 VSUBS 0.28901f
C80 B.n28 VSUBS 0.095474f
C81 B.n29 VSUBS 0.076226f
C82 B.n30 VSUBS 0.022666f
C83 B.n31 VSUBS 0.009783f
C84 B.n32 VSUBS 0.009783f
C85 B.n33 VSUBS 0.009783f
C86 B.n34 VSUBS 0.009783f
C87 B.n35 VSUBS 0.023455f
C88 B.n36 VSUBS 0.009783f
C89 B.n37 VSUBS 0.009783f
C90 B.n38 VSUBS 0.009783f
C91 B.n39 VSUBS 0.009783f
C92 B.n40 VSUBS 0.009783f
C93 B.n41 VSUBS 0.009783f
C94 B.n42 VSUBS 0.009783f
C95 B.n43 VSUBS 0.009783f
C96 B.n44 VSUBS 0.009783f
C97 B.n45 VSUBS 0.009783f
C98 B.n46 VSUBS 0.009783f
C99 B.n47 VSUBS 0.009783f
C100 B.n48 VSUBS 0.009783f
C101 B.n49 VSUBS 0.009783f
C102 B.n50 VSUBS 0.009783f
C103 B.n51 VSUBS 0.009783f
C104 B.n52 VSUBS 0.009783f
C105 B.n53 VSUBS 0.009783f
C106 B.n54 VSUBS 0.009783f
C107 B.n55 VSUBS 0.009783f
C108 B.n56 VSUBS 0.009783f
C109 B.n57 VSUBS 0.009783f
C110 B.n58 VSUBS 0.009783f
C111 B.n59 VSUBS 0.009783f
C112 B.n60 VSUBS 0.024884f
C113 B.n61 VSUBS 0.009783f
C114 B.n62 VSUBS 0.009783f
C115 B.n63 VSUBS 0.009783f
C116 B.n64 VSUBS 0.009783f
C117 B.n65 VSUBS 0.009207f
C118 B.n66 VSUBS 0.009783f
C119 B.n67 VSUBS 0.009783f
C120 B.n68 VSUBS 0.009783f
C121 B.n69 VSUBS 0.009783f
C122 B.n70 VSUBS 0.009783f
C123 B.t2 VSUBS 0.048104f
C124 B.t1 VSUBS 0.059295f
C125 B.t0 VSUBS 0.28901f
C126 B.n71 VSUBS 0.095474f
C127 B.n72 VSUBS 0.076226f
C128 B.n73 VSUBS 0.009783f
C129 B.n74 VSUBS 0.009783f
C130 B.n75 VSUBS 0.009783f
C131 B.n76 VSUBS 0.009783f
C132 B.n77 VSUBS 0.009783f
C133 B.n78 VSUBS 0.023455f
C134 B.n79 VSUBS 0.009783f
C135 B.n80 VSUBS 0.009783f
C136 B.n81 VSUBS 0.009783f
C137 B.n82 VSUBS 0.009783f
C138 B.n83 VSUBS 0.009783f
C139 B.n84 VSUBS 0.009783f
C140 B.n85 VSUBS 0.009783f
C141 B.n86 VSUBS 0.009783f
C142 B.n87 VSUBS 0.009783f
C143 B.n88 VSUBS 0.009783f
C144 B.n89 VSUBS 0.009783f
C145 B.n90 VSUBS 0.009783f
C146 B.n91 VSUBS 0.009783f
C147 B.n92 VSUBS 0.009783f
C148 B.n93 VSUBS 0.009783f
C149 B.n94 VSUBS 0.009783f
C150 B.n95 VSUBS 0.009783f
C151 B.n96 VSUBS 0.009783f
C152 B.n97 VSUBS 0.009783f
C153 B.n98 VSUBS 0.009783f
C154 B.n99 VSUBS 0.009783f
C155 B.n100 VSUBS 0.009783f
C156 B.n101 VSUBS 0.009783f
C157 B.n102 VSUBS 0.009783f
C158 B.n103 VSUBS 0.009783f
C159 B.n104 VSUBS 0.009783f
C160 B.n105 VSUBS 0.009783f
C161 B.n106 VSUBS 0.009783f
C162 B.n107 VSUBS 0.009783f
C163 B.n108 VSUBS 0.009783f
C164 B.n109 VSUBS 0.009783f
C165 B.n110 VSUBS 0.009783f
C166 B.n111 VSUBS 0.009783f
C167 B.n112 VSUBS 0.009783f
C168 B.n113 VSUBS 0.009783f
C169 B.n114 VSUBS 0.009783f
C170 B.n115 VSUBS 0.009783f
C171 B.n116 VSUBS 0.009783f
C172 B.n117 VSUBS 0.009783f
C173 B.n118 VSUBS 0.009783f
C174 B.n119 VSUBS 0.009783f
C175 B.n120 VSUBS 0.009783f
C176 B.n121 VSUBS 0.009783f
C177 B.n122 VSUBS 0.009783f
C178 B.n123 VSUBS 0.023455f
C179 B.n124 VSUBS 0.024884f
C180 B.n125 VSUBS 0.024884f
C181 B.n126 VSUBS 0.009783f
C182 B.n127 VSUBS 0.009783f
C183 B.n128 VSUBS 0.009783f
C184 B.n129 VSUBS 0.009783f
C185 B.n130 VSUBS 0.009783f
C186 B.n131 VSUBS 0.009783f
C187 B.n132 VSUBS 0.009783f
C188 B.n133 VSUBS 0.009783f
C189 B.n134 VSUBS 0.009783f
C190 B.n135 VSUBS 0.009783f
C191 B.n136 VSUBS 0.009783f
C192 B.n137 VSUBS 0.009783f
C193 B.n138 VSUBS 0.009783f
C194 B.n139 VSUBS 0.009783f
C195 B.n140 VSUBS 0.009207f
C196 B.n141 VSUBS 0.022666f
C197 B.n142 VSUBS 0.005467f
C198 B.n143 VSUBS 0.009783f
C199 B.n144 VSUBS 0.009783f
C200 B.n145 VSUBS 0.009783f
C201 B.n146 VSUBS 0.009783f
C202 B.n147 VSUBS 0.009783f
C203 B.n148 VSUBS 0.009783f
C204 B.n149 VSUBS 0.009783f
C205 B.n150 VSUBS 0.009783f
C206 B.n151 VSUBS 0.009783f
C207 B.n152 VSUBS 0.009783f
C208 B.n153 VSUBS 0.009783f
C209 B.n154 VSUBS 0.009783f
C210 B.t11 VSUBS 0.048104f
C211 B.t10 VSUBS 0.059295f
C212 B.t9 VSUBS 0.28901f
C213 B.n155 VSUBS 0.095474f
C214 B.n156 VSUBS 0.076226f
C215 B.n157 VSUBS 0.022666f
C216 B.n158 VSUBS 0.005467f
C217 B.n159 VSUBS 0.009783f
C218 B.n160 VSUBS 0.009783f
C219 B.n161 VSUBS 0.009783f
C220 B.n162 VSUBS 0.009783f
C221 B.n163 VSUBS 0.009783f
C222 B.n164 VSUBS 0.009783f
C223 B.n165 VSUBS 0.009783f
C224 B.n166 VSUBS 0.009783f
C225 B.n167 VSUBS 0.009783f
C226 B.n168 VSUBS 0.009783f
C227 B.n169 VSUBS 0.009783f
C228 B.n170 VSUBS 0.009783f
C229 B.n171 VSUBS 0.009783f
C230 B.n172 VSUBS 0.009783f
C231 B.n173 VSUBS 0.009783f
C232 B.n174 VSUBS 0.009783f
C233 B.n175 VSUBS 0.023818f
C234 B.n176 VSUBS 0.02452f
C235 B.n177 VSUBS 0.023455f
C236 B.n178 VSUBS 0.009783f
C237 B.n179 VSUBS 0.009783f
C238 B.n180 VSUBS 0.009783f
C239 B.n181 VSUBS 0.009783f
C240 B.n182 VSUBS 0.009783f
C241 B.n183 VSUBS 0.009783f
C242 B.n184 VSUBS 0.009783f
C243 B.n185 VSUBS 0.009783f
C244 B.n186 VSUBS 0.009783f
C245 B.n187 VSUBS 0.009783f
C246 B.n188 VSUBS 0.009783f
C247 B.n189 VSUBS 0.009783f
C248 B.n190 VSUBS 0.009783f
C249 B.n191 VSUBS 0.009783f
C250 B.n192 VSUBS 0.009783f
C251 B.n193 VSUBS 0.009783f
C252 B.n194 VSUBS 0.009783f
C253 B.n195 VSUBS 0.009783f
C254 B.n196 VSUBS 0.009783f
C255 B.n197 VSUBS 0.009783f
C256 B.n198 VSUBS 0.009783f
C257 B.n199 VSUBS 0.009783f
C258 B.n200 VSUBS 0.009783f
C259 B.n201 VSUBS 0.009783f
C260 B.n202 VSUBS 0.009783f
C261 B.n203 VSUBS 0.009783f
C262 B.n204 VSUBS 0.009783f
C263 B.n205 VSUBS 0.009783f
C264 B.n206 VSUBS 0.009783f
C265 B.n207 VSUBS 0.009783f
C266 B.n208 VSUBS 0.009783f
C267 B.n209 VSUBS 0.009783f
C268 B.n210 VSUBS 0.009783f
C269 B.n211 VSUBS 0.009783f
C270 B.n212 VSUBS 0.009783f
C271 B.n213 VSUBS 0.009783f
C272 B.n214 VSUBS 0.009783f
C273 B.n215 VSUBS 0.009783f
C274 B.n216 VSUBS 0.009783f
C275 B.n217 VSUBS 0.009783f
C276 B.n218 VSUBS 0.009783f
C277 B.n219 VSUBS 0.009783f
C278 B.n220 VSUBS 0.009783f
C279 B.n221 VSUBS 0.009783f
C280 B.n222 VSUBS 0.009783f
C281 B.n223 VSUBS 0.009783f
C282 B.n224 VSUBS 0.009783f
C283 B.n225 VSUBS 0.009783f
C284 B.n226 VSUBS 0.009783f
C285 B.n227 VSUBS 0.009783f
C286 B.n228 VSUBS 0.009783f
C287 B.n229 VSUBS 0.009783f
C288 B.n230 VSUBS 0.009783f
C289 B.n231 VSUBS 0.009783f
C290 B.n232 VSUBS 0.009783f
C291 B.n233 VSUBS 0.009783f
C292 B.n234 VSUBS 0.009783f
C293 B.n235 VSUBS 0.009783f
C294 B.n236 VSUBS 0.009783f
C295 B.n237 VSUBS 0.009783f
C296 B.n238 VSUBS 0.009783f
C297 B.n239 VSUBS 0.009783f
C298 B.n240 VSUBS 0.009783f
C299 B.n241 VSUBS 0.009783f
C300 B.n242 VSUBS 0.009783f
C301 B.n243 VSUBS 0.009783f
C302 B.n244 VSUBS 0.009783f
C303 B.n245 VSUBS 0.009783f
C304 B.n246 VSUBS 0.009783f
C305 B.n247 VSUBS 0.009783f
C306 B.n248 VSUBS 0.009783f
C307 B.n249 VSUBS 0.009783f
C308 B.n250 VSUBS 0.023455f
C309 B.n251 VSUBS 0.024884f
C310 B.n252 VSUBS 0.024884f
C311 B.n253 VSUBS 0.009783f
C312 B.n254 VSUBS 0.009783f
C313 B.n255 VSUBS 0.009783f
C314 B.n256 VSUBS 0.009783f
C315 B.n257 VSUBS 0.009783f
C316 B.n258 VSUBS 0.009783f
C317 B.n259 VSUBS 0.009783f
C318 B.n260 VSUBS 0.009783f
C319 B.n261 VSUBS 0.009783f
C320 B.n262 VSUBS 0.009783f
C321 B.n263 VSUBS 0.009783f
C322 B.n264 VSUBS 0.009783f
C323 B.n265 VSUBS 0.009783f
C324 B.n266 VSUBS 0.009207f
C325 B.n267 VSUBS 0.009783f
C326 B.n268 VSUBS 0.009783f
C327 B.n269 VSUBS 0.009783f
C328 B.n270 VSUBS 0.009783f
C329 B.n271 VSUBS 0.009783f
C330 B.n272 VSUBS 0.009783f
C331 B.n273 VSUBS 0.009783f
C332 B.n274 VSUBS 0.009783f
C333 B.n275 VSUBS 0.009783f
C334 B.n276 VSUBS 0.009783f
C335 B.n277 VSUBS 0.009783f
C336 B.n278 VSUBS 0.009783f
C337 B.n279 VSUBS 0.009783f
C338 B.n280 VSUBS 0.009783f
C339 B.n281 VSUBS 0.009783f
C340 B.n282 VSUBS 0.005467f
C341 B.n283 VSUBS 0.022666f
C342 B.n284 VSUBS 0.009207f
C343 B.n285 VSUBS 0.009783f
C344 B.n286 VSUBS 0.009783f
C345 B.n287 VSUBS 0.009783f
C346 B.n288 VSUBS 0.009783f
C347 B.n289 VSUBS 0.009783f
C348 B.n290 VSUBS 0.009783f
C349 B.n291 VSUBS 0.009783f
C350 B.n292 VSUBS 0.009783f
C351 B.n293 VSUBS 0.009783f
C352 B.n294 VSUBS 0.009783f
C353 B.n295 VSUBS 0.009783f
C354 B.n296 VSUBS 0.009783f
C355 B.n297 VSUBS 0.009783f
C356 B.n298 VSUBS 0.009783f
C357 B.n299 VSUBS 0.024884f
C358 B.n300 VSUBS 0.023455f
C359 B.n301 VSUBS 0.023455f
C360 B.n302 VSUBS 0.009783f
C361 B.n303 VSUBS 0.009783f
C362 B.n304 VSUBS 0.009783f
C363 B.n305 VSUBS 0.009783f
C364 B.n306 VSUBS 0.009783f
C365 B.n307 VSUBS 0.009783f
C366 B.n308 VSUBS 0.009783f
C367 B.n309 VSUBS 0.009783f
C368 B.n310 VSUBS 0.009783f
C369 B.n311 VSUBS 0.009783f
C370 B.n312 VSUBS 0.009783f
C371 B.n313 VSUBS 0.009783f
C372 B.n314 VSUBS 0.009783f
C373 B.n315 VSUBS 0.009783f
C374 B.n316 VSUBS 0.009783f
C375 B.n317 VSUBS 0.009783f
C376 B.n318 VSUBS 0.009783f
C377 B.n319 VSUBS 0.009783f
C378 B.n320 VSUBS 0.009783f
C379 B.n321 VSUBS 0.009783f
C380 B.n322 VSUBS 0.009783f
C381 B.n323 VSUBS 0.009783f
C382 B.n324 VSUBS 0.009783f
C383 B.n325 VSUBS 0.009783f
C384 B.n326 VSUBS 0.009783f
C385 B.n327 VSUBS 0.009783f
C386 B.n328 VSUBS 0.009783f
C387 B.n329 VSUBS 0.009783f
C388 B.n330 VSUBS 0.009783f
C389 B.n331 VSUBS 0.009783f
C390 B.n332 VSUBS 0.009783f
C391 B.n333 VSUBS 0.009783f
C392 B.n334 VSUBS 0.009783f
C393 B.n335 VSUBS 0.012766f
C394 B.n336 VSUBS 0.013599f
C395 B.n337 VSUBS 0.027043f
.ends

