* NGSPICE file created from diff_pair_sample_1370.ext - technology: sky130A

.subckt diff_pair_sample_1370 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2278_n2956# sky130_fd_pr__pfet_01v8 ad=3.8766 pd=20.66 as=0 ps=0 w=9.94 l=0.76
X1 VTAIL.t19 VN.t0 VDD2.t4 w_n2278_n2956# sky130_fd_pr__pfet_01v8 ad=1.6401 pd=10.27 as=1.6401 ps=10.27 w=9.94 l=0.76
X2 VDD1.t9 VP.t0 VTAIL.t8 w_n2278_n2956# sky130_fd_pr__pfet_01v8 ad=3.8766 pd=20.66 as=1.6401 ps=10.27 w=9.94 l=0.76
X3 VDD2.t9 VN.t1 VTAIL.t18 w_n2278_n2956# sky130_fd_pr__pfet_01v8 ad=1.6401 pd=10.27 as=3.8766 ps=20.66 w=9.94 l=0.76
X4 VTAIL.t17 VN.t2 VDD2.t8 w_n2278_n2956# sky130_fd_pr__pfet_01v8 ad=1.6401 pd=10.27 as=1.6401 ps=10.27 w=9.94 l=0.76
X5 VTAIL.t16 VN.t3 VDD2.t6 w_n2278_n2956# sky130_fd_pr__pfet_01v8 ad=1.6401 pd=10.27 as=1.6401 ps=10.27 w=9.94 l=0.76
X6 VDD2.t2 VN.t4 VTAIL.t15 w_n2278_n2956# sky130_fd_pr__pfet_01v8 ad=1.6401 pd=10.27 as=1.6401 ps=10.27 w=9.94 l=0.76
X7 VDD2.t5 VN.t5 VTAIL.t14 w_n2278_n2956# sky130_fd_pr__pfet_01v8 ad=1.6401 pd=10.27 as=3.8766 ps=20.66 w=9.94 l=0.76
X8 B.t8 B.t6 B.t7 w_n2278_n2956# sky130_fd_pr__pfet_01v8 ad=3.8766 pd=20.66 as=0 ps=0 w=9.94 l=0.76
X9 VDD1.t8 VP.t1 VTAIL.t9 w_n2278_n2956# sky130_fd_pr__pfet_01v8 ad=1.6401 pd=10.27 as=3.8766 ps=20.66 w=9.94 l=0.76
X10 VDD1.t7 VP.t2 VTAIL.t0 w_n2278_n2956# sky130_fd_pr__pfet_01v8 ad=1.6401 pd=10.27 as=1.6401 ps=10.27 w=9.94 l=0.76
X11 VTAIL.t6 VP.t3 VDD1.t6 w_n2278_n2956# sky130_fd_pr__pfet_01v8 ad=1.6401 pd=10.27 as=1.6401 ps=10.27 w=9.94 l=0.76
X12 B.t5 B.t3 B.t4 w_n2278_n2956# sky130_fd_pr__pfet_01v8 ad=3.8766 pd=20.66 as=0 ps=0 w=9.94 l=0.76
X13 VDD2.t3 VN.t6 VTAIL.t13 w_n2278_n2956# sky130_fd_pr__pfet_01v8 ad=1.6401 pd=10.27 as=1.6401 ps=10.27 w=9.94 l=0.76
X14 VDD1.t5 VP.t4 VTAIL.t2 w_n2278_n2956# sky130_fd_pr__pfet_01v8 ad=1.6401 pd=10.27 as=3.8766 ps=20.66 w=9.94 l=0.76
X15 VTAIL.t3 VP.t5 VDD1.t4 w_n2278_n2956# sky130_fd_pr__pfet_01v8 ad=1.6401 pd=10.27 as=1.6401 ps=10.27 w=9.94 l=0.76
X16 VDD1.t3 VP.t6 VTAIL.t5 w_n2278_n2956# sky130_fd_pr__pfet_01v8 ad=1.6401 pd=10.27 as=1.6401 ps=10.27 w=9.94 l=0.76
X17 VDD1.t2 VP.t7 VTAIL.t1 w_n2278_n2956# sky130_fd_pr__pfet_01v8 ad=3.8766 pd=20.66 as=1.6401 ps=10.27 w=9.94 l=0.76
X18 B.t2 B.t0 B.t1 w_n2278_n2956# sky130_fd_pr__pfet_01v8 ad=3.8766 pd=20.66 as=0 ps=0 w=9.94 l=0.76
X19 VTAIL.t7 VP.t8 VDD1.t1 w_n2278_n2956# sky130_fd_pr__pfet_01v8 ad=1.6401 pd=10.27 as=1.6401 ps=10.27 w=9.94 l=0.76
X20 VDD2.t1 VN.t7 VTAIL.t12 w_n2278_n2956# sky130_fd_pr__pfet_01v8 ad=3.8766 pd=20.66 as=1.6401 ps=10.27 w=9.94 l=0.76
X21 VDD2.t0 VN.t8 VTAIL.t11 w_n2278_n2956# sky130_fd_pr__pfet_01v8 ad=3.8766 pd=20.66 as=1.6401 ps=10.27 w=9.94 l=0.76
X22 VTAIL.t4 VP.t9 VDD1.t0 w_n2278_n2956# sky130_fd_pr__pfet_01v8 ad=1.6401 pd=10.27 as=1.6401 ps=10.27 w=9.94 l=0.76
X23 VTAIL.t10 VN.t9 VDD2.t7 w_n2278_n2956# sky130_fd_pr__pfet_01v8 ad=1.6401 pd=10.27 as=1.6401 ps=10.27 w=9.94 l=0.76
R0 B.n308 B.n307 585
R1 B.n306 B.n89 585
R2 B.n305 B.n304 585
R3 B.n303 B.n90 585
R4 B.n302 B.n301 585
R5 B.n300 B.n91 585
R6 B.n299 B.n298 585
R7 B.n297 B.n92 585
R8 B.n296 B.n295 585
R9 B.n294 B.n93 585
R10 B.n293 B.n292 585
R11 B.n291 B.n94 585
R12 B.n290 B.n289 585
R13 B.n288 B.n95 585
R14 B.n287 B.n286 585
R15 B.n285 B.n96 585
R16 B.n284 B.n283 585
R17 B.n282 B.n97 585
R18 B.n281 B.n280 585
R19 B.n279 B.n98 585
R20 B.n278 B.n277 585
R21 B.n276 B.n99 585
R22 B.n275 B.n274 585
R23 B.n273 B.n100 585
R24 B.n272 B.n271 585
R25 B.n270 B.n101 585
R26 B.n269 B.n268 585
R27 B.n267 B.n102 585
R28 B.n266 B.n265 585
R29 B.n264 B.n103 585
R30 B.n263 B.n262 585
R31 B.n261 B.n104 585
R32 B.n260 B.n259 585
R33 B.n258 B.n105 585
R34 B.n257 B.n256 585
R35 B.n255 B.n106 585
R36 B.n254 B.n253 585
R37 B.n249 B.n107 585
R38 B.n248 B.n247 585
R39 B.n246 B.n108 585
R40 B.n245 B.n244 585
R41 B.n243 B.n109 585
R42 B.n242 B.n241 585
R43 B.n240 B.n110 585
R44 B.n239 B.n238 585
R45 B.n236 B.n111 585
R46 B.n235 B.n234 585
R47 B.n233 B.n114 585
R48 B.n232 B.n231 585
R49 B.n230 B.n115 585
R50 B.n229 B.n228 585
R51 B.n227 B.n116 585
R52 B.n226 B.n225 585
R53 B.n224 B.n117 585
R54 B.n223 B.n222 585
R55 B.n221 B.n118 585
R56 B.n220 B.n219 585
R57 B.n218 B.n119 585
R58 B.n217 B.n216 585
R59 B.n215 B.n120 585
R60 B.n214 B.n213 585
R61 B.n212 B.n121 585
R62 B.n211 B.n210 585
R63 B.n209 B.n122 585
R64 B.n208 B.n207 585
R65 B.n206 B.n123 585
R66 B.n205 B.n204 585
R67 B.n203 B.n124 585
R68 B.n202 B.n201 585
R69 B.n200 B.n125 585
R70 B.n199 B.n198 585
R71 B.n197 B.n126 585
R72 B.n196 B.n195 585
R73 B.n194 B.n127 585
R74 B.n193 B.n192 585
R75 B.n191 B.n128 585
R76 B.n190 B.n189 585
R77 B.n188 B.n129 585
R78 B.n187 B.n186 585
R79 B.n185 B.n130 585
R80 B.n184 B.n183 585
R81 B.n309 B.n88 585
R82 B.n311 B.n310 585
R83 B.n312 B.n87 585
R84 B.n314 B.n313 585
R85 B.n315 B.n86 585
R86 B.n317 B.n316 585
R87 B.n318 B.n85 585
R88 B.n320 B.n319 585
R89 B.n321 B.n84 585
R90 B.n323 B.n322 585
R91 B.n324 B.n83 585
R92 B.n326 B.n325 585
R93 B.n327 B.n82 585
R94 B.n329 B.n328 585
R95 B.n330 B.n81 585
R96 B.n332 B.n331 585
R97 B.n333 B.n80 585
R98 B.n335 B.n334 585
R99 B.n336 B.n79 585
R100 B.n338 B.n337 585
R101 B.n339 B.n78 585
R102 B.n341 B.n340 585
R103 B.n342 B.n77 585
R104 B.n344 B.n343 585
R105 B.n345 B.n76 585
R106 B.n347 B.n346 585
R107 B.n348 B.n75 585
R108 B.n350 B.n349 585
R109 B.n351 B.n74 585
R110 B.n353 B.n352 585
R111 B.n354 B.n73 585
R112 B.n356 B.n355 585
R113 B.n357 B.n72 585
R114 B.n359 B.n358 585
R115 B.n360 B.n71 585
R116 B.n362 B.n361 585
R117 B.n363 B.n70 585
R118 B.n365 B.n364 585
R119 B.n366 B.n69 585
R120 B.n368 B.n367 585
R121 B.n369 B.n68 585
R122 B.n371 B.n370 585
R123 B.n372 B.n67 585
R124 B.n374 B.n373 585
R125 B.n375 B.n66 585
R126 B.n377 B.n376 585
R127 B.n378 B.n65 585
R128 B.n380 B.n379 585
R129 B.n381 B.n64 585
R130 B.n383 B.n382 585
R131 B.n384 B.n63 585
R132 B.n386 B.n385 585
R133 B.n387 B.n62 585
R134 B.n389 B.n388 585
R135 B.n390 B.n61 585
R136 B.n392 B.n391 585
R137 B.n515 B.n514 585
R138 B.n513 B.n16 585
R139 B.n512 B.n511 585
R140 B.n510 B.n17 585
R141 B.n509 B.n508 585
R142 B.n507 B.n18 585
R143 B.n506 B.n505 585
R144 B.n504 B.n19 585
R145 B.n503 B.n502 585
R146 B.n501 B.n20 585
R147 B.n500 B.n499 585
R148 B.n498 B.n21 585
R149 B.n497 B.n496 585
R150 B.n495 B.n22 585
R151 B.n494 B.n493 585
R152 B.n492 B.n23 585
R153 B.n491 B.n490 585
R154 B.n489 B.n24 585
R155 B.n488 B.n487 585
R156 B.n486 B.n25 585
R157 B.n485 B.n484 585
R158 B.n483 B.n26 585
R159 B.n482 B.n481 585
R160 B.n480 B.n27 585
R161 B.n479 B.n478 585
R162 B.n477 B.n28 585
R163 B.n476 B.n475 585
R164 B.n474 B.n29 585
R165 B.n473 B.n472 585
R166 B.n471 B.n30 585
R167 B.n470 B.n469 585
R168 B.n468 B.n31 585
R169 B.n467 B.n466 585
R170 B.n465 B.n32 585
R171 B.n464 B.n463 585
R172 B.n462 B.n33 585
R173 B.n460 B.n459 585
R174 B.n458 B.n36 585
R175 B.n457 B.n456 585
R176 B.n455 B.n37 585
R177 B.n454 B.n453 585
R178 B.n452 B.n38 585
R179 B.n451 B.n450 585
R180 B.n449 B.n39 585
R181 B.n448 B.n447 585
R182 B.n446 B.n445 585
R183 B.n444 B.n43 585
R184 B.n443 B.n442 585
R185 B.n441 B.n44 585
R186 B.n440 B.n439 585
R187 B.n438 B.n45 585
R188 B.n437 B.n436 585
R189 B.n435 B.n46 585
R190 B.n434 B.n433 585
R191 B.n432 B.n47 585
R192 B.n431 B.n430 585
R193 B.n429 B.n48 585
R194 B.n428 B.n427 585
R195 B.n426 B.n49 585
R196 B.n425 B.n424 585
R197 B.n423 B.n50 585
R198 B.n422 B.n421 585
R199 B.n420 B.n51 585
R200 B.n419 B.n418 585
R201 B.n417 B.n52 585
R202 B.n416 B.n415 585
R203 B.n414 B.n53 585
R204 B.n413 B.n412 585
R205 B.n411 B.n54 585
R206 B.n410 B.n409 585
R207 B.n408 B.n55 585
R208 B.n407 B.n406 585
R209 B.n405 B.n56 585
R210 B.n404 B.n403 585
R211 B.n402 B.n57 585
R212 B.n401 B.n400 585
R213 B.n399 B.n58 585
R214 B.n398 B.n397 585
R215 B.n396 B.n59 585
R216 B.n395 B.n394 585
R217 B.n393 B.n60 585
R218 B.n516 B.n15 585
R219 B.n518 B.n517 585
R220 B.n519 B.n14 585
R221 B.n521 B.n520 585
R222 B.n522 B.n13 585
R223 B.n524 B.n523 585
R224 B.n525 B.n12 585
R225 B.n527 B.n526 585
R226 B.n528 B.n11 585
R227 B.n530 B.n529 585
R228 B.n531 B.n10 585
R229 B.n533 B.n532 585
R230 B.n534 B.n9 585
R231 B.n536 B.n535 585
R232 B.n537 B.n8 585
R233 B.n539 B.n538 585
R234 B.n540 B.n7 585
R235 B.n542 B.n541 585
R236 B.n543 B.n6 585
R237 B.n545 B.n544 585
R238 B.n546 B.n5 585
R239 B.n548 B.n547 585
R240 B.n549 B.n4 585
R241 B.n551 B.n550 585
R242 B.n552 B.n3 585
R243 B.n554 B.n553 585
R244 B.n555 B.n0 585
R245 B.n2 B.n1 585
R246 B.n145 B.n144 585
R247 B.n146 B.n143 585
R248 B.n148 B.n147 585
R249 B.n149 B.n142 585
R250 B.n151 B.n150 585
R251 B.n152 B.n141 585
R252 B.n154 B.n153 585
R253 B.n155 B.n140 585
R254 B.n157 B.n156 585
R255 B.n158 B.n139 585
R256 B.n160 B.n159 585
R257 B.n161 B.n138 585
R258 B.n163 B.n162 585
R259 B.n164 B.n137 585
R260 B.n166 B.n165 585
R261 B.n167 B.n136 585
R262 B.n169 B.n168 585
R263 B.n170 B.n135 585
R264 B.n172 B.n171 585
R265 B.n173 B.n134 585
R266 B.n175 B.n174 585
R267 B.n176 B.n133 585
R268 B.n178 B.n177 585
R269 B.n179 B.n132 585
R270 B.n181 B.n180 585
R271 B.n182 B.n131 585
R272 B.n112 B.t0 517.489
R273 B.n250 B.t6 517.489
R274 B.n40 B.t3 517.489
R275 B.n34 B.t9 517.489
R276 B.n184 B.n131 449.257
R277 B.n309 B.n308 449.257
R278 B.n393 B.n392 449.257
R279 B.n514 B.n15 449.257
R280 B.n250 B.t7 359.553
R281 B.n40 B.t5 359.553
R282 B.n112 B.t1 359.551
R283 B.n34 B.t11 359.551
R284 B.n251 B.t8 338.413
R285 B.n41 B.t4 338.413
R286 B.n113 B.t2 338.413
R287 B.n35 B.t10 338.413
R288 B.n557 B.n556 256.663
R289 B.n556 B.n555 235.042
R290 B.n556 B.n2 235.042
R291 B.n185 B.n184 163.367
R292 B.n186 B.n185 163.367
R293 B.n186 B.n129 163.367
R294 B.n190 B.n129 163.367
R295 B.n191 B.n190 163.367
R296 B.n192 B.n191 163.367
R297 B.n192 B.n127 163.367
R298 B.n196 B.n127 163.367
R299 B.n197 B.n196 163.367
R300 B.n198 B.n197 163.367
R301 B.n198 B.n125 163.367
R302 B.n202 B.n125 163.367
R303 B.n203 B.n202 163.367
R304 B.n204 B.n203 163.367
R305 B.n204 B.n123 163.367
R306 B.n208 B.n123 163.367
R307 B.n209 B.n208 163.367
R308 B.n210 B.n209 163.367
R309 B.n210 B.n121 163.367
R310 B.n214 B.n121 163.367
R311 B.n215 B.n214 163.367
R312 B.n216 B.n215 163.367
R313 B.n216 B.n119 163.367
R314 B.n220 B.n119 163.367
R315 B.n221 B.n220 163.367
R316 B.n222 B.n221 163.367
R317 B.n222 B.n117 163.367
R318 B.n226 B.n117 163.367
R319 B.n227 B.n226 163.367
R320 B.n228 B.n227 163.367
R321 B.n228 B.n115 163.367
R322 B.n232 B.n115 163.367
R323 B.n233 B.n232 163.367
R324 B.n234 B.n233 163.367
R325 B.n234 B.n111 163.367
R326 B.n239 B.n111 163.367
R327 B.n240 B.n239 163.367
R328 B.n241 B.n240 163.367
R329 B.n241 B.n109 163.367
R330 B.n245 B.n109 163.367
R331 B.n246 B.n245 163.367
R332 B.n247 B.n246 163.367
R333 B.n247 B.n107 163.367
R334 B.n254 B.n107 163.367
R335 B.n255 B.n254 163.367
R336 B.n256 B.n255 163.367
R337 B.n256 B.n105 163.367
R338 B.n260 B.n105 163.367
R339 B.n261 B.n260 163.367
R340 B.n262 B.n261 163.367
R341 B.n262 B.n103 163.367
R342 B.n266 B.n103 163.367
R343 B.n267 B.n266 163.367
R344 B.n268 B.n267 163.367
R345 B.n268 B.n101 163.367
R346 B.n272 B.n101 163.367
R347 B.n273 B.n272 163.367
R348 B.n274 B.n273 163.367
R349 B.n274 B.n99 163.367
R350 B.n278 B.n99 163.367
R351 B.n279 B.n278 163.367
R352 B.n280 B.n279 163.367
R353 B.n280 B.n97 163.367
R354 B.n284 B.n97 163.367
R355 B.n285 B.n284 163.367
R356 B.n286 B.n285 163.367
R357 B.n286 B.n95 163.367
R358 B.n290 B.n95 163.367
R359 B.n291 B.n290 163.367
R360 B.n292 B.n291 163.367
R361 B.n292 B.n93 163.367
R362 B.n296 B.n93 163.367
R363 B.n297 B.n296 163.367
R364 B.n298 B.n297 163.367
R365 B.n298 B.n91 163.367
R366 B.n302 B.n91 163.367
R367 B.n303 B.n302 163.367
R368 B.n304 B.n303 163.367
R369 B.n304 B.n89 163.367
R370 B.n308 B.n89 163.367
R371 B.n392 B.n61 163.367
R372 B.n388 B.n61 163.367
R373 B.n388 B.n387 163.367
R374 B.n387 B.n386 163.367
R375 B.n386 B.n63 163.367
R376 B.n382 B.n63 163.367
R377 B.n382 B.n381 163.367
R378 B.n381 B.n380 163.367
R379 B.n380 B.n65 163.367
R380 B.n376 B.n65 163.367
R381 B.n376 B.n375 163.367
R382 B.n375 B.n374 163.367
R383 B.n374 B.n67 163.367
R384 B.n370 B.n67 163.367
R385 B.n370 B.n369 163.367
R386 B.n369 B.n368 163.367
R387 B.n368 B.n69 163.367
R388 B.n364 B.n69 163.367
R389 B.n364 B.n363 163.367
R390 B.n363 B.n362 163.367
R391 B.n362 B.n71 163.367
R392 B.n358 B.n71 163.367
R393 B.n358 B.n357 163.367
R394 B.n357 B.n356 163.367
R395 B.n356 B.n73 163.367
R396 B.n352 B.n73 163.367
R397 B.n352 B.n351 163.367
R398 B.n351 B.n350 163.367
R399 B.n350 B.n75 163.367
R400 B.n346 B.n75 163.367
R401 B.n346 B.n345 163.367
R402 B.n345 B.n344 163.367
R403 B.n344 B.n77 163.367
R404 B.n340 B.n77 163.367
R405 B.n340 B.n339 163.367
R406 B.n339 B.n338 163.367
R407 B.n338 B.n79 163.367
R408 B.n334 B.n79 163.367
R409 B.n334 B.n333 163.367
R410 B.n333 B.n332 163.367
R411 B.n332 B.n81 163.367
R412 B.n328 B.n81 163.367
R413 B.n328 B.n327 163.367
R414 B.n327 B.n326 163.367
R415 B.n326 B.n83 163.367
R416 B.n322 B.n83 163.367
R417 B.n322 B.n321 163.367
R418 B.n321 B.n320 163.367
R419 B.n320 B.n85 163.367
R420 B.n316 B.n85 163.367
R421 B.n316 B.n315 163.367
R422 B.n315 B.n314 163.367
R423 B.n314 B.n87 163.367
R424 B.n310 B.n87 163.367
R425 B.n310 B.n309 163.367
R426 B.n514 B.n513 163.367
R427 B.n513 B.n512 163.367
R428 B.n512 B.n17 163.367
R429 B.n508 B.n17 163.367
R430 B.n508 B.n507 163.367
R431 B.n507 B.n506 163.367
R432 B.n506 B.n19 163.367
R433 B.n502 B.n19 163.367
R434 B.n502 B.n501 163.367
R435 B.n501 B.n500 163.367
R436 B.n500 B.n21 163.367
R437 B.n496 B.n21 163.367
R438 B.n496 B.n495 163.367
R439 B.n495 B.n494 163.367
R440 B.n494 B.n23 163.367
R441 B.n490 B.n23 163.367
R442 B.n490 B.n489 163.367
R443 B.n489 B.n488 163.367
R444 B.n488 B.n25 163.367
R445 B.n484 B.n25 163.367
R446 B.n484 B.n483 163.367
R447 B.n483 B.n482 163.367
R448 B.n482 B.n27 163.367
R449 B.n478 B.n27 163.367
R450 B.n478 B.n477 163.367
R451 B.n477 B.n476 163.367
R452 B.n476 B.n29 163.367
R453 B.n472 B.n29 163.367
R454 B.n472 B.n471 163.367
R455 B.n471 B.n470 163.367
R456 B.n470 B.n31 163.367
R457 B.n466 B.n31 163.367
R458 B.n466 B.n465 163.367
R459 B.n465 B.n464 163.367
R460 B.n464 B.n33 163.367
R461 B.n459 B.n33 163.367
R462 B.n459 B.n458 163.367
R463 B.n458 B.n457 163.367
R464 B.n457 B.n37 163.367
R465 B.n453 B.n37 163.367
R466 B.n453 B.n452 163.367
R467 B.n452 B.n451 163.367
R468 B.n451 B.n39 163.367
R469 B.n447 B.n39 163.367
R470 B.n447 B.n446 163.367
R471 B.n446 B.n43 163.367
R472 B.n442 B.n43 163.367
R473 B.n442 B.n441 163.367
R474 B.n441 B.n440 163.367
R475 B.n440 B.n45 163.367
R476 B.n436 B.n45 163.367
R477 B.n436 B.n435 163.367
R478 B.n435 B.n434 163.367
R479 B.n434 B.n47 163.367
R480 B.n430 B.n47 163.367
R481 B.n430 B.n429 163.367
R482 B.n429 B.n428 163.367
R483 B.n428 B.n49 163.367
R484 B.n424 B.n49 163.367
R485 B.n424 B.n423 163.367
R486 B.n423 B.n422 163.367
R487 B.n422 B.n51 163.367
R488 B.n418 B.n51 163.367
R489 B.n418 B.n417 163.367
R490 B.n417 B.n416 163.367
R491 B.n416 B.n53 163.367
R492 B.n412 B.n53 163.367
R493 B.n412 B.n411 163.367
R494 B.n411 B.n410 163.367
R495 B.n410 B.n55 163.367
R496 B.n406 B.n55 163.367
R497 B.n406 B.n405 163.367
R498 B.n405 B.n404 163.367
R499 B.n404 B.n57 163.367
R500 B.n400 B.n57 163.367
R501 B.n400 B.n399 163.367
R502 B.n399 B.n398 163.367
R503 B.n398 B.n59 163.367
R504 B.n394 B.n59 163.367
R505 B.n394 B.n393 163.367
R506 B.n518 B.n15 163.367
R507 B.n519 B.n518 163.367
R508 B.n520 B.n519 163.367
R509 B.n520 B.n13 163.367
R510 B.n524 B.n13 163.367
R511 B.n525 B.n524 163.367
R512 B.n526 B.n525 163.367
R513 B.n526 B.n11 163.367
R514 B.n530 B.n11 163.367
R515 B.n531 B.n530 163.367
R516 B.n532 B.n531 163.367
R517 B.n532 B.n9 163.367
R518 B.n536 B.n9 163.367
R519 B.n537 B.n536 163.367
R520 B.n538 B.n537 163.367
R521 B.n538 B.n7 163.367
R522 B.n542 B.n7 163.367
R523 B.n543 B.n542 163.367
R524 B.n544 B.n543 163.367
R525 B.n544 B.n5 163.367
R526 B.n548 B.n5 163.367
R527 B.n549 B.n548 163.367
R528 B.n550 B.n549 163.367
R529 B.n550 B.n3 163.367
R530 B.n554 B.n3 163.367
R531 B.n555 B.n554 163.367
R532 B.n144 B.n2 163.367
R533 B.n144 B.n143 163.367
R534 B.n148 B.n143 163.367
R535 B.n149 B.n148 163.367
R536 B.n150 B.n149 163.367
R537 B.n150 B.n141 163.367
R538 B.n154 B.n141 163.367
R539 B.n155 B.n154 163.367
R540 B.n156 B.n155 163.367
R541 B.n156 B.n139 163.367
R542 B.n160 B.n139 163.367
R543 B.n161 B.n160 163.367
R544 B.n162 B.n161 163.367
R545 B.n162 B.n137 163.367
R546 B.n166 B.n137 163.367
R547 B.n167 B.n166 163.367
R548 B.n168 B.n167 163.367
R549 B.n168 B.n135 163.367
R550 B.n172 B.n135 163.367
R551 B.n173 B.n172 163.367
R552 B.n174 B.n173 163.367
R553 B.n174 B.n133 163.367
R554 B.n178 B.n133 163.367
R555 B.n179 B.n178 163.367
R556 B.n180 B.n179 163.367
R557 B.n180 B.n131 163.367
R558 B.n237 B.n113 59.5399
R559 B.n252 B.n251 59.5399
R560 B.n42 B.n41 59.5399
R561 B.n461 B.n35 59.5399
R562 B.n516 B.n515 29.1907
R563 B.n391 B.n60 29.1907
R564 B.n307 B.n88 29.1907
R565 B.n183 B.n182 29.1907
R566 B.n113 B.n112 21.1399
R567 B.n251 B.n250 21.1399
R568 B.n41 B.n40 21.1399
R569 B.n35 B.n34 21.1399
R570 B B.n557 18.0485
R571 B.n517 B.n516 10.6151
R572 B.n517 B.n14 10.6151
R573 B.n521 B.n14 10.6151
R574 B.n522 B.n521 10.6151
R575 B.n523 B.n522 10.6151
R576 B.n523 B.n12 10.6151
R577 B.n527 B.n12 10.6151
R578 B.n528 B.n527 10.6151
R579 B.n529 B.n528 10.6151
R580 B.n529 B.n10 10.6151
R581 B.n533 B.n10 10.6151
R582 B.n534 B.n533 10.6151
R583 B.n535 B.n534 10.6151
R584 B.n535 B.n8 10.6151
R585 B.n539 B.n8 10.6151
R586 B.n540 B.n539 10.6151
R587 B.n541 B.n540 10.6151
R588 B.n541 B.n6 10.6151
R589 B.n545 B.n6 10.6151
R590 B.n546 B.n545 10.6151
R591 B.n547 B.n546 10.6151
R592 B.n547 B.n4 10.6151
R593 B.n551 B.n4 10.6151
R594 B.n552 B.n551 10.6151
R595 B.n553 B.n552 10.6151
R596 B.n553 B.n0 10.6151
R597 B.n515 B.n16 10.6151
R598 B.n511 B.n16 10.6151
R599 B.n511 B.n510 10.6151
R600 B.n510 B.n509 10.6151
R601 B.n509 B.n18 10.6151
R602 B.n505 B.n18 10.6151
R603 B.n505 B.n504 10.6151
R604 B.n504 B.n503 10.6151
R605 B.n503 B.n20 10.6151
R606 B.n499 B.n20 10.6151
R607 B.n499 B.n498 10.6151
R608 B.n498 B.n497 10.6151
R609 B.n497 B.n22 10.6151
R610 B.n493 B.n22 10.6151
R611 B.n493 B.n492 10.6151
R612 B.n492 B.n491 10.6151
R613 B.n491 B.n24 10.6151
R614 B.n487 B.n24 10.6151
R615 B.n487 B.n486 10.6151
R616 B.n486 B.n485 10.6151
R617 B.n485 B.n26 10.6151
R618 B.n481 B.n26 10.6151
R619 B.n481 B.n480 10.6151
R620 B.n480 B.n479 10.6151
R621 B.n479 B.n28 10.6151
R622 B.n475 B.n28 10.6151
R623 B.n475 B.n474 10.6151
R624 B.n474 B.n473 10.6151
R625 B.n473 B.n30 10.6151
R626 B.n469 B.n30 10.6151
R627 B.n469 B.n468 10.6151
R628 B.n468 B.n467 10.6151
R629 B.n467 B.n32 10.6151
R630 B.n463 B.n32 10.6151
R631 B.n463 B.n462 10.6151
R632 B.n460 B.n36 10.6151
R633 B.n456 B.n36 10.6151
R634 B.n456 B.n455 10.6151
R635 B.n455 B.n454 10.6151
R636 B.n454 B.n38 10.6151
R637 B.n450 B.n38 10.6151
R638 B.n450 B.n449 10.6151
R639 B.n449 B.n448 10.6151
R640 B.n445 B.n444 10.6151
R641 B.n444 B.n443 10.6151
R642 B.n443 B.n44 10.6151
R643 B.n439 B.n44 10.6151
R644 B.n439 B.n438 10.6151
R645 B.n438 B.n437 10.6151
R646 B.n437 B.n46 10.6151
R647 B.n433 B.n46 10.6151
R648 B.n433 B.n432 10.6151
R649 B.n432 B.n431 10.6151
R650 B.n431 B.n48 10.6151
R651 B.n427 B.n48 10.6151
R652 B.n427 B.n426 10.6151
R653 B.n426 B.n425 10.6151
R654 B.n425 B.n50 10.6151
R655 B.n421 B.n50 10.6151
R656 B.n421 B.n420 10.6151
R657 B.n420 B.n419 10.6151
R658 B.n419 B.n52 10.6151
R659 B.n415 B.n52 10.6151
R660 B.n415 B.n414 10.6151
R661 B.n414 B.n413 10.6151
R662 B.n413 B.n54 10.6151
R663 B.n409 B.n54 10.6151
R664 B.n409 B.n408 10.6151
R665 B.n408 B.n407 10.6151
R666 B.n407 B.n56 10.6151
R667 B.n403 B.n56 10.6151
R668 B.n403 B.n402 10.6151
R669 B.n402 B.n401 10.6151
R670 B.n401 B.n58 10.6151
R671 B.n397 B.n58 10.6151
R672 B.n397 B.n396 10.6151
R673 B.n396 B.n395 10.6151
R674 B.n395 B.n60 10.6151
R675 B.n391 B.n390 10.6151
R676 B.n390 B.n389 10.6151
R677 B.n389 B.n62 10.6151
R678 B.n385 B.n62 10.6151
R679 B.n385 B.n384 10.6151
R680 B.n384 B.n383 10.6151
R681 B.n383 B.n64 10.6151
R682 B.n379 B.n64 10.6151
R683 B.n379 B.n378 10.6151
R684 B.n378 B.n377 10.6151
R685 B.n377 B.n66 10.6151
R686 B.n373 B.n66 10.6151
R687 B.n373 B.n372 10.6151
R688 B.n372 B.n371 10.6151
R689 B.n371 B.n68 10.6151
R690 B.n367 B.n68 10.6151
R691 B.n367 B.n366 10.6151
R692 B.n366 B.n365 10.6151
R693 B.n365 B.n70 10.6151
R694 B.n361 B.n70 10.6151
R695 B.n361 B.n360 10.6151
R696 B.n360 B.n359 10.6151
R697 B.n359 B.n72 10.6151
R698 B.n355 B.n72 10.6151
R699 B.n355 B.n354 10.6151
R700 B.n354 B.n353 10.6151
R701 B.n353 B.n74 10.6151
R702 B.n349 B.n74 10.6151
R703 B.n349 B.n348 10.6151
R704 B.n348 B.n347 10.6151
R705 B.n347 B.n76 10.6151
R706 B.n343 B.n76 10.6151
R707 B.n343 B.n342 10.6151
R708 B.n342 B.n341 10.6151
R709 B.n341 B.n78 10.6151
R710 B.n337 B.n78 10.6151
R711 B.n337 B.n336 10.6151
R712 B.n336 B.n335 10.6151
R713 B.n335 B.n80 10.6151
R714 B.n331 B.n80 10.6151
R715 B.n331 B.n330 10.6151
R716 B.n330 B.n329 10.6151
R717 B.n329 B.n82 10.6151
R718 B.n325 B.n82 10.6151
R719 B.n325 B.n324 10.6151
R720 B.n324 B.n323 10.6151
R721 B.n323 B.n84 10.6151
R722 B.n319 B.n84 10.6151
R723 B.n319 B.n318 10.6151
R724 B.n318 B.n317 10.6151
R725 B.n317 B.n86 10.6151
R726 B.n313 B.n86 10.6151
R727 B.n313 B.n312 10.6151
R728 B.n312 B.n311 10.6151
R729 B.n311 B.n88 10.6151
R730 B.n145 B.n1 10.6151
R731 B.n146 B.n145 10.6151
R732 B.n147 B.n146 10.6151
R733 B.n147 B.n142 10.6151
R734 B.n151 B.n142 10.6151
R735 B.n152 B.n151 10.6151
R736 B.n153 B.n152 10.6151
R737 B.n153 B.n140 10.6151
R738 B.n157 B.n140 10.6151
R739 B.n158 B.n157 10.6151
R740 B.n159 B.n158 10.6151
R741 B.n159 B.n138 10.6151
R742 B.n163 B.n138 10.6151
R743 B.n164 B.n163 10.6151
R744 B.n165 B.n164 10.6151
R745 B.n165 B.n136 10.6151
R746 B.n169 B.n136 10.6151
R747 B.n170 B.n169 10.6151
R748 B.n171 B.n170 10.6151
R749 B.n171 B.n134 10.6151
R750 B.n175 B.n134 10.6151
R751 B.n176 B.n175 10.6151
R752 B.n177 B.n176 10.6151
R753 B.n177 B.n132 10.6151
R754 B.n181 B.n132 10.6151
R755 B.n182 B.n181 10.6151
R756 B.n183 B.n130 10.6151
R757 B.n187 B.n130 10.6151
R758 B.n188 B.n187 10.6151
R759 B.n189 B.n188 10.6151
R760 B.n189 B.n128 10.6151
R761 B.n193 B.n128 10.6151
R762 B.n194 B.n193 10.6151
R763 B.n195 B.n194 10.6151
R764 B.n195 B.n126 10.6151
R765 B.n199 B.n126 10.6151
R766 B.n200 B.n199 10.6151
R767 B.n201 B.n200 10.6151
R768 B.n201 B.n124 10.6151
R769 B.n205 B.n124 10.6151
R770 B.n206 B.n205 10.6151
R771 B.n207 B.n206 10.6151
R772 B.n207 B.n122 10.6151
R773 B.n211 B.n122 10.6151
R774 B.n212 B.n211 10.6151
R775 B.n213 B.n212 10.6151
R776 B.n213 B.n120 10.6151
R777 B.n217 B.n120 10.6151
R778 B.n218 B.n217 10.6151
R779 B.n219 B.n218 10.6151
R780 B.n219 B.n118 10.6151
R781 B.n223 B.n118 10.6151
R782 B.n224 B.n223 10.6151
R783 B.n225 B.n224 10.6151
R784 B.n225 B.n116 10.6151
R785 B.n229 B.n116 10.6151
R786 B.n230 B.n229 10.6151
R787 B.n231 B.n230 10.6151
R788 B.n231 B.n114 10.6151
R789 B.n235 B.n114 10.6151
R790 B.n236 B.n235 10.6151
R791 B.n238 B.n110 10.6151
R792 B.n242 B.n110 10.6151
R793 B.n243 B.n242 10.6151
R794 B.n244 B.n243 10.6151
R795 B.n244 B.n108 10.6151
R796 B.n248 B.n108 10.6151
R797 B.n249 B.n248 10.6151
R798 B.n253 B.n249 10.6151
R799 B.n257 B.n106 10.6151
R800 B.n258 B.n257 10.6151
R801 B.n259 B.n258 10.6151
R802 B.n259 B.n104 10.6151
R803 B.n263 B.n104 10.6151
R804 B.n264 B.n263 10.6151
R805 B.n265 B.n264 10.6151
R806 B.n265 B.n102 10.6151
R807 B.n269 B.n102 10.6151
R808 B.n270 B.n269 10.6151
R809 B.n271 B.n270 10.6151
R810 B.n271 B.n100 10.6151
R811 B.n275 B.n100 10.6151
R812 B.n276 B.n275 10.6151
R813 B.n277 B.n276 10.6151
R814 B.n277 B.n98 10.6151
R815 B.n281 B.n98 10.6151
R816 B.n282 B.n281 10.6151
R817 B.n283 B.n282 10.6151
R818 B.n283 B.n96 10.6151
R819 B.n287 B.n96 10.6151
R820 B.n288 B.n287 10.6151
R821 B.n289 B.n288 10.6151
R822 B.n289 B.n94 10.6151
R823 B.n293 B.n94 10.6151
R824 B.n294 B.n293 10.6151
R825 B.n295 B.n294 10.6151
R826 B.n295 B.n92 10.6151
R827 B.n299 B.n92 10.6151
R828 B.n300 B.n299 10.6151
R829 B.n301 B.n300 10.6151
R830 B.n301 B.n90 10.6151
R831 B.n305 B.n90 10.6151
R832 B.n306 B.n305 10.6151
R833 B.n307 B.n306 10.6151
R834 B.n557 B.n0 8.11757
R835 B.n557 B.n1 8.11757
R836 B.n461 B.n460 6.5566
R837 B.n448 B.n42 6.5566
R838 B.n238 B.n237 6.5566
R839 B.n253 B.n252 6.5566
R840 B.n462 B.n461 4.05904
R841 B.n445 B.n42 4.05904
R842 B.n237 B.n236 4.05904
R843 B.n252 B.n106 4.05904
R844 VN.n3 VN.t7 387.705
R845 VN.n13 VN.t5 387.705
R846 VN.n2 VN.t2 366.892
R847 VN.n1 VN.t4 366.892
R848 VN.n6 VN.t3 366.892
R849 VN.n8 VN.t1 366.892
R850 VN.n12 VN.t9 366.892
R851 VN.n11 VN.t6 366.892
R852 VN.n16 VN.t0 366.892
R853 VN.n18 VN.t8 366.892
R854 VN.n9 VN.n8 161.3
R855 VN.n19 VN.n18 161.3
R856 VN.n17 VN.n10 161.3
R857 VN.n7 VN.n0 161.3
R858 VN.n16 VN.n15 80.6037
R859 VN.n14 VN.n11 80.6037
R860 VN.n6 VN.n5 80.6037
R861 VN.n4 VN.n1 80.6037
R862 VN.n2 VN.n1 48.2005
R863 VN.n6 VN.n1 48.2005
R864 VN.n12 VN.n11 48.2005
R865 VN.n16 VN.n11 48.2005
R866 VN VN.n19 41.8471
R867 VN.n7 VN.n6 40.8975
R868 VN.n17 VN.n16 40.8975
R869 VN.n14 VN.n13 31.6317
R870 VN.n4 VN.n3 31.6317
R871 VN.n3 VN.n2 17.5473
R872 VN.n13 VN.n12 17.5473
R873 VN.n8 VN.n7 7.30353
R874 VN.n18 VN.n17 7.30353
R875 VN.n15 VN.n14 0.380177
R876 VN.n5 VN.n4 0.380177
R877 VN.n15 VN.n10 0.285035
R878 VN.n5 VN.n0 0.285035
R879 VN.n19 VN.n10 0.189894
R880 VN.n9 VN.n0 0.189894
R881 VN VN.n9 0.0516364
R882 VDD2.n105 VDD2.n57 756.745
R883 VDD2.n48 VDD2.n0 756.745
R884 VDD2.n106 VDD2.n105 585
R885 VDD2.n104 VDD2.n103 585
R886 VDD2.n61 VDD2.n60 585
R887 VDD2.n98 VDD2.n97 585
R888 VDD2.n96 VDD2.n63 585
R889 VDD2.n95 VDD2.n94 585
R890 VDD2.n66 VDD2.n64 585
R891 VDD2.n89 VDD2.n88 585
R892 VDD2.n87 VDD2.n86 585
R893 VDD2.n70 VDD2.n69 585
R894 VDD2.n81 VDD2.n80 585
R895 VDD2.n79 VDD2.n78 585
R896 VDD2.n74 VDD2.n73 585
R897 VDD2.n16 VDD2.n15 585
R898 VDD2.n21 VDD2.n20 585
R899 VDD2.n23 VDD2.n22 585
R900 VDD2.n12 VDD2.n11 585
R901 VDD2.n29 VDD2.n28 585
R902 VDD2.n31 VDD2.n30 585
R903 VDD2.n8 VDD2.n7 585
R904 VDD2.n38 VDD2.n37 585
R905 VDD2.n39 VDD2.n6 585
R906 VDD2.n41 VDD2.n40 585
R907 VDD2.n4 VDD2.n3 585
R908 VDD2.n47 VDD2.n46 585
R909 VDD2.n49 VDD2.n48 585
R910 VDD2.n17 VDD2.t1 329.038
R911 VDD2.n75 VDD2.t0 329.038
R912 VDD2.n105 VDD2.n104 171.744
R913 VDD2.n104 VDD2.n60 171.744
R914 VDD2.n97 VDD2.n60 171.744
R915 VDD2.n97 VDD2.n96 171.744
R916 VDD2.n96 VDD2.n95 171.744
R917 VDD2.n95 VDD2.n64 171.744
R918 VDD2.n88 VDD2.n64 171.744
R919 VDD2.n88 VDD2.n87 171.744
R920 VDD2.n87 VDD2.n69 171.744
R921 VDD2.n80 VDD2.n69 171.744
R922 VDD2.n80 VDD2.n79 171.744
R923 VDD2.n79 VDD2.n73 171.744
R924 VDD2.n21 VDD2.n15 171.744
R925 VDD2.n22 VDD2.n21 171.744
R926 VDD2.n22 VDD2.n11 171.744
R927 VDD2.n29 VDD2.n11 171.744
R928 VDD2.n30 VDD2.n29 171.744
R929 VDD2.n30 VDD2.n7 171.744
R930 VDD2.n38 VDD2.n7 171.744
R931 VDD2.n39 VDD2.n38 171.744
R932 VDD2.n40 VDD2.n39 171.744
R933 VDD2.n40 VDD2.n3 171.744
R934 VDD2.n47 VDD2.n3 171.744
R935 VDD2.n48 VDD2.n47 171.744
R936 VDD2.t0 VDD2.n73 85.8723
R937 VDD2.t1 VDD2.n15 85.8723
R938 VDD2.n56 VDD2.n55 77.3803
R939 VDD2 VDD2.n113 77.3775
R940 VDD2.n112 VDD2.n111 76.7311
R941 VDD2.n54 VDD2.n53 76.7309
R942 VDD2.n54 VDD2.n52 49.4159
R943 VDD2.n110 VDD2.n109 48.4763
R944 VDD2.n110 VDD2.n56 36.7476
R945 VDD2.n98 VDD2.n63 13.1884
R946 VDD2.n41 VDD2.n6 13.1884
R947 VDD2.n99 VDD2.n61 12.8005
R948 VDD2.n94 VDD2.n65 12.8005
R949 VDD2.n37 VDD2.n36 12.8005
R950 VDD2.n42 VDD2.n4 12.8005
R951 VDD2.n103 VDD2.n102 12.0247
R952 VDD2.n93 VDD2.n66 12.0247
R953 VDD2.n35 VDD2.n8 12.0247
R954 VDD2.n46 VDD2.n45 12.0247
R955 VDD2.n106 VDD2.n59 11.249
R956 VDD2.n90 VDD2.n89 11.249
R957 VDD2.n32 VDD2.n31 11.249
R958 VDD2.n49 VDD2.n2 11.249
R959 VDD2.n75 VDD2.n74 10.7239
R960 VDD2.n17 VDD2.n16 10.7239
R961 VDD2.n107 VDD2.n57 10.4732
R962 VDD2.n86 VDD2.n68 10.4732
R963 VDD2.n28 VDD2.n10 10.4732
R964 VDD2.n50 VDD2.n0 10.4732
R965 VDD2.n85 VDD2.n70 9.69747
R966 VDD2.n27 VDD2.n12 9.69747
R967 VDD2.n109 VDD2.n108 9.45567
R968 VDD2.n52 VDD2.n51 9.45567
R969 VDD2.n77 VDD2.n76 9.3005
R970 VDD2.n72 VDD2.n71 9.3005
R971 VDD2.n83 VDD2.n82 9.3005
R972 VDD2.n85 VDD2.n84 9.3005
R973 VDD2.n68 VDD2.n67 9.3005
R974 VDD2.n91 VDD2.n90 9.3005
R975 VDD2.n93 VDD2.n92 9.3005
R976 VDD2.n65 VDD2.n62 9.3005
R977 VDD2.n108 VDD2.n107 9.3005
R978 VDD2.n59 VDD2.n58 9.3005
R979 VDD2.n102 VDD2.n101 9.3005
R980 VDD2.n100 VDD2.n99 9.3005
R981 VDD2.n51 VDD2.n50 9.3005
R982 VDD2.n2 VDD2.n1 9.3005
R983 VDD2.n45 VDD2.n44 9.3005
R984 VDD2.n43 VDD2.n42 9.3005
R985 VDD2.n19 VDD2.n18 9.3005
R986 VDD2.n14 VDD2.n13 9.3005
R987 VDD2.n25 VDD2.n24 9.3005
R988 VDD2.n27 VDD2.n26 9.3005
R989 VDD2.n10 VDD2.n9 9.3005
R990 VDD2.n33 VDD2.n32 9.3005
R991 VDD2.n35 VDD2.n34 9.3005
R992 VDD2.n36 VDD2.n5 9.3005
R993 VDD2.n82 VDD2.n81 8.92171
R994 VDD2.n24 VDD2.n23 8.92171
R995 VDD2.n78 VDD2.n72 8.14595
R996 VDD2.n20 VDD2.n14 8.14595
R997 VDD2.n77 VDD2.n74 7.3702
R998 VDD2.n19 VDD2.n16 7.3702
R999 VDD2.n78 VDD2.n77 5.81868
R1000 VDD2.n20 VDD2.n19 5.81868
R1001 VDD2.n81 VDD2.n72 5.04292
R1002 VDD2.n23 VDD2.n14 5.04292
R1003 VDD2.n82 VDD2.n70 4.26717
R1004 VDD2.n24 VDD2.n12 4.26717
R1005 VDD2.n109 VDD2.n57 3.49141
R1006 VDD2.n86 VDD2.n85 3.49141
R1007 VDD2.n28 VDD2.n27 3.49141
R1008 VDD2.n52 VDD2.n0 3.49141
R1009 VDD2.n113 VDD2.t7 3.27062
R1010 VDD2.n113 VDD2.t5 3.27062
R1011 VDD2.n111 VDD2.t4 3.27062
R1012 VDD2.n111 VDD2.t3 3.27062
R1013 VDD2.n55 VDD2.t6 3.27062
R1014 VDD2.n55 VDD2.t9 3.27062
R1015 VDD2.n53 VDD2.t8 3.27062
R1016 VDD2.n53 VDD2.t2 3.27062
R1017 VDD2.n107 VDD2.n106 2.71565
R1018 VDD2.n89 VDD2.n68 2.71565
R1019 VDD2.n31 VDD2.n10 2.71565
R1020 VDD2.n50 VDD2.n49 2.71565
R1021 VDD2.n76 VDD2.n75 2.41283
R1022 VDD2.n18 VDD2.n17 2.41283
R1023 VDD2.n103 VDD2.n59 1.93989
R1024 VDD2.n90 VDD2.n66 1.93989
R1025 VDD2.n32 VDD2.n8 1.93989
R1026 VDD2.n46 VDD2.n2 1.93989
R1027 VDD2.n102 VDD2.n61 1.16414
R1028 VDD2.n94 VDD2.n93 1.16414
R1029 VDD2.n37 VDD2.n35 1.16414
R1030 VDD2.n45 VDD2.n4 1.16414
R1031 VDD2.n112 VDD2.n110 0.940155
R1032 VDD2.n99 VDD2.n98 0.388379
R1033 VDD2.n65 VDD2.n63 0.388379
R1034 VDD2.n36 VDD2.n6 0.388379
R1035 VDD2.n42 VDD2.n41 0.388379
R1036 VDD2 VDD2.n112 0.293603
R1037 VDD2.n56 VDD2.n54 0.180068
R1038 VDD2.n108 VDD2.n58 0.155672
R1039 VDD2.n101 VDD2.n58 0.155672
R1040 VDD2.n101 VDD2.n100 0.155672
R1041 VDD2.n100 VDD2.n62 0.155672
R1042 VDD2.n92 VDD2.n62 0.155672
R1043 VDD2.n92 VDD2.n91 0.155672
R1044 VDD2.n91 VDD2.n67 0.155672
R1045 VDD2.n84 VDD2.n67 0.155672
R1046 VDD2.n84 VDD2.n83 0.155672
R1047 VDD2.n83 VDD2.n71 0.155672
R1048 VDD2.n76 VDD2.n71 0.155672
R1049 VDD2.n18 VDD2.n13 0.155672
R1050 VDD2.n25 VDD2.n13 0.155672
R1051 VDD2.n26 VDD2.n25 0.155672
R1052 VDD2.n26 VDD2.n9 0.155672
R1053 VDD2.n33 VDD2.n9 0.155672
R1054 VDD2.n34 VDD2.n33 0.155672
R1055 VDD2.n34 VDD2.n5 0.155672
R1056 VDD2.n43 VDD2.n5 0.155672
R1057 VDD2.n44 VDD2.n43 0.155672
R1058 VDD2.n44 VDD2.n1 0.155672
R1059 VDD2.n51 VDD2.n1 0.155672
R1060 VTAIL.n224 VTAIL.n176 756.745
R1061 VTAIL.n50 VTAIL.n2 756.745
R1062 VTAIL.n170 VTAIL.n122 756.745
R1063 VTAIL.n112 VTAIL.n64 756.745
R1064 VTAIL.n192 VTAIL.n191 585
R1065 VTAIL.n197 VTAIL.n196 585
R1066 VTAIL.n199 VTAIL.n198 585
R1067 VTAIL.n188 VTAIL.n187 585
R1068 VTAIL.n205 VTAIL.n204 585
R1069 VTAIL.n207 VTAIL.n206 585
R1070 VTAIL.n184 VTAIL.n183 585
R1071 VTAIL.n214 VTAIL.n213 585
R1072 VTAIL.n215 VTAIL.n182 585
R1073 VTAIL.n217 VTAIL.n216 585
R1074 VTAIL.n180 VTAIL.n179 585
R1075 VTAIL.n223 VTAIL.n222 585
R1076 VTAIL.n225 VTAIL.n224 585
R1077 VTAIL.n18 VTAIL.n17 585
R1078 VTAIL.n23 VTAIL.n22 585
R1079 VTAIL.n25 VTAIL.n24 585
R1080 VTAIL.n14 VTAIL.n13 585
R1081 VTAIL.n31 VTAIL.n30 585
R1082 VTAIL.n33 VTAIL.n32 585
R1083 VTAIL.n10 VTAIL.n9 585
R1084 VTAIL.n40 VTAIL.n39 585
R1085 VTAIL.n41 VTAIL.n8 585
R1086 VTAIL.n43 VTAIL.n42 585
R1087 VTAIL.n6 VTAIL.n5 585
R1088 VTAIL.n49 VTAIL.n48 585
R1089 VTAIL.n51 VTAIL.n50 585
R1090 VTAIL.n171 VTAIL.n170 585
R1091 VTAIL.n169 VTAIL.n168 585
R1092 VTAIL.n126 VTAIL.n125 585
R1093 VTAIL.n163 VTAIL.n162 585
R1094 VTAIL.n161 VTAIL.n128 585
R1095 VTAIL.n160 VTAIL.n159 585
R1096 VTAIL.n131 VTAIL.n129 585
R1097 VTAIL.n154 VTAIL.n153 585
R1098 VTAIL.n152 VTAIL.n151 585
R1099 VTAIL.n135 VTAIL.n134 585
R1100 VTAIL.n146 VTAIL.n145 585
R1101 VTAIL.n144 VTAIL.n143 585
R1102 VTAIL.n139 VTAIL.n138 585
R1103 VTAIL.n113 VTAIL.n112 585
R1104 VTAIL.n111 VTAIL.n110 585
R1105 VTAIL.n68 VTAIL.n67 585
R1106 VTAIL.n105 VTAIL.n104 585
R1107 VTAIL.n103 VTAIL.n70 585
R1108 VTAIL.n102 VTAIL.n101 585
R1109 VTAIL.n73 VTAIL.n71 585
R1110 VTAIL.n96 VTAIL.n95 585
R1111 VTAIL.n94 VTAIL.n93 585
R1112 VTAIL.n77 VTAIL.n76 585
R1113 VTAIL.n88 VTAIL.n87 585
R1114 VTAIL.n86 VTAIL.n85 585
R1115 VTAIL.n81 VTAIL.n80 585
R1116 VTAIL.n193 VTAIL.t18 329.038
R1117 VTAIL.n19 VTAIL.t2 329.038
R1118 VTAIL.n140 VTAIL.t9 329.038
R1119 VTAIL.n82 VTAIL.t14 329.038
R1120 VTAIL.n197 VTAIL.n191 171.744
R1121 VTAIL.n198 VTAIL.n197 171.744
R1122 VTAIL.n198 VTAIL.n187 171.744
R1123 VTAIL.n205 VTAIL.n187 171.744
R1124 VTAIL.n206 VTAIL.n205 171.744
R1125 VTAIL.n206 VTAIL.n183 171.744
R1126 VTAIL.n214 VTAIL.n183 171.744
R1127 VTAIL.n215 VTAIL.n214 171.744
R1128 VTAIL.n216 VTAIL.n215 171.744
R1129 VTAIL.n216 VTAIL.n179 171.744
R1130 VTAIL.n223 VTAIL.n179 171.744
R1131 VTAIL.n224 VTAIL.n223 171.744
R1132 VTAIL.n23 VTAIL.n17 171.744
R1133 VTAIL.n24 VTAIL.n23 171.744
R1134 VTAIL.n24 VTAIL.n13 171.744
R1135 VTAIL.n31 VTAIL.n13 171.744
R1136 VTAIL.n32 VTAIL.n31 171.744
R1137 VTAIL.n32 VTAIL.n9 171.744
R1138 VTAIL.n40 VTAIL.n9 171.744
R1139 VTAIL.n41 VTAIL.n40 171.744
R1140 VTAIL.n42 VTAIL.n41 171.744
R1141 VTAIL.n42 VTAIL.n5 171.744
R1142 VTAIL.n49 VTAIL.n5 171.744
R1143 VTAIL.n50 VTAIL.n49 171.744
R1144 VTAIL.n170 VTAIL.n169 171.744
R1145 VTAIL.n169 VTAIL.n125 171.744
R1146 VTAIL.n162 VTAIL.n125 171.744
R1147 VTAIL.n162 VTAIL.n161 171.744
R1148 VTAIL.n161 VTAIL.n160 171.744
R1149 VTAIL.n160 VTAIL.n129 171.744
R1150 VTAIL.n153 VTAIL.n129 171.744
R1151 VTAIL.n153 VTAIL.n152 171.744
R1152 VTAIL.n152 VTAIL.n134 171.744
R1153 VTAIL.n145 VTAIL.n134 171.744
R1154 VTAIL.n145 VTAIL.n144 171.744
R1155 VTAIL.n144 VTAIL.n138 171.744
R1156 VTAIL.n112 VTAIL.n111 171.744
R1157 VTAIL.n111 VTAIL.n67 171.744
R1158 VTAIL.n104 VTAIL.n67 171.744
R1159 VTAIL.n104 VTAIL.n103 171.744
R1160 VTAIL.n103 VTAIL.n102 171.744
R1161 VTAIL.n102 VTAIL.n71 171.744
R1162 VTAIL.n95 VTAIL.n71 171.744
R1163 VTAIL.n95 VTAIL.n94 171.744
R1164 VTAIL.n94 VTAIL.n76 171.744
R1165 VTAIL.n87 VTAIL.n76 171.744
R1166 VTAIL.n87 VTAIL.n86 171.744
R1167 VTAIL.n86 VTAIL.n80 171.744
R1168 VTAIL.t18 VTAIL.n191 85.8723
R1169 VTAIL.t2 VTAIL.n17 85.8723
R1170 VTAIL.t9 VTAIL.n138 85.8723
R1171 VTAIL.t14 VTAIL.n80 85.8723
R1172 VTAIL.n121 VTAIL.n120 60.0523
R1173 VTAIL.n119 VTAIL.n118 60.0523
R1174 VTAIL.n63 VTAIL.n62 60.0523
R1175 VTAIL.n61 VTAIL.n60 60.0523
R1176 VTAIL.n231 VTAIL.n230 60.0521
R1177 VTAIL.n1 VTAIL.n0 60.0521
R1178 VTAIL.n57 VTAIL.n56 60.0521
R1179 VTAIL.n59 VTAIL.n58 60.0521
R1180 VTAIL.n229 VTAIL.n228 31.7975
R1181 VTAIL.n55 VTAIL.n54 31.7975
R1182 VTAIL.n175 VTAIL.n174 31.7975
R1183 VTAIL.n117 VTAIL.n116 31.7975
R1184 VTAIL.n61 VTAIL.n59 22.8152
R1185 VTAIL.n229 VTAIL.n175 21.8755
R1186 VTAIL.n217 VTAIL.n182 13.1884
R1187 VTAIL.n43 VTAIL.n8 13.1884
R1188 VTAIL.n163 VTAIL.n128 13.1884
R1189 VTAIL.n105 VTAIL.n70 13.1884
R1190 VTAIL.n213 VTAIL.n212 12.8005
R1191 VTAIL.n218 VTAIL.n180 12.8005
R1192 VTAIL.n39 VTAIL.n38 12.8005
R1193 VTAIL.n44 VTAIL.n6 12.8005
R1194 VTAIL.n164 VTAIL.n126 12.8005
R1195 VTAIL.n159 VTAIL.n130 12.8005
R1196 VTAIL.n106 VTAIL.n68 12.8005
R1197 VTAIL.n101 VTAIL.n72 12.8005
R1198 VTAIL.n211 VTAIL.n184 12.0247
R1199 VTAIL.n222 VTAIL.n221 12.0247
R1200 VTAIL.n37 VTAIL.n10 12.0247
R1201 VTAIL.n48 VTAIL.n47 12.0247
R1202 VTAIL.n168 VTAIL.n167 12.0247
R1203 VTAIL.n158 VTAIL.n131 12.0247
R1204 VTAIL.n110 VTAIL.n109 12.0247
R1205 VTAIL.n100 VTAIL.n73 12.0247
R1206 VTAIL.n208 VTAIL.n207 11.249
R1207 VTAIL.n225 VTAIL.n178 11.249
R1208 VTAIL.n34 VTAIL.n33 11.249
R1209 VTAIL.n51 VTAIL.n4 11.249
R1210 VTAIL.n171 VTAIL.n124 11.249
R1211 VTAIL.n155 VTAIL.n154 11.249
R1212 VTAIL.n113 VTAIL.n66 11.249
R1213 VTAIL.n97 VTAIL.n96 11.249
R1214 VTAIL.n193 VTAIL.n192 10.7239
R1215 VTAIL.n19 VTAIL.n18 10.7239
R1216 VTAIL.n140 VTAIL.n139 10.7239
R1217 VTAIL.n82 VTAIL.n81 10.7239
R1218 VTAIL.n204 VTAIL.n186 10.4732
R1219 VTAIL.n226 VTAIL.n176 10.4732
R1220 VTAIL.n30 VTAIL.n12 10.4732
R1221 VTAIL.n52 VTAIL.n2 10.4732
R1222 VTAIL.n172 VTAIL.n122 10.4732
R1223 VTAIL.n151 VTAIL.n133 10.4732
R1224 VTAIL.n114 VTAIL.n64 10.4732
R1225 VTAIL.n93 VTAIL.n75 10.4732
R1226 VTAIL.n203 VTAIL.n188 9.69747
R1227 VTAIL.n29 VTAIL.n14 9.69747
R1228 VTAIL.n150 VTAIL.n135 9.69747
R1229 VTAIL.n92 VTAIL.n77 9.69747
R1230 VTAIL.n228 VTAIL.n227 9.45567
R1231 VTAIL.n54 VTAIL.n53 9.45567
R1232 VTAIL.n174 VTAIL.n173 9.45567
R1233 VTAIL.n116 VTAIL.n115 9.45567
R1234 VTAIL.n227 VTAIL.n226 9.3005
R1235 VTAIL.n178 VTAIL.n177 9.3005
R1236 VTAIL.n221 VTAIL.n220 9.3005
R1237 VTAIL.n219 VTAIL.n218 9.3005
R1238 VTAIL.n195 VTAIL.n194 9.3005
R1239 VTAIL.n190 VTAIL.n189 9.3005
R1240 VTAIL.n201 VTAIL.n200 9.3005
R1241 VTAIL.n203 VTAIL.n202 9.3005
R1242 VTAIL.n186 VTAIL.n185 9.3005
R1243 VTAIL.n209 VTAIL.n208 9.3005
R1244 VTAIL.n211 VTAIL.n210 9.3005
R1245 VTAIL.n212 VTAIL.n181 9.3005
R1246 VTAIL.n53 VTAIL.n52 9.3005
R1247 VTAIL.n4 VTAIL.n3 9.3005
R1248 VTAIL.n47 VTAIL.n46 9.3005
R1249 VTAIL.n45 VTAIL.n44 9.3005
R1250 VTAIL.n21 VTAIL.n20 9.3005
R1251 VTAIL.n16 VTAIL.n15 9.3005
R1252 VTAIL.n27 VTAIL.n26 9.3005
R1253 VTAIL.n29 VTAIL.n28 9.3005
R1254 VTAIL.n12 VTAIL.n11 9.3005
R1255 VTAIL.n35 VTAIL.n34 9.3005
R1256 VTAIL.n37 VTAIL.n36 9.3005
R1257 VTAIL.n38 VTAIL.n7 9.3005
R1258 VTAIL.n142 VTAIL.n141 9.3005
R1259 VTAIL.n137 VTAIL.n136 9.3005
R1260 VTAIL.n148 VTAIL.n147 9.3005
R1261 VTAIL.n150 VTAIL.n149 9.3005
R1262 VTAIL.n133 VTAIL.n132 9.3005
R1263 VTAIL.n156 VTAIL.n155 9.3005
R1264 VTAIL.n158 VTAIL.n157 9.3005
R1265 VTAIL.n130 VTAIL.n127 9.3005
R1266 VTAIL.n173 VTAIL.n172 9.3005
R1267 VTAIL.n124 VTAIL.n123 9.3005
R1268 VTAIL.n167 VTAIL.n166 9.3005
R1269 VTAIL.n165 VTAIL.n164 9.3005
R1270 VTAIL.n84 VTAIL.n83 9.3005
R1271 VTAIL.n79 VTAIL.n78 9.3005
R1272 VTAIL.n90 VTAIL.n89 9.3005
R1273 VTAIL.n92 VTAIL.n91 9.3005
R1274 VTAIL.n75 VTAIL.n74 9.3005
R1275 VTAIL.n98 VTAIL.n97 9.3005
R1276 VTAIL.n100 VTAIL.n99 9.3005
R1277 VTAIL.n72 VTAIL.n69 9.3005
R1278 VTAIL.n115 VTAIL.n114 9.3005
R1279 VTAIL.n66 VTAIL.n65 9.3005
R1280 VTAIL.n109 VTAIL.n108 9.3005
R1281 VTAIL.n107 VTAIL.n106 9.3005
R1282 VTAIL.n200 VTAIL.n199 8.92171
R1283 VTAIL.n26 VTAIL.n25 8.92171
R1284 VTAIL.n147 VTAIL.n146 8.92171
R1285 VTAIL.n89 VTAIL.n88 8.92171
R1286 VTAIL.n196 VTAIL.n190 8.14595
R1287 VTAIL.n22 VTAIL.n16 8.14595
R1288 VTAIL.n143 VTAIL.n137 8.14595
R1289 VTAIL.n85 VTAIL.n79 8.14595
R1290 VTAIL.n195 VTAIL.n192 7.3702
R1291 VTAIL.n21 VTAIL.n18 7.3702
R1292 VTAIL.n142 VTAIL.n139 7.3702
R1293 VTAIL.n84 VTAIL.n81 7.3702
R1294 VTAIL.n196 VTAIL.n195 5.81868
R1295 VTAIL.n22 VTAIL.n21 5.81868
R1296 VTAIL.n143 VTAIL.n142 5.81868
R1297 VTAIL.n85 VTAIL.n84 5.81868
R1298 VTAIL.n199 VTAIL.n190 5.04292
R1299 VTAIL.n25 VTAIL.n16 5.04292
R1300 VTAIL.n146 VTAIL.n137 5.04292
R1301 VTAIL.n88 VTAIL.n79 5.04292
R1302 VTAIL.n200 VTAIL.n188 4.26717
R1303 VTAIL.n26 VTAIL.n14 4.26717
R1304 VTAIL.n147 VTAIL.n135 4.26717
R1305 VTAIL.n89 VTAIL.n77 4.26717
R1306 VTAIL.n204 VTAIL.n203 3.49141
R1307 VTAIL.n228 VTAIL.n176 3.49141
R1308 VTAIL.n30 VTAIL.n29 3.49141
R1309 VTAIL.n54 VTAIL.n2 3.49141
R1310 VTAIL.n174 VTAIL.n122 3.49141
R1311 VTAIL.n151 VTAIL.n150 3.49141
R1312 VTAIL.n116 VTAIL.n64 3.49141
R1313 VTAIL.n93 VTAIL.n92 3.49141
R1314 VTAIL.n230 VTAIL.t15 3.27062
R1315 VTAIL.n230 VTAIL.t16 3.27062
R1316 VTAIL.n0 VTAIL.t12 3.27062
R1317 VTAIL.n0 VTAIL.t17 3.27062
R1318 VTAIL.n56 VTAIL.t5 3.27062
R1319 VTAIL.n56 VTAIL.t6 3.27062
R1320 VTAIL.n58 VTAIL.t1 3.27062
R1321 VTAIL.n58 VTAIL.t3 3.27062
R1322 VTAIL.n120 VTAIL.t0 3.27062
R1323 VTAIL.n120 VTAIL.t4 3.27062
R1324 VTAIL.n118 VTAIL.t8 3.27062
R1325 VTAIL.n118 VTAIL.t7 3.27062
R1326 VTAIL.n62 VTAIL.t13 3.27062
R1327 VTAIL.n62 VTAIL.t10 3.27062
R1328 VTAIL.n60 VTAIL.t11 3.27062
R1329 VTAIL.n60 VTAIL.t19 3.27062
R1330 VTAIL.n207 VTAIL.n186 2.71565
R1331 VTAIL.n226 VTAIL.n225 2.71565
R1332 VTAIL.n33 VTAIL.n12 2.71565
R1333 VTAIL.n52 VTAIL.n51 2.71565
R1334 VTAIL.n172 VTAIL.n171 2.71565
R1335 VTAIL.n154 VTAIL.n133 2.71565
R1336 VTAIL.n114 VTAIL.n113 2.71565
R1337 VTAIL.n96 VTAIL.n75 2.71565
R1338 VTAIL.n194 VTAIL.n193 2.41283
R1339 VTAIL.n20 VTAIL.n19 2.41283
R1340 VTAIL.n141 VTAIL.n140 2.41283
R1341 VTAIL.n83 VTAIL.n82 2.41283
R1342 VTAIL.n208 VTAIL.n184 1.93989
R1343 VTAIL.n222 VTAIL.n178 1.93989
R1344 VTAIL.n34 VTAIL.n10 1.93989
R1345 VTAIL.n48 VTAIL.n4 1.93989
R1346 VTAIL.n168 VTAIL.n124 1.93989
R1347 VTAIL.n155 VTAIL.n131 1.93989
R1348 VTAIL.n110 VTAIL.n66 1.93989
R1349 VTAIL.n97 VTAIL.n73 1.93989
R1350 VTAIL.n213 VTAIL.n211 1.16414
R1351 VTAIL.n221 VTAIL.n180 1.16414
R1352 VTAIL.n39 VTAIL.n37 1.16414
R1353 VTAIL.n47 VTAIL.n6 1.16414
R1354 VTAIL.n167 VTAIL.n126 1.16414
R1355 VTAIL.n159 VTAIL.n158 1.16414
R1356 VTAIL.n109 VTAIL.n68 1.16414
R1357 VTAIL.n101 VTAIL.n100 1.16414
R1358 VTAIL.n63 VTAIL.n61 0.940155
R1359 VTAIL.n117 VTAIL.n63 0.940155
R1360 VTAIL.n119 VTAIL.n117 0.940155
R1361 VTAIL.n121 VTAIL.n119 0.940155
R1362 VTAIL.n175 VTAIL.n121 0.940155
R1363 VTAIL.n59 VTAIL.n57 0.940155
R1364 VTAIL.n57 VTAIL.n55 0.940155
R1365 VTAIL.n55 VTAIL.n1 0.940155
R1366 VTAIL.n231 VTAIL.n229 0.940155
R1367 VTAIL VTAIL.n1 0.763431
R1368 VTAIL.n212 VTAIL.n182 0.388379
R1369 VTAIL.n218 VTAIL.n217 0.388379
R1370 VTAIL.n38 VTAIL.n8 0.388379
R1371 VTAIL.n44 VTAIL.n43 0.388379
R1372 VTAIL.n164 VTAIL.n163 0.388379
R1373 VTAIL.n130 VTAIL.n128 0.388379
R1374 VTAIL.n106 VTAIL.n105 0.388379
R1375 VTAIL.n72 VTAIL.n70 0.388379
R1376 VTAIL VTAIL.n231 0.177224
R1377 VTAIL.n194 VTAIL.n189 0.155672
R1378 VTAIL.n201 VTAIL.n189 0.155672
R1379 VTAIL.n202 VTAIL.n201 0.155672
R1380 VTAIL.n202 VTAIL.n185 0.155672
R1381 VTAIL.n209 VTAIL.n185 0.155672
R1382 VTAIL.n210 VTAIL.n209 0.155672
R1383 VTAIL.n210 VTAIL.n181 0.155672
R1384 VTAIL.n219 VTAIL.n181 0.155672
R1385 VTAIL.n220 VTAIL.n219 0.155672
R1386 VTAIL.n220 VTAIL.n177 0.155672
R1387 VTAIL.n227 VTAIL.n177 0.155672
R1388 VTAIL.n20 VTAIL.n15 0.155672
R1389 VTAIL.n27 VTAIL.n15 0.155672
R1390 VTAIL.n28 VTAIL.n27 0.155672
R1391 VTAIL.n28 VTAIL.n11 0.155672
R1392 VTAIL.n35 VTAIL.n11 0.155672
R1393 VTAIL.n36 VTAIL.n35 0.155672
R1394 VTAIL.n36 VTAIL.n7 0.155672
R1395 VTAIL.n45 VTAIL.n7 0.155672
R1396 VTAIL.n46 VTAIL.n45 0.155672
R1397 VTAIL.n46 VTAIL.n3 0.155672
R1398 VTAIL.n53 VTAIL.n3 0.155672
R1399 VTAIL.n173 VTAIL.n123 0.155672
R1400 VTAIL.n166 VTAIL.n123 0.155672
R1401 VTAIL.n166 VTAIL.n165 0.155672
R1402 VTAIL.n165 VTAIL.n127 0.155672
R1403 VTAIL.n157 VTAIL.n127 0.155672
R1404 VTAIL.n157 VTAIL.n156 0.155672
R1405 VTAIL.n156 VTAIL.n132 0.155672
R1406 VTAIL.n149 VTAIL.n132 0.155672
R1407 VTAIL.n149 VTAIL.n148 0.155672
R1408 VTAIL.n148 VTAIL.n136 0.155672
R1409 VTAIL.n141 VTAIL.n136 0.155672
R1410 VTAIL.n115 VTAIL.n65 0.155672
R1411 VTAIL.n108 VTAIL.n65 0.155672
R1412 VTAIL.n108 VTAIL.n107 0.155672
R1413 VTAIL.n107 VTAIL.n69 0.155672
R1414 VTAIL.n99 VTAIL.n69 0.155672
R1415 VTAIL.n99 VTAIL.n98 0.155672
R1416 VTAIL.n98 VTAIL.n74 0.155672
R1417 VTAIL.n91 VTAIL.n74 0.155672
R1418 VTAIL.n91 VTAIL.n90 0.155672
R1419 VTAIL.n90 VTAIL.n78 0.155672
R1420 VTAIL.n83 VTAIL.n78 0.155672
R1421 VP.n6 VP.t0 387.705
R1422 VP.n14 VP.t7 366.892
R1423 VP.n16 VP.t5 366.892
R1424 VP.n1 VP.t6 366.892
R1425 VP.n20 VP.t3 366.892
R1426 VP.n22 VP.t4 366.892
R1427 VP.n11 VP.t1 366.892
R1428 VP.n9 VP.t9 366.892
R1429 VP.n8 VP.t2 366.892
R1430 VP.n7 VP.t8 366.892
R1431 VP.n23 VP.n22 161.3
R1432 VP.n10 VP.n3 161.3
R1433 VP.n12 VP.n11 161.3
R1434 VP.n21 VP.n0 161.3
R1435 VP.n15 VP.n2 161.3
R1436 VP.n14 VP.n13 161.3
R1437 VP.n8 VP.n5 80.6037
R1438 VP.n9 VP.n4 80.6037
R1439 VP.n20 VP.n19 80.6037
R1440 VP.n18 VP.n1 80.6037
R1441 VP.n17 VP.n16 80.6037
R1442 VP.n16 VP.n1 48.2005
R1443 VP.n20 VP.n1 48.2005
R1444 VP.n9 VP.n8 48.2005
R1445 VP.n8 VP.n7 48.2005
R1446 VP.n13 VP.n12 41.4664
R1447 VP.n16 VP.n15 40.8975
R1448 VP.n21 VP.n20 40.8975
R1449 VP.n10 VP.n9 40.8975
R1450 VP.n6 VP.n5 31.6317
R1451 VP.n7 VP.n6 17.5473
R1452 VP.n15 VP.n14 7.30353
R1453 VP.n22 VP.n21 7.30353
R1454 VP.n11 VP.n10 7.30353
R1455 VP.n5 VP.n4 0.380177
R1456 VP.n18 VP.n17 0.380177
R1457 VP.n19 VP.n18 0.380177
R1458 VP.n4 VP.n3 0.285035
R1459 VP.n17 VP.n2 0.285035
R1460 VP.n19 VP.n0 0.285035
R1461 VP.n12 VP.n3 0.189894
R1462 VP.n13 VP.n2 0.189894
R1463 VP.n23 VP.n0 0.189894
R1464 VP VP.n23 0.0516364
R1465 VDD1.n48 VDD1.n0 756.745
R1466 VDD1.n103 VDD1.n55 756.745
R1467 VDD1.n49 VDD1.n48 585
R1468 VDD1.n47 VDD1.n46 585
R1469 VDD1.n4 VDD1.n3 585
R1470 VDD1.n41 VDD1.n40 585
R1471 VDD1.n39 VDD1.n6 585
R1472 VDD1.n38 VDD1.n37 585
R1473 VDD1.n9 VDD1.n7 585
R1474 VDD1.n32 VDD1.n31 585
R1475 VDD1.n30 VDD1.n29 585
R1476 VDD1.n13 VDD1.n12 585
R1477 VDD1.n24 VDD1.n23 585
R1478 VDD1.n22 VDD1.n21 585
R1479 VDD1.n17 VDD1.n16 585
R1480 VDD1.n71 VDD1.n70 585
R1481 VDD1.n76 VDD1.n75 585
R1482 VDD1.n78 VDD1.n77 585
R1483 VDD1.n67 VDD1.n66 585
R1484 VDD1.n84 VDD1.n83 585
R1485 VDD1.n86 VDD1.n85 585
R1486 VDD1.n63 VDD1.n62 585
R1487 VDD1.n93 VDD1.n92 585
R1488 VDD1.n94 VDD1.n61 585
R1489 VDD1.n96 VDD1.n95 585
R1490 VDD1.n59 VDD1.n58 585
R1491 VDD1.n102 VDD1.n101 585
R1492 VDD1.n104 VDD1.n103 585
R1493 VDD1.n72 VDD1.t2 329.038
R1494 VDD1.n18 VDD1.t9 329.038
R1495 VDD1.n48 VDD1.n47 171.744
R1496 VDD1.n47 VDD1.n3 171.744
R1497 VDD1.n40 VDD1.n3 171.744
R1498 VDD1.n40 VDD1.n39 171.744
R1499 VDD1.n39 VDD1.n38 171.744
R1500 VDD1.n38 VDD1.n7 171.744
R1501 VDD1.n31 VDD1.n7 171.744
R1502 VDD1.n31 VDD1.n30 171.744
R1503 VDD1.n30 VDD1.n12 171.744
R1504 VDD1.n23 VDD1.n12 171.744
R1505 VDD1.n23 VDD1.n22 171.744
R1506 VDD1.n22 VDD1.n16 171.744
R1507 VDD1.n76 VDD1.n70 171.744
R1508 VDD1.n77 VDD1.n76 171.744
R1509 VDD1.n77 VDD1.n66 171.744
R1510 VDD1.n84 VDD1.n66 171.744
R1511 VDD1.n85 VDD1.n84 171.744
R1512 VDD1.n85 VDD1.n62 171.744
R1513 VDD1.n93 VDD1.n62 171.744
R1514 VDD1.n94 VDD1.n93 171.744
R1515 VDD1.n95 VDD1.n94 171.744
R1516 VDD1.n95 VDD1.n58 171.744
R1517 VDD1.n102 VDD1.n58 171.744
R1518 VDD1.n103 VDD1.n102 171.744
R1519 VDD1.t9 VDD1.n16 85.8723
R1520 VDD1.t2 VDD1.n70 85.8723
R1521 VDD1.n111 VDD1.n110 77.3803
R1522 VDD1.n54 VDD1.n53 76.7311
R1523 VDD1.n113 VDD1.n112 76.7309
R1524 VDD1.n109 VDD1.n108 76.7309
R1525 VDD1.n54 VDD1.n52 49.4159
R1526 VDD1.n109 VDD1.n107 49.4159
R1527 VDD1.n113 VDD1.n111 37.8005
R1528 VDD1.n41 VDD1.n6 13.1884
R1529 VDD1.n96 VDD1.n61 13.1884
R1530 VDD1.n42 VDD1.n4 12.8005
R1531 VDD1.n37 VDD1.n8 12.8005
R1532 VDD1.n92 VDD1.n91 12.8005
R1533 VDD1.n97 VDD1.n59 12.8005
R1534 VDD1.n46 VDD1.n45 12.0247
R1535 VDD1.n36 VDD1.n9 12.0247
R1536 VDD1.n90 VDD1.n63 12.0247
R1537 VDD1.n101 VDD1.n100 12.0247
R1538 VDD1.n49 VDD1.n2 11.249
R1539 VDD1.n33 VDD1.n32 11.249
R1540 VDD1.n87 VDD1.n86 11.249
R1541 VDD1.n104 VDD1.n57 11.249
R1542 VDD1.n18 VDD1.n17 10.7239
R1543 VDD1.n72 VDD1.n71 10.7239
R1544 VDD1.n50 VDD1.n0 10.4732
R1545 VDD1.n29 VDD1.n11 10.4732
R1546 VDD1.n83 VDD1.n65 10.4732
R1547 VDD1.n105 VDD1.n55 10.4732
R1548 VDD1.n28 VDD1.n13 9.69747
R1549 VDD1.n82 VDD1.n67 9.69747
R1550 VDD1.n52 VDD1.n51 9.45567
R1551 VDD1.n107 VDD1.n106 9.45567
R1552 VDD1.n20 VDD1.n19 9.3005
R1553 VDD1.n15 VDD1.n14 9.3005
R1554 VDD1.n26 VDD1.n25 9.3005
R1555 VDD1.n28 VDD1.n27 9.3005
R1556 VDD1.n11 VDD1.n10 9.3005
R1557 VDD1.n34 VDD1.n33 9.3005
R1558 VDD1.n36 VDD1.n35 9.3005
R1559 VDD1.n8 VDD1.n5 9.3005
R1560 VDD1.n51 VDD1.n50 9.3005
R1561 VDD1.n2 VDD1.n1 9.3005
R1562 VDD1.n45 VDD1.n44 9.3005
R1563 VDD1.n43 VDD1.n42 9.3005
R1564 VDD1.n106 VDD1.n105 9.3005
R1565 VDD1.n57 VDD1.n56 9.3005
R1566 VDD1.n100 VDD1.n99 9.3005
R1567 VDD1.n98 VDD1.n97 9.3005
R1568 VDD1.n74 VDD1.n73 9.3005
R1569 VDD1.n69 VDD1.n68 9.3005
R1570 VDD1.n80 VDD1.n79 9.3005
R1571 VDD1.n82 VDD1.n81 9.3005
R1572 VDD1.n65 VDD1.n64 9.3005
R1573 VDD1.n88 VDD1.n87 9.3005
R1574 VDD1.n90 VDD1.n89 9.3005
R1575 VDD1.n91 VDD1.n60 9.3005
R1576 VDD1.n25 VDD1.n24 8.92171
R1577 VDD1.n79 VDD1.n78 8.92171
R1578 VDD1.n21 VDD1.n15 8.14595
R1579 VDD1.n75 VDD1.n69 8.14595
R1580 VDD1.n20 VDD1.n17 7.3702
R1581 VDD1.n74 VDD1.n71 7.3702
R1582 VDD1.n21 VDD1.n20 5.81868
R1583 VDD1.n75 VDD1.n74 5.81868
R1584 VDD1.n24 VDD1.n15 5.04292
R1585 VDD1.n78 VDD1.n69 5.04292
R1586 VDD1.n25 VDD1.n13 4.26717
R1587 VDD1.n79 VDD1.n67 4.26717
R1588 VDD1.n52 VDD1.n0 3.49141
R1589 VDD1.n29 VDD1.n28 3.49141
R1590 VDD1.n83 VDD1.n82 3.49141
R1591 VDD1.n107 VDD1.n55 3.49141
R1592 VDD1.n112 VDD1.t0 3.27062
R1593 VDD1.n112 VDD1.t8 3.27062
R1594 VDD1.n53 VDD1.t1 3.27062
R1595 VDD1.n53 VDD1.t7 3.27062
R1596 VDD1.n110 VDD1.t6 3.27062
R1597 VDD1.n110 VDD1.t5 3.27062
R1598 VDD1.n108 VDD1.t4 3.27062
R1599 VDD1.n108 VDD1.t3 3.27062
R1600 VDD1.n50 VDD1.n49 2.71565
R1601 VDD1.n32 VDD1.n11 2.71565
R1602 VDD1.n86 VDD1.n65 2.71565
R1603 VDD1.n105 VDD1.n104 2.71565
R1604 VDD1.n19 VDD1.n18 2.41283
R1605 VDD1.n73 VDD1.n72 2.41283
R1606 VDD1.n46 VDD1.n2 1.93989
R1607 VDD1.n33 VDD1.n9 1.93989
R1608 VDD1.n87 VDD1.n63 1.93989
R1609 VDD1.n101 VDD1.n57 1.93989
R1610 VDD1.n45 VDD1.n4 1.16414
R1611 VDD1.n37 VDD1.n36 1.16414
R1612 VDD1.n92 VDD1.n90 1.16414
R1613 VDD1.n100 VDD1.n59 1.16414
R1614 VDD1 VDD1.n113 0.647052
R1615 VDD1.n42 VDD1.n41 0.388379
R1616 VDD1.n8 VDD1.n6 0.388379
R1617 VDD1.n91 VDD1.n61 0.388379
R1618 VDD1.n97 VDD1.n96 0.388379
R1619 VDD1 VDD1.n54 0.293603
R1620 VDD1.n111 VDD1.n109 0.180068
R1621 VDD1.n51 VDD1.n1 0.155672
R1622 VDD1.n44 VDD1.n1 0.155672
R1623 VDD1.n44 VDD1.n43 0.155672
R1624 VDD1.n43 VDD1.n5 0.155672
R1625 VDD1.n35 VDD1.n5 0.155672
R1626 VDD1.n35 VDD1.n34 0.155672
R1627 VDD1.n34 VDD1.n10 0.155672
R1628 VDD1.n27 VDD1.n10 0.155672
R1629 VDD1.n27 VDD1.n26 0.155672
R1630 VDD1.n26 VDD1.n14 0.155672
R1631 VDD1.n19 VDD1.n14 0.155672
R1632 VDD1.n73 VDD1.n68 0.155672
R1633 VDD1.n80 VDD1.n68 0.155672
R1634 VDD1.n81 VDD1.n80 0.155672
R1635 VDD1.n81 VDD1.n64 0.155672
R1636 VDD1.n88 VDD1.n64 0.155672
R1637 VDD1.n89 VDD1.n88 0.155672
R1638 VDD1.n89 VDD1.n60 0.155672
R1639 VDD1.n98 VDD1.n60 0.155672
R1640 VDD1.n99 VDD1.n98 0.155672
R1641 VDD1.n99 VDD1.n56 0.155672
R1642 VDD1.n106 VDD1.n56 0.155672
C0 VP w_n2278_n2956# 4.56728f
C1 VTAIL B 2.40071f
C2 VTAIL VDD2 11.845901f
C3 VN VP 5.30475f
C4 B w_n2278_n2956# 6.87722f
C5 VDD2 w_n2278_n2956# 1.96427f
C6 VN B 0.791923f
C7 VN VDD2 5.85425f
C8 VTAIL w_n2278_n2956# 2.6989f
C9 VDD1 VP 6.05005f
C10 VTAIL VN 5.80212f
C11 VDD1 B 1.57903f
C12 VDD1 VDD2 1.00973f
C13 VN w_n2278_n2956# 4.27637f
C14 VTAIL VDD1 11.8099f
C15 VDD1 w_n2278_n2956# 1.91657f
C16 VP B 1.27095f
C17 VDD1 VN 0.149518f
C18 VP VDD2 0.349262f
C19 VDD2 B 1.62561f
C20 VTAIL VP 5.81662f
C21 VDD2 VSUBS 1.326265f
C22 VDD1 VSUBS 1.113464f
C23 VTAIL VSUBS 0.740993f
C24 VN VSUBS 4.848f
C25 VP VSUBS 1.815084f
C26 B VSUBS 2.910527f
C27 w_n2278_n2956# VSUBS 83.183395f
C28 VDD1.n0 VSUBS 0.02517f
C29 VDD1.n1 VSUBS 0.024313f
C30 VDD1.n2 VSUBS 0.013065f
C31 VDD1.n3 VSUBS 0.03088f
C32 VDD1.n4 VSUBS 0.013833f
C33 VDD1.n5 VSUBS 0.024313f
C34 VDD1.n6 VSUBS 0.013449f
C35 VDD1.n7 VSUBS 0.03088f
C36 VDD1.n8 VSUBS 0.013065f
C37 VDD1.n9 VSUBS 0.013833f
C38 VDD1.n10 VSUBS 0.024313f
C39 VDD1.n11 VSUBS 0.013065f
C40 VDD1.n12 VSUBS 0.03088f
C41 VDD1.n13 VSUBS 0.013833f
C42 VDD1.n14 VSUBS 0.024313f
C43 VDD1.n15 VSUBS 0.013065f
C44 VDD1.n16 VSUBS 0.02316f
C45 VDD1.n17 VSUBS 0.02323f
C46 VDD1.t9 VSUBS 0.066389f
C47 VDD1.n18 VSUBS 0.168846f
C48 VDD1.n19 VSUBS 0.975096f
C49 VDD1.n20 VSUBS 0.013065f
C50 VDD1.n21 VSUBS 0.013833f
C51 VDD1.n22 VSUBS 0.03088f
C52 VDD1.n23 VSUBS 0.03088f
C53 VDD1.n24 VSUBS 0.013833f
C54 VDD1.n25 VSUBS 0.013065f
C55 VDD1.n26 VSUBS 0.024313f
C56 VDD1.n27 VSUBS 0.024313f
C57 VDD1.n28 VSUBS 0.013065f
C58 VDD1.n29 VSUBS 0.013833f
C59 VDD1.n30 VSUBS 0.03088f
C60 VDD1.n31 VSUBS 0.03088f
C61 VDD1.n32 VSUBS 0.013833f
C62 VDD1.n33 VSUBS 0.013065f
C63 VDD1.n34 VSUBS 0.024313f
C64 VDD1.n35 VSUBS 0.024313f
C65 VDD1.n36 VSUBS 0.013065f
C66 VDD1.n37 VSUBS 0.013833f
C67 VDD1.n38 VSUBS 0.03088f
C68 VDD1.n39 VSUBS 0.03088f
C69 VDD1.n40 VSUBS 0.03088f
C70 VDD1.n41 VSUBS 0.013449f
C71 VDD1.n42 VSUBS 0.013065f
C72 VDD1.n43 VSUBS 0.024313f
C73 VDD1.n44 VSUBS 0.024313f
C74 VDD1.n45 VSUBS 0.013065f
C75 VDD1.n46 VSUBS 0.013833f
C76 VDD1.n47 VSUBS 0.03088f
C77 VDD1.n48 VSUBS 0.069497f
C78 VDD1.n49 VSUBS 0.013833f
C79 VDD1.n50 VSUBS 0.013065f
C80 VDD1.n51 VSUBS 0.055534f
C81 VDD1.n52 VSUBS 0.053771f
C82 VDD1.t1 VSUBS 0.190976f
C83 VDD1.t7 VSUBS 0.190976f
C84 VDD1.n53 VSUBS 1.43899f
C85 VDD1.n54 VSUBS 0.654383f
C86 VDD1.n55 VSUBS 0.02517f
C87 VDD1.n56 VSUBS 0.024313f
C88 VDD1.n57 VSUBS 0.013065f
C89 VDD1.n58 VSUBS 0.03088f
C90 VDD1.n59 VSUBS 0.013833f
C91 VDD1.n60 VSUBS 0.024313f
C92 VDD1.n61 VSUBS 0.013449f
C93 VDD1.n62 VSUBS 0.03088f
C94 VDD1.n63 VSUBS 0.013833f
C95 VDD1.n64 VSUBS 0.024313f
C96 VDD1.n65 VSUBS 0.013065f
C97 VDD1.n66 VSUBS 0.03088f
C98 VDD1.n67 VSUBS 0.013833f
C99 VDD1.n68 VSUBS 0.024313f
C100 VDD1.n69 VSUBS 0.013065f
C101 VDD1.n70 VSUBS 0.02316f
C102 VDD1.n71 VSUBS 0.02323f
C103 VDD1.t2 VSUBS 0.066389f
C104 VDD1.n72 VSUBS 0.168846f
C105 VDD1.n73 VSUBS 0.975096f
C106 VDD1.n74 VSUBS 0.013065f
C107 VDD1.n75 VSUBS 0.013833f
C108 VDD1.n76 VSUBS 0.03088f
C109 VDD1.n77 VSUBS 0.03088f
C110 VDD1.n78 VSUBS 0.013833f
C111 VDD1.n79 VSUBS 0.013065f
C112 VDD1.n80 VSUBS 0.024313f
C113 VDD1.n81 VSUBS 0.024313f
C114 VDD1.n82 VSUBS 0.013065f
C115 VDD1.n83 VSUBS 0.013833f
C116 VDD1.n84 VSUBS 0.03088f
C117 VDD1.n85 VSUBS 0.03088f
C118 VDD1.n86 VSUBS 0.013833f
C119 VDD1.n87 VSUBS 0.013065f
C120 VDD1.n88 VSUBS 0.024313f
C121 VDD1.n89 VSUBS 0.024313f
C122 VDD1.n90 VSUBS 0.013065f
C123 VDD1.n91 VSUBS 0.013065f
C124 VDD1.n92 VSUBS 0.013833f
C125 VDD1.n93 VSUBS 0.03088f
C126 VDD1.n94 VSUBS 0.03088f
C127 VDD1.n95 VSUBS 0.03088f
C128 VDD1.n96 VSUBS 0.013449f
C129 VDD1.n97 VSUBS 0.013065f
C130 VDD1.n98 VSUBS 0.024313f
C131 VDD1.n99 VSUBS 0.024313f
C132 VDD1.n100 VSUBS 0.013065f
C133 VDD1.n101 VSUBS 0.013833f
C134 VDD1.n102 VSUBS 0.03088f
C135 VDD1.n103 VSUBS 0.069497f
C136 VDD1.n104 VSUBS 0.013833f
C137 VDD1.n105 VSUBS 0.013065f
C138 VDD1.n106 VSUBS 0.055534f
C139 VDD1.n107 VSUBS 0.053771f
C140 VDD1.t4 VSUBS 0.190976f
C141 VDD1.t3 VSUBS 0.190976f
C142 VDD1.n108 VSUBS 1.43899f
C143 VDD1.n109 VSUBS 0.648634f
C144 VDD1.t6 VSUBS 0.190976f
C145 VDD1.t5 VSUBS 0.190976f
C146 VDD1.n110 VSUBS 1.44381f
C147 VDD1.n111 VSUBS 2.07506f
C148 VDD1.t0 VSUBS 0.190976f
C149 VDD1.t8 VSUBS 0.190976f
C150 VDD1.n112 VSUBS 1.43899f
C151 VDD1.n113 VSUBS 2.42868f
C152 VP.n0 VSUBS 0.071551f
C153 VP.t6 VSUBS 1.1592f
C154 VP.n1 VSUBS 0.489917f
C155 VP.n2 VSUBS 0.071551f
C156 VP.n3 VSUBS 0.071551f
C157 VP.t1 VSUBS 1.1592f
C158 VP.t9 VSUBS 1.1592f
C159 VP.n4 VSUBS 0.089313f
C160 VP.t2 VSUBS 1.1592f
C161 VP.n5 VSUBS 0.322547f
C162 VP.t8 VSUBS 1.1592f
C163 VP.t0 VSUBS 1.18487f
C164 VP.n6 VSUBS 0.457158f
C165 VP.n7 VSUBS 0.489241f
C166 VP.n8 VSUBS 0.489917f
C167 VP.n9 VSUBS 0.488264f
C168 VP.n10 VSUBS 0.012168f
C169 VP.n11 VSUBS 0.468493f
C170 VP.n12 VSUBS 2.16638f
C171 VP.n13 VSUBS 2.213f
C172 VP.t7 VSUBS 1.1592f
C173 VP.n14 VSUBS 0.468493f
C174 VP.n15 VSUBS 0.012168f
C175 VP.t5 VSUBS 1.1592f
C176 VP.n16 VSUBS 0.488264f
C177 VP.n17 VSUBS 0.089313f
C178 VP.n18 VSUBS 0.107242f
C179 VP.n19 VSUBS 0.089313f
C180 VP.t3 VSUBS 1.1592f
C181 VP.n20 VSUBS 0.488264f
C182 VP.n21 VSUBS 0.012168f
C183 VP.t4 VSUBS 1.1592f
C184 VP.n22 VSUBS 0.468493f
C185 VP.n23 VSUBS 0.041554f
C186 VTAIL.t12 VSUBS 0.23174f
C187 VTAIL.t17 VSUBS 0.23174f
C188 VTAIL.n0 VSUBS 1.59939f
C189 VTAIL.n1 VSUBS 0.802473f
C190 VTAIL.n2 VSUBS 0.030543f
C191 VTAIL.n3 VSUBS 0.029503f
C192 VTAIL.n4 VSUBS 0.015853f
C193 VTAIL.n5 VSUBS 0.037472f
C194 VTAIL.n6 VSUBS 0.016786f
C195 VTAIL.n7 VSUBS 0.029503f
C196 VTAIL.n8 VSUBS 0.01632f
C197 VTAIL.n9 VSUBS 0.037472f
C198 VTAIL.n10 VSUBS 0.016786f
C199 VTAIL.n11 VSUBS 0.029503f
C200 VTAIL.n12 VSUBS 0.015853f
C201 VTAIL.n13 VSUBS 0.037472f
C202 VTAIL.n14 VSUBS 0.016786f
C203 VTAIL.n15 VSUBS 0.029503f
C204 VTAIL.n16 VSUBS 0.015853f
C205 VTAIL.n17 VSUBS 0.028104f
C206 VTAIL.n18 VSUBS 0.028188f
C207 VTAIL.t2 VSUBS 0.08056f
C208 VTAIL.n19 VSUBS 0.204886f
C209 VTAIL.n20 VSUBS 1.18323f
C210 VTAIL.n21 VSUBS 0.015853f
C211 VTAIL.n22 VSUBS 0.016786f
C212 VTAIL.n23 VSUBS 0.037472f
C213 VTAIL.n24 VSUBS 0.037472f
C214 VTAIL.n25 VSUBS 0.016786f
C215 VTAIL.n26 VSUBS 0.015853f
C216 VTAIL.n27 VSUBS 0.029503f
C217 VTAIL.n28 VSUBS 0.029503f
C218 VTAIL.n29 VSUBS 0.015853f
C219 VTAIL.n30 VSUBS 0.016786f
C220 VTAIL.n31 VSUBS 0.037472f
C221 VTAIL.n32 VSUBS 0.037472f
C222 VTAIL.n33 VSUBS 0.016786f
C223 VTAIL.n34 VSUBS 0.015853f
C224 VTAIL.n35 VSUBS 0.029503f
C225 VTAIL.n36 VSUBS 0.029503f
C226 VTAIL.n37 VSUBS 0.015853f
C227 VTAIL.n38 VSUBS 0.015853f
C228 VTAIL.n39 VSUBS 0.016786f
C229 VTAIL.n40 VSUBS 0.037472f
C230 VTAIL.n41 VSUBS 0.037472f
C231 VTAIL.n42 VSUBS 0.037472f
C232 VTAIL.n43 VSUBS 0.01632f
C233 VTAIL.n44 VSUBS 0.015853f
C234 VTAIL.n45 VSUBS 0.029503f
C235 VTAIL.n46 VSUBS 0.029503f
C236 VTAIL.n47 VSUBS 0.015853f
C237 VTAIL.n48 VSUBS 0.016786f
C238 VTAIL.n49 VSUBS 0.037472f
C239 VTAIL.n50 VSUBS 0.084331f
C240 VTAIL.n51 VSUBS 0.016786f
C241 VTAIL.n52 VSUBS 0.015853f
C242 VTAIL.n53 VSUBS 0.067388f
C243 VTAIL.n54 VSUBS 0.042101f
C244 VTAIL.n55 VSUBS 0.203397f
C245 VTAIL.t5 VSUBS 0.23174f
C246 VTAIL.t6 VSUBS 0.23174f
C247 VTAIL.n56 VSUBS 1.59939f
C248 VTAIL.n57 VSUBS 0.819273f
C249 VTAIL.t1 VSUBS 0.23174f
C250 VTAIL.t3 VSUBS 0.23174f
C251 VTAIL.n58 VSUBS 1.59939f
C252 VTAIL.n59 VSUBS 2.12396f
C253 VTAIL.t11 VSUBS 0.23174f
C254 VTAIL.t19 VSUBS 0.23174f
C255 VTAIL.n60 VSUBS 1.5994f
C256 VTAIL.n61 VSUBS 2.12395f
C257 VTAIL.t13 VSUBS 0.23174f
C258 VTAIL.t10 VSUBS 0.23174f
C259 VTAIL.n62 VSUBS 1.5994f
C260 VTAIL.n63 VSUBS 0.819262f
C261 VTAIL.n64 VSUBS 0.030543f
C262 VTAIL.n65 VSUBS 0.029503f
C263 VTAIL.n66 VSUBS 0.015853f
C264 VTAIL.n67 VSUBS 0.037472f
C265 VTAIL.n68 VSUBS 0.016786f
C266 VTAIL.n69 VSUBS 0.029503f
C267 VTAIL.n70 VSUBS 0.01632f
C268 VTAIL.n71 VSUBS 0.037472f
C269 VTAIL.n72 VSUBS 0.015853f
C270 VTAIL.n73 VSUBS 0.016786f
C271 VTAIL.n74 VSUBS 0.029503f
C272 VTAIL.n75 VSUBS 0.015853f
C273 VTAIL.n76 VSUBS 0.037472f
C274 VTAIL.n77 VSUBS 0.016786f
C275 VTAIL.n78 VSUBS 0.029503f
C276 VTAIL.n79 VSUBS 0.015853f
C277 VTAIL.n80 VSUBS 0.028104f
C278 VTAIL.n81 VSUBS 0.028188f
C279 VTAIL.t14 VSUBS 0.08056f
C280 VTAIL.n82 VSUBS 0.204886f
C281 VTAIL.n83 VSUBS 1.18323f
C282 VTAIL.n84 VSUBS 0.015853f
C283 VTAIL.n85 VSUBS 0.016786f
C284 VTAIL.n86 VSUBS 0.037472f
C285 VTAIL.n87 VSUBS 0.037472f
C286 VTAIL.n88 VSUBS 0.016786f
C287 VTAIL.n89 VSUBS 0.015853f
C288 VTAIL.n90 VSUBS 0.029503f
C289 VTAIL.n91 VSUBS 0.029503f
C290 VTAIL.n92 VSUBS 0.015853f
C291 VTAIL.n93 VSUBS 0.016786f
C292 VTAIL.n94 VSUBS 0.037472f
C293 VTAIL.n95 VSUBS 0.037472f
C294 VTAIL.n96 VSUBS 0.016786f
C295 VTAIL.n97 VSUBS 0.015853f
C296 VTAIL.n98 VSUBS 0.029503f
C297 VTAIL.n99 VSUBS 0.029503f
C298 VTAIL.n100 VSUBS 0.015853f
C299 VTAIL.n101 VSUBS 0.016786f
C300 VTAIL.n102 VSUBS 0.037472f
C301 VTAIL.n103 VSUBS 0.037472f
C302 VTAIL.n104 VSUBS 0.037472f
C303 VTAIL.n105 VSUBS 0.01632f
C304 VTAIL.n106 VSUBS 0.015853f
C305 VTAIL.n107 VSUBS 0.029503f
C306 VTAIL.n108 VSUBS 0.029503f
C307 VTAIL.n109 VSUBS 0.015853f
C308 VTAIL.n110 VSUBS 0.016786f
C309 VTAIL.n111 VSUBS 0.037472f
C310 VTAIL.n112 VSUBS 0.084331f
C311 VTAIL.n113 VSUBS 0.016786f
C312 VTAIL.n114 VSUBS 0.015853f
C313 VTAIL.n115 VSUBS 0.067388f
C314 VTAIL.n116 VSUBS 0.042101f
C315 VTAIL.n117 VSUBS 0.203397f
C316 VTAIL.t8 VSUBS 0.23174f
C317 VTAIL.t7 VSUBS 0.23174f
C318 VTAIL.n118 VSUBS 1.5994f
C319 VTAIL.n119 VSUBS 0.819262f
C320 VTAIL.t0 VSUBS 0.23174f
C321 VTAIL.t4 VSUBS 0.23174f
C322 VTAIL.n120 VSUBS 1.5994f
C323 VTAIL.n121 VSUBS 0.819262f
C324 VTAIL.n122 VSUBS 0.030543f
C325 VTAIL.n123 VSUBS 0.029503f
C326 VTAIL.n124 VSUBS 0.015853f
C327 VTAIL.n125 VSUBS 0.037472f
C328 VTAIL.n126 VSUBS 0.016786f
C329 VTAIL.n127 VSUBS 0.029503f
C330 VTAIL.n128 VSUBS 0.01632f
C331 VTAIL.n129 VSUBS 0.037472f
C332 VTAIL.n130 VSUBS 0.015853f
C333 VTAIL.n131 VSUBS 0.016786f
C334 VTAIL.n132 VSUBS 0.029503f
C335 VTAIL.n133 VSUBS 0.015853f
C336 VTAIL.n134 VSUBS 0.037472f
C337 VTAIL.n135 VSUBS 0.016786f
C338 VTAIL.n136 VSUBS 0.029503f
C339 VTAIL.n137 VSUBS 0.015853f
C340 VTAIL.n138 VSUBS 0.028104f
C341 VTAIL.n139 VSUBS 0.028188f
C342 VTAIL.t9 VSUBS 0.08056f
C343 VTAIL.n140 VSUBS 0.204886f
C344 VTAIL.n141 VSUBS 1.18323f
C345 VTAIL.n142 VSUBS 0.015853f
C346 VTAIL.n143 VSUBS 0.016786f
C347 VTAIL.n144 VSUBS 0.037472f
C348 VTAIL.n145 VSUBS 0.037472f
C349 VTAIL.n146 VSUBS 0.016786f
C350 VTAIL.n147 VSUBS 0.015853f
C351 VTAIL.n148 VSUBS 0.029503f
C352 VTAIL.n149 VSUBS 0.029503f
C353 VTAIL.n150 VSUBS 0.015853f
C354 VTAIL.n151 VSUBS 0.016786f
C355 VTAIL.n152 VSUBS 0.037472f
C356 VTAIL.n153 VSUBS 0.037472f
C357 VTAIL.n154 VSUBS 0.016786f
C358 VTAIL.n155 VSUBS 0.015853f
C359 VTAIL.n156 VSUBS 0.029503f
C360 VTAIL.n157 VSUBS 0.029503f
C361 VTAIL.n158 VSUBS 0.015853f
C362 VTAIL.n159 VSUBS 0.016786f
C363 VTAIL.n160 VSUBS 0.037472f
C364 VTAIL.n161 VSUBS 0.037472f
C365 VTAIL.n162 VSUBS 0.037472f
C366 VTAIL.n163 VSUBS 0.01632f
C367 VTAIL.n164 VSUBS 0.015853f
C368 VTAIL.n165 VSUBS 0.029503f
C369 VTAIL.n166 VSUBS 0.029503f
C370 VTAIL.n167 VSUBS 0.015853f
C371 VTAIL.n168 VSUBS 0.016786f
C372 VTAIL.n169 VSUBS 0.037472f
C373 VTAIL.n170 VSUBS 0.084331f
C374 VTAIL.n171 VSUBS 0.016786f
C375 VTAIL.n172 VSUBS 0.015853f
C376 VTAIL.n173 VSUBS 0.067388f
C377 VTAIL.n174 VSUBS 0.042101f
C378 VTAIL.n175 VSUBS 1.41876f
C379 VTAIL.n176 VSUBS 0.030543f
C380 VTAIL.n177 VSUBS 0.029503f
C381 VTAIL.n178 VSUBS 0.015853f
C382 VTAIL.n179 VSUBS 0.037472f
C383 VTAIL.n180 VSUBS 0.016786f
C384 VTAIL.n181 VSUBS 0.029503f
C385 VTAIL.n182 VSUBS 0.01632f
C386 VTAIL.n183 VSUBS 0.037472f
C387 VTAIL.n184 VSUBS 0.016786f
C388 VTAIL.n185 VSUBS 0.029503f
C389 VTAIL.n186 VSUBS 0.015853f
C390 VTAIL.n187 VSUBS 0.037472f
C391 VTAIL.n188 VSUBS 0.016786f
C392 VTAIL.n189 VSUBS 0.029503f
C393 VTAIL.n190 VSUBS 0.015853f
C394 VTAIL.n191 VSUBS 0.028104f
C395 VTAIL.n192 VSUBS 0.028188f
C396 VTAIL.t18 VSUBS 0.08056f
C397 VTAIL.n193 VSUBS 0.204886f
C398 VTAIL.n194 VSUBS 1.18323f
C399 VTAIL.n195 VSUBS 0.015853f
C400 VTAIL.n196 VSUBS 0.016786f
C401 VTAIL.n197 VSUBS 0.037472f
C402 VTAIL.n198 VSUBS 0.037472f
C403 VTAIL.n199 VSUBS 0.016786f
C404 VTAIL.n200 VSUBS 0.015853f
C405 VTAIL.n201 VSUBS 0.029503f
C406 VTAIL.n202 VSUBS 0.029503f
C407 VTAIL.n203 VSUBS 0.015853f
C408 VTAIL.n204 VSUBS 0.016786f
C409 VTAIL.n205 VSUBS 0.037472f
C410 VTAIL.n206 VSUBS 0.037472f
C411 VTAIL.n207 VSUBS 0.016786f
C412 VTAIL.n208 VSUBS 0.015853f
C413 VTAIL.n209 VSUBS 0.029503f
C414 VTAIL.n210 VSUBS 0.029503f
C415 VTAIL.n211 VSUBS 0.015853f
C416 VTAIL.n212 VSUBS 0.015853f
C417 VTAIL.n213 VSUBS 0.016786f
C418 VTAIL.n214 VSUBS 0.037472f
C419 VTAIL.n215 VSUBS 0.037472f
C420 VTAIL.n216 VSUBS 0.037472f
C421 VTAIL.n217 VSUBS 0.01632f
C422 VTAIL.n218 VSUBS 0.015853f
C423 VTAIL.n219 VSUBS 0.029503f
C424 VTAIL.n220 VSUBS 0.029503f
C425 VTAIL.n221 VSUBS 0.015853f
C426 VTAIL.n222 VSUBS 0.016786f
C427 VTAIL.n223 VSUBS 0.037472f
C428 VTAIL.n224 VSUBS 0.084331f
C429 VTAIL.n225 VSUBS 0.016786f
C430 VTAIL.n226 VSUBS 0.015853f
C431 VTAIL.n227 VSUBS 0.067388f
C432 VTAIL.n228 VSUBS 0.042101f
C433 VTAIL.n229 VSUBS 1.41876f
C434 VTAIL.t15 VSUBS 0.23174f
C435 VTAIL.t16 VSUBS 0.23174f
C436 VTAIL.n230 VSUBS 1.59939f
C437 VTAIL.n231 VSUBS 0.746746f
C438 VDD2.n0 VSUBS 0.025014f
C439 VDD2.n1 VSUBS 0.024163f
C440 VDD2.n2 VSUBS 0.012984f
C441 VDD2.n3 VSUBS 0.030689f
C442 VDD2.n4 VSUBS 0.013748f
C443 VDD2.n5 VSUBS 0.024163f
C444 VDD2.n6 VSUBS 0.013366f
C445 VDD2.n7 VSUBS 0.030689f
C446 VDD2.n8 VSUBS 0.013748f
C447 VDD2.n9 VSUBS 0.024163f
C448 VDD2.n10 VSUBS 0.012984f
C449 VDD2.n11 VSUBS 0.030689f
C450 VDD2.n12 VSUBS 0.013748f
C451 VDD2.n13 VSUBS 0.024163f
C452 VDD2.n14 VSUBS 0.012984f
C453 VDD2.n15 VSUBS 0.023017f
C454 VDD2.n16 VSUBS 0.023086f
C455 VDD2.t1 VSUBS 0.065979f
C456 VDD2.n17 VSUBS 0.167801f
C457 VDD2.n18 VSUBS 0.969062f
C458 VDD2.n19 VSUBS 0.012984f
C459 VDD2.n20 VSUBS 0.013748f
C460 VDD2.n21 VSUBS 0.030689f
C461 VDD2.n22 VSUBS 0.030689f
C462 VDD2.n23 VSUBS 0.013748f
C463 VDD2.n24 VSUBS 0.012984f
C464 VDD2.n25 VSUBS 0.024163f
C465 VDD2.n26 VSUBS 0.024163f
C466 VDD2.n27 VSUBS 0.012984f
C467 VDD2.n28 VSUBS 0.013748f
C468 VDD2.n29 VSUBS 0.030689f
C469 VDD2.n30 VSUBS 0.030689f
C470 VDD2.n31 VSUBS 0.013748f
C471 VDD2.n32 VSUBS 0.012984f
C472 VDD2.n33 VSUBS 0.024163f
C473 VDD2.n34 VSUBS 0.024163f
C474 VDD2.n35 VSUBS 0.012984f
C475 VDD2.n36 VSUBS 0.012984f
C476 VDD2.n37 VSUBS 0.013748f
C477 VDD2.n38 VSUBS 0.030689f
C478 VDD2.n39 VSUBS 0.030689f
C479 VDD2.n40 VSUBS 0.030689f
C480 VDD2.n41 VSUBS 0.013366f
C481 VDD2.n42 VSUBS 0.012984f
C482 VDD2.n43 VSUBS 0.024163f
C483 VDD2.n44 VSUBS 0.024163f
C484 VDD2.n45 VSUBS 0.012984f
C485 VDD2.n46 VSUBS 0.013748f
C486 VDD2.n47 VSUBS 0.030689f
C487 VDD2.n48 VSUBS 0.069067f
C488 VDD2.n49 VSUBS 0.013748f
C489 VDD2.n50 VSUBS 0.012984f
C490 VDD2.n51 VSUBS 0.05519f
C491 VDD2.n52 VSUBS 0.053438f
C492 VDD2.t8 VSUBS 0.189794f
C493 VDD2.t2 VSUBS 0.189794f
C494 VDD2.n53 VSUBS 1.43008f
C495 VDD2.n54 VSUBS 0.644621f
C496 VDD2.t6 VSUBS 0.189794f
C497 VDD2.t9 VSUBS 0.189794f
C498 VDD2.n55 VSUBS 1.43488f
C499 VDD2.n56 VSUBS 1.98716f
C500 VDD2.n57 VSUBS 0.025014f
C501 VDD2.n58 VSUBS 0.024163f
C502 VDD2.n59 VSUBS 0.012984f
C503 VDD2.n60 VSUBS 0.030689f
C504 VDD2.n61 VSUBS 0.013748f
C505 VDD2.n62 VSUBS 0.024163f
C506 VDD2.n63 VSUBS 0.013366f
C507 VDD2.n64 VSUBS 0.030689f
C508 VDD2.n65 VSUBS 0.012984f
C509 VDD2.n66 VSUBS 0.013748f
C510 VDD2.n67 VSUBS 0.024163f
C511 VDD2.n68 VSUBS 0.012984f
C512 VDD2.n69 VSUBS 0.030689f
C513 VDD2.n70 VSUBS 0.013748f
C514 VDD2.n71 VSUBS 0.024163f
C515 VDD2.n72 VSUBS 0.012984f
C516 VDD2.n73 VSUBS 0.023017f
C517 VDD2.n74 VSUBS 0.023086f
C518 VDD2.t0 VSUBS 0.065979f
C519 VDD2.n75 VSUBS 0.167801f
C520 VDD2.n76 VSUBS 0.969062f
C521 VDD2.n77 VSUBS 0.012984f
C522 VDD2.n78 VSUBS 0.013748f
C523 VDD2.n79 VSUBS 0.030689f
C524 VDD2.n80 VSUBS 0.030689f
C525 VDD2.n81 VSUBS 0.013748f
C526 VDD2.n82 VSUBS 0.012984f
C527 VDD2.n83 VSUBS 0.024163f
C528 VDD2.n84 VSUBS 0.024163f
C529 VDD2.n85 VSUBS 0.012984f
C530 VDD2.n86 VSUBS 0.013748f
C531 VDD2.n87 VSUBS 0.030689f
C532 VDD2.n88 VSUBS 0.030689f
C533 VDD2.n89 VSUBS 0.013748f
C534 VDD2.n90 VSUBS 0.012984f
C535 VDD2.n91 VSUBS 0.024163f
C536 VDD2.n92 VSUBS 0.024163f
C537 VDD2.n93 VSUBS 0.012984f
C538 VDD2.n94 VSUBS 0.013748f
C539 VDD2.n95 VSUBS 0.030689f
C540 VDD2.n96 VSUBS 0.030689f
C541 VDD2.n97 VSUBS 0.030689f
C542 VDD2.n98 VSUBS 0.013366f
C543 VDD2.n99 VSUBS 0.012984f
C544 VDD2.n100 VSUBS 0.024163f
C545 VDD2.n101 VSUBS 0.024163f
C546 VDD2.n102 VSUBS 0.012984f
C547 VDD2.n103 VSUBS 0.013748f
C548 VDD2.n104 VSUBS 0.030689f
C549 VDD2.n105 VSUBS 0.069067f
C550 VDD2.n106 VSUBS 0.013748f
C551 VDD2.n107 VSUBS 0.012984f
C552 VDD2.n108 VSUBS 0.05519f
C553 VDD2.n109 VSUBS 0.05117f
C554 VDD2.n110 VSUBS 1.94823f
C555 VDD2.t4 VSUBS 0.189794f
C556 VDD2.t3 VSUBS 0.189794f
C557 VDD2.n111 VSUBS 1.43009f
C558 VDD2.n112 VSUBS 0.533294f
C559 VDD2.t7 VSUBS 0.189794f
C560 VDD2.t5 VSUBS 0.189794f
C561 VDD2.n113 VSUBS 1.43485f
C562 VN.n0 VSUBS 0.069669f
C563 VN.t4 VSUBS 1.12871f
C564 VN.n1 VSUBS 0.477031f
C565 VN.t7 VSUBS 1.1537f
C566 VN.t2 VSUBS 1.12871f
C567 VN.n2 VSUBS 0.476373f
C568 VN.n3 VSUBS 0.445134f
C569 VN.n4 VSUBS 0.314064f
C570 VN.n5 VSUBS 0.086964f
C571 VN.t3 VSUBS 1.12871f
C572 VN.n6 VSUBS 0.475422f
C573 VN.n7 VSUBS 0.011848f
C574 VN.t1 VSUBS 1.12871f
C575 VN.n8 VSUBS 0.45617f
C576 VN.n9 VSUBS 0.040461f
C577 VN.n10 VSUBS 0.069669f
C578 VN.t6 VSUBS 1.12871f
C579 VN.n11 VSUBS 0.477031f
C580 VN.t0 VSUBS 1.12871f
C581 VN.t5 VSUBS 1.1537f
C582 VN.t9 VSUBS 1.12871f
C583 VN.n12 VSUBS 0.476373f
C584 VN.n13 VSUBS 0.445134f
C585 VN.n14 VSUBS 0.314064f
C586 VN.n15 VSUBS 0.086964f
C587 VN.n16 VSUBS 0.475422f
C588 VN.n17 VSUBS 0.011848f
C589 VN.t8 VSUBS 1.12871f
C590 VN.n18 VSUBS 0.45617f
C591 VN.n19 VSUBS 2.14371f
C592 B.n0 VSUBS 0.006669f
C593 B.n1 VSUBS 0.006669f
C594 B.n2 VSUBS 0.009864f
C595 B.n3 VSUBS 0.007559f
C596 B.n4 VSUBS 0.007559f
C597 B.n5 VSUBS 0.007559f
C598 B.n6 VSUBS 0.007559f
C599 B.n7 VSUBS 0.007559f
C600 B.n8 VSUBS 0.007559f
C601 B.n9 VSUBS 0.007559f
C602 B.n10 VSUBS 0.007559f
C603 B.n11 VSUBS 0.007559f
C604 B.n12 VSUBS 0.007559f
C605 B.n13 VSUBS 0.007559f
C606 B.n14 VSUBS 0.007559f
C607 B.n15 VSUBS 0.015976f
C608 B.n16 VSUBS 0.007559f
C609 B.n17 VSUBS 0.007559f
C610 B.n18 VSUBS 0.007559f
C611 B.n19 VSUBS 0.007559f
C612 B.n20 VSUBS 0.007559f
C613 B.n21 VSUBS 0.007559f
C614 B.n22 VSUBS 0.007559f
C615 B.n23 VSUBS 0.007559f
C616 B.n24 VSUBS 0.007559f
C617 B.n25 VSUBS 0.007559f
C618 B.n26 VSUBS 0.007559f
C619 B.n27 VSUBS 0.007559f
C620 B.n28 VSUBS 0.007559f
C621 B.n29 VSUBS 0.007559f
C622 B.n30 VSUBS 0.007559f
C623 B.n31 VSUBS 0.007559f
C624 B.n32 VSUBS 0.007559f
C625 B.n33 VSUBS 0.007559f
C626 B.t10 VSUBS 0.179377f
C627 B.t11 VSUBS 0.19237f
C628 B.t9 VSUBS 0.342613f
C629 B.n34 VSUBS 0.290651f
C630 B.n35 VSUBS 0.231765f
C631 B.n36 VSUBS 0.007559f
C632 B.n37 VSUBS 0.007559f
C633 B.n38 VSUBS 0.007559f
C634 B.n39 VSUBS 0.007559f
C635 B.t4 VSUBS 0.17938f
C636 B.t5 VSUBS 0.192373f
C637 B.t3 VSUBS 0.342613f
C638 B.n40 VSUBS 0.290649f
C639 B.n41 VSUBS 0.231762f
C640 B.n42 VSUBS 0.017513f
C641 B.n43 VSUBS 0.007559f
C642 B.n44 VSUBS 0.007559f
C643 B.n45 VSUBS 0.007559f
C644 B.n46 VSUBS 0.007559f
C645 B.n47 VSUBS 0.007559f
C646 B.n48 VSUBS 0.007559f
C647 B.n49 VSUBS 0.007559f
C648 B.n50 VSUBS 0.007559f
C649 B.n51 VSUBS 0.007559f
C650 B.n52 VSUBS 0.007559f
C651 B.n53 VSUBS 0.007559f
C652 B.n54 VSUBS 0.007559f
C653 B.n55 VSUBS 0.007559f
C654 B.n56 VSUBS 0.007559f
C655 B.n57 VSUBS 0.007559f
C656 B.n58 VSUBS 0.007559f
C657 B.n59 VSUBS 0.007559f
C658 B.n60 VSUBS 0.016926f
C659 B.n61 VSUBS 0.007559f
C660 B.n62 VSUBS 0.007559f
C661 B.n63 VSUBS 0.007559f
C662 B.n64 VSUBS 0.007559f
C663 B.n65 VSUBS 0.007559f
C664 B.n66 VSUBS 0.007559f
C665 B.n67 VSUBS 0.007559f
C666 B.n68 VSUBS 0.007559f
C667 B.n69 VSUBS 0.007559f
C668 B.n70 VSUBS 0.007559f
C669 B.n71 VSUBS 0.007559f
C670 B.n72 VSUBS 0.007559f
C671 B.n73 VSUBS 0.007559f
C672 B.n74 VSUBS 0.007559f
C673 B.n75 VSUBS 0.007559f
C674 B.n76 VSUBS 0.007559f
C675 B.n77 VSUBS 0.007559f
C676 B.n78 VSUBS 0.007559f
C677 B.n79 VSUBS 0.007559f
C678 B.n80 VSUBS 0.007559f
C679 B.n81 VSUBS 0.007559f
C680 B.n82 VSUBS 0.007559f
C681 B.n83 VSUBS 0.007559f
C682 B.n84 VSUBS 0.007559f
C683 B.n85 VSUBS 0.007559f
C684 B.n86 VSUBS 0.007559f
C685 B.n87 VSUBS 0.007559f
C686 B.n88 VSUBS 0.016975f
C687 B.n89 VSUBS 0.007559f
C688 B.n90 VSUBS 0.007559f
C689 B.n91 VSUBS 0.007559f
C690 B.n92 VSUBS 0.007559f
C691 B.n93 VSUBS 0.007559f
C692 B.n94 VSUBS 0.007559f
C693 B.n95 VSUBS 0.007559f
C694 B.n96 VSUBS 0.007559f
C695 B.n97 VSUBS 0.007559f
C696 B.n98 VSUBS 0.007559f
C697 B.n99 VSUBS 0.007559f
C698 B.n100 VSUBS 0.007559f
C699 B.n101 VSUBS 0.007559f
C700 B.n102 VSUBS 0.007559f
C701 B.n103 VSUBS 0.007559f
C702 B.n104 VSUBS 0.007559f
C703 B.n105 VSUBS 0.007559f
C704 B.n106 VSUBS 0.005224f
C705 B.n107 VSUBS 0.007559f
C706 B.n108 VSUBS 0.007559f
C707 B.n109 VSUBS 0.007559f
C708 B.n110 VSUBS 0.007559f
C709 B.n111 VSUBS 0.007559f
C710 B.t2 VSUBS 0.179377f
C711 B.t1 VSUBS 0.19237f
C712 B.t0 VSUBS 0.342613f
C713 B.n112 VSUBS 0.290651f
C714 B.n113 VSUBS 0.231765f
C715 B.n114 VSUBS 0.007559f
C716 B.n115 VSUBS 0.007559f
C717 B.n116 VSUBS 0.007559f
C718 B.n117 VSUBS 0.007559f
C719 B.n118 VSUBS 0.007559f
C720 B.n119 VSUBS 0.007559f
C721 B.n120 VSUBS 0.007559f
C722 B.n121 VSUBS 0.007559f
C723 B.n122 VSUBS 0.007559f
C724 B.n123 VSUBS 0.007559f
C725 B.n124 VSUBS 0.007559f
C726 B.n125 VSUBS 0.007559f
C727 B.n126 VSUBS 0.007559f
C728 B.n127 VSUBS 0.007559f
C729 B.n128 VSUBS 0.007559f
C730 B.n129 VSUBS 0.007559f
C731 B.n130 VSUBS 0.007559f
C732 B.n131 VSUBS 0.015976f
C733 B.n132 VSUBS 0.007559f
C734 B.n133 VSUBS 0.007559f
C735 B.n134 VSUBS 0.007559f
C736 B.n135 VSUBS 0.007559f
C737 B.n136 VSUBS 0.007559f
C738 B.n137 VSUBS 0.007559f
C739 B.n138 VSUBS 0.007559f
C740 B.n139 VSUBS 0.007559f
C741 B.n140 VSUBS 0.007559f
C742 B.n141 VSUBS 0.007559f
C743 B.n142 VSUBS 0.007559f
C744 B.n143 VSUBS 0.007559f
C745 B.n144 VSUBS 0.007559f
C746 B.n145 VSUBS 0.007559f
C747 B.n146 VSUBS 0.007559f
C748 B.n147 VSUBS 0.007559f
C749 B.n148 VSUBS 0.007559f
C750 B.n149 VSUBS 0.007559f
C751 B.n150 VSUBS 0.007559f
C752 B.n151 VSUBS 0.007559f
C753 B.n152 VSUBS 0.007559f
C754 B.n153 VSUBS 0.007559f
C755 B.n154 VSUBS 0.007559f
C756 B.n155 VSUBS 0.007559f
C757 B.n156 VSUBS 0.007559f
C758 B.n157 VSUBS 0.007559f
C759 B.n158 VSUBS 0.007559f
C760 B.n159 VSUBS 0.007559f
C761 B.n160 VSUBS 0.007559f
C762 B.n161 VSUBS 0.007559f
C763 B.n162 VSUBS 0.007559f
C764 B.n163 VSUBS 0.007559f
C765 B.n164 VSUBS 0.007559f
C766 B.n165 VSUBS 0.007559f
C767 B.n166 VSUBS 0.007559f
C768 B.n167 VSUBS 0.007559f
C769 B.n168 VSUBS 0.007559f
C770 B.n169 VSUBS 0.007559f
C771 B.n170 VSUBS 0.007559f
C772 B.n171 VSUBS 0.007559f
C773 B.n172 VSUBS 0.007559f
C774 B.n173 VSUBS 0.007559f
C775 B.n174 VSUBS 0.007559f
C776 B.n175 VSUBS 0.007559f
C777 B.n176 VSUBS 0.007559f
C778 B.n177 VSUBS 0.007559f
C779 B.n178 VSUBS 0.007559f
C780 B.n179 VSUBS 0.007559f
C781 B.n180 VSUBS 0.007559f
C782 B.n181 VSUBS 0.007559f
C783 B.n182 VSUBS 0.015976f
C784 B.n183 VSUBS 0.016926f
C785 B.n184 VSUBS 0.016926f
C786 B.n185 VSUBS 0.007559f
C787 B.n186 VSUBS 0.007559f
C788 B.n187 VSUBS 0.007559f
C789 B.n188 VSUBS 0.007559f
C790 B.n189 VSUBS 0.007559f
C791 B.n190 VSUBS 0.007559f
C792 B.n191 VSUBS 0.007559f
C793 B.n192 VSUBS 0.007559f
C794 B.n193 VSUBS 0.007559f
C795 B.n194 VSUBS 0.007559f
C796 B.n195 VSUBS 0.007559f
C797 B.n196 VSUBS 0.007559f
C798 B.n197 VSUBS 0.007559f
C799 B.n198 VSUBS 0.007559f
C800 B.n199 VSUBS 0.007559f
C801 B.n200 VSUBS 0.007559f
C802 B.n201 VSUBS 0.007559f
C803 B.n202 VSUBS 0.007559f
C804 B.n203 VSUBS 0.007559f
C805 B.n204 VSUBS 0.007559f
C806 B.n205 VSUBS 0.007559f
C807 B.n206 VSUBS 0.007559f
C808 B.n207 VSUBS 0.007559f
C809 B.n208 VSUBS 0.007559f
C810 B.n209 VSUBS 0.007559f
C811 B.n210 VSUBS 0.007559f
C812 B.n211 VSUBS 0.007559f
C813 B.n212 VSUBS 0.007559f
C814 B.n213 VSUBS 0.007559f
C815 B.n214 VSUBS 0.007559f
C816 B.n215 VSUBS 0.007559f
C817 B.n216 VSUBS 0.007559f
C818 B.n217 VSUBS 0.007559f
C819 B.n218 VSUBS 0.007559f
C820 B.n219 VSUBS 0.007559f
C821 B.n220 VSUBS 0.007559f
C822 B.n221 VSUBS 0.007559f
C823 B.n222 VSUBS 0.007559f
C824 B.n223 VSUBS 0.007559f
C825 B.n224 VSUBS 0.007559f
C826 B.n225 VSUBS 0.007559f
C827 B.n226 VSUBS 0.007559f
C828 B.n227 VSUBS 0.007559f
C829 B.n228 VSUBS 0.007559f
C830 B.n229 VSUBS 0.007559f
C831 B.n230 VSUBS 0.007559f
C832 B.n231 VSUBS 0.007559f
C833 B.n232 VSUBS 0.007559f
C834 B.n233 VSUBS 0.007559f
C835 B.n234 VSUBS 0.007559f
C836 B.n235 VSUBS 0.007559f
C837 B.n236 VSUBS 0.005224f
C838 B.n237 VSUBS 0.017513f
C839 B.n238 VSUBS 0.006114f
C840 B.n239 VSUBS 0.007559f
C841 B.n240 VSUBS 0.007559f
C842 B.n241 VSUBS 0.007559f
C843 B.n242 VSUBS 0.007559f
C844 B.n243 VSUBS 0.007559f
C845 B.n244 VSUBS 0.007559f
C846 B.n245 VSUBS 0.007559f
C847 B.n246 VSUBS 0.007559f
C848 B.n247 VSUBS 0.007559f
C849 B.n248 VSUBS 0.007559f
C850 B.n249 VSUBS 0.007559f
C851 B.t8 VSUBS 0.17938f
C852 B.t7 VSUBS 0.192373f
C853 B.t6 VSUBS 0.342613f
C854 B.n250 VSUBS 0.290649f
C855 B.n251 VSUBS 0.231762f
C856 B.n252 VSUBS 0.017513f
C857 B.n253 VSUBS 0.006114f
C858 B.n254 VSUBS 0.007559f
C859 B.n255 VSUBS 0.007559f
C860 B.n256 VSUBS 0.007559f
C861 B.n257 VSUBS 0.007559f
C862 B.n258 VSUBS 0.007559f
C863 B.n259 VSUBS 0.007559f
C864 B.n260 VSUBS 0.007559f
C865 B.n261 VSUBS 0.007559f
C866 B.n262 VSUBS 0.007559f
C867 B.n263 VSUBS 0.007559f
C868 B.n264 VSUBS 0.007559f
C869 B.n265 VSUBS 0.007559f
C870 B.n266 VSUBS 0.007559f
C871 B.n267 VSUBS 0.007559f
C872 B.n268 VSUBS 0.007559f
C873 B.n269 VSUBS 0.007559f
C874 B.n270 VSUBS 0.007559f
C875 B.n271 VSUBS 0.007559f
C876 B.n272 VSUBS 0.007559f
C877 B.n273 VSUBS 0.007559f
C878 B.n274 VSUBS 0.007559f
C879 B.n275 VSUBS 0.007559f
C880 B.n276 VSUBS 0.007559f
C881 B.n277 VSUBS 0.007559f
C882 B.n278 VSUBS 0.007559f
C883 B.n279 VSUBS 0.007559f
C884 B.n280 VSUBS 0.007559f
C885 B.n281 VSUBS 0.007559f
C886 B.n282 VSUBS 0.007559f
C887 B.n283 VSUBS 0.007559f
C888 B.n284 VSUBS 0.007559f
C889 B.n285 VSUBS 0.007559f
C890 B.n286 VSUBS 0.007559f
C891 B.n287 VSUBS 0.007559f
C892 B.n288 VSUBS 0.007559f
C893 B.n289 VSUBS 0.007559f
C894 B.n290 VSUBS 0.007559f
C895 B.n291 VSUBS 0.007559f
C896 B.n292 VSUBS 0.007559f
C897 B.n293 VSUBS 0.007559f
C898 B.n294 VSUBS 0.007559f
C899 B.n295 VSUBS 0.007559f
C900 B.n296 VSUBS 0.007559f
C901 B.n297 VSUBS 0.007559f
C902 B.n298 VSUBS 0.007559f
C903 B.n299 VSUBS 0.007559f
C904 B.n300 VSUBS 0.007559f
C905 B.n301 VSUBS 0.007559f
C906 B.n302 VSUBS 0.007559f
C907 B.n303 VSUBS 0.007559f
C908 B.n304 VSUBS 0.007559f
C909 B.n305 VSUBS 0.007559f
C910 B.n306 VSUBS 0.007559f
C911 B.n307 VSUBS 0.015927f
C912 B.n308 VSUBS 0.016926f
C913 B.n309 VSUBS 0.015976f
C914 B.n310 VSUBS 0.007559f
C915 B.n311 VSUBS 0.007559f
C916 B.n312 VSUBS 0.007559f
C917 B.n313 VSUBS 0.007559f
C918 B.n314 VSUBS 0.007559f
C919 B.n315 VSUBS 0.007559f
C920 B.n316 VSUBS 0.007559f
C921 B.n317 VSUBS 0.007559f
C922 B.n318 VSUBS 0.007559f
C923 B.n319 VSUBS 0.007559f
C924 B.n320 VSUBS 0.007559f
C925 B.n321 VSUBS 0.007559f
C926 B.n322 VSUBS 0.007559f
C927 B.n323 VSUBS 0.007559f
C928 B.n324 VSUBS 0.007559f
C929 B.n325 VSUBS 0.007559f
C930 B.n326 VSUBS 0.007559f
C931 B.n327 VSUBS 0.007559f
C932 B.n328 VSUBS 0.007559f
C933 B.n329 VSUBS 0.007559f
C934 B.n330 VSUBS 0.007559f
C935 B.n331 VSUBS 0.007559f
C936 B.n332 VSUBS 0.007559f
C937 B.n333 VSUBS 0.007559f
C938 B.n334 VSUBS 0.007559f
C939 B.n335 VSUBS 0.007559f
C940 B.n336 VSUBS 0.007559f
C941 B.n337 VSUBS 0.007559f
C942 B.n338 VSUBS 0.007559f
C943 B.n339 VSUBS 0.007559f
C944 B.n340 VSUBS 0.007559f
C945 B.n341 VSUBS 0.007559f
C946 B.n342 VSUBS 0.007559f
C947 B.n343 VSUBS 0.007559f
C948 B.n344 VSUBS 0.007559f
C949 B.n345 VSUBS 0.007559f
C950 B.n346 VSUBS 0.007559f
C951 B.n347 VSUBS 0.007559f
C952 B.n348 VSUBS 0.007559f
C953 B.n349 VSUBS 0.007559f
C954 B.n350 VSUBS 0.007559f
C955 B.n351 VSUBS 0.007559f
C956 B.n352 VSUBS 0.007559f
C957 B.n353 VSUBS 0.007559f
C958 B.n354 VSUBS 0.007559f
C959 B.n355 VSUBS 0.007559f
C960 B.n356 VSUBS 0.007559f
C961 B.n357 VSUBS 0.007559f
C962 B.n358 VSUBS 0.007559f
C963 B.n359 VSUBS 0.007559f
C964 B.n360 VSUBS 0.007559f
C965 B.n361 VSUBS 0.007559f
C966 B.n362 VSUBS 0.007559f
C967 B.n363 VSUBS 0.007559f
C968 B.n364 VSUBS 0.007559f
C969 B.n365 VSUBS 0.007559f
C970 B.n366 VSUBS 0.007559f
C971 B.n367 VSUBS 0.007559f
C972 B.n368 VSUBS 0.007559f
C973 B.n369 VSUBS 0.007559f
C974 B.n370 VSUBS 0.007559f
C975 B.n371 VSUBS 0.007559f
C976 B.n372 VSUBS 0.007559f
C977 B.n373 VSUBS 0.007559f
C978 B.n374 VSUBS 0.007559f
C979 B.n375 VSUBS 0.007559f
C980 B.n376 VSUBS 0.007559f
C981 B.n377 VSUBS 0.007559f
C982 B.n378 VSUBS 0.007559f
C983 B.n379 VSUBS 0.007559f
C984 B.n380 VSUBS 0.007559f
C985 B.n381 VSUBS 0.007559f
C986 B.n382 VSUBS 0.007559f
C987 B.n383 VSUBS 0.007559f
C988 B.n384 VSUBS 0.007559f
C989 B.n385 VSUBS 0.007559f
C990 B.n386 VSUBS 0.007559f
C991 B.n387 VSUBS 0.007559f
C992 B.n388 VSUBS 0.007559f
C993 B.n389 VSUBS 0.007559f
C994 B.n390 VSUBS 0.007559f
C995 B.n391 VSUBS 0.015976f
C996 B.n392 VSUBS 0.015976f
C997 B.n393 VSUBS 0.016926f
C998 B.n394 VSUBS 0.007559f
C999 B.n395 VSUBS 0.007559f
C1000 B.n396 VSUBS 0.007559f
C1001 B.n397 VSUBS 0.007559f
C1002 B.n398 VSUBS 0.007559f
C1003 B.n399 VSUBS 0.007559f
C1004 B.n400 VSUBS 0.007559f
C1005 B.n401 VSUBS 0.007559f
C1006 B.n402 VSUBS 0.007559f
C1007 B.n403 VSUBS 0.007559f
C1008 B.n404 VSUBS 0.007559f
C1009 B.n405 VSUBS 0.007559f
C1010 B.n406 VSUBS 0.007559f
C1011 B.n407 VSUBS 0.007559f
C1012 B.n408 VSUBS 0.007559f
C1013 B.n409 VSUBS 0.007559f
C1014 B.n410 VSUBS 0.007559f
C1015 B.n411 VSUBS 0.007559f
C1016 B.n412 VSUBS 0.007559f
C1017 B.n413 VSUBS 0.007559f
C1018 B.n414 VSUBS 0.007559f
C1019 B.n415 VSUBS 0.007559f
C1020 B.n416 VSUBS 0.007559f
C1021 B.n417 VSUBS 0.007559f
C1022 B.n418 VSUBS 0.007559f
C1023 B.n419 VSUBS 0.007559f
C1024 B.n420 VSUBS 0.007559f
C1025 B.n421 VSUBS 0.007559f
C1026 B.n422 VSUBS 0.007559f
C1027 B.n423 VSUBS 0.007559f
C1028 B.n424 VSUBS 0.007559f
C1029 B.n425 VSUBS 0.007559f
C1030 B.n426 VSUBS 0.007559f
C1031 B.n427 VSUBS 0.007559f
C1032 B.n428 VSUBS 0.007559f
C1033 B.n429 VSUBS 0.007559f
C1034 B.n430 VSUBS 0.007559f
C1035 B.n431 VSUBS 0.007559f
C1036 B.n432 VSUBS 0.007559f
C1037 B.n433 VSUBS 0.007559f
C1038 B.n434 VSUBS 0.007559f
C1039 B.n435 VSUBS 0.007559f
C1040 B.n436 VSUBS 0.007559f
C1041 B.n437 VSUBS 0.007559f
C1042 B.n438 VSUBS 0.007559f
C1043 B.n439 VSUBS 0.007559f
C1044 B.n440 VSUBS 0.007559f
C1045 B.n441 VSUBS 0.007559f
C1046 B.n442 VSUBS 0.007559f
C1047 B.n443 VSUBS 0.007559f
C1048 B.n444 VSUBS 0.007559f
C1049 B.n445 VSUBS 0.005224f
C1050 B.n446 VSUBS 0.007559f
C1051 B.n447 VSUBS 0.007559f
C1052 B.n448 VSUBS 0.006114f
C1053 B.n449 VSUBS 0.007559f
C1054 B.n450 VSUBS 0.007559f
C1055 B.n451 VSUBS 0.007559f
C1056 B.n452 VSUBS 0.007559f
C1057 B.n453 VSUBS 0.007559f
C1058 B.n454 VSUBS 0.007559f
C1059 B.n455 VSUBS 0.007559f
C1060 B.n456 VSUBS 0.007559f
C1061 B.n457 VSUBS 0.007559f
C1062 B.n458 VSUBS 0.007559f
C1063 B.n459 VSUBS 0.007559f
C1064 B.n460 VSUBS 0.006114f
C1065 B.n461 VSUBS 0.017513f
C1066 B.n462 VSUBS 0.005224f
C1067 B.n463 VSUBS 0.007559f
C1068 B.n464 VSUBS 0.007559f
C1069 B.n465 VSUBS 0.007559f
C1070 B.n466 VSUBS 0.007559f
C1071 B.n467 VSUBS 0.007559f
C1072 B.n468 VSUBS 0.007559f
C1073 B.n469 VSUBS 0.007559f
C1074 B.n470 VSUBS 0.007559f
C1075 B.n471 VSUBS 0.007559f
C1076 B.n472 VSUBS 0.007559f
C1077 B.n473 VSUBS 0.007559f
C1078 B.n474 VSUBS 0.007559f
C1079 B.n475 VSUBS 0.007559f
C1080 B.n476 VSUBS 0.007559f
C1081 B.n477 VSUBS 0.007559f
C1082 B.n478 VSUBS 0.007559f
C1083 B.n479 VSUBS 0.007559f
C1084 B.n480 VSUBS 0.007559f
C1085 B.n481 VSUBS 0.007559f
C1086 B.n482 VSUBS 0.007559f
C1087 B.n483 VSUBS 0.007559f
C1088 B.n484 VSUBS 0.007559f
C1089 B.n485 VSUBS 0.007559f
C1090 B.n486 VSUBS 0.007559f
C1091 B.n487 VSUBS 0.007559f
C1092 B.n488 VSUBS 0.007559f
C1093 B.n489 VSUBS 0.007559f
C1094 B.n490 VSUBS 0.007559f
C1095 B.n491 VSUBS 0.007559f
C1096 B.n492 VSUBS 0.007559f
C1097 B.n493 VSUBS 0.007559f
C1098 B.n494 VSUBS 0.007559f
C1099 B.n495 VSUBS 0.007559f
C1100 B.n496 VSUBS 0.007559f
C1101 B.n497 VSUBS 0.007559f
C1102 B.n498 VSUBS 0.007559f
C1103 B.n499 VSUBS 0.007559f
C1104 B.n500 VSUBS 0.007559f
C1105 B.n501 VSUBS 0.007559f
C1106 B.n502 VSUBS 0.007559f
C1107 B.n503 VSUBS 0.007559f
C1108 B.n504 VSUBS 0.007559f
C1109 B.n505 VSUBS 0.007559f
C1110 B.n506 VSUBS 0.007559f
C1111 B.n507 VSUBS 0.007559f
C1112 B.n508 VSUBS 0.007559f
C1113 B.n509 VSUBS 0.007559f
C1114 B.n510 VSUBS 0.007559f
C1115 B.n511 VSUBS 0.007559f
C1116 B.n512 VSUBS 0.007559f
C1117 B.n513 VSUBS 0.007559f
C1118 B.n514 VSUBS 0.016926f
C1119 B.n515 VSUBS 0.016926f
C1120 B.n516 VSUBS 0.015976f
C1121 B.n517 VSUBS 0.007559f
C1122 B.n518 VSUBS 0.007559f
C1123 B.n519 VSUBS 0.007559f
C1124 B.n520 VSUBS 0.007559f
C1125 B.n521 VSUBS 0.007559f
C1126 B.n522 VSUBS 0.007559f
C1127 B.n523 VSUBS 0.007559f
C1128 B.n524 VSUBS 0.007559f
C1129 B.n525 VSUBS 0.007559f
C1130 B.n526 VSUBS 0.007559f
C1131 B.n527 VSUBS 0.007559f
C1132 B.n528 VSUBS 0.007559f
C1133 B.n529 VSUBS 0.007559f
C1134 B.n530 VSUBS 0.007559f
C1135 B.n531 VSUBS 0.007559f
C1136 B.n532 VSUBS 0.007559f
C1137 B.n533 VSUBS 0.007559f
C1138 B.n534 VSUBS 0.007559f
C1139 B.n535 VSUBS 0.007559f
C1140 B.n536 VSUBS 0.007559f
C1141 B.n537 VSUBS 0.007559f
C1142 B.n538 VSUBS 0.007559f
C1143 B.n539 VSUBS 0.007559f
C1144 B.n540 VSUBS 0.007559f
C1145 B.n541 VSUBS 0.007559f
C1146 B.n542 VSUBS 0.007559f
C1147 B.n543 VSUBS 0.007559f
C1148 B.n544 VSUBS 0.007559f
C1149 B.n545 VSUBS 0.007559f
C1150 B.n546 VSUBS 0.007559f
C1151 B.n547 VSUBS 0.007559f
C1152 B.n548 VSUBS 0.007559f
C1153 B.n549 VSUBS 0.007559f
C1154 B.n550 VSUBS 0.007559f
C1155 B.n551 VSUBS 0.007559f
C1156 B.n552 VSUBS 0.007559f
C1157 B.n553 VSUBS 0.007559f
C1158 B.n554 VSUBS 0.007559f
C1159 B.n555 VSUBS 0.009864f
C1160 B.n556 VSUBS 0.010507f
C1161 B.n557 VSUBS 0.020895f
.ends

