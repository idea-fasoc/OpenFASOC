* NGSPICE file created from diff_pair_sample_1057.ext - technology: sky130A

.subckt diff_pair_sample_1057 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1874_n1432# sky130_fd_pr__pfet_01v8 ad=0.9048 pd=5.42 as=0 ps=0 w=2.32 l=0.8
X1 B.t8 B.t6 B.t7 w_n1874_n1432# sky130_fd_pr__pfet_01v8 ad=0.9048 pd=5.42 as=0 ps=0 w=2.32 l=0.8
X2 B.t5 B.t3 B.t4 w_n1874_n1432# sky130_fd_pr__pfet_01v8 ad=0.9048 pd=5.42 as=0 ps=0 w=2.32 l=0.8
X3 VDD2.t5 VN.t0 VTAIL.t11 w_n1874_n1432# sky130_fd_pr__pfet_01v8 ad=0.9048 pd=5.42 as=0.3828 ps=2.65 w=2.32 l=0.8
X4 VDD2.t4 VN.t1 VTAIL.t10 w_n1874_n1432# sky130_fd_pr__pfet_01v8 ad=0.3828 pd=2.65 as=0.9048 ps=5.42 w=2.32 l=0.8
X5 VDD1.t5 VP.t0 VTAIL.t3 w_n1874_n1432# sky130_fd_pr__pfet_01v8 ad=0.3828 pd=2.65 as=0.9048 ps=5.42 w=2.32 l=0.8
X6 VDD2.t3 VN.t2 VTAIL.t9 w_n1874_n1432# sky130_fd_pr__pfet_01v8 ad=0.9048 pd=5.42 as=0.3828 ps=2.65 w=2.32 l=0.8
X7 VDD1.t4 VP.t1 VTAIL.t0 w_n1874_n1432# sky130_fd_pr__pfet_01v8 ad=0.9048 pd=5.42 as=0.3828 ps=2.65 w=2.32 l=0.8
X8 VTAIL.t7 VN.t3 VDD2.t2 w_n1874_n1432# sky130_fd_pr__pfet_01v8 ad=0.3828 pd=2.65 as=0.3828 ps=2.65 w=2.32 l=0.8
X9 VDD2.t1 VN.t4 VTAIL.t6 w_n1874_n1432# sky130_fd_pr__pfet_01v8 ad=0.3828 pd=2.65 as=0.9048 ps=5.42 w=2.32 l=0.8
X10 VTAIL.t8 VN.t5 VDD2.t0 w_n1874_n1432# sky130_fd_pr__pfet_01v8 ad=0.3828 pd=2.65 as=0.3828 ps=2.65 w=2.32 l=0.8
X11 VDD1.t3 VP.t2 VTAIL.t5 w_n1874_n1432# sky130_fd_pr__pfet_01v8 ad=0.3828 pd=2.65 as=0.9048 ps=5.42 w=2.32 l=0.8
X12 VTAIL.t1 VP.t3 VDD1.t2 w_n1874_n1432# sky130_fd_pr__pfet_01v8 ad=0.3828 pd=2.65 as=0.3828 ps=2.65 w=2.32 l=0.8
X13 VTAIL.t2 VP.t4 VDD1.t1 w_n1874_n1432# sky130_fd_pr__pfet_01v8 ad=0.3828 pd=2.65 as=0.3828 ps=2.65 w=2.32 l=0.8
X14 VDD1.t0 VP.t5 VTAIL.t4 w_n1874_n1432# sky130_fd_pr__pfet_01v8 ad=0.9048 pd=5.42 as=0.3828 ps=2.65 w=2.32 l=0.8
X15 B.t2 B.t0 B.t1 w_n1874_n1432# sky130_fd_pr__pfet_01v8 ad=0.9048 pd=5.42 as=0 ps=0 w=2.32 l=0.8
R0 B.n174 B.n57 585
R1 B.n173 B.n172 585
R2 B.n171 B.n58 585
R3 B.n170 B.n169 585
R4 B.n168 B.n59 585
R5 B.n167 B.n166 585
R6 B.n165 B.n60 585
R7 B.n164 B.n163 585
R8 B.n162 B.n61 585
R9 B.n161 B.n160 585
R10 B.n159 B.n62 585
R11 B.n158 B.n157 585
R12 B.n156 B.n63 585
R13 B.n154 B.n153 585
R14 B.n152 B.n66 585
R15 B.n151 B.n150 585
R16 B.n149 B.n67 585
R17 B.n148 B.n147 585
R18 B.n146 B.n68 585
R19 B.n145 B.n144 585
R20 B.n143 B.n69 585
R21 B.n142 B.n141 585
R22 B.n140 B.n70 585
R23 B.n139 B.n138 585
R24 B.n134 B.n71 585
R25 B.n133 B.n132 585
R26 B.n131 B.n72 585
R27 B.n130 B.n129 585
R28 B.n128 B.n73 585
R29 B.n127 B.n126 585
R30 B.n125 B.n74 585
R31 B.n124 B.n123 585
R32 B.n122 B.n75 585
R33 B.n121 B.n120 585
R34 B.n119 B.n76 585
R35 B.n118 B.n117 585
R36 B.n176 B.n175 585
R37 B.n177 B.n56 585
R38 B.n179 B.n178 585
R39 B.n180 B.n55 585
R40 B.n182 B.n181 585
R41 B.n183 B.n54 585
R42 B.n185 B.n184 585
R43 B.n186 B.n53 585
R44 B.n188 B.n187 585
R45 B.n189 B.n52 585
R46 B.n191 B.n190 585
R47 B.n192 B.n51 585
R48 B.n194 B.n193 585
R49 B.n195 B.n50 585
R50 B.n197 B.n196 585
R51 B.n198 B.n49 585
R52 B.n200 B.n199 585
R53 B.n201 B.n48 585
R54 B.n203 B.n202 585
R55 B.n204 B.n47 585
R56 B.n206 B.n205 585
R57 B.n207 B.n46 585
R58 B.n209 B.n208 585
R59 B.n210 B.n45 585
R60 B.n212 B.n211 585
R61 B.n213 B.n44 585
R62 B.n215 B.n214 585
R63 B.n216 B.n43 585
R64 B.n218 B.n217 585
R65 B.n219 B.n42 585
R66 B.n221 B.n220 585
R67 B.n222 B.n41 585
R68 B.n224 B.n223 585
R69 B.n225 B.n40 585
R70 B.n227 B.n226 585
R71 B.n228 B.n39 585
R72 B.n230 B.n229 585
R73 B.n231 B.n38 585
R74 B.n233 B.n232 585
R75 B.n234 B.n37 585
R76 B.n236 B.n235 585
R77 B.n237 B.n36 585
R78 B.n239 B.n238 585
R79 B.n240 B.n35 585
R80 B.n296 B.n295 585
R81 B.n294 B.n13 585
R82 B.n293 B.n292 585
R83 B.n291 B.n14 585
R84 B.n290 B.n289 585
R85 B.n288 B.n15 585
R86 B.n287 B.n286 585
R87 B.n285 B.n16 585
R88 B.n284 B.n283 585
R89 B.n282 B.n17 585
R90 B.n281 B.n280 585
R91 B.n279 B.n18 585
R92 B.n278 B.n277 585
R93 B.n275 B.n19 585
R94 B.n274 B.n273 585
R95 B.n272 B.n22 585
R96 B.n271 B.n270 585
R97 B.n269 B.n23 585
R98 B.n268 B.n267 585
R99 B.n266 B.n24 585
R100 B.n265 B.n264 585
R101 B.n263 B.n25 585
R102 B.n262 B.n261 585
R103 B.n260 B.n259 585
R104 B.n258 B.n29 585
R105 B.n257 B.n256 585
R106 B.n255 B.n30 585
R107 B.n254 B.n253 585
R108 B.n252 B.n31 585
R109 B.n251 B.n250 585
R110 B.n249 B.n32 585
R111 B.n248 B.n247 585
R112 B.n246 B.n33 585
R113 B.n245 B.n244 585
R114 B.n243 B.n34 585
R115 B.n242 B.n241 585
R116 B.n297 B.n12 585
R117 B.n299 B.n298 585
R118 B.n300 B.n11 585
R119 B.n302 B.n301 585
R120 B.n303 B.n10 585
R121 B.n305 B.n304 585
R122 B.n306 B.n9 585
R123 B.n308 B.n307 585
R124 B.n309 B.n8 585
R125 B.n311 B.n310 585
R126 B.n312 B.n7 585
R127 B.n314 B.n313 585
R128 B.n315 B.n6 585
R129 B.n317 B.n316 585
R130 B.n318 B.n5 585
R131 B.n320 B.n319 585
R132 B.n321 B.n4 585
R133 B.n323 B.n322 585
R134 B.n324 B.n3 585
R135 B.n326 B.n325 585
R136 B.n327 B.n0 585
R137 B.n2 B.n1 585
R138 B.n88 B.n87 585
R139 B.n89 B.n86 585
R140 B.n91 B.n90 585
R141 B.n92 B.n85 585
R142 B.n94 B.n93 585
R143 B.n95 B.n84 585
R144 B.n97 B.n96 585
R145 B.n98 B.n83 585
R146 B.n100 B.n99 585
R147 B.n101 B.n82 585
R148 B.n103 B.n102 585
R149 B.n104 B.n81 585
R150 B.n106 B.n105 585
R151 B.n107 B.n80 585
R152 B.n109 B.n108 585
R153 B.n110 B.n79 585
R154 B.n112 B.n111 585
R155 B.n113 B.n78 585
R156 B.n115 B.n114 585
R157 B.n116 B.n77 585
R158 B.n118 B.n77 473.281
R159 B.n176 B.n57 473.281
R160 B.n242 B.n35 473.281
R161 B.n297 B.n296 473.281
R162 B.n135 B.t9 271.779
R163 B.n64 B.t6 271.779
R164 B.n26 B.t0 271.779
R165 B.n20 B.t3 271.779
R166 B.n329 B.n328 256.663
R167 B.n328 B.n327 235.042
R168 B.n328 B.n2 235.042
R169 B.n64 B.t7 196.327
R170 B.n26 B.t2 196.327
R171 B.n135 B.t10 196.327
R172 B.n20 B.t5 196.327
R173 B.n65 B.t8 174.411
R174 B.n27 B.t1 174.411
R175 B.n136 B.t11 174.411
R176 B.n21 B.t4 174.411
R177 B.n119 B.n118 163.367
R178 B.n120 B.n119 163.367
R179 B.n120 B.n75 163.367
R180 B.n124 B.n75 163.367
R181 B.n125 B.n124 163.367
R182 B.n126 B.n125 163.367
R183 B.n126 B.n73 163.367
R184 B.n130 B.n73 163.367
R185 B.n131 B.n130 163.367
R186 B.n132 B.n131 163.367
R187 B.n132 B.n71 163.367
R188 B.n139 B.n71 163.367
R189 B.n140 B.n139 163.367
R190 B.n141 B.n140 163.367
R191 B.n141 B.n69 163.367
R192 B.n145 B.n69 163.367
R193 B.n146 B.n145 163.367
R194 B.n147 B.n146 163.367
R195 B.n147 B.n67 163.367
R196 B.n151 B.n67 163.367
R197 B.n152 B.n151 163.367
R198 B.n153 B.n152 163.367
R199 B.n153 B.n63 163.367
R200 B.n158 B.n63 163.367
R201 B.n159 B.n158 163.367
R202 B.n160 B.n159 163.367
R203 B.n160 B.n61 163.367
R204 B.n164 B.n61 163.367
R205 B.n165 B.n164 163.367
R206 B.n166 B.n165 163.367
R207 B.n166 B.n59 163.367
R208 B.n170 B.n59 163.367
R209 B.n171 B.n170 163.367
R210 B.n172 B.n171 163.367
R211 B.n172 B.n57 163.367
R212 B.n238 B.n35 163.367
R213 B.n238 B.n237 163.367
R214 B.n237 B.n236 163.367
R215 B.n236 B.n37 163.367
R216 B.n232 B.n37 163.367
R217 B.n232 B.n231 163.367
R218 B.n231 B.n230 163.367
R219 B.n230 B.n39 163.367
R220 B.n226 B.n39 163.367
R221 B.n226 B.n225 163.367
R222 B.n225 B.n224 163.367
R223 B.n224 B.n41 163.367
R224 B.n220 B.n41 163.367
R225 B.n220 B.n219 163.367
R226 B.n219 B.n218 163.367
R227 B.n218 B.n43 163.367
R228 B.n214 B.n43 163.367
R229 B.n214 B.n213 163.367
R230 B.n213 B.n212 163.367
R231 B.n212 B.n45 163.367
R232 B.n208 B.n45 163.367
R233 B.n208 B.n207 163.367
R234 B.n207 B.n206 163.367
R235 B.n206 B.n47 163.367
R236 B.n202 B.n47 163.367
R237 B.n202 B.n201 163.367
R238 B.n201 B.n200 163.367
R239 B.n200 B.n49 163.367
R240 B.n196 B.n49 163.367
R241 B.n196 B.n195 163.367
R242 B.n195 B.n194 163.367
R243 B.n194 B.n51 163.367
R244 B.n190 B.n51 163.367
R245 B.n190 B.n189 163.367
R246 B.n189 B.n188 163.367
R247 B.n188 B.n53 163.367
R248 B.n184 B.n53 163.367
R249 B.n184 B.n183 163.367
R250 B.n183 B.n182 163.367
R251 B.n182 B.n55 163.367
R252 B.n178 B.n55 163.367
R253 B.n178 B.n177 163.367
R254 B.n177 B.n176 163.367
R255 B.n296 B.n13 163.367
R256 B.n292 B.n13 163.367
R257 B.n292 B.n291 163.367
R258 B.n291 B.n290 163.367
R259 B.n290 B.n15 163.367
R260 B.n286 B.n15 163.367
R261 B.n286 B.n285 163.367
R262 B.n285 B.n284 163.367
R263 B.n284 B.n17 163.367
R264 B.n280 B.n17 163.367
R265 B.n280 B.n279 163.367
R266 B.n279 B.n278 163.367
R267 B.n278 B.n19 163.367
R268 B.n273 B.n19 163.367
R269 B.n273 B.n272 163.367
R270 B.n272 B.n271 163.367
R271 B.n271 B.n23 163.367
R272 B.n267 B.n23 163.367
R273 B.n267 B.n266 163.367
R274 B.n266 B.n265 163.367
R275 B.n265 B.n25 163.367
R276 B.n261 B.n25 163.367
R277 B.n261 B.n260 163.367
R278 B.n260 B.n29 163.367
R279 B.n256 B.n29 163.367
R280 B.n256 B.n255 163.367
R281 B.n255 B.n254 163.367
R282 B.n254 B.n31 163.367
R283 B.n250 B.n31 163.367
R284 B.n250 B.n249 163.367
R285 B.n249 B.n248 163.367
R286 B.n248 B.n33 163.367
R287 B.n244 B.n33 163.367
R288 B.n244 B.n243 163.367
R289 B.n243 B.n242 163.367
R290 B.n298 B.n297 163.367
R291 B.n298 B.n11 163.367
R292 B.n302 B.n11 163.367
R293 B.n303 B.n302 163.367
R294 B.n304 B.n303 163.367
R295 B.n304 B.n9 163.367
R296 B.n308 B.n9 163.367
R297 B.n309 B.n308 163.367
R298 B.n310 B.n309 163.367
R299 B.n310 B.n7 163.367
R300 B.n314 B.n7 163.367
R301 B.n315 B.n314 163.367
R302 B.n316 B.n315 163.367
R303 B.n316 B.n5 163.367
R304 B.n320 B.n5 163.367
R305 B.n321 B.n320 163.367
R306 B.n322 B.n321 163.367
R307 B.n322 B.n3 163.367
R308 B.n326 B.n3 163.367
R309 B.n327 B.n326 163.367
R310 B.n88 B.n2 163.367
R311 B.n89 B.n88 163.367
R312 B.n90 B.n89 163.367
R313 B.n90 B.n85 163.367
R314 B.n94 B.n85 163.367
R315 B.n95 B.n94 163.367
R316 B.n96 B.n95 163.367
R317 B.n96 B.n83 163.367
R318 B.n100 B.n83 163.367
R319 B.n101 B.n100 163.367
R320 B.n102 B.n101 163.367
R321 B.n102 B.n81 163.367
R322 B.n106 B.n81 163.367
R323 B.n107 B.n106 163.367
R324 B.n108 B.n107 163.367
R325 B.n108 B.n79 163.367
R326 B.n112 B.n79 163.367
R327 B.n113 B.n112 163.367
R328 B.n114 B.n113 163.367
R329 B.n114 B.n77 163.367
R330 B.n137 B.n136 59.5399
R331 B.n155 B.n65 59.5399
R332 B.n28 B.n27 59.5399
R333 B.n276 B.n21 59.5399
R334 B.n295 B.n12 30.7517
R335 B.n241 B.n240 30.7517
R336 B.n175 B.n174 30.7517
R337 B.n117 B.n116 30.7517
R338 B.n136 B.n135 21.9157
R339 B.n65 B.n64 21.9157
R340 B.n27 B.n26 21.9157
R341 B.n21 B.n20 21.9157
R342 B B.n329 18.0485
R343 B.n299 B.n12 10.6151
R344 B.n300 B.n299 10.6151
R345 B.n301 B.n300 10.6151
R346 B.n301 B.n10 10.6151
R347 B.n305 B.n10 10.6151
R348 B.n306 B.n305 10.6151
R349 B.n307 B.n306 10.6151
R350 B.n307 B.n8 10.6151
R351 B.n311 B.n8 10.6151
R352 B.n312 B.n311 10.6151
R353 B.n313 B.n312 10.6151
R354 B.n313 B.n6 10.6151
R355 B.n317 B.n6 10.6151
R356 B.n318 B.n317 10.6151
R357 B.n319 B.n318 10.6151
R358 B.n319 B.n4 10.6151
R359 B.n323 B.n4 10.6151
R360 B.n324 B.n323 10.6151
R361 B.n325 B.n324 10.6151
R362 B.n325 B.n0 10.6151
R363 B.n295 B.n294 10.6151
R364 B.n294 B.n293 10.6151
R365 B.n293 B.n14 10.6151
R366 B.n289 B.n14 10.6151
R367 B.n289 B.n288 10.6151
R368 B.n288 B.n287 10.6151
R369 B.n287 B.n16 10.6151
R370 B.n283 B.n16 10.6151
R371 B.n283 B.n282 10.6151
R372 B.n282 B.n281 10.6151
R373 B.n281 B.n18 10.6151
R374 B.n277 B.n18 10.6151
R375 B.n275 B.n274 10.6151
R376 B.n274 B.n22 10.6151
R377 B.n270 B.n22 10.6151
R378 B.n270 B.n269 10.6151
R379 B.n269 B.n268 10.6151
R380 B.n268 B.n24 10.6151
R381 B.n264 B.n24 10.6151
R382 B.n264 B.n263 10.6151
R383 B.n263 B.n262 10.6151
R384 B.n259 B.n258 10.6151
R385 B.n258 B.n257 10.6151
R386 B.n257 B.n30 10.6151
R387 B.n253 B.n30 10.6151
R388 B.n253 B.n252 10.6151
R389 B.n252 B.n251 10.6151
R390 B.n251 B.n32 10.6151
R391 B.n247 B.n32 10.6151
R392 B.n247 B.n246 10.6151
R393 B.n246 B.n245 10.6151
R394 B.n245 B.n34 10.6151
R395 B.n241 B.n34 10.6151
R396 B.n240 B.n239 10.6151
R397 B.n239 B.n36 10.6151
R398 B.n235 B.n36 10.6151
R399 B.n235 B.n234 10.6151
R400 B.n234 B.n233 10.6151
R401 B.n233 B.n38 10.6151
R402 B.n229 B.n38 10.6151
R403 B.n229 B.n228 10.6151
R404 B.n228 B.n227 10.6151
R405 B.n227 B.n40 10.6151
R406 B.n223 B.n40 10.6151
R407 B.n223 B.n222 10.6151
R408 B.n222 B.n221 10.6151
R409 B.n221 B.n42 10.6151
R410 B.n217 B.n42 10.6151
R411 B.n217 B.n216 10.6151
R412 B.n216 B.n215 10.6151
R413 B.n215 B.n44 10.6151
R414 B.n211 B.n44 10.6151
R415 B.n211 B.n210 10.6151
R416 B.n210 B.n209 10.6151
R417 B.n209 B.n46 10.6151
R418 B.n205 B.n46 10.6151
R419 B.n205 B.n204 10.6151
R420 B.n204 B.n203 10.6151
R421 B.n203 B.n48 10.6151
R422 B.n199 B.n48 10.6151
R423 B.n199 B.n198 10.6151
R424 B.n198 B.n197 10.6151
R425 B.n197 B.n50 10.6151
R426 B.n193 B.n50 10.6151
R427 B.n193 B.n192 10.6151
R428 B.n192 B.n191 10.6151
R429 B.n191 B.n52 10.6151
R430 B.n187 B.n52 10.6151
R431 B.n187 B.n186 10.6151
R432 B.n186 B.n185 10.6151
R433 B.n185 B.n54 10.6151
R434 B.n181 B.n54 10.6151
R435 B.n181 B.n180 10.6151
R436 B.n180 B.n179 10.6151
R437 B.n179 B.n56 10.6151
R438 B.n175 B.n56 10.6151
R439 B.n87 B.n1 10.6151
R440 B.n87 B.n86 10.6151
R441 B.n91 B.n86 10.6151
R442 B.n92 B.n91 10.6151
R443 B.n93 B.n92 10.6151
R444 B.n93 B.n84 10.6151
R445 B.n97 B.n84 10.6151
R446 B.n98 B.n97 10.6151
R447 B.n99 B.n98 10.6151
R448 B.n99 B.n82 10.6151
R449 B.n103 B.n82 10.6151
R450 B.n104 B.n103 10.6151
R451 B.n105 B.n104 10.6151
R452 B.n105 B.n80 10.6151
R453 B.n109 B.n80 10.6151
R454 B.n110 B.n109 10.6151
R455 B.n111 B.n110 10.6151
R456 B.n111 B.n78 10.6151
R457 B.n115 B.n78 10.6151
R458 B.n116 B.n115 10.6151
R459 B.n117 B.n76 10.6151
R460 B.n121 B.n76 10.6151
R461 B.n122 B.n121 10.6151
R462 B.n123 B.n122 10.6151
R463 B.n123 B.n74 10.6151
R464 B.n127 B.n74 10.6151
R465 B.n128 B.n127 10.6151
R466 B.n129 B.n128 10.6151
R467 B.n129 B.n72 10.6151
R468 B.n133 B.n72 10.6151
R469 B.n134 B.n133 10.6151
R470 B.n138 B.n134 10.6151
R471 B.n142 B.n70 10.6151
R472 B.n143 B.n142 10.6151
R473 B.n144 B.n143 10.6151
R474 B.n144 B.n68 10.6151
R475 B.n148 B.n68 10.6151
R476 B.n149 B.n148 10.6151
R477 B.n150 B.n149 10.6151
R478 B.n150 B.n66 10.6151
R479 B.n154 B.n66 10.6151
R480 B.n157 B.n156 10.6151
R481 B.n157 B.n62 10.6151
R482 B.n161 B.n62 10.6151
R483 B.n162 B.n161 10.6151
R484 B.n163 B.n162 10.6151
R485 B.n163 B.n60 10.6151
R486 B.n167 B.n60 10.6151
R487 B.n168 B.n167 10.6151
R488 B.n169 B.n168 10.6151
R489 B.n169 B.n58 10.6151
R490 B.n173 B.n58 10.6151
R491 B.n174 B.n173 10.6151
R492 B.n277 B.n276 9.36635
R493 B.n259 B.n28 9.36635
R494 B.n138 B.n137 9.36635
R495 B.n156 B.n155 9.36635
R496 B.n329 B.n0 8.11757
R497 B.n329 B.n1 8.11757
R498 B.n276 B.n275 1.24928
R499 B.n262 B.n28 1.24928
R500 B.n137 B.n70 1.24928
R501 B.n155 B.n154 1.24928
R502 VN.n5 VN.n4 161.3
R503 VN.n11 VN.n10 161.3
R504 VN.n9 VN.n6 161.3
R505 VN.n3 VN.n0 161.3
R506 VN.n1 VN.t0 142.481
R507 VN.n7 VN.t4 142.481
R508 VN.n2 VN.t5 118.995
R509 VN.n4 VN.t1 118.995
R510 VN.n8 VN.t3 118.995
R511 VN.n10 VN.t2 118.995
R512 VN.n7 VN.n6 44.8973
R513 VN.n1 VN.n0 44.8973
R514 VN VN.n11 34.741
R515 VN.n4 VN.n3 33.5944
R516 VN.n10 VN.n9 33.5944
R517 VN.n2 VN.n1 18.1882
R518 VN.n8 VN.n7 18.1882
R519 VN.n3 VN.n2 14.6066
R520 VN.n9 VN.n8 14.6066
R521 VN.n11 VN.n6 0.189894
R522 VN.n5 VN.n0 0.189894
R523 VN VN.n5 0.0516364
R524 VTAIL.n7 VTAIL.t6 168.297
R525 VTAIL.n10 VTAIL.t5 168.297
R526 VTAIL.n11 VTAIL.t10 168.297
R527 VTAIL.n2 VTAIL.t3 168.297
R528 VTAIL.n9 VTAIL.n8 154.286
R529 VTAIL.n6 VTAIL.n5 154.286
R530 VTAIL.n1 VTAIL.n0 154.286
R531 VTAIL.n4 VTAIL.n3 154.286
R532 VTAIL.n6 VTAIL.n4 16.3152
R533 VTAIL.n11 VTAIL.n10 15.341
R534 VTAIL.n0 VTAIL.t11 14.0113
R535 VTAIL.n0 VTAIL.t8 14.0113
R536 VTAIL.n3 VTAIL.t0 14.0113
R537 VTAIL.n3 VTAIL.t1 14.0113
R538 VTAIL.n8 VTAIL.t4 14.0113
R539 VTAIL.n8 VTAIL.t2 14.0113
R540 VTAIL.n5 VTAIL.t9 14.0113
R541 VTAIL.n5 VTAIL.t7 14.0113
R542 VTAIL.n7 VTAIL.n6 0.974638
R543 VTAIL.n10 VTAIL.n9 0.974638
R544 VTAIL.n4 VTAIL.n2 0.974638
R545 VTAIL.n9 VTAIL.n7 0.957397
R546 VTAIL.n2 VTAIL.n1 0.957397
R547 VTAIL VTAIL.n11 0.672914
R548 VTAIL VTAIL.n1 0.302224
R549 VDD2.n1 VDD2.t5 185.65
R550 VDD2.n2 VDD2.t3 184.975
R551 VDD2.n1 VDD2.n0 171.153
R552 VDD2 VDD2.n3 171.149
R553 VDD2.n2 VDD2.n1 28.8812
R554 VDD2.n3 VDD2.t2 14.0113
R555 VDD2.n3 VDD2.t1 14.0113
R556 VDD2.n0 VDD2.t0 14.0113
R557 VDD2.n0 VDD2.t4 14.0113
R558 VDD2 VDD2.n2 0.789293
R559 VP.n15 VP.n14 161.3
R560 VP.n5 VP.n2 161.3
R561 VP.n7 VP.n6 161.3
R562 VP.n13 VP.n0 161.3
R563 VP.n12 VP.n11 161.3
R564 VP.n10 VP.n1 161.3
R565 VP.n9 VP.n8 161.3
R566 VP.n3 VP.t5 142.481
R567 VP.n8 VP.t1 118.995
R568 VP.n12 VP.t3 118.995
R569 VP.n14 VP.t0 118.995
R570 VP.n6 VP.t2 118.995
R571 VP.n4 VP.t4 118.995
R572 VP.n3 VP.n2 44.8973
R573 VP.n9 VP.n7 34.3603
R574 VP.n8 VP.n1 33.5944
R575 VP.n14 VP.n13 33.5944
R576 VP.n6 VP.n5 33.5944
R577 VP.n4 VP.n3 18.1882
R578 VP.n12 VP.n1 14.6066
R579 VP.n13 VP.n12 14.6066
R580 VP.n5 VP.n4 14.6066
R581 VP.n7 VP.n2 0.189894
R582 VP.n10 VP.n9 0.189894
R583 VP.n11 VP.n10 0.189894
R584 VP.n11 VP.n0 0.189894
R585 VP.n15 VP.n0 0.189894
R586 VP VP.n15 0.0516364
R587 VDD1 VDD1.t0 185.763
R588 VDD1.n1 VDD1.t4 185.65
R589 VDD1.n1 VDD1.n0 171.153
R590 VDD1.n3 VDD1.n2 170.964
R591 VDD1.n3 VDD1.n1 29.9513
R592 VDD1.n2 VDD1.t1 14.0113
R593 VDD1.n2 VDD1.t3 14.0113
R594 VDD1.n0 VDD1.t2 14.0113
R595 VDD1.n0 VDD1.t5 14.0113
R596 VDD1 VDD1.n3 0.185845
C0 VDD2 VTAIL 3.44199f
C1 VP VTAIL 1.3943f
C2 VP VDD2 0.311419f
C3 VTAIL VDD1 3.40177f
C4 VDD2 VDD1 0.743611f
C5 VTAIL VN 1.3801f
C6 VDD2 VN 1.17068f
C7 w_n1874_n1432# VTAIL 1.37107f
C8 w_n1874_n1432# VDD2 1.14697f
C9 VP VDD1 1.32584f
C10 B VTAIL 0.977978f
C11 B VDD2 0.910602f
C12 VP VN 3.38594f
C13 w_n1874_n1432# VP 3.13106f
C14 VDD1 VN 0.154419f
C15 B VP 1.0503f
C16 w_n1874_n1432# VDD1 1.12033f
C17 w_n1874_n1432# VN 2.89738f
C18 B VDD1 0.879133f
C19 B VN 0.663852f
C20 B w_n1874_n1432# 4.47148f
C21 VDD2 VSUBS 0.732818f
C22 VDD1 VSUBS 0.986498f
C23 VTAIL VSUBS 0.320546f
C24 VN VSUBS 3.30242f
C25 VP VSUBS 1.085994f
C26 B VSUBS 1.939325f
C27 w_n1874_n1432# VSUBS 34.1593f
C28 VDD1.t0 VSUBS 0.209128f
C29 VDD1.t4 VSUBS 0.208947f
C30 VDD1.t2 VSUBS 0.03086f
C31 VDD1.t5 VSUBS 0.03086f
C32 VDD1.n0 VSUBS 0.138665f
C33 VDD1.n1 VSUBS 1.19329f
C34 VDD1.t1 VSUBS 0.03086f
C35 VDD1.t3 VSUBS 0.03086f
C36 VDD1.n2 VSUBS 0.138369f
C37 VDD1.n3 VSUBS 1.07426f
C38 VP.n0 VSUBS 0.052505f
C39 VP.n1 VSUBS 0.011915f
C40 VP.n2 VSUBS 0.227009f
C41 VP.t2 VSUBS 0.29782f
C42 VP.t4 VSUBS 0.29782f
C43 VP.t5 VSUBS 0.329439f
C44 VP.n3 VSUBS 0.164926f
C45 VP.n4 VSUBS 0.194673f
C46 VP.n5 VSUBS 0.011915f
C47 VP.n6 VSUBS 0.189567f
C48 VP.n7 VSUBS 1.50929f
C49 VP.t1 VSUBS 0.29782f
C50 VP.n8 VSUBS 0.189567f
C51 VP.n9 VSUBS 1.56437f
C52 VP.n10 VSUBS 0.052505f
C53 VP.n11 VSUBS 0.052505f
C54 VP.t3 VSUBS 0.29782f
C55 VP.n12 VSUBS 0.188596f
C56 VP.n13 VSUBS 0.011915f
C57 VP.t0 VSUBS 0.29782f
C58 VP.n14 VSUBS 0.189567f
C59 VP.n15 VSUBS 0.04069f
C60 VDD2.t5 VSUBS 0.212839f
C61 VDD2.t0 VSUBS 0.031435f
C62 VDD2.t4 VSUBS 0.031435f
C63 VDD2.n0 VSUBS 0.141248f
C64 VDD2.n1 VSUBS 1.16465f
C65 VDD2.t3 VSUBS 0.211889f
C66 VDD2.n2 VSUBS 1.07611f
C67 VDD2.t2 VSUBS 0.031435f
C68 VDD2.t1 VSUBS 0.031435f
C69 VDD2.n3 VSUBS 0.141242f
C70 VTAIL.t11 VSUBS 0.038947f
C71 VTAIL.t8 VSUBS 0.038947f
C72 VTAIL.n0 VSUBS 0.148036f
C73 VTAIL.n1 VSUBS 0.333883f
C74 VTAIL.t3 VSUBS 0.23633f
C75 VTAIL.n2 VSUBS 0.397835f
C76 VTAIL.t0 VSUBS 0.038947f
C77 VTAIL.t1 VSUBS 0.038947f
C78 VTAIL.n3 VSUBS 0.148036f
C79 VTAIL.n4 VSUBS 0.873246f
C80 VTAIL.t9 VSUBS 0.038947f
C81 VTAIL.t7 VSUBS 0.038947f
C82 VTAIL.n5 VSUBS 0.148037f
C83 VTAIL.n6 VSUBS 0.873245f
C84 VTAIL.t6 VSUBS 0.236331f
C85 VTAIL.n7 VSUBS 0.397835f
C86 VTAIL.t4 VSUBS 0.038947f
C87 VTAIL.t2 VSUBS 0.038947f
C88 VTAIL.n8 VSUBS 0.148037f
C89 VTAIL.n9 VSUBS 0.37991f
C90 VTAIL.t5 VSUBS 0.236331f
C91 VTAIL.n10 VSUBS 0.824488f
C92 VTAIL.t10 VSUBS 0.23633f
C93 VTAIL.n11 VSUBS 0.803835f
C94 VN.n0 VSUBS 0.217554f
C95 VN.t0 VSUBS 0.315717f
C96 VN.n1 VSUBS 0.158057f
C97 VN.t5 VSUBS 0.285416f
C98 VN.n2 VSUBS 0.186564f
C99 VN.n3 VSUBS 0.011418f
C100 VN.t1 VSUBS 0.285416f
C101 VN.n4 VSUBS 0.181671f
C102 VN.n5 VSUBS 0.038995f
C103 VN.n6 VSUBS 0.217554f
C104 VN.t4 VSUBS 0.315717f
C105 VN.n7 VSUBS 0.158057f
C106 VN.t3 VSUBS 0.285416f
C107 VN.n8 VSUBS 0.186564f
C108 VN.n9 VSUBS 0.011418f
C109 VN.t2 VSUBS 0.285416f
C110 VN.n10 VSUBS 0.181671f
C111 VN.n11 VSUBS 1.47992f
C112 B.n0 VSUBS 0.007555f
C113 B.n1 VSUBS 0.007555f
C114 B.n2 VSUBS 0.011173f
C115 B.n3 VSUBS 0.008562f
C116 B.n4 VSUBS 0.008562f
C117 B.n5 VSUBS 0.008562f
C118 B.n6 VSUBS 0.008562f
C119 B.n7 VSUBS 0.008562f
C120 B.n8 VSUBS 0.008562f
C121 B.n9 VSUBS 0.008562f
C122 B.n10 VSUBS 0.008562f
C123 B.n11 VSUBS 0.008562f
C124 B.n12 VSUBS 0.01878f
C125 B.n13 VSUBS 0.008562f
C126 B.n14 VSUBS 0.008562f
C127 B.n15 VSUBS 0.008562f
C128 B.n16 VSUBS 0.008562f
C129 B.n17 VSUBS 0.008562f
C130 B.n18 VSUBS 0.008562f
C131 B.n19 VSUBS 0.008562f
C132 B.t4 VSUBS 0.06319f
C133 B.t5 VSUBS 0.069167f
C134 B.t3 VSUBS 0.107057f
C135 B.n20 VSUBS 0.072648f
C136 B.n21 VSUBS 0.065759f
C137 B.n22 VSUBS 0.008562f
C138 B.n23 VSUBS 0.008562f
C139 B.n24 VSUBS 0.008562f
C140 B.n25 VSUBS 0.008562f
C141 B.t1 VSUBS 0.06319f
C142 B.t2 VSUBS 0.069167f
C143 B.t0 VSUBS 0.107057f
C144 B.n26 VSUBS 0.072648f
C145 B.n27 VSUBS 0.065759f
C146 B.n28 VSUBS 0.019838f
C147 B.n29 VSUBS 0.008562f
C148 B.n30 VSUBS 0.008562f
C149 B.n31 VSUBS 0.008562f
C150 B.n32 VSUBS 0.008562f
C151 B.n33 VSUBS 0.008562f
C152 B.n34 VSUBS 0.008562f
C153 B.n35 VSUBS 0.01878f
C154 B.n36 VSUBS 0.008562f
C155 B.n37 VSUBS 0.008562f
C156 B.n38 VSUBS 0.008562f
C157 B.n39 VSUBS 0.008562f
C158 B.n40 VSUBS 0.008562f
C159 B.n41 VSUBS 0.008562f
C160 B.n42 VSUBS 0.008562f
C161 B.n43 VSUBS 0.008562f
C162 B.n44 VSUBS 0.008562f
C163 B.n45 VSUBS 0.008562f
C164 B.n46 VSUBS 0.008562f
C165 B.n47 VSUBS 0.008562f
C166 B.n48 VSUBS 0.008562f
C167 B.n49 VSUBS 0.008562f
C168 B.n50 VSUBS 0.008562f
C169 B.n51 VSUBS 0.008562f
C170 B.n52 VSUBS 0.008562f
C171 B.n53 VSUBS 0.008562f
C172 B.n54 VSUBS 0.008562f
C173 B.n55 VSUBS 0.008562f
C174 B.n56 VSUBS 0.008562f
C175 B.n57 VSUBS 0.01975f
C176 B.n58 VSUBS 0.008562f
C177 B.n59 VSUBS 0.008562f
C178 B.n60 VSUBS 0.008562f
C179 B.n61 VSUBS 0.008562f
C180 B.n62 VSUBS 0.008562f
C181 B.n63 VSUBS 0.008562f
C182 B.t8 VSUBS 0.06319f
C183 B.t7 VSUBS 0.069167f
C184 B.t6 VSUBS 0.107057f
C185 B.n64 VSUBS 0.072648f
C186 B.n65 VSUBS 0.065759f
C187 B.n66 VSUBS 0.008562f
C188 B.n67 VSUBS 0.008562f
C189 B.n68 VSUBS 0.008562f
C190 B.n69 VSUBS 0.008562f
C191 B.n70 VSUBS 0.004785f
C192 B.n71 VSUBS 0.008562f
C193 B.n72 VSUBS 0.008562f
C194 B.n73 VSUBS 0.008562f
C195 B.n74 VSUBS 0.008562f
C196 B.n75 VSUBS 0.008562f
C197 B.n76 VSUBS 0.008562f
C198 B.n77 VSUBS 0.01878f
C199 B.n78 VSUBS 0.008562f
C200 B.n79 VSUBS 0.008562f
C201 B.n80 VSUBS 0.008562f
C202 B.n81 VSUBS 0.008562f
C203 B.n82 VSUBS 0.008562f
C204 B.n83 VSUBS 0.008562f
C205 B.n84 VSUBS 0.008562f
C206 B.n85 VSUBS 0.008562f
C207 B.n86 VSUBS 0.008562f
C208 B.n87 VSUBS 0.008562f
C209 B.n88 VSUBS 0.008562f
C210 B.n89 VSUBS 0.008562f
C211 B.n90 VSUBS 0.008562f
C212 B.n91 VSUBS 0.008562f
C213 B.n92 VSUBS 0.008562f
C214 B.n93 VSUBS 0.008562f
C215 B.n94 VSUBS 0.008562f
C216 B.n95 VSUBS 0.008562f
C217 B.n96 VSUBS 0.008562f
C218 B.n97 VSUBS 0.008562f
C219 B.n98 VSUBS 0.008562f
C220 B.n99 VSUBS 0.008562f
C221 B.n100 VSUBS 0.008562f
C222 B.n101 VSUBS 0.008562f
C223 B.n102 VSUBS 0.008562f
C224 B.n103 VSUBS 0.008562f
C225 B.n104 VSUBS 0.008562f
C226 B.n105 VSUBS 0.008562f
C227 B.n106 VSUBS 0.008562f
C228 B.n107 VSUBS 0.008562f
C229 B.n108 VSUBS 0.008562f
C230 B.n109 VSUBS 0.008562f
C231 B.n110 VSUBS 0.008562f
C232 B.n111 VSUBS 0.008562f
C233 B.n112 VSUBS 0.008562f
C234 B.n113 VSUBS 0.008562f
C235 B.n114 VSUBS 0.008562f
C236 B.n115 VSUBS 0.008562f
C237 B.n116 VSUBS 0.01878f
C238 B.n117 VSUBS 0.01975f
C239 B.n118 VSUBS 0.01975f
C240 B.n119 VSUBS 0.008562f
C241 B.n120 VSUBS 0.008562f
C242 B.n121 VSUBS 0.008562f
C243 B.n122 VSUBS 0.008562f
C244 B.n123 VSUBS 0.008562f
C245 B.n124 VSUBS 0.008562f
C246 B.n125 VSUBS 0.008562f
C247 B.n126 VSUBS 0.008562f
C248 B.n127 VSUBS 0.008562f
C249 B.n128 VSUBS 0.008562f
C250 B.n129 VSUBS 0.008562f
C251 B.n130 VSUBS 0.008562f
C252 B.n131 VSUBS 0.008562f
C253 B.n132 VSUBS 0.008562f
C254 B.n133 VSUBS 0.008562f
C255 B.n134 VSUBS 0.008562f
C256 B.t11 VSUBS 0.06319f
C257 B.t10 VSUBS 0.069167f
C258 B.t9 VSUBS 0.107057f
C259 B.n135 VSUBS 0.072648f
C260 B.n136 VSUBS 0.065759f
C261 B.n137 VSUBS 0.019838f
C262 B.n138 VSUBS 0.008059f
C263 B.n139 VSUBS 0.008562f
C264 B.n140 VSUBS 0.008562f
C265 B.n141 VSUBS 0.008562f
C266 B.n142 VSUBS 0.008562f
C267 B.n143 VSUBS 0.008562f
C268 B.n144 VSUBS 0.008562f
C269 B.n145 VSUBS 0.008562f
C270 B.n146 VSUBS 0.008562f
C271 B.n147 VSUBS 0.008562f
C272 B.n148 VSUBS 0.008562f
C273 B.n149 VSUBS 0.008562f
C274 B.n150 VSUBS 0.008562f
C275 B.n151 VSUBS 0.008562f
C276 B.n152 VSUBS 0.008562f
C277 B.n153 VSUBS 0.008562f
C278 B.n154 VSUBS 0.004785f
C279 B.n155 VSUBS 0.019838f
C280 B.n156 VSUBS 0.008059f
C281 B.n157 VSUBS 0.008562f
C282 B.n158 VSUBS 0.008562f
C283 B.n159 VSUBS 0.008562f
C284 B.n160 VSUBS 0.008562f
C285 B.n161 VSUBS 0.008562f
C286 B.n162 VSUBS 0.008562f
C287 B.n163 VSUBS 0.008562f
C288 B.n164 VSUBS 0.008562f
C289 B.n165 VSUBS 0.008562f
C290 B.n166 VSUBS 0.008562f
C291 B.n167 VSUBS 0.008562f
C292 B.n168 VSUBS 0.008562f
C293 B.n169 VSUBS 0.008562f
C294 B.n170 VSUBS 0.008562f
C295 B.n171 VSUBS 0.008562f
C296 B.n172 VSUBS 0.008562f
C297 B.n173 VSUBS 0.008562f
C298 B.n174 VSUBS 0.018675f
C299 B.n175 VSUBS 0.019855f
C300 B.n176 VSUBS 0.01878f
C301 B.n177 VSUBS 0.008562f
C302 B.n178 VSUBS 0.008562f
C303 B.n179 VSUBS 0.008562f
C304 B.n180 VSUBS 0.008562f
C305 B.n181 VSUBS 0.008562f
C306 B.n182 VSUBS 0.008562f
C307 B.n183 VSUBS 0.008562f
C308 B.n184 VSUBS 0.008562f
C309 B.n185 VSUBS 0.008562f
C310 B.n186 VSUBS 0.008562f
C311 B.n187 VSUBS 0.008562f
C312 B.n188 VSUBS 0.008562f
C313 B.n189 VSUBS 0.008562f
C314 B.n190 VSUBS 0.008562f
C315 B.n191 VSUBS 0.008562f
C316 B.n192 VSUBS 0.008562f
C317 B.n193 VSUBS 0.008562f
C318 B.n194 VSUBS 0.008562f
C319 B.n195 VSUBS 0.008562f
C320 B.n196 VSUBS 0.008562f
C321 B.n197 VSUBS 0.008562f
C322 B.n198 VSUBS 0.008562f
C323 B.n199 VSUBS 0.008562f
C324 B.n200 VSUBS 0.008562f
C325 B.n201 VSUBS 0.008562f
C326 B.n202 VSUBS 0.008562f
C327 B.n203 VSUBS 0.008562f
C328 B.n204 VSUBS 0.008562f
C329 B.n205 VSUBS 0.008562f
C330 B.n206 VSUBS 0.008562f
C331 B.n207 VSUBS 0.008562f
C332 B.n208 VSUBS 0.008562f
C333 B.n209 VSUBS 0.008562f
C334 B.n210 VSUBS 0.008562f
C335 B.n211 VSUBS 0.008562f
C336 B.n212 VSUBS 0.008562f
C337 B.n213 VSUBS 0.008562f
C338 B.n214 VSUBS 0.008562f
C339 B.n215 VSUBS 0.008562f
C340 B.n216 VSUBS 0.008562f
C341 B.n217 VSUBS 0.008562f
C342 B.n218 VSUBS 0.008562f
C343 B.n219 VSUBS 0.008562f
C344 B.n220 VSUBS 0.008562f
C345 B.n221 VSUBS 0.008562f
C346 B.n222 VSUBS 0.008562f
C347 B.n223 VSUBS 0.008562f
C348 B.n224 VSUBS 0.008562f
C349 B.n225 VSUBS 0.008562f
C350 B.n226 VSUBS 0.008562f
C351 B.n227 VSUBS 0.008562f
C352 B.n228 VSUBS 0.008562f
C353 B.n229 VSUBS 0.008562f
C354 B.n230 VSUBS 0.008562f
C355 B.n231 VSUBS 0.008562f
C356 B.n232 VSUBS 0.008562f
C357 B.n233 VSUBS 0.008562f
C358 B.n234 VSUBS 0.008562f
C359 B.n235 VSUBS 0.008562f
C360 B.n236 VSUBS 0.008562f
C361 B.n237 VSUBS 0.008562f
C362 B.n238 VSUBS 0.008562f
C363 B.n239 VSUBS 0.008562f
C364 B.n240 VSUBS 0.01878f
C365 B.n241 VSUBS 0.01975f
C366 B.n242 VSUBS 0.01975f
C367 B.n243 VSUBS 0.008562f
C368 B.n244 VSUBS 0.008562f
C369 B.n245 VSUBS 0.008562f
C370 B.n246 VSUBS 0.008562f
C371 B.n247 VSUBS 0.008562f
C372 B.n248 VSUBS 0.008562f
C373 B.n249 VSUBS 0.008562f
C374 B.n250 VSUBS 0.008562f
C375 B.n251 VSUBS 0.008562f
C376 B.n252 VSUBS 0.008562f
C377 B.n253 VSUBS 0.008562f
C378 B.n254 VSUBS 0.008562f
C379 B.n255 VSUBS 0.008562f
C380 B.n256 VSUBS 0.008562f
C381 B.n257 VSUBS 0.008562f
C382 B.n258 VSUBS 0.008562f
C383 B.n259 VSUBS 0.008059f
C384 B.n260 VSUBS 0.008562f
C385 B.n261 VSUBS 0.008562f
C386 B.n262 VSUBS 0.004785f
C387 B.n263 VSUBS 0.008562f
C388 B.n264 VSUBS 0.008562f
C389 B.n265 VSUBS 0.008562f
C390 B.n266 VSUBS 0.008562f
C391 B.n267 VSUBS 0.008562f
C392 B.n268 VSUBS 0.008562f
C393 B.n269 VSUBS 0.008562f
C394 B.n270 VSUBS 0.008562f
C395 B.n271 VSUBS 0.008562f
C396 B.n272 VSUBS 0.008562f
C397 B.n273 VSUBS 0.008562f
C398 B.n274 VSUBS 0.008562f
C399 B.n275 VSUBS 0.004785f
C400 B.n276 VSUBS 0.019838f
C401 B.n277 VSUBS 0.008059f
C402 B.n278 VSUBS 0.008562f
C403 B.n279 VSUBS 0.008562f
C404 B.n280 VSUBS 0.008562f
C405 B.n281 VSUBS 0.008562f
C406 B.n282 VSUBS 0.008562f
C407 B.n283 VSUBS 0.008562f
C408 B.n284 VSUBS 0.008562f
C409 B.n285 VSUBS 0.008562f
C410 B.n286 VSUBS 0.008562f
C411 B.n287 VSUBS 0.008562f
C412 B.n288 VSUBS 0.008562f
C413 B.n289 VSUBS 0.008562f
C414 B.n290 VSUBS 0.008562f
C415 B.n291 VSUBS 0.008562f
C416 B.n292 VSUBS 0.008562f
C417 B.n293 VSUBS 0.008562f
C418 B.n294 VSUBS 0.008562f
C419 B.n295 VSUBS 0.01975f
C420 B.n296 VSUBS 0.01975f
C421 B.n297 VSUBS 0.01878f
C422 B.n298 VSUBS 0.008562f
C423 B.n299 VSUBS 0.008562f
C424 B.n300 VSUBS 0.008562f
C425 B.n301 VSUBS 0.008562f
C426 B.n302 VSUBS 0.008562f
C427 B.n303 VSUBS 0.008562f
C428 B.n304 VSUBS 0.008562f
C429 B.n305 VSUBS 0.008562f
C430 B.n306 VSUBS 0.008562f
C431 B.n307 VSUBS 0.008562f
C432 B.n308 VSUBS 0.008562f
C433 B.n309 VSUBS 0.008562f
C434 B.n310 VSUBS 0.008562f
C435 B.n311 VSUBS 0.008562f
C436 B.n312 VSUBS 0.008562f
C437 B.n313 VSUBS 0.008562f
C438 B.n314 VSUBS 0.008562f
C439 B.n315 VSUBS 0.008562f
C440 B.n316 VSUBS 0.008562f
C441 B.n317 VSUBS 0.008562f
C442 B.n318 VSUBS 0.008562f
C443 B.n319 VSUBS 0.008562f
C444 B.n320 VSUBS 0.008562f
C445 B.n321 VSUBS 0.008562f
C446 B.n322 VSUBS 0.008562f
C447 B.n323 VSUBS 0.008562f
C448 B.n324 VSUBS 0.008562f
C449 B.n325 VSUBS 0.008562f
C450 B.n326 VSUBS 0.008562f
C451 B.n327 VSUBS 0.011173f
C452 B.n328 VSUBS 0.011902f
C453 B.n329 VSUBS 0.023669f
.ends

