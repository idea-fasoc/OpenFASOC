* NGSPICE file created from diff_pair_sample_1475.ext - technology: sky130A

.subckt diff_pair_sample_1475 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t3 VN.t0 VTAIL.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=0.1221 pd=1.07 as=0.2886 ps=2.26 w=0.74 l=2.26
X1 VTAIL.t3 VP.t0 VDD1.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.2886 pd=2.26 as=0.1221 ps=1.07 w=0.74 l=2.26
X2 VDD1.t2 VP.t1 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.1221 pd=1.07 as=0.2886 ps=2.26 w=0.74 l=2.26
X3 VTAIL.t5 VN.t1 VDD2.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=0.2886 pd=2.26 as=0.1221 ps=1.07 w=0.74 l=2.26
X4 VTAIL.t0 VP.t2 VDD1.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=0.2886 pd=2.26 as=0.1221 ps=1.07 w=0.74 l=2.26
X5 VDD1.t0 VP.t3 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.1221 pd=1.07 as=0.2886 ps=2.26 w=0.74 l=2.26
X6 B.t17 B.t15 B.t16 B.t5 sky130_fd_pr__nfet_01v8 ad=0.2886 pd=2.26 as=0 ps=0 w=0.74 l=2.26
X7 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=0.2886 pd=2.26 as=0 ps=0 w=0.74 l=2.26
X8 VTAIL.t6 VN.t2 VDD2.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=0.2886 pd=2.26 as=0.1221 ps=1.07 w=0.74 l=2.26
X9 VDD2.t0 VN.t3 VTAIL.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=0.1221 pd=1.07 as=0.2886 ps=2.26 w=0.74 l=2.26
X10 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=0.2886 pd=2.26 as=0 ps=0 w=0.74 l=2.26
X11 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=0.2886 pd=2.26 as=0 ps=0 w=0.74 l=2.26
R0 VN.n0 VN.t2 44.0585
R1 VN.n1 VN.t3 44.0585
R2 VN.n0 VN.t0 43.4112
R3 VN.n1 VN.t1 43.4112
R4 VN VN.n1 42.642
R5 VN VN.n0 5.66096
R6 VTAIL.n7 VTAIL.t7 246.657
R7 VTAIL.n0 VTAIL.t6 246.657
R8 VTAIL.n1 VTAIL.t1 246.657
R9 VTAIL.n2 VTAIL.t3 246.657
R10 VTAIL.n6 VTAIL.t2 246.657
R11 VTAIL.n5 VTAIL.t0 246.657
R12 VTAIL.n4 VTAIL.t4 246.657
R13 VTAIL.n3 VTAIL.t5 246.657
R14 VTAIL.n7 VTAIL.n6 15.2376
R15 VTAIL.n3 VTAIL.n2 15.2376
R16 VTAIL.n4 VTAIL.n3 2.23326
R17 VTAIL.n6 VTAIL.n5 2.23326
R18 VTAIL.n2 VTAIL.n1 2.23326
R19 VTAIL VTAIL.n0 1.17507
R20 VTAIL VTAIL.n7 1.05869
R21 VTAIL.n5 VTAIL.n4 0.470328
R22 VTAIL.n1 VTAIL.n0 0.470328
R23 VDD2.n2 VDD2.n0 267.63
R24 VDD2.n2 VDD2.n1 236.579
R25 VDD2.n1 VDD2.t2 26.7573
R26 VDD2.n1 VDD2.t0 26.7573
R27 VDD2.n0 VDD2.t1 26.7573
R28 VDD2.n0 VDD2.t3 26.7573
R29 VDD2 VDD2.n2 0.0586897
R30 B.n394 B.n393 585
R31 B.n395 B.n394 585
R32 B.n127 B.n73 585
R33 B.n126 B.n125 585
R34 B.n124 B.n123 585
R35 B.n122 B.n121 585
R36 B.n120 B.n119 585
R37 B.n118 B.n117 585
R38 B.n116 B.n115 585
R39 B.n114 B.n113 585
R40 B.n112 B.n111 585
R41 B.n110 B.n109 585
R42 B.n108 B.n107 585
R43 B.n106 B.n105 585
R44 B.n104 B.n103 585
R45 B.n102 B.n101 585
R46 B.n100 B.n99 585
R47 B.n98 B.n97 585
R48 B.n96 B.n95 585
R49 B.n93 B.n92 585
R50 B.n91 B.n90 585
R51 B.n89 B.n88 585
R52 B.n87 B.n86 585
R53 B.n85 B.n84 585
R54 B.n83 B.n82 585
R55 B.n81 B.n80 585
R56 B.n60 B.n59 585
R57 B.n398 B.n397 585
R58 B.n392 B.n74 585
R59 B.n74 B.n57 585
R60 B.n391 B.n56 585
R61 B.n402 B.n56 585
R62 B.n390 B.n55 585
R63 B.n403 B.n55 585
R64 B.n389 B.n54 585
R65 B.n404 B.n54 585
R66 B.n388 B.n387 585
R67 B.n387 B.n50 585
R68 B.n386 B.n49 585
R69 B.n410 B.n49 585
R70 B.n385 B.n48 585
R71 B.n411 B.n48 585
R72 B.n384 B.n47 585
R73 B.n412 B.n47 585
R74 B.n383 B.n382 585
R75 B.n382 B.n43 585
R76 B.n381 B.n42 585
R77 B.n418 B.n42 585
R78 B.n380 B.n41 585
R79 B.n419 B.n41 585
R80 B.n379 B.n40 585
R81 B.n420 B.n40 585
R82 B.n378 B.n377 585
R83 B.n377 B.n36 585
R84 B.n376 B.n35 585
R85 B.n426 B.n35 585
R86 B.n375 B.n34 585
R87 B.n427 B.n34 585
R88 B.n374 B.n33 585
R89 B.n428 B.n33 585
R90 B.n373 B.n372 585
R91 B.n372 B.n29 585
R92 B.n371 B.n28 585
R93 B.n434 B.n28 585
R94 B.n370 B.n27 585
R95 B.n435 B.n27 585
R96 B.n369 B.n26 585
R97 B.n436 B.n26 585
R98 B.n368 B.n367 585
R99 B.n367 B.n22 585
R100 B.n366 B.n21 585
R101 B.n442 B.n21 585
R102 B.n365 B.n20 585
R103 B.n443 B.n20 585
R104 B.n364 B.n19 585
R105 B.n444 B.n19 585
R106 B.n363 B.n362 585
R107 B.n362 B.n15 585
R108 B.n361 B.n14 585
R109 B.n450 B.n14 585
R110 B.n360 B.n13 585
R111 B.n451 B.n13 585
R112 B.n359 B.n12 585
R113 B.n452 B.n12 585
R114 B.n358 B.n357 585
R115 B.n357 B.n8 585
R116 B.n356 B.n7 585
R117 B.n458 B.n7 585
R118 B.n355 B.n6 585
R119 B.n459 B.n6 585
R120 B.n354 B.n5 585
R121 B.n460 B.n5 585
R122 B.n353 B.n352 585
R123 B.n352 B.n4 585
R124 B.n351 B.n128 585
R125 B.n351 B.n350 585
R126 B.n341 B.n129 585
R127 B.n130 B.n129 585
R128 B.n343 B.n342 585
R129 B.n344 B.n343 585
R130 B.n340 B.n135 585
R131 B.n135 B.n134 585
R132 B.n339 B.n338 585
R133 B.n338 B.n337 585
R134 B.n137 B.n136 585
R135 B.n138 B.n137 585
R136 B.n330 B.n329 585
R137 B.n331 B.n330 585
R138 B.n328 B.n143 585
R139 B.n143 B.n142 585
R140 B.n327 B.n326 585
R141 B.n326 B.n325 585
R142 B.n145 B.n144 585
R143 B.n146 B.n145 585
R144 B.n318 B.n317 585
R145 B.n319 B.n318 585
R146 B.n316 B.n151 585
R147 B.n151 B.n150 585
R148 B.n315 B.n314 585
R149 B.n314 B.n313 585
R150 B.n153 B.n152 585
R151 B.n154 B.n153 585
R152 B.n306 B.n305 585
R153 B.n307 B.n306 585
R154 B.n304 B.n159 585
R155 B.n159 B.n158 585
R156 B.n303 B.n302 585
R157 B.n302 B.n301 585
R158 B.n161 B.n160 585
R159 B.n162 B.n161 585
R160 B.n294 B.n293 585
R161 B.n295 B.n294 585
R162 B.n292 B.n167 585
R163 B.n167 B.n166 585
R164 B.n291 B.n290 585
R165 B.n290 B.n289 585
R166 B.n169 B.n168 585
R167 B.n170 B.n169 585
R168 B.n282 B.n281 585
R169 B.n283 B.n282 585
R170 B.n280 B.n175 585
R171 B.n175 B.n174 585
R172 B.n279 B.n278 585
R173 B.n278 B.n277 585
R174 B.n177 B.n176 585
R175 B.n178 B.n177 585
R176 B.n270 B.n269 585
R177 B.n271 B.n270 585
R178 B.n268 B.n183 585
R179 B.n183 B.n182 585
R180 B.n267 B.n266 585
R181 B.n266 B.n265 585
R182 B.n185 B.n184 585
R183 B.n186 B.n185 585
R184 B.n261 B.n260 585
R185 B.n189 B.n188 585
R186 B.n257 B.n256 585
R187 B.n258 B.n257 585
R188 B.n255 B.n202 585
R189 B.n254 B.n253 585
R190 B.n252 B.n251 585
R191 B.n250 B.n249 585
R192 B.n248 B.n247 585
R193 B.n246 B.n245 585
R194 B.n244 B.n243 585
R195 B.n242 B.n241 585
R196 B.n240 B.n239 585
R197 B.n238 B.n237 585
R198 B.n236 B.n235 585
R199 B.n234 B.n233 585
R200 B.n232 B.n231 585
R201 B.n230 B.n229 585
R202 B.n228 B.n227 585
R203 B.n225 B.n224 585
R204 B.n223 B.n222 585
R205 B.n221 B.n220 585
R206 B.n219 B.n218 585
R207 B.n217 B.n216 585
R208 B.n215 B.n214 585
R209 B.n213 B.n212 585
R210 B.n211 B.n210 585
R211 B.n209 B.n208 585
R212 B.n262 B.n187 585
R213 B.n187 B.n186 585
R214 B.n264 B.n263 585
R215 B.n265 B.n264 585
R216 B.n181 B.n180 585
R217 B.n182 B.n181 585
R218 B.n273 B.n272 585
R219 B.n272 B.n271 585
R220 B.n274 B.n179 585
R221 B.n179 B.n178 585
R222 B.n276 B.n275 585
R223 B.n277 B.n276 585
R224 B.n173 B.n172 585
R225 B.n174 B.n173 585
R226 B.n285 B.n284 585
R227 B.n284 B.n283 585
R228 B.n286 B.n171 585
R229 B.n171 B.n170 585
R230 B.n288 B.n287 585
R231 B.n289 B.n288 585
R232 B.n165 B.n164 585
R233 B.n166 B.n165 585
R234 B.n297 B.n296 585
R235 B.n296 B.n295 585
R236 B.n298 B.n163 585
R237 B.n163 B.n162 585
R238 B.n300 B.n299 585
R239 B.n301 B.n300 585
R240 B.n157 B.n156 585
R241 B.n158 B.n157 585
R242 B.n309 B.n308 585
R243 B.n308 B.n307 585
R244 B.n310 B.n155 585
R245 B.n155 B.n154 585
R246 B.n312 B.n311 585
R247 B.n313 B.n312 585
R248 B.n149 B.n148 585
R249 B.n150 B.n149 585
R250 B.n321 B.n320 585
R251 B.n320 B.n319 585
R252 B.n322 B.n147 585
R253 B.n147 B.n146 585
R254 B.n324 B.n323 585
R255 B.n325 B.n324 585
R256 B.n141 B.n140 585
R257 B.n142 B.n141 585
R258 B.n333 B.n332 585
R259 B.n332 B.n331 585
R260 B.n334 B.n139 585
R261 B.n139 B.n138 585
R262 B.n336 B.n335 585
R263 B.n337 B.n336 585
R264 B.n133 B.n132 585
R265 B.n134 B.n133 585
R266 B.n346 B.n345 585
R267 B.n345 B.n344 585
R268 B.n347 B.n131 585
R269 B.n131 B.n130 585
R270 B.n349 B.n348 585
R271 B.n350 B.n349 585
R272 B.n2 B.n0 585
R273 B.n4 B.n2 585
R274 B.n3 B.n1 585
R275 B.n459 B.n3 585
R276 B.n457 B.n456 585
R277 B.n458 B.n457 585
R278 B.n455 B.n9 585
R279 B.n9 B.n8 585
R280 B.n454 B.n453 585
R281 B.n453 B.n452 585
R282 B.n11 B.n10 585
R283 B.n451 B.n11 585
R284 B.n449 B.n448 585
R285 B.n450 B.n449 585
R286 B.n447 B.n16 585
R287 B.n16 B.n15 585
R288 B.n446 B.n445 585
R289 B.n445 B.n444 585
R290 B.n18 B.n17 585
R291 B.n443 B.n18 585
R292 B.n441 B.n440 585
R293 B.n442 B.n441 585
R294 B.n439 B.n23 585
R295 B.n23 B.n22 585
R296 B.n438 B.n437 585
R297 B.n437 B.n436 585
R298 B.n25 B.n24 585
R299 B.n435 B.n25 585
R300 B.n433 B.n432 585
R301 B.n434 B.n433 585
R302 B.n431 B.n30 585
R303 B.n30 B.n29 585
R304 B.n430 B.n429 585
R305 B.n429 B.n428 585
R306 B.n32 B.n31 585
R307 B.n427 B.n32 585
R308 B.n425 B.n424 585
R309 B.n426 B.n425 585
R310 B.n423 B.n37 585
R311 B.n37 B.n36 585
R312 B.n422 B.n421 585
R313 B.n421 B.n420 585
R314 B.n39 B.n38 585
R315 B.n419 B.n39 585
R316 B.n417 B.n416 585
R317 B.n418 B.n417 585
R318 B.n415 B.n44 585
R319 B.n44 B.n43 585
R320 B.n414 B.n413 585
R321 B.n413 B.n412 585
R322 B.n46 B.n45 585
R323 B.n411 B.n46 585
R324 B.n409 B.n408 585
R325 B.n410 B.n409 585
R326 B.n407 B.n51 585
R327 B.n51 B.n50 585
R328 B.n406 B.n405 585
R329 B.n405 B.n404 585
R330 B.n53 B.n52 585
R331 B.n403 B.n53 585
R332 B.n401 B.n400 585
R333 B.n402 B.n401 585
R334 B.n399 B.n58 585
R335 B.n58 B.n57 585
R336 B.n462 B.n461 585
R337 B.n461 B.n460 585
R338 B.n260 B.n187 458.866
R339 B.n397 B.n58 458.866
R340 B.n208 B.n185 458.866
R341 B.n394 B.n74 458.866
R342 B.n206 B.t11 286.036
R343 B.n203 B.t14 286.036
R344 B.n78 B.t16 286.036
R345 B.n75 B.t6 286.036
R346 B.n395 B.n72 256.663
R347 B.n395 B.n71 256.663
R348 B.n395 B.n70 256.663
R349 B.n395 B.n69 256.663
R350 B.n395 B.n68 256.663
R351 B.n395 B.n67 256.663
R352 B.n395 B.n66 256.663
R353 B.n395 B.n65 256.663
R354 B.n395 B.n64 256.663
R355 B.n395 B.n63 256.663
R356 B.n395 B.n62 256.663
R357 B.n395 B.n61 256.663
R358 B.n396 B.n395 256.663
R359 B.n259 B.n258 256.663
R360 B.n258 B.n190 256.663
R361 B.n258 B.n191 256.663
R362 B.n258 B.n192 256.663
R363 B.n258 B.n193 256.663
R364 B.n258 B.n194 256.663
R365 B.n258 B.n195 256.663
R366 B.n258 B.n196 256.663
R367 B.n258 B.n197 256.663
R368 B.n258 B.n198 256.663
R369 B.n258 B.n199 256.663
R370 B.n258 B.n200 256.663
R371 B.n258 B.n201 256.663
R372 B.n207 B.t10 235.805
R373 B.n204 B.t13 235.805
R374 B.n79 B.t17 235.805
R375 B.n76 B.t7 235.805
R376 B.n258 B.n186 221.28
R377 B.n395 B.n57 221.28
R378 B.n206 B.t8 208.733
R379 B.n203 B.t12 208.733
R380 B.n78 B.t15 208.733
R381 B.n75 B.t4 208.733
R382 B.n264 B.n187 163.367
R383 B.n264 B.n181 163.367
R384 B.n272 B.n181 163.367
R385 B.n272 B.n179 163.367
R386 B.n276 B.n179 163.367
R387 B.n276 B.n173 163.367
R388 B.n284 B.n173 163.367
R389 B.n284 B.n171 163.367
R390 B.n288 B.n171 163.367
R391 B.n288 B.n165 163.367
R392 B.n296 B.n165 163.367
R393 B.n296 B.n163 163.367
R394 B.n300 B.n163 163.367
R395 B.n300 B.n157 163.367
R396 B.n308 B.n157 163.367
R397 B.n308 B.n155 163.367
R398 B.n312 B.n155 163.367
R399 B.n312 B.n149 163.367
R400 B.n320 B.n149 163.367
R401 B.n320 B.n147 163.367
R402 B.n324 B.n147 163.367
R403 B.n324 B.n141 163.367
R404 B.n332 B.n141 163.367
R405 B.n332 B.n139 163.367
R406 B.n336 B.n139 163.367
R407 B.n336 B.n133 163.367
R408 B.n345 B.n133 163.367
R409 B.n345 B.n131 163.367
R410 B.n349 B.n131 163.367
R411 B.n349 B.n2 163.367
R412 B.n461 B.n2 163.367
R413 B.n461 B.n3 163.367
R414 B.n457 B.n3 163.367
R415 B.n457 B.n9 163.367
R416 B.n453 B.n9 163.367
R417 B.n453 B.n11 163.367
R418 B.n449 B.n11 163.367
R419 B.n449 B.n16 163.367
R420 B.n445 B.n16 163.367
R421 B.n445 B.n18 163.367
R422 B.n441 B.n18 163.367
R423 B.n441 B.n23 163.367
R424 B.n437 B.n23 163.367
R425 B.n437 B.n25 163.367
R426 B.n433 B.n25 163.367
R427 B.n433 B.n30 163.367
R428 B.n429 B.n30 163.367
R429 B.n429 B.n32 163.367
R430 B.n425 B.n32 163.367
R431 B.n425 B.n37 163.367
R432 B.n421 B.n37 163.367
R433 B.n421 B.n39 163.367
R434 B.n417 B.n39 163.367
R435 B.n417 B.n44 163.367
R436 B.n413 B.n44 163.367
R437 B.n413 B.n46 163.367
R438 B.n409 B.n46 163.367
R439 B.n409 B.n51 163.367
R440 B.n405 B.n51 163.367
R441 B.n405 B.n53 163.367
R442 B.n401 B.n53 163.367
R443 B.n401 B.n58 163.367
R444 B.n257 B.n189 163.367
R445 B.n257 B.n202 163.367
R446 B.n253 B.n252 163.367
R447 B.n249 B.n248 163.367
R448 B.n245 B.n244 163.367
R449 B.n241 B.n240 163.367
R450 B.n237 B.n236 163.367
R451 B.n233 B.n232 163.367
R452 B.n229 B.n228 163.367
R453 B.n224 B.n223 163.367
R454 B.n220 B.n219 163.367
R455 B.n216 B.n215 163.367
R456 B.n212 B.n211 163.367
R457 B.n266 B.n185 163.367
R458 B.n266 B.n183 163.367
R459 B.n270 B.n183 163.367
R460 B.n270 B.n177 163.367
R461 B.n278 B.n177 163.367
R462 B.n278 B.n175 163.367
R463 B.n282 B.n175 163.367
R464 B.n282 B.n169 163.367
R465 B.n290 B.n169 163.367
R466 B.n290 B.n167 163.367
R467 B.n294 B.n167 163.367
R468 B.n294 B.n161 163.367
R469 B.n302 B.n161 163.367
R470 B.n302 B.n159 163.367
R471 B.n306 B.n159 163.367
R472 B.n306 B.n153 163.367
R473 B.n314 B.n153 163.367
R474 B.n314 B.n151 163.367
R475 B.n318 B.n151 163.367
R476 B.n318 B.n145 163.367
R477 B.n326 B.n145 163.367
R478 B.n326 B.n143 163.367
R479 B.n330 B.n143 163.367
R480 B.n330 B.n137 163.367
R481 B.n338 B.n137 163.367
R482 B.n338 B.n135 163.367
R483 B.n343 B.n135 163.367
R484 B.n343 B.n129 163.367
R485 B.n351 B.n129 163.367
R486 B.n352 B.n351 163.367
R487 B.n352 B.n5 163.367
R488 B.n6 B.n5 163.367
R489 B.n7 B.n6 163.367
R490 B.n357 B.n7 163.367
R491 B.n357 B.n12 163.367
R492 B.n13 B.n12 163.367
R493 B.n14 B.n13 163.367
R494 B.n362 B.n14 163.367
R495 B.n362 B.n19 163.367
R496 B.n20 B.n19 163.367
R497 B.n21 B.n20 163.367
R498 B.n367 B.n21 163.367
R499 B.n367 B.n26 163.367
R500 B.n27 B.n26 163.367
R501 B.n28 B.n27 163.367
R502 B.n372 B.n28 163.367
R503 B.n372 B.n33 163.367
R504 B.n34 B.n33 163.367
R505 B.n35 B.n34 163.367
R506 B.n377 B.n35 163.367
R507 B.n377 B.n40 163.367
R508 B.n41 B.n40 163.367
R509 B.n42 B.n41 163.367
R510 B.n382 B.n42 163.367
R511 B.n382 B.n47 163.367
R512 B.n48 B.n47 163.367
R513 B.n49 B.n48 163.367
R514 B.n387 B.n49 163.367
R515 B.n387 B.n54 163.367
R516 B.n55 B.n54 163.367
R517 B.n56 B.n55 163.367
R518 B.n74 B.n56 163.367
R519 B.n80 B.n60 163.367
R520 B.n84 B.n83 163.367
R521 B.n88 B.n87 163.367
R522 B.n92 B.n91 163.367
R523 B.n97 B.n96 163.367
R524 B.n101 B.n100 163.367
R525 B.n105 B.n104 163.367
R526 B.n109 B.n108 163.367
R527 B.n113 B.n112 163.367
R528 B.n117 B.n116 163.367
R529 B.n121 B.n120 163.367
R530 B.n125 B.n124 163.367
R531 B.n394 B.n73 163.367
R532 B.n265 B.n186 124.356
R533 B.n265 B.n182 124.356
R534 B.n271 B.n182 124.356
R535 B.n271 B.n178 124.356
R536 B.n277 B.n178 124.356
R537 B.n277 B.n174 124.356
R538 B.n283 B.n174 124.356
R539 B.n289 B.n170 124.356
R540 B.n289 B.n166 124.356
R541 B.n295 B.n166 124.356
R542 B.n295 B.n162 124.356
R543 B.n301 B.n162 124.356
R544 B.n301 B.n158 124.356
R545 B.n307 B.n158 124.356
R546 B.n307 B.n154 124.356
R547 B.n313 B.n154 124.356
R548 B.n319 B.n150 124.356
R549 B.n319 B.n146 124.356
R550 B.n325 B.n146 124.356
R551 B.n325 B.n142 124.356
R552 B.n331 B.n142 124.356
R553 B.n331 B.n138 124.356
R554 B.n337 B.n138 124.356
R555 B.n344 B.n134 124.356
R556 B.n344 B.n130 124.356
R557 B.n350 B.n130 124.356
R558 B.n350 B.n4 124.356
R559 B.n460 B.n4 124.356
R560 B.n460 B.n459 124.356
R561 B.n459 B.n458 124.356
R562 B.n458 B.n8 124.356
R563 B.n452 B.n8 124.356
R564 B.n452 B.n451 124.356
R565 B.n450 B.n15 124.356
R566 B.n444 B.n15 124.356
R567 B.n444 B.n443 124.356
R568 B.n443 B.n442 124.356
R569 B.n442 B.n22 124.356
R570 B.n436 B.n22 124.356
R571 B.n436 B.n435 124.356
R572 B.n434 B.n29 124.356
R573 B.n428 B.n29 124.356
R574 B.n428 B.n427 124.356
R575 B.n427 B.n426 124.356
R576 B.n426 B.n36 124.356
R577 B.n420 B.n36 124.356
R578 B.n420 B.n419 124.356
R579 B.n419 B.n418 124.356
R580 B.n418 B.n43 124.356
R581 B.n412 B.n411 124.356
R582 B.n411 B.n410 124.356
R583 B.n410 B.n50 124.356
R584 B.n404 B.n50 124.356
R585 B.n404 B.n403 124.356
R586 B.n403 B.n402 124.356
R587 B.n402 B.n57 124.356
R588 B.n313 B.t3 120.698
R589 B.t2 B.n434 120.698
R590 B.t9 B.n170 106.069
R591 B.t5 B.n43 106.069
R592 B.n337 B.t1 73.151
R593 B.t0 B.n450 73.151
R594 B.n260 B.n259 71.676
R595 B.n202 B.n190 71.676
R596 B.n252 B.n191 71.676
R597 B.n248 B.n192 71.676
R598 B.n244 B.n193 71.676
R599 B.n240 B.n194 71.676
R600 B.n236 B.n195 71.676
R601 B.n232 B.n196 71.676
R602 B.n228 B.n197 71.676
R603 B.n223 B.n198 71.676
R604 B.n219 B.n199 71.676
R605 B.n215 B.n200 71.676
R606 B.n211 B.n201 71.676
R607 B.n397 B.n396 71.676
R608 B.n80 B.n61 71.676
R609 B.n84 B.n62 71.676
R610 B.n88 B.n63 71.676
R611 B.n92 B.n64 71.676
R612 B.n97 B.n65 71.676
R613 B.n101 B.n66 71.676
R614 B.n105 B.n67 71.676
R615 B.n109 B.n68 71.676
R616 B.n113 B.n69 71.676
R617 B.n117 B.n70 71.676
R618 B.n121 B.n71 71.676
R619 B.n125 B.n72 71.676
R620 B.n73 B.n72 71.676
R621 B.n124 B.n71 71.676
R622 B.n120 B.n70 71.676
R623 B.n116 B.n69 71.676
R624 B.n112 B.n68 71.676
R625 B.n108 B.n67 71.676
R626 B.n104 B.n66 71.676
R627 B.n100 B.n65 71.676
R628 B.n96 B.n64 71.676
R629 B.n91 B.n63 71.676
R630 B.n87 B.n62 71.676
R631 B.n83 B.n61 71.676
R632 B.n396 B.n60 71.676
R633 B.n259 B.n189 71.676
R634 B.n253 B.n190 71.676
R635 B.n249 B.n191 71.676
R636 B.n245 B.n192 71.676
R637 B.n241 B.n193 71.676
R638 B.n237 B.n194 71.676
R639 B.n233 B.n195 71.676
R640 B.n229 B.n196 71.676
R641 B.n224 B.n197 71.676
R642 B.n220 B.n198 71.676
R643 B.n216 B.n199 71.676
R644 B.n212 B.n200 71.676
R645 B.n208 B.n201 71.676
R646 B.n226 B.n207 59.5399
R647 B.n205 B.n204 59.5399
R648 B.n94 B.n79 59.5399
R649 B.n77 B.n76 59.5399
R650 B.t1 B.n134 51.2058
R651 B.n451 B.t0 51.2058
R652 B.n207 B.n206 50.2308
R653 B.n204 B.n203 50.2308
R654 B.n79 B.n78 50.2308
R655 B.n76 B.n75 50.2308
R656 B.n393 B.n392 29.8151
R657 B.n399 B.n398 29.8151
R658 B.n209 B.n184 29.8151
R659 B.n262 B.n261 29.8151
R660 B.n283 B.t9 18.2881
R661 B.n412 B.t5 18.2881
R662 B B.n462 18.0485
R663 B.n398 B.n59 10.6151
R664 B.n81 B.n59 10.6151
R665 B.n82 B.n81 10.6151
R666 B.n85 B.n82 10.6151
R667 B.n86 B.n85 10.6151
R668 B.n89 B.n86 10.6151
R669 B.n90 B.n89 10.6151
R670 B.n93 B.n90 10.6151
R671 B.n98 B.n95 10.6151
R672 B.n99 B.n98 10.6151
R673 B.n102 B.n99 10.6151
R674 B.n103 B.n102 10.6151
R675 B.n106 B.n103 10.6151
R676 B.n107 B.n106 10.6151
R677 B.n110 B.n107 10.6151
R678 B.n111 B.n110 10.6151
R679 B.n115 B.n114 10.6151
R680 B.n118 B.n115 10.6151
R681 B.n119 B.n118 10.6151
R682 B.n122 B.n119 10.6151
R683 B.n123 B.n122 10.6151
R684 B.n126 B.n123 10.6151
R685 B.n127 B.n126 10.6151
R686 B.n393 B.n127 10.6151
R687 B.n267 B.n184 10.6151
R688 B.n268 B.n267 10.6151
R689 B.n269 B.n268 10.6151
R690 B.n269 B.n176 10.6151
R691 B.n279 B.n176 10.6151
R692 B.n280 B.n279 10.6151
R693 B.n281 B.n280 10.6151
R694 B.n281 B.n168 10.6151
R695 B.n291 B.n168 10.6151
R696 B.n292 B.n291 10.6151
R697 B.n293 B.n292 10.6151
R698 B.n293 B.n160 10.6151
R699 B.n303 B.n160 10.6151
R700 B.n304 B.n303 10.6151
R701 B.n305 B.n304 10.6151
R702 B.n305 B.n152 10.6151
R703 B.n315 B.n152 10.6151
R704 B.n316 B.n315 10.6151
R705 B.n317 B.n316 10.6151
R706 B.n317 B.n144 10.6151
R707 B.n327 B.n144 10.6151
R708 B.n328 B.n327 10.6151
R709 B.n329 B.n328 10.6151
R710 B.n329 B.n136 10.6151
R711 B.n339 B.n136 10.6151
R712 B.n340 B.n339 10.6151
R713 B.n342 B.n340 10.6151
R714 B.n342 B.n341 10.6151
R715 B.n341 B.n128 10.6151
R716 B.n353 B.n128 10.6151
R717 B.n354 B.n353 10.6151
R718 B.n355 B.n354 10.6151
R719 B.n356 B.n355 10.6151
R720 B.n358 B.n356 10.6151
R721 B.n359 B.n358 10.6151
R722 B.n360 B.n359 10.6151
R723 B.n361 B.n360 10.6151
R724 B.n363 B.n361 10.6151
R725 B.n364 B.n363 10.6151
R726 B.n365 B.n364 10.6151
R727 B.n366 B.n365 10.6151
R728 B.n368 B.n366 10.6151
R729 B.n369 B.n368 10.6151
R730 B.n370 B.n369 10.6151
R731 B.n371 B.n370 10.6151
R732 B.n373 B.n371 10.6151
R733 B.n374 B.n373 10.6151
R734 B.n375 B.n374 10.6151
R735 B.n376 B.n375 10.6151
R736 B.n378 B.n376 10.6151
R737 B.n379 B.n378 10.6151
R738 B.n380 B.n379 10.6151
R739 B.n381 B.n380 10.6151
R740 B.n383 B.n381 10.6151
R741 B.n384 B.n383 10.6151
R742 B.n385 B.n384 10.6151
R743 B.n386 B.n385 10.6151
R744 B.n388 B.n386 10.6151
R745 B.n389 B.n388 10.6151
R746 B.n390 B.n389 10.6151
R747 B.n391 B.n390 10.6151
R748 B.n392 B.n391 10.6151
R749 B.n261 B.n188 10.6151
R750 B.n256 B.n188 10.6151
R751 B.n256 B.n255 10.6151
R752 B.n255 B.n254 10.6151
R753 B.n254 B.n251 10.6151
R754 B.n251 B.n250 10.6151
R755 B.n250 B.n247 10.6151
R756 B.n247 B.n246 10.6151
R757 B.n243 B.n242 10.6151
R758 B.n242 B.n239 10.6151
R759 B.n239 B.n238 10.6151
R760 B.n238 B.n235 10.6151
R761 B.n235 B.n234 10.6151
R762 B.n234 B.n231 10.6151
R763 B.n231 B.n230 10.6151
R764 B.n230 B.n227 10.6151
R765 B.n225 B.n222 10.6151
R766 B.n222 B.n221 10.6151
R767 B.n221 B.n218 10.6151
R768 B.n218 B.n217 10.6151
R769 B.n217 B.n214 10.6151
R770 B.n214 B.n213 10.6151
R771 B.n213 B.n210 10.6151
R772 B.n210 B.n209 10.6151
R773 B.n263 B.n262 10.6151
R774 B.n263 B.n180 10.6151
R775 B.n273 B.n180 10.6151
R776 B.n274 B.n273 10.6151
R777 B.n275 B.n274 10.6151
R778 B.n275 B.n172 10.6151
R779 B.n285 B.n172 10.6151
R780 B.n286 B.n285 10.6151
R781 B.n287 B.n286 10.6151
R782 B.n287 B.n164 10.6151
R783 B.n297 B.n164 10.6151
R784 B.n298 B.n297 10.6151
R785 B.n299 B.n298 10.6151
R786 B.n299 B.n156 10.6151
R787 B.n309 B.n156 10.6151
R788 B.n310 B.n309 10.6151
R789 B.n311 B.n310 10.6151
R790 B.n311 B.n148 10.6151
R791 B.n321 B.n148 10.6151
R792 B.n322 B.n321 10.6151
R793 B.n323 B.n322 10.6151
R794 B.n323 B.n140 10.6151
R795 B.n333 B.n140 10.6151
R796 B.n334 B.n333 10.6151
R797 B.n335 B.n334 10.6151
R798 B.n335 B.n132 10.6151
R799 B.n346 B.n132 10.6151
R800 B.n347 B.n346 10.6151
R801 B.n348 B.n347 10.6151
R802 B.n348 B.n0 10.6151
R803 B.n456 B.n1 10.6151
R804 B.n456 B.n455 10.6151
R805 B.n455 B.n454 10.6151
R806 B.n454 B.n10 10.6151
R807 B.n448 B.n10 10.6151
R808 B.n448 B.n447 10.6151
R809 B.n447 B.n446 10.6151
R810 B.n446 B.n17 10.6151
R811 B.n440 B.n17 10.6151
R812 B.n440 B.n439 10.6151
R813 B.n439 B.n438 10.6151
R814 B.n438 B.n24 10.6151
R815 B.n432 B.n24 10.6151
R816 B.n432 B.n431 10.6151
R817 B.n431 B.n430 10.6151
R818 B.n430 B.n31 10.6151
R819 B.n424 B.n31 10.6151
R820 B.n424 B.n423 10.6151
R821 B.n423 B.n422 10.6151
R822 B.n422 B.n38 10.6151
R823 B.n416 B.n38 10.6151
R824 B.n416 B.n415 10.6151
R825 B.n415 B.n414 10.6151
R826 B.n414 B.n45 10.6151
R827 B.n408 B.n45 10.6151
R828 B.n408 B.n407 10.6151
R829 B.n407 B.n406 10.6151
R830 B.n406 B.n52 10.6151
R831 B.n400 B.n52 10.6151
R832 B.n400 B.n399 10.6151
R833 B.n95 B.n94 6.5566
R834 B.n111 B.n77 6.5566
R835 B.n243 B.n205 6.5566
R836 B.n227 B.n226 6.5566
R837 B.n94 B.n93 4.05904
R838 B.n114 B.n77 4.05904
R839 B.n246 B.n205 4.05904
R840 B.n226 B.n225 4.05904
R841 B.t3 B.n150 3.65802
R842 B.n435 B.t2 3.65802
R843 B.n462 B.n0 2.81026
R844 B.n462 B.n1 2.81026
R845 VP.n12 VP.n0 161.3
R846 VP.n11 VP.n10 161.3
R847 VP.n9 VP.n1 161.3
R848 VP.n8 VP.n7 161.3
R849 VP.n6 VP.n2 161.3
R850 VP.n5 VP.n4 96.3991
R851 VP.n14 VP.n13 96.3991
R852 VP.n3 VP.t2 44.0585
R853 VP.n3 VP.t1 43.4112
R854 VP.n4 VP.n3 42.3632
R855 VP.n7 VP.n1 40.577
R856 VP.n11 VP.n1 40.577
R857 VP.n7 VP.n6 24.5923
R858 VP.n12 VP.n11 24.5923
R859 VP.n6 VP.n5 14.5097
R860 VP.n13 VP.n12 14.5097
R861 VP.n5 VP.t0 7.89165
R862 VP.n13 VP.t3 7.89165
R863 VP.n4 VP.n2 0.278335
R864 VP.n14 VP.n0 0.278335
R865 VP.n8 VP.n2 0.189894
R866 VP.n9 VP.n8 0.189894
R867 VP.n10 VP.n9 0.189894
R868 VP.n10 VP.n0 0.189894
R869 VP VP.n14 0.153485
R870 VDD1 VDD1.n1 268.156
R871 VDD1 VDD1.n0 236.637
R872 VDD1.n0 VDD1.t1 26.7573
R873 VDD1.n0 VDD1.t2 26.7573
R874 VDD1.n1 VDD1.t3 26.7573
R875 VDD1.n1 VDD1.t0 26.7573
C0 VP VN 3.86761f
C1 VDD2 VTAIL 2.59309f
C2 VDD1 VTAIL 2.54117f
C3 VTAIL VP 1.25455f
C4 VTAIL VN 1.24044f
C5 VDD2 VDD1 0.947428f
C6 VDD2 VP 0.38183f
C7 VDD1 VP 0.817578f
C8 VDD2 VN 0.594445f
C9 VDD1 VN 0.156305f
C10 VDD2 B 2.669709f
C11 VDD1 B 5.023839f
C12 VTAIL B 2.724209f
C13 VN B 8.7191f
C14 VP B 7.188066f
C15 VDD1.t1 B 0.014088f
C16 VDD1.t2 B 0.014088f
C17 VDD1.n0 B 0.034519f
C18 VDD1.t3 B 0.014088f
C19 VDD1.t0 B 0.014088f
C20 VDD1.n1 B 0.122005f
C21 VP.n0 B 0.038564f
C22 VP.t3 B 0.075344f
C23 VP.n1 B 0.023626f
C24 VP.n2 B 0.038564f
C25 VP.t0 B 0.075344f
C26 VP.t1 B 0.269866f
C27 VP.t2 B 0.273379f
C28 VP.n3 B 1.23387f
C29 VP.n4 B 1.17845f
C30 VP.n5 B 0.163615f
C31 VP.n6 B 0.043266f
C32 VP.n7 B 0.057832f
C33 VP.n8 B 0.029252f
C34 VP.n9 B 0.029252f
C35 VP.n10 B 0.029252f
C36 VP.n11 B 0.057832f
C37 VP.n12 B 0.043266f
C38 VP.n13 B 0.163615f
C39 VP.n14 B 0.041391f
C40 VDD2.t1 B 0.015193f
C41 VDD2.t3 B 0.015193f
C42 VDD2.n0 B 0.124037f
C43 VDD2.t2 B 0.015193f
C44 VDD2.t0 B 0.015193f
C45 VDD2.n1 B 0.037158f
C46 VDD2.n2 B 2.18552f
C47 VTAIL.t6 B 0.070218f
C48 VTAIL.n0 B 0.187246f
C49 VTAIL.t1 B 0.070218f
C50 VTAIL.n1 B 0.279346f
C51 VTAIL.t3 B 0.070218f
C52 VTAIL.n2 B 0.855218f
C53 VTAIL.t5 B 0.070218f
C54 VTAIL.n3 B 0.855218f
C55 VTAIL.t4 B 0.070218f
C56 VTAIL.n4 B 0.279346f
C57 VTAIL.t0 B 0.070218f
C58 VTAIL.n5 B 0.279346f
C59 VTAIL.t2 B 0.070218f
C60 VTAIL.n6 B 0.855218f
C61 VTAIL.t7 B 0.070218f
C62 VTAIL.n7 B 0.752989f
C63 VN.t2 B 0.270527f
C64 VN.t0 B 0.26705f
C65 VN.n0 B 0.178097f
C66 VN.t3 B 0.270527f
C67 VN.t1 B 0.26705f
C68 VN.n1 B 1.23634f
.ends

