* NGSPICE file created from diff_pair_sample_1568.ext - technology: sky130A

.subckt diff_pair_sample_1568 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t18 VP.t0 VDD1.t4 w_n2842_n4408# sky130_fd_pr__pfet_01v8 ad=2.838 pd=17.53 as=2.838 ps=17.53 w=17.2 l=1.23
X1 VDD2.t9 VN.t0 VTAIL.t2 w_n2842_n4408# sky130_fd_pr__pfet_01v8 ad=2.838 pd=17.53 as=6.708 ps=35.18 w=17.2 l=1.23
X2 VTAIL.t19 VN.t1 VDD2.t8 w_n2842_n4408# sky130_fd_pr__pfet_01v8 ad=2.838 pd=17.53 as=2.838 ps=17.53 w=17.2 l=1.23
X3 VDD1.t7 VP.t1 VTAIL.t17 w_n2842_n4408# sky130_fd_pr__pfet_01v8 ad=2.838 pd=17.53 as=6.708 ps=35.18 w=17.2 l=1.23
X4 B.t11 B.t9 B.t10 w_n2842_n4408# sky130_fd_pr__pfet_01v8 ad=6.708 pd=35.18 as=0 ps=0 w=17.2 l=1.23
X5 VTAIL.t1 VN.t2 VDD2.t7 w_n2842_n4408# sky130_fd_pr__pfet_01v8 ad=2.838 pd=17.53 as=2.838 ps=17.53 w=17.2 l=1.23
X6 VDD1.t6 VP.t2 VTAIL.t16 w_n2842_n4408# sky130_fd_pr__pfet_01v8 ad=6.708 pd=35.18 as=2.838 ps=17.53 w=17.2 l=1.23
X7 VDD2.t6 VN.t3 VTAIL.t5 w_n2842_n4408# sky130_fd_pr__pfet_01v8 ad=6.708 pd=35.18 as=2.838 ps=17.53 w=17.2 l=1.23
X8 B.t8 B.t6 B.t7 w_n2842_n4408# sky130_fd_pr__pfet_01v8 ad=6.708 pd=35.18 as=0 ps=0 w=17.2 l=1.23
X9 VDD1.t1 VP.t3 VTAIL.t15 w_n2842_n4408# sky130_fd_pr__pfet_01v8 ad=2.838 pd=17.53 as=2.838 ps=17.53 w=17.2 l=1.23
X10 VDD2.t5 VN.t4 VTAIL.t6 w_n2842_n4408# sky130_fd_pr__pfet_01v8 ad=2.838 pd=17.53 as=2.838 ps=17.53 w=17.2 l=1.23
X11 VTAIL.t3 VN.t5 VDD2.t4 w_n2842_n4408# sky130_fd_pr__pfet_01v8 ad=2.838 pd=17.53 as=2.838 ps=17.53 w=17.2 l=1.23
X12 VDD2.t3 VN.t6 VTAIL.t4 w_n2842_n4408# sky130_fd_pr__pfet_01v8 ad=2.838 pd=17.53 as=6.708 ps=35.18 w=17.2 l=1.23
X13 B.t5 B.t3 B.t4 w_n2842_n4408# sky130_fd_pr__pfet_01v8 ad=6.708 pd=35.18 as=0 ps=0 w=17.2 l=1.23
X14 VTAIL.t14 VP.t4 VDD1.t0 w_n2842_n4408# sky130_fd_pr__pfet_01v8 ad=2.838 pd=17.53 as=2.838 ps=17.53 w=17.2 l=1.23
X15 VDD2.t2 VN.t7 VTAIL.t7 w_n2842_n4408# sky130_fd_pr__pfet_01v8 ad=6.708 pd=35.18 as=2.838 ps=17.53 w=17.2 l=1.23
X16 VTAIL.t8 VN.t8 VDD2.t1 w_n2842_n4408# sky130_fd_pr__pfet_01v8 ad=2.838 pd=17.53 as=2.838 ps=17.53 w=17.2 l=1.23
X17 VTAIL.t13 VP.t5 VDD1.t3 w_n2842_n4408# sky130_fd_pr__pfet_01v8 ad=2.838 pd=17.53 as=2.838 ps=17.53 w=17.2 l=1.23
X18 VDD1.t2 VP.t6 VTAIL.t12 w_n2842_n4408# sky130_fd_pr__pfet_01v8 ad=2.838 pd=17.53 as=6.708 ps=35.18 w=17.2 l=1.23
X19 VDD1.t9 VP.t7 VTAIL.t11 w_n2842_n4408# sky130_fd_pr__pfet_01v8 ad=6.708 pd=35.18 as=2.838 ps=17.53 w=17.2 l=1.23
X20 VDD2.t0 VN.t9 VTAIL.t0 w_n2842_n4408# sky130_fd_pr__pfet_01v8 ad=2.838 pd=17.53 as=2.838 ps=17.53 w=17.2 l=1.23
X21 B.t2 B.t0 B.t1 w_n2842_n4408# sky130_fd_pr__pfet_01v8 ad=6.708 pd=35.18 as=0 ps=0 w=17.2 l=1.23
X22 VDD1.t8 VP.t8 VTAIL.t10 w_n2842_n4408# sky130_fd_pr__pfet_01v8 ad=2.838 pd=17.53 as=2.838 ps=17.53 w=17.2 l=1.23
X23 VTAIL.t9 VP.t9 VDD1.t5 w_n2842_n4408# sky130_fd_pr__pfet_01v8 ad=2.838 pd=17.53 as=2.838 ps=17.53 w=17.2 l=1.23
R0 VP.n13 VP.t7 389.293
R1 VP.n30 VP.t2 368.947
R2 VP.n47 VP.t1 368.947
R3 VP.n27 VP.t6 368.947
R4 VP.n5 VP.t5 337.009
R5 VP.n3 VP.t8 337.009
R6 VP.n1 VP.t0 337.009
R7 VP.n8 VP.t4 337.009
R8 VP.n10 VP.t3 337.009
R9 VP.n12 VP.t9 337.009
R10 VP.n15 VP.n14 161.3
R11 VP.n16 VP.n11 161.3
R12 VP.n18 VP.n17 161.3
R13 VP.n20 VP.n19 161.3
R14 VP.n21 VP.n9 161.3
R15 VP.n23 VP.n22 161.3
R16 VP.n25 VP.n24 161.3
R17 VP.n26 VP.n7 161.3
R18 VP.n46 VP.n0 161.3
R19 VP.n45 VP.n44 161.3
R20 VP.n43 VP.n42 161.3
R21 VP.n41 VP.n2 161.3
R22 VP.n40 VP.n39 161.3
R23 VP.n38 VP.n37 161.3
R24 VP.n36 VP.n4 161.3
R25 VP.n35 VP.n34 161.3
R26 VP.n33 VP.n32 161.3
R27 VP.n31 VP.n6 161.3
R28 VP.n28 VP.n27 80.6037
R29 VP.n48 VP.n47 80.6037
R30 VP.n30 VP.n29 80.6037
R31 VP.n29 VP.n28 49.7817
R32 VP.n36 VP.n35 43.4833
R33 VP.n42 VP.n41 43.4833
R34 VP.n22 VP.n21 43.4833
R35 VP.n16 VP.n15 43.4833
R36 VP.n13 VP.n12 42.2534
R37 VP.n37 VP.n36 37.6707
R38 VP.n41 VP.n40 37.6707
R39 VP.n21 VP.n20 37.6707
R40 VP.n17 VP.n16 37.6707
R41 VP.n31 VP.n30 37.246
R42 VP.n47 VP.n46 37.246
R43 VP.n27 VP.n26 37.246
R44 VP.n32 VP.n31 31.8581
R45 VP.n46 VP.n45 31.8581
R46 VP.n26 VP.n25 31.8581
R47 VP.n14 VP.n13 29.1038
R48 VP.n35 VP.n5 15.2474
R49 VP.n42 VP.n1 15.2474
R50 VP.n22 VP.n8 15.2474
R51 VP.n15 VP.n12 15.2474
R52 VP.n37 VP.n3 12.2964
R53 VP.n40 VP.n3 12.2964
R54 VP.n17 VP.n10 12.2964
R55 VP.n20 VP.n10 12.2964
R56 VP.n32 VP.n5 9.3454
R57 VP.n45 VP.n1 9.3454
R58 VP.n25 VP.n8 9.3454
R59 VP.n28 VP.n7 0.285035
R60 VP.n29 VP.n6 0.285035
R61 VP.n48 VP.n0 0.285035
R62 VP.n14 VP.n11 0.189894
R63 VP.n18 VP.n11 0.189894
R64 VP.n19 VP.n18 0.189894
R65 VP.n19 VP.n9 0.189894
R66 VP.n23 VP.n9 0.189894
R67 VP.n24 VP.n23 0.189894
R68 VP.n24 VP.n7 0.189894
R69 VP.n33 VP.n6 0.189894
R70 VP.n34 VP.n33 0.189894
R71 VP.n34 VP.n4 0.189894
R72 VP.n38 VP.n4 0.189894
R73 VP.n39 VP.n38 0.189894
R74 VP.n39 VP.n2 0.189894
R75 VP.n43 VP.n2 0.189894
R76 VP.n44 VP.n43 0.189894
R77 VP.n44 VP.n0 0.189894
R78 VP VP.n48 0.146778
R79 VDD1.n1 VDD1.t9 73.2125
R80 VDD1.n3 VDD1.t6 73.2124
R81 VDD1.n5 VDD1.n4 70.931
R82 VDD1.n1 VDD1.n0 69.978
R83 VDD1.n7 VDD1.n6 69.9778
R84 VDD1.n3 VDD1.n2 69.9777
R85 VDD1.n7 VDD1.n5 46.1862
R86 VDD1.n6 VDD1.t0 1.89033
R87 VDD1.n6 VDD1.t2 1.89033
R88 VDD1.n0 VDD1.t5 1.89033
R89 VDD1.n0 VDD1.t1 1.89033
R90 VDD1.n4 VDD1.t4 1.89033
R91 VDD1.n4 VDD1.t7 1.89033
R92 VDD1.n2 VDD1.t3 1.89033
R93 VDD1.n2 VDD1.t8 1.89033
R94 VDD1 VDD1.n7 0.950931
R95 VDD1 VDD1.n1 0.394897
R96 VDD1.n5 VDD1.n3 0.281361
R97 VTAIL.n11 VTAIL.t4 55.1889
R98 VTAIL.n17 VTAIL.t2 55.1888
R99 VTAIL.n2 VTAIL.t17 55.1888
R100 VTAIL.n16 VTAIL.t12 55.1888
R101 VTAIL.n15 VTAIL.n14 53.2992
R102 VTAIL.n13 VTAIL.n12 53.2992
R103 VTAIL.n10 VTAIL.n9 53.2992
R104 VTAIL.n8 VTAIL.n7 53.2992
R105 VTAIL.n19 VTAIL.n18 53.2989
R106 VTAIL.n1 VTAIL.n0 53.2989
R107 VTAIL.n4 VTAIL.n3 53.2989
R108 VTAIL.n6 VTAIL.n5 53.2989
R109 VTAIL.n8 VTAIL.n6 29.8841
R110 VTAIL.n17 VTAIL.n16 28.5393
R111 VTAIL.n18 VTAIL.t6 1.89033
R112 VTAIL.n18 VTAIL.t1 1.89033
R113 VTAIL.n0 VTAIL.t7 1.89033
R114 VTAIL.n0 VTAIL.t3 1.89033
R115 VTAIL.n3 VTAIL.t10 1.89033
R116 VTAIL.n3 VTAIL.t18 1.89033
R117 VTAIL.n5 VTAIL.t16 1.89033
R118 VTAIL.n5 VTAIL.t13 1.89033
R119 VTAIL.n14 VTAIL.t15 1.89033
R120 VTAIL.n14 VTAIL.t14 1.89033
R121 VTAIL.n12 VTAIL.t11 1.89033
R122 VTAIL.n12 VTAIL.t9 1.89033
R123 VTAIL.n9 VTAIL.t0 1.89033
R124 VTAIL.n9 VTAIL.t8 1.89033
R125 VTAIL.n7 VTAIL.t5 1.89033
R126 VTAIL.n7 VTAIL.t19 1.89033
R127 VTAIL.n10 VTAIL.n8 1.34533
R128 VTAIL.n11 VTAIL.n10 1.34533
R129 VTAIL.n15 VTAIL.n13 1.34533
R130 VTAIL.n16 VTAIL.n15 1.34533
R131 VTAIL.n6 VTAIL.n4 1.34533
R132 VTAIL.n4 VTAIL.n2 1.34533
R133 VTAIL.n19 VTAIL.n17 1.34533
R134 VTAIL.n13 VTAIL.n11 1.14274
R135 VTAIL.n2 VTAIL.n1 1.14274
R136 VTAIL VTAIL.n1 1.06731
R137 VTAIL VTAIL.n19 0.278517
R138 VN.n6 VN.t7 389.293
R139 VN.n28 VN.t6 389.293
R140 VN.n20 VN.t0 368.947
R141 VN.n42 VN.t3 368.947
R142 VN.n5 VN.t5 337.009
R143 VN.n3 VN.t4 337.009
R144 VN.n1 VN.t2 337.009
R145 VN.n27 VN.t8 337.009
R146 VN.n25 VN.t9 337.009
R147 VN.n23 VN.t1 337.009
R148 VN.n41 VN.n22 161.3
R149 VN.n40 VN.n39 161.3
R150 VN.n38 VN.n37 161.3
R151 VN.n36 VN.n24 161.3
R152 VN.n35 VN.n34 161.3
R153 VN.n33 VN.n32 161.3
R154 VN.n31 VN.n26 161.3
R155 VN.n30 VN.n29 161.3
R156 VN.n19 VN.n0 161.3
R157 VN.n18 VN.n17 161.3
R158 VN.n16 VN.n15 161.3
R159 VN.n14 VN.n2 161.3
R160 VN.n13 VN.n12 161.3
R161 VN.n11 VN.n10 161.3
R162 VN.n9 VN.n4 161.3
R163 VN.n8 VN.n7 161.3
R164 VN.n43 VN.n42 80.6037
R165 VN.n21 VN.n20 80.6037
R166 VN VN.n43 50.0672
R167 VN.n9 VN.n8 43.4833
R168 VN.n15 VN.n14 43.4833
R169 VN.n31 VN.n30 43.4833
R170 VN.n37 VN.n36 43.4833
R171 VN.n6 VN.n5 42.2534
R172 VN.n28 VN.n27 42.2534
R173 VN.n10 VN.n9 37.6707
R174 VN.n14 VN.n13 37.6707
R175 VN.n32 VN.n31 37.6707
R176 VN.n36 VN.n35 37.6707
R177 VN.n20 VN.n19 37.246
R178 VN.n42 VN.n41 37.246
R179 VN.n19 VN.n18 31.8581
R180 VN.n41 VN.n40 31.8581
R181 VN.n29 VN.n28 29.1038
R182 VN.n7 VN.n6 29.1038
R183 VN.n8 VN.n5 15.2474
R184 VN.n15 VN.n1 15.2474
R185 VN.n30 VN.n27 15.2474
R186 VN.n37 VN.n23 15.2474
R187 VN.n10 VN.n3 12.2964
R188 VN.n13 VN.n3 12.2964
R189 VN.n35 VN.n25 12.2964
R190 VN.n32 VN.n25 12.2964
R191 VN.n18 VN.n1 9.3454
R192 VN.n40 VN.n23 9.3454
R193 VN.n43 VN.n22 0.285035
R194 VN.n21 VN.n0 0.285035
R195 VN.n39 VN.n22 0.189894
R196 VN.n39 VN.n38 0.189894
R197 VN.n38 VN.n24 0.189894
R198 VN.n34 VN.n24 0.189894
R199 VN.n34 VN.n33 0.189894
R200 VN.n33 VN.n26 0.189894
R201 VN.n29 VN.n26 0.189894
R202 VN.n7 VN.n4 0.189894
R203 VN.n11 VN.n4 0.189894
R204 VN.n12 VN.n11 0.189894
R205 VN.n12 VN.n2 0.189894
R206 VN.n16 VN.n2 0.189894
R207 VN.n17 VN.n16 0.189894
R208 VN.n17 VN.n0 0.189894
R209 VN VN.n21 0.146778
R210 VDD2.n1 VDD2.t2 73.2124
R211 VDD2.n4 VDD2.t6 71.8677
R212 VDD2.n3 VDD2.n2 70.931
R213 VDD2 VDD2.n7 70.9282
R214 VDD2.n6 VDD2.n5 69.978
R215 VDD2.n1 VDD2.n0 69.9777
R216 VDD2.n4 VDD2.n3 44.9308
R217 VDD2.n7 VDD2.t1 1.89033
R218 VDD2.n7 VDD2.t3 1.89033
R219 VDD2.n5 VDD2.t8 1.89033
R220 VDD2.n5 VDD2.t0 1.89033
R221 VDD2.n2 VDD2.t7 1.89033
R222 VDD2.n2 VDD2.t9 1.89033
R223 VDD2.n0 VDD2.t4 1.89033
R224 VDD2.n0 VDD2.t5 1.89033
R225 VDD2.n6 VDD2.n4 1.34533
R226 VDD2 VDD2.n6 0.394897
R227 VDD2.n3 VDD2.n1 0.281361
R228 B.n441 B.n440 585
R229 B.n439 B.n122 585
R230 B.n438 B.n437 585
R231 B.n436 B.n123 585
R232 B.n435 B.n434 585
R233 B.n433 B.n124 585
R234 B.n432 B.n431 585
R235 B.n430 B.n125 585
R236 B.n429 B.n428 585
R237 B.n427 B.n126 585
R238 B.n426 B.n425 585
R239 B.n424 B.n127 585
R240 B.n423 B.n422 585
R241 B.n421 B.n128 585
R242 B.n420 B.n419 585
R243 B.n418 B.n129 585
R244 B.n417 B.n416 585
R245 B.n415 B.n130 585
R246 B.n414 B.n413 585
R247 B.n412 B.n131 585
R248 B.n411 B.n410 585
R249 B.n409 B.n132 585
R250 B.n408 B.n407 585
R251 B.n406 B.n133 585
R252 B.n405 B.n404 585
R253 B.n403 B.n134 585
R254 B.n402 B.n401 585
R255 B.n400 B.n135 585
R256 B.n399 B.n398 585
R257 B.n397 B.n136 585
R258 B.n396 B.n395 585
R259 B.n394 B.n137 585
R260 B.n393 B.n392 585
R261 B.n391 B.n138 585
R262 B.n390 B.n389 585
R263 B.n388 B.n139 585
R264 B.n387 B.n386 585
R265 B.n385 B.n140 585
R266 B.n384 B.n383 585
R267 B.n382 B.n141 585
R268 B.n381 B.n380 585
R269 B.n379 B.n142 585
R270 B.n378 B.n377 585
R271 B.n376 B.n143 585
R272 B.n375 B.n374 585
R273 B.n373 B.n144 585
R274 B.n372 B.n371 585
R275 B.n370 B.n145 585
R276 B.n369 B.n368 585
R277 B.n367 B.n146 585
R278 B.n366 B.n365 585
R279 B.n364 B.n147 585
R280 B.n363 B.n362 585
R281 B.n361 B.n148 585
R282 B.n360 B.n359 585
R283 B.n358 B.n149 585
R284 B.n357 B.n356 585
R285 B.n355 B.n354 585
R286 B.n353 B.n153 585
R287 B.n352 B.n351 585
R288 B.n350 B.n154 585
R289 B.n349 B.n348 585
R290 B.n347 B.n155 585
R291 B.n346 B.n345 585
R292 B.n344 B.n156 585
R293 B.n343 B.n342 585
R294 B.n340 B.n157 585
R295 B.n339 B.n338 585
R296 B.n337 B.n160 585
R297 B.n336 B.n335 585
R298 B.n334 B.n161 585
R299 B.n333 B.n332 585
R300 B.n331 B.n162 585
R301 B.n330 B.n329 585
R302 B.n328 B.n163 585
R303 B.n327 B.n326 585
R304 B.n325 B.n164 585
R305 B.n324 B.n323 585
R306 B.n322 B.n165 585
R307 B.n321 B.n320 585
R308 B.n319 B.n166 585
R309 B.n318 B.n317 585
R310 B.n316 B.n167 585
R311 B.n315 B.n314 585
R312 B.n313 B.n168 585
R313 B.n312 B.n311 585
R314 B.n310 B.n169 585
R315 B.n309 B.n308 585
R316 B.n307 B.n170 585
R317 B.n306 B.n305 585
R318 B.n304 B.n171 585
R319 B.n303 B.n302 585
R320 B.n301 B.n172 585
R321 B.n300 B.n299 585
R322 B.n298 B.n173 585
R323 B.n297 B.n296 585
R324 B.n295 B.n174 585
R325 B.n294 B.n293 585
R326 B.n292 B.n175 585
R327 B.n291 B.n290 585
R328 B.n289 B.n176 585
R329 B.n288 B.n287 585
R330 B.n286 B.n177 585
R331 B.n285 B.n284 585
R332 B.n283 B.n178 585
R333 B.n282 B.n281 585
R334 B.n280 B.n179 585
R335 B.n279 B.n278 585
R336 B.n277 B.n180 585
R337 B.n276 B.n275 585
R338 B.n274 B.n181 585
R339 B.n273 B.n272 585
R340 B.n271 B.n182 585
R341 B.n270 B.n269 585
R342 B.n268 B.n183 585
R343 B.n267 B.n266 585
R344 B.n265 B.n184 585
R345 B.n264 B.n263 585
R346 B.n262 B.n185 585
R347 B.n261 B.n260 585
R348 B.n259 B.n186 585
R349 B.n258 B.n257 585
R350 B.n256 B.n187 585
R351 B.n442 B.n121 585
R352 B.n444 B.n443 585
R353 B.n445 B.n120 585
R354 B.n447 B.n446 585
R355 B.n448 B.n119 585
R356 B.n450 B.n449 585
R357 B.n451 B.n118 585
R358 B.n453 B.n452 585
R359 B.n454 B.n117 585
R360 B.n456 B.n455 585
R361 B.n457 B.n116 585
R362 B.n459 B.n458 585
R363 B.n460 B.n115 585
R364 B.n462 B.n461 585
R365 B.n463 B.n114 585
R366 B.n465 B.n464 585
R367 B.n466 B.n113 585
R368 B.n468 B.n467 585
R369 B.n469 B.n112 585
R370 B.n471 B.n470 585
R371 B.n472 B.n111 585
R372 B.n474 B.n473 585
R373 B.n475 B.n110 585
R374 B.n477 B.n476 585
R375 B.n478 B.n109 585
R376 B.n480 B.n479 585
R377 B.n481 B.n108 585
R378 B.n483 B.n482 585
R379 B.n484 B.n107 585
R380 B.n486 B.n485 585
R381 B.n487 B.n106 585
R382 B.n489 B.n488 585
R383 B.n490 B.n105 585
R384 B.n492 B.n491 585
R385 B.n493 B.n104 585
R386 B.n495 B.n494 585
R387 B.n496 B.n103 585
R388 B.n498 B.n497 585
R389 B.n499 B.n102 585
R390 B.n501 B.n500 585
R391 B.n502 B.n101 585
R392 B.n504 B.n503 585
R393 B.n505 B.n100 585
R394 B.n507 B.n506 585
R395 B.n508 B.n99 585
R396 B.n510 B.n509 585
R397 B.n511 B.n98 585
R398 B.n513 B.n512 585
R399 B.n514 B.n97 585
R400 B.n516 B.n515 585
R401 B.n517 B.n96 585
R402 B.n519 B.n518 585
R403 B.n520 B.n95 585
R404 B.n522 B.n521 585
R405 B.n523 B.n94 585
R406 B.n525 B.n524 585
R407 B.n526 B.n93 585
R408 B.n528 B.n527 585
R409 B.n529 B.n92 585
R410 B.n531 B.n530 585
R411 B.n532 B.n91 585
R412 B.n534 B.n533 585
R413 B.n535 B.n90 585
R414 B.n537 B.n536 585
R415 B.n538 B.n89 585
R416 B.n540 B.n539 585
R417 B.n541 B.n88 585
R418 B.n543 B.n542 585
R419 B.n544 B.n87 585
R420 B.n546 B.n545 585
R421 B.n547 B.n86 585
R422 B.n549 B.n548 585
R423 B.n735 B.n734 585
R424 B.n733 B.n20 585
R425 B.n732 B.n731 585
R426 B.n730 B.n21 585
R427 B.n729 B.n728 585
R428 B.n727 B.n22 585
R429 B.n726 B.n725 585
R430 B.n724 B.n23 585
R431 B.n723 B.n722 585
R432 B.n721 B.n24 585
R433 B.n720 B.n719 585
R434 B.n718 B.n25 585
R435 B.n717 B.n716 585
R436 B.n715 B.n26 585
R437 B.n714 B.n713 585
R438 B.n712 B.n27 585
R439 B.n711 B.n710 585
R440 B.n709 B.n28 585
R441 B.n708 B.n707 585
R442 B.n706 B.n29 585
R443 B.n705 B.n704 585
R444 B.n703 B.n30 585
R445 B.n702 B.n701 585
R446 B.n700 B.n31 585
R447 B.n699 B.n698 585
R448 B.n697 B.n32 585
R449 B.n696 B.n695 585
R450 B.n694 B.n33 585
R451 B.n693 B.n692 585
R452 B.n691 B.n34 585
R453 B.n690 B.n689 585
R454 B.n688 B.n35 585
R455 B.n687 B.n686 585
R456 B.n685 B.n36 585
R457 B.n684 B.n683 585
R458 B.n682 B.n37 585
R459 B.n681 B.n680 585
R460 B.n679 B.n38 585
R461 B.n678 B.n677 585
R462 B.n676 B.n39 585
R463 B.n675 B.n674 585
R464 B.n673 B.n40 585
R465 B.n672 B.n671 585
R466 B.n670 B.n41 585
R467 B.n669 B.n668 585
R468 B.n667 B.n42 585
R469 B.n666 B.n665 585
R470 B.n664 B.n43 585
R471 B.n663 B.n662 585
R472 B.n661 B.n44 585
R473 B.n660 B.n659 585
R474 B.n658 B.n45 585
R475 B.n657 B.n656 585
R476 B.n655 B.n46 585
R477 B.n654 B.n653 585
R478 B.n652 B.n47 585
R479 B.n651 B.n650 585
R480 B.n649 B.n648 585
R481 B.n647 B.n51 585
R482 B.n646 B.n645 585
R483 B.n644 B.n52 585
R484 B.n643 B.n642 585
R485 B.n641 B.n53 585
R486 B.n640 B.n639 585
R487 B.n638 B.n54 585
R488 B.n637 B.n636 585
R489 B.n634 B.n55 585
R490 B.n633 B.n632 585
R491 B.n631 B.n58 585
R492 B.n630 B.n629 585
R493 B.n628 B.n59 585
R494 B.n627 B.n626 585
R495 B.n625 B.n60 585
R496 B.n624 B.n623 585
R497 B.n622 B.n61 585
R498 B.n621 B.n620 585
R499 B.n619 B.n62 585
R500 B.n618 B.n617 585
R501 B.n616 B.n63 585
R502 B.n615 B.n614 585
R503 B.n613 B.n64 585
R504 B.n612 B.n611 585
R505 B.n610 B.n65 585
R506 B.n609 B.n608 585
R507 B.n607 B.n66 585
R508 B.n606 B.n605 585
R509 B.n604 B.n67 585
R510 B.n603 B.n602 585
R511 B.n601 B.n68 585
R512 B.n600 B.n599 585
R513 B.n598 B.n69 585
R514 B.n597 B.n596 585
R515 B.n595 B.n70 585
R516 B.n594 B.n593 585
R517 B.n592 B.n71 585
R518 B.n591 B.n590 585
R519 B.n589 B.n72 585
R520 B.n588 B.n587 585
R521 B.n586 B.n73 585
R522 B.n585 B.n584 585
R523 B.n583 B.n74 585
R524 B.n582 B.n581 585
R525 B.n580 B.n75 585
R526 B.n579 B.n578 585
R527 B.n577 B.n76 585
R528 B.n576 B.n575 585
R529 B.n574 B.n77 585
R530 B.n573 B.n572 585
R531 B.n571 B.n78 585
R532 B.n570 B.n569 585
R533 B.n568 B.n79 585
R534 B.n567 B.n566 585
R535 B.n565 B.n80 585
R536 B.n564 B.n563 585
R537 B.n562 B.n81 585
R538 B.n561 B.n560 585
R539 B.n559 B.n82 585
R540 B.n558 B.n557 585
R541 B.n556 B.n83 585
R542 B.n555 B.n554 585
R543 B.n553 B.n84 585
R544 B.n552 B.n551 585
R545 B.n550 B.n85 585
R546 B.n736 B.n19 585
R547 B.n738 B.n737 585
R548 B.n739 B.n18 585
R549 B.n741 B.n740 585
R550 B.n742 B.n17 585
R551 B.n744 B.n743 585
R552 B.n745 B.n16 585
R553 B.n747 B.n746 585
R554 B.n748 B.n15 585
R555 B.n750 B.n749 585
R556 B.n751 B.n14 585
R557 B.n753 B.n752 585
R558 B.n754 B.n13 585
R559 B.n756 B.n755 585
R560 B.n757 B.n12 585
R561 B.n759 B.n758 585
R562 B.n760 B.n11 585
R563 B.n762 B.n761 585
R564 B.n763 B.n10 585
R565 B.n765 B.n764 585
R566 B.n766 B.n9 585
R567 B.n768 B.n767 585
R568 B.n769 B.n8 585
R569 B.n771 B.n770 585
R570 B.n772 B.n7 585
R571 B.n774 B.n773 585
R572 B.n775 B.n6 585
R573 B.n777 B.n776 585
R574 B.n778 B.n5 585
R575 B.n780 B.n779 585
R576 B.n781 B.n4 585
R577 B.n783 B.n782 585
R578 B.n784 B.n3 585
R579 B.n786 B.n785 585
R580 B.n787 B.n0 585
R581 B.n2 B.n1 585
R582 B.n205 B.n204 585
R583 B.n207 B.n206 585
R584 B.n208 B.n203 585
R585 B.n210 B.n209 585
R586 B.n211 B.n202 585
R587 B.n213 B.n212 585
R588 B.n214 B.n201 585
R589 B.n216 B.n215 585
R590 B.n217 B.n200 585
R591 B.n219 B.n218 585
R592 B.n220 B.n199 585
R593 B.n222 B.n221 585
R594 B.n223 B.n198 585
R595 B.n225 B.n224 585
R596 B.n226 B.n197 585
R597 B.n228 B.n227 585
R598 B.n229 B.n196 585
R599 B.n231 B.n230 585
R600 B.n232 B.n195 585
R601 B.n234 B.n233 585
R602 B.n235 B.n194 585
R603 B.n237 B.n236 585
R604 B.n238 B.n193 585
R605 B.n240 B.n239 585
R606 B.n241 B.n192 585
R607 B.n243 B.n242 585
R608 B.n244 B.n191 585
R609 B.n246 B.n245 585
R610 B.n247 B.n190 585
R611 B.n249 B.n248 585
R612 B.n250 B.n189 585
R613 B.n252 B.n251 585
R614 B.n253 B.n188 585
R615 B.n255 B.n254 585
R616 B.n254 B.n187 554.963
R617 B.n440 B.n121 554.963
R618 B.n548 B.n85 554.963
R619 B.n734 B.n19 554.963
R620 B.n158 B.t9 541.279
R621 B.n150 B.t0 541.279
R622 B.n56 B.t3 541.279
R623 B.n48 B.t6 541.279
R624 B.n789 B.n788 256.663
R625 B.n788 B.n787 235.042
R626 B.n788 B.n2 235.042
R627 B.n258 B.n187 163.367
R628 B.n259 B.n258 163.367
R629 B.n260 B.n259 163.367
R630 B.n260 B.n185 163.367
R631 B.n264 B.n185 163.367
R632 B.n265 B.n264 163.367
R633 B.n266 B.n265 163.367
R634 B.n266 B.n183 163.367
R635 B.n270 B.n183 163.367
R636 B.n271 B.n270 163.367
R637 B.n272 B.n271 163.367
R638 B.n272 B.n181 163.367
R639 B.n276 B.n181 163.367
R640 B.n277 B.n276 163.367
R641 B.n278 B.n277 163.367
R642 B.n278 B.n179 163.367
R643 B.n282 B.n179 163.367
R644 B.n283 B.n282 163.367
R645 B.n284 B.n283 163.367
R646 B.n284 B.n177 163.367
R647 B.n288 B.n177 163.367
R648 B.n289 B.n288 163.367
R649 B.n290 B.n289 163.367
R650 B.n290 B.n175 163.367
R651 B.n294 B.n175 163.367
R652 B.n295 B.n294 163.367
R653 B.n296 B.n295 163.367
R654 B.n296 B.n173 163.367
R655 B.n300 B.n173 163.367
R656 B.n301 B.n300 163.367
R657 B.n302 B.n301 163.367
R658 B.n302 B.n171 163.367
R659 B.n306 B.n171 163.367
R660 B.n307 B.n306 163.367
R661 B.n308 B.n307 163.367
R662 B.n308 B.n169 163.367
R663 B.n312 B.n169 163.367
R664 B.n313 B.n312 163.367
R665 B.n314 B.n313 163.367
R666 B.n314 B.n167 163.367
R667 B.n318 B.n167 163.367
R668 B.n319 B.n318 163.367
R669 B.n320 B.n319 163.367
R670 B.n320 B.n165 163.367
R671 B.n324 B.n165 163.367
R672 B.n325 B.n324 163.367
R673 B.n326 B.n325 163.367
R674 B.n326 B.n163 163.367
R675 B.n330 B.n163 163.367
R676 B.n331 B.n330 163.367
R677 B.n332 B.n331 163.367
R678 B.n332 B.n161 163.367
R679 B.n336 B.n161 163.367
R680 B.n337 B.n336 163.367
R681 B.n338 B.n337 163.367
R682 B.n338 B.n157 163.367
R683 B.n343 B.n157 163.367
R684 B.n344 B.n343 163.367
R685 B.n345 B.n344 163.367
R686 B.n345 B.n155 163.367
R687 B.n349 B.n155 163.367
R688 B.n350 B.n349 163.367
R689 B.n351 B.n350 163.367
R690 B.n351 B.n153 163.367
R691 B.n355 B.n153 163.367
R692 B.n356 B.n355 163.367
R693 B.n356 B.n149 163.367
R694 B.n360 B.n149 163.367
R695 B.n361 B.n360 163.367
R696 B.n362 B.n361 163.367
R697 B.n362 B.n147 163.367
R698 B.n366 B.n147 163.367
R699 B.n367 B.n366 163.367
R700 B.n368 B.n367 163.367
R701 B.n368 B.n145 163.367
R702 B.n372 B.n145 163.367
R703 B.n373 B.n372 163.367
R704 B.n374 B.n373 163.367
R705 B.n374 B.n143 163.367
R706 B.n378 B.n143 163.367
R707 B.n379 B.n378 163.367
R708 B.n380 B.n379 163.367
R709 B.n380 B.n141 163.367
R710 B.n384 B.n141 163.367
R711 B.n385 B.n384 163.367
R712 B.n386 B.n385 163.367
R713 B.n386 B.n139 163.367
R714 B.n390 B.n139 163.367
R715 B.n391 B.n390 163.367
R716 B.n392 B.n391 163.367
R717 B.n392 B.n137 163.367
R718 B.n396 B.n137 163.367
R719 B.n397 B.n396 163.367
R720 B.n398 B.n397 163.367
R721 B.n398 B.n135 163.367
R722 B.n402 B.n135 163.367
R723 B.n403 B.n402 163.367
R724 B.n404 B.n403 163.367
R725 B.n404 B.n133 163.367
R726 B.n408 B.n133 163.367
R727 B.n409 B.n408 163.367
R728 B.n410 B.n409 163.367
R729 B.n410 B.n131 163.367
R730 B.n414 B.n131 163.367
R731 B.n415 B.n414 163.367
R732 B.n416 B.n415 163.367
R733 B.n416 B.n129 163.367
R734 B.n420 B.n129 163.367
R735 B.n421 B.n420 163.367
R736 B.n422 B.n421 163.367
R737 B.n422 B.n127 163.367
R738 B.n426 B.n127 163.367
R739 B.n427 B.n426 163.367
R740 B.n428 B.n427 163.367
R741 B.n428 B.n125 163.367
R742 B.n432 B.n125 163.367
R743 B.n433 B.n432 163.367
R744 B.n434 B.n433 163.367
R745 B.n434 B.n123 163.367
R746 B.n438 B.n123 163.367
R747 B.n439 B.n438 163.367
R748 B.n440 B.n439 163.367
R749 B.n548 B.n547 163.367
R750 B.n547 B.n546 163.367
R751 B.n546 B.n87 163.367
R752 B.n542 B.n87 163.367
R753 B.n542 B.n541 163.367
R754 B.n541 B.n540 163.367
R755 B.n540 B.n89 163.367
R756 B.n536 B.n89 163.367
R757 B.n536 B.n535 163.367
R758 B.n535 B.n534 163.367
R759 B.n534 B.n91 163.367
R760 B.n530 B.n91 163.367
R761 B.n530 B.n529 163.367
R762 B.n529 B.n528 163.367
R763 B.n528 B.n93 163.367
R764 B.n524 B.n93 163.367
R765 B.n524 B.n523 163.367
R766 B.n523 B.n522 163.367
R767 B.n522 B.n95 163.367
R768 B.n518 B.n95 163.367
R769 B.n518 B.n517 163.367
R770 B.n517 B.n516 163.367
R771 B.n516 B.n97 163.367
R772 B.n512 B.n97 163.367
R773 B.n512 B.n511 163.367
R774 B.n511 B.n510 163.367
R775 B.n510 B.n99 163.367
R776 B.n506 B.n99 163.367
R777 B.n506 B.n505 163.367
R778 B.n505 B.n504 163.367
R779 B.n504 B.n101 163.367
R780 B.n500 B.n101 163.367
R781 B.n500 B.n499 163.367
R782 B.n499 B.n498 163.367
R783 B.n498 B.n103 163.367
R784 B.n494 B.n103 163.367
R785 B.n494 B.n493 163.367
R786 B.n493 B.n492 163.367
R787 B.n492 B.n105 163.367
R788 B.n488 B.n105 163.367
R789 B.n488 B.n487 163.367
R790 B.n487 B.n486 163.367
R791 B.n486 B.n107 163.367
R792 B.n482 B.n107 163.367
R793 B.n482 B.n481 163.367
R794 B.n481 B.n480 163.367
R795 B.n480 B.n109 163.367
R796 B.n476 B.n109 163.367
R797 B.n476 B.n475 163.367
R798 B.n475 B.n474 163.367
R799 B.n474 B.n111 163.367
R800 B.n470 B.n111 163.367
R801 B.n470 B.n469 163.367
R802 B.n469 B.n468 163.367
R803 B.n468 B.n113 163.367
R804 B.n464 B.n113 163.367
R805 B.n464 B.n463 163.367
R806 B.n463 B.n462 163.367
R807 B.n462 B.n115 163.367
R808 B.n458 B.n115 163.367
R809 B.n458 B.n457 163.367
R810 B.n457 B.n456 163.367
R811 B.n456 B.n117 163.367
R812 B.n452 B.n117 163.367
R813 B.n452 B.n451 163.367
R814 B.n451 B.n450 163.367
R815 B.n450 B.n119 163.367
R816 B.n446 B.n119 163.367
R817 B.n446 B.n445 163.367
R818 B.n445 B.n444 163.367
R819 B.n444 B.n121 163.367
R820 B.n734 B.n733 163.367
R821 B.n733 B.n732 163.367
R822 B.n732 B.n21 163.367
R823 B.n728 B.n21 163.367
R824 B.n728 B.n727 163.367
R825 B.n727 B.n726 163.367
R826 B.n726 B.n23 163.367
R827 B.n722 B.n23 163.367
R828 B.n722 B.n721 163.367
R829 B.n721 B.n720 163.367
R830 B.n720 B.n25 163.367
R831 B.n716 B.n25 163.367
R832 B.n716 B.n715 163.367
R833 B.n715 B.n714 163.367
R834 B.n714 B.n27 163.367
R835 B.n710 B.n27 163.367
R836 B.n710 B.n709 163.367
R837 B.n709 B.n708 163.367
R838 B.n708 B.n29 163.367
R839 B.n704 B.n29 163.367
R840 B.n704 B.n703 163.367
R841 B.n703 B.n702 163.367
R842 B.n702 B.n31 163.367
R843 B.n698 B.n31 163.367
R844 B.n698 B.n697 163.367
R845 B.n697 B.n696 163.367
R846 B.n696 B.n33 163.367
R847 B.n692 B.n33 163.367
R848 B.n692 B.n691 163.367
R849 B.n691 B.n690 163.367
R850 B.n690 B.n35 163.367
R851 B.n686 B.n35 163.367
R852 B.n686 B.n685 163.367
R853 B.n685 B.n684 163.367
R854 B.n684 B.n37 163.367
R855 B.n680 B.n37 163.367
R856 B.n680 B.n679 163.367
R857 B.n679 B.n678 163.367
R858 B.n678 B.n39 163.367
R859 B.n674 B.n39 163.367
R860 B.n674 B.n673 163.367
R861 B.n673 B.n672 163.367
R862 B.n672 B.n41 163.367
R863 B.n668 B.n41 163.367
R864 B.n668 B.n667 163.367
R865 B.n667 B.n666 163.367
R866 B.n666 B.n43 163.367
R867 B.n662 B.n43 163.367
R868 B.n662 B.n661 163.367
R869 B.n661 B.n660 163.367
R870 B.n660 B.n45 163.367
R871 B.n656 B.n45 163.367
R872 B.n656 B.n655 163.367
R873 B.n655 B.n654 163.367
R874 B.n654 B.n47 163.367
R875 B.n650 B.n47 163.367
R876 B.n650 B.n649 163.367
R877 B.n649 B.n51 163.367
R878 B.n645 B.n51 163.367
R879 B.n645 B.n644 163.367
R880 B.n644 B.n643 163.367
R881 B.n643 B.n53 163.367
R882 B.n639 B.n53 163.367
R883 B.n639 B.n638 163.367
R884 B.n638 B.n637 163.367
R885 B.n637 B.n55 163.367
R886 B.n632 B.n55 163.367
R887 B.n632 B.n631 163.367
R888 B.n631 B.n630 163.367
R889 B.n630 B.n59 163.367
R890 B.n626 B.n59 163.367
R891 B.n626 B.n625 163.367
R892 B.n625 B.n624 163.367
R893 B.n624 B.n61 163.367
R894 B.n620 B.n61 163.367
R895 B.n620 B.n619 163.367
R896 B.n619 B.n618 163.367
R897 B.n618 B.n63 163.367
R898 B.n614 B.n63 163.367
R899 B.n614 B.n613 163.367
R900 B.n613 B.n612 163.367
R901 B.n612 B.n65 163.367
R902 B.n608 B.n65 163.367
R903 B.n608 B.n607 163.367
R904 B.n607 B.n606 163.367
R905 B.n606 B.n67 163.367
R906 B.n602 B.n67 163.367
R907 B.n602 B.n601 163.367
R908 B.n601 B.n600 163.367
R909 B.n600 B.n69 163.367
R910 B.n596 B.n69 163.367
R911 B.n596 B.n595 163.367
R912 B.n595 B.n594 163.367
R913 B.n594 B.n71 163.367
R914 B.n590 B.n71 163.367
R915 B.n590 B.n589 163.367
R916 B.n589 B.n588 163.367
R917 B.n588 B.n73 163.367
R918 B.n584 B.n73 163.367
R919 B.n584 B.n583 163.367
R920 B.n583 B.n582 163.367
R921 B.n582 B.n75 163.367
R922 B.n578 B.n75 163.367
R923 B.n578 B.n577 163.367
R924 B.n577 B.n576 163.367
R925 B.n576 B.n77 163.367
R926 B.n572 B.n77 163.367
R927 B.n572 B.n571 163.367
R928 B.n571 B.n570 163.367
R929 B.n570 B.n79 163.367
R930 B.n566 B.n79 163.367
R931 B.n566 B.n565 163.367
R932 B.n565 B.n564 163.367
R933 B.n564 B.n81 163.367
R934 B.n560 B.n81 163.367
R935 B.n560 B.n559 163.367
R936 B.n559 B.n558 163.367
R937 B.n558 B.n83 163.367
R938 B.n554 B.n83 163.367
R939 B.n554 B.n553 163.367
R940 B.n553 B.n552 163.367
R941 B.n552 B.n85 163.367
R942 B.n738 B.n19 163.367
R943 B.n739 B.n738 163.367
R944 B.n740 B.n739 163.367
R945 B.n740 B.n17 163.367
R946 B.n744 B.n17 163.367
R947 B.n745 B.n744 163.367
R948 B.n746 B.n745 163.367
R949 B.n746 B.n15 163.367
R950 B.n750 B.n15 163.367
R951 B.n751 B.n750 163.367
R952 B.n752 B.n751 163.367
R953 B.n752 B.n13 163.367
R954 B.n756 B.n13 163.367
R955 B.n757 B.n756 163.367
R956 B.n758 B.n757 163.367
R957 B.n758 B.n11 163.367
R958 B.n762 B.n11 163.367
R959 B.n763 B.n762 163.367
R960 B.n764 B.n763 163.367
R961 B.n764 B.n9 163.367
R962 B.n768 B.n9 163.367
R963 B.n769 B.n768 163.367
R964 B.n770 B.n769 163.367
R965 B.n770 B.n7 163.367
R966 B.n774 B.n7 163.367
R967 B.n775 B.n774 163.367
R968 B.n776 B.n775 163.367
R969 B.n776 B.n5 163.367
R970 B.n780 B.n5 163.367
R971 B.n781 B.n780 163.367
R972 B.n782 B.n781 163.367
R973 B.n782 B.n3 163.367
R974 B.n786 B.n3 163.367
R975 B.n787 B.n786 163.367
R976 B.n205 B.n2 163.367
R977 B.n206 B.n205 163.367
R978 B.n206 B.n203 163.367
R979 B.n210 B.n203 163.367
R980 B.n211 B.n210 163.367
R981 B.n212 B.n211 163.367
R982 B.n212 B.n201 163.367
R983 B.n216 B.n201 163.367
R984 B.n217 B.n216 163.367
R985 B.n218 B.n217 163.367
R986 B.n218 B.n199 163.367
R987 B.n222 B.n199 163.367
R988 B.n223 B.n222 163.367
R989 B.n224 B.n223 163.367
R990 B.n224 B.n197 163.367
R991 B.n228 B.n197 163.367
R992 B.n229 B.n228 163.367
R993 B.n230 B.n229 163.367
R994 B.n230 B.n195 163.367
R995 B.n234 B.n195 163.367
R996 B.n235 B.n234 163.367
R997 B.n236 B.n235 163.367
R998 B.n236 B.n193 163.367
R999 B.n240 B.n193 163.367
R1000 B.n241 B.n240 163.367
R1001 B.n242 B.n241 163.367
R1002 B.n242 B.n191 163.367
R1003 B.n246 B.n191 163.367
R1004 B.n247 B.n246 163.367
R1005 B.n248 B.n247 163.367
R1006 B.n248 B.n189 163.367
R1007 B.n252 B.n189 163.367
R1008 B.n253 B.n252 163.367
R1009 B.n254 B.n253 163.367
R1010 B.n150 B.t1 140.421
R1011 B.n56 B.t5 140.421
R1012 B.n158 B.t10 140.399
R1013 B.n48 B.t8 140.399
R1014 B.n151 B.t2 110.165
R1015 B.n57 B.t4 110.165
R1016 B.n159 B.t11 110.144
R1017 B.n49 B.t7 110.144
R1018 B.n341 B.n159 59.5399
R1019 B.n152 B.n151 59.5399
R1020 B.n635 B.n57 59.5399
R1021 B.n50 B.n49 59.5399
R1022 B.n736 B.n735 36.059
R1023 B.n550 B.n549 36.059
R1024 B.n256 B.n255 36.059
R1025 B.n442 B.n441 36.059
R1026 B.n159 B.n158 30.255
R1027 B.n151 B.n150 30.255
R1028 B.n57 B.n56 30.255
R1029 B.n49 B.n48 30.255
R1030 B B.n789 18.0485
R1031 B.n737 B.n736 10.6151
R1032 B.n737 B.n18 10.6151
R1033 B.n741 B.n18 10.6151
R1034 B.n742 B.n741 10.6151
R1035 B.n743 B.n742 10.6151
R1036 B.n743 B.n16 10.6151
R1037 B.n747 B.n16 10.6151
R1038 B.n748 B.n747 10.6151
R1039 B.n749 B.n748 10.6151
R1040 B.n749 B.n14 10.6151
R1041 B.n753 B.n14 10.6151
R1042 B.n754 B.n753 10.6151
R1043 B.n755 B.n754 10.6151
R1044 B.n755 B.n12 10.6151
R1045 B.n759 B.n12 10.6151
R1046 B.n760 B.n759 10.6151
R1047 B.n761 B.n760 10.6151
R1048 B.n761 B.n10 10.6151
R1049 B.n765 B.n10 10.6151
R1050 B.n766 B.n765 10.6151
R1051 B.n767 B.n766 10.6151
R1052 B.n767 B.n8 10.6151
R1053 B.n771 B.n8 10.6151
R1054 B.n772 B.n771 10.6151
R1055 B.n773 B.n772 10.6151
R1056 B.n773 B.n6 10.6151
R1057 B.n777 B.n6 10.6151
R1058 B.n778 B.n777 10.6151
R1059 B.n779 B.n778 10.6151
R1060 B.n779 B.n4 10.6151
R1061 B.n783 B.n4 10.6151
R1062 B.n784 B.n783 10.6151
R1063 B.n785 B.n784 10.6151
R1064 B.n785 B.n0 10.6151
R1065 B.n735 B.n20 10.6151
R1066 B.n731 B.n20 10.6151
R1067 B.n731 B.n730 10.6151
R1068 B.n730 B.n729 10.6151
R1069 B.n729 B.n22 10.6151
R1070 B.n725 B.n22 10.6151
R1071 B.n725 B.n724 10.6151
R1072 B.n724 B.n723 10.6151
R1073 B.n723 B.n24 10.6151
R1074 B.n719 B.n24 10.6151
R1075 B.n719 B.n718 10.6151
R1076 B.n718 B.n717 10.6151
R1077 B.n717 B.n26 10.6151
R1078 B.n713 B.n26 10.6151
R1079 B.n713 B.n712 10.6151
R1080 B.n712 B.n711 10.6151
R1081 B.n711 B.n28 10.6151
R1082 B.n707 B.n28 10.6151
R1083 B.n707 B.n706 10.6151
R1084 B.n706 B.n705 10.6151
R1085 B.n705 B.n30 10.6151
R1086 B.n701 B.n30 10.6151
R1087 B.n701 B.n700 10.6151
R1088 B.n700 B.n699 10.6151
R1089 B.n699 B.n32 10.6151
R1090 B.n695 B.n32 10.6151
R1091 B.n695 B.n694 10.6151
R1092 B.n694 B.n693 10.6151
R1093 B.n693 B.n34 10.6151
R1094 B.n689 B.n34 10.6151
R1095 B.n689 B.n688 10.6151
R1096 B.n688 B.n687 10.6151
R1097 B.n687 B.n36 10.6151
R1098 B.n683 B.n36 10.6151
R1099 B.n683 B.n682 10.6151
R1100 B.n682 B.n681 10.6151
R1101 B.n681 B.n38 10.6151
R1102 B.n677 B.n38 10.6151
R1103 B.n677 B.n676 10.6151
R1104 B.n676 B.n675 10.6151
R1105 B.n675 B.n40 10.6151
R1106 B.n671 B.n40 10.6151
R1107 B.n671 B.n670 10.6151
R1108 B.n670 B.n669 10.6151
R1109 B.n669 B.n42 10.6151
R1110 B.n665 B.n42 10.6151
R1111 B.n665 B.n664 10.6151
R1112 B.n664 B.n663 10.6151
R1113 B.n663 B.n44 10.6151
R1114 B.n659 B.n44 10.6151
R1115 B.n659 B.n658 10.6151
R1116 B.n658 B.n657 10.6151
R1117 B.n657 B.n46 10.6151
R1118 B.n653 B.n46 10.6151
R1119 B.n653 B.n652 10.6151
R1120 B.n652 B.n651 10.6151
R1121 B.n648 B.n647 10.6151
R1122 B.n647 B.n646 10.6151
R1123 B.n646 B.n52 10.6151
R1124 B.n642 B.n52 10.6151
R1125 B.n642 B.n641 10.6151
R1126 B.n641 B.n640 10.6151
R1127 B.n640 B.n54 10.6151
R1128 B.n636 B.n54 10.6151
R1129 B.n634 B.n633 10.6151
R1130 B.n633 B.n58 10.6151
R1131 B.n629 B.n58 10.6151
R1132 B.n629 B.n628 10.6151
R1133 B.n628 B.n627 10.6151
R1134 B.n627 B.n60 10.6151
R1135 B.n623 B.n60 10.6151
R1136 B.n623 B.n622 10.6151
R1137 B.n622 B.n621 10.6151
R1138 B.n621 B.n62 10.6151
R1139 B.n617 B.n62 10.6151
R1140 B.n617 B.n616 10.6151
R1141 B.n616 B.n615 10.6151
R1142 B.n615 B.n64 10.6151
R1143 B.n611 B.n64 10.6151
R1144 B.n611 B.n610 10.6151
R1145 B.n610 B.n609 10.6151
R1146 B.n609 B.n66 10.6151
R1147 B.n605 B.n66 10.6151
R1148 B.n605 B.n604 10.6151
R1149 B.n604 B.n603 10.6151
R1150 B.n603 B.n68 10.6151
R1151 B.n599 B.n68 10.6151
R1152 B.n599 B.n598 10.6151
R1153 B.n598 B.n597 10.6151
R1154 B.n597 B.n70 10.6151
R1155 B.n593 B.n70 10.6151
R1156 B.n593 B.n592 10.6151
R1157 B.n592 B.n591 10.6151
R1158 B.n591 B.n72 10.6151
R1159 B.n587 B.n72 10.6151
R1160 B.n587 B.n586 10.6151
R1161 B.n586 B.n585 10.6151
R1162 B.n585 B.n74 10.6151
R1163 B.n581 B.n74 10.6151
R1164 B.n581 B.n580 10.6151
R1165 B.n580 B.n579 10.6151
R1166 B.n579 B.n76 10.6151
R1167 B.n575 B.n76 10.6151
R1168 B.n575 B.n574 10.6151
R1169 B.n574 B.n573 10.6151
R1170 B.n573 B.n78 10.6151
R1171 B.n569 B.n78 10.6151
R1172 B.n569 B.n568 10.6151
R1173 B.n568 B.n567 10.6151
R1174 B.n567 B.n80 10.6151
R1175 B.n563 B.n80 10.6151
R1176 B.n563 B.n562 10.6151
R1177 B.n562 B.n561 10.6151
R1178 B.n561 B.n82 10.6151
R1179 B.n557 B.n82 10.6151
R1180 B.n557 B.n556 10.6151
R1181 B.n556 B.n555 10.6151
R1182 B.n555 B.n84 10.6151
R1183 B.n551 B.n84 10.6151
R1184 B.n551 B.n550 10.6151
R1185 B.n549 B.n86 10.6151
R1186 B.n545 B.n86 10.6151
R1187 B.n545 B.n544 10.6151
R1188 B.n544 B.n543 10.6151
R1189 B.n543 B.n88 10.6151
R1190 B.n539 B.n88 10.6151
R1191 B.n539 B.n538 10.6151
R1192 B.n538 B.n537 10.6151
R1193 B.n537 B.n90 10.6151
R1194 B.n533 B.n90 10.6151
R1195 B.n533 B.n532 10.6151
R1196 B.n532 B.n531 10.6151
R1197 B.n531 B.n92 10.6151
R1198 B.n527 B.n92 10.6151
R1199 B.n527 B.n526 10.6151
R1200 B.n526 B.n525 10.6151
R1201 B.n525 B.n94 10.6151
R1202 B.n521 B.n94 10.6151
R1203 B.n521 B.n520 10.6151
R1204 B.n520 B.n519 10.6151
R1205 B.n519 B.n96 10.6151
R1206 B.n515 B.n96 10.6151
R1207 B.n515 B.n514 10.6151
R1208 B.n514 B.n513 10.6151
R1209 B.n513 B.n98 10.6151
R1210 B.n509 B.n98 10.6151
R1211 B.n509 B.n508 10.6151
R1212 B.n508 B.n507 10.6151
R1213 B.n507 B.n100 10.6151
R1214 B.n503 B.n100 10.6151
R1215 B.n503 B.n502 10.6151
R1216 B.n502 B.n501 10.6151
R1217 B.n501 B.n102 10.6151
R1218 B.n497 B.n102 10.6151
R1219 B.n497 B.n496 10.6151
R1220 B.n496 B.n495 10.6151
R1221 B.n495 B.n104 10.6151
R1222 B.n491 B.n104 10.6151
R1223 B.n491 B.n490 10.6151
R1224 B.n490 B.n489 10.6151
R1225 B.n489 B.n106 10.6151
R1226 B.n485 B.n106 10.6151
R1227 B.n485 B.n484 10.6151
R1228 B.n484 B.n483 10.6151
R1229 B.n483 B.n108 10.6151
R1230 B.n479 B.n108 10.6151
R1231 B.n479 B.n478 10.6151
R1232 B.n478 B.n477 10.6151
R1233 B.n477 B.n110 10.6151
R1234 B.n473 B.n110 10.6151
R1235 B.n473 B.n472 10.6151
R1236 B.n472 B.n471 10.6151
R1237 B.n471 B.n112 10.6151
R1238 B.n467 B.n112 10.6151
R1239 B.n467 B.n466 10.6151
R1240 B.n466 B.n465 10.6151
R1241 B.n465 B.n114 10.6151
R1242 B.n461 B.n114 10.6151
R1243 B.n461 B.n460 10.6151
R1244 B.n460 B.n459 10.6151
R1245 B.n459 B.n116 10.6151
R1246 B.n455 B.n116 10.6151
R1247 B.n455 B.n454 10.6151
R1248 B.n454 B.n453 10.6151
R1249 B.n453 B.n118 10.6151
R1250 B.n449 B.n118 10.6151
R1251 B.n449 B.n448 10.6151
R1252 B.n448 B.n447 10.6151
R1253 B.n447 B.n120 10.6151
R1254 B.n443 B.n120 10.6151
R1255 B.n443 B.n442 10.6151
R1256 B.n204 B.n1 10.6151
R1257 B.n207 B.n204 10.6151
R1258 B.n208 B.n207 10.6151
R1259 B.n209 B.n208 10.6151
R1260 B.n209 B.n202 10.6151
R1261 B.n213 B.n202 10.6151
R1262 B.n214 B.n213 10.6151
R1263 B.n215 B.n214 10.6151
R1264 B.n215 B.n200 10.6151
R1265 B.n219 B.n200 10.6151
R1266 B.n220 B.n219 10.6151
R1267 B.n221 B.n220 10.6151
R1268 B.n221 B.n198 10.6151
R1269 B.n225 B.n198 10.6151
R1270 B.n226 B.n225 10.6151
R1271 B.n227 B.n226 10.6151
R1272 B.n227 B.n196 10.6151
R1273 B.n231 B.n196 10.6151
R1274 B.n232 B.n231 10.6151
R1275 B.n233 B.n232 10.6151
R1276 B.n233 B.n194 10.6151
R1277 B.n237 B.n194 10.6151
R1278 B.n238 B.n237 10.6151
R1279 B.n239 B.n238 10.6151
R1280 B.n239 B.n192 10.6151
R1281 B.n243 B.n192 10.6151
R1282 B.n244 B.n243 10.6151
R1283 B.n245 B.n244 10.6151
R1284 B.n245 B.n190 10.6151
R1285 B.n249 B.n190 10.6151
R1286 B.n250 B.n249 10.6151
R1287 B.n251 B.n250 10.6151
R1288 B.n251 B.n188 10.6151
R1289 B.n255 B.n188 10.6151
R1290 B.n257 B.n256 10.6151
R1291 B.n257 B.n186 10.6151
R1292 B.n261 B.n186 10.6151
R1293 B.n262 B.n261 10.6151
R1294 B.n263 B.n262 10.6151
R1295 B.n263 B.n184 10.6151
R1296 B.n267 B.n184 10.6151
R1297 B.n268 B.n267 10.6151
R1298 B.n269 B.n268 10.6151
R1299 B.n269 B.n182 10.6151
R1300 B.n273 B.n182 10.6151
R1301 B.n274 B.n273 10.6151
R1302 B.n275 B.n274 10.6151
R1303 B.n275 B.n180 10.6151
R1304 B.n279 B.n180 10.6151
R1305 B.n280 B.n279 10.6151
R1306 B.n281 B.n280 10.6151
R1307 B.n281 B.n178 10.6151
R1308 B.n285 B.n178 10.6151
R1309 B.n286 B.n285 10.6151
R1310 B.n287 B.n286 10.6151
R1311 B.n287 B.n176 10.6151
R1312 B.n291 B.n176 10.6151
R1313 B.n292 B.n291 10.6151
R1314 B.n293 B.n292 10.6151
R1315 B.n293 B.n174 10.6151
R1316 B.n297 B.n174 10.6151
R1317 B.n298 B.n297 10.6151
R1318 B.n299 B.n298 10.6151
R1319 B.n299 B.n172 10.6151
R1320 B.n303 B.n172 10.6151
R1321 B.n304 B.n303 10.6151
R1322 B.n305 B.n304 10.6151
R1323 B.n305 B.n170 10.6151
R1324 B.n309 B.n170 10.6151
R1325 B.n310 B.n309 10.6151
R1326 B.n311 B.n310 10.6151
R1327 B.n311 B.n168 10.6151
R1328 B.n315 B.n168 10.6151
R1329 B.n316 B.n315 10.6151
R1330 B.n317 B.n316 10.6151
R1331 B.n317 B.n166 10.6151
R1332 B.n321 B.n166 10.6151
R1333 B.n322 B.n321 10.6151
R1334 B.n323 B.n322 10.6151
R1335 B.n323 B.n164 10.6151
R1336 B.n327 B.n164 10.6151
R1337 B.n328 B.n327 10.6151
R1338 B.n329 B.n328 10.6151
R1339 B.n329 B.n162 10.6151
R1340 B.n333 B.n162 10.6151
R1341 B.n334 B.n333 10.6151
R1342 B.n335 B.n334 10.6151
R1343 B.n335 B.n160 10.6151
R1344 B.n339 B.n160 10.6151
R1345 B.n340 B.n339 10.6151
R1346 B.n342 B.n156 10.6151
R1347 B.n346 B.n156 10.6151
R1348 B.n347 B.n346 10.6151
R1349 B.n348 B.n347 10.6151
R1350 B.n348 B.n154 10.6151
R1351 B.n352 B.n154 10.6151
R1352 B.n353 B.n352 10.6151
R1353 B.n354 B.n353 10.6151
R1354 B.n358 B.n357 10.6151
R1355 B.n359 B.n358 10.6151
R1356 B.n359 B.n148 10.6151
R1357 B.n363 B.n148 10.6151
R1358 B.n364 B.n363 10.6151
R1359 B.n365 B.n364 10.6151
R1360 B.n365 B.n146 10.6151
R1361 B.n369 B.n146 10.6151
R1362 B.n370 B.n369 10.6151
R1363 B.n371 B.n370 10.6151
R1364 B.n371 B.n144 10.6151
R1365 B.n375 B.n144 10.6151
R1366 B.n376 B.n375 10.6151
R1367 B.n377 B.n376 10.6151
R1368 B.n377 B.n142 10.6151
R1369 B.n381 B.n142 10.6151
R1370 B.n382 B.n381 10.6151
R1371 B.n383 B.n382 10.6151
R1372 B.n383 B.n140 10.6151
R1373 B.n387 B.n140 10.6151
R1374 B.n388 B.n387 10.6151
R1375 B.n389 B.n388 10.6151
R1376 B.n389 B.n138 10.6151
R1377 B.n393 B.n138 10.6151
R1378 B.n394 B.n393 10.6151
R1379 B.n395 B.n394 10.6151
R1380 B.n395 B.n136 10.6151
R1381 B.n399 B.n136 10.6151
R1382 B.n400 B.n399 10.6151
R1383 B.n401 B.n400 10.6151
R1384 B.n401 B.n134 10.6151
R1385 B.n405 B.n134 10.6151
R1386 B.n406 B.n405 10.6151
R1387 B.n407 B.n406 10.6151
R1388 B.n407 B.n132 10.6151
R1389 B.n411 B.n132 10.6151
R1390 B.n412 B.n411 10.6151
R1391 B.n413 B.n412 10.6151
R1392 B.n413 B.n130 10.6151
R1393 B.n417 B.n130 10.6151
R1394 B.n418 B.n417 10.6151
R1395 B.n419 B.n418 10.6151
R1396 B.n419 B.n128 10.6151
R1397 B.n423 B.n128 10.6151
R1398 B.n424 B.n423 10.6151
R1399 B.n425 B.n424 10.6151
R1400 B.n425 B.n126 10.6151
R1401 B.n429 B.n126 10.6151
R1402 B.n430 B.n429 10.6151
R1403 B.n431 B.n430 10.6151
R1404 B.n431 B.n124 10.6151
R1405 B.n435 B.n124 10.6151
R1406 B.n436 B.n435 10.6151
R1407 B.n437 B.n436 10.6151
R1408 B.n437 B.n122 10.6151
R1409 B.n441 B.n122 10.6151
R1410 B.n789 B.n0 8.11757
R1411 B.n789 B.n1 8.11757
R1412 B.n648 B.n50 6.5566
R1413 B.n636 B.n635 6.5566
R1414 B.n342 B.n341 6.5566
R1415 B.n354 B.n152 6.5566
R1416 B.n651 B.n50 4.05904
R1417 B.n635 B.n634 4.05904
R1418 B.n341 B.n340 4.05904
R1419 B.n357 B.n152 4.05904
C0 B VDD2 2.38543f
C1 VTAIL VN 12.050401f
C2 VN VP 7.33584f
C3 w_n2842_n4408# VDD2 2.7054f
C4 w_n2842_n4408# B 9.70067f
C5 VDD1 VTAIL 15.1167f
C6 VDD1 VP 12.4392f
C7 VDD1 VN 0.150308f
C8 VTAIL VDD2 15.154f
C9 B VTAIL 4.07836f
C10 VP VDD2 0.409718f
C11 B VP 1.60578f
C12 VN VDD2 12.1855f
C13 w_n2842_n4408# VTAIL 3.81865f
C14 B VN 0.998244f
C15 w_n2842_n4408# VP 6.11903f
C16 w_n2842_n4408# VN 5.75324f
C17 VDD1 VDD2 1.29864f
C18 B VDD1 2.32083f
C19 w_n2842_n4408# VDD1 2.63304f
C20 VTAIL VP 12.0651f
C21 VDD2 VSUBS 1.810184f
C22 VDD1 VSUBS 1.537686f
C23 VTAIL VSUBS 1.120711f
C24 VN VSUBS 5.90959f
C25 VP VSUBS 2.698792f
C26 B VSUBS 4.107967f
C27 w_n2842_n4408# VSUBS 0.153297p
C28 B.n0 VSUBS 0.007549f
C29 B.n1 VSUBS 0.007549f
C30 B.n2 VSUBS 0.011165f
C31 B.n3 VSUBS 0.008556f
C32 B.n4 VSUBS 0.008556f
C33 B.n5 VSUBS 0.008556f
C34 B.n6 VSUBS 0.008556f
C35 B.n7 VSUBS 0.008556f
C36 B.n8 VSUBS 0.008556f
C37 B.n9 VSUBS 0.008556f
C38 B.n10 VSUBS 0.008556f
C39 B.n11 VSUBS 0.008556f
C40 B.n12 VSUBS 0.008556f
C41 B.n13 VSUBS 0.008556f
C42 B.n14 VSUBS 0.008556f
C43 B.n15 VSUBS 0.008556f
C44 B.n16 VSUBS 0.008556f
C45 B.n17 VSUBS 0.008556f
C46 B.n18 VSUBS 0.008556f
C47 B.n19 VSUBS 0.020999f
C48 B.n20 VSUBS 0.008556f
C49 B.n21 VSUBS 0.008556f
C50 B.n22 VSUBS 0.008556f
C51 B.n23 VSUBS 0.008556f
C52 B.n24 VSUBS 0.008556f
C53 B.n25 VSUBS 0.008556f
C54 B.n26 VSUBS 0.008556f
C55 B.n27 VSUBS 0.008556f
C56 B.n28 VSUBS 0.008556f
C57 B.n29 VSUBS 0.008556f
C58 B.n30 VSUBS 0.008556f
C59 B.n31 VSUBS 0.008556f
C60 B.n32 VSUBS 0.008556f
C61 B.n33 VSUBS 0.008556f
C62 B.n34 VSUBS 0.008556f
C63 B.n35 VSUBS 0.008556f
C64 B.n36 VSUBS 0.008556f
C65 B.n37 VSUBS 0.008556f
C66 B.n38 VSUBS 0.008556f
C67 B.n39 VSUBS 0.008556f
C68 B.n40 VSUBS 0.008556f
C69 B.n41 VSUBS 0.008556f
C70 B.n42 VSUBS 0.008556f
C71 B.n43 VSUBS 0.008556f
C72 B.n44 VSUBS 0.008556f
C73 B.n45 VSUBS 0.008556f
C74 B.n46 VSUBS 0.008556f
C75 B.n47 VSUBS 0.008556f
C76 B.t7 VSUBS 0.707435f
C77 B.t8 VSUBS 0.722292f
C78 B.t6 VSUBS 1.08638f
C79 B.n48 VSUBS 0.288656f
C80 B.n49 VSUBS 0.081149f
C81 B.n50 VSUBS 0.019823f
C82 B.n51 VSUBS 0.008556f
C83 B.n52 VSUBS 0.008556f
C84 B.n53 VSUBS 0.008556f
C85 B.n54 VSUBS 0.008556f
C86 B.n55 VSUBS 0.008556f
C87 B.t4 VSUBS 0.707411f
C88 B.t5 VSUBS 0.722271f
C89 B.t3 VSUBS 1.08638f
C90 B.n56 VSUBS 0.288677f
C91 B.n57 VSUBS 0.081173f
C92 B.n58 VSUBS 0.008556f
C93 B.n59 VSUBS 0.008556f
C94 B.n60 VSUBS 0.008556f
C95 B.n61 VSUBS 0.008556f
C96 B.n62 VSUBS 0.008556f
C97 B.n63 VSUBS 0.008556f
C98 B.n64 VSUBS 0.008556f
C99 B.n65 VSUBS 0.008556f
C100 B.n66 VSUBS 0.008556f
C101 B.n67 VSUBS 0.008556f
C102 B.n68 VSUBS 0.008556f
C103 B.n69 VSUBS 0.008556f
C104 B.n70 VSUBS 0.008556f
C105 B.n71 VSUBS 0.008556f
C106 B.n72 VSUBS 0.008556f
C107 B.n73 VSUBS 0.008556f
C108 B.n74 VSUBS 0.008556f
C109 B.n75 VSUBS 0.008556f
C110 B.n76 VSUBS 0.008556f
C111 B.n77 VSUBS 0.008556f
C112 B.n78 VSUBS 0.008556f
C113 B.n79 VSUBS 0.008556f
C114 B.n80 VSUBS 0.008556f
C115 B.n81 VSUBS 0.008556f
C116 B.n82 VSUBS 0.008556f
C117 B.n83 VSUBS 0.008556f
C118 B.n84 VSUBS 0.008556f
C119 B.n85 VSUBS 0.02178f
C120 B.n86 VSUBS 0.008556f
C121 B.n87 VSUBS 0.008556f
C122 B.n88 VSUBS 0.008556f
C123 B.n89 VSUBS 0.008556f
C124 B.n90 VSUBS 0.008556f
C125 B.n91 VSUBS 0.008556f
C126 B.n92 VSUBS 0.008556f
C127 B.n93 VSUBS 0.008556f
C128 B.n94 VSUBS 0.008556f
C129 B.n95 VSUBS 0.008556f
C130 B.n96 VSUBS 0.008556f
C131 B.n97 VSUBS 0.008556f
C132 B.n98 VSUBS 0.008556f
C133 B.n99 VSUBS 0.008556f
C134 B.n100 VSUBS 0.008556f
C135 B.n101 VSUBS 0.008556f
C136 B.n102 VSUBS 0.008556f
C137 B.n103 VSUBS 0.008556f
C138 B.n104 VSUBS 0.008556f
C139 B.n105 VSUBS 0.008556f
C140 B.n106 VSUBS 0.008556f
C141 B.n107 VSUBS 0.008556f
C142 B.n108 VSUBS 0.008556f
C143 B.n109 VSUBS 0.008556f
C144 B.n110 VSUBS 0.008556f
C145 B.n111 VSUBS 0.008556f
C146 B.n112 VSUBS 0.008556f
C147 B.n113 VSUBS 0.008556f
C148 B.n114 VSUBS 0.008556f
C149 B.n115 VSUBS 0.008556f
C150 B.n116 VSUBS 0.008556f
C151 B.n117 VSUBS 0.008556f
C152 B.n118 VSUBS 0.008556f
C153 B.n119 VSUBS 0.008556f
C154 B.n120 VSUBS 0.008556f
C155 B.n121 VSUBS 0.020999f
C156 B.n122 VSUBS 0.008556f
C157 B.n123 VSUBS 0.008556f
C158 B.n124 VSUBS 0.008556f
C159 B.n125 VSUBS 0.008556f
C160 B.n126 VSUBS 0.008556f
C161 B.n127 VSUBS 0.008556f
C162 B.n128 VSUBS 0.008556f
C163 B.n129 VSUBS 0.008556f
C164 B.n130 VSUBS 0.008556f
C165 B.n131 VSUBS 0.008556f
C166 B.n132 VSUBS 0.008556f
C167 B.n133 VSUBS 0.008556f
C168 B.n134 VSUBS 0.008556f
C169 B.n135 VSUBS 0.008556f
C170 B.n136 VSUBS 0.008556f
C171 B.n137 VSUBS 0.008556f
C172 B.n138 VSUBS 0.008556f
C173 B.n139 VSUBS 0.008556f
C174 B.n140 VSUBS 0.008556f
C175 B.n141 VSUBS 0.008556f
C176 B.n142 VSUBS 0.008556f
C177 B.n143 VSUBS 0.008556f
C178 B.n144 VSUBS 0.008556f
C179 B.n145 VSUBS 0.008556f
C180 B.n146 VSUBS 0.008556f
C181 B.n147 VSUBS 0.008556f
C182 B.n148 VSUBS 0.008556f
C183 B.n149 VSUBS 0.008556f
C184 B.t2 VSUBS 0.707411f
C185 B.t1 VSUBS 0.722271f
C186 B.t0 VSUBS 1.08638f
C187 B.n150 VSUBS 0.288677f
C188 B.n151 VSUBS 0.081173f
C189 B.n152 VSUBS 0.019823f
C190 B.n153 VSUBS 0.008556f
C191 B.n154 VSUBS 0.008556f
C192 B.n155 VSUBS 0.008556f
C193 B.n156 VSUBS 0.008556f
C194 B.n157 VSUBS 0.008556f
C195 B.t11 VSUBS 0.707435f
C196 B.t10 VSUBS 0.722292f
C197 B.t9 VSUBS 1.08638f
C198 B.n158 VSUBS 0.288656f
C199 B.n159 VSUBS 0.081149f
C200 B.n160 VSUBS 0.008556f
C201 B.n161 VSUBS 0.008556f
C202 B.n162 VSUBS 0.008556f
C203 B.n163 VSUBS 0.008556f
C204 B.n164 VSUBS 0.008556f
C205 B.n165 VSUBS 0.008556f
C206 B.n166 VSUBS 0.008556f
C207 B.n167 VSUBS 0.008556f
C208 B.n168 VSUBS 0.008556f
C209 B.n169 VSUBS 0.008556f
C210 B.n170 VSUBS 0.008556f
C211 B.n171 VSUBS 0.008556f
C212 B.n172 VSUBS 0.008556f
C213 B.n173 VSUBS 0.008556f
C214 B.n174 VSUBS 0.008556f
C215 B.n175 VSUBS 0.008556f
C216 B.n176 VSUBS 0.008556f
C217 B.n177 VSUBS 0.008556f
C218 B.n178 VSUBS 0.008556f
C219 B.n179 VSUBS 0.008556f
C220 B.n180 VSUBS 0.008556f
C221 B.n181 VSUBS 0.008556f
C222 B.n182 VSUBS 0.008556f
C223 B.n183 VSUBS 0.008556f
C224 B.n184 VSUBS 0.008556f
C225 B.n185 VSUBS 0.008556f
C226 B.n186 VSUBS 0.008556f
C227 B.n187 VSUBS 0.02178f
C228 B.n188 VSUBS 0.008556f
C229 B.n189 VSUBS 0.008556f
C230 B.n190 VSUBS 0.008556f
C231 B.n191 VSUBS 0.008556f
C232 B.n192 VSUBS 0.008556f
C233 B.n193 VSUBS 0.008556f
C234 B.n194 VSUBS 0.008556f
C235 B.n195 VSUBS 0.008556f
C236 B.n196 VSUBS 0.008556f
C237 B.n197 VSUBS 0.008556f
C238 B.n198 VSUBS 0.008556f
C239 B.n199 VSUBS 0.008556f
C240 B.n200 VSUBS 0.008556f
C241 B.n201 VSUBS 0.008556f
C242 B.n202 VSUBS 0.008556f
C243 B.n203 VSUBS 0.008556f
C244 B.n204 VSUBS 0.008556f
C245 B.n205 VSUBS 0.008556f
C246 B.n206 VSUBS 0.008556f
C247 B.n207 VSUBS 0.008556f
C248 B.n208 VSUBS 0.008556f
C249 B.n209 VSUBS 0.008556f
C250 B.n210 VSUBS 0.008556f
C251 B.n211 VSUBS 0.008556f
C252 B.n212 VSUBS 0.008556f
C253 B.n213 VSUBS 0.008556f
C254 B.n214 VSUBS 0.008556f
C255 B.n215 VSUBS 0.008556f
C256 B.n216 VSUBS 0.008556f
C257 B.n217 VSUBS 0.008556f
C258 B.n218 VSUBS 0.008556f
C259 B.n219 VSUBS 0.008556f
C260 B.n220 VSUBS 0.008556f
C261 B.n221 VSUBS 0.008556f
C262 B.n222 VSUBS 0.008556f
C263 B.n223 VSUBS 0.008556f
C264 B.n224 VSUBS 0.008556f
C265 B.n225 VSUBS 0.008556f
C266 B.n226 VSUBS 0.008556f
C267 B.n227 VSUBS 0.008556f
C268 B.n228 VSUBS 0.008556f
C269 B.n229 VSUBS 0.008556f
C270 B.n230 VSUBS 0.008556f
C271 B.n231 VSUBS 0.008556f
C272 B.n232 VSUBS 0.008556f
C273 B.n233 VSUBS 0.008556f
C274 B.n234 VSUBS 0.008556f
C275 B.n235 VSUBS 0.008556f
C276 B.n236 VSUBS 0.008556f
C277 B.n237 VSUBS 0.008556f
C278 B.n238 VSUBS 0.008556f
C279 B.n239 VSUBS 0.008556f
C280 B.n240 VSUBS 0.008556f
C281 B.n241 VSUBS 0.008556f
C282 B.n242 VSUBS 0.008556f
C283 B.n243 VSUBS 0.008556f
C284 B.n244 VSUBS 0.008556f
C285 B.n245 VSUBS 0.008556f
C286 B.n246 VSUBS 0.008556f
C287 B.n247 VSUBS 0.008556f
C288 B.n248 VSUBS 0.008556f
C289 B.n249 VSUBS 0.008556f
C290 B.n250 VSUBS 0.008556f
C291 B.n251 VSUBS 0.008556f
C292 B.n252 VSUBS 0.008556f
C293 B.n253 VSUBS 0.008556f
C294 B.n254 VSUBS 0.020999f
C295 B.n255 VSUBS 0.020999f
C296 B.n256 VSUBS 0.02178f
C297 B.n257 VSUBS 0.008556f
C298 B.n258 VSUBS 0.008556f
C299 B.n259 VSUBS 0.008556f
C300 B.n260 VSUBS 0.008556f
C301 B.n261 VSUBS 0.008556f
C302 B.n262 VSUBS 0.008556f
C303 B.n263 VSUBS 0.008556f
C304 B.n264 VSUBS 0.008556f
C305 B.n265 VSUBS 0.008556f
C306 B.n266 VSUBS 0.008556f
C307 B.n267 VSUBS 0.008556f
C308 B.n268 VSUBS 0.008556f
C309 B.n269 VSUBS 0.008556f
C310 B.n270 VSUBS 0.008556f
C311 B.n271 VSUBS 0.008556f
C312 B.n272 VSUBS 0.008556f
C313 B.n273 VSUBS 0.008556f
C314 B.n274 VSUBS 0.008556f
C315 B.n275 VSUBS 0.008556f
C316 B.n276 VSUBS 0.008556f
C317 B.n277 VSUBS 0.008556f
C318 B.n278 VSUBS 0.008556f
C319 B.n279 VSUBS 0.008556f
C320 B.n280 VSUBS 0.008556f
C321 B.n281 VSUBS 0.008556f
C322 B.n282 VSUBS 0.008556f
C323 B.n283 VSUBS 0.008556f
C324 B.n284 VSUBS 0.008556f
C325 B.n285 VSUBS 0.008556f
C326 B.n286 VSUBS 0.008556f
C327 B.n287 VSUBS 0.008556f
C328 B.n288 VSUBS 0.008556f
C329 B.n289 VSUBS 0.008556f
C330 B.n290 VSUBS 0.008556f
C331 B.n291 VSUBS 0.008556f
C332 B.n292 VSUBS 0.008556f
C333 B.n293 VSUBS 0.008556f
C334 B.n294 VSUBS 0.008556f
C335 B.n295 VSUBS 0.008556f
C336 B.n296 VSUBS 0.008556f
C337 B.n297 VSUBS 0.008556f
C338 B.n298 VSUBS 0.008556f
C339 B.n299 VSUBS 0.008556f
C340 B.n300 VSUBS 0.008556f
C341 B.n301 VSUBS 0.008556f
C342 B.n302 VSUBS 0.008556f
C343 B.n303 VSUBS 0.008556f
C344 B.n304 VSUBS 0.008556f
C345 B.n305 VSUBS 0.008556f
C346 B.n306 VSUBS 0.008556f
C347 B.n307 VSUBS 0.008556f
C348 B.n308 VSUBS 0.008556f
C349 B.n309 VSUBS 0.008556f
C350 B.n310 VSUBS 0.008556f
C351 B.n311 VSUBS 0.008556f
C352 B.n312 VSUBS 0.008556f
C353 B.n313 VSUBS 0.008556f
C354 B.n314 VSUBS 0.008556f
C355 B.n315 VSUBS 0.008556f
C356 B.n316 VSUBS 0.008556f
C357 B.n317 VSUBS 0.008556f
C358 B.n318 VSUBS 0.008556f
C359 B.n319 VSUBS 0.008556f
C360 B.n320 VSUBS 0.008556f
C361 B.n321 VSUBS 0.008556f
C362 B.n322 VSUBS 0.008556f
C363 B.n323 VSUBS 0.008556f
C364 B.n324 VSUBS 0.008556f
C365 B.n325 VSUBS 0.008556f
C366 B.n326 VSUBS 0.008556f
C367 B.n327 VSUBS 0.008556f
C368 B.n328 VSUBS 0.008556f
C369 B.n329 VSUBS 0.008556f
C370 B.n330 VSUBS 0.008556f
C371 B.n331 VSUBS 0.008556f
C372 B.n332 VSUBS 0.008556f
C373 B.n333 VSUBS 0.008556f
C374 B.n334 VSUBS 0.008556f
C375 B.n335 VSUBS 0.008556f
C376 B.n336 VSUBS 0.008556f
C377 B.n337 VSUBS 0.008556f
C378 B.n338 VSUBS 0.008556f
C379 B.n339 VSUBS 0.008556f
C380 B.n340 VSUBS 0.005914f
C381 B.n341 VSUBS 0.019823f
C382 B.n342 VSUBS 0.00692f
C383 B.n343 VSUBS 0.008556f
C384 B.n344 VSUBS 0.008556f
C385 B.n345 VSUBS 0.008556f
C386 B.n346 VSUBS 0.008556f
C387 B.n347 VSUBS 0.008556f
C388 B.n348 VSUBS 0.008556f
C389 B.n349 VSUBS 0.008556f
C390 B.n350 VSUBS 0.008556f
C391 B.n351 VSUBS 0.008556f
C392 B.n352 VSUBS 0.008556f
C393 B.n353 VSUBS 0.008556f
C394 B.n354 VSUBS 0.00692f
C395 B.n355 VSUBS 0.008556f
C396 B.n356 VSUBS 0.008556f
C397 B.n357 VSUBS 0.005914f
C398 B.n358 VSUBS 0.008556f
C399 B.n359 VSUBS 0.008556f
C400 B.n360 VSUBS 0.008556f
C401 B.n361 VSUBS 0.008556f
C402 B.n362 VSUBS 0.008556f
C403 B.n363 VSUBS 0.008556f
C404 B.n364 VSUBS 0.008556f
C405 B.n365 VSUBS 0.008556f
C406 B.n366 VSUBS 0.008556f
C407 B.n367 VSUBS 0.008556f
C408 B.n368 VSUBS 0.008556f
C409 B.n369 VSUBS 0.008556f
C410 B.n370 VSUBS 0.008556f
C411 B.n371 VSUBS 0.008556f
C412 B.n372 VSUBS 0.008556f
C413 B.n373 VSUBS 0.008556f
C414 B.n374 VSUBS 0.008556f
C415 B.n375 VSUBS 0.008556f
C416 B.n376 VSUBS 0.008556f
C417 B.n377 VSUBS 0.008556f
C418 B.n378 VSUBS 0.008556f
C419 B.n379 VSUBS 0.008556f
C420 B.n380 VSUBS 0.008556f
C421 B.n381 VSUBS 0.008556f
C422 B.n382 VSUBS 0.008556f
C423 B.n383 VSUBS 0.008556f
C424 B.n384 VSUBS 0.008556f
C425 B.n385 VSUBS 0.008556f
C426 B.n386 VSUBS 0.008556f
C427 B.n387 VSUBS 0.008556f
C428 B.n388 VSUBS 0.008556f
C429 B.n389 VSUBS 0.008556f
C430 B.n390 VSUBS 0.008556f
C431 B.n391 VSUBS 0.008556f
C432 B.n392 VSUBS 0.008556f
C433 B.n393 VSUBS 0.008556f
C434 B.n394 VSUBS 0.008556f
C435 B.n395 VSUBS 0.008556f
C436 B.n396 VSUBS 0.008556f
C437 B.n397 VSUBS 0.008556f
C438 B.n398 VSUBS 0.008556f
C439 B.n399 VSUBS 0.008556f
C440 B.n400 VSUBS 0.008556f
C441 B.n401 VSUBS 0.008556f
C442 B.n402 VSUBS 0.008556f
C443 B.n403 VSUBS 0.008556f
C444 B.n404 VSUBS 0.008556f
C445 B.n405 VSUBS 0.008556f
C446 B.n406 VSUBS 0.008556f
C447 B.n407 VSUBS 0.008556f
C448 B.n408 VSUBS 0.008556f
C449 B.n409 VSUBS 0.008556f
C450 B.n410 VSUBS 0.008556f
C451 B.n411 VSUBS 0.008556f
C452 B.n412 VSUBS 0.008556f
C453 B.n413 VSUBS 0.008556f
C454 B.n414 VSUBS 0.008556f
C455 B.n415 VSUBS 0.008556f
C456 B.n416 VSUBS 0.008556f
C457 B.n417 VSUBS 0.008556f
C458 B.n418 VSUBS 0.008556f
C459 B.n419 VSUBS 0.008556f
C460 B.n420 VSUBS 0.008556f
C461 B.n421 VSUBS 0.008556f
C462 B.n422 VSUBS 0.008556f
C463 B.n423 VSUBS 0.008556f
C464 B.n424 VSUBS 0.008556f
C465 B.n425 VSUBS 0.008556f
C466 B.n426 VSUBS 0.008556f
C467 B.n427 VSUBS 0.008556f
C468 B.n428 VSUBS 0.008556f
C469 B.n429 VSUBS 0.008556f
C470 B.n430 VSUBS 0.008556f
C471 B.n431 VSUBS 0.008556f
C472 B.n432 VSUBS 0.008556f
C473 B.n433 VSUBS 0.008556f
C474 B.n434 VSUBS 0.008556f
C475 B.n435 VSUBS 0.008556f
C476 B.n436 VSUBS 0.008556f
C477 B.n437 VSUBS 0.008556f
C478 B.n438 VSUBS 0.008556f
C479 B.n439 VSUBS 0.008556f
C480 B.n440 VSUBS 0.02178f
C481 B.n441 VSUBS 0.020865f
C482 B.n442 VSUBS 0.021914f
C483 B.n443 VSUBS 0.008556f
C484 B.n444 VSUBS 0.008556f
C485 B.n445 VSUBS 0.008556f
C486 B.n446 VSUBS 0.008556f
C487 B.n447 VSUBS 0.008556f
C488 B.n448 VSUBS 0.008556f
C489 B.n449 VSUBS 0.008556f
C490 B.n450 VSUBS 0.008556f
C491 B.n451 VSUBS 0.008556f
C492 B.n452 VSUBS 0.008556f
C493 B.n453 VSUBS 0.008556f
C494 B.n454 VSUBS 0.008556f
C495 B.n455 VSUBS 0.008556f
C496 B.n456 VSUBS 0.008556f
C497 B.n457 VSUBS 0.008556f
C498 B.n458 VSUBS 0.008556f
C499 B.n459 VSUBS 0.008556f
C500 B.n460 VSUBS 0.008556f
C501 B.n461 VSUBS 0.008556f
C502 B.n462 VSUBS 0.008556f
C503 B.n463 VSUBS 0.008556f
C504 B.n464 VSUBS 0.008556f
C505 B.n465 VSUBS 0.008556f
C506 B.n466 VSUBS 0.008556f
C507 B.n467 VSUBS 0.008556f
C508 B.n468 VSUBS 0.008556f
C509 B.n469 VSUBS 0.008556f
C510 B.n470 VSUBS 0.008556f
C511 B.n471 VSUBS 0.008556f
C512 B.n472 VSUBS 0.008556f
C513 B.n473 VSUBS 0.008556f
C514 B.n474 VSUBS 0.008556f
C515 B.n475 VSUBS 0.008556f
C516 B.n476 VSUBS 0.008556f
C517 B.n477 VSUBS 0.008556f
C518 B.n478 VSUBS 0.008556f
C519 B.n479 VSUBS 0.008556f
C520 B.n480 VSUBS 0.008556f
C521 B.n481 VSUBS 0.008556f
C522 B.n482 VSUBS 0.008556f
C523 B.n483 VSUBS 0.008556f
C524 B.n484 VSUBS 0.008556f
C525 B.n485 VSUBS 0.008556f
C526 B.n486 VSUBS 0.008556f
C527 B.n487 VSUBS 0.008556f
C528 B.n488 VSUBS 0.008556f
C529 B.n489 VSUBS 0.008556f
C530 B.n490 VSUBS 0.008556f
C531 B.n491 VSUBS 0.008556f
C532 B.n492 VSUBS 0.008556f
C533 B.n493 VSUBS 0.008556f
C534 B.n494 VSUBS 0.008556f
C535 B.n495 VSUBS 0.008556f
C536 B.n496 VSUBS 0.008556f
C537 B.n497 VSUBS 0.008556f
C538 B.n498 VSUBS 0.008556f
C539 B.n499 VSUBS 0.008556f
C540 B.n500 VSUBS 0.008556f
C541 B.n501 VSUBS 0.008556f
C542 B.n502 VSUBS 0.008556f
C543 B.n503 VSUBS 0.008556f
C544 B.n504 VSUBS 0.008556f
C545 B.n505 VSUBS 0.008556f
C546 B.n506 VSUBS 0.008556f
C547 B.n507 VSUBS 0.008556f
C548 B.n508 VSUBS 0.008556f
C549 B.n509 VSUBS 0.008556f
C550 B.n510 VSUBS 0.008556f
C551 B.n511 VSUBS 0.008556f
C552 B.n512 VSUBS 0.008556f
C553 B.n513 VSUBS 0.008556f
C554 B.n514 VSUBS 0.008556f
C555 B.n515 VSUBS 0.008556f
C556 B.n516 VSUBS 0.008556f
C557 B.n517 VSUBS 0.008556f
C558 B.n518 VSUBS 0.008556f
C559 B.n519 VSUBS 0.008556f
C560 B.n520 VSUBS 0.008556f
C561 B.n521 VSUBS 0.008556f
C562 B.n522 VSUBS 0.008556f
C563 B.n523 VSUBS 0.008556f
C564 B.n524 VSUBS 0.008556f
C565 B.n525 VSUBS 0.008556f
C566 B.n526 VSUBS 0.008556f
C567 B.n527 VSUBS 0.008556f
C568 B.n528 VSUBS 0.008556f
C569 B.n529 VSUBS 0.008556f
C570 B.n530 VSUBS 0.008556f
C571 B.n531 VSUBS 0.008556f
C572 B.n532 VSUBS 0.008556f
C573 B.n533 VSUBS 0.008556f
C574 B.n534 VSUBS 0.008556f
C575 B.n535 VSUBS 0.008556f
C576 B.n536 VSUBS 0.008556f
C577 B.n537 VSUBS 0.008556f
C578 B.n538 VSUBS 0.008556f
C579 B.n539 VSUBS 0.008556f
C580 B.n540 VSUBS 0.008556f
C581 B.n541 VSUBS 0.008556f
C582 B.n542 VSUBS 0.008556f
C583 B.n543 VSUBS 0.008556f
C584 B.n544 VSUBS 0.008556f
C585 B.n545 VSUBS 0.008556f
C586 B.n546 VSUBS 0.008556f
C587 B.n547 VSUBS 0.008556f
C588 B.n548 VSUBS 0.020999f
C589 B.n549 VSUBS 0.020999f
C590 B.n550 VSUBS 0.02178f
C591 B.n551 VSUBS 0.008556f
C592 B.n552 VSUBS 0.008556f
C593 B.n553 VSUBS 0.008556f
C594 B.n554 VSUBS 0.008556f
C595 B.n555 VSUBS 0.008556f
C596 B.n556 VSUBS 0.008556f
C597 B.n557 VSUBS 0.008556f
C598 B.n558 VSUBS 0.008556f
C599 B.n559 VSUBS 0.008556f
C600 B.n560 VSUBS 0.008556f
C601 B.n561 VSUBS 0.008556f
C602 B.n562 VSUBS 0.008556f
C603 B.n563 VSUBS 0.008556f
C604 B.n564 VSUBS 0.008556f
C605 B.n565 VSUBS 0.008556f
C606 B.n566 VSUBS 0.008556f
C607 B.n567 VSUBS 0.008556f
C608 B.n568 VSUBS 0.008556f
C609 B.n569 VSUBS 0.008556f
C610 B.n570 VSUBS 0.008556f
C611 B.n571 VSUBS 0.008556f
C612 B.n572 VSUBS 0.008556f
C613 B.n573 VSUBS 0.008556f
C614 B.n574 VSUBS 0.008556f
C615 B.n575 VSUBS 0.008556f
C616 B.n576 VSUBS 0.008556f
C617 B.n577 VSUBS 0.008556f
C618 B.n578 VSUBS 0.008556f
C619 B.n579 VSUBS 0.008556f
C620 B.n580 VSUBS 0.008556f
C621 B.n581 VSUBS 0.008556f
C622 B.n582 VSUBS 0.008556f
C623 B.n583 VSUBS 0.008556f
C624 B.n584 VSUBS 0.008556f
C625 B.n585 VSUBS 0.008556f
C626 B.n586 VSUBS 0.008556f
C627 B.n587 VSUBS 0.008556f
C628 B.n588 VSUBS 0.008556f
C629 B.n589 VSUBS 0.008556f
C630 B.n590 VSUBS 0.008556f
C631 B.n591 VSUBS 0.008556f
C632 B.n592 VSUBS 0.008556f
C633 B.n593 VSUBS 0.008556f
C634 B.n594 VSUBS 0.008556f
C635 B.n595 VSUBS 0.008556f
C636 B.n596 VSUBS 0.008556f
C637 B.n597 VSUBS 0.008556f
C638 B.n598 VSUBS 0.008556f
C639 B.n599 VSUBS 0.008556f
C640 B.n600 VSUBS 0.008556f
C641 B.n601 VSUBS 0.008556f
C642 B.n602 VSUBS 0.008556f
C643 B.n603 VSUBS 0.008556f
C644 B.n604 VSUBS 0.008556f
C645 B.n605 VSUBS 0.008556f
C646 B.n606 VSUBS 0.008556f
C647 B.n607 VSUBS 0.008556f
C648 B.n608 VSUBS 0.008556f
C649 B.n609 VSUBS 0.008556f
C650 B.n610 VSUBS 0.008556f
C651 B.n611 VSUBS 0.008556f
C652 B.n612 VSUBS 0.008556f
C653 B.n613 VSUBS 0.008556f
C654 B.n614 VSUBS 0.008556f
C655 B.n615 VSUBS 0.008556f
C656 B.n616 VSUBS 0.008556f
C657 B.n617 VSUBS 0.008556f
C658 B.n618 VSUBS 0.008556f
C659 B.n619 VSUBS 0.008556f
C660 B.n620 VSUBS 0.008556f
C661 B.n621 VSUBS 0.008556f
C662 B.n622 VSUBS 0.008556f
C663 B.n623 VSUBS 0.008556f
C664 B.n624 VSUBS 0.008556f
C665 B.n625 VSUBS 0.008556f
C666 B.n626 VSUBS 0.008556f
C667 B.n627 VSUBS 0.008556f
C668 B.n628 VSUBS 0.008556f
C669 B.n629 VSUBS 0.008556f
C670 B.n630 VSUBS 0.008556f
C671 B.n631 VSUBS 0.008556f
C672 B.n632 VSUBS 0.008556f
C673 B.n633 VSUBS 0.008556f
C674 B.n634 VSUBS 0.005914f
C675 B.n635 VSUBS 0.019823f
C676 B.n636 VSUBS 0.00692f
C677 B.n637 VSUBS 0.008556f
C678 B.n638 VSUBS 0.008556f
C679 B.n639 VSUBS 0.008556f
C680 B.n640 VSUBS 0.008556f
C681 B.n641 VSUBS 0.008556f
C682 B.n642 VSUBS 0.008556f
C683 B.n643 VSUBS 0.008556f
C684 B.n644 VSUBS 0.008556f
C685 B.n645 VSUBS 0.008556f
C686 B.n646 VSUBS 0.008556f
C687 B.n647 VSUBS 0.008556f
C688 B.n648 VSUBS 0.00692f
C689 B.n649 VSUBS 0.008556f
C690 B.n650 VSUBS 0.008556f
C691 B.n651 VSUBS 0.005914f
C692 B.n652 VSUBS 0.008556f
C693 B.n653 VSUBS 0.008556f
C694 B.n654 VSUBS 0.008556f
C695 B.n655 VSUBS 0.008556f
C696 B.n656 VSUBS 0.008556f
C697 B.n657 VSUBS 0.008556f
C698 B.n658 VSUBS 0.008556f
C699 B.n659 VSUBS 0.008556f
C700 B.n660 VSUBS 0.008556f
C701 B.n661 VSUBS 0.008556f
C702 B.n662 VSUBS 0.008556f
C703 B.n663 VSUBS 0.008556f
C704 B.n664 VSUBS 0.008556f
C705 B.n665 VSUBS 0.008556f
C706 B.n666 VSUBS 0.008556f
C707 B.n667 VSUBS 0.008556f
C708 B.n668 VSUBS 0.008556f
C709 B.n669 VSUBS 0.008556f
C710 B.n670 VSUBS 0.008556f
C711 B.n671 VSUBS 0.008556f
C712 B.n672 VSUBS 0.008556f
C713 B.n673 VSUBS 0.008556f
C714 B.n674 VSUBS 0.008556f
C715 B.n675 VSUBS 0.008556f
C716 B.n676 VSUBS 0.008556f
C717 B.n677 VSUBS 0.008556f
C718 B.n678 VSUBS 0.008556f
C719 B.n679 VSUBS 0.008556f
C720 B.n680 VSUBS 0.008556f
C721 B.n681 VSUBS 0.008556f
C722 B.n682 VSUBS 0.008556f
C723 B.n683 VSUBS 0.008556f
C724 B.n684 VSUBS 0.008556f
C725 B.n685 VSUBS 0.008556f
C726 B.n686 VSUBS 0.008556f
C727 B.n687 VSUBS 0.008556f
C728 B.n688 VSUBS 0.008556f
C729 B.n689 VSUBS 0.008556f
C730 B.n690 VSUBS 0.008556f
C731 B.n691 VSUBS 0.008556f
C732 B.n692 VSUBS 0.008556f
C733 B.n693 VSUBS 0.008556f
C734 B.n694 VSUBS 0.008556f
C735 B.n695 VSUBS 0.008556f
C736 B.n696 VSUBS 0.008556f
C737 B.n697 VSUBS 0.008556f
C738 B.n698 VSUBS 0.008556f
C739 B.n699 VSUBS 0.008556f
C740 B.n700 VSUBS 0.008556f
C741 B.n701 VSUBS 0.008556f
C742 B.n702 VSUBS 0.008556f
C743 B.n703 VSUBS 0.008556f
C744 B.n704 VSUBS 0.008556f
C745 B.n705 VSUBS 0.008556f
C746 B.n706 VSUBS 0.008556f
C747 B.n707 VSUBS 0.008556f
C748 B.n708 VSUBS 0.008556f
C749 B.n709 VSUBS 0.008556f
C750 B.n710 VSUBS 0.008556f
C751 B.n711 VSUBS 0.008556f
C752 B.n712 VSUBS 0.008556f
C753 B.n713 VSUBS 0.008556f
C754 B.n714 VSUBS 0.008556f
C755 B.n715 VSUBS 0.008556f
C756 B.n716 VSUBS 0.008556f
C757 B.n717 VSUBS 0.008556f
C758 B.n718 VSUBS 0.008556f
C759 B.n719 VSUBS 0.008556f
C760 B.n720 VSUBS 0.008556f
C761 B.n721 VSUBS 0.008556f
C762 B.n722 VSUBS 0.008556f
C763 B.n723 VSUBS 0.008556f
C764 B.n724 VSUBS 0.008556f
C765 B.n725 VSUBS 0.008556f
C766 B.n726 VSUBS 0.008556f
C767 B.n727 VSUBS 0.008556f
C768 B.n728 VSUBS 0.008556f
C769 B.n729 VSUBS 0.008556f
C770 B.n730 VSUBS 0.008556f
C771 B.n731 VSUBS 0.008556f
C772 B.n732 VSUBS 0.008556f
C773 B.n733 VSUBS 0.008556f
C774 B.n734 VSUBS 0.02178f
C775 B.n735 VSUBS 0.02178f
C776 B.n736 VSUBS 0.020999f
C777 B.n737 VSUBS 0.008556f
C778 B.n738 VSUBS 0.008556f
C779 B.n739 VSUBS 0.008556f
C780 B.n740 VSUBS 0.008556f
C781 B.n741 VSUBS 0.008556f
C782 B.n742 VSUBS 0.008556f
C783 B.n743 VSUBS 0.008556f
C784 B.n744 VSUBS 0.008556f
C785 B.n745 VSUBS 0.008556f
C786 B.n746 VSUBS 0.008556f
C787 B.n747 VSUBS 0.008556f
C788 B.n748 VSUBS 0.008556f
C789 B.n749 VSUBS 0.008556f
C790 B.n750 VSUBS 0.008556f
C791 B.n751 VSUBS 0.008556f
C792 B.n752 VSUBS 0.008556f
C793 B.n753 VSUBS 0.008556f
C794 B.n754 VSUBS 0.008556f
C795 B.n755 VSUBS 0.008556f
C796 B.n756 VSUBS 0.008556f
C797 B.n757 VSUBS 0.008556f
C798 B.n758 VSUBS 0.008556f
C799 B.n759 VSUBS 0.008556f
C800 B.n760 VSUBS 0.008556f
C801 B.n761 VSUBS 0.008556f
C802 B.n762 VSUBS 0.008556f
C803 B.n763 VSUBS 0.008556f
C804 B.n764 VSUBS 0.008556f
C805 B.n765 VSUBS 0.008556f
C806 B.n766 VSUBS 0.008556f
C807 B.n767 VSUBS 0.008556f
C808 B.n768 VSUBS 0.008556f
C809 B.n769 VSUBS 0.008556f
C810 B.n770 VSUBS 0.008556f
C811 B.n771 VSUBS 0.008556f
C812 B.n772 VSUBS 0.008556f
C813 B.n773 VSUBS 0.008556f
C814 B.n774 VSUBS 0.008556f
C815 B.n775 VSUBS 0.008556f
C816 B.n776 VSUBS 0.008556f
C817 B.n777 VSUBS 0.008556f
C818 B.n778 VSUBS 0.008556f
C819 B.n779 VSUBS 0.008556f
C820 B.n780 VSUBS 0.008556f
C821 B.n781 VSUBS 0.008556f
C822 B.n782 VSUBS 0.008556f
C823 B.n783 VSUBS 0.008556f
C824 B.n784 VSUBS 0.008556f
C825 B.n785 VSUBS 0.008556f
C826 B.n786 VSUBS 0.008556f
C827 B.n787 VSUBS 0.011165f
C828 B.n788 VSUBS 0.011893f
C829 B.n789 VSUBS 0.023651f
C830 VDD2.t2 VSUBS 3.9549f
C831 VDD2.t4 VSUBS 0.367181f
C832 VDD2.t5 VSUBS 0.367181f
C833 VDD2.n0 VSUBS 3.03623f
C834 VDD2.n1 VSUBS 1.40701f
C835 VDD2.t7 VSUBS 0.367181f
C836 VDD2.t9 VSUBS 0.367181f
C837 VDD2.n2 VSUBS 3.04615f
C838 VDD2.n3 VSUBS 3.01011f
C839 VDD2.t6 VSUBS 3.94113f
C840 VDD2.n4 VSUBS 3.56284f
C841 VDD2.t8 VSUBS 0.367181f
C842 VDD2.t0 VSUBS 0.367181f
C843 VDD2.n5 VSUBS 3.03623f
C844 VDD2.n6 VSUBS 0.677685f
C845 VDD2.t1 VSUBS 0.367181f
C846 VDD2.t3 VSUBS 0.367181f
C847 VDD2.n7 VSUBS 3.0461f
C848 VN.n0 VSUBS 0.051764f
C849 VN.t2 VSUBS 2.25543f
C850 VN.n1 VSUBS 0.80218f
C851 VN.n2 VSUBS 0.038793f
C852 VN.t4 VSUBS 2.25543f
C853 VN.n3 VSUBS 0.80218f
C854 VN.n4 VSUBS 0.038793f
C855 VN.t5 VSUBS 2.25543f
C856 VN.n5 VSUBS 0.854823f
C857 VN.t7 VSUBS 2.37436f
C858 VN.n6 VSUBS 0.864968f
C859 VN.n7 VSUBS 0.203347f
C860 VN.n8 VSUBS 0.061837f
C861 VN.n9 VSUBS 0.031779f
C862 VN.n10 VSUBS 0.059853f
C863 VN.n11 VSUBS 0.038793f
C864 VN.n12 VSUBS 0.038793f
C865 VN.n13 VSUBS 0.059853f
C866 VN.n14 VSUBS 0.031779f
C867 VN.n15 VSUBS 0.061837f
C868 VN.n16 VSUBS 0.038793f
C869 VN.n17 VSUBS 0.038793f
C870 VN.n18 VSUBS 0.055589f
C871 VN.n19 VSUBS 0.029787f
C872 VN.t0 VSUBS 2.32808f
C873 VN.n20 VSUBS 0.876659f
C874 VN.n21 VSUBS 0.036331f
C875 VN.n22 VSUBS 0.051764f
C876 VN.t1 VSUBS 2.25543f
C877 VN.n23 VSUBS 0.80218f
C878 VN.n24 VSUBS 0.038793f
C879 VN.t9 VSUBS 2.25543f
C880 VN.n25 VSUBS 0.80218f
C881 VN.n26 VSUBS 0.038793f
C882 VN.t8 VSUBS 2.25543f
C883 VN.n27 VSUBS 0.854823f
C884 VN.t6 VSUBS 2.37436f
C885 VN.n28 VSUBS 0.864968f
C886 VN.n29 VSUBS 0.203347f
C887 VN.n30 VSUBS 0.061837f
C888 VN.n31 VSUBS 0.031779f
C889 VN.n32 VSUBS 0.059853f
C890 VN.n33 VSUBS 0.038793f
C891 VN.n34 VSUBS 0.038793f
C892 VN.n35 VSUBS 0.059853f
C893 VN.n36 VSUBS 0.031779f
C894 VN.n37 VSUBS 0.061837f
C895 VN.n38 VSUBS 0.038793f
C896 VN.n39 VSUBS 0.038793f
C897 VN.n40 VSUBS 0.055589f
C898 VN.n41 VSUBS 0.029787f
C899 VN.t3 VSUBS 2.32808f
C900 VN.n42 VSUBS 0.876659f
C901 VN.n43 VSUBS 2.13014f
C902 VTAIL.t7 VSUBS 0.370782f
C903 VTAIL.t3 VSUBS 0.370782f
C904 VTAIL.n0 VSUBS 2.90132f
C905 VTAIL.n1 VSUBS 0.85324f
C906 VTAIL.t17 VSUBS 3.79126f
C907 VTAIL.n2 VSUBS 0.998971f
C908 VTAIL.t10 VSUBS 0.370782f
C909 VTAIL.t18 VSUBS 0.370782f
C910 VTAIL.n3 VSUBS 2.90132f
C911 VTAIL.n4 VSUBS 0.895486f
C912 VTAIL.t16 VSUBS 0.370782f
C913 VTAIL.t13 VSUBS 0.370782f
C914 VTAIL.n5 VSUBS 2.90132f
C915 VTAIL.n6 VSUBS 2.68761f
C916 VTAIL.t5 VSUBS 0.370782f
C917 VTAIL.t19 VSUBS 0.370782f
C918 VTAIL.n7 VSUBS 2.90133f
C919 VTAIL.n8 VSUBS 2.68761f
C920 VTAIL.t0 VSUBS 0.370782f
C921 VTAIL.t8 VSUBS 0.370782f
C922 VTAIL.n9 VSUBS 2.90133f
C923 VTAIL.n10 VSUBS 0.89548f
C924 VTAIL.t4 VSUBS 3.79129f
C925 VTAIL.n11 VSUBS 0.998943f
C926 VTAIL.t11 VSUBS 0.370782f
C927 VTAIL.t9 VSUBS 0.370782f
C928 VTAIL.n12 VSUBS 2.90133f
C929 VTAIL.n13 VSUBS 0.877672f
C930 VTAIL.t15 VSUBS 0.370782f
C931 VTAIL.t14 VSUBS 0.370782f
C932 VTAIL.n14 VSUBS 2.90133f
C933 VTAIL.n15 VSUBS 0.89548f
C934 VTAIL.t12 VSUBS 3.79126f
C935 VTAIL.n16 VSUBS 2.6907f
C936 VTAIL.t2 VSUBS 3.79126f
C937 VTAIL.n17 VSUBS 2.6907f
C938 VTAIL.t6 VSUBS 0.370782f
C939 VTAIL.t1 VSUBS 0.370782f
C940 VTAIL.n18 VSUBS 2.90132f
C941 VTAIL.n19 VSUBS 0.801713f
C942 VDD1.t9 VSUBS 3.93068f
C943 VDD1.t5 VSUBS 0.364931f
C944 VDD1.t1 VSUBS 0.364931f
C945 VDD1.n0 VSUBS 3.01763f
C946 VDD1.n1 VSUBS 1.40597f
C947 VDD1.t6 VSUBS 3.93066f
C948 VDD1.t3 VSUBS 0.364931f
C949 VDD1.t8 VSUBS 0.364931f
C950 VDD1.n2 VSUBS 3.01762f
C951 VDD1.n3 VSUBS 1.39839f
C952 VDD1.t4 VSUBS 0.364931f
C953 VDD1.t7 VSUBS 0.364931f
C954 VDD1.n4 VSUBS 3.02748f
C955 VDD1.n5 VSUBS 3.09019f
C956 VDD1.t0 VSUBS 0.364931f
C957 VDD1.t2 VSUBS 0.364931f
C958 VDD1.n6 VSUBS 3.01762f
C959 VDD1.n7 VSUBS 3.52797f
C960 VP.n0 VSUBS 0.052533f
C961 VP.t0 VSUBS 2.28892f
C962 VP.n1 VSUBS 0.814091f
C963 VP.n2 VSUBS 0.039369f
C964 VP.t8 VSUBS 2.28892f
C965 VP.n3 VSUBS 0.814091f
C966 VP.n4 VSUBS 0.039369f
C967 VP.t5 VSUBS 2.28892f
C968 VP.n5 VSUBS 0.814091f
C969 VP.n6 VSUBS 0.052533f
C970 VP.n7 VSUBS 0.052533f
C971 VP.t6 VSUBS 2.36265f
C972 VP.t4 VSUBS 2.28892f
C973 VP.n8 VSUBS 0.814091f
C974 VP.n9 VSUBS 0.039369f
C975 VP.t3 VSUBS 2.28892f
C976 VP.n10 VSUBS 0.814091f
C977 VP.n11 VSUBS 0.039369f
C978 VP.t9 VSUBS 2.28892f
C979 VP.n12 VSUBS 0.867516f
C980 VP.t7 VSUBS 2.40962f
C981 VP.n13 VSUBS 0.877812f
C982 VP.n14 VSUBS 0.206367f
C983 VP.n15 VSUBS 0.062755f
C984 VP.n16 VSUBS 0.032251f
C985 VP.n17 VSUBS 0.060741f
C986 VP.n18 VSUBS 0.039369f
C987 VP.n19 VSUBS 0.039369f
C988 VP.n20 VSUBS 0.060741f
C989 VP.n21 VSUBS 0.032251f
C990 VP.n22 VSUBS 0.062755f
C991 VP.n23 VSUBS 0.039369f
C992 VP.n24 VSUBS 0.039369f
C993 VP.n25 VSUBS 0.056415f
C994 VP.n26 VSUBS 0.030229f
C995 VP.n27 VSUBS 0.889676f
C996 VP.n28 VSUBS 2.14029f
C997 VP.n29 VSUBS 2.1688f
C998 VP.t2 VSUBS 2.36265f
C999 VP.n30 VSUBS 0.889676f
C1000 VP.n31 VSUBS 0.030229f
C1001 VP.n32 VSUBS 0.056415f
C1002 VP.n33 VSUBS 0.039369f
C1003 VP.n34 VSUBS 0.039369f
C1004 VP.n35 VSUBS 0.062755f
C1005 VP.n36 VSUBS 0.032251f
C1006 VP.n37 VSUBS 0.060741f
C1007 VP.n38 VSUBS 0.039369f
C1008 VP.n39 VSUBS 0.039369f
C1009 VP.n40 VSUBS 0.060741f
C1010 VP.n41 VSUBS 0.032251f
C1011 VP.n42 VSUBS 0.062755f
C1012 VP.n43 VSUBS 0.039369f
C1013 VP.n44 VSUBS 0.039369f
C1014 VP.n45 VSUBS 0.056415f
C1015 VP.n46 VSUBS 0.030229f
C1016 VP.t1 VSUBS 2.36265f
C1017 VP.n47 VSUBS 0.889676f
C1018 VP.n48 VSUBS 0.036871f
.ends

