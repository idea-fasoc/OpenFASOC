* NGSPICE file created from diff_pair_sample_0013.ext - technology: sky130A

.subckt diff_pair_sample_0013 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=2.8197 pd=15.24 as=0 ps=0 w=7.23 l=3.92
X1 VDD1.t1 VP.t0 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=2.8197 pd=15.24 as=2.8197 ps=15.24 w=7.23 l=3.92
X2 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=2.8197 pd=15.24 as=0 ps=0 w=7.23 l=3.92
X3 VDD2.t1 VN.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.8197 pd=15.24 as=2.8197 ps=15.24 w=7.23 l=3.92
X4 VDD2.t0 VN.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.8197 pd=15.24 as=2.8197 ps=15.24 w=7.23 l=3.92
X5 VDD1.t0 VP.t1 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=2.8197 pd=15.24 as=2.8197 ps=15.24 w=7.23 l=3.92
X6 B.t8 B.t6 B.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=2.8197 pd=15.24 as=0 ps=0 w=7.23 l=3.92
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=2.8197 pd=15.24 as=0 ps=0 w=7.23 l=3.92
R0 B.n603 B.n602 585
R1 B.n604 B.n603 585
R2 B.n228 B.n95 585
R3 B.n227 B.n226 585
R4 B.n225 B.n224 585
R5 B.n223 B.n222 585
R6 B.n221 B.n220 585
R7 B.n219 B.n218 585
R8 B.n217 B.n216 585
R9 B.n215 B.n214 585
R10 B.n213 B.n212 585
R11 B.n211 B.n210 585
R12 B.n209 B.n208 585
R13 B.n207 B.n206 585
R14 B.n205 B.n204 585
R15 B.n203 B.n202 585
R16 B.n201 B.n200 585
R17 B.n199 B.n198 585
R18 B.n197 B.n196 585
R19 B.n195 B.n194 585
R20 B.n193 B.n192 585
R21 B.n191 B.n190 585
R22 B.n189 B.n188 585
R23 B.n187 B.n186 585
R24 B.n185 B.n184 585
R25 B.n183 B.n182 585
R26 B.n181 B.n180 585
R27 B.n179 B.n178 585
R28 B.n177 B.n176 585
R29 B.n174 B.n173 585
R30 B.n172 B.n171 585
R31 B.n170 B.n169 585
R32 B.n168 B.n167 585
R33 B.n166 B.n165 585
R34 B.n164 B.n163 585
R35 B.n162 B.n161 585
R36 B.n160 B.n159 585
R37 B.n158 B.n157 585
R38 B.n156 B.n155 585
R39 B.n154 B.n153 585
R40 B.n152 B.n151 585
R41 B.n150 B.n149 585
R42 B.n148 B.n147 585
R43 B.n146 B.n145 585
R44 B.n144 B.n143 585
R45 B.n142 B.n141 585
R46 B.n140 B.n139 585
R47 B.n138 B.n137 585
R48 B.n136 B.n135 585
R49 B.n134 B.n133 585
R50 B.n132 B.n131 585
R51 B.n130 B.n129 585
R52 B.n128 B.n127 585
R53 B.n126 B.n125 585
R54 B.n124 B.n123 585
R55 B.n122 B.n121 585
R56 B.n120 B.n119 585
R57 B.n118 B.n117 585
R58 B.n116 B.n115 585
R59 B.n114 B.n113 585
R60 B.n112 B.n111 585
R61 B.n110 B.n109 585
R62 B.n108 B.n107 585
R63 B.n106 B.n105 585
R64 B.n104 B.n103 585
R65 B.n102 B.n101 585
R66 B.n601 B.n62 585
R67 B.n605 B.n62 585
R68 B.n600 B.n61 585
R69 B.n606 B.n61 585
R70 B.n599 B.n598 585
R71 B.n598 B.n57 585
R72 B.n597 B.n56 585
R73 B.n612 B.n56 585
R74 B.n596 B.n55 585
R75 B.n613 B.n55 585
R76 B.n595 B.n54 585
R77 B.n614 B.n54 585
R78 B.n594 B.n593 585
R79 B.n593 B.n50 585
R80 B.n592 B.n49 585
R81 B.n620 B.n49 585
R82 B.n591 B.n48 585
R83 B.n621 B.n48 585
R84 B.n590 B.n47 585
R85 B.n622 B.n47 585
R86 B.n589 B.n588 585
R87 B.n588 B.n43 585
R88 B.n587 B.n42 585
R89 B.n628 B.n42 585
R90 B.n586 B.n41 585
R91 B.n629 B.n41 585
R92 B.n585 B.n40 585
R93 B.n630 B.n40 585
R94 B.n584 B.n583 585
R95 B.n583 B.n36 585
R96 B.n582 B.n35 585
R97 B.n636 B.n35 585
R98 B.n581 B.n34 585
R99 B.n637 B.n34 585
R100 B.n580 B.n33 585
R101 B.n638 B.n33 585
R102 B.n579 B.n578 585
R103 B.n578 B.n29 585
R104 B.n577 B.n28 585
R105 B.n644 B.n28 585
R106 B.n576 B.n27 585
R107 B.n645 B.n27 585
R108 B.n575 B.n26 585
R109 B.n646 B.n26 585
R110 B.n574 B.n573 585
R111 B.n573 B.n22 585
R112 B.n572 B.n21 585
R113 B.n652 B.n21 585
R114 B.n571 B.n20 585
R115 B.n653 B.n20 585
R116 B.n570 B.n19 585
R117 B.n654 B.n19 585
R118 B.n569 B.n568 585
R119 B.n568 B.n15 585
R120 B.n567 B.n14 585
R121 B.n660 B.n14 585
R122 B.n566 B.n13 585
R123 B.n661 B.n13 585
R124 B.n565 B.n12 585
R125 B.n662 B.n12 585
R126 B.n564 B.n563 585
R127 B.n563 B.n8 585
R128 B.n562 B.n7 585
R129 B.n668 B.n7 585
R130 B.n561 B.n6 585
R131 B.n669 B.n6 585
R132 B.n560 B.n5 585
R133 B.n670 B.n5 585
R134 B.n559 B.n558 585
R135 B.n558 B.n4 585
R136 B.n557 B.n229 585
R137 B.n557 B.n556 585
R138 B.n547 B.n230 585
R139 B.n231 B.n230 585
R140 B.n549 B.n548 585
R141 B.n550 B.n549 585
R142 B.n546 B.n236 585
R143 B.n236 B.n235 585
R144 B.n545 B.n544 585
R145 B.n544 B.n543 585
R146 B.n238 B.n237 585
R147 B.n239 B.n238 585
R148 B.n536 B.n535 585
R149 B.n537 B.n536 585
R150 B.n534 B.n244 585
R151 B.n244 B.n243 585
R152 B.n533 B.n532 585
R153 B.n532 B.n531 585
R154 B.n246 B.n245 585
R155 B.n247 B.n246 585
R156 B.n524 B.n523 585
R157 B.n525 B.n524 585
R158 B.n522 B.n252 585
R159 B.n252 B.n251 585
R160 B.n521 B.n520 585
R161 B.n520 B.n519 585
R162 B.n254 B.n253 585
R163 B.n255 B.n254 585
R164 B.n512 B.n511 585
R165 B.n513 B.n512 585
R166 B.n510 B.n260 585
R167 B.n260 B.n259 585
R168 B.n509 B.n508 585
R169 B.n508 B.n507 585
R170 B.n262 B.n261 585
R171 B.n263 B.n262 585
R172 B.n500 B.n499 585
R173 B.n501 B.n500 585
R174 B.n498 B.n268 585
R175 B.n268 B.n267 585
R176 B.n497 B.n496 585
R177 B.n496 B.n495 585
R178 B.n270 B.n269 585
R179 B.n271 B.n270 585
R180 B.n488 B.n487 585
R181 B.n489 B.n488 585
R182 B.n486 B.n276 585
R183 B.n276 B.n275 585
R184 B.n485 B.n484 585
R185 B.n484 B.n483 585
R186 B.n278 B.n277 585
R187 B.n279 B.n278 585
R188 B.n476 B.n475 585
R189 B.n477 B.n476 585
R190 B.n474 B.n284 585
R191 B.n284 B.n283 585
R192 B.n473 B.n472 585
R193 B.n472 B.n471 585
R194 B.n286 B.n285 585
R195 B.n287 B.n286 585
R196 B.n464 B.n463 585
R197 B.n465 B.n464 585
R198 B.n462 B.n292 585
R199 B.n292 B.n291 585
R200 B.n456 B.n455 585
R201 B.n454 B.n326 585
R202 B.n453 B.n325 585
R203 B.n458 B.n325 585
R204 B.n452 B.n451 585
R205 B.n450 B.n449 585
R206 B.n448 B.n447 585
R207 B.n446 B.n445 585
R208 B.n444 B.n443 585
R209 B.n442 B.n441 585
R210 B.n440 B.n439 585
R211 B.n438 B.n437 585
R212 B.n436 B.n435 585
R213 B.n434 B.n433 585
R214 B.n432 B.n431 585
R215 B.n430 B.n429 585
R216 B.n428 B.n427 585
R217 B.n426 B.n425 585
R218 B.n424 B.n423 585
R219 B.n422 B.n421 585
R220 B.n420 B.n419 585
R221 B.n418 B.n417 585
R222 B.n416 B.n415 585
R223 B.n414 B.n413 585
R224 B.n412 B.n411 585
R225 B.n410 B.n409 585
R226 B.n408 B.n407 585
R227 B.n406 B.n405 585
R228 B.n404 B.n403 585
R229 B.n401 B.n400 585
R230 B.n399 B.n398 585
R231 B.n397 B.n396 585
R232 B.n395 B.n394 585
R233 B.n393 B.n392 585
R234 B.n391 B.n390 585
R235 B.n389 B.n388 585
R236 B.n387 B.n386 585
R237 B.n385 B.n384 585
R238 B.n383 B.n382 585
R239 B.n381 B.n380 585
R240 B.n379 B.n378 585
R241 B.n377 B.n376 585
R242 B.n375 B.n374 585
R243 B.n373 B.n372 585
R244 B.n371 B.n370 585
R245 B.n369 B.n368 585
R246 B.n367 B.n366 585
R247 B.n365 B.n364 585
R248 B.n363 B.n362 585
R249 B.n361 B.n360 585
R250 B.n359 B.n358 585
R251 B.n357 B.n356 585
R252 B.n355 B.n354 585
R253 B.n353 B.n352 585
R254 B.n351 B.n350 585
R255 B.n349 B.n348 585
R256 B.n347 B.n346 585
R257 B.n345 B.n344 585
R258 B.n343 B.n342 585
R259 B.n341 B.n340 585
R260 B.n339 B.n338 585
R261 B.n337 B.n336 585
R262 B.n335 B.n334 585
R263 B.n333 B.n332 585
R264 B.n294 B.n293 585
R265 B.n461 B.n460 585
R266 B.n290 B.n289 585
R267 B.n291 B.n290 585
R268 B.n467 B.n466 585
R269 B.n466 B.n465 585
R270 B.n468 B.n288 585
R271 B.n288 B.n287 585
R272 B.n470 B.n469 585
R273 B.n471 B.n470 585
R274 B.n282 B.n281 585
R275 B.n283 B.n282 585
R276 B.n479 B.n478 585
R277 B.n478 B.n477 585
R278 B.n480 B.n280 585
R279 B.n280 B.n279 585
R280 B.n482 B.n481 585
R281 B.n483 B.n482 585
R282 B.n274 B.n273 585
R283 B.n275 B.n274 585
R284 B.n491 B.n490 585
R285 B.n490 B.n489 585
R286 B.n492 B.n272 585
R287 B.n272 B.n271 585
R288 B.n494 B.n493 585
R289 B.n495 B.n494 585
R290 B.n266 B.n265 585
R291 B.n267 B.n266 585
R292 B.n503 B.n502 585
R293 B.n502 B.n501 585
R294 B.n504 B.n264 585
R295 B.n264 B.n263 585
R296 B.n506 B.n505 585
R297 B.n507 B.n506 585
R298 B.n258 B.n257 585
R299 B.n259 B.n258 585
R300 B.n515 B.n514 585
R301 B.n514 B.n513 585
R302 B.n516 B.n256 585
R303 B.n256 B.n255 585
R304 B.n518 B.n517 585
R305 B.n519 B.n518 585
R306 B.n250 B.n249 585
R307 B.n251 B.n250 585
R308 B.n527 B.n526 585
R309 B.n526 B.n525 585
R310 B.n528 B.n248 585
R311 B.n248 B.n247 585
R312 B.n530 B.n529 585
R313 B.n531 B.n530 585
R314 B.n242 B.n241 585
R315 B.n243 B.n242 585
R316 B.n539 B.n538 585
R317 B.n538 B.n537 585
R318 B.n540 B.n240 585
R319 B.n240 B.n239 585
R320 B.n542 B.n541 585
R321 B.n543 B.n542 585
R322 B.n234 B.n233 585
R323 B.n235 B.n234 585
R324 B.n552 B.n551 585
R325 B.n551 B.n550 585
R326 B.n553 B.n232 585
R327 B.n232 B.n231 585
R328 B.n555 B.n554 585
R329 B.n556 B.n555 585
R330 B.n2 B.n0 585
R331 B.n4 B.n2 585
R332 B.n3 B.n1 585
R333 B.n669 B.n3 585
R334 B.n667 B.n666 585
R335 B.n668 B.n667 585
R336 B.n665 B.n9 585
R337 B.n9 B.n8 585
R338 B.n664 B.n663 585
R339 B.n663 B.n662 585
R340 B.n11 B.n10 585
R341 B.n661 B.n11 585
R342 B.n659 B.n658 585
R343 B.n660 B.n659 585
R344 B.n657 B.n16 585
R345 B.n16 B.n15 585
R346 B.n656 B.n655 585
R347 B.n655 B.n654 585
R348 B.n18 B.n17 585
R349 B.n653 B.n18 585
R350 B.n651 B.n650 585
R351 B.n652 B.n651 585
R352 B.n649 B.n23 585
R353 B.n23 B.n22 585
R354 B.n648 B.n647 585
R355 B.n647 B.n646 585
R356 B.n25 B.n24 585
R357 B.n645 B.n25 585
R358 B.n643 B.n642 585
R359 B.n644 B.n643 585
R360 B.n641 B.n30 585
R361 B.n30 B.n29 585
R362 B.n640 B.n639 585
R363 B.n639 B.n638 585
R364 B.n32 B.n31 585
R365 B.n637 B.n32 585
R366 B.n635 B.n634 585
R367 B.n636 B.n635 585
R368 B.n633 B.n37 585
R369 B.n37 B.n36 585
R370 B.n632 B.n631 585
R371 B.n631 B.n630 585
R372 B.n39 B.n38 585
R373 B.n629 B.n39 585
R374 B.n627 B.n626 585
R375 B.n628 B.n627 585
R376 B.n625 B.n44 585
R377 B.n44 B.n43 585
R378 B.n624 B.n623 585
R379 B.n623 B.n622 585
R380 B.n46 B.n45 585
R381 B.n621 B.n46 585
R382 B.n619 B.n618 585
R383 B.n620 B.n619 585
R384 B.n617 B.n51 585
R385 B.n51 B.n50 585
R386 B.n616 B.n615 585
R387 B.n615 B.n614 585
R388 B.n53 B.n52 585
R389 B.n613 B.n53 585
R390 B.n611 B.n610 585
R391 B.n612 B.n611 585
R392 B.n609 B.n58 585
R393 B.n58 B.n57 585
R394 B.n608 B.n607 585
R395 B.n607 B.n606 585
R396 B.n60 B.n59 585
R397 B.n605 B.n60 585
R398 B.n672 B.n671 585
R399 B.n671 B.n670 585
R400 B.n456 B.n290 497.305
R401 B.n101 B.n60 497.305
R402 B.n460 B.n292 497.305
R403 B.n603 B.n62 497.305
R404 B.n329 B.t5 282.264
R405 B.n96 B.t11 282.264
R406 B.n327 B.t8 282.264
R407 B.n98 B.t14 282.264
R408 B.n604 B.n94 256.663
R409 B.n604 B.n93 256.663
R410 B.n604 B.n92 256.663
R411 B.n604 B.n91 256.663
R412 B.n604 B.n90 256.663
R413 B.n604 B.n89 256.663
R414 B.n604 B.n88 256.663
R415 B.n604 B.n87 256.663
R416 B.n604 B.n86 256.663
R417 B.n604 B.n85 256.663
R418 B.n604 B.n84 256.663
R419 B.n604 B.n83 256.663
R420 B.n604 B.n82 256.663
R421 B.n604 B.n81 256.663
R422 B.n604 B.n80 256.663
R423 B.n604 B.n79 256.663
R424 B.n604 B.n78 256.663
R425 B.n604 B.n77 256.663
R426 B.n604 B.n76 256.663
R427 B.n604 B.n75 256.663
R428 B.n604 B.n74 256.663
R429 B.n604 B.n73 256.663
R430 B.n604 B.n72 256.663
R431 B.n604 B.n71 256.663
R432 B.n604 B.n70 256.663
R433 B.n604 B.n69 256.663
R434 B.n604 B.n68 256.663
R435 B.n604 B.n67 256.663
R436 B.n604 B.n66 256.663
R437 B.n604 B.n65 256.663
R438 B.n604 B.n64 256.663
R439 B.n604 B.n63 256.663
R440 B.n458 B.n457 256.663
R441 B.n458 B.n295 256.663
R442 B.n458 B.n296 256.663
R443 B.n458 B.n297 256.663
R444 B.n458 B.n298 256.663
R445 B.n458 B.n299 256.663
R446 B.n458 B.n300 256.663
R447 B.n458 B.n301 256.663
R448 B.n458 B.n302 256.663
R449 B.n458 B.n303 256.663
R450 B.n458 B.n304 256.663
R451 B.n458 B.n305 256.663
R452 B.n458 B.n306 256.663
R453 B.n458 B.n307 256.663
R454 B.n458 B.n308 256.663
R455 B.n458 B.n309 256.663
R456 B.n458 B.n310 256.663
R457 B.n458 B.n311 256.663
R458 B.n458 B.n312 256.663
R459 B.n458 B.n313 256.663
R460 B.n458 B.n314 256.663
R461 B.n458 B.n315 256.663
R462 B.n458 B.n316 256.663
R463 B.n458 B.n317 256.663
R464 B.n458 B.n318 256.663
R465 B.n458 B.n319 256.663
R466 B.n458 B.n320 256.663
R467 B.n458 B.n321 256.663
R468 B.n458 B.n322 256.663
R469 B.n458 B.n323 256.663
R470 B.n458 B.n324 256.663
R471 B.n459 B.n458 256.663
R472 B.n329 B.t2 253.883
R473 B.n327 B.t6 253.883
R474 B.n98 B.t13 253.883
R475 B.n96 B.t9 253.883
R476 B.n330 B.t4 199.84
R477 B.n97 B.t12 199.84
R478 B.n328 B.t7 199.84
R479 B.n99 B.t15 199.84
R480 B.n466 B.n290 163.367
R481 B.n466 B.n288 163.367
R482 B.n470 B.n288 163.367
R483 B.n470 B.n282 163.367
R484 B.n478 B.n282 163.367
R485 B.n478 B.n280 163.367
R486 B.n482 B.n280 163.367
R487 B.n482 B.n274 163.367
R488 B.n490 B.n274 163.367
R489 B.n490 B.n272 163.367
R490 B.n494 B.n272 163.367
R491 B.n494 B.n266 163.367
R492 B.n502 B.n266 163.367
R493 B.n502 B.n264 163.367
R494 B.n506 B.n264 163.367
R495 B.n506 B.n258 163.367
R496 B.n514 B.n258 163.367
R497 B.n514 B.n256 163.367
R498 B.n518 B.n256 163.367
R499 B.n518 B.n250 163.367
R500 B.n526 B.n250 163.367
R501 B.n526 B.n248 163.367
R502 B.n530 B.n248 163.367
R503 B.n530 B.n242 163.367
R504 B.n538 B.n242 163.367
R505 B.n538 B.n240 163.367
R506 B.n542 B.n240 163.367
R507 B.n542 B.n234 163.367
R508 B.n551 B.n234 163.367
R509 B.n551 B.n232 163.367
R510 B.n555 B.n232 163.367
R511 B.n555 B.n2 163.367
R512 B.n671 B.n2 163.367
R513 B.n671 B.n3 163.367
R514 B.n667 B.n3 163.367
R515 B.n667 B.n9 163.367
R516 B.n663 B.n9 163.367
R517 B.n663 B.n11 163.367
R518 B.n659 B.n11 163.367
R519 B.n659 B.n16 163.367
R520 B.n655 B.n16 163.367
R521 B.n655 B.n18 163.367
R522 B.n651 B.n18 163.367
R523 B.n651 B.n23 163.367
R524 B.n647 B.n23 163.367
R525 B.n647 B.n25 163.367
R526 B.n643 B.n25 163.367
R527 B.n643 B.n30 163.367
R528 B.n639 B.n30 163.367
R529 B.n639 B.n32 163.367
R530 B.n635 B.n32 163.367
R531 B.n635 B.n37 163.367
R532 B.n631 B.n37 163.367
R533 B.n631 B.n39 163.367
R534 B.n627 B.n39 163.367
R535 B.n627 B.n44 163.367
R536 B.n623 B.n44 163.367
R537 B.n623 B.n46 163.367
R538 B.n619 B.n46 163.367
R539 B.n619 B.n51 163.367
R540 B.n615 B.n51 163.367
R541 B.n615 B.n53 163.367
R542 B.n611 B.n53 163.367
R543 B.n611 B.n58 163.367
R544 B.n607 B.n58 163.367
R545 B.n607 B.n60 163.367
R546 B.n326 B.n325 163.367
R547 B.n451 B.n325 163.367
R548 B.n449 B.n448 163.367
R549 B.n445 B.n444 163.367
R550 B.n441 B.n440 163.367
R551 B.n437 B.n436 163.367
R552 B.n433 B.n432 163.367
R553 B.n429 B.n428 163.367
R554 B.n425 B.n424 163.367
R555 B.n421 B.n420 163.367
R556 B.n417 B.n416 163.367
R557 B.n413 B.n412 163.367
R558 B.n409 B.n408 163.367
R559 B.n405 B.n404 163.367
R560 B.n400 B.n399 163.367
R561 B.n396 B.n395 163.367
R562 B.n392 B.n391 163.367
R563 B.n388 B.n387 163.367
R564 B.n384 B.n383 163.367
R565 B.n380 B.n379 163.367
R566 B.n376 B.n375 163.367
R567 B.n372 B.n371 163.367
R568 B.n368 B.n367 163.367
R569 B.n364 B.n363 163.367
R570 B.n360 B.n359 163.367
R571 B.n356 B.n355 163.367
R572 B.n352 B.n351 163.367
R573 B.n348 B.n347 163.367
R574 B.n344 B.n343 163.367
R575 B.n340 B.n339 163.367
R576 B.n336 B.n335 163.367
R577 B.n332 B.n294 163.367
R578 B.n464 B.n292 163.367
R579 B.n464 B.n286 163.367
R580 B.n472 B.n286 163.367
R581 B.n472 B.n284 163.367
R582 B.n476 B.n284 163.367
R583 B.n476 B.n278 163.367
R584 B.n484 B.n278 163.367
R585 B.n484 B.n276 163.367
R586 B.n488 B.n276 163.367
R587 B.n488 B.n270 163.367
R588 B.n496 B.n270 163.367
R589 B.n496 B.n268 163.367
R590 B.n500 B.n268 163.367
R591 B.n500 B.n262 163.367
R592 B.n508 B.n262 163.367
R593 B.n508 B.n260 163.367
R594 B.n512 B.n260 163.367
R595 B.n512 B.n254 163.367
R596 B.n520 B.n254 163.367
R597 B.n520 B.n252 163.367
R598 B.n524 B.n252 163.367
R599 B.n524 B.n246 163.367
R600 B.n532 B.n246 163.367
R601 B.n532 B.n244 163.367
R602 B.n536 B.n244 163.367
R603 B.n536 B.n238 163.367
R604 B.n544 B.n238 163.367
R605 B.n544 B.n236 163.367
R606 B.n549 B.n236 163.367
R607 B.n549 B.n230 163.367
R608 B.n557 B.n230 163.367
R609 B.n558 B.n557 163.367
R610 B.n558 B.n5 163.367
R611 B.n6 B.n5 163.367
R612 B.n7 B.n6 163.367
R613 B.n563 B.n7 163.367
R614 B.n563 B.n12 163.367
R615 B.n13 B.n12 163.367
R616 B.n14 B.n13 163.367
R617 B.n568 B.n14 163.367
R618 B.n568 B.n19 163.367
R619 B.n20 B.n19 163.367
R620 B.n21 B.n20 163.367
R621 B.n573 B.n21 163.367
R622 B.n573 B.n26 163.367
R623 B.n27 B.n26 163.367
R624 B.n28 B.n27 163.367
R625 B.n578 B.n28 163.367
R626 B.n578 B.n33 163.367
R627 B.n34 B.n33 163.367
R628 B.n35 B.n34 163.367
R629 B.n583 B.n35 163.367
R630 B.n583 B.n40 163.367
R631 B.n41 B.n40 163.367
R632 B.n42 B.n41 163.367
R633 B.n588 B.n42 163.367
R634 B.n588 B.n47 163.367
R635 B.n48 B.n47 163.367
R636 B.n49 B.n48 163.367
R637 B.n593 B.n49 163.367
R638 B.n593 B.n54 163.367
R639 B.n55 B.n54 163.367
R640 B.n56 B.n55 163.367
R641 B.n598 B.n56 163.367
R642 B.n598 B.n61 163.367
R643 B.n62 B.n61 163.367
R644 B.n105 B.n104 163.367
R645 B.n109 B.n108 163.367
R646 B.n113 B.n112 163.367
R647 B.n117 B.n116 163.367
R648 B.n121 B.n120 163.367
R649 B.n125 B.n124 163.367
R650 B.n129 B.n128 163.367
R651 B.n133 B.n132 163.367
R652 B.n137 B.n136 163.367
R653 B.n141 B.n140 163.367
R654 B.n145 B.n144 163.367
R655 B.n149 B.n148 163.367
R656 B.n153 B.n152 163.367
R657 B.n157 B.n156 163.367
R658 B.n161 B.n160 163.367
R659 B.n165 B.n164 163.367
R660 B.n169 B.n168 163.367
R661 B.n173 B.n172 163.367
R662 B.n178 B.n177 163.367
R663 B.n182 B.n181 163.367
R664 B.n186 B.n185 163.367
R665 B.n190 B.n189 163.367
R666 B.n194 B.n193 163.367
R667 B.n198 B.n197 163.367
R668 B.n202 B.n201 163.367
R669 B.n206 B.n205 163.367
R670 B.n210 B.n209 163.367
R671 B.n214 B.n213 163.367
R672 B.n218 B.n217 163.367
R673 B.n222 B.n221 163.367
R674 B.n226 B.n225 163.367
R675 B.n603 B.n95 163.367
R676 B.n458 B.n291 115.234
R677 B.n605 B.n604 115.234
R678 B.n330 B.n329 82.4247
R679 B.n328 B.n327 82.4247
R680 B.n99 B.n98 82.4247
R681 B.n97 B.n96 82.4247
R682 B.n457 B.n456 71.676
R683 B.n451 B.n295 71.676
R684 B.n448 B.n296 71.676
R685 B.n444 B.n297 71.676
R686 B.n440 B.n298 71.676
R687 B.n436 B.n299 71.676
R688 B.n432 B.n300 71.676
R689 B.n428 B.n301 71.676
R690 B.n424 B.n302 71.676
R691 B.n420 B.n303 71.676
R692 B.n416 B.n304 71.676
R693 B.n412 B.n305 71.676
R694 B.n408 B.n306 71.676
R695 B.n404 B.n307 71.676
R696 B.n399 B.n308 71.676
R697 B.n395 B.n309 71.676
R698 B.n391 B.n310 71.676
R699 B.n387 B.n311 71.676
R700 B.n383 B.n312 71.676
R701 B.n379 B.n313 71.676
R702 B.n375 B.n314 71.676
R703 B.n371 B.n315 71.676
R704 B.n367 B.n316 71.676
R705 B.n363 B.n317 71.676
R706 B.n359 B.n318 71.676
R707 B.n355 B.n319 71.676
R708 B.n351 B.n320 71.676
R709 B.n347 B.n321 71.676
R710 B.n343 B.n322 71.676
R711 B.n339 B.n323 71.676
R712 B.n335 B.n324 71.676
R713 B.n459 B.n294 71.676
R714 B.n101 B.n63 71.676
R715 B.n105 B.n64 71.676
R716 B.n109 B.n65 71.676
R717 B.n113 B.n66 71.676
R718 B.n117 B.n67 71.676
R719 B.n121 B.n68 71.676
R720 B.n125 B.n69 71.676
R721 B.n129 B.n70 71.676
R722 B.n133 B.n71 71.676
R723 B.n137 B.n72 71.676
R724 B.n141 B.n73 71.676
R725 B.n145 B.n74 71.676
R726 B.n149 B.n75 71.676
R727 B.n153 B.n76 71.676
R728 B.n157 B.n77 71.676
R729 B.n161 B.n78 71.676
R730 B.n165 B.n79 71.676
R731 B.n169 B.n80 71.676
R732 B.n173 B.n81 71.676
R733 B.n178 B.n82 71.676
R734 B.n182 B.n83 71.676
R735 B.n186 B.n84 71.676
R736 B.n190 B.n85 71.676
R737 B.n194 B.n86 71.676
R738 B.n198 B.n87 71.676
R739 B.n202 B.n88 71.676
R740 B.n206 B.n89 71.676
R741 B.n210 B.n90 71.676
R742 B.n214 B.n91 71.676
R743 B.n218 B.n92 71.676
R744 B.n222 B.n93 71.676
R745 B.n226 B.n94 71.676
R746 B.n95 B.n94 71.676
R747 B.n225 B.n93 71.676
R748 B.n221 B.n92 71.676
R749 B.n217 B.n91 71.676
R750 B.n213 B.n90 71.676
R751 B.n209 B.n89 71.676
R752 B.n205 B.n88 71.676
R753 B.n201 B.n87 71.676
R754 B.n197 B.n86 71.676
R755 B.n193 B.n85 71.676
R756 B.n189 B.n84 71.676
R757 B.n185 B.n83 71.676
R758 B.n181 B.n82 71.676
R759 B.n177 B.n81 71.676
R760 B.n172 B.n80 71.676
R761 B.n168 B.n79 71.676
R762 B.n164 B.n78 71.676
R763 B.n160 B.n77 71.676
R764 B.n156 B.n76 71.676
R765 B.n152 B.n75 71.676
R766 B.n148 B.n74 71.676
R767 B.n144 B.n73 71.676
R768 B.n140 B.n72 71.676
R769 B.n136 B.n71 71.676
R770 B.n132 B.n70 71.676
R771 B.n128 B.n69 71.676
R772 B.n124 B.n68 71.676
R773 B.n120 B.n67 71.676
R774 B.n116 B.n66 71.676
R775 B.n112 B.n65 71.676
R776 B.n108 B.n64 71.676
R777 B.n104 B.n63 71.676
R778 B.n457 B.n326 71.676
R779 B.n449 B.n295 71.676
R780 B.n445 B.n296 71.676
R781 B.n441 B.n297 71.676
R782 B.n437 B.n298 71.676
R783 B.n433 B.n299 71.676
R784 B.n429 B.n300 71.676
R785 B.n425 B.n301 71.676
R786 B.n421 B.n302 71.676
R787 B.n417 B.n303 71.676
R788 B.n413 B.n304 71.676
R789 B.n409 B.n305 71.676
R790 B.n405 B.n306 71.676
R791 B.n400 B.n307 71.676
R792 B.n396 B.n308 71.676
R793 B.n392 B.n309 71.676
R794 B.n388 B.n310 71.676
R795 B.n384 B.n311 71.676
R796 B.n380 B.n312 71.676
R797 B.n376 B.n313 71.676
R798 B.n372 B.n314 71.676
R799 B.n368 B.n315 71.676
R800 B.n364 B.n316 71.676
R801 B.n360 B.n317 71.676
R802 B.n356 B.n318 71.676
R803 B.n352 B.n319 71.676
R804 B.n348 B.n320 71.676
R805 B.n344 B.n321 71.676
R806 B.n340 B.n322 71.676
R807 B.n336 B.n323 71.676
R808 B.n332 B.n324 71.676
R809 B.n460 B.n459 71.676
R810 B.n465 B.n291 59.8166
R811 B.n465 B.n287 59.8166
R812 B.n471 B.n287 59.8166
R813 B.n471 B.n283 59.8166
R814 B.n477 B.n283 59.8166
R815 B.n477 B.n279 59.8166
R816 B.n483 B.n279 59.8166
R817 B.n483 B.n275 59.8166
R818 B.n489 B.n275 59.8166
R819 B.n495 B.n271 59.8166
R820 B.n495 B.n267 59.8166
R821 B.n501 B.n267 59.8166
R822 B.n501 B.n263 59.8166
R823 B.n507 B.n263 59.8166
R824 B.n507 B.n259 59.8166
R825 B.n513 B.n259 59.8166
R826 B.n513 B.n255 59.8166
R827 B.n519 B.n255 59.8166
R828 B.n519 B.n251 59.8166
R829 B.n525 B.n251 59.8166
R830 B.n525 B.n247 59.8166
R831 B.n531 B.n247 59.8166
R832 B.n531 B.n243 59.8166
R833 B.n537 B.n243 59.8166
R834 B.n543 B.n239 59.8166
R835 B.n543 B.n235 59.8166
R836 B.n550 B.n235 59.8166
R837 B.n550 B.n231 59.8166
R838 B.n556 B.n231 59.8166
R839 B.n556 B.n4 59.8166
R840 B.n670 B.n4 59.8166
R841 B.n670 B.n669 59.8166
R842 B.n669 B.n668 59.8166
R843 B.n668 B.n8 59.8166
R844 B.n662 B.n8 59.8166
R845 B.n662 B.n661 59.8166
R846 B.n661 B.n660 59.8166
R847 B.n660 B.n15 59.8166
R848 B.n654 B.n653 59.8166
R849 B.n653 B.n652 59.8166
R850 B.n652 B.n22 59.8166
R851 B.n646 B.n22 59.8166
R852 B.n646 B.n645 59.8166
R853 B.n645 B.n644 59.8166
R854 B.n644 B.n29 59.8166
R855 B.n638 B.n29 59.8166
R856 B.n638 B.n637 59.8166
R857 B.n637 B.n636 59.8166
R858 B.n636 B.n36 59.8166
R859 B.n630 B.n36 59.8166
R860 B.n630 B.n629 59.8166
R861 B.n629 B.n628 59.8166
R862 B.n628 B.n43 59.8166
R863 B.n622 B.n621 59.8166
R864 B.n621 B.n620 59.8166
R865 B.n620 B.n50 59.8166
R866 B.n614 B.n50 59.8166
R867 B.n614 B.n613 59.8166
R868 B.n613 B.n612 59.8166
R869 B.n612 B.n57 59.8166
R870 B.n606 B.n57 59.8166
R871 B.n606 B.n605 59.8166
R872 B.n331 B.n330 59.5399
R873 B.n402 B.n328 59.5399
R874 B.n100 B.n99 59.5399
R875 B.n175 B.n97 59.5399
R876 B.t0 B.n239 51.0201
R877 B.t1 B.n15 51.0201
R878 B.t3 B.n271 33.4271
R879 B.t10 B.n43 33.4271
R880 B.n102 B.n59 32.3127
R881 B.n602 B.n601 32.3127
R882 B.n462 B.n461 32.3127
R883 B.n455 B.n289 32.3127
R884 B.n489 B.t3 26.3899
R885 B.n622 B.t10 26.3899
R886 B B.n672 18.0485
R887 B.n103 B.n102 10.6151
R888 B.n106 B.n103 10.6151
R889 B.n107 B.n106 10.6151
R890 B.n110 B.n107 10.6151
R891 B.n111 B.n110 10.6151
R892 B.n114 B.n111 10.6151
R893 B.n115 B.n114 10.6151
R894 B.n118 B.n115 10.6151
R895 B.n119 B.n118 10.6151
R896 B.n122 B.n119 10.6151
R897 B.n123 B.n122 10.6151
R898 B.n126 B.n123 10.6151
R899 B.n127 B.n126 10.6151
R900 B.n130 B.n127 10.6151
R901 B.n131 B.n130 10.6151
R902 B.n134 B.n131 10.6151
R903 B.n135 B.n134 10.6151
R904 B.n138 B.n135 10.6151
R905 B.n139 B.n138 10.6151
R906 B.n142 B.n139 10.6151
R907 B.n143 B.n142 10.6151
R908 B.n146 B.n143 10.6151
R909 B.n147 B.n146 10.6151
R910 B.n150 B.n147 10.6151
R911 B.n151 B.n150 10.6151
R912 B.n154 B.n151 10.6151
R913 B.n155 B.n154 10.6151
R914 B.n159 B.n158 10.6151
R915 B.n162 B.n159 10.6151
R916 B.n163 B.n162 10.6151
R917 B.n166 B.n163 10.6151
R918 B.n167 B.n166 10.6151
R919 B.n170 B.n167 10.6151
R920 B.n171 B.n170 10.6151
R921 B.n174 B.n171 10.6151
R922 B.n179 B.n176 10.6151
R923 B.n180 B.n179 10.6151
R924 B.n183 B.n180 10.6151
R925 B.n184 B.n183 10.6151
R926 B.n187 B.n184 10.6151
R927 B.n188 B.n187 10.6151
R928 B.n191 B.n188 10.6151
R929 B.n192 B.n191 10.6151
R930 B.n195 B.n192 10.6151
R931 B.n196 B.n195 10.6151
R932 B.n199 B.n196 10.6151
R933 B.n200 B.n199 10.6151
R934 B.n203 B.n200 10.6151
R935 B.n204 B.n203 10.6151
R936 B.n207 B.n204 10.6151
R937 B.n208 B.n207 10.6151
R938 B.n211 B.n208 10.6151
R939 B.n212 B.n211 10.6151
R940 B.n215 B.n212 10.6151
R941 B.n216 B.n215 10.6151
R942 B.n219 B.n216 10.6151
R943 B.n220 B.n219 10.6151
R944 B.n223 B.n220 10.6151
R945 B.n224 B.n223 10.6151
R946 B.n227 B.n224 10.6151
R947 B.n228 B.n227 10.6151
R948 B.n602 B.n228 10.6151
R949 B.n463 B.n462 10.6151
R950 B.n463 B.n285 10.6151
R951 B.n473 B.n285 10.6151
R952 B.n474 B.n473 10.6151
R953 B.n475 B.n474 10.6151
R954 B.n475 B.n277 10.6151
R955 B.n485 B.n277 10.6151
R956 B.n486 B.n485 10.6151
R957 B.n487 B.n486 10.6151
R958 B.n487 B.n269 10.6151
R959 B.n497 B.n269 10.6151
R960 B.n498 B.n497 10.6151
R961 B.n499 B.n498 10.6151
R962 B.n499 B.n261 10.6151
R963 B.n509 B.n261 10.6151
R964 B.n510 B.n509 10.6151
R965 B.n511 B.n510 10.6151
R966 B.n511 B.n253 10.6151
R967 B.n521 B.n253 10.6151
R968 B.n522 B.n521 10.6151
R969 B.n523 B.n522 10.6151
R970 B.n523 B.n245 10.6151
R971 B.n533 B.n245 10.6151
R972 B.n534 B.n533 10.6151
R973 B.n535 B.n534 10.6151
R974 B.n535 B.n237 10.6151
R975 B.n545 B.n237 10.6151
R976 B.n546 B.n545 10.6151
R977 B.n548 B.n546 10.6151
R978 B.n548 B.n547 10.6151
R979 B.n547 B.n229 10.6151
R980 B.n559 B.n229 10.6151
R981 B.n560 B.n559 10.6151
R982 B.n561 B.n560 10.6151
R983 B.n562 B.n561 10.6151
R984 B.n564 B.n562 10.6151
R985 B.n565 B.n564 10.6151
R986 B.n566 B.n565 10.6151
R987 B.n567 B.n566 10.6151
R988 B.n569 B.n567 10.6151
R989 B.n570 B.n569 10.6151
R990 B.n571 B.n570 10.6151
R991 B.n572 B.n571 10.6151
R992 B.n574 B.n572 10.6151
R993 B.n575 B.n574 10.6151
R994 B.n576 B.n575 10.6151
R995 B.n577 B.n576 10.6151
R996 B.n579 B.n577 10.6151
R997 B.n580 B.n579 10.6151
R998 B.n581 B.n580 10.6151
R999 B.n582 B.n581 10.6151
R1000 B.n584 B.n582 10.6151
R1001 B.n585 B.n584 10.6151
R1002 B.n586 B.n585 10.6151
R1003 B.n587 B.n586 10.6151
R1004 B.n589 B.n587 10.6151
R1005 B.n590 B.n589 10.6151
R1006 B.n591 B.n590 10.6151
R1007 B.n592 B.n591 10.6151
R1008 B.n594 B.n592 10.6151
R1009 B.n595 B.n594 10.6151
R1010 B.n596 B.n595 10.6151
R1011 B.n597 B.n596 10.6151
R1012 B.n599 B.n597 10.6151
R1013 B.n600 B.n599 10.6151
R1014 B.n601 B.n600 10.6151
R1015 B.n455 B.n454 10.6151
R1016 B.n454 B.n453 10.6151
R1017 B.n453 B.n452 10.6151
R1018 B.n452 B.n450 10.6151
R1019 B.n450 B.n447 10.6151
R1020 B.n447 B.n446 10.6151
R1021 B.n446 B.n443 10.6151
R1022 B.n443 B.n442 10.6151
R1023 B.n442 B.n439 10.6151
R1024 B.n439 B.n438 10.6151
R1025 B.n438 B.n435 10.6151
R1026 B.n435 B.n434 10.6151
R1027 B.n434 B.n431 10.6151
R1028 B.n431 B.n430 10.6151
R1029 B.n430 B.n427 10.6151
R1030 B.n427 B.n426 10.6151
R1031 B.n426 B.n423 10.6151
R1032 B.n423 B.n422 10.6151
R1033 B.n422 B.n419 10.6151
R1034 B.n419 B.n418 10.6151
R1035 B.n418 B.n415 10.6151
R1036 B.n415 B.n414 10.6151
R1037 B.n414 B.n411 10.6151
R1038 B.n411 B.n410 10.6151
R1039 B.n410 B.n407 10.6151
R1040 B.n407 B.n406 10.6151
R1041 B.n406 B.n403 10.6151
R1042 B.n401 B.n398 10.6151
R1043 B.n398 B.n397 10.6151
R1044 B.n397 B.n394 10.6151
R1045 B.n394 B.n393 10.6151
R1046 B.n393 B.n390 10.6151
R1047 B.n390 B.n389 10.6151
R1048 B.n389 B.n386 10.6151
R1049 B.n386 B.n385 10.6151
R1050 B.n382 B.n381 10.6151
R1051 B.n381 B.n378 10.6151
R1052 B.n378 B.n377 10.6151
R1053 B.n377 B.n374 10.6151
R1054 B.n374 B.n373 10.6151
R1055 B.n373 B.n370 10.6151
R1056 B.n370 B.n369 10.6151
R1057 B.n369 B.n366 10.6151
R1058 B.n366 B.n365 10.6151
R1059 B.n365 B.n362 10.6151
R1060 B.n362 B.n361 10.6151
R1061 B.n361 B.n358 10.6151
R1062 B.n358 B.n357 10.6151
R1063 B.n357 B.n354 10.6151
R1064 B.n354 B.n353 10.6151
R1065 B.n353 B.n350 10.6151
R1066 B.n350 B.n349 10.6151
R1067 B.n349 B.n346 10.6151
R1068 B.n346 B.n345 10.6151
R1069 B.n345 B.n342 10.6151
R1070 B.n342 B.n341 10.6151
R1071 B.n341 B.n338 10.6151
R1072 B.n338 B.n337 10.6151
R1073 B.n337 B.n334 10.6151
R1074 B.n334 B.n333 10.6151
R1075 B.n333 B.n293 10.6151
R1076 B.n461 B.n293 10.6151
R1077 B.n467 B.n289 10.6151
R1078 B.n468 B.n467 10.6151
R1079 B.n469 B.n468 10.6151
R1080 B.n469 B.n281 10.6151
R1081 B.n479 B.n281 10.6151
R1082 B.n480 B.n479 10.6151
R1083 B.n481 B.n480 10.6151
R1084 B.n481 B.n273 10.6151
R1085 B.n491 B.n273 10.6151
R1086 B.n492 B.n491 10.6151
R1087 B.n493 B.n492 10.6151
R1088 B.n493 B.n265 10.6151
R1089 B.n503 B.n265 10.6151
R1090 B.n504 B.n503 10.6151
R1091 B.n505 B.n504 10.6151
R1092 B.n505 B.n257 10.6151
R1093 B.n515 B.n257 10.6151
R1094 B.n516 B.n515 10.6151
R1095 B.n517 B.n516 10.6151
R1096 B.n517 B.n249 10.6151
R1097 B.n527 B.n249 10.6151
R1098 B.n528 B.n527 10.6151
R1099 B.n529 B.n528 10.6151
R1100 B.n529 B.n241 10.6151
R1101 B.n539 B.n241 10.6151
R1102 B.n540 B.n539 10.6151
R1103 B.n541 B.n540 10.6151
R1104 B.n541 B.n233 10.6151
R1105 B.n552 B.n233 10.6151
R1106 B.n553 B.n552 10.6151
R1107 B.n554 B.n553 10.6151
R1108 B.n554 B.n0 10.6151
R1109 B.n666 B.n1 10.6151
R1110 B.n666 B.n665 10.6151
R1111 B.n665 B.n664 10.6151
R1112 B.n664 B.n10 10.6151
R1113 B.n658 B.n10 10.6151
R1114 B.n658 B.n657 10.6151
R1115 B.n657 B.n656 10.6151
R1116 B.n656 B.n17 10.6151
R1117 B.n650 B.n17 10.6151
R1118 B.n650 B.n649 10.6151
R1119 B.n649 B.n648 10.6151
R1120 B.n648 B.n24 10.6151
R1121 B.n642 B.n24 10.6151
R1122 B.n642 B.n641 10.6151
R1123 B.n641 B.n640 10.6151
R1124 B.n640 B.n31 10.6151
R1125 B.n634 B.n31 10.6151
R1126 B.n634 B.n633 10.6151
R1127 B.n633 B.n632 10.6151
R1128 B.n632 B.n38 10.6151
R1129 B.n626 B.n38 10.6151
R1130 B.n626 B.n625 10.6151
R1131 B.n625 B.n624 10.6151
R1132 B.n624 B.n45 10.6151
R1133 B.n618 B.n45 10.6151
R1134 B.n618 B.n617 10.6151
R1135 B.n617 B.n616 10.6151
R1136 B.n616 B.n52 10.6151
R1137 B.n610 B.n52 10.6151
R1138 B.n610 B.n609 10.6151
R1139 B.n609 B.n608 10.6151
R1140 B.n608 B.n59 10.6151
R1141 B.n537 B.t0 8.79698
R1142 B.n654 B.t1 8.79698
R1143 B.n158 B.n100 6.5566
R1144 B.n175 B.n174 6.5566
R1145 B.n402 B.n401 6.5566
R1146 B.n385 B.n331 6.5566
R1147 B.n155 B.n100 4.05904
R1148 B.n176 B.n175 4.05904
R1149 B.n403 B.n402 4.05904
R1150 B.n382 B.n331 4.05904
R1151 B.n672 B.n0 2.81026
R1152 B.n672 B.n1 2.81026
R1153 VP.n0 VP.t0 124.031
R1154 VP.n0 VP.t1 79.4874
R1155 VP VP.n0 0.621237
R1156 VTAIL.n138 VTAIL.n108 214.453
R1157 VTAIL.n30 VTAIL.n0 214.453
R1158 VTAIL.n102 VTAIL.n72 214.453
R1159 VTAIL.n66 VTAIL.n36 214.453
R1160 VTAIL.n121 VTAIL.n120 185
R1161 VTAIL.n123 VTAIL.n122 185
R1162 VTAIL.n116 VTAIL.n115 185
R1163 VTAIL.n129 VTAIL.n128 185
R1164 VTAIL.n131 VTAIL.n130 185
R1165 VTAIL.n112 VTAIL.n111 185
R1166 VTAIL.n137 VTAIL.n136 185
R1167 VTAIL.n139 VTAIL.n138 185
R1168 VTAIL.n13 VTAIL.n12 185
R1169 VTAIL.n15 VTAIL.n14 185
R1170 VTAIL.n8 VTAIL.n7 185
R1171 VTAIL.n21 VTAIL.n20 185
R1172 VTAIL.n23 VTAIL.n22 185
R1173 VTAIL.n4 VTAIL.n3 185
R1174 VTAIL.n29 VTAIL.n28 185
R1175 VTAIL.n31 VTAIL.n30 185
R1176 VTAIL.n103 VTAIL.n102 185
R1177 VTAIL.n101 VTAIL.n100 185
R1178 VTAIL.n76 VTAIL.n75 185
R1179 VTAIL.n95 VTAIL.n94 185
R1180 VTAIL.n93 VTAIL.n92 185
R1181 VTAIL.n80 VTAIL.n79 185
R1182 VTAIL.n87 VTAIL.n86 185
R1183 VTAIL.n85 VTAIL.n84 185
R1184 VTAIL.n67 VTAIL.n66 185
R1185 VTAIL.n65 VTAIL.n64 185
R1186 VTAIL.n40 VTAIL.n39 185
R1187 VTAIL.n59 VTAIL.n58 185
R1188 VTAIL.n57 VTAIL.n56 185
R1189 VTAIL.n44 VTAIL.n43 185
R1190 VTAIL.n51 VTAIL.n50 185
R1191 VTAIL.n49 VTAIL.n48 185
R1192 VTAIL.n119 VTAIL.t1 149.524
R1193 VTAIL.n11 VTAIL.t3 149.524
R1194 VTAIL.n83 VTAIL.t2 149.524
R1195 VTAIL.n47 VTAIL.t0 149.524
R1196 VTAIL.n122 VTAIL.n121 104.615
R1197 VTAIL.n122 VTAIL.n115 104.615
R1198 VTAIL.n129 VTAIL.n115 104.615
R1199 VTAIL.n130 VTAIL.n129 104.615
R1200 VTAIL.n130 VTAIL.n111 104.615
R1201 VTAIL.n137 VTAIL.n111 104.615
R1202 VTAIL.n138 VTAIL.n137 104.615
R1203 VTAIL.n14 VTAIL.n13 104.615
R1204 VTAIL.n14 VTAIL.n7 104.615
R1205 VTAIL.n21 VTAIL.n7 104.615
R1206 VTAIL.n22 VTAIL.n21 104.615
R1207 VTAIL.n22 VTAIL.n3 104.615
R1208 VTAIL.n29 VTAIL.n3 104.615
R1209 VTAIL.n30 VTAIL.n29 104.615
R1210 VTAIL.n102 VTAIL.n101 104.615
R1211 VTAIL.n101 VTAIL.n75 104.615
R1212 VTAIL.n94 VTAIL.n75 104.615
R1213 VTAIL.n94 VTAIL.n93 104.615
R1214 VTAIL.n93 VTAIL.n79 104.615
R1215 VTAIL.n86 VTAIL.n79 104.615
R1216 VTAIL.n86 VTAIL.n85 104.615
R1217 VTAIL.n66 VTAIL.n65 104.615
R1218 VTAIL.n65 VTAIL.n39 104.615
R1219 VTAIL.n58 VTAIL.n39 104.615
R1220 VTAIL.n58 VTAIL.n57 104.615
R1221 VTAIL.n57 VTAIL.n43 104.615
R1222 VTAIL.n50 VTAIL.n43 104.615
R1223 VTAIL.n50 VTAIL.n49 104.615
R1224 VTAIL.n121 VTAIL.t1 52.3082
R1225 VTAIL.n13 VTAIL.t3 52.3082
R1226 VTAIL.n85 VTAIL.t2 52.3082
R1227 VTAIL.n49 VTAIL.t0 52.3082
R1228 VTAIL.n143 VTAIL.n142 35.0944
R1229 VTAIL.n35 VTAIL.n34 35.0944
R1230 VTAIL.n107 VTAIL.n106 35.0944
R1231 VTAIL.n71 VTAIL.n70 35.0944
R1232 VTAIL.n71 VTAIL.n35 25.9272
R1233 VTAIL.n143 VTAIL.n107 22.2634
R1234 VTAIL.n140 VTAIL.n139 12.8005
R1235 VTAIL.n32 VTAIL.n31 12.8005
R1236 VTAIL.n104 VTAIL.n103 12.8005
R1237 VTAIL.n68 VTAIL.n67 12.8005
R1238 VTAIL.n136 VTAIL.n110 12.0247
R1239 VTAIL.n28 VTAIL.n2 12.0247
R1240 VTAIL.n100 VTAIL.n74 12.0247
R1241 VTAIL.n64 VTAIL.n38 12.0247
R1242 VTAIL.n135 VTAIL.n112 11.249
R1243 VTAIL.n27 VTAIL.n4 11.249
R1244 VTAIL.n99 VTAIL.n76 11.249
R1245 VTAIL.n63 VTAIL.n40 11.249
R1246 VTAIL.n132 VTAIL.n131 10.4732
R1247 VTAIL.n24 VTAIL.n23 10.4732
R1248 VTAIL.n96 VTAIL.n95 10.4732
R1249 VTAIL.n60 VTAIL.n59 10.4732
R1250 VTAIL.n120 VTAIL.n119 10.2747
R1251 VTAIL.n12 VTAIL.n11 10.2747
R1252 VTAIL.n84 VTAIL.n83 10.2747
R1253 VTAIL.n48 VTAIL.n47 10.2747
R1254 VTAIL.n128 VTAIL.n114 9.69747
R1255 VTAIL.n20 VTAIL.n6 9.69747
R1256 VTAIL.n92 VTAIL.n78 9.69747
R1257 VTAIL.n56 VTAIL.n42 9.69747
R1258 VTAIL.n142 VTAIL.n141 9.45567
R1259 VTAIL.n34 VTAIL.n33 9.45567
R1260 VTAIL.n106 VTAIL.n105 9.45567
R1261 VTAIL.n70 VTAIL.n69 9.45567
R1262 VTAIL.n118 VTAIL.n117 9.3005
R1263 VTAIL.n125 VTAIL.n124 9.3005
R1264 VTAIL.n127 VTAIL.n126 9.3005
R1265 VTAIL.n114 VTAIL.n113 9.3005
R1266 VTAIL.n133 VTAIL.n132 9.3005
R1267 VTAIL.n135 VTAIL.n134 9.3005
R1268 VTAIL.n110 VTAIL.n109 9.3005
R1269 VTAIL.n141 VTAIL.n140 9.3005
R1270 VTAIL.n10 VTAIL.n9 9.3005
R1271 VTAIL.n17 VTAIL.n16 9.3005
R1272 VTAIL.n19 VTAIL.n18 9.3005
R1273 VTAIL.n6 VTAIL.n5 9.3005
R1274 VTAIL.n25 VTAIL.n24 9.3005
R1275 VTAIL.n27 VTAIL.n26 9.3005
R1276 VTAIL.n2 VTAIL.n1 9.3005
R1277 VTAIL.n33 VTAIL.n32 9.3005
R1278 VTAIL.n82 VTAIL.n81 9.3005
R1279 VTAIL.n89 VTAIL.n88 9.3005
R1280 VTAIL.n91 VTAIL.n90 9.3005
R1281 VTAIL.n78 VTAIL.n77 9.3005
R1282 VTAIL.n97 VTAIL.n96 9.3005
R1283 VTAIL.n99 VTAIL.n98 9.3005
R1284 VTAIL.n74 VTAIL.n73 9.3005
R1285 VTAIL.n105 VTAIL.n104 9.3005
R1286 VTAIL.n46 VTAIL.n45 9.3005
R1287 VTAIL.n53 VTAIL.n52 9.3005
R1288 VTAIL.n55 VTAIL.n54 9.3005
R1289 VTAIL.n42 VTAIL.n41 9.3005
R1290 VTAIL.n61 VTAIL.n60 9.3005
R1291 VTAIL.n63 VTAIL.n62 9.3005
R1292 VTAIL.n38 VTAIL.n37 9.3005
R1293 VTAIL.n69 VTAIL.n68 9.3005
R1294 VTAIL.n127 VTAIL.n116 8.92171
R1295 VTAIL.n19 VTAIL.n8 8.92171
R1296 VTAIL.n91 VTAIL.n80 8.92171
R1297 VTAIL.n55 VTAIL.n44 8.92171
R1298 VTAIL.n142 VTAIL.n108 8.2187
R1299 VTAIL.n34 VTAIL.n0 8.2187
R1300 VTAIL.n106 VTAIL.n72 8.2187
R1301 VTAIL.n70 VTAIL.n36 8.2187
R1302 VTAIL.n124 VTAIL.n123 8.14595
R1303 VTAIL.n16 VTAIL.n15 8.14595
R1304 VTAIL.n88 VTAIL.n87 8.14595
R1305 VTAIL.n52 VTAIL.n51 8.14595
R1306 VTAIL.n120 VTAIL.n118 7.3702
R1307 VTAIL.n12 VTAIL.n10 7.3702
R1308 VTAIL.n84 VTAIL.n82 7.3702
R1309 VTAIL.n48 VTAIL.n46 7.3702
R1310 VTAIL.n123 VTAIL.n118 5.81868
R1311 VTAIL.n15 VTAIL.n10 5.81868
R1312 VTAIL.n87 VTAIL.n82 5.81868
R1313 VTAIL.n51 VTAIL.n46 5.81868
R1314 VTAIL.n140 VTAIL.n108 5.3904
R1315 VTAIL.n32 VTAIL.n0 5.3904
R1316 VTAIL.n104 VTAIL.n72 5.3904
R1317 VTAIL.n68 VTAIL.n36 5.3904
R1318 VTAIL.n124 VTAIL.n116 5.04292
R1319 VTAIL.n16 VTAIL.n8 5.04292
R1320 VTAIL.n88 VTAIL.n80 5.04292
R1321 VTAIL.n52 VTAIL.n44 5.04292
R1322 VTAIL.n128 VTAIL.n127 4.26717
R1323 VTAIL.n20 VTAIL.n19 4.26717
R1324 VTAIL.n92 VTAIL.n91 4.26717
R1325 VTAIL.n56 VTAIL.n55 4.26717
R1326 VTAIL.n131 VTAIL.n114 3.49141
R1327 VTAIL.n23 VTAIL.n6 3.49141
R1328 VTAIL.n95 VTAIL.n78 3.49141
R1329 VTAIL.n59 VTAIL.n42 3.49141
R1330 VTAIL.n119 VTAIL.n117 2.84305
R1331 VTAIL.n11 VTAIL.n9 2.84305
R1332 VTAIL.n83 VTAIL.n81 2.84305
R1333 VTAIL.n47 VTAIL.n45 2.84305
R1334 VTAIL.n132 VTAIL.n112 2.71565
R1335 VTAIL.n24 VTAIL.n4 2.71565
R1336 VTAIL.n96 VTAIL.n76 2.71565
R1337 VTAIL.n60 VTAIL.n40 2.71565
R1338 VTAIL.n107 VTAIL.n71 2.30222
R1339 VTAIL.n136 VTAIL.n135 1.93989
R1340 VTAIL.n28 VTAIL.n27 1.93989
R1341 VTAIL.n100 VTAIL.n99 1.93989
R1342 VTAIL.n64 VTAIL.n63 1.93989
R1343 VTAIL VTAIL.n35 1.44447
R1344 VTAIL.n139 VTAIL.n110 1.16414
R1345 VTAIL.n31 VTAIL.n2 1.16414
R1346 VTAIL.n103 VTAIL.n74 1.16414
R1347 VTAIL.n67 VTAIL.n38 1.16414
R1348 VTAIL VTAIL.n143 0.858259
R1349 VTAIL.n125 VTAIL.n117 0.155672
R1350 VTAIL.n126 VTAIL.n125 0.155672
R1351 VTAIL.n126 VTAIL.n113 0.155672
R1352 VTAIL.n133 VTAIL.n113 0.155672
R1353 VTAIL.n134 VTAIL.n133 0.155672
R1354 VTAIL.n134 VTAIL.n109 0.155672
R1355 VTAIL.n141 VTAIL.n109 0.155672
R1356 VTAIL.n17 VTAIL.n9 0.155672
R1357 VTAIL.n18 VTAIL.n17 0.155672
R1358 VTAIL.n18 VTAIL.n5 0.155672
R1359 VTAIL.n25 VTAIL.n5 0.155672
R1360 VTAIL.n26 VTAIL.n25 0.155672
R1361 VTAIL.n26 VTAIL.n1 0.155672
R1362 VTAIL.n33 VTAIL.n1 0.155672
R1363 VTAIL.n105 VTAIL.n73 0.155672
R1364 VTAIL.n98 VTAIL.n73 0.155672
R1365 VTAIL.n98 VTAIL.n97 0.155672
R1366 VTAIL.n97 VTAIL.n77 0.155672
R1367 VTAIL.n90 VTAIL.n77 0.155672
R1368 VTAIL.n90 VTAIL.n89 0.155672
R1369 VTAIL.n89 VTAIL.n81 0.155672
R1370 VTAIL.n69 VTAIL.n37 0.155672
R1371 VTAIL.n62 VTAIL.n37 0.155672
R1372 VTAIL.n62 VTAIL.n61 0.155672
R1373 VTAIL.n61 VTAIL.n41 0.155672
R1374 VTAIL.n54 VTAIL.n41 0.155672
R1375 VTAIL.n54 VTAIL.n53 0.155672
R1376 VTAIL.n53 VTAIL.n45 0.155672
R1377 VDD1.n30 VDD1.n0 214.453
R1378 VDD1.n65 VDD1.n35 214.453
R1379 VDD1.n31 VDD1.n30 185
R1380 VDD1.n29 VDD1.n28 185
R1381 VDD1.n4 VDD1.n3 185
R1382 VDD1.n23 VDD1.n22 185
R1383 VDD1.n21 VDD1.n20 185
R1384 VDD1.n8 VDD1.n7 185
R1385 VDD1.n15 VDD1.n14 185
R1386 VDD1.n13 VDD1.n12 185
R1387 VDD1.n48 VDD1.n47 185
R1388 VDD1.n50 VDD1.n49 185
R1389 VDD1.n43 VDD1.n42 185
R1390 VDD1.n56 VDD1.n55 185
R1391 VDD1.n58 VDD1.n57 185
R1392 VDD1.n39 VDD1.n38 185
R1393 VDD1.n64 VDD1.n63 185
R1394 VDD1.n66 VDD1.n65 185
R1395 VDD1.n46 VDD1.t0 149.524
R1396 VDD1.n11 VDD1.t1 149.524
R1397 VDD1.n30 VDD1.n29 104.615
R1398 VDD1.n29 VDD1.n3 104.615
R1399 VDD1.n22 VDD1.n3 104.615
R1400 VDD1.n22 VDD1.n21 104.615
R1401 VDD1.n21 VDD1.n7 104.615
R1402 VDD1.n14 VDD1.n7 104.615
R1403 VDD1.n14 VDD1.n13 104.615
R1404 VDD1.n49 VDD1.n48 104.615
R1405 VDD1.n49 VDD1.n42 104.615
R1406 VDD1.n56 VDD1.n42 104.615
R1407 VDD1.n57 VDD1.n56 104.615
R1408 VDD1.n57 VDD1.n38 104.615
R1409 VDD1.n64 VDD1.n38 104.615
R1410 VDD1.n65 VDD1.n64 104.615
R1411 VDD1 VDD1.n69 90.4338
R1412 VDD1 VDD1.n34 52.7474
R1413 VDD1.n13 VDD1.t1 52.3082
R1414 VDD1.n48 VDD1.t0 52.3082
R1415 VDD1.n32 VDD1.n31 12.8005
R1416 VDD1.n67 VDD1.n66 12.8005
R1417 VDD1.n28 VDD1.n2 12.0247
R1418 VDD1.n63 VDD1.n37 12.0247
R1419 VDD1.n27 VDD1.n4 11.249
R1420 VDD1.n62 VDD1.n39 11.249
R1421 VDD1.n24 VDD1.n23 10.4732
R1422 VDD1.n59 VDD1.n58 10.4732
R1423 VDD1.n12 VDD1.n11 10.2747
R1424 VDD1.n47 VDD1.n46 10.2747
R1425 VDD1.n20 VDD1.n6 9.69747
R1426 VDD1.n55 VDD1.n41 9.69747
R1427 VDD1.n34 VDD1.n33 9.45567
R1428 VDD1.n69 VDD1.n68 9.45567
R1429 VDD1.n10 VDD1.n9 9.3005
R1430 VDD1.n17 VDD1.n16 9.3005
R1431 VDD1.n19 VDD1.n18 9.3005
R1432 VDD1.n6 VDD1.n5 9.3005
R1433 VDD1.n25 VDD1.n24 9.3005
R1434 VDD1.n27 VDD1.n26 9.3005
R1435 VDD1.n2 VDD1.n1 9.3005
R1436 VDD1.n33 VDD1.n32 9.3005
R1437 VDD1.n45 VDD1.n44 9.3005
R1438 VDD1.n52 VDD1.n51 9.3005
R1439 VDD1.n54 VDD1.n53 9.3005
R1440 VDD1.n41 VDD1.n40 9.3005
R1441 VDD1.n60 VDD1.n59 9.3005
R1442 VDD1.n62 VDD1.n61 9.3005
R1443 VDD1.n37 VDD1.n36 9.3005
R1444 VDD1.n68 VDD1.n67 9.3005
R1445 VDD1.n19 VDD1.n8 8.92171
R1446 VDD1.n54 VDD1.n43 8.92171
R1447 VDD1.n34 VDD1.n0 8.2187
R1448 VDD1.n69 VDD1.n35 8.2187
R1449 VDD1.n16 VDD1.n15 8.14595
R1450 VDD1.n51 VDD1.n50 8.14595
R1451 VDD1.n12 VDD1.n10 7.3702
R1452 VDD1.n47 VDD1.n45 7.3702
R1453 VDD1.n15 VDD1.n10 5.81868
R1454 VDD1.n50 VDD1.n45 5.81868
R1455 VDD1.n32 VDD1.n0 5.3904
R1456 VDD1.n67 VDD1.n35 5.3904
R1457 VDD1.n16 VDD1.n8 5.04292
R1458 VDD1.n51 VDD1.n43 5.04292
R1459 VDD1.n20 VDD1.n19 4.26717
R1460 VDD1.n55 VDD1.n54 4.26717
R1461 VDD1.n23 VDD1.n6 3.49141
R1462 VDD1.n58 VDD1.n41 3.49141
R1463 VDD1.n11 VDD1.n9 2.84305
R1464 VDD1.n46 VDD1.n44 2.84305
R1465 VDD1.n24 VDD1.n4 2.71565
R1466 VDD1.n59 VDD1.n39 2.71565
R1467 VDD1.n28 VDD1.n27 1.93989
R1468 VDD1.n63 VDD1.n62 1.93989
R1469 VDD1.n31 VDD1.n2 1.16414
R1470 VDD1.n66 VDD1.n37 1.16414
R1471 VDD1.n33 VDD1.n1 0.155672
R1472 VDD1.n26 VDD1.n1 0.155672
R1473 VDD1.n26 VDD1.n25 0.155672
R1474 VDD1.n25 VDD1.n5 0.155672
R1475 VDD1.n18 VDD1.n5 0.155672
R1476 VDD1.n18 VDD1.n17 0.155672
R1477 VDD1.n17 VDD1.n9 0.155672
R1478 VDD1.n52 VDD1.n44 0.155672
R1479 VDD1.n53 VDD1.n52 0.155672
R1480 VDD1.n53 VDD1.n40 0.155672
R1481 VDD1.n60 VDD1.n40 0.155672
R1482 VDD1.n61 VDD1.n60 0.155672
R1483 VDD1.n61 VDD1.n36 0.155672
R1484 VDD1.n68 VDD1.n36 0.155672
R1485 VN VN.t1 123.843
R1486 VN VN.t0 80.1081
R1487 VDD2.n65 VDD2.n35 214.453
R1488 VDD2.n30 VDD2.n0 214.453
R1489 VDD2.n66 VDD2.n65 185
R1490 VDD2.n64 VDD2.n63 185
R1491 VDD2.n39 VDD2.n38 185
R1492 VDD2.n58 VDD2.n57 185
R1493 VDD2.n56 VDD2.n55 185
R1494 VDD2.n43 VDD2.n42 185
R1495 VDD2.n50 VDD2.n49 185
R1496 VDD2.n48 VDD2.n47 185
R1497 VDD2.n13 VDD2.n12 185
R1498 VDD2.n15 VDD2.n14 185
R1499 VDD2.n8 VDD2.n7 185
R1500 VDD2.n21 VDD2.n20 185
R1501 VDD2.n23 VDD2.n22 185
R1502 VDD2.n4 VDD2.n3 185
R1503 VDD2.n29 VDD2.n28 185
R1504 VDD2.n31 VDD2.n30 185
R1505 VDD2.n11 VDD2.t1 149.524
R1506 VDD2.n46 VDD2.t0 149.524
R1507 VDD2.n65 VDD2.n64 104.615
R1508 VDD2.n64 VDD2.n38 104.615
R1509 VDD2.n57 VDD2.n38 104.615
R1510 VDD2.n57 VDD2.n56 104.615
R1511 VDD2.n56 VDD2.n42 104.615
R1512 VDD2.n49 VDD2.n42 104.615
R1513 VDD2.n49 VDD2.n48 104.615
R1514 VDD2.n14 VDD2.n13 104.615
R1515 VDD2.n14 VDD2.n7 104.615
R1516 VDD2.n21 VDD2.n7 104.615
R1517 VDD2.n22 VDD2.n21 104.615
R1518 VDD2.n22 VDD2.n3 104.615
R1519 VDD2.n29 VDD2.n3 104.615
R1520 VDD2.n30 VDD2.n29 104.615
R1521 VDD2.n70 VDD2.n34 88.993
R1522 VDD2.n48 VDD2.t0 52.3082
R1523 VDD2.n13 VDD2.t1 52.3082
R1524 VDD2.n70 VDD2.n69 51.7732
R1525 VDD2.n67 VDD2.n66 12.8005
R1526 VDD2.n32 VDD2.n31 12.8005
R1527 VDD2.n63 VDD2.n37 12.0247
R1528 VDD2.n28 VDD2.n2 12.0247
R1529 VDD2.n62 VDD2.n39 11.249
R1530 VDD2.n27 VDD2.n4 11.249
R1531 VDD2.n59 VDD2.n58 10.4732
R1532 VDD2.n24 VDD2.n23 10.4732
R1533 VDD2.n47 VDD2.n46 10.2747
R1534 VDD2.n12 VDD2.n11 10.2747
R1535 VDD2.n55 VDD2.n41 9.69747
R1536 VDD2.n20 VDD2.n6 9.69747
R1537 VDD2.n69 VDD2.n68 9.45567
R1538 VDD2.n34 VDD2.n33 9.45567
R1539 VDD2.n45 VDD2.n44 9.3005
R1540 VDD2.n52 VDD2.n51 9.3005
R1541 VDD2.n54 VDD2.n53 9.3005
R1542 VDD2.n41 VDD2.n40 9.3005
R1543 VDD2.n60 VDD2.n59 9.3005
R1544 VDD2.n62 VDD2.n61 9.3005
R1545 VDD2.n37 VDD2.n36 9.3005
R1546 VDD2.n68 VDD2.n67 9.3005
R1547 VDD2.n10 VDD2.n9 9.3005
R1548 VDD2.n17 VDD2.n16 9.3005
R1549 VDD2.n19 VDD2.n18 9.3005
R1550 VDD2.n6 VDD2.n5 9.3005
R1551 VDD2.n25 VDD2.n24 9.3005
R1552 VDD2.n27 VDD2.n26 9.3005
R1553 VDD2.n2 VDD2.n1 9.3005
R1554 VDD2.n33 VDD2.n32 9.3005
R1555 VDD2.n54 VDD2.n43 8.92171
R1556 VDD2.n19 VDD2.n8 8.92171
R1557 VDD2.n69 VDD2.n35 8.2187
R1558 VDD2.n34 VDD2.n0 8.2187
R1559 VDD2.n51 VDD2.n50 8.14595
R1560 VDD2.n16 VDD2.n15 8.14595
R1561 VDD2.n47 VDD2.n45 7.3702
R1562 VDD2.n12 VDD2.n10 7.3702
R1563 VDD2.n50 VDD2.n45 5.81868
R1564 VDD2.n15 VDD2.n10 5.81868
R1565 VDD2.n67 VDD2.n35 5.3904
R1566 VDD2.n32 VDD2.n0 5.3904
R1567 VDD2.n51 VDD2.n43 5.04292
R1568 VDD2.n16 VDD2.n8 5.04292
R1569 VDD2.n55 VDD2.n54 4.26717
R1570 VDD2.n20 VDD2.n19 4.26717
R1571 VDD2.n58 VDD2.n41 3.49141
R1572 VDD2.n23 VDD2.n6 3.49141
R1573 VDD2.n46 VDD2.n44 2.84305
R1574 VDD2.n11 VDD2.n9 2.84305
R1575 VDD2.n59 VDD2.n39 2.71565
R1576 VDD2.n24 VDD2.n4 2.71565
R1577 VDD2.n63 VDD2.n62 1.93989
R1578 VDD2.n28 VDD2.n27 1.93989
R1579 VDD2.n66 VDD2.n37 1.16414
R1580 VDD2.n31 VDD2.n2 1.16414
R1581 VDD2 VDD2.n70 0.974638
R1582 VDD2.n68 VDD2.n36 0.155672
R1583 VDD2.n61 VDD2.n36 0.155672
R1584 VDD2.n61 VDD2.n60 0.155672
R1585 VDD2.n60 VDD2.n40 0.155672
R1586 VDD2.n53 VDD2.n40 0.155672
R1587 VDD2.n53 VDD2.n52 0.155672
R1588 VDD2.n52 VDD2.n44 0.155672
R1589 VDD2.n17 VDD2.n9 0.155672
R1590 VDD2.n18 VDD2.n17 0.155672
R1591 VDD2.n18 VDD2.n5 0.155672
R1592 VDD2.n25 VDD2.n5 0.155672
R1593 VDD2.n26 VDD2.n25 0.155672
R1594 VDD2.n26 VDD2.n1 0.155672
R1595 VDD2.n33 VDD2.n1 0.155672
C0 VDD1 VN 0.148729f
C1 VDD2 VP 0.387878f
C2 VDD2 VTAIL 4.22205f
C3 VDD2 VDD1 0.822843f
C4 VDD2 VN 1.86724f
C5 VP VTAIL 1.86415f
C6 VP VDD1 2.10531f
C7 VTAIL VDD1 4.16084f
C8 VP VN 5.19214f
C9 VTAIL VN 1.84957f
C10 VDD2 B 3.999734f
C11 VDD1 B 6.79048f
C12 VTAIL B 5.951669f
C13 VN B 9.680889f
C14 VP B 7.697283f
C15 VDD2.n0 B 0.019966f
C16 VDD2.n1 B 0.014607f
C17 VDD2.n2 B 0.007849f
C18 VDD2.n3 B 0.018552f
C19 VDD2.n4 B 0.008311f
C20 VDD2.n5 B 0.014607f
C21 VDD2.n6 B 0.007849f
C22 VDD2.n7 B 0.018552f
C23 VDD2.n8 B 0.008311f
C24 VDD2.n9 B 0.426927f
C25 VDD2.n10 B 0.007849f
C26 VDD2.t1 B 0.030978f
C27 VDD2.n11 B 0.078598f
C28 VDD2.n12 B 0.013115f
C29 VDD2.n13 B 0.013914f
C30 VDD2.n14 B 0.018552f
C31 VDD2.n15 B 0.008311f
C32 VDD2.n16 B 0.007849f
C33 VDD2.n17 B 0.014607f
C34 VDD2.n18 B 0.014607f
C35 VDD2.n19 B 0.007849f
C36 VDD2.n20 B 0.008311f
C37 VDD2.n21 B 0.018552f
C38 VDD2.n22 B 0.018552f
C39 VDD2.n23 B 0.008311f
C40 VDD2.n24 B 0.007849f
C41 VDD2.n25 B 0.014607f
C42 VDD2.n26 B 0.014607f
C43 VDD2.n27 B 0.007849f
C44 VDD2.n28 B 0.008311f
C45 VDD2.n29 B 0.018552f
C46 VDD2.n30 B 0.037962f
C47 VDD2.n31 B 0.008311f
C48 VDD2.n32 B 0.015347f
C49 VDD2.n33 B 0.036756f
C50 VDD2.n34 B 0.388646f
C51 VDD2.n35 B 0.019966f
C52 VDD2.n36 B 0.014607f
C53 VDD2.n37 B 0.007849f
C54 VDD2.n38 B 0.018552f
C55 VDD2.n39 B 0.008311f
C56 VDD2.n40 B 0.014607f
C57 VDD2.n41 B 0.007849f
C58 VDD2.n42 B 0.018552f
C59 VDD2.n43 B 0.008311f
C60 VDD2.n44 B 0.426927f
C61 VDD2.n45 B 0.007849f
C62 VDD2.t0 B 0.030978f
C63 VDD2.n46 B 0.078598f
C64 VDD2.n47 B 0.013115f
C65 VDD2.n48 B 0.013914f
C66 VDD2.n49 B 0.018552f
C67 VDD2.n50 B 0.008311f
C68 VDD2.n51 B 0.007849f
C69 VDD2.n52 B 0.014607f
C70 VDD2.n53 B 0.014607f
C71 VDD2.n54 B 0.007849f
C72 VDD2.n55 B 0.008311f
C73 VDD2.n56 B 0.018552f
C74 VDD2.n57 B 0.018552f
C75 VDD2.n58 B 0.008311f
C76 VDD2.n59 B 0.007849f
C77 VDD2.n60 B 0.014607f
C78 VDD2.n61 B 0.014607f
C79 VDD2.n62 B 0.007849f
C80 VDD2.n63 B 0.008311f
C81 VDD2.n64 B 0.018552f
C82 VDD2.n65 B 0.037962f
C83 VDD2.n66 B 0.008311f
C84 VDD2.n67 B 0.015347f
C85 VDD2.n68 B 0.036756f
C86 VDD2.n69 B 0.049246f
C87 VDD2.n70 B 1.65837f
C88 VN.t0 B 1.42175f
C89 VN.t1 B 1.8356f
C90 VDD1.n0 B 0.029569f
C91 VDD1.n1 B 0.021632f
C92 VDD1.n2 B 0.011624f
C93 VDD1.n3 B 0.027475f
C94 VDD1.n4 B 0.012308f
C95 VDD1.n5 B 0.021632f
C96 VDD1.n6 B 0.011624f
C97 VDD1.n7 B 0.027475f
C98 VDD1.n8 B 0.012308f
C99 VDD1.n9 B 0.632269f
C100 VDD1.n10 B 0.011624f
C101 VDD1.t1 B 0.045878f
C102 VDD1.n11 B 0.116402f
C103 VDD1.n12 B 0.019423f
C104 VDD1.n13 B 0.020606f
C105 VDD1.n14 B 0.027475f
C106 VDD1.n15 B 0.012308f
C107 VDD1.n16 B 0.011624f
C108 VDD1.n17 B 0.021632f
C109 VDD1.n18 B 0.021632f
C110 VDD1.n19 B 0.011624f
C111 VDD1.n20 B 0.012308f
C112 VDD1.n21 B 0.027475f
C113 VDD1.n22 B 0.027475f
C114 VDD1.n23 B 0.012308f
C115 VDD1.n24 B 0.011624f
C116 VDD1.n25 B 0.021632f
C117 VDD1.n26 B 0.021632f
C118 VDD1.n27 B 0.011624f
C119 VDD1.n28 B 0.012308f
C120 VDD1.n29 B 0.027475f
C121 VDD1.n30 B 0.056221f
C122 VDD1.n31 B 0.012308f
C123 VDD1.n32 B 0.022729f
C124 VDD1.n33 B 0.054434f
C125 VDD1.n34 B 0.075002f
C126 VDD1.n35 B 0.029569f
C127 VDD1.n36 B 0.021632f
C128 VDD1.n37 B 0.011624f
C129 VDD1.n38 B 0.027475f
C130 VDD1.n39 B 0.012308f
C131 VDD1.n40 B 0.021632f
C132 VDD1.n41 B 0.011624f
C133 VDD1.n42 B 0.027475f
C134 VDD1.n43 B 0.012308f
C135 VDD1.n44 B 0.632269f
C136 VDD1.n45 B 0.011624f
C137 VDD1.t0 B 0.045878f
C138 VDD1.n46 B 0.116402f
C139 VDD1.n47 B 0.019423f
C140 VDD1.n48 B 0.020606f
C141 VDD1.n49 B 0.027475f
C142 VDD1.n50 B 0.012308f
C143 VDD1.n51 B 0.011624f
C144 VDD1.n52 B 0.021632f
C145 VDD1.n53 B 0.021632f
C146 VDD1.n54 B 0.011624f
C147 VDD1.n55 B 0.012308f
C148 VDD1.n56 B 0.027475f
C149 VDD1.n57 B 0.027475f
C150 VDD1.n58 B 0.012308f
C151 VDD1.n59 B 0.011624f
C152 VDD1.n60 B 0.021632f
C153 VDD1.n61 B 0.021632f
C154 VDD1.n62 B 0.011624f
C155 VDD1.n63 B 0.012308f
C156 VDD1.n64 B 0.027475f
C157 VDD1.n65 B 0.056221f
C158 VDD1.n66 B 0.012308f
C159 VDD1.n67 B 0.022729f
C160 VDD1.n68 B 0.054434f
C161 VDD1.n69 B 0.622728f
C162 VTAIL.n0 B 0.022094f
C163 VTAIL.n1 B 0.016163f
C164 VTAIL.n2 B 0.008686f
C165 VTAIL.n3 B 0.020529f
C166 VTAIL.n4 B 0.009196f
C167 VTAIL.n5 B 0.016163f
C168 VTAIL.n6 B 0.008686f
C169 VTAIL.n7 B 0.020529f
C170 VTAIL.n8 B 0.009196f
C171 VTAIL.n9 B 0.472428f
C172 VTAIL.n10 B 0.008686f
C173 VTAIL.t3 B 0.034279f
C174 VTAIL.n11 B 0.086975f
C175 VTAIL.n12 B 0.014513f
C176 VTAIL.n13 B 0.015397f
C177 VTAIL.n14 B 0.020529f
C178 VTAIL.n15 B 0.009196f
C179 VTAIL.n16 B 0.008686f
C180 VTAIL.n17 B 0.016163f
C181 VTAIL.n18 B 0.016163f
C182 VTAIL.n19 B 0.008686f
C183 VTAIL.n20 B 0.009196f
C184 VTAIL.n21 B 0.020529f
C185 VTAIL.n22 B 0.020529f
C186 VTAIL.n23 B 0.009196f
C187 VTAIL.n24 B 0.008686f
C188 VTAIL.n25 B 0.016163f
C189 VTAIL.n26 B 0.016163f
C190 VTAIL.n27 B 0.008686f
C191 VTAIL.n28 B 0.009196f
C192 VTAIL.n29 B 0.020529f
C193 VTAIL.n30 B 0.042008f
C194 VTAIL.n31 B 0.009196f
C195 VTAIL.n32 B 0.016983f
C196 VTAIL.n33 B 0.040673f
C197 VTAIL.n34 B 0.043358f
C198 VTAIL.n35 B 1.0167f
C199 VTAIL.n36 B 0.022094f
C200 VTAIL.n37 B 0.016163f
C201 VTAIL.n38 B 0.008686f
C202 VTAIL.n39 B 0.020529f
C203 VTAIL.n40 B 0.009196f
C204 VTAIL.n41 B 0.016163f
C205 VTAIL.n42 B 0.008686f
C206 VTAIL.n43 B 0.020529f
C207 VTAIL.n44 B 0.009196f
C208 VTAIL.n45 B 0.472428f
C209 VTAIL.n46 B 0.008686f
C210 VTAIL.t0 B 0.034279f
C211 VTAIL.n47 B 0.086975f
C212 VTAIL.n48 B 0.014513f
C213 VTAIL.n49 B 0.015397f
C214 VTAIL.n50 B 0.020529f
C215 VTAIL.n51 B 0.009196f
C216 VTAIL.n52 B 0.008686f
C217 VTAIL.n53 B 0.016163f
C218 VTAIL.n54 B 0.016163f
C219 VTAIL.n55 B 0.008686f
C220 VTAIL.n56 B 0.009196f
C221 VTAIL.n57 B 0.020529f
C222 VTAIL.n58 B 0.020529f
C223 VTAIL.n59 B 0.009196f
C224 VTAIL.n60 B 0.008686f
C225 VTAIL.n61 B 0.016163f
C226 VTAIL.n62 B 0.016163f
C227 VTAIL.n63 B 0.008686f
C228 VTAIL.n64 B 0.009196f
C229 VTAIL.n65 B 0.020529f
C230 VTAIL.n66 B 0.042008f
C231 VTAIL.n67 B 0.009196f
C232 VTAIL.n68 B 0.016983f
C233 VTAIL.n69 B 0.040673f
C234 VTAIL.n70 B 0.043358f
C235 VTAIL.n71 B 1.06137f
C236 VTAIL.n72 B 0.022094f
C237 VTAIL.n73 B 0.016163f
C238 VTAIL.n74 B 0.008686f
C239 VTAIL.n75 B 0.020529f
C240 VTAIL.n76 B 0.009196f
C241 VTAIL.n77 B 0.016163f
C242 VTAIL.n78 B 0.008686f
C243 VTAIL.n79 B 0.020529f
C244 VTAIL.n80 B 0.009196f
C245 VTAIL.n81 B 0.472428f
C246 VTAIL.n82 B 0.008686f
C247 VTAIL.t2 B 0.034279f
C248 VTAIL.n83 B 0.086975f
C249 VTAIL.n84 B 0.014513f
C250 VTAIL.n85 B 0.015397f
C251 VTAIL.n86 B 0.020529f
C252 VTAIL.n87 B 0.009196f
C253 VTAIL.n88 B 0.008686f
C254 VTAIL.n89 B 0.016163f
C255 VTAIL.n90 B 0.016163f
C256 VTAIL.n91 B 0.008686f
C257 VTAIL.n92 B 0.009196f
C258 VTAIL.n93 B 0.020529f
C259 VTAIL.n94 B 0.020529f
C260 VTAIL.n95 B 0.009196f
C261 VTAIL.n96 B 0.008686f
C262 VTAIL.n97 B 0.016163f
C263 VTAIL.n98 B 0.016163f
C264 VTAIL.n99 B 0.008686f
C265 VTAIL.n100 B 0.009196f
C266 VTAIL.n101 B 0.020529f
C267 VTAIL.n102 B 0.042008f
C268 VTAIL.n103 B 0.009196f
C269 VTAIL.n104 B 0.016983f
C270 VTAIL.n105 B 0.040673f
C271 VTAIL.n106 B 0.043358f
C272 VTAIL.n107 B 0.870552f
C273 VTAIL.n108 B 0.022094f
C274 VTAIL.n109 B 0.016163f
C275 VTAIL.n110 B 0.008686f
C276 VTAIL.n111 B 0.020529f
C277 VTAIL.n112 B 0.009196f
C278 VTAIL.n113 B 0.016163f
C279 VTAIL.n114 B 0.008686f
C280 VTAIL.n115 B 0.020529f
C281 VTAIL.n116 B 0.009196f
C282 VTAIL.n117 B 0.472428f
C283 VTAIL.n118 B 0.008686f
C284 VTAIL.t1 B 0.034279f
C285 VTAIL.n119 B 0.086975f
C286 VTAIL.n120 B 0.014513f
C287 VTAIL.n121 B 0.015397f
C288 VTAIL.n122 B 0.020529f
C289 VTAIL.n123 B 0.009196f
C290 VTAIL.n124 B 0.008686f
C291 VTAIL.n125 B 0.016163f
C292 VTAIL.n126 B 0.016163f
C293 VTAIL.n127 B 0.008686f
C294 VTAIL.n128 B 0.009196f
C295 VTAIL.n129 B 0.020529f
C296 VTAIL.n130 B 0.020529f
C297 VTAIL.n131 B 0.009196f
C298 VTAIL.n132 B 0.008686f
C299 VTAIL.n133 B 0.016163f
C300 VTAIL.n134 B 0.016163f
C301 VTAIL.n135 B 0.008686f
C302 VTAIL.n136 B 0.009196f
C303 VTAIL.n137 B 0.020529f
C304 VTAIL.n138 B 0.042008f
C305 VTAIL.n139 B 0.009196f
C306 VTAIL.n140 B 0.016983f
C307 VTAIL.n141 B 0.040673f
C308 VTAIL.n142 B 0.043358f
C309 VTAIL.n143 B 0.795347f
C310 VP.t0 B 2.58909f
C311 VP.t1 B 1.99951f
C312 VP.n0 B 2.61511f
.ends

