* NGSPICE file created from diff_pair_sample_1702.ext - technology: sky130A

.subckt diff_pair_sample_1702 VTAIL VN VP B VDD2 VDD1
X0 B.t23 B.t21 B.t22 B.t18 sky130_fd_pr__nfet_01v8 ad=7.1136 pd=37.26 as=0 ps=0 w=18.24 l=1.87
X1 VDD2.t9 VN.t0 VTAIL.t16 B.t8 sky130_fd_pr__nfet_01v8 ad=3.0096 pd=18.57 as=7.1136 ps=37.26 w=18.24 l=1.87
X2 VDD2.t8 VN.t1 VTAIL.t10 B.t6 sky130_fd_pr__nfet_01v8 ad=7.1136 pd=37.26 as=3.0096 ps=18.57 w=18.24 l=1.87
X3 VDD1.t9 VP.t0 VTAIL.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=3.0096 pd=18.57 as=3.0096 ps=18.57 w=18.24 l=1.87
X4 VDD1.t8 VP.t1 VTAIL.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=3.0096 pd=18.57 as=3.0096 ps=18.57 w=18.24 l=1.87
X5 VTAIL.t0 VP.t2 VDD1.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=3.0096 pd=18.57 as=3.0096 ps=18.57 w=18.24 l=1.87
X6 VTAIL.t12 VN.t2 VDD2.t7 B.t0 sky130_fd_pr__nfet_01v8 ad=3.0096 pd=18.57 as=3.0096 ps=18.57 w=18.24 l=1.87
X7 VDD2.t6 VN.t3 VTAIL.t18 B.t5 sky130_fd_pr__nfet_01v8 ad=7.1136 pd=37.26 as=3.0096 ps=18.57 w=18.24 l=1.87
X8 B.t20 B.t17 B.t19 B.t18 sky130_fd_pr__nfet_01v8 ad=7.1136 pd=37.26 as=0 ps=0 w=18.24 l=1.87
X9 VTAIL.t15 VN.t4 VDD2.t5 B.t9 sky130_fd_pr__nfet_01v8 ad=3.0096 pd=18.57 as=3.0096 ps=18.57 w=18.24 l=1.87
X10 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=7.1136 pd=37.26 as=0 ps=0 w=18.24 l=1.87
X11 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=7.1136 pd=37.26 as=0 ps=0 w=18.24 l=1.87
X12 VTAIL.t9 VP.t3 VDD1.t6 B.t9 sky130_fd_pr__nfet_01v8 ad=3.0096 pd=18.57 as=3.0096 ps=18.57 w=18.24 l=1.87
X13 VDD2.t4 VN.t5 VTAIL.t14 B.t4 sky130_fd_pr__nfet_01v8 ad=3.0096 pd=18.57 as=3.0096 ps=18.57 w=18.24 l=1.87
X14 VTAIL.t8 VP.t4 VDD1.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=3.0096 pd=18.57 as=3.0096 ps=18.57 w=18.24 l=1.87
X15 VTAIL.t19 VN.t6 VDD2.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=3.0096 pd=18.57 as=3.0096 ps=18.57 w=18.24 l=1.87
X16 VDD2.t2 VN.t7 VTAIL.t17 B.t2 sky130_fd_pr__nfet_01v8 ad=3.0096 pd=18.57 as=3.0096 ps=18.57 w=18.24 l=1.87
X17 VDD2.t1 VN.t8 VTAIL.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=3.0096 pd=18.57 as=7.1136 ps=37.26 w=18.24 l=1.87
X18 VDD1.t4 VP.t5 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=7.1136 pd=37.26 as=3.0096 ps=18.57 w=18.24 l=1.87
X19 VDD1.t3 VP.t6 VTAIL.t3 B.t7 sky130_fd_pr__nfet_01v8 ad=3.0096 pd=18.57 as=7.1136 ps=37.26 w=18.24 l=1.87
X20 VDD1.t2 VP.t7 VTAIL.t4 B.t8 sky130_fd_pr__nfet_01v8 ad=3.0096 pd=18.57 as=7.1136 ps=37.26 w=18.24 l=1.87
X21 VTAIL.t13 VN.t9 VDD2.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=3.0096 pd=18.57 as=3.0096 ps=18.57 w=18.24 l=1.87
X22 VTAIL.t2 VP.t8 VDD1.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=3.0096 pd=18.57 as=3.0096 ps=18.57 w=18.24 l=1.87
X23 VDD1.t0 VP.t9 VTAIL.t7 B.t5 sky130_fd_pr__nfet_01v8 ad=7.1136 pd=37.26 as=3.0096 ps=18.57 w=18.24 l=1.87
R0 B.n1036 B.n1035 585
R1 B.n412 B.n152 585
R2 B.n411 B.n410 585
R3 B.n409 B.n408 585
R4 B.n407 B.n406 585
R5 B.n405 B.n404 585
R6 B.n403 B.n402 585
R7 B.n401 B.n400 585
R8 B.n399 B.n398 585
R9 B.n397 B.n396 585
R10 B.n395 B.n394 585
R11 B.n393 B.n392 585
R12 B.n391 B.n390 585
R13 B.n389 B.n388 585
R14 B.n387 B.n386 585
R15 B.n385 B.n384 585
R16 B.n383 B.n382 585
R17 B.n381 B.n380 585
R18 B.n379 B.n378 585
R19 B.n377 B.n376 585
R20 B.n375 B.n374 585
R21 B.n373 B.n372 585
R22 B.n371 B.n370 585
R23 B.n369 B.n368 585
R24 B.n367 B.n366 585
R25 B.n365 B.n364 585
R26 B.n363 B.n362 585
R27 B.n361 B.n360 585
R28 B.n359 B.n358 585
R29 B.n357 B.n356 585
R30 B.n355 B.n354 585
R31 B.n353 B.n352 585
R32 B.n351 B.n350 585
R33 B.n349 B.n348 585
R34 B.n347 B.n346 585
R35 B.n345 B.n344 585
R36 B.n343 B.n342 585
R37 B.n341 B.n340 585
R38 B.n339 B.n338 585
R39 B.n337 B.n336 585
R40 B.n335 B.n334 585
R41 B.n333 B.n332 585
R42 B.n331 B.n330 585
R43 B.n329 B.n328 585
R44 B.n327 B.n326 585
R45 B.n325 B.n324 585
R46 B.n323 B.n322 585
R47 B.n321 B.n320 585
R48 B.n319 B.n318 585
R49 B.n317 B.n316 585
R50 B.n315 B.n314 585
R51 B.n313 B.n312 585
R52 B.n311 B.n310 585
R53 B.n309 B.n308 585
R54 B.n307 B.n306 585
R55 B.n305 B.n304 585
R56 B.n303 B.n302 585
R57 B.n301 B.n300 585
R58 B.n299 B.n298 585
R59 B.n297 B.n296 585
R60 B.n295 B.n294 585
R61 B.n293 B.n292 585
R62 B.n291 B.n290 585
R63 B.n289 B.n288 585
R64 B.n287 B.n286 585
R65 B.n285 B.n284 585
R66 B.n283 B.n282 585
R67 B.n281 B.n280 585
R68 B.n279 B.n278 585
R69 B.n277 B.n276 585
R70 B.n275 B.n274 585
R71 B.n273 B.n272 585
R72 B.n271 B.n270 585
R73 B.n269 B.n268 585
R74 B.n267 B.n266 585
R75 B.n265 B.n264 585
R76 B.n263 B.n262 585
R77 B.n261 B.n260 585
R78 B.n259 B.n258 585
R79 B.n257 B.n256 585
R80 B.n255 B.n254 585
R81 B.n253 B.n252 585
R82 B.n251 B.n250 585
R83 B.n249 B.n248 585
R84 B.n247 B.n246 585
R85 B.n245 B.n244 585
R86 B.n243 B.n242 585
R87 B.n241 B.n240 585
R88 B.n239 B.n238 585
R89 B.n237 B.n236 585
R90 B.n235 B.n234 585
R91 B.n233 B.n232 585
R92 B.n231 B.n230 585
R93 B.n229 B.n228 585
R94 B.n227 B.n226 585
R95 B.n225 B.n224 585
R96 B.n223 B.n222 585
R97 B.n221 B.n220 585
R98 B.n219 B.n218 585
R99 B.n217 B.n216 585
R100 B.n215 B.n214 585
R101 B.n213 B.n212 585
R102 B.n211 B.n210 585
R103 B.n209 B.n208 585
R104 B.n207 B.n206 585
R105 B.n205 B.n204 585
R106 B.n203 B.n202 585
R107 B.n201 B.n200 585
R108 B.n199 B.n198 585
R109 B.n197 B.n196 585
R110 B.n195 B.n194 585
R111 B.n193 B.n192 585
R112 B.n191 B.n190 585
R113 B.n189 B.n188 585
R114 B.n187 B.n186 585
R115 B.n185 B.n184 585
R116 B.n183 B.n182 585
R117 B.n181 B.n180 585
R118 B.n179 B.n178 585
R119 B.n177 B.n176 585
R120 B.n175 B.n174 585
R121 B.n173 B.n172 585
R122 B.n171 B.n170 585
R123 B.n169 B.n168 585
R124 B.n167 B.n166 585
R125 B.n165 B.n164 585
R126 B.n163 B.n162 585
R127 B.n161 B.n160 585
R128 B.n88 B.n87 585
R129 B.n1041 B.n1040 585
R130 B.n1034 B.n153 585
R131 B.n153 B.n85 585
R132 B.n1033 B.n84 585
R133 B.n1045 B.n84 585
R134 B.n1032 B.n83 585
R135 B.n1046 B.n83 585
R136 B.n1031 B.n82 585
R137 B.n1047 B.n82 585
R138 B.n1030 B.n1029 585
R139 B.n1029 B.n78 585
R140 B.n1028 B.n77 585
R141 B.n1053 B.n77 585
R142 B.n1027 B.n76 585
R143 B.n1054 B.n76 585
R144 B.n1026 B.n75 585
R145 B.n1055 B.n75 585
R146 B.n1025 B.n1024 585
R147 B.n1024 B.n71 585
R148 B.n1023 B.n70 585
R149 B.n1061 B.n70 585
R150 B.n1022 B.n69 585
R151 B.n1062 B.n69 585
R152 B.n1021 B.n68 585
R153 B.n1063 B.n68 585
R154 B.n1020 B.n1019 585
R155 B.n1019 B.n64 585
R156 B.n1018 B.n63 585
R157 B.n1069 B.n63 585
R158 B.n1017 B.n62 585
R159 B.n1070 B.n62 585
R160 B.n1016 B.n61 585
R161 B.n1071 B.n61 585
R162 B.n1015 B.n1014 585
R163 B.n1014 B.n60 585
R164 B.n1013 B.n56 585
R165 B.n1077 B.n56 585
R166 B.n1012 B.n55 585
R167 B.n1078 B.n55 585
R168 B.n1011 B.n54 585
R169 B.n1079 B.n54 585
R170 B.n1010 B.n1009 585
R171 B.n1009 B.n50 585
R172 B.n1008 B.n49 585
R173 B.n1085 B.n49 585
R174 B.n1007 B.n48 585
R175 B.n1086 B.n48 585
R176 B.n1006 B.n47 585
R177 B.n1087 B.n47 585
R178 B.n1005 B.n1004 585
R179 B.n1004 B.n43 585
R180 B.n1003 B.n42 585
R181 B.n1093 B.n42 585
R182 B.n1002 B.n41 585
R183 B.n1094 B.n41 585
R184 B.n1001 B.n40 585
R185 B.n1095 B.n40 585
R186 B.n1000 B.n999 585
R187 B.n999 B.n36 585
R188 B.n998 B.n35 585
R189 B.n1101 B.n35 585
R190 B.n997 B.n34 585
R191 B.n1102 B.n34 585
R192 B.n996 B.n33 585
R193 B.n1103 B.n33 585
R194 B.n995 B.n994 585
R195 B.n994 B.n29 585
R196 B.n993 B.n28 585
R197 B.n1109 B.n28 585
R198 B.n992 B.n27 585
R199 B.n1110 B.n27 585
R200 B.n991 B.n26 585
R201 B.n1111 B.n26 585
R202 B.n990 B.n989 585
R203 B.n989 B.n22 585
R204 B.n988 B.n21 585
R205 B.n1117 B.n21 585
R206 B.n987 B.n20 585
R207 B.n1118 B.n20 585
R208 B.n986 B.n19 585
R209 B.n1119 B.n19 585
R210 B.n985 B.n984 585
R211 B.n984 B.n15 585
R212 B.n983 B.n14 585
R213 B.n1125 B.n14 585
R214 B.n982 B.n13 585
R215 B.n1126 B.n13 585
R216 B.n981 B.n12 585
R217 B.n1127 B.n12 585
R218 B.n980 B.n979 585
R219 B.n979 B.n8 585
R220 B.n978 B.n7 585
R221 B.n1133 B.n7 585
R222 B.n977 B.n6 585
R223 B.n1134 B.n6 585
R224 B.n976 B.n5 585
R225 B.n1135 B.n5 585
R226 B.n975 B.n974 585
R227 B.n974 B.n4 585
R228 B.n973 B.n413 585
R229 B.n973 B.n972 585
R230 B.n963 B.n414 585
R231 B.n415 B.n414 585
R232 B.n965 B.n964 585
R233 B.n966 B.n965 585
R234 B.n962 B.n419 585
R235 B.n423 B.n419 585
R236 B.n961 B.n960 585
R237 B.n960 B.n959 585
R238 B.n421 B.n420 585
R239 B.n422 B.n421 585
R240 B.n952 B.n951 585
R241 B.n953 B.n952 585
R242 B.n950 B.n428 585
R243 B.n428 B.n427 585
R244 B.n949 B.n948 585
R245 B.n948 B.n947 585
R246 B.n430 B.n429 585
R247 B.n431 B.n430 585
R248 B.n940 B.n939 585
R249 B.n941 B.n940 585
R250 B.n938 B.n436 585
R251 B.n436 B.n435 585
R252 B.n937 B.n936 585
R253 B.n936 B.n935 585
R254 B.n438 B.n437 585
R255 B.n439 B.n438 585
R256 B.n928 B.n927 585
R257 B.n929 B.n928 585
R258 B.n926 B.n444 585
R259 B.n444 B.n443 585
R260 B.n925 B.n924 585
R261 B.n924 B.n923 585
R262 B.n446 B.n445 585
R263 B.n447 B.n446 585
R264 B.n916 B.n915 585
R265 B.n917 B.n916 585
R266 B.n914 B.n452 585
R267 B.n452 B.n451 585
R268 B.n913 B.n912 585
R269 B.n912 B.n911 585
R270 B.n454 B.n453 585
R271 B.n455 B.n454 585
R272 B.n904 B.n903 585
R273 B.n905 B.n904 585
R274 B.n902 B.n459 585
R275 B.n463 B.n459 585
R276 B.n901 B.n900 585
R277 B.n900 B.n899 585
R278 B.n461 B.n460 585
R279 B.n462 B.n461 585
R280 B.n892 B.n891 585
R281 B.n893 B.n892 585
R282 B.n890 B.n468 585
R283 B.n468 B.n467 585
R284 B.n889 B.n888 585
R285 B.n888 B.n887 585
R286 B.n470 B.n469 585
R287 B.n880 B.n470 585
R288 B.n879 B.n878 585
R289 B.n881 B.n879 585
R290 B.n877 B.n475 585
R291 B.n475 B.n474 585
R292 B.n876 B.n875 585
R293 B.n875 B.n874 585
R294 B.n477 B.n476 585
R295 B.n478 B.n477 585
R296 B.n867 B.n866 585
R297 B.n868 B.n867 585
R298 B.n865 B.n483 585
R299 B.n483 B.n482 585
R300 B.n864 B.n863 585
R301 B.n863 B.n862 585
R302 B.n485 B.n484 585
R303 B.n486 B.n485 585
R304 B.n855 B.n854 585
R305 B.n856 B.n855 585
R306 B.n853 B.n490 585
R307 B.n494 B.n490 585
R308 B.n852 B.n851 585
R309 B.n851 B.n850 585
R310 B.n492 B.n491 585
R311 B.n493 B.n492 585
R312 B.n843 B.n842 585
R313 B.n844 B.n843 585
R314 B.n841 B.n499 585
R315 B.n499 B.n498 585
R316 B.n840 B.n839 585
R317 B.n839 B.n838 585
R318 B.n501 B.n500 585
R319 B.n502 B.n501 585
R320 B.n834 B.n833 585
R321 B.n505 B.n504 585
R322 B.n830 B.n829 585
R323 B.n831 B.n830 585
R324 B.n828 B.n570 585
R325 B.n827 B.n826 585
R326 B.n825 B.n824 585
R327 B.n823 B.n822 585
R328 B.n821 B.n820 585
R329 B.n819 B.n818 585
R330 B.n817 B.n816 585
R331 B.n815 B.n814 585
R332 B.n813 B.n812 585
R333 B.n811 B.n810 585
R334 B.n809 B.n808 585
R335 B.n807 B.n806 585
R336 B.n805 B.n804 585
R337 B.n803 B.n802 585
R338 B.n801 B.n800 585
R339 B.n799 B.n798 585
R340 B.n797 B.n796 585
R341 B.n795 B.n794 585
R342 B.n793 B.n792 585
R343 B.n791 B.n790 585
R344 B.n789 B.n788 585
R345 B.n787 B.n786 585
R346 B.n785 B.n784 585
R347 B.n783 B.n782 585
R348 B.n781 B.n780 585
R349 B.n779 B.n778 585
R350 B.n777 B.n776 585
R351 B.n775 B.n774 585
R352 B.n773 B.n772 585
R353 B.n771 B.n770 585
R354 B.n769 B.n768 585
R355 B.n767 B.n766 585
R356 B.n765 B.n764 585
R357 B.n763 B.n762 585
R358 B.n761 B.n760 585
R359 B.n759 B.n758 585
R360 B.n757 B.n756 585
R361 B.n755 B.n754 585
R362 B.n753 B.n752 585
R363 B.n751 B.n750 585
R364 B.n749 B.n748 585
R365 B.n747 B.n746 585
R366 B.n745 B.n744 585
R367 B.n743 B.n742 585
R368 B.n741 B.n740 585
R369 B.n739 B.n738 585
R370 B.n737 B.n736 585
R371 B.n735 B.n734 585
R372 B.n733 B.n732 585
R373 B.n731 B.n730 585
R374 B.n729 B.n728 585
R375 B.n727 B.n726 585
R376 B.n725 B.n724 585
R377 B.n723 B.n722 585
R378 B.n721 B.n720 585
R379 B.n719 B.n718 585
R380 B.n717 B.n716 585
R381 B.n714 B.n713 585
R382 B.n712 B.n711 585
R383 B.n710 B.n709 585
R384 B.n708 B.n707 585
R385 B.n706 B.n705 585
R386 B.n704 B.n703 585
R387 B.n702 B.n701 585
R388 B.n700 B.n699 585
R389 B.n698 B.n697 585
R390 B.n696 B.n695 585
R391 B.n693 B.n692 585
R392 B.n691 B.n690 585
R393 B.n689 B.n688 585
R394 B.n687 B.n686 585
R395 B.n685 B.n684 585
R396 B.n683 B.n682 585
R397 B.n681 B.n680 585
R398 B.n679 B.n678 585
R399 B.n677 B.n676 585
R400 B.n675 B.n674 585
R401 B.n673 B.n672 585
R402 B.n671 B.n670 585
R403 B.n669 B.n668 585
R404 B.n667 B.n666 585
R405 B.n665 B.n664 585
R406 B.n663 B.n662 585
R407 B.n661 B.n660 585
R408 B.n659 B.n658 585
R409 B.n657 B.n656 585
R410 B.n655 B.n654 585
R411 B.n653 B.n652 585
R412 B.n651 B.n650 585
R413 B.n649 B.n648 585
R414 B.n647 B.n646 585
R415 B.n645 B.n644 585
R416 B.n643 B.n642 585
R417 B.n641 B.n640 585
R418 B.n639 B.n638 585
R419 B.n637 B.n636 585
R420 B.n635 B.n634 585
R421 B.n633 B.n632 585
R422 B.n631 B.n630 585
R423 B.n629 B.n628 585
R424 B.n627 B.n626 585
R425 B.n625 B.n624 585
R426 B.n623 B.n622 585
R427 B.n621 B.n620 585
R428 B.n619 B.n618 585
R429 B.n617 B.n616 585
R430 B.n615 B.n614 585
R431 B.n613 B.n612 585
R432 B.n611 B.n610 585
R433 B.n609 B.n608 585
R434 B.n607 B.n606 585
R435 B.n605 B.n604 585
R436 B.n603 B.n602 585
R437 B.n601 B.n600 585
R438 B.n599 B.n598 585
R439 B.n597 B.n596 585
R440 B.n595 B.n594 585
R441 B.n593 B.n592 585
R442 B.n591 B.n590 585
R443 B.n589 B.n588 585
R444 B.n587 B.n586 585
R445 B.n585 B.n584 585
R446 B.n583 B.n582 585
R447 B.n581 B.n580 585
R448 B.n579 B.n578 585
R449 B.n577 B.n576 585
R450 B.n575 B.n569 585
R451 B.n831 B.n569 585
R452 B.n835 B.n503 585
R453 B.n503 B.n502 585
R454 B.n837 B.n836 585
R455 B.n838 B.n837 585
R456 B.n497 B.n496 585
R457 B.n498 B.n497 585
R458 B.n846 B.n845 585
R459 B.n845 B.n844 585
R460 B.n847 B.n495 585
R461 B.n495 B.n493 585
R462 B.n849 B.n848 585
R463 B.n850 B.n849 585
R464 B.n489 B.n488 585
R465 B.n494 B.n489 585
R466 B.n858 B.n857 585
R467 B.n857 B.n856 585
R468 B.n859 B.n487 585
R469 B.n487 B.n486 585
R470 B.n861 B.n860 585
R471 B.n862 B.n861 585
R472 B.n481 B.n480 585
R473 B.n482 B.n481 585
R474 B.n870 B.n869 585
R475 B.n869 B.n868 585
R476 B.n871 B.n479 585
R477 B.n479 B.n478 585
R478 B.n873 B.n872 585
R479 B.n874 B.n873 585
R480 B.n473 B.n472 585
R481 B.n474 B.n473 585
R482 B.n883 B.n882 585
R483 B.n882 B.n881 585
R484 B.n884 B.n471 585
R485 B.n880 B.n471 585
R486 B.n886 B.n885 585
R487 B.n887 B.n886 585
R488 B.n466 B.n465 585
R489 B.n467 B.n466 585
R490 B.n895 B.n894 585
R491 B.n894 B.n893 585
R492 B.n896 B.n464 585
R493 B.n464 B.n462 585
R494 B.n898 B.n897 585
R495 B.n899 B.n898 585
R496 B.n458 B.n457 585
R497 B.n463 B.n458 585
R498 B.n907 B.n906 585
R499 B.n906 B.n905 585
R500 B.n908 B.n456 585
R501 B.n456 B.n455 585
R502 B.n910 B.n909 585
R503 B.n911 B.n910 585
R504 B.n450 B.n449 585
R505 B.n451 B.n450 585
R506 B.n919 B.n918 585
R507 B.n918 B.n917 585
R508 B.n920 B.n448 585
R509 B.n448 B.n447 585
R510 B.n922 B.n921 585
R511 B.n923 B.n922 585
R512 B.n442 B.n441 585
R513 B.n443 B.n442 585
R514 B.n931 B.n930 585
R515 B.n930 B.n929 585
R516 B.n932 B.n440 585
R517 B.n440 B.n439 585
R518 B.n934 B.n933 585
R519 B.n935 B.n934 585
R520 B.n434 B.n433 585
R521 B.n435 B.n434 585
R522 B.n943 B.n942 585
R523 B.n942 B.n941 585
R524 B.n944 B.n432 585
R525 B.n432 B.n431 585
R526 B.n946 B.n945 585
R527 B.n947 B.n946 585
R528 B.n426 B.n425 585
R529 B.n427 B.n426 585
R530 B.n955 B.n954 585
R531 B.n954 B.n953 585
R532 B.n956 B.n424 585
R533 B.n424 B.n422 585
R534 B.n958 B.n957 585
R535 B.n959 B.n958 585
R536 B.n418 B.n417 585
R537 B.n423 B.n418 585
R538 B.n968 B.n967 585
R539 B.n967 B.n966 585
R540 B.n969 B.n416 585
R541 B.n416 B.n415 585
R542 B.n971 B.n970 585
R543 B.n972 B.n971 585
R544 B.n2 B.n0 585
R545 B.n4 B.n2 585
R546 B.n3 B.n1 585
R547 B.n1134 B.n3 585
R548 B.n1132 B.n1131 585
R549 B.n1133 B.n1132 585
R550 B.n1130 B.n9 585
R551 B.n9 B.n8 585
R552 B.n1129 B.n1128 585
R553 B.n1128 B.n1127 585
R554 B.n11 B.n10 585
R555 B.n1126 B.n11 585
R556 B.n1124 B.n1123 585
R557 B.n1125 B.n1124 585
R558 B.n1122 B.n16 585
R559 B.n16 B.n15 585
R560 B.n1121 B.n1120 585
R561 B.n1120 B.n1119 585
R562 B.n18 B.n17 585
R563 B.n1118 B.n18 585
R564 B.n1116 B.n1115 585
R565 B.n1117 B.n1116 585
R566 B.n1114 B.n23 585
R567 B.n23 B.n22 585
R568 B.n1113 B.n1112 585
R569 B.n1112 B.n1111 585
R570 B.n25 B.n24 585
R571 B.n1110 B.n25 585
R572 B.n1108 B.n1107 585
R573 B.n1109 B.n1108 585
R574 B.n1106 B.n30 585
R575 B.n30 B.n29 585
R576 B.n1105 B.n1104 585
R577 B.n1104 B.n1103 585
R578 B.n32 B.n31 585
R579 B.n1102 B.n32 585
R580 B.n1100 B.n1099 585
R581 B.n1101 B.n1100 585
R582 B.n1098 B.n37 585
R583 B.n37 B.n36 585
R584 B.n1097 B.n1096 585
R585 B.n1096 B.n1095 585
R586 B.n39 B.n38 585
R587 B.n1094 B.n39 585
R588 B.n1092 B.n1091 585
R589 B.n1093 B.n1092 585
R590 B.n1090 B.n44 585
R591 B.n44 B.n43 585
R592 B.n1089 B.n1088 585
R593 B.n1088 B.n1087 585
R594 B.n46 B.n45 585
R595 B.n1086 B.n46 585
R596 B.n1084 B.n1083 585
R597 B.n1085 B.n1084 585
R598 B.n1082 B.n51 585
R599 B.n51 B.n50 585
R600 B.n1081 B.n1080 585
R601 B.n1080 B.n1079 585
R602 B.n53 B.n52 585
R603 B.n1078 B.n53 585
R604 B.n1076 B.n1075 585
R605 B.n1077 B.n1076 585
R606 B.n1074 B.n57 585
R607 B.n60 B.n57 585
R608 B.n1073 B.n1072 585
R609 B.n1072 B.n1071 585
R610 B.n59 B.n58 585
R611 B.n1070 B.n59 585
R612 B.n1068 B.n1067 585
R613 B.n1069 B.n1068 585
R614 B.n1066 B.n65 585
R615 B.n65 B.n64 585
R616 B.n1065 B.n1064 585
R617 B.n1064 B.n1063 585
R618 B.n67 B.n66 585
R619 B.n1062 B.n67 585
R620 B.n1060 B.n1059 585
R621 B.n1061 B.n1060 585
R622 B.n1058 B.n72 585
R623 B.n72 B.n71 585
R624 B.n1057 B.n1056 585
R625 B.n1056 B.n1055 585
R626 B.n74 B.n73 585
R627 B.n1054 B.n74 585
R628 B.n1052 B.n1051 585
R629 B.n1053 B.n1052 585
R630 B.n1050 B.n79 585
R631 B.n79 B.n78 585
R632 B.n1049 B.n1048 585
R633 B.n1048 B.n1047 585
R634 B.n81 B.n80 585
R635 B.n1046 B.n81 585
R636 B.n1044 B.n1043 585
R637 B.n1045 B.n1044 585
R638 B.n1042 B.n86 585
R639 B.n86 B.n85 585
R640 B.n1137 B.n1136 585
R641 B.n1136 B.n1135 585
R642 B.n833 B.n503 449.257
R643 B.n1040 B.n86 449.257
R644 B.n569 B.n501 449.257
R645 B.n1036 B.n153 449.257
R646 B.n573 B.t10 441.668
R647 B.n571 B.t14 441.668
R648 B.n157 B.t17 441.668
R649 B.n154 B.t21 441.668
R650 B.n573 B.t13 432.413
R651 B.n154 B.t22 432.413
R652 B.n571 B.t16 432.413
R653 B.n157 B.t19 432.413
R654 B.n574 B.t12 389.748
R655 B.n155 B.t23 389.748
R656 B.n572 B.t15 389.748
R657 B.n158 B.t20 389.748
R658 B.n1038 B.n1037 256.663
R659 B.n1038 B.n151 256.663
R660 B.n1038 B.n150 256.663
R661 B.n1038 B.n149 256.663
R662 B.n1038 B.n148 256.663
R663 B.n1038 B.n147 256.663
R664 B.n1038 B.n146 256.663
R665 B.n1038 B.n145 256.663
R666 B.n1038 B.n144 256.663
R667 B.n1038 B.n143 256.663
R668 B.n1038 B.n142 256.663
R669 B.n1038 B.n141 256.663
R670 B.n1038 B.n140 256.663
R671 B.n1038 B.n139 256.663
R672 B.n1038 B.n138 256.663
R673 B.n1038 B.n137 256.663
R674 B.n1038 B.n136 256.663
R675 B.n1038 B.n135 256.663
R676 B.n1038 B.n134 256.663
R677 B.n1038 B.n133 256.663
R678 B.n1038 B.n132 256.663
R679 B.n1038 B.n131 256.663
R680 B.n1038 B.n130 256.663
R681 B.n1038 B.n129 256.663
R682 B.n1038 B.n128 256.663
R683 B.n1038 B.n127 256.663
R684 B.n1038 B.n126 256.663
R685 B.n1038 B.n125 256.663
R686 B.n1038 B.n124 256.663
R687 B.n1038 B.n123 256.663
R688 B.n1038 B.n122 256.663
R689 B.n1038 B.n121 256.663
R690 B.n1038 B.n120 256.663
R691 B.n1038 B.n119 256.663
R692 B.n1038 B.n118 256.663
R693 B.n1038 B.n117 256.663
R694 B.n1038 B.n116 256.663
R695 B.n1038 B.n115 256.663
R696 B.n1038 B.n114 256.663
R697 B.n1038 B.n113 256.663
R698 B.n1038 B.n112 256.663
R699 B.n1038 B.n111 256.663
R700 B.n1038 B.n110 256.663
R701 B.n1038 B.n109 256.663
R702 B.n1038 B.n108 256.663
R703 B.n1038 B.n107 256.663
R704 B.n1038 B.n106 256.663
R705 B.n1038 B.n105 256.663
R706 B.n1038 B.n104 256.663
R707 B.n1038 B.n103 256.663
R708 B.n1038 B.n102 256.663
R709 B.n1038 B.n101 256.663
R710 B.n1038 B.n100 256.663
R711 B.n1038 B.n99 256.663
R712 B.n1038 B.n98 256.663
R713 B.n1038 B.n97 256.663
R714 B.n1038 B.n96 256.663
R715 B.n1038 B.n95 256.663
R716 B.n1038 B.n94 256.663
R717 B.n1038 B.n93 256.663
R718 B.n1038 B.n92 256.663
R719 B.n1038 B.n91 256.663
R720 B.n1038 B.n90 256.663
R721 B.n1038 B.n89 256.663
R722 B.n1039 B.n1038 256.663
R723 B.n832 B.n831 256.663
R724 B.n831 B.n506 256.663
R725 B.n831 B.n507 256.663
R726 B.n831 B.n508 256.663
R727 B.n831 B.n509 256.663
R728 B.n831 B.n510 256.663
R729 B.n831 B.n511 256.663
R730 B.n831 B.n512 256.663
R731 B.n831 B.n513 256.663
R732 B.n831 B.n514 256.663
R733 B.n831 B.n515 256.663
R734 B.n831 B.n516 256.663
R735 B.n831 B.n517 256.663
R736 B.n831 B.n518 256.663
R737 B.n831 B.n519 256.663
R738 B.n831 B.n520 256.663
R739 B.n831 B.n521 256.663
R740 B.n831 B.n522 256.663
R741 B.n831 B.n523 256.663
R742 B.n831 B.n524 256.663
R743 B.n831 B.n525 256.663
R744 B.n831 B.n526 256.663
R745 B.n831 B.n527 256.663
R746 B.n831 B.n528 256.663
R747 B.n831 B.n529 256.663
R748 B.n831 B.n530 256.663
R749 B.n831 B.n531 256.663
R750 B.n831 B.n532 256.663
R751 B.n831 B.n533 256.663
R752 B.n831 B.n534 256.663
R753 B.n831 B.n535 256.663
R754 B.n831 B.n536 256.663
R755 B.n831 B.n537 256.663
R756 B.n831 B.n538 256.663
R757 B.n831 B.n539 256.663
R758 B.n831 B.n540 256.663
R759 B.n831 B.n541 256.663
R760 B.n831 B.n542 256.663
R761 B.n831 B.n543 256.663
R762 B.n831 B.n544 256.663
R763 B.n831 B.n545 256.663
R764 B.n831 B.n546 256.663
R765 B.n831 B.n547 256.663
R766 B.n831 B.n548 256.663
R767 B.n831 B.n549 256.663
R768 B.n831 B.n550 256.663
R769 B.n831 B.n551 256.663
R770 B.n831 B.n552 256.663
R771 B.n831 B.n553 256.663
R772 B.n831 B.n554 256.663
R773 B.n831 B.n555 256.663
R774 B.n831 B.n556 256.663
R775 B.n831 B.n557 256.663
R776 B.n831 B.n558 256.663
R777 B.n831 B.n559 256.663
R778 B.n831 B.n560 256.663
R779 B.n831 B.n561 256.663
R780 B.n831 B.n562 256.663
R781 B.n831 B.n563 256.663
R782 B.n831 B.n564 256.663
R783 B.n831 B.n565 256.663
R784 B.n831 B.n566 256.663
R785 B.n831 B.n567 256.663
R786 B.n831 B.n568 256.663
R787 B.n837 B.n503 163.367
R788 B.n837 B.n497 163.367
R789 B.n845 B.n497 163.367
R790 B.n845 B.n495 163.367
R791 B.n849 B.n495 163.367
R792 B.n849 B.n489 163.367
R793 B.n857 B.n489 163.367
R794 B.n857 B.n487 163.367
R795 B.n861 B.n487 163.367
R796 B.n861 B.n481 163.367
R797 B.n869 B.n481 163.367
R798 B.n869 B.n479 163.367
R799 B.n873 B.n479 163.367
R800 B.n873 B.n473 163.367
R801 B.n882 B.n473 163.367
R802 B.n882 B.n471 163.367
R803 B.n886 B.n471 163.367
R804 B.n886 B.n466 163.367
R805 B.n894 B.n466 163.367
R806 B.n894 B.n464 163.367
R807 B.n898 B.n464 163.367
R808 B.n898 B.n458 163.367
R809 B.n906 B.n458 163.367
R810 B.n906 B.n456 163.367
R811 B.n910 B.n456 163.367
R812 B.n910 B.n450 163.367
R813 B.n918 B.n450 163.367
R814 B.n918 B.n448 163.367
R815 B.n922 B.n448 163.367
R816 B.n922 B.n442 163.367
R817 B.n930 B.n442 163.367
R818 B.n930 B.n440 163.367
R819 B.n934 B.n440 163.367
R820 B.n934 B.n434 163.367
R821 B.n942 B.n434 163.367
R822 B.n942 B.n432 163.367
R823 B.n946 B.n432 163.367
R824 B.n946 B.n426 163.367
R825 B.n954 B.n426 163.367
R826 B.n954 B.n424 163.367
R827 B.n958 B.n424 163.367
R828 B.n958 B.n418 163.367
R829 B.n967 B.n418 163.367
R830 B.n967 B.n416 163.367
R831 B.n971 B.n416 163.367
R832 B.n971 B.n2 163.367
R833 B.n1136 B.n2 163.367
R834 B.n1136 B.n3 163.367
R835 B.n1132 B.n3 163.367
R836 B.n1132 B.n9 163.367
R837 B.n1128 B.n9 163.367
R838 B.n1128 B.n11 163.367
R839 B.n1124 B.n11 163.367
R840 B.n1124 B.n16 163.367
R841 B.n1120 B.n16 163.367
R842 B.n1120 B.n18 163.367
R843 B.n1116 B.n18 163.367
R844 B.n1116 B.n23 163.367
R845 B.n1112 B.n23 163.367
R846 B.n1112 B.n25 163.367
R847 B.n1108 B.n25 163.367
R848 B.n1108 B.n30 163.367
R849 B.n1104 B.n30 163.367
R850 B.n1104 B.n32 163.367
R851 B.n1100 B.n32 163.367
R852 B.n1100 B.n37 163.367
R853 B.n1096 B.n37 163.367
R854 B.n1096 B.n39 163.367
R855 B.n1092 B.n39 163.367
R856 B.n1092 B.n44 163.367
R857 B.n1088 B.n44 163.367
R858 B.n1088 B.n46 163.367
R859 B.n1084 B.n46 163.367
R860 B.n1084 B.n51 163.367
R861 B.n1080 B.n51 163.367
R862 B.n1080 B.n53 163.367
R863 B.n1076 B.n53 163.367
R864 B.n1076 B.n57 163.367
R865 B.n1072 B.n57 163.367
R866 B.n1072 B.n59 163.367
R867 B.n1068 B.n59 163.367
R868 B.n1068 B.n65 163.367
R869 B.n1064 B.n65 163.367
R870 B.n1064 B.n67 163.367
R871 B.n1060 B.n67 163.367
R872 B.n1060 B.n72 163.367
R873 B.n1056 B.n72 163.367
R874 B.n1056 B.n74 163.367
R875 B.n1052 B.n74 163.367
R876 B.n1052 B.n79 163.367
R877 B.n1048 B.n79 163.367
R878 B.n1048 B.n81 163.367
R879 B.n1044 B.n81 163.367
R880 B.n1044 B.n86 163.367
R881 B.n830 B.n505 163.367
R882 B.n830 B.n570 163.367
R883 B.n826 B.n825 163.367
R884 B.n822 B.n821 163.367
R885 B.n818 B.n817 163.367
R886 B.n814 B.n813 163.367
R887 B.n810 B.n809 163.367
R888 B.n806 B.n805 163.367
R889 B.n802 B.n801 163.367
R890 B.n798 B.n797 163.367
R891 B.n794 B.n793 163.367
R892 B.n790 B.n789 163.367
R893 B.n786 B.n785 163.367
R894 B.n782 B.n781 163.367
R895 B.n778 B.n777 163.367
R896 B.n774 B.n773 163.367
R897 B.n770 B.n769 163.367
R898 B.n766 B.n765 163.367
R899 B.n762 B.n761 163.367
R900 B.n758 B.n757 163.367
R901 B.n754 B.n753 163.367
R902 B.n750 B.n749 163.367
R903 B.n746 B.n745 163.367
R904 B.n742 B.n741 163.367
R905 B.n738 B.n737 163.367
R906 B.n734 B.n733 163.367
R907 B.n730 B.n729 163.367
R908 B.n726 B.n725 163.367
R909 B.n722 B.n721 163.367
R910 B.n718 B.n717 163.367
R911 B.n713 B.n712 163.367
R912 B.n709 B.n708 163.367
R913 B.n705 B.n704 163.367
R914 B.n701 B.n700 163.367
R915 B.n697 B.n696 163.367
R916 B.n692 B.n691 163.367
R917 B.n688 B.n687 163.367
R918 B.n684 B.n683 163.367
R919 B.n680 B.n679 163.367
R920 B.n676 B.n675 163.367
R921 B.n672 B.n671 163.367
R922 B.n668 B.n667 163.367
R923 B.n664 B.n663 163.367
R924 B.n660 B.n659 163.367
R925 B.n656 B.n655 163.367
R926 B.n652 B.n651 163.367
R927 B.n648 B.n647 163.367
R928 B.n644 B.n643 163.367
R929 B.n640 B.n639 163.367
R930 B.n636 B.n635 163.367
R931 B.n632 B.n631 163.367
R932 B.n628 B.n627 163.367
R933 B.n624 B.n623 163.367
R934 B.n620 B.n619 163.367
R935 B.n616 B.n615 163.367
R936 B.n612 B.n611 163.367
R937 B.n608 B.n607 163.367
R938 B.n604 B.n603 163.367
R939 B.n600 B.n599 163.367
R940 B.n596 B.n595 163.367
R941 B.n592 B.n591 163.367
R942 B.n588 B.n587 163.367
R943 B.n584 B.n583 163.367
R944 B.n580 B.n579 163.367
R945 B.n576 B.n569 163.367
R946 B.n839 B.n501 163.367
R947 B.n839 B.n499 163.367
R948 B.n843 B.n499 163.367
R949 B.n843 B.n492 163.367
R950 B.n851 B.n492 163.367
R951 B.n851 B.n490 163.367
R952 B.n855 B.n490 163.367
R953 B.n855 B.n485 163.367
R954 B.n863 B.n485 163.367
R955 B.n863 B.n483 163.367
R956 B.n867 B.n483 163.367
R957 B.n867 B.n477 163.367
R958 B.n875 B.n477 163.367
R959 B.n875 B.n475 163.367
R960 B.n879 B.n475 163.367
R961 B.n879 B.n470 163.367
R962 B.n888 B.n470 163.367
R963 B.n888 B.n468 163.367
R964 B.n892 B.n468 163.367
R965 B.n892 B.n461 163.367
R966 B.n900 B.n461 163.367
R967 B.n900 B.n459 163.367
R968 B.n904 B.n459 163.367
R969 B.n904 B.n454 163.367
R970 B.n912 B.n454 163.367
R971 B.n912 B.n452 163.367
R972 B.n916 B.n452 163.367
R973 B.n916 B.n446 163.367
R974 B.n924 B.n446 163.367
R975 B.n924 B.n444 163.367
R976 B.n928 B.n444 163.367
R977 B.n928 B.n438 163.367
R978 B.n936 B.n438 163.367
R979 B.n936 B.n436 163.367
R980 B.n940 B.n436 163.367
R981 B.n940 B.n430 163.367
R982 B.n948 B.n430 163.367
R983 B.n948 B.n428 163.367
R984 B.n952 B.n428 163.367
R985 B.n952 B.n421 163.367
R986 B.n960 B.n421 163.367
R987 B.n960 B.n419 163.367
R988 B.n965 B.n419 163.367
R989 B.n965 B.n414 163.367
R990 B.n973 B.n414 163.367
R991 B.n974 B.n973 163.367
R992 B.n974 B.n5 163.367
R993 B.n6 B.n5 163.367
R994 B.n7 B.n6 163.367
R995 B.n979 B.n7 163.367
R996 B.n979 B.n12 163.367
R997 B.n13 B.n12 163.367
R998 B.n14 B.n13 163.367
R999 B.n984 B.n14 163.367
R1000 B.n984 B.n19 163.367
R1001 B.n20 B.n19 163.367
R1002 B.n21 B.n20 163.367
R1003 B.n989 B.n21 163.367
R1004 B.n989 B.n26 163.367
R1005 B.n27 B.n26 163.367
R1006 B.n28 B.n27 163.367
R1007 B.n994 B.n28 163.367
R1008 B.n994 B.n33 163.367
R1009 B.n34 B.n33 163.367
R1010 B.n35 B.n34 163.367
R1011 B.n999 B.n35 163.367
R1012 B.n999 B.n40 163.367
R1013 B.n41 B.n40 163.367
R1014 B.n42 B.n41 163.367
R1015 B.n1004 B.n42 163.367
R1016 B.n1004 B.n47 163.367
R1017 B.n48 B.n47 163.367
R1018 B.n49 B.n48 163.367
R1019 B.n1009 B.n49 163.367
R1020 B.n1009 B.n54 163.367
R1021 B.n55 B.n54 163.367
R1022 B.n56 B.n55 163.367
R1023 B.n1014 B.n56 163.367
R1024 B.n1014 B.n61 163.367
R1025 B.n62 B.n61 163.367
R1026 B.n63 B.n62 163.367
R1027 B.n1019 B.n63 163.367
R1028 B.n1019 B.n68 163.367
R1029 B.n69 B.n68 163.367
R1030 B.n70 B.n69 163.367
R1031 B.n1024 B.n70 163.367
R1032 B.n1024 B.n75 163.367
R1033 B.n76 B.n75 163.367
R1034 B.n77 B.n76 163.367
R1035 B.n1029 B.n77 163.367
R1036 B.n1029 B.n82 163.367
R1037 B.n83 B.n82 163.367
R1038 B.n84 B.n83 163.367
R1039 B.n153 B.n84 163.367
R1040 B.n160 B.n88 163.367
R1041 B.n164 B.n163 163.367
R1042 B.n168 B.n167 163.367
R1043 B.n172 B.n171 163.367
R1044 B.n176 B.n175 163.367
R1045 B.n180 B.n179 163.367
R1046 B.n184 B.n183 163.367
R1047 B.n188 B.n187 163.367
R1048 B.n192 B.n191 163.367
R1049 B.n196 B.n195 163.367
R1050 B.n200 B.n199 163.367
R1051 B.n204 B.n203 163.367
R1052 B.n208 B.n207 163.367
R1053 B.n212 B.n211 163.367
R1054 B.n216 B.n215 163.367
R1055 B.n220 B.n219 163.367
R1056 B.n224 B.n223 163.367
R1057 B.n228 B.n227 163.367
R1058 B.n232 B.n231 163.367
R1059 B.n236 B.n235 163.367
R1060 B.n240 B.n239 163.367
R1061 B.n244 B.n243 163.367
R1062 B.n248 B.n247 163.367
R1063 B.n252 B.n251 163.367
R1064 B.n256 B.n255 163.367
R1065 B.n260 B.n259 163.367
R1066 B.n264 B.n263 163.367
R1067 B.n268 B.n267 163.367
R1068 B.n272 B.n271 163.367
R1069 B.n276 B.n275 163.367
R1070 B.n280 B.n279 163.367
R1071 B.n284 B.n283 163.367
R1072 B.n288 B.n287 163.367
R1073 B.n292 B.n291 163.367
R1074 B.n296 B.n295 163.367
R1075 B.n300 B.n299 163.367
R1076 B.n304 B.n303 163.367
R1077 B.n308 B.n307 163.367
R1078 B.n312 B.n311 163.367
R1079 B.n316 B.n315 163.367
R1080 B.n320 B.n319 163.367
R1081 B.n324 B.n323 163.367
R1082 B.n328 B.n327 163.367
R1083 B.n332 B.n331 163.367
R1084 B.n336 B.n335 163.367
R1085 B.n340 B.n339 163.367
R1086 B.n344 B.n343 163.367
R1087 B.n348 B.n347 163.367
R1088 B.n352 B.n351 163.367
R1089 B.n356 B.n355 163.367
R1090 B.n360 B.n359 163.367
R1091 B.n364 B.n363 163.367
R1092 B.n368 B.n367 163.367
R1093 B.n372 B.n371 163.367
R1094 B.n376 B.n375 163.367
R1095 B.n380 B.n379 163.367
R1096 B.n384 B.n383 163.367
R1097 B.n388 B.n387 163.367
R1098 B.n392 B.n391 163.367
R1099 B.n396 B.n395 163.367
R1100 B.n400 B.n399 163.367
R1101 B.n404 B.n403 163.367
R1102 B.n408 B.n407 163.367
R1103 B.n410 B.n152 163.367
R1104 B.n833 B.n832 71.676
R1105 B.n570 B.n506 71.676
R1106 B.n825 B.n507 71.676
R1107 B.n821 B.n508 71.676
R1108 B.n817 B.n509 71.676
R1109 B.n813 B.n510 71.676
R1110 B.n809 B.n511 71.676
R1111 B.n805 B.n512 71.676
R1112 B.n801 B.n513 71.676
R1113 B.n797 B.n514 71.676
R1114 B.n793 B.n515 71.676
R1115 B.n789 B.n516 71.676
R1116 B.n785 B.n517 71.676
R1117 B.n781 B.n518 71.676
R1118 B.n777 B.n519 71.676
R1119 B.n773 B.n520 71.676
R1120 B.n769 B.n521 71.676
R1121 B.n765 B.n522 71.676
R1122 B.n761 B.n523 71.676
R1123 B.n757 B.n524 71.676
R1124 B.n753 B.n525 71.676
R1125 B.n749 B.n526 71.676
R1126 B.n745 B.n527 71.676
R1127 B.n741 B.n528 71.676
R1128 B.n737 B.n529 71.676
R1129 B.n733 B.n530 71.676
R1130 B.n729 B.n531 71.676
R1131 B.n725 B.n532 71.676
R1132 B.n721 B.n533 71.676
R1133 B.n717 B.n534 71.676
R1134 B.n712 B.n535 71.676
R1135 B.n708 B.n536 71.676
R1136 B.n704 B.n537 71.676
R1137 B.n700 B.n538 71.676
R1138 B.n696 B.n539 71.676
R1139 B.n691 B.n540 71.676
R1140 B.n687 B.n541 71.676
R1141 B.n683 B.n542 71.676
R1142 B.n679 B.n543 71.676
R1143 B.n675 B.n544 71.676
R1144 B.n671 B.n545 71.676
R1145 B.n667 B.n546 71.676
R1146 B.n663 B.n547 71.676
R1147 B.n659 B.n548 71.676
R1148 B.n655 B.n549 71.676
R1149 B.n651 B.n550 71.676
R1150 B.n647 B.n551 71.676
R1151 B.n643 B.n552 71.676
R1152 B.n639 B.n553 71.676
R1153 B.n635 B.n554 71.676
R1154 B.n631 B.n555 71.676
R1155 B.n627 B.n556 71.676
R1156 B.n623 B.n557 71.676
R1157 B.n619 B.n558 71.676
R1158 B.n615 B.n559 71.676
R1159 B.n611 B.n560 71.676
R1160 B.n607 B.n561 71.676
R1161 B.n603 B.n562 71.676
R1162 B.n599 B.n563 71.676
R1163 B.n595 B.n564 71.676
R1164 B.n591 B.n565 71.676
R1165 B.n587 B.n566 71.676
R1166 B.n583 B.n567 71.676
R1167 B.n579 B.n568 71.676
R1168 B.n1040 B.n1039 71.676
R1169 B.n160 B.n89 71.676
R1170 B.n164 B.n90 71.676
R1171 B.n168 B.n91 71.676
R1172 B.n172 B.n92 71.676
R1173 B.n176 B.n93 71.676
R1174 B.n180 B.n94 71.676
R1175 B.n184 B.n95 71.676
R1176 B.n188 B.n96 71.676
R1177 B.n192 B.n97 71.676
R1178 B.n196 B.n98 71.676
R1179 B.n200 B.n99 71.676
R1180 B.n204 B.n100 71.676
R1181 B.n208 B.n101 71.676
R1182 B.n212 B.n102 71.676
R1183 B.n216 B.n103 71.676
R1184 B.n220 B.n104 71.676
R1185 B.n224 B.n105 71.676
R1186 B.n228 B.n106 71.676
R1187 B.n232 B.n107 71.676
R1188 B.n236 B.n108 71.676
R1189 B.n240 B.n109 71.676
R1190 B.n244 B.n110 71.676
R1191 B.n248 B.n111 71.676
R1192 B.n252 B.n112 71.676
R1193 B.n256 B.n113 71.676
R1194 B.n260 B.n114 71.676
R1195 B.n264 B.n115 71.676
R1196 B.n268 B.n116 71.676
R1197 B.n272 B.n117 71.676
R1198 B.n276 B.n118 71.676
R1199 B.n280 B.n119 71.676
R1200 B.n284 B.n120 71.676
R1201 B.n288 B.n121 71.676
R1202 B.n292 B.n122 71.676
R1203 B.n296 B.n123 71.676
R1204 B.n300 B.n124 71.676
R1205 B.n304 B.n125 71.676
R1206 B.n308 B.n126 71.676
R1207 B.n312 B.n127 71.676
R1208 B.n316 B.n128 71.676
R1209 B.n320 B.n129 71.676
R1210 B.n324 B.n130 71.676
R1211 B.n328 B.n131 71.676
R1212 B.n332 B.n132 71.676
R1213 B.n336 B.n133 71.676
R1214 B.n340 B.n134 71.676
R1215 B.n344 B.n135 71.676
R1216 B.n348 B.n136 71.676
R1217 B.n352 B.n137 71.676
R1218 B.n356 B.n138 71.676
R1219 B.n360 B.n139 71.676
R1220 B.n364 B.n140 71.676
R1221 B.n368 B.n141 71.676
R1222 B.n372 B.n142 71.676
R1223 B.n376 B.n143 71.676
R1224 B.n380 B.n144 71.676
R1225 B.n384 B.n145 71.676
R1226 B.n388 B.n146 71.676
R1227 B.n392 B.n147 71.676
R1228 B.n396 B.n148 71.676
R1229 B.n400 B.n149 71.676
R1230 B.n404 B.n150 71.676
R1231 B.n408 B.n151 71.676
R1232 B.n1037 B.n152 71.676
R1233 B.n1037 B.n1036 71.676
R1234 B.n410 B.n151 71.676
R1235 B.n407 B.n150 71.676
R1236 B.n403 B.n149 71.676
R1237 B.n399 B.n148 71.676
R1238 B.n395 B.n147 71.676
R1239 B.n391 B.n146 71.676
R1240 B.n387 B.n145 71.676
R1241 B.n383 B.n144 71.676
R1242 B.n379 B.n143 71.676
R1243 B.n375 B.n142 71.676
R1244 B.n371 B.n141 71.676
R1245 B.n367 B.n140 71.676
R1246 B.n363 B.n139 71.676
R1247 B.n359 B.n138 71.676
R1248 B.n355 B.n137 71.676
R1249 B.n351 B.n136 71.676
R1250 B.n347 B.n135 71.676
R1251 B.n343 B.n134 71.676
R1252 B.n339 B.n133 71.676
R1253 B.n335 B.n132 71.676
R1254 B.n331 B.n131 71.676
R1255 B.n327 B.n130 71.676
R1256 B.n323 B.n129 71.676
R1257 B.n319 B.n128 71.676
R1258 B.n315 B.n127 71.676
R1259 B.n311 B.n126 71.676
R1260 B.n307 B.n125 71.676
R1261 B.n303 B.n124 71.676
R1262 B.n299 B.n123 71.676
R1263 B.n295 B.n122 71.676
R1264 B.n291 B.n121 71.676
R1265 B.n287 B.n120 71.676
R1266 B.n283 B.n119 71.676
R1267 B.n279 B.n118 71.676
R1268 B.n275 B.n117 71.676
R1269 B.n271 B.n116 71.676
R1270 B.n267 B.n115 71.676
R1271 B.n263 B.n114 71.676
R1272 B.n259 B.n113 71.676
R1273 B.n255 B.n112 71.676
R1274 B.n251 B.n111 71.676
R1275 B.n247 B.n110 71.676
R1276 B.n243 B.n109 71.676
R1277 B.n239 B.n108 71.676
R1278 B.n235 B.n107 71.676
R1279 B.n231 B.n106 71.676
R1280 B.n227 B.n105 71.676
R1281 B.n223 B.n104 71.676
R1282 B.n219 B.n103 71.676
R1283 B.n215 B.n102 71.676
R1284 B.n211 B.n101 71.676
R1285 B.n207 B.n100 71.676
R1286 B.n203 B.n99 71.676
R1287 B.n199 B.n98 71.676
R1288 B.n195 B.n97 71.676
R1289 B.n191 B.n96 71.676
R1290 B.n187 B.n95 71.676
R1291 B.n183 B.n94 71.676
R1292 B.n179 B.n93 71.676
R1293 B.n175 B.n92 71.676
R1294 B.n171 B.n91 71.676
R1295 B.n167 B.n90 71.676
R1296 B.n163 B.n89 71.676
R1297 B.n1039 B.n88 71.676
R1298 B.n832 B.n505 71.676
R1299 B.n826 B.n506 71.676
R1300 B.n822 B.n507 71.676
R1301 B.n818 B.n508 71.676
R1302 B.n814 B.n509 71.676
R1303 B.n810 B.n510 71.676
R1304 B.n806 B.n511 71.676
R1305 B.n802 B.n512 71.676
R1306 B.n798 B.n513 71.676
R1307 B.n794 B.n514 71.676
R1308 B.n790 B.n515 71.676
R1309 B.n786 B.n516 71.676
R1310 B.n782 B.n517 71.676
R1311 B.n778 B.n518 71.676
R1312 B.n774 B.n519 71.676
R1313 B.n770 B.n520 71.676
R1314 B.n766 B.n521 71.676
R1315 B.n762 B.n522 71.676
R1316 B.n758 B.n523 71.676
R1317 B.n754 B.n524 71.676
R1318 B.n750 B.n525 71.676
R1319 B.n746 B.n526 71.676
R1320 B.n742 B.n527 71.676
R1321 B.n738 B.n528 71.676
R1322 B.n734 B.n529 71.676
R1323 B.n730 B.n530 71.676
R1324 B.n726 B.n531 71.676
R1325 B.n722 B.n532 71.676
R1326 B.n718 B.n533 71.676
R1327 B.n713 B.n534 71.676
R1328 B.n709 B.n535 71.676
R1329 B.n705 B.n536 71.676
R1330 B.n701 B.n537 71.676
R1331 B.n697 B.n538 71.676
R1332 B.n692 B.n539 71.676
R1333 B.n688 B.n540 71.676
R1334 B.n684 B.n541 71.676
R1335 B.n680 B.n542 71.676
R1336 B.n676 B.n543 71.676
R1337 B.n672 B.n544 71.676
R1338 B.n668 B.n545 71.676
R1339 B.n664 B.n546 71.676
R1340 B.n660 B.n547 71.676
R1341 B.n656 B.n548 71.676
R1342 B.n652 B.n549 71.676
R1343 B.n648 B.n550 71.676
R1344 B.n644 B.n551 71.676
R1345 B.n640 B.n552 71.676
R1346 B.n636 B.n553 71.676
R1347 B.n632 B.n554 71.676
R1348 B.n628 B.n555 71.676
R1349 B.n624 B.n556 71.676
R1350 B.n620 B.n557 71.676
R1351 B.n616 B.n558 71.676
R1352 B.n612 B.n559 71.676
R1353 B.n608 B.n560 71.676
R1354 B.n604 B.n561 71.676
R1355 B.n600 B.n562 71.676
R1356 B.n596 B.n563 71.676
R1357 B.n592 B.n564 71.676
R1358 B.n588 B.n565 71.676
R1359 B.n584 B.n566 71.676
R1360 B.n580 B.n567 71.676
R1361 B.n576 B.n568 71.676
R1362 B.n694 B.n574 59.5399
R1363 B.n715 B.n572 59.5399
R1364 B.n159 B.n158 59.5399
R1365 B.n156 B.n155 59.5399
R1366 B.n831 B.n502 55.6671
R1367 B.n1038 B.n85 55.6671
R1368 B.n574 B.n573 42.6672
R1369 B.n572 B.n571 42.6672
R1370 B.n158 B.n157 42.6672
R1371 B.n155 B.n154 42.6672
R1372 B.n838 B.n502 31.81
R1373 B.n838 B.n498 31.81
R1374 B.n844 B.n498 31.81
R1375 B.n844 B.n493 31.81
R1376 B.n850 B.n493 31.81
R1377 B.n850 B.n494 31.81
R1378 B.n856 B.n486 31.81
R1379 B.n862 B.n486 31.81
R1380 B.n862 B.n482 31.81
R1381 B.n868 B.n482 31.81
R1382 B.n868 B.n478 31.81
R1383 B.n874 B.n478 31.81
R1384 B.n874 B.n474 31.81
R1385 B.n881 B.n474 31.81
R1386 B.n881 B.n880 31.81
R1387 B.n887 B.n467 31.81
R1388 B.n893 B.n467 31.81
R1389 B.n893 B.n462 31.81
R1390 B.n899 B.n462 31.81
R1391 B.n899 B.n463 31.81
R1392 B.n905 B.n455 31.81
R1393 B.n911 B.n455 31.81
R1394 B.n911 B.n451 31.81
R1395 B.n917 B.n451 31.81
R1396 B.n917 B.n447 31.81
R1397 B.n923 B.n447 31.81
R1398 B.n929 B.n443 31.81
R1399 B.n929 B.n439 31.81
R1400 B.n935 B.n439 31.81
R1401 B.n935 B.n435 31.81
R1402 B.n941 B.n435 31.81
R1403 B.n947 B.n431 31.81
R1404 B.n947 B.n427 31.81
R1405 B.n953 B.n427 31.81
R1406 B.n953 B.n422 31.81
R1407 B.n959 B.n422 31.81
R1408 B.n959 B.n423 31.81
R1409 B.n966 B.n415 31.81
R1410 B.n972 B.n415 31.81
R1411 B.n972 B.n4 31.81
R1412 B.n1135 B.n4 31.81
R1413 B.n1135 B.n1134 31.81
R1414 B.n1134 B.n1133 31.81
R1415 B.n1133 B.n8 31.81
R1416 B.n1127 B.n8 31.81
R1417 B.n1126 B.n1125 31.81
R1418 B.n1125 B.n15 31.81
R1419 B.n1119 B.n15 31.81
R1420 B.n1119 B.n1118 31.81
R1421 B.n1118 B.n1117 31.81
R1422 B.n1117 B.n22 31.81
R1423 B.n1111 B.n1110 31.81
R1424 B.n1110 B.n1109 31.81
R1425 B.n1109 B.n29 31.81
R1426 B.n1103 B.n29 31.81
R1427 B.n1103 B.n1102 31.81
R1428 B.n1101 B.n36 31.81
R1429 B.n1095 B.n36 31.81
R1430 B.n1095 B.n1094 31.81
R1431 B.n1094 B.n1093 31.81
R1432 B.n1093 B.n43 31.81
R1433 B.n1087 B.n43 31.81
R1434 B.n1086 B.n1085 31.81
R1435 B.n1085 B.n50 31.81
R1436 B.n1079 B.n50 31.81
R1437 B.n1079 B.n1078 31.81
R1438 B.n1078 B.n1077 31.81
R1439 B.n1071 B.n60 31.81
R1440 B.n1071 B.n1070 31.81
R1441 B.n1070 B.n1069 31.81
R1442 B.n1069 B.n64 31.81
R1443 B.n1063 B.n64 31.81
R1444 B.n1063 B.n1062 31.81
R1445 B.n1062 B.n1061 31.81
R1446 B.n1061 B.n71 31.81
R1447 B.n1055 B.n71 31.81
R1448 B.n1054 B.n1053 31.81
R1449 B.n1053 B.n78 31.81
R1450 B.n1047 B.n78 31.81
R1451 B.n1047 B.n1046 31.81
R1452 B.n1046 B.n1045 31.81
R1453 B.n1045 B.n85 31.81
R1454 B.n1035 B.n1034 29.1907
R1455 B.n1042 B.n1041 29.1907
R1456 B.n575 B.n500 29.1907
R1457 B.n835 B.n834 29.1907
R1458 B.n966 B.t7 26.6643
R1459 B.n1127 B.t6 26.6643
R1460 B.t4 B.n443 24.7932
R1461 B.n1102 B.t2 24.7932
R1462 B.n463 B.t0 23.8576
R1463 B.t1 B.n1086 23.8576
R1464 B.n887 B.t5 22.922
R1465 B.n1077 B.t8 22.922
R1466 B.n941 B.t9 21.9865
R1467 B.n1111 B.t3 21.9865
R1468 B.n494 B.t11 19.1797
R1469 B.t18 B.n1054 19.1797
R1470 B B.n1137 18.0485
R1471 B.n856 B.t11 12.6307
R1472 B.n1055 B.t18 12.6307
R1473 B.n1041 B.n87 10.6151
R1474 B.n161 B.n87 10.6151
R1475 B.n162 B.n161 10.6151
R1476 B.n165 B.n162 10.6151
R1477 B.n166 B.n165 10.6151
R1478 B.n169 B.n166 10.6151
R1479 B.n170 B.n169 10.6151
R1480 B.n173 B.n170 10.6151
R1481 B.n174 B.n173 10.6151
R1482 B.n177 B.n174 10.6151
R1483 B.n178 B.n177 10.6151
R1484 B.n181 B.n178 10.6151
R1485 B.n182 B.n181 10.6151
R1486 B.n185 B.n182 10.6151
R1487 B.n186 B.n185 10.6151
R1488 B.n189 B.n186 10.6151
R1489 B.n190 B.n189 10.6151
R1490 B.n193 B.n190 10.6151
R1491 B.n194 B.n193 10.6151
R1492 B.n197 B.n194 10.6151
R1493 B.n198 B.n197 10.6151
R1494 B.n201 B.n198 10.6151
R1495 B.n202 B.n201 10.6151
R1496 B.n205 B.n202 10.6151
R1497 B.n206 B.n205 10.6151
R1498 B.n209 B.n206 10.6151
R1499 B.n210 B.n209 10.6151
R1500 B.n213 B.n210 10.6151
R1501 B.n214 B.n213 10.6151
R1502 B.n217 B.n214 10.6151
R1503 B.n218 B.n217 10.6151
R1504 B.n221 B.n218 10.6151
R1505 B.n222 B.n221 10.6151
R1506 B.n225 B.n222 10.6151
R1507 B.n226 B.n225 10.6151
R1508 B.n229 B.n226 10.6151
R1509 B.n230 B.n229 10.6151
R1510 B.n233 B.n230 10.6151
R1511 B.n234 B.n233 10.6151
R1512 B.n237 B.n234 10.6151
R1513 B.n238 B.n237 10.6151
R1514 B.n241 B.n238 10.6151
R1515 B.n242 B.n241 10.6151
R1516 B.n245 B.n242 10.6151
R1517 B.n246 B.n245 10.6151
R1518 B.n249 B.n246 10.6151
R1519 B.n250 B.n249 10.6151
R1520 B.n253 B.n250 10.6151
R1521 B.n254 B.n253 10.6151
R1522 B.n257 B.n254 10.6151
R1523 B.n258 B.n257 10.6151
R1524 B.n261 B.n258 10.6151
R1525 B.n262 B.n261 10.6151
R1526 B.n265 B.n262 10.6151
R1527 B.n266 B.n265 10.6151
R1528 B.n269 B.n266 10.6151
R1529 B.n270 B.n269 10.6151
R1530 B.n273 B.n270 10.6151
R1531 B.n274 B.n273 10.6151
R1532 B.n278 B.n277 10.6151
R1533 B.n281 B.n278 10.6151
R1534 B.n282 B.n281 10.6151
R1535 B.n285 B.n282 10.6151
R1536 B.n286 B.n285 10.6151
R1537 B.n289 B.n286 10.6151
R1538 B.n290 B.n289 10.6151
R1539 B.n293 B.n290 10.6151
R1540 B.n294 B.n293 10.6151
R1541 B.n298 B.n297 10.6151
R1542 B.n301 B.n298 10.6151
R1543 B.n302 B.n301 10.6151
R1544 B.n305 B.n302 10.6151
R1545 B.n306 B.n305 10.6151
R1546 B.n309 B.n306 10.6151
R1547 B.n310 B.n309 10.6151
R1548 B.n313 B.n310 10.6151
R1549 B.n314 B.n313 10.6151
R1550 B.n317 B.n314 10.6151
R1551 B.n318 B.n317 10.6151
R1552 B.n321 B.n318 10.6151
R1553 B.n322 B.n321 10.6151
R1554 B.n325 B.n322 10.6151
R1555 B.n326 B.n325 10.6151
R1556 B.n329 B.n326 10.6151
R1557 B.n330 B.n329 10.6151
R1558 B.n333 B.n330 10.6151
R1559 B.n334 B.n333 10.6151
R1560 B.n337 B.n334 10.6151
R1561 B.n338 B.n337 10.6151
R1562 B.n341 B.n338 10.6151
R1563 B.n342 B.n341 10.6151
R1564 B.n345 B.n342 10.6151
R1565 B.n346 B.n345 10.6151
R1566 B.n349 B.n346 10.6151
R1567 B.n350 B.n349 10.6151
R1568 B.n353 B.n350 10.6151
R1569 B.n354 B.n353 10.6151
R1570 B.n357 B.n354 10.6151
R1571 B.n358 B.n357 10.6151
R1572 B.n361 B.n358 10.6151
R1573 B.n362 B.n361 10.6151
R1574 B.n365 B.n362 10.6151
R1575 B.n366 B.n365 10.6151
R1576 B.n369 B.n366 10.6151
R1577 B.n370 B.n369 10.6151
R1578 B.n373 B.n370 10.6151
R1579 B.n374 B.n373 10.6151
R1580 B.n377 B.n374 10.6151
R1581 B.n378 B.n377 10.6151
R1582 B.n381 B.n378 10.6151
R1583 B.n382 B.n381 10.6151
R1584 B.n385 B.n382 10.6151
R1585 B.n386 B.n385 10.6151
R1586 B.n389 B.n386 10.6151
R1587 B.n390 B.n389 10.6151
R1588 B.n393 B.n390 10.6151
R1589 B.n394 B.n393 10.6151
R1590 B.n397 B.n394 10.6151
R1591 B.n398 B.n397 10.6151
R1592 B.n401 B.n398 10.6151
R1593 B.n402 B.n401 10.6151
R1594 B.n405 B.n402 10.6151
R1595 B.n406 B.n405 10.6151
R1596 B.n409 B.n406 10.6151
R1597 B.n411 B.n409 10.6151
R1598 B.n412 B.n411 10.6151
R1599 B.n1035 B.n412 10.6151
R1600 B.n840 B.n500 10.6151
R1601 B.n841 B.n840 10.6151
R1602 B.n842 B.n841 10.6151
R1603 B.n842 B.n491 10.6151
R1604 B.n852 B.n491 10.6151
R1605 B.n853 B.n852 10.6151
R1606 B.n854 B.n853 10.6151
R1607 B.n854 B.n484 10.6151
R1608 B.n864 B.n484 10.6151
R1609 B.n865 B.n864 10.6151
R1610 B.n866 B.n865 10.6151
R1611 B.n866 B.n476 10.6151
R1612 B.n876 B.n476 10.6151
R1613 B.n877 B.n876 10.6151
R1614 B.n878 B.n877 10.6151
R1615 B.n878 B.n469 10.6151
R1616 B.n889 B.n469 10.6151
R1617 B.n890 B.n889 10.6151
R1618 B.n891 B.n890 10.6151
R1619 B.n891 B.n460 10.6151
R1620 B.n901 B.n460 10.6151
R1621 B.n902 B.n901 10.6151
R1622 B.n903 B.n902 10.6151
R1623 B.n903 B.n453 10.6151
R1624 B.n913 B.n453 10.6151
R1625 B.n914 B.n913 10.6151
R1626 B.n915 B.n914 10.6151
R1627 B.n915 B.n445 10.6151
R1628 B.n925 B.n445 10.6151
R1629 B.n926 B.n925 10.6151
R1630 B.n927 B.n926 10.6151
R1631 B.n927 B.n437 10.6151
R1632 B.n937 B.n437 10.6151
R1633 B.n938 B.n937 10.6151
R1634 B.n939 B.n938 10.6151
R1635 B.n939 B.n429 10.6151
R1636 B.n949 B.n429 10.6151
R1637 B.n950 B.n949 10.6151
R1638 B.n951 B.n950 10.6151
R1639 B.n951 B.n420 10.6151
R1640 B.n961 B.n420 10.6151
R1641 B.n962 B.n961 10.6151
R1642 B.n964 B.n962 10.6151
R1643 B.n964 B.n963 10.6151
R1644 B.n963 B.n413 10.6151
R1645 B.n975 B.n413 10.6151
R1646 B.n976 B.n975 10.6151
R1647 B.n977 B.n976 10.6151
R1648 B.n978 B.n977 10.6151
R1649 B.n980 B.n978 10.6151
R1650 B.n981 B.n980 10.6151
R1651 B.n982 B.n981 10.6151
R1652 B.n983 B.n982 10.6151
R1653 B.n985 B.n983 10.6151
R1654 B.n986 B.n985 10.6151
R1655 B.n987 B.n986 10.6151
R1656 B.n988 B.n987 10.6151
R1657 B.n990 B.n988 10.6151
R1658 B.n991 B.n990 10.6151
R1659 B.n992 B.n991 10.6151
R1660 B.n993 B.n992 10.6151
R1661 B.n995 B.n993 10.6151
R1662 B.n996 B.n995 10.6151
R1663 B.n997 B.n996 10.6151
R1664 B.n998 B.n997 10.6151
R1665 B.n1000 B.n998 10.6151
R1666 B.n1001 B.n1000 10.6151
R1667 B.n1002 B.n1001 10.6151
R1668 B.n1003 B.n1002 10.6151
R1669 B.n1005 B.n1003 10.6151
R1670 B.n1006 B.n1005 10.6151
R1671 B.n1007 B.n1006 10.6151
R1672 B.n1008 B.n1007 10.6151
R1673 B.n1010 B.n1008 10.6151
R1674 B.n1011 B.n1010 10.6151
R1675 B.n1012 B.n1011 10.6151
R1676 B.n1013 B.n1012 10.6151
R1677 B.n1015 B.n1013 10.6151
R1678 B.n1016 B.n1015 10.6151
R1679 B.n1017 B.n1016 10.6151
R1680 B.n1018 B.n1017 10.6151
R1681 B.n1020 B.n1018 10.6151
R1682 B.n1021 B.n1020 10.6151
R1683 B.n1022 B.n1021 10.6151
R1684 B.n1023 B.n1022 10.6151
R1685 B.n1025 B.n1023 10.6151
R1686 B.n1026 B.n1025 10.6151
R1687 B.n1027 B.n1026 10.6151
R1688 B.n1028 B.n1027 10.6151
R1689 B.n1030 B.n1028 10.6151
R1690 B.n1031 B.n1030 10.6151
R1691 B.n1032 B.n1031 10.6151
R1692 B.n1033 B.n1032 10.6151
R1693 B.n1034 B.n1033 10.6151
R1694 B.n834 B.n504 10.6151
R1695 B.n829 B.n504 10.6151
R1696 B.n829 B.n828 10.6151
R1697 B.n828 B.n827 10.6151
R1698 B.n827 B.n824 10.6151
R1699 B.n824 B.n823 10.6151
R1700 B.n823 B.n820 10.6151
R1701 B.n820 B.n819 10.6151
R1702 B.n819 B.n816 10.6151
R1703 B.n816 B.n815 10.6151
R1704 B.n815 B.n812 10.6151
R1705 B.n812 B.n811 10.6151
R1706 B.n811 B.n808 10.6151
R1707 B.n808 B.n807 10.6151
R1708 B.n807 B.n804 10.6151
R1709 B.n804 B.n803 10.6151
R1710 B.n803 B.n800 10.6151
R1711 B.n800 B.n799 10.6151
R1712 B.n799 B.n796 10.6151
R1713 B.n796 B.n795 10.6151
R1714 B.n795 B.n792 10.6151
R1715 B.n792 B.n791 10.6151
R1716 B.n791 B.n788 10.6151
R1717 B.n788 B.n787 10.6151
R1718 B.n787 B.n784 10.6151
R1719 B.n784 B.n783 10.6151
R1720 B.n783 B.n780 10.6151
R1721 B.n780 B.n779 10.6151
R1722 B.n779 B.n776 10.6151
R1723 B.n776 B.n775 10.6151
R1724 B.n775 B.n772 10.6151
R1725 B.n772 B.n771 10.6151
R1726 B.n771 B.n768 10.6151
R1727 B.n768 B.n767 10.6151
R1728 B.n767 B.n764 10.6151
R1729 B.n764 B.n763 10.6151
R1730 B.n763 B.n760 10.6151
R1731 B.n760 B.n759 10.6151
R1732 B.n759 B.n756 10.6151
R1733 B.n756 B.n755 10.6151
R1734 B.n755 B.n752 10.6151
R1735 B.n752 B.n751 10.6151
R1736 B.n751 B.n748 10.6151
R1737 B.n748 B.n747 10.6151
R1738 B.n747 B.n744 10.6151
R1739 B.n744 B.n743 10.6151
R1740 B.n743 B.n740 10.6151
R1741 B.n740 B.n739 10.6151
R1742 B.n739 B.n736 10.6151
R1743 B.n736 B.n735 10.6151
R1744 B.n735 B.n732 10.6151
R1745 B.n732 B.n731 10.6151
R1746 B.n731 B.n728 10.6151
R1747 B.n728 B.n727 10.6151
R1748 B.n727 B.n724 10.6151
R1749 B.n724 B.n723 10.6151
R1750 B.n723 B.n720 10.6151
R1751 B.n720 B.n719 10.6151
R1752 B.n719 B.n716 10.6151
R1753 B.n714 B.n711 10.6151
R1754 B.n711 B.n710 10.6151
R1755 B.n710 B.n707 10.6151
R1756 B.n707 B.n706 10.6151
R1757 B.n706 B.n703 10.6151
R1758 B.n703 B.n702 10.6151
R1759 B.n702 B.n699 10.6151
R1760 B.n699 B.n698 10.6151
R1761 B.n698 B.n695 10.6151
R1762 B.n693 B.n690 10.6151
R1763 B.n690 B.n689 10.6151
R1764 B.n689 B.n686 10.6151
R1765 B.n686 B.n685 10.6151
R1766 B.n685 B.n682 10.6151
R1767 B.n682 B.n681 10.6151
R1768 B.n681 B.n678 10.6151
R1769 B.n678 B.n677 10.6151
R1770 B.n677 B.n674 10.6151
R1771 B.n674 B.n673 10.6151
R1772 B.n673 B.n670 10.6151
R1773 B.n670 B.n669 10.6151
R1774 B.n669 B.n666 10.6151
R1775 B.n666 B.n665 10.6151
R1776 B.n665 B.n662 10.6151
R1777 B.n662 B.n661 10.6151
R1778 B.n661 B.n658 10.6151
R1779 B.n658 B.n657 10.6151
R1780 B.n657 B.n654 10.6151
R1781 B.n654 B.n653 10.6151
R1782 B.n653 B.n650 10.6151
R1783 B.n650 B.n649 10.6151
R1784 B.n649 B.n646 10.6151
R1785 B.n646 B.n645 10.6151
R1786 B.n645 B.n642 10.6151
R1787 B.n642 B.n641 10.6151
R1788 B.n641 B.n638 10.6151
R1789 B.n638 B.n637 10.6151
R1790 B.n637 B.n634 10.6151
R1791 B.n634 B.n633 10.6151
R1792 B.n633 B.n630 10.6151
R1793 B.n630 B.n629 10.6151
R1794 B.n629 B.n626 10.6151
R1795 B.n626 B.n625 10.6151
R1796 B.n625 B.n622 10.6151
R1797 B.n622 B.n621 10.6151
R1798 B.n621 B.n618 10.6151
R1799 B.n618 B.n617 10.6151
R1800 B.n617 B.n614 10.6151
R1801 B.n614 B.n613 10.6151
R1802 B.n613 B.n610 10.6151
R1803 B.n610 B.n609 10.6151
R1804 B.n609 B.n606 10.6151
R1805 B.n606 B.n605 10.6151
R1806 B.n605 B.n602 10.6151
R1807 B.n602 B.n601 10.6151
R1808 B.n601 B.n598 10.6151
R1809 B.n598 B.n597 10.6151
R1810 B.n597 B.n594 10.6151
R1811 B.n594 B.n593 10.6151
R1812 B.n593 B.n590 10.6151
R1813 B.n590 B.n589 10.6151
R1814 B.n589 B.n586 10.6151
R1815 B.n586 B.n585 10.6151
R1816 B.n585 B.n582 10.6151
R1817 B.n582 B.n581 10.6151
R1818 B.n581 B.n578 10.6151
R1819 B.n578 B.n577 10.6151
R1820 B.n577 B.n575 10.6151
R1821 B.n836 B.n835 10.6151
R1822 B.n836 B.n496 10.6151
R1823 B.n846 B.n496 10.6151
R1824 B.n847 B.n846 10.6151
R1825 B.n848 B.n847 10.6151
R1826 B.n848 B.n488 10.6151
R1827 B.n858 B.n488 10.6151
R1828 B.n859 B.n858 10.6151
R1829 B.n860 B.n859 10.6151
R1830 B.n860 B.n480 10.6151
R1831 B.n870 B.n480 10.6151
R1832 B.n871 B.n870 10.6151
R1833 B.n872 B.n871 10.6151
R1834 B.n872 B.n472 10.6151
R1835 B.n883 B.n472 10.6151
R1836 B.n884 B.n883 10.6151
R1837 B.n885 B.n884 10.6151
R1838 B.n885 B.n465 10.6151
R1839 B.n895 B.n465 10.6151
R1840 B.n896 B.n895 10.6151
R1841 B.n897 B.n896 10.6151
R1842 B.n897 B.n457 10.6151
R1843 B.n907 B.n457 10.6151
R1844 B.n908 B.n907 10.6151
R1845 B.n909 B.n908 10.6151
R1846 B.n909 B.n449 10.6151
R1847 B.n919 B.n449 10.6151
R1848 B.n920 B.n919 10.6151
R1849 B.n921 B.n920 10.6151
R1850 B.n921 B.n441 10.6151
R1851 B.n931 B.n441 10.6151
R1852 B.n932 B.n931 10.6151
R1853 B.n933 B.n932 10.6151
R1854 B.n933 B.n433 10.6151
R1855 B.n943 B.n433 10.6151
R1856 B.n944 B.n943 10.6151
R1857 B.n945 B.n944 10.6151
R1858 B.n945 B.n425 10.6151
R1859 B.n955 B.n425 10.6151
R1860 B.n956 B.n955 10.6151
R1861 B.n957 B.n956 10.6151
R1862 B.n957 B.n417 10.6151
R1863 B.n968 B.n417 10.6151
R1864 B.n969 B.n968 10.6151
R1865 B.n970 B.n969 10.6151
R1866 B.n970 B.n0 10.6151
R1867 B.n1131 B.n1 10.6151
R1868 B.n1131 B.n1130 10.6151
R1869 B.n1130 B.n1129 10.6151
R1870 B.n1129 B.n10 10.6151
R1871 B.n1123 B.n10 10.6151
R1872 B.n1123 B.n1122 10.6151
R1873 B.n1122 B.n1121 10.6151
R1874 B.n1121 B.n17 10.6151
R1875 B.n1115 B.n17 10.6151
R1876 B.n1115 B.n1114 10.6151
R1877 B.n1114 B.n1113 10.6151
R1878 B.n1113 B.n24 10.6151
R1879 B.n1107 B.n24 10.6151
R1880 B.n1107 B.n1106 10.6151
R1881 B.n1106 B.n1105 10.6151
R1882 B.n1105 B.n31 10.6151
R1883 B.n1099 B.n31 10.6151
R1884 B.n1099 B.n1098 10.6151
R1885 B.n1098 B.n1097 10.6151
R1886 B.n1097 B.n38 10.6151
R1887 B.n1091 B.n38 10.6151
R1888 B.n1091 B.n1090 10.6151
R1889 B.n1090 B.n1089 10.6151
R1890 B.n1089 B.n45 10.6151
R1891 B.n1083 B.n45 10.6151
R1892 B.n1083 B.n1082 10.6151
R1893 B.n1082 B.n1081 10.6151
R1894 B.n1081 B.n52 10.6151
R1895 B.n1075 B.n52 10.6151
R1896 B.n1075 B.n1074 10.6151
R1897 B.n1074 B.n1073 10.6151
R1898 B.n1073 B.n58 10.6151
R1899 B.n1067 B.n58 10.6151
R1900 B.n1067 B.n1066 10.6151
R1901 B.n1066 B.n1065 10.6151
R1902 B.n1065 B.n66 10.6151
R1903 B.n1059 B.n66 10.6151
R1904 B.n1059 B.n1058 10.6151
R1905 B.n1058 B.n1057 10.6151
R1906 B.n1057 B.n73 10.6151
R1907 B.n1051 B.n73 10.6151
R1908 B.n1051 B.n1050 10.6151
R1909 B.n1050 B.n1049 10.6151
R1910 B.n1049 B.n80 10.6151
R1911 B.n1043 B.n80 10.6151
R1912 B.n1043 B.n1042 10.6151
R1913 B.t9 B.n431 9.82402
R1914 B.t3 B.n22 9.82402
R1915 B.n274 B.n159 9.36635
R1916 B.n297 B.n156 9.36635
R1917 B.n716 B.n715 9.36635
R1918 B.n694 B.n693 9.36635
R1919 B.n880 B.t5 8.88844
R1920 B.n60 B.t8 8.88844
R1921 B.n905 B.t0 7.95287
R1922 B.n1087 B.t1 7.95287
R1923 B.n923 B.t4 7.0173
R1924 B.t2 B.n1101 7.0173
R1925 B.n423 B.t7 5.14615
R1926 B.t6 B.n1126 5.14615
R1927 B.n1137 B.n0 2.81026
R1928 B.n1137 B.n1 2.81026
R1929 B.n277 B.n159 1.24928
R1930 B.n294 B.n156 1.24928
R1931 B.n715 B.n714 1.24928
R1932 B.n695 B.n694 1.24928
R1933 VN.n7 VN.t1 265.42
R1934 VN.n38 VN.t8 265.42
R1935 VN.n15 VN.t7 235.072
R1936 VN.n8 VN.t9 235.072
R1937 VN.n22 VN.t6 235.072
R1938 VN.n29 VN.t0 235.072
R1939 VN.n46 VN.t5 235.072
R1940 VN.n39 VN.t4 235.072
R1941 VN.n53 VN.t2 235.072
R1942 VN.n60 VN.t3 235.072
R1943 VN.n59 VN.n31 161.3
R1944 VN.n58 VN.n57 161.3
R1945 VN.n56 VN.n32 161.3
R1946 VN.n55 VN.n54 161.3
R1947 VN.n52 VN.n33 161.3
R1948 VN.n51 VN.n50 161.3
R1949 VN.n49 VN.n34 161.3
R1950 VN.n48 VN.n47 161.3
R1951 VN.n46 VN.n35 161.3
R1952 VN.n45 VN.n44 161.3
R1953 VN.n43 VN.n36 161.3
R1954 VN.n42 VN.n41 161.3
R1955 VN.n40 VN.n37 161.3
R1956 VN.n28 VN.n0 161.3
R1957 VN.n27 VN.n26 161.3
R1958 VN.n25 VN.n1 161.3
R1959 VN.n24 VN.n23 161.3
R1960 VN.n21 VN.n2 161.3
R1961 VN.n20 VN.n19 161.3
R1962 VN.n18 VN.n3 161.3
R1963 VN.n17 VN.n16 161.3
R1964 VN.n15 VN.n4 161.3
R1965 VN.n14 VN.n13 161.3
R1966 VN.n12 VN.n5 161.3
R1967 VN.n11 VN.n10 161.3
R1968 VN.n9 VN.n6 161.3
R1969 VN.n30 VN.n29 91.2348
R1970 VN.n61 VN.n60 91.2348
R1971 VN.n8 VN.n7 60.1239
R1972 VN.n39 VN.n38 60.1239
R1973 VN.n27 VN.n1 56.5617
R1974 VN.n58 VN.n32 56.5617
R1975 VN VN.n61 54.1421
R1976 VN.n10 VN.n5 50.2647
R1977 VN.n20 VN.n3 50.2647
R1978 VN.n41 VN.n36 50.2647
R1979 VN.n51 VN.n34 50.2647
R1980 VN.n14 VN.n5 30.8893
R1981 VN.n16 VN.n3 30.8893
R1982 VN.n45 VN.n36 30.8893
R1983 VN.n47 VN.n34 30.8893
R1984 VN.n10 VN.n9 24.5923
R1985 VN.n15 VN.n14 24.5923
R1986 VN.n16 VN.n15 24.5923
R1987 VN.n21 VN.n20 24.5923
R1988 VN.n23 VN.n1 24.5923
R1989 VN.n28 VN.n27 24.5923
R1990 VN.n41 VN.n40 24.5923
R1991 VN.n47 VN.n46 24.5923
R1992 VN.n46 VN.n45 24.5923
R1993 VN.n54 VN.n32 24.5923
R1994 VN.n52 VN.n51 24.5923
R1995 VN.n59 VN.n58 24.5923
R1996 VN.n29 VN.n28 19.674
R1997 VN.n60 VN.n59 19.674
R1998 VN.n23 VN.n22 14.7556
R1999 VN.n54 VN.n53 14.7556
R2000 VN.n38 VN.n37 13.3418
R2001 VN.n7 VN.n6 13.3418
R2002 VN.n9 VN.n8 9.83723
R2003 VN.n22 VN.n21 9.83723
R2004 VN.n40 VN.n39 9.83723
R2005 VN.n53 VN.n52 9.83723
R2006 VN.n61 VN.n31 0.278335
R2007 VN.n30 VN.n0 0.278335
R2008 VN.n57 VN.n31 0.189894
R2009 VN.n57 VN.n56 0.189894
R2010 VN.n56 VN.n55 0.189894
R2011 VN.n55 VN.n33 0.189894
R2012 VN.n50 VN.n33 0.189894
R2013 VN.n50 VN.n49 0.189894
R2014 VN.n49 VN.n48 0.189894
R2015 VN.n48 VN.n35 0.189894
R2016 VN.n44 VN.n35 0.189894
R2017 VN.n44 VN.n43 0.189894
R2018 VN.n43 VN.n42 0.189894
R2019 VN.n42 VN.n37 0.189894
R2020 VN.n11 VN.n6 0.189894
R2021 VN.n12 VN.n11 0.189894
R2022 VN.n13 VN.n12 0.189894
R2023 VN.n13 VN.n4 0.189894
R2024 VN.n17 VN.n4 0.189894
R2025 VN.n18 VN.n17 0.189894
R2026 VN.n19 VN.n18 0.189894
R2027 VN.n19 VN.n2 0.189894
R2028 VN.n24 VN.n2 0.189894
R2029 VN.n25 VN.n24 0.189894
R2030 VN.n26 VN.n25 0.189894
R2031 VN.n26 VN.n0 0.189894
R2032 VN VN.n30 0.153485
R2033 VTAIL.n416 VTAIL.n320 289.615
R2034 VTAIL.n98 VTAIL.n2 289.615
R2035 VTAIL.n314 VTAIL.n218 289.615
R2036 VTAIL.n208 VTAIL.n112 289.615
R2037 VTAIL.n352 VTAIL.n351 185
R2038 VTAIL.n357 VTAIL.n356 185
R2039 VTAIL.n359 VTAIL.n358 185
R2040 VTAIL.n348 VTAIL.n347 185
R2041 VTAIL.n365 VTAIL.n364 185
R2042 VTAIL.n367 VTAIL.n366 185
R2043 VTAIL.n344 VTAIL.n343 185
R2044 VTAIL.n373 VTAIL.n372 185
R2045 VTAIL.n375 VTAIL.n374 185
R2046 VTAIL.n340 VTAIL.n339 185
R2047 VTAIL.n381 VTAIL.n380 185
R2048 VTAIL.n383 VTAIL.n382 185
R2049 VTAIL.n336 VTAIL.n335 185
R2050 VTAIL.n389 VTAIL.n388 185
R2051 VTAIL.n391 VTAIL.n390 185
R2052 VTAIL.n332 VTAIL.n331 185
R2053 VTAIL.n398 VTAIL.n397 185
R2054 VTAIL.n399 VTAIL.n330 185
R2055 VTAIL.n401 VTAIL.n400 185
R2056 VTAIL.n328 VTAIL.n327 185
R2057 VTAIL.n407 VTAIL.n406 185
R2058 VTAIL.n409 VTAIL.n408 185
R2059 VTAIL.n324 VTAIL.n323 185
R2060 VTAIL.n415 VTAIL.n414 185
R2061 VTAIL.n417 VTAIL.n416 185
R2062 VTAIL.n34 VTAIL.n33 185
R2063 VTAIL.n39 VTAIL.n38 185
R2064 VTAIL.n41 VTAIL.n40 185
R2065 VTAIL.n30 VTAIL.n29 185
R2066 VTAIL.n47 VTAIL.n46 185
R2067 VTAIL.n49 VTAIL.n48 185
R2068 VTAIL.n26 VTAIL.n25 185
R2069 VTAIL.n55 VTAIL.n54 185
R2070 VTAIL.n57 VTAIL.n56 185
R2071 VTAIL.n22 VTAIL.n21 185
R2072 VTAIL.n63 VTAIL.n62 185
R2073 VTAIL.n65 VTAIL.n64 185
R2074 VTAIL.n18 VTAIL.n17 185
R2075 VTAIL.n71 VTAIL.n70 185
R2076 VTAIL.n73 VTAIL.n72 185
R2077 VTAIL.n14 VTAIL.n13 185
R2078 VTAIL.n80 VTAIL.n79 185
R2079 VTAIL.n81 VTAIL.n12 185
R2080 VTAIL.n83 VTAIL.n82 185
R2081 VTAIL.n10 VTAIL.n9 185
R2082 VTAIL.n89 VTAIL.n88 185
R2083 VTAIL.n91 VTAIL.n90 185
R2084 VTAIL.n6 VTAIL.n5 185
R2085 VTAIL.n97 VTAIL.n96 185
R2086 VTAIL.n99 VTAIL.n98 185
R2087 VTAIL.n315 VTAIL.n314 185
R2088 VTAIL.n313 VTAIL.n312 185
R2089 VTAIL.n222 VTAIL.n221 185
R2090 VTAIL.n307 VTAIL.n306 185
R2091 VTAIL.n305 VTAIL.n304 185
R2092 VTAIL.n226 VTAIL.n225 185
R2093 VTAIL.n299 VTAIL.n298 185
R2094 VTAIL.n297 VTAIL.n228 185
R2095 VTAIL.n296 VTAIL.n295 185
R2096 VTAIL.n231 VTAIL.n229 185
R2097 VTAIL.n290 VTAIL.n289 185
R2098 VTAIL.n288 VTAIL.n287 185
R2099 VTAIL.n235 VTAIL.n234 185
R2100 VTAIL.n282 VTAIL.n281 185
R2101 VTAIL.n280 VTAIL.n279 185
R2102 VTAIL.n239 VTAIL.n238 185
R2103 VTAIL.n274 VTAIL.n273 185
R2104 VTAIL.n272 VTAIL.n271 185
R2105 VTAIL.n243 VTAIL.n242 185
R2106 VTAIL.n266 VTAIL.n265 185
R2107 VTAIL.n264 VTAIL.n263 185
R2108 VTAIL.n247 VTAIL.n246 185
R2109 VTAIL.n258 VTAIL.n257 185
R2110 VTAIL.n256 VTAIL.n255 185
R2111 VTAIL.n251 VTAIL.n250 185
R2112 VTAIL.n209 VTAIL.n208 185
R2113 VTAIL.n207 VTAIL.n206 185
R2114 VTAIL.n116 VTAIL.n115 185
R2115 VTAIL.n201 VTAIL.n200 185
R2116 VTAIL.n199 VTAIL.n198 185
R2117 VTAIL.n120 VTAIL.n119 185
R2118 VTAIL.n193 VTAIL.n192 185
R2119 VTAIL.n191 VTAIL.n122 185
R2120 VTAIL.n190 VTAIL.n189 185
R2121 VTAIL.n125 VTAIL.n123 185
R2122 VTAIL.n184 VTAIL.n183 185
R2123 VTAIL.n182 VTAIL.n181 185
R2124 VTAIL.n129 VTAIL.n128 185
R2125 VTAIL.n176 VTAIL.n175 185
R2126 VTAIL.n174 VTAIL.n173 185
R2127 VTAIL.n133 VTAIL.n132 185
R2128 VTAIL.n168 VTAIL.n167 185
R2129 VTAIL.n166 VTAIL.n165 185
R2130 VTAIL.n137 VTAIL.n136 185
R2131 VTAIL.n160 VTAIL.n159 185
R2132 VTAIL.n158 VTAIL.n157 185
R2133 VTAIL.n141 VTAIL.n140 185
R2134 VTAIL.n152 VTAIL.n151 185
R2135 VTAIL.n150 VTAIL.n149 185
R2136 VTAIL.n145 VTAIL.n144 185
R2137 VTAIL.n353 VTAIL.t16 147.659
R2138 VTAIL.n35 VTAIL.t3 147.659
R2139 VTAIL.n252 VTAIL.t4 147.659
R2140 VTAIL.n146 VTAIL.t11 147.659
R2141 VTAIL.n357 VTAIL.n351 104.615
R2142 VTAIL.n358 VTAIL.n357 104.615
R2143 VTAIL.n358 VTAIL.n347 104.615
R2144 VTAIL.n365 VTAIL.n347 104.615
R2145 VTAIL.n366 VTAIL.n365 104.615
R2146 VTAIL.n366 VTAIL.n343 104.615
R2147 VTAIL.n373 VTAIL.n343 104.615
R2148 VTAIL.n374 VTAIL.n373 104.615
R2149 VTAIL.n374 VTAIL.n339 104.615
R2150 VTAIL.n381 VTAIL.n339 104.615
R2151 VTAIL.n382 VTAIL.n381 104.615
R2152 VTAIL.n382 VTAIL.n335 104.615
R2153 VTAIL.n389 VTAIL.n335 104.615
R2154 VTAIL.n390 VTAIL.n389 104.615
R2155 VTAIL.n390 VTAIL.n331 104.615
R2156 VTAIL.n398 VTAIL.n331 104.615
R2157 VTAIL.n399 VTAIL.n398 104.615
R2158 VTAIL.n400 VTAIL.n399 104.615
R2159 VTAIL.n400 VTAIL.n327 104.615
R2160 VTAIL.n407 VTAIL.n327 104.615
R2161 VTAIL.n408 VTAIL.n407 104.615
R2162 VTAIL.n408 VTAIL.n323 104.615
R2163 VTAIL.n415 VTAIL.n323 104.615
R2164 VTAIL.n416 VTAIL.n415 104.615
R2165 VTAIL.n39 VTAIL.n33 104.615
R2166 VTAIL.n40 VTAIL.n39 104.615
R2167 VTAIL.n40 VTAIL.n29 104.615
R2168 VTAIL.n47 VTAIL.n29 104.615
R2169 VTAIL.n48 VTAIL.n47 104.615
R2170 VTAIL.n48 VTAIL.n25 104.615
R2171 VTAIL.n55 VTAIL.n25 104.615
R2172 VTAIL.n56 VTAIL.n55 104.615
R2173 VTAIL.n56 VTAIL.n21 104.615
R2174 VTAIL.n63 VTAIL.n21 104.615
R2175 VTAIL.n64 VTAIL.n63 104.615
R2176 VTAIL.n64 VTAIL.n17 104.615
R2177 VTAIL.n71 VTAIL.n17 104.615
R2178 VTAIL.n72 VTAIL.n71 104.615
R2179 VTAIL.n72 VTAIL.n13 104.615
R2180 VTAIL.n80 VTAIL.n13 104.615
R2181 VTAIL.n81 VTAIL.n80 104.615
R2182 VTAIL.n82 VTAIL.n81 104.615
R2183 VTAIL.n82 VTAIL.n9 104.615
R2184 VTAIL.n89 VTAIL.n9 104.615
R2185 VTAIL.n90 VTAIL.n89 104.615
R2186 VTAIL.n90 VTAIL.n5 104.615
R2187 VTAIL.n97 VTAIL.n5 104.615
R2188 VTAIL.n98 VTAIL.n97 104.615
R2189 VTAIL.n314 VTAIL.n313 104.615
R2190 VTAIL.n313 VTAIL.n221 104.615
R2191 VTAIL.n306 VTAIL.n221 104.615
R2192 VTAIL.n306 VTAIL.n305 104.615
R2193 VTAIL.n305 VTAIL.n225 104.615
R2194 VTAIL.n298 VTAIL.n225 104.615
R2195 VTAIL.n298 VTAIL.n297 104.615
R2196 VTAIL.n297 VTAIL.n296 104.615
R2197 VTAIL.n296 VTAIL.n229 104.615
R2198 VTAIL.n289 VTAIL.n229 104.615
R2199 VTAIL.n289 VTAIL.n288 104.615
R2200 VTAIL.n288 VTAIL.n234 104.615
R2201 VTAIL.n281 VTAIL.n234 104.615
R2202 VTAIL.n281 VTAIL.n280 104.615
R2203 VTAIL.n280 VTAIL.n238 104.615
R2204 VTAIL.n273 VTAIL.n238 104.615
R2205 VTAIL.n273 VTAIL.n272 104.615
R2206 VTAIL.n272 VTAIL.n242 104.615
R2207 VTAIL.n265 VTAIL.n242 104.615
R2208 VTAIL.n265 VTAIL.n264 104.615
R2209 VTAIL.n264 VTAIL.n246 104.615
R2210 VTAIL.n257 VTAIL.n246 104.615
R2211 VTAIL.n257 VTAIL.n256 104.615
R2212 VTAIL.n256 VTAIL.n250 104.615
R2213 VTAIL.n208 VTAIL.n207 104.615
R2214 VTAIL.n207 VTAIL.n115 104.615
R2215 VTAIL.n200 VTAIL.n115 104.615
R2216 VTAIL.n200 VTAIL.n199 104.615
R2217 VTAIL.n199 VTAIL.n119 104.615
R2218 VTAIL.n192 VTAIL.n119 104.615
R2219 VTAIL.n192 VTAIL.n191 104.615
R2220 VTAIL.n191 VTAIL.n190 104.615
R2221 VTAIL.n190 VTAIL.n123 104.615
R2222 VTAIL.n183 VTAIL.n123 104.615
R2223 VTAIL.n183 VTAIL.n182 104.615
R2224 VTAIL.n182 VTAIL.n128 104.615
R2225 VTAIL.n175 VTAIL.n128 104.615
R2226 VTAIL.n175 VTAIL.n174 104.615
R2227 VTAIL.n174 VTAIL.n132 104.615
R2228 VTAIL.n167 VTAIL.n132 104.615
R2229 VTAIL.n167 VTAIL.n166 104.615
R2230 VTAIL.n166 VTAIL.n136 104.615
R2231 VTAIL.n159 VTAIL.n136 104.615
R2232 VTAIL.n159 VTAIL.n158 104.615
R2233 VTAIL.n158 VTAIL.n140 104.615
R2234 VTAIL.n151 VTAIL.n140 104.615
R2235 VTAIL.n151 VTAIL.n150 104.615
R2236 VTAIL.n150 VTAIL.n144 104.615
R2237 VTAIL.t16 VTAIL.n351 52.3082
R2238 VTAIL.t3 VTAIL.n33 52.3082
R2239 VTAIL.t4 VTAIL.n250 52.3082
R2240 VTAIL.t11 VTAIL.n144 52.3082
R2241 VTAIL.n217 VTAIL.n216 43.9695
R2242 VTAIL.n215 VTAIL.n214 43.9695
R2243 VTAIL.n111 VTAIL.n110 43.9695
R2244 VTAIL.n109 VTAIL.n108 43.9695
R2245 VTAIL.n423 VTAIL.n422 43.9693
R2246 VTAIL.n1 VTAIL.n0 43.9693
R2247 VTAIL.n105 VTAIL.n104 43.9693
R2248 VTAIL.n107 VTAIL.n106 43.9693
R2249 VTAIL.n421 VTAIL.n420 32.1853
R2250 VTAIL.n103 VTAIL.n102 32.1853
R2251 VTAIL.n319 VTAIL.n318 32.1853
R2252 VTAIL.n213 VTAIL.n212 32.1853
R2253 VTAIL.n109 VTAIL.n107 31.8841
R2254 VTAIL.n421 VTAIL.n319 29.9876
R2255 VTAIL.n353 VTAIL.n352 15.6677
R2256 VTAIL.n35 VTAIL.n34 15.6677
R2257 VTAIL.n252 VTAIL.n251 15.6677
R2258 VTAIL.n146 VTAIL.n145 15.6677
R2259 VTAIL.n401 VTAIL.n330 13.1884
R2260 VTAIL.n83 VTAIL.n12 13.1884
R2261 VTAIL.n299 VTAIL.n228 13.1884
R2262 VTAIL.n193 VTAIL.n122 13.1884
R2263 VTAIL.n356 VTAIL.n355 12.8005
R2264 VTAIL.n397 VTAIL.n396 12.8005
R2265 VTAIL.n402 VTAIL.n328 12.8005
R2266 VTAIL.n38 VTAIL.n37 12.8005
R2267 VTAIL.n79 VTAIL.n78 12.8005
R2268 VTAIL.n84 VTAIL.n10 12.8005
R2269 VTAIL.n300 VTAIL.n226 12.8005
R2270 VTAIL.n295 VTAIL.n230 12.8005
R2271 VTAIL.n255 VTAIL.n254 12.8005
R2272 VTAIL.n194 VTAIL.n120 12.8005
R2273 VTAIL.n189 VTAIL.n124 12.8005
R2274 VTAIL.n149 VTAIL.n148 12.8005
R2275 VTAIL.n359 VTAIL.n350 12.0247
R2276 VTAIL.n395 VTAIL.n332 12.0247
R2277 VTAIL.n406 VTAIL.n405 12.0247
R2278 VTAIL.n41 VTAIL.n32 12.0247
R2279 VTAIL.n77 VTAIL.n14 12.0247
R2280 VTAIL.n88 VTAIL.n87 12.0247
R2281 VTAIL.n304 VTAIL.n303 12.0247
R2282 VTAIL.n294 VTAIL.n231 12.0247
R2283 VTAIL.n258 VTAIL.n249 12.0247
R2284 VTAIL.n198 VTAIL.n197 12.0247
R2285 VTAIL.n188 VTAIL.n125 12.0247
R2286 VTAIL.n152 VTAIL.n143 12.0247
R2287 VTAIL.n360 VTAIL.n348 11.249
R2288 VTAIL.n392 VTAIL.n391 11.249
R2289 VTAIL.n409 VTAIL.n326 11.249
R2290 VTAIL.n42 VTAIL.n30 11.249
R2291 VTAIL.n74 VTAIL.n73 11.249
R2292 VTAIL.n91 VTAIL.n8 11.249
R2293 VTAIL.n307 VTAIL.n224 11.249
R2294 VTAIL.n291 VTAIL.n290 11.249
R2295 VTAIL.n259 VTAIL.n247 11.249
R2296 VTAIL.n201 VTAIL.n118 11.249
R2297 VTAIL.n185 VTAIL.n184 11.249
R2298 VTAIL.n153 VTAIL.n141 11.249
R2299 VTAIL.n364 VTAIL.n363 10.4732
R2300 VTAIL.n388 VTAIL.n334 10.4732
R2301 VTAIL.n410 VTAIL.n324 10.4732
R2302 VTAIL.n46 VTAIL.n45 10.4732
R2303 VTAIL.n70 VTAIL.n16 10.4732
R2304 VTAIL.n92 VTAIL.n6 10.4732
R2305 VTAIL.n308 VTAIL.n222 10.4732
R2306 VTAIL.n287 VTAIL.n233 10.4732
R2307 VTAIL.n263 VTAIL.n262 10.4732
R2308 VTAIL.n202 VTAIL.n116 10.4732
R2309 VTAIL.n181 VTAIL.n127 10.4732
R2310 VTAIL.n157 VTAIL.n156 10.4732
R2311 VTAIL.n367 VTAIL.n346 9.69747
R2312 VTAIL.n387 VTAIL.n336 9.69747
R2313 VTAIL.n414 VTAIL.n413 9.69747
R2314 VTAIL.n49 VTAIL.n28 9.69747
R2315 VTAIL.n69 VTAIL.n18 9.69747
R2316 VTAIL.n96 VTAIL.n95 9.69747
R2317 VTAIL.n312 VTAIL.n311 9.69747
R2318 VTAIL.n286 VTAIL.n235 9.69747
R2319 VTAIL.n266 VTAIL.n245 9.69747
R2320 VTAIL.n206 VTAIL.n205 9.69747
R2321 VTAIL.n180 VTAIL.n129 9.69747
R2322 VTAIL.n160 VTAIL.n139 9.69747
R2323 VTAIL.n420 VTAIL.n419 9.45567
R2324 VTAIL.n102 VTAIL.n101 9.45567
R2325 VTAIL.n318 VTAIL.n317 9.45567
R2326 VTAIL.n212 VTAIL.n211 9.45567
R2327 VTAIL.n419 VTAIL.n418 9.3005
R2328 VTAIL.n322 VTAIL.n321 9.3005
R2329 VTAIL.n413 VTAIL.n412 9.3005
R2330 VTAIL.n411 VTAIL.n410 9.3005
R2331 VTAIL.n326 VTAIL.n325 9.3005
R2332 VTAIL.n405 VTAIL.n404 9.3005
R2333 VTAIL.n403 VTAIL.n402 9.3005
R2334 VTAIL.n342 VTAIL.n341 9.3005
R2335 VTAIL.n371 VTAIL.n370 9.3005
R2336 VTAIL.n369 VTAIL.n368 9.3005
R2337 VTAIL.n346 VTAIL.n345 9.3005
R2338 VTAIL.n363 VTAIL.n362 9.3005
R2339 VTAIL.n361 VTAIL.n360 9.3005
R2340 VTAIL.n350 VTAIL.n349 9.3005
R2341 VTAIL.n355 VTAIL.n354 9.3005
R2342 VTAIL.n377 VTAIL.n376 9.3005
R2343 VTAIL.n379 VTAIL.n378 9.3005
R2344 VTAIL.n338 VTAIL.n337 9.3005
R2345 VTAIL.n385 VTAIL.n384 9.3005
R2346 VTAIL.n387 VTAIL.n386 9.3005
R2347 VTAIL.n334 VTAIL.n333 9.3005
R2348 VTAIL.n393 VTAIL.n392 9.3005
R2349 VTAIL.n395 VTAIL.n394 9.3005
R2350 VTAIL.n396 VTAIL.n329 9.3005
R2351 VTAIL.n101 VTAIL.n100 9.3005
R2352 VTAIL.n4 VTAIL.n3 9.3005
R2353 VTAIL.n95 VTAIL.n94 9.3005
R2354 VTAIL.n93 VTAIL.n92 9.3005
R2355 VTAIL.n8 VTAIL.n7 9.3005
R2356 VTAIL.n87 VTAIL.n86 9.3005
R2357 VTAIL.n85 VTAIL.n84 9.3005
R2358 VTAIL.n24 VTAIL.n23 9.3005
R2359 VTAIL.n53 VTAIL.n52 9.3005
R2360 VTAIL.n51 VTAIL.n50 9.3005
R2361 VTAIL.n28 VTAIL.n27 9.3005
R2362 VTAIL.n45 VTAIL.n44 9.3005
R2363 VTAIL.n43 VTAIL.n42 9.3005
R2364 VTAIL.n32 VTAIL.n31 9.3005
R2365 VTAIL.n37 VTAIL.n36 9.3005
R2366 VTAIL.n59 VTAIL.n58 9.3005
R2367 VTAIL.n61 VTAIL.n60 9.3005
R2368 VTAIL.n20 VTAIL.n19 9.3005
R2369 VTAIL.n67 VTAIL.n66 9.3005
R2370 VTAIL.n69 VTAIL.n68 9.3005
R2371 VTAIL.n16 VTAIL.n15 9.3005
R2372 VTAIL.n75 VTAIL.n74 9.3005
R2373 VTAIL.n77 VTAIL.n76 9.3005
R2374 VTAIL.n78 VTAIL.n11 9.3005
R2375 VTAIL.n278 VTAIL.n277 9.3005
R2376 VTAIL.n237 VTAIL.n236 9.3005
R2377 VTAIL.n284 VTAIL.n283 9.3005
R2378 VTAIL.n286 VTAIL.n285 9.3005
R2379 VTAIL.n233 VTAIL.n232 9.3005
R2380 VTAIL.n292 VTAIL.n291 9.3005
R2381 VTAIL.n294 VTAIL.n293 9.3005
R2382 VTAIL.n230 VTAIL.n227 9.3005
R2383 VTAIL.n317 VTAIL.n316 9.3005
R2384 VTAIL.n220 VTAIL.n219 9.3005
R2385 VTAIL.n311 VTAIL.n310 9.3005
R2386 VTAIL.n309 VTAIL.n308 9.3005
R2387 VTAIL.n224 VTAIL.n223 9.3005
R2388 VTAIL.n303 VTAIL.n302 9.3005
R2389 VTAIL.n301 VTAIL.n300 9.3005
R2390 VTAIL.n276 VTAIL.n275 9.3005
R2391 VTAIL.n241 VTAIL.n240 9.3005
R2392 VTAIL.n270 VTAIL.n269 9.3005
R2393 VTAIL.n268 VTAIL.n267 9.3005
R2394 VTAIL.n245 VTAIL.n244 9.3005
R2395 VTAIL.n262 VTAIL.n261 9.3005
R2396 VTAIL.n260 VTAIL.n259 9.3005
R2397 VTAIL.n249 VTAIL.n248 9.3005
R2398 VTAIL.n254 VTAIL.n253 9.3005
R2399 VTAIL.n172 VTAIL.n171 9.3005
R2400 VTAIL.n131 VTAIL.n130 9.3005
R2401 VTAIL.n178 VTAIL.n177 9.3005
R2402 VTAIL.n180 VTAIL.n179 9.3005
R2403 VTAIL.n127 VTAIL.n126 9.3005
R2404 VTAIL.n186 VTAIL.n185 9.3005
R2405 VTAIL.n188 VTAIL.n187 9.3005
R2406 VTAIL.n124 VTAIL.n121 9.3005
R2407 VTAIL.n211 VTAIL.n210 9.3005
R2408 VTAIL.n114 VTAIL.n113 9.3005
R2409 VTAIL.n205 VTAIL.n204 9.3005
R2410 VTAIL.n203 VTAIL.n202 9.3005
R2411 VTAIL.n118 VTAIL.n117 9.3005
R2412 VTAIL.n197 VTAIL.n196 9.3005
R2413 VTAIL.n195 VTAIL.n194 9.3005
R2414 VTAIL.n170 VTAIL.n169 9.3005
R2415 VTAIL.n135 VTAIL.n134 9.3005
R2416 VTAIL.n164 VTAIL.n163 9.3005
R2417 VTAIL.n162 VTAIL.n161 9.3005
R2418 VTAIL.n139 VTAIL.n138 9.3005
R2419 VTAIL.n156 VTAIL.n155 9.3005
R2420 VTAIL.n154 VTAIL.n153 9.3005
R2421 VTAIL.n143 VTAIL.n142 9.3005
R2422 VTAIL.n148 VTAIL.n147 9.3005
R2423 VTAIL.n368 VTAIL.n344 8.92171
R2424 VTAIL.n384 VTAIL.n383 8.92171
R2425 VTAIL.n417 VTAIL.n322 8.92171
R2426 VTAIL.n50 VTAIL.n26 8.92171
R2427 VTAIL.n66 VTAIL.n65 8.92171
R2428 VTAIL.n99 VTAIL.n4 8.92171
R2429 VTAIL.n315 VTAIL.n220 8.92171
R2430 VTAIL.n283 VTAIL.n282 8.92171
R2431 VTAIL.n267 VTAIL.n243 8.92171
R2432 VTAIL.n209 VTAIL.n114 8.92171
R2433 VTAIL.n177 VTAIL.n176 8.92171
R2434 VTAIL.n161 VTAIL.n137 8.92171
R2435 VTAIL.n372 VTAIL.n371 8.14595
R2436 VTAIL.n380 VTAIL.n338 8.14595
R2437 VTAIL.n418 VTAIL.n320 8.14595
R2438 VTAIL.n54 VTAIL.n53 8.14595
R2439 VTAIL.n62 VTAIL.n20 8.14595
R2440 VTAIL.n100 VTAIL.n2 8.14595
R2441 VTAIL.n316 VTAIL.n218 8.14595
R2442 VTAIL.n279 VTAIL.n237 8.14595
R2443 VTAIL.n271 VTAIL.n270 8.14595
R2444 VTAIL.n210 VTAIL.n112 8.14595
R2445 VTAIL.n173 VTAIL.n131 8.14595
R2446 VTAIL.n165 VTAIL.n164 8.14595
R2447 VTAIL.n375 VTAIL.n342 7.3702
R2448 VTAIL.n379 VTAIL.n340 7.3702
R2449 VTAIL.n57 VTAIL.n24 7.3702
R2450 VTAIL.n61 VTAIL.n22 7.3702
R2451 VTAIL.n278 VTAIL.n239 7.3702
R2452 VTAIL.n274 VTAIL.n241 7.3702
R2453 VTAIL.n172 VTAIL.n133 7.3702
R2454 VTAIL.n168 VTAIL.n135 7.3702
R2455 VTAIL.n376 VTAIL.n375 6.59444
R2456 VTAIL.n376 VTAIL.n340 6.59444
R2457 VTAIL.n58 VTAIL.n57 6.59444
R2458 VTAIL.n58 VTAIL.n22 6.59444
R2459 VTAIL.n275 VTAIL.n239 6.59444
R2460 VTAIL.n275 VTAIL.n274 6.59444
R2461 VTAIL.n169 VTAIL.n133 6.59444
R2462 VTAIL.n169 VTAIL.n168 6.59444
R2463 VTAIL.n372 VTAIL.n342 5.81868
R2464 VTAIL.n380 VTAIL.n379 5.81868
R2465 VTAIL.n420 VTAIL.n320 5.81868
R2466 VTAIL.n54 VTAIL.n24 5.81868
R2467 VTAIL.n62 VTAIL.n61 5.81868
R2468 VTAIL.n102 VTAIL.n2 5.81868
R2469 VTAIL.n318 VTAIL.n218 5.81868
R2470 VTAIL.n279 VTAIL.n278 5.81868
R2471 VTAIL.n271 VTAIL.n241 5.81868
R2472 VTAIL.n212 VTAIL.n112 5.81868
R2473 VTAIL.n173 VTAIL.n172 5.81868
R2474 VTAIL.n165 VTAIL.n135 5.81868
R2475 VTAIL.n371 VTAIL.n344 5.04292
R2476 VTAIL.n383 VTAIL.n338 5.04292
R2477 VTAIL.n418 VTAIL.n417 5.04292
R2478 VTAIL.n53 VTAIL.n26 5.04292
R2479 VTAIL.n65 VTAIL.n20 5.04292
R2480 VTAIL.n100 VTAIL.n99 5.04292
R2481 VTAIL.n316 VTAIL.n315 5.04292
R2482 VTAIL.n282 VTAIL.n237 5.04292
R2483 VTAIL.n270 VTAIL.n243 5.04292
R2484 VTAIL.n210 VTAIL.n209 5.04292
R2485 VTAIL.n176 VTAIL.n131 5.04292
R2486 VTAIL.n164 VTAIL.n137 5.04292
R2487 VTAIL.n354 VTAIL.n353 4.38563
R2488 VTAIL.n36 VTAIL.n35 4.38563
R2489 VTAIL.n253 VTAIL.n252 4.38563
R2490 VTAIL.n147 VTAIL.n146 4.38563
R2491 VTAIL.n368 VTAIL.n367 4.26717
R2492 VTAIL.n384 VTAIL.n336 4.26717
R2493 VTAIL.n414 VTAIL.n322 4.26717
R2494 VTAIL.n50 VTAIL.n49 4.26717
R2495 VTAIL.n66 VTAIL.n18 4.26717
R2496 VTAIL.n96 VTAIL.n4 4.26717
R2497 VTAIL.n312 VTAIL.n220 4.26717
R2498 VTAIL.n283 VTAIL.n235 4.26717
R2499 VTAIL.n267 VTAIL.n266 4.26717
R2500 VTAIL.n206 VTAIL.n114 4.26717
R2501 VTAIL.n177 VTAIL.n129 4.26717
R2502 VTAIL.n161 VTAIL.n160 4.26717
R2503 VTAIL.n364 VTAIL.n346 3.49141
R2504 VTAIL.n388 VTAIL.n387 3.49141
R2505 VTAIL.n413 VTAIL.n324 3.49141
R2506 VTAIL.n46 VTAIL.n28 3.49141
R2507 VTAIL.n70 VTAIL.n69 3.49141
R2508 VTAIL.n95 VTAIL.n6 3.49141
R2509 VTAIL.n311 VTAIL.n222 3.49141
R2510 VTAIL.n287 VTAIL.n286 3.49141
R2511 VTAIL.n263 VTAIL.n245 3.49141
R2512 VTAIL.n205 VTAIL.n116 3.49141
R2513 VTAIL.n181 VTAIL.n180 3.49141
R2514 VTAIL.n157 VTAIL.n139 3.49141
R2515 VTAIL.n363 VTAIL.n348 2.71565
R2516 VTAIL.n391 VTAIL.n334 2.71565
R2517 VTAIL.n410 VTAIL.n409 2.71565
R2518 VTAIL.n45 VTAIL.n30 2.71565
R2519 VTAIL.n73 VTAIL.n16 2.71565
R2520 VTAIL.n92 VTAIL.n91 2.71565
R2521 VTAIL.n308 VTAIL.n307 2.71565
R2522 VTAIL.n290 VTAIL.n233 2.71565
R2523 VTAIL.n262 VTAIL.n247 2.71565
R2524 VTAIL.n202 VTAIL.n201 2.71565
R2525 VTAIL.n184 VTAIL.n127 2.71565
R2526 VTAIL.n156 VTAIL.n141 2.71565
R2527 VTAIL.n360 VTAIL.n359 1.93989
R2528 VTAIL.n392 VTAIL.n332 1.93989
R2529 VTAIL.n406 VTAIL.n326 1.93989
R2530 VTAIL.n42 VTAIL.n41 1.93989
R2531 VTAIL.n74 VTAIL.n14 1.93989
R2532 VTAIL.n88 VTAIL.n8 1.93989
R2533 VTAIL.n304 VTAIL.n224 1.93989
R2534 VTAIL.n291 VTAIL.n231 1.93989
R2535 VTAIL.n259 VTAIL.n258 1.93989
R2536 VTAIL.n198 VTAIL.n118 1.93989
R2537 VTAIL.n185 VTAIL.n125 1.93989
R2538 VTAIL.n153 VTAIL.n152 1.93989
R2539 VTAIL.n111 VTAIL.n109 1.89705
R2540 VTAIL.n213 VTAIL.n111 1.89705
R2541 VTAIL.n217 VTAIL.n215 1.89705
R2542 VTAIL.n319 VTAIL.n217 1.89705
R2543 VTAIL.n107 VTAIL.n105 1.89705
R2544 VTAIL.n105 VTAIL.n103 1.89705
R2545 VTAIL.n423 VTAIL.n421 1.89705
R2546 VTAIL VTAIL.n1 1.4811
R2547 VTAIL.n215 VTAIL.n213 1.4186
R2548 VTAIL.n103 VTAIL.n1 1.4186
R2549 VTAIL.n356 VTAIL.n350 1.16414
R2550 VTAIL.n397 VTAIL.n395 1.16414
R2551 VTAIL.n405 VTAIL.n328 1.16414
R2552 VTAIL.n38 VTAIL.n32 1.16414
R2553 VTAIL.n79 VTAIL.n77 1.16414
R2554 VTAIL.n87 VTAIL.n10 1.16414
R2555 VTAIL.n303 VTAIL.n226 1.16414
R2556 VTAIL.n295 VTAIL.n294 1.16414
R2557 VTAIL.n255 VTAIL.n249 1.16414
R2558 VTAIL.n197 VTAIL.n120 1.16414
R2559 VTAIL.n189 VTAIL.n188 1.16414
R2560 VTAIL.n149 VTAIL.n143 1.16414
R2561 VTAIL.n422 VTAIL.t17 1.08603
R2562 VTAIL.n422 VTAIL.t19 1.08603
R2563 VTAIL.n0 VTAIL.t10 1.08603
R2564 VTAIL.n0 VTAIL.t13 1.08603
R2565 VTAIL.n104 VTAIL.t1 1.08603
R2566 VTAIL.n104 VTAIL.t9 1.08603
R2567 VTAIL.n106 VTAIL.t7 1.08603
R2568 VTAIL.n106 VTAIL.t2 1.08603
R2569 VTAIL.n216 VTAIL.t5 1.08603
R2570 VTAIL.n216 VTAIL.t0 1.08603
R2571 VTAIL.n214 VTAIL.t6 1.08603
R2572 VTAIL.n214 VTAIL.t8 1.08603
R2573 VTAIL.n110 VTAIL.t14 1.08603
R2574 VTAIL.n110 VTAIL.t15 1.08603
R2575 VTAIL.n108 VTAIL.t18 1.08603
R2576 VTAIL.n108 VTAIL.t12 1.08603
R2577 VTAIL VTAIL.n423 0.416448
R2578 VTAIL.n355 VTAIL.n352 0.388379
R2579 VTAIL.n396 VTAIL.n330 0.388379
R2580 VTAIL.n402 VTAIL.n401 0.388379
R2581 VTAIL.n37 VTAIL.n34 0.388379
R2582 VTAIL.n78 VTAIL.n12 0.388379
R2583 VTAIL.n84 VTAIL.n83 0.388379
R2584 VTAIL.n300 VTAIL.n299 0.388379
R2585 VTAIL.n230 VTAIL.n228 0.388379
R2586 VTAIL.n254 VTAIL.n251 0.388379
R2587 VTAIL.n194 VTAIL.n193 0.388379
R2588 VTAIL.n124 VTAIL.n122 0.388379
R2589 VTAIL.n148 VTAIL.n145 0.388379
R2590 VTAIL.n354 VTAIL.n349 0.155672
R2591 VTAIL.n361 VTAIL.n349 0.155672
R2592 VTAIL.n362 VTAIL.n361 0.155672
R2593 VTAIL.n362 VTAIL.n345 0.155672
R2594 VTAIL.n369 VTAIL.n345 0.155672
R2595 VTAIL.n370 VTAIL.n369 0.155672
R2596 VTAIL.n370 VTAIL.n341 0.155672
R2597 VTAIL.n377 VTAIL.n341 0.155672
R2598 VTAIL.n378 VTAIL.n377 0.155672
R2599 VTAIL.n378 VTAIL.n337 0.155672
R2600 VTAIL.n385 VTAIL.n337 0.155672
R2601 VTAIL.n386 VTAIL.n385 0.155672
R2602 VTAIL.n386 VTAIL.n333 0.155672
R2603 VTAIL.n393 VTAIL.n333 0.155672
R2604 VTAIL.n394 VTAIL.n393 0.155672
R2605 VTAIL.n394 VTAIL.n329 0.155672
R2606 VTAIL.n403 VTAIL.n329 0.155672
R2607 VTAIL.n404 VTAIL.n403 0.155672
R2608 VTAIL.n404 VTAIL.n325 0.155672
R2609 VTAIL.n411 VTAIL.n325 0.155672
R2610 VTAIL.n412 VTAIL.n411 0.155672
R2611 VTAIL.n412 VTAIL.n321 0.155672
R2612 VTAIL.n419 VTAIL.n321 0.155672
R2613 VTAIL.n36 VTAIL.n31 0.155672
R2614 VTAIL.n43 VTAIL.n31 0.155672
R2615 VTAIL.n44 VTAIL.n43 0.155672
R2616 VTAIL.n44 VTAIL.n27 0.155672
R2617 VTAIL.n51 VTAIL.n27 0.155672
R2618 VTAIL.n52 VTAIL.n51 0.155672
R2619 VTAIL.n52 VTAIL.n23 0.155672
R2620 VTAIL.n59 VTAIL.n23 0.155672
R2621 VTAIL.n60 VTAIL.n59 0.155672
R2622 VTAIL.n60 VTAIL.n19 0.155672
R2623 VTAIL.n67 VTAIL.n19 0.155672
R2624 VTAIL.n68 VTAIL.n67 0.155672
R2625 VTAIL.n68 VTAIL.n15 0.155672
R2626 VTAIL.n75 VTAIL.n15 0.155672
R2627 VTAIL.n76 VTAIL.n75 0.155672
R2628 VTAIL.n76 VTAIL.n11 0.155672
R2629 VTAIL.n85 VTAIL.n11 0.155672
R2630 VTAIL.n86 VTAIL.n85 0.155672
R2631 VTAIL.n86 VTAIL.n7 0.155672
R2632 VTAIL.n93 VTAIL.n7 0.155672
R2633 VTAIL.n94 VTAIL.n93 0.155672
R2634 VTAIL.n94 VTAIL.n3 0.155672
R2635 VTAIL.n101 VTAIL.n3 0.155672
R2636 VTAIL.n317 VTAIL.n219 0.155672
R2637 VTAIL.n310 VTAIL.n219 0.155672
R2638 VTAIL.n310 VTAIL.n309 0.155672
R2639 VTAIL.n309 VTAIL.n223 0.155672
R2640 VTAIL.n302 VTAIL.n223 0.155672
R2641 VTAIL.n302 VTAIL.n301 0.155672
R2642 VTAIL.n301 VTAIL.n227 0.155672
R2643 VTAIL.n293 VTAIL.n227 0.155672
R2644 VTAIL.n293 VTAIL.n292 0.155672
R2645 VTAIL.n292 VTAIL.n232 0.155672
R2646 VTAIL.n285 VTAIL.n232 0.155672
R2647 VTAIL.n285 VTAIL.n284 0.155672
R2648 VTAIL.n284 VTAIL.n236 0.155672
R2649 VTAIL.n277 VTAIL.n236 0.155672
R2650 VTAIL.n277 VTAIL.n276 0.155672
R2651 VTAIL.n276 VTAIL.n240 0.155672
R2652 VTAIL.n269 VTAIL.n240 0.155672
R2653 VTAIL.n269 VTAIL.n268 0.155672
R2654 VTAIL.n268 VTAIL.n244 0.155672
R2655 VTAIL.n261 VTAIL.n244 0.155672
R2656 VTAIL.n261 VTAIL.n260 0.155672
R2657 VTAIL.n260 VTAIL.n248 0.155672
R2658 VTAIL.n253 VTAIL.n248 0.155672
R2659 VTAIL.n211 VTAIL.n113 0.155672
R2660 VTAIL.n204 VTAIL.n113 0.155672
R2661 VTAIL.n204 VTAIL.n203 0.155672
R2662 VTAIL.n203 VTAIL.n117 0.155672
R2663 VTAIL.n196 VTAIL.n117 0.155672
R2664 VTAIL.n196 VTAIL.n195 0.155672
R2665 VTAIL.n195 VTAIL.n121 0.155672
R2666 VTAIL.n187 VTAIL.n121 0.155672
R2667 VTAIL.n187 VTAIL.n186 0.155672
R2668 VTAIL.n186 VTAIL.n126 0.155672
R2669 VTAIL.n179 VTAIL.n126 0.155672
R2670 VTAIL.n179 VTAIL.n178 0.155672
R2671 VTAIL.n178 VTAIL.n130 0.155672
R2672 VTAIL.n171 VTAIL.n130 0.155672
R2673 VTAIL.n171 VTAIL.n170 0.155672
R2674 VTAIL.n170 VTAIL.n134 0.155672
R2675 VTAIL.n163 VTAIL.n134 0.155672
R2676 VTAIL.n163 VTAIL.n162 0.155672
R2677 VTAIL.n162 VTAIL.n138 0.155672
R2678 VTAIL.n155 VTAIL.n138 0.155672
R2679 VTAIL.n155 VTAIL.n154 0.155672
R2680 VTAIL.n154 VTAIL.n142 0.155672
R2681 VTAIL.n147 VTAIL.n142 0.155672
R2682 VDD2.n201 VDD2.n105 289.615
R2683 VDD2.n96 VDD2.n0 289.615
R2684 VDD2.n202 VDD2.n201 185
R2685 VDD2.n200 VDD2.n199 185
R2686 VDD2.n109 VDD2.n108 185
R2687 VDD2.n194 VDD2.n193 185
R2688 VDD2.n192 VDD2.n191 185
R2689 VDD2.n113 VDD2.n112 185
R2690 VDD2.n186 VDD2.n185 185
R2691 VDD2.n184 VDD2.n115 185
R2692 VDD2.n183 VDD2.n182 185
R2693 VDD2.n118 VDD2.n116 185
R2694 VDD2.n177 VDD2.n176 185
R2695 VDD2.n175 VDD2.n174 185
R2696 VDD2.n122 VDD2.n121 185
R2697 VDD2.n169 VDD2.n168 185
R2698 VDD2.n167 VDD2.n166 185
R2699 VDD2.n126 VDD2.n125 185
R2700 VDD2.n161 VDD2.n160 185
R2701 VDD2.n159 VDD2.n158 185
R2702 VDD2.n130 VDD2.n129 185
R2703 VDD2.n153 VDD2.n152 185
R2704 VDD2.n151 VDD2.n150 185
R2705 VDD2.n134 VDD2.n133 185
R2706 VDD2.n145 VDD2.n144 185
R2707 VDD2.n143 VDD2.n142 185
R2708 VDD2.n138 VDD2.n137 185
R2709 VDD2.n32 VDD2.n31 185
R2710 VDD2.n37 VDD2.n36 185
R2711 VDD2.n39 VDD2.n38 185
R2712 VDD2.n28 VDD2.n27 185
R2713 VDD2.n45 VDD2.n44 185
R2714 VDD2.n47 VDD2.n46 185
R2715 VDD2.n24 VDD2.n23 185
R2716 VDD2.n53 VDD2.n52 185
R2717 VDD2.n55 VDD2.n54 185
R2718 VDD2.n20 VDD2.n19 185
R2719 VDD2.n61 VDD2.n60 185
R2720 VDD2.n63 VDD2.n62 185
R2721 VDD2.n16 VDD2.n15 185
R2722 VDD2.n69 VDD2.n68 185
R2723 VDD2.n71 VDD2.n70 185
R2724 VDD2.n12 VDD2.n11 185
R2725 VDD2.n78 VDD2.n77 185
R2726 VDD2.n79 VDD2.n10 185
R2727 VDD2.n81 VDD2.n80 185
R2728 VDD2.n8 VDD2.n7 185
R2729 VDD2.n87 VDD2.n86 185
R2730 VDD2.n89 VDD2.n88 185
R2731 VDD2.n4 VDD2.n3 185
R2732 VDD2.n95 VDD2.n94 185
R2733 VDD2.n97 VDD2.n96 185
R2734 VDD2.n139 VDD2.t6 147.659
R2735 VDD2.n33 VDD2.t8 147.659
R2736 VDD2.n201 VDD2.n200 104.615
R2737 VDD2.n200 VDD2.n108 104.615
R2738 VDD2.n193 VDD2.n108 104.615
R2739 VDD2.n193 VDD2.n192 104.615
R2740 VDD2.n192 VDD2.n112 104.615
R2741 VDD2.n185 VDD2.n112 104.615
R2742 VDD2.n185 VDD2.n184 104.615
R2743 VDD2.n184 VDD2.n183 104.615
R2744 VDD2.n183 VDD2.n116 104.615
R2745 VDD2.n176 VDD2.n116 104.615
R2746 VDD2.n176 VDD2.n175 104.615
R2747 VDD2.n175 VDD2.n121 104.615
R2748 VDD2.n168 VDD2.n121 104.615
R2749 VDD2.n168 VDD2.n167 104.615
R2750 VDD2.n167 VDD2.n125 104.615
R2751 VDD2.n160 VDD2.n125 104.615
R2752 VDD2.n160 VDD2.n159 104.615
R2753 VDD2.n159 VDD2.n129 104.615
R2754 VDD2.n152 VDD2.n129 104.615
R2755 VDD2.n152 VDD2.n151 104.615
R2756 VDD2.n151 VDD2.n133 104.615
R2757 VDD2.n144 VDD2.n133 104.615
R2758 VDD2.n144 VDD2.n143 104.615
R2759 VDD2.n143 VDD2.n137 104.615
R2760 VDD2.n37 VDD2.n31 104.615
R2761 VDD2.n38 VDD2.n37 104.615
R2762 VDD2.n38 VDD2.n27 104.615
R2763 VDD2.n45 VDD2.n27 104.615
R2764 VDD2.n46 VDD2.n45 104.615
R2765 VDD2.n46 VDD2.n23 104.615
R2766 VDD2.n53 VDD2.n23 104.615
R2767 VDD2.n54 VDD2.n53 104.615
R2768 VDD2.n54 VDD2.n19 104.615
R2769 VDD2.n61 VDD2.n19 104.615
R2770 VDD2.n62 VDD2.n61 104.615
R2771 VDD2.n62 VDD2.n15 104.615
R2772 VDD2.n69 VDD2.n15 104.615
R2773 VDD2.n70 VDD2.n69 104.615
R2774 VDD2.n70 VDD2.n11 104.615
R2775 VDD2.n78 VDD2.n11 104.615
R2776 VDD2.n79 VDD2.n78 104.615
R2777 VDD2.n80 VDD2.n79 104.615
R2778 VDD2.n80 VDD2.n7 104.615
R2779 VDD2.n87 VDD2.n7 104.615
R2780 VDD2.n88 VDD2.n87 104.615
R2781 VDD2.n88 VDD2.n3 104.615
R2782 VDD2.n95 VDD2.n3 104.615
R2783 VDD2.n96 VDD2.n95 104.615
R2784 VDD2.n104 VDD2.n103 62.0152
R2785 VDD2 VDD2.n209 62.0123
R2786 VDD2.n208 VDD2.n207 60.6483
R2787 VDD2.n102 VDD2.n101 60.6481
R2788 VDD2.t6 VDD2.n137 52.3082
R2789 VDD2.t8 VDD2.n31 52.3082
R2790 VDD2.n102 VDD2.n100 50.7607
R2791 VDD2.n206 VDD2.n205 48.8641
R2792 VDD2.n206 VDD2.n104 48.4481
R2793 VDD2.n139 VDD2.n138 15.6677
R2794 VDD2.n33 VDD2.n32 15.6677
R2795 VDD2.n186 VDD2.n115 13.1884
R2796 VDD2.n81 VDD2.n10 13.1884
R2797 VDD2.n187 VDD2.n113 12.8005
R2798 VDD2.n182 VDD2.n117 12.8005
R2799 VDD2.n142 VDD2.n141 12.8005
R2800 VDD2.n36 VDD2.n35 12.8005
R2801 VDD2.n77 VDD2.n76 12.8005
R2802 VDD2.n82 VDD2.n8 12.8005
R2803 VDD2.n191 VDD2.n190 12.0247
R2804 VDD2.n181 VDD2.n118 12.0247
R2805 VDD2.n145 VDD2.n136 12.0247
R2806 VDD2.n39 VDD2.n30 12.0247
R2807 VDD2.n75 VDD2.n12 12.0247
R2808 VDD2.n86 VDD2.n85 12.0247
R2809 VDD2.n194 VDD2.n111 11.249
R2810 VDD2.n178 VDD2.n177 11.249
R2811 VDD2.n146 VDD2.n134 11.249
R2812 VDD2.n40 VDD2.n28 11.249
R2813 VDD2.n72 VDD2.n71 11.249
R2814 VDD2.n89 VDD2.n6 11.249
R2815 VDD2.n195 VDD2.n109 10.4732
R2816 VDD2.n174 VDD2.n120 10.4732
R2817 VDD2.n150 VDD2.n149 10.4732
R2818 VDD2.n44 VDD2.n43 10.4732
R2819 VDD2.n68 VDD2.n14 10.4732
R2820 VDD2.n90 VDD2.n4 10.4732
R2821 VDD2.n199 VDD2.n198 9.69747
R2822 VDD2.n173 VDD2.n122 9.69747
R2823 VDD2.n153 VDD2.n132 9.69747
R2824 VDD2.n47 VDD2.n26 9.69747
R2825 VDD2.n67 VDD2.n16 9.69747
R2826 VDD2.n94 VDD2.n93 9.69747
R2827 VDD2.n205 VDD2.n204 9.45567
R2828 VDD2.n100 VDD2.n99 9.45567
R2829 VDD2.n165 VDD2.n164 9.3005
R2830 VDD2.n124 VDD2.n123 9.3005
R2831 VDD2.n171 VDD2.n170 9.3005
R2832 VDD2.n173 VDD2.n172 9.3005
R2833 VDD2.n120 VDD2.n119 9.3005
R2834 VDD2.n179 VDD2.n178 9.3005
R2835 VDD2.n181 VDD2.n180 9.3005
R2836 VDD2.n117 VDD2.n114 9.3005
R2837 VDD2.n204 VDD2.n203 9.3005
R2838 VDD2.n107 VDD2.n106 9.3005
R2839 VDD2.n198 VDD2.n197 9.3005
R2840 VDD2.n196 VDD2.n195 9.3005
R2841 VDD2.n111 VDD2.n110 9.3005
R2842 VDD2.n190 VDD2.n189 9.3005
R2843 VDD2.n188 VDD2.n187 9.3005
R2844 VDD2.n163 VDD2.n162 9.3005
R2845 VDD2.n128 VDD2.n127 9.3005
R2846 VDD2.n157 VDD2.n156 9.3005
R2847 VDD2.n155 VDD2.n154 9.3005
R2848 VDD2.n132 VDD2.n131 9.3005
R2849 VDD2.n149 VDD2.n148 9.3005
R2850 VDD2.n147 VDD2.n146 9.3005
R2851 VDD2.n136 VDD2.n135 9.3005
R2852 VDD2.n141 VDD2.n140 9.3005
R2853 VDD2.n99 VDD2.n98 9.3005
R2854 VDD2.n2 VDD2.n1 9.3005
R2855 VDD2.n93 VDD2.n92 9.3005
R2856 VDD2.n91 VDD2.n90 9.3005
R2857 VDD2.n6 VDD2.n5 9.3005
R2858 VDD2.n85 VDD2.n84 9.3005
R2859 VDD2.n83 VDD2.n82 9.3005
R2860 VDD2.n22 VDD2.n21 9.3005
R2861 VDD2.n51 VDD2.n50 9.3005
R2862 VDD2.n49 VDD2.n48 9.3005
R2863 VDD2.n26 VDD2.n25 9.3005
R2864 VDD2.n43 VDD2.n42 9.3005
R2865 VDD2.n41 VDD2.n40 9.3005
R2866 VDD2.n30 VDD2.n29 9.3005
R2867 VDD2.n35 VDD2.n34 9.3005
R2868 VDD2.n57 VDD2.n56 9.3005
R2869 VDD2.n59 VDD2.n58 9.3005
R2870 VDD2.n18 VDD2.n17 9.3005
R2871 VDD2.n65 VDD2.n64 9.3005
R2872 VDD2.n67 VDD2.n66 9.3005
R2873 VDD2.n14 VDD2.n13 9.3005
R2874 VDD2.n73 VDD2.n72 9.3005
R2875 VDD2.n75 VDD2.n74 9.3005
R2876 VDD2.n76 VDD2.n9 9.3005
R2877 VDD2.n202 VDD2.n107 8.92171
R2878 VDD2.n170 VDD2.n169 8.92171
R2879 VDD2.n154 VDD2.n130 8.92171
R2880 VDD2.n48 VDD2.n24 8.92171
R2881 VDD2.n64 VDD2.n63 8.92171
R2882 VDD2.n97 VDD2.n2 8.92171
R2883 VDD2.n203 VDD2.n105 8.14595
R2884 VDD2.n166 VDD2.n124 8.14595
R2885 VDD2.n158 VDD2.n157 8.14595
R2886 VDD2.n52 VDD2.n51 8.14595
R2887 VDD2.n60 VDD2.n18 8.14595
R2888 VDD2.n98 VDD2.n0 8.14595
R2889 VDD2.n165 VDD2.n126 7.3702
R2890 VDD2.n161 VDD2.n128 7.3702
R2891 VDD2.n55 VDD2.n22 7.3702
R2892 VDD2.n59 VDD2.n20 7.3702
R2893 VDD2.n162 VDD2.n126 6.59444
R2894 VDD2.n162 VDD2.n161 6.59444
R2895 VDD2.n56 VDD2.n55 6.59444
R2896 VDD2.n56 VDD2.n20 6.59444
R2897 VDD2.n205 VDD2.n105 5.81868
R2898 VDD2.n166 VDD2.n165 5.81868
R2899 VDD2.n158 VDD2.n128 5.81868
R2900 VDD2.n52 VDD2.n22 5.81868
R2901 VDD2.n60 VDD2.n59 5.81868
R2902 VDD2.n100 VDD2.n0 5.81868
R2903 VDD2.n203 VDD2.n202 5.04292
R2904 VDD2.n169 VDD2.n124 5.04292
R2905 VDD2.n157 VDD2.n130 5.04292
R2906 VDD2.n51 VDD2.n24 5.04292
R2907 VDD2.n63 VDD2.n18 5.04292
R2908 VDD2.n98 VDD2.n97 5.04292
R2909 VDD2.n140 VDD2.n139 4.38563
R2910 VDD2.n34 VDD2.n33 4.38563
R2911 VDD2.n199 VDD2.n107 4.26717
R2912 VDD2.n170 VDD2.n122 4.26717
R2913 VDD2.n154 VDD2.n153 4.26717
R2914 VDD2.n48 VDD2.n47 4.26717
R2915 VDD2.n64 VDD2.n16 4.26717
R2916 VDD2.n94 VDD2.n2 4.26717
R2917 VDD2.n198 VDD2.n109 3.49141
R2918 VDD2.n174 VDD2.n173 3.49141
R2919 VDD2.n150 VDD2.n132 3.49141
R2920 VDD2.n44 VDD2.n26 3.49141
R2921 VDD2.n68 VDD2.n67 3.49141
R2922 VDD2.n93 VDD2.n4 3.49141
R2923 VDD2.n195 VDD2.n194 2.71565
R2924 VDD2.n177 VDD2.n120 2.71565
R2925 VDD2.n149 VDD2.n134 2.71565
R2926 VDD2.n43 VDD2.n28 2.71565
R2927 VDD2.n71 VDD2.n14 2.71565
R2928 VDD2.n90 VDD2.n89 2.71565
R2929 VDD2.n191 VDD2.n111 1.93989
R2930 VDD2.n178 VDD2.n118 1.93989
R2931 VDD2.n146 VDD2.n145 1.93989
R2932 VDD2.n40 VDD2.n39 1.93989
R2933 VDD2.n72 VDD2.n12 1.93989
R2934 VDD2.n86 VDD2.n6 1.93989
R2935 VDD2.n208 VDD2.n206 1.89705
R2936 VDD2.n190 VDD2.n113 1.16414
R2937 VDD2.n182 VDD2.n181 1.16414
R2938 VDD2.n142 VDD2.n136 1.16414
R2939 VDD2.n36 VDD2.n30 1.16414
R2940 VDD2.n77 VDD2.n75 1.16414
R2941 VDD2.n85 VDD2.n8 1.16414
R2942 VDD2.n209 VDD2.t5 1.08603
R2943 VDD2.n209 VDD2.t1 1.08603
R2944 VDD2.n207 VDD2.t7 1.08603
R2945 VDD2.n207 VDD2.t4 1.08603
R2946 VDD2.n103 VDD2.t3 1.08603
R2947 VDD2.n103 VDD2.t9 1.08603
R2948 VDD2.n101 VDD2.t0 1.08603
R2949 VDD2.n101 VDD2.t2 1.08603
R2950 VDD2 VDD2.n208 0.532828
R2951 VDD2.n104 VDD2.n102 0.419292
R2952 VDD2.n187 VDD2.n186 0.388379
R2953 VDD2.n117 VDD2.n115 0.388379
R2954 VDD2.n141 VDD2.n138 0.388379
R2955 VDD2.n35 VDD2.n32 0.388379
R2956 VDD2.n76 VDD2.n10 0.388379
R2957 VDD2.n82 VDD2.n81 0.388379
R2958 VDD2.n204 VDD2.n106 0.155672
R2959 VDD2.n197 VDD2.n106 0.155672
R2960 VDD2.n197 VDD2.n196 0.155672
R2961 VDD2.n196 VDD2.n110 0.155672
R2962 VDD2.n189 VDD2.n110 0.155672
R2963 VDD2.n189 VDD2.n188 0.155672
R2964 VDD2.n188 VDD2.n114 0.155672
R2965 VDD2.n180 VDD2.n114 0.155672
R2966 VDD2.n180 VDD2.n179 0.155672
R2967 VDD2.n179 VDD2.n119 0.155672
R2968 VDD2.n172 VDD2.n119 0.155672
R2969 VDD2.n172 VDD2.n171 0.155672
R2970 VDD2.n171 VDD2.n123 0.155672
R2971 VDD2.n164 VDD2.n123 0.155672
R2972 VDD2.n164 VDD2.n163 0.155672
R2973 VDD2.n163 VDD2.n127 0.155672
R2974 VDD2.n156 VDD2.n127 0.155672
R2975 VDD2.n156 VDD2.n155 0.155672
R2976 VDD2.n155 VDD2.n131 0.155672
R2977 VDD2.n148 VDD2.n131 0.155672
R2978 VDD2.n148 VDD2.n147 0.155672
R2979 VDD2.n147 VDD2.n135 0.155672
R2980 VDD2.n140 VDD2.n135 0.155672
R2981 VDD2.n34 VDD2.n29 0.155672
R2982 VDD2.n41 VDD2.n29 0.155672
R2983 VDD2.n42 VDD2.n41 0.155672
R2984 VDD2.n42 VDD2.n25 0.155672
R2985 VDD2.n49 VDD2.n25 0.155672
R2986 VDD2.n50 VDD2.n49 0.155672
R2987 VDD2.n50 VDD2.n21 0.155672
R2988 VDD2.n57 VDD2.n21 0.155672
R2989 VDD2.n58 VDD2.n57 0.155672
R2990 VDD2.n58 VDD2.n17 0.155672
R2991 VDD2.n65 VDD2.n17 0.155672
R2992 VDD2.n66 VDD2.n65 0.155672
R2993 VDD2.n66 VDD2.n13 0.155672
R2994 VDD2.n73 VDD2.n13 0.155672
R2995 VDD2.n74 VDD2.n73 0.155672
R2996 VDD2.n74 VDD2.n9 0.155672
R2997 VDD2.n83 VDD2.n9 0.155672
R2998 VDD2.n84 VDD2.n83 0.155672
R2999 VDD2.n84 VDD2.n5 0.155672
R3000 VDD2.n91 VDD2.n5 0.155672
R3001 VDD2.n92 VDD2.n91 0.155672
R3002 VDD2.n92 VDD2.n1 0.155672
R3003 VDD2.n99 VDD2.n1 0.155672
R3004 VP.n16 VP.t5 265.42
R3005 VP.n55 VP.t1 235.072
R3006 VP.n41 VP.t9 235.072
R3007 VP.n48 VP.t8 235.072
R3008 VP.n62 VP.t3 235.072
R3009 VP.n69 VP.t6 235.072
R3010 VP.n24 VP.t0 235.072
R3011 VP.n38 VP.t7 235.072
R3012 VP.n31 VP.t2 235.072
R3013 VP.n17 VP.t4 235.072
R3014 VP.n18 VP.n15 161.3
R3015 VP.n20 VP.n19 161.3
R3016 VP.n21 VP.n14 161.3
R3017 VP.n23 VP.n22 161.3
R3018 VP.n24 VP.n13 161.3
R3019 VP.n26 VP.n25 161.3
R3020 VP.n27 VP.n12 161.3
R3021 VP.n29 VP.n28 161.3
R3022 VP.n30 VP.n11 161.3
R3023 VP.n33 VP.n32 161.3
R3024 VP.n34 VP.n10 161.3
R3025 VP.n36 VP.n35 161.3
R3026 VP.n37 VP.n9 161.3
R3027 VP.n68 VP.n0 161.3
R3028 VP.n67 VP.n66 161.3
R3029 VP.n65 VP.n1 161.3
R3030 VP.n64 VP.n63 161.3
R3031 VP.n61 VP.n2 161.3
R3032 VP.n60 VP.n59 161.3
R3033 VP.n58 VP.n3 161.3
R3034 VP.n57 VP.n56 161.3
R3035 VP.n55 VP.n4 161.3
R3036 VP.n54 VP.n53 161.3
R3037 VP.n52 VP.n5 161.3
R3038 VP.n51 VP.n50 161.3
R3039 VP.n49 VP.n6 161.3
R3040 VP.n47 VP.n46 161.3
R3041 VP.n45 VP.n7 161.3
R3042 VP.n44 VP.n43 161.3
R3043 VP.n42 VP.n8 161.3
R3044 VP.n41 VP.n40 91.2348
R3045 VP.n70 VP.n69 91.2348
R3046 VP.n39 VP.n38 91.2348
R3047 VP.n17 VP.n16 60.1239
R3048 VP.n43 VP.n7 56.5617
R3049 VP.n67 VP.n1 56.5617
R3050 VP.n36 VP.n10 56.5617
R3051 VP.n40 VP.n39 53.8633
R3052 VP.n50 VP.n5 50.2647
R3053 VP.n60 VP.n3 50.2647
R3054 VP.n29 VP.n12 50.2647
R3055 VP.n19 VP.n14 50.2647
R3056 VP.n54 VP.n5 30.8893
R3057 VP.n56 VP.n3 30.8893
R3058 VP.n25 VP.n12 30.8893
R3059 VP.n23 VP.n14 30.8893
R3060 VP.n43 VP.n42 24.5923
R3061 VP.n47 VP.n7 24.5923
R3062 VP.n50 VP.n49 24.5923
R3063 VP.n55 VP.n54 24.5923
R3064 VP.n56 VP.n55 24.5923
R3065 VP.n61 VP.n60 24.5923
R3066 VP.n63 VP.n1 24.5923
R3067 VP.n68 VP.n67 24.5923
R3068 VP.n37 VP.n36 24.5923
R3069 VP.n30 VP.n29 24.5923
R3070 VP.n32 VP.n10 24.5923
R3071 VP.n24 VP.n23 24.5923
R3072 VP.n25 VP.n24 24.5923
R3073 VP.n19 VP.n18 24.5923
R3074 VP.n42 VP.n41 19.674
R3075 VP.n69 VP.n68 19.674
R3076 VP.n38 VP.n37 19.674
R3077 VP.n48 VP.n47 14.7556
R3078 VP.n63 VP.n62 14.7556
R3079 VP.n32 VP.n31 14.7556
R3080 VP.n16 VP.n15 13.3418
R3081 VP.n49 VP.n48 9.83723
R3082 VP.n62 VP.n61 9.83723
R3083 VP.n31 VP.n30 9.83723
R3084 VP.n18 VP.n17 9.83723
R3085 VP.n39 VP.n9 0.278335
R3086 VP.n40 VP.n8 0.278335
R3087 VP.n70 VP.n0 0.278335
R3088 VP.n20 VP.n15 0.189894
R3089 VP.n21 VP.n20 0.189894
R3090 VP.n22 VP.n21 0.189894
R3091 VP.n22 VP.n13 0.189894
R3092 VP.n26 VP.n13 0.189894
R3093 VP.n27 VP.n26 0.189894
R3094 VP.n28 VP.n27 0.189894
R3095 VP.n28 VP.n11 0.189894
R3096 VP.n33 VP.n11 0.189894
R3097 VP.n34 VP.n33 0.189894
R3098 VP.n35 VP.n34 0.189894
R3099 VP.n35 VP.n9 0.189894
R3100 VP.n44 VP.n8 0.189894
R3101 VP.n45 VP.n44 0.189894
R3102 VP.n46 VP.n45 0.189894
R3103 VP.n46 VP.n6 0.189894
R3104 VP.n51 VP.n6 0.189894
R3105 VP.n52 VP.n51 0.189894
R3106 VP.n53 VP.n52 0.189894
R3107 VP.n53 VP.n4 0.189894
R3108 VP.n57 VP.n4 0.189894
R3109 VP.n58 VP.n57 0.189894
R3110 VP.n59 VP.n58 0.189894
R3111 VP.n59 VP.n2 0.189894
R3112 VP.n64 VP.n2 0.189894
R3113 VP.n65 VP.n64 0.189894
R3114 VP.n66 VP.n65 0.189894
R3115 VP.n66 VP.n0 0.189894
R3116 VP VP.n70 0.153485
R3117 VDD1.n96 VDD1.n0 289.615
R3118 VDD1.n199 VDD1.n103 289.615
R3119 VDD1.n97 VDD1.n96 185
R3120 VDD1.n95 VDD1.n94 185
R3121 VDD1.n4 VDD1.n3 185
R3122 VDD1.n89 VDD1.n88 185
R3123 VDD1.n87 VDD1.n86 185
R3124 VDD1.n8 VDD1.n7 185
R3125 VDD1.n81 VDD1.n80 185
R3126 VDD1.n79 VDD1.n10 185
R3127 VDD1.n78 VDD1.n77 185
R3128 VDD1.n13 VDD1.n11 185
R3129 VDD1.n72 VDD1.n71 185
R3130 VDD1.n70 VDD1.n69 185
R3131 VDD1.n17 VDD1.n16 185
R3132 VDD1.n64 VDD1.n63 185
R3133 VDD1.n62 VDD1.n61 185
R3134 VDD1.n21 VDD1.n20 185
R3135 VDD1.n56 VDD1.n55 185
R3136 VDD1.n54 VDD1.n53 185
R3137 VDD1.n25 VDD1.n24 185
R3138 VDD1.n48 VDD1.n47 185
R3139 VDD1.n46 VDD1.n45 185
R3140 VDD1.n29 VDD1.n28 185
R3141 VDD1.n40 VDD1.n39 185
R3142 VDD1.n38 VDD1.n37 185
R3143 VDD1.n33 VDD1.n32 185
R3144 VDD1.n135 VDD1.n134 185
R3145 VDD1.n140 VDD1.n139 185
R3146 VDD1.n142 VDD1.n141 185
R3147 VDD1.n131 VDD1.n130 185
R3148 VDD1.n148 VDD1.n147 185
R3149 VDD1.n150 VDD1.n149 185
R3150 VDD1.n127 VDD1.n126 185
R3151 VDD1.n156 VDD1.n155 185
R3152 VDD1.n158 VDD1.n157 185
R3153 VDD1.n123 VDD1.n122 185
R3154 VDD1.n164 VDD1.n163 185
R3155 VDD1.n166 VDD1.n165 185
R3156 VDD1.n119 VDD1.n118 185
R3157 VDD1.n172 VDD1.n171 185
R3158 VDD1.n174 VDD1.n173 185
R3159 VDD1.n115 VDD1.n114 185
R3160 VDD1.n181 VDD1.n180 185
R3161 VDD1.n182 VDD1.n113 185
R3162 VDD1.n184 VDD1.n183 185
R3163 VDD1.n111 VDD1.n110 185
R3164 VDD1.n190 VDD1.n189 185
R3165 VDD1.n192 VDD1.n191 185
R3166 VDD1.n107 VDD1.n106 185
R3167 VDD1.n198 VDD1.n197 185
R3168 VDD1.n200 VDD1.n199 185
R3169 VDD1.n34 VDD1.t4 147.659
R3170 VDD1.n136 VDD1.t0 147.659
R3171 VDD1.n96 VDD1.n95 104.615
R3172 VDD1.n95 VDD1.n3 104.615
R3173 VDD1.n88 VDD1.n3 104.615
R3174 VDD1.n88 VDD1.n87 104.615
R3175 VDD1.n87 VDD1.n7 104.615
R3176 VDD1.n80 VDD1.n7 104.615
R3177 VDD1.n80 VDD1.n79 104.615
R3178 VDD1.n79 VDD1.n78 104.615
R3179 VDD1.n78 VDD1.n11 104.615
R3180 VDD1.n71 VDD1.n11 104.615
R3181 VDD1.n71 VDD1.n70 104.615
R3182 VDD1.n70 VDD1.n16 104.615
R3183 VDD1.n63 VDD1.n16 104.615
R3184 VDD1.n63 VDD1.n62 104.615
R3185 VDD1.n62 VDD1.n20 104.615
R3186 VDD1.n55 VDD1.n20 104.615
R3187 VDD1.n55 VDD1.n54 104.615
R3188 VDD1.n54 VDD1.n24 104.615
R3189 VDD1.n47 VDD1.n24 104.615
R3190 VDD1.n47 VDD1.n46 104.615
R3191 VDD1.n46 VDD1.n28 104.615
R3192 VDD1.n39 VDD1.n28 104.615
R3193 VDD1.n39 VDD1.n38 104.615
R3194 VDD1.n38 VDD1.n32 104.615
R3195 VDD1.n140 VDD1.n134 104.615
R3196 VDD1.n141 VDD1.n140 104.615
R3197 VDD1.n141 VDD1.n130 104.615
R3198 VDD1.n148 VDD1.n130 104.615
R3199 VDD1.n149 VDD1.n148 104.615
R3200 VDD1.n149 VDD1.n126 104.615
R3201 VDD1.n156 VDD1.n126 104.615
R3202 VDD1.n157 VDD1.n156 104.615
R3203 VDD1.n157 VDD1.n122 104.615
R3204 VDD1.n164 VDD1.n122 104.615
R3205 VDD1.n165 VDD1.n164 104.615
R3206 VDD1.n165 VDD1.n118 104.615
R3207 VDD1.n172 VDD1.n118 104.615
R3208 VDD1.n173 VDD1.n172 104.615
R3209 VDD1.n173 VDD1.n114 104.615
R3210 VDD1.n181 VDD1.n114 104.615
R3211 VDD1.n182 VDD1.n181 104.615
R3212 VDD1.n183 VDD1.n182 104.615
R3213 VDD1.n183 VDD1.n110 104.615
R3214 VDD1.n190 VDD1.n110 104.615
R3215 VDD1.n191 VDD1.n190 104.615
R3216 VDD1.n191 VDD1.n106 104.615
R3217 VDD1.n198 VDD1.n106 104.615
R3218 VDD1.n199 VDD1.n198 104.615
R3219 VDD1.n207 VDD1.n206 62.0152
R3220 VDD1.n102 VDD1.n101 60.6483
R3221 VDD1.n209 VDD1.n208 60.6481
R3222 VDD1.n205 VDD1.n204 60.6481
R3223 VDD1.t4 VDD1.n32 52.3082
R3224 VDD1.t0 VDD1.n134 52.3082
R3225 VDD1.n102 VDD1.n100 50.7607
R3226 VDD1.n205 VDD1.n203 50.7607
R3227 VDD1.n209 VDD1.n207 49.9793
R3228 VDD1.n34 VDD1.n33 15.6677
R3229 VDD1.n136 VDD1.n135 15.6677
R3230 VDD1.n81 VDD1.n10 13.1884
R3231 VDD1.n184 VDD1.n113 13.1884
R3232 VDD1.n82 VDD1.n8 12.8005
R3233 VDD1.n77 VDD1.n12 12.8005
R3234 VDD1.n37 VDD1.n36 12.8005
R3235 VDD1.n139 VDD1.n138 12.8005
R3236 VDD1.n180 VDD1.n179 12.8005
R3237 VDD1.n185 VDD1.n111 12.8005
R3238 VDD1.n86 VDD1.n85 12.0247
R3239 VDD1.n76 VDD1.n13 12.0247
R3240 VDD1.n40 VDD1.n31 12.0247
R3241 VDD1.n142 VDD1.n133 12.0247
R3242 VDD1.n178 VDD1.n115 12.0247
R3243 VDD1.n189 VDD1.n188 12.0247
R3244 VDD1.n89 VDD1.n6 11.249
R3245 VDD1.n73 VDD1.n72 11.249
R3246 VDD1.n41 VDD1.n29 11.249
R3247 VDD1.n143 VDD1.n131 11.249
R3248 VDD1.n175 VDD1.n174 11.249
R3249 VDD1.n192 VDD1.n109 11.249
R3250 VDD1.n90 VDD1.n4 10.4732
R3251 VDD1.n69 VDD1.n15 10.4732
R3252 VDD1.n45 VDD1.n44 10.4732
R3253 VDD1.n147 VDD1.n146 10.4732
R3254 VDD1.n171 VDD1.n117 10.4732
R3255 VDD1.n193 VDD1.n107 10.4732
R3256 VDD1.n94 VDD1.n93 9.69747
R3257 VDD1.n68 VDD1.n17 9.69747
R3258 VDD1.n48 VDD1.n27 9.69747
R3259 VDD1.n150 VDD1.n129 9.69747
R3260 VDD1.n170 VDD1.n119 9.69747
R3261 VDD1.n197 VDD1.n196 9.69747
R3262 VDD1.n100 VDD1.n99 9.45567
R3263 VDD1.n203 VDD1.n202 9.45567
R3264 VDD1.n60 VDD1.n59 9.3005
R3265 VDD1.n19 VDD1.n18 9.3005
R3266 VDD1.n66 VDD1.n65 9.3005
R3267 VDD1.n68 VDD1.n67 9.3005
R3268 VDD1.n15 VDD1.n14 9.3005
R3269 VDD1.n74 VDD1.n73 9.3005
R3270 VDD1.n76 VDD1.n75 9.3005
R3271 VDD1.n12 VDD1.n9 9.3005
R3272 VDD1.n99 VDD1.n98 9.3005
R3273 VDD1.n2 VDD1.n1 9.3005
R3274 VDD1.n93 VDD1.n92 9.3005
R3275 VDD1.n91 VDD1.n90 9.3005
R3276 VDD1.n6 VDD1.n5 9.3005
R3277 VDD1.n85 VDD1.n84 9.3005
R3278 VDD1.n83 VDD1.n82 9.3005
R3279 VDD1.n58 VDD1.n57 9.3005
R3280 VDD1.n23 VDD1.n22 9.3005
R3281 VDD1.n52 VDD1.n51 9.3005
R3282 VDD1.n50 VDD1.n49 9.3005
R3283 VDD1.n27 VDD1.n26 9.3005
R3284 VDD1.n44 VDD1.n43 9.3005
R3285 VDD1.n42 VDD1.n41 9.3005
R3286 VDD1.n31 VDD1.n30 9.3005
R3287 VDD1.n36 VDD1.n35 9.3005
R3288 VDD1.n202 VDD1.n201 9.3005
R3289 VDD1.n105 VDD1.n104 9.3005
R3290 VDD1.n196 VDD1.n195 9.3005
R3291 VDD1.n194 VDD1.n193 9.3005
R3292 VDD1.n109 VDD1.n108 9.3005
R3293 VDD1.n188 VDD1.n187 9.3005
R3294 VDD1.n186 VDD1.n185 9.3005
R3295 VDD1.n125 VDD1.n124 9.3005
R3296 VDD1.n154 VDD1.n153 9.3005
R3297 VDD1.n152 VDD1.n151 9.3005
R3298 VDD1.n129 VDD1.n128 9.3005
R3299 VDD1.n146 VDD1.n145 9.3005
R3300 VDD1.n144 VDD1.n143 9.3005
R3301 VDD1.n133 VDD1.n132 9.3005
R3302 VDD1.n138 VDD1.n137 9.3005
R3303 VDD1.n160 VDD1.n159 9.3005
R3304 VDD1.n162 VDD1.n161 9.3005
R3305 VDD1.n121 VDD1.n120 9.3005
R3306 VDD1.n168 VDD1.n167 9.3005
R3307 VDD1.n170 VDD1.n169 9.3005
R3308 VDD1.n117 VDD1.n116 9.3005
R3309 VDD1.n176 VDD1.n175 9.3005
R3310 VDD1.n178 VDD1.n177 9.3005
R3311 VDD1.n179 VDD1.n112 9.3005
R3312 VDD1.n97 VDD1.n2 8.92171
R3313 VDD1.n65 VDD1.n64 8.92171
R3314 VDD1.n49 VDD1.n25 8.92171
R3315 VDD1.n151 VDD1.n127 8.92171
R3316 VDD1.n167 VDD1.n166 8.92171
R3317 VDD1.n200 VDD1.n105 8.92171
R3318 VDD1.n98 VDD1.n0 8.14595
R3319 VDD1.n61 VDD1.n19 8.14595
R3320 VDD1.n53 VDD1.n52 8.14595
R3321 VDD1.n155 VDD1.n154 8.14595
R3322 VDD1.n163 VDD1.n121 8.14595
R3323 VDD1.n201 VDD1.n103 8.14595
R3324 VDD1.n60 VDD1.n21 7.3702
R3325 VDD1.n56 VDD1.n23 7.3702
R3326 VDD1.n158 VDD1.n125 7.3702
R3327 VDD1.n162 VDD1.n123 7.3702
R3328 VDD1.n57 VDD1.n21 6.59444
R3329 VDD1.n57 VDD1.n56 6.59444
R3330 VDD1.n159 VDD1.n158 6.59444
R3331 VDD1.n159 VDD1.n123 6.59444
R3332 VDD1.n100 VDD1.n0 5.81868
R3333 VDD1.n61 VDD1.n60 5.81868
R3334 VDD1.n53 VDD1.n23 5.81868
R3335 VDD1.n155 VDD1.n125 5.81868
R3336 VDD1.n163 VDD1.n162 5.81868
R3337 VDD1.n203 VDD1.n103 5.81868
R3338 VDD1.n98 VDD1.n97 5.04292
R3339 VDD1.n64 VDD1.n19 5.04292
R3340 VDD1.n52 VDD1.n25 5.04292
R3341 VDD1.n154 VDD1.n127 5.04292
R3342 VDD1.n166 VDD1.n121 5.04292
R3343 VDD1.n201 VDD1.n200 5.04292
R3344 VDD1.n35 VDD1.n34 4.38563
R3345 VDD1.n137 VDD1.n136 4.38563
R3346 VDD1.n94 VDD1.n2 4.26717
R3347 VDD1.n65 VDD1.n17 4.26717
R3348 VDD1.n49 VDD1.n48 4.26717
R3349 VDD1.n151 VDD1.n150 4.26717
R3350 VDD1.n167 VDD1.n119 4.26717
R3351 VDD1.n197 VDD1.n105 4.26717
R3352 VDD1.n93 VDD1.n4 3.49141
R3353 VDD1.n69 VDD1.n68 3.49141
R3354 VDD1.n45 VDD1.n27 3.49141
R3355 VDD1.n147 VDD1.n129 3.49141
R3356 VDD1.n171 VDD1.n170 3.49141
R3357 VDD1.n196 VDD1.n107 3.49141
R3358 VDD1.n90 VDD1.n89 2.71565
R3359 VDD1.n72 VDD1.n15 2.71565
R3360 VDD1.n44 VDD1.n29 2.71565
R3361 VDD1.n146 VDD1.n131 2.71565
R3362 VDD1.n174 VDD1.n117 2.71565
R3363 VDD1.n193 VDD1.n192 2.71565
R3364 VDD1.n86 VDD1.n6 1.93989
R3365 VDD1.n73 VDD1.n13 1.93989
R3366 VDD1.n41 VDD1.n40 1.93989
R3367 VDD1.n143 VDD1.n142 1.93989
R3368 VDD1.n175 VDD1.n115 1.93989
R3369 VDD1.n189 VDD1.n109 1.93989
R3370 VDD1 VDD1.n209 1.36472
R3371 VDD1.n85 VDD1.n8 1.16414
R3372 VDD1.n77 VDD1.n76 1.16414
R3373 VDD1.n37 VDD1.n31 1.16414
R3374 VDD1.n139 VDD1.n133 1.16414
R3375 VDD1.n180 VDD1.n178 1.16414
R3376 VDD1.n188 VDD1.n111 1.16414
R3377 VDD1.n208 VDD1.t7 1.08603
R3378 VDD1.n208 VDD1.t2 1.08603
R3379 VDD1.n101 VDD1.t5 1.08603
R3380 VDD1.n101 VDD1.t9 1.08603
R3381 VDD1.n206 VDD1.t6 1.08603
R3382 VDD1.n206 VDD1.t3 1.08603
R3383 VDD1.n204 VDD1.t1 1.08603
R3384 VDD1.n204 VDD1.t8 1.08603
R3385 VDD1 VDD1.n102 0.532828
R3386 VDD1.n207 VDD1.n205 0.419292
R3387 VDD1.n82 VDD1.n81 0.388379
R3388 VDD1.n12 VDD1.n10 0.388379
R3389 VDD1.n36 VDD1.n33 0.388379
R3390 VDD1.n138 VDD1.n135 0.388379
R3391 VDD1.n179 VDD1.n113 0.388379
R3392 VDD1.n185 VDD1.n184 0.388379
R3393 VDD1.n99 VDD1.n1 0.155672
R3394 VDD1.n92 VDD1.n1 0.155672
R3395 VDD1.n92 VDD1.n91 0.155672
R3396 VDD1.n91 VDD1.n5 0.155672
R3397 VDD1.n84 VDD1.n5 0.155672
R3398 VDD1.n84 VDD1.n83 0.155672
R3399 VDD1.n83 VDD1.n9 0.155672
R3400 VDD1.n75 VDD1.n9 0.155672
R3401 VDD1.n75 VDD1.n74 0.155672
R3402 VDD1.n74 VDD1.n14 0.155672
R3403 VDD1.n67 VDD1.n14 0.155672
R3404 VDD1.n67 VDD1.n66 0.155672
R3405 VDD1.n66 VDD1.n18 0.155672
R3406 VDD1.n59 VDD1.n18 0.155672
R3407 VDD1.n59 VDD1.n58 0.155672
R3408 VDD1.n58 VDD1.n22 0.155672
R3409 VDD1.n51 VDD1.n22 0.155672
R3410 VDD1.n51 VDD1.n50 0.155672
R3411 VDD1.n50 VDD1.n26 0.155672
R3412 VDD1.n43 VDD1.n26 0.155672
R3413 VDD1.n43 VDD1.n42 0.155672
R3414 VDD1.n42 VDD1.n30 0.155672
R3415 VDD1.n35 VDD1.n30 0.155672
R3416 VDD1.n137 VDD1.n132 0.155672
R3417 VDD1.n144 VDD1.n132 0.155672
R3418 VDD1.n145 VDD1.n144 0.155672
R3419 VDD1.n145 VDD1.n128 0.155672
R3420 VDD1.n152 VDD1.n128 0.155672
R3421 VDD1.n153 VDD1.n152 0.155672
R3422 VDD1.n153 VDD1.n124 0.155672
R3423 VDD1.n160 VDD1.n124 0.155672
R3424 VDD1.n161 VDD1.n160 0.155672
R3425 VDD1.n161 VDD1.n120 0.155672
R3426 VDD1.n168 VDD1.n120 0.155672
R3427 VDD1.n169 VDD1.n168 0.155672
R3428 VDD1.n169 VDD1.n116 0.155672
R3429 VDD1.n176 VDD1.n116 0.155672
R3430 VDD1.n177 VDD1.n176 0.155672
R3431 VDD1.n177 VDD1.n112 0.155672
R3432 VDD1.n186 VDD1.n112 0.155672
R3433 VDD1.n187 VDD1.n186 0.155672
R3434 VDD1.n187 VDD1.n108 0.155672
R3435 VDD1.n194 VDD1.n108 0.155672
R3436 VDD1.n195 VDD1.n194 0.155672
R3437 VDD1.n195 VDD1.n104 0.155672
R3438 VDD1.n202 VDD1.n104 0.155672
C0 VP VDD1 15.095599f
C1 VP VDD2 0.491485f
C2 VP VN 8.476139f
C3 VP VTAIL 14.8564f
C4 VDD1 VDD2 1.70069f
C5 VN VDD1 0.152047f
C6 VN VDD2 14.7615f
C7 VTAIL VDD1 13.9357f
C8 VTAIL VDD2 13.9788f
C9 VN VTAIL 14.841901f
C10 VDD2 B 7.446495f
C11 VDD1 B 7.430696f
C12 VTAIL B 10.06076f
C13 VN B 15.294451f
C14 VP B 13.575357f
C15 VDD1.n0 B 0.031231f
C16 VDD1.n1 B 0.022219f
C17 VDD1.n2 B 0.01194f
C18 VDD1.n3 B 0.028221f
C19 VDD1.n4 B 0.012642f
C20 VDD1.n5 B 0.022219f
C21 VDD1.n6 B 0.01194f
C22 VDD1.n7 B 0.028221f
C23 VDD1.n8 B 0.012642f
C24 VDD1.n9 B 0.022219f
C25 VDD1.n10 B 0.012291f
C26 VDD1.n11 B 0.028221f
C27 VDD1.n12 B 0.01194f
C28 VDD1.n13 B 0.012642f
C29 VDD1.n14 B 0.022219f
C30 VDD1.n15 B 0.01194f
C31 VDD1.n16 B 0.028221f
C32 VDD1.n17 B 0.012642f
C33 VDD1.n18 B 0.022219f
C34 VDD1.n19 B 0.01194f
C35 VDD1.n20 B 0.028221f
C36 VDD1.n21 B 0.012642f
C37 VDD1.n22 B 0.022219f
C38 VDD1.n23 B 0.01194f
C39 VDD1.n24 B 0.028221f
C40 VDD1.n25 B 0.012642f
C41 VDD1.n26 B 0.022219f
C42 VDD1.n27 B 0.01194f
C43 VDD1.n28 B 0.028221f
C44 VDD1.n29 B 0.012642f
C45 VDD1.n30 B 0.022219f
C46 VDD1.n31 B 0.01194f
C47 VDD1.n32 B 0.021166f
C48 VDD1.n33 B 0.016671f
C49 VDD1.t4 B 0.04678f
C50 VDD1.n34 B 0.162969f
C51 VDD1.n35 B 1.77556f
C52 VDD1.n36 B 0.01194f
C53 VDD1.n37 B 0.012642f
C54 VDD1.n38 B 0.028221f
C55 VDD1.n39 B 0.028221f
C56 VDD1.n40 B 0.012642f
C57 VDD1.n41 B 0.01194f
C58 VDD1.n42 B 0.022219f
C59 VDD1.n43 B 0.022219f
C60 VDD1.n44 B 0.01194f
C61 VDD1.n45 B 0.012642f
C62 VDD1.n46 B 0.028221f
C63 VDD1.n47 B 0.028221f
C64 VDD1.n48 B 0.012642f
C65 VDD1.n49 B 0.01194f
C66 VDD1.n50 B 0.022219f
C67 VDD1.n51 B 0.022219f
C68 VDD1.n52 B 0.01194f
C69 VDD1.n53 B 0.012642f
C70 VDD1.n54 B 0.028221f
C71 VDD1.n55 B 0.028221f
C72 VDD1.n56 B 0.012642f
C73 VDD1.n57 B 0.01194f
C74 VDD1.n58 B 0.022219f
C75 VDD1.n59 B 0.022219f
C76 VDD1.n60 B 0.01194f
C77 VDD1.n61 B 0.012642f
C78 VDD1.n62 B 0.028221f
C79 VDD1.n63 B 0.028221f
C80 VDD1.n64 B 0.012642f
C81 VDD1.n65 B 0.01194f
C82 VDD1.n66 B 0.022219f
C83 VDD1.n67 B 0.022219f
C84 VDD1.n68 B 0.01194f
C85 VDD1.n69 B 0.012642f
C86 VDD1.n70 B 0.028221f
C87 VDD1.n71 B 0.028221f
C88 VDD1.n72 B 0.012642f
C89 VDD1.n73 B 0.01194f
C90 VDD1.n74 B 0.022219f
C91 VDD1.n75 B 0.022219f
C92 VDD1.n76 B 0.01194f
C93 VDD1.n77 B 0.012642f
C94 VDD1.n78 B 0.028221f
C95 VDD1.n79 B 0.028221f
C96 VDD1.n80 B 0.028221f
C97 VDD1.n81 B 0.012291f
C98 VDD1.n82 B 0.01194f
C99 VDD1.n83 B 0.022219f
C100 VDD1.n84 B 0.022219f
C101 VDD1.n85 B 0.01194f
C102 VDD1.n86 B 0.012642f
C103 VDD1.n87 B 0.028221f
C104 VDD1.n88 B 0.028221f
C105 VDD1.n89 B 0.012642f
C106 VDD1.n90 B 0.01194f
C107 VDD1.n91 B 0.022219f
C108 VDD1.n92 B 0.022219f
C109 VDD1.n93 B 0.01194f
C110 VDD1.n94 B 0.012642f
C111 VDD1.n95 B 0.028221f
C112 VDD1.n96 B 0.061094f
C113 VDD1.n97 B 0.012642f
C114 VDD1.n98 B 0.01194f
C115 VDD1.n99 B 0.051359f
C116 VDD1.n100 B 0.056198f
C117 VDD1.t5 B 0.320265f
C118 VDD1.t9 B 0.320265f
C119 VDD1.n101 B 2.91884f
C120 VDD1.n102 B 0.530871f
C121 VDD1.n103 B 0.031231f
C122 VDD1.n104 B 0.022219f
C123 VDD1.n105 B 0.01194f
C124 VDD1.n106 B 0.028221f
C125 VDD1.n107 B 0.012642f
C126 VDD1.n108 B 0.022219f
C127 VDD1.n109 B 0.01194f
C128 VDD1.n110 B 0.028221f
C129 VDD1.n111 B 0.012642f
C130 VDD1.n112 B 0.022219f
C131 VDD1.n113 B 0.012291f
C132 VDD1.n114 B 0.028221f
C133 VDD1.n115 B 0.012642f
C134 VDD1.n116 B 0.022219f
C135 VDD1.n117 B 0.01194f
C136 VDD1.n118 B 0.028221f
C137 VDD1.n119 B 0.012642f
C138 VDD1.n120 B 0.022219f
C139 VDD1.n121 B 0.01194f
C140 VDD1.n122 B 0.028221f
C141 VDD1.n123 B 0.012642f
C142 VDD1.n124 B 0.022219f
C143 VDD1.n125 B 0.01194f
C144 VDD1.n126 B 0.028221f
C145 VDD1.n127 B 0.012642f
C146 VDD1.n128 B 0.022219f
C147 VDD1.n129 B 0.01194f
C148 VDD1.n130 B 0.028221f
C149 VDD1.n131 B 0.012642f
C150 VDD1.n132 B 0.022219f
C151 VDD1.n133 B 0.01194f
C152 VDD1.n134 B 0.021166f
C153 VDD1.n135 B 0.016671f
C154 VDD1.t0 B 0.04678f
C155 VDD1.n136 B 0.162969f
C156 VDD1.n137 B 1.77556f
C157 VDD1.n138 B 0.01194f
C158 VDD1.n139 B 0.012642f
C159 VDD1.n140 B 0.028221f
C160 VDD1.n141 B 0.028221f
C161 VDD1.n142 B 0.012642f
C162 VDD1.n143 B 0.01194f
C163 VDD1.n144 B 0.022219f
C164 VDD1.n145 B 0.022219f
C165 VDD1.n146 B 0.01194f
C166 VDD1.n147 B 0.012642f
C167 VDD1.n148 B 0.028221f
C168 VDD1.n149 B 0.028221f
C169 VDD1.n150 B 0.012642f
C170 VDD1.n151 B 0.01194f
C171 VDD1.n152 B 0.022219f
C172 VDD1.n153 B 0.022219f
C173 VDD1.n154 B 0.01194f
C174 VDD1.n155 B 0.012642f
C175 VDD1.n156 B 0.028221f
C176 VDD1.n157 B 0.028221f
C177 VDD1.n158 B 0.012642f
C178 VDD1.n159 B 0.01194f
C179 VDD1.n160 B 0.022219f
C180 VDD1.n161 B 0.022219f
C181 VDD1.n162 B 0.01194f
C182 VDD1.n163 B 0.012642f
C183 VDD1.n164 B 0.028221f
C184 VDD1.n165 B 0.028221f
C185 VDD1.n166 B 0.012642f
C186 VDD1.n167 B 0.01194f
C187 VDD1.n168 B 0.022219f
C188 VDD1.n169 B 0.022219f
C189 VDD1.n170 B 0.01194f
C190 VDD1.n171 B 0.012642f
C191 VDD1.n172 B 0.028221f
C192 VDD1.n173 B 0.028221f
C193 VDD1.n174 B 0.012642f
C194 VDD1.n175 B 0.01194f
C195 VDD1.n176 B 0.022219f
C196 VDD1.n177 B 0.022219f
C197 VDD1.n178 B 0.01194f
C198 VDD1.n179 B 0.01194f
C199 VDD1.n180 B 0.012642f
C200 VDD1.n181 B 0.028221f
C201 VDD1.n182 B 0.028221f
C202 VDD1.n183 B 0.028221f
C203 VDD1.n184 B 0.012291f
C204 VDD1.n185 B 0.01194f
C205 VDD1.n186 B 0.022219f
C206 VDD1.n187 B 0.022219f
C207 VDD1.n188 B 0.01194f
C208 VDD1.n189 B 0.012642f
C209 VDD1.n190 B 0.028221f
C210 VDD1.n191 B 0.028221f
C211 VDD1.n192 B 0.012642f
C212 VDD1.n193 B 0.01194f
C213 VDD1.n194 B 0.022219f
C214 VDD1.n195 B 0.022219f
C215 VDD1.n196 B 0.01194f
C216 VDD1.n197 B 0.012642f
C217 VDD1.n198 B 0.028221f
C218 VDD1.n199 B 0.061094f
C219 VDD1.n200 B 0.012642f
C220 VDD1.n201 B 0.01194f
C221 VDD1.n202 B 0.051359f
C222 VDD1.n203 B 0.056198f
C223 VDD1.t1 B 0.320265f
C224 VDD1.t8 B 0.320265f
C225 VDD1.n204 B 2.91883f
C226 VDD1.n205 B 0.523982f
C227 VDD1.t6 B 0.320265f
C228 VDD1.t3 B 0.320265f
C229 VDD1.n206 B 2.92826f
C230 VDD1.n207 B 2.6869f
C231 VDD1.t7 B 0.320265f
C232 VDD1.t2 B 0.320265f
C233 VDD1.n208 B 2.91883f
C234 VDD1.n209 B 2.97519f
C235 VP.n0 B 0.034033f
C236 VP.t6 B 2.42259f
C237 VP.n1 B 0.041098f
C238 VP.n2 B 0.025816f
C239 VP.t3 B 2.42259f
C240 VP.n3 B 0.02434f
C241 VP.n4 B 0.025816f
C242 VP.t1 B 2.42259f
C243 VP.n5 B 0.02434f
C244 VP.n6 B 0.025816f
C245 VP.t8 B 2.42259f
C246 VP.n7 B 0.041098f
C247 VP.n8 B 0.034033f
C248 VP.t9 B 2.42259f
C249 VP.n9 B 0.034033f
C250 VP.t7 B 2.42259f
C251 VP.n10 B 0.041098f
C252 VP.n11 B 0.025816f
C253 VP.t2 B 2.42259f
C254 VP.n12 B 0.02434f
C255 VP.n13 B 0.025816f
C256 VP.t0 B 2.42259f
C257 VP.n14 B 0.02434f
C258 VP.n15 B 0.190189f
C259 VP.t4 B 2.42259f
C260 VP.t5 B 2.53291f
C261 VP.n16 B 0.914437f
C262 VP.n17 B 0.90236f
C263 VP.n18 B 0.033693f
C264 VP.n19 B 0.047148f
C265 VP.n20 B 0.025816f
C266 VP.n21 B 0.025816f
C267 VP.n22 B 0.025816f
C268 VP.n23 B 0.051438f
C269 VP.n24 B 0.870436f
C270 VP.n25 B 0.051438f
C271 VP.n26 B 0.025816f
C272 VP.n27 B 0.025816f
C273 VP.n28 B 0.025816f
C274 VP.n29 B 0.047148f
C275 VP.n30 B 0.033693f
C276 VP.n31 B 0.846197f
C277 VP.n32 B 0.038419f
C278 VP.n33 B 0.025816f
C279 VP.n34 B 0.025816f
C280 VP.n35 B 0.025816f
C281 VP.n36 B 0.033956f
C282 VP.n37 B 0.043146f
C283 VP.n38 B 0.919498f
C284 VP.n39 B 1.5871f
C285 VP.n40 B 1.60438f
C286 VP.n41 B 0.919498f
C287 VP.n42 B 0.043146f
C288 VP.n43 B 0.033956f
C289 VP.n44 B 0.025816f
C290 VP.n45 B 0.025816f
C291 VP.n46 B 0.025816f
C292 VP.n47 B 0.038419f
C293 VP.n48 B 0.846197f
C294 VP.n49 B 0.033693f
C295 VP.n50 B 0.047148f
C296 VP.n51 B 0.025816f
C297 VP.n52 B 0.025816f
C298 VP.n53 B 0.025816f
C299 VP.n54 B 0.051438f
C300 VP.n55 B 0.870436f
C301 VP.n56 B 0.051438f
C302 VP.n57 B 0.025816f
C303 VP.n58 B 0.025816f
C304 VP.n59 B 0.025816f
C305 VP.n60 B 0.047148f
C306 VP.n61 B 0.033693f
C307 VP.n62 B 0.846197f
C308 VP.n63 B 0.038419f
C309 VP.n64 B 0.025816f
C310 VP.n65 B 0.025816f
C311 VP.n66 B 0.025816f
C312 VP.n67 B 0.033956f
C313 VP.n68 B 0.043146f
C314 VP.n69 B 0.919498f
C315 VP.n70 B 0.030934f
C316 VDD2.n0 B 0.031104f
C317 VDD2.n1 B 0.022129f
C318 VDD2.n2 B 0.011891f
C319 VDD2.n3 B 0.028106f
C320 VDD2.n4 B 0.01259f
C321 VDD2.n5 B 0.022129f
C322 VDD2.n6 B 0.011891f
C323 VDD2.n7 B 0.028106f
C324 VDD2.n8 B 0.01259f
C325 VDD2.n9 B 0.022129f
C326 VDD2.n10 B 0.012241f
C327 VDD2.n11 B 0.028106f
C328 VDD2.n12 B 0.01259f
C329 VDD2.n13 B 0.022129f
C330 VDD2.n14 B 0.011891f
C331 VDD2.n15 B 0.028106f
C332 VDD2.n16 B 0.01259f
C333 VDD2.n17 B 0.022129f
C334 VDD2.n18 B 0.011891f
C335 VDD2.n19 B 0.028106f
C336 VDD2.n20 B 0.01259f
C337 VDD2.n21 B 0.022129f
C338 VDD2.n22 B 0.011891f
C339 VDD2.n23 B 0.028106f
C340 VDD2.n24 B 0.01259f
C341 VDD2.n25 B 0.022129f
C342 VDD2.n26 B 0.011891f
C343 VDD2.n27 B 0.028106f
C344 VDD2.n28 B 0.01259f
C345 VDD2.n29 B 0.022129f
C346 VDD2.n30 B 0.011891f
C347 VDD2.n31 B 0.021079f
C348 VDD2.n32 B 0.016603f
C349 VDD2.t8 B 0.046589f
C350 VDD2.n33 B 0.162305f
C351 VDD2.n34 B 1.76832f
C352 VDD2.n35 B 0.011891f
C353 VDD2.n36 B 0.01259f
C354 VDD2.n37 B 0.028106f
C355 VDD2.n38 B 0.028106f
C356 VDD2.n39 B 0.01259f
C357 VDD2.n40 B 0.011891f
C358 VDD2.n41 B 0.022129f
C359 VDD2.n42 B 0.022129f
C360 VDD2.n43 B 0.011891f
C361 VDD2.n44 B 0.01259f
C362 VDD2.n45 B 0.028106f
C363 VDD2.n46 B 0.028106f
C364 VDD2.n47 B 0.01259f
C365 VDD2.n48 B 0.011891f
C366 VDD2.n49 B 0.022129f
C367 VDD2.n50 B 0.022129f
C368 VDD2.n51 B 0.011891f
C369 VDD2.n52 B 0.01259f
C370 VDD2.n53 B 0.028106f
C371 VDD2.n54 B 0.028106f
C372 VDD2.n55 B 0.01259f
C373 VDD2.n56 B 0.011891f
C374 VDD2.n57 B 0.022129f
C375 VDD2.n58 B 0.022129f
C376 VDD2.n59 B 0.011891f
C377 VDD2.n60 B 0.01259f
C378 VDD2.n61 B 0.028106f
C379 VDD2.n62 B 0.028106f
C380 VDD2.n63 B 0.01259f
C381 VDD2.n64 B 0.011891f
C382 VDD2.n65 B 0.022129f
C383 VDD2.n66 B 0.022129f
C384 VDD2.n67 B 0.011891f
C385 VDD2.n68 B 0.01259f
C386 VDD2.n69 B 0.028106f
C387 VDD2.n70 B 0.028106f
C388 VDD2.n71 B 0.01259f
C389 VDD2.n72 B 0.011891f
C390 VDD2.n73 B 0.022129f
C391 VDD2.n74 B 0.022129f
C392 VDD2.n75 B 0.011891f
C393 VDD2.n76 B 0.011891f
C394 VDD2.n77 B 0.01259f
C395 VDD2.n78 B 0.028106f
C396 VDD2.n79 B 0.028106f
C397 VDD2.n80 B 0.028106f
C398 VDD2.n81 B 0.012241f
C399 VDD2.n82 B 0.011891f
C400 VDD2.n83 B 0.022129f
C401 VDD2.n84 B 0.022129f
C402 VDD2.n85 B 0.011891f
C403 VDD2.n86 B 0.01259f
C404 VDD2.n87 B 0.028106f
C405 VDD2.n88 B 0.028106f
C406 VDD2.n89 B 0.01259f
C407 VDD2.n90 B 0.011891f
C408 VDD2.n91 B 0.022129f
C409 VDD2.n92 B 0.022129f
C410 VDD2.n93 B 0.011891f
C411 VDD2.n94 B 0.01259f
C412 VDD2.n95 B 0.028106f
C413 VDD2.n96 B 0.060845f
C414 VDD2.n97 B 0.01259f
C415 VDD2.n98 B 0.011891f
C416 VDD2.n99 B 0.05115f
C417 VDD2.n100 B 0.055969f
C418 VDD2.t0 B 0.318959f
C419 VDD2.t2 B 0.318959f
C420 VDD2.n101 B 2.90692f
C421 VDD2.n102 B 0.521845f
C422 VDD2.t3 B 0.318959f
C423 VDD2.t9 B 0.318959f
C424 VDD2.n103 B 2.91632f
C425 VDD2.n104 B 2.57953f
C426 VDD2.n105 B 0.031104f
C427 VDD2.n106 B 0.022129f
C428 VDD2.n107 B 0.011891f
C429 VDD2.n108 B 0.028106f
C430 VDD2.n109 B 0.01259f
C431 VDD2.n110 B 0.022129f
C432 VDD2.n111 B 0.011891f
C433 VDD2.n112 B 0.028106f
C434 VDD2.n113 B 0.01259f
C435 VDD2.n114 B 0.022129f
C436 VDD2.n115 B 0.012241f
C437 VDD2.n116 B 0.028106f
C438 VDD2.n117 B 0.011891f
C439 VDD2.n118 B 0.01259f
C440 VDD2.n119 B 0.022129f
C441 VDD2.n120 B 0.011891f
C442 VDD2.n121 B 0.028106f
C443 VDD2.n122 B 0.01259f
C444 VDD2.n123 B 0.022129f
C445 VDD2.n124 B 0.011891f
C446 VDD2.n125 B 0.028106f
C447 VDD2.n126 B 0.01259f
C448 VDD2.n127 B 0.022129f
C449 VDD2.n128 B 0.011891f
C450 VDD2.n129 B 0.028106f
C451 VDD2.n130 B 0.01259f
C452 VDD2.n131 B 0.022129f
C453 VDD2.n132 B 0.011891f
C454 VDD2.n133 B 0.028106f
C455 VDD2.n134 B 0.01259f
C456 VDD2.n135 B 0.022129f
C457 VDD2.n136 B 0.011891f
C458 VDD2.n137 B 0.021079f
C459 VDD2.n138 B 0.016603f
C460 VDD2.t6 B 0.046589f
C461 VDD2.n139 B 0.162305f
C462 VDD2.n140 B 1.76832f
C463 VDD2.n141 B 0.011891f
C464 VDD2.n142 B 0.01259f
C465 VDD2.n143 B 0.028106f
C466 VDD2.n144 B 0.028106f
C467 VDD2.n145 B 0.01259f
C468 VDD2.n146 B 0.011891f
C469 VDD2.n147 B 0.022129f
C470 VDD2.n148 B 0.022129f
C471 VDD2.n149 B 0.011891f
C472 VDD2.n150 B 0.01259f
C473 VDD2.n151 B 0.028106f
C474 VDD2.n152 B 0.028106f
C475 VDD2.n153 B 0.01259f
C476 VDD2.n154 B 0.011891f
C477 VDD2.n155 B 0.022129f
C478 VDD2.n156 B 0.022129f
C479 VDD2.n157 B 0.011891f
C480 VDD2.n158 B 0.01259f
C481 VDD2.n159 B 0.028106f
C482 VDD2.n160 B 0.028106f
C483 VDD2.n161 B 0.01259f
C484 VDD2.n162 B 0.011891f
C485 VDD2.n163 B 0.022129f
C486 VDD2.n164 B 0.022129f
C487 VDD2.n165 B 0.011891f
C488 VDD2.n166 B 0.01259f
C489 VDD2.n167 B 0.028106f
C490 VDD2.n168 B 0.028106f
C491 VDD2.n169 B 0.01259f
C492 VDD2.n170 B 0.011891f
C493 VDD2.n171 B 0.022129f
C494 VDD2.n172 B 0.022129f
C495 VDD2.n173 B 0.011891f
C496 VDD2.n174 B 0.01259f
C497 VDD2.n175 B 0.028106f
C498 VDD2.n176 B 0.028106f
C499 VDD2.n177 B 0.01259f
C500 VDD2.n178 B 0.011891f
C501 VDD2.n179 B 0.022129f
C502 VDD2.n180 B 0.022129f
C503 VDD2.n181 B 0.011891f
C504 VDD2.n182 B 0.01259f
C505 VDD2.n183 B 0.028106f
C506 VDD2.n184 B 0.028106f
C507 VDD2.n185 B 0.028106f
C508 VDD2.n186 B 0.012241f
C509 VDD2.n187 B 0.011891f
C510 VDD2.n188 B 0.022129f
C511 VDD2.n189 B 0.022129f
C512 VDD2.n190 B 0.011891f
C513 VDD2.n191 B 0.01259f
C514 VDD2.n192 B 0.028106f
C515 VDD2.n193 B 0.028106f
C516 VDD2.n194 B 0.01259f
C517 VDD2.n195 B 0.011891f
C518 VDD2.n196 B 0.022129f
C519 VDD2.n197 B 0.022129f
C520 VDD2.n198 B 0.011891f
C521 VDD2.n199 B 0.01259f
C522 VDD2.n200 B 0.028106f
C523 VDD2.n201 B 0.060845f
C524 VDD2.n202 B 0.01259f
C525 VDD2.n203 B 0.011891f
C526 VDD2.n204 B 0.05115f
C527 VDD2.n205 B 0.049324f
C528 VDD2.n206 B 2.72983f
C529 VDD2.t7 B 0.318959f
C530 VDD2.t4 B 0.318959f
C531 VDD2.n207 B 2.90693f
C532 VDD2.n208 B 0.357509f
C533 VDD2.t5 B 0.318959f
C534 VDD2.t1 B 0.318959f
C535 VDD2.n209 B 2.91629f
C536 VTAIL.t10 B 0.337823f
C537 VTAIL.t13 B 0.337823f
C538 VTAIL.n0 B 3.00648f
C539 VTAIL.n1 B 0.454653f
C540 VTAIL.n2 B 0.032943f
C541 VTAIL.n3 B 0.023438f
C542 VTAIL.n4 B 0.012594f
C543 VTAIL.n5 B 0.029768f
C544 VTAIL.n6 B 0.013335f
C545 VTAIL.n7 B 0.023438f
C546 VTAIL.n8 B 0.012594f
C547 VTAIL.n9 B 0.029768f
C548 VTAIL.n10 B 0.013335f
C549 VTAIL.n11 B 0.023438f
C550 VTAIL.n12 B 0.012965f
C551 VTAIL.n13 B 0.029768f
C552 VTAIL.n14 B 0.013335f
C553 VTAIL.n15 B 0.023438f
C554 VTAIL.n16 B 0.012594f
C555 VTAIL.n17 B 0.029768f
C556 VTAIL.n18 B 0.013335f
C557 VTAIL.n19 B 0.023438f
C558 VTAIL.n20 B 0.012594f
C559 VTAIL.n21 B 0.029768f
C560 VTAIL.n22 B 0.013335f
C561 VTAIL.n23 B 0.023438f
C562 VTAIL.n24 B 0.012594f
C563 VTAIL.n25 B 0.029768f
C564 VTAIL.n26 B 0.013335f
C565 VTAIL.n27 B 0.023438f
C566 VTAIL.n28 B 0.012594f
C567 VTAIL.n29 B 0.029768f
C568 VTAIL.n30 B 0.013335f
C569 VTAIL.n31 B 0.023438f
C570 VTAIL.n32 B 0.012594f
C571 VTAIL.n33 B 0.022326f
C572 VTAIL.n34 B 0.017585f
C573 VTAIL.t3 B 0.049345f
C574 VTAIL.n35 B 0.171903f
C575 VTAIL.n36 B 1.8729f
C576 VTAIL.n37 B 0.012594f
C577 VTAIL.n38 B 0.013335f
C578 VTAIL.n39 B 0.029768f
C579 VTAIL.n40 B 0.029768f
C580 VTAIL.n41 B 0.013335f
C581 VTAIL.n42 B 0.012594f
C582 VTAIL.n43 B 0.023438f
C583 VTAIL.n44 B 0.023438f
C584 VTAIL.n45 B 0.012594f
C585 VTAIL.n46 B 0.013335f
C586 VTAIL.n47 B 0.029768f
C587 VTAIL.n48 B 0.029768f
C588 VTAIL.n49 B 0.013335f
C589 VTAIL.n50 B 0.012594f
C590 VTAIL.n51 B 0.023438f
C591 VTAIL.n52 B 0.023438f
C592 VTAIL.n53 B 0.012594f
C593 VTAIL.n54 B 0.013335f
C594 VTAIL.n55 B 0.029768f
C595 VTAIL.n56 B 0.029768f
C596 VTAIL.n57 B 0.013335f
C597 VTAIL.n58 B 0.012594f
C598 VTAIL.n59 B 0.023438f
C599 VTAIL.n60 B 0.023438f
C600 VTAIL.n61 B 0.012594f
C601 VTAIL.n62 B 0.013335f
C602 VTAIL.n63 B 0.029768f
C603 VTAIL.n64 B 0.029768f
C604 VTAIL.n65 B 0.013335f
C605 VTAIL.n66 B 0.012594f
C606 VTAIL.n67 B 0.023438f
C607 VTAIL.n68 B 0.023438f
C608 VTAIL.n69 B 0.012594f
C609 VTAIL.n70 B 0.013335f
C610 VTAIL.n71 B 0.029768f
C611 VTAIL.n72 B 0.029768f
C612 VTAIL.n73 B 0.013335f
C613 VTAIL.n74 B 0.012594f
C614 VTAIL.n75 B 0.023438f
C615 VTAIL.n76 B 0.023438f
C616 VTAIL.n77 B 0.012594f
C617 VTAIL.n78 B 0.012594f
C618 VTAIL.n79 B 0.013335f
C619 VTAIL.n80 B 0.029768f
C620 VTAIL.n81 B 0.029768f
C621 VTAIL.n82 B 0.029768f
C622 VTAIL.n83 B 0.012965f
C623 VTAIL.n84 B 0.012594f
C624 VTAIL.n85 B 0.023438f
C625 VTAIL.n86 B 0.023438f
C626 VTAIL.n87 B 0.012594f
C627 VTAIL.n88 B 0.013335f
C628 VTAIL.n89 B 0.029768f
C629 VTAIL.n90 B 0.029768f
C630 VTAIL.n91 B 0.013335f
C631 VTAIL.n92 B 0.012594f
C632 VTAIL.n93 B 0.023438f
C633 VTAIL.n94 B 0.023438f
C634 VTAIL.n95 B 0.012594f
C635 VTAIL.n96 B 0.013335f
C636 VTAIL.n97 B 0.029768f
C637 VTAIL.n98 B 0.064443f
C638 VTAIL.n99 B 0.013335f
C639 VTAIL.n100 B 0.012594f
C640 VTAIL.n101 B 0.054175f
C641 VTAIL.n102 B 0.036059f
C642 VTAIL.n103 B 0.270342f
C643 VTAIL.t1 B 0.337823f
C644 VTAIL.t9 B 0.337823f
C645 VTAIL.n104 B 3.00648f
C646 VTAIL.n105 B 0.522198f
C647 VTAIL.t7 B 0.337823f
C648 VTAIL.t2 B 0.337823f
C649 VTAIL.n106 B 3.00648f
C650 VTAIL.n107 B 2.1713f
C651 VTAIL.t18 B 0.337823f
C652 VTAIL.t12 B 0.337823f
C653 VTAIL.n108 B 3.00649f
C654 VTAIL.n109 B 2.17128f
C655 VTAIL.t14 B 0.337823f
C656 VTAIL.t15 B 0.337823f
C657 VTAIL.n110 B 3.00649f
C658 VTAIL.n111 B 0.522185f
C659 VTAIL.n112 B 0.032943f
C660 VTAIL.n113 B 0.023438f
C661 VTAIL.n114 B 0.012594f
C662 VTAIL.n115 B 0.029768f
C663 VTAIL.n116 B 0.013335f
C664 VTAIL.n117 B 0.023438f
C665 VTAIL.n118 B 0.012594f
C666 VTAIL.n119 B 0.029768f
C667 VTAIL.n120 B 0.013335f
C668 VTAIL.n121 B 0.023438f
C669 VTAIL.n122 B 0.012965f
C670 VTAIL.n123 B 0.029768f
C671 VTAIL.n124 B 0.012594f
C672 VTAIL.n125 B 0.013335f
C673 VTAIL.n126 B 0.023438f
C674 VTAIL.n127 B 0.012594f
C675 VTAIL.n128 B 0.029768f
C676 VTAIL.n129 B 0.013335f
C677 VTAIL.n130 B 0.023438f
C678 VTAIL.n131 B 0.012594f
C679 VTAIL.n132 B 0.029768f
C680 VTAIL.n133 B 0.013335f
C681 VTAIL.n134 B 0.023438f
C682 VTAIL.n135 B 0.012594f
C683 VTAIL.n136 B 0.029768f
C684 VTAIL.n137 B 0.013335f
C685 VTAIL.n138 B 0.023438f
C686 VTAIL.n139 B 0.012594f
C687 VTAIL.n140 B 0.029768f
C688 VTAIL.n141 B 0.013335f
C689 VTAIL.n142 B 0.023438f
C690 VTAIL.n143 B 0.012594f
C691 VTAIL.n144 B 0.022326f
C692 VTAIL.n145 B 0.017585f
C693 VTAIL.t11 B 0.049345f
C694 VTAIL.n146 B 0.171903f
C695 VTAIL.n147 B 1.8729f
C696 VTAIL.n148 B 0.012594f
C697 VTAIL.n149 B 0.013335f
C698 VTAIL.n150 B 0.029768f
C699 VTAIL.n151 B 0.029768f
C700 VTAIL.n152 B 0.013335f
C701 VTAIL.n153 B 0.012594f
C702 VTAIL.n154 B 0.023438f
C703 VTAIL.n155 B 0.023438f
C704 VTAIL.n156 B 0.012594f
C705 VTAIL.n157 B 0.013335f
C706 VTAIL.n158 B 0.029768f
C707 VTAIL.n159 B 0.029768f
C708 VTAIL.n160 B 0.013335f
C709 VTAIL.n161 B 0.012594f
C710 VTAIL.n162 B 0.023438f
C711 VTAIL.n163 B 0.023438f
C712 VTAIL.n164 B 0.012594f
C713 VTAIL.n165 B 0.013335f
C714 VTAIL.n166 B 0.029768f
C715 VTAIL.n167 B 0.029768f
C716 VTAIL.n168 B 0.013335f
C717 VTAIL.n169 B 0.012594f
C718 VTAIL.n170 B 0.023438f
C719 VTAIL.n171 B 0.023438f
C720 VTAIL.n172 B 0.012594f
C721 VTAIL.n173 B 0.013335f
C722 VTAIL.n174 B 0.029768f
C723 VTAIL.n175 B 0.029768f
C724 VTAIL.n176 B 0.013335f
C725 VTAIL.n177 B 0.012594f
C726 VTAIL.n178 B 0.023438f
C727 VTAIL.n179 B 0.023438f
C728 VTAIL.n180 B 0.012594f
C729 VTAIL.n181 B 0.013335f
C730 VTAIL.n182 B 0.029768f
C731 VTAIL.n183 B 0.029768f
C732 VTAIL.n184 B 0.013335f
C733 VTAIL.n185 B 0.012594f
C734 VTAIL.n186 B 0.023438f
C735 VTAIL.n187 B 0.023438f
C736 VTAIL.n188 B 0.012594f
C737 VTAIL.n189 B 0.013335f
C738 VTAIL.n190 B 0.029768f
C739 VTAIL.n191 B 0.029768f
C740 VTAIL.n192 B 0.029768f
C741 VTAIL.n193 B 0.012965f
C742 VTAIL.n194 B 0.012594f
C743 VTAIL.n195 B 0.023438f
C744 VTAIL.n196 B 0.023438f
C745 VTAIL.n197 B 0.012594f
C746 VTAIL.n198 B 0.013335f
C747 VTAIL.n199 B 0.029768f
C748 VTAIL.n200 B 0.029768f
C749 VTAIL.n201 B 0.013335f
C750 VTAIL.n202 B 0.012594f
C751 VTAIL.n203 B 0.023438f
C752 VTAIL.n204 B 0.023438f
C753 VTAIL.n205 B 0.012594f
C754 VTAIL.n206 B 0.013335f
C755 VTAIL.n207 B 0.029768f
C756 VTAIL.n208 B 0.064443f
C757 VTAIL.n209 B 0.013335f
C758 VTAIL.n210 B 0.012594f
C759 VTAIL.n211 B 0.054175f
C760 VTAIL.n212 B 0.036059f
C761 VTAIL.n213 B 0.270342f
C762 VTAIL.t6 B 0.337823f
C763 VTAIL.t8 B 0.337823f
C764 VTAIL.n214 B 3.00649f
C765 VTAIL.n215 B 0.486052f
C766 VTAIL.t5 B 0.337823f
C767 VTAIL.t0 B 0.337823f
C768 VTAIL.n216 B 3.00649f
C769 VTAIL.n217 B 0.522185f
C770 VTAIL.n218 B 0.032943f
C771 VTAIL.n219 B 0.023438f
C772 VTAIL.n220 B 0.012594f
C773 VTAIL.n221 B 0.029768f
C774 VTAIL.n222 B 0.013335f
C775 VTAIL.n223 B 0.023438f
C776 VTAIL.n224 B 0.012594f
C777 VTAIL.n225 B 0.029768f
C778 VTAIL.n226 B 0.013335f
C779 VTAIL.n227 B 0.023438f
C780 VTAIL.n228 B 0.012965f
C781 VTAIL.n229 B 0.029768f
C782 VTAIL.n230 B 0.012594f
C783 VTAIL.n231 B 0.013335f
C784 VTAIL.n232 B 0.023438f
C785 VTAIL.n233 B 0.012594f
C786 VTAIL.n234 B 0.029768f
C787 VTAIL.n235 B 0.013335f
C788 VTAIL.n236 B 0.023438f
C789 VTAIL.n237 B 0.012594f
C790 VTAIL.n238 B 0.029768f
C791 VTAIL.n239 B 0.013335f
C792 VTAIL.n240 B 0.023438f
C793 VTAIL.n241 B 0.012594f
C794 VTAIL.n242 B 0.029768f
C795 VTAIL.n243 B 0.013335f
C796 VTAIL.n244 B 0.023438f
C797 VTAIL.n245 B 0.012594f
C798 VTAIL.n246 B 0.029768f
C799 VTAIL.n247 B 0.013335f
C800 VTAIL.n248 B 0.023438f
C801 VTAIL.n249 B 0.012594f
C802 VTAIL.n250 B 0.022326f
C803 VTAIL.n251 B 0.017585f
C804 VTAIL.t4 B 0.049345f
C805 VTAIL.n252 B 0.171903f
C806 VTAIL.n253 B 1.8729f
C807 VTAIL.n254 B 0.012594f
C808 VTAIL.n255 B 0.013335f
C809 VTAIL.n256 B 0.029768f
C810 VTAIL.n257 B 0.029768f
C811 VTAIL.n258 B 0.013335f
C812 VTAIL.n259 B 0.012594f
C813 VTAIL.n260 B 0.023438f
C814 VTAIL.n261 B 0.023438f
C815 VTAIL.n262 B 0.012594f
C816 VTAIL.n263 B 0.013335f
C817 VTAIL.n264 B 0.029768f
C818 VTAIL.n265 B 0.029768f
C819 VTAIL.n266 B 0.013335f
C820 VTAIL.n267 B 0.012594f
C821 VTAIL.n268 B 0.023438f
C822 VTAIL.n269 B 0.023438f
C823 VTAIL.n270 B 0.012594f
C824 VTAIL.n271 B 0.013335f
C825 VTAIL.n272 B 0.029768f
C826 VTAIL.n273 B 0.029768f
C827 VTAIL.n274 B 0.013335f
C828 VTAIL.n275 B 0.012594f
C829 VTAIL.n276 B 0.023438f
C830 VTAIL.n277 B 0.023438f
C831 VTAIL.n278 B 0.012594f
C832 VTAIL.n279 B 0.013335f
C833 VTAIL.n280 B 0.029768f
C834 VTAIL.n281 B 0.029768f
C835 VTAIL.n282 B 0.013335f
C836 VTAIL.n283 B 0.012594f
C837 VTAIL.n284 B 0.023438f
C838 VTAIL.n285 B 0.023438f
C839 VTAIL.n286 B 0.012594f
C840 VTAIL.n287 B 0.013335f
C841 VTAIL.n288 B 0.029768f
C842 VTAIL.n289 B 0.029768f
C843 VTAIL.n290 B 0.013335f
C844 VTAIL.n291 B 0.012594f
C845 VTAIL.n292 B 0.023438f
C846 VTAIL.n293 B 0.023438f
C847 VTAIL.n294 B 0.012594f
C848 VTAIL.n295 B 0.013335f
C849 VTAIL.n296 B 0.029768f
C850 VTAIL.n297 B 0.029768f
C851 VTAIL.n298 B 0.029768f
C852 VTAIL.n299 B 0.012965f
C853 VTAIL.n300 B 0.012594f
C854 VTAIL.n301 B 0.023438f
C855 VTAIL.n302 B 0.023438f
C856 VTAIL.n303 B 0.012594f
C857 VTAIL.n304 B 0.013335f
C858 VTAIL.n305 B 0.029768f
C859 VTAIL.n306 B 0.029768f
C860 VTAIL.n307 B 0.013335f
C861 VTAIL.n308 B 0.012594f
C862 VTAIL.n309 B 0.023438f
C863 VTAIL.n310 B 0.023438f
C864 VTAIL.n311 B 0.012594f
C865 VTAIL.n312 B 0.013335f
C866 VTAIL.n313 B 0.029768f
C867 VTAIL.n314 B 0.064443f
C868 VTAIL.n315 B 0.013335f
C869 VTAIL.n316 B 0.012594f
C870 VTAIL.n317 B 0.054175f
C871 VTAIL.n318 B 0.036059f
C872 VTAIL.n319 B 1.81234f
C873 VTAIL.n320 B 0.032943f
C874 VTAIL.n321 B 0.023438f
C875 VTAIL.n322 B 0.012594f
C876 VTAIL.n323 B 0.029768f
C877 VTAIL.n324 B 0.013335f
C878 VTAIL.n325 B 0.023438f
C879 VTAIL.n326 B 0.012594f
C880 VTAIL.n327 B 0.029768f
C881 VTAIL.n328 B 0.013335f
C882 VTAIL.n329 B 0.023438f
C883 VTAIL.n330 B 0.012965f
C884 VTAIL.n331 B 0.029768f
C885 VTAIL.n332 B 0.013335f
C886 VTAIL.n333 B 0.023438f
C887 VTAIL.n334 B 0.012594f
C888 VTAIL.n335 B 0.029768f
C889 VTAIL.n336 B 0.013335f
C890 VTAIL.n337 B 0.023438f
C891 VTAIL.n338 B 0.012594f
C892 VTAIL.n339 B 0.029768f
C893 VTAIL.n340 B 0.013335f
C894 VTAIL.n341 B 0.023438f
C895 VTAIL.n342 B 0.012594f
C896 VTAIL.n343 B 0.029768f
C897 VTAIL.n344 B 0.013335f
C898 VTAIL.n345 B 0.023438f
C899 VTAIL.n346 B 0.012594f
C900 VTAIL.n347 B 0.029768f
C901 VTAIL.n348 B 0.013335f
C902 VTAIL.n349 B 0.023438f
C903 VTAIL.n350 B 0.012594f
C904 VTAIL.n351 B 0.022326f
C905 VTAIL.n352 B 0.017585f
C906 VTAIL.t16 B 0.049345f
C907 VTAIL.n353 B 0.171903f
C908 VTAIL.n354 B 1.8729f
C909 VTAIL.n355 B 0.012594f
C910 VTAIL.n356 B 0.013335f
C911 VTAIL.n357 B 0.029768f
C912 VTAIL.n358 B 0.029768f
C913 VTAIL.n359 B 0.013335f
C914 VTAIL.n360 B 0.012594f
C915 VTAIL.n361 B 0.023438f
C916 VTAIL.n362 B 0.023438f
C917 VTAIL.n363 B 0.012594f
C918 VTAIL.n364 B 0.013335f
C919 VTAIL.n365 B 0.029768f
C920 VTAIL.n366 B 0.029768f
C921 VTAIL.n367 B 0.013335f
C922 VTAIL.n368 B 0.012594f
C923 VTAIL.n369 B 0.023438f
C924 VTAIL.n370 B 0.023438f
C925 VTAIL.n371 B 0.012594f
C926 VTAIL.n372 B 0.013335f
C927 VTAIL.n373 B 0.029768f
C928 VTAIL.n374 B 0.029768f
C929 VTAIL.n375 B 0.013335f
C930 VTAIL.n376 B 0.012594f
C931 VTAIL.n377 B 0.023438f
C932 VTAIL.n378 B 0.023438f
C933 VTAIL.n379 B 0.012594f
C934 VTAIL.n380 B 0.013335f
C935 VTAIL.n381 B 0.029768f
C936 VTAIL.n382 B 0.029768f
C937 VTAIL.n383 B 0.013335f
C938 VTAIL.n384 B 0.012594f
C939 VTAIL.n385 B 0.023438f
C940 VTAIL.n386 B 0.023438f
C941 VTAIL.n387 B 0.012594f
C942 VTAIL.n388 B 0.013335f
C943 VTAIL.n389 B 0.029768f
C944 VTAIL.n390 B 0.029768f
C945 VTAIL.n391 B 0.013335f
C946 VTAIL.n392 B 0.012594f
C947 VTAIL.n393 B 0.023438f
C948 VTAIL.n394 B 0.023438f
C949 VTAIL.n395 B 0.012594f
C950 VTAIL.n396 B 0.012594f
C951 VTAIL.n397 B 0.013335f
C952 VTAIL.n398 B 0.029768f
C953 VTAIL.n399 B 0.029768f
C954 VTAIL.n400 B 0.029768f
C955 VTAIL.n401 B 0.012965f
C956 VTAIL.n402 B 0.012594f
C957 VTAIL.n403 B 0.023438f
C958 VTAIL.n404 B 0.023438f
C959 VTAIL.n405 B 0.012594f
C960 VTAIL.n406 B 0.013335f
C961 VTAIL.n407 B 0.029768f
C962 VTAIL.n408 B 0.029768f
C963 VTAIL.n409 B 0.013335f
C964 VTAIL.n410 B 0.012594f
C965 VTAIL.n411 B 0.023438f
C966 VTAIL.n412 B 0.023438f
C967 VTAIL.n413 B 0.012594f
C968 VTAIL.n414 B 0.013335f
C969 VTAIL.n415 B 0.029768f
C970 VTAIL.n416 B 0.064443f
C971 VTAIL.n417 B 0.013335f
C972 VTAIL.n418 B 0.012594f
C973 VTAIL.n419 B 0.054175f
C974 VTAIL.n420 B 0.036059f
C975 VTAIL.n421 B 1.81234f
C976 VTAIL.t17 B 0.337823f
C977 VTAIL.t19 B 0.337823f
C978 VTAIL.n422 B 3.00648f
C979 VTAIL.n423 B 0.410382f
C980 VN.n0 B 0.033648f
C981 VN.t0 B 2.39517f
C982 VN.n1 B 0.040633f
C983 VN.n2 B 0.025523f
C984 VN.t6 B 2.39517f
C985 VN.n3 B 0.024065f
C986 VN.n4 B 0.025523f
C987 VN.t7 B 2.39517f
C988 VN.n5 B 0.024065f
C989 VN.n6 B 0.188035f
C990 VN.t9 B 2.39517f
C991 VN.t1 B 2.50423f
C992 VN.n7 B 0.904084f
C993 VN.n8 B 0.892144f
C994 VN.n9 B 0.033311f
C995 VN.n10 B 0.046615f
C996 VN.n11 B 0.025523f
C997 VN.n12 B 0.025523f
C998 VN.n13 B 0.025523f
C999 VN.n14 B 0.050856f
C1000 VN.n15 B 0.860581f
C1001 VN.n16 B 0.050856f
C1002 VN.n17 B 0.025523f
C1003 VN.n18 B 0.025523f
C1004 VN.n19 B 0.025523f
C1005 VN.n20 B 0.046615f
C1006 VN.n21 B 0.033311f
C1007 VN.n22 B 0.836616f
C1008 VN.n23 B 0.037984f
C1009 VN.n24 B 0.025523f
C1010 VN.n25 B 0.025523f
C1011 VN.n26 B 0.025523f
C1012 VN.n27 B 0.033571f
C1013 VN.n28 B 0.042658f
C1014 VN.n29 B 0.909088f
C1015 VN.n30 B 0.030584f
C1016 VN.n31 B 0.033648f
C1017 VN.t3 B 2.39517f
C1018 VN.n32 B 0.040633f
C1019 VN.n33 B 0.025523f
C1020 VN.t2 B 2.39517f
C1021 VN.n34 B 0.024065f
C1022 VN.n35 B 0.025523f
C1023 VN.t5 B 2.39517f
C1024 VN.n36 B 0.024065f
C1025 VN.n37 B 0.188035f
C1026 VN.t4 B 2.39517f
C1027 VN.t8 B 2.50423f
C1028 VN.n38 B 0.904084f
C1029 VN.n39 B 0.892144f
C1030 VN.n40 B 0.033311f
C1031 VN.n41 B 0.046615f
C1032 VN.n42 B 0.025523f
C1033 VN.n43 B 0.025523f
C1034 VN.n44 B 0.025523f
C1035 VN.n45 B 0.050856f
C1036 VN.n46 B 0.860581f
C1037 VN.n47 B 0.050856f
C1038 VN.n48 B 0.025523f
C1039 VN.n49 B 0.025523f
C1040 VN.n50 B 0.025523f
C1041 VN.n51 B 0.046615f
C1042 VN.n52 B 0.033311f
C1043 VN.n53 B 0.836616f
C1044 VN.n54 B 0.037984f
C1045 VN.n55 B 0.025523f
C1046 VN.n56 B 0.025523f
C1047 VN.n57 B 0.025523f
C1048 VN.n58 B 0.033571f
C1049 VN.n59 B 0.042658f
C1050 VN.n60 B 0.909088f
C1051 VN.n61 B 1.58269f
.ends

