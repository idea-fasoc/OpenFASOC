* NGSPICE file created from diff_pair_sample_1473.ext - technology: sky130A

.subckt diff_pair_sample_1473 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=2.925 pd=15.78 as=2.925 ps=15.78 w=7.5 l=0.82
X1 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=2.925 pd=15.78 as=0 ps=0 w=7.5 l=0.82
X2 VDD2.t1 VN.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.925 pd=15.78 as=2.925 ps=15.78 w=7.5 l=0.82
X3 VDD1.t0 VP.t1 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=2.925 pd=15.78 as=2.925 ps=15.78 w=7.5 l=0.82
X4 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=2.925 pd=15.78 as=0 ps=0 w=7.5 l=0.82
X5 B.t8 B.t6 B.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=2.925 pd=15.78 as=0 ps=0 w=7.5 l=0.82
X6 VDD2.t0 VN.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.925 pd=15.78 as=2.925 ps=15.78 w=7.5 l=0.82
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=2.925 pd=15.78 as=0 ps=0 w=7.5 l=0.82
R0 VP.n0 VP.t1 466.175
R1 VP.n0 VP.t0 429.634
R2 VP VP.n0 0.0516364
R3 VTAIL.n1 VTAIL.t0 51.4161
R4 VTAIL.n3 VTAIL.t1 51.4159
R5 VTAIL.n0 VTAIL.t2 51.4159
R6 VTAIL.n2 VTAIL.t3 51.4159
R7 VTAIL.n1 VTAIL.n0 20.8324
R8 VTAIL.n3 VTAIL.n2 19.841
R9 VTAIL.n2 VTAIL.n1 0.966017
R10 VTAIL VTAIL.n0 0.776362
R11 VTAIL VTAIL.n3 0.190155
R12 VDD1 VDD1.t1 100.993
R13 VDD1 VDD1.t0 68.4008
R14 B.n460 B.n459 585
R15 B.n196 B.n64 585
R16 B.n195 B.n194 585
R17 B.n193 B.n192 585
R18 B.n191 B.n190 585
R19 B.n189 B.n188 585
R20 B.n187 B.n186 585
R21 B.n185 B.n184 585
R22 B.n183 B.n182 585
R23 B.n181 B.n180 585
R24 B.n179 B.n178 585
R25 B.n177 B.n176 585
R26 B.n175 B.n174 585
R27 B.n173 B.n172 585
R28 B.n171 B.n170 585
R29 B.n169 B.n168 585
R30 B.n167 B.n166 585
R31 B.n165 B.n164 585
R32 B.n163 B.n162 585
R33 B.n161 B.n160 585
R34 B.n159 B.n158 585
R35 B.n157 B.n156 585
R36 B.n155 B.n154 585
R37 B.n153 B.n152 585
R38 B.n151 B.n150 585
R39 B.n149 B.n148 585
R40 B.n147 B.n146 585
R41 B.n145 B.n144 585
R42 B.n143 B.n142 585
R43 B.n141 B.n140 585
R44 B.n139 B.n138 585
R45 B.n137 B.n136 585
R46 B.n135 B.n134 585
R47 B.n133 B.n132 585
R48 B.n131 B.n130 585
R49 B.n129 B.n128 585
R50 B.n127 B.n126 585
R51 B.n125 B.n124 585
R52 B.n123 B.n122 585
R53 B.n121 B.n120 585
R54 B.n119 B.n118 585
R55 B.n117 B.n116 585
R56 B.n115 B.n114 585
R57 B.n113 B.n112 585
R58 B.n111 B.n110 585
R59 B.n109 B.n108 585
R60 B.n107 B.n106 585
R61 B.n105 B.n104 585
R62 B.n103 B.n102 585
R63 B.n101 B.n100 585
R64 B.n99 B.n98 585
R65 B.n97 B.n96 585
R66 B.n95 B.n94 585
R67 B.n93 B.n92 585
R68 B.n91 B.n90 585
R69 B.n89 B.n88 585
R70 B.n87 B.n86 585
R71 B.n85 B.n84 585
R72 B.n83 B.n82 585
R73 B.n81 B.n80 585
R74 B.n79 B.n78 585
R75 B.n77 B.n76 585
R76 B.n75 B.n74 585
R77 B.n73 B.n72 585
R78 B.n32 B.n31 585
R79 B.n465 B.n464 585
R80 B.n458 B.n65 585
R81 B.n65 B.n29 585
R82 B.n457 B.n28 585
R83 B.n469 B.n28 585
R84 B.n456 B.n27 585
R85 B.n470 B.n27 585
R86 B.n455 B.n26 585
R87 B.n471 B.n26 585
R88 B.n454 B.n453 585
R89 B.n453 B.n22 585
R90 B.n452 B.n21 585
R91 B.n477 B.n21 585
R92 B.n451 B.n20 585
R93 B.n478 B.n20 585
R94 B.n450 B.n19 585
R95 B.n479 B.n19 585
R96 B.n449 B.n448 585
R97 B.n448 B.n15 585
R98 B.n447 B.n14 585
R99 B.n485 B.n14 585
R100 B.n446 B.n13 585
R101 B.n486 B.n13 585
R102 B.n445 B.n12 585
R103 B.n487 B.n12 585
R104 B.n444 B.n443 585
R105 B.n443 B.n8 585
R106 B.n442 B.n7 585
R107 B.n493 B.n7 585
R108 B.n441 B.n6 585
R109 B.n494 B.n6 585
R110 B.n440 B.n5 585
R111 B.n495 B.n5 585
R112 B.n439 B.n438 585
R113 B.n438 B.n4 585
R114 B.n437 B.n197 585
R115 B.n437 B.n436 585
R116 B.n427 B.n198 585
R117 B.n199 B.n198 585
R118 B.n429 B.n428 585
R119 B.n430 B.n429 585
R120 B.n426 B.n204 585
R121 B.n204 B.n203 585
R122 B.n425 B.n424 585
R123 B.n424 B.n423 585
R124 B.n206 B.n205 585
R125 B.n207 B.n206 585
R126 B.n416 B.n415 585
R127 B.n417 B.n416 585
R128 B.n414 B.n212 585
R129 B.n212 B.n211 585
R130 B.n413 B.n412 585
R131 B.n412 B.n411 585
R132 B.n214 B.n213 585
R133 B.n215 B.n214 585
R134 B.n404 B.n403 585
R135 B.n405 B.n404 585
R136 B.n402 B.n220 585
R137 B.n220 B.n219 585
R138 B.n401 B.n400 585
R139 B.n400 B.n399 585
R140 B.n222 B.n221 585
R141 B.n223 B.n222 585
R142 B.n395 B.n394 585
R143 B.n226 B.n225 585
R144 B.n391 B.n390 585
R145 B.n392 B.n391 585
R146 B.n389 B.n259 585
R147 B.n388 B.n387 585
R148 B.n386 B.n385 585
R149 B.n384 B.n383 585
R150 B.n382 B.n381 585
R151 B.n380 B.n379 585
R152 B.n378 B.n377 585
R153 B.n376 B.n375 585
R154 B.n374 B.n373 585
R155 B.n372 B.n371 585
R156 B.n370 B.n369 585
R157 B.n368 B.n367 585
R158 B.n366 B.n365 585
R159 B.n364 B.n363 585
R160 B.n362 B.n361 585
R161 B.n360 B.n359 585
R162 B.n358 B.n357 585
R163 B.n356 B.n355 585
R164 B.n354 B.n353 585
R165 B.n352 B.n351 585
R166 B.n350 B.n349 585
R167 B.n348 B.n347 585
R168 B.n346 B.n345 585
R169 B.n344 B.n343 585
R170 B.n342 B.n341 585
R171 B.n339 B.n338 585
R172 B.n337 B.n336 585
R173 B.n335 B.n334 585
R174 B.n333 B.n332 585
R175 B.n331 B.n330 585
R176 B.n329 B.n328 585
R177 B.n327 B.n326 585
R178 B.n325 B.n324 585
R179 B.n323 B.n322 585
R180 B.n321 B.n320 585
R181 B.n318 B.n317 585
R182 B.n316 B.n315 585
R183 B.n314 B.n313 585
R184 B.n312 B.n311 585
R185 B.n310 B.n309 585
R186 B.n308 B.n307 585
R187 B.n306 B.n305 585
R188 B.n304 B.n303 585
R189 B.n302 B.n301 585
R190 B.n300 B.n299 585
R191 B.n298 B.n297 585
R192 B.n296 B.n295 585
R193 B.n294 B.n293 585
R194 B.n292 B.n291 585
R195 B.n290 B.n289 585
R196 B.n288 B.n287 585
R197 B.n286 B.n285 585
R198 B.n284 B.n283 585
R199 B.n282 B.n281 585
R200 B.n280 B.n279 585
R201 B.n278 B.n277 585
R202 B.n276 B.n275 585
R203 B.n274 B.n273 585
R204 B.n272 B.n271 585
R205 B.n270 B.n269 585
R206 B.n268 B.n267 585
R207 B.n266 B.n265 585
R208 B.n264 B.n258 585
R209 B.n392 B.n258 585
R210 B.n396 B.n224 585
R211 B.n224 B.n223 585
R212 B.n398 B.n397 585
R213 B.n399 B.n398 585
R214 B.n218 B.n217 585
R215 B.n219 B.n218 585
R216 B.n407 B.n406 585
R217 B.n406 B.n405 585
R218 B.n408 B.n216 585
R219 B.n216 B.n215 585
R220 B.n410 B.n409 585
R221 B.n411 B.n410 585
R222 B.n210 B.n209 585
R223 B.n211 B.n210 585
R224 B.n419 B.n418 585
R225 B.n418 B.n417 585
R226 B.n420 B.n208 585
R227 B.n208 B.n207 585
R228 B.n422 B.n421 585
R229 B.n423 B.n422 585
R230 B.n202 B.n201 585
R231 B.n203 B.n202 585
R232 B.n432 B.n431 585
R233 B.n431 B.n430 585
R234 B.n433 B.n200 585
R235 B.n200 B.n199 585
R236 B.n435 B.n434 585
R237 B.n436 B.n435 585
R238 B.n2 B.n0 585
R239 B.n4 B.n2 585
R240 B.n3 B.n1 585
R241 B.n494 B.n3 585
R242 B.n492 B.n491 585
R243 B.n493 B.n492 585
R244 B.n490 B.n9 585
R245 B.n9 B.n8 585
R246 B.n489 B.n488 585
R247 B.n488 B.n487 585
R248 B.n11 B.n10 585
R249 B.n486 B.n11 585
R250 B.n484 B.n483 585
R251 B.n485 B.n484 585
R252 B.n482 B.n16 585
R253 B.n16 B.n15 585
R254 B.n481 B.n480 585
R255 B.n480 B.n479 585
R256 B.n18 B.n17 585
R257 B.n478 B.n18 585
R258 B.n476 B.n475 585
R259 B.n477 B.n476 585
R260 B.n474 B.n23 585
R261 B.n23 B.n22 585
R262 B.n473 B.n472 585
R263 B.n472 B.n471 585
R264 B.n25 B.n24 585
R265 B.n470 B.n25 585
R266 B.n468 B.n467 585
R267 B.n469 B.n468 585
R268 B.n466 B.n30 585
R269 B.n30 B.n29 585
R270 B.n497 B.n496 585
R271 B.n496 B.n495 585
R272 B.n394 B.n224 516.524
R273 B.n464 B.n30 516.524
R274 B.n258 B.n222 516.524
R275 B.n460 B.n65 516.524
R276 B.n262 B.t13 422.087
R277 B.n260 B.t9 422.087
R278 B.n69 B.t6 422.087
R279 B.n66 B.t2 422.087
R280 B.n462 B.n461 256.663
R281 B.n462 B.n63 256.663
R282 B.n462 B.n62 256.663
R283 B.n462 B.n61 256.663
R284 B.n462 B.n60 256.663
R285 B.n462 B.n59 256.663
R286 B.n462 B.n58 256.663
R287 B.n462 B.n57 256.663
R288 B.n462 B.n56 256.663
R289 B.n462 B.n55 256.663
R290 B.n462 B.n54 256.663
R291 B.n462 B.n53 256.663
R292 B.n462 B.n52 256.663
R293 B.n462 B.n51 256.663
R294 B.n462 B.n50 256.663
R295 B.n462 B.n49 256.663
R296 B.n462 B.n48 256.663
R297 B.n462 B.n47 256.663
R298 B.n462 B.n46 256.663
R299 B.n462 B.n45 256.663
R300 B.n462 B.n44 256.663
R301 B.n462 B.n43 256.663
R302 B.n462 B.n42 256.663
R303 B.n462 B.n41 256.663
R304 B.n462 B.n40 256.663
R305 B.n462 B.n39 256.663
R306 B.n462 B.n38 256.663
R307 B.n462 B.n37 256.663
R308 B.n462 B.n36 256.663
R309 B.n462 B.n35 256.663
R310 B.n462 B.n34 256.663
R311 B.n462 B.n33 256.663
R312 B.n463 B.n462 256.663
R313 B.n393 B.n392 256.663
R314 B.n392 B.n227 256.663
R315 B.n392 B.n228 256.663
R316 B.n392 B.n229 256.663
R317 B.n392 B.n230 256.663
R318 B.n392 B.n231 256.663
R319 B.n392 B.n232 256.663
R320 B.n392 B.n233 256.663
R321 B.n392 B.n234 256.663
R322 B.n392 B.n235 256.663
R323 B.n392 B.n236 256.663
R324 B.n392 B.n237 256.663
R325 B.n392 B.n238 256.663
R326 B.n392 B.n239 256.663
R327 B.n392 B.n240 256.663
R328 B.n392 B.n241 256.663
R329 B.n392 B.n242 256.663
R330 B.n392 B.n243 256.663
R331 B.n392 B.n244 256.663
R332 B.n392 B.n245 256.663
R333 B.n392 B.n246 256.663
R334 B.n392 B.n247 256.663
R335 B.n392 B.n248 256.663
R336 B.n392 B.n249 256.663
R337 B.n392 B.n250 256.663
R338 B.n392 B.n251 256.663
R339 B.n392 B.n252 256.663
R340 B.n392 B.n253 256.663
R341 B.n392 B.n254 256.663
R342 B.n392 B.n255 256.663
R343 B.n392 B.n256 256.663
R344 B.n392 B.n257 256.663
R345 B.n398 B.n224 163.367
R346 B.n398 B.n218 163.367
R347 B.n406 B.n218 163.367
R348 B.n406 B.n216 163.367
R349 B.n410 B.n216 163.367
R350 B.n410 B.n210 163.367
R351 B.n418 B.n210 163.367
R352 B.n418 B.n208 163.367
R353 B.n422 B.n208 163.367
R354 B.n422 B.n202 163.367
R355 B.n431 B.n202 163.367
R356 B.n431 B.n200 163.367
R357 B.n435 B.n200 163.367
R358 B.n435 B.n2 163.367
R359 B.n496 B.n2 163.367
R360 B.n496 B.n3 163.367
R361 B.n492 B.n3 163.367
R362 B.n492 B.n9 163.367
R363 B.n488 B.n9 163.367
R364 B.n488 B.n11 163.367
R365 B.n484 B.n11 163.367
R366 B.n484 B.n16 163.367
R367 B.n480 B.n16 163.367
R368 B.n480 B.n18 163.367
R369 B.n476 B.n18 163.367
R370 B.n476 B.n23 163.367
R371 B.n472 B.n23 163.367
R372 B.n472 B.n25 163.367
R373 B.n468 B.n25 163.367
R374 B.n468 B.n30 163.367
R375 B.n391 B.n226 163.367
R376 B.n391 B.n259 163.367
R377 B.n387 B.n386 163.367
R378 B.n383 B.n382 163.367
R379 B.n379 B.n378 163.367
R380 B.n375 B.n374 163.367
R381 B.n371 B.n370 163.367
R382 B.n367 B.n366 163.367
R383 B.n363 B.n362 163.367
R384 B.n359 B.n358 163.367
R385 B.n355 B.n354 163.367
R386 B.n351 B.n350 163.367
R387 B.n347 B.n346 163.367
R388 B.n343 B.n342 163.367
R389 B.n338 B.n337 163.367
R390 B.n334 B.n333 163.367
R391 B.n330 B.n329 163.367
R392 B.n326 B.n325 163.367
R393 B.n322 B.n321 163.367
R394 B.n317 B.n316 163.367
R395 B.n313 B.n312 163.367
R396 B.n309 B.n308 163.367
R397 B.n305 B.n304 163.367
R398 B.n301 B.n300 163.367
R399 B.n297 B.n296 163.367
R400 B.n293 B.n292 163.367
R401 B.n289 B.n288 163.367
R402 B.n285 B.n284 163.367
R403 B.n281 B.n280 163.367
R404 B.n277 B.n276 163.367
R405 B.n273 B.n272 163.367
R406 B.n269 B.n268 163.367
R407 B.n265 B.n258 163.367
R408 B.n400 B.n222 163.367
R409 B.n400 B.n220 163.367
R410 B.n404 B.n220 163.367
R411 B.n404 B.n214 163.367
R412 B.n412 B.n214 163.367
R413 B.n412 B.n212 163.367
R414 B.n416 B.n212 163.367
R415 B.n416 B.n206 163.367
R416 B.n424 B.n206 163.367
R417 B.n424 B.n204 163.367
R418 B.n429 B.n204 163.367
R419 B.n429 B.n198 163.367
R420 B.n437 B.n198 163.367
R421 B.n438 B.n437 163.367
R422 B.n438 B.n5 163.367
R423 B.n6 B.n5 163.367
R424 B.n7 B.n6 163.367
R425 B.n443 B.n7 163.367
R426 B.n443 B.n12 163.367
R427 B.n13 B.n12 163.367
R428 B.n14 B.n13 163.367
R429 B.n448 B.n14 163.367
R430 B.n448 B.n19 163.367
R431 B.n20 B.n19 163.367
R432 B.n21 B.n20 163.367
R433 B.n453 B.n21 163.367
R434 B.n453 B.n26 163.367
R435 B.n27 B.n26 163.367
R436 B.n28 B.n27 163.367
R437 B.n65 B.n28 163.367
R438 B.n72 B.n32 163.367
R439 B.n76 B.n75 163.367
R440 B.n80 B.n79 163.367
R441 B.n84 B.n83 163.367
R442 B.n88 B.n87 163.367
R443 B.n92 B.n91 163.367
R444 B.n96 B.n95 163.367
R445 B.n100 B.n99 163.367
R446 B.n104 B.n103 163.367
R447 B.n108 B.n107 163.367
R448 B.n112 B.n111 163.367
R449 B.n116 B.n115 163.367
R450 B.n120 B.n119 163.367
R451 B.n124 B.n123 163.367
R452 B.n128 B.n127 163.367
R453 B.n132 B.n131 163.367
R454 B.n136 B.n135 163.367
R455 B.n140 B.n139 163.367
R456 B.n144 B.n143 163.367
R457 B.n148 B.n147 163.367
R458 B.n152 B.n151 163.367
R459 B.n156 B.n155 163.367
R460 B.n160 B.n159 163.367
R461 B.n164 B.n163 163.367
R462 B.n168 B.n167 163.367
R463 B.n172 B.n171 163.367
R464 B.n176 B.n175 163.367
R465 B.n180 B.n179 163.367
R466 B.n184 B.n183 163.367
R467 B.n188 B.n187 163.367
R468 B.n192 B.n191 163.367
R469 B.n194 B.n64 163.367
R470 B.n392 B.n223 98.8672
R471 B.n462 B.n29 98.8672
R472 B.n262 B.t15 91.4657
R473 B.n66 B.t4 91.4657
R474 B.n260 B.t12 91.457
R475 B.n69 B.t7 91.457
R476 B.n394 B.n393 71.676
R477 B.n259 B.n227 71.676
R478 B.n386 B.n228 71.676
R479 B.n382 B.n229 71.676
R480 B.n378 B.n230 71.676
R481 B.n374 B.n231 71.676
R482 B.n370 B.n232 71.676
R483 B.n366 B.n233 71.676
R484 B.n362 B.n234 71.676
R485 B.n358 B.n235 71.676
R486 B.n354 B.n236 71.676
R487 B.n350 B.n237 71.676
R488 B.n346 B.n238 71.676
R489 B.n342 B.n239 71.676
R490 B.n337 B.n240 71.676
R491 B.n333 B.n241 71.676
R492 B.n329 B.n242 71.676
R493 B.n325 B.n243 71.676
R494 B.n321 B.n244 71.676
R495 B.n316 B.n245 71.676
R496 B.n312 B.n246 71.676
R497 B.n308 B.n247 71.676
R498 B.n304 B.n248 71.676
R499 B.n300 B.n249 71.676
R500 B.n296 B.n250 71.676
R501 B.n292 B.n251 71.676
R502 B.n288 B.n252 71.676
R503 B.n284 B.n253 71.676
R504 B.n280 B.n254 71.676
R505 B.n276 B.n255 71.676
R506 B.n272 B.n256 71.676
R507 B.n268 B.n257 71.676
R508 B.n464 B.n463 71.676
R509 B.n72 B.n33 71.676
R510 B.n76 B.n34 71.676
R511 B.n80 B.n35 71.676
R512 B.n84 B.n36 71.676
R513 B.n88 B.n37 71.676
R514 B.n92 B.n38 71.676
R515 B.n96 B.n39 71.676
R516 B.n100 B.n40 71.676
R517 B.n104 B.n41 71.676
R518 B.n108 B.n42 71.676
R519 B.n112 B.n43 71.676
R520 B.n116 B.n44 71.676
R521 B.n120 B.n45 71.676
R522 B.n124 B.n46 71.676
R523 B.n128 B.n47 71.676
R524 B.n132 B.n48 71.676
R525 B.n136 B.n49 71.676
R526 B.n140 B.n50 71.676
R527 B.n144 B.n51 71.676
R528 B.n148 B.n52 71.676
R529 B.n152 B.n53 71.676
R530 B.n156 B.n54 71.676
R531 B.n160 B.n55 71.676
R532 B.n164 B.n56 71.676
R533 B.n168 B.n57 71.676
R534 B.n172 B.n58 71.676
R535 B.n176 B.n59 71.676
R536 B.n180 B.n60 71.676
R537 B.n184 B.n61 71.676
R538 B.n188 B.n62 71.676
R539 B.n192 B.n63 71.676
R540 B.n461 B.n64 71.676
R541 B.n461 B.n460 71.676
R542 B.n194 B.n63 71.676
R543 B.n191 B.n62 71.676
R544 B.n187 B.n61 71.676
R545 B.n183 B.n60 71.676
R546 B.n179 B.n59 71.676
R547 B.n175 B.n58 71.676
R548 B.n171 B.n57 71.676
R549 B.n167 B.n56 71.676
R550 B.n163 B.n55 71.676
R551 B.n159 B.n54 71.676
R552 B.n155 B.n53 71.676
R553 B.n151 B.n52 71.676
R554 B.n147 B.n51 71.676
R555 B.n143 B.n50 71.676
R556 B.n139 B.n49 71.676
R557 B.n135 B.n48 71.676
R558 B.n131 B.n47 71.676
R559 B.n127 B.n46 71.676
R560 B.n123 B.n45 71.676
R561 B.n119 B.n44 71.676
R562 B.n115 B.n43 71.676
R563 B.n111 B.n42 71.676
R564 B.n107 B.n41 71.676
R565 B.n103 B.n40 71.676
R566 B.n99 B.n39 71.676
R567 B.n95 B.n38 71.676
R568 B.n91 B.n37 71.676
R569 B.n87 B.n36 71.676
R570 B.n83 B.n35 71.676
R571 B.n79 B.n34 71.676
R572 B.n75 B.n33 71.676
R573 B.n463 B.n32 71.676
R574 B.n393 B.n226 71.676
R575 B.n387 B.n227 71.676
R576 B.n383 B.n228 71.676
R577 B.n379 B.n229 71.676
R578 B.n375 B.n230 71.676
R579 B.n371 B.n231 71.676
R580 B.n367 B.n232 71.676
R581 B.n363 B.n233 71.676
R582 B.n359 B.n234 71.676
R583 B.n355 B.n235 71.676
R584 B.n351 B.n236 71.676
R585 B.n347 B.n237 71.676
R586 B.n343 B.n238 71.676
R587 B.n338 B.n239 71.676
R588 B.n334 B.n240 71.676
R589 B.n330 B.n241 71.676
R590 B.n326 B.n242 71.676
R591 B.n322 B.n243 71.676
R592 B.n317 B.n244 71.676
R593 B.n313 B.n245 71.676
R594 B.n309 B.n246 71.676
R595 B.n305 B.n247 71.676
R596 B.n301 B.n248 71.676
R597 B.n297 B.n249 71.676
R598 B.n293 B.n250 71.676
R599 B.n289 B.n251 71.676
R600 B.n285 B.n252 71.676
R601 B.n281 B.n253 71.676
R602 B.n277 B.n254 71.676
R603 B.n273 B.n255 71.676
R604 B.n269 B.n256 71.676
R605 B.n265 B.n257 71.676
R606 B.n263 B.t14 69.1627
R607 B.n67 B.t5 69.1627
R608 B.n261 B.t11 69.1539
R609 B.n70 B.t8 69.1539
R610 B.n319 B.n263 59.5399
R611 B.n340 B.n261 59.5399
R612 B.n71 B.n70 59.5399
R613 B.n68 B.n67 59.5399
R614 B.n399 B.n223 58.4608
R615 B.n399 B.n219 58.4608
R616 B.n405 B.n219 58.4608
R617 B.n405 B.n215 58.4608
R618 B.n411 B.n215 58.4608
R619 B.n417 B.n211 58.4608
R620 B.n417 B.n207 58.4608
R621 B.n423 B.n207 58.4608
R622 B.n423 B.n203 58.4608
R623 B.n430 B.n203 58.4608
R624 B.n436 B.n199 58.4608
R625 B.n436 B.n4 58.4608
R626 B.n495 B.n4 58.4608
R627 B.n495 B.n494 58.4608
R628 B.n494 B.n493 58.4608
R629 B.n493 B.n8 58.4608
R630 B.n487 B.n486 58.4608
R631 B.n486 B.n485 58.4608
R632 B.n485 B.n15 58.4608
R633 B.n479 B.n15 58.4608
R634 B.n479 B.n478 58.4608
R635 B.n477 B.n22 58.4608
R636 B.n471 B.n22 58.4608
R637 B.n471 B.n470 58.4608
R638 B.n470 B.n469 58.4608
R639 B.n469 B.n29 58.4608
R640 B.t10 B.n211 51.5831
R641 B.n478 B.t3 51.5831
R642 B.n430 B.t0 41.2666
R643 B.n487 B.t1 41.2666
R644 B.n466 B.n465 33.5615
R645 B.n459 B.n458 33.5615
R646 B.n264 B.n221 33.5615
R647 B.n396 B.n395 33.5615
R648 B.n263 B.n262 22.3035
R649 B.n261 B.n260 22.3035
R650 B.n70 B.n69 22.3035
R651 B.n67 B.n66 22.3035
R652 B B.n497 18.0485
R653 B.t0 B.n199 17.1947
R654 B.t1 B.n8 17.1947
R655 B.n465 B.n31 10.6151
R656 B.n73 B.n31 10.6151
R657 B.n74 B.n73 10.6151
R658 B.n77 B.n74 10.6151
R659 B.n78 B.n77 10.6151
R660 B.n81 B.n78 10.6151
R661 B.n82 B.n81 10.6151
R662 B.n85 B.n82 10.6151
R663 B.n86 B.n85 10.6151
R664 B.n89 B.n86 10.6151
R665 B.n90 B.n89 10.6151
R666 B.n93 B.n90 10.6151
R667 B.n94 B.n93 10.6151
R668 B.n97 B.n94 10.6151
R669 B.n98 B.n97 10.6151
R670 B.n101 B.n98 10.6151
R671 B.n102 B.n101 10.6151
R672 B.n105 B.n102 10.6151
R673 B.n106 B.n105 10.6151
R674 B.n109 B.n106 10.6151
R675 B.n110 B.n109 10.6151
R676 B.n113 B.n110 10.6151
R677 B.n114 B.n113 10.6151
R678 B.n117 B.n114 10.6151
R679 B.n118 B.n117 10.6151
R680 B.n121 B.n118 10.6151
R681 B.n122 B.n121 10.6151
R682 B.n126 B.n125 10.6151
R683 B.n129 B.n126 10.6151
R684 B.n130 B.n129 10.6151
R685 B.n133 B.n130 10.6151
R686 B.n134 B.n133 10.6151
R687 B.n137 B.n134 10.6151
R688 B.n138 B.n137 10.6151
R689 B.n141 B.n138 10.6151
R690 B.n142 B.n141 10.6151
R691 B.n146 B.n145 10.6151
R692 B.n149 B.n146 10.6151
R693 B.n150 B.n149 10.6151
R694 B.n153 B.n150 10.6151
R695 B.n154 B.n153 10.6151
R696 B.n157 B.n154 10.6151
R697 B.n158 B.n157 10.6151
R698 B.n161 B.n158 10.6151
R699 B.n162 B.n161 10.6151
R700 B.n165 B.n162 10.6151
R701 B.n166 B.n165 10.6151
R702 B.n169 B.n166 10.6151
R703 B.n170 B.n169 10.6151
R704 B.n173 B.n170 10.6151
R705 B.n174 B.n173 10.6151
R706 B.n177 B.n174 10.6151
R707 B.n178 B.n177 10.6151
R708 B.n181 B.n178 10.6151
R709 B.n182 B.n181 10.6151
R710 B.n185 B.n182 10.6151
R711 B.n186 B.n185 10.6151
R712 B.n189 B.n186 10.6151
R713 B.n190 B.n189 10.6151
R714 B.n193 B.n190 10.6151
R715 B.n195 B.n193 10.6151
R716 B.n196 B.n195 10.6151
R717 B.n459 B.n196 10.6151
R718 B.n401 B.n221 10.6151
R719 B.n402 B.n401 10.6151
R720 B.n403 B.n402 10.6151
R721 B.n403 B.n213 10.6151
R722 B.n413 B.n213 10.6151
R723 B.n414 B.n413 10.6151
R724 B.n415 B.n414 10.6151
R725 B.n415 B.n205 10.6151
R726 B.n425 B.n205 10.6151
R727 B.n426 B.n425 10.6151
R728 B.n428 B.n426 10.6151
R729 B.n428 B.n427 10.6151
R730 B.n427 B.n197 10.6151
R731 B.n439 B.n197 10.6151
R732 B.n440 B.n439 10.6151
R733 B.n441 B.n440 10.6151
R734 B.n442 B.n441 10.6151
R735 B.n444 B.n442 10.6151
R736 B.n445 B.n444 10.6151
R737 B.n446 B.n445 10.6151
R738 B.n447 B.n446 10.6151
R739 B.n449 B.n447 10.6151
R740 B.n450 B.n449 10.6151
R741 B.n451 B.n450 10.6151
R742 B.n452 B.n451 10.6151
R743 B.n454 B.n452 10.6151
R744 B.n455 B.n454 10.6151
R745 B.n456 B.n455 10.6151
R746 B.n457 B.n456 10.6151
R747 B.n458 B.n457 10.6151
R748 B.n395 B.n225 10.6151
R749 B.n390 B.n225 10.6151
R750 B.n390 B.n389 10.6151
R751 B.n389 B.n388 10.6151
R752 B.n388 B.n385 10.6151
R753 B.n385 B.n384 10.6151
R754 B.n384 B.n381 10.6151
R755 B.n381 B.n380 10.6151
R756 B.n380 B.n377 10.6151
R757 B.n377 B.n376 10.6151
R758 B.n376 B.n373 10.6151
R759 B.n373 B.n372 10.6151
R760 B.n372 B.n369 10.6151
R761 B.n369 B.n368 10.6151
R762 B.n368 B.n365 10.6151
R763 B.n365 B.n364 10.6151
R764 B.n364 B.n361 10.6151
R765 B.n361 B.n360 10.6151
R766 B.n360 B.n357 10.6151
R767 B.n357 B.n356 10.6151
R768 B.n356 B.n353 10.6151
R769 B.n353 B.n352 10.6151
R770 B.n352 B.n349 10.6151
R771 B.n349 B.n348 10.6151
R772 B.n348 B.n345 10.6151
R773 B.n345 B.n344 10.6151
R774 B.n344 B.n341 10.6151
R775 B.n339 B.n336 10.6151
R776 B.n336 B.n335 10.6151
R777 B.n335 B.n332 10.6151
R778 B.n332 B.n331 10.6151
R779 B.n331 B.n328 10.6151
R780 B.n328 B.n327 10.6151
R781 B.n327 B.n324 10.6151
R782 B.n324 B.n323 10.6151
R783 B.n323 B.n320 10.6151
R784 B.n318 B.n315 10.6151
R785 B.n315 B.n314 10.6151
R786 B.n314 B.n311 10.6151
R787 B.n311 B.n310 10.6151
R788 B.n310 B.n307 10.6151
R789 B.n307 B.n306 10.6151
R790 B.n306 B.n303 10.6151
R791 B.n303 B.n302 10.6151
R792 B.n302 B.n299 10.6151
R793 B.n299 B.n298 10.6151
R794 B.n298 B.n295 10.6151
R795 B.n295 B.n294 10.6151
R796 B.n294 B.n291 10.6151
R797 B.n291 B.n290 10.6151
R798 B.n290 B.n287 10.6151
R799 B.n287 B.n286 10.6151
R800 B.n286 B.n283 10.6151
R801 B.n283 B.n282 10.6151
R802 B.n282 B.n279 10.6151
R803 B.n279 B.n278 10.6151
R804 B.n278 B.n275 10.6151
R805 B.n275 B.n274 10.6151
R806 B.n274 B.n271 10.6151
R807 B.n271 B.n270 10.6151
R808 B.n270 B.n267 10.6151
R809 B.n267 B.n266 10.6151
R810 B.n266 B.n264 10.6151
R811 B.n397 B.n396 10.6151
R812 B.n397 B.n217 10.6151
R813 B.n407 B.n217 10.6151
R814 B.n408 B.n407 10.6151
R815 B.n409 B.n408 10.6151
R816 B.n409 B.n209 10.6151
R817 B.n419 B.n209 10.6151
R818 B.n420 B.n419 10.6151
R819 B.n421 B.n420 10.6151
R820 B.n421 B.n201 10.6151
R821 B.n432 B.n201 10.6151
R822 B.n433 B.n432 10.6151
R823 B.n434 B.n433 10.6151
R824 B.n434 B.n0 10.6151
R825 B.n491 B.n1 10.6151
R826 B.n491 B.n490 10.6151
R827 B.n490 B.n489 10.6151
R828 B.n489 B.n10 10.6151
R829 B.n483 B.n10 10.6151
R830 B.n483 B.n482 10.6151
R831 B.n482 B.n481 10.6151
R832 B.n481 B.n17 10.6151
R833 B.n475 B.n17 10.6151
R834 B.n475 B.n474 10.6151
R835 B.n474 B.n473 10.6151
R836 B.n473 B.n24 10.6151
R837 B.n467 B.n24 10.6151
R838 B.n467 B.n466 10.6151
R839 B.n122 B.n71 8.74196
R840 B.n145 B.n68 8.74196
R841 B.n341 B.n340 8.74196
R842 B.n319 B.n318 8.74196
R843 B.n411 B.t10 6.87819
R844 B.t3 B.n477 6.87819
R845 B.n497 B.n0 2.81026
R846 B.n497 B.n1 2.81026
R847 B.n125 B.n71 1.87367
R848 B.n142 B.n68 1.87367
R849 B.n340 B.n339 1.87367
R850 B.n320 B.n319 1.87367
R851 VN VN.t0 466.555
R852 VN VN.t1 429.685
R853 VDD2.n0 VDD2.t0 100.219
R854 VDD2.n0 VDD2.t1 68.0947
R855 VDD2 VDD2.n0 0.306534
C0 VP VDD1 1.50596f
C1 VP VDD2 0.259664f
C2 VP VTAIL 1.12335f
C3 VDD1 VDD2 0.472666f
C4 VDD1 VTAIL 3.90311f
C5 VTAIL VDD2 3.94056f
C6 VN VP 3.78051f
C7 VN VDD1 0.148977f
C8 VN VDD2 1.39795f
C9 VN VTAIL 1.10895f
C10 VDD2 B 2.974867f
C11 VDD1 B 4.755401f
C12 VTAIL B 4.713236f
C13 VN B 6.3296f
C14 VP B 3.865474f
C15 VDD2.t0 B 1.24038f
C16 VDD2.t1 B 0.988916f
C17 VDD2.n0 B 1.63087f
C18 VN.t1 B 0.661973f
C19 VN.t0 B 0.758554f
C20 VDD1.t0 B 0.975616f
C21 VDD1.t1 B 1.23907f
C22 VTAIL.t2 B 1.03353f
C23 VTAIL.n0 B 0.933035f
C24 VTAIL.t0 B 1.03353f
C25 VTAIL.n1 B 0.943295f
C26 VTAIL.t3 B 1.03352f
C27 VTAIL.n2 B 0.889652f
C28 VTAIL.t1 B 1.03353f
C29 VTAIL.n3 B 0.847669f
C30 VP.t1 B 0.765082f
C31 VP.t0 B 0.669938f
C32 VP.n0 B 2.35121f
.ends

