* NGSPICE file created from diff_pair_sample_1018.ext - technology: sky130A

.subckt diff_pair_sample_1018 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t11 VN.t0 VDD2.t0 w_n2994_n1320# sky130_fd_pr__pfet_01v8 ad=0.2904 pd=2.09 as=0.2904 ps=2.09 w=1.76 l=2.2
X1 VDD1.t5 VP.t0 VTAIL.t4 w_n2994_n1320# sky130_fd_pr__pfet_01v8 ad=0.6864 pd=4.3 as=0.2904 ps=2.09 w=1.76 l=2.2
X2 VDD1.t4 VP.t1 VTAIL.t5 w_n2994_n1320# sky130_fd_pr__pfet_01v8 ad=0.2904 pd=2.09 as=0.6864 ps=4.3 w=1.76 l=2.2
X3 VTAIL.t0 VP.t2 VDD1.t3 w_n2994_n1320# sky130_fd_pr__pfet_01v8 ad=0.2904 pd=2.09 as=0.2904 ps=2.09 w=1.76 l=2.2
X4 VTAIL.t10 VN.t1 VDD2.t2 w_n2994_n1320# sky130_fd_pr__pfet_01v8 ad=0.2904 pd=2.09 as=0.2904 ps=2.09 w=1.76 l=2.2
X5 B.t11 B.t9 B.t10 w_n2994_n1320# sky130_fd_pr__pfet_01v8 ad=0.6864 pd=4.3 as=0 ps=0 w=1.76 l=2.2
X6 B.t8 B.t6 B.t7 w_n2994_n1320# sky130_fd_pr__pfet_01v8 ad=0.6864 pd=4.3 as=0 ps=0 w=1.76 l=2.2
X7 VDD2.t1 VN.t2 VTAIL.t9 w_n2994_n1320# sky130_fd_pr__pfet_01v8 ad=0.2904 pd=2.09 as=0.6864 ps=4.3 w=1.76 l=2.2
X8 B.t5 B.t3 B.t4 w_n2994_n1320# sky130_fd_pr__pfet_01v8 ad=0.6864 pd=4.3 as=0 ps=0 w=1.76 l=2.2
X9 VTAIL.t2 VP.t3 VDD1.t2 w_n2994_n1320# sky130_fd_pr__pfet_01v8 ad=0.2904 pd=2.09 as=0.2904 ps=2.09 w=1.76 l=2.2
X10 VDD2.t3 VN.t3 VTAIL.t8 w_n2994_n1320# sky130_fd_pr__pfet_01v8 ad=0.6864 pd=4.3 as=0.2904 ps=2.09 w=1.76 l=2.2
X11 VDD1.t1 VP.t4 VTAIL.t1 w_n2994_n1320# sky130_fd_pr__pfet_01v8 ad=0.6864 pd=4.3 as=0.2904 ps=2.09 w=1.76 l=2.2
X12 B.t2 B.t0 B.t1 w_n2994_n1320# sky130_fd_pr__pfet_01v8 ad=0.6864 pd=4.3 as=0 ps=0 w=1.76 l=2.2
X13 VDD2.t5 VN.t4 VTAIL.t7 w_n2994_n1320# sky130_fd_pr__pfet_01v8 ad=0.2904 pd=2.09 as=0.6864 ps=4.3 w=1.76 l=2.2
X14 VDD2.t4 VN.t5 VTAIL.t6 w_n2994_n1320# sky130_fd_pr__pfet_01v8 ad=0.6864 pd=4.3 as=0.2904 ps=2.09 w=1.76 l=2.2
X15 VDD1.t0 VP.t5 VTAIL.t3 w_n2994_n1320# sky130_fd_pr__pfet_01v8 ad=0.2904 pd=2.09 as=0.6864 ps=4.3 w=1.76 l=2.2
R0 VN.n25 VN.n14 161.3
R1 VN.n24 VN.n23 161.3
R2 VN.n22 VN.n15 161.3
R3 VN.n21 VN.n20 161.3
R4 VN.n19 VN.n16 161.3
R5 VN.n11 VN.n0 161.3
R6 VN.n10 VN.n9 161.3
R7 VN.n8 VN.n1 161.3
R8 VN.n7 VN.n6 161.3
R9 VN.n5 VN.n2 161.3
R10 VN.n13 VN.n12 97.1368
R11 VN.n27 VN.n26 97.1368
R12 VN.n4 VN.n3 59.4181
R13 VN.n18 VN.n17 59.4181
R14 VN.n3 VN.t5 51.7897
R15 VN.n17 VN.t2 51.7897
R16 VN.n10 VN.n1 42.0302
R17 VN.n24 VN.n15 42.0302
R18 VN VN.n27 39.608
R19 VN.n6 VN.n1 39.1239
R20 VN.n20 VN.n15 39.1239
R21 VN.n6 VN.n5 24.5923
R22 VN.n11 VN.n10 24.5923
R23 VN.n20 VN.n19 24.5923
R24 VN.n25 VN.n24 24.5923
R25 VN.n4 VN.t1 19.2805
R26 VN.n12 VN.t4 19.2805
R27 VN.n18 VN.t0 19.2805
R28 VN.n26 VN.t3 19.2805
R29 VN.n12 VN.n11 13.7719
R30 VN.n26 VN.n25 13.7719
R31 VN.n5 VN.n4 12.2964
R32 VN.n19 VN.n18 12.2964
R33 VN.n17 VN.n16 9.56133
R34 VN.n3 VN.n2 9.56133
R35 VN.n27 VN.n14 0.278335
R36 VN.n13 VN.n0 0.278335
R37 VN.n23 VN.n14 0.189894
R38 VN.n23 VN.n22 0.189894
R39 VN.n22 VN.n21 0.189894
R40 VN.n21 VN.n16 0.189894
R41 VN.n7 VN.n2 0.189894
R42 VN.n8 VN.n7 0.189894
R43 VN.n9 VN.n8 0.189894
R44 VN.n9 VN.n0 0.189894
R45 VN VN.n13 0.153485
R46 VDD2.n11 VDD2.n9 756.745
R47 VDD2.n2 VDD2.n0 756.745
R48 VDD2.n12 VDD2.n11 585
R49 VDD2.n3 VDD2.n2 585
R50 VDD2.t4 VDD2.n1 415.613
R51 VDD2.t3 VDD2.n10 415.613
R52 VDD2.n8 VDD2.n7 201.601
R53 VDD2 VDD2.n17 201.597
R54 VDD2.n11 VDD2.t3 85.8723
R55 VDD2.n2 VDD2.t4 85.8723
R56 VDD2.n8 VDD2.n6 51.9961
R57 VDD2.n16 VDD2.n15 50.4157
R58 VDD2.n16 VDD2.n8 32.3209
R59 VDD2.n17 VDD2.t0 18.4693
R60 VDD2.n17 VDD2.t1 18.4693
R61 VDD2.n7 VDD2.t2 18.4693
R62 VDD2.n7 VDD2.t5 18.4693
R63 VDD2.n12 VDD2.n10 14.9339
R64 VDD2.n3 VDD2.n1 14.9339
R65 VDD2.n13 VDD2.n9 12.8005
R66 VDD2.n4 VDD2.n0 12.8005
R67 VDD2.n15 VDD2.n14 9.45567
R68 VDD2.n6 VDD2.n5 9.45567
R69 VDD2.n14 VDD2.n13 9.3005
R70 VDD2.n5 VDD2.n4 9.3005
R71 VDD2.n14 VDD2.n10 5.44463
R72 VDD2.n5 VDD2.n1 5.44463
R73 VDD2 VDD2.n16 1.69447
R74 VDD2.n15 VDD2.n9 1.16414
R75 VDD2.n6 VDD2.n0 1.16414
R76 VDD2.n13 VDD2.n12 0.388379
R77 VDD2.n4 VDD2.n3 0.388379
R78 VTAIL.n34 VTAIL.n32 756.745
R79 VTAIL.n4 VTAIL.n2 756.745
R80 VTAIL.n26 VTAIL.n24 756.745
R81 VTAIL.n16 VTAIL.n14 756.745
R82 VTAIL.n35 VTAIL.n34 585
R83 VTAIL.n5 VTAIL.n4 585
R84 VTAIL.n27 VTAIL.n26 585
R85 VTAIL.n17 VTAIL.n16 585
R86 VTAIL.t7 VTAIL.n33 415.613
R87 VTAIL.t3 VTAIL.n3 415.613
R88 VTAIL.t5 VTAIL.n25 415.613
R89 VTAIL.t9 VTAIL.n15 415.613
R90 VTAIL.n23 VTAIL.n22 184.431
R91 VTAIL.n13 VTAIL.n12 184.431
R92 VTAIL.n1 VTAIL.n0 184.431
R93 VTAIL.n11 VTAIL.n10 184.431
R94 VTAIL.n34 VTAIL.t7 85.8723
R95 VTAIL.n4 VTAIL.t3 85.8723
R96 VTAIL.n26 VTAIL.t5 85.8723
R97 VTAIL.n16 VTAIL.t9 85.8723
R98 VTAIL.n39 VTAIL.n38 33.7369
R99 VTAIL.n9 VTAIL.n8 33.7369
R100 VTAIL.n31 VTAIL.n30 33.7369
R101 VTAIL.n21 VTAIL.n20 33.7369
R102 VTAIL.n0 VTAIL.t6 18.4693
R103 VTAIL.n0 VTAIL.t10 18.4693
R104 VTAIL.n10 VTAIL.t1 18.4693
R105 VTAIL.n10 VTAIL.t0 18.4693
R106 VTAIL.n22 VTAIL.t4 18.4693
R107 VTAIL.n22 VTAIL.t2 18.4693
R108 VTAIL.n12 VTAIL.t8 18.4693
R109 VTAIL.n12 VTAIL.t11 18.4693
R110 VTAIL.n13 VTAIL.n11 18.2462
R111 VTAIL.n39 VTAIL.n31 16.0652
R112 VTAIL.n35 VTAIL.n33 14.9339
R113 VTAIL.n5 VTAIL.n3 14.9339
R114 VTAIL.n27 VTAIL.n25 14.9339
R115 VTAIL.n17 VTAIL.n15 14.9339
R116 VTAIL.n36 VTAIL.n32 12.8005
R117 VTAIL.n6 VTAIL.n2 12.8005
R118 VTAIL.n28 VTAIL.n24 12.8005
R119 VTAIL.n18 VTAIL.n14 12.8005
R120 VTAIL.n38 VTAIL.n37 9.45567
R121 VTAIL.n8 VTAIL.n7 9.45567
R122 VTAIL.n30 VTAIL.n29 9.45567
R123 VTAIL.n20 VTAIL.n19 9.45567
R124 VTAIL.n37 VTAIL.n36 9.3005
R125 VTAIL.n7 VTAIL.n6 9.3005
R126 VTAIL.n29 VTAIL.n28 9.3005
R127 VTAIL.n19 VTAIL.n18 9.3005
R128 VTAIL.n37 VTAIL.n33 5.44463
R129 VTAIL.n7 VTAIL.n3 5.44463
R130 VTAIL.n29 VTAIL.n25 5.44463
R131 VTAIL.n19 VTAIL.n15 5.44463
R132 VTAIL.n21 VTAIL.n13 2.18153
R133 VTAIL.n31 VTAIL.n23 2.18153
R134 VTAIL.n11 VTAIL.n9 2.18153
R135 VTAIL VTAIL.n39 1.57809
R136 VTAIL.n23 VTAIL.n21 1.56084
R137 VTAIL.n9 VTAIL.n1 1.56084
R138 VTAIL.n38 VTAIL.n32 1.16414
R139 VTAIL.n8 VTAIL.n2 1.16414
R140 VTAIL.n30 VTAIL.n24 1.16414
R141 VTAIL.n20 VTAIL.n14 1.16414
R142 VTAIL VTAIL.n1 0.603948
R143 VTAIL.n36 VTAIL.n35 0.388379
R144 VTAIL.n6 VTAIL.n5 0.388379
R145 VTAIL.n28 VTAIL.n27 0.388379
R146 VTAIL.n18 VTAIL.n17 0.388379
R147 VP.n11 VP.n8 161.3
R148 VP.n13 VP.n12 161.3
R149 VP.n14 VP.n7 161.3
R150 VP.n16 VP.n15 161.3
R151 VP.n17 VP.n6 161.3
R152 VP.n36 VP.n0 161.3
R153 VP.n35 VP.n34 161.3
R154 VP.n33 VP.n1 161.3
R155 VP.n32 VP.n31 161.3
R156 VP.n30 VP.n2 161.3
R157 VP.n28 VP.n27 161.3
R158 VP.n26 VP.n3 161.3
R159 VP.n25 VP.n24 161.3
R160 VP.n23 VP.n4 161.3
R161 VP.n22 VP.n21 161.3
R162 VP.n20 VP.n5 97.1368
R163 VP.n38 VP.n37 97.1368
R164 VP.n19 VP.n18 97.1368
R165 VP.n10 VP.n9 59.4181
R166 VP.n9 VP.t0 51.7897
R167 VP.n24 VP.n23 42.0302
R168 VP.n35 VP.n1 42.0302
R169 VP.n16 VP.n7 42.0302
R170 VP.n20 VP.n19 39.3292
R171 VP.n24 VP.n3 39.1239
R172 VP.n31 VP.n1 39.1239
R173 VP.n12 VP.n7 39.1239
R174 VP.n23 VP.n22 24.5923
R175 VP.n28 VP.n3 24.5923
R176 VP.n31 VP.n30 24.5923
R177 VP.n36 VP.n35 24.5923
R178 VP.n17 VP.n16 24.5923
R179 VP.n12 VP.n11 24.5923
R180 VP.n5 VP.t4 19.2805
R181 VP.n29 VP.t2 19.2805
R182 VP.n37 VP.t5 19.2805
R183 VP.n18 VP.t1 19.2805
R184 VP.n10 VP.t3 19.2805
R185 VP.n22 VP.n5 13.7719
R186 VP.n37 VP.n36 13.7719
R187 VP.n18 VP.n17 13.7719
R188 VP.n29 VP.n28 12.2964
R189 VP.n30 VP.n29 12.2964
R190 VP.n11 VP.n10 12.2964
R191 VP.n9 VP.n8 9.56133
R192 VP.n19 VP.n6 0.278335
R193 VP.n21 VP.n20 0.278335
R194 VP.n38 VP.n0 0.278335
R195 VP.n13 VP.n8 0.189894
R196 VP.n14 VP.n13 0.189894
R197 VP.n15 VP.n14 0.189894
R198 VP.n15 VP.n6 0.189894
R199 VP.n21 VP.n4 0.189894
R200 VP.n25 VP.n4 0.189894
R201 VP.n26 VP.n25 0.189894
R202 VP.n27 VP.n26 0.189894
R203 VP.n27 VP.n2 0.189894
R204 VP.n32 VP.n2 0.189894
R205 VP.n33 VP.n32 0.189894
R206 VP.n34 VP.n33 0.189894
R207 VP.n34 VP.n0 0.189894
R208 VP VP.n38 0.153485
R209 VDD1.n2 VDD1.n0 756.745
R210 VDD1.n9 VDD1.n7 756.745
R211 VDD1.n3 VDD1.n2 585
R212 VDD1.n10 VDD1.n9 585
R213 VDD1.t1 VDD1.n8 415.613
R214 VDD1.t5 VDD1.n1 415.613
R215 VDD1.n15 VDD1.n14 201.601
R216 VDD1.n17 VDD1.n16 201.111
R217 VDD1.n2 VDD1.t5 85.8723
R218 VDD1.n9 VDD1.t1 85.8723
R219 VDD1 VDD1.n6 52.1096
R220 VDD1.n15 VDD1.n13 51.9961
R221 VDD1.n17 VDD1.n15 33.9944
R222 VDD1.n16 VDD1.t2 18.4693
R223 VDD1.n16 VDD1.t4 18.4693
R224 VDD1.n14 VDD1.t3 18.4693
R225 VDD1.n14 VDD1.t0 18.4693
R226 VDD1.n3 VDD1.n1 14.9339
R227 VDD1.n10 VDD1.n8 14.9339
R228 VDD1.n4 VDD1.n0 12.8005
R229 VDD1.n11 VDD1.n7 12.8005
R230 VDD1.n6 VDD1.n5 9.45567
R231 VDD1.n13 VDD1.n12 9.45567
R232 VDD1.n5 VDD1.n4 9.3005
R233 VDD1.n12 VDD1.n11 9.3005
R234 VDD1.n5 VDD1.n1 5.44463
R235 VDD1.n12 VDD1.n8 5.44463
R236 VDD1.n6 VDD1.n0 1.16414
R237 VDD1.n13 VDD1.n7 1.16414
R238 VDD1 VDD1.n17 0.487569
R239 VDD1.n4 VDD1.n3 0.388379
R240 VDD1.n11 VDD1.n10 0.388379
R241 B.n342 B.n41 585
R242 B.n344 B.n343 585
R243 B.n345 B.n40 585
R244 B.n347 B.n346 585
R245 B.n348 B.n39 585
R246 B.n350 B.n349 585
R247 B.n351 B.n38 585
R248 B.n353 B.n352 585
R249 B.n354 B.n37 585
R250 B.n356 B.n355 585
R251 B.n357 B.n36 585
R252 B.n359 B.n358 585
R253 B.n361 B.n33 585
R254 B.n363 B.n362 585
R255 B.n364 B.n32 585
R256 B.n366 B.n365 585
R257 B.n367 B.n31 585
R258 B.n369 B.n368 585
R259 B.n370 B.n30 585
R260 B.n372 B.n371 585
R261 B.n373 B.n27 585
R262 B.n376 B.n375 585
R263 B.n377 B.n26 585
R264 B.n379 B.n378 585
R265 B.n380 B.n25 585
R266 B.n382 B.n381 585
R267 B.n383 B.n24 585
R268 B.n385 B.n384 585
R269 B.n386 B.n23 585
R270 B.n388 B.n387 585
R271 B.n389 B.n22 585
R272 B.n391 B.n390 585
R273 B.n392 B.n21 585
R274 B.n341 B.n340 585
R275 B.n339 B.n42 585
R276 B.n338 B.n337 585
R277 B.n336 B.n43 585
R278 B.n335 B.n334 585
R279 B.n333 B.n44 585
R280 B.n332 B.n331 585
R281 B.n330 B.n45 585
R282 B.n329 B.n328 585
R283 B.n327 B.n46 585
R284 B.n326 B.n325 585
R285 B.n324 B.n47 585
R286 B.n323 B.n322 585
R287 B.n321 B.n48 585
R288 B.n320 B.n319 585
R289 B.n318 B.n49 585
R290 B.n317 B.n316 585
R291 B.n315 B.n50 585
R292 B.n314 B.n313 585
R293 B.n312 B.n51 585
R294 B.n311 B.n310 585
R295 B.n309 B.n52 585
R296 B.n308 B.n307 585
R297 B.n306 B.n53 585
R298 B.n305 B.n304 585
R299 B.n303 B.n54 585
R300 B.n302 B.n301 585
R301 B.n300 B.n55 585
R302 B.n299 B.n298 585
R303 B.n297 B.n56 585
R304 B.n296 B.n295 585
R305 B.n294 B.n57 585
R306 B.n293 B.n292 585
R307 B.n291 B.n58 585
R308 B.n290 B.n289 585
R309 B.n288 B.n59 585
R310 B.n287 B.n286 585
R311 B.n285 B.n60 585
R312 B.n284 B.n283 585
R313 B.n282 B.n61 585
R314 B.n281 B.n280 585
R315 B.n279 B.n62 585
R316 B.n278 B.n277 585
R317 B.n276 B.n63 585
R318 B.n275 B.n274 585
R319 B.n273 B.n64 585
R320 B.n272 B.n271 585
R321 B.n270 B.n65 585
R322 B.n269 B.n268 585
R323 B.n267 B.n66 585
R324 B.n266 B.n265 585
R325 B.n264 B.n67 585
R326 B.n263 B.n262 585
R327 B.n261 B.n68 585
R328 B.n260 B.n259 585
R329 B.n258 B.n69 585
R330 B.n257 B.n256 585
R331 B.n255 B.n70 585
R332 B.n254 B.n253 585
R333 B.n252 B.n71 585
R334 B.n251 B.n250 585
R335 B.n249 B.n72 585
R336 B.n248 B.n247 585
R337 B.n246 B.n73 585
R338 B.n245 B.n244 585
R339 B.n243 B.n74 585
R340 B.n242 B.n241 585
R341 B.n240 B.n75 585
R342 B.n239 B.n238 585
R343 B.n237 B.n76 585
R344 B.n236 B.n235 585
R345 B.n234 B.n77 585
R346 B.n233 B.n232 585
R347 B.n231 B.n78 585
R348 B.n230 B.n229 585
R349 B.n228 B.n79 585
R350 B.n227 B.n226 585
R351 B.n176 B.n175 585
R352 B.n177 B.n100 585
R353 B.n179 B.n178 585
R354 B.n180 B.n99 585
R355 B.n182 B.n181 585
R356 B.n183 B.n98 585
R357 B.n185 B.n184 585
R358 B.n186 B.n97 585
R359 B.n188 B.n187 585
R360 B.n189 B.n96 585
R361 B.n191 B.n190 585
R362 B.n192 B.n93 585
R363 B.n195 B.n194 585
R364 B.n196 B.n92 585
R365 B.n198 B.n197 585
R366 B.n199 B.n91 585
R367 B.n201 B.n200 585
R368 B.n202 B.n90 585
R369 B.n204 B.n203 585
R370 B.n205 B.n89 585
R371 B.n207 B.n206 585
R372 B.n209 B.n208 585
R373 B.n210 B.n85 585
R374 B.n212 B.n211 585
R375 B.n213 B.n84 585
R376 B.n215 B.n214 585
R377 B.n216 B.n83 585
R378 B.n218 B.n217 585
R379 B.n219 B.n82 585
R380 B.n221 B.n220 585
R381 B.n222 B.n81 585
R382 B.n224 B.n223 585
R383 B.n225 B.n80 585
R384 B.n174 B.n101 585
R385 B.n173 B.n172 585
R386 B.n171 B.n102 585
R387 B.n170 B.n169 585
R388 B.n168 B.n103 585
R389 B.n167 B.n166 585
R390 B.n165 B.n104 585
R391 B.n164 B.n163 585
R392 B.n162 B.n105 585
R393 B.n161 B.n160 585
R394 B.n159 B.n106 585
R395 B.n158 B.n157 585
R396 B.n156 B.n107 585
R397 B.n155 B.n154 585
R398 B.n153 B.n108 585
R399 B.n152 B.n151 585
R400 B.n150 B.n109 585
R401 B.n149 B.n148 585
R402 B.n147 B.n110 585
R403 B.n146 B.n145 585
R404 B.n144 B.n111 585
R405 B.n143 B.n142 585
R406 B.n141 B.n112 585
R407 B.n140 B.n139 585
R408 B.n138 B.n113 585
R409 B.n137 B.n136 585
R410 B.n135 B.n114 585
R411 B.n134 B.n133 585
R412 B.n132 B.n115 585
R413 B.n131 B.n130 585
R414 B.n129 B.n116 585
R415 B.n128 B.n127 585
R416 B.n126 B.n117 585
R417 B.n125 B.n124 585
R418 B.n123 B.n118 585
R419 B.n122 B.n121 585
R420 B.n120 B.n119 585
R421 B.n2 B.n0 585
R422 B.n449 B.n1 585
R423 B.n448 B.n447 585
R424 B.n446 B.n3 585
R425 B.n445 B.n444 585
R426 B.n443 B.n4 585
R427 B.n442 B.n441 585
R428 B.n440 B.n5 585
R429 B.n439 B.n438 585
R430 B.n437 B.n6 585
R431 B.n436 B.n435 585
R432 B.n434 B.n7 585
R433 B.n433 B.n432 585
R434 B.n431 B.n8 585
R435 B.n430 B.n429 585
R436 B.n428 B.n9 585
R437 B.n427 B.n426 585
R438 B.n425 B.n10 585
R439 B.n424 B.n423 585
R440 B.n422 B.n11 585
R441 B.n421 B.n420 585
R442 B.n419 B.n12 585
R443 B.n418 B.n417 585
R444 B.n416 B.n13 585
R445 B.n415 B.n414 585
R446 B.n413 B.n14 585
R447 B.n412 B.n411 585
R448 B.n410 B.n15 585
R449 B.n409 B.n408 585
R450 B.n407 B.n16 585
R451 B.n406 B.n405 585
R452 B.n404 B.n17 585
R453 B.n403 B.n402 585
R454 B.n401 B.n18 585
R455 B.n400 B.n399 585
R456 B.n398 B.n19 585
R457 B.n397 B.n396 585
R458 B.n395 B.n20 585
R459 B.n394 B.n393 585
R460 B.n451 B.n450 585
R461 B.n176 B.n101 444.452
R462 B.n394 B.n21 444.452
R463 B.n226 B.n225 444.452
R464 B.n340 B.n41 444.452
R465 B.n86 B.t8 292.75
R466 B.n34 B.t4 292.75
R467 B.n94 B.t2 292.75
R468 B.n28 B.t10 292.75
R469 B.n87 B.t7 243.684
R470 B.n35 B.t5 243.684
R471 B.n95 B.t1 243.683
R472 B.n29 B.t11 243.683
R473 B.n86 B.t6 226.631
R474 B.n94 B.t0 226.631
R475 B.n28 B.t9 226.631
R476 B.n34 B.t3 226.631
R477 B.n172 B.n101 163.367
R478 B.n172 B.n171 163.367
R479 B.n171 B.n170 163.367
R480 B.n170 B.n103 163.367
R481 B.n166 B.n103 163.367
R482 B.n166 B.n165 163.367
R483 B.n165 B.n164 163.367
R484 B.n164 B.n105 163.367
R485 B.n160 B.n105 163.367
R486 B.n160 B.n159 163.367
R487 B.n159 B.n158 163.367
R488 B.n158 B.n107 163.367
R489 B.n154 B.n107 163.367
R490 B.n154 B.n153 163.367
R491 B.n153 B.n152 163.367
R492 B.n152 B.n109 163.367
R493 B.n148 B.n109 163.367
R494 B.n148 B.n147 163.367
R495 B.n147 B.n146 163.367
R496 B.n146 B.n111 163.367
R497 B.n142 B.n111 163.367
R498 B.n142 B.n141 163.367
R499 B.n141 B.n140 163.367
R500 B.n140 B.n113 163.367
R501 B.n136 B.n113 163.367
R502 B.n136 B.n135 163.367
R503 B.n135 B.n134 163.367
R504 B.n134 B.n115 163.367
R505 B.n130 B.n115 163.367
R506 B.n130 B.n129 163.367
R507 B.n129 B.n128 163.367
R508 B.n128 B.n117 163.367
R509 B.n124 B.n117 163.367
R510 B.n124 B.n123 163.367
R511 B.n123 B.n122 163.367
R512 B.n122 B.n119 163.367
R513 B.n119 B.n2 163.367
R514 B.n450 B.n2 163.367
R515 B.n450 B.n449 163.367
R516 B.n449 B.n448 163.367
R517 B.n448 B.n3 163.367
R518 B.n444 B.n3 163.367
R519 B.n444 B.n443 163.367
R520 B.n443 B.n442 163.367
R521 B.n442 B.n5 163.367
R522 B.n438 B.n5 163.367
R523 B.n438 B.n437 163.367
R524 B.n437 B.n436 163.367
R525 B.n436 B.n7 163.367
R526 B.n432 B.n7 163.367
R527 B.n432 B.n431 163.367
R528 B.n431 B.n430 163.367
R529 B.n430 B.n9 163.367
R530 B.n426 B.n9 163.367
R531 B.n426 B.n425 163.367
R532 B.n425 B.n424 163.367
R533 B.n424 B.n11 163.367
R534 B.n420 B.n11 163.367
R535 B.n420 B.n419 163.367
R536 B.n419 B.n418 163.367
R537 B.n418 B.n13 163.367
R538 B.n414 B.n13 163.367
R539 B.n414 B.n413 163.367
R540 B.n413 B.n412 163.367
R541 B.n412 B.n15 163.367
R542 B.n408 B.n15 163.367
R543 B.n408 B.n407 163.367
R544 B.n407 B.n406 163.367
R545 B.n406 B.n17 163.367
R546 B.n402 B.n17 163.367
R547 B.n402 B.n401 163.367
R548 B.n401 B.n400 163.367
R549 B.n400 B.n19 163.367
R550 B.n396 B.n19 163.367
R551 B.n396 B.n395 163.367
R552 B.n395 B.n394 163.367
R553 B.n177 B.n176 163.367
R554 B.n178 B.n177 163.367
R555 B.n178 B.n99 163.367
R556 B.n182 B.n99 163.367
R557 B.n183 B.n182 163.367
R558 B.n184 B.n183 163.367
R559 B.n184 B.n97 163.367
R560 B.n188 B.n97 163.367
R561 B.n189 B.n188 163.367
R562 B.n190 B.n189 163.367
R563 B.n190 B.n93 163.367
R564 B.n195 B.n93 163.367
R565 B.n196 B.n195 163.367
R566 B.n197 B.n196 163.367
R567 B.n197 B.n91 163.367
R568 B.n201 B.n91 163.367
R569 B.n202 B.n201 163.367
R570 B.n203 B.n202 163.367
R571 B.n203 B.n89 163.367
R572 B.n207 B.n89 163.367
R573 B.n208 B.n207 163.367
R574 B.n208 B.n85 163.367
R575 B.n212 B.n85 163.367
R576 B.n213 B.n212 163.367
R577 B.n214 B.n213 163.367
R578 B.n214 B.n83 163.367
R579 B.n218 B.n83 163.367
R580 B.n219 B.n218 163.367
R581 B.n220 B.n219 163.367
R582 B.n220 B.n81 163.367
R583 B.n224 B.n81 163.367
R584 B.n225 B.n224 163.367
R585 B.n226 B.n79 163.367
R586 B.n230 B.n79 163.367
R587 B.n231 B.n230 163.367
R588 B.n232 B.n231 163.367
R589 B.n232 B.n77 163.367
R590 B.n236 B.n77 163.367
R591 B.n237 B.n236 163.367
R592 B.n238 B.n237 163.367
R593 B.n238 B.n75 163.367
R594 B.n242 B.n75 163.367
R595 B.n243 B.n242 163.367
R596 B.n244 B.n243 163.367
R597 B.n244 B.n73 163.367
R598 B.n248 B.n73 163.367
R599 B.n249 B.n248 163.367
R600 B.n250 B.n249 163.367
R601 B.n250 B.n71 163.367
R602 B.n254 B.n71 163.367
R603 B.n255 B.n254 163.367
R604 B.n256 B.n255 163.367
R605 B.n256 B.n69 163.367
R606 B.n260 B.n69 163.367
R607 B.n261 B.n260 163.367
R608 B.n262 B.n261 163.367
R609 B.n262 B.n67 163.367
R610 B.n266 B.n67 163.367
R611 B.n267 B.n266 163.367
R612 B.n268 B.n267 163.367
R613 B.n268 B.n65 163.367
R614 B.n272 B.n65 163.367
R615 B.n273 B.n272 163.367
R616 B.n274 B.n273 163.367
R617 B.n274 B.n63 163.367
R618 B.n278 B.n63 163.367
R619 B.n279 B.n278 163.367
R620 B.n280 B.n279 163.367
R621 B.n280 B.n61 163.367
R622 B.n284 B.n61 163.367
R623 B.n285 B.n284 163.367
R624 B.n286 B.n285 163.367
R625 B.n286 B.n59 163.367
R626 B.n290 B.n59 163.367
R627 B.n291 B.n290 163.367
R628 B.n292 B.n291 163.367
R629 B.n292 B.n57 163.367
R630 B.n296 B.n57 163.367
R631 B.n297 B.n296 163.367
R632 B.n298 B.n297 163.367
R633 B.n298 B.n55 163.367
R634 B.n302 B.n55 163.367
R635 B.n303 B.n302 163.367
R636 B.n304 B.n303 163.367
R637 B.n304 B.n53 163.367
R638 B.n308 B.n53 163.367
R639 B.n309 B.n308 163.367
R640 B.n310 B.n309 163.367
R641 B.n310 B.n51 163.367
R642 B.n314 B.n51 163.367
R643 B.n315 B.n314 163.367
R644 B.n316 B.n315 163.367
R645 B.n316 B.n49 163.367
R646 B.n320 B.n49 163.367
R647 B.n321 B.n320 163.367
R648 B.n322 B.n321 163.367
R649 B.n322 B.n47 163.367
R650 B.n326 B.n47 163.367
R651 B.n327 B.n326 163.367
R652 B.n328 B.n327 163.367
R653 B.n328 B.n45 163.367
R654 B.n332 B.n45 163.367
R655 B.n333 B.n332 163.367
R656 B.n334 B.n333 163.367
R657 B.n334 B.n43 163.367
R658 B.n338 B.n43 163.367
R659 B.n339 B.n338 163.367
R660 B.n340 B.n339 163.367
R661 B.n390 B.n21 163.367
R662 B.n390 B.n389 163.367
R663 B.n389 B.n388 163.367
R664 B.n388 B.n23 163.367
R665 B.n384 B.n23 163.367
R666 B.n384 B.n383 163.367
R667 B.n383 B.n382 163.367
R668 B.n382 B.n25 163.367
R669 B.n378 B.n25 163.367
R670 B.n378 B.n377 163.367
R671 B.n377 B.n376 163.367
R672 B.n376 B.n27 163.367
R673 B.n371 B.n27 163.367
R674 B.n371 B.n370 163.367
R675 B.n370 B.n369 163.367
R676 B.n369 B.n31 163.367
R677 B.n365 B.n31 163.367
R678 B.n365 B.n364 163.367
R679 B.n364 B.n363 163.367
R680 B.n363 B.n33 163.367
R681 B.n358 B.n33 163.367
R682 B.n358 B.n357 163.367
R683 B.n357 B.n356 163.367
R684 B.n356 B.n37 163.367
R685 B.n352 B.n37 163.367
R686 B.n352 B.n351 163.367
R687 B.n351 B.n350 163.367
R688 B.n350 B.n39 163.367
R689 B.n346 B.n39 163.367
R690 B.n346 B.n345 163.367
R691 B.n345 B.n344 163.367
R692 B.n344 B.n41 163.367
R693 B.n88 B.n87 59.5399
R694 B.n193 B.n95 59.5399
R695 B.n374 B.n29 59.5399
R696 B.n360 B.n35 59.5399
R697 B.n87 B.n86 49.0672
R698 B.n95 B.n94 49.0672
R699 B.n29 B.n28 49.0672
R700 B.n35 B.n34 49.0672
R701 B.n342 B.n341 28.8785
R702 B.n393 B.n392 28.8785
R703 B.n227 B.n80 28.8785
R704 B.n175 B.n174 28.8785
R705 B B.n451 18.0485
R706 B.n392 B.n391 10.6151
R707 B.n391 B.n22 10.6151
R708 B.n387 B.n22 10.6151
R709 B.n387 B.n386 10.6151
R710 B.n386 B.n385 10.6151
R711 B.n385 B.n24 10.6151
R712 B.n381 B.n24 10.6151
R713 B.n381 B.n380 10.6151
R714 B.n380 B.n379 10.6151
R715 B.n379 B.n26 10.6151
R716 B.n375 B.n26 10.6151
R717 B.n373 B.n372 10.6151
R718 B.n372 B.n30 10.6151
R719 B.n368 B.n30 10.6151
R720 B.n368 B.n367 10.6151
R721 B.n367 B.n366 10.6151
R722 B.n366 B.n32 10.6151
R723 B.n362 B.n32 10.6151
R724 B.n362 B.n361 10.6151
R725 B.n359 B.n36 10.6151
R726 B.n355 B.n36 10.6151
R727 B.n355 B.n354 10.6151
R728 B.n354 B.n353 10.6151
R729 B.n353 B.n38 10.6151
R730 B.n349 B.n38 10.6151
R731 B.n349 B.n348 10.6151
R732 B.n348 B.n347 10.6151
R733 B.n347 B.n40 10.6151
R734 B.n343 B.n40 10.6151
R735 B.n343 B.n342 10.6151
R736 B.n228 B.n227 10.6151
R737 B.n229 B.n228 10.6151
R738 B.n229 B.n78 10.6151
R739 B.n233 B.n78 10.6151
R740 B.n234 B.n233 10.6151
R741 B.n235 B.n234 10.6151
R742 B.n235 B.n76 10.6151
R743 B.n239 B.n76 10.6151
R744 B.n240 B.n239 10.6151
R745 B.n241 B.n240 10.6151
R746 B.n241 B.n74 10.6151
R747 B.n245 B.n74 10.6151
R748 B.n246 B.n245 10.6151
R749 B.n247 B.n246 10.6151
R750 B.n247 B.n72 10.6151
R751 B.n251 B.n72 10.6151
R752 B.n252 B.n251 10.6151
R753 B.n253 B.n252 10.6151
R754 B.n253 B.n70 10.6151
R755 B.n257 B.n70 10.6151
R756 B.n258 B.n257 10.6151
R757 B.n259 B.n258 10.6151
R758 B.n259 B.n68 10.6151
R759 B.n263 B.n68 10.6151
R760 B.n264 B.n263 10.6151
R761 B.n265 B.n264 10.6151
R762 B.n265 B.n66 10.6151
R763 B.n269 B.n66 10.6151
R764 B.n270 B.n269 10.6151
R765 B.n271 B.n270 10.6151
R766 B.n271 B.n64 10.6151
R767 B.n275 B.n64 10.6151
R768 B.n276 B.n275 10.6151
R769 B.n277 B.n276 10.6151
R770 B.n277 B.n62 10.6151
R771 B.n281 B.n62 10.6151
R772 B.n282 B.n281 10.6151
R773 B.n283 B.n282 10.6151
R774 B.n283 B.n60 10.6151
R775 B.n287 B.n60 10.6151
R776 B.n288 B.n287 10.6151
R777 B.n289 B.n288 10.6151
R778 B.n289 B.n58 10.6151
R779 B.n293 B.n58 10.6151
R780 B.n294 B.n293 10.6151
R781 B.n295 B.n294 10.6151
R782 B.n295 B.n56 10.6151
R783 B.n299 B.n56 10.6151
R784 B.n300 B.n299 10.6151
R785 B.n301 B.n300 10.6151
R786 B.n301 B.n54 10.6151
R787 B.n305 B.n54 10.6151
R788 B.n306 B.n305 10.6151
R789 B.n307 B.n306 10.6151
R790 B.n307 B.n52 10.6151
R791 B.n311 B.n52 10.6151
R792 B.n312 B.n311 10.6151
R793 B.n313 B.n312 10.6151
R794 B.n313 B.n50 10.6151
R795 B.n317 B.n50 10.6151
R796 B.n318 B.n317 10.6151
R797 B.n319 B.n318 10.6151
R798 B.n319 B.n48 10.6151
R799 B.n323 B.n48 10.6151
R800 B.n324 B.n323 10.6151
R801 B.n325 B.n324 10.6151
R802 B.n325 B.n46 10.6151
R803 B.n329 B.n46 10.6151
R804 B.n330 B.n329 10.6151
R805 B.n331 B.n330 10.6151
R806 B.n331 B.n44 10.6151
R807 B.n335 B.n44 10.6151
R808 B.n336 B.n335 10.6151
R809 B.n337 B.n336 10.6151
R810 B.n337 B.n42 10.6151
R811 B.n341 B.n42 10.6151
R812 B.n175 B.n100 10.6151
R813 B.n179 B.n100 10.6151
R814 B.n180 B.n179 10.6151
R815 B.n181 B.n180 10.6151
R816 B.n181 B.n98 10.6151
R817 B.n185 B.n98 10.6151
R818 B.n186 B.n185 10.6151
R819 B.n187 B.n186 10.6151
R820 B.n187 B.n96 10.6151
R821 B.n191 B.n96 10.6151
R822 B.n192 B.n191 10.6151
R823 B.n194 B.n92 10.6151
R824 B.n198 B.n92 10.6151
R825 B.n199 B.n198 10.6151
R826 B.n200 B.n199 10.6151
R827 B.n200 B.n90 10.6151
R828 B.n204 B.n90 10.6151
R829 B.n205 B.n204 10.6151
R830 B.n206 B.n205 10.6151
R831 B.n210 B.n209 10.6151
R832 B.n211 B.n210 10.6151
R833 B.n211 B.n84 10.6151
R834 B.n215 B.n84 10.6151
R835 B.n216 B.n215 10.6151
R836 B.n217 B.n216 10.6151
R837 B.n217 B.n82 10.6151
R838 B.n221 B.n82 10.6151
R839 B.n222 B.n221 10.6151
R840 B.n223 B.n222 10.6151
R841 B.n223 B.n80 10.6151
R842 B.n174 B.n173 10.6151
R843 B.n173 B.n102 10.6151
R844 B.n169 B.n102 10.6151
R845 B.n169 B.n168 10.6151
R846 B.n168 B.n167 10.6151
R847 B.n167 B.n104 10.6151
R848 B.n163 B.n104 10.6151
R849 B.n163 B.n162 10.6151
R850 B.n162 B.n161 10.6151
R851 B.n161 B.n106 10.6151
R852 B.n157 B.n106 10.6151
R853 B.n157 B.n156 10.6151
R854 B.n156 B.n155 10.6151
R855 B.n155 B.n108 10.6151
R856 B.n151 B.n108 10.6151
R857 B.n151 B.n150 10.6151
R858 B.n150 B.n149 10.6151
R859 B.n149 B.n110 10.6151
R860 B.n145 B.n110 10.6151
R861 B.n145 B.n144 10.6151
R862 B.n144 B.n143 10.6151
R863 B.n143 B.n112 10.6151
R864 B.n139 B.n112 10.6151
R865 B.n139 B.n138 10.6151
R866 B.n138 B.n137 10.6151
R867 B.n137 B.n114 10.6151
R868 B.n133 B.n114 10.6151
R869 B.n133 B.n132 10.6151
R870 B.n132 B.n131 10.6151
R871 B.n131 B.n116 10.6151
R872 B.n127 B.n116 10.6151
R873 B.n127 B.n126 10.6151
R874 B.n126 B.n125 10.6151
R875 B.n125 B.n118 10.6151
R876 B.n121 B.n118 10.6151
R877 B.n121 B.n120 10.6151
R878 B.n120 B.n0 10.6151
R879 B.n447 B.n1 10.6151
R880 B.n447 B.n446 10.6151
R881 B.n446 B.n445 10.6151
R882 B.n445 B.n4 10.6151
R883 B.n441 B.n4 10.6151
R884 B.n441 B.n440 10.6151
R885 B.n440 B.n439 10.6151
R886 B.n439 B.n6 10.6151
R887 B.n435 B.n6 10.6151
R888 B.n435 B.n434 10.6151
R889 B.n434 B.n433 10.6151
R890 B.n433 B.n8 10.6151
R891 B.n429 B.n8 10.6151
R892 B.n429 B.n428 10.6151
R893 B.n428 B.n427 10.6151
R894 B.n427 B.n10 10.6151
R895 B.n423 B.n10 10.6151
R896 B.n423 B.n422 10.6151
R897 B.n422 B.n421 10.6151
R898 B.n421 B.n12 10.6151
R899 B.n417 B.n12 10.6151
R900 B.n417 B.n416 10.6151
R901 B.n416 B.n415 10.6151
R902 B.n415 B.n14 10.6151
R903 B.n411 B.n14 10.6151
R904 B.n411 B.n410 10.6151
R905 B.n410 B.n409 10.6151
R906 B.n409 B.n16 10.6151
R907 B.n405 B.n16 10.6151
R908 B.n405 B.n404 10.6151
R909 B.n404 B.n403 10.6151
R910 B.n403 B.n18 10.6151
R911 B.n399 B.n18 10.6151
R912 B.n399 B.n398 10.6151
R913 B.n398 B.n397 10.6151
R914 B.n397 B.n20 10.6151
R915 B.n393 B.n20 10.6151
R916 B.n374 B.n373 6.5566
R917 B.n361 B.n360 6.5566
R918 B.n194 B.n193 6.5566
R919 B.n206 B.n88 6.5566
R920 B.n375 B.n374 4.05904
R921 B.n360 B.n359 4.05904
R922 B.n193 B.n192 4.05904
R923 B.n209 B.n88 4.05904
R924 B.n451 B.n0 2.81026
R925 B.n451 B.n1 2.81026
C0 B w_n2994_n1320# 6.28628f
C1 VDD1 w_n2994_n1320# 1.46712f
C2 VP w_n2994_n1320# 5.75961f
C3 VTAIL VDD2 3.78631f
C4 VTAIL VN 2.02328f
C5 VN VDD2 1.28273f
C6 VTAIL B 1.202f
C7 B VDD2 1.25011f
C8 VDD1 VTAIL 3.73586f
C9 VDD1 VDD2 1.24846f
C10 VTAIL VP 2.03742f
C11 VP VDD2 0.431448f
C12 B VN 0.946818f
C13 VTAIL w_n2994_n1320# 1.43347f
C14 VDD2 w_n2994_n1320# 1.53866f
C15 VDD1 VN 0.157061f
C16 VP VN 4.64768f
C17 VDD1 B 1.18526f
C18 VP B 1.58837f
C19 VN w_n2994_n1320# 5.37907f
C20 VDD1 VP 1.55455f
C21 VDD2 VSUBS 0.967329f
C22 VDD1 VSUBS 1.211298f
C23 VTAIL VSUBS 0.475804f
C24 VN VSUBS 5.2247f
C25 VP VSUBS 2.064043f
C26 B VSUBS 3.182658f
C27 w_n2994_n1320# VSUBS 50.5507f
C28 B.n0 VSUBS 0.005756f
C29 B.n1 VSUBS 0.005756f
C30 B.n2 VSUBS 0.009102f
C31 B.n3 VSUBS 0.009102f
C32 B.n4 VSUBS 0.009102f
C33 B.n5 VSUBS 0.009102f
C34 B.n6 VSUBS 0.009102f
C35 B.n7 VSUBS 0.009102f
C36 B.n8 VSUBS 0.009102f
C37 B.n9 VSUBS 0.009102f
C38 B.n10 VSUBS 0.009102f
C39 B.n11 VSUBS 0.009102f
C40 B.n12 VSUBS 0.009102f
C41 B.n13 VSUBS 0.009102f
C42 B.n14 VSUBS 0.009102f
C43 B.n15 VSUBS 0.009102f
C44 B.n16 VSUBS 0.009102f
C45 B.n17 VSUBS 0.009102f
C46 B.n18 VSUBS 0.009102f
C47 B.n19 VSUBS 0.009102f
C48 B.n20 VSUBS 0.009102f
C49 B.n21 VSUBS 0.020345f
C50 B.n22 VSUBS 0.009102f
C51 B.n23 VSUBS 0.009102f
C52 B.n24 VSUBS 0.009102f
C53 B.n25 VSUBS 0.009102f
C54 B.n26 VSUBS 0.009102f
C55 B.n27 VSUBS 0.009102f
C56 B.t11 VSUBS 0.038745f
C57 B.t10 VSUBS 0.049903f
C58 B.t9 VSUBS 0.248579f
C59 B.n28 VSUBS 0.094035f
C60 B.n29 VSUBS 0.079554f
C61 B.n30 VSUBS 0.009102f
C62 B.n31 VSUBS 0.009102f
C63 B.n32 VSUBS 0.009102f
C64 B.n33 VSUBS 0.009102f
C65 B.t5 VSUBS 0.038745f
C66 B.t4 VSUBS 0.049903f
C67 B.t3 VSUBS 0.248579f
C68 B.n34 VSUBS 0.094034f
C69 B.n35 VSUBS 0.079554f
C70 B.n36 VSUBS 0.009102f
C71 B.n37 VSUBS 0.009102f
C72 B.n38 VSUBS 0.009102f
C73 B.n39 VSUBS 0.009102f
C74 B.n40 VSUBS 0.009102f
C75 B.n41 VSUBS 0.020345f
C76 B.n42 VSUBS 0.009102f
C77 B.n43 VSUBS 0.009102f
C78 B.n44 VSUBS 0.009102f
C79 B.n45 VSUBS 0.009102f
C80 B.n46 VSUBS 0.009102f
C81 B.n47 VSUBS 0.009102f
C82 B.n48 VSUBS 0.009102f
C83 B.n49 VSUBS 0.009102f
C84 B.n50 VSUBS 0.009102f
C85 B.n51 VSUBS 0.009102f
C86 B.n52 VSUBS 0.009102f
C87 B.n53 VSUBS 0.009102f
C88 B.n54 VSUBS 0.009102f
C89 B.n55 VSUBS 0.009102f
C90 B.n56 VSUBS 0.009102f
C91 B.n57 VSUBS 0.009102f
C92 B.n58 VSUBS 0.009102f
C93 B.n59 VSUBS 0.009102f
C94 B.n60 VSUBS 0.009102f
C95 B.n61 VSUBS 0.009102f
C96 B.n62 VSUBS 0.009102f
C97 B.n63 VSUBS 0.009102f
C98 B.n64 VSUBS 0.009102f
C99 B.n65 VSUBS 0.009102f
C100 B.n66 VSUBS 0.009102f
C101 B.n67 VSUBS 0.009102f
C102 B.n68 VSUBS 0.009102f
C103 B.n69 VSUBS 0.009102f
C104 B.n70 VSUBS 0.009102f
C105 B.n71 VSUBS 0.009102f
C106 B.n72 VSUBS 0.009102f
C107 B.n73 VSUBS 0.009102f
C108 B.n74 VSUBS 0.009102f
C109 B.n75 VSUBS 0.009102f
C110 B.n76 VSUBS 0.009102f
C111 B.n77 VSUBS 0.009102f
C112 B.n78 VSUBS 0.009102f
C113 B.n79 VSUBS 0.009102f
C114 B.n80 VSUBS 0.020345f
C115 B.n81 VSUBS 0.009102f
C116 B.n82 VSUBS 0.009102f
C117 B.n83 VSUBS 0.009102f
C118 B.n84 VSUBS 0.009102f
C119 B.n85 VSUBS 0.009102f
C120 B.t7 VSUBS 0.038745f
C121 B.t8 VSUBS 0.049903f
C122 B.t6 VSUBS 0.248579f
C123 B.n86 VSUBS 0.094034f
C124 B.n87 VSUBS 0.079554f
C125 B.n88 VSUBS 0.021089f
C126 B.n89 VSUBS 0.009102f
C127 B.n90 VSUBS 0.009102f
C128 B.n91 VSUBS 0.009102f
C129 B.n92 VSUBS 0.009102f
C130 B.n93 VSUBS 0.009102f
C131 B.t1 VSUBS 0.038745f
C132 B.t2 VSUBS 0.049903f
C133 B.t0 VSUBS 0.248579f
C134 B.n94 VSUBS 0.094035f
C135 B.n95 VSUBS 0.079554f
C136 B.n96 VSUBS 0.009102f
C137 B.n97 VSUBS 0.009102f
C138 B.n98 VSUBS 0.009102f
C139 B.n99 VSUBS 0.009102f
C140 B.n100 VSUBS 0.009102f
C141 B.n101 VSUBS 0.01901f
C142 B.n102 VSUBS 0.009102f
C143 B.n103 VSUBS 0.009102f
C144 B.n104 VSUBS 0.009102f
C145 B.n105 VSUBS 0.009102f
C146 B.n106 VSUBS 0.009102f
C147 B.n107 VSUBS 0.009102f
C148 B.n108 VSUBS 0.009102f
C149 B.n109 VSUBS 0.009102f
C150 B.n110 VSUBS 0.009102f
C151 B.n111 VSUBS 0.009102f
C152 B.n112 VSUBS 0.009102f
C153 B.n113 VSUBS 0.009102f
C154 B.n114 VSUBS 0.009102f
C155 B.n115 VSUBS 0.009102f
C156 B.n116 VSUBS 0.009102f
C157 B.n117 VSUBS 0.009102f
C158 B.n118 VSUBS 0.009102f
C159 B.n119 VSUBS 0.009102f
C160 B.n120 VSUBS 0.009102f
C161 B.n121 VSUBS 0.009102f
C162 B.n122 VSUBS 0.009102f
C163 B.n123 VSUBS 0.009102f
C164 B.n124 VSUBS 0.009102f
C165 B.n125 VSUBS 0.009102f
C166 B.n126 VSUBS 0.009102f
C167 B.n127 VSUBS 0.009102f
C168 B.n128 VSUBS 0.009102f
C169 B.n129 VSUBS 0.009102f
C170 B.n130 VSUBS 0.009102f
C171 B.n131 VSUBS 0.009102f
C172 B.n132 VSUBS 0.009102f
C173 B.n133 VSUBS 0.009102f
C174 B.n134 VSUBS 0.009102f
C175 B.n135 VSUBS 0.009102f
C176 B.n136 VSUBS 0.009102f
C177 B.n137 VSUBS 0.009102f
C178 B.n138 VSUBS 0.009102f
C179 B.n139 VSUBS 0.009102f
C180 B.n140 VSUBS 0.009102f
C181 B.n141 VSUBS 0.009102f
C182 B.n142 VSUBS 0.009102f
C183 B.n143 VSUBS 0.009102f
C184 B.n144 VSUBS 0.009102f
C185 B.n145 VSUBS 0.009102f
C186 B.n146 VSUBS 0.009102f
C187 B.n147 VSUBS 0.009102f
C188 B.n148 VSUBS 0.009102f
C189 B.n149 VSUBS 0.009102f
C190 B.n150 VSUBS 0.009102f
C191 B.n151 VSUBS 0.009102f
C192 B.n152 VSUBS 0.009102f
C193 B.n153 VSUBS 0.009102f
C194 B.n154 VSUBS 0.009102f
C195 B.n155 VSUBS 0.009102f
C196 B.n156 VSUBS 0.009102f
C197 B.n157 VSUBS 0.009102f
C198 B.n158 VSUBS 0.009102f
C199 B.n159 VSUBS 0.009102f
C200 B.n160 VSUBS 0.009102f
C201 B.n161 VSUBS 0.009102f
C202 B.n162 VSUBS 0.009102f
C203 B.n163 VSUBS 0.009102f
C204 B.n164 VSUBS 0.009102f
C205 B.n165 VSUBS 0.009102f
C206 B.n166 VSUBS 0.009102f
C207 B.n167 VSUBS 0.009102f
C208 B.n168 VSUBS 0.009102f
C209 B.n169 VSUBS 0.009102f
C210 B.n170 VSUBS 0.009102f
C211 B.n171 VSUBS 0.009102f
C212 B.n172 VSUBS 0.009102f
C213 B.n173 VSUBS 0.009102f
C214 B.n174 VSUBS 0.01901f
C215 B.n175 VSUBS 0.020345f
C216 B.n176 VSUBS 0.020345f
C217 B.n177 VSUBS 0.009102f
C218 B.n178 VSUBS 0.009102f
C219 B.n179 VSUBS 0.009102f
C220 B.n180 VSUBS 0.009102f
C221 B.n181 VSUBS 0.009102f
C222 B.n182 VSUBS 0.009102f
C223 B.n183 VSUBS 0.009102f
C224 B.n184 VSUBS 0.009102f
C225 B.n185 VSUBS 0.009102f
C226 B.n186 VSUBS 0.009102f
C227 B.n187 VSUBS 0.009102f
C228 B.n188 VSUBS 0.009102f
C229 B.n189 VSUBS 0.009102f
C230 B.n190 VSUBS 0.009102f
C231 B.n191 VSUBS 0.009102f
C232 B.n192 VSUBS 0.006291f
C233 B.n193 VSUBS 0.021089f
C234 B.n194 VSUBS 0.007362f
C235 B.n195 VSUBS 0.009102f
C236 B.n196 VSUBS 0.009102f
C237 B.n197 VSUBS 0.009102f
C238 B.n198 VSUBS 0.009102f
C239 B.n199 VSUBS 0.009102f
C240 B.n200 VSUBS 0.009102f
C241 B.n201 VSUBS 0.009102f
C242 B.n202 VSUBS 0.009102f
C243 B.n203 VSUBS 0.009102f
C244 B.n204 VSUBS 0.009102f
C245 B.n205 VSUBS 0.009102f
C246 B.n206 VSUBS 0.007362f
C247 B.n207 VSUBS 0.009102f
C248 B.n208 VSUBS 0.009102f
C249 B.n209 VSUBS 0.006291f
C250 B.n210 VSUBS 0.009102f
C251 B.n211 VSUBS 0.009102f
C252 B.n212 VSUBS 0.009102f
C253 B.n213 VSUBS 0.009102f
C254 B.n214 VSUBS 0.009102f
C255 B.n215 VSUBS 0.009102f
C256 B.n216 VSUBS 0.009102f
C257 B.n217 VSUBS 0.009102f
C258 B.n218 VSUBS 0.009102f
C259 B.n219 VSUBS 0.009102f
C260 B.n220 VSUBS 0.009102f
C261 B.n221 VSUBS 0.009102f
C262 B.n222 VSUBS 0.009102f
C263 B.n223 VSUBS 0.009102f
C264 B.n224 VSUBS 0.009102f
C265 B.n225 VSUBS 0.020345f
C266 B.n226 VSUBS 0.01901f
C267 B.n227 VSUBS 0.01901f
C268 B.n228 VSUBS 0.009102f
C269 B.n229 VSUBS 0.009102f
C270 B.n230 VSUBS 0.009102f
C271 B.n231 VSUBS 0.009102f
C272 B.n232 VSUBS 0.009102f
C273 B.n233 VSUBS 0.009102f
C274 B.n234 VSUBS 0.009102f
C275 B.n235 VSUBS 0.009102f
C276 B.n236 VSUBS 0.009102f
C277 B.n237 VSUBS 0.009102f
C278 B.n238 VSUBS 0.009102f
C279 B.n239 VSUBS 0.009102f
C280 B.n240 VSUBS 0.009102f
C281 B.n241 VSUBS 0.009102f
C282 B.n242 VSUBS 0.009102f
C283 B.n243 VSUBS 0.009102f
C284 B.n244 VSUBS 0.009102f
C285 B.n245 VSUBS 0.009102f
C286 B.n246 VSUBS 0.009102f
C287 B.n247 VSUBS 0.009102f
C288 B.n248 VSUBS 0.009102f
C289 B.n249 VSUBS 0.009102f
C290 B.n250 VSUBS 0.009102f
C291 B.n251 VSUBS 0.009102f
C292 B.n252 VSUBS 0.009102f
C293 B.n253 VSUBS 0.009102f
C294 B.n254 VSUBS 0.009102f
C295 B.n255 VSUBS 0.009102f
C296 B.n256 VSUBS 0.009102f
C297 B.n257 VSUBS 0.009102f
C298 B.n258 VSUBS 0.009102f
C299 B.n259 VSUBS 0.009102f
C300 B.n260 VSUBS 0.009102f
C301 B.n261 VSUBS 0.009102f
C302 B.n262 VSUBS 0.009102f
C303 B.n263 VSUBS 0.009102f
C304 B.n264 VSUBS 0.009102f
C305 B.n265 VSUBS 0.009102f
C306 B.n266 VSUBS 0.009102f
C307 B.n267 VSUBS 0.009102f
C308 B.n268 VSUBS 0.009102f
C309 B.n269 VSUBS 0.009102f
C310 B.n270 VSUBS 0.009102f
C311 B.n271 VSUBS 0.009102f
C312 B.n272 VSUBS 0.009102f
C313 B.n273 VSUBS 0.009102f
C314 B.n274 VSUBS 0.009102f
C315 B.n275 VSUBS 0.009102f
C316 B.n276 VSUBS 0.009102f
C317 B.n277 VSUBS 0.009102f
C318 B.n278 VSUBS 0.009102f
C319 B.n279 VSUBS 0.009102f
C320 B.n280 VSUBS 0.009102f
C321 B.n281 VSUBS 0.009102f
C322 B.n282 VSUBS 0.009102f
C323 B.n283 VSUBS 0.009102f
C324 B.n284 VSUBS 0.009102f
C325 B.n285 VSUBS 0.009102f
C326 B.n286 VSUBS 0.009102f
C327 B.n287 VSUBS 0.009102f
C328 B.n288 VSUBS 0.009102f
C329 B.n289 VSUBS 0.009102f
C330 B.n290 VSUBS 0.009102f
C331 B.n291 VSUBS 0.009102f
C332 B.n292 VSUBS 0.009102f
C333 B.n293 VSUBS 0.009102f
C334 B.n294 VSUBS 0.009102f
C335 B.n295 VSUBS 0.009102f
C336 B.n296 VSUBS 0.009102f
C337 B.n297 VSUBS 0.009102f
C338 B.n298 VSUBS 0.009102f
C339 B.n299 VSUBS 0.009102f
C340 B.n300 VSUBS 0.009102f
C341 B.n301 VSUBS 0.009102f
C342 B.n302 VSUBS 0.009102f
C343 B.n303 VSUBS 0.009102f
C344 B.n304 VSUBS 0.009102f
C345 B.n305 VSUBS 0.009102f
C346 B.n306 VSUBS 0.009102f
C347 B.n307 VSUBS 0.009102f
C348 B.n308 VSUBS 0.009102f
C349 B.n309 VSUBS 0.009102f
C350 B.n310 VSUBS 0.009102f
C351 B.n311 VSUBS 0.009102f
C352 B.n312 VSUBS 0.009102f
C353 B.n313 VSUBS 0.009102f
C354 B.n314 VSUBS 0.009102f
C355 B.n315 VSUBS 0.009102f
C356 B.n316 VSUBS 0.009102f
C357 B.n317 VSUBS 0.009102f
C358 B.n318 VSUBS 0.009102f
C359 B.n319 VSUBS 0.009102f
C360 B.n320 VSUBS 0.009102f
C361 B.n321 VSUBS 0.009102f
C362 B.n322 VSUBS 0.009102f
C363 B.n323 VSUBS 0.009102f
C364 B.n324 VSUBS 0.009102f
C365 B.n325 VSUBS 0.009102f
C366 B.n326 VSUBS 0.009102f
C367 B.n327 VSUBS 0.009102f
C368 B.n328 VSUBS 0.009102f
C369 B.n329 VSUBS 0.009102f
C370 B.n330 VSUBS 0.009102f
C371 B.n331 VSUBS 0.009102f
C372 B.n332 VSUBS 0.009102f
C373 B.n333 VSUBS 0.009102f
C374 B.n334 VSUBS 0.009102f
C375 B.n335 VSUBS 0.009102f
C376 B.n336 VSUBS 0.009102f
C377 B.n337 VSUBS 0.009102f
C378 B.n338 VSUBS 0.009102f
C379 B.n339 VSUBS 0.009102f
C380 B.n340 VSUBS 0.01901f
C381 B.n341 VSUBS 0.020226f
C382 B.n342 VSUBS 0.019128f
C383 B.n343 VSUBS 0.009102f
C384 B.n344 VSUBS 0.009102f
C385 B.n345 VSUBS 0.009102f
C386 B.n346 VSUBS 0.009102f
C387 B.n347 VSUBS 0.009102f
C388 B.n348 VSUBS 0.009102f
C389 B.n349 VSUBS 0.009102f
C390 B.n350 VSUBS 0.009102f
C391 B.n351 VSUBS 0.009102f
C392 B.n352 VSUBS 0.009102f
C393 B.n353 VSUBS 0.009102f
C394 B.n354 VSUBS 0.009102f
C395 B.n355 VSUBS 0.009102f
C396 B.n356 VSUBS 0.009102f
C397 B.n357 VSUBS 0.009102f
C398 B.n358 VSUBS 0.009102f
C399 B.n359 VSUBS 0.006291f
C400 B.n360 VSUBS 0.021089f
C401 B.n361 VSUBS 0.007362f
C402 B.n362 VSUBS 0.009102f
C403 B.n363 VSUBS 0.009102f
C404 B.n364 VSUBS 0.009102f
C405 B.n365 VSUBS 0.009102f
C406 B.n366 VSUBS 0.009102f
C407 B.n367 VSUBS 0.009102f
C408 B.n368 VSUBS 0.009102f
C409 B.n369 VSUBS 0.009102f
C410 B.n370 VSUBS 0.009102f
C411 B.n371 VSUBS 0.009102f
C412 B.n372 VSUBS 0.009102f
C413 B.n373 VSUBS 0.007362f
C414 B.n374 VSUBS 0.021089f
C415 B.n375 VSUBS 0.006291f
C416 B.n376 VSUBS 0.009102f
C417 B.n377 VSUBS 0.009102f
C418 B.n378 VSUBS 0.009102f
C419 B.n379 VSUBS 0.009102f
C420 B.n380 VSUBS 0.009102f
C421 B.n381 VSUBS 0.009102f
C422 B.n382 VSUBS 0.009102f
C423 B.n383 VSUBS 0.009102f
C424 B.n384 VSUBS 0.009102f
C425 B.n385 VSUBS 0.009102f
C426 B.n386 VSUBS 0.009102f
C427 B.n387 VSUBS 0.009102f
C428 B.n388 VSUBS 0.009102f
C429 B.n389 VSUBS 0.009102f
C430 B.n390 VSUBS 0.009102f
C431 B.n391 VSUBS 0.009102f
C432 B.n392 VSUBS 0.020345f
C433 B.n393 VSUBS 0.01901f
C434 B.n394 VSUBS 0.01901f
C435 B.n395 VSUBS 0.009102f
C436 B.n396 VSUBS 0.009102f
C437 B.n397 VSUBS 0.009102f
C438 B.n398 VSUBS 0.009102f
C439 B.n399 VSUBS 0.009102f
C440 B.n400 VSUBS 0.009102f
C441 B.n401 VSUBS 0.009102f
C442 B.n402 VSUBS 0.009102f
C443 B.n403 VSUBS 0.009102f
C444 B.n404 VSUBS 0.009102f
C445 B.n405 VSUBS 0.009102f
C446 B.n406 VSUBS 0.009102f
C447 B.n407 VSUBS 0.009102f
C448 B.n408 VSUBS 0.009102f
C449 B.n409 VSUBS 0.009102f
C450 B.n410 VSUBS 0.009102f
C451 B.n411 VSUBS 0.009102f
C452 B.n412 VSUBS 0.009102f
C453 B.n413 VSUBS 0.009102f
C454 B.n414 VSUBS 0.009102f
C455 B.n415 VSUBS 0.009102f
C456 B.n416 VSUBS 0.009102f
C457 B.n417 VSUBS 0.009102f
C458 B.n418 VSUBS 0.009102f
C459 B.n419 VSUBS 0.009102f
C460 B.n420 VSUBS 0.009102f
C461 B.n421 VSUBS 0.009102f
C462 B.n422 VSUBS 0.009102f
C463 B.n423 VSUBS 0.009102f
C464 B.n424 VSUBS 0.009102f
C465 B.n425 VSUBS 0.009102f
C466 B.n426 VSUBS 0.009102f
C467 B.n427 VSUBS 0.009102f
C468 B.n428 VSUBS 0.009102f
C469 B.n429 VSUBS 0.009102f
C470 B.n430 VSUBS 0.009102f
C471 B.n431 VSUBS 0.009102f
C472 B.n432 VSUBS 0.009102f
C473 B.n433 VSUBS 0.009102f
C474 B.n434 VSUBS 0.009102f
C475 B.n435 VSUBS 0.009102f
C476 B.n436 VSUBS 0.009102f
C477 B.n437 VSUBS 0.009102f
C478 B.n438 VSUBS 0.009102f
C479 B.n439 VSUBS 0.009102f
C480 B.n440 VSUBS 0.009102f
C481 B.n441 VSUBS 0.009102f
C482 B.n442 VSUBS 0.009102f
C483 B.n443 VSUBS 0.009102f
C484 B.n444 VSUBS 0.009102f
C485 B.n445 VSUBS 0.009102f
C486 B.n446 VSUBS 0.009102f
C487 B.n447 VSUBS 0.009102f
C488 B.n448 VSUBS 0.009102f
C489 B.n449 VSUBS 0.009102f
C490 B.n450 VSUBS 0.009102f
C491 B.n451 VSUBS 0.020611f
C492 VDD1.n0 VSUBS 0.016776f
C493 VDD1.n1 VSUBS 0.044577f
C494 VDD1.t5 VSUBS 0.043083f
C495 VDD1.n2 VSUBS 0.041042f
C496 VDD1.n3 VSUBS 0.011021f
C497 VDD1.n4 VSUBS 0.00878f
C498 VDD1.n5 VSUBS 0.094191f
C499 VDD1.n6 VSUBS 0.038348f
C500 VDD1.n7 VSUBS 0.016776f
C501 VDD1.n8 VSUBS 0.044577f
C502 VDD1.t1 VSUBS 0.043083f
C503 VDD1.n9 VSUBS 0.041042f
C504 VDD1.n10 VSUBS 0.011021f
C505 VDD1.n11 VSUBS 0.00878f
C506 VDD1.n12 VSUBS 0.094191f
C507 VDD1.n13 VSUBS 0.037916f
C508 VDD1.t3 VSUBS 0.022723f
C509 VDD1.t0 VSUBS 0.022723f
C510 VDD1.n14 VSUBS 0.096424f
C511 VDD1.n15 VSUBS 1.33814f
C512 VDD1.t2 VSUBS 0.022723f
C513 VDD1.t4 VSUBS 0.022723f
C514 VDD1.n16 VSUBS 0.095671f
C515 VDD1.n17 VSUBS 1.25114f
C516 VP.n0 VSUBS 0.072502f
C517 VP.t5 VSUBS 0.483742f
C518 VP.n1 VSUBS 0.044576f
C519 VP.n2 VSUBS 0.054995f
C520 VP.t2 VSUBS 0.483742f
C521 VP.n3 VSUBS 0.109464f
C522 VP.n4 VSUBS 0.054995f
C523 VP.t4 VSUBS 0.483742f
C524 VP.n5 VSUBS 0.41366f
C525 VP.n6 VSUBS 0.072502f
C526 VP.t1 VSUBS 0.483742f
C527 VP.n7 VSUBS 0.044576f
C528 VP.n8 VSUBS 0.468074f
C529 VP.t3 VSUBS 0.483742f
C530 VP.t0 VSUBS 0.824021f
C531 VP.n9 VSUBS 0.369134f
C532 VP.n10 VSUBS 0.3903f
C533 VP.n11 VSUBS 0.076811f
C534 VP.n12 VSUBS 0.109464f
C535 VP.n13 VSUBS 0.054995f
C536 VP.n14 VSUBS 0.054995f
C537 VP.n15 VSUBS 0.054995f
C538 VP.n16 VSUBS 0.107833f
C539 VP.n17 VSUBS 0.079831f
C540 VP.n18 VSUBS 0.41366f
C541 VP.n19 VSUBS 2.08612f
C542 VP.n20 VSUBS 2.13653f
C543 VP.n21 VSUBS 0.072502f
C544 VP.n22 VSUBS 0.079831f
C545 VP.n23 VSUBS 0.107833f
C546 VP.n24 VSUBS 0.044576f
C547 VP.n25 VSUBS 0.054995f
C548 VP.n26 VSUBS 0.054995f
C549 VP.n27 VSUBS 0.054995f
C550 VP.n28 VSUBS 0.076811f
C551 VP.n29 VSUBS 0.249269f
C552 VP.n30 VSUBS 0.076811f
C553 VP.n31 VSUBS 0.109464f
C554 VP.n32 VSUBS 0.054995f
C555 VP.n33 VSUBS 0.054995f
C556 VP.n34 VSUBS 0.054995f
C557 VP.n35 VSUBS 0.107833f
C558 VP.n36 VSUBS 0.079831f
C559 VP.n37 VSUBS 0.41366f
C560 VP.n38 VSUBS 0.07801f
C561 VTAIL.t6 VSUBS 0.047881f
C562 VTAIL.t10 VSUBS 0.047881f
C563 VTAIL.n0 VSUBS 0.171288f
C564 VTAIL.n1 VSUBS 0.565145f
C565 VTAIL.n2 VSUBS 0.035349f
C566 VTAIL.n3 VSUBS 0.093928f
C567 VTAIL.t3 VSUBS 0.090781f
C568 VTAIL.n4 VSUBS 0.086481f
C569 VTAIL.n5 VSUBS 0.023223f
C570 VTAIL.n6 VSUBS 0.0185f
C571 VTAIL.n7 VSUBS 0.19847f
C572 VTAIL.n8 VSUBS 0.048726f
C573 VTAIL.n9 VSUBS 0.446563f
C574 VTAIL.t1 VSUBS 0.047881f
C575 VTAIL.t0 VSUBS 0.047881f
C576 VTAIL.n10 VSUBS 0.171288f
C577 VTAIL.n11 VSUBS 1.6869f
C578 VTAIL.t8 VSUBS 0.047881f
C579 VTAIL.t11 VSUBS 0.047881f
C580 VTAIL.n12 VSUBS 0.171289f
C581 VTAIL.n13 VSUBS 1.6869f
C582 VTAIL.n14 VSUBS 0.035349f
C583 VTAIL.n15 VSUBS 0.093928f
C584 VTAIL.t9 VSUBS 0.090781f
C585 VTAIL.n16 VSUBS 0.086481f
C586 VTAIL.n17 VSUBS 0.023223f
C587 VTAIL.n18 VSUBS 0.0185f
C588 VTAIL.n19 VSUBS 0.19847f
C589 VTAIL.n20 VSUBS 0.048726f
C590 VTAIL.n21 VSUBS 0.446563f
C591 VTAIL.t4 VSUBS 0.047881f
C592 VTAIL.t2 VSUBS 0.047881f
C593 VTAIL.n22 VSUBS 0.171289f
C594 VTAIL.n23 VSUBS 0.740148f
C595 VTAIL.n24 VSUBS 0.035349f
C596 VTAIL.n25 VSUBS 0.093928f
C597 VTAIL.t5 VSUBS 0.090781f
C598 VTAIL.n26 VSUBS 0.086481f
C599 VTAIL.n27 VSUBS 0.023223f
C600 VTAIL.n28 VSUBS 0.0185f
C601 VTAIL.n29 VSUBS 0.19847f
C602 VTAIL.n30 VSUBS 0.048726f
C603 VTAIL.n31 VSUBS 1.15137f
C604 VTAIL.n32 VSUBS 0.035349f
C605 VTAIL.n33 VSUBS 0.093928f
C606 VTAIL.t7 VSUBS 0.090781f
C607 VTAIL.n34 VSUBS 0.086481f
C608 VTAIL.n35 VSUBS 0.023223f
C609 VTAIL.n36 VSUBS 0.0185f
C610 VTAIL.n37 VSUBS 0.19847f
C611 VTAIL.n38 VSUBS 0.048726f
C612 VTAIL.n39 VSUBS 1.08443f
C613 VDD2.n0 VSUBS 0.017515f
C614 VDD2.n1 VSUBS 0.046541f
C615 VDD2.t4 VSUBS 0.044981f
C616 VDD2.n2 VSUBS 0.04285f
C617 VDD2.n3 VSUBS 0.011507f
C618 VDD2.n4 VSUBS 0.009166f
C619 VDD2.n5 VSUBS 0.09834f
C620 VDD2.n6 VSUBS 0.039586f
C621 VDD2.t2 VSUBS 0.023725f
C622 VDD2.t5 VSUBS 0.023725f
C623 VDD2.n7 VSUBS 0.100672f
C624 VDD2.n8 VSUBS 1.32637f
C625 VDD2.n9 VSUBS 0.017515f
C626 VDD2.n10 VSUBS 0.046541f
C627 VDD2.t3 VSUBS 0.044981f
C628 VDD2.n11 VSUBS 0.04285f
C629 VDD2.n12 VSUBS 0.011507f
C630 VDD2.n13 VSUBS 0.009166f
C631 VDD2.n14 VSUBS 0.09834f
C632 VDD2.n15 VSUBS 0.035908f
C633 VDD2.n16 VSUBS 1.11821f
C634 VDD2.t0 VSUBS 0.023725f
C635 VDD2.t1 VSUBS 0.023725f
C636 VDD2.n17 VSUBS 0.100665f
C637 VN.n0 VSUBS 0.069728f
C638 VN.t4 VSUBS 0.465237f
C639 VN.n1 VSUBS 0.042871f
C640 VN.n2 VSUBS 0.450168f
C641 VN.t1 VSUBS 0.465237f
C642 VN.t5 VSUBS 0.792499f
C643 VN.n3 VSUBS 0.355013f
C644 VN.n4 VSUBS 0.375369f
C645 VN.n5 VSUBS 0.073872f
C646 VN.n6 VSUBS 0.105277f
C647 VN.n7 VSUBS 0.052892f
C648 VN.n8 VSUBS 0.052892f
C649 VN.n9 VSUBS 0.052892f
C650 VN.n10 VSUBS 0.103708f
C651 VN.n11 VSUBS 0.076778f
C652 VN.n12 VSUBS 0.397836f
C653 VN.n13 VSUBS 0.075026f
C654 VN.n14 VSUBS 0.069728f
C655 VN.t3 VSUBS 0.465237f
C656 VN.n15 VSUBS 0.042871f
C657 VN.n16 VSUBS 0.450168f
C658 VN.t0 VSUBS 0.465237f
C659 VN.t2 VSUBS 0.792499f
C660 VN.n17 VSUBS 0.355013f
C661 VN.n18 VSUBS 0.375369f
C662 VN.n19 VSUBS 0.073872f
C663 VN.n20 VSUBS 0.105277f
C664 VN.n21 VSUBS 0.052892f
C665 VN.n22 VSUBS 0.052892f
C666 VN.n23 VSUBS 0.052892f
C667 VN.n24 VSUBS 0.103708f
C668 VN.n25 VSUBS 0.076778f
C669 VN.n26 VSUBS 0.397836f
C670 VN.n27 VSUBS 2.03596f
.ends

