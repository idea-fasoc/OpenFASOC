* NGSPICE file created from diff_pair_sample_0179.ext - technology: sky130A

.subckt diff_pair_sample_0179 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n3490_n4058# sky130_fd_pr__pfet_01v8 ad=6.0255 pd=31.68 as=0 ps=0 w=15.45 l=2.82
X1 B.t8 B.t6 B.t7 w_n3490_n4058# sky130_fd_pr__pfet_01v8 ad=6.0255 pd=31.68 as=0 ps=0 w=15.45 l=2.82
X2 VDD1.t5 VP.t0 VTAIL.t10 w_n3490_n4058# sky130_fd_pr__pfet_01v8 ad=2.54925 pd=15.78 as=6.0255 ps=31.68 w=15.45 l=2.82
X3 VTAIL.t3 VN.t0 VDD2.t5 w_n3490_n4058# sky130_fd_pr__pfet_01v8 ad=2.54925 pd=15.78 as=2.54925 ps=15.78 w=15.45 l=2.82
X4 VDD1.t4 VP.t1 VTAIL.t8 w_n3490_n4058# sky130_fd_pr__pfet_01v8 ad=6.0255 pd=31.68 as=2.54925 ps=15.78 w=15.45 l=2.82
X5 B.t5 B.t3 B.t4 w_n3490_n4058# sky130_fd_pr__pfet_01v8 ad=6.0255 pd=31.68 as=0 ps=0 w=15.45 l=2.82
X6 VDD2.t4 VN.t1 VTAIL.t5 w_n3490_n4058# sky130_fd_pr__pfet_01v8 ad=6.0255 pd=31.68 as=2.54925 ps=15.78 w=15.45 l=2.82
X7 VDD2.t3 VN.t2 VTAIL.t1 w_n3490_n4058# sky130_fd_pr__pfet_01v8 ad=2.54925 pd=15.78 as=6.0255 ps=31.68 w=15.45 l=2.82
X8 VDD1.t3 VP.t2 VTAIL.t6 w_n3490_n4058# sky130_fd_pr__pfet_01v8 ad=6.0255 pd=31.68 as=2.54925 ps=15.78 w=15.45 l=2.82
X9 VTAIL.t7 VP.t3 VDD1.t2 w_n3490_n4058# sky130_fd_pr__pfet_01v8 ad=2.54925 pd=15.78 as=2.54925 ps=15.78 w=15.45 l=2.82
X10 VTAIL.t11 VP.t4 VDD1.t1 w_n3490_n4058# sky130_fd_pr__pfet_01v8 ad=2.54925 pd=15.78 as=2.54925 ps=15.78 w=15.45 l=2.82
X11 VDD2.t2 VN.t3 VTAIL.t0 w_n3490_n4058# sky130_fd_pr__pfet_01v8 ad=6.0255 pd=31.68 as=2.54925 ps=15.78 w=15.45 l=2.82
X12 B.t2 B.t0 B.t1 w_n3490_n4058# sky130_fd_pr__pfet_01v8 ad=6.0255 pd=31.68 as=0 ps=0 w=15.45 l=2.82
X13 VDD2.t1 VN.t4 VTAIL.t2 w_n3490_n4058# sky130_fd_pr__pfet_01v8 ad=2.54925 pd=15.78 as=6.0255 ps=31.68 w=15.45 l=2.82
X14 VTAIL.t4 VN.t5 VDD2.t0 w_n3490_n4058# sky130_fd_pr__pfet_01v8 ad=2.54925 pd=15.78 as=2.54925 ps=15.78 w=15.45 l=2.82
X15 VDD1.t0 VP.t5 VTAIL.t9 w_n3490_n4058# sky130_fd_pr__pfet_01v8 ad=2.54925 pd=15.78 as=6.0255 ps=31.68 w=15.45 l=2.82
R0 B.n589 B.n588 585
R1 B.n590 B.n85 585
R2 B.n592 B.n591 585
R3 B.n593 B.n84 585
R4 B.n595 B.n594 585
R5 B.n596 B.n83 585
R6 B.n598 B.n597 585
R7 B.n599 B.n82 585
R8 B.n601 B.n600 585
R9 B.n602 B.n81 585
R10 B.n604 B.n603 585
R11 B.n605 B.n80 585
R12 B.n607 B.n606 585
R13 B.n608 B.n79 585
R14 B.n610 B.n609 585
R15 B.n611 B.n78 585
R16 B.n613 B.n612 585
R17 B.n614 B.n77 585
R18 B.n616 B.n615 585
R19 B.n617 B.n76 585
R20 B.n619 B.n618 585
R21 B.n620 B.n75 585
R22 B.n622 B.n621 585
R23 B.n623 B.n74 585
R24 B.n625 B.n624 585
R25 B.n626 B.n73 585
R26 B.n628 B.n627 585
R27 B.n629 B.n72 585
R28 B.n631 B.n630 585
R29 B.n632 B.n71 585
R30 B.n634 B.n633 585
R31 B.n635 B.n70 585
R32 B.n637 B.n636 585
R33 B.n638 B.n69 585
R34 B.n640 B.n639 585
R35 B.n641 B.n68 585
R36 B.n643 B.n642 585
R37 B.n644 B.n67 585
R38 B.n646 B.n645 585
R39 B.n647 B.n66 585
R40 B.n649 B.n648 585
R41 B.n650 B.n65 585
R42 B.n652 B.n651 585
R43 B.n653 B.n64 585
R44 B.n655 B.n654 585
R45 B.n656 B.n63 585
R46 B.n658 B.n657 585
R47 B.n659 B.n62 585
R48 B.n661 B.n660 585
R49 B.n662 B.n61 585
R50 B.n664 B.n663 585
R51 B.n665 B.n58 585
R52 B.n668 B.n667 585
R53 B.n669 B.n57 585
R54 B.n671 B.n670 585
R55 B.n672 B.n56 585
R56 B.n674 B.n673 585
R57 B.n675 B.n55 585
R58 B.n677 B.n676 585
R59 B.n678 B.n51 585
R60 B.n680 B.n679 585
R61 B.n681 B.n50 585
R62 B.n683 B.n682 585
R63 B.n684 B.n49 585
R64 B.n686 B.n685 585
R65 B.n687 B.n48 585
R66 B.n689 B.n688 585
R67 B.n690 B.n47 585
R68 B.n692 B.n691 585
R69 B.n693 B.n46 585
R70 B.n695 B.n694 585
R71 B.n696 B.n45 585
R72 B.n698 B.n697 585
R73 B.n699 B.n44 585
R74 B.n701 B.n700 585
R75 B.n702 B.n43 585
R76 B.n704 B.n703 585
R77 B.n705 B.n42 585
R78 B.n707 B.n706 585
R79 B.n708 B.n41 585
R80 B.n710 B.n709 585
R81 B.n711 B.n40 585
R82 B.n713 B.n712 585
R83 B.n714 B.n39 585
R84 B.n716 B.n715 585
R85 B.n717 B.n38 585
R86 B.n719 B.n718 585
R87 B.n720 B.n37 585
R88 B.n722 B.n721 585
R89 B.n723 B.n36 585
R90 B.n725 B.n724 585
R91 B.n726 B.n35 585
R92 B.n728 B.n727 585
R93 B.n729 B.n34 585
R94 B.n731 B.n730 585
R95 B.n732 B.n33 585
R96 B.n734 B.n733 585
R97 B.n735 B.n32 585
R98 B.n737 B.n736 585
R99 B.n738 B.n31 585
R100 B.n740 B.n739 585
R101 B.n741 B.n30 585
R102 B.n743 B.n742 585
R103 B.n744 B.n29 585
R104 B.n746 B.n745 585
R105 B.n747 B.n28 585
R106 B.n749 B.n748 585
R107 B.n750 B.n27 585
R108 B.n752 B.n751 585
R109 B.n753 B.n26 585
R110 B.n755 B.n754 585
R111 B.n756 B.n25 585
R112 B.n758 B.n757 585
R113 B.n587 B.n86 585
R114 B.n586 B.n585 585
R115 B.n584 B.n87 585
R116 B.n583 B.n582 585
R117 B.n581 B.n88 585
R118 B.n580 B.n579 585
R119 B.n578 B.n89 585
R120 B.n577 B.n576 585
R121 B.n575 B.n90 585
R122 B.n574 B.n573 585
R123 B.n572 B.n91 585
R124 B.n571 B.n570 585
R125 B.n569 B.n92 585
R126 B.n568 B.n567 585
R127 B.n566 B.n93 585
R128 B.n565 B.n564 585
R129 B.n563 B.n94 585
R130 B.n562 B.n561 585
R131 B.n560 B.n95 585
R132 B.n559 B.n558 585
R133 B.n557 B.n96 585
R134 B.n556 B.n555 585
R135 B.n554 B.n97 585
R136 B.n553 B.n552 585
R137 B.n551 B.n98 585
R138 B.n550 B.n549 585
R139 B.n548 B.n99 585
R140 B.n547 B.n546 585
R141 B.n545 B.n100 585
R142 B.n544 B.n543 585
R143 B.n542 B.n101 585
R144 B.n541 B.n540 585
R145 B.n539 B.n102 585
R146 B.n538 B.n537 585
R147 B.n536 B.n103 585
R148 B.n535 B.n534 585
R149 B.n533 B.n104 585
R150 B.n532 B.n531 585
R151 B.n530 B.n105 585
R152 B.n529 B.n528 585
R153 B.n527 B.n106 585
R154 B.n526 B.n525 585
R155 B.n524 B.n107 585
R156 B.n523 B.n522 585
R157 B.n521 B.n108 585
R158 B.n520 B.n519 585
R159 B.n518 B.n109 585
R160 B.n517 B.n516 585
R161 B.n515 B.n110 585
R162 B.n514 B.n513 585
R163 B.n512 B.n111 585
R164 B.n511 B.n510 585
R165 B.n509 B.n112 585
R166 B.n508 B.n507 585
R167 B.n506 B.n113 585
R168 B.n505 B.n504 585
R169 B.n503 B.n114 585
R170 B.n502 B.n501 585
R171 B.n500 B.n115 585
R172 B.n499 B.n498 585
R173 B.n497 B.n116 585
R174 B.n496 B.n495 585
R175 B.n494 B.n117 585
R176 B.n493 B.n492 585
R177 B.n491 B.n118 585
R178 B.n490 B.n489 585
R179 B.n488 B.n119 585
R180 B.n487 B.n486 585
R181 B.n485 B.n120 585
R182 B.n484 B.n483 585
R183 B.n482 B.n121 585
R184 B.n481 B.n480 585
R185 B.n479 B.n122 585
R186 B.n478 B.n477 585
R187 B.n476 B.n123 585
R188 B.n475 B.n474 585
R189 B.n473 B.n124 585
R190 B.n472 B.n471 585
R191 B.n470 B.n125 585
R192 B.n469 B.n468 585
R193 B.n467 B.n126 585
R194 B.n466 B.n465 585
R195 B.n464 B.n127 585
R196 B.n463 B.n462 585
R197 B.n461 B.n128 585
R198 B.n460 B.n459 585
R199 B.n458 B.n129 585
R200 B.n457 B.n456 585
R201 B.n455 B.n130 585
R202 B.n454 B.n453 585
R203 B.n452 B.n131 585
R204 B.n279 B.n278 585
R205 B.n280 B.n189 585
R206 B.n282 B.n281 585
R207 B.n283 B.n188 585
R208 B.n285 B.n284 585
R209 B.n286 B.n187 585
R210 B.n288 B.n287 585
R211 B.n289 B.n186 585
R212 B.n291 B.n290 585
R213 B.n292 B.n185 585
R214 B.n294 B.n293 585
R215 B.n295 B.n184 585
R216 B.n297 B.n296 585
R217 B.n298 B.n183 585
R218 B.n300 B.n299 585
R219 B.n301 B.n182 585
R220 B.n303 B.n302 585
R221 B.n304 B.n181 585
R222 B.n306 B.n305 585
R223 B.n307 B.n180 585
R224 B.n309 B.n308 585
R225 B.n310 B.n179 585
R226 B.n312 B.n311 585
R227 B.n313 B.n178 585
R228 B.n315 B.n314 585
R229 B.n316 B.n177 585
R230 B.n318 B.n317 585
R231 B.n319 B.n176 585
R232 B.n321 B.n320 585
R233 B.n322 B.n175 585
R234 B.n324 B.n323 585
R235 B.n325 B.n174 585
R236 B.n327 B.n326 585
R237 B.n328 B.n173 585
R238 B.n330 B.n329 585
R239 B.n331 B.n172 585
R240 B.n333 B.n332 585
R241 B.n334 B.n171 585
R242 B.n336 B.n335 585
R243 B.n337 B.n170 585
R244 B.n339 B.n338 585
R245 B.n340 B.n169 585
R246 B.n342 B.n341 585
R247 B.n343 B.n168 585
R248 B.n345 B.n344 585
R249 B.n346 B.n167 585
R250 B.n348 B.n347 585
R251 B.n349 B.n166 585
R252 B.n351 B.n350 585
R253 B.n352 B.n165 585
R254 B.n354 B.n353 585
R255 B.n355 B.n162 585
R256 B.n358 B.n357 585
R257 B.n359 B.n161 585
R258 B.n361 B.n360 585
R259 B.n362 B.n160 585
R260 B.n364 B.n363 585
R261 B.n365 B.n159 585
R262 B.n367 B.n366 585
R263 B.n368 B.n158 585
R264 B.n373 B.n372 585
R265 B.n374 B.n157 585
R266 B.n376 B.n375 585
R267 B.n377 B.n156 585
R268 B.n379 B.n378 585
R269 B.n380 B.n155 585
R270 B.n382 B.n381 585
R271 B.n383 B.n154 585
R272 B.n385 B.n384 585
R273 B.n386 B.n153 585
R274 B.n388 B.n387 585
R275 B.n389 B.n152 585
R276 B.n391 B.n390 585
R277 B.n392 B.n151 585
R278 B.n394 B.n393 585
R279 B.n395 B.n150 585
R280 B.n397 B.n396 585
R281 B.n398 B.n149 585
R282 B.n400 B.n399 585
R283 B.n401 B.n148 585
R284 B.n403 B.n402 585
R285 B.n404 B.n147 585
R286 B.n406 B.n405 585
R287 B.n407 B.n146 585
R288 B.n409 B.n408 585
R289 B.n410 B.n145 585
R290 B.n412 B.n411 585
R291 B.n413 B.n144 585
R292 B.n415 B.n414 585
R293 B.n416 B.n143 585
R294 B.n418 B.n417 585
R295 B.n419 B.n142 585
R296 B.n421 B.n420 585
R297 B.n422 B.n141 585
R298 B.n424 B.n423 585
R299 B.n425 B.n140 585
R300 B.n427 B.n426 585
R301 B.n428 B.n139 585
R302 B.n430 B.n429 585
R303 B.n431 B.n138 585
R304 B.n433 B.n432 585
R305 B.n434 B.n137 585
R306 B.n436 B.n435 585
R307 B.n437 B.n136 585
R308 B.n439 B.n438 585
R309 B.n440 B.n135 585
R310 B.n442 B.n441 585
R311 B.n443 B.n134 585
R312 B.n445 B.n444 585
R313 B.n446 B.n133 585
R314 B.n448 B.n447 585
R315 B.n449 B.n132 585
R316 B.n451 B.n450 585
R317 B.n277 B.n190 585
R318 B.n276 B.n275 585
R319 B.n274 B.n191 585
R320 B.n273 B.n272 585
R321 B.n271 B.n192 585
R322 B.n270 B.n269 585
R323 B.n268 B.n193 585
R324 B.n267 B.n266 585
R325 B.n265 B.n194 585
R326 B.n264 B.n263 585
R327 B.n262 B.n195 585
R328 B.n261 B.n260 585
R329 B.n259 B.n196 585
R330 B.n258 B.n257 585
R331 B.n256 B.n197 585
R332 B.n255 B.n254 585
R333 B.n253 B.n198 585
R334 B.n252 B.n251 585
R335 B.n250 B.n199 585
R336 B.n249 B.n248 585
R337 B.n247 B.n200 585
R338 B.n246 B.n245 585
R339 B.n244 B.n201 585
R340 B.n243 B.n242 585
R341 B.n241 B.n202 585
R342 B.n240 B.n239 585
R343 B.n238 B.n203 585
R344 B.n237 B.n236 585
R345 B.n235 B.n204 585
R346 B.n234 B.n233 585
R347 B.n232 B.n205 585
R348 B.n231 B.n230 585
R349 B.n229 B.n206 585
R350 B.n228 B.n227 585
R351 B.n226 B.n207 585
R352 B.n225 B.n224 585
R353 B.n223 B.n208 585
R354 B.n222 B.n221 585
R355 B.n220 B.n209 585
R356 B.n219 B.n218 585
R357 B.n217 B.n210 585
R358 B.n216 B.n215 585
R359 B.n214 B.n211 585
R360 B.n213 B.n212 585
R361 B.n2 B.n0 585
R362 B.n825 B.n1 585
R363 B.n824 B.n823 585
R364 B.n822 B.n3 585
R365 B.n821 B.n820 585
R366 B.n819 B.n4 585
R367 B.n818 B.n817 585
R368 B.n816 B.n5 585
R369 B.n815 B.n814 585
R370 B.n813 B.n6 585
R371 B.n812 B.n811 585
R372 B.n810 B.n7 585
R373 B.n809 B.n808 585
R374 B.n807 B.n8 585
R375 B.n806 B.n805 585
R376 B.n804 B.n9 585
R377 B.n803 B.n802 585
R378 B.n801 B.n10 585
R379 B.n800 B.n799 585
R380 B.n798 B.n11 585
R381 B.n797 B.n796 585
R382 B.n795 B.n12 585
R383 B.n794 B.n793 585
R384 B.n792 B.n13 585
R385 B.n791 B.n790 585
R386 B.n789 B.n14 585
R387 B.n788 B.n787 585
R388 B.n786 B.n15 585
R389 B.n785 B.n784 585
R390 B.n783 B.n16 585
R391 B.n782 B.n781 585
R392 B.n780 B.n17 585
R393 B.n779 B.n778 585
R394 B.n777 B.n18 585
R395 B.n776 B.n775 585
R396 B.n774 B.n19 585
R397 B.n773 B.n772 585
R398 B.n771 B.n20 585
R399 B.n770 B.n769 585
R400 B.n768 B.n21 585
R401 B.n767 B.n766 585
R402 B.n765 B.n22 585
R403 B.n764 B.n763 585
R404 B.n762 B.n23 585
R405 B.n761 B.n760 585
R406 B.n759 B.n24 585
R407 B.n827 B.n826 585
R408 B.n279 B.n190 535.745
R409 B.n759 B.n758 535.745
R410 B.n452 B.n451 535.745
R411 B.n589 B.n86 535.745
R412 B.n369 B.t11 498.829
R413 B.n59 B.t1 498.829
R414 B.n163 B.t5 498.829
R415 B.n52 B.t7 498.829
R416 B.n370 B.t10 437.738
R417 B.n60 B.t2 437.738
R418 B.n164 B.t4 437.738
R419 B.n53 B.t8 437.738
R420 B.n369 B.t9 340.394
R421 B.n163 B.t3 340.394
R422 B.n52 B.t6 340.394
R423 B.n59 B.t0 340.394
R424 B.n275 B.n190 163.367
R425 B.n275 B.n274 163.367
R426 B.n274 B.n273 163.367
R427 B.n273 B.n192 163.367
R428 B.n269 B.n192 163.367
R429 B.n269 B.n268 163.367
R430 B.n268 B.n267 163.367
R431 B.n267 B.n194 163.367
R432 B.n263 B.n194 163.367
R433 B.n263 B.n262 163.367
R434 B.n262 B.n261 163.367
R435 B.n261 B.n196 163.367
R436 B.n257 B.n196 163.367
R437 B.n257 B.n256 163.367
R438 B.n256 B.n255 163.367
R439 B.n255 B.n198 163.367
R440 B.n251 B.n198 163.367
R441 B.n251 B.n250 163.367
R442 B.n250 B.n249 163.367
R443 B.n249 B.n200 163.367
R444 B.n245 B.n200 163.367
R445 B.n245 B.n244 163.367
R446 B.n244 B.n243 163.367
R447 B.n243 B.n202 163.367
R448 B.n239 B.n202 163.367
R449 B.n239 B.n238 163.367
R450 B.n238 B.n237 163.367
R451 B.n237 B.n204 163.367
R452 B.n233 B.n204 163.367
R453 B.n233 B.n232 163.367
R454 B.n232 B.n231 163.367
R455 B.n231 B.n206 163.367
R456 B.n227 B.n206 163.367
R457 B.n227 B.n226 163.367
R458 B.n226 B.n225 163.367
R459 B.n225 B.n208 163.367
R460 B.n221 B.n208 163.367
R461 B.n221 B.n220 163.367
R462 B.n220 B.n219 163.367
R463 B.n219 B.n210 163.367
R464 B.n215 B.n210 163.367
R465 B.n215 B.n214 163.367
R466 B.n214 B.n213 163.367
R467 B.n213 B.n2 163.367
R468 B.n826 B.n2 163.367
R469 B.n826 B.n825 163.367
R470 B.n825 B.n824 163.367
R471 B.n824 B.n3 163.367
R472 B.n820 B.n3 163.367
R473 B.n820 B.n819 163.367
R474 B.n819 B.n818 163.367
R475 B.n818 B.n5 163.367
R476 B.n814 B.n5 163.367
R477 B.n814 B.n813 163.367
R478 B.n813 B.n812 163.367
R479 B.n812 B.n7 163.367
R480 B.n808 B.n7 163.367
R481 B.n808 B.n807 163.367
R482 B.n807 B.n806 163.367
R483 B.n806 B.n9 163.367
R484 B.n802 B.n9 163.367
R485 B.n802 B.n801 163.367
R486 B.n801 B.n800 163.367
R487 B.n800 B.n11 163.367
R488 B.n796 B.n11 163.367
R489 B.n796 B.n795 163.367
R490 B.n795 B.n794 163.367
R491 B.n794 B.n13 163.367
R492 B.n790 B.n13 163.367
R493 B.n790 B.n789 163.367
R494 B.n789 B.n788 163.367
R495 B.n788 B.n15 163.367
R496 B.n784 B.n15 163.367
R497 B.n784 B.n783 163.367
R498 B.n783 B.n782 163.367
R499 B.n782 B.n17 163.367
R500 B.n778 B.n17 163.367
R501 B.n778 B.n777 163.367
R502 B.n777 B.n776 163.367
R503 B.n776 B.n19 163.367
R504 B.n772 B.n19 163.367
R505 B.n772 B.n771 163.367
R506 B.n771 B.n770 163.367
R507 B.n770 B.n21 163.367
R508 B.n766 B.n21 163.367
R509 B.n766 B.n765 163.367
R510 B.n765 B.n764 163.367
R511 B.n764 B.n23 163.367
R512 B.n760 B.n23 163.367
R513 B.n760 B.n759 163.367
R514 B.n280 B.n279 163.367
R515 B.n281 B.n280 163.367
R516 B.n281 B.n188 163.367
R517 B.n285 B.n188 163.367
R518 B.n286 B.n285 163.367
R519 B.n287 B.n286 163.367
R520 B.n287 B.n186 163.367
R521 B.n291 B.n186 163.367
R522 B.n292 B.n291 163.367
R523 B.n293 B.n292 163.367
R524 B.n293 B.n184 163.367
R525 B.n297 B.n184 163.367
R526 B.n298 B.n297 163.367
R527 B.n299 B.n298 163.367
R528 B.n299 B.n182 163.367
R529 B.n303 B.n182 163.367
R530 B.n304 B.n303 163.367
R531 B.n305 B.n304 163.367
R532 B.n305 B.n180 163.367
R533 B.n309 B.n180 163.367
R534 B.n310 B.n309 163.367
R535 B.n311 B.n310 163.367
R536 B.n311 B.n178 163.367
R537 B.n315 B.n178 163.367
R538 B.n316 B.n315 163.367
R539 B.n317 B.n316 163.367
R540 B.n317 B.n176 163.367
R541 B.n321 B.n176 163.367
R542 B.n322 B.n321 163.367
R543 B.n323 B.n322 163.367
R544 B.n323 B.n174 163.367
R545 B.n327 B.n174 163.367
R546 B.n328 B.n327 163.367
R547 B.n329 B.n328 163.367
R548 B.n329 B.n172 163.367
R549 B.n333 B.n172 163.367
R550 B.n334 B.n333 163.367
R551 B.n335 B.n334 163.367
R552 B.n335 B.n170 163.367
R553 B.n339 B.n170 163.367
R554 B.n340 B.n339 163.367
R555 B.n341 B.n340 163.367
R556 B.n341 B.n168 163.367
R557 B.n345 B.n168 163.367
R558 B.n346 B.n345 163.367
R559 B.n347 B.n346 163.367
R560 B.n347 B.n166 163.367
R561 B.n351 B.n166 163.367
R562 B.n352 B.n351 163.367
R563 B.n353 B.n352 163.367
R564 B.n353 B.n162 163.367
R565 B.n358 B.n162 163.367
R566 B.n359 B.n358 163.367
R567 B.n360 B.n359 163.367
R568 B.n360 B.n160 163.367
R569 B.n364 B.n160 163.367
R570 B.n365 B.n364 163.367
R571 B.n366 B.n365 163.367
R572 B.n366 B.n158 163.367
R573 B.n373 B.n158 163.367
R574 B.n374 B.n373 163.367
R575 B.n375 B.n374 163.367
R576 B.n375 B.n156 163.367
R577 B.n379 B.n156 163.367
R578 B.n380 B.n379 163.367
R579 B.n381 B.n380 163.367
R580 B.n381 B.n154 163.367
R581 B.n385 B.n154 163.367
R582 B.n386 B.n385 163.367
R583 B.n387 B.n386 163.367
R584 B.n387 B.n152 163.367
R585 B.n391 B.n152 163.367
R586 B.n392 B.n391 163.367
R587 B.n393 B.n392 163.367
R588 B.n393 B.n150 163.367
R589 B.n397 B.n150 163.367
R590 B.n398 B.n397 163.367
R591 B.n399 B.n398 163.367
R592 B.n399 B.n148 163.367
R593 B.n403 B.n148 163.367
R594 B.n404 B.n403 163.367
R595 B.n405 B.n404 163.367
R596 B.n405 B.n146 163.367
R597 B.n409 B.n146 163.367
R598 B.n410 B.n409 163.367
R599 B.n411 B.n410 163.367
R600 B.n411 B.n144 163.367
R601 B.n415 B.n144 163.367
R602 B.n416 B.n415 163.367
R603 B.n417 B.n416 163.367
R604 B.n417 B.n142 163.367
R605 B.n421 B.n142 163.367
R606 B.n422 B.n421 163.367
R607 B.n423 B.n422 163.367
R608 B.n423 B.n140 163.367
R609 B.n427 B.n140 163.367
R610 B.n428 B.n427 163.367
R611 B.n429 B.n428 163.367
R612 B.n429 B.n138 163.367
R613 B.n433 B.n138 163.367
R614 B.n434 B.n433 163.367
R615 B.n435 B.n434 163.367
R616 B.n435 B.n136 163.367
R617 B.n439 B.n136 163.367
R618 B.n440 B.n439 163.367
R619 B.n441 B.n440 163.367
R620 B.n441 B.n134 163.367
R621 B.n445 B.n134 163.367
R622 B.n446 B.n445 163.367
R623 B.n447 B.n446 163.367
R624 B.n447 B.n132 163.367
R625 B.n451 B.n132 163.367
R626 B.n453 B.n452 163.367
R627 B.n453 B.n130 163.367
R628 B.n457 B.n130 163.367
R629 B.n458 B.n457 163.367
R630 B.n459 B.n458 163.367
R631 B.n459 B.n128 163.367
R632 B.n463 B.n128 163.367
R633 B.n464 B.n463 163.367
R634 B.n465 B.n464 163.367
R635 B.n465 B.n126 163.367
R636 B.n469 B.n126 163.367
R637 B.n470 B.n469 163.367
R638 B.n471 B.n470 163.367
R639 B.n471 B.n124 163.367
R640 B.n475 B.n124 163.367
R641 B.n476 B.n475 163.367
R642 B.n477 B.n476 163.367
R643 B.n477 B.n122 163.367
R644 B.n481 B.n122 163.367
R645 B.n482 B.n481 163.367
R646 B.n483 B.n482 163.367
R647 B.n483 B.n120 163.367
R648 B.n487 B.n120 163.367
R649 B.n488 B.n487 163.367
R650 B.n489 B.n488 163.367
R651 B.n489 B.n118 163.367
R652 B.n493 B.n118 163.367
R653 B.n494 B.n493 163.367
R654 B.n495 B.n494 163.367
R655 B.n495 B.n116 163.367
R656 B.n499 B.n116 163.367
R657 B.n500 B.n499 163.367
R658 B.n501 B.n500 163.367
R659 B.n501 B.n114 163.367
R660 B.n505 B.n114 163.367
R661 B.n506 B.n505 163.367
R662 B.n507 B.n506 163.367
R663 B.n507 B.n112 163.367
R664 B.n511 B.n112 163.367
R665 B.n512 B.n511 163.367
R666 B.n513 B.n512 163.367
R667 B.n513 B.n110 163.367
R668 B.n517 B.n110 163.367
R669 B.n518 B.n517 163.367
R670 B.n519 B.n518 163.367
R671 B.n519 B.n108 163.367
R672 B.n523 B.n108 163.367
R673 B.n524 B.n523 163.367
R674 B.n525 B.n524 163.367
R675 B.n525 B.n106 163.367
R676 B.n529 B.n106 163.367
R677 B.n530 B.n529 163.367
R678 B.n531 B.n530 163.367
R679 B.n531 B.n104 163.367
R680 B.n535 B.n104 163.367
R681 B.n536 B.n535 163.367
R682 B.n537 B.n536 163.367
R683 B.n537 B.n102 163.367
R684 B.n541 B.n102 163.367
R685 B.n542 B.n541 163.367
R686 B.n543 B.n542 163.367
R687 B.n543 B.n100 163.367
R688 B.n547 B.n100 163.367
R689 B.n548 B.n547 163.367
R690 B.n549 B.n548 163.367
R691 B.n549 B.n98 163.367
R692 B.n553 B.n98 163.367
R693 B.n554 B.n553 163.367
R694 B.n555 B.n554 163.367
R695 B.n555 B.n96 163.367
R696 B.n559 B.n96 163.367
R697 B.n560 B.n559 163.367
R698 B.n561 B.n560 163.367
R699 B.n561 B.n94 163.367
R700 B.n565 B.n94 163.367
R701 B.n566 B.n565 163.367
R702 B.n567 B.n566 163.367
R703 B.n567 B.n92 163.367
R704 B.n571 B.n92 163.367
R705 B.n572 B.n571 163.367
R706 B.n573 B.n572 163.367
R707 B.n573 B.n90 163.367
R708 B.n577 B.n90 163.367
R709 B.n578 B.n577 163.367
R710 B.n579 B.n578 163.367
R711 B.n579 B.n88 163.367
R712 B.n583 B.n88 163.367
R713 B.n584 B.n583 163.367
R714 B.n585 B.n584 163.367
R715 B.n585 B.n86 163.367
R716 B.n758 B.n25 163.367
R717 B.n754 B.n25 163.367
R718 B.n754 B.n753 163.367
R719 B.n753 B.n752 163.367
R720 B.n752 B.n27 163.367
R721 B.n748 B.n27 163.367
R722 B.n748 B.n747 163.367
R723 B.n747 B.n746 163.367
R724 B.n746 B.n29 163.367
R725 B.n742 B.n29 163.367
R726 B.n742 B.n741 163.367
R727 B.n741 B.n740 163.367
R728 B.n740 B.n31 163.367
R729 B.n736 B.n31 163.367
R730 B.n736 B.n735 163.367
R731 B.n735 B.n734 163.367
R732 B.n734 B.n33 163.367
R733 B.n730 B.n33 163.367
R734 B.n730 B.n729 163.367
R735 B.n729 B.n728 163.367
R736 B.n728 B.n35 163.367
R737 B.n724 B.n35 163.367
R738 B.n724 B.n723 163.367
R739 B.n723 B.n722 163.367
R740 B.n722 B.n37 163.367
R741 B.n718 B.n37 163.367
R742 B.n718 B.n717 163.367
R743 B.n717 B.n716 163.367
R744 B.n716 B.n39 163.367
R745 B.n712 B.n39 163.367
R746 B.n712 B.n711 163.367
R747 B.n711 B.n710 163.367
R748 B.n710 B.n41 163.367
R749 B.n706 B.n41 163.367
R750 B.n706 B.n705 163.367
R751 B.n705 B.n704 163.367
R752 B.n704 B.n43 163.367
R753 B.n700 B.n43 163.367
R754 B.n700 B.n699 163.367
R755 B.n699 B.n698 163.367
R756 B.n698 B.n45 163.367
R757 B.n694 B.n45 163.367
R758 B.n694 B.n693 163.367
R759 B.n693 B.n692 163.367
R760 B.n692 B.n47 163.367
R761 B.n688 B.n47 163.367
R762 B.n688 B.n687 163.367
R763 B.n687 B.n686 163.367
R764 B.n686 B.n49 163.367
R765 B.n682 B.n49 163.367
R766 B.n682 B.n681 163.367
R767 B.n681 B.n680 163.367
R768 B.n680 B.n51 163.367
R769 B.n676 B.n51 163.367
R770 B.n676 B.n675 163.367
R771 B.n675 B.n674 163.367
R772 B.n674 B.n56 163.367
R773 B.n670 B.n56 163.367
R774 B.n670 B.n669 163.367
R775 B.n669 B.n668 163.367
R776 B.n668 B.n58 163.367
R777 B.n663 B.n58 163.367
R778 B.n663 B.n662 163.367
R779 B.n662 B.n661 163.367
R780 B.n661 B.n62 163.367
R781 B.n657 B.n62 163.367
R782 B.n657 B.n656 163.367
R783 B.n656 B.n655 163.367
R784 B.n655 B.n64 163.367
R785 B.n651 B.n64 163.367
R786 B.n651 B.n650 163.367
R787 B.n650 B.n649 163.367
R788 B.n649 B.n66 163.367
R789 B.n645 B.n66 163.367
R790 B.n645 B.n644 163.367
R791 B.n644 B.n643 163.367
R792 B.n643 B.n68 163.367
R793 B.n639 B.n68 163.367
R794 B.n639 B.n638 163.367
R795 B.n638 B.n637 163.367
R796 B.n637 B.n70 163.367
R797 B.n633 B.n70 163.367
R798 B.n633 B.n632 163.367
R799 B.n632 B.n631 163.367
R800 B.n631 B.n72 163.367
R801 B.n627 B.n72 163.367
R802 B.n627 B.n626 163.367
R803 B.n626 B.n625 163.367
R804 B.n625 B.n74 163.367
R805 B.n621 B.n74 163.367
R806 B.n621 B.n620 163.367
R807 B.n620 B.n619 163.367
R808 B.n619 B.n76 163.367
R809 B.n615 B.n76 163.367
R810 B.n615 B.n614 163.367
R811 B.n614 B.n613 163.367
R812 B.n613 B.n78 163.367
R813 B.n609 B.n78 163.367
R814 B.n609 B.n608 163.367
R815 B.n608 B.n607 163.367
R816 B.n607 B.n80 163.367
R817 B.n603 B.n80 163.367
R818 B.n603 B.n602 163.367
R819 B.n602 B.n601 163.367
R820 B.n601 B.n82 163.367
R821 B.n597 B.n82 163.367
R822 B.n597 B.n596 163.367
R823 B.n596 B.n595 163.367
R824 B.n595 B.n84 163.367
R825 B.n591 B.n84 163.367
R826 B.n591 B.n590 163.367
R827 B.n590 B.n589 163.367
R828 B.n370 B.n369 61.0914
R829 B.n164 B.n163 61.0914
R830 B.n53 B.n52 61.0914
R831 B.n60 B.n59 61.0914
R832 B.n371 B.n370 59.5399
R833 B.n356 B.n164 59.5399
R834 B.n54 B.n53 59.5399
R835 B.n666 B.n60 59.5399
R836 B.n588 B.n587 34.8103
R837 B.n757 B.n24 34.8103
R838 B.n450 B.n131 34.8103
R839 B.n278 B.n277 34.8103
R840 B B.n827 18.0485
R841 B.n757 B.n756 10.6151
R842 B.n756 B.n755 10.6151
R843 B.n755 B.n26 10.6151
R844 B.n751 B.n26 10.6151
R845 B.n751 B.n750 10.6151
R846 B.n750 B.n749 10.6151
R847 B.n749 B.n28 10.6151
R848 B.n745 B.n28 10.6151
R849 B.n745 B.n744 10.6151
R850 B.n744 B.n743 10.6151
R851 B.n743 B.n30 10.6151
R852 B.n739 B.n30 10.6151
R853 B.n739 B.n738 10.6151
R854 B.n738 B.n737 10.6151
R855 B.n737 B.n32 10.6151
R856 B.n733 B.n32 10.6151
R857 B.n733 B.n732 10.6151
R858 B.n732 B.n731 10.6151
R859 B.n731 B.n34 10.6151
R860 B.n727 B.n34 10.6151
R861 B.n727 B.n726 10.6151
R862 B.n726 B.n725 10.6151
R863 B.n725 B.n36 10.6151
R864 B.n721 B.n36 10.6151
R865 B.n721 B.n720 10.6151
R866 B.n720 B.n719 10.6151
R867 B.n719 B.n38 10.6151
R868 B.n715 B.n38 10.6151
R869 B.n715 B.n714 10.6151
R870 B.n714 B.n713 10.6151
R871 B.n713 B.n40 10.6151
R872 B.n709 B.n40 10.6151
R873 B.n709 B.n708 10.6151
R874 B.n708 B.n707 10.6151
R875 B.n707 B.n42 10.6151
R876 B.n703 B.n42 10.6151
R877 B.n703 B.n702 10.6151
R878 B.n702 B.n701 10.6151
R879 B.n701 B.n44 10.6151
R880 B.n697 B.n44 10.6151
R881 B.n697 B.n696 10.6151
R882 B.n696 B.n695 10.6151
R883 B.n695 B.n46 10.6151
R884 B.n691 B.n46 10.6151
R885 B.n691 B.n690 10.6151
R886 B.n690 B.n689 10.6151
R887 B.n689 B.n48 10.6151
R888 B.n685 B.n48 10.6151
R889 B.n685 B.n684 10.6151
R890 B.n684 B.n683 10.6151
R891 B.n683 B.n50 10.6151
R892 B.n679 B.n678 10.6151
R893 B.n678 B.n677 10.6151
R894 B.n677 B.n55 10.6151
R895 B.n673 B.n55 10.6151
R896 B.n673 B.n672 10.6151
R897 B.n672 B.n671 10.6151
R898 B.n671 B.n57 10.6151
R899 B.n667 B.n57 10.6151
R900 B.n665 B.n664 10.6151
R901 B.n664 B.n61 10.6151
R902 B.n660 B.n61 10.6151
R903 B.n660 B.n659 10.6151
R904 B.n659 B.n658 10.6151
R905 B.n658 B.n63 10.6151
R906 B.n654 B.n63 10.6151
R907 B.n654 B.n653 10.6151
R908 B.n653 B.n652 10.6151
R909 B.n652 B.n65 10.6151
R910 B.n648 B.n65 10.6151
R911 B.n648 B.n647 10.6151
R912 B.n647 B.n646 10.6151
R913 B.n646 B.n67 10.6151
R914 B.n642 B.n67 10.6151
R915 B.n642 B.n641 10.6151
R916 B.n641 B.n640 10.6151
R917 B.n640 B.n69 10.6151
R918 B.n636 B.n69 10.6151
R919 B.n636 B.n635 10.6151
R920 B.n635 B.n634 10.6151
R921 B.n634 B.n71 10.6151
R922 B.n630 B.n71 10.6151
R923 B.n630 B.n629 10.6151
R924 B.n629 B.n628 10.6151
R925 B.n628 B.n73 10.6151
R926 B.n624 B.n73 10.6151
R927 B.n624 B.n623 10.6151
R928 B.n623 B.n622 10.6151
R929 B.n622 B.n75 10.6151
R930 B.n618 B.n75 10.6151
R931 B.n618 B.n617 10.6151
R932 B.n617 B.n616 10.6151
R933 B.n616 B.n77 10.6151
R934 B.n612 B.n77 10.6151
R935 B.n612 B.n611 10.6151
R936 B.n611 B.n610 10.6151
R937 B.n610 B.n79 10.6151
R938 B.n606 B.n79 10.6151
R939 B.n606 B.n605 10.6151
R940 B.n605 B.n604 10.6151
R941 B.n604 B.n81 10.6151
R942 B.n600 B.n81 10.6151
R943 B.n600 B.n599 10.6151
R944 B.n599 B.n598 10.6151
R945 B.n598 B.n83 10.6151
R946 B.n594 B.n83 10.6151
R947 B.n594 B.n593 10.6151
R948 B.n593 B.n592 10.6151
R949 B.n592 B.n85 10.6151
R950 B.n588 B.n85 10.6151
R951 B.n454 B.n131 10.6151
R952 B.n455 B.n454 10.6151
R953 B.n456 B.n455 10.6151
R954 B.n456 B.n129 10.6151
R955 B.n460 B.n129 10.6151
R956 B.n461 B.n460 10.6151
R957 B.n462 B.n461 10.6151
R958 B.n462 B.n127 10.6151
R959 B.n466 B.n127 10.6151
R960 B.n467 B.n466 10.6151
R961 B.n468 B.n467 10.6151
R962 B.n468 B.n125 10.6151
R963 B.n472 B.n125 10.6151
R964 B.n473 B.n472 10.6151
R965 B.n474 B.n473 10.6151
R966 B.n474 B.n123 10.6151
R967 B.n478 B.n123 10.6151
R968 B.n479 B.n478 10.6151
R969 B.n480 B.n479 10.6151
R970 B.n480 B.n121 10.6151
R971 B.n484 B.n121 10.6151
R972 B.n485 B.n484 10.6151
R973 B.n486 B.n485 10.6151
R974 B.n486 B.n119 10.6151
R975 B.n490 B.n119 10.6151
R976 B.n491 B.n490 10.6151
R977 B.n492 B.n491 10.6151
R978 B.n492 B.n117 10.6151
R979 B.n496 B.n117 10.6151
R980 B.n497 B.n496 10.6151
R981 B.n498 B.n497 10.6151
R982 B.n498 B.n115 10.6151
R983 B.n502 B.n115 10.6151
R984 B.n503 B.n502 10.6151
R985 B.n504 B.n503 10.6151
R986 B.n504 B.n113 10.6151
R987 B.n508 B.n113 10.6151
R988 B.n509 B.n508 10.6151
R989 B.n510 B.n509 10.6151
R990 B.n510 B.n111 10.6151
R991 B.n514 B.n111 10.6151
R992 B.n515 B.n514 10.6151
R993 B.n516 B.n515 10.6151
R994 B.n516 B.n109 10.6151
R995 B.n520 B.n109 10.6151
R996 B.n521 B.n520 10.6151
R997 B.n522 B.n521 10.6151
R998 B.n522 B.n107 10.6151
R999 B.n526 B.n107 10.6151
R1000 B.n527 B.n526 10.6151
R1001 B.n528 B.n527 10.6151
R1002 B.n528 B.n105 10.6151
R1003 B.n532 B.n105 10.6151
R1004 B.n533 B.n532 10.6151
R1005 B.n534 B.n533 10.6151
R1006 B.n534 B.n103 10.6151
R1007 B.n538 B.n103 10.6151
R1008 B.n539 B.n538 10.6151
R1009 B.n540 B.n539 10.6151
R1010 B.n540 B.n101 10.6151
R1011 B.n544 B.n101 10.6151
R1012 B.n545 B.n544 10.6151
R1013 B.n546 B.n545 10.6151
R1014 B.n546 B.n99 10.6151
R1015 B.n550 B.n99 10.6151
R1016 B.n551 B.n550 10.6151
R1017 B.n552 B.n551 10.6151
R1018 B.n552 B.n97 10.6151
R1019 B.n556 B.n97 10.6151
R1020 B.n557 B.n556 10.6151
R1021 B.n558 B.n557 10.6151
R1022 B.n558 B.n95 10.6151
R1023 B.n562 B.n95 10.6151
R1024 B.n563 B.n562 10.6151
R1025 B.n564 B.n563 10.6151
R1026 B.n564 B.n93 10.6151
R1027 B.n568 B.n93 10.6151
R1028 B.n569 B.n568 10.6151
R1029 B.n570 B.n569 10.6151
R1030 B.n570 B.n91 10.6151
R1031 B.n574 B.n91 10.6151
R1032 B.n575 B.n574 10.6151
R1033 B.n576 B.n575 10.6151
R1034 B.n576 B.n89 10.6151
R1035 B.n580 B.n89 10.6151
R1036 B.n581 B.n580 10.6151
R1037 B.n582 B.n581 10.6151
R1038 B.n582 B.n87 10.6151
R1039 B.n586 B.n87 10.6151
R1040 B.n587 B.n586 10.6151
R1041 B.n278 B.n189 10.6151
R1042 B.n282 B.n189 10.6151
R1043 B.n283 B.n282 10.6151
R1044 B.n284 B.n283 10.6151
R1045 B.n284 B.n187 10.6151
R1046 B.n288 B.n187 10.6151
R1047 B.n289 B.n288 10.6151
R1048 B.n290 B.n289 10.6151
R1049 B.n290 B.n185 10.6151
R1050 B.n294 B.n185 10.6151
R1051 B.n295 B.n294 10.6151
R1052 B.n296 B.n295 10.6151
R1053 B.n296 B.n183 10.6151
R1054 B.n300 B.n183 10.6151
R1055 B.n301 B.n300 10.6151
R1056 B.n302 B.n301 10.6151
R1057 B.n302 B.n181 10.6151
R1058 B.n306 B.n181 10.6151
R1059 B.n307 B.n306 10.6151
R1060 B.n308 B.n307 10.6151
R1061 B.n308 B.n179 10.6151
R1062 B.n312 B.n179 10.6151
R1063 B.n313 B.n312 10.6151
R1064 B.n314 B.n313 10.6151
R1065 B.n314 B.n177 10.6151
R1066 B.n318 B.n177 10.6151
R1067 B.n319 B.n318 10.6151
R1068 B.n320 B.n319 10.6151
R1069 B.n320 B.n175 10.6151
R1070 B.n324 B.n175 10.6151
R1071 B.n325 B.n324 10.6151
R1072 B.n326 B.n325 10.6151
R1073 B.n326 B.n173 10.6151
R1074 B.n330 B.n173 10.6151
R1075 B.n331 B.n330 10.6151
R1076 B.n332 B.n331 10.6151
R1077 B.n332 B.n171 10.6151
R1078 B.n336 B.n171 10.6151
R1079 B.n337 B.n336 10.6151
R1080 B.n338 B.n337 10.6151
R1081 B.n338 B.n169 10.6151
R1082 B.n342 B.n169 10.6151
R1083 B.n343 B.n342 10.6151
R1084 B.n344 B.n343 10.6151
R1085 B.n344 B.n167 10.6151
R1086 B.n348 B.n167 10.6151
R1087 B.n349 B.n348 10.6151
R1088 B.n350 B.n349 10.6151
R1089 B.n350 B.n165 10.6151
R1090 B.n354 B.n165 10.6151
R1091 B.n355 B.n354 10.6151
R1092 B.n357 B.n161 10.6151
R1093 B.n361 B.n161 10.6151
R1094 B.n362 B.n361 10.6151
R1095 B.n363 B.n362 10.6151
R1096 B.n363 B.n159 10.6151
R1097 B.n367 B.n159 10.6151
R1098 B.n368 B.n367 10.6151
R1099 B.n372 B.n368 10.6151
R1100 B.n376 B.n157 10.6151
R1101 B.n377 B.n376 10.6151
R1102 B.n378 B.n377 10.6151
R1103 B.n378 B.n155 10.6151
R1104 B.n382 B.n155 10.6151
R1105 B.n383 B.n382 10.6151
R1106 B.n384 B.n383 10.6151
R1107 B.n384 B.n153 10.6151
R1108 B.n388 B.n153 10.6151
R1109 B.n389 B.n388 10.6151
R1110 B.n390 B.n389 10.6151
R1111 B.n390 B.n151 10.6151
R1112 B.n394 B.n151 10.6151
R1113 B.n395 B.n394 10.6151
R1114 B.n396 B.n395 10.6151
R1115 B.n396 B.n149 10.6151
R1116 B.n400 B.n149 10.6151
R1117 B.n401 B.n400 10.6151
R1118 B.n402 B.n401 10.6151
R1119 B.n402 B.n147 10.6151
R1120 B.n406 B.n147 10.6151
R1121 B.n407 B.n406 10.6151
R1122 B.n408 B.n407 10.6151
R1123 B.n408 B.n145 10.6151
R1124 B.n412 B.n145 10.6151
R1125 B.n413 B.n412 10.6151
R1126 B.n414 B.n413 10.6151
R1127 B.n414 B.n143 10.6151
R1128 B.n418 B.n143 10.6151
R1129 B.n419 B.n418 10.6151
R1130 B.n420 B.n419 10.6151
R1131 B.n420 B.n141 10.6151
R1132 B.n424 B.n141 10.6151
R1133 B.n425 B.n424 10.6151
R1134 B.n426 B.n425 10.6151
R1135 B.n426 B.n139 10.6151
R1136 B.n430 B.n139 10.6151
R1137 B.n431 B.n430 10.6151
R1138 B.n432 B.n431 10.6151
R1139 B.n432 B.n137 10.6151
R1140 B.n436 B.n137 10.6151
R1141 B.n437 B.n436 10.6151
R1142 B.n438 B.n437 10.6151
R1143 B.n438 B.n135 10.6151
R1144 B.n442 B.n135 10.6151
R1145 B.n443 B.n442 10.6151
R1146 B.n444 B.n443 10.6151
R1147 B.n444 B.n133 10.6151
R1148 B.n448 B.n133 10.6151
R1149 B.n449 B.n448 10.6151
R1150 B.n450 B.n449 10.6151
R1151 B.n277 B.n276 10.6151
R1152 B.n276 B.n191 10.6151
R1153 B.n272 B.n191 10.6151
R1154 B.n272 B.n271 10.6151
R1155 B.n271 B.n270 10.6151
R1156 B.n270 B.n193 10.6151
R1157 B.n266 B.n193 10.6151
R1158 B.n266 B.n265 10.6151
R1159 B.n265 B.n264 10.6151
R1160 B.n264 B.n195 10.6151
R1161 B.n260 B.n195 10.6151
R1162 B.n260 B.n259 10.6151
R1163 B.n259 B.n258 10.6151
R1164 B.n258 B.n197 10.6151
R1165 B.n254 B.n197 10.6151
R1166 B.n254 B.n253 10.6151
R1167 B.n253 B.n252 10.6151
R1168 B.n252 B.n199 10.6151
R1169 B.n248 B.n199 10.6151
R1170 B.n248 B.n247 10.6151
R1171 B.n247 B.n246 10.6151
R1172 B.n246 B.n201 10.6151
R1173 B.n242 B.n201 10.6151
R1174 B.n242 B.n241 10.6151
R1175 B.n241 B.n240 10.6151
R1176 B.n240 B.n203 10.6151
R1177 B.n236 B.n203 10.6151
R1178 B.n236 B.n235 10.6151
R1179 B.n235 B.n234 10.6151
R1180 B.n234 B.n205 10.6151
R1181 B.n230 B.n205 10.6151
R1182 B.n230 B.n229 10.6151
R1183 B.n229 B.n228 10.6151
R1184 B.n228 B.n207 10.6151
R1185 B.n224 B.n207 10.6151
R1186 B.n224 B.n223 10.6151
R1187 B.n223 B.n222 10.6151
R1188 B.n222 B.n209 10.6151
R1189 B.n218 B.n209 10.6151
R1190 B.n218 B.n217 10.6151
R1191 B.n217 B.n216 10.6151
R1192 B.n216 B.n211 10.6151
R1193 B.n212 B.n211 10.6151
R1194 B.n212 B.n0 10.6151
R1195 B.n823 B.n1 10.6151
R1196 B.n823 B.n822 10.6151
R1197 B.n822 B.n821 10.6151
R1198 B.n821 B.n4 10.6151
R1199 B.n817 B.n4 10.6151
R1200 B.n817 B.n816 10.6151
R1201 B.n816 B.n815 10.6151
R1202 B.n815 B.n6 10.6151
R1203 B.n811 B.n6 10.6151
R1204 B.n811 B.n810 10.6151
R1205 B.n810 B.n809 10.6151
R1206 B.n809 B.n8 10.6151
R1207 B.n805 B.n8 10.6151
R1208 B.n805 B.n804 10.6151
R1209 B.n804 B.n803 10.6151
R1210 B.n803 B.n10 10.6151
R1211 B.n799 B.n10 10.6151
R1212 B.n799 B.n798 10.6151
R1213 B.n798 B.n797 10.6151
R1214 B.n797 B.n12 10.6151
R1215 B.n793 B.n12 10.6151
R1216 B.n793 B.n792 10.6151
R1217 B.n792 B.n791 10.6151
R1218 B.n791 B.n14 10.6151
R1219 B.n787 B.n14 10.6151
R1220 B.n787 B.n786 10.6151
R1221 B.n786 B.n785 10.6151
R1222 B.n785 B.n16 10.6151
R1223 B.n781 B.n16 10.6151
R1224 B.n781 B.n780 10.6151
R1225 B.n780 B.n779 10.6151
R1226 B.n779 B.n18 10.6151
R1227 B.n775 B.n18 10.6151
R1228 B.n775 B.n774 10.6151
R1229 B.n774 B.n773 10.6151
R1230 B.n773 B.n20 10.6151
R1231 B.n769 B.n20 10.6151
R1232 B.n769 B.n768 10.6151
R1233 B.n768 B.n767 10.6151
R1234 B.n767 B.n22 10.6151
R1235 B.n763 B.n22 10.6151
R1236 B.n763 B.n762 10.6151
R1237 B.n762 B.n761 10.6151
R1238 B.n761 B.n24 10.6151
R1239 B.n679 B.n54 6.5566
R1240 B.n667 B.n666 6.5566
R1241 B.n357 B.n356 6.5566
R1242 B.n372 B.n371 6.5566
R1243 B.n54 B.n50 4.05904
R1244 B.n666 B.n665 4.05904
R1245 B.n356 B.n355 4.05904
R1246 B.n371 B.n157 4.05904
R1247 B.n827 B.n0 2.81026
R1248 B.n827 B.n1 2.81026
R1249 VP.n11 VP.t1 163.718
R1250 VP.n13 VP.n10 161.3
R1251 VP.n15 VP.n14 161.3
R1252 VP.n16 VP.n9 161.3
R1253 VP.n18 VP.n17 161.3
R1254 VP.n19 VP.n8 161.3
R1255 VP.n21 VP.n20 161.3
R1256 VP.n43 VP.n42 161.3
R1257 VP.n41 VP.n1 161.3
R1258 VP.n40 VP.n39 161.3
R1259 VP.n38 VP.n2 161.3
R1260 VP.n37 VP.n36 161.3
R1261 VP.n35 VP.n3 161.3
R1262 VP.n33 VP.n32 161.3
R1263 VP.n31 VP.n4 161.3
R1264 VP.n30 VP.n29 161.3
R1265 VP.n28 VP.n5 161.3
R1266 VP.n27 VP.n26 161.3
R1267 VP.n25 VP.n6 161.3
R1268 VP.n23 VP.t2 132.037
R1269 VP.n34 VP.t3 132.037
R1270 VP.n0 VP.t5 132.037
R1271 VP.n7 VP.t0 132.037
R1272 VP.n12 VP.t4 132.037
R1273 VP.n24 VP.n23 70.4938
R1274 VP.n44 VP.n0 70.4938
R1275 VP.n22 VP.n7 70.4938
R1276 VP.n12 VP.n11 61.3922
R1277 VP.n29 VP.n28 56.5193
R1278 VP.n40 VP.n2 56.5193
R1279 VP.n18 VP.n9 56.5193
R1280 VP.n24 VP.n22 52.2228
R1281 VP.n27 VP.n6 24.4675
R1282 VP.n28 VP.n27 24.4675
R1283 VP.n29 VP.n4 24.4675
R1284 VP.n33 VP.n4 24.4675
R1285 VP.n36 VP.n35 24.4675
R1286 VP.n36 VP.n2 24.4675
R1287 VP.n41 VP.n40 24.4675
R1288 VP.n42 VP.n41 24.4675
R1289 VP.n19 VP.n18 24.4675
R1290 VP.n20 VP.n19 24.4675
R1291 VP.n14 VP.n13 24.4675
R1292 VP.n14 VP.n9 24.4675
R1293 VP.n23 VP.n6 19.5741
R1294 VP.n42 VP.n0 19.5741
R1295 VP.n20 VP.n7 19.5741
R1296 VP.n34 VP.n33 12.234
R1297 VP.n35 VP.n34 12.234
R1298 VP.n13 VP.n12 12.234
R1299 VP.n11 VP.n10 5.58426
R1300 VP.n22 VP.n21 0.354971
R1301 VP.n25 VP.n24 0.354971
R1302 VP.n44 VP.n43 0.354971
R1303 VP VP.n44 0.26696
R1304 VP.n15 VP.n10 0.189894
R1305 VP.n16 VP.n15 0.189894
R1306 VP.n17 VP.n16 0.189894
R1307 VP.n17 VP.n8 0.189894
R1308 VP.n21 VP.n8 0.189894
R1309 VP.n26 VP.n25 0.189894
R1310 VP.n26 VP.n5 0.189894
R1311 VP.n30 VP.n5 0.189894
R1312 VP.n31 VP.n30 0.189894
R1313 VP.n32 VP.n31 0.189894
R1314 VP.n32 VP.n3 0.189894
R1315 VP.n37 VP.n3 0.189894
R1316 VP.n38 VP.n37 0.189894
R1317 VP.n39 VP.n38 0.189894
R1318 VP.n39 VP.n1 0.189894
R1319 VP.n43 VP.n1 0.189894
R1320 VTAIL.n346 VTAIL.n266 756.745
R1321 VTAIL.n82 VTAIL.n2 756.745
R1322 VTAIL.n260 VTAIL.n180 756.745
R1323 VTAIL.n172 VTAIL.n92 756.745
R1324 VTAIL.n295 VTAIL.n294 585
R1325 VTAIL.n297 VTAIL.n296 585
R1326 VTAIL.n290 VTAIL.n289 585
R1327 VTAIL.n303 VTAIL.n302 585
R1328 VTAIL.n305 VTAIL.n304 585
R1329 VTAIL.n286 VTAIL.n285 585
R1330 VTAIL.n311 VTAIL.n310 585
R1331 VTAIL.n313 VTAIL.n312 585
R1332 VTAIL.n282 VTAIL.n281 585
R1333 VTAIL.n319 VTAIL.n318 585
R1334 VTAIL.n321 VTAIL.n320 585
R1335 VTAIL.n278 VTAIL.n277 585
R1336 VTAIL.n327 VTAIL.n326 585
R1337 VTAIL.n329 VTAIL.n328 585
R1338 VTAIL.n274 VTAIL.n273 585
R1339 VTAIL.n336 VTAIL.n335 585
R1340 VTAIL.n337 VTAIL.n272 585
R1341 VTAIL.n339 VTAIL.n338 585
R1342 VTAIL.n270 VTAIL.n269 585
R1343 VTAIL.n345 VTAIL.n344 585
R1344 VTAIL.n347 VTAIL.n346 585
R1345 VTAIL.n31 VTAIL.n30 585
R1346 VTAIL.n33 VTAIL.n32 585
R1347 VTAIL.n26 VTAIL.n25 585
R1348 VTAIL.n39 VTAIL.n38 585
R1349 VTAIL.n41 VTAIL.n40 585
R1350 VTAIL.n22 VTAIL.n21 585
R1351 VTAIL.n47 VTAIL.n46 585
R1352 VTAIL.n49 VTAIL.n48 585
R1353 VTAIL.n18 VTAIL.n17 585
R1354 VTAIL.n55 VTAIL.n54 585
R1355 VTAIL.n57 VTAIL.n56 585
R1356 VTAIL.n14 VTAIL.n13 585
R1357 VTAIL.n63 VTAIL.n62 585
R1358 VTAIL.n65 VTAIL.n64 585
R1359 VTAIL.n10 VTAIL.n9 585
R1360 VTAIL.n72 VTAIL.n71 585
R1361 VTAIL.n73 VTAIL.n8 585
R1362 VTAIL.n75 VTAIL.n74 585
R1363 VTAIL.n6 VTAIL.n5 585
R1364 VTAIL.n81 VTAIL.n80 585
R1365 VTAIL.n83 VTAIL.n82 585
R1366 VTAIL.n261 VTAIL.n260 585
R1367 VTAIL.n259 VTAIL.n258 585
R1368 VTAIL.n184 VTAIL.n183 585
R1369 VTAIL.n188 VTAIL.n186 585
R1370 VTAIL.n253 VTAIL.n252 585
R1371 VTAIL.n251 VTAIL.n250 585
R1372 VTAIL.n190 VTAIL.n189 585
R1373 VTAIL.n245 VTAIL.n244 585
R1374 VTAIL.n243 VTAIL.n242 585
R1375 VTAIL.n194 VTAIL.n193 585
R1376 VTAIL.n237 VTAIL.n236 585
R1377 VTAIL.n235 VTAIL.n234 585
R1378 VTAIL.n198 VTAIL.n197 585
R1379 VTAIL.n229 VTAIL.n228 585
R1380 VTAIL.n227 VTAIL.n226 585
R1381 VTAIL.n202 VTAIL.n201 585
R1382 VTAIL.n221 VTAIL.n220 585
R1383 VTAIL.n219 VTAIL.n218 585
R1384 VTAIL.n206 VTAIL.n205 585
R1385 VTAIL.n213 VTAIL.n212 585
R1386 VTAIL.n211 VTAIL.n210 585
R1387 VTAIL.n173 VTAIL.n172 585
R1388 VTAIL.n171 VTAIL.n170 585
R1389 VTAIL.n96 VTAIL.n95 585
R1390 VTAIL.n100 VTAIL.n98 585
R1391 VTAIL.n165 VTAIL.n164 585
R1392 VTAIL.n163 VTAIL.n162 585
R1393 VTAIL.n102 VTAIL.n101 585
R1394 VTAIL.n157 VTAIL.n156 585
R1395 VTAIL.n155 VTAIL.n154 585
R1396 VTAIL.n106 VTAIL.n105 585
R1397 VTAIL.n149 VTAIL.n148 585
R1398 VTAIL.n147 VTAIL.n146 585
R1399 VTAIL.n110 VTAIL.n109 585
R1400 VTAIL.n141 VTAIL.n140 585
R1401 VTAIL.n139 VTAIL.n138 585
R1402 VTAIL.n114 VTAIL.n113 585
R1403 VTAIL.n133 VTAIL.n132 585
R1404 VTAIL.n131 VTAIL.n130 585
R1405 VTAIL.n118 VTAIL.n117 585
R1406 VTAIL.n125 VTAIL.n124 585
R1407 VTAIL.n123 VTAIL.n122 585
R1408 VTAIL.n293 VTAIL.t2 327.466
R1409 VTAIL.n29 VTAIL.t9 327.466
R1410 VTAIL.n209 VTAIL.t10 327.466
R1411 VTAIL.n121 VTAIL.t1 327.466
R1412 VTAIL.n296 VTAIL.n295 171.744
R1413 VTAIL.n296 VTAIL.n289 171.744
R1414 VTAIL.n303 VTAIL.n289 171.744
R1415 VTAIL.n304 VTAIL.n303 171.744
R1416 VTAIL.n304 VTAIL.n285 171.744
R1417 VTAIL.n311 VTAIL.n285 171.744
R1418 VTAIL.n312 VTAIL.n311 171.744
R1419 VTAIL.n312 VTAIL.n281 171.744
R1420 VTAIL.n319 VTAIL.n281 171.744
R1421 VTAIL.n320 VTAIL.n319 171.744
R1422 VTAIL.n320 VTAIL.n277 171.744
R1423 VTAIL.n327 VTAIL.n277 171.744
R1424 VTAIL.n328 VTAIL.n327 171.744
R1425 VTAIL.n328 VTAIL.n273 171.744
R1426 VTAIL.n336 VTAIL.n273 171.744
R1427 VTAIL.n337 VTAIL.n336 171.744
R1428 VTAIL.n338 VTAIL.n337 171.744
R1429 VTAIL.n338 VTAIL.n269 171.744
R1430 VTAIL.n345 VTAIL.n269 171.744
R1431 VTAIL.n346 VTAIL.n345 171.744
R1432 VTAIL.n32 VTAIL.n31 171.744
R1433 VTAIL.n32 VTAIL.n25 171.744
R1434 VTAIL.n39 VTAIL.n25 171.744
R1435 VTAIL.n40 VTAIL.n39 171.744
R1436 VTAIL.n40 VTAIL.n21 171.744
R1437 VTAIL.n47 VTAIL.n21 171.744
R1438 VTAIL.n48 VTAIL.n47 171.744
R1439 VTAIL.n48 VTAIL.n17 171.744
R1440 VTAIL.n55 VTAIL.n17 171.744
R1441 VTAIL.n56 VTAIL.n55 171.744
R1442 VTAIL.n56 VTAIL.n13 171.744
R1443 VTAIL.n63 VTAIL.n13 171.744
R1444 VTAIL.n64 VTAIL.n63 171.744
R1445 VTAIL.n64 VTAIL.n9 171.744
R1446 VTAIL.n72 VTAIL.n9 171.744
R1447 VTAIL.n73 VTAIL.n72 171.744
R1448 VTAIL.n74 VTAIL.n73 171.744
R1449 VTAIL.n74 VTAIL.n5 171.744
R1450 VTAIL.n81 VTAIL.n5 171.744
R1451 VTAIL.n82 VTAIL.n81 171.744
R1452 VTAIL.n260 VTAIL.n259 171.744
R1453 VTAIL.n259 VTAIL.n183 171.744
R1454 VTAIL.n188 VTAIL.n183 171.744
R1455 VTAIL.n252 VTAIL.n188 171.744
R1456 VTAIL.n252 VTAIL.n251 171.744
R1457 VTAIL.n251 VTAIL.n189 171.744
R1458 VTAIL.n244 VTAIL.n189 171.744
R1459 VTAIL.n244 VTAIL.n243 171.744
R1460 VTAIL.n243 VTAIL.n193 171.744
R1461 VTAIL.n236 VTAIL.n193 171.744
R1462 VTAIL.n236 VTAIL.n235 171.744
R1463 VTAIL.n235 VTAIL.n197 171.744
R1464 VTAIL.n228 VTAIL.n197 171.744
R1465 VTAIL.n228 VTAIL.n227 171.744
R1466 VTAIL.n227 VTAIL.n201 171.744
R1467 VTAIL.n220 VTAIL.n201 171.744
R1468 VTAIL.n220 VTAIL.n219 171.744
R1469 VTAIL.n219 VTAIL.n205 171.744
R1470 VTAIL.n212 VTAIL.n205 171.744
R1471 VTAIL.n212 VTAIL.n211 171.744
R1472 VTAIL.n172 VTAIL.n171 171.744
R1473 VTAIL.n171 VTAIL.n95 171.744
R1474 VTAIL.n100 VTAIL.n95 171.744
R1475 VTAIL.n164 VTAIL.n100 171.744
R1476 VTAIL.n164 VTAIL.n163 171.744
R1477 VTAIL.n163 VTAIL.n101 171.744
R1478 VTAIL.n156 VTAIL.n101 171.744
R1479 VTAIL.n156 VTAIL.n155 171.744
R1480 VTAIL.n155 VTAIL.n105 171.744
R1481 VTAIL.n148 VTAIL.n105 171.744
R1482 VTAIL.n148 VTAIL.n147 171.744
R1483 VTAIL.n147 VTAIL.n109 171.744
R1484 VTAIL.n140 VTAIL.n109 171.744
R1485 VTAIL.n140 VTAIL.n139 171.744
R1486 VTAIL.n139 VTAIL.n113 171.744
R1487 VTAIL.n132 VTAIL.n113 171.744
R1488 VTAIL.n132 VTAIL.n131 171.744
R1489 VTAIL.n131 VTAIL.n117 171.744
R1490 VTAIL.n124 VTAIL.n117 171.744
R1491 VTAIL.n124 VTAIL.n123 171.744
R1492 VTAIL.n295 VTAIL.t2 85.8723
R1493 VTAIL.n31 VTAIL.t9 85.8723
R1494 VTAIL.n211 VTAIL.t10 85.8723
R1495 VTAIL.n123 VTAIL.t1 85.8723
R1496 VTAIL.n179 VTAIL.n178 55.3248
R1497 VTAIL.n91 VTAIL.n90 55.3248
R1498 VTAIL.n1 VTAIL.n0 55.3246
R1499 VTAIL.n89 VTAIL.n88 55.3246
R1500 VTAIL.n351 VTAIL.n350 33.9308
R1501 VTAIL.n87 VTAIL.n86 33.9308
R1502 VTAIL.n265 VTAIL.n264 33.9308
R1503 VTAIL.n177 VTAIL.n176 33.9308
R1504 VTAIL.n91 VTAIL.n89 31.1169
R1505 VTAIL.n351 VTAIL.n265 28.4014
R1506 VTAIL.n294 VTAIL.n293 16.3895
R1507 VTAIL.n30 VTAIL.n29 16.3895
R1508 VTAIL.n210 VTAIL.n209 16.3895
R1509 VTAIL.n122 VTAIL.n121 16.3895
R1510 VTAIL.n339 VTAIL.n270 13.1884
R1511 VTAIL.n75 VTAIL.n6 13.1884
R1512 VTAIL.n186 VTAIL.n184 13.1884
R1513 VTAIL.n98 VTAIL.n96 13.1884
R1514 VTAIL.n297 VTAIL.n292 12.8005
R1515 VTAIL.n340 VTAIL.n272 12.8005
R1516 VTAIL.n344 VTAIL.n343 12.8005
R1517 VTAIL.n33 VTAIL.n28 12.8005
R1518 VTAIL.n76 VTAIL.n8 12.8005
R1519 VTAIL.n80 VTAIL.n79 12.8005
R1520 VTAIL.n258 VTAIL.n257 12.8005
R1521 VTAIL.n254 VTAIL.n253 12.8005
R1522 VTAIL.n213 VTAIL.n208 12.8005
R1523 VTAIL.n170 VTAIL.n169 12.8005
R1524 VTAIL.n166 VTAIL.n165 12.8005
R1525 VTAIL.n125 VTAIL.n120 12.8005
R1526 VTAIL.n298 VTAIL.n290 12.0247
R1527 VTAIL.n335 VTAIL.n334 12.0247
R1528 VTAIL.n347 VTAIL.n268 12.0247
R1529 VTAIL.n34 VTAIL.n26 12.0247
R1530 VTAIL.n71 VTAIL.n70 12.0247
R1531 VTAIL.n83 VTAIL.n4 12.0247
R1532 VTAIL.n261 VTAIL.n182 12.0247
R1533 VTAIL.n250 VTAIL.n187 12.0247
R1534 VTAIL.n214 VTAIL.n206 12.0247
R1535 VTAIL.n173 VTAIL.n94 12.0247
R1536 VTAIL.n162 VTAIL.n99 12.0247
R1537 VTAIL.n126 VTAIL.n118 12.0247
R1538 VTAIL.n302 VTAIL.n301 11.249
R1539 VTAIL.n333 VTAIL.n274 11.249
R1540 VTAIL.n348 VTAIL.n266 11.249
R1541 VTAIL.n38 VTAIL.n37 11.249
R1542 VTAIL.n69 VTAIL.n10 11.249
R1543 VTAIL.n84 VTAIL.n2 11.249
R1544 VTAIL.n262 VTAIL.n180 11.249
R1545 VTAIL.n249 VTAIL.n190 11.249
R1546 VTAIL.n218 VTAIL.n217 11.249
R1547 VTAIL.n174 VTAIL.n92 11.249
R1548 VTAIL.n161 VTAIL.n102 11.249
R1549 VTAIL.n130 VTAIL.n129 11.249
R1550 VTAIL.n305 VTAIL.n288 10.4732
R1551 VTAIL.n330 VTAIL.n329 10.4732
R1552 VTAIL.n41 VTAIL.n24 10.4732
R1553 VTAIL.n66 VTAIL.n65 10.4732
R1554 VTAIL.n246 VTAIL.n245 10.4732
R1555 VTAIL.n221 VTAIL.n204 10.4732
R1556 VTAIL.n158 VTAIL.n157 10.4732
R1557 VTAIL.n133 VTAIL.n116 10.4732
R1558 VTAIL.n306 VTAIL.n286 9.69747
R1559 VTAIL.n326 VTAIL.n276 9.69747
R1560 VTAIL.n42 VTAIL.n22 9.69747
R1561 VTAIL.n62 VTAIL.n12 9.69747
R1562 VTAIL.n242 VTAIL.n192 9.69747
R1563 VTAIL.n222 VTAIL.n202 9.69747
R1564 VTAIL.n154 VTAIL.n104 9.69747
R1565 VTAIL.n134 VTAIL.n114 9.69747
R1566 VTAIL.n350 VTAIL.n349 9.45567
R1567 VTAIL.n86 VTAIL.n85 9.45567
R1568 VTAIL.n264 VTAIL.n263 9.45567
R1569 VTAIL.n176 VTAIL.n175 9.45567
R1570 VTAIL.n349 VTAIL.n348 9.3005
R1571 VTAIL.n268 VTAIL.n267 9.3005
R1572 VTAIL.n343 VTAIL.n342 9.3005
R1573 VTAIL.n315 VTAIL.n314 9.3005
R1574 VTAIL.n284 VTAIL.n283 9.3005
R1575 VTAIL.n309 VTAIL.n308 9.3005
R1576 VTAIL.n307 VTAIL.n306 9.3005
R1577 VTAIL.n288 VTAIL.n287 9.3005
R1578 VTAIL.n301 VTAIL.n300 9.3005
R1579 VTAIL.n299 VTAIL.n298 9.3005
R1580 VTAIL.n292 VTAIL.n291 9.3005
R1581 VTAIL.n317 VTAIL.n316 9.3005
R1582 VTAIL.n280 VTAIL.n279 9.3005
R1583 VTAIL.n323 VTAIL.n322 9.3005
R1584 VTAIL.n325 VTAIL.n324 9.3005
R1585 VTAIL.n276 VTAIL.n275 9.3005
R1586 VTAIL.n331 VTAIL.n330 9.3005
R1587 VTAIL.n333 VTAIL.n332 9.3005
R1588 VTAIL.n334 VTAIL.n271 9.3005
R1589 VTAIL.n341 VTAIL.n340 9.3005
R1590 VTAIL.n85 VTAIL.n84 9.3005
R1591 VTAIL.n4 VTAIL.n3 9.3005
R1592 VTAIL.n79 VTAIL.n78 9.3005
R1593 VTAIL.n51 VTAIL.n50 9.3005
R1594 VTAIL.n20 VTAIL.n19 9.3005
R1595 VTAIL.n45 VTAIL.n44 9.3005
R1596 VTAIL.n43 VTAIL.n42 9.3005
R1597 VTAIL.n24 VTAIL.n23 9.3005
R1598 VTAIL.n37 VTAIL.n36 9.3005
R1599 VTAIL.n35 VTAIL.n34 9.3005
R1600 VTAIL.n28 VTAIL.n27 9.3005
R1601 VTAIL.n53 VTAIL.n52 9.3005
R1602 VTAIL.n16 VTAIL.n15 9.3005
R1603 VTAIL.n59 VTAIL.n58 9.3005
R1604 VTAIL.n61 VTAIL.n60 9.3005
R1605 VTAIL.n12 VTAIL.n11 9.3005
R1606 VTAIL.n67 VTAIL.n66 9.3005
R1607 VTAIL.n69 VTAIL.n68 9.3005
R1608 VTAIL.n70 VTAIL.n7 9.3005
R1609 VTAIL.n77 VTAIL.n76 9.3005
R1610 VTAIL.n196 VTAIL.n195 9.3005
R1611 VTAIL.n239 VTAIL.n238 9.3005
R1612 VTAIL.n241 VTAIL.n240 9.3005
R1613 VTAIL.n192 VTAIL.n191 9.3005
R1614 VTAIL.n247 VTAIL.n246 9.3005
R1615 VTAIL.n249 VTAIL.n248 9.3005
R1616 VTAIL.n187 VTAIL.n185 9.3005
R1617 VTAIL.n255 VTAIL.n254 9.3005
R1618 VTAIL.n263 VTAIL.n262 9.3005
R1619 VTAIL.n182 VTAIL.n181 9.3005
R1620 VTAIL.n257 VTAIL.n256 9.3005
R1621 VTAIL.n233 VTAIL.n232 9.3005
R1622 VTAIL.n231 VTAIL.n230 9.3005
R1623 VTAIL.n200 VTAIL.n199 9.3005
R1624 VTAIL.n225 VTAIL.n224 9.3005
R1625 VTAIL.n223 VTAIL.n222 9.3005
R1626 VTAIL.n204 VTAIL.n203 9.3005
R1627 VTAIL.n217 VTAIL.n216 9.3005
R1628 VTAIL.n215 VTAIL.n214 9.3005
R1629 VTAIL.n208 VTAIL.n207 9.3005
R1630 VTAIL.n108 VTAIL.n107 9.3005
R1631 VTAIL.n151 VTAIL.n150 9.3005
R1632 VTAIL.n153 VTAIL.n152 9.3005
R1633 VTAIL.n104 VTAIL.n103 9.3005
R1634 VTAIL.n159 VTAIL.n158 9.3005
R1635 VTAIL.n161 VTAIL.n160 9.3005
R1636 VTAIL.n99 VTAIL.n97 9.3005
R1637 VTAIL.n167 VTAIL.n166 9.3005
R1638 VTAIL.n175 VTAIL.n174 9.3005
R1639 VTAIL.n94 VTAIL.n93 9.3005
R1640 VTAIL.n169 VTAIL.n168 9.3005
R1641 VTAIL.n145 VTAIL.n144 9.3005
R1642 VTAIL.n143 VTAIL.n142 9.3005
R1643 VTAIL.n112 VTAIL.n111 9.3005
R1644 VTAIL.n137 VTAIL.n136 9.3005
R1645 VTAIL.n135 VTAIL.n134 9.3005
R1646 VTAIL.n116 VTAIL.n115 9.3005
R1647 VTAIL.n129 VTAIL.n128 9.3005
R1648 VTAIL.n127 VTAIL.n126 9.3005
R1649 VTAIL.n120 VTAIL.n119 9.3005
R1650 VTAIL.n310 VTAIL.n309 8.92171
R1651 VTAIL.n325 VTAIL.n278 8.92171
R1652 VTAIL.n46 VTAIL.n45 8.92171
R1653 VTAIL.n61 VTAIL.n14 8.92171
R1654 VTAIL.n241 VTAIL.n194 8.92171
R1655 VTAIL.n226 VTAIL.n225 8.92171
R1656 VTAIL.n153 VTAIL.n106 8.92171
R1657 VTAIL.n138 VTAIL.n137 8.92171
R1658 VTAIL.n313 VTAIL.n284 8.14595
R1659 VTAIL.n322 VTAIL.n321 8.14595
R1660 VTAIL.n49 VTAIL.n20 8.14595
R1661 VTAIL.n58 VTAIL.n57 8.14595
R1662 VTAIL.n238 VTAIL.n237 8.14595
R1663 VTAIL.n229 VTAIL.n200 8.14595
R1664 VTAIL.n150 VTAIL.n149 8.14595
R1665 VTAIL.n141 VTAIL.n112 8.14595
R1666 VTAIL.n314 VTAIL.n282 7.3702
R1667 VTAIL.n318 VTAIL.n280 7.3702
R1668 VTAIL.n50 VTAIL.n18 7.3702
R1669 VTAIL.n54 VTAIL.n16 7.3702
R1670 VTAIL.n234 VTAIL.n196 7.3702
R1671 VTAIL.n230 VTAIL.n198 7.3702
R1672 VTAIL.n146 VTAIL.n108 7.3702
R1673 VTAIL.n142 VTAIL.n110 7.3702
R1674 VTAIL.n317 VTAIL.n282 6.59444
R1675 VTAIL.n318 VTAIL.n317 6.59444
R1676 VTAIL.n53 VTAIL.n18 6.59444
R1677 VTAIL.n54 VTAIL.n53 6.59444
R1678 VTAIL.n234 VTAIL.n233 6.59444
R1679 VTAIL.n233 VTAIL.n198 6.59444
R1680 VTAIL.n146 VTAIL.n145 6.59444
R1681 VTAIL.n145 VTAIL.n110 6.59444
R1682 VTAIL.n314 VTAIL.n313 5.81868
R1683 VTAIL.n321 VTAIL.n280 5.81868
R1684 VTAIL.n50 VTAIL.n49 5.81868
R1685 VTAIL.n57 VTAIL.n16 5.81868
R1686 VTAIL.n237 VTAIL.n196 5.81868
R1687 VTAIL.n230 VTAIL.n229 5.81868
R1688 VTAIL.n149 VTAIL.n108 5.81868
R1689 VTAIL.n142 VTAIL.n141 5.81868
R1690 VTAIL.n310 VTAIL.n284 5.04292
R1691 VTAIL.n322 VTAIL.n278 5.04292
R1692 VTAIL.n46 VTAIL.n20 5.04292
R1693 VTAIL.n58 VTAIL.n14 5.04292
R1694 VTAIL.n238 VTAIL.n194 5.04292
R1695 VTAIL.n226 VTAIL.n200 5.04292
R1696 VTAIL.n150 VTAIL.n106 5.04292
R1697 VTAIL.n138 VTAIL.n112 5.04292
R1698 VTAIL.n309 VTAIL.n286 4.26717
R1699 VTAIL.n326 VTAIL.n325 4.26717
R1700 VTAIL.n45 VTAIL.n22 4.26717
R1701 VTAIL.n62 VTAIL.n61 4.26717
R1702 VTAIL.n242 VTAIL.n241 4.26717
R1703 VTAIL.n225 VTAIL.n202 4.26717
R1704 VTAIL.n154 VTAIL.n153 4.26717
R1705 VTAIL.n137 VTAIL.n114 4.26717
R1706 VTAIL.n293 VTAIL.n291 3.70982
R1707 VTAIL.n29 VTAIL.n27 3.70982
R1708 VTAIL.n209 VTAIL.n207 3.70982
R1709 VTAIL.n121 VTAIL.n119 3.70982
R1710 VTAIL.n306 VTAIL.n305 3.49141
R1711 VTAIL.n329 VTAIL.n276 3.49141
R1712 VTAIL.n42 VTAIL.n41 3.49141
R1713 VTAIL.n65 VTAIL.n12 3.49141
R1714 VTAIL.n245 VTAIL.n192 3.49141
R1715 VTAIL.n222 VTAIL.n221 3.49141
R1716 VTAIL.n157 VTAIL.n104 3.49141
R1717 VTAIL.n134 VTAIL.n133 3.49141
R1718 VTAIL.n177 VTAIL.n91 2.71602
R1719 VTAIL.n265 VTAIL.n179 2.71602
R1720 VTAIL.n89 VTAIL.n87 2.71602
R1721 VTAIL.n302 VTAIL.n288 2.71565
R1722 VTAIL.n330 VTAIL.n274 2.71565
R1723 VTAIL.n350 VTAIL.n266 2.71565
R1724 VTAIL.n38 VTAIL.n24 2.71565
R1725 VTAIL.n66 VTAIL.n10 2.71565
R1726 VTAIL.n86 VTAIL.n2 2.71565
R1727 VTAIL.n264 VTAIL.n180 2.71565
R1728 VTAIL.n246 VTAIL.n190 2.71565
R1729 VTAIL.n218 VTAIL.n204 2.71565
R1730 VTAIL.n176 VTAIL.n92 2.71565
R1731 VTAIL.n158 VTAIL.n102 2.71565
R1732 VTAIL.n130 VTAIL.n116 2.71565
R1733 VTAIL.n0 VTAIL.t5 2.10438
R1734 VTAIL.n0 VTAIL.t3 2.10438
R1735 VTAIL.n88 VTAIL.t6 2.10438
R1736 VTAIL.n88 VTAIL.t7 2.10438
R1737 VTAIL.n178 VTAIL.t8 2.10438
R1738 VTAIL.n178 VTAIL.t11 2.10438
R1739 VTAIL.n90 VTAIL.t0 2.10438
R1740 VTAIL.n90 VTAIL.t4 2.10438
R1741 VTAIL VTAIL.n351 1.97895
R1742 VTAIL.n301 VTAIL.n290 1.93989
R1743 VTAIL.n335 VTAIL.n333 1.93989
R1744 VTAIL.n348 VTAIL.n347 1.93989
R1745 VTAIL.n37 VTAIL.n26 1.93989
R1746 VTAIL.n71 VTAIL.n69 1.93989
R1747 VTAIL.n84 VTAIL.n83 1.93989
R1748 VTAIL.n262 VTAIL.n261 1.93989
R1749 VTAIL.n250 VTAIL.n249 1.93989
R1750 VTAIL.n217 VTAIL.n206 1.93989
R1751 VTAIL.n174 VTAIL.n173 1.93989
R1752 VTAIL.n162 VTAIL.n161 1.93989
R1753 VTAIL.n129 VTAIL.n118 1.93989
R1754 VTAIL.n179 VTAIL.n177 1.82809
R1755 VTAIL.n87 VTAIL.n1 1.82809
R1756 VTAIL.n298 VTAIL.n297 1.16414
R1757 VTAIL.n334 VTAIL.n272 1.16414
R1758 VTAIL.n344 VTAIL.n268 1.16414
R1759 VTAIL.n34 VTAIL.n33 1.16414
R1760 VTAIL.n70 VTAIL.n8 1.16414
R1761 VTAIL.n80 VTAIL.n4 1.16414
R1762 VTAIL.n258 VTAIL.n182 1.16414
R1763 VTAIL.n253 VTAIL.n187 1.16414
R1764 VTAIL.n214 VTAIL.n213 1.16414
R1765 VTAIL.n170 VTAIL.n94 1.16414
R1766 VTAIL.n165 VTAIL.n99 1.16414
R1767 VTAIL.n126 VTAIL.n125 1.16414
R1768 VTAIL VTAIL.n1 0.737569
R1769 VTAIL.n294 VTAIL.n292 0.388379
R1770 VTAIL.n340 VTAIL.n339 0.388379
R1771 VTAIL.n343 VTAIL.n270 0.388379
R1772 VTAIL.n30 VTAIL.n28 0.388379
R1773 VTAIL.n76 VTAIL.n75 0.388379
R1774 VTAIL.n79 VTAIL.n6 0.388379
R1775 VTAIL.n257 VTAIL.n184 0.388379
R1776 VTAIL.n254 VTAIL.n186 0.388379
R1777 VTAIL.n210 VTAIL.n208 0.388379
R1778 VTAIL.n169 VTAIL.n96 0.388379
R1779 VTAIL.n166 VTAIL.n98 0.388379
R1780 VTAIL.n122 VTAIL.n120 0.388379
R1781 VTAIL.n299 VTAIL.n291 0.155672
R1782 VTAIL.n300 VTAIL.n299 0.155672
R1783 VTAIL.n300 VTAIL.n287 0.155672
R1784 VTAIL.n307 VTAIL.n287 0.155672
R1785 VTAIL.n308 VTAIL.n307 0.155672
R1786 VTAIL.n308 VTAIL.n283 0.155672
R1787 VTAIL.n315 VTAIL.n283 0.155672
R1788 VTAIL.n316 VTAIL.n315 0.155672
R1789 VTAIL.n316 VTAIL.n279 0.155672
R1790 VTAIL.n323 VTAIL.n279 0.155672
R1791 VTAIL.n324 VTAIL.n323 0.155672
R1792 VTAIL.n324 VTAIL.n275 0.155672
R1793 VTAIL.n331 VTAIL.n275 0.155672
R1794 VTAIL.n332 VTAIL.n331 0.155672
R1795 VTAIL.n332 VTAIL.n271 0.155672
R1796 VTAIL.n341 VTAIL.n271 0.155672
R1797 VTAIL.n342 VTAIL.n341 0.155672
R1798 VTAIL.n342 VTAIL.n267 0.155672
R1799 VTAIL.n349 VTAIL.n267 0.155672
R1800 VTAIL.n35 VTAIL.n27 0.155672
R1801 VTAIL.n36 VTAIL.n35 0.155672
R1802 VTAIL.n36 VTAIL.n23 0.155672
R1803 VTAIL.n43 VTAIL.n23 0.155672
R1804 VTAIL.n44 VTAIL.n43 0.155672
R1805 VTAIL.n44 VTAIL.n19 0.155672
R1806 VTAIL.n51 VTAIL.n19 0.155672
R1807 VTAIL.n52 VTAIL.n51 0.155672
R1808 VTAIL.n52 VTAIL.n15 0.155672
R1809 VTAIL.n59 VTAIL.n15 0.155672
R1810 VTAIL.n60 VTAIL.n59 0.155672
R1811 VTAIL.n60 VTAIL.n11 0.155672
R1812 VTAIL.n67 VTAIL.n11 0.155672
R1813 VTAIL.n68 VTAIL.n67 0.155672
R1814 VTAIL.n68 VTAIL.n7 0.155672
R1815 VTAIL.n77 VTAIL.n7 0.155672
R1816 VTAIL.n78 VTAIL.n77 0.155672
R1817 VTAIL.n78 VTAIL.n3 0.155672
R1818 VTAIL.n85 VTAIL.n3 0.155672
R1819 VTAIL.n263 VTAIL.n181 0.155672
R1820 VTAIL.n256 VTAIL.n181 0.155672
R1821 VTAIL.n256 VTAIL.n255 0.155672
R1822 VTAIL.n255 VTAIL.n185 0.155672
R1823 VTAIL.n248 VTAIL.n185 0.155672
R1824 VTAIL.n248 VTAIL.n247 0.155672
R1825 VTAIL.n247 VTAIL.n191 0.155672
R1826 VTAIL.n240 VTAIL.n191 0.155672
R1827 VTAIL.n240 VTAIL.n239 0.155672
R1828 VTAIL.n239 VTAIL.n195 0.155672
R1829 VTAIL.n232 VTAIL.n195 0.155672
R1830 VTAIL.n232 VTAIL.n231 0.155672
R1831 VTAIL.n231 VTAIL.n199 0.155672
R1832 VTAIL.n224 VTAIL.n199 0.155672
R1833 VTAIL.n224 VTAIL.n223 0.155672
R1834 VTAIL.n223 VTAIL.n203 0.155672
R1835 VTAIL.n216 VTAIL.n203 0.155672
R1836 VTAIL.n216 VTAIL.n215 0.155672
R1837 VTAIL.n215 VTAIL.n207 0.155672
R1838 VTAIL.n175 VTAIL.n93 0.155672
R1839 VTAIL.n168 VTAIL.n93 0.155672
R1840 VTAIL.n168 VTAIL.n167 0.155672
R1841 VTAIL.n167 VTAIL.n97 0.155672
R1842 VTAIL.n160 VTAIL.n97 0.155672
R1843 VTAIL.n160 VTAIL.n159 0.155672
R1844 VTAIL.n159 VTAIL.n103 0.155672
R1845 VTAIL.n152 VTAIL.n103 0.155672
R1846 VTAIL.n152 VTAIL.n151 0.155672
R1847 VTAIL.n151 VTAIL.n107 0.155672
R1848 VTAIL.n144 VTAIL.n107 0.155672
R1849 VTAIL.n144 VTAIL.n143 0.155672
R1850 VTAIL.n143 VTAIL.n111 0.155672
R1851 VTAIL.n136 VTAIL.n111 0.155672
R1852 VTAIL.n136 VTAIL.n135 0.155672
R1853 VTAIL.n135 VTAIL.n115 0.155672
R1854 VTAIL.n128 VTAIL.n115 0.155672
R1855 VTAIL.n128 VTAIL.n127 0.155672
R1856 VTAIL.n127 VTAIL.n119 0.155672
R1857 VDD1.n80 VDD1.n0 756.745
R1858 VDD1.n165 VDD1.n85 756.745
R1859 VDD1.n81 VDD1.n80 585
R1860 VDD1.n79 VDD1.n78 585
R1861 VDD1.n4 VDD1.n3 585
R1862 VDD1.n8 VDD1.n6 585
R1863 VDD1.n73 VDD1.n72 585
R1864 VDD1.n71 VDD1.n70 585
R1865 VDD1.n10 VDD1.n9 585
R1866 VDD1.n65 VDD1.n64 585
R1867 VDD1.n63 VDD1.n62 585
R1868 VDD1.n14 VDD1.n13 585
R1869 VDD1.n57 VDD1.n56 585
R1870 VDD1.n55 VDD1.n54 585
R1871 VDD1.n18 VDD1.n17 585
R1872 VDD1.n49 VDD1.n48 585
R1873 VDD1.n47 VDD1.n46 585
R1874 VDD1.n22 VDD1.n21 585
R1875 VDD1.n41 VDD1.n40 585
R1876 VDD1.n39 VDD1.n38 585
R1877 VDD1.n26 VDD1.n25 585
R1878 VDD1.n33 VDD1.n32 585
R1879 VDD1.n31 VDD1.n30 585
R1880 VDD1.n114 VDD1.n113 585
R1881 VDD1.n116 VDD1.n115 585
R1882 VDD1.n109 VDD1.n108 585
R1883 VDD1.n122 VDD1.n121 585
R1884 VDD1.n124 VDD1.n123 585
R1885 VDD1.n105 VDD1.n104 585
R1886 VDD1.n130 VDD1.n129 585
R1887 VDD1.n132 VDD1.n131 585
R1888 VDD1.n101 VDD1.n100 585
R1889 VDD1.n138 VDD1.n137 585
R1890 VDD1.n140 VDD1.n139 585
R1891 VDD1.n97 VDD1.n96 585
R1892 VDD1.n146 VDD1.n145 585
R1893 VDD1.n148 VDD1.n147 585
R1894 VDD1.n93 VDD1.n92 585
R1895 VDD1.n155 VDD1.n154 585
R1896 VDD1.n156 VDD1.n91 585
R1897 VDD1.n158 VDD1.n157 585
R1898 VDD1.n89 VDD1.n88 585
R1899 VDD1.n164 VDD1.n163 585
R1900 VDD1.n166 VDD1.n165 585
R1901 VDD1.n29 VDD1.t4 327.466
R1902 VDD1.n112 VDD1.t3 327.466
R1903 VDD1.n80 VDD1.n79 171.744
R1904 VDD1.n79 VDD1.n3 171.744
R1905 VDD1.n8 VDD1.n3 171.744
R1906 VDD1.n72 VDD1.n8 171.744
R1907 VDD1.n72 VDD1.n71 171.744
R1908 VDD1.n71 VDD1.n9 171.744
R1909 VDD1.n64 VDD1.n9 171.744
R1910 VDD1.n64 VDD1.n63 171.744
R1911 VDD1.n63 VDD1.n13 171.744
R1912 VDD1.n56 VDD1.n13 171.744
R1913 VDD1.n56 VDD1.n55 171.744
R1914 VDD1.n55 VDD1.n17 171.744
R1915 VDD1.n48 VDD1.n17 171.744
R1916 VDD1.n48 VDD1.n47 171.744
R1917 VDD1.n47 VDD1.n21 171.744
R1918 VDD1.n40 VDD1.n21 171.744
R1919 VDD1.n40 VDD1.n39 171.744
R1920 VDD1.n39 VDD1.n25 171.744
R1921 VDD1.n32 VDD1.n25 171.744
R1922 VDD1.n32 VDD1.n31 171.744
R1923 VDD1.n115 VDD1.n114 171.744
R1924 VDD1.n115 VDD1.n108 171.744
R1925 VDD1.n122 VDD1.n108 171.744
R1926 VDD1.n123 VDD1.n122 171.744
R1927 VDD1.n123 VDD1.n104 171.744
R1928 VDD1.n130 VDD1.n104 171.744
R1929 VDD1.n131 VDD1.n130 171.744
R1930 VDD1.n131 VDD1.n100 171.744
R1931 VDD1.n138 VDD1.n100 171.744
R1932 VDD1.n139 VDD1.n138 171.744
R1933 VDD1.n139 VDD1.n96 171.744
R1934 VDD1.n146 VDD1.n96 171.744
R1935 VDD1.n147 VDD1.n146 171.744
R1936 VDD1.n147 VDD1.n92 171.744
R1937 VDD1.n155 VDD1.n92 171.744
R1938 VDD1.n156 VDD1.n155 171.744
R1939 VDD1.n157 VDD1.n156 171.744
R1940 VDD1.n157 VDD1.n88 171.744
R1941 VDD1.n164 VDD1.n88 171.744
R1942 VDD1.n165 VDD1.n164 171.744
R1943 VDD1.n31 VDD1.t4 85.8723
R1944 VDD1.n114 VDD1.t3 85.8723
R1945 VDD1.n171 VDD1.n170 72.6269
R1946 VDD1.n173 VDD1.n172 72.0034
R1947 VDD1 VDD1.n84 52.7044
R1948 VDD1.n171 VDD1.n169 52.5909
R1949 VDD1.n173 VDD1.n171 47.8005
R1950 VDD1.n30 VDD1.n29 16.3895
R1951 VDD1.n113 VDD1.n112 16.3895
R1952 VDD1.n6 VDD1.n4 13.1884
R1953 VDD1.n158 VDD1.n89 13.1884
R1954 VDD1.n78 VDD1.n77 12.8005
R1955 VDD1.n74 VDD1.n73 12.8005
R1956 VDD1.n33 VDD1.n28 12.8005
R1957 VDD1.n116 VDD1.n111 12.8005
R1958 VDD1.n159 VDD1.n91 12.8005
R1959 VDD1.n163 VDD1.n162 12.8005
R1960 VDD1.n81 VDD1.n2 12.0247
R1961 VDD1.n70 VDD1.n7 12.0247
R1962 VDD1.n34 VDD1.n26 12.0247
R1963 VDD1.n117 VDD1.n109 12.0247
R1964 VDD1.n154 VDD1.n153 12.0247
R1965 VDD1.n166 VDD1.n87 12.0247
R1966 VDD1.n82 VDD1.n0 11.249
R1967 VDD1.n69 VDD1.n10 11.249
R1968 VDD1.n38 VDD1.n37 11.249
R1969 VDD1.n121 VDD1.n120 11.249
R1970 VDD1.n152 VDD1.n93 11.249
R1971 VDD1.n167 VDD1.n85 11.249
R1972 VDD1.n66 VDD1.n65 10.4732
R1973 VDD1.n41 VDD1.n24 10.4732
R1974 VDD1.n124 VDD1.n107 10.4732
R1975 VDD1.n149 VDD1.n148 10.4732
R1976 VDD1.n62 VDD1.n12 9.69747
R1977 VDD1.n42 VDD1.n22 9.69747
R1978 VDD1.n125 VDD1.n105 9.69747
R1979 VDD1.n145 VDD1.n95 9.69747
R1980 VDD1.n84 VDD1.n83 9.45567
R1981 VDD1.n169 VDD1.n168 9.45567
R1982 VDD1.n16 VDD1.n15 9.3005
R1983 VDD1.n59 VDD1.n58 9.3005
R1984 VDD1.n61 VDD1.n60 9.3005
R1985 VDD1.n12 VDD1.n11 9.3005
R1986 VDD1.n67 VDD1.n66 9.3005
R1987 VDD1.n69 VDD1.n68 9.3005
R1988 VDD1.n7 VDD1.n5 9.3005
R1989 VDD1.n75 VDD1.n74 9.3005
R1990 VDD1.n83 VDD1.n82 9.3005
R1991 VDD1.n2 VDD1.n1 9.3005
R1992 VDD1.n77 VDD1.n76 9.3005
R1993 VDD1.n53 VDD1.n52 9.3005
R1994 VDD1.n51 VDD1.n50 9.3005
R1995 VDD1.n20 VDD1.n19 9.3005
R1996 VDD1.n45 VDD1.n44 9.3005
R1997 VDD1.n43 VDD1.n42 9.3005
R1998 VDD1.n24 VDD1.n23 9.3005
R1999 VDD1.n37 VDD1.n36 9.3005
R2000 VDD1.n35 VDD1.n34 9.3005
R2001 VDD1.n28 VDD1.n27 9.3005
R2002 VDD1.n168 VDD1.n167 9.3005
R2003 VDD1.n87 VDD1.n86 9.3005
R2004 VDD1.n162 VDD1.n161 9.3005
R2005 VDD1.n134 VDD1.n133 9.3005
R2006 VDD1.n103 VDD1.n102 9.3005
R2007 VDD1.n128 VDD1.n127 9.3005
R2008 VDD1.n126 VDD1.n125 9.3005
R2009 VDD1.n107 VDD1.n106 9.3005
R2010 VDD1.n120 VDD1.n119 9.3005
R2011 VDD1.n118 VDD1.n117 9.3005
R2012 VDD1.n111 VDD1.n110 9.3005
R2013 VDD1.n136 VDD1.n135 9.3005
R2014 VDD1.n99 VDD1.n98 9.3005
R2015 VDD1.n142 VDD1.n141 9.3005
R2016 VDD1.n144 VDD1.n143 9.3005
R2017 VDD1.n95 VDD1.n94 9.3005
R2018 VDD1.n150 VDD1.n149 9.3005
R2019 VDD1.n152 VDD1.n151 9.3005
R2020 VDD1.n153 VDD1.n90 9.3005
R2021 VDD1.n160 VDD1.n159 9.3005
R2022 VDD1.n61 VDD1.n14 8.92171
R2023 VDD1.n46 VDD1.n45 8.92171
R2024 VDD1.n129 VDD1.n128 8.92171
R2025 VDD1.n144 VDD1.n97 8.92171
R2026 VDD1.n58 VDD1.n57 8.14595
R2027 VDD1.n49 VDD1.n20 8.14595
R2028 VDD1.n132 VDD1.n103 8.14595
R2029 VDD1.n141 VDD1.n140 8.14595
R2030 VDD1.n54 VDD1.n16 7.3702
R2031 VDD1.n50 VDD1.n18 7.3702
R2032 VDD1.n133 VDD1.n101 7.3702
R2033 VDD1.n137 VDD1.n99 7.3702
R2034 VDD1.n54 VDD1.n53 6.59444
R2035 VDD1.n53 VDD1.n18 6.59444
R2036 VDD1.n136 VDD1.n101 6.59444
R2037 VDD1.n137 VDD1.n136 6.59444
R2038 VDD1.n57 VDD1.n16 5.81868
R2039 VDD1.n50 VDD1.n49 5.81868
R2040 VDD1.n133 VDD1.n132 5.81868
R2041 VDD1.n140 VDD1.n99 5.81868
R2042 VDD1.n58 VDD1.n14 5.04292
R2043 VDD1.n46 VDD1.n20 5.04292
R2044 VDD1.n129 VDD1.n103 5.04292
R2045 VDD1.n141 VDD1.n97 5.04292
R2046 VDD1.n62 VDD1.n61 4.26717
R2047 VDD1.n45 VDD1.n22 4.26717
R2048 VDD1.n128 VDD1.n105 4.26717
R2049 VDD1.n145 VDD1.n144 4.26717
R2050 VDD1.n29 VDD1.n27 3.70982
R2051 VDD1.n112 VDD1.n110 3.70982
R2052 VDD1.n65 VDD1.n12 3.49141
R2053 VDD1.n42 VDD1.n41 3.49141
R2054 VDD1.n125 VDD1.n124 3.49141
R2055 VDD1.n148 VDD1.n95 3.49141
R2056 VDD1.n84 VDD1.n0 2.71565
R2057 VDD1.n66 VDD1.n10 2.71565
R2058 VDD1.n38 VDD1.n24 2.71565
R2059 VDD1.n121 VDD1.n107 2.71565
R2060 VDD1.n149 VDD1.n93 2.71565
R2061 VDD1.n169 VDD1.n85 2.71565
R2062 VDD1.n172 VDD1.t1 2.10438
R2063 VDD1.n172 VDD1.t5 2.10438
R2064 VDD1.n170 VDD1.t2 2.10438
R2065 VDD1.n170 VDD1.t0 2.10438
R2066 VDD1.n82 VDD1.n81 1.93989
R2067 VDD1.n70 VDD1.n69 1.93989
R2068 VDD1.n37 VDD1.n26 1.93989
R2069 VDD1.n120 VDD1.n109 1.93989
R2070 VDD1.n154 VDD1.n152 1.93989
R2071 VDD1.n167 VDD1.n166 1.93989
R2072 VDD1.n78 VDD1.n2 1.16414
R2073 VDD1.n73 VDD1.n7 1.16414
R2074 VDD1.n34 VDD1.n33 1.16414
R2075 VDD1.n117 VDD1.n116 1.16414
R2076 VDD1.n153 VDD1.n91 1.16414
R2077 VDD1.n163 VDD1.n87 1.16414
R2078 VDD1 VDD1.n173 0.62119
R2079 VDD1.n77 VDD1.n4 0.388379
R2080 VDD1.n74 VDD1.n6 0.388379
R2081 VDD1.n30 VDD1.n28 0.388379
R2082 VDD1.n113 VDD1.n111 0.388379
R2083 VDD1.n159 VDD1.n158 0.388379
R2084 VDD1.n162 VDD1.n89 0.388379
R2085 VDD1.n83 VDD1.n1 0.155672
R2086 VDD1.n76 VDD1.n1 0.155672
R2087 VDD1.n76 VDD1.n75 0.155672
R2088 VDD1.n75 VDD1.n5 0.155672
R2089 VDD1.n68 VDD1.n5 0.155672
R2090 VDD1.n68 VDD1.n67 0.155672
R2091 VDD1.n67 VDD1.n11 0.155672
R2092 VDD1.n60 VDD1.n11 0.155672
R2093 VDD1.n60 VDD1.n59 0.155672
R2094 VDD1.n59 VDD1.n15 0.155672
R2095 VDD1.n52 VDD1.n15 0.155672
R2096 VDD1.n52 VDD1.n51 0.155672
R2097 VDD1.n51 VDD1.n19 0.155672
R2098 VDD1.n44 VDD1.n19 0.155672
R2099 VDD1.n44 VDD1.n43 0.155672
R2100 VDD1.n43 VDD1.n23 0.155672
R2101 VDD1.n36 VDD1.n23 0.155672
R2102 VDD1.n36 VDD1.n35 0.155672
R2103 VDD1.n35 VDD1.n27 0.155672
R2104 VDD1.n118 VDD1.n110 0.155672
R2105 VDD1.n119 VDD1.n118 0.155672
R2106 VDD1.n119 VDD1.n106 0.155672
R2107 VDD1.n126 VDD1.n106 0.155672
R2108 VDD1.n127 VDD1.n126 0.155672
R2109 VDD1.n127 VDD1.n102 0.155672
R2110 VDD1.n134 VDD1.n102 0.155672
R2111 VDD1.n135 VDD1.n134 0.155672
R2112 VDD1.n135 VDD1.n98 0.155672
R2113 VDD1.n142 VDD1.n98 0.155672
R2114 VDD1.n143 VDD1.n142 0.155672
R2115 VDD1.n143 VDD1.n94 0.155672
R2116 VDD1.n150 VDD1.n94 0.155672
R2117 VDD1.n151 VDD1.n150 0.155672
R2118 VDD1.n151 VDD1.n90 0.155672
R2119 VDD1.n160 VDD1.n90 0.155672
R2120 VDD1.n161 VDD1.n160 0.155672
R2121 VDD1.n161 VDD1.n86 0.155672
R2122 VDD1.n168 VDD1.n86 0.155672
R2123 VN.n4 VN.t1 163.718
R2124 VN.n20 VN.t2 163.718
R2125 VN.n30 VN.n29 161.3
R2126 VN.n28 VN.n17 161.3
R2127 VN.n27 VN.n26 161.3
R2128 VN.n25 VN.n18 161.3
R2129 VN.n24 VN.n23 161.3
R2130 VN.n22 VN.n19 161.3
R2131 VN.n14 VN.n13 161.3
R2132 VN.n12 VN.n1 161.3
R2133 VN.n11 VN.n10 161.3
R2134 VN.n9 VN.n2 161.3
R2135 VN.n8 VN.n7 161.3
R2136 VN.n6 VN.n3 161.3
R2137 VN.n5 VN.t0 132.037
R2138 VN.n0 VN.t4 132.037
R2139 VN.n21 VN.t5 132.037
R2140 VN.n16 VN.t3 132.037
R2141 VN.n15 VN.n0 70.4938
R2142 VN.n31 VN.n16 70.4938
R2143 VN.n5 VN.n4 61.3921
R2144 VN.n21 VN.n20 61.3921
R2145 VN.n11 VN.n2 56.5193
R2146 VN.n27 VN.n18 56.5193
R2147 VN VN.n31 52.3882
R2148 VN.n7 VN.n6 24.4675
R2149 VN.n7 VN.n2 24.4675
R2150 VN.n12 VN.n11 24.4675
R2151 VN.n13 VN.n12 24.4675
R2152 VN.n23 VN.n18 24.4675
R2153 VN.n23 VN.n22 24.4675
R2154 VN.n29 VN.n28 24.4675
R2155 VN.n28 VN.n27 24.4675
R2156 VN.n13 VN.n0 19.5741
R2157 VN.n29 VN.n16 19.5741
R2158 VN.n6 VN.n5 12.234
R2159 VN.n22 VN.n21 12.234
R2160 VN.n20 VN.n19 5.5843
R2161 VN.n4 VN.n3 5.5843
R2162 VN.n31 VN.n30 0.354971
R2163 VN.n15 VN.n14 0.354971
R2164 VN VN.n15 0.26696
R2165 VN.n30 VN.n17 0.189894
R2166 VN.n26 VN.n17 0.189894
R2167 VN.n26 VN.n25 0.189894
R2168 VN.n25 VN.n24 0.189894
R2169 VN.n24 VN.n19 0.189894
R2170 VN.n8 VN.n3 0.189894
R2171 VN.n9 VN.n8 0.189894
R2172 VN.n10 VN.n9 0.189894
R2173 VN.n10 VN.n1 0.189894
R2174 VN.n14 VN.n1 0.189894
R2175 VDD2.n167 VDD2.n87 756.745
R2176 VDD2.n80 VDD2.n0 756.745
R2177 VDD2.n168 VDD2.n167 585
R2178 VDD2.n166 VDD2.n165 585
R2179 VDD2.n91 VDD2.n90 585
R2180 VDD2.n95 VDD2.n93 585
R2181 VDD2.n160 VDD2.n159 585
R2182 VDD2.n158 VDD2.n157 585
R2183 VDD2.n97 VDD2.n96 585
R2184 VDD2.n152 VDD2.n151 585
R2185 VDD2.n150 VDD2.n149 585
R2186 VDD2.n101 VDD2.n100 585
R2187 VDD2.n144 VDD2.n143 585
R2188 VDD2.n142 VDD2.n141 585
R2189 VDD2.n105 VDD2.n104 585
R2190 VDD2.n136 VDD2.n135 585
R2191 VDD2.n134 VDD2.n133 585
R2192 VDD2.n109 VDD2.n108 585
R2193 VDD2.n128 VDD2.n127 585
R2194 VDD2.n126 VDD2.n125 585
R2195 VDD2.n113 VDD2.n112 585
R2196 VDD2.n120 VDD2.n119 585
R2197 VDD2.n118 VDD2.n117 585
R2198 VDD2.n29 VDD2.n28 585
R2199 VDD2.n31 VDD2.n30 585
R2200 VDD2.n24 VDD2.n23 585
R2201 VDD2.n37 VDD2.n36 585
R2202 VDD2.n39 VDD2.n38 585
R2203 VDD2.n20 VDD2.n19 585
R2204 VDD2.n45 VDD2.n44 585
R2205 VDD2.n47 VDD2.n46 585
R2206 VDD2.n16 VDD2.n15 585
R2207 VDD2.n53 VDD2.n52 585
R2208 VDD2.n55 VDD2.n54 585
R2209 VDD2.n12 VDD2.n11 585
R2210 VDD2.n61 VDD2.n60 585
R2211 VDD2.n63 VDD2.n62 585
R2212 VDD2.n8 VDD2.n7 585
R2213 VDD2.n70 VDD2.n69 585
R2214 VDD2.n71 VDD2.n6 585
R2215 VDD2.n73 VDD2.n72 585
R2216 VDD2.n4 VDD2.n3 585
R2217 VDD2.n79 VDD2.n78 585
R2218 VDD2.n81 VDD2.n80 585
R2219 VDD2.n116 VDD2.t2 327.466
R2220 VDD2.n27 VDD2.t4 327.466
R2221 VDD2.n167 VDD2.n166 171.744
R2222 VDD2.n166 VDD2.n90 171.744
R2223 VDD2.n95 VDD2.n90 171.744
R2224 VDD2.n159 VDD2.n95 171.744
R2225 VDD2.n159 VDD2.n158 171.744
R2226 VDD2.n158 VDD2.n96 171.744
R2227 VDD2.n151 VDD2.n96 171.744
R2228 VDD2.n151 VDD2.n150 171.744
R2229 VDD2.n150 VDD2.n100 171.744
R2230 VDD2.n143 VDD2.n100 171.744
R2231 VDD2.n143 VDD2.n142 171.744
R2232 VDD2.n142 VDD2.n104 171.744
R2233 VDD2.n135 VDD2.n104 171.744
R2234 VDD2.n135 VDD2.n134 171.744
R2235 VDD2.n134 VDD2.n108 171.744
R2236 VDD2.n127 VDD2.n108 171.744
R2237 VDD2.n127 VDD2.n126 171.744
R2238 VDD2.n126 VDD2.n112 171.744
R2239 VDD2.n119 VDD2.n112 171.744
R2240 VDD2.n119 VDD2.n118 171.744
R2241 VDD2.n30 VDD2.n29 171.744
R2242 VDD2.n30 VDD2.n23 171.744
R2243 VDD2.n37 VDD2.n23 171.744
R2244 VDD2.n38 VDD2.n37 171.744
R2245 VDD2.n38 VDD2.n19 171.744
R2246 VDD2.n45 VDD2.n19 171.744
R2247 VDD2.n46 VDD2.n45 171.744
R2248 VDD2.n46 VDD2.n15 171.744
R2249 VDD2.n53 VDD2.n15 171.744
R2250 VDD2.n54 VDD2.n53 171.744
R2251 VDD2.n54 VDD2.n11 171.744
R2252 VDD2.n61 VDD2.n11 171.744
R2253 VDD2.n62 VDD2.n61 171.744
R2254 VDD2.n62 VDD2.n7 171.744
R2255 VDD2.n70 VDD2.n7 171.744
R2256 VDD2.n71 VDD2.n70 171.744
R2257 VDD2.n72 VDD2.n71 171.744
R2258 VDD2.n72 VDD2.n3 171.744
R2259 VDD2.n79 VDD2.n3 171.744
R2260 VDD2.n80 VDD2.n79 171.744
R2261 VDD2.n118 VDD2.t2 85.8723
R2262 VDD2.n29 VDD2.t4 85.8723
R2263 VDD2.n86 VDD2.n85 72.6269
R2264 VDD2 VDD2.n173 72.6241
R2265 VDD2.n86 VDD2.n84 52.5909
R2266 VDD2.n172 VDD2.n171 50.6096
R2267 VDD2.n172 VDD2.n86 45.8597
R2268 VDD2.n117 VDD2.n116 16.3895
R2269 VDD2.n28 VDD2.n27 16.3895
R2270 VDD2.n93 VDD2.n91 13.1884
R2271 VDD2.n73 VDD2.n4 13.1884
R2272 VDD2.n165 VDD2.n164 12.8005
R2273 VDD2.n161 VDD2.n160 12.8005
R2274 VDD2.n120 VDD2.n115 12.8005
R2275 VDD2.n31 VDD2.n26 12.8005
R2276 VDD2.n74 VDD2.n6 12.8005
R2277 VDD2.n78 VDD2.n77 12.8005
R2278 VDD2.n168 VDD2.n89 12.0247
R2279 VDD2.n157 VDD2.n94 12.0247
R2280 VDD2.n121 VDD2.n113 12.0247
R2281 VDD2.n32 VDD2.n24 12.0247
R2282 VDD2.n69 VDD2.n68 12.0247
R2283 VDD2.n81 VDD2.n2 12.0247
R2284 VDD2.n169 VDD2.n87 11.249
R2285 VDD2.n156 VDD2.n97 11.249
R2286 VDD2.n125 VDD2.n124 11.249
R2287 VDD2.n36 VDD2.n35 11.249
R2288 VDD2.n67 VDD2.n8 11.249
R2289 VDD2.n82 VDD2.n0 11.249
R2290 VDD2.n153 VDD2.n152 10.4732
R2291 VDD2.n128 VDD2.n111 10.4732
R2292 VDD2.n39 VDD2.n22 10.4732
R2293 VDD2.n64 VDD2.n63 10.4732
R2294 VDD2.n149 VDD2.n99 9.69747
R2295 VDD2.n129 VDD2.n109 9.69747
R2296 VDD2.n40 VDD2.n20 9.69747
R2297 VDD2.n60 VDD2.n10 9.69747
R2298 VDD2.n171 VDD2.n170 9.45567
R2299 VDD2.n84 VDD2.n83 9.45567
R2300 VDD2.n103 VDD2.n102 9.3005
R2301 VDD2.n146 VDD2.n145 9.3005
R2302 VDD2.n148 VDD2.n147 9.3005
R2303 VDD2.n99 VDD2.n98 9.3005
R2304 VDD2.n154 VDD2.n153 9.3005
R2305 VDD2.n156 VDD2.n155 9.3005
R2306 VDD2.n94 VDD2.n92 9.3005
R2307 VDD2.n162 VDD2.n161 9.3005
R2308 VDD2.n170 VDD2.n169 9.3005
R2309 VDD2.n89 VDD2.n88 9.3005
R2310 VDD2.n164 VDD2.n163 9.3005
R2311 VDD2.n140 VDD2.n139 9.3005
R2312 VDD2.n138 VDD2.n137 9.3005
R2313 VDD2.n107 VDD2.n106 9.3005
R2314 VDD2.n132 VDD2.n131 9.3005
R2315 VDD2.n130 VDD2.n129 9.3005
R2316 VDD2.n111 VDD2.n110 9.3005
R2317 VDD2.n124 VDD2.n123 9.3005
R2318 VDD2.n122 VDD2.n121 9.3005
R2319 VDD2.n115 VDD2.n114 9.3005
R2320 VDD2.n83 VDD2.n82 9.3005
R2321 VDD2.n2 VDD2.n1 9.3005
R2322 VDD2.n77 VDD2.n76 9.3005
R2323 VDD2.n49 VDD2.n48 9.3005
R2324 VDD2.n18 VDD2.n17 9.3005
R2325 VDD2.n43 VDD2.n42 9.3005
R2326 VDD2.n41 VDD2.n40 9.3005
R2327 VDD2.n22 VDD2.n21 9.3005
R2328 VDD2.n35 VDD2.n34 9.3005
R2329 VDD2.n33 VDD2.n32 9.3005
R2330 VDD2.n26 VDD2.n25 9.3005
R2331 VDD2.n51 VDD2.n50 9.3005
R2332 VDD2.n14 VDD2.n13 9.3005
R2333 VDD2.n57 VDD2.n56 9.3005
R2334 VDD2.n59 VDD2.n58 9.3005
R2335 VDD2.n10 VDD2.n9 9.3005
R2336 VDD2.n65 VDD2.n64 9.3005
R2337 VDD2.n67 VDD2.n66 9.3005
R2338 VDD2.n68 VDD2.n5 9.3005
R2339 VDD2.n75 VDD2.n74 9.3005
R2340 VDD2.n148 VDD2.n101 8.92171
R2341 VDD2.n133 VDD2.n132 8.92171
R2342 VDD2.n44 VDD2.n43 8.92171
R2343 VDD2.n59 VDD2.n12 8.92171
R2344 VDD2.n145 VDD2.n144 8.14595
R2345 VDD2.n136 VDD2.n107 8.14595
R2346 VDD2.n47 VDD2.n18 8.14595
R2347 VDD2.n56 VDD2.n55 8.14595
R2348 VDD2.n141 VDD2.n103 7.3702
R2349 VDD2.n137 VDD2.n105 7.3702
R2350 VDD2.n48 VDD2.n16 7.3702
R2351 VDD2.n52 VDD2.n14 7.3702
R2352 VDD2.n141 VDD2.n140 6.59444
R2353 VDD2.n140 VDD2.n105 6.59444
R2354 VDD2.n51 VDD2.n16 6.59444
R2355 VDD2.n52 VDD2.n51 6.59444
R2356 VDD2.n144 VDD2.n103 5.81868
R2357 VDD2.n137 VDD2.n136 5.81868
R2358 VDD2.n48 VDD2.n47 5.81868
R2359 VDD2.n55 VDD2.n14 5.81868
R2360 VDD2.n145 VDD2.n101 5.04292
R2361 VDD2.n133 VDD2.n107 5.04292
R2362 VDD2.n44 VDD2.n18 5.04292
R2363 VDD2.n56 VDD2.n12 5.04292
R2364 VDD2.n149 VDD2.n148 4.26717
R2365 VDD2.n132 VDD2.n109 4.26717
R2366 VDD2.n43 VDD2.n20 4.26717
R2367 VDD2.n60 VDD2.n59 4.26717
R2368 VDD2.n116 VDD2.n114 3.70982
R2369 VDD2.n27 VDD2.n25 3.70982
R2370 VDD2.n152 VDD2.n99 3.49141
R2371 VDD2.n129 VDD2.n128 3.49141
R2372 VDD2.n40 VDD2.n39 3.49141
R2373 VDD2.n63 VDD2.n10 3.49141
R2374 VDD2.n171 VDD2.n87 2.71565
R2375 VDD2.n153 VDD2.n97 2.71565
R2376 VDD2.n125 VDD2.n111 2.71565
R2377 VDD2.n36 VDD2.n22 2.71565
R2378 VDD2.n64 VDD2.n8 2.71565
R2379 VDD2.n84 VDD2.n0 2.71565
R2380 VDD2.n173 VDD2.t0 2.10438
R2381 VDD2.n173 VDD2.t3 2.10438
R2382 VDD2.n85 VDD2.t5 2.10438
R2383 VDD2.n85 VDD2.t1 2.10438
R2384 VDD2 VDD2.n172 2.09533
R2385 VDD2.n169 VDD2.n168 1.93989
R2386 VDD2.n157 VDD2.n156 1.93989
R2387 VDD2.n124 VDD2.n113 1.93989
R2388 VDD2.n35 VDD2.n24 1.93989
R2389 VDD2.n69 VDD2.n67 1.93989
R2390 VDD2.n82 VDD2.n81 1.93989
R2391 VDD2.n165 VDD2.n89 1.16414
R2392 VDD2.n160 VDD2.n94 1.16414
R2393 VDD2.n121 VDD2.n120 1.16414
R2394 VDD2.n32 VDD2.n31 1.16414
R2395 VDD2.n68 VDD2.n6 1.16414
R2396 VDD2.n78 VDD2.n2 1.16414
R2397 VDD2.n164 VDD2.n91 0.388379
R2398 VDD2.n161 VDD2.n93 0.388379
R2399 VDD2.n117 VDD2.n115 0.388379
R2400 VDD2.n28 VDD2.n26 0.388379
R2401 VDD2.n74 VDD2.n73 0.388379
R2402 VDD2.n77 VDD2.n4 0.388379
R2403 VDD2.n170 VDD2.n88 0.155672
R2404 VDD2.n163 VDD2.n88 0.155672
R2405 VDD2.n163 VDD2.n162 0.155672
R2406 VDD2.n162 VDD2.n92 0.155672
R2407 VDD2.n155 VDD2.n92 0.155672
R2408 VDD2.n155 VDD2.n154 0.155672
R2409 VDD2.n154 VDD2.n98 0.155672
R2410 VDD2.n147 VDD2.n98 0.155672
R2411 VDD2.n147 VDD2.n146 0.155672
R2412 VDD2.n146 VDD2.n102 0.155672
R2413 VDD2.n139 VDD2.n102 0.155672
R2414 VDD2.n139 VDD2.n138 0.155672
R2415 VDD2.n138 VDD2.n106 0.155672
R2416 VDD2.n131 VDD2.n106 0.155672
R2417 VDD2.n131 VDD2.n130 0.155672
R2418 VDD2.n130 VDD2.n110 0.155672
R2419 VDD2.n123 VDD2.n110 0.155672
R2420 VDD2.n123 VDD2.n122 0.155672
R2421 VDD2.n122 VDD2.n114 0.155672
R2422 VDD2.n33 VDD2.n25 0.155672
R2423 VDD2.n34 VDD2.n33 0.155672
R2424 VDD2.n34 VDD2.n21 0.155672
R2425 VDD2.n41 VDD2.n21 0.155672
R2426 VDD2.n42 VDD2.n41 0.155672
R2427 VDD2.n42 VDD2.n17 0.155672
R2428 VDD2.n49 VDD2.n17 0.155672
R2429 VDD2.n50 VDD2.n49 0.155672
R2430 VDD2.n50 VDD2.n13 0.155672
R2431 VDD2.n57 VDD2.n13 0.155672
R2432 VDD2.n58 VDD2.n57 0.155672
R2433 VDD2.n58 VDD2.n9 0.155672
R2434 VDD2.n65 VDD2.n9 0.155672
R2435 VDD2.n66 VDD2.n65 0.155672
R2436 VDD2.n66 VDD2.n5 0.155672
R2437 VDD2.n75 VDD2.n5 0.155672
R2438 VDD2.n76 VDD2.n75 0.155672
R2439 VDD2.n76 VDD2.n1 0.155672
R2440 VDD2.n83 VDD2.n1 0.155672
C0 VDD2 B 2.50408f
C1 VDD1 VP 8.99642f
C2 VTAIL w_n3490_n4058# 3.47285f
C3 VN VDD2 8.67394f
C4 w_n3490_n4058# B 10.9474f
C5 VDD2 VP 0.477313f
C6 VN w_n3490_n4058# 6.73971f
C7 w_n3490_n4058# VP 7.19153f
C8 VDD1 VDD2 1.49372f
C9 VDD1 w_n3490_n4058# 2.58483f
C10 VTAIL B 4.56645f
C11 VDD2 w_n3490_n4058# 2.6769f
C12 VN VTAIL 8.72908f
C13 VTAIL VP 8.743401f
C14 VN B 1.25405f
C15 B VP 2.00952f
C16 VN VP 7.784709f
C17 VTAIL VDD1 8.990581f
C18 VDD1 B 2.42471f
C19 VTAIL VDD2 9.04237f
C20 VN VDD1 0.151124f
C21 VDD2 VSUBS 2.054896f
C22 VDD1 VSUBS 2.001587f
C23 VTAIL VSUBS 1.358085f
C24 VN VSUBS 6.18083f
C25 VP VSUBS 3.243813f
C26 B VSUBS 5.147926f
C27 w_n3490_n4058# VSUBS 0.173593p
C28 VDD2.n0 VSUBS 0.029228f
C29 VDD2.n1 VSUBS 0.027445f
C30 VDD2.n2 VSUBS 0.014748f
C31 VDD2.n3 VSUBS 0.034859f
C32 VDD2.n4 VSUBS 0.015182f
C33 VDD2.n5 VSUBS 0.027445f
C34 VDD2.n6 VSUBS 0.015616f
C35 VDD2.n7 VSUBS 0.034859f
C36 VDD2.n8 VSUBS 0.015616f
C37 VDD2.n9 VSUBS 0.027445f
C38 VDD2.n10 VSUBS 0.014748f
C39 VDD2.n11 VSUBS 0.034859f
C40 VDD2.n12 VSUBS 0.015616f
C41 VDD2.n13 VSUBS 0.027445f
C42 VDD2.n14 VSUBS 0.014748f
C43 VDD2.n15 VSUBS 0.034859f
C44 VDD2.n16 VSUBS 0.015616f
C45 VDD2.n17 VSUBS 0.027445f
C46 VDD2.n18 VSUBS 0.014748f
C47 VDD2.n19 VSUBS 0.034859f
C48 VDD2.n20 VSUBS 0.015616f
C49 VDD2.n21 VSUBS 0.027445f
C50 VDD2.n22 VSUBS 0.014748f
C51 VDD2.n23 VSUBS 0.034859f
C52 VDD2.n24 VSUBS 0.015616f
C53 VDD2.n25 VSUBS 1.80852f
C54 VDD2.n26 VSUBS 0.014748f
C55 VDD2.t4 VSUBS 0.074657f
C56 VDD2.n27 VSUBS 0.19711f
C57 VDD2.n28 VSUBS 0.022176f
C58 VDD2.n29 VSUBS 0.026144f
C59 VDD2.n30 VSUBS 0.034859f
C60 VDD2.n31 VSUBS 0.015616f
C61 VDD2.n32 VSUBS 0.014748f
C62 VDD2.n33 VSUBS 0.027445f
C63 VDD2.n34 VSUBS 0.027445f
C64 VDD2.n35 VSUBS 0.014748f
C65 VDD2.n36 VSUBS 0.015616f
C66 VDD2.n37 VSUBS 0.034859f
C67 VDD2.n38 VSUBS 0.034859f
C68 VDD2.n39 VSUBS 0.015616f
C69 VDD2.n40 VSUBS 0.014748f
C70 VDD2.n41 VSUBS 0.027445f
C71 VDD2.n42 VSUBS 0.027445f
C72 VDD2.n43 VSUBS 0.014748f
C73 VDD2.n44 VSUBS 0.015616f
C74 VDD2.n45 VSUBS 0.034859f
C75 VDD2.n46 VSUBS 0.034859f
C76 VDD2.n47 VSUBS 0.015616f
C77 VDD2.n48 VSUBS 0.014748f
C78 VDD2.n49 VSUBS 0.027445f
C79 VDD2.n50 VSUBS 0.027445f
C80 VDD2.n51 VSUBS 0.014748f
C81 VDD2.n52 VSUBS 0.015616f
C82 VDD2.n53 VSUBS 0.034859f
C83 VDD2.n54 VSUBS 0.034859f
C84 VDD2.n55 VSUBS 0.015616f
C85 VDD2.n56 VSUBS 0.014748f
C86 VDD2.n57 VSUBS 0.027445f
C87 VDD2.n58 VSUBS 0.027445f
C88 VDD2.n59 VSUBS 0.014748f
C89 VDD2.n60 VSUBS 0.015616f
C90 VDD2.n61 VSUBS 0.034859f
C91 VDD2.n62 VSUBS 0.034859f
C92 VDD2.n63 VSUBS 0.015616f
C93 VDD2.n64 VSUBS 0.014748f
C94 VDD2.n65 VSUBS 0.027445f
C95 VDD2.n66 VSUBS 0.027445f
C96 VDD2.n67 VSUBS 0.014748f
C97 VDD2.n68 VSUBS 0.014748f
C98 VDD2.n69 VSUBS 0.015616f
C99 VDD2.n70 VSUBS 0.034859f
C100 VDD2.n71 VSUBS 0.034859f
C101 VDD2.n72 VSUBS 0.034859f
C102 VDD2.n73 VSUBS 0.015182f
C103 VDD2.n74 VSUBS 0.014748f
C104 VDD2.n75 VSUBS 0.027445f
C105 VDD2.n76 VSUBS 0.027445f
C106 VDD2.n77 VSUBS 0.014748f
C107 VDD2.n78 VSUBS 0.015616f
C108 VDD2.n79 VSUBS 0.034859f
C109 VDD2.n80 VSUBS 0.081225f
C110 VDD2.n81 VSUBS 0.015616f
C111 VDD2.n82 VSUBS 0.014748f
C112 VDD2.n83 VSUBS 0.066813f
C113 VDD2.n84 VSUBS 0.06841f
C114 VDD2.t5 VSUBS 0.335084f
C115 VDD2.t1 VSUBS 0.335084f
C116 VDD2.n85 VSUBS 2.74402f
C117 VDD2.n86 VSUBS 3.57568f
C118 VDD2.n87 VSUBS 0.029228f
C119 VDD2.n88 VSUBS 0.027445f
C120 VDD2.n89 VSUBS 0.014748f
C121 VDD2.n90 VSUBS 0.034859f
C122 VDD2.n91 VSUBS 0.015182f
C123 VDD2.n92 VSUBS 0.027445f
C124 VDD2.n93 VSUBS 0.015182f
C125 VDD2.n94 VSUBS 0.014748f
C126 VDD2.n95 VSUBS 0.034859f
C127 VDD2.n96 VSUBS 0.034859f
C128 VDD2.n97 VSUBS 0.015616f
C129 VDD2.n98 VSUBS 0.027445f
C130 VDD2.n99 VSUBS 0.014748f
C131 VDD2.n100 VSUBS 0.034859f
C132 VDD2.n101 VSUBS 0.015616f
C133 VDD2.n102 VSUBS 0.027445f
C134 VDD2.n103 VSUBS 0.014748f
C135 VDD2.n104 VSUBS 0.034859f
C136 VDD2.n105 VSUBS 0.015616f
C137 VDD2.n106 VSUBS 0.027445f
C138 VDD2.n107 VSUBS 0.014748f
C139 VDD2.n108 VSUBS 0.034859f
C140 VDD2.n109 VSUBS 0.015616f
C141 VDD2.n110 VSUBS 0.027445f
C142 VDD2.n111 VSUBS 0.014748f
C143 VDD2.n112 VSUBS 0.034859f
C144 VDD2.n113 VSUBS 0.015616f
C145 VDD2.n114 VSUBS 1.80852f
C146 VDD2.n115 VSUBS 0.014748f
C147 VDD2.t2 VSUBS 0.074657f
C148 VDD2.n116 VSUBS 0.19711f
C149 VDD2.n117 VSUBS 0.022176f
C150 VDD2.n118 VSUBS 0.026144f
C151 VDD2.n119 VSUBS 0.034859f
C152 VDD2.n120 VSUBS 0.015616f
C153 VDD2.n121 VSUBS 0.014748f
C154 VDD2.n122 VSUBS 0.027445f
C155 VDD2.n123 VSUBS 0.027445f
C156 VDD2.n124 VSUBS 0.014748f
C157 VDD2.n125 VSUBS 0.015616f
C158 VDD2.n126 VSUBS 0.034859f
C159 VDD2.n127 VSUBS 0.034859f
C160 VDD2.n128 VSUBS 0.015616f
C161 VDD2.n129 VSUBS 0.014748f
C162 VDD2.n130 VSUBS 0.027445f
C163 VDD2.n131 VSUBS 0.027445f
C164 VDD2.n132 VSUBS 0.014748f
C165 VDD2.n133 VSUBS 0.015616f
C166 VDD2.n134 VSUBS 0.034859f
C167 VDD2.n135 VSUBS 0.034859f
C168 VDD2.n136 VSUBS 0.015616f
C169 VDD2.n137 VSUBS 0.014748f
C170 VDD2.n138 VSUBS 0.027445f
C171 VDD2.n139 VSUBS 0.027445f
C172 VDD2.n140 VSUBS 0.014748f
C173 VDD2.n141 VSUBS 0.015616f
C174 VDD2.n142 VSUBS 0.034859f
C175 VDD2.n143 VSUBS 0.034859f
C176 VDD2.n144 VSUBS 0.015616f
C177 VDD2.n145 VSUBS 0.014748f
C178 VDD2.n146 VSUBS 0.027445f
C179 VDD2.n147 VSUBS 0.027445f
C180 VDD2.n148 VSUBS 0.014748f
C181 VDD2.n149 VSUBS 0.015616f
C182 VDD2.n150 VSUBS 0.034859f
C183 VDD2.n151 VSUBS 0.034859f
C184 VDD2.n152 VSUBS 0.015616f
C185 VDD2.n153 VSUBS 0.014748f
C186 VDD2.n154 VSUBS 0.027445f
C187 VDD2.n155 VSUBS 0.027445f
C188 VDD2.n156 VSUBS 0.014748f
C189 VDD2.n157 VSUBS 0.015616f
C190 VDD2.n158 VSUBS 0.034859f
C191 VDD2.n159 VSUBS 0.034859f
C192 VDD2.n160 VSUBS 0.015616f
C193 VDD2.n161 VSUBS 0.014748f
C194 VDD2.n162 VSUBS 0.027445f
C195 VDD2.n163 VSUBS 0.027445f
C196 VDD2.n164 VSUBS 0.014748f
C197 VDD2.n165 VSUBS 0.015616f
C198 VDD2.n166 VSUBS 0.034859f
C199 VDD2.n167 VSUBS 0.081225f
C200 VDD2.n168 VSUBS 0.015616f
C201 VDD2.n169 VSUBS 0.014748f
C202 VDD2.n170 VSUBS 0.066813f
C203 VDD2.n171 VSUBS 0.059733f
C204 VDD2.n172 VSUBS 3.17015f
C205 VDD2.t0 VSUBS 0.335084f
C206 VDD2.t3 VSUBS 0.335084f
C207 VDD2.n173 VSUBS 2.74398f
C208 VN.t4 VSUBS 3.23901f
C209 VN.n0 VSUBS 1.22909f
C210 VN.n1 VSUBS 0.027112f
C211 VN.n2 VSUBS 0.045248f
C212 VN.n3 VSUBS 0.287683f
C213 VN.t0 VSUBS 3.23901f
C214 VN.t1 VSUBS 3.49095f
C215 VN.n4 VSUBS 1.1801f
C216 VN.n5 VSUBS 1.2117f
C217 VN.n6 VSUBS 0.038057f
C218 VN.n7 VSUBS 0.05053f
C219 VN.n8 VSUBS 0.027112f
C220 VN.n9 VSUBS 0.027112f
C221 VN.n10 VSUBS 0.027112f
C222 VN.n11 VSUBS 0.033915f
C223 VN.n12 VSUBS 0.05053f
C224 VN.n13 VSUBS 0.045541f
C225 VN.n14 VSUBS 0.043759f
C226 VN.n15 VSUBS 0.055307f
C227 VN.t3 VSUBS 3.23901f
C228 VN.n16 VSUBS 1.22909f
C229 VN.n17 VSUBS 0.027112f
C230 VN.n18 VSUBS 0.045248f
C231 VN.n19 VSUBS 0.287683f
C232 VN.t5 VSUBS 3.23901f
C233 VN.t2 VSUBS 3.49095f
C234 VN.n20 VSUBS 1.1801f
C235 VN.n21 VSUBS 1.2117f
C236 VN.n22 VSUBS 0.038057f
C237 VN.n23 VSUBS 0.05053f
C238 VN.n24 VSUBS 0.027112f
C239 VN.n25 VSUBS 0.027112f
C240 VN.n26 VSUBS 0.027112f
C241 VN.n27 VSUBS 0.033915f
C242 VN.n28 VSUBS 0.05053f
C243 VN.n29 VSUBS 0.045541f
C244 VN.n30 VSUBS 0.043759f
C245 VN.n31 VSUBS 1.63899f
C246 VDD1.n0 VSUBS 0.029226f
C247 VDD1.n1 VSUBS 0.027444f
C248 VDD1.n2 VSUBS 0.014747f
C249 VDD1.n3 VSUBS 0.034857f
C250 VDD1.n4 VSUBS 0.015181f
C251 VDD1.n5 VSUBS 0.027444f
C252 VDD1.n6 VSUBS 0.015181f
C253 VDD1.n7 VSUBS 0.014747f
C254 VDD1.n8 VSUBS 0.034857f
C255 VDD1.n9 VSUBS 0.034857f
C256 VDD1.n10 VSUBS 0.015615f
C257 VDD1.n11 VSUBS 0.027444f
C258 VDD1.n12 VSUBS 0.014747f
C259 VDD1.n13 VSUBS 0.034857f
C260 VDD1.n14 VSUBS 0.015615f
C261 VDD1.n15 VSUBS 0.027444f
C262 VDD1.n16 VSUBS 0.014747f
C263 VDD1.n17 VSUBS 0.034857f
C264 VDD1.n18 VSUBS 0.015615f
C265 VDD1.n19 VSUBS 0.027444f
C266 VDD1.n20 VSUBS 0.014747f
C267 VDD1.n21 VSUBS 0.034857f
C268 VDD1.n22 VSUBS 0.015615f
C269 VDD1.n23 VSUBS 0.027444f
C270 VDD1.n24 VSUBS 0.014747f
C271 VDD1.n25 VSUBS 0.034857f
C272 VDD1.n26 VSUBS 0.015615f
C273 VDD1.n27 VSUBS 1.80841f
C274 VDD1.n28 VSUBS 0.014747f
C275 VDD1.t4 VSUBS 0.074652f
C276 VDD1.n29 VSUBS 0.197098f
C277 VDD1.n30 VSUBS 0.022174f
C278 VDD1.n31 VSUBS 0.026143f
C279 VDD1.n32 VSUBS 0.034857f
C280 VDD1.n33 VSUBS 0.015615f
C281 VDD1.n34 VSUBS 0.014747f
C282 VDD1.n35 VSUBS 0.027444f
C283 VDD1.n36 VSUBS 0.027444f
C284 VDD1.n37 VSUBS 0.014747f
C285 VDD1.n38 VSUBS 0.015615f
C286 VDD1.n39 VSUBS 0.034857f
C287 VDD1.n40 VSUBS 0.034857f
C288 VDD1.n41 VSUBS 0.015615f
C289 VDD1.n42 VSUBS 0.014747f
C290 VDD1.n43 VSUBS 0.027444f
C291 VDD1.n44 VSUBS 0.027444f
C292 VDD1.n45 VSUBS 0.014747f
C293 VDD1.n46 VSUBS 0.015615f
C294 VDD1.n47 VSUBS 0.034857f
C295 VDD1.n48 VSUBS 0.034857f
C296 VDD1.n49 VSUBS 0.015615f
C297 VDD1.n50 VSUBS 0.014747f
C298 VDD1.n51 VSUBS 0.027444f
C299 VDD1.n52 VSUBS 0.027444f
C300 VDD1.n53 VSUBS 0.014747f
C301 VDD1.n54 VSUBS 0.015615f
C302 VDD1.n55 VSUBS 0.034857f
C303 VDD1.n56 VSUBS 0.034857f
C304 VDD1.n57 VSUBS 0.015615f
C305 VDD1.n58 VSUBS 0.014747f
C306 VDD1.n59 VSUBS 0.027444f
C307 VDD1.n60 VSUBS 0.027444f
C308 VDD1.n61 VSUBS 0.014747f
C309 VDD1.n62 VSUBS 0.015615f
C310 VDD1.n63 VSUBS 0.034857f
C311 VDD1.n64 VSUBS 0.034857f
C312 VDD1.n65 VSUBS 0.015615f
C313 VDD1.n66 VSUBS 0.014747f
C314 VDD1.n67 VSUBS 0.027444f
C315 VDD1.n68 VSUBS 0.027444f
C316 VDD1.n69 VSUBS 0.014747f
C317 VDD1.n70 VSUBS 0.015615f
C318 VDD1.n71 VSUBS 0.034857f
C319 VDD1.n72 VSUBS 0.034857f
C320 VDD1.n73 VSUBS 0.015615f
C321 VDD1.n74 VSUBS 0.014747f
C322 VDD1.n75 VSUBS 0.027444f
C323 VDD1.n76 VSUBS 0.027444f
C324 VDD1.n77 VSUBS 0.014747f
C325 VDD1.n78 VSUBS 0.015615f
C326 VDD1.n79 VSUBS 0.034857f
C327 VDD1.n80 VSUBS 0.08122f
C328 VDD1.n81 VSUBS 0.015615f
C329 VDD1.n82 VSUBS 0.014747f
C330 VDD1.n83 VSUBS 0.066809f
C331 VDD1.n84 VSUBS 0.06927f
C332 VDD1.n85 VSUBS 0.029226f
C333 VDD1.n86 VSUBS 0.027444f
C334 VDD1.n87 VSUBS 0.014747f
C335 VDD1.n88 VSUBS 0.034857f
C336 VDD1.n89 VSUBS 0.015181f
C337 VDD1.n90 VSUBS 0.027444f
C338 VDD1.n91 VSUBS 0.015615f
C339 VDD1.n92 VSUBS 0.034857f
C340 VDD1.n93 VSUBS 0.015615f
C341 VDD1.n94 VSUBS 0.027444f
C342 VDD1.n95 VSUBS 0.014747f
C343 VDD1.n96 VSUBS 0.034857f
C344 VDD1.n97 VSUBS 0.015615f
C345 VDD1.n98 VSUBS 0.027444f
C346 VDD1.n99 VSUBS 0.014747f
C347 VDD1.n100 VSUBS 0.034857f
C348 VDD1.n101 VSUBS 0.015615f
C349 VDD1.n102 VSUBS 0.027444f
C350 VDD1.n103 VSUBS 0.014747f
C351 VDD1.n104 VSUBS 0.034857f
C352 VDD1.n105 VSUBS 0.015615f
C353 VDD1.n106 VSUBS 0.027444f
C354 VDD1.n107 VSUBS 0.014747f
C355 VDD1.n108 VSUBS 0.034857f
C356 VDD1.n109 VSUBS 0.015615f
C357 VDD1.n110 VSUBS 1.80841f
C358 VDD1.n111 VSUBS 0.014747f
C359 VDD1.t3 VSUBS 0.074652f
C360 VDD1.n112 VSUBS 0.197098f
C361 VDD1.n113 VSUBS 0.022174f
C362 VDD1.n114 VSUBS 0.026143f
C363 VDD1.n115 VSUBS 0.034857f
C364 VDD1.n116 VSUBS 0.015615f
C365 VDD1.n117 VSUBS 0.014747f
C366 VDD1.n118 VSUBS 0.027444f
C367 VDD1.n119 VSUBS 0.027444f
C368 VDD1.n120 VSUBS 0.014747f
C369 VDD1.n121 VSUBS 0.015615f
C370 VDD1.n122 VSUBS 0.034857f
C371 VDD1.n123 VSUBS 0.034857f
C372 VDD1.n124 VSUBS 0.015615f
C373 VDD1.n125 VSUBS 0.014747f
C374 VDD1.n126 VSUBS 0.027444f
C375 VDD1.n127 VSUBS 0.027444f
C376 VDD1.n128 VSUBS 0.014747f
C377 VDD1.n129 VSUBS 0.015615f
C378 VDD1.n130 VSUBS 0.034857f
C379 VDD1.n131 VSUBS 0.034857f
C380 VDD1.n132 VSUBS 0.015615f
C381 VDD1.n133 VSUBS 0.014747f
C382 VDD1.n134 VSUBS 0.027444f
C383 VDD1.n135 VSUBS 0.027444f
C384 VDD1.n136 VSUBS 0.014747f
C385 VDD1.n137 VSUBS 0.015615f
C386 VDD1.n138 VSUBS 0.034857f
C387 VDD1.n139 VSUBS 0.034857f
C388 VDD1.n140 VSUBS 0.015615f
C389 VDD1.n141 VSUBS 0.014747f
C390 VDD1.n142 VSUBS 0.027444f
C391 VDD1.n143 VSUBS 0.027444f
C392 VDD1.n144 VSUBS 0.014747f
C393 VDD1.n145 VSUBS 0.015615f
C394 VDD1.n146 VSUBS 0.034857f
C395 VDD1.n147 VSUBS 0.034857f
C396 VDD1.n148 VSUBS 0.015615f
C397 VDD1.n149 VSUBS 0.014747f
C398 VDD1.n150 VSUBS 0.027444f
C399 VDD1.n151 VSUBS 0.027444f
C400 VDD1.n152 VSUBS 0.014747f
C401 VDD1.n153 VSUBS 0.014747f
C402 VDD1.n154 VSUBS 0.015615f
C403 VDD1.n155 VSUBS 0.034857f
C404 VDD1.n156 VSUBS 0.034857f
C405 VDD1.n157 VSUBS 0.034857f
C406 VDD1.n158 VSUBS 0.015181f
C407 VDD1.n159 VSUBS 0.014747f
C408 VDD1.n160 VSUBS 0.027444f
C409 VDD1.n161 VSUBS 0.027444f
C410 VDD1.n162 VSUBS 0.014747f
C411 VDD1.n163 VSUBS 0.015615f
C412 VDD1.n164 VSUBS 0.034857f
C413 VDD1.n165 VSUBS 0.08122f
C414 VDD1.n166 VSUBS 0.015615f
C415 VDD1.n167 VSUBS 0.014747f
C416 VDD1.n168 VSUBS 0.066809f
C417 VDD1.n169 VSUBS 0.068406f
C418 VDD1.t2 VSUBS 0.335064f
C419 VDD1.t0 VSUBS 0.335064f
C420 VDD1.n170 VSUBS 2.74386f
C421 VDD1.n171 VSUBS 3.72085f
C422 VDD1.t1 VSUBS 0.335064f
C423 VDD1.t5 VSUBS 0.335064f
C424 VDD1.n172 VSUBS 2.73674f
C425 VDD1.n173 VSUBS 3.71326f
C426 VTAIL.t5 VSUBS 0.34447f
C427 VTAIL.t3 VSUBS 0.34447f
C428 VTAIL.n0 VSUBS 2.65363f
C429 VTAIL.n1 VSUBS 0.89066f
C430 VTAIL.n2 VSUBS 0.030046f
C431 VTAIL.n3 VSUBS 0.028214f
C432 VTAIL.n4 VSUBS 0.015161f
C433 VTAIL.n5 VSUBS 0.035835f
C434 VTAIL.n6 VSUBS 0.015607f
C435 VTAIL.n7 VSUBS 0.028214f
C436 VTAIL.n8 VSUBS 0.016053f
C437 VTAIL.n9 VSUBS 0.035835f
C438 VTAIL.n10 VSUBS 0.016053f
C439 VTAIL.n11 VSUBS 0.028214f
C440 VTAIL.n12 VSUBS 0.015161f
C441 VTAIL.n13 VSUBS 0.035835f
C442 VTAIL.n14 VSUBS 0.016053f
C443 VTAIL.n15 VSUBS 0.028214f
C444 VTAIL.n16 VSUBS 0.015161f
C445 VTAIL.n17 VSUBS 0.035835f
C446 VTAIL.n18 VSUBS 0.016053f
C447 VTAIL.n19 VSUBS 0.028214f
C448 VTAIL.n20 VSUBS 0.015161f
C449 VTAIL.n21 VSUBS 0.035835f
C450 VTAIL.n22 VSUBS 0.016053f
C451 VTAIL.n23 VSUBS 0.028214f
C452 VTAIL.n24 VSUBS 0.015161f
C453 VTAIL.n25 VSUBS 0.035835f
C454 VTAIL.n26 VSUBS 0.016053f
C455 VTAIL.n27 VSUBS 1.85918f
C456 VTAIL.n28 VSUBS 0.015161f
C457 VTAIL.t9 VSUBS 0.076748f
C458 VTAIL.n29 VSUBS 0.202631f
C459 VTAIL.n30 VSUBS 0.022797f
C460 VTAIL.n31 VSUBS 0.026877f
C461 VTAIL.n32 VSUBS 0.035835f
C462 VTAIL.n33 VSUBS 0.016053f
C463 VTAIL.n34 VSUBS 0.015161f
C464 VTAIL.n35 VSUBS 0.028214f
C465 VTAIL.n36 VSUBS 0.028214f
C466 VTAIL.n37 VSUBS 0.015161f
C467 VTAIL.n38 VSUBS 0.016053f
C468 VTAIL.n39 VSUBS 0.035835f
C469 VTAIL.n40 VSUBS 0.035835f
C470 VTAIL.n41 VSUBS 0.016053f
C471 VTAIL.n42 VSUBS 0.015161f
C472 VTAIL.n43 VSUBS 0.028214f
C473 VTAIL.n44 VSUBS 0.028214f
C474 VTAIL.n45 VSUBS 0.015161f
C475 VTAIL.n46 VSUBS 0.016053f
C476 VTAIL.n47 VSUBS 0.035835f
C477 VTAIL.n48 VSUBS 0.035835f
C478 VTAIL.n49 VSUBS 0.016053f
C479 VTAIL.n50 VSUBS 0.015161f
C480 VTAIL.n51 VSUBS 0.028214f
C481 VTAIL.n52 VSUBS 0.028214f
C482 VTAIL.n53 VSUBS 0.015161f
C483 VTAIL.n54 VSUBS 0.016053f
C484 VTAIL.n55 VSUBS 0.035835f
C485 VTAIL.n56 VSUBS 0.035835f
C486 VTAIL.n57 VSUBS 0.016053f
C487 VTAIL.n58 VSUBS 0.015161f
C488 VTAIL.n59 VSUBS 0.028214f
C489 VTAIL.n60 VSUBS 0.028214f
C490 VTAIL.n61 VSUBS 0.015161f
C491 VTAIL.n62 VSUBS 0.016053f
C492 VTAIL.n63 VSUBS 0.035835f
C493 VTAIL.n64 VSUBS 0.035835f
C494 VTAIL.n65 VSUBS 0.016053f
C495 VTAIL.n66 VSUBS 0.015161f
C496 VTAIL.n67 VSUBS 0.028214f
C497 VTAIL.n68 VSUBS 0.028214f
C498 VTAIL.n69 VSUBS 0.015161f
C499 VTAIL.n70 VSUBS 0.015161f
C500 VTAIL.n71 VSUBS 0.016053f
C501 VTAIL.n72 VSUBS 0.035835f
C502 VTAIL.n73 VSUBS 0.035835f
C503 VTAIL.n74 VSUBS 0.035835f
C504 VTAIL.n75 VSUBS 0.015607f
C505 VTAIL.n76 VSUBS 0.015161f
C506 VTAIL.n77 VSUBS 0.028214f
C507 VTAIL.n78 VSUBS 0.028214f
C508 VTAIL.n79 VSUBS 0.015161f
C509 VTAIL.n80 VSUBS 0.016053f
C510 VTAIL.n81 VSUBS 0.035835f
C511 VTAIL.n82 VSUBS 0.0835f
C512 VTAIL.n83 VSUBS 0.016053f
C513 VTAIL.n84 VSUBS 0.015161f
C514 VTAIL.n85 VSUBS 0.068685f
C515 VTAIL.n86 VSUBS 0.041951f
C516 VTAIL.n87 VSUBS 0.439084f
C517 VTAIL.t6 VSUBS 0.34447f
C518 VTAIL.t7 VSUBS 0.34447f
C519 VTAIL.n88 VSUBS 2.65363f
C520 VTAIL.n89 VSUBS 2.99225f
C521 VTAIL.t0 VSUBS 0.34447f
C522 VTAIL.t4 VSUBS 0.34447f
C523 VTAIL.n90 VSUBS 2.65365f
C524 VTAIL.n91 VSUBS 2.99223f
C525 VTAIL.n92 VSUBS 0.030046f
C526 VTAIL.n93 VSUBS 0.028214f
C527 VTAIL.n94 VSUBS 0.015161f
C528 VTAIL.n95 VSUBS 0.035835f
C529 VTAIL.n96 VSUBS 0.015607f
C530 VTAIL.n97 VSUBS 0.028214f
C531 VTAIL.n98 VSUBS 0.015607f
C532 VTAIL.n99 VSUBS 0.015161f
C533 VTAIL.n100 VSUBS 0.035835f
C534 VTAIL.n101 VSUBS 0.035835f
C535 VTAIL.n102 VSUBS 0.016053f
C536 VTAIL.n103 VSUBS 0.028214f
C537 VTAIL.n104 VSUBS 0.015161f
C538 VTAIL.n105 VSUBS 0.035835f
C539 VTAIL.n106 VSUBS 0.016053f
C540 VTAIL.n107 VSUBS 0.028214f
C541 VTAIL.n108 VSUBS 0.015161f
C542 VTAIL.n109 VSUBS 0.035835f
C543 VTAIL.n110 VSUBS 0.016053f
C544 VTAIL.n111 VSUBS 0.028214f
C545 VTAIL.n112 VSUBS 0.015161f
C546 VTAIL.n113 VSUBS 0.035835f
C547 VTAIL.n114 VSUBS 0.016053f
C548 VTAIL.n115 VSUBS 0.028214f
C549 VTAIL.n116 VSUBS 0.015161f
C550 VTAIL.n117 VSUBS 0.035835f
C551 VTAIL.n118 VSUBS 0.016053f
C552 VTAIL.n119 VSUBS 1.85918f
C553 VTAIL.n120 VSUBS 0.015161f
C554 VTAIL.t1 VSUBS 0.076748f
C555 VTAIL.n121 VSUBS 0.202631f
C556 VTAIL.n122 VSUBS 0.022797f
C557 VTAIL.n123 VSUBS 0.026877f
C558 VTAIL.n124 VSUBS 0.035835f
C559 VTAIL.n125 VSUBS 0.016053f
C560 VTAIL.n126 VSUBS 0.015161f
C561 VTAIL.n127 VSUBS 0.028214f
C562 VTAIL.n128 VSUBS 0.028214f
C563 VTAIL.n129 VSUBS 0.015161f
C564 VTAIL.n130 VSUBS 0.016053f
C565 VTAIL.n131 VSUBS 0.035835f
C566 VTAIL.n132 VSUBS 0.035835f
C567 VTAIL.n133 VSUBS 0.016053f
C568 VTAIL.n134 VSUBS 0.015161f
C569 VTAIL.n135 VSUBS 0.028214f
C570 VTAIL.n136 VSUBS 0.028214f
C571 VTAIL.n137 VSUBS 0.015161f
C572 VTAIL.n138 VSUBS 0.016053f
C573 VTAIL.n139 VSUBS 0.035835f
C574 VTAIL.n140 VSUBS 0.035835f
C575 VTAIL.n141 VSUBS 0.016053f
C576 VTAIL.n142 VSUBS 0.015161f
C577 VTAIL.n143 VSUBS 0.028214f
C578 VTAIL.n144 VSUBS 0.028214f
C579 VTAIL.n145 VSUBS 0.015161f
C580 VTAIL.n146 VSUBS 0.016053f
C581 VTAIL.n147 VSUBS 0.035835f
C582 VTAIL.n148 VSUBS 0.035835f
C583 VTAIL.n149 VSUBS 0.016053f
C584 VTAIL.n150 VSUBS 0.015161f
C585 VTAIL.n151 VSUBS 0.028214f
C586 VTAIL.n152 VSUBS 0.028214f
C587 VTAIL.n153 VSUBS 0.015161f
C588 VTAIL.n154 VSUBS 0.016053f
C589 VTAIL.n155 VSUBS 0.035835f
C590 VTAIL.n156 VSUBS 0.035835f
C591 VTAIL.n157 VSUBS 0.016053f
C592 VTAIL.n158 VSUBS 0.015161f
C593 VTAIL.n159 VSUBS 0.028214f
C594 VTAIL.n160 VSUBS 0.028214f
C595 VTAIL.n161 VSUBS 0.015161f
C596 VTAIL.n162 VSUBS 0.016053f
C597 VTAIL.n163 VSUBS 0.035835f
C598 VTAIL.n164 VSUBS 0.035835f
C599 VTAIL.n165 VSUBS 0.016053f
C600 VTAIL.n166 VSUBS 0.015161f
C601 VTAIL.n167 VSUBS 0.028214f
C602 VTAIL.n168 VSUBS 0.028214f
C603 VTAIL.n169 VSUBS 0.015161f
C604 VTAIL.n170 VSUBS 0.016053f
C605 VTAIL.n171 VSUBS 0.035835f
C606 VTAIL.n172 VSUBS 0.0835f
C607 VTAIL.n173 VSUBS 0.016053f
C608 VTAIL.n174 VSUBS 0.015161f
C609 VTAIL.n175 VSUBS 0.068685f
C610 VTAIL.n176 VSUBS 0.041951f
C611 VTAIL.n177 VSUBS 0.439084f
C612 VTAIL.t8 VSUBS 0.34447f
C613 VTAIL.t11 VSUBS 0.34447f
C614 VTAIL.n178 VSUBS 2.65365f
C615 VTAIL.n179 VSUBS 1.07051f
C616 VTAIL.n180 VSUBS 0.030046f
C617 VTAIL.n181 VSUBS 0.028214f
C618 VTAIL.n182 VSUBS 0.015161f
C619 VTAIL.n183 VSUBS 0.035835f
C620 VTAIL.n184 VSUBS 0.015607f
C621 VTAIL.n185 VSUBS 0.028214f
C622 VTAIL.n186 VSUBS 0.015607f
C623 VTAIL.n187 VSUBS 0.015161f
C624 VTAIL.n188 VSUBS 0.035835f
C625 VTAIL.n189 VSUBS 0.035835f
C626 VTAIL.n190 VSUBS 0.016053f
C627 VTAIL.n191 VSUBS 0.028214f
C628 VTAIL.n192 VSUBS 0.015161f
C629 VTAIL.n193 VSUBS 0.035835f
C630 VTAIL.n194 VSUBS 0.016053f
C631 VTAIL.n195 VSUBS 0.028214f
C632 VTAIL.n196 VSUBS 0.015161f
C633 VTAIL.n197 VSUBS 0.035835f
C634 VTAIL.n198 VSUBS 0.016053f
C635 VTAIL.n199 VSUBS 0.028214f
C636 VTAIL.n200 VSUBS 0.015161f
C637 VTAIL.n201 VSUBS 0.035835f
C638 VTAIL.n202 VSUBS 0.016053f
C639 VTAIL.n203 VSUBS 0.028214f
C640 VTAIL.n204 VSUBS 0.015161f
C641 VTAIL.n205 VSUBS 0.035835f
C642 VTAIL.n206 VSUBS 0.016053f
C643 VTAIL.n207 VSUBS 1.85918f
C644 VTAIL.n208 VSUBS 0.015161f
C645 VTAIL.t10 VSUBS 0.076748f
C646 VTAIL.n209 VSUBS 0.202631f
C647 VTAIL.n210 VSUBS 0.022797f
C648 VTAIL.n211 VSUBS 0.026877f
C649 VTAIL.n212 VSUBS 0.035835f
C650 VTAIL.n213 VSUBS 0.016053f
C651 VTAIL.n214 VSUBS 0.015161f
C652 VTAIL.n215 VSUBS 0.028214f
C653 VTAIL.n216 VSUBS 0.028214f
C654 VTAIL.n217 VSUBS 0.015161f
C655 VTAIL.n218 VSUBS 0.016053f
C656 VTAIL.n219 VSUBS 0.035835f
C657 VTAIL.n220 VSUBS 0.035835f
C658 VTAIL.n221 VSUBS 0.016053f
C659 VTAIL.n222 VSUBS 0.015161f
C660 VTAIL.n223 VSUBS 0.028214f
C661 VTAIL.n224 VSUBS 0.028214f
C662 VTAIL.n225 VSUBS 0.015161f
C663 VTAIL.n226 VSUBS 0.016053f
C664 VTAIL.n227 VSUBS 0.035835f
C665 VTAIL.n228 VSUBS 0.035835f
C666 VTAIL.n229 VSUBS 0.016053f
C667 VTAIL.n230 VSUBS 0.015161f
C668 VTAIL.n231 VSUBS 0.028214f
C669 VTAIL.n232 VSUBS 0.028214f
C670 VTAIL.n233 VSUBS 0.015161f
C671 VTAIL.n234 VSUBS 0.016053f
C672 VTAIL.n235 VSUBS 0.035835f
C673 VTAIL.n236 VSUBS 0.035835f
C674 VTAIL.n237 VSUBS 0.016053f
C675 VTAIL.n238 VSUBS 0.015161f
C676 VTAIL.n239 VSUBS 0.028214f
C677 VTAIL.n240 VSUBS 0.028214f
C678 VTAIL.n241 VSUBS 0.015161f
C679 VTAIL.n242 VSUBS 0.016053f
C680 VTAIL.n243 VSUBS 0.035835f
C681 VTAIL.n244 VSUBS 0.035835f
C682 VTAIL.n245 VSUBS 0.016053f
C683 VTAIL.n246 VSUBS 0.015161f
C684 VTAIL.n247 VSUBS 0.028214f
C685 VTAIL.n248 VSUBS 0.028214f
C686 VTAIL.n249 VSUBS 0.015161f
C687 VTAIL.n250 VSUBS 0.016053f
C688 VTAIL.n251 VSUBS 0.035835f
C689 VTAIL.n252 VSUBS 0.035835f
C690 VTAIL.n253 VSUBS 0.016053f
C691 VTAIL.n254 VSUBS 0.015161f
C692 VTAIL.n255 VSUBS 0.028214f
C693 VTAIL.n256 VSUBS 0.028214f
C694 VTAIL.n257 VSUBS 0.015161f
C695 VTAIL.n258 VSUBS 0.016053f
C696 VTAIL.n259 VSUBS 0.035835f
C697 VTAIL.n260 VSUBS 0.0835f
C698 VTAIL.n261 VSUBS 0.016053f
C699 VTAIL.n262 VSUBS 0.015161f
C700 VTAIL.n263 VSUBS 0.068685f
C701 VTAIL.n264 VSUBS 0.041951f
C702 VTAIL.n265 VSUBS 2.11393f
C703 VTAIL.n266 VSUBS 0.030046f
C704 VTAIL.n267 VSUBS 0.028214f
C705 VTAIL.n268 VSUBS 0.015161f
C706 VTAIL.n269 VSUBS 0.035835f
C707 VTAIL.n270 VSUBS 0.015607f
C708 VTAIL.n271 VSUBS 0.028214f
C709 VTAIL.n272 VSUBS 0.016053f
C710 VTAIL.n273 VSUBS 0.035835f
C711 VTAIL.n274 VSUBS 0.016053f
C712 VTAIL.n275 VSUBS 0.028214f
C713 VTAIL.n276 VSUBS 0.015161f
C714 VTAIL.n277 VSUBS 0.035835f
C715 VTAIL.n278 VSUBS 0.016053f
C716 VTAIL.n279 VSUBS 0.028214f
C717 VTAIL.n280 VSUBS 0.015161f
C718 VTAIL.n281 VSUBS 0.035835f
C719 VTAIL.n282 VSUBS 0.016053f
C720 VTAIL.n283 VSUBS 0.028214f
C721 VTAIL.n284 VSUBS 0.015161f
C722 VTAIL.n285 VSUBS 0.035835f
C723 VTAIL.n286 VSUBS 0.016053f
C724 VTAIL.n287 VSUBS 0.028214f
C725 VTAIL.n288 VSUBS 0.015161f
C726 VTAIL.n289 VSUBS 0.035835f
C727 VTAIL.n290 VSUBS 0.016053f
C728 VTAIL.n291 VSUBS 1.85918f
C729 VTAIL.n292 VSUBS 0.015161f
C730 VTAIL.t2 VSUBS 0.076748f
C731 VTAIL.n293 VSUBS 0.202631f
C732 VTAIL.n294 VSUBS 0.022797f
C733 VTAIL.n295 VSUBS 0.026877f
C734 VTAIL.n296 VSUBS 0.035835f
C735 VTAIL.n297 VSUBS 0.016053f
C736 VTAIL.n298 VSUBS 0.015161f
C737 VTAIL.n299 VSUBS 0.028214f
C738 VTAIL.n300 VSUBS 0.028214f
C739 VTAIL.n301 VSUBS 0.015161f
C740 VTAIL.n302 VSUBS 0.016053f
C741 VTAIL.n303 VSUBS 0.035835f
C742 VTAIL.n304 VSUBS 0.035835f
C743 VTAIL.n305 VSUBS 0.016053f
C744 VTAIL.n306 VSUBS 0.015161f
C745 VTAIL.n307 VSUBS 0.028214f
C746 VTAIL.n308 VSUBS 0.028214f
C747 VTAIL.n309 VSUBS 0.015161f
C748 VTAIL.n310 VSUBS 0.016053f
C749 VTAIL.n311 VSUBS 0.035835f
C750 VTAIL.n312 VSUBS 0.035835f
C751 VTAIL.n313 VSUBS 0.016053f
C752 VTAIL.n314 VSUBS 0.015161f
C753 VTAIL.n315 VSUBS 0.028214f
C754 VTAIL.n316 VSUBS 0.028214f
C755 VTAIL.n317 VSUBS 0.015161f
C756 VTAIL.n318 VSUBS 0.016053f
C757 VTAIL.n319 VSUBS 0.035835f
C758 VTAIL.n320 VSUBS 0.035835f
C759 VTAIL.n321 VSUBS 0.016053f
C760 VTAIL.n322 VSUBS 0.015161f
C761 VTAIL.n323 VSUBS 0.028214f
C762 VTAIL.n324 VSUBS 0.028214f
C763 VTAIL.n325 VSUBS 0.015161f
C764 VTAIL.n326 VSUBS 0.016053f
C765 VTAIL.n327 VSUBS 0.035835f
C766 VTAIL.n328 VSUBS 0.035835f
C767 VTAIL.n329 VSUBS 0.016053f
C768 VTAIL.n330 VSUBS 0.015161f
C769 VTAIL.n331 VSUBS 0.028214f
C770 VTAIL.n332 VSUBS 0.028214f
C771 VTAIL.n333 VSUBS 0.015161f
C772 VTAIL.n334 VSUBS 0.015161f
C773 VTAIL.n335 VSUBS 0.016053f
C774 VTAIL.n336 VSUBS 0.035835f
C775 VTAIL.n337 VSUBS 0.035835f
C776 VTAIL.n338 VSUBS 0.035835f
C777 VTAIL.n339 VSUBS 0.015607f
C778 VTAIL.n340 VSUBS 0.015161f
C779 VTAIL.n341 VSUBS 0.028214f
C780 VTAIL.n342 VSUBS 0.028214f
C781 VTAIL.n343 VSUBS 0.015161f
C782 VTAIL.n344 VSUBS 0.016053f
C783 VTAIL.n345 VSUBS 0.035835f
C784 VTAIL.n346 VSUBS 0.0835f
C785 VTAIL.n347 VSUBS 0.016053f
C786 VTAIL.n348 VSUBS 0.015161f
C787 VTAIL.n349 VSUBS 0.068685f
C788 VTAIL.n350 VSUBS 0.041951f
C789 VTAIL.n351 VSUBS 2.04692f
C790 VP.t5 VSUBS 3.52753f
C791 VP.n0 VSUBS 1.33857f
C792 VP.n1 VSUBS 0.029527f
C793 VP.n2 VSUBS 0.049278f
C794 VP.n3 VSUBS 0.029527f
C795 VP.t3 VSUBS 3.52753f
C796 VP.n4 VSUBS 0.055032f
C797 VP.n5 VSUBS 0.029527f
C798 VP.n6 VSUBS 0.049598f
C799 VP.t0 VSUBS 3.52753f
C800 VP.n7 VSUBS 1.33857f
C801 VP.n8 VSUBS 0.029527f
C802 VP.n9 VSUBS 0.049278f
C803 VP.n10 VSUBS 0.313309f
C804 VP.t4 VSUBS 3.52753f
C805 VP.t1 VSUBS 3.8019f
C806 VP.n11 VSUBS 1.28522f
C807 VP.n12 VSUBS 1.31964f
C808 VP.n13 VSUBS 0.041447f
C809 VP.n14 VSUBS 0.055032f
C810 VP.n15 VSUBS 0.029527f
C811 VP.n16 VSUBS 0.029527f
C812 VP.n17 VSUBS 0.029527f
C813 VP.n18 VSUBS 0.036936f
C814 VP.n19 VSUBS 0.055032f
C815 VP.n20 VSUBS 0.049598f
C816 VP.n21 VSUBS 0.047657f
C817 VP.n22 VSUBS 1.77306f
C818 VP.t2 VSUBS 3.52753f
C819 VP.n23 VSUBS 1.33857f
C820 VP.n24 VSUBS 1.79339f
C821 VP.n25 VSUBS 0.047657f
C822 VP.n26 VSUBS 0.029527f
C823 VP.n27 VSUBS 0.055032f
C824 VP.n28 VSUBS 0.036936f
C825 VP.n29 VSUBS 0.049278f
C826 VP.n30 VSUBS 0.029527f
C827 VP.n31 VSUBS 0.029527f
C828 VP.n32 VSUBS 0.029527f
C829 VP.n33 VSUBS 0.041447f
C830 VP.n34 VSUBS 1.22894f
C831 VP.n35 VSUBS 0.041447f
C832 VP.n36 VSUBS 0.055032f
C833 VP.n37 VSUBS 0.029527f
C834 VP.n38 VSUBS 0.029527f
C835 VP.n39 VSUBS 0.029527f
C836 VP.n40 VSUBS 0.036936f
C837 VP.n41 VSUBS 0.055032f
C838 VP.n42 VSUBS 0.049598f
C839 VP.n43 VSUBS 0.047657f
C840 VP.n44 VSUBS 0.060233f
C841 B.n0 VSUBS 0.005089f
C842 B.n1 VSUBS 0.005089f
C843 B.n2 VSUBS 0.008048f
C844 B.n3 VSUBS 0.008048f
C845 B.n4 VSUBS 0.008048f
C846 B.n5 VSUBS 0.008048f
C847 B.n6 VSUBS 0.008048f
C848 B.n7 VSUBS 0.008048f
C849 B.n8 VSUBS 0.008048f
C850 B.n9 VSUBS 0.008048f
C851 B.n10 VSUBS 0.008048f
C852 B.n11 VSUBS 0.008048f
C853 B.n12 VSUBS 0.008048f
C854 B.n13 VSUBS 0.008048f
C855 B.n14 VSUBS 0.008048f
C856 B.n15 VSUBS 0.008048f
C857 B.n16 VSUBS 0.008048f
C858 B.n17 VSUBS 0.008048f
C859 B.n18 VSUBS 0.008048f
C860 B.n19 VSUBS 0.008048f
C861 B.n20 VSUBS 0.008048f
C862 B.n21 VSUBS 0.008048f
C863 B.n22 VSUBS 0.008048f
C864 B.n23 VSUBS 0.008048f
C865 B.n24 VSUBS 0.019136f
C866 B.n25 VSUBS 0.008048f
C867 B.n26 VSUBS 0.008048f
C868 B.n27 VSUBS 0.008048f
C869 B.n28 VSUBS 0.008048f
C870 B.n29 VSUBS 0.008048f
C871 B.n30 VSUBS 0.008048f
C872 B.n31 VSUBS 0.008048f
C873 B.n32 VSUBS 0.008048f
C874 B.n33 VSUBS 0.008048f
C875 B.n34 VSUBS 0.008048f
C876 B.n35 VSUBS 0.008048f
C877 B.n36 VSUBS 0.008048f
C878 B.n37 VSUBS 0.008048f
C879 B.n38 VSUBS 0.008048f
C880 B.n39 VSUBS 0.008048f
C881 B.n40 VSUBS 0.008048f
C882 B.n41 VSUBS 0.008048f
C883 B.n42 VSUBS 0.008048f
C884 B.n43 VSUBS 0.008048f
C885 B.n44 VSUBS 0.008048f
C886 B.n45 VSUBS 0.008048f
C887 B.n46 VSUBS 0.008048f
C888 B.n47 VSUBS 0.008048f
C889 B.n48 VSUBS 0.008048f
C890 B.n49 VSUBS 0.008048f
C891 B.n50 VSUBS 0.005563f
C892 B.n51 VSUBS 0.008048f
C893 B.t8 VSUBS 0.3336f
C894 B.t7 VSUBS 0.374205f
C895 B.t6 VSUBS 2.25807f
C896 B.n52 VSUBS 0.584627f
C897 B.n53 VSUBS 0.343033f
C898 B.n54 VSUBS 0.018647f
C899 B.n55 VSUBS 0.008048f
C900 B.n56 VSUBS 0.008048f
C901 B.n57 VSUBS 0.008048f
C902 B.n58 VSUBS 0.008048f
C903 B.t2 VSUBS 0.333604f
C904 B.t1 VSUBS 0.374208f
C905 B.t0 VSUBS 2.25807f
C906 B.n59 VSUBS 0.584624f
C907 B.n60 VSUBS 0.343029f
C908 B.n61 VSUBS 0.008048f
C909 B.n62 VSUBS 0.008048f
C910 B.n63 VSUBS 0.008048f
C911 B.n64 VSUBS 0.008048f
C912 B.n65 VSUBS 0.008048f
C913 B.n66 VSUBS 0.008048f
C914 B.n67 VSUBS 0.008048f
C915 B.n68 VSUBS 0.008048f
C916 B.n69 VSUBS 0.008048f
C917 B.n70 VSUBS 0.008048f
C918 B.n71 VSUBS 0.008048f
C919 B.n72 VSUBS 0.008048f
C920 B.n73 VSUBS 0.008048f
C921 B.n74 VSUBS 0.008048f
C922 B.n75 VSUBS 0.008048f
C923 B.n76 VSUBS 0.008048f
C924 B.n77 VSUBS 0.008048f
C925 B.n78 VSUBS 0.008048f
C926 B.n79 VSUBS 0.008048f
C927 B.n80 VSUBS 0.008048f
C928 B.n81 VSUBS 0.008048f
C929 B.n82 VSUBS 0.008048f
C930 B.n83 VSUBS 0.008048f
C931 B.n84 VSUBS 0.008048f
C932 B.n85 VSUBS 0.008048f
C933 B.n86 VSUBS 0.019136f
C934 B.n87 VSUBS 0.008048f
C935 B.n88 VSUBS 0.008048f
C936 B.n89 VSUBS 0.008048f
C937 B.n90 VSUBS 0.008048f
C938 B.n91 VSUBS 0.008048f
C939 B.n92 VSUBS 0.008048f
C940 B.n93 VSUBS 0.008048f
C941 B.n94 VSUBS 0.008048f
C942 B.n95 VSUBS 0.008048f
C943 B.n96 VSUBS 0.008048f
C944 B.n97 VSUBS 0.008048f
C945 B.n98 VSUBS 0.008048f
C946 B.n99 VSUBS 0.008048f
C947 B.n100 VSUBS 0.008048f
C948 B.n101 VSUBS 0.008048f
C949 B.n102 VSUBS 0.008048f
C950 B.n103 VSUBS 0.008048f
C951 B.n104 VSUBS 0.008048f
C952 B.n105 VSUBS 0.008048f
C953 B.n106 VSUBS 0.008048f
C954 B.n107 VSUBS 0.008048f
C955 B.n108 VSUBS 0.008048f
C956 B.n109 VSUBS 0.008048f
C957 B.n110 VSUBS 0.008048f
C958 B.n111 VSUBS 0.008048f
C959 B.n112 VSUBS 0.008048f
C960 B.n113 VSUBS 0.008048f
C961 B.n114 VSUBS 0.008048f
C962 B.n115 VSUBS 0.008048f
C963 B.n116 VSUBS 0.008048f
C964 B.n117 VSUBS 0.008048f
C965 B.n118 VSUBS 0.008048f
C966 B.n119 VSUBS 0.008048f
C967 B.n120 VSUBS 0.008048f
C968 B.n121 VSUBS 0.008048f
C969 B.n122 VSUBS 0.008048f
C970 B.n123 VSUBS 0.008048f
C971 B.n124 VSUBS 0.008048f
C972 B.n125 VSUBS 0.008048f
C973 B.n126 VSUBS 0.008048f
C974 B.n127 VSUBS 0.008048f
C975 B.n128 VSUBS 0.008048f
C976 B.n129 VSUBS 0.008048f
C977 B.n130 VSUBS 0.008048f
C978 B.n131 VSUBS 0.019136f
C979 B.n132 VSUBS 0.008048f
C980 B.n133 VSUBS 0.008048f
C981 B.n134 VSUBS 0.008048f
C982 B.n135 VSUBS 0.008048f
C983 B.n136 VSUBS 0.008048f
C984 B.n137 VSUBS 0.008048f
C985 B.n138 VSUBS 0.008048f
C986 B.n139 VSUBS 0.008048f
C987 B.n140 VSUBS 0.008048f
C988 B.n141 VSUBS 0.008048f
C989 B.n142 VSUBS 0.008048f
C990 B.n143 VSUBS 0.008048f
C991 B.n144 VSUBS 0.008048f
C992 B.n145 VSUBS 0.008048f
C993 B.n146 VSUBS 0.008048f
C994 B.n147 VSUBS 0.008048f
C995 B.n148 VSUBS 0.008048f
C996 B.n149 VSUBS 0.008048f
C997 B.n150 VSUBS 0.008048f
C998 B.n151 VSUBS 0.008048f
C999 B.n152 VSUBS 0.008048f
C1000 B.n153 VSUBS 0.008048f
C1001 B.n154 VSUBS 0.008048f
C1002 B.n155 VSUBS 0.008048f
C1003 B.n156 VSUBS 0.008048f
C1004 B.n157 VSUBS 0.005563f
C1005 B.n158 VSUBS 0.008048f
C1006 B.n159 VSUBS 0.008048f
C1007 B.n160 VSUBS 0.008048f
C1008 B.n161 VSUBS 0.008048f
C1009 B.n162 VSUBS 0.008048f
C1010 B.t4 VSUBS 0.3336f
C1011 B.t5 VSUBS 0.374205f
C1012 B.t3 VSUBS 2.25807f
C1013 B.n163 VSUBS 0.584627f
C1014 B.n164 VSUBS 0.343033f
C1015 B.n165 VSUBS 0.008048f
C1016 B.n166 VSUBS 0.008048f
C1017 B.n167 VSUBS 0.008048f
C1018 B.n168 VSUBS 0.008048f
C1019 B.n169 VSUBS 0.008048f
C1020 B.n170 VSUBS 0.008048f
C1021 B.n171 VSUBS 0.008048f
C1022 B.n172 VSUBS 0.008048f
C1023 B.n173 VSUBS 0.008048f
C1024 B.n174 VSUBS 0.008048f
C1025 B.n175 VSUBS 0.008048f
C1026 B.n176 VSUBS 0.008048f
C1027 B.n177 VSUBS 0.008048f
C1028 B.n178 VSUBS 0.008048f
C1029 B.n179 VSUBS 0.008048f
C1030 B.n180 VSUBS 0.008048f
C1031 B.n181 VSUBS 0.008048f
C1032 B.n182 VSUBS 0.008048f
C1033 B.n183 VSUBS 0.008048f
C1034 B.n184 VSUBS 0.008048f
C1035 B.n185 VSUBS 0.008048f
C1036 B.n186 VSUBS 0.008048f
C1037 B.n187 VSUBS 0.008048f
C1038 B.n188 VSUBS 0.008048f
C1039 B.n189 VSUBS 0.008048f
C1040 B.n190 VSUBS 0.019136f
C1041 B.n191 VSUBS 0.008048f
C1042 B.n192 VSUBS 0.008048f
C1043 B.n193 VSUBS 0.008048f
C1044 B.n194 VSUBS 0.008048f
C1045 B.n195 VSUBS 0.008048f
C1046 B.n196 VSUBS 0.008048f
C1047 B.n197 VSUBS 0.008048f
C1048 B.n198 VSUBS 0.008048f
C1049 B.n199 VSUBS 0.008048f
C1050 B.n200 VSUBS 0.008048f
C1051 B.n201 VSUBS 0.008048f
C1052 B.n202 VSUBS 0.008048f
C1053 B.n203 VSUBS 0.008048f
C1054 B.n204 VSUBS 0.008048f
C1055 B.n205 VSUBS 0.008048f
C1056 B.n206 VSUBS 0.008048f
C1057 B.n207 VSUBS 0.008048f
C1058 B.n208 VSUBS 0.008048f
C1059 B.n209 VSUBS 0.008048f
C1060 B.n210 VSUBS 0.008048f
C1061 B.n211 VSUBS 0.008048f
C1062 B.n212 VSUBS 0.008048f
C1063 B.n213 VSUBS 0.008048f
C1064 B.n214 VSUBS 0.008048f
C1065 B.n215 VSUBS 0.008048f
C1066 B.n216 VSUBS 0.008048f
C1067 B.n217 VSUBS 0.008048f
C1068 B.n218 VSUBS 0.008048f
C1069 B.n219 VSUBS 0.008048f
C1070 B.n220 VSUBS 0.008048f
C1071 B.n221 VSUBS 0.008048f
C1072 B.n222 VSUBS 0.008048f
C1073 B.n223 VSUBS 0.008048f
C1074 B.n224 VSUBS 0.008048f
C1075 B.n225 VSUBS 0.008048f
C1076 B.n226 VSUBS 0.008048f
C1077 B.n227 VSUBS 0.008048f
C1078 B.n228 VSUBS 0.008048f
C1079 B.n229 VSUBS 0.008048f
C1080 B.n230 VSUBS 0.008048f
C1081 B.n231 VSUBS 0.008048f
C1082 B.n232 VSUBS 0.008048f
C1083 B.n233 VSUBS 0.008048f
C1084 B.n234 VSUBS 0.008048f
C1085 B.n235 VSUBS 0.008048f
C1086 B.n236 VSUBS 0.008048f
C1087 B.n237 VSUBS 0.008048f
C1088 B.n238 VSUBS 0.008048f
C1089 B.n239 VSUBS 0.008048f
C1090 B.n240 VSUBS 0.008048f
C1091 B.n241 VSUBS 0.008048f
C1092 B.n242 VSUBS 0.008048f
C1093 B.n243 VSUBS 0.008048f
C1094 B.n244 VSUBS 0.008048f
C1095 B.n245 VSUBS 0.008048f
C1096 B.n246 VSUBS 0.008048f
C1097 B.n247 VSUBS 0.008048f
C1098 B.n248 VSUBS 0.008048f
C1099 B.n249 VSUBS 0.008048f
C1100 B.n250 VSUBS 0.008048f
C1101 B.n251 VSUBS 0.008048f
C1102 B.n252 VSUBS 0.008048f
C1103 B.n253 VSUBS 0.008048f
C1104 B.n254 VSUBS 0.008048f
C1105 B.n255 VSUBS 0.008048f
C1106 B.n256 VSUBS 0.008048f
C1107 B.n257 VSUBS 0.008048f
C1108 B.n258 VSUBS 0.008048f
C1109 B.n259 VSUBS 0.008048f
C1110 B.n260 VSUBS 0.008048f
C1111 B.n261 VSUBS 0.008048f
C1112 B.n262 VSUBS 0.008048f
C1113 B.n263 VSUBS 0.008048f
C1114 B.n264 VSUBS 0.008048f
C1115 B.n265 VSUBS 0.008048f
C1116 B.n266 VSUBS 0.008048f
C1117 B.n267 VSUBS 0.008048f
C1118 B.n268 VSUBS 0.008048f
C1119 B.n269 VSUBS 0.008048f
C1120 B.n270 VSUBS 0.008048f
C1121 B.n271 VSUBS 0.008048f
C1122 B.n272 VSUBS 0.008048f
C1123 B.n273 VSUBS 0.008048f
C1124 B.n274 VSUBS 0.008048f
C1125 B.n275 VSUBS 0.008048f
C1126 B.n276 VSUBS 0.008048f
C1127 B.n277 VSUBS 0.019136f
C1128 B.n278 VSUBS 0.020159f
C1129 B.n279 VSUBS 0.020159f
C1130 B.n280 VSUBS 0.008048f
C1131 B.n281 VSUBS 0.008048f
C1132 B.n282 VSUBS 0.008048f
C1133 B.n283 VSUBS 0.008048f
C1134 B.n284 VSUBS 0.008048f
C1135 B.n285 VSUBS 0.008048f
C1136 B.n286 VSUBS 0.008048f
C1137 B.n287 VSUBS 0.008048f
C1138 B.n288 VSUBS 0.008048f
C1139 B.n289 VSUBS 0.008048f
C1140 B.n290 VSUBS 0.008048f
C1141 B.n291 VSUBS 0.008048f
C1142 B.n292 VSUBS 0.008048f
C1143 B.n293 VSUBS 0.008048f
C1144 B.n294 VSUBS 0.008048f
C1145 B.n295 VSUBS 0.008048f
C1146 B.n296 VSUBS 0.008048f
C1147 B.n297 VSUBS 0.008048f
C1148 B.n298 VSUBS 0.008048f
C1149 B.n299 VSUBS 0.008048f
C1150 B.n300 VSUBS 0.008048f
C1151 B.n301 VSUBS 0.008048f
C1152 B.n302 VSUBS 0.008048f
C1153 B.n303 VSUBS 0.008048f
C1154 B.n304 VSUBS 0.008048f
C1155 B.n305 VSUBS 0.008048f
C1156 B.n306 VSUBS 0.008048f
C1157 B.n307 VSUBS 0.008048f
C1158 B.n308 VSUBS 0.008048f
C1159 B.n309 VSUBS 0.008048f
C1160 B.n310 VSUBS 0.008048f
C1161 B.n311 VSUBS 0.008048f
C1162 B.n312 VSUBS 0.008048f
C1163 B.n313 VSUBS 0.008048f
C1164 B.n314 VSUBS 0.008048f
C1165 B.n315 VSUBS 0.008048f
C1166 B.n316 VSUBS 0.008048f
C1167 B.n317 VSUBS 0.008048f
C1168 B.n318 VSUBS 0.008048f
C1169 B.n319 VSUBS 0.008048f
C1170 B.n320 VSUBS 0.008048f
C1171 B.n321 VSUBS 0.008048f
C1172 B.n322 VSUBS 0.008048f
C1173 B.n323 VSUBS 0.008048f
C1174 B.n324 VSUBS 0.008048f
C1175 B.n325 VSUBS 0.008048f
C1176 B.n326 VSUBS 0.008048f
C1177 B.n327 VSUBS 0.008048f
C1178 B.n328 VSUBS 0.008048f
C1179 B.n329 VSUBS 0.008048f
C1180 B.n330 VSUBS 0.008048f
C1181 B.n331 VSUBS 0.008048f
C1182 B.n332 VSUBS 0.008048f
C1183 B.n333 VSUBS 0.008048f
C1184 B.n334 VSUBS 0.008048f
C1185 B.n335 VSUBS 0.008048f
C1186 B.n336 VSUBS 0.008048f
C1187 B.n337 VSUBS 0.008048f
C1188 B.n338 VSUBS 0.008048f
C1189 B.n339 VSUBS 0.008048f
C1190 B.n340 VSUBS 0.008048f
C1191 B.n341 VSUBS 0.008048f
C1192 B.n342 VSUBS 0.008048f
C1193 B.n343 VSUBS 0.008048f
C1194 B.n344 VSUBS 0.008048f
C1195 B.n345 VSUBS 0.008048f
C1196 B.n346 VSUBS 0.008048f
C1197 B.n347 VSUBS 0.008048f
C1198 B.n348 VSUBS 0.008048f
C1199 B.n349 VSUBS 0.008048f
C1200 B.n350 VSUBS 0.008048f
C1201 B.n351 VSUBS 0.008048f
C1202 B.n352 VSUBS 0.008048f
C1203 B.n353 VSUBS 0.008048f
C1204 B.n354 VSUBS 0.008048f
C1205 B.n355 VSUBS 0.005563f
C1206 B.n356 VSUBS 0.018647f
C1207 B.n357 VSUBS 0.00651f
C1208 B.n358 VSUBS 0.008048f
C1209 B.n359 VSUBS 0.008048f
C1210 B.n360 VSUBS 0.008048f
C1211 B.n361 VSUBS 0.008048f
C1212 B.n362 VSUBS 0.008048f
C1213 B.n363 VSUBS 0.008048f
C1214 B.n364 VSUBS 0.008048f
C1215 B.n365 VSUBS 0.008048f
C1216 B.n366 VSUBS 0.008048f
C1217 B.n367 VSUBS 0.008048f
C1218 B.n368 VSUBS 0.008048f
C1219 B.t10 VSUBS 0.333604f
C1220 B.t11 VSUBS 0.374208f
C1221 B.t9 VSUBS 2.25807f
C1222 B.n369 VSUBS 0.584624f
C1223 B.n370 VSUBS 0.343029f
C1224 B.n371 VSUBS 0.018647f
C1225 B.n372 VSUBS 0.00651f
C1226 B.n373 VSUBS 0.008048f
C1227 B.n374 VSUBS 0.008048f
C1228 B.n375 VSUBS 0.008048f
C1229 B.n376 VSUBS 0.008048f
C1230 B.n377 VSUBS 0.008048f
C1231 B.n378 VSUBS 0.008048f
C1232 B.n379 VSUBS 0.008048f
C1233 B.n380 VSUBS 0.008048f
C1234 B.n381 VSUBS 0.008048f
C1235 B.n382 VSUBS 0.008048f
C1236 B.n383 VSUBS 0.008048f
C1237 B.n384 VSUBS 0.008048f
C1238 B.n385 VSUBS 0.008048f
C1239 B.n386 VSUBS 0.008048f
C1240 B.n387 VSUBS 0.008048f
C1241 B.n388 VSUBS 0.008048f
C1242 B.n389 VSUBS 0.008048f
C1243 B.n390 VSUBS 0.008048f
C1244 B.n391 VSUBS 0.008048f
C1245 B.n392 VSUBS 0.008048f
C1246 B.n393 VSUBS 0.008048f
C1247 B.n394 VSUBS 0.008048f
C1248 B.n395 VSUBS 0.008048f
C1249 B.n396 VSUBS 0.008048f
C1250 B.n397 VSUBS 0.008048f
C1251 B.n398 VSUBS 0.008048f
C1252 B.n399 VSUBS 0.008048f
C1253 B.n400 VSUBS 0.008048f
C1254 B.n401 VSUBS 0.008048f
C1255 B.n402 VSUBS 0.008048f
C1256 B.n403 VSUBS 0.008048f
C1257 B.n404 VSUBS 0.008048f
C1258 B.n405 VSUBS 0.008048f
C1259 B.n406 VSUBS 0.008048f
C1260 B.n407 VSUBS 0.008048f
C1261 B.n408 VSUBS 0.008048f
C1262 B.n409 VSUBS 0.008048f
C1263 B.n410 VSUBS 0.008048f
C1264 B.n411 VSUBS 0.008048f
C1265 B.n412 VSUBS 0.008048f
C1266 B.n413 VSUBS 0.008048f
C1267 B.n414 VSUBS 0.008048f
C1268 B.n415 VSUBS 0.008048f
C1269 B.n416 VSUBS 0.008048f
C1270 B.n417 VSUBS 0.008048f
C1271 B.n418 VSUBS 0.008048f
C1272 B.n419 VSUBS 0.008048f
C1273 B.n420 VSUBS 0.008048f
C1274 B.n421 VSUBS 0.008048f
C1275 B.n422 VSUBS 0.008048f
C1276 B.n423 VSUBS 0.008048f
C1277 B.n424 VSUBS 0.008048f
C1278 B.n425 VSUBS 0.008048f
C1279 B.n426 VSUBS 0.008048f
C1280 B.n427 VSUBS 0.008048f
C1281 B.n428 VSUBS 0.008048f
C1282 B.n429 VSUBS 0.008048f
C1283 B.n430 VSUBS 0.008048f
C1284 B.n431 VSUBS 0.008048f
C1285 B.n432 VSUBS 0.008048f
C1286 B.n433 VSUBS 0.008048f
C1287 B.n434 VSUBS 0.008048f
C1288 B.n435 VSUBS 0.008048f
C1289 B.n436 VSUBS 0.008048f
C1290 B.n437 VSUBS 0.008048f
C1291 B.n438 VSUBS 0.008048f
C1292 B.n439 VSUBS 0.008048f
C1293 B.n440 VSUBS 0.008048f
C1294 B.n441 VSUBS 0.008048f
C1295 B.n442 VSUBS 0.008048f
C1296 B.n443 VSUBS 0.008048f
C1297 B.n444 VSUBS 0.008048f
C1298 B.n445 VSUBS 0.008048f
C1299 B.n446 VSUBS 0.008048f
C1300 B.n447 VSUBS 0.008048f
C1301 B.n448 VSUBS 0.008048f
C1302 B.n449 VSUBS 0.008048f
C1303 B.n450 VSUBS 0.020159f
C1304 B.n451 VSUBS 0.020159f
C1305 B.n452 VSUBS 0.019136f
C1306 B.n453 VSUBS 0.008048f
C1307 B.n454 VSUBS 0.008048f
C1308 B.n455 VSUBS 0.008048f
C1309 B.n456 VSUBS 0.008048f
C1310 B.n457 VSUBS 0.008048f
C1311 B.n458 VSUBS 0.008048f
C1312 B.n459 VSUBS 0.008048f
C1313 B.n460 VSUBS 0.008048f
C1314 B.n461 VSUBS 0.008048f
C1315 B.n462 VSUBS 0.008048f
C1316 B.n463 VSUBS 0.008048f
C1317 B.n464 VSUBS 0.008048f
C1318 B.n465 VSUBS 0.008048f
C1319 B.n466 VSUBS 0.008048f
C1320 B.n467 VSUBS 0.008048f
C1321 B.n468 VSUBS 0.008048f
C1322 B.n469 VSUBS 0.008048f
C1323 B.n470 VSUBS 0.008048f
C1324 B.n471 VSUBS 0.008048f
C1325 B.n472 VSUBS 0.008048f
C1326 B.n473 VSUBS 0.008048f
C1327 B.n474 VSUBS 0.008048f
C1328 B.n475 VSUBS 0.008048f
C1329 B.n476 VSUBS 0.008048f
C1330 B.n477 VSUBS 0.008048f
C1331 B.n478 VSUBS 0.008048f
C1332 B.n479 VSUBS 0.008048f
C1333 B.n480 VSUBS 0.008048f
C1334 B.n481 VSUBS 0.008048f
C1335 B.n482 VSUBS 0.008048f
C1336 B.n483 VSUBS 0.008048f
C1337 B.n484 VSUBS 0.008048f
C1338 B.n485 VSUBS 0.008048f
C1339 B.n486 VSUBS 0.008048f
C1340 B.n487 VSUBS 0.008048f
C1341 B.n488 VSUBS 0.008048f
C1342 B.n489 VSUBS 0.008048f
C1343 B.n490 VSUBS 0.008048f
C1344 B.n491 VSUBS 0.008048f
C1345 B.n492 VSUBS 0.008048f
C1346 B.n493 VSUBS 0.008048f
C1347 B.n494 VSUBS 0.008048f
C1348 B.n495 VSUBS 0.008048f
C1349 B.n496 VSUBS 0.008048f
C1350 B.n497 VSUBS 0.008048f
C1351 B.n498 VSUBS 0.008048f
C1352 B.n499 VSUBS 0.008048f
C1353 B.n500 VSUBS 0.008048f
C1354 B.n501 VSUBS 0.008048f
C1355 B.n502 VSUBS 0.008048f
C1356 B.n503 VSUBS 0.008048f
C1357 B.n504 VSUBS 0.008048f
C1358 B.n505 VSUBS 0.008048f
C1359 B.n506 VSUBS 0.008048f
C1360 B.n507 VSUBS 0.008048f
C1361 B.n508 VSUBS 0.008048f
C1362 B.n509 VSUBS 0.008048f
C1363 B.n510 VSUBS 0.008048f
C1364 B.n511 VSUBS 0.008048f
C1365 B.n512 VSUBS 0.008048f
C1366 B.n513 VSUBS 0.008048f
C1367 B.n514 VSUBS 0.008048f
C1368 B.n515 VSUBS 0.008048f
C1369 B.n516 VSUBS 0.008048f
C1370 B.n517 VSUBS 0.008048f
C1371 B.n518 VSUBS 0.008048f
C1372 B.n519 VSUBS 0.008048f
C1373 B.n520 VSUBS 0.008048f
C1374 B.n521 VSUBS 0.008048f
C1375 B.n522 VSUBS 0.008048f
C1376 B.n523 VSUBS 0.008048f
C1377 B.n524 VSUBS 0.008048f
C1378 B.n525 VSUBS 0.008048f
C1379 B.n526 VSUBS 0.008048f
C1380 B.n527 VSUBS 0.008048f
C1381 B.n528 VSUBS 0.008048f
C1382 B.n529 VSUBS 0.008048f
C1383 B.n530 VSUBS 0.008048f
C1384 B.n531 VSUBS 0.008048f
C1385 B.n532 VSUBS 0.008048f
C1386 B.n533 VSUBS 0.008048f
C1387 B.n534 VSUBS 0.008048f
C1388 B.n535 VSUBS 0.008048f
C1389 B.n536 VSUBS 0.008048f
C1390 B.n537 VSUBS 0.008048f
C1391 B.n538 VSUBS 0.008048f
C1392 B.n539 VSUBS 0.008048f
C1393 B.n540 VSUBS 0.008048f
C1394 B.n541 VSUBS 0.008048f
C1395 B.n542 VSUBS 0.008048f
C1396 B.n543 VSUBS 0.008048f
C1397 B.n544 VSUBS 0.008048f
C1398 B.n545 VSUBS 0.008048f
C1399 B.n546 VSUBS 0.008048f
C1400 B.n547 VSUBS 0.008048f
C1401 B.n548 VSUBS 0.008048f
C1402 B.n549 VSUBS 0.008048f
C1403 B.n550 VSUBS 0.008048f
C1404 B.n551 VSUBS 0.008048f
C1405 B.n552 VSUBS 0.008048f
C1406 B.n553 VSUBS 0.008048f
C1407 B.n554 VSUBS 0.008048f
C1408 B.n555 VSUBS 0.008048f
C1409 B.n556 VSUBS 0.008048f
C1410 B.n557 VSUBS 0.008048f
C1411 B.n558 VSUBS 0.008048f
C1412 B.n559 VSUBS 0.008048f
C1413 B.n560 VSUBS 0.008048f
C1414 B.n561 VSUBS 0.008048f
C1415 B.n562 VSUBS 0.008048f
C1416 B.n563 VSUBS 0.008048f
C1417 B.n564 VSUBS 0.008048f
C1418 B.n565 VSUBS 0.008048f
C1419 B.n566 VSUBS 0.008048f
C1420 B.n567 VSUBS 0.008048f
C1421 B.n568 VSUBS 0.008048f
C1422 B.n569 VSUBS 0.008048f
C1423 B.n570 VSUBS 0.008048f
C1424 B.n571 VSUBS 0.008048f
C1425 B.n572 VSUBS 0.008048f
C1426 B.n573 VSUBS 0.008048f
C1427 B.n574 VSUBS 0.008048f
C1428 B.n575 VSUBS 0.008048f
C1429 B.n576 VSUBS 0.008048f
C1430 B.n577 VSUBS 0.008048f
C1431 B.n578 VSUBS 0.008048f
C1432 B.n579 VSUBS 0.008048f
C1433 B.n580 VSUBS 0.008048f
C1434 B.n581 VSUBS 0.008048f
C1435 B.n582 VSUBS 0.008048f
C1436 B.n583 VSUBS 0.008048f
C1437 B.n584 VSUBS 0.008048f
C1438 B.n585 VSUBS 0.008048f
C1439 B.n586 VSUBS 0.008048f
C1440 B.n587 VSUBS 0.020028f
C1441 B.n588 VSUBS 0.019266f
C1442 B.n589 VSUBS 0.020159f
C1443 B.n590 VSUBS 0.008048f
C1444 B.n591 VSUBS 0.008048f
C1445 B.n592 VSUBS 0.008048f
C1446 B.n593 VSUBS 0.008048f
C1447 B.n594 VSUBS 0.008048f
C1448 B.n595 VSUBS 0.008048f
C1449 B.n596 VSUBS 0.008048f
C1450 B.n597 VSUBS 0.008048f
C1451 B.n598 VSUBS 0.008048f
C1452 B.n599 VSUBS 0.008048f
C1453 B.n600 VSUBS 0.008048f
C1454 B.n601 VSUBS 0.008048f
C1455 B.n602 VSUBS 0.008048f
C1456 B.n603 VSUBS 0.008048f
C1457 B.n604 VSUBS 0.008048f
C1458 B.n605 VSUBS 0.008048f
C1459 B.n606 VSUBS 0.008048f
C1460 B.n607 VSUBS 0.008048f
C1461 B.n608 VSUBS 0.008048f
C1462 B.n609 VSUBS 0.008048f
C1463 B.n610 VSUBS 0.008048f
C1464 B.n611 VSUBS 0.008048f
C1465 B.n612 VSUBS 0.008048f
C1466 B.n613 VSUBS 0.008048f
C1467 B.n614 VSUBS 0.008048f
C1468 B.n615 VSUBS 0.008048f
C1469 B.n616 VSUBS 0.008048f
C1470 B.n617 VSUBS 0.008048f
C1471 B.n618 VSUBS 0.008048f
C1472 B.n619 VSUBS 0.008048f
C1473 B.n620 VSUBS 0.008048f
C1474 B.n621 VSUBS 0.008048f
C1475 B.n622 VSUBS 0.008048f
C1476 B.n623 VSUBS 0.008048f
C1477 B.n624 VSUBS 0.008048f
C1478 B.n625 VSUBS 0.008048f
C1479 B.n626 VSUBS 0.008048f
C1480 B.n627 VSUBS 0.008048f
C1481 B.n628 VSUBS 0.008048f
C1482 B.n629 VSUBS 0.008048f
C1483 B.n630 VSUBS 0.008048f
C1484 B.n631 VSUBS 0.008048f
C1485 B.n632 VSUBS 0.008048f
C1486 B.n633 VSUBS 0.008048f
C1487 B.n634 VSUBS 0.008048f
C1488 B.n635 VSUBS 0.008048f
C1489 B.n636 VSUBS 0.008048f
C1490 B.n637 VSUBS 0.008048f
C1491 B.n638 VSUBS 0.008048f
C1492 B.n639 VSUBS 0.008048f
C1493 B.n640 VSUBS 0.008048f
C1494 B.n641 VSUBS 0.008048f
C1495 B.n642 VSUBS 0.008048f
C1496 B.n643 VSUBS 0.008048f
C1497 B.n644 VSUBS 0.008048f
C1498 B.n645 VSUBS 0.008048f
C1499 B.n646 VSUBS 0.008048f
C1500 B.n647 VSUBS 0.008048f
C1501 B.n648 VSUBS 0.008048f
C1502 B.n649 VSUBS 0.008048f
C1503 B.n650 VSUBS 0.008048f
C1504 B.n651 VSUBS 0.008048f
C1505 B.n652 VSUBS 0.008048f
C1506 B.n653 VSUBS 0.008048f
C1507 B.n654 VSUBS 0.008048f
C1508 B.n655 VSUBS 0.008048f
C1509 B.n656 VSUBS 0.008048f
C1510 B.n657 VSUBS 0.008048f
C1511 B.n658 VSUBS 0.008048f
C1512 B.n659 VSUBS 0.008048f
C1513 B.n660 VSUBS 0.008048f
C1514 B.n661 VSUBS 0.008048f
C1515 B.n662 VSUBS 0.008048f
C1516 B.n663 VSUBS 0.008048f
C1517 B.n664 VSUBS 0.008048f
C1518 B.n665 VSUBS 0.005563f
C1519 B.n666 VSUBS 0.018647f
C1520 B.n667 VSUBS 0.00651f
C1521 B.n668 VSUBS 0.008048f
C1522 B.n669 VSUBS 0.008048f
C1523 B.n670 VSUBS 0.008048f
C1524 B.n671 VSUBS 0.008048f
C1525 B.n672 VSUBS 0.008048f
C1526 B.n673 VSUBS 0.008048f
C1527 B.n674 VSUBS 0.008048f
C1528 B.n675 VSUBS 0.008048f
C1529 B.n676 VSUBS 0.008048f
C1530 B.n677 VSUBS 0.008048f
C1531 B.n678 VSUBS 0.008048f
C1532 B.n679 VSUBS 0.00651f
C1533 B.n680 VSUBS 0.008048f
C1534 B.n681 VSUBS 0.008048f
C1535 B.n682 VSUBS 0.008048f
C1536 B.n683 VSUBS 0.008048f
C1537 B.n684 VSUBS 0.008048f
C1538 B.n685 VSUBS 0.008048f
C1539 B.n686 VSUBS 0.008048f
C1540 B.n687 VSUBS 0.008048f
C1541 B.n688 VSUBS 0.008048f
C1542 B.n689 VSUBS 0.008048f
C1543 B.n690 VSUBS 0.008048f
C1544 B.n691 VSUBS 0.008048f
C1545 B.n692 VSUBS 0.008048f
C1546 B.n693 VSUBS 0.008048f
C1547 B.n694 VSUBS 0.008048f
C1548 B.n695 VSUBS 0.008048f
C1549 B.n696 VSUBS 0.008048f
C1550 B.n697 VSUBS 0.008048f
C1551 B.n698 VSUBS 0.008048f
C1552 B.n699 VSUBS 0.008048f
C1553 B.n700 VSUBS 0.008048f
C1554 B.n701 VSUBS 0.008048f
C1555 B.n702 VSUBS 0.008048f
C1556 B.n703 VSUBS 0.008048f
C1557 B.n704 VSUBS 0.008048f
C1558 B.n705 VSUBS 0.008048f
C1559 B.n706 VSUBS 0.008048f
C1560 B.n707 VSUBS 0.008048f
C1561 B.n708 VSUBS 0.008048f
C1562 B.n709 VSUBS 0.008048f
C1563 B.n710 VSUBS 0.008048f
C1564 B.n711 VSUBS 0.008048f
C1565 B.n712 VSUBS 0.008048f
C1566 B.n713 VSUBS 0.008048f
C1567 B.n714 VSUBS 0.008048f
C1568 B.n715 VSUBS 0.008048f
C1569 B.n716 VSUBS 0.008048f
C1570 B.n717 VSUBS 0.008048f
C1571 B.n718 VSUBS 0.008048f
C1572 B.n719 VSUBS 0.008048f
C1573 B.n720 VSUBS 0.008048f
C1574 B.n721 VSUBS 0.008048f
C1575 B.n722 VSUBS 0.008048f
C1576 B.n723 VSUBS 0.008048f
C1577 B.n724 VSUBS 0.008048f
C1578 B.n725 VSUBS 0.008048f
C1579 B.n726 VSUBS 0.008048f
C1580 B.n727 VSUBS 0.008048f
C1581 B.n728 VSUBS 0.008048f
C1582 B.n729 VSUBS 0.008048f
C1583 B.n730 VSUBS 0.008048f
C1584 B.n731 VSUBS 0.008048f
C1585 B.n732 VSUBS 0.008048f
C1586 B.n733 VSUBS 0.008048f
C1587 B.n734 VSUBS 0.008048f
C1588 B.n735 VSUBS 0.008048f
C1589 B.n736 VSUBS 0.008048f
C1590 B.n737 VSUBS 0.008048f
C1591 B.n738 VSUBS 0.008048f
C1592 B.n739 VSUBS 0.008048f
C1593 B.n740 VSUBS 0.008048f
C1594 B.n741 VSUBS 0.008048f
C1595 B.n742 VSUBS 0.008048f
C1596 B.n743 VSUBS 0.008048f
C1597 B.n744 VSUBS 0.008048f
C1598 B.n745 VSUBS 0.008048f
C1599 B.n746 VSUBS 0.008048f
C1600 B.n747 VSUBS 0.008048f
C1601 B.n748 VSUBS 0.008048f
C1602 B.n749 VSUBS 0.008048f
C1603 B.n750 VSUBS 0.008048f
C1604 B.n751 VSUBS 0.008048f
C1605 B.n752 VSUBS 0.008048f
C1606 B.n753 VSUBS 0.008048f
C1607 B.n754 VSUBS 0.008048f
C1608 B.n755 VSUBS 0.008048f
C1609 B.n756 VSUBS 0.008048f
C1610 B.n757 VSUBS 0.020159f
C1611 B.n758 VSUBS 0.020159f
C1612 B.n759 VSUBS 0.019136f
C1613 B.n760 VSUBS 0.008048f
C1614 B.n761 VSUBS 0.008048f
C1615 B.n762 VSUBS 0.008048f
C1616 B.n763 VSUBS 0.008048f
C1617 B.n764 VSUBS 0.008048f
C1618 B.n765 VSUBS 0.008048f
C1619 B.n766 VSUBS 0.008048f
C1620 B.n767 VSUBS 0.008048f
C1621 B.n768 VSUBS 0.008048f
C1622 B.n769 VSUBS 0.008048f
C1623 B.n770 VSUBS 0.008048f
C1624 B.n771 VSUBS 0.008048f
C1625 B.n772 VSUBS 0.008048f
C1626 B.n773 VSUBS 0.008048f
C1627 B.n774 VSUBS 0.008048f
C1628 B.n775 VSUBS 0.008048f
C1629 B.n776 VSUBS 0.008048f
C1630 B.n777 VSUBS 0.008048f
C1631 B.n778 VSUBS 0.008048f
C1632 B.n779 VSUBS 0.008048f
C1633 B.n780 VSUBS 0.008048f
C1634 B.n781 VSUBS 0.008048f
C1635 B.n782 VSUBS 0.008048f
C1636 B.n783 VSUBS 0.008048f
C1637 B.n784 VSUBS 0.008048f
C1638 B.n785 VSUBS 0.008048f
C1639 B.n786 VSUBS 0.008048f
C1640 B.n787 VSUBS 0.008048f
C1641 B.n788 VSUBS 0.008048f
C1642 B.n789 VSUBS 0.008048f
C1643 B.n790 VSUBS 0.008048f
C1644 B.n791 VSUBS 0.008048f
C1645 B.n792 VSUBS 0.008048f
C1646 B.n793 VSUBS 0.008048f
C1647 B.n794 VSUBS 0.008048f
C1648 B.n795 VSUBS 0.008048f
C1649 B.n796 VSUBS 0.008048f
C1650 B.n797 VSUBS 0.008048f
C1651 B.n798 VSUBS 0.008048f
C1652 B.n799 VSUBS 0.008048f
C1653 B.n800 VSUBS 0.008048f
C1654 B.n801 VSUBS 0.008048f
C1655 B.n802 VSUBS 0.008048f
C1656 B.n803 VSUBS 0.008048f
C1657 B.n804 VSUBS 0.008048f
C1658 B.n805 VSUBS 0.008048f
C1659 B.n806 VSUBS 0.008048f
C1660 B.n807 VSUBS 0.008048f
C1661 B.n808 VSUBS 0.008048f
C1662 B.n809 VSUBS 0.008048f
C1663 B.n810 VSUBS 0.008048f
C1664 B.n811 VSUBS 0.008048f
C1665 B.n812 VSUBS 0.008048f
C1666 B.n813 VSUBS 0.008048f
C1667 B.n814 VSUBS 0.008048f
C1668 B.n815 VSUBS 0.008048f
C1669 B.n816 VSUBS 0.008048f
C1670 B.n817 VSUBS 0.008048f
C1671 B.n818 VSUBS 0.008048f
C1672 B.n819 VSUBS 0.008048f
C1673 B.n820 VSUBS 0.008048f
C1674 B.n821 VSUBS 0.008048f
C1675 B.n822 VSUBS 0.008048f
C1676 B.n823 VSUBS 0.008048f
C1677 B.n824 VSUBS 0.008048f
C1678 B.n825 VSUBS 0.008048f
C1679 B.n826 VSUBS 0.008048f
C1680 B.n827 VSUBS 0.018224f
.ends

