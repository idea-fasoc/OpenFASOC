* NGSPICE file created from diff_pair_sample_1624.ext - technology: sky130A

.subckt diff_pair_sample_1624 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t6 VN.t0 VDD2.t2 w_n2770_n4732# sky130_fd_pr__pfet_01v8 ad=7.3398 pd=38.42 as=3.1053 ps=19.15 w=18.82 l=2.67
X1 VDD1.t3 VP.t0 VTAIL.t7 w_n2770_n4732# sky130_fd_pr__pfet_01v8 ad=3.1053 pd=19.15 as=7.3398 ps=38.42 w=18.82 l=2.67
X2 B.t11 B.t9 B.t10 w_n2770_n4732# sky130_fd_pr__pfet_01v8 ad=7.3398 pd=38.42 as=0 ps=0 w=18.82 l=2.67
X3 VDD2.t0 VN.t1 VTAIL.t5 w_n2770_n4732# sky130_fd_pr__pfet_01v8 ad=3.1053 pd=19.15 as=7.3398 ps=38.42 w=18.82 l=2.67
X4 B.t8 B.t6 B.t7 w_n2770_n4732# sky130_fd_pr__pfet_01v8 ad=7.3398 pd=38.42 as=0 ps=0 w=18.82 l=2.67
X5 VTAIL.t4 VN.t2 VDD2.t3 w_n2770_n4732# sky130_fd_pr__pfet_01v8 ad=7.3398 pd=38.42 as=3.1053 ps=19.15 w=18.82 l=2.67
X6 VDD2.t1 VN.t3 VTAIL.t3 w_n2770_n4732# sky130_fd_pr__pfet_01v8 ad=3.1053 pd=19.15 as=7.3398 ps=38.42 w=18.82 l=2.67
X7 VTAIL.t2 VP.t1 VDD1.t2 w_n2770_n4732# sky130_fd_pr__pfet_01v8 ad=7.3398 pd=38.42 as=3.1053 ps=19.15 w=18.82 l=2.67
X8 VTAIL.t0 VP.t2 VDD1.t1 w_n2770_n4732# sky130_fd_pr__pfet_01v8 ad=7.3398 pd=38.42 as=3.1053 ps=19.15 w=18.82 l=2.67
X9 VDD1.t0 VP.t3 VTAIL.t1 w_n2770_n4732# sky130_fd_pr__pfet_01v8 ad=3.1053 pd=19.15 as=7.3398 ps=38.42 w=18.82 l=2.67
X10 B.t5 B.t3 B.t4 w_n2770_n4732# sky130_fd_pr__pfet_01v8 ad=7.3398 pd=38.42 as=0 ps=0 w=18.82 l=2.67
X11 B.t2 B.t0 B.t1 w_n2770_n4732# sky130_fd_pr__pfet_01v8 ad=7.3398 pd=38.42 as=0 ps=0 w=18.82 l=2.67
R0 VN.n0 VN.t0 203.659
R1 VN.n1 VN.t1 203.659
R2 VN.n0 VN.t3 202.793
R3 VN.n1 VN.t2 202.793
R4 VN VN.n1 55.538
R5 VN VN.n0 3.68577
R6 VDD2.n2 VDD2.n0 120.05
R7 VDD2.n2 VDD2.n1 72.3529
R8 VDD2.n1 VDD2.t3 1.72765
R9 VDD2.n1 VDD2.t0 1.72765
R10 VDD2.n0 VDD2.t2 1.72765
R11 VDD2.n0 VDD2.t1 1.72765
R12 VDD2 VDD2.n2 0.0586897
R13 VTAIL.n830 VTAIL.n829 756.745
R14 VTAIL.n102 VTAIL.n101 756.745
R15 VTAIL.n206 VTAIL.n205 756.745
R16 VTAIL.n310 VTAIL.n309 756.745
R17 VTAIL.n726 VTAIL.n725 756.745
R18 VTAIL.n622 VTAIL.n621 756.745
R19 VTAIL.n518 VTAIL.n517 756.745
R20 VTAIL.n414 VTAIL.n413 756.745
R21 VTAIL.n763 VTAIL.n762 585
R22 VTAIL.n765 VTAIL.n764 585
R23 VTAIL.n758 VTAIL.n757 585
R24 VTAIL.n771 VTAIL.n770 585
R25 VTAIL.n773 VTAIL.n772 585
R26 VTAIL.n754 VTAIL.n753 585
R27 VTAIL.n780 VTAIL.n779 585
R28 VTAIL.n781 VTAIL.n752 585
R29 VTAIL.n783 VTAIL.n782 585
R30 VTAIL.n750 VTAIL.n749 585
R31 VTAIL.n789 VTAIL.n788 585
R32 VTAIL.n791 VTAIL.n790 585
R33 VTAIL.n746 VTAIL.n745 585
R34 VTAIL.n797 VTAIL.n796 585
R35 VTAIL.n799 VTAIL.n798 585
R36 VTAIL.n742 VTAIL.n741 585
R37 VTAIL.n805 VTAIL.n804 585
R38 VTAIL.n807 VTAIL.n806 585
R39 VTAIL.n738 VTAIL.n737 585
R40 VTAIL.n813 VTAIL.n812 585
R41 VTAIL.n815 VTAIL.n814 585
R42 VTAIL.n734 VTAIL.n733 585
R43 VTAIL.n821 VTAIL.n820 585
R44 VTAIL.n823 VTAIL.n822 585
R45 VTAIL.n730 VTAIL.n729 585
R46 VTAIL.n829 VTAIL.n828 585
R47 VTAIL.n35 VTAIL.n34 585
R48 VTAIL.n37 VTAIL.n36 585
R49 VTAIL.n30 VTAIL.n29 585
R50 VTAIL.n43 VTAIL.n42 585
R51 VTAIL.n45 VTAIL.n44 585
R52 VTAIL.n26 VTAIL.n25 585
R53 VTAIL.n52 VTAIL.n51 585
R54 VTAIL.n53 VTAIL.n24 585
R55 VTAIL.n55 VTAIL.n54 585
R56 VTAIL.n22 VTAIL.n21 585
R57 VTAIL.n61 VTAIL.n60 585
R58 VTAIL.n63 VTAIL.n62 585
R59 VTAIL.n18 VTAIL.n17 585
R60 VTAIL.n69 VTAIL.n68 585
R61 VTAIL.n71 VTAIL.n70 585
R62 VTAIL.n14 VTAIL.n13 585
R63 VTAIL.n77 VTAIL.n76 585
R64 VTAIL.n79 VTAIL.n78 585
R65 VTAIL.n10 VTAIL.n9 585
R66 VTAIL.n85 VTAIL.n84 585
R67 VTAIL.n87 VTAIL.n86 585
R68 VTAIL.n6 VTAIL.n5 585
R69 VTAIL.n93 VTAIL.n92 585
R70 VTAIL.n95 VTAIL.n94 585
R71 VTAIL.n2 VTAIL.n1 585
R72 VTAIL.n101 VTAIL.n100 585
R73 VTAIL.n139 VTAIL.n138 585
R74 VTAIL.n141 VTAIL.n140 585
R75 VTAIL.n134 VTAIL.n133 585
R76 VTAIL.n147 VTAIL.n146 585
R77 VTAIL.n149 VTAIL.n148 585
R78 VTAIL.n130 VTAIL.n129 585
R79 VTAIL.n156 VTAIL.n155 585
R80 VTAIL.n157 VTAIL.n128 585
R81 VTAIL.n159 VTAIL.n158 585
R82 VTAIL.n126 VTAIL.n125 585
R83 VTAIL.n165 VTAIL.n164 585
R84 VTAIL.n167 VTAIL.n166 585
R85 VTAIL.n122 VTAIL.n121 585
R86 VTAIL.n173 VTAIL.n172 585
R87 VTAIL.n175 VTAIL.n174 585
R88 VTAIL.n118 VTAIL.n117 585
R89 VTAIL.n181 VTAIL.n180 585
R90 VTAIL.n183 VTAIL.n182 585
R91 VTAIL.n114 VTAIL.n113 585
R92 VTAIL.n189 VTAIL.n188 585
R93 VTAIL.n191 VTAIL.n190 585
R94 VTAIL.n110 VTAIL.n109 585
R95 VTAIL.n197 VTAIL.n196 585
R96 VTAIL.n199 VTAIL.n198 585
R97 VTAIL.n106 VTAIL.n105 585
R98 VTAIL.n205 VTAIL.n204 585
R99 VTAIL.n243 VTAIL.n242 585
R100 VTAIL.n245 VTAIL.n244 585
R101 VTAIL.n238 VTAIL.n237 585
R102 VTAIL.n251 VTAIL.n250 585
R103 VTAIL.n253 VTAIL.n252 585
R104 VTAIL.n234 VTAIL.n233 585
R105 VTAIL.n260 VTAIL.n259 585
R106 VTAIL.n261 VTAIL.n232 585
R107 VTAIL.n263 VTAIL.n262 585
R108 VTAIL.n230 VTAIL.n229 585
R109 VTAIL.n269 VTAIL.n268 585
R110 VTAIL.n271 VTAIL.n270 585
R111 VTAIL.n226 VTAIL.n225 585
R112 VTAIL.n277 VTAIL.n276 585
R113 VTAIL.n279 VTAIL.n278 585
R114 VTAIL.n222 VTAIL.n221 585
R115 VTAIL.n285 VTAIL.n284 585
R116 VTAIL.n287 VTAIL.n286 585
R117 VTAIL.n218 VTAIL.n217 585
R118 VTAIL.n293 VTAIL.n292 585
R119 VTAIL.n295 VTAIL.n294 585
R120 VTAIL.n214 VTAIL.n213 585
R121 VTAIL.n301 VTAIL.n300 585
R122 VTAIL.n303 VTAIL.n302 585
R123 VTAIL.n210 VTAIL.n209 585
R124 VTAIL.n309 VTAIL.n308 585
R125 VTAIL.n725 VTAIL.n724 585
R126 VTAIL.n626 VTAIL.n625 585
R127 VTAIL.n719 VTAIL.n718 585
R128 VTAIL.n717 VTAIL.n716 585
R129 VTAIL.n630 VTAIL.n629 585
R130 VTAIL.n711 VTAIL.n710 585
R131 VTAIL.n709 VTAIL.n708 585
R132 VTAIL.n634 VTAIL.n633 585
R133 VTAIL.n703 VTAIL.n702 585
R134 VTAIL.n701 VTAIL.n700 585
R135 VTAIL.n638 VTAIL.n637 585
R136 VTAIL.n695 VTAIL.n694 585
R137 VTAIL.n693 VTAIL.n692 585
R138 VTAIL.n642 VTAIL.n641 585
R139 VTAIL.n687 VTAIL.n686 585
R140 VTAIL.n685 VTAIL.n684 585
R141 VTAIL.n646 VTAIL.n645 585
R142 VTAIL.n650 VTAIL.n648 585
R143 VTAIL.n679 VTAIL.n678 585
R144 VTAIL.n677 VTAIL.n676 585
R145 VTAIL.n652 VTAIL.n651 585
R146 VTAIL.n671 VTAIL.n670 585
R147 VTAIL.n669 VTAIL.n668 585
R148 VTAIL.n656 VTAIL.n655 585
R149 VTAIL.n663 VTAIL.n662 585
R150 VTAIL.n661 VTAIL.n660 585
R151 VTAIL.n621 VTAIL.n620 585
R152 VTAIL.n522 VTAIL.n521 585
R153 VTAIL.n615 VTAIL.n614 585
R154 VTAIL.n613 VTAIL.n612 585
R155 VTAIL.n526 VTAIL.n525 585
R156 VTAIL.n607 VTAIL.n606 585
R157 VTAIL.n605 VTAIL.n604 585
R158 VTAIL.n530 VTAIL.n529 585
R159 VTAIL.n599 VTAIL.n598 585
R160 VTAIL.n597 VTAIL.n596 585
R161 VTAIL.n534 VTAIL.n533 585
R162 VTAIL.n591 VTAIL.n590 585
R163 VTAIL.n589 VTAIL.n588 585
R164 VTAIL.n538 VTAIL.n537 585
R165 VTAIL.n583 VTAIL.n582 585
R166 VTAIL.n581 VTAIL.n580 585
R167 VTAIL.n542 VTAIL.n541 585
R168 VTAIL.n546 VTAIL.n544 585
R169 VTAIL.n575 VTAIL.n574 585
R170 VTAIL.n573 VTAIL.n572 585
R171 VTAIL.n548 VTAIL.n547 585
R172 VTAIL.n567 VTAIL.n566 585
R173 VTAIL.n565 VTAIL.n564 585
R174 VTAIL.n552 VTAIL.n551 585
R175 VTAIL.n559 VTAIL.n558 585
R176 VTAIL.n557 VTAIL.n556 585
R177 VTAIL.n517 VTAIL.n516 585
R178 VTAIL.n418 VTAIL.n417 585
R179 VTAIL.n511 VTAIL.n510 585
R180 VTAIL.n509 VTAIL.n508 585
R181 VTAIL.n422 VTAIL.n421 585
R182 VTAIL.n503 VTAIL.n502 585
R183 VTAIL.n501 VTAIL.n500 585
R184 VTAIL.n426 VTAIL.n425 585
R185 VTAIL.n495 VTAIL.n494 585
R186 VTAIL.n493 VTAIL.n492 585
R187 VTAIL.n430 VTAIL.n429 585
R188 VTAIL.n487 VTAIL.n486 585
R189 VTAIL.n485 VTAIL.n484 585
R190 VTAIL.n434 VTAIL.n433 585
R191 VTAIL.n479 VTAIL.n478 585
R192 VTAIL.n477 VTAIL.n476 585
R193 VTAIL.n438 VTAIL.n437 585
R194 VTAIL.n442 VTAIL.n440 585
R195 VTAIL.n471 VTAIL.n470 585
R196 VTAIL.n469 VTAIL.n468 585
R197 VTAIL.n444 VTAIL.n443 585
R198 VTAIL.n463 VTAIL.n462 585
R199 VTAIL.n461 VTAIL.n460 585
R200 VTAIL.n448 VTAIL.n447 585
R201 VTAIL.n455 VTAIL.n454 585
R202 VTAIL.n453 VTAIL.n452 585
R203 VTAIL.n413 VTAIL.n412 585
R204 VTAIL.n314 VTAIL.n313 585
R205 VTAIL.n407 VTAIL.n406 585
R206 VTAIL.n405 VTAIL.n404 585
R207 VTAIL.n318 VTAIL.n317 585
R208 VTAIL.n399 VTAIL.n398 585
R209 VTAIL.n397 VTAIL.n396 585
R210 VTAIL.n322 VTAIL.n321 585
R211 VTAIL.n391 VTAIL.n390 585
R212 VTAIL.n389 VTAIL.n388 585
R213 VTAIL.n326 VTAIL.n325 585
R214 VTAIL.n383 VTAIL.n382 585
R215 VTAIL.n381 VTAIL.n380 585
R216 VTAIL.n330 VTAIL.n329 585
R217 VTAIL.n375 VTAIL.n374 585
R218 VTAIL.n373 VTAIL.n372 585
R219 VTAIL.n334 VTAIL.n333 585
R220 VTAIL.n338 VTAIL.n336 585
R221 VTAIL.n367 VTAIL.n366 585
R222 VTAIL.n365 VTAIL.n364 585
R223 VTAIL.n340 VTAIL.n339 585
R224 VTAIL.n359 VTAIL.n358 585
R225 VTAIL.n357 VTAIL.n356 585
R226 VTAIL.n344 VTAIL.n343 585
R227 VTAIL.n351 VTAIL.n350 585
R228 VTAIL.n349 VTAIL.n348 585
R229 VTAIL.n761 VTAIL.t3 329.036
R230 VTAIL.n33 VTAIL.t6 329.036
R231 VTAIL.n137 VTAIL.t7 329.036
R232 VTAIL.n241 VTAIL.t0 329.036
R233 VTAIL.n659 VTAIL.t1 329.036
R234 VTAIL.n555 VTAIL.t2 329.036
R235 VTAIL.n451 VTAIL.t5 329.036
R236 VTAIL.n347 VTAIL.t4 329.036
R237 VTAIL.n764 VTAIL.n763 171.744
R238 VTAIL.n764 VTAIL.n757 171.744
R239 VTAIL.n771 VTAIL.n757 171.744
R240 VTAIL.n772 VTAIL.n771 171.744
R241 VTAIL.n772 VTAIL.n753 171.744
R242 VTAIL.n780 VTAIL.n753 171.744
R243 VTAIL.n781 VTAIL.n780 171.744
R244 VTAIL.n782 VTAIL.n781 171.744
R245 VTAIL.n782 VTAIL.n749 171.744
R246 VTAIL.n789 VTAIL.n749 171.744
R247 VTAIL.n790 VTAIL.n789 171.744
R248 VTAIL.n790 VTAIL.n745 171.744
R249 VTAIL.n797 VTAIL.n745 171.744
R250 VTAIL.n798 VTAIL.n797 171.744
R251 VTAIL.n798 VTAIL.n741 171.744
R252 VTAIL.n805 VTAIL.n741 171.744
R253 VTAIL.n806 VTAIL.n805 171.744
R254 VTAIL.n806 VTAIL.n737 171.744
R255 VTAIL.n813 VTAIL.n737 171.744
R256 VTAIL.n814 VTAIL.n813 171.744
R257 VTAIL.n814 VTAIL.n733 171.744
R258 VTAIL.n821 VTAIL.n733 171.744
R259 VTAIL.n822 VTAIL.n821 171.744
R260 VTAIL.n822 VTAIL.n729 171.744
R261 VTAIL.n829 VTAIL.n729 171.744
R262 VTAIL.n36 VTAIL.n35 171.744
R263 VTAIL.n36 VTAIL.n29 171.744
R264 VTAIL.n43 VTAIL.n29 171.744
R265 VTAIL.n44 VTAIL.n43 171.744
R266 VTAIL.n44 VTAIL.n25 171.744
R267 VTAIL.n52 VTAIL.n25 171.744
R268 VTAIL.n53 VTAIL.n52 171.744
R269 VTAIL.n54 VTAIL.n53 171.744
R270 VTAIL.n54 VTAIL.n21 171.744
R271 VTAIL.n61 VTAIL.n21 171.744
R272 VTAIL.n62 VTAIL.n61 171.744
R273 VTAIL.n62 VTAIL.n17 171.744
R274 VTAIL.n69 VTAIL.n17 171.744
R275 VTAIL.n70 VTAIL.n69 171.744
R276 VTAIL.n70 VTAIL.n13 171.744
R277 VTAIL.n77 VTAIL.n13 171.744
R278 VTAIL.n78 VTAIL.n77 171.744
R279 VTAIL.n78 VTAIL.n9 171.744
R280 VTAIL.n85 VTAIL.n9 171.744
R281 VTAIL.n86 VTAIL.n85 171.744
R282 VTAIL.n86 VTAIL.n5 171.744
R283 VTAIL.n93 VTAIL.n5 171.744
R284 VTAIL.n94 VTAIL.n93 171.744
R285 VTAIL.n94 VTAIL.n1 171.744
R286 VTAIL.n101 VTAIL.n1 171.744
R287 VTAIL.n140 VTAIL.n139 171.744
R288 VTAIL.n140 VTAIL.n133 171.744
R289 VTAIL.n147 VTAIL.n133 171.744
R290 VTAIL.n148 VTAIL.n147 171.744
R291 VTAIL.n148 VTAIL.n129 171.744
R292 VTAIL.n156 VTAIL.n129 171.744
R293 VTAIL.n157 VTAIL.n156 171.744
R294 VTAIL.n158 VTAIL.n157 171.744
R295 VTAIL.n158 VTAIL.n125 171.744
R296 VTAIL.n165 VTAIL.n125 171.744
R297 VTAIL.n166 VTAIL.n165 171.744
R298 VTAIL.n166 VTAIL.n121 171.744
R299 VTAIL.n173 VTAIL.n121 171.744
R300 VTAIL.n174 VTAIL.n173 171.744
R301 VTAIL.n174 VTAIL.n117 171.744
R302 VTAIL.n181 VTAIL.n117 171.744
R303 VTAIL.n182 VTAIL.n181 171.744
R304 VTAIL.n182 VTAIL.n113 171.744
R305 VTAIL.n189 VTAIL.n113 171.744
R306 VTAIL.n190 VTAIL.n189 171.744
R307 VTAIL.n190 VTAIL.n109 171.744
R308 VTAIL.n197 VTAIL.n109 171.744
R309 VTAIL.n198 VTAIL.n197 171.744
R310 VTAIL.n198 VTAIL.n105 171.744
R311 VTAIL.n205 VTAIL.n105 171.744
R312 VTAIL.n244 VTAIL.n243 171.744
R313 VTAIL.n244 VTAIL.n237 171.744
R314 VTAIL.n251 VTAIL.n237 171.744
R315 VTAIL.n252 VTAIL.n251 171.744
R316 VTAIL.n252 VTAIL.n233 171.744
R317 VTAIL.n260 VTAIL.n233 171.744
R318 VTAIL.n261 VTAIL.n260 171.744
R319 VTAIL.n262 VTAIL.n261 171.744
R320 VTAIL.n262 VTAIL.n229 171.744
R321 VTAIL.n269 VTAIL.n229 171.744
R322 VTAIL.n270 VTAIL.n269 171.744
R323 VTAIL.n270 VTAIL.n225 171.744
R324 VTAIL.n277 VTAIL.n225 171.744
R325 VTAIL.n278 VTAIL.n277 171.744
R326 VTAIL.n278 VTAIL.n221 171.744
R327 VTAIL.n285 VTAIL.n221 171.744
R328 VTAIL.n286 VTAIL.n285 171.744
R329 VTAIL.n286 VTAIL.n217 171.744
R330 VTAIL.n293 VTAIL.n217 171.744
R331 VTAIL.n294 VTAIL.n293 171.744
R332 VTAIL.n294 VTAIL.n213 171.744
R333 VTAIL.n301 VTAIL.n213 171.744
R334 VTAIL.n302 VTAIL.n301 171.744
R335 VTAIL.n302 VTAIL.n209 171.744
R336 VTAIL.n309 VTAIL.n209 171.744
R337 VTAIL.n725 VTAIL.n625 171.744
R338 VTAIL.n718 VTAIL.n625 171.744
R339 VTAIL.n718 VTAIL.n717 171.744
R340 VTAIL.n717 VTAIL.n629 171.744
R341 VTAIL.n710 VTAIL.n629 171.744
R342 VTAIL.n710 VTAIL.n709 171.744
R343 VTAIL.n709 VTAIL.n633 171.744
R344 VTAIL.n702 VTAIL.n633 171.744
R345 VTAIL.n702 VTAIL.n701 171.744
R346 VTAIL.n701 VTAIL.n637 171.744
R347 VTAIL.n694 VTAIL.n637 171.744
R348 VTAIL.n694 VTAIL.n693 171.744
R349 VTAIL.n693 VTAIL.n641 171.744
R350 VTAIL.n686 VTAIL.n641 171.744
R351 VTAIL.n686 VTAIL.n685 171.744
R352 VTAIL.n685 VTAIL.n645 171.744
R353 VTAIL.n650 VTAIL.n645 171.744
R354 VTAIL.n678 VTAIL.n650 171.744
R355 VTAIL.n678 VTAIL.n677 171.744
R356 VTAIL.n677 VTAIL.n651 171.744
R357 VTAIL.n670 VTAIL.n651 171.744
R358 VTAIL.n670 VTAIL.n669 171.744
R359 VTAIL.n669 VTAIL.n655 171.744
R360 VTAIL.n662 VTAIL.n655 171.744
R361 VTAIL.n662 VTAIL.n661 171.744
R362 VTAIL.n621 VTAIL.n521 171.744
R363 VTAIL.n614 VTAIL.n521 171.744
R364 VTAIL.n614 VTAIL.n613 171.744
R365 VTAIL.n613 VTAIL.n525 171.744
R366 VTAIL.n606 VTAIL.n525 171.744
R367 VTAIL.n606 VTAIL.n605 171.744
R368 VTAIL.n605 VTAIL.n529 171.744
R369 VTAIL.n598 VTAIL.n529 171.744
R370 VTAIL.n598 VTAIL.n597 171.744
R371 VTAIL.n597 VTAIL.n533 171.744
R372 VTAIL.n590 VTAIL.n533 171.744
R373 VTAIL.n590 VTAIL.n589 171.744
R374 VTAIL.n589 VTAIL.n537 171.744
R375 VTAIL.n582 VTAIL.n537 171.744
R376 VTAIL.n582 VTAIL.n581 171.744
R377 VTAIL.n581 VTAIL.n541 171.744
R378 VTAIL.n546 VTAIL.n541 171.744
R379 VTAIL.n574 VTAIL.n546 171.744
R380 VTAIL.n574 VTAIL.n573 171.744
R381 VTAIL.n573 VTAIL.n547 171.744
R382 VTAIL.n566 VTAIL.n547 171.744
R383 VTAIL.n566 VTAIL.n565 171.744
R384 VTAIL.n565 VTAIL.n551 171.744
R385 VTAIL.n558 VTAIL.n551 171.744
R386 VTAIL.n558 VTAIL.n557 171.744
R387 VTAIL.n517 VTAIL.n417 171.744
R388 VTAIL.n510 VTAIL.n417 171.744
R389 VTAIL.n510 VTAIL.n509 171.744
R390 VTAIL.n509 VTAIL.n421 171.744
R391 VTAIL.n502 VTAIL.n421 171.744
R392 VTAIL.n502 VTAIL.n501 171.744
R393 VTAIL.n501 VTAIL.n425 171.744
R394 VTAIL.n494 VTAIL.n425 171.744
R395 VTAIL.n494 VTAIL.n493 171.744
R396 VTAIL.n493 VTAIL.n429 171.744
R397 VTAIL.n486 VTAIL.n429 171.744
R398 VTAIL.n486 VTAIL.n485 171.744
R399 VTAIL.n485 VTAIL.n433 171.744
R400 VTAIL.n478 VTAIL.n433 171.744
R401 VTAIL.n478 VTAIL.n477 171.744
R402 VTAIL.n477 VTAIL.n437 171.744
R403 VTAIL.n442 VTAIL.n437 171.744
R404 VTAIL.n470 VTAIL.n442 171.744
R405 VTAIL.n470 VTAIL.n469 171.744
R406 VTAIL.n469 VTAIL.n443 171.744
R407 VTAIL.n462 VTAIL.n443 171.744
R408 VTAIL.n462 VTAIL.n461 171.744
R409 VTAIL.n461 VTAIL.n447 171.744
R410 VTAIL.n454 VTAIL.n447 171.744
R411 VTAIL.n454 VTAIL.n453 171.744
R412 VTAIL.n413 VTAIL.n313 171.744
R413 VTAIL.n406 VTAIL.n313 171.744
R414 VTAIL.n406 VTAIL.n405 171.744
R415 VTAIL.n405 VTAIL.n317 171.744
R416 VTAIL.n398 VTAIL.n317 171.744
R417 VTAIL.n398 VTAIL.n397 171.744
R418 VTAIL.n397 VTAIL.n321 171.744
R419 VTAIL.n390 VTAIL.n321 171.744
R420 VTAIL.n390 VTAIL.n389 171.744
R421 VTAIL.n389 VTAIL.n325 171.744
R422 VTAIL.n382 VTAIL.n325 171.744
R423 VTAIL.n382 VTAIL.n381 171.744
R424 VTAIL.n381 VTAIL.n329 171.744
R425 VTAIL.n374 VTAIL.n329 171.744
R426 VTAIL.n374 VTAIL.n373 171.744
R427 VTAIL.n373 VTAIL.n333 171.744
R428 VTAIL.n338 VTAIL.n333 171.744
R429 VTAIL.n366 VTAIL.n338 171.744
R430 VTAIL.n366 VTAIL.n365 171.744
R431 VTAIL.n365 VTAIL.n339 171.744
R432 VTAIL.n358 VTAIL.n339 171.744
R433 VTAIL.n358 VTAIL.n357 171.744
R434 VTAIL.n357 VTAIL.n343 171.744
R435 VTAIL.n350 VTAIL.n343 171.744
R436 VTAIL.n350 VTAIL.n349 171.744
R437 VTAIL.n763 VTAIL.t3 85.8723
R438 VTAIL.n35 VTAIL.t6 85.8723
R439 VTAIL.n139 VTAIL.t7 85.8723
R440 VTAIL.n243 VTAIL.t0 85.8723
R441 VTAIL.n661 VTAIL.t1 85.8723
R442 VTAIL.n557 VTAIL.t2 85.8723
R443 VTAIL.n453 VTAIL.t5 85.8723
R444 VTAIL.n349 VTAIL.t4 85.8723
R445 VTAIL.n831 VTAIL.n830 36.0641
R446 VTAIL.n103 VTAIL.n102 36.0641
R447 VTAIL.n207 VTAIL.n206 36.0641
R448 VTAIL.n311 VTAIL.n310 36.0641
R449 VTAIL.n727 VTAIL.n726 36.0641
R450 VTAIL.n623 VTAIL.n622 36.0641
R451 VTAIL.n519 VTAIL.n518 36.0641
R452 VTAIL.n415 VTAIL.n414 36.0641
R453 VTAIL.n831 VTAIL.n727 31.1772
R454 VTAIL.n415 VTAIL.n311 31.1772
R455 VTAIL.n783 VTAIL.n750 13.1884
R456 VTAIL.n55 VTAIL.n22 13.1884
R457 VTAIL.n159 VTAIL.n126 13.1884
R458 VTAIL.n263 VTAIL.n230 13.1884
R459 VTAIL.n648 VTAIL.n646 13.1884
R460 VTAIL.n544 VTAIL.n542 13.1884
R461 VTAIL.n440 VTAIL.n438 13.1884
R462 VTAIL.n336 VTAIL.n334 13.1884
R463 VTAIL.n784 VTAIL.n752 12.8005
R464 VTAIL.n788 VTAIL.n787 12.8005
R465 VTAIL.n828 VTAIL.n728 12.8005
R466 VTAIL.n56 VTAIL.n24 12.8005
R467 VTAIL.n60 VTAIL.n59 12.8005
R468 VTAIL.n100 VTAIL.n0 12.8005
R469 VTAIL.n160 VTAIL.n128 12.8005
R470 VTAIL.n164 VTAIL.n163 12.8005
R471 VTAIL.n204 VTAIL.n104 12.8005
R472 VTAIL.n264 VTAIL.n232 12.8005
R473 VTAIL.n268 VTAIL.n267 12.8005
R474 VTAIL.n308 VTAIL.n208 12.8005
R475 VTAIL.n724 VTAIL.n624 12.8005
R476 VTAIL.n684 VTAIL.n683 12.8005
R477 VTAIL.n680 VTAIL.n679 12.8005
R478 VTAIL.n620 VTAIL.n520 12.8005
R479 VTAIL.n580 VTAIL.n579 12.8005
R480 VTAIL.n576 VTAIL.n575 12.8005
R481 VTAIL.n516 VTAIL.n416 12.8005
R482 VTAIL.n476 VTAIL.n475 12.8005
R483 VTAIL.n472 VTAIL.n471 12.8005
R484 VTAIL.n412 VTAIL.n312 12.8005
R485 VTAIL.n372 VTAIL.n371 12.8005
R486 VTAIL.n368 VTAIL.n367 12.8005
R487 VTAIL.n779 VTAIL.n778 12.0247
R488 VTAIL.n791 VTAIL.n748 12.0247
R489 VTAIL.n827 VTAIL.n730 12.0247
R490 VTAIL.n51 VTAIL.n50 12.0247
R491 VTAIL.n63 VTAIL.n20 12.0247
R492 VTAIL.n99 VTAIL.n2 12.0247
R493 VTAIL.n155 VTAIL.n154 12.0247
R494 VTAIL.n167 VTAIL.n124 12.0247
R495 VTAIL.n203 VTAIL.n106 12.0247
R496 VTAIL.n259 VTAIL.n258 12.0247
R497 VTAIL.n271 VTAIL.n228 12.0247
R498 VTAIL.n307 VTAIL.n210 12.0247
R499 VTAIL.n723 VTAIL.n626 12.0247
R500 VTAIL.n687 VTAIL.n644 12.0247
R501 VTAIL.n676 VTAIL.n649 12.0247
R502 VTAIL.n619 VTAIL.n522 12.0247
R503 VTAIL.n583 VTAIL.n540 12.0247
R504 VTAIL.n572 VTAIL.n545 12.0247
R505 VTAIL.n515 VTAIL.n418 12.0247
R506 VTAIL.n479 VTAIL.n436 12.0247
R507 VTAIL.n468 VTAIL.n441 12.0247
R508 VTAIL.n411 VTAIL.n314 12.0247
R509 VTAIL.n375 VTAIL.n332 12.0247
R510 VTAIL.n364 VTAIL.n337 12.0247
R511 VTAIL.n777 VTAIL.n754 11.249
R512 VTAIL.n792 VTAIL.n746 11.249
R513 VTAIL.n824 VTAIL.n823 11.249
R514 VTAIL.n49 VTAIL.n26 11.249
R515 VTAIL.n64 VTAIL.n18 11.249
R516 VTAIL.n96 VTAIL.n95 11.249
R517 VTAIL.n153 VTAIL.n130 11.249
R518 VTAIL.n168 VTAIL.n122 11.249
R519 VTAIL.n200 VTAIL.n199 11.249
R520 VTAIL.n257 VTAIL.n234 11.249
R521 VTAIL.n272 VTAIL.n226 11.249
R522 VTAIL.n304 VTAIL.n303 11.249
R523 VTAIL.n720 VTAIL.n719 11.249
R524 VTAIL.n688 VTAIL.n642 11.249
R525 VTAIL.n675 VTAIL.n652 11.249
R526 VTAIL.n616 VTAIL.n615 11.249
R527 VTAIL.n584 VTAIL.n538 11.249
R528 VTAIL.n571 VTAIL.n548 11.249
R529 VTAIL.n512 VTAIL.n511 11.249
R530 VTAIL.n480 VTAIL.n434 11.249
R531 VTAIL.n467 VTAIL.n444 11.249
R532 VTAIL.n408 VTAIL.n407 11.249
R533 VTAIL.n376 VTAIL.n330 11.249
R534 VTAIL.n363 VTAIL.n340 11.249
R535 VTAIL.n762 VTAIL.n761 10.7239
R536 VTAIL.n34 VTAIL.n33 10.7239
R537 VTAIL.n138 VTAIL.n137 10.7239
R538 VTAIL.n242 VTAIL.n241 10.7239
R539 VTAIL.n660 VTAIL.n659 10.7239
R540 VTAIL.n556 VTAIL.n555 10.7239
R541 VTAIL.n452 VTAIL.n451 10.7239
R542 VTAIL.n348 VTAIL.n347 10.7239
R543 VTAIL.n774 VTAIL.n773 10.4732
R544 VTAIL.n796 VTAIL.n795 10.4732
R545 VTAIL.n820 VTAIL.n732 10.4732
R546 VTAIL.n46 VTAIL.n45 10.4732
R547 VTAIL.n68 VTAIL.n67 10.4732
R548 VTAIL.n92 VTAIL.n4 10.4732
R549 VTAIL.n150 VTAIL.n149 10.4732
R550 VTAIL.n172 VTAIL.n171 10.4732
R551 VTAIL.n196 VTAIL.n108 10.4732
R552 VTAIL.n254 VTAIL.n253 10.4732
R553 VTAIL.n276 VTAIL.n275 10.4732
R554 VTAIL.n300 VTAIL.n212 10.4732
R555 VTAIL.n716 VTAIL.n628 10.4732
R556 VTAIL.n692 VTAIL.n691 10.4732
R557 VTAIL.n672 VTAIL.n671 10.4732
R558 VTAIL.n612 VTAIL.n524 10.4732
R559 VTAIL.n588 VTAIL.n587 10.4732
R560 VTAIL.n568 VTAIL.n567 10.4732
R561 VTAIL.n508 VTAIL.n420 10.4732
R562 VTAIL.n484 VTAIL.n483 10.4732
R563 VTAIL.n464 VTAIL.n463 10.4732
R564 VTAIL.n404 VTAIL.n316 10.4732
R565 VTAIL.n380 VTAIL.n379 10.4732
R566 VTAIL.n360 VTAIL.n359 10.4732
R567 VTAIL.n770 VTAIL.n756 9.69747
R568 VTAIL.n799 VTAIL.n744 9.69747
R569 VTAIL.n819 VTAIL.n734 9.69747
R570 VTAIL.n42 VTAIL.n28 9.69747
R571 VTAIL.n71 VTAIL.n16 9.69747
R572 VTAIL.n91 VTAIL.n6 9.69747
R573 VTAIL.n146 VTAIL.n132 9.69747
R574 VTAIL.n175 VTAIL.n120 9.69747
R575 VTAIL.n195 VTAIL.n110 9.69747
R576 VTAIL.n250 VTAIL.n236 9.69747
R577 VTAIL.n279 VTAIL.n224 9.69747
R578 VTAIL.n299 VTAIL.n214 9.69747
R579 VTAIL.n715 VTAIL.n630 9.69747
R580 VTAIL.n695 VTAIL.n640 9.69747
R581 VTAIL.n668 VTAIL.n654 9.69747
R582 VTAIL.n611 VTAIL.n526 9.69747
R583 VTAIL.n591 VTAIL.n536 9.69747
R584 VTAIL.n564 VTAIL.n550 9.69747
R585 VTAIL.n507 VTAIL.n422 9.69747
R586 VTAIL.n487 VTAIL.n432 9.69747
R587 VTAIL.n460 VTAIL.n446 9.69747
R588 VTAIL.n403 VTAIL.n318 9.69747
R589 VTAIL.n383 VTAIL.n328 9.69747
R590 VTAIL.n356 VTAIL.n342 9.69747
R591 VTAIL.n826 VTAIL.n728 9.45567
R592 VTAIL.n98 VTAIL.n0 9.45567
R593 VTAIL.n202 VTAIL.n104 9.45567
R594 VTAIL.n306 VTAIL.n208 9.45567
R595 VTAIL.n722 VTAIL.n624 9.45567
R596 VTAIL.n618 VTAIL.n520 9.45567
R597 VTAIL.n514 VTAIL.n416 9.45567
R598 VTAIL.n410 VTAIL.n312 9.45567
R599 VTAIL.n809 VTAIL.n808 9.3005
R600 VTAIL.n811 VTAIL.n810 9.3005
R601 VTAIL.n736 VTAIL.n735 9.3005
R602 VTAIL.n817 VTAIL.n816 9.3005
R603 VTAIL.n819 VTAIL.n818 9.3005
R604 VTAIL.n732 VTAIL.n731 9.3005
R605 VTAIL.n825 VTAIL.n824 9.3005
R606 VTAIL.n827 VTAIL.n826 9.3005
R607 VTAIL.n803 VTAIL.n802 9.3005
R608 VTAIL.n801 VTAIL.n800 9.3005
R609 VTAIL.n744 VTAIL.n743 9.3005
R610 VTAIL.n795 VTAIL.n794 9.3005
R611 VTAIL.n793 VTAIL.n792 9.3005
R612 VTAIL.n748 VTAIL.n747 9.3005
R613 VTAIL.n787 VTAIL.n786 9.3005
R614 VTAIL.n760 VTAIL.n759 9.3005
R615 VTAIL.n767 VTAIL.n766 9.3005
R616 VTAIL.n769 VTAIL.n768 9.3005
R617 VTAIL.n756 VTAIL.n755 9.3005
R618 VTAIL.n775 VTAIL.n774 9.3005
R619 VTAIL.n777 VTAIL.n776 9.3005
R620 VTAIL.n778 VTAIL.n751 9.3005
R621 VTAIL.n785 VTAIL.n784 9.3005
R622 VTAIL.n740 VTAIL.n739 9.3005
R623 VTAIL.n81 VTAIL.n80 9.3005
R624 VTAIL.n83 VTAIL.n82 9.3005
R625 VTAIL.n8 VTAIL.n7 9.3005
R626 VTAIL.n89 VTAIL.n88 9.3005
R627 VTAIL.n91 VTAIL.n90 9.3005
R628 VTAIL.n4 VTAIL.n3 9.3005
R629 VTAIL.n97 VTAIL.n96 9.3005
R630 VTAIL.n99 VTAIL.n98 9.3005
R631 VTAIL.n75 VTAIL.n74 9.3005
R632 VTAIL.n73 VTAIL.n72 9.3005
R633 VTAIL.n16 VTAIL.n15 9.3005
R634 VTAIL.n67 VTAIL.n66 9.3005
R635 VTAIL.n65 VTAIL.n64 9.3005
R636 VTAIL.n20 VTAIL.n19 9.3005
R637 VTAIL.n59 VTAIL.n58 9.3005
R638 VTAIL.n32 VTAIL.n31 9.3005
R639 VTAIL.n39 VTAIL.n38 9.3005
R640 VTAIL.n41 VTAIL.n40 9.3005
R641 VTAIL.n28 VTAIL.n27 9.3005
R642 VTAIL.n47 VTAIL.n46 9.3005
R643 VTAIL.n49 VTAIL.n48 9.3005
R644 VTAIL.n50 VTAIL.n23 9.3005
R645 VTAIL.n57 VTAIL.n56 9.3005
R646 VTAIL.n12 VTAIL.n11 9.3005
R647 VTAIL.n185 VTAIL.n184 9.3005
R648 VTAIL.n187 VTAIL.n186 9.3005
R649 VTAIL.n112 VTAIL.n111 9.3005
R650 VTAIL.n193 VTAIL.n192 9.3005
R651 VTAIL.n195 VTAIL.n194 9.3005
R652 VTAIL.n108 VTAIL.n107 9.3005
R653 VTAIL.n201 VTAIL.n200 9.3005
R654 VTAIL.n203 VTAIL.n202 9.3005
R655 VTAIL.n179 VTAIL.n178 9.3005
R656 VTAIL.n177 VTAIL.n176 9.3005
R657 VTAIL.n120 VTAIL.n119 9.3005
R658 VTAIL.n171 VTAIL.n170 9.3005
R659 VTAIL.n169 VTAIL.n168 9.3005
R660 VTAIL.n124 VTAIL.n123 9.3005
R661 VTAIL.n163 VTAIL.n162 9.3005
R662 VTAIL.n136 VTAIL.n135 9.3005
R663 VTAIL.n143 VTAIL.n142 9.3005
R664 VTAIL.n145 VTAIL.n144 9.3005
R665 VTAIL.n132 VTAIL.n131 9.3005
R666 VTAIL.n151 VTAIL.n150 9.3005
R667 VTAIL.n153 VTAIL.n152 9.3005
R668 VTAIL.n154 VTAIL.n127 9.3005
R669 VTAIL.n161 VTAIL.n160 9.3005
R670 VTAIL.n116 VTAIL.n115 9.3005
R671 VTAIL.n289 VTAIL.n288 9.3005
R672 VTAIL.n291 VTAIL.n290 9.3005
R673 VTAIL.n216 VTAIL.n215 9.3005
R674 VTAIL.n297 VTAIL.n296 9.3005
R675 VTAIL.n299 VTAIL.n298 9.3005
R676 VTAIL.n212 VTAIL.n211 9.3005
R677 VTAIL.n305 VTAIL.n304 9.3005
R678 VTAIL.n307 VTAIL.n306 9.3005
R679 VTAIL.n283 VTAIL.n282 9.3005
R680 VTAIL.n281 VTAIL.n280 9.3005
R681 VTAIL.n224 VTAIL.n223 9.3005
R682 VTAIL.n275 VTAIL.n274 9.3005
R683 VTAIL.n273 VTAIL.n272 9.3005
R684 VTAIL.n228 VTAIL.n227 9.3005
R685 VTAIL.n267 VTAIL.n266 9.3005
R686 VTAIL.n240 VTAIL.n239 9.3005
R687 VTAIL.n247 VTAIL.n246 9.3005
R688 VTAIL.n249 VTAIL.n248 9.3005
R689 VTAIL.n236 VTAIL.n235 9.3005
R690 VTAIL.n255 VTAIL.n254 9.3005
R691 VTAIL.n257 VTAIL.n256 9.3005
R692 VTAIL.n258 VTAIL.n231 9.3005
R693 VTAIL.n265 VTAIL.n264 9.3005
R694 VTAIL.n220 VTAIL.n219 9.3005
R695 VTAIL.n723 VTAIL.n722 9.3005
R696 VTAIL.n721 VTAIL.n720 9.3005
R697 VTAIL.n628 VTAIL.n627 9.3005
R698 VTAIL.n715 VTAIL.n714 9.3005
R699 VTAIL.n713 VTAIL.n712 9.3005
R700 VTAIL.n632 VTAIL.n631 9.3005
R701 VTAIL.n707 VTAIL.n706 9.3005
R702 VTAIL.n705 VTAIL.n704 9.3005
R703 VTAIL.n636 VTAIL.n635 9.3005
R704 VTAIL.n699 VTAIL.n698 9.3005
R705 VTAIL.n697 VTAIL.n696 9.3005
R706 VTAIL.n640 VTAIL.n639 9.3005
R707 VTAIL.n691 VTAIL.n690 9.3005
R708 VTAIL.n689 VTAIL.n688 9.3005
R709 VTAIL.n644 VTAIL.n643 9.3005
R710 VTAIL.n683 VTAIL.n682 9.3005
R711 VTAIL.n681 VTAIL.n680 9.3005
R712 VTAIL.n649 VTAIL.n647 9.3005
R713 VTAIL.n675 VTAIL.n674 9.3005
R714 VTAIL.n673 VTAIL.n672 9.3005
R715 VTAIL.n654 VTAIL.n653 9.3005
R716 VTAIL.n667 VTAIL.n666 9.3005
R717 VTAIL.n665 VTAIL.n664 9.3005
R718 VTAIL.n658 VTAIL.n657 9.3005
R719 VTAIL.n554 VTAIL.n553 9.3005
R720 VTAIL.n561 VTAIL.n560 9.3005
R721 VTAIL.n563 VTAIL.n562 9.3005
R722 VTAIL.n550 VTAIL.n549 9.3005
R723 VTAIL.n569 VTAIL.n568 9.3005
R724 VTAIL.n571 VTAIL.n570 9.3005
R725 VTAIL.n545 VTAIL.n543 9.3005
R726 VTAIL.n577 VTAIL.n576 9.3005
R727 VTAIL.n603 VTAIL.n602 9.3005
R728 VTAIL.n528 VTAIL.n527 9.3005
R729 VTAIL.n609 VTAIL.n608 9.3005
R730 VTAIL.n611 VTAIL.n610 9.3005
R731 VTAIL.n524 VTAIL.n523 9.3005
R732 VTAIL.n617 VTAIL.n616 9.3005
R733 VTAIL.n619 VTAIL.n618 9.3005
R734 VTAIL.n601 VTAIL.n600 9.3005
R735 VTAIL.n532 VTAIL.n531 9.3005
R736 VTAIL.n595 VTAIL.n594 9.3005
R737 VTAIL.n593 VTAIL.n592 9.3005
R738 VTAIL.n536 VTAIL.n535 9.3005
R739 VTAIL.n587 VTAIL.n586 9.3005
R740 VTAIL.n585 VTAIL.n584 9.3005
R741 VTAIL.n540 VTAIL.n539 9.3005
R742 VTAIL.n579 VTAIL.n578 9.3005
R743 VTAIL.n450 VTAIL.n449 9.3005
R744 VTAIL.n457 VTAIL.n456 9.3005
R745 VTAIL.n459 VTAIL.n458 9.3005
R746 VTAIL.n446 VTAIL.n445 9.3005
R747 VTAIL.n465 VTAIL.n464 9.3005
R748 VTAIL.n467 VTAIL.n466 9.3005
R749 VTAIL.n441 VTAIL.n439 9.3005
R750 VTAIL.n473 VTAIL.n472 9.3005
R751 VTAIL.n499 VTAIL.n498 9.3005
R752 VTAIL.n424 VTAIL.n423 9.3005
R753 VTAIL.n505 VTAIL.n504 9.3005
R754 VTAIL.n507 VTAIL.n506 9.3005
R755 VTAIL.n420 VTAIL.n419 9.3005
R756 VTAIL.n513 VTAIL.n512 9.3005
R757 VTAIL.n515 VTAIL.n514 9.3005
R758 VTAIL.n497 VTAIL.n496 9.3005
R759 VTAIL.n428 VTAIL.n427 9.3005
R760 VTAIL.n491 VTAIL.n490 9.3005
R761 VTAIL.n489 VTAIL.n488 9.3005
R762 VTAIL.n432 VTAIL.n431 9.3005
R763 VTAIL.n483 VTAIL.n482 9.3005
R764 VTAIL.n481 VTAIL.n480 9.3005
R765 VTAIL.n436 VTAIL.n435 9.3005
R766 VTAIL.n475 VTAIL.n474 9.3005
R767 VTAIL.n346 VTAIL.n345 9.3005
R768 VTAIL.n353 VTAIL.n352 9.3005
R769 VTAIL.n355 VTAIL.n354 9.3005
R770 VTAIL.n342 VTAIL.n341 9.3005
R771 VTAIL.n361 VTAIL.n360 9.3005
R772 VTAIL.n363 VTAIL.n362 9.3005
R773 VTAIL.n337 VTAIL.n335 9.3005
R774 VTAIL.n369 VTAIL.n368 9.3005
R775 VTAIL.n395 VTAIL.n394 9.3005
R776 VTAIL.n320 VTAIL.n319 9.3005
R777 VTAIL.n401 VTAIL.n400 9.3005
R778 VTAIL.n403 VTAIL.n402 9.3005
R779 VTAIL.n316 VTAIL.n315 9.3005
R780 VTAIL.n409 VTAIL.n408 9.3005
R781 VTAIL.n411 VTAIL.n410 9.3005
R782 VTAIL.n393 VTAIL.n392 9.3005
R783 VTAIL.n324 VTAIL.n323 9.3005
R784 VTAIL.n387 VTAIL.n386 9.3005
R785 VTAIL.n385 VTAIL.n384 9.3005
R786 VTAIL.n328 VTAIL.n327 9.3005
R787 VTAIL.n379 VTAIL.n378 9.3005
R788 VTAIL.n377 VTAIL.n376 9.3005
R789 VTAIL.n332 VTAIL.n331 9.3005
R790 VTAIL.n371 VTAIL.n370 9.3005
R791 VTAIL.n769 VTAIL.n758 8.92171
R792 VTAIL.n800 VTAIL.n742 8.92171
R793 VTAIL.n816 VTAIL.n815 8.92171
R794 VTAIL.n41 VTAIL.n30 8.92171
R795 VTAIL.n72 VTAIL.n14 8.92171
R796 VTAIL.n88 VTAIL.n87 8.92171
R797 VTAIL.n145 VTAIL.n134 8.92171
R798 VTAIL.n176 VTAIL.n118 8.92171
R799 VTAIL.n192 VTAIL.n191 8.92171
R800 VTAIL.n249 VTAIL.n238 8.92171
R801 VTAIL.n280 VTAIL.n222 8.92171
R802 VTAIL.n296 VTAIL.n295 8.92171
R803 VTAIL.n712 VTAIL.n711 8.92171
R804 VTAIL.n696 VTAIL.n638 8.92171
R805 VTAIL.n667 VTAIL.n656 8.92171
R806 VTAIL.n608 VTAIL.n607 8.92171
R807 VTAIL.n592 VTAIL.n534 8.92171
R808 VTAIL.n563 VTAIL.n552 8.92171
R809 VTAIL.n504 VTAIL.n503 8.92171
R810 VTAIL.n488 VTAIL.n430 8.92171
R811 VTAIL.n459 VTAIL.n448 8.92171
R812 VTAIL.n400 VTAIL.n399 8.92171
R813 VTAIL.n384 VTAIL.n326 8.92171
R814 VTAIL.n355 VTAIL.n344 8.92171
R815 VTAIL.n766 VTAIL.n765 8.14595
R816 VTAIL.n804 VTAIL.n803 8.14595
R817 VTAIL.n812 VTAIL.n736 8.14595
R818 VTAIL.n38 VTAIL.n37 8.14595
R819 VTAIL.n76 VTAIL.n75 8.14595
R820 VTAIL.n84 VTAIL.n8 8.14595
R821 VTAIL.n142 VTAIL.n141 8.14595
R822 VTAIL.n180 VTAIL.n179 8.14595
R823 VTAIL.n188 VTAIL.n112 8.14595
R824 VTAIL.n246 VTAIL.n245 8.14595
R825 VTAIL.n284 VTAIL.n283 8.14595
R826 VTAIL.n292 VTAIL.n216 8.14595
R827 VTAIL.n708 VTAIL.n632 8.14595
R828 VTAIL.n700 VTAIL.n699 8.14595
R829 VTAIL.n664 VTAIL.n663 8.14595
R830 VTAIL.n604 VTAIL.n528 8.14595
R831 VTAIL.n596 VTAIL.n595 8.14595
R832 VTAIL.n560 VTAIL.n559 8.14595
R833 VTAIL.n500 VTAIL.n424 8.14595
R834 VTAIL.n492 VTAIL.n491 8.14595
R835 VTAIL.n456 VTAIL.n455 8.14595
R836 VTAIL.n396 VTAIL.n320 8.14595
R837 VTAIL.n388 VTAIL.n387 8.14595
R838 VTAIL.n352 VTAIL.n351 8.14595
R839 VTAIL.n762 VTAIL.n760 7.3702
R840 VTAIL.n807 VTAIL.n740 7.3702
R841 VTAIL.n811 VTAIL.n738 7.3702
R842 VTAIL.n34 VTAIL.n32 7.3702
R843 VTAIL.n79 VTAIL.n12 7.3702
R844 VTAIL.n83 VTAIL.n10 7.3702
R845 VTAIL.n138 VTAIL.n136 7.3702
R846 VTAIL.n183 VTAIL.n116 7.3702
R847 VTAIL.n187 VTAIL.n114 7.3702
R848 VTAIL.n242 VTAIL.n240 7.3702
R849 VTAIL.n287 VTAIL.n220 7.3702
R850 VTAIL.n291 VTAIL.n218 7.3702
R851 VTAIL.n707 VTAIL.n634 7.3702
R852 VTAIL.n703 VTAIL.n636 7.3702
R853 VTAIL.n660 VTAIL.n658 7.3702
R854 VTAIL.n603 VTAIL.n530 7.3702
R855 VTAIL.n599 VTAIL.n532 7.3702
R856 VTAIL.n556 VTAIL.n554 7.3702
R857 VTAIL.n499 VTAIL.n426 7.3702
R858 VTAIL.n495 VTAIL.n428 7.3702
R859 VTAIL.n452 VTAIL.n450 7.3702
R860 VTAIL.n395 VTAIL.n322 7.3702
R861 VTAIL.n391 VTAIL.n324 7.3702
R862 VTAIL.n348 VTAIL.n346 7.3702
R863 VTAIL.n808 VTAIL.n807 6.59444
R864 VTAIL.n808 VTAIL.n738 6.59444
R865 VTAIL.n80 VTAIL.n79 6.59444
R866 VTAIL.n80 VTAIL.n10 6.59444
R867 VTAIL.n184 VTAIL.n183 6.59444
R868 VTAIL.n184 VTAIL.n114 6.59444
R869 VTAIL.n288 VTAIL.n287 6.59444
R870 VTAIL.n288 VTAIL.n218 6.59444
R871 VTAIL.n704 VTAIL.n634 6.59444
R872 VTAIL.n704 VTAIL.n703 6.59444
R873 VTAIL.n600 VTAIL.n530 6.59444
R874 VTAIL.n600 VTAIL.n599 6.59444
R875 VTAIL.n496 VTAIL.n426 6.59444
R876 VTAIL.n496 VTAIL.n495 6.59444
R877 VTAIL.n392 VTAIL.n322 6.59444
R878 VTAIL.n392 VTAIL.n391 6.59444
R879 VTAIL.n765 VTAIL.n760 5.81868
R880 VTAIL.n804 VTAIL.n740 5.81868
R881 VTAIL.n812 VTAIL.n811 5.81868
R882 VTAIL.n37 VTAIL.n32 5.81868
R883 VTAIL.n76 VTAIL.n12 5.81868
R884 VTAIL.n84 VTAIL.n83 5.81868
R885 VTAIL.n141 VTAIL.n136 5.81868
R886 VTAIL.n180 VTAIL.n116 5.81868
R887 VTAIL.n188 VTAIL.n187 5.81868
R888 VTAIL.n245 VTAIL.n240 5.81868
R889 VTAIL.n284 VTAIL.n220 5.81868
R890 VTAIL.n292 VTAIL.n291 5.81868
R891 VTAIL.n708 VTAIL.n707 5.81868
R892 VTAIL.n700 VTAIL.n636 5.81868
R893 VTAIL.n663 VTAIL.n658 5.81868
R894 VTAIL.n604 VTAIL.n603 5.81868
R895 VTAIL.n596 VTAIL.n532 5.81868
R896 VTAIL.n559 VTAIL.n554 5.81868
R897 VTAIL.n500 VTAIL.n499 5.81868
R898 VTAIL.n492 VTAIL.n428 5.81868
R899 VTAIL.n455 VTAIL.n450 5.81868
R900 VTAIL.n396 VTAIL.n395 5.81868
R901 VTAIL.n388 VTAIL.n324 5.81868
R902 VTAIL.n351 VTAIL.n346 5.81868
R903 VTAIL.n766 VTAIL.n758 5.04292
R904 VTAIL.n803 VTAIL.n742 5.04292
R905 VTAIL.n815 VTAIL.n736 5.04292
R906 VTAIL.n38 VTAIL.n30 5.04292
R907 VTAIL.n75 VTAIL.n14 5.04292
R908 VTAIL.n87 VTAIL.n8 5.04292
R909 VTAIL.n142 VTAIL.n134 5.04292
R910 VTAIL.n179 VTAIL.n118 5.04292
R911 VTAIL.n191 VTAIL.n112 5.04292
R912 VTAIL.n246 VTAIL.n238 5.04292
R913 VTAIL.n283 VTAIL.n222 5.04292
R914 VTAIL.n295 VTAIL.n216 5.04292
R915 VTAIL.n711 VTAIL.n632 5.04292
R916 VTAIL.n699 VTAIL.n638 5.04292
R917 VTAIL.n664 VTAIL.n656 5.04292
R918 VTAIL.n607 VTAIL.n528 5.04292
R919 VTAIL.n595 VTAIL.n534 5.04292
R920 VTAIL.n560 VTAIL.n552 5.04292
R921 VTAIL.n503 VTAIL.n424 5.04292
R922 VTAIL.n491 VTAIL.n430 5.04292
R923 VTAIL.n456 VTAIL.n448 5.04292
R924 VTAIL.n399 VTAIL.n320 5.04292
R925 VTAIL.n387 VTAIL.n326 5.04292
R926 VTAIL.n352 VTAIL.n344 5.04292
R927 VTAIL.n770 VTAIL.n769 4.26717
R928 VTAIL.n800 VTAIL.n799 4.26717
R929 VTAIL.n816 VTAIL.n734 4.26717
R930 VTAIL.n42 VTAIL.n41 4.26717
R931 VTAIL.n72 VTAIL.n71 4.26717
R932 VTAIL.n88 VTAIL.n6 4.26717
R933 VTAIL.n146 VTAIL.n145 4.26717
R934 VTAIL.n176 VTAIL.n175 4.26717
R935 VTAIL.n192 VTAIL.n110 4.26717
R936 VTAIL.n250 VTAIL.n249 4.26717
R937 VTAIL.n280 VTAIL.n279 4.26717
R938 VTAIL.n296 VTAIL.n214 4.26717
R939 VTAIL.n712 VTAIL.n630 4.26717
R940 VTAIL.n696 VTAIL.n695 4.26717
R941 VTAIL.n668 VTAIL.n667 4.26717
R942 VTAIL.n608 VTAIL.n526 4.26717
R943 VTAIL.n592 VTAIL.n591 4.26717
R944 VTAIL.n564 VTAIL.n563 4.26717
R945 VTAIL.n504 VTAIL.n422 4.26717
R946 VTAIL.n488 VTAIL.n487 4.26717
R947 VTAIL.n460 VTAIL.n459 4.26717
R948 VTAIL.n400 VTAIL.n318 4.26717
R949 VTAIL.n384 VTAIL.n383 4.26717
R950 VTAIL.n356 VTAIL.n355 4.26717
R951 VTAIL.n773 VTAIL.n756 3.49141
R952 VTAIL.n796 VTAIL.n744 3.49141
R953 VTAIL.n820 VTAIL.n819 3.49141
R954 VTAIL.n45 VTAIL.n28 3.49141
R955 VTAIL.n68 VTAIL.n16 3.49141
R956 VTAIL.n92 VTAIL.n91 3.49141
R957 VTAIL.n149 VTAIL.n132 3.49141
R958 VTAIL.n172 VTAIL.n120 3.49141
R959 VTAIL.n196 VTAIL.n195 3.49141
R960 VTAIL.n253 VTAIL.n236 3.49141
R961 VTAIL.n276 VTAIL.n224 3.49141
R962 VTAIL.n300 VTAIL.n299 3.49141
R963 VTAIL.n716 VTAIL.n715 3.49141
R964 VTAIL.n692 VTAIL.n640 3.49141
R965 VTAIL.n671 VTAIL.n654 3.49141
R966 VTAIL.n612 VTAIL.n611 3.49141
R967 VTAIL.n588 VTAIL.n536 3.49141
R968 VTAIL.n567 VTAIL.n550 3.49141
R969 VTAIL.n508 VTAIL.n507 3.49141
R970 VTAIL.n484 VTAIL.n432 3.49141
R971 VTAIL.n463 VTAIL.n446 3.49141
R972 VTAIL.n404 VTAIL.n403 3.49141
R973 VTAIL.n380 VTAIL.n328 3.49141
R974 VTAIL.n359 VTAIL.n342 3.49141
R975 VTAIL.n774 VTAIL.n754 2.71565
R976 VTAIL.n795 VTAIL.n746 2.71565
R977 VTAIL.n823 VTAIL.n732 2.71565
R978 VTAIL.n46 VTAIL.n26 2.71565
R979 VTAIL.n67 VTAIL.n18 2.71565
R980 VTAIL.n95 VTAIL.n4 2.71565
R981 VTAIL.n150 VTAIL.n130 2.71565
R982 VTAIL.n171 VTAIL.n122 2.71565
R983 VTAIL.n199 VTAIL.n108 2.71565
R984 VTAIL.n254 VTAIL.n234 2.71565
R985 VTAIL.n275 VTAIL.n226 2.71565
R986 VTAIL.n303 VTAIL.n212 2.71565
R987 VTAIL.n719 VTAIL.n628 2.71565
R988 VTAIL.n691 VTAIL.n642 2.71565
R989 VTAIL.n672 VTAIL.n652 2.71565
R990 VTAIL.n615 VTAIL.n524 2.71565
R991 VTAIL.n587 VTAIL.n538 2.71565
R992 VTAIL.n568 VTAIL.n548 2.71565
R993 VTAIL.n511 VTAIL.n420 2.71565
R994 VTAIL.n483 VTAIL.n434 2.71565
R995 VTAIL.n464 VTAIL.n444 2.71565
R996 VTAIL.n407 VTAIL.n316 2.71565
R997 VTAIL.n379 VTAIL.n330 2.71565
R998 VTAIL.n360 VTAIL.n340 2.71565
R999 VTAIL.n519 VTAIL.n415 2.58671
R1000 VTAIL.n727 VTAIL.n623 2.58671
R1001 VTAIL.n311 VTAIL.n207 2.58671
R1002 VTAIL.n659 VTAIL.n657 2.41282
R1003 VTAIL.n555 VTAIL.n553 2.41282
R1004 VTAIL.n451 VTAIL.n449 2.41282
R1005 VTAIL.n347 VTAIL.n345 2.41282
R1006 VTAIL.n761 VTAIL.n759 2.41282
R1007 VTAIL.n33 VTAIL.n31 2.41282
R1008 VTAIL.n137 VTAIL.n135 2.41282
R1009 VTAIL.n241 VTAIL.n239 2.41282
R1010 VTAIL.n779 VTAIL.n777 1.93989
R1011 VTAIL.n792 VTAIL.n791 1.93989
R1012 VTAIL.n824 VTAIL.n730 1.93989
R1013 VTAIL.n51 VTAIL.n49 1.93989
R1014 VTAIL.n64 VTAIL.n63 1.93989
R1015 VTAIL.n96 VTAIL.n2 1.93989
R1016 VTAIL.n155 VTAIL.n153 1.93989
R1017 VTAIL.n168 VTAIL.n167 1.93989
R1018 VTAIL.n200 VTAIL.n106 1.93989
R1019 VTAIL.n259 VTAIL.n257 1.93989
R1020 VTAIL.n272 VTAIL.n271 1.93989
R1021 VTAIL.n304 VTAIL.n210 1.93989
R1022 VTAIL.n720 VTAIL.n626 1.93989
R1023 VTAIL.n688 VTAIL.n687 1.93989
R1024 VTAIL.n676 VTAIL.n675 1.93989
R1025 VTAIL.n616 VTAIL.n522 1.93989
R1026 VTAIL.n584 VTAIL.n583 1.93989
R1027 VTAIL.n572 VTAIL.n571 1.93989
R1028 VTAIL.n512 VTAIL.n418 1.93989
R1029 VTAIL.n480 VTAIL.n479 1.93989
R1030 VTAIL.n468 VTAIL.n467 1.93989
R1031 VTAIL.n408 VTAIL.n314 1.93989
R1032 VTAIL.n376 VTAIL.n375 1.93989
R1033 VTAIL.n364 VTAIL.n363 1.93989
R1034 VTAIL VTAIL.n103 1.35179
R1035 VTAIL VTAIL.n831 1.23541
R1036 VTAIL.n778 VTAIL.n752 1.16414
R1037 VTAIL.n788 VTAIL.n748 1.16414
R1038 VTAIL.n828 VTAIL.n827 1.16414
R1039 VTAIL.n50 VTAIL.n24 1.16414
R1040 VTAIL.n60 VTAIL.n20 1.16414
R1041 VTAIL.n100 VTAIL.n99 1.16414
R1042 VTAIL.n154 VTAIL.n128 1.16414
R1043 VTAIL.n164 VTAIL.n124 1.16414
R1044 VTAIL.n204 VTAIL.n203 1.16414
R1045 VTAIL.n258 VTAIL.n232 1.16414
R1046 VTAIL.n268 VTAIL.n228 1.16414
R1047 VTAIL.n308 VTAIL.n307 1.16414
R1048 VTAIL.n724 VTAIL.n723 1.16414
R1049 VTAIL.n684 VTAIL.n644 1.16414
R1050 VTAIL.n679 VTAIL.n649 1.16414
R1051 VTAIL.n620 VTAIL.n619 1.16414
R1052 VTAIL.n580 VTAIL.n540 1.16414
R1053 VTAIL.n575 VTAIL.n545 1.16414
R1054 VTAIL.n516 VTAIL.n515 1.16414
R1055 VTAIL.n476 VTAIL.n436 1.16414
R1056 VTAIL.n471 VTAIL.n441 1.16414
R1057 VTAIL.n412 VTAIL.n411 1.16414
R1058 VTAIL.n372 VTAIL.n332 1.16414
R1059 VTAIL.n367 VTAIL.n337 1.16414
R1060 VTAIL.n623 VTAIL.n519 0.470328
R1061 VTAIL.n207 VTAIL.n103 0.470328
R1062 VTAIL.n784 VTAIL.n783 0.388379
R1063 VTAIL.n787 VTAIL.n750 0.388379
R1064 VTAIL.n830 VTAIL.n728 0.388379
R1065 VTAIL.n56 VTAIL.n55 0.388379
R1066 VTAIL.n59 VTAIL.n22 0.388379
R1067 VTAIL.n102 VTAIL.n0 0.388379
R1068 VTAIL.n160 VTAIL.n159 0.388379
R1069 VTAIL.n163 VTAIL.n126 0.388379
R1070 VTAIL.n206 VTAIL.n104 0.388379
R1071 VTAIL.n264 VTAIL.n263 0.388379
R1072 VTAIL.n267 VTAIL.n230 0.388379
R1073 VTAIL.n310 VTAIL.n208 0.388379
R1074 VTAIL.n726 VTAIL.n624 0.388379
R1075 VTAIL.n683 VTAIL.n646 0.388379
R1076 VTAIL.n680 VTAIL.n648 0.388379
R1077 VTAIL.n622 VTAIL.n520 0.388379
R1078 VTAIL.n579 VTAIL.n542 0.388379
R1079 VTAIL.n576 VTAIL.n544 0.388379
R1080 VTAIL.n518 VTAIL.n416 0.388379
R1081 VTAIL.n475 VTAIL.n438 0.388379
R1082 VTAIL.n472 VTAIL.n440 0.388379
R1083 VTAIL.n414 VTAIL.n312 0.388379
R1084 VTAIL.n371 VTAIL.n334 0.388379
R1085 VTAIL.n368 VTAIL.n336 0.388379
R1086 VTAIL.n767 VTAIL.n759 0.155672
R1087 VTAIL.n768 VTAIL.n767 0.155672
R1088 VTAIL.n768 VTAIL.n755 0.155672
R1089 VTAIL.n775 VTAIL.n755 0.155672
R1090 VTAIL.n776 VTAIL.n775 0.155672
R1091 VTAIL.n776 VTAIL.n751 0.155672
R1092 VTAIL.n785 VTAIL.n751 0.155672
R1093 VTAIL.n786 VTAIL.n785 0.155672
R1094 VTAIL.n786 VTAIL.n747 0.155672
R1095 VTAIL.n793 VTAIL.n747 0.155672
R1096 VTAIL.n794 VTAIL.n793 0.155672
R1097 VTAIL.n794 VTAIL.n743 0.155672
R1098 VTAIL.n801 VTAIL.n743 0.155672
R1099 VTAIL.n802 VTAIL.n801 0.155672
R1100 VTAIL.n802 VTAIL.n739 0.155672
R1101 VTAIL.n809 VTAIL.n739 0.155672
R1102 VTAIL.n810 VTAIL.n809 0.155672
R1103 VTAIL.n810 VTAIL.n735 0.155672
R1104 VTAIL.n817 VTAIL.n735 0.155672
R1105 VTAIL.n818 VTAIL.n817 0.155672
R1106 VTAIL.n818 VTAIL.n731 0.155672
R1107 VTAIL.n825 VTAIL.n731 0.155672
R1108 VTAIL.n826 VTAIL.n825 0.155672
R1109 VTAIL.n39 VTAIL.n31 0.155672
R1110 VTAIL.n40 VTAIL.n39 0.155672
R1111 VTAIL.n40 VTAIL.n27 0.155672
R1112 VTAIL.n47 VTAIL.n27 0.155672
R1113 VTAIL.n48 VTAIL.n47 0.155672
R1114 VTAIL.n48 VTAIL.n23 0.155672
R1115 VTAIL.n57 VTAIL.n23 0.155672
R1116 VTAIL.n58 VTAIL.n57 0.155672
R1117 VTAIL.n58 VTAIL.n19 0.155672
R1118 VTAIL.n65 VTAIL.n19 0.155672
R1119 VTAIL.n66 VTAIL.n65 0.155672
R1120 VTAIL.n66 VTAIL.n15 0.155672
R1121 VTAIL.n73 VTAIL.n15 0.155672
R1122 VTAIL.n74 VTAIL.n73 0.155672
R1123 VTAIL.n74 VTAIL.n11 0.155672
R1124 VTAIL.n81 VTAIL.n11 0.155672
R1125 VTAIL.n82 VTAIL.n81 0.155672
R1126 VTAIL.n82 VTAIL.n7 0.155672
R1127 VTAIL.n89 VTAIL.n7 0.155672
R1128 VTAIL.n90 VTAIL.n89 0.155672
R1129 VTAIL.n90 VTAIL.n3 0.155672
R1130 VTAIL.n97 VTAIL.n3 0.155672
R1131 VTAIL.n98 VTAIL.n97 0.155672
R1132 VTAIL.n143 VTAIL.n135 0.155672
R1133 VTAIL.n144 VTAIL.n143 0.155672
R1134 VTAIL.n144 VTAIL.n131 0.155672
R1135 VTAIL.n151 VTAIL.n131 0.155672
R1136 VTAIL.n152 VTAIL.n151 0.155672
R1137 VTAIL.n152 VTAIL.n127 0.155672
R1138 VTAIL.n161 VTAIL.n127 0.155672
R1139 VTAIL.n162 VTAIL.n161 0.155672
R1140 VTAIL.n162 VTAIL.n123 0.155672
R1141 VTAIL.n169 VTAIL.n123 0.155672
R1142 VTAIL.n170 VTAIL.n169 0.155672
R1143 VTAIL.n170 VTAIL.n119 0.155672
R1144 VTAIL.n177 VTAIL.n119 0.155672
R1145 VTAIL.n178 VTAIL.n177 0.155672
R1146 VTAIL.n178 VTAIL.n115 0.155672
R1147 VTAIL.n185 VTAIL.n115 0.155672
R1148 VTAIL.n186 VTAIL.n185 0.155672
R1149 VTAIL.n186 VTAIL.n111 0.155672
R1150 VTAIL.n193 VTAIL.n111 0.155672
R1151 VTAIL.n194 VTAIL.n193 0.155672
R1152 VTAIL.n194 VTAIL.n107 0.155672
R1153 VTAIL.n201 VTAIL.n107 0.155672
R1154 VTAIL.n202 VTAIL.n201 0.155672
R1155 VTAIL.n247 VTAIL.n239 0.155672
R1156 VTAIL.n248 VTAIL.n247 0.155672
R1157 VTAIL.n248 VTAIL.n235 0.155672
R1158 VTAIL.n255 VTAIL.n235 0.155672
R1159 VTAIL.n256 VTAIL.n255 0.155672
R1160 VTAIL.n256 VTAIL.n231 0.155672
R1161 VTAIL.n265 VTAIL.n231 0.155672
R1162 VTAIL.n266 VTAIL.n265 0.155672
R1163 VTAIL.n266 VTAIL.n227 0.155672
R1164 VTAIL.n273 VTAIL.n227 0.155672
R1165 VTAIL.n274 VTAIL.n273 0.155672
R1166 VTAIL.n274 VTAIL.n223 0.155672
R1167 VTAIL.n281 VTAIL.n223 0.155672
R1168 VTAIL.n282 VTAIL.n281 0.155672
R1169 VTAIL.n282 VTAIL.n219 0.155672
R1170 VTAIL.n289 VTAIL.n219 0.155672
R1171 VTAIL.n290 VTAIL.n289 0.155672
R1172 VTAIL.n290 VTAIL.n215 0.155672
R1173 VTAIL.n297 VTAIL.n215 0.155672
R1174 VTAIL.n298 VTAIL.n297 0.155672
R1175 VTAIL.n298 VTAIL.n211 0.155672
R1176 VTAIL.n305 VTAIL.n211 0.155672
R1177 VTAIL.n306 VTAIL.n305 0.155672
R1178 VTAIL.n722 VTAIL.n721 0.155672
R1179 VTAIL.n721 VTAIL.n627 0.155672
R1180 VTAIL.n714 VTAIL.n627 0.155672
R1181 VTAIL.n714 VTAIL.n713 0.155672
R1182 VTAIL.n713 VTAIL.n631 0.155672
R1183 VTAIL.n706 VTAIL.n631 0.155672
R1184 VTAIL.n706 VTAIL.n705 0.155672
R1185 VTAIL.n705 VTAIL.n635 0.155672
R1186 VTAIL.n698 VTAIL.n635 0.155672
R1187 VTAIL.n698 VTAIL.n697 0.155672
R1188 VTAIL.n697 VTAIL.n639 0.155672
R1189 VTAIL.n690 VTAIL.n639 0.155672
R1190 VTAIL.n690 VTAIL.n689 0.155672
R1191 VTAIL.n689 VTAIL.n643 0.155672
R1192 VTAIL.n682 VTAIL.n643 0.155672
R1193 VTAIL.n682 VTAIL.n681 0.155672
R1194 VTAIL.n681 VTAIL.n647 0.155672
R1195 VTAIL.n674 VTAIL.n647 0.155672
R1196 VTAIL.n674 VTAIL.n673 0.155672
R1197 VTAIL.n673 VTAIL.n653 0.155672
R1198 VTAIL.n666 VTAIL.n653 0.155672
R1199 VTAIL.n666 VTAIL.n665 0.155672
R1200 VTAIL.n665 VTAIL.n657 0.155672
R1201 VTAIL.n618 VTAIL.n617 0.155672
R1202 VTAIL.n617 VTAIL.n523 0.155672
R1203 VTAIL.n610 VTAIL.n523 0.155672
R1204 VTAIL.n610 VTAIL.n609 0.155672
R1205 VTAIL.n609 VTAIL.n527 0.155672
R1206 VTAIL.n602 VTAIL.n527 0.155672
R1207 VTAIL.n602 VTAIL.n601 0.155672
R1208 VTAIL.n601 VTAIL.n531 0.155672
R1209 VTAIL.n594 VTAIL.n531 0.155672
R1210 VTAIL.n594 VTAIL.n593 0.155672
R1211 VTAIL.n593 VTAIL.n535 0.155672
R1212 VTAIL.n586 VTAIL.n535 0.155672
R1213 VTAIL.n586 VTAIL.n585 0.155672
R1214 VTAIL.n585 VTAIL.n539 0.155672
R1215 VTAIL.n578 VTAIL.n539 0.155672
R1216 VTAIL.n578 VTAIL.n577 0.155672
R1217 VTAIL.n577 VTAIL.n543 0.155672
R1218 VTAIL.n570 VTAIL.n543 0.155672
R1219 VTAIL.n570 VTAIL.n569 0.155672
R1220 VTAIL.n569 VTAIL.n549 0.155672
R1221 VTAIL.n562 VTAIL.n549 0.155672
R1222 VTAIL.n562 VTAIL.n561 0.155672
R1223 VTAIL.n561 VTAIL.n553 0.155672
R1224 VTAIL.n514 VTAIL.n513 0.155672
R1225 VTAIL.n513 VTAIL.n419 0.155672
R1226 VTAIL.n506 VTAIL.n419 0.155672
R1227 VTAIL.n506 VTAIL.n505 0.155672
R1228 VTAIL.n505 VTAIL.n423 0.155672
R1229 VTAIL.n498 VTAIL.n423 0.155672
R1230 VTAIL.n498 VTAIL.n497 0.155672
R1231 VTAIL.n497 VTAIL.n427 0.155672
R1232 VTAIL.n490 VTAIL.n427 0.155672
R1233 VTAIL.n490 VTAIL.n489 0.155672
R1234 VTAIL.n489 VTAIL.n431 0.155672
R1235 VTAIL.n482 VTAIL.n431 0.155672
R1236 VTAIL.n482 VTAIL.n481 0.155672
R1237 VTAIL.n481 VTAIL.n435 0.155672
R1238 VTAIL.n474 VTAIL.n435 0.155672
R1239 VTAIL.n474 VTAIL.n473 0.155672
R1240 VTAIL.n473 VTAIL.n439 0.155672
R1241 VTAIL.n466 VTAIL.n439 0.155672
R1242 VTAIL.n466 VTAIL.n465 0.155672
R1243 VTAIL.n465 VTAIL.n445 0.155672
R1244 VTAIL.n458 VTAIL.n445 0.155672
R1245 VTAIL.n458 VTAIL.n457 0.155672
R1246 VTAIL.n457 VTAIL.n449 0.155672
R1247 VTAIL.n410 VTAIL.n409 0.155672
R1248 VTAIL.n409 VTAIL.n315 0.155672
R1249 VTAIL.n402 VTAIL.n315 0.155672
R1250 VTAIL.n402 VTAIL.n401 0.155672
R1251 VTAIL.n401 VTAIL.n319 0.155672
R1252 VTAIL.n394 VTAIL.n319 0.155672
R1253 VTAIL.n394 VTAIL.n393 0.155672
R1254 VTAIL.n393 VTAIL.n323 0.155672
R1255 VTAIL.n386 VTAIL.n323 0.155672
R1256 VTAIL.n386 VTAIL.n385 0.155672
R1257 VTAIL.n385 VTAIL.n327 0.155672
R1258 VTAIL.n378 VTAIL.n327 0.155672
R1259 VTAIL.n378 VTAIL.n377 0.155672
R1260 VTAIL.n377 VTAIL.n331 0.155672
R1261 VTAIL.n370 VTAIL.n331 0.155672
R1262 VTAIL.n370 VTAIL.n369 0.155672
R1263 VTAIL.n369 VTAIL.n335 0.155672
R1264 VTAIL.n362 VTAIL.n335 0.155672
R1265 VTAIL.n362 VTAIL.n361 0.155672
R1266 VTAIL.n361 VTAIL.n341 0.155672
R1267 VTAIL.n354 VTAIL.n341 0.155672
R1268 VTAIL.n354 VTAIL.n353 0.155672
R1269 VTAIL.n353 VTAIL.n345 0.155672
R1270 VP.n3 VP.t1 203.659
R1271 VP.n3 VP.t3 202.793
R1272 VP.n0 VP.t0 169.874
R1273 VP.n5 VP.t2 169.874
R1274 VP.n13 VP.n12 161.3
R1275 VP.n11 VP.n1 161.3
R1276 VP.n10 VP.n9 161.3
R1277 VP.n8 VP.n2 161.3
R1278 VP.n7 VP.n6 161.3
R1279 VP.n14 VP.n0 65.6537
R1280 VP.n5 VP.n4 65.6537
R1281 VP.n4 VP.n3 55.3724
R1282 VP.n10 VP.n2 40.577
R1283 VP.n11 VP.n10 40.577
R1284 VP.n6 VP.n5 24.5923
R1285 VP.n6 VP.n2 24.5923
R1286 VP.n12 VP.n11 24.5923
R1287 VP.n12 VP.n0 24.5923
R1288 VP.n7 VP.n4 0.354861
R1289 VP.n14 VP.n13 0.354861
R1290 VP VP.n14 0.267071
R1291 VP.n8 VP.n7 0.189894
R1292 VP.n9 VP.n8 0.189894
R1293 VP.n9 VP.n1 0.189894
R1294 VP.n13 VP.n1 0.189894
R1295 VDD1 VDD1.n1 120.576
R1296 VDD1 VDD1.n0 72.4111
R1297 VDD1.n0 VDD1.t2 1.72765
R1298 VDD1.n0 VDD1.t0 1.72765
R1299 VDD1.n1 VDD1.t1 1.72765
R1300 VDD1.n1 VDD1.t3 1.72765
R1301 B.n462 B.n125 585
R1302 B.n461 B.n460 585
R1303 B.n459 B.n126 585
R1304 B.n458 B.n457 585
R1305 B.n456 B.n127 585
R1306 B.n455 B.n454 585
R1307 B.n453 B.n128 585
R1308 B.n452 B.n451 585
R1309 B.n450 B.n129 585
R1310 B.n449 B.n448 585
R1311 B.n447 B.n130 585
R1312 B.n446 B.n445 585
R1313 B.n444 B.n131 585
R1314 B.n443 B.n442 585
R1315 B.n441 B.n132 585
R1316 B.n440 B.n439 585
R1317 B.n438 B.n133 585
R1318 B.n437 B.n436 585
R1319 B.n435 B.n134 585
R1320 B.n434 B.n433 585
R1321 B.n432 B.n135 585
R1322 B.n431 B.n430 585
R1323 B.n429 B.n136 585
R1324 B.n428 B.n427 585
R1325 B.n426 B.n137 585
R1326 B.n425 B.n424 585
R1327 B.n423 B.n138 585
R1328 B.n422 B.n421 585
R1329 B.n420 B.n139 585
R1330 B.n419 B.n418 585
R1331 B.n417 B.n140 585
R1332 B.n416 B.n415 585
R1333 B.n414 B.n141 585
R1334 B.n413 B.n412 585
R1335 B.n411 B.n142 585
R1336 B.n410 B.n409 585
R1337 B.n408 B.n143 585
R1338 B.n407 B.n406 585
R1339 B.n405 B.n144 585
R1340 B.n404 B.n403 585
R1341 B.n402 B.n145 585
R1342 B.n401 B.n400 585
R1343 B.n399 B.n146 585
R1344 B.n398 B.n397 585
R1345 B.n396 B.n147 585
R1346 B.n395 B.n394 585
R1347 B.n393 B.n148 585
R1348 B.n392 B.n391 585
R1349 B.n390 B.n149 585
R1350 B.n389 B.n388 585
R1351 B.n387 B.n150 585
R1352 B.n386 B.n385 585
R1353 B.n384 B.n151 585
R1354 B.n383 B.n382 585
R1355 B.n381 B.n152 585
R1356 B.n380 B.n379 585
R1357 B.n378 B.n153 585
R1358 B.n377 B.n376 585
R1359 B.n375 B.n154 585
R1360 B.n374 B.n373 585
R1361 B.n372 B.n155 585
R1362 B.n371 B.n370 585
R1363 B.n369 B.n368 585
R1364 B.n367 B.n159 585
R1365 B.n366 B.n365 585
R1366 B.n364 B.n160 585
R1367 B.n363 B.n362 585
R1368 B.n361 B.n161 585
R1369 B.n360 B.n359 585
R1370 B.n358 B.n162 585
R1371 B.n357 B.n356 585
R1372 B.n354 B.n163 585
R1373 B.n353 B.n352 585
R1374 B.n351 B.n166 585
R1375 B.n350 B.n349 585
R1376 B.n348 B.n167 585
R1377 B.n347 B.n346 585
R1378 B.n345 B.n168 585
R1379 B.n344 B.n343 585
R1380 B.n342 B.n169 585
R1381 B.n341 B.n340 585
R1382 B.n339 B.n170 585
R1383 B.n338 B.n337 585
R1384 B.n336 B.n171 585
R1385 B.n335 B.n334 585
R1386 B.n333 B.n172 585
R1387 B.n332 B.n331 585
R1388 B.n330 B.n173 585
R1389 B.n329 B.n328 585
R1390 B.n327 B.n174 585
R1391 B.n326 B.n325 585
R1392 B.n324 B.n175 585
R1393 B.n323 B.n322 585
R1394 B.n321 B.n176 585
R1395 B.n320 B.n319 585
R1396 B.n318 B.n177 585
R1397 B.n317 B.n316 585
R1398 B.n315 B.n178 585
R1399 B.n314 B.n313 585
R1400 B.n312 B.n179 585
R1401 B.n311 B.n310 585
R1402 B.n309 B.n180 585
R1403 B.n308 B.n307 585
R1404 B.n306 B.n181 585
R1405 B.n305 B.n304 585
R1406 B.n303 B.n182 585
R1407 B.n302 B.n301 585
R1408 B.n300 B.n183 585
R1409 B.n299 B.n298 585
R1410 B.n297 B.n184 585
R1411 B.n296 B.n295 585
R1412 B.n294 B.n185 585
R1413 B.n293 B.n292 585
R1414 B.n291 B.n186 585
R1415 B.n290 B.n289 585
R1416 B.n288 B.n187 585
R1417 B.n287 B.n286 585
R1418 B.n285 B.n188 585
R1419 B.n284 B.n283 585
R1420 B.n282 B.n189 585
R1421 B.n281 B.n280 585
R1422 B.n279 B.n190 585
R1423 B.n278 B.n277 585
R1424 B.n276 B.n191 585
R1425 B.n275 B.n274 585
R1426 B.n273 B.n192 585
R1427 B.n272 B.n271 585
R1428 B.n270 B.n193 585
R1429 B.n269 B.n268 585
R1430 B.n267 B.n194 585
R1431 B.n266 B.n265 585
R1432 B.n264 B.n195 585
R1433 B.n263 B.n262 585
R1434 B.n464 B.n463 585
R1435 B.n465 B.n124 585
R1436 B.n467 B.n466 585
R1437 B.n468 B.n123 585
R1438 B.n470 B.n469 585
R1439 B.n471 B.n122 585
R1440 B.n473 B.n472 585
R1441 B.n474 B.n121 585
R1442 B.n476 B.n475 585
R1443 B.n477 B.n120 585
R1444 B.n479 B.n478 585
R1445 B.n480 B.n119 585
R1446 B.n482 B.n481 585
R1447 B.n483 B.n118 585
R1448 B.n485 B.n484 585
R1449 B.n486 B.n117 585
R1450 B.n488 B.n487 585
R1451 B.n489 B.n116 585
R1452 B.n491 B.n490 585
R1453 B.n492 B.n115 585
R1454 B.n494 B.n493 585
R1455 B.n495 B.n114 585
R1456 B.n497 B.n496 585
R1457 B.n498 B.n113 585
R1458 B.n500 B.n499 585
R1459 B.n501 B.n112 585
R1460 B.n503 B.n502 585
R1461 B.n504 B.n111 585
R1462 B.n506 B.n505 585
R1463 B.n507 B.n110 585
R1464 B.n509 B.n508 585
R1465 B.n510 B.n109 585
R1466 B.n512 B.n511 585
R1467 B.n513 B.n108 585
R1468 B.n515 B.n514 585
R1469 B.n516 B.n107 585
R1470 B.n518 B.n517 585
R1471 B.n519 B.n106 585
R1472 B.n521 B.n520 585
R1473 B.n522 B.n105 585
R1474 B.n524 B.n523 585
R1475 B.n525 B.n104 585
R1476 B.n527 B.n526 585
R1477 B.n528 B.n103 585
R1478 B.n530 B.n529 585
R1479 B.n531 B.n102 585
R1480 B.n533 B.n532 585
R1481 B.n534 B.n101 585
R1482 B.n536 B.n535 585
R1483 B.n537 B.n100 585
R1484 B.n539 B.n538 585
R1485 B.n540 B.n99 585
R1486 B.n542 B.n541 585
R1487 B.n543 B.n98 585
R1488 B.n545 B.n544 585
R1489 B.n546 B.n97 585
R1490 B.n548 B.n547 585
R1491 B.n549 B.n96 585
R1492 B.n551 B.n550 585
R1493 B.n552 B.n95 585
R1494 B.n554 B.n553 585
R1495 B.n555 B.n94 585
R1496 B.n557 B.n556 585
R1497 B.n558 B.n93 585
R1498 B.n560 B.n559 585
R1499 B.n561 B.n92 585
R1500 B.n563 B.n562 585
R1501 B.n564 B.n91 585
R1502 B.n566 B.n565 585
R1503 B.n567 B.n90 585
R1504 B.n768 B.n19 585
R1505 B.n767 B.n766 585
R1506 B.n765 B.n20 585
R1507 B.n764 B.n763 585
R1508 B.n762 B.n21 585
R1509 B.n761 B.n760 585
R1510 B.n759 B.n22 585
R1511 B.n758 B.n757 585
R1512 B.n756 B.n23 585
R1513 B.n755 B.n754 585
R1514 B.n753 B.n24 585
R1515 B.n752 B.n751 585
R1516 B.n750 B.n25 585
R1517 B.n749 B.n748 585
R1518 B.n747 B.n26 585
R1519 B.n746 B.n745 585
R1520 B.n744 B.n27 585
R1521 B.n743 B.n742 585
R1522 B.n741 B.n28 585
R1523 B.n740 B.n739 585
R1524 B.n738 B.n29 585
R1525 B.n737 B.n736 585
R1526 B.n735 B.n30 585
R1527 B.n734 B.n733 585
R1528 B.n732 B.n31 585
R1529 B.n731 B.n730 585
R1530 B.n729 B.n32 585
R1531 B.n728 B.n727 585
R1532 B.n726 B.n33 585
R1533 B.n725 B.n724 585
R1534 B.n723 B.n34 585
R1535 B.n722 B.n721 585
R1536 B.n720 B.n35 585
R1537 B.n719 B.n718 585
R1538 B.n717 B.n36 585
R1539 B.n716 B.n715 585
R1540 B.n714 B.n37 585
R1541 B.n713 B.n712 585
R1542 B.n711 B.n38 585
R1543 B.n710 B.n709 585
R1544 B.n708 B.n39 585
R1545 B.n707 B.n706 585
R1546 B.n705 B.n40 585
R1547 B.n704 B.n703 585
R1548 B.n702 B.n41 585
R1549 B.n701 B.n700 585
R1550 B.n699 B.n42 585
R1551 B.n698 B.n697 585
R1552 B.n696 B.n43 585
R1553 B.n695 B.n694 585
R1554 B.n693 B.n44 585
R1555 B.n692 B.n691 585
R1556 B.n690 B.n45 585
R1557 B.n689 B.n688 585
R1558 B.n687 B.n46 585
R1559 B.n686 B.n685 585
R1560 B.n684 B.n47 585
R1561 B.n683 B.n682 585
R1562 B.n681 B.n48 585
R1563 B.n680 B.n679 585
R1564 B.n678 B.n49 585
R1565 B.n677 B.n676 585
R1566 B.n675 B.n674 585
R1567 B.n673 B.n53 585
R1568 B.n672 B.n671 585
R1569 B.n670 B.n54 585
R1570 B.n669 B.n668 585
R1571 B.n667 B.n55 585
R1572 B.n666 B.n665 585
R1573 B.n664 B.n56 585
R1574 B.n663 B.n662 585
R1575 B.n660 B.n57 585
R1576 B.n659 B.n658 585
R1577 B.n657 B.n60 585
R1578 B.n656 B.n655 585
R1579 B.n654 B.n61 585
R1580 B.n653 B.n652 585
R1581 B.n651 B.n62 585
R1582 B.n650 B.n649 585
R1583 B.n648 B.n63 585
R1584 B.n647 B.n646 585
R1585 B.n645 B.n64 585
R1586 B.n644 B.n643 585
R1587 B.n642 B.n65 585
R1588 B.n641 B.n640 585
R1589 B.n639 B.n66 585
R1590 B.n638 B.n637 585
R1591 B.n636 B.n67 585
R1592 B.n635 B.n634 585
R1593 B.n633 B.n68 585
R1594 B.n632 B.n631 585
R1595 B.n630 B.n69 585
R1596 B.n629 B.n628 585
R1597 B.n627 B.n70 585
R1598 B.n626 B.n625 585
R1599 B.n624 B.n71 585
R1600 B.n623 B.n622 585
R1601 B.n621 B.n72 585
R1602 B.n620 B.n619 585
R1603 B.n618 B.n73 585
R1604 B.n617 B.n616 585
R1605 B.n615 B.n74 585
R1606 B.n614 B.n613 585
R1607 B.n612 B.n75 585
R1608 B.n611 B.n610 585
R1609 B.n609 B.n76 585
R1610 B.n608 B.n607 585
R1611 B.n606 B.n77 585
R1612 B.n605 B.n604 585
R1613 B.n603 B.n78 585
R1614 B.n602 B.n601 585
R1615 B.n600 B.n79 585
R1616 B.n599 B.n598 585
R1617 B.n597 B.n80 585
R1618 B.n596 B.n595 585
R1619 B.n594 B.n81 585
R1620 B.n593 B.n592 585
R1621 B.n591 B.n82 585
R1622 B.n590 B.n589 585
R1623 B.n588 B.n83 585
R1624 B.n587 B.n586 585
R1625 B.n585 B.n84 585
R1626 B.n584 B.n583 585
R1627 B.n582 B.n85 585
R1628 B.n581 B.n580 585
R1629 B.n579 B.n86 585
R1630 B.n578 B.n577 585
R1631 B.n576 B.n87 585
R1632 B.n575 B.n574 585
R1633 B.n573 B.n88 585
R1634 B.n572 B.n571 585
R1635 B.n570 B.n89 585
R1636 B.n569 B.n568 585
R1637 B.n770 B.n769 585
R1638 B.n771 B.n18 585
R1639 B.n773 B.n772 585
R1640 B.n774 B.n17 585
R1641 B.n776 B.n775 585
R1642 B.n777 B.n16 585
R1643 B.n779 B.n778 585
R1644 B.n780 B.n15 585
R1645 B.n782 B.n781 585
R1646 B.n783 B.n14 585
R1647 B.n785 B.n784 585
R1648 B.n786 B.n13 585
R1649 B.n788 B.n787 585
R1650 B.n789 B.n12 585
R1651 B.n791 B.n790 585
R1652 B.n792 B.n11 585
R1653 B.n794 B.n793 585
R1654 B.n795 B.n10 585
R1655 B.n797 B.n796 585
R1656 B.n798 B.n9 585
R1657 B.n800 B.n799 585
R1658 B.n801 B.n8 585
R1659 B.n803 B.n802 585
R1660 B.n804 B.n7 585
R1661 B.n806 B.n805 585
R1662 B.n807 B.n6 585
R1663 B.n809 B.n808 585
R1664 B.n810 B.n5 585
R1665 B.n812 B.n811 585
R1666 B.n813 B.n4 585
R1667 B.n815 B.n814 585
R1668 B.n816 B.n3 585
R1669 B.n818 B.n817 585
R1670 B.n819 B.n0 585
R1671 B.n2 B.n1 585
R1672 B.n213 B.n212 585
R1673 B.n215 B.n214 585
R1674 B.n216 B.n211 585
R1675 B.n218 B.n217 585
R1676 B.n219 B.n210 585
R1677 B.n221 B.n220 585
R1678 B.n222 B.n209 585
R1679 B.n224 B.n223 585
R1680 B.n225 B.n208 585
R1681 B.n227 B.n226 585
R1682 B.n228 B.n207 585
R1683 B.n230 B.n229 585
R1684 B.n231 B.n206 585
R1685 B.n233 B.n232 585
R1686 B.n234 B.n205 585
R1687 B.n236 B.n235 585
R1688 B.n237 B.n204 585
R1689 B.n239 B.n238 585
R1690 B.n240 B.n203 585
R1691 B.n242 B.n241 585
R1692 B.n243 B.n202 585
R1693 B.n245 B.n244 585
R1694 B.n246 B.n201 585
R1695 B.n248 B.n247 585
R1696 B.n249 B.n200 585
R1697 B.n251 B.n250 585
R1698 B.n252 B.n199 585
R1699 B.n254 B.n253 585
R1700 B.n255 B.n198 585
R1701 B.n257 B.n256 585
R1702 B.n258 B.n197 585
R1703 B.n260 B.n259 585
R1704 B.n261 B.n196 585
R1705 B.n156 B.t4 556.58
R1706 B.n58 B.t2 556.58
R1707 B.n164 B.t10 556.58
R1708 B.n50 B.t8 556.58
R1709 B.n262 B.n261 506.916
R1710 B.n464 B.n125 506.916
R1711 B.n568 B.n567 506.916
R1712 B.n770 B.n19 506.916
R1713 B.n157 B.t5 498.397
R1714 B.n59 B.t1 498.397
R1715 B.n165 B.t11 498.397
R1716 B.n51 B.t7 498.397
R1717 B.n164 B.t9 378.024
R1718 B.n156 B.t3 378.024
R1719 B.n58 B.t0 378.024
R1720 B.n50 B.t6 378.024
R1721 B.n821 B.n820 256.663
R1722 B.n820 B.n819 235.042
R1723 B.n820 B.n2 235.042
R1724 B.n262 B.n195 163.367
R1725 B.n266 B.n195 163.367
R1726 B.n267 B.n266 163.367
R1727 B.n268 B.n267 163.367
R1728 B.n268 B.n193 163.367
R1729 B.n272 B.n193 163.367
R1730 B.n273 B.n272 163.367
R1731 B.n274 B.n273 163.367
R1732 B.n274 B.n191 163.367
R1733 B.n278 B.n191 163.367
R1734 B.n279 B.n278 163.367
R1735 B.n280 B.n279 163.367
R1736 B.n280 B.n189 163.367
R1737 B.n284 B.n189 163.367
R1738 B.n285 B.n284 163.367
R1739 B.n286 B.n285 163.367
R1740 B.n286 B.n187 163.367
R1741 B.n290 B.n187 163.367
R1742 B.n291 B.n290 163.367
R1743 B.n292 B.n291 163.367
R1744 B.n292 B.n185 163.367
R1745 B.n296 B.n185 163.367
R1746 B.n297 B.n296 163.367
R1747 B.n298 B.n297 163.367
R1748 B.n298 B.n183 163.367
R1749 B.n302 B.n183 163.367
R1750 B.n303 B.n302 163.367
R1751 B.n304 B.n303 163.367
R1752 B.n304 B.n181 163.367
R1753 B.n308 B.n181 163.367
R1754 B.n309 B.n308 163.367
R1755 B.n310 B.n309 163.367
R1756 B.n310 B.n179 163.367
R1757 B.n314 B.n179 163.367
R1758 B.n315 B.n314 163.367
R1759 B.n316 B.n315 163.367
R1760 B.n316 B.n177 163.367
R1761 B.n320 B.n177 163.367
R1762 B.n321 B.n320 163.367
R1763 B.n322 B.n321 163.367
R1764 B.n322 B.n175 163.367
R1765 B.n326 B.n175 163.367
R1766 B.n327 B.n326 163.367
R1767 B.n328 B.n327 163.367
R1768 B.n328 B.n173 163.367
R1769 B.n332 B.n173 163.367
R1770 B.n333 B.n332 163.367
R1771 B.n334 B.n333 163.367
R1772 B.n334 B.n171 163.367
R1773 B.n338 B.n171 163.367
R1774 B.n339 B.n338 163.367
R1775 B.n340 B.n339 163.367
R1776 B.n340 B.n169 163.367
R1777 B.n344 B.n169 163.367
R1778 B.n345 B.n344 163.367
R1779 B.n346 B.n345 163.367
R1780 B.n346 B.n167 163.367
R1781 B.n350 B.n167 163.367
R1782 B.n351 B.n350 163.367
R1783 B.n352 B.n351 163.367
R1784 B.n352 B.n163 163.367
R1785 B.n357 B.n163 163.367
R1786 B.n358 B.n357 163.367
R1787 B.n359 B.n358 163.367
R1788 B.n359 B.n161 163.367
R1789 B.n363 B.n161 163.367
R1790 B.n364 B.n363 163.367
R1791 B.n365 B.n364 163.367
R1792 B.n365 B.n159 163.367
R1793 B.n369 B.n159 163.367
R1794 B.n370 B.n369 163.367
R1795 B.n370 B.n155 163.367
R1796 B.n374 B.n155 163.367
R1797 B.n375 B.n374 163.367
R1798 B.n376 B.n375 163.367
R1799 B.n376 B.n153 163.367
R1800 B.n380 B.n153 163.367
R1801 B.n381 B.n380 163.367
R1802 B.n382 B.n381 163.367
R1803 B.n382 B.n151 163.367
R1804 B.n386 B.n151 163.367
R1805 B.n387 B.n386 163.367
R1806 B.n388 B.n387 163.367
R1807 B.n388 B.n149 163.367
R1808 B.n392 B.n149 163.367
R1809 B.n393 B.n392 163.367
R1810 B.n394 B.n393 163.367
R1811 B.n394 B.n147 163.367
R1812 B.n398 B.n147 163.367
R1813 B.n399 B.n398 163.367
R1814 B.n400 B.n399 163.367
R1815 B.n400 B.n145 163.367
R1816 B.n404 B.n145 163.367
R1817 B.n405 B.n404 163.367
R1818 B.n406 B.n405 163.367
R1819 B.n406 B.n143 163.367
R1820 B.n410 B.n143 163.367
R1821 B.n411 B.n410 163.367
R1822 B.n412 B.n411 163.367
R1823 B.n412 B.n141 163.367
R1824 B.n416 B.n141 163.367
R1825 B.n417 B.n416 163.367
R1826 B.n418 B.n417 163.367
R1827 B.n418 B.n139 163.367
R1828 B.n422 B.n139 163.367
R1829 B.n423 B.n422 163.367
R1830 B.n424 B.n423 163.367
R1831 B.n424 B.n137 163.367
R1832 B.n428 B.n137 163.367
R1833 B.n429 B.n428 163.367
R1834 B.n430 B.n429 163.367
R1835 B.n430 B.n135 163.367
R1836 B.n434 B.n135 163.367
R1837 B.n435 B.n434 163.367
R1838 B.n436 B.n435 163.367
R1839 B.n436 B.n133 163.367
R1840 B.n440 B.n133 163.367
R1841 B.n441 B.n440 163.367
R1842 B.n442 B.n441 163.367
R1843 B.n442 B.n131 163.367
R1844 B.n446 B.n131 163.367
R1845 B.n447 B.n446 163.367
R1846 B.n448 B.n447 163.367
R1847 B.n448 B.n129 163.367
R1848 B.n452 B.n129 163.367
R1849 B.n453 B.n452 163.367
R1850 B.n454 B.n453 163.367
R1851 B.n454 B.n127 163.367
R1852 B.n458 B.n127 163.367
R1853 B.n459 B.n458 163.367
R1854 B.n460 B.n459 163.367
R1855 B.n460 B.n125 163.367
R1856 B.n567 B.n566 163.367
R1857 B.n566 B.n91 163.367
R1858 B.n562 B.n91 163.367
R1859 B.n562 B.n561 163.367
R1860 B.n561 B.n560 163.367
R1861 B.n560 B.n93 163.367
R1862 B.n556 B.n93 163.367
R1863 B.n556 B.n555 163.367
R1864 B.n555 B.n554 163.367
R1865 B.n554 B.n95 163.367
R1866 B.n550 B.n95 163.367
R1867 B.n550 B.n549 163.367
R1868 B.n549 B.n548 163.367
R1869 B.n548 B.n97 163.367
R1870 B.n544 B.n97 163.367
R1871 B.n544 B.n543 163.367
R1872 B.n543 B.n542 163.367
R1873 B.n542 B.n99 163.367
R1874 B.n538 B.n99 163.367
R1875 B.n538 B.n537 163.367
R1876 B.n537 B.n536 163.367
R1877 B.n536 B.n101 163.367
R1878 B.n532 B.n101 163.367
R1879 B.n532 B.n531 163.367
R1880 B.n531 B.n530 163.367
R1881 B.n530 B.n103 163.367
R1882 B.n526 B.n103 163.367
R1883 B.n526 B.n525 163.367
R1884 B.n525 B.n524 163.367
R1885 B.n524 B.n105 163.367
R1886 B.n520 B.n105 163.367
R1887 B.n520 B.n519 163.367
R1888 B.n519 B.n518 163.367
R1889 B.n518 B.n107 163.367
R1890 B.n514 B.n107 163.367
R1891 B.n514 B.n513 163.367
R1892 B.n513 B.n512 163.367
R1893 B.n512 B.n109 163.367
R1894 B.n508 B.n109 163.367
R1895 B.n508 B.n507 163.367
R1896 B.n507 B.n506 163.367
R1897 B.n506 B.n111 163.367
R1898 B.n502 B.n111 163.367
R1899 B.n502 B.n501 163.367
R1900 B.n501 B.n500 163.367
R1901 B.n500 B.n113 163.367
R1902 B.n496 B.n113 163.367
R1903 B.n496 B.n495 163.367
R1904 B.n495 B.n494 163.367
R1905 B.n494 B.n115 163.367
R1906 B.n490 B.n115 163.367
R1907 B.n490 B.n489 163.367
R1908 B.n489 B.n488 163.367
R1909 B.n488 B.n117 163.367
R1910 B.n484 B.n117 163.367
R1911 B.n484 B.n483 163.367
R1912 B.n483 B.n482 163.367
R1913 B.n482 B.n119 163.367
R1914 B.n478 B.n119 163.367
R1915 B.n478 B.n477 163.367
R1916 B.n477 B.n476 163.367
R1917 B.n476 B.n121 163.367
R1918 B.n472 B.n121 163.367
R1919 B.n472 B.n471 163.367
R1920 B.n471 B.n470 163.367
R1921 B.n470 B.n123 163.367
R1922 B.n466 B.n123 163.367
R1923 B.n466 B.n465 163.367
R1924 B.n465 B.n464 163.367
R1925 B.n766 B.n19 163.367
R1926 B.n766 B.n765 163.367
R1927 B.n765 B.n764 163.367
R1928 B.n764 B.n21 163.367
R1929 B.n760 B.n21 163.367
R1930 B.n760 B.n759 163.367
R1931 B.n759 B.n758 163.367
R1932 B.n758 B.n23 163.367
R1933 B.n754 B.n23 163.367
R1934 B.n754 B.n753 163.367
R1935 B.n753 B.n752 163.367
R1936 B.n752 B.n25 163.367
R1937 B.n748 B.n25 163.367
R1938 B.n748 B.n747 163.367
R1939 B.n747 B.n746 163.367
R1940 B.n746 B.n27 163.367
R1941 B.n742 B.n27 163.367
R1942 B.n742 B.n741 163.367
R1943 B.n741 B.n740 163.367
R1944 B.n740 B.n29 163.367
R1945 B.n736 B.n29 163.367
R1946 B.n736 B.n735 163.367
R1947 B.n735 B.n734 163.367
R1948 B.n734 B.n31 163.367
R1949 B.n730 B.n31 163.367
R1950 B.n730 B.n729 163.367
R1951 B.n729 B.n728 163.367
R1952 B.n728 B.n33 163.367
R1953 B.n724 B.n33 163.367
R1954 B.n724 B.n723 163.367
R1955 B.n723 B.n722 163.367
R1956 B.n722 B.n35 163.367
R1957 B.n718 B.n35 163.367
R1958 B.n718 B.n717 163.367
R1959 B.n717 B.n716 163.367
R1960 B.n716 B.n37 163.367
R1961 B.n712 B.n37 163.367
R1962 B.n712 B.n711 163.367
R1963 B.n711 B.n710 163.367
R1964 B.n710 B.n39 163.367
R1965 B.n706 B.n39 163.367
R1966 B.n706 B.n705 163.367
R1967 B.n705 B.n704 163.367
R1968 B.n704 B.n41 163.367
R1969 B.n700 B.n41 163.367
R1970 B.n700 B.n699 163.367
R1971 B.n699 B.n698 163.367
R1972 B.n698 B.n43 163.367
R1973 B.n694 B.n43 163.367
R1974 B.n694 B.n693 163.367
R1975 B.n693 B.n692 163.367
R1976 B.n692 B.n45 163.367
R1977 B.n688 B.n45 163.367
R1978 B.n688 B.n687 163.367
R1979 B.n687 B.n686 163.367
R1980 B.n686 B.n47 163.367
R1981 B.n682 B.n47 163.367
R1982 B.n682 B.n681 163.367
R1983 B.n681 B.n680 163.367
R1984 B.n680 B.n49 163.367
R1985 B.n676 B.n49 163.367
R1986 B.n676 B.n675 163.367
R1987 B.n675 B.n53 163.367
R1988 B.n671 B.n53 163.367
R1989 B.n671 B.n670 163.367
R1990 B.n670 B.n669 163.367
R1991 B.n669 B.n55 163.367
R1992 B.n665 B.n55 163.367
R1993 B.n665 B.n664 163.367
R1994 B.n664 B.n663 163.367
R1995 B.n663 B.n57 163.367
R1996 B.n658 B.n57 163.367
R1997 B.n658 B.n657 163.367
R1998 B.n657 B.n656 163.367
R1999 B.n656 B.n61 163.367
R2000 B.n652 B.n61 163.367
R2001 B.n652 B.n651 163.367
R2002 B.n651 B.n650 163.367
R2003 B.n650 B.n63 163.367
R2004 B.n646 B.n63 163.367
R2005 B.n646 B.n645 163.367
R2006 B.n645 B.n644 163.367
R2007 B.n644 B.n65 163.367
R2008 B.n640 B.n65 163.367
R2009 B.n640 B.n639 163.367
R2010 B.n639 B.n638 163.367
R2011 B.n638 B.n67 163.367
R2012 B.n634 B.n67 163.367
R2013 B.n634 B.n633 163.367
R2014 B.n633 B.n632 163.367
R2015 B.n632 B.n69 163.367
R2016 B.n628 B.n69 163.367
R2017 B.n628 B.n627 163.367
R2018 B.n627 B.n626 163.367
R2019 B.n626 B.n71 163.367
R2020 B.n622 B.n71 163.367
R2021 B.n622 B.n621 163.367
R2022 B.n621 B.n620 163.367
R2023 B.n620 B.n73 163.367
R2024 B.n616 B.n73 163.367
R2025 B.n616 B.n615 163.367
R2026 B.n615 B.n614 163.367
R2027 B.n614 B.n75 163.367
R2028 B.n610 B.n75 163.367
R2029 B.n610 B.n609 163.367
R2030 B.n609 B.n608 163.367
R2031 B.n608 B.n77 163.367
R2032 B.n604 B.n77 163.367
R2033 B.n604 B.n603 163.367
R2034 B.n603 B.n602 163.367
R2035 B.n602 B.n79 163.367
R2036 B.n598 B.n79 163.367
R2037 B.n598 B.n597 163.367
R2038 B.n597 B.n596 163.367
R2039 B.n596 B.n81 163.367
R2040 B.n592 B.n81 163.367
R2041 B.n592 B.n591 163.367
R2042 B.n591 B.n590 163.367
R2043 B.n590 B.n83 163.367
R2044 B.n586 B.n83 163.367
R2045 B.n586 B.n585 163.367
R2046 B.n585 B.n584 163.367
R2047 B.n584 B.n85 163.367
R2048 B.n580 B.n85 163.367
R2049 B.n580 B.n579 163.367
R2050 B.n579 B.n578 163.367
R2051 B.n578 B.n87 163.367
R2052 B.n574 B.n87 163.367
R2053 B.n574 B.n573 163.367
R2054 B.n573 B.n572 163.367
R2055 B.n572 B.n89 163.367
R2056 B.n568 B.n89 163.367
R2057 B.n771 B.n770 163.367
R2058 B.n772 B.n771 163.367
R2059 B.n772 B.n17 163.367
R2060 B.n776 B.n17 163.367
R2061 B.n777 B.n776 163.367
R2062 B.n778 B.n777 163.367
R2063 B.n778 B.n15 163.367
R2064 B.n782 B.n15 163.367
R2065 B.n783 B.n782 163.367
R2066 B.n784 B.n783 163.367
R2067 B.n784 B.n13 163.367
R2068 B.n788 B.n13 163.367
R2069 B.n789 B.n788 163.367
R2070 B.n790 B.n789 163.367
R2071 B.n790 B.n11 163.367
R2072 B.n794 B.n11 163.367
R2073 B.n795 B.n794 163.367
R2074 B.n796 B.n795 163.367
R2075 B.n796 B.n9 163.367
R2076 B.n800 B.n9 163.367
R2077 B.n801 B.n800 163.367
R2078 B.n802 B.n801 163.367
R2079 B.n802 B.n7 163.367
R2080 B.n806 B.n7 163.367
R2081 B.n807 B.n806 163.367
R2082 B.n808 B.n807 163.367
R2083 B.n808 B.n5 163.367
R2084 B.n812 B.n5 163.367
R2085 B.n813 B.n812 163.367
R2086 B.n814 B.n813 163.367
R2087 B.n814 B.n3 163.367
R2088 B.n818 B.n3 163.367
R2089 B.n819 B.n818 163.367
R2090 B.n213 B.n2 163.367
R2091 B.n214 B.n213 163.367
R2092 B.n214 B.n211 163.367
R2093 B.n218 B.n211 163.367
R2094 B.n219 B.n218 163.367
R2095 B.n220 B.n219 163.367
R2096 B.n220 B.n209 163.367
R2097 B.n224 B.n209 163.367
R2098 B.n225 B.n224 163.367
R2099 B.n226 B.n225 163.367
R2100 B.n226 B.n207 163.367
R2101 B.n230 B.n207 163.367
R2102 B.n231 B.n230 163.367
R2103 B.n232 B.n231 163.367
R2104 B.n232 B.n205 163.367
R2105 B.n236 B.n205 163.367
R2106 B.n237 B.n236 163.367
R2107 B.n238 B.n237 163.367
R2108 B.n238 B.n203 163.367
R2109 B.n242 B.n203 163.367
R2110 B.n243 B.n242 163.367
R2111 B.n244 B.n243 163.367
R2112 B.n244 B.n201 163.367
R2113 B.n248 B.n201 163.367
R2114 B.n249 B.n248 163.367
R2115 B.n250 B.n249 163.367
R2116 B.n250 B.n199 163.367
R2117 B.n254 B.n199 163.367
R2118 B.n255 B.n254 163.367
R2119 B.n256 B.n255 163.367
R2120 B.n256 B.n197 163.367
R2121 B.n260 B.n197 163.367
R2122 B.n261 B.n260 163.367
R2123 B.n355 B.n165 59.5399
R2124 B.n158 B.n157 59.5399
R2125 B.n661 B.n59 59.5399
R2126 B.n52 B.n51 59.5399
R2127 B.n165 B.n164 58.1823
R2128 B.n157 B.n156 58.1823
R2129 B.n59 B.n58 58.1823
R2130 B.n51 B.n50 58.1823
R2131 B.n769 B.n768 32.9371
R2132 B.n569 B.n90 32.9371
R2133 B.n463 B.n462 32.9371
R2134 B.n263 B.n196 32.9371
R2135 B B.n821 18.0485
R2136 B.n769 B.n18 10.6151
R2137 B.n773 B.n18 10.6151
R2138 B.n774 B.n773 10.6151
R2139 B.n775 B.n774 10.6151
R2140 B.n775 B.n16 10.6151
R2141 B.n779 B.n16 10.6151
R2142 B.n780 B.n779 10.6151
R2143 B.n781 B.n780 10.6151
R2144 B.n781 B.n14 10.6151
R2145 B.n785 B.n14 10.6151
R2146 B.n786 B.n785 10.6151
R2147 B.n787 B.n786 10.6151
R2148 B.n787 B.n12 10.6151
R2149 B.n791 B.n12 10.6151
R2150 B.n792 B.n791 10.6151
R2151 B.n793 B.n792 10.6151
R2152 B.n793 B.n10 10.6151
R2153 B.n797 B.n10 10.6151
R2154 B.n798 B.n797 10.6151
R2155 B.n799 B.n798 10.6151
R2156 B.n799 B.n8 10.6151
R2157 B.n803 B.n8 10.6151
R2158 B.n804 B.n803 10.6151
R2159 B.n805 B.n804 10.6151
R2160 B.n805 B.n6 10.6151
R2161 B.n809 B.n6 10.6151
R2162 B.n810 B.n809 10.6151
R2163 B.n811 B.n810 10.6151
R2164 B.n811 B.n4 10.6151
R2165 B.n815 B.n4 10.6151
R2166 B.n816 B.n815 10.6151
R2167 B.n817 B.n816 10.6151
R2168 B.n817 B.n0 10.6151
R2169 B.n768 B.n767 10.6151
R2170 B.n767 B.n20 10.6151
R2171 B.n763 B.n20 10.6151
R2172 B.n763 B.n762 10.6151
R2173 B.n762 B.n761 10.6151
R2174 B.n761 B.n22 10.6151
R2175 B.n757 B.n22 10.6151
R2176 B.n757 B.n756 10.6151
R2177 B.n756 B.n755 10.6151
R2178 B.n755 B.n24 10.6151
R2179 B.n751 B.n24 10.6151
R2180 B.n751 B.n750 10.6151
R2181 B.n750 B.n749 10.6151
R2182 B.n749 B.n26 10.6151
R2183 B.n745 B.n26 10.6151
R2184 B.n745 B.n744 10.6151
R2185 B.n744 B.n743 10.6151
R2186 B.n743 B.n28 10.6151
R2187 B.n739 B.n28 10.6151
R2188 B.n739 B.n738 10.6151
R2189 B.n738 B.n737 10.6151
R2190 B.n737 B.n30 10.6151
R2191 B.n733 B.n30 10.6151
R2192 B.n733 B.n732 10.6151
R2193 B.n732 B.n731 10.6151
R2194 B.n731 B.n32 10.6151
R2195 B.n727 B.n32 10.6151
R2196 B.n727 B.n726 10.6151
R2197 B.n726 B.n725 10.6151
R2198 B.n725 B.n34 10.6151
R2199 B.n721 B.n34 10.6151
R2200 B.n721 B.n720 10.6151
R2201 B.n720 B.n719 10.6151
R2202 B.n719 B.n36 10.6151
R2203 B.n715 B.n36 10.6151
R2204 B.n715 B.n714 10.6151
R2205 B.n714 B.n713 10.6151
R2206 B.n713 B.n38 10.6151
R2207 B.n709 B.n38 10.6151
R2208 B.n709 B.n708 10.6151
R2209 B.n708 B.n707 10.6151
R2210 B.n707 B.n40 10.6151
R2211 B.n703 B.n40 10.6151
R2212 B.n703 B.n702 10.6151
R2213 B.n702 B.n701 10.6151
R2214 B.n701 B.n42 10.6151
R2215 B.n697 B.n42 10.6151
R2216 B.n697 B.n696 10.6151
R2217 B.n696 B.n695 10.6151
R2218 B.n695 B.n44 10.6151
R2219 B.n691 B.n44 10.6151
R2220 B.n691 B.n690 10.6151
R2221 B.n690 B.n689 10.6151
R2222 B.n689 B.n46 10.6151
R2223 B.n685 B.n46 10.6151
R2224 B.n685 B.n684 10.6151
R2225 B.n684 B.n683 10.6151
R2226 B.n683 B.n48 10.6151
R2227 B.n679 B.n48 10.6151
R2228 B.n679 B.n678 10.6151
R2229 B.n678 B.n677 10.6151
R2230 B.n674 B.n673 10.6151
R2231 B.n673 B.n672 10.6151
R2232 B.n672 B.n54 10.6151
R2233 B.n668 B.n54 10.6151
R2234 B.n668 B.n667 10.6151
R2235 B.n667 B.n666 10.6151
R2236 B.n666 B.n56 10.6151
R2237 B.n662 B.n56 10.6151
R2238 B.n660 B.n659 10.6151
R2239 B.n659 B.n60 10.6151
R2240 B.n655 B.n60 10.6151
R2241 B.n655 B.n654 10.6151
R2242 B.n654 B.n653 10.6151
R2243 B.n653 B.n62 10.6151
R2244 B.n649 B.n62 10.6151
R2245 B.n649 B.n648 10.6151
R2246 B.n648 B.n647 10.6151
R2247 B.n647 B.n64 10.6151
R2248 B.n643 B.n64 10.6151
R2249 B.n643 B.n642 10.6151
R2250 B.n642 B.n641 10.6151
R2251 B.n641 B.n66 10.6151
R2252 B.n637 B.n66 10.6151
R2253 B.n637 B.n636 10.6151
R2254 B.n636 B.n635 10.6151
R2255 B.n635 B.n68 10.6151
R2256 B.n631 B.n68 10.6151
R2257 B.n631 B.n630 10.6151
R2258 B.n630 B.n629 10.6151
R2259 B.n629 B.n70 10.6151
R2260 B.n625 B.n70 10.6151
R2261 B.n625 B.n624 10.6151
R2262 B.n624 B.n623 10.6151
R2263 B.n623 B.n72 10.6151
R2264 B.n619 B.n72 10.6151
R2265 B.n619 B.n618 10.6151
R2266 B.n618 B.n617 10.6151
R2267 B.n617 B.n74 10.6151
R2268 B.n613 B.n74 10.6151
R2269 B.n613 B.n612 10.6151
R2270 B.n612 B.n611 10.6151
R2271 B.n611 B.n76 10.6151
R2272 B.n607 B.n76 10.6151
R2273 B.n607 B.n606 10.6151
R2274 B.n606 B.n605 10.6151
R2275 B.n605 B.n78 10.6151
R2276 B.n601 B.n78 10.6151
R2277 B.n601 B.n600 10.6151
R2278 B.n600 B.n599 10.6151
R2279 B.n599 B.n80 10.6151
R2280 B.n595 B.n80 10.6151
R2281 B.n595 B.n594 10.6151
R2282 B.n594 B.n593 10.6151
R2283 B.n593 B.n82 10.6151
R2284 B.n589 B.n82 10.6151
R2285 B.n589 B.n588 10.6151
R2286 B.n588 B.n587 10.6151
R2287 B.n587 B.n84 10.6151
R2288 B.n583 B.n84 10.6151
R2289 B.n583 B.n582 10.6151
R2290 B.n582 B.n581 10.6151
R2291 B.n581 B.n86 10.6151
R2292 B.n577 B.n86 10.6151
R2293 B.n577 B.n576 10.6151
R2294 B.n576 B.n575 10.6151
R2295 B.n575 B.n88 10.6151
R2296 B.n571 B.n88 10.6151
R2297 B.n571 B.n570 10.6151
R2298 B.n570 B.n569 10.6151
R2299 B.n565 B.n90 10.6151
R2300 B.n565 B.n564 10.6151
R2301 B.n564 B.n563 10.6151
R2302 B.n563 B.n92 10.6151
R2303 B.n559 B.n92 10.6151
R2304 B.n559 B.n558 10.6151
R2305 B.n558 B.n557 10.6151
R2306 B.n557 B.n94 10.6151
R2307 B.n553 B.n94 10.6151
R2308 B.n553 B.n552 10.6151
R2309 B.n552 B.n551 10.6151
R2310 B.n551 B.n96 10.6151
R2311 B.n547 B.n96 10.6151
R2312 B.n547 B.n546 10.6151
R2313 B.n546 B.n545 10.6151
R2314 B.n545 B.n98 10.6151
R2315 B.n541 B.n98 10.6151
R2316 B.n541 B.n540 10.6151
R2317 B.n540 B.n539 10.6151
R2318 B.n539 B.n100 10.6151
R2319 B.n535 B.n100 10.6151
R2320 B.n535 B.n534 10.6151
R2321 B.n534 B.n533 10.6151
R2322 B.n533 B.n102 10.6151
R2323 B.n529 B.n102 10.6151
R2324 B.n529 B.n528 10.6151
R2325 B.n528 B.n527 10.6151
R2326 B.n527 B.n104 10.6151
R2327 B.n523 B.n104 10.6151
R2328 B.n523 B.n522 10.6151
R2329 B.n522 B.n521 10.6151
R2330 B.n521 B.n106 10.6151
R2331 B.n517 B.n106 10.6151
R2332 B.n517 B.n516 10.6151
R2333 B.n516 B.n515 10.6151
R2334 B.n515 B.n108 10.6151
R2335 B.n511 B.n108 10.6151
R2336 B.n511 B.n510 10.6151
R2337 B.n510 B.n509 10.6151
R2338 B.n509 B.n110 10.6151
R2339 B.n505 B.n110 10.6151
R2340 B.n505 B.n504 10.6151
R2341 B.n504 B.n503 10.6151
R2342 B.n503 B.n112 10.6151
R2343 B.n499 B.n112 10.6151
R2344 B.n499 B.n498 10.6151
R2345 B.n498 B.n497 10.6151
R2346 B.n497 B.n114 10.6151
R2347 B.n493 B.n114 10.6151
R2348 B.n493 B.n492 10.6151
R2349 B.n492 B.n491 10.6151
R2350 B.n491 B.n116 10.6151
R2351 B.n487 B.n116 10.6151
R2352 B.n487 B.n486 10.6151
R2353 B.n486 B.n485 10.6151
R2354 B.n485 B.n118 10.6151
R2355 B.n481 B.n118 10.6151
R2356 B.n481 B.n480 10.6151
R2357 B.n480 B.n479 10.6151
R2358 B.n479 B.n120 10.6151
R2359 B.n475 B.n120 10.6151
R2360 B.n475 B.n474 10.6151
R2361 B.n474 B.n473 10.6151
R2362 B.n473 B.n122 10.6151
R2363 B.n469 B.n122 10.6151
R2364 B.n469 B.n468 10.6151
R2365 B.n468 B.n467 10.6151
R2366 B.n467 B.n124 10.6151
R2367 B.n463 B.n124 10.6151
R2368 B.n212 B.n1 10.6151
R2369 B.n215 B.n212 10.6151
R2370 B.n216 B.n215 10.6151
R2371 B.n217 B.n216 10.6151
R2372 B.n217 B.n210 10.6151
R2373 B.n221 B.n210 10.6151
R2374 B.n222 B.n221 10.6151
R2375 B.n223 B.n222 10.6151
R2376 B.n223 B.n208 10.6151
R2377 B.n227 B.n208 10.6151
R2378 B.n228 B.n227 10.6151
R2379 B.n229 B.n228 10.6151
R2380 B.n229 B.n206 10.6151
R2381 B.n233 B.n206 10.6151
R2382 B.n234 B.n233 10.6151
R2383 B.n235 B.n234 10.6151
R2384 B.n235 B.n204 10.6151
R2385 B.n239 B.n204 10.6151
R2386 B.n240 B.n239 10.6151
R2387 B.n241 B.n240 10.6151
R2388 B.n241 B.n202 10.6151
R2389 B.n245 B.n202 10.6151
R2390 B.n246 B.n245 10.6151
R2391 B.n247 B.n246 10.6151
R2392 B.n247 B.n200 10.6151
R2393 B.n251 B.n200 10.6151
R2394 B.n252 B.n251 10.6151
R2395 B.n253 B.n252 10.6151
R2396 B.n253 B.n198 10.6151
R2397 B.n257 B.n198 10.6151
R2398 B.n258 B.n257 10.6151
R2399 B.n259 B.n258 10.6151
R2400 B.n259 B.n196 10.6151
R2401 B.n264 B.n263 10.6151
R2402 B.n265 B.n264 10.6151
R2403 B.n265 B.n194 10.6151
R2404 B.n269 B.n194 10.6151
R2405 B.n270 B.n269 10.6151
R2406 B.n271 B.n270 10.6151
R2407 B.n271 B.n192 10.6151
R2408 B.n275 B.n192 10.6151
R2409 B.n276 B.n275 10.6151
R2410 B.n277 B.n276 10.6151
R2411 B.n277 B.n190 10.6151
R2412 B.n281 B.n190 10.6151
R2413 B.n282 B.n281 10.6151
R2414 B.n283 B.n282 10.6151
R2415 B.n283 B.n188 10.6151
R2416 B.n287 B.n188 10.6151
R2417 B.n288 B.n287 10.6151
R2418 B.n289 B.n288 10.6151
R2419 B.n289 B.n186 10.6151
R2420 B.n293 B.n186 10.6151
R2421 B.n294 B.n293 10.6151
R2422 B.n295 B.n294 10.6151
R2423 B.n295 B.n184 10.6151
R2424 B.n299 B.n184 10.6151
R2425 B.n300 B.n299 10.6151
R2426 B.n301 B.n300 10.6151
R2427 B.n301 B.n182 10.6151
R2428 B.n305 B.n182 10.6151
R2429 B.n306 B.n305 10.6151
R2430 B.n307 B.n306 10.6151
R2431 B.n307 B.n180 10.6151
R2432 B.n311 B.n180 10.6151
R2433 B.n312 B.n311 10.6151
R2434 B.n313 B.n312 10.6151
R2435 B.n313 B.n178 10.6151
R2436 B.n317 B.n178 10.6151
R2437 B.n318 B.n317 10.6151
R2438 B.n319 B.n318 10.6151
R2439 B.n319 B.n176 10.6151
R2440 B.n323 B.n176 10.6151
R2441 B.n324 B.n323 10.6151
R2442 B.n325 B.n324 10.6151
R2443 B.n325 B.n174 10.6151
R2444 B.n329 B.n174 10.6151
R2445 B.n330 B.n329 10.6151
R2446 B.n331 B.n330 10.6151
R2447 B.n331 B.n172 10.6151
R2448 B.n335 B.n172 10.6151
R2449 B.n336 B.n335 10.6151
R2450 B.n337 B.n336 10.6151
R2451 B.n337 B.n170 10.6151
R2452 B.n341 B.n170 10.6151
R2453 B.n342 B.n341 10.6151
R2454 B.n343 B.n342 10.6151
R2455 B.n343 B.n168 10.6151
R2456 B.n347 B.n168 10.6151
R2457 B.n348 B.n347 10.6151
R2458 B.n349 B.n348 10.6151
R2459 B.n349 B.n166 10.6151
R2460 B.n353 B.n166 10.6151
R2461 B.n354 B.n353 10.6151
R2462 B.n356 B.n162 10.6151
R2463 B.n360 B.n162 10.6151
R2464 B.n361 B.n360 10.6151
R2465 B.n362 B.n361 10.6151
R2466 B.n362 B.n160 10.6151
R2467 B.n366 B.n160 10.6151
R2468 B.n367 B.n366 10.6151
R2469 B.n368 B.n367 10.6151
R2470 B.n372 B.n371 10.6151
R2471 B.n373 B.n372 10.6151
R2472 B.n373 B.n154 10.6151
R2473 B.n377 B.n154 10.6151
R2474 B.n378 B.n377 10.6151
R2475 B.n379 B.n378 10.6151
R2476 B.n379 B.n152 10.6151
R2477 B.n383 B.n152 10.6151
R2478 B.n384 B.n383 10.6151
R2479 B.n385 B.n384 10.6151
R2480 B.n385 B.n150 10.6151
R2481 B.n389 B.n150 10.6151
R2482 B.n390 B.n389 10.6151
R2483 B.n391 B.n390 10.6151
R2484 B.n391 B.n148 10.6151
R2485 B.n395 B.n148 10.6151
R2486 B.n396 B.n395 10.6151
R2487 B.n397 B.n396 10.6151
R2488 B.n397 B.n146 10.6151
R2489 B.n401 B.n146 10.6151
R2490 B.n402 B.n401 10.6151
R2491 B.n403 B.n402 10.6151
R2492 B.n403 B.n144 10.6151
R2493 B.n407 B.n144 10.6151
R2494 B.n408 B.n407 10.6151
R2495 B.n409 B.n408 10.6151
R2496 B.n409 B.n142 10.6151
R2497 B.n413 B.n142 10.6151
R2498 B.n414 B.n413 10.6151
R2499 B.n415 B.n414 10.6151
R2500 B.n415 B.n140 10.6151
R2501 B.n419 B.n140 10.6151
R2502 B.n420 B.n419 10.6151
R2503 B.n421 B.n420 10.6151
R2504 B.n421 B.n138 10.6151
R2505 B.n425 B.n138 10.6151
R2506 B.n426 B.n425 10.6151
R2507 B.n427 B.n426 10.6151
R2508 B.n427 B.n136 10.6151
R2509 B.n431 B.n136 10.6151
R2510 B.n432 B.n431 10.6151
R2511 B.n433 B.n432 10.6151
R2512 B.n433 B.n134 10.6151
R2513 B.n437 B.n134 10.6151
R2514 B.n438 B.n437 10.6151
R2515 B.n439 B.n438 10.6151
R2516 B.n439 B.n132 10.6151
R2517 B.n443 B.n132 10.6151
R2518 B.n444 B.n443 10.6151
R2519 B.n445 B.n444 10.6151
R2520 B.n445 B.n130 10.6151
R2521 B.n449 B.n130 10.6151
R2522 B.n450 B.n449 10.6151
R2523 B.n451 B.n450 10.6151
R2524 B.n451 B.n128 10.6151
R2525 B.n455 B.n128 10.6151
R2526 B.n456 B.n455 10.6151
R2527 B.n457 B.n456 10.6151
R2528 B.n457 B.n126 10.6151
R2529 B.n461 B.n126 10.6151
R2530 B.n462 B.n461 10.6151
R2531 B.n821 B.n0 8.11757
R2532 B.n821 B.n1 8.11757
R2533 B.n674 B.n52 6.5566
R2534 B.n662 B.n661 6.5566
R2535 B.n356 B.n355 6.5566
R2536 B.n368 B.n158 6.5566
R2537 B.n677 B.n52 4.05904
R2538 B.n661 B.n660 4.05904
R2539 B.n355 B.n354 4.05904
R2540 B.n371 B.n158 4.05904
C0 VDD1 VN 0.149233f
C1 w_n2770_n4732# VDD2 1.70469f
C2 VDD2 B 1.51029f
C3 VDD2 VN 7.31073f
C4 VDD1 VTAIL 7.02481f
C5 VDD2 VTAIL 7.07948f
C6 w_n2770_n4732# VP 5.1957f
C7 B VP 1.79741f
C8 VDD1 VDD2 1.03629f
C9 VN VP 7.50455f
C10 w_n2770_n4732# B 11.244499f
C11 VTAIL VP 6.93426f
C12 w_n2770_n4732# VN 4.83943f
C13 VN B 1.20587f
C14 VDD1 VP 7.55967f
C15 VDD2 VP 0.398929f
C16 w_n2770_n4732# VTAIL 5.50547f
C17 VTAIL B 7.22531f
C18 VN VTAIL 6.92016f
C19 w_n2770_n4732# VDD1 1.64702f
C20 VDD1 B 1.45699f
C21 VDD2 VSUBS 1.127475f
C22 VDD1 VSUBS 6.63304f
C23 VTAIL VSUBS 1.545952f
C24 VN VSUBS 5.74516f
C25 VP VSUBS 2.585169f
C26 B VSUBS 4.913567f
C27 w_n2770_n4732# VSUBS 0.160184p
C28 B.n0 VSUBS 0.005225f
C29 B.n1 VSUBS 0.005225f
C30 B.n2 VSUBS 0.007727f
C31 B.n3 VSUBS 0.005922f
C32 B.n4 VSUBS 0.005922f
C33 B.n5 VSUBS 0.005922f
C34 B.n6 VSUBS 0.005922f
C35 B.n7 VSUBS 0.005922f
C36 B.n8 VSUBS 0.005922f
C37 B.n9 VSUBS 0.005922f
C38 B.n10 VSUBS 0.005922f
C39 B.n11 VSUBS 0.005922f
C40 B.n12 VSUBS 0.005922f
C41 B.n13 VSUBS 0.005922f
C42 B.n14 VSUBS 0.005922f
C43 B.n15 VSUBS 0.005922f
C44 B.n16 VSUBS 0.005922f
C45 B.n17 VSUBS 0.005922f
C46 B.n18 VSUBS 0.005922f
C47 B.n19 VSUBS 0.014331f
C48 B.n20 VSUBS 0.005922f
C49 B.n21 VSUBS 0.005922f
C50 B.n22 VSUBS 0.005922f
C51 B.n23 VSUBS 0.005922f
C52 B.n24 VSUBS 0.005922f
C53 B.n25 VSUBS 0.005922f
C54 B.n26 VSUBS 0.005922f
C55 B.n27 VSUBS 0.005922f
C56 B.n28 VSUBS 0.005922f
C57 B.n29 VSUBS 0.005922f
C58 B.n30 VSUBS 0.005922f
C59 B.n31 VSUBS 0.005922f
C60 B.n32 VSUBS 0.005922f
C61 B.n33 VSUBS 0.005922f
C62 B.n34 VSUBS 0.005922f
C63 B.n35 VSUBS 0.005922f
C64 B.n36 VSUBS 0.005922f
C65 B.n37 VSUBS 0.005922f
C66 B.n38 VSUBS 0.005922f
C67 B.n39 VSUBS 0.005922f
C68 B.n40 VSUBS 0.005922f
C69 B.n41 VSUBS 0.005922f
C70 B.n42 VSUBS 0.005922f
C71 B.n43 VSUBS 0.005922f
C72 B.n44 VSUBS 0.005922f
C73 B.n45 VSUBS 0.005922f
C74 B.n46 VSUBS 0.005922f
C75 B.n47 VSUBS 0.005922f
C76 B.n48 VSUBS 0.005922f
C77 B.n49 VSUBS 0.005922f
C78 B.t7 VSUBS 0.313756f
C79 B.t8 VSUBS 0.342835f
C80 B.t6 VSUBS 1.88355f
C81 B.n50 VSUBS 0.52572f
C82 B.n51 VSUBS 0.286621f
C83 B.n52 VSUBS 0.013719f
C84 B.n53 VSUBS 0.005922f
C85 B.n54 VSUBS 0.005922f
C86 B.n55 VSUBS 0.005922f
C87 B.n56 VSUBS 0.005922f
C88 B.n57 VSUBS 0.005922f
C89 B.t1 VSUBS 0.313759f
C90 B.t2 VSUBS 0.342838f
C91 B.t0 VSUBS 1.88355f
C92 B.n58 VSUBS 0.525717f
C93 B.n59 VSUBS 0.286617f
C94 B.n60 VSUBS 0.005922f
C95 B.n61 VSUBS 0.005922f
C96 B.n62 VSUBS 0.005922f
C97 B.n63 VSUBS 0.005922f
C98 B.n64 VSUBS 0.005922f
C99 B.n65 VSUBS 0.005922f
C100 B.n66 VSUBS 0.005922f
C101 B.n67 VSUBS 0.005922f
C102 B.n68 VSUBS 0.005922f
C103 B.n69 VSUBS 0.005922f
C104 B.n70 VSUBS 0.005922f
C105 B.n71 VSUBS 0.005922f
C106 B.n72 VSUBS 0.005922f
C107 B.n73 VSUBS 0.005922f
C108 B.n74 VSUBS 0.005922f
C109 B.n75 VSUBS 0.005922f
C110 B.n76 VSUBS 0.005922f
C111 B.n77 VSUBS 0.005922f
C112 B.n78 VSUBS 0.005922f
C113 B.n79 VSUBS 0.005922f
C114 B.n80 VSUBS 0.005922f
C115 B.n81 VSUBS 0.005922f
C116 B.n82 VSUBS 0.005922f
C117 B.n83 VSUBS 0.005922f
C118 B.n84 VSUBS 0.005922f
C119 B.n85 VSUBS 0.005922f
C120 B.n86 VSUBS 0.005922f
C121 B.n87 VSUBS 0.005922f
C122 B.n88 VSUBS 0.005922f
C123 B.n89 VSUBS 0.005922f
C124 B.n90 VSUBS 0.013535f
C125 B.n91 VSUBS 0.005922f
C126 B.n92 VSUBS 0.005922f
C127 B.n93 VSUBS 0.005922f
C128 B.n94 VSUBS 0.005922f
C129 B.n95 VSUBS 0.005922f
C130 B.n96 VSUBS 0.005922f
C131 B.n97 VSUBS 0.005922f
C132 B.n98 VSUBS 0.005922f
C133 B.n99 VSUBS 0.005922f
C134 B.n100 VSUBS 0.005922f
C135 B.n101 VSUBS 0.005922f
C136 B.n102 VSUBS 0.005922f
C137 B.n103 VSUBS 0.005922f
C138 B.n104 VSUBS 0.005922f
C139 B.n105 VSUBS 0.005922f
C140 B.n106 VSUBS 0.005922f
C141 B.n107 VSUBS 0.005922f
C142 B.n108 VSUBS 0.005922f
C143 B.n109 VSUBS 0.005922f
C144 B.n110 VSUBS 0.005922f
C145 B.n111 VSUBS 0.005922f
C146 B.n112 VSUBS 0.005922f
C147 B.n113 VSUBS 0.005922f
C148 B.n114 VSUBS 0.005922f
C149 B.n115 VSUBS 0.005922f
C150 B.n116 VSUBS 0.005922f
C151 B.n117 VSUBS 0.005922f
C152 B.n118 VSUBS 0.005922f
C153 B.n119 VSUBS 0.005922f
C154 B.n120 VSUBS 0.005922f
C155 B.n121 VSUBS 0.005922f
C156 B.n122 VSUBS 0.005922f
C157 B.n123 VSUBS 0.005922f
C158 B.n124 VSUBS 0.005922f
C159 B.n125 VSUBS 0.014331f
C160 B.n126 VSUBS 0.005922f
C161 B.n127 VSUBS 0.005922f
C162 B.n128 VSUBS 0.005922f
C163 B.n129 VSUBS 0.005922f
C164 B.n130 VSUBS 0.005922f
C165 B.n131 VSUBS 0.005922f
C166 B.n132 VSUBS 0.005922f
C167 B.n133 VSUBS 0.005922f
C168 B.n134 VSUBS 0.005922f
C169 B.n135 VSUBS 0.005922f
C170 B.n136 VSUBS 0.005922f
C171 B.n137 VSUBS 0.005922f
C172 B.n138 VSUBS 0.005922f
C173 B.n139 VSUBS 0.005922f
C174 B.n140 VSUBS 0.005922f
C175 B.n141 VSUBS 0.005922f
C176 B.n142 VSUBS 0.005922f
C177 B.n143 VSUBS 0.005922f
C178 B.n144 VSUBS 0.005922f
C179 B.n145 VSUBS 0.005922f
C180 B.n146 VSUBS 0.005922f
C181 B.n147 VSUBS 0.005922f
C182 B.n148 VSUBS 0.005922f
C183 B.n149 VSUBS 0.005922f
C184 B.n150 VSUBS 0.005922f
C185 B.n151 VSUBS 0.005922f
C186 B.n152 VSUBS 0.005922f
C187 B.n153 VSUBS 0.005922f
C188 B.n154 VSUBS 0.005922f
C189 B.n155 VSUBS 0.005922f
C190 B.t5 VSUBS 0.313759f
C191 B.t4 VSUBS 0.342838f
C192 B.t3 VSUBS 1.88355f
C193 B.n156 VSUBS 0.525717f
C194 B.n157 VSUBS 0.286617f
C195 B.n158 VSUBS 0.013719f
C196 B.n159 VSUBS 0.005922f
C197 B.n160 VSUBS 0.005922f
C198 B.n161 VSUBS 0.005922f
C199 B.n162 VSUBS 0.005922f
C200 B.n163 VSUBS 0.005922f
C201 B.t11 VSUBS 0.313756f
C202 B.t10 VSUBS 0.342835f
C203 B.t9 VSUBS 1.88355f
C204 B.n164 VSUBS 0.52572f
C205 B.n165 VSUBS 0.286621f
C206 B.n166 VSUBS 0.005922f
C207 B.n167 VSUBS 0.005922f
C208 B.n168 VSUBS 0.005922f
C209 B.n169 VSUBS 0.005922f
C210 B.n170 VSUBS 0.005922f
C211 B.n171 VSUBS 0.005922f
C212 B.n172 VSUBS 0.005922f
C213 B.n173 VSUBS 0.005922f
C214 B.n174 VSUBS 0.005922f
C215 B.n175 VSUBS 0.005922f
C216 B.n176 VSUBS 0.005922f
C217 B.n177 VSUBS 0.005922f
C218 B.n178 VSUBS 0.005922f
C219 B.n179 VSUBS 0.005922f
C220 B.n180 VSUBS 0.005922f
C221 B.n181 VSUBS 0.005922f
C222 B.n182 VSUBS 0.005922f
C223 B.n183 VSUBS 0.005922f
C224 B.n184 VSUBS 0.005922f
C225 B.n185 VSUBS 0.005922f
C226 B.n186 VSUBS 0.005922f
C227 B.n187 VSUBS 0.005922f
C228 B.n188 VSUBS 0.005922f
C229 B.n189 VSUBS 0.005922f
C230 B.n190 VSUBS 0.005922f
C231 B.n191 VSUBS 0.005922f
C232 B.n192 VSUBS 0.005922f
C233 B.n193 VSUBS 0.005922f
C234 B.n194 VSUBS 0.005922f
C235 B.n195 VSUBS 0.005922f
C236 B.n196 VSUBS 0.013535f
C237 B.n197 VSUBS 0.005922f
C238 B.n198 VSUBS 0.005922f
C239 B.n199 VSUBS 0.005922f
C240 B.n200 VSUBS 0.005922f
C241 B.n201 VSUBS 0.005922f
C242 B.n202 VSUBS 0.005922f
C243 B.n203 VSUBS 0.005922f
C244 B.n204 VSUBS 0.005922f
C245 B.n205 VSUBS 0.005922f
C246 B.n206 VSUBS 0.005922f
C247 B.n207 VSUBS 0.005922f
C248 B.n208 VSUBS 0.005922f
C249 B.n209 VSUBS 0.005922f
C250 B.n210 VSUBS 0.005922f
C251 B.n211 VSUBS 0.005922f
C252 B.n212 VSUBS 0.005922f
C253 B.n213 VSUBS 0.005922f
C254 B.n214 VSUBS 0.005922f
C255 B.n215 VSUBS 0.005922f
C256 B.n216 VSUBS 0.005922f
C257 B.n217 VSUBS 0.005922f
C258 B.n218 VSUBS 0.005922f
C259 B.n219 VSUBS 0.005922f
C260 B.n220 VSUBS 0.005922f
C261 B.n221 VSUBS 0.005922f
C262 B.n222 VSUBS 0.005922f
C263 B.n223 VSUBS 0.005922f
C264 B.n224 VSUBS 0.005922f
C265 B.n225 VSUBS 0.005922f
C266 B.n226 VSUBS 0.005922f
C267 B.n227 VSUBS 0.005922f
C268 B.n228 VSUBS 0.005922f
C269 B.n229 VSUBS 0.005922f
C270 B.n230 VSUBS 0.005922f
C271 B.n231 VSUBS 0.005922f
C272 B.n232 VSUBS 0.005922f
C273 B.n233 VSUBS 0.005922f
C274 B.n234 VSUBS 0.005922f
C275 B.n235 VSUBS 0.005922f
C276 B.n236 VSUBS 0.005922f
C277 B.n237 VSUBS 0.005922f
C278 B.n238 VSUBS 0.005922f
C279 B.n239 VSUBS 0.005922f
C280 B.n240 VSUBS 0.005922f
C281 B.n241 VSUBS 0.005922f
C282 B.n242 VSUBS 0.005922f
C283 B.n243 VSUBS 0.005922f
C284 B.n244 VSUBS 0.005922f
C285 B.n245 VSUBS 0.005922f
C286 B.n246 VSUBS 0.005922f
C287 B.n247 VSUBS 0.005922f
C288 B.n248 VSUBS 0.005922f
C289 B.n249 VSUBS 0.005922f
C290 B.n250 VSUBS 0.005922f
C291 B.n251 VSUBS 0.005922f
C292 B.n252 VSUBS 0.005922f
C293 B.n253 VSUBS 0.005922f
C294 B.n254 VSUBS 0.005922f
C295 B.n255 VSUBS 0.005922f
C296 B.n256 VSUBS 0.005922f
C297 B.n257 VSUBS 0.005922f
C298 B.n258 VSUBS 0.005922f
C299 B.n259 VSUBS 0.005922f
C300 B.n260 VSUBS 0.005922f
C301 B.n261 VSUBS 0.013535f
C302 B.n262 VSUBS 0.014331f
C303 B.n263 VSUBS 0.014331f
C304 B.n264 VSUBS 0.005922f
C305 B.n265 VSUBS 0.005922f
C306 B.n266 VSUBS 0.005922f
C307 B.n267 VSUBS 0.005922f
C308 B.n268 VSUBS 0.005922f
C309 B.n269 VSUBS 0.005922f
C310 B.n270 VSUBS 0.005922f
C311 B.n271 VSUBS 0.005922f
C312 B.n272 VSUBS 0.005922f
C313 B.n273 VSUBS 0.005922f
C314 B.n274 VSUBS 0.005922f
C315 B.n275 VSUBS 0.005922f
C316 B.n276 VSUBS 0.005922f
C317 B.n277 VSUBS 0.005922f
C318 B.n278 VSUBS 0.005922f
C319 B.n279 VSUBS 0.005922f
C320 B.n280 VSUBS 0.005922f
C321 B.n281 VSUBS 0.005922f
C322 B.n282 VSUBS 0.005922f
C323 B.n283 VSUBS 0.005922f
C324 B.n284 VSUBS 0.005922f
C325 B.n285 VSUBS 0.005922f
C326 B.n286 VSUBS 0.005922f
C327 B.n287 VSUBS 0.005922f
C328 B.n288 VSUBS 0.005922f
C329 B.n289 VSUBS 0.005922f
C330 B.n290 VSUBS 0.005922f
C331 B.n291 VSUBS 0.005922f
C332 B.n292 VSUBS 0.005922f
C333 B.n293 VSUBS 0.005922f
C334 B.n294 VSUBS 0.005922f
C335 B.n295 VSUBS 0.005922f
C336 B.n296 VSUBS 0.005922f
C337 B.n297 VSUBS 0.005922f
C338 B.n298 VSUBS 0.005922f
C339 B.n299 VSUBS 0.005922f
C340 B.n300 VSUBS 0.005922f
C341 B.n301 VSUBS 0.005922f
C342 B.n302 VSUBS 0.005922f
C343 B.n303 VSUBS 0.005922f
C344 B.n304 VSUBS 0.005922f
C345 B.n305 VSUBS 0.005922f
C346 B.n306 VSUBS 0.005922f
C347 B.n307 VSUBS 0.005922f
C348 B.n308 VSUBS 0.005922f
C349 B.n309 VSUBS 0.005922f
C350 B.n310 VSUBS 0.005922f
C351 B.n311 VSUBS 0.005922f
C352 B.n312 VSUBS 0.005922f
C353 B.n313 VSUBS 0.005922f
C354 B.n314 VSUBS 0.005922f
C355 B.n315 VSUBS 0.005922f
C356 B.n316 VSUBS 0.005922f
C357 B.n317 VSUBS 0.005922f
C358 B.n318 VSUBS 0.005922f
C359 B.n319 VSUBS 0.005922f
C360 B.n320 VSUBS 0.005922f
C361 B.n321 VSUBS 0.005922f
C362 B.n322 VSUBS 0.005922f
C363 B.n323 VSUBS 0.005922f
C364 B.n324 VSUBS 0.005922f
C365 B.n325 VSUBS 0.005922f
C366 B.n326 VSUBS 0.005922f
C367 B.n327 VSUBS 0.005922f
C368 B.n328 VSUBS 0.005922f
C369 B.n329 VSUBS 0.005922f
C370 B.n330 VSUBS 0.005922f
C371 B.n331 VSUBS 0.005922f
C372 B.n332 VSUBS 0.005922f
C373 B.n333 VSUBS 0.005922f
C374 B.n334 VSUBS 0.005922f
C375 B.n335 VSUBS 0.005922f
C376 B.n336 VSUBS 0.005922f
C377 B.n337 VSUBS 0.005922f
C378 B.n338 VSUBS 0.005922f
C379 B.n339 VSUBS 0.005922f
C380 B.n340 VSUBS 0.005922f
C381 B.n341 VSUBS 0.005922f
C382 B.n342 VSUBS 0.005922f
C383 B.n343 VSUBS 0.005922f
C384 B.n344 VSUBS 0.005922f
C385 B.n345 VSUBS 0.005922f
C386 B.n346 VSUBS 0.005922f
C387 B.n347 VSUBS 0.005922f
C388 B.n348 VSUBS 0.005922f
C389 B.n349 VSUBS 0.005922f
C390 B.n350 VSUBS 0.005922f
C391 B.n351 VSUBS 0.005922f
C392 B.n352 VSUBS 0.005922f
C393 B.n353 VSUBS 0.005922f
C394 B.n354 VSUBS 0.004093f
C395 B.n355 VSUBS 0.013719f
C396 B.n356 VSUBS 0.004789f
C397 B.n357 VSUBS 0.005922f
C398 B.n358 VSUBS 0.005922f
C399 B.n359 VSUBS 0.005922f
C400 B.n360 VSUBS 0.005922f
C401 B.n361 VSUBS 0.005922f
C402 B.n362 VSUBS 0.005922f
C403 B.n363 VSUBS 0.005922f
C404 B.n364 VSUBS 0.005922f
C405 B.n365 VSUBS 0.005922f
C406 B.n366 VSUBS 0.005922f
C407 B.n367 VSUBS 0.005922f
C408 B.n368 VSUBS 0.004789f
C409 B.n369 VSUBS 0.005922f
C410 B.n370 VSUBS 0.005922f
C411 B.n371 VSUBS 0.004093f
C412 B.n372 VSUBS 0.005922f
C413 B.n373 VSUBS 0.005922f
C414 B.n374 VSUBS 0.005922f
C415 B.n375 VSUBS 0.005922f
C416 B.n376 VSUBS 0.005922f
C417 B.n377 VSUBS 0.005922f
C418 B.n378 VSUBS 0.005922f
C419 B.n379 VSUBS 0.005922f
C420 B.n380 VSUBS 0.005922f
C421 B.n381 VSUBS 0.005922f
C422 B.n382 VSUBS 0.005922f
C423 B.n383 VSUBS 0.005922f
C424 B.n384 VSUBS 0.005922f
C425 B.n385 VSUBS 0.005922f
C426 B.n386 VSUBS 0.005922f
C427 B.n387 VSUBS 0.005922f
C428 B.n388 VSUBS 0.005922f
C429 B.n389 VSUBS 0.005922f
C430 B.n390 VSUBS 0.005922f
C431 B.n391 VSUBS 0.005922f
C432 B.n392 VSUBS 0.005922f
C433 B.n393 VSUBS 0.005922f
C434 B.n394 VSUBS 0.005922f
C435 B.n395 VSUBS 0.005922f
C436 B.n396 VSUBS 0.005922f
C437 B.n397 VSUBS 0.005922f
C438 B.n398 VSUBS 0.005922f
C439 B.n399 VSUBS 0.005922f
C440 B.n400 VSUBS 0.005922f
C441 B.n401 VSUBS 0.005922f
C442 B.n402 VSUBS 0.005922f
C443 B.n403 VSUBS 0.005922f
C444 B.n404 VSUBS 0.005922f
C445 B.n405 VSUBS 0.005922f
C446 B.n406 VSUBS 0.005922f
C447 B.n407 VSUBS 0.005922f
C448 B.n408 VSUBS 0.005922f
C449 B.n409 VSUBS 0.005922f
C450 B.n410 VSUBS 0.005922f
C451 B.n411 VSUBS 0.005922f
C452 B.n412 VSUBS 0.005922f
C453 B.n413 VSUBS 0.005922f
C454 B.n414 VSUBS 0.005922f
C455 B.n415 VSUBS 0.005922f
C456 B.n416 VSUBS 0.005922f
C457 B.n417 VSUBS 0.005922f
C458 B.n418 VSUBS 0.005922f
C459 B.n419 VSUBS 0.005922f
C460 B.n420 VSUBS 0.005922f
C461 B.n421 VSUBS 0.005922f
C462 B.n422 VSUBS 0.005922f
C463 B.n423 VSUBS 0.005922f
C464 B.n424 VSUBS 0.005922f
C465 B.n425 VSUBS 0.005922f
C466 B.n426 VSUBS 0.005922f
C467 B.n427 VSUBS 0.005922f
C468 B.n428 VSUBS 0.005922f
C469 B.n429 VSUBS 0.005922f
C470 B.n430 VSUBS 0.005922f
C471 B.n431 VSUBS 0.005922f
C472 B.n432 VSUBS 0.005922f
C473 B.n433 VSUBS 0.005922f
C474 B.n434 VSUBS 0.005922f
C475 B.n435 VSUBS 0.005922f
C476 B.n436 VSUBS 0.005922f
C477 B.n437 VSUBS 0.005922f
C478 B.n438 VSUBS 0.005922f
C479 B.n439 VSUBS 0.005922f
C480 B.n440 VSUBS 0.005922f
C481 B.n441 VSUBS 0.005922f
C482 B.n442 VSUBS 0.005922f
C483 B.n443 VSUBS 0.005922f
C484 B.n444 VSUBS 0.005922f
C485 B.n445 VSUBS 0.005922f
C486 B.n446 VSUBS 0.005922f
C487 B.n447 VSUBS 0.005922f
C488 B.n448 VSUBS 0.005922f
C489 B.n449 VSUBS 0.005922f
C490 B.n450 VSUBS 0.005922f
C491 B.n451 VSUBS 0.005922f
C492 B.n452 VSUBS 0.005922f
C493 B.n453 VSUBS 0.005922f
C494 B.n454 VSUBS 0.005922f
C495 B.n455 VSUBS 0.005922f
C496 B.n456 VSUBS 0.005922f
C497 B.n457 VSUBS 0.005922f
C498 B.n458 VSUBS 0.005922f
C499 B.n459 VSUBS 0.005922f
C500 B.n460 VSUBS 0.005922f
C501 B.n461 VSUBS 0.005922f
C502 B.n462 VSUBS 0.013637f
C503 B.n463 VSUBS 0.014229f
C504 B.n464 VSUBS 0.013535f
C505 B.n465 VSUBS 0.005922f
C506 B.n466 VSUBS 0.005922f
C507 B.n467 VSUBS 0.005922f
C508 B.n468 VSUBS 0.005922f
C509 B.n469 VSUBS 0.005922f
C510 B.n470 VSUBS 0.005922f
C511 B.n471 VSUBS 0.005922f
C512 B.n472 VSUBS 0.005922f
C513 B.n473 VSUBS 0.005922f
C514 B.n474 VSUBS 0.005922f
C515 B.n475 VSUBS 0.005922f
C516 B.n476 VSUBS 0.005922f
C517 B.n477 VSUBS 0.005922f
C518 B.n478 VSUBS 0.005922f
C519 B.n479 VSUBS 0.005922f
C520 B.n480 VSUBS 0.005922f
C521 B.n481 VSUBS 0.005922f
C522 B.n482 VSUBS 0.005922f
C523 B.n483 VSUBS 0.005922f
C524 B.n484 VSUBS 0.005922f
C525 B.n485 VSUBS 0.005922f
C526 B.n486 VSUBS 0.005922f
C527 B.n487 VSUBS 0.005922f
C528 B.n488 VSUBS 0.005922f
C529 B.n489 VSUBS 0.005922f
C530 B.n490 VSUBS 0.005922f
C531 B.n491 VSUBS 0.005922f
C532 B.n492 VSUBS 0.005922f
C533 B.n493 VSUBS 0.005922f
C534 B.n494 VSUBS 0.005922f
C535 B.n495 VSUBS 0.005922f
C536 B.n496 VSUBS 0.005922f
C537 B.n497 VSUBS 0.005922f
C538 B.n498 VSUBS 0.005922f
C539 B.n499 VSUBS 0.005922f
C540 B.n500 VSUBS 0.005922f
C541 B.n501 VSUBS 0.005922f
C542 B.n502 VSUBS 0.005922f
C543 B.n503 VSUBS 0.005922f
C544 B.n504 VSUBS 0.005922f
C545 B.n505 VSUBS 0.005922f
C546 B.n506 VSUBS 0.005922f
C547 B.n507 VSUBS 0.005922f
C548 B.n508 VSUBS 0.005922f
C549 B.n509 VSUBS 0.005922f
C550 B.n510 VSUBS 0.005922f
C551 B.n511 VSUBS 0.005922f
C552 B.n512 VSUBS 0.005922f
C553 B.n513 VSUBS 0.005922f
C554 B.n514 VSUBS 0.005922f
C555 B.n515 VSUBS 0.005922f
C556 B.n516 VSUBS 0.005922f
C557 B.n517 VSUBS 0.005922f
C558 B.n518 VSUBS 0.005922f
C559 B.n519 VSUBS 0.005922f
C560 B.n520 VSUBS 0.005922f
C561 B.n521 VSUBS 0.005922f
C562 B.n522 VSUBS 0.005922f
C563 B.n523 VSUBS 0.005922f
C564 B.n524 VSUBS 0.005922f
C565 B.n525 VSUBS 0.005922f
C566 B.n526 VSUBS 0.005922f
C567 B.n527 VSUBS 0.005922f
C568 B.n528 VSUBS 0.005922f
C569 B.n529 VSUBS 0.005922f
C570 B.n530 VSUBS 0.005922f
C571 B.n531 VSUBS 0.005922f
C572 B.n532 VSUBS 0.005922f
C573 B.n533 VSUBS 0.005922f
C574 B.n534 VSUBS 0.005922f
C575 B.n535 VSUBS 0.005922f
C576 B.n536 VSUBS 0.005922f
C577 B.n537 VSUBS 0.005922f
C578 B.n538 VSUBS 0.005922f
C579 B.n539 VSUBS 0.005922f
C580 B.n540 VSUBS 0.005922f
C581 B.n541 VSUBS 0.005922f
C582 B.n542 VSUBS 0.005922f
C583 B.n543 VSUBS 0.005922f
C584 B.n544 VSUBS 0.005922f
C585 B.n545 VSUBS 0.005922f
C586 B.n546 VSUBS 0.005922f
C587 B.n547 VSUBS 0.005922f
C588 B.n548 VSUBS 0.005922f
C589 B.n549 VSUBS 0.005922f
C590 B.n550 VSUBS 0.005922f
C591 B.n551 VSUBS 0.005922f
C592 B.n552 VSUBS 0.005922f
C593 B.n553 VSUBS 0.005922f
C594 B.n554 VSUBS 0.005922f
C595 B.n555 VSUBS 0.005922f
C596 B.n556 VSUBS 0.005922f
C597 B.n557 VSUBS 0.005922f
C598 B.n558 VSUBS 0.005922f
C599 B.n559 VSUBS 0.005922f
C600 B.n560 VSUBS 0.005922f
C601 B.n561 VSUBS 0.005922f
C602 B.n562 VSUBS 0.005922f
C603 B.n563 VSUBS 0.005922f
C604 B.n564 VSUBS 0.005922f
C605 B.n565 VSUBS 0.005922f
C606 B.n566 VSUBS 0.005922f
C607 B.n567 VSUBS 0.013535f
C608 B.n568 VSUBS 0.014331f
C609 B.n569 VSUBS 0.014331f
C610 B.n570 VSUBS 0.005922f
C611 B.n571 VSUBS 0.005922f
C612 B.n572 VSUBS 0.005922f
C613 B.n573 VSUBS 0.005922f
C614 B.n574 VSUBS 0.005922f
C615 B.n575 VSUBS 0.005922f
C616 B.n576 VSUBS 0.005922f
C617 B.n577 VSUBS 0.005922f
C618 B.n578 VSUBS 0.005922f
C619 B.n579 VSUBS 0.005922f
C620 B.n580 VSUBS 0.005922f
C621 B.n581 VSUBS 0.005922f
C622 B.n582 VSUBS 0.005922f
C623 B.n583 VSUBS 0.005922f
C624 B.n584 VSUBS 0.005922f
C625 B.n585 VSUBS 0.005922f
C626 B.n586 VSUBS 0.005922f
C627 B.n587 VSUBS 0.005922f
C628 B.n588 VSUBS 0.005922f
C629 B.n589 VSUBS 0.005922f
C630 B.n590 VSUBS 0.005922f
C631 B.n591 VSUBS 0.005922f
C632 B.n592 VSUBS 0.005922f
C633 B.n593 VSUBS 0.005922f
C634 B.n594 VSUBS 0.005922f
C635 B.n595 VSUBS 0.005922f
C636 B.n596 VSUBS 0.005922f
C637 B.n597 VSUBS 0.005922f
C638 B.n598 VSUBS 0.005922f
C639 B.n599 VSUBS 0.005922f
C640 B.n600 VSUBS 0.005922f
C641 B.n601 VSUBS 0.005922f
C642 B.n602 VSUBS 0.005922f
C643 B.n603 VSUBS 0.005922f
C644 B.n604 VSUBS 0.005922f
C645 B.n605 VSUBS 0.005922f
C646 B.n606 VSUBS 0.005922f
C647 B.n607 VSUBS 0.005922f
C648 B.n608 VSUBS 0.005922f
C649 B.n609 VSUBS 0.005922f
C650 B.n610 VSUBS 0.005922f
C651 B.n611 VSUBS 0.005922f
C652 B.n612 VSUBS 0.005922f
C653 B.n613 VSUBS 0.005922f
C654 B.n614 VSUBS 0.005922f
C655 B.n615 VSUBS 0.005922f
C656 B.n616 VSUBS 0.005922f
C657 B.n617 VSUBS 0.005922f
C658 B.n618 VSUBS 0.005922f
C659 B.n619 VSUBS 0.005922f
C660 B.n620 VSUBS 0.005922f
C661 B.n621 VSUBS 0.005922f
C662 B.n622 VSUBS 0.005922f
C663 B.n623 VSUBS 0.005922f
C664 B.n624 VSUBS 0.005922f
C665 B.n625 VSUBS 0.005922f
C666 B.n626 VSUBS 0.005922f
C667 B.n627 VSUBS 0.005922f
C668 B.n628 VSUBS 0.005922f
C669 B.n629 VSUBS 0.005922f
C670 B.n630 VSUBS 0.005922f
C671 B.n631 VSUBS 0.005922f
C672 B.n632 VSUBS 0.005922f
C673 B.n633 VSUBS 0.005922f
C674 B.n634 VSUBS 0.005922f
C675 B.n635 VSUBS 0.005922f
C676 B.n636 VSUBS 0.005922f
C677 B.n637 VSUBS 0.005922f
C678 B.n638 VSUBS 0.005922f
C679 B.n639 VSUBS 0.005922f
C680 B.n640 VSUBS 0.005922f
C681 B.n641 VSUBS 0.005922f
C682 B.n642 VSUBS 0.005922f
C683 B.n643 VSUBS 0.005922f
C684 B.n644 VSUBS 0.005922f
C685 B.n645 VSUBS 0.005922f
C686 B.n646 VSUBS 0.005922f
C687 B.n647 VSUBS 0.005922f
C688 B.n648 VSUBS 0.005922f
C689 B.n649 VSUBS 0.005922f
C690 B.n650 VSUBS 0.005922f
C691 B.n651 VSUBS 0.005922f
C692 B.n652 VSUBS 0.005922f
C693 B.n653 VSUBS 0.005922f
C694 B.n654 VSUBS 0.005922f
C695 B.n655 VSUBS 0.005922f
C696 B.n656 VSUBS 0.005922f
C697 B.n657 VSUBS 0.005922f
C698 B.n658 VSUBS 0.005922f
C699 B.n659 VSUBS 0.005922f
C700 B.n660 VSUBS 0.004093f
C701 B.n661 VSUBS 0.013719f
C702 B.n662 VSUBS 0.004789f
C703 B.n663 VSUBS 0.005922f
C704 B.n664 VSUBS 0.005922f
C705 B.n665 VSUBS 0.005922f
C706 B.n666 VSUBS 0.005922f
C707 B.n667 VSUBS 0.005922f
C708 B.n668 VSUBS 0.005922f
C709 B.n669 VSUBS 0.005922f
C710 B.n670 VSUBS 0.005922f
C711 B.n671 VSUBS 0.005922f
C712 B.n672 VSUBS 0.005922f
C713 B.n673 VSUBS 0.005922f
C714 B.n674 VSUBS 0.004789f
C715 B.n675 VSUBS 0.005922f
C716 B.n676 VSUBS 0.005922f
C717 B.n677 VSUBS 0.004093f
C718 B.n678 VSUBS 0.005922f
C719 B.n679 VSUBS 0.005922f
C720 B.n680 VSUBS 0.005922f
C721 B.n681 VSUBS 0.005922f
C722 B.n682 VSUBS 0.005922f
C723 B.n683 VSUBS 0.005922f
C724 B.n684 VSUBS 0.005922f
C725 B.n685 VSUBS 0.005922f
C726 B.n686 VSUBS 0.005922f
C727 B.n687 VSUBS 0.005922f
C728 B.n688 VSUBS 0.005922f
C729 B.n689 VSUBS 0.005922f
C730 B.n690 VSUBS 0.005922f
C731 B.n691 VSUBS 0.005922f
C732 B.n692 VSUBS 0.005922f
C733 B.n693 VSUBS 0.005922f
C734 B.n694 VSUBS 0.005922f
C735 B.n695 VSUBS 0.005922f
C736 B.n696 VSUBS 0.005922f
C737 B.n697 VSUBS 0.005922f
C738 B.n698 VSUBS 0.005922f
C739 B.n699 VSUBS 0.005922f
C740 B.n700 VSUBS 0.005922f
C741 B.n701 VSUBS 0.005922f
C742 B.n702 VSUBS 0.005922f
C743 B.n703 VSUBS 0.005922f
C744 B.n704 VSUBS 0.005922f
C745 B.n705 VSUBS 0.005922f
C746 B.n706 VSUBS 0.005922f
C747 B.n707 VSUBS 0.005922f
C748 B.n708 VSUBS 0.005922f
C749 B.n709 VSUBS 0.005922f
C750 B.n710 VSUBS 0.005922f
C751 B.n711 VSUBS 0.005922f
C752 B.n712 VSUBS 0.005922f
C753 B.n713 VSUBS 0.005922f
C754 B.n714 VSUBS 0.005922f
C755 B.n715 VSUBS 0.005922f
C756 B.n716 VSUBS 0.005922f
C757 B.n717 VSUBS 0.005922f
C758 B.n718 VSUBS 0.005922f
C759 B.n719 VSUBS 0.005922f
C760 B.n720 VSUBS 0.005922f
C761 B.n721 VSUBS 0.005922f
C762 B.n722 VSUBS 0.005922f
C763 B.n723 VSUBS 0.005922f
C764 B.n724 VSUBS 0.005922f
C765 B.n725 VSUBS 0.005922f
C766 B.n726 VSUBS 0.005922f
C767 B.n727 VSUBS 0.005922f
C768 B.n728 VSUBS 0.005922f
C769 B.n729 VSUBS 0.005922f
C770 B.n730 VSUBS 0.005922f
C771 B.n731 VSUBS 0.005922f
C772 B.n732 VSUBS 0.005922f
C773 B.n733 VSUBS 0.005922f
C774 B.n734 VSUBS 0.005922f
C775 B.n735 VSUBS 0.005922f
C776 B.n736 VSUBS 0.005922f
C777 B.n737 VSUBS 0.005922f
C778 B.n738 VSUBS 0.005922f
C779 B.n739 VSUBS 0.005922f
C780 B.n740 VSUBS 0.005922f
C781 B.n741 VSUBS 0.005922f
C782 B.n742 VSUBS 0.005922f
C783 B.n743 VSUBS 0.005922f
C784 B.n744 VSUBS 0.005922f
C785 B.n745 VSUBS 0.005922f
C786 B.n746 VSUBS 0.005922f
C787 B.n747 VSUBS 0.005922f
C788 B.n748 VSUBS 0.005922f
C789 B.n749 VSUBS 0.005922f
C790 B.n750 VSUBS 0.005922f
C791 B.n751 VSUBS 0.005922f
C792 B.n752 VSUBS 0.005922f
C793 B.n753 VSUBS 0.005922f
C794 B.n754 VSUBS 0.005922f
C795 B.n755 VSUBS 0.005922f
C796 B.n756 VSUBS 0.005922f
C797 B.n757 VSUBS 0.005922f
C798 B.n758 VSUBS 0.005922f
C799 B.n759 VSUBS 0.005922f
C800 B.n760 VSUBS 0.005922f
C801 B.n761 VSUBS 0.005922f
C802 B.n762 VSUBS 0.005922f
C803 B.n763 VSUBS 0.005922f
C804 B.n764 VSUBS 0.005922f
C805 B.n765 VSUBS 0.005922f
C806 B.n766 VSUBS 0.005922f
C807 B.n767 VSUBS 0.005922f
C808 B.n768 VSUBS 0.014331f
C809 B.n769 VSUBS 0.013535f
C810 B.n770 VSUBS 0.013535f
C811 B.n771 VSUBS 0.005922f
C812 B.n772 VSUBS 0.005922f
C813 B.n773 VSUBS 0.005922f
C814 B.n774 VSUBS 0.005922f
C815 B.n775 VSUBS 0.005922f
C816 B.n776 VSUBS 0.005922f
C817 B.n777 VSUBS 0.005922f
C818 B.n778 VSUBS 0.005922f
C819 B.n779 VSUBS 0.005922f
C820 B.n780 VSUBS 0.005922f
C821 B.n781 VSUBS 0.005922f
C822 B.n782 VSUBS 0.005922f
C823 B.n783 VSUBS 0.005922f
C824 B.n784 VSUBS 0.005922f
C825 B.n785 VSUBS 0.005922f
C826 B.n786 VSUBS 0.005922f
C827 B.n787 VSUBS 0.005922f
C828 B.n788 VSUBS 0.005922f
C829 B.n789 VSUBS 0.005922f
C830 B.n790 VSUBS 0.005922f
C831 B.n791 VSUBS 0.005922f
C832 B.n792 VSUBS 0.005922f
C833 B.n793 VSUBS 0.005922f
C834 B.n794 VSUBS 0.005922f
C835 B.n795 VSUBS 0.005922f
C836 B.n796 VSUBS 0.005922f
C837 B.n797 VSUBS 0.005922f
C838 B.n798 VSUBS 0.005922f
C839 B.n799 VSUBS 0.005922f
C840 B.n800 VSUBS 0.005922f
C841 B.n801 VSUBS 0.005922f
C842 B.n802 VSUBS 0.005922f
C843 B.n803 VSUBS 0.005922f
C844 B.n804 VSUBS 0.005922f
C845 B.n805 VSUBS 0.005922f
C846 B.n806 VSUBS 0.005922f
C847 B.n807 VSUBS 0.005922f
C848 B.n808 VSUBS 0.005922f
C849 B.n809 VSUBS 0.005922f
C850 B.n810 VSUBS 0.005922f
C851 B.n811 VSUBS 0.005922f
C852 B.n812 VSUBS 0.005922f
C853 B.n813 VSUBS 0.005922f
C854 B.n814 VSUBS 0.005922f
C855 B.n815 VSUBS 0.005922f
C856 B.n816 VSUBS 0.005922f
C857 B.n817 VSUBS 0.005922f
C858 B.n818 VSUBS 0.005922f
C859 B.n819 VSUBS 0.007727f
C860 B.n820 VSUBS 0.008231f
C861 B.n821 VSUBS 0.016369f
C862 VDD1.t2 VSUBS 0.396828f
C863 VDD1.t0 VSUBS 0.396828f
C864 VDD1.n0 VSUBS 3.34265f
C865 VDD1.t1 VSUBS 0.396828f
C866 VDD1.t3 VSUBS 0.396828f
C867 VDD1.n1 VSUBS 4.32733f
C868 VP.t0 VSUBS 4.10695f
C869 VP.n0 VSUBS 1.535f
C870 VP.n1 VSUBS 0.02969f
C871 VP.n2 VSUBS 0.058698f
C872 VP.t3 VSUBS 4.36845f
C873 VP.t1 VSUBS 4.37523f
C874 VP.n3 VSUBS 4.72055f
C875 VP.n4 VSUBS 1.90844f
C876 VP.t2 VSUBS 4.10695f
C877 VP.n5 VSUBS 1.535f
C878 VP.n6 VSUBS 0.055057f
C879 VP.n7 VSUBS 0.047911f
C880 VP.n8 VSUBS 0.02969f
C881 VP.n9 VSUBS 0.02969f
C882 VP.n10 VSUBS 0.023979f
C883 VP.n11 VSUBS 0.058698f
C884 VP.n12 VSUBS 0.055057f
C885 VP.n13 VSUBS 0.047911f
C886 VP.n14 VSUBS 0.052686f
C887 VTAIL.n0 VSUBS 0.012481f
C888 VTAIL.n1 VSUBS 0.028093f
C889 VTAIL.n2 VSUBS 0.012585f
C890 VTAIL.n3 VSUBS 0.022119f
C891 VTAIL.n4 VSUBS 0.011886f
C892 VTAIL.n5 VSUBS 0.028093f
C893 VTAIL.n6 VSUBS 0.012585f
C894 VTAIL.n7 VSUBS 0.022119f
C895 VTAIL.n8 VSUBS 0.011886f
C896 VTAIL.n9 VSUBS 0.028093f
C897 VTAIL.n10 VSUBS 0.012585f
C898 VTAIL.n11 VSUBS 0.022119f
C899 VTAIL.n12 VSUBS 0.011886f
C900 VTAIL.n13 VSUBS 0.028093f
C901 VTAIL.n14 VSUBS 0.012585f
C902 VTAIL.n15 VSUBS 0.022119f
C903 VTAIL.n16 VSUBS 0.011886f
C904 VTAIL.n17 VSUBS 0.028093f
C905 VTAIL.n18 VSUBS 0.012585f
C906 VTAIL.n19 VSUBS 0.022119f
C907 VTAIL.n20 VSUBS 0.011886f
C908 VTAIL.n21 VSUBS 0.028093f
C909 VTAIL.n22 VSUBS 0.012235f
C910 VTAIL.n23 VSUBS 0.022119f
C911 VTAIL.n24 VSUBS 0.012585f
C912 VTAIL.n25 VSUBS 0.028093f
C913 VTAIL.n26 VSUBS 0.012585f
C914 VTAIL.n27 VSUBS 0.022119f
C915 VTAIL.n28 VSUBS 0.011886f
C916 VTAIL.n29 VSUBS 0.028093f
C917 VTAIL.n30 VSUBS 0.012585f
C918 VTAIL.n31 VSUBS 1.74773f
C919 VTAIL.n32 VSUBS 0.011886f
C920 VTAIL.t6 VSUBS 0.061047f
C921 VTAIL.n33 VSUBS 0.242405f
C922 VTAIL.n34 VSUBS 0.021133f
C923 VTAIL.n35 VSUBS 0.02107f
C924 VTAIL.n36 VSUBS 0.028093f
C925 VTAIL.n37 VSUBS 0.012585f
C926 VTAIL.n38 VSUBS 0.011886f
C927 VTAIL.n39 VSUBS 0.022119f
C928 VTAIL.n40 VSUBS 0.022119f
C929 VTAIL.n41 VSUBS 0.011886f
C930 VTAIL.n42 VSUBS 0.012585f
C931 VTAIL.n43 VSUBS 0.028093f
C932 VTAIL.n44 VSUBS 0.028093f
C933 VTAIL.n45 VSUBS 0.012585f
C934 VTAIL.n46 VSUBS 0.011886f
C935 VTAIL.n47 VSUBS 0.022119f
C936 VTAIL.n48 VSUBS 0.022119f
C937 VTAIL.n49 VSUBS 0.011886f
C938 VTAIL.n50 VSUBS 0.011886f
C939 VTAIL.n51 VSUBS 0.012585f
C940 VTAIL.n52 VSUBS 0.028093f
C941 VTAIL.n53 VSUBS 0.028093f
C942 VTAIL.n54 VSUBS 0.028093f
C943 VTAIL.n55 VSUBS 0.012235f
C944 VTAIL.n56 VSUBS 0.011886f
C945 VTAIL.n57 VSUBS 0.022119f
C946 VTAIL.n58 VSUBS 0.022119f
C947 VTAIL.n59 VSUBS 0.011886f
C948 VTAIL.n60 VSUBS 0.012585f
C949 VTAIL.n61 VSUBS 0.028093f
C950 VTAIL.n62 VSUBS 0.028093f
C951 VTAIL.n63 VSUBS 0.012585f
C952 VTAIL.n64 VSUBS 0.011886f
C953 VTAIL.n65 VSUBS 0.022119f
C954 VTAIL.n66 VSUBS 0.022119f
C955 VTAIL.n67 VSUBS 0.011886f
C956 VTAIL.n68 VSUBS 0.012585f
C957 VTAIL.n69 VSUBS 0.028093f
C958 VTAIL.n70 VSUBS 0.028093f
C959 VTAIL.n71 VSUBS 0.012585f
C960 VTAIL.n72 VSUBS 0.011886f
C961 VTAIL.n73 VSUBS 0.022119f
C962 VTAIL.n74 VSUBS 0.022119f
C963 VTAIL.n75 VSUBS 0.011886f
C964 VTAIL.n76 VSUBS 0.012585f
C965 VTAIL.n77 VSUBS 0.028093f
C966 VTAIL.n78 VSUBS 0.028093f
C967 VTAIL.n79 VSUBS 0.012585f
C968 VTAIL.n80 VSUBS 0.011886f
C969 VTAIL.n81 VSUBS 0.022119f
C970 VTAIL.n82 VSUBS 0.022119f
C971 VTAIL.n83 VSUBS 0.011886f
C972 VTAIL.n84 VSUBS 0.012585f
C973 VTAIL.n85 VSUBS 0.028093f
C974 VTAIL.n86 VSUBS 0.028093f
C975 VTAIL.n87 VSUBS 0.012585f
C976 VTAIL.n88 VSUBS 0.011886f
C977 VTAIL.n89 VSUBS 0.022119f
C978 VTAIL.n90 VSUBS 0.022119f
C979 VTAIL.n91 VSUBS 0.011886f
C980 VTAIL.n92 VSUBS 0.012585f
C981 VTAIL.n93 VSUBS 0.028093f
C982 VTAIL.n94 VSUBS 0.028093f
C983 VTAIL.n95 VSUBS 0.012585f
C984 VTAIL.n96 VSUBS 0.011886f
C985 VTAIL.n97 VSUBS 0.022119f
C986 VTAIL.n98 VSUBS 0.057774f
C987 VTAIL.n99 VSUBS 0.011886f
C988 VTAIL.n100 VSUBS 0.012585f
C989 VTAIL.n101 VSUBS 0.064502f
C990 VTAIL.n102 VSUBS 0.042912f
C991 VTAIL.n103 VSUBS 0.152105f
C992 VTAIL.n104 VSUBS 0.012481f
C993 VTAIL.n105 VSUBS 0.028093f
C994 VTAIL.n106 VSUBS 0.012585f
C995 VTAIL.n107 VSUBS 0.022119f
C996 VTAIL.n108 VSUBS 0.011886f
C997 VTAIL.n109 VSUBS 0.028093f
C998 VTAIL.n110 VSUBS 0.012585f
C999 VTAIL.n111 VSUBS 0.022119f
C1000 VTAIL.n112 VSUBS 0.011886f
C1001 VTAIL.n113 VSUBS 0.028093f
C1002 VTAIL.n114 VSUBS 0.012585f
C1003 VTAIL.n115 VSUBS 0.022119f
C1004 VTAIL.n116 VSUBS 0.011886f
C1005 VTAIL.n117 VSUBS 0.028093f
C1006 VTAIL.n118 VSUBS 0.012585f
C1007 VTAIL.n119 VSUBS 0.022119f
C1008 VTAIL.n120 VSUBS 0.011886f
C1009 VTAIL.n121 VSUBS 0.028093f
C1010 VTAIL.n122 VSUBS 0.012585f
C1011 VTAIL.n123 VSUBS 0.022119f
C1012 VTAIL.n124 VSUBS 0.011886f
C1013 VTAIL.n125 VSUBS 0.028093f
C1014 VTAIL.n126 VSUBS 0.012235f
C1015 VTAIL.n127 VSUBS 0.022119f
C1016 VTAIL.n128 VSUBS 0.012585f
C1017 VTAIL.n129 VSUBS 0.028093f
C1018 VTAIL.n130 VSUBS 0.012585f
C1019 VTAIL.n131 VSUBS 0.022119f
C1020 VTAIL.n132 VSUBS 0.011886f
C1021 VTAIL.n133 VSUBS 0.028093f
C1022 VTAIL.n134 VSUBS 0.012585f
C1023 VTAIL.n135 VSUBS 1.74773f
C1024 VTAIL.n136 VSUBS 0.011886f
C1025 VTAIL.t7 VSUBS 0.061047f
C1026 VTAIL.n137 VSUBS 0.242405f
C1027 VTAIL.n138 VSUBS 0.021133f
C1028 VTAIL.n139 VSUBS 0.02107f
C1029 VTAIL.n140 VSUBS 0.028093f
C1030 VTAIL.n141 VSUBS 0.012585f
C1031 VTAIL.n142 VSUBS 0.011886f
C1032 VTAIL.n143 VSUBS 0.022119f
C1033 VTAIL.n144 VSUBS 0.022119f
C1034 VTAIL.n145 VSUBS 0.011886f
C1035 VTAIL.n146 VSUBS 0.012585f
C1036 VTAIL.n147 VSUBS 0.028093f
C1037 VTAIL.n148 VSUBS 0.028093f
C1038 VTAIL.n149 VSUBS 0.012585f
C1039 VTAIL.n150 VSUBS 0.011886f
C1040 VTAIL.n151 VSUBS 0.022119f
C1041 VTAIL.n152 VSUBS 0.022119f
C1042 VTAIL.n153 VSUBS 0.011886f
C1043 VTAIL.n154 VSUBS 0.011886f
C1044 VTAIL.n155 VSUBS 0.012585f
C1045 VTAIL.n156 VSUBS 0.028093f
C1046 VTAIL.n157 VSUBS 0.028093f
C1047 VTAIL.n158 VSUBS 0.028093f
C1048 VTAIL.n159 VSUBS 0.012235f
C1049 VTAIL.n160 VSUBS 0.011886f
C1050 VTAIL.n161 VSUBS 0.022119f
C1051 VTAIL.n162 VSUBS 0.022119f
C1052 VTAIL.n163 VSUBS 0.011886f
C1053 VTAIL.n164 VSUBS 0.012585f
C1054 VTAIL.n165 VSUBS 0.028093f
C1055 VTAIL.n166 VSUBS 0.028093f
C1056 VTAIL.n167 VSUBS 0.012585f
C1057 VTAIL.n168 VSUBS 0.011886f
C1058 VTAIL.n169 VSUBS 0.022119f
C1059 VTAIL.n170 VSUBS 0.022119f
C1060 VTAIL.n171 VSUBS 0.011886f
C1061 VTAIL.n172 VSUBS 0.012585f
C1062 VTAIL.n173 VSUBS 0.028093f
C1063 VTAIL.n174 VSUBS 0.028093f
C1064 VTAIL.n175 VSUBS 0.012585f
C1065 VTAIL.n176 VSUBS 0.011886f
C1066 VTAIL.n177 VSUBS 0.022119f
C1067 VTAIL.n178 VSUBS 0.022119f
C1068 VTAIL.n179 VSUBS 0.011886f
C1069 VTAIL.n180 VSUBS 0.012585f
C1070 VTAIL.n181 VSUBS 0.028093f
C1071 VTAIL.n182 VSUBS 0.028093f
C1072 VTAIL.n183 VSUBS 0.012585f
C1073 VTAIL.n184 VSUBS 0.011886f
C1074 VTAIL.n185 VSUBS 0.022119f
C1075 VTAIL.n186 VSUBS 0.022119f
C1076 VTAIL.n187 VSUBS 0.011886f
C1077 VTAIL.n188 VSUBS 0.012585f
C1078 VTAIL.n189 VSUBS 0.028093f
C1079 VTAIL.n190 VSUBS 0.028093f
C1080 VTAIL.n191 VSUBS 0.012585f
C1081 VTAIL.n192 VSUBS 0.011886f
C1082 VTAIL.n193 VSUBS 0.022119f
C1083 VTAIL.n194 VSUBS 0.022119f
C1084 VTAIL.n195 VSUBS 0.011886f
C1085 VTAIL.n196 VSUBS 0.012585f
C1086 VTAIL.n197 VSUBS 0.028093f
C1087 VTAIL.n198 VSUBS 0.028093f
C1088 VTAIL.n199 VSUBS 0.012585f
C1089 VTAIL.n200 VSUBS 0.011886f
C1090 VTAIL.n201 VSUBS 0.022119f
C1091 VTAIL.n202 VSUBS 0.057774f
C1092 VTAIL.n203 VSUBS 0.011886f
C1093 VTAIL.n204 VSUBS 0.012585f
C1094 VTAIL.n205 VSUBS 0.064502f
C1095 VTAIL.n206 VSUBS 0.042912f
C1096 VTAIL.n207 VSUBS 0.240119f
C1097 VTAIL.n208 VSUBS 0.012481f
C1098 VTAIL.n209 VSUBS 0.028093f
C1099 VTAIL.n210 VSUBS 0.012585f
C1100 VTAIL.n211 VSUBS 0.022119f
C1101 VTAIL.n212 VSUBS 0.011886f
C1102 VTAIL.n213 VSUBS 0.028093f
C1103 VTAIL.n214 VSUBS 0.012585f
C1104 VTAIL.n215 VSUBS 0.022119f
C1105 VTAIL.n216 VSUBS 0.011886f
C1106 VTAIL.n217 VSUBS 0.028093f
C1107 VTAIL.n218 VSUBS 0.012585f
C1108 VTAIL.n219 VSUBS 0.022119f
C1109 VTAIL.n220 VSUBS 0.011886f
C1110 VTAIL.n221 VSUBS 0.028093f
C1111 VTAIL.n222 VSUBS 0.012585f
C1112 VTAIL.n223 VSUBS 0.022119f
C1113 VTAIL.n224 VSUBS 0.011886f
C1114 VTAIL.n225 VSUBS 0.028093f
C1115 VTAIL.n226 VSUBS 0.012585f
C1116 VTAIL.n227 VSUBS 0.022119f
C1117 VTAIL.n228 VSUBS 0.011886f
C1118 VTAIL.n229 VSUBS 0.028093f
C1119 VTAIL.n230 VSUBS 0.012235f
C1120 VTAIL.n231 VSUBS 0.022119f
C1121 VTAIL.n232 VSUBS 0.012585f
C1122 VTAIL.n233 VSUBS 0.028093f
C1123 VTAIL.n234 VSUBS 0.012585f
C1124 VTAIL.n235 VSUBS 0.022119f
C1125 VTAIL.n236 VSUBS 0.011886f
C1126 VTAIL.n237 VSUBS 0.028093f
C1127 VTAIL.n238 VSUBS 0.012585f
C1128 VTAIL.n239 VSUBS 1.74773f
C1129 VTAIL.n240 VSUBS 0.011886f
C1130 VTAIL.t0 VSUBS 0.061047f
C1131 VTAIL.n241 VSUBS 0.242405f
C1132 VTAIL.n242 VSUBS 0.021133f
C1133 VTAIL.n243 VSUBS 0.02107f
C1134 VTAIL.n244 VSUBS 0.028093f
C1135 VTAIL.n245 VSUBS 0.012585f
C1136 VTAIL.n246 VSUBS 0.011886f
C1137 VTAIL.n247 VSUBS 0.022119f
C1138 VTAIL.n248 VSUBS 0.022119f
C1139 VTAIL.n249 VSUBS 0.011886f
C1140 VTAIL.n250 VSUBS 0.012585f
C1141 VTAIL.n251 VSUBS 0.028093f
C1142 VTAIL.n252 VSUBS 0.028093f
C1143 VTAIL.n253 VSUBS 0.012585f
C1144 VTAIL.n254 VSUBS 0.011886f
C1145 VTAIL.n255 VSUBS 0.022119f
C1146 VTAIL.n256 VSUBS 0.022119f
C1147 VTAIL.n257 VSUBS 0.011886f
C1148 VTAIL.n258 VSUBS 0.011886f
C1149 VTAIL.n259 VSUBS 0.012585f
C1150 VTAIL.n260 VSUBS 0.028093f
C1151 VTAIL.n261 VSUBS 0.028093f
C1152 VTAIL.n262 VSUBS 0.028093f
C1153 VTAIL.n263 VSUBS 0.012235f
C1154 VTAIL.n264 VSUBS 0.011886f
C1155 VTAIL.n265 VSUBS 0.022119f
C1156 VTAIL.n266 VSUBS 0.022119f
C1157 VTAIL.n267 VSUBS 0.011886f
C1158 VTAIL.n268 VSUBS 0.012585f
C1159 VTAIL.n269 VSUBS 0.028093f
C1160 VTAIL.n270 VSUBS 0.028093f
C1161 VTAIL.n271 VSUBS 0.012585f
C1162 VTAIL.n272 VSUBS 0.011886f
C1163 VTAIL.n273 VSUBS 0.022119f
C1164 VTAIL.n274 VSUBS 0.022119f
C1165 VTAIL.n275 VSUBS 0.011886f
C1166 VTAIL.n276 VSUBS 0.012585f
C1167 VTAIL.n277 VSUBS 0.028093f
C1168 VTAIL.n278 VSUBS 0.028093f
C1169 VTAIL.n279 VSUBS 0.012585f
C1170 VTAIL.n280 VSUBS 0.011886f
C1171 VTAIL.n281 VSUBS 0.022119f
C1172 VTAIL.n282 VSUBS 0.022119f
C1173 VTAIL.n283 VSUBS 0.011886f
C1174 VTAIL.n284 VSUBS 0.012585f
C1175 VTAIL.n285 VSUBS 0.028093f
C1176 VTAIL.n286 VSUBS 0.028093f
C1177 VTAIL.n287 VSUBS 0.012585f
C1178 VTAIL.n288 VSUBS 0.011886f
C1179 VTAIL.n289 VSUBS 0.022119f
C1180 VTAIL.n290 VSUBS 0.022119f
C1181 VTAIL.n291 VSUBS 0.011886f
C1182 VTAIL.n292 VSUBS 0.012585f
C1183 VTAIL.n293 VSUBS 0.028093f
C1184 VTAIL.n294 VSUBS 0.028093f
C1185 VTAIL.n295 VSUBS 0.012585f
C1186 VTAIL.n296 VSUBS 0.011886f
C1187 VTAIL.n297 VSUBS 0.022119f
C1188 VTAIL.n298 VSUBS 0.022119f
C1189 VTAIL.n299 VSUBS 0.011886f
C1190 VTAIL.n300 VSUBS 0.012585f
C1191 VTAIL.n301 VSUBS 0.028093f
C1192 VTAIL.n302 VSUBS 0.028093f
C1193 VTAIL.n303 VSUBS 0.012585f
C1194 VTAIL.n304 VSUBS 0.011886f
C1195 VTAIL.n305 VSUBS 0.022119f
C1196 VTAIL.n306 VSUBS 0.057774f
C1197 VTAIL.n307 VSUBS 0.011886f
C1198 VTAIL.n308 VSUBS 0.012585f
C1199 VTAIL.n309 VSUBS 0.064502f
C1200 VTAIL.n310 VSUBS 0.042912f
C1201 VTAIL.n311 VSUBS 1.84773f
C1202 VTAIL.n312 VSUBS 0.012481f
C1203 VTAIL.n313 VSUBS 0.028093f
C1204 VTAIL.n314 VSUBS 0.012585f
C1205 VTAIL.n315 VSUBS 0.022119f
C1206 VTAIL.n316 VSUBS 0.011886f
C1207 VTAIL.n317 VSUBS 0.028093f
C1208 VTAIL.n318 VSUBS 0.012585f
C1209 VTAIL.n319 VSUBS 0.022119f
C1210 VTAIL.n320 VSUBS 0.011886f
C1211 VTAIL.n321 VSUBS 0.028093f
C1212 VTAIL.n322 VSUBS 0.012585f
C1213 VTAIL.n323 VSUBS 0.022119f
C1214 VTAIL.n324 VSUBS 0.011886f
C1215 VTAIL.n325 VSUBS 0.028093f
C1216 VTAIL.n326 VSUBS 0.012585f
C1217 VTAIL.n327 VSUBS 0.022119f
C1218 VTAIL.n328 VSUBS 0.011886f
C1219 VTAIL.n329 VSUBS 0.028093f
C1220 VTAIL.n330 VSUBS 0.012585f
C1221 VTAIL.n331 VSUBS 0.022119f
C1222 VTAIL.n332 VSUBS 0.011886f
C1223 VTAIL.n333 VSUBS 0.028093f
C1224 VTAIL.n334 VSUBS 0.012235f
C1225 VTAIL.n335 VSUBS 0.022119f
C1226 VTAIL.n336 VSUBS 0.012235f
C1227 VTAIL.n337 VSUBS 0.011886f
C1228 VTAIL.n338 VSUBS 0.028093f
C1229 VTAIL.n339 VSUBS 0.028093f
C1230 VTAIL.n340 VSUBS 0.012585f
C1231 VTAIL.n341 VSUBS 0.022119f
C1232 VTAIL.n342 VSUBS 0.011886f
C1233 VTAIL.n343 VSUBS 0.028093f
C1234 VTAIL.n344 VSUBS 0.012585f
C1235 VTAIL.n345 VSUBS 1.74773f
C1236 VTAIL.n346 VSUBS 0.011886f
C1237 VTAIL.t4 VSUBS 0.061047f
C1238 VTAIL.n347 VSUBS 0.242405f
C1239 VTAIL.n348 VSUBS 0.021133f
C1240 VTAIL.n349 VSUBS 0.02107f
C1241 VTAIL.n350 VSUBS 0.028093f
C1242 VTAIL.n351 VSUBS 0.012585f
C1243 VTAIL.n352 VSUBS 0.011886f
C1244 VTAIL.n353 VSUBS 0.022119f
C1245 VTAIL.n354 VSUBS 0.022119f
C1246 VTAIL.n355 VSUBS 0.011886f
C1247 VTAIL.n356 VSUBS 0.012585f
C1248 VTAIL.n357 VSUBS 0.028093f
C1249 VTAIL.n358 VSUBS 0.028093f
C1250 VTAIL.n359 VSUBS 0.012585f
C1251 VTAIL.n360 VSUBS 0.011886f
C1252 VTAIL.n361 VSUBS 0.022119f
C1253 VTAIL.n362 VSUBS 0.022119f
C1254 VTAIL.n363 VSUBS 0.011886f
C1255 VTAIL.n364 VSUBS 0.012585f
C1256 VTAIL.n365 VSUBS 0.028093f
C1257 VTAIL.n366 VSUBS 0.028093f
C1258 VTAIL.n367 VSUBS 0.012585f
C1259 VTAIL.n368 VSUBS 0.011886f
C1260 VTAIL.n369 VSUBS 0.022119f
C1261 VTAIL.n370 VSUBS 0.022119f
C1262 VTAIL.n371 VSUBS 0.011886f
C1263 VTAIL.n372 VSUBS 0.012585f
C1264 VTAIL.n373 VSUBS 0.028093f
C1265 VTAIL.n374 VSUBS 0.028093f
C1266 VTAIL.n375 VSUBS 0.012585f
C1267 VTAIL.n376 VSUBS 0.011886f
C1268 VTAIL.n377 VSUBS 0.022119f
C1269 VTAIL.n378 VSUBS 0.022119f
C1270 VTAIL.n379 VSUBS 0.011886f
C1271 VTAIL.n380 VSUBS 0.012585f
C1272 VTAIL.n381 VSUBS 0.028093f
C1273 VTAIL.n382 VSUBS 0.028093f
C1274 VTAIL.n383 VSUBS 0.012585f
C1275 VTAIL.n384 VSUBS 0.011886f
C1276 VTAIL.n385 VSUBS 0.022119f
C1277 VTAIL.n386 VSUBS 0.022119f
C1278 VTAIL.n387 VSUBS 0.011886f
C1279 VTAIL.n388 VSUBS 0.012585f
C1280 VTAIL.n389 VSUBS 0.028093f
C1281 VTAIL.n390 VSUBS 0.028093f
C1282 VTAIL.n391 VSUBS 0.012585f
C1283 VTAIL.n392 VSUBS 0.011886f
C1284 VTAIL.n393 VSUBS 0.022119f
C1285 VTAIL.n394 VSUBS 0.022119f
C1286 VTAIL.n395 VSUBS 0.011886f
C1287 VTAIL.n396 VSUBS 0.012585f
C1288 VTAIL.n397 VSUBS 0.028093f
C1289 VTAIL.n398 VSUBS 0.028093f
C1290 VTAIL.n399 VSUBS 0.012585f
C1291 VTAIL.n400 VSUBS 0.011886f
C1292 VTAIL.n401 VSUBS 0.022119f
C1293 VTAIL.n402 VSUBS 0.022119f
C1294 VTAIL.n403 VSUBS 0.011886f
C1295 VTAIL.n404 VSUBS 0.012585f
C1296 VTAIL.n405 VSUBS 0.028093f
C1297 VTAIL.n406 VSUBS 0.028093f
C1298 VTAIL.n407 VSUBS 0.012585f
C1299 VTAIL.n408 VSUBS 0.011886f
C1300 VTAIL.n409 VSUBS 0.022119f
C1301 VTAIL.n410 VSUBS 0.057774f
C1302 VTAIL.n411 VSUBS 0.011886f
C1303 VTAIL.n412 VSUBS 0.012585f
C1304 VTAIL.n413 VSUBS 0.064502f
C1305 VTAIL.n414 VSUBS 0.042912f
C1306 VTAIL.n415 VSUBS 1.84773f
C1307 VTAIL.n416 VSUBS 0.012481f
C1308 VTAIL.n417 VSUBS 0.028093f
C1309 VTAIL.n418 VSUBS 0.012585f
C1310 VTAIL.n419 VSUBS 0.022119f
C1311 VTAIL.n420 VSUBS 0.011886f
C1312 VTAIL.n421 VSUBS 0.028093f
C1313 VTAIL.n422 VSUBS 0.012585f
C1314 VTAIL.n423 VSUBS 0.022119f
C1315 VTAIL.n424 VSUBS 0.011886f
C1316 VTAIL.n425 VSUBS 0.028093f
C1317 VTAIL.n426 VSUBS 0.012585f
C1318 VTAIL.n427 VSUBS 0.022119f
C1319 VTAIL.n428 VSUBS 0.011886f
C1320 VTAIL.n429 VSUBS 0.028093f
C1321 VTAIL.n430 VSUBS 0.012585f
C1322 VTAIL.n431 VSUBS 0.022119f
C1323 VTAIL.n432 VSUBS 0.011886f
C1324 VTAIL.n433 VSUBS 0.028093f
C1325 VTAIL.n434 VSUBS 0.012585f
C1326 VTAIL.n435 VSUBS 0.022119f
C1327 VTAIL.n436 VSUBS 0.011886f
C1328 VTAIL.n437 VSUBS 0.028093f
C1329 VTAIL.n438 VSUBS 0.012235f
C1330 VTAIL.n439 VSUBS 0.022119f
C1331 VTAIL.n440 VSUBS 0.012235f
C1332 VTAIL.n441 VSUBS 0.011886f
C1333 VTAIL.n442 VSUBS 0.028093f
C1334 VTAIL.n443 VSUBS 0.028093f
C1335 VTAIL.n444 VSUBS 0.012585f
C1336 VTAIL.n445 VSUBS 0.022119f
C1337 VTAIL.n446 VSUBS 0.011886f
C1338 VTAIL.n447 VSUBS 0.028093f
C1339 VTAIL.n448 VSUBS 0.012585f
C1340 VTAIL.n449 VSUBS 1.74773f
C1341 VTAIL.n450 VSUBS 0.011886f
C1342 VTAIL.t5 VSUBS 0.061047f
C1343 VTAIL.n451 VSUBS 0.242405f
C1344 VTAIL.n452 VSUBS 0.021133f
C1345 VTAIL.n453 VSUBS 0.02107f
C1346 VTAIL.n454 VSUBS 0.028093f
C1347 VTAIL.n455 VSUBS 0.012585f
C1348 VTAIL.n456 VSUBS 0.011886f
C1349 VTAIL.n457 VSUBS 0.022119f
C1350 VTAIL.n458 VSUBS 0.022119f
C1351 VTAIL.n459 VSUBS 0.011886f
C1352 VTAIL.n460 VSUBS 0.012585f
C1353 VTAIL.n461 VSUBS 0.028093f
C1354 VTAIL.n462 VSUBS 0.028093f
C1355 VTAIL.n463 VSUBS 0.012585f
C1356 VTAIL.n464 VSUBS 0.011886f
C1357 VTAIL.n465 VSUBS 0.022119f
C1358 VTAIL.n466 VSUBS 0.022119f
C1359 VTAIL.n467 VSUBS 0.011886f
C1360 VTAIL.n468 VSUBS 0.012585f
C1361 VTAIL.n469 VSUBS 0.028093f
C1362 VTAIL.n470 VSUBS 0.028093f
C1363 VTAIL.n471 VSUBS 0.012585f
C1364 VTAIL.n472 VSUBS 0.011886f
C1365 VTAIL.n473 VSUBS 0.022119f
C1366 VTAIL.n474 VSUBS 0.022119f
C1367 VTAIL.n475 VSUBS 0.011886f
C1368 VTAIL.n476 VSUBS 0.012585f
C1369 VTAIL.n477 VSUBS 0.028093f
C1370 VTAIL.n478 VSUBS 0.028093f
C1371 VTAIL.n479 VSUBS 0.012585f
C1372 VTAIL.n480 VSUBS 0.011886f
C1373 VTAIL.n481 VSUBS 0.022119f
C1374 VTAIL.n482 VSUBS 0.022119f
C1375 VTAIL.n483 VSUBS 0.011886f
C1376 VTAIL.n484 VSUBS 0.012585f
C1377 VTAIL.n485 VSUBS 0.028093f
C1378 VTAIL.n486 VSUBS 0.028093f
C1379 VTAIL.n487 VSUBS 0.012585f
C1380 VTAIL.n488 VSUBS 0.011886f
C1381 VTAIL.n489 VSUBS 0.022119f
C1382 VTAIL.n490 VSUBS 0.022119f
C1383 VTAIL.n491 VSUBS 0.011886f
C1384 VTAIL.n492 VSUBS 0.012585f
C1385 VTAIL.n493 VSUBS 0.028093f
C1386 VTAIL.n494 VSUBS 0.028093f
C1387 VTAIL.n495 VSUBS 0.012585f
C1388 VTAIL.n496 VSUBS 0.011886f
C1389 VTAIL.n497 VSUBS 0.022119f
C1390 VTAIL.n498 VSUBS 0.022119f
C1391 VTAIL.n499 VSUBS 0.011886f
C1392 VTAIL.n500 VSUBS 0.012585f
C1393 VTAIL.n501 VSUBS 0.028093f
C1394 VTAIL.n502 VSUBS 0.028093f
C1395 VTAIL.n503 VSUBS 0.012585f
C1396 VTAIL.n504 VSUBS 0.011886f
C1397 VTAIL.n505 VSUBS 0.022119f
C1398 VTAIL.n506 VSUBS 0.022119f
C1399 VTAIL.n507 VSUBS 0.011886f
C1400 VTAIL.n508 VSUBS 0.012585f
C1401 VTAIL.n509 VSUBS 0.028093f
C1402 VTAIL.n510 VSUBS 0.028093f
C1403 VTAIL.n511 VSUBS 0.012585f
C1404 VTAIL.n512 VSUBS 0.011886f
C1405 VTAIL.n513 VSUBS 0.022119f
C1406 VTAIL.n514 VSUBS 0.057774f
C1407 VTAIL.n515 VSUBS 0.011886f
C1408 VTAIL.n516 VSUBS 0.012585f
C1409 VTAIL.n517 VSUBS 0.064502f
C1410 VTAIL.n518 VSUBS 0.042912f
C1411 VTAIL.n519 VSUBS 0.240119f
C1412 VTAIL.n520 VSUBS 0.012481f
C1413 VTAIL.n521 VSUBS 0.028093f
C1414 VTAIL.n522 VSUBS 0.012585f
C1415 VTAIL.n523 VSUBS 0.022119f
C1416 VTAIL.n524 VSUBS 0.011886f
C1417 VTAIL.n525 VSUBS 0.028093f
C1418 VTAIL.n526 VSUBS 0.012585f
C1419 VTAIL.n527 VSUBS 0.022119f
C1420 VTAIL.n528 VSUBS 0.011886f
C1421 VTAIL.n529 VSUBS 0.028093f
C1422 VTAIL.n530 VSUBS 0.012585f
C1423 VTAIL.n531 VSUBS 0.022119f
C1424 VTAIL.n532 VSUBS 0.011886f
C1425 VTAIL.n533 VSUBS 0.028093f
C1426 VTAIL.n534 VSUBS 0.012585f
C1427 VTAIL.n535 VSUBS 0.022119f
C1428 VTAIL.n536 VSUBS 0.011886f
C1429 VTAIL.n537 VSUBS 0.028093f
C1430 VTAIL.n538 VSUBS 0.012585f
C1431 VTAIL.n539 VSUBS 0.022119f
C1432 VTAIL.n540 VSUBS 0.011886f
C1433 VTAIL.n541 VSUBS 0.028093f
C1434 VTAIL.n542 VSUBS 0.012235f
C1435 VTAIL.n543 VSUBS 0.022119f
C1436 VTAIL.n544 VSUBS 0.012235f
C1437 VTAIL.n545 VSUBS 0.011886f
C1438 VTAIL.n546 VSUBS 0.028093f
C1439 VTAIL.n547 VSUBS 0.028093f
C1440 VTAIL.n548 VSUBS 0.012585f
C1441 VTAIL.n549 VSUBS 0.022119f
C1442 VTAIL.n550 VSUBS 0.011886f
C1443 VTAIL.n551 VSUBS 0.028093f
C1444 VTAIL.n552 VSUBS 0.012585f
C1445 VTAIL.n553 VSUBS 1.74773f
C1446 VTAIL.n554 VSUBS 0.011886f
C1447 VTAIL.t2 VSUBS 0.061047f
C1448 VTAIL.n555 VSUBS 0.242405f
C1449 VTAIL.n556 VSUBS 0.021133f
C1450 VTAIL.n557 VSUBS 0.02107f
C1451 VTAIL.n558 VSUBS 0.028093f
C1452 VTAIL.n559 VSUBS 0.012585f
C1453 VTAIL.n560 VSUBS 0.011886f
C1454 VTAIL.n561 VSUBS 0.022119f
C1455 VTAIL.n562 VSUBS 0.022119f
C1456 VTAIL.n563 VSUBS 0.011886f
C1457 VTAIL.n564 VSUBS 0.012585f
C1458 VTAIL.n565 VSUBS 0.028093f
C1459 VTAIL.n566 VSUBS 0.028093f
C1460 VTAIL.n567 VSUBS 0.012585f
C1461 VTAIL.n568 VSUBS 0.011886f
C1462 VTAIL.n569 VSUBS 0.022119f
C1463 VTAIL.n570 VSUBS 0.022119f
C1464 VTAIL.n571 VSUBS 0.011886f
C1465 VTAIL.n572 VSUBS 0.012585f
C1466 VTAIL.n573 VSUBS 0.028093f
C1467 VTAIL.n574 VSUBS 0.028093f
C1468 VTAIL.n575 VSUBS 0.012585f
C1469 VTAIL.n576 VSUBS 0.011886f
C1470 VTAIL.n577 VSUBS 0.022119f
C1471 VTAIL.n578 VSUBS 0.022119f
C1472 VTAIL.n579 VSUBS 0.011886f
C1473 VTAIL.n580 VSUBS 0.012585f
C1474 VTAIL.n581 VSUBS 0.028093f
C1475 VTAIL.n582 VSUBS 0.028093f
C1476 VTAIL.n583 VSUBS 0.012585f
C1477 VTAIL.n584 VSUBS 0.011886f
C1478 VTAIL.n585 VSUBS 0.022119f
C1479 VTAIL.n586 VSUBS 0.022119f
C1480 VTAIL.n587 VSUBS 0.011886f
C1481 VTAIL.n588 VSUBS 0.012585f
C1482 VTAIL.n589 VSUBS 0.028093f
C1483 VTAIL.n590 VSUBS 0.028093f
C1484 VTAIL.n591 VSUBS 0.012585f
C1485 VTAIL.n592 VSUBS 0.011886f
C1486 VTAIL.n593 VSUBS 0.022119f
C1487 VTAIL.n594 VSUBS 0.022119f
C1488 VTAIL.n595 VSUBS 0.011886f
C1489 VTAIL.n596 VSUBS 0.012585f
C1490 VTAIL.n597 VSUBS 0.028093f
C1491 VTAIL.n598 VSUBS 0.028093f
C1492 VTAIL.n599 VSUBS 0.012585f
C1493 VTAIL.n600 VSUBS 0.011886f
C1494 VTAIL.n601 VSUBS 0.022119f
C1495 VTAIL.n602 VSUBS 0.022119f
C1496 VTAIL.n603 VSUBS 0.011886f
C1497 VTAIL.n604 VSUBS 0.012585f
C1498 VTAIL.n605 VSUBS 0.028093f
C1499 VTAIL.n606 VSUBS 0.028093f
C1500 VTAIL.n607 VSUBS 0.012585f
C1501 VTAIL.n608 VSUBS 0.011886f
C1502 VTAIL.n609 VSUBS 0.022119f
C1503 VTAIL.n610 VSUBS 0.022119f
C1504 VTAIL.n611 VSUBS 0.011886f
C1505 VTAIL.n612 VSUBS 0.012585f
C1506 VTAIL.n613 VSUBS 0.028093f
C1507 VTAIL.n614 VSUBS 0.028093f
C1508 VTAIL.n615 VSUBS 0.012585f
C1509 VTAIL.n616 VSUBS 0.011886f
C1510 VTAIL.n617 VSUBS 0.022119f
C1511 VTAIL.n618 VSUBS 0.057774f
C1512 VTAIL.n619 VSUBS 0.011886f
C1513 VTAIL.n620 VSUBS 0.012585f
C1514 VTAIL.n621 VSUBS 0.064502f
C1515 VTAIL.n622 VSUBS 0.042912f
C1516 VTAIL.n623 VSUBS 0.240119f
C1517 VTAIL.n624 VSUBS 0.012481f
C1518 VTAIL.n625 VSUBS 0.028093f
C1519 VTAIL.n626 VSUBS 0.012585f
C1520 VTAIL.n627 VSUBS 0.022119f
C1521 VTAIL.n628 VSUBS 0.011886f
C1522 VTAIL.n629 VSUBS 0.028093f
C1523 VTAIL.n630 VSUBS 0.012585f
C1524 VTAIL.n631 VSUBS 0.022119f
C1525 VTAIL.n632 VSUBS 0.011886f
C1526 VTAIL.n633 VSUBS 0.028093f
C1527 VTAIL.n634 VSUBS 0.012585f
C1528 VTAIL.n635 VSUBS 0.022119f
C1529 VTAIL.n636 VSUBS 0.011886f
C1530 VTAIL.n637 VSUBS 0.028093f
C1531 VTAIL.n638 VSUBS 0.012585f
C1532 VTAIL.n639 VSUBS 0.022119f
C1533 VTAIL.n640 VSUBS 0.011886f
C1534 VTAIL.n641 VSUBS 0.028093f
C1535 VTAIL.n642 VSUBS 0.012585f
C1536 VTAIL.n643 VSUBS 0.022119f
C1537 VTAIL.n644 VSUBS 0.011886f
C1538 VTAIL.n645 VSUBS 0.028093f
C1539 VTAIL.n646 VSUBS 0.012235f
C1540 VTAIL.n647 VSUBS 0.022119f
C1541 VTAIL.n648 VSUBS 0.012235f
C1542 VTAIL.n649 VSUBS 0.011886f
C1543 VTAIL.n650 VSUBS 0.028093f
C1544 VTAIL.n651 VSUBS 0.028093f
C1545 VTAIL.n652 VSUBS 0.012585f
C1546 VTAIL.n653 VSUBS 0.022119f
C1547 VTAIL.n654 VSUBS 0.011886f
C1548 VTAIL.n655 VSUBS 0.028093f
C1549 VTAIL.n656 VSUBS 0.012585f
C1550 VTAIL.n657 VSUBS 1.74773f
C1551 VTAIL.n658 VSUBS 0.011886f
C1552 VTAIL.t1 VSUBS 0.061047f
C1553 VTAIL.n659 VSUBS 0.242405f
C1554 VTAIL.n660 VSUBS 0.021133f
C1555 VTAIL.n661 VSUBS 0.02107f
C1556 VTAIL.n662 VSUBS 0.028093f
C1557 VTAIL.n663 VSUBS 0.012585f
C1558 VTAIL.n664 VSUBS 0.011886f
C1559 VTAIL.n665 VSUBS 0.022119f
C1560 VTAIL.n666 VSUBS 0.022119f
C1561 VTAIL.n667 VSUBS 0.011886f
C1562 VTAIL.n668 VSUBS 0.012585f
C1563 VTAIL.n669 VSUBS 0.028093f
C1564 VTAIL.n670 VSUBS 0.028093f
C1565 VTAIL.n671 VSUBS 0.012585f
C1566 VTAIL.n672 VSUBS 0.011886f
C1567 VTAIL.n673 VSUBS 0.022119f
C1568 VTAIL.n674 VSUBS 0.022119f
C1569 VTAIL.n675 VSUBS 0.011886f
C1570 VTAIL.n676 VSUBS 0.012585f
C1571 VTAIL.n677 VSUBS 0.028093f
C1572 VTAIL.n678 VSUBS 0.028093f
C1573 VTAIL.n679 VSUBS 0.012585f
C1574 VTAIL.n680 VSUBS 0.011886f
C1575 VTAIL.n681 VSUBS 0.022119f
C1576 VTAIL.n682 VSUBS 0.022119f
C1577 VTAIL.n683 VSUBS 0.011886f
C1578 VTAIL.n684 VSUBS 0.012585f
C1579 VTAIL.n685 VSUBS 0.028093f
C1580 VTAIL.n686 VSUBS 0.028093f
C1581 VTAIL.n687 VSUBS 0.012585f
C1582 VTAIL.n688 VSUBS 0.011886f
C1583 VTAIL.n689 VSUBS 0.022119f
C1584 VTAIL.n690 VSUBS 0.022119f
C1585 VTAIL.n691 VSUBS 0.011886f
C1586 VTAIL.n692 VSUBS 0.012585f
C1587 VTAIL.n693 VSUBS 0.028093f
C1588 VTAIL.n694 VSUBS 0.028093f
C1589 VTAIL.n695 VSUBS 0.012585f
C1590 VTAIL.n696 VSUBS 0.011886f
C1591 VTAIL.n697 VSUBS 0.022119f
C1592 VTAIL.n698 VSUBS 0.022119f
C1593 VTAIL.n699 VSUBS 0.011886f
C1594 VTAIL.n700 VSUBS 0.012585f
C1595 VTAIL.n701 VSUBS 0.028093f
C1596 VTAIL.n702 VSUBS 0.028093f
C1597 VTAIL.n703 VSUBS 0.012585f
C1598 VTAIL.n704 VSUBS 0.011886f
C1599 VTAIL.n705 VSUBS 0.022119f
C1600 VTAIL.n706 VSUBS 0.022119f
C1601 VTAIL.n707 VSUBS 0.011886f
C1602 VTAIL.n708 VSUBS 0.012585f
C1603 VTAIL.n709 VSUBS 0.028093f
C1604 VTAIL.n710 VSUBS 0.028093f
C1605 VTAIL.n711 VSUBS 0.012585f
C1606 VTAIL.n712 VSUBS 0.011886f
C1607 VTAIL.n713 VSUBS 0.022119f
C1608 VTAIL.n714 VSUBS 0.022119f
C1609 VTAIL.n715 VSUBS 0.011886f
C1610 VTAIL.n716 VSUBS 0.012585f
C1611 VTAIL.n717 VSUBS 0.028093f
C1612 VTAIL.n718 VSUBS 0.028093f
C1613 VTAIL.n719 VSUBS 0.012585f
C1614 VTAIL.n720 VSUBS 0.011886f
C1615 VTAIL.n721 VSUBS 0.022119f
C1616 VTAIL.n722 VSUBS 0.057774f
C1617 VTAIL.n723 VSUBS 0.011886f
C1618 VTAIL.n724 VSUBS 0.012585f
C1619 VTAIL.n725 VSUBS 0.064502f
C1620 VTAIL.n726 VSUBS 0.042912f
C1621 VTAIL.n727 VSUBS 1.84773f
C1622 VTAIL.n728 VSUBS 0.012481f
C1623 VTAIL.n729 VSUBS 0.028093f
C1624 VTAIL.n730 VSUBS 0.012585f
C1625 VTAIL.n731 VSUBS 0.022119f
C1626 VTAIL.n732 VSUBS 0.011886f
C1627 VTAIL.n733 VSUBS 0.028093f
C1628 VTAIL.n734 VSUBS 0.012585f
C1629 VTAIL.n735 VSUBS 0.022119f
C1630 VTAIL.n736 VSUBS 0.011886f
C1631 VTAIL.n737 VSUBS 0.028093f
C1632 VTAIL.n738 VSUBS 0.012585f
C1633 VTAIL.n739 VSUBS 0.022119f
C1634 VTAIL.n740 VSUBS 0.011886f
C1635 VTAIL.n741 VSUBS 0.028093f
C1636 VTAIL.n742 VSUBS 0.012585f
C1637 VTAIL.n743 VSUBS 0.022119f
C1638 VTAIL.n744 VSUBS 0.011886f
C1639 VTAIL.n745 VSUBS 0.028093f
C1640 VTAIL.n746 VSUBS 0.012585f
C1641 VTAIL.n747 VSUBS 0.022119f
C1642 VTAIL.n748 VSUBS 0.011886f
C1643 VTAIL.n749 VSUBS 0.028093f
C1644 VTAIL.n750 VSUBS 0.012235f
C1645 VTAIL.n751 VSUBS 0.022119f
C1646 VTAIL.n752 VSUBS 0.012585f
C1647 VTAIL.n753 VSUBS 0.028093f
C1648 VTAIL.n754 VSUBS 0.012585f
C1649 VTAIL.n755 VSUBS 0.022119f
C1650 VTAIL.n756 VSUBS 0.011886f
C1651 VTAIL.n757 VSUBS 0.028093f
C1652 VTAIL.n758 VSUBS 0.012585f
C1653 VTAIL.n759 VSUBS 1.74773f
C1654 VTAIL.n760 VSUBS 0.011886f
C1655 VTAIL.t3 VSUBS 0.061047f
C1656 VTAIL.n761 VSUBS 0.242405f
C1657 VTAIL.n762 VSUBS 0.021133f
C1658 VTAIL.n763 VSUBS 0.02107f
C1659 VTAIL.n764 VSUBS 0.028093f
C1660 VTAIL.n765 VSUBS 0.012585f
C1661 VTAIL.n766 VSUBS 0.011886f
C1662 VTAIL.n767 VSUBS 0.022119f
C1663 VTAIL.n768 VSUBS 0.022119f
C1664 VTAIL.n769 VSUBS 0.011886f
C1665 VTAIL.n770 VSUBS 0.012585f
C1666 VTAIL.n771 VSUBS 0.028093f
C1667 VTAIL.n772 VSUBS 0.028093f
C1668 VTAIL.n773 VSUBS 0.012585f
C1669 VTAIL.n774 VSUBS 0.011886f
C1670 VTAIL.n775 VSUBS 0.022119f
C1671 VTAIL.n776 VSUBS 0.022119f
C1672 VTAIL.n777 VSUBS 0.011886f
C1673 VTAIL.n778 VSUBS 0.011886f
C1674 VTAIL.n779 VSUBS 0.012585f
C1675 VTAIL.n780 VSUBS 0.028093f
C1676 VTAIL.n781 VSUBS 0.028093f
C1677 VTAIL.n782 VSUBS 0.028093f
C1678 VTAIL.n783 VSUBS 0.012235f
C1679 VTAIL.n784 VSUBS 0.011886f
C1680 VTAIL.n785 VSUBS 0.022119f
C1681 VTAIL.n786 VSUBS 0.022119f
C1682 VTAIL.n787 VSUBS 0.011886f
C1683 VTAIL.n788 VSUBS 0.012585f
C1684 VTAIL.n789 VSUBS 0.028093f
C1685 VTAIL.n790 VSUBS 0.028093f
C1686 VTAIL.n791 VSUBS 0.012585f
C1687 VTAIL.n792 VSUBS 0.011886f
C1688 VTAIL.n793 VSUBS 0.022119f
C1689 VTAIL.n794 VSUBS 0.022119f
C1690 VTAIL.n795 VSUBS 0.011886f
C1691 VTAIL.n796 VSUBS 0.012585f
C1692 VTAIL.n797 VSUBS 0.028093f
C1693 VTAIL.n798 VSUBS 0.028093f
C1694 VTAIL.n799 VSUBS 0.012585f
C1695 VTAIL.n800 VSUBS 0.011886f
C1696 VTAIL.n801 VSUBS 0.022119f
C1697 VTAIL.n802 VSUBS 0.022119f
C1698 VTAIL.n803 VSUBS 0.011886f
C1699 VTAIL.n804 VSUBS 0.012585f
C1700 VTAIL.n805 VSUBS 0.028093f
C1701 VTAIL.n806 VSUBS 0.028093f
C1702 VTAIL.n807 VSUBS 0.012585f
C1703 VTAIL.n808 VSUBS 0.011886f
C1704 VTAIL.n809 VSUBS 0.022119f
C1705 VTAIL.n810 VSUBS 0.022119f
C1706 VTAIL.n811 VSUBS 0.011886f
C1707 VTAIL.n812 VSUBS 0.012585f
C1708 VTAIL.n813 VSUBS 0.028093f
C1709 VTAIL.n814 VSUBS 0.028093f
C1710 VTAIL.n815 VSUBS 0.012585f
C1711 VTAIL.n816 VSUBS 0.011886f
C1712 VTAIL.n817 VSUBS 0.022119f
C1713 VTAIL.n818 VSUBS 0.022119f
C1714 VTAIL.n819 VSUBS 0.011886f
C1715 VTAIL.n820 VSUBS 0.012585f
C1716 VTAIL.n821 VSUBS 0.028093f
C1717 VTAIL.n822 VSUBS 0.028093f
C1718 VTAIL.n823 VSUBS 0.012585f
C1719 VTAIL.n824 VSUBS 0.011886f
C1720 VTAIL.n825 VSUBS 0.022119f
C1721 VTAIL.n826 VSUBS 0.057774f
C1722 VTAIL.n827 VSUBS 0.011886f
C1723 VTAIL.n828 VSUBS 0.012585f
C1724 VTAIL.n829 VSUBS 0.064502f
C1725 VTAIL.n830 VSUBS 0.042912f
C1726 VTAIL.n831 VSUBS 1.75142f
C1727 VDD2.t2 VSUBS 0.394052f
C1728 VDD2.t1 VSUBS 0.394052f
C1729 VDD2.n0 VSUBS 4.26998f
C1730 VDD2.t3 VSUBS 0.394052f
C1731 VDD2.t0 VSUBS 0.394052f
C1732 VDD2.n1 VSUBS 3.31867f
C1733 VDD2.n2 VSUBS 5.00863f
C1734 VN.t3 VSUBS 4.2495f
C1735 VN.t0 VSUBS 4.2561f
C1736 VN.n0 VSUBS 2.75969f
C1737 VN.t2 VSUBS 4.2495f
C1738 VN.t1 VSUBS 4.2561f
C1739 VN.n1 VSUBS 4.60332f
.ends

