* NGSPICE file created from diff_pair_sample_0876.ext - technology: sky130A

.subckt diff_pair_sample_0876 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t5 VN.t0 VTAIL.t10 w_n2674_n4626# sky130_fd_pr__pfet_01v8 ad=7.1331 pd=37.36 as=3.01785 ps=18.62 w=18.29 l=1.8
X1 VDD1.t5 VP.t0 VTAIL.t2 w_n2674_n4626# sky130_fd_pr__pfet_01v8 ad=7.1331 pd=37.36 as=3.01785 ps=18.62 w=18.29 l=1.8
X2 VDD2.t4 VN.t1 VTAIL.t9 w_n2674_n4626# sky130_fd_pr__pfet_01v8 ad=7.1331 pd=37.36 as=3.01785 ps=18.62 w=18.29 l=1.8
X3 B.t11 B.t9 B.t10 w_n2674_n4626# sky130_fd_pr__pfet_01v8 ad=7.1331 pd=37.36 as=0 ps=0 w=18.29 l=1.8
X4 VDD1.t4 VP.t1 VTAIL.t3 w_n2674_n4626# sky130_fd_pr__pfet_01v8 ad=3.01785 pd=18.62 as=7.1331 ps=37.36 w=18.29 l=1.8
X5 B.t8 B.t6 B.t7 w_n2674_n4626# sky130_fd_pr__pfet_01v8 ad=7.1331 pd=37.36 as=0 ps=0 w=18.29 l=1.8
X6 VDD2.t3 VN.t2 VTAIL.t8 w_n2674_n4626# sky130_fd_pr__pfet_01v8 ad=3.01785 pd=18.62 as=7.1331 ps=37.36 w=18.29 l=1.8
X7 VTAIL.t0 VP.t2 VDD1.t3 w_n2674_n4626# sky130_fd_pr__pfet_01v8 ad=3.01785 pd=18.62 as=3.01785 ps=18.62 w=18.29 l=1.8
X8 VTAIL.t11 VN.t3 VDD2.t2 w_n2674_n4626# sky130_fd_pr__pfet_01v8 ad=3.01785 pd=18.62 as=3.01785 ps=18.62 w=18.29 l=1.8
X9 B.t5 B.t3 B.t4 w_n2674_n4626# sky130_fd_pr__pfet_01v8 ad=7.1331 pd=37.36 as=0 ps=0 w=18.29 l=1.8
X10 VDD2.t1 VN.t4 VTAIL.t6 w_n2674_n4626# sky130_fd_pr__pfet_01v8 ad=3.01785 pd=18.62 as=7.1331 ps=37.36 w=18.29 l=1.8
X11 VTAIL.t1 VP.t3 VDD1.t2 w_n2674_n4626# sky130_fd_pr__pfet_01v8 ad=3.01785 pd=18.62 as=3.01785 ps=18.62 w=18.29 l=1.8
X12 VDD1.t1 VP.t4 VTAIL.t4 w_n2674_n4626# sky130_fd_pr__pfet_01v8 ad=3.01785 pd=18.62 as=7.1331 ps=37.36 w=18.29 l=1.8
X13 VDD1.t0 VP.t5 VTAIL.t5 w_n2674_n4626# sky130_fd_pr__pfet_01v8 ad=7.1331 pd=37.36 as=3.01785 ps=18.62 w=18.29 l=1.8
X14 VTAIL.t7 VN.t5 VDD2.t0 w_n2674_n4626# sky130_fd_pr__pfet_01v8 ad=3.01785 pd=18.62 as=3.01785 ps=18.62 w=18.29 l=1.8
X15 B.t2 B.t0 B.t1 w_n2674_n4626# sky130_fd_pr__pfet_01v8 ad=7.1331 pd=37.36 as=0 ps=0 w=18.29 l=1.8
R0 VN.n2 VN.t1 281.091
R1 VN.n14 VN.t2 281.091
R2 VN.n3 VN.t3 244.883
R3 VN.n10 VN.t4 244.883
R4 VN.n15 VN.t5 244.883
R5 VN.n22 VN.t0 244.883
R6 VN.n11 VN.n10 179.406
R7 VN.n23 VN.n22 179.406
R8 VN.n21 VN.n12 161.3
R9 VN.n20 VN.n19 161.3
R10 VN.n18 VN.n13 161.3
R11 VN.n17 VN.n16 161.3
R12 VN.n9 VN.n0 161.3
R13 VN.n8 VN.n7 161.3
R14 VN.n6 VN.n1 161.3
R15 VN.n5 VN.n4 161.3
R16 VN VN.n23 50.6274
R17 VN.n8 VN.n1 46.8066
R18 VN.n20 VN.n13 46.8066
R19 VN.n15 VN.n14 44.4618
R20 VN.n3 VN.n2 44.4618
R21 VN.n4 VN.n1 34.1802
R22 VN.n16 VN.n13 34.1802
R23 VN.n4 VN.n3 24.4675
R24 VN.n9 VN.n8 24.4675
R25 VN.n16 VN.n15 24.4675
R26 VN.n21 VN.n20 24.4675
R27 VN.n17 VN.n14 12.1055
R28 VN.n5 VN.n2 12.1055
R29 VN.n10 VN.n9 6.36192
R30 VN.n22 VN.n21 6.36192
R31 VN.n23 VN.n12 0.189894
R32 VN.n19 VN.n12 0.189894
R33 VN.n19 VN.n18 0.189894
R34 VN.n18 VN.n17 0.189894
R35 VN.n6 VN.n5 0.189894
R36 VN.n7 VN.n6 0.189894
R37 VN.n7 VN.n0 0.189894
R38 VN.n11 VN.n0 0.189894
R39 VN VN.n11 0.0516364
R40 VTAIL.n410 VTAIL.n314 756.745
R41 VTAIL.n98 VTAIL.n2 756.745
R42 VTAIL.n308 VTAIL.n212 756.745
R43 VTAIL.n204 VTAIL.n108 756.745
R44 VTAIL.n346 VTAIL.n345 585
R45 VTAIL.n351 VTAIL.n350 585
R46 VTAIL.n353 VTAIL.n352 585
R47 VTAIL.n342 VTAIL.n341 585
R48 VTAIL.n359 VTAIL.n358 585
R49 VTAIL.n361 VTAIL.n360 585
R50 VTAIL.n338 VTAIL.n337 585
R51 VTAIL.n367 VTAIL.n366 585
R52 VTAIL.n369 VTAIL.n368 585
R53 VTAIL.n334 VTAIL.n333 585
R54 VTAIL.n375 VTAIL.n374 585
R55 VTAIL.n377 VTAIL.n376 585
R56 VTAIL.n330 VTAIL.n329 585
R57 VTAIL.n383 VTAIL.n382 585
R58 VTAIL.n385 VTAIL.n384 585
R59 VTAIL.n326 VTAIL.n325 585
R60 VTAIL.n392 VTAIL.n391 585
R61 VTAIL.n393 VTAIL.n324 585
R62 VTAIL.n395 VTAIL.n394 585
R63 VTAIL.n322 VTAIL.n321 585
R64 VTAIL.n401 VTAIL.n400 585
R65 VTAIL.n403 VTAIL.n402 585
R66 VTAIL.n318 VTAIL.n317 585
R67 VTAIL.n409 VTAIL.n408 585
R68 VTAIL.n411 VTAIL.n410 585
R69 VTAIL.n34 VTAIL.n33 585
R70 VTAIL.n39 VTAIL.n38 585
R71 VTAIL.n41 VTAIL.n40 585
R72 VTAIL.n30 VTAIL.n29 585
R73 VTAIL.n47 VTAIL.n46 585
R74 VTAIL.n49 VTAIL.n48 585
R75 VTAIL.n26 VTAIL.n25 585
R76 VTAIL.n55 VTAIL.n54 585
R77 VTAIL.n57 VTAIL.n56 585
R78 VTAIL.n22 VTAIL.n21 585
R79 VTAIL.n63 VTAIL.n62 585
R80 VTAIL.n65 VTAIL.n64 585
R81 VTAIL.n18 VTAIL.n17 585
R82 VTAIL.n71 VTAIL.n70 585
R83 VTAIL.n73 VTAIL.n72 585
R84 VTAIL.n14 VTAIL.n13 585
R85 VTAIL.n80 VTAIL.n79 585
R86 VTAIL.n81 VTAIL.n12 585
R87 VTAIL.n83 VTAIL.n82 585
R88 VTAIL.n10 VTAIL.n9 585
R89 VTAIL.n89 VTAIL.n88 585
R90 VTAIL.n91 VTAIL.n90 585
R91 VTAIL.n6 VTAIL.n5 585
R92 VTAIL.n97 VTAIL.n96 585
R93 VTAIL.n99 VTAIL.n98 585
R94 VTAIL.n309 VTAIL.n308 585
R95 VTAIL.n307 VTAIL.n306 585
R96 VTAIL.n216 VTAIL.n215 585
R97 VTAIL.n301 VTAIL.n300 585
R98 VTAIL.n299 VTAIL.n298 585
R99 VTAIL.n220 VTAIL.n219 585
R100 VTAIL.n293 VTAIL.n292 585
R101 VTAIL.n291 VTAIL.n222 585
R102 VTAIL.n290 VTAIL.n289 585
R103 VTAIL.n225 VTAIL.n223 585
R104 VTAIL.n284 VTAIL.n283 585
R105 VTAIL.n282 VTAIL.n281 585
R106 VTAIL.n229 VTAIL.n228 585
R107 VTAIL.n276 VTAIL.n275 585
R108 VTAIL.n274 VTAIL.n273 585
R109 VTAIL.n233 VTAIL.n232 585
R110 VTAIL.n268 VTAIL.n267 585
R111 VTAIL.n266 VTAIL.n265 585
R112 VTAIL.n237 VTAIL.n236 585
R113 VTAIL.n260 VTAIL.n259 585
R114 VTAIL.n258 VTAIL.n257 585
R115 VTAIL.n241 VTAIL.n240 585
R116 VTAIL.n252 VTAIL.n251 585
R117 VTAIL.n250 VTAIL.n249 585
R118 VTAIL.n245 VTAIL.n244 585
R119 VTAIL.n205 VTAIL.n204 585
R120 VTAIL.n203 VTAIL.n202 585
R121 VTAIL.n112 VTAIL.n111 585
R122 VTAIL.n197 VTAIL.n196 585
R123 VTAIL.n195 VTAIL.n194 585
R124 VTAIL.n116 VTAIL.n115 585
R125 VTAIL.n189 VTAIL.n188 585
R126 VTAIL.n187 VTAIL.n118 585
R127 VTAIL.n186 VTAIL.n185 585
R128 VTAIL.n121 VTAIL.n119 585
R129 VTAIL.n180 VTAIL.n179 585
R130 VTAIL.n178 VTAIL.n177 585
R131 VTAIL.n125 VTAIL.n124 585
R132 VTAIL.n172 VTAIL.n171 585
R133 VTAIL.n170 VTAIL.n169 585
R134 VTAIL.n129 VTAIL.n128 585
R135 VTAIL.n164 VTAIL.n163 585
R136 VTAIL.n162 VTAIL.n161 585
R137 VTAIL.n133 VTAIL.n132 585
R138 VTAIL.n156 VTAIL.n155 585
R139 VTAIL.n154 VTAIL.n153 585
R140 VTAIL.n137 VTAIL.n136 585
R141 VTAIL.n148 VTAIL.n147 585
R142 VTAIL.n146 VTAIL.n145 585
R143 VTAIL.n141 VTAIL.n140 585
R144 VTAIL.n347 VTAIL.t6 327.466
R145 VTAIL.n35 VTAIL.t3 327.466
R146 VTAIL.n246 VTAIL.t4 327.466
R147 VTAIL.n142 VTAIL.t8 327.466
R148 VTAIL.n351 VTAIL.n345 171.744
R149 VTAIL.n352 VTAIL.n351 171.744
R150 VTAIL.n352 VTAIL.n341 171.744
R151 VTAIL.n359 VTAIL.n341 171.744
R152 VTAIL.n360 VTAIL.n359 171.744
R153 VTAIL.n360 VTAIL.n337 171.744
R154 VTAIL.n367 VTAIL.n337 171.744
R155 VTAIL.n368 VTAIL.n367 171.744
R156 VTAIL.n368 VTAIL.n333 171.744
R157 VTAIL.n375 VTAIL.n333 171.744
R158 VTAIL.n376 VTAIL.n375 171.744
R159 VTAIL.n376 VTAIL.n329 171.744
R160 VTAIL.n383 VTAIL.n329 171.744
R161 VTAIL.n384 VTAIL.n383 171.744
R162 VTAIL.n384 VTAIL.n325 171.744
R163 VTAIL.n392 VTAIL.n325 171.744
R164 VTAIL.n393 VTAIL.n392 171.744
R165 VTAIL.n394 VTAIL.n393 171.744
R166 VTAIL.n394 VTAIL.n321 171.744
R167 VTAIL.n401 VTAIL.n321 171.744
R168 VTAIL.n402 VTAIL.n401 171.744
R169 VTAIL.n402 VTAIL.n317 171.744
R170 VTAIL.n409 VTAIL.n317 171.744
R171 VTAIL.n410 VTAIL.n409 171.744
R172 VTAIL.n39 VTAIL.n33 171.744
R173 VTAIL.n40 VTAIL.n39 171.744
R174 VTAIL.n40 VTAIL.n29 171.744
R175 VTAIL.n47 VTAIL.n29 171.744
R176 VTAIL.n48 VTAIL.n47 171.744
R177 VTAIL.n48 VTAIL.n25 171.744
R178 VTAIL.n55 VTAIL.n25 171.744
R179 VTAIL.n56 VTAIL.n55 171.744
R180 VTAIL.n56 VTAIL.n21 171.744
R181 VTAIL.n63 VTAIL.n21 171.744
R182 VTAIL.n64 VTAIL.n63 171.744
R183 VTAIL.n64 VTAIL.n17 171.744
R184 VTAIL.n71 VTAIL.n17 171.744
R185 VTAIL.n72 VTAIL.n71 171.744
R186 VTAIL.n72 VTAIL.n13 171.744
R187 VTAIL.n80 VTAIL.n13 171.744
R188 VTAIL.n81 VTAIL.n80 171.744
R189 VTAIL.n82 VTAIL.n81 171.744
R190 VTAIL.n82 VTAIL.n9 171.744
R191 VTAIL.n89 VTAIL.n9 171.744
R192 VTAIL.n90 VTAIL.n89 171.744
R193 VTAIL.n90 VTAIL.n5 171.744
R194 VTAIL.n97 VTAIL.n5 171.744
R195 VTAIL.n98 VTAIL.n97 171.744
R196 VTAIL.n308 VTAIL.n307 171.744
R197 VTAIL.n307 VTAIL.n215 171.744
R198 VTAIL.n300 VTAIL.n215 171.744
R199 VTAIL.n300 VTAIL.n299 171.744
R200 VTAIL.n299 VTAIL.n219 171.744
R201 VTAIL.n292 VTAIL.n219 171.744
R202 VTAIL.n292 VTAIL.n291 171.744
R203 VTAIL.n291 VTAIL.n290 171.744
R204 VTAIL.n290 VTAIL.n223 171.744
R205 VTAIL.n283 VTAIL.n223 171.744
R206 VTAIL.n283 VTAIL.n282 171.744
R207 VTAIL.n282 VTAIL.n228 171.744
R208 VTAIL.n275 VTAIL.n228 171.744
R209 VTAIL.n275 VTAIL.n274 171.744
R210 VTAIL.n274 VTAIL.n232 171.744
R211 VTAIL.n267 VTAIL.n232 171.744
R212 VTAIL.n267 VTAIL.n266 171.744
R213 VTAIL.n266 VTAIL.n236 171.744
R214 VTAIL.n259 VTAIL.n236 171.744
R215 VTAIL.n259 VTAIL.n258 171.744
R216 VTAIL.n258 VTAIL.n240 171.744
R217 VTAIL.n251 VTAIL.n240 171.744
R218 VTAIL.n251 VTAIL.n250 171.744
R219 VTAIL.n250 VTAIL.n244 171.744
R220 VTAIL.n204 VTAIL.n203 171.744
R221 VTAIL.n203 VTAIL.n111 171.744
R222 VTAIL.n196 VTAIL.n111 171.744
R223 VTAIL.n196 VTAIL.n195 171.744
R224 VTAIL.n195 VTAIL.n115 171.744
R225 VTAIL.n188 VTAIL.n115 171.744
R226 VTAIL.n188 VTAIL.n187 171.744
R227 VTAIL.n187 VTAIL.n186 171.744
R228 VTAIL.n186 VTAIL.n119 171.744
R229 VTAIL.n179 VTAIL.n119 171.744
R230 VTAIL.n179 VTAIL.n178 171.744
R231 VTAIL.n178 VTAIL.n124 171.744
R232 VTAIL.n171 VTAIL.n124 171.744
R233 VTAIL.n171 VTAIL.n170 171.744
R234 VTAIL.n170 VTAIL.n128 171.744
R235 VTAIL.n163 VTAIL.n128 171.744
R236 VTAIL.n163 VTAIL.n162 171.744
R237 VTAIL.n162 VTAIL.n132 171.744
R238 VTAIL.n155 VTAIL.n132 171.744
R239 VTAIL.n155 VTAIL.n154 171.744
R240 VTAIL.n154 VTAIL.n136 171.744
R241 VTAIL.n147 VTAIL.n136 171.744
R242 VTAIL.n147 VTAIL.n146 171.744
R243 VTAIL.n146 VTAIL.n140 171.744
R244 VTAIL.t6 VTAIL.n345 85.8723
R245 VTAIL.t3 VTAIL.n33 85.8723
R246 VTAIL.t4 VTAIL.n244 85.8723
R247 VTAIL.t8 VTAIL.n140 85.8723
R248 VTAIL.n211 VTAIL.n210 52.9788
R249 VTAIL.n107 VTAIL.n106 52.9788
R250 VTAIL.n1 VTAIL.n0 52.9786
R251 VTAIL.n105 VTAIL.n104 52.9786
R252 VTAIL.n415 VTAIL.n414 33.155
R253 VTAIL.n103 VTAIL.n102 33.155
R254 VTAIL.n313 VTAIL.n312 33.155
R255 VTAIL.n209 VTAIL.n208 33.155
R256 VTAIL.n107 VTAIL.n105 31.8065
R257 VTAIL.n415 VTAIL.n313 29.9703
R258 VTAIL.n347 VTAIL.n346 16.3895
R259 VTAIL.n35 VTAIL.n34 16.3895
R260 VTAIL.n246 VTAIL.n245 16.3895
R261 VTAIL.n142 VTAIL.n141 16.3895
R262 VTAIL.n395 VTAIL.n324 13.1884
R263 VTAIL.n83 VTAIL.n12 13.1884
R264 VTAIL.n293 VTAIL.n222 13.1884
R265 VTAIL.n189 VTAIL.n118 13.1884
R266 VTAIL.n350 VTAIL.n349 12.8005
R267 VTAIL.n391 VTAIL.n390 12.8005
R268 VTAIL.n396 VTAIL.n322 12.8005
R269 VTAIL.n38 VTAIL.n37 12.8005
R270 VTAIL.n79 VTAIL.n78 12.8005
R271 VTAIL.n84 VTAIL.n10 12.8005
R272 VTAIL.n294 VTAIL.n220 12.8005
R273 VTAIL.n289 VTAIL.n224 12.8005
R274 VTAIL.n249 VTAIL.n248 12.8005
R275 VTAIL.n190 VTAIL.n116 12.8005
R276 VTAIL.n185 VTAIL.n120 12.8005
R277 VTAIL.n145 VTAIL.n144 12.8005
R278 VTAIL.n353 VTAIL.n344 12.0247
R279 VTAIL.n389 VTAIL.n326 12.0247
R280 VTAIL.n400 VTAIL.n399 12.0247
R281 VTAIL.n41 VTAIL.n32 12.0247
R282 VTAIL.n77 VTAIL.n14 12.0247
R283 VTAIL.n88 VTAIL.n87 12.0247
R284 VTAIL.n298 VTAIL.n297 12.0247
R285 VTAIL.n288 VTAIL.n225 12.0247
R286 VTAIL.n252 VTAIL.n243 12.0247
R287 VTAIL.n194 VTAIL.n193 12.0247
R288 VTAIL.n184 VTAIL.n121 12.0247
R289 VTAIL.n148 VTAIL.n139 12.0247
R290 VTAIL.n354 VTAIL.n342 11.249
R291 VTAIL.n386 VTAIL.n385 11.249
R292 VTAIL.n403 VTAIL.n320 11.249
R293 VTAIL.n42 VTAIL.n30 11.249
R294 VTAIL.n74 VTAIL.n73 11.249
R295 VTAIL.n91 VTAIL.n8 11.249
R296 VTAIL.n301 VTAIL.n218 11.249
R297 VTAIL.n285 VTAIL.n284 11.249
R298 VTAIL.n253 VTAIL.n241 11.249
R299 VTAIL.n197 VTAIL.n114 11.249
R300 VTAIL.n181 VTAIL.n180 11.249
R301 VTAIL.n149 VTAIL.n137 11.249
R302 VTAIL.n358 VTAIL.n357 10.4732
R303 VTAIL.n382 VTAIL.n328 10.4732
R304 VTAIL.n404 VTAIL.n318 10.4732
R305 VTAIL.n46 VTAIL.n45 10.4732
R306 VTAIL.n70 VTAIL.n16 10.4732
R307 VTAIL.n92 VTAIL.n6 10.4732
R308 VTAIL.n302 VTAIL.n216 10.4732
R309 VTAIL.n281 VTAIL.n227 10.4732
R310 VTAIL.n257 VTAIL.n256 10.4732
R311 VTAIL.n198 VTAIL.n112 10.4732
R312 VTAIL.n177 VTAIL.n123 10.4732
R313 VTAIL.n153 VTAIL.n152 10.4732
R314 VTAIL.n361 VTAIL.n340 9.69747
R315 VTAIL.n381 VTAIL.n330 9.69747
R316 VTAIL.n408 VTAIL.n407 9.69747
R317 VTAIL.n49 VTAIL.n28 9.69747
R318 VTAIL.n69 VTAIL.n18 9.69747
R319 VTAIL.n96 VTAIL.n95 9.69747
R320 VTAIL.n306 VTAIL.n305 9.69747
R321 VTAIL.n280 VTAIL.n229 9.69747
R322 VTAIL.n260 VTAIL.n239 9.69747
R323 VTAIL.n202 VTAIL.n201 9.69747
R324 VTAIL.n176 VTAIL.n125 9.69747
R325 VTAIL.n156 VTAIL.n135 9.69747
R326 VTAIL.n414 VTAIL.n413 9.45567
R327 VTAIL.n102 VTAIL.n101 9.45567
R328 VTAIL.n312 VTAIL.n311 9.45567
R329 VTAIL.n208 VTAIL.n207 9.45567
R330 VTAIL.n413 VTAIL.n412 9.3005
R331 VTAIL.n316 VTAIL.n315 9.3005
R332 VTAIL.n407 VTAIL.n406 9.3005
R333 VTAIL.n405 VTAIL.n404 9.3005
R334 VTAIL.n320 VTAIL.n319 9.3005
R335 VTAIL.n399 VTAIL.n398 9.3005
R336 VTAIL.n397 VTAIL.n396 9.3005
R337 VTAIL.n336 VTAIL.n335 9.3005
R338 VTAIL.n365 VTAIL.n364 9.3005
R339 VTAIL.n363 VTAIL.n362 9.3005
R340 VTAIL.n340 VTAIL.n339 9.3005
R341 VTAIL.n357 VTAIL.n356 9.3005
R342 VTAIL.n355 VTAIL.n354 9.3005
R343 VTAIL.n344 VTAIL.n343 9.3005
R344 VTAIL.n349 VTAIL.n348 9.3005
R345 VTAIL.n371 VTAIL.n370 9.3005
R346 VTAIL.n373 VTAIL.n372 9.3005
R347 VTAIL.n332 VTAIL.n331 9.3005
R348 VTAIL.n379 VTAIL.n378 9.3005
R349 VTAIL.n381 VTAIL.n380 9.3005
R350 VTAIL.n328 VTAIL.n327 9.3005
R351 VTAIL.n387 VTAIL.n386 9.3005
R352 VTAIL.n389 VTAIL.n388 9.3005
R353 VTAIL.n390 VTAIL.n323 9.3005
R354 VTAIL.n101 VTAIL.n100 9.3005
R355 VTAIL.n4 VTAIL.n3 9.3005
R356 VTAIL.n95 VTAIL.n94 9.3005
R357 VTAIL.n93 VTAIL.n92 9.3005
R358 VTAIL.n8 VTAIL.n7 9.3005
R359 VTAIL.n87 VTAIL.n86 9.3005
R360 VTAIL.n85 VTAIL.n84 9.3005
R361 VTAIL.n24 VTAIL.n23 9.3005
R362 VTAIL.n53 VTAIL.n52 9.3005
R363 VTAIL.n51 VTAIL.n50 9.3005
R364 VTAIL.n28 VTAIL.n27 9.3005
R365 VTAIL.n45 VTAIL.n44 9.3005
R366 VTAIL.n43 VTAIL.n42 9.3005
R367 VTAIL.n32 VTAIL.n31 9.3005
R368 VTAIL.n37 VTAIL.n36 9.3005
R369 VTAIL.n59 VTAIL.n58 9.3005
R370 VTAIL.n61 VTAIL.n60 9.3005
R371 VTAIL.n20 VTAIL.n19 9.3005
R372 VTAIL.n67 VTAIL.n66 9.3005
R373 VTAIL.n69 VTAIL.n68 9.3005
R374 VTAIL.n16 VTAIL.n15 9.3005
R375 VTAIL.n75 VTAIL.n74 9.3005
R376 VTAIL.n77 VTAIL.n76 9.3005
R377 VTAIL.n78 VTAIL.n11 9.3005
R378 VTAIL.n272 VTAIL.n271 9.3005
R379 VTAIL.n231 VTAIL.n230 9.3005
R380 VTAIL.n278 VTAIL.n277 9.3005
R381 VTAIL.n280 VTAIL.n279 9.3005
R382 VTAIL.n227 VTAIL.n226 9.3005
R383 VTAIL.n286 VTAIL.n285 9.3005
R384 VTAIL.n288 VTAIL.n287 9.3005
R385 VTAIL.n224 VTAIL.n221 9.3005
R386 VTAIL.n311 VTAIL.n310 9.3005
R387 VTAIL.n214 VTAIL.n213 9.3005
R388 VTAIL.n305 VTAIL.n304 9.3005
R389 VTAIL.n303 VTAIL.n302 9.3005
R390 VTAIL.n218 VTAIL.n217 9.3005
R391 VTAIL.n297 VTAIL.n296 9.3005
R392 VTAIL.n295 VTAIL.n294 9.3005
R393 VTAIL.n270 VTAIL.n269 9.3005
R394 VTAIL.n235 VTAIL.n234 9.3005
R395 VTAIL.n264 VTAIL.n263 9.3005
R396 VTAIL.n262 VTAIL.n261 9.3005
R397 VTAIL.n239 VTAIL.n238 9.3005
R398 VTAIL.n256 VTAIL.n255 9.3005
R399 VTAIL.n254 VTAIL.n253 9.3005
R400 VTAIL.n243 VTAIL.n242 9.3005
R401 VTAIL.n248 VTAIL.n247 9.3005
R402 VTAIL.n168 VTAIL.n167 9.3005
R403 VTAIL.n127 VTAIL.n126 9.3005
R404 VTAIL.n174 VTAIL.n173 9.3005
R405 VTAIL.n176 VTAIL.n175 9.3005
R406 VTAIL.n123 VTAIL.n122 9.3005
R407 VTAIL.n182 VTAIL.n181 9.3005
R408 VTAIL.n184 VTAIL.n183 9.3005
R409 VTAIL.n120 VTAIL.n117 9.3005
R410 VTAIL.n207 VTAIL.n206 9.3005
R411 VTAIL.n110 VTAIL.n109 9.3005
R412 VTAIL.n201 VTAIL.n200 9.3005
R413 VTAIL.n199 VTAIL.n198 9.3005
R414 VTAIL.n114 VTAIL.n113 9.3005
R415 VTAIL.n193 VTAIL.n192 9.3005
R416 VTAIL.n191 VTAIL.n190 9.3005
R417 VTAIL.n166 VTAIL.n165 9.3005
R418 VTAIL.n131 VTAIL.n130 9.3005
R419 VTAIL.n160 VTAIL.n159 9.3005
R420 VTAIL.n158 VTAIL.n157 9.3005
R421 VTAIL.n135 VTAIL.n134 9.3005
R422 VTAIL.n152 VTAIL.n151 9.3005
R423 VTAIL.n150 VTAIL.n149 9.3005
R424 VTAIL.n139 VTAIL.n138 9.3005
R425 VTAIL.n144 VTAIL.n143 9.3005
R426 VTAIL.n362 VTAIL.n338 8.92171
R427 VTAIL.n378 VTAIL.n377 8.92171
R428 VTAIL.n411 VTAIL.n316 8.92171
R429 VTAIL.n50 VTAIL.n26 8.92171
R430 VTAIL.n66 VTAIL.n65 8.92171
R431 VTAIL.n99 VTAIL.n4 8.92171
R432 VTAIL.n309 VTAIL.n214 8.92171
R433 VTAIL.n277 VTAIL.n276 8.92171
R434 VTAIL.n261 VTAIL.n237 8.92171
R435 VTAIL.n205 VTAIL.n110 8.92171
R436 VTAIL.n173 VTAIL.n172 8.92171
R437 VTAIL.n157 VTAIL.n133 8.92171
R438 VTAIL.n366 VTAIL.n365 8.14595
R439 VTAIL.n374 VTAIL.n332 8.14595
R440 VTAIL.n412 VTAIL.n314 8.14595
R441 VTAIL.n54 VTAIL.n53 8.14595
R442 VTAIL.n62 VTAIL.n20 8.14595
R443 VTAIL.n100 VTAIL.n2 8.14595
R444 VTAIL.n310 VTAIL.n212 8.14595
R445 VTAIL.n273 VTAIL.n231 8.14595
R446 VTAIL.n265 VTAIL.n264 8.14595
R447 VTAIL.n206 VTAIL.n108 8.14595
R448 VTAIL.n169 VTAIL.n127 8.14595
R449 VTAIL.n161 VTAIL.n160 8.14595
R450 VTAIL.n369 VTAIL.n336 7.3702
R451 VTAIL.n373 VTAIL.n334 7.3702
R452 VTAIL.n57 VTAIL.n24 7.3702
R453 VTAIL.n61 VTAIL.n22 7.3702
R454 VTAIL.n272 VTAIL.n233 7.3702
R455 VTAIL.n268 VTAIL.n235 7.3702
R456 VTAIL.n168 VTAIL.n129 7.3702
R457 VTAIL.n164 VTAIL.n131 7.3702
R458 VTAIL.n370 VTAIL.n369 6.59444
R459 VTAIL.n370 VTAIL.n334 6.59444
R460 VTAIL.n58 VTAIL.n57 6.59444
R461 VTAIL.n58 VTAIL.n22 6.59444
R462 VTAIL.n269 VTAIL.n233 6.59444
R463 VTAIL.n269 VTAIL.n268 6.59444
R464 VTAIL.n165 VTAIL.n129 6.59444
R465 VTAIL.n165 VTAIL.n164 6.59444
R466 VTAIL.n366 VTAIL.n336 5.81868
R467 VTAIL.n374 VTAIL.n373 5.81868
R468 VTAIL.n414 VTAIL.n314 5.81868
R469 VTAIL.n54 VTAIL.n24 5.81868
R470 VTAIL.n62 VTAIL.n61 5.81868
R471 VTAIL.n102 VTAIL.n2 5.81868
R472 VTAIL.n312 VTAIL.n212 5.81868
R473 VTAIL.n273 VTAIL.n272 5.81868
R474 VTAIL.n265 VTAIL.n235 5.81868
R475 VTAIL.n208 VTAIL.n108 5.81868
R476 VTAIL.n169 VTAIL.n168 5.81868
R477 VTAIL.n161 VTAIL.n131 5.81868
R478 VTAIL.n365 VTAIL.n338 5.04292
R479 VTAIL.n377 VTAIL.n332 5.04292
R480 VTAIL.n412 VTAIL.n411 5.04292
R481 VTAIL.n53 VTAIL.n26 5.04292
R482 VTAIL.n65 VTAIL.n20 5.04292
R483 VTAIL.n100 VTAIL.n99 5.04292
R484 VTAIL.n310 VTAIL.n309 5.04292
R485 VTAIL.n276 VTAIL.n231 5.04292
R486 VTAIL.n264 VTAIL.n237 5.04292
R487 VTAIL.n206 VTAIL.n205 5.04292
R488 VTAIL.n172 VTAIL.n127 5.04292
R489 VTAIL.n160 VTAIL.n133 5.04292
R490 VTAIL.n362 VTAIL.n361 4.26717
R491 VTAIL.n378 VTAIL.n330 4.26717
R492 VTAIL.n408 VTAIL.n316 4.26717
R493 VTAIL.n50 VTAIL.n49 4.26717
R494 VTAIL.n66 VTAIL.n18 4.26717
R495 VTAIL.n96 VTAIL.n4 4.26717
R496 VTAIL.n306 VTAIL.n214 4.26717
R497 VTAIL.n277 VTAIL.n229 4.26717
R498 VTAIL.n261 VTAIL.n260 4.26717
R499 VTAIL.n202 VTAIL.n110 4.26717
R500 VTAIL.n173 VTAIL.n125 4.26717
R501 VTAIL.n157 VTAIL.n156 4.26717
R502 VTAIL.n348 VTAIL.n347 3.70982
R503 VTAIL.n36 VTAIL.n35 3.70982
R504 VTAIL.n247 VTAIL.n246 3.70982
R505 VTAIL.n143 VTAIL.n142 3.70982
R506 VTAIL.n358 VTAIL.n340 3.49141
R507 VTAIL.n382 VTAIL.n381 3.49141
R508 VTAIL.n407 VTAIL.n318 3.49141
R509 VTAIL.n46 VTAIL.n28 3.49141
R510 VTAIL.n70 VTAIL.n69 3.49141
R511 VTAIL.n95 VTAIL.n6 3.49141
R512 VTAIL.n305 VTAIL.n216 3.49141
R513 VTAIL.n281 VTAIL.n280 3.49141
R514 VTAIL.n257 VTAIL.n239 3.49141
R515 VTAIL.n201 VTAIL.n112 3.49141
R516 VTAIL.n177 VTAIL.n176 3.49141
R517 VTAIL.n153 VTAIL.n135 3.49141
R518 VTAIL.n357 VTAIL.n342 2.71565
R519 VTAIL.n385 VTAIL.n328 2.71565
R520 VTAIL.n404 VTAIL.n403 2.71565
R521 VTAIL.n45 VTAIL.n30 2.71565
R522 VTAIL.n73 VTAIL.n16 2.71565
R523 VTAIL.n92 VTAIL.n91 2.71565
R524 VTAIL.n302 VTAIL.n301 2.71565
R525 VTAIL.n284 VTAIL.n227 2.71565
R526 VTAIL.n256 VTAIL.n241 2.71565
R527 VTAIL.n198 VTAIL.n197 2.71565
R528 VTAIL.n180 VTAIL.n123 2.71565
R529 VTAIL.n152 VTAIL.n137 2.71565
R530 VTAIL.n354 VTAIL.n353 1.93989
R531 VTAIL.n386 VTAIL.n326 1.93989
R532 VTAIL.n400 VTAIL.n320 1.93989
R533 VTAIL.n42 VTAIL.n41 1.93989
R534 VTAIL.n74 VTAIL.n14 1.93989
R535 VTAIL.n88 VTAIL.n8 1.93989
R536 VTAIL.n298 VTAIL.n218 1.93989
R537 VTAIL.n285 VTAIL.n225 1.93989
R538 VTAIL.n253 VTAIL.n252 1.93989
R539 VTAIL.n194 VTAIL.n114 1.93989
R540 VTAIL.n181 VTAIL.n121 1.93989
R541 VTAIL.n149 VTAIL.n148 1.93989
R542 VTAIL.n209 VTAIL.n107 1.83671
R543 VTAIL.n313 VTAIL.n211 1.83671
R544 VTAIL.n105 VTAIL.n103 1.83671
R545 VTAIL.n0 VTAIL.t9 1.7777
R546 VTAIL.n0 VTAIL.t11 1.7777
R547 VTAIL.n104 VTAIL.t5 1.7777
R548 VTAIL.n104 VTAIL.t1 1.7777
R549 VTAIL.n210 VTAIL.t2 1.7777
R550 VTAIL.n210 VTAIL.t0 1.7777
R551 VTAIL.n106 VTAIL.t10 1.7777
R552 VTAIL.n106 VTAIL.t7 1.7777
R553 VTAIL.n211 VTAIL.n209 1.38843
R554 VTAIL.n103 VTAIL.n1 1.38843
R555 VTAIL VTAIL.n415 1.31947
R556 VTAIL.n350 VTAIL.n344 1.16414
R557 VTAIL.n391 VTAIL.n389 1.16414
R558 VTAIL.n399 VTAIL.n322 1.16414
R559 VTAIL.n38 VTAIL.n32 1.16414
R560 VTAIL.n79 VTAIL.n77 1.16414
R561 VTAIL.n87 VTAIL.n10 1.16414
R562 VTAIL.n297 VTAIL.n220 1.16414
R563 VTAIL.n289 VTAIL.n288 1.16414
R564 VTAIL.n249 VTAIL.n243 1.16414
R565 VTAIL.n193 VTAIL.n116 1.16414
R566 VTAIL.n185 VTAIL.n184 1.16414
R567 VTAIL.n145 VTAIL.n139 1.16414
R568 VTAIL VTAIL.n1 0.517741
R569 VTAIL.n349 VTAIL.n346 0.388379
R570 VTAIL.n390 VTAIL.n324 0.388379
R571 VTAIL.n396 VTAIL.n395 0.388379
R572 VTAIL.n37 VTAIL.n34 0.388379
R573 VTAIL.n78 VTAIL.n12 0.388379
R574 VTAIL.n84 VTAIL.n83 0.388379
R575 VTAIL.n294 VTAIL.n293 0.388379
R576 VTAIL.n224 VTAIL.n222 0.388379
R577 VTAIL.n248 VTAIL.n245 0.388379
R578 VTAIL.n190 VTAIL.n189 0.388379
R579 VTAIL.n120 VTAIL.n118 0.388379
R580 VTAIL.n144 VTAIL.n141 0.388379
R581 VTAIL.n348 VTAIL.n343 0.155672
R582 VTAIL.n355 VTAIL.n343 0.155672
R583 VTAIL.n356 VTAIL.n355 0.155672
R584 VTAIL.n356 VTAIL.n339 0.155672
R585 VTAIL.n363 VTAIL.n339 0.155672
R586 VTAIL.n364 VTAIL.n363 0.155672
R587 VTAIL.n364 VTAIL.n335 0.155672
R588 VTAIL.n371 VTAIL.n335 0.155672
R589 VTAIL.n372 VTAIL.n371 0.155672
R590 VTAIL.n372 VTAIL.n331 0.155672
R591 VTAIL.n379 VTAIL.n331 0.155672
R592 VTAIL.n380 VTAIL.n379 0.155672
R593 VTAIL.n380 VTAIL.n327 0.155672
R594 VTAIL.n387 VTAIL.n327 0.155672
R595 VTAIL.n388 VTAIL.n387 0.155672
R596 VTAIL.n388 VTAIL.n323 0.155672
R597 VTAIL.n397 VTAIL.n323 0.155672
R598 VTAIL.n398 VTAIL.n397 0.155672
R599 VTAIL.n398 VTAIL.n319 0.155672
R600 VTAIL.n405 VTAIL.n319 0.155672
R601 VTAIL.n406 VTAIL.n405 0.155672
R602 VTAIL.n406 VTAIL.n315 0.155672
R603 VTAIL.n413 VTAIL.n315 0.155672
R604 VTAIL.n36 VTAIL.n31 0.155672
R605 VTAIL.n43 VTAIL.n31 0.155672
R606 VTAIL.n44 VTAIL.n43 0.155672
R607 VTAIL.n44 VTAIL.n27 0.155672
R608 VTAIL.n51 VTAIL.n27 0.155672
R609 VTAIL.n52 VTAIL.n51 0.155672
R610 VTAIL.n52 VTAIL.n23 0.155672
R611 VTAIL.n59 VTAIL.n23 0.155672
R612 VTAIL.n60 VTAIL.n59 0.155672
R613 VTAIL.n60 VTAIL.n19 0.155672
R614 VTAIL.n67 VTAIL.n19 0.155672
R615 VTAIL.n68 VTAIL.n67 0.155672
R616 VTAIL.n68 VTAIL.n15 0.155672
R617 VTAIL.n75 VTAIL.n15 0.155672
R618 VTAIL.n76 VTAIL.n75 0.155672
R619 VTAIL.n76 VTAIL.n11 0.155672
R620 VTAIL.n85 VTAIL.n11 0.155672
R621 VTAIL.n86 VTAIL.n85 0.155672
R622 VTAIL.n86 VTAIL.n7 0.155672
R623 VTAIL.n93 VTAIL.n7 0.155672
R624 VTAIL.n94 VTAIL.n93 0.155672
R625 VTAIL.n94 VTAIL.n3 0.155672
R626 VTAIL.n101 VTAIL.n3 0.155672
R627 VTAIL.n311 VTAIL.n213 0.155672
R628 VTAIL.n304 VTAIL.n213 0.155672
R629 VTAIL.n304 VTAIL.n303 0.155672
R630 VTAIL.n303 VTAIL.n217 0.155672
R631 VTAIL.n296 VTAIL.n217 0.155672
R632 VTAIL.n296 VTAIL.n295 0.155672
R633 VTAIL.n295 VTAIL.n221 0.155672
R634 VTAIL.n287 VTAIL.n221 0.155672
R635 VTAIL.n287 VTAIL.n286 0.155672
R636 VTAIL.n286 VTAIL.n226 0.155672
R637 VTAIL.n279 VTAIL.n226 0.155672
R638 VTAIL.n279 VTAIL.n278 0.155672
R639 VTAIL.n278 VTAIL.n230 0.155672
R640 VTAIL.n271 VTAIL.n230 0.155672
R641 VTAIL.n271 VTAIL.n270 0.155672
R642 VTAIL.n270 VTAIL.n234 0.155672
R643 VTAIL.n263 VTAIL.n234 0.155672
R644 VTAIL.n263 VTAIL.n262 0.155672
R645 VTAIL.n262 VTAIL.n238 0.155672
R646 VTAIL.n255 VTAIL.n238 0.155672
R647 VTAIL.n255 VTAIL.n254 0.155672
R648 VTAIL.n254 VTAIL.n242 0.155672
R649 VTAIL.n247 VTAIL.n242 0.155672
R650 VTAIL.n207 VTAIL.n109 0.155672
R651 VTAIL.n200 VTAIL.n109 0.155672
R652 VTAIL.n200 VTAIL.n199 0.155672
R653 VTAIL.n199 VTAIL.n113 0.155672
R654 VTAIL.n192 VTAIL.n113 0.155672
R655 VTAIL.n192 VTAIL.n191 0.155672
R656 VTAIL.n191 VTAIL.n117 0.155672
R657 VTAIL.n183 VTAIL.n117 0.155672
R658 VTAIL.n183 VTAIL.n182 0.155672
R659 VTAIL.n182 VTAIL.n122 0.155672
R660 VTAIL.n175 VTAIL.n122 0.155672
R661 VTAIL.n175 VTAIL.n174 0.155672
R662 VTAIL.n174 VTAIL.n126 0.155672
R663 VTAIL.n167 VTAIL.n126 0.155672
R664 VTAIL.n167 VTAIL.n166 0.155672
R665 VTAIL.n166 VTAIL.n130 0.155672
R666 VTAIL.n159 VTAIL.n130 0.155672
R667 VTAIL.n159 VTAIL.n158 0.155672
R668 VTAIL.n158 VTAIL.n134 0.155672
R669 VTAIL.n151 VTAIL.n134 0.155672
R670 VTAIL.n151 VTAIL.n150 0.155672
R671 VTAIL.n150 VTAIL.n138 0.155672
R672 VTAIL.n143 VTAIL.n138 0.155672
R673 VDD2.n199 VDD2.n103 756.745
R674 VDD2.n96 VDD2.n0 756.745
R675 VDD2.n200 VDD2.n199 585
R676 VDD2.n198 VDD2.n197 585
R677 VDD2.n107 VDD2.n106 585
R678 VDD2.n192 VDD2.n191 585
R679 VDD2.n190 VDD2.n189 585
R680 VDD2.n111 VDD2.n110 585
R681 VDD2.n184 VDD2.n183 585
R682 VDD2.n182 VDD2.n113 585
R683 VDD2.n181 VDD2.n180 585
R684 VDD2.n116 VDD2.n114 585
R685 VDD2.n175 VDD2.n174 585
R686 VDD2.n173 VDD2.n172 585
R687 VDD2.n120 VDD2.n119 585
R688 VDD2.n167 VDD2.n166 585
R689 VDD2.n165 VDD2.n164 585
R690 VDD2.n124 VDD2.n123 585
R691 VDD2.n159 VDD2.n158 585
R692 VDD2.n157 VDD2.n156 585
R693 VDD2.n128 VDD2.n127 585
R694 VDD2.n151 VDD2.n150 585
R695 VDD2.n149 VDD2.n148 585
R696 VDD2.n132 VDD2.n131 585
R697 VDD2.n143 VDD2.n142 585
R698 VDD2.n141 VDD2.n140 585
R699 VDD2.n136 VDD2.n135 585
R700 VDD2.n32 VDD2.n31 585
R701 VDD2.n37 VDD2.n36 585
R702 VDD2.n39 VDD2.n38 585
R703 VDD2.n28 VDD2.n27 585
R704 VDD2.n45 VDD2.n44 585
R705 VDD2.n47 VDD2.n46 585
R706 VDD2.n24 VDD2.n23 585
R707 VDD2.n53 VDD2.n52 585
R708 VDD2.n55 VDD2.n54 585
R709 VDD2.n20 VDD2.n19 585
R710 VDD2.n61 VDD2.n60 585
R711 VDD2.n63 VDD2.n62 585
R712 VDD2.n16 VDD2.n15 585
R713 VDD2.n69 VDD2.n68 585
R714 VDD2.n71 VDD2.n70 585
R715 VDD2.n12 VDD2.n11 585
R716 VDD2.n78 VDD2.n77 585
R717 VDD2.n79 VDD2.n10 585
R718 VDD2.n81 VDD2.n80 585
R719 VDD2.n8 VDD2.n7 585
R720 VDD2.n87 VDD2.n86 585
R721 VDD2.n89 VDD2.n88 585
R722 VDD2.n4 VDD2.n3 585
R723 VDD2.n95 VDD2.n94 585
R724 VDD2.n97 VDD2.n96 585
R725 VDD2.n137 VDD2.t5 327.466
R726 VDD2.n33 VDD2.t4 327.466
R727 VDD2.n199 VDD2.n198 171.744
R728 VDD2.n198 VDD2.n106 171.744
R729 VDD2.n191 VDD2.n106 171.744
R730 VDD2.n191 VDD2.n190 171.744
R731 VDD2.n190 VDD2.n110 171.744
R732 VDD2.n183 VDD2.n110 171.744
R733 VDD2.n183 VDD2.n182 171.744
R734 VDD2.n182 VDD2.n181 171.744
R735 VDD2.n181 VDD2.n114 171.744
R736 VDD2.n174 VDD2.n114 171.744
R737 VDD2.n174 VDD2.n173 171.744
R738 VDD2.n173 VDD2.n119 171.744
R739 VDD2.n166 VDD2.n119 171.744
R740 VDD2.n166 VDD2.n165 171.744
R741 VDD2.n165 VDD2.n123 171.744
R742 VDD2.n158 VDD2.n123 171.744
R743 VDD2.n158 VDD2.n157 171.744
R744 VDD2.n157 VDD2.n127 171.744
R745 VDD2.n150 VDD2.n127 171.744
R746 VDD2.n150 VDD2.n149 171.744
R747 VDD2.n149 VDD2.n131 171.744
R748 VDD2.n142 VDD2.n131 171.744
R749 VDD2.n142 VDD2.n141 171.744
R750 VDD2.n141 VDD2.n135 171.744
R751 VDD2.n37 VDD2.n31 171.744
R752 VDD2.n38 VDD2.n37 171.744
R753 VDD2.n38 VDD2.n27 171.744
R754 VDD2.n45 VDD2.n27 171.744
R755 VDD2.n46 VDD2.n45 171.744
R756 VDD2.n46 VDD2.n23 171.744
R757 VDD2.n53 VDD2.n23 171.744
R758 VDD2.n54 VDD2.n53 171.744
R759 VDD2.n54 VDD2.n19 171.744
R760 VDD2.n61 VDD2.n19 171.744
R761 VDD2.n62 VDD2.n61 171.744
R762 VDD2.n62 VDD2.n15 171.744
R763 VDD2.n69 VDD2.n15 171.744
R764 VDD2.n70 VDD2.n69 171.744
R765 VDD2.n70 VDD2.n11 171.744
R766 VDD2.n78 VDD2.n11 171.744
R767 VDD2.n79 VDD2.n78 171.744
R768 VDD2.n80 VDD2.n79 171.744
R769 VDD2.n80 VDD2.n7 171.744
R770 VDD2.n87 VDD2.n7 171.744
R771 VDD2.n88 VDD2.n87 171.744
R772 VDD2.n88 VDD2.n3 171.744
R773 VDD2.n95 VDD2.n3 171.744
R774 VDD2.n96 VDD2.n95 171.744
R775 VDD2.t5 VDD2.n135 85.8723
R776 VDD2.t4 VDD2.n31 85.8723
R777 VDD2.n102 VDD2.n101 70.0611
R778 VDD2 VDD2.n205 70.0583
R779 VDD2.n102 VDD2.n100 51.1556
R780 VDD2.n204 VDD2.n203 49.8338
R781 VDD2.n204 VDD2.n102 45.4502
R782 VDD2.n137 VDD2.n136 16.3895
R783 VDD2.n33 VDD2.n32 16.3895
R784 VDD2.n184 VDD2.n113 13.1884
R785 VDD2.n81 VDD2.n10 13.1884
R786 VDD2.n185 VDD2.n111 12.8005
R787 VDD2.n180 VDD2.n115 12.8005
R788 VDD2.n140 VDD2.n139 12.8005
R789 VDD2.n36 VDD2.n35 12.8005
R790 VDD2.n77 VDD2.n76 12.8005
R791 VDD2.n82 VDD2.n8 12.8005
R792 VDD2.n189 VDD2.n188 12.0247
R793 VDD2.n179 VDD2.n116 12.0247
R794 VDD2.n143 VDD2.n134 12.0247
R795 VDD2.n39 VDD2.n30 12.0247
R796 VDD2.n75 VDD2.n12 12.0247
R797 VDD2.n86 VDD2.n85 12.0247
R798 VDD2.n192 VDD2.n109 11.249
R799 VDD2.n176 VDD2.n175 11.249
R800 VDD2.n144 VDD2.n132 11.249
R801 VDD2.n40 VDD2.n28 11.249
R802 VDD2.n72 VDD2.n71 11.249
R803 VDD2.n89 VDD2.n6 11.249
R804 VDD2.n193 VDD2.n107 10.4732
R805 VDD2.n172 VDD2.n118 10.4732
R806 VDD2.n148 VDD2.n147 10.4732
R807 VDD2.n44 VDD2.n43 10.4732
R808 VDD2.n68 VDD2.n14 10.4732
R809 VDD2.n90 VDD2.n4 10.4732
R810 VDD2.n197 VDD2.n196 9.69747
R811 VDD2.n171 VDD2.n120 9.69747
R812 VDD2.n151 VDD2.n130 9.69747
R813 VDD2.n47 VDD2.n26 9.69747
R814 VDD2.n67 VDD2.n16 9.69747
R815 VDD2.n94 VDD2.n93 9.69747
R816 VDD2.n203 VDD2.n202 9.45567
R817 VDD2.n100 VDD2.n99 9.45567
R818 VDD2.n163 VDD2.n162 9.3005
R819 VDD2.n122 VDD2.n121 9.3005
R820 VDD2.n169 VDD2.n168 9.3005
R821 VDD2.n171 VDD2.n170 9.3005
R822 VDD2.n118 VDD2.n117 9.3005
R823 VDD2.n177 VDD2.n176 9.3005
R824 VDD2.n179 VDD2.n178 9.3005
R825 VDD2.n115 VDD2.n112 9.3005
R826 VDD2.n202 VDD2.n201 9.3005
R827 VDD2.n105 VDD2.n104 9.3005
R828 VDD2.n196 VDD2.n195 9.3005
R829 VDD2.n194 VDD2.n193 9.3005
R830 VDD2.n109 VDD2.n108 9.3005
R831 VDD2.n188 VDD2.n187 9.3005
R832 VDD2.n186 VDD2.n185 9.3005
R833 VDD2.n161 VDD2.n160 9.3005
R834 VDD2.n126 VDD2.n125 9.3005
R835 VDD2.n155 VDD2.n154 9.3005
R836 VDD2.n153 VDD2.n152 9.3005
R837 VDD2.n130 VDD2.n129 9.3005
R838 VDD2.n147 VDD2.n146 9.3005
R839 VDD2.n145 VDD2.n144 9.3005
R840 VDD2.n134 VDD2.n133 9.3005
R841 VDD2.n139 VDD2.n138 9.3005
R842 VDD2.n99 VDD2.n98 9.3005
R843 VDD2.n2 VDD2.n1 9.3005
R844 VDD2.n93 VDD2.n92 9.3005
R845 VDD2.n91 VDD2.n90 9.3005
R846 VDD2.n6 VDD2.n5 9.3005
R847 VDD2.n85 VDD2.n84 9.3005
R848 VDD2.n83 VDD2.n82 9.3005
R849 VDD2.n22 VDD2.n21 9.3005
R850 VDD2.n51 VDD2.n50 9.3005
R851 VDD2.n49 VDD2.n48 9.3005
R852 VDD2.n26 VDD2.n25 9.3005
R853 VDD2.n43 VDD2.n42 9.3005
R854 VDD2.n41 VDD2.n40 9.3005
R855 VDD2.n30 VDD2.n29 9.3005
R856 VDD2.n35 VDD2.n34 9.3005
R857 VDD2.n57 VDD2.n56 9.3005
R858 VDD2.n59 VDD2.n58 9.3005
R859 VDD2.n18 VDD2.n17 9.3005
R860 VDD2.n65 VDD2.n64 9.3005
R861 VDD2.n67 VDD2.n66 9.3005
R862 VDD2.n14 VDD2.n13 9.3005
R863 VDD2.n73 VDD2.n72 9.3005
R864 VDD2.n75 VDD2.n74 9.3005
R865 VDD2.n76 VDD2.n9 9.3005
R866 VDD2.n200 VDD2.n105 8.92171
R867 VDD2.n168 VDD2.n167 8.92171
R868 VDD2.n152 VDD2.n128 8.92171
R869 VDD2.n48 VDD2.n24 8.92171
R870 VDD2.n64 VDD2.n63 8.92171
R871 VDD2.n97 VDD2.n2 8.92171
R872 VDD2.n201 VDD2.n103 8.14595
R873 VDD2.n164 VDD2.n122 8.14595
R874 VDD2.n156 VDD2.n155 8.14595
R875 VDD2.n52 VDD2.n51 8.14595
R876 VDD2.n60 VDD2.n18 8.14595
R877 VDD2.n98 VDD2.n0 8.14595
R878 VDD2.n163 VDD2.n124 7.3702
R879 VDD2.n159 VDD2.n126 7.3702
R880 VDD2.n55 VDD2.n22 7.3702
R881 VDD2.n59 VDD2.n20 7.3702
R882 VDD2.n160 VDD2.n124 6.59444
R883 VDD2.n160 VDD2.n159 6.59444
R884 VDD2.n56 VDD2.n55 6.59444
R885 VDD2.n56 VDD2.n20 6.59444
R886 VDD2.n203 VDD2.n103 5.81868
R887 VDD2.n164 VDD2.n163 5.81868
R888 VDD2.n156 VDD2.n126 5.81868
R889 VDD2.n52 VDD2.n22 5.81868
R890 VDD2.n60 VDD2.n59 5.81868
R891 VDD2.n100 VDD2.n0 5.81868
R892 VDD2.n201 VDD2.n200 5.04292
R893 VDD2.n167 VDD2.n122 5.04292
R894 VDD2.n155 VDD2.n128 5.04292
R895 VDD2.n51 VDD2.n24 5.04292
R896 VDD2.n63 VDD2.n18 5.04292
R897 VDD2.n98 VDD2.n97 5.04292
R898 VDD2.n197 VDD2.n105 4.26717
R899 VDD2.n168 VDD2.n120 4.26717
R900 VDD2.n152 VDD2.n151 4.26717
R901 VDD2.n48 VDD2.n47 4.26717
R902 VDD2.n64 VDD2.n16 4.26717
R903 VDD2.n94 VDD2.n2 4.26717
R904 VDD2.n138 VDD2.n137 3.70982
R905 VDD2.n34 VDD2.n33 3.70982
R906 VDD2.n196 VDD2.n107 3.49141
R907 VDD2.n172 VDD2.n171 3.49141
R908 VDD2.n148 VDD2.n130 3.49141
R909 VDD2.n44 VDD2.n26 3.49141
R910 VDD2.n68 VDD2.n67 3.49141
R911 VDD2.n93 VDD2.n4 3.49141
R912 VDD2.n193 VDD2.n192 2.71565
R913 VDD2.n175 VDD2.n118 2.71565
R914 VDD2.n147 VDD2.n132 2.71565
R915 VDD2.n43 VDD2.n28 2.71565
R916 VDD2.n71 VDD2.n14 2.71565
R917 VDD2.n90 VDD2.n89 2.71565
R918 VDD2.n189 VDD2.n109 1.93989
R919 VDD2.n176 VDD2.n116 1.93989
R920 VDD2.n144 VDD2.n143 1.93989
R921 VDD2.n40 VDD2.n39 1.93989
R922 VDD2.n72 VDD2.n12 1.93989
R923 VDD2.n86 VDD2.n6 1.93989
R924 VDD2.n205 VDD2.t0 1.7777
R925 VDD2.n205 VDD2.t3 1.7777
R926 VDD2.n101 VDD2.t2 1.7777
R927 VDD2.n101 VDD2.t1 1.7777
R928 VDD2 VDD2.n204 1.43584
R929 VDD2.n188 VDD2.n111 1.16414
R930 VDD2.n180 VDD2.n179 1.16414
R931 VDD2.n140 VDD2.n134 1.16414
R932 VDD2.n36 VDD2.n30 1.16414
R933 VDD2.n77 VDD2.n75 1.16414
R934 VDD2.n85 VDD2.n8 1.16414
R935 VDD2.n185 VDD2.n184 0.388379
R936 VDD2.n115 VDD2.n113 0.388379
R937 VDD2.n139 VDD2.n136 0.388379
R938 VDD2.n35 VDD2.n32 0.388379
R939 VDD2.n76 VDD2.n10 0.388379
R940 VDD2.n82 VDD2.n81 0.388379
R941 VDD2.n202 VDD2.n104 0.155672
R942 VDD2.n195 VDD2.n104 0.155672
R943 VDD2.n195 VDD2.n194 0.155672
R944 VDD2.n194 VDD2.n108 0.155672
R945 VDD2.n187 VDD2.n108 0.155672
R946 VDD2.n187 VDD2.n186 0.155672
R947 VDD2.n186 VDD2.n112 0.155672
R948 VDD2.n178 VDD2.n112 0.155672
R949 VDD2.n178 VDD2.n177 0.155672
R950 VDD2.n177 VDD2.n117 0.155672
R951 VDD2.n170 VDD2.n117 0.155672
R952 VDD2.n170 VDD2.n169 0.155672
R953 VDD2.n169 VDD2.n121 0.155672
R954 VDD2.n162 VDD2.n121 0.155672
R955 VDD2.n162 VDD2.n161 0.155672
R956 VDD2.n161 VDD2.n125 0.155672
R957 VDD2.n154 VDD2.n125 0.155672
R958 VDD2.n154 VDD2.n153 0.155672
R959 VDD2.n153 VDD2.n129 0.155672
R960 VDD2.n146 VDD2.n129 0.155672
R961 VDD2.n146 VDD2.n145 0.155672
R962 VDD2.n145 VDD2.n133 0.155672
R963 VDD2.n138 VDD2.n133 0.155672
R964 VDD2.n34 VDD2.n29 0.155672
R965 VDD2.n41 VDD2.n29 0.155672
R966 VDD2.n42 VDD2.n41 0.155672
R967 VDD2.n42 VDD2.n25 0.155672
R968 VDD2.n49 VDD2.n25 0.155672
R969 VDD2.n50 VDD2.n49 0.155672
R970 VDD2.n50 VDD2.n21 0.155672
R971 VDD2.n57 VDD2.n21 0.155672
R972 VDD2.n58 VDD2.n57 0.155672
R973 VDD2.n58 VDD2.n17 0.155672
R974 VDD2.n65 VDD2.n17 0.155672
R975 VDD2.n66 VDD2.n65 0.155672
R976 VDD2.n66 VDD2.n13 0.155672
R977 VDD2.n73 VDD2.n13 0.155672
R978 VDD2.n74 VDD2.n73 0.155672
R979 VDD2.n74 VDD2.n9 0.155672
R980 VDD2.n83 VDD2.n9 0.155672
R981 VDD2.n84 VDD2.n83 0.155672
R982 VDD2.n84 VDD2.n5 0.155672
R983 VDD2.n91 VDD2.n5 0.155672
R984 VDD2.n92 VDD2.n91 0.155672
R985 VDD2.n92 VDD2.n1 0.155672
R986 VDD2.n99 VDD2.n1 0.155672
R987 VP.n7 VP.t0 281.091
R988 VP.n25 VP.t3 244.883
R989 VP.n18 VP.t5 244.883
R990 VP.n32 VP.t1 244.883
R991 VP.n8 VP.t2 244.883
R992 VP.n15 VP.t4 244.883
R993 VP.n18 VP.n17 179.406
R994 VP.n33 VP.n32 179.406
R995 VP.n16 VP.n15 179.406
R996 VP.n10 VP.n9 161.3
R997 VP.n11 VP.n6 161.3
R998 VP.n13 VP.n12 161.3
R999 VP.n14 VP.n5 161.3
R1000 VP.n31 VP.n0 161.3
R1001 VP.n30 VP.n29 161.3
R1002 VP.n28 VP.n1 161.3
R1003 VP.n27 VP.n26 161.3
R1004 VP.n25 VP.n2 161.3
R1005 VP.n24 VP.n23 161.3
R1006 VP.n22 VP.n3 161.3
R1007 VP.n21 VP.n20 161.3
R1008 VP.n19 VP.n4 161.3
R1009 VP.n17 VP.n16 50.2467
R1010 VP.n20 VP.n3 46.8066
R1011 VP.n30 VP.n1 46.8066
R1012 VP.n13 VP.n6 46.8066
R1013 VP.n8 VP.n7 44.4618
R1014 VP.n24 VP.n3 34.1802
R1015 VP.n26 VP.n1 34.1802
R1016 VP.n9 VP.n6 34.1802
R1017 VP.n20 VP.n19 24.4675
R1018 VP.n25 VP.n24 24.4675
R1019 VP.n26 VP.n25 24.4675
R1020 VP.n31 VP.n30 24.4675
R1021 VP.n14 VP.n13 24.4675
R1022 VP.n9 VP.n8 24.4675
R1023 VP.n10 VP.n7 12.1055
R1024 VP.n19 VP.n18 6.36192
R1025 VP.n32 VP.n31 6.36192
R1026 VP.n15 VP.n14 6.36192
R1027 VP.n11 VP.n10 0.189894
R1028 VP.n12 VP.n11 0.189894
R1029 VP.n12 VP.n5 0.189894
R1030 VP.n16 VP.n5 0.189894
R1031 VP.n17 VP.n4 0.189894
R1032 VP.n21 VP.n4 0.189894
R1033 VP.n22 VP.n21 0.189894
R1034 VP.n23 VP.n22 0.189894
R1035 VP.n23 VP.n2 0.189894
R1036 VP.n27 VP.n2 0.189894
R1037 VP.n28 VP.n27 0.189894
R1038 VP.n29 VP.n28 0.189894
R1039 VP.n29 VP.n0 0.189894
R1040 VP.n33 VP.n0 0.189894
R1041 VP VP.n33 0.0516364
R1042 VDD1.n96 VDD1.n0 756.745
R1043 VDD1.n197 VDD1.n101 756.745
R1044 VDD1.n97 VDD1.n96 585
R1045 VDD1.n95 VDD1.n94 585
R1046 VDD1.n4 VDD1.n3 585
R1047 VDD1.n89 VDD1.n88 585
R1048 VDD1.n87 VDD1.n86 585
R1049 VDD1.n8 VDD1.n7 585
R1050 VDD1.n81 VDD1.n80 585
R1051 VDD1.n79 VDD1.n10 585
R1052 VDD1.n78 VDD1.n77 585
R1053 VDD1.n13 VDD1.n11 585
R1054 VDD1.n72 VDD1.n71 585
R1055 VDD1.n70 VDD1.n69 585
R1056 VDD1.n17 VDD1.n16 585
R1057 VDD1.n64 VDD1.n63 585
R1058 VDD1.n62 VDD1.n61 585
R1059 VDD1.n21 VDD1.n20 585
R1060 VDD1.n56 VDD1.n55 585
R1061 VDD1.n54 VDD1.n53 585
R1062 VDD1.n25 VDD1.n24 585
R1063 VDD1.n48 VDD1.n47 585
R1064 VDD1.n46 VDD1.n45 585
R1065 VDD1.n29 VDD1.n28 585
R1066 VDD1.n40 VDD1.n39 585
R1067 VDD1.n38 VDD1.n37 585
R1068 VDD1.n33 VDD1.n32 585
R1069 VDD1.n133 VDD1.n132 585
R1070 VDD1.n138 VDD1.n137 585
R1071 VDD1.n140 VDD1.n139 585
R1072 VDD1.n129 VDD1.n128 585
R1073 VDD1.n146 VDD1.n145 585
R1074 VDD1.n148 VDD1.n147 585
R1075 VDD1.n125 VDD1.n124 585
R1076 VDD1.n154 VDD1.n153 585
R1077 VDD1.n156 VDD1.n155 585
R1078 VDD1.n121 VDD1.n120 585
R1079 VDD1.n162 VDD1.n161 585
R1080 VDD1.n164 VDD1.n163 585
R1081 VDD1.n117 VDD1.n116 585
R1082 VDD1.n170 VDD1.n169 585
R1083 VDD1.n172 VDD1.n171 585
R1084 VDD1.n113 VDD1.n112 585
R1085 VDD1.n179 VDD1.n178 585
R1086 VDD1.n180 VDD1.n111 585
R1087 VDD1.n182 VDD1.n181 585
R1088 VDD1.n109 VDD1.n108 585
R1089 VDD1.n188 VDD1.n187 585
R1090 VDD1.n190 VDD1.n189 585
R1091 VDD1.n105 VDD1.n104 585
R1092 VDD1.n196 VDD1.n195 585
R1093 VDD1.n198 VDD1.n197 585
R1094 VDD1.n34 VDD1.t5 327.466
R1095 VDD1.n134 VDD1.t0 327.466
R1096 VDD1.n96 VDD1.n95 171.744
R1097 VDD1.n95 VDD1.n3 171.744
R1098 VDD1.n88 VDD1.n3 171.744
R1099 VDD1.n88 VDD1.n87 171.744
R1100 VDD1.n87 VDD1.n7 171.744
R1101 VDD1.n80 VDD1.n7 171.744
R1102 VDD1.n80 VDD1.n79 171.744
R1103 VDD1.n79 VDD1.n78 171.744
R1104 VDD1.n78 VDD1.n11 171.744
R1105 VDD1.n71 VDD1.n11 171.744
R1106 VDD1.n71 VDD1.n70 171.744
R1107 VDD1.n70 VDD1.n16 171.744
R1108 VDD1.n63 VDD1.n16 171.744
R1109 VDD1.n63 VDD1.n62 171.744
R1110 VDD1.n62 VDD1.n20 171.744
R1111 VDD1.n55 VDD1.n20 171.744
R1112 VDD1.n55 VDD1.n54 171.744
R1113 VDD1.n54 VDD1.n24 171.744
R1114 VDD1.n47 VDD1.n24 171.744
R1115 VDD1.n47 VDD1.n46 171.744
R1116 VDD1.n46 VDD1.n28 171.744
R1117 VDD1.n39 VDD1.n28 171.744
R1118 VDD1.n39 VDD1.n38 171.744
R1119 VDD1.n38 VDD1.n32 171.744
R1120 VDD1.n138 VDD1.n132 171.744
R1121 VDD1.n139 VDD1.n138 171.744
R1122 VDD1.n139 VDD1.n128 171.744
R1123 VDD1.n146 VDD1.n128 171.744
R1124 VDD1.n147 VDD1.n146 171.744
R1125 VDD1.n147 VDD1.n124 171.744
R1126 VDD1.n154 VDD1.n124 171.744
R1127 VDD1.n155 VDD1.n154 171.744
R1128 VDD1.n155 VDD1.n120 171.744
R1129 VDD1.n162 VDD1.n120 171.744
R1130 VDD1.n163 VDD1.n162 171.744
R1131 VDD1.n163 VDD1.n116 171.744
R1132 VDD1.n170 VDD1.n116 171.744
R1133 VDD1.n171 VDD1.n170 171.744
R1134 VDD1.n171 VDD1.n112 171.744
R1135 VDD1.n179 VDD1.n112 171.744
R1136 VDD1.n180 VDD1.n179 171.744
R1137 VDD1.n181 VDD1.n180 171.744
R1138 VDD1.n181 VDD1.n108 171.744
R1139 VDD1.n188 VDD1.n108 171.744
R1140 VDD1.n189 VDD1.n188 171.744
R1141 VDD1.n189 VDD1.n104 171.744
R1142 VDD1.n196 VDD1.n104 171.744
R1143 VDD1.n197 VDD1.n196 171.744
R1144 VDD1.t5 VDD1.n32 85.8723
R1145 VDD1.t0 VDD1.n132 85.8723
R1146 VDD1.n203 VDD1.n202 70.0611
R1147 VDD1.n205 VDD1.n204 69.6574
R1148 VDD1 VDD1.n100 51.2692
R1149 VDD1.n203 VDD1.n201 51.1556
R1150 VDD1.n205 VDD1.n203 46.9513
R1151 VDD1.n34 VDD1.n33 16.3895
R1152 VDD1.n134 VDD1.n133 16.3895
R1153 VDD1.n81 VDD1.n10 13.1884
R1154 VDD1.n182 VDD1.n111 13.1884
R1155 VDD1.n82 VDD1.n8 12.8005
R1156 VDD1.n77 VDD1.n12 12.8005
R1157 VDD1.n37 VDD1.n36 12.8005
R1158 VDD1.n137 VDD1.n136 12.8005
R1159 VDD1.n178 VDD1.n177 12.8005
R1160 VDD1.n183 VDD1.n109 12.8005
R1161 VDD1.n86 VDD1.n85 12.0247
R1162 VDD1.n76 VDD1.n13 12.0247
R1163 VDD1.n40 VDD1.n31 12.0247
R1164 VDD1.n140 VDD1.n131 12.0247
R1165 VDD1.n176 VDD1.n113 12.0247
R1166 VDD1.n187 VDD1.n186 12.0247
R1167 VDD1.n89 VDD1.n6 11.249
R1168 VDD1.n73 VDD1.n72 11.249
R1169 VDD1.n41 VDD1.n29 11.249
R1170 VDD1.n141 VDD1.n129 11.249
R1171 VDD1.n173 VDD1.n172 11.249
R1172 VDD1.n190 VDD1.n107 11.249
R1173 VDD1.n90 VDD1.n4 10.4732
R1174 VDD1.n69 VDD1.n15 10.4732
R1175 VDD1.n45 VDD1.n44 10.4732
R1176 VDD1.n145 VDD1.n144 10.4732
R1177 VDD1.n169 VDD1.n115 10.4732
R1178 VDD1.n191 VDD1.n105 10.4732
R1179 VDD1.n94 VDD1.n93 9.69747
R1180 VDD1.n68 VDD1.n17 9.69747
R1181 VDD1.n48 VDD1.n27 9.69747
R1182 VDD1.n148 VDD1.n127 9.69747
R1183 VDD1.n168 VDD1.n117 9.69747
R1184 VDD1.n195 VDD1.n194 9.69747
R1185 VDD1.n100 VDD1.n99 9.45567
R1186 VDD1.n201 VDD1.n200 9.45567
R1187 VDD1.n60 VDD1.n59 9.3005
R1188 VDD1.n19 VDD1.n18 9.3005
R1189 VDD1.n66 VDD1.n65 9.3005
R1190 VDD1.n68 VDD1.n67 9.3005
R1191 VDD1.n15 VDD1.n14 9.3005
R1192 VDD1.n74 VDD1.n73 9.3005
R1193 VDD1.n76 VDD1.n75 9.3005
R1194 VDD1.n12 VDD1.n9 9.3005
R1195 VDD1.n99 VDD1.n98 9.3005
R1196 VDD1.n2 VDD1.n1 9.3005
R1197 VDD1.n93 VDD1.n92 9.3005
R1198 VDD1.n91 VDD1.n90 9.3005
R1199 VDD1.n6 VDD1.n5 9.3005
R1200 VDD1.n85 VDD1.n84 9.3005
R1201 VDD1.n83 VDD1.n82 9.3005
R1202 VDD1.n58 VDD1.n57 9.3005
R1203 VDD1.n23 VDD1.n22 9.3005
R1204 VDD1.n52 VDD1.n51 9.3005
R1205 VDD1.n50 VDD1.n49 9.3005
R1206 VDD1.n27 VDD1.n26 9.3005
R1207 VDD1.n44 VDD1.n43 9.3005
R1208 VDD1.n42 VDD1.n41 9.3005
R1209 VDD1.n31 VDD1.n30 9.3005
R1210 VDD1.n36 VDD1.n35 9.3005
R1211 VDD1.n200 VDD1.n199 9.3005
R1212 VDD1.n103 VDD1.n102 9.3005
R1213 VDD1.n194 VDD1.n193 9.3005
R1214 VDD1.n192 VDD1.n191 9.3005
R1215 VDD1.n107 VDD1.n106 9.3005
R1216 VDD1.n186 VDD1.n185 9.3005
R1217 VDD1.n184 VDD1.n183 9.3005
R1218 VDD1.n123 VDD1.n122 9.3005
R1219 VDD1.n152 VDD1.n151 9.3005
R1220 VDD1.n150 VDD1.n149 9.3005
R1221 VDD1.n127 VDD1.n126 9.3005
R1222 VDD1.n144 VDD1.n143 9.3005
R1223 VDD1.n142 VDD1.n141 9.3005
R1224 VDD1.n131 VDD1.n130 9.3005
R1225 VDD1.n136 VDD1.n135 9.3005
R1226 VDD1.n158 VDD1.n157 9.3005
R1227 VDD1.n160 VDD1.n159 9.3005
R1228 VDD1.n119 VDD1.n118 9.3005
R1229 VDD1.n166 VDD1.n165 9.3005
R1230 VDD1.n168 VDD1.n167 9.3005
R1231 VDD1.n115 VDD1.n114 9.3005
R1232 VDD1.n174 VDD1.n173 9.3005
R1233 VDD1.n176 VDD1.n175 9.3005
R1234 VDD1.n177 VDD1.n110 9.3005
R1235 VDD1.n97 VDD1.n2 8.92171
R1236 VDD1.n65 VDD1.n64 8.92171
R1237 VDD1.n49 VDD1.n25 8.92171
R1238 VDD1.n149 VDD1.n125 8.92171
R1239 VDD1.n165 VDD1.n164 8.92171
R1240 VDD1.n198 VDD1.n103 8.92171
R1241 VDD1.n98 VDD1.n0 8.14595
R1242 VDD1.n61 VDD1.n19 8.14595
R1243 VDD1.n53 VDD1.n52 8.14595
R1244 VDD1.n153 VDD1.n152 8.14595
R1245 VDD1.n161 VDD1.n119 8.14595
R1246 VDD1.n199 VDD1.n101 8.14595
R1247 VDD1.n60 VDD1.n21 7.3702
R1248 VDD1.n56 VDD1.n23 7.3702
R1249 VDD1.n156 VDD1.n123 7.3702
R1250 VDD1.n160 VDD1.n121 7.3702
R1251 VDD1.n57 VDD1.n21 6.59444
R1252 VDD1.n57 VDD1.n56 6.59444
R1253 VDD1.n157 VDD1.n156 6.59444
R1254 VDD1.n157 VDD1.n121 6.59444
R1255 VDD1.n100 VDD1.n0 5.81868
R1256 VDD1.n61 VDD1.n60 5.81868
R1257 VDD1.n53 VDD1.n23 5.81868
R1258 VDD1.n153 VDD1.n123 5.81868
R1259 VDD1.n161 VDD1.n160 5.81868
R1260 VDD1.n201 VDD1.n101 5.81868
R1261 VDD1.n98 VDD1.n97 5.04292
R1262 VDD1.n64 VDD1.n19 5.04292
R1263 VDD1.n52 VDD1.n25 5.04292
R1264 VDD1.n152 VDD1.n125 5.04292
R1265 VDD1.n164 VDD1.n119 5.04292
R1266 VDD1.n199 VDD1.n198 5.04292
R1267 VDD1.n94 VDD1.n2 4.26717
R1268 VDD1.n65 VDD1.n17 4.26717
R1269 VDD1.n49 VDD1.n48 4.26717
R1270 VDD1.n149 VDD1.n148 4.26717
R1271 VDD1.n165 VDD1.n117 4.26717
R1272 VDD1.n195 VDD1.n103 4.26717
R1273 VDD1.n35 VDD1.n34 3.70982
R1274 VDD1.n135 VDD1.n134 3.70982
R1275 VDD1.n93 VDD1.n4 3.49141
R1276 VDD1.n69 VDD1.n68 3.49141
R1277 VDD1.n45 VDD1.n27 3.49141
R1278 VDD1.n145 VDD1.n127 3.49141
R1279 VDD1.n169 VDD1.n168 3.49141
R1280 VDD1.n194 VDD1.n105 3.49141
R1281 VDD1.n90 VDD1.n89 2.71565
R1282 VDD1.n72 VDD1.n15 2.71565
R1283 VDD1.n44 VDD1.n29 2.71565
R1284 VDD1.n144 VDD1.n129 2.71565
R1285 VDD1.n172 VDD1.n115 2.71565
R1286 VDD1.n191 VDD1.n190 2.71565
R1287 VDD1.n86 VDD1.n6 1.93989
R1288 VDD1.n73 VDD1.n13 1.93989
R1289 VDD1.n41 VDD1.n40 1.93989
R1290 VDD1.n141 VDD1.n140 1.93989
R1291 VDD1.n173 VDD1.n113 1.93989
R1292 VDD1.n187 VDD1.n107 1.93989
R1293 VDD1.n204 VDD1.t3 1.7777
R1294 VDD1.n204 VDD1.t1 1.7777
R1295 VDD1.n202 VDD1.t2 1.7777
R1296 VDD1.n202 VDD1.t4 1.7777
R1297 VDD1.n85 VDD1.n8 1.16414
R1298 VDD1.n77 VDD1.n76 1.16414
R1299 VDD1.n37 VDD1.n31 1.16414
R1300 VDD1.n137 VDD1.n131 1.16414
R1301 VDD1.n178 VDD1.n176 1.16414
R1302 VDD1.n186 VDD1.n109 1.16414
R1303 VDD1 VDD1.n205 0.401362
R1304 VDD1.n82 VDD1.n81 0.388379
R1305 VDD1.n12 VDD1.n10 0.388379
R1306 VDD1.n36 VDD1.n33 0.388379
R1307 VDD1.n136 VDD1.n133 0.388379
R1308 VDD1.n177 VDD1.n111 0.388379
R1309 VDD1.n183 VDD1.n182 0.388379
R1310 VDD1.n99 VDD1.n1 0.155672
R1311 VDD1.n92 VDD1.n1 0.155672
R1312 VDD1.n92 VDD1.n91 0.155672
R1313 VDD1.n91 VDD1.n5 0.155672
R1314 VDD1.n84 VDD1.n5 0.155672
R1315 VDD1.n84 VDD1.n83 0.155672
R1316 VDD1.n83 VDD1.n9 0.155672
R1317 VDD1.n75 VDD1.n9 0.155672
R1318 VDD1.n75 VDD1.n74 0.155672
R1319 VDD1.n74 VDD1.n14 0.155672
R1320 VDD1.n67 VDD1.n14 0.155672
R1321 VDD1.n67 VDD1.n66 0.155672
R1322 VDD1.n66 VDD1.n18 0.155672
R1323 VDD1.n59 VDD1.n18 0.155672
R1324 VDD1.n59 VDD1.n58 0.155672
R1325 VDD1.n58 VDD1.n22 0.155672
R1326 VDD1.n51 VDD1.n22 0.155672
R1327 VDD1.n51 VDD1.n50 0.155672
R1328 VDD1.n50 VDD1.n26 0.155672
R1329 VDD1.n43 VDD1.n26 0.155672
R1330 VDD1.n43 VDD1.n42 0.155672
R1331 VDD1.n42 VDD1.n30 0.155672
R1332 VDD1.n35 VDD1.n30 0.155672
R1333 VDD1.n135 VDD1.n130 0.155672
R1334 VDD1.n142 VDD1.n130 0.155672
R1335 VDD1.n143 VDD1.n142 0.155672
R1336 VDD1.n143 VDD1.n126 0.155672
R1337 VDD1.n150 VDD1.n126 0.155672
R1338 VDD1.n151 VDD1.n150 0.155672
R1339 VDD1.n151 VDD1.n122 0.155672
R1340 VDD1.n158 VDD1.n122 0.155672
R1341 VDD1.n159 VDD1.n158 0.155672
R1342 VDD1.n159 VDD1.n118 0.155672
R1343 VDD1.n166 VDD1.n118 0.155672
R1344 VDD1.n167 VDD1.n166 0.155672
R1345 VDD1.n167 VDD1.n114 0.155672
R1346 VDD1.n174 VDD1.n114 0.155672
R1347 VDD1.n175 VDD1.n174 0.155672
R1348 VDD1.n175 VDD1.n110 0.155672
R1349 VDD1.n184 VDD1.n110 0.155672
R1350 VDD1.n185 VDD1.n184 0.155672
R1351 VDD1.n185 VDD1.n106 0.155672
R1352 VDD1.n192 VDD1.n106 0.155672
R1353 VDD1.n193 VDD1.n192 0.155672
R1354 VDD1.n193 VDD1.n102 0.155672
R1355 VDD1.n200 VDD1.n102 0.155672
R1356 B.n553 B.n88 585
R1357 B.n555 B.n554 585
R1358 B.n556 B.n87 585
R1359 B.n558 B.n557 585
R1360 B.n559 B.n86 585
R1361 B.n561 B.n560 585
R1362 B.n562 B.n85 585
R1363 B.n564 B.n563 585
R1364 B.n565 B.n84 585
R1365 B.n567 B.n566 585
R1366 B.n568 B.n83 585
R1367 B.n570 B.n569 585
R1368 B.n571 B.n82 585
R1369 B.n573 B.n572 585
R1370 B.n574 B.n81 585
R1371 B.n576 B.n575 585
R1372 B.n577 B.n80 585
R1373 B.n579 B.n578 585
R1374 B.n580 B.n79 585
R1375 B.n582 B.n581 585
R1376 B.n583 B.n78 585
R1377 B.n585 B.n584 585
R1378 B.n586 B.n77 585
R1379 B.n588 B.n587 585
R1380 B.n589 B.n76 585
R1381 B.n591 B.n590 585
R1382 B.n592 B.n75 585
R1383 B.n594 B.n593 585
R1384 B.n595 B.n74 585
R1385 B.n597 B.n596 585
R1386 B.n598 B.n73 585
R1387 B.n600 B.n599 585
R1388 B.n601 B.n72 585
R1389 B.n603 B.n602 585
R1390 B.n604 B.n71 585
R1391 B.n606 B.n605 585
R1392 B.n607 B.n70 585
R1393 B.n609 B.n608 585
R1394 B.n610 B.n69 585
R1395 B.n612 B.n611 585
R1396 B.n613 B.n68 585
R1397 B.n615 B.n614 585
R1398 B.n616 B.n67 585
R1399 B.n618 B.n617 585
R1400 B.n619 B.n66 585
R1401 B.n621 B.n620 585
R1402 B.n622 B.n65 585
R1403 B.n624 B.n623 585
R1404 B.n625 B.n64 585
R1405 B.n627 B.n626 585
R1406 B.n628 B.n63 585
R1407 B.n630 B.n629 585
R1408 B.n631 B.n62 585
R1409 B.n633 B.n632 585
R1410 B.n634 B.n61 585
R1411 B.n636 B.n635 585
R1412 B.n637 B.n60 585
R1413 B.n639 B.n638 585
R1414 B.n640 B.n59 585
R1415 B.n642 B.n641 585
R1416 B.n644 B.n56 585
R1417 B.n646 B.n645 585
R1418 B.n647 B.n55 585
R1419 B.n649 B.n648 585
R1420 B.n650 B.n54 585
R1421 B.n652 B.n651 585
R1422 B.n653 B.n53 585
R1423 B.n655 B.n654 585
R1424 B.n656 B.n49 585
R1425 B.n658 B.n657 585
R1426 B.n659 B.n48 585
R1427 B.n661 B.n660 585
R1428 B.n662 B.n47 585
R1429 B.n664 B.n663 585
R1430 B.n665 B.n46 585
R1431 B.n667 B.n666 585
R1432 B.n668 B.n45 585
R1433 B.n670 B.n669 585
R1434 B.n671 B.n44 585
R1435 B.n673 B.n672 585
R1436 B.n674 B.n43 585
R1437 B.n676 B.n675 585
R1438 B.n677 B.n42 585
R1439 B.n679 B.n678 585
R1440 B.n680 B.n41 585
R1441 B.n682 B.n681 585
R1442 B.n683 B.n40 585
R1443 B.n685 B.n684 585
R1444 B.n686 B.n39 585
R1445 B.n688 B.n687 585
R1446 B.n689 B.n38 585
R1447 B.n691 B.n690 585
R1448 B.n692 B.n37 585
R1449 B.n694 B.n693 585
R1450 B.n695 B.n36 585
R1451 B.n697 B.n696 585
R1452 B.n698 B.n35 585
R1453 B.n700 B.n699 585
R1454 B.n701 B.n34 585
R1455 B.n703 B.n702 585
R1456 B.n704 B.n33 585
R1457 B.n706 B.n705 585
R1458 B.n707 B.n32 585
R1459 B.n709 B.n708 585
R1460 B.n710 B.n31 585
R1461 B.n712 B.n711 585
R1462 B.n713 B.n30 585
R1463 B.n715 B.n714 585
R1464 B.n716 B.n29 585
R1465 B.n718 B.n717 585
R1466 B.n719 B.n28 585
R1467 B.n721 B.n720 585
R1468 B.n722 B.n27 585
R1469 B.n724 B.n723 585
R1470 B.n725 B.n26 585
R1471 B.n727 B.n726 585
R1472 B.n728 B.n25 585
R1473 B.n730 B.n729 585
R1474 B.n731 B.n24 585
R1475 B.n733 B.n732 585
R1476 B.n734 B.n23 585
R1477 B.n736 B.n735 585
R1478 B.n737 B.n22 585
R1479 B.n739 B.n738 585
R1480 B.n740 B.n21 585
R1481 B.n742 B.n741 585
R1482 B.n743 B.n20 585
R1483 B.n745 B.n744 585
R1484 B.n746 B.n19 585
R1485 B.n748 B.n747 585
R1486 B.n552 B.n551 585
R1487 B.n550 B.n89 585
R1488 B.n549 B.n548 585
R1489 B.n547 B.n90 585
R1490 B.n546 B.n545 585
R1491 B.n544 B.n91 585
R1492 B.n543 B.n542 585
R1493 B.n541 B.n92 585
R1494 B.n540 B.n539 585
R1495 B.n538 B.n93 585
R1496 B.n537 B.n536 585
R1497 B.n535 B.n94 585
R1498 B.n534 B.n533 585
R1499 B.n532 B.n95 585
R1500 B.n531 B.n530 585
R1501 B.n529 B.n96 585
R1502 B.n528 B.n527 585
R1503 B.n526 B.n97 585
R1504 B.n525 B.n524 585
R1505 B.n523 B.n98 585
R1506 B.n522 B.n521 585
R1507 B.n520 B.n99 585
R1508 B.n519 B.n518 585
R1509 B.n517 B.n100 585
R1510 B.n516 B.n515 585
R1511 B.n514 B.n101 585
R1512 B.n513 B.n512 585
R1513 B.n511 B.n102 585
R1514 B.n510 B.n509 585
R1515 B.n508 B.n103 585
R1516 B.n507 B.n506 585
R1517 B.n505 B.n104 585
R1518 B.n504 B.n503 585
R1519 B.n502 B.n105 585
R1520 B.n501 B.n500 585
R1521 B.n499 B.n106 585
R1522 B.n498 B.n497 585
R1523 B.n496 B.n107 585
R1524 B.n495 B.n494 585
R1525 B.n493 B.n108 585
R1526 B.n492 B.n491 585
R1527 B.n490 B.n109 585
R1528 B.n489 B.n488 585
R1529 B.n487 B.n110 585
R1530 B.n486 B.n485 585
R1531 B.n484 B.n111 585
R1532 B.n483 B.n482 585
R1533 B.n481 B.n112 585
R1534 B.n480 B.n479 585
R1535 B.n478 B.n113 585
R1536 B.n477 B.n476 585
R1537 B.n475 B.n114 585
R1538 B.n474 B.n473 585
R1539 B.n472 B.n115 585
R1540 B.n471 B.n470 585
R1541 B.n469 B.n116 585
R1542 B.n468 B.n467 585
R1543 B.n466 B.n117 585
R1544 B.n465 B.n464 585
R1545 B.n463 B.n118 585
R1546 B.n462 B.n461 585
R1547 B.n460 B.n119 585
R1548 B.n459 B.n458 585
R1549 B.n457 B.n120 585
R1550 B.n456 B.n455 585
R1551 B.n454 B.n121 585
R1552 B.n453 B.n452 585
R1553 B.n256 B.n191 585
R1554 B.n258 B.n257 585
R1555 B.n259 B.n190 585
R1556 B.n261 B.n260 585
R1557 B.n262 B.n189 585
R1558 B.n264 B.n263 585
R1559 B.n265 B.n188 585
R1560 B.n267 B.n266 585
R1561 B.n268 B.n187 585
R1562 B.n270 B.n269 585
R1563 B.n271 B.n186 585
R1564 B.n273 B.n272 585
R1565 B.n274 B.n185 585
R1566 B.n276 B.n275 585
R1567 B.n277 B.n184 585
R1568 B.n279 B.n278 585
R1569 B.n280 B.n183 585
R1570 B.n282 B.n281 585
R1571 B.n283 B.n182 585
R1572 B.n285 B.n284 585
R1573 B.n286 B.n181 585
R1574 B.n288 B.n287 585
R1575 B.n289 B.n180 585
R1576 B.n291 B.n290 585
R1577 B.n292 B.n179 585
R1578 B.n294 B.n293 585
R1579 B.n295 B.n178 585
R1580 B.n297 B.n296 585
R1581 B.n298 B.n177 585
R1582 B.n300 B.n299 585
R1583 B.n301 B.n176 585
R1584 B.n303 B.n302 585
R1585 B.n304 B.n175 585
R1586 B.n306 B.n305 585
R1587 B.n307 B.n174 585
R1588 B.n309 B.n308 585
R1589 B.n310 B.n173 585
R1590 B.n312 B.n311 585
R1591 B.n313 B.n172 585
R1592 B.n315 B.n314 585
R1593 B.n316 B.n171 585
R1594 B.n318 B.n317 585
R1595 B.n319 B.n170 585
R1596 B.n321 B.n320 585
R1597 B.n322 B.n169 585
R1598 B.n324 B.n323 585
R1599 B.n325 B.n168 585
R1600 B.n327 B.n326 585
R1601 B.n328 B.n167 585
R1602 B.n330 B.n329 585
R1603 B.n331 B.n166 585
R1604 B.n333 B.n332 585
R1605 B.n334 B.n165 585
R1606 B.n336 B.n335 585
R1607 B.n337 B.n164 585
R1608 B.n339 B.n338 585
R1609 B.n340 B.n163 585
R1610 B.n342 B.n341 585
R1611 B.n343 B.n162 585
R1612 B.n345 B.n344 585
R1613 B.n347 B.n346 585
R1614 B.n348 B.n158 585
R1615 B.n350 B.n349 585
R1616 B.n351 B.n157 585
R1617 B.n353 B.n352 585
R1618 B.n354 B.n156 585
R1619 B.n356 B.n355 585
R1620 B.n357 B.n155 585
R1621 B.n359 B.n358 585
R1622 B.n360 B.n152 585
R1623 B.n363 B.n362 585
R1624 B.n364 B.n151 585
R1625 B.n366 B.n365 585
R1626 B.n367 B.n150 585
R1627 B.n369 B.n368 585
R1628 B.n370 B.n149 585
R1629 B.n372 B.n371 585
R1630 B.n373 B.n148 585
R1631 B.n375 B.n374 585
R1632 B.n376 B.n147 585
R1633 B.n378 B.n377 585
R1634 B.n379 B.n146 585
R1635 B.n381 B.n380 585
R1636 B.n382 B.n145 585
R1637 B.n384 B.n383 585
R1638 B.n385 B.n144 585
R1639 B.n387 B.n386 585
R1640 B.n388 B.n143 585
R1641 B.n390 B.n389 585
R1642 B.n391 B.n142 585
R1643 B.n393 B.n392 585
R1644 B.n394 B.n141 585
R1645 B.n396 B.n395 585
R1646 B.n397 B.n140 585
R1647 B.n399 B.n398 585
R1648 B.n400 B.n139 585
R1649 B.n402 B.n401 585
R1650 B.n403 B.n138 585
R1651 B.n405 B.n404 585
R1652 B.n406 B.n137 585
R1653 B.n408 B.n407 585
R1654 B.n409 B.n136 585
R1655 B.n411 B.n410 585
R1656 B.n412 B.n135 585
R1657 B.n414 B.n413 585
R1658 B.n415 B.n134 585
R1659 B.n417 B.n416 585
R1660 B.n418 B.n133 585
R1661 B.n420 B.n419 585
R1662 B.n421 B.n132 585
R1663 B.n423 B.n422 585
R1664 B.n424 B.n131 585
R1665 B.n426 B.n425 585
R1666 B.n427 B.n130 585
R1667 B.n429 B.n428 585
R1668 B.n430 B.n129 585
R1669 B.n432 B.n431 585
R1670 B.n433 B.n128 585
R1671 B.n435 B.n434 585
R1672 B.n436 B.n127 585
R1673 B.n438 B.n437 585
R1674 B.n439 B.n126 585
R1675 B.n441 B.n440 585
R1676 B.n442 B.n125 585
R1677 B.n444 B.n443 585
R1678 B.n445 B.n124 585
R1679 B.n447 B.n446 585
R1680 B.n448 B.n123 585
R1681 B.n450 B.n449 585
R1682 B.n451 B.n122 585
R1683 B.n255 B.n254 585
R1684 B.n253 B.n192 585
R1685 B.n252 B.n251 585
R1686 B.n250 B.n193 585
R1687 B.n249 B.n248 585
R1688 B.n247 B.n194 585
R1689 B.n246 B.n245 585
R1690 B.n244 B.n195 585
R1691 B.n243 B.n242 585
R1692 B.n241 B.n196 585
R1693 B.n240 B.n239 585
R1694 B.n238 B.n197 585
R1695 B.n237 B.n236 585
R1696 B.n235 B.n198 585
R1697 B.n234 B.n233 585
R1698 B.n232 B.n199 585
R1699 B.n231 B.n230 585
R1700 B.n229 B.n200 585
R1701 B.n228 B.n227 585
R1702 B.n226 B.n201 585
R1703 B.n225 B.n224 585
R1704 B.n223 B.n202 585
R1705 B.n222 B.n221 585
R1706 B.n220 B.n203 585
R1707 B.n219 B.n218 585
R1708 B.n217 B.n204 585
R1709 B.n216 B.n215 585
R1710 B.n214 B.n205 585
R1711 B.n213 B.n212 585
R1712 B.n211 B.n206 585
R1713 B.n210 B.n209 585
R1714 B.n208 B.n207 585
R1715 B.n2 B.n0 585
R1716 B.n797 B.n1 585
R1717 B.n796 B.n795 585
R1718 B.n794 B.n3 585
R1719 B.n793 B.n792 585
R1720 B.n791 B.n4 585
R1721 B.n790 B.n789 585
R1722 B.n788 B.n5 585
R1723 B.n787 B.n786 585
R1724 B.n785 B.n6 585
R1725 B.n784 B.n783 585
R1726 B.n782 B.n7 585
R1727 B.n781 B.n780 585
R1728 B.n779 B.n8 585
R1729 B.n778 B.n777 585
R1730 B.n776 B.n9 585
R1731 B.n775 B.n774 585
R1732 B.n773 B.n10 585
R1733 B.n772 B.n771 585
R1734 B.n770 B.n11 585
R1735 B.n769 B.n768 585
R1736 B.n767 B.n12 585
R1737 B.n766 B.n765 585
R1738 B.n764 B.n13 585
R1739 B.n763 B.n762 585
R1740 B.n761 B.n14 585
R1741 B.n760 B.n759 585
R1742 B.n758 B.n15 585
R1743 B.n757 B.n756 585
R1744 B.n755 B.n16 585
R1745 B.n754 B.n753 585
R1746 B.n752 B.n17 585
R1747 B.n751 B.n750 585
R1748 B.n749 B.n18 585
R1749 B.n799 B.n798 585
R1750 B.n153 B.t11 530.367
R1751 B.n57 B.t1 530.367
R1752 B.n159 B.t8 530.367
R1753 B.n50 B.t4 530.367
R1754 B.n256 B.n255 511.721
R1755 B.n749 B.n748 511.721
R1756 B.n453 B.n122 511.721
R1757 B.n551 B.n88 511.721
R1758 B.n154 B.t10 489.058
R1759 B.n58 B.t2 489.058
R1760 B.n160 B.t7 489.058
R1761 B.n51 B.t5 489.058
R1762 B.n153 B.t9 451.289
R1763 B.n159 B.t6 451.289
R1764 B.n50 B.t3 451.289
R1765 B.n57 B.t0 451.289
R1766 B.n255 B.n192 163.367
R1767 B.n251 B.n192 163.367
R1768 B.n251 B.n250 163.367
R1769 B.n250 B.n249 163.367
R1770 B.n249 B.n194 163.367
R1771 B.n245 B.n194 163.367
R1772 B.n245 B.n244 163.367
R1773 B.n244 B.n243 163.367
R1774 B.n243 B.n196 163.367
R1775 B.n239 B.n196 163.367
R1776 B.n239 B.n238 163.367
R1777 B.n238 B.n237 163.367
R1778 B.n237 B.n198 163.367
R1779 B.n233 B.n198 163.367
R1780 B.n233 B.n232 163.367
R1781 B.n232 B.n231 163.367
R1782 B.n231 B.n200 163.367
R1783 B.n227 B.n200 163.367
R1784 B.n227 B.n226 163.367
R1785 B.n226 B.n225 163.367
R1786 B.n225 B.n202 163.367
R1787 B.n221 B.n202 163.367
R1788 B.n221 B.n220 163.367
R1789 B.n220 B.n219 163.367
R1790 B.n219 B.n204 163.367
R1791 B.n215 B.n204 163.367
R1792 B.n215 B.n214 163.367
R1793 B.n214 B.n213 163.367
R1794 B.n213 B.n206 163.367
R1795 B.n209 B.n206 163.367
R1796 B.n209 B.n208 163.367
R1797 B.n208 B.n2 163.367
R1798 B.n798 B.n2 163.367
R1799 B.n798 B.n797 163.367
R1800 B.n797 B.n796 163.367
R1801 B.n796 B.n3 163.367
R1802 B.n792 B.n3 163.367
R1803 B.n792 B.n791 163.367
R1804 B.n791 B.n790 163.367
R1805 B.n790 B.n5 163.367
R1806 B.n786 B.n5 163.367
R1807 B.n786 B.n785 163.367
R1808 B.n785 B.n784 163.367
R1809 B.n784 B.n7 163.367
R1810 B.n780 B.n7 163.367
R1811 B.n780 B.n779 163.367
R1812 B.n779 B.n778 163.367
R1813 B.n778 B.n9 163.367
R1814 B.n774 B.n9 163.367
R1815 B.n774 B.n773 163.367
R1816 B.n773 B.n772 163.367
R1817 B.n772 B.n11 163.367
R1818 B.n768 B.n11 163.367
R1819 B.n768 B.n767 163.367
R1820 B.n767 B.n766 163.367
R1821 B.n766 B.n13 163.367
R1822 B.n762 B.n13 163.367
R1823 B.n762 B.n761 163.367
R1824 B.n761 B.n760 163.367
R1825 B.n760 B.n15 163.367
R1826 B.n756 B.n15 163.367
R1827 B.n756 B.n755 163.367
R1828 B.n755 B.n754 163.367
R1829 B.n754 B.n17 163.367
R1830 B.n750 B.n17 163.367
R1831 B.n750 B.n749 163.367
R1832 B.n257 B.n256 163.367
R1833 B.n257 B.n190 163.367
R1834 B.n261 B.n190 163.367
R1835 B.n262 B.n261 163.367
R1836 B.n263 B.n262 163.367
R1837 B.n263 B.n188 163.367
R1838 B.n267 B.n188 163.367
R1839 B.n268 B.n267 163.367
R1840 B.n269 B.n268 163.367
R1841 B.n269 B.n186 163.367
R1842 B.n273 B.n186 163.367
R1843 B.n274 B.n273 163.367
R1844 B.n275 B.n274 163.367
R1845 B.n275 B.n184 163.367
R1846 B.n279 B.n184 163.367
R1847 B.n280 B.n279 163.367
R1848 B.n281 B.n280 163.367
R1849 B.n281 B.n182 163.367
R1850 B.n285 B.n182 163.367
R1851 B.n286 B.n285 163.367
R1852 B.n287 B.n286 163.367
R1853 B.n287 B.n180 163.367
R1854 B.n291 B.n180 163.367
R1855 B.n292 B.n291 163.367
R1856 B.n293 B.n292 163.367
R1857 B.n293 B.n178 163.367
R1858 B.n297 B.n178 163.367
R1859 B.n298 B.n297 163.367
R1860 B.n299 B.n298 163.367
R1861 B.n299 B.n176 163.367
R1862 B.n303 B.n176 163.367
R1863 B.n304 B.n303 163.367
R1864 B.n305 B.n304 163.367
R1865 B.n305 B.n174 163.367
R1866 B.n309 B.n174 163.367
R1867 B.n310 B.n309 163.367
R1868 B.n311 B.n310 163.367
R1869 B.n311 B.n172 163.367
R1870 B.n315 B.n172 163.367
R1871 B.n316 B.n315 163.367
R1872 B.n317 B.n316 163.367
R1873 B.n317 B.n170 163.367
R1874 B.n321 B.n170 163.367
R1875 B.n322 B.n321 163.367
R1876 B.n323 B.n322 163.367
R1877 B.n323 B.n168 163.367
R1878 B.n327 B.n168 163.367
R1879 B.n328 B.n327 163.367
R1880 B.n329 B.n328 163.367
R1881 B.n329 B.n166 163.367
R1882 B.n333 B.n166 163.367
R1883 B.n334 B.n333 163.367
R1884 B.n335 B.n334 163.367
R1885 B.n335 B.n164 163.367
R1886 B.n339 B.n164 163.367
R1887 B.n340 B.n339 163.367
R1888 B.n341 B.n340 163.367
R1889 B.n341 B.n162 163.367
R1890 B.n345 B.n162 163.367
R1891 B.n346 B.n345 163.367
R1892 B.n346 B.n158 163.367
R1893 B.n350 B.n158 163.367
R1894 B.n351 B.n350 163.367
R1895 B.n352 B.n351 163.367
R1896 B.n352 B.n156 163.367
R1897 B.n356 B.n156 163.367
R1898 B.n357 B.n356 163.367
R1899 B.n358 B.n357 163.367
R1900 B.n358 B.n152 163.367
R1901 B.n363 B.n152 163.367
R1902 B.n364 B.n363 163.367
R1903 B.n365 B.n364 163.367
R1904 B.n365 B.n150 163.367
R1905 B.n369 B.n150 163.367
R1906 B.n370 B.n369 163.367
R1907 B.n371 B.n370 163.367
R1908 B.n371 B.n148 163.367
R1909 B.n375 B.n148 163.367
R1910 B.n376 B.n375 163.367
R1911 B.n377 B.n376 163.367
R1912 B.n377 B.n146 163.367
R1913 B.n381 B.n146 163.367
R1914 B.n382 B.n381 163.367
R1915 B.n383 B.n382 163.367
R1916 B.n383 B.n144 163.367
R1917 B.n387 B.n144 163.367
R1918 B.n388 B.n387 163.367
R1919 B.n389 B.n388 163.367
R1920 B.n389 B.n142 163.367
R1921 B.n393 B.n142 163.367
R1922 B.n394 B.n393 163.367
R1923 B.n395 B.n394 163.367
R1924 B.n395 B.n140 163.367
R1925 B.n399 B.n140 163.367
R1926 B.n400 B.n399 163.367
R1927 B.n401 B.n400 163.367
R1928 B.n401 B.n138 163.367
R1929 B.n405 B.n138 163.367
R1930 B.n406 B.n405 163.367
R1931 B.n407 B.n406 163.367
R1932 B.n407 B.n136 163.367
R1933 B.n411 B.n136 163.367
R1934 B.n412 B.n411 163.367
R1935 B.n413 B.n412 163.367
R1936 B.n413 B.n134 163.367
R1937 B.n417 B.n134 163.367
R1938 B.n418 B.n417 163.367
R1939 B.n419 B.n418 163.367
R1940 B.n419 B.n132 163.367
R1941 B.n423 B.n132 163.367
R1942 B.n424 B.n423 163.367
R1943 B.n425 B.n424 163.367
R1944 B.n425 B.n130 163.367
R1945 B.n429 B.n130 163.367
R1946 B.n430 B.n429 163.367
R1947 B.n431 B.n430 163.367
R1948 B.n431 B.n128 163.367
R1949 B.n435 B.n128 163.367
R1950 B.n436 B.n435 163.367
R1951 B.n437 B.n436 163.367
R1952 B.n437 B.n126 163.367
R1953 B.n441 B.n126 163.367
R1954 B.n442 B.n441 163.367
R1955 B.n443 B.n442 163.367
R1956 B.n443 B.n124 163.367
R1957 B.n447 B.n124 163.367
R1958 B.n448 B.n447 163.367
R1959 B.n449 B.n448 163.367
R1960 B.n449 B.n122 163.367
R1961 B.n454 B.n453 163.367
R1962 B.n455 B.n454 163.367
R1963 B.n455 B.n120 163.367
R1964 B.n459 B.n120 163.367
R1965 B.n460 B.n459 163.367
R1966 B.n461 B.n460 163.367
R1967 B.n461 B.n118 163.367
R1968 B.n465 B.n118 163.367
R1969 B.n466 B.n465 163.367
R1970 B.n467 B.n466 163.367
R1971 B.n467 B.n116 163.367
R1972 B.n471 B.n116 163.367
R1973 B.n472 B.n471 163.367
R1974 B.n473 B.n472 163.367
R1975 B.n473 B.n114 163.367
R1976 B.n477 B.n114 163.367
R1977 B.n478 B.n477 163.367
R1978 B.n479 B.n478 163.367
R1979 B.n479 B.n112 163.367
R1980 B.n483 B.n112 163.367
R1981 B.n484 B.n483 163.367
R1982 B.n485 B.n484 163.367
R1983 B.n485 B.n110 163.367
R1984 B.n489 B.n110 163.367
R1985 B.n490 B.n489 163.367
R1986 B.n491 B.n490 163.367
R1987 B.n491 B.n108 163.367
R1988 B.n495 B.n108 163.367
R1989 B.n496 B.n495 163.367
R1990 B.n497 B.n496 163.367
R1991 B.n497 B.n106 163.367
R1992 B.n501 B.n106 163.367
R1993 B.n502 B.n501 163.367
R1994 B.n503 B.n502 163.367
R1995 B.n503 B.n104 163.367
R1996 B.n507 B.n104 163.367
R1997 B.n508 B.n507 163.367
R1998 B.n509 B.n508 163.367
R1999 B.n509 B.n102 163.367
R2000 B.n513 B.n102 163.367
R2001 B.n514 B.n513 163.367
R2002 B.n515 B.n514 163.367
R2003 B.n515 B.n100 163.367
R2004 B.n519 B.n100 163.367
R2005 B.n520 B.n519 163.367
R2006 B.n521 B.n520 163.367
R2007 B.n521 B.n98 163.367
R2008 B.n525 B.n98 163.367
R2009 B.n526 B.n525 163.367
R2010 B.n527 B.n526 163.367
R2011 B.n527 B.n96 163.367
R2012 B.n531 B.n96 163.367
R2013 B.n532 B.n531 163.367
R2014 B.n533 B.n532 163.367
R2015 B.n533 B.n94 163.367
R2016 B.n537 B.n94 163.367
R2017 B.n538 B.n537 163.367
R2018 B.n539 B.n538 163.367
R2019 B.n539 B.n92 163.367
R2020 B.n543 B.n92 163.367
R2021 B.n544 B.n543 163.367
R2022 B.n545 B.n544 163.367
R2023 B.n545 B.n90 163.367
R2024 B.n549 B.n90 163.367
R2025 B.n550 B.n549 163.367
R2026 B.n551 B.n550 163.367
R2027 B.n748 B.n19 163.367
R2028 B.n744 B.n19 163.367
R2029 B.n744 B.n743 163.367
R2030 B.n743 B.n742 163.367
R2031 B.n742 B.n21 163.367
R2032 B.n738 B.n21 163.367
R2033 B.n738 B.n737 163.367
R2034 B.n737 B.n736 163.367
R2035 B.n736 B.n23 163.367
R2036 B.n732 B.n23 163.367
R2037 B.n732 B.n731 163.367
R2038 B.n731 B.n730 163.367
R2039 B.n730 B.n25 163.367
R2040 B.n726 B.n25 163.367
R2041 B.n726 B.n725 163.367
R2042 B.n725 B.n724 163.367
R2043 B.n724 B.n27 163.367
R2044 B.n720 B.n27 163.367
R2045 B.n720 B.n719 163.367
R2046 B.n719 B.n718 163.367
R2047 B.n718 B.n29 163.367
R2048 B.n714 B.n29 163.367
R2049 B.n714 B.n713 163.367
R2050 B.n713 B.n712 163.367
R2051 B.n712 B.n31 163.367
R2052 B.n708 B.n31 163.367
R2053 B.n708 B.n707 163.367
R2054 B.n707 B.n706 163.367
R2055 B.n706 B.n33 163.367
R2056 B.n702 B.n33 163.367
R2057 B.n702 B.n701 163.367
R2058 B.n701 B.n700 163.367
R2059 B.n700 B.n35 163.367
R2060 B.n696 B.n35 163.367
R2061 B.n696 B.n695 163.367
R2062 B.n695 B.n694 163.367
R2063 B.n694 B.n37 163.367
R2064 B.n690 B.n37 163.367
R2065 B.n690 B.n689 163.367
R2066 B.n689 B.n688 163.367
R2067 B.n688 B.n39 163.367
R2068 B.n684 B.n39 163.367
R2069 B.n684 B.n683 163.367
R2070 B.n683 B.n682 163.367
R2071 B.n682 B.n41 163.367
R2072 B.n678 B.n41 163.367
R2073 B.n678 B.n677 163.367
R2074 B.n677 B.n676 163.367
R2075 B.n676 B.n43 163.367
R2076 B.n672 B.n43 163.367
R2077 B.n672 B.n671 163.367
R2078 B.n671 B.n670 163.367
R2079 B.n670 B.n45 163.367
R2080 B.n666 B.n45 163.367
R2081 B.n666 B.n665 163.367
R2082 B.n665 B.n664 163.367
R2083 B.n664 B.n47 163.367
R2084 B.n660 B.n47 163.367
R2085 B.n660 B.n659 163.367
R2086 B.n659 B.n658 163.367
R2087 B.n658 B.n49 163.367
R2088 B.n654 B.n49 163.367
R2089 B.n654 B.n653 163.367
R2090 B.n653 B.n652 163.367
R2091 B.n652 B.n54 163.367
R2092 B.n648 B.n54 163.367
R2093 B.n648 B.n647 163.367
R2094 B.n647 B.n646 163.367
R2095 B.n646 B.n56 163.367
R2096 B.n641 B.n56 163.367
R2097 B.n641 B.n640 163.367
R2098 B.n640 B.n639 163.367
R2099 B.n639 B.n60 163.367
R2100 B.n635 B.n60 163.367
R2101 B.n635 B.n634 163.367
R2102 B.n634 B.n633 163.367
R2103 B.n633 B.n62 163.367
R2104 B.n629 B.n62 163.367
R2105 B.n629 B.n628 163.367
R2106 B.n628 B.n627 163.367
R2107 B.n627 B.n64 163.367
R2108 B.n623 B.n64 163.367
R2109 B.n623 B.n622 163.367
R2110 B.n622 B.n621 163.367
R2111 B.n621 B.n66 163.367
R2112 B.n617 B.n66 163.367
R2113 B.n617 B.n616 163.367
R2114 B.n616 B.n615 163.367
R2115 B.n615 B.n68 163.367
R2116 B.n611 B.n68 163.367
R2117 B.n611 B.n610 163.367
R2118 B.n610 B.n609 163.367
R2119 B.n609 B.n70 163.367
R2120 B.n605 B.n70 163.367
R2121 B.n605 B.n604 163.367
R2122 B.n604 B.n603 163.367
R2123 B.n603 B.n72 163.367
R2124 B.n599 B.n72 163.367
R2125 B.n599 B.n598 163.367
R2126 B.n598 B.n597 163.367
R2127 B.n597 B.n74 163.367
R2128 B.n593 B.n74 163.367
R2129 B.n593 B.n592 163.367
R2130 B.n592 B.n591 163.367
R2131 B.n591 B.n76 163.367
R2132 B.n587 B.n76 163.367
R2133 B.n587 B.n586 163.367
R2134 B.n586 B.n585 163.367
R2135 B.n585 B.n78 163.367
R2136 B.n581 B.n78 163.367
R2137 B.n581 B.n580 163.367
R2138 B.n580 B.n579 163.367
R2139 B.n579 B.n80 163.367
R2140 B.n575 B.n80 163.367
R2141 B.n575 B.n574 163.367
R2142 B.n574 B.n573 163.367
R2143 B.n573 B.n82 163.367
R2144 B.n569 B.n82 163.367
R2145 B.n569 B.n568 163.367
R2146 B.n568 B.n567 163.367
R2147 B.n567 B.n84 163.367
R2148 B.n563 B.n84 163.367
R2149 B.n563 B.n562 163.367
R2150 B.n562 B.n561 163.367
R2151 B.n561 B.n86 163.367
R2152 B.n557 B.n86 163.367
R2153 B.n557 B.n556 163.367
R2154 B.n556 B.n555 163.367
R2155 B.n555 B.n88 163.367
R2156 B.n361 B.n154 59.5399
R2157 B.n161 B.n160 59.5399
R2158 B.n52 B.n51 59.5399
R2159 B.n643 B.n58 59.5399
R2160 B.n154 B.n153 41.3096
R2161 B.n160 B.n159 41.3096
R2162 B.n51 B.n50 41.3096
R2163 B.n58 B.n57 41.3096
R2164 B.n747 B.n18 33.2493
R2165 B.n553 B.n552 33.2493
R2166 B.n452 B.n451 33.2493
R2167 B.n254 B.n191 33.2493
R2168 B B.n799 18.0485
R2169 B.n747 B.n746 10.6151
R2170 B.n746 B.n745 10.6151
R2171 B.n745 B.n20 10.6151
R2172 B.n741 B.n20 10.6151
R2173 B.n741 B.n740 10.6151
R2174 B.n740 B.n739 10.6151
R2175 B.n739 B.n22 10.6151
R2176 B.n735 B.n22 10.6151
R2177 B.n735 B.n734 10.6151
R2178 B.n734 B.n733 10.6151
R2179 B.n733 B.n24 10.6151
R2180 B.n729 B.n24 10.6151
R2181 B.n729 B.n728 10.6151
R2182 B.n728 B.n727 10.6151
R2183 B.n727 B.n26 10.6151
R2184 B.n723 B.n26 10.6151
R2185 B.n723 B.n722 10.6151
R2186 B.n722 B.n721 10.6151
R2187 B.n721 B.n28 10.6151
R2188 B.n717 B.n28 10.6151
R2189 B.n717 B.n716 10.6151
R2190 B.n716 B.n715 10.6151
R2191 B.n715 B.n30 10.6151
R2192 B.n711 B.n30 10.6151
R2193 B.n711 B.n710 10.6151
R2194 B.n710 B.n709 10.6151
R2195 B.n709 B.n32 10.6151
R2196 B.n705 B.n32 10.6151
R2197 B.n705 B.n704 10.6151
R2198 B.n704 B.n703 10.6151
R2199 B.n703 B.n34 10.6151
R2200 B.n699 B.n34 10.6151
R2201 B.n699 B.n698 10.6151
R2202 B.n698 B.n697 10.6151
R2203 B.n697 B.n36 10.6151
R2204 B.n693 B.n36 10.6151
R2205 B.n693 B.n692 10.6151
R2206 B.n692 B.n691 10.6151
R2207 B.n691 B.n38 10.6151
R2208 B.n687 B.n38 10.6151
R2209 B.n687 B.n686 10.6151
R2210 B.n686 B.n685 10.6151
R2211 B.n685 B.n40 10.6151
R2212 B.n681 B.n40 10.6151
R2213 B.n681 B.n680 10.6151
R2214 B.n680 B.n679 10.6151
R2215 B.n679 B.n42 10.6151
R2216 B.n675 B.n42 10.6151
R2217 B.n675 B.n674 10.6151
R2218 B.n674 B.n673 10.6151
R2219 B.n673 B.n44 10.6151
R2220 B.n669 B.n44 10.6151
R2221 B.n669 B.n668 10.6151
R2222 B.n668 B.n667 10.6151
R2223 B.n667 B.n46 10.6151
R2224 B.n663 B.n46 10.6151
R2225 B.n663 B.n662 10.6151
R2226 B.n662 B.n661 10.6151
R2227 B.n661 B.n48 10.6151
R2228 B.n657 B.n656 10.6151
R2229 B.n656 B.n655 10.6151
R2230 B.n655 B.n53 10.6151
R2231 B.n651 B.n53 10.6151
R2232 B.n651 B.n650 10.6151
R2233 B.n650 B.n649 10.6151
R2234 B.n649 B.n55 10.6151
R2235 B.n645 B.n55 10.6151
R2236 B.n645 B.n644 10.6151
R2237 B.n642 B.n59 10.6151
R2238 B.n638 B.n59 10.6151
R2239 B.n638 B.n637 10.6151
R2240 B.n637 B.n636 10.6151
R2241 B.n636 B.n61 10.6151
R2242 B.n632 B.n61 10.6151
R2243 B.n632 B.n631 10.6151
R2244 B.n631 B.n630 10.6151
R2245 B.n630 B.n63 10.6151
R2246 B.n626 B.n63 10.6151
R2247 B.n626 B.n625 10.6151
R2248 B.n625 B.n624 10.6151
R2249 B.n624 B.n65 10.6151
R2250 B.n620 B.n65 10.6151
R2251 B.n620 B.n619 10.6151
R2252 B.n619 B.n618 10.6151
R2253 B.n618 B.n67 10.6151
R2254 B.n614 B.n67 10.6151
R2255 B.n614 B.n613 10.6151
R2256 B.n613 B.n612 10.6151
R2257 B.n612 B.n69 10.6151
R2258 B.n608 B.n69 10.6151
R2259 B.n608 B.n607 10.6151
R2260 B.n607 B.n606 10.6151
R2261 B.n606 B.n71 10.6151
R2262 B.n602 B.n71 10.6151
R2263 B.n602 B.n601 10.6151
R2264 B.n601 B.n600 10.6151
R2265 B.n600 B.n73 10.6151
R2266 B.n596 B.n73 10.6151
R2267 B.n596 B.n595 10.6151
R2268 B.n595 B.n594 10.6151
R2269 B.n594 B.n75 10.6151
R2270 B.n590 B.n75 10.6151
R2271 B.n590 B.n589 10.6151
R2272 B.n589 B.n588 10.6151
R2273 B.n588 B.n77 10.6151
R2274 B.n584 B.n77 10.6151
R2275 B.n584 B.n583 10.6151
R2276 B.n583 B.n582 10.6151
R2277 B.n582 B.n79 10.6151
R2278 B.n578 B.n79 10.6151
R2279 B.n578 B.n577 10.6151
R2280 B.n577 B.n576 10.6151
R2281 B.n576 B.n81 10.6151
R2282 B.n572 B.n81 10.6151
R2283 B.n572 B.n571 10.6151
R2284 B.n571 B.n570 10.6151
R2285 B.n570 B.n83 10.6151
R2286 B.n566 B.n83 10.6151
R2287 B.n566 B.n565 10.6151
R2288 B.n565 B.n564 10.6151
R2289 B.n564 B.n85 10.6151
R2290 B.n560 B.n85 10.6151
R2291 B.n560 B.n559 10.6151
R2292 B.n559 B.n558 10.6151
R2293 B.n558 B.n87 10.6151
R2294 B.n554 B.n87 10.6151
R2295 B.n554 B.n553 10.6151
R2296 B.n452 B.n121 10.6151
R2297 B.n456 B.n121 10.6151
R2298 B.n457 B.n456 10.6151
R2299 B.n458 B.n457 10.6151
R2300 B.n458 B.n119 10.6151
R2301 B.n462 B.n119 10.6151
R2302 B.n463 B.n462 10.6151
R2303 B.n464 B.n463 10.6151
R2304 B.n464 B.n117 10.6151
R2305 B.n468 B.n117 10.6151
R2306 B.n469 B.n468 10.6151
R2307 B.n470 B.n469 10.6151
R2308 B.n470 B.n115 10.6151
R2309 B.n474 B.n115 10.6151
R2310 B.n475 B.n474 10.6151
R2311 B.n476 B.n475 10.6151
R2312 B.n476 B.n113 10.6151
R2313 B.n480 B.n113 10.6151
R2314 B.n481 B.n480 10.6151
R2315 B.n482 B.n481 10.6151
R2316 B.n482 B.n111 10.6151
R2317 B.n486 B.n111 10.6151
R2318 B.n487 B.n486 10.6151
R2319 B.n488 B.n487 10.6151
R2320 B.n488 B.n109 10.6151
R2321 B.n492 B.n109 10.6151
R2322 B.n493 B.n492 10.6151
R2323 B.n494 B.n493 10.6151
R2324 B.n494 B.n107 10.6151
R2325 B.n498 B.n107 10.6151
R2326 B.n499 B.n498 10.6151
R2327 B.n500 B.n499 10.6151
R2328 B.n500 B.n105 10.6151
R2329 B.n504 B.n105 10.6151
R2330 B.n505 B.n504 10.6151
R2331 B.n506 B.n505 10.6151
R2332 B.n506 B.n103 10.6151
R2333 B.n510 B.n103 10.6151
R2334 B.n511 B.n510 10.6151
R2335 B.n512 B.n511 10.6151
R2336 B.n512 B.n101 10.6151
R2337 B.n516 B.n101 10.6151
R2338 B.n517 B.n516 10.6151
R2339 B.n518 B.n517 10.6151
R2340 B.n518 B.n99 10.6151
R2341 B.n522 B.n99 10.6151
R2342 B.n523 B.n522 10.6151
R2343 B.n524 B.n523 10.6151
R2344 B.n524 B.n97 10.6151
R2345 B.n528 B.n97 10.6151
R2346 B.n529 B.n528 10.6151
R2347 B.n530 B.n529 10.6151
R2348 B.n530 B.n95 10.6151
R2349 B.n534 B.n95 10.6151
R2350 B.n535 B.n534 10.6151
R2351 B.n536 B.n535 10.6151
R2352 B.n536 B.n93 10.6151
R2353 B.n540 B.n93 10.6151
R2354 B.n541 B.n540 10.6151
R2355 B.n542 B.n541 10.6151
R2356 B.n542 B.n91 10.6151
R2357 B.n546 B.n91 10.6151
R2358 B.n547 B.n546 10.6151
R2359 B.n548 B.n547 10.6151
R2360 B.n548 B.n89 10.6151
R2361 B.n552 B.n89 10.6151
R2362 B.n258 B.n191 10.6151
R2363 B.n259 B.n258 10.6151
R2364 B.n260 B.n259 10.6151
R2365 B.n260 B.n189 10.6151
R2366 B.n264 B.n189 10.6151
R2367 B.n265 B.n264 10.6151
R2368 B.n266 B.n265 10.6151
R2369 B.n266 B.n187 10.6151
R2370 B.n270 B.n187 10.6151
R2371 B.n271 B.n270 10.6151
R2372 B.n272 B.n271 10.6151
R2373 B.n272 B.n185 10.6151
R2374 B.n276 B.n185 10.6151
R2375 B.n277 B.n276 10.6151
R2376 B.n278 B.n277 10.6151
R2377 B.n278 B.n183 10.6151
R2378 B.n282 B.n183 10.6151
R2379 B.n283 B.n282 10.6151
R2380 B.n284 B.n283 10.6151
R2381 B.n284 B.n181 10.6151
R2382 B.n288 B.n181 10.6151
R2383 B.n289 B.n288 10.6151
R2384 B.n290 B.n289 10.6151
R2385 B.n290 B.n179 10.6151
R2386 B.n294 B.n179 10.6151
R2387 B.n295 B.n294 10.6151
R2388 B.n296 B.n295 10.6151
R2389 B.n296 B.n177 10.6151
R2390 B.n300 B.n177 10.6151
R2391 B.n301 B.n300 10.6151
R2392 B.n302 B.n301 10.6151
R2393 B.n302 B.n175 10.6151
R2394 B.n306 B.n175 10.6151
R2395 B.n307 B.n306 10.6151
R2396 B.n308 B.n307 10.6151
R2397 B.n308 B.n173 10.6151
R2398 B.n312 B.n173 10.6151
R2399 B.n313 B.n312 10.6151
R2400 B.n314 B.n313 10.6151
R2401 B.n314 B.n171 10.6151
R2402 B.n318 B.n171 10.6151
R2403 B.n319 B.n318 10.6151
R2404 B.n320 B.n319 10.6151
R2405 B.n320 B.n169 10.6151
R2406 B.n324 B.n169 10.6151
R2407 B.n325 B.n324 10.6151
R2408 B.n326 B.n325 10.6151
R2409 B.n326 B.n167 10.6151
R2410 B.n330 B.n167 10.6151
R2411 B.n331 B.n330 10.6151
R2412 B.n332 B.n331 10.6151
R2413 B.n332 B.n165 10.6151
R2414 B.n336 B.n165 10.6151
R2415 B.n337 B.n336 10.6151
R2416 B.n338 B.n337 10.6151
R2417 B.n338 B.n163 10.6151
R2418 B.n342 B.n163 10.6151
R2419 B.n343 B.n342 10.6151
R2420 B.n344 B.n343 10.6151
R2421 B.n348 B.n347 10.6151
R2422 B.n349 B.n348 10.6151
R2423 B.n349 B.n157 10.6151
R2424 B.n353 B.n157 10.6151
R2425 B.n354 B.n353 10.6151
R2426 B.n355 B.n354 10.6151
R2427 B.n355 B.n155 10.6151
R2428 B.n359 B.n155 10.6151
R2429 B.n360 B.n359 10.6151
R2430 B.n362 B.n151 10.6151
R2431 B.n366 B.n151 10.6151
R2432 B.n367 B.n366 10.6151
R2433 B.n368 B.n367 10.6151
R2434 B.n368 B.n149 10.6151
R2435 B.n372 B.n149 10.6151
R2436 B.n373 B.n372 10.6151
R2437 B.n374 B.n373 10.6151
R2438 B.n374 B.n147 10.6151
R2439 B.n378 B.n147 10.6151
R2440 B.n379 B.n378 10.6151
R2441 B.n380 B.n379 10.6151
R2442 B.n380 B.n145 10.6151
R2443 B.n384 B.n145 10.6151
R2444 B.n385 B.n384 10.6151
R2445 B.n386 B.n385 10.6151
R2446 B.n386 B.n143 10.6151
R2447 B.n390 B.n143 10.6151
R2448 B.n391 B.n390 10.6151
R2449 B.n392 B.n391 10.6151
R2450 B.n392 B.n141 10.6151
R2451 B.n396 B.n141 10.6151
R2452 B.n397 B.n396 10.6151
R2453 B.n398 B.n397 10.6151
R2454 B.n398 B.n139 10.6151
R2455 B.n402 B.n139 10.6151
R2456 B.n403 B.n402 10.6151
R2457 B.n404 B.n403 10.6151
R2458 B.n404 B.n137 10.6151
R2459 B.n408 B.n137 10.6151
R2460 B.n409 B.n408 10.6151
R2461 B.n410 B.n409 10.6151
R2462 B.n410 B.n135 10.6151
R2463 B.n414 B.n135 10.6151
R2464 B.n415 B.n414 10.6151
R2465 B.n416 B.n415 10.6151
R2466 B.n416 B.n133 10.6151
R2467 B.n420 B.n133 10.6151
R2468 B.n421 B.n420 10.6151
R2469 B.n422 B.n421 10.6151
R2470 B.n422 B.n131 10.6151
R2471 B.n426 B.n131 10.6151
R2472 B.n427 B.n426 10.6151
R2473 B.n428 B.n427 10.6151
R2474 B.n428 B.n129 10.6151
R2475 B.n432 B.n129 10.6151
R2476 B.n433 B.n432 10.6151
R2477 B.n434 B.n433 10.6151
R2478 B.n434 B.n127 10.6151
R2479 B.n438 B.n127 10.6151
R2480 B.n439 B.n438 10.6151
R2481 B.n440 B.n439 10.6151
R2482 B.n440 B.n125 10.6151
R2483 B.n444 B.n125 10.6151
R2484 B.n445 B.n444 10.6151
R2485 B.n446 B.n445 10.6151
R2486 B.n446 B.n123 10.6151
R2487 B.n450 B.n123 10.6151
R2488 B.n451 B.n450 10.6151
R2489 B.n254 B.n253 10.6151
R2490 B.n253 B.n252 10.6151
R2491 B.n252 B.n193 10.6151
R2492 B.n248 B.n193 10.6151
R2493 B.n248 B.n247 10.6151
R2494 B.n247 B.n246 10.6151
R2495 B.n246 B.n195 10.6151
R2496 B.n242 B.n195 10.6151
R2497 B.n242 B.n241 10.6151
R2498 B.n241 B.n240 10.6151
R2499 B.n240 B.n197 10.6151
R2500 B.n236 B.n197 10.6151
R2501 B.n236 B.n235 10.6151
R2502 B.n235 B.n234 10.6151
R2503 B.n234 B.n199 10.6151
R2504 B.n230 B.n199 10.6151
R2505 B.n230 B.n229 10.6151
R2506 B.n229 B.n228 10.6151
R2507 B.n228 B.n201 10.6151
R2508 B.n224 B.n201 10.6151
R2509 B.n224 B.n223 10.6151
R2510 B.n223 B.n222 10.6151
R2511 B.n222 B.n203 10.6151
R2512 B.n218 B.n203 10.6151
R2513 B.n218 B.n217 10.6151
R2514 B.n217 B.n216 10.6151
R2515 B.n216 B.n205 10.6151
R2516 B.n212 B.n205 10.6151
R2517 B.n212 B.n211 10.6151
R2518 B.n211 B.n210 10.6151
R2519 B.n210 B.n207 10.6151
R2520 B.n207 B.n0 10.6151
R2521 B.n795 B.n1 10.6151
R2522 B.n795 B.n794 10.6151
R2523 B.n794 B.n793 10.6151
R2524 B.n793 B.n4 10.6151
R2525 B.n789 B.n4 10.6151
R2526 B.n789 B.n788 10.6151
R2527 B.n788 B.n787 10.6151
R2528 B.n787 B.n6 10.6151
R2529 B.n783 B.n6 10.6151
R2530 B.n783 B.n782 10.6151
R2531 B.n782 B.n781 10.6151
R2532 B.n781 B.n8 10.6151
R2533 B.n777 B.n8 10.6151
R2534 B.n777 B.n776 10.6151
R2535 B.n776 B.n775 10.6151
R2536 B.n775 B.n10 10.6151
R2537 B.n771 B.n10 10.6151
R2538 B.n771 B.n770 10.6151
R2539 B.n770 B.n769 10.6151
R2540 B.n769 B.n12 10.6151
R2541 B.n765 B.n12 10.6151
R2542 B.n765 B.n764 10.6151
R2543 B.n764 B.n763 10.6151
R2544 B.n763 B.n14 10.6151
R2545 B.n759 B.n14 10.6151
R2546 B.n759 B.n758 10.6151
R2547 B.n758 B.n757 10.6151
R2548 B.n757 B.n16 10.6151
R2549 B.n753 B.n16 10.6151
R2550 B.n753 B.n752 10.6151
R2551 B.n752 B.n751 10.6151
R2552 B.n751 B.n18 10.6151
R2553 B.n52 B.n48 9.36635
R2554 B.n643 B.n642 9.36635
R2555 B.n344 B.n161 9.36635
R2556 B.n362 B.n361 9.36635
R2557 B.n799 B.n0 2.81026
R2558 B.n799 B.n1 2.81026
R2559 B.n657 B.n52 1.24928
R2560 B.n644 B.n643 1.24928
R2561 B.n347 B.n161 1.24928
R2562 B.n361 B.n360 1.24928
C0 VN VDD1 0.14953f
C1 w_n2674_n4626# VDD2 2.59856f
C2 VP VTAIL 8.97348f
C3 w_n2674_n4626# VDD1 2.53908f
C4 VP VDD2 0.39109f
C5 VDD2 VTAIL 10.490499f
C6 B VN 1.07192f
C7 VP VDD1 9.48183f
C8 VTAIL VDD1 10.4482f
C9 w_n2674_n4626# B 10.334599f
C10 VDD2 VDD1 1.1209f
C11 B VP 1.64137f
C12 B VTAIL 4.65411f
C13 B VDD2 2.41876f
C14 w_n2674_n4626# VN 4.98529f
C15 B VDD1 2.36382f
C16 VP VN 7.31151f
C17 VN VTAIL 8.95897f
C18 w_n2674_n4626# VP 5.32877f
C19 VN VDD2 9.24521f
C20 w_n2674_n4626# VTAIL 3.82459f
C21 VDD2 VSUBS 1.869946f
C22 VDD1 VSUBS 1.715343f
C23 VTAIL VSUBS 1.271041f
C24 VN VSUBS 5.44107f
C25 VP VSUBS 2.534878f
C26 B VSUBS 4.378794f
C27 w_n2674_n4626# VSUBS 0.151231p
C28 B.n0 VSUBS 0.004898f
C29 B.n1 VSUBS 0.004898f
C30 B.n2 VSUBS 0.007746f
C31 B.n3 VSUBS 0.007746f
C32 B.n4 VSUBS 0.007746f
C33 B.n5 VSUBS 0.007746f
C34 B.n6 VSUBS 0.007746f
C35 B.n7 VSUBS 0.007746f
C36 B.n8 VSUBS 0.007746f
C37 B.n9 VSUBS 0.007746f
C38 B.n10 VSUBS 0.007746f
C39 B.n11 VSUBS 0.007746f
C40 B.n12 VSUBS 0.007746f
C41 B.n13 VSUBS 0.007746f
C42 B.n14 VSUBS 0.007746f
C43 B.n15 VSUBS 0.007746f
C44 B.n16 VSUBS 0.007746f
C45 B.n17 VSUBS 0.007746f
C46 B.n18 VSUBS 0.017714f
C47 B.n19 VSUBS 0.007746f
C48 B.n20 VSUBS 0.007746f
C49 B.n21 VSUBS 0.007746f
C50 B.n22 VSUBS 0.007746f
C51 B.n23 VSUBS 0.007746f
C52 B.n24 VSUBS 0.007746f
C53 B.n25 VSUBS 0.007746f
C54 B.n26 VSUBS 0.007746f
C55 B.n27 VSUBS 0.007746f
C56 B.n28 VSUBS 0.007746f
C57 B.n29 VSUBS 0.007746f
C58 B.n30 VSUBS 0.007746f
C59 B.n31 VSUBS 0.007746f
C60 B.n32 VSUBS 0.007746f
C61 B.n33 VSUBS 0.007746f
C62 B.n34 VSUBS 0.007746f
C63 B.n35 VSUBS 0.007746f
C64 B.n36 VSUBS 0.007746f
C65 B.n37 VSUBS 0.007746f
C66 B.n38 VSUBS 0.007746f
C67 B.n39 VSUBS 0.007746f
C68 B.n40 VSUBS 0.007746f
C69 B.n41 VSUBS 0.007746f
C70 B.n42 VSUBS 0.007746f
C71 B.n43 VSUBS 0.007746f
C72 B.n44 VSUBS 0.007746f
C73 B.n45 VSUBS 0.007746f
C74 B.n46 VSUBS 0.007746f
C75 B.n47 VSUBS 0.007746f
C76 B.n48 VSUBS 0.00729f
C77 B.n49 VSUBS 0.007746f
C78 B.t5 VSUBS 0.396408f
C79 B.t4 VSUBS 0.423879f
C80 B.t3 VSUBS 1.56944f
C81 B.n50 VSUBS 0.610689f
C82 B.n51 VSUBS 0.363743f
C83 B.n52 VSUBS 0.017946f
C84 B.n53 VSUBS 0.007746f
C85 B.n54 VSUBS 0.007746f
C86 B.n55 VSUBS 0.007746f
C87 B.n56 VSUBS 0.007746f
C88 B.t2 VSUBS 0.396412f
C89 B.t1 VSUBS 0.423882f
C90 B.t0 VSUBS 1.56944f
C91 B.n57 VSUBS 0.610685f
C92 B.n58 VSUBS 0.363739f
C93 B.n59 VSUBS 0.007746f
C94 B.n60 VSUBS 0.007746f
C95 B.n61 VSUBS 0.007746f
C96 B.n62 VSUBS 0.007746f
C97 B.n63 VSUBS 0.007746f
C98 B.n64 VSUBS 0.007746f
C99 B.n65 VSUBS 0.007746f
C100 B.n66 VSUBS 0.007746f
C101 B.n67 VSUBS 0.007746f
C102 B.n68 VSUBS 0.007746f
C103 B.n69 VSUBS 0.007746f
C104 B.n70 VSUBS 0.007746f
C105 B.n71 VSUBS 0.007746f
C106 B.n72 VSUBS 0.007746f
C107 B.n73 VSUBS 0.007746f
C108 B.n74 VSUBS 0.007746f
C109 B.n75 VSUBS 0.007746f
C110 B.n76 VSUBS 0.007746f
C111 B.n77 VSUBS 0.007746f
C112 B.n78 VSUBS 0.007746f
C113 B.n79 VSUBS 0.007746f
C114 B.n80 VSUBS 0.007746f
C115 B.n81 VSUBS 0.007746f
C116 B.n82 VSUBS 0.007746f
C117 B.n83 VSUBS 0.007746f
C118 B.n84 VSUBS 0.007746f
C119 B.n85 VSUBS 0.007746f
C120 B.n86 VSUBS 0.007746f
C121 B.n87 VSUBS 0.007746f
C122 B.n88 VSUBS 0.018964f
C123 B.n89 VSUBS 0.007746f
C124 B.n90 VSUBS 0.007746f
C125 B.n91 VSUBS 0.007746f
C126 B.n92 VSUBS 0.007746f
C127 B.n93 VSUBS 0.007746f
C128 B.n94 VSUBS 0.007746f
C129 B.n95 VSUBS 0.007746f
C130 B.n96 VSUBS 0.007746f
C131 B.n97 VSUBS 0.007746f
C132 B.n98 VSUBS 0.007746f
C133 B.n99 VSUBS 0.007746f
C134 B.n100 VSUBS 0.007746f
C135 B.n101 VSUBS 0.007746f
C136 B.n102 VSUBS 0.007746f
C137 B.n103 VSUBS 0.007746f
C138 B.n104 VSUBS 0.007746f
C139 B.n105 VSUBS 0.007746f
C140 B.n106 VSUBS 0.007746f
C141 B.n107 VSUBS 0.007746f
C142 B.n108 VSUBS 0.007746f
C143 B.n109 VSUBS 0.007746f
C144 B.n110 VSUBS 0.007746f
C145 B.n111 VSUBS 0.007746f
C146 B.n112 VSUBS 0.007746f
C147 B.n113 VSUBS 0.007746f
C148 B.n114 VSUBS 0.007746f
C149 B.n115 VSUBS 0.007746f
C150 B.n116 VSUBS 0.007746f
C151 B.n117 VSUBS 0.007746f
C152 B.n118 VSUBS 0.007746f
C153 B.n119 VSUBS 0.007746f
C154 B.n120 VSUBS 0.007746f
C155 B.n121 VSUBS 0.007746f
C156 B.n122 VSUBS 0.018964f
C157 B.n123 VSUBS 0.007746f
C158 B.n124 VSUBS 0.007746f
C159 B.n125 VSUBS 0.007746f
C160 B.n126 VSUBS 0.007746f
C161 B.n127 VSUBS 0.007746f
C162 B.n128 VSUBS 0.007746f
C163 B.n129 VSUBS 0.007746f
C164 B.n130 VSUBS 0.007746f
C165 B.n131 VSUBS 0.007746f
C166 B.n132 VSUBS 0.007746f
C167 B.n133 VSUBS 0.007746f
C168 B.n134 VSUBS 0.007746f
C169 B.n135 VSUBS 0.007746f
C170 B.n136 VSUBS 0.007746f
C171 B.n137 VSUBS 0.007746f
C172 B.n138 VSUBS 0.007746f
C173 B.n139 VSUBS 0.007746f
C174 B.n140 VSUBS 0.007746f
C175 B.n141 VSUBS 0.007746f
C176 B.n142 VSUBS 0.007746f
C177 B.n143 VSUBS 0.007746f
C178 B.n144 VSUBS 0.007746f
C179 B.n145 VSUBS 0.007746f
C180 B.n146 VSUBS 0.007746f
C181 B.n147 VSUBS 0.007746f
C182 B.n148 VSUBS 0.007746f
C183 B.n149 VSUBS 0.007746f
C184 B.n150 VSUBS 0.007746f
C185 B.n151 VSUBS 0.007746f
C186 B.n152 VSUBS 0.007746f
C187 B.t10 VSUBS 0.396412f
C188 B.t11 VSUBS 0.423882f
C189 B.t9 VSUBS 1.56944f
C190 B.n153 VSUBS 0.610685f
C191 B.n154 VSUBS 0.363739f
C192 B.n155 VSUBS 0.007746f
C193 B.n156 VSUBS 0.007746f
C194 B.n157 VSUBS 0.007746f
C195 B.n158 VSUBS 0.007746f
C196 B.t7 VSUBS 0.396408f
C197 B.t8 VSUBS 0.423879f
C198 B.t6 VSUBS 1.56944f
C199 B.n159 VSUBS 0.610689f
C200 B.n160 VSUBS 0.363743f
C201 B.n161 VSUBS 0.017946f
C202 B.n162 VSUBS 0.007746f
C203 B.n163 VSUBS 0.007746f
C204 B.n164 VSUBS 0.007746f
C205 B.n165 VSUBS 0.007746f
C206 B.n166 VSUBS 0.007746f
C207 B.n167 VSUBS 0.007746f
C208 B.n168 VSUBS 0.007746f
C209 B.n169 VSUBS 0.007746f
C210 B.n170 VSUBS 0.007746f
C211 B.n171 VSUBS 0.007746f
C212 B.n172 VSUBS 0.007746f
C213 B.n173 VSUBS 0.007746f
C214 B.n174 VSUBS 0.007746f
C215 B.n175 VSUBS 0.007746f
C216 B.n176 VSUBS 0.007746f
C217 B.n177 VSUBS 0.007746f
C218 B.n178 VSUBS 0.007746f
C219 B.n179 VSUBS 0.007746f
C220 B.n180 VSUBS 0.007746f
C221 B.n181 VSUBS 0.007746f
C222 B.n182 VSUBS 0.007746f
C223 B.n183 VSUBS 0.007746f
C224 B.n184 VSUBS 0.007746f
C225 B.n185 VSUBS 0.007746f
C226 B.n186 VSUBS 0.007746f
C227 B.n187 VSUBS 0.007746f
C228 B.n188 VSUBS 0.007746f
C229 B.n189 VSUBS 0.007746f
C230 B.n190 VSUBS 0.007746f
C231 B.n191 VSUBS 0.018964f
C232 B.n192 VSUBS 0.007746f
C233 B.n193 VSUBS 0.007746f
C234 B.n194 VSUBS 0.007746f
C235 B.n195 VSUBS 0.007746f
C236 B.n196 VSUBS 0.007746f
C237 B.n197 VSUBS 0.007746f
C238 B.n198 VSUBS 0.007746f
C239 B.n199 VSUBS 0.007746f
C240 B.n200 VSUBS 0.007746f
C241 B.n201 VSUBS 0.007746f
C242 B.n202 VSUBS 0.007746f
C243 B.n203 VSUBS 0.007746f
C244 B.n204 VSUBS 0.007746f
C245 B.n205 VSUBS 0.007746f
C246 B.n206 VSUBS 0.007746f
C247 B.n207 VSUBS 0.007746f
C248 B.n208 VSUBS 0.007746f
C249 B.n209 VSUBS 0.007746f
C250 B.n210 VSUBS 0.007746f
C251 B.n211 VSUBS 0.007746f
C252 B.n212 VSUBS 0.007746f
C253 B.n213 VSUBS 0.007746f
C254 B.n214 VSUBS 0.007746f
C255 B.n215 VSUBS 0.007746f
C256 B.n216 VSUBS 0.007746f
C257 B.n217 VSUBS 0.007746f
C258 B.n218 VSUBS 0.007746f
C259 B.n219 VSUBS 0.007746f
C260 B.n220 VSUBS 0.007746f
C261 B.n221 VSUBS 0.007746f
C262 B.n222 VSUBS 0.007746f
C263 B.n223 VSUBS 0.007746f
C264 B.n224 VSUBS 0.007746f
C265 B.n225 VSUBS 0.007746f
C266 B.n226 VSUBS 0.007746f
C267 B.n227 VSUBS 0.007746f
C268 B.n228 VSUBS 0.007746f
C269 B.n229 VSUBS 0.007746f
C270 B.n230 VSUBS 0.007746f
C271 B.n231 VSUBS 0.007746f
C272 B.n232 VSUBS 0.007746f
C273 B.n233 VSUBS 0.007746f
C274 B.n234 VSUBS 0.007746f
C275 B.n235 VSUBS 0.007746f
C276 B.n236 VSUBS 0.007746f
C277 B.n237 VSUBS 0.007746f
C278 B.n238 VSUBS 0.007746f
C279 B.n239 VSUBS 0.007746f
C280 B.n240 VSUBS 0.007746f
C281 B.n241 VSUBS 0.007746f
C282 B.n242 VSUBS 0.007746f
C283 B.n243 VSUBS 0.007746f
C284 B.n244 VSUBS 0.007746f
C285 B.n245 VSUBS 0.007746f
C286 B.n246 VSUBS 0.007746f
C287 B.n247 VSUBS 0.007746f
C288 B.n248 VSUBS 0.007746f
C289 B.n249 VSUBS 0.007746f
C290 B.n250 VSUBS 0.007746f
C291 B.n251 VSUBS 0.007746f
C292 B.n252 VSUBS 0.007746f
C293 B.n253 VSUBS 0.007746f
C294 B.n254 VSUBS 0.017714f
C295 B.n255 VSUBS 0.017714f
C296 B.n256 VSUBS 0.018964f
C297 B.n257 VSUBS 0.007746f
C298 B.n258 VSUBS 0.007746f
C299 B.n259 VSUBS 0.007746f
C300 B.n260 VSUBS 0.007746f
C301 B.n261 VSUBS 0.007746f
C302 B.n262 VSUBS 0.007746f
C303 B.n263 VSUBS 0.007746f
C304 B.n264 VSUBS 0.007746f
C305 B.n265 VSUBS 0.007746f
C306 B.n266 VSUBS 0.007746f
C307 B.n267 VSUBS 0.007746f
C308 B.n268 VSUBS 0.007746f
C309 B.n269 VSUBS 0.007746f
C310 B.n270 VSUBS 0.007746f
C311 B.n271 VSUBS 0.007746f
C312 B.n272 VSUBS 0.007746f
C313 B.n273 VSUBS 0.007746f
C314 B.n274 VSUBS 0.007746f
C315 B.n275 VSUBS 0.007746f
C316 B.n276 VSUBS 0.007746f
C317 B.n277 VSUBS 0.007746f
C318 B.n278 VSUBS 0.007746f
C319 B.n279 VSUBS 0.007746f
C320 B.n280 VSUBS 0.007746f
C321 B.n281 VSUBS 0.007746f
C322 B.n282 VSUBS 0.007746f
C323 B.n283 VSUBS 0.007746f
C324 B.n284 VSUBS 0.007746f
C325 B.n285 VSUBS 0.007746f
C326 B.n286 VSUBS 0.007746f
C327 B.n287 VSUBS 0.007746f
C328 B.n288 VSUBS 0.007746f
C329 B.n289 VSUBS 0.007746f
C330 B.n290 VSUBS 0.007746f
C331 B.n291 VSUBS 0.007746f
C332 B.n292 VSUBS 0.007746f
C333 B.n293 VSUBS 0.007746f
C334 B.n294 VSUBS 0.007746f
C335 B.n295 VSUBS 0.007746f
C336 B.n296 VSUBS 0.007746f
C337 B.n297 VSUBS 0.007746f
C338 B.n298 VSUBS 0.007746f
C339 B.n299 VSUBS 0.007746f
C340 B.n300 VSUBS 0.007746f
C341 B.n301 VSUBS 0.007746f
C342 B.n302 VSUBS 0.007746f
C343 B.n303 VSUBS 0.007746f
C344 B.n304 VSUBS 0.007746f
C345 B.n305 VSUBS 0.007746f
C346 B.n306 VSUBS 0.007746f
C347 B.n307 VSUBS 0.007746f
C348 B.n308 VSUBS 0.007746f
C349 B.n309 VSUBS 0.007746f
C350 B.n310 VSUBS 0.007746f
C351 B.n311 VSUBS 0.007746f
C352 B.n312 VSUBS 0.007746f
C353 B.n313 VSUBS 0.007746f
C354 B.n314 VSUBS 0.007746f
C355 B.n315 VSUBS 0.007746f
C356 B.n316 VSUBS 0.007746f
C357 B.n317 VSUBS 0.007746f
C358 B.n318 VSUBS 0.007746f
C359 B.n319 VSUBS 0.007746f
C360 B.n320 VSUBS 0.007746f
C361 B.n321 VSUBS 0.007746f
C362 B.n322 VSUBS 0.007746f
C363 B.n323 VSUBS 0.007746f
C364 B.n324 VSUBS 0.007746f
C365 B.n325 VSUBS 0.007746f
C366 B.n326 VSUBS 0.007746f
C367 B.n327 VSUBS 0.007746f
C368 B.n328 VSUBS 0.007746f
C369 B.n329 VSUBS 0.007746f
C370 B.n330 VSUBS 0.007746f
C371 B.n331 VSUBS 0.007746f
C372 B.n332 VSUBS 0.007746f
C373 B.n333 VSUBS 0.007746f
C374 B.n334 VSUBS 0.007746f
C375 B.n335 VSUBS 0.007746f
C376 B.n336 VSUBS 0.007746f
C377 B.n337 VSUBS 0.007746f
C378 B.n338 VSUBS 0.007746f
C379 B.n339 VSUBS 0.007746f
C380 B.n340 VSUBS 0.007746f
C381 B.n341 VSUBS 0.007746f
C382 B.n342 VSUBS 0.007746f
C383 B.n343 VSUBS 0.007746f
C384 B.n344 VSUBS 0.00729f
C385 B.n345 VSUBS 0.007746f
C386 B.n346 VSUBS 0.007746f
C387 B.n347 VSUBS 0.004329f
C388 B.n348 VSUBS 0.007746f
C389 B.n349 VSUBS 0.007746f
C390 B.n350 VSUBS 0.007746f
C391 B.n351 VSUBS 0.007746f
C392 B.n352 VSUBS 0.007746f
C393 B.n353 VSUBS 0.007746f
C394 B.n354 VSUBS 0.007746f
C395 B.n355 VSUBS 0.007746f
C396 B.n356 VSUBS 0.007746f
C397 B.n357 VSUBS 0.007746f
C398 B.n358 VSUBS 0.007746f
C399 B.n359 VSUBS 0.007746f
C400 B.n360 VSUBS 0.004329f
C401 B.n361 VSUBS 0.017946f
C402 B.n362 VSUBS 0.00729f
C403 B.n363 VSUBS 0.007746f
C404 B.n364 VSUBS 0.007746f
C405 B.n365 VSUBS 0.007746f
C406 B.n366 VSUBS 0.007746f
C407 B.n367 VSUBS 0.007746f
C408 B.n368 VSUBS 0.007746f
C409 B.n369 VSUBS 0.007746f
C410 B.n370 VSUBS 0.007746f
C411 B.n371 VSUBS 0.007746f
C412 B.n372 VSUBS 0.007746f
C413 B.n373 VSUBS 0.007746f
C414 B.n374 VSUBS 0.007746f
C415 B.n375 VSUBS 0.007746f
C416 B.n376 VSUBS 0.007746f
C417 B.n377 VSUBS 0.007746f
C418 B.n378 VSUBS 0.007746f
C419 B.n379 VSUBS 0.007746f
C420 B.n380 VSUBS 0.007746f
C421 B.n381 VSUBS 0.007746f
C422 B.n382 VSUBS 0.007746f
C423 B.n383 VSUBS 0.007746f
C424 B.n384 VSUBS 0.007746f
C425 B.n385 VSUBS 0.007746f
C426 B.n386 VSUBS 0.007746f
C427 B.n387 VSUBS 0.007746f
C428 B.n388 VSUBS 0.007746f
C429 B.n389 VSUBS 0.007746f
C430 B.n390 VSUBS 0.007746f
C431 B.n391 VSUBS 0.007746f
C432 B.n392 VSUBS 0.007746f
C433 B.n393 VSUBS 0.007746f
C434 B.n394 VSUBS 0.007746f
C435 B.n395 VSUBS 0.007746f
C436 B.n396 VSUBS 0.007746f
C437 B.n397 VSUBS 0.007746f
C438 B.n398 VSUBS 0.007746f
C439 B.n399 VSUBS 0.007746f
C440 B.n400 VSUBS 0.007746f
C441 B.n401 VSUBS 0.007746f
C442 B.n402 VSUBS 0.007746f
C443 B.n403 VSUBS 0.007746f
C444 B.n404 VSUBS 0.007746f
C445 B.n405 VSUBS 0.007746f
C446 B.n406 VSUBS 0.007746f
C447 B.n407 VSUBS 0.007746f
C448 B.n408 VSUBS 0.007746f
C449 B.n409 VSUBS 0.007746f
C450 B.n410 VSUBS 0.007746f
C451 B.n411 VSUBS 0.007746f
C452 B.n412 VSUBS 0.007746f
C453 B.n413 VSUBS 0.007746f
C454 B.n414 VSUBS 0.007746f
C455 B.n415 VSUBS 0.007746f
C456 B.n416 VSUBS 0.007746f
C457 B.n417 VSUBS 0.007746f
C458 B.n418 VSUBS 0.007746f
C459 B.n419 VSUBS 0.007746f
C460 B.n420 VSUBS 0.007746f
C461 B.n421 VSUBS 0.007746f
C462 B.n422 VSUBS 0.007746f
C463 B.n423 VSUBS 0.007746f
C464 B.n424 VSUBS 0.007746f
C465 B.n425 VSUBS 0.007746f
C466 B.n426 VSUBS 0.007746f
C467 B.n427 VSUBS 0.007746f
C468 B.n428 VSUBS 0.007746f
C469 B.n429 VSUBS 0.007746f
C470 B.n430 VSUBS 0.007746f
C471 B.n431 VSUBS 0.007746f
C472 B.n432 VSUBS 0.007746f
C473 B.n433 VSUBS 0.007746f
C474 B.n434 VSUBS 0.007746f
C475 B.n435 VSUBS 0.007746f
C476 B.n436 VSUBS 0.007746f
C477 B.n437 VSUBS 0.007746f
C478 B.n438 VSUBS 0.007746f
C479 B.n439 VSUBS 0.007746f
C480 B.n440 VSUBS 0.007746f
C481 B.n441 VSUBS 0.007746f
C482 B.n442 VSUBS 0.007746f
C483 B.n443 VSUBS 0.007746f
C484 B.n444 VSUBS 0.007746f
C485 B.n445 VSUBS 0.007746f
C486 B.n446 VSUBS 0.007746f
C487 B.n447 VSUBS 0.007746f
C488 B.n448 VSUBS 0.007746f
C489 B.n449 VSUBS 0.007746f
C490 B.n450 VSUBS 0.007746f
C491 B.n451 VSUBS 0.018964f
C492 B.n452 VSUBS 0.017714f
C493 B.n453 VSUBS 0.017714f
C494 B.n454 VSUBS 0.007746f
C495 B.n455 VSUBS 0.007746f
C496 B.n456 VSUBS 0.007746f
C497 B.n457 VSUBS 0.007746f
C498 B.n458 VSUBS 0.007746f
C499 B.n459 VSUBS 0.007746f
C500 B.n460 VSUBS 0.007746f
C501 B.n461 VSUBS 0.007746f
C502 B.n462 VSUBS 0.007746f
C503 B.n463 VSUBS 0.007746f
C504 B.n464 VSUBS 0.007746f
C505 B.n465 VSUBS 0.007746f
C506 B.n466 VSUBS 0.007746f
C507 B.n467 VSUBS 0.007746f
C508 B.n468 VSUBS 0.007746f
C509 B.n469 VSUBS 0.007746f
C510 B.n470 VSUBS 0.007746f
C511 B.n471 VSUBS 0.007746f
C512 B.n472 VSUBS 0.007746f
C513 B.n473 VSUBS 0.007746f
C514 B.n474 VSUBS 0.007746f
C515 B.n475 VSUBS 0.007746f
C516 B.n476 VSUBS 0.007746f
C517 B.n477 VSUBS 0.007746f
C518 B.n478 VSUBS 0.007746f
C519 B.n479 VSUBS 0.007746f
C520 B.n480 VSUBS 0.007746f
C521 B.n481 VSUBS 0.007746f
C522 B.n482 VSUBS 0.007746f
C523 B.n483 VSUBS 0.007746f
C524 B.n484 VSUBS 0.007746f
C525 B.n485 VSUBS 0.007746f
C526 B.n486 VSUBS 0.007746f
C527 B.n487 VSUBS 0.007746f
C528 B.n488 VSUBS 0.007746f
C529 B.n489 VSUBS 0.007746f
C530 B.n490 VSUBS 0.007746f
C531 B.n491 VSUBS 0.007746f
C532 B.n492 VSUBS 0.007746f
C533 B.n493 VSUBS 0.007746f
C534 B.n494 VSUBS 0.007746f
C535 B.n495 VSUBS 0.007746f
C536 B.n496 VSUBS 0.007746f
C537 B.n497 VSUBS 0.007746f
C538 B.n498 VSUBS 0.007746f
C539 B.n499 VSUBS 0.007746f
C540 B.n500 VSUBS 0.007746f
C541 B.n501 VSUBS 0.007746f
C542 B.n502 VSUBS 0.007746f
C543 B.n503 VSUBS 0.007746f
C544 B.n504 VSUBS 0.007746f
C545 B.n505 VSUBS 0.007746f
C546 B.n506 VSUBS 0.007746f
C547 B.n507 VSUBS 0.007746f
C548 B.n508 VSUBS 0.007746f
C549 B.n509 VSUBS 0.007746f
C550 B.n510 VSUBS 0.007746f
C551 B.n511 VSUBS 0.007746f
C552 B.n512 VSUBS 0.007746f
C553 B.n513 VSUBS 0.007746f
C554 B.n514 VSUBS 0.007746f
C555 B.n515 VSUBS 0.007746f
C556 B.n516 VSUBS 0.007746f
C557 B.n517 VSUBS 0.007746f
C558 B.n518 VSUBS 0.007746f
C559 B.n519 VSUBS 0.007746f
C560 B.n520 VSUBS 0.007746f
C561 B.n521 VSUBS 0.007746f
C562 B.n522 VSUBS 0.007746f
C563 B.n523 VSUBS 0.007746f
C564 B.n524 VSUBS 0.007746f
C565 B.n525 VSUBS 0.007746f
C566 B.n526 VSUBS 0.007746f
C567 B.n527 VSUBS 0.007746f
C568 B.n528 VSUBS 0.007746f
C569 B.n529 VSUBS 0.007746f
C570 B.n530 VSUBS 0.007746f
C571 B.n531 VSUBS 0.007746f
C572 B.n532 VSUBS 0.007746f
C573 B.n533 VSUBS 0.007746f
C574 B.n534 VSUBS 0.007746f
C575 B.n535 VSUBS 0.007746f
C576 B.n536 VSUBS 0.007746f
C577 B.n537 VSUBS 0.007746f
C578 B.n538 VSUBS 0.007746f
C579 B.n539 VSUBS 0.007746f
C580 B.n540 VSUBS 0.007746f
C581 B.n541 VSUBS 0.007746f
C582 B.n542 VSUBS 0.007746f
C583 B.n543 VSUBS 0.007746f
C584 B.n544 VSUBS 0.007746f
C585 B.n545 VSUBS 0.007746f
C586 B.n546 VSUBS 0.007746f
C587 B.n547 VSUBS 0.007746f
C588 B.n548 VSUBS 0.007746f
C589 B.n549 VSUBS 0.007746f
C590 B.n550 VSUBS 0.007746f
C591 B.n551 VSUBS 0.017714f
C592 B.n552 VSUBS 0.018613f
C593 B.n553 VSUBS 0.018065f
C594 B.n554 VSUBS 0.007746f
C595 B.n555 VSUBS 0.007746f
C596 B.n556 VSUBS 0.007746f
C597 B.n557 VSUBS 0.007746f
C598 B.n558 VSUBS 0.007746f
C599 B.n559 VSUBS 0.007746f
C600 B.n560 VSUBS 0.007746f
C601 B.n561 VSUBS 0.007746f
C602 B.n562 VSUBS 0.007746f
C603 B.n563 VSUBS 0.007746f
C604 B.n564 VSUBS 0.007746f
C605 B.n565 VSUBS 0.007746f
C606 B.n566 VSUBS 0.007746f
C607 B.n567 VSUBS 0.007746f
C608 B.n568 VSUBS 0.007746f
C609 B.n569 VSUBS 0.007746f
C610 B.n570 VSUBS 0.007746f
C611 B.n571 VSUBS 0.007746f
C612 B.n572 VSUBS 0.007746f
C613 B.n573 VSUBS 0.007746f
C614 B.n574 VSUBS 0.007746f
C615 B.n575 VSUBS 0.007746f
C616 B.n576 VSUBS 0.007746f
C617 B.n577 VSUBS 0.007746f
C618 B.n578 VSUBS 0.007746f
C619 B.n579 VSUBS 0.007746f
C620 B.n580 VSUBS 0.007746f
C621 B.n581 VSUBS 0.007746f
C622 B.n582 VSUBS 0.007746f
C623 B.n583 VSUBS 0.007746f
C624 B.n584 VSUBS 0.007746f
C625 B.n585 VSUBS 0.007746f
C626 B.n586 VSUBS 0.007746f
C627 B.n587 VSUBS 0.007746f
C628 B.n588 VSUBS 0.007746f
C629 B.n589 VSUBS 0.007746f
C630 B.n590 VSUBS 0.007746f
C631 B.n591 VSUBS 0.007746f
C632 B.n592 VSUBS 0.007746f
C633 B.n593 VSUBS 0.007746f
C634 B.n594 VSUBS 0.007746f
C635 B.n595 VSUBS 0.007746f
C636 B.n596 VSUBS 0.007746f
C637 B.n597 VSUBS 0.007746f
C638 B.n598 VSUBS 0.007746f
C639 B.n599 VSUBS 0.007746f
C640 B.n600 VSUBS 0.007746f
C641 B.n601 VSUBS 0.007746f
C642 B.n602 VSUBS 0.007746f
C643 B.n603 VSUBS 0.007746f
C644 B.n604 VSUBS 0.007746f
C645 B.n605 VSUBS 0.007746f
C646 B.n606 VSUBS 0.007746f
C647 B.n607 VSUBS 0.007746f
C648 B.n608 VSUBS 0.007746f
C649 B.n609 VSUBS 0.007746f
C650 B.n610 VSUBS 0.007746f
C651 B.n611 VSUBS 0.007746f
C652 B.n612 VSUBS 0.007746f
C653 B.n613 VSUBS 0.007746f
C654 B.n614 VSUBS 0.007746f
C655 B.n615 VSUBS 0.007746f
C656 B.n616 VSUBS 0.007746f
C657 B.n617 VSUBS 0.007746f
C658 B.n618 VSUBS 0.007746f
C659 B.n619 VSUBS 0.007746f
C660 B.n620 VSUBS 0.007746f
C661 B.n621 VSUBS 0.007746f
C662 B.n622 VSUBS 0.007746f
C663 B.n623 VSUBS 0.007746f
C664 B.n624 VSUBS 0.007746f
C665 B.n625 VSUBS 0.007746f
C666 B.n626 VSUBS 0.007746f
C667 B.n627 VSUBS 0.007746f
C668 B.n628 VSUBS 0.007746f
C669 B.n629 VSUBS 0.007746f
C670 B.n630 VSUBS 0.007746f
C671 B.n631 VSUBS 0.007746f
C672 B.n632 VSUBS 0.007746f
C673 B.n633 VSUBS 0.007746f
C674 B.n634 VSUBS 0.007746f
C675 B.n635 VSUBS 0.007746f
C676 B.n636 VSUBS 0.007746f
C677 B.n637 VSUBS 0.007746f
C678 B.n638 VSUBS 0.007746f
C679 B.n639 VSUBS 0.007746f
C680 B.n640 VSUBS 0.007746f
C681 B.n641 VSUBS 0.007746f
C682 B.n642 VSUBS 0.00729f
C683 B.n643 VSUBS 0.017946f
C684 B.n644 VSUBS 0.004329f
C685 B.n645 VSUBS 0.007746f
C686 B.n646 VSUBS 0.007746f
C687 B.n647 VSUBS 0.007746f
C688 B.n648 VSUBS 0.007746f
C689 B.n649 VSUBS 0.007746f
C690 B.n650 VSUBS 0.007746f
C691 B.n651 VSUBS 0.007746f
C692 B.n652 VSUBS 0.007746f
C693 B.n653 VSUBS 0.007746f
C694 B.n654 VSUBS 0.007746f
C695 B.n655 VSUBS 0.007746f
C696 B.n656 VSUBS 0.007746f
C697 B.n657 VSUBS 0.004329f
C698 B.n658 VSUBS 0.007746f
C699 B.n659 VSUBS 0.007746f
C700 B.n660 VSUBS 0.007746f
C701 B.n661 VSUBS 0.007746f
C702 B.n662 VSUBS 0.007746f
C703 B.n663 VSUBS 0.007746f
C704 B.n664 VSUBS 0.007746f
C705 B.n665 VSUBS 0.007746f
C706 B.n666 VSUBS 0.007746f
C707 B.n667 VSUBS 0.007746f
C708 B.n668 VSUBS 0.007746f
C709 B.n669 VSUBS 0.007746f
C710 B.n670 VSUBS 0.007746f
C711 B.n671 VSUBS 0.007746f
C712 B.n672 VSUBS 0.007746f
C713 B.n673 VSUBS 0.007746f
C714 B.n674 VSUBS 0.007746f
C715 B.n675 VSUBS 0.007746f
C716 B.n676 VSUBS 0.007746f
C717 B.n677 VSUBS 0.007746f
C718 B.n678 VSUBS 0.007746f
C719 B.n679 VSUBS 0.007746f
C720 B.n680 VSUBS 0.007746f
C721 B.n681 VSUBS 0.007746f
C722 B.n682 VSUBS 0.007746f
C723 B.n683 VSUBS 0.007746f
C724 B.n684 VSUBS 0.007746f
C725 B.n685 VSUBS 0.007746f
C726 B.n686 VSUBS 0.007746f
C727 B.n687 VSUBS 0.007746f
C728 B.n688 VSUBS 0.007746f
C729 B.n689 VSUBS 0.007746f
C730 B.n690 VSUBS 0.007746f
C731 B.n691 VSUBS 0.007746f
C732 B.n692 VSUBS 0.007746f
C733 B.n693 VSUBS 0.007746f
C734 B.n694 VSUBS 0.007746f
C735 B.n695 VSUBS 0.007746f
C736 B.n696 VSUBS 0.007746f
C737 B.n697 VSUBS 0.007746f
C738 B.n698 VSUBS 0.007746f
C739 B.n699 VSUBS 0.007746f
C740 B.n700 VSUBS 0.007746f
C741 B.n701 VSUBS 0.007746f
C742 B.n702 VSUBS 0.007746f
C743 B.n703 VSUBS 0.007746f
C744 B.n704 VSUBS 0.007746f
C745 B.n705 VSUBS 0.007746f
C746 B.n706 VSUBS 0.007746f
C747 B.n707 VSUBS 0.007746f
C748 B.n708 VSUBS 0.007746f
C749 B.n709 VSUBS 0.007746f
C750 B.n710 VSUBS 0.007746f
C751 B.n711 VSUBS 0.007746f
C752 B.n712 VSUBS 0.007746f
C753 B.n713 VSUBS 0.007746f
C754 B.n714 VSUBS 0.007746f
C755 B.n715 VSUBS 0.007746f
C756 B.n716 VSUBS 0.007746f
C757 B.n717 VSUBS 0.007746f
C758 B.n718 VSUBS 0.007746f
C759 B.n719 VSUBS 0.007746f
C760 B.n720 VSUBS 0.007746f
C761 B.n721 VSUBS 0.007746f
C762 B.n722 VSUBS 0.007746f
C763 B.n723 VSUBS 0.007746f
C764 B.n724 VSUBS 0.007746f
C765 B.n725 VSUBS 0.007746f
C766 B.n726 VSUBS 0.007746f
C767 B.n727 VSUBS 0.007746f
C768 B.n728 VSUBS 0.007746f
C769 B.n729 VSUBS 0.007746f
C770 B.n730 VSUBS 0.007746f
C771 B.n731 VSUBS 0.007746f
C772 B.n732 VSUBS 0.007746f
C773 B.n733 VSUBS 0.007746f
C774 B.n734 VSUBS 0.007746f
C775 B.n735 VSUBS 0.007746f
C776 B.n736 VSUBS 0.007746f
C777 B.n737 VSUBS 0.007746f
C778 B.n738 VSUBS 0.007746f
C779 B.n739 VSUBS 0.007746f
C780 B.n740 VSUBS 0.007746f
C781 B.n741 VSUBS 0.007746f
C782 B.n742 VSUBS 0.007746f
C783 B.n743 VSUBS 0.007746f
C784 B.n744 VSUBS 0.007746f
C785 B.n745 VSUBS 0.007746f
C786 B.n746 VSUBS 0.007746f
C787 B.n747 VSUBS 0.018964f
C788 B.n748 VSUBS 0.018964f
C789 B.n749 VSUBS 0.017714f
C790 B.n750 VSUBS 0.007746f
C791 B.n751 VSUBS 0.007746f
C792 B.n752 VSUBS 0.007746f
C793 B.n753 VSUBS 0.007746f
C794 B.n754 VSUBS 0.007746f
C795 B.n755 VSUBS 0.007746f
C796 B.n756 VSUBS 0.007746f
C797 B.n757 VSUBS 0.007746f
C798 B.n758 VSUBS 0.007746f
C799 B.n759 VSUBS 0.007746f
C800 B.n760 VSUBS 0.007746f
C801 B.n761 VSUBS 0.007746f
C802 B.n762 VSUBS 0.007746f
C803 B.n763 VSUBS 0.007746f
C804 B.n764 VSUBS 0.007746f
C805 B.n765 VSUBS 0.007746f
C806 B.n766 VSUBS 0.007746f
C807 B.n767 VSUBS 0.007746f
C808 B.n768 VSUBS 0.007746f
C809 B.n769 VSUBS 0.007746f
C810 B.n770 VSUBS 0.007746f
C811 B.n771 VSUBS 0.007746f
C812 B.n772 VSUBS 0.007746f
C813 B.n773 VSUBS 0.007746f
C814 B.n774 VSUBS 0.007746f
C815 B.n775 VSUBS 0.007746f
C816 B.n776 VSUBS 0.007746f
C817 B.n777 VSUBS 0.007746f
C818 B.n778 VSUBS 0.007746f
C819 B.n779 VSUBS 0.007746f
C820 B.n780 VSUBS 0.007746f
C821 B.n781 VSUBS 0.007746f
C822 B.n782 VSUBS 0.007746f
C823 B.n783 VSUBS 0.007746f
C824 B.n784 VSUBS 0.007746f
C825 B.n785 VSUBS 0.007746f
C826 B.n786 VSUBS 0.007746f
C827 B.n787 VSUBS 0.007746f
C828 B.n788 VSUBS 0.007746f
C829 B.n789 VSUBS 0.007746f
C830 B.n790 VSUBS 0.007746f
C831 B.n791 VSUBS 0.007746f
C832 B.n792 VSUBS 0.007746f
C833 B.n793 VSUBS 0.007746f
C834 B.n794 VSUBS 0.007746f
C835 B.n795 VSUBS 0.007746f
C836 B.n796 VSUBS 0.007746f
C837 B.n797 VSUBS 0.007746f
C838 B.n798 VSUBS 0.007746f
C839 B.n799 VSUBS 0.017539f
C840 VDD1.n0 VSUBS 0.029913f
C841 VDD1.n1 VSUBS 0.026809f
C842 VDD1.n2 VSUBS 0.014406f
C843 VDD1.n3 VSUBS 0.03405f
C844 VDD1.n4 VSUBS 0.015253f
C845 VDD1.n5 VSUBS 0.026809f
C846 VDD1.n6 VSUBS 0.014406f
C847 VDD1.n7 VSUBS 0.03405f
C848 VDD1.n8 VSUBS 0.015253f
C849 VDD1.n9 VSUBS 0.026809f
C850 VDD1.n10 VSUBS 0.01483f
C851 VDD1.n11 VSUBS 0.03405f
C852 VDD1.n12 VSUBS 0.014406f
C853 VDD1.n13 VSUBS 0.015253f
C854 VDD1.n14 VSUBS 0.026809f
C855 VDD1.n15 VSUBS 0.014406f
C856 VDD1.n16 VSUBS 0.03405f
C857 VDD1.n17 VSUBS 0.015253f
C858 VDD1.n18 VSUBS 0.026809f
C859 VDD1.n19 VSUBS 0.014406f
C860 VDD1.n20 VSUBS 0.03405f
C861 VDD1.n21 VSUBS 0.015253f
C862 VDD1.n22 VSUBS 0.026809f
C863 VDD1.n23 VSUBS 0.014406f
C864 VDD1.n24 VSUBS 0.03405f
C865 VDD1.n25 VSUBS 0.015253f
C866 VDD1.n26 VSUBS 0.026809f
C867 VDD1.n27 VSUBS 0.014406f
C868 VDD1.n28 VSUBS 0.03405f
C869 VDD1.n29 VSUBS 0.015253f
C870 VDD1.n30 VSUBS 0.026809f
C871 VDD1.n31 VSUBS 0.014406f
C872 VDD1.n32 VSUBS 0.025538f
C873 VDD1.n33 VSUBS 0.021661f
C874 VDD1.t5 VSUBS 0.073114f
C875 VDD1.n34 VSUBS 0.214994f
C876 VDD1.n35 VSUBS 2.1122f
C877 VDD1.n36 VSUBS 0.014406f
C878 VDD1.n37 VSUBS 0.015253f
C879 VDD1.n38 VSUBS 0.03405f
C880 VDD1.n39 VSUBS 0.03405f
C881 VDD1.n40 VSUBS 0.015253f
C882 VDD1.n41 VSUBS 0.014406f
C883 VDD1.n42 VSUBS 0.026809f
C884 VDD1.n43 VSUBS 0.026809f
C885 VDD1.n44 VSUBS 0.014406f
C886 VDD1.n45 VSUBS 0.015253f
C887 VDD1.n46 VSUBS 0.03405f
C888 VDD1.n47 VSUBS 0.03405f
C889 VDD1.n48 VSUBS 0.015253f
C890 VDD1.n49 VSUBS 0.014406f
C891 VDD1.n50 VSUBS 0.026809f
C892 VDD1.n51 VSUBS 0.026809f
C893 VDD1.n52 VSUBS 0.014406f
C894 VDD1.n53 VSUBS 0.015253f
C895 VDD1.n54 VSUBS 0.03405f
C896 VDD1.n55 VSUBS 0.03405f
C897 VDD1.n56 VSUBS 0.015253f
C898 VDD1.n57 VSUBS 0.014406f
C899 VDD1.n58 VSUBS 0.026809f
C900 VDD1.n59 VSUBS 0.026809f
C901 VDD1.n60 VSUBS 0.014406f
C902 VDD1.n61 VSUBS 0.015253f
C903 VDD1.n62 VSUBS 0.03405f
C904 VDD1.n63 VSUBS 0.03405f
C905 VDD1.n64 VSUBS 0.015253f
C906 VDD1.n65 VSUBS 0.014406f
C907 VDD1.n66 VSUBS 0.026809f
C908 VDD1.n67 VSUBS 0.026809f
C909 VDD1.n68 VSUBS 0.014406f
C910 VDD1.n69 VSUBS 0.015253f
C911 VDD1.n70 VSUBS 0.03405f
C912 VDD1.n71 VSUBS 0.03405f
C913 VDD1.n72 VSUBS 0.015253f
C914 VDD1.n73 VSUBS 0.014406f
C915 VDD1.n74 VSUBS 0.026809f
C916 VDD1.n75 VSUBS 0.026809f
C917 VDD1.n76 VSUBS 0.014406f
C918 VDD1.n77 VSUBS 0.015253f
C919 VDD1.n78 VSUBS 0.03405f
C920 VDD1.n79 VSUBS 0.03405f
C921 VDD1.n80 VSUBS 0.03405f
C922 VDD1.n81 VSUBS 0.01483f
C923 VDD1.n82 VSUBS 0.014406f
C924 VDD1.n83 VSUBS 0.026809f
C925 VDD1.n84 VSUBS 0.026809f
C926 VDD1.n85 VSUBS 0.014406f
C927 VDD1.n86 VSUBS 0.015253f
C928 VDD1.n87 VSUBS 0.03405f
C929 VDD1.n88 VSUBS 0.03405f
C930 VDD1.n89 VSUBS 0.015253f
C931 VDD1.n90 VSUBS 0.014406f
C932 VDD1.n91 VSUBS 0.026809f
C933 VDD1.n92 VSUBS 0.026809f
C934 VDD1.n93 VSUBS 0.014406f
C935 VDD1.n94 VSUBS 0.015253f
C936 VDD1.n95 VSUBS 0.03405f
C937 VDD1.n96 VSUBS 0.083985f
C938 VDD1.n97 VSUBS 0.015253f
C939 VDD1.n98 VSUBS 0.014406f
C940 VDD1.n99 VSUBS 0.063798f
C941 VDD1.n100 VSUBS 0.065803f
C942 VDD1.n101 VSUBS 0.029913f
C943 VDD1.n102 VSUBS 0.026809f
C944 VDD1.n103 VSUBS 0.014406f
C945 VDD1.n104 VSUBS 0.03405f
C946 VDD1.n105 VSUBS 0.015253f
C947 VDD1.n106 VSUBS 0.026809f
C948 VDD1.n107 VSUBS 0.014406f
C949 VDD1.n108 VSUBS 0.03405f
C950 VDD1.n109 VSUBS 0.015253f
C951 VDD1.n110 VSUBS 0.026809f
C952 VDD1.n111 VSUBS 0.01483f
C953 VDD1.n112 VSUBS 0.03405f
C954 VDD1.n113 VSUBS 0.015253f
C955 VDD1.n114 VSUBS 0.026809f
C956 VDD1.n115 VSUBS 0.014406f
C957 VDD1.n116 VSUBS 0.03405f
C958 VDD1.n117 VSUBS 0.015253f
C959 VDD1.n118 VSUBS 0.026809f
C960 VDD1.n119 VSUBS 0.014406f
C961 VDD1.n120 VSUBS 0.03405f
C962 VDD1.n121 VSUBS 0.015253f
C963 VDD1.n122 VSUBS 0.026809f
C964 VDD1.n123 VSUBS 0.014406f
C965 VDD1.n124 VSUBS 0.03405f
C966 VDD1.n125 VSUBS 0.015253f
C967 VDD1.n126 VSUBS 0.026809f
C968 VDD1.n127 VSUBS 0.014406f
C969 VDD1.n128 VSUBS 0.03405f
C970 VDD1.n129 VSUBS 0.015253f
C971 VDD1.n130 VSUBS 0.026809f
C972 VDD1.n131 VSUBS 0.014406f
C973 VDD1.n132 VSUBS 0.025538f
C974 VDD1.n133 VSUBS 0.021661f
C975 VDD1.t0 VSUBS 0.073114f
C976 VDD1.n134 VSUBS 0.214994f
C977 VDD1.n135 VSUBS 2.1122f
C978 VDD1.n136 VSUBS 0.014406f
C979 VDD1.n137 VSUBS 0.015253f
C980 VDD1.n138 VSUBS 0.03405f
C981 VDD1.n139 VSUBS 0.03405f
C982 VDD1.n140 VSUBS 0.015253f
C983 VDD1.n141 VSUBS 0.014406f
C984 VDD1.n142 VSUBS 0.026809f
C985 VDD1.n143 VSUBS 0.026809f
C986 VDD1.n144 VSUBS 0.014406f
C987 VDD1.n145 VSUBS 0.015253f
C988 VDD1.n146 VSUBS 0.03405f
C989 VDD1.n147 VSUBS 0.03405f
C990 VDD1.n148 VSUBS 0.015253f
C991 VDD1.n149 VSUBS 0.014406f
C992 VDD1.n150 VSUBS 0.026809f
C993 VDD1.n151 VSUBS 0.026809f
C994 VDD1.n152 VSUBS 0.014406f
C995 VDD1.n153 VSUBS 0.015253f
C996 VDD1.n154 VSUBS 0.03405f
C997 VDD1.n155 VSUBS 0.03405f
C998 VDD1.n156 VSUBS 0.015253f
C999 VDD1.n157 VSUBS 0.014406f
C1000 VDD1.n158 VSUBS 0.026809f
C1001 VDD1.n159 VSUBS 0.026809f
C1002 VDD1.n160 VSUBS 0.014406f
C1003 VDD1.n161 VSUBS 0.015253f
C1004 VDD1.n162 VSUBS 0.03405f
C1005 VDD1.n163 VSUBS 0.03405f
C1006 VDD1.n164 VSUBS 0.015253f
C1007 VDD1.n165 VSUBS 0.014406f
C1008 VDD1.n166 VSUBS 0.026809f
C1009 VDD1.n167 VSUBS 0.026809f
C1010 VDD1.n168 VSUBS 0.014406f
C1011 VDD1.n169 VSUBS 0.015253f
C1012 VDD1.n170 VSUBS 0.03405f
C1013 VDD1.n171 VSUBS 0.03405f
C1014 VDD1.n172 VSUBS 0.015253f
C1015 VDD1.n173 VSUBS 0.014406f
C1016 VDD1.n174 VSUBS 0.026809f
C1017 VDD1.n175 VSUBS 0.026809f
C1018 VDD1.n176 VSUBS 0.014406f
C1019 VDD1.n177 VSUBS 0.014406f
C1020 VDD1.n178 VSUBS 0.015253f
C1021 VDD1.n179 VSUBS 0.03405f
C1022 VDD1.n180 VSUBS 0.03405f
C1023 VDD1.n181 VSUBS 0.03405f
C1024 VDD1.n182 VSUBS 0.01483f
C1025 VDD1.n183 VSUBS 0.014406f
C1026 VDD1.n184 VSUBS 0.026809f
C1027 VDD1.n185 VSUBS 0.026809f
C1028 VDD1.n186 VSUBS 0.014406f
C1029 VDD1.n187 VSUBS 0.015253f
C1030 VDD1.n188 VSUBS 0.03405f
C1031 VDD1.n189 VSUBS 0.03405f
C1032 VDD1.n190 VSUBS 0.015253f
C1033 VDD1.n191 VSUBS 0.014406f
C1034 VDD1.n192 VSUBS 0.026809f
C1035 VDD1.n193 VSUBS 0.026809f
C1036 VDD1.n194 VSUBS 0.014406f
C1037 VDD1.n195 VSUBS 0.015253f
C1038 VDD1.n196 VSUBS 0.03405f
C1039 VDD1.n197 VSUBS 0.083985f
C1040 VDD1.n198 VSUBS 0.015253f
C1041 VDD1.n199 VSUBS 0.014406f
C1042 VDD1.n200 VSUBS 0.063798f
C1043 VDD1.n201 VSUBS 0.06518f
C1044 VDD1.t2 VSUBS 0.387475f
C1045 VDD1.t4 VSUBS 0.387475f
C1046 VDD1.n202 VSUBS 3.23315f
C1047 VDD1.n203 VSUBS 3.33996f
C1048 VDD1.t3 VSUBS 0.387475f
C1049 VDD1.t1 VSUBS 0.387475f
C1050 VDD1.n204 VSUBS 3.22894f
C1051 VDD1.n205 VSUBS 3.5685f
C1052 VP.n0 VSUBS 0.034523f
C1053 VP.t1 VSUBS 3.12712f
C1054 VP.n1 VSUBS 0.02983f
C1055 VP.n2 VSUBS 0.034523f
C1056 VP.t3 VSUBS 3.12712f
C1057 VP.n3 VSUBS 0.02983f
C1058 VP.n4 VSUBS 0.034523f
C1059 VP.t5 VSUBS 3.12712f
C1060 VP.n5 VSUBS 0.034523f
C1061 VP.t4 VSUBS 3.12712f
C1062 VP.n6 VSUBS 0.02983f
C1063 VP.t0 VSUBS 3.28922f
C1064 VP.n7 VSUBS 1.16626f
C1065 VP.t2 VSUBS 3.12712f
C1066 VP.n8 VSUBS 1.18684f
C1067 VP.n9 VSUBS 0.069758f
C1068 VP.n10 VSUBS 0.255574f
C1069 VP.n11 VSUBS 0.034523f
C1070 VP.n12 VSUBS 0.034523f
C1071 VP.n13 VSUBS 0.065555f
C1072 VP.n14 VSUBS 0.040835f
C1073 VP.n15 VSUBS 1.1759f
C1074 VP.n16 VSUBS 1.90007f
C1075 VP.n17 VSUBS 1.92477f
C1076 VP.n18 VSUBS 1.1759f
C1077 VP.n19 VSUBS 0.040835f
C1078 VP.n20 VSUBS 0.065555f
C1079 VP.n21 VSUBS 0.034523f
C1080 VP.n22 VSUBS 0.034523f
C1081 VP.n23 VSUBS 0.034523f
C1082 VP.n24 VSUBS 0.069758f
C1083 VP.n25 VSUBS 1.12607f
C1084 VP.n26 VSUBS 0.069758f
C1085 VP.n27 VSUBS 0.034523f
C1086 VP.n28 VSUBS 0.034523f
C1087 VP.n29 VSUBS 0.034523f
C1088 VP.n30 VSUBS 0.065555f
C1089 VP.n31 VSUBS 0.040835f
C1090 VP.n32 VSUBS 1.1759f
C1091 VP.n33 VSUBS 0.036004f
C1092 VDD2.n0 VSUBS 0.029912f
C1093 VDD2.n1 VSUBS 0.026808f
C1094 VDD2.n2 VSUBS 0.014405f
C1095 VDD2.n3 VSUBS 0.034049f
C1096 VDD2.n4 VSUBS 0.015253f
C1097 VDD2.n5 VSUBS 0.026808f
C1098 VDD2.n6 VSUBS 0.014405f
C1099 VDD2.n7 VSUBS 0.034049f
C1100 VDD2.n8 VSUBS 0.015253f
C1101 VDD2.n9 VSUBS 0.026808f
C1102 VDD2.n10 VSUBS 0.014829f
C1103 VDD2.n11 VSUBS 0.034049f
C1104 VDD2.n12 VSUBS 0.015253f
C1105 VDD2.n13 VSUBS 0.026808f
C1106 VDD2.n14 VSUBS 0.014405f
C1107 VDD2.n15 VSUBS 0.034049f
C1108 VDD2.n16 VSUBS 0.015253f
C1109 VDD2.n17 VSUBS 0.026808f
C1110 VDD2.n18 VSUBS 0.014405f
C1111 VDD2.n19 VSUBS 0.034049f
C1112 VDD2.n20 VSUBS 0.015253f
C1113 VDD2.n21 VSUBS 0.026808f
C1114 VDD2.n22 VSUBS 0.014405f
C1115 VDD2.n23 VSUBS 0.034049f
C1116 VDD2.n24 VSUBS 0.015253f
C1117 VDD2.n25 VSUBS 0.026808f
C1118 VDD2.n26 VSUBS 0.014405f
C1119 VDD2.n27 VSUBS 0.034049f
C1120 VDD2.n28 VSUBS 0.015253f
C1121 VDD2.n29 VSUBS 0.026808f
C1122 VDD2.n30 VSUBS 0.014405f
C1123 VDD2.n31 VSUBS 0.025537f
C1124 VDD2.n32 VSUBS 0.02166f
C1125 VDD2.t4 VSUBS 0.073111f
C1126 VDD2.n33 VSUBS 0.214985f
C1127 VDD2.n34 VSUBS 2.11211f
C1128 VDD2.n35 VSUBS 0.014405f
C1129 VDD2.n36 VSUBS 0.015253f
C1130 VDD2.n37 VSUBS 0.034049f
C1131 VDD2.n38 VSUBS 0.034049f
C1132 VDD2.n39 VSUBS 0.015253f
C1133 VDD2.n40 VSUBS 0.014405f
C1134 VDD2.n41 VSUBS 0.026808f
C1135 VDD2.n42 VSUBS 0.026808f
C1136 VDD2.n43 VSUBS 0.014405f
C1137 VDD2.n44 VSUBS 0.015253f
C1138 VDD2.n45 VSUBS 0.034049f
C1139 VDD2.n46 VSUBS 0.034049f
C1140 VDD2.n47 VSUBS 0.015253f
C1141 VDD2.n48 VSUBS 0.014405f
C1142 VDD2.n49 VSUBS 0.026808f
C1143 VDD2.n50 VSUBS 0.026808f
C1144 VDD2.n51 VSUBS 0.014405f
C1145 VDD2.n52 VSUBS 0.015253f
C1146 VDD2.n53 VSUBS 0.034049f
C1147 VDD2.n54 VSUBS 0.034049f
C1148 VDD2.n55 VSUBS 0.015253f
C1149 VDD2.n56 VSUBS 0.014405f
C1150 VDD2.n57 VSUBS 0.026808f
C1151 VDD2.n58 VSUBS 0.026808f
C1152 VDD2.n59 VSUBS 0.014405f
C1153 VDD2.n60 VSUBS 0.015253f
C1154 VDD2.n61 VSUBS 0.034049f
C1155 VDD2.n62 VSUBS 0.034049f
C1156 VDD2.n63 VSUBS 0.015253f
C1157 VDD2.n64 VSUBS 0.014405f
C1158 VDD2.n65 VSUBS 0.026808f
C1159 VDD2.n66 VSUBS 0.026808f
C1160 VDD2.n67 VSUBS 0.014405f
C1161 VDD2.n68 VSUBS 0.015253f
C1162 VDD2.n69 VSUBS 0.034049f
C1163 VDD2.n70 VSUBS 0.034049f
C1164 VDD2.n71 VSUBS 0.015253f
C1165 VDD2.n72 VSUBS 0.014405f
C1166 VDD2.n73 VSUBS 0.026808f
C1167 VDD2.n74 VSUBS 0.026808f
C1168 VDD2.n75 VSUBS 0.014405f
C1169 VDD2.n76 VSUBS 0.014405f
C1170 VDD2.n77 VSUBS 0.015253f
C1171 VDD2.n78 VSUBS 0.034049f
C1172 VDD2.n79 VSUBS 0.034049f
C1173 VDD2.n80 VSUBS 0.034049f
C1174 VDD2.n81 VSUBS 0.014829f
C1175 VDD2.n82 VSUBS 0.014405f
C1176 VDD2.n83 VSUBS 0.026808f
C1177 VDD2.n84 VSUBS 0.026808f
C1178 VDD2.n85 VSUBS 0.014405f
C1179 VDD2.n86 VSUBS 0.015253f
C1180 VDD2.n87 VSUBS 0.034049f
C1181 VDD2.n88 VSUBS 0.034049f
C1182 VDD2.n89 VSUBS 0.015253f
C1183 VDD2.n90 VSUBS 0.014405f
C1184 VDD2.n91 VSUBS 0.026808f
C1185 VDD2.n92 VSUBS 0.026808f
C1186 VDD2.n93 VSUBS 0.014405f
C1187 VDD2.n94 VSUBS 0.015253f
C1188 VDD2.n95 VSUBS 0.034049f
C1189 VDD2.n96 VSUBS 0.083982f
C1190 VDD2.n97 VSUBS 0.015253f
C1191 VDD2.n98 VSUBS 0.014405f
C1192 VDD2.n99 VSUBS 0.063796f
C1193 VDD2.n100 VSUBS 0.065178f
C1194 VDD2.t2 VSUBS 0.387459f
C1195 VDD2.t1 VSUBS 0.387459f
C1196 VDD2.n101 VSUBS 3.23302f
C1197 VDD2.n102 VSUBS 3.22516f
C1198 VDD2.n103 VSUBS 0.029912f
C1199 VDD2.n104 VSUBS 0.026808f
C1200 VDD2.n105 VSUBS 0.014405f
C1201 VDD2.n106 VSUBS 0.034049f
C1202 VDD2.n107 VSUBS 0.015253f
C1203 VDD2.n108 VSUBS 0.026808f
C1204 VDD2.n109 VSUBS 0.014405f
C1205 VDD2.n110 VSUBS 0.034049f
C1206 VDD2.n111 VSUBS 0.015253f
C1207 VDD2.n112 VSUBS 0.026808f
C1208 VDD2.n113 VSUBS 0.014829f
C1209 VDD2.n114 VSUBS 0.034049f
C1210 VDD2.n115 VSUBS 0.014405f
C1211 VDD2.n116 VSUBS 0.015253f
C1212 VDD2.n117 VSUBS 0.026808f
C1213 VDD2.n118 VSUBS 0.014405f
C1214 VDD2.n119 VSUBS 0.034049f
C1215 VDD2.n120 VSUBS 0.015253f
C1216 VDD2.n121 VSUBS 0.026808f
C1217 VDD2.n122 VSUBS 0.014405f
C1218 VDD2.n123 VSUBS 0.034049f
C1219 VDD2.n124 VSUBS 0.015253f
C1220 VDD2.n125 VSUBS 0.026808f
C1221 VDD2.n126 VSUBS 0.014405f
C1222 VDD2.n127 VSUBS 0.034049f
C1223 VDD2.n128 VSUBS 0.015253f
C1224 VDD2.n129 VSUBS 0.026808f
C1225 VDD2.n130 VSUBS 0.014405f
C1226 VDD2.n131 VSUBS 0.034049f
C1227 VDD2.n132 VSUBS 0.015253f
C1228 VDD2.n133 VSUBS 0.026808f
C1229 VDD2.n134 VSUBS 0.014405f
C1230 VDD2.n135 VSUBS 0.025537f
C1231 VDD2.n136 VSUBS 0.02166f
C1232 VDD2.t5 VSUBS 0.073111f
C1233 VDD2.n137 VSUBS 0.214985f
C1234 VDD2.n138 VSUBS 2.11211f
C1235 VDD2.n139 VSUBS 0.014405f
C1236 VDD2.n140 VSUBS 0.015253f
C1237 VDD2.n141 VSUBS 0.034049f
C1238 VDD2.n142 VSUBS 0.034049f
C1239 VDD2.n143 VSUBS 0.015253f
C1240 VDD2.n144 VSUBS 0.014405f
C1241 VDD2.n145 VSUBS 0.026808f
C1242 VDD2.n146 VSUBS 0.026808f
C1243 VDD2.n147 VSUBS 0.014405f
C1244 VDD2.n148 VSUBS 0.015253f
C1245 VDD2.n149 VSUBS 0.034049f
C1246 VDD2.n150 VSUBS 0.034049f
C1247 VDD2.n151 VSUBS 0.015253f
C1248 VDD2.n152 VSUBS 0.014405f
C1249 VDD2.n153 VSUBS 0.026808f
C1250 VDD2.n154 VSUBS 0.026808f
C1251 VDD2.n155 VSUBS 0.014405f
C1252 VDD2.n156 VSUBS 0.015253f
C1253 VDD2.n157 VSUBS 0.034049f
C1254 VDD2.n158 VSUBS 0.034049f
C1255 VDD2.n159 VSUBS 0.015253f
C1256 VDD2.n160 VSUBS 0.014405f
C1257 VDD2.n161 VSUBS 0.026808f
C1258 VDD2.n162 VSUBS 0.026808f
C1259 VDD2.n163 VSUBS 0.014405f
C1260 VDD2.n164 VSUBS 0.015253f
C1261 VDD2.n165 VSUBS 0.034049f
C1262 VDD2.n166 VSUBS 0.034049f
C1263 VDD2.n167 VSUBS 0.015253f
C1264 VDD2.n168 VSUBS 0.014405f
C1265 VDD2.n169 VSUBS 0.026808f
C1266 VDD2.n170 VSUBS 0.026808f
C1267 VDD2.n171 VSUBS 0.014405f
C1268 VDD2.n172 VSUBS 0.015253f
C1269 VDD2.n173 VSUBS 0.034049f
C1270 VDD2.n174 VSUBS 0.034049f
C1271 VDD2.n175 VSUBS 0.015253f
C1272 VDD2.n176 VSUBS 0.014405f
C1273 VDD2.n177 VSUBS 0.026808f
C1274 VDD2.n178 VSUBS 0.026808f
C1275 VDD2.n179 VSUBS 0.014405f
C1276 VDD2.n180 VSUBS 0.015253f
C1277 VDD2.n181 VSUBS 0.034049f
C1278 VDD2.n182 VSUBS 0.034049f
C1279 VDD2.n183 VSUBS 0.034049f
C1280 VDD2.n184 VSUBS 0.014829f
C1281 VDD2.n185 VSUBS 0.014405f
C1282 VDD2.n186 VSUBS 0.026808f
C1283 VDD2.n187 VSUBS 0.026808f
C1284 VDD2.n188 VSUBS 0.014405f
C1285 VDD2.n189 VSUBS 0.015253f
C1286 VDD2.n190 VSUBS 0.034049f
C1287 VDD2.n191 VSUBS 0.034049f
C1288 VDD2.n192 VSUBS 0.015253f
C1289 VDD2.n193 VSUBS 0.014405f
C1290 VDD2.n194 VSUBS 0.026808f
C1291 VDD2.n195 VSUBS 0.026808f
C1292 VDD2.n196 VSUBS 0.014405f
C1293 VDD2.n197 VSUBS 0.015253f
C1294 VDD2.n198 VSUBS 0.034049f
C1295 VDD2.n199 VSUBS 0.083982f
C1296 VDD2.n200 VSUBS 0.015253f
C1297 VDD2.n201 VSUBS 0.014405f
C1298 VDD2.n202 VSUBS 0.063796f
C1299 VDD2.n203 VSUBS 0.060854f
C1300 VDD2.n204 VSUBS 3.03048f
C1301 VDD2.t0 VSUBS 0.387459f
C1302 VDD2.t3 VSUBS 0.387459f
C1303 VDD2.n205 VSUBS 3.23298f
C1304 VTAIL.t9 VSUBS 0.393442f
C1305 VTAIL.t11 VSUBS 0.393442f
C1306 VTAIL.n0 VSUBS 3.11209f
C1307 VTAIL.n1 VSUBS 0.830946f
C1308 VTAIL.n2 VSUBS 0.030374f
C1309 VTAIL.n3 VSUBS 0.027222f
C1310 VTAIL.n4 VSUBS 0.014628f
C1311 VTAIL.n5 VSUBS 0.034575f
C1312 VTAIL.n6 VSUBS 0.015488f
C1313 VTAIL.n7 VSUBS 0.027222f
C1314 VTAIL.n8 VSUBS 0.014628f
C1315 VTAIL.n9 VSUBS 0.034575f
C1316 VTAIL.n10 VSUBS 0.015488f
C1317 VTAIL.n11 VSUBS 0.027222f
C1318 VTAIL.n12 VSUBS 0.015058f
C1319 VTAIL.n13 VSUBS 0.034575f
C1320 VTAIL.n14 VSUBS 0.015488f
C1321 VTAIL.n15 VSUBS 0.027222f
C1322 VTAIL.n16 VSUBS 0.014628f
C1323 VTAIL.n17 VSUBS 0.034575f
C1324 VTAIL.n18 VSUBS 0.015488f
C1325 VTAIL.n19 VSUBS 0.027222f
C1326 VTAIL.n20 VSUBS 0.014628f
C1327 VTAIL.n21 VSUBS 0.034575f
C1328 VTAIL.n22 VSUBS 0.015488f
C1329 VTAIL.n23 VSUBS 0.027222f
C1330 VTAIL.n24 VSUBS 0.014628f
C1331 VTAIL.n25 VSUBS 0.034575f
C1332 VTAIL.n26 VSUBS 0.015488f
C1333 VTAIL.n27 VSUBS 0.027222f
C1334 VTAIL.n28 VSUBS 0.014628f
C1335 VTAIL.n29 VSUBS 0.034575f
C1336 VTAIL.n30 VSUBS 0.015488f
C1337 VTAIL.n31 VSUBS 0.027222f
C1338 VTAIL.n32 VSUBS 0.014628f
C1339 VTAIL.n33 VSUBS 0.025931f
C1340 VTAIL.n34 VSUBS 0.021995f
C1341 VTAIL.t3 VSUBS 0.07424f
C1342 VTAIL.n35 VSUBS 0.218305f
C1343 VTAIL.n36 VSUBS 2.14473f
C1344 VTAIL.n37 VSUBS 0.014628f
C1345 VTAIL.n38 VSUBS 0.015488f
C1346 VTAIL.n39 VSUBS 0.034575f
C1347 VTAIL.n40 VSUBS 0.034575f
C1348 VTAIL.n41 VSUBS 0.015488f
C1349 VTAIL.n42 VSUBS 0.014628f
C1350 VTAIL.n43 VSUBS 0.027222f
C1351 VTAIL.n44 VSUBS 0.027222f
C1352 VTAIL.n45 VSUBS 0.014628f
C1353 VTAIL.n46 VSUBS 0.015488f
C1354 VTAIL.n47 VSUBS 0.034575f
C1355 VTAIL.n48 VSUBS 0.034575f
C1356 VTAIL.n49 VSUBS 0.015488f
C1357 VTAIL.n50 VSUBS 0.014628f
C1358 VTAIL.n51 VSUBS 0.027222f
C1359 VTAIL.n52 VSUBS 0.027222f
C1360 VTAIL.n53 VSUBS 0.014628f
C1361 VTAIL.n54 VSUBS 0.015488f
C1362 VTAIL.n55 VSUBS 0.034575f
C1363 VTAIL.n56 VSUBS 0.034575f
C1364 VTAIL.n57 VSUBS 0.015488f
C1365 VTAIL.n58 VSUBS 0.014628f
C1366 VTAIL.n59 VSUBS 0.027222f
C1367 VTAIL.n60 VSUBS 0.027222f
C1368 VTAIL.n61 VSUBS 0.014628f
C1369 VTAIL.n62 VSUBS 0.015488f
C1370 VTAIL.n63 VSUBS 0.034575f
C1371 VTAIL.n64 VSUBS 0.034575f
C1372 VTAIL.n65 VSUBS 0.015488f
C1373 VTAIL.n66 VSUBS 0.014628f
C1374 VTAIL.n67 VSUBS 0.027222f
C1375 VTAIL.n68 VSUBS 0.027222f
C1376 VTAIL.n69 VSUBS 0.014628f
C1377 VTAIL.n70 VSUBS 0.015488f
C1378 VTAIL.n71 VSUBS 0.034575f
C1379 VTAIL.n72 VSUBS 0.034575f
C1380 VTAIL.n73 VSUBS 0.015488f
C1381 VTAIL.n74 VSUBS 0.014628f
C1382 VTAIL.n75 VSUBS 0.027222f
C1383 VTAIL.n76 VSUBS 0.027222f
C1384 VTAIL.n77 VSUBS 0.014628f
C1385 VTAIL.n78 VSUBS 0.014628f
C1386 VTAIL.n79 VSUBS 0.015488f
C1387 VTAIL.n80 VSUBS 0.034575f
C1388 VTAIL.n81 VSUBS 0.034575f
C1389 VTAIL.n82 VSUBS 0.034575f
C1390 VTAIL.n83 VSUBS 0.015058f
C1391 VTAIL.n84 VSUBS 0.014628f
C1392 VTAIL.n85 VSUBS 0.027222f
C1393 VTAIL.n86 VSUBS 0.027222f
C1394 VTAIL.n87 VSUBS 0.014628f
C1395 VTAIL.n88 VSUBS 0.015488f
C1396 VTAIL.n89 VSUBS 0.034575f
C1397 VTAIL.n90 VSUBS 0.034575f
C1398 VTAIL.n91 VSUBS 0.015488f
C1399 VTAIL.n92 VSUBS 0.014628f
C1400 VTAIL.n93 VSUBS 0.027222f
C1401 VTAIL.n94 VSUBS 0.027222f
C1402 VTAIL.n95 VSUBS 0.014628f
C1403 VTAIL.n96 VSUBS 0.015488f
C1404 VTAIL.n97 VSUBS 0.034575f
C1405 VTAIL.n98 VSUBS 0.085279f
C1406 VTAIL.n99 VSUBS 0.015488f
C1407 VTAIL.n100 VSUBS 0.014628f
C1408 VTAIL.n101 VSUBS 0.064781f
C1409 VTAIL.n102 VSUBS 0.043012f
C1410 VTAIL.n103 VSUBS 0.307101f
C1411 VTAIL.t5 VSUBS 0.393442f
C1412 VTAIL.t1 VSUBS 0.393442f
C1413 VTAIL.n104 VSUBS 3.11209f
C1414 VTAIL.n105 VSUBS 2.8998f
C1415 VTAIL.t10 VSUBS 0.393442f
C1416 VTAIL.t7 VSUBS 0.393442f
C1417 VTAIL.n106 VSUBS 3.11211f
C1418 VTAIL.n107 VSUBS 2.89978f
C1419 VTAIL.n108 VSUBS 0.030374f
C1420 VTAIL.n109 VSUBS 0.027222f
C1421 VTAIL.n110 VSUBS 0.014628f
C1422 VTAIL.n111 VSUBS 0.034575f
C1423 VTAIL.n112 VSUBS 0.015488f
C1424 VTAIL.n113 VSUBS 0.027222f
C1425 VTAIL.n114 VSUBS 0.014628f
C1426 VTAIL.n115 VSUBS 0.034575f
C1427 VTAIL.n116 VSUBS 0.015488f
C1428 VTAIL.n117 VSUBS 0.027222f
C1429 VTAIL.n118 VSUBS 0.015058f
C1430 VTAIL.n119 VSUBS 0.034575f
C1431 VTAIL.n120 VSUBS 0.014628f
C1432 VTAIL.n121 VSUBS 0.015488f
C1433 VTAIL.n122 VSUBS 0.027222f
C1434 VTAIL.n123 VSUBS 0.014628f
C1435 VTAIL.n124 VSUBS 0.034575f
C1436 VTAIL.n125 VSUBS 0.015488f
C1437 VTAIL.n126 VSUBS 0.027222f
C1438 VTAIL.n127 VSUBS 0.014628f
C1439 VTAIL.n128 VSUBS 0.034575f
C1440 VTAIL.n129 VSUBS 0.015488f
C1441 VTAIL.n130 VSUBS 0.027222f
C1442 VTAIL.n131 VSUBS 0.014628f
C1443 VTAIL.n132 VSUBS 0.034575f
C1444 VTAIL.n133 VSUBS 0.015488f
C1445 VTAIL.n134 VSUBS 0.027222f
C1446 VTAIL.n135 VSUBS 0.014628f
C1447 VTAIL.n136 VSUBS 0.034575f
C1448 VTAIL.n137 VSUBS 0.015488f
C1449 VTAIL.n138 VSUBS 0.027222f
C1450 VTAIL.n139 VSUBS 0.014628f
C1451 VTAIL.n140 VSUBS 0.025931f
C1452 VTAIL.n141 VSUBS 0.021995f
C1453 VTAIL.t8 VSUBS 0.07424f
C1454 VTAIL.n142 VSUBS 0.218305f
C1455 VTAIL.n143 VSUBS 2.14473f
C1456 VTAIL.n144 VSUBS 0.014628f
C1457 VTAIL.n145 VSUBS 0.015488f
C1458 VTAIL.n146 VSUBS 0.034575f
C1459 VTAIL.n147 VSUBS 0.034575f
C1460 VTAIL.n148 VSUBS 0.015488f
C1461 VTAIL.n149 VSUBS 0.014628f
C1462 VTAIL.n150 VSUBS 0.027222f
C1463 VTAIL.n151 VSUBS 0.027222f
C1464 VTAIL.n152 VSUBS 0.014628f
C1465 VTAIL.n153 VSUBS 0.015488f
C1466 VTAIL.n154 VSUBS 0.034575f
C1467 VTAIL.n155 VSUBS 0.034575f
C1468 VTAIL.n156 VSUBS 0.015488f
C1469 VTAIL.n157 VSUBS 0.014628f
C1470 VTAIL.n158 VSUBS 0.027222f
C1471 VTAIL.n159 VSUBS 0.027222f
C1472 VTAIL.n160 VSUBS 0.014628f
C1473 VTAIL.n161 VSUBS 0.015488f
C1474 VTAIL.n162 VSUBS 0.034575f
C1475 VTAIL.n163 VSUBS 0.034575f
C1476 VTAIL.n164 VSUBS 0.015488f
C1477 VTAIL.n165 VSUBS 0.014628f
C1478 VTAIL.n166 VSUBS 0.027222f
C1479 VTAIL.n167 VSUBS 0.027222f
C1480 VTAIL.n168 VSUBS 0.014628f
C1481 VTAIL.n169 VSUBS 0.015488f
C1482 VTAIL.n170 VSUBS 0.034575f
C1483 VTAIL.n171 VSUBS 0.034575f
C1484 VTAIL.n172 VSUBS 0.015488f
C1485 VTAIL.n173 VSUBS 0.014628f
C1486 VTAIL.n174 VSUBS 0.027222f
C1487 VTAIL.n175 VSUBS 0.027222f
C1488 VTAIL.n176 VSUBS 0.014628f
C1489 VTAIL.n177 VSUBS 0.015488f
C1490 VTAIL.n178 VSUBS 0.034575f
C1491 VTAIL.n179 VSUBS 0.034575f
C1492 VTAIL.n180 VSUBS 0.015488f
C1493 VTAIL.n181 VSUBS 0.014628f
C1494 VTAIL.n182 VSUBS 0.027222f
C1495 VTAIL.n183 VSUBS 0.027222f
C1496 VTAIL.n184 VSUBS 0.014628f
C1497 VTAIL.n185 VSUBS 0.015488f
C1498 VTAIL.n186 VSUBS 0.034575f
C1499 VTAIL.n187 VSUBS 0.034575f
C1500 VTAIL.n188 VSUBS 0.034575f
C1501 VTAIL.n189 VSUBS 0.015058f
C1502 VTAIL.n190 VSUBS 0.014628f
C1503 VTAIL.n191 VSUBS 0.027222f
C1504 VTAIL.n192 VSUBS 0.027222f
C1505 VTAIL.n193 VSUBS 0.014628f
C1506 VTAIL.n194 VSUBS 0.015488f
C1507 VTAIL.n195 VSUBS 0.034575f
C1508 VTAIL.n196 VSUBS 0.034575f
C1509 VTAIL.n197 VSUBS 0.015488f
C1510 VTAIL.n198 VSUBS 0.014628f
C1511 VTAIL.n199 VSUBS 0.027222f
C1512 VTAIL.n200 VSUBS 0.027222f
C1513 VTAIL.n201 VSUBS 0.014628f
C1514 VTAIL.n202 VSUBS 0.015488f
C1515 VTAIL.n203 VSUBS 0.034575f
C1516 VTAIL.n204 VSUBS 0.085279f
C1517 VTAIL.n205 VSUBS 0.015488f
C1518 VTAIL.n206 VSUBS 0.014628f
C1519 VTAIL.n207 VSUBS 0.064781f
C1520 VTAIL.n208 VSUBS 0.043012f
C1521 VTAIL.n209 VSUBS 0.307101f
C1522 VTAIL.t2 VSUBS 0.393442f
C1523 VTAIL.t0 VSUBS 0.393442f
C1524 VTAIL.n210 VSUBS 3.11211f
C1525 VTAIL.n211 VSUBS 0.946619f
C1526 VTAIL.n212 VSUBS 0.030374f
C1527 VTAIL.n213 VSUBS 0.027222f
C1528 VTAIL.n214 VSUBS 0.014628f
C1529 VTAIL.n215 VSUBS 0.034575f
C1530 VTAIL.n216 VSUBS 0.015488f
C1531 VTAIL.n217 VSUBS 0.027222f
C1532 VTAIL.n218 VSUBS 0.014628f
C1533 VTAIL.n219 VSUBS 0.034575f
C1534 VTAIL.n220 VSUBS 0.015488f
C1535 VTAIL.n221 VSUBS 0.027222f
C1536 VTAIL.n222 VSUBS 0.015058f
C1537 VTAIL.n223 VSUBS 0.034575f
C1538 VTAIL.n224 VSUBS 0.014628f
C1539 VTAIL.n225 VSUBS 0.015488f
C1540 VTAIL.n226 VSUBS 0.027222f
C1541 VTAIL.n227 VSUBS 0.014628f
C1542 VTAIL.n228 VSUBS 0.034575f
C1543 VTAIL.n229 VSUBS 0.015488f
C1544 VTAIL.n230 VSUBS 0.027222f
C1545 VTAIL.n231 VSUBS 0.014628f
C1546 VTAIL.n232 VSUBS 0.034575f
C1547 VTAIL.n233 VSUBS 0.015488f
C1548 VTAIL.n234 VSUBS 0.027222f
C1549 VTAIL.n235 VSUBS 0.014628f
C1550 VTAIL.n236 VSUBS 0.034575f
C1551 VTAIL.n237 VSUBS 0.015488f
C1552 VTAIL.n238 VSUBS 0.027222f
C1553 VTAIL.n239 VSUBS 0.014628f
C1554 VTAIL.n240 VSUBS 0.034575f
C1555 VTAIL.n241 VSUBS 0.015488f
C1556 VTAIL.n242 VSUBS 0.027222f
C1557 VTAIL.n243 VSUBS 0.014628f
C1558 VTAIL.n244 VSUBS 0.025931f
C1559 VTAIL.n245 VSUBS 0.021995f
C1560 VTAIL.t4 VSUBS 0.07424f
C1561 VTAIL.n246 VSUBS 0.218305f
C1562 VTAIL.n247 VSUBS 2.14473f
C1563 VTAIL.n248 VSUBS 0.014628f
C1564 VTAIL.n249 VSUBS 0.015488f
C1565 VTAIL.n250 VSUBS 0.034575f
C1566 VTAIL.n251 VSUBS 0.034575f
C1567 VTAIL.n252 VSUBS 0.015488f
C1568 VTAIL.n253 VSUBS 0.014628f
C1569 VTAIL.n254 VSUBS 0.027222f
C1570 VTAIL.n255 VSUBS 0.027222f
C1571 VTAIL.n256 VSUBS 0.014628f
C1572 VTAIL.n257 VSUBS 0.015488f
C1573 VTAIL.n258 VSUBS 0.034575f
C1574 VTAIL.n259 VSUBS 0.034575f
C1575 VTAIL.n260 VSUBS 0.015488f
C1576 VTAIL.n261 VSUBS 0.014628f
C1577 VTAIL.n262 VSUBS 0.027222f
C1578 VTAIL.n263 VSUBS 0.027222f
C1579 VTAIL.n264 VSUBS 0.014628f
C1580 VTAIL.n265 VSUBS 0.015488f
C1581 VTAIL.n266 VSUBS 0.034575f
C1582 VTAIL.n267 VSUBS 0.034575f
C1583 VTAIL.n268 VSUBS 0.015488f
C1584 VTAIL.n269 VSUBS 0.014628f
C1585 VTAIL.n270 VSUBS 0.027222f
C1586 VTAIL.n271 VSUBS 0.027222f
C1587 VTAIL.n272 VSUBS 0.014628f
C1588 VTAIL.n273 VSUBS 0.015488f
C1589 VTAIL.n274 VSUBS 0.034575f
C1590 VTAIL.n275 VSUBS 0.034575f
C1591 VTAIL.n276 VSUBS 0.015488f
C1592 VTAIL.n277 VSUBS 0.014628f
C1593 VTAIL.n278 VSUBS 0.027222f
C1594 VTAIL.n279 VSUBS 0.027222f
C1595 VTAIL.n280 VSUBS 0.014628f
C1596 VTAIL.n281 VSUBS 0.015488f
C1597 VTAIL.n282 VSUBS 0.034575f
C1598 VTAIL.n283 VSUBS 0.034575f
C1599 VTAIL.n284 VSUBS 0.015488f
C1600 VTAIL.n285 VSUBS 0.014628f
C1601 VTAIL.n286 VSUBS 0.027222f
C1602 VTAIL.n287 VSUBS 0.027222f
C1603 VTAIL.n288 VSUBS 0.014628f
C1604 VTAIL.n289 VSUBS 0.015488f
C1605 VTAIL.n290 VSUBS 0.034575f
C1606 VTAIL.n291 VSUBS 0.034575f
C1607 VTAIL.n292 VSUBS 0.034575f
C1608 VTAIL.n293 VSUBS 0.015058f
C1609 VTAIL.n294 VSUBS 0.014628f
C1610 VTAIL.n295 VSUBS 0.027222f
C1611 VTAIL.n296 VSUBS 0.027222f
C1612 VTAIL.n297 VSUBS 0.014628f
C1613 VTAIL.n298 VSUBS 0.015488f
C1614 VTAIL.n299 VSUBS 0.034575f
C1615 VTAIL.n300 VSUBS 0.034575f
C1616 VTAIL.n301 VSUBS 0.015488f
C1617 VTAIL.n302 VSUBS 0.014628f
C1618 VTAIL.n303 VSUBS 0.027222f
C1619 VTAIL.n304 VSUBS 0.027222f
C1620 VTAIL.n305 VSUBS 0.014628f
C1621 VTAIL.n306 VSUBS 0.015488f
C1622 VTAIL.n307 VSUBS 0.034575f
C1623 VTAIL.n308 VSUBS 0.085279f
C1624 VTAIL.n309 VSUBS 0.015488f
C1625 VTAIL.n310 VSUBS 0.014628f
C1626 VTAIL.n311 VSUBS 0.064781f
C1627 VTAIL.n312 VSUBS 0.043012f
C1628 VTAIL.n313 VSUBS 2.0992f
C1629 VTAIL.n314 VSUBS 0.030374f
C1630 VTAIL.n315 VSUBS 0.027222f
C1631 VTAIL.n316 VSUBS 0.014628f
C1632 VTAIL.n317 VSUBS 0.034575f
C1633 VTAIL.n318 VSUBS 0.015488f
C1634 VTAIL.n319 VSUBS 0.027222f
C1635 VTAIL.n320 VSUBS 0.014628f
C1636 VTAIL.n321 VSUBS 0.034575f
C1637 VTAIL.n322 VSUBS 0.015488f
C1638 VTAIL.n323 VSUBS 0.027222f
C1639 VTAIL.n324 VSUBS 0.015058f
C1640 VTAIL.n325 VSUBS 0.034575f
C1641 VTAIL.n326 VSUBS 0.015488f
C1642 VTAIL.n327 VSUBS 0.027222f
C1643 VTAIL.n328 VSUBS 0.014628f
C1644 VTAIL.n329 VSUBS 0.034575f
C1645 VTAIL.n330 VSUBS 0.015488f
C1646 VTAIL.n331 VSUBS 0.027222f
C1647 VTAIL.n332 VSUBS 0.014628f
C1648 VTAIL.n333 VSUBS 0.034575f
C1649 VTAIL.n334 VSUBS 0.015488f
C1650 VTAIL.n335 VSUBS 0.027222f
C1651 VTAIL.n336 VSUBS 0.014628f
C1652 VTAIL.n337 VSUBS 0.034575f
C1653 VTAIL.n338 VSUBS 0.015488f
C1654 VTAIL.n339 VSUBS 0.027222f
C1655 VTAIL.n340 VSUBS 0.014628f
C1656 VTAIL.n341 VSUBS 0.034575f
C1657 VTAIL.n342 VSUBS 0.015488f
C1658 VTAIL.n343 VSUBS 0.027222f
C1659 VTAIL.n344 VSUBS 0.014628f
C1660 VTAIL.n345 VSUBS 0.025931f
C1661 VTAIL.n346 VSUBS 0.021995f
C1662 VTAIL.t6 VSUBS 0.07424f
C1663 VTAIL.n347 VSUBS 0.218305f
C1664 VTAIL.n348 VSUBS 2.14473f
C1665 VTAIL.n349 VSUBS 0.014628f
C1666 VTAIL.n350 VSUBS 0.015488f
C1667 VTAIL.n351 VSUBS 0.034575f
C1668 VTAIL.n352 VSUBS 0.034575f
C1669 VTAIL.n353 VSUBS 0.015488f
C1670 VTAIL.n354 VSUBS 0.014628f
C1671 VTAIL.n355 VSUBS 0.027222f
C1672 VTAIL.n356 VSUBS 0.027222f
C1673 VTAIL.n357 VSUBS 0.014628f
C1674 VTAIL.n358 VSUBS 0.015488f
C1675 VTAIL.n359 VSUBS 0.034575f
C1676 VTAIL.n360 VSUBS 0.034575f
C1677 VTAIL.n361 VSUBS 0.015488f
C1678 VTAIL.n362 VSUBS 0.014628f
C1679 VTAIL.n363 VSUBS 0.027222f
C1680 VTAIL.n364 VSUBS 0.027222f
C1681 VTAIL.n365 VSUBS 0.014628f
C1682 VTAIL.n366 VSUBS 0.015488f
C1683 VTAIL.n367 VSUBS 0.034575f
C1684 VTAIL.n368 VSUBS 0.034575f
C1685 VTAIL.n369 VSUBS 0.015488f
C1686 VTAIL.n370 VSUBS 0.014628f
C1687 VTAIL.n371 VSUBS 0.027222f
C1688 VTAIL.n372 VSUBS 0.027222f
C1689 VTAIL.n373 VSUBS 0.014628f
C1690 VTAIL.n374 VSUBS 0.015488f
C1691 VTAIL.n375 VSUBS 0.034575f
C1692 VTAIL.n376 VSUBS 0.034575f
C1693 VTAIL.n377 VSUBS 0.015488f
C1694 VTAIL.n378 VSUBS 0.014628f
C1695 VTAIL.n379 VSUBS 0.027222f
C1696 VTAIL.n380 VSUBS 0.027222f
C1697 VTAIL.n381 VSUBS 0.014628f
C1698 VTAIL.n382 VSUBS 0.015488f
C1699 VTAIL.n383 VSUBS 0.034575f
C1700 VTAIL.n384 VSUBS 0.034575f
C1701 VTAIL.n385 VSUBS 0.015488f
C1702 VTAIL.n386 VSUBS 0.014628f
C1703 VTAIL.n387 VSUBS 0.027222f
C1704 VTAIL.n388 VSUBS 0.027222f
C1705 VTAIL.n389 VSUBS 0.014628f
C1706 VTAIL.n390 VSUBS 0.014628f
C1707 VTAIL.n391 VSUBS 0.015488f
C1708 VTAIL.n392 VSUBS 0.034575f
C1709 VTAIL.n393 VSUBS 0.034575f
C1710 VTAIL.n394 VSUBS 0.034575f
C1711 VTAIL.n395 VSUBS 0.015058f
C1712 VTAIL.n396 VSUBS 0.014628f
C1713 VTAIL.n397 VSUBS 0.027222f
C1714 VTAIL.n398 VSUBS 0.027222f
C1715 VTAIL.n399 VSUBS 0.014628f
C1716 VTAIL.n400 VSUBS 0.015488f
C1717 VTAIL.n401 VSUBS 0.034575f
C1718 VTAIL.n402 VSUBS 0.034575f
C1719 VTAIL.n403 VSUBS 0.015488f
C1720 VTAIL.n404 VSUBS 0.014628f
C1721 VTAIL.n405 VSUBS 0.027222f
C1722 VTAIL.n406 VSUBS 0.027222f
C1723 VTAIL.n407 VSUBS 0.014628f
C1724 VTAIL.n408 VSUBS 0.015488f
C1725 VTAIL.n409 VSUBS 0.034575f
C1726 VTAIL.n410 VSUBS 0.085279f
C1727 VTAIL.n411 VSUBS 0.015488f
C1728 VTAIL.n412 VSUBS 0.014628f
C1729 VTAIL.n413 VSUBS 0.064781f
C1730 VTAIL.n414 VSUBS 0.043012f
C1731 VTAIL.n415 VSUBS 2.05383f
C1732 VN.n0 VSUBS 0.033804f
C1733 VN.t4 VSUBS 3.06201f
C1734 VN.n1 VSUBS 0.029209f
C1735 VN.t1 VSUBS 3.22073f
C1736 VN.n2 VSUBS 1.14198f
C1737 VN.t3 VSUBS 3.06201f
C1738 VN.n3 VSUBS 1.16213f
C1739 VN.n4 VSUBS 0.068305f
C1740 VN.n5 VSUBS 0.250252f
C1741 VN.n6 VSUBS 0.033804f
C1742 VN.n7 VSUBS 0.033804f
C1743 VN.n8 VSUBS 0.06419f
C1744 VN.n9 VSUBS 0.039985f
C1745 VN.n10 VSUBS 1.15142f
C1746 VN.n11 VSUBS 0.035255f
C1747 VN.n12 VSUBS 0.033804f
C1748 VN.t0 VSUBS 3.06201f
C1749 VN.n13 VSUBS 0.029209f
C1750 VN.t2 VSUBS 3.22073f
C1751 VN.n14 VSUBS 1.14198f
C1752 VN.t5 VSUBS 3.06201f
C1753 VN.n15 VSUBS 1.16213f
C1754 VN.n16 VSUBS 0.068305f
C1755 VN.n17 VSUBS 0.250252f
C1756 VN.n18 VSUBS 0.033804f
C1757 VN.n19 VSUBS 0.033804f
C1758 VN.n20 VSUBS 0.06419f
C1759 VN.n21 VSUBS 0.039985f
C1760 VN.n22 VSUBS 1.15142f
C1761 VN.n23 VSUBS 1.88248f
.ends

