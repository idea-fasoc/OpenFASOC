* NGSPICE file created from diff_pair_sample_1207.ext - technology: sky130A

.subckt diff_pair_sample_1207 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t19 VP.t0 VDD1.t1 B.t7 sky130_fd_pr__nfet_01v8 ad=2.0163 pd=12.55 as=2.0163 ps=12.55 w=12.22 l=2.4
X1 VDD2.t9 VN.t0 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.0163 pd=12.55 as=2.0163 ps=12.55 w=12.22 l=2.4
X2 VDD1.t0 VP.t1 VTAIL.t18 B.t3 sky130_fd_pr__nfet_01v8 ad=2.0163 pd=12.55 as=4.7658 ps=25.22 w=12.22 l=2.4
X3 VTAIL.t17 VP.t2 VDD1.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=2.0163 pd=12.55 as=2.0163 ps=12.55 w=12.22 l=2.4
X4 VDD1.t2 VP.t3 VTAIL.t16 B.t4 sky130_fd_pr__nfet_01v8 ad=4.7658 pd=25.22 as=2.0163 ps=12.55 w=12.22 l=2.4
X5 VTAIL.t15 VP.t4 VDD1.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=2.0163 pd=12.55 as=2.0163 ps=12.55 w=12.22 l=2.4
X6 VDD2.t8 VN.t1 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=4.7658 pd=25.22 as=2.0163 ps=12.55 w=12.22 l=2.4
X7 B.t23 B.t21 B.t22 B.t15 sky130_fd_pr__nfet_01v8 ad=4.7658 pd=25.22 as=0 ps=0 w=12.22 l=2.4
X8 VTAIL.t7 VN.t2 VDD2.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=2.0163 pd=12.55 as=2.0163 ps=12.55 w=12.22 l=2.4
X9 VTAIL.t9 VN.t3 VDD2.t6 B.t9 sky130_fd_pr__nfet_01v8 ad=2.0163 pd=12.55 as=2.0163 ps=12.55 w=12.22 l=2.4
X10 VDD2.t5 VN.t4 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=4.7658 pd=25.22 as=2.0163 ps=12.55 w=12.22 l=2.4
X11 B.t20 B.t18 B.t19 B.t11 sky130_fd_pr__nfet_01v8 ad=4.7658 pd=25.22 as=0 ps=0 w=12.22 l=2.4
X12 VDD2.t4 VN.t5 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.0163 pd=12.55 as=4.7658 ps=25.22 w=12.22 l=2.4
X13 VDD1.t4 VP.t5 VTAIL.t14 B.t2 sky130_fd_pr__nfet_01v8 ad=2.0163 pd=12.55 as=2.0163 ps=12.55 w=12.22 l=2.4
X14 VDD1.t9 VP.t6 VTAIL.t13 B.t6 sky130_fd_pr__nfet_01v8 ad=4.7658 pd=25.22 as=2.0163 ps=12.55 w=12.22 l=2.4
X15 VTAIL.t1 VN.t6 VDD2.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=2.0163 pd=12.55 as=2.0163 ps=12.55 w=12.22 l=2.4
X16 VDD2.t2 VN.t7 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.0163 pd=12.55 as=4.7658 ps=25.22 w=12.22 l=2.4
X17 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=4.7658 pd=25.22 as=0 ps=0 w=12.22 l=2.4
X18 VTAIL.t0 VN.t8 VDD2.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=2.0163 pd=12.55 as=2.0163 ps=12.55 w=12.22 l=2.4
X19 VDD1.t8 VP.t7 VTAIL.t12 B.t8 sky130_fd_pr__nfet_01v8 ad=2.0163 pd=12.55 as=2.0163 ps=12.55 w=12.22 l=2.4
X20 VTAIL.t11 VP.t8 VDD1.t7 B.t9 sky130_fd_pr__nfet_01v8 ad=2.0163 pd=12.55 as=2.0163 ps=12.55 w=12.22 l=2.4
X21 VDD1.t6 VP.t9 VTAIL.t10 B.t5 sky130_fd_pr__nfet_01v8 ad=2.0163 pd=12.55 as=4.7658 ps=25.22 w=12.22 l=2.4
X22 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=4.7658 pd=25.22 as=0 ps=0 w=12.22 l=2.4
X23 VDD2.t0 VN.t9 VTAIL.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=2.0163 pd=12.55 as=2.0163 ps=12.55 w=12.22 l=2.4
R0 VP.n23 VP.n20 161.3
R1 VP.n25 VP.n24 161.3
R2 VP.n26 VP.n19 161.3
R3 VP.n28 VP.n27 161.3
R4 VP.n29 VP.n18 161.3
R5 VP.n32 VP.n31 161.3
R6 VP.n33 VP.n17 161.3
R7 VP.n35 VP.n34 161.3
R8 VP.n36 VP.n16 161.3
R9 VP.n38 VP.n37 161.3
R10 VP.n40 VP.n39 161.3
R11 VP.n41 VP.n14 161.3
R12 VP.n43 VP.n42 161.3
R13 VP.n44 VP.n13 161.3
R14 VP.n46 VP.n45 161.3
R15 VP.n47 VP.n12 161.3
R16 VP.n86 VP.n0 161.3
R17 VP.n85 VP.n84 161.3
R18 VP.n83 VP.n1 161.3
R19 VP.n82 VP.n81 161.3
R20 VP.n80 VP.n2 161.3
R21 VP.n79 VP.n78 161.3
R22 VP.n77 VP.n76 161.3
R23 VP.n75 VP.n4 161.3
R24 VP.n74 VP.n73 161.3
R25 VP.n72 VP.n5 161.3
R26 VP.n71 VP.n70 161.3
R27 VP.n68 VP.n6 161.3
R28 VP.n67 VP.n66 161.3
R29 VP.n65 VP.n7 161.3
R30 VP.n64 VP.n63 161.3
R31 VP.n62 VP.n8 161.3
R32 VP.n60 VP.n59 161.3
R33 VP.n58 VP.n9 161.3
R34 VP.n57 VP.n56 161.3
R35 VP.n55 VP.n10 161.3
R36 VP.n54 VP.n53 161.3
R37 VP.n52 VP.n11 161.3
R38 VP.n21 VP.t6 156.357
R39 VP.n50 VP.t3 122.71
R40 VP.n61 VP.t2 122.71
R41 VP.n69 VP.t5 122.71
R42 VP.n3 VP.t8 122.71
R43 VP.n87 VP.t1 122.71
R44 VP.n48 VP.t9 122.71
R45 VP.n15 VP.t4 122.71
R46 VP.n30 VP.t7 122.71
R47 VP.n22 VP.t0 122.71
R48 VP.n51 VP.n50 100.382
R49 VP.n88 VP.n87 100.382
R50 VP.n49 VP.n48 100.382
R51 VP.n56 VP.n55 55.5035
R52 VP.n81 VP.n1 55.5035
R53 VP.n42 VP.n13 55.5035
R54 VP.n51 VP.n49 52.17
R55 VP.n63 VP.n7 51.6086
R56 VP.n75 VP.n74 51.6086
R57 VP.n36 VP.n35 51.6086
R58 VP.n24 VP.n19 51.6086
R59 VP.n22 VP.n21 48.8439
R60 VP.n67 VP.n7 29.2126
R61 VP.n74 VP.n5 29.2126
R62 VP.n35 VP.n17 29.2126
R63 VP.n28 VP.n19 29.2126
R64 VP.n55 VP.n54 25.3177
R65 VP.n85 VP.n1 25.3177
R66 VP.n46 VP.n13 25.3177
R67 VP.n54 VP.n11 24.3439
R68 VP.n56 VP.n9 24.3439
R69 VP.n60 VP.n9 24.3439
R70 VP.n63 VP.n62 24.3439
R71 VP.n68 VP.n67 24.3439
R72 VP.n70 VP.n5 24.3439
R73 VP.n76 VP.n75 24.3439
R74 VP.n80 VP.n79 24.3439
R75 VP.n81 VP.n80 24.3439
R76 VP.n86 VP.n85 24.3439
R77 VP.n47 VP.n46 24.3439
R78 VP.n37 VP.n36 24.3439
R79 VP.n41 VP.n40 24.3439
R80 VP.n42 VP.n41 24.3439
R81 VP.n29 VP.n28 24.3439
R82 VP.n31 VP.n17 24.3439
R83 VP.n24 VP.n23 24.3439
R84 VP.n62 VP.n61 23.3702
R85 VP.n76 VP.n3 23.3702
R86 VP.n37 VP.n15 23.3702
R87 VP.n23 VP.n22 23.3702
R88 VP.n69 VP.n68 12.1722
R89 VP.n70 VP.n69 12.1722
R90 VP.n30 VP.n29 12.1722
R91 VP.n31 VP.n30 12.1722
R92 VP.n50 VP.n11 10.2247
R93 VP.n87 VP.n86 10.2247
R94 VP.n48 VP.n47 10.2247
R95 VP.n21 VP.n20 6.8468
R96 VP.n61 VP.n60 0.974237
R97 VP.n79 VP.n3 0.974237
R98 VP.n40 VP.n15 0.974237
R99 VP.n49 VP.n12 0.278398
R100 VP.n52 VP.n51 0.278398
R101 VP.n88 VP.n0 0.278398
R102 VP.n25 VP.n20 0.189894
R103 VP.n26 VP.n25 0.189894
R104 VP.n27 VP.n26 0.189894
R105 VP.n27 VP.n18 0.189894
R106 VP.n32 VP.n18 0.189894
R107 VP.n33 VP.n32 0.189894
R108 VP.n34 VP.n33 0.189894
R109 VP.n34 VP.n16 0.189894
R110 VP.n38 VP.n16 0.189894
R111 VP.n39 VP.n38 0.189894
R112 VP.n39 VP.n14 0.189894
R113 VP.n43 VP.n14 0.189894
R114 VP.n44 VP.n43 0.189894
R115 VP.n45 VP.n44 0.189894
R116 VP.n45 VP.n12 0.189894
R117 VP.n53 VP.n52 0.189894
R118 VP.n53 VP.n10 0.189894
R119 VP.n57 VP.n10 0.189894
R120 VP.n58 VP.n57 0.189894
R121 VP.n59 VP.n58 0.189894
R122 VP.n59 VP.n8 0.189894
R123 VP.n64 VP.n8 0.189894
R124 VP.n65 VP.n64 0.189894
R125 VP.n66 VP.n65 0.189894
R126 VP.n66 VP.n6 0.189894
R127 VP.n71 VP.n6 0.189894
R128 VP.n72 VP.n71 0.189894
R129 VP.n73 VP.n72 0.189894
R130 VP.n73 VP.n4 0.189894
R131 VP.n77 VP.n4 0.189894
R132 VP.n78 VP.n77 0.189894
R133 VP.n78 VP.n2 0.189894
R134 VP.n82 VP.n2 0.189894
R135 VP.n83 VP.n82 0.189894
R136 VP.n84 VP.n83 0.189894
R137 VP.n84 VP.n0 0.189894
R138 VP VP.n88 0.153422
R139 VDD1.n60 VDD1.n0 289.615
R140 VDD1.n127 VDD1.n67 289.615
R141 VDD1.n61 VDD1.n60 185
R142 VDD1.n59 VDD1.n58 185
R143 VDD1.n4 VDD1.n3 185
R144 VDD1.n53 VDD1.n52 185
R145 VDD1.n51 VDD1.n50 185
R146 VDD1.n8 VDD1.n7 185
R147 VDD1.n45 VDD1.n44 185
R148 VDD1.n43 VDD1.n10 185
R149 VDD1.n42 VDD1.n41 185
R150 VDD1.n13 VDD1.n11 185
R151 VDD1.n36 VDD1.n35 185
R152 VDD1.n34 VDD1.n33 185
R153 VDD1.n17 VDD1.n16 185
R154 VDD1.n28 VDD1.n27 185
R155 VDD1.n26 VDD1.n25 185
R156 VDD1.n21 VDD1.n20 185
R157 VDD1.n87 VDD1.n86 185
R158 VDD1.n92 VDD1.n91 185
R159 VDD1.n94 VDD1.n93 185
R160 VDD1.n83 VDD1.n82 185
R161 VDD1.n100 VDD1.n99 185
R162 VDD1.n102 VDD1.n101 185
R163 VDD1.n79 VDD1.n78 185
R164 VDD1.n109 VDD1.n108 185
R165 VDD1.n110 VDD1.n77 185
R166 VDD1.n112 VDD1.n111 185
R167 VDD1.n75 VDD1.n74 185
R168 VDD1.n118 VDD1.n117 185
R169 VDD1.n120 VDD1.n119 185
R170 VDD1.n71 VDD1.n70 185
R171 VDD1.n126 VDD1.n125 185
R172 VDD1.n128 VDD1.n127 185
R173 VDD1.n22 VDD1.t9 149.524
R174 VDD1.n88 VDD1.t2 149.524
R175 VDD1.n60 VDD1.n59 104.615
R176 VDD1.n59 VDD1.n3 104.615
R177 VDD1.n52 VDD1.n3 104.615
R178 VDD1.n52 VDD1.n51 104.615
R179 VDD1.n51 VDD1.n7 104.615
R180 VDD1.n44 VDD1.n7 104.615
R181 VDD1.n44 VDD1.n43 104.615
R182 VDD1.n43 VDD1.n42 104.615
R183 VDD1.n42 VDD1.n11 104.615
R184 VDD1.n35 VDD1.n11 104.615
R185 VDD1.n35 VDD1.n34 104.615
R186 VDD1.n34 VDD1.n16 104.615
R187 VDD1.n27 VDD1.n16 104.615
R188 VDD1.n27 VDD1.n26 104.615
R189 VDD1.n26 VDD1.n20 104.615
R190 VDD1.n92 VDD1.n86 104.615
R191 VDD1.n93 VDD1.n92 104.615
R192 VDD1.n93 VDD1.n82 104.615
R193 VDD1.n100 VDD1.n82 104.615
R194 VDD1.n101 VDD1.n100 104.615
R195 VDD1.n101 VDD1.n78 104.615
R196 VDD1.n109 VDD1.n78 104.615
R197 VDD1.n110 VDD1.n109 104.615
R198 VDD1.n111 VDD1.n110 104.615
R199 VDD1.n111 VDD1.n74 104.615
R200 VDD1.n118 VDD1.n74 104.615
R201 VDD1.n119 VDD1.n118 104.615
R202 VDD1.n119 VDD1.n70 104.615
R203 VDD1.n126 VDD1.n70 104.615
R204 VDD1.n127 VDD1.n126 104.615
R205 VDD1.n135 VDD1.n134 65.5289
R206 VDD1.n66 VDD1.n65 63.8193
R207 VDD1.n137 VDD1.n136 63.8192
R208 VDD1.n133 VDD1.n132 63.8192
R209 VDD1.n66 VDD1.n64 53.157
R210 VDD1.n133 VDD1.n131 53.157
R211 VDD1.t9 VDD1.n20 52.3082
R212 VDD1.t2 VDD1.n86 52.3082
R213 VDD1.n137 VDD1.n135 47.1884
R214 VDD1.n45 VDD1.n10 13.1884
R215 VDD1.n112 VDD1.n77 13.1884
R216 VDD1.n46 VDD1.n8 12.8005
R217 VDD1.n41 VDD1.n12 12.8005
R218 VDD1.n108 VDD1.n107 12.8005
R219 VDD1.n113 VDD1.n75 12.8005
R220 VDD1.n50 VDD1.n49 12.0247
R221 VDD1.n40 VDD1.n13 12.0247
R222 VDD1.n106 VDD1.n79 12.0247
R223 VDD1.n117 VDD1.n116 12.0247
R224 VDD1.n53 VDD1.n6 11.249
R225 VDD1.n37 VDD1.n36 11.249
R226 VDD1.n103 VDD1.n102 11.249
R227 VDD1.n120 VDD1.n73 11.249
R228 VDD1.n54 VDD1.n4 10.4732
R229 VDD1.n33 VDD1.n15 10.4732
R230 VDD1.n99 VDD1.n81 10.4732
R231 VDD1.n121 VDD1.n71 10.4732
R232 VDD1.n22 VDD1.n21 10.2747
R233 VDD1.n88 VDD1.n87 10.2747
R234 VDD1.n58 VDD1.n57 9.69747
R235 VDD1.n32 VDD1.n17 9.69747
R236 VDD1.n98 VDD1.n83 9.69747
R237 VDD1.n125 VDD1.n124 9.69747
R238 VDD1.n64 VDD1.n63 9.45567
R239 VDD1.n131 VDD1.n130 9.45567
R240 VDD1.n24 VDD1.n23 9.3005
R241 VDD1.n19 VDD1.n18 9.3005
R242 VDD1.n30 VDD1.n29 9.3005
R243 VDD1.n32 VDD1.n31 9.3005
R244 VDD1.n15 VDD1.n14 9.3005
R245 VDD1.n38 VDD1.n37 9.3005
R246 VDD1.n40 VDD1.n39 9.3005
R247 VDD1.n12 VDD1.n9 9.3005
R248 VDD1.n63 VDD1.n62 9.3005
R249 VDD1.n2 VDD1.n1 9.3005
R250 VDD1.n57 VDD1.n56 9.3005
R251 VDD1.n55 VDD1.n54 9.3005
R252 VDD1.n6 VDD1.n5 9.3005
R253 VDD1.n49 VDD1.n48 9.3005
R254 VDD1.n47 VDD1.n46 9.3005
R255 VDD1.n130 VDD1.n129 9.3005
R256 VDD1.n69 VDD1.n68 9.3005
R257 VDD1.n124 VDD1.n123 9.3005
R258 VDD1.n122 VDD1.n121 9.3005
R259 VDD1.n73 VDD1.n72 9.3005
R260 VDD1.n116 VDD1.n115 9.3005
R261 VDD1.n114 VDD1.n113 9.3005
R262 VDD1.n90 VDD1.n89 9.3005
R263 VDD1.n85 VDD1.n84 9.3005
R264 VDD1.n96 VDD1.n95 9.3005
R265 VDD1.n98 VDD1.n97 9.3005
R266 VDD1.n81 VDD1.n80 9.3005
R267 VDD1.n104 VDD1.n103 9.3005
R268 VDD1.n106 VDD1.n105 9.3005
R269 VDD1.n107 VDD1.n76 9.3005
R270 VDD1.n61 VDD1.n2 8.92171
R271 VDD1.n29 VDD1.n28 8.92171
R272 VDD1.n95 VDD1.n94 8.92171
R273 VDD1.n128 VDD1.n69 8.92171
R274 VDD1.n62 VDD1.n0 8.14595
R275 VDD1.n25 VDD1.n19 8.14595
R276 VDD1.n91 VDD1.n85 8.14595
R277 VDD1.n129 VDD1.n67 8.14595
R278 VDD1.n24 VDD1.n21 7.3702
R279 VDD1.n90 VDD1.n87 7.3702
R280 VDD1.n64 VDD1.n0 5.81868
R281 VDD1.n25 VDD1.n24 5.81868
R282 VDD1.n91 VDD1.n90 5.81868
R283 VDD1.n131 VDD1.n67 5.81868
R284 VDD1.n62 VDD1.n61 5.04292
R285 VDD1.n28 VDD1.n19 5.04292
R286 VDD1.n94 VDD1.n85 5.04292
R287 VDD1.n129 VDD1.n128 5.04292
R288 VDD1.n58 VDD1.n2 4.26717
R289 VDD1.n29 VDD1.n17 4.26717
R290 VDD1.n95 VDD1.n83 4.26717
R291 VDD1.n125 VDD1.n69 4.26717
R292 VDD1.n57 VDD1.n4 3.49141
R293 VDD1.n33 VDD1.n32 3.49141
R294 VDD1.n99 VDD1.n98 3.49141
R295 VDD1.n124 VDD1.n71 3.49141
R296 VDD1.n23 VDD1.n22 2.84303
R297 VDD1.n89 VDD1.n88 2.84303
R298 VDD1.n54 VDD1.n53 2.71565
R299 VDD1.n36 VDD1.n15 2.71565
R300 VDD1.n102 VDD1.n81 2.71565
R301 VDD1.n121 VDD1.n120 2.71565
R302 VDD1.n50 VDD1.n6 1.93989
R303 VDD1.n37 VDD1.n13 1.93989
R304 VDD1.n103 VDD1.n79 1.93989
R305 VDD1.n117 VDD1.n73 1.93989
R306 VDD1 VDD1.n137 1.7074
R307 VDD1.n136 VDD1.t5 1.62079
R308 VDD1.n136 VDD1.t6 1.62079
R309 VDD1.n65 VDD1.t1 1.62079
R310 VDD1.n65 VDD1.t8 1.62079
R311 VDD1.n134 VDD1.t7 1.62079
R312 VDD1.n134 VDD1.t0 1.62079
R313 VDD1.n132 VDD1.t3 1.62079
R314 VDD1.n132 VDD1.t4 1.62079
R315 VDD1.n49 VDD1.n8 1.16414
R316 VDD1.n41 VDD1.n40 1.16414
R317 VDD1.n108 VDD1.n106 1.16414
R318 VDD1.n116 VDD1.n75 1.16414
R319 VDD1 VDD1.n66 0.647052
R320 VDD1.n135 VDD1.n133 0.533516
R321 VDD1.n46 VDD1.n45 0.388379
R322 VDD1.n12 VDD1.n10 0.388379
R323 VDD1.n107 VDD1.n77 0.388379
R324 VDD1.n113 VDD1.n112 0.388379
R325 VDD1.n63 VDD1.n1 0.155672
R326 VDD1.n56 VDD1.n1 0.155672
R327 VDD1.n56 VDD1.n55 0.155672
R328 VDD1.n55 VDD1.n5 0.155672
R329 VDD1.n48 VDD1.n5 0.155672
R330 VDD1.n48 VDD1.n47 0.155672
R331 VDD1.n47 VDD1.n9 0.155672
R332 VDD1.n39 VDD1.n9 0.155672
R333 VDD1.n39 VDD1.n38 0.155672
R334 VDD1.n38 VDD1.n14 0.155672
R335 VDD1.n31 VDD1.n14 0.155672
R336 VDD1.n31 VDD1.n30 0.155672
R337 VDD1.n30 VDD1.n18 0.155672
R338 VDD1.n23 VDD1.n18 0.155672
R339 VDD1.n89 VDD1.n84 0.155672
R340 VDD1.n96 VDD1.n84 0.155672
R341 VDD1.n97 VDD1.n96 0.155672
R342 VDD1.n97 VDD1.n80 0.155672
R343 VDD1.n104 VDD1.n80 0.155672
R344 VDD1.n105 VDD1.n104 0.155672
R345 VDD1.n105 VDD1.n76 0.155672
R346 VDD1.n114 VDD1.n76 0.155672
R347 VDD1.n115 VDD1.n114 0.155672
R348 VDD1.n115 VDD1.n72 0.155672
R349 VDD1.n122 VDD1.n72 0.155672
R350 VDD1.n123 VDD1.n122 0.155672
R351 VDD1.n123 VDD1.n68 0.155672
R352 VDD1.n130 VDD1.n68 0.155672
R353 VTAIL.n272 VTAIL.n212 289.615
R354 VTAIL.n62 VTAIL.n2 289.615
R355 VTAIL.n206 VTAIL.n146 289.615
R356 VTAIL.n136 VTAIL.n76 289.615
R357 VTAIL.n232 VTAIL.n231 185
R358 VTAIL.n237 VTAIL.n236 185
R359 VTAIL.n239 VTAIL.n238 185
R360 VTAIL.n228 VTAIL.n227 185
R361 VTAIL.n245 VTAIL.n244 185
R362 VTAIL.n247 VTAIL.n246 185
R363 VTAIL.n224 VTAIL.n223 185
R364 VTAIL.n254 VTAIL.n253 185
R365 VTAIL.n255 VTAIL.n222 185
R366 VTAIL.n257 VTAIL.n256 185
R367 VTAIL.n220 VTAIL.n219 185
R368 VTAIL.n263 VTAIL.n262 185
R369 VTAIL.n265 VTAIL.n264 185
R370 VTAIL.n216 VTAIL.n215 185
R371 VTAIL.n271 VTAIL.n270 185
R372 VTAIL.n273 VTAIL.n272 185
R373 VTAIL.n22 VTAIL.n21 185
R374 VTAIL.n27 VTAIL.n26 185
R375 VTAIL.n29 VTAIL.n28 185
R376 VTAIL.n18 VTAIL.n17 185
R377 VTAIL.n35 VTAIL.n34 185
R378 VTAIL.n37 VTAIL.n36 185
R379 VTAIL.n14 VTAIL.n13 185
R380 VTAIL.n44 VTAIL.n43 185
R381 VTAIL.n45 VTAIL.n12 185
R382 VTAIL.n47 VTAIL.n46 185
R383 VTAIL.n10 VTAIL.n9 185
R384 VTAIL.n53 VTAIL.n52 185
R385 VTAIL.n55 VTAIL.n54 185
R386 VTAIL.n6 VTAIL.n5 185
R387 VTAIL.n61 VTAIL.n60 185
R388 VTAIL.n63 VTAIL.n62 185
R389 VTAIL.n207 VTAIL.n206 185
R390 VTAIL.n205 VTAIL.n204 185
R391 VTAIL.n150 VTAIL.n149 185
R392 VTAIL.n199 VTAIL.n198 185
R393 VTAIL.n197 VTAIL.n196 185
R394 VTAIL.n154 VTAIL.n153 185
R395 VTAIL.n191 VTAIL.n190 185
R396 VTAIL.n189 VTAIL.n156 185
R397 VTAIL.n188 VTAIL.n187 185
R398 VTAIL.n159 VTAIL.n157 185
R399 VTAIL.n182 VTAIL.n181 185
R400 VTAIL.n180 VTAIL.n179 185
R401 VTAIL.n163 VTAIL.n162 185
R402 VTAIL.n174 VTAIL.n173 185
R403 VTAIL.n172 VTAIL.n171 185
R404 VTAIL.n167 VTAIL.n166 185
R405 VTAIL.n137 VTAIL.n136 185
R406 VTAIL.n135 VTAIL.n134 185
R407 VTAIL.n80 VTAIL.n79 185
R408 VTAIL.n129 VTAIL.n128 185
R409 VTAIL.n127 VTAIL.n126 185
R410 VTAIL.n84 VTAIL.n83 185
R411 VTAIL.n121 VTAIL.n120 185
R412 VTAIL.n119 VTAIL.n86 185
R413 VTAIL.n118 VTAIL.n117 185
R414 VTAIL.n89 VTAIL.n87 185
R415 VTAIL.n112 VTAIL.n111 185
R416 VTAIL.n110 VTAIL.n109 185
R417 VTAIL.n93 VTAIL.n92 185
R418 VTAIL.n104 VTAIL.n103 185
R419 VTAIL.n102 VTAIL.n101 185
R420 VTAIL.n97 VTAIL.n96 185
R421 VTAIL.n233 VTAIL.t5 149.524
R422 VTAIL.n23 VTAIL.t18 149.524
R423 VTAIL.n168 VTAIL.t10 149.524
R424 VTAIL.n98 VTAIL.t3 149.524
R425 VTAIL.n237 VTAIL.n231 104.615
R426 VTAIL.n238 VTAIL.n237 104.615
R427 VTAIL.n238 VTAIL.n227 104.615
R428 VTAIL.n245 VTAIL.n227 104.615
R429 VTAIL.n246 VTAIL.n245 104.615
R430 VTAIL.n246 VTAIL.n223 104.615
R431 VTAIL.n254 VTAIL.n223 104.615
R432 VTAIL.n255 VTAIL.n254 104.615
R433 VTAIL.n256 VTAIL.n255 104.615
R434 VTAIL.n256 VTAIL.n219 104.615
R435 VTAIL.n263 VTAIL.n219 104.615
R436 VTAIL.n264 VTAIL.n263 104.615
R437 VTAIL.n264 VTAIL.n215 104.615
R438 VTAIL.n271 VTAIL.n215 104.615
R439 VTAIL.n272 VTAIL.n271 104.615
R440 VTAIL.n27 VTAIL.n21 104.615
R441 VTAIL.n28 VTAIL.n27 104.615
R442 VTAIL.n28 VTAIL.n17 104.615
R443 VTAIL.n35 VTAIL.n17 104.615
R444 VTAIL.n36 VTAIL.n35 104.615
R445 VTAIL.n36 VTAIL.n13 104.615
R446 VTAIL.n44 VTAIL.n13 104.615
R447 VTAIL.n45 VTAIL.n44 104.615
R448 VTAIL.n46 VTAIL.n45 104.615
R449 VTAIL.n46 VTAIL.n9 104.615
R450 VTAIL.n53 VTAIL.n9 104.615
R451 VTAIL.n54 VTAIL.n53 104.615
R452 VTAIL.n54 VTAIL.n5 104.615
R453 VTAIL.n61 VTAIL.n5 104.615
R454 VTAIL.n62 VTAIL.n61 104.615
R455 VTAIL.n206 VTAIL.n205 104.615
R456 VTAIL.n205 VTAIL.n149 104.615
R457 VTAIL.n198 VTAIL.n149 104.615
R458 VTAIL.n198 VTAIL.n197 104.615
R459 VTAIL.n197 VTAIL.n153 104.615
R460 VTAIL.n190 VTAIL.n153 104.615
R461 VTAIL.n190 VTAIL.n189 104.615
R462 VTAIL.n189 VTAIL.n188 104.615
R463 VTAIL.n188 VTAIL.n157 104.615
R464 VTAIL.n181 VTAIL.n157 104.615
R465 VTAIL.n181 VTAIL.n180 104.615
R466 VTAIL.n180 VTAIL.n162 104.615
R467 VTAIL.n173 VTAIL.n162 104.615
R468 VTAIL.n173 VTAIL.n172 104.615
R469 VTAIL.n172 VTAIL.n166 104.615
R470 VTAIL.n136 VTAIL.n135 104.615
R471 VTAIL.n135 VTAIL.n79 104.615
R472 VTAIL.n128 VTAIL.n79 104.615
R473 VTAIL.n128 VTAIL.n127 104.615
R474 VTAIL.n127 VTAIL.n83 104.615
R475 VTAIL.n120 VTAIL.n83 104.615
R476 VTAIL.n120 VTAIL.n119 104.615
R477 VTAIL.n119 VTAIL.n118 104.615
R478 VTAIL.n118 VTAIL.n87 104.615
R479 VTAIL.n111 VTAIL.n87 104.615
R480 VTAIL.n111 VTAIL.n110 104.615
R481 VTAIL.n110 VTAIL.n92 104.615
R482 VTAIL.n103 VTAIL.n92 104.615
R483 VTAIL.n103 VTAIL.n102 104.615
R484 VTAIL.n102 VTAIL.n96 104.615
R485 VTAIL.t5 VTAIL.n231 52.3082
R486 VTAIL.t18 VTAIL.n21 52.3082
R487 VTAIL.t10 VTAIL.n166 52.3082
R488 VTAIL.t3 VTAIL.n96 52.3082
R489 VTAIL.n145 VTAIL.n144 47.1406
R490 VTAIL.n143 VTAIL.n142 47.1406
R491 VTAIL.n75 VTAIL.n74 47.1406
R492 VTAIL.n73 VTAIL.n72 47.1406
R493 VTAIL.n279 VTAIL.n278 47.1404
R494 VTAIL.n1 VTAIL.n0 47.1404
R495 VTAIL.n69 VTAIL.n68 47.1404
R496 VTAIL.n71 VTAIL.n70 47.1404
R497 VTAIL.n277 VTAIL.n276 34.1247
R498 VTAIL.n67 VTAIL.n66 34.1247
R499 VTAIL.n211 VTAIL.n210 34.1247
R500 VTAIL.n141 VTAIL.n140 34.1247
R501 VTAIL.n73 VTAIL.n71 27.6083
R502 VTAIL.n277 VTAIL.n211 25.2548
R503 VTAIL.n257 VTAIL.n222 13.1884
R504 VTAIL.n47 VTAIL.n12 13.1884
R505 VTAIL.n191 VTAIL.n156 13.1884
R506 VTAIL.n121 VTAIL.n86 13.1884
R507 VTAIL.n253 VTAIL.n252 12.8005
R508 VTAIL.n258 VTAIL.n220 12.8005
R509 VTAIL.n43 VTAIL.n42 12.8005
R510 VTAIL.n48 VTAIL.n10 12.8005
R511 VTAIL.n192 VTAIL.n154 12.8005
R512 VTAIL.n187 VTAIL.n158 12.8005
R513 VTAIL.n122 VTAIL.n84 12.8005
R514 VTAIL.n117 VTAIL.n88 12.8005
R515 VTAIL.n251 VTAIL.n224 12.0247
R516 VTAIL.n262 VTAIL.n261 12.0247
R517 VTAIL.n41 VTAIL.n14 12.0247
R518 VTAIL.n52 VTAIL.n51 12.0247
R519 VTAIL.n196 VTAIL.n195 12.0247
R520 VTAIL.n186 VTAIL.n159 12.0247
R521 VTAIL.n126 VTAIL.n125 12.0247
R522 VTAIL.n116 VTAIL.n89 12.0247
R523 VTAIL.n248 VTAIL.n247 11.249
R524 VTAIL.n265 VTAIL.n218 11.249
R525 VTAIL.n38 VTAIL.n37 11.249
R526 VTAIL.n55 VTAIL.n8 11.249
R527 VTAIL.n199 VTAIL.n152 11.249
R528 VTAIL.n183 VTAIL.n182 11.249
R529 VTAIL.n129 VTAIL.n82 11.249
R530 VTAIL.n113 VTAIL.n112 11.249
R531 VTAIL.n244 VTAIL.n226 10.4732
R532 VTAIL.n266 VTAIL.n216 10.4732
R533 VTAIL.n34 VTAIL.n16 10.4732
R534 VTAIL.n56 VTAIL.n6 10.4732
R535 VTAIL.n200 VTAIL.n150 10.4732
R536 VTAIL.n179 VTAIL.n161 10.4732
R537 VTAIL.n130 VTAIL.n80 10.4732
R538 VTAIL.n109 VTAIL.n91 10.4732
R539 VTAIL.n233 VTAIL.n232 10.2747
R540 VTAIL.n23 VTAIL.n22 10.2747
R541 VTAIL.n168 VTAIL.n167 10.2747
R542 VTAIL.n98 VTAIL.n97 10.2747
R543 VTAIL.n243 VTAIL.n228 9.69747
R544 VTAIL.n270 VTAIL.n269 9.69747
R545 VTAIL.n33 VTAIL.n18 9.69747
R546 VTAIL.n60 VTAIL.n59 9.69747
R547 VTAIL.n204 VTAIL.n203 9.69747
R548 VTAIL.n178 VTAIL.n163 9.69747
R549 VTAIL.n134 VTAIL.n133 9.69747
R550 VTAIL.n108 VTAIL.n93 9.69747
R551 VTAIL.n276 VTAIL.n275 9.45567
R552 VTAIL.n66 VTAIL.n65 9.45567
R553 VTAIL.n210 VTAIL.n209 9.45567
R554 VTAIL.n140 VTAIL.n139 9.45567
R555 VTAIL.n275 VTAIL.n274 9.3005
R556 VTAIL.n214 VTAIL.n213 9.3005
R557 VTAIL.n269 VTAIL.n268 9.3005
R558 VTAIL.n267 VTAIL.n266 9.3005
R559 VTAIL.n218 VTAIL.n217 9.3005
R560 VTAIL.n261 VTAIL.n260 9.3005
R561 VTAIL.n259 VTAIL.n258 9.3005
R562 VTAIL.n235 VTAIL.n234 9.3005
R563 VTAIL.n230 VTAIL.n229 9.3005
R564 VTAIL.n241 VTAIL.n240 9.3005
R565 VTAIL.n243 VTAIL.n242 9.3005
R566 VTAIL.n226 VTAIL.n225 9.3005
R567 VTAIL.n249 VTAIL.n248 9.3005
R568 VTAIL.n251 VTAIL.n250 9.3005
R569 VTAIL.n252 VTAIL.n221 9.3005
R570 VTAIL.n65 VTAIL.n64 9.3005
R571 VTAIL.n4 VTAIL.n3 9.3005
R572 VTAIL.n59 VTAIL.n58 9.3005
R573 VTAIL.n57 VTAIL.n56 9.3005
R574 VTAIL.n8 VTAIL.n7 9.3005
R575 VTAIL.n51 VTAIL.n50 9.3005
R576 VTAIL.n49 VTAIL.n48 9.3005
R577 VTAIL.n25 VTAIL.n24 9.3005
R578 VTAIL.n20 VTAIL.n19 9.3005
R579 VTAIL.n31 VTAIL.n30 9.3005
R580 VTAIL.n33 VTAIL.n32 9.3005
R581 VTAIL.n16 VTAIL.n15 9.3005
R582 VTAIL.n39 VTAIL.n38 9.3005
R583 VTAIL.n41 VTAIL.n40 9.3005
R584 VTAIL.n42 VTAIL.n11 9.3005
R585 VTAIL.n170 VTAIL.n169 9.3005
R586 VTAIL.n165 VTAIL.n164 9.3005
R587 VTAIL.n176 VTAIL.n175 9.3005
R588 VTAIL.n178 VTAIL.n177 9.3005
R589 VTAIL.n161 VTAIL.n160 9.3005
R590 VTAIL.n184 VTAIL.n183 9.3005
R591 VTAIL.n186 VTAIL.n185 9.3005
R592 VTAIL.n158 VTAIL.n155 9.3005
R593 VTAIL.n209 VTAIL.n208 9.3005
R594 VTAIL.n148 VTAIL.n147 9.3005
R595 VTAIL.n203 VTAIL.n202 9.3005
R596 VTAIL.n201 VTAIL.n200 9.3005
R597 VTAIL.n152 VTAIL.n151 9.3005
R598 VTAIL.n195 VTAIL.n194 9.3005
R599 VTAIL.n193 VTAIL.n192 9.3005
R600 VTAIL.n100 VTAIL.n99 9.3005
R601 VTAIL.n95 VTAIL.n94 9.3005
R602 VTAIL.n106 VTAIL.n105 9.3005
R603 VTAIL.n108 VTAIL.n107 9.3005
R604 VTAIL.n91 VTAIL.n90 9.3005
R605 VTAIL.n114 VTAIL.n113 9.3005
R606 VTAIL.n116 VTAIL.n115 9.3005
R607 VTAIL.n88 VTAIL.n85 9.3005
R608 VTAIL.n139 VTAIL.n138 9.3005
R609 VTAIL.n78 VTAIL.n77 9.3005
R610 VTAIL.n133 VTAIL.n132 9.3005
R611 VTAIL.n131 VTAIL.n130 9.3005
R612 VTAIL.n82 VTAIL.n81 9.3005
R613 VTAIL.n125 VTAIL.n124 9.3005
R614 VTAIL.n123 VTAIL.n122 9.3005
R615 VTAIL.n240 VTAIL.n239 8.92171
R616 VTAIL.n273 VTAIL.n214 8.92171
R617 VTAIL.n30 VTAIL.n29 8.92171
R618 VTAIL.n63 VTAIL.n4 8.92171
R619 VTAIL.n207 VTAIL.n148 8.92171
R620 VTAIL.n175 VTAIL.n174 8.92171
R621 VTAIL.n137 VTAIL.n78 8.92171
R622 VTAIL.n105 VTAIL.n104 8.92171
R623 VTAIL.n236 VTAIL.n230 8.14595
R624 VTAIL.n274 VTAIL.n212 8.14595
R625 VTAIL.n26 VTAIL.n20 8.14595
R626 VTAIL.n64 VTAIL.n2 8.14595
R627 VTAIL.n208 VTAIL.n146 8.14595
R628 VTAIL.n171 VTAIL.n165 8.14595
R629 VTAIL.n138 VTAIL.n76 8.14595
R630 VTAIL.n101 VTAIL.n95 8.14595
R631 VTAIL.n235 VTAIL.n232 7.3702
R632 VTAIL.n25 VTAIL.n22 7.3702
R633 VTAIL.n170 VTAIL.n167 7.3702
R634 VTAIL.n100 VTAIL.n97 7.3702
R635 VTAIL.n236 VTAIL.n235 5.81868
R636 VTAIL.n276 VTAIL.n212 5.81868
R637 VTAIL.n26 VTAIL.n25 5.81868
R638 VTAIL.n66 VTAIL.n2 5.81868
R639 VTAIL.n210 VTAIL.n146 5.81868
R640 VTAIL.n171 VTAIL.n170 5.81868
R641 VTAIL.n140 VTAIL.n76 5.81868
R642 VTAIL.n101 VTAIL.n100 5.81868
R643 VTAIL.n239 VTAIL.n230 5.04292
R644 VTAIL.n274 VTAIL.n273 5.04292
R645 VTAIL.n29 VTAIL.n20 5.04292
R646 VTAIL.n64 VTAIL.n63 5.04292
R647 VTAIL.n208 VTAIL.n207 5.04292
R648 VTAIL.n174 VTAIL.n165 5.04292
R649 VTAIL.n138 VTAIL.n137 5.04292
R650 VTAIL.n104 VTAIL.n95 5.04292
R651 VTAIL.n240 VTAIL.n228 4.26717
R652 VTAIL.n270 VTAIL.n214 4.26717
R653 VTAIL.n30 VTAIL.n18 4.26717
R654 VTAIL.n60 VTAIL.n4 4.26717
R655 VTAIL.n204 VTAIL.n148 4.26717
R656 VTAIL.n175 VTAIL.n163 4.26717
R657 VTAIL.n134 VTAIL.n78 4.26717
R658 VTAIL.n105 VTAIL.n93 4.26717
R659 VTAIL.n244 VTAIL.n243 3.49141
R660 VTAIL.n269 VTAIL.n216 3.49141
R661 VTAIL.n34 VTAIL.n33 3.49141
R662 VTAIL.n59 VTAIL.n6 3.49141
R663 VTAIL.n203 VTAIL.n150 3.49141
R664 VTAIL.n179 VTAIL.n178 3.49141
R665 VTAIL.n133 VTAIL.n80 3.49141
R666 VTAIL.n109 VTAIL.n108 3.49141
R667 VTAIL.n234 VTAIL.n233 2.84303
R668 VTAIL.n24 VTAIL.n23 2.84303
R669 VTAIL.n169 VTAIL.n168 2.84303
R670 VTAIL.n99 VTAIL.n98 2.84303
R671 VTAIL.n247 VTAIL.n226 2.71565
R672 VTAIL.n266 VTAIL.n265 2.71565
R673 VTAIL.n37 VTAIL.n16 2.71565
R674 VTAIL.n56 VTAIL.n55 2.71565
R675 VTAIL.n200 VTAIL.n199 2.71565
R676 VTAIL.n182 VTAIL.n161 2.71565
R677 VTAIL.n130 VTAIL.n129 2.71565
R678 VTAIL.n112 VTAIL.n91 2.71565
R679 VTAIL.n75 VTAIL.n73 2.35395
R680 VTAIL.n141 VTAIL.n75 2.35395
R681 VTAIL.n145 VTAIL.n143 2.35395
R682 VTAIL.n211 VTAIL.n145 2.35395
R683 VTAIL.n71 VTAIL.n69 2.35395
R684 VTAIL.n69 VTAIL.n67 2.35395
R685 VTAIL.n279 VTAIL.n277 2.35395
R686 VTAIL.n248 VTAIL.n224 1.93989
R687 VTAIL.n262 VTAIL.n218 1.93989
R688 VTAIL.n38 VTAIL.n14 1.93989
R689 VTAIL.n52 VTAIL.n8 1.93989
R690 VTAIL.n196 VTAIL.n152 1.93989
R691 VTAIL.n183 VTAIL.n159 1.93989
R692 VTAIL.n126 VTAIL.n82 1.93989
R693 VTAIL.n113 VTAIL.n89 1.93989
R694 VTAIL VTAIL.n1 1.82378
R695 VTAIL.n143 VTAIL.n141 1.64705
R696 VTAIL.n67 VTAIL.n1 1.64705
R697 VTAIL.n278 VTAIL.t8 1.62079
R698 VTAIL.n278 VTAIL.t0 1.62079
R699 VTAIL.n0 VTAIL.t6 1.62079
R700 VTAIL.n0 VTAIL.t7 1.62079
R701 VTAIL.n68 VTAIL.t14 1.62079
R702 VTAIL.n68 VTAIL.t11 1.62079
R703 VTAIL.n70 VTAIL.t16 1.62079
R704 VTAIL.n70 VTAIL.t17 1.62079
R705 VTAIL.n144 VTAIL.t12 1.62079
R706 VTAIL.n144 VTAIL.t15 1.62079
R707 VTAIL.n142 VTAIL.t13 1.62079
R708 VTAIL.n142 VTAIL.t19 1.62079
R709 VTAIL.n74 VTAIL.t2 1.62079
R710 VTAIL.n74 VTAIL.t9 1.62079
R711 VTAIL.n72 VTAIL.t4 1.62079
R712 VTAIL.n72 VTAIL.t1 1.62079
R713 VTAIL.n253 VTAIL.n251 1.16414
R714 VTAIL.n261 VTAIL.n220 1.16414
R715 VTAIL.n43 VTAIL.n41 1.16414
R716 VTAIL.n51 VTAIL.n10 1.16414
R717 VTAIL.n195 VTAIL.n154 1.16414
R718 VTAIL.n187 VTAIL.n186 1.16414
R719 VTAIL.n125 VTAIL.n84 1.16414
R720 VTAIL.n117 VTAIL.n116 1.16414
R721 VTAIL VTAIL.n279 0.530672
R722 VTAIL.n252 VTAIL.n222 0.388379
R723 VTAIL.n258 VTAIL.n257 0.388379
R724 VTAIL.n42 VTAIL.n12 0.388379
R725 VTAIL.n48 VTAIL.n47 0.388379
R726 VTAIL.n192 VTAIL.n191 0.388379
R727 VTAIL.n158 VTAIL.n156 0.388379
R728 VTAIL.n122 VTAIL.n121 0.388379
R729 VTAIL.n88 VTAIL.n86 0.388379
R730 VTAIL.n234 VTAIL.n229 0.155672
R731 VTAIL.n241 VTAIL.n229 0.155672
R732 VTAIL.n242 VTAIL.n241 0.155672
R733 VTAIL.n242 VTAIL.n225 0.155672
R734 VTAIL.n249 VTAIL.n225 0.155672
R735 VTAIL.n250 VTAIL.n249 0.155672
R736 VTAIL.n250 VTAIL.n221 0.155672
R737 VTAIL.n259 VTAIL.n221 0.155672
R738 VTAIL.n260 VTAIL.n259 0.155672
R739 VTAIL.n260 VTAIL.n217 0.155672
R740 VTAIL.n267 VTAIL.n217 0.155672
R741 VTAIL.n268 VTAIL.n267 0.155672
R742 VTAIL.n268 VTAIL.n213 0.155672
R743 VTAIL.n275 VTAIL.n213 0.155672
R744 VTAIL.n24 VTAIL.n19 0.155672
R745 VTAIL.n31 VTAIL.n19 0.155672
R746 VTAIL.n32 VTAIL.n31 0.155672
R747 VTAIL.n32 VTAIL.n15 0.155672
R748 VTAIL.n39 VTAIL.n15 0.155672
R749 VTAIL.n40 VTAIL.n39 0.155672
R750 VTAIL.n40 VTAIL.n11 0.155672
R751 VTAIL.n49 VTAIL.n11 0.155672
R752 VTAIL.n50 VTAIL.n49 0.155672
R753 VTAIL.n50 VTAIL.n7 0.155672
R754 VTAIL.n57 VTAIL.n7 0.155672
R755 VTAIL.n58 VTAIL.n57 0.155672
R756 VTAIL.n58 VTAIL.n3 0.155672
R757 VTAIL.n65 VTAIL.n3 0.155672
R758 VTAIL.n209 VTAIL.n147 0.155672
R759 VTAIL.n202 VTAIL.n147 0.155672
R760 VTAIL.n202 VTAIL.n201 0.155672
R761 VTAIL.n201 VTAIL.n151 0.155672
R762 VTAIL.n194 VTAIL.n151 0.155672
R763 VTAIL.n194 VTAIL.n193 0.155672
R764 VTAIL.n193 VTAIL.n155 0.155672
R765 VTAIL.n185 VTAIL.n155 0.155672
R766 VTAIL.n185 VTAIL.n184 0.155672
R767 VTAIL.n184 VTAIL.n160 0.155672
R768 VTAIL.n177 VTAIL.n160 0.155672
R769 VTAIL.n177 VTAIL.n176 0.155672
R770 VTAIL.n176 VTAIL.n164 0.155672
R771 VTAIL.n169 VTAIL.n164 0.155672
R772 VTAIL.n139 VTAIL.n77 0.155672
R773 VTAIL.n132 VTAIL.n77 0.155672
R774 VTAIL.n132 VTAIL.n131 0.155672
R775 VTAIL.n131 VTAIL.n81 0.155672
R776 VTAIL.n124 VTAIL.n81 0.155672
R777 VTAIL.n124 VTAIL.n123 0.155672
R778 VTAIL.n123 VTAIL.n85 0.155672
R779 VTAIL.n115 VTAIL.n85 0.155672
R780 VTAIL.n115 VTAIL.n114 0.155672
R781 VTAIL.n114 VTAIL.n90 0.155672
R782 VTAIL.n107 VTAIL.n90 0.155672
R783 VTAIL.n107 VTAIL.n106 0.155672
R784 VTAIL.n106 VTAIL.n94 0.155672
R785 VTAIL.n99 VTAIL.n94 0.155672
R786 B.n933 B.n932 585
R787 B.n340 B.n151 585
R788 B.n339 B.n338 585
R789 B.n337 B.n336 585
R790 B.n335 B.n334 585
R791 B.n333 B.n332 585
R792 B.n331 B.n330 585
R793 B.n329 B.n328 585
R794 B.n327 B.n326 585
R795 B.n325 B.n324 585
R796 B.n323 B.n322 585
R797 B.n321 B.n320 585
R798 B.n319 B.n318 585
R799 B.n317 B.n316 585
R800 B.n315 B.n314 585
R801 B.n313 B.n312 585
R802 B.n311 B.n310 585
R803 B.n309 B.n308 585
R804 B.n307 B.n306 585
R805 B.n305 B.n304 585
R806 B.n303 B.n302 585
R807 B.n301 B.n300 585
R808 B.n299 B.n298 585
R809 B.n297 B.n296 585
R810 B.n295 B.n294 585
R811 B.n293 B.n292 585
R812 B.n291 B.n290 585
R813 B.n289 B.n288 585
R814 B.n287 B.n286 585
R815 B.n285 B.n284 585
R816 B.n283 B.n282 585
R817 B.n281 B.n280 585
R818 B.n279 B.n278 585
R819 B.n277 B.n276 585
R820 B.n275 B.n274 585
R821 B.n273 B.n272 585
R822 B.n271 B.n270 585
R823 B.n269 B.n268 585
R824 B.n267 B.n266 585
R825 B.n265 B.n264 585
R826 B.n263 B.n262 585
R827 B.n261 B.n260 585
R828 B.n259 B.n258 585
R829 B.n257 B.n256 585
R830 B.n255 B.n254 585
R831 B.n253 B.n252 585
R832 B.n251 B.n250 585
R833 B.n249 B.n248 585
R834 B.n247 B.n246 585
R835 B.n245 B.n244 585
R836 B.n243 B.n242 585
R837 B.n241 B.n240 585
R838 B.n239 B.n238 585
R839 B.n237 B.n236 585
R840 B.n235 B.n234 585
R841 B.n233 B.n232 585
R842 B.n231 B.n230 585
R843 B.n229 B.n228 585
R844 B.n227 B.n226 585
R845 B.n225 B.n224 585
R846 B.n223 B.n222 585
R847 B.n221 B.n220 585
R848 B.n219 B.n218 585
R849 B.n217 B.n216 585
R850 B.n215 B.n214 585
R851 B.n213 B.n212 585
R852 B.n211 B.n210 585
R853 B.n209 B.n208 585
R854 B.n207 B.n206 585
R855 B.n205 B.n204 585
R856 B.n203 B.n202 585
R857 B.n201 B.n200 585
R858 B.n199 B.n198 585
R859 B.n197 B.n196 585
R860 B.n195 B.n194 585
R861 B.n193 B.n192 585
R862 B.n191 B.n190 585
R863 B.n189 B.n188 585
R864 B.n187 B.n186 585
R865 B.n185 B.n184 585
R866 B.n183 B.n182 585
R867 B.n181 B.n180 585
R868 B.n179 B.n178 585
R869 B.n177 B.n176 585
R870 B.n175 B.n174 585
R871 B.n173 B.n172 585
R872 B.n171 B.n170 585
R873 B.n169 B.n168 585
R874 B.n167 B.n166 585
R875 B.n165 B.n164 585
R876 B.n163 B.n162 585
R877 B.n161 B.n160 585
R878 B.n159 B.n158 585
R879 B.n103 B.n102 585
R880 B.n931 B.n104 585
R881 B.n936 B.n104 585
R882 B.n930 B.n929 585
R883 B.n929 B.n100 585
R884 B.n928 B.n99 585
R885 B.n942 B.n99 585
R886 B.n927 B.n98 585
R887 B.n943 B.n98 585
R888 B.n926 B.n97 585
R889 B.n944 B.n97 585
R890 B.n925 B.n924 585
R891 B.n924 B.n93 585
R892 B.n923 B.n92 585
R893 B.n950 B.n92 585
R894 B.n922 B.n91 585
R895 B.n951 B.n91 585
R896 B.n921 B.n90 585
R897 B.n952 B.n90 585
R898 B.n920 B.n919 585
R899 B.n919 B.n86 585
R900 B.n918 B.n85 585
R901 B.n958 B.n85 585
R902 B.n917 B.n84 585
R903 B.n959 B.n84 585
R904 B.n916 B.n83 585
R905 B.n960 B.n83 585
R906 B.n915 B.n914 585
R907 B.n914 B.n79 585
R908 B.n913 B.n78 585
R909 B.n966 B.n78 585
R910 B.n912 B.n77 585
R911 B.n967 B.n77 585
R912 B.n911 B.n76 585
R913 B.n968 B.n76 585
R914 B.n910 B.n909 585
R915 B.n909 B.n72 585
R916 B.n908 B.n71 585
R917 B.n974 B.n71 585
R918 B.n907 B.n70 585
R919 B.n975 B.n70 585
R920 B.n906 B.n69 585
R921 B.n976 B.n69 585
R922 B.n905 B.n904 585
R923 B.n904 B.n65 585
R924 B.n903 B.n64 585
R925 B.n982 B.n64 585
R926 B.n902 B.n63 585
R927 B.n983 B.n63 585
R928 B.n901 B.n62 585
R929 B.n984 B.n62 585
R930 B.n900 B.n899 585
R931 B.n899 B.n58 585
R932 B.n898 B.n57 585
R933 B.n990 B.n57 585
R934 B.n897 B.n56 585
R935 B.n991 B.n56 585
R936 B.n896 B.n55 585
R937 B.n992 B.n55 585
R938 B.n895 B.n894 585
R939 B.n894 B.n51 585
R940 B.n893 B.n50 585
R941 B.n998 B.n50 585
R942 B.n892 B.n49 585
R943 B.n999 B.n49 585
R944 B.n891 B.n48 585
R945 B.n1000 B.n48 585
R946 B.n890 B.n889 585
R947 B.n889 B.n44 585
R948 B.n888 B.n43 585
R949 B.n1006 B.n43 585
R950 B.n887 B.n42 585
R951 B.n1007 B.n42 585
R952 B.n886 B.n41 585
R953 B.n1008 B.n41 585
R954 B.n885 B.n884 585
R955 B.n884 B.n37 585
R956 B.n883 B.n36 585
R957 B.n1014 B.n36 585
R958 B.n882 B.n35 585
R959 B.n1015 B.n35 585
R960 B.n881 B.n34 585
R961 B.n1016 B.n34 585
R962 B.n880 B.n879 585
R963 B.n879 B.n30 585
R964 B.n878 B.n29 585
R965 B.n1022 B.n29 585
R966 B.n877 B.n28 585
R967 B.n1023 B.n28 585
R968 B.n876 B.n27 585
R969 B.n1024 B.n27 585
R970 B.n875 B.n874 585
R971 B.n874 B.n23 585
R972 B.n873 B.n22 585
R973 B.n1030 B.n22 585
R974 B.n872 B.n21 585
R975 B.n1031 B.n21 585
R976 B.n871 B.n20 585
R977 B.n1032 B.n20 585
R978 B.n870 B.n869 585
R979 B.n869 B.n16 585
R980 B.n868 B.n15 585
R981 B.n1038 B.n15 585
R982 B.n867 B.n14 585
R983 B.n1039 B.n14 585
R984 B.n866 B.n13 585
R985 B.n1040 B.n13 585
R986 B.n865 B.n864 585
R987 B.n864 B.n12 585
R988 B.n863 B.n862 585
R989 B.n863 B.n8 585
R990 B.n861 B.n7 585
R991 B.n1047 B.n7 585
R992 B.n860 B.n6 585
R993 B.n1048 B.n6 585
R994 B.n859 B.n5 585
R995 B.n1049 B.n5 585
R996 B.n858 B.n857 585
R997 B.n857 B.n4 585
R998 B.n856 B.n341 585
R999 B.n856 B.n855 585
R1000 B.n846 B.n342 585
R1001 B.n343 B.n342 585
R1002 B.n848 B.n847 585
R1003 B.n849 B.n848 585
R1004 B.n845 B.n348 585
R1005 B.n348 B.n347 585
R1006 B.n844 B.n843 585
R1007 B.n843 B.n842 585
R1008 B.n350 B.n349 585
R1009 B.n351 B.n350 585
R1010 B.n835 B.n834 585
R1011 B.n836 B.n835 585
R1012 B.n833 B.n356 585
R1013 B.n356 B.n355 585
R1014 B.n832 B.n831 585
R1015 B.n831 B.n830 585
R1016 B.n358 B.n357 585
R1017 B.n359 B.n358 585
R1018 B.n823 B.n822 585
R1019 B.n824 B.n823 585
R1020 B.n821 B.n364 585
R1021 B.n364 B.n363 585
R1022 B.n820 B.n819 585
R1023 B.n819 B.n818 585
R1024 B.n366 B.n365 585
R1025 B.n367 B.n366 585
R1026 B.n811 B.n810 585
R1027 B.n812 B.n811 585
R1028 B.n809 B.n372 585
R1029 B.n372 B.n371 585
R1030 B.n808 B.n807 585
R1031 B.n807 B.n806 585
R1032 B.n374 B.n373 585
R1033 B.n375 B.n374 585
R1034 B.n799 B.n798 585
R1035 B.n800 B.n799 585
R1036 B.n797 B.n380 585
R1037 B.n380 B.n379 585
R1038 B.n796 B.n795 585
R1039 B.n795 B.n794 585
R1040 B.n382 B.n381 585
R1041 B.n383 B.n382 585
R1042 B.n787 B.n786 585
R1043 B.n788 B.n787 585
R1044 B.n785 B.n388 585
R1045 B.n388 B.n387 585
R1046 B.n784 B.n783 585
R1047 B.n783 B.n782 585
R1048 B.n390 B.n389 585
R1049 B.n391 B.n390 585
R1050 B.n775 B.n774 585
R1051 B.n776 B.n775 585
R1052 B.n773 B.n396 585
R1053 B.n396 B.n395 585
R1054 B.n772 B.n771 585
R1055 B.n771 B.n770 585
R1056 B.n398 B.n397 585
R1057 B.n399 B.n398 585
R1058 B.n763 B.n762 585
R1059 B.n764 B.n763 585
R1060 B.n761 B.n404 585
R1061 B.n404 B.n403 585
R1062 B.n760 B.n759 585
R1063 B.n759 B.n758 585
R1064 B.n406 B.n405 585
R1065 B.n407 B.n406 585
R1066 B.n751 B.n750 585
R1067 B.n752 B.n751 585
R1068 B.n749 B.n412 585
R1069 B.n412 B.n411 585
R1070 B.n748 B.n747 585
R1071 B.n747 B.n746 585
R1072 B.n414 B.n413 585
R1073 B.n415 B.n414 585
R1074 B.n739 B.n738 585
R1075 B.n740 B.n739 585
R1076 B.n737 B.n420 585
R1077 B.n420 B.n419 585
R1078 B.n736 B.n735 585
R1079 B.n735 B.n734 585
R1080 B.n422 B.n421 585
R1081 B.n423 B.n422 585
R1082 B.n727 B.n726 585
R1083 B.n728 B.n727 585
R1084 B.n725 B.n428 585
R1085 B.n428 B.n427 585
R1086 B.n724 B.n723 585
R1087 B.n723 B.n722 585
R1088 B.n430 B.n429 585
R1089 B.n431 B.n430 585
R1090 B.n715 B.n714 585
R1091 B.n716 B.n715 585
R1092 B.n713 B.n435 585
R1093 B.n439 B.n435 585
R1094 B.n712 B.n711 585
R1095 B.n711 B.n710 585
R1096 B.n437 B.n436 585
R1097 B.n438 B.n437 585
R1098 B.n703 B.n702 585
R1099 B.n704 B.n703 585
R1100 B.n701 B.n444 585
R1101 B.n444 B.n443 585
R1102 B.n700 B.n699 585
R1103 B.n699 B.n698 585
R1104 B.n446 B.n445 585
R1105 B.n447 B.n446 585
R1106 B.n691 B.n690 585
R1107 B.n692 B.n691 585
R1108 B.n450 B.n449 585
R1109 B.n503 B.n501 585
R1110 B.n504 B.n500 585
R1111 B.n504 B.n451 585
R1112 B.n507 B.n506 585
R1113 B.n508 B.n499 585
R1114 B.n510 B.n509 585
R1115 B.n512 B.n498 585
R1116 B.n515 B.n514 585
R1117 B.n516 B.n497 585
R1118 B.n518 B.n517 585
R1119 B.n520 B.n496 585
R1120 B.n523 B.n522 585
R1121 B.n524 B.n495 585
R1122 B.n526 B.n525 585
R1123 B.n528 B.n494 585
R1124 B.n531 B.n530 585
R1125 B.n532 B.n493 585
R1126 B.n534 B.n533 585
R1127 B.n536 B.n492 585
R1128 B.n539 B.n538 585
R1129 B.n540 B.n491 585
R1130 B.n542 B.n541 585
R1131 B.n544 B.n490 585
R1132 B.n547 B.n546 585
R1133 B.n548 B.n489 585
R1134 B.n550 B.n549 585
R1135 B.n552 B.n488 585
R1136 B.n555 B.n554 585
R1137 B.n556 B.n487 585
R1138 B.n558 B.n557 585
R1139 B.n560 B.n486 585
R1140 B.n563 B.n562 585
R1141 B.n564 B.n485 585
R1142 B.n566 B.n565 585
R1143 B.n568 B.n484 585
R1144 B.n571 B.n570 585
R1145 B.n572 B.n483 585
R1146 B.n574 B.n573 585
R1147 B.n576 B.n482 585
R1148 B.n579 B.n578 585
R1149 B.n580 B.n481 585
R1150 B.n585 B.n584 585
R1151 B.n587 B.n480 585
R1152 B.n590 B.n589 585
R1153 B.n591 B.n479 585
R1154 B.n593 B.n592 585
R1155 B.n595 B.n478 585
R1156 B.n598 B.n597 585
R1157 B.n599 B.n477 585
R1158 B.n601 B.n600 585
R1159 B.n603 B.n476 585
R1160 B.n606 B.n605 585
R1161 B.n608 B.n473 585
R1162 B.n610 B.n609 585
R1163 B.n612 B.n472 585
R1164 B.n615 B.n614 585
R1165 B.n616 B.n471 585
R1166 B.n618 B.n617 585
R1167 B.n620 B.n470 585
R1168 B.n623 B.n622 585
R1169 B.n624 B.n469 585
R1170 B.n626 B.n625 585
R1171 B.n628 B.n468 585
R1172 B.n631 B.n630 585
R1173 B.n632 B.n467 585
R1174 B.n634 B.n633 585
R1175 B.n636 B.n466 585
R1176 B.n639 B.n638 585
R1177 B.n640 B.n465 585
R1178 B.n642 B.n641 585
R1179 B.n644 B.n464 585
R1180 B.n647 B.n646 585
R1181 B.n648 B.n463 585
R1182 B.n650 B.n649 585
R1183 B.n652 B.n462 585
R1184 B.n655 B.n654 585
R1185 B.n656 B.n461 585
R1186 B.n658 B.n657 585
R1187 B.n660 B.n460 585
R1188 B.n663 B.n662 585
R1189 B.n664 B.n459 585
R1190 B.n666 B.n665 585
R1191 B.n668 B.n458 585
R1192 B.n671 B.n670 585
R1193 B.n672 B.n457 585
R1194 B.n674 B.n673 585
R1195 B.n676 B.n456 585
R1196 B.n679 B.n678 585
R1197 B.n680 B.n455 585
R1198 B.n682 B.n681 585
R1199 B.n684 B.n454 585
R1200 B.n685 B.n453 585
R1201 B.n688 B.n687 585
R1202 B.n689 B.n452 585
R1203 B.n452 B.n451 585
R1204 B.n694 B.n693 585
R1205 B.n693 B.n692 585
R1206 B.n695 B.n448 585
R1207 B.n448 B.n447 585
R1208 B.n697 B.n696 585
R1209 B.n698 B.n697 585
R1210 B.n442 B.n441 585
R1211 B.n443 B.n442 585
R1212 B.n706 B.n705 585
R1213 B.n705 B.n704 585
R1214 B.n707 B.n440 585
R1215 B.n440 B.n438 585
R1216 B.n709 B.n708 585
R1217 B.n710 B.n709 585
R1218 B.n434 B.n433 585
R1219 B.n439 B.n434 585
R1220 B.n718 B.n717 585
R1221 B.n717 B.n716 585
R1222 B.n719 B.n432 585
R1223 B.n432 B.n431 585
R1224 B.n721 B.n720 585
R1225 B.n722 B.n721 585
R1226 B.n426 B.n425 585
R1227 B.n427 B.n426 585
R1228 B.n730 B.n729 585
R1229 B.n729 B.n728 585
R1230 B.n731 B.n424 585
R1231 B.n424 B.n423 585
R1232 B.n733 B.n732 585
R1233 B.n734 B.n733 585
R1234 B.n418 B.n417 585
R1235 B.n419 B.n418 585
R1236 B.n742 B.n741 585
R1237 B.n741 B.n740 585
R1238 B.n743 B.n416 585
R1239 B.n416 B.n415 585
R1240 B.n745 B.n744 585
R1241 B.n746 B.n745 585
R1242 B.n410 B.n409 585
R1243 B.n411 B.n410 585
R1244 B.n754 B.n753 585
R1245 B.n753 B.n752 585
R1246 B.n755 B.n408 585
R1247 B.n408 B.n407 585
R1248 B.n757 B.n756 585
R1249 B.n758 B.n757 585
R1250 B.n402 B.n401 585
R1251 B.n403 B.n402 585
R1252 B.n766 B.n765 585
R1253 B.n765 B.n764 585
R1254 B.n767 B.n400 585
R1255 B.n400 B.n399 585
R1256 B.n769 B.n768 585
R1257 B.n770 B.n769 585
R1258 B.n394 B.n393 585
R1259 B.n395 B.n394 585
R1260 B.n778 B.n777 585
R1261 B.n777 B.n776 585
R1262 B.n779 B.n392 585
R1263 B.n392 B.n391 585
R1264 B.n781 B.n780 585
R1265 B.n782 B.n781 585
R1266 B.n386 B.n385 585
R1267 B.n387 B.n386 585
R1268 B.n790 B.n789 585
R1269 B.n789 B.n788 585
R1270 B.n791 B.n384 585
R1271 B.n384 B.n383 585
R1272 B.n793 B.n792 585
R1273 B.n794 B.n793 585
R1274 B.n378 B.n377 585
R1275 B.n379 B.n378 585
R1276 B.n802 B.n801 585
R1277 B.n801 B.n800 585
R1278 B.n803 B.n376 585
R1279 B.n376 B.n375 585
R1280 B.n805 B.n804 585
R1281 B.n806 B.n805 585
R1282 B.n370 B.n369 585
R1283 B.n371 B.n370 585
R1284 B.n814 B.n813 585
R1285 B.n813 B.n812 585
R1286 B.n815 B.n368 585
R1287 B.n368 B.n367 585
R1288 B.n817 B.n816 585
R1289 B.n818 B.n817 585
R1290 B.n362 B.n361 585
R1291 B.n363 B.n362 585
R1292 B.n826 B.n825 585
R1293 B.n825 B.n824 585
R1294 B.n827 B.n360 585
R1295 B.n360 B.n359 585
R1296 B.n829 B.n828 585
R1297 B.n830 B.n829 585
R1298 B.n354 B.n353 585
R1299 B.n355 B.n354 585
R1300 B.n838 B.n837 585
R1301 B.n837 B.n836 585
R1302 B.n839 B.n352 585
R1303 B.n352 B.n351 585
R1304 B.n841 B.n840 585
R1305 B.n842 B.n841 585
R1306 B.n346 B.n345 585
R1307 B.n347 B.n346 585
R1308 B.n851 B.n850 585
R1309 B.n850 B.n849 585
R1310 B.n852 B.n344 585
R1311 B.n344 B.n343 585
R1312 B.n854 B.n853 585
R1313 B.n855 B.n854 585
R1314 B.n3 B.n0 585
R1315 B.n4 B.n3 585
R1316 B.n1046 B.n1 585
R1317 B.n1047 B.n1046 585
R1318 B.n1045 B.n1044 585
R1319 B.n1045 B.n8 585
R1320 B.n1043 B.n9 585
R1321 B.n12 B.n9 585
R1322 B.n1042 B.n1041 585
R1323 B.n1041 B.n1040 585
R1324 B.n11 B.n10 585
R1325 B.n1039 B.n11 585
R1326 B.n1037 B.n1036 585
R1327 B.n1038 B.n1037 585
R1328 B.n1035 B.n17 585
R1329 B.n17 B.n16 585
R1330 B.n1034 B.n1033 585
R1331 B.n1033 B.n1032 585
R1332 B.n19 B.n18 585
R1333 B.n1031 B.n19 585
R1334 B.n1029 B.n1028 585
R1335 B.n1030 B.n1029 585
R1336 B.n1027 B.n24 585
R1337 B.n24 B.n23 585
R1338 B.n1026 B.n1025 585
R1339 B.n1025 B.n1024 585
R1340 B.n26 B.n25 585
R1341 B.n1023 B.n26 585
R1342 B.n1021 B.n1020 585
R1343 B.n1022 B.n1021 585
R1344 B.n1019 B.n31 585
R1345 B.n31 B.n30 585
R1346 B.n1018 B.n1017 585
R1347 B.n1017 B.n1016 585
R1348 B.n33 B.n32 585
R1349 B.n1015 B.n33 585
R1350 B.n1013 B.n1012 585
R1351 B.n1014 B.n1013 585
R1352 B.n1011 B.n38 585
R1353 B.n38 B.n37 585
R1354 B.n1010 B.n1009 585
R1355 B.n1009 B.n1008 585
R1356 B.n40 B.n39 585
R1357 B.n1007 B.n40 585
R1358 B.n1005 B.n1004 585
R1359 B.n1006 B.n1005 585
R1360 B.n1003 B.n45 585
R1361 B.n45 B.n44 585
R1362 B.n1002 B.n1001 585
R1363 B.n1001 B.n1000 585
R1364 B.n47 B.n46 585
R1365 B.n999 B.n47 585
R1366 B.n997 B.n996 585
R1367 B.n998 B.n997 585
R1368 B.n995 B.n52 585
R1369 B.n52 B.n51 585
R1370 B.n994 B.n993 585
R1371 B.n993 B.n992 585
R1372 B.n54 B.n53 585
R1373 B.n991 B.n54 585
R1374 B.n989 B.n988 585
R1375 B.n990 B.n989 585
R1376 B.n987 B.n59 585
R1377 B.n59 B.n58 585
R1378 B.n986 B.n985 585
R1379 B.n985 B.n984 585
R1380 B.n61 B.n60 585
R1381 B.n983 B.n61 585
R1382 B.n981 B.n980 585
R1383 B.n982 B.n981 585
R1384 B.n979 B.n66 585
R1385 B.n66 B.n65 585
R1386 B.n978 B.n977 585
R1387 B.n977 B.n976 585
R1388 B.n68 B.n67 585
R1389 B.n975 B.n68 585
R1390 B.n973 B.n972 585
R1391 B.n974 B.n973 585
R1392 B.n971 B.n73 585
R1393 B.n73 B.n72 585
R1394 B.n970 B.n969 585
R1395 B.n969 B.n968 585
R1396 B.n75 B.n74 585
R1397 B.n967 B.n75 585
R1398 B.n965 B.n964 585
R1399 B.n966 B.n965 585
R1400 B.n963 B.n80 585
R1401 B.n80 B.n79 585
R1402 B.n962 B.n961 585
R1403 B.n961 B.n960 585
R1404 B.n82 B.n81 585
R1405 B.n959 B.n82 585
R1406 B.n957 B.n956 585
R1407 B.n958 B.n957 585
R1408 B.n955 B.n87 585
R1409 B.n87 B.n86 585
R1410 B.n954 B.n953 585
R1411 B.n953 B.n952 585
R1412 B.n89 B.n88 585
R1413 B.n951 B.n89 585
R1414 B.n949 B.n948 585
R1415 B.n950 B.n949 585
R1416 B.n947 B.n94 585
R1417 B.n94 B.n93 585
R1418 B.n946 B.n945 585
R1419 B.n945 B.n944 585
R1420 B.n96 B.n95 585
R1421 B.n943 B.n96 585
R1422 B.n941 B.n940 585
R1423 B.n942 B.n941 585
R1424 B.n939 B.n101 585
R1425 B.n101 B.n100 585
R1426 B.n938 B.n937 585
R1427 B.n937 B.n936 585
R1428 B.n1050 B.n1049 585
R1429 B.n1048 B.n2 585
R1430 B.n937 B.n103 473.281
R1431 B.n933 B.n104 473.281
R1432 B.n691 B.n452 473.281
R1433 B.n693 B.n450 473.281
R1434 B.n152 B.t22 339.221
R1435 B.n474 B.t20 339.221
R1436 B.n155 B.t16 339.221
R1437 B.n581 B.t13 339.221
R1438 B.n155 B.t14 330.433
R1439 B.n152 B.t21 330.433
R1440 B.n474 B.t18 330.433
R1441 B.n581 B.t10 330.433
R1442 B.n153 B.t23 286.274
R1443 B.n475 B.t19 286.274
R1444 B.n156 B.t17 286.274
R1445 B.n582 B.t12 286.274
R1446 B.n935 B.n934 256.663
R1447 B.n935 B.n150 256.663
R1448 B.n935 B.n149 256.663
R1449 B.n935 B.n148 256.663
R1450 B.n935 B.n147 256.663
R1451 B.n935 B.n146 256.663
R1452 B.n935 B.n145 256.663
R1453 B.n935 B.n144 256.663
R1454 B.n935 B.n143 256.663
R1455 B.n935 B.n142 256.663
R1456 B.n935 B.n141 256.663
R1457 B.n935 B.n140 256.663
R1458 B.n935 B.n139 256.663
R1459 B.n935 B.n138 256.663
R1460 B.n935 B.n137 256.663
R1461 B.n935 B.n136 256.663
R1462 B.n935 B.n135 256.663
R1463 B.n935 B.n134 256.663
R1464 B.n935 B.n133 256.663
R1465 B.n935 B.n132 256.663
R1466 B.n935 B.n131 256.663
R1467 B.n935 B.n130 256.663
R1468 B.n935 B.n129 256.663
R1469 B.n935 B.n128 256.663
R1470 B.n935 B.n127 256.663
R1471 B.n935 B.n126 256.663
R1472 B.n935 B.n125 256.663
R1473 B.n935 B.n124 256.663
R1474 B.n935 B.n123 256.663
R1475 B.n935 B.n122 256.663
R1476 B.n935 B.n121 256.663
R1477 B.n935 B.n120 256.663
R1478 B.n935 B.n119 256.663
R1479 B.n935 B.n118 256.663
R1480 B.n935 B.n117 256.663
R1481 B.n935 B.n116 256.663
R1482 B.n935 B.n115 256.663
R1483 B.n935 B.n114 256.663
R1484 B.n935 B.n113 256.663
R1485 B.n935 B.n112 256.663
R1486 B.n935 B.n111 256.663
R1487 B.n935 B.n110 256.663
R1488 B.n935 B.n109 256.663
R1489 B.n935 B.n108 256.663
R1490 B.n935 B.n107 256.663
R1491 B.n935 B.n106 256.663
R1492 B.n935 B.n105 256.663
R1493 B.n502 B.n451 256.663
R1494 B.n505 B.n451 256.663
R1495 B.n511 B.n451 256.663
R1496 B.n513 B.n451 256.663
R1497 B.n519 B.n451 256.663
R1498 B.n521 B.n451 256.663
R1499 B.n527 B.n451 256.663
R1500 B.n529 B.n451 256.663
R1501 B.n535 B.n451 256.663
R1502 B.n537 B.n451 256.663
R1503 B.n543 B.n451 256.663
R1504 B.n545 B.n451 256.663
R1505 B.n551 B.n451 256.663
R1506 B.n553 B.n451 256.663
R1507 B.n559 B.n451 256.663
R1508 B.n561 B.n451 256.663
R1509 B.n567 B.n451 256.663
R1510 B.n569 B.n451 256.663
R1511 B.n575 B.n451 256.663
R1512 B.n577 B.n451 256.663
R1513 B.n586 B.n451 256.663
R1514 B.n588 B.n451 256.663
R1515 B.n594 B.n451 256.663
R1516 B.n596 B.n451 256.663
R1517 B.n602 B.n451 256.663
R1518 B.n604 B.n451 256.663
R1519 B.n611 B.n451 256.663
R1520 B.n613 B.n451 256.663
R1521 B.n619 B.n451 256.663
R1522 B.n621 B.n451 256.663
R1523 B.n627 B.n451 256.663
R1524 B.n629 B.n451 256.663
R1525 B.n635 B.n451 256.663
R1526 B.n637 B.n451 256.663
R1527 B.n643 B.n451 256.663
R1528 B.n645 B.n451 256.663
R1529 B.n651 B.n451 256.663
R1530 B.n653 B.n451 256.663
R1531 B.n659 B.n451 256.663
R1532 B.n661 B.n451 256.663
R1533 B.n667 B.n451 256.663
R1534 B.n669 B.n451 256.663
R1535 B.n675 B.n451 256.663
R1536 B.n677 B.n451 256.663
R1537 B.n683 B.n451 256.663
R1538 B.n686 B.n451 256.663
R1539 B.n1052 B.n1051 256.663
R1540 B.n160 B.n159 163.367
R1541 B.n164 B.n163 163.367
R1542 B.n168 B.n167 163.367
R1543 B.n172 B.n171 163.367
R1544 B.n176 B.n175 163.367
R1545 B.n180 B.n179 163.367
R1546 B.n184 B.n183 163.367
R1547 B.n188 B.n187 163.367
R1548 B.n192 B.n191 163.367
R1549 B.n196 B.n195 163.367
R1550 B.n200 B.n199 163.367
R1551 B.n204 B.n203 163.367
R1552 B.n208 B.n207 163.367
R1553 B.n212 B.n211 163.367
R1554 B.n216 B.n215 163.367
R1555 B.n220 B.n219 163.367
R1556 B.n224 B.n223 163.367
R1557 B.n228 B.n227 163.367
R1558 B.n232 B.n231 163.367
R1559 B.n236 B.n235 163.367
R1560 B.n240 B.n239 163.367
R1561 B.n244 B.n243 163.367
R1562 B.n248 B.n247 163.367
R1563 B.n252 B.n251 163.367
R1564 B.n256 B.n255 163.367
R1565 B.n260 B.n259 163.367
R1566 B.n264 B.n263 163.367
R1567 B.n268 B.n267 163.367
R1568 B.n272 B.n271 163.367
R1569 B.n276 B.n275 163.367
R1570 B.n280 B.n279 163.367
R1571 B.n284 B.n283 163.367
R1572 B.n288 B.n287 163.367
R1573 B.n292 B.n291 163.367
R1574 B.n296 B.n295 163.367
R1575 B.n300 B.n299 163.367
R1576 B.n304 B.n303 163.367
R1577 B.n308 B.n307 163.367
R1578 B.n312 B.n311 163.367
R1579 B.n316 B.n315 163.367
R1580 B.n320 B.n319 163.367
R1581 B.n324 B.n323 163.367
R1582 B.n328 B.n327 163.367
R1583 B.n332 B.n331 163.367
R1584 B.n336 B.n335 163.367
R1585 B.n338 B.n151 163.367
R1586 B.n691 B.n446 163.367
R1587 B.n699 B.n446 163.367
R1588 B.n699 B.n444 163.367
R1589 B.n703 B.n444 163.367
R1590 B.n703 B.n437 163.367
R1591 B.n711 B.n437 163.367
R1592 B.n711 B.n435 163.367
R1593 B.n715 B.n435 163.367
R1594 B.n715 B.n430 163.367
R1595 B.n723 B.n430 163.367
R1596 B.n723 B.n428 163.367
R1597 B.n727 B.n428 163.367
R1598 B.n727 B.n422 163.367
R1599 B.n735 B.n422 163.367
R1600 B.n735 B.n420 163.367
R1601 B.n739 B.n420 163.367
R1602 B.n739 B.n414 163.367
R1603 B.n747 B.n414 163.367
R1604 B.n747 B.n412 163.367
R1605 B.n751 B.n412 163.367
R1606 B.n751 B.n406 163.367
R1607 B.n759 B.n406 163.367
R1608 B.n759 B.n404 163.367
R1609 B.n763 B.n404 163.367
R1610 B.n763 B.n398 163.367
R1611 B.n771 B.n398 163.367
R1612 B.n771 B.n396 163.367
R1613 B.n775 B.n396 163.367
R1614 B.n775 B.n390 163.367
R1615 B.n783 B.n390 163.367
R1616 B.n783 B.n388 163.367
R1617 B.n787 B.n388 163.367
R1618 B.n787 B.n382 163.367
R1619 B.n795 B.n382 163.367
R1620 B.n795 B.n380 163.367
R1621 B.n799 B.n380 163.367
R1622 B.n799 B.n374 163.367
R1623 B.n807 B.n374 163.367
R1624 B.n807 B.n372 163.367
R1625 B.n811 B.n372 163.367
R1626 B.n811 B.n366 163.367
R1627 B.n819 B.n366 163.367
R1628 B.n819 B.n364 163.367
R1629 B.n823 B.n364 163.367
R1630 B.n823 B.n358 163.367
R1631 B.n831 B.n358 163.367
R1632 B.n831 B.n356 163.367
R1633 B.n835 B.n356 163.367
R1634 B.n835 B.n350 163.367
R1635 B.n843 B.n350 163.367
R1636 B.n843 B.n348 163.367
R1637 B.n848 B.n348 163.367
R1638 B.n848 B.n342 163.367
R1639 B.n856 B.n342 163.367
R1640 B.n857 B.n856 163.367
R1641 B.n857 B.n5 163.367
R1642 B.n6 B.n5 163.367
R1643 B.n7 B.n6 163.367
R1644 B.n863 B.n7 163.367
R1645 B.n864 B.n863 163.367
R1646 B.n864 B.n13 163.367
R1647 B.n14 B.n13 163.367
R1648 B.n15 B.n14 163.367
R1649 B.n869 B.n15 163.367
R1650 B.n869 B.n20 163.367
R1651 B.n21 B.n20 163.367
R1652 B.n22 B.n21 163.367
R1653 B.n874 B.n22 163.367
R1654 B.n874 B.n27 163.367
R1655 B.n28 B.n27 163.367
R1656 B.n29 B.n28 163.367
R1657 B.n879 B.n29 163.367
R1658 B.n879 B.n34 163.367
R1659 B.n35 B.n34 163.367
R1660 B.n36 B.n35 163.367
R1661 B.n884 B.n36 163.367
R1662 B.n884 B.n41 163.367
R1663 B.n42 B.n41 163.367
R1664 B.n43 B.n42 163.367
R1665 B.n889 B.n43 163.367
R1666 B.n889 B.n48 163.367
R1667 B.n49 B.n48 163.367
R1668 B.n50 B.n49 163.367
R1669 B.n894 B.n50 163.367
R1670 B.n894 B.n55 163.367
R1671 B.n56 B.n55 163.367
R1672 B.n57 B.n56 163.367
R1673 B.n899 B.n57 163.367
R1674 B.n899 B.n62 163.367
R1675 B.n63 B.n62 163.367
R1676 B.n64 B.n63 163.367
R1677 B.n904 B.n64 163.367
R1678 B.n904 B.n69 163.367
R1679 B.n70 B.n69 163.367
R1680 B.n71 B.n70 163.367
R1681 B.n909 B.n71 163.367
R1682 B.n909 B.n76 163.367
R1683 B.n77 B.n76 163.367
R1684 B.n78 B.n77 163.367
R1685 B.n914 B.n78 163.367
R1686 B.n914 B.n83 163.367
R1687 B.n84 B.n83 163.367
R1688 B.n85 B.n84 163.367
R1689 B.n919 B.n85 163.367
R1690 B.n919 B.n90 163.367
R1691 B.n91 B.n90 163.367
R1692 B.n92 B.n91 163.367
R1693 B.n924 B.n92 163.367
R1694 B.n924 B.n97 163.367
R1695 B.n98 B.n97 163.367
R1696 B.n99 B.n98 163.367
R1697 B.n929 B.n99 163.367
R1698 B.n929 B.n104 163.367
R1699 B.n504 B.n503 163.367
R1700 B.n506 B.n504 163.367
R1701 B.n510 B.n499 163.367
R1702 B.n514 B.n512 163.367
R1703 B.n518 B.n497 163.367
R1704 B.n522 B.n520 163.367
R1705 B.n526 B.n495 163.367
R1706 B.n530 B.n528 163.367
R1707 B.n534 B.n493 163.367
R1708 B.n538 B.n536 163.367
R1709 B.n542 B.n491 163.367
R1710 B.n546 B.n544 163.367
R1711 B.n550 B.n489 163.367
R1712 B.n554 B.n552 163.367
R1713 B.n558 B.n487 163.367
R1714 B.n562 B.n560 163.367
R1715 B.n566 B.n485 163.367
R1716 B.n570 B.n568 163.367
R1717 B.n574 B.n483 163.367
R1718 B.n578 B.n576 163.367
R1719 B.n585 B.n481 163.367
R1720 B.n589 B.n587 163.367
R1721 B.n593 B.n479 163.367
R1722 B.n597 B.n595 163.367
R1723 B.n601 B.n477 163.367
R1724 B.n605 B.n603 163.367
R1725 B.n610 B.n473 163.367
R1726 B.n614 B.n612 163.367
R1727 B.n618 B.n471 163.367
R1728 B.n622 B.n620 163.367
R1729 B.n626 B.n469 163.367
R1730 B.n630 B.n628 163.367
R1731 B.n634 B.n467 163.367
R1732 B.n638 B.n636 163.367
R1733 B.n642 B.n465 163.367
R1734 B.n646 B.n644 163.367
R1735 B.n650 B.n463 163.367
R1736 B.n654 B.n652 163.367
R1737 B.n658 B.n461 163.367
R1738 B.n662 B.n660 163.367
R1739 B.n666 B.n459 163.367
R1740 B.n670 B.n668 163.367
R1741 B.n674 B.n457 163.367
R1742 B.n678 B.n676 163.367
R1743 B.n682 B.n455 163.367
R1744 B.n685 B.n684 163.367
R1745 B.n687 B.n452 163.367
R1746 B.n693 B.n448 163.367
R1747 B.n697 B.n448 163.367
R1748 B.n697 B.n442 163.367
R1749 B.n705 B.n442 163.367
R1750 B.n705 B.n440 163.367
R1751 B.n709 B.n440 163.367
R1752 B.n709 B.n434 163.367
R1753 B.n717 B.n434 163.367
R1754 B.n717 B.n432 163.367
R1755 B.n721 B.n432 163.367
R1756 B.n721 B.n426 163.367
R1757 B.n729 B.n426 163.367
R1758 B.n729 B.n424 163.367
R1759 B.n733 B.n424 163.367
R1760 B.n733 B.n418 163.367
R1761 B.n741 B.n418 163.367
R1762 B.n741 B.n416 163.367
R1763 B.n745 B.n416 163.367
R1764 B.n745 B.n410 163.367
R1765 B.n753 B.n410 163.367
R1766 B.n753 B.n408 163.367
R1767 B.n757 B.n408 163.367
R1768 B.n757 B.n402 163.367
R1769 B.n765 B.n402 163.367
R1770 B.n765 B.n400 163.367
R1771 B.n769 B.n400 163.367
R1772 B.n769 B.n394 163.367
R1773 B.n777 B.n394 163.367
R1774 B.n777 B.n392 163.367
R1775 B.n781 B.n392 163.367
R1776 B.n781 B.n386 163.367
R1777 B.n789 B.n386 163.367
R1778 B.n789 B.n384 163.367
R1779 B.n793 B.n384 163.367
R1780 B.n793 B.n378 163.367
R1781 B.n801 B.n378 163.367
R1782 B.n801 B.n376 163.367
R1783 B.n805 B.n376 163.367
R1784 B.n805 B.n370 163.367
R1785 B.n813 B.n370 163.367
R1786 B.n813 B.n368 163.367
R1787 B.n817 B.n368 163.367
R1788 B.n817 B.n362 163.367
R1789 B.n825 B.n362 163.367
R1790 B.n825 B.n360 163.367
R1791 B.n829 B.n360 163.367
R1792 B.n829 B.n354 163.367
R1793 B.n837 B.n354 163.367
R1794 B.n837 B.n352 163.367
R1795 B.n841 B.n352 163.367
R1796 B.n841 B.n346 163.367
R1797 B.n850 B.n346 163.367
R1798 B.n850 B.n344 163.367
R1799 B.n854 B.n344 163.367
R1800 B.n854 B.n3 163.367
R1801 B.n1050 B.n3 163.367
R1802 B.n1046 B.n2 163.367
R1803 B.n1046 B.n1045 163.367
R1804 B.n1045 B.n9 163.367
R1805 B.n1041 B.n9 163.367
R1806 B.n1041 B.n11 163.367
R1807 B.n1037 B.n11 163.367
R1808 B.n1037 B.n17 163.367
R1809 B.n1033 B.n17 163.367
R1810 B.n1033 B.n19 163.367
R1811 B.n1029 B.n19 163.367
R1812 B.n1029 B.n24 163.367
R1813 B.n1025 B.n24 163.367
R1814 B.n1025 B.n26 163.367
R1815 B.n1021 B.n26 163.367
R1816 B.n1021 B.n31 163.367
R1817 B.n1017 B.n31 163.367
R1818 B.n1017 B.n33 163.367
R1819 B.n1013 B.n33 163.367
R1820 B.n1013 B.n38 163.367
R1821 B.n1009 B.n38 163.367
R1822 B.n1009 B.n40 163.367
R1823 B.n1005 B.n40 163.367
R1824 B.n1005 B.n45 163.367
R1825 B.n1001 B.n45 163.367
R1826 B.n1001 B.n47 163.367
R1827 B.n997 B.n47 163.367
R1828 B.n997 B.n52 163.367
R1829 B.n993 B.n52 163.367
R1830 B.n993 B.n54 163.367
R1831 B.n989 B.n54 163.367
R1832 B.n989 B.n59 163.367
R1833 B.n985 B.n59 163.367
R1834 B.n985 B.n61 163.367
R1835 B.n981 B.n61 163.367
R1836 B.n981 B.n66 163.367
R1837 B.n977 B.n66 163.367
R1838 B.n977 B.n68 163.367
R1839 B.n973 B.n68 163.367
R1840 B.n973 B.n73 163.367
R1841 B.n969 B.n73 163.367
R1842 B.n969 B.n75 163.367
R1843 B.n965 B.n75 163.367
R1844 B.n965 B.n80 163.367
R1845 B.n961 B.n80 163.367
R1846 B.n961 B.n82 163.367
R1847 B.n957 B.n82 163.367
R1848 B.n957 B.n87 163.367
R1849 B.n953 B.n87 163.367
R1850 B.n953 B.n89 163.367
R1851 B.n949 B.n89 163.367
R1852 B.n949 B.n94 163.367
R1853 B.n945 B.n94 163.367
R1854 B.n945 B.n96 163.367
R1855 B.n941 B.n96 163.367
R1856 B.n941 B.n101 163.367
R1857 B.n937 B.n101 163.367
R1858 B.n105 B.n103 71.676
R1859 B.n160 B.n106 71.676
R1860 B.n164 B.n107 71.676
R1861 B.n168 B.n108 71.676
R1862 B.n172 B.n109 71.676
R1863 B.n176 B.n110 71.676
R1864 B.n180 B.n111 71.676
R1865 B.n184 B.n112 71.676
R1866 B.n188 B.n113 71.676
R1867 B.n192 B.n114 71.676
R1868 B.n196 B.n115 71.676
R1869 B.n200 B.n116 71.676
R1870 B.n204 B.n117 71.676
R1871 B.n208 B.n118 71.676
R1872 B.n212 B.n119 71.676
R1873 B.n216 B.n120 71.676
R1874 B.n220 B.n121 71.676
R1875 B.n224 B.n122 71.676
R1876 B.n228 B.n123 71.676
R1877 B.n232 B.n124 71.676
R1878 B.n236 B.n125 71.676
R1879 B.n240 B.n126 71.676
R1880 B.n244 B.n127 71.676
R1881 B.n248 B.n128 71.676
R1882 B.n252 B.n129 71.676
R1883 B.n256 B.n130 71.676
R1884 B.n260 B.n131 71.676
R1885 B.n264 B.n132 71.676
R1886 B.n268 B.n133 71.676
R1887 B.n272 B.n134 71.676
R1888 B.n276 B.n135 71.676
R1889 B.n280 B.n136 71.676
R1890 B.n284 B.n137 71.676
R1891 B.n288 B.n138 71.676
R1892 B.n292 B.n139 71.676
R1893 B.n296 B.n140 71.676
R1894 B.n300 B.n141 71.676
R1895 B.n304 B.n142 71.676
R1896 B.n308 B.n143 71.676
R1897 B.n312 B.n144 71.676
R1898 B.n316 B.n145 71.676
R1899 B.n320 B.n146 71.676
R1900 B.n324 B.n147 71.676
R1901 B.n328 B.n148 71.676
R1902 B.n332 B.n149 71.676
R1903 B.n336 B.n150 71.676
R1904 B.n934 B.n151 71.676
R1905 B.n934 B.n933 71.676
R1906 B.n338 B.n150 71.676
R1907 B.n335 B.n149 71.676
R1908 B.n331 B.n148 71.676
R1909 B.n327 B.n147 71.676
R1910 B.n323 B.n146 71.676
R1911 B.n319 B.n145 71.676
R1912 B.n315 B.n144 71.676
R1913 B.n311 B.n143 71.676
R1914 B.n307 B.n142 71.676
R1915 B.n303 B.n141 71.676
R1916 B.n299 B.n140 71.676
R1917 B.n295 B.n139 71.676
R1918 B.n291 B.n138 71.676
R1919 B.n287 B.n137 71.676
R1920 B.n283 B.n136 71.676
R1921 B.n279 B.n135 71.676
R1922 B.n275 B.n134 71.676
R1923 B.n271 B.n133 71.676
R1924 B.n267 B.n132 71.676
R1925 B.n263 B.n131 71.676
R1926 B.n259 B.n130 71.676
R1927 B.n255 B.n129 71.676
R1928 B.n251 B.n128 71.676
R1929 B.n247 B.n127 71.676
R1930 B.n243 B.n126 71.676
R1931 B.n239 B.n125 71.676
R1932 B.n235 B.n124 71.676
R1933 B.n231 B.n123 71.676
R1934 B.n227 B.n122 71.676
R1935 B.n223 B.n121 71.676
R1936 B.n219 B.n120 71.676
R1937 B.n215 B.n119 71.676
R1938 B.n211 B.n118 71.676
R1939 B.n207 B.n117 71.676
R1940 B.n203 B.n116 71.676
R1941 B.n199 B.n115 71.676
R1942 B.n195 B.n114 71.676
R1943 B.n191 B.n113 71.676
R1944 B.n187 B.n112 71.676
R1945 B.n183 B.n111 71.676
R1946 B.n179 B.n110 71.676
R1947 B.n175 B.n109 71.676
R1948 B.n171 B.n108 71.676
R1949 B.n167 B.n107 71.676
R1950 B.n163 B.n106 71.676
R1951 B.n159 B.n105 71.676
R1952 B.n502 B.n450 71.676
R1953 B.n506 B.n505 71.676
R1954 B.n511 B.n510 71.676
R1955 B.n514 B.n513 71.676
R1956 B.n519 B.n518 71.676
R1957 B.n522 B.n521 71.676
R1958 B.n527 B.n526 71.676
R1959 B.n530 B.n529 71.676
R1960 B.n535 B.n534 71.676
R1961 B.n538 B.n537 71.676
R1962 B.n543 B.n542 71.676
R1963 B.n546 B.n545 71.676
R1964 B.n551 B.n550 71.676
R1965 B.n554 B.n553 71.676
R1966 B.n559 B.n558 71.676
R1967 B.n562 B.n561 71.676
R1968 B.n567 B.n566 71.676
R1969 B.n570 B.n569 71.676
R1970 B.n575 B.n574 71.676
R1971 B.n578 B.n577 71.676
R1972 B.n586 B.n585 71.676
R1973 B.n589 B.n588 71.676
R1974 B.n594 B.n593 71.676
R1975 B.n597 B.n596 71.676
R1976 B.n602 B.n601 71.676
R1977 B.n605 B.n604 71.676
R1978 B.n611 B.n610 71.676
R1979 B.n614 B.n613 71.676
R1980 B.n619 B.n618 71.676
R1981 B.n622 B.n621 71.676
R1982 B.n627 B.n626 71.676
R1983 B.n630 B.n629 71.676
R1984 B.n635 B.n634 71.676
R1985 B.n638 B.n637 71.676
R1986 B.n643 B.n642 71.676
R1987 B.n646 B.n645 71.676
R1988 B.n651 B.n650 71.676
R1989 B.n654 B.n653 71.676
R1990 B.n659 B.n658 71.676
R1991 B.n662 B.n661 71.676
R1992 B.n667 B.n666 71.676
R1993 B.n670 B.n669 71.676
R1994 B.n675 B.n674 71.676
R1995 B.n678 B.n677 71.676
R1996 B.n683 B.n682 71.676
R1997 B.n686 B.n685 71.676
R1998 B.n503 B.n502 71.676
R1999 B.n505 B.n499 71.676
R2000 B.n512 B.n511 71.676
R2001 B.n513 B.n497 71.676
R2002 B.n520 B.n519 71.676
R2003 B.n521 B.n495 71.676
R2004 B.n528 B.n527 71.676
R2005 B.n529 B.n493 71.676
R2006 B.n536 B.n535 71.676
R2007 B.n537 B.n491 71.676
R2008 B.n544 B.n543 71.676
R2009 B.n545 B.n489 71.676
R2010 B.n552 B.n551 71.676
R2011 B.n553 B.n487 71.676
R2012 B.n560 B.n559 71.676
R2013 B.n561 B.n485 71.676
R2014 B.n568 B.n567 71.676
R2015 B.n569 B.n483 71.676
R2016 B.n576 B.n575 71.676
R2017 B.n577 B.n481 71.676
R2018 B.n587 B.n586 71.676
R2019 B.n588 B.n479 71.676
R2020 B.n595 B.n594 71.676
R2021 B.n596 B.n477 71.676
R2022 B.n603 B.n602 71.676
R2023 B.n604 B.n473 71.676
R2024 B.n612 B.n611 71.676
R2025 B.n613 B.n471 71.676
R2026 B.n620 B.n619 71.676
R2027 B.n621 B.n469 71.676
R2028 B.n628 B.n627 71.676
R2029 B.n629 B.n467 71.676
R2030 B.n636 B.n635 71.676
R2031 B.n637 B.n465 71.676
R2032 B.n644 B.n643 71.676
R2033 B.n645 B.n463 71.676
R2034 B.n652 B.n651 71.676
R2035 B.n653 B.n461 71.676
R2036 B.n660 B.n659 71.676
R2037 B.n661 B.n459 71.676
R2038 B.n668 B.n667 71.676
R2039 B.n669 B.n457 71.676
R2040 B.n676 B.n675 71.676
R2041 B.n677 B.n455 71.676
R2042 B.n684 B.n683 71.676
R2043 B.n687 B.n686 71.676
R2044 B.n1051 B.n1050 71.676
R2045 B.n1051 B.n2 71.676
R2046 B.n692 B.n451 68.5344
R2047 B.n936 B.n935 68.5344
R2048 B.n157 B.n156 59.5399
R2049 B.n154 B.n153 59.5399
R2050 B.n607 B.n475 59.5399
R2051 B.n583 B.n582 59.5399
R2052 B.n156 B.n155 52.946
R2053 B.n153 B.n152 52.946
R2054 B.n475 B.n474 52.946
R2055 B.n582 B.n581 52.946
R2056 B.n692 B.n447 42.7556
R2057 B.n698 B.n447 42.7556
R2058 B.n698 B.n443 42.7556
R2059 B.n704 B.n443 42.7556
R2060 B.n704 B.n438 42.7556
R2061 B.n710 B.n438 42.7556
R2062 B.n710 B.n439 42.7556
R2063 B.n716 B.n431 42.7556
R2064 B.n722 B.n431 42.7556
R2065 B.n722 B.n427 42.7556
R2066 B.n728 B.n427 42.7556
R2067 B.n728 B.n423 42.7556
R2068 B.n734 B.n423 42.7556
R2069 B.n734 B.n419 42.7556
R2070 B.n740 B.n419 42.7556
R2071 B.n740 B.n415 42.7556
R2072 B.n746 B.n415 42.7556
R2073 B.n752 B.n411 42.7556
R2074 B.n752 B.n407 42.7556
R2075 B.n758 B.n407 42.7556
R2076 B.n758 B.n403 42.7556
R2077 B.n764 B.n403 42.7556
R2078 B.n764 B.n399 42.7556
R2079 B.n770 B.n399 42.7556
R2080 B.n776 B.n395 42.7556
R2081 B.n776 B.n391 42.7556
R2082 B.n782 B.n391 42.7556
R2083 B.n782 B.n387 42.7556
R2084 B.n788 B.n387 42.7556
R2085 B.n788 B.n383 42.7556
R2086 B.n794 B.n383 42.7556
R2087 B.n800 B.n379 42.7556
R2088 B.n800 B.n375 42.7556
R2089 B.n806 B.n375 42.7556
R2090 B.n806 B.n371 42.7556
R2091 B.n812 B.n371 42.7556
R2092 B.n812 B.n367 42.7556
R2093 B.n818 B.n367 42.7556
R2094 B.n824 B.n363 42.7556
R2095 B.n824 B.n359 42.7556
R2096 B.n830 B.n359 42.7556
R2097 B.n830 B.n355 42.7556
R2098 B.n836 B.n355 42.7556
R2099 B.n836 B.n351 42.7556
R2100 B.n842 B.n351 42.7556
R2101 B.n849 B.n347 42.7556
R2102 B.n849 B.n343 42.7556
R2103 B.n855 B.n343 42.7556
R2104 B.n855 B.n4 42.7556
R2105 B.n1049 B.n4 42.7556
R2106 B.n1049 B.n1048 42.7556
R2107 B.n1048 B.n1047 42.7556
R2108 B.n1047 B.n8 42.7556
R2109 B.n12 B.n8 42.7556
R2110 B.n1040 B.n12 42.7556
R2111 B.n1040 B.n1039 42.7556
R2112 B.n1038 B.n16 42.7556
R2113 B.n1032 B.n16 42.7556
R2114 B.n1032 B.n1031 42.7556
R2115 B.n1031 B.n1030 42.7556
R2116 B.n1030 B.n23 42.7556
R2117 B.n1024 B.n23 42.7556
R2118 B.n1024 B.n1023 42.7556
R2119 B.n1022 B.n30 42.7556
R2120 B.n1016 B.n30 42.7556
R2121 B.n1016 B.n1015 42.7556
R2122 B.n1015 B.n1014 42.7556
R2123 B.n1014 B.n37 42.7556
R2124 B.n1008 B.n37 42.7556
R2125 B.n1008 B.n1007 42.7556
R2126 B.n1006 B.n44 42.7556
R2127 B.n1000 B.n44 42.7556
R2128 B.n1000 B.n999 42.7556
R2129 B.n999 B.n998 42.7556
R2130 B.n998 B.n51 42.7556
R2131 B.n992 B.n51 42.7556
R2132 B.n992 B.n991 42.7556
R2133 B.n990 B.n58 42.7556
R2134 B.n984 B.n58 42.7556
R2135 B.n984 B.n983 42.7556
R2136 B.n983 B.n982 42.7556
R2137 B.n982 B.n65 42.7556
R2138 B.n976 B.n65 42.7556
R2139 B.n976 B.n975 42.7556
R2140 B.n974 B.n72 42.7556
R2141 B.n968 B.n72 42.7556
R2142 B.n968 B.n967 42.7556
R2143 B.n967 B.n966 42.7556
R2144 B.n966 B.n79 42.7556
R2145 B.n960 B.n79 42.7556
R2146 B.n960 B.n959 42.7556
R2147 B.n959 B.n958 42.7556
R2148 B.n958 B.n86 42.7556
R2149 B.n952 B.n86 42.7556
R2150 B.n951 B.n950 42.7556
R2151 B.n950 B.n93 42.7556
R2152 B.n944 B.n93 42.7556
R2153 B.n944 B.n943 42.7556
R2154 B.n943 B.n942 42.7556
R2155 B.n942 B.n100 42.7556
R2156 B.n936 B.n100 42.7556
R2157 B.n842 B.t3 37.7256
R2158 B.t6 B.n1038 37.7256
R2159 B.n818 B.t9 36.4681
R2160 B.t7 B.n1022 36.4681
R2161 B.n794 B.t2 35.2106
R2162 B.t8 B.n1006 35.2106
R2163 B.n770 B.t1 33.9531
R2164 B.t0 B.n990 33.9531
R2165 B.n746 B.t4 32.6956
R2166 B.t5 B.n974 32.6956
R2167 B.n694 B.n449 30.7517
R2168 B.n690 B.n689 30.7517
R2169 B.n932 B.n931 30.7517
R2170 B.n938 B.n102 30.7517
R2171 B.n439 B.t11 22.6355
R2172 B.t15 B.n951 22.6355
R2173 B.n716 B.t11 20.1205
R2174 B.n952 B.t15 20.1205
R2175 B B.n1052 18.0485
R2176 B.n695 B.n694 10.6151
R2177 B.n696 B.n695 10.6151
R2178 B.n696 B.n441 10.6151
R2179 B.n706 B.n441 10.6151
R2180 B.n707 B.n706 10.6151
R2181 B.n708 B.n707 10.6151
R2182 B.n708 B.n433 10.6151
R2183 B.n718 B.n433 10.6151
R2184 B.n719 B.n718 10.6151
R2185 B.n720 B.n719 10.6151
R2186 B.n720 B.n425 10.6151
R2187 B.n730 B.n425 10.6151
R2188 B.n731 B.n730 10.6151
R2189 B.n732 B.n731 10.6151
R2190 B.n732 B.n417 10.6151
R2191 B.n742 B.n417 10.6151
R2192 B.n743 B.n742 10.6151
R2193 B.n744 B.n743 10.6151
R2194 B.n744 B.n409 10.6151
R2195 B.n754 B.n409 10.6151
R2196 B.n755 B.n754 10.6151
R2197 B.n756 B.n755 10.6151
R2198 B.n756 B.n401 10.6151
R2199 B.n766 B.n401 10.6151
R2200 B.n767 B.n766 10.6151
R2201 B.n768 B.n767 10.6151
R2202 B.n768 B.n393 10.6151
R2203 B.n778 B.n393 10.6151
R2204 B.n779 B.n778 10.6151
R2205 B.n780 B.n779 10.6151
R2206 B.n780 B.n385 10.6151
R2207 B.n790 B.n385 10.6151
R2208 B.n791 B.n790 10.6151
R2209 B.n792 B.n791 10.6151
R2210 B.n792 B.n377 10.6151
R2211 B.n802 B.n377 10.6151
R2212 B.n803 B.n802 10.6151
R2213 B.n804 B.n803 10.6151
R2214 B.n804 B.n369 10.6151
R2215 B.n814 B.n369 10.6151
R2216 B.n815 B.n814 10.6151
R2217 B.n816 B.n815 10.6151
R2218 B.n816 B.n361 10.6151
R2219 B.n826 B.n361 10.6151
R2220 B.n827 B.n826 10.6151
R2221 B.n828 B.n827 10.6151
R2222 B.n828 B.n353 10.6151
R2223 B.n838 B.n353 10.6151
R2224 B.n839 B.n838 10.6151
R2225 B.n840 B.n839 10.6151
R2226 B.n840 B.n345 10.6151
R2227 B.n851 B.n345 10.6151
R2228 B.n852 B.n851 10.6151
R2229 B.n853 B.n852 10.6151
R2230 B.n853 B.n0 10.6151
R2231 B.n501 B.n449 10.6151
R2232 B.n501 B.n500 10.6151
R2233 B.n507 B.n500 10.6151
R2234 B.n508 B.n507 10.6151
R2235 B.n509 B.n508 10.6151
R2236 B.n509 B.n498 10.6151
R2237 B.n515 B.n498 10.6151
R2238 B.n516 B.n515 10.6151
R2239 B.n517 B.n516 10.6151
R2240 B.n517 B.n496 10.6151
R2241 B.n523 B.n496 10.6151
R2242 B.n524 B.n523 10.6151
R2243 B.n525 B.n524 10.6151
R2244 B.n525 B.n494 10.6151
R2245 B.n531 B.n494 10.6151
R2246 B.n532 B.n531 10.6151
R2247 B.n533 B.n532 10.6151
R2248 B.n533 B.n492 10.6151
R2249 B.n539 B.n492 10.6151
R2250 B.n540 B.n539 10.6151
R2251 B.n541 B.n540 10.6151
R2252 B.n541 B.n490 10.6151
R2253 B.n547 B.n490 10.6151
R2254 B.n548 B.n547 10.6151
R2255 B.n549 B.n548 10.6151
R2256 B.n549 B.n488 10.6151
R2257 B.n555 B.n488 10.6151
R2258 B.n556 B.n555 10.6151
R2259 B.n557 B.n556 10.6151
R2260 B.n557 B.n486 10.6151
R2261 B.n563 B.n486 10.6151
R2262 B.n564 B.n563 10.6151
R2263 B.n565 B.n564 10.6151
R2264 B.n565 B.n484 10.6151
R2265 B.n571 B.n484 10.6151
R2266 B.n572 B.n571 10.6151
R2267 B.n573 B.n572 10.6151
R2268 B.n573 B.n482 10.6151
R2269 B.n579 B.n482 10.6151
R2270 B.n580 B.n579 10.6151
R2271 B.n584 B.n580 10.6151
R2272 B.n590 B.n480 10.6151
R2273 B.n591 B.n590 10.6151
R2274 B.n592 B.n591 10.6151
R2275 B.n592 B.n478 10.6151
R2276 B.n598 B.n478 10.6151
R2277 B.n599 B.n598 10.6151
R2278 B.n600 B.n599 10.6151
R2279 B.n600 B.n476 10.6151
R2280 B.n606 B.n476 10.6151
R2281 B.n609 B.n608 10.6151
R2282 B.n609 B.n472 10.6151
R2283 B.n615 B.n472 10.6151
R2284 B.n616 B.n615 10.6151
R2285 B.n617 B.n616 10.6151
R2286 B.n617 B.n470 10.6151
R2287 B.n623 B.n470 10.6151
R2288 B.n624 B.n623 10.6151
R2289 B.n625 B.n624 10.6151
R2290 B.n625 B.n468 10.6151
R2291 B.n631 B.n468 10.6151
R2292 B.n632 B.n631 10.6151
R2293 B.n633 B.n632 10.6151
R2294 B.n633 B.n466 10.6151
R2295 B.n639 B.n466 10.6151
R2296 B.n640 B.n639 10.6151
R2297 B.n641 B.n640 10.6151
R2298 B.n641 B.n464 10.6151
R2299 B.n647 B.n464 10.6151
R2300 B.n648 B.n647 10.6151
R2301 B.n649 B.n648 10.6151
R2302 B.n649 B.n462 10.6151
R2303 B.n655 B.n462 10.6151
R2304 B.n656 B.n655 10.6151
R2305 B.n657 B.n656 10.6151
R2306 B.n657 B.n460 10.6151
R2307 B.n663 B.n460 10.6151
R2308 B.n664 B.n663 10.6151
R2309 B.n665 B.n664 10.6151
R2310 B.n665 B.n458 10.6151
R2311 B.n671 B.n458 10.6151
R2312 B.n672 B.n671 10.6151
R2313 B.n673 B.n672 10.6151
R2314 B.n673 B.n456 10.6151
R2315 B.n679 B.n456 10.6151
R2316 B.n680 B.n679 10.6151
R2317 B.n681 B.n680 10.6151
R2318 B.n681 B.n454 10.6151
R2319 B.n454 B.n453 10.6151
R2320 B.n688 B.n453 10.6151
R2321 B.n689 B.n688 10.6151
R2322 B.n690 B.n445 10.6151
R2323 B.n700 B.n445 10.6151
R2324 B.n701 B.n700 10.6151
R2325 B.n702 B.n701 10.6151
R2326 B.n702 B.n436 10.6151
R2327 B.n712 B.n436 10.6151
R2328 B.n713 B.n712 10.6151
R2329 B.n714 B.n713 10.6151
R2330 B.n714 B.n429 10.6151
R2331 B.n724 B.n429 10.6151
R2332 B.n725 B.n724 10.6151
R2333 B.n726 B.n725 10.6151
R2334 B.n726 B.n421 10.6151
R2335 B.n736 B.n421 10.6151
R2336 B.n737 B.n736 10.6151
R2337 B.n738 B.n737 10.6151
R2338 B.n738 B.n413 10.6151
R2339 B.n748 B.n413 10.6151
R2340 B.n749 B.n748 10.6151
R2341 B.n750 B.n749 10.6151
R2342 B.n750 B.n405 10.6151
R2343 B.n760 B.n405 10.6151
R2344 B.n761 B.n760 10.6151
R2345 B.n762 B.n761 10.6151
R2346 B.n762 B.n397 10.6151
R2347 B.n772 B.n397 10.6151
R2348 B.n773 B.n772 10.6151
R2349 B.n774 B.n773 10.6151
R2350 B.n774 B.n389 10.6151
R2351 B.n784 B.n389 10.6151
R2352 B.n785 B.n784 10.6151
R2353 B.n786 B.n785 10.6151
R2354 B.n786 B.n381 10.6151
R2355 B.n796 B.n381 10.6151
R2356 B.n797 B.n796 10.6151
R2357 B.n798 B.n797 10.6151
R2358 B.n798 B.n373 10.6151
R2359 B.n808 B.n373 10.6151
R2360 B.n809 B.n808 10.6151
R2361 B.n810 B.n809 10.6151
R2362 B.n810 B.n365 10.6151
R2363 B.n820 B.n365 10.6151
R2364 B.n821 B.n820 10.6151
R2365 B.n822 B.n821 10.6151
R2366 B.n822 B.n357 10.6151
R2367 B.n832 B.n357 10.6151
R2368 B.n833 B.n832 10.6151
R2369 B.n834 B.n833 10.6151
R2370 B.n834 B.n349 10.6151
R2371 B.n844 B.n349 10.6151
R2372 B.n845 B.n844 10.6151
R2373 B.n847 B.n845 10.6151
R2374 B.n847 B.n846 10.6151
R2375 B.n846 B.n341 10.6151
R2376 B.n858 B.n341 10.6151
R2377 B.n859 B.n858 10.6151
R2378 B.n860 B.n859 10.6151
R2379 B.n861 B.n860 10.6151
R2380 B.n862 B.n861 10.6151
R2381 B.n865 B.n862 10.6151
R2382 B.n866 B.n865 10.6151
R2383 B.n867 B.n866 10.6151
R2384 B.n868 B.n867 10.6151
R2385 B.n870 B.n868 10.6151
R2386 B.n871 B.n870 10.6151
R2387 B.n872 B.n871 10.6151
R2388 B.n873 B.n872 10.6151
R2389 B.n875 B.n873 10.6151
R2390 B.n876 B.n875 10.6151
R2391 B.n877 B.n876 10.6151
R2392 B.n878 B.n877 10.6151
R2393 B.n880 B.n878 10.6151
R2394 B.n881 B.n880 10.6151
R2395 B.n882 B.n881 10.6151
R2396 B.n883 B.n882 10.6151
R2397 B.n885 B.n883 10.6151
R2398 B.n886 B.n885 10.6151
R2399 B.n887 B.n886 10.6151
R2400 B.n888 B.n887 10.6151
R2401 B.n890 B.n888 10.6151
R2402 B.n891 B.n890 10.6151
R2403 B.n892 B.n891 10.6151
R2404 B.n893 B.n892 10.6151
R2405 B.n895 B.n893 10.6151
R2406 B.n896 B.n895 10.6151
R2407 B.n897 B.n896 10.6151
R2408 B.n898 B.n897 10.6151
R2409 B.n900 B.n898 10.6151
R2410 B.n901 B.n900 10.6151
R2411 B.n902 B.n901 10.6151
R2412 B.n903 B.n902 10.6151
R2413 B.n905 B.n903 10.6151
R2414 B.n906 B.n905 10.6151
R2415 B.n907 B.n906 10.6151
R2416 B.n908 B.n907 10.6151
R2417 B.n910 B.n908 10.6151
R2418 B.n911 B.n910 10.6151
R2419 B.n912 B.n911 10.6151
R2420 B.n913 B.n912 10.6151
R2421 B.n915 B.n913 10.6151
R2422 B.n916 B.n915 10.6151
R2423 B.n917 B.n916 10.6151
R2424 B.n918 B.n917 10.6151
R2425 B.n920 B.n918 10.6151
R2426 B.n921 B.n920 10.6151
R2427 B.n922 B.n921 10.6151
R2428 B.n923 B.n922 10.6151
R2429 B.n925 B.n923 10.6151
R2430 B.n926 B.n925 10.6151
R2431 B.n927 B.n926 10.6151
R2432 B.n928 B.n927 10.6151
R2433 B.n930 B.n928 10.6151
R2434 B.n931 B.n930 10.6151
R2435 B.n1044 B.n1 10.6151
R2436 B.n1044 B.n1043 10.6151
R2437 B.n1043 B.n1042 10.6151
R2438 B.n1042 B.n10 10.6151
R2439 B.n1036 B.n10 10.6151
R2440 B.n1036 B.n1035 10.6151
R2441 B.n1035 B.n1034 10.6151
R2442 B.n1034 B.n18 10.6151
R2443 B.n1028 B.n18 10.6151
R2444 B.n1028 B.n1027 10.6151
R2445 B.n1027 B.n1026 10.6151
R2446 B.n1026 B.n25 10.6151
R2447 B.n1020 B.n25 10.6151
R2448 B.n1020 B.n1019 10.6151
R2449 B.n1019 B.n1018 10.6151
R2450 B.n1018 B.n32 10.6151
R2451 B.n1012 B.n32 10.6151
R2452 B.n1012 B.n1011 10.6151
R2453 B.n1011 B.n1010 10.6151
R2454 B.n1010 B.n39 10.6151
R2455 B.n1004 B.n39 10.6151
R2456 B.n1004 B.n1003 10.6151
R2457 B.n1003 B.n1002 10.6151
R2458 B.n1002 B.n46 10.6151
R2459 B.n996 B.n46 10.6151
R2460 B.n996 B.n995 10.6151
R2461 B.n995 B.n994 10.6151
R2462 B.n994 B.n53 10.6151
R2463 B.n988 B.n53 10.6151
R2464 B.n988 B.n987 10.6151
R2465 B.n987 B.n986 10.6151
R2466 B.n986 B.n60 10.6151
R2467 B.n980 B.n60 10.6151
R2468 B.n980 B.n979 10.6151
R2469 B.n979 B.n978 10.6151
R2470 B.n978 B.n67 10.6151
R2471 B.n972 B.n67 10.6151
R2472 B.n972 B.n971 10.6151
R2473 B.n971 B.n970 10.6151
R2474 B.n970 B.n74 10.6151
R2475 B.n964 B.n74 10.6151
R2476 B.n964 B.n963 10.6151
R2477 B.n963 B.n962 10.6151
R2478 B.n962 B.n81 10.6151
R2479 B.n956 B.n81 10.6151
R2480 B.n956 B.n955 10.6151
R2481 B.n955 B.n954 10.6151
R2482 B.n954 B.n88 10.6151
R2483 B.n948 B.n88 10.6151
R2484 B.n948 B.n947 10.6151
R2485 B.n947 B.n946 10.6151
R2486 B.n946 B.n95 10.6151
R2487 B.n940 B.n95 10.6151
R2488 B.n940 B.n939 10.6151
R2489 B.n939 B.n938 10.6151
R2490 B.n158 B.n102 10.6151
R2491 B.n161 B.n158 10.6151
R2492 B.n162 B.n161 10.6151
R2493 B.n165 B.n162 10.6151
R2494 B.n166 B.n165 10.6151
R2495 B.n169 B.n166 10.6151
R2496 B.n170 B.n169 10.6151
R2497 B.n173 B.n170 10.6151
R2498 B.n174 B.n173 10.6151
R2499 B.n177 B.n174 10.6151
R2500 B.n178 B.n177 10.6151
R2501 B.n181 B.n178 10.6151
R2502 B.n182 B.n181 10.6151
R2503 B.n185 B.n182 10.6151
R2504 B.n186 B.n185 10.6151
R2505 B.n189 B.n186 10.6151
R2506 B.n190 B.n189 10.6151
R2507 B.n193 B.n190 10.6151
R2508 B.n194 B.n193 10.6151
R2509 B.n197 B.n194 10.6151
R2510 B.n198 B.n197 10.6151
R2511 B.n201 B.n198 10.6151
R2512 B.n202 B.n201 10.6151
R2513 B.n205 B.n202 10.6151
R2514 B.n206 B.n205 10.6151
R2515 B.n209 B.n206 10.6151
R2516 B.n210 B.n209 10.6151
R2517 B.n213 B.n210 10.6151
R2518 B.n214 B.n213 10.6151
R2519 B.n217 B.n214 10.6151
R2520 B.n218 B.n217 10.6151
R2521 B.n221 B.n218 10.6151
R2522 B.n222 B.n221 10.6151
R2523 B.n225 B.n222 10.6151
R2524 B.n226 B.n225 10.6151
R2525 B.n229 B.n226 10.6151
R2526 B.n230 B.n229 10.6151
R2527 B.n233 B.n230 10.6151
R2528 B.n234 B.n233 10.6151
R2529 B.n237 B.n234 10.6151
R2530 B.n238 B.n237 10.6151
R2531 B.n242 B.n241 10.6151
R2532 B.n245 B.n242 10.6151
R2533 B.n246 B.n245 10.6151
R2534 B.n249 B.n246 10.6151
R2535 B.n250 B.n249 10.6151
R2536 B.n253 B.n250 10.6151
R2537 B.n254 B.n253 10.6151
R2538 B.n257 B.n254 10.6151
R2539 B.n258 B.n257 10.6151
R2540 B.n262 B.n261 10.6151
R2541 B.n265 B.n262 10.6151
R2542 B.n266 B.n265 10.6151
R2543 B.n269 B.n266 10.6151
R2544 B.n270 B.n269 10.6151
R2545 B.n273 B.n270 10.6151
R2546 B.n274 B.n273 10.6151
R2547 B.n277 B.n274 10.6151
R2548 B.n278 B.n277 10.6151
R2549 B.n281 B.n278 10.6151
R2550 B.n282 B.n281 10.6151
R2551 B.n285 B.n282 10.6151
R2552 B.n286 B.n285 10.6151
R2553 B.n289 B.n286 10.6151
R2554 B.n290 B.n289 10.6151
R2555 B.n293 B.n290 10.6151
R2556 B.n294 B.n293 10.6151
R2557 B.n297 B.n294 10.6151
R2558 B.n298 B.n297 10.6151
R2559 B.n301 B.n298 10.6151
R2560 B.n302 B.n301 10.6151
R2561 B.n305 B.n302 10.6151
R2562 B.n306 B.n305 10.6151
R2563 B.n309 B.n306 10.6151
R2564 B.n310 B.n309 10.6151
R2565 B.n313 B.n310 10.6151
R2566 B.n314 B.n313 10.6151
R2567 B.n317 B.n314 10.6151
R2568 B.n318 B.n317 10.6151
R2569 B.n321 B.n318 10.6151
R2570 B.n322 B.n321 10.6151
R2571 B.n325 B.n322 10.6151
R2572 B.n326 B.n325 10.6151
R2573 B.n329 B.n326 10.6151
R2574 B.n330 B.n329 10.6151
R2575 B.n333 B.n330 10.6151
R2576 B.n334 B.n333 10.6151
R2577 B.n337 B.n334 10.6151
R2578 B.n339 B.n337 10.6151
R2579 B.n340 B.n339 10.6151
R2580 B.n932 B.n340 10.6151
R2581 B.t4 B.n411 10.0605
R2582 B.n975 B.t5 10.0605
R2583 B.n584 B.n583 9.36635
R2584 B.n608 B.n607 9.36635
R2585 B.n238 B.n157 9.36635
R2586 B.n261 B.n154 9.36635
R2587 B.t1 B.n395 8.80302
R2588 B.n991 B.t0 8.80302
R2589 B.n1052 B.n0 8.11757
R2590 B.n1052 B.n1 8.11757
R2591 B.t2 B.n379 7.54551
R2592 B.n1007 B.t8 7.54551
R2593 B.t9 B.n363 6.28801
R2594 B.n1023 B.t7 6.28801
R2595 B.t3 B.n347 5.03051
R2596 B.n1039 B.t6 5.03051
R2597 B.n583 B.n480 1.24928
R2598 B.n607 B.n606 1.24928
R2599 B.n241 B.n157 1.24928
R2600 B.n258 B.n154 1.24928
R2601 VN.n73 VN.n38 161.3
R2602 VN.n72 VN.n71 161.3
R2603 VN.n70 VN.n39 161.3
R2604 VN.n69 VN.n68 161.3
R2605 VN.n67 VN.n40 161.3
R2606 VN.n66 VN.n65 161.3
R2607 VN.n64 VN.n63 161.3
R2608 VN.n62 VN.n42 161.3
R2609 VN.n61 VN.n60 161.3
R2610 VN.n59 VN.n43 161.3
R2611 VN.n58 VN.n57 161.3
R2612 VN.n55 VN.n44 161.3
R2613 VN.n54 VN.n53 161.3
R2614 VN.n52 VN.n45 161.3
R2615 VN.n51 VN.n50 161.3
R2616 VN.n49 VN.n46 161.3
R2617 VN.n35 VN.n0 161.3
R2618 VN.n34 VN.n33 161.3
R2619 VN.n32 VN.n1 161.3
R2620 VN.n31 VN.n30 161.3
R2621 VN.n29 VN.n2 161.3
R2622 VN.n28 VN.n27 161.3
R2623 VN.n26 VN.n25 161.3
R2624 VN.n24 VN.n4 161.3
R2625 VN.n23 VN.n22 161.3
R2626 VN.n21 VN.n5 161.3
R2627 VN.n20 VN.n19 161.3
R2628 VN.n17 VN.n6 161.3
R2629 VN.n16 VN.n15 161.3
R2630 VN.n14 VN.n7 161.3
R2631 VN.n13 VN.n12 161.3
R2632 VN.n11 VN.n8 161.3
R2633 VN.n9 VN.t4 156.357
R2634 VN.n47 VN.t7 156.357
R2635 VN.n10 VN.t2 122.71
R2636 VN.n18 VN.t9 122.71
R2637 VN.n3 VN.t8 122.71
R2638 VN.n36 VN.t5 122.71
R2639 VN.n48 VN.t3 122.71
R2640 VN.n56 VN.t0 122.71
R2641 VN.n41 VN.t6 122.71
R2642 VN.n74 VN.t1 122.71
R2643 VN.n37 VN.n36 100.382
R2644 VN.n75 VN.n74 100.382
R2645 VN.n30 VN.n1 55.5035
R2646 VN.n68 VN.n39 55.5035
R2647 VN VN.n75 52.4489
R2648 VN.n12 VN.n7 51.6086
R2649 VN.n24 VN.n23 51.6086
R2650 VN.n50 VN.n45 51.6086
R2651 VN.n62 VN.n61 51.6086
R2652 VN.n10 VN.n9 48.8439
R2653 VN.n48 VN.n47 48.8439
R2654 VN.n16 VN.n7 29.2126
R2655 VN.n23 VN.n5 29.2126
R2656 VN.n54 VN.n45 29.2126
R2657 VN.n61 VN.n43 29.2126
R2658 VN.n34 VN.n1 25.3177
R2659 VN.n72 VN.n39 25.3177
R2660 VN.n12 VN.n11 24.3439
R2661 VN.n17 VN.n16 24.3439
R2662 VN.n19 VN.n5 24.3439
R2663 VN.n25 VN.n24 24.3439
R2664 VN.n29 VN.n28 24.3439
R2665 VN.n30 VN.n29 24.3439
R2666 VN.n35 VN.n34 24.3439
R2667 VN.n50 VN.n49 24.3439
R2668 VN.n57 VN.n43 24.3439
R2669 VN.n55 VN.n54 24.3439
R2670 VN.n68 VN.n67 24.3439
R2671 VN.n67 VN.n66 24.3439
R2672 VN.n63 VN.n62 24.3439
R2673 VN.n73 VN.n72 24.3439
R2674 VN.n11 VN.n10 23.3702
R2675 VN.n25 VN.n3 23.3702
R2676 VN.n49 VN.n48 23.3702
R2677 VN.n63 VN.n41 23.3702
R2678 VN.n18 VN.n17 12.1722
R2679 VN.n19 VN.n18 12.1722
R2680 VN.n57 VN.n56 12.1722
R2681 VN.n56 VN.n55 12.1722
R2682 VN.n36 VN.n35 10.2247
R2683 VN.n74 VN.n73 10.2247
R2684 VN.n47 VN.n46 6.8468
R2685 VN.n9 VN.n8 6.8468
R2686 VN.n28 VN.n3 0.974237
R2687 VN.n66 VN.n41 0.974237
R2688 VN.n75 VN.n38 0.278398
R2689 VN.n37 VN.n0 0.278398
R2690 VN.n71 VN.n38 0.189894
R2691 VN.n71 VN.n70 0.189894
R2692 VN.n70 VN.n69 0.189894
R2693 VN.n69 VN.n40 0.189894
R2694 VN.n65 VN.n40 0.189894
R2695 VN.n65 VN.n64 0.189894
R2696 VN.n64 VN.n42 0.189894
R2697 VN.n60 VN.n42 0.189894
R2698 VN.n60 VN.n59 0.189894
R2699 VN.n59 VN.n58 0.189894
R2700 VN.n58 VN.n44 0.189894
R2701 VN.n53 VN.n44 0.189894
R2702 VN.n53 VN.n52 0.189894
R2703 VN.n52 VN.n51 0.189894
R2704 VN.n51 VN.n46 0.189894
R2705 VN.n13 VN.n8 0.189894
R2706 VN.n14 VN.n13 0.189894
R2707 VN.n15 VN.n14 0.189894
R2708 VN.n15 VN.n6 0.189894
R2709 VN.n20 VN.n6 0.189894
R2710 VN.n21 VN.n20 0.189894
R2711 VN.n22 VN.n21 0.189894
R2712 VN.n22 VN.n4 0.189894
R2713 VN.n26 VN.n4 0.189894
R2714 VN.n27 VN.n26 0.189894
R2715 VN.n27 VN.n2 0.189894
R2716 VN.n31 VN.n2 0.189894
R2717 VN.n32 VN.n31 0.189894
R2718 VN.n33 VN.n32 0.189894
R2719 VN.n33 VN.n0 0.189894
R2720 VN VN.n37 0.153422
R2721 VDD2.n129 VDD2.n69 289.615
R2722 VDD2.n60 VDD2.n0 289.615
R2723 VDD2.n130 VDD2.n129 185
R2724 VDD2.n128 VDD2.n127 185
R2725 VDD2.n73 VDD2.n72 185
R2726 VDD2.n122 VDD2.n121 185
R2727 VDD2.n120 VDD2.n119 185
R2728 VDD2.n77 VDD2.n76 185
R2729 VDD2.n114 VDD2.n113 185
R2730 VDD2.n112 VDD2.n79 185
R2731 VDD2.n111 VDD2.n110 185
R2732 VDD2.n82 VDD2.n80 185
R2733 VDD2.n105 VDD2.n104 185
R2734 VDD2.n103 VDD2.n102 185
R2735 VDD2.n86 VDD2.n85 185
R2736 VDD2.n97 VDD2.n96 185
R2737 VDD2.n95 VDD2.n94 185
R2738 VDD2.n90 VDD2.n89 185
R2739 VDD2.n20 VDD2.n19 185
R2740 VDD2.n25 VDD2.n24 185
R2741 VDD2.n27 VDD2.n26 185
R2742 VDD2.n16 VDD2.n15 185
R2743 VDD2.n33 VDD2.n32 185
R2744 VDD2.n35 VDD2.n34 185
R2745 VDD2.n12 VDD2.n11 185
R2746 VDD2.n42 VDD2.n41 185
R2747 VDD2.n43 VDD2.n10 185
R2748 VDD2.n45 VDD2.n44 185
R2749 VDD2.n8 VDD2.n7 185
R2750 VDD2.n51 VDD2.n50 185
R2751 VDD2.n53 VDD2.n52 185
R2752 VDD2.n4 VDD2.n3 185
R2753 VDD2.n59 VDD2.n58 185
R2754 VDD2.n61 VDD2.n60 185
R2755 VDD2.n91 VDD2.t8 149.524
R2756 VDD2.n21 VDD2.t5 149.524
R2757 VDD2.n129 VDD2.n128 104.615
R2758 VDD2.n128 VDD2.n72 104.615
R2759 VDD2.n121 VDD2.n72 104.615
R2760 VDD2.n121 VDD2.n120 104.615
R2761 VDD2.n120 VDD2.n76 104.615
R2762 VDD2.n113 VDD2.n76 104.615
R2763 VDD2.n113 VDD2.n112 104.615
R2764 VDD2.n112 VDD2.n111 104.615
R2765 VDD2.n111 VDD2.n80 104.615
R2766 VDD2.n104 VDD2.n80 104.615
R2767 VDD2.n104 VDD2.n103 104.615
R2768 VDD2.n103 VDD2.n85 104.615
R2769 VDD2.n96 VDD2.n85 104.615
R2770 VDD2.n96 VDD2.n95 104.615
R2771 VDD2.n95 VDD2.n89 104.615
R2772 VDD2.n25 VDD2.n19 104.615
R2773 VDD2.n26 VDD2.n25 104.615
R2774 VDD2.n26 VDD2.n15 104.615
R2775 VDD2.n33 VDD2.n15 104.615
R2776 VDD2.n34 VDD2.n33 104.615
R2777 VDD2.n34 VDD2.n11 104.615
R2778 VDD2.n42 VDD2.n11 104.615
R2779 VDD2.n43 VDD2.n42 104.615
R2780 VDD2.n44 VDD2.n43 104.615
R2781 VDD2.n44 VDD2.n7 104.615
R2782 VDD2.n51 VDD2.n7 104.615
R2783 VDD2.n52 VDD2.n51 104.615
R2784 VDD2.n52 VDD2.n3 104.615
R2785 VDD2.n59 VDD2.n3 104.615
R2786 VDD2.n60 VDD2.n59 104.615
R2787 VDD2.n68 VDD2.n67 65.5289
R2788 VDD2 VDD2.n137 65.5261
R2789 VDD2.n136 VDD2.n135 63.8193
R2790 VDD2.n66 VDD2.n65 63.8192
R2791 VDD2.n66 VDD2.n64 53.157
R2792 VDD2.t8 VDD2.n89 52.3082
R2793 VDD2.t5 VDD2.n19 52.3082
R2794 VDD2.n134 VDD2.n133 50.8035
R2795 VDD2.n134 VDD2.n68 45.4287
R2796 VDD2.n114 VDD2.n79 13.1884
R2797 VDD2.n45 VDD2.n10 13.1884
R2798 VDD2.n115 VDD2.n77 12.8005
R2799 VDD2.n110 VDD2.n81 12.8005
R2800 VDD2.n41 VDD2.n40 12.8005
R2801 VDD2.n46 VDD2.n8 12.8005
R2802 VDD2.n119 VDD2.n118 12.0247
R2803 VDD2.n109 VDD2.n82 12.0247
R2804 VDD2.n39 VDD2.n12 12.0247
R2805 VDD2.n50 VDD2.n49 12.0247
R2806 VDD2.n122 VDD2.n75 11.249
R2807 VDD2.n106 VDD2.n105 11.249
R2808 VDD2.n36 VDD2.n35 11.249
R2809 VDD2.n53 VDD2.n6 11.249
R2810 VDD2.n123 VDD2.n73 10.4732
R2811 VDD2.n102 VDD2.n84 10.4732
R2812 VDD2.n32 VDD2.n14 10.4732
R2813 VDD2.n54 VDD2.n4 10.4732
R2814 VDD2.n91 VDD2.n90 10.2747
R2815 VDD2.n21 VDD2.n20 10.2747
R2816 VDD2.n127 VDD2.n126 9.69747
R2817 VDD2.n101 VDD2.n86 9.69747
R2818 VDD2.n31 VDD2.n16 9.69747
R2819 VDD2.n58 VDD2.n57 9.69747
R2820 VDD2.n133 VDD2.n132 9.45567
R2821 VDD2.n64 VDD2.n63 9.45567
R2822 VDD2.n93 VDD2.n92 9.3005
R2823 VDD2.n88 VDD2.n87 9.3005
R2824 VDD2.n99 VDD2.n98 9.3005
R2825 VDD2.n101 VDD2.n100 9.3005
R2826 VDD2.n84 VDD2.n83 9.3005
R2827 VDD2.n107 VDD2.n106 9.3005
R2828 VDD2.n109 VDD2.n108 9.3005
R2829 VDD2.n81 VDD2.n78 9.3005
R2830 VDD2.n132 VDD2.n131 9.3005
R2831 VDD2.n71 VDD2.n70 9.3005
R2832 VDD2.n126 VDD2.n125 9.3005
R2833 VDD2.n124 VDD2.n123 9.3005
R2834 VDD2.n75 VDD2.n74 9.3005
R2835 VDD2.n118 VDD2.n117 9.3005
R2836 VDD2.n116 VDD2.n115 9.3005
R2837 VDD2.n63 VDD2.n62 9.3005
R2838 VDD2.n2 VDD2.n1 9.3005
R2839 VDD2.n57 VDD2.n56 9.3005
R2840 VDD2.n55 VDD2.n54 9.3005
R2841 VDD2.n6 VDD2.n5 9.3005
R2842 VDD2.n49 VDD2.n48 9.3005
R2843 VDD2.n47 VDD2.n46 9.3005
R2844 VDD2.n23 VDD2.n22 9.3005
R2845 VDD2.n18 VDD2.n17 9.3005
R2846 VDD2.n29 VDD2.n28 9.3005
R2847 VDD2.n31 VDD2.n30 9.3005
R2848 VDD2.n14 VDD2.n13 9.3005
R2849 VDD2.n37 VDD2.n36 9.3005
R2850 VDD2.n39 VDD2.n38 9.3005
R2851 VDD2.n40 VDD2.n9 9.3005
R2852 VDD2.n130 VDD2.n71 8.92171
R2853 VDD2.n98 VDD2.n97 8.92171
R2854 VDD2.n28 VDD2.n27 8.92171
R2855 VDD2.n61 VDD2.n2 8.92171
R2856 VDD2.n131 VDD2.n69 8.14595
R2857 VDD2.n94 VDD2.n88 8.14595
R2858 VDD2.n24 VDD2.n18 8.14595
R2859 VDD2.n62 VDD2.n0 8.14595
R2860 VDD2.n93 VDD2.n90 7.3702
R2861 VDD2.n23 VDD2.n20 7.3702
R2862 VDD2.n133 VDD2.n69 5.81868
R2863 VDD2.n94 VDD2.n93 5.81868
R2864 VDD2.n24 VDD2.n23 5.81868
R2865 VDD2.n64 VDD2.n0 5.81868
R2866 VDD2.n131 VDD2.n130 5.04292
R2867 VDD2.n97 VDD2.n88 5.04292
R2868 VDD2.n27 VDD2.n18 5.04292
R2869 VDD2.n62 VDD2.n61 5.04292
R2870 VDD2.n127 VDD2.n71 4.26717
R2871 VDD2.n98 VDD2.n86 4.26717
R2872 VDD2.n28 VDD2.n16 4.26717
R2873 VDD2.n58 VDD2.n2 4.26717
R2874 VDD2.n126 VDD2.n73 3.49141
R2875 VDD2.n102 VDD2.n101 3.49141
R2876 VDD2.n32 VDD2.n31 3.49141
R2877 VDD2.n57 VDD2.n4 3.49141
R2878 VDD2.n92 VDD2.n91 2.84303
R2879 VDD2.n22 VDD2.n21 2.84303
R2880 VDD2.n123 VDD2.n122 2.71565
R2881 VDD2.n105 VDD2.n84 2.71565
R2882 VDD2.n35 VDD2.n14 2.71565
R2883 VDD2.n54 VDD2.n53 2.71565
R2884 VDD2.n136 VDD2.n134 2.35395
R2885 VDD2.n119 VDD2.n75 1.93989
R2886 VDD2.n106 VDD2.n82 1.93989
R2887 VDD2.n36 VDD2.n12 1.93989
R2888 VDD2.n50 VDD2.n6 1.93989
R2889 VDD2.n137 VDD2.t6 1.62079
R2890 VDD2.n137 VDD2.t2 1.62079
R2891 VDD2.n135 VDD2.t3 1.62079
R2892 VDD2.n135 VDD2.t9 1.62079
R2893 VDD2.n67 VDD2.t1 1.62079
R2894 VDD2.n67 VDD2.t4 1.62079
R2895 VDD2.n65 VDD2.t7 1.62079
R2896 VDD2.n65 VDD2.t0 1.62079
R2897 VDD2.n118 VDD2.n77 1.16414
R2898 VDD2.n110 VDD2.n109 1.16414
R2899 VDD2.n41 VDD2.n39 1.16414
R2900 VDD2.n49 VDD2.n8 1.16414
R2901 VDD2 VDD2.n136 0.647052
R2902 VDD2.n68 VDD2.n66 0.533516
R2903 VDD2.n115 VDD2.n114 0.388379
R2904 VDD2.n81 VDD2.n79 0.388379
R2905 VDD2.n40 VDD2.n10 0.388379
R2906 VDD2.n46 VDD2.n45 0.388379
R2907 VDD2.n132 VDD2.n70 0.155672
R2908 VDD2.n125 VDD2.n70 0.155672
R2909 VDD2.n125 VDD2.n124 0.155672
R2910 VDD2.n124 VDD2.n74 0.155672
R2911 VDD2.n117 VDD2.n74 0.155672
R2912 VDD2.n117 VDD2.n116 0.155672
R2913 VDD2.n116 VDD2.n78 0.155672
R2914 VDD2.n108 VDD2.n78 0.155672
R2915 VDD2.n108 VDD2.n107 0.155672
R2916 VDD2.n107 VDD2.n83 0.155672
R2917 VDD2.n100 VDD2.n83 0.155672
R2918 VDD2.n100 VDD2.n99 0.155672
R2919 VDD2.n99 VDD2.n87 0.155672
R2920 VDD2.n92 VDD2.n87 0.155672
R2921 VDD2.n22 VDD2.n17 0.155672
R2922 VDD2.n29 VDD2.n17 0.155672
R2923 VDD2.n30 VDD2.n29 0.155672
R2924 VDD2.n30 VDD2.n13 0.155672
R2925 VDD2.n37 VDD2.n13 0.155672
R2926 VDD2.n38 VDD2.n37 0.155672
R2927 VDD2.n38 VDD2.n9 0.155672
R2928 VDD2.n47 VDD2.n9 0.155672
R2929 VDD2.n48 VDD2.n47 0.155672
R2930 VDD2.n48 VDD2.n5 0.155672
R2931 VDD2.n55 VDD2.n5 0.155672
R2932 VDD2.n56 VDD2.n55 0.155672
R2933 VDD2.n56 VDD2.n1 0.155672
R2934 VDD2.n63 VDD2.n1 0.155672
C0 VP VDD1 11.074201f
C1 VP VDD2 0.55779f
C2 VN VTAIL 11.2205f
C3 VN VDD1 0.152602f
C4 VN VDD2 10.6729f
C5 VTAIL VDD1 10.4751f
C6 VN VP 8.15274f
C7 VTAIL VDD2 10.524401f
C8 VDD1 VDD2 2.04452f
C9 VTAIL VP 11.2348f
C10 VDD2 B 7.031544f
C11 VDD1 B 6.99155f
C12 VTAIL B 8.140217f
C13 VN B 17.224209f
C14 VP B 15.729388f
C15 VDD2.n0 B 0.035557f
C16 VDD2.n1 B 0.024138f
C17 VDD2.n2 B 0.012971f
C18 VDD2.n3 B 0.030658f
C19 VDD2.n4 B 0.013734f
C20 VDD2.n5 B 0.024138f
C21 VDD2.n6 B 0.012971f
C22 VDD2.n7 B 0.030658f
C23 VDD2.n8 B 0.013734f
C24 VDD2.n9 B 0.024138f
C25 VDD2.n10 B 0.013352f
C26 VDD2.n11 B 0.030658f
C27 VDD2.n12 B 0.013734f
C28 VDD2.n13 B 0.024138f
C29 VDD2.n14 B 0.012971f
C30 VDD2.n15 B 0.030658f
C31 VDD2.n16 B 0.013734f
C32 VDD2.n17 B 0.024138f
C33 VDD2.n18 B 0.012971f
C34 VDD2.n19 B 0.022993f
C35 VDD2.n20 B 0.021673f
C36 VDD2.t5 B 0.051808f
C37 VDD2.n21 B 0.176071f
C38 VDD2.n22 B 1.24134f
C39 VDD2.n23 B 0.012971f
C40 VDD2.n24 B 0.013734f
C41 VDD2.n25 B 0.030658f
C42 VDD2.n26 B 0.030658f
C43 VDD2.n27 B 0.013734f
C44 VDD2.n28 B 0.012971f
C45 VDD2.n29 B 0.024138f
C46 VDD2.n30 B 0.024138f
C47 VDD2.n31 B 0.012971f
C48 VDD2.n32 B 0.013734f
C49 VDD2.n33 B 0.030658f
C50 VDD2.n34 B 0.030658f
C51 VDD2.n35 B 0.013734f
C52 VDD2.n36 B 0.012971f
C53 VDD2.n37 B 0.024138f
C54 VDD2.n38 B 0.024138f
C55 VDD2.n39 B 0.012971f
C56 VDD2.n40 B 0.012971f
C57 VDD2.n41 B 0.013734f
C58 VDD2.n42 B 0.030658f
C59 VDD2.n43 B 0.030658f
C60 VDD2.n44 B 0.030658f
C61 VDD2.n45 B 0.013352f
C62 VDD2.n46 B 0.012971f
C63 VDD2.n47 B 0.024138f
C64 VDD2.n48 B 0.024138f
C65 VDD2.n49 B 0.012971f
C66 VDD2.n50 B 0.013734f
C67 VDD2.n51 B 0.030658f
C68 VDD2.n52 B 0.030658f
C69 VDD2.n53 B 0.013734f
C70 VDD2.n54 B 0.012971f
C71 VDD2.n55 B 0.024138f
C72 VDD2.n56 B 0.024138f
C73 VDD2.n57 B 0.012971f
C74 VDD2.n58 B 0.013734f
C75 VDD2.n59 B 0.030658f
C76 VDD2.n60 B 0.069249f
C77 VDD2.n61 B 0.013734f
C78 VDD2.n62 B 0.012971f
C79 VDD2.n63 B 0.059091f
C80 VDD2.n64 B 0.06603f
C81 VDD2.t7 B 0.233091f
C82 VDD2.t0 B 0.233091f
C83 VDD2.n65 B 2.08096f
C84 VDD2.n66 B 0.645078f
C85 VDD2.t1 B 0.233091f
C86 VDD2.t4 B 0.233091f
C87 VDD2.n67 B 2.09464f
C88 VDD2.n68 B 2.71734f
C89 VDD2.n69 B 0.035557f
C90 VDD2.n70 B 0.024138f
C91 VDD2.n71 B 0.012971f
C92 VDD2.n72 B 0.030658f
C93 VDD2.n73 B 0.013734f
C94 VDD2.n74 B 0.024138f
C95 VDD2.n75 B 0.012971f
C96 VDD2.n76 B 0.030658f
C97 VDD2.n77 B 0.013734f
C98 VDD2.n78 B 0.024138f
C99 VDD2.n79 B 0.013352f
C100 VDD2.n80 B 0.030658f
C101 VDD2.n81 B 0.012971f
C102 VDD2.n82 B 0.013734f
C103 VDD2.n83 B 0.024138f
C104 VDD2.n84 B 0.012971f
C105 VDD2.n85 B 0.030658f
C106 VDD2.n86 B 0.013734f
C107 VDD2.n87 B 0.024138f
C108 VDD2.n88 B 0.012971f
C109 VDD2.n89 B 0.022993f
C110 VDD2.n90 B 0.021673f
C111 VDD2.t8 B 0.051808f
C112 VDD2.n91 B 0.176071f
C113 VDD2.n92 B 1.24134f
C114 VDD2.n93 B 0.012971f
C115 VDD2.n94 B 0.013734f
C116 VDD2.n95 B 0.030658f
C117 VDD2.n96 B 0.030658f
C118 VDD2.n97 B 0.013734f
C119 VDD2.n98 B 0.012971f
C120 VDD2.n99 B 0.024138f
C121 VDD2.n100 B 0.024138f
C122 VDD2.n101 B 0.012971f
C123 VDD2.n102 B 0.013734f
C124 VDD2.n103 B 0.030658f
C125 VDD2.n104 B 0.030658f
C126 VDD2.n105 B 0.013734f
C127 VDD2.n106 B 0.012971f
C128 VDD2.n107 B 0.024138f
C129 VDD2.n108 B 0.024138f
C130 VDD2.n109 B 0.012971f
C131 VDD2.n110 B 0.013734f
C132 VDD2.n111 B 0.030658f
C133 VDD2.n112 B 0.030658f
C134 VDD2.n113 B 0.030658f
C135 VDD2.n114 B 0.013352f
C136 VDD2.n115 B 0.012971f
C137 VDD2.n116 B 0.024138f
C138 VDD2.n117 B 0.024138f
C139 VDD2.n118 B 0.012971f
C140 VDD2.n119 B 0.013734f
C141 VDD2.n120 B 0.030658f
C142 VDD2.n121 B 0.030658f
C143 VDD2.n122 B 0.013734f
C144 VDD2.n123 B 0.012971f
C145 VDD2.n124 B 0.024138f
C146 VDD2.n125 B 0.024138f
C147 VDD2.n126 B 0.012971f
C148 VDD2.n127 B 0.013734f
C149 VDD2.n128 B 0.030658f
C150 VDD2.n129 B 0.069249f
C151 VDD2.n130 B 0.013734f
C152 VDD2.n131 B 0.012971f
C153 VDD2.n132 B 0.059091f
C154 VDD2.n133 B 0.055785f
C155 VDD2.n134 B 2.73371f
C156 VDD2.t3 B 0.233091f
C157 VDD2.t9 B 0.233091f
C158 VDD2.n135 B 2.08097f
C159 VDD2.n136 B 0.431683f
C160 VDD2.t6 B 0.233091f
C161 VDD2.t2 B 0.233091f
C162 VDD2.n137 B 2.09461f
C163 VN.n0 B 0.029742f
C164 VN.t5 B 1.80344f
C165 VN.n1 B 0.026403f
C166 VN.n2 B 0.022558f
C167 VN.t8 B 1.80344f
C168 VN.n3 B 0.638867f
C169 VN.n4 B 0.022558f
C170 VN.n5 B 0.045034f
C171 VN.n6 B 0.022558f
C172 VN.t9 B 1.80344f
C173 VN.n7 B 0.022435f
C174 VN.n8 B 0.213555f
C175 VN.t2 B 1.80344f
C176 VN.t4 B 1.96959f
C177 VN.n9 B 0.68514f
C178 VN.n10 B 0.71248f
C179 VN.n11 B 0.041418f
C180 VN.n12 B 0.04093f
C181 VN.n13 B 0.022558f
C182 VN.n14 B 0.022558f
C183 VN.n15 B 0.022558f
C184 VN.n16 B 0.045034f
C185 VN.n17 B 0.031821f
C186 VN.n18 B 0.638867f
C187 VN.n19 B 0.031821f
C188 VN.n20 B 0.022558f
C189 VN.n21 B 0.022558f
C190 VN.n22 B 0.022558f
C191 VN.n23 B 0.022435f
C192 VN.n24 B 0.04093f
C193 VN.n25 B 0.041418f
C194 VN.n26 B 0.022558f
C195 VN.n27 B 0.022558f
C196 VN.n28 B 0.022225f
C197 VN.n29 B 0.042252f
C198 VN.n30 B 0.038973f
C199 VN.n31 B 0.022558f
C200 VN.n32 B 0.022558f
C201 VN.n33 B 0.022558f
C202 VN.n34 B 0.043022f
C203 VN.n35 B 0.030152f
C204 VN.n36 B 0.709163f
C205 VN.n37 B 0.035163f
C206 VN.n38 B 0.029742f
C207 VN.t1 B 1.80344f
C208 VN.n39 B 0.026403f
C209 VN.n40 B 0.022558f
C210 VN.t6 B 1.80344f
C211 VN.n41 B 0.638867f
C212 VN.n42 B 0.022558f
C213 VN.n43 B 0.045034f
C214 VN.n44 B 0.022558f
C215 VN.t0 B 1.80344f
C216 VN.n45 B 0.022435f
C217 VN.n46 B 0.213555f
C218 VN.t3 B 1.80344f
C219 VN.t7 B 1.96959f
C220 VN.n47 B 0.68514f
C221 VN.n48 B 0.71248f
C222 VN.n49 B 0.041418f
C223 VN.n50 B 0.04093f
C224 VN.n51 B 0.022558f
C225 VN.n52 B 0.022558f
C226 VN.n53 B 0.022558f
C227 VN.n54 B 0.045034f
C228 VN.n55 B 0.031821f
C229 VN.n56 B 0.638867f
C230 VN.n57 B 0.031821f
C231 VN.n58 B 0.022558f
C232 VN.n59 B 0.022558f
C233 VN.n60 B 0.022558f
C234 VN.n61 B 0.022435f
C235 VN.n62 B 0.04093f
C236 VN.n63 B 0.041418f
C237 VN.n64 B 0.022558f
C238 VN.n65 B 0.022558f
C239 VN.n66 B 0.022225f
C240 VN.n67 B 0.042252f
C241 VN.n68 B 0.038973f
C242 VN.n69 B 0.022558f
C243 VN.n70 B 0.022558f
C244 VN.n71 B 0.022558f
C245 VN.n72 B 0.043022f
C246 VN.n73 B 0.030152f
C247 VN.n74 B 0.709163f
C248 VN.n75 B 1.34515f
C249 VTAIL.t6 B 0.238822f
C250 VTAIL.t7 B 0.238822f
C251 VTAIL.n0 B 2.06188f
C252 VTAIL.n1 B 0.516371f
C253 VTAIL.n2 B 0.036431f
C254 VTAIL.n3 B 0.024731f
C255 VTAIL.n4 B 0.01329f
C256 VTAIL.n5 B 0.031412f
C257 VTAIL.n6 B 0.014071f
C258 VTAIL.n7 B 0.024731f
C259 VTAIL.n8 B 0.01329f
C260 VTAIL.n9 B 0.031412f
C261 VTAIL.n10 B 0.014071f
C262 VTAIL.n11 B 0.024731f
C263 VTAIL.n12 B 0.01368f
C264 VTAIL.n13 B 0.031412f
C265 VTAIL.n14 B 0.014071f
C266 VTAIL.n15 B 0.024731f
C267 VTAIL.n16 B 0.01329f
C268 VTAIL.n17 B 0.031412f
C269 VTAIL.n18 B 0.014071f
C270 VTAIL.n19 B 0.024731f
C271 VTAIL.n20 B 0.01329f
C272 VTAIL.n21 B 0.023559f
C273 VTAIL.n22 B 0.022206f
C274 VTAIL.t18 B 0.053082f
C275 VTAIL.n23 B 0.1804f
C276 VTAIL.n24 B 1.27186f
C277 VTAIL.n25 B 0.01329f
C278 VTAIL.n26 B 0.014071f
C279 VTAIL.n27 B 0.031412f
C280 VTAIL.n28 B 0.031412f
C281 VTAIL.n29 B 0.014071f
C282 VTAIL.n30 B 0.01329f
C283 VTAIL.n31 B 0.024731f
C284 VTAIL.n32 B 0.024731f
C285 VTAIL.n33 B 0.01329f
C286 VTAIL.n34 B 0.014071f
C287 VTAIL.n35 B 0.031412f
C288 VTAIL.n36 B 0.031412f
C289 VTAIL.n37 B 0.014071f
C290 VTAIL.n38 B 0.01329f
C291 VTAIL.n39 B 0.024731f
C292 VTAIL.n40 B 0.024731f
C293 VTAIL.n41 B 0.01329f
C294 VTAIL.n42 B 0.01329f
C295 VTAIL.n43 B 0.014071f
C296 VTAIL.n44 B 0.031412f
C297 VTAIL.n45 B 0.031412f
C298 VTAIL.n46 B 0.031412f
C299 VTAIL.n47 B 0.01368f
C300 VTAIL.n48 B 0.01329f
C301 VTAIL.n49 B 0.024731f
C302 VTAIL.n50 B 0.024731f
C303 VTAIL.n51 B 0.01329f
C304 VTAIL.n52 B 0.014071f
C305 VTAIL.n53 B 0.031412f
C306 VTAIL.n54 B 0.031412f
C307 VTAIL.n55 B 0.014071f
C308 VTAIL.n56 B 0.01329f
C309 VTAIL.n57 B 0.024731f
C310 VTAIL.n58 B 0.024731f
C311 VTAIL.n59 B 0.01329f
C312 VTAIL.n60 B 0.014071f
C313 VTAIL.n61 B 0.031412f
C314 VTAIL.n62 B 0.070952f
C315 VTAIL.n63 B 0.014071f
C316 VTAIL.n64 B 0.01329f
C317 VTAIL.n65 B 0.060544f
C318 VTAIL.n66 B 0.040105f
C319 VTAIL.n67 B 0.341793f
C320 VTAIL.t14 B 0.238822f
C321 VTAIL.t11 B 0.238822f
C322 VTAIL.n68 B 2.06188f
C323 VTAIL.n69 B 0.614953f
C324 VTAIL.t16 B 0.238822f
C325 VTAIL.t17 B 0.238822f
C326 VTAIL.n70 B 2.06188f
C327 VTAIL.n71 B 1.97794f
C328 VTAIL.t4 B 0.238822f
C329 VTAIL.t1 B 0.238822f
C330 VTAIL.n72 B 2.06189f
C331 VTAIL.n73 B 1.97793f
C332 VTAIL.t2 B 0.238822f
C333 VTAIL.t9 B 0.238822f
C334 VTAIL.n74 B 2.06189f
C335 VTAIL.n75 B 0.614942f
C336 VTAIL.n76 B 0.036431f
C337 VTAIL.n77 B 0.024731f
C338 VTAIL.n78 B 0.01329f
C339 VTAIL.n79 B 0.031412f
C340 VTAIL.n80 B 0.014071f
C341 VTAIL.n81 B 0.024731f
C342 VTAIL.n82 B 0.01329f
C343 VTAIL.n83 B 0.031412f
C344 VTAIL.n84 B 0.014071f
C345 VTAIL.n85 B 0.024731f
C346 VTAIL.n86 B 0.01368f
C347 VTAIL.n87 B 0.031412f
C348 VTAIL.n88 B 0.01329f
C349 VTAIL.n89 B 0.014071f
C350 VTAIL.n90 B 0.024731f
C351 VTAIL.n91 B 0.01329f
C352 VTAIL.n92 B 0.031412f
C353 VTAIL.n93 B 0.014071f
C354 VTAIL.n94 B 0.024731f
C355 VTAIL.n95 B 0.01329f
C356 VTAIL.n96 B 0.023559f
C357 VTAIL.n97 B 0.022206f
C358 VTAIL.t3 B 0.053082f
C359 VTAIL.n98 B 0.1804f
C360 VTAIL.n99 B 1.27186f
C361 VTAIL.n100 B 0.01329f
C362 VTAIL.n101 B 0.014071f
C363 VTAIL.n102 B 0.031412f
C364 VTAIL.n103 B 0.031412f
C365 VTAIL.n104 B 0.014071f
C366 VTAIL.n105 B 0.01329f
C367 VTAIL.n106 B 0.024731f
C368 VTAIL.n107 B 0.024731f
C369 VTAIL.n108 B 0.01329f
C370 VTAIL.n109 B 0.014071f
C371 VTAIL.n110 B 0.031412f
C372 VTAIL.n111 B 0.031412f
C373 VTAIL.n112 B 0.014071f
C374 VTAIL.n113 B 0.01329f
C375 VTAIL.n114 B 0.024731f
C376 VTAIL.n115 B 0.024731f
C377 VTAIL.n116 B 0.01329f
C378 VTAIL.n117 B 0.014071f
C379 VTAIL.n118 B 0.031412f
C380 VTAIL.n119 B 0.031412f
C381 VTAIL.n120 B 0.031412f
C382 VTAIL.n121 B 0.01368f
C383 VTAIL.n122 B 0.01329f
C384 VTAIL.n123 B 0.024731f
C385 VTAIL.n124 B 0.024731f
C386 VTAIL.n125 B 0.01329f
C387 VTAIL.n126 B 0.014071f
C388 VTAIL.n127 B 0.031412f
C389 VTAIL.n128 B 0.031412f
C390 VTAIL.n129 B 0.014071f
C391 VTAIL.n130 B 0.01329f
C392 VTAIL.n131 B 0.024731f
C393 VTAIL.n132 B 0.024731f
C394 VTAIL.n133 B 0.01329f
C395 VTAIL.n134 B 0.014071f
C396 VTAIL.n135 B 0.031412f
C397 VTAIL.n136 B 0.070952f
C398 VTAIL.n137 B 0.014071f
C399 VTAIL.n138 B 0.01329f
C400 VTAIL.n139 B 0.060544f
C401 VTAIL.n140 B 0.040105f
C402 VTAIL.n141 B 0.341793f
C403 VTAIL.t13 B 0.238822f
C404 VTAIL.t19 B 0.238822f
C405 VTAIL.n142 B 2.06189f
C406 VTAIL.n143 B 0.558609f
C407 VTAIL.t12 B 0.238822f
C408 VTAIL.t15 B 0.238822f
C409 VTAIL.n144 B 2.06189f
C410 VTAIL.n145 B 0.614942f
C411 VTAIL.n146 B 0.036431f
C412 VTAIL.n147 B 0.024731f
C413 VTAIL.n148 B 0.01329f
C414 VTAIL.n149 B 0.031412f
C415 VTAIL.n150 B 0.014071f
C416 VTAIL.n151 B 0.024731f
C417 VTAIL.n152 B 0.01329f
C418 VTAIL.n153 B 0.031412f
C419 VTAIL.n154 B 0.014071f
C420 VTAIL.n155 B 0.024731f
C421 VTAIL.n156 B 0.01368f
C422 VTAIL.n157 B 0.031412f
C423 VTAIL.n158 B 0.01329f
C424 VTAIL.n159 B 0.014071f
C425 VTAIL.n160 B 0.024731f
C426 VTAIL.n161 B 0.01329f
C427 VTAIL.n162 B 0.031412f
C428 VTAIL.n163 B 0.014071f
C429 VTAIL.n164 B 0.024731f
C430 VTAIL.n165 B 0.01329f
C431 VTAIL.n166 B 0.023559f
C432 VTAIL.n167 B 0.022206f
C433 VTAIL.t10 B 0.053082f
C434 VTAIL.n168 B 0.1804f
C435 VTAIL.n169 B 1.27186f
C436 VTAIL.n170 B 0.01329f
C437 VTAIL.n171 B 0.014071f
C438 VTAIL.n172 B 0.031412f
C439 VTAIL.n173 B 0.031412f
C440 VTAIL.n174 B 0.014071f
C441 VTAIL.n175 B 0.01329f
C442 VTAIL.n176 B 0.024731f
C443 VTAIL.n177 B 0.024731f
C444 VTAIL.n178 B 0.01329f
C445 VTAIL.n179 B 0.014071f
C446 VTAIL.n180 B 0.031412f
C447 VTAIL.n181 B 0.031412f
C448 VTAIL.n182 B 0.014071f
C449 VTAIL.n183 B 0.01329f
C450 VTAIL.n184 B 0.024731f
C451 VTAIL.n185 B 0.024731f
C452 VTAIL.n186 B 0.01329f
C453 VTAIL.n187 B 0.014071f
C454 VTAIL.n188 B 0.031412f
C455 VTAIL.n189 B 0.031412f
C456 VTAIL.n190 B 0.031412f
C457 VTAIL.n191 B 0.01368f
C458 VTAIL.n192 B 0.01329f
C459 VTAIL.n193 B 0.024731f
C460 VTAIL.n194 B 0.024731f
C461 VTAIL.n195 B 0.01329f
C462 VTAIL.n196 B 0.014071f
C463 VTAIL.n197 B 0.031412f
C464 VTAIL.n198 B 0.031412f
C465 VTAIL.n199 B 0.014071f
C466 VTAIL.n200 B 0.01329f
C467 VTAIL.n201 B 0.024731f
C468 VTAIL.n202 B 0.024731f
C469 VTAIL.n203 B 0.01329f
C470 VTAIL.n204 B 0.014071f
C471 VTAIL.n205 B 0.031412f
C472 VTAIL.n206 B 0.070952f
C473 VTAIL.n207 B 0.014071f
C474 VTAIL.n208 B 0.01329f
C475 VTAIL.n209 B 0.060544f
C476 VTAIL.n210 B 0.040105f
C477 VTAIL.n211 B 1.57357f
C478 VTAIL.n212 B 0.036431f
C479 VTAIL.n213 B 0.024731f
C480 VTAIL.n214 B 0.01329f
C481 VTAIL.n215 B 0.031412f
C482 VTAIL.n216 B 0.014071f
C483 VTAIL.n217 B 0.024731f
C484 VTAIL.n218 B 0.01329f
C485 VTAIL.n219 B 0.031412f
C486 VTAIL.n220 B 0.014071f
C487 VTAIL.n221 B 0.024731f
C488 VTAIL.n222 B 0.01368f
C489 VTAIL.n223 B 0.031412f
C490 VTAIL.n224 B 0.014071f
C491 VTAIL.n225 B 0.024731f
C492 VTAIL.n226 B 0.01329f
C493 VTAIL.n227 B 0.031412f
C494 VTAIL.n228 B 0.014071f
C495 VTAIL.n229 B 0.024731f
C496 VTAIL.n230 B 0.01329f
C497 VTAIL.n231 B 0.023559f
C498 VTAIL.n232 B 0.022206f
C499 VTAIL.t5 B 0.053082f
C500 VTAIL.n233 B 0.1804f
C501 VTAIL.n234 B 1.27186f
C502 VTAIL.n235 B 0.01329f
C503 VTAIL.n236 B 0.014071f
C504 VTAIL.n237 B 0.031412f
C505 VTAIL.n238 B 0.031412f
C506 VTAIL.n239 B 0.014071f
C507 VTAIL.n240 B 0.01329f
C508 VTAIL.n241 B 0.024731f
C509 VTAIL.n242 B 0.024731f
C510 VTAIL.n243 B 0.01329f
C511 VTAIL.n244 B 0.014071f
C512 VTAIL.n245 B 0.031412f
C513 VTAIL.n246 B 0.031412f
C514 VTAIL.n247 B 0.014071f
C515 VTAIL.n248 B 0.01329f
C516 VTAIL.n249 B 0.024731f
C517 VTAIL.n250 B 0.024731f
C518 VTAIL.n251 B 0.01329f
C519 VTAIL.n252 B 0.01329f
C520 VTAIL.n253 B 0.014071f
C521 VTAIL.n254 B 0.031412f
C522 VTAIL.n255 B 0.031412f
C523 VTAIL.n256 B 0.031412f
C524 VTAIL.n257 B 0.01368f
C525 VTAIL.n258 B 0.01329f
C526 VTAIL.n259 B 0.024731f
C527 VTAIL.n260 B 0.024731f
C528 VTAIL.n261 B 0.01329f
C529 VTAIL.n262 B 0.014071f
C530 VTAIL.n263 B 0.031412f
C531 VTAIL.n264 B 0.031412f
C532 VTAIL.n265 B 0.014071f
C533 VTAIL.n266 B 0.01329f
C534 VTAIL.n267 B 0.024731f
C535 VTAIL.n268 B 0.024731f
C536 VTAIL.n269 B 0.01329f
C537 VTAIL.n270 B 0.014071f
C538 VTAIL.n271 B 0.031412f
C539 VTAIL.n272 B 0.070952f
C540 VTAIL.n273 B 0.014071f
C541 VTAIL.n274 B 0.01329f
C542 VTAIL.n275 B 0.060544f
C543 VTAIL.n276 B 0.040105f
C544 VTAIL.n277 B 1.57357f
C545 VTAIL.t8 B 0.238822f
C546 VTAIL.t0 B 0.238822f
C547 VTAIL.n278 B 2.06188f
C548 VTAIL.n279 B 0.469656f
C549 VDD1.n0 B 0.036031f
C550 VDD1.n1 B 0.02446f
C551 VDD1.n2 B 0.013144f
C552 VDD1.n3 B 0.031067f
C553 VDD1.n4 B 0.013917f
C554 VDD1.n5 B 0.02446f
C555 VDD1.n6 B 0.013144f
C556 VDD1.n7 B 0.031067f
C557 VDD1.n8 B 0.013917f
C558 VDD1.n9 B 0.02446f
C559 VDD1.n10 B 0.01353f
C560 VDD1.n11 B 0.031067f
C561 VDD1.n12 B 0.013144f
C562 VDD1.n13 B 0.013917f
C563 VDD1.n14 B 0.02446f
C564 VDD1.n15 B 0.013144f
C565 VDD1.n16 B 0.031067f
C566 VDD1.n17 B 0.013917f
C567 VDD1.n18 B 0.02446f
C568 VDD1.n19 B 0.013144f
C569 VDD1.n20 B 0.0233f
C570 VDD1.n21 B 0.021962f
C571 VDD1.t9 B 0.0525f
C572 VDD1.n22 B 0.178421f
C573 VDD1.n23 B 1.25791f
C574 VDD1.n24 B 0.013144f
C575 VDD1.n25 B 0.013917f
C576 VDD1.n26 B 0.031067f
C577 VDD1.n27 B 0.031067f
C578 VDD1.n28 B 0.013917f
C579 VDD1.n29 B 0.013144f
C580 VDD1.n30 B 0.02446f
C581 VDD1.n31 B 0.02446f
C582 VDD1.n32 B 0.013144f
C583 VDD1.n33 B 0.013917f
C584 VDD1.n34 B 0.031067f
C585 VDD1.n35 B 0.031067f
C586 VDD1.n36 B 0.013917f
C587 VDD1.n37 B 0.013144f
C588 VDD1.n38 B 0.02446f
C589 VDD1.n39 B 0.02446f
C590 VDD1.n40 B 0.013144f
C591 VDD1.n41 B 0.013917f
C592 VDD1.n42 B 0.031067f
C593 VDD1.n43 B 0.031067f
C594 VDD1.n44 B 0.031067f
C595 VDD1.n45 B 0.01353f
C596 VDD1.n46 B 0.013144f
C597 VDD1.n47 B 0.02446f
C598 VDD1.n48 B 0.02446f
C599 VDD1.n49 B 0.013144f
C600 VDD1.n50 B 0.013917f
C601 VDD1.n51 B 0.031067f
C602 VDD1.n52 B 0.031067f
C603 VDD1.n53 B 0.013917f
C604 VDD1.n54 B 0.013144f
C605 VDD1.n55 B 0.02446f
C606 VDD1.n56 B 0.02446f
C607 VDD1.n57 B 0.013144f
C608 VDD1.n58 B 0.013917f
C609 VDD1.n59 B 0.031067f
C610 VDD1.n60 B 0.070174f
C611 VDD1.n61 B 0.013917f
C612 VDD1.n62 B 0.013144f
C613 VDD1.n63 B 0.05988f
C614 VDD1.n64 B 0.066912f
C615 VDD1.t1 B 0.236202f
C616 VDD1.t8 B 0.236202f
C617 VDD1.n65 B 2.10874f
C618 VDD1.n66 B 0.661565f
C619 VDD1.n67 B 0.036031f
C620 VDD1.n68 B 0.02446f
C621 VDD1.n69 B 0.013144f
C622 VDD1.n70 B 0.031067f
C623 VDD1.n71 B 0.013917f
C624 VDD1.n72 B 0.02446f
C625 VDD1.n73 B 0.013144f
C626 VDD1.n74 B 0.031067f
C627 VDD1.n75 B 0.013917f
C628 VDD1.n76 B 0.02446f
C629 VDD1.n77 B 0.01353f
C630 VDD1.n78 B 0.031067f
C631 VDD1.n79 B 0.013917f
C632 VDD1.n80 B 0.02446f
C633 VDD1.n81 B 0.013144f
C634 VDD1.n82 B 0.031067f
C635 VDD1.n83 B 0.013917f
C636 VDD1.n84 B 0.02446f
C637 VDD1.n85 B 0.013144f
C638 VDD1.n86 B 0.0233f
C639 VDD1.n87 B 0.021962f
C640 VDD1.t2 B 0.0525f
C641 VDD1.n88 B 0.178421f
C642 VDD1.n89 B 1.25791f
C643 VDD1.n90 B 0.013144f
C644 VDD1.n91 B 0.013917f
C645 VDD1.n92 B 0.031067f
C646 VDD1.n93 B 0.031067f
C647 VDD1.n94 B 0.013917f
C648 VDD1.n95 B 0.013144f
C649 VDD1.n96 B 0.02446f
C650 VDD1.n97 B 0.02446f
C651 VDD1.n98 B 0.013144f
C652 VDD1.n99 B 0.013917f
C653 VDD1.n100 B 0.031067f
C654 VDD1.n101 B 0.031067f
C655 VDD1.n102 B 0.013917f
C656 VDD1.n103 B 0.013144f
C657 VDD1.n104 B 0.02446f
C658 VDD1.n105 B 0.02446f
C659 VDD1.n106 B 0.013144f
C660 VDD1.n107 B 0.013144f
C661 VDD1.n108 B 0.013917f
C662 VDD1.n109 B 0.031067f
C663 VDD1.n110 B 0.031067f
C664 VDD1.n111 B 0.031067f
C665 VDD1.n112 B 0.01353f
C666 VDD1.n113 B 0.013144f
C667 VDD1.n114 B 0.02446f
C668 VDD1.n115 B 0.02446f
C669 VDD1.n116 B 0.013144f
C670 VDD1.n117 B 0.013917f
C671 VDD1.n118 B 0.031067f
C672 VDD1.n119 B 0.031067f
C673 VDD1.n120 B 0.013917f
C674 VDD1.n121 B 0.013144f
C675 VDD1.n122 B 0.02446f
C676 VDD1.n123 B 0.02446f
C677 VDD1.n124 B 0.013144f
C678 VDD1.n125 B 0.013917f
C679 VDD1.n126 B 0.031067f
C680 VDD1.n127 B 0.070174f
C681 VDD1.n128 B 0.013917f
C682 VDD1.n129 B 0.013144f
C683 VDD1.n130 B 0.05988f
C684 VDD1.n131 B 0.066912f
C685 VDD1.t3 B 0.236202f
C686 VDD1.t4 B 0.236202f
C687 VDD1.n132 B 2.10874f
C688 VDD1.n133 B 0.653688f
C689 VDD1.t7 B 0.236202f
C690 VDD1.t0 B 0.236202f
C691 VDD1.n134 B 2.1226f
C692 VDD1.n135 B 2.87089f
C693 VDD1.t5 B 0.236202f
C694 VDD1.t6 B 0.236202f
C695 VDD1.n136 B 2.10874f
C696 VDD1.n137 B 3.03963f
C697 VP.n0 B 0.030169f
C698 VP.t1 B 1.82934f
C699 VP.n1 B 0.026782f
C700 VP.n2 B 0.022881f
C701 VP.t8 B 1.82934f
C702 VP.n3 B 0.64804f
C703 VP.n4 B 0.022881f
C704 VP.n5 B 0.04568f
C705 VP.n6 B 0.022881f
C706 VP.t5 B 1.82934f
C707 VP.n7 B 0.022757f
C708 VP.n8 B 0.022881f
C709 VP.t2 B 1.82934f
C710 VP.n9 B 0.042859f
C711 VP.n10 B 0.022881f
C712 VP.n11 B 0.030585f
C713 VP.n12 B 0.030169f
C714 VP.t9 B 1.82934f
C715 VP.n13 B 0.026782f
C716 VP.n14 B 0.022881f
C717 VP.t4 B 1.82934f
C718 VP.n15 B 0.64804f
C719 VP.n16 B 0.022881f
C720 VP.n17 B 0.04568f
C721 VP.n18 B 0.022881f
C722 VP.t7 B 1.82934f
C723 VP.n19 B 0.022757f
C724 VP.n20 B 0.216622f
C725 VP.t0 B 1.82934f
C726 VP.t6 B 1.99787f
C727 VP.n21 B 0.694977f
C728 VP.n22 B 0.72271f
C729 VP.n23 B 0.042012f
C730 VP.n24 B 0.041517f
C731 VP.n25 B 0.022881f
C732 VP.n26 B 0.022881f
C733 VP.n27 B 0.022881f
C734 VP.n28 B 0.04568f
C735 VP.n29 B 0.032278f
C736 VP.n30 B 0.64804f
C737 VP.n31 B 0.032278f
C738 VP.n32 B 0.022881f
C739 VP.n33 B 0.022881f
C740 VP.n34 B 0.022881f
C741 VP.n35 B 0.022757f
C742 VP.n36 B 0.041517f
C743 VP.n37 B 0.042012f
C744 VP.n38 B 0.022881f
C745 VP.n39 B 0.022881f
C746 VP.n40 B 0.022544f
C747 VP.n41 B 0.042859f
C748 VP.n42 B 0.039533f
C749 VP.n43 B 0.022881f
C750 VP.n44 B 0.022881f
C751 VP.n45 B 0.022881f
C752 VP.n46 B 0.04364f
C753 VP.n47 B 0.030585f
C754 VP.n48 B 0.719345f
C755 VP.n49 B 1.35225f
C756 VP.t3 B 1.82934f
C757 VP.n50 B 0.719345f
C758 VP.n51 B 1.36797f
C759 VP.n52 B 0.030169f
C760 VP.n53 B 0.022881f
C761 VP.n54 B 0.04364f
C762 VP.n55 B 0.026782f
C763 VP.n56 B 0.039533f
C764 VP.n57 B 0.022881f
C765 VP.n58 B 0.022881f
C766 VP.n59 B 0.022881f
C767 VP.n60 B 0.022544f
C768 VP.n61 B 0.64804f
C769 VP.n62 B 0.042012f
C770 VP.n63 B 0.041517f
C771 VP.n64 B 0.022881f
C772 VP.n65 B 0.022881f
C773 VP.n66 B 0.022881f
C774 VP.n67 B 0.04568f
C775 VP.n68 B 0.032278f
C776 VP.n69 B 0.64804f
C777 VP.n70 B 0.032278f
C778 VP.n71 B 0.022881f
C779 VP.n72 B 0.022881f
C780 VP.n73 B 0.022881f
C781 VP.n74 B 0.022757f
C782 VP.n75 B 0.041517f
C783 VP.n76 B 0.042012f
C784 VP.n77 B 0.022881f
C785 VP.n78 B 0.022881f
C786 VP.n79 B 0.022544f
C787 VP.n80 B 0.042859f
C788 VP.n81 B 0.039533f
C789 VP.n82 B 0.022881f
C790 VP.n83 B 0.022881f
C791 VP.n84 B 0.022881f
C792 VP.n85 B 0.04364f
C793 VP.n86 B 0.030585f
C794 VP.n87 B 0.719345f
C795 VP.n88 B 0.035668f
.ends

