* NGSPICE file created from diff_pair_sample_0798.ext - technology: sky130A

.subckt diff_pair_sample_0798 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t3 w_n1554_n1418# sky130_fd_pr__pfet_01v8 ad=0.8775 pd=5.28 as=0.8775 ps=5.28 w=2.25 l=1.13
X1 VDD2.t1 VN.t0 VTAIL.t1 w_n1554_n1418# sky130_fd_pr__pfet_01v8 ad=0.8775 pd=5.28 as=0.8775 ps=5.28 w=2.25 l=1.13
X2 B.t11 B.t9 B.t10 w_n1554_n1418# sky130_fd_pr__pfet_01v8 ad=0.8775 pd=5.28 as=0 ps=0 w=2.25 l=1.13
X3 VDD2.t0 VN.t1 VTAIL.t0 w_n1554_n1418# sky130_fd_pr__pfet_01v8 ad=0.8775 pd=5.28 as=0.8775 ps=5.28 w=2.25 l=1.13
X4 B.t8 B.t6 B.t7 w_n1554_n1418# sky130_fd_pr__pfet_01v8 ad=0.8775 pd=5.28 as=0 ps=0 w=2.25 l=1.13
X5 B.t5 B.t3 B.t4 w_n1554_n1418# sky130_fd_pr__pfet_01v8 ad=0.8775 pd=5.28 as=0 ps=0 w=2.25 l=1.13
X6 VDD1.t0 VP.t1 VTAIL.t2 w_n1554_n1418# sky130_fd_pr__pfet_01v8 ad=0.8775 pd=5.28 as=0.8775 ps=5.28 w=2.25 l=1.13
X7 B.t2 B.t0 B.t1 w_n1554_n1418# sky130_fd_pr__pfet_01v8 ad=0.8775 pd=5.28 as=0 ps=0 w=2.25 l=1.13
R0 VP.n0 VP.t0 196.94
R1 VP.n0 VP.t1 163.567
R2 VP VP.n0 0.146778
R3 VTAIL.n3 VTAIL.t0 172.679
R4 VTAIL.n0 VTAIL.t2 172.679
R5 VTAIL.n2 VTAIL.t3 172.679
R6 VTAIL.n1 VTAIL.t1 172.679
R7 VTAIL.n1 VTAIL.n0 16.8238
R8 VTAIL.n3 VTAIL.n2 15.5652
R9 VTAIL.n2 VTAIL.n1 1.09964
R10 VTAIL VTAIL.n0 0.843172
R11 VTAIL VTAIL.n3 0.256966
R12 VDD1 VDD1.t0 218.315
R13 VDD1 VDD1.t1 189.732
R14 VN VN.t0 197.226
R15 VN VN.t1 163.714
R16 VDD2.n0 VDD2.t0 217.476
R17 VDD2.n0 VDD2.t1 189.358
R18 VDD2 VDD2.n0 0.373345
R19 B.n155 B.n154 585
R20 B.n153 B.n50 585
R21 B.n152 B.n151 585
R22 B.n150 B.n51 585
R23 B.n149 B.n148 585
R24 B.n147 B.n52 585
R25 B.n146 B.n145 585
R26 B.n144 B.n53 585
R27 B.n143 B.n142 585
R28 B.n141 B.n54 585
R29 B.n140 B.n139 585
R30 B.n138 B.n55 585
R31 B.n137 B.n136 585
R32 B.n134 B.n56 585
R33 B.n133 B.n132 585
R34 B.n131 B.n59 585
R35 B.n130 B.n129 585
R36 B.n128 B.n60 585
R37 B.n127 B.n126 585
R38 B.n125 B.n61 585
R39 B.n124 B.n123 585
R40 B.n122 B.n62 585
R41 B.n120 B.n119 585
R42 B.n118 B.n65 585
R43 B.n117 B.n116 585
R44 B.n115 B.n66 585
R45 B.n114 B.n113 585
R46 B.n112 B.n67 585
R47 B.n111 B.n110 585
R48 B.n109 B.n68 585
R49 B.n108 B.n107 585
R50 B.n106 B.n69 585
R51 B.n105 B.n104 585
R52 B.n103 B.n70 585
R53 B.n102 B.n101 585
R54 B.n156 B.n49 585
R55 B.n158 B.n157 585
R56 B.n159 B.n48 585
R57 B.n161 B.n160 585
R58 B.n162 B.n47 585
R59 B.n164 B.n163 585
R60 B.n165 B.n46 585
R61 B.n167 B.n166 585
R62 B.n168 B.n45 585
R63 B.n170 B.n169 585
R64 B.n171 B.n44 585
R65 B.n173 B.n172 585
R66 B.n174 B.n43 585
R67 B.n176 B.n175 585
R68 B.n177 B.n42 585
R69 B.n179 B.n178 585
R70 B.n180 B.n41 585
R71 B.n182 B.n181 585
R72 B.n183 B.n40 585
R73 B.n185 B.n184 585
R74 B.n186 B.n39 585
R75 B.n188 B.n187 585
R76 B.n189 B.n38 585
R77 B.n191 B.n190 585
R78 B.n192 B.n37 585
R79 B.n194 B.n193 585
R80 B.n195 B.n36 585
R81 B.n197 B.n196 585
R82 B.n198 B.n35 585
R83 B.n200 B.n199 585
R84 B.n201 B.n34 585
R85 B.n203 B.n202 585
R86 B.n204 B.n33 585
R87 B.n206 B.n205 585
R88 B.n259 B.n10 585
R89 B.n258 B.n257 585
R90 B.n256 B.n11 585
R91 B.n255 B.n254 585
R92 B.n253 B.n12 585
R93 B.n252 B.n251 585
R94 B.n250 B.n13 585
R95 B.n249 B.n248 585
R96 B.n247 B.n14 585
R97 B.n246 B.n245 585
R98 B.n244 B.n15 585
R99 B.n243 B.n242 585
R100 B.n241 B.n16 585
R101 B.n240 B.n239 585
R102 B.n238 B.n17 585
R103 B.n237 B.n236 585
R104 B.n235 B.n21 585
R105 B.n234 B.n233 585
R106 B.n232 B.n22 585
R107 B.n231 B.n230 585
R108 B.n229 B.n23 585
R109 B.n228 B.n227 585
R110 B.n225 B.n24 585
R111 B.n224 B.n223 585
R112 B.n222 B.n27 585
R113 B.n221 B.n220 585
R114 B.n219 B.n28 585
R115 B.n218 B.n217 585
R116 B.n216 B.n29 585
R117 B.n215 B.n214 585
R118 B.n213 B.n30 585
R119 B.n212 B.n211 585
R120 B.n210 B.n31 585
R121 B.n209 B.n208 585
R122 B.n207 B.n32 585
R123 B.n261 B.n260 585
R124 B.n262 B.n9 585
R125 B.n264 B.n263 585
R126 B.n265 B.n8 585
R127 B.n267 B.n266 585
R128 B.n268 B.n7 585
R129 B.n270 B.n269 585
R130 B.n271 B.n6 585
R131 B.n273 B.n272 585
R132 B.n274 B.n5 585
R133 B.n276 B.n275 585
R134 B.n277 B.n4 585
R135 B.n279 B.n278 585
R136 B.n280 B.n3 585
R137 B.n282 B.n281 585
R138 B.n283 B.n0 585
R139 B.n2 B.n1 585
R140 B.n79 B.n78 585
R141 B.n81 B.n80 585
R142 B.n82 B.n77 585
R143 B.n84 B.n83 585
R144 B.n85 B.n76 585
R145 B.n87 B.n86 585
R146 B.n88 B.n75 585
R147 B.n90 B.n89 585
R148 B.n91 B.n74 585
R149 B.n93 B.n92 585
R150 B.n94 B.n73 585
R151 B.n96 B.n95 585
R152 B.n97 B.n72 585
R153 B.n99 B.n98 585
R154 B.n100 B.n71 585
R155 B.n101 B.n100 569.379
R156 B.n156 B.n155 569.379
R157 B.n205 B.n32 569.379
R158 B.n260 B.n259 569.379
R159 B.n285 B.n284 256.663
R160 B.n63 B.t6 251.722
R161 B.n57 B.t0 251.722
R162 B.n25 B.t9 251.722
R163 B.n18 B.t3 251.722
R164 B.n284 B.n283 235.042
R165 B.n284 B.n2 235.042
R166 B.n57 B.t1 201.804
R167 B.n25 B.t11 201.804
R168 B.n63 B.t7 201.804
R169 B.n18 B.t5 201.804
R170 B.n58 B.t2 173.489
R171 B.n26 B.t10 173.489
R172 B.n64 B.t8 173.489
R173 B.n19 B.t4 173.489
R174 B.n101 B.n70 163.367
R175 B.n105 B.n70 163.367
R176 B.n106 B.n105 163.367
R177 B.n107 B.n106 163.367
R178 B.n107 B.n68 163.367
R179 B.n111 B.n68 163.367
R180 B.n112 B.n111 163.367
R181 B.n113 B.n112 163.367
R182 B.n113 B.n66 163.367
R183 B.n117 B.n66 163.367
R184 B.n118 B.n117 163.367
R185 B.n119 B.n118 163.367
R186 B.n119 B.n62 163.367
R187 B.n124 B.n62 163.367
R188 B.n125 B.n124 163.367
R189 B.n126 B.n125 163.367
R190 B.n126 B.n60 163.367
R191 B.n130 B.n60 163.367
R192 B.n131 B.n130 163.367
R193 B.n132 B.n131 163.367
R194 B.n132 B.n56 163.367
R195 B.n137 B.n56 163.367
R196 B.n138 B.n137 163.367
R197 B.n139 B.n138 163.367
R198 B.n139 B.n54 163.367
R199 B.n143 B.n54 163.367
R200 B.n144 B.n143 163.367
R201 B.n145 B.n144 163.367
R202 B.n145 B.n52 163.367
R203 B.n149 B.n52 163.367
R204 B.n150 B.n149 163.367
R205 B.n151 B.n150 163.367
R206 B.n151 B.n50 163.367
R207 B.n155 B.n50 163.367
R208 B.n205 B.n204 163.367
R209 B.n204 B.n203 163.367
R210 B.n203 B.n34 163.367
R211 B.n199 B.n34 163.367
R212 B.n199 B.n198 163.367
R213 B.n198 B.n197 163.367
R214 B.n197 B.n36 163.367
R215 B.n193 B.n36 163.367
R216 B.n193 B.n192 163.367
R217 B.n192 B.n191 163.367
R218 B.n191 B.n38 163.367
R219 B.n187 B.n38 163.367
R220 B.n187 B.n186 163.367
R221 B.n186 B.n185 163.367
R222 B.n185 B.n40 163.367
R223 B.n181 B.n40 163.367
R224 B.n181 B.n180 163.367
R225 B.n180 B.n179 163.367
R226 B.n179 B.n42 163.367
R227 B.n175 B.n42 163.367
R228 B.n175 B.n174 163.367
R229 B.n174 B.n173 163.367
R230 B.n173 B.n44 163.367
R231 B.n169 B.n44 163.367
R232 B.n169 B.n168 163.367
R233 B.n168 B.n167 163.367
R234 B.n167 B.n46 163.367
R235 B.n163 B.n46 163.367
R236 B.n163 B.n162 163.367
R237 B.n162 B.n161 163.367
R238 B.n161 B.n48 163.367
R239 B.n157 B.n48 163.367
R240 B.n157 B.n156 163.367
R241 B.n259 B.n258 163.367
R242 B.n258 B.n11 163.367
R243 B.n254 B.n11 163.367
R244 B.n254 B.n253 163.367
R245 B.n253 B.n252 163.367
R246 B.n252 B.n13 163.367
R247 B.n248 B.n13 163.367
R248 B.n248 B.n247 163.367
R249 B.n247 B.n246 163.367
R250 B.n246 B.n15 163.367
R251 B.n242 B.n15 163.367
R252 B.n242 B.n241 163.367
R253 B.n241 B.n240 163.367
R254 B.n240 B.n17 163.367
R255 B.n236 B.n17 163.367
R256 B.n236 B.n235 163.367
R257 B.n235 B.n234 163.367
R258 B.n234 B.n22 163.367
R259 B.n230 B.n22 163.367
R260 B.n230 B.n229 163.367
R261 B.n229 B.n228 163.367
R262 B.n228 B.n24 163.367
R263 B.n223 B.n24 163.367
R264 B.n223 B.n222 163.367
R265 B.n222 B.n221 163.367
R266 B.n221 B.n28 163.367
R267 B.n217 B.n28 163.367
R268 B.n217 B.n216 163.367
R269 B.n216 B.n215 163.367
R270 B.n215 B.n30 163.367
R271 B.n211 B.n30 163.367
R272 B.n211 B.n210 163.367
R273 B.n210 B.n209 163.367
R274 B.n209 B.n32 163.367
R275 B.n260 B.n9 163.367
R276 B.n264 B.n9 163.367
R277 B.n265 B.n264 163.367
R278 B.n266 B.n265 163.367
R279 B.n266 B.n7 163.367
R280 B.n270 B.n7 163.367
R281 B.n271 B.n270 163.367
R282 B.n272 B.n271 163.367
R283 B.n272 B.n5 163.367
R284 B.n276 B.n5 163.367
R285 B.n277 B.n276 163.367
R286 B.n278 B.n277 163.367
R287 B.n278 B.n3 163.367
R288 B.n282 B.n3 163.367
R289 B.n283 B.n282 163.367
R290 B.n78 B.n2 163.367
R291 B.n81 B.n78 163.367
R292 B.n82 B.n81 163.367
R293 B.n83 B.n82 163.367
R294 B.n83 B.n76 163.367
R295 B.n87 B.n76 163.367
R296 B.n88 B.n87 163.367
R297 B.n89 B.n88 163.367
R298 B.n89 B.n74 163.367
R299 B.n93 B.n74 163.367
R300 B.n94 B.n93 163.367
R301 B.n95 B.n94 163.367
R302 B.n95 B.n72 163.367
R303 B.n99 B.n72 163.367
R304 B.n100 B.n99 163.367
R305 B.n121 B.n64 59.5399
R306 B.n135 B.n58 59.5399
R307 B.n226 B.n26 59.5399
R308 B.n20 B.n19 59.5399
R309 B.n261 B.n10 36.9956
R310 B.n207 B.n206 36.9956
R311 B.n154 B.n49 36.9956
R312 B.n102 B.n71 36.9956
R313 B.n64 B.n63 28.3157
R314 B.n58 B.n57 28.3157
R315 B.n26 B.n25 28.3157
R316 B.n19 B.n18 28.3157
R317 B B.n285 18.0485
R318 B.n262 B.n261 10.6151
R319 B.n263 B.n262 10.6151
R320 B.n263 B.n8 10.6151
R321 B.n267 B.n8 10.6151
R322 B.n268 B.n267 10.6151
R323 B.n269 B.n268 10.6151
R324 B.n269 B.n6 10.6151
R325 B.n273 B.n6 10.6151
R326 B.n274 B.n273 10.6151
R327 B.n275 B.n274 10.6151
R328 B.n275 B.n4 10.6151
R329 B.n279 B.n4 10.6151
R330 B.n280 B.n279 10.6151
R331 B.n281 B.n280 10.6151
R332 B.n281 B.n0 10.6151
R333 B.n257 B.n10 10.6151
R334 B.n257 B.n256 10.6151
R335 B.n256 B.n255 10.6151
R336 B.n255 B.n12 10.6151
R337 B.n251 B.n12 10.6151
R338 B.n251 B.n250 10.6151
R339 B.n250 B.n249 10.6151
R340 B.n249 B.n14 10.6151
R341 B.n245 B.n14 10.6151
R342 B.n245 B.n244 10.6151
R343 B.n244 B.n243 10.6151
R344 B.n243 B.n16 10.6151
R345 B.n239 B.n238 10.6151
R346 B.n238 B.n237 10.6151
R347 B.n237 B.n21 10.6151
R348 B.n233 B.n21 10.6151
R349 B.n233 B.n232 10.6151
R350 B.n232 B.n231 10.6151
R351 B.n231 B.n23 10.6151
R352 B.n227 B.n23 10.6151
R353 B.n225 B.n224 10.6151
R354 B.n224 B.n27 10.6151
R355 B.n220 B.n27 10.6151
R356 B.n220 B.n219 10.6151
R357 B.n219 B.n218 10.6151
R358 B.n218 B.n29 10.6151
R359 B.n214 B.n29 10.6151
R360 B.n214 B.n213 10.6151
R361 B.n213 B.n212 10.6151
R362 B.n212 B.n31 10.6151
R363 B.n208 B.n31 10.6151
R364 B.n208 B.n207 10.6151
R365 B.n206 B.n33 10.6151
R366 B.n202 B.n33 10.6151
R367 B.n202 B.n201 10.6151
R368 B.n201 B.n200 10.6151
R369 B.n200 B.n35 10.6151
R370 B.n196 B.n35 10.6151
R371 B.n196 B.n195 10.6151
R372 B.n195 B.n194 10.6151
R373 B.n194 B.n37 10.6151
R374 B.n190 B.n37 10.6151
R375 B.n190 B.n189 10.6151
R376 B.n189 B.n188 10.6151
R377 B.n188 B.n39 10.6151
R378 B.n184 B.n39 10.6151
R379 B.n184 B.n183 10.6151
R380 B.n183 B.n182 10.6151
R381 B.n182 B.n41 10.6151
R382 B.n178 B.n41 10.6151
R383 B.n178 B.n177 10.6151
R384 B.n177 B.n176 10.6151
R385 B.n176 B.n43 10.6151
R386 B.n172 B.n43 10.6151
R387 B.n172 B.n171 10.6151
R388 B.n171 B.n170 10.6151
R389 B.n170 B.n45 10.6151
R390 B.n166 B.n45 10.6151
R391 B.n166 B.n165 10.6151
R392 B.n165 B.n164 10.6151
R393 B.n164 B.n47 10.6151
R394 B.n160 B.n47 10.6151
R395 B.n160 B.n159 10.6151
R396 B.n159 B.n158 10.6151
R397 B.n158 B.n49 10.6151
R398 B.n79 B.n1 10.6151
R399 B.n80 B.n79 10.6151
R400 B.n80 B.n77 10.6151
R401 B.n84 B.n77 10.6151
R402 B.n85 B.n84 10.6151
R403 B.n86 B.n85 10.6151
R404 B.n86 B.n75 10.6151
R405 B.n90 B.n75 10.6151
R406 B.n91 B.n90 10.6151
R407 B.n92 B.n91 10.6151
R408 B.n92 B.n73 10.6151
R409 B.n96 B.n73 10.6151
R410 B.n97 B.n96 10.6151
R411 B.n98 B.n97 10.6151
R412 B.n98 B.n71 10.6151
R413 B.n103 B.n102 10.6151
R414 B.n104 B.n103 10.6151
R415 B.n104 B.n69 10.6151
R416 B.n108 B.n69 10.6151
R417 B.n109 B.n108 10.6151
R418 B.n110 B.n109 10.6151
R419 B.n110 B.n67 10.6151
R420 B.n114 B.n67 10.6151
R421 B.n115 B.n114 10.6151
R422 B.n116 B.n115 10.6151
R423 B.n116 B.n65 10.6151
R424 B.n120 B.n65 10.6151
R425 B.n123 B.n122 10.6151
R426 B.n123 B.n61 10.6151
R427 B.n127 B.n61 10.6151
R428 B.n128 B.n127 10.6151
R429 B.n129 B.n128 10.6151
R430 B.n129 B.n59 10.6151
R431 B.n133 B.n59 10.6151
R432 B.n134 B.n133 10.6151
R433 B.n136 B.n55 10.6151
R434 B.n140 B.n55 10.6151
R435 B.n141 B.n140 10.6151
R436 B.n142 B.n141 10.6151
R437 B.n142 B.n53 10.6151
R438 B.n146 B.n53 10.6151
R439 B.n147 B.n146 10.6151
R440 B.n148 B.n147 10.6151
R441 B.n148 B.n51 10.6151
R442 B.n152 B.n51 10.6151
R443 B.n153 B.n152 10.6151
R444 B.n154 B.n153 10.6151
R445 B.n285 B.n0 8.11757
R446 B.n285 B.n1 8.11757
R447 B.n239 B.n20 6.5566
R448 B.n227 B.n226 6.5566
R449 B.n122 B.n121 6.5566
R450 B.n135 B.n134 6.5566
R451 B.n20 B.n16 4.05904
R452 B.n226 B.n225 4.05904
R453 B.n121 B.n120 4.05904
R454 B.n136 B.n135 4.05904
C0 VDD1 VP 0.754784f
C1 w_n1554_n1418# VP 2.00341f
C2 w_n1554_n1418# VDD1 0.90649f
C3 VDD2 VP 0.276872f
C4 VDD2 VDD1 0.503661f
C5 VP VTAIL 0.721149f
C6 w_n1554_n1418# VDD2 0.914784f
C7 VDD1 VTAIL 2.09341f
C8 VP VN 2.97067f
C9 B VP 0.982725f
C10 VDD1 VN 0.153407f
C11 VDD1 B 0.758134f
C12 w_n1554_n1418# VTAIL 1.26849f
C13 w_n1554_n1418# VN 1.8124f
C14 w_n1554_n1418# B 4.47924f
C15 VDD2 VTAIL 2.13589f
C16 VDD2 VN 0.632877f
C17 VDD2 B 0.77593f
C18 VN VTAIL 0.70697f
C19 B VTAIL 1.03023f
C20 B VN 0.669051f
C21 VDD2 VSUBS 0.434421f
C22 VDD1 VSUBS 2.169918f
C23 VTAIL VSUBS 0.324224f
C24 VN VSUBS 3.45707f
C25 VP VSUBS 0.795627f
C26 B VSUBS 1.88854f
C27 w_n1554_n1418# VSUBS 28.0652f
C28 B.n0 VSUBS 0.007844f
C29 B.n1 VSUBS 0.007844f
C30 B.n2 VSUBS 0.0116f
C31 B.n3 VSUBS 0.00889f
C32 B.n4 VSUBS 0.00889f
C33 B.n5 VSUBS 0.00889f
C34 B.n6 VSUBS 0.00889f
C35 B.n7 VSUBS 0.00889f
C36 B.n8 VSUBS 0.00889f
C37 B.n9 VSUBS 0.00889f
C38 B.n10 VSUBS 0.023035f
C39 B.n11 VSUBS 0.00889f
C40 B.n12 VSUBS 0.00889f
C41 B.n13 VSUBS 0.00889f
C42 B.n14 VSUBS 0.00889f
C43 B.n15 VSUBS 0.00889f
C44 B.n16 VSUBS 0.006144f
C45 B.n17 VSUBS 0.00889f
C46 B.t4 VSUBS 0.063267f
C47 B.t5 VSUBS 0.071188f
C48 B.t3 VSUBS 0.154974f
C49 B.n18 VSUBS 0.078005f
C50 B.n19 VSUBS 0.069136f
C51 B.n20 VSUBS 0.020596f
C52 B.n21 VSUBS 0.00889f
C53 B.n22 VSUBS 0.00889f
C54 B.n23 VSUBS 0.00889f
C55 B.n24 VSUBS 0.00889f
C56 B.t10 VSUBS 0.063267f
C57 B.t11 VSUBS 0.071188f
C58 B.t9 VSUBS 0.154974f
C59 B.n25 VSUBS 0.078005f
C60 B.n26 VSUBS 0.069136f
C61 B.n27 VSUBS 0.00889f
C62 B.n28 VSUBS 0.00889f
C63 B.n29 VSUBS 0.00889f
C64 B.n30 VSUBS 0.00889f
C65 B.n31 VSUBS 0.00889f
C66 B.n32 VSUBS 0.023035f
C67 B.n33 VSUBS 0.00889f
C68 B.n34 VSUBS 0.00889f
C69 B.n35 VSUBS 0.00889f
C70 B.n36 VSUBS 0.00889f
C71 B.n37 VSUBS 0.00889f
C72 B.n38 VSUBS 0.00889f
C73 B.n39 VSUBS 0.00889f
C74 B.n40 VSUBS 0.00889f
C75 B.n41 VSUBS 0.00889f
C76 B.n42 VSUBS 0.00889f
C77 B.n43 VSUBS 0.00889f
C78 B.n44 VSUBS 0.00889f
C79 B.n45 VSUBS 0.00889f
C80 B.n46 VSUBS 0.00889f
C81 B.n47 VSUBS 0.00889f
C82 B.n48 VSUBS 0.00889f
C83 B.n49 VSUBS 0.023125f
C84 B.n50 VSUBS 0.00889f
C85 B.n51 VSUBS 0.00889f
C86 B.n52 VSUBS 0.00889f
C87 B.n53 VSUBS 0.00889f
C88 B.n54 VSUBS 0.00889f
C89 B.n55 VSUBS 0.00889f
C90 B.n56 VSUBS 0.00889f
C91 B.t2 VSUBS 0.063267f
C92 B.t1 VSUBS 0.071188f
C93 B.t0 VSUBS 0.154974f
C94 B.n57 VSUBS 0.078005f
C95 B.n58 VSUBS 0.069136f
C96 B.n59 VSUBS 0.00889f
C97 B.n60 VSUBS 0.00889f
C98 B.n61 VSUBS 0.00889f
C99 B.n62 VSUBS 0.00889f
C100 B.t8 VSUBS 0.063267f
C101 B.t7 VSUBS 0.071188f
C102 B.t6 VSUBS 0.154974f
C103 B.n63 VSUBS 0.078005f
C104 B.n64 VSUBS 0.069136f
C105 B.n65 VSUBS 0.00889f
C106 B.n66 VSUBS 0.00889f
C107 B.n67 VSUBS 0.00889f
C108 B.n68 VSUBS 0.00889f
C109 B.n69 VSUBS 0.00889f
C110 B.n70 VSUBS 0.00889f
C111 B.n71 VSUBS 0.022198f
C112 B.n72 VSUBS 0.00889f
C113 B.n73 VSUBS 0.00889f
C114 B.n74 VSUBS 0.00889f
C115 B.n75 VSUBS 0.00889f
C116 B.n76 VSUBS 0.00889f
C117 B.n77 VSUBS 0.00889f
C118 B.n78 VSUBS 0.00889f
C119 B.n79 VSUBS 0.00889f
C120 B.n80 VSUBS 0.00889f
C121 B.n81 VSUBS 0.00889f
C122 B.n82 VSUBS 0.00889f
C123 B.n83 VSUBS 0.00889f
C124 B.n84 VSUBS 0.00889f
C125 B.n85 VSUBS 0.00889f
C126 B.n86 VSUBS 0.00889f
C127 B.n87 VSUBS 0.00889f
C128 B.n88 VSUBS 0.00889f
C129 B.n89 VSUBS 0.00889f
C130 B.n90 VSUBS 0.00889f
C131 B.n91 VSUBS 0.00889f
C132 B.n92 VSUBS 0.00889f
C133 B.n93 VSUBS 0.00889f
C134 B.n94 VSUBS 0.00889f
C135 B.n95 VSUBS 0.00889f
C136 B.n96 VSUBS 0.00889f
C137 B.n97 VSUBS 0.00889f
C138 B.n98 VSUBS 0.00889f
C139 B.n99 VSUBS 0.00889f
C140 B.n100 VSUBS 0.022198f
C141 B.n101 VSUBS 0.023035f
C142 B.n102 VSUBS 0.023035f
C143 B.n103 VSUBS 0.00889f
C144 B.n104 VSUBS 0.00889f
C145 B.n105 VSUBS 0.00889f
C146 B.n106 VSUBS 0.00889f
C147 B.n107 VSUBS 0.00889f
C148 B.n108 VSUBS 0.00889f
C149 B.n109 VSUBS 0.00889f
C150 B.n110 VSUBS 0.00889f
C151 B.n111 VSUBS 0.00889f
C152 B.n112 VSUBS 0.00889f
C153 B.n113 VSUBS 0.00889f
C154 B.n114 VSUBS 0.00889f
C155 B.n115 VSUBS 0.00889f
C156 B.n116 VSUBS 0.00889f
C157 B.n117 VSUBS 0.00889f
C158 B.n118 VSUBS 0.00889f
C159 B.n119 VSUBS 0.00889f
C160 B.n120 VSUBS 0.006144f
C161 B.n121 VSUBS 0.020596f
C162 B.n122 VSUBS 0.00719f
C163 B.n123 VSUBS 0.00889f
C164 B.n124 VSUBS 0.00889f
C165 B.n125 VSUBS 0.00889f
C166 B.n126 VSUBS 0.00889f
C167 B.n127 VSUBS 0.00889f
C168 B.n128 VSUBS 0.00889f
C169 B.n129 VSUBS 0.00889f
C170 B.n130 VSUBS 0.00889f
C171 B.n131 VSUBS 0.00889f
C172 B.n132 VSUBS 0.00889f
C173 B.n133 VSUBS 0.00889f
C174 B.n134 VSUBS 0.00719f
C175 B.n135 VSUBS 0.020596f
C176 B.n136 VSUBS 0.006144f
C177 B.n137 VSUBS 0.00889f
C178 B.n138 VSUBS 0.00889f
C179 B.n139 VSUBS 0.00889f
C180 B.n140 VSUBS 0.00889f
C181 B.n141 VSUBS 0.00889f
C182 B.n142 VSUBS 0.00889f
C183 B.n143 VSUBS 0.00889f
C184 B.n144 VSUBS 0.00889f
C185 B.n145 VSUBS 0.00889f
C186 B.n146 VSUBS 0.00889f
C187 B.n147 VSUBS 0.00889f
C188 B.n148 VSUBS 0.00889f
C189 B.n149 VSUBS 0.00889f
C190 B.n150 VSUBS 0.00889f
C191 B.n151 VSUBS 0.00889f
C192 B.n152 VSUBS 0.00889f
C193 B.n153 VSUBS 0.00889f
C194 B.n154 VSUBS 0.022108f
C195 B.n155 VSUBS 0.023035f
C196 B.n156 VSUBS 0.022198f
C197 B.n157 VSUBS 0.00889f
C198 B.n158 VSUBS 0.00889f
C199 B.n159 VSUBS 0.00889f
C200 B.n160 VSUBS 0.00889f
C201 B.n161 VSUBS 0.00889f
C202 B.n162 VSUBS 0.00889f
C203 B.n163 VSUBS 0.00889f
C204 B.n164 VSUBS 0.00889f
C205 B.n165 VSUBS 0.00889f
C206 B.n166 VSUBS 0.00889f
C207 B.n167 VSUBS 0.00889f
C208 B.n168 VSUBS 0.00889f
C209 B.n169 VSUBS 0.00889f
C210 B.n170 VSUBS 0.00889f
C211 B.n171 VSUBS 0.00889f
C212 B.n172 VSUBS 0.00889f
C213 B.n173 VSUBS 0.00889f
C214 B.n174 VSUBS 0.00889f
C215 B.n175 VSUBS 0.00889f
C216 B.n176 VSUBS 0.00889f
C217 B.n177 VSUBS 0.00889f
C218 B.n178 VSUBS 0.00889f
C219 B.n179 VSUBS 0.00889f
C220 B.n180 VSUBS 0.00889f
C221 B.n181 VSUBS 0.00889f
C222 B.n182 VSUBS 0.00889f
C223 B.n183 VSUBS 0.00889f
C224 B.n184 VSUBS 0.00889f
C225 B.n185 VSUBS 0.00889f
C226 B.n186 VSUBS 0.00889f
C227 B.n187 VSUBS 0.00889f
C228 B.n188 VSUBS 0.00889f
C229 B.n189 VSUBS 0.00889f
C230 B.n190 VSUBS 0.00889f
C231 B.n191 VSUBS 0.00889f
C232 B.n192 VSUBS 0.00889f
C233 B.n193 VSUBS 0.00889f
C234 B.n194 VSUBS 0.00889f
C235 B.n195 VSUBS 0.00889f
C236 B.n196 VSUBS 0.00889f
C237 B.n197 VSUBS 0.00889f
C238 B.n198 VSUBS 0.00889f
C239 B.n199 VSUBS 0.00889f
C240 B.n200 VSUBS 0.00889f
C241 B.n201 VSUBS 0.00889f
C242 B.n202 VSUBS 0.00889f
C243 B.n203 VSUBS 0.00889f
C244 B.n204 VSUBS 0.00889f
C245 B.n205 VSUBS 0.022198f
C246 B.n206 VSUBS 0.022198f
C247 B.n207 VSUBS 0.023035f
C248 B.n208 VSUBS 0.00889f
C249 B.n209 VSUBS 0.00889f
C250 B.n210 VSUBS 0.00889f
C251 B.n211 VSUBS 0.00889f
C252 B.n212 VSUBS 0.00889f
C253 B.n213 VSUBS 0.00889f
C254 B.n214 VSUBS 0.00889f
C255 B.n215 VSUBS 0.00889f
C256 B.n216 VSUBS 0.00889f
C257 B.n217 VSUBS 0.00889f
C258 B.n218 VSUBS 0.00889f
C259 B.n219 VSUBS 0.00889f
C260 B.n220 VSUBS 0.00889f
C261 B.n221 VSUBS 0.00889f
C262 B.n222 VSUBS 0.00889f
C263 B.n223 VSUBS 0.00889f
C264 B.n224 VSUBS 0.00889f
C265 B.n225 VSUBS 0.006144f
C266 B.n226 VSUBS 0.020596f
C267 B.n227 VSUBS 0.00719f
C268 B.n228 VSUBS 0.00889f
C269 B.n229 VSUBS 0.00889f
C270 B.n230 VSUBS 0.00889f
C271 B.n231 VSUBS 0.00889f
C272 B.n232 VSUBS 0.00889f
C273 B.n233 VSUBS 0.00889f
C274 B.n234 VSUBS 0.00889f
C275 B.n235 VSUBS 0.00889f
C276 B.n236 VSUBS 0.00889f
C277 B.n237 VSUBS 0.00889f
C278 B.n238 VSUBS 0.00889f
C279 B.n239 VSUBS 0.00719f
C280 B.n240 VSUBS 0.00889f
C281 B.n241 VSUBS 0.00889f
C282 B.n242 VSUBS 0.00889f
C283 B.n243 VSUBS 0.00889f
C284 B.n244 VSUBS 0.00889f
C285 B.n245 VSUBS 0.00889f
C286 B.n246 VSUBS 0.00889f
C287 B.n247 VSUBS 0.00889f
C288 B.n248 VSUBS 0.00889f
C289 B.n249 VSUBS 0.00889f
C290 B.n250 VSUBS 0.00889f
C291 B.n251 VSUBS 0.00889f
C292 B.n252 VSUBS 0.00889f
C293 B.n253 VSUBS 0.00889f
C294 B.n254 VSUBS 0.00889f
C295 B.n255 VSUBS 0.00889f
C296 B.n256 VSUBS 0.00889f
C297 B.n257 VSUBS 0.00889f
C298 B.n258 VSUBS 0.00889f
C299 B.n259 VSUBS 0.023035f
C300 B.n260 VSUBS 0.022198f
C301 B.n261 VSUBS 0.022198f
C302 B.n262 VSUBS 0.00889f
C303 B.n263 VSUBS 0.00889f
C304 B.n264 VSUBS 0.00889f
C305 B.n265 VSUBS 0.00889f
C306 B.n266 VSUBS 0.00889f
C307 B.n267 VSUBS 0.00889f
C308 B.n268 VSUBS 0.00889f
C309 B.n269 VSUBS 0.00889f
C310 B.n270 VSUBS 0.00889f
C311 B.n271 VSUBS 0.00889f
C312 B.n272 VSUBS 0.00889f
C313 B.n273 VSUBS 0.00889f
C314 B.n274 VSUBS 0.00889f
C315 B.n275 VSUBS 0.00889f
C316 B.n276 VSUBS 0.00889f
C317 B.n277 VSUBS 0.00889f
C318 B.n278 VSUBS 0.00889f
C319 B.n279 VSUBS 0.00889f
C320 B.n280 VSUBS 0.00889f
C321 B.n281 VSUBS 0.00889f
C322 B.n282 VSUBS 0.00889f
C323 B.n283 VSUBS 0.0116f
C324 B.n284 VSUBS 0.012358f
C325 B.n285 VSUBS 0.024574f
C326 VDD2.t0 VSUBS 0.289107f
C327 VDD2.t1 VSUBS 0.199108f
C328 VDD2.n0 VSUBS 1.55862f
C329 VN.t1 VSUBS 0.365941f
C330 VN.t0 VSUBS 0.555363f
C331 VDD1.t1 VSUBS 0.193979f
C332 VDD1.t0 VSUBS 0.288712f
C333 VTAIL.t2 VSUBS 0.221277f
C334 VTAIL.n0 VSUBS 0.852791f
C335 VTAIL.t1 VSUBS 0.221278f
C336 VTAIL.n1 VSUBS 0.869346f
C337 VTAIL.t3 VSUBS 0.221277f
C338 VTAIL.n2 VSUBS 0.788098f
C339 VTAIL.t0 VSUBS 0.221277f
C340 VTAIL.n3 VSUBS 0.733701f
C341 VP.t0 VSUBS 0.933127f
C342 VP.t1 VSUBS 0.620128f
C343 VP.n0 VSUBS 3.3975f
.ends

