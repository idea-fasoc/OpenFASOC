* NGSPICE file created from diff_pair_sample_0775.ext - technology: sky130A

.subckt diff_pair_sample_0775 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t19 VP.t0 VDD1.t8 B.t5 sky130_fd_pr__nfet_01v8 ad=0.35475 pd=2.48 as=0.35475 ps=2.48 w=2.15 l=3.74
X1 B.t23 B.t21 B.t22 B.t11 sky130_fd_pr__nfet_01v8 ad=0.8385 pd=5.08 as=0 ps=0 w=2.15 l=3.74
X2 VTAIL.t4 VN.t0 VDD2.t9 B.t4 sky130_fd_pr__nfet_01v8 ad=0.35475 pd=2.48 as=0.35475 ps=2.48 w=2.15 l=3.74
X3 VDD2.t8 VN.t1 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=0.35475 pd=2.48 as=0.8385 ps=5.08 w=2.15 l=3.74
X4 VDD1.t5 VP.t1 VTAIL.t18 B.t7 sky130_fd_pr__nfet_01v8 ad=0.35475 pd=2.48 as=0.8385 ps=5.08 w=2.15 l=3.74
X5 VDD2.t7 VN.t2 VTAIL.t9 B.t9 sky130_fd_pr__nfet_01v8 ad=0.8385 pd=5.08 as=0.35475 ps=2.48 w=2.15 l=3.74
X6 VDD1.t3 VP.t2 VTAIL.t17 B.t6 sky130_fd_pr__nfet_01v8 ad=0.35475 pd=2.48 as=0.35475 ps=2.48 w=2.15 l=3.74
X7 VTAIL.t16 VP.t3 VDD1.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=0.35475 pd=2.48 as=0.35475 ps=2.48 w=2.15 l=3.74
X8 VTAIL.t15 VP.t4 VDD1.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.35475 pd=2.48 as=0.35475 ps=2.48 w=2.15 l=3.74
X9 VTAIL.t14 VP.t5 VDD1.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.35475 pd=2.48 as=0.35475 ps=2.48 w=2.15 l=3.74
X10 VTAIL.t2 VN.t3 VDD2.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=0.35475 pd=2.48 as=0.35475 ps=2.48 w=2.15 l=3.74
X11 VDD1.t9 VP.t6 VTAIL.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=0.8385 pd=5.08 as=0.35475 ps=2.48 w=2.15 l=3.74
X12 VDD2.t5 VN.t4 VTAIL.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=0.35475 pd=2.48 as=0.8385 ps=5.08 w=2.15 l=3.74
X13 VTAIL.t3 VN.t5 VDD2.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=0.35475 pd=2.48 as=0.35475 ps=2.48 w=2.15 l=3.74
X14 B.t20 B.t18 B.t19 B.t15 sky130_fd_pr__nfet_01v8 ad=0.8385 pd=5.08 as=0 ps=0 w=2.15 l=3.74
X15 VTAIL.t5 VN.t6 VDD2.t3 B.t5 sky130_fd_pr__nfet_01v8 ad=0.35475 pd=2.48 as=0.35475 ps=2.48 w=2.15 l=3.74
X16 VDD1.t0 VP.t7 VTAIL.t12 B.t8 sky130_fd_pr__nfet_01v8 ad=0.35475 pd=2.48 as=0.8385 ps=5.08 w=2.15 l=3.74
X17 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=0.8385 pd=5.08 as=0 ps=0 w=2.15 l=3.74
X18 VDD2.t2 VN.t7 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=0.35475 pd=2.48 as=0.35475 ps=2.48 w=2.15 l=3.74
X19 VDD1.t1 VP.t8 VTAIL.t11 B.t0 sky130_fd_pr__nfet_01v8 ad=0.8385 pd=5.08 as=0.35475 ps=2.48 w=2.15 l=3.74
X20 VDD1.t7 VP.t9 VTAIL.t10 B.t1 sky130_fd_pr__nfet_01v8 ad=0.35475 pd=2.48 as=0.35475 ps=2.48 w=2.15 l=3.74
X21 VDD2.t1 VN.t8 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.35475 pd=2.48 as=0.35475 ps=2.48 w=2.15 l=3.74
X22 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=0.8385 pd=5.08 as=0 ps=0 w=2.15 l=3.74
X23 VDD2.t0 VN.t9 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.8385 pd=5.08 as=0.35475 ps=2.48 w=2.15 l=3.74
R0 VP.n33 VP.n32 161.3
R1 VP.n34 VP.n29 161.3
R2 VP.n36 VP.n35 161.3
R3 VP.n37 VP.n28 161.3
R4 VP.n39 VP.n38 161.3
R5 VP.n40 VP.n27 161.3
R6 VP.n42 VP.n41 161.3
R7 VP.n43 VP.n26 161.3
R8 VP.n45 VP.n44 161.3
R9 VP.n46 VP.n25 161.3
R10 VP.n48 VP.n47 161.3
R11 VP.n49 VP.n24 161.3
R12 VP.n51 VP.n50 161.3
R13 VP.n52 VP.n23 161.3
R14 VP.n54 VP.n53 161.3
R15 VP.n55 VP.n22 161.3
R16 VP.n58 VP.n57 161.3
R17 VP.n59 VP.n21 161.3
R18 VP.n61 VP.n60 161.3
R19 VP.n62 VP.n20 161.3
R20 VP.n64 VP.n63 161.3
R21 VP.n65 VP.n19 161.3
R22 VP.n67 VP.n66 161.3
R23 VP.n68 VP.n18 161.3
R24 VP.n70 VP.n69 161.3
R25 VP.n125 VP.n124 161.3
R26 VP.n123 VP.n1 161.3
R27 VP.n122 VP.n121 161.3
R28 VP.n120 VP.n2 161.3
R29 VP.n119 VP.n118 161.3
R30 VP.n117 VP.n3 161.3
R31 VP.n116 VP.n115 161.3
R32 VP.n114 VP.n4 161.3
R33 VP.n113 VP.n112 161.3
R34 VP.n110 VP.n5 161.3
R35 VP.n109 VP.n108 161.3
R36 VP.n107 VP.n6 161.3
R37 VP.n106 VP.n105 161.3
R38 VP.n104 VP.n7 161.3
R39 VP.n103 VP.n102 161.3
R40 VP.n101 VP.n8 161.3
R41 VP.n100 VP.n99 161.3
R42 VP.n98 VP.n9 161.3
R43 VP.n97 VP.n96 161.3
R44 VP.n95 VP.n10 161.3
R45 VP.n94 VP.n93 161.3
R46 VP.n92 VP.n11 161.3
R47 VP.n91 VP.n90 161.3
R48 VP.n89 VP.n12 161.3
R49 VP.n88 VP.n87 161.3
R50 VP.n85 VP.n13 161.3
R51 VP.n84 VP.n83 161.3
R52 VP.n82 VP.n14 161.3
R53 VP.n81 VP.n80 161.3
R54 VP.n79 VP.n15 161.3
R55 VP.n78 VP.n77 161.3
R56 VP.n76 VP.n16 161.3
R57 VP.n75 VP.n74 161.3
R58 VP.n73 VP.n72 83.2166
R59 VP.n126 VP.n0 83.2166
R60 VP.n71 VP.n17 83.2166
R61 VP.n31 VP.n30 71.3788
R62 VP.n72 VP.n71 51.9501
R63 VP.n80 VP.n79 50.6917
R64 VP.n118 VP.n2 50.6917
R65 VP.n63 VP.n19 50.6917
R66 VP.n30 VP.t8 46.66
R67 VP.n93 VP.n92 43.8928
R68 VP.n105 VP.n6 43.8928
R69 VP.n50 VP.n23 43.8928
R70 VP.n38 VP.n37 43.8928
R71 VP.n93 VP.n10 37.094
R72 VP.n105 VP.n104 37.094
R73 VP.n50 VP.n49 37.094
R74 VP.n38 VP.n27 37.094
R75 VP.n80 VP.n14 30.2951
R76 VP.n118 VP.n117 30.2951
R77 VP.n63 VP.n62 30.2951
R78 VP.n74 VP.n16 24.4675
R79 VP.n78 VP.n16 24.4675
R80 VP.n79 VP.n78 24.4675
R81 VP.n84 VP.n14 24.4675
R82 VP.n85 VP.n84 24.4675
R83 VP.n87 VP.n12 24.4675
R84 VP.n91 VP.n12 24.4675
R85 VP.n92 VP.n91 24.4675
R86 VP.n97 VP.n10 24.4675
R87 VP.n98 VP.n97 24.4675
R88 VP.n99 VP.n98 24.4675
R89 VP.n99 VP.n8 24.4675
R90 VP.n103 VP.n8 24.4675
R91 VP.n104 VP.n103 24.4675
R92 VP.n109 VP.n6 24.4675
R93 VP.n110 VP.n109 24.4675
R94 VP.n112 VP.n110 24.4675
R95 VP.n116 VP.n4 24.4675
R96 VP.n117 VP.n116 24.4675
R97 VP.n122 VP.n2 24.4675
R98 VP.n123 VP.n122 24.4675
R99 VP.n124 VP.n123 24.4675
R100 VP.n67 VP.n19 24.4675
R101 VP.n68 VP.n67 24.4675
R102 VP.n69 VP.n68 24.4675
R103 VP.n54 VP.n23 24.4675
R104 VP.n55 VP.n54 24.4675
R105 VP.n57 VP.n55 24.4675
R106 VP.n61 VP.n21 24.4675
R107 VP.n62 VP.n61 24.4675
R108 VP.n42 VP.n27 24.4675
R109 VP.n43 VP.n42 24.4675
R110 VP.n44 VP.n43 24.4675
R111 VP.n44 VP.n25 24.4675
R112 VP.n48 VP.n25 24.4675
R113 VP.n49 VP.n48 24.4675
R114 VP.n32 VP.n29 24.4675
R115 VP.n36 VP.n29 24.4675
R116 VP.n37 VP.n36 24.4675
R117 VP.n86 VP.n85 21.0421
R118 VP.n111 VP.n4 21.0421
R119 VP.n56 VP.n21 21.0421
R120 VP.n99 VP.t2 13.8548
R121 VP.n73 VP.t6 13.8548
R122 VP.n86 VP.t4 13.8548
R123 VP.n111 VP.t3 13.8548
R124 VP.n0 VP.t7 13.8548
R125 VP.n44 VP.t9 13.8548
R126 VP.n17 VP.t1 13.8548
R127 VP.n56 VP.t5 13.8548
R128 VP.n31 VP.t0 13.8548
R129 VP.n74 VP.n73 6.85126
R130 VP.n124 VP.n0 6.85126
R131 VP.n69 VP.n17 6.85126
R132 VP.n87 VP.n86 3.42588
R133 VP.n112 VP.n111 3.42588
R134 VP.n57 VP.n56 3.42588
R135 VP.n32 VP.n31 3.42588
R136 VP.n33 VP.n30 3.25232
R137 VP.n71 VP.n70 0.354971
R138 VP.n75 VP.n72 0.354971
R139 VP.n126 VP.n125 0.354971
R140 VP VP.n126 0.26696
R141 VP.n34 VP.n33 0.189894
R142 VP.n35 VP.n34 0.189894
R143 VP.n35 VP.n28 0.189894
R144 VP.n39 VP.n28 0.189894
R145 VP.n40 VP.n39 0.189894
R146 VP.n41 VP.n40 0.189894
R147 VP.n41 VP.n26 0.189894
R148 VP.n45 VP.n26 0.189894
R149 VP.n46 VP.n45 0.189894
R150 VP.n47 VP.n46 0.189894
R151 VP.n47 VP.n24 0.189894
R152 VP.n51 VP.n24 0.189894
R153 VP.n52 VP.n51 0.189894
R154 VP.n53 VP.n52 0.189894
R155 VP.n53 VP.n22 0.189894
R156 VP.n58 VP.n22 0.189894
R157 VP.n59 VP.n58 0.189894
R158 VP.n60 VP.n59 0.189894
R159 VP.n60 VP.n20 0.189894
R160 VP.n64 VP.n20 0.189894
R161 VP.n65 VP.n64 0.189894
R162 VP.n66 VP.n65 0.189894
R163 VP.n66 VP.n18 0.189894
R164 VP.n70 VP.n18 0.189894
R165 VP.n76 VP.n75 0.189894
R166 VP.n77 VP.n76 0.189894
R167 VP.n77 VP.n15 0.189894
R168 VP.n81 VP.n15 0.189894
R169 VP.n82 VP.n81 0.189894
R170 VP.n83 VP.n82 0.189894
R171 VP.n83 VP.n13 0.189894
R172 VP.n88 VP.n13 0.189894
R173 VP.n89 VP.n88 0.189894
R174 VP.n90 VP.n89 0.189894
R175 VP.n90 VP.n11 0.189894
R176 VP.n94 VP.n11 0.189894
R177 VP.n95 VP.n94 0.189894
R178 VP.n96 VP.n95 0.189894
R179 VP.n96 VP.n9 0.189894
R180 VP.n100 VP.n9 0.189894
R181 VP.n101 VP.n100 0.189894
R182 VP.n102 VP.n101 0.189894
R183 VP.n102 VP.n7 0.189894
R184 VP.n106 VP.n7 0.189894
R185 VP.n107 VP.n106 0.189894
R186 VP.n108 VP.n107 0.189894
R187 VP.n108 VP.n5 0.189894
R188 VP.n113 VP.n5 0.189894
R189 VP.n114 VP.n113 0.189894
R190 VP.n115 VP.n114 0.189894
R191 VP.n115 VP.n3 0.189894
R192 VP.n119 VP.n3 0.189894
R193 VP.n120 VP.n119 0.189894
R194 VP.n121 VP.n120 0.189894
R195 VP.n121 VP.n1 0.189894
R196 VP.n125 VP.n1 0.189894
R197 VDD1.n3 VDD1.t9 105.603
R198 VDD1.n1 VDD1.t1 105.603
R199 VDD1.n5 VDD1.n4 95.4617
R200 VDD1.n1 VDD1.n0 92.8859
R201 VDD1.n7 VDD1.n6 92.8858
R202 VDD1.n3 VDD1.n2 92.8856
R203 VDD1.n7 VDD1.n5 44.572
R204 VDD1.n6 VDD1.t4 9.2098
R205 VDD1.n6 VDD1.t5 9.2098
R206 VDD1.n0 VDD1.t8 9.2098
R207 VDD1.n0 VDD1.t7 9.2098
R208 VDD1.n4 VDD1.t6 9.2098
R209 VDD1.n4 VDD1.t0 9.2098
R210 VDD1.n2 VDD1.t2 9.2098
R211 VDD1.n2 VDD1.t3 9.2098
R212 VDD1 VDD1.n7 2.57378
R213 VDD1 VDD1.n1 0.935845
R214 VDD1.n5 VDD1.n3 0.822309
R215 VTAIL.n17 VTAIL.t7 85.4163
R216 VTAIL.n2 VTAIL.t12 85.4163
R217 VTAIL.n16 VTAIL.t18 85.4163
R218 VTAIL.n11 VTAIL.t8 85.4162
R219 VTAIL.n15 VTAIL.n14 76.2071
R220 VTAIL.n13 VTAIL.n12 76.2071
R221 VTAIL.n10 VTAIL.n9 76.2071
R222 VTAIL.n8 VTAIL.n7 76.2071
R223 VTAIL.n19 VTAIL.n18 76.2068
R224 VTAIL.n1 VTAIL.n0 76.2068
R225 VTAIL.n4 VTAIL.n3 76.2068
R226 VTAIL.n6 VTAIL.n5 76.2068
R227 VTAIL.n8 VTAIL.n6 21.2376
R228 VTAIL.n17 VTAIL.n16 17.7289
R229 VTAIL.n18 VTAIL.t1 9.2098
R230 VTAIL.n18 VTAIL.t4 9.2098
R231 VTAIL.n0 VTAIL.t0 9.2098
R232 VTAIL.n0 VTAIL.t5 9.2098
R233 VTAIL.n3 VTAIL.t17 9.2098
R234 VTAIL.n3 VTAIL.t16 9.2098
R235 VTAIL.n5 VTAIL.t13 9.2098
R236 VTAIL.n5 VTAIL.t15 9.2098
R237 VTAIL.n14 VTAIL.t10 9.2098
R238 VTAIL.n14 VTAIL.t14 9.2098
R239 VTAIL.n12 VTAIL.t11 9.2098
R240 VTAIL.n12 VTAIL.t19 9.2098
R241 VTAIL.n9 VTAIL.t6 9.2098
R242 VTAIL.n9 VTAIL.t3 9.2098
R243 VTAIL.n7 VTAIL.t9 9.2098
R244 VTAIL.n7 VTAIL.t2 9.2098
R245 VTAIL.n10 VTAIL.n8 3.50912
R246 VTAIL.n11 VTAIL.n10 3.50912
R247 VTAIL.n15 VTAIL.n13 3.50912
R248 VTAIL.n16 VTAIL.n15 3.50912
R249 VTAIL.n6 VTAIL.n4 3.50912
R250 VTAIL.n4 VTAIL.n2 3.50912
R251 VTAIL.n19 VTAIL.n17 3.50912
R252 VTAIL VTAIL.n1 2.69016
R253 VTAIL.n13 VTAIL.n11 2.22464
R254 VTAIL.n2 VTAIL.n1 2.22464
R255 VTAIL VTAIL.n19 0.819465
R256 B.n828 B.n827 585
R257 B.n829 B.n828 585
R258 B.n234 B.n163 585
R259 B.n233 B.n232 585
R260 B.n231 B.n230 585
R261 B.n229 B.n228 585
R262 B.n227 B.n226 585
R263 B.n225 B.n224 585
R264 B.n223 B.n222 585
R265 B.n221 B.n220 585
R266 B.n219 B.n218 585
R267 B.n217 B.n216 585
R268 B.n215 B.n214 585
R269 B.n213 B.n212 585
R270 B.n211 B.n210 585
R271 B.n209 B.n208 585
R272 B.n207 B.n206 585
R273 B.n205 B.n204 585
R274 B.n203 B.n202 585
R275 B.n201 B.n200 585
R276 B.n199 B.n198 585
R277 B.n197 B.n196 585
R278 B.n195 B.n194 585
R279 B.n192 B.n191 585
R280 B.n190 B.n189 585
R281 B.n188 B.n187 585
R282 B.n186 B.n185 585
R283 B.n184 B.n183 585
R284 B.n182 B.n181 585
R285 B.n180 B.n179 585
R286 B.n178 B.n177 585
R287 B.n176 B.n175 585
R288 B.n174 B.n173 585
R289 B.n172 B.n171 585
R290 B.n170 B.n169 585
R291 B.n144 B.n143 585
R292 B.n826 B.n145 585
R293 B.n830 B.n145 585
R294 B.n825 B.n824 585
R295 B.n824 B.n141 585
R296 B.n823 B.n140 585
R297 B.n836 B.n140 585
R298 B.n822 B.n139 585
R299 B.n837 B.n139 585
R300 B.n821 B.n138 585
R301 B.n838 B.n138 585
R302 B.n820 B.n819 585
R303 B.n819 B.n134 585
R304 B.n818 B.n133 585
R305 B.n844 B.n133 585
R306 B.n817 B.n132 585
R307 B.n845 B.n132 585
R308 B.n816 B.n131 585
R309 B.n846 B.n131 585
R310 B.n815 B.n814 585
R311 B.n814 B.n130 585
R312 B.n813 B.n126 585
R313 B.n852 B.n126 585
R314 B.n812 B.n125 585
R315 B.n853 B.n125 585
R316 B.n811 B.n124 585
R317 B.n854 B.n124 585
R318 B.n810 B.n809 585
R319 B.n809 B.n120 585
R320 B.n808 B.n119 585
R321 B.n860 B.n119 585
R322 B.n807 B.n118 585
R323 B.n861 B.n118 585
R324 B.n806 B.n117 585
R325 B.n862 B.n117 585
R326 B.n805 B.n804 585
R327 B.n804 B.n113 585
R328 B.n803 B.n112 585
R329 B.n868 B.n112 585
R330 B.n802 B.n111 585
R331 B.n869 B.n111 585
R332 B.n801 B.n110 585
R333 B.n870 B.n110 585
R334 B.n800 B.n799 585
R335 B.n799 B.n106 585
R336 B.n798 B.n105 585
R337 B.n876 B.n105 585
R338 B.n797 B.n104 585
R339 B.n877 B.n104 585
R340 B.n796 B.n103 585
R341 B.n878 B.n103 585
R342 B.n795 B.n794 585
R343 B.n794 B.n99 585
R344 B.n793 B.n98 585
R345 B.n884 B.n98 585
R346 B.n792 B.n97 585
R347 B.n885 B.n97 585
R348 B.n791 B.n96 585
R349 B.n886 B.n96 585
R350 B.n790 B.n789 585
R351 B.n789 B.n92 585
R352 B.n788 B.n91 585
R353 B.n892 B.n91 585
R354 B.n787 B.n90 585
R355 B.n893 B.n90 585
R356 B.n786 B.n89 585
R357 B.n894 B.n89 585
R358 B.n785 B.n784 585
R359 B.n784 B.n85 585
R360 B.n783 B.n84 585
R361 B.n900 B.n84 585
R362 B.n782 B.n83 585
R363 B.n901 B.n83 585
R364 B.n781 B.n82 585
R365 B.n902 B.n82 585
R366 B.n780 B.n779 585
R367 B.n779 B.n78 585
R368 B.n778 B.n77 585
R369 B.n908 B.n77 585
R370 B.n777 B.n76 585
R371 B.n909 B.n76 585
R372 B.n776 B.n75 585
R373 B.n910 B.n75 585
R374 B.n775 B.n774 585
R375 B.n774 B.n71 585
R376 B.n773 B.n70 585
R377 B.n916 B.n70 585
R378 B.n772 B.n69 585
R379 B.n917 B.n69 585
R380 B.n771 B.n68 585
R381 B.n918 B.n68 585
R382 B.n770 B.n769 585
R383 B.n769 B.n64 585
R384 B.n768 B.n63 585
R385 B.n924 B.n63 585
R386 B.n767 B.n62 585
R387 B.n925 B.n62 585
R388 B.n766 B.n61 585
R389 B.n926 B.n61 585
R390 B.n765 B.n764 585
R391 B.n764 B.n57 585
R392 B.n763 B.n56 585
R393 B.n932 B.n56 585
R394 B.n762 B.n55 585
R395 B.n933 B.n55 585
R396 B.n761 B.n54 585
R397 B.n934 B.n54 585
R398 B.n760 B.n759 585
R399 B.n759 B.n50 585
R400 B.n758 B.n49 585
R401 B.n940 B.n49 585
R402 B.n757 B.n48 585
R403 B.n941 B.n48 585
R404 B.n756 B.n47 585
R405 B.n942 B.n47 585
R406 B.n755 B.n754 585
R407 B.n754 B.n43 585
R408 B.n753 B.n42 585
R409 B.n948 B.n42 585
R410 B.n752 B.n41 585
R411 B.n949 B.n41 585
R412 B.n751 B.n40 585
R413 B.n950 B.n40 585
R414 B.n750 B.n749 585
R415 B.n749 B.n36 585
R416 B.n748 B.n35 585
R417 B.n956 B.n35 585
R418 B.n747 B.n34 585
R419 B.n957 B.n34 585
R420 B.n746 B.n33 585
R421 B.n958 B.n33 585
R422 B.n745 B.n744 585
R423 B.n744 B.n29 585
R424 B.n743 B.n28 585
R425 B.n964 B.n28 585
R426 B.n742 B.n27 585
R427 B.n965 B.n27 585
R428 B.n741 B.n26 585
R429 B.n966 B.n26 585
R430 B.n740 B.n739 585
R431 B.n739 B.n22 585
R432 B.n738 B.n21 585
R433 B.n972 B.n21 585
R434 B.n737 B.n20 585
R435 B.n973 B.n20 585
R436 B.n736 B.n19 585
R437 B.n974 B.n19 585
R438 B.n735 B.n734 585
R439 B.n734 B.n15 585
R440 B.n733 B.n14 585
R441 B.n980 B.n14 585
R442 B.n732 B.n13 585
R443 B.n981 B.n13 585
R444 B.n731 B.n12 585
R445 B.n982 B.n12 585
R446 B.n730 B.n729 585
R447 B.n729 B.n8 585
R448 B.n728 B.n7 585
R449 B.n988 B.n7 585
R450 B.n727 B.n6 585
R451 B.n989 B.n6 585
R452 B.n726 B.n5 585
R453 B.n990 B.n5 585
R454 B.n725 B.n724 585
R455 B.n724 B.n4 585
R456 B.n723 B.n235 585
R457 B.n723 B.n722 585
R458 B.n713 B.n236 585
R459 B.n237 B.n236 585
R460 B.n715 B.n714 585
R461 B.n716 B.n715 585
R462 B.n712 B.n242 585
R463 B.n242 B.n241 585
R464 B.n711 B.n710 585
R465 B.n710 B.n709 585
R466 B.n244 B.n243 585
R467 B.n245 B.n244 585
R468 B.n702 B.n701 585
R469 B.n703 B.n702 585
R470 B.n700 B.n250 585
R471 B.n250 B.n249 585
R472 B.n699 B.n698 585
R473 B.n698 B.n697 585
R474 B.n252 B.n251 585
R475 B.n253 B.n252 585
R476 B.n690 B.n689 585
R477 B.n691 B.n690 585
R478 B.n688 B.n258 585
R479 B.n258 B.n257 585
R480 B.n687 B.n686 585
R481 B.n686 B.n685 585
R482 B.n260 B.n259 585
R483 B.n261 B.n260 585
R484 B.n678 B.n677 585
R485 B.n679 B.n678 585
R486 B.n676 B.n266 585
R487 B.n266 B.n265 585
R488 B.n675 B.n674 585
R489 B.n674 B.n673 585
R490 B.n268 B.n267 585
R491 B.n269 B.n268 585
R492 B.n666 B.n665 585
R493 B.n667 B.n666 585
R494 B.n664 B.n274 585
R495 B.n274 B.n273 585
R496 B.n663 B.n662 585
R497 B.n662 B.n661 585
R498 B.n276 B.n275 585
R499 B.n277 B.n276 585
R500 B.n654 B.n653 585
R501 B.n655 B.n654 585
R502 B.n652 B.n282 585
R503 B.n282 B.n281 585
R504 B.n651 B.n650 585
R505 B.n650 B.n649 585
R506 B.n284 B.n283 585
R507 B.n285 B.n284 585
R508 B.n642 B.n641 585
R509 B.n643 B.n642 585
R510 B.n640 B.n290 585
R511 B.n290 B.n289 585
R512 B.n639 B.n638 585
R513 B.n638 B.n637 585
R514 B.n292 B.n291 585
R515 B.n293 B.n292 585
R516 B.n630 B.n629 585
R517 B.n631 B.n630 585
R518 B.n628 B.n298 585
R519 B.n298 B.n297 585
R520 B.n627 B.n626 585
R521 B.n626 B.n625 585
R522 B.n300 B.n299 585
R523 B.n301 B.n300 585
R524 B.n618 B.n617 585
R525 B.n619 B.n618 585
R526 B.n616 B.n306 585
R527 B.n306 B.n305 585
R528 B.n615 B.n614 585
R529 B.n614 B.n613 585
R530 B.n308 B.n307 585
R531 B.n309 B.n308 585
R532 B.n606 B.n605 585
R533 B.n607 B.n606 585
R534 B.n604 B.n314 585
R535 B.n314 B.n313 585
R536 B.n603 B.n602 585
R537 B.n602 B.n601 585
R538 B.n316 B.n315 585
R539 B.n317 B.n316 585
R540 B.n594 B.n593 585
R541 B.n595 B.n594 585
R542 B.n592 B.n322 585
R543 B.n322 B.n321 585
R544 B.n591 B.n590 585
R545 B.n590 B.n589 585
R546 B.n324 B.n323 585
R547 B.n325 B.n324 585
R548 B.n582 B.n581 585
R549 B.n583 B.n582 585
R550 B.n580 B.n330 585
R551 B.n330 B.n329 585
R552 B.n579 B.n578 585
R553 B.n578 B.n577 585
R554 B.n332 B.n331 585
R555 B.n333 B.n332 585
R556 B.n570 B.n569 585
R557 B.n571 B.n570 585
R558 B.n568 B.n338 585
R559 B.n338 B.n337 585
R560 B.n567 B.n566 585
R561 B.n566 B.n565 585
R562 B.n340 B.n339 585
R563 B.n341 B.n340 585
R564 B.n558 B.n557 585
R565 B.n559 B.n558 585
R566 B.n556 B.n346 585
R567 B.n346 B.n345 585
R568 B.n555 B.n554 585
R569 B.n554 B.n553 585
R570 B.n348 B.n347 585
R571 B.n349 B.n348 585
R572 B.n546 B.n545 585
R573 B.n547 B.n546 585
R574 B.n544 B.n354 585
R575 B.n354 B.n353 585
R576 B.n543 B.n542 585
R577 B.n542 B.n541 585
R578 B.n356 B.n355 585
R579 B.n357 B.n356 585
R580 B.n534 B.n533 585
R581 B.n535 B.n534 585
R582 B.n532 B.n362 585
R583 B.n362 B.n361 585
R584 B.n531 B.n530 585
R585 B.n530 B.n529 585
R586 B.n364 B.n363 585
R587 B.n365 B.n364 585
R588 B.n522 B.n521 585
R589 B.n523 B.n522 585
R590 B.n520 B.n370 585
R591 B.n370 B.n369 585
R592 B.n519 B.n518 585
R593 B.n518 B.n517 585
R594 B.n372 B.n371 585
R595 B.n510 B.n372 585
R596 B.n509 B.n508 585
R597 B.n511 B.n509 585
R598 B.n507 B.n377 585
R599 B.n377 B.n376 585
R600 B.n506 B.n505 585
R601 B.n505 B.n504 585
R602 B.n379 B.n378 585
R603 B.n380 B.n379 585
R604 B.n497 B.n496 585
R605 B.n498 B.n497 585
R606 B.n495 B.n385 585
R607 B.n385 B.n384 585
R608 B.n494 B.n493 585
R609 B.n493 B.n492 585
R610 B.n387 B.n386 585
R611 B.n388 B.n387 585
R612 B.n485 B.n484 585
R613 B.n486 B.n485 585
R614 B.n391 B.n390 585
R615 B.n417 B.n416 585
R616 B.n418 B.n414 585
R617 B.n414 B.n392 585
R618 B.n420 B.n419 585
R619 B.n422 B.n413 585
R620 B.n425 B.n424 585
R621 B.n426 B.n412 585
R622 B.n428 B.n427 585
R623 B.n430 B.n411 585
R624 B.n433 B.n432 585
R625 B.n434 B.n410 585
R626 B.n436 B.n435 585
R627 B.n438 B.n409 585
R628 B.n441 B.n440 585
R629 B.n442 B.n405 585
R630 B.n444 B.n443 585
R631 B.n446 B.n404 585
R632 B.n449 B.n448 585
R633 B.n450 B.n403 585
R634 B.n452 B.n451 585
R635 B.n454 B.n402 585
R636 B.n457 B.n456 585
R637 B.n459 B.n399 585
R638 B.n461 B.n460 585
R639 B.n463 B.n398 585
R640 B.n466 B.n465 585
R641 B.n467 B.n397 585
R642 B.n469 B.n468 585
R643 B.n471 B.n396 585
R644 B.n474 B.n473 585
R645 B.n475 B.n395 585
R646 B.n477 B.n476 585
R647 B.n479 B.n394 585
R648 B.n482 B.n481 585
R649 B.n483 B.n393 585
R650 B.n488 B.n487 585
R651 B.n487 B.n486 585
R652 B.n489 B.n389 585
R653 B.n389 B.n388 585
R654 B.n491 B.n490 585
R655 B.n492 B.n491 585
R656 B.n383 B.n382 585
R657 B.n384 B.n383 585
R658 B.n500 B.n499 585
R659 B.n499 B.n498 585
R660 B.n501 B.n381 585
R661 B.n381 B.n380 585
R662 B.n503 B.n502 585
R663 B.n504 B.n503 585
R664 B.n375 B.n374 585
R665 B.n376 B.n375 585
R666 B.n513 B.n512 585
R667 B.n512 B.n511 585
R668 B.n514 B.n373 585
R669 B.n510 B.n373 585
R670 B.n516 B.n515 585
R671 B.n517 B.n516 585
R672 B.n368 B.n367 585
R673 B.n369 B.n368 585
R674 B.n525 B.n524 585
R675 B.n524 B.n523 585
R676 B.n526 B.n366 585
R677 B.n366 B.n365 585
R678 B.n528 B.n527 585
R679 B.n529 B.n528 585
R680 B.n360 B.n359 585
R681 B.n361 B.n360 585
R682 B.n537 B.n536 585
R683 B.n536 B.n535 585
R684 B.n538 B.n358 585
R685 B.n358 B.n357 585
R686 B.n540 B.n539 585
R687 B.n541 B.n540 585
R688 B.n352 B.n351 585
R689 B.n353 B.n352 585
R690 B.n549 B.n548 585
R691 B.n548 B.n547 585
R692 B.n550 B.n350 585
R693 B.n350 B.n349 585
R694 B.n552 B.n551 585
R695 B.n553 B.n552 585
R696 B.n344 B.n343 585
R697 B.n345 B.n344 585
R698 B.n561 B.n560 585
R699 B.n560 B.n559 585
R700 B.n562 B.n342 585
R701 B.n342 B.n341 585
R702 B.n564 B.n563 585
R703 B.n565 B.n564 585
R704 B.n336 B.n335 585
R705 B.n337 B.n336 585
R706 B.n573 B.n572 585
R707 B.n572 B.n571 585
R708 B.n574 B.n334 585
R709 B.n334 B.n333 585
R710 B.n576 B.n575 585
R711 B.n577 B.n576 585
R712 B.n328 B.n327 585
R713 B.n329 B.n328 585
R714 B.n585 B.n584 585
R715 B.n584 B.n583 585
R716 B.n586 B.n326 585
R717 B.n326 B.n325 585
R718 B.n588 B.n587 585
R719 B.n589 B.n588 585
R720 B.n320 B.n319 585
R721 B.n321 B.n320 585
R722 B.n597 B.n596 585
R723 B.n596 B.n595 585
R724 B.n598 B.n318 585
R725 B.n318 B.n317 585
R726 B.n600 B.n599 585
R727 B.n601 B.n600 585
R728 B.n312 B.n311 585
R729 B.n313 B.n312 585
R730 B.n609 B.n608 585
R731 B.n608 B.n607 585
R732 B.n610 B.n310 585
R733 B.n310 B.n309 585
R734 B.n612 B.n611 585
R735 B.n613 B.n612 585
R736 B.n304 B.n303 585
R737 B.n305 B.n304 585
R738 B.n621 B.n620 585
R739 B.n620 B.n619 585
R740 B.n622 B.n302 585
R741 B.n302 B.n301 585
R742 B.n624 B.n623 585
R743 B.n625 B.n624 585
R744 B.n296 B.n295 585
R745 B.n297 B.n296 585
R746 B.n633 B.n632 585
R747 B.n632 B.n631 585
R748 B.n634 B.n294 585
R749 B.n294 B.n293 585
R750 B.n636 B.n635 585
R751 B.n637 B.n636 585
R752 B.n288 B.n287 585
R753 B.n289 B.n288 585
R754 B.n645 B.n644 585
R755 B.n644 B.n643 585
R756 B.n646 B.n286 585
R757 B.n286 B.n285 585
R758 B.n648 B.n647 585
R759 B.n649 B.n648 585
R760 B.n280 B.n279 585
R761 B.n281 B.n280 585
R762 B.n657 B.n656 585
R763 B.n656 B.n655 585
R764 B.n658 B.n278 585
R765 B.n278 B.n277 585
R766 B.n660 B.n659 585
R767 B.n661 B.n660 585
R768 B.n272 B.n271 585
R769 B.n273 B.n272 585
R770 B.n669 B.n668 585
R771 B.n668 B.n667 585
R772 B.n670 B.n270 585
R773 B.n270 B.n269 585
R774 B.n672 B.n671 585
R775 B.n673 B.n672 585
R776 B.n264 B.n263 585
R777 B.n265 B.n264 585
R778 B.n681 B.n680 585
R779 B.n680 B.n679 585
R780 B.n682 B.n262 585
R781 B.n262 B.n261 585
R782 B.n684 B.n683 585
R783 B.n685 B.n684 585
R784 B.n256 B.n255 585
R785 B.n257 B.n256 585
R786 B.n693 B.n692 585
R787 B.n692 B.n691 585
R788 B.n694 B.n254 585
R789 B.n254 B.n253 585
R790 B.n696 B.n695 585
R791 B.n697 B.n696 585
R792 B.n248 B.n247 585
R793 B.n249 B.n248 585
R794 B.n705 B.n704 585
R795 B.n704 B.n703 585
R796 B.n706 B.n246 585
R797 B.n246 B.n245 585
R798 B.n708 B.n707 585
R799 B.n709 B.n708 585
R800 B.n240 B.n239 585
R801 B.n241 B.n240 585
R802 B.n718 B.n717 585
R803 B.n717 B.n716 585
R804 B.n719 B.n238 585
R805 B.n238 B.n237 585
R806 B.n721 B.n720 585
R807 B.n722 B.n721 585
R808 B.n2 B.n0 585
R809 B.n4 B.n2 585
R810 B.n3 B.n1 585
R811 B.n989 B.n3 585
R812 B.n987 B.n986 585
R813 B.n988 B.n987 585
R814 B.n985 B.n9 585
R815 B.n9 B.n8 585
R816 B.n984 B.n983 585
R817 B.n983 B.n982 585
R818 B.n11 B.n10 585
R819 B.n981 B.n11 585
R820 B.n979 B.n978 585
R821 B.n980 B.n979 585
R822 B.n977 B.n16 585
R823 B.n16 B.n15 585
R824 B.n976 B.n975 585
R825 B.n975 B.n974 585
R826 B.n18 B.n17 585
R827 B.n973 B.n18 585
R828 B.n971 B.n970 585
R829 B.n972 B.n971 585
R830 B.n969 B.n23 585
R831 B.n23 B.n22 585
R832 B.n968 B.n967 585
R833 B.n967 B.n966 585
R834 B.n25 B.n24 585
R835 B.n965 B.n25 585
R836 B.n963 B.n962 585
R837 B.n964 B.n963 585
R838 B.n961 B.n30 585
R839 B.n30 B.n29 585
R840 B.n960 B.n959 585
R841 B.n959 B.n958 585
R842 B.n32 B.n31 585
R843 B.n957 B.n32 585
R844 B.n955 B.n954 585
R845 B.n956 B.n955 585
R846 B.n953 B.n37 585
R847 B.n37 B.n36 585
R848 B.n952 B.n951 585
R849 B.n951 B.n950 585
R850 B.n39 B.n38 585
R851 B.n949 B.n39 585
R852 B.n947 B.n946 585
R853 B.n948 B.n947 585
R854 B.n945 B.n44 585
R855 B.n44 B.n43 585
R856 B.n944 B.n943 585
R857 B.n943 B.n942 585
R858 B.n46 B.n45 585
R859 B.n941 B.n46 585
R860 B.n939 B.n938 585
R861 B.n940 B.n939 585
R862 B.n937 B.n51 585
R863 B.n51 B.n50 585
R864 B.n936 B.n935 585
R865 B.n935 B.n934 585
R866 B.n53 B.n52 585
R867 B.n933 B.n53 585
R868 B.n931 B.n930 585
R869 B.n932 B.n931 585
R870 B.n929 B.n58 585
R871 B.n58 B.n57 585
R872 B.n928 B.n927 585
R873 B.n927 B.n926 585
R874 B.n60 B.n59 585
R875 B.n925 B.n60 585
R876 B.n923 B.n922 585
R877 B.n924 B.n923 585
R878 B.n921 B.n65 585
R879 B.n65 B.n64 585
R880 B.n920 B.n919 585
R881 B.n919 B.n918 585
R882 B.n67 B.n66 585
R883 B.n917 B.n67 585
R884 B.n915 B.n914 585
R885 B.n916 B.n915 585
R886 B.n913 B.n72 585
R887 B.n72 B.n71 585
R888 B.n912 B.n911 585
R889 B.n911 B.n910 585
R890 B.n74 B.n73 585
R891 B.n909 B.n74 585
R892 B.n907 B.n906 585
R893 B.n908 B.n907 585
R894 B.n905 B.n79 585
R895 B.n79 B.n78 585
R896 B.n904 B.n903 585
R897 B.n903 B.n902 585
R898 B.n81 B.n80 585
R899 B.n901 B.n81 585
R900 B.n899 B.n898 585
R901 B.n900 B.n899 585
R902 B.n897 B.n86 585
R903 B.n86 B.n85 585
R904 B.n896 B.n895 585
R905 B.n895 B.n894 585
R906 B.n88 B.n87 585
R907 B.n893 B.n88 585
R908 B.n891 B.n890 585
R909 B.n892 B.n891 585
R910 B.n889 B.n93 585
R911 B.n93 B.n92 585
R912 B.n888 B.n887 585
R913 B.n887 B.n886 585
R914 B.n95 B.n94 585
R915 B.n885 B.n95 585
R916 B.n883 B.n882 585
R917 B.n884 B.n883 585
R918 B.n881 B.n100 585
R919 B.n100 B.n99 585
R920 B.n880 B.n879 585
R921 B.n879 B.n878 585
R922 B.n102 B.n101 585
R923 B.n877 B.n102 585
R924 B.n875 B.n874 585
R925 B.n876 B.n875 585
R926 B.n873 B.n107 585
R927 B.n107 B.n106 585
R928 B.n872 B.n871 585
R929 B.n871 B.n870 585
R930 B.n109 B.n108 585
R931 B.n869 B.n109 585
R932 B.n867 B.n866 585
R933 B.n868 B.n867 585
R934 B.n865 B.n114 585
R935 B.n114 B.n113 585
R936 B.n864 B.n863 585
R937 B.n863 B.n862 585
R938 B.n116 B.n115 585
R939 B.n861 B.n116 585
R940 B.n859 B.n858 585
R941 B.n860 B.n859 585
R942 B.n857 B.n121 585
R943 B.n121 B.n120 585
R944 B.n856 B.n855 585
R945 B.n855 B.n854 585
R946 B.n123 B.n122 585
R947 B.n853 B.n123 585
R948 B.n851 B.n850 585
R949 B.n852 B.n851 585
R950 B.n849 B.n127 585
R951 B.n130 B.n127 585
R952 B.n848 B.n847 585
R953 B.n847 B.n846 585
R954 B.n129 B.n128 585
R955 B.n845 B.n129 585
R956 B.n843 B.n842 585
R957 B.n844 B.n843 585
R958 B.n841 B.n135 585
R959 B.n135 B.n134 585
R960 B.n840 B.n839 585
R961 B.n839 B.n838 585
R962 B.n137 B.n136 585
R963 B.n837 B.n137 585
R964 B.n835 B.n834 585
R965 B.n836 B.n835 585
R966 B.n833 B.n142 585
R967 B.n142 B.n141 585
R968 B.n832 B.n831 585
R969 B.n831 B.n830 585
R970 B.n992 B.n991 585
R971 B.n991 B.n990 585
R972 B.n487 B.n391 478.086
R973 B.n831 B.n144 478.086
R974 B.n485 B.n393 478.086
R975 B.n828 B.n145 478.086
R976 B.n829 B.n162 256.663
R977 B.n829 B.n161 256.663
R978 B.n829 B.n160 256.663
R979 B.n829 B.n159 256.663
R980 B.n829 B.n158 256.663
R981 B.n829 B.n157 256.663
R982 B.n829 B.n156 256.663
R983 B.n829 B.n155 256.663
R984 B.n829 B.n154 256.663
R985 B.n829 B.n153 256.663
R986 B.n829 B.n152 256.663
R987 B.n829 B.n151 256.663
R988 B.n829 B.n150 256.663
R989 B.n829 B.n149 256.663
R990 B.n829 B.n148 256.663
R991 B.n829 B.n147 256.663
R992 B.n829 B.n146 256.663
R993 B.n415 B.n392 256.663
R994 B.n421 B.n392 256.663
R995 B.n423 B.n392 256.663
R996 B.n429 B.n392 256.663
R997 B.n431 B.n392 256.663
R998 B.n437 B.n392 256.663
R999 B.n439 B.n392 256.663
R1000 B.n445 B.n392 256.663
R1001 B.n447 B.n392 256.663
R1002 B.n453 B.n392 256.663
R1003 B.n455 B.n392 256.663
R1004 B.n462 B.n392 256.663
R1005 B.n464 B.n392 256.663
R1006 B.n470 B.n392 256.663
R1007 B.n472 B.n392 256.663
R1008 B.n478 B.n392 256.663
R1009 B.n480 B.n392 256.663
R1010 B.n400 B.t21 223.151
R1011 B.n406 B.t10 223.151
R1012 B.n167 B.t14 223.151
R1013 B.n164 B.t18 223.151
R1014 B.n486 B.n392 176.297
R1015 B.n830 B.n829 176.297
R1016 B.n400 B.t23 163.881
R1017 B.n164 B.t19 163.881
R1018 B.n406 B.t13 163.881
R1019 B.n167 B.t16 163.881
R1020 B.n487 B.n389 163.367
R1021 B.n491 B.n389 163.367
R1022 B.n491 B.n383 163.367
R1023 B.n499 B.n383 163.367
R1024 B.n499 B.n381 163.367
R1025 B.n503 B.n381 163.367
R1026 B.n503 B.n375 163.367
R1027 B.n512 B.n375 163.367
R1028 B.n512 B.n373 163.367
R1029 B.n516 B.n373 163.367
R1030 B.n516 B.n368 163.367
R1031 B.n524 B.n368 163.367
R1032 B.n524 B.n366 163.367
R1033 B.n528 B.n366 163.367
R1034 B.n528 B.n360 163.367
R1035 B.n536 B.n360 163.367
R1036 B.n536 B.n358 163.367
R1037 B.n540 B.n358 163.367
R1038 B.n540 B.n352 163.367
R1039 B.n548 B.n352 163.367
R1040 B.n548 B.n350 163.367
R1041 B.n552 B.n350 163.367
R1042 B.n552 B.n344 163.367
R1043 B.n560 B.n344 163.367
R1044 B.n560 B.n342 163.367
R1045 B.n564 B.n342 163.367
R1046 B.n564 B.n336 163.367
R1047 B.n572 B.n336 163.367
R1048 B.n572 B.n334 163.367
R1049 B.n576 B.n334 163.367
R1050 B.n576 B.n328 163.367
R1051 B.n584 B.n328 163.367
R1052 B.n584 B.n326 163.367
R1053 B.n588 B.n326 163.367
R1054 B.n588 B.n320 163.367
R1055 B.n596 B.n320 163.367
R1056 B.n596 B.n318 163.367
R1057 B.n600 B.n318 163.367
R1058 B.n600 B.n312 163.367
R1059 B.n608 B.n312 163.367
R1060 B.n608 B.n310 163.367
R1061 B.n612 B.n310 163.367
R1062 B.n612 B.n304 163.367
R1063 B.n620 B.n304 163.367
R1064 B.n620 B.n302 163.367
R1065 B.n624 B.n302 163.367
R1066 B.n624 B.n296 163.367
R1067 B.n632 B.n296 163.367
R1068 B.n632 B.n294 163.367
R1069 B.n636 B.n294 163.367
R1070 B.n636 B.n288 163.367
R1071 B.n644 B.n288 163.367
R1072 B.n644 B.n286 163.367
R1073 B.n648 B.n286 163.367
R1074 B.n648 B.n280 163.367
R1075 B.n656 B.n280 163.367
R1076 B.n656 B.n278 163.367
R1077 B.n660 B.n278 163.367
R1078 B.n660 B.n272 163.367
R1079 B.n668 B.n272 163.367
R1080 B.n668 B.n270 163.367
R1081 B.n672 B.n270 163.367
R1082 B.n672 B.n264 163.367
R1083 B.n680 B.n264 163.367
R1084 B.n680 B.n262 163.367
R1085 B.n684 B.n262 163.367
R1086 B.n684 B.n256 163.367
R1087 B.n692 B.n256 163.367
R1088 B.n692 B.n254 163.367
R1089 B.n696 B.n254 163.367
R1090 B.n696 B.n248 163.367
R1091 B.n704 B.n248 163.367
R1092 B.n704 B.n246 163.367
R1093 B.n708 B.n246 163.367
R1094 B.n708 B.n240 163.367
R1095 B.n717 B.n240 163.367
R1096 B.n717 B.n238 163.367
R1097 B.n721 B.n238 163.367
R1098 B.n721 B.n2 163.367
R1099 B.n991 B.n2 163.367
R1100 B.n991 B.n3 163.367
R1101 B.n987 B.n3 163.367
R1102 B.n987 B.n9 163.367
R1103 B.n983 B.n9 163.367
R1104 B.n983 B.n11 163.367
R1105 B.n979 B.n11 163.367
R1106 B.n979 B.n16 163.367
R1107 B.n975 B.n16 163.367
R1108 B.n975 B.n18 163.367
R1109 B.n971 B.n18 163.367
R1110 B.n971 B.n23 163.367
R1111 B.n967 B.n23 163.367
R1112 B.n967 B.n25 163.367
R1113 B.n963 B.n25 163.367
R1114 B.n963 B.n30 163.367
R1115 B.n959 B.n30 163.367
R1116 B.n959 B.n32 163.367
R1117 B.n955 B.n32 163.367
R1118 B.n955 B.n37 163.367
R1119 B.n951 B.n37 163.367
R1120 B.n951 B.n39 163.367
R1121 B.n947 B.n39 163.367
R1122 B.n947 B.n44 163.367
R1123 B.n943 B.n44 163.367
R1124 B.n943 B.n46 163.367
R1125 B.n939 B.n46 163.367
R1126 B.n939 B.n51 163.367
R1127 B.n935 B.n51 163.367
R1128 B.n935 B.n53 163.367
R1129 B.n931 B.n53 163.367
R1130 B.n931 B.n58 163.367
R1131 B.n927 B.n58 163.367
R1132 B.n927 B.n60 163.367
R1133 B.n923 B.n60 163.367
R1134 B.n923 B.n65 163.367
R1135 B.n919 B.n65 163.367
R1136 B.n919 B.n67 163.367
R1137 B.n915 B.n67 163.367
R1138 B.n915 B.n72 163.367
R1139 B.n911 B.n72 163.367
R1140 B.n911 B.n74 163.367
R1141 B.n907 B.n74 163.367
R1142 B.n907 B.n79 163.367
R1143 B.n903 B.n79 163.367
R1144 B.n903 B.n81 163.367
R1145 B.n899 B.n81 163.367
R1146 B.n899 B.n86 163.367
R1147 B.n895 B.n86 163.367
R1148 B.n895 B.n88 163.367
R1149 B.n891 B.n88 163.367
R1150 B.n891 B.n93 163.367
R1151 B.n887 B.n93 163.367
R1152 B.n887 B.n95 163.367
R1153 B.n883 B.n95 163.367
R1154 B.n883 B.n100 163.367
R1155 B.n879 B.n100 163.367
R1156 B.n879 B.n102 163.367
R1157 B.n875 B.n102 163.367
R1158 B.n875 B.n107 163.367
R1159 B.n871 B.n107 163.367
R1160 B.n871 B.n109 163.367
R1161 B.n867 B.n109 163.367
R1162 B.n867 B.n114 163.367
R1163 B.n863 B.n114 163.367
R1164 B.n863 B.n116 163.367
R1165 B.n859 B.n116 163.367
R1166 B.n859 B.n121 163.367
R1167 B.n855 B.n121 163.367
R1168 B.n855 B.n123 163.367
R1169 B.n851 B.n123 163.367
R1170 B.n851 B.n127 163.367
R1171 B.n847 B.n127 163.367
R1172 B.n847 B.n129 163.367
R1173 B.n843 B.n129 163.367
R1174 B.n843 B.n135 163.367
R1175 B.n839 B.n135 163.367
R1176 B.n839 B.n137 163.367
R1177 B.n835 B.n137 163.367
R1178 B.n835 B.n142 163.367
R1179 B.n831 B.n142 163.367
R1180 B.n416 B.n414 163.367
R1181 B.n420 B.n414 163.367
R1182 B.n424 B.n422 163.367
R1183 B.n428 B.n412 163.367
R1184 B.n432 B.n430 163.367
R1185 B.n436 B.n410 163.367
R1186 B.n440 B.n438 163.367
R1187 B.n444 B.n405 163.367
R1188 B.n448 B.n446 163.367
R1189 B.n452 B.n403 163.367
R1190 B.n456 B.n454 163.367
R1191 B.n461 B.n399 163.367
R1192 B.n465 B.n463 163.367
R1193 B.n469 B.n397 163.367
R1194 B.n473 B.n471 163.367
R1195 B.n477 B.n395 163.367
R1196 B.n481 B.n479 163.367
R1197 B.n485 B.n387 163.367
R1198 B.n493 B.n387 163.367
R1199 B.n493 B.n385 163.367
R1200 B.n497 B.n385 163.367
R1201 B.n497 B.n379 163.367
R1202 B.n505 B.n379 163.367
R1203 B.n505 B.n377 163.367
R1204 B.n509 B.n377 163.367
R1205 B.n509 B.n372 163.367
R1206 B.n518 B.n372 163.367
R1207 B.n518 B.n370 163.367
R1208 B.n522 B.n370 163.367
R1209 B.n522 B.n364 163.367
R1210 B.n530 B.n364 163.367
R1211 B.n530 B.n362 163.367
R1212 B.n534 B.n362 163.367
R1213 B.n534 B.n356 163.367
R1214 B.n542 B.n356 163.367
R1215 B.n542 B.n354 163.367
R1216 B.n546 B.n354 163.367
R1217 B.n546 B.n348 163.367
R1218 B.n554 B.n348 163.367
R1219 B.n554 B.n346 163.367
R1220 B.n558 B.n346 163.367
R1221 B.n558 B.n340 163.367
R1222 B.n566 B.n340 163.367
R1223 B.n566 B.n338 163.367
R1224 B.n570 B.n338 163.367
R1225 B.n570 B.n332 163.367
R1226 B.n578 B.n332 163.367
R1227 B.n578 B.n330 163.367
R1228 B.n582 B.n330 163.367
R1229 B.n582 B.n324 163.367
R1230 B.n590 B.n324 163.367
R1231 B.n590 B.n322 163.367
R1232 B.n594 B.n322 163.367
R1233 B.n594 B.n316 163.367
R1234 B.n602 B.n316 163.367
R1235 B.n602 B.n314 163.367
R1236 B.n606 B.n314 163.367
R1237 B.n606 B.n308 163.367
R1238 B.n614 B.n308 163.367
R1239 B.n614 B.n306 163.367
R1240 B.n618 B.n306 163.367
R1241 B.n618 B.n300 163.367
R1242 B.n626 B.n300 163.367
R1243 B.n626 B.n298 163.367
R1244 B.n630 B.n298 163.367
R1245 B.n630 B.n292 163.367
R1246 B.n638 B.n292 163.367
R1247 B.n638 B.n290 163.367
R1248 B.n642 B.n290 163.367
R1249 B.n642 B.n284 163.367
R1250 B.n650 B.n284 163.367
R1251 B.n650 B.n282 163.367
R1252 B.n654 B.n282 163.367
R1253 B.n654 B.n276 163.367
R1254 B.n662 B.n276 163.367
R1255 B.n662 B.n274 163.367
R1256 B.n666 B.n274 163.367
R1257 B.n666 B.n268 163.367
R1258 B.n674 B.n268 163.367
R1259 B.n674 B.n266 163.367
R1260 B.n678 B.n266 163.367
R1261 B.n678 B.n260 163.367
R1262 B.n686 B.n260 163.367
R1263 B.n686 B.n258 163.367
R1264 B.n690 B.n258 163.367
R1265 B.n690 B.n252 163.367
R1266 B.n698 B.n252 163.367
R1267 B.n698 B.n250 163.367
R1268 B.n702 B.n250 163.367
R1269 B.n702 B.n244 163.367
R1270 B.n710 B.n244 163.367
R1271 B.n710 B.n242 163.367
R1272 B.n715 B.n242 163.367
R1273 B.n715 B.n236 163.367
R1274 B.n723 B.n236 163.367
R1275 B.n724 B.n723 163.367
R1276 B.n724 B.n5 163.367
R1277 B.n6 B.n5 163.367
R1278 B.n7 B.n6 163.367
R1279 B.n729 B.n7 163.367
R1280 B.n729 B.n12 163.367
R1281 B.n13 B.n12 163.367
R1282 B.n14 B.n13 163.367
R1283 B.n734 B.n14 163.367
R1284 B.n734 B.n19 163.367
R1285 B.n20 B.n19 163.367
R1286 B.n21 B.n20 163.367
R1287 B.n739 B.n21 163.367
R1288 B.n739 B.n26 163.367
R1289 B.n27 B.n26 163.367
R1290 B.n28 B.n27 163.367
R1291 B.n744 B.n28 163.367
R1292 B.n744 B.n33 163.367
R1293 B.n34 B.n33 163.367
R1294 B.n35 B.n34 163.367
R1295 B.n749 B.n35 163.367
R1296 B.n749 B.n40 163.367
R1297 B.n41 B.n40 163.367
R1298 B.n42 B.n41 163.367
R1299 B.n754 B.n42 163.367
R1300 B.n754 B.n47 163.367
R1301 B.n48 B.n47 163.367
R1302 B.n49 B.n48 163.367
R1303 B.n759 B.n49 163.367
R1304 B.n759 B.n54 163.367
R1305 B.n55 B.n54 163.367
R1306 B.n56 B.n55 163.367
R1307 B.n764 B.n56 163.367
R1308 B.n764 B.n61 163.367
R1309 B.n62 B.n61 163.367
R1310 B.n63 B.n62 163.367
R1311 B.n769 B.n63 163.367
R1312 B.n769 B.n68 163.367
R1313 B.n69 B.n68 163.367
R1314 B.n70 B.n69 163.367
R1315 B.n774 B.n70 163.367
R1316 B.n774 B.n75 163.367
R1317 B.n76 B.n75 163.367
R1318 B.n77 B.n76 163.367
R1319 B.n779 B.n77 163.367
R1320 B.n779 B.n82 163.367
R1321 B.n83 B.n82 163.367
R1322 B.n84 B.n83 163.367
R1323 B.n784 B.n84 163.367
R1324 B.n784 B.n89 163.367
R1325 B.n90 B.n89 163.367
R1326 B.n91 B.n90 163.367
R1327 B.n789 B.n91 163.367
R1328 B.n789 B.n96 163.367
R1329 B.n97 B.n96 163.367
R1330 B.n98 B.n97 163.367
R1331 B.n794 B.n98 163.367
R1332 B.n794 B.n103 163.367
R1333 B.n104 B.n103 163.367
R1334 B.n105 B.n104 163.367
R1335 B.n799 B.n105 163.367
R1336 B.n799 B.n110 163.367
R1337 B.n111 B.n110 163.367
R1338 B.n112 B.n111 163.367
R1339 B.n804 B.n112 163.367
R1340 B.n804 B.n117 163.367
R1341 B.n118 B.n117 163.367
R1342 B.n119 B.n118 163.367
R1343 B.n809 B.n119 163.367
R1344 B.n809 B.n124 163.367
R1345 B.n125 B.n124 163.367
R1346 B.n126 B.n125 163.367
R1347 B.n814 B.n126 163.367
R1348 B.n814 B.n131 163.367
R1349 B.n132 B.n131 163.367
R1350 B.n133 B.n132 163.367
R1351 B.n819 B.n133 163.367
R1352 B.n819 B.n138 163.367
R1353 B.n139 B.n138 163.367
R1354 B.n140 B.n139 163.367
R1355 B.n824 B.n140 163.367
R1356 B.n824 B.n145 163.367
R1357 B.n171 B.n170 163.367
R1358 B.n175 B.n174 163.367
R1359 B.n179 B.n178 163.367
R1360 B.n183 B.n182 163.367
R1361 B.n187 B.n186 163.367
R1362 B.n191 B.n190 163.367
R1363 B.n196 B.n195 163.367
R1364 B.n200 B.n199 163.367
R1365 B.n204 B.n203 163.367
R1366 B.n208 B.n207 163.367
R1367 B.n212 B.n211 163.367
R1368 B.n216 B.n215 163.367
R1369 B.n220 B.n219 163.367
R1370 B.n224 B.n223 163.367
R1371 B.n228 B.n227 163.367
R1372 B.n232 B.n231 163.367
R1373 B.n828 B.n163 163.367
R1374 B.n486 B.n388 100.742
R1375 B.n492 B.n388 100.742
R1376 B.n492 B.n384 100.742
R1377 B.n498 B.n384 100.742
R1378 B.n498 B.n380 100.742
R1379 B.n504 B.n380 100.742
R1380 B.n504 B.n376 100.742
R1381 B.n511 B.n376 100.742
R1382 B.n511 B.n510 100.742
R1383 B.n517 B.n369 100.742
R1384 B.n523 B.n369 100.742
R1385 B.n523 B.n365 100.742
R1386 B.n529 B.n365 100.742
R1387 B.n529 B.n361 100.742
R1388 B.n535 B.n361 100.742
R1389 B.n535 B.n357 100.742
R1390 B.n541 B.n357 100.742
R1391 B.n541 B.n353 100.742
R1392 B.n547 B.n353 100.742
R1393 B.n547 B.n349 100.742
R1394 B.n553 B.n349 100.742
R1395 B.n553 B.n345 100.742
R1396 B.n559 B.n345 100.742
R1397 B.n565 B.n341 100.742
R1398 B.n565 B.n337 100.742
R1399 B.n571 B.n337 100.742
R1400 B.n571 B.n333 100.742
R1401 B.n577 B.n333 100.742
R1402 B.n577 B.n329 100.742
R1403 B.n583 B.n329 100.742
R1404 B.n583 B.n325 100.742
R1405 B.n589 B.n325 100.742
R1406 B.n589 B.n321 100.742
R1407 B.n595 B.n321 100.742
R1408 B.n601 B.n317 100.742
R1409 B.n601 B.n313 100.742
R1410 B.n607 B.n313 100.742
R1411 B.n607 B.n309 100.742
R1412 B.n613 B.n309 100.742
R1413 B.n613 B.n305 100.742
R1414 B.n619 B.n305 100.742
R1415 B.n619 B.n301 100.742
R1416 B.n625 B.n301 100.742
R1417 B.n625 B.n297 100.742
R1418 B.n631 B.n297 100.742
R1419 B.n637 B.n293 100.742
R1420 B.n637 B.n289 100.742
R1421 B.n643 B.n289 100.742
R1422 B.n643 B.n285 100.742
R1423 B.n649 B.n285 100.742
R1424 B.n649 B.n281 100.742
R1425 B.n655 B.n281 100.742
R1426 B.n655 B.n277 100.742
R1427 B.n661 B.n277 100.742
R1428 B.n661 B.n273 100.742
R1429 B.n667 B.n273 100.742
R1430 B.n673 B.n269 100.742
R1431 B.n673 B.n265 100.742
R1432 B.n679 B.n265 100.742
R1433 B.n679 B.n261 100.742
R1434 B.n685 B.n261 100.742
R1435 B.n685 B.n257 100.742
R1436 B.n691 B.n257 100.742
R1437 B.n691 B.n253 100.742
R1438 B.n697 B.n253 100.742
R1439 B.n697 B.n249 100.742
R1440 B.n703 B.n249 100.742
R1441 B.n709 B.n245 100.742
R1442 B.n709 B.n241 100.742
R1443 B.n716 B.n241 100.742
R1444 B.n716 B.n237 100.742
R1445 B.n722 B.n237 100.742
R1446 B.n722 B.n4 100.742
R1447 B.n990 B.n4 100.742
R1448 B.n990 B.n989 100.742
R1449 B.n989 B.n988 100.742
R1450 B.n988 B.n8 100.742
R1451 B.n982 B.n8 100.742
R1452 B.n982 B.n981 100.742
R1453 B.n981 B.n980 100.742
R1454 B.n980 B.n15 100.742
R1455 B.n974 B.n973 100.742
R1456 B.n973 B.n972 100.742
R1457 B.n972 B.n22 100.742
R1458 B.n966 B.n22 100.742
R1459 B.n966 B.n965 100.742
R1460 B.n965 B.n964 100.742
R1461 B.n964 B.n29 100.742
R1462 B.n958 B.n29 100.742
R1463 B.n958 B.n957 100.742
R1464 B.n957 B.n956 100.742
R1465 B.n956 B.n36 100.742
R1466 B.n950 B.n949 100.742
R1467 B.n949 B.n948 100.742
R1468 B.n948 B.n43 100.742
R1469 B.n942 B.n43 100.742
R1470 B.n942 B.n941 100.742
R1471 B.n941 B.n940 100.742
R1472 B.n940 B.n50 100.742
R1473 B.n934 B.n50 100.742
R1474 B.n934 B.n933 100.742
R1475 B.n933 B.n932 100.742
R1476 B.n932 B.n57 100.742
R1477 B.n926 B.n925 100.742
R1478 B.n925 B.n924 100.742
R1479 B.n924 B.n64 100.742
R1480 B.n918 B.n64 100.742
R1481 B.n918 B.n917 100.742
R1482 B.n917 B.n916 100.742
R1483 B.n916 B.n71 100.742
R1484 B.n910 B.n71 100.742
R1485 B.n910 B.n909 100.742
R1486 B.n909 B.n908 100.742
R1487 B.n908 B.n78 100.742
R1488 B.n902 B.n901 100.742
R1489 B.n901 B.n900 100.742
R1490 B.n900 B.n85 100.742
R1491 B.n894 B.n85 100.742
R1492 B.n894 B.n893 100.742
R1493 B.n893 B.n892 100.742
R1494 B.n892 B.n92 100.742
R1495 B.n886 B.n92 100.742
R1496 B.n886 B.n885 100.742
R1497 B.n885 B.n884 100.742
R1498 B.n884 B.n99 100.742
R1499 B.n878 B.n877 100.742
R1500 B.n877 B.n876 100.742
R1501 B.n876 B.n106 100.742
R1502 B.n870 B.n106 100.742
R1503 B.n870 B.n869 100.742
R1504 B.n869 B.n868 100.742
R1505 B.n868 B.n113 100.742
R1506 B.n862 B.n113 100.742
R1507 B.n862 B.n861 100.742
R1508 B.n861 B.n860 100.742
R1509 B.n860 B.n120 100.742
R1510 B.n854 B.n120 100.742
R1511 B.n854 B.n853 100.742
R1512 B.n853 B.n852 100.742
R1513 B.n846 B.n130 100.742
R1514 B.n846 B.n845 100.742
R1515 B.n845 B.n844 100.742
R1516 B.n844 B.n134 100.742
R1517 B.n838 B.n134 100.742
R1518 B.n838 B.n837 100.742
R1519 B.n837 B.n836 100.742
R1520 B.n836 B.n141 100.742
R1521 B.n830 B.n141 100.742
R1522 B.n401 B.t22 84.9474
R1523 B.n165 B.t20 84.9474
R1524 B.n407 B.t12 84.9471
R1525 B.n168 B.t17 84.9471
R1526 B.n401 B.n400 78.9338
R1527 B.n407 B.n406 78.9338
R1528 B.n168 B.n167 78.9338
R1529 B.n165 B.n164 78.9338
R1530 B.n415 B.n391 71.676
R1531 B.n421 B.n420 71.676
R1532 B.n424 B.n423 71.676
R1533 B.n429 B.n428 71.676
R1534 B.n432 B.n431 71.676
R1535 B.n437 B.n436 71.676
R1536 B.n440 B.n439 71.676
R1537 B.n445 B.n444 71.676
R1538 B.n448 B.n447 71.676
R1539 B.n453 B.n452 71.676
R1540 B.n456 B.n455 71.676
R1541 B.n462 B.n461 71.676
R1542 B.n465 B.n464 71.676
R1543 B.n470 B.n469 71.676
R1544 B.n473 B.n472 71.676
R1545 B.n478 B.n477 71.676
R1546 B.n481 B.n480 71.676
R1547 B.n146 B.n144 71.676
R1548 B.n171 B.n147 71.676
R1549 B.n175 B.n148 71.676
R1550 B.n179 B.n149 71.676
R1551 B.n183 B.n150 71.676
R1552 B.n187 B.n151 71.676
R1553 B.n191 B.n152 71.676
R1554 B.n196 B.n153 71.676
R1555 B.n200 B.n154 71.676
R1556 B.n204 B.n155 71.676
R1557 B.n208 B.n156 71.676
R1558 B.n212 B.n157 71.676
R1559 B.n216 B.n158 71.676
R1560 B.n220 B.n159 71.676
R1561 B.n224 B.n160 71.676
R1562 B.n228 B.n161 71.676
R1563 B.n232 B.n162 71.676
R1564 B.n163 B.n162 71.676
R1565 B.n231 B.n161 71.676
R1566 B.n227 B.n160 71.676
R1567 B.n223 B.n159 71.676
R1568 B.n219 B.n158 71.676
R1569 B.n215 B.n157 71.676
R1570 B.n211 B.n156 71.676
R1571 B.n207 B.n155 71.676
R1572 B.n203 B.n154 71.676
R1573 B.n199 B.n153 71.676
R1574 B.n195 B.n152 71.676
R1575 B.n190 B.n151 71.676
R1576 B.n186 B.n150 71.676
R1577 B.n182 B.n149 71.676
R1578 B.n178 B.n148 71.676
R1579 B.n174 B.n147 71.676
R1580 B.n170 B.n146 71.676
R1581 B.n416 B.n415 71.676
R1582 B.n422 B.n421 71.676
R1583 B.n423 B.n412 71.676
R1584 B.n430 B.n429 71.676
R1585 B.n431 B.n410 71.676
R1586 B.n438 B.n437 71.676
R1587 B.n439 B.n405 71.676
R1588 B.n446 B.n445 71.676
R1589 B.n447 B.n403 71.676
R1590 B.n454 B.n453 71.676
R1591 B.n455 B.n399 71.676
R1592 B.n463 B.n462 71.676
R1593 B.n464 B.n397 71.676
R1594 B.n471 B.n470 71.676
R1595 B.n472 B.n395 71.676
R1596 B.n479 B.n478 71.676
R1597 B.n480 B.n393 71.676
R1598 B.n517 B.t11 65.1857
R1599 B.n852 B.t15 65.1857
R1600 B.n458 B.n401 59.5399
R1601 B.n408 B.n407 59.5399
R1602 B.n193 B.n168 59.5399
R1603 B.n166 B.n165 59.5399
R1604 B.t8 B.n245 59.2598
R1605 B.t0 B.n15 59.2598
R1606 B.t3 B.n269 56.2968
R1607 B.t5 B.n36 56.2968
R1608 B.n559 B.t9 53.3338
R1609 B.t6 B.n293 53.3338
R1610 B.t1 B.n57 53.3338
R1611 B.n878 B.t7 53.3338
R1612 B.n595 B.t2 50.3709
R1613 B.t2 B.n317 50.3709
R1614 B.t4 B.n78 50.3709
R1615 B.n902 B.t4 50.3709
R1616 B.t9 B.n341 47.4079
R1617 B.n631 B.t6 47.4079
R1618 B.n926 B.t1 47.4079
R1619 B.t7 B.n99 47.4079
R1620 B.n667 B.t3 44.4449
R1621 B.n950 B.t5 44.4449
R1622 B.n703 B.t8 41.482
R1623 B.n974 B.t0 41.482
R1624 B.n510 B.t11 35.5561
R1625 B.n130 B.t15 35.5561
R1626 B.n832 B.n143 31.0639
R1627 B.n827 B.n826 31.0639
R1628 B.n484 B.n483 31.0639
R1629 B.n488 B.n390 31.0639
R1630 B B.n992 18.0485
R1631 B.n169 B.n143 10.6151
R1632 B.n172 B.n169 10.6151
R1633 B.n173 B.n172 10.6151
R1634 B.n176 B.n173 10.6151
R1635 B.n177 B.n176 10.6151
R1636 B.n180 B.n177 10.6151
R1637 B.n181 B.n180 10.6151
R1638 B.n184 B.n181 10.6151
R1639 B.n185 B.n184 10.6151
R1640 B.n188 B.n185 10.6151
R1641 B.n189 B.n188 10.6151
R1642 B.n192 B.n189 10.6151
R1643 B.n197 B.n194 10.6151
R1644 B.n198 B.n197 10.6151
R1645 B.n201 B.n198 10.6151
R1646 B.n202 B.n201 10.6151
R1647 B.n205 B.n202 10.6151
R1648 B.n206 B.n205 10.6151
R1649 B.n209 B.n206 10.6151
R1650 B.n210 B.n209 10.6151
R1651 B.n214 B.n213 10.6151
R1652 B.n217 B.n214 10.6151
R1653 B.n218 B.n217 10.6151
R1654 B.n221 B.n218 10.6151
R1655 B.n222 B.n221 10.6151
R1656 B.n225 B.n222 10.6151
R1657 B.n226 B.n225 10.6151
R1658 B.n229 B.n226 10.6151
R1659 B.n230 B.n229 10.6151
R1660 B.n233 B.n230 10.6151
R1661 B.n234 B.n233 10.6151
R1662 B.n827 B.n234 10.6151
R1663 B.n484 B.n386 10.6151
R1664 B.n494 B.n386 10.6151
R1665 B.n495 B.n494 10.6151
R1666 B.n496 B.n495 10.6151
R1667 B.n496 B.n378 10.6151
R1668 B.n506 B.n378 10.6151
R1669 B.n507 B.n506 10.6151
R1670 B.n508 B.n507 10.6151
R1671 B.n508 B.n371 10.6151
R1672 B.n519 B.n371 10.6151
R1673 B.n520 B.n519 10.6151
R1674 B.n521 B.n520 10.6151
R1675 B.n521 B.n363 10.6151
R1676 B.n531 B.n363 10.6151
R1677 B.n532 B.n531 10.6151
R1678 B.n533 B.n532 10.6151
R1679 B.n533 B.n355 10.6151
R1680 B.n543 B.n355 10.6151
R1681 B.n544 B.n543 10.6151
R1682 B.n545 B.n544 10.6151
R1683 B.n545 B.n347 10.6151
R1684 B.n555 B.n347 10.6151
R1685 B.n556 B.n555 10.6151
R1686 B.n557 B.n556 10.6151
R1687 B.n557 B.n339 10.6151
R1688 B.n567 B.n339 10.6151
R1689 B.n568 B.n567 10.6151
R1690 B.n569 B.n568 10.6151
R1691 B.n569 B.n331 10.6151
R1692 B.n579 B.n331 10.6151
R1693 B.n580 B.n579 10.6151
R1694 B.n581 B.n580 10.6151
R1695 B.n581 B.n323 10.6151
R1696 B.n591 B.n323 10.6151
R1697 B.n592 B.n591 10.6151
R1698 B.n593 B.n592 10.6151
R1699 B.n593 B.n315 10.6151
R1700 B.n603 B.n315 10.6151
R1701 B.n604 B.n603 10.6151
R1702 B.n605 B.n604 10.6151
R1703 B.n605 B.n307 10.6151
R1704 B.n615 B.n307 10.6151
R1705 B.n616 B.n615 10.6151
R1706 B.n617 B.n616 10.6151
R1707 B.n617 B.n299 10.6151
R1708 B.n627 B.n299 10.6151
R1709 B.n628 B.n627 10.6151
R1710 B.n629 B.n628 10.6151
R1711 B.n629 B.n291 10.6151
R1712 B.n639 B.n291 10.6151
R1713 B.n640 B.n639 10.6151
R1714 B.n641 B.n640 10.6151
R1715 B.n641 B.n283 10.6151
R1716 B.n651 B.n283 10.6151
R1717 B.n652 B.n651 10.6151
R1718 B.n653 B.n652 10.6151
R1719 B.n653 B.n275 10.6151
R1720 B.n663 B.n275 10.6151
R1721 B.n664 B.n663 10.6151
R1722 B.n665 B.n664 10.6151
R1723 B.n665 B.n267 10.6151
R1724 B.n675 B.n267 10.6151
R1725 B.n676 B.n675 10.6151
R1726 B.n677 B.n676 10.6151
R1727 B.n677 B.n259 10.6151
R1728 B.n687 B.n259 10.6151
R1729 B.n688 B.n687 10.6151
R1730 B.n689 B.n688 10.6151
R1731 B.n689 B.n251 10.6151
R1732 B.n699 B.n251 10.6151
R1733 B.n700 B.n699 10.6151
R1734 B.n701 B.n700 10.6151
R1735 B.n701 B.n243 10.6151
R1736 B.n711 B.n243 10.6151
R1737 B.n712 B.n711 10.6151
R1738 B.n714 B.n712 10.6151
R1739 B.n714 B.n713 10.6151
R1740 B.n713 B.n235 10.6151
R1741 B.n725 B.n235 10.6151
R1742 B.n726 B.n725 10.6151
R1743 B.n727 B.n726 10.6151
R1744 B.n728 B.n727 10.6151
R1745 B.n730 B.n728 10.6151
R1746 B.n731 B.n730 10.6151
R1747 B.n732 B.n731 10.6151
R1748 B.n733 B.n732 10.6151
R1749 B.n735 B.n733 10.6151
R1750 B.n736 B.n735 10.6151
R1751 B.n737 B.n736 10.6151
R1752 B.n738 B.n737 10.6151
R1753 B.n740 B.n738 10.6151
R1754 B.n741 B.n740 10.6151
R1755 B.n742 B.n741 10.6151
R1756 B.n743 B.n742 10.6151
R1757 B.n745 B.n743 10.6151
R1758 B.n746 B.n745 10.6151
R1759 B.n747 B.n746 10.6151
R1760 B.n748 B.n747 10.6151
R1761 B.n750 B.n748 10.6151
R1762 B.n751 B.n750 10.6151
R1763 B.n752 B.n751 10.6151
R1764 B.n753 B.n752 10.6151
R1765 B.n755 B.n753 10.6151
R1766 B.n756 B.n755 10.6151
R1767 B.n757 B.n756 10.6151
R1768 B.n758 B.n757 10.6151
R1769 B.n760 B.n758 10.6151
R1770 B.n761 B.n760 10.6151
R1771 B.n762 B.n761 10.6151
R1772 B.n763 B.n762 10.6151
R1773 B.n765 B.n763 10.6151
R1774 B.n766 B.n765 10.6151
R1775 B.n767 B.n766 10.6151
R1776 B.n768 B.n767 10.6151
R1777 B.n770 B.n768 10.6151
R1778 B.n771 B.n770 10.6151
R1779 B.n772 B.n771 10.6151
R1780 B.n773 B.n772 10.6151
R1781 B.n775 B.n773 10.6151
R1782 B.n776 B.n775 10.6151
R1783 B.n777 B.n776 10.6151
R1784 B.n778 B.n777 10.6151
R1785 B.n780 B.n778 10.6151
R1786 B.n781 B.n780 10.6151
R1787 B.n782 B.n781 10.6151
R1788 B.n783 B.n782 10.6151
R1789 B.n785 B.n783 10.6151
R1790 B.n786 B.n785 10.6151
R1791 B.n787 B.n786 10.6151
R1792 B.n788 B.n787 10.6151
R1793 B.n790 B.n788 10.6151
R1794 B.n791 B.n790 10.6151
R1795 B.n792 B.n791 10.6151
R1796 B.n793 B.n792 10.6151
R1797 B.n795 B.n793 10.6151
R1798 B.n796 B.n795 10.6151
R1799 B.n797 B.n796 10.6151
R1800 B.n798 B.n797 10.6151
R1801 B.n800 B.n798 10.6151
R1802 B.n801 B.n800 10.6151
R1803 B.n802 B.n801 10.6151
R1804 B.n803 B.n802 10.6151
R1805 B.n805 B.n803 10.6151
R1806 B.n806 B.n805 10.6151
R1807 B.n807 B.n806 10.6151
R1808 B.n808 B.n807 10.6151
R1809 B.n810 B.n808 10.6151
R1810 B.n811 B.n810 10.6151
R1811 B.n812 B.n811 10.6151
R1812 B.n813 B.n812 10.6151
R1813 B.n815 B.n813 10.6151
R1814 B.n816 B.n815 10.6151
R1815 B.n817 B.n816 10.6151
R1816 B.n818 B.n817 10.6151
R1817 B.n820 B.n818 10.6151
R1818 B.n821 B.n820 10.6151
R1819 B.n822 B.n821 10.6151
R1820 B.n823 B.n822 10.6151
R1821 B.n825 B.n823 10.6151
R1822 B.n826 B.n825 10.6151
R1823 B.n417 B.n390 10.6151
R1824 B.n418 B.n417 10.6151
R1825 B.n419 B.n418 10.6151
R1826 B.n419 B.n413 10.6151
R1827 B.n425 B.n413 10.6151
R1828 B.n426 B.n425 10.6151
R1829 B.n427 B.n426 10.6151
R1830 B.n427 B.n411 10.6151
R1831 B.n433 B.n411 10.6151
R1832 B.n434 B.n433 10.6151
R1833 B.n435 B.n434 10.6151
R1834 B.n435 B.n409 10.6151
R1835 B.n442 B.n441 10.6151
R1836 B.n443 B.n442 10.6151
R1837 B.n443 B.n404 10.6151
R1838 B.n449 B.n404 10.6151
R1839 B.n450 B.n449 10.6151
R1840 B.n451 B.n450 10.6151
R1841 B.n451 B.n402 10.6151
R1842 B.n457 B.n402 10.6151
R1843 B.n460 B.n459 10.6151
R1844 B.n460 B.n398 10.6151
R1845 B.n466 B.n398 10.6151
R1846 B.n467 B.n466 10.6151
R1847 B.n468 B.n467 10.6151
R1848 B.n468 B.n396 10.6151
R1849 B.n474 B.n396 10.6151
R1850 B.n475 B.n474 10.6151
R1851 B.n476 B.n475 10.6151
R1852 B.n476 B.n394 10.6151
R1853 B.n482 B.n394 10.6151
R1854 B.n483 B.n482 10.6151
R1855 B.n489 B.n488 10.6151
R1856 B.n490 B.n489 10.6151
R1857 B.n490 B.n382 10.6151
R1858 B.n500 B.n382 10.6151
R1859 B.n501 B.n500 10.6151
R1860 B.n502 B.n501 10.6151
R1861 B.n502 B.n374 10.6151
R1862 B.n513 B.n374 10.6151
R1863 B.n514 B.n513 10.6151
R1864 B.n515 B.n514 10.6151
R1865 B.n515 B.n367 10.6151
R1866 B.n525 B.n367 10.6151
R1867 B.n526 B.n525 10.6151
R1868 B.n527 B.n526 10.6151
R1869 B.n527 B.n359 10.6151
R1870 B.n537 B.n359 10.6151
R1871 B.n538 B.n537 10.6151
R1872 B.n539 B.n538 10.6151
R1873 B.n539 B.n351 10.6151
R1874 B.n549 B.n351 10.6151
R1875 B.n550 B.n549 10.6151
R1876 B.n551 B.n550 10.6151
R1877 B.n551 B.n343 10.6151
R1878 B.n561 B.n343 10.6151
R1879 B.n562 B.n561 10.6151
R1880 B.n563 B.n562 10.6151
R1881 B.n563 B.n335 10.6151
R1882 B.n573 B.n335 10.6151
R1883 B.n574 B.n573 10.6151
R1884 B.n575 B.n574 10.6151
R1885 B.n575 B.n327 10.6151
R1886 B.n585 B.n327 10.6151
R1887 B.n586 B.n585 10.6151
R1888 B.n587 B.n586 10.6151
R1889 B.n587 B.n319 10.6151
R1890 B.n597 B.n319 10.6151
R1891 B.n598 B.n597 10.6151
R1892 B.n599 B.n598 10.6151
R1893 B.n599 B.n311 10.6151
R1894 B.n609 B.n311 10.6151
R1895 B.n610 B.n609 10.6151
R1896 B.n611 B.n610 10.6151
R1897 B.n611 B.n303 10.6151
R1898 B.n621 B.n303 10.6151
R1899 B.n622 B.n621 10.6151
R1900 B.n623 B.n622 10.6151
R1901 B.n623 B.n295 10.6151
R1902 B.n633 B.n295 10.6151
R1903 B.n634 B.n633 10.6151
R1904 B.n635 B.n634 10.6151
R1905 B.n635 B.n287 10.6151
R1906 B.n645 B.n287 10.6151
R1907 B.n646 B.n645 10.6151
R1908 B.n647 B.n646 10.6151
R1909 B.n647 B.n279 10.6151
R1910 B.n657 B.n279 10.6151
R1911 B.n658 B.n657 10.6151
R1912 B.n659 B.n658 10.6151
R1913 B.n659 B.n271 10.6151
R1914 B.n669 B.n271 10.6151
R1915 B.n670 B.n669 10.6151
R1916 B.n671 B.n670 10.6151
R1917 B.n671 B.n263 10.6151
R1918 B.n681 B.n263 10.6151
R1919 B.n682 B.n681 10.6151
R1920 B.n683 B.n682 10.6151
R1921 B.n683 B.n255 10.6151
R1922 B.n693 B.n255 10.6151
R1923 B.n694 B.n693 10.6151
R1924 B.n695 B.n694 10.6151
R1925 B.n695 B.n247 10.6151
R1926 B.n705 B.n247 10.6151
R1927 B.n706 B.n705 10.6151
R1928 B.n707 B.n706 10.6151
R1929 B.n707 B.n239 10.6151
R1930 B.n718 B.n239 10.6151
R1931 B.n719 B.n718 10.6151
R1932 B.n720 B.n719 10.6151
R1933 B.n720 B.n0 10.6151
R1934 B.n986 B.n1 10.6151
R1935 B.n986 B.n985 10.6151
R1936 B.n985 B.n984 10.6151
R1937 B.n984 B.n10 10.6151
R1938 B.n978 B.n10 10.6151
R1939 B.n978 B.n977 10.6151
R1940 B.n977 B.n976 10.6151
R1941 B.n976 B.n17 10.6151
R1942 B.n970 B.n17 10.6151
R1943 B.n970 B.n969 10.6151
R1944 B.n969 B.n968 10.6151
R1945 B.n968 B.n24 10.6151
R1946 B.n962 B.n24 10.6151
R1947 B.n962 B.n961 10.6151
R1948 B.n961 B.n960 10.6151
R1949 B.n960 B.n31 10.6151
R1950 B.n954 B.n31 10.6151
R1951 B.n954 B.n953 10.6151
R1952 B.n953 B.n952 10.6151
R1953 B.n952 B.n38 10.6151
R1954 B.n946 B.n38 10.6151
R1955 B.n946 B.n945 10.6151
R1956 B.n945 B.n944 10.6151
R1957 B.n944 B.n45 10.6151
R1958 B.n938 B.n45 10.6151
R1959 B.n938 B.n937 10.6151
R1960 B.n937 B.n936 10.6151
R1961 B.n936 B.n52 10.6151
R1962 B.n930 B.n52 10.6151
R1963 B.n930 B.n929 10.6151
R1964 B.n929 B.n928 10.6151
R1965 B.n928 B.n59 10.6151
R1966 B.n922 B.n59 10.6151
R1967 B.n922 B.n921 10.6151
R1968 B.n921 B.n920 10.6151
R1969 B.n920 B.n66 10.6151
R1970 B.n914 B.n66 10.6151
R1971 B.n914 B.n913 10.6151
R1972 B.n913 B.n912 10.6151
R1973 B.n912 B.n73 10.6151
R1974 B.n906 B.n73 10.6151
R1975 B.n906 B.n905 10.6151
R1976 B.n905 B.n904 10.6151
R1977 B.n904 B.n80 10.6151
R1978 B.n898 B.n80 10.6151
R1979 B.n898 B.n897 10.6151
R1980 B.n897 B.n896 10.6151
R1981 B.n896 B.n87 10.6151
R1982 B.n890 B.n87 10.6151
R1983 B.n890 B.n889 10.6151
R1984 B.n889 B.n888 10.6151
R1985 B.n888 B.n94 10.6151
R1986 B.n882 B.n94 10.6151
R1987 B.n882 B.n881 10.6151
R1988 B.n881 B.n880 10.6151
R1989 B.n880 B.n101 10.6151
R1990 B.n874 B.n101 10.6151
R1991 B.n874 B.n873 10.6151
R1992 B.n873 B.n872 10.6151
R1993 B.n872 B.n108 10.6151
R1994 B.n866 B.n108 10.6151
R1995 B.n866 B.n865 10.6151
R1996 B.n865 B.n864 10.6151
R1997 B.n864 B.n115 10.6151
R1998 B.n858 B.n115 10.6151
R1999 B.n858 B.n857 10.6151
R2000 B.n857 B.n856 10.6151
R2001 B.n856 B.n122 10.6151
R2002 B.n850 B.n122 10.6151
R2003 B.n850 B.n849 10.6151
R2004 B.n849 B.n848 10.6151
R2005 B.n848 B.n128 10.6151
R2006 B.n842 B.n128 10.6151
R2007 B.n842 B.n841 10.6151
R2008 B.n841 B.n840 10.6151
R2009 B.n840 B.n136 10.6151
R2010 B.n834 B.n136 10.6151
R2011 B.n834 B.n833 10.6151
R2012 B.n833 B.n832 10.6151
R2013 B.n194 B.n193 6.5566
R2014 B.n210 B.n166 6.5566
R2015 B.n441 B.n408 6.5566
R2016 B.n458 B.n457 6.5566
R2017 B.n193 B.n192 4.05904
R2018 B.n213 B.n166 4.05904
R2019 B.n409 B.n408 4.05904
R2020 B.n459 B.n458 4.05904
R2021 B.n992 B.n0 2.81026
R2022 B.n992 B.n1 2.81026
R2023 VN.n108 VN.n107 161.3
R2024 VN.n106 VN.n56 161.3
R2025 VN.n105 VN.n104 161.3
R2026 VN.n103 VN.n57 161.3
R2027 VN.n102 VN.n101 161.3
R2028 VN.n100 VN.n58 161.3
R2029 VN.n99 VN.n98 161.3
R2030 VN.n97 VN.n59 161.3
R2031 VN.n96 VN.n95 161.3
R2032 VN.n94 VN.n60 161.3
R2033 VN.n93 VN.n92 161.3
R2034 VN.n91 VN.n62 161.3
R2035 VN.n90 VN.n89 161.3
R2036 VN.n88 VN.n63 161.3
R2037 VN.n87 VN.n86 161.3
R2038 VN.n85 VN.n64 161.3
R2039 VN.n84 VN.n83 161.3
R2040 VN.n82 VN.n65 161.3
R2041 VN.n81 VN.n80 161.3
R2042 VN.n79 VN.n66 161.3
R2043 VN.n78 VN.n77 161.3
R2044 VN.n76 VN.n67 161.3
R2045 VN.n75 VN.n74 161.3
R2046 VN.n73 VN.n68 161.3
R2047 VN.n72 VN.n71 161.3
R2048 VN.n53 VN.n52 161.3
R2049 VN.n51 VN.n1 161.3
R2050 VN.n50 VN.n49 161.3
R2051 VN.n48 VN.n2 161.3
R2052 VN.n47 VN.n46 161.3
R2053 VN.n45 VN.n3 161.3
R2054 VN.n44 VN.n43 161.3
R2055 VN.n42 VN.n4 161.3
R2056 VN.n41 VN.n40 161.3
R2057 VN.n38 VN.n5 161.3
R2058 VN.n37 VN.n36 161.3
R2059 VN.n35 VN.n6 161.3
R2060 VN.n34 VN.n33 161.3
R2061 VN.n32 VN.n7 161.3
R2062 VN.n31 VN.n30 161.3
R2063 VN.n29 VN.n8 161.3
R2064 VN.n28 VN.n27 161.3
R2065 VN.n26 VN.n9 161.3
R2066 VN.n25 VN.n24 161.3
R2067 VN.n23 VN.n10 161.3
R2068 VN.n22 VN.n21 161.3
R2069 VN.n20 VN.n11 161.3
R2070 VN.n19 VN.n18 161.3
R2071 VN.n17 VN.n12 161.3
R2072 VN.n16 VN.n15 161.3
R2073 VN.n54 VN.n0 83.2166
R2074 VN.n109 VN.n55 83.2166
R2075 VN.n14 VN.n13 71.3788
R2076 VN.n70 VN.n69 71.3788
R2077 VN VN.n109 52.1154
R2078 VN.n46 VN.n2 50.6917
R2079 VN.n101 VN.n57 50.6917
R2080 VN.n13 VN.t9 46.6601
R2081 VN.n69 VN.t4 46.6601
R2082 VN.n21 VN.n20 43.8928
R2083 VN.n33 VN.n6 43.8928
R2084 VN.n77 VN.n76 43.8928
R2085 VN.n89 VN.n62 43.8928
R2086 VN.n21 VN.n10 37.094
R2087 VN.n33 VN.n32 37.094
R2088 VN.n77 VN.n66 37.094
R2089 VN.n89 VN.n88 37.094
R2090 VN.n46 VN.n45 30.2951
R2091 VN.n101 VN.n100 30.2951
R2092 VN.n15 VN.n12 24.4675
R2093 VN.n19 VN.n12 24.4675
R2094 VN.n20 VN.n19 24.4675
R2095 VN.n25 VN.n10 24.4675
R2096 VN.n26 VN.n25 24.4675
R2097 VN.n27 VN.n26 24.4675
R2098 VN.n27 VN.n8 24.4675
R2099 VN.n31 VN.n8 24.4675
R2100 VN.n32 VN.n31 24.4675
R2101 VN.n37 VN.n6 24.4675
R2102 VN.n38 VN.n37 24.4675
R2103 VN.n40 VN.n38 24.4675
R2104 VN.n44 VN.n4 24.4675
R2105 VN.n45 VN.n44 24.4675
R2106 VN.n50 VN.n2 24.4675
R2107 VN.n51 VN.n50 24.4675
R2108 VN.n52 VN.n51 24.4675
R2109 VN.n76 VN.n75 24.4675
R2110 VN.n75 VN.n68 24.4675
R2111 VN.n71 VN.n68 24.4675
R2112 VN.n88 VN.n87 24.4675
R2113 VN.n87 VN.n64 24.4675
R2114 VN.n83 VN.n64 24.4675
R2115 VN.n83 VN.n82 24.4675
R2116 VN.n82 VN.n81 24.4675
R2117 VN.n81 VN.n66 24.4675
R2118 VN.n100 VN.n99 24.4675
R2119 VN.n99 VN.n59 24.4675
R2120 VN.n95 VN.n94 24.4675
R2121 VN.n94 VN.n93 24.4675
R2122 VN.n93 VN.n62 24.4675
R2123 VN.n107 VN.n106 24.4675
R2124 VN.n106 VN.n105 24.4675
R2125 VN.n105 VN.n57 24.4675
R2126 VN.n39 VN.n4 21.0421
R2127 VN.n61 VN.n59 21.0421
R2128 VN.n27 VN.t8 13.8548
R2129 VN.n14 VN.t6 13.8548
R2130 VN.n39 VN.t0 13.8548
R2131 VN.n0 VN.t1 13.8548
R2132 VN.n83 VN.t7 13.8548
R2133 VN.n70 VN.t5 13.8548
R2134 VN.n61 VN.t3 13.8548
R2135 VN.n55 VN.t2 13.8548
R2136 VN.n52 VN.n0 6.85126
R2137 VN.n107 VN.n55 6.85126
R2138 VN.n15 VN.n14 3.42588
R2139 VN.n40 VN.n39 3.42588
R2140 VN.n71 VN.n70 3.42588
R2141 VN.n95 VN.n61 3.42588
R2142 VN.n16 VN.n13 3.25233
R2143 VN.n72 VN.n69 3.25233
R2144 VN.n109 VN.n108 0.354971
R2145 VN.n54 VN.n53 0.354971
R2146 VN VN.n54 0.26696
R2147 VN.n108 VN.n56 0.189894
R2148 VN.n104 VN.n56 0.189894
R2149 VN.n104 VN.n103 0.189894
R2150 VN.n103 VN.n102 0.189894
R2151 VN.n102 VN.n58 0.189894
R2152 VN.n98 VN.n58 0.189894
R2153 VN.n98 VN.n97 0.189894
R2154 VN.n97 VN.n96 0.189894
R2155 VN.n96 VN.n60 0.189894
R2156 VN.n92 VN.n60 0.189894
R2157 VN.n92 VN.n91 0.189894
R2158 VN.n91 VN.n90 0.189894
R2159 VN.n90 VN.n63 0.189894
R2160 VN.n86 VN.n63 0.189894
R2161 VN.n86 VN.n85 0.189894
R2162 VN.n85 VN.n84 0.189894
R2163 VN.n84 VN.n65 0.189894
R2164 VN.n80 VN.n65 0.189894
R2165 VN.n80 VN.n79 0.189894
R2166 VN.n79 VN.n78 0.189894
R2167 VN.n78 VN.n67 0.189894
R2168 VN.n74 VN.n67 0.189894
R2169 VN.n74 VN.n73 0.189894
R2170 VN.n73 VN.n72 0.189894
R2171 VN.n17 VN.n16 0.189894
R2172 VN.n18 VN.n17 0.189894
R2173 VN.n18 VN.n11 0.189894
R2174 VN.n22 VN.n11 0.189894
R2175 VN.n23 VN.n22 0.189894
R2176 VN.n24 VN.n23 0.189894
R2177 VN.n24 VN.n9 0.189894
R2178 VN.n28 VN.n9 0.189894
R2179 VN.n29 VN.n28 0.189894
R2180 VN.n30 VN.n29 0.189894
R2181 VN.n30 VN.n7 0.189894
R2182 VN.n34 VN.n7 0.189894
R2183 VN.n35 VN.n34 0.189894
R2184 VN.n36 VN.n35 0.189894
R2185 VN.n36 VN.n5 0.189894
R2186 VN.n41 VN.n5 0.189894
R2187 VN.n42 VN.n41 0.189894
R2188 VN.n43 VN.n42 0.189894
R2189 VN.n43 VN.n3 0.189894
R2190 VN.n47 VN.n3 0.189894
R2191 VN.n48 VN.n47 0.189894
R2192 VN.n49 VN.n48 0.189894
R2193 VN.n49 VN.n1 0.189894
R2194 VN.n53 VN.n1 0.189894
R2195 VDD2.n1 VDD2.t0 105.603
R2196 VDD2.n4 VDD2.t7 102.094
R2197 VDD2.n3 VDD2.n2 95.4617
R2198 VDD2 VDD2.n7 95.4591
R2199 VDD2.n6 VDD2.n5 92.8859
R2200 VDD2.n1 VDD2.n0 92.8856
R2201 VDD2.n4 VDD2.n3 42.2347
R2202 VDD2.n7 VDD2.t4 9.2098
R2203 VDD2.n7 VDD2.t5 9.2098
R2204 VDD2.n5 VDD2.t6 9.2098
R2205 VDD2.n5 VDD2.t2 9.2098
R2206 VDD2.n2 VDD2.t9 9.2098
R2207 VDD2.n2 VDD2.t8 9.2098
R2208 VDD2.n0 VDD2.t3 9.2098
R2209 VDD2.n0 VDD2.t1 9.2098
R2210 VDD2.n6 VDD2.n4 3.50912
R2211 VDD2 VDD2.n6 0.935845
R2212 VDD2.n3 VDD2.n1 0.822309
C0 VTAIL VN 4.52498f
C1 VP VDD1 3.06386f
C2 VTAIL VDD2 7.18606f
C3 VDD2 VN 2.49456f
C4 VP VTAIL 4.53917f
C5 VP VN 8.26186f
C6 VP VDD2 0.735988f
C7 VTAIL VDD1 7.12499f
C8 VN VDD1 0.162017f
C9 VDD2 VDD1 2.91513f
C10 VDD2 B 6.96253f
C11 VDD1 B 6.812512f
C12 VTAIL B 4.391224f
C13 VN B 22.872288f
C14 VP B 21.152428f
C15 VDD2.t0 B 0.47024f
C16 VDD2.t3 B 0.05141f
C17 VDD2.t1 B 0.05141f
C18 VDD2.n0 B 0.349256f
C19 VDD2.n1 B 1.2304f
C20 VDD2.t9 B 0.05141f
C21 VDD2.t8 B 0.05141f
C22 VDD2.n2 B 0.371455f
C23 VDD2.n3 B 3.48663f
C24 VDD2.t7 B 0.449951f
C25 VDD2.n4 B 3.31789f
C26 VDD2.t6 B 0.05141f
C27 VDD2.t2 B 0.05141f
C28 VDD2.n5 B 0.349256f
C29 VDD2.n6 B 0.650202f
C30 VDD2.t4 B 0.05141f
C31 VDD2.t5 B 0.05141f
C32 VDD2.n7 B 0.371416f
C33 VN.t1 B 0.48497f
C34 VN.n0 B 0.314468f
C35 VN.n1 B 0.02547f
C36 VN.n2 B 0.0465f
C37 VN.n3 B 0.02547f
C38 VN.n4 B 0.044188f
C39 VN.n5 B 0.02547f
C40 VN.n6 B 0.049544f
C41 VN.n7 B 0.02547f
C42 VN.n8 B 0.04747f
C43 VN.n9 B 0.02547f
C44 VN.t8 B 0.48497f
C45 VN.n10 B 0.051299f
C46 VN.n11 B 0.02547f
C47 VN.n12 B 0.04747f
C48 VN.t9 B 0.774223f
C49 VN.n13 B 0.33234f
C50 VN.t6 B 0.48497f
C51 VN.n14 B 0.297404f
C52 VN.n15 B 0.027315f
C53 VN.n16 B 0.323567f
C54 VN.n17 B 0.02547f
C55 VN.n18 B 0.02547f
C56 VN.n19 B 0.04747f
C57 VN.n20 B 0.049544f
C58 VN.n21 B 0.020995f
C59 VN.n22 B 0.02547f
C60 VN.n23 B 0.02547f
C61 VN.n24 B 0.02547f
C62 VN.n25 B 0.04747f
C63 VN.n26 B 0.04747f
C64 VN.n27 B 0.238788f
C65 VN.n28 B 0.02547f
C66 VN.n29 B 0.02547f
C67 VN.n30 B 0.02547f
C68 VN.n31 B 0.04747f
C69 VN.n32 B 0.051299f
C70 VN.n33 B 0.020995f
C71 VN.n34 B 0.02547f
C72 VN.n35 B 0.02547f
C73 VN.n36 B 0.02547f
C74 VN.n37 B 0.04747f
C75 VN.n38 B 0.04747f
C76 VN.t0 B 0.48497f
C77 VN.n39 B 0.214755f
C78 VN.n40 B 0.027315f
C79 VN.n41 B 0.02547f
C80 VN.n42 B 0.02547f
C81 VN.n43 B 0.02547f
C82 VN.n44 B 0.04747f
C83 VN.n45 B 0.050896f
C84 VN.n46 B 0.024442f
C85 VN.n47 B 0.02547f
C86 VN.n48 B 0.02547f
C87 VN.n49 B 0.02547f
C88 VN.n50 B 0.04747f
C89 VN.n51 B 0.04747f
C90 VN.n52 B 0.030596f
C91 VN.n53 B 0.041108f
C92 VN.n54 B 0.074217f
C93 VN.t2 B 0.48497f
C94 VN.n55 B 0.314468f
C95 VN.n56 B 0.02547f
C96 VN.n57 B 0.0465f
C97 VN.n58 B 0.02547f
C98 VN.n59 B 0.044188f
C99 VN.n60 B 0.02547f
C100 VN.t3 B 0.48497f
C101 VN.n61 B 0.214755f
C102 VN.n62 B 0.049544f
C103 VN.n63 B 0.02547f
C104 VN.n64 B 0.04747f
C105 VN.n65 B 0.02547f
C106 VN.t7 B 0.48497f
C107 VN.n66 B 0.051299f
C108 VN.n67 B 0.02547f
C109 VN.n68 B 0.04747f
C110 VN.t4 B 0.774223f
C111 VN.n69 B 0.33234f
C112 VN.t5 B 0.48497f
C113 VN.n70 B 0.297404f
C114 VN.n71 B 0.027315f
C115 VN.n72 B 0.323567f
C116 VN.n73 B 0.02547f
C117 VN.n74 B 0.02547f
C118 VN.n75 B 0.04747f
C119 VN.n76 B 0.049544f
C120 VN.n77 B 0.020995f
C121 VN.n78 B 0.02547f
C122 VN.n79 B 0.02547f
C123 VN.n80 B 0.02547f
C124 VN.n81 B 0.04747f
C125 VN.n82 B 0.04747f
C126 VN.n83 B 0.238788f
C127 VN.n84 B 0.02547f
C128 VN.n85 B 0.02547f
C129 VN.n86 B 0.02547f
C130 VN.n87 B 0.04747f
C131 VN.n88 B 0.051299f
C132 VN.n89 B 0.020995f
C133 VN.n90 B 0.02547f
C134 VN.n91 B 0.02547f
C135 VN.n92 B 0.02547f
C136 VN.n93 B 0.04747f
C137 VN.n94 B 0.04747f
C138 VN.n95 B 0.027315f
C139 VN.n96 B 0.02547f
C140 VN.n97 B 0.02547f
C141 VN.n98 B 0.02547f
C142 VN.n99 B 0.04747f
C143 VN.n100 B 0.050896f
C144 VN.n101 B 0.024442f
C145 VN.n102 B 0.02547f
C146 VN.n103 B 0.02547f
C147 VN.n104 B 0.02547f
C148 VN.n105 B 0.04747f
C149 VN.n106 B 0.04747f
C150 VN.n107 B 0.030596f
C151 VN.n108 B 0.041108f
C152 VN.n109 B 1.55414f
C153 VTAIL.t0 B 0.064944f
C154 VTAIL.t5 B 0.064944f
C155 VTAIL.n0 B 0.382822f
C156 VTAIL.n1 B 0.885668f
C157 VTAIL.t12 B 0.506571f
C158 VTAIL.n2 B 1.03991f
C159 VTAIL.t17 B 0.064944f
C160 VTAIL.t16 B 0.064944f
C161 VTAIL.n3 B 0.382822f
C162 VTAIL.n4 B 1.14475f
C163 VTAIL.t13 B 0.064944f
C164 VTAIL.t15 B 0.064944f
C165 VTAIL.n5 B 0.382822f
C166 VTAIL.n6 B 2.32443f
C167 VTAIL.t9 B 0.064944f
C168 VTAIL.t2 B 0.064944f
C169 VTAIL.n7 B 0.382823f
C170 VTAIL.n8 B 2.32443f
C171 VTAIL.t6 B 0.064944f
C172 VTAIL.t3 B 0.064944f
C173 VTAIL.n9 B 0.382823f
C174 VTAIL.n10 B 1.14475f
C175 VTAIL.t8 B 0.506574f
C176 VTAIL.n11 B 1.03991f
C177 VTAIL.t11 B 0.064944f
C178 VTAIL.t19 B 0.064944f
C179 VTAIL.n12 B 0.382823f
C180 VTAIL.n13 B 0.986538f
C181 VTAIL.t10 B 0.064944f
C182 VTAIL.t14 B 0.064944f
C183 VTAIL.n14 B 0.382823f
C184 VTAIL.n15 B 1.14475f
C185 VTAIL.t18 B 0.506571f
C186 VTAIL.n16 B 1.94565f
C187 VTAIL.t7 B 0.506571f
C188 VTAIL.n17 B 1.94565f
C189 VTAIL.t1 B 0.064944f
C190 VTAIL.t4 B 0.064944f
C191 VTAIL.n18 B 0.382822f
C192 VTAIL.n19 B 0.813465f
C193 VDD1.t1 B 0.484604f
C194 VDD1.t8 B 0.05298f
C195 VDD1.t7 B 0.05298f
C196 VDD1.n0 B 0.359923f
C197 VDD1.n1 B 1.27851f
C198 VDD1.t9 B 0.484602f
C199 VDD1.t2 B 0.05298f
C200 VDD1.t3 B 0.05298f
C201 VDD1.n2 B 0.359923f
C202 VDD1.n3 B 1.26798f
C203 VDD1.t6 B 0.05298f
C204 VDD1.t0 B 0.05298f
C205 VDD1.n4 B 0.3828f
C206 VDD1.n5 B 3.77569f
C207 VDD1.t4 B 0.05298f
C208 VDD1.t5 B 0.05298f
C209 VDD1.n6 B 0.359922f
C210 VDD1.n7 B 3.56966f
C211 VP.t7 B 0.505171f
C212 VP.n0 B 0.327567f
C213 VP.n1 B 0.026531f
C214 VP.n2 B 0.048437f
C215 VP.n3 B 0.026531f
C216 VP.n4 B 0.046029f
C217 VP.n5 B 0.026531f
C218 VP.n6 B 0.051608f
C219 VP.n7 B 0.026531f
C220 VP.n8 B 0.049447f
C221 VP.n9 B 0.026531f
C222 VP.t2 B 0.505171f
C223 VP.n10 B 0.053436f
C224 VP.n11 B 0.026531f
C225 VP.n12 B 0.049447f
C226 VP.n13 B 0.026531f
C227 VP.t4 B 0.505171f
C228 VP.n14 B 0.053016f
C229 VP.n15 B 0.026531f
C230 VP.n16 B 0.049447f
C231 VP.t1 B 0.505171f
C232 VP.n17 B 0.327567f
C233 VP.n18 B 0.026531f
C234 VP.n19 B 0.048437f
C235 VP.n20 B 0.026531f
C236 VP.n21 B 0.046029f
C237 VP.n22 B 0.026531f
C238 VP.n23 B 0.051608f
C239 VP.n24 B 0.026531f
C240 VP.n25 B 0.049447f
C241 VP.n26 B 0.026531f
C242 VP.t9 B 0.505171f
C243 VP.n27 B 0.053436f
C244 VP.n28 B 0.026531f
C245 VP.n29 B 0.049447f
C246 VP.t8 B 0.806471f
C247 VP.n30 B 0.346184f
C248 VP.t0 B 0.505171f
C249 VP.n31 B 0.309792f
C250 VP.n32 B 0.028452f
C251 VP.n33 B 0.337045f
C252 VP.n34 B 0.026531f
C253 VP.n35 B 0.026531f
C254 VP.n36 B 0.049447f
C255 VP.n37 B 0.051608f
C256 VP.n38 B 0.021869f
C257 VP.n39 B 0.026531f
C258 VP.n40 B 0.026531f
C259 VP.n41 B 0.026531f
C260 VP.n42 B 0.049447f
C261 VP.n43 B 0.049447f
C262 VP.n44 B 0.248734f
C263 VP.n45 B 0.026531f
C264 VP.n46 B 0.026531f
C265 VP.n47 B 0.026531f
C266 VP.n48 B 0.049447f
C267 VP.n49 B 0.053436f
C268 VP.n50 B 0.021869f
C269 VP.n51 B 0.026531f
C270 VP.n52 B 0.026531f
C271 VP.n53 B 0.026531f
C272 VP.n54 B 0.049447f
C273 VP.n55 B 0.049447f
C274 VP.t5 B 0.505171f
C275 VP.n56 B 0.2237f
C276 VP.n57 B 0.028452f
C277 VP.n58 B 0.026531f
C278 VP.n59 B 0.026531f
C279 VP.n60 B 0.026531f
C280 VP.n61 B 0.049447f
C281 VP.n62 B 0.053016f
C282 VP.n63 B 0.02546f
C283 VP.n64 B 0.026531f
C284 VP.n65 B 0.026531f
C285 VP.n66 B 0.026531f
C286 VP.n67 B 0.049447f
C287 VP.n68 B 0.049447f
C288 VP.n69 B 0.03187f
C289 VP.n70 B 0.04282f
C290 VP.n71 B 1.60817f
C291 VP.n72 B 1.62652f
C292 VP.t6 B 0.505171f
C293 VP.n73 B 0.327567f
C294 VP.n74 B 0.03187f
C295 VP.n75 B 0.04282f
C296 VP.n76 B 0.026531f
C297 VP.n77 B 0.026531f
C298 VP.n78 B 0.049447f
C299 VP.n79 B 0.048437f
C300 VP.n80 B 0.02546f
C301 VP.n81 B 0.026531f
C302 VP.n82 B 0.026531f
C303 VP.n83 B 0.026531f
C304 VP.n84 B 0.049447f
C305 VP.n85 B 0.046029f
C306 VP.n86 B 0.2237f
C307 VP.n87 B 0.028452f
C308 VP.n88 B 0.026531f
C309 VP.n89 B 0.026531f
C310 VP.n90 B 0.026531f
C311 VP.n91 B 0.049447f
C312 VP.n92 B 0.051608f
C313 VP.n93 B 0.021869f
C314 VP.n94 B 0.026531f
C315 VP.n95 B 0.026531f
C316 VP.n96 B 0.026531f
C317 VP.n97 B 0.049447f
C318 VP.n98 B 0.049447f
C319 VP.n99 B 0.248734f
C320 VP.n100 B 0.026531f
C321 VP.n101 B 0.026531f
C322 VP.n102 B 0.026531f
C323 VP.n103 B 0.049447f
C324 VP.n104 B 0.053436f
C325 VP.n105 B 0.021869f
C326 VP.n106 B 0.026531f
C327 VP.n107 B 0.026531f
C328 VP.n108 B 0.026531f
C329 VP.n109 B 0.049447f
C330 VP.n110 B 0.049447f
C331 VP.t3 B 0.505171f
C332 VP.n111 B 0.2237f
C333 VP.n112 B 0.028452f
C334 VP.n113 B 0.026531f
C335 VP.n114 B 0.026531f
C336 VP.n115 B 0.026531f
C337 VP.n116 B 0.049447f
C338 VP.n117 B 0.053016f
C339 VP.n118 B 0.02546f
C340 VP.n119 B 0.026531f
C341 VP.n120 B 0.026531f
C342 VP.n121 B 0.026531f
C343 VP.n122 B 0.049447f
C344 VP.n123 B 0.049447f
C345 VP.n124 B 0.03187f
C346 VP.n125 B 0.04282f
C347 VP.n126 B 0.077309f
.ends

