* NGSPICE file created from diff_pair_sample_0761.ext - technology: sky130A

.subckt diff_pair_sample_0761 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t9 VN.t0 VTAIL.t11 w_n2794_n4356# sky130_fd_pr__pfet_01v8 ad=2.7951 pd=17.27 as=2.7951 ps=17.27 w=16.94 l=1.19
X1 B.t11 B.t9 B.t10 w_n2794_n4356# sky130_fd_pr__pfet_01v8 ad=6.6066 pd=34.66 as=0 ps=0 w=16.94 l=1.19
X2 VDD2.t8 VN.t1 VTAIL.t9 w_n2794_n4356# sky130_fd_pr__pfet_01v8 ad=2.7951 pd=17.27 as=2.7951 ps=17.27 w=16.94 l=1.19
X3 VDD1.t9 VP.t0 VTAIL.t5 w_n2794_n4356# sky130_fd_pr__pfet_01v8 ad=2.7951 pd=17.27 as=2.7951 ps=17.27 w=16.94 l=1.19
X4 B.t8 B.t6 B.t7 w_n2794_n4356# sky130_fd_pr__pfet_01v8 ad=6.6066 pd=34.66 as=0 ps=0 w=16.94 l=1.19
X5 VTAIL.t7 VP.t1 VDD1.t8 w_n2794_n4356# sky130_fd_pr__pfet_01v8 ad=2.7951 pd=17.27 as=2.7951 ps=17.27 w=16.94 l=1.19
X6 VTAIL.t10 VN.t2 VDD2.t7 w_n2794_n4356# sky130_fd_pr__pfet_01v8 ad=2.7951 pd=17.27 as=2.7951 ps=17.27 w=16.94 l=1.19
X7 VDD2.t6 VN.t3 VTAIL.t12 w_n2794_n4356# sky130_fd_pr__pfet_01v8 ad=6.6066 pd=34.66 as=2.7951 ps=17.27 w=16.94 l=1.19
X8 VDD1.t7 VP.t2 VTAIL.t4 w_n2794_n4356# sky130_fd_pr__pfet_01v8 ad=2.7951 pd=17.27 as=6.6066 ps=34.66 w=16.94 l=1.19
X9 VTAIL.t13 VN.t4 VDD2.t5 w_n2794_n4356# sky130_fd_pr__pfet_01v8 ad=2.7951 pd=17.27 as=2.7951 ps=17.27 w=16.94 l=1.19
X10 VDD1.t6 VP.t3 VTAIL.t0 w_n2794_n4356# sky130_fd_pr__pfet_01v8 ad=6.6066 pd=34.66 as=2.7951 ps=17.27 w=16.94 l=1.19
X11 VDD2.t4 VN.t5 VTAIL.t16 w_n2794_n4356# sky130_fd_pr__pfet_01v8 ad=2.7951 pd=17.27 as=6.6066 ps=34.66 w=16.94 l=1.19
X12 VTAIL.t18 VP.t4 VDD1.t5 w_n2794_n4356# sky130_fd_pr__pfet_01v8 ad=2.7951 pd=17.27 as=2.7951 ps=17.27 w=16.94 l=1.19
X13 VDD1.t4 VP.t5 VTAIL.t6 w_n2794_n4356# sky130_fd_pr__pfet_01v8 ad=2.7951 pd=17.27 as=6.6066 ps=34.66 w=16.94 l=1.19
X14 VTAIL.t8 VN.t6 VDD2.t3 w_n2794_n4356# sky130_fd_pr__pfet_01v8 ad=2.7951 pd=17.27 as=2.7951 ps=17.27 w=16.94 l=1.19
X15 B.t5 B.t3 B.t4 w_n2794_n4356# sky130_fd_pr__pfet_01v8 ad=6.6066 pd=34.66 as=0 ps=0 w=16.94 l=1.19
X16 VTAIL.t2 VP.t6 VDD1.t3 w_n2794_n4356# sky130_fd_pr__pfet_01v8 ad=2.7951 pd=17.27 as=2.7951 ps=17.27 w=16.94 l=1.19
X17 VDD2.t2 VN.t7 VTAIL.t17 w_n2794_n4356# sky130_fd_pr__pfet_01v8 ad=6.6066 pd=34.66 as=2.7951 ps=17.27 w=16.94 l=1.19
X18 VTAIL.t19 VP.t7 VDD1.t2 w_n2794_n4356# sky130_fd_pr__pfet_01v8 ad=2.7951 pd=17.27 as=2.7951 ps=17.27 w=16.94 l=1.19
X19 B.t2 B.t0 B.t1 w_n2794_n4356# sky130_fd_pr__pfet_01v8 ad=6.6066 pd=34.66 as=0 ps=0 w=16.94 l=1.19
X20 VDD2.t1 VN.t8 VTAIL.t15 w_n2794_n4356# sky130_fd_pr__pfet_01v8 ad=2.7951 pd=17.27 as=6.6066 ps=34.66 w=16.94 l=1.19
X21 VTAIL.t14 VN.t9 VDD2.t0 w_n2794_n4356# sky130_fd_pr__pfet_01v8 ad=2.7951 pd=17.27 as=2.7951 ps=17.27 w=16.94 l=1.19
X22 VDD1.t1 VP.t8 VTAIL.t3 w_n2794_n4356# sky130_fd_pr__pfet_01v8 ad=6.6066 pd=34.66 as=2.7951 ps=17.27 w=16.94 l=1.19
X23 VDD1.t0 VP.t9 VTAIL.t1 w_n2794_n4356# sky130_fd_pr__pfet_01v8 ad=2.7951 pd=17.27 as=2.7951 ps=17.27 w=16.94 l=1.19
R0 VN.n6 VN.t3 394.978
R1 VN.n28 VN.t5 394.978
R2 VN.n20 VN.t8 376.488
R3 VN.n42 VN.t7 376.488
R4 VN.n5 VN.t6 343.072
R5 VN.n3 VN.t1 343.072
R6 VN.n1 VN.t4 343.072
R7 VN.n27 VN.t2 343.072
R8 VN.n25 VN.t0 343.072
R9 VN.n23 VN.t9 343.072
R10 VN.n41 VN.n22 161.3
R11 VN.n40 VN.n39 161.3
R12 VN.n38 VN.n37 161.3
R13 VN.n36 VN.n24 161.3
R14 VN.n35 VN.n34 161.3
R15 VN.n33 VN.n32 161.3
R16 VN.n31 VN.n26 161.3
R17 VN.n30 VN.n29 161.3
R18 VN.n19 VN.n0 161.3
R19 VN.n18 VN.n17 161.3
R20 VN.n16 VN.n15 161.3
R21 VN.n14 VN.n2 161.3
R22 VN.n13 VN.n12 161.3
R23 VN.n11 VN.n10 161.3
R24 VN.n9 VN.n4 161.3
R25 VN.n8 VN.n7 161.3
R26 VN.n43 VN.n42 80.6037
R27 VN.n21 VN.n20 80.6037
R28 VN VN.n43 49.5824
R29 VN.n6 VN.n5 44.4551
R30 VN.n28 VN.n27 44.4551
R31 VN.n9 VN.n8 41.3843
R32 VN.n15 VN.n14 41.3843
R33 VN.n31 VN.n30 41.3843
R34 VN.n37 VN.n36 41.3843
R35 VN.n10 VN.n9 39.4369
R36 VN.n14 VN.n13 39.4369
R37 VN.n32 VN.n31 39.4369
R38 VN.n36 VN.n35 39.4369
R39 VN.n19 VN.n18 37.4894
R40 VN.n41 VN.n40 37.4894
R41 VN.n29 VN.n28 29.7405
R42 VN.n7 VN.n6 29.7405
R43 VN.n20 VN.n19 28.4823
R44 VN.n42 VN.n41 28.4823
R45 VN.n8 VN.n5 13.146
R46 VN.n15 VN.n1 13.146
R47 VN.n30 VN.n27 13.146
R48 VN.n37 VN.n23 13.146
R49 VN.n10 VN.n3 12.1722
R50 VN.n13 VN.n3 12.1722
R51 VN.n35 VN.n25 12.1722
R52 VN.n32 VN.n25 12.1722
R53 VN.n18 VN.n1 11.1985
R54 VN.n40 VN.n23 11.1985
R55 VN.n43 VN.n22 0.285035
R56 VN.n21 VN.n0 0.285035
R57 VN.n39 VN.n22 0.189894
R58 VN.n39 VN.n38 0.189894
R59 VN.n38 VN.n24 0.189894
R60 VN.n34 VN.n24 0.189894
R61 VN.n34 VN.n33 0.189894
R62 VN.n33 VN.n26 0.189894
R63 VN.n29 VN.n26 0.189894
R64 VN.n7 VN.n4 0.189894
R65 VN.n11 VN.n4 0.189894
R66 VN.n12 VN.n11 0.189894
R67 VN.n12 VN.n2 0.189894
R68 VN.n16 VN.n2 0.189894
R69 VN.n17 VN.n16 0.189894
R70 VN.n17 VN.n0 0.189894
R71 VN VN.n21 0.146778
R72 VTAIL.n384 VTAIL.n296 756.745
R73 VTAIL.n90 VTAIL.n2 756.745
R74 VTAIL.n290 VTAIL.n202 756.745
R75 VTAIL.n192 VTAIL.n104 756.745
R76 VTAIL.n327 VTAIL.n326 585
R77 VTAIL.n324 VTAIL.n323 585
R78 VTAIL.n333 VTAIL.n332 585
R79 VTAIL.n335 VTAIL.n334 585
R80 VTAIL.n320 VTAIL.n319 585
R81 VTAIL.n341 VTAIL.n340 585
R82 VTAIL.n343 VTAIL.n342 585
R83 VTAIL.n316 VTAIL.n315 585
R84 VTAIL.n349 VTAIL.n348 585
R85 VTAIL.n351 VTAIL.n350 585
R86 VTAIL.n312 VTAIL.n311 585
R87 VTAIL.n357 VTAIL.n356 585
R88 VTAIL.n359 VTAIL.n358 585
R89 VTAIL.n308 VTAIL.n307 585
R90 VTAIL.n365 VTAIL.n364 585
R91 VTAIL.n368 VTAIL.n367 585
R92 VTAIL.n366 VTAIL.n304 585
R93 VTAIL.n373 VTAIL.n303 585
R94 VTAIL.n375 VTAIL.n374 585
R95 VTAIL.n377 VTAIL.n376 585
R96 VTAIL.n300 VTAIL.n299 585
R97 VTAIL.n383 VTAIL.n382 585
R98 VTAIL.n385 VTAIL.n384 585
R99 VTAIL.n33 VTAIL.n32 585
R100 VTAIL.n30 VTAIL.n29 585
R101 VTAIL.n39 VTAIL.n38 585
R102 VTAIL.n41 VTAIL.n40 585
R103 VTAIL.n26 VTAIL.n25 585
R104 VTAIL.n47 VTAIL.n46 585
R105 VTAIL.n49 VTAIL.n48 585
R106 VTAIL.n22 VTAIL.n21 585
R107 VTAIL.n55 VTAIL.n54 585
R108 VTAIL.n57 VTAIL.n56 585
R109 VTAIL.n18 VTAIL.n17 585
R110 VTAIL.n63 VTAIL.n62 585
R111 VTAIL.n65 VTAIL.n64 585
R112 VTAIL.n14 VTAIL.n13 585
R113 VTAIL.n71 VTAIL.n70 585
R114 VTAIL.n74 VTAIL.n73 585
R115 VTAIL.n72 VTAIL.n10 585
R116 VTAIL.n79 VTAIL.n9 585
R117 VTAIL.n81 VTAIL.n80 585
R118 VTAIL.n83 VTAIL.n82 585
R119 VTAIL.n6 VTAIL.n5 585
R120 VTAIL.n89 VTAIL.n88 585
R121 VTAIL.n91 VTAIL.n90 585
R122 VTAIL.n291 VTAIL.n290 585
R123 VTAIL.n289 VTAIL.n288 585
R124 VTAIL.n206 VTAIL.n205 585
R125 VTAIL.n283 VTAIL.n282 585
R126 VTAIL.n281 VTAIL.n280 585
R127 VTAIL.n279 VTAIL.n209 585
R128 VTAIL.n213 VTAIL.n210 585
R129 VTAIL.n274 VTAIL.n273 585
R130 VTAIL.n272 VTAIL.n271 585
R131 VTAIL.n215 VTAIL.n214 585
R132 VTAIL.n266 VTAIL.n265 585
R133 VTAIL.n264 VTAIL.n263 585
R134 VTAIL.n219 VTAIL.n218 585
R135 VTAIL.n258 VTAIL.n257 585
R136 VTAIL.n256 VTAIL.n255 585
R137 VTAIL.n223 VTAIL.n222 585
R138 VTAIL.n250 VTAIL.n249 585
R139 VTAIL.n248 VTAIL.n247 585
R140 VTAIL.n227 VTAIL.n226 585
R141 VTAIL.n242 VTAIL.n241 585
R142 VTAIL.n240 VTAIL.n239 585
R143 VTAIL.n231 VTAIL.n230 585
R144 VTAIL.n234 VTAIL.n233 585
R145 VTAIL.n193 VTAIL.n192 585
R146 VTAIL.n191 VTAIL.n190 585
R147 VTAIL.n108 VTAIL.n107 585
R148 VTAIL.n185 VTAIL.n184 585
R149 VTAIL.n183 VTAIL.n182 585
R150 VTAIL.n181 VTAIL.n111 585
R151 VTAIL.n115 VTAIL.n112 585
R152 VTAIL.n176 VTAIL.n175 585
R153 VTAIL.n174 VTAIL.n173 585
R154 VTAIL.n117 VTAIL.n116 585
R155 VTAIL.n168 VTAIL.n167 585
R156 VTAIL.n166 VTAIL.n165 585
R157 VTAIL.n121 VTAIL.n120 585
R158 VTAIL.n160 VTAIL.n159 585
R159 VTAIL.n158 VTAIL.n157 585
R160 VTAIL.n125 VTAIL.n124 585
R161 VTAIL.n152 VTAIL.n151 585
R162 VTAIL.n150 VTAIL.n149 585
R163 VTAIL.n129 VTAIL.n128 585
R164 VTAIL.n144 VTAIL.n143 585
R165 VTAIL.n142 VTAIL.n141 585
R166 VTAIL.n133 VTAIL.n132 585
R167 VTAIL.n136 VTAIL.n135 585
R168 VTAIL.t6 VTAIL.n232 327.466
R169 VTAIL.t16 VTAIL.n134 327.466
R170 VTAIL.t15 VTAIL.n325 327.466
R171 VTAIL.t4 VTAIL.n31 327.466
R172 VTAIL.n326 VTAIL.n323 171.744
R173 VTAIL.n333 VTAIL.n323 171.744
R174 VTAIL.n334 VTAIL.n333 171.744
R175 VTAIL.n334 VTAIL.n319 171.744
R176 VTAIL.n341 VTAIL.n319 171.744
R177 VTAIL.n342 VTAIL.n341 171.744
R178 VTAIL.n342 VTAIL.n315 171.744
R179 VTAIL.n349 VTAIL.n315 171.744
R180 VTAIL.n350 VTAIL.n349 171.744
R181 VTAIL.n350 VTAIL.n311 171.744
R182 VTAIL.n357 VTAIL.n311 171.744
R183 VTAIL.n358 VTAIL.n357 171.744
R184 VTAIL.n358 VTAIL.n307 171.744
R185 VTAIL.n365 VTAIL.n307 171.744
R186 VTAIL.n367 VTAIL.n365 171.744
R187 VTAIL.n367 VTAIL.n366 171.744
R188 VTAIL.n366 VTAIL.n303 171.744
R189 VTAIL.n375 VTAIL.n303 171.744
R190 VTAIL.n376 VTAIL.n375 171.744
R191 VTAIL.n376 VTAIL.n299 171.744
R192 VTAIL.n383 VTAIL.n299 171.744
R193 VTAIL.n384 VTAIL.n383 171.744
R194 VTAIL.n32 VTAIL.n29 171.744
R195 VTAIL.n39 VTAIL.n29 171.744
R196 VTAIL.n40 VTAIL.n39 171.744
R197 VTAIL.n40 VTAIL.n25 171.744
R198 VTAIL.n47 VTAIL.n25 171.744
R199 VTAIL.n48 VTAIL.n47 171.744
R200 VTAIL.n48 VTAIL.n21 171.744
R201 VTAIL.n55 VTAIL.n21 171.744
R202 VTAIL.n56 VTAIL.n55 171.744
R203 VTAIL.n56 VTAIL.n17 171.744
R204 VTAIL.n63 VTAIL.n17 171.744
R205 VTAIL.n64 VTAIL.n63 171.744
R206 VTAIL.n64 VTAIL.n13 171.744
R207 VTAIL.n71 VTAIL.n13 171.744
R208 VTAIL.n73 VTAIL.n71 171.744
R209 VTAIL.n73 VTAIL.n72 171.744
R210 VTAIL.n72 VTAIL.n9 171.744
R211 VTAIL.n81 VTAIL.n9 171.744
R212 VTAIL.n82 VTAIL.n81 171.744
R213 VTAIL.n82 VTAIL.n5 171.744
R214 VTAIL.n89 VTAIL.n5 171.744
R215 VTAIL.n90 VTAIL.n89 171.744
R216 VTAIL.n290 VTAIL.n289 171.744
R217 VTAIL.n289 VTAIL.n205 171.744
R218 VTAIL.n282 VTAIL.n205 171.744
R219 VTAIL.n282 VTAIL.n281 171.744
R220 VTAIL.n281 VTAIL.n209 171.744
R221 VTAIL.n213 VTAIL.n209 171.744
R222 VTAIL.n273 VTAIL.n213 171.744
R223 VTAIL.n273 VTAIL.n272 171.744
R224 VTAIL.n272 VTAIL.n214 171.744
R225 VTAIL.n265 VTAIL.n214 171.744
R226 VTAIL.n265 VTAIL.n264 171.744
R227 VTAIL.n264 VTAIL.n218 171.744
R228 VTAIL.n257 VTAIL.n218 171.744
R229 VTAIL.n257 VTAIL.n256 171.744
R230 VTAIL.n256 VTAIL.n222 171.744
R231 VTAIL.n249 VTAIL.n222 171.744
R232 VTAIL.n249 VTAIL.n248 171.744
R233 VTAIL.n248 VTAIL.n226 171.744
R234 VTAIL.n241 VTAIL.n226 171.744
R235 VTAIL.n241 VTAIL.n240 171.744
R236 VTAIL.n240 VTAIL.n230 171.744
R237 VTAIL.n233 VTAIL.n230 171.744
R238 VTAIL.n192 VTAIL.n191 171.744
R239 VTAIL.n191 VTAIL.n107 171.744
R240 VTAIL.n184 VTAIL.n107 171.744
R241 VTAIL.n184 VTAIL.n183 171.744
R242 VTAIL.n183 VTAIL.n111 171.744
R243 VTAIL.n115 VTAIL.n111 171.744
R244 VTAIL.n175 VTAIL.n115 171.744
R245 VTAIL.n175 VTAIL.n174 171.744
R246 VTAIL.n174 VTAIL.n116 171.744
R247 VTAIL.n167 VTAIL.n116 171.744
R248 VTAIL.n167 VTAIL.n166 171.744
R249 VTAIL.n166 VTAIL.n120 171.744
R250 VTAIL.n159 VTAIL.n120 171.744
R251 VTAIL.n159 VTAIL.n158 171.744
R252 VTAIL.n158 VTAIL.n124 171.744
R253 VTAIL.n151 VTAIL.n124 171.744
R254 VTAIL.n151 VTAIL.n150 171.744
R255 VTAIL.n150 VTAIL.n128 171.744
R256 VTAIL.n143 VTAIL.n128 171.744
R257 VTAIL.n143 VTAIL.n142 171.744
R258 VTAIL.n142 VTAIL.n132 171.744
R259 VTAIL.n135 VTAIL.n132 171.744
R260 VTAIL.n326 VTAIL.t15 85.8723
R261 VTAIL.n32 VTAIL.t4 85.8723
R262 VTAIL.n233 VTAIL.t6 85.8723
R263 VTAIL.n135 VTAIL.t16 85.8723
R264 VTAIL.n201 VTAIL.n200 55.4284
R265 VTAIL.n199 VTAIL.n198 55.4284
R266 VTAIL.n103 VTAIL.n102 55.4284
R267 VTAIL.n101 VTAIL.n100 55.4284
R268 VTAIL.n391 VTAIL.n390 55.4282
R269 VTAIL.n1 VTAIL.n0 55.4282
R270 VTAIL.n97 VTAIL.n96 55.4282
R271 VTAIL.n99 VTAIL.n98 55.4282
R272 VTAIL.n389 VTAIL.n388 34.9005
R273 VTAIL.n95 VTAIL.n94 34.9005
R274 VTAIL.n295 VTAIL.n294 34.9005
R275 VTAIL.n197 VTAIL.n196 34.9005
R276 VTAIL.n101 VTAIL.n99 29.591
R277 VTAIL.n389 VTAIL.n295 28.2807
R278 VTAIL.n327 VTAIL.n325 16.3895
R279 VTAIL.n33 VTAIL.n31 16.3895
R280 VTAIL.n234 VTAIL.n232 16.3895
R281 VTAIL.n136 VTAIL.n134 16.3895
R282 VTAIL.n374 VTAIL.n373 13.1884
R283 VTAIL.n80 VTAIL.n79 13.1884
R284 VTAIL.n280 VTAIL.n279 13.1884
R285 VTAIL.n182 VTAIL.n181 13.1884
R286 VTAIL.n328 VTAIL.n324 12.8005
R287 VTAIL.n372 VTAIL.n304 12.8005
R288 VTAIL.n377 VTAIL.n302 12.8005
R289 VTAIL.n34 VTAIL.n30 12.8005
R290 VTAIL.n78 VTAIL.n10 12.8005
R291 VTAIL.n83 VTAIL.n8 12.8005
R292 VTAIL.n283 VTAIL.n208 12.8005
R293 VTAIL.n278 VTAIL.n210 12.8005
R294 VTAIL.n235 VTAIL.n231 12.8005
R295 VTAIL.n185 VTAIL.n110 12.8005
R296 VTAIL.n180 VTAIL.n112 12.8005
R297 VTAIL.n137 VTAIL.n133 12.8005
R298 VTAIL.n332 VTAIL.n331 12.0247
R299 VTAIL.n369 VTAIL.n368 12.0247
R300 VTAIL.n378 VTAIL.n300 12.0247
R301 VTAIL.n38 VTAIL.n37 12.0247
R302 VTAIL.n75 VTAIL.n74 12.0247
R303 VTAIL.n84 VTAIL.n6 12.0247
R304 VTAIL.n284 VTAIL.n206 12.0247
R305 VTAIL.n275 VTAIL.n274 12.0247
R306 VTAIL.n239 VTAIL.n238 12.0247
R307 VTAIL.n186 VTAIL.n108 12.0247
R308 VTAIL.n177 VTAIL.n176 12.0247
R309 VTAIL.n141 VTAIL.n140 12.0247
R310 VTAIL.n335 VTAIL.n322 11.249
R311 VTAIL.n364 VTAIL.n306 11.249
R312 VTAIL.n382 VTAIL.n381 11.249
R313 VTAIL.n41 VTAIL.n28 11.249
R314 VTAIL.n70 VTAIL.n12 11.249
R315 VTAIL.n88 VTAIL.n87 11.249
R316 VTAIL.n288 VTAIL.n287 11.249
R317 VTAIL.n271 VTAIL.n212 11.249
R318 VTAIL.n242 VTAIL.n229 11.249
R319 VTAIL.n190 VTAIL.n189 11.249
R320 VTAIL.n173 VTAIL.n114 11.249
R321 VTAIL.n144 VTAIL.n131 11.249
R322 VTAIL.n336 VTAIL.n320 10.4732
R323 VTAIL.n363 VTAIL.n308 10.4732
R324 VTAIL.n385 VTAIL.n298 10.4732
R325 VTAIL.n42 VTAIL.n26 10.4732
R326 VTAIL.n69 VTAIL.n14 10.4732
R327 VTAIL.n91 VTAIL.n4 10.4732
R328 VTAIL.n291 VTAIL.n204 10.4732
R329 VTAIL.n270 VTAIL.n215 10.4732
R330 VTAIL.n243 VTAIL.n227 10.4732
R331 VTAIL.n193 VTAIL.n106 10.4732
R332 VTAIL.n172 VTAIL.n117 10.4732
R333 VTAIL.n145 VTAIL.n129 10.4732
R334 VTAIL.n340 VTAIL.n339 9.69747
R335 VTAIL.n360 VTAIL.n359 9.69747
R336 VTAIL.n386 VTAIL.n296 9.69747
R337 VTAIL.n46 VTAIL.n45 9.69747
R338 VTAIL.n66 VTAIL.n65 9.69747
R339 VTAIL.n92 VTAIL.n2 9.69747
R340 VTAIL.n292 VTAIL.n202 9.69747
R341 VTAIL.n267 VTAIL.n266 9.69747
R342 VTAIL.n247 VTAIL.n246 9.69747
R343 VTAIL.n194 VTAIL.n104 9.69747
R344 VTAIL.n169 VTAIL.n168 9.69747
R345 VTAIL.n149 VTAIL.n148 9.69747
R346 VTAIL.n388 VTAIL.n387 9.45567
R347 VTAIL.n94 VTAIL.n93 9.45567
R348 VTAIL.n294 VTAIL.n293 9.45567
R349 VTAIL.n196 VTAIL.n195 9.45567
R350 VTAIL.n387 VTAIL.n386 9.3005
R351 VTAIL.n298 VTAIL.n297 9.3005
R352 VTAIL.n381 VTAIL.n380 9.3005
R353 VTAIL.n379 VTAIL.n378 9.3005
R354 VTAIL.n302 VTAIL.n301 9.3005
R355 VTAIL.n347 VTAIL.n346 9.3005
R356 VTAIL.n345 VTAIL.n344 9.3005
R357 VTAIL.n318 VTAIL.n317 9.3005
R358 VTAIL.n339 VTAIL.n338 9.3005
R359 VTAIL.n337 VTAIL.n336 9.3005
R360 VTAIL.n322 VTAIL.n321 9.3005
R361 VTAIL.n331 VTAIL.n330 9.3005
R362 VTAIL.n329 VTAIL.n328 9.3005
R363 VTAIL.n314 VTAIL.n313 9.3005
R364 VTAIL.n353 VTAIL.n352 9.3005
R365 VTAIL.n355 VTAIL.n354 9.3005
R366 VTAIL.n310 VTAIL.n309 9.3005
R367 VTAIL.n361 VTAIL.n360 9.3005
R368 VTAIL.n363 VTAIL.n362 9.3005
R369 VTAIL.n306 VTAIL.n305 9.3005
R370 VTAIL.n370 VTAIL.n369 9.3005
R371 VTAIL.n372 VTAIL.n371 9.3005
R372 VTAIL.n93 VTAIL.n92 9.3005
R373 VTAIL.n4 VTAIL.n3 9.3005
R374 VTAIL.n87 VTAIL.n86 9.3005
R375 VTAIL.n85 VTAIL.n84 9.3005
R376 VTAIL.n8 VTAIL.n7 9.3005
R377 VTAIL.n53 VTAIL.n52 9.3005
R378 VTAIL.n51 VTAIL.n50 9.3005
R379 VTAIL.n24 VTAIL.n23 9.3005
R380 VTAIL.n45 VTAIL.n44 9.3005
R381 VTAIL.n43 VTAIL.n42 9.3005
R382 VTAIL.n28 VTAIL.n27 9.3005
R383 VTAIL.n37 VTAIL.n36 9.3005
R384 VTAIL.n35 VTAIL.n34 9.3005
R385 VTAIL.n20 VTAIL.n19 9.3005
R386 VTAIL.n59 VTAIL.n58 9.3005
R387 VTAIL.n61 VTAIL.n60 9.3005
R388 VTAIL.n16 VTAIL.n15 9.3005
R389 VTAIL.n67 VTAIL.n66 9.3005
R390 VTAIL.n69 VTAIL.n68 9.3005
R391 VTAIL.n12 VTAIL.n11 9.3005
R392 VTAIL.n76 VTAIL.n75 9.3005
R393 VTAIL.n78 VTAIL.n77 9.3005
R394 VTAIL.n260 VTAIL.n259 9.3005
R395 VTAIL.n262 VTAIL.n261 9.3005
R396 VTAIL.n217 VTAIL.n216 9.3005
R397 VTAIL.n268 VTAIL.n267 9.3005
R398 VTAIL.n270 VTAIL.n269 9.3005
R399 VTAIL.n212 VTAIL.n211 9.3005
R400 VTAIL.n276 VTAIL.n275 9.3005
R401 VTAIL.n278 VTAIL.n277 9.3005
R402 VTAIL.n293 VTAIL.n292 9.3005
R403 VTAIL.n204 VTAIL.n203 9.3005
R404 VTAIL.n287 VTAIL.n286 9.3005
R405 VTAIL.n285 VTAIL.n284 9.3005
R406 VTAIL.n208 VTAIL.n207 9.3005
R407 VTAIL.n221 VTAIL.n220 9.3005
R408 VTAIL.n254 VTAIL.n253 9.3005
R409 VTAIL.n252 VTAIL.n251 9.3005
R410 VTAIL.n225 VTAIL.n224 9.3005
R411 VTAIL.n246 VTAIL.n245 9.3005
R412 VTAIL.n244 VTAIL.n243 9.3005
R413 VTAIL.n229 VTAIL.n228 9.3005
R414 VTAIL.n238 VTAIL.n237 9.3005
R415 VTAIL.n236 VTAIL.n235 9.3005
R416 VTAIL.n162 VTAIL.n161 9.3005
R417 VTAIL.n164 VTAIL.n163 9.3005
R418 VTAIL.n119 VTAIL.n118 9.3005
R419 VTAIL.n170 VTAIL.n169 9.3005
R420 VTAIL.n172 VTAIL.n171 9.3005
R421 VTAIL.n114 VTAIL.n113 9.3005
R422 VTAIL.n178 VTAIL.n177 9.3005
R423 VTAIL.n180 VTAIL.n179 9.3005
R424 VTAIL.n195 VTAIL.n194 9.3005
R425 VTAIL.n106 VTAIL.n105 9.3005
R426 VTAIL.n189 VTAIL.n188 9.3005
R427 VTAIL.n187 VTAIL.n186 9.3005
R428 VTAIL.n110 VTAIL.n109 9.3005
R429 VTAIL.n123 VTAIL.n122 9.3005
R430 VTAIL.n156 VTAIL.n155 9.3005
R431 VTAIL.n154 VTAIL.n153 9.3005
R432 VTAIL.n127 VTAIL.n126 9.3005
R433 VTAIL.n148 VTAIL.n147 9.3005
R434 VTAIL.n146 VTAIL.n145 9.3005
R435 VTAIL.n131 VTAIL.n130 9.3005
R436 VTAIL.n140 VTAIL.n139 9.3005
R437 VTAIL.n138 VTAIL.n137 9.3005
R438 VTAIL.n343 VTAIL.n318 8.92171
R439 VTAIL.n356 VTAIL.n310 8.92171
R440 VTAIL.n49 VTAIL.n24 8.92171
R441 VTAIL.n62 VTAIL.n16 8.92171
R442 VTAIL.n263 VTAIL.n217 8.92171
R443 VTAIL.n250 VTAIL.n225 8.92171
R444 VTAIL.n165 VTAIL.n119 8.92171
R445 VTAIL.n152 VTAIL.n127 8.92171
R446 VTAIL.n344 VTAIL.n316 8.14595
R447 VTAIL.n355 VTAIL.n312 8.14595
R448 VTAIL.n50 VTAIL.n22 8.14595
R449 VTAIL.n61 VTAIL.n18 8.14595
R450 VTAIL.n262 VTAIL.n219 8.14595
R451 VTAIL.n251 VTAIL.n223 8.14595
R452 VTAIL.n164 VTAIL.n121 8.14595
R453 VTAIL.n153 VTAIL.n125 8.14595
R454 VTAIL.n348 VTAIL.n347 7.3702
R455 VTAIL.n352 VTAIL.n351 7.3702
R456 VTAIL.n54 VTAIL.n53 7.3702
R457 VTAIL.n58 VTAIL.n57 7.3702
R458 VTAIL.n259 VTAIL.n258 7.3702
R459 VTAIL.n255 VTAIL.n254 7.3702
R460 VTAIL.n161 VTAIL.n160 7.3702
R461 VTAIL.n157 VTAIL.n156 7.3702
R462 VTAIL.n348 VTAIL.n314 6.59444
R463 VTAIL.n351 VTAIL.n314 6.59444
R464 VTAIL.n54 VTAIL.n20 6.59444
R465 VTAIL.n57 VTAIL.n20 6.59444
R466 VTAIL.n258 VTAIL.n221 6.59444
R467 VTAIL.n255 VTAIL.n221 6.59444
R468 VTAIL.n160 VTAIL.n123 6.59444
R469 VTAIL.n157 VTAIL.n123 6.59444
R470 VTAIL.n347 VTAIL.n316 5.81868
R471 VTAIL.n352 VTAIL.n312 5.81868
R472 VTAIL.n53 VTAIL.n22 5.81868
R473 VTAIL.n58 VTAIL.n18 5.81868
R474 VTAIL.n259 VTAIL.n219 5.81868
R475 VTAIL.n254 VTAIL.n223 5.81868
R476 VTAIL.n161 VTAIL.n121 5.81868
R477 VTAIL.n156 VTAIL.n125 5.81868
R478 VTAIL.n344 VTAIL.n343 5.04292
R479 VTAIL.n356 VTAIL.n355 5.04292
R480 VTAIL.n50 VTAIL.n49 5.04292
R481 VTAIL.n62 VTAIL.n61 5.04292
R482 VTAIL.n263 VTAIL.n262 5.04292
R483 VTAIL.n251 VTAIL.n250 5.04292
R484 VTAIL.n165 VTAIL.n164 5.04292
R485 VTAIL.n153 VTAIL.n152 5.04292
R486 VTAIL.n340 VTAIL.n318 4.26717
R487 VTAIL.n359 VTAIL.n310 4.26717
R488 VTAIL.n388 VTAIL.n296 4.26717
R489 VTAIL.n46 VTAIL.n24 4.26717
R490 VTAIL.n65 VTAIL.n16 4.26717
R491 VTAIL.n94 VTAIL.n2 4.26717
R492 VTAIL.n294 VTAIL.n202 4.26717
R493 VTAIL.n266 VTAIL.n217 4.26717
R494 VTAIL.n247 VTAIL.n225 4.26717
R495 VTAIL.n196 VTAIL.n104 4.26717
R496 VTAIL.n168 VTAIL.n119 4.26717
R497 VTAIL.n149 VTAIL.n127 4.26717
R498 VTAIL.n329 VTAIL.n325 3.70982
R499 VTAIL.n35 VTAIL.n31 3.70982
R500 VTAIL.n236 VTAIL.n232 3.70982
R501 VTAIL.n138 VTAIL.n134 3.70982
R502 VTAIL.n339 VTAIL.n320 3.49141
R503 VTAIL.n360 VTAIL.n308 3.49141
R504 VTAIL.n386 VTAIL.n385 3.49141
R505 VTAIL.n45 VTAIL.n26 3.49141
R506 VTAIL.n66 VTAIL.n14 3.49141
R507 VTAIL.n92 VTAIL.n91 3.49141
R508 VTAIL.n292 VTAIL.n291 3.49141
R509 VTAIL.n267 VTAIL.n215 3.49141
R510 VTAIL.n246 VTAIL.n227 3.49141
R511 VTAIL.n194 VTAIL.n193 3.49141
R512 VTAIL.n169 VTAIL.n117 3.49141
R513 VTAIL.n148 VTAIL.n129 3.49141
R514 VTAIL.n336 VTAIL.n335 2.71565
R515 VTAIL.n364 VTAIL.n363 2.71565
R516 VTAIL.n382 VTAIL.n298 2.71565
R517 VTAIL.n42 VTAIL.n41 2.71565
R518 VTAIL.n70 VTAIL.n69 2.71565
R519 VTAIL.n88 VTAIL.n4 2.71565
R520 VTAIL.n288 VTAIL.n204 2.71565
R521 VTAIL.n271 VTAIL.n270 2.71565
R522 VTAIL.n243 VTAIL.n242 2.71565
R523 VTAIL.n190 VTAIL.n106 2.71565
R524 VTAIL.n173 VTAIL.n172 2.71565
R525 VTAIL.n145 VTAIL.n144 2.71565
R526 VTAIL.n332 VTAIL.n322 1.93989
R527 VTAIL.n368 VTAIL.n306 1.93989
R528 VTAIL.n381 VTAIL.n300 1.93989
R529 VTAIL.n38 VTAIL.n28 1.93989
R530 VTAIL.n74 VTAIL.n12 1.93989
R531 VTAIL.n87 VTAIL.n6 1.93989
R532 VTAIL.n287 VTAIL.n206 1.93989
R533 VTAIL.n274 VTAIL.n212 1.93989
R534 VTAIL.n239 VTAIL.n229 1.93989
R535 VTAIL.n189 VTAIL.n108 1.93989
R536 VTAIL.n176 VTAIL.n114 1.93989
R537 VTAIL.n141 VTAIL.n131 1.93989
R538 VTAIL.n390 VTAIL.t9 1.91933
R539 VTAIL.n390 VTAIL.t13 1.91933
R540 VTAIL.n0 VTAIL.t12 1.91933
R541 VTAIL.n0 VTAIL.t8 1.91933
R542 VTAIL.n96 VTAIL.t5 1.91933
R543 VTAIL.n96 VTAIL.t19 1.91933
R544 VTAIL.n98 VTAIL.t3 1.91933
R545 VTAIL.n98 VTAIL.t18 1.91933
R546 VTAIL.n200 VTAIL.t1 1.91933
R547 VTAIL.n200 VTAIL.t2 1.91933
R548 VTAIL.n198 VTAIL.t0 1.91933
R549 VTAIL.n198 VTAIL.t7 1.91933
R550 VTAIL.n102 VTAIL.t11 1.91933
R551 VTAIL.n102 VTAIL.t10 1.91933
R552 VTAIL.n100 VTAIL.t17 1.91933
R553 VTAIL.n100 VTAIL.t14 1.91933
R554 VTAIL.n103 VTAIL.n101 1.31084
R555 VTAIL.n197 VTAIL.n103 1.31084
R556 VTAIL.n201 VTAIL.n199 1.31084
R557 VTAIL.n295 VTAIL.n201 1.31084
R558 VTAIL.n99 VTAIL.n97 1.31084
R559 VTAIL.n97 VTAIL.n95 1.31084
R560 VTAIL.n391 VTAIL.n389 1.31084
R561 VTAIL.n331 VTAIL.n324 1.16414
R562 VTAIL.n369 VTAIL.n304 1.16414
R563 VTAIL.n378 VTAIL.n377 1.16414
R564 VTAIL.n37 VTAIL.n30 1.16414
R565 VTAIL.n75 VTAIL.n10 1.16414
R566 VTAIL.n84 VTAIL.n83 1.16414
R567 VTAIL.n284 VTAIL.n283 1.16414
R568 VTAIL.n275 VTAIL.n210 1.16414
R569 VTAIL.n238 VTAIL.n231 1.16414
R570 VTAIL.n186 VTAIL.n185 1.16414
R571 VTAIL.n177 VTAIL.n112 1.16414
R572 VTAIL.n140 VTAIL.n133 1.16414
R573 VTAIL.n199 VTAIL.n197 1.1255
R574 VTAIL.n95 VTAIL.n1 1.1255
R575 VTAIL VTAIL.n1 1.04145
R576 VTAIL.n328 VTAIL.n327 0.388379
R577 VTAIL.n373 VTAIL.n372 0.388379
R578 VTAIL.n374 VTAIL.n302 0.388379
R579 VTAIL.n34 VTAIL.n33 0.388379
R580 VTAIL.n79 VTAIL.n78 0.388379
R581 VTAIL.n80 VTAIL.n8 0.388379
R582 VTAIL.n280 VTAIL.n208 0.388379
R583 VTAIL.n279 VTAIL.n278 0.388379
R584 VTAIL.n235 VTAIL.n234 0.388379
R585 VTAIL.n182 VTAIL.n110 0.388379
R586 VTAIL.n181 VTAIL.n180 0.388379
R587 VTAIL.n137 VTAIL.n136 0.388379
R588 VTAIL VTAIL.n391 0.269897
R589 VTAIL.n330 VTAIL.n329 0.155672
R590 VTAIL.n330 VTAIL.n321 0.155672
R591 VTAIL.n337 VTAIL.n321 0.155672
R592 VTAIL.n338 VTAIL.n337 0.155672
R593 VTAIL.n338 VTAIL.n317 0.155672
R594 VTAIL.n345 VTAIL.n317 0.155672
R595 VTAIL.n346 VTAIL.n345 0.155672
R596 VTAIL.n346 VTAIL.n313 0.155672
R597 VTAIL.n353 VTAIL.n313 0.155672
R598 VTAIL.n354 VTAIL.n353 0.155672
R599 VTAIL.n354 VTAIL.n309 0.155672
R600 VTAIL.n361 VTAIL.n309 0.155672
R601 VTAIL.n362 VTAIL.n361 0.155672
R602 VTAIL.n362 VTAIL.n305 0.155672
R603 VTAIL.n370 VTAIL.n305 0.155672
R604 VTAIL.n371 VTAIL.n370 0.155672
R605 VTAIL.n371 VTAIL.n301 0.155672
R606 VTAIL.n379 VTAIL.n301 0.155672
R607 VTAIL.n380 VTAIL.n379 0.155672
R608 VTAIL.n380 VTAIL.n297 0.155672
R609 VTAIL.n387 VTAIL.n297 0.155672
R610 VTAIL.n36 VTAIL.n35 0.155672
R611 VTAIL.n36 VTAIL.n27 0.155672
R612 VTAIL.n43 VTAIL.n27 0.155672
R613 VTAIL.n44 VTAIL.n43 0.155672
R614 VTAIL.n44 VTAIL.n23 0.155672
R615 VTAIL.n51 VTAIL.n23 0.155672
R616 VTAIL.n52 VTAIL.n51 0.155672
R617 VTAIL.n52 VTAIL.n19 0.155672
R618 VTAIL.n59 VTAIL.n19 0.155672
R619 VTAIL.n60 VTAIL.n59 0.155672
R620 VTAIL.n60 VTAIL.n15 0.155672
R621 VTAIL.n67 VTAIL.n15 0.155672
R622 VTAIL.n68 VTAIL.n67 0.155672
R623 VTAIL.n68 VTAIL.n11 0.155672
R624 VTAIL.n76 VTAIL.n11 0.155672
R625 VTAIL.n77 VTAIL.n76 0.155672
R626 VTAIL.n77 VTAIL.n7 0.155672
R627 VTAIL.n85 VTAIL.n7 0.155672
R628 VTAIL.n86 VTAIL.n85 0.155672
R629 VTAIL.n86 VTAIL.n3 0.155672
R630 VTAIL.n93 VTAIL.n3 0.155672
R631 VTAIL.n293 VTAIL.n203 0.155672
R632 VTAIL.n286 VTAIL.n203 0.155672
R633 VTAIL.n286 VTAIL.n285 0.155672
R634 VTAIL.n285 VTAIL.n207 0.155672
R635 VTAIL.n277 VTAIL.n207 0.155672
R636 VTAIL.n277 VTAIL.n276 0.155672
R637 VTAIL.n276 VTAIL.n211 0.155672
R638 VTAIL.n269 VTAIL.n211 0.155672
R639 VTAIL.n269 VTAIL.n268 0.155672
R640 VTAIL.n268 VTAIL.n216 0.155672
R641 VTAIL.n261 VTAIL.n216 0.155672
R642 VTAIL.n261 VTAIL.n260 0.155672
R643 VTAIL.n260 VTAIL.n220 0.155672
R644 VTAIL.n253 VTAIL.n220 0.155672
R645 VTAIL.n253 VTAIL.n252 0.155672
R646 VTAIL.n252 VTAIL.n224 0.155672
R647 VTAIL.n245 VTAIL.n224 0.155672
R648 VTAIL.n245 VTAIL.n244 0.155672
R649 VTAIL.n244 VTAIL.n228 0.155672
R650 VTAIL.n237 VTAIL.n228 0.155672
R651 VTAIL.n237 VTAIL.n236 0.155672
R652 VTAIL.n195 VTAIL.n105 0.155672
R653 VTAIL.n188 VTAIL.n105 0.155672
R654 VTAIL.n188 VTAIL.n187 0.155672
R655 VTAIL.n187 VTAIL.n109 0.155672
R656 VTAIL.n179 VTAIL.n109 0.155672
R657 VTAIL.n179 VTAIL.n178 0.155672
R658 VTAIL.n178 VTAIL.n113 0.155672
R659 VTAIL.n171 VTAIL.n113 0.155672
R660 VTAIL.n171 VTAIL.n170 0.155672
R661 VTAIL.n170 VTAIL.n118 0.155672
R662 VTAIL.n163 VTAIL.n118 0.155672
R663 VTAIL.n163 VTAIL.n162 0.155672
R664 VTAIL.n162 VTAIL.n122 0.155672
R665 VTAIL.n155 VTAIL.n122 0.155672
R666 VTAIL.n155 VTAIL.n154 0.155672
R667 VTAIL.n154 VTAIL.n126 0.155672
R668 VTAIL.n147 VTAIL.n126 0.155672
R669 VTAIL.n147 VTAIL.n146 0.155672
R670 VTAIL.n146 VTAIL.n130 0.155672
R671 VTAIL.n139 VTAIL.n130 0.155672
R672 VTAIL.n139 VTAIL.n138 0.155672
R673 VDD2.n185 VDD2.n97 756.745
R674 VDD2.n88 VDD2.n0 756.745
R675 VDD2.n186 VDD2.n185 585
R676 VDD2.n184 VDD2.n183 585
R677 VDD2.n101 VDD2.n100 585
R678 VDD2.n178 VDD2.n177 585
R679 VDD2.n176 VDD2.n175 585
R680 VDD2.n174 VDD2.n104 585
R681 VDD2.n108 VDD2.n105 585
R682 VDD2.n169 VDD2.n168 585
R683 VDD2.n167 VDD2.n166 585
R684 VDD2.n110 VDD2.n109 585
R685 VDD2.n161 VDD2.n160 585
R686 VDD2.n159 VDD2.n158 585
R687 VDD2.n114 VDD2.n113 585
R688 VDD2.n153 VDD2.n152 585
R689 VDD2.n151 VDD2.n150 585
R690 VDD2.n118 VDD2.n117 585
R691 VDD2.n145 VDD2.n144 585
R692 VDD2.n143 VDD2.n142 585
R693 VDD2.n122 VDD2.n121 585
R694 VDD2.n137 VDD2.n136 585
R695 VDD2.n135 VDD2.n134 585
R696 VDD2.n126 VDD2.n125 585
R697 VDD2.n129 VDD2.n128 585
R698 VDD2.n31 VDD2.n30 585
R699 VDD2.n28 VDD2.n27 585
R700 VDD2.n37 VDD2.n36 585
R701 VDD2.n39 VDD2.n38 585
R702 VDD2.n24 VDD2.n23 585
R703 VDD2.n45 VDD2.n44 585
R704 VDD2.n47 VDD2.n46 585
R705 VDD2.n20 VDD2.n19 585
R706 VDD2.n53 VDD2.n52 585
R707 VDD2.n55 VDD2.n54 585
R708 VDD2.n16 VDD2.n15 585
R709 VDD2.n61 VDD2.n60 585
R710 VDD2.n63 VDD2.n62 585
R711 VDD2.n12 VDD2.n11 585
R712 VDD2.n69 VDD2.n68 585
R713 VDD2.n72 VDD2.n71 585
R714 VDD2.n70 VDD2.n8 585
R715 VDD2.n77 VDD2.n7 585
R716 VDD2.n79 VDD2.n78 585
R717 VDD2.n81 VDD2.n80 585
R718 VDD2.n4 VDD2.n3 585
R719 VDD2.n87 VDD2.n86 585
R720 VDD2.n89 VDD2.n88 585
R721 VDD2.t2 VDD2.n127 327.466
R722 VDD2.t6 VDD2.n29 327.466
R723 VDD2.n185 VDD2.n184 171.744
R724 VDD2.n184 VDD2.n100 171.744
R725 VDD2.n177 VDD2.n100 171.744
R726 VDD2.n177 VDD2.n176 171.744
R727 VDD2.n176 VDD2.n104 171.744
R728 VDD2.n108 VDD2.n104 171.744
R729 VDD2.n168 VDD2.n108 171.744
R730 VDD2.n168 VDD2.n167 171.744
R731 VDD2.n167 VDD2.n109 171.744
R732 VDD2.n160 VDD2.n109 171.744
R733 VDD2.n160 VDD2.n159 171.744
R734 VDD2.n159 VDD2.n113 171.744
R735 VDD2.n152 VDD2.n113 171.744
R736 VDD2.n152 VDD2.n151 171.744
R737 VDD2.n151 VDD2.n117 171.744
R738 VDD2.n144 VDD2.n117 171.744
R739 VDD2.n144 VDD2.n143 171.744
R740 VDD2.n143 VDD2.n121 171.744
R741 VDD2.n136 VDD2.n121 171.744
R742 VDD2.n136 VDD2.n135 171.744
R743 VDD2.n135 VDD2.n125 171.744
R744 VDD2.n128 VDD2.n125 171.744
R745 VDD2.n30 VDD2.n27 171.744
R746 VDD2.n37 VDD2.n27 171.744
R747 VDD2.n38 VDD2.n37 171.744
R748 VDD2.n38 VDD2.n23 171.744
R749 VDD2.n45 VDD2.n23 171.744
R750 VDD2.n46 VDD2.n45 171.744
R751 VDD2.n46 VDD2.n19 171.744
R752 VDD2.n53 VDD2.n19 171.744
R753 VDD2.n54 VDD2.n53 171.744
R754 VDD2.n54 VDD2.n15 171.744
R755 VDD2.n61 VDD2.n15 171.744
R756 VDD2.n62 VDD2.n61 171.744
R757 VDD2.n62 VDD2.n11 171.744
R758 VDD2.n69 VDD2.n11 171.744
R759 VDD2.n71 VDD2.n69 171.744
R760 VDD2.n71 VDD2.n70 171.744
R761 VDD2.n70 VDD2.n7 171.744
R762 VDD2.n79 VDD2.n7 171.744
R763 VDD2.n80 VDD2.n79 171.744
R764 VDD2.n80 VDD2.n3 171.744
R765 VDD2.n87 VDD2.n3 171.744
R766 VDD2.n88 VDD2.n87 171.744
R767 VDD2.n128 VDD2.t2 85.8723
R768 VDD2.n30 VDD2.t6 85.8723
R769 VDD2.n96 VDD2.n95 73.0344
R770 VDD2 VDD2.n193 73.0316
R771 VDD2.n192 VDD2.n191 72.1072
R772 VDD2.n94 VDD2.n93 72.107
R773 VDD2.n94 VDD2.n92 52.8896
R774 VDD2.n190 VDD2.n189 51.5793
R775 VDD2.n190 VDD2.n96 44.5429
R776 VDD2.n129 VDD2.n127 16.3895
R777 VDD2.n31 VDD2.n29 16.3895
R778 VDD2.n175 VDD2.n174 13.1884
R779 VDD2.n78 VDD2.n77 13.1884
R780 VDD2.n178 VDD2.n103 12.8005
R781 VDD2.n173 VDD2.n105 12.8005
R782 VDD2.n130 VDD2.n126 12.8005
R783 VDD2.n32 VDD2.n28 12.8005
R784 VDD2.n76 VDD2.n8 12.8005
R785 VDD2.n81 VDD2.n6 12.8005
R786 VDD2.n179 VDD2.n101 12.0247
R787 VDD2.n170 VDD2.n169 12.0247
R788 VDD2.n134 VDD2.n133 12.0247
R789 VDD2.n36 VDD2.n35 12.0247
R790 VDD2.n73 VDD2.n72 12.0247
R791 VDD2.n82 VDD2.n4 12.0247
R792 VDD2.n183 VDD2.n182 11.249
R793 VDD2.n166 VDD2.n107 11.249
R794 VDD2.n137 VDD2.n124 11.249
R795 VDD2.n39 VDD2.n26 11.249
R796 VDD2.n68 VDD2.n10 11.249
R797 VDD2.n86 VDD2.n85 11.249
R798 VDD2.n186 VDD2.n99 10.4732
R799 VDD2.n165 VDD2.n110 10.4732
R800 VDD2.n138 VDD2.n122 10.4732
R801 VDD2.n40 VDD2.n24 10.4732
R802 VDD2.n67 VDD2.n12 10.4732
R803 VDD2.n89 VDD2.n2 10.4732
R804 VDD2.n187 VDD2.n97 9.69747
R805 VDD2.n162 VDD2.n161 9.69747
R806 VDD2.n142 VDD2.n141 9.69747
R807 VDD2.n44 VDD2.n43 9.69747
R808 VDD2.n64 VDD2.n63 9.69747
R809 VDD2.n90 VDD2.n0 9.69747
R810 VDD2.n189 VDD2.n188 9.45567
R811 VDD2.n92 VDD2.n91 9.45567
R812 VDD2.n155 VDD2.n154 9.3005
R813 VDD2.n157 VDD2.n156 9.3005
R814 VDD2.n112 VDD2.n111 9.3005
R815 VDD2.n163 VDD2.n162 9.3005
R816 VDD2.n165 VDD2.n164 9.3005
R817 VDD2.n107 VDD2.n106 9.3005
R818 VDD2.n171 VDD2.n170 9.3005
R819 VDD2.n173 VDD2.n172 9.3005
R820 VDD2.n188 VDD2.n187 9.3005
R821 VDD2.n99 VDD2.n98 9.3005
R822 VDD2.n182 VDD2.n181 9.3005
R823 VDD2.n180 VDD2.n179 9.3005
R824 VDD2.n103 VDD2.n102 9.3005
R825 VDD2.n116 VDD2.n115 9.3005
R826 VDD2.n149 VDD2.n148 9.3005
R827 VDD2.n147 VDD2.n146 9.3005
R828 VDD2.n120 VDD2.n119 9.3005
R829 VDD2.n141 VDD2.n140 9.3005
R830 VDD2.n139 VDD2.n138 9.3005
R831 VDD2.n124 VDD2.n123 9.3005
R832 VDD2.n133 VDD2.n132 9.3005
R833 VDD2.n131 VDD2.n130 9.3005
R834 VDD2.n91 VDD2.n90 9.3005
R835 VDD2.n2 VDD2.n1 9.3005
R836 VDD2.n85 VDD2.n84 9.3005
R837 VDD2.n83 VDD2.n82 9.3005
R838 VDD2.n6 VDD2.n5 9.3005
R839 VDD2.n51 VDD2.n50 9.3005
R840 VDD2.n49 VDD2.n48 9.3005
R841 VDD2.n22 VDD2.n21 9.3005
R842 VDD2.n43 VDD2.n42 9.3005
R843 VDD2.n41 VDD2.n40 9.3005
R844 VDD2.n26 VDD2.n25 9.3005
R845 VDD2.n35 VDD2.n34 9.3005
R846 VDD2.n33 VDD2.n32 9.3005
R847 VDD2.n18 VDD2.n17 9.3005
R848 VDD2.n57 VDD2.n56 9.3005
R849 VDD2.n59 VDD2.n58 9.3005
R850 VDD2.n14 VDD2.n13 9.3005
R851 VDD2.n65 VDD2.n64 9.3005
R852 VDD2.n67 VDD2.n66 9.3005
R853 VDD2.n10 VDD2.n9 9.3005
R854 VDD2.n74 VDD2.n73 9.3005
R855 VDD2.n76 VDD2.n75 9.3005
R856 VDD2.n158 VDD2.n112 8.92171
R857 VDD2.n145 VDD2.n120 8.92171
R858 VDD2.n47 VDD2.n22 8.92171
R859 VDD2.n60 VDD2.n14 8.92171
R860 VDD2.n157 VDD2.n114 8.14595
R861 VDD2.n146 VDD2.n118 8.14595
R862 VDD2.n48 VDD2.n20 8.14595
R863 VDD2.n59 VDD2.n16 8.14595
R864 VDD2.n154 VDD2.n153 7.3702
R865 VDD2.n150 VDD2.n149 7.3702
R866 VDD2.n52 VDD2.n51 7.3702
R867 VDD2.n56 VDD2.n55 7.3702
R868 VDD2.n153 VDD2.n116 6.59444
R869 VDD2.n150 VDD2.n116 6.59444
R870 VDD2.n52 VDD2.n18 6.59444
R871 VDD2.n55 VDD2.n18 6.59444
R872 VDD2.n154 VDD2.n114 5.81868
R873 VDD2.n149 VDD2.n118 5.81868
R874 VDD2.n51 VDD2.n20 5.81868
R875 VDD2.n56 VDD2.n16 5.81868
R876 VDD2.n158 VDD2.n157 5.04292
R877 VDD2.n146 VDD2.n145 5.04292
R878 VDD2.n48 VDD2.n47 5.04292
R879 VDD2.n60 VDD2.n59 5.04292
R880 VDD2.n189 VDD2.n97 4.26717
R881 VDD2.n161 VDD2.n112 4.26717
R882 VDD2.n142 VDD2.n120 4.26717
R883 VDD2.n44 VDD2.n22 4.26717
R884 VDD2.n63 VDD2.n14 4.26717
R885 VDD2.n92 VDD2.n0 4.26717
R886 VDD2.n131 VDD2.n127 3.70982
R887 VDD2.n33 VDD2.n29 3.70982
R888 VDD2.n187 VDD2.n186 3.49141
R889 VDD2.n162 VDD2.n110 3.49141
R890 VDD2.n141 VDD2.n122 3.49141
R891 VDD2.n43 VDD2.n24 3.49141
R892 VDD2.n64 VDD2.n12 3.49141
R893 VDD2.n90 VDD2.n89 3.49141
R894 VDD2.n183 VDD2.n99 2.71565
R895 VDD2.n166 VDD2.n165 2.71565
R896 VDD2.n138 VDD2.n137 2.71565
R897 VDD2.n40 VDD2.n39 2.71565
R898 VDD2.n68 VDD2.n67 2.71565
R899 VDD2.n86 VDD2.n2 2.71565
R900 VDD2.n182 VDD2.n101 1.93989
R901 VDD2.n169 VDD2.n107 1.93989
R902 VDD2.n134 VDD2.n124 1.93989
R903 VDD2.n36 VDD2.n26 1.93989
R904 VDD2.n72 VDD2.n10 1.93989
R905 VDD2.n85 VDD2.n4 1.93989
R906 VDD2.n193 VDD2.t7 1.91933
R907 VDD2.n193 VDD2.t4 1.91933
R908 VDD2.n191 VDD2.t0 1.91933
R909 VDD2.n191 VDD2.t9 1.91933
R910 VDD2.n95 VDD2.t5 1.91933
R911 VDD2.n95 VDD2.t1 1.91933
R912 VDD2.n93 VDD2.t3 1.91933
R913 VDD2.n93 VDD2.t8 1.91933
R914 VDD2.n192 VDD2.n190 1.31084
R915 VDD2.n179 VDD2.n178 1.16414
R916 VDD2.n170 VDD2.n105 1.16414
R917 VDD2.n133 VDD2.n126 1.16414
R918 VDD2.n35 VDD2.n28 1.16414
R919 VDD2.n73 VDD2.n8 1.16414
R920 VDD2.n82 VDD2.n81 1.16414
R921 VDD2.n175 VDD2.n103 0.388379
R922 VDD2.n174 VDD2.n173 0.388379
R923 VDD2.n130 VDD2.n129 0.388379
R924 VDD2.n32 VDD2.n31 0.388379
R925 VDD2.n77 VDD2.n76 0.388379
R926 VDD2.n78 VDD2.n6 0.388379
R927 VDD2 VDD2.n192 0.386276
R928 VDD2.n96 VDD2.n94 0.27274
R929 VDD2.n188 VDD2.n98 0.155672
R930 VDD2.n181 VDD2.n98 0.155672
R931 VDD2.n181 VDD2.n180 0.155672
R932 VDD2.n180 VDD2.n102 0.155672
R933 VDD2.n172 VDD2.n102 0.155672
R934 VDD2.n172 VDD2.n171 0.155672
R935 VDD2.n171 VDD2.n106 0.155672
R936 VDD2.n164 VDD2.n106 0.155672
R937 VDD2.n164 VDD2.n163 0.155672
R938 VDD2.n163 VDD2.n111 0.155672
R939 VDD2.n156 VDD2.n111 0.155672
R940 VDD2.n156 VDD2.n155 0.155672
R941 VDD2.n155 VDD2.n115 0.155672
R942 VDD2.n148 VDD2.n115 0.155672
R943 VDD2.n148 VDD2.n147 0.155672
R944 VDD2.n147 VDD2.n119 0.155672
R945 VDD2.n140 VDD2.n119 0.155672
R946 VDD2.n140 VDD2.n139 0.155672
R947 VDD2.n139 VDD2.n123 0.155672
R948 VDD2.n132 VDD2.n123 0.155672
R949 VDD2.n132 VDD2.n131 0.155672
R950 VDD2.n34 VDD2.n33 0.155672
R951 VDD2.n34 VDD2.n25 0.155672
R952 VDD2.n41 VDD2.n25 0.155672
R953 VDD2.n42 VDD2.n41 0.155672
R954 VDD2.n42 VDD2.n21 0.155672
R955 VDD2.n49 VDD2.n21 0.155672
R956 VDD2.n50 VDD2.n49 0.155672
R957 VDD2.n50 VDD2.n17 0.155672
R958 VDD2.n57 VDD2.n17 0.155672
R959 VDD2.n58 VDD2.n57 0.155672
R960 VDD2.n58 VDD2.n13 0.155672
R961 VDD2.n65 VDD2.n13 0.155672
R962 VDD2.n66 VDD2.n65 0.155672
R963 VDD2.n66 VDD2.n9 0.155672
R964 VDD2.n74 VDD2.n9 0.155672
R965 VDD2.n75 VDD2.n74 0.155672
R966 VDD2.n75 VDD2.n5 0.155672
R967 VDD2.n83 VDD2.n5 0.155672
R968 VDD2.n84 VDD2.n83 0.155672
R969 VDD2.n84 VDD2.n1 0.155672
R970 VDD2.n91 VDD2.n1 0.155672
R971 B.n546 B.n85 585
R972 B.n548 B.n547 585
R973 B.n549 B.n84 585
R974 B.n551 B.n550 585
R975 B.n552 B.n83 585
R976 B.n554 B.n553 585
R977 B.n555 B.n82 585
R978 B.n557 B.n556 585
R979 B.n558 B.n81 585
R980 B.n560 B.n559 585
R981 B.n561 B.n80 585
R982 B.n563 B.n562 585
R983 B.n564 B.n79 585
R984 B.n566 B.n565 585
R985 B.n567 B.n78 585
R986 B.n569 B.n568 585
R987 B.n570 B.n77 585
R988 B.n572 B.n571 585
R989 B.n573 B.n76 585
R990 B.n575 B.n574 585
R991 B.n576 B.n75 585
R992 B.n578 B.n577 585
R993 B.n579 B.n74 585
R994 B.n581 B.n580 585
R995 B.n582 B.n73 585
R996 B.n584 B.n583 585
R997 B.n585 B.n72 585
R998 B.n587 B.n586 585
R999 B.n588 B.n71 585
R1000 B.n590 B.n589 585
R1001 B.n591 B.n70 585
R1002 B.n593 B.n592 585
R1003 B.n594 B.n69 585
R1004 B.n596 B.n595 585
R1005 B.n597 B.n68 585
R1006 B.n599 B.n598 585
R1007 B.n600 B.n67 585
R1008 B.n602 B.n601 585
R1009 B.n603 B.n66 585
R1010 B.n605 B.n604 585
R1011 B.n606 B.n65 585
R1012 B.n608 B.n607 585
R1013 B.n609 B.n64 585
R1014 B.n611 B.n610 585
R1015 B.n612 B.n63 585
R1016 B.n614 B.n613 585
R1017 B.n615 B.n62 585
R1018 B.n617 B.n616 585
R1019 B.n618 B.n61 585
R1020 B.n620 B.n619 585
R1021 B.n621 B.n60 585
R1022 B.n623 B.n622 585
R1023 B.n624 B.n59 585
R1024 B.n626 B.n625 585
R1025 B.n627 B.n55 585
R1026 B.n629 B.n628 585
R1027 B.n630 B.n54 585
R1028 B.n632 B.n631 585
R1029 B.n633 B.n53 585
R1030 B.n635 B.n634 585
R1031 B.n636 B.n52 585
R1032 B.n638 B.n637 585
R1033 B.n639 B.n51 585
R1034 B.n641 B.n640 585
R1035 B.n642 B.n50 585
R1036 B.n644 B.n643 585
R1037 B.n646 B.n47 585
R1038 B.n648 B.n647 585
R1039 B.n649 B.n46 585
R1040 B.n651 B.n650 585
R1041 B.n652 B.n45 585
R1042 B.n654 B.n653 585
R1043 B.n655 B.n44 585
R1044 B.n657 B.n656 585
R1045 B.n658 B.n43 585
R1046 B.n660 B.n659 585
R1047 B.n661 B.n42 585
R1048 B.n663 B.n662 585
R1049 B.n664 B.n41 585
R1050 B.n666 B.n665 585
R1051 B.n667 B.n40 585
R1052 B.n669 B.n668 585
R1053 B.n670 B.n39 585
R1054 B.n672 B.n671 585
R1055 B.n673 B.n38 585
R1056 B.n675 B.n674 585
R1057 B.n676 B.n37 585
R1058 B.n678 B.n677 585
R1059 B.n679 B.n36 585
R1060 B.n681 B.n680 585
R1061 B.n682 B.n35 585
R1062 B.n684 B.n683 585
R1063 B.n685 B.n34 585
R1064 B.n687 B.n686 585
R1065 B.n688 B.n33 585
R1066 B.n690 B.n689 585
R1067 B.n691 B.n32 585
R1068 B.n693 B.n692 585
R1069 B.n694 B.n31 585
R1070 B.n696 B.n695 585
R1071 B.n697 B.n30 585
R1072 B.n699 B.n698 585
R1073 B.n700 B.n29 585
R1074 B.n702 B.n701 585
R1075 B.n703 B.n28 585
R1076 B.n705 B.n704 585
R1077 B.n706 B.n27 585
R1078 B.n708 B.n707 585
R1079 B.n709 B.n26 585
R1080 B.n711 B.n710 585
R1081 B.n712 B.n25 585
R1082 B.n714 B.n713 585
R1083 B.n715 B.n24 585
R1084 B.n717 B.n716 585
R1085 B.n718 B.n23 585
R1086 B.n720 B.n719 585
R1087 B.n721 B.n22 585
R1088 B.n723 B.n722 585
R1089 B.n724 B.n21 585
R1090 B.n726 B.n725 585
R1091 B.n727 B.n20 585
R1092 B.n729 B.n728 585
R1093 B.n545 B.n544 585
R1094 B.n543 B.n86 585
R1095 B.n542 B.n541 585
R1096 B.n540 B.n87 585
R1097 B.n539 B.n538 585
R1098 B.n537 B.n88 585
R1099 B.n536 B.n535 585
R1100 B.n534 B.n89 585
R1101 B.n533 B.n532 585
R1102 B.n531 B.n90 585
R1103 B.n530 B.n529 585
R1104 B.n528 B.n91 585
R1105 B.n527 B.n526 585
R1106 B.n525 B.n92 585
R1107 B.n524 B.n523 585
R1108 B.n522 B.n93 585
R1109 B.n521 B.n520 585
R1110 B.n519 B.n94 585
R1111 B.n518 B.n517 585
R1112 B.n516 B.n95 585
R1113 B.n515 B.n514 585
R1114 B.n513 B.n96 585
R1115 B.n512 B.n511 585
R1116 B.n510 B.n97 585
R1117 B.n509 B.n508 585
R1118 B.n507 B.n98 585
R1119 B.n506 B.n505 585
R1120 B.n504 B.n99 585
R1121 B.n503 B.n502 585
R1122 B.n501 B.n100 585
R1123 B.n500 B.n499 585
R1124 B.n498 B.n101 585
R1125 B.n497 B.n496 585
R1126 B.n495 B.n102 585
R1127 B.n494 B.n493 585
R1128 B.n492 B.n103 585
R1129 B.n491 B.n490 585
R1130 B.n489 B.n104 585
R1131 B.n488 B.n487 585
R1132 B.n486 B.n105 585
R1133 B.n485 B.n484 585
R1134 B.n483 B.n106 585
R1135 B.n482 B.n481 585
R1136 B.n480 B.n107 585
R1137 B.n479 B.n478 585
R1138 B.n477 B.n108 585
R1139 B.n476 B.n475 585
R1140 B.n474 B.n109 585
R1141 B.n473 B.n472 585
R1142 B.n471 B.n110 585
R1143 B.n470 B.n469 585
R1144 B.n468 B.n111 585
R1145 B.n467 B.n466 585
R1146 B.n465 B.n112 585
R1147 B.n464 B.n463 585
R1148 B.n462 B.n113 585
R1149 B.n461 B.n460 585
R1150 B.n459 B.n114 585
R1151 B.n458 B.n457 585
R1152 B.n456 B.n115 585
R1153 B.n455 B.n454 585
R1154 B.n453 B.n116 585
R1155 B.n452 B.n451 585
R1156 B.n450 B.n117 585
R1157 B.n449 B.n448 585
R1158 B.n447 B.n118 585
R1159 B.n446 B.n445 585
R1160 B.n444 B.n119 585
R1161 B.n443 B.n442 585
R1162 B.n441 B.n120 585
R1163 B.n440 B.n439 585
R1164 B.n255 B.n186 585
R1165 B.n257 B.n256 585
R1166 B.n258 B.n185 585
R1167 B.n260 B.n259 585
R1168 B.n261 B.n184 585
R1169 B.n263 B.n262 585
R1170 B.n264 B.n183 585
R1171 B.n266 B.n265 585
R1172 B.n267 B.n182 585
R1173 B.n269 B.n268 585
R1174 B.n270 B.n181 585
R1175 B.n272 B.n271 585
R1176 B.n273 B.n180 585
R1177 B.n275 B.n274 585
R1178 B.n276 B.n179 585
R1179 B.n278 B.n277 585
R1180 B.n279 B.n178 585
R1181 B.n281 B.n280 585
R1182 B.n282 B.n177 585
R1183 B.n284 B.n283 585
R1184 B.n285 B.n176 585
R1185 B.n287 B.n286 585
R1186 B.n288 B.n175 585
R1187 B.n290 B.n289 585
R1188 B.n291 B.n174 585
R1189 B.n293 B.n292 585
R1190 B.n294 B.n173 585
R1191 B.n296 B.n295 585
R1192 B.n297 B.n172 585
R1193 B.n299 B.n298 585
R1194 B.n300 B.n171 585
R1195 B.n302 B.n301 585
R1196 B.n303 B.n170 585
R1197 B.n305 B.n304 585
R1198 B.n306 B.n169 585
R1199 B.n308 B.n307 585
R1200 B.n309 B.n168 585
R1201 B.n311 B.n310 585
R1202 B.n312 B.n167 585
R1203 B.n314 B.n313 585
R1204 B.n315 B.n166 585
R1205 B.n317 B.n316 585
R1206 B.n318 B.n165 585
R1207 B.n320 B.n319 585
R1208 B.n321 B.n164 585
R1209 B.n323 B.n322 585
R1210 B.n324 B.n163 585
R1211 B.n326 B.n325 585
R1212 B.n327 B.n162 585
R1213 B.n329 B.n328 585
R1214 B.n330 B.n161 585
R1215 B.n332 B.n331 585
R1216 B.n333 B.n160 585
R1217 B.n335 B.n334 585
R1218 B.n336 B.n159 585
R1219 B.n338 B.n337 585
R1220 B.n340 B.n156 585
R1221 B.n342 B.n341 585
R1222 B.n343 B.n155 585
R1223 B.n345 B.n344 585
R1224 B.n346 B.n154 585
R1225 B.n348 B.n347 585
R1226 B.n349 B.n153 585
R1227 B.n351 B.n350 585
R1228 B.n352 B.n152 585
R1229 B.n354 B.n353 585
R1230 B.n356 B.n355 585
R1231 B.n357 B.n148 585
R1232 B.n359 B.n358 585
R1233 B.n360 B.n147 585
R1234 B.n362 B.n361 585
R1235 B.n363 B.n146 585
R1236 B.n365 B.n364 585
R1237 B.n366 B.n145 585
R1238 B.n368 B.n367 585
R1239 B.n369 B.n144 585
R1240 B.n371 B.n370 585
R1241 B.n372 B.n143 585
R1242 B.n374 B.n373 585
R1243 B.n375 B.n142 585
R1244 B.n377 B.n376 585
R1245 B.n378 B.n141 585
R1246 B.n380 B.n379 585
R1247 B.n381 B.n140 585
R1248 B.n383 B.n382 585
R1249 B.n384 B.n139 585
R1250 B.n386 B.n385 585
R1251 B.n387 B.n138 585
R1252 B.n389 B.n388 585
R1253 B.n390 B.n137 585
R1254 B.n392 B.n391 585
R1255 B.n393 B.n136 585
R1256 B.n395 B.n394 585
R1257 B.n396 B.n135 585
R1258 B.n398 B.n397 585
R1259 B.n399 B.n134 585
R1260 B.n401 B.n400 585
R1261 B.n402 B.n133 585
R1262 B.n404 B.n403 585
R1263 B.n405 B.n132 585
R1264 B.n407 B.n406 585
R1265 B.n408 B.n131 585
R1266 B.n410 B.n409 585
R1267 B.n411 B.n130 585
R1268 B.n413 B.n412 585
R1269 B.n414 B.n129 585
R1270 B.n416 B.n415 585
R1271 B.n417 B.n128 585
R1272 B.n419 B.n418 585
R1273 B.n420 B.n127 585
R1274 B.n422 B.n421 585
R1275 B.n423 B.n126 585
R1276 B.n425 B.n424 585
R1277 B.n426 B.n125 585
R1278 B.n428 B.n427 585
R1279 B.n429 B.n124 585
R1280 B.n431 B.n430 585
R1281 B.n432 B.n123 585
R1282 B.n434 B.n433 585
R1283 B.n435 B.n122 585
R1284 B.n437 B.n436 585
R1285 B.n438 B.n121 585
R1286 B.n254 B.n253 585
R1287 B.n252 B.n187 585
R1288 B.n251 B.n250 585
R1289 B.n249 B.n188 585
R1290 B.n248 B.n247 585
R1291 B.n246 B.n189 585
R1292 B.n245 B.n244 585
R1293 B.n243 B.n190 585
R1294 B.n242 B.n241 585
R1295 B.n240 B.n191 585
R1296 B.n239 B.n238 585
R1297 B.n237 B.n192 585
R1298 B.n236 B.n235 585
R1299 B.n234 B.n193 585
R1300 B.n233 B.n232 585
R1301 B.n231 B.n194 585
R1302 B.n230 B.n229 585
R1303 B.n228 B.n195 585
R1304 B.n227 B.n226 585
R1305 B.n225 B.n196 585
R1306 B.n224 B.n223 585
R1307 B.n222 B.n197 585
R1308 B.n221 B.n220 585
R1309 B.n219 B.n198 585
R1310 B.n218 B.n217 585
R1311 B.n216 B.n199 585
R1312 B.n215 B.n214 585
R1313 B.n213 B.n200 585
R1314 B.n212 B.n211 585
R1315 B.n210 B.n201 585
R1316 B.n209 B.n208 585
R1317 B.n207 B.n202 585
R1318 B.n206 B.n205 585
R1319 B.n204 B.n203 585
R1320 B.n2 B.n0 585
R1321 B.n781 B.n1 585
R1322 B.n780 B.n779 585
R1323 B.n778 B.n3 585
R1324 B.n777 B.n776 585
R1325 B.n775 B.n4 585
R1326 B.n774 B.n773 585
R1327 B.n772 B.n5 585
R1328 B.n771 B.n770 585
R1329 B.n769 B.n6 585
R1330 B.n768 B.n767 585
R1331 B.n766 B.n7 585
R1332 B.n765 B.n764 585
R1333 B.n763 B.n8 585
R1334 B.n762 B.n761 585
R1335 B.n760 B.n9 585
R1336 B.n759 B.n758 585
R1337 B.n757 B.n10 585
R1338 B.n756 B.n755 585
R1339 B.n754 B.n11 585
R1340 B.n753 B.n752 585
R1341 B.n751 B.n12 585
R1342 B.n750 B.n749 585
R1343 B.n748 B.n13 585
R1344 B.n747 B.n746 585
R1345 B.n745 B.n14 585
R1346 B.n744 B.n743 585
R1347 B.n742 B.n15 585
R1348 B.n741 B.n740 585
R1349 B.n739 B.n16 585
R1350 B.n738 B.n737 585
R1351 B.n736 B.n17 585
R1352 B.n735 B.n734 585
R1353 B.n733 B.n18 585
R1354 B.n732 B.n731 585
R1355 B.n730 B.n19 585
R1356 B.n783 B.n782 585
R1357 B.n149 B.t6 547.135
R1358 B.n157 B.t9 547.135
R1359 B.n48 B.t0 547.135
R1360 B.n56 B.t3 547.135
R1361 B.n149 B.t8 494.235
R1362 B.n56 B.t4 494.235
R1363 B.n157 B.t11 494.235
R1364 B.n48 B.t1 494.235
R1365 B.n253 B.n186 478.086
R1366 B.n728 B.n19 478.086
R1367 B.n439 B.n438 478.086
R1368 B.n546 B.n545 478.086
R1369 B.n150 B.t7 464.755
R1370 B.n57 B.t5 464.755
R1371 B.n158 B.t10 464.755
R1372 B.n49 B.t2 464.755
R1373 B.n253 B.n252 163.367
R1374 B.n252 B.n251 163.367
R1375 B.n251 B.n188 163.367
R1376 B.n247 B.n188 163.367
R1377 B.n247 B.n246 163.367
R1378 B.n246 B.n245 163.367
R1379 B.n245 B.n190 163.367
R1380 B.n241 B.n190 163.367
R1381 B.n241 B.n240 163.367
R1382 B.n240 B.n239 163.367
R1383 B.n239 B.n192 163.367
R1384 B.n235 B.n192 163.367
R1385 B.n235 B.n234 163.367
R1386 B.n234 B.n233 163.367
R1387 B.n233 B.n194 163.367
R1388 B.n229 B.n194 163.367
R1389 B.n229 B.n228 163.367
R1390 B.n228 B.n227 163.367
R1391 B.n227 B.n196 163.367
R1392 B.n223 B.n196 163.367
R1393 B.n223 B.n222 163.367
R1394 B.n222 B.n221 163.367
R1395 B.n221 B.n198 163.367
R1396 B.n217 B.n198 163.367
R1397 B.n217 B.n216 163.367
R1398 B.n216 B.n215 163.367
R1399 B.n215 B.n200 163.367
R1400 B.n211 B.n200 163.367
R1401 B.n211 B.n210 163.367
R1402 B.n210 B.n209 163.367
R1403 B.n209 B.n202 163.367
R1404 B.n205 B.n202 163.367
R1405 B.n205 B.n204 163.367
R1406 B.n204 B.n2 163.367
R1407 B.n782 B.n2 163.367
R1408 B.n782 B.n781 163.367
R1409 B.n781 B.n780 163.367
R1410 B.n780 B.n3 163.367
R1411 B.n776 B.n3 163.367
R1412 B.n776 B.n775 163.367
R1413 B.n775 B.n774 163.367
R1414 B.n774 B.n5 163.367
R1415 B.n770 B.n5 163.367
R1416 B.n770 B.n769 163.367
R1417 B.n769 B.n768 163.367
R1418 B.n768 B.n7 163.367
R1419 B.n764 B.n7 163.367
R1420 B.n764 B.n763 163.367
R1421 B.n763 B.n762 163.367
R1422 B.n762 B.n9 163.367
R1423 B.n758 B.n9 163.367
R1424 B.n758 B.n757 163.367
R1425 B.n757 B.n756 163.367
R1426 B.n756 B.n11 163.367
R1427 B.n752 B.n11 163.367
R1428 B.n752 B.n751 163.367
R1429 B.n751 B.n750 163.367
R1430 B.n750 B.n13 163.367
R1431 B.n746 B.n13 163.367
R1432 B.n746 B.n745 163.367
R1433 B.n745 B.n744 163.367
R1434 B.n744 B.n15 163.367
R1435 B.n740 B.n15 163.367
R1436 B.n740 B.n739 163.367
R1437 B.n739 B.n738 163.367
R1438 B.n738 B.n17 163.367
R1439 B.n734 B.n17 163.367
R1440 B.n734 B.n733 163.367
R1441 B.n733 B.n732 163.367
R1442 B.n732 B.n19 163.367
R1443 B.n257 B.n186 163.367
R1444 B.n258 B.n257 163.367
R1445 B.n259 B.n258 163.367
R1446 B.n259 B.n184 163.367
R1447 B.n263 B.n184 163.367
R1448 B.n264 B.n263 163.367
R1449 B.n265 B.n264 163.367
R1450 B.n265 B.n182 163.367
R1451 B.n269 B.n182 163.367
R1452 B.n270 B.n269 163.367
R1453 B.n271 B.n270 163.367
R1454 B.n271 B.n180 163.367
R1455 B.n275 B.n180 163.367
R1456 B.n276 B.n275 163.367
R1457 B.n277 B.n276 163.367
R1458 B.n277 B.n178 163.367
R1459 B.n281 B.n178 163.367
R1460 B.n282 B.n281 163.367
R1461 B.n283 B.n282 163.367
R1462 B.n283 B.n176 163.367
R1463 B.n287 B.n176 163.367
R1464 B.n288 B.n287 163.367
R1465 B.n289 B.n288 163.367
R1466 B.n289 B.n174 163.367
R1467 B.n293 B.n174 163.367
R1468 B.n294 B.n293 163.367
R1469 B.n295 B.n294 163.367
R1470 B.n295 B.n172 163.367
R1471 B.n299 B.n172 163.367
R1472 B.n300 B.n299 163.367
R1473 B.n301 B.n300 163.367
R1474 B.n301 B.n170 163.367
R1475 B.n305 B.n170 163.367
R1476 B.n306 B.n305 163.367
R1477 B.n307 B.n306 163.367
R1478 B.n307 B.n168 163.367
R1479 B.n311 B.n168 163.367
R1480 B.n312 B.n311 163.367
R1481 B.n313 B.n312 163.367
R1482 B.n313 B.n166 163.367
R1483 B.n317 B.n166 163.367
R1484 B.n318 B.n317 163.367
R1485 B.n319 B.n318 163.367
R1486 B.n319 B.n164 163.367
R1487 B.n323 B.n164 163.367
R1488 B.n324 B.n323 163.367
R1489 B.n325 B.n324 163.367
R1490 B.n325 B.n162 163.367
R1491 B.n329 B.n162 163.367
R1492 B.n330 B.n329 163.367
R1493 B.n331 B.n330 163.367
R1494 B.n331 B.n160 163.367
R1495 B.n335 B.n160 163.367
R1496 B.n336 B.n335 163.367
R1497 B.n337 B.n336 163.367
R1498 B.n337 B.n156 163.367
R1499 B.n342 B.n156 163.367
R1500 B.n343 B.n342 163.367
R1501 B.n344 B.n343 163.367
R1502 B.n344 B.n154 163.367
R1503 B.n348 B.n154 163.367
R1504 B.n349 B.n348 163.367
R1505 B.n350 B.n349 163.367
R1506 B.n350 B.n152 163.367
R1507 B.n354 B.n152 163.367
R1508 B.n355 B.n354 163.367
R1509 B.n355 B.n148 163.367
R1510 B.n359 B.n148 163.367
R1511 B.n360 B.n359 163.367
R1512 B.n361 B.n360 163.367
R1513 B.n361 B.n146 163.367
R1514 B.n365 B.n146 163.367
R1515 B.n366 B.n365 163.367
R1516 B.n367 B.n366 163.367
R1517 B.n367 B.n144 163.367
R1518 B.n371 B.n144 163.367
R1519 B.n372 B.n371 163.367
R1520 B.n373 B.n372 163.367
R1521 B.n373 B.n142 163.367
R1522 B.n377 B.n142 163.367
R1523 B.n378 B.n377 163.367
R1524 B.n379 B.n378 163.367
R1525 B.n379 B.n140 163.367
R1526 B.n383 B.n140 163.367
R1527 B.n384 B.n383 163.367
R1528 B.n385 B.n384 163.367
R1529 B.n385 B.n138 163.367
R1530 B.n389 B.n138 163.367
R1531 B.n390 B.n389 163.367
R1532 B.n391 B.n390 163.367
R1533 B.n391 B.n136 163.367
R1534 B.n395 B.n136 163.367
R1535 B.n396 B.n395 163.367
R1536 B.n397 B.n396 163.367
R1537 B.n397 B.n134 163.367
R1538 B.n401 B.n134 163.367
R1539 B.n402 B.n401 163.367
R1540 B.n403 B.n402 163.367
R1541 B.n403 B.n132 163.367
R1542 B.n407 B.n132 163.367
R1543 B.n408 B.n407 163.367
R1544 B.n409 B.n408 163.367
R1545 B.n409 B.n130 163.367
R1546 B.n413 B.n130 163.367
R1547 B.n414 B.n413 163.367
R1548 B.n415 B.n414 163.367
R1549 B.n415 B.n128 163.367
R1550 B.n419 B.n128 163.367
R1551 B.n420 B.n419 163.367
R1552 B.n421 B.n420 163.367
R1553 B.n421 B.n126 163.367
R1554 B.n425 B.n126 163.367
R1555 B.n426 B.n425 163.367
R1556 B.n427 B.n426 163.367
R1557 B.n427 B.n124 163.367
R1558 B.n431 B.n124 163.367
R1559 B.n432 B.n431 163.367
R1560 B.n433 B.n432 163.367
R1561 B.n433 B.n122 163.367
R1562 B.n437 B.n122 163.367
R1563 B.n438 B.n437 163.367
R1564 B.n439 B.n120 163.367
R1565 B.n443 B.n120 163.367
R1566 B.n444 B.n443 163.367
R1567 B.n445 B.n444 163.367
R1568 B.n445 B.n118 163.367
R1569 B.n449 B.n118 163.367
R1570 B.n450 B.n449 163.367
R1571 B.n451 B.n450 163.367
R1572 B.n451 B.n116 163.367
R1573 B.n455 B.n116 163.367
R1574 B.n456 B.n455 163.367
R1575 B.n457 B.n456 163.367
R1576 B.n457 B.n114 163.367
R1577 B.n461 B.n114 163.367
R1578 B.n462 B.n461 163.367
R1579 B.n463 B.n462 163.367
R1580 B.n463 B.n112 163.367
R1581 B.n467 B.n112 163.367
R1582 B.n468 B.n467 163.367
R1583 B.n469 B.n468 163.367
R1584 B.n469 B.n110 163.367
R1585 B.n473 B.n110 163.367
R1586 B.n474 B.n473 163.367
R1587 B.n475 B.n474 163.367
R1588 B.n475 B.n108 163.367
R1589 B.n479 B.n108 163.367
R1590 B.n480 B.n479 163.367
R1591 B.n481 B.n480 163.367
R1592 B.n481 B.n106 163.367
R1593 B.n485 B.n106 163.367
R1594 B.n486 B.n485 163.367
R1595 B.n487 B.n486 163.367
R1596 B.n487 B.n104 163.367
R1597 B.n491 B.n104 163.367
R1598 B.n492 B.n491 163.367
R1599 B.n493 B.n492 163.367
R1600 B.n493 B.n102 163.367
R1601 B.n497 B.n102 163.367
R1602 B.n498 B.n497 163.367
R1603 B.n499 B.n498 163.367
R1604 B.n499 B.n100 163.367
R1605 B.n503 B.n100 163.367
R1606 B.n504 B.n503 163.367
R1607 B.n505 B.n504 163.367
R1608 B.n505 B.n98 163.367
R1609 B.n509 B.n98 163.367
R1610 B.n510 B.n509 163.367
R1611 B.n511 B.n510 163.367
R1612 B.n511 B.n96 163.367
R1613 B.n515 B.n96 163.367
R1614 B.n516 B.n515 163.367
R1615 B.n517 B.n516 163.367
R1616 B.n517 B.n94 163.367
R1617 B.n521 B.n94 163.367
R1618 B.n522 B.n521 163.367
R1619 B.n523 B.n522 163.367
R1620 B.n523 B.n92 163.367
R1621 B.n527 B.n92 163.367
R1622 B.n528 B.n527 163.367
R1623 B.n529 B.n528 163.367
R1624 B.n529 B.n90 163.367
R1625 B.n533 B.n90 163.367
R1626 B.n534 B.n533 163.367
R1627 B.n535 B.n534 163.367
R1628 B.n535 B.n88 163.367
R1629 B.n539 B.n88 163.367
R1630 B.n540 B.n539 163.367
R1631 B.n541 B.n540 163.367
R1632 B.n541 B.n86 163.367
R1633 B.n545 B.n86 163.367
R1634 B.n728 B.n727 163.367
R1635 B.n727 B.n726 163.367
R1636 B.n726 B.n21 163.367
R1637 B.n722 B.n21 163.367
R1638 B.n722 B.n721 163.367
R1639 B.n721 B.n720 163.367
R1640 B.n720 B.n23 163.367
R1641 B.n716 B.n23 163.367
R1642 B.n716 B.n715 163.367
R1643 B.n715 B.n714 163.367
R1644 B.n714 B.n25 163.367
R1645 B.n710 B.n25 163.367
R1646 B.n710 B.n709 163.367
R1647 B.n709 B.n708 163.367
R1648 B.n708 B.n27 163.367
R1649 B.n704 B.n27 163.367
R1650 B.n704 B.n703 163.367
R1651 B.n703 B.n702 163.367
R1652 B.n702 B.n29 163.367
R1653 B.n698 B.n29 163.367
R1654 B.n698 B.n697 163.367
R1655 B.n697 B.n696 163.367
R1656 B.n696 B.n31 163.367
R1657 B.n692 B.n31 163.367
R1658 B.n692 B.n691 163.367
R1659 B.n691 B.n690 163.367
R1660 B.n690 B.n33 163.367
R1661 B.n686 B.n33 163.367
R1662 B.n686 B.n685 163.367
R1663 B.n685 B.n684 163.367
R1664 B.n684 B.n35 163.367
R1665 B.n680 B.n35 163.367
R1666 B.n680 B.n679 163.367
R1667 B.n679 B.n678 163.367
R1668 B.n678 B.n37 163.367
R1669 B.n674 B.n37 163.367
R1670 B.n674 B.n673 163.367
R1671 B.n673 B.n672 163.367
R1672 B.n672 B.n39 163.367
R1673 B.n668 B.n39 163.367
R1674 B.n668 B.n667 163.367
R1675 B.n667 B.n666 163.367
R1676 B.n666 B.n41 163.367
R1677 B.n662 B.n41 163.367
R1678 B.n662 B.n661 163.367
R1679 B.n661 B.n660 163.367
R1680 B.n660 B.n43 163.367
R1681 B.n656 B.n43 163.367
R1682 B.n656 B.n655 163.367
R1683 B.n655 B.n654 163.367
R1684 B.n654 B.n45 163.367
R1685 B.n650 B.n45 163.367
R1686 B.n650 B.n649 163.367
R1687 B.n649 B.n648 163.367
R1688 B.n648 B.n47 163.367
R1689 B.n643 B.n47 163.367
R1690 B.n643 B.n642 163.367
R1691 B.n642 B.n641 163.367
R1692 B.n641 B.n51 163.367
R1693 B.n637 B.n51 163.367
R1694 B.n637 B.n636 163.367
R1695 B.n636 B.n635 163.367
R1696 B.n635 B.n53 163.367
R1697 B.n631 B.n53 163.367
R1698 B.n631 B.n630 163.367
R1699 B.n630 B.n629 163.367
R1700 B.n629 B.n55 163.367
R1701 B.n625 B.n55 163.367
R1702 B.n625 B.n624 163.367
R1703 B.n624 B.n623 163.367
R1704 B.n623 B.n60 163.367
R1705 B.n619 B.n60 163.367
R1706 B.n619 B.n618 163.367
R1707 B.n618 B.n617 163.367
R1708 B.n617 B.n62 163.367
R1709 B.n613 B.n62 163.367
R1710 B.n613 B.n612 163.367
R1711 B.n612 B.n611 163.367
R1712 B.n611 B.n64 163.367
R1713 B.n607 B.n64 163.367
R1714 B.n607 B.n606 163.367
R1715 B.n606 B.n605 163.367
R1716 B.n605 B.n66 163.367
R1717 B.n601 B.n66 163.367
R1718 B.n601 B.n600 163.367
R1719 B.n600 B.n599 163.367
R1720 B.n599 B.n68 163.367
R1721 B.n595 B.n68 163.367
R1722 B.n595 B.n594 163.367
R1723 B.n594 B.n593 163.367
R1724 B.n593 B.n70 163.367
R1725 B.n589 B.n70 163.367
R1726 B.n589 B.n588 163.367
R1727 B.n588 B.n587 163.367
R1728 B.n587 B.n72 163.367
R1729 B.n583 B.n72 163.367
R1730 B.n583 B.n582 163.367
R1731 B.n582 B.n581 163.367
R1732 B.n581 B.n74 163.367
R1733 B.n577 B.n74 163.367
R1734 B.n577 B.n576 163.367
R1735 B.n576 B.n575 163.367
R1736 B.n575 B.n76 163.367
R1737 B.n571 B.n76 163.367
R1738 B.n571 B.n570 163.367
R1739 B.n570 B.n569 163.367
R1740 B.n569 B.n78 163.367
R1741 B.n565 B.n78 163.367
R1742 B.n565 B.n564 163.367
R1743 B.n564 B.n563 163.367
R1744 B.n563 B.n80 163.367
R1745 B.n559 B.n80 163.367
R1746 B.n559 B.n558 163.367
R1747 B.n558 B.n557 163.367
R1748 B.n557 B.n82 163.367
R1749 B.n553 B.n82 163.367
R1750 B.n553 B.n552 163.367
R1751 B.n552 B.n551 163.367
R1752 B.n551 B.n84 163.367
R1753 B.n547 B.n84 163.367
R1754 B.n547 B.n546 163.367
R1755 B.n151 B.n150 59.5399
R1756 B.n339 B.n158 59.5399
R1757 B.n645 B.n49 59.5399
R1758 B.n58 B.n57 59.5399
R1759 B.n730 B.n729 31.0639
R1760 B.n544 B.n85 31.0639
R1761 B.n440 B.n121 31.0639
R1762 B.n255 B.n254 31.0639
R1763 B.n150 B.n149 29.4793
R1764 B.n158 B.n157 29.4793
R1765 B.n49 B.n48 29.4793
R1766 B.n57 B.n56 29.4793
R1767 B B.n783 18.0485
R1768 B.n729 B.n20 10.6151
R1769 B.n725 B.n20 10.6151
R1770 B.n725 B.n724 10.6151
R1771 B.n724 B.n723 10.6151
R1772 B.n723 B.n22 10.6151
R1773 B.n719 B.n22 10.6151
R1774 B.n719 B.n718 10.6151
R1775 B.n718 B.n717 10.6151
R1776 B.n717 B.n24 10.6151
R1777 B.n713 B.n24 10.6151
R1778 B.n713 B.n712 10.6151
R1779 B.n712 B.n711 10.6151
R1780 B.n711 B.n26 10.6151
R1781 B.n707 B.n26 10.6151
R1782 B.n707 B.n706 10.6151
R1783 B.n706 B.n705 10.6151
R1784 B.n705 B.n28 10.6151
R1785 B.n701 B.n28 10.6151
R1786 B.n701 B.n700 10.6151
R1787 B.n700 B.n699 10.6151
R1788 B.n699 B.n30 10.6151
R1789 B.n695 B.n30 10.6151
R1790 B.n695 B.n694 10.6151
R1791 B.n694 B.n693 10.6151
R1792 B.n693 B.n32 10.6151
R1793 B.n689 B.n32 10.6151
R1794 B.n689 B.n688 10.6151
R1795 B.n688 B.n687 10.6151
R1796 B.n687 B.n34 10.6151
R1797 B.n683 B.n34 10.6151
R1798 B.n683 B.n682 10.6151
R1799 B.n682 B.n681 10.6151
R1800 B.n681 B.n36 10.6151
R1801 B.n677 B.n36 10.6151
R1802 B.n677 B.n676 10.6151
R1803 B.n676 B.n675 10.6151
R1804 B.n675 B.n38 10.6151
R1805 B.n671 B.n38 10.6151
R1806 B.n671 B.n670 10.6151
R1807 B.n670 B.n669 10.6151
R1808 B.n669 B.n40 10.6151
R1809 B.n665 B.n40 10.6151
R1810 B.n665 B.n664 10.6151
R1811 B.n664 B.n663 10.6151
R1812 B.n663 B.n42 10.6151
R1813 B.n659 B.n42 10.6151
R1814 B.n659 B.n658 10.6151
R1815 B.n658 B.n657 10.6151
R1816 B.n657 B.n44 10.6151
R1817 B.n653 B.n44 10.6151
R1818 B.n653 B.n652 10.6151
R1819 B.n652 B.n651 10.6151
R1820 B.n651 B.n46 10.6151
R1821 B.n647 B.n46 10.6151
R1822 B.n647 B.n646 10.6151
R1823 B.n644 B.n50 10.6151
R1824 B.n640 B.n50 10.6151
R1825 B.n640 B.n639 10.6151
R1826 B.n639 B.n638 10.6151
R1827 B.n638 B.n52 10.6151
R1828 B.n634 B.n52 10.6151
R1829 B.n634 B.n633 10.6151
R1830 B.n633 B.n632 10.6151
R1831 B.n632 B.n54 10.6151
R1832 B.n628 B.n627 10.6151
R1833 B.n627 B.n626 10.6151
R1834 B.n626 B.n59 10.6151
R1835 B.n622 B.n59 10.6151
R1836 B.n622 B.n621 10.6151
R1837 B.n621 B.n620 10.6151
R1838 B.n620 B.n61 10.6151
R1839 B.n616 B.n61 10.6151
R1840 B.n616 B.n615 10.6151
R1841 B.n615 B.n614 10.6151
R1842 B.n614 B.n63 10.6151
R1843 B.n610 B.n63 10.6151
R1844 B.n610 B.n609 10.6151
R1845 B.n609 B.n608 10.6151
R1846 B.n608 B.n65 10.6151
R1847 B.n604 B.n65 10.6151
R1848 B.n604 B.n603 10.6151
R1849 B.n603 B.n602 10.6151
R1850 B.n602 B.n67 10.6151
R1851 B.n598 B.n67 10.6151
R1852 B.n598 B.n597 10.6151
R1853 B.n597 B.n596 10.6151
R1854 B.n596 B.n69 10.6151
R1855 B.n592 B.n69 10.6151
R1856 B.n592 B.n591 10.6151
R1857 B.n591 B.n590 10.6151
R1858 B.n590 B.n71 10.6151
R1859 B.n586 B.n71 10.6151
R1860 B.n586 B.n585 10.6151
R1861 B.n585 B.n584 10.6151
R1862 B.n584 B.n73 10.6151
R1863 B.n580 B.n73 10.6151
R1864 B.n580 B.n579 10.6151
R1865 B.n579 B.n578 10.6151
R1866 B.n578 B.n75 10.6151
R1867 B.n574 B.n75 10.6151
R1868 B.n574 B.n573 10.6151
R1869 B.n573 B.n572 10.6151
R1870 B.n572 B.n77 10.6151
R1871 B.n568 B.n77 10.6151
R1872 B.n568 B.n567 10.6151
R1873 B.n567 B.n566 10.6151
R1874 B.n566 B.n79 10.6151
R1875 B.n562 B.n79 10.6151
R1876 B.n562 B.n561 10.6151
R1877 B.n561 B.n560 10.6151
R1878 B.n560 B.n81 10.6151
R1879 B.n556 B.n81 10.6151
R1880 B.n556 B.n555 10.6151
R1881 B.n555 B.n554 10.6151
R1882 B.n554 B.n83 10.6151
R1883 B.n550 B.n83 10.6151
R1884 B.n550 B.n549 10.6151
R1885 B.n549 B.n548 10.6151
R1886 B.n548 B.n85 10.6151
R1887 B.n441 B.n440 10.6151
R1888 B.n442 B.n441 10.6151
R1889 B.n442 B.n119 10.6151
R1890 B.n446 B.n119 10.6151
R1891 B.n447 B.n446 10.6151
R1892 B.n448 B.n447 10.6151
R1893 B.n448 B.n117 10.6151
R1894 B.n452 B.n117 10.6151
R1895 B.n453 B.n452 10.6151
R1896 B.n454 B.n453 10.6151
R1897 B.n454 B.n115 10.6151
R1898 B.n458 B.n115 10.6151
R1899 B.n459 B.n458 10.6151
R1900 B.n460 B.n459 10.6151
R1901 B.n460 B.n113 10.6151
R1902 B.n464 B.n113 10.6151
R1903 B.n465 B.n464 10.6151
R1904 B.n466 B.n465 10.6151
R1905 B.n466 B.n111 10.6151
R1906 B.n470 B.n111 10.6151
R1907 B.n471 B.n470 10.6151
R1908 B.n472 B.n471 10.6151
R1909 B.n472 B.n109 10.6151
R1910 B.n476 B.n109 10.6151
R1911 B.n477 B.n476 10.6151
R1912 B.n478 B.n477 10.6151
R1913 B.n478 B.n107 10.6151
R1914 B.n482 B.n107 10.6151
R1915 B.n483 B.n482 10.6151
R1916 B.n484 B.n483 10.6151
R1917 B.n484 B.n105 10.6151
R1918 B.n488 B.n105 10.6151
R1919 B.n489 B.n488 10.6151
R1920 B.n490 B.n489 10.6151
R1921 B.n490 B.n103 10.6151
R1922 B.n494 B.n103 10.6151
R1923 B.n495 B.n494 10.6151
R1924 B.n496 B.n495 10.6151
R1925 B.n496 B.n101 10.6151
R1926 B.n500 B.n101 10.6151
R1927 B.n501 B.n500 10.6151
R1928 B.n502 B.n501 10.6151
R1929 B.n502 B.n99 10.6151
R1930 B.n506 B.n99 10.6151
R1931 B.n507 B.n506 10.6151
R1932 B.n508 B.n507 10.6151
R1933 B.n508 B.n97 10.6151
R1934 B.n512 B.n97 10.6151
R1935 B.n513 B.n512 10.6151
R1936 B.n514 B.n513 10.6151
R1937 B.n514 B.n95 10.6151
R1938 B.n518 B.n95 10.6151
R1939 B.n519 B.n518 10.6151
R1940 B.n520 B.n519 10.6151
R1941 B.n520 B.n93 10.6151
R1942 B.n524 B.n93 10.6151
R1943 B.n525 B.n524 10.6151
R1944 B.n526 B.n525 10.6151
R1945 B.n526 B.n91 10.6151
R1946 B.n530 B.n91 10.6151
R1947 B.n531 B.n530 10.6151
R1948 B.n532 B.n531 10.6151
R1949 B.n532 B.n89 10.6151
R1950 B.n536 B.n89 10.6151
R1951 B.n537 B.n536 10.6151
R1952 B.n538 B.n537 10.6151
R1953 B.n538 B.n87 10.6151
R1954 B.n542 B.n87 10.6151
R1955 B.n543 B.n542 10.6151
R1956 B.n544 B.n543 10.6151
R1957 B.n256 B.n255 10.6151
R1958 B.n256 B.n185 10.6151
R1959 B.n260 B.n185 10.6151
R1960 B.n261 B.n260 10.6151
R1961 B.n262 B.n261 10.6151
R1962 B.n262 B.n183 10.6151
R1963 B.n266 B.n183 10.6151
R1964 B.n267 B.n266 10.6151
R1965 B.n268 B.n267 10.6151
R1966 B.n268 B.n181 10.6151
R1967 B.n272 B.n181 10.6151
R1968 B.n273 B.n272 10.6151
R1969 B.n274 B.n273 10.6151
R1970 B.n274 B.n179 10.6151
R1971 B.n278 B.n179 10.6151
R1972 B.n279 B.n278 10.6151
R1973 B.n280 B.n279 10.6151
R1974 B.n280 B.n177 10.6151
R1975 B.n284 B.n177 10.6151
R1976 B.n285 B.n284 10.6151
R1977 B.n286 B.n285 10.6151
R1978 B.n286 B.n175 10.6151
R1979 B.n290 B.n175 10.6151
R1980 B.n291 B.n290 10.6151
R1981 B.n292 B.n291 10.6151
R1982 B.n292 B.n173 10.6151
R1983 B.n296 B.n173 10.6151
R1984 B.n297 B.n296 10.6151
R1985 B.n298 B.n297 10.6151
R1986 B.n298 B.n171 10.6151
R1987 B.n302 B.n171 10.6151
R1988 B.n303 B.n302 10.6151
R1989 B.n304 B.n303 10.6151
R1990 B.n304 B.n169 10.6151
R1991 B.n308 B.n169 10.6151
R1992 B.n309 B.n308 10.6151
R1993 B.n310 B.n309 10.6151
R1994 B.n310 B.n167 10.6151
R1995 B.n314 B.n167 10.6151
R1996 B.n315 B.n314 10.6151
R1997 B.n316 B.n315 10.6151
R1998 B.n316 B.n165 10.6151
R1999 B.n320 B.n165 10.6151
R2000 B.n321 B.n320 10.6151
R2001 B.n322 B.n321 10.6151
R2002 B.n322 B.n163 10.6151
R2003 B.n326 B.n163 10.6151
R2004 B.n327 B.n326 10.6151
R2005 B.n328 B.n327 10.6151
R2006 B.n328 B.n161 10.6151
R2007 B.n332 B.n161 10.6151
R2008 B.n333 B.n332 10.6151
R2009 B.n334 B.n333 10.6151
R2010 B.n334 B.n159 10.6151
R2011 B.n338 B.n159 10.6151
R2012 B.n341 B.n340 10.6151
R2013 B.n341 B.n155 10.6151
R2014 B.n345 B.n155 10.6151
R2015 B.n346 B.n345 10.6151
R2016 B.n347 B.n346 10.6151
R2017 B.n347 B.n153 10.6151
R2018 B.n351 B.n153 10.6151
R2019 B.n352 B.n351 10.6151
R2020 B.n353 B.n352 10.6151
R2021 B.n357 B.n356 10.6151
R2022 B.n358 B.n357 10.6151
R2023 B.n358 B.n147 10.6151
R2024 B.n362 B.n147 10.6151
R2025 B.n363 B.n362 10.6151
R2026 B.n364 B.n363 10.6151
R2027 B.n364 B.n145 10.6151
R2028 B.n368 B.n145 10.6151
R2029 B.n369 B.n368 10.6151
R2030 B.n370 B.n369 10.6151
R2031 B.n370 B.n143 10.6151
R2032 B.n374 B.n143 10.6151
R2033 B.n375 B.n374 10.6151
R2034 B.n376 B.n375 10.6151
R2035 B.n376 B.n141 10.6151
R2036 B.n380 B.n141 10.6151
R2037 B.n381 B.n380 10.6151
R2038 B.n382 B.n381 10.6151
R2039 B.n382 B.n139 10.6151
R2040 B.n386 B.n139 10.6151
R2041 B.n387 B.n386 10.6151
R2042 B.n388 B.n387 10.6151
R2043 B.n388 B.n137 10.6151
R2044 B.n392 B.n137 10.6151
R2045 B.n393 B.n392 10.6151
R2046 B.n394 B.n393 10.6151
R2047 B.n394 B.n135 10.6151
R2048 B.n398 B.n135 10.6151
R2049 B.n399 B.n398 10.6151
R2050 B.n400 B.n399 10.6151
R2051 B.n400 B.n133 10.6151
R2052 B.n404 B.n133 10.6151
R2053 B.n405 B.n404 10.6151
R2054 B.n406 B.n405 10.6151
R2055 B.n406 B.n131 10.6151
R2056 B.n410 B.n131 10.6151
R2057 B.n411 B.n410 10.6151
R2058 B.n412 B.n411 10.6151
R2059 B.n412 B.n129 10.6151
R2060 B.n416 B.n129 10.6151
R2061 B.n417 B.n416 10.6151
R2062 B.n418 B.n417 10.6151
R2063 B.n418 B.n127 10.6151
R2064 B.n422 B.n127 10.6151
R2065 B.n423 B.n422 10.6151
R2066 B.n424 B.n423 10.6151
R2067 B.n424 B.n125 10.6151
R2068 B.n428 B.n125 10.6151
R2069 B.n429 B.n428 10.6151
R2070 B.n430 B.n429 10.6151
R2071 B.n430 B.n123 10.6151
R2072 B.n434 B.n123 10.6151
R2073 B.n435 B.n434 10.6151
R2074 B.n436 B.n435 10.6151
R2075 B.n436 B.n121 10.6151
R2076 B.n254 B.n187 10.6151
R2077 B.n250 B.n187 10.6151
R2078 B.n250 B.n249 10.6151
R2079 B.n249 B.n248 10.6151
R2080 B.n248 B.n189 10.6151
R2081 B.n244 B.n189 10.6151
R2082 B.n244 B.n243 10.6151
R2083 B.n243 B.n242 10.6151
R2084 B.n242 B.n191 10.6151
R2085 B.n238 B.n191 10.6151
R2086 B.n238 B.n237 10.6151
R2087 B.n237 B.n236 10.6151
R2088 B.n236 B.n193 10.6151
R2089 B.n232 B.n193 10.6151
R2090 B.n232 B.n231 10.6151
R2091 B.n231 B.n230 10.6151
R2092 B.n230 B.n195 10.6151
R2093 B.n226 B.n195 10.6151
R2094 B.n226 B.n225 10.6151
R2095 B.n225 B.n224 10.6151
R2096 B.n224 B.n197 10.6151
R2097 B.n220 B.n197 10.6151
R2098 B.n220 B.n219 10.6151
R2099 B.n219 B.n218 10.6151
R2100 B.n218 B.n199 10.6151
R2101 B.n214 B.n199 10.6151
R2102 B.n214 B.n213 10.6151
R2103 B.n213 B.n212 10.6151
R2104 B.n212 B.n201 10.6151
R2105 B.n208 B.n201 10.6151
R2106 B.n208 B.n207 10.6151
R2107 B.n207 B.n206 10.6151
R2108 B.n206 B.n203 10.6151
R2109 B.n203 B.n0 10.6151
R2110 B.n779 B.n1 10.6151
R2111 B.n779 B.n778 10.6151
R2112 B.n778 B.n777 10.6151
R2113 B.n777 B.n4 10.6151
R2114 B.n773 B.n4 10.6151
R2115 B.n773 B.n772 10.6151
R2116 B.n772 B.n771 10.6151
R2117 B.n771 B.n6 10.6151
R2118 B.n767 B.n6 10.6151
R2119 B.n767 B.n766 10.6151
R2120 B.n766 B.n765 10.6151
R2121 B.n765 B.n8 10.6151
R2122 B.n761 B.n8 10.6151
R2123 B.n761 B.n760 10.6151
R2124 B.n760 B.n759 10.6151
R2125 B.n759 B.n10 10.6151
R2126 B.n755 B.n10 10.6151
R2127 B.n755 B.n754 10.6151
R2128 B.n754 B.n753 10.6151
R2129 B.n753 B.n12 10.6151
R2130 B.n749 B.n12 10.6151
R2131 B.n749 B.n748 10.6151
R2132 B.n748 B.n747 10.6151
R2133 B.n747 B.n14 10.6151
R2134 B.n743 B.n14 10.6151
R2135 B.n743 B.n742 10.6151
R2136 B.n742 B.n741 10.6151
R2137 B.n741 B.n16 10.6151
R2138 B.n737 B.n16 10.6151
R2139 B.n737 B.n736 10.6151
R2140 B.n736 B.n735 10.6151
R2141 B.n735 B.n18 10.6151
R2142 B.n731 B.n18 10.6151
R2143 B.n731 B.n730 10.6151
R2144 B.n646 B.n645 9.36635
R2145 B.n628 B.n58 9.36635
R2146 B.n339 B.n338 9.36635
R2147 B.n356 B.n151 9.36635
R2148 B.n783 B.n0 2.81026
R2149 B.n783 B.n1 2.81026
R2150 B.n645 B.n644 1.24928
R2151 B.n58 B.n54 1.24928
R2152 B.n340 B.n339 1.24928
R2153 B.n353 B.n151 1.24928
R2154 VP.n13 VP.t3 394.978
R2155 VP.n30 VP.t8 376.488
R2156 VP.n47 VP.t2 376.488
R2157 VP.n27 VP.t5 376.488
R2158 VP.n5 VP.t4 343.072
R2159 VP.n3 VP.t0 343.072
R2160 VP.n1 VP.t7 343.072
R2161 VP.n8 VP.t6 343.072
R2162 VP.n10 VP.t9 343.072
R2163 VP.n12 VP.t1 343.072
R2164 VP.n15 VP.n14 161.3
R2165 VP.n16 VP.n11 161.3
R2166 VP.n18 VP.n17 161.3
R2167 VP.n20 VP.n19 161.3
R2168 VP.n21 VP.n9 161.3
R2169 VP.n23 VP.n22 161.3
R2170 VP.n25 VP.n24 161.3
R2171 VP.n26 VP.n7 161.3
R2172 VP.n46 VP.n0 161.3
R2173 VP.n45 VP.n44 161.3
R2174 VP.n43 VP.n42 161.3
R2175 VP.n41 VP.n2 161.3
R2176 VP.n40 VP.n39 161.3
R2177 VP.n38 VP.n37 161.3
R2178 VP.n36 VP.n4 161.3
R2179 VP.n35 VP.n34 161.3
R2180 VP.n33 VP.n32 161.3
R2181 VP.n31 VP.n6 161.3
R2182 VP.n28 VP.n27 80.6037
R2183 VP.n48 VP.n47 80.6037
R2184 VP.n30 VP.n29 80.6037
R2185 VP.n29 VP.n28 49.2968
R2186 VP.n13 VP.n12 44.4551
R2187 VP.n36 VP.n35 41.3843
R2188 VP.n42 VP.n41 41.3843
R2189 VP.n22 VP.n21 41.3843
R2190 VP.n16 VP.n15 41.3843
R2191 VP.n37 VP.n36 39.4369
R2192 VP.n41 VP.n40 39.4369
R2193 VP.n21 VP.n20 39.4369
R2194 VP.n17 VP.n16 39.4369
R2195 VP.n32 VP.n31 37.4894
R2196 VP.n46 VP.n45 37.4894
R2197 VP.n26 VP.n25 37.4894
R2198 VP.n14 VP.n13 29.7405
R2199 VP.n31 VP.n30 28.4823
R2200 VP.n47 VP.n46 28.4823
R2201 VP.n27 VP.n26 28.4823
R2202 VP.n35 VP.n5 13.146
R2203 VP.n42 VP.n1 13.146
R2204 VP.n22 VP.n8 13.146
R2205 VP.n15 VP.n12 13.146
R2206 VP.n37 VP.n3 12.1722
R2207 VP.n40 VP.n3 12.1722
R2208 VP.n17 VP.n10 12.1722
R2209 VP.n20 VP.n10 12.1722
R2210 VP.n32 VP.n5 11.1985
R2211 VP.n45 VP.n1 11.1985
R2212 VP.n25 VP.n8 11.1985
R2213 VP.n28 VP.n7 0.285035
R2214 VP.n29 VP.n6 0.285035
R2215 VP.n48 VP.n0 0.285035
R2216 VP.n14 VP.n11 0.189894
R2217 VP.n18 VP.n11 0.189894
R2218 VP.n19 VP.n18 0.189894
R2219 VP.n19 VP.n9 0.189894
R2220 VP.n23 VP.n9 0.189894
R2221 VP.n24 VP.n23 0.189894
R2222 VP.n24 VP.n7 0.189894
R2223 VP.n33 VP.n6 0.189894
R2224 VP.n34 VP.n33 0.189894
R2225 VP.n34 VP.n4 0.189894
R2226 VP.n38 VP.n4 0.189894
R2227 VP.n39 VP.n38 0.189894
R2228 VP.n39 VP.n2 0.189894
R2229 VP.n43 VP.n2 0.189894
R2230 VP.n44 VP.n43 0.189894
R2231 VP.n44 VP.n0 0.189894
R2232 VP VP.n48 0.146778
R2233 VDD1.n88 VDD1.n0 756.745
R2234 VDD1.n183 VDD1.n95 756.745
R2235 VDD1.n89 VDD1.n88 585
R2236 VDD1.n87 VDD1.n86 585
R2237 VDD1.n4 VDD1.n3 585
R2238 VDD1.n81 VDD1.n80 585
R2239 VDD1.n79 VDD1.n78 585
R2240 VDD1.n77 VDD1.n7 585
R2241 VDD1.n11 VDD1.n8 585
R2242 VDD1.n72 VDD1.n71 585
R2243 VDD1.n70 VDD1.n69 585
R2244 VDD1.n13 VDD1.n12 585
R2245 VDD1.n64 VDD1.n63 585
R2246 VDD1.n62 VDD1.n61 585
R2247 VDD1.n17 VDD1.n16 585
R2248 VDD1.n56 VDD1.n55 585
R2249 VDD1.n54 VDD1.n53 585
R2250 VDD1.n21 VDD1.n20 585
R2251 VDD1.n48 VDD1.n47 585
R2252 VDD1.n46 VDD1.n45 585
R2253 VDD1.n25 VDD1.n24 585
R2254 VDD1.n40 VDD1.n39 585
R2255 VDD1.n38 VDD1.n37 585
R2256 VDD1.n29 VDD1.n28 585
R2257 VDD1.n32 VDD1.n31 585
R2258 VDD1.n126 VDD1.n125 585
R2259 VDD1.n123 VDD1.n122 585
R2260 VDD1.n132 VDD1.n131 585
R2261 VDD1.n134 VDD1.n133 585
R2262 VDD1.n119 VDD1.n118 585
R2263 VDD1.n140 VDD1.n139 585
R2264 VDD1.n142 VDD1.n141 585
R2265 VDD1.n115 VDD1.n114 585
R2266 VDD1.n148 VDD1.n147 585
R2267 VDD1.n150 VDD1.n149 585
R2268 VDD1.n111 VDD1.n110 585
R2269 VDD1.n156 VDD1.n155 585
R2270 VDD1.n158 VDD1.n157 585
R2271 VDD1.n107 VDD1.n106 585
R2272 VDD1.n164 VDD1.n163 585
R2273 VDD1.n167 VDD1.n166 585
R2274 VDD1.n165 VDD1.n103 585
R2275 VDD1.n172 VDD1.n102 585
R2276 VDD1.n174 VDD1.n173 585
R2277 VDD1.n176 VDD1.n175 585
R2278 VDD1.n99 VDD1.n98 585
R2279 VDD1.n182 VDD1.n181 585
R2280 VDD1.n184 VDD1.n183 585
R2281 VDD1.t6 VDD1.n30 327.466
R2282 VDD1.t1 VDD1.n124 327.466
R2283 VDD1.n88 VDD1.n87 171.744
R2284 VDD1.n87 VDD1.n3 171.744
R2285 VDD1.n80 VDD1.n3 171.744
R2286 VDD1.n80 VDD1.n79 171.744
R2287 VDD1.n79 VDD1.n7 171.744
R2288 VDD1.n11 VDD1.n7 171.744
R2289 VDD1.n71 VDD1.n11 171.744
R2290 VDD1.n71 VDD1.n70 171.744
R2291 VDD1.n70 VDD1.n12 171.744
R2292 VDD1.n63 VDD1.n12 171.744
R2293 VDD1.n63 VDD1.n62 171.744
R2294 VDD1.n62 VDD1.n16 171.744
R2295 VDD1.n55 VDD1.n16 171.744
R2296 VDD1.n55 VDD1.n54 171.744
R2297 VDD1.n54 VDD1.n20 171.744
R2298 VDD1.n47 VDD1.n20 171.744
R2299 VDD1.n47 VDD1.n46 171.744
R2300 VDD1.n46 VDD1.n24 171.744
R2301 VDD1.n39 VDD1.n24 171.744
R2302 VDD1.n39 VDD1.n38 171.744
R2303 VDD1.n38 VDD1.n28 171.744
R2304 VDD1.n31 VDD1.n28 171.744
R2305 VDD1.n125 VDD1.n122 171.744
R2306 VDD1.n132 VDD1.n122 171.744
R2307 VDD1.n133 VDD1.n132 171.744
R2308 VDD1.n133 VDD1.n118 171.744
R2309 VDD1.n140 VDD1.n118 171.744
R2310 VDD1.n141 VDD1.n140 171.744
R2311 VDD1.n141 VDD1.n114 171.744
R2312 VDD1.n148 VDD1.n114 171.744
R2313 VDD1.n149 VDD1.n148 171.744
R2314 VDD1.n149 VDD1.n110 171.744
R2315 VDD1.n156 VDD1.n110 171.744
R2316 VDD1.n157 VDD1.n156 171.744
R2317 VDD1.n157 VDD1.n106 171.744
R2318 VDD1.n164 VDD1.n106 171.744
R2319 VDD1.n166 VDD1.n164 171.744
R2320 VDD1.n166 VDD1.n165 171.744
R2321 VDD1.n165 VDD1.n102 171.744
R2322 VDD1.n174 VDD1.n102 171.744
R2323 VDD1.n175 VDD1.n174 171.744
R2324 VDD1.n175 VDD1.n98 171.744
R2325 VDD1.n182 VDD1.n98 171.744
R2326 VDD1.n183 VDD1.n182 171.744
R2327 VDD1.n31 VDD1.t6 85.8723
R2328 VDD1.n125 VDD1.t1 85.8723
R2329 VDD1.n191 VDD1.n190 73.0344
R2330 VDD1.n94 VDD1.n93 72.1072
R2331 VDD1.n193 VDD1.n192 72.107
R2332 VDD1.n189 VDD1.n188 72.107
R2333 VDD1.n94 VDD1.n92 52.8896
R2334 VDD1.n189 VDD1.n187 52.8896
R2335 VDD1.n193 VDD1.n191 45.7811
R2336 VDD1.n32 VDD1.n30 16.3895
R2337 VDD1.n126 VDD1.n124 16.3895
R2338 VDD1.n78 VDD1.n77 13.1884
R2339 VDD1.n173 VDD1.n172 13.1884
R2340 VDD1.n81 VDD1.n6 12.8005
R2341 VDD1.n76 VDD1.n8 12.8005
R2342 VDD1.n33 VDD1.n29 12.8005
R2343 VDD1.n127 VDD1.n123 12.8005
R2344 VDD1.n171 VDD1.n103 12.8005
R2345 VDD1.n176 VDD1.n101 12.8005
R2346 VDD1.n82 VDD1.n4 12.0247
R2347 VDD1.n73 VDD1.n72 12.0247
R2348 VDD1.n37 VDD1.n36 12.0247
R2349 VDD1.n131 VDD1.n130 12.0247
R2350 VDD1.n168 VDD1.n167 12.0247
R2351 VDD1.n177 VDD1.n99 12.0247
R2352 VDD1.n86 VDD1.n85 11.249
R2353 VDD1.n69 VDD1.n10 11.249
R2354 VDD1.n40 VDD1.n27 11.249
R2355 VDD1.n134 VDD1.n121 11.249
R2356 VDD1.n163 VDD1.n105 11.249
R2357 VDD1.n181 VDD1.n180 11.249
R2358 VDD1.n89 VDD1.n2 10.4732
R2359 VDD1.n68 VDD1.n13 10.4732
R2360 VDD1.n41 VDD1.n25 10.4732
R2361 VDD1.n135 VDD1.n119 10.4732
R2362 VDD1.n162 VDD1.n107 10.4732
R2363 VDD1.n184 VDD1.n97 10.4732
R2364 VDD1.n90 VDD1.n0 9.69747
R2365 VDD1.n65 VDD1.n64 9.69747
R2366 VDD1.n45 VDD1.n44 9.69747
R2367 VDD1.n139 VDD1.n138 9.69747
R2368 VDD1.n159 VDD1.n158 9.69747
R2369 VDD1.n185 VDD1.n95 9.69747
R2370 VDD1.n92 VDD1.n91 9.45567
R2371 VDD1.n187 VDD1.n186 9.45567
R2372 VDD1.n58 VDD1.n57 9.3005
R2373 VDD1.n60 VDD1.n59 9.3005
R2374 VDD1.n15 VDD1.n14 9.3005
R2375 VDD1.n66 VDD1.n65 9.3005
R2376 VDD1.n68 VDD1.n67 9.3005
R2377 VDD1.n10 VDD1.n9 9.3005
R2378 VDD1.n74 VDD1.n73 9.3005
R2379 VDD1.n76 VDD1.n75 9.3005
R2380 VDD1.n91 VDD1.n90 9.3005
R2381 VDD1.n2 VDD1.n1 9.3005
R2382 VDD1.n85 VDD1.n84 9.3005
R2383 VDD1.n83 VDD1.n82 9.3005
R2384 VDD1.n6 VDD1.n5 9.3005
R2385 VDD1.n19 VDD1.n18 9.3005
R2386 VDD1.n52 VDD1.n51 9.3005
R2387 VDD1.n50 VDD1.n49 9.3005
R2388 VDD1.n23 VDD1.n22 9.3005
R2389 VDD1.n44 VDD1.n43 9.3005
R2390 VDD1.n42 VDD1.n41 9.3005
R2391 VDD1.n27 VDD1.n26 9.3005
R2392 VDD1.n36 VDD1.n35 9.3005
R2393 VDD1.n34 VDD1.n33 9.3005
R2394 VDD1.n186 VDD1.n185 9.3005
R2395 VDD1.n97 VDD1.n96 9.3005
R2396 VDD1.n180 VDD1.n179 9.3005
R2397 VDD1.n178 VDD1.n177 9.3005
R2398 VDD1.n101 VDD1.n100 9.3005
R2399 VDD1.n146 VDD1.n145 9.3005
R2400 VDD1.n144 VDD1.n143 9.3005
R2401 VDD1.n117 VDD1.n116 9.3005
R2402 VDD1.n138 VDD1.n137 9.3005
R2403 VDD1.n136 VDD1.n135 9.3005
R2404 VDD1.n121 VDD1.n120 9.3005
R2405 VDD1.n130 VDD1.n129 9.3005
R2406 VDD1.n128 VDD1.n127 9.3005
R2407 VDD1.n113 VDD1.n112 9.3005
R2408 VDD1.n152 VDD1.n151 9.3005
R2409 VDD1.n154 VDD1.n153 9.3005
R2410 VDD1.n109 VDD1.n108 9.3005
R2411 VDD1.n160 VDD1.n159 9.3005
R2412 VDD1.n162 VDD1.n161 9.3005
R2413 VDD1.n105 VDD1.n104 9.3005
R2414 VDD1.n169 VDD1.n168 9.3005
R2415 VDD1.n171 VDD1.n170 9.3005
R2416 VDD1.n61 VDD1.n15 8.92171
R2417 VDD1.n48 VDD1.n23 8.92171
R2418 VDD1.n142 VDD1.n117 8.92171
R2419 VDD1.n155 VDD1.n109 8.92171
R2420 VDD1.n60 VDD1.n17 8.14595
R2421 VDD1.n49 VDD1.n21 8.14595
R2422 VDD1.n143 VDD1.n115 8.14595
R2423 VDD1.n154 VDD1.n111 8.14595
R2424 VDD1.n57 VDD1.n56 7.3702
R2425 VDD1.n53 VDD1.n52 7.3702
R2426 VDD1.n147 VDD1.n146 7.3702
R2427 VDD1.n151 VDD1.n150 7.3702
R2428 VDD1.n56 VDD1.n19 6.59444
R2429 VDD1.n53 VDD1.n19 6.59444
R2430 VDD1.n147 VDD1.n113 6.59444
R2431 VDD1.n150 VDD1.n113 6.59444
R2432 VDD1.n57 VDD1.n17 5.81868
R2433 VDD1.n52 VDD1.n21 5.81868
R2434 VDD1.n146 VDD1.n115 5.81868
R2435 VDD1.n151 VDD1.n111 5.81868
R2436 VDD1.n61 VDD1.n60 5.04292
R2437 VDD1.n49 VDD1.n48 5.04292
R2438 VDD1.n143 VDD1.n142 5.04292
R2439 VDD1.n155 VDD1.n154 5.04292
R2440 VDD1.n92 VDD1.n0 4.26717
R2441 VDD1.n64 VDD1.n15 4.26717
R2442 VDD1.n45 VDD1.n23 4.26717
R2443 VDD1.n139 VDD1.n117 4.26717
R2444 VDD1.n158 VDD1.n109 4.26717
R2445 VDD1.n187 VDD1.n95 4.26717
R2446 VDD1.n34 VDD1.n30 3.70982
R2447 VDD1.n128 VDD1.n124 3.70982
R2448 VDD1.n90 VDD1.n89 3.49141
R2449 VDD1.n65 VDD1.n13 3.49141
R2450 VDD1.n44 VDD1.n25 3.49141
R2451 VDD1.n138 VDD1.n119 3.49141
R2452 VDD1.n159 VDD1.n107 3.49141
R2453 VDD1.n185 VDD1.n184 3.49141
R2454 VDD1.n86 VDD1.n2 2.71565
R2455 VDD1.n69 VDD1.n68 2.71565
R2456 VDD1.n41 VDD1.n40 2.71565
R2457 VDD1.n135 VDD1.n134 2.71565
R2458 VDD1.n163 VDD1.n162 2.71565
R2459 VDD1.n181 VDD1.n97 2.71565
R2460 VDD1.n85 VDD1.n4 1.93989
R2461 VDD1.n72 VDD1.n10 1.93989
R2462 VDD1.n37 VDD1.n27 1.93989
R2463 VDD1.n131 VDD1.n121 1.93989
R2464 VDD1.n167 VDD1.n105 1.93989
R2465 VDD1.n180 VDD1.n99 1.93989
R2466 VDD1.n192 VDD1.t3 1.91933
R2467 VDD1.n192 VDD1.t4 1.91933
R2468 VDD1.n93 VDD1.t8 1.91933
R2469 VDD1.n93 VDD1.t0 1.91933
R2470 VDD1.n190 VDD1.t2 1.91933
R2471 VDD1.n190 VDD1.t7 1.91933
R2472 VDD1.n188 VDD1.t5 1.91933
R2473 VDD1.n188 VDD1.t9 1.91933
R2474 VDD1.n82 VDD1.n81 1.16414
R2475 VDD1.n73 VDD1.n8 1.16414
R2476 VDD1.n36 VDD1.n29 1.16414
R2477 VDD1.n130 VDD1.n123 1.16414
R2478 VDD1.n168 VDD1.n103 1.16414
R2479 VDD1.n177 VDD1.n176 1.16414
R2480 VDD1 VDD1.n193 0.925069
R2481 VDD1.n78 VDD1.n6 0.388379
R2482 VDD1.n77 VDD1.n76 0.388379
R2483 VDD1.n33 VDD1.n32 0.388379
R2484 VDD1.n127 VDD1.n126 0.388379
R2485 VDD1.n172 VDD1.n171 0.388379
R2486 VDD1.n173 VDD1.n101 0.388379
R2487 VDD1 VDD1.n94 0.386276
R2488 VDD1.n191 VDD1.n189 0.27274
R2489 VDD1.n91 VDD1.n1 0.155672
R2490 VDD1.n84 VDD1.n1 0.155672
R2491 VDD1.n84 VDD1.n83 0.155672
R2492 VDD1.n83 VDD1.n5 0.155672
R2493 VDD1.n75 VDD1.n5 0.155672
R2494 VDD1.n75 VDD1.n74 0.155672
R2495 VDD1.n74 VDD1.n9 0.155672
R2496 VDD1.n67 VDD1.n9 0.155672
R2497 VDD1.n67 VDD1.n66 0.155672
R2498 VDD1.n66 VDD1.n14 0.155672
R2499 VDD1.n59 VDD1.n14 0.155672
R2500 VDD1.n59 VDD1.n58 0.155672
R2501 VDD1.n58 VDD1.n18 0.155672
R2502 VDD1.n51 VDD1.n18 0.155672
R2503 VDD1.n51 VDD1.n50 0.155672
R2504 VDD1.n50 VDD1.n22 0.155672
R2505 VDD1.n43 VDD1.n22 0.155672
R2506 VDD1.n43 VDD1.n42 0.155672
R2507 VDD1.n42 VDD1.n26 0.155672
R2508 VDD1.n35 VDD1.n26 0.155672
R2509 VDD1.n35 VDD1.n34 0.155672
R2510 VDD1.n129 VDD1.n128 0.155672
R2511 VDD1.n129 VDD1.n120 0.155672
R2512 VDD1.n136 VDD1.n120 0.155672
R2513 VDD1.n137 VDD1.n136 0.155672
R2514 VDD1.n137 VDD1.n116 0.155672
R2515 VDD1.n144 VDD1.n116 0.155672
R2516 VDD1.n145 VDD1.n144 0.155672
R2517 VDD1.n145 VDD1.n112 0.155672
R2518 VDD1.n152 VDD1.n112 0.155672
R2519 VDD1.n153 VDD1.n152 0.155672
R2520 VDD1.n153 VDD1.n108 0.155672
R2521 VDD1.n160 VDD1.n108 0.155672
R2522 VDD1.n161 VDD1.n160 0.155672
R2523 VDD1.n161 VDD1.n104 0.155672
R2524 VDD1.n169 VDD1.n104 0.155672
R2525 VDD1.n170 VDD1.n169 0.155672
R2526 VDD1.n170 VDD1.n100 0.155672
R2527 VDD1.n178 VDD1.n100 0.155672
R2528 VDD1.n179 VDD1.n178 0.155672
R2529 VDD1.n179 VDD1.n96 0.155672
R2530 VDD1.n186 VDD1.n96 0.155672
C0 VDD2 w_n2794_n4356# 2.66697f
C1 VP VTAIL 11.7306f
C2 B VN 0.979773f
C3 VP VN 7.24078f
C4 w_n2794_n4356# VTAIL 3.77399f
C5 B VP 1.57637f
C6 w_n2794_n4356# VN 5.65984f
C7 w_n2794_n4356# B 9.56036f
C8 VDD1 VDD2 1.27196f
C9 w_n2794_n4356# VP 6.01925f
C10 VDD1 VTAIL 15.119501f
C11 VDD2 VTAIL 15.156499f
C12 VDD1 VN 0.149408f
C13 VDD1 B 2.28379f
C14 VDD2 VN 11.8593f
C15 VDD2 B 2.34686f
C16 VDD1 VP 12.1081f
C17 VN VTAIL 11.716f
C18 VDD2 VP 0.403795f
C19 VDD1 w_n2794_n4356# 2.59673f
C20 B VTAIL 3.99873f
C21 VDD2 VSUBS 1.783807f
C22 VDD1 VSUBS 1.515424f
C23 VTAIL VSUBS 1.095286f
C24 VN VSUBS 5.83704f
C25 VP VSUBS 2.633802f
C26 B VSUBS 4.036532f
C27 w_n2794_n4356# VSUBS 0.148965p
C28 VDD1.n0 VSUBS 0.030247f
C29 VDD1.n1 VSUBS 0.027006f
C30 VDD1.n2 VSUBS 0.014512f
C31 VDD1.n3 VSUBS 0.0343f
C32 VDD1.n4 VSUBS 0.015365f
C33 VDD1.n5 VSUBS 0.027006f
C34 VDD1.n6 VSUBS 0.014512f
C35 VDD1.n7 VSUBS 0.0343f
C36 VDD1.n8 VSUBS 0.015365f
C37 VDD1.n9 VSUBS 0.027006f
C38 VDD1.n10 VSUBS 0.014512f
C39 VDD1.n11 VSUBS 0.0343f
C40 VDD1.n12 VSUBS 0.0343f
C41 VDD1.n13 VSUBS 0.015365f
C42 VDD1.n14 VSUBS 0.027006f
C43 VDD1.n15 VSUBS 0.014512f
C44 VDD1.n16 VSUBS 0.0343f
C45 VDD1.n17 VSUBS 0.015365f
C46 VDD1.n18 VSUBS 0.027006f
C47 VDD1.n19 VSUBS 0.014512f
C48 VDD1.n20 VSUBS 0.0343f
C49 VDD1.n21 VSUBS 0.015365f
C50 VDD1.n22 VSUBS 0.027006f
C51 VDD1.n23 VSUBS 0.014512f
C52 VDD1.n24 VSUBS 0.0343f
C53 VDD1.n25 VSUBS 0.015365f
C54 VDD1.n26 VSUBS 0.027006f
C55 VDD1.n27 VSUBS 0.014512f
C56 VDD1.n28 VSUBS 0.0343f
C57 VDD1.n29 VSUBS 0.015365f
C58 VDD1.n30 VSUBS 0.205819f
C59 VDD1.t6 VSUBS 0.07356f
C60 VDD1.n31 VSUBS 0.025725f
C61 VDD1.n32 VSUBS 0.02182f
C62 VDD1.n33 VSUBS 0.014512f
C63 VDD1.n34 VSUBS 1.9622f
C64 VDD1.n35 VSUBS 0.027006f
C65 VDD1.n36 VSUBS 0.014512f
C66 VDD1.n37 VSUBS 0.015365f
C67 VDD1.n38 VSUBS 0.0343f
C68 VDD1.n39 VSUBS 0.0343f
C69 VDD1.n40 VSUBS 0.015365f
C70 VDD1.n41 VSUBS 0.014512f
C71 VDD1.n42 VSUBS 0.027006f
C72 VDD1.n43 VSUBS 0.027006f
C73 VDD1.n44 VSUBS 0.014512f
C74 VDD1.n45 VSUBS 0.015365f
C75 VDD1.n46 VSUBS 0.0343f
C76 VDD1.n47 VSUBS 0.0343f
C77 VDD1.n48 VSUBS 0.015365f
C78 VDD1.n49 VSUBS 0.014512f
C79 VDD1.n50 VSUBS 0.027006f
C80 VDD1.n51 VSUBS 0.027006f
C81 VDD1.n52 VSUBS 0.014512f
C82 VDD1.n53 VSUBS 0.015365f
C83 VDD1.n54 VSUBS 0.0343f
C84 VDD1.n55 VSUBS 0.0343f
C85 VDD1.n56 VSUBS 0.015365f
C86 VDD1.n57 VSUBS 0.014512f
C87 VDD1.n58 VSUBS 0.027006f
C88 VDD1.n59 VSUBS 0.027006f
C89 VDD1.n60 VSUBS 0.014512f
C90 VDD1.n61 VSUBS 0.015365f
C91 VDD1.n62 VSUBS 0.0343f
C92 VDD1.n63 VSUBS 0.0343f
C93 VDD1.n64 VSUBS 0.015365f
C94 VDD1.n65 VSUBS 0.014512f
C95 VDD1.n66 VSUBS 0.027006f
C96 VDD1.n67 VSUBS 0.027006f
C97 VDD1.n68 VSUBS 0.014512f
C98 VDD1.n69 VSUBS 0.015365f
C99 VDD1.n70 VSUBS 0.0343f
C100 VDD1.n71 VSUBS 0.0343f
C101 VDD1.n72 VSUBS 0.015365f
C102 VDD1.n73 VSUBS 0.014512f
C103 VDD1.n74 VSUBS 0.027006f
C104 VDD1.n75 VSUBS 0.027006f
C105 VDD1.n76 VSUBS 0.014512f
C106 VDD1.n77 VSUBS 0.014938f
C107 VDD1.n78 VSUBS 0.014938f
C108 VDD1.n79 VSUBS 0.0343f
C109 VDD1.n80 VSUBS 0.0343f
C110 VDD1.n81 VSUBS 0.015365f
C111 VDD1.n82 VSUBS 0.014512f
C112 VDD1.n83 VSUBS 0.027006f
C113 VDD1.n84 VSUBS 0.027006f
C114 VDD1.n85 VSUBS 0.014512f
C115 VDD1.n86 VSUBS 0.015365f
C116 VDD1.n87 VSUBS 0.0343f
C117 VDD1.n88 VSUBS 0.084992f
C118 VDD1.n89 VSUBS 0.015365f
C119 VDD1.n90 VSUBS 0.014512f
C120 VDD1.n91 VSUBS 0.067587f
C121 VDD1.n92 VSUBS 0.065778f
C122 VDD1.t8 VSUBS 0.361511f
C123 VDD1.t0 VSUBS 0.361511f
C124 VDD1.n93 VSUBS 2.9924f
C125 VDD1.n94 VSUBS 0.828534f
C126 VDD1.n95 VSUBS 0.030247f
C127 VDD1.n96 VSUBS 0.027006f
C128 VDD1.n97 VSUBS 0.014512f
C129 VDD1.n98 VSUBS 0.0343f
C130 VDD1.n99 VSUBS 0.015365f
C131 VDD1.n100 VSUBS 0.027006f
C132 VDD1.n101 VSUBS 0.014512f
C133 VDD1.n102 VSUBS 0.0343f
C134 VDD1.n103 VSUBS 0.015365f
C135 VDD1.n104 VSUBS 0.027006f
C136 VDD1.n105 VSUBS 0.014512f
C137 VDD1.n106 VSUBS 0.0343f
C138 VDD1.n107 VSUBS 0.015365f
C139 VDD1.n108 VSUBS 0.027006f
C140 VDD1.n109 VSUBS 0.014512f
C141 VDD1.n110 VSUBS 0.0343f
C142 VDD1.n111 VSUBS 0.015365f
C143 VDD1.n112 VSUBS 0.027006f
C144 VDD1.n113 VSUBS 0.014512f
C145 VDD1.n114 VSUBS 0.0343f
C146 VDD1.n115 VSUBS 0.015365f
C147 VDD1.n116 VSUBS 0.027006f
C148 VDD1.n117 VSUBS 0.014512f
C149 VDD1.n118 VSUBS 0.0343f
C150 VDD1.n119 VSUBS 0.015365f
C151 VDD1.n120 VSUBS 0.027006f
C152 VDD1.n121 VSUBS 0.014512f
C153 VDD1.n122 VSUBS 0.0343f
C154 VDD1.n123 VSUBS 0.015365f
C155 VDD1.n124 VSUBS 0.205819f
C156 VDD1.t1 VSUBS 0.07356f
C157 VDD1.n125 VSUBS 0.025725f
C158 VDD1.n126 VSUBS 0.02182f
C159 VDD1.n127 VSUBS 0.014512f
C160 VDD1.n128 VSUBS 1.9622f
C161 VDD1.n129 VSUBS 0.027006f
C162 VDD1.n130 VSUBS 0.014512f
C163 VDD1.n131 VSUBS 0.015365f
C164 VDD1.n132 VSUBS 0.0343f
C165 VDD1.n133 VSUBS 0.0343f
C166 VDD1.n134 VSUBS 0.015365f
C167 VDD1.n135 VSUBS 0.014512f
C168 VDD1.n136 VSUBS 0.027006f
C169 VDD1.n137 VSUBS 0.027006f
C170 VDD1.n138 VSUBS 0.014512f
C171 VDD1.n139 VSUBS 0.015365f
C172 VDD1.n140 VSUBS 0.0343f
C173 VDD1.n141 VSUBS 0.0343f
C174 VDD1.n142 VSUBS 0.015365f
C175 VDD1.n143 VSUBS 0.014512f
C176 VDD1.n144 VSUBS 0.027006f
C177 VDD1.n145 VSUBS 0.027006f
C178 VDD1.n146 VSUBS 0.014512f
C179 VDD1.n147 VSUBS 0.015365f
C180 VDD1.n148 VSUBS 0.0343f
C181 VDD1.n149 VSUBS 0.0343f
C182 VDD1.n150 VSUBS 0.015365f
C183 VDD1.n151 VSUBS 0.014512f
C184 VDD1.n152 VSUBS 0.027006f
C185 VDD1.n153 VSUBS 0.027006f
C186 VDD1.n154 VSUBS 0.014512f
C187 VDD1.n155 VSUBS 0.015365f
C188 VDD1.n156 VSUBS 0.0343f
C189 VDD1.n157 VSUBS 0.0343f
C190 VDD1.n158 VSUBS 0.015365f
C191 VDD1.n159 VSUBS 0.014512f
C192 VDD1.n160 VSUBS 0.027006f
C193 VDD1.n161 VSUBS 0.027006f
C194 VDD1.n162 VSUBS 0.014512f
C195 VDD1.n163 VSUBS 0.015365f
C196 VDD1.n164 VSUBS 0.0343f
C197 VDD1.n165 VSUBS 0.0343f
C198 VDD1.n166 VSUBS 0.0343f
C199 VDD1.n167 VSUBS 0.015365f
C200 VDD1.n168 VSUBS 0.014512f
C201 VDD1.n169 VSUBS 0.027006f
C202 VDD1.n170 VSUBS 0.027006f
C203 VDD1.n171 VSUBS 0.014512f
C204 VDD1.n172 VSUBS 0.014938f
C205 VDD1.n173 VSUBS 0.014938f
C206 VDD1.n174 VSUBS 0.0343f
C207 VDD1.n175 VSUBS 0.0343f
C208 VDD1.n176 VSUBS 0.015365f
C209 VDD1.n177 VSUBS 0.014512f
C210 VDD1.n178 VSUBS 0.027006f
C211 VDD1.n179 VSUBS 0.027006f
C212 VDD1.n180 VSUBS 0.014512f
C213 VDD1.n181 VSUBS 0.015365f
C214 VDD1.n182 VSUBS 0.0343f
C215 VDD1.n183 VSUBS 0.084992f
C216 VDD1.n184 VSUBS 0.015365f
C217 VDD1.n185 VSUBS 0.014512f
C218 VDD1.n186 VSUBS 0.067587f
C219 VDD1.n187 VSUBS 0.065778f
C220 VDD1.t5 VSUBS 0.361511f
C221 VDD1.t9 VSUBS 0.361511f
C222 VDD1.n188 VSUBS 2.99239f
C223 VDD1.n189 VSUBS 0.820966f
C224 VDD1.t2 VSUBS 0.361511f
C225 VDD1.t7 VSUBS 0.361511f
C226 VDD1.n190 VSUBS 3.00156f
C227 VDD1.n191 VSUBS 3.05694f
C228 VDD1.t3 VSUBS 0.361511f
C229 VDD1.t4 VSUBS 0.361511f
C230 VDD1.n192 VSUBS 2.99239f
C231 VDD1.n193 VSUBS 3.49952f
C232 VP.n0 VSUBS 0.053494f
C233 VP.t7 VSUBS 2.22022f
C234 VP.n1 VSUBS 0.792003f
C235 VP.n2 VSUBS 0.040089f
C236 VP.t0 VSUBS 2.22022f
C237 VP.n3 VSUBS 0.792003f
C238 VP.n4 VSUBS 0.040089f
C239 VP.t4 VSUBS 2.22022f
C240 VP.n5 VSUBS 0.792003f
C241 VP.n6 VSUBS 0.053494f
C242 VP.n7 VSUBS 0.053494f
C243 VP.t5 VSUBS 2.29375f
C244 VP.t6 VSUBS 2.22022f
C245 VP.n8 VSUBS 0.792003f
C246 VP.n9 VSUBS 0.040089f
C247 VP.t9 VSUBS 2.22022f
C248 VP.n10 VSUBS 0.792003f
C249 VP.n11 VSUBS 0.040089f
C250 VP.t1 VSUBS 2.22022f
C251 VP.n12 VSUBS 0.843156f
C252 VP.t3 VSUBS 2.33466f
C253 VP.n13 VSUBS 0.858885f
C254 VP.n14 VSUBS 0.205306f
C255 VP.n15 VSUBS 0.062616f
C256 VP.n16 VSUBS 0.032493f
C257 VP.n17 VSUBS 0.061945f
C258 VP.n18 VSUBS 0.040089f
C259 VP.n19 VSUBS 0.040089f
C260 VP.n20 VSUBS 0.061945f
C261 VP.n21 VSUBS 0.032493f
C262 VP.n22 VSUBS 0.062616f
C263 VP.n23 VSUBS 0.040089f
C264 VP.n24 VSUBS 0.040089f
C265 VP.n25 VSUBS 0.06105f
C266 VP.n26 VSUBS 0.023508f
C267 VP.n27 VSUBS 0.864574f
C268 VP.n28 VSUBS 2.14773f
C269 VP.n29 VSUBS 2.17688f
C270 VP.t8 VSUBS 2.29375f
C271 VP.n30 VSUBS 0.864574f
C272 VP.n31 VSUBS 0.023508f
C273 VP.n32 VSUBS 0.06105f
C274 VP.n33 VSUBS 0.040089f
C275 VP.n34 VSUBS 0.040089f
C276 VP.n35 VSUBS 0.062616f
C277 VP.n36 VSUBS 0.032493f
C278 VP.n37 VSUBS 0.061945f
C279 VP.n38 VSUBS 0.040089f
C280 VP.n39 VSUBS 0.040089f
C281 VP.n40 VSUBS 0.061945f
C282 VP.n41 VSUBS 0.032493f
C283 VP.n42 VSUBS 0.062616f
C284 VP.n43 VSUBS 0.040089f
C285 VP.n44 VSUBS 0.040089f
C286 VP.n45 VSUBS 0.06105f
C287 VP.n46 VSUBS 0.023508f
C288 VP.t2 VSUBS 2.29375f
C289 VP.n47 VSUBS 0.864574f
C290 VP.n48 VSUBS 0.037545f
C291 B.n0 VSUBS 0.005452f
C292 B.n1 VSUBS 0.005452f
C293 B.n2 VSUBS 0.008622f
C294 B.n3 VSUBS 0.008622f
C295 B.n4 VSUBS 0.008622f
C296 B.n5 VSUBS 0.008622f
C297 B.n6 VSUBS 0.008622f
C298 B.n7 VSUBS 0.008622f
C299 B.n8 VSUBS 0.008622f
C300 B.n9 VSUBS 0.008622f
C301 B.n10 VSUBS 0.008622f
C302 B.n11 VSUBS 0.008622f
C303 B.n12 VSUBS 0.008622f
C304 B.n13 VSUBS 0.008622f
C305 B.n14 VSUBS 0.008622f
C306 B.n15 VSUBS 0.008622f
C307 B.n16 VSUBS 0.008622f
C308 B.n17 VSUBS 0.008622f
C309 B.n18 VSUBS 0.008622f
C310 B.n19 VSUBS 0.019018f
C311 B.n20 VSUBS 0.008622f
C312 B.n21 VSUBS 0.008622f
C313 B.n22 VSUBS 0.008622f
C314 B.n23 VSUBS 0.008622f
C315 B.n24 VSUBS 0.008622f
C316 B.n25 VSUBS 0.008622f
C317 B.n26 VSUBS 0.008622f
C318 B.n27 VSUBS 0.008622f
C319 B.n28 VSUBS 0.008622f
C320 B.n29 VSUBS 0.008622f
C321 B.n30 VSUBS 0.008622f
C322 B.n31 VSUBS 0.008622f
C323 B.n32 VSUBS 0.008622f
C324 B.n33 VSUBS 0.008622f
C325 B.n34 VSUBS 0.008622f
C326 B.n35 VSUBS 0.008622f
C327 B.n36 VSUBS 0.008622f
C328 B.n37 VSUBS 0.008622f
C329 B.n38 VSUBS 0.008622f
C330 B.n39 VSUBS 0.008622f
C331 B.n40 VSUBS 0.008622f
C332 B.n41 VSUBS 0.008622f
C333 B.n42 VSUBS 0.008622f
C334 B.n43 VSUBS 0.008622f
C335 B.n44 VSUBS 0.008622f
C336 B.n45 VSUBS 0.008622f
C337 B.n46 VSUBS 0.008622f
C338 B.n47 VSUBS 0.008622f
C339 B.t2 VSUBS 0.40122f
C340 B.t1 VSUBS 0.423255f
C341 B.t0 VSUBS 1.04166f
C342 B.n48 VSUBS 0.574861f
C343 B.n49 VSUBS 0.381723f
C344 B.n50 VSUBS 0.008622f
C345 B.n51 VSUBS 0.008622f
C346 B.n52 VSUBS 0.008622f
C347 B.n53 VSUBS 0.008622f
C348 B.n54 VSUBS 0.004818f
C349 B.n55 VSUBS 0.008622f
C350 B.t5 VSUBS 0.401225f
C351 B.t4 VSUBS 0.423259f
C352 B.t3 VSUBS 1.04166f
C353 B.n56 VSUBS 0.574857f
C354 B.n57 VSUBS 0.381719f
C355 B.n58 VSUBS 0.019977f
C356 B.n59 VSUBS 0.008622f
C357 B.n60 VSUBS 0.008622f
C358 B.n61 VSUBS 0.008622f
C359 B.n62 VSUBS 0.008622f
C360 B.n63 VSUBS 0.008622f
C361 B.n64 VSUBS 0.008622f
C362 B.n65 VSUBS 0.008622f
C363 B.n66 VSUBS 0.008622f
C364 B.n67 VSUBS 0.008622f
C365 B.n68 VSUBS 0.008622f
C366 B.n69 VSUBS 0.008622f
C367 B.n70 VSUBS 0.008622f
C368 B.n71 VSUBS 0.008622f
C369 B.n72 VSUBS 0.008622f
C370 B.n73 VSUBS 0.008622f
C371 B.n74 VSUBS 0.008622f
C372 B.n75 VSUBS 0.008622f
C373 B.n76 VSUBS 0.008622f
C374 B.n77 VSUBS 0.008622f
C375 B.n78 VSUBS 0.008622f
C376 B.n79 VSUBS 0.008622f
C377 B.n80 VSUBS 0.008622f
C378 B.n81 VSUBS 0.008622f
C379 B.n82 VSUBS 0.008622f
C380 B.n83 VSUBS 0.008622f
C381 B.n84 VSUBS 0.008622f
C382 B.n85 VSUBS 0.018966f
C383 B.n86 VSUBS 0.008622f
C384 B.n87 VSUBS 0.008622f
C385 B.n88 VSUBS 0.008622f
C386 B.n89 VSUBS 0.008622f
C387 B.n90 VSUBS 0.008622f
C388 B.n91 VSUBS 0.008622f
C389 B.n92 VSUBS 0.008622f
C390 B.n93 VSUBS 0.008622f
C391 B.n94 VSUBS 0.008622f
C392 B.n95 VSUBS 0.008622f
C393 B.n96 VSUBS 0.008622f
C394 B.n97 VSUBS 0.008622f
C395 B.n98 VSUBS 0.008622f
C396 B.n99 VSUBS 0.008622f
C397 B.n100 VSUBS 0.008622f
C398 B.n101 VSUBS 0.008622f
C399 B.n102 VSUBS 0.008622f
C400 B.n103 VSUBS 0.008622f
C401 B.n104 VSUBS 0.008622f
C402 B.n105 VSUBS 0.008622f
C403 B.n106 VSUBS 0.008622f
C404 B.n107 VSUBS 0.008622f
C405 B.n108 VSUBS 0.008622f
C406 B.n109 VSUBS 0.008622f
C407 B.n110 VSUBS 0.008622f
C408 B.n111 VSUBS 0.008622f
C409 B.n112 VSUBS 0.008622f
C410 B.n113 VSUBS 0.008622f
C411 B.n114 VSUBS 0.008622f
C412 B.n115 VSUBS 0.008622f
C413 B.n116 VSUBS 0.008622f
C414 B.n117 VSUBS 0.008622f
C415 B.n118 VSUBS 0.008622f
C416 B.n119 VSUBS 0.008622f
C417 B.n120 VSUBS 0.008622f
C418 B.n121 VSUBS 0.020037f
C419 B.n122 VSUBS 0.008622f
C420 B.n123 VSUBS 0.008622f
C421 B.n124 VSUBS 0.008622f
C422 B.n125 VSUBS 0.008622f
C423 B.n126 VSUBS 0.008622f
C424 B.n127 VSUBS 0.008622f
C425 B.n128 VSUBS 0.008622f
C426 B.n129 VSUBS 0.008622f
C427 B.n130 VSUBS 0.008622f
C428 B.n131 VSUBS 0.008622f
C429 B.n132 VSUBS 0.008622f
C430 B.n133 VSUBS 0.008622f
C431 B.n134 VSUBS 0.008622f
C432 B.n135 VSUBS 0.008622f
C433 B.n136 VSUBS 0.008622f
C434 B.n137 VSUBS 0.008622f
C435 B.n138 VSUBS 0.008622f
C436 B.n139 VSUBS 0.008622f
C437 B.n140 VSUBS 0.008622f
C438 B.n141 VSUBS 0.008622f
C439 B.n142 VSUBS 0.008622f
C440 B.n143 VSUBS 0.008622f
C441 B.n144 VSUBS 0.008622f
C442 B.n145 VSUBS 0.008622f
C443 B.n146 VSUBS 0.008622f
C444 B.n147 VSUBS 0.008622f
C445 B.n148 VSUBS 0.008622f
C446 B.t7 VSUBS 0.401225f
C447 B.t8 VSUBS 0.423259f
C448 B.t6 VSUBS 1.04166f
C449 B.n149 VSUBS 0.574857f
C450 B.n150 VSUBS 0.381719f
C451 B.n151 VSUBS 0.019977f
C452 B.n152 VSUBS 0.008622f
C453 B.n153 VSUBS 0.008622f
C454 B.n154 VSUBS 0.008622f
C455 B.n155 VSUBS 0.008622f
C456 B.n156 VSUBS 0.008622f
C457 B.t10 VSUBS 0.40122f
C458 B.t11 VSUBS 0.423255f
C459 B.t9 VSUBS 1.04166f
C460 B.n157 VSUBS 0.574861f
C461 B.n158 VSUBS 0.381723f
C462 B.n159 VSUBS 0.008622f
C463 B.n160 VSUBS 0.008622f
C464 B.n161 VSUBS 0.008622f
C465 B.n162 VSUBS 0.008622f
C466 B.n163 VSUBS 0.008622f
C467 B.n164 VSUBS 0.008622f
C468 B.n165 VSUBS 0.008622f
C469 B.n166 VSUBS 0.008622f
C470 B.n167 VSUBS 0.008622f
C471 B.n168 VSUBS 0.008622f
C472 B.n169 VSUBS 0.008622f
C473 B.n170 VSUBS 0.008622f
C474 B.n171 VSUBS 0.008622f
C475 B.n172 VSUBS 0.008622f
C476 B.n173 VSUBS 0.008622f
C477 B.n174 VSUBS 0.008622f
C478 B.n175 VSUBS 0.008622f
C479 B.n176 VSUBS 0.008622f
C480 B.n177 VSUBS 0.008622f
C481 B.n178 VSUBS 0.008622f
C482 B.n179 VSUBS 0.008622f
C483 B.n180 VSUBS 0.008622f
C484 B.n181 VSUBS 0.008622f
C485 B.n182 VSUBS 0.008622f
C486 B.n183 VSUBS 0.008622f
C487 B.n184 VSUBS 0.008622f
C488 B.n185 VSUBS 0.008622f
C489 B.n186 VSUBS 0.020037f
C490 B.n187 VSUBS 0.008622f
C491 B.n188 VSUBS 0.008622f
C492 B.n189 VSUBS 0.008622f
C493 B.n190 VSUBS 0.008622f
C494 B.n191 VSUBS 0.008622f
C495 B.n192 VSUBS 0.008622f
C496 B.n193 VSUBS 0.008622f
C497 B.n194 VSUBS 0.008622f
C498 B.n195 VSUBS 0.008622f
C499 B.n196 VSUBS 0.008622f
C500 B.n197 VSUBS 0.008622f
C501 B.n198 VSUBS 0.008622f
C502 B.n199 VSUBS 0.008622f
C503 B.n200 VSUBS 0.008622f
C504 B.n201 VSUBS 0.008622f
C505 B.n202 VSUBS 0.008622f
C506 B.n203 VSUBS 0.008622f
C507 B.n204 VSUBS 0.008622f
C508 B.n205 VSUBS 0.008622f
C509 B.n206 VSUBS 0.008622f
C510 B.n207 VSUBS 0.008622f
C511 B.n208 VSUBS 0.008622f
C512 B.n209 VSUBS 0.008622f
C513 B.n210 VSUBS 0.008622f
C514 B.n211 VSUBS 0.008622f
C515 B.n212 VSUBS 0.008622f
C516 B.n213 VSUBS 0.008622f
C517 B.n214 VSUBS 0.008622f
C518 B.n215 VSUBS 0.008622f
C519 B.n216 VSUBS 0.008622f
C520 B.n217 VSUBS 0.008622f
C521 B.n218 VSUBS 0.008622f
C522 B.n219 VSUBS 0.008622f
C523 B.n220 VSUBS 0.008622f
C524 B.n221 VSUBS 0.008622f
C525 B.n222 VSUBS 0.008622f
C526 B.n223 VSUBS 0.008622f
C527 B.n224 VSUBS 0.008622f
C528 B.n225 VSUBS 0.008622f
C529 B.n226 VSUBS 0.008622f
C530 B.n227 VSUBS 0.008622f
C531 B.n228 VSUBS 0.008622f
C532 B.n229 VSUBS 0.008622f
C533 B.n230 VSUBS 0.008622f
C534 B.n231 VSUBS 0.008622f
C535 B.n232 VSUBS 0.008622f
C536 B.n233 VSUBS 0.008622f
C537 B.n234 VSUBS 0.008622f
C538 B.n235 VSUBS 0.008622f
C539 B.n236 VSUBS 0.008622f
C540 B.n237 VSUBS 0.008622f
C541 B.n238 VSUBS 0.008622f
C542 B.n239 VSUBS 0.008622f
C543 B.n240 VSUBS 0.008622f
C544 B.n241 VSUBS 0.008622f
C545 B.n242 VSUBS 0.008622f
C546 B.n243 VSUBS 0.008622f
C547 B.n244 VSUBS 0.008622f
C548 B.n245 VSUBS 0.008622f
C549 B.n246 VSUBS 0.008622f
C550 B.n247 VSUBS 0.008622f
C551 B.n248 VSUBS 0.008622f
C552 B.n249 VSUBS 0.008622f
C553 B.n250 VSUBS 0.008622f
C554 B.n251 VSUBS 0.008622f
C555 B.n252 VSUBS 0.008622f
C556 B.n253 VSUBS 0.019018f
C557 B.n254 VSUBS 0.019018f
C558 B.n255 VSUBS 0.020037f
C559 B.n256 VSUBS 0.008622f
C560 B.n257 VSUBS 0.008622f
C561 B.n258 VSUBS 0.008622f
C562 B.n259 VSUBS 0.008622f
C563 B.n260 VSUBS 0.008622f
C564 B.n261 VSUBS 0.008622f
C565 B.n262 VSUBS 0.008622f
C566 B.n263 VSUBS 0.008622f
C567 B.n264 VSUBS 0.008622f
C568 B.n265 VSUBS 0.008622f
C569 B.n266 VSUBS 0.008622f
C570 B.n267 VSUBS 0.008622f
C571 B.n268 VSUBS 0.008622f
C572 B.n269 VSUBS 0.008622f
C573 B.n270 VSUBS 0.008622f
C574 B.n271 VSUBS 0.008622f
C575 B.n272 VSUBS 0.008622f
C576 B.n273 VSUBS 0.008622f
C577 B.n274 VSUBS 0.008622f
C578 B.n275 VSUBS 0.008622f
C579 B.n276 VSUBS 0.008622f
C580 B.n277 VSUBS 0.008622f
C581 B.n278 VSUBS 0.008622f
C582 B.n279 VSUBS 0.008622f
C583 B.n280 VSUBS 0.008622f
C584 B.n281 VSUBS 0.008622f
C585 B.n282 VSUBS 0.008622f
C586 B.n283 VSUBS 0.008622f
C587 B.n284 VSUBS 0.008622f
C588 B.n285 VSUBS 0.008622f
C589 B.n286 VSUBS 0.008622f
C590 B.n287 VSUBS 0.008622f
C591 B.n288 VSUBS 0.008622f
C592 B.n289 VSUBS 0.008622f
C593 B.n290 VSUBS 0.008622f
C594 B.n291 VSUBS 0.008622f
C595 B.n292 VSUBS 0.008622f
C596 B.n293 VSUBS 0.008622f
C597 B.n294 VSUBS 0.008622f
C598 B.n295 VSUBS 0.008622f
C599 B.n296 VSUBS 0.008622f
C600 B.n297 VSUBS 0.008622f
C601 B.n298 VSUBS 0.008622f
C602 B.n299 VSUBS 0.008622f
C603 B.n300 VSUBS 0.008622f
C604 B.n301 VSUBS 0.008622f
C605 B.n302 VSUBS 0.008622f
C606 B.n303 VSUBS 0.008622f
C607 B.n304 VSUBS 0.008622f
C608 B.n305 VSUBS 0.008622f
C609 B.n306 VSUBS 0.008622f
C610 B.n307 VSUBS 0.008622f
C611 B.n308 VSUBS 0.008622f
C612 B.n309 VSUBS 0.008622f
C613 B.n310 VSUBS 0.008622f
C614 B.n311 VSUBS 0.008622f
C615 B.n312 VSUBS 0.008622f
C616 B.n313 VSUBS 0.008622f
C617 B.n314 VSUBS 0.008622f
C618 B.n315 VSUBS 0.008622f
C619 B.n316 VSUBS 0.008622f
C620 B.n317 VSUBS 0.008622f
C621 B.n318 VSUBS 0.008622f
C622 B.n319 VSUBS 0.008622f
C623 B.n320 VSUBS 0.008622f
C624 B.n321 VSUBS 0.008622f
C625 B.n322 VSUBS 0.008622f
C626 B.n323 VSUBS 0.008622f
C627 B.n324 VSUBS 0.008622f
C628 B.n325 VSUBS 0.008622f
C629 B.n326 VSUBS 0.008622f
C630 B.n327 VSUBS 0.008622f
C631 B.n328 VSUBS 0.008622f
C632 B.n329 VSUBS 0.008622f
C633 B.n330 VSUBS 0.008622f
C634 B.n331 VSUBS 0.008622f
C635 B.n332 VSUBS 0.008622f
C636 B.n333 VSUBS 0.008622f
C637 B.n334 VSUBS 0.008622f
C638 B.n335 VSUBS 0.008622f
C639 B.n336 VSUBS 0.008622f
C640 B.n337 VSUBS 0.008622f
C641 B.n338 VSUBS 0.008115f
C642 B.n339 VSUBS 0.019977f
C643 B.n340 VSUBS 0.004818f
C644 B.n341 VSUBS 0.008622f
C645 B.n342 VSUBS 0.008622f
C646 B.n343 VSUBS 0.008622f
C647 B.n344 VSUBS 0.008622f
C648 B.n345 VSUBS 0.008622f
C649 B.n346 VSUBS 0.008622f
C650 B.n347 VSUBS 0.008622f
C651 B.n348 VSUBS 0.008622f
C652 B.n349 VSUBS 0.008622f
C653 B.n350 VSUBS 0.008622f
C654 B.n351 VSUBS 0.008622f
C655 B.n352 VSUBS 0.008622f
C656 B.n353 VSUBS 0.004818f
C657 B.n354 VSUBS 0.008622f
C658 B.n355 VSUBS 0.008622f
C659 B.n356 VSUBS 0.008115f
C660 B.n357 VSUBS 0.008622f
C661 B.n358 VSUBS 0.008622f
C662 B.n359 VSUBS 0.008622f
C663 B.n360 VSUBS 0.008622f
C664 B.n361 VSUBS 0.008622f
C665 B.n362 VSUBS 0.008622f
C666 B.n363 VSUBS 0.008622f
C667 B.n364 VSUBS 0.008622f
C668 B.n365 VSUBS 0.008622f
C669 B.n366 VSUBS 0.008622f
C670 B.n367 VSUBS 0.008622f
C671 B.n368 VSUBS 0.008622f
C672 B.n369 VSUBS 0.008622f
C673 B.n370 VSUBS 0.008622f
C674 B.n371 VSUBS 0.008622f
C675 B.n372 VSUBS 0.008622f
C676 B.n373 VSUBS 0.008622f
C677 B.n374 VSUBS 0.008622f
C678 B.n375 VSUBS 0.008622f
C679 B.n376 VSUBS 0.008622f
C680 B.n377 VSUBS 0.008622f
C681 B.n378 VSUBS 0.008622f
C682 B.n379 VSUBS 0.008622f
C683 B.n380 VSUBS 0.008622f
C684 B.n381 VSUBS 0.008622f
C685 B.n382 VSUBS 0.008622f
C686 B.n383 VSUBS 0.008622f
C687 B.n384 VSUBS 0.008622f
C688 B.n385 VSUBS 0.008622f
C689 B.n386 VSUBS 0.008622f
C690 B.n387 VSUBS 0.008622f
C691 B.n388 VSUBS 0.008622f
C692 B.n389 VSUBS 0.008622f
C693 B.n390 VSUBS 0.008622f
C694 B.n391 VSUBS 0.008622f
C695 B.n392 VSUBS 0.008622f
C696 B.n393 VSUBS 0.008622f
C697 B.n394 VSUBS 0.008622f
C698 B.n395 VSUBS 0.008622f
C699 B.n396 VSUBS 0.008622f
C700 B.n397 VSUBS 0.008622f
C701 B.n398 VSUBS 0.008622f
C702 B.n399 VSUBS 0.008622f
C703 B.n400 VSUBS 0.008622f
C704 B.n401 VSUBS 0.008622f
C705 B.n402 VSUBS 0.008622f
C706 B.n403 VSUBS 0.008622f
C707 B.n404 VSUBS 0.008622f
C708 B.n405 VSUBS 0.008622f
C709 B.n406 VSUBS 0.008622f
C710 B.n407 VSUBS 0.008622f
C711 B.n408 VSUBS 0.008622f
C712 B.n409 VSUBS 0.008622f
C713 B.n410 VSUBS 0.008622f
C714 B.n411 VSUBS 0.008622f
C715 B.n412 VSUBS 0.008622f
C716 B.n413 VSUBS 0.008622f
C717 B.n414 VSUBS 0.008622f
C718 B.n415 VSUBS 0.008622f
C719 B.n416 VSUBS 0.008622f
C720 B.n417 VSUBS 0.008622f
C721 B.n418 VSUBS 0.008622f
C722 B.n419 VSUBS 0.008622f
C723 B.n420 VSUBS 0.008622f
C724 B.n421 VSUBS 0.008622f
C725 B.n422 VSUBS 0.008622f
C726 B.n423 VSUBS 0.008622f
C727 B.n424 VSUBS 0.008622f
C728 B.n425 VSUBS 0.008622f
C729 B.n426 VSUBS 0.008622f
C730 B.n427 VSUBS 0.008622f
C731 B.n428 VSUBS 0.008622f
C732 B.n429 VSUBS 0.008622f
C733 B.n430 VSUBS 0.008622f
C734 B.n431 VSUBS 0.008622f
C735 B.n432 VSUBS 0.008622f
C736 B.n433 VSUBS 0.008622f
C737 B.n434 VSUBS 0.008622f
C738 B.n435 VSUBS 0.008622f
C739 B.n436 VSUBS 0.008622f
C740 B.n437 VSUBS 0.008622f
C741 B.n438 VSUBS 0.020037f
C742 B.n439 VSUBS 0.019018f
C743 B.n440 VSUBS 0.019018f
C744 B.n441 VSUBS 0.008622f
C745 B.n442 VSUBS 0.008622f
C746 B.n443 VSUBS 0.008622f
C747 B.n444 VSUBS 0.008622f
C748 B.n445 VSUBS 0.008622f
C749 B.n446 VSUBS 0.008622f
C750 B.n447 VSUBS 0.008622f
C751 B.n448 VSUBS 0.008622f
C752 B.n449 VSUBS 0.008622f
C753 B.n450 VSUBS 0.008622f
C754 B.n451 VSUBS 0.008622f
C755 B.n452 VSUBS 0.008622f
C756 B.n453 VSUBS 0.008622f
C757 B.n454 VSUBS 0.008622f
C758 B.n455 VSUBS 0.008622f
C759 B.n456 VSUBS 0.008622f
C760 B.n457 VSUBS 0.008622f
C761 B.n458 VSUBS 0.008622f
C762 B.n459 VSUBS 0.008622f
C763 B.n460 VSUBS 0.008622f
C764 B.n461 VSUBS 0.008622f
C765 B.n462 VSUBS 0.008622f
C766 B.n463 VSUBS 0.008622f
C767 B.n464 VSUBS 0.008622f
C768 B.n465 VSUBS 0.008622f
C769 B.n466 VSUBS 0.008622f
C770 B.n467 VSUBS 0.008622f
C771 B.n468 VSUBS 0.008622f
C772 B.n469 VSUBS 0.008622f
C773 B.n470 VSUBS 0.008622f
C774 B.n471 VSUBS 0.008622f
C775 B.n472 VSUBS 0.008622f
C776 B.n473 VSUBS 0.008622f
C777 B.n474 VSUBS 0.008622f
C778 B.n475 VSUBS 0.008622f
C779 B.n476 VSUBS 0.008622f
C780 B.n477 VSUBS 0.008622f
C781 B.n478 VSUBS 0.008622f
C782 B.n479 VSUBS 0.008622f
C783 B.n480 VSUBS 0.008622f
C784 B.n481 VSUBS 0.008622f
C785 B.n482 VSUBS 0.008622f
C786 B.n483 VSUBS 0.008622f
C787 B.n484 VSUBS 0.008622f
C788 B.n485 VSUBS 0.008622f
C789 B.n486 VSUBS 0.008622f
C790 B.n487 VSUBS 0.008622f
C791 B.n488 VSUBS 0.008622f
C792 B.n489 VSUBS 0.008622f
C793 B.n490 VSUBS 0.008622f
C794 B.n491 VSUBS 0.008622f
C795 B.n492 VSUBS 0.008622f
C796 B.n493 VSUBS 0.008622f
C797 B.n494 VSUBS 0.008622f
C798 B.n495 VSUBS 0.008622f
C799 B.n496 VSUBS 0.008622f
C800 B.n497 VSUBS 0.008622f
C801 B.n498 VSUBS 0.008622f
C802 B.n499 VSUBS 0.008622f
C803 B.n500 VSUBS 0.008622f
C804 B.n501 VSUBS 0.008622f
C805 B.n502 VSUBS 0.008622f
C806 B.n503 VSUBS 0.008622f
C807 B.n504 VSUBS 0.008622f
C808 B.n505 VSUBS 0.008622f
C809 B.n506 VSUBS 0.008622f
C810 B.n507 VSUBS 0.008622f
C811 B.n508 VSUBS 0.008622f
C812 B.n509 VSUBS 0.008622f
C813 B.n510 VSUBS 0.008622f
C814 B.n511 VSUBS 0.008622f
C815 B.n512 VSUBS 0.008622f
C816 B.n513 VSUBS 0.008622f
C817 B.n514 VSUBS 0.008622f
C818 B.n515 VSUBS 0.008622f
C819 B.n516 VSUBS 0.008622f
C820 B.n517 VSUBS 0.008622f
C821 B.n518 VSUBS 0.008622f
C822 B.n519 VSUBS 0.008622f
C823 B.n520 VSUBS 0.008622f
C824 B.n521 VSUBS 0.008622f
C825 B.n522 VSUBS 0.008622f
C826 B.n523 VSUBS 0.008622f
C827 B.n524 VSUBS 0.008622f
C828 B.n525 VSUBS 0.008622f
C829 B.n526 VSUBS 0.008622f
C830 B.n527 VSUBS 0.008622f
C831 B.n528 VSUBS 0.008622f
C832 B.n529 VSUBS 0.008622f
C833 B.n530 VSUBS 0.008622f
C834 B.n531 VSUBS 0.008622f
C835 B.n532 VSUBS 0.008622f
C836 B.n533 VSUBS 0.008622f
C837 B.n534 VSUBS 0.008622f
C838 B.n535 VSUBS 0.008622f
C839 B.n536 VSUBS 0.008622f
C840 B.n537 VSUBS 0.008622f
C841 B.n538 VSUBS 0.008622f
C842 B.n539 VSUBS 0.008622f
C843 B.n540 VSUBS 0.008622f
C844 B.n541 VSUBS 0.008622f
C845 B.n542 VSUBS 0.008622f
C846 B.n543 VSUBS 0.008622f
C847 B.n544 VSUBS 0.020089f
C848 B.n545 VSUBS 0.019018f
C849 B.n546 VSUBS 0.020037f
C850 B.n547 VSUBS 0.008622f
C851 B.n548 VSUBS 0.008622f
C852 B.n549 VSUBS 0.008622f
C853 B.n550 VSUBS 0.008622f
C854 B.n551 VSUBS 0.008622f
C855 B.n552 VSUBS 0.008622f
C856 B.n553 VSUBS 0.008622f
C857 B.n554 VSUBS 0.008622f
C858 B.n555 VSUBS 0.008622f
C859 B.n556 VSUBS 0.008622f
C860 B.n557 VSUBS 0.008622f
C861 B.n558 VSUBS 0.008622f
C862 B.n559 VSUBS 0.008622f
C863 B.n560 VSUBS 0.008622f
C864 B.n561 VSUBS 0.008622f
C865 B.n562 VSUBS 0.008622f
C866 B.n563 VSUBS 0.008622f
C867 B.n564 VSUBS 0.008622f
C868 B.n565 VSUBS 0.008622f
C869 B.n566 VSUBS 0.008622f
C870 B.n567 VSUBS 0.008622f
C871 B.n568 VSUBS 0.008622f
C872 B.n569 VSUBS 0.008622f
C873 B.n570 VSUBS 0.008622f
C874 B.n571 VSUBS 0.008622f
C875 B.n572 VSUBS 0.008622f
C876 B.n573 VSUBS 0.008622f
C877 B.n574 VSUBS 0.008622f
C878 B.n575 VSUBS 0.008622f
C879 B.n576 VSUBS 0.008622f
C880 B.n577 VSUBS 0.008622f
C881 B.n578 VSUBS 0.008622f
C882 B.n579 VSUBS 0.008622f
C883 B.n580 VSUBS 0.008622f
C884 B.n581 VSUBS 0.008622f
C885 B.n582 VSUBS 0.008622f
C886 B.n583 VSUBS 0.008622f
C887 B.n584 VSUBS 0.008622f
C888 B.n585 VSUBS 0.008622f
C889 B.n586 VSUBS 0.008622f
C890 B.n587 VSUBS 0.008622f
C891 B.n588 VSUBS 0.008622f
C892 B.n589 VSUBS 0.008622f
C893 B.n590 VSUBS 0.008622f
C894 B.n591 VSUBS 0.008622f
C895 B.n592 VSUBS 0.008622f
C896 B.n593 VSUBS 0.008622f
C897 B.n594 VSUBS 0.008622f
C898 B.n595 VSUBS 0.008622f
C899 B.n596 VSUBS 0.008622f
C900 B.n597 VSUBS 0.008622f
C901 B.n598 VSUBS 0.008622f
C902 B.n599 VSUBS 0.008622f
C903 B.n600 VSUBS 0.008622f
C904 B.n601 VSUBS 0.008622f
C905 B.n602 VSUBS 0.008622f
C906 B.n603 VSUBS 0.008622f
C907 B.n604 VSUBS 0.008622f
C908 B.n605 VSUBS 0.008622f
C909 B.n606 VSUBS 0.008622f
C910 B.n607 VSUBS 0.008622f
C911 B.n608 VSUBS 0.008622f
C912 B.n609 VSUBS 0.008622f
C913 B.n610 VSUBS 0.008622f
C914 B.n611 VSUBS 0.008622f
C915 B.n612 VSUBS 0.008622f
C916 B.n613 VSUBS 0.008622f
C917 B.n614 VSUBS 0.008622f
C918 B.n615 VSUBS 0.008622f
C919 B.n616 VSUBS 0.008622f
C920 B.n617 VSUBS 0.008622f
C921 B.n618 VSUBS 0.008622f
C922 B.n619 VSUBS 0.008622f
C923 B.n620 VSUBS 0.008622f
C924 B.n621 VSUBS 0.008622f
C925 B.n622 VSUBS 0.008622f
C926 B.n623 VSUBS 0.008622f
C927 B.n624 VSUBS 0.008622f
C928 B.n625 VSUBS 0.008622f
C929 B.n626 VSUBS 0.008622f
C930 B.n627 VSUBS 0.008622f
C931 B.n628 VSUBS 0.008115f
C932 B.n629 VSUBS 0.008622f
C933 B.n630 VSUBS 0.008622f
C934 B.n631 VSUBS 0.008622f
C935 B.n632 VSUBS 0.008622f
C936 B.n633 VSUBS 0.008622f
C937 B.n634 VSUBS 0.008622f
C938 B.n635 VSUBS 0.008622f
C939 B.n636 VSUBS 0.008622f
C940 B.n637 VSUBS 0.008622f
C941 B.n638 VSUBS 0.008622f
C942 B.n639 VSUBS 0.008622f
C943 B.n640 VSUBS 0.008622f
C944 B.n641 VSUBS 0.008622f
C945 B.n642 VSUBS 0.008622f
C946 B.n643 VSUBS 0.008622f
C947 B.n644 VSUBS 0.004818f
C948 B.n645 VSUBS 0.019977f
C949 B.n646 VSUBS 0.008115f
C950 B.n647 VSUBS 0.008622f
C951 B.n648 VSUBS 0.008622f
C952 B.n649 VSUBS 0.008622f
C953 B.n650 VSUBS 0.008622f
C954 B.n651 VSUBS 0.008622f
C955 B.n652 VSUBS 0.008622f
C956 B.n653 VSUBS 0.008622f
C957 B.n654 VSUBS 0.008622f
C958 B.n655 VSUBS 0.008622f
C959 B.n656 VSUBS 0.008622f
C960 B.n657 VSUBS 0.008622f
C961 B.n658 VSUBS 0.008622f
C962 B.n659 VSUBS 0.008622f
C963 B.n660 VSUBS 0.008622f
C964 B.n661 VSUBS 0.008622f
C965 B.n662 VSUBS 0.008622f
C966 B.n663 VSUBS 0.008622f
C967 B.n664 VSUBS 0.008622f
C968 B.n665 VSUBS 0.008622f
C969 B.n666 VSUBS 0.008622f
C970 B.n667 VSUBS 0.008622f
C971 B.n668 VSUBS 0.008622f
C972 B.n669 VSUBS 0.008622f
C973 B.n670 VSUBS 0.008622f
C974 B.n671 VSUBS 0.008622f
C975 B.n672 VSUBS 0.008622f
C976 B.n673 VSUBS 0.008622f
C977 B.n674 VSUBS 0.008622f
C978 B.n675 VSUBS 0.008622f
C979 B.n676 VSUBS 0.008622f
C980 B.n677 VSUBS 0.008622f
C981 B.n678 VSUBS 0.008622f
C982 B.n679 VSUBS 0.008622f
C983 B.n680 VSUBS 0.008622f
C984 B.n681 VSUBS 0.008622f
C985 B.n682 VSUBS 0.008622f
C986 B.n683 VSUBS 0.008622f
C987 B.n684 VSUBS 0.008622f
C988 B.n685 VSUBS 0.008622f
C989 B.n686 VSUBS 0.008622f
C990 B.n687 VSUBS 0.008622f
C991 B.n688 VSUBS 0.008622f
C992 B.n689 VSUBS 0.008622f
C993 B.n690 VSUBS 0.008622f
C994 B.n691 VSUBS 0.008622f
C995 B.n692 VSUBS 0.008622f
C996 B.n693 VSUBS 0.008622f
C997 B.n694 VSUBS 0.008622f
C998 B.n695 VSUBS 0.008622f
C999 B.n696 VSUBS 0.008622f
C1000 B.n697 VSUBS 0.008622f
C1001 B.n698 VSUBS 0.008622f
C1002 B.n699 VSUBS 0.008622f
C1003 B.n700 VSUBS 0.008622f
C1004 B.n701 VSUBS 0.008622f
C1005 B.n702 VSUBS 0.008622f
C1006 B.n703 VSUBS 0.008622f
C1007 B.n704 VSUBS 0.008622f
C1008 B.n705 VSUBS 0.008622f
C1009 B.n706 VSUBS 0.008622f
C1010 B.n707 VSUBS 0.008622f
C1011 B.n708 VSUBS 0.008622f
C1012 B.n709 VSUBS 0.008622f
C1013 B.n710 VSUBS 0.008622f
C1014 B.n711 VSUBS 0.008622f
C1015 B.n712 VSUBS 0.008622f
C1016 B.n713 VSUBS 0.008622f
C1017 B.n714 VSUBS 0.008622f
C1018 B.n715 VSUBS 0.008622f
C1019 B.n716 VSUBS 0.008622f
C1020 B.n717 VSUBS 0.008622f
C1021 B.n718 VSUBS 0.008622f
C1022 B.n719 VSUBS 0.008622f
C1023 B.n720 VSUBS 0.008622f
C1024 B.n721 VSUBS 0.008622f
C1025 B.n722 VSUBS 0.008622f
C1026 B.n723 VSUBS 0.008622f
C1027 B.n724 VSUBS 0.008622f
C1028 B.n725 VSUBS 0.008622f
C1029 B.n726 VSUBS 0.008622f
C1030 B.n727 VSUBS 0.008622f
C1031 B.n728 VSUBS 0.020037f
C1032 B.n729 VSUBS 0.020037f
C1033 B.n730 VSUBS 0.019018f
C1034 B.n731 VSUBS 0.008622f
C1035 B.n732 VSUBS 0.008622f
C1036 B.n733 VSUBS 0.008622f
C1037 B.n734 VSUBS 0.008622f
C1038 B.n735 VSUBS 0.008622f
C1039 B.n736 VSUBS 0.008622f
C1040 B.n737 VSUBS 0.008622f
C1041 B.n738 VSUBS 0.008622f
C1042 B.n739 VSUBS 0.008622f
C1043 B.n740 VSUBS 0.008622f
C1044 B.n741 VSUBS 0.008622f
C1045 B.n742 VSUBS 0.008622f
C1046 B.n743 VSUBS 0.008622f
C1047 B.n744 VSUBS 0.008622f
C1048 B.n745 VSUBS 0.008622f
C1049 B.n746 VSUBS 0.008622f
C1050 B.n747 VSUBS 0.008622f
C1051 B.n748 VSUBS 0.008622f
C1052 B.n749 VSUBS 0.008622f
C1053 B.n750 VSUBS 0.008622f
C1054 B.n751 VSUBS 0.008622f
C1055 B.n752 VSUBS 0.008622f
C1056 B.n753 VSUBS 0.008622f
C1057 B.n754 VSUBS 0.008622f
C1058 B.n755 VSUBS 0.008622f
C1059 B.n756 VSUBS 0.008622f
C1060 B.n757 VSUBS 0.008622f
C1061 B.n758 VSUBS 0.008622f
C1062 B.n759 VSUBS 0.008622f
C1063 B.n760 VSUBS 0.008622f
C1064 B.n761 VSUBS 0.008622f
C1065 B.n762 VSUBS 0.008622f
C1066 B.n763 VSUBS 0.008622f
C1067 B.n764 VSUBS 0.008622f
C1068 B.n765 VSUBS 0.008622f
C1069 B.n766 VSUBS 0.008622f
C1070 B.n767 VSUBS 0.008622f
C1071 B.n768 VSUBS 0.008622f
C1072 B.n769 VSUBS 0.008622f
C1073 B.n770 VSUBS 0.008622f
C1074 B.n771 VSUBS 0.008622f
C1075 B.n772 VSUBS 0.008622f
C1076 B.n773 VSUBS 0.008622f
C1077 B.n774 VSUBS 0.008622f
C1078 B.n775 VSUBS 0.008622f
C1079 B.n776 VSUBS 0.008622f
C1080 B.n777 VSUBS 0.008622f
C1081 B.n778 VSUBS 0.008622f
C1082 B.n779 VSUBS 0.008622f
C1083 B.n780 VSUBS 0.008622f
C1084 B.n781 VSUBS 0.008622f
C1085 B.n782 VSUBS 0.008622f
C1086 B.n783 VSUBS 0.019524f
C1087 VDD2.n0 VSUBS 0.030342f
C1088 VDD2.n1 VSUBS 0.02709f
C1089 VDD2.n2 VSUBS 0.014557f
C1090 VDD2.n3 VSUBS 0.034407f
C1091 VDD2.n4 VSUBS 0.015413f
C1092 VDD2.n5 VSUBS 0.02709f
C1093 VDD2.n6 VSUBS 0.014557f
C1094 VDD2.n7 VSUBS 0.034407f
C1095 VDD2.n8 VSUBS 0.015413f
C1096 VDD2.n9 VSUBS 0.02709f
C1097 VDD2.n10 VSUBS 0.014557f
C1098 VDD2.n11 VSUBS 0.034407f
C1099 VDD2.n12 VSUBS 0.015413f
C1100 VDD2.n13 VSUBS 0.02709f
C1101 VDD2.n14 VSUBS 0.014557f
C1102 VDD2.n15 VSUBS 0.034407f
C1103 VDD2.n16 VSUBS 0.015413f
C1104 VDD2.n17 VSUBS 0.02709f
C1105 VDD2.n18 VSUBS 0.014557f
C1106 VDD2.n19 VSUBS 0.034407f
C1107 VDD2.n20 VSUBS 0.015413f
C1108 VDD2.n21 VSUBS 0.02709f
C1109 VDD2.n22 VSUBS 0.014557f
C1110 VDD2.n23 VSUBS 0.034407f
C1111 VDD2.n24 VSUBS 0.015413f
C1112 VDD2.n25 VSUBS 0.02709f
C1113 VDD2.n26 VSUBS 0.014557f
C1114 VDD2.n27 VSUBS 0.034407f
C1115 VDD2.n28 VSUBS 0.015413f
C1116 VDD2.n29 VSUBS 0.206461f
C1117 VDD2.t6 VSUBS 0.073789f
C1118 VDD2.n30 VSUBS 0.025805f
C1119 VDD2.n31 VSUBS 0.021888f
C1120 VDD2.n32 VSUBS 0.014557f
C1121 VDD2.n33 VSUBS 1.96832f
C1122 VDD2.n34 VSUBS 0.02709f
C1123 VDD2.n35 VSUBS 0.014557f
C1124 VDD2.n36 VSUBS 0.015413f
C1125 VDD2.n37 VSUBS 0.034407f
C1126 VDD2.n38 VSUBS 0.034407f
C1127 VDD2.n39 VSUBS 0.015413f
C1128 VDD2.n40 VSUBS 0.014557f
C1129 VDD2.n41 VSUBS 0.02709f
C1130 VDD2.n42 VSUBS 0.02709f
C1131 VDD2.n43 VSUBS 0.014557f
C1132 VDD2.n44 VSUBS 0.015413f
C1133 VDD2.n45 VSUBS 0.034407f
C1134 VDD2.n46 VSUBS 0.034407f
C1135 VDD2.n47 VSUBS 0.015413f
C1136 VDD2.n48 VSUBS 0.014557f
C1137 VDD2.n49 VSUBS 0.02709f
C1138 VDD2.n50 VSUBS 0.02709f
C1139 VDD2.n51 VSUBS 0.014557f
C1140 VDD2.n52 VSUBS 0.015413f
C1141 VDD2.n53 VSUBS 0.034407f
C1142 VDD2.n54 VSUBS 0.034407f
C1143 VDD2.n55 VSUBS 0.015413f
C1144 VDD2.n56 VSUBS 0.014557f
C1145 VDD2.n57 VSUBS 0.02709f
C1146 VDD2.n58 VSUBS 0.02709f
C1147 VDD2.n59 VSUBS 0.014557f
C1148 VDD2.n60 VSUBS 0.015413f
C1149 VDD2.n61 VSUBS 0.034407f
C1150 VDD2.n62 VSUBS 0.034407f
C1151 VDD2.n63 VSUBS 0.015413f
C1152 VDD2.n64 VSUBS 0.014557f
C1153 VDD2.n65 VSUBS 0.02709f
C1154 VDD2.n66 VSUBS 0.02709f
C1155 VDD2.n67 VSUBS 0.014557f
C1156 VDD2.n68 VSUBS 0.015413f
C1157 VDD2.n69 VSUBS 0.034407f
C1158 VDD2.n70 VSUBS 0.034407f
C1159 VDD2.n71 VSUBS 0.034407f
C1160 VDD2.n72 VSUBS 0.015413f
C1161 VDD2.n73 VSUBS 0.014557f
C1162 VDD2.n74 VSUBS 0.02709f
C1163 VDD2.n75 VSUBS 0.02709f
C1164 VDD2.n76 VSUBS 0.014557f
C1165 VDD2.n77 VSUBS 0.014985f
C1166 VDD2.n78 VSUBS 0.014985f
C1167 VDD2.n79 VSUBS 0.034407f
C1168 VDD2.n80 VSUBS 0.034407f
C1169 VDD2.n81 VSUBS 0.015413f
C1170 VDD2.n82 VSUBS 0.014557f
C1171 VDD2.n83 VSUBS 0.02709f
C1172 VDD2.n84 VSUBS 0.02709f
C1173 VDD2.n85 VSUBS 0.014557f
C1174 VDD2.n86 VSUBS 0.015413f
C1175 VDD2.n87 VSUBS 0.034407f
C1176 VDD2.n88 VSUBS 0.085257f
C1177 VDD2.n89 VSUBS 0.015413f
C1178 VDD2.n90 VSUBS 0.014557f
C1179 VDD2.n91 VSUBS 0.067798f
C1180 VDD2.n92 VSUBS 0.065983f
C1181 VDD2.t3 VSUBS 0.362638f
C1182 VDD2.t8 VSUBS 0.362638f
C1183 VDD2.n93 VSUBS 3.00172f
C1184 VDD2.n94 VSUBS 0.823525f
C1185 VDD2.t5 VSUBS 0.362638f
C1186 VDD2.t1 VSUBS 0.362638f
C1187 VDD2.n95 VSUBS 3.01092f
C1188 VDD2.n96 VSUBS 2.96827f
C1189 VDD2.n97 VSUBS 0.030342f
C1190 VDD2.n98 VSUBS 0.02709f
C1191 VDD2.n99 VSUBS 0.014557f
C1192 VDD2.n100 VSUBS 0.034407f
C1193 VDD2.n101 VSUBS 0.015413f
C1194 VDD2.n102 VSUBS 0.02709f
C1195 VDD2.n103 VSUBS 0.014557f
C1196 VDD2.n104 VSUBS 0.034407f
C1197 VDD2.n105 VSUBS 0.015413f
C1198 VDD2.n106 VSUBS 0.02709f
C1199 VDD2.n107 VSUBS 0.014557f
C1200 VDD2.n108 VSUBS 0.034407f
C1201 VDD2.n109 VSUBS 0.034407f
C1202 VDD2.n110 VSUBS 0.015413f
C1203 VDD2.n111 VSUBS 0.02709f
C1204 VDD2.n112 VSUBS 0.014557f
C1205 VDD2.n113 VSUBS 0.034407f
C1206 VDD2.n114 VSUBS 0.015413f
C1207 VDD2.n115 VSUBS 0.02709f
C1208 VDD2.n116 VSUBS 0.014557f
C1209 VDD2.n117 VSUBS 0.034407f
C1210 VDD2.n118 VSUBS 0.015413f
C1211 VDD2.n119 VSUBS 0.02709f
C1212 VDD2.n120 VSUBS 0.014557f
C1213 VDD2.n121 VSUBS 0.034407f
C1214 VDD2.n122 VSUBS 0.015413f
C1215 VDD2.n123 VSUBS 0.02709f
C1216 VDD2.n124 VSUBS 0.014557f
C1217 VDD2.n125 VSUBS 0.034407f
C1218 VDD2.n126 VSUBS 0.015413f
C1219 VDD2.n127 VSUBS 0.206461f
C1220 VDD2.t2 VSUBS 0.073789f
C1221 VDD2.n128 VSUBS 0.025805f
C1222 VDD2.n129 VSUBS 0.021888f
C1223 VDD2.n130 VSUBS 0.014557f
C1224 VDD2.n131 VSUBS 1.96832f
C1225 VDD2.n132 VSUBS 0.02709f
C1226 VDD2.n133 VSUBS 0.014557f
C1227 VDD2.n134 VSUBS 0.015413f
C1228 VDD2.n135 VSUBS 0.034407f
C1229 VDD2.n136 VSUBS 0.034407f
C1230 VDD2.n137 VSUBS 0.015413f
C1231 VDD2.n138 VSUBS 0.014557f
C1232 VDD2.n139 VSUBS 0.02709f
C1233 VDD2.n140 VSUBS 0.02709f
C1234 VDD2.n141 VSUBS 0.014557f
C1235 VDD2.n142 VSUBS 0.015413f
C1236 VDD2.n143 VSUBS 0.034407f
C1237 VDD2.n144 VSUBS 0.034407f
C1238 VDD2.n145 VSUBS 0.015413f
C1239 VDD2.n146 VSUBS 0.014557f
C1240 VDD2.n147 VSUBS 0.02709f
C1241 VDD2.n148 VSUBS 0.02709f
C1242 VDD2.n149 VSUBS 0.014557f
C1243 VDD2.n150 VSUBS 0.015413f
C1244 VDD2.n151 VSUBS 0.034407f
C1245 VDD2.n152 VSUBS 0.034407f
C1246 VDD2.n153 VSUBS 0.015413f
C1247 VDD2.n154 VSUBS 0.014557f
C1248 VDD2.n155 VSUBS 0.02709f
C1249 VDD2.n156 VSUBS 0.02709f
C1250 VDD2.n157 VSUBS 0.014557f
C1251 VDD2.n158 VSUBS 0.015413f
C1252 VDD2.n159 VSUBS 0.034407f
C1253 VDD2.n160 VSUBS 0.034407f
C1254 VDD2.n161 VSUBS 0.015413f
C1255 VDD2.n162 VSUBS 0.014557f
C1256 VDD2.n163 VSUBS 0.02709f
C1257 VDD2.n164 VSUBS 0.02709f
C1258 VDD2.n165 VSUBS 0.014557f
C1259 VDD2.n166 VSUBS 0.015413f
C1260 VDD2.n167 VSUBS 0.034407f
C1261 VDD2.n168 VSUBS 0.034407f
C1262 VDD2.n169 VSUBS 0.015413f
C1263 VDD2.n170 VSUBS 0.014557f
C1264 VDD2.n171 VSUBS 0.02709f
C1265 VDD2.n172 VSUBS 0.02709f
C1266 VDD2.n173 VSUBS 0.014557f
C1267 VDD2.n174 VSUBS 0.014985f
C1268 VDD2.n175 VSUBS 0.014985f
C1269 VDD2.n176 VSUBS 0.034407f
C1270 VDD2.n177 VSUBS 0.034407f
C1271 VDD2.n178 VSUBS 0.015413f
C1272 VDD2.n179 VSUBS 0.014557f
C1273 VDD2.n180 VSUBS 0.02709f
C1274 VDD2.n181 VSUBS 0.02709f
C1275 VDD2.n182 VSUBS 0.014557f
C1276 VDD2.n183 VSUBS 0.015413f
C1277 VDD2.n184 VSUBS 0.034407f
C1278 VDD2.n185 VSUBS 0.085257f
C1279 VDD2.n186 VSUBS 0.015413f
C1280 VDD2.n187 VSUBS 0.014557f
C1281 VDD2.n188 VSUBS 0.067798f
C1282 VDD2.n189 VSUBS 0.061783f
C1283 VDD2.n190 VSUBS 2.95432f
C1284 VDD2.t0 VSUBS 0.362638f
C1285 VDD2.t9 VSUBS 0.362638f
C1286 VDD2.n191 VSUBS 3.00173f
C1287 VDD2.n192 VSUBS 0.665806f
C1288 VDD2.t7 VSUBS 0.362638f
C1289 VDD2.t4 VSUBS 0.362638f
C1290 VDD2.n193 VSUBS 3.01088f
C1291 VTAIL.t12 VSUBS 0.365429f
C1292 VTAIL.t8 VSUBS 0.365429f
C1293 VTAIL.n0 VSUBS 2.86939f
C1294 VTAIL.n1 VSUBS 0.830604f
C1295 VTAIL.n2 VSUBS 0.030575f
C1296 VTAIL.n3 VSUBS 0.027298f
C1297 VTAIL.n4 VSUBS 0.014669f
C1298 VTAIL.n5 VSUBS 0.034672f
C1299 VTAIL.n6 VSUBS 0.015532f
C1300 VTAIL.n7 VSUBS 0.027298f
C1301 VTAIL.n8 VSUBS 0.014669f
C1302 VTAIL.n9 VSUBS 0.034672f
C1303 VTAIL.n10 VSUBS 0.015532f
C1304 VTAIL.n11 VSUBS 0.027298f
C1305 VTAIL.n12 VSUBS 0.014669f
C1306 VTAIL.n13 VSUBS 0.034672f
C1307 VTAIL.n14 VSUBS 0.015532f
C1308 VTAIL.n15 VSUBS 0.027298f
C1309 VTAIL.n16 VSUBS 0.014669f
C1310 VTAIL.n17 VSUBS 0.034672f
C1311 VTAIL.n18 VSUBS 0.015532f
C1312 VTAIL.n19 VSUBS 0.027298f
C1313 VTAIL.n20 VSUBS 0.014669f
C1314 VTAIL.n21 VSUBS 0.034672f
C1315 VTAIL.n22 VSUBS 0.015532f
C1316 VTAIL.n23 VSUBS 0.027298f
C1317 VTAIL.n24 VSUBS 0.014669f
C1318 VTAIL.n25 VSUBS 0.034672f
C1319 VTAIL.n26 VSUBS 0.015532f
C1320 VTAIL.n27 VSUBS 0.027298f
C1321 VTAIL.n28 VSUBS 0.014669f
C1322 VTAIL.n29 VSUBS 0.034672f
C1323 VTAIL.n30 VSUBS 0.015532f
C1324 VTAIL.n31 VSUBS 0.20805f
C1325 VTAIL.t4 VSUBS 0.074357f
C1326 VTAIL.n32 VSUBS 0.026004f
C1327 VTAIL.n33 VSUBS 0.022057f
C1328 VTAIL.n34 VSUBS 0.014669f
C1329 VTAIL.n35 VSUBS 1.98347f
C1330 VTAIL.n36 VSUBS 0.027298f
C1331 VTAIL.n37 VSUBS 0.014669f
C1332 VTAIL.n38 VSUBS 0.015532f
C1333 VTAIL.n39 VSUBS 0.034672f
C1334 VTAIL.n40 VSUBS 0.034672f
C1335 VTAIL.n41 VSUBS 0.015532f
C1336 VTAIL.n42 VSUBS 0.014669f
C1337 VTAIL.n43 VSUBS 0.027298f
C1338 VTAIL.n44 VSUBS 0.027298f
C1339 VTAIL.n45 VSUBS 0.014669f
C1340 VTAIL.n46 VSUBS 0.015532f
C1341 VTAIL.n47 VSUBS 0.034672f
C1342 VTAIL.n48 VSUBS 0.034672f
C1343 VTAIL.n49 VSUBS 0.015532f
C1344 VTAIL.n50 VSUBS 0.014669f
C1345 VTAIL.n51 VSUBS 0.027298f
C1346 VTAIL.n52 VSUBS 0.027298f
C1347 VTAIL.n53 VSUBS 0.014669f
C1348 VTAIL.n54 VSUBS 0.015532f
C1349 VTAIL.n55 VSUBS 0.034672f
C1350 VTAIL.n56 VSUBS 0.034672f
C1351 VTAIL.n57 VSUBS 0.015532f
C1352 VTAIL.n58 VSUBS 0.014669f
C1353 VTAIL.n59 VSUBS 0.027298f
C1354 VTAIL.n60 VSUBS 0.027298f
C1355 VTAIL.n61 VSUBS 0.014669f
C1356 VTAIL.n62 VSUBS 0.015532f
C1357 VTAIL.n63 VSUBS 0.034672f
C1358 VTAIL.n64 VSUBS 0.034672f
C1359 VTAIL.n65 VSUBS 0.015532f
C1360 VTAIL.n66 VSUBS 0.014669f
C1361 VTAIL.n67 VSUBS 0.027298f
C1362 VTAIL.n68 VSUBS 0.027298f
C1363 VTAIL.n69 VSUBS 0.014669f
C1364 VTAIL.n70 VSUBS 0.015532f
C1365 VTAIL.n71 VSUBS 0.034672f
C1366 VTAIL.n72 VSUBS 0.034672f
C1367 VTAIL.n73 VSUBS 0.034672f
C1368 VTAIL.n74 VSUBS 0.015532f
C1369 VTAIL.n75 VSUBS 0.014669f
C1370 VTAIL.n76 VSUBS 0.027298f
C1371 VTAIL.n77 VSUBS 0.027298f
C1372 VTAIL.n78 VSUBS 0.014669f
C1373 VTAIL.n79 VSUBS 0.0151f
C1374 VTAIL.n80 VSUBS 0.0151f
C1375 VTAIL.n81 VSUBS 0.034672f
C1376 VTAIL.n82 VSUBS 0.034672f
C1377 VTAIL.n83 VSUBS 0.015532f
C1378 VTAIL.n84 VSUBS 0.014669f
C1379 VTAIL.n85 VSUBS 0.027298f
C1380 VTAIL.n86 VSUBS 0.027298f
C1381 VTAIL.n87 VSUBS 0.014669f
C1382 VTAIL.n88 VSUBS 0.015532f
C1383 VTAIL.n89 VSUBS 0.034672f
C1384 VTAIL.n90 VSUBS 0.085913f
C1385 VTAIL.n91 VSUBS 0.015532f
C1386 VTAIL.n92 VSUBS 0.014669f
C1387 VTAIL.n93 VSUBS 0.06832f
C1388 VTAIL.n94 VSUBS 0.043448f
C1389 VTAIL.n95 VSUBS 0.240483f
C1390 VTAIL.t5 VSUBS 0.365429f
C1391 VTAIL.t19 VSUBS 0.365429f
C1392 VTAIL.n96 VSUBS 2.86939f
C1393 VTAIL.n97 VSUBS 0.870603f
C1394 VTAIL.t3 VSUBS 0.365429f
C1395 VTAIL.t18 VSUBS 0.365429f
C1396 VTAIL.n98 VSUBS 2.86939f
C1397 VTAIL.n99 VSUBS 2.64122f
C1398 VTAIL.t17 VSUBS 0.365429f
C1399 VTAIL.t14 VSUBS 0.365429f
C1400 VTAIL.n100 VSUBS 2.86941f
C1401 VTAIL.n101 VSUBS 2.6412f
C1402 VTAIL.t11 VSUBS 0.365429f
C1403 VTAIL.t10 VSUBS 0.365429f
C1404 VTAIL.n102 VSUBS 2.86941f
C1405 VTAIL.n103 VSUBS 0.870586f
C1406 VTAIL.n104 VSUBS 0.030575f
C1407 VTAIL.n105 VSUBS 0.027298f
C1408 VTAIL.n106 VSUBS 0.014669f
C1409 VTAIL.n107 VSUBS 0.034672f
C1410 VTAIL.n108 VSUBS 0.015532f
C1411 VTAIL.n109 VSUBS 0.027298f
C1412 VTAIL.n110 VSUBS 0.014669f
C1413 VTAIL.n111 VSUBS 0.034672f
C1414 VTAIL.n112 VSUBS 0.015532f
C1415 VTAIL.n113 VSUBS 0.027298f
C1416 VTAIL.n114 VSUBS 0.014669f
C1417 VTAIL.n115 VSUBS 0.034672f
C1418 VTAIL.n116 VSUBS 0.034672f
C1419 VTAIL.n117 VSUBS 0.015532f
C1420 VTAIL.n118 VSUBS 0.027298f
C1421 VTAIL.n119 VSUBS 0.014669f
C1422 VTAIL.n120 VSUBS 0.034672f
C1423 VTAIL.n121 VSUBS 0.015532f
C1424 VTAIL.n122 VSUBS 0.027298f
C1425 VTAIL.n123 VSUBS 0.014669f
C1426 VTAIL.n124 VSUBS 0.034672f
C1427 VTAIL.n125 VSUBS 0.015532f
C1428 VTAIL.n126 VSUBS 0.027298f
C1429 VTAIL.n127 VSUBS 0.014669f
C1430 VTAIL.n128 VSUBS 0.034672f
C1431 VTAIL.n129 VSUBS 0.015532f
C1432 VTAIL.n130 VSUBS 0.027298f
C1433 VTAIL.n131 VSUBS 0.014669f
C1434 VTAIL.n132 VSUBS 0.034672f
C1435 VTAIL.n133 VSUBS 0.015532f
C1436 VTAIL.n134 VSUBS 0.20805f
C1437 VTAIL.t16 VSUBS 0.074357f
C1438 VTAIL.n135 VSUBS 0.026004f
C1439 VTAIL.n136 VSUBS 0.022057f
C1440 VTAIL.n137 VSUBS 0.014669f
C1441 VTAIL.n138 VSUBS 1.98347f
C1442 VTAIL.n139 VSUBS 0.027298f
C1443 VTAIL.n140 VSUBS 0.014669f
C1444 VTAIL.n141 VSUBS 0.015532f
C1445 VTAIL.n142 VSUBS 0.034672f
C1446 VTAIL.n143 VSUBS 0.034672f
C1447 VTAIL.n144 VSUBS 0.015532f
C1448 VTAIL.n145 VSUBS 0.014669f
C1449 VTAIL.n146 VSUBS 0.027298f
C1450 VTAIL.n147 VSUBS 0.027298f
C1451 VTAIL.n148 VSUBS 0.014669f
C1452 VTAIL.n149 VSUBS 0.015532f
C1453 VTAIL.n150 VSUBS 0.034672f
C1454 VTAIL.n151 VSUBS 0.034672f
C1455 VTAIL.n152 VSUBS 0.015532f
C1456 VTAIL.n153 VSUBS 0.014669f
C1457 VTAIL.n154 VSUBS 0.027298f
C1458 VTAIL.n155 VSUBS 0.027298f
C1459 VTAIL.n156 VSUBS 0.014669f
C1460 VTAIL.n157 VSUBS 0.015532f
C1461 VTAIL.n158 VSUBS 0.034672f
C1462 VTAIL.n159 VSUBS 0.034672f
C1463 VTAIL.n160 VSUBS 0.015532f
C1464 VTAIL.n161 VSUBS 0.014669f
C1465 VTAIL.n162 VSUBS 0.027298f
C1466 VTAIL.n163 VSUBS 0.027298f
C1467 VTAIL.n164 VSUBS 0.014669f
C1468 VTAIL.n165 VSUBS 0.015532f
C1469 VTAIL.n166 VSUBS 0.034672f
C1470 VTAIL.n167 VSUBS 0.034672f
C1471 VTAIL.n168 VSUBS 0.015532f
C1472 VTAIL.n169 VSUBS 0.014669f
C1473 VTAIL.n170 VSUBS 0.027298f
C1474 VTAIL.n171 VSUBS 0.027298f
C1475 VTAIL.n172 VSUBS 0.014669f
C1476 VTAIL.n173 VSUBS 0.015532f
C1477 VTAIL.n174 VSUBS 0.034672f
C1478 VTAIL.n175 VSUBS 0.034672f
C1479 VTAIL.n176 VSUBS 0.015532f
C1480 VTAIL.n177 VSUBS 0.014669f
C1481 VTAIL.n178 VSUBS 0.027298f
C1482 VTAIL.n179 VSUBS 0.027298f
C1483 VTAIL.n180 VSUBS 0.014669f
C1484 VTAIL.n181 VSUBS 0.0151f
C1485 VTAIL.n182 VSUBS 0.0151f
C1486 VTAIL.n183 VSUBS 0.034672f
C1487 VTAIL.n184 VSUBS 0.034672f
C1488 VTAIL.n185 VSUBS 0.015532f
C1489 VTAIL.n186 VSUBS 0.014669f
C1490 VTAIL.n187 VSUBS 0.027298f
C1491 VTAIL.n188 VSUBS 0.027298f
C1492 VTAIL.n189 VSUBS 0.014669f
C1493 VTAIL.n190 VSUBS 0.015532f
C1494 VTAIL.n191 VSUBS 0.034672f
C1495 VTAIL.n192 VSUBS 0.085913f
C1496 VTAIL.n193 VSUBS 0.015532f
C1497 VTAIL.n194 VSUBS 0.014669f
C1498 VTAIL.n195 VSUBS 0.06832f
C1499 VTAIL.n196 VSUBS 0.043448f
C1500 VTAIL.n197 VSUBS 0.240483f
C1501 VTAIL.t0 VSUBS 0.365429f
C1502 VTAIL.t7 VSUBS 0.365429f
C1503 VTAIL.n198 VSUBS 2.86941f
C1504 VTAIL.n199 VSUBS 0.854283f
C1505 VTAIL.t1 VSUBS 0.365429f
C1506 VTAIL.t2 VSUBS 0.365429f
C1507 VTAIL.n200 VSUBS 2.86941f
C1508 VTAIL.n201 VSUBS 0.870586f
C1509 VTAIL.n202 VSUBS 0.030575f
C1510 VTAIL.n203 VSUBS 0.027298f
C1511 VTAIL.n204 VSUBS 0.014669f
C1512 VTAIL.n205 VSUBS 0.034672f
C1513 VTAIL.n206 VSUBS 0.015532f
C1514 VTAIL.n207 VSUBS 0.027298f
C1515 VTAIL.n208 VSUBS 0.014669f
C1516 VTAIL.n209 VSUBS 0.034672f
C1517 VTAIL.n210 VSUBS 0.015532f
C1518 VTAIL.n211 VSUBS 0.027298f
C1519 VTAIL.n212 VSUBS 0.014669f
C1520 VTAIL.n213 VSUBS 0.034672f
C1521 VTAIL.n214 VSUBS 0.034672f
C1522 VTAIL.n215 VSUBS 0.015532f
C1523 VTAIL.n216 VSUBS 0.027298f
C1524 VTAIL.n217 VSUBS 0.014669f
C1525 VTAIL.n218 VSUBS 0.034672f
C1526 VTAIL.n219 VSUBS 0.015532f
C1527 VTAIL.n220 VSUBS 0.027298f
C1528 VTAIL.n221 VSUBS 0.014669f
C1529 VTAIL.n222 VSUBS 0.034672f
C1530 VTAIL.n223 VSUBS 0.015532f
C1531 VTAIL.n224 VSUBS 0.027298f
C1532 VTAIL.n225 VSUBS 0.014669f
C1533 VTAIL.n226 VSUBS 0.034672f
C1534 VTAIL.n227 VSUBS 0.015532f
C1535 VTAIL.n228 VSUBS 0.027298f
C1536 VTAIL.n229 VSUBS 0.014669f
C1537 VTAIL.n230 VSUBS 0.034672f
C1538 VTAIL.n231 VSUBS 0.015532f
C1539 VTAIL.n232 VSUBS 0.20805f
C1540 VTAIL.t6 VSUBS 0.074357f
C1541 VTAIL.n233 VSUBS 0.026004f
C1542 VTAIL.n234 VSUBS 0.022057f
C1543 VTAIL.n235 VSUBS 0.014669f
C1544 VTAIL.n236 VSUBS 1.98347f
C1545 VTAIL.n237 VSUBS 0.027298f
C1546 VTAIL.n238 VSUBS 0.014669f
C1547 VTAIL.n239 VSUBS 0.015532f
C1548 VTAIL.n240 VSUBS 0.034672f
C1549 VTAIL.n241 VSUBS 0.034672f
C1550 VTAIL.n242 VSUBS 0.015532f
C1551 VTAIL.n243 VSUBS 0.014669f
C1552 VTAIL.n244 VSUBS 0.027298f
C1553 VTAIL.n245 VSUBS 0.027298f
C1554 VTAIL.n246 VSUBS 0.014669f
C1555 VTAIL.n247 VSUBS 0.015532f
C1556 VTAIL.n248 VSUBS 0.034672f
C1557 VTAIL.n249 VSUBS 0.034672f
C1558 VTAIL.n250 VSUBS 0.015532f
C1559 VTAIL.n251 VSUBS 0.014669f
C1560 VTAIL.n252 VSUBS 0.027298f
C1561 VTAIL.n253 VSUBS 0.027298f
C1562 VTAIL.n254 VSUBS 0.014669f
C1563 VTAIL.n255 VSUBS 0.015532f
C1564 VTAIL.n256 VSUBS 0.034672f
C1565 VTAIL.n257 VSUBS 0.034672f
C1566 VTAIL.n258 VSUBS 0.015532f
C1567 VTAIL.n259 VSUBS 0.014669f
C1568 VTAIL.n260 VSUBS 0.027298f
C1569 VTAIL.n261 VSUBS 0.027298f
C1570 VTAIL.n262 VSUBS 0.014669f
C1571 VTAIL.n263 VSUBS 0.015532f
C1572 VTAIL.n264 VSUBS 0.034672f
C1573 VTAIL.n265 VSUBS 0.034672f
C1574 VTAIL.n266 VSUBS 0.015532f
C1575 VTAIL.n267 VSUBS 0.014669f
C1576 VTAIL.n268 VSUBS 0.027298f
C1577 VTAIL.n269 VSUBS 0.027298f
C1578 VTAIL.n270 VSUBS 0.014669f
C1579 VTAIL.n271 VSUBS 0.015532f
C1580 VTAIL.n272 VSUBS 0.034672f
C1581 VTAIL.n273 VSUBS 0.034672f
C1582 VTAIL.n274 VSUBS 0.015532f
C1583 VTAIL.n275 VSUBS 0.014669f
C1584 VTAIL.n276 VSUBS 0.027298f
C1585 VTAIL.n277 VSUBS 0.027298f
C1586 VTAIL.n278 VSUBS 0.014669f
C1587 VTAIL.n279 VSUBS 0.0151f
C1588 VTAIL.n280 VSUBS 0.0151f
C1589 VTAIL.n281 VSUBS 0.034672f
C1590 VTAIL.n282 VSUBS 0.034672f
C1591 VTAIL.n283 VSUBS 0.015532f
C1592 VTAIL.n284 VSUBS 0.014669f
C1593 VTAIL.n285 VSUBS 0.027298f
C1594 VTAIL.n286 VSUBS 0.027298f
C1595 VTAIL.n287 VSUBS 0.014669f
C1596 VTAIL.n288 VSUBS 0.015532f
C1597 VTAIL.n289 VSUBS 0.034672f
C1598 VTAIL.n290 VSUBS 0.085913f
C1599 VTAIL.n291 VSUBS 0.015532f
C1600 VTAIL.n292 VSUBS 0.014669f
C1601 VTAIL.n293 VSUBS 0.06832f
C1602 VTAIL.n294 VSUBS 0.043448f
C1603 VTAIL.n295 VSUBS 1.91214f
C1604 VTAIL.n296 VSUBS 0.030575f
C1605 VTAIL.n297 VSUBS 0.027298f
C1606 VTAIL.n298 VSUBS 0.014669f
C1607 VTAIL.n299 VSUBS 0.034672f
C1608 VTAIL.n300 VSUBS 0.015532f
C1609 VTAIL.n301 VSUBS 0.027298f
C1610 VTAIL.n302 VSUBS 0.014669f
C1611 VTAIL.n303 VSUBS 0.034672f
C1612 VTAIL.n304 VSUBS 0.015532f
C1613 VTAIL.n305 VSUBS 0.027298f
C1614 VTAIL.n306 VSUBS 0.014669f
C1615 VTAIL.n307 VSUBS 0.034672f
C1616 VTAIL.n308 VSUBS 0.015532f
C1617 VTAIL.n309 VSUBS 0.027298f
C1618 VTAIL.n310 VSUBS 0.014669f
C1619 VTAIL.n311 VSUBS 0.034672f
C1620 VTAIL.n312 VSUBS 0.015532f
C1621 VTAIL.n313 VSUBS 0.027298f
C1622 VTAIL.n314 VSUBS 0.014669f
C1623 VTAIL.n315 VSUBS 0.034672f
C1624 VTAIL.n316 VSUBS 0.015532f
C1625 VTAIL.n317 VSUBS 0.027298f
C1626 VTAIL.n318 VSUBS 0.014669f
C1627 VTAIL.n319 VSUBS 0.034672f
C1628 VTAIL.n320 VSUBS 0.015532f
C1629 VTAIL.n321 VSUBS 0.027298f
C1630 VTAIL.n322 VSUBS 0.014669f
C1631 VTAIL.n323 VSUBS 0.034672f
C1632 VTAIL.n324 VSUBS 0.015532f
C1633 VTAIL.n325 VSUBS 0.20805f
C1634 VTAIL.t15 VSUBS 0.074357f
C1635 VTAIL.n326 VSUBS 0.026004f
C1636 VTAIL.n327 VSUBS 0.022057f
C1637 VTAIL.n328 VSUBS 0.014669f
C1638 VTAIL.n329 VSUBS 1.98347f
C1639 VTAIL.n330 VSUBS 0.027298f
C1640 VTAIL.n331 VSUBS 0.014669f
C1641 VTAIL.n332 VSUBS 0.015532f
C1642 VTAIL.n333 VSUBS 0.034672f
C1643 VTAIL.n334 VSUBS 0.034672f
C1644 VTAIL.n335 VSUBS 0.015532f
C1645 VTAIL.n336 VSUBS 0.014669f
C1646 VTAIL.n337 VSUBS 0.027298f
C1647 VTAIL.n338 VSUBS 0.027298f
C1648 VTAIL.n339 VSUBS 0.014669f
C1649 VTAIL.n340 VSUBS 0.015532f
C1650 VTAIL.n341 VSUBS 0.034672f
C1651 VTAIL.n342 VSUBS 0.034672f
C1652 VTAIL.n343 VSUBS 0.015532f
C1653 VTAIL.n344 VSUBS 0.014669f
C1654 VTAIL.n345 VSUBS 0.027298f
C1655 VTAIL.n346 VSUBS 0.027298f
C1656 VTAIL.n347 VSUBS 0.014669f
C1657 VTAIL.n348 VSUBS 0.015532f
C1658 VTAIL.n349 VSUBS 0.034672f
C1659 VTAIL.n350 VSUBS 0.034672f
C1660 VTAIL.n351 VSUBS 0.015532f
C1661 VTAIL.n352 VSUBS 0.014669f
C1662 VTAIL.n353 VSUBS 0.027298f
C1663 VTAIL.n354 VSUBS 0.027298f
C1664 VTAIL.n355 VSUBS 0.014669f
C1665 VTAIL.n356 VSUBS 0.015532f
C1666 VTAIL.n357 VSUBS 0.034672f
C1667 VTAIL.n358 VSUBS 0.034672f
C1668 VTAIL.n359 VSUBS 0.015532f
C1669 VTAIL.n360 VSUBS 0.014669f
C1670 VTAIL.n361 VSUBS 0.027298f
C1671 VTAIL.n362 VSUBS 0.027298f
C1672 VTAIL.n363 VSUBS 0.014669f
C1673 VTAIL.n364 VSUBS 0.015532f
C1674 VTAIL.n365 VSUBS 0.034672f
C1675 VTAIL.n366 VSUBS 0.034672f
C1676 VTAIL.n367 VSUBS 0.034672f
C1677 VTAIL.n368 VSUBS 0.015532f
C1678 VTAIL.n369 VSUBS 0.014669f
C1679 VTAIL.n370 VSUBS 0.027298f
C1680 VTAIL.n371 VSUBS 0.027298f
C1681 VTAIL.n372 VSUBS 0.014669f
C1682 VTAIL.n373 VSUBS 0.0151f
C1683 VTAIL.n374 VSUBS 0.0151f
C1684 VTAIL.n375 VSUBS 0.034672f
C1685 VTAIL.n376 VSUBS 0.034672f
C1686 VTAIL.n377 VSUBS 0.015532f
C1687 VTAIL.n378 VSUBS 0.014669f
C1688 VTAIL.n379 VSUBS 0.027298f
C1689 VTAIL.n380 VSUBS 0.027298f
C1690 VTAIL.n381 VSUBS 0.014669f
C1691 VTAIL.n382 VSUBS 0.015532f
C1692 VTAIL.n383 VSUBS 0.034672f
C1693 VTAIL.n384 VSUBS 0.085913f
C1694 VTAIL.n385 VSUBS 0.015532f
C1695 VTAIL.n386 VSUBS 0.014669f
C1696 VTAIL.n387 VSUBS 0.06832f
C1697 VTAIL.n388 VSUBS 0.043448f
C1698 VTAIL.n389 VSUBS 1.91214f
C1699 VTAIL.t9 VSUBS 0.365429f
C1700 VTAIL.t13 VSUBS 0.365429f
C1701 VTAIL.n390 VSUBS 2.86939f
C1702 VTAIL.n391 VSUBS 0.77904f
C1703 VN.n0 VSUBS 0.052691f
C1704 VN.t4 VSUBS 2.18689f
C1705 VN.n1 VSUBS 0.780112f
C1706 VN.n2 VSUBS 0.039487f
C1707 VN.t1 VSUBS 2.18689f
C1708 VN.n3 VSUBS 0.780112f
C1709 VN.n4 VSUBS 0.039487f
C1710 VN.t6 VSUBS 2.18689f
C1711 VN.n5 VSUBS 0.830497f
C1712 VN.t3 VSUBS 2.29961f
C1713 VN.n6 VSUBS 0.84599f
C1714 VN.n7 VSUBS 0.202223f
C1715 VN.n8 VSUBS 0.061676f
C1716 VN.n9 VSUBS 0.032005f
C1717 VN.n10 VSUBS 0.061015f
C1718 VN.n11 VSUBS 0.039487f
C1719 VN.n12 VSUBS 0.039487f
C1720 VN.n13 VSUBS 0.061015f
C1721 VN.n14 VSUBS 0.032005f
C1722 VN.n15 VSUBS 0.061676f
C1723 VN.n16 VSUBS 0.039487f
C1724 VN.n17 VSUBS 0.039487f
C1725 VN.n18 VSUBS 0.060133f
C1726 VN.n19 VSUBS 0.023155f
C1727 VN.t8 VSUBS 2.25931f
C1728 VN.n20 VSUBS 0.851593f
C1729 VN.n21 VSUBS 0.036981f
C1730 VN.n22 VSUBS 0.052691f
C1731 VN.t9 VSUBS 2.18689f
C1732 VN.n23 VSUBS 0.780112f
C1733 VN.n24 VSUBS 0.039487f
C1734 VN.t0 VSUBS 2.18689f
C1735 VN.n25 VSUBS 0.780112f
C1736 VN.n26 VSUBS 0.039487f
C1737 VN.t2 VSUBS 2.18689f
C1738 VN.n27 VSUBS 0.830497f
C1739 VN.t5 VSUBS 2.29961f
C1740 VN.n28 VSUBS 0.84599f
C1741 VN.n29 VSUBS 0.202223f
C1742 VN.n30 VSUBS 0.061676f
C1743 VN.n31 VSUBS 0.032005f
C1744 VN.n32 VSUBS 0.061015f
C1745 VN.n33 VSUBS 0.039487f
C1746 VN.n34 VSUBS 0.039487f
C1747 VN.n35 VSUBS 0.061015f
C1748 VN.n36 VSUBS 0.032005f
C1749 VN.n37 VSUBS 0.061676f
C1750 VN.n38 VSUBS 0.039487f
C1751 VN.n39 VSUBS 0.039487f
C1752 VN.n40 VSUBS 0.060133f
C1753 VN.n41 VSUBS 0.023155f
C1754 VN.t7 VSUBS 2.25931f
C1755 VN.n42 VSUBS 0.851593f
C1756 VN.n43 VSUBS 2.13707f
.ends

