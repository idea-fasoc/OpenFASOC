* NGSPICE file created from diff_pair_sample_0241.ext - technology: sky130A

.subckt diff_pair_sample_0241 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t14 w_n4510_n2178# sky130_fd_pr__pfet_01v8 ad=0.99825 pd=6.38 as=0.99825 ps=6.38 w=6.05 l=3.21
X1 B.t11 B.t9 B.t10 w_n4510_n2178# sky130_fd_pr__pfet_01v8 ad=2.3595 pd=12.88 as=0 ps=0 w=6.05 l=3.21
X2 VDD2.t7 VN.t0 VTAIL.t4 w_n4510_n2178# sky130_fd_pr__pfet_01v8 ad=0.99825 pd=6.38 as=0.99825 ps=6.38 w=6.05 l=3.21
X3 VTAIL.t15 VP.t1 VDD1.t6 w_n4510_n2178# sky130_fd_pr__pfet_01v8 ad=0.99825 pd=6.38 as=0.99825 ps=6.38 w=6.05 l=3.21
X4 VTAIL.t2 VN.t1 VDD2.t6 w_n4510_n2178# sky130_fd_pr__pfet_01v8 ad=2.3595 pd=12.88 as=0.99825 ps=6.38 w=6.05 l=3.21
X5 VDD1.t5 VP.t2 VTAIL.t12 w_n4510_n2178# sky130_fd_pr__pfet_01v8 ad=0.99825 pd=6.38 as=0.99825 ps=6.38 w=6.05 l=3.21
X6 B.t8 B.t6 B.t7 w_n4510_n2178# sky130_fd_pr__pfet_01v8 ad=2.3595 pd=12.88 as=0 ps=0 w=6.05 l=3.21
X7 VDD2.t5 VN.t2 VTAIL.t7 w_n4510_n2178# sky130_fd_pr__pfet_01v8 ad=0.99825 pd=6.38 as=2.3595 ps=12.88 w=6.05 l=3.21
X8 B.t5 B.t3 B.t4 w_n4510_n2178# sky130_fd_pr__pfet_01v8 ad=2.3595 pd=12.88 as=0 ps=0 w=6.05 l=3.21
X9 VTAIL.t8 VP.t3 VDD1.t4 w_n4510_n2178# sky130_fd_pr__pfet_01v8 ad=0.99825 pd=6.38 as=0.99825 ps=6.38 w=6.05 l=3.21
X10 VTAIL.t5 VN.t3 VDD2.t4 w_n4510_n2178# sky130_fd_pr__pfet_01v8 ad=0.99825 pd=6.38 as=0.99825 ps=6.38 w=6.05 l=3.21
X11 VDD2.t3 VN.t4 VTAIL.t1 w_n4510_n2178# sky130_fd_pr__pfet_01v8 ad=0.99825 pd=6.38 as=2.3595 ps=12.88 w=6.05 l=3.21
X12 VDD2.t2 VN.t5 VTAIL.t3 w_n4510_n2178# sky130_fd_pr__pfet_01v8 ad=0.99825 pd=6.38 as=0.99825 ps=6.38 w=6.05 l=3.21
X13 VDD1.t3 VP.t4 VTAIL.t10 w_n4510_n2178# sky130_fd_pr__pfet_01v8 ad=0.99825 pd=6.38 as=2.3595 ps=12.88 w=6.05 l=3.21
X14 VTAIL.t6 VN.t6 VDD2.t1 w_n4510_n2178# sky130_fd_pr__pfet_01v8 ad=0.99825 pd=6.38 as=0.99825 ps=6.38 w=6.05 l=3.21
X15 B.t2 B.t0 B.t1 w_n4510_n2178# sky130_fd_pr__pfet_01v8 ad=2.3595 pd=12.88 as=0 ps=0 w=6.05 l=3.21
X16 VDD1.t2 VP.t5 VTAIL.t9 w_n4510_n2178# sky130_fd_pr__pfet_01v8 ad=0.99825 pd=6.38 as=2.3595 ps=12.88 w=6.05 l=3.21
X17 VTAIL.t13 VP.t6 VDD1.t1 w_n4510_n2178# sky130_fd_pr__pfet_01v8 ad=2.3595 pd=12.88 as=0.99825 ps=6.38 w=6.05 l=3.21
X18 VTAIL.t11 VP.t7 VDD1.t0 w_n4510_n2178# sky130_fd_pr__pfet_01v8 ad=2.3595 pd=12.88 as=0.99825 ps=6.38 w=6.05 l=3.21
X19 VTAIL.t0 VN.t7 VDD2.t0 w_n4510_n2178# sky130_fd_pr__pfet_01v8 ad=2.3595 pd=12.88 as=0.99825 ps=6.38 w=6.05 l=3.21
R0 VP.n24 VP.n23 161.3
R1 VP.n25 VP.n20 161.3
R2 VP.n27 VP.n26 161.3
R3 VP.n28 VP.n19 161.3
R4 VP.n30 VP.n29 161.3
R5 VP.n31 VP.n18 161.3
R6 VP.n33 VP.n32 161.3
R7 VP.n35 VP.n34 161.3
R8 VP.n36 VP.n16 161.3
R9 VP.n38 VP.n37 161.3
R10 VP.n39 VP.n15 161.3
R11 VP.n41 VP.n40 161.3
R12 VP.n42 VP.n14 161.3
R13 VP.n44 VP.n43 161.3
R14 VP.n79 VP.n78 161.3
R15 VP.n77 VP.n1 161.3
R16 VP.n76 VP.n75 161.3
R17 VP.n74 VP.n2 161.3
R18 VP.n73 VP.n72 161.3
R19 VP.n71 VP.n3 161.3
R20 VP.n70 VP.n69 161.3
R21 VP.n68 VP.n67 161.3
R22 VP.n66 VP.n5 161.3
R23 VP.n65 VP.n64 161.3
R24 VP.n63 VP.n6 161.3
R25 VP.n62 VP.n61 161.3
R26 VP.n60 VP.n7 161.3
R27 VP.n59 VP.n58 161.3
R28 VP.n57 VP.n56 161.3
R29 VP.n55 VP.n9 161.3
R30 VP.n54 VP.n53 161.3
R31 VP.n52 VP.n10 161.3
R32 VP.n51 VP.n50 161.3
R33 VP.n49 VP.n11 161.3
R34 VP.n48 VP.n47 161.3
R35 VP.n22 VP.t6 78.4386
R36 VP.n46 VP.n12 74.8979
R37 VP.n80 VP.n0 74.8979
R38 VP.n45 VP.n13 74.8979
R39 VP.n22 VP.n21 61.0251
R40 VP.n46 VP.n45 49.3402
R41 VP.n12 VP.t7 45.4226
R42 VP.n8 VP.t2 45.4226
R43 VP.n4 VP.t3 45.4226
R44 VP.n0 VP.t5 45.4226
R45 VP.n13 VP.t4 45.4226
R46 VP.n17 VP.t1 45.4226
R47 VP.n21 VP.t0 45.4226
R48 VP.n50 VP.n10 44.3785
R49 VP.n76 VP.n2 44.3785
R50 VP.n41 VP.n15 44.3785
R51 VP.n61 VP.n6 40.4934
R52 VP.n65 VP.n6 40.4934
R53 VP.n30 VP.n19 40.4934
R54 VP.n26 VP.n19 40.4934
R55 VP.n54 VP.n10 36.6083
R56 VP.n72 VP.n2 36.6083
R57 VP.n37 VP.n15 36.6083
R58 VP.n49 VP.n48 24.4675
R59 VP.n50 VP.n49 24.4675
R60 VP.n55 VP.n54 24.4675
R61 VP.n56 VP.n55 24.4675
R62 VP.n60 VP.n59 24.4675
R63 VP.n61 VP.n60 24.4675
R64 VP.n66 VP.n65 24.4675
R65 VP.n67 VP.n66 24.4675
R66 VP.n71 VP.n70 24.4675
R67 VP.n72 VP.n71 24.4675
R68 VP.n77 VP.n76 24.4675
R69 VP.n78 VP.n77 24.4675
R70 VP.n42 VP.n41 24.4675
R71 VP.n43 VP.n42 24.4675
R72 VP.n31 VP.n30 24.4675
R73 VP.n32 VP.n31 24.4675
R74 VP.n36 VP.n35 24.4675
R75 VP.n37 VP.n36 24.4675
R76 VP.n25 VP.n24 24.4675
R77 VP.n26 VP.n25 24.4675
R78 VP.n48 VP.n12 15.17
R79 VP.n78 VP.n0 15.17
R80 VP.n43 VP.n13 15.17
R81 VP.n59 VP.n8 13.2127
R82 VP.n67 VP.n4 13.2127
R83 VP.n32 VP.n17 13.2127
R84 VP.n24 VP.n21 13.2127
R85 VP.n56 VP.n8 11.2553
R86 VP.n70 VP.n4 11.2553
R87 VP.n35 VP.n17 11.2553
R88 VP.n23 VP.n22 4.13479
R89 VP.n45 VP.n44 0.354971
R90 VP.n47 VP.n46 0.354971
R91 VP.n80 VP.n79 0.354971
R92 VP VP.n80 0.26696
R93 VP.n23 VP.n20 0.189894
R94 VP.n27 VP.n20 0.189894
R95 VP.n28 VP.n27 0.189894
R96 VP.n29 VP.n28 0.189894
R97 VP.n29 VP.n18 0.189894
R98 VP.n33 VP.n18 0.189894
R99 VP.n34 VP.n33 0.189894
R100 VP.n34 VP.n16 0.189894
R101 VP.n38 VP.n16 0.189894
R102 VP.n39 VP.n38 0.189894
R103 VP.n40 VP.n39 0.189894
R104 VP.n40 VP.n14 0.189894
R105 VP.n44 VP.n14 0.189894
R106 VP.n47 VP.n11 0.189894
R107 VP.n51 VP.n11 0.189894
R108 VP.n52 VP.n51 0.189894
R109 VP.n53 VP.n52 0.189894
R110 VP.n53 VP.n9 0.189894
R111 VP.n57 VP.n9 0.189894
R112 VP.n58 VP.n57 0.189894
R113 VP.n58 VP.n7 0.189894
R114 VP.n62 VP.n7 0.189894
R115 VP.n63 VP.n62 0.189894
R116 VP.n64 VP.n63 0.189894
R117 VP.n64 VP.n5 0.189894
R118 VP.n68 VP.n5 0.189894
R119 VP.n69 VP.n68 0.189894
R120 VP.n69 VP.n3 0.189894
R121 VP.n73 VP.n3 0.189894
R122 VP.n74 VP.n73 0.189894
R123 VP.n75 VP.n74 0.189894
R124 VP.n75 VP.n1 0.189894
R125 VP.n79 VP.n1 0.189894
R126 VTAIL.n258 VTAIL.n232 756.745
R127 VTAIL.n28 VTAIL.n2 756.745
R128 VTAIL.n60 VTAIL.n34 756.745
R129 VTAIL.n94 VTAIL.n68 756.745
R130 VTAIL.n226 VTAIL.n200 756.745
R131 VTAIL.n192 VTAIL.n166 756.745
R132 VTAIL.n160 VTAIL.n134 756.745
R133 VTAIL.n126 VTAIL.n100 756.745
R134 VTAIL.n243 VTAIL.n242 585
R135 VTAIL.n240 VTAIL.n239 585
R136 VTAIL.n249 VTAIL.n248 585
R137 VTAIL.n251 VTAIL.n250 585
R138 VTAIL.n236 VTAIL.n235 585
R139 VTAIL.n257 VTAIL.n256 585
R140 VTAIL.n259 VTAIL.n258 585
R141 VTAIL.n13 VTAIL.n12 585
R142 VTAIL.n10 VTAIL.n9 585
R143 VTAIL.n19 VTAIL.n18 585
R144 VTAIL.n21 VTAIL.n20 585
R145 VTAIL.n6 VTAIL.n5 585
R146 VTAIL.n27 VTAIL.n26 585
R147 VTAIL.n29 VTAIL.n28 585
R148 VTAIL.n45 VTAIL.n44 585
R149 VTAIL.n42 VTAIL.n41 585
R150 VTAIL.n51 VTAIL.n50 585
R151 VTAIL.n53 VTAIL.n52 585
R152 VTAIL.n38 VTAIL.n37 585
R153 VTAIL.n59 VTAIL.n58 585
R154 VTAIL.n61 VTAIL.n60 585
R155 VTAIL.n79 VTAIL.n78 585
R156 VTAIL.n76 VTAIL.n75 585
R157 VTAIL.n85 VTAIL.n84 585
R158 VTAIL.n87 VTAIL.n86 585
R159 VTAIL.n72 VTAIL.n71 585
R160 VTAIL.n93 VTAIL.n92 585
R161 VTAIL.n95 VTAIL.n94 585
R162 VTAIL.n227 VTAIL.n226 585
R163 VTAIL.n225 VTAIL.n224 585
R164 VTAIL.n204 VTAIL.n203 585
R165 VTAIL.n219 VTAIL.n218 585
R166 VTAIL.n217 VTAIL.n216 585
R167 VTAIL.n208 VTAIL.n207 585
R168 VTAIL.n211 VTAIL.n210 585
R169 VTAIL.n193 VTAIL.n192 585
R170 VTAIL.n191 VTAIL.n190 585
R171 VTAIL.n170 VTAIL.n169 585
R172 VTAIL.n185 VTAIL.n184 585
R173 VTAIL.n183 VTAIL.n182 585
R174 VTAIL.n174 VTAIL.n173 585
R175 VTAIL.n177 VTAIL.n176 585
R176 VTAIL.n161 VTAIL.n160 585
R177 VTAIL.n159 VTAIL.n158 585
R178 VTAIL.n138 VTAIL.n137 585
R179 VTAIL.n153 VTAIL.n152 585
R180 VTAIL.n151 VTAIL.n150 585
R181 VTAIL.n142 VTAIL.n141 585
R182 VTAIL.n145 VTAIL.n144 585
R183 VTAIL.n127 VTAIL.n126 585
R184 VTAIL.n125 VTAIL.n124 585
R185 VTAIL.n104 VTAIL.n103 585
R186 VTAIL.n119 VTAIL.n118 585
R187 VTAIL.n117 VTAIL.n116 585
R188 VTAIL.n108 VTAIL.n107 585
R189 VTAIL.n111 VTAIL.n110 585
R190 VTAIL.t1 VTAIL.n241 327.601
R191 VTAIL.t0 VTAIL.n11 327.601
R192 VTAIL.t9 VTAIL.n43 327.601
R193 VTAIL.t11 VTAIL.n77 327.601
R194 VTAIL.t10 VTAIL.n209 327.601
R195 VTAIL.t13 VTAIL.n175 327.601
R196 VTAIL.t7 VTAIL.n143 327.601
R197 VTAIL.t2 VTAIL.n109 327.601
R198 VTAIL.n242 VTAIL.n239 171.744
R199 VTAIL.n249 VTAIL.n239 171.744
R200 VTAIL.n250 VTAIL.n249 171.744
R201 VTAIL.n250 VTAIL.n235 171.744
R202 VTAIL.n257 VTAIL.n235 171.744
R203 VTAIL.n258 VTAIL.n257 171.744
R204 VTAIL.n12 VTAIL.n9 171.744
R205 VTAIL.n19 VTAIL.n9 171.744
R206 VTAIL.n20 VTAIL.n19 171.744
R207 VTAIL.n20 VTAIL.n5 171.744
R208 VTAIL.n27 VTAIL.n5 171.744
R209 VTAIL.n28 VTAIL.n27 171.744
R210 VTAIL.n44 VTAIL.n41 171.744
R211 VTAIL.n51 VTAIL.n41 171.744
R212 VTAIL.n52 VTAIL.n51 171.744
R213 VTAIL.n52 VTAIL.n37 171.744
R214 VTAIL.n59 VTAIL.n37 171.744
R215 VTAIL.n60 VTAIL.n59 171.744
R216 VTAIL.n78 VTAIL.n75 171.744
R217 VTAIL.n85 VTAIL.n75 171.744
R218 VTAIL.n86 VTAIL.n85 171.744
R219 VTAIL.n86 VTAIL.n71 171.744
R220 VTAIL.n93 VTAIL.n71 171.744
R221 VTAIL.n94 VTAIL.n93 171.744
R222 VTAIL.n226 VTAIL.n225 171.744
R223 VTAIL.n225 VTAIL.n203 171.744
R224 VTAIL.n218 VTAIL.n203 171.744
R225 VTAIL.n218 VTAIL.n217 171.744
R226 VTAIL.n217 VTAIL.n207 171.744
R227 VTAIL.n210 VTAIL.n207 171.744
R228 VTAIL.n192 VTAIL.n191 171.744
R229 VTAIL.n191 VTAIL.n169 171.744
R230 VTAIL.n184 VTAIL.n169 171.744
R231 VTAIL.n184 VTAIL.n183 171.744
R232 VTAIL.n183 VTAIL.n173 171.744
R233 VTAIL.n176 VTAIL.n173 171.744
R234 VTAIL.n160 VTAIL.n159 171.744
R235 VTAIL.n159 VTAIL.n137 171.744
R236 VTAIL.n152 VTAIL.n137 171.744
R237 VTAIL.n152 VTAIL.n151 171.744
R238 VTAIL.n151 VTAIL.n141 171.744
R239 VTAIL.n144 VTAIL.n141 171.744
R240 VTAIL.n126 VTAIL.n125 171.744
R241 VTAIL.n125 VTAIL.n103 171.744
R242 VTAIL.n118 VTAIL.n103 171.744
R243 VTAIL.n118 VTAIL.n117 171.744
R244 VTAIL.n117 VTAIL.n107 171.744
R245 VTAIL.n110 VTAIL.n107 171.744
R246 VTAIL.n242 VTAIL.t1 85.8723
R247 VTAIL.n12 VTAIL.t0 85.8723
R248 VTAIL.n44 VTAIL.t9 85.8723
R249 VTAIL.n78 VTAIL.t11 85.8723
R250 VTAIL.n210 VTAIL.t10 85.8723
R251 VTAIL.n176 VTAIL.t13 85.8723
R252 VTAIL.n144 VTAIL.t7 85.8723
R253 VTAIL.n110 VTAIL.t2 85.8723
R254 VTAIL.n199 VTAIL.n198 76.5852
R255 VTAIL.n133 VTAIL.n132 76.5852
R256 VTAIL.n1 VTAIL.n0 76.585
R257 VTAIL.n67 VTAIL.n66 76.585
R258 VTAIL.n263 VTAIL.n262 33.155
R259 VTAIL.n33 VTAIL.n32 33.155
R260 VTAIL.n65 VTAIL.n64 33.155
R261 VTAIL.n99 VTAIL.n98 33.155
R262 VTAIL.n231 VTAIL.n230 33.155
R263 VTAIL.n197 VTAIL.n196 33.155
R264 VTAIL.n165 VTAIL.n164 33.155
R265 VTAIL.n131 VTAIL.n130 33.155
R266 VTAIL.n263 VTAIL.n231 20.6341
R267 VTAIL.n131 VTAIL.n99 20.6341
R268 VTAIL.n243 VTAIL.n241 16.3865
R269 VTAIL.n13 VTAIL.n11 16.3865
R270 VTAIL.n45 VTAIL.n43 16.3865
R271 VTAIL.n79 VTAIL.n77 16.3865
R272 VTAIL.n211 VTAIL.n209 16.3865
R273 VTAIL.n177 VTAIL.n175 16.3865
R274 VTAIL.n145 VTAIL.n143 16.3865
R275 VTAIL.n111 VTAIL.n109 16.3865
R276 VTAIL.n244 VTAIL.n240 12.8005
R277 VTAIL.n14 VTAIL.n10 12.8005
R278 VTAIL.n46 VTAIL.n42 12.8005
R279 VTAIL.n80 VTAIL.n76 12.8005
R280 VTAIL.n212 VTAIL.n208 12.8005
R281 VTAIL.n178 VTAIL.n174 12.8005
R282 VTAIL.n146 VTAIL.n142 12.8005
R283 VTAIL.n112 VTAIL.n108 12.8005
R284 VTAIL.n248 VTAIL.n247 12.0247
R285 VTAIL.n18 VTAIL.n17 12.0247
R286 VTAIL.n50 VTAIL.n49 12.0247
R287 VTAIL.n84 VTAIL.n83 12.0247
R288 VTAIL.n216 VTAIL.n215 12.0247
R289 VTAIL.n182 VTAIL.n181 12.0247
R290 VTAIL.n150 VTAIL.n149 12.0247
R291 VTAIL.n116 VTAIL.n115 12.0247
R292 VTAIL.n251 VTAIL.n238 11.249
R293 VTAIL.n21 VTAIL.n8 11.249
R294 VTAIL.n53 VTAIL.n40 11.249
R295 VTAIL.n87 VTAIL.n74 11.249
R296 VTAIL.n219 VTAIL.n206 11.249
R297 VTAIL.n185 VTAIL.n172 11.249
R298 VTAIL.n153 VTAIL.n140 11.249
R299 VTAIL.n119 VTAIL.n106 11.249
R300 VTAIL.n252 VTAIL.n236 10.4732
R301 VTAIL.n22 VTAIL.n6 10.4732
R302 VTAIL.n54 VTAIL.n38 10.4732
R303 VTAIL.n88 VTAIL.n72 10.4732
R304 VTAIL.n220 VTAIL.n204 10.4732
R305 VTAIL.n186 VTAIL.n170 10.4732
R306 VTAIL.n154 VTAIL.n138 10.4732
R307 VTAIL.n120 VTAIL.n104 10.4732
R308 VTAIL.n256 VTAIL.n255 9.69747
R309 VTAIL.n26 VTAIL.n25 9.69747
R310 VTAIL.n58 VTAIL.n57 9.69747
R311 VTAIL.n92 VTAIL.n91 9.69747
R312 VTAIL.n224 VTAIL.n223 9.69747
R313 VTAIL.n190 VTAIL.n189 9.69747
R314 VTAIL.n158 VTAIL.n157 9.69747
R315 VTAIL.n124 VTAIL.n123 9.69747
R316 VTAIL.n262 VTAIL.n261 9.45567
R317 VTAIL.n32 VTAIL.n31 9.45567
R318 VTAIL.n64 VTAIL.n63 9.45567
R319 VTAIL.n98 VTAIL.n97 9.45567
R320 VTAIL.n230 VTAIL.n229 9.45567
R321 VTAIL.n196 VTAIL.n195 9.45567
R322 VTAIL.n164 VTAIL.n163 9.45567
R323 VTAIL.n130 VTAIL.n129 9.45567
R324 VTAIL.n261 VTAIL.n260 9.3005
R325 VTAIL.n234 VTAIL.n233 9.3005
R326 VTAIL.n255 VTAIL.n254 9.3005
R327 VTAIL.n253 VTAIL.n252 9.3005
R328 VTAIL.n238 VTAIL.n237 9.3005
R329 VTAIL.n247 VTAIL.n246 9.3005
R330 VTAIL.n245 VTAIL.n244 9.3005
R331 VTAIL.n31 VTAIL.n30 9.3005
R332 VTAIL.n4 VTAIL.n3 9.3005
R333 VTAIL.n25 VTAIL.n24 9.3005
R334 VTAIL.n23 VTAIL.n22 9.3005
R335 VTAIL.n8 VTAIL.n7 9.3005
R336 VTAIL.n17 VTAIL.n16 9.3005
R337 VTAIL.n15 VTAIL.n14 9.3005
R338 VTAIL.n63 VTAIL.n62 9.3005
R339 VTAIL.n36 VTAIL.n35 9.3005
R340 VTAIL.n57 VTAIL.n56 9.3005
R341 VTAIL.n55 VTAIL.n54 9.3005
R342 VTAIL.n40 VTAIL.n39 9.3005
R343 VTAIL.n49 VTAIL.n48 9.3005
R344 VTAIL.n47 VTAIL.n46 9.3005
R345 VTAIL.n97 VTAIL.n96 9.3005
R346 VTAIL.n70 VTAIL.n69 9.3005
R347 VTAIL.n91 VTAIL.n90 9.3005
R348 VTAIL.n89 VTAIL.n88 9.3005
R349 VTAIL.n74 VTAIL.n73 9.3005
R350 VTAIL.n83 VTAIL.n82 9.3005
R351 VTAIL.n81 VTAIL.n80 9.3005
R352 VTAIL.n229 VTAIL.n228 9.3005
R353 VTAIL.n202 VTAIL.n201 9.3005
R354 VTAIL.n223 VTAIL.n222 9.3005
R355 VTAIL.n221 VTAIL.n220 9.3005
R356 VTAIL.n206 VTAIL.n205 9.3005
R357 VTAIL.n215 VTAIL.n214 9.3005
R358 VTAIL.n213 VTAIL.n212 9.3005
R359 VTAIL.n195 VTAIL.n194 9.3005
R360 VTAIL.n168 VTAIL.n167 9.3005
R361 VTAIL.n189 VTAIL.n188 9.3005
R362 VTAIL.n187 VTAIL.n186 9.3005
R363 VTAIL.n172 VTAIL.n171 9.3005
R364 VTAIL.n181 VTAIL.n180 9.3005
R365 VTAIL.n179 VTAIL.n178 9.3005
R366 VTAIL.n163 VTAIL.n162 9.3005
R367 VTAIL.n136 VTAIL.n135 9.3005
R368 VTAIL.n157 VTAIL.n156 9.3005
R369 VTAIL.n155 VTAIL.n154 9.3005
R370 VTAIL.n140 VTAIL.n139 9.3005
R371 VTAIL.n149 VTAIL.n148 9.3005
R372 VTAIL.n147 VTAIL.n146 9.3005
R373 VTAIL.n129 VTAIL.n128 9.3005
R374 VTAIL.n102 VTAIL.n101 9.3005
R375 VTAIL.n123 VTAIL.n122 9.3005
R376 VTAIL.n121 VTAIL.n120 9.3005
R377 VTAIL.n106 VTAIL.n105 9.3005
R378 VTAIL.n115 VTAIL.n114 9.3005
R379 VTAIL.n113 VTAIL.n112 9.3005
R380 VTAIL.n259 VTAIL.n234 8.92171
R381 VTAIL.n29 VTAIL.n4 8.92171
R382 VTAIL.n61 VTAIL.n36 8.92171
R383 VTAIL.n95 VTAIL.n70 8.92171
R384 VTAIL.n227 VTAIL.n202 8.92171
R385 VTAIL.n193 VTAIL.n168 8.92171
R386 VTAIL.n161 VTAIL.n136 8.92171
R387 VTAIL.n127 VTAIL.n102 8.92171
R388 VTAIL.n260 VTAIL.n232 8.14595
R389 VTAIL.n30 VTAIL.n2 8.14595
R390 VTAIL.n62 VTAIL.n34 8.14595
R391 VTAIL.n96 VTAIL.n68 8.14595
R392 VTAIL.n228 VTAIL.n200 8.14595
R393 VTAIL.n194 VTAIL.n166 8.14595
R394 VTAIL.n162 VTAIL.n134 8.14595
R395 VTAIL.n128 VTAIL.n100 8.14595
R396 VTAIL.n262 VTAIL.n232 5.81868
R397 VTAIL.n32 VTAIL.n2 5.81868
R398 VTAIL.n64 VTAIL.n34 5.81868
R399 VTAIL.n98 VTAIL.n68 5.81868
R400 VTAIL.n230 VTAIL.n200 5.81868
R401 VTAIL.n196 VTAIL.n166 5.81868
R402 VTAIL.n164 VTAIL.n134 5.81868
R403 VTAIL.n130 VTAIL.n100 5.81868
R404 VTAIL.n0 VTAIL.t3 5.37323
R405 VTAIL.n0 VTAIL.t5 5.37323
R406 VTAIL.n66 VTAIL.t12 5.37323
R407 VTAIL.n66 VTAIL.t8 5.37323
R408 VTAIL.n198 VTAIL.t14 5.37323
R409 VTAIL.n198 VTAIL.t15 5.37323
R410 VTAIL.n132 VTAIL.t4 5.37323
R411 VTAIL.n132 VTAIL.t6 5.37323
R412 VTAIL.n260 VTAIL.n259 5.04292
R413 VTAIL.n30 VTAIL.n29 5.04292
R414 VTAIL.n62 VTAIL.n61 5.04292
R415 VTAIL.n96 VTAIL.n95 5.04292
R416 VTAIL.n228 VTAIL.n227 5.04292
R417 VTAIL.n194 VTAIL.n193 5.04292
R418 VTAIL.n162 VTAIL.n161 5.04292
R419 VTAIL.n128 VTAIL.n127 5.04292
R420 VTAIL.n256 VTAIL.n234 4.26717
R421 VTAIL.n26 VTAIL.n4 4.26717
R422 VTAIL.n58 VTAIL.n36 4.26717
R423 VTAIL.n92 VTAIL.n70 4.26717
R424 VTAIL.n224 VTAIL.n202 4.26717
R425 VTAIL.n190 VTAIL.n168 4.26717
R426 VTAIL.n158 VTAIL.n136 4.26717
R427 VTAIL.n124 VTAIL.n102 4.26717
R428 VTAIL.n213 VTAIL.n209 3.71286
R429 VTAIL.n179 VTAIL.n175 3.71286
R430 VTAIL.n147 VTAIL.n143 3.71286
R431 VTAIL.n113 VTAIL.n109 3.71286
R432 VTAIL.n245 VTAIL.n241 3.71286
R433 VTAIL.n15 VTAIL.n11 3.71286
R434 VTAIL.n47 VTAIL.n43 3.71286
R435 VTAIL.n81 VTAIL.n77 3.71286
R436 VTAIL.n255 VTAIL.n236 3.49141
R437 VTAIL.n25 VTAIL.n6 3.49141
R438 VTAIL.n57 VTAIL.n38 3.49141
R439 VTAIL.n91 VTAIL.n72 3.49141
R440 VTAIL.n223 VTAIL.n204 3.49141
R441 VTAIL.n189 VTAIL.n170 3.49141
R442 VTAIL.n157 VTAIL.n138 3.49141
R443 VTAIL.n123 VTAIL.n104 3.49141
R444 VTAIL.n133 VTAIL.n131 3.05222
R445 VTAIL.n165 VTAIL.n133 3.05222
R446 VTAIL.n199 VTAIL.n197 3.05222
R447 VTAIL.n231 VTAIL.n199 3.05222
R448 VTAIL.n99 VTAIL.n67 3.05222
R449 VTAIL.n67 VTAIL.n65 3.05222
R450 VTAIL.n33 VTAIL.n1 3.05222
R451 VTAIL VTAIL.n263 2.99403
R452 VTAIL.n252 VTAIL.n251 2.71565
R453 VTAIL.n22 VTAIL.n21 2.71565
R454 VTAIL.n54 VTAIL.n53 2.71565
R455 VTAIL.n88 VTAIL.n87 2.71565
R456 VTAIL.n220 VTAIL.n219 2.71565
R457 VTAIL.n186 VTAIL.n185 2.71565
R458 VTAIL.n154 VTAIL.n153 2.71565
R459 VTAIL.n120 VTAIL.n119 2.71565
R460 VTAIL.n248 VTAIL.n238 1.93989
R461 VTAIL.n18 VTAIL.n8 1.93989
R462 VTAIL.n50 VTAIL.n40 1.93989
R463 VTAIL.n84 VTAIL.n74 1.93989
R464 VTAIL.n216 VTAIL.n206 1.93989
R465 VTAIL.n182 VTAIL.n172 1.93989
R466 VTAIL.n150 VTAIL.n140 1.93989
R467 VTAIL.n116 VTAIL.n106 1.93989
R468 VTAIL.n247 VTAIL.n240 1.16414
R469 VTAIL.n17 VTAIL.n10 1.16414
R470 VTAIL.n49 VTAIL.n42 1.16414
R471 VTAIL.n83 VTAIL.n76 1.16414
R472 VTAIL.n215 VTAIL.n208 1.16414
R473 VTAIL.n181 VTAIL.n174 1.16414
R474 VTAIL.n149 VTAIL.n142 1.16414
R475 VTAIL.n115 VTAIL.n108 1.16414
R476 VTAIL.n197 VTAIL.n165 0.470328
R477 VTAIL.n65 VTAIL.n33 0.470328
R478 VTAIL.n244 VTAIL.n243 0.388379
R479 VTAIL.n14 VTAIL.n13 0.388379
R480 VTAIL.n46 VTAIL.n45 0.388379
R481 VTAIL.n80 VTAIL.n79 0.388379
R482 VTAIL.n212 VTAIL.n211 0.388379
R483 VTAIL.n178 VTAIL.n177 0.388379
R484 VTAIL.n146 VTAIL.n145 0.388379
R485 VTAIL.n112 VTAIL.n111 0.388379
R486 VTAIL.n246 VTAIL.n245 0.155672
R487 VTAIL.n246 VTAIL.n237 0.155672
R488 VTAIL.n253 VTAIL.n237 0.155672
R489 VTAIL.n254 VTAIL.n253 0.155672
R490 VTAIL.n254 VTAIL.n233 0.155672
R491 VTAIL.n261 VTAIL.n233 0.155672
R492 VTAIL.n16 VTAIL.n15 0.155672
R493 VTAIL.n16 VTAIL.n7 0.155672
R494 VTAIL.n23 VTAIL.n7 0.155672
R495 VTAIL.n24 VTAIL.n23 0.155672
R496 VTAIL.n24 VTAIL.n3 0.155672
R497 VTAIL.n31 VTAIL.n3 0.155672
R498 VTAIL.n48 VTAIL.n47 0.155672
R499 VTAIL.n48 VTAIL.n39 0.155672
R500 VTAIL.n55 VTAIL.n39 0.155672
R501 VTAIL.n56 VTAIL.n55 0.155672
R502 VTAIL.n56 VTAIL.n35 0.155672
R503 VTAIL.n63 VTAIL.n35 0.155672
R504 VTAIL.n82 VTAIL.n81 0.155672
R505 VTAIL.n82 VTAIL.n73 0.155672
R506 VTAIL.n89 VTAIL.n73 0.155672
R507 VTAIL.n90 VTAIL.n89 0.155672
R508 VTAIL.n90 VTAIL.n69 0.155672
R509 VTAIL.n97 VTAIL.n69 0.155672
R510 VTAIL.n229 VTAIL.n201 0.155672
R511 VTAIL.n222 VTAIL.n201 0.155672
R512 VTAIL.n222 VTAIL.n221 0.155672
R513 VTAIL.n221 VTAIL.n205 0.155672
R514 VTAIL.n214 VTAIL.n205 0.155672
R515 VTAIL.n214 VTAIL.n213 0.155672
R516 VTAIL.n195 VTAIL.n167 0.155672
R517 VTAIL.n188 VTAIL.n167 0.155672
R518 VTAIL.n188 VTAIL.n187 0.155672
R519 VTAIL.n187 VTAIL.n171 0.155672
R520 VTAIL.n180 VTAIL.n171 0.155672
R521 VTAIL.n180 VTAIL.n179 0.155672
R522 VTAIL.n163 VTAIL.n135 0.155672
R523 VTAIL.n156 VTAIL.n135 0.155672
R524 VTAIL.n156 VTAIL.n155 0.155672
R525 VTAIL.n155 VTAIL.n139 0.155672
R526 VTAIL.n148 VTAIL.n139 0.155672
R527 VTAIL.n148 VTAIL.n147 0.155672
R528 VTAIL.n129 VTAIL.n101 0.155672
R529 VTAIL.n122 VTAIL.n101 0.155672
R530 VTAIL.n122 VTAIL.n121 0.155672
R531 VTAIL.n121 VTAIL.n105 0.155672
R532 VTAIL.n114 VTAIL.n105 0.155672
R533 VTAIL.n114 VTAIL.n113 0.155672
R534 VTAIL VTAIL.n1 0.0586897
R535 VDD1 VDD1.n0 94.848
R536 VDD1.n3 VDD1.n2 94.7343
R537 VDD1.n3 VDD1.n1 94.7343
R538 VDD1.n5 VDD1.n4 93.2638
R539 VDD1.n5 VDD1.n3 43.2466
R540 VDD1.n4 VDD1.t6 5.37323
R541 VDD1.n4 VDD1.t3 5.37323
R542 VDD1.n0 VDD1.t1 5.37323
R543 VDD1.n0 VDD1.t7 5.37323
R544 VDD1.n2 VDD1.t4 5.37323
R545 VDD1.n2 VDD1.t2 5.37323
R546 VDD1.n1 VDD1.t0 5.37323
R547 VDD1.n1 VDD1.t5 5.37323
R548 VDD1 VDD1.n5 1.46817
R549 B.n548 B.n65 585
R550 B.n550 B.n549 585
R551 B.n551 B.n64 585
R552 B.n553 B.n552 585
R553 B.n554 B.n63 585
R554 B.n556 B.n555 585
R555 B.n557 B.n62 585
R556 B.n559 B.n558 585
R557 B.n560 B.n61 585
R558 B.n562 B.n561 585
R559 B.n563 B.n60 585
R560 B.n565 B.n564 585
R561 B.n566 B.n59 585
R562 B.n568 B.n567 585
R563 B.n569 B.n58 585
R564 B.n571 B.n570 585
R565 B.n572 B.n57 585
R566 B.n574 B.n573 585
R567 B.n575 B.n56 585
R568 B.n577 B.n576 585
R569 B.n578 B.n55 585
R570 B.n580 B.n579 585
R571 B.n581 B.n54 585
R572 B.n583 B.n582 585
R573 B.n585 B.n51 585
R574 B.n587 B.n586 585
R575 B.n588 B.n50 585
R576 B.n590 B.n589 585
R577 B.n591 B.n49 585
R578 B.n593 B.n592 585
R579 B.n594 B.n48 585
R580 B.n596 B.n595 585
R581 B.n597 B.n47 585
R582 B.n599 B.n598 585
R583 B.n601 B.n600 585
R584 B.n602 B.n43 585
R585 B.n604 B.n603 585
R586 B.n605 B.n42 585
R587 B.n607 B.n606 585
R588 B.n608 B.n41 585
R589 B.n610 B.n609 585
R590 B.n611 B.n40 585
R591 B.n613 B.n612 585
R592 B.n614 B.n39 585
R593 B.n616 B.n615 585
R594 B.n617 B.n38 585
R595 B.n619 B.n618 585
R596 B.n620 B.n37 585
R597 B.n622 B.n621 585
R598 B.n623 B.n36 585
R599 B.n625 B.n624 585
R600 B.n626 B.n35 585
R601 B.n628 B.n627 585
R602 B.n629 B.n34 585
R603 B.n631 B.n630 585
R604 B.n632 B.n33 585
R605 B.n634 B.n633 585
R606 B.n635 B.n32 585
R607 B.n547 B.n546 585
R608 B.n545 B.n66 585
R609 B.n544 B.n543 585
R610 B.n542 B.n67 585
R611 B.n541 B.n540 585
R612 B.n539 B.n68 585
R613 B.n538 B.n537 585
R614 B.n536 B.n69 585
R615 B.n535 B.n534 585
R616 B.n533 B.n70 585
R617 B.n532 B.n531 585
R618 B.n530 B.n71 585
R619 B.n529 B.n528 585
R620 B.n527 B.n72 585
R621 B.n526 B.n525 585
R622 B.n524 B.n73 585
R623 B.n523 B.n522 585
R624 B.n521 B.n74 585
R625 B.n520 B.n519 585
R626 B.n518 B.n75 585
R627 B.n517 B.n516 585
R628 B.n515 B.n76 585
R629 B.n514 B.n513 585
R630 B.n512 B.n77 585
R631 B.n511 B.n510 585
R632 B.n509 B.n78 585
R633 B.n508 B.n507 585
R634 B.n506 B.n79 585
R635 B.n505 B.n504 585
R636 B.n503 B.n80 585
R637 B.n502 B.n501 585
R638 B.n500 B.n81 585
R639 B.n499 B.n498 585
R640 B.n497 B.n82 585
R641 B.n496 B.n495 585
R642 B.n494 B.n83 585
R643 B.n493 B.n492 585
R644 B.n491 B.n84 585
R645 B.n490 B.n489 585
R646 B.n488 B.n85 585
R647 B.n487 B.n486 585
R648 B.n485 B.n86 585
R649 B.n484 B.n483 585
R650 B.n482 B.n87 585
R651 B.n481 B.n480 585
R652 B.n479 B.n88 585
R653 B.n478 B.n477 585
R654 B.n476 B.n89 585
R655 B.n475 B.n474 585
R656 B.n473 B.n90 585
R657 B.n472 B.n471 585
R658 B.n470 B.n91 585
R659 B.n469 B.n468 585
R660 B.n467 B.n92 585
R661 B.n466 B.n465 585
R662 B.n464 B.n93 585
R663 B.n463 B.n462 585
R664 B.n461 B.n94 585
R665 B.n460 B.n459 585
R666 B.n458 B.n95 585
R667 B.n457 B.n456 585
R668 B.n455 B.n96 585
R669 B.n454 B.n453 585
R670 B.n452 B.n97 585
R671 B.n451 B.n450 585
R672 B.n449 B.n98 585
R673 B.n448 B.n447 585
R674 B.n446 B.n99 585
R675 B.n445 B.n444 585
R676 B.n443 B.n100 585
R677 B.n442 B.n441 585
R678 B.n440 B.n101 585
R679 B.n439 B.n438 585
R680 B.n437 B.n102 585
R681 B.n436 B.n435 585
R682 B.n434 B.n103 585
R683 B.n433 B.n432 585
R684 B.n431 B.n104 585
R685 B.n430 B.n429 585
R686 B.n428 B.n105 585
R687 B.n427 B.n426 585
R688 B.n425 B.n106 585
R689 B.n424 B.n423 585
R690 B.n422 B.n107 585
R691 B.n421 B.n420 585
R692 B.n419 B.n108 585
R693 B.n418 B.n417 585
R694 B.n416 B.n109 585
R695 B.n415 B.n414 585
R696 B.n413 B.n110 585
R697 B.n412 B.n411 585
R698 B.n410 B.n111 585
R699 B.n409 B.n408 585
R700 B.n407 B.n112 585
R701 B.n406 B.n405 585
R702 B.n404 B.n113 585
R703 B.n403 B.n402 585
R704 B.n401 B.n114 585
R705 B.n400 B.n399 585
R706 B.n398 B.n115 585
R707 B.n397 B.n396 585
R708 B.n395 B.n116 585
R709 B.n394 B.n393 585
R710 B.n392 B.n117 585
R711 B.n391 B.n390 585
R712 B.n389 B.n118 585
R713 B.n388 B.n387 585
R714 B.n386 B.n119 585
R715 B.n385 B.n384 585
R716 B.n383 B.n120 585
R717 B.n382 B.n381 585
R718 B.n380 B.n121 585
R719 B.n379 B.n378 585
R720 B.n377 B.n122 585
R721 B.n376 B.n375 585
R722 B.n374 B.n123 585
R723 B.n373 B.n372 585
R724 B.n371 B.n124 585
R725 B.n370 B.n369 585
R726 B.n368 B.n125 585
R727 B.n367 B.n366 585
R728 B.n278 B.n159 585
R729 B.n280 B.n279 585
R730 B.n281 B.n158 585
R731 B.n283 B.n282 585
R732 B.n284 B.n157 585
R733 B.n286 B.n285 585
R734 B.n287 B.n156 585
R735 B.n289 B.n288 585
R736 B.n290 B.n155 585
R737 B.n292 B.n291 585
R738 B.n293 B.n154 585
R739 B.n295 B.n294 585
R740 B.n296 B.n153 585
R741 B.n298 B.n297 585
R742 B.n299 B.n152 585
R743 B.n301 B.n300 585
R744 B.n302 B.n151 585
R745 B.n304 B.n303 585
R746 B.n305 B.n150 585
R747 B.n307 B.n306 585
R748 B.n308 B.n149 585
R749 B.n310 B.n309 585
R750 B.n311 B.n148 585
R751 B.n313 B.n312 585
R752 B.n315 B.n145 585
R753 B.n317 B.n316 585
R754 B.n318 B.n144 585
R755 B.n320 B.n319 585
R756 B.n321 B.n143 585
R757 B.n323 B.n322 585
R758 B.n324 B.n142 585
R759 B.n326 B.n325 585
R760 B.n327 B.n141 585
R761 B.n329 B.n328 585
R762 B.n331 B.n330 585
R763 B.n332 B.n137 585
R764 B.n334 B.n333 585
R765 B.n335 B.n136 585
R766 B.n337 B.n336 585
R767 B.n338 B.n135 585
R768 B.n340 B.n339 585
R769 B.n341 B.n134 585
R770 B.n343 B.n342 585
R771 B.n344 B.n133 585
R772 B.n346 B.n345 585
R773 B.n347 B.n132 585
R774 B.n349 B.n348 585
R775 B.n350 B.n131 585
R776 B.n352 B.n351 585
R777 B.n353 B.n130 585
R778 B.n355 B.n354 585
R779 B.n356 B.n129 585
R780 B.n358 B.n357 585
R781 B.n359 B.n128 585
R782 B.n361 B.n360 585
R783 B.n362 B.n127 585
R784 B.n364 B.n363 585
R785 B.n365 B.n126 585
R786 B.n277 B.n276 585
R787 B.n275 B.n160 585
R788 B.n274 B.n273 585
R789 B.n272 B.n161 585
R790 B.n271 B.n270 585
R791 B.n269 B.n162 585
R792 B.n268 B.n267 585
R793 B.n266 B.n163 585
R794 B.n265 B.n264 585
R795 B.n263 B.n164 585
R796 B.n262 B.n261 585
R797 B.n260 B.n165 585
R798 B.n259 B.n258 585
R799 B.n257 B.n166 585
R800 B.n256 B.n255 585
R801 B.n254 B.n167 585
R802 B.n253 B.n252 585
R803 B.n251 B.n168 585
R804 B.n250 B.n249 585
R805 B.n248 B.n169 585
R806 B.n247 B.n246 585
R807 B.n245 B.n170 585
R808 B.n244 B.n243 585
R809 B.n242 B.n171 585
R810 B.n241 B.n240 585
R811 B.n239 B.n172 585
R812 B.n238 B.n237 585
R813 B.n236 B.n173 585
R814 B.n235 B.n234 585
R815 B.n233 B.n174 585
R816 B.n232 B.n231 585
R817 B.n230 B.n175 585
R818 B.n229 B.n228 585
R819 B.n227 B.n176 585
R820 B.n226 B.n225 585
R821 B.n224 B.n177 585
R822 B.n223 B.n222 585
R823 B.n221 B.n178 585
R824 B.n220 B.n219 585
R825 B.n218 B.n179 585
R826 B.n217 B.n216 585
R827 B.n215 B.n180 585
R828 B.n214 B.n213 585
R829 B.n212 B.n181 585
R830 B.n211 B.n210 585
R831 B.n209 B.n182 585
R832 B.n208 B.n207 585
R833 B.n206 B.n183 585
R834 B.n205 B.n204 585
R835 B.n203 B.n184 585
R836 B.n202 B.n201 585
R837 B.n200 B.n185 585
R838 B.n199 B.n198 585
R839 B.n197 B.n186 585
R840 B.n196 B.n195 585
R841 B.n194 B.n187 585
R842 B.n193 B.n192 585
R843 B.n191 B.n188 585
R844 B.n190 B.n189 585
R845 B.n2 B.n0 585
R846 B.n725 B.n1 585
R847 B.n724 B.n723 585
R848 B.n722 B.n3 585
R849 B.n721 B.n720 585
R850 B.n719 B.n4 585
R851 B.n718 B.n717 585
R852 B.n716 B.n5 585
R853 B.n715 B.n714 585
R854 B.n713 B.n6 585
R855 B.n712 B.n711 585
R856 B.n710 B.n7 585
R857 B.n709 B.n708 585
R858 B.n707 B.n8 585
R859 B.n706 B.n705 585
R860 B.n704 B.n9 585
R861 B.n703 B.n702 585
R862 B.n701 B.n10 585
R863 B.n700 B.n699 585
R864 B.n698 B.n11 585
R865 B.n697 B.n696 585
R866 B.n695 B.n12 585
R867 B.n694 B.n693 585
R868 B.n692 B.n13 585
R869 B.n691 B.n690 585
R870 B.n689 B.n14 585
R871 B.n688 B.n687 585
R872 B.n686 B.n15 585
R873 B.n685 B.n684 585
R874 B.n683 B.n16 585
R875 B.n682 B.n681 585
R876 B.n680 B.n17 585
R877 B.n679 B.n678 585
R878 B.n677 B.n18 585
R879 B.n676 B.n675 585
R880 B.n674 B.n19 585
R881 B.n673 B.n672 585
R882 B.n671 B.n20 585
R883 B.n670 B.n669 585
R884 B.n668 B.n21 585
R885 B.n667 B.n666 585
R886 B.n665 B.n22 585
R887 B.n664 B.n663 585
R888 B.n662 B.n23 585
R889 B.n661 B.n660 585
R890 B.n659 B.n24 585
R891 B.n658 B.n657 585
R892 B.n656 B.n25 585
R893 B.n655 B.n654 585
R894 B.n653 B.n26 585
R895 B.n652 B.n651 585
R896 B.n650 B.n27 585
R897 B.n649 B.n648 585
R898 B.n647 B.n28 585
R899 B.n646 B.n645 585
R900 B.n644 B.n29 585
R901 B.n643 B.n642 585
R902 B.n641 B.n30 585
R903 B.n640 B.n639 585
R904 B.n638 B.n31 585
R905 B.n637 B.n636 585
R906 B.n727 B.n726 585
R907 B.n276 B.n159 511.721
R908 B.n636 B.n635 511.721
R909 B.n366 B.n365 511.721
R910 B.n546 B.n65 511.721
R911 B.n138 B.t5 337.817
R912 B.n52 B.t10 337.817
R913 B.n146 B.t2 337.817
R914 B.n44 B.t7 337.817
R915 B.n139 B.t4 269.163
R916 B.n53 B.t11 269.163
R917 B.n147 B.t1 269.163
R918 B.n45 B.t8 269.163
R919 B.n138 B.t3 254.236
R920 B.n146 B.t0 254.236
R921 B.n44 B.t6 254.236
R922 B.n52 B.t9 254.236
R923 B.n276 B.n275 163.367
R924 B.n275 B.n274 163.367
R925 B.n274 B.n161 163.367
R926 B.n270 B.n161 163.367
R927 B.n270 B.n269 163.367
R928 B.n269 B.n268 163.367
R929 B.n268 B.n163 163.367
R930 B.n264 B.n163 163.367
R931 B.n264 B.n263 163.367
R932 B.n263 B.n262 163.367
R933 B.n262 B.n165 163.367
R934 B.n258 B.n165 163.367
R935 B.n258 B.n257 163.367
R936 B.n257 B.n256 163.367
R937 B.n256 B.n167 163.367
R938 B.n252 B.n167 163.367
R939 B.n252 B.n251 163.367
R940 B.n251 B.n250 163.367
R941 B.n250 B.n169 163.367
R942 B.n246 B.n169 163.367
R943 B.n246 B.n245 163.367
R944 B.n245 B.n244 163.367
R945 B.n244 B.n171 163.367
R946 B.n240 B.n171 163.367
R947 B.n240 B.n239 163.367
R948 B.n239 B.n238 163.367
R949 B.n238 B.n173 163.367
R950 B.n234 B.n173 163.367
R951 B.n234 B.n233 163.367
R952 B.n233 B.n232 163.367
R953 B.n232 B.n175 163.367
R954 B.n228 B.n175 163.367
R955 B.n228 B.n227 163.367
R956 B.n227 B.n226 163.367
R957 B.n226 B.n177 163.367
R958 B.n222 B.n177 163.367
R959 B.n222 B.n221 163.367
R960 B.n221 B.n220 163.367
R961 B.n220 B.n179 163.367
R962 B.n216 B.n179 163.367
R963 B.n216 B.n215 163.367
R964 B.n215 B.n214 163.367
R965 B.n214 B.n181 163.367
R966 B.n210 B.n181 163.367
R967 B.n210 B.n209 163.367
R968 B.n209 B.n208 163.367
R969 B.n208 B.n183 163.367
R970 B.n204 B.n183 163.367
R971 B.n204 B.n203 163.367
R972 B.n203 B.n202 163.367
R973 B.n202 B.n185 163.367
R974 B.n198 B.n185 163.367
R975 B.n198 B.n197 163.367
R976 B.n197 B.n196 163.367
R977 B.n196 B.n187 163.367
R978 B.n192 B.n187 163.367
R979 B.n192 B.n191 163.367
R980 B.n191 B.n190 163.367
R981 B.n190 B.n2 163.367
R982 B.n726 B.n2 163.367
R983 B.n726 B.n725 163.367
R984 B.n725 B.n724 163.367
R985 B.n724 B.n3 163.367
R986 B.n720 B.n3 163.367
R987 B.n720 B.n719 163.367
R988 B.n719 B.n718 163.367
R989 B.n718 B.n5 163.367
R990 B.n714 B.n5 163.367
R991 B.n714 B.n713 163.367
R992 B.n713 B.n712 163.367
R993 B.n712 B.n7 163.367
R994 B.n708 B.n7 163.367
R995 B.n708 B.n707 163.367
R996 B.n707 B.n706 163.367
R997 B.n706 B.n9 163.367
R998 B.n702 B.n9 163.367
R999 B.n702 B.n701 163.367
R1000 B.n701 B.n700 163.367
R1001 B.n700 B.n11 163.367
R1002 B.n696 B.n11 163.367
R1003 B.n696 B.n695 163.367
R1004 B.n695 B.n694 163.367
R1005 B.n694 B.n13 163.367
R1006 B.n690 B.n13 163.367
R1007 B.n690 B.n689 163.367
R1008 B.n689 B.n688 163.367
R1009 B.n688 B.n15 163.367
R1010 B.n684 B.n15 163.367
R1011 B.n684 B.n683 163.367
R1012 B.n683 B.n682 163.367
R1013 B.n682 B.n17 163.367
R1014 B.n678 B.n17 163.367
R1015 B.n678 B.n677 163.367
R1016 B.n677 B.n676 163.367
R1017 B.n676 B.n19 163.367
R1018 B.n672 B.n19 163.367
R1019 B.n672 B.n671 163.367
R1020 B.n671 B.n670 163.367
R1021 B.n670 B.n21 163.367
R1022 B.n666 B.n21 163.367
R1023 B.n666 B.n665 163.367
R1024 B.n665 B.n664 163.367
R1025 B.n664 B.n23 163.367
R1026 B.n660 B.n23 163.367
R1027 B.n660 B.n659 163.367
R1028 B.n659 B.n658 163.367
R1029 B.n658 B.n25 163.367
R1030 B.n654 B.n25 163.367
R1031 B.n654 B.n653 163.367
R1032 B.n653 B.n652 163.367
R1033 B.n652 B.n27 163.367
R1034 B.n648 B.n27 163.367
R1035 B.n648 B.n647 163.367
R1036 B.n647 B.n646 163.367
R1037 B.n646 B.n29 163.367
R1038 B.n642 B.n29 163.367
R1039 B.n642 B.n641 163.367
R1040 B.n641 B.n640 163.367
R1041 B.n640 B.n31 163.367
R1042 B.n636 B.n31 163.367
R1043 B.n280 B.n159 163.367
R1044 B.n281 B.n280 163.367
R1045 B.n282 B.n281 163.367
R1046 B.n282 B.n157 163.367
R1047 B.n286 B.n157 163.367
R1048 B.n287 B.n286 163.367
R1049 B.n288 B.n287 163.367
R1050 B.n288 B.n155 163.367
R1051 B.n292 B.n155 163.367
R1052 B.n293 B.n292 163.367
R1053 B.n294 B.n293 163.367
R1054 B.n294 B.n153 163.367
R1055 B.n298 B.n153 163.367
R1056 B.n299 B.n298 163.367
R1057 B.n300 B.n299 163.367
R1058 B.n300 B.n151 163.367
R1059 B.n304 B.n151 163.367
R1060 B.n305 B.n304 163.367
R1061 B.n306 B.n305 163.367
R1062 B.n306 B.n149 163.367
R1063 B.n310 B.n149 163.367
R1064 B.n311 B.n310 163.367
R1065 B.n312 B.n311 163.367
R1066 B.n312 B.n145 163.367
R1067 B.n317 B.n145 163.367
R1068 B.n318 B.n317 163.367
R1069 B.n319 B.n318 163.367
R1070 B.n319 B.n143 163.367
R1071 B.n323 B.n143 163.367
R1072 B.n324 B.n323 163.367
R1073 B.n325 B.n324 163.367
R1074 B.n325 B.n141 163.367
R1075 B.n329 B.n141 163.367
R1076 B.n330 B.n329 163.367
R1077 B.n330 B.n137 163.367
R1078 B.n334 B.n137 163.367
R1079 B.n335 B.n334 163.367
R1080 B.n336 B.n335 163.367
R1081 B.n336 B.n135 163.367
R1082 B.n340 B.n135 163.367
R1083 B.n341 B.n340 163.367
R1084 B.n342 B.n341 163.367
R1085 B.n342 B.n133 163.367
R1086 B.n346 B.n133 163.367
R1087 B.n347 B.n346 163.367
R1088 B.n348 B.n347 163.367
R1089 B.n348 B.n131 163.367
R1090 B.n352 B.n131 163.367
R1091 B.n353 B.n352 163.367
R1092 B.n354 B.n353 163.367
R1093 B.n354 B.n129 163.367
R1094 B.n358 B.n129 163.367
R1095 B.n359 B.n358 163.367
R1096 B.n360 B.n359 163.367
R1097 B.n360 B.n127 163.367
R1098 B.n364 B.n127 163.367
R1099 B.n365 B.n364 163.367
R1100 B.n366 B.n125 163.367
R1101 B.n370 B.n125 163.367
R1102 B.n371 B.n370 163.367
R1103 B.n372 B.n371 163.367
R1104 B.n372 B.n123 163.367
R1105 B.n376 B.n123 163.367
R1106 B.n377 B.n376 163.367
R1107 B.n378 B.n377 163.367
R1108 B.n378 B.n121 163.367
R1109 B.n382 B.n121 163.367
R1110 B.n383 B.n382 163.367
R1111 B.n384 B.n383 163.367
R1112 B.n384 B.n119 163.367
R1113 B.n388 B.n119 163.367
R1114 B.n389 B.n388 163.367
R1115 B.n390 B.n389 163.367
R1116 B.n390 B.n117 163.367
R1117 B.n394 B.n117 163.367
R1118 B.n395 B.n394 163.367
R1119 B.n396 B.n395 163.367
R1120 B.n396 B.n115 163.367
R1121 B.n400 B.n115 163.367
R1122 B.n401 B.n400 163.367
R1123 B.n402 B.n401 163.367
R1124 B.n402 B.n113 163.367
R1125 B.n406 B.n113 163.367
R1126 B.n407 B.n406 163.367
R1127 B.n408 B.n407 163.367
R1128 B.n408 B.n111 163.367
R1129 B.n412 B.n111 163.367
R1130 B.n413 B.n412 163.367
R1131 B.n414 B.n413 163.367
R1132 B.n414 B.n109 163.367
R1133 B.n418 B.n109 163.367
R1134 B.n419 B.n418 163.367
R1135 B.n420 B.n419 163.367
R1136 B.n420 B.n107 163.367
R1137 B.n424 B.n107 163.367
R1138 B.n425 B.n424 163.367
R1139 B.n426 B.n425 163.367
R1140 B.n426 B.n105 163.367
R1141 B.n430 B.n105 163.367
R1142 B.n431 B.n430 163.367
R1143 B.n432 B.n431 163.367
R1144 B.n432 B.n103 163.367
R1145 B.n436 B.n103 163.367
R1146 B.n437 B.n436 163.367
R1147 B.n438 B.n437 163.367
R1148 B.n438 B.n101 163.367
R1149 B.n442 B.n101 163.367
R1150 B.n443 B.n442 163.367
R1151 B.n444 B.n443 163.367
R1152 B.n444 B.n99 163.367
R1153 B.n448 B.n99 163.367
R1154 B.n449 B.n448 163.367
R1155 B.n450 B.n449 163.367
R1156 B.n450 B.n97 163.367
R1157 B.n454 B.n97 163.367
R1158 B.n455 B.n454 163.367
R1159 B.n456 B.n455 163.367
R1160 B.n456 B.n95 163.367
R1161 B.n460 B.n95 163.367
R1162 B.n461 B.n460 163.367
R1163 B.n462 B.n461 163.367
R1164 B.n462 B.n93 163.367
R1165 B.n466 B.n93 163.367
R1166 B.n467 B.n466 163.367
R1167 B.n468 B.n467 163.367
R1168 B.n468 B.n91 163.367
R1169 B.n472 B.n91 163.367
R1170 B.n473 B.n472 163.367
R1171 B.n474 B.n473 163.367
R1172 B.n474 B.n89 163.367
R1173 B.n478 B.n89 163.367
R1174 B.n479 B.n478 163.367
R1175 B.n480 B.n479 163.367
R1176 B.n480 B.n87 163.367
R1177 B.n484 B.n87 163.367
R1178 B.n485 B.n484 163.367
R1179 B.n486 B.n485 163.367
R1180 B.n486 B.n85 163.367
R1181 B.n490 B.n85 163.367
R1182 B.n491 B.n490 163.367
R1183 B.n492 B.n491 163.367
R1184 B.n492 B.n83 163.367
R1185 B.n496 B.n83 163.367
R1186 B.n497 B.n496 163.367
R1187 B.n498 B.n497 163.367
R1188 B.n498 B.n81 163.367
R1189 B.n502 B.n81 163.367
R1190 B.n503 B.n502 163.367
R1191 B.n504 B.n503 163.367
R1192 B.n504 B.n79 163.367
R1193 B.n508 B.n79 163.367
R1194 B.n509 B.n508 163.367
R1195 B.n510 B.n509 163.367
R1196 B.n510 B.n77 163.367
R1197 B.n514 B.n77 163.367
R1198 B.n515 B.n514 163.367
R1199 B.n516 B.n515 163.367
R1200 B.n516 B.n75 163.367
R1201 B.n520 B.n75 163.367
R1202 B.n521 B.n520 163.367
R1203 B.n522 B.n521 163.367
R1204 B.n522 B.n73 163.367
R1205 B.n526 B.n73 163.367
R1206 B.n527 B.n526 163.367
R1207 B.n528 B.n527 163.367
R1208 B.n528 B.n71 163.367
R1209 B.n532 B.n71 163.367
R1210 B.n533 B.n532 163.367
R1211 B.n534 B.n533 163.367
R1212 B.n534 B.n69 163.367
R1213 B.n538 B.n69 163.367
R1214 B.n539 B.n538 163.367
R1215 B.n540 B.n539 163.367
R1216 B.n540 B.n67 163.367
R1217 B.n544 B.n67 163.367
R1218 B.n545 B.n544 163.367
R1219 B.n546 B.n545 163.367
R1220 B.n635 B.n634 163.367
R1221 B.n634 B.n33 163.367
R1222 B.n630 B.n33 163.367
R1223 B.n630 B.n629 163.367
R1224 B.n629 B.n628 163.367
R1225 B.n628 B.n35 163.367
R1226 B.n624 B.n35 163.367
R1227 B.n624 B.n623 163.367
R1228 B.n623 B.n622 163.367
R1229 B.n622 B.n37 163.367
R1230 B.n618 B.n37 163.367
R1231 B.n618 B.n617 163.367
R1232 B.n617 B.n616 163.367
R1233 B.n616 B.n39 163.367
R1234 B.n612 B.n39 163.367
R1235 B.n612 B.n611 163.367
R1236 B.n611 B.n610 163.367
R1237 B.n610 B.n41 163.367
R1238 B.n606 B.n41 163.367
R1239 B.n606 B.n605 163.367
R1240 B.n605 B.n604 163.367
R1241 B.n604 B.n43 163.367
R1242 B.n600 B.n43 163.367
R1243 B.n600 B.n599 163.367
R1244 B.n599 B.n47 163.367
R1245 B.n595 B.n47 163.367
R1246 B.n595 B.n594 163.367
R1247 B.n594 B.n593 163.367
R1248 B.n593 B.n49 163.367
R1249 B.n589 B.n49 163.367
R1250 B.n589 B.n588 163.367
R1251 B.n588 B.n587 163.367
R1252 B.n587 B.n51 163.367
R1253 B.n582 B.n51 163.367
R1254 B.n582 B.n581 163.367
R1255 B.n581 B.n580 163.367
R1256 B.n580 B.n55 163.367
R1257 B.n576 B.n55 163.367
R1258 B.n576 B.n575 163.367
R1259 B.n575 B.n574 163.367
R1260 B.n574 B.n57 163.367
R1261 B.n570 B.n57 163.367
R1262 B.n570 B.n569 163.367
R1263 B.n569 B.n568 163.367
R1264 B.n568 B.n59 163.367
R1265 B.n564 B.n59 163.367
R1266 B.n564 B.n563 163.367
R1267 B.n563 B.n562 163.367
R1268 B.n562 B.n61 163.367
R1269 B.n558 B.n61 163.367
R1270 B.n558 B.n557 163.367
R1271 B.n557 B.n556 163.367
R1272 B.n556 B.n63 163.367
R1273 B.n552 B.n63 163.367
R1274 B.n552 B.n551 163.367
R1275 B.n551 B.n550 163.367
R1276 B.n550 B.n65 163.367
R1277 B.n139 B.n138 68.655
R1278 B.n147 B.n146 68.655
R1279 B.n45 B.n44 68.655
R1280 B.n53 B.n52 68.655
R1281 B.n140 B.n139 59.5399
R1282 B.n314 B.n147 59.5399
R1283 B.n46 B.n45 59.5399
R1284 B.n584 B.n53 59.5399
R1285 B.n637 B.n32 33.2493
R1286 B.n548 B.n547 33.2493
R1287 B.n367 B.n126 33.2493
R1288 B.n278 B.n277 33.2493
R1289 B B.n727 18.0485
R1290 B.n633 B.n32 10.6151
R1291 B.n633 B.n632 10.6151
R1292 B.n632 B.n631 10.6151
R1293 B.n631 B.n34 10.6151
R1294 B.n627 B.n34 10.6151
R1295 B.n627 B.n626 10.6151
R1296 B.n626 B.n625 10.6151
R1297 B.n625 B.n36 10.6151
R1298 B.n621 B.n36 10.6151
R1299 B.n621 B.n620 10.6151
R1300 B.n620 B.n619 10.6151
R1301 B.n619 B.n38 10.6151
R1302 B.n615 B.n38 10.6151
R1303 B.n615 B.n614 10.6151
R1304 B.n614 B.n613 10.6151
R1305 B.n613 B.n40 10.6151
R1306 B.n609 B.n40 10.6151
R1307 B.n609 B.n608 10.6151
R1308 B.n608 B.n607 10.6151
R1309 B.n607 B.n42 10.6151
R1310 B.n603 B.n42 10.6151
R1311 B.n603 B.n602 10.6151
R1312 B.n602 B.n601 10.6151
R1313 B.n598 B.n597 10.6151
R1314 B.n597 B.n596 10.6151
R1315 B.n596 B.n48 10.6151
R1316 B.n592 B.n48 10.6151
R1317 B.n592 B.n591 10.6151
R1318 B.n591 B.n590 10.6151
R1319 B.n590 B.n50 10.6151
R1320 B.n586 B.n50 10.6151
R1321 B.n586 B.n585 10.6151
R1322 B.n583 B.n54 10.6151
R1323 B.n579 B.n54 10.6151
R1324 B.n579 B.n578 10.6151
R1325 B.n578 B.n577 10.6151
R1326 B.n577 B.n56 10.6151
R1327 B.n573 B.n56 10.6151
R1328 B.n573 B.n572 10.6151
R1329 B.n572 B.n571 10.6151
R1330 B.n571 B.n58 10.6151
R1331 B.n567 B.n58 10.6151
R1332 B.n567 B.n566 10.6151
R1333 B.n566 B.n565 10.6151
R1334 B.n565 B.n60 10.6151
R1335 B.n561 B.n60 10.6151
R1336 B.n561 B.n560 10.6151
R1337 B.n560 B.n559 10.6151
R1338 B.n559 B.n62 10.6151
R1339 B.n555 B.n62 10.6151
R1340 B.n555 B.n554 10.6151
R1341 B.n554 B.n553 10.6151
R1342 B.n553 B.n64 10.6151
R1343 B.n549 B.n64 10.6151
R1344 B.n549 B.n548 10.6151
R1345 B.n368 B.n367 10.6151
R1346 B.n369 B.n368 10.6151
R1347 B.n369 B.n124 10.6151
R1348 B.n373 B.n124 10.6151
R1349 B.n374 B.n373 10.6151
R1350 B.n375 B.n374 10.6151
R1351 B.n375 B.n122 10.6151
R1352 B.n379 B.n122 10.6151
R1353 B.n380 B.n379 10.6151
R1354 B.n381 B.n380 10.6151
R1355 B.n381 B.n120 10.6151
R1356 B.n385 B.n120 10.6151
R1357 B.n386 B.n385 10.6151
R1358 B.n387 B.n386 10.6151
R1359 B.n387 B.n118 10.6151
R1360 B.n391 B.n118 10.6151
R1361 B.n392 B.n391 10.6151
R1362 B.n393 B.n392 10.6151
R1363 B.n393 B.n116 10.6151
R1364 B.n397 B.n116 10.6151
R1365 B.n398 B.n397 10.6151
R1366 B.n399 B.n398 10.6151
R1367 B.n399 B.n114 10.6151
R1368 B.n403 B.n114 10.6151
R1369 B.n404 B.n403 10.6151
R1370 B.n405 B.n404 10.6151
R1371 B.n405 B.n112 10.6151
R1372 B.n409 B.n112 10.6151
R1373 B.n410 B.n409 10.6151
R1374 B.n411 B.n410 10.6151
R1375 B.n411 B.n110 10.6151
R1376 B.n415 B.n110 10.6151
R1377 B.n416 B.n415 10.6151
R1378 B.n417 B.n416 10.6151
R1379 B.n417 B.n108 10.6151
R1380 B.n421 B.n108 10.6151
R1381 B.n422 B.n421 10.6151
R1382 B.n423 B.n422 10.6151
R1383 B.n423 B.n106 10.6151
R1384 B.n427 B.n106 10.6151
R1385 B.n428 B.n427 10.6151
R1386 B.n429 B.n428 10.6151
R1387 B.n429 B.n104 10.6151
R1388 B.n433 B.n104 10.6151
R1389 B.n434 B.n433 10.6151
R1390 B.n435 B.n434 10.6151
R1391 B.n435 B.n102 10.6151
R1392 B.n439 B.n102 10.6151
R1393 B.n440 B.n439 10.6151
R1394 B.n441 B.n440 10.6151
R1395 B.n441 B.n100 10.6151
R1396 B.n445 B.n100 10.6151
R1397 B.n446 B.n445 10.6151
R1398 B.n447 B.n446 10.6151
R1399 B.n447 B.n98 10.6151
R1400 B.n451 B.n98 10.6151
R1401 B.n452 B.n451 10.6151
R1402 B.n453 B.n452 10.6151
R1403 B.n453 B.n96 10.6151
R1404 B.n457 B.n96 10.6151
R1405 B.n458 B.n457 10.6151
R1406 B.n459 B.n458 10.6151
R1407 B.n459 B.n94 10.6151
R1408 B.n463 B.n94 10.6151
R1409 B.n464 B.n463 10.6151
R1410 B.n465 B.n464 10.6151
R1411 B.n465 B.n92 10.6151
R1412 B.n469 B.n92 10.6151
R1413 B.n470 B.n469 10.6151
R1414 B.n471 B.n470 10.6151
R1415 B.n471 B.n90 10.6151
R1416 B.n475 B.n90 10.6151
R1417 B.n476 B.n475 10.6151
R1418 B.n477 B.n476 10.6151
R1419 B.n477 B.n88 10.6151
R1420 B.n481 B.n88 10.6151
R1421 B.n482 B.n481 10.6151
R1422 B.n483 B.n482 10.6151
R1423 B.n483 B.n86 10.6151
R1424 B.n487 B.n86 10.6151
R1425 B.n488 B.n487 10.6151
R1426 B.n489 B.n488 10.6151
R1427 B.n489 B.n84 10.6151
R1428 B.n493 B.n84 10.6151
R1429 B.n494 B.n493 10.6151
R1430 B.n495 B.n494 10.6151
R1431 B.n495 B.n82 10.6151
R1432 B.n499 B.n82 10.6151
R1433 B.n500 B.n499 10.6151
R1434 B.n501 B.n500 10.6151
R1435 B.n501 B.n80 10.6151
R1436 B.n505 B.n80 10.6151
R1437 B.n506 B.n505 10.6151
R1438 B.n507 B.n506 10.6151
R1439 B.n507 B.n78 10.6151
R1440 B.n511 B.n78 10.6151
R1441 B.n512 B.n511 10.6151
R1442 B.n513 B.n512 10.6151
R1443 B.n513 B.n76 10.6151
R1444 B.n517 B.n76 10.6151
R1445 B.n518 B.n517 10.6151
R1446 B.n519 B.n518 10.6151
R1447 B.n519 B.n74 10.6151
R1448 B.n523 B.n74 10.6151
R1449 B.n524 B.n523 10.6151
R1450 B.n525 B.n524 10.6151
R1451 B.n525 B.n72 10.6151
R1452 B.n529 B.n72 10.6151
R1453 B.n530 B.n529 10.6151
R1454 B.n531 B.n530 10.6151
R1455 B.n531 B.n70 10.6151
R1456 B.n535 B.n70 10.6151
R1457 B.n536 B.n535 10.6151
R1458 B.n537 B.n536 10.6151
R1459 B.n537 B.n68 10.6151
R1460 B.n541 B.n68 10.6151
R1461 B.n542 B.n541 10.6151
R1462 B.n543 B.n542 10.6151
R1463 B.n543 B.n66 10.6151
R1464 B.n547 B.n66 10.6151
R1465 B.n279 B.n278 10.6151
R1466 B.n279 B.n158 10.6151
R1467 B.n283 B.n158 10.6151
R1468 B.n284 B.n283 10.6151
R1469 B.n285 B.n284 10.6151
R1470 B.n285 B.n156 10.6151
R1471 B.n289 B.n156 10.6151
R1472 B.n290 B.n289 10.6151
R1473 B.n291 B.n290 10.6151
R1474 B.n291 B.n154 10.6151
R1475 B.n295 B.n154 10.6151
R1476 B.n296 B.n295 10.6151
R1477 B.n297 B.n296 10.6151
R1478 B.n297 B.n152 10.6151
R1479 B.n301 B.n152 10.6151
R1480 B.n302 B.n301 10.6151
R1481 B.n303 B.n302 10.6151
R1482 B.n303 B.n150 10.6151
R1483 B.n307 B.n150 10.6151
R1484 B.n308 B.n307 10.6151
R1485 B.n309 B.n308 10.6151
R1486 B.n309 B.n148 10.6151
R1487 B.n313 B.n148 10.6151
R1488 B.n316 B.n315 10.6151
R1489 B.n316 B.n144 10.6151
R1490 B.n320 B.n144 10.6151
R1491 B.n321 B.n320 10.6151
R1492 B.n322 B.n321 10.6151
R1493 B.n322 B.n142 10.6151
R1494 B.n326 B.n142 10.6151
R1495 B.n327 B.n326 10.6151
R1496 B.n328 B.n327 10.6151
R1497 B.n332 B.n331 10.6151
R1498 B.n333 B.n332 10.6151
R1499 B.n333 B.n136 10.6151
R1500 B.n337 B.n136 10.6151
R1501 B.n338 B.n337 10.6151
R1502 B.n339 B.n338 10.6151
R1503 B.n339 B.n134 10.6151
R1504 B.n343 B.n134 10.6151
R1505 B.n344 B.n343 10.6151
R1506 B.n345 B.n344 10.6151
R1507 B.n345 B.n132 10.6151
R1508 B.n349 B.n132 10.6151
R1509 B.n350 B.n349 10.6151
R1510 B.n351 B.n350 10.6151
R1511 B.n351 B.n130 10.6151
R1512 B.n355 B.n130 10.6151
R1513 B.n356 B.n355 10.6151
R1514 B.n357 B.n356 10.6151
R1515 B.n357 B.n128 10.6151
R1516 B.n361 B.n128 10.6151
R1517 B.n362 B.n361 10.6151
R1518 B.n363 B.n362 10.6151
R1519 B.n363 B.n126 10.6151
R1520 B.n277 B.n160 10.6151
R1521 B.n273 B.n160 10.6151
R1522 B.n273 B.n272 10.6151
R1523 B.n272 B.n271 10.6151
R1524 B.n271 B.n162 10.6151
R1525 B.n267 B.n162 10.6151
R1526 B.n267 B.n266 10.6151
R1527 B.n266 B.n265 10.6151
R1528 B.n265 B.n164 10.6151
R1529 B.n261 B.n164 10.6151
R1530 B.n261 B.n260 10.6151
R1531 B.n260 B.n259 10.6151
R1532 B.n259 B.n166 10.6151
R1533 B.n255 B.n166 10.6151
R1534 B.n255 B.n254 10.6151
R1535 B.n254 B.n253 10.6151
R1536 B.n253 B.n168 10.6151
R1537 B.n249 B.n168 10.6151
R1538 B.n249 B.n248 10.6151
R1539 B.n248 B.n247 10.6151
R1540 B.n247 B.n170 10.6151
R1541 B.n243 B.n170 10.6151
R1542 B.n243 B.n242 10.6151
R1543 B.n242 B.n241 10.6151
R1544 B.n241 B.n172 10.6151
R1545 B.n237 B.n172 10.6151
R1546 B.n237 B.n236 10.6151
R1547 B.n236 B.n235 10.6151
R1548 B.n235 B.n174 10.6151
R1549 B.n231 B.n174 10.6151
R1550 B.n231 B.n230 10.6151
R1551 B.n230 B.n229 10.6151
R1552 B.n229 B.n176 10.6151
R1553 B.n225 B.n176 10.6151
R1554 B.n225 B.n224 10.6151
R1555 B.n224 B.n223 10.6151
R1556 B.n223 B.n178 10.6151
R1557 B.n219 B.n178 10.6151
R1558 B.n219 B.n218 10.6151
R1559 B.n218 B.n217 10.6151
R1560 B.n217 B.n180 10.6151
R1561 B.n213 B.n180 10.6151
R1562 B.n213 B.n212 10.6151
R1563 B.n212 B.n211 10.6151
R1564 B.n211 B.n182 10.6151
R1565 B.n207 B.n182 10.6151
R1566 B.n207 B.n206 10.6151
R1567 B.n206 B.n205 10.6151
R1568 B.n205 B.n184 10.6151
R1569 B.n201 B.n184 10.6151
R1570 B.n201 B.n200 10.6151
R1571 B.n200 B.n199 10.6151
R1572 B.n199 B.n186 10.6151
R1573 B.n195 B.n186 10.6151
R1574 B.n195 B.n194 10.6151
R1575 B.n194 B.n193 10.6151
R1576 B.n193 B.n188 10.6151
R1577 B.n189 B.n188 10.6151
R1578 B.n189 B.n0 10.6151
R1579 B.n723 B.n1 10.6151
R1580 B.n723 B.n722 10.6151
R1581 B.n722 B.n721 10.6151
R1582 B.n721 B.n4 10.6151
R1583 B.n717 B.n4 10.6151
R1584 B.n717 B.n716 10.6151
R1585 B.n716 B.n715 10.6151
R1586 B.n715 B.n6 10.6151
R1587 B.n711 B.n6 10.6151
R1588 B.n711 B.n710 10.6151
R1589 B.n710 B.n709 10.6151
R1590 B.n709 B.n8 10.6151
R1591 B.n705 B.n8 10.6151
R1592 B.n705 B.n704 10.6151
R1593 B.n704 B.n703 10.6151
R1594 B.n703 B.n10 10.6151
R1595 B.n699 B.n10 10.6151
R1596 B.n699 B.n698 10.6151
R1597 B.n698 B.n697 10.6151
R1598 B.n697 B.n12 10.6151
R1599 B.n693 B.n12 10.6151
R1600 B.n693 B.n692 10.6151
R1601 B.n692 B.n691 10.6151
R1602 B.n691 B.n14 10.6151
R1603 B.n687 B.n14 10.6151
R1604 B.n687 B.n686 10.6151
R1605 B.n686 B.n685 10.6151
R1606 B.n685 B.n16 10.6151
R1607 B.n681 B.n16 10.6151
R1608 B.n681 B.n680 10.6151
R1609 B.n680 B.n679 10.6151
R1610 B.n679 B.n18 10.6151
R1611 B.n675 B.n18 10.6151
R1612 B.n675 B.n674 10.6151
R1613 B.n674 B.n673 10.6151
R1614 B.n673 B.n20 10.6151
R1615 B.n669 B.n20 10.6151
R1616 B.n669 B.n668 10.6151
R1617 B.n668 B.n667 10.6151
R1618 B.n667 B.n22 10.6151
R1619 B.n663 B.n22 10.6151
R1620 B.n663 B.n662 10.6151
R1621 B.n662 B.n661 10.6151
R1622 B.n661 B.n24 10.6151
R1623 B.n657 B.n24 10.6151
R1624 B.n657 B.n656 10.6151
R1625 B.n656 B.n655 10.6151
R1626 B.n655 B.n26 10.6151
R1627 B.n651 B.n26 10.6151
R1628 B.n651 B.n650 10.6151
R1629 B.n650 B.n649 10.6151
R1630 B.n649 B.n28 10.6151
R1631 B.n645 B.n28 10.6151
R1632 B.n645 B.n644 10.6151
R1633 B.n644 B.n643 10.6151
R1634 B.n643 B.n30 10.6151
R1635 B.n639 B.n30 10.6151
R1636 B.n639 B.n638 10.6151
R1637 B.n638 B.n637 10.6151
R1638 B.n601 B.n46 9.36635
R1639 B.n584 B.n583 9.36635
R1640 B.n314 B.n313 9.36635
R1641 B.n331 B.n140 9.36635
R1642 B.n727 B.n0 2.81026
R1643 B.n727 B.n1 2.81026
R1644 B.n598 B.n46 1.24928
R1645 B.n585 B.n584 1.24928
R1646 B.n315 B.n314 1.24928
R1647 B.n328 B.n140 1.24928
R1648 VN.n64 VN.n63 161.3
R1649 VN.n62 VN.n34 161.3
R1650 VN.n61 VN.n60 161.3
R1651 VN.n59 VN.n35 161.3
R1652 VN.n58 VN.n57 161.3
R1653 VN.n56 VN.n36 161.3
R1654 VN.n55 VN.n54 161.3
R1655 VN.n53 VN.n52 161.3
R1656 VN.n51 VN.n38 161.3
R1657 VN.n50 VN.n49 161.3
R1658 VN.n48 VN.n39 161.3
R1659 VN.n47 VN.n46 161.3
R1660 VN.n45 VN.n40 161.3
R1661 VN.n44 VN.n43 161.3
R1662 VN.n31 VN.n30 161.3
R1663 VN.n29 VN.n1 161.3
R1664 VN.n28 VN.n27 161.3
R1665 VN.n26 VN.n2 161.3
R1666 VN.n25 VN.n24 161.3
R1667 VN.n23 VN.n3 161.3
R1668 VN.n22 VN.n21 161.3
R1669 VN.n20 VN.n19 161.3
R1670 VN.n18 VN.n5 161.3
R1671 VN.n17 VN.n16 161.3
R1672 VN.n15 VN.n6 161.3
R1673 VN.n14 VN.n13 161.3
R1674 VN.n12 VN.n7 161.3
R1675 VN.n11 VN.n10 161.3
R1676 VN.n42 VN.t2 78.4388
R1677 VN.n9 VN.t7 78.4388
R1678 VN.n32 VN.n0 74.8979
R1679 VN.n65 VN.n33 74.8979
R1680 VN.n9 VN.n8 61.0251
R1681 VN.n42 VN.n41 61.0251
R1682 VN VN.n65 49.5056
R1683 VN.n8 VN.t5 45.4226
R1684 VN.n4 VN.t3 45.4226
R1685 VN.n0 VN.t4 45.4226
R1686 VN.n41 VN.t6 45.4226
R1687 VN.n37 VN.t0 45.4226
R1688 VN.n33 VN.t1 45.4226
R1689 VN.n28 VN.n2 44.3785
R1690 VN.n61 VN.n35 44.3785
R1691 VN.n13 VN.n6 40.4934
R1692 VN.n17 VN.n6 40.4934
R1693 VN.n46 VN.n39 40.4934
R1694 VN.n50 VN.n39 40.4934
R1695 VN.n24 VN.n2 36.6083
R1696 VN.n57 VN.n35 36.6083
R1697 VN.n12 VN.n11 24.4675
R1698 VN.n13 VN.n12 24.4675
R1699 VN.n18 VN.n17 24.4675
R1700 VN.n19 VN.n18 24.4675
R1701 VN.n23 VN.n22 24.4675
R1702 VN.n24 VN.n23 24.4675
R1703 VN.n29 VN.n28 24.4675
R1704 VN.n30 VN.n29 24.4675
R1705 VN.n46 VN.n45 24.4675
R1706 VN.n45 VN.n44 24.4675
R1707 VN.n57 VN.n56 24.4675
R1708 VN.n56 VN.n55 24.4675
R1709 VN.n52 VN.n51 24.4675
R1710 VN.n51 VN.n50 24.4675
R1711 VN.n63 VN.n62 24.4675
R1712 VN.n62 VN.n61 24.4675
R1713 VN.n30 VN.n0 15.17
R1714 VN.n63 VN.n33 15.17
R1715 VN.n11 VN.n8 13.2127
R1716 VN.n19 VN.n4 13.2127
R1717 VN.n44 VN.n41 13.2127
R1718 VN.n52 VN.n37 13.2127
R1719 VN.n22 VN.n4 11.2553
R1720 VN.n55 VN.n37 11.2553
R1721 VN.n43 VN.n42 4.13482
R1722 VN.n10 VN.n9 4.13482
R1723 VN.n65 VN.n64 0.354971
R1724 VN.n32 VN.n31 0.354971
R1725 VN VN.n32 0.26696
R1726 VN.n64 VN.n34 0.189894
R1727 VN.n60 VN.n34 0.189894
R1728 VN.n60 VN.n59 0.189894
R1729 VN.n59 VN.n58 0.189894
R1730 VN.n58 VN.n36 0.189894
R1731 VN.n54 VN.n36 0.189894
R1732 VN.n54 VN.n53 0.189894
R1733 VN.n53 VN.n38 0.189894
R1734 VN.n49 VN.n38 0.189894
R1735 VN.n49 VN.n48 0.189894
R1736 VN.n48 VN.n47 0.189894
R1737 VN.n47 VN.n40 0.189894
R1738 VN.n43 VN.n40 0.189894
R1739 VN.n10 VN.n7 0.189894
R1740 VN.n14 VN.n7 0.189894
R1741 VN.n15 VN.n14 0.189894
R1742 VN.n16 VN.n15 0.189894
R1743 VN.n16 VN.n5 0.189894
R1744 VN.n20 VN.n5 0.189894
R1745 VN.n21 VN.n20 0.189894
R1746 VN.n21 VN.n3 0.189894
R1747 VN.n25 VN.n3 0.189894
R1748 VN.n26 VN.n25 0.189894
R1749 VN.n27 VN.n26 0.189894
R1750 VN.n27 VN.n1 0.189894
R1751 VN.n31 VN.n1 0.189894
R1752 VDD2.n2 VDD2.n1 94.7343
R1753 VDD2.n2 VDD2.n0 94.7343
R1754 VDD2 VDD2.n5 94.7314
R1755 VDD2.n4 VDD2.n3 93.264
R1756 VDD2.n4 VDD2.n2 42.6636
R1757 VDD2.n5 VDD2.t1 5.37323
R1758 VDD2.n5 VDD2.t5 5.37323
R1759 VDD2.n3 VDD2.t6 5.37323
R1760 VDD2.n3 VDD2.t7 5.37323
R1761 VDD2.n1 VDD2.t4 5.37323
R1762 VDD2.n1 VDD2.t3 5.37323
R1763 VDD2.n0 VDD2.t0 5.37323
R1764 VDD2.n0 VDD2.t2 5.37323
R1765 VDD2 VDD2.n4 1.58455
C0 VP VN 7.30896f
C1 VN VTAIL 5.86989f
C2 VP B 2.27993f
C3 VDD1 VN 0.152498f
C4 VN w_n4510_n2178# 9.254741f
C5 VTAIL B 3.21889f
C6 VDD1 B 1.6751f
C7 w_n4510_n2178# B 9.39347f
C8 VP VTAIL 5.884f
C9 VP VDD1 5.22031f
C10 VP w_n4510_n2178# 9.84203f
C11 VDD1 VTAIL 6.490779f
C12 w_n4510_n2178# VTAIL 2.93962f
C13 VDD1 w_n4510_n2178# 1.98651f
C14 VDD2 VN 4.79026f
C15 VDD2 B 1.79032f
C16 VDD2 VP 0.584248f
C17 VDD2 VTAIL 6.54929f
C18 VDD2 VDD1 2.09286f
C19 VDD2 w_n4510_n2178# 2.12681f
C20 VN B 1.29218f
C21 VDD2 VSUBS 2.092965f
C22 VDD1 VSUBS 2.68518f
C23 VTAIL VSUBS 0.761395f
C24 VN VSUBS 7.32498f
C25 VP VSUBS 3.781534f
C26 B VSUBS 5.183002f
C27 w_n4510_n2178# VSUBS 0.122582p
C28 VDD2.t0 VSUBS 0.157596f
C29 VDD2.t2 VSUBS 0.157596f
C30 VDD2.n0 VSUBS 1.06396f
C31 VDD2.t4 VSUBS 0.157596f
C32 VDD2.t3 VSUBS 0.157596f
C33 VDD2.n1 VSUBS 1.06396f
C34 VDD2.n2 VSUBS 4.83194f
C35 VDD2.t6 VSUBS 0.157596f
C36 VDD2.t7 VSUBS 0.157596f
C37 VDD2.n3 VSUBS 1.04798f
C38 VDD2.n4 VSUBS 3.83051f
C39 VDD2.t1 VSUBS 0.157596f
C40 VDD2.t5 VSUBS 0.157596f
C41 VDD2.n5 VSUBS 1.06391f
C42 VN.t4 VSUBS 1.72372f
C43 VN.n0 VSUBS 0.768585f
C44 VN.n1 VSUBS 0.033518f
C45 VN.n2 VSUBS 0.027791f
C46 VN.n3 VSUBS 0.033518f
C47 VN.t3 VSUBS 1.72372f
C48 VN.n4 VSUBS 0.638917f
C49 VN.n5 VSUBS 0.033518f
C50 VN.n6 VSUBS 0.027096f
C51 VN.n7 VSUBS 0.033518f
C52 VN.t5 VSUBS 1.72372f
C53 VN.n8 VSUBS 0.750517f
C54 VN.t7 VSUBS 2.09222f
C55 VN.n9 VSUBS 0.714892f
C56 VN.n10 VSUBS 0.389916f
C57 VN.n11 VSUBS 0.048282f
C58 VN.n12 VSUBS 0.062469f
C59 VN.n13 VSUBS 0.066617f
C60 VN.n14 VSUBS 0.033518f
C61 VN.n15 VSUBS 0.033518f
C62 VN.n16 VSUBS 0.033518f
C63 VN.n17 VSUBS 0.066617f
C64 VN.n18 VSUBS 0.062469f
C65 VN.n19 VSUBS 0.048282f
C66 VN.n20 VSUBS 0.033518f
C67 VN.n21 VSUBS 0.033518f
C68 VN.n22 VSUBS 0.045815f
C69 VN.n23 VSUBS 0.062469f
C70 VN.n24 VSUBS 0.067581f
C71 VN.n25 VSUBS 0.033518f
C72 VN.n26 VSUBS 0.033518f
C73 VN.n27 VSUBS 0.033518f
C74 VN.n28 VSUBS 0.064957f
C75 VN.n29 VSUBS 0.062469f
C76 VN.n30 VSUBS 0.050749f
C77 VN.n31 VSUBS 0.054097f
C78 VN.n32 VSUBS 0.079222f
C79 VN.t1 VSUBS 1.72372f
C80 VN.n33 VSUBS 0.768585f
C81 VN.n34 VSUBS 0.033518f
C82 VN.n35 VSUBS 0.027791f
C83 VN.n36 VSUBS 0.033518f
C84 VN.t0 VSUBS 1.72372f
C85 VN.n37 VSUBS 0.638917f
C86 VN.n38 VSUBS 0.033518f
C87 VN.n39 VSUBS 0.027096f
C88 VN.n40 VSUBS 0.033518f
C89 VN.t6 VSUBS 1.72372f
C90 VN.n41 VSUBS 0.750517f
C91 VN.t2 VSUBS 2.09222f
C92 VN.n42 VSUBS 0.714892f
C93 VN.n43 VSUBS 0.389916f
C94 VN.n44 VSUBS 0.048282f
C95 VN.n45 VSUBS 0.062469f
C96 VN.n46 VSUBS 0.066617f
C97 VN.n47 VSUBS 0.033518f
C98 VN.n48 VSUBS 0.033518f
C99 VN.n49 VSUBS 0.033518f
C100 VN.n50 VSUBS 0.066617f
C101 VN.n51 VSUBS 0.062469f
C102 VN.n52 VSUBS 0.048282f
C103 VN.n53 VSUBS 0.033518f
C104 VN.n54 VSUBS 0.033518f
C105 VN.n55 VSUBS 0.045815f
C106 VN.n56 VSUBS 0.062469f
C107 VN.n57 VSUBS 0.067581f
C108 VN.n58 VSUBS 0.033518f
C109 VN.n59 VSUBS 0.033518f
C110 VN.n60 VSUBS 0.033518f
C111 VN.n61 VSUBS 0.064957f
C112 VN.n62 VSUBS 0.062469f
C113 VN.n63 VSUBS 0.050749f
C114 VN.n64 VSUBS 0.054097f
C115 VN.n65 VSUBS 1.88182f
C116 B.n0 VSUBS 0.005873f
C117 B.n1 VSUBS 0.005873f
C118 B.n2 VSUBS 0.009287f
C119 B.n3 VSUBS 0.009287f
C120 B.n4 VSUBS 0.009287f
C121 B.n5 VSUBS 0.009287f
C122 B.n6 VSUBS 0.009287f
C123 B.n7 VSUBS 0.009287f
C124 B.n8 VSUBS 0.009287f
C125 B.n9 VSUBS 0.009287f
C126 B.n10 VSUBS 0.009287f
C127 B.n11 VSUBS 0.009287f
C128 B.n12 VSUBS 0.009287f
C129 B.n13 VSUBS 0.009287f
C130 B.n14 VSUBS 0.009287f
C131 B.n15 VSUBS 0.009287f
C132 B.n16 VSUBS 0.009287f
C133 B.n17 VSUBS 0.009287f
C134 B.n18 VSUBS 0.009287f
C135 B.n19 VSUBS 0.009287f
C136 B.n20 VSUBS 0.009287f
C137 B.n21 VSUBS 0.009287f
C138 B.n22 VSUBS 0.009287f
C139 B.n23 VSUBS 0.009287f
C140 B.n24 VSUBS 0.009287f
C141 B.n25 VSUBS 0.009287f
C142 B.n26 VSUBS 0.009287f
C143 B.n27 VSUBS 0.009287f
C144 B.n28 VSUBS 0.009287f
C145 B.n29 VSUBS 0.009287f
C146 B.n30 VSUBS 0.009287f
C147 B.n31 VSUBS 0.009287f
C148 B.n32 VSUBS 0.022737f
C149 B.n33 VSUBS 0.009287f
C150 B.n34 VSUBS 0.009287f
C151 B.n35 VSUBS 0.009287f
C152 B.n36 VSUBS 0.009287f
C153 B.n37 VSUBS 0.009287f
C154 B.n38 VSUBS 0.009287f
C155 B.n39 VSUBS 0.009287f
C156 B.n40 VSUBS 0.009287f
C157 B.n41 VSUBS 0.009287f
C158 B.n42 VSUBS 0.009287f
C159 B.n43 VSUBS 0.009287f
C160 B.t8 VSUBS 0.120037f
C161 B.t7 VSUBS 0.160428f
C162 B.t6 VSUBS 1.22997f
C163 B.n44 VSUBS 0.268368f
C164 B.n45 VSUBS 0.211991f
C165 B.n46 VSUBS 0.021517f
C166 B.n47 VSUBS 0.009287f
C167 B.n48 VSUBS 0.009287f
C168 B.n49 VSUBS 0.009287f
C169 B.n50 VSUBS 0.009287f
C170 B.n51 VSUBS 0.009287f
C171 B.t11 VSUBS 0.120039f
C172 B.t10 VSUBS 0.160429f
C173 B.t9 VSUBS 1.22997f
C174 B.n52 VSUBS 0.268366f
C175 B.n53 VSUBS 0.211988f
C176 B.n54 VSUBS 0.009287f
C177 B.n55 VSUBS 0.009287f
C178 B.n56 VSUBS 0.009287f
C179 B.n57 VSUBS 0.009287f
C180 B.n58 VSUBS 0.009287f
C181 B.n59 VSUBS 0.009287f
C182 B.n60 VSUBS 0.009287f
C183 B.n61 VSUBS 0.009287f
C184 B.n62 VSUBS 0.009287f
C185 B.n63 VSUBS 0.009287f
C186 B.n64 VSUBS 0.009287f
C187 B.n65 VSUBS 0.022737f
C188 B.n66 VSUBS 0.009287f
C189 B.n67 VSUBS 0.009287f
C190 B.n68 VSUBS 0.009287f
C191 B.n69 VSUBS 0.009287f
C192 B.n70 VSUBS 0.009287f
C193 B.n71 VSUBS 0.009287f
C194 B.n72 VSUBS 0.009287f
C195 B.n73 VSUBS 0.009287f
C196 B.n74 VSUBS 0.009287f
C197 B.n75 VSUBS 0.009287f
C198 B.n76 VSUBS 0.009287f
C199 B.n77 VSUBS 0.009287f
C200 B.n78 VSUBS 0.009287f
C201 B.n79 VSUBS 0.009287f
C202 B.n80 VSUBS 0.009287f
C203 B.n81 VSUBS 0.009287f
C204 B.n82 VSUBS 0.009287f
C205 B.n83 VSUBS 0.009287f
C206 B.n84 VSUBS 0.009287f
C207 B.n85 VSUBS 0.009287f
C208 B.n86 VSUBS 0.009287f
C209 B.n87 VSUBS 0.009287f
C210 B.n88 VSUBS 0.009287f
C211 B.n89 VSUBS 0.009287f
C212 B.n90 VSUBS 0.009287f
C213 B.n91 VSUBS 0.009287f
C214 B.n92 VSUBS 0.009287f
C215 B.n93 VSUBS 0.009287f
C216 B.n94 VSUBS 0.009287f
C217 B.n95 VSUBS 0.009287f
C218 B.n96 VSUBS 0.009287f
C219 B.n97 VSUBS 0.009287f
C220 B.n98 VSUBS 0.009287f
C221 B.n99 VSUBS 0.009287f
C222 B.n100 VSUBS 0.009287f
C223 B.n101 VSUBS 0.009287f
C224 B.n102 VSUBS 0.009287f
C225 B.n103 VSUBS 0.009287f
C226 B.n104 VSUBS 0.009287f
C227 B.n105 VSUBS 0.009287f
C228 B.n106 VSUBS 0.009287f
C229 B.n107 VSUBS 0.009287f
C230 B.n108 VSUBS 0.009287f
C231 B.n109 VSUBS 0.009287f
C232 B.n110 VSUBS 0.009287f
C233 B.n111 VSUBS 0.009287f
C234 B.n112 VSUBS 0.009287f
C235 B.n113 VSUBS 0.009287f
C236 B.n114 VSUBS 0.009287f
C237 B.n115 VSUBS 0.009287f
C238 B.n116 VSUBS 0.009287f
C239 B.n117 VSUBS 0.009287f
C240 B.n118 VSUBS 0.009287f
C241 B.n119 VSUBS 0.009287f
C242 B.n120 VSUBS 0.009287f
C243 B.n121 VSUBS 0.009287f
C244 B.n122 VSUBS 0.009287f
C245 B.n123 VSUBS 0.009287f
C246 B.n124 VSUBS 0.009287f
C247 B.n125 VSUBS 0.009287f
C248 B.n126 VSUBS 0.022737f
C249 B.n127 VSUBS 0.009287f
C250 B.n128 VSUBS 0.009287f
C251 B.n129 VSUBS 0.009287f
C252 B.n130 VSUBS 0.009287f
C253 B.n131 VSUBS 0.009287f
C254 B.n132 VSUBS 0.009287f
C255 B.n133 VSUBS 0.009287f
C256 B.n134 VSUBS 0.009287f
C257 B.n135 VSUBS 0.009287f
C258 B.n136 VSUBS 0.009287f
C259 B.n137 VSUBS 0.009287f
C260 B.t4 VSUBS 0.120039f
C261 B.t5 VSUBS 0.160429f
C262 B.t3 VSUBS 1.22997f
C263 B.n138 VSUBS 0.268366f
C264 B.n139 VSUBS 0.211988f
C265 B.n140 VSUBS 0.021517f
C266 B.n141 VSUBS 0.009287f
C267 B.n142 VSUBS 0.009287f
C268 B.n143 VSUBS 0.009287f
C269 B.n144 VSUBS 0.009287f
C270 B.n145 VSUBS 0.009287f
C271 B.t1 VSUBS 0.120037f
C272 B.t2 VSUBS 0.160428f
C273 B.t0 VSUBS 1.22997f
C274 B.n146 VSUBS 0.268368f
C275 B.n147 VSUBS 0.211991f
C276 B.n148 VSUBS 0.009287f
C277 B.n149 VSUBS 0.009287f
C278 B.n150 VSUBS 0.009287f
C279 B.n151 VSUBS 0.009287f
C280 B.n152 VSUBS 0.009287f
C281 B.n153 VSUBS 0.009287f
C282 B.n154 VSUBS 0.009287f
C283 B.n155 VSUBS 0.009287f
C284 B.n156 VSUBS 0.009287f
C285 B.n157 VSUBS 0.009287f
C286 B.n158 VSUBS 0.009287f
C287 B.n159 VSUBS 0.022737f
C288 B.n160 VSUBS 0.009287f
C289 B.n161 VSUBS 0.009287f
C290 B.n162 VSUBS 0.009287f
C291 B.n163 VSUBS 0.009287f
C292 B.n164 VSUBS 0.009287f
C293 B.n165 VSUBS 0.009287f
C294 B.n166 VSUBS 0.009287f
C295 B.n167 VSUBS 0.009287f
C296 B.n168 VSUBS 0.009287f
C297 B.n169 VSUBS 0.009287f
C298 B.n170 VSUBS 0.009287f
C299 B.n171 VSUBS 0.009287f
C300 B.n172 VSUBS 0.009287f
C301 B.n173 VSUBS 0.009287f
C302 B.n174 VSUBS 0.009287f
C303 B.n175 VSUBS 0.009287f
C304 B.n176 VSUBS 0.009287f
C305 B.n177 VSUBS 0.009287f
C306 B.n178 VSUBS 0.009287f
C307 B.n179 VSUBS 0.009287f
C308 B.n180 VSUBS 0.009287f
C309 B.n181 VSUBS 0.009287f
C310 B.n182 VSUBS 0.009287f
C311 B.n183 VSUBS 0.009287f
C312 B.n184 VSUBS 0.009287f
C313 B.n185 VSUBS 0.009287f
C314 B.n186 VSUBS 0.009287f
C315 B.n187 VSUBS 0.009287f
C316 B.n188 VSUBS 0.009287f
C317 B.n189 VSUBS 0.009287f
C318 B.n190 VSUBS 0.009287f
C319 B.n191 VSUBS 0.009287f
C320 B.n192 VSUBS 0.009287f
C321 B.n193 VSUBS 0.009287f
C322 B.n194 VSUBS 0.009287f
C323 B.n195 VSUBS 0.009287f
C324 B.n196 VSUBS 0.009287f
C325 B.n197 VSUBS 0.009287f
C326 B.n198 VSUBS 0.009287f
C327 B.n199 VSUBS 0.009287f
C328 B.n200 VSUBS 0.009287f
C329 B.n201 VSUBS 0.009287f
C330 B.n202 VSUBS 0.009287f
C331 B.n203 VSUBS 0.009287f
C332 B.n204 VSUBS 0.009287f
C333 B.n205 VSUBS 0.009287f
C334 B.n206 VSUBS 0.009287f
C335 B.n207 VSUBS 0.009287f
C336 B.n208 VSUBS 0.009287f
C337 B.n209 VSUBS 0.009287f
C338 B.n210 VSUBS 0.009287f
C339 B.n211 VSUBS 0.009287f
C340 B.n212 VSUBS 0.009287f
C341 B.n213 VSUBS 0.009287f
C342 B.n214 VSUBS 0.009287f
C343 B.n215 VSUBS 0.009287f
C344 B.n216 VSUBS 0.009287f
C345 B.n217 VSUBS 0.009287f
C346 B.n218 VSUBS 0.009287f
C347 B.n219 VSUBS 0.009287f
C348 B.n220 VSUBS 0.009287f
C349 B.n221 VSUBS 0.009287f
C350 B.n222 VSUBS 0.009287f
C351 B.n223 VSUBS 0.009287f
C352 B.n224 VSUBS 0.009287f
C353 B.n225 VSUBS 0.009287f
C354 B.n226 VSUBS 0.009287f
C355 B.n227 VSUBS 0.009287f
C356 B.n228 VSUBS 0.009287f
C357 B.n229 VSUBS 0.009287f
C358 B.n230 VSUBS 0.009287f
C359 B.n231 VSUBS 0.009287f
C360 B.n232 VSUBS 0.009287f
C361 B.n233 VSUBS 0.009287f
C362 B.n234 VSUBS 0.009287f
C363 B.n235 VSUBS 0.009287f
C364 B.n236 VSUBS 0.009287f
C365 B.n237 VSUBS 0.009287f
C366 B.n238 VSUBS 0.009287f
C367 B.n239 VSUBS 0.009287f
C368 B.n240 VSUBS 0.009287f
C369 B.n241 VSUBS 0.009287f
C370 B.n242 VSUBS 0.009287f
C371 B.n243 VSUBS 0.009287f
C372 B.n244 VSUBS 0.009287f
C373 B.n245 VSUBS 0.009287f
C374 B.n246 VSUBS 0.009287f
C375 B.n247 VSUBS 0.009287f
C376 B.n248 VSUBS 0.009287f
C377 B.n249 VSUBS 0.009287f
C378 B.n250 VSUBS 0.009287f
C379 B.n251 VSUBS 0.009287f
C380 B.n252 VSUBS 0.009287f
C381 B.n253 VSUBS 0.009287f
C382 B.n254 VSUBS 0.009287f
C383 B.n255 VSUBS 0.009287f
C384 B.n256 VSUBS 0.009287f
C385 B.n257 VSUBS 0.009287f
C386 B.n258 VSUBS 0.009287f
C387 B.n259 VSUBS 0.009287f
C388 B.n260 VSUBS 0.009287f
C389 B.n261 VSUBS 0.009287f
C390 B.n262 VSUBS 0.009287f
C391 B.n263 VSUBS 0.009287f
C392 B.n264 VSUBS 0.009287f
C393 B.n265 VSUBS 0.009287f
C394 B.n266 VSUBS 0.009287f
C395 B.n267 VSUBS 0.009287f
C396 B.n268 VSUBS 0.009287f
C397 B.n269 VSUBS 0.009287f
C398 B.n270 VSUBS 0.009287f
C399 B.n271 VSUBS 0.009287f
C400 B.n272 VSUBS 0.009287f
C401 B.n273 VSUBS 0.009287f
C402 B.n274 VSUBS 0.009287f
C403 B.n275 VSUBS 0.009287f
C404 B.n276 VSUBS 0.021239f
C405 B.n277 VSUBS 0.021239f
C406 B.n278 VSUBS 0.022737f
C407 B.n279 VSUBS 0.009287f
C408 B.n280 VSUBS 0.009287f
C409 B.n281 VSUBS 0.009287f
C410 B.n282 VSUBS 0.009287f
C411 B.n283 VSUBS 0.009287f
C412 B.n284 VSUBS 0.009287f
C413 B.n285 VSUBS 0.009287f
C414 B.n286 VSUBS 0.009287f
C415 B.n287 VSUBS 0.009287f
C416 B.n288 VSUBS 0.009287f
C417 B.n289 VSUBS 0.009287f
C418 B.n290 VSUBS 0.009287f
C419 B.n291 VSUBS 0.009287f
C420 B.n292 VSUBS 0.009287f
C421 B.n293 VSUBS 0.009287f
C422 B.n294 VSUBS 0.009287f
C423 B.n295 VSUBS 0.009287f
C424 B.n296 VSUBS 0.009287f
C425 B.n297 VSUBS 0.009287f
C426 B.n298 VSUBS 0.009287f
C427 B.n299 VSUBS 0.009287f
C428 B.n300 VSUBS 0.009287f
C429 B.n301 VSUBS 0.009287f
C430 B.n302 VSUBS 0.009287f
C431 B.n303 VSUBS 0.009287f
C432 B.n304 VSUBS 0.009287f
C433 B.n305 VSUBS 0.009287f
C434 B.n306 VSUBS 0.009287f
C435 B.n307 VSUBS 0.009287f
C436 B.n308 VSUBS 0.009287f
C437 B.n309 VSUBS 0.009287f
C438 B.n310 VSUBS 0.009287f
C439 B.n311 VSUBS 0.009287f
C440 B.n312 VSUBS 0.009287f
C441 B.n313 VSUBS 0.008741f
C442 B.n314 VSUBS 0.021517f
C443 B.n315 VSUBS 0.00519f
C444 B.n316 VSUBS 0.009287f
C445 B.n317 VSUBS 0.009287f
C446 B.n318 VSUBS 0.009287f
C447 B.n319 VSUBS 0.009287f
C448 B.n320 VSUBS 0.009287f
C449 B.n321 VSUBS 0.009287f
C450 B.n322 VSUBS 0.009287f
C451 B.n323 VSUBS 0.009287f
C452 B.n324 VSUBS 0.009287f
C453 B.n325 VSUBS 0.009287f
C454 B.n326 VSUBS 0.009287f
C455 B.n327 VSUBS 0.009287f
C456 B.n328 VSUBS 0.00519f
C457 B.n329 VSUBS 0.009287f
C458 B.n330 VSUBS 0.009287f
C459 B.n331 VSUBS 0.008741f
C460 B.n332 VSUBS 0.009287f
C461 B.n333 VSUBS 0.009287f
C462 B.n334 VSUBS 0.009287f
C463 B.n335 VSUBS 0.009287f
C464 B.n336 VSUBS 0.009287f
C465 B.n337 VSUBS 0.009287f
C466 B.n338 VSUBS 0.009287f
C467 B.n339 VSUBS 0.009287f
C468 B.n340 VSUBS 0.009287f
C469 B.n341 VSUBS 0.009287f
C470 B.n342 VSUBS 0.009287f
C471 B.n343 VSUBS 0.009287f
C472 B.n344 VSUBS 0.009287f
C473 B.n345 VSUBS 0.009287f
C474 B.n346 VSUBS 0.009287f
C475 B.n347 VSUBS 0.009287f
C476 B.n348 VSUBS 0.009287f
C477 B.n349 VSUBS 0.009287f
C478 B.n350 VSUBS 0.009287f
C479 B.n351 VSUBS 0.009287f
C480 B.n352 VSUBS 0.009287f
C481 B.n353 VSUBS 0.009287f
C482 B.n354 VSUBS 0.009287f
C483 B.n355 VSUBS 0.009287f
C484 B.n356 VSUBS 0.009287f
C485 B.n357 VSUBS 0.009287f
C486 B.n358 VSUBS 0.009287f
C487 B.n359 VSUBS 0.009287f
C488 B.n360 VSUBS 0.009287f
C489 B.n361 VSUBS 0.009287f
C490 B.n362 VSUBS 0.009287f
C491 B.n363 VSUBS 0.009287f
C492 B.n364 VSUBS 0.009287f
C493 B.n365 VSUBS 0.022737f
C494 B.n366 VSUBS 0.021239f
C495 B.n367 VSUBS 0.021239f
C496 B.n368 VSUBS 0.009287f
C497 B.n369 VSUBS 0.009287f
C498 B.n370 VSUBS 0.009287f
C499 B.n371 VSUBS 0.009287f
C500 B.n372 VSUBS 0.009287f
C501 B.n373 VSUBS 0.009287f
C502 B.n374 VSUBS 0.009287f
C503 B.n375 VSUBS 0.009287f
C504 B.n376 VSUBS 0.009287f
C505 B.n377 VSUBS 0.009287f
C506 B.n378 VSUBS 0.009287f
C507 B.n379 VSUBS 0.009287f
C508 B.n380 VSUBS 0.009287f
C509 B.n381 VSUBS 0.009287f
C510 B.n382 VSUBS 0.009287f
C511 B.n383 VSUBS 0.009287f
C512 B.n384 VSUBS 0.009287f
C513 B.n385 VSUBS 0.009287f
C514 B.n386 VSUBS 0.009287f
C515 B.n387 VSUBS 0.009287f
C516 B.n388 VSUBS 0.009287f
C517 B.n389 VSUBS 0.009287f
C518 B.n390 VSUBS 0.009287f
C519 B.n391 VSUBS 0.009287f
C520 B.n392 VSUBS 0.009287f
C521 B.n393 VSUBS 0.009287f
C522 B.n394 VSUBS 0.009287f
C523 B.n395 VSUBS 0.009287f
C524 B.n396 VSUBS 0.009287f
C525 B.n397 VSUBS 0.009287f
C526 B.n398 VSUBS 0.009287f
C527 B.n399 VSUBS 0.009287f
C528 B.n400 VSUBS 0.009287f
C529 B.n401 VSUBS 0.009287f
C530 B.n402 VSUBS 0.009287f
C531 B.n403 VSUBS 0.009287f
C532 B.n404 VSUBS 0.009287f
C533 B.n405 VSUBS 0.009287f
C534 B.n406 VSUBS 0.009287f
C535 B.n407 VSUBS 0.009287f
C536 B.n408 VSUBS 0.009287f
C537 B.n409 VSUBS 0.009287f
C538 B.n410 VSUBS 0.009287f
C539 B.n411 VSUBS 0.009287f
C540 B.n412 VSUBS 0.009287f
C541 B.n413 VSUBS 0.009287f
C542 B.n414 VSUBS 0.009287f
C543 B.n415 VSUBS 0.009287f
C544 B.n416 VSUBS 0.009287f
C545 B.n417 VSUBS 0.009287f
C546 B.n418 VSUBS 0.009287f
C547 B.n419 VSUBS 0.009287f
C548 B.n420 VSUBS 0.009287f
C549 B.n421 VSUBS 0.009287f
C550 B.n422 VSUBS 0.009287f
C551 B.n423 VSUBS 0.009287f
C552 B.n424 VSUBS 0.009287f
C553 B.n425 VSUBS 0.009287f
C554 B.n426 VSUBS 0.009287f
C555 B.n427 VSUBS 0.009287f
C556 B.n428 VSUBS 0.009287f
C557 B.n429 VSUBS 0.009287f
C558 B.n430 VSUBS 0.009287f
C559 B.n431 VSUBS 0.009287f
C560 B.n432 VSUBS 0.009287f
C561 B.n433 VSUBS 0.009287f
C562 B.n434 VSUBS 0.009287f
C563 B.n435 VSUBS 0.009287f
C564 B.n436 VSUBS 0.009287f
C565 B.n437 VSUBS 0.009287f
C566 B.n438 VSUBS 0.009287f
C567 B.n439 VSUBS 0.009287f
C568 B.n440 VSUBS 0.009287f
C569 B.n441 VSUBS 0.009287f
C570 B.n442 VSUBS 0.009287f
C571 B.n443 VSUBS 0.009287f
C572 B.n444 VSUBS 0.009287f
C573 B.n445 VSUBS 0.009287f
C574 B.n446 VSUBS 0.009287f
C575 B.n447 VSUBS 0.009287f
C576 B.n448 VSUBS 0.009287f
C577 B.n449 VSUBS 0.009287f
C578 B.n450 VSUBS 0.009287f
C579 B.n451 VSUBS 0.009287f
C580 B.n452 VSUBS 0.009287f
C581 B.n453 VSUBS 0.009287f
C582 B.n454 VSUBS 0.009287f
C583 B.n455 VSUBS 0.009287f
C584 B.n456 VSUBS 0.009287f
C585 B.n457 VSUBS 0.009287f
C586 B.n458 VSUBS 0.009287f
C587 B.n459 VSUBS 0.009287f
C588 B.n460 VSUBS 0.009287f
C589 B.n461 VSUBS 0.009287f
C590 B.n462 VSUBS 0.009287f
C591 B.n463 VSUBS 0.009287f
C592 B.n464 VSUBS 0.009287f
C593 B.n465 VSUBS 0.009287f
C594 B.n466 VSUBS 0.009287f
C595 B.n467 VSUBS 0.009287f
C596 B.n468 VSUBS 0.009287f
C597 B.n469 VSUBS 0.009287f
C598 B.n470 VSUBS 0.009287f
C599 B.n471 VSUBS 0.009287f
C600 B.n472 VSUBS 0.009287f
C601 B.n473 VSUBS 0.009287f
C602 B.n474 VSUBS 0.009287f
C603 B.n475 VSUBS 0.009287f
C604 B.n476 VSUBS 0.009287f
C605 B.n477 VSUBS 0.009287f
C606 B.n478 VSUBS 0.009287f
C607 B.n479 VSUBS 0.009287f
C608 B.n480 VSUBS 0.009287f
C609 B.n481 VSUBS 0.009287f
C610 B.n482 VSUBS 0.009287f
C611 B.n483 VSUBS 0.009287f
C612 B.n484 VSUBS 0.009287f
C613 B.n485 VSUBS 0.009287f
C614 B.n486 VSUBS 0.009287f
C615 B.n487 VSUBS 0.009287f
C616 B.n488 VSUBS 0.009287f
C617 B.n489 VSUBS 0.009287f
C618 B.n490 VSUBS 0.009287f
C619 B.n491 VSUBS 0.009287f
C620 B.n492 VSUBS 0.009287f
C621 B.n493 VSUBS 0.009287f
C622 B.n494 VSUBS 0.009287f
C623 B.n495 VSUBS 0.009287f
C624 B.n496 VSUBS 0.009287f
C625 B.n497 VSUBS 0.009287f
C626 B.n498 VSUBS 0.009287f
C627 B.n499 VSUBS 0.009287f
C628 B.n500 VSUBS 0.009287f
C629 B.n501 VSUBS 0.009287f
C630 B.n502 VSUBS 0.009287f
C631 B.n503 VSUBS 0.009287f
C632 B.n504 VSUBS 0.009287f
C633 B.n505 VSUBS 0.009287f
C634 B.n506 VSUBS 0.009287f
C635 B.n507 VSUBS 0.009287f
C636 B.n508 VSUBS 0.009287f
C637 B.n509 VSUBS 0.009287f
C638 B.n510 VSUBS 0.009287f
C639 B.n511 VSUBS 0.009287f
C640 B.n512 VSUBS 0.009287f
C641 B.n513 VSUBS 0.009287f
C642 B.n514 VSUBS 0.009287f
C643 B.n515 VSUBS 0.009287f
C644 B.n516 VSUBS 0.009287f
C645 B.n517 VSUBS 0.009287f
C646 B.n518 VSUBS 0.009287f
C647 B.n519 VSUBS 0.009287f
C648 B.n520 VSUBS 0.009287f
C649 B.n521 VSUBS 0.009287f
C650 B.n522 VSUBS 0.009287f
C651 B.n523 VSUBS 0.009287f
C652 B.n524 VSUBS 0.009287f
C653 B.n525 VSUBS 0.009287f
C654 B.n526 VSUBS 0.009287f
C655 B.n527 VSUBS 0.009287f
C656 B.n528 VSUBS 0.009287f
C657 B.n529 VSUBS 0.009287f
C658 B.n530 VSUBS 0.009287f
C659 B.n531 VSUBS 0.009287f
C660 B.n532 VSUBS 0.009287f
C661 B.n533 VSUBS 0.009287f
C662 B.n534 VSUBS 0.009287f
C663 B.n535 VSUBS 0.009287f
C664 B.n536 VSUBS 0.009287f
C665 B.n537 VSUBS 0.009287f
C666 B.n538 VSUBS 0.009287f
C667 B.n539 VSUBS 0.009287f
C668 B.n540 VSUBS 0.009287f
C669 B.n541 VSUBS 0.009287f
C670 B.n542 VSUBS 0.009287f
C671 B.n543 VSUBS 0.009287f
C672 B.n544 VSUBS 0.009287f
C673 B.n545 VSUBS 0.009287f
C674 B.n546 VSUBS 0.021239f
C675 B.n547 VSUBS 0.022317f
C676 B.n548 VSUBS 0.02166f
C677 B.n549 VSUBS 0.009287f
C678 B.n550 VSUBS 0.009287f
C679 B.n551 VSUBS 0.009287f
C680 B.n552 VSUBS 0.009287f
C681 B.n553 VSUBS 0.009287f
C682 B.n554 VSUBS 0.009287f
C683 B.n555 VSUBS 0.009287f
C684 B.n556 VSUBS 0.009287f
C685 B.n557 VSUBS 0.009287f
C686 B.n558 VSUBS 0.009287f
C687 B.n559 VSUBS 0.009287f
C688 B.n560 VSUBS 0.009287f
C689 B.n561 VSUBS 0.009287f
C690 B.n562 VSUBS 0.009287f
C691 B.n563 VSUBS 0.009287f
C692 B.n564 VSUBS 0.009287f
C693 B.n565 VSUBS 0.009287f
C694 B.n566 VSUBS 0.009287f
C695 B.n567 VSUBS 0.009287f
C696 B.n568 VSUBS 0.009287f
C697 B.n569 VSUBS 0.009287f
C698 B.n570 VSUBS 0.009287f
C699 B.n571 VSUBS 0.009287f
C700 B.n572 VSUBS 0.009287f
C701 B.n573 VSUBS 0.009287f
C702 B.n574 VSUBS 0.009287f
C703 B.n575 VSUBS 0.009287f
C704 B.n576 VSUBS 0.009287f
C705 B.n577 VSUBS 0.009287f
C706 B.n578 VSUBS 0.009287f
C707 B.n579 VSUBS 0.009287f
C708 B.n580 VSUBS 0.009287f
C709 B.n581 VSUBS 0.009287f
C710 B.n582 VSUBS 0.009287f
C711 B.n583 VSUBS 0.008741f
C712 B.n584 VSUBS 0.021517f
C713 B.n585 VSUBS 0.00519f
C714 B.n586 VSUBS 0.009287f
C715 B.n587 VSUBS 0.009287f
C716 B.n588 VSUBS 0.009287f
C717 B.n589 VSUBS 0.009287f
C718 B.n590 VSUBS 0.009287f
C719 B.n591 VSUBS 0.009287f
C720 B.n592 VSUBS 0.009287f
C721 B.n593 VSUBS 0.009287f
C722 B.n594 VSUBS 0.009287f
C723 B.n595 VSUBS 0.009287f
C724 B.n596 VSUBS 0.009287f
C725 B.n597 VSUBS 0.009287f
C726 B.n598 VSUBS 0.00519f
C727 B.n599 VSUBS 0.009287f
C728 B.n600 VSUBS 0.009287f
C729 B.n601 VSUBS 0.008741f
C730 B.n602 VSUBS 0.009287f
C731 B.n603 VSUBS 0.009287f
C732 B.n604 VSUBS 0.009287f
C733 B.n605 VSUBS 0.009287f
C734 B.n606 VSUBS 0.009287f
C735 B.n607 VSUBS 0.009287f
C736 B.n608 VSUBS 0.009287f
C737 B.n609 VSUBS 0.009287f
C738 B.n610 VSUBS 0.009287f
C739 B.n611 VSUBS 0.009287f
C740 B.n612 VSUBS 0.009287f
C741 B.n613 VSUBS 0.009287f
C742 B.n614 VSUBS 0.009287f
C743 B.n615 VSUBS 0.009287f
C744 B.n616 VSUBS 0.009287f
C745 B.n617 VSUBS 0.009287f
C746 B.n618 VSUBS 0.009287f
C747 B.n619 VSUBS 0.009287f
C748 B.n620 VSUBS 0.009287f
C749 B.n621 VSUBS 0.009287f
C750 B.n622 VSUBS 0.009287f
C751 B.n623 VSUBS 0.009287f
C752 B.n624 VSUBS 0.009287f
C753 B.n625 VSUBS 0.009287f
C754 B.n626 VSUBS 0.009287f
C755 B.n627 VSUBS 0.009287f
C756 B.n628 VSUBS 0.009287f
C757 B.n629 VSUBS 0.009287f
C758 B.n630 VSUBS 0.009287f
C759 B.n631 VSUBS 0.009287f
C760 B.n632 VSUBS 0.009287f
C761 B.n633 VSUBS 0.009287f
C762 B.n634 VSUBS 0.009287f
C763 B.n635 VSUBS 0.022737f
C764 B.n636 VSUBS 0.021239f
C765 B.n637 VSUBS 0.021239f
C766 B.n638 VSUBS 0.009287f
C767 B.n639 VSUBS 0.009287f
C768 B.n640 VSUBS 0.009287f
C769 B.n641 VSUBS 0.009287f
C770 B.n642 VSUBS 0.009287f
C771 B.n643 VSUBS 0.009287f
C772 B.n644 VSUBS 0.009287f
C773 B.n645 VSUBS 0.009287f
C774 B.n646 VSUBS 0.009287f
C775 B.n647 VSUBS 0.009287f
C776 B.n648 VSUBS 0.009287f
C777 B.n649 VSUBS 0.009287f
C778 B.n650 VSUBS 0.009287f
C779 B.n651 VSUBS 0.009287f
C780 B.n652 VSUBS 0.009287f
C781 B.n653 VSUBS 0.009287f
C782 B.n654 VSUBS 0.009287f
C783 B.n655 VSUBS 0.009287f
C784 B.n656 VSUBS 0.009287f
C785 B.n657 VSUBS 0.009287f
C786 B.n658 VSUBS 0.009287f
C787 B.n659 VSUBS 0.009287f
C788 B.n660 VSUBS 0.009287f
C789 B.n661 VSUBS 0.009287f
C790 B.n662 VSUBS 0.009287f
C791 B.n663 VSUBS 0.009287f
C792 B.n664 VSUBS 0.009287f
C793 B.n665 VSUBS 0.009287f
C794 B.n666 VSUBS 0.009287f
C795 B.n667 VSUBS 0.009287f
C796 B.n668 VSUBS 0.009287f
C797 B.n669 VSUBS 0.009287f
C798 B.n670 VSUBS 0.009287f
C799 B.n671 VSUBS 0.009287f
C800 B.n672 VSUBS 0.009287f
C801 B.n673 VSUBS 0.009287f
C802 B.n674 VSUBS 0.009287f
C803 B.n675 VSUBS 0.009287f
C804 B.n676 VSUBS 0.009287f
C805 B.n677 VSUBS 0.009287f
C806 B.n678 VSUBS 0.009287f
C807 B.n679 VSUBS 0.009287f
C808 B.n680 VSUBS 0.009287f
C809 B.n681 VSUBS 0.009287f
C810 B.n682 VSUBS 0.009287f
C811 B.n683 VSUBS 0.009287f
C812 B.n684 VSUBS 0.009287f
C813 B.n685 VSUBS 0.009287f
C814 B.n686 VSUBS 0.009287f
C815 B.n687 VSUBS 0.009287f
C816 B.n688 VSUBS 0.009287f
C817 B.n689 VSUBS 0.009287f
C818 B.n690 VSUBS 0.009287f
C819 B.n691 VSUBS 0.009287f
C820 B.n692 VSUBS 0.009287f
C821 B.n693 VSUBS 0.009287f
C822 B.n694 VSUBS 0.009287f
C823 B.n695 VSUBS 0.009287f
C824 B.n696 VSUBS 0.009287f
C825 B.n697 VSUBS 0.009287f
C826 B.n698 VSUBS 0.009287f
C827 B.n699 VSUBS 0.009287f
C828 B.n700 VSUBS 0.009287f
C829 B.n701 VSUBS 0.009287f
C830 B.n702 VSUBS 0.009287f
C831 B.n703 VSUBS 0.009287f
C832 B.n704 VSUBS 0.009287f
C833 B.n705 VSUBS 0.009287f
C834 B.n706 VSUBS 0.009287f
C835 B.n707 VSUBS 0.009287f
C836 B.n708 VSUBS 0.009287f
C837 B.n709 VSUBS 0.009287f
C838 B.n710 VSUBS 0.009287f
C839 B.n711 VSUBS 0.009287f
C840 B.n712 VSUBS 0.009287f
C841 B.n713 VSUBS 0.009287f
C842 B.n714 VSUBS 0.009287f
C843 B.n715 VSUBS 0.009287f
C844 B.n716 VSUBS 0.009287f
C845 B.n717 VSUBS 0.009287f
C846 B.n718 VSUBS 0.009287f
C847 B.n719 VSUBS 0.009287f
C848 B.n720 VSUBS 0.009287f
C849 B.n721 VSUBS 0.009287f
C850 B.n722 VSUBS 0.009287f
C851 B.n723 VSUBS 0.009287f
C852 B.n724 VSUBS 0.009287f
C853 B.n725 VSUBS 0.009287f
C854 B.n726 VSUBS 0.009287f
C855 B.n727 VSUBS 0.021029f
C856 VDD1.t1 VSUBS 0.139218f
C857 VDD1.t7 VSUBS 0.139218f
C858 VDD1.n0 VSUBS 0.941128f
C859 VDD1.t0 VSUBS 0.139218f
C860 VDD1.t5 VSUBS 0.139218f
C861 VDD1.n1 VSUBS 0.939881f
C862 VDD1.t4 VSUBS 0.139218f
C863 VDD1.t2 VSUBS 0.139218f
C864 VDD1.n2 VSUBS 0.939881f
C865 VDD1.n3 VSUBS 4.32892f
C866 VDD1.t6 VSUBS 0.139218f
C867 VDD1.t3 VSUBS 0.139218f
C868 VDD1.n4 VSUBS 0.925763f
C869 VDD1.n5 VSUBS 3.41998f
C870 VTAIL.t3 VSUBS 0.143852f
C871 VTAIL.t5 VSUBS 0.143852f
C872 VTAIL.n0 VSUBS 0.851384f
C873 VTAIL.n1 VSUBS 0.854576f
C874 VTAIL.n2 VSUBS 0.033573f
C875 VTAIL.n3 VSUBS 0.030089f
C876 VTAIL.n4 VSUBS 0.016169f
C877 VTAIL.n5 VSUBS 0.038216f
C878 VTAIL.n6 VSUBS 0.01712f
C879 VTAIL.n7 VSUBS 0.030089f
C880 VTAIL.n8 VSUBS 0.016169f
C881 VTAIL.n9 VSUBS 0.038216f
C882 VTAIL.n10 VSUBS 0.01712f
C883 VTAIL.n11 VSUBS 0.133563f
C884 VTAIL.t0 VSUBS 0.082088f
C885 VTAIL.n12 VSUBS 0.028662f
C886 VTAIL.n13 VSUBS 0.024299f
C887 VTAIL.n14 VSUBS 0.016169f
C888 VTAIL.n15 VSUBS 0.696889f
C889 VTAIL.n16 VSUBS 0.030089f
C890 VTAIL.n17 VSUBS 0.016169f
C891 VTAIL.n18 VSUBS 0.01712f
C892 VTAIL.n19 VSUBS 0.038216f
C893 VTAIL.n20 VSUBS 0.038216f
C894 VTAIL.n21 VSUBS 0.01712f
C895 VTAIL.n22 VSUBS 0.016169f
C896 VTAIL.n23 VSUBS 0.030089f
C897 VTAIL.n24 VSUBS 0.030089f
C898 VTAIL.n25 VSUBS 0.016169f
C899 VTAIL.n26 VSUBS 0.01712f
C900 VTAIL.n27 VSUBS 0.038216f
C901 VTAIL.n28 VSUBS 0.094262f
C902 VTAIL.n29 VSUBS 0.01712f
C903 VTAIL.n30 VSUBS 0.016169f
C904 VTAIL.n31 VSUBS 0.071605f
C905 VTAIL.n32 VSUBS 0.047543f
C906 VTAIL.n33 VSUBS 0.368286f
C907 VTAIL.n34 VSUBS 0.033573f
C908 VTAIL.n35 VSUBS 0.030089f
C909 VTAIL.n36 VSUBS 0.016169f
C910 VTAIL.n37 VSUBS 0.038216f
C911 VTAIL.n38 VSUBS 0.01712f
C912 VTAIL.n39 VSUBS 0.030089f
C913 VTAIL.n40 VSUBS 0.016169f
C914 VTAIL.n41 VSUBS 0.038216f
C915 VTAIL.n42 VSUBS 0.01712f
C916 VTAIL.n43 VSUBS 0.133563f
C917 VTAIL.t9 VSUBS 0.082088f
C918 VTAIL.n44 VSUBS 0.028662f
C919 VTAIL.n45 VSUBS 0.024299f
C920 VTAIL.n46 VSUBS 0.016169f
C921 VTAIL.n47 VSUBS 0.696889f
C922 VTAIL.n48 VSUBS 0.030089f
C923 VTAIL.n49 VSUBS 0.016169f
C924 VTAIL.n50 VSUBS 0.01712f
C925 VTAIL.n51 VSUBS 0.038216f
C926 VTAIL.n52 VSUBS 0.038216f
C927 VTAIL.n53 VSUBS 0.01712f
C928 VTAIL.n54 VSUBS 0.016169f
C929 VTAIL.n55 VSUBS 0.030089f
C930 VTAIL.n56 VSUBS 0.030089f
C931 VTAIL.n57 VSUBS 0.016169f
C932 VTAIL.n58 VSUBS 0.01712f
C933 VTAIL.n59 VSUBS 0.038216f
C934 VTAIL.n60 VSUBS 0.094262f
C935 VTAIL.n61 VSUBS 0.01712f
C936 VTAIL.n62 VSUBS 0.016169f
C937 VTAIL.n63 VSUBS 0.071605f
C938 VTAIL.n64 VSUBS 0.047543f
C939 VTAIL.n65 VSUBS 0.368286f
C940 VTAIL.t12 VSUBS 0.143852f
C941 VTAIL.t8 VSUBS 0.143852f
C942 VTAIL.n66 VSUBS 0.851384f
C943 VTAIL.n67 VSUBS 1.14481f
C944 VTAIL.n68 VSUBS 0.033573f
C945 VTAIL.n69 VSUBS 0.030089f
C946 VTAIL.n70 VSUBS 0.016169f
C947 VTAIL.n71 VSUBS 0.038216f
C948 VTAIL.n72 VSUBS 0.01712f
C949 VTAIL.n73 VSUBS 0.030089f
C950 VTAIL.n74 VSUBS 0.016169f
C951 VTAIL.n75 VSUBS 0.038216f
C952 VTAIL.n76 VSUBS 0.01712f
C953 VTAIL.n77 VSUBS 0.133563f
C954 VTAIL.t11 VSUBS 0.082088f
C955 VTAIL.n78 VSUBS 0.028662f
C956 VTAIL.n79 VSUBS 0.024299f
C957 VTAIL.n80 VSUBS 0.016169f
C958 VTAIL.n81 VSUBS 0.696889f
C959 VTAIL.n82 VSUBS 0.030089f
C960 VTAIL.n83 VSUBS 0.016169f
C961 VTAIL.n84 VSUBS 0.01712f
C962 VTAIL.n85 VSUBS 0.038216f
C963 VTAIL.n86 VSUBS 0.038216f
C964 VTAIL.n87 VSUBS 0.01712f
C965 VTAIL.n88 VSUBS 0.016169f
C966 VTAIL.n89 VSUBS 0.030089f
C967 VTAIL.n90 VSUBS 0.030089f
C968 VTAIL.n91 VSUBS 0.016169f
C969 VTAIL.n92 VSUBS 0.01712f
C970 VTAIL.n93 VSUBS 0.038216f
C971 VTAIL.n94 VSUBS 0.094262f
C972 VTAIL.n95 VSUBS 0.01712f
C973 VTAIL.n96 VSUBS 0.016169f
C974 VTAIL.n97 VSUBS 0.071605f
C975 VTAIL.n98 VSUBS 0.047543f
C976 VTAIL.n99 VSUBS 1.533f
C977 VTAIL.n100 VSUBS 0.033573f
C978 VTAIL.n101 VSUBS 0.030089f
C979 VTAIL.n102 VSUBS 0.016169f
C980 VTAIL.n103 VSUBS 0.038216f
C981 VTAIL.n104 VSUBS 0.01712f
C982 VTAIL.n105 VSUBS 0.030089f
C983 VTAIL.n106 VSUBS 0.016169f
C984 VTAIL.n107 VSUBS 0.038216f
C985 VTAIL.n108 VSUBS 0.01712f
C986 VTAIL.n109 VSUBS 0.133563f
C987 VTAIL.t2 VSUBS 0.082088f
C988 VTAIL.n110 VSUBS 0.028662f
C989 VTAIL.n111 VSUBS 0.024299f
C990 VTAIL.n112 VSUBS 0.016169f
C991 VTAIL.n113 VSUBS 0.696889f
C992 VTAIL.n114 VSUBS 0.030089f
C993 VTAIL.n115 VSUBS 0.016169f
C994 VTAIL.n116 VSUBS 0.01712f
C995 VTAIL.n117 VSUBS 0.038216f
C996 VTAIL.n118 VSUBS 0.038216f
C997 VTAIL.n119 VSUBS 0.01712f
C998 VTAIL.n120 VSUBS 0.016169f
C999 VTAIL.n121 VSUBS 0.030089f
C1000 VTAIL.n122 VSUBS 0.030089f
C1001 VTAIL.n123 VSUBS 0.016169f
C1002 VTAIL.n124 VSUBS 0.01712f
C1003 VTAIL.n125 VSUBS 0.038216f
C1004 VTAIL.n126 VSUBS 0.094262f
C1005 VTAIL.n127 VSUBS 0.01712f
C1006 VTAIL.n128 VSUBS 0.016169f
C1007 VTAIL.n129 VSUBS 0.071605f
C1008 VTAIL.n130 VSUBS 0.047543f
C1009 VTAIL.n131 VSUBS 1.533f
C1010 VTAIL.t4 VSUBS 0.143852f
C1011 VTAIL.t6 VSUBS 0.143852f
C1012 VTAIL.n132 VSUBS 0.85139f
C1013 VTAIL.n133 VSUBS 1.1448f
C1014 VTAIL.n134 VSUBS 0.033573f
C1015 VTAIL.n135 VSUBS 0.030089f
C1016 VTAIL.n136 VSUBS 0.016169f
C1017 VTAIL.n137 VSUBS 0.038216f
C1018 VTAIL.n138 VSUBS 0.01712f
C1019 VTAIL.n139 VSUBS 0.030089f
C1020 VTAIL.n140 VSUBS 0.016169f
C1021 VTAIL.n141 VSUBS 0.038216f
C1022 VTAIL.n142 VSUBS 0.01712f
C1023 VTAIL.n143 VSUBS 0.133563f
C1024 VTAIL.t7 VSUBS 0.082088f
C1025 VTAIL.n144 VSUBS 0.028662f
C1026 VTAIL.n145 VSUBS 0.024299f
C1027 VTAIL.n146 VSUBS 0.016169f
C1028 VTAIL.n147 VSUBS 0.696889f
C1029 VTAIL.n148 VSUBS 0.030089f
C1030 VTAIL.n149 VSUBS 0.016169f
C1031 VTAIL.n150 VSUBS 0.01712f
C1032 VTAIL.n151 VSUBS 0.038216f
C1033 VTAIL.n152 VSUBS 0.038216f
C1034 VTAIL.n153 VSUBS 0.01712f
C1035 VTAIL.n154 VSUBS 0.016169f
C1036 VTAIL.n155 VSUBS 0.030089f
C1037 VTAIL.n156 VSUBS 0.030089f
C1038 VTAIL.n157 VSUBS 0.016169f
C1039 VTAIL.n158 VSUBS 0.01712f
C1040 VTAIL.n159 VSUBS 0.038216f
C1041 VTAIL.n160 VSUBS 0.094262f
C1042 VTAIL.n161 VSUBS 0.01712f
C1043 VTAIL.n162 VSUBS 0.016169f
C1044 VTAIL.n163 VSUBS 0.071605f
C1045 VTAIL.n164 VSUBS 0.047543f
C1046 VTAIL.n165 VSUBS 0.368286f
C1047 VTAIL.n166 VSUBS 0.033573f
C1048 VTAIL.n167 VSUBS 0.030089f
C1049 VTAIL.n168 VSUBS 0.016169f
C1050 VTAIL.n169 VSUBS 0.038216f
C1051 VTAIL.n170 VSUBS 0.01712f
C1052 VTAIL.n171 VSUBS 0.030089f
C1053 VTAIL.n172 VSUBS 0.016169f
C1054 VTAIL.n173 VSUBS 0.038216f
C1055 VTAIL.n174 VSUBS 0.01712f
C1056 VTAIL.n175 VSUBS 0.133563f
C1057 VTAIL.t13 VSUBS 0.082088f
C1058 VTAIL.n176 VSUBS 0.028662f
C1059 VTAIL.n177 VSUBS 0.024299f
C1060 VTAIL.n178 VSUBS 0.016169f
C1061 VTAIL.n179 VSUBS 0.696889f
C1062 VTAIL.n180 VSUBS 0.030089f
C1063 VTAIL.n181 VSUBS 0.016169f
C1064 VTAIL.n182 VSUBS 0.01712f
C1065 VTAIL.n183 VSUBS 0.038216f
C1066 VTAIL.n184 VSUBS 0.038216f
C1067 VTAIL.n185 VSUBS 0.01712f
C1068 VTAIL.n186 VSUBS 0.016169f
C1069 VTAIL.n187 VSUBS 0.030089f
C1070 VTAIL.n188 VSUBS 0.030089f
C1071 VTAIL.n189 VSUBS 0.016169f
C1072 VTAIL.n190 VSUBS 0.01712f
C1073 VTAIL.n191 VSUBS 0.038216f
C1074 VTAIL.n192 VSUBS 0.094262f
C1075 VTAIL.n193 VSUBS 0.01712f
C1076 VTAIL.n194 VSUBS 0.016169f
C1077 VTAIL.n195 VSUBS 0.071605f
C1078 VTAIL.n196 VSUBS 0.047543f
C1079 VTAIL.n197 VSUBS 0.368286f
C1080 VTAIL.t14 VSUBS 0.143852f
C1081 VTAIL.t15 VSUBS 0.143852f
C1082 VTAIL.n198 VSUBS 0.85139f
C1083 VTAIL.n199 VSUBS 1.1448f
C1084 VTAIL.n200 VSUBS 0.033573f
C1085 VTAIL.n201 VSUBS 0.030089f
C1086 VTAIL.n202 VSUBS 0.016169f
C1087 VTAIL.n203 VSUBS 0.038216f
C1088 VTAIL.n204 VSUBS 0.01712f
C1089 VTAIL.n205 VSUBS 0.030089f
C1090 VTAIL.n206 VSUBS 0.016169f
C1091 VTAIL.n207 VSUBS 0.038216f
C1092 VTAIL.n208 VSUBS 0.01712f
C1093 VTAIL.n209 VSUBS 0.133563f
C1094 VTAIL.t10 VSUBS 0.082088f
C1095 VTAIL.n210 VSUBS 0.028662f
C1096 VTAIL.n211 VSUBS 0.024299f
C1097 VTAIL.n212 VSUBS 0.016169f
C1098 VTAIL.n213 VSUBS 0.696889f
C1099 VTAIL.n214 VSUBS 0.030089f
C1100 VTAIL.n215 VSUBS 0.016169f
C1101 VTAIL.n216 VSUBS 0.01712f
C1102 VTAIL.n217 VSUBS 0.038216f
C1103 VTAIL.n218 VSUBS 0.038216f
C1104 VTAIL.n219 VSUBS 0.01712f
C1105 VTAIL.n220 VSUBS 0.016169f
C1106 VTAIL.n221 VSUBS 0.030089f
C1107 VTAIL.n222 VSUBS 0.030089f
C1108 VTAIL.n223 VSUBS 0.016169f
C1109 VTAIL.n224 VSUBS 0.01712f
C1110 VTAIL.n225 VSUBS 0.038216f
C1111 VTAIL.n226 VSUBS 0.094262f
C1112 VTAIL.n227 VSUBS 0.01712f
C1113 VTAIL.n228 VSUBS 0.016169f
C1114 VTAIL.n229 VSUBS 0.071605f
C1115 VTAIL.n230 VSUBS 0.047543f
C1116 VTAIL.n231 VSUBS 1.533f
C1117 VTAIL.n232 VSUBS 0.033573f
C1118 VTAIL.n233 VSUBS 0.030089f
C1119 VTAIL.n234 VSUBS 0.016169f
C1120 VTAIL.n235 VSUBS 0.038216f
C1121 VTAIL.n236 VSUBS 0.01712f
C1122 VTAIL.n237 VSUBS 0.030089f
C1123 VTAIL.n238 VSUBS 0.016169f
C1124 VTAIL.n239 VSUBS 0.038216f
C1125 VTAIL.n240 VSUBS 0.01712f
C1126 VTAIL.n241 VSUBS 0.133563f
C1127 VTAIL.t1 VSUBS 0.082088f
C1128 VTAIL.n242 VSUBS 0.028662f
C1129 VTAIL.n243 VSUBS 0.024299f
C1130 VTAIL.n244 VSUBS 0.016169f
C1131 VTAIL.n245 VSUBS 0.696889f
C1132 VTAIL.n246 VSUBS 0.030089f
C1133 VTAIL.n247 VSUBS 0.016169f
C1134 VTAIL.n248 VSUBS 0.01712f
C1135 VTAIL.n249 VSUBS 0.038216f
C1136 VTAIL.n250 VSUBS 0.038216f
C1137 VTAIL.n251 VSUBS 0.01712f
C1138 VTAIL.n252 VSUBS 0.016169f
C1139 VTAIL.n253 VSUBS 0.030089f
C1140 VTAIL.n254 VSUBS 0.030089f
C1141 VTAIL.n255 VSUBS 0.016169f
C1142 VTAIL.n256 VSUBS 0.01712f
C1143 VTAIL.n257 VSUBS 0.038216f
C1144 VTAIL.n258 VSUBS 0.094262f
C1145 VTAIL.n259 VSUBS 0.01712f
C1146 VTAIL.n260 VSUBS 0.016169f
C1147 VTAIL.n261 VSUBS 0.071605f
C1148 VTAIL.n262 VSUBS 0.047543f
C1149 VTAIL.n263 VSUBS 1.52736f
C1150 VP.t5 VSUBS 1.9291f
C1151 VP.n0 VSUBS 0.86016f
C1152 VP.n1 VSUBS 0.037512f
C1153 VP.n2 VSUBS 0.031103f
C1154 VP.n3 VSUBS 0.037512f
C1155 VP.t3 VSUBS 1.9291f
C1156 VP.n4 VSUBS 0.715043f
C1157 VP.n5 VSUBS 0.037512f
C1158 VP.n6 VSUBS 0.030325f
C1159 VP.n7 VSUBS 0.037512f
C1160 VP.t2 VSUBS 1.9291f
C1161 VP.n8 VSUBS 0.715043f
C1162 VP.n9 VSUBS 0.037512f
C1163 VP.n10 VSUBS 0.031103f
C1164 VP.n11 VSUBS 0.037512f
C1165 VP.t7 VSUBS 1.9291f
C1166 VP.n12 VSUBS 0.86016f
C1167 VP.t4 VSUBS 1.9291f
C1168 VP.n13 VSUBS 0.86016f
C1169 VP.n14 VSUBS 0.037512f
C1170 VP.n15 VSUBS 0.031103f
C1171 VP.n16 VSUBS 0.037512f
C1172 VP.t1 VSUBS 1.9291f
C1173 VP.n17 VSUBS 0.715043f
C1174 VP.n18 VSUBS 0.037512f
C1175 VP.n19 VSUBS 0.030325f
C1176 VP.n20 VSUBS 0.037512f
C1177 VP.t0 VSUBS 1.9291f
C1178 VP.n21 VSUBS 0.839939f
C1179 VP.t6 VSUBS 2.3415f
C1180 VP.n22 VSUBS 0.800071f
C1181 VP.n23 VSUBS 0.436375f
C1182 VP.n24 VSUBS 0.054035f
C1183 VP.n25 VSUBS 0.069912f
C1184 VP.n26 VSUBS 0.074554f
C1185 VP.n27 VSUBS 0.037512f
C1186 VP.n28 VSUBS 0.037512f
C1187 VP.n29 VSUBS 0.037512f
C1188 VP.n30 VSUBS 0.074554f
C1189 VP.n31 VSUBS 0.069912f
C1190 VP.n32 VSUBS 0.054035f
C1191 VP.n33 VSUBS 0.037512f
C1192 VP.n34 VSUBS 0.037512f
C1193 VP.n35 VSUBS 0.051273f
C1194 VP.n36 VSUBS 0.069912f
C1195 VP.n37 VSUBS 0.075633f
C1196 VP.n38 VSUBS 0.037512f
C1197 VP.n39 VSUBS 0.037512f
C1198 VP.n40 VSUBS 0.037512f
C1199 VP.n41 VSUBS 0.072697f
C1200 VP.n42 VSUBS 0.069912f
C1201 VP.n43 VSUBS 0.056796f
C1202 VP.n44 VSUBS 0.060543f
C1203 VP.n45 VSUBS 2.09062f
C1204 VP.n46 VSUBS 2.11795f
C1205 VP.n47 VSUBS 0.060543f
C1206 VP.n48 VSUBS 0.056796f
C1207 VP.n49 VSUBS 0.069912f
C1208 VP.n50 VSUBS 0.072697f
C1209 VP.n51 VSUBS 0.037512f
C1210 VP.n52 VSUBS 0.037512f
C1211 VP.n53 VSUBS 0.037512f
C1212 VP.n54 VSUBS 0.075633f
C1213 VP.n55 VSUBS 0.069912f
C1214 VP.n56 VSUBS 0.051273f
C1215 VP.n57 VSUBS 0.037512f
C1216 VP.n58 VSUBS 0.037512f
C1217 VP.n59 VSUBS 0.054035f
C1218 VP.n60 VSUBS 0.069912f
C1219 VP.n61 VSUBS 0.074554f
C1220 VP.n62 VSUBS 0.037512f
C1221 VP.n63 VSUBS 0.037512f
C1222 VP.n64 VSUBS 0.037512f
C1223 VP.n65 VSUBS 0.074554f
C1224 VP.n66 VSUBS 0.069912f
C1225 VP.n67 VSUBS 0.054035f
C1226 VP.n68 VSUBS 0.037512f
C1227 VP.n69 VSUBS 0.037512f
C1228 VP.n70 VSUBS 0.051273f
C1229 VP.n71 VSUBS 0.069912f
C1230 VP.n72 VSUBS 0.075633f
C1231 VP.n73 VSUBS 0.037512f
C1232 VP.n74 VSUBS 0.037512f
C1233 VP.n75 VSUBS 0.037512f
C1234 VP.n76 VSUBS 0.072697f
C1235 VP.n77 VSUBS 0.069912f
C1236 VP.n78 VSUBS 0.056796f
C1237 VP.n79 VSUBS 0.060543f
C1238 VP.n80 VSUBS 0.088661f
.ends

