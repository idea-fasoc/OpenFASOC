* NGSPICE file created from opamp_sample_0001.ext - technology: sky130A

.subckt opamp_sample_0001 GND VOUT VDD VN VP CS_BIAS DIFFPAIR_BIAS
X0 GND.t129 GND.t127 GND.t128 GND.t12 sky130_fd_pr__nfet_01v8 ad=1.6263 pd=9.12 as=0 ps=0 w=4.17 l=2.04
X1 VDD.t174 a_n14320_7092.t8 VOUT.t5 VDD.t135 sky130_fd_pr__pfet_01v8 ad=0.9555 pd=5.68 as=0.40425 ps=2.78 w=2.45 l=5.22
X2 VDD.t1 a_n6573_8708.t22 a_n6651_8904.t7 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.8415 pd=5.43 as=1.989 ps=10.98 w=5.1 l=3.3
X3 VOUT.t48 a_n5180_7124.t0 sky130_fd_pr__cap_mim_m3_1 l=7.69 w=9.42
X4 a_n6651_8904.t17 a_n6573_8708.t2 a_n6573_8708.t3 VDD.t18 sky130_fd_pr__pfet_01v8 ad=0.8415 pd=5.43 as=1.989 ps=10.98 w=5.1 l=3.3
X5 GND.t126 GND.t124 GND.t125 GND.t32 sky130_fd_pr__nfet_01v8 ad=1.6263 pd=9.12 as=0 ps=0 w=4.17 l=2.04
X6 VN.t5 GND.t121 GND.t123 GND.t122 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X7 GND.t120 GND.t118 GND.t119 GND.t52 sky130_fd_pr__nfet_01v8 ad=1.6263 pd=9.12 as=0 ps=0 w=4.17 l=2.04
X8 a_n14320_7092.t1 a_n6573_8708.t23 a_n5180_7124.t18 VDD.t5 sky130_fd_pr__pfet_01v8 ad=0.8415 pd=5.43 as=0.8415 ps=5.43 w=5.1 l=3.3
X9 VOUT.t4 a_n14320_7092.t9 VDD.t173 VDD.t141 sky130_fd_pr__pfet_01v8 ad=0.40425 pd=2.78 as=0.9555 ps=5.68 w=2.45 l=5.22
X10 VDD.t172 a_n14320_7092.t10 VOUT.t35 VDD.t148 sky130_fd_pr__pfet_01v8 ad=0.40425 pd=2.78 as=0.40425 ps=2.78 w=2.45 l=5.22
X11 VDD.t8 a_n6573_8708.t24 a_n6651_8904.t6 VDD.t7 sky130_fd_pr__pfet_01v8 ad=0.8415 pd=5.43 as=0.8415 ps=5.43 w=5.1 l=3.3
X12 VOUT.t34 a_n14320_7092.t11 VDD.t171 VDD.t131 sky130_fd_pr__pfet_01v8 ad=0.40425 pd=2.78 as=0.9555 ps=5.68 w=2.45 l=5.22
X13 GND.t117 GND.t115 GND.t116 GND.t16 sky130_fd_pr__nfet_01v8 ad=1.6263 pd=9.12 as=0 ps=0 w=4.17 l=2.04
X14 a_n874_n120.t4 DIFFPAIR_BIAS.t6 a_n1379_n2440.t0 GND.t134 sky130_fd_pr__nfet_01v8 ad=1.5522 pd=8.74 as=1.5522 ps=8.74 w=3.98 l=2.27
X15 GND.t114 GND.t112 GND.t113 GND.t16 sky130_fd_pr__nfet_01v8 ad=1.6263 pd=9.12 as=0 ps=0 w=4.17 l=2.04
X16 VOUT.t47 CS_BIAS.t4 GND.t140 GND.t1 sky130_fd_pr__nfet_01v8 ad=1.6263 pd=9.12 as=1.6263 ps=9.12 w=4.17 l=2.04
X17 VOUT.t46 CS_BIAS.t5 GND.t139 GND.t130 sky130_fd_pr__nfet_01v8 ad=1.6263 pd=9.12 as=1.6263 ps=9.12 w=4.17 l=2.04
X18 VDD.t124 VDD.t122 VDD.t123 VDD.t113 sky130_fd_pr__pfet_01v8 ad=1.989 pd=10.98 as=0 ps=0 w=5.1 l=3.3
X19 a_n6651_8904.t5 a_n6573_8708.t25 VDD.t28 VDD.t27 sky130_fd_pr__pfet_01v8 ad=0.8415 pd=5.43 as=0.8415 ps=5.43 w=5.1 l=3.3
X20 GND.t111 GND.t109 GND.t110 GND.t52 sky130_fd_pr__nfet_01v8 ad=1.6263 pd=9.12 as=0 ps=0 w=4.17 l=2.04
X21 VDD.t170 a_n14320_7092.t12 VOUT.t33 VDD.t138 sky130_fd_pr__pfet_01v8 ad=0.40425 pd=2.78 as=0.40425 ps=2.78 w=2.45 l=5.22
X22 VDD.t121 VDD.t119 VDD.t120 VDD.t42 sky130_fd_pr__pfet_01v8 ad=0.9555 pd=5.68 as=0 ps=0 w=2.45 l=5.22
X23 VDD.t118 VDD.t116 VDD.t117 VDD.t81 sky130_fd_pr__pfet_01v8 ad=1.989 pd=10.98 as=0 ps=0 w=5.1 l=3.3
X24 VOUT.t9 a_n14320_7092.t13 VDD.t169 VDD.t143 sky130_fd_pr__pfet_01v8 ad=0.40425 pd=2.78 as=0.40425 ps=2.78 w=2.45 l=5.22
X25 VOUT.t8 a_n14320_7092.t14 VDD.t168 VDD.t143 sky130_fd_pr__pfet_01v8 ad=0.40425 pd=2.78 as=0.40425 ps=2.78 w=2.45 l=5.22
X26 a_n6573_8708.t13 a_n6573_8708.t12 a_n6651_8904.t16 VDD.t12 sky130_fd_pr__pfet_01v8 ad=0.8415 pd=5.43 as=0.8415 ps=5.43 w=5.1 l=3.3
X27 VN.t4 GND.t106 GND.t108 GND.t107 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X28 VP.t5 GND.t103 GND.t105 GND.t104 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X29 GND.t102 GND.t100 GND.t101 GND.t32 sky130_fd_pr__nfet_01v8 ad=1.6263 pd=9.12 as=0 ps=0 w=4.17 l=2.04
X30 a_n874_n120.t3 DIFFPAIR_BIAS.t7 a_n1379_n2440.t2 GND.t4 sky130_fd_pr__nfet_01v8 ad=1.5522 pd=8.74 as=1.5522 ps=8.74 w=3.98 l=2.27
X31 VOUT.t7 a_n14320_7092.t15 VDD.t167 VDD.t141 sky130_fd_pr__pfet_01v8 ad=0.40425 pd=2.78 as=0.9555 ps=5.68 w=2.45 l=5.22
X32 VDD.t166 a_n14320_7092.t16 VOUT.t15 VDD.t129 sky130_fd_pr__pfet_01v8 ad=0.9555 pd=5.68 as=0.40425 ps=2.78 w=2.45 l=5.22
X33 GND.t99 GND.t97 GND.t98 GND.t16 sky130_fd_pr__nfet_01v8 ad=1.6263 pd=9.12 as=0 ps=0 w=4.17 l=2.04
X34 a_n6651_8904.t4 a_n6573_8708.t26 VDD.t126 VDD.t125 sky130_fd_pr__pfet_01v8 ad=1.989 pd=10.98 as=0.8415 ps=5.43 w=5.1 l=3.3
X35 GND.t96 GND.t94 GND.t95 GND.t12 sky130_fd_pr__nfet_01v8 ad=1.6263 pd=9.12 as=0 ps=0 w=4.17 l=2.04
X36 a_n6651_8904.t15 a_n6573_8708.t8 a_n6573_8708.t9 VDD.t13 sky130_fd_pr__pfet_01v8 ad=0.8415 pd=5.43 as=0.8415 ps=5.43 w=5.1 l=3.3
X37 VDD.t165 a_n14320_7092.t17 VOUT.t14 VDD.t135 sky130_fd_pr__pfet_01v8 ad=0.9555 pd=5.68 as=0.40425 ps=2.78 w=2.45 l=5.22
X38 a_n6651_8904.t14 a_n6573_8708.t6 a_n6573_8708.t7 VDD.t4 sky130_fd_pr__pfet_01v8 ad=0.8415 pd=5.43 as=1.989 ps=10.98 w=5.1 l=3.3
X39 a_n6651_8904.t13 a_n6573_8708.t4 a_n6573_8708.t5 VDD.t20 sky130_fd_pr__pfet_01v8 ad=1.989 pd=10.98 as=0.8415 ps=5.43 w=5.1 l=3.3
X40 VDD.t179 a_n6573_8708.t27 a_n5180_7124.t8 VDD.t178 sky130_fd_pr__pfet_01v8 ad=0.8415 pd=5.43 as=1.989 ps=10.98 w=5.1 l=3.3
X41 VOUT.t45 CS_BIAS.t6 GND.t138 GND.t1 sky130_fd_pr__nfet_01v8 ad=1.6263 pd=9.12 as=1.6263 ps=9.12 w=4.17 l=2.04
X42 a_n6651_8904.t3 a_n6573_8708.t28 VDD.t32 VDD.t31 sky130_fd_pr__pfet_01v8 ad=0.8415 pd=5.43 as=0.8415 ps=5.43 w=5.1 l=3.3
X43 a_n14320_7092.t7 VN.t6 a_n874_n120.t6 GND.t133 sky130_fd_pr__nfet_01v8 ad=1.0647 pd=6.24 as=1.0647 ps=6.24 w=2.73 l=3.27
X44 VDD.t115 VDD.t112 VDD.t114 VDD.t113 sky130_fd_pr__pfet_01v8 ad=1.989 pd=10.98 as=0 ps=0 w=5.1 l=3.3
X45 VP.t4 GND.t91 GND.t93 GND.t92 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X46 VDD.t164 a_n14320_7092.t18 VOUT.t13 VDD.t148 sky130_fd_pr__pfet_01v8 ad=0.40425 pd=2.78 as=0.40425 ps=2.78 w=2.45 l=5.22
X47 VDD.t163 a_n14320_7092.t19 VOUT.t22 VDD.t138 sky130_fd_pr__pfet_01v8 ad=0.40425 pd=2.78 as=0.40425 ps=2.78 w=2.45 l=5.22
X48 VDD.t111 VDD.t109 VDD.t110 VDD.t42 sky130_fd_pr__pfet_01v8 ad=0.9555 pd=5.68 as=0 ps=0 w=2.45 l=5.22
X49 GND.t90 GND.t87 GND.t89 GND.t88 sky130_fd_pr__nfet_01v8 ad=1.5522 pd=8.74 as=0 ps=0 w=3.98 l=2.27
X50 VOUT.t0 CS_BIAS.t7 GND.t2 GND.t1 sky130_fd_pr__nfet_01v8 ad=1.6263 pd=9.12 as=1.6263 ps=9.12 w=4.17 l=2.04
X51 VP.t3 GND.t84 GND.t86 GND.t85 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X52 DIFFPAIR_BIAS.t3 DIFFPAIR_BIAS.t2 a_n2095_n2440.t2 GND.t0 sky130_fd_pr__nfet_01v8 ad=1.5522 pd=8.74 as=1.5522 ps=8.74 w=3.98 l=2.27
X53 a_n6651_8904.t12 a_n6573_8708.t18 a_n6573_8708.t19 VDD.t177 sky130_fd_pr__pfet_01v8 ad=1.989 pd=10.98 as=0.8415 ps=5.43 w=5.1 l=3.3
X54 a_n14320_7092.t0 a_n6573_8708.t29 a_n5180_7124.t17 VDD.t4 sky130_fd_pr__pfet_01v8 ad=0.8415 pd=5.43 as=1.989 ps=10.98 w=5.1 l=3.3
X55 VOUT.t49 a_n5180_7124.t0 sky130_fd_pr__cap_mim_m3_1 l=7.69 w=9.42
X56 VOUT.t21 a_n14320_7092.t20 VDD.t162 VDD.t127 sky130_fd_pr__pfet_01v8 ad=0.40425 pd=2.78 as=0.40425 ps=2.78 w=2.45 l=5.22
X57 GND.t83 GND.t81 GND.t82 GND.t52 sky130_fd_pr__nfet_01v8 ad=1.6263 pd=9.12 as=0 ps=0 w=4.17 l=2.04
X58 VDD.t161 a_n14320_7092.t21 VOUT.t20 VDD.t129 sky130_fd_pr__pfet_01v8 ad=0.9555 pd=5.68 as=0.40425 ps=2.78 w=2.45 l=5.22
X59 VDD.t108 VDD.t106 VDD.t107 VDD.t52 sky130_fd_pr__pfet_01v8 ad=0.9555 pd=5.68 as=0 ps=0 w=2.45 l=5.22
X60 GND.t80 GND.t78 GND.t79 GND.t32 sky130_fd_pr__nfet_01v8 ad=1.6263 pd=9.12 as=0 ps=0 w=4.17 l=2.04
X61 GND.t77 GND.t75 GND.t76 GND.t63 sky130_fd_pr__nfet_01v8 ad=1.0647 pd=6.24 as=0 ps=0 w=2.73 l=3.27
X62 VDD.t105 VDD.t103 VDD.t104 VDD.t34 sky130_fd_pr__pfet_01v8 ad=0.9555 pd=5.68 as=0 ps=0 w=2.45 l=5.22
X63 a_n14320_7092.t6 a_n6573_8708.t30 a_n5180_7124.t16 VDD.t177 sky130_fd_pr__pfet_01v8 ad=1.989 pd=10.98 as=0.8415 ps=5.43 w=5.1 l=3.3
X64 VDD.t102 VDD.t100 VDD.t101 VDD.t38 sky130_fd_pr__pfet_01v8 ad=0.9555 pd=5.68 as=0 ps=0 w=2.45 l=5.22
X65 GND.t74 GND.t72 GND.t73 GND.t56 sky130_fd_pr__nfet_01v8 ad=1.0647 pd=6.24 as=0 ps=0 w=2.73 l=3.27
X66 VOUT.t44 CS_BIAS.t8 GND.t137 GND.t130 sky130_fd_pr__nfet_01v8 ad=1.6263 pd=9.12 as=1.6263 ps=9.12 w=4.17 l=2.04
X67 VOUT.t28 a_n14320_7092.t22 VDD.t160 VDD.t141 sky130_fd_pr__pfet_01v8 ad=0.40425 pd=2.78 as=0.9555 ps=5.68 w=2.45 l=5.22
X68 VDD.t99 VDD.t97 VDD.t98 VDD.t42 sky130_fd_pr__pfet_01v8 ad=0.9555 pd=5.68 as=0 ps=0 w=2.45 l=5.22
X69 VDD.t96 VDD.t94 VDD.t95 VDD.t34 sky130_fd_pr__pfet_01v8 ad=0.9555 pd=5.68 as=0 ps=0 w=2.45 l=5.22
X70 a_n874_n120.t2 DIFFPAIR_BIAS.t8 a_n1379_n2440.t1 GND.t3 sky130_fd_pr__nfet_01v8 ad=1.5522 pd=8.74 as=1.5522 ps=8.74 w=3.98 l=2.27
X71 VDD.t93 VDD.t91 VDD.t92 VDD.t88 sky130_fd_pr__pfet_01v8 ad=1.989 pd=10.98 as=0 ps=0 w=5.1 l=3.3
X72 VDD.t90 VDD.t87 VDD.t89 VDD.t88 sky130_fd_pr__pfet_01v8 ad=1.989 pd=10.98 as=0 ps=0 w=5.1 l=3.3
X73 VOUT.t50 a_n5180_7124.t0 sky130_fd_pr__cap_mim_m3_1 l=7.69 w=9.42
X74 a_n6573_8708.t1 VP.t6 a_n874_n120.t1 GND.t7 sky130_fd_pr__nfet_01v8 ad=1.0647 pd=6.24 as=1.0647 ps=6.24 w=2.73 l=3.27
X75 a_n6573_8708.t0 VP.t7 a_n874_n120.t0 GND.t133 sky130_fd_pr__nfet_01v8 ad=1.0647 pd=6.24 as=1.0647 ps=6.24 w=2.73 l=3.27
X76 VOUT.t27 a_n14320_7092.t23 VDD.t159 VDD.t127 sky130_fd_pr__pfet_01v8 ad=0.40425 pd=2.78 as=0.40425 ps=2.78 w=2.45 l=5.22
X77 VDD.t86 VDD.t84 VDD.t85 VDD.t38 sky130_fd_pr__pfet_01v8 ad=0.9555 pd=5.68 as=0 ps=0 w=2.45 l=5.22
X78 CS_BIAS.t3 CS_BIAS.t2 GND.t6 GND.t1 sky130_fd_pr__nfet_01v8 ad=1.6263 pd=9.12 as=1.6263 ps=9.12 w=4.17 l=2.04
X79 a_n6651_8904.t11 a_n6573_8708.t16 a_n6573_8708.t17 VDD.t5 sky130_fd_pr__pfet_01v8 ad=0.8415 pd=5.43 as=0.8415 ps=5.43 w=5.1 l=3.3
X80 VDD.t83 VDD.t80 VDD.t82 VDD.t81 sky130_fd_pr__pfet_01v8 ad=1.989 pd=10.98 as=0 ps=0 w=5.1 l=3.3
X81 VDD.t158 a_n14320_7092.t24 VOUT.t26 VDD.t135 sky130_fd_pr__pfet_01v8 ad=0.9555 pd=5.68 as=0.40425 ps=2.78 w=2.45 l=5.22
X82 a_n6573_8708.t15 a_n6573_8708.t14 a_n6651_8904.t10 VDD.t9 sky130_fd_pr__pfet_01v8 ad=0.8415 pd=5.43 as=0.8415 ps=5.43 w=5.1 l=3.3
X83 VDD.t157 a_n14320_7092.t25 VOUT.t38 VDD.t148 sky130_fd_pr__pfet_01v8 ad=0.40425 pd=2.78 as=0.40425 ps=2.78 w=2.45 l=5.22
X84 GND.t71 GND.t69 VN.t3 GND.t70 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X85 VDD.t79 VDD.t77 VDD.t78 VDD.t52 sky130_fd_pr__pfet_01v8 ad=0.9555 pd=5.68 as=0 ps=0 w=2.45 l=5.22
X86 GND.t68 GND.t66 VP.t2 GND.t67 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X87 a_n6573_8708.t11 a_n6573_8708.t10 a_n6651_8904.t9 VDD.t19 sky130_fd_pr__pfet_01v8 ad=0.8415 pd=5.43 as=0.8415 ps=5.43 w=5.1 l=3.3
X88 VDD.t76 VDD.t74 VDD.t75 VDD.t34 sky130_fd_pr__pfet_01v8 ad=0.9555 pd=5.68 as=0 ps=0 w=2.45 l=5.22
X89 VDD.t17 a_n6573_8708.t31 a_n5180_7124.t7 VDD.t16 sky130_fd_pr__pfet_01v8 ad=0.8415 pd=5.43 as=1.989 ps=10.98 w=5.1 l=3.3
X90 VDD.t176 a_n6573_8708.t32 a_n5180_7124.t6 VDD.t175 sky130_fd_pr__pfet_01v8 ad=0.8415 pd=5.43 as=0.8415 ps=5.43 w=5.1 l=3.3
X91 DIFFPAIR_BIAS.t1 DIFFPAIR_BIAS.t0 a_n2095_n2440.t1 GND.t136 sky130_fd_pr__nfet_01v8 ad=1.5522 pd=8.74 as=1.5522 ps=8.74 w=3.98 l=2.27
X92 a_n14320_7092.t2 a_n6573_8708.t33 a_n5180_7124.t15 VDD.t13 sky130_fd_pr__pfet_01v8 ad=0.8415 pd=5.43 as=0.8415 ps=5.43 w=5.1 l=3.3
X93 GND.t65 GND.t62 GND.t64 GND.t63 sky130_fd_pr__nfet_01v8 ad=1.0647 pd=6.24 as=0 ps=0 w=2.73 l=3.27
X94 GND.t61 GND.t59 GND.t60 GND.t52 sky130_fd_pr__nfet_01v8 ad=1.6263 pd=9.12 as=0 ps=0 w=4.17 l=2.04
X95 a_n5180_7124.t14 a_n6573_8708.t34 a_n14320_7092.t1 VDD.t19 sky130_fd_pr__pfet_01v8 ad=0.8415 pd=5.43 as=0.8415 ps=5.43 w=5.1 l=3.3
X96 a_n14320_7092.t5 a_n6573_8708.t35 a_n5180_7124.t13 VDD.t20 sky130_fd_pr__pfet_01v8 ad=1.989 pd=10.98 as=0.8415 ps=5.43 w=5.1 l=3.3
X97 GND.t47 GND.t45 GND.t46 GND.t32 sky130_fd_pr__nfet_01v8 ad=1.6263 pd=9.12 as=0 ps=0 w=4.17 l=2.04
X98 GND.t58 GND.t55 GND.t57 GND.t56 sky130_fd_pr__nfet_01v8 ad=1.0647 pd=6.24 as=0 ps=0 w=2.73 l=3.27
X99 VOUT.t37 a_n14320_7092.t26 VDD.t156 VDD.t131 sky130_fd_pr__pfet_01v8 ad=0.40425 pd=2.78 as=0.9555 ps=5.68 w=2.45 l=5.22
X100 VOUT.t36 a_n14320_7092.t27 VDD.t155 VDD.t131 sky130_fd_pr__pfet_01v8 ad=0.40425 pd=2.78 as=0.9555 ps=5.68 w=2.45 l=5.22
X101 VDD.t154 a_n14320_7092.t28 VOUT.t12 VDD.t129 sky130_fd_pr__pfet_01v8 ad=0.9555 pd=5.68 as=0.40425 ps=2.78 w=2.45 l=5.22
X102 a_n6651_8904.t2 a_n6573_8708.t36 VDD.t15 VDD.t14 sky130_fd_pr__pfet_01v8 ad=1.989 pd=10.98 as=0.8415 ps=5.43 w=5.1 l=3.3
X103 a_n5180_7124.t5 a_n6573_8708.t37 VDD.t11 VDD.t10 sky130_fd_pr__pfet_01v8 ad=1.989 pd=10.98 as=0.8415 ps=5.43 w=5.1 l=3.3
X104 GND.t54 GND.t51 GND.t53 GND.t52 sky130_fd_pr__nfet_01v8 ad=1.6263 pd=9.12 as=0 ps=0 w=4.17 l=2.04
X105 VOUT.t11 a_n14320_7092.t29 VDD.t153 VDD.t143 sky130_fd_pr__pfet_01v8 ad=0.40425 pd=2.78 as=0.40425 ps=2.78 w=2.45 l=5.22
X106 VOUT.t51 a_n5180_7124.t0 sky130_fd_pr__cap_mim_m3_1 l=7.69 w=9.42
X107 GND.t50 GND.t48 VN.t2 GND.t49 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X108 VDD.t152 a_n14320_7092.t30 VOUT.t10 VDD.t148 sky130_fd_pr__pfet_01v8 ad=0.40425 pd=2.78 as=0.40425 ps=2.78 w=2.45 l=5.22
X109 a_6779_8904# a_6779_8904# a_6779_8904# VDD.t26 sky130_fd_pr__pfet_01v8 ad=1.989 pd=10.98 as=3.978 ps=21.96 w=5.1 l=3.3
X110 GND.t44 GND.t42 VP.t1 GND.t43 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X111 VOUT.t3 CS_BIAS.t9 GND.t135 GND.t1 sky130_fd_pr__nfet_01v8 ad=1.6263 pd=9.12 as=1.6263 ps=9.12 w=4.17 l=2.04
X112 GND.t41 GND.t38 GND.t40 GND.t39 sky130_fd_pr__nfet_01v8 ad=1.5522 pd=8.74 as=0 ps=0 w=3.98 l=2.27
X113 VOUT.t2 CS_BIAS.t10 GND.t132 GND.t130 sky130_fd_pr__nfet_01v8 ad=1.6263 pd=9.12 as=1.6263 ps=9.12 w=4.17 l=2.04
X114 a_n14320_7092.t4 VN.t7 a_n874_n120.t5 GND.t7 sky130_fd_pr__nfet_01v8 ad=1.0647 pd=6.24 as=1.0647 ps=6.24 w=2.73 l=3.27
X115 VDD.t151 a_n14320_7092.t31 VOUT.t18 VDD.t135 sky130_fd_pr__pfet_01v8 ad=0.9555 pd=5.68 as=0.40425 ps=2.78 w=2.45 l=5.22
X116 VDD.t30 a_n6573_8708.t38 a_n6651_8904.t1 VDD.t29 sky130_fd_pr__pfet_01v8 ad=0.8415 pd=5.43 as=0.8415 ps=5.43 w=5.1 l=3.3
X117 VOUT.t17 a_n14320_7092.t32 VDD.t150 VDD.t141 sky130_fd_pr__pfet_01v8 ad=0.40425 pd=2.78 as=0.9555 ps=5.68 w=2.45 l=5.22
X118 a_n5180_7124.t4 a_n6573_8708.t39 VDD.t183 VDD.t182 sky130_fd_pr__pfet_01v8 ad=1.989 pd=10.98 as=0.8415 ps=5.43 w=5.1 l=3.3
X119 GND.t37 GND.t35 VP.t0 GND.t36 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X120 VDD.t149 a_n14320_7092.t33 VOUT.t16 VDD.t148 sky130_fd_pr__pfet_01v8 ad=0.40425 pd=2.78 as=0.40425 ps=2.78 w=2.45 l=5.22
X121 VDD.t147 a_n14320_7092.t34 VOUT.t43 VDD.t138 sky130_fd_pr__pfet_01v8 ad=0.40425 pd=2.78 as=0.40425 ps=2.78 w=2.45 l=5.22
X122 GND.t34 GND.t31 GND.t33 GND.t32 sky130_fd_pr__nfet_01v8 ad=1.6263 pd=9.12 as=0 ps=0 w=4.17 l=2.04
X123 a_n7595_8904# a_n7595_8904# a_n7595_8904# VDD.t25 sky130_fd_pr__pfet_01v8 ad=1.989 pd=10.98 as=3.978 ps=21.96 w=5.1 l=3.3
X124 a_n5180_7124.t12 a_n6573_8708.t40 a_n14320_7092.t3 VDD.t6 sky130_fd_pr__pfet_01v8 ad=0.8415 pd=5.43 as=0.8415 ps=5.43 w=5.1 l=3.3
X125 GND.t30 GND.t28 GND.t29 GND.t16 sky130_fd_pr__nfet_01v8 ad=1.6263 pd=9.12 as=0 ps=0 w=4.17 l=2.04
X126 DIFFPAIR_BIAS.t5 DIFFPAIR_BIAS.t4 a_n2095_n2440.t0 GND.t5 sky130_fd_pr__nfet_01v8 ad=1.5522 pd=8.74 as=1.5522 ps=8.74 w=3.98 l=2.27
X127 GND.t27 GND.t25 GND.t26 GND.t12 sky130_fd_pr__nfet_01v8 ad=1.6263 pd=9.12 as=0 ps=0 w=4.17 l=2.04
X128 VOUT.t42 a_n14320_7092.t35 VDD.t146 VDD.t143 sky130_fd_pr__pfet_01v8 ad=0.40425 pd=2.78 as=0.40425 ps=2.78 w=2.45 l=5.22
X129 VDD.t73 VDD.t71 VDD.t72 VDD.t62 sky130_fd_pr__pfet_01v8 ad=1.989 pd=10.98 as=0 ps=0 w=5.1 l=3.3
X130 VDD.t145 a_n14320_7092.t36 VOUT.t30 VDD.t138 sky130_fd_pr__pfet_01v8 ad=0.40425 pd=2.78 as=0.40425 ps=2.78 w=2.45 l=5.22
X131 VDD.t70 VDD.t68 VDD.t69 VDD.t52 sky130_fd_pr__pfet_01v8 ad=0.9555 pd=5.68 as=0 ps=0 w=2.45 l=5.22
X132 VOUT.t52 a_n5180_7124.t0 sky130_fd_pr__cap_mim_m3_1 l=7.69 w=9.42
X133 GND.t24 GND.t22 VN.t1 GND.t23 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X134 VDD.t67 VDD.t65 VDD.t66 VDD.t42 sky130_fd_pr__pfet_01v8 ad=0.9555 pd=5.68 as=0 ps=0 w=2.45 l=5.22
X135 VOUT.t29 a_n14320_7092.t37 VDD.t144 VDD.t143 sky130_fd_pr__pfet_01v8 ad=0.40425 pd=2.78 as=0.40425 ps=2.78 w=2.45 l=5.22
X136 VOUT.t24 a_n14320_7092.t38 VDD.t142 VDD.t141 sky130_fd_pr__pfet_01v8 ad=0.40425 pd=2.78 as=0.9555 ps=5.68 w=2.45 l=5.22
X137 VOUT.t1 CS_BIAS.t11 GND.t131 GND.t130 sky130_fd_pr__nfet_01v8 ad=1.6263 pd=9.12 as=1.6263 ps=9.12 w=4.17 l=2.04
X138 a_n6573_8708.t21 a_n6573_8708.t20 a_n6651_8904.t8 VDD.t6 sky130_fd_pr__pfet_01v8 ad=0.8415 pd=5.43 as=0.8415 ps=5.43 w=5.1 l=3.3
X139 GND.t21 GND.t19 GND.t20 GND.t12 sky130_fd_pr__nfet_01v8 ad=1.6263 pd=9.12 as=0 ps=0 w=4.17 l=2.04
X140 VDD.t140 a_n14320_7092.t39 VOUT.t23 VDD.t129 sky130_fd_pr__pfet_01v8 ad=0.9555 pd=5.68 as=0.40425 ps=2.78 w=2.45 l=5.22
X141 a_n5180_7124.t11 a_n6573_8708.t41 a_n14320_7092.t0 VDD.t12 sky130_fd_pr__pfet_01v8 ad=0.8415 pd=5.43 as=0.8415 ps=5.43 w=5.1 l=3.3
X142 VDD.t24 a_n6573_8708.t42 a_n5180_7124.t3 VDD.t23 sky130_fd_pr__pfet_01v8 ad=0.8415 pd=5.43 as=0.8415 ps=5.43 w=5.1 l=3.3
X143 VDD.t64 VDD.t61 VDD.t63 VDD.t62 sky130_fd_pr__pfet_01v8 ad=1.989 pd=10.98 as=0 ps=0 w=5.1 l=3.3
X144 VDD.t139 a_n14320_7092.t40 VOUT.t19 VDD.t138 sky130_fd_pr__pfet_01v8 ad=0.40425 pd=2.78 as=0.40425 ps=2.78 w=2.45 l=5.22
X145 a_n5180_7124.t10 a_n6573_8708.t43 a_n14320_7092.t2 VDD.t9 sky130_fd_pr__pfet_01v8 ad=0.8415 pd=5.43 as=0.8415 ps=5.43 w=5.1 l=3.3
X146 VOUT.t40 a_n14320_7092.t41 VDD.t137 VDD.t127 sky130_fd_pr__pfet_01v8 ad=0.40425 pd=2.78 as=0.40425 ps=2.78 w=2.45 l=5.22
X147 VDD.t60 VDD.t58 VDD.t59 VDD.t38 sky130_fd_pr__pfet_01v8 ad=0.9555 pd=5.68 as=0 ps=0 w=2.45 l=5.22
X148 VDD.t136 a_n14320_7092.t42 VOUT.t39 VDD.t135 sky130_fd_pr__pfet_01v8 ad=0.9555 pd=5.68 as=0.40425 ps=2.78 w=2.45 l=5.22
X149 VDD.t57 VDD.t55 VDD.t56 VDD.t52 sky130_fd_pr__pfet_01v8 ad=0.9555 pd=5.68 as=0 ps=0 w=2.45 l=5.22
X150 VDD.t54 VDD.t51 VDD.t53 VDD.t52 sky130_fd_pr__pfet_01v8 ad=0.9555 pd=5.68 as=0 ps=0 w=2.45 l=5.22
X151 a_n5180_7124.t2 a_n6573_8708.t44 VDD.t3 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0.8415 pd=5.43 as=0.8415 ps=5.43 w=5.1 l=3.3
X152 GND.t18 GND.t15 GND.t17 GND.t16 sky130_fd_pr__nfet_01v8 ad=1.6263 pd=9.12 as=0 ps=0 w=4.17 l=2.04
X153 VDD.t181 a_n6573_8708.t45 a_n6651_8904.t0 VDD.t180 sky130_fd_pr__pfet_01v8 ad=0.8415 pd=5.43 as=1.989 ps=10.98 w=5.1 l=3.3
X154 GND.t14 GND.t11 GND.t13 GND.t12 sky130_fd_pr__nfet_01v8 ad=1.6263 pd=9.12 as=0 ps=0 w=4.17 l=2.04
X155 VN.t0 GND.t8 GND.t10 GND.t9 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X156 VOUT.t32 a_n14320_7092.t43 VDD.t134 VDD.t127 sky130_fd_pr__pfet_01v8 ad=0.40425 pd=2.78 as=0.40425 ps=2.78 w=2.45 l=5.22
X157 VOUT.t31 a_n14320_7092.t44 VDD.t133 VDD.t131 sky130_fd_pr__pfet_01v8 ad=0.40425 pd=2.78 as=0.9555 ps=5.68 w=2.45 l=5.22
X158 VDD.t50 VDD.t48 VDD.t49 VDD.t34 sky130_fd_pr__pfet_01v8 ad=0.9555 pd=5.68 as=0 ps=0 w=2.45 l=5.22
X159 VOUT.t6 a_n14320_7092.t45 VDD.t132 VDD.t131 sky130_fd_pr__pfet_01v8 ad=0.40425 pd=2.78 as=0.9555 ps=5.68 w=2.45 l=5.22
X160 VDD.t47 VDD.t45 VDD.t46 VDD.t38 sky130_fd_pr__pfet_01v8 ad=0.9555 pd=5.68 as=0 ps=0 w=2.45 l=5.22
X161 VDD.t130 a_n14320_7092.t46 VOUT.t25 VDD.t129 sky130_fd_pr__pfet_01v8 ad=0.9555 pd=5.68 as=0.40425 ps=2.78 w=2.45 l=5.22
X162 VOUT.t41 a_n14320_7092.t47 VDD.t128 VDD.t127 sky130_fd_pr__pfet_01v8 ad=0.40425 pd=2.78 as=0.40425 ps=2.78 w=2.45 l=5.22
X163 a_n14320_7092.t3 a_n6573_8708.t46 a_n5180_7124.t9 VDD.t18 sky130_fd_pr__pfet_01v8 ad=0.8415 pd=5.43 as=1.989 ps=10.98 w=5.1 l=3.3
X164 VDD.t44 VDD.t41 VDD.t43 VDD.t42 sky130_fd_pr__pfet_01v8 ad=0.9555 pd=5.68 as=0 ps=0 w=2.45 l=5.22
X165 VDD.t40 VDD.t37 VDD.t39 VDD.t38 sky130_fd_pr__pfet_01v8 ad=0.9555 pd=5.68 as=0 ps=0 w=2.45 l=5.22
X166 VDD.t36 VDD.t33 VDD.t35 VDD.t34 sky130_fd_pr__pfet_01v8 ad=0.9555 pd=5.68 as=0 ps=0 w=2.45 l=5.22
X167 a_n5180_7124.t1 a_n6573_8708.t47 VDD.t22 VDD.t21 sky130_fd_pr__pfet_01v8 ad=0.8415 pd=5.43 as=0.8415 ps=5.43 w=5.1 l=3.3
X168 VOUT.t53 a_n5180_7124.t0 sky130_fd_pr__cap_mim_m3_1 l=7.69 w=9.42
X169 CS_BIAS.t1 CS_BIAS.t0 GND.t141 GND.t130 sky130_fd_pr__nfet_01v8 ad=1.6263 pd=9.12 as=1.6263 ps=9.12 w=4.17 l=2.04
R0 GND.n5117 GND.n5116 2197.03
R1 GND.n4204 GND.n4203 1258.16
R2 GND.n3289 GND.n55 857.672
R3 GND.n3318 GND.n60 857.672
R4 GND.n3232 GND.n2147 857.672
R5 GND.n3400 GND.n2149 857.672
R6 GND.n2536 GND.n1360 857.672
R7 GND.n2755 GND.n1358 857.672
R8 GND.n1535 GND.n1415 857.672
R9 GND.n2846 GND.n1412 857.672
R10 GND.n257 GND.n50 833.646
R11 GND.n5475 GND.n59 833.646
R12 GND.n3403 GND.n3402 833.646
R13 GND.n3498 GND.n1979 833.646
R14 GND.n3949 GND.n1417 833.646
R15 GND.n3951 GND.n1410 833.646
R16 GND.n2722 GND.n1357 833.646
R17 GND.n3986 GND.n1361 833.646
R18 GND.n3546 GND.n1899 718.33
R19 GND.n3511 GND.n3510 718.33
R20 GND.n3852 GND.n1541 718.33
R21 GND.n3848 GND.n1554 718.33
R22 GND.n4313 GND.n1028 701.513
R23 GND.n5118 GND.n548 701.513
R24 GND.n5260 GND.n465 701.513
R25 GND.n4201 GND.n1139 701.513
R26 GND.n4313 GND.n4312 585
R27 GND.n4314 GND.n4313 585
R28 GND.n4311 GND.n1030 585
R29 GND.n1030 GND.n1029 585
R30 GND.n4310 GND.n4309 585
R31 GND.n4309 GND.n4308 585
R32 GND.n1035 GND.n1034 585
R33 GND.n4307 GND.n1035 585
R34 GND.n4305 GND.n4304 585
R35 GND.n4306 GND.n4305 585
R36 GND.n4303 GND.n1037 585
R37 GND.n1037 GND.n1036 585
R38 GND.n4302 GND.n4301 585
R39 GND.n4301 GND.n4300 585
R40 GND.n1043 GND.n1042 585
R41 GND.n4299 GND.n1043 585
R42 GND.n4297 GND.n4296 585
R43 GND.n4298 GND.n4297 585
R44 GND.n4295 GND.n1045 585
R45 GND.n1045 GND.n1044 585
R46 GND.n4294 GND.n4293 585
R47 GND.n4293 GND.n4292 585
R48 GND.n1051 GND.n1050 585
R49 GND.n4291 GND.n1051 585
R50 GND.n4289 GND.n4288 585
R51 GND.n4290 GND.n4289 585
R52 GND.n4287 GND.n1053 585
R53 GND.n1053 GND.n1052 585
R54 GND.n4286 GND.n4285 585
R55 GND.n4285 GND.n4284 585
R56 GND.n1059 GND.n1058 585
R57 GND.n4283 GND.n1059 585
R58 GND.n4281 GND.n4280 585
R59 GND.n4282 GND.n4281 585
R60 GND.n4279 GND.n1061 585
R61 GND.n1061 GND.n1060 585
R62 GND.n4278 GND.n4277 585
R63 GND.n4277 GND.n4276 585
R64 GND.n1067 GND.n1066 585
R65 GND.n4275 GND.n1067 585
R66 GND.n4273 GND.n4272 585
R67 GND.n4274 GND.n4273 585
R68 GND.n4271 GND.n1069 585
R69 GND.n1069 GND.n1068 585
R70 GND.n4270 GND.n4269 585
R71 GND.n4269 GND.n4268 585
R72 GND.n1075 GND.n1074 585
R73 GND.n4267 GND.n1075 585
R74 GND.n4265 GND.n4264 585
R75 GND.n4266 GND.n4265 585
R76 GND.n4263 GND.n1077 585
R77 GND.n1077 GND.n1076 585
R78 GND.n4262 GND.n4261 585
R79 GND.n4261 GND.n4260 585
R80 GND.n1083 GND.n1082 585
R81 GND.n4259 GND.n1083 585
R82 GND.n4257 GND.n4256 585
R83 GND.n4258 GND.n4257 585
R84 GND.n4255 GND.n1085 585
R85 GND.n1085 GND.n1084 585
R86 GND.n4254 GND.n4253 585
R87 GND.n4253 GND.n4252 585
R88 GND.n1091 GND.n1090 585
R89 GND.n4251 GND.n1091 585
R90 GND.n4249 GND.n4248 585
R91 GND.n4250 GND.n4249 585
R92 GND.n4247 GND.n1093 585
R93 GND.n1093 GND.n1092 585
R94 GND.n4246 GND.n4245 585
R95 GND.n4245 GND.n4244 585
R96 GND.n1099 GND.n1098 585
R97 GND.n4243 GND.n1099 585
R98 GND.n4241 GND.n4240 585
R99 GND.n4242 GND.n4241 585
R100 GND.n4239 GND.n1101 585
R101 GND.n1101 GND.n1100 585
R102 GND.n4238 GND.n4237 585
R103 GND.n4237 GND.n4236 585
R104 GND.n1107 GND.n1106 585
R105 GND.n4235 GND.n1107 585
R106 GND.n4233 GND.n4232 585
R107 GND.n4234 GND.n4233 585
R108 GND.n4231 GND.n1109 585
R109 GND.n1109 GND.n1108 585
R110 GND.n4230 GND.n4229 585
R111 GND.n4229 GND.n4228 585
R112 GND.n1115 GND.n1114 585
R113 GND.n4227 GND.n1115 585
R114 GND.n4225 GND.n4224 585
R115 GND.n4226 GND.n4225 585
R116 GND.n4223 GND.n1117 585
R117 GND.n1117 GND.n1116 585
R118 GND.n4222 GND.n4221 585
R119 GND.n4221 GND.n4220 585
R120 GND.n1123 GND.n1122 585
R121 GND.n4219 GND.n1123 585
R122 GND.n4217 GND.n4216 585
R123 GND.n4218 GND.n4217 585
R124 GND.n4215 GND.n1125 585
R125 GND.n1125 GND.n1124 585
R126 GND.n4214 GND.n4213 585
R127 GND.n4213 GND.n4212 585
R128 GND.n1131 GND.n1130 585
R129 GND.n4211 GND.n1131 585
R130 GND.n4209 GND.n4208 585
R131 GND.n4210 GND.n4209 585
R132 GND.n4207 GND.n1133 585
R133 GND.n1133 GND.n1132 585
R134 GND.n4206 GND.n4205 585
R135 GND.n4205 GND.n4204 585
R136 GND.n1028 GND.n1027 585
R137 GND.n4315 GND.n1028 585
R138 GND.n4318 GND.n4317 585
R139 GND.n4317 GND.n4316 585
R140 GND.n1025 GND.n1024 585
R141 GND.n1024 GND.n1023 585
R142 GND.n4323 GND.n4322 585
R143 GND.n4324 GND.n4323 585
R144 GND.n1022 GND.n1021 585
R145 GND.n4325 GND.n1022 585
R146 GND.n4328 GND.n4327 585
R147 GND.n4327 GND.n4326 585
R148 GND.n1019 GND.n1018 585
R149 GND.n1018 GND.n1017 585
R150 GND.n4333 GND.n4332 585
R151 GND.n4334 GND.n4333 585
R152 GND.n1016 GND.n1015 585
R153 GND.n4335 GND.n1016 585
R154 GND.n4338 GND.n4337 585
R155 GND.n4337 GND.n4336 585
R156 GND.n1013 GND.n1012 585
R157 GND.n1012 GND.n1011 585
R158 GND.n4343 GND.n4342 585
R159 GND.n4344 GND.n4343 585
R160 GND.n1010 GND.n1009 585
R161 GND.n4345 GND.n1010 585
R162 GND.n4348 GND.n4347 585
R163 GND.n4347 GND.n4346 585
R164 GND.n1007 GND.n1006 585
R165 GND.n1006 GND.n1005 585
R166 GND.n4353 GND.n4352 585
R167 GND.n4354 GND.n4353 585
R168 GND.n1004 GND.n1003 585
R169 GND.n4355 GND.n1004 585
R170 GND.n4358 GND.n4357 585
R171 GND.n4357 GND.n4356 585
R172 GND.n1001 GND.n1000 585
R173 GND.n1000 GND.n999 585
R174 GND.n4363 GND.n4362 585
R175 GND.n4364 GND.n4363 585
R176 GND.n998 GND.n997 585
R177 GND.n4365 GND.n998 585
R178 GND.n4368 GND.n4367 585
R179 GND.n4367 GND.n4366 585
R180 GND.n995 GND.n994 585
R181 GND.n994 GND.n993 585
R182 GND.n4373 GND.n4372 585
R183 GND.n4374 GND.n4373 585
R184 GND.n992 GND.n991 585
R185 GND.n4375 GND.n992 585
R186 GND.n4378 GND.n4377 585
R187 GND.n4377 GND.n4376 585
R188 GND.n989 GND.n988 585
R189 GND.n988 GND.n987 585
R190 GND.n4383 GND.n4382 585
R191 GND.n4384 GND.n4383 585
R192 GND.n986 GND.n985 585
R193 GND.n4385 GND.n986 585
R194 GND.n4388 GND.n4387 585
R195 GND.n4387 GND.n4386 585
R196 GND.n983 GND.n982 585
R197 GND.n982 GND.n981 585
R198 GND.n4393 GND.n4392 585
R199 GND.n4394 GND.n4393 585
R200 GND.n980 GND.n979 585
R201 GND.n4395 GND.n980 585
R202 GND.n4398 GND.n4397 585
R203 GND.n4397 GND.n4396 585
R204 GND.n977 GND.n976 585
R205 GND.n976 GND.n975 585
R206 GND.n4403 GND.n4402 585
R207 GND.n4404 GND.n4403 585
R208 GND.n974 GND.n973 585
R209 GND.n4405 GND.n974 585
R210 GND.n4408 GND.n4407 585
R211 GND.n4407 GND.n4406 585
R212 GND.n971 GND.n970 585
R213 GND.n970 GND.n969 585
R214 GND.n4413 GND.n4412 585
R215 GND.n4414 GND.n4413 585
R216 GND.n968 GND.n967 585
R217 GND.n4415 GND.n968 585
R218 GND.n4418 GND.n4417 585
R219 GND.n4417 GND.n4416 585
R220 GND.n965 GND.n964 585
R221 GND.n964 GND.n963 585
R222 GND.n4423 GND.n4422 585
R223 GND.n4424 GND.n4423 585
R224 GND.n962 GND.n961 585
R225 GND.n4425 GND.n962 585
R226 GND.n4428 GND.n4427 585
R227 GND.n4427 GND.n4426 585
R228 GND.n959 GND.n958 585
R229 GND.n958 GND.n957 585
R230 GND.n4433 GND.n4432 585
R231 GND.n4434 GND.n4433 585
R232 GND.n956 GND.n955 585
R233 GND.n4435 GND.n956 585
R234 GND.n4438 GND.n4437 585
R235 GND.n4437 GND.n4436 585
R236 GND.n953 GND.n952 585
R237 GND.n952 GND.n951 585
R238 GND.n4443 GND.n4442 585
R239 GND.n4444 GND.n4443 585
R240 GND.n950 GND.n949 585
R241 GND.n4445 GND.n950 585
R242 GND.n4448 GND.n4447 585
R243 GND.n4447 GND.n4446 585
R244 GND.n947 GND.n946 585
R245 GND.n946 GND.n945 585
R246 GND.n4453 GND.n4452 585
R247 GND.n4454 GND.n4453 585
R248 GND.n944 GND.n943 585
R249 GND.n4455 GND.n944 585
R250 GND.n4458 GND.n4457 585
R251 GND.n4457 GND.n4456 585
R252 GND.n941 GND.n940 585
R253 GND.n940 GND.n939 585
R254 GND.n4463 GND.n4462 585
R255 GND.n4464 GND.n4463 585
R256 GND.n938 GND.n937 585
R257 GND.n4465 GND.n938 585
R258 GND.n4468 GND.n4467 585
R259 GND.n4467 GND.n4466 585
R260 GND.n935 GND.n934 585
R261 GND.n934 GND.n933 585
R262 GND.n4473 GND.n4472 585
R263 GND.n4474 GND.n4473 585
R264 GND.n932 GND.n931 585
R265 GND.n4475 GND.n932 585
R266 GND.n4478 GND.n4477 585
R267 GND.n4477 GND.n4476 585
R268 GND.n929 GND.n928 585
R269 GND.n928 GND.n927 585
R270 GND.n4483 GND.n4482 585
R271 GND.n4484 GND.n4483 585
R272 GND.n926 GND.n925 585
R273 GND.n4485 GND.n926 585
R274 GND.n4488 GND.n4487 585
R275 GND.n4487 GND.n4486 585
R276 GND.n923 GND.n922 585
R277 GND.n922 GND.n921 585
R278 GND.n4493 GND.n4492 585
R279 GND.n4494 GND.n4493 585
R280 GND.n920 GND.n919 585
R281 GND.n4495 GND.n920 585
R282 GND.n4498 GND.n4497 585
R283 GND.n4497 GND.n4496 585
R284 GND.n917 GND.n916 585
R285 GND.n916 GND.n915 585
R286 GND.n4503 GND.n4502 585
R287 GND.n4504 GND.n4503 585
R288 GND.n914 GND.n913 585
R289 GND.n4505 GND.n914 585
R290 GND.n4508 GND.n4507 585
R291 GND.n4507 GND.n4506 585
R292 GND.n911 GND.n910 585
R293 GND.n910 GND.n909 585
R294 GND.n4513 GND.n4512 585
R295 GND.n4514 GND.n4513 585
R296 GND.n908 GND.n907 585
R297 GND.n4515 GND.n908 585
R298 GND.n4518 GND.n4517 585
R299 GND.n4517 GND.n4516 585
R300 GND.n905 GND.n904 585
R301 GND.n904 GND.n903 585
R302 GND.n4523 GND.n4522 585
R303 GND.n4524 GND.n4523 585
R304 GND.n902 GND.n901 585
R305 GND.n4525 GND.n902 585
R306 GND.n4528 GND.n4527 585
R307 GND.n4527 GND.n4526 585
R308 GND.n899 GND.n898 585
R309 GND.n898 GND.n897 585
R310 GND.n4533 GND.n4532 585
R311 GND.n4534 GND.n4533 585
R312 GND.n896 GND.n895 585
R313 GND.n4535 GND.n896 585
R314 GND.n4538 GND.n4537 585
R315 GND.n4537 GND.n4536 585
R316 GND.n893 GND.n892 585
R317 GND.n892 GND.n891 585
R318 GND.n4543 GND.n4542 585
R319 GND.n4544 GND.n4543 585
R320 GND.n890 GND.n889 585
R321 GND.n4545 GND.n890 585
R322 GND.n4548 GND.n4547 585
R323 GND.n4547 GND.n4546 585
R324 GND.n887 GND.n886 585
R325 GND.n886 GND.n885 585
R326 GND.n4553 GND.n4552 585
R327 GND.n4554 GND.n4553 585
R328 GND.n884 GND.n883 585
R329 GND.n4555 GND.n884 585
R330 GND.n4558 GND.n4557 585
R331 GND.n4557 GND.n4556 585
R332 GND.n881 GND.n880 585
R333 GND.n880 GND.n879 585
R334 GND.n4563 GND.n4562 585
R335 GND.n4564 GND.n4563 585
R336 GND.n878 GND.n877 585
R337 GND.n4565 GND.n878 585
R338 GND.n4568 GND.n4567 585
R339 GND.n4567 GND.n4566 585
R340 GND.n875 GND.n874 585
R341 GND.n874 GND.n873 585
R342 GND.n4573 GND.n4572 585
R343 GND.n4574 GND.n4573 585
R344 GND.n872 GND.n871 585
R345 GND.n4575 GND.n872 585
R346 GND.n4578 GND.n4577 585
R347 GND.n4577 GND.n4576 585
R348 GND.n869 GND.n868 585
R349 GND.n868 GND.n867 585
R350 GND.n4583 GND.n4582 585
R351 GND.n4584 GND.n4583 585
R352 GND.n866 GND.n865 585
R353 GND.n4585 GND.n866 585
R354 GND.n4588 GND.n4587 585
R355 GND.n4587 GND.n4586 585
R356 GND.n863 GND.n862 585
R357 GND.n862 GND.n861 585
R358 GND.n4593 GND.n4592 585
R359 GND.n4594 GND.n4593 585
R360 GND.n860 GND.n859 585
R361 GND.n4595 GND.n860 585
R362 GND.n4598 GND.n4597 585
R363 GND.n4597 GND.n4596 585
R364 GND.n857 GND.n856 585
R365 GND.n856 GND.n855 585
R366 GND.n4603 GND.n4602 585
R367 GND.n4604 GND.n4603 585
R368 GND.n854 GND.n853 585
R369 GND.n4605 GND.n854 585
R370 GND.n4608 GND.n4607 585
R371 GND.n4607 GND.n4606 585
R372 GND.n851 GND.n850 585
R373 GND.n850 GND.n849 585
R374 GND.n4613 GND.n4612 585
R375 GND.n4614 GND.n4613 585
R376 GND.n848 GND.n847 585
R377 GND.n4615 GND.n848 585
R378 GND.n4618 GND.n4617 585
R379 GND.n4617 GND.n4616 585
R380 GND.n845 GND.n844 585
R381 GND.n844 GND.n843 585
R382 GND.n4623 GND.n4622 585
R383 GND.n4624 GND.n4623 585
R384 GND.n842 GND.n841 585
R385 GND.n4625 GND.n842 585
R386 GND.n4628 GND.n4627 585
R387 GND.n4627 GND.n4626 585
R388 GND.n839 GND.n838 585
R389 GND.n838 GND.n837 585
R390 GND.n4633 GND.n4632 585
R391 GND.n4634 GND.n4633 585
R392 GND.n836 GND.n835 585
R393 GND.n4635 GND.n836 585
R394 GND.n4638 GND.n4637 585
R395 GND.n4637 GND.n4636 585
R396 GND.n833 GND.n832 585
R397 GND.n832 GND.n831 585
R398 GND.n4643 GND.n4642 585
R399 GND.n4644 GND.n4643 585
R400 GND.n830 GND.n829 585
R401 GND.n4645 GND.n830 585
R402 GND.n4648 GND.n4647 585
R403 GND.n4647 GND.n4646 585
R404 GND.n827 GND.n826 585
R405 GND.n826 GND.n825 585
R406 GND.n4653 GND.n4652 585
R407 GND.n4654 GND.n4653 585
R408 GND.n824 GND.n823 585
R409 GND.n4655 GND.n824 585
R410 GND.n4658 GND.n4657 585
R411 GND.n4657 GND.n4656 585
R412 GND.n821 GND.n820 585
R413 GND.n820 GND.n819 585
R414 GND.n4663 GND.n4662 585
R415 GND.n4664 GND.n4663 585
R416 GND.n818 GND.n817 585
R417 GND.n4665 GND.n818 585
R418 GND.n4668 GND.n4667 585
R419 GND.n4667 GND.n4666 585
R420 GND.n815 GND.n814 585
R421 GND.n814 GND.n813 585
R422 GND.n4673 GND.n4672 585
R423 GND.n4674 GND.n4673 585
R424 GND.n812 GND.n811 585
R425 GND.n4675 GND.n812 585
R426 GND.n4678 GND.n4677 585
R427 GND.n4677 GND.n4676 585
R428 GND.n809 GND.n808 585
R429 GND.n808 GND.n807 585
R430 GND.n4683 GND.n4682 585
R431 GND.n4684 GND.n4683 585
R432 GND.n806 GND.n805 585
R433 GND.n4685 GND.n806 585
R434 GND.n4688 GND.n4687 585
R435 GND.n4687 GND.n4686 585
R436 GND.n803 GND.n802 585
R437 GND.n802 GND.n801 585
R438 GND.n4693 GND.n4692 585
R439 GND.n4694 GND.n4693 585
R440 GND.n800 GND.n799 585
R441 GND.n4695 GND.n800 585
R442 GND.n4698 GND.n4697 585
R443 GND.n4697 GND.n4696 585
R444 GND.n797 GND.n796 585
R445 GND.n796 GND.n795 585
R446 GND.n4703 GND.n4702 585
R447 GND.n4704 GND.n4703 585
R448 GND.n794 GND.n793 585
R449 GND.n4705 GND.n794 585
R450 GND.n4708 GND.n4707 585
R451 GND.n4707 GND.n4706 585
R452 GND.n791 GND.n790 585
R453 GND.n790 GND.n789 585
R454 GND.n4713 GND.n4712 585
R455 GND.n4714 GND.n4713 585
R456 GND.n788 GND.n787 585
R457 GND.n4715 GND.n788 585
R458 GND.n4718 GND.n4717 585
R459 GND.n4717 GND.n4716 585
R460 GND.n785 GND.n784 585
R461 GND.n784 GND.n783 585
R462 GND.n4723 GND.n4722 585
R463 GND.n4724 GND.n4723 585
R464 GND.n782 GND.n781 585
R465 GND.n4725 GND.n782 585
R466 GND.n4728 GND.n4727 585
R467 GND.n4727 GND.n4726 585
R468 GND.n779 GND.n778 585
R469 GND.n778 GND.n777 585
R470 GND.n4733 GND.n4732 585
R471 GND.n4734 GND.n4733 585
R472 GND.n776 GND.n775 585
R473 GND.n4735 GND.n776 585
R474 GND.n4738 GND.n4737 585
R475 GND.n4737 GND.n4736 585
R476 GND.n773 GND.n772 585
R477 GND.n772 GND.n771 585
R478 GND.n4743 GND.n4742 585
R479 GND.n4744 GND.n4743 585
R480 GND.n770 GND.n769 585
R481 GND.n4745 GND.n770 585
R482 GND.n4748 GND.n4747 585
R483 GND.n4747 GND.n4746 585
R484 GND.n767 GND.n766 585
R485 GND.n766 GND.n765 585
R486 GND.n4753 GND.n4752 585
R487 GND.n4754 GND.n4753 585
R488 GND.n764 GND.n763 585
R489 GND.n4755 GND.n764 585
R490 GND.n4758 GND.n4757 585
R491 GND.n4757 GND.n4756 585
R492 GND.n761 GND.n760 585
R493 GND.n760 GND.n759 585
R494 GND.n4763 GND.n4762 585
R495 GND.n4764 GND.n4763 585
R496 GND.n758 GND.n757 585
R497 GND.n4765 GND.n758 585
R498 GND.n4768 GND.n4767 585
R499 GND.n4767 GND.n4766 585
R500 GND.n755 GND.n754 585
R501 GND.n754 GND.n753 585
R502 GND.n4773 GND.n4772 585
R503 GND.n4774 GND.n4773 585
R504 GND.n752 GND.n751 585
R505 GND.n4775 GND.n752 585
R506 GND.n4778 GND.n4777 585
R507 GND.n4777 GND.n4776 585
R508 GND.n749 GND.n748 585
R509 GND.n748 GND.n747 585
R510 GND.n4783 GND.n4782 585
R511 GND.n4784 GND.n4783 585
R512 GND.n746 GND.n745 585
R513 GND.n4785 GND.n746 585
R514 GND.n4788 GND.n4787 585
R515 GND.n4787 GND.n4786 585
R516 GND.n743 GND.n742 585
R517 GND.n742 GND.n741 585
R518 GND.n4793 GND.n4792 585
R519 GND.n4794 GND.n4793 585
R520 GND.n740 GND.n739 585
R521 GND.n4795 GND.n740 585
R522 GND.n4798 GND.n4797 585
R523 GND.n4797 GND.n4796 585
R524 GND.n737 GND.n736 585
R525 GND.n736 GND.n735 585
R526 GND.n4803 GND.n4802 585
R527 GND.n4804 GND.n4803 585
R528 GND.n734 GND.n733 585
R529 GND.n4805 GND.n734 585
R530 GND.n4808 GND.n4807 585
R531 GND.n4807 GND.n4806 585
R532 GND.n731 GND.n730 585
R533 GND.n730 GND.n729 585
R534 GND.n4813 GND.n4812 585
R535 GND.n4814 GND.n4813 585
R536 GND.n728 GND.n727 585
R537 GND.n4815 GND.n728 585
R538 GND.n4818 GND.n4817 585
R539 GND.n4817 GND.n4816 585
R540 GND.n725 GND.n724 585
R541 GND.n724 GND.n723 585
R542 GND.n4823 GND.n4822 585
R543 GND.n4824 GND.n4823 585
R544 GND.n722 GND.n721 585
R545 GND.n4825 GND.n722 585
R546 GND.n4828 GND.n4827 585
R547 GND.n4827 GND.n4826 585
R548 GND.n719 GND.n718 585
R549 GND.n718 GND.n717 585
R550 GND.n4833 GND.n4832 585
R551 GND.n4834 GND.n4833 585
R552 GND.n716 GND.n715 585
R553 GND.n4835 GND.n716 585
R554 GND.n4838 GND.n4837 585
R555 GND.n4837 GND.n4836 585
R556 GND.n713 GND.n712 585
R557 GND.n712 GND.n711 585
R558 GND.n4843 GND.n4842 585
R559 GND.n4844 GND.n4843 585
R560 GND.n710 GND.n709 585
R561 GND.n4845 GND.n710 585
R562 GND.n4848 GND.n4847 585
R563 GND.n4847 GND.n4846 585
R564 GND.n707 GND.n706 585
R565 GND.n706 GND.n705 585
R566 GND.n4853 GND.n4852 585
R567 GND.n4854 GND.n4853 585
R568 GND.n704 GND.n703 585
R569 GND.n4855 GND.n704 585
R570 GND.n4858 GND.n4857 585
R571 GND.n4857 GND.n4856 585
R572 GND.n701 GND.n700 585
R573 GND.n700 GND.n699 585
R574 GND.n4863 GND.n4862 585
R575 GND.n4864 GND.n4863 585
R576 GND.n698 GND.n697 585
R577 GND.n4865 GND.n698 585
R578 GND.n4868 GND.n4867 585
R579 GND.n4867 GND.n4866 585
R580 GND.n695 GND.n694 585
R581 GND.n694 GND.n693 585
R582 GND.n4873 GND.n4872 585
R583 GND.n4874 GND.n4873 585
R584 GND.n692 GND.n691 585
R585 GND.n4875 GND.n692 585
R586 GND.n4878 GND.n4877 585
R587 GND.n4877 GND.n4876 585
R588 GND.n689 GND.n688 585
R589 GND.n688 GND.n687 585
R590 GND.n4883 GND.n4882 585
R591 GND.n4884 GND.n4883 585
R592 GND.n686 GND.n685 585
R593 GND.n4885 GND.n686 585
R594 GND.n4888 GND.n4887 585
R595 GND.n4887 GND.n4886 585
R596 GND.n683 GND.n682 585
R597 GND.n682 GND.n681 585
R598 GND.n4893 GND.n4892 585
R599 GND.n4894 GND.n4893 585
R600 GND.n680 GND.n679 585
R601 GND.n4895 GND.n680 585
R602 GND.n4898 GND.n4897 585
R603 GND.n4897 GND.n4896 585
R604 GND.n677 GND.n676 585
R605 GND.n676 GND.n675 585
R606 GND.n4903 GND.n4902 585
R607 GND.n4904 GND.n4903 585
R608 GND.n674 GND.n673 585
R609 GND.n4905 GND.n674 585
R610 GND.n4908 GND.n4907 585
R611 GND.n4907 GND.n4906 585
R612 GND.n671 GND.n670 585
R613 GND.n670 GND.n669 585
R614 GND.n4913 GND.n4912 585
R615 GND.n4914 GND.n4913 585
R616 GND.n668 GND.n667 585
R617 GND.n4915 GND.n668 585
R618 GND.n4918 GND.n4917 585
R619 GND.n4917 GND.n4916 585
R620 GND.n665 GND.n664 585
R621 GND.n664 GND.n663 585
R622 GND.n4923 GND.n4922 585
R623 GND.n4924 GND.n4923 585
R624 GND.n662 GND.n661 585
R625 GND.n4925 GND.n662 585
R626 GND.n4928 GND.n4927 585
R627 GND.n4927 GND.n4926 585
R628 GND.n659 GND.n658 585
R629 GND.n658 GND.n657 585
R630 GND.n4933 GND.n4932 585
R631 GND.n4934 GND.n4933 585
R632 GND.n656 GND.n655 585
R633 GND.n4935 GND.n656 585
R634 GND.n4938 GND.n4937 585
R635 GND.n4937 GND.n4936 585
R636 GND.n653 GND.n652 585
R637 GND.n652 GND.n651 585
R638 GND.n4943 GND.n4942 585
R639 GND.n4944 GND.n4943 585
R640 GND.n650 GND.n649 585
R641 GND.n4945 GND.n650 585
R642 GND.n4948 GND.n4947 585
R643 GND.n4947 GND.n4946 585
R644 GND.n647 GND.n646 585
R645 GND.n646 GND.n645 585
R646 GND.n4953 GND.n4952 585
R647 GND.n4954 GND.n4953 585
R648 GND.n644 GND.n643 585
R649 GND.n4955 GND.n644 585
R650 GND.n4958 GND.n4957 585
R651 GND.n4957 GND.n4956 585
R652 GND.n641 GND.n640 585
R653 GND.n640 GND.n639 585
R654 GND.n4963 GND.n4962 585
R655 GND.n4964 GND.n4963 585
R656 GND.n638 GND.n637 585
R657 GND.n4965 GND.n638 585
R658 GND.n4968 GND.n4967 585
R659 GND.n4967 GND.n4966 585
R660 GND.n635 GND.n634 585
R661 GND.n634 GND.n633 585
R662 GND.n4973 GND.n4972 585
R663 GND.n4974 GND.n4973 585
R664 GND.n632 GND.n631 585
R665 GND.n4975 GND.n632 585
R666 GND.n4978 GND.n4977 585
R667 GND.n4977 GND.n4976 585
R668 GND.n629 GND.n628 585
R669 GND.n628 GND.n627 585
R670 GND.n4983 GND.n4982 585
R671 GND.n4984 GND.n4983 585
R672 GND.n626 GND.n625 585
R673 GND.n4985 GND.n626 585
R674 GND.n4988 GND.n4987 585
R675 GND.n4987 GND.n4986 585
R676 GND.n623 GND.n622 585
R677 GND.n622 GND.n621 585
R678 GND.n4993 GND.n4992 585
R679 GND.n4994 GND.n4993 585
R680 GND.n620 GND.n619 585
R681 GND.n4995 GND.n620 585
R682 GND.n4998 GND.n4997 585
R683 GND.n4997 GND.n4996 585
R684 GND.n617 GND.n616 585
R685 GND.n616 GND.n615 585
R686 GND.n5003 GND.n5002 585
R687 GND.n5004 GND.n5003 585
R688 GND.n614 GND.n613 585
R689 GND.n5005 GND.n614 585
R690 GND.n5008 GND.n5007 585
R691 GND.n5007 GND.n5006 585
R692 GND.n611 GND.n610 585
R693 GND.n610 GND.n609 585
R694 GND.n5013 GND.n5012 585
R695 GND.n5014 GND.n5013 585
R696 GND.n608 GND.n607 585
R697 GND.n5015 GND.n608 585
R698 GND.n5018 GND.n5017 585
R699 GND.n5017 GND.n5016 585
R700 GND.n605 GND.n604 585
R701 GND.n604 GND.n603 585
R702 GND.n5023 GND.n5022 585
R703 GND.n5024 GND.n5023 585
R704 GND.n602 GND.n601 585
R705 GND.n5025 GND.n602 585
R706 GND.n5028 GND.n5027 585
R707 GND.n5027 GND.n5026 585
R708 GND.n599 GND.n598 585
R709 GND.n598 GND.n597 585
R710 GND.n5033 GND.n5032 585
R711 GND.n5034 GND.n5033 585
R712 GND.n596 GND.n595 585
R713 GND.n5035 GND.n596 585
R714 GND.n5038 GND.n5037 585
R715 GND.n5037 GND.n5036 585
R716 GND.n593 GND.n592 585
R717 GND.n592 GND.n591 585
R718 GND.n5043 GND.n5042 585
R719 GND.n5044 GND.n5043 585
R720 GND.n590 GND.n589 585
R721 GND.n5045 GND.n590 585
R722 GND.n5048 GND.n5047 585
R723 GND.n5047 GND.n5046 585
R724 GND.n587 GND.n586 585
R725 GND.n586 GND.n585 585
R726 GND.n5053 GND.n5052 585
R727 GND.n5054 GND.n5053 585
R728 GND.n584 GND.n583 585
R729 GND.n5055 GND.n584 585
R730 GND.n5058 GND.n5057 585
R731 GND.n5057 GND.n5056 585
R732 GND.n581 GND.n580 585
R733 GND.n580 GND.n579 585
R734 GND.n5063 GND.n5062 585
R735 GND.n5064 GND.n5063 585
R736 GND.n578 GND.n577 585
R737 GND.n5065 GND.n578 585
R738 GND.n5068 GND.n5067 585
R739 GND.n5067 GND.n5066 585
R740 GND.n575 GND.n574 585
R741 GND.n574 GND.n573 585
R742 GND.n5073 GND.n5072 585
R743 GND.n5074 GND.n5073 585
R744 GND.n572 GND.n571 585
R745 GND.n5075 GND.n572 585
R746 GND.n5078 GND.n5077 585
R747 GND.n5077 GND.n5076 585
R748 GND.n569 GND.n568 585
R749 GND.n568 GND.n567 585
R750 GND.n5083 GND.n5082 585
R751 GND.n5084 GND.n5083 585
R752 GND.n566 GND.n565 585
R753 GND.n5085 GND.n566 585
R754 GND.n5088 GND.n5087 585
R755 GND.n5087 GND.n5086 585
R756 GND.n563 GND.n562 585
R757 GND.n562 GND.n561 585
R758 GND.n5093 GND.n5092 585
R759 GND.n5094 GND.n5093 585
R760 GND.n560 GND.n559 585
R761 GND.n5095 GND.n560 585
R762 GND.n5098 GND.n5097 585
R763 GND.n5097 GND.n5096 585
R764 GND.n557 GND.n556 585
R765 GND.n556 GND.n555 585
R766 GND.n5103 GND.n5102 585
R767 GND.n5104 GND.n5103 585
R768 GND.n554 GND.n553 585
R769 GND.n5105 GND.n554 585
R770 GND.n5108 GND.n5107 585
R771 GND.n5107 GND.n5106 585
R772 GND.n551 GND.n550 585
R773 GND.n550 GND.n549 585
R774 GND.n5114 GND.n5113 585
R775 GND.n5115 GND.n5114 585
R776 GND.n5112 GND.n548 585
R777 GND.n5116 GND.n548 585
R778 GND.n5256 GND.n5255 585
R779 GND.n5257 GND.n5256 585
R780 GND.n468 GND.n467 585
R781 GND.n467 GND.n466 585
R782 GND.n5249 GND.n5248 585
R783 GND.n5248 GND.n5247 585
R784 GND.n471 GND.n470 585
R785 GND.n5246 GND.n471 585
R786 GND.n5244 GND.n5243 585
R787 GND.n5245 GND.n5244 585
R788 GND.n474 GND.n473 585
R789 GND.n473 GND.n472 585
R790 GND.n5239 GND.n5238 585
R791 GND.n5238 GND.n5237 585
R792 GND.n477 GND.n476 585
R793 GND.n5236 GND.n477 585
R794 GND.n5234 GND.n5233 585
R795 GND.n5235 GND.n5234 585
R796 GND.n480 GND.n479 585
R797 GND.n479 GND.n478 585
R798 GND.n5229 GND.n5228 585
R799 GND.n5228 GND.n5227 585
R800 GND.n483 GND.n482 585
R801 GND.n5226 GND.n483 585
R802 GND.n5224 GND.n5223 585
R803 GND.n5225 GND.n5224 585
R804 GND.n486 GND.n485 585
R805 GND.n485 GND.n484 585
R806 GND.n5219 GND.n5218 585
R807 GND.n5218 GND.n5217 585
R808 GND.n489 GND.n488 585
R809 GND.n5216 GND.n489 585
R810 GND.n5214 GND.n5213 585
R811 GND.n5215 GND.n5214 585
R812 GND.n492 GND.n491 585
R813 GND.n491 GND.n490 585
R814 GND.n5209 GND.n5208 585
R815 GND.n5208 GND.n5207 585
R816 GND.n495 GND.n494 585
R817 GND.n5206 GND.n495 585
R818 GND.n5204 GND.n5203 585
R819 GND.n5205 GND.n5204 585
R820 GND.n498 GND.n497 585
R821 GND.n497 GND.n496 585
R822 GND.n5199 GND.n5198 585
R823 GND.n5198 GND.n5197 585
R824 GND.n501 GND.n500 585
R825 GND.n5196 GND.n501 585
R826 GND.n5194 GND.n5193 585
R827 GND.n5195 GND.n5194 585
R828 GND.n504 GND.n503 585
R829 GND.n503 GND.n502 585
R830 GND.n5189 GND.n5188 585
R831 GND.n5188 GND.n5187 585
R832 GND.n507 GND.n506 585
R833 GND.n5186 GND.n507 585
R834 GND.n5184 GND.n5183 585
R835 GND.n5185 GND.n5184 585
R836 GND.n510 GND.n509 585
R837 GND.n509 GND.n508 585
R838 GND.n5179 GND.n5178 585
R839 GND.n5178 GND.n5177 585
R840 GND.n513 GND.n512 585
R841 GND.n5176 GND.n513 585
R842 GND.n5174 GND.n5173 585
R843 GND.n5175 GND.n5174 585
R844 GND.n516 GND.n515 585
R845 GND.n515 GND.n514 585
R846 GND.n5169 GND.n5168 585
R847 GND.n5168 GND.n5167 585
R848 GND.n519 GND.n518 585
R849 GND.n5166 GND.n519 585
R850 GND.n5164 GND.n5163 585
R851 GND.n5165 GND.n5164 585
R852 GND.n522 GND.n521 585
R853 GND.n521 GND.n520 585
R854 GND.n5159 GND.n5158 585
R855 GND.n5158 GND.n5157 585
R856 GND.n525 GND.n524 585
R857 GND.n5156 GND.n525 585
R858 GND.n5154 GND.n5153 585
R859 GND.n5155 GND.n5154 585
R860 GND.n528 GND.n527 585
R861 GND.n527 GND.n526 585
R862 GND.n5149 GND.n5148 585
R863 GND.n5148 GND.n5147 585
R864 GND.n531 GND.n530 585
R865 GND.n5146 GND.n531 585
R866 GND.n5144 GND.n5143 585
R867 GND.n5145 GND.n5144 585
R868 GND.n534 GND.n533 585
R869 GND.n533 GND.n532 585
R870 GND.n5139 GND.n5138 585
R871 GND.n5138 GND.n5137 585
R872 GND.n537 GND.n536 585
R873 GND.n5136 GND.n537 585
R874 GND.n5134 GND.n5133 585
R875 GND.n5135 GND.n5134 585
R876 GND.n540 GND.n539 585
R877 GND.n539 GND.n538 585
R878 GND.n5129 GND.n5128 585
R879 GND.n5128 GND.n5127 585
R880 GND.n543 GND.n542 585
R881 GND.n5126 GND.n543 585
R882 GND.n5124 GND.n5123 585
R883 GND.n5125 GND.n5124 585
R884 GND.n546 GND.n545 585
R885 GND.n545 GND.n544 585
R886 GND.n5119 GND.n5118 585
R887 GND.n5118 GND.n5117 585
R888 GND.n5478 GND.n55 585
R889 GND.n5474 GND.n55 585
R890 GND.n5480 GND.n5479 585
R891 GND.n5481 GND.n5480 585
R892 GND.n40 GND.n39 585
R893 GND.n3326 GND.n40 585
R894 GND.n5489 GND.n5488 585
R895 GND.n5488 GND.n5487 585
R896 GND.n5490 GND.n34 585
R897 GND.n3332 GND.n34 585
R898 GND.n5492 GND.n5491 585
R899 GND.n5493 GND.n5492 585
R900 GND.n35 GND.n33 585
R901 GND.n3338 GND.n33 585
R902 GND.n2229 GND.n2228 585
R903 GND.n2233 GND.n2229 585
R904 GND.n3364 GND.n3363 585
R905 GND.n3363 GND.n3362 585
R906 GND.n3365 GND.n13 585
R907 GND.n5500 GND.n13 585
R908 GND.n3367 GND.n3366 585
R909 GND.n3368 GND.n3367 585
R910 GND.n2224 GND.n2223 585
R911 GND.n2223 GND.n2191 585
R912 GND.n2182 GND.n2181 585
R913 GND.n3377 GND.n2182 585
R914 GND.n3383 GND.n3382 585
R915 GND.n3382 GND.n3381 585
R916 GND.n3384 GND.n2175 585
R917 GND.n3254 GND.n2175 585
R918 GND.n3386 GND.n3385 585
R919 GND.n3387 GND.n3386 585
R920 GND.n2176 GND.n2174 585
R921 GND.n3239 GND.n2174 585
R922 GND.n2159 GND.n2152 585
R923 GND.n3393 GND.n2159 585
R924 GND.n3398 GND.n2150 585
R925 GND.n2246 GND.n2150 585
R926 GND.n3400 GND.n3399 585
R927 GND.n3401 GND.n3400 585
R928 GND.n3203 GND.n2149 585
R929 GND.n3207 GND.n3205 585
R930 GND.n3209 GND.n3208 585
R931 GND.n3212 GND.n3211 585
R932 GND.n3210 GND.n2253 585
R933 GND.n3218 GND.n3217 585
R934 GND.n3220 GND.n3219 585
R935 GND.n3223 GND.n3222 585
R936 GND.n3221 GND.n2251 585
R937 GND.n3228 GND.n3227 585
R938 GND.n3230 GND.n3229 585
R939 GND.n3233 GND.n3232 585
R940 GND.n3319 GND.n3318 585
R941 GND.n3316 GND.n3315 585
R942 GND.n3314 GND.n3280 585
R943 GND.n3308 GND.n3281 585
R944 GND.n3310 GND.n3309 585
R945 GND.n3305 GND.n3283 585
R946 GND.n3304 GND.n3303 585
R947 GND.n3297 GND.n3285 585
R948 GND.n3299 GND.n3298 585
R949 GND.n3295 GND.n3287 585
R950 GND.n3294 GND.n3293 585
R951 GND.n3290 GND.n3289 585
R952 GND.n3322 GND.n60 585
R953 GND.n5474 GND.n60 585
R954 GND.n3323 GND.n53 585
R955 GND.n5481 GND.n53 585
R956 GND.n3325 GND.n3324 585
R957 GND.n3326 GND.n3325 585
R958 GND.n2241 GND.n43 585
R959 GND.n5487 GND.n43 585
R960 GND.n3334 GND.n3333 585
R961 GND.n3333 GND.n3332 585
R962 GND.n3335 GND.n31 585
R963 GND.n5493 GND.n31 585
R964 GND.n3337 GND.n3336 585
R965 GND.n3338 GND.n3337 585
R966 GND.n2236 GND.n2235 585
R967 GND.n2235 GND.n2233 585
R968 GND.n10 GND.n8 585
R969 GND.n3362 GND.n10 585
R970 GND.n5502 GND.n5501 585
R971 GND.n5501 GND.n5500 585
R972 GND.n9 GND.n7 585
R973 GND.n3368 GND.n9 585
R974 GND.n3249 GND.n3248 585
R975 GND.n3248 GND.n2191 585
R976 GND.n3250 GND.n2190 585
R977 GND.n3377 GND.n2190 585
R978 GND.n3251 GND.n2185 585
R979 GND.n3381 GND.n2185 585
R980 GND.n3253 GND.n3252 585
R981 GND.n3254 GND.n3253 585
R982 GND.n2243 GND.n2172 585
R983 GND.n3387 GND.n2172 585
R984 GND.n3241 GND.n3240 585
R985 GND.n3240 GND.n3239 585
R986 GND.n3238 GND.n2157 585
R987 GND.n3393 GND.n2157 585
R988 GND.n3237 GND.n2247 585
R989 GND.n2247 GND.n2246 585
R990 GND.n2245 GND.n2147 585
R991 GND.n3401 GND.n2147 585
R992 GND.n3550 GND.n1899 585
R993 GND.n3509 GND.n1899 585
R994 GND.n3552 GND.n3551 585
R995 GND.n3553 GND.n3552 585
R996 GND.n1900 GND.n1898 585
R997 GND.n1898 GND.n1895 585
R998 GND.n1882 GND.n1881 585
R999 GND.n3195 GND.n1882 585
R1000 GND.n3563 GND.n3562 585
R1001 GND.n3562 GND.n3561 585
R1002 GND.n3564 GND.n1876 585
R1003 GND.n3187 GND.n1876 585
R1004 GND.n3566 GND.n3565 585
R1005 GND.n3567 GND.n3566 585
R1006 GND.n1877 GND.n1875 585
R1007 GND.n1875 GND.n1872 585
R1008 GND.n3178 GND.n3162 585
R1009 GND.n3162 GND.n1861 585
R1010 GND.n3180 GND.n3179 585
R1011 GND.n3181 GND.n3180 585
R1012 GND.n3163 GND.n3161 585
R1013 GND.n3161 GND.n1829 585
R1014 GND.n3172 GND.n3171 585
R1015 GND.n3171 GND.n1822 585
R1016 GND.n3170 GND.n3165 585
R1017 GND.n3170 GND.n1820 585
R1018 GND.n3169 GND.n3168 585
R1019 GND.n3169 GND.n1806 585
R1020 GND.n1796 GND.n1795 585
R1021 GND.n3134 GND.n1796 585
R1022 GND.n3603 GND.n3602 585
R1023 GND.n3602 GND.n3601 585
R1024 GND.n3604 GND.n1790 585
R1025 GND.n3142 GND.n1790 585
R1026 GND.n3606 GND.n3605 585
R1027 GND.n3607 GND.n3606 585
R1028 GND.n1791 GND.n1789 585
R1029 GND.n3111 GND.n1789 585
R1030 GND.n3094 GND.n3093 585
R1031 GND.n3094 GND.n1778 585
R1032 GND.n3096 GND.n3095 585
R1033 GND.n3095 GND.n1776 585
R1034 GND.n3097 GND.n2287 585
R1035 GND.n2287 GND.n1770 585
R1036 GND.n3099 GND.n3098 585
R1037 GND.n3100 GND.n3099 585
R1038 GND.n2288 GND.n2286 585
R1039 GND.n2286 GND.n2285 585
R1040 GND.n3085 GND.n3084 585
R1041 GND.n3084 GND.n3083 585
R1042 GND.n2291 GND.n2290 585
R1043 GND.n2291 GND.n1753 585
R1044 GND.n3071 GND.n3070 585
R1045 GND.n3072 GND.n3071 585
R1046 GND.n2305 GND.n2304 585
R1047 GND.n2304 GND.n2303 585
R1048 GND.n3066 GND.n3065 585
R1049 GND.n3065 GND.n1741 585
R1050 GND.n3064 GND.n2307 585
R1051 GND.n3064 GND.n1735 585
R1052 GND.n3063 GND.n2309 585
R1053 GND.n3063 GND.n3062 585
R1054 GND.n3044 GND.n2308 585
R1055 GND.n3016 GND.n2308 585
R1056 GND.n3045 GND.n2320 585
R1057 GND.n2320 GND.n1723 585
R1058 GND.n3047 GND.n3046 585
R1059 GND.n3048 GND.n3047 585
R1060 GND.n2321 GND.n2319 585
R1061 GND.n3030 GND.n2319 585
R1062 GND.n3037 GND.n3036 585
R1063 GND.n3036 GND.n3035 585
R1064 GND.n2331 GND.n2323 585
R1065 GND.n2331 GND.n1706 585
R1066 GND.n2330 GND.n2329 585
R1067 GND.n2330 GND.n1700 585
R1068 GND.n2325 GND.n2324 585
R1069 GND.n2324 GND.n1698 585
R1070 GND.n1681 GND.n1680 585
R1071 GND.n2337 GND.n1681 585
R1072 GND.n3687 GND.n3686 585
R1073 GND.n3686 GND.n3685 585
R1074 GND.n3688 GND.n1675 585
R1075 GND.n2340 GND.n1675 585
R1076 GND.n3690 GND.n3689 585
R1077 GND.n3691 GND.n3690 585
R1078 GND.n1676 GND.n1674 585
R1079 GND.n1674 GND.n1664 585
R1080 GND.n2949 GND.n2948 585
R1081 GND.n2950 GND.n2949 585
R1082 GND.n1650 GND.n1649 585
R1083 GND.n2903 GND.n1650 585
R1084 GND.n3708 GND.n3707 585
R1085 GND.n3707 GND.n3706 585
R1086 GND.n3709 GND.n1644 585
R1087 GND.t70 GND.n1644 585
R1088 GND.n3711 GND.n3710 585
R1089 GND.n3712 GND.n3711 585
R1090 GND.n1584 GND.n1583 585
R1091 GND.n2351 GND.n1584 585
R1092 GND.n3793 GND.n3792 585
R1093 GND.n3792 GND.n3791 585
R1094 GND.n3794 GND.n1576 585
R1095 GND.n2870 GND.n1576 585
R1096 GND.n3796 GND.n3795 585
R1097 GND.n3797 GND.n3796 585
R1098 GND.n1577 GND.n1575 585
R1099 GND.n1575 GND.n1572 585
R1100 GND.n1559 GND.n1558 585
R1101 GND.n1562 GND.n1559 585
R1102 GND.n3807 GND.n3806 585
R1103 GND.n3806 GND.n3805 585
R1104 GND.n3808 GND.n1556 585
R1105 GND.n2473 GND.n1556 585
R1106 GND.n3809 GND.n1554 585
R1107 GND.n2475 GND.n1554 585
R1108 GND.n3848 GND.n3847 585
R1109 GND.n3846 GND.n1553 585
R1110 GND.n3845 GND.n1552 585
R1111 GND.n3850 GND.n1552 585
R1112 GND.n3844 GND.n3843 585
R1113 GND.n3842 GND.n3841 585
R1114 GND.n3840 GND.n3839 585
R1115 GND.n3838 GND.n3837 585
R1116 GND.n3836 GND.n3835 585
R1117 GND.n3834 GND.n3833 585
R1118 GND.n3832 GND.n3831 585
R1119 GND.n3830 GND.n3829 585
R1120 GND.n3828 GND.n3827 585
R1121 GND.n3826 GND.n3825 585
R1122 GND.n3824 GND.n1527 585
R1123 GND.n3865 GND.n1528 585
R1124 GND.n3861 GND.n1529 585
R1125 GND.n3860 GND.n1530 585
R1126 GND.n1542 GND.n1531 585
R1127 GND.n3853 GND.n3852 585
R1128 GND.n3512 GND.n3511 585
R1129 GND.n3514 GND.n3513 585
R1130 GND.n3516 GND.n3515 585
R1131 GND.n3518 GND.n3517 585
R1132 GND.n3520 GND.n3519 585
R1133 GND.n3522 GND.n3521 585
R1134 GND.n3524 GND.n3523 585
R1135 GND.n3526 GND.n3525 585
R1136 GND.n3528 GND.n3527 585
R1137 GND.n3530 GND.n3529 585
R1138 GND.n3532 GND.n3531 585
R1139 GND.n3534 GND.n3533 585
R1140 GND.n3536 GND.n3535 585
R1141 GND.n3538 GND.n3537 585
R1142 GND.n3540 GND.n3539 585
R1143 GND.n3541 GND.n1917 585
R1144 GND.n3543 GND.n3542 585
R1145 GND.n1906 GND.n1905 585
R1146 GND.n3547 GND.n3546 585
R1147 GND.n3546 GND.n3545 585
R1148 GND.n3510 GND.n1938 585
R1149 GND.n3510 GND.n3509 585
R1150 GND.n3199 GND.n1896 585
R1151 GND.n3553 GND.n1896 585
R1152 GND.n3198 GND.n3197 585
R1153 GND.n3197 GND.n1895 585
R1154 GND.n3196 GND.n3193 585
R1155 GND.n3196 GND.n3195 585
R1156 GND.n2255 GND.n1884 585
R1157 GND.n3561 GND.n1884 585
R1158 GND.n3189 GND.n3188 585
R1159 GND.n3188 GND.n3187 585
R1160 GND.n3186 GND.n1873 585
R1161 GND.n3567 GND.n1873 585
R1162 GND.n3185 GND.n3184 585
R1163 GND.n3184 GND.n1872 585
R1164 GND.n3183 GND.n2257 585
R1165 GND.n3183 GND.n1861 585
R1166 GND.n3182 GND.n3158 585
R1167 GND.n3182 GND.n3181 585
R1168 GND.n2260 GND.n2259 585
R1169 GND.n2259 GND.n1829 585
R1170 GND.n3153 GND.n3152 585
R1171 GND.n3152 GND.n1822 585
R1172 GND.n3151 GND.n2262 585
R1173 GND.n3151 GND.n1820 585
R1174 GND.n3150 GND.n3149 585
R1175 GND.n3150 GND.n1806 585
R1176 GND.n2264 GND.n2263 585
R1177 GND.n3134 GND.n2263 585
R1178 GND.n3145 GND.n1797 585
R1179 GND.n3601 GND.n1797 585
R1180 GND.n3144 GND.n3143 585
R1181 GND.n3143 GND.n3142 585
R1182 GND.n2266 GND.n1787 585
R1183 GND.n3607 GND.n1787 585
R1184 GND.n3110 GND.n3109 585
R1185 GND.n3111 GND.n3110 585
R1186 GND.n2276 GND.n2275 585
R1187 GND.n2275 GND.n1778 585
R1188 GND.n3104 GND.n3103 585
R1189 GND.n3103 GND.n1776 585
R1190 GND.n3102 GND.n2278 585
R1191 GND.n3102 GND.n1770 585
R1192 GND.n3101 GND.n2280 585
R1193 GND.n3101 GND.n3100 585
R1194 GND.n3080 GND.n2279 585
R1195 GND.n2285 GND.n2279 585
R1196 GND.n3082 GND.n3081 585
R1197 GND.n3083 GND.n3082 585
R1198 GND.n2295 GND.n2294 585
R1199 GND.n2294 GND.n1753 585
R1200 GND.n3074 GND.n3073 585
R1201 GND.n3073 GND.n3072 585
R1202 GND.n2298 GND.n2297 585
R1203 GND.n2303 GND.n2298 585
R1204 GND.n3058 GND.n3057 585
R1205 GND.n3057 GND.n1741 585
R1206 GND.n3059 GND.n2312 585
R1207 GND.n2312 GND.n1735 585
R1208 GND.n3061 GND.n3060 585
R1209 GND.n3062 GND.n3061 585
R1210 GND.n2313 GND.n2311 585
R1211 GND.n3016 GND.n2311 585
R1212 GND.n3051 GND.n3050 585
R1213 GND.n3050 GND.n1723 585
R1214 GND.n3049 GND.n2315 585
R1215 GND.n3049 GND.n3048 585
R1216 GND.n2930 GND.n2316 585
R1217 GND.n3030 GND.n2316 585
R1218 GND.n2931 GND.n2332 585
R1219 GND.n3035 GND.n2332 585
R1220 GND.n2932 GND.n2924 585
R1221 GND.n2924 GND.n1706 585
R1222 GND.n2934 GND.n2933 585
R1223 GND.n2934 GND.n1700 585
R1224 GND.n2935 GND.n2923 585
R1225 GND.n2935 GND.n1698 585
R1226 GND.n2937 GND.n2936 585
R1227 GND.n2936 GND.n2337 585
R1228 GND.n2938 GND.n1683 585
R1229 GND.n3685 GND.n1683 585
R1230 GND.n2940 GND.n2939 585
R1231 GND.n2939 GND.n2340 585
R1232 GND.n2941 GND.n1672 585
R1233 GND.n3691 GND.n1672 585
R1234 GND.n2942 GND.n2348 585
R1235 GND.n2348 GND.n1664 585
R1236 GND.n2944 GND.n2943 585
R1237 GND.n2950 GND.n2944 585
R1238 GND.n2349 GND.n2347 585
R1239 GND.n2903 GND.n2347 585
R1240 GND.n2914 GND.n1652 585
R1241 GND.n3706 GND.n1652 585
R1242 GND.n2913 GND.n2912 585
R1243 GND.n2912 GND.t70 585
R1244 GND.n2877 GND.n1642 585
R1245 GND.n3712 GND.n1642 585
R1246 GND.n2353 GND.n2352 585
R1247 GND.n2352 GND.n2351 585
R1248 GND.n2873 GND.n1586 585
R1249 GND.n3791 GND.n1586 585
R1250 GND.n2872 GND.n2871 585
R1251 GND.n2871 GND.n2870 585
R1252 GND.n2869 GND.n1573 585
R1253 GND.n3797 GND.n1573 585
R1254 GND.n2863 GND.n2355 585
R1255 GND.n2863 GND.n1572 585
R1256 GND.n2865 GND.n2864 585
R1257 GND.n2864 GND.n1562 585
R1258 GND.n2862 GND.n1561 585
R1259 GND.n3805 GND.n1561 585
R1260 GND.n2861 GND.n2358 585
R1261 GND.n2473 GND.n2358 585
R1262 GND.n2357 GND.n1541 585
R1263 GND.n2475 GND.n1541 585
R1264 GND.n3577 GND.n3576 585
R1265 GND.n3576 GND.n3575 585
R1266 GND.n3578 GND.n1832 585
R1267 GND.n3160 GND.n1832 585
R1268 GND.n3580 GND.n3579 585
R1269 GND.n3581 GND.n3580 585
R1270 GND.n1833 GND.n1831 585
R1271 GND.n1831 GND.n1830 585
R1272 GND.n3126 GND.n1821 585
R1273 GND.n3587 GND.n1821 585
R1274 GND.n3128 GND.n3127 585
R1275 GND.t85 GND.n3128 585
R1276 GND.n1804 GND.n1803 585
R1277 GND.n3130 GND.n1804 585
R1278 GND.n3596 GND.n3595 585
R1279 GND.n3595 GND.n3594 585
R1280 GND.n3597 GND.n1801 585
R1281 GND.n3135 GND.n1801 585
R1282 GND.n3599 GND.n3598 585
R1283 GND.n3600 GND.n3599 585
R1284 GND.n1802 GND.n1800 585
R1285 GND.n3141 GND.n1800 585
R1286 GND.n3114 GND.n3113 585
R1287 GND.n3114 GND.n2268 585
R1288 GND.n3116 GND.n3115 585
R1289 GND.n3115 GND.n1788 585
R1290 GND.n3117 GND.n3112 585
R1291 GND.n3112 GND.n1786 585
R1292 GND.n3119 GND.n3118 585
R1293 GND.n3120 GND.n3119 585
R1294 GND.n1775 GND.n1774 585
R1295 GND.n2273 GND.n1775 585
R1296 GND.n3617 GND.n3616 585
R1297 GND.n3616 GND.n3615 585
R1298 GND.n3618 GND.n1772 585
R1299 GND.n2991 GND.n1772 585
R1300 GND.n3620 GND.n3619 585
R1301 GND.n3621 GND.n3620 585
R1302 GND.n1773 GND.n1771 585
R1303 GND.n1771 GND.n1768 585
R1304 GND.n2282 GND.n2281 585
R1305 GND.n2283 GND.n2282 585
R1306 GND.n1758 GND.n1757 585
R1307 GND.n1760 GND.n1758 585
R1308 GND.n3631 GND.n3630 585
R1309 GND.n3630 GND.n3629 585
R1310 GND.n3632 GND.n1755 585
R1311 GND.n2293 GND.n1755 585
R1312 GND.n3634 GND.n3633 585
R1313 GND.n3635 GND.n3634 585
R1314 GND.n1756 GND.n1754 585
R1315 GND.n1754 GND.n1751 585
R1316 GND.n2300 GND.n2299 585
R1317 GND.n2301 GND.n2300 585
R1318 GND.n1740 GND.n1739 585
R1319 GND.n1743 GND.n1740 585
R1320 GND.n3645 GND.n3644 585
R1321 GND.n3644 GND.n3643 585
R1322 GND.n3646 GND.n1737 585
R1323 GND.n3010 GND.n1737 585
R1324 GND.n3648 GND.n3647 585
R1325 GND.n3649 GND.n3648 585
R1326 GND.n1738 GND.n1736 585
R1327 GND.n1736 GND.n1733 585
R1328 GND.n3018 GND.n3017 585
R1329 GND.n3019 GND.n3018 585
R1330 GND.n1722 GND.n1721 585
R1331 GND.n1725 GND.n1722 585
R1332 GND.n3659 GND.n3658 585
R1333 GND.n3658 GND.n3657 585
R1334 GND.n3660 GND.n1719 585
R1335 GND.n2318 GND.n1719 585
R1336 GND.n3662 GND.n3661 585
R1337 GND.n3663 GND.n3662 585
R1338 GND.n1720 GND.n1718 585
R1339 GND.n1718 GND.n1716 585
R1340 GND.n3033 GND.n3032 585
R1341 GND.n3034 GND.n3033 585
R1342 GND.n1705 GND.n1704 585
R1343 GND.n1708 GND.n1705 585
R1344 GND.n3673 GND.n3672 585
R1345 GND.n3672 GND.n3671 585
R1346 GND.n3674 GND.n1702 585
R1347 GND.n2980 GND.n1702 585
R1348 GND.n3676 GND.n3675 585
R1349 GND.n3677 GND.n3676 585
R1350 GND.n1703 GND.n1701 585
R1351 GND.n2975 GND.n1701 585
R1352 GND.n2972 GND.n2971 585
R1353 GND.n2973 GND.n2972 585
R1354 GND.n2970 GND.n2338 585
R1355 GND.n2338 GND.n1684 585
R1356 GND.n2969 GND.n2968 585
R1357 GND.n2968 GND.n1682 585
R1358 GND.n2967 GND.n2339 585
R1359 GND.n2967 GND.n2966 585
R1360 GND.n1669 GND.n1668 585
R1361 GND.n2341 GND.n1669 585
R1362 GND.n3694 GND.n3693 585
R1363 GND.n3693 GND.n3692 585
R1364 GND.n3695 GND.n1666 585
R1365 GND.n2955 GND.n1666 585
R1366 GND.n3697 GND.n3696 585
R1367 GND.n3698 GND.n3697 585
R1368 GND.n1667 GND.n1665 585
R1369 GND.n2951 GND.n1665 585
R1370 GND.n2906 GND.n2905 585
R1371 GND.n2905 GND.n2904 585
R1372 GND.n2907 GND.n1653 585
R1373 GND.n3705 GND.n1653 585
R1374 GND.n2908 GND.n2900 585
R1375 GND.n2900 GND.n1651 585
R1376 GND.n2910 GND.n2909 585
R1377 GND.n2911 GND.n2910 585
R1378 GND.n2902 GND.n2899 585
R1379 GND.n2899 GND.n1643 585
R1380 GND.n2901 GND.n1608 585
R1381 GND.n3713 GND.n1608 585
R1382 GND.n3788 GND.n3787 585
R1383 GND.n3786 GND.n1607 585
R1384 GND.n3785 GND.n1606 585
R1385 GND.n3790 GND.n1606 585
R1386 GND.n3784 GND.n3783 585
R1387 GND.n3782 GND.n3781 585
R1388 GND.n3780 GND.n3779 585
R1389 GND.n3778 GND.n3777 585
R1390 GND.n3776 GND.n3775 585
R1391 GND.n3774 GND.n3773 585
R1392 GND.n3772 GND.n3771 585
R1393 GND.n3770 GND.n3769 585
R1394 GND.n3768 GND.n3767 585
R1395 GND.n3766 GND.n3765 585
R1396 GND.n3764 GND.n3763 585
R1397 GND.n3761 GND.n3760 585
R1398 GND.n3759 GND.n3758 585
R1399 GND.n3757 GND.n3756 585
R1400 GND.n3755 GND.n3754 585
R1401 GND.n3751 GND.n3750 585
R1402 GND.n3749 GND.n3748 585
R1403 GND.n3747 GND.n3746 585
R1404 GND.n3745 GND.n3744 585
R1405 GND.n3742 GND.n3741 585
R1406 GND.n3740 GND.n3739 585
R1407 GND.n3738 GND.n3737 585
R1408 GND.n3736 GND.n3735 585
R1409 GND.n3734 GND.n3733 585
R1410 GND.n3732 GND.n3731 585
R1411 GND.n3730 GND.n3729 585
R1412 GND.n3728 GND.n3727 585
R1413 GND.n3726 GND.n3725 585
R1414 GND.n3724 GND.n3723 585
R1415 GND.n3722 GND.n3721 585
R1416 GND.n3720 GND.n3719 585
R1417 GND.n3718 GND.n3717 585
R1418 GND.n3716 GND.n1604 585
R1419 GND.n3790 GND.n1604 585
R1420 GND.n2055 GND.n2054 585
R1421 GND.n2052 GND.n2018 585
R1422 GND.n2051 GND.n2050 585
R1423 GND.n2049 GND.n2048 585
R1424 GND.n2047 GND.n2046 585
R1425 GND.n2045 GND.n2044 585
R1426 GND.n2043 GND.n2042 585
R1427 GND.n2041 GND.n2040 585
R1428 GND.n2039 GND.n2038 585
R1429 GND.n2037 GND.n2036 585
R1430 GND.n2035 GND.n2034 585
R1431 GND.n2033 GND.n2032 585
R1432 GND.n2031 GND.n2030 585
R1433 GND.n2029 GND.n2028 585
R1434 GND.n2027 GND.n2026 585
R1435 GND.n2025 GND.n2024 585
R1436 GND.n2023 GND.n2022 585
R1437 GND.n2008 GND.n2005 585
R1438 GND.n2103 GND.n2102 585
R1439 GND.n2070 GND.n2006 585
R1440 GND.n2072 GND.n2071 585
R1441 GND.n2074 GND.n2073 585
R1442 GND.n2076 GND.n2075 585
R1443 GND.n2079 GND.n2078 585
R1444 GND.n2081 GND.n2080 585
R1445 GND.n2083 GND.n2082 585
R1446 GND.n2085 GND.n2084 585
R1447 GND.n2087 GND.n2086 585
R1448 GND.n2089 GND.n2088 585
R1449 GND.n2091 GND.n2090 585
R1450 GND.n2093 GND.n2092 585
R1451 GND.n2095 GND.n2094 585
R1452 GND.n2097 GND.n2096 585
R1453 GND.n2098 GND.n2065 585
R1454 GND.n2100 GND.n2099 585
R1455 GND.n2067 GND.n2064 585
R1456 GND.n2066 GND.n1859 585
R1457 GND.n2102 GND.n1859 585
R1458 GND.n2053 GND.n1860 585
R1459 GND.n3575 GND.n1860 585
R1460 GND.n1827 GND.n1826 585
R1461 GND.n3160 GND.n1827 585
R1462 GND.n3583 GND.n3582 585
R1463 GND.n3582 GND.n3581 585
R1464 GND.n3584 GND.n1824 585
R1465 GND.n1830 GND.n1824 585
R1466 GND.n3586 GND.n3585 585
R1467 GND.n3587 GND.n3586 585
R1468 GND.n1825 GND.n1823 585
R1469 GND.t85 GND.n1823 585
R1470 GND.n3132 GND.n3131 585
R1471 GND.n3131 GND.n3130 585
R1472 GND.n3133 GND.n1805 585
R1473 GND.n3594 GND.n1805 585
R1474 GND.n3137 GND.n3136 585
R1475 GND.n3136 GND.n3135 585
R1476 GND.n3138 GND.n1798 585
R1477 GND.n3600 GND.n1798 585
R1478 GND.n3140 GND.n3139 585
R1479 GND.n3141 GND.n3140 585
R1480 GND.n3125 GND.n2269 585
R1481 GND.n2269 GND.n2268 585
R1482 GND.n3124 GND.n3123 585
R1483 GND.n3123 GND.n1788 585
R1484 GND.n3122 GND.n2270 585
R1485 GND.n3122 GND.n1786 585
R1486 GND.n3121 GND.n2272 585
R1487 GND.n3121 GND.n3120 585
R1488 GND.n2988 GND.n2271 585
R1489 GND.n2273 GND.n2271 585
R1490 GND.n2989 GND.n1777 585
R1491 GND.n3615 GND.n1777 585
R1492 GND.n2993 GND.n2992 585
R1493 GND.n2992 GND.n2991 585
R1494 GND.n2994 GND.n1769 585
R1495 GND.n3621 GND.n1769 585
R1496 GND.n2996 GND.n2995 585
R1497 GND.n2996 GND.n1768 585
R1498 GND.n2997 GND.n2987 585
R1499 GND.n2997 GND.n2283 585
R1500 GND.n2999 GND.n2998 585
R1501 GND.n2998 GND.n1760 585
R1502 GND.n3000 GND.n1759 585
R1503 GND.n3629 GND.n1759 585
R1504 GND.n3002 GND.n3001 585
R1505 GND.n3001 GND.n2293 585
R1506 GND.n3003 GND.n1752 585
R1507 GND.n3635 GND.n1752 585
R1508 GND.n3005 GND.n3004 585
R1509 GND.n3005 GND.n1751 585
R1510 GND.n3006 GND.n2986 585
R1511 GND.n3006 GND.n2301 585
R1512 GND.n3008 GND.n3007 585
R1513 GND.n3007 GND.n1743 585
R1514 GND.n3009 GND.n1742 585
R1515 GND.n3643 GND.n1742 585
R1516 GND.n3012 GND.n3011 585
R1517 GND.n3011 GND.n3010 585
R1518 GND.n3013 GND.n1734 585
R1519 GND.n3649 GND.n1734 585
R1520 GND.n3015 GND.n3014 585
R1521 GND.n3015 GND.n1733 585
R1522 GND.n3020 GND.n2985 585
R1523 GND.n3020 GND.n3019 585
R1524 GND.n3022 GND.n3021 585
R1525 GND.n3021 GND.n1725 585
R1526 GND.n3023 GND.n1724 585
R1527 GND.n3657 GND.n1724 585
R1528 GND.n3025 GND.n3024 585
R1529 GND.n3024 GND.n2318 585
R1530 GND.n3026 GND.n1717 585
R1531 GND.n3663 GND.n1717 585
R1532 GND.n3027 GND.n2334 585
R1533 GND.n2334 GND.n1716 585
R1534 GND.n3029 GND.n3028 585
R1535 GND.n3034 GND.n3029 585
R1536 GND.n2984 GND.n2333 585
R1537 GND.n2333 GND.n1708 585
R1538 GND.n2983 GND.n1707 585
R1539 GND.n3671 GND.n1707 585
R1540 GND.n2982 GND.n2981 585
R1541 GND.n2981 GND.n2980 585
R1542 GND.n2978 GND.n1699 585
R1543 GND.n3677 GND.n1699 585
R1544 GND.n2977 GND.n2976 585
R1545 GND.n2976 GND.n2975 585
R1546 GND.n2336 GND.n2335 585
R1547 GND.n2973 GND.n2336 585
R1548 GND.n2961 GND.n2960 585
R1549 GND.n2960 GND.n1684 585
R1550 GND.n2962 GND.n2343 585
R1551 GND.n2343 GND.n1682 585
R1552 GND.n2964 GND.n2963 585
R1553 GND.n2966 GND.n2964 585
R1554 GND.n2959 GND.n2342 585
R1555 GND.n2342 GND.n2341 585
R1556 GND.n2958 GND.n1671 585
R1557 GND.n3692 GND.n1671 585
R1558 GND.n2957 GND.n2956 585
R1559 GND.n2956 GND.n2955 585
R1560 GND.n2954 GND.n1663 585
R1561 GND.n3698 GND.n1663 585
R1562 GND.n2953 GND.n2952 585
R1563 GND.n2952 GND.n2951 585
R1564 GND.n2345 GND.n2344 585
R1565 GND.n2904 GND.n2345 585
R1566 GND.n2894 GND.n1654 585
R1567 GND.n3705 GND.n1654 585
R1568 GND.n2895 GND.n2893 585
R1569 GND.n2893 GND.n1651 585
R1570 GND.n2897 GND.n2896 585
R1571 GND.n2911 GND.n2897 585
R1572 GND.n1640 GND.n1639 585
R1573 GND.n1643 GND.n1640 585
R1574 GND.n3715 GND.n3714 585
R1575 GND.n3714 GND.n3713 585
R1576 GND.n3949 GND.n3948 585
R1577 GND.n3950 GND.n3949 585
R1578 GND.n1418 GND.n1416 585
R1579 GND.n2839 GND.n1416 585
R1580 GND.n2835 GND.n2834 585
R1581 GND.n2836 GND.n2835 585
R1582 GND.n2386 GND.n2385 585
R1583 GND.n2816 GND.n2385 585
R1584 GND.n2830 GND.n2829 585
R1585 GND.n2829 GND.n2828 585
R1586 GND.n2389 GND.n2388 585
R1587 GND.n2824 GND.n2389 585
R1588 GND.n2806 GND.n2407 585
R1589 GND.n2407 GND.n2406 585
R1590 GND.n2809 GND.n2808 585
R1591 GND.n2810 GND.n2809 585
R1592 GND.n2805 GND.n2404 585
R1593 GND.n2798 GND.n2404 585
R1594 GND.n2803 GND.n2802 585
R1595 GND.n2802 GND.n2801 585
R1596 GND.n2409 GND.n2408 585
R1597 GND.n2795 GND.n2409 585
R1598 GND.n2782 GND.n2428 585
R1599 GND.n2428 GND.n2427 585
R1600 GND.n2784 GND.n2783 585
R1601 GND.n2785 GND.n2784 585
R1602 GND.n2780 GND.n2426 585
R1603 GND.n2773 GND.n2426 585
R1604 GND.n2778 GND.n2777 585
R1605 GND.n2777 GND.n2776 585
R1606 GND.n2432 GND.n2431 585
R1607 GND.n2771 GND.n2432 585
R1608 GND.n1367 GND.n1366 585
R1609 GND.n2518 GND.n1367 585
R1610 GND.n3983 GND.n3982 585
R1611 GND.n3982 GND.n3981 585
R1612 GND.n3984 GND.n1362 585
R1613 GND.n2761 GND.n1362 585
R1614 GND.n3986 GND.n3985 585
R1615 GND.n3987 GND.n3986 585
R1616 GND.n2595 GND.n1361 585
R1617 GND.n2598 GND.n2596 585
R1618 GND.n2601 GND.n2600 585
R1619 GND.n2592 GND.n2591 585
R1620 GND.n2606 GND.n2605 585
R1621 GND.n2608 GND.n2590 585
R1622 GND.n2611 GND.n2610 585
R1623 GND.n2588 GND.n2587 585
R1624 GND.n2616 GND.n2615 585
R1625 GND.n2618 GND.n2583 585
R1626 GND.n2621 GND.n2620 585
R1627 GND.n2581 GND.n2580 585
R1628 GND.n2626 GND.n2625 585
R1629 GND.n2628 GND.n2579 585
R1630 GND.n2631 GND.n2630 585
R1631 GND.n2577 GND.n2576 585
R1632 GND.n2636 GND.n2635 585
R1633 GND.n2638 GND.n2575 585
R1634 GND.n2641 GND.n2640 585
R1635 GND.n2573 GND.n2572 585
R1636 GND.n2647 GND.n2646 585
R1637 GND.n2649 GND.n2571 585
R1638 GND.n2652 GND.n2651 585
R1639 GND.n2653 GND.n2566 585
R1640 GND.n2657 GND.n2656 585
R1641 GND.n2659 GND.n2565 585
R1642 GND.n2662 GND.n2661 585
R1643 GND.n2563 GND.n2562 585
R1644 GND.n2667 GND.n2666 585
R1645 GND.n2669 GND.n2561 585
R1646 GND.n2672 GND.n2671 585
R1647 GND.n2559 GND.n2558 585
R1648 GND.n2677 GND.n2676 585
R1649 GND.n2679 GND.n2557 585
R1650 GND.n2682 GND.n2681 585
R1651 GND.n2555 GND.n2554 585
R1652 GND.n2689 GND.n2688 585
R1653 GND.n2691 GND.n2553 585
R1654 GND.n2694 GND.n2693 585
R1655 GND.n2551 GND.n2550 585
R1656 GND.n2699 GND.n2698 585
R1657 GND.n2701 GND.n2549 585
R1658 GND.n2704 GND.n2703 585
R1659 GND.n2547 GND.n2546 585
R1660 GND.n2709 GND.n2708 585
R1661 GND.n2711 GND.n2545 585
R1662 GND.n2714 GND.n2713 585
R1663 GND.n2543 GND.n2542 585
R1664 GND.n2719 GND.n2718 585
R1665 GND.n2721 GND.n2541 585
R1666 GND.n2723 GND.n2722 585
R1667 GND.n2722 GND.n1348 585
R1668 GND.n3870 GND.n1410 585
R1669 GND.n3871 GND.n1524 585
R1670 GND.n3872 GND.n1519 585
R1671 GND.n3873 GND.n1517 585
R1672 GND.n1516 GND.n1513 585
R1673 GND.n3877 GND.n1512 585
R1674 GND.n3878 GND.n1511 585
R1675 GND.n3879 GND.n1509 585
R1676 GND.n1508 GND.n1505 585
R1677 GND.n3883 GND.n1504 585
R1678 GND.n3884 GND.n1503 585
R1679 GND.n3885 GND.n1501 585
R1680 GND.n1500 GND.n1497 585
R1681 GND.n3889 GND.n1496 585
R1682 GND.n3890 GND.n1495 585
R1683 GND.n3891 GND.n1490 585
R1684 GND.n3892 GND.n1489 585
R1685 GND.n1487 GND.n1485 585
R1686 GND.n3896 GND.n1484 585
R1687 GND.n3897 GND.n1482 585
R1688 GND.n3898 GND.n1481 585
R1689 GND.n1479 GND.n1477 585
R1690 GND.n3902 GND.n1476 585
R1691 GND.n3903 GND.n1474 585
R1692 GND.n3904 GND.n1473 585
R1693 GND.n1469 GND.n1468 585
R1694 GND.n3909 GND.n3908 585
R1695 GND.n3914 GND.n3913 585
R1696 GND.n3915 GND.n1448 585
R1697 GND.n3916 GND.n1447 585
R1698 GND.n1454 GND.n1445 585
R1699 GND.n3920 GND.n1444 585
R1700 GND.n3921 GND.n1443 585
R1701 GND.n3922 GND.n1442 585
R1702 GND.n1457 GND.n1440 585
R1703 GND.n3926 GND.n1439 585
R1704 GND.n3927 GND.n1438 585
R1705 GND.n3928 GND.n1437 585
R1706 GND.n3931 GND.n1432 585
R1707 GND.n3932 GND.n1431 585
R1708 GND.n3933 GND.n1430 585
R1709 GND.n1461 GND.n1428 585
R1710 GND.n3937 GND.n1427 585
R1711 GND.n3938 GND.n1426 585
R1712 GND.n3939 GND.n1425 585
R1713 GND.n1464 GND.n1423 585
R1714 GND.n3943 GND.n1422 585
R1715 GND.n3944 GND.n1421 585
R1716 GND.n3945 GND.n1417 585
R1717 GND.n1467 GND.n1417 585
R1718 GND.n3952 GND.n3951 585
R1719 GND.n3951 GND.n3950 585
R1720 GND.n3953 GND.n1409 585
R1721 GND.n2839 GND.n1409 585
R1722 GND.n2384 GND.n1404 585
R1723 GND.n2836 GND.n2384 585
R1724 GND.n3957 GND.n1403 585
R1725 GND.n2816 GND.n1403 585
R1726 GND.n3958 GND.n1402 585
R1727 GND.n2828 GND.n1402 585
R1728 GND.n3959 GND.n1401 585
R1729 GND.n2824 GND.n1401 585
R1730 GND.n2405 GND.n1396 585
R1731 GND.n2406 GND.n2405 585
R1732 GND.n3963 GND.n1395 585
R1733 GND.n2810 GND.n1395 585
R1734 GND.n3964 GND.n1394 585
R1735 GND.n2798 GND.n1394 585
R1736 GND.n3965 GND.n1393 585
R1737 GND.n2801 GND.n1393 585
R1738 GND.n2415 GND.n1388 585
R1739 GND.n2795 GND.n2415 585
R1740 GND.n3969 GND.n1387 585
R1741 GND.n2427 GND.n1387 585
R1742 GND.n3970 GND.n1386 585
R1743 GND.n2785 GND.n1386 585
R1744 GND.n3971 GND.n1385 585
R1745 GND.n2773 GND.n1385 585
R1746 GND.n2434 GND.n1380 585
R1747 GND.n2776 GND.n2434 585
R1748 GND.n3975 GND.n1379 585
R1749 GND.n2771 GND.n1379 585
R1750 GND.n3976 GND.n1378 585
R1751 GND.n2518 GND.n1378 585
R1752 GND.n3977 GND.n1369 585
R1753 GND.n3981 GND.n1369 585
R1754 GND.n2760 GND.n1377 585
R1755 GND.n2761 GND.n2760 585
R1756 GND.n2726 GND.n1357 585
R1757 GND.n3987 GND.n1357 585
R1758 GND.n50 GND.n49 585
R1759 GND.n5474 GND.n50 585
R1760 GND.n5483 GND.n5482 585
R1761 GND.n5482 GND.n5481 585
R1762 GND.n5484 GND.n45 585
R1763 GND.n3326 GND.n45 585
R1764 GND.n5486 GND.n5485 585
R1765 GND.n5487 GND.n5486 585
R1766 GND.n28 GND.n26 585
R1767 GND.n3332 GND.n28 585
R1768 GND.n5495 GND.n5494 585
R1769 GND.n5494 GND.n5493 585
R1770 GND.n27 GND.n25 585
R1771 GND.n3338 GND.n27 585
R1772 GND.n2232 GND.n2231 585
R1773 GND.n2233 GND.n2232 585
R1774 GND.n17 GND.n15 585
R1775 GND.n3362 GND.n15 585
R1776 GND.n5499 GND.n5498 585
R1777 GND.n5500 GND.n5499 585
R1778 GND.n16 GND.n14 585
R1779 GND.n3368 GND.n14 585
R1780 GND.n2188 GND.n2187 585
R1781 GND.n2191 GND.n2188 585
R1782 GND.n3378 GND.n23 585
R1783 GND.n3378 GND.n3377 585
R1784 GND.n3380 GND.n3379 585
R1785 GND.n3381 GND.n3380 585
R1786 GND.n2169 GND.n2168 585
R1787 GND.n3254 GND.n2169 585
R1788 GND.n3389 GND.n3388 585
R1789 GND.n3388 GND.n3387 585
R1790 GND.n3390 GND.n2161 585
R1791 GND.n3239 GND.n2161 585
R1792 GND.n3392 GND.n3391 585
R1793 GND.n3393 GND.n3392 585
R1794 GND.n2162 GND.n2160 585
R1795 GND.n2246 GND.n2160 585
R1796 GND.n2163 GND.n1979 585
R1797 GND.n3401 GND.n1979 585
R1798 GND.n3498 GND.n3497 585
R1799 GND.n3496 GND.n1978 585
R1800 GND.n3495 GND.n1977 585
R1801 GND.n3500 GND.n1977 585
R1802 GND.n3494 GND.n3493 585
R1803 GND.n3492 GND.n3491 585
R1804 GND.n3490 GND.n3489 585
R1805 GND.n3488 GND.n3487 585
R1806 GND.n3486 GND.n3485 585
R1807 GND.n3484 GND.n3483 585
R1808 GND.n3482 GND.n3481 585
R1809 GND.n3480 GND.n3479 585
R1810 GND.n3478 GND.n3477 585
R1811 GND.n3476 GND.n3475 585
R1812 GND.n3474 GND.n3473 585
R1813 GND.n3472 GND.n3471 585
R1814 GND.n3470 GND.n3469 585
R1815 GND.n3468 GND.n3467 585
R1816 GND.n3466 GND.n3465 585
R1817 GND.n3464 GND.n3463 585
R1818 GND.n3462 GND.n3461 585
R1819 GND.n3460 GND.n3459 585
R1820 GND.n3458 GND.n3457 585
R1821 GND.n3455 GND.n3454 585
R1822 GND.n3453 GND.n3452 585
R1823 GND.n3451 GND.n3450 585
R1824 GND.n3449 GND.n3448 585
R1825 GND.n3447 GND.n3446 585
R1826 GND.n3445 GND.n3444 585
R1827 GND.n3443 GND.n3442 585
R1828 GND.n3441 GND.n3440 585
R1829 GND.n3439 GND.n3438 585
R1830 GND.n3437 GND.n3436 585
R1831 GND.n3435 GND.n3434 585
R1832 GND.n3433 GND.n3432 585
R1833 GND.n3431 GND.n2122 585
R1834 GND.n3430 GND.n3429 585
R1835 GND.n3428 GND.n3427 585
R1836 GND.n3426 GND.n3425 585
R1837 GND.n3424 GND.n3423 585
R1838 GND.n3422 GND.n3421 585
R1839 GND.n3420 GND.n3419 585
R1840 GND.n3418 GND.n3417 585
R1841 GND.n3416 GND.n3415 585
R1842 GND.n3414 GND.n3413 585
R1843 GND.n3412 GND.n3411 585
R1844 GND.n3410 GND.n3409 585
R1845 GND.n3408 GND.n2137 585
R1846 GND.n2141 GND.n2138 585
R1847 GND.n3404 GND.n3403 585
R1848 GND.n149 GND.n59 585
R1849 GND.n155 GND.n154 585
R1850 GND.n157 GND.n156 585
R1851 GND.n159 GND.n158 585
R1852 GND.n161 GND.n160 585
R1853 GND.n163 GND.n162 585
R1854 GND.n165 GND.n164 585
R1855 GND.n167 GND.n166 585
R1856 GND.n169 GND.n168 585
R1857 GND.n171 GND.n170 585
R1858 GND.n173 GND.n172 585
R1859 GND.n175 GND.n174 585
R1860 GND.n177 GND.n176 585
R1861 GND.n137 GND.n134 585
R1862 GND.n181 GND.n138 585
R1863 GND.n183 GND.n182 585
R1864 GND.n185 GND.n184 585
R1865 GND.n187 GND.n186 585
R1866 GND.n189 GND.n188 585
R1867 GND.n191 GND.n190 585
R1868 GND.n193 GND.n192 585
R1869 GND.n195 GND.n194 585
R1870 GND.n197 GND.n196 585
R1871 GND.n199 GND.n198 585
R1872 GND.n201 GND.n200 585
R1873 GND.n203 GND.n202 585
R1874 GND.n205 GND.n204 585
R1875 GND.n210 GND.n209 585
R1876 GND.n212 GND.n211 585
R1877 GND.n214 GND.n213 585
R1878 GND.n216 GND.n215 585
R1879 GND.n218 GND.n217 585
R1880 GND.n220 GND.n219 585
R1881 GND.n222 GND.n221 585
R1882 GND.n224 GND.n223 585
R1883 GND.n226 GND.n225 585
R1884 GND.n228 GND.n227 585
R1885 GND.n230 GND.n229 585
R1886 GND.n232 GND.n231 585
R1887 GND.n234 GND.n233 585
R1888 GND.n236 GND.n235 585
R1889 GND.n238 GND.n237 585
R1890 GND.n240 GND.n239 585
R1891 GND.n242 GND.n241 585
R1892 GND.n244 GND.n243 585
R1893 GND.n246 GND.n245 585
R1894 GND.n248 GND.n247 585
R1895 GND.n251 GND.n250 585
R1896 GND.n249 GND.n98 585
R1897 GND.n255 GND.n95 585
R1898 GND.n257 GND.n256 585
R1899 GND.n258 GND.n257 585
R1900 GND.n5476 GND.n5475 585
R1901 GND.n5475 GND.n5474 585
R1902 GND.n58 GND.n52 585
R1903 GND.n5481 GND.n52 585
R1904 GND.n3328 GND.n3327 585
R1905 GND.n3327 GND.n3326 585
R1906 GND.n3329 GND.n42 585
R1907 GND.n5487 GND.n42 585
R1908 GND.n3331 GND.n3330 585
R1909 GND.n3332 GND.n3331 585
R1910 GND.n3271 GND.n30 585
R1911 GND.n5493 GND.n30 585
R1912 GND.n3270 GND.n2234 585
R1913 GND.n3338 GND.n2234 585
R1914 GND.n3267 GND.n3266 585
R1915 GND.n3266 GND.n2233 585
R1916 GND.n3265 GND.n2230 585
R1917 GND.n3362 GND.n2230 585
R1918 GND.n3264 GND.n11 585
R1919 GND.n5500 GND.n11 585
R1920 GND.n3263 GND.n2222 585
R1921 GND.n3368 GND.n2222 585
R1922 GND.n3262 GND.n3261 585
R1923 GND.n3261 GND.n2191 585
R1924 GND.n3258 GND.n2189 585
R1925 GND.n3377 GND.n2189 585
R1926 GND.n3257 GND.n2184 585
R1927 GND.n3381 GND.n2184 585
R1928 GND.n3256 GND.n3255 585
R1929 GND.n3255 GND.n3254 585
R1930 GND.n2242 GND.n2171 585
R1931 GND.n3387 GND.n2171 585
R1932 GND.n2155 GND.n2154 585
R1933 GND.n3239 GND.n2155 585
R1934 GND.n3395 GND.n3394 585
R1935 GND.n3394 GND.n3393 585
R1936 GND.n3396 GND.n2144 585
R1937 GND.n2246 GND.n2144 585
R1938 GND.n3402 GND.n2145 585
R1939 GND.n3402 GND.n3401 585
R1940 GND.n1139 GND.n1138 585
R1941 GND.n4203 GND.n1139 585
R1942 GND.n5254 GND.n465 585
R1943 GND.n5258 GND.n465 585
R1944 GND.n5261 GND.n5260 585
R1945 GND.n5260 GND.n5259 585
R1946 GND.n5262 GND.n460 585
R1947 GND.n460 GND.n459 585
R1948 GND.n5264 GND.n5263 585
R1949 GND.n5265 GND.n5264 585
R1950 GND.n458 GND.n457 585
R1951 GND.n5266 GND.n458 585
R1952 GND.n5269 GND.n5268 585
R1953 GND.n5268 GND.n5267 585
R1954 GND.n5270 GND.n452 585
R1955 GND.n452 GND.n451 585
R1956 GND.n5272 GND.n5271 585
R1957 GND.n5273 GND.n5272 585
R1958 GND.n450 GND.n449 585
R1959 GND.n5274 GND.n450 585
R1960 GND.n5277 GND.n5276 585
R1961 GND.n5276 GND.n5275 585
R1962 GND.n5278 GND.n444 585
R1963 GND.n444 GND.n443 585
R1964 GND.n5280 GND.n5279 585
R1965 GND.n5281 GND.n5280 585
R1966 GND.n442 GND.n441 585
R1967 GND.n5282 GND.n442 585
R1968 GND.n5285 GND.n5284 585
R1969 GND.n5284 GND.n5283 585
R1970 GND.n5286 GND.n436 585
R1971 GND.n436 GND.n435 585
R1972 GND.n5288 GND.n5287 585
R1973 GND.n5289 GND.n5288 585
R1974 GND.n434 GND.n433 585
R1975 GND.n5290 GND.n434 585
R1976 GND.n5293 GND.n5292 585
R1977 GND.n5292 GND.n5291 585
R1978 GND.n5294 GND.n428 585
R1979 GND.n428 GND.n427 585
R1980 GND.n5296 GND.n5295 585
R1981 GND.n5297 GND.n5296 585
R1982 GND.n426 GND.n425 585
R1983 GND.n5298 GND.n426 585
R1984 GND.n5301 GND.n5300 585
R1985 GND.n5300 GND.n5299 585
R1986 GND.n5302 GND.n420 585
R1987 GND.n420 GND.n419 585
R1988 GND.n5304 GND.n5303 585
R1989 GND.n5305 GND.n5304 585
R1990 GND.n418 GND.n417 585
R1991 GND.n5306 GND.n418 585
R1992 GND.n5309 GND.n5308 585
R1993 GND.n5308 GND.n5307 585
R1994 GND.n5310 GND.n412 585
R1995 GND.n412 GND.n411 585
R1996 GND.n5312 GND.n5311 585
R1997 GND.n5313 GND.n5312 585
R1998 GND.n410 GND.n409 585
R1999 GND.n5314 GND.n410 585
R2000 GND.n5317 GND.n5316 585
R2001 GND.n5316 GND.n5315 585
R2002 GND.n5318 GND.n404 585
R2003 GND.n404 GND.n403 585
R2004 GND.n5320 GND.n5319 585
R2005 GND.n5321 GND.n5320 585
R2006 GND.n402 GND.n401 585
R2007 GND.n5322 GND.n402 585
R2008 GND.n5325 GND.n5324 585
R2009 GND.n5324 GND.n5323 585
R2010 GND.n5326 GND.n396 585
R2011 GND.n396 GND.n395 585
R2012 GND.n5328 GND.n5327 585
R2013 GND.n5329 GND.n5328 585
R2014 GND.n394 GND.n393 585
R2015 GND.n5330 GND.n394 585
R2016 GND.n5333 GND.n5332 585
R2017 GND.n5332 GND.n5331 585
R2018 GND.n5334 GND.n388 585
R2019 GND.n388 GND.n387 585
R2020 GND.n5336 GND.n5335 585
R2021 GND.n5337 GND.n5336 585
R2022 GND.n386 GND.n385 585
R2023 GND.n5338 GND.n386 585
R2024 GND.n5341 GND.n5340 585
R2025 GND.n5340 GND.n5339 585
R2026 GND.n5342 GND.n380 585
R2027 GND.n380 GND.n379 585
R2028 GND.n5344 GND.n5343 585
R2029 GND.n5345 GND.n5344 585
R2030 GND.n378 GND.n377 585
R2031 GND.n5346 GND.n378 585
R2032 GND.n5349 GND.n5348 585
R2033 GND.n5348 GND.n5347 585
R2034 GND.n5350 GND.n372 585
R2035 GND.n372 GND.n371 585
R2036 GND.n5352 GND.n5351 585
R2037 GND.n5353 GND.n5352 585
R2038 GND.n370 GND.n369 585
R2039 GND.n5354 GND.n370 585
R2040 GND.n5357 GND.n5356 585
R2041 GND.n5356 GND.n5355 585
R2042 GND.n5358 GND.n364 585
R2043 GND.n364 GND.n363 585
R2044 GND.n5360 GND.n5359 585
R2045 GND.n5361 GND.n5360 585
R2046 GND.n362 GND.n361 585
R2047 GND.n5362 GND.n362 585
R2048 GND.n5365 GND.n5364 585
R2049 GND.n5364 GND.n5363 585
R2050 GND.n5366 GND.n356 585
R2051 GND.n356 GND.n355 585
R2052 GND.n5368 GND.n5367 585
R2053 GND.n5369 GND.n5368 585
R2054 GND.n354 GND.n353 585
R2055 GND.n5370 GND.n354 585
R2056 GND.n5373 GND.n5372 585
R2057 GND.n5372 GND.n5371 585
R2058 GND.n5374 GND.n348 585
R2059 GND.n348 GND.n347 585
R2060 GND.n5376 GND.n5375 585
R2061 GND.n5377 GND.n5376 585
R2062 GND.n346 GND.n345 585
R2063 GND.n5378 GND.n346 585
R2064 GND.n5381 GND.n5380 585
R2065 GND.n5380 GND.n5379 585
R2066 GND.n5382 GND.n340 585
R2067 GND.n340 GND.n339 585
R2068 GND.n5384 GND.n5383 585
R2069 GND.n5385 GND.n5384 585
R2070 GND.n338 GND.n337 585
R2071 GND.n5386 GND.n338 585
R2072 GND.n5389 GND.n5388 585
R2073 GND.n5388 GND.n5387 585
R2074 GND.n5390 GND.n332 585
R2075 GND.n332 GND.n331 585
R2076 GND.n5392 GND.n5391 585
R2077 GND.n5393 GND.n5392 585
R2078 GND.n330 GND.n329 585
R2079 GND.n5394 GND.n330 585
R2080 GND.n5397 GND.n5396 585
R2081 GND.n5396 GND.n5395 585
R2082 GND.n5398 GND.n324 585
R2083 GND.n324 GND.n323 585
R2084 GND.n5400 GND.n5399 585
R2085 GND.n5401 GND.n5400 585
R2086 GND.n322 GND.n321 585
R2087 GND.n5402 GND.n322 585
R2088 GND.n5405 GND.n5404 585
R2089 GND.n5404 GND.n5403 585
R2090 GND.n5406 GND.n316 585
R2091 GND.n316 GND.n315 585
R2092 GND.n5408 GND.n5407 585
R2093 GND.n5409 GND.n5408 585
R2094 GND.n314 GND.n313 585
R2095 GND.n5410 GND.n314 585
R2096 GND.n5413 GND.n5412 585
R2097 GND.n5412 GND.n5411 585
R2098 GND.n5414 GND.n308 585
R2099 GND.n308 GND.n307 585
R2100 GND.n5416 GND.n5415 585
R2101 GND.n5417 GND.n5416 585
R2102 GND.n306 GND.n305 585
R2103 GND.n5418 GND.n306 585
R2104 GND.n5421 GND.n5420 585
R2105 GND.n5420 GND.n5419 585
R2106 GND.n5422 GND.n300 585
R2107 GND.n300 GND.n299 585
R2108 GND.n5424 GND.n5423 585
R2109 GND.n5425 GND.n5424 585
R2110 GND.n298 GND.n297 585
R2111 GND.n5426 GND.n298 585
R2112 GND.n5429 GND.n5428 585
R2113 GND.n5428 GND.n5427 585
R2114 GND.n5430 GND.n292 585
R2115 GND.n292 GND.n291 585
R2116 GND.n5432 GND.n5431 585
R2117 GND.n5433 GND.n5432 585
R2118 GND.n290 GND.n289 585
R2119 GND.n5434 GND.n290 585
R2120 GND.n5437 GND.n5436 585
R2121 GND.n5436 GND.n5435 585
R2122 GND.n5438 GND.n284 585
R2123 GND.n284 GND.n283 585
R2124 GND.n5440 GND.n5439 585
R2125 GND.n5441 GND.n5440 585
R2126 GND.n282 GND.n281 585
R2127 GND.n5442 GND.n282 585
R2128 GND.n5445 GND.n5444 585
R2129 GND.n5444 GND.n5443 585
R2130 GND.n5446 GND.n276 585
R2131 GND.n276 GND.n275 585
R2132 GND.n5448 GND.n5447 585
R2133 GND.n5449 GND.n5448 585
R2134 GND.n274 GND.n273 585
R2135 GND.n5450 GND.n274 585
R2136 GND.n5453 GND.n5452 585
R2137 GND.n5452 GND.n5451 585
R2138 GND.n5454 GND.n268 585
R2139 GND.n268 GND.n267 585
R2140 GND.n5456 GND.n5455 585
R2141 GND.n5457 GND.n5456 585
R2142 GND.n266 GND.n265 585
R2143 GND.n5458 GND.n266 585
R2144 GND.n5461 GND.n5460 585
R2145 GND.n5460 GND.n5459 585
R2146 GND.n5462 GND.n260 585
R2147 GND.n260 GND.n259 585
R2148 GND.n5464 GND.n5463 585
R2149 GND.n5465 GND.n5464 585
R2150 GND.n69 GND.n68 585
R2151 GND.n5466 GND.n69 585
R2152 GND.n5469 GND.n5468 585
R2153 GND.n5468 GND.n5467 585
R2154 GND.n5470 GND.n63 585
R2155 GND.n63 GND.n61 585
R2156 GND.n5472 GND.n5471 585
R2157 GND.n5473 GND.n5472 585
R2158 GND.n64 GND.n62 585
R2159 GND.n62 GND.n54 585
R2160 GND.n3349 GND.n3348 585
R2161 GND.n3349 GND.n51 585
R2162 GND.n3351 GND.n3350 585
R2163 GND.n3350 GND.n44 585
R2164 GND.n3352 GND.n3343 585
R2165 GND.n3343 GND.n41 585
R2166 GND.n3354 GND.n3353 585
R2167 GND.n3354 GND.n32 585
R2168 GND.n3356 GND.n3355 585
R2169 GND.n3355 GND.n29 585
R2170 GND.n3357 GND.n3340 585
R2171 GND.n3340 GND.n3339 585
R2172 GND.n3360 GND.n3359 585
R2173 GND.n3361 GND.n3360 585
R2174 GND.n3341 GND.n2220 585
R2175 GND.n2220 GND.n12 585
R2176 GND.n3371 GND.n3370 585
R2177 GND.n3370 GND.n3369 585
R2178 GND.n3372 GND.n2193 585
R2179 GND.n2221 GND.n2193 585
R2180 GND.n3375 GND.n3374 585
R2181 GND.n3376 GND.n3375 585
R2182 GND.n2218 GND.n2192 585
R2183 GND.n2192 GND.n2186 585
R2184 GND.n2216 GND.n2215 585
R2185 GND.n2215 GND.n2183 585
R2186 GND.n2214 GND.n2194 585
R2187 GND.n2214 GND.n2173 585
R2188 GND.n2213 GND.n2212 585
R2189 GND.n2213 GND.n2170 585
R2190 GND.n2196 GND.n2195 585
R2191 GND.n2195 GND.n2158 585
R2192 GND.n2207 GND.n2206 585
R2193 GND.n2206 GND.n2156 585
R2194 GND.n2205 GND.n2198 585
R2195 GND.n2205 GND.n2148 585
R2196 GND.n2204 GND.n2203 585
R2197 GND.n2204 GND.n2146 585
R2198 GND.n2199 GND.n1945 585
R2199 GND.n1976 GND.n1945 585
R2200 GND.n3502 GND.n1944 585
R2201 GND.n3502 GND.n3501 585
R2202 GND.n3504 GND.n3503 585
R2203 GND.n3503 GND.n1908 585
R2204 GND.n3505 GND.n1939 585
R2205 GND.n1939 GND.n1907 585
R2206 GND.n3507 GND.n3506 585
R2207 GND.n3508 GND.n3507 585
R2208 GND.n1894 GND.n1893 585
R2209 GND.n1897 GND.n1894 585
R2210 GND.n3556 GND.n3555 585
R2211 GND.n3555 GND.n3554 585
R2212 GND.n3557 GND.n1886 585
R2213 GND.n3194 GND.n1886 585
R2214 GND.n3559 GND.n3558 585
R2215 GND.n3560 GND.n3559 585
R2216 GND.n1887 GND.n1885 585
R2217 GND.n1885 GND.n1883 585
R2218 GND.n1871 GND.n1870 585
R2219 GND.n1874 GND.n1871 585
R2220 GND.n3570 GND.n3569 585
R2221 GND.n3569 GND.n3568 585
R2222 GND.n3571 GND.n1863 585
R2223 GND.n2009 GND.n1863 585
R2224 GND.n3573 GND.n3572 585
R2225 GND.n3574 GND.n3573 585
R2226 GND.n1864 GND.n1862 585
R2227 GND.n3159 GND.n1862 585
R2228 GND.n1819 GND.n1818 585
R2229 GND.n1828 GND.n1819 585
R2230 GND.n3589 GND.n3588 585
R2231 GND.n3588 GND.n3587 585
R2232 GND.n3590 GND.n1808 585
R2233 GND.n3129 GND.n1808 585
R2234 GND.n3592 GND.n3591 585
R2235 GND.n3593 GND.n3592 585
R2236 GND.n1809 GND.n1807 585
R2237 GND.n1807 GND.n1799 585
R2238 GND.n1812 GND.n1811 585
R2239 GND.n1811 GND.t104 585
R2240 GND.n1785 GND.n1784 585
R2241 GND.n2267 GND.n1785 585
R2242 GND.n3610 GND.n3609 585
R2243 GND.n3609 GND.n3608 585
R2244 GND.n3611 GND.n1779 585
R2245 GND.n2274 GND.n1779 585
R2246 GND.n3613 GND.n3612 585
R2247 GND.n3614 GND.n3613 585
R2248 GND.n1767 GND.n1766 585
R2249 GND.n2990 GND.n1767 585
R2250 GND.n3624 GND.n3623 585
R2251 GND.n3623 GND.n3622 585
R2252 GND.n3625 GND.n1761 585
R2253 GND.n2284 GND.n1761 585
R2254 GND.n3627 GND.n3626 585
R2255 GND.n3628 GND.n3627 585
R2256 GND.n1750 GND.n1749 585
R2257 GND.n2292 GND.n1750 585
R2258 GND.n3638 GND.n3637 585
R2259 GND.n3637 GND.n3636 585
R2260 GND.n3639 GND.n1744 585
R2261 GND.n2302 GND.n1744 585
R2262 GND.n3641 GND.n3640 585
R2263 GND.n3642 GND.n3641 585
R2264 GND.n1732 GND.n1731 585
R2265 GND.n3010 GND.n1732 585
R2266 GND.n3652 GND.n3651 585
R2267 GND.n3651 GND.n3650 585
R2268 GND.n3653 GND.n1726 585
R2269 GND.n2310 GND.n1726 585
R2270 GND.n3655 GND.n3654 585
R2271 GND.n3656 GND.n3655 585
R2272 GND.n1715 GND.n1714 585
R2273 GND.n2317 GND.n1715 585
R2274 GND.n3666 GND.n3665 585
R2275 GND.n3665 GND.n3664 585
R2276 GND.n3667 GND.n1709 585
R2277 GND.n3031 GND.n1709 585
R2278 GND.n3669 GND.n3668 585
R2279 GND.n3670 GND.n3669 585
R2280 GND.n1697 GND.n1696 585
R2281 GND.n2979 GND.n1697 585
R2282 GND.n3680 GND.n3679 585
R2283 GND.n3679 GND.n3678 585
R2284 GND.n3681 GND.n1686 585
R2285 GND.n2974 GND.n1686 585
R2286 GND.n3683 GND.n3682 585
R2287 GND.n3684 GND.n3683 585
R2288 GND.n1687 GND.n1685 585
R2289 GND.n2965 GND.n1685 585
R2290 GND.n1690 GND.n1689 585
R2291 GND.n1689 GND.n1673 585
R2292 GND.n1662 GND.n1661 585
R2293 GND.n1670 GND.n1662 585
R2294 GND.n3701 GND.n3700 585
R2295 GND.n3700 GND.n3699 585
R2296 GND.n3702 GND.n1656 585
R2297 GND.n2346 GND.n1656 585
R2298 GND.n3704 GND.n3703 585
R2299 GND.n3705 GND.n3704 585
R2300 GND.n1657 GND.n1655 585
R2301 GND.n2898 GND.n1655 585
R2302 GND.n2891 GND.n2890 585
R2303 GND.n2892 GND.n2891 585
R2304 GND.n2879 GND.n2878 585
R2305 GND.n2878 GND.n1641 585
R2306 GND.n2885 GND.n2884 585
R2307 GND.n2884 GND.n1605 585
R2308 GND.n2883 GND.n2882 585
R2309 GND.n2883 GND.n1585 585
R2310 GND.n1570 GND.n1569 585
R2311 GND.n1574 GND.n1570 585
R2312 GND.n3800 GND.n3799 585
R2313 GND.n3799 GND.n3798 585
R2314 GND.n3801 GND.n1564 585
R2315 GND.n1571 GND.n1564 585
R2316 GND.n3803 GND.n3802 585
R2317 GND.n3804 GND.n3803 585
R2318 GND.n1565 GND.n1563 585
R2319 GND.n1563 GND.n1560 585
R2320 GND.n2472 GND.n2471 585
R2321 GND.n2474 GND.n2472 585
R2322 GND.n2477 GND.n2467 585
R2323 GND.n2477 GND.n2476 585
R2324 GND.n2479 GND.n2478 585
R2325 GND.n2478 GND.n1551 585
R2326 GND.n2480 GND.n2462 585
R2327 GND.n2462 GND.n1543 585
R2328 GND.n2483 GND.n2481 585
R2329 GND.n2483 GND.n2482 585
R2330 GND.n2485 GND.n2461 585
R2331 GND.n2485 GND.n2484 585
R2332 GND.n2487 GND.n2486 585
R2333 GND.n2486 GND.n1413 585
R2334 GND.n2488 GND.n2456 585
R2335 GND.n2456 GND.n1411 585
R2336 GND.n2490 GND.n2489 585
R2337 GND.n2490 GND.n2381 585
R2338 GND.n2491 GND.n2455 585
R2339 GND.n2491 GND.n2383 585
R2340 GND.n2493 GND.n2492 585
R2341 GND.n2492 GND.n2392 585
R2342 GND.n2494 GND.n2453 585
R2343 GND.n2453 GND.n2390 585
R2344 GND.n2496 GND.n2495 585
R2345 GND.n2496 GND.n2394 585
R2346 GND.n2498 GND.n2497 585
R2347 GND.n2497 GND.n2402 585
R2348 GND.n2500 GND.n2499 585
R2349 GND.n2500 GND.n2401 585
R2350 GND.n2502 GND.n2501 585
R2351 GND.n2501 GND.n2412 585
R2352 GND.n2504 GND.n2503 585
R2353 GND.n2504 GND.n2410 585
R2354 GND.n2506 GND.n2505 585
R2355 GND.n2506 GND.n2414 585
R2356 GND.n2507 GND.n2451 585
R2357 GND.n2507 GND.n2423 585
R2358 GND.n2509 GND.n2508 585
R2359 GND.n2508 GND.n2422 585
R2360 GND.n2452 GND.n2446 585
R2361 GND.n2452 GND.n2436 585
R2362 GND.n2513 GND.n2445 585
R2363 GND.n2445 GND.n2433 585
R2364 GND.n2514 GND.n2439 585
R2365 GND.n2439 GND.n2437 585
R2366 GND.n2516 GND.n2515 585
R2367 GND.n2517 GND.n2516 585
R2368 GND.n2440 GND.n2438 585
R2369 GND.n2438 GND.n1368 585
R2370 GND.n1355 GND.n1354 585
R2371 GND.n1359 GND.n1355 585
R2372 GND.n3990 GND.n3989 585
R2373 GND.n3989 GND.n3988 585
R2374 GND.n3991 GND.n1349 585
R2375 GND.n1356 GND.n1349 585
R2376 GND.n3993 GND.n3992 585
R2377 GND.n3994 GND.n3993 585
R2378 GND.n1347 GND.n1346 585
R2379 GND.n3995 GND.n1347 585
R2380 GND.n3998 GND.n3997 585
R2381 GND.n3997 GND.n3996 585
R2382 GND.n3999 GND.n1341 585
R2383 GND.n1341 GND.n1340 585
R2384 GND.n4001 GND.n4000 585
R2385 GND.n4002 GND.n4001 585
R2386 GND.n1339 GND.n1338 585
R2387 GND.n4003 GND.n1339 585
R2388 GND.n4006 GND.n4005 585
R2389 GND.n4005 GND.n4004 585
R2390 GND.n4007 GND.n1333 585
R2391 GND.n1333 GND.n1332 585
R2392 GND.n4009 GND.n4008 585
R2393 GND.n4010 GND.n4009 585
R2394 GND.n1331 GND.n1330 585
R2395 GND.n4011 GND.n1331 585
R2396 GND.n4014 GND.n4013 585
R2397 GND.n4013 GND.n4012 585
R2398 GND.n4015 GND.n1325 585
R2399 GND.n1325 GND.n1324 585
R2400 GND.n4017 GND.n4016 585
R2401 GND.n4018 GND.n4017 585
R2402 GND.n1323 GND.n1322 585
R2403 GND.n4019 GND.n1323 585
R2404 GND.n4022 GND.n4021 585
R2405 GND.n4021 GND.n4020 585
R2406 GND.n4023 GND.n1317 585
R2407 GND.n1317 GND.n1316 585
R2408 GND.n4025 GND.n4024 585
R2409 GND.n4026 GND.n4025 585
R2410 GND.n1315 GND.n1314 585
R2411 GND.n4027 GND.n1315 585
R2412 GND.n4030 GND.n4029 585
R2413 GND.n4029 GND.n4028 585
R2414 GND.n4031 GND.n1309 585
R2415 GND.n1309 GND.n1308 585
R2416 GND.n4033 GND.n4032 585
R2417 GND.n4034 GND.n4033 585
R2418 GND.n1307 GND.n1306 585
R2419 GND.n4035 GND.n1307 585
R2420 GND.n4038 GND.n4037 585
R2421 GND.n4037 GND.n4036 585
R2422 GND.n4039 GND.n1301 585
R2423 GND.n1301 GND.n1300 585
R2424 GND.n4041 GND.n4040 585
R2425 GND.n4042 GND.n4041 585
R2426 GND.n1299 GND.n1298 585
R2427 GND.n4043 GND.n1299 585
R2428 GND.n4046 GND.n4045 585
R2429 GND.n4045 GND.n4044 585
R2430 GND.n4047 GND.n1293 585
R2431 GND.n1293 GND.n1292 585
R2432 GND.n4049 GND.n4048 585
R2433 GND.n4050 GND.n4049 585
R2434 GND.n1291 GND.n1290 585
R2435 GND.n4051 GND.n1291 585
R2436 GND.n4054 GND.n4053 585
R2437 GND.n4053 GND.n4052 585
R2438 GND.n4055 GND.n1285 585
R2439 GND.n1285 GND.n1284 585
R2440 GND.n4057 GND.n4056 585
R2441 GND.n4058 GND.n4057 585
R2442 GND.n1283 GND.n1282 585
R2443 GND.n4059 GND.n1283 585
R2444 GND.n4062 GND.n4061 585
R2445 GND.n4061 GND.n4060 585
R2446 GND.n4063 GND.n1277 585
R2447 GND.n1277 GND.n1276 585
R2448 GND.n4065 GND.n4064 585
R2449 GND.n4066 GND.n4065 585
R2450 GND.n1275 GND.n1274 585
R2451 GND.n4067 GND.n1275 585
R2452 GND.n4070 GND.n4069 585
R2453 GND.n4069 GND.n4068 585
R2454 GND.n4071 GND.n1269 585
R2455 GND.n1269 GND.n1268 585
R2456 GND.n4073 GND.n4072 585
R2457 GND.n4074 GND.n4073 585
R2458 GND.n1267 GND.n1266 585
R2459 GND.n4075 GND.n1267 585
R2460 GND.n4078 GND.n4077 585
R2461 GND.n4077 GND.n4076 585
R2462 GND.n4079 GND.n1261 585
R2463 GND.n1261 GND.n1260 585
R2464 GND.n4081 GND.n4080 585
R2465 GND.n4082 GND.n4081 585
R2466 GND.n1259 GND.n1258 585
R2467 GND.n4083 GND.n1259 585
R2468 GND.n4086 GND.n4085 585
R2469 GND.n4085 GND.n4084 585
R2470 GND.n4087 GND.n1253 585
R2471 GND.n1253 GND.n1252 585
R2472 GND.n4089 GND.n4088 585
R2473 GND.n4090 GND.n4089 585
R2474 GND.n1251 GND.n1250 585
R2475 GND.n4091 GND.n1251 585
R2476 GND.n4094 GND.n4093 585
R2477 GND.n4093 GND.n4092 585
R2478 GND.n4095 GND.n1245 585
R2479 GND.n1245 GND.n1244 585
R2480 GND.n4097 GND.n4096 585
R2481 GND.n4098 GND.n4097 585
R2482 GND.n1243 GND.n1242 585
R2483 GND.n4099 GND.n1243 585
R2484 GND.n4102 GND.n4101 585
R2485 GND.n4101 GND.n4100 585
R2486 GND.n4103 GND.n1237 585
R2487 GND.n1237 GND.n1236 585
R2488 GND.n4105 GND.n4104 585
R2489 GND.n4106 GND.n4105 585
R2490 GND.n1235 GND.n1234 585
R2491 GND.n4107 GND.n1235 585
R2492 GND.n4110 GND.n4109 585
R2493 GND.n4109 GND.n4108 585
R2494 GND.n4111 GND.n1229 585
R2495 GND.n1229 GND.n1228 585
R2496 GND.n4113 GND.n4112 585
R2497 GND.n4114 GND.n4113 585
R2498 GND.n1227 GND.n1226 585
R2499 GND.n4115 GND.n1227 585
R2500 GND.n4118 GND.n4117 585
R2501 GND.n4117 GND.n4116 585
R2502 GND.n4119 GND.n1221 585
R2503 GND.n1221 GND.n1220 585
R2504 GND.n4121 GND.n4120 585
R2505 GND.n4122 GND.n4121 585
R2506 GND.n1219 GND.n1218 585
R2507 GND.n4123 GND.n1219 585
R2508 GND.n4126 GND.n4125 585
R2509 GND.n4125 GND.n4124 585
R2510 GND.n4127 GND.n1213 585
R2511 GND.n1213 GND.n1212 585
R2512 GND.n4129 GND.n4128 585
R2513 GND.n4130 GND.n4129 585
R2514 GND.n1211 GND.n1210 585
R2515 GND.n4131 GND.n1211 585
R2516 GND.n4134 GND.n4133 585
R2517 GND.n4133 GND.n4132 585
R2518 GND.n4135 GND.n1205 585
R2519 GND.n1205 GND.n1204 585
R2520 GND.n4137 GND.n4136 585
R2521 GND.n4138 GND.n4137 585
R2522 GND.n1203 GND.n1202 585
R2523 GND.n4139 GND.n1203 585
R2524 GND.n4142 GND.n4141 585
R2525 GND.n4141 GND.n4140 585
R2526 GND.n4143 GND.n1197 585
R2527 GND.n1197 GND.n1196 585
R2528 GND.n4145 GND.n4144 585
R2529 GND.n4146 GND.n4145 585
R2530 GND.n1195 GND.n1194 585
R2531 GND.n4147 GND.n1195 585
R2532 GND.n4150 GND.n4149 585
R2533 GND.n4149 GND.n4148 585
R2534 GND.n4151 GND.n1189 585
R2535 GND.n1189 GND.n1188 585
R2536 GND.n4153 GND.n4152 585
R2537 GND.n4154 GND.n4153 585
R2538 GND.n1187 GND.n1186 585
R2539 GND.n4155 GND.n1187 585
R2540 GND.n4158 GND.n4157 585
R2541 GND.n4157 GND.n4156 585
R2542 GND.n4159 GND.n1181 585
R2543 GND.n1181 GND.n1180 585
R2544 GND.n4161 GND.n4160 585
R2545 GND.n4162 GND.n4161 585
R2546 GND.n1179 GND.n1178 585
R2547 GND.n4163 GND.n1179 585
R2548 GND.n4166 GND.n4165 585
R2549 GND.n4165 GND.n4164 585
R2550 GND.n4167 GND.n1173 585
R2551 GND.n1173 GND.n1172 585
R2552 GND.n4169 GND.n4168 585
R2553 GND.n4170 GND.n4169 585
R2554 GND.n1171 GND.n1170 585
R2555 GND.n4171 GND.n1171 585
R2556 GND.n4174 GND.n4173 585
R2557 GND.n4173 GND.n4172 585
R2558 GND.n4175 GND.n1165 585
R2559 GND.n1165 GND.n1164 585
R2560 GND.n4177 GND.n4176 585
R2561 GND.n4178 GND.n4177 585
R2562 GND.n1163 GND.n1162 585
R2563 GND.n4179 GND.n1163 585
R2564 GND.n4182 GND.n4181 585
R2565 GND.n4181 GND.n4180 585
R2566 GND.n4183 GND.n1157 585
R2567 GND.n1157 GND.n1156 585
R2568 GND.n4185 GND.n4184 585
R2569 GND.n4186 GND.n4185 585
R2570 GND.n1155 GND.n1154 585
R2571 GND.n4187 GND.n1155 585
R2572 GND.n4190 GND.n4189 585
R2573 GND.n4189 GND.n4188 585
R2574 GND.n4191 GND.n1149 585
R2575 GND.n1149 GND.n1148 585
R2576 GND.n4193 GND.n4192 585
R2577 GND.n4194 GND.n4193 585
R2578 GND.n1147 GND.n1146 585
R2579 GND.n4195 GND.n1147 585
R2580 GND.n4198 GND.n4197 585
R2581 GND.n4197 GND.n4196 585
R2582 GND.n4199 GND.n1141 585
R2583 GND.n1141 GND.n1140 585
R2584 GND.n4201 GND.n4200 585
R2585 GND.n4202 GND.n4201 585
R2586 GND.n2537 GND.n2536 585
R2587 GND.n2536 GND.n1348 585
R2588 GND.n2732 GND.n2731 585
R2589 GND.n2734 GND.n2535 585
R2590 GND.n2737 GND.n2736 585
R2591 GND.n2533 GND.n2532 585
R2592 GND.n2742 GND.n2741 585
R2593 GND.n2744 GND.n2531 585
R2594 GND.n2747 GND.n2746 585
R2595 GND.n2529 GND.n2528 585
R2596 GND.n2752 GND.n2751 585
R2597 GND.n2754 GND.n2527 585
R2598 GND.n2756 GND.n2755 585
R2599 GND.n2755 GND.n1348 585
R2600 GND.n1415 GND.n1414 585
R2601 GND.n3950 GND.n1415 585
R2602 GND.n2838 GND.n1407 585
R2603 GND.n2839 GND.n2838 585
R2604 GND.n2837 GND.n1406 585
R2605 GND.n2837 GND.n2836 585
R2606 GND.n2382 GND.n1405 585
R2607 GND.n2816 GND.n2382 585
R2608 GND.n2827 GND.n2826 585
R2609 GND.n2828 GND.n2827 585
R2610 GND.n2825 GND.n1399 585
R2611 GND.n2825 GND.n2824 585
R2612 GND.n2393 GND.n1398 585
R2613 GND.n2406 GND.n2393 585
R2614 GND.n2403 GND.n1397 585
R2615 GND.n2810 GND.n2403 585
R2616 GND.n2799 GND.n2797 585
R2617 GND.n2799 GND.n2798 585
R2618 GND.n2800 GND.n1391 585
R2619 GND.n2801 GND.n2800 585
R2620 GND.n2796 GND.n1390 585
R2621 GND.n2796 GND.n2795 585
R2622 GND.n2413 GND.n1389 585
R2623 GND.n2427 GND.n2413 585
R2624 GND.n2425 GND.n2424 585
R2625 GND.n2785 GND.n2425 585
R2626 GND.n2774 GND.n1383 585
R2627 GND.n2774 GND.n2773 585
R2628 GND.n2775 GND.n1382 585
R2629 GND.n2776 GND.n2775 585
R2630 GND.n2772 GND.n1381 585
R2631 GND.n2772 GND.n2771 585
R2632 GND.n1374 GND.n1372 585
R2633 GND.n2518 GND.n1372 585
R2634 GND.n3980 GND.n3979 585
R2635 GND.n3981 GND.n3980 585
R2636 GND.n1373 GND.n1371 585
R2637 GND.n2761 GND.n1371 585
R2638 GND.n2725 GND.n1360 585
R2639 GND.n3987 GND.n1360 585
R2640 GND.n2847 GND.n2846 585
R2641 GND.n2849 GND.n2375 585
R2642 GND.n2850 GND.n2374 585
R2643 GND.n2372 GND.n2370 585
R2644 GND.n2854 GND.n2369 585
R2645 GND.n2855 GND.n2367 585
R2646 GND.n2856 GND.n2366 585
R2647 GND.n2364 GND.n2361 585
R2648 GND.n2363 GND.n1539 585
R2649 GND.n3856 GND.n1538 585
R2650 GND.n3857 GND.n1537 585
R2651 GND.n1535 GND.n1534 585
R2652 GND.n2842 GND.n1412 585
R2653 GND.n3950 GND.n1412 585
R2654 GND.n2841 GND.n2840 585
R2655 GND.n2840 GND.n2839 585
R2656 GND.n2380 GND.n2379 585
R2657 GND.n2836 GND.n2380 585
R2658 GND.n2818 GND.n2817 585
R2659 GND.n2817 GND.n2816 585
R2660 GND.n2397 GND.n2391 585
R2661 GND.n2828 GND.n2391 585
R2662 GND.n2823 GND.n2822 585
R2663 GND.n2824 GND.n2823 585
R2664 GND.n2396 GND.n2395 585
R2665 GND.n2406 GND.n2395 585
R2666 GND.n2812 GND.n2811 585
R2667 GND.n2811 GND.n2810 585
R2668 GND.n2400 GND.n2399 585
R2669 GND.n2798 GND.n2400 585
R2670 GND.n2418 GND.n2411 585
R2671 GND.n2801 GND.n2411 585
R2672 GND.n2794 GND.n2793 585
R2673 GND.n2795 GND.n2794 585
R2674 GND.n2417 GND.n2416 585
R2675 GND.n2427 GND.n2416 585
R2676 GND.n2787 GND.n2786 585
R2677 GND.n2786 GND.n2785 585
R2678 GND.n2421 GND.n2420 585
R2679 GND.n2773 GND.n2421 585
R2680 GND.n2521 GND.n2435 585
R2681 GND.n2776 GND.n2435 585
R2682 GND.n2770 GND.n2769 585
R2683 GND.n2771 GND.n2770 585
R2684 GND.n2520 GND.n2519 585
R2685 GND.n2519 GND.n2518 585
R2686 GND.n2764 GND.n1370 585
R2687 GND.n3981 GND.n1370 585
R2688 GND.n2763 GND.n2762 585
R2689 GND.n2762 GND.n2761 585
R2690 GND.n2759 GND.n1358 585
R2691 GND.n3987 GND.n1358 585
R2692 GND.n3576 GND.n1859 569.379
R2693 GND.n2055 GND.n1860 569.379
R2694 GND.n3714 GND.n1604 569.379
R2695 GND.n3788 GND.n1608 569.379
R2696 GND.n4315 GND.n4314 545.866
R2697 GND.n5117 GND.n544 301.784
R2698 GND.n5125 GND.n544 301.784
R2699 GND.n5126 GND.n5125 301.784
R2700 GND.n5127 GND.n5126 301.784
R2701 GND.n5127 GND.n538 301.784
R2702 GND.n5135 GND.n538 301.784
R2703 GND.n5136 GND.n5135 301.784
R2704 GND.n5137 GND.n5136 301.784
R2705 GND.n5137 GND.n532 301.784
R2706 GND.n5145 GND.n532 301.784
R2707 GND.n5146 GND.n5145 301.784
R2708 GND.n5147 GND.n5146 301.784
R2709 GND.n5147 GND.n526 301.784
R2710 GND.n5155 GND.n526 301.784
R2711 GND.n5156 GND.n5155 301.784
R2712 GND.n5157 GND.n5156 301.784
R2713 GND.n5157 GND.n520 301.784
R2714 GND.n5165 GND.n520 301.784
R2715 GND.n5166 GND.n5165 301.784
R2716 GND.n5167 GND.n5166 301.784
R2717 GND.n5167 GND.n514 301.784
R2718 GND.n5175 GND.n514 301.784
R2719 GND.n5176 GND.n5175 301.784
R2720 GND.n5177 GND.n5176 301.784
R2721 GND.n5177 GND.n508 301.784
R2722 GND.n5185 GND.n508 301.784
R2723 GND.n5186 GND.n5185 301.784
R2724 GND.n5187 GND.n5186 301.784
R2725 GND.n5187 GND.n502 301.784
R2726 GND.n5195 GND.n502 301.784
R2727 GND.n5196 GND.n5195 301.784
R2728 GND.n5197 GND.n5196 301.784
R2729 GND.n5197 GND.n496 301.784
R2730 GND.n5205 GND.n496 301.784
R2731 GND.n5206 GND.n5205 301.784
R2732 GND.n5207 GND.n5206 301.784
R2733 GND.n5207 GND.n490 301.784
R2734 GND.n5215 GND.n490 301.784
R2735 GND.n5216 GND.n5215 301.784
R2736 GND.n5217 GND.n5216 301.784
R2737 GND.n5217 GND.n484 301.784
R2738 GND.n5225 GND.n484 301.784
R2739 GND.n5226 GND.n5225 301.784
R2740 GND.n5227 GND.n5226 301.784
R2741 GND.n5227 GND.n478 301.784
R2742 GND.n5235 GND.n478 301.784
R2743 GND.n5236 GND.n5235 301.784
R2744 GND.n5237 GND.n5236 301.784
R2745 GND.n5237 GND.n472 301.784
R2746 GND.n5245 GND.n472 301.784
R2747 GND.n5246 GND.n5245 301.784
R2748 GND.n5247 GND.n5246 301.784
R2749 GND.n5247 GND.n466 301.784
R2750 GND.n5257 GND.n466 301.784
R2751 GND.n4316 GND.n4315 280.613
R2752 GND.n4316 GND.n1023 280.613
R2753 GND.n4324 GND.n1023 280.613
R2754 GND.n4325 GND.n4324 280.613
R2755 GND.n4326 GND.n4325 280.613
R2756 GND.n4326 GND.n1017 280.613
R2757 GND.n4334 GND.n1017 280.613
R2758 GND.n4335 GND.n4334 280.613
R2759 GND.n4336 GND.n4335 280.613
R2760 GND.n4336 GND.n1011 280.613
R2761 GND.n4344 GND.n1011 280.613
R2762 GND.n4345 GND.n4344 280.613
R2763 GND.n4346 GND.n4345 280.613
R2764 GND.n4346 GND.n1005 280.613
R2765 GND.n4354 GND.n1005 280.613
R2766 GND.n4355 GND.n4354 280.613
R2767 GND.n4356 GND.n4355 280.613
R2768 GND.n4356 GND.n999 280.613
R2769 GND.n4364 GND.n999 280.613
R2770 GND.n4365 GND.n4364 280.613
R2771 GND.n4366 GND.n4365 280.613
R2772 GND.n4366 GND.n993 280.613
R2773 GND.n4374 GND.n993 280.613
R2774 GND.n4375 GND.n4374 280.613
R2775 GND.n4376 GND.n4375 280.613
R2776 GND.n4376 GND.n987 280.613
R2777 GND.n4384 GND.n987 280.613
R2778 GND.n4385 GND.n4384 280.613
R2779 GND.n4386 GND.n4385 280.613
R2780 GND.n4386 GND.n981 280.613
R2781 GND.n4394 GND.n981 280.613
R2782 GND.n4395 GND.n4394 280.613
R2783 GND.n4396 GND.n4395 280.613
R2784 GND.n4396 GND.n975 280.613
R2785 GND.n4404 GND.n975 280.613
R2786 GND.n4405 GND.n4404 280.613
R2787 GND.n4406 GND.n4405 280.613
R2788 GND.n4406 GND.n969 280.613
R2789 GND.n4414 GND.n969 280.613
R2790 GND.n4415 GND.n4414 280.613
R2791 GND.n4416 GND.n4415 280.613
R2792 GND.n4416 GND.n963 280.613
R2793 GND.n4424 GND.n963 280.613
R2794 GND.n4425 GND.n4424 280.613
R2795 GND.n4426 GND.n4425 280.613
R2796 GND.n4426 GND.n957 280.613
R2797 GND.n4434 GND.n957 280.613
R2798 GND.n4435 GND.n4434 280.613
R2799 GND.n4436 GND.n4435 280.613
R2800 GND.n4436 GND.n951 280.613
R2801 GND.n4444 GND.n951 280.613
R2802 GND.n4445 GND.n4444 280.613
R2803 GND.n4446 GND.n4445 280.613
R2804 GND.n4446 GND.n945 280.613
R2805 GND.n4454 GND.n945 280.613
R2806 GND.n4455 GND.n4454 280.613
R2807 GND.n4456 GND.n4455 280.613
R2808 GND.n4456 GND.n939 280.613
R2809 GND.n4464 GND.n939 280.613
R2810 GND.n4465 GND.n4464 280.613
R2811 GND.n4466 GND.n4465 280.613
R2812 GND.n4466 GND.n933 280.613
R2813 GND.n4474 GND.n933 280.613
R2814 GND.n4475 GND.n4474 280.613
R2815 GND.n4476 GND.n4475 280.613
R2816 GND.n4476 GND.n927 280.613
R2817 GND.n4484 GND.n927 280.613
R2818 GND.n4485 GND.n4484 280.613
R2819 GND.n4486 GND.n4485 280.613
R2820 GND.n4486 GND.n921 280.613
R2821 GND.n4494 GND.n921 280.613
R2822 GND.n4495 GND.n4494 280.613
R2823 GND.n4496 GND.n4495 280.613
R2824 GND.n4496 GND.n915 280.613
R2825 GND.n4504 GND.n915 280.613
R2826 GND.n4505 GND.n4504 280.613
R2827 GND.n4506 GND.n4505 280.613
R2828 GND.n4506 GND.n909 280.613
R2829 GND.n4514 GND.n909 280.613
R2830 GND.n4515 GND.n4514 280.613
R2831 GND.n4516 GND.n4515 280.613
R2832 GND.n4516 GND.n903 280.613
R2833 GND.n4524 GND.n903 280.613
R2834 GND.n4525 GND.n4524 280.613
R2835 GND.n4526 GND.n4525 280.613
R2836 GND.n4526 GND.n897 280.613
R2837 GND.n4534 GND.n897 280.613
R2838 GND.n4535 GND.n4534 280.613
R2839 GND.n4536 GND.n4535 280.613
R2840 GND.n4536 GND.n891 280.613
R2841 GND.n4544 GND.n891 280.613
R2842 GND.n4545 GND.n4544 280.613
R2843 GND.n4546 GND.n4545 280.613
R2844 GND.n4546 GND.n885 280.613
R2845 GND.n4554 GND.n885 280.613
R2846 GND.n4555 GND.n4554 280.613
R2847 GND.n4556 GND.n4555 280.613
R2848 GND.n4556 GND.n879 280.613
R2849 GND.n4564 GND.n879 280.613
R2850 GND.n4565 GND.n4564 280.613
R2851 GND.n4566 GND.n4565 280.613
R2852 GND.n4566 GND.n873 280.613
R2853 GND.n4574 GND.n873 280.613
R2854 GND.n4575 GND.n4574 280.613
R2855 GND.n4576 GND.n4575 280.613
R2856 GND.n4576 GND.n867 280.613
R2857 GND.n4584 GND.n867 280.613
R2858 GND.n4585 GND.n4584 280.613
R2859 GND.n4586 GND.n4585 280.613
R2860 GND.n4586 GND.n861 280.613
R2861 GND.n4594 GND.n861 280.613
R2862 GND.n4595 GND.n4594 280.613
R2863 GND.n4596 GND.n4595 280.613
R2864 GND.n4596 GND.n855 280.613
R2865 GND.n4604 GND.n855 280.613
R2866 GND.n4605 GND.n4604 280.613
R2867 GND.n4606 GND.n4605 280.613
R2868 GND.n4606 GND.n849 280.613
R2869 GND.n4614 GND.n849 280.613
R2870 GND.n4615 GND.n4614 280.613
R2871 GND.n4616 GND.n4615 280.613
R2872 GND.n4616 GND.n843 280.613
R2873 GND.n4624 GND.n843 280.613
R2874 GND.n4625 GND.n4624 280.613
R2875 GND.n4626 GND.n4625 280.613
R2876 GND.n4626 GND.n837 280.613
R2877 GND.n4634 GND.n837 280.613
R2878 GND.n4635 GND.n4634 280.613
R2879 GND.n4636 GND.n4635 280.613
R2880 GND.n4636 GND.n831 280.613
R2881 GND.n4644 GND.n831 280.613
R2882 GND.n4645 GND.n4644 280.613
R2883 GND.n4646 GND.n4645 280.613
R2884 GND.n4646 GND.n825 280.613
R2885 GND.n4654 GND.n825 280.613
R2886 GND.n4655 GND.n4654 280.613
R2887 GND.n4656 GND.n4655 280.613
R2888 GND.n4656 GND.n819 280.613
R2889 GND.n4664 GND.n819 280.613
R2890 GND.n4665 GND.n4664 280.613
R2891 GND.n4666 GND.n4665 280.613
R2892 GND.n4666 GND.n813 280.613
R2893 GND.n4674 GND.n813 280.613
R2894 GND.n4675 GND.n4674 280.613
R2895 GND.n4676 GND.n4675 280.613
R2896 GND.n4676 GND.n807 280.613
R2897 GND.n4684 GND.n807 280.613
R2898 GND.n4685 GND.n4684 280.613
R2899 GND.n4686 GND.n4685 280.613
R2900 GND.n4686 GND.n801 280.613
R2901 GND.n4694 GND.n801 280.613
R2902 GND.n4695 GND.n4694 280.613
R2903 GND.n4696 GND.n4695 280.613
R2904 GND.n4696 GND.n795 280.613
R2905 GND.n4704 GND.n795 280.613
R2906 GND.n4705 GND.n4704 280.613
R2907 GND.n4706 GND.n4705 280.613
R2908 GND.n4706 GND.n789 280.613
R2909 GND.n4714 GND.n789 280.613
R2910 GND.n4715 GND.n4714 280.613
R2911 GND.n4716 GND.n4715 280.613
R2912 GND.n4716 GND.n783 280.613
R2913 GND.n4724 GND.n783 280.613
R2914 GND.n4725 GND.n4724 280.613
R2915 GND.n4726 GND.n4725 280.613
R2916 GND.n4726 GND.n777 280.613
R2917 GND.n4734 GND.n777 280.613
R2918 GND.n4735 GND.n4734 280.613
R2919 GND.n4736 GND.n4735 280.613
R2920 GND.n4736 GND.n771 280.613
R2921 GND.n4744 GND.n771 280.613
R2922 GND.n4745 GND.n4744 280.613
R2923 GND.n4746 GND.n4745 280.613
R2924 GND.n4746 GND.n765 280.613
R2925 GND.n4754 GND.n765 280.613
R2926 GND.n4755 GND.n4754 280.613
R2927 GND.n4756 GND.n4755 280.613
R2928 GND.n4756 GND.n759 280.613
R2929 GND.n4764 GND.n759 280.613
R2930 GND.n4765 GND.n4764 280.613
R2931 GND.n4766 GND.n4765 280.613
R2932 GND.n4766 GND.n753 280.613
R2933 GND.n4774 GND.n753 280.613
R2934 GND.n4775 GND.n4774 280.613
R2935 GND.n4776 GND.n4775 280.613
R2936 GND.n4776 GND.n747 280.613
R2937 GND.n4784 GND.n747 280.613
R2938 GND.n4785 GND.n4784 280.613
R2939 GND.n4786 GND.n4785 280.613
R2940 GND.n4786 GND.n741 280.613
R2941 GND.n4794 GND.n741 280.613
R2942 GND.n4795 GND.n4794 280.613
R2943 GND.n4796 GND.n4795 280.613
R2944 GND.n4796 GND.n735 280.613
R2945 GND.n4804 GND.n735 280.613
R2946 GND.n4805 GND.n4804 280.613
R2947 GND.n4806 GND.n4805 280.613
R2948 GND.n4806 GND.n729 280.613
R2949 GND.n4814 GND.n729 280.613
R2950 GND.n4815 GND.n4814 280.613
R2951 GND.n4816 GND.n4815 280.613
R2952 GND.n4816 GND.n723 280.613
R2953 GND.n4824 GND.n723 280.613
R2954 GND.n4825 GND.n4824 280.613
R2955 GND.n4826 GND.n4825 280.613
R2956 GND.n4826 GND.n717 280.613
R2957 GND.n4834 GND.n717 280.613
R2958 GND.n4835 GND.n4834 280.613
R2959 GND.n4836 GND.n4835 280.613
R2960 GND.n4836 GND.n711 280.613
R2961 GND.n4844 GND.n711 280.613
R2962 GND.n4845 GND.n4844 280.613
R2963 GND.n4846 GND.n4845 280.613
R2964 GND.n4846 GND.n705 280.613
R2965 GND.n4854 GND.n705 280.613
R2966 GND.n4855 GND.n4854 280.613
R2967 GND.n4856 GND.n4855 280.613
R2968 GND.n4856 GND.n699 280.613
R2969 GND.n4864 GND.n699 280.613
R2970 GND.n4865 GND.n4864 280.613
R2971 GND.n4866 GND.n4865 280.613
R2972 GND.n4866 GND.n693 280.613
R2973 GND.n4874 GND.n693 280.613
R2974 GND.n4875 GND.n4874 280.613
R2975 GND.n4876 GND.n4875 280.613
R2976 GND.n4876 GND.n687 280.613
R2977 GND.n4884 GND.n687 280.613
R2978 GND.n4885 GND.n4884 280.613
R2979 GND.n4886 GND.n4885 280.613
R2980 GND.n4886 GND.n681 280.613
R2981 GND.n4894 GND.n681 280.613
R2982 GND.n4895 GND.n4894 280.613
R2983 GND.n4896 GND.n4895 280.613
R2984 GND.n4896 GND.n675 280.613
R2985 GND.n4904 GND.n675 280.613
R2986 GND.n4905 GND.n4904 280.613
R2987 GND.n4906 GND.n4905 280.613
R2988 GND.n4906 GND.n669 280.613
R2989 GND.n4914 GND.n669 280.613
R2990 GND.n4915 GND.n4914 280.613
R2991 GND.n4916 GND.n4915 280.613
R2992 GND.n4916 GND.n663 280.613
R2993 GND.n4924 GND.n663 280.613
R2994 GND.n4925 GND.n4924 280.613
R2995 GND.n4926 GND.n4925 280.613
R2996 GND.n4926 GND.n657 280.613
R2997 GND.n4934 GND.n657 280.613
R2998 GND.n4935 GND.n4934 280.613
R2999 GND.n4936 GND.n4935 280.613
R3000 GND.n4936 GND.n651 280.613
R3001 GND.n4944 GND.n651 280.613
R3002 GND.n4945 GND.n4944 280.613
R3003 GND.n4946 GND.n4945 280.613
R3004 GND.n4946 GND.n645 280.613
R3005 GND.n4954 GND.n645 280.613
R3006 GND.n4955 GND.n4954 280.613
R3007 GND.n4956 GND.n4955 280.613
R3008 GND.n4956 GND.n639 280.613
R3009 GND.n4964 GND.n639 280.613
R3010 GND.n4965 GND.n4964 280.613
R3011 GND.n4966 GND.n4965 280.613
R3012 GND.n4966 GND.n633 280.613
R3013 GND.n4974 GND.n633 280.613
R3014 GND.n4975 GND.n4974 280.613
R3015 GND.n4976 GND.n4975 280.613
R3016 GND.n4976 GND.n627 280.613
R3017 GND.n4984 GND.n627 280.613
R3018 GND.n4985 GND.n4984 280.613
R3019 GND.n4986 GND.n4985 280.613
R3020 GND.n4986 GND.n621 280.613
R3021 GND.n4994 GND.n621 280.613
R3022 GND.n4995 GND.n4994 280.613
R3023 GND.n4996 GND.n4995 280.613
R3024 GND.n4996 GND.n615 280.613
R3025 GND.n5004 GND.n615 280.613
R3026 GND.n5005 GND.n5004 280.613
R3027 GND.n5006 GND.n5005 280.613
R3028 GND.n5006 GND.n609 280.613
R3029 GND.n5014 GND.n609 280.613
R3030 GND.n5015 GND.n5014 280.613
R3031 GND.n5016 GND.n5015 280.613
R3032 GND.n5016 GND.n603 280.613
R3033 GND.n5024 GND.n603 280.613
R3034 GND.n5025 GND.n5024 280.613
R3035 GND.n5026 GND.n5025 280.613
R3036 GND.n5026 GND.n597 280.613
R3037 GND.n5034 GND.n597 280.613
R3038 GND.n5035 GND.n5034 280.613
R3039 GND.n5036 GND.n5035 280.613
R3040 GND.n5036 GND.n591 280.613
R3041 GND.n5044 GND.n591 280.613
R3042 GND.n5045 GND.n5044 280.613
R3043 GND.n5046 GND.n5045 280.613
R3044 GND.n5046 GND.n585 280.613
R3045 GND.n5054 GND.n585 280.613
R3046 GND.n5055 GND.n5054 280.613
R3047 GND.n5056 GND.n5055 280.613
R3048 GND.n5056 GND.n579 280.613
R3049 GND.n5064 GND.n579 280.613
R3050 GND.n5065 GND.n5064 280.613
R3051 GND.n5066 GND.n5065 280.613
R3052 GND.n5066 GND.n573 280.613
R3053 GND.n5074 GND.n573 280.613
R3054 GND.n5075 GND.n5074 280.613
R3055 GND.n5076 GND.n5075 280.613
R3056 GND.n5076 GND.n567 280.613
R3057 GND.n5084 GND.n567 280.613
R3058 GND.n5085 GND.n5084 280.613
R3059 GND.n5086 GND.n5085 280.613
R3060 GND.n5086 GND.n561 280.613
R3061 GND.n5094 GND.n561 280.613
R3062 GND.n5095 GND.n5094 280.613
R3063 GND.n5096 GND.n5095 280.613
R3064 GND.n5096 GND.n555 280.613
R3065 GND.n5104 GND.n555 280.613
R3066 GND.n5105 GND.n5104 280.613
R3067 GND.n5106 GND.n5105 280.613
R3068 GND.n5106 GND.n549 280.613
R3069 GND.n5115 GND.n549 280.613
R3070 GND.n5116 GND.n5115 280.613
R3071 GND.n5258 GND.n5257 279.082
R3072 GND.n3790 GND.n3789 256.663
R3073 GND.n3790 GND.n1587 256.663
R3074 GND.n3790 GND.n1588 256.663
R3075 GND.n3790 GND.n1589 256.663
R3076 GND.n3790 GND.n1590 256.663
R3077 GND.n3790 GND.n1591 256.663
R3078 GND.n3790 GND.n1592 256.663
R3079 GND.n3790 GND.n1593 256.663
R3080 GND.n3790 GND.n1594 256.663
R3081 GND.n3753 GND.n3752 256.663
R3082 GND.n3790 GND.n1595 256.663
R3083 GND.n3790 GND.n1596 256.663
R3084 GND.n3790 GND.n1597 256.663
R3085 GND.n3790 GND.n1598 256.663
R3086 GND.n3790 GND.n1599 256.663
R3087 GND.n3790 GND.n1600 256.663
R3088 GND.n3790 GND.n1601 256.663
R3089 GND.n3790 GND.n1602 256.663
R3090 GND.n3790 GND.n1603 256.663
R3091 GND.n2102 GND.n2056 256.663
R3092 GND.n2102 GND.n2017 256.663
R3093 GND.n2102 GND.n2016 256.663
R3094 GND.n2102 GND.n2015 256.663
R3095 GND.n2102 GND.n2014 256.663
R3096 GND.n2102 GND.n2013 256.663
R3097 GND.n2102 GND.n2012 256.663
R3098 GND.n2102 GND.n2011 256.663
R3099 GND.n2102 GND.n2010 256.663
R3100 GND.n2105 GND.n2104 256.663
R3101 GND.n2102 GND.n2007 256.663
R3102 GND.n2102 GND.n2057 256.663
R3103 GND.n2102 GND.n2058 256.663
R3104 GND.n2102 GND.n2059 256.663
R3105 GND.n2102 GND.n2060 256.663
R3106 GND.n2102 GND.n2061 256.663
R3107 GND.n2102 GND.n2062 256.663
R3108 GND.n2102 GND.n2063 256.663
R3109 GND.n2102 GND.n2101 256.663
R3110 GND.n2376 GND.t115 256.274
R3111 GND.n1433 GND.t28 256.274
R3112 GND.n1491 GND.t97 256.274
R3113 GND.n1520 GND.t15 256.274
R3114 GND.n1450 GND.t112 256.274
R3115 GND.n1991 GND.t100 256.274
R3116 GND.n2108 GND.t124 256.274
R3117 GND.n2124 GND.t31 256.274
R3118 GND.n2139 GND.t78 256.274
R3119 GND.n150 GND.t109 256.274
R3120 GND.n135 GND.t59 256.274
R3121 GND.n206 GND.t51 256.274
R3122 GND.n106 GND.t118 256.274
R3123 GND.n3277 GND.t81 256.274
R3124 GND.n2249 GND.t45 256.274
R3125 GND.n2584 GND.t94 256.274
R3126 GND.n2567 GND.t11 256.274
R3127 GND.n2686 GND.t25 256.274
R3128 GND.n2539 GND.t19 256.274
R3129 GND.n2524 GND.t127 256.274
R3130 GND.n1931 GND.t87 249.743
R3131 GND.n3862 GND.t38 249.743
R3132 GND.n3500 GND.n1970 242.672
R3133 GND.n3500 GND.n1971 242.672
R3134 GND.n3500 GND.n1972 242.672
R3135 GND.n3500 GND.n1973 242.672
R3136 GND.n3500 GND.n1974 242.672
R3137 GND.n3500 GND.n1975 242.672
R3138 GND.n3317 GND.n258 242.672
R3139 GND.n3307 GND.n258 242.672
R3140 GND.n3306 GND.n258 242.672
R3141 GND.n3284 GND.n258 242.672
R3142 GND.n3296 GND.n258 242.672
R3143 GND.n3288 GND.n258 242.672
R3144 GND.n3850 GND.n3849 242.672
R3145 GND.n3850 GND.n1544 242.672
R3146 GND.n3850 GND.n1545 242.672
R3147 GND.n3850 GND.n1546 242.672
R3148 GND.n3850 GND.n1547 242.672
R3149 GND.n3850 GND.n1548 242.672
R3150 GND.n3850 GND.n1549 242.672
R3151 GND.n3850 GND.n1550 242.672
R3152 GND.n3851 GND.n3850 242.672
R3153 GND.n3545 GND.n1909 242.672
R3154 GND.n3545 GND.n1910 242.672
R3155 GND.n3545 GND.n1911 242.672
R3156 GND.n3545 GND.n1912 242.672
R3157 GND.n3545 GND.n1913 242.672
R3158 GND.n3545 GND.n1914 242.672
R3159 GND.n3545 GND.n1915 242.672
R3160 GND.n3545 GND.n1916 242.672
R3161 GND.n3545 GND.n3544 242.672
R3162 GND.n2597 GND.n1348 242.672
R3163 GND.n2599 GND.n1348 242.672
R3164 GND.n2607 GND.n1348 242.672
R3165 GND.n2609 GND.n1348 242.672
R3166 GND.n2617 GND.n1348 242.672
R3167 GND.n2619 GND.n1348 242.672
R3168 GND.n2627 GND.n1348 242.672
R3169 GND.n2629 GND.n1348 242.672
R3170 GND.n2637 GND.n1348 242.672
R3171 GND.n2639 GND.n1348 242.672
R3172 GND.n2648 GND.n1348 242.672
R3173 GND.n2650 GND.n1348 242.672
R3174 GND.n2658 GND.n1348 242.672
R3175 GND.n2660 GND.n1348 242.672
R3176 GND.n2668 GND.n1348 242.672
R3177 GND.n2670 GND.n1348 242.672
R3178 GND.n2678 GND.n1348 242.672
R3179 GND.n2680 GND.n1348 242.672
R3180 GND.n2690 GND.n1348 242.672
R3181 GND.n2692 GND.n1348 242.672
R3182 GND.n2700 GND.n1348 242.672
R3183 GND.n2702 GND.n1348 242.672
R3184 GND.n2710 GND.n1348 242.672
R3185 GND.n2712 GND.n1348 242.672
R3186 GND.n2720 GND.n1348 242.672
R3187 GND.n1523 GND.n1467 242.672
R3188 GND.n1518 GND.n1467 242.672
R3189 GND.n1515 GND.n1467 242.672
R3190 GND.n1510 GND.n1467 242.672
R3191 GND.n1507 GND.n1467 242.672
R3192 GND.n1502 GND.n1467 242.672
R3193 GND.n1499 GND.n1467 242.672
R3194 GND.n1494 GND.n1467 242.672
R3195 GND.n1488 GND.n1467 242.672
R3196 GND.n1483 GND.n1467 242.672
R3197 GND.n1480 GND.n1467 242.672
R3198 GND.n1475 GND.n1467 242.672
R3199 GND.n1472 GND.n1467 242.672
R3200 GND.n3910 GND.n1467 242.672
R3201 GND.n3911 GND.n1452 242.672
R3202 GND.n3912 GND.n1467 242.672
R3203 GND.n1467 GND.n1453 242.672
R3204 GND.n1467 GND.n1455 242.672
R3205 GND.n1467 GND.n1456 242.672
R3206 GND.n1467 GND.n1458 242.672
R3207 GND.n1467 GND.n1459 242.672
R3208 GND.n1467 GND.n1460 242.672
R3209 GND.n1467 GND.n1462 242.672
R3210 GND.n1467 GND.n1463 242.672
R3211 GND.n1467 GND.n1465 242.672
R3212 GND.n1467 GND.n1466 242.672
R3213 GND.n3500 GND.n3499 242.672
R3214 GND.n3500 GND.n1946 242.672
R3215 GND.n3500 GND.n1947 242.672
R3216 GND.n3500 GND.n1948 242.672
R3217 GND.n3500 GND.n1949 242.672
R3218 GND.n3500 GND.n1950 242.672
R3219 GND.n3500 GND.n1951 242.672
R3220 GND.n3500 GND.n1952 242.672
R3221 GND.n3500 GND.n1953 242.672
R3222 GND.n3500 GND.n1954 242.672
R3223 GND.n3500 GND.n1955 242.672
R3224 GND.n3456 GND.n2106 242.672
R3225 GND.n3500 GND.n1956 242.672
R3226 GND.n3500 GND.n1957 242.672
R3227 GND.n3500 GND.n1958 242.672
R3228 GND.n3500 GND.n1959 242.672
R3229 GND.n3500 GND.n1960 242.672
R3230 GND.n3500 GND.n1961 242.672
R3231 GND.n3500 GND.n1962 242.672
R3232 GND.n3500 GND.n1963 242.672
R3233 GND.n3500 GND.n1964 242.672
R3234 GND.n3500 GND.n1965 242.672
R3235 GND.n3500 GND.n1966 242.672
R3236 GND.n3500 GND.n1967 242.672
R3237 GND.n3500 GND.n1968 242.672
R3238 GND.n3500 GND.n1969 242.672
R3239 GND.n258 GND.n70 242.672
R3240 GND.n258 GND.n71 242.672
R3241 GND.n258 GND.n72 242.672
R3242 GND.n258 GND.n73 242.672
R3243 GND.n258 GND.n74 242.672
R3244 GND.n258 GND.n75 242.672
R3245 GND.n258 GND.n76 242.672
R3246 GND.n258 GND.n77 242.672
R3247 GND.n258 GND.n78 242.672
R3248 GND.n258 GND.n79 242.672
R3249 GND.n258 GND.n80 242.672
R3250 GND.n258 GND.n81 242.672
R3251 GND.n258 GND.n82 242.672
R3252 GND.n258 GND.n83 242.672
R3253 GND.n258 GND.n84 242.672
R3254 GND.n258 GND.n85 242.672
R3255 GND.n258 GND.n86 242.672
R3256 GND.n258 GND.n87 242.672
R3257 GND.n258 GND.n88 242.672
R3258 GND.n258 GND.n89 242.672
R3259 GND.n258 GND.n90 242.672
R3260 GND.n258 GND.n91 242.672
R3261 GND.n258 GND.n92 242.672
R3262 GND.n258 GND.n93 242.672
R3263 GND.n258 GND.n94 242.672
R3264 GND.n2733 GND.n1348 242.672
R3265 GND.n2735 GND.n1348 242.672
R3266 GND.n2743 GND.n1348 242.672
R3267 GND.n2745 GND.n1348 242.672
R3268 GND.n2753 GND.n1348 242.672
R3269 GND.n2845 GND.n1467 242.672
R3270 GND.n2373 GND.n1467 242.672
R3271 GND.n2368 GND.n1467 242.672
R3272 GND.n2365 GND.n1467 242.672
R3273 GND.n2362 GND.n1467 242.672
R3274 GND.n1536 GND.n1467 242.672
R3275 GND.n1617 GND.n1615 240.849
R3276 GND.n1850 GND.n1848 240.849
R3277 GND.n257 GND.n95 240.244
R3278 GND.n250 GND.n249 240.244
R3279 GND.n247 GND.n246 240.244
R3280 GND.n243 GND.n242 240.244
R3281 GND.n239 GND.n238 240.244
R3282 GND.n235 GND.n234 240.244
R3283 GND.n231 GND.n230 240.244
R3284 GND.n227 GND.n226 240.244
R3285 GND.n223 GND.n222 240.244
R3286 GND.n219 GND.n218 240.244
R3287 GND.n215 GND.n214 240.244
R3288 GND.n211 GND.n210 240.244
R3289 GND.n204 GND.n203 240.244
R3290 GND.n200 GND.n199 240.244
R3291 GND.n196 GND.n195 240.244
R3292 GND.n192 GND.n191 240.244
R3293 GND.n188 GND.n187 240.244
R3294 GND.n184 GND.n183 240.244
R3295 GND.n138 GND.n137 240.244
R3296 GND.n176 GND.n175 240.244
R3297 GND.n172 GND.n171 240.244
R3298 GND.n168 GND.n167 240.244
R3299 GND.n164 GND.n163 240.244
R3300 GND.n160 GND.n159 240.244
R3301 GND.n156 GND.n155 240.244
R3302 GND.n3402 GND.n2144 240.244
R3303 GND.n3394 GND.n2144 240.244
R3304 GND.n3394 GND.n2155 240.244
R3305 GND.n2171 GND.n2155 240.244
R3306 GND.n3255 GND.n2171 240.244
R3307 GND.n3255 GND.n2184 240.244
R3308 GND.n2189 GND.n2184 240.244
R3309 GND.n3261 GND.n2189 240.244
R3310 GND.n3261 GND.n2222 240.244
R3311 GND.n2222 GND.n11 240.244
R3312 GND.n2230 GND.n11 240.244
R3313 GND.n3266 GND.n2230 240.244
R3314 GND.n3266 GND.n2234 240.244
R3315 GND.n2234 GND.n30 240.244
R3316 GND.n3331 GND.n30 240.244
R3317 GND.n3331 GND.n42 240.244
R3318 GND.n3327 GND.n42 240.244
R3319 GND.n3327 GND.n52 240.244
R3320 GND.n5475 GND.n52 240.244
R3321 GND.n1978 GND.n1977 240.244
R3322 GND.n3493 GND.n1977 240.244
R3323 GND.n3491 GND.n3490 240.244
R3324 GND.n3487 GND.n3486 240.244
R3325 GND.n3483 GND.n3482 240.244
R3326 GND.n3479 GND.n3478 240.244
R3327 GND.n3475 GND.n3474 240.244
R3328 GND.n3471 GND.n3470 240.244
R3329 GND.n3467 GND.n3466 240.244
R3330 GND.n3463 GND.n3462 240.244
R3331 GND.n3459 GND.n3458 240.244
R3332 GND.n3454 GND.n3453 240.244
R3333 GND.n3450 GND.n3449 240.244
R3334 GND.n3446 GND.n3445 240.244
R3335 GND.n3442 GND.n3441 240.244
R3336 GND.n3438 GND.n3437 240.244
R3337 GND.n3434 GND.n3433 240.244
R3338 GND.n3429 GND.n2122 240.244
R3339 GND.n3427 GND.n3426 240.244
R3340 GND.n3423 GND.n3422 240.244
R3341 GND.n3419 GND.n3418 240.244
R3342 GND.n3415 GND.n3414 240.244
R3343 GND.n3411 GND.n3410 240.244
R3344 GND.n2138 GND.n2137 240.244
R3345 GND.n2160 GND.n1979 240.244
R3346 GND.n3392 GND.n2160 240.244
R3347 GND.n3392 GND.n2161 240.244
R3348 GND.n3388 GND.n2161 240.244
R3349 GND.n3388 GND.n2169 240.244
R3350 GND.n3380 GND.n2169 240.244
R3351 GND.n3380 GND.n3378 240.244
R3352 GND.n3378 GND.n2188 240.244
R3353 GND.n2188 GND.n14 240.244
R3354 GND.n5499 GND.n14 240.244
R3355 GND.n5499 GND.n15 240.244
R3356 GND.n2232 GND.n15 240.244
R3357 GND.n2232 GND.n27 240.244
R3358 GND.n5494 GND.n27 240.244
R3359 GND.n5494 GND.n28 240.244
R3360 GND.n5486 GND.n28 240.244
R3361 GND.n5486 GND.n45 240.244
R3362 GND.n5482 GND.n45 240.244
R3363 GND.n5482 GND.n50 240.244
R3364 GND.n1421 GND.n1417 240.244
R3365 GND.n1464 GND.n1422 240.244
R3366 GND.n1426 GND.n1425 240.244
R3367 GND.n1461 GND.n1427 240.244
R3368 GND.n1431 GND.n1430 240.244
R3369 GND.n1437 GND.n1432 240.244
R3370 GND.n1439 GND.n1438 240.244
R3371 GND.n1457 GND.n1442 240.244
R3372 GND.n1444 GND.n1443 240.244
R3373 GND.n1454 GND.n1447 240.244
R3374 GND.n3913 GND.n1448 240.244
R3375 GND.n3909 GND.n1468 240.244
R3376 GND.n1474 GND.n1473 240.244
R3377 GND.n1479 GND.n1476 240.244
R3378 GND.n1482 GND.n1481 240.244
R3379 GND.n1487 GND.n1484 240.244
R3380 GND.n1490 GND.n1489 240.244
R3381 GND.n1496 GND.n1495 240.244
R3382 GND.n1501 GND.n1500 240.244
R3383 GND.n1504 GND.n1503 240.244
R3384 GND.n1509 GND.n1508 240.244
R3385 GND.n1512 GND.n1511 240.244
R3386 GND.n1517 GND.n1516 240.244
R3387 GND.n1524 GND.n1519 240.244
R3388 GND.n2760 GND.n1357 240.244
R3389 GND.n2760 GND.n1369 240.244
R3390 GND.n1378 GND.n1369 240.244
R3391 GND.n1379 GND.n1378 240.244
R3392 GND.n2434 GND.n1379 240.244
R3393 GND.n2434 GND.n1385 240.244
R3394 GND.n1386 GND.n1385 240.244
R3395 GND.n1387 GND.n1386 240.244
R3396 GND.n2415 GND.n1387 240.244
R3397 GND.n2415 GND.n1393 240.244
R3398 GND.n1394 GND.n1393 240.244
R3399 GND.n1395 GND.n1394 240.244
R3400 GND.n2405 GND.n1395 240.244
R3401 GND.n2405 GND.n1401 240.244
R3402 GND.n1402 GND.n1401 240.244
R3403 GND.n1403 GND.n1402 240.244
R3404 GND.n2384 GND.n1403 240.244
R3405 GND.n2384 GND.n1409 240.244
R3406 GND.n3951 GND.n1409 240.244
R3407 GND.n2600 GND.n2598 240.244
R3408 GND.n2606 GND.n2591 240.244
R3409 GND.n2610 GND.n2608 240.244
R3410 GND.n2616 GND.n2587 240.244
R3411 GND.n2620 GND.n2618 240.244
R3412 GND.n2626 GND.n2580 240.244
R3413 GND.n2630 GND.n2628 240.244
R3414 GND.n2636 GND.n2576 240.244
R3415 GND.n2640 GND.n2638 240.244
R3416 GND.n2647 GND.n2572 240.244
R3417 GND.n2651 GND.n2649 240.244
R3418 GND.n2657 GND.n2566 240.244
R3419 GND.n2661 GND.n2659 240.244
R3420 GND.n2667 GND.n2562 240.244
R3421 GND.n2671 GND.n2669 240.244
R3422 GND.n2677 GND.n2558 240.244
R3423 GND.n2681 GND.n2679 240.244
R3424 GND.n2689 GND.n2554 240.244
R3425 GND.n2693 GND.n2691 240.244
R3426 GND.n2699 GND.n2550 240.244
R3427 GND.n2703 GND.n2701 240.244
R3428 GND.n2709 GND.n2546 240.244
R3429 GND.n2713 GND.n2711 240.244
R3430 GND.n2719 GND.n2542 240.244
R3431 GND.n2722 GND.n2721 240.244
R3432 GND.n3986 GND.n1362 240.244
R3433 GND.n3982 GND.n1362 240.244
R3434 GND.n3982 GND.n1367 240.244
R3435 GND.n2432 GND.n1367 240.244
R3436 GND.n2777 GND.n2432 240.244
R3437 GND.n2777 GND.n2426 240.244
R3438 GND.n2784 GND.n2426 240.244
R3439 GND.n2784 GND.n2428 240.244
R3440 GND.n2428 GND.n2409 240.244
R3441 GND.n2802 GND.n2409 240.244
R3442 GND.n2802 GND.n2404 240.244
R3443 GND.n2809 GND.n2404 240.244
R3444 GND.n2809 GND.n2407 240.244
R3445 GND.n2407 GND.n2389 240.244
R3446 GND.n2829 GND.n2389 240.244
R3447 GND.n2829 GND.n2385 240.244
R3448 GND.n2835 GND.n2385 240.244
R3449 GND.n2835 GND.n1416 240.244
R3450 GND.n3949 GND.n1416 240.244
R3451 GND.n3546 GND.n1906 240.244
R3452 GND.n3543 GND.n1917 240.244
R3453 GND.n3539 GND.n3538 240.244
R3454 GND.n3535 GND.n3534 240.244
R3455 GND.n3531 GND.n3530 240.244
R3456 GND.n3527 GND.n3526 240.244
R3457 GND.n3523 GND.n3522 240.244
R3458 GND.n3519 GND.n3518 240.244
R3459 GND.n3515 GND.n3514 240.244
R3460 GND.n2358 GND.n1541 240.244
R3461 GND.n2358 GND.n1561 240.244
R3462 GND.n2864 GND.n1561 240.244
R3463 GND.n2864 GND.n2863 240.244
R3464 GND.n2863 GND.n1573 240.244
R3465 GND.n2871 GND.n1573 240.244
R3466 GND.n2871 GND.n1586 240.244
R3467 GND.n2352 GND.n1586 240.244
R3468 GND.n2352 GND.n1642 240.244
R3469 GND.n2912 GND.n1642 240.244
R3470 GND.n2912 GND.n1652 240.244
R3471 GND.n2347 GND.n1652 240.244
R3472 GND.n2944 GND.n2347 240.244
R3473 GND.n2944 GND.n2348 240.244
R3474 GND.n2348 GND.n1672 240.244
R3475 GND.n2939 GND.n1672 240.244
R3476 GND.n2939 GND.n1683 240.244
R3477 GND.n2936 GND.n1683 240.244
R3478 GND.n2936 GND.n2935 240.244
R3479 GND.n2935 GND.n2934 240.244
R3480 GND.n2934 GND.n2924 240.244
R3481 GND.n2924 GND.n2332 240.244
R3482 GND.n2332 GND.n2316 240.244
R3483 GND.n3049 GND.n2316 240.244
R3484 GND.n3050 GND.n3049 240.244
R3485 GND.n3050 GND.n2311 240.244
R3486 GND.n3061 GND.n2311 240.244
R3487 GND.n3061 GND.n2312 240.244
R3488 GND.n3057 GND.n2312 240.244
R3489 GND.n3057 GND.n2298 240.244
R3490 GND.n3073 GND.n2298 240.244
R3491 GND.n3073 GND.n2294 240.244
R3492 GND.n3082 GND.n2294 240.244
R3493 GND.n3082 GND.n2279 240.244
R3494 GND.n3101 GND.n2279 240.244
R3495 GND.n3102 GND.n3101 240.244
R3496 GND.n3103 GND.n3102 240.244
R3497 GND.n3103 GND.n2275 240.244
R3498 GND.n3110 GND.n2275 240.244
R3499 GND.n3110 GND.n1787 240.244
R3500 GND.n3143 GND.n1787 240.244
R3501 GND.n3143 GND.n1797 240.244
R3502 GND.n2263 GND.n1797 240.244
R3503 GND.n3150 GND.n2263 240.244
R3504 GND.n3151 GND.n3150 240.244
R3505 GND.n3152 GND.n3151 240.244
R3506 GND.n3152 GND.n2259 240.244
R3507 GND.n3182 GND.n2259 240.244
R3508 GND.n3183 GND.n3182 240.244
R3509 GND.n3184 GND.n3183 240.244
R3510 GND.n3184 GND.n1873 240.244
R3511 GND.n3188 GND.n1873 240.244
R3512 GND.n3188 GND.n1884 240.244
R3513 GND.n3196 GND.n1884 240.244
R3514 GND.n3197 GND.n3196 240.244
R3515 GND.n3197 GND.n1896 240.244
R3516 GND.n3510 GND.n1896 240.244
R3517 GND.n1553 GND.n1552 240.244
R3518 GND.n3843 GND.n1552 240.244
R3519 GND.n3841 GND.n3840 240.244
R3520 GND.n3837 GND.n3836 240.244
R3521 GND.n3833 GND.n3832 240.244
R3522 GND.n3829 GND.n3828 240.244
R3523 GND.n3825 GND.n3824 240.244
R3524 GND.n1529 GND.n1528 240.244
R3525 GND.n1542 GND.n1530 240.244
R3526 GND.n1556 GND.n1554 240.244
R3527 GND.n3806 GND.n1556 240.244
R3528 GND.n3806 GND.n1559 240.244
R3529 GND.n1575 GND.n1559 240.244
R3530 GND.n3796 GND.n1575 240.244
R3531 GND.n3796 GND.n1576 240.244
R3532 GND.n3792 GND.n1576 240.244
R3533 GND.n3792 GND.n1584 240.244
R3534 GND.n3711 GND.n1584 240.244
R3535 GND.n3711 GND.n1644 240.244
R3536 GND.n3707 GND.n1644 240.244
R3537 GND.n3707 GND.n1650 240.244
R3538 GND.n2949 GND.n1650 240.244
R3539 GND.n2949 GND.n1674 240.244
R3540 GND.n3690 GND.n1674 240.244
R3541 GND.n3690 GND.n1675 240.244
R3542 GND.n3686 GND.n1675 240.244
R3543 GND.n3686 GND.n1681 240.244
R3544 GND.n2324 GND.n1681 240.244
R3545 GND.n2330 GND.n2324 240.244
R3546 GND.n2331 GND.n2330 240.244
R3547 GND.n3036 GND.n2331 240.244
R3548 GND.n3036 GND.n2319 240.244
R3549 GND.n3047 GND.n2319 240.244
R3550 GND.n3047 GND.n2320 240.244
R3551 GND.n2320 GND.n2308 240.244
R3552 GND.n3063 GND.n2308 240.244
R3553 GND.n3064 GND.n3063 240.244
R3554 GND.n3065 GND.n3064 240.244
R3555 GND.n3065 GND.n2304 240.244
R3556 GND.n3071 GND.n2304 240.244
R3557 GND.n3071 GND.n2291 240.244
R3558 GND.n3084 GND.n2291 240.244
R3559 GND.n3084 GND.n2286 240.244
R3560 GND.n3099 GND.n2286 240.244
R3561 GND.n3099 GND.n2287 240.244
R3562 GND.n3095 GND.n2287 240.244
R3563 GND.n3095 GND.n3094 240.244
R3564 GND.n3094 GND.n1789 240.244
R3565 GND.n3606 GND.n1789 240.244
R3566 GND.n3606 GND.n1790 240.244
R3567 GND.n3602 GND.n1790 240.244
R3568 GND.n3602 GND.n1796 240.244
R3569 GND.n3169 GND.n1796 240.244
R3570 GND.n3170 GND.n3169 240.244
R3571 GND.n3171 GND.n3170 240.244
R3572 GND.n3171 GND.n3161 240.244
R3573 GND.n3180 GND.n3161 240.244
R3574 GND.n3180 GND.n3162 240.244
R3575 GND.n3162 GND.n1875 240.244
R3576 GND.n3566 GND.n1875 240.244
R3577 GND.n3566 GND.n1876 240.244
R3578 GND.n3562 GND.n1876 240.244
R3579 GND.n3562 GND.n1882 240.244
R3580 GND.n1898 GND.n1882 240.244
R3581 GND.n3552 GND.n1898 240.244
R3582 GND.n3552 GND.n1899 240.244
R3583 GND.n3295 GND.n3294 240.244
R3584 GND.n3298 GND.n3297 240.244
R3585 GND.n3305 GND.n3304 240.244
R3586 GND.n3309 GND.n3308 240.244
R3587 GND.n3316 GND.n3280 240.244
R3588 GND.n2247 GND.n2147 240.244
R3589 GND.n2247 GND.n2157 240.244
R3590 GND.n3240 GND.n2157 240.244
R3591 GND.n3240 GND.n2172 240.244
R3592 GND.n3253 GND.n2172 240.244
R3593 GND.n3253 GND.n2185 240.244
R3594 GND.n2190 GND.n2185 240.244
R3595 GND.n3248 GND.n2190 240.244
R3596 GND.n3248 GND.n9 240.244
R3597 GND.n5501 GND.n9 240.244
R3598 GND.n5501 GND.n10 240.244
R3599 GND.n2235 GND.n10 240.244
R3600 GND.n3337 GND.n2235 240.244
R3601 GND.n3337 GND.n31 240.244
R3602 GND.n3333 GND.n31 240.244
R3603 GND.n3333 GND.n43 240.244
R3604 GND.n3325 GND.n43 240.244
R3605 GND.n3325 GND.n53 240.244
R3606 GND.n60 GND.n53 240.244
R3607 GND.n3208 GND.n3207 240.244
R3608 GND.n3211 GND.n3210 240.244
R3609 GND.n3219 GND.n3218 240.244
R3610 GND.n3222 GND.n3221 240.244
R3611 GND.n3229 GND.n3228 240.244
R3612 GND.n3400 GND.n2150 240.244
R3613 GND.n2159 GND.n2150 240.244
R3614 GND.n2174 GND.n2159 240.244
R3615 GND.n3386 GND.n2174 240.244
R3616 GND.n3386 GND.n2175 240.244
R3617 GND.n3382 GND.n2175 240.244
R3618 GND.n3382 GND.n2182 240.244
R3619 GND.n2223 GND.n2182 240.244
R3620 GND.n3367 GND.n2223 240.244
R3621 GND.n3367 GND.n13 240.244
R3622 GND.n3363 GND.n13 240.244
R3623 GND.n3363 GND.n2229 240.244
R3624 GND.n2229 GND.n33 240.244
R3625 GND.n5492 GND.n33 240.244
R3626 GND.n5492 GND.n34 240.244
R3627 GND.n5488 GND.n34 240.244
R3628 GND.n5488 GND.n40 240.244
R3629 GND.n5480 GND.n40 240.244
R3630 GND.n5480 GND.n55 240.244
R3631 GND.n4317 GND.n1028 240.244
R3632 GND.n4317 GND.n1024 240.244
R3633 GND.n4323 GND.n1024 240.244
R3634 GND.n4323 GND.n1022 240.244
R3635 GND.n4327 GND.n1022 240.244
R3636 GND.n4327 GND.n1018 240.244
R3637 GND.n4333 GND.n1018 240.244
R3638 GND.n4333 GND.n1016 240.244
R3639 GND.n4337 GND.n1016 240.244
R3640 GND.n4337 GND.n1012 240.244
R3641 GND.n4343 GND.n1012 240.244
R3642 GND.n4343 GND.n1010 240.244
R3643 GND.n4347 GND.n1010 240.244
R3644 GND.n4347 GND.n1006 240.244
R3645 GND.n4353 GND.n1006 240.244
R3646 GND.n4353 GND.n1004 240.244
R3647 GND.n4357 GND.n1004 240.244
R3648 GND.n4357 GND.n1000 240.244
R3649 GND.n4363 GND.n1000 240.244
R3650 GND.n4363 GND.n998 240.244
R3651 GND.n4367 GND.n998 240.244
R3652 GND.n4367 GND.n994 240.244
R3653 GND.n4373 GND.n994 240.244
R3654 GND.n4373 GND.n992 240.244
R3655 GND.n4377 GND.n992 240.244
R3656 GND.n4377 GND.n988 240.244
R3657 GND.n4383 GND.n988 240.244
R3658 GND.n4383 GND.n986 240.244
R3659 GND.n4387 GND.n986 240.244
R3660 GND.n4387 GND.n982 240.244
R3661 GND.n4393 GND.n982 240.244
R3662 GND.n4393 GND.n980 240.244
R3663 GND.n4397 GND.n980 240.244
R3664 GND.n4397 GND.n976 240.244
R3665 GND.n4403 GND.n976 240.244
R3666 GND.n4403 GND.n974 240.244
R3667 GND.n4407 GND.n974 240.244
R3668 GND.n4407 GND.n970 240.244
R3669 GND.n4413 GND.n970 240.244
R3670 GND.n4413 GND.n968 240.244
R3671 GND.n4417 GND.n968 240.244
R3672 GND.n4417 GND.n964 240.244
R3673 GND.n4423 GND.n964 240.244
R3674 GND.n4423 GND.n962 240.244
R3675 GND.n4427 GND.n962 240.244
R3676 GND.n4427 GND.n958 240.244
R3677 GND.n4433 GND.n958 240.244
R3678 GND.n4433 GND.n956 240.244
R3679 GND.n4437 GND.n956 240.244
R3680 GND.n4437 GND.n952 240.244
R3681 GND.n4443 GND.n952 240.244
R3682 GND.n4443 GND.n950 240.244
R3683 GND.n4447 GND.n950 240.244
R3684 GND.n4447 GND.n946 240.244
R3685 GND.n4453 GND.n946 240.244
R3686 GND.n4453 GND.n944 240.244
R3687 GND.n4457 GND.n944 240.244
R3688 GND.n4457 GND.n940 240.244
R3689 GND.n4463 GND.n940 240.244
R3690 GND.n4463 GND.n938 240.244
R3691 GND.n4467 GND.n938 240.244
R3692 GND.n4467 GND.n934 240.244
R3693 GND.n4473 GND.n934 240.244
R3694 GND.n4473 GND.n932 240.244
R3695 GND.n4477 GND.n932 240.244
R3696 GND.n4477 GND.n928 240.244
R3697 GND.n4483 GND.n928 240.244
R3698 GND.n4483 GND.n926 240.244
R3699 GND.n4487 GND.n926 240.244
R3700 GND.n4487 GND.n922 240.244
R3701 GND.n4493 GND.n922 240.244
R3702 GND.n4493 GND.n920 240.244
R3703 GND.n4497 GND.n920 240.244
R3704 GND.n4497 GND.n916 240.244
R3705 GND.n4503 GND.n916 240.244
R3706 GND.n4503 GND.n914 240.244
R3707 GND.n4507 GND.n914 240.244
R3708 GND.n4507 GND.n910 240.244
R3709 GND.n4513 GND.n910 240.244
R3710 GND.n4513 GND.n908 240.244
R3711 GND.n4517 GND.n908 240.244
R3712 GND.n4517 GND.n904 240.244
R3713 GND.n4523 GND.n904 240.244
R3714 GND.n4523 GND.n902 240.244
R3715 GND.n4527 GND.n902 240.244
R3716 GND.n4527 GND.n898 240.244
R3717 GND.n4533 GND.n898 240.244
R3718 GND.n4533 GND.n896 240.244
R3719 GND.n4537 GND.n896 240.244
R3720 GND.n4537 GND.n892 240.244
R3721 GND.n4543 GND.n892 240.244
R3722 GND.n4543 GND.n890 240.244
R3723 GND.n4547 GND.n890 240.244
R3724 GND.n4547 GND.n886 240.244
R3725 GND.n4553 GND.n886 240.244
R3726 GND.n4553 GND.n884 240.244
R3727 GND.n4557 GND.n884 240.244
R3728 GND.n4557 GND.n880 240.244
R3729 GND.n4563 GND.n880 240.244
R3730 GND.n4563 GND.n878 240.244
R3731 GND.n4567 GND.n878 240.244
R3732 GND.n4567 GND.n874 240.244
R3733 GND.n4573 GND.n874 240.244
R3734 GND.n4573 GND.n872 240.244
R3735 GND.n4577 GND.n872 240.244
R3736 GND.n4577 GND.n868 240.244
R3737 GND.n4583 GND.n868 240.244
R3738 GND.n4583 GND.n866 240.244
R3739 GND.n4587 GND.n866 240.244
R3740 GND.n4587 GND.n862 240.244
R3741 GND.n4593 GND.n862 240.244
R3742 GND.n4593 GND.n860 240.244
R3743 GND.n4597 GND.n860 240.244
R3744 GND.n4597 GND.n856 240.244
R3745 GND.n4603 GND.n856 240.244
R3746 GND.n4603 GND.n854 240.244
R3747 GND.n4607 GND.n854 240.244
R3748 GND.n4607 GND.n850 240.244
R3749 GND.n4613 GND.n850 240.244
R3750 GND.n4613 GND.n848 240.244
R3751 GND.n4617 GND.n848 240.244
R3752 GND.n4617 GND.n844 240.244
R3753 GND.n4623 GND.n844 240.244
R3754 GND.n4623 GND.n842 240.244
R3755 GND.n4627 GND.n842 240.244
R3756 GND.n4627 GND.n838 240.244
R3757 GND.n4633 GND.n838 240.244
R3758 GND.n4633 GND.n836 240.244
R3759 GND.n4637 GND.n836 240.244
R3760 GND.n4637 GND.n832 240.244
R3761 GND.n4643 GND.n832 240.244
R3762 GND.n4643 GND.n830 240.244
R3763 GND.n4647 GND.n830 240.244
R3764 GND.n4647 GND.n826 240.244
R3765 GND.n4653 GND.n826 240.244
R3766 GND.n4653 GND.n824 240.244
R3767 GND.n4657 GND.n824 240.244
R3768 GND.n4657 GND.n820 240.244
R3769 GND.n4663 GND.n820 240.244
R3770 GND.n4663 GND.n818 240.244
R3771 GND.n4667 GND.n818 240.244
R3772 GND.n4667 GND.n814 240.244
R3773 GND.n4673 GND.n814 240.244
R3774 GND.n4673 GND.n812 240.244
R3775 GND.n4677 GND.n812 240.244
R3776 GND.n4677 GND.n808 240.244
R3777 GND.n4683 GND.n808 240.244
R3778 GND.n4683 GND.n806 240.244
R3779 GND.n4687 GND.n806 240.244
R3780 GND.n4687 GND.n802 240.244
R3781 GND.n4693 GND.n802 240.244
R3782 GND.n4693 GND.n800 240.244
R3783 GND.n4697 GND.n800 240.244
R3784 GND.n4697 GND.n796 240.244
R3785 GND.n4703 GND.n796 240.244
R3786 GND.n4703 GND.n794 240.244
R3787 GND.n4707 GND.n794 240.244
R3788 GND.n4707 GND.n790 240.244
R3789 GND.n4713 GND.n790 240.244
R3790 GND.n4713 GND.n788 240.244
R3791 GND.n4717 GND.n788 240.244
R3792 GND.n4717 GND.n784 240.244
R3793 GND.n4723 GND.n784 240.244
R3794 GND.n4723 GND.n782 240.244
R3795 GND.n4727 GND.n782 240.244
R3796 GND.n4727 GND.n778 240.244
R3797 GND.n4733 GND.n778 240.244
R3798 GND.n4733 GND.n776 240.244
R3799 GND.n4737 GND.n776 240.244
R3800 GND.n4737 GND.n772 240.244
R3801 GND.n4743 GND.n772 240.244
R3802 GND.n4743 GND.n770 240.244
R3803 GND.n4747 GND.n770 240.244
R3804 GND.n4747 GND.n766 240.244
R3805 GND.n4753 GND.n766 240.244
R3806 GND.n4753 GND.n764 240.244
R3807 GND.n4757 GND.n764 240.244
R3808 GND.n4757 GND.n760 240.244
R3809 GND.n4763 GND.n760 240.244
R3810 GND.n4763 GND.n758 240.244
R3811 GND.n4767 GND.n758 240.244
R3812 GND.n4767 GND.n754 240.244
R3813 GND.n4773 GND.n754 240.244
R3814 GND.n4773 GND.n752 240.244
R3815 GND.n4777 GND.n752 240.244
R3816 GND.n4777 GND.n748 240.244
R3817 GND.n4783 GND.n748 240.244
R3818 GND.n4783 GND.n746 240.244
R3819 GND.n4787 GND.n746 240.244
R3820 GND.n4787 GND.n742 240.244
R3821 GND.n4793 GND.n742 240.244
R3822 GND.n4793 GND.n740 240.244
R3823 GND.n4797 GND.n740 240.244
R3824 GND.n4797 GND.n736 240.244
R3825 GND.n4803 GND.n736 240.244
R3826 GND.n4803 GND.n734 240.244
R3827 GND.n4807 GND.n734 240.244
R3828 GND.n4807 GND.n730 240.244
R3829 GND.n4813 GND.n730 240.244
R3830 GND.n4813 GND.n728 240.244
R3831 GND.n4817 GND.n728 240.244
R3832 GND.n4817 GND.n724 240.244
R3833 GND.n4823 GND.n724 240.244
R3834 GND.n4823 GND.n722 240.244
R3835 GND.n4827 GND.n722 240.244
R3836 GND.n4827 GND.n718 240.244
R3837 GND.n4833 GND.n718 240.244
R3838 GND.n4833 GND.n716 240.244
R3839 GND.n4837 GND.n716 240.244
R3840 GND.n4837 GND.n712 240.244
R3841 GND.n4843 GND.n712 240.244
R3842 GND.n4843 GND.n710 240.244
R3843 GND.n4847 GND.n710 240.244
R3844 GND.n4847 GND.n706 240.244
R3845 GND.n4853 GND.n706 240.244
R3846 GND.n4853 GND.n704 240.244
R3847 GND.n4857 GND.n704 240.244
R3848 GND.n4857 GND.n700 240.244
R3849 GND.n4863 GND.n700 240.244
R3850 GND.n4863 GND.n698 240.244
R3851 GND.n4867 GND.n698 240.244
R3852 GND.n4867 GND.n694 240.244
R3853 GND.n4873 GND.n694 240.244
R3854 GND.n4873 GND.n692 240.244
R3855 GND.n4877 GND.n692 240.244
R3856 GND.n4877 GND.n688 240.244
R3857 GND.n4883 GND.n688 240.244
R3858 GND.n4883 GND.n686 240.244
R3859 GND.n4887 GND.n686 240.244
R3860 GND.n4887 GND.n682 240.244
R3861 GND.n4893 GND.n682 240.244
R3862 GND.n4893 GND.n680 240.244
R3863 GND.n4897 GND.n680 240.244
R3864 GND.n4897 GND.n676 240.244
R3865 GND.n4903 GND.n676 240.244
R3866 GND.n4903 GND.n674 240.244
R3867 GND.n4907 GND.n674 240.244
R3868 GND.n4907 GND.n670 240.244
R3869 GND.n4913 GND.n670 240.244
R3870 GND.n4913 GND.n668 240.244
R3871 GND.n4917 GND.n668 240.244
R3872 GND.n4917 GND.n664 240.244
R3873 GND.n4923 GND.n664 240.244
R3874 GND.n4923 GND.n662 240.244
R3875 GND.n4927 GND.n662 240.244
R3876 GND.n4927 GND.n658 240.244
R3877 GND.n4933 GND.n658 240.244
R3878 GND.n4933 GND.n656 240.244
R3879 GND.n4937 GND.n656 240.244
R3880 GND.n4937 GND.n652 240.244
R3881 GND.n4943 GND.n652 240.244
R3882 GND.n4943 GND.n650 240.244
R3883 GND.n4947 GND.n650 240.244
R3884 GND.n4947 GND.n646 240.244
R3885 GND.n4953 GND.n646 240.244
R3886 GND.n4953 GND.n644 240.244
R3887 GND.n4957 GND.n644 240.244
R3888 GND.n4957 GND.n640 240.244
R3889 GND.n4963 GND.n640 240.244
R3890 GND.n4963 GND.n638 240.244
R3891 GND.n4967 GND.n638 240.244
R3892 GND.n4967 GND.n634 240.244
R3893 GND.n4973 GND.n634 240.244
R3894 GND.n4973 GND.n632 240.244
R3895 GND.n4977 GND.n632 240.244
R3896 GND.n4977 GND.n628 240.244
R3897 GND.n4983 GND.n628 240.244
R3898 GND.n4983 GND.n626 240.244
R3899 GND.n4987 GND.n626 240.244
R3900 GND.n4987 GND.n622 240.244
R3901 GND.n4993 GND.n622 240.244
R3902 GND.n4993 GND.n620 240.244
R3903 GND.n4997 GND.n620 240.244
R3904 GND.n4997 GND.n616 240.244
R3905 GND.n5003 GND.n616 240.244
R3906 GND.n5003 GND.n614 240.244
R3907 GND.n5007 GND.n614 240.244
R3908 GND.n5007 GND.n610 240.244
R3909 GND.n5013 GND.n610 240.244
R3910 GND.n5013 GND.n608 240.244
R3911 GND.n5017 GND.n608 240.244
R3912 GND.n5017 GND.n604 240.244
R3913 GND.n5023 GND.n604 240.244
R3914 GND.n5023 GND.n602 240.244
R3915 GND.n5027 GND.n602 240.244
R3916 GND.n5027 GND.n598 240.244
R3917 GND.n5033 GND.n598 240.244
R3918 GND.n5033 GND.n596 240.244
R3919 GND.n5037 GND.n596 240.244
R3920 GND.n5037 GND.n592 240.244
R3921 GND.n5043 GND.n592 240.244
R3922 GND.n5043 GND.n590 240.244
R3923 GND.n5047 GND.n590 240.244
R3924 GND.n5047 GND.n586 240.244
R3925 GND.n5053 GND.n586 240.244
R3926 GND.n5053 GND.n584 240.244
R3927 GND.n5057 GND.n584 240.244
R3928 GND.n5057 GND.n580 240.244
R3929 GND.n5063 GND.n580 240.244
R3930 GND.n5063 GND.n578 240.244
R3931 GND.n5067 GND.n578 240.244
R3932 GND.n5067 GND.n574 240.244
R3933 GND.n5073 GND.n574 240.244
R3934 GND.n5073 GND.n572 240.244
R3935 GND.n5077 GND.n572 240.244
R3936 GND.n5077 GND.n568 240.244
R3937 GND.n5083 GND.n568 240.244
R3938 GND.n5083 GND.n566 240.244
R3939 GND.n5087 GND.n566 240.244
R3940 GND.n5087 GND.n562 240.244
R3941 GND.n5093 GND.n562 240.244
R3942 GND.n5093 GND.n560 240.244
R3943 GND.n5097 GND.n560 240.244
R3944 GND.n5097 GND.n556 240.244
R3945 GND.n5103 GND.n556 240.244
R3946 GND.n5103 GND.n554 240.244
R3947 GND.n5107 GND.n554 240.244
R3948 GND.n5107 GND.n550 240.244
R3949 GND.n5114 GND.n550 240.244
R3950 GND.n5114 GND.n548 240.244
R3951 GND.n5118 GND.n545 240.244
R3952 GND.n5124 GND.n545 240.244
R3953 GND.n5124 GND.n543 240.244
R3954 GND.n5128 GND.n543 240.244
R3955 GND.n5128 GND.n539 240.244
R3956 GND.n5134 GND.n539 240.244
R3957 GND.n5134 GND.n537 240.244
R3958 GND.n5138 GND.n537 240.244
R3959 GND.n5138 GND.n533 240.244
R3960 GND.n5144 GND.n533 240.244
R3961 GND.n5144 GND.n531 240.244
R3962 GND.n5148 GND.n531 240.244
R3963 GND.n5148 GND.n527 240.244
R3964 GND.n5154 GND.n527 240.244
R3965 GND.n5154 GND.n525 240.244
R3966 GND.n5158 GND.n525 240.244
R3967 GND.n5158 GND.n521 240.244
R3968 GND.n5164 GND.n521 240.244
R3969 GND.n5164 GND.n519 240.244
R3970 GND.n5168 GND.n519 240.244
R3971 GND.n5168 GND.n515 240.244
R3972 GND.n5174 GND.n515 240.244
R3973 GND.n5174 GND.n513 240.244
R3974 GND.n5178 GND.n513 240.244
R3975 GND.n5178 GND.n509 240.244
R3976 GND.n5184 GND.n509 240.244
R3977 GND.n5184 GND.n507 240.244
R3978 GND.n5188 GND.n507 240.244
R3979 GND.n5188 GND.n503 240.244
R3980 GND.n5194 GND.n503 240.244
R3981 GND.n5194 GND.n501 240.244
R3982 GND.n5198 GND.n501 240.244
R3983 GND.n5198 GND.n497 240.244
R3984 GND.n5204 GND.n497 240.244
R3985 GND.n5204 GND.n495 240.244
R3986 GND.n5208 GND.n495 240.244
R3987 GND.n5208 GND.n491 240.244
R3988 GND.n5214 GND.n491 240.244
R3989 GND.n5214 GND.n489 240.244
R3990 GND.n5218 GND.n489 240.244
R3991 GND.n5218 GND.n485 240.244
R3992 GND.n5224 GND.n485 240.244
R3993 GND.n5224 GND.n483 240.244
R3994 GND.n5228 GND.n483 240.244
R3995 GND.n5228 GND.n479 240.244
R3996 GND.n5234 GND.n479 240.244
R3997 GND.n5234 GND.n477 240.244
R3998 GND.n5238 GND.n477 240.244
R3999 GND.n5238 GND.n473 240.244
R4000 GND.n5244 GND.n473 240.244
R4001 GND.n5244 GND.n471 240.244
R4002 GND.n5248 GND.n471 240.244
R4003 GND.n5248 GND.n467 240.244
R4004 GND.n5256 GND.n467 240.244
R4005 GND.n5256 GND.n465 240.244
R4006 GND.n4201 GND.n1141 240.244
R4007 GND.n4197 GND.n1141 240.244
R4008 GND.n4197 GND.n1147 240.244
R4009 GND.n4193 GND.n1147 240.244
R4010 GND.n4193 GND.n1149 240.244
R4011 GND.n4189 GND.n1149 240.244
R4012 GND.n4189 GND.n1155 240.244
R4013 GND.n4185 GND.n1155 240.244
R4014 GND.n4185 GND.n1157 240.244
R4015 GND.n4181 GND.n1157 240.244
R4016 GND.n4181 GND.n1163 240.244
R4017 GND.n4177 GND.n1163 240.244
R4018 GND.n4177 GND.n1165 240.244
R4019 GND.n4173 GND.n1165 240.244
R4020 GND.n4173 GND.n1171 240.244
R4021 GND.n4169 GND.n1171 240.244
R4022 GND.n4169 GND.n1173 240.244
R4023 GND.n4165 GND.n1173 240.244
R4024 GND.n4165 GND.n1179 240.244
R4025 GND.n4161 GND.n1179 240.244
R4026 GND.n4161 GND.n1181 240.244
R4027 GND.n4157 GND.n1181 240.244
R4028 GND.n4157 GND.n1187 240.244
R4029 GND.n4153 GND.n1187 240.244
R4030 GND.n4153 GND.n1189 240.244
R4031 GND.n4149 GND.n1189 240.244
R4032 GND.n4149 GND.n1195 240.244
R4033 GND.n4145 GND.n1195 240.244
R4034 GND.n4145 GND.n1197 240.244
R4035 GND.n4141 GND.n1197 240.244
R4036 GND.n4141 GND.n1203 240.244
R4037 GND.n4137 GND.n1203 240.244
R4038 GND.n4137 GND.n1205 240.244
R4039 GND.n4133 GND.n1205 240.244
R4040 GND.n4133 GND.n1211 240.244
R4041 GND.n4129 GND.n1211 240.244
R4042 GND.n4129 GND.n1213 240.244
R4043 GND.n4125 GND.n1213 240.244
R4044 GND.n4125 GND.n1219 240.244
R4045 GND.n4121 GND.n1219 240.244
R4046 GND.n4121 GND.n1221 240.244
R4047 GND.n4117 GND.n1221 240.244
R4048 GND.n4117 GND.n1227 240.244
R4049 GND.n4113 GND.n1227 240.244
R4050 GND.n4113 GND.n1229 240.244
R4051 GND.n4109 GND.n1229 240.244
R4052 GND.n4109 GND.n1235 240.244
R4053 GND.n4105 GND.n1235 240.244
R4054 GND.n4105 GND.n1237 240.244
R4055 GND.n4101 GND.n1237 240.244
R4056 GND.n4101 GND.n1243 240.244
R4057 GND.n4097 GND.n1243 240.244
R4058 GND.n4097 GND.n1245 240.244
R4059 GND.n4093 GND.n1245 240.244
R4060 GND.n4093 GND.n1251 240.244
R4061 GND.n4089 GND.n1251 240.244
R4062 GND.n4089 GND.n1253 240.244
R4063 GND.n4085 GND.n1253 240.244
R4064 GND.n4085 GND.n1259 240.244
R4065 GND.n4081 GND.n1259 240.244
R4066 GND.n4081 GND.n1261 240.244
R4067 GND.n4077 GND.n1261 240.244
R4068 GND.n4077 GND.n1267 240.244
R4069 GND.n4073 GND.n1267 240.244
R4070 GND.n4073 GND.n1269 240.244
R4071 GND.n4069 GND.n1269 240.244
R4072 GND.n4069 GND.n1275 240.244
R4073 GND.n4065 GND.n1275 240.244
R4074 GND.n4065 GND.n1277 240.244
R4075 GND.n4061 GND.n1277 240.244
R4076 GND.n4061 GND.n1283 240.244
R4077 GND.n4057 GND.n1283 240.244
R4078 GND.n4057 GND.n1285 240.244
R4079 GND.n4053 GND.n1285 240.244
R4080 GND.n4053 GND.n1291 240.244
R4081 GND.n4049 GND.n1291 240.244
R4082 GND.n4049 GND.n1293 240.244
R4083 GND.n4045 GND.n1293 240.244
R4084 GND.n4045 GND.n1299 240.244
R4085 GND.n4041 GND.n1299 240.244
R4086 GND.n4041 GND.n1301 240.244
R4087 GND.n4037 GND.n1301 240.244
R4088 GND.n4037 GND.n1307 240.244
R4089 GND.n4033 GND.n1307 240.244
R4090 GND.n4033 GND.n1309 240.244
R4091 GND.n4029 GND.n1309 240.244
R4092 GND.n4029 GND.n1315 240.244
R4093 GND.n4025 GND.n1315 240.244
R4094 GND.n4025 GND.n1317 240.244
R4095 GND.n4021 GND.n1317 240.244
R4096 GND.n4021 GND.n1323 240.244
R4097 GND.n4017 GND.n1323 240.244
R4098 GND.n4017 GND.n1325 240.244
R4099 GND.n4013 GND.n1325 240.244
R4100 GND.n4013 GND.n1331 240.244
R4101 GND.n4009 GND.n1331 240.244
R4102 GND.n4009 GND.n1333 240.244
R4103 GND.n4005 GND.n1333 240.244
R4104 GND.n4005 GND.n1339 240.244
R4105 GND.n4001 GND.n1339 240.244
R4106 GND.n4001 GND.n1341 240.244
R4107 GND.n3997 GND.n1341 240.244
R4108 GND.n3997 GND.n1347 240.244
R4109 GND.n3993 GND.n1347 240.244
R4110 GND.n3993 GND.n1349 240.244
R4111 GND.n3989 GND.n1349 240.244
R4112 GND.n3989 GND.n1355 240.244
R4113 GND.n2438 GND.n1355 240.244
R4114 GND.n2516 GND.n2438 240.244
R4115 GND.n2516 GND.n2439 240.244
R4116 GND.n2445 GND.n2439 240.244
R4117 GND.n2452 GND.n2445 240.244
R4118 GND.n2508 GND.n2452 240.244
R4119 GND.n2508 GND.n2507 240.244
R4120 GND.n2507 GND.n2506 240.244
R4121 GND.n2506 GND.n2504 240.244
R4122 GND.n2504 GND.n2501 240.244
R4123 GND.n2501 GND.n2500 240.244
R4124 GND.n2500 GND.n2497 240.244
R4125 GND.n2497 GND.n2496 240.244
R4126 GND.n2496 GND.n2453 240.244
R4127 GND.n2492 GND.n2453 240.244
R4128 GND.n2492 GND.n2491 240.244
R4129 GND.n2491 GND.n2490 240.244
R4130 GND.n2490 GND.n2456 240.244
R4131 GND.n2486 GND.n2456 240.244
R4132 GND.n2486 GND.n2485 240.244
R4133 GND.n2485 GND.n2483 240.244
R4134 GND.n2483 GND.n2462 240.244
R4135 GND.n2478 GND.n2462 240.244
R4136 GND.n2478 GND.n2477 240.244
R4137 GND.n2477 GND.n2472 240.244
R4138 GND.n2472 GND.n1563 240.244
R4139 GND.n3803 GND.n1563 240.244
R4140 GND.n3803 GND.n1564 240.244
R4141 GND.n3799 GND.n1564 240.244
R4142 GND.n3799 GND.n1570 240.244
R4143 GND.n2883 GND.n1570 240.244
R4144 GND.n2884 GND.n2883 240.244
R4145 GND.n2884 GND.n2878 240.244
R4146 GND.n2891 GND.n2878 240.244
R4147 GND.n2891 GND.n1655 240.244
R4148 GND.n3704 GND.n1655 240.244
R4149 GND.n3704 GND.n1656 240.244
R4150 GND.n3700 GND.n1656 240.244
R4151 GND.n3700 GND.n1662 240.244
R4152 GND.n1689 GND.n1662 240.244
R4153 GND.n1689 GND.n1685 240.244
R4154 GND.n3683 GND.n1685 240.244
R4155 GND.n3683 GND.n1686 240.244
R4156 GND.n3679 GND.n1686 240.244
R4157 GND.n3679 GND.n1697 240.244
R4158 GND.n3669 GND.n1697 240.244
R4159 GND.n3669 GND.n1709 240.244
R4160 GND.n3665 GND.n1709 240.244
R4161 GND.n3665 GND.n1715 240.244
R4162 GND.n3655 GND.n1715 240.244
R4163 GND.n3655 GND.n1726 240.244
R4164 GND.n3651 GND.n1726 240.244
R4165 GND.n3651 GND.n1732 240.244
R4166 GND.n3641 GND.n1732 240.244
R4167 GND.n3641 GND.n1744 240.244
R4168 GND.n3637 GND.n1744 240.244
R4169 GND.n3637 GND.n1750 240.244
R4170 GND.n3627 GND.n1750 240.244
R4171 GND.n3627 GND.n1761 240.244
R4172 GND.n3623 GND.n1761 240.244
R4173 GND.n3623 GND.n1767 240.244
R4174 GND.n3613 GND.n1767 240.244
R4175 GND.n3613 GND.n1779 240.244
R4176 GND.n3609 GND.n1779 240.244
R4177 GND.n3609 GND.n1785 240.244
R4178 GND.n1811 GND.n1785 240.244
R4179 GND.n1811 GND.n1807 240.244
R4180 GND.n3592 GND.n1807 240.244
R4181 GND.n3592 GND.n1808 240.244
R4182 GND.n3588 GND.n1808 240.244
R4183 GND.n3588 GND.n1819 240.244
R4184 GND.n1862 GND.n1819 240.244
R4185 GND.n3573 GND.n1862 240.244
R4186 GND.n3573 GND.n1863 240.244
R4187 GND.n3569 GND.n1863 240.244
R4188 GND.n3569 GND.n1871 240.244
R4189 GND.n1885 GND.n1871 240.244
R4190 GND.n3559 GND.n1885 240.244
R4191 GND.n3559 GND.n1886 240.244
R4192 GND.n3555 GND.n1886 240.244
R4193 GND.n3555 GND.n1894 240.244
R4194 GND.n3507 GND.n1894 240.244
R4195 GND.n3507 GND.n1939 240.244
R4196 GND.n3503 GND.n1939 240.244
R4197 GND.n3503 GND.n3502 240.244
R4198 GND.n3502 GND.n1945 240.244
R4199 GND.n2204 GND.n1945 240.244
R4200 GND.n2205 GND.n2204 240.244
R4201 GND.n2206 GND.n2205 240.244
R4202 GND.n2206 GND.n2195 240.244
R4203 GND.n2213 GND.n2195 240.244
R4204 GND.n2214 GND.n2213 240.244
R4205 GND.n2215 GND.n2214 240.244
R4206 GND.n2215 GND.n2192 240.244
R4207 GND.n3375 GND.n2192 240.244
R4208 GND.n3375 GND.n2193 240.244
R4209 GND.n3370 GND.n2193 240.244
R4210 GND.n3370 GND.n2220 240.244
R4211 GND.n3360 GND.n2220 240.244
R4212 GND.n3360 GND.n3340 240.244
R4213 GND.n3355 GND.n3340 240.244
R4214 GND.n3355 GND.n3354 240.244
R4215 GND.n3354 GND.n3343 240.244
R4216 GND.n3350 GND.n3343 240.244
R4217 GND.n3350 GND.n3349 240.244
R4218 GND.n3349 GND.n62 240.244
R4219 GND.n5472 GND.n62 240.244
R4220 GND.n5472 GND.n63 240.244
R4221 GND.n5468 GND.n63 240.244
R4222 GND.n5468 GND.n69 240.244
R4223 GND.n5464 GND.n69 240.244
R4224 GND.n5464 GND.n260 240.244
R4225 GND.n5460 GND.n260 240.244
R4226 GND.n5460 GND.n266 240.244
R4227 GND.n5456 GND.n266 240.244
R4228 GND.n5456 GND.n268 240.244
R4229 GND.n5452 GND.n268 240.244
R4230 GND.n5452 GND.n274 240.244
R4231 GND.n5448 GND.n274 240.244
R4232 GND.n5448 GND.n276 240.244
R4233 GND.n5444 GND.n276 240.244
R4234 GND.n5444 GND.n282 240.244
R4235 GND.n5440 GND.n282 240.244
R4236 GND.n5440 GND.n284 240.244
R4237 GND.n5436 GND.n284 240.244
R4238 GND.n5436 GND.n290 240.244
R4239 GND.n5432 GND.n290 240.244
R4240 GND.n5432 GND.n292 240.244
R4241 GND.n5428 GND.n292 240.244
R4242 GND.n5428 GND.n298 240.244
R4243 GND.n5424 GND.n298 240.244
R4244 GND.n5424 GND.n300 240.244
R4245 GND.n5420 GND.n300 240.244
R4246 GND.n5420 GND.n306 240.244
R4247 GND.n5416 GND.n306 240.244
R4248 GND.n5416 GND.n308 240.244
R4249 GND.n5412 GND.n308 240.244
R4250 GND.n5412 GND.n314 240.244
R4251 GND.n5408 GND.n314 240.244
R4252 GND.n5408 GND.n316 240.244
R4253 GND.n5404 GND.n316 240.244
R4254 GND.n5404 GND.n322 240.244
R4255 GND.n5400 GND.n322 240.244
R4256 GND.n5400 GND.n324 240.244
R4257 GND.n5396 GND.n324 240.244
R4258 GND.n5396 GND.n330 240.244
R4259 GND.n5392 GND.n330 240.244
R4260 GND.n5392 GND.n332 240.244
R4261 GND.n5388 GND.n332 240.244
R4262 GND.n5388 GND.n338 240.244
R4263 GND.n5384 GND.n338 240.244
R4264 GND.n5384 GND.n340 240.244
R4265 GND.n5380 GND.n340 240.244
R4266 GND.n5380 GND.n346 240.244
R4267 GND.n5376 GND.n346 240.244
R4268 GND.n5376 GND.n348 240.244
R4269 GND.n5372 GND.n348 240.244
R4270 GND.n5372 GND.n354 240.244
R4271 GND.n5368 GND.n354 240.244
R4272 GND.n5368 GND.n356 240.244
R4273 GND.n5364 GND.n356 240.244
R4274 GND.n5364 GND.n362 240.244
R4275 GND.n5360 GND.n362 240.244
R4276 GND.n5360 GND.n364 240.244
R4277 GND.n5356 GND.n364 240.244
R4278 GND.n5356 GND.n370 240.244
R4279 GND.n5352 GND.n370 240.244
R4280 GND.n5352 GND.n372 240.244
R4281 GND.n5348 GND.n372 240.244
R4282 GND.n5348 GND.n378 240.244
R4283 GND.n5344 GND.n378 240.244
R4284 GND.n5344 GND.n380 240.244
R4285 GND.n5340 GND.n380 240.244
R4286 GND.n5340 GND.n386 240.244
R4287 GND.n5336 GND.n386 240.244
R4288 GND.n5336 GND.n388 240.244
R4289 GND.n5332 GND.n388 240.244
R4290 GND.n5332 GND.n394 240.244
R4291 GND.n5328 GND.n394 240.244
R4292 GND.n5328 GND.n396 240.244
R4293 GND.n5324 GND.n396 240.244
R4294 GND.n5324 GND.n402 240.244
R4295 GND.n5320 GND.n402 240.244
R4296 GND.n5320 GND.n404 240.244
R4297 GND.n5316 GND.n404 240.244
R4298 GND.n5316 GND.n410 240.244
R4299 GND.n5312 GND.n410 240.244
R4300 GND.n5312 GND.n412 240.244
R4301 GND.n5308 GND.n412 240.244
R4302 GND.n5308 GND.n418 240.244
R4303 GND.n5304 GND.n418 240.244
R4304 GND.n5304 GND.n420 240.244
R4305 GND.n5300 GND.n420 240.244
R4306 GND.n5300 GND.n426 240.244
R4307 GND.n5296 GND.n426 240.244
R4308 GND.n5296 GND.n428 240.244
R4309 GND.n5292 GND.n428 240.244
R4310 GND.n5292 GND.n434 240.244
R4311 GND.n5288 GND.n434 240.244
R4312 GND.n5288 GND.n436 240.244
R4313 GND.n5284 GND.n436 240.244
R4314 GND.n5284 GND.n442 240.244
R4315 GND.n5280 GND.n442 240.244
R4316 GND.n5280 GND.n444 240.244
R4317 GND.n5276 GND.n444 240.244
R4318 GND.n5276 GND.n450 240.244
R4319 GND.n5272 GND.n450 240.244
R4320 GND.n5272 GND.n452 240.244
R4321 GND.n5268 GND.n452 240.244
R4322 GND.n5268 GND.n458 240.244
R4323 GND.n5264 GND.n458 240.244
R4324 GND.n5264 GND.n460 240.244
R4325 GND.n5260 GND.n460 240.244
R4326 GND.n4313 GND.n1030 240.244
R4327 GND.n4309 GND.n1030 240.244
R4328 GND.n4309 GND.n1035 240.244
R4329 GND.n4305 GND.n1035 240.244
R4330 GND.n4305 GND.n1037 240.244
R4331 GND.n4301 GND.n1037 240.244
R4332 GND.n4301 GND.n1043 240.244
R4333 GND.n4297 GND.n1043 240.244
R4334 GND.n4297 GND.n1045 240.244
R4335 GND.n4293 GND.n1045 240.244
R4336 GND.n4293 GND.n1051 240.244
R4337 GND.n4289 GND.n1051 240.244
R4338 GND.n4289 GND.n1053 240.244
R4339 GND.n4285 GND.n1053 240.244
R4340 GND.n4285 GND.n1059 240.244
R4341 GND.n4281 GND.n1059 240.244
R4342 GND.n4281 GND.n1061 240.244
R4343 GND.n4277 GND.n1061 240.244
R4344 GND.n4277 GND.n1067 240.244
R4345 GND.n4273 GND.n1067 240.244
R4346 GND.n4273 GND.n1069 240.244
R4347 GND.n4269 GND.n1069 240.244
R4348 GND.n4269 GND.n1075 240.244
R4349 GND.n4265 GND.n1075 240.244
R4350 GND.n4265 GND.n1077 240.244
R4351 GND.n4261 GND.n1077 240.244
R4352 GND.n4261 GND.n1083 240.244
R4353 GND.n4257 GND.n1083 240.244
R4354 GND.n4257 GND.n1085 240.244
R4355 GND.n4253 GND.n1085 240.244
R4356 GND.n4253 GND.n1091 240.244
R4357 GND.n4249 GND.n1091 240.244
R4358 GND.n4249 GND.n1093 240.244
R4359 GND.n4245 GND.n1093 240.244
R4360 GND.n4245 GND.n1099 240.244
R4361 GND.n4241 GND.n1099 240.244
R4362 GND.n4241 GND.n1101 240.244
R4363 GND.n4237 GND.n1101 240.244
R4364 GND.n4237 GND.n1107 240.244
R4365 GND.n4233 GND.n1107 240.244
R4366 GND.n4233 GND.n1109 240.244
R4367 GND.n4229 GND.n1109 240.244
R4368 GND.n4229 GND.n1115 240.244
R4369 GND.n4225 GND.n1115 240.244
R4370 GND.n4225 GND.n1117 240.244
R4371 GND.n4221 GND.n1117 240.244
R4372 GND.n4221 GND.n1123 240.244
R4373 GND.n4217 GND.n1123 240.244
R4374 GND.n4217 GND.n1125 240.244
R4375 GND.n4213 GND.n1125 240.244
R4376 GND.n4213 GND.n1131 240.244
R4377 GND.n4209 GND.n1131 240.244
R4378 GND.n4209 GND.n1133 240.244
R4379 GND.n4205 GND.n1133 240.244
R4380 GND.n4205 GND.n1139 240.244
R4381 GND.n2732 GND.n2536 240.244
R4382 GND.n2736 GND.n2734 240.244
R4383 GND.n2742 GND.n2532 240.244
R4384 GND.n2746 GND.n2744 240.244
R4385 GND.n2752 GND.n2528 240.244
R4386 GND.n2755 GND.n2754 240.244
R4387 GND.n1371 GND.n1360 240.244
R4388 GND.n3980 GND.n1371 240.244
R4389 GND.n3980 GND.n1372 240.244
R4390 GND.n2772 GND.n1372 240.244
R4391 GND.n2775 GND.n2772 240.244
R4392 GND.n2775 GND.n2774 240.244
R4393 GND.n2774 GND.n2425 240.244
R4394 GND.n2425 GND.n2413 240.244
R4395 GND.n2796 GND.n2413 240.244
R4396 GND.n2800 GND.n2796 240.244
R4397 GND.n2800 GND.n2799 240.244
R4398 GND.n2799 GND.n2403 240.244
R4399 GND.n2403 GND.n2393 240.244
R4400 GND.n2825 GND.n2393 240.244
R4401 GND.n2827 GND.n2825 240.244
R4402 GND.n2827 GND.n2382 240.244
R4403 GND.n2837 GND.n2382 240.244
R4404 GND.n2838 GND.n2837 240.244
R4405 GND.n2838 GND.n1415 240.244
R4406 GND.n1538 GND.n1537 240.244
R4407 GND.n2364 GND.n2363 240.244
R4408 GND.n2367 GND.n2366 240.244
R4409 GND.n2372 GND.n2369 240.244
R4410 GND.n2375 GND.n2374 240.244
R4411 GND.n2762 GND.n1358 240.244
R4412 GND.n2762 GND.n1370 240.244
R4413 GND.n2519 GND.n1370 240.244
R4414 GND.n2770 GND.n2519 240.244
R4415 GND.n2770 GND.n2435 240.244
R4416 GND.n2435 GND.n2421 240.244
R4417 GND.n2786 GND.n2421 240.244
R4418 GND.n2786 GND.n2416 240.244
R4419 GND.n2794 GND.n2416 240.244
R4420 GND.n2794 GND.n2411 240.244
R4421 GND.n2411 GND.n2400 240.244
R4422 GND.n2811 GND.n2400 240.244
R4423 GND.n2811 GND.n2395 240.244
R4424 GND.n2823 GND.n2395 240.244
R4425 GND.n2823 GND.n2391 240.244
R4426 GND.n2817 GND.n2391 240.244
R4427 GND.n2817 GND.n2380 240.244
R4428 GND.n2840 GND.n2380 240.244
R4429 GND.n2840 GND.n1412 240.244
R4430 GND.n1617 GND.n1616 240.132
R4431 GND.n1850 GND.n1849 240.132
R4432 GND.n1635 GND.t62 228.995
R4433 GND.n1637 GND.t75 228.995
R4434 GND.n2019 GND.t72 228.995
R4435 GND.n2068 GND.t55 228.995
R4436 GND.n2106 GND.n1955 199.319
R4437 GND.n2106 GND.n1956 199.319
R4438 GND.n3912 GND.n3911 199.319
R4439 GND.n3911 GND.n3910 199.319
R4440 GND.n1931 GND.t89 195.297
R4441 GND.n3862 GND.t41 195.297
R4442 GND.n1618 GND.n1614 186.49
R4443 GND.n1851 GND.n1847 186.49
R4444 GND.n2064 GND.n1859 163.367
R4445 GND.n2100 GND.n2065 163.367
R4446 GND.n2096 GND.n2095 163.367
R4447 GND.n2092 GND.n2091 163.367
R4448 GND.n2088 GND.n2087 163.367
R4449 GND.n2084 GND.n2083 163.367
R4450 GND.n2080 GND.n2079 163.367
R4451 GND.n2075 GND.n2074 163.367
R4452 GND.n2071 GND.n2070 163.367
R4453 GND.n2103 GND.n2008 163.367
R4454 GND.n2024 GND.n2023 163.367
R4455 GND.n2028 GND.n2027 163.367
R4456 GND.n2032 GND.n2031 163.367
R4457 GND.n2036 GND.n2035 163.367
R4458 GND.n2040 GND.n2039 163.367
R4459 GND.n2044 GND.n2043 163.367
R4460 GND.n2048 GND.n2047 163.367
R4461 GND.n2050 GND.n2018 163.367
R4462 GND.n3714 GND.n1640 163.367
R4463 GND.n2897 GND.n1640 163.367
R4464 GND.n2897 GND.n2893 163.367
R4465 GND.n2893 GND.n1654 163.367
R4466 GND.n2345 GND.n1654 163.367
R4467 GND.n2952 GND.n2345 163.367
R4468 GND.n2952 GND.n1663 163.367
R4469 GND.n2956 GND.n1663 163.367
R4470 GND.n2956 GND.n1671 163.367
R4471 GND.n2342 GND.n1671 163.367
R4472 GND.n2964 GND.n2342 163.367
R4473 GND.n2964 GND.n2343 163.367
R4474 GND.n2960 GND.n2343 163.367
R4475 GND.n2960 GND.n2336 163.367
R4476 GND.n2976 GND.n2336 163.367
R4477 GND.n2976 GND.n1699 163.367
R4478 GND.n2981 GND.n1699 163.367
R4479 GND.n2981 GND.n1707 163.367
R4480 GND.n2333 GND.n1707 163.367
R4481 GND.n3029 GND.n2333 163.367
R4482 GND.n3029 GND.n2334 163.367
R4483 GND.n2334 GND.n1717 163.367
R4484 GND.n3024 GND.n1717 163.367
R4485 GND.n3024 GND.n1724 163.367
R4486 GND.n3021 GND.n1724 163.367
R4487 GND.n3021 GND.n3020 163.367
R4488 GND.n3020 GND.n3015 163.367
R4489 GND.n3015 GND.n1734 163.367
R4490 GND.n3011 GND.n1734 163.367
R4491 GND.n3011 GND.n1742 163.367
R4492 GND.n3007 GND.n1742 163.367
R4493 GND.n3007 GND.n3006 163.367
R4494 GND.n3006 GND.n3005 163.367
R4495 GND.n3005 GND.n1752 163.367
R4496 GND.n3001 GND.n1752 163.367
R4497 GND.n3001 GND.n1759 163.367
R4498 GND.n2998 GND.n1759 163.367
R4499 GND.n2998 GND.n2997 163.367
R4500 GND.n2997 GND.n2996 163.367
R4501 GND.n2996 GND.n1769 163.367
R4502 GND.n2992 GND.n1769 163.367
R4503 GND.n2992 GND.n1777 163.367
R4504 GND.n2271 GND.n1777 163.367
R4505 GND.n3121 GND.n2271 163.367
R4506 GND.n3122 GND.n3121 163.367
R4507 GND.n3123 GND.n3122 163.367
R4508 GND.n3123 GND.n2269 163.367
R4509 GND.n3140 GND.n2269 163.367
R4510 GND.n3140 GND.n1798 163.367
R4511 GND.n3136 GND.n1798 163.367
R4512 GND.n3136 GND.n1805 163.367
R4513 GND.n3131 GND.n1805 163.367
R4514 GND.n3131 GND.n1823 163.367
R4515 GND.n3586 GND.n1823 163.367
R4516 GND.n3586 GND.n1824 163.367
R4517 GND.n3582 GND.n1824 163.367
R4518 GND.n3582 GND.n1827 163.367
R4519 GND.n1860 GND.n1827 163.367
R4520 GND.n1607 GND.n1606 163.367
R4521 GND.n3783 GND.n1606 163.367
R4522 GND.n3781 GND.n3780 163.367
R4523 GND.n3777 GND.n3776 163.367
R4524 GND.n3773 GND.n3772 163.367
R4525 GND.n3769 GND.n3768 163.367
R4526 GND.n3765 GND.n3764 163.367
R4527 GND.n3760 GND.n3759 163.367
R4528 GND.n3756 GND.n3755 163.367
R4529 GND.n3750 GND.n3749 163.367
R4530 GND.n3746 GND.n3745 163.367
R4531 GND.n3741 GND.n3740 163.367
R4532 GND.n3737 GND.n3736 163.367
R4533 GND.n3733 GND.n3732 163.367
R4534 GND.n3729 GND.n3728 163.367
R4535 GND.n3725 GND.n3724 163.367
R4536 GND.n3721 GND.n3720 163.367
R4537 GND.n3717 GND.n1604 163.367
R4538 GND.n2899 GND.n1608 163.367
R4539 GND.n2910 GND.n2899 163.367
R4540 GND.n2910 GND.n2900 163.367
R4541 GND.n2900 GND.n1653 163.367
R4542 GND.n2905 GND.n1653 163.367
R4543 GND.n2905 GND.n1665 163.367
R4544 GND.n3697 GND.n1665 163.367
R4545 GND.n3697 GND.n1666 163.367
R4546 GND.n3693 GND.n1666 163.367
R4547 GND.n3693 GND.n1669 163.367
R4548 GND.n2967 GND.n1669 163.367
R4549 GND.n2968 GND.n2967 163.367
R4550 GND.n2968 GND.n2338 163.367
R4551 GND.n2972 GND.n2338 163.367
R4552 GND.n2972 GND.n1701 163.367
R4553 GND.n3676 GND.n1701 163.367
R4554 GND.n3676 GND.n1702 163.367
R4555 GND.n3672 GND.n1702 163.367
R4556 GND.n3672 GND.n1705 163.367
R4557 GND.n3033 GND.n1705 163.367
R4558 GND.n3033 GND.n1718 163.367
R4559 GND.n3662 GND.n1718 163.367
R4560 GND.n3662 GND.n1719 163.367
R4561 GND.n3658 GND.n1719 163.367
R4562 GND.n3658 GND.n1722 163.367
R4563 GND.n3018 GND.n1722 163.367
R4564 GND.n3018 GND.n1736 163.367
R4565 GND.n3648 GND.n1736 163.367
R4566 GND.n3648 GND.n1737 163.367
R4567 GND.n3644 GND.n1737 163.367
R4568 GND.n3644 GND.n1740 163.367
R4569 GND.n2300 GND.n1740 163.367
R4570 GND.n2300 GND.n1754 163.367
R4571 GND.n3634 GND.n1754 163.367
R4572 GND.n3634 GND.n1755 163.367
R4573 GND.n3630 GND.n1755 163.367
R4574 GND.n3630 GND.n1758 163.367
R4575 GND.n2282 GND.n1758 163.367
R4576 GND.n2282 GND.n1771 163.367
R4577 GND.n3620 GND.n1771 163.367
R4578 GND.n3620 GND.n1772 163.367
R4579 GND.n3616 GND.n1772 163.367
R4580 GND.n3616 GND.n1775 163.367
R4581 GND.n3119 GND.n1775 163.367
R4582 GND.n3119 GND.n3112 163.367
R4583 GND.n3115 GND.n3112 163.367
R4584 GND.n3115 GND.n3114 163.367
R4585 GND.n3114 GND.n1800 163.367
R4586 GND.n3599 GND.n1800 163.367
R4587 GND.n3599 GND.n1801 163.367
R4588 GND.n3595 GND.n1801 163.367
R4589 GND.n3595 GND.n1804 163.367
R4590 GND.n3128 GND.n1804 163.367
R4591 GND.n3128 GND.n1821 163.367
R4592 GND.n1831 GND.n1821 163.367
R4593 GND.n3580 GND.n1831 163.367
R4594 GND.n3580 GND.n1832 163.367
R4595 GND.n3576 GND.n1832 163.367
R4596 GND.n1857 GND.n1856 153.553
R4597 GND.n1839 GND.t103 153.314
R4598 GND.n1623 GND.n1622 152
R4599 GND.n1624 GND.n1612 152
R4600 GND.n1626 GND.n1625 152
R4601 GND.n1627 GND.n1611 152
R4602 GND.n1629 GND.n1628 152
R4603 GND.n1631 GND.n1609 152
R4604 GND.n1633 GND.n1632 152
R4605 GND.n1855 GND.n1834 152
R4606 GND.n1846 GND.n1835 152
R4607 GND.n1845 GND.n1844 152
R4608 GND.n1843 GND.n1836 152
R4609 GND.n1842 GND.n1841 152
R4610 GND.n1840 GND.n1837 152
R4611 GND.n1637 GND.t77 145.85
R4612 GND.n2019 GND.t73 145.85
R4613 GND.n1635 GND.t65 145.847
R4614 GND.n2068 GND.t57 145.847
R4615 GND.n1932 GND.t90 144.873
R4616 GND.n3863 GND.t40 144.873
R4617 GND.n2104 GND.n2007 143.351
R4618 GND.n3752 GND.n1594 143.351
R4619 GND.n3752 GND.n1595 143.351
R4620 GND.n1619 GND.t22 135.757
R4621 GND.n1632 GND.t8 126.766
R4622 GND.n1630 GND.t69 126.766
R4623 GND.n1611 GND.t121 126.766
R4624 GND.n1624 GND.t48 126.766
R4625 GND.n1613 GND.t106 126.766
R4626 GND.n1838 GND.t42 126.766
R4627 GND.n1842 GND.t84 126.766
R4628 GND.n1844 GND.t66 126.766
R4629 GND.n1854 GND.t91 126.766
R4630 GND.n1856 GND.t35 126.766
R4631 GND.n2376 GND.t116 118.868
R4632 GND.n1433 GND.t29 118.868
R4633 GND.n1491 GND.t98 118.868
R4634 GND.n1520 GND.t17 118.868
R4635 GND.n1450 GND.t113 118.868
R4636 GND.n1991 GND.t102 118.868
R4637 GND.n2108 GND.t126 118.868
R4638 GND.n2124 GND.t34 118.868
R4639 GND.n2139 GND.t80 118.868
R4640 GND.n150 GND.t110 118.868
R4641 GND.n135 GND.t60 118.868
R4642 GND.n206 GND.t53 118.868
R4643 GND.n106 GND.t119 118.868
R4644 GND.n3277 GND.t82 118.868
R4645 GND.n2249 GND.t47 118.868
R4646 GND.n2584 GND.t96 118.868
R4647 GND.n2567 GND.t14 118.868
R4648 GND.n2686 GND.t27 118.868
R4649 GND.n2539 GND.t21 118.868
R4650 GND.n2524 GND.t129 118.868
R4651 GND.n249 GND.n94 99.6594
R4652 GND.n247 GND.n93 99.6594
R4653 GND.n243 GND.n92 99.6594
R4654 GND.n239 GND.n91 99.6594
R4655 GND.n235 GND.n90 99.6594
R4656 GND.n231 GND.n89 99.6594
R4657 GND.n227 GND.n88 99.6594
R4658 GND.n223 GND.n87 99.6594
R4659 GND.n219 GND.n86 99.6594
R4660 GND.n215 GND.n85 99.6594
R4661 GND.n211 GND.n84 99.6594
R4662 GND.n204 GND.n83 99.6594
R4663 GND.n200 GND.n82 99.6594
R4664 GND.n196 GND.n81 99.6594
R4665 GND.n192 GND.n80 99.6594
R4666 GND.n188 GND.n79 99.6594
R4667 GND.n184 GND.n78 99.6594
R4668 GND.n138 GND.n77 99.6594
R4669 GND.n176 GND.n76 99.6594
R4670 GND.n172 GND.n75 99.6594
R4671 GND.n168 GND.n74 99.6594
R4672 GND.n164 GND.n73 99.6594
R4673 GND.n160 GND.n72 99.6594
R4674 GND.n156 GND.n71 99.6594
R4675 GND.n70 GND.n59 99.6594
R4676 GND.n3499 GND.n3498 99.6594
R4677 GND.n3493 GND.n1946 99.6594
R4678 GND.n3490 GND.n1947 99.6594
R4679 GND.n3486 GND.n1948 99.6594
R4680 GND.n3482 GND.n1949 99.6594
R4681 GND.n3478 GND.n1950 99.6594
R4682 GND.n3474 GND.n1951 99.6594
R4683 GND.n3470 GND.n1952 99.6594
R4684 GND.n3466 GND.n1953 99.6594
R4685 GND.n3462 GND.n1954 99.6594
R4686 GND.n3458 GND.n1955 99.6594
R4687 GND.n3453 GND.n1957 99.6594
R4688 GND.n3449 GND.n1958 99.6594
R4689 GND.n3445 GND.n1959 99.6594
R4690 GND.n3441 GND.n1960 99.6594
R4691 GND.n3437 GND.n1961 99.6594
R4692 GND.n3433 GND.n1962 99.6594
R4693 GND.n3429 GND.n1963 99.6594
R4694 GND.n3426 GND.n1964 99.6594
R4695 GND.n3422 GND.n1965 99.6594
R4696 GND.n3418 GND.n1966 99.6594
R4697 GND.n3414 GND.n1967 99.6594
R4698 GND.n3410 GND.n1968 99.6594
R4699 GND.n2138 GND.n1969 99.6594
R4700 GND.n1466 GND.n1422 99.6594
R4701 GND.n1465 GND.n1425 99.6594
R4702 GND.n1463 GND.n1427 99.6594
R4703 GND.n1462 GND.n1430 99.6594
R4704 GND.n1460 GND.n1432 99.6594
R4705 GND.n1459 GND.n1438 99.6594
R4706 GND.n1458 GND.n1457 99.6594
R4707 GND.n1456 GND.n1443 99.6594
R4708 GND.n1455 GND.n1454 99.6594
R4709 GND.n1453 GND.n1448 99.6594
R4710 GND.n3910 GND.n3909 99.6594
R4711 GND.n1473 GND.n1472 99.6594
R4712 GND.n1476 GND.n1475 99.6594
R4713 GND.n1481 GND.n1480 99.6594
R4714 GND.n1484 GND.n1483 99.6594
R4715 GND.n1489 GND.n1488 99.6594
R4716 GND.n1495 GND.n1494 99.6594
R4717 GND.n1500 GND.n1499 99.6594
R4718 GND.n1503 GND.n1502 99.6594
R4719 GND.n1508 GND.n1507 99.6594
R4720 GND.n1511 GND.n1510 99.6594
R4721 GND.n1516 GND.n1515 99.6594
R4722 GND.n1519 GND.n1518 99.6594
R4723 GND.n1523 GND.n1410 99.6594
R4724 GND.n2597 GND.n1361 99.6594
R4725 GND.n2600 GND.n2599 99.6594
R4726 GND.n2607 GND.n2606 99.6594
R4727 GND.n2610 GND.n2609 99.6594
R4728 GND.n2617 GND.n2616 99.6594
R4729 GND.n2620 GND.n2619 99.6594
R4730 GND.n2627 GND.n2626 99.6594
R4731 GND.n2630 GND.n2629 99.6594
R4732 GND.n2637 GND.n2636 99.6594
R4733 GND.n2640 GND.n2639 99.6594
R4734 GND.n2648 GND.n2647 99.6594
R4735 GND.n2651 GND.n2650 99.6594
R4736 GND.n2658 GND.n2657 99.6594
R4737 GND.n2661 GND.n2660 99.6594
R4738 GND.n2668 GND.n2667 99.6594
R4739 GND.n2671 GND.n2670 99.6594
R4740 GND.n2678 GND.n2677 99.6594
R4741 GND.n2681 GND.n2680 99.6594
R4742 GND.n2690 GND.n2689 99.6594
R4743 GND.n2693 GND.n2692 99.6594
R4744 GND.n2700 GND.n2699 99.6594
R4745 GND.n2703 GND.n2702 99.6594
R4746 GND.n2710 GND.n2709 99.6594
R4747 GND.n2713 GND.n2712 99.6594
R4748 GND.n2720 GND.n2719 99.6594
R4749 GND.n3544 GND.n3543 99.6594
R4750 GND.n3539 GND.n1916 99.6594
R4751 GND.n3535 GND.n1915 99.6594
R4752 GND.n3531 GND.n1914 99.6594
R4753 GND.n3527 GND.n1913 99.6594
R4754 GND.n3523 GND.n1912 99.6594
R4755 GND.n3519 GND.n1911 99.6594
R4756 GND.n3515 GND.n1910 99.6594
R4757 GND.n3511 GND.n1909 99.6594
R4758 GND.n3849 GND.n3848 99.6594
R4759 GND.n3843 GND.n1544 99.6594
R4760 GND.n3840 GND.n1545 99.6594
R4761 GND.n3836 GND.n1546 99.6594
R4762 GND.n3832 GND.n1547 99.6594
R4763 GND.n3828 GND.n1548 99.6594
R4764 GND.n3824 GND.n1549 99.6594
R4765 GND.n1550 GND.n1529 99.6594
R4766 GND.n3851 GND.n1542 99.6594
R4767 GND.n3294 GND.n3288 99.6594
R4768 GND.n3298 GND.n3296 99.6594
R4769 GND.n3304 GND.n3284 99.6594
R4770 GND.n3309 GND.n3306 99.6594
R4771 GND.n3307 GND.n3280 99.6594
R4772 GND.n3318 GND.n3317 99.6594
R4773 GND.n2149 GND.n1970 99.6594
R4774 GND.n3208 GND.n1971 99.6594
R4775 GND.n3210 GND.n1972 99.6594
R4776 GND.n3219 GND.n1973 99.6594
R4777 GND.n3221 GND.n1974 99.6594
R4778 GND.n3229 GND.n1975 99.6594
R4779 GND.n3207 GND.n1970 99.6594
R4780 GND.n3211 GND.n1971 99.6594
R4781 GND.n3218 GND.n1972 99.6594
R4782 GND.n3222 GND.n1973 99.6594
R4783 GND.n3228 GND.n1974 99.6594
R4784 GND.n3232 GND.n1975 99.6594
R4785 GND.n3317 GND.n3316 99.6594
R4786 GND.n3308 GND.n3307 99.6594
R4787 GND.n3306 GND.n3305 99.6594
R4788 GND.n3297 GND.n3284 99.6594
R4789 GND.n3296 GND.n3295 99.6594
R4790 GND.n3289 GND.n3288 99.6594
R4791 GND.n3849 GND.n1553 99.6594
R4792 GND.n3841 GND.n1544 99.6594
R4793 GND.n3837 GND.n1545 99.6594
R4794 GND.n3833 GND.n1546 99.6594
R4795 GND.n3829 GND.n1547 99.6594
R4796 GND.n3825 GND.n1548 99.6594
R4797 GND.n1549 GND.n1528 99.6594
R4798 GND.n1550 GND.n1530 99.6594
R4799 GND.n3852 GND.n3851 99.6594
R4800 GND.n3514 GND.n1909 99.6594
R4801 GND.n3518 GND.n1910 99.6594
R4802 GND.n3522 GND.n1911 99.6594
R4803 GND.n3526 GND.n1912 99.6594
R4804 GND.n3530 GND.n1913 99.6594
R4805 GND.n3534 GND.n1914 99.6594
R4806 GND.n3538 GND.n1915 99.6594
R4807 GND.n1917 GND.n1916 99.6594
R4808 GND.n3544 GND.n1906 99.6594
R4809 GND.n2598 GND.n2597 99.6594
R4810 GND.n2599 GND.n2591 99.6594
R4811 GND.n2608 GND.n2607 99.6594
R4812 GND.n2609 GND.n2587 99.6594
R4813 GND.n2618 GND.n2617 99.6594
R4814 GND.n2619 GND.n2580 99.6594
R4815 GND.n2628 GND.n2627 99.6594
R4816 GND.n2629 GND.n2576 99.6594
R4817 GND.n2638 GND.n2637 99.6594
R4818 GND.n2639 GND.n2572 99.6594
R4819 GND.n2649 GND.n2648 99.6594
R4820 GND.n2650 GND.n2566 99.6594
R4821 GND.n2659 GND.n2658 99.6594
R4822 GND.n2660 GND.n2562 99.6594
R4823 GND.n2669 GND.n2668 99.6594
R4824 GND.n2670 GND.n2558 99.6594
R4825 GND.n2679 GND.n2678 99.6594
R4826 GND.n2680 GND.n2554 99.6594
R4827 GND.n2691 GND.n2690 99.6594
R4828 GND.n2692 GND.n2550 99.6594
R4829 GND.n2701 GND.n2700 99.6594
R4830 GND.n2702 GND.n2546 99.6594
R4831 GND.n2711 GND.n2710 99.6594
R4832 GND.n2712 GND.n2542 99.6594
R4833 GND.n2721 GND.n2720 99.6594
R4834 GND.n1524 GND.n1523 99.6594
R4835 GND.n1518 GND.n1517 99.6594
R4836 GND.n1515 GND.n1512 99.6594
R4837 GND.n1510 GND.n1509 99.6594
R4838 GND.n1507 GND.n1504 99.6594
R4839 GND.n1502 GND.n1501 99.6594
R4840 GND.n1499 GND.n1496 99.6594
R4841 GND.n1494 GND.n1490 99.6594
R4842 GND.n1488 GND.n1487 99.6594
R4843 GND.n1483 GND.n1482 99.6594
R4844 GND.n1480 GND.n1479 99.6594
R4845 GND.n1475 GND.n1474 99.6594
R4846 GND.n1472 GND.n1468 99.6594
R4847 GND.n3913 GND.n3912 99.6594
R4848 GND.n1453 GND.n1447 99.6594
R4849 GND.n1455 GND.n1444 99.6594
R4850 GND.n1456 GND.n1442 99.6594
R4851 GND.n1458 GND.n1439 99.6594
R4852 GND.n1459 GND.n1437 99.6594
R4853 GND.n1460 GND.n1431 99.6594
R4854 GND.n1462 GND.n1461 99.6594
R4855 GND.n1463 GND.n1426 99.6594
R4856 GND.n1465 GND.n1464 99.6594
R4857 GND.n1466 GND.n1421 99.6594
R4858 GND.n3499 GND.n1978 99.6594
R4859 GND.n3491 GND.n1946 99.6594
R4860 GND.n3487 GND.n1947 99.6594
R4861 GND.n3483 GND.n1948 99.6594
R4862 GND.n3479 GND.n1949 99.6594
R4863 GND.n3475 GND.n1950 99.6594
R4864 GND.n3471 GND.n1951 99.6594
R4865 GND.n3467 GND.n1952 99.6594
R4866 GND.n3463 GND.n1953 99.6594
R4867 GND.n3459 GND.n1954 99.6594
R4868 GND.n3454 GND.n1956 99.6594
R4869 GND.n3450 GND.n1957 99.6594
R4870 GND.n3446 GND.n1958 99.6594
R4871 GND.n3442 GND.n1959 99.6594
R4872 GND.n3438 GND.n1960 99.6594
R4873 GND.n3434 GND.n1961 99.6594
R4874 GND.n2122 GND.n1962 99.6594
R4875 GND.n3427 GND.n1963 99.6594
R4876 GND.n3423 GND.n1964 99.6594
R4877 GND.n3419 GND.n1965 99.6594
R4878 GND.n3415 GND.n1966 99.6594
R4879 GND.n3411 GND.n1967 99.6594
R4880 GND.n2137 GND.n1968 99.6594
R4881 GND.n3403 GND.n1969 99.6594
R4882 GND.n155 GND.n70 99.6594
R4883 GND.n159 GND.n71 99.6594
R4884 GND.n163 GND.n72 99.6594
R4885 GND.n167 GND.n73 99.6594
R4886 GND.n171 GND.n74 99.6594
R4887 GND.n175 GND.n75 99.6594
R4888 GND.n137 GND.n76 99.6594
R4889 GND.n183 GND.n77 99.6594
R4890 GND.n187 GND.n78 99.6594
R4891 GND.n191 GND.n79 99.6594
R4892 GND.n195 GND.n80 99.6594
R4893 GND.n199 GND.n81 99.6594
R4894 GND.n203 GND.n82 99.6594
R4895 GND.n210 GND.n83 99.6594
R4896 GND.n214 GND.n84 99.6594
R4897 GND.n218 GND.n85 99.6594
R4898 GND.n222 GND.n86 99.6594
R4899 GND.n226 GND.n87 99.6594
R4900 GND.n230 GND.n88 99.6594
R4901 GND.n234 GND.n89 99.6594
R4902 GND.n238 GND.n90 99.6594
R4903 GND.n242 GND.n91 99.6594
R4904 GND.n246 GND.n92 99.6594
R4905 GND.n250 GND.n93 99.6594
R4906 GND.n95 GND.n94 99.6594
R4907 GND.n2733 GND.n2732 99.6594
R4908 GND.n2736 GND.n2735 99.6594
R4909 GND.n2743 GND.n2742 99.6594
R4910 GND.n2746 GND.n2745 99.6594
R4911 GND.n2753 GND.n2752 99.6594
R4912 GND.n2734 GND.n2733 99.6594
R4913 GND.n2735 GND.n2532 99.6594
R4914 GND.n2744 GND.n2743 99.6594
R4915 GND.n2745 GND.n2528 99.6594
R4916 GND.n2754 GND.n2753 99.6594
R4917 GND.n1536 GND.n1535 99.6594
R4918 GND.n2362 GND.n1538 99.6594
R4919 GND.n2365 GND.n2364 99.6594
R4920 GND.n2368 GND.n2367 99.6594
R4921 GND.n2373 GND.n2372 99.6594
R4922 GND.n2845 GND.n2375 99.6594
R4923 GND.n2846 GND.n2845 99.6594
R4924 GND.n2374 GND.n2373 99.6594
R4925 GND.n2369 GND.n2368 99.6594
R4926 GND.n2366 GND.n2365 99.6594
R4927 GND.n2363 GND.n2362 99.6594
R4928 GND.n1537 GND.n1536 99.6594
R4929 GND.n1620 GND.n1619 76.4039
R4930 GND.n1638 GND.t76 76.0312
R4931 GND.n2020 GND.t74 76.0312
R4932 GND.n1636 GND.t64 76.0294
R4933 GND.n2069 GND.t58 76.0294
R4934 GND.n3753 GND.n1452 75.3925
R4935 GND.n3456 GND.n2105 75.3925
R4936 GND.n2377 GND.t117 72.9043
R4937 GND.n1434 GND.t30 72.9043
R4938 GND.n1492 GND.t99 72.9043
R4939 GND.n1521 GND.t18 72.9043
R4940 GND.n1451 GND.t114 72.9043
R4941 GND.n1992 GND.t101 72.9043
R4942 GND.n2109 GND.t125 72.9043
R4943 GND.n2125 GND.t33 72.9043
R4944 GND.n2140 GND.t79 72.9043
R4945 GND.n151 GND.t111 72.9043
R4946 GND.n136 GND.t61 72.9043
R4947 GND.n207 GND.t54 72.9043
R4948 GND.n107 GND.t120 72.9043
R4949 GND.n3278 GND.t83 72.9043
R4950 GND.n2250 GND.t46 72.9043
R4951 GND.n2585 GND.t95 72.9043
R4952 GND.n2568 GND.t13 72.9043
R4953 GND.n2687 GND.t26 72.9043
R4954 GND.n2540 GND.t20 72.9043
R4955 GND.n2525 GND.t128 72.9043
R4956 GND.n1621 GND.n1613 72.8411
R4957 GND.n1630 GND.n1610 72.8411
R4958 GND.n1854 GND.n1853 72.8411
R4959 GND.n2101 GND.n2100 71.676
R4960 GND.n2096 GND.n2063 71.676
R4961 GND.n2092 GND.n2062 71.676
R4962 GND.n2088 GND.n2061 71.676
R4963 GND.n2084 GND.n2060 71.676
R4964 GND.n2080 GND.n2059 71.676
R4965 GND.n2075 GND.n2058 71.676
R4966 GND.n2071 GND.n2057 71.676
R4967 GND.n2104 GND.n2103 71.676
R4968 GND.n2023 GND.n2010 71.676
R4969 GND.n2027 GND.n2011 71.676
R4970 GND.n2031 GND.n2012 71.676
R4971 GND.n2035 GND.n2013 71.676
R4972 GND.n2039 GND.n2014 71.676
R4973 GND.n2043 GND.n2015 71.676
R4974 GND.n2047 GND.n2016 71.676
R4975 GND.n2050 GND.n2017 71.676
R4976 GND.n2056 GND.n2055 71.676
R4977 GND.n3789 GND.n3788 71.676
R4978 GND.n3783 GND.n1587 71.676
R4979 GND.n3780 GND.n1588 71.676
R4980 GND.n3776 GND.n1589 71.676
R4981 GND.n3772 GND.n1590 71.676
R4982 GND.n3768 GND.n1591 71.676
R4983 GND.n3764 GND.n1592 71.676
R4984 GND.n3759 GND.n1593 71.676
R4985 GND.n3755 GND.n1594 71.676
R4986 GND.n3749 GND.n1596 71.676
R4987 GND.n3745 GND.n1597 71.676
R4988 GND.n3740 GND.n1598 71.676
R4989 GND.n3736 GND.n1599 71.676
R4990 GND.n3732 GND.n1600 71.676
R4991 GND.n3728 GND.n1601 71.676
R4992 GND.n3724 GND.n1602 71.676
R4993 GND.n3720 GND.n1603 71.676
R4994 GND.n3789 GND.n1607 71.676
R4995 GND.n3781 GND.n1587 71.676
R4996 GND.n3777 GND.n1588 71.676
R4997 GND.n3773 GND.n1589 71.676
R4998 GND.n3769 GND.n1590 71.676
R4999 GND.n3765 GND.n1591 71.676
R5000 GND.n3760 GND.n1592 71.676
R5001 GND.n3756 GND.n1593 71.676
R5002 GND.n3750 GND.n1595 71.676
R5003 GND.n3746 GND.n1596 71.676
R5004 GND.n3741 GND.n1597 71.676
R5005 GND.n3737 GND.n1598 71.676
R5006 GND.n3733 GND.n1599 71.676
R5007 GND.n3729 GND.n1600 71.676
R5008 GND.n3725 GND.n1601 71.676
R5009 GND.n3721 GND.n1602 71.676
R5010 GND.n3717 GND.n1603 71.676
R5011 GND.n2056 GND.n2018 71.676
R5012 GND.n2048 GND.n2017 71.676
R5013 GND.n2044 GND.n2016 71.676
R5014 GND.n2040 GND.n2015 71.676
R5015 GND.n2036 GND.n2014 71.676
R5016 GND.n2032 GND.n2013 71.676
R5017 GND.n2028 GND.n2012 71.676
R5018 GND.n2024 GND.n2011 71.676
R5019 GND.n2010 GND.n2008 71.676
R5020 GND.n2070 GND.n2007 71.676
R5021 GND.n2074 GND.n2057 71.676
R5022 GND.n2079 GND.n2058 71.676
R5023 GND.n2083 GND.n2059 71.676
R5024 GND.n2087 GND.n2060 71.676
R5025 GND.n2091 GND.n2061 71.676
R5026 GND.n2095 GND.n2062 71.676
R5027 GND.n2065 GND.n2063 71.676
R5028 GND.n2101 GND.n2064 71.676
R5029 GND.n1636 GND.n1635 69.8187
R5030 GND.n1638 GND.n1637 69.8187
R5031 GND.n2020 GND.n2019 69.8187
R5032 GND.n2069 GND.n2068 69.8187
R5033 GND.n0 GND.t139 68.0267
R5034 GND.n5505 GND.t135 67.0052
R5035 GND.n3 GND.t141 65.3737
R5036 GND.n2 GND.t131 65.3112
R5037 GND.n1 GND.t132 65.3112
R5038 GND.n0 GND.t137 65.3112
R5039 GND.n5508 GND.t6 64.3522
R5040 GND.n5507 GND.t138 64.2897
R5041 GND.n5506 GND.t140 64.2897
R5042 GND.n5505 GND.t2 64.2897
R5043 GND.n4314 GND.n1029 62.2353
R5044 GND.n4308 GND.n1029 62.2353
R5045 GND.n4308 GND.n4307 62.2353
R5046 GND.n4307 GND.n4306 62.2353
R5047 GND.n4306 GND.n1036 62.2353
R5048 GND.n4300 GND.n1036 62.2353
R5049 GND.n4300 GND.n4299 62.2353
R5050 GND.n4299 GND.n4298 62.2353
R5051 GND.n4298 GND.n1044 62.2353
R5052 GND.n4292 GND.n1044 62.2353
R5053 GND.n4292 GND.n4291 62.2353
R5054 GND.n4291 GND.n4290 62.2353
R5055 GND.n4290 GND.n1052 62.2353
R5056 GND.n4284 GND.n1052 62.2353
R5057 GND.n4284 GND.n4283 62.2353
R5058 GND.n4283 GND.n4282 62.2353
R5059 GND.n4282 GND.n1060 62.2353
R5060 GND.n4276 GND.n1060 62.2353
R5061 GND.n4276 GND.n4275 62.2353
R5062 GND.n4275 GND.n4274 62.2353
R5063 GND.n4274 GND.n1068 62.2353
R5064 GND.n4268 GND.n1068 62.2353
R5065 GND.n4268 GND.n4267 62.2353
R5066 GND.n4267 GND.n4266 62.2353
R5067 GND.n4266 GND.n1076 62.2353
R5068 GND.n4260 GND.n1076 62.2353
R5069 GND.n4260 GND.n4259 62.2353
R5070 GND.n4259 GND.n4258 62.2353
R5071 GND.n4258 GND.n1084 62.2353
R5072 GND.n4252 GND.n1084 62.2353
R5073 GND.n4252 GND.n4251 62.2353
R5074 GND.n4251 GND.n4250 62.2353
R5075 GND.n4250 GND.n1092 62.2353
R5076 GND.n4244 GND.n1092 62.2353
R5077 GND.n4244 GND.n4243 62.2353
R5078 GND.n4243 GND.n4242 62.2353
R5079 GND.n4242 GND.n1100 62.2353
R5080 GND.n4236 GND.n1100 62.2353
R5081 GND.n4236 GND.n4235 62.2353
R5082 GND.n4235 GND.n4234 62.2353
R5083 GND.n4234 GND.n1108 62.2353
R5084 GND.n4228 GND.n1108 62.2353
R5085 GND.n4228 GND.n4227 62.2353
R5086 GND.n4227 GND.n4226 62.2353
R5087 GND.n4226 GND.n1116 62.2353
R5088 GND.n4220 GND.n1116 62.2353
R5089 GND.n4220 GND.n4219 62.2353
R5090 GND.n4219 GND.n4218 62.2353
R5091 GND.n4218 GND.n1124 62.2353
R5092 GND.n4212 GND.n1124 62.2353
R5093 GND.n4212 GND.n4211 62.2353
R5094 GND.n4211 GND.n4210 62.2353
R5095 GND.n4210 GND.n1132 62.2353
R5096 GND.n4204 GND.n1132 62.2353
R5097 GND.n1634 GND.n1633 62.0895
R5098 GND.n3762 GND.n1636 59.5399
R5099 GND.n3743 GND.n1638 59.5399
R5100 GND.n2021 GND.n2020 59.5399
R5101 GND.n2077 GND.n2069 59.5399
R5102 GND.n4203 GND.n4202 56.1286
R5103 GND.n5259 GND.n5258 56.1286
R5104 GND.n1618 GND.n1617 54.358
R5105 GND.n1851 GND.n1850 54.358
R5106 GND.n1840 GND.n1839 52.9692
R5107 GND.n1932 GND.n1931 50.4247
R5108 GND.n3863 GND.n3862 50.4247
R5109 GND.n1630 GND.n1629 46.0096
R5110 GND.n1623 GND.n1613 46.0096
R5111 GND.n1838 GND.n1837 46.0096
R5112 GND.n1854 GND.n1835 46.0096
R5113 GND.n2377 GND.n2376 45.9641
R5114 GND.n1434 GND.n1433 45.9641
R5115 GND.n1492 GND.n1491 45.9641
R5116 GND.n1521 GND.n1520 45.9641
R5117 GND.n1451 GND.n1450 45.9641
R5118 GND.n1992 GND.n1991 45.9641
R5119 GND.n2109 GND.n2108 45.9641
R5120 GND.n2125 GND.n2124 45.9641
R5121 GND.n2140 GND.n2139 45.9641
R5122 GND.n151 GND.n150 45.9641
R5123 GND.n136 GND.n135 45.9641
R5124 GND.n207 GND.n206 45.9641
R5125 GND.n107 GND.n106 45.9641
R5126 GND.n3278 GND.n3277 45.9641
R5127 GND.n2250 GND.n2249 45.9641
R5128 GND.n2585 GND.n2584 45.9641
R5129 GND.n2568 GND.n2567 45.9641
R5130 GND.n2687 GND.n2686 45.9641
R5131 GND.n2540 GND.n2539 45.9641
R5132 GND.n2525 GND.n2524 45.9641
R5133 GND.n1858 GND.n1857 44.3322
R5134 GND.n2848 GND.n2377 42.2793
R5135 GND.n1435 GND.n1434 42.2793
R5136 GND.n3890 GND.n1492 42.2793
R5137 GND.n3871 GND.n1521 42.2793
R5138 GND.n1993 GND.n1992 42.2793
R5139 GND.n3431 GND.n2125 42.2793
R5140 GND.n2141 GND.n2140 42.2793
R5141 GND.n154 GND.n151 42.2793
R5142 GND.n181 GND.n136 42.2793
R5143 GND.n208 GND.n207 42.2793
R5144 GND.n108 GND.n107 42.2793
R5145 GND.n3279 GND.n3278 42.2793
R5146 GND.n3231 GND.n2250 42.2793
R5147 GND.n1933 GND.n1932 42.2793
R5148 GND.n3864 GND.n3863 42.2793
R5149 GND.n2586 GND.n2585 42.2793
R5150 GND.n2569 GND.n2568 42.2793
R5151 GND.n2688 GND.n2687 42.2793
R5152 GND.n2541 GND.n2540 42.2793
R5153 GND.n2526 GND.n2525 42.2793
R5154 GND.n1620 GND.n1618 41.6274
R5155 GND.n1852 GND.n1851 41.6274
R5156 GND.n1619 GND.n1613 38.2165
R5157 GND.n2054 GND.n2053 36.9956
R5158 GND.n3716 GND.n3715 36.9956
R5159 GND.n1452 GND.n1451 36.9518
R5160 GND.n3456 GND.n2109 36.9518
R5161 GND.n4202 GND.n1140 36.6855
R5162 GND.n4196 GND.n1140 36.6855
R5163 GND.n4196 GND.n4195 36.6855
R5164 GND.n4195 GND.n4194 36.6855
R5165 GND.n4194 GND.n1148 36.6855
R5166 GND.n4188 GND.n1148 36.6855
R5167 GND.n4188 GND.n4187 36.6855
R5168 GND.n4187 GND.n4186 36.6855
R5169 GND.n4186 GND.n1156 36.6855
R5170 GND.n4180 GND.n1156 36.6855
R5171 GND.n4180 GND.n4179 36.6855
R5172 GND.n4179 GND.n4178 36.6855
R5173 GND.n4178 GND.n1164 36.6855
R5174 GND.n4172 GND.n1164 36.6855
R5175 GND.n4172 GND.n4171 36.6855
R5176 GND.n4171 GND.n4170 36.6855
R5177 GND.n4170 GND.n1172 36.6855
R5178 GND.n4164 GND.n1172 36.6855
R5179 GND.n4164 GND.n4163 36.6855
R5180 GND.n4163 GND.n4162 36.6855
R5181 GND.n4162 GND.n1180 36.6855
R5182 GND.n4156 GND.n1180 36.6855
R5183 GND.n4156 GND.n4155 36.6855
R5184 GND.n4155 GND.n4154 36.6855
R5185 GND.n4154 GND.n1188 36.6855
R5186 GND.n4148 GND.n1188 36.6855
R5187 GND.n4148 GND.n4147 36.6855
R5188 GND.n4147 GND.n4146 36.6855
R5189 GND.n4146 GND.n1196 36.6855
R5190 GND.n4140 GND.n1196 36.6855
R5191 GND.n4140 GND.n4139 36.6855
R5192 GND.n4139 GND.n4138 36.6855
R5193 GND.n4138 GND.n1204 36.6855
R5194 GND.n4132 GND.n1204 36.6855
R5195 GND.n4132 GND.n4131 36.6855
R5196 GND.n4131 GND.n4130 36.6855
R5197 GND.n4130 GND.n1212 36.6855
R5198 GND.n4124 GND.n1212 36.6855
R5199 GND.n4124 GND.n4123 36.6855
R5200 GND.n4123 GND.n4122 36.6855
R5201 GND.n4122 GND.n1220 36.6855
R5202 GND.n4116 GND.n1220 36.6855
R5203 GND.n4116 GND.n4115 36.6855
R5204 GND.n4115 GND.n4114 36.6855
R5205 GND.n4114 GND.n1228 36.6855
R5206 GND.n4108 GND.n1228 36.6855
R5207 GND.n4108 GND.n4107 36.6855
R5208 GND.n4107 GND.n4106 36.6855
R5209 GND.n4106 GND.n1236 36.6855
R5210 GND.n4100 GND.n1236 36.6855
R5211 GND.n4100 GND.n4099 36.6855
R5212 GND.n4099 GND.n4098 36.6855
R5213 GND.n4098 GND.n1244 36.6855
R5214 GND.n4092 GND.n1244 36.6855
R5215 GND.n4092 GND.n4091 36.6855
R5216 GND.n4091 GND.n4090 36.6855
R5217 GND.n4090 GND.n1252 36.6855
R5218 GND.n4084 GND.n1252 36.6855
R5219 GND.n4084 GND.n4083 36.6855
R5220 GND.n4083 GND.n4082 36.6855
R5221 GND.n4082 GND.n1260 36.6855
R5222 GND.n4076 GND.n1260 36.6855
R5223 GND.n4076 GND.n4075 36.6855
R5224 GND.n4075 GND.n4074 36.6855
R5225 GND.n4074 GND.n1268 36.6855
R5226 GND.n4068 GND.n1268 36.6855
R5227 GND.n4068 GND.n4067 36.6855
R5228 GND.n4067 GND.n4066 36.6855
R5229 GND.n4066 GND.n1276 36.6855
R5230 GND.n4060 GND.n1276 36.6855
R5231 GND.n4060 GND.n4059 36.6855
R5232 GND.n4059 GND.n4058 36.6855
R5233 GND.n4058 GND.n1284 36.6855
R5234 GND.n4052 GND.n1284 36.6855
R5235 GND.n4052 GND.n4051 36.6855
R5236 GND.n4051 GND.n4050 36.6855
R5237 GND.n4050 GND.n1292 36.6855
R5238 GND.n4044 GND.n1292 36.6855
R5239 GND.n4044 GND.n4043 36.6855
R5240 GND.n4043 GND.n4042 36.6855
R5241 GND.n4042 GND.n1300 36.6855
R5242 GND.n4036 GND.n1300 36.6855
R5243 GND.n4036 GND.n4035 36.6855
R5244 GND.n4035 GND.n4034 36.6855
R5245 GND.n4034 GND.n1308 36.6855
R5246 GND.n4028 GND.n1308 36.6855
R5247 GND.n4028 GND.n4027 36.6855
R5248 GND.n4027 GND.n4026 36.6855
R5249 GND.n4026 GND.n1316 36.6855
R5250 GND.n4020 GND.n1316 36.6855
R5251 GND.n4020 GND.n4019 36.6855
R5252 GND.n4019 GND.n4018 36.6855
R5253 GND.n4018 GND.n1324 36.6855
R5254 GND.n4012 GND.n1324 36.6855
R5255 GND.n4012 GND.n4011 36.6855
R5256 GND.n4011 GND.n4010 36.6855
R5257 GND.n4010 GND.n1332 36.6855
R5258 GND.n4004 GND.n1332 36.6855
R5259 GND.n4004 GND.n4003 36.6855
R5260 GND.n4003 GND.n4002 36.6855
R5261 GND.n4002 GND.n1340 36.6855
R5262 GND.n3996 GND.n1340 36.6855
R5263 GND.n3996 GND.n3995 36.6855
R5264 GND.n3995 GND.n3994 36.6855
R5265 GND.n3988 GND.n1356 36.6855
R5266 GND.n2484 GND.n1413 36.6855
R5267 GND.n2482 GND.n1543 36.6855
R5268 GND.n2476 GND.n1551 36.6855
R5269 GND.n3508 GND.n1907 36.6855
R5270 GND.n3501 GND.n1908 36.6855
R5271 GND.n2146 GND.n1976 36.6855
R5272 GND.n5473 GND.n61 36.6855
R5273 GND.n5467 GND.n5466 36.6855
R5274 GND.n5466 GND.n5465 36.6855
R5275 GND.n5465 GND.n259 36.6855
R5276 GND.n5459 GND.n259 36.6855
R5277 GND.n5459 GND.n5458 36.6855
R5278 GND.n5458 GND.n5457 36.6855
R5279 GND.n5457 GND.n267 36.6855
R5280 GND.n5451 GND.n267 36.6855
R5281 GND.n5451 GND.n5450 36.6855
R5282 GND.n5450 GND.n5449 36.6855
R5283 GND.n5449 GND.n275 36.6855
R5284 GND.n5443 GND.n275 36.6855
R5285 GND.n5443 GND.n5442 36.6855
R5286 GND.n5442 GND.n5441 36.6855
R5287 GND.n5441 GND.n283 36.6855
R5288 GND.n5435 GND.n283 36.6855
R5289 GND.n5435 GND.n5434 36.6855
R5290 GND.n5434 GND.n5433 36.6855
R5291 GND.n5433 GND.n291 36.6855
R5292 GND.n5427 GND.n291 36.6855
R5293 GND.n5427 GND.n5426 36.6855
R5294 GND.n5426 GND.n5425 36.6855
R5295 GND.n5425 GND.n299 36.6855
R5296 GND.n5419 GND.n299 36.6855
R5297 GND.n5419 GND.n5418 36.6855
R5298 GND.n5418 GND.n5417 36.6855
R5299 GND.n5417 GND.n307 36.6855
R5300 GND.n5411 GND.n307 36.6855
R5301 GND.n5411 GND.n5410 36.6855
R5302 GND.n5410 GND.n5409 36.6855
R5303 GND.n5409 GND.n315 36.6855
R5304 GND.n5403 GND.n315 36.6855
R5305 GND.n5403 GND.n5402 36.6855
R5306 GND.n5402 GND.n5401 36.6855
R5307 GND.n5401 GND.n323 36.6855
R5308 GND.n5395 GND.n323 36.6855
R5309 GND.n5395 GND.n5394 36.6855
R5310 GND.n5394 GND.n5393 36.6855
R5311 GND.n5393 GND.n331 36.6855
R5312 GND.n5387 GND.n331 36.6855
R5313 GND.n5387 GND.n5386 36.6855
R5314 GND.n5386 GND.n5385 36.6855
R5315 GND.n5385 GND.n339 36.6855
R5316 GND.n5379 GND.n339 36.6855
R5317 GND.n5379 GND.n5378 36.6855
R5318 GND.n5378 GND.n5377 36.6855
R5319 GND.n5377 GND.n347 36.6855
R5320 GND.n5371 GND.n347 36.6855
R5321 GND.n5371 GND.n5370 36.6855
R5322 GND.n5370 GND.n5369 36.6855
R5323 GND.n5369 GND.n355 36.6855
R5324 GND.n5363 GND.n355 36.6855
R5325 GND.n5363 GND.n5362 36.6855
R5326 GND.n5362 GND.n5361 36.6855
R5327 GND.n5361 GND.n363 36.6855
R5328 GND.n5355 GND.n363 36.6855
R5329 GND.n5355 GND.n5354 36.6855
R5330 GND.n5354 GND.n5353 36.6855
R5331 GND.n5353 GND.n371 36.6855
R5332 GND.n5347 GND.n371 36.6855
R5333 GND.n5347 GND.n5346 36.6855
R5334 GND.n5346 GND.n5345 36.6855
R5335 GND.n5345 GND.n379 36.6855
R5336 GND.n5339 GND.n379 36.6855
R5337 GND.n5339 GND.n5338 36.6855
R5338 GND.n5338 GND.n5337 36.6855
R5339 GND.n5337 GND.n387 36.6855
R5340 GND.n5331 GND.n387 36.6855
R5341 GND.n5331 GND.n5330 36.6855
R5342 GND.n5330 GND.n5329 36.6855
R5343 GND.n5329 GND.n395 36.6855
R5344 GND.n5323 GND.n395 36.6855
R5345 GND.n5323 GND.n5322 36.6855
R5346 GND.n5322 GND.n5321 36.6855
R5347 GND.n5321 GND.n403 36.6855
R5348 GND.n5315 GND.n403 36.6855
R5349 GND.n5315 GND.n5314 36.6855
R5350 GND.n5314 GND.n5313 36.6855
R5351 GND.n5313 GND.n411 36.6855
R5352 GND.n5307 GND.n411 36.6855
R5353 GND.n5307 GND.n5306 36.6855
R5354 GND.n5306 GND.n5305 36.6855
R5355 GND.n5305 GND.n419 36.6855
R5356 GND.n5299 GND.n419 36.6855
R5357 GND.n5299 GND.n5298 36.6855
R5358 GND.n5298 GND.n5297 36.6855
R5359 GND.n5297 GND.n427 36.6855
R5360 GND.n5291 GND.n427 36.6855
R5361 GND.n5291 GND.n5290 36.6855
R5362 GND.n5290 GND.n5289 36.6855
R5363 GND.n5289 GND.n435 36.6855
R5364 GND.n5283 GND.n435 36.6855
R5365 GND.n5283 GND.n5282 36.6855
R5366 GND.n5282 GND.n5281 36.6855
R5367 GND.n5281 GND.n443 36.6855
R5368 GND.n5275 GND.n443 36.6855
R5369 GND.n5275 GND.n5274 36.6855
R5370 GND.n5274 GND.n5273 36.6855
R5371 GND.n5273 GND.n451 36.6855
R5372 GND.n5267 GND.n451 36.6855
R5373 GND.n5267 GND.n5266 36.6855
R5374 GND.n5266 GND.n5265 36.6855
R5375 GND.n5265 GND.n459 36.6855
R5376 GND.n5259 GND.n459 36.6855
R5377 GND.n3850 GND.n1543 34.4844
R5378 GND.n3545 GND.n1908 34.4844
R5379 GND.n2482 GND.n1467 34.1176
R5380 GND.n3501 GND.n3500 34.1176
R5381 GND.n3987 GND.n1359 33.017
R5382 GND.n2761 GND.n1368 33.017
R5383 GND.n2518 GND.n2437 33.017
R5384 GND.n2771 GND.n2433 33.017
R5385 GND.n2776 GND.n2436 33.017
R5386 GND.n2773 GND.n2422 33.017
R5387 GND.n2785 GND.n2423 33.017
R5388 GND.n2427 GND.n2414 33.017
R5389 GND.n2801 GND.n2412 33.017
R5390 GND.n2798 GND.n2401 33.017
R5391 GND.n2810 GND.n2402 33.017
R5392 GND.n2406 GND.n2394 33.017
R5393 GND.n2824 GND.n2390 33.017
R5394 GND.n2828 GND.n2392 33.017
R5395 GND.n2836 GND.n2381 33.017
R5396 GND.n2839 GND.n1411 33.017
R5397 GND.n3950 GND.n1413 33.017
R5398 GND.n3401 GND.n2146 33.017
R5399 GND.n2246 GND.n2148 33.017
R5400 GND.n3393 GND.n2156 33.017
R5401 GND.n3387 GND.n2170 33.017
R5402 GND.n3254 GND.n2173 33.017
R5403 GND.n3381 GND.n2183 33.017
R5404 GND.n3377 GND.n2186 33.017
R5405 GND.n3376 GND.n2191 33.017
R5406 GND.n3368 GND.n2221 33.017
R5407 GND.n3362 GND.n12 33.017
R5408 GND.n3361 GND.n2233 33.017
R5409 GND.n3339 GND.n3338 33.017
R5410 GND.n5493 GND.n29 33.017
R5411 GND.n3332 GND.n32 33.017
R5412 GND.n5487 GND.n41 33.017
R5413 GND.n5481 GND.n51 33.017
R5414 GND.n5474 GND.n54 33.017
R5415 GND.n1356 GND.n1348 31.9165
R5416 GND.n258 GND.n61 31.9165
R5417 GND.n1631 GND.n1630 29.9429
R5418 GND.n1855 GND.n1854 29.9429
R5419 GND.n1625 GND.n1611 24.1005
R5420 GND.n1625 GND.n1624 24.1005
R5421 GND.n1843 GND.n1842 24.1005
R5422 GND.n1844 GND.n1843 24.1005
R5423 GND.n2901 GND.n1634 22.3225
R5424 GND.n3577 GND.n1858 22.3225
R5425 GND.n3981 GND.t12 21.2778
R5426 GND.n3326 GND.t52 21.2778
R5427 GND.n1616 GND.t123 19.8005
R5428 GND.n1616 GND.t50 19.8005
R5429 GND.n1615 GND.t10 19.8005
R5430 GND.n1615 GND.t71 19.8005
R5431 GND.n1614 GND.t108 19.8005
R5432 GND.n1614 GND.t24 19.8005
R5433 GND.n1849 GND.t86 19.8005
R5434 GND.n1849 GND.t68 19.8005
R5435 GND.n1848 GND.t105 19.8005
R5436 GND.n1848 GND.t44 19.8005
R5437 GND.n1847 GND.t93 19.8005
R5438 GND.n1847 GND.t37 19.8005
R5439 GND.n1610 GND.n1609 19.5087
R5440 GND.n1628 GND.n1610 19.5087
R5441 GND.n1622 GND.n1621 19.5087
R5442 GND.n1853 GND.n1846 19.5087
R5443 GND.n3857 GND.n1534 19.3944
R5444 GND.n3857 GND.n3856 19.3944
R5445 GND.n3856 GND.n1539 19.3944
R5446 GND.n2361 GND.n1539 19.3944
R5447 GND.n2856 GND.n2361 19.3944
R5448 GND.n2856 GND.n2855 19.3944
R5449 GND.n2855 GND.n2854 19.3944
R5450 GND.n2854 GND.n2370 19.3944
R5451 GND.n2850 GND.n2370 19.3944
R5452 GND.n2850 GND.n2849 19.3944
R5453 GND.n2725 GND.n1373 19.3944
R5454 GND.n3979 GND.n1373 19.3944
R5455 GND.n3979 GND.n1374 19.3944
R5456 GND.n1381 GND.n1374 19.3944
R5457 GND.n1382 GND.n1381 19.3944
R5458 GND.n1383 GND.n1382 19.3944
R5459 GND.n2424 GND.n1383 19.3944
R5460 GND.n2424 GND.n1389 19.3944
R5461 GND.n1390 GND.n1389 19.3944
R5462 GND.n1391 GND.n1390 19.3944
R5463 GND.n2797 GND.n1391 19.3944
R5464 GND.n2797 GND.n1397 19.3944
R5465 GND.n1398 GND.n1397 19.3944
R5466 GND.n1399 GND.n1398 19.3944
R5467 GND.n2826 GND.n1399 19.3944
R5468 GND.n2826 GND.n1405 19.3944
R5469 GND.n1406 GND.n1405 19.3944
R5470 GND.n1407 GND.n1406 19.3944
R5471 GND.n1414 GND.n1407 19.3944
R5472 GND.n2726 GND.n1377 19.3944
R5473 GND.n3977 GND.n1377 19.3944
R5474 GND.n3977 GND.n3976 19.3944
R5475 GND.n3976 GND.n3975 19.3944
R5476 GND.n3975 GND.n1380 19.3944
R5477 GND.n3971 GND.n1380 19.3944
R5478 GND.n3971 GND.n3970 19.3944
R5479 GND.n3970 GND.n3969 19.3944
R5480 GND.n3969 GND.n1388 19.3944
R5481 GND.n3965 GND.n1388 19.3944
R5482 GND.n3965 GND.n3964 19.3944
R5483 GND.n3964 GND.n3963 19.3944
R5484 GND.n3963 GND.n1396 19.3944
R5485 GND.n3959 GND.n1396 19.3944
R5486 GND.n3959 GND.n3958 19.3944
R5487 GND.n3958 GND.n3957 19.3944
R5488 GND.n3957 GND.n1404 19.3944
R5489 GND.n3953 GND.n1404 19.3944
R5490 GND.n3953 GND.n3952 19.3944
R5491 GND.n3945 GND.n3944 19.3944
R5492 GND.n3944 GND.n3943 19.3944
R5493 GND.n3943 GND.n1423 19.3944
R5494 GND.n3939 GND.n1423 19.3944
R5495 GND.n3939 GND.n3938 19.3944
R5496 GND.n3938 GND.n3937 19.3944
R5497 GND.n3937 GND.n1428 19.3944
R5498 GND.n3933 GND.n1428 19.3944
R5499 GND.n3933 GND.n3932 19.3944
R5500 GND.n3932 GND.n3931 19.3944
R5501 GND.n3928 GND.n3927 19.3944
R5502 GND.n3927 GND.n3926 19.3944
R5503 GND.n3926 GND.n1440 19.3944
R5504 GND.n3922 GND.n1440 19.3944
R5505 GND.n3922 GND.n3921 19.3944
R5506 GND.n3921 GND.n3920 19.3944
R5507 GND.n3920 GND.n1445 19.3944
R5508 GND.n3916 GND.n1445 19.3944
R5509 GND.n3916 GND.n3915 19.3944
R5510 GND.n3915 GND.n3914 19.3944
R5511 GND.n3908 GND.n1469 19.3944
R5512 GND.n3904 GND.n1469 19.3944
R5513 GND.n3904 GND.n3903 19.3944
R5514 GND.n3903 GND.n3902 19.3944
R5515 GND.n3902 GND.n1477 19.3944
R5516 GND.n3898 GND.n1477 19.3944
R5517 GND.n3898 GND.n3897 19.3944
R5518 GND.n3897 GND.n3896 19.3944
R5519 GND.n3896 GND.n1485 19.3944
R5520 GND.n3892 GND.n1485 19.3944
R5521 GND.n3892 GND.n3891 19.3944
R5522 GND.n3889 GND.n1497 19.3944
R5523 GND.n3885 GND.n1497 19.3944
R5524 GND.n3885 GND.n3884 19.3944
R5525 GND.n3884 GND.n3883 19.3944
R5526 GND.n3883 GND.n1505 19.3944
R5527 GND.n3879 GND.n1505 19.3944
R5528 GND.n3879 GND.n3878 19.3944
R5529 GND.n3878 GND.n3877 19.3944
R5530 GND.n3877 GND.n1513 19.3944
R5531 GND.n3873 GND.n1513 19.3944
R5532 GND.n3873 GND.n3872 19.3944
R5533 GND.n5119 GND.n546 19.3944
R5534 GND.n5123 GND.n546 19.3944
R5535 GND.n5123 GND.n542 19.3944
R5536 GND.n5129 GND.n542 19.3944
R5537 GND.n5129 GND.n540 19.3944
R5538 GND.n5133 GND.n540 19.3944
R5539 GND.n5133 GND.n536 19.3944
R5540 GND.n5139 GND.n536 19.3944
R5541 GND.n5139 GND.n534 19.3944
R5542 GND.n5143 GND.n534 19.3944
R5543 GND.n5143 GND.n530 19.3944
R5544 GND.n5149 GND.n530 19.3944
R5545 GND.n5149 GND.n528 19.3944
R5546 GND.n5153 GND.n528 19.3944
R5547 GND.n5153 GND.n524 19.3944
R5548 GND.n5159 GND.n524 19.3944
R5549 GND.n5159 GND.n522 19.3944
R5550 GND.n5163 GND.n522 19.3944
R5551 GND.n5163 GND.n518 19.3944
R5552 GND.n5169 GND.n518 19.3944
R5553 GND.n5169 GND.n516 19.3944
R5554 GND.n5173 GND.n516 19.3944
R5555 GND.n5173 GND.n512 19.3944
R5556 GND.n5179 GND.n512 19.3944
R5557 GND.n5179 GND.n510 19.3944
R5558 GND.n5183 GND.n510 19.3944
R5559 GND.n5183 GND.n506 19.3944
R5560 GND.n5189 GND.n506 19.3944
R5561 GND.n5189 GND.n504 19.3944
R5562 GND.n5193 GND.n504 19.3944
R5563 GND.n5193 GND.n500 19.3944
R5564 GND.n5199 GND.n500 19.3944
R5565 GND.n5199 GND.n498 19.3944
R5566 GND.n5203 GND.n498 19.3944
R5567 GND.n5203 GND.n494 19.3944
R5568 GND.n5209 GND.n494 19.3944
R5569 GND.n5209 GND.n492 19.3944
R5570 GND.n5213 GND.n492 19.3944
R5571 GND.n5213 GND.n488 19.3944
R5572 GND.n5219 GND.n488 19.3944
R5573 GND.n5219 GND.n486 19.3944
R5574 GND.n5223 GND.n486 19.3944
R5575 GND.n5223 GND.n482 19.3944
R5576 GND.n5229 GND.n482 19.3944
R5577 GND.n5229 GND.n480 19.3944
R5578 GND.n5233 GND.n480 19.3944
R5579 GND.n5233 GND.n476 19.3944
R5580 GND.n5239 GND.n476 19.3944
R5581 GND.n5239 GND.n474 19.3944
R5582 GND.n5243 GND.n474 19.3944
R5583 GND.n5243 GND.n470 19.3944
R5584 GND.n5249 GND.n470 19.3944
R5585 GND.n5249 GND.n468 19.3944
R5586 GND.n5255 GND.n468 19.3944
R5587 GND.n5255 GND.n5254 19.3944
R5588 GND.n4318 GND.n1027 19.3944
R5589 GND.n4318 GND.n1025 19.3944
R5590 GND.n4322 GND.n1025 19.3944
R5591 GND.n4322 GND.n1021 19.3944
R5592 GND.n4328 GND.n1021 19.3944
R5593 GND.n4328 GND.n1019 19.3944
R5594 GND.n4332 GND.n1019 19.3944
R5595 GND.n4332 GND.n1015 19.3944
R5596 GND.n4338 GND.n1015 19.3944
R5597 GND.n4338 GND.n1013 19.3944
R5598 GND.n4342 GND.n1013 19.3944
R5599 GND.n4342 GND.n1009 19.3944
R5600 GND.n4348 GND.n1009 19.3944
R5601 GND.n4348 GND.n1007 19.3944
R5602 GND.n4352 GND.n1007 19.3944
R5603 GND.n4352 GND.n1003 19.3944
R5604 GND.n4358 GND.n1003 19.3944
R5605 GND.n4358 GND.n1001 19.3944
R5606 GND.n4362 GND.n1001 19.3944
R5607 GND.n4362 GND.n997 19.3944
R5608 GND.n4368 GND.n997 19.3944
R5609 GND.n4368 GND.n995 19.3944
R5610 GND.n4372 GND.n995 19.3944
R5611 GND.n4372 GND.n991 19.3944
R5612 GND.n4378 GND.n991 19.3944
R5613 GND.n4378 GND.n989 19.3944
R5614 GND.n4382 GND.n989 19.3944
R5615 GND.n4382 GND.n985 19.3944
R5616 GND.n4388 GND.n985 19.3944
R5617 GND.n4388 GND.n983 19.3944
R5618 GND.n4392 GND.n983 19.3944
R5619 GND.n4392 GND.n979 19.3944
R5620 GND.n4398 GND.n979 19.3944
R5621 GND.n4398 GND.n977 19.3944
R5622 GND.n4402 GND.n977 19.3944
R5623 GND.n4402 GND.n973 19.3944
R5624 GND.n4408 GND.n973 19.3944
R5625 GND.n4408 GND.n971 19.3944
R5626 GND.n4412 GND.n971 19.3944
R5627 GND.n4412 GND.n967 19.3944
R5628 GND.n4418 GND.n967 19.3944
R5629 GND.n4418 GND.n965 19.3944
R5630 GND.n4422 GND.n965 19.3944
R5631 GND.n4422 GND.n961 19.3944
R5632 GND.n4428 GND.n961 19.3944
R5633 GND.n4428 GND.n959 19.3944
R5634 GND.n4432 GND.n959 19.3944
R5635 GND.n4432 GND.n955 19.3944
R5636 GND.n4438 GND.n955 19.3944
R5637 GND.n4438 GND.n953 19.3944
R5638 GND.n4442 GND.n953 19.3944
R5639 GND.n4442 GND.n949 19.3944
R5640 GND.n4448 GND.n949 19.3944
R5641 GND.n4448 GND.n947 19.3944
R5642 GND.n4452 GND.n947 19.3944
R5643 GND.n4452 GND.n943 19.3944
R5644 GND.n4458 GND.n943 19.3944
R5645 GND.n4458 GND.n941 19.3944
R5646 GND.n4462 GND.n941 19.3944
R5647 GND.n4462 GND.n937 19.3944
R5648 GND.n4468 GND.n937 19.3944
R5649 GND.n4468 GND.n935 19.3944
R5650 GND.n4472 GND.n935 19.3944
R5651 GND.n4472 GND.n931 19.3944
R5652 GND.n4478 GND.n931 19.3944
R5653 GND.n4478 GND.n929 19.3944
R5654 GND.n4482 GND.n929 19.3944
R5655 GND.n4482 GND.n925 19.3944
R5656 GND.n4488 GND.n925 19.3944
R5657 GND.n4488 GND.n923 19.3944
R5658 GND.n4492 GND.n923 19.3944
R5659 GND.n4492 GND.n919 19.3944
R5660 GND.n4498 GND.n919 19.3944
R5661 GND.n4498 GND.n917 19.3944
R5662 GND.n4502 GND.n917 19.3944
R5663 GND.n4502 GND.n913 19.3944
R5664 GND.n4508 GND.n913 19.3944
R5665 GND.n4508 GND.n911 19.3944
R5666 GND.n4512 GND.n911 19.3944
R5667 GND.n4512 GND.n907 19.3944
R5668 GND.n4518 GND.n907 19.3944
R5669 GND.n4518 GND.n905 19.3944
R5670 GND.n4522 GND.n905 19.3944
R5671 GND.n4522 GND.n901 19.3944
R5672 GND.n4528 GND.n901 19.3944
R5673 GND.n4528 GND.n899 19.3944
R5674 GND.n4532 GND.n899 19.3944
R5675 GND.n4532 GND.n895 19.3944
R5676 GND.n4538 GND.n895 19.3944
R5677 GND.n4538 GND.n893 19.3944
R5678 GND.n4542 GND.n893 19.3944
R5679 GND.n4542 GND.n889 19.3944
R5680 GND.n4548 GND.n889 19.3944
R5681 GND.n4548 GND.n887 19.3944
R5682 GND.n4552 GND.n887 19.3944
R5683 GND.n4552 GND.n883 19.3944
R5684 GND.n4558 GND.n883 19.3944
R5685 GND.n4558 GND.n881 19.3944
R5686 GND.n4562 GND.n881 19.3944
R5687 GND.n4562 GND.n877 19.3944
R5688 GND.n4568 GND.n877 19.3944
R5689 GND.n4568 GND.n875 19.3944
R5690 GND.n4572 GND.n875 19.3944
R5691 GND.n4572 GND.n871 19.3944
R5692 GND.n4578 GND.n871 19.3944
R5693 GND.n4578 GND.n869 19.3944
R5694 GND.n4582 GND.n869 19.3944
R5695 GND.n4582 GND.n865 19.3944
R5696 GND.n4588 GND.n865 19.3944
R5697 GND.n4588 GND.n863 19.3944
R5698 GND.n4592 GND.n863 19.3944
R5699 GND.n4592 GND.n859 19.3944
R5700 GND.n4598 GND.n859 19.3944
R5701 GND.n4598 GND.n857 19.3944
R5702 GND.n4602 GND.n857 19.3944
R5703 GND.n4602 GND.n853 19.3944
R5704 GND.n4608 GND.n853 19.3944
R5705 GND.n4608 GND.n851 19.3944
R5706 GND.n4612 GND.n851 19.3944
R5707 GND.n4612 GND.n847 19.3944
R5708 GND.n4618 GND.n847 19.3944
R5709 GND.n4618 GND.n845 19.3944
R5710 GND.n4622 GND.n845 19.3944
R5711 GND.n4622 GND.n841 19.3944
R5712 GND.n4628 GND.n841 19.3944
R5713 GND.n4628 GND.n839 19.3944
R5714 GND.n4632 GND.n839 19.3944
R5715 GND.n4632 GND.n835 19.3944
R5716 GND.n4638 GND.n835 19.3944
R5717 GND.n4638 GND.n833 19.3944
R5718 GND.n4642 GND.n833 19.3944
R5719 GND.n4642 GND.n829 19.3944
R5720 GND.n4648 GND.n829 19.3944
R5721 GND.n4648 GND.n827 19.3944
R5722 GND.n4652 GND.n827 19.3944
R5723 GND.n4652 GND.n823 19.3944
R5724 GND.n4658 GND.n823 19.3944
R5725 GND.n4658 GND.n821 19.3944
R5726 GND.n4662 GND.n821 19.3944
R5727 GND.n4662 GND.n817 19.3944
R5728 GND.n4668 GND.n817 19.3944
R5729 GND.n4668 GND.n815 19.3944
R5730 GND.n4672 GND.n815 19.3944
R5731 GND.n4672 GND.n811 19.3944
R5732 GND.n4678 GND.n811 19.3944
R5733 GND.n4678 GND.n809 19.3944
R5734 GND.n4682 GND.n809 19.3944
R5735 GND.n4682 GND.n805 19.3944
R5736 GND.n4688 GND.n805 19.3944
R5737 GND.n4688 GND.n803 19.3944
R5738 GND.n4692 GND.n803 19.3944
R5739 GND.n4692 GND.n799 19.3944
R5740 GND.n4698 GND.n799 19.3944
R5741 GND.n4698 GND.n797 19.3944
R5742 GND.n4702 GND.n797 19.3944
R5743 GND.n4702 GND.n793 19.3944
R5744 GND.n4708 GND.n793 19.3944
R5745 GND.n4708 GND.n791 19.3944
R5746 GND.n4712 GND.n791 19.3944
R5747 GND.n4712 GND.n787 19.3944
R5748 GND.n4718 GND.n787 19.3944
R5749 GND.n4718 GND.n785 19.3944
R5750 GND.n4722 GND.n785 19.3944
R5751 GND.n4722 GND.n781 19.3944
R5752 GND.n4728 GND.n781 19.3944
R5753 GND.n4728 GND.n779 19.3944
R5754 GND.n4732 GND.n779 19.3944
R5755 GND.n4732 GND.n775 19.3944
R5756 GND.n4738 GND.n775 19.3944
R5757 GND.n4738 GND.n773 19.3944
R5758 GND.n4742 GND.n773 19.3944
R5759 GND.n4742 GND.n769 19.3944
R5760 GND.n4748 GND.n769 19.3944
R5761 GND.n4748 GND.n767 19.3944
R5762 GND.n4752 GND.n767 19.3944
R5763 GND.n4752 GND.n763 19.3944
R5764 GND.n4758 GND.n763 19.3944
R5765 GND.n4758 GND.n761 19.3944
R5766 GND.n4762 GND.n761 19.3944
R5767 GND.n4762 GND.n757 19.3944
R5768 GND.n4768 GND.n757 19.3944
R5769 GND.n4768 GND.n755 19.3944
R5770 GND.n4772 GND.n755 19.3944
R5771 GND.n4772 GND.n751 19.3944
R5772 GND.n4778 GND.n751 19.3944
R5773 GND.n4778 GND.n749 19.3944
R5774 GND.n4782 GND.n749 19.3944
R5775 GND.n4782 GND.n745 19.3944
R5776 GND.n4788 GND.n745 19.3944
R5777 GND.n4788 GND.n743 19.3944
R5778 GND.n4792 GND.n743 19.3944
R5779 GND.n4792 GND.n739 19.3944
R5780 GND.n4798 GND.n739 19.3944
R5781 GND.n4798 GND.n737 19.3944
R5782 GND.n4802 GND.n737 19.3944
R5783 GND.n4802 GND.n733 19.3944
R5784 GND.n4808 GND.n733 19.3944
R5785 GND.n4808 GND.n731 19.3944
R5786 GND.n4812 GND.n731 19.3944
R5787 GND.n4812 GND.n727 19.3944
R5788 GND.n4818 GND.n727 19.3944
R5789 GND.n4818 GND.n725 19.3944
R5790 GND.n4822 GND.n725 19.3944
R5791 GND.n4822 GND.n721 19.3944
R5792 GND.n4828 GND.n721 19.3944
R5793 GND.n4828 GND.n719 19.3944
R5794 GND.n4832 GND.n719 19.3944
R5795 GND.n4832 GND.n715 19.3944
R5796 GND.n4838 GND.n715 19.3944
R5797 GND.n4838 GND.n713 19.3944
R5798 GND.n4842 GND.n713 19.3944
R5799 GND.n4842 GND.n709 19.3944
R5800 GND.n4848 GND.n709 19.3944
R5801 GND.n4848 GND.n707 19.3944
R5802 GND.n4852 GND.n707 19.3944
R5803 GND.n4852 GND.n703 19.3944
R5804 GND.n4858 GND.n703 19.3944
R5805 GND.n4858 GND.n701 19.3944
R5806 GND.n4862 GND.n701 19.3944
R5807 GND.n4862 GND.n697 19.3944
R5808 GND.n4868 GND.n697 19.3944
R5809 GND.n4868 GND.n695 19.3944
R5810 GND.n4872 GND.n695 19.3944
R5811 GND.n4872 GND.n691 19.3944
R5812 GND.n4878 GND.n691 19.3944
R5813 GND.n4878 GND.n689 19.3944
R5814 GND.n4882 GND.n689 19.3944
R5815 GND.n4882 GND.n685 19.3944
R5816 GND.n4888 GND.n685 19.3944
R5817 GND.n4888 GND.n683 19.3944
R5818 GND.n4892 GND.n683 19.3944
R5819 GND.n4892 GND.n679 19.3944
R5820 GND.n4898 GND.n679 19.3944
R5821 GND.n4898 GND.n677 19.3944
R5822 GND.n4902 GND.n677 19.3944
R5823 GND.n4902 GND.n673 19.3944
R5824 GND.n4908 GND.n673 19.3944
R5825 GND.n4908 GND.n671 19.3944
R5826 GND.n4912 GND.n671 19.3944
R5827 GND.n4912 GND.n667 19.3944
R5828 GND.n4918 GND.n667 19.3944
R5829 GND.n4918 GND.n665 19.3944
R5830 GND.n4922 GND.n665 19.3944
R5831 GND.n4922 GND.n661 19.3944
R5832 GND.n4928 GND.n661 19.3944
R5833 GND.n4928 GND.n659 19.3944
R5834 GND.n4932 GND.n659 19.3944
R5835 GND.n4932 GND.n655 19.3944
R5836 GND.n4938 GND.n655 19.3944
R5837 GND.n4938 GND.n653 19.3944
R5838 GND.n4942 GND.n653 19.3944
R5839 GND.n4942 GND.n649 19.3944
R5840 GND.n4948 GND.n649 19.3944
R5841 GND.n4948 GND.n647 19.3944
R5842 GND.n4952 GND.n647 19.3944
R5843 GND.n4952 GND.n643 19.3944
R5844 GND.n4958 GND.n643 19.3944
R5845 GND.n4958 GND.n641 19.3944
R5846 GND.n4962 GND.n641 19.3944
R5847 GND.n4962 GND.n637 19.3944
R5848 GND.n4968 GND.n637 19.3944
R5849 GND.n4968 GND.n635 19.3944
R5850 GND.n4972 GND.n635 19.3944
R5851 GND.n4972 GND.n631 19.3944
R5852 GND.n4978 GND.n631 19.3944
R5853 GND.n4978 GND.n629 19.3944
R5854 GND.n4982 GND.n629 19.3944
R5855 GND.n4982 GND.n625 19.3944
R5856 GND.n4988 GND.n625 19.3944
R5857 GND.n4988 GND.n623 19.3944
R5858 GND.n4992 GND.n623 19.3944
R5859 GND.n4992 GND.n619 19.3944
R5860 GND.n4998 GND.n619 19.3944
R5861 GND.n4998 GND.n617 19.3944
R5862 GND.n5002 GND.n617 19.3944
R5863 GND.n5002 GND.n613 19.3944
R5864 GND.n5008 GND.n613 19.3944
R5865 GND.n5008 GND.n611 19.3944
R5866 GND.n5012 GND.n611 19.3944
R5867 GND.n5012 GND.n607 19.3944
R5868 GND.n5018 GND.n607 19.3944
R5869 GND.n5018 GND.n605 19.3944
R5870 GND.n5022 GND.n605 19.3944
R5871 GND.n5022 GND.n601 19.3944
R5872 GND.n5028 GND.n601 19.3944
R5873 GND.n5028 GND.n599 19.3944
R5874 GND.n5032 GND.n599 19.3944
R5875 GND.n5032 GND.n595 19.3944
R5876 GND.n5038 GND.n595 19.3944
R5877 GND.n5038 GND.n593 19.3944
R5878 GND.n5042 GND.n593 19.3944
R5879 GND.n5042 GND.n589 19.3944
R5880 GND.n5048 GND.n589 19.3944
R5881 GND.n5048 GND.n587 19.3944
R5882 GND.n5052 GND.n587 19.3944
R5883 GND.n5052 GND.n583 19.3944
R5884 GND.n5058 GND.n583 19.3944
R5885 GND.n5058 GND.n581 19.3944
R5886 GND.n5062 GND.n581 19.3944
R5887 GND.n5062 GND.n577 19.3944
R5888 GND.n5068 GND.n577 19.3944
R5889 GND.n5068 GND.n575 19.3944
R5890 GND.n5072 GND.n575 19.3944
R5891 GND.n5072 GND.n571 19.3944
R5892 GND.n5078 GND.n571 19.3944
R5893 GND.n5078 GND.n569 19.3944
R5894 GND.n5082 GND.n569 19.3944
R5895 GND.n5082 GND.n565 19.3944
R5896 GND.n5088 GND.n565 19.3944
R5897 GND.n5088 GND.n563 19.3944
R5898 GND.n5092 GND.n563 19.3944
R5899 GND.n5092 GND.n559 19.3944
R5900 GND.n5098 GND.n559 19.3944
R5901 GND.n5098 GND.n557 19.3944
R5902 GND.n5102 GND.n557 19.3944
R5903 GND.n5102 GND.n553 19.3944
R5904 GND.n5108 GND.n553 19.3944
R5905 GND.n5108 GND.n551 19.3944
R5906 GND.n5113 GND.n551 19.3944
R5907 GND.n5113 GND.n5112 19.3944
R5908 GND.n3497 GND.n3496 19.3944
R5909 GND.n3496 GND.n3495 19.3944
R5910 GND.n3495 GND.n3494 19.3944
R5911 GND.n3494 GND.n3492 19.3944
R5912 GND.n3492 GND.n3489 19.3944
R5913 GND.n3489 GND.n3488 19.3944
R5914 GND.n3488 GND.n3485 19.3944
R5915 GND.n3485 GND.n3484 19.3944
R5916 GND.n3484 GND.n3481 19.3944
R5917 GND.n3481 GND.n3480 19.3944
R5918 GND.n3477 GND.n3476 19.3944
R5919 GND.n3476 GND.n3473 19.3944
R5920 GND.n3473 GND.n3472 19.3944
R5921 GND.n3472 GND.n3469 19.3944
R5922 GND.n3469 GND.n3468 19.3944
R5923 GND.n3468 GND.n3465 19.3944
R5924 GND.n3465 GND.n3464 19.3944
R5925 GND.n3464 GND.n3461 19.3944
R5926 GND.n3461 GND.n3460 19.3944
R5927 GND.n3460 GND.n3457 19.3944
R5928 GND.n3455 GND.n3452 19.3944
R5929 GND.n3452 GND.n3451 19.3944
R5930 GND.n3451 GND.n3448 19.3944
R5931 GND.n3448 GND.n3447 19.3944
R5932 GND.n3447 GND.n3444 19.3944
R5933 GND.n3444 GND.n3443 19.3944
R5934 GND.n3443 GND.n3440 19.3944
R5935 GND.n3440 GND.n3439 19.3944
R5936 GND.n3439 GND.n3436 19.3944
R5937 GND.n3436 GND.n3435 19.3944
R5938 GND.n3435 GND.n3432 19.3944
R5939 GND.n3430 GND.n3428 19.3944
R5940 GND.n3428 GND.n3425 19.3944
R5941 GND.n3425 GND.n3424 19.3944
R5942 GND.n3424 GND.n3421 19.3944
R5943 GND.n3421 GND.n3420 19.3944
R5944 GND.n3420 GND.n3417 19.3944
R5945 GND.n3417 GND.n3416 19.3944
R5946 GND.n3416 GND.n3413 19.3944
R5947 GND.n3413 GND.n3412 19.3944
R5948 GND.n3412 GND.n3409 19.3944
R5949 GND.n3409 GND.n3408 19.3944
R5950 GND.n3396 GND.n2145 19.3944
R5951 GND.n3396 GND.n3395 19.3944
R5952 GND.n3395 GND.n2154 19.3944
R5953 GND.n2242 GND.n2154 19.3944
R5954 GND.n3256 GND.n2242 19.3944
R5955 GND.n3257 GND.n3256 19.3944
R5956 GND.n3258 GND.n3257 19.3944
R5957 GND.n3262 GND.n3258 19.3944
R5958 GND.n3263 GND.n3262 19.3944
R5959 GND.n3264 GND.n3263 19.3944
R5960 GND.n3265 GND.n3264 19.3944
R5961 GND.n3267 GND.n3265 19.3944
R5962 GND.n3270 GND.n3267 19.3944
R5963 GND.n3271 GND.n3270 19.3944
R5964 GND.n3330 GND.n3271 19.3944
R5965 GND.n3330 GND.n3329 19.3944
R5966 GND.n3329 GND.n3328 19.3944
R5967 GND.n3328 GND.n58 19.3944
R5968 GND.n5476 GND.n58 19.3944
R5969 GND.n3399 GND.n3398 19.3944
R5970 GND.n3398 GND.n2152 19.3944
R5971 GND.n2176 GND.n2152 19.3944
R5972 GND.n3385 GND.n2176 19.3944
R5973 GND.n3385 GND.n3384 19.3944
R5974 GND.n3384 GND.n3383 19.3944
R5975 GND.n3383 GND.n2181 19.3944
R5976 GND.n2224 GND.n2181 19.3944
R5977 GND.n3366 GND.n2224 19.3944
R5978 GND.n3366 GND.n3365 19.3944
R5979 GND.n3365 GND.n3364 19.3944
R5980 GND.n3364 GND.n2228 19.3944
R5981 GND.n2228 GND.n35 19.3944
R5982 GND.n5491 GND.n35 19.3944
R5983 GND.n5491 GND.n5490 19.3944
R5984 GND.n5490 GND.n5489 19.3944
R5985 GND.n5489 GND.n39 19.3944
R5986 GND.n5479 GND.n39 19.3944
R5987 GND.n5479 GND.n5478 19.3944
R5988 GND.n177 GND.n134 19.3944
R5989 GND.n177 GND.n174 19.3944
R5990 GND.n174 GND.n173 19.3944
R5991 GND.n173 GND.n170 19.3944
R5992 GND.n170 GND.n169 19.3944
R5993 GND.n169 GND.n166 19.3944
R5994 GND.n166 GND.n165 19.3944
R5995 GND.n165 GND.n162 19.3944
R5996 GND.n162 GND.n161 19.3944
R5997 GND.n161 GND.n158 19.3944
R5998 GND.n158 GND.n157 19.3944
R5999 GND.n205 GND.n202 19.3944
R6000 GND.n202 GND.n201 19.3944
R6001 GND.n201 GND.n198 19.3944
R6002 GND.n198 GND.n197 19.3944
R6003 GND.n197 GND.n194 19.3944
R6004 GND.n194 GND.n193 19.3944
R6005 GND.n193 GND.n190 19.3944
R6006 GND.n190 GND.n189 19.3944
R6007 GND.n189 GND.n186 19.3944
R6008 GND.n186 GND.n185 19.3944
R6009 GND.n185 GND.n182 19.3944
R6010 GND.n233 GND.n232 19.3944
R6011 GND.n232 GND.n229 19.3944
R6012 GND.n229 GND.n228 19.3944
R6013 GND.n228 GND.n225 19.3944
R6014 GND.n225 GND.n224 19.3944
R6015 GND.n224 GND.n221 19.3944
R6016 GND.n221 GND.n220 19.3944
R6017 GND.n220 GND.n217 19.3944
R6018 GND.n217 GND.n216 19.3944
R6019 GND.n216 GND.n213 19.3944
R6020 GND.n213 GND.n212 19.3944
R6021 GND.n212 GND.n209 19.3944
R6022 GND.n256 GND.n255 19.3944
R6023 GND.n255 GND.n98 19.3944
R6024 GND.n251 GND.n98 19.3944
R6025 GND.n251 GND.n248 19.3944
R6026 GND.n248 GND.n245 19.3944
R6027 GND.n245 GND.n244 19.3944
R6028 GND.n244 GND.n241 19.3944
R6029 GND.n241 GND.n240 19.3944
R6030 GND.n240 GND.n237 19.3944
R6031 GND.n237 GND.n236 19.3944
R6032 GND.n3293 GND.n3290 19.3944
R6033 GND.n3293 GND.n3287 19.3944
R6034 GND.n3299 GND.n3287 19.3944
R6035 GND.n3299 GND.n3285 19.3944
R6036 GND.n3303 GND.n3285 19.3944
R6037 GND.n3303 GND.n3283 19.3944
R6038 GND.n3310 GND.n3283 19.3944
R6039 GND.n3310 GND.n3281 19.3944
R6040 GND.n3314 GND.n3281 19.3944
R6041 GND.n3315 GND.n3314 19.3944
R6042 GND.n3237 GND.n2245 19.3944
R6043 GND.n3238 GND.n3237 19.3944
R6044 GND.n3241 GND.n3238 19.3944
R6045 GND.n3241 GND.n2243 19.3944
R6046 GND.n3252 GND.n2243 19.3944
R6047 GND.n3252 GND.n3251 19.3944
R6048 GND.n3251 GND.n3250 19.3944
R6049 GND.n3250 GND.n3249 19.3944
R6050 GND.n3249 GND.n7 19.3944
R6051 GND.n5502 GND.n7 19.3944
R6052 GND.n5502 GND.n8 19.3944
R6053 GND.n2236 GND.n8 19.3944
R6054 GND.n3336 GND.n2236 19.3944
R6055 GND.n3336 GND.n3335 19.3944
R6056 GND.n3335 GND.n3334 19.3944
R6057 GND.n3334 GND.n2241 19.3944
R6058 GND.n3324 GND.n2241 19.3944
R6059 GND.n3324 GND.n3323 19.3944
R6060 GND.n3323 GND.n3322 19.3944
R6061 GND.n3205 GND.n3203 19.3944
R6062 GND.n3209 GND.n3205 19.3944
R6063 GND.n3212 GND.n3209 19.3944
R6064 GND.n3212 GND.n2253 19.3944
R6065 GND.n3217 GND.n2253 19.3944
R6066 GND.n3220 GND.n3217 19.3944
R6067 GND.n3223 GND.n3220 19.3944
R6068 GND.n3223 GND.n2251 19.3944
R6069 GND.n3227 GND.n2251 19.3944
R6070 GND.n3230 GND.n3227 19.3944
R6071 GND.n2861 GND.n2357 19.3944
R6072 GND.n2862 GND.n2861 19.3944
R6073 GND.n2865 GND.n2862 19.3944
R6074 GND.n2865 GND.n2355 19.3944
R6075 GND.n2869 GND.n2355 19.3944
R6076 GND.n2872 GND.n2869 19.3944
R6077 GND.n2873 GND.n2872 19.3944
R6078 GND.n2873 GND.n2353 19.3944
R6079 GND.n2877 GND.n2353 19.3944
R6080 GND.n2913 GND.n2877 19.3944
R6081 GND.n2914 GND.n2913 19.3944
R6082 GND.n2914 GND.n2349 19.3944
R6083 GND.n2943 GND.n2349 19.3944
R6084 GND.n2943 GND.n2942 19.3944
R6085 GND.n2942 GND.n2941 19.3944
R6086 GND.n2941 GND.n2940 19.3944
R6087 GND.n2940 GND.n2938 19.3944
R6088 GND.n2938 GND.n2937 19.3944
R6089 GND.n2937 GND.n2923 19.3944
R6090 GND.n2933 GND.n2923 19.3944
R6091 GND.n2933 GND.n2932 19.3944
R6092 GND.n2932 GND.n2931 19.3944
R6093 GND.n2931 GND.n2930 19.3944
R6094 GND.n2930 GND.n2315 19.3944
R6095 GND.n3051 GND.n2315 19.3944
R6096 GND.n3051 GND.n2313 19.3944
R6097 GND.n3060 GND.n2313 19.3944
R6098 GND.n3060 GND.n3059 19.3944
R6099 GND.n3059 GND.n3058 19.3944
R6100 GND.n3058 GND.n2297 19.3944
R6101 GND.n3074 GND.n2297 19.3944
R6102 GND.n3074 GND.n2295 19.3944
R6103 GND.n3081 GND.n2295 19.3944
R6104 GND.n3081 GND.n3080 19.3944
R6105 GND.n3080 GND.n2280 19.3944
R6106 GND.n2280 GND.n2278 19.3944
R6107 GND.n3104 GND.n2278 19.3944
R6108 GND.n3104 GND.n2276 19.3944
R6109 GND.n3109 GND.n2276 19.3944
R6110 GND.n3109 GND.n2266 19.3944
R6111 GND.n3144 GND.n2266 19.3944
R6112 GND.n3145 GND.n3144 19.3944
R6113 GND.n3145 GND.n2264 19.3944
R6114 GND.n3149 GND.n2264 19.3944
R6115 GND.n3149 GND.n2262 19.3944
R6116 GND.n3153 GND.n2262 19.3944
R6117 GND.n3153 GND.n2260 19.3944
R6118 GND.n3158 GND.n2260 19.3944
R6119 GND.n3158 GND.n2257 19.3944
R6120 GND.n3185 GND.n2257 19.3944
R6121 GND.n3186 GND.n3185 19.3944
R6122 GND.n3189 GND.n3186 19.3944
R6123 GND.n3189 GND.n2255 19.3944
R6124 GND.n3193 GND.n2255 19.3944
R6125 GND.n3198 GND.n3193 19.3944
R6126 GND.n3199 GND.n3198 19.3944
R6127 GND.n3199 GND.n1938 19.3944
R6128 GND.n3517 GND.n3516 19.3944
R6129 GND.n3516 GND.n3513 19.3944
R6130 GND.n3513 GND.n3512 19.3944
R6131 GND.n3547 GND.n1905 19.3944
R6132 GND.n3542 GND.n1905 19.3944
R6133 GND.n3542 GND.n3541 19.3944
R6134 GND.n3541 GND.n3540 19.3944
R6135 GND.n3540 GND.n3537 19.3944
R6136 GND.n3537 GND.n3536 19.3944
R6137 GND.n3536 GND.n3533 19.3944
R6138 GND.n3533 GND.n3532 19.3944
R6139 GND.n3532 GND.n3529 19.3944
R6140 GND.n3529 GND.n3528 19.3944
R6141 GND.n3528 GND.n3525 19.3944
R6142 GND.n3525 GND.n3524 19.3944
R6143 GND.n3524 GND.n3521 19.3944
R6144 GND.n3521 GND.n3520 19.3944
R6145 GND.n3809 GND.n3808 19.3944
R6146 GND.n3808 GND.n3807 19.3944
R6147 GND.n3807 GND.n1558 19.3944
R6148 GND.n1577 GND.n1558 19.3944
R6149 GND.n3795 GND.n1577 19.3944
R6150 GND.n3795 GND.n3794 19.3944
R6151 GND.n3794 GND.n3793 19.3944
R6152 GND.n3793 GND.n1583 19.3944
R6153 GND.n3710 GND.n1583 19.3944
R6154 GND.n3710 GND.n3709 19.3944
R6155 GND.n3709 GND.n3708 19.3944
R6156 GND.n3708 GND.n1649 19.3944
R6157 GND.n2948 GND.n1649 19.3944
R6158 GND.n2948 GND.n1676 19.3944
R6159 GND.n3689 GND.n1676 19.3944
R6160 GND.n3689 GND.n3688 19.3944
R6161 GND.n3688 GND.n3687 19.3944
R6162 GND.n3687 GND.n1680 19.3944
R6163 GND.n2325 GND.n1680 19.3944
R6164 GND.n2329 GND.n2325 19.3944
R6165 GND.n2329 GND.n2323 19.3944
R6166 GND.n3037 GND.n2323 19.3944
R6167 GND.n3037 GND.n2321 19.3944
R6168 GND.n3046 GND.n2321 19.3944
R6169 GND.n3046 GND.n3045 19.3944
R6170 GND.n3045 GND.n3044 19.3944
R6171 GND.n3044 GND.n2309 19.3944
R6172 GND.n2309 GND.n2307 19.3944
R6173 GND.n3066 GND.n2307 19.3944
R6174 GND.n3066 GND.n2305 19.3944
R6175 GND.n3070 GND.n2305 19.3944
R6176 GND.n3070 GND.n2290 19.3944
R6177 GND.n3085 GND.n2290 19.3944
R6178 GND.n3085 GND.n2288 19.3944
R6179 GND.n3098 GND.n2288 19.3944
R6180 GND.n3098 GND.n3097 19.3944
R6181 GND.n3097 GND.n3096 19.3944
R6182 GND.n3096 GND.n3093 19.3944
R6183 GND.n3093 GND.n1791 19.3944
R6184 GND.n3605 GND.n1791 19.3944
R6185 GND.n3605 GND.n3604 19.3944
R6186 GND.n3604 GND.n3603 19.3944
R6187 GND.n3603 GND.n1795 19.3944
R6188 GND.n3168 GND.n1795 19.3944
R6189 GND.n3168 GND.n3165 19.3944
R6190 GND.n3172 GND.n3165 19.3944
R6191 GND.n3172 GND.n3163 19.3944
R6192 GND.n3179 GND.n3163 19.3944
R6193 GND.n3179 GND.n3178 19.3944
R6194 GND.n3178 GND.n1877 19.3944
R6195 GND.n3565 GND.n1877 19.3944
R6196 GND.n3565 GND.n3564 19.3944
R6197 GND.n3564 GND.n3563 19.3944
R6198 GND.n3563 GND.n1881 19.3944
R6199 GND.n1900 GND.n1881 19.3944
R6200 GND.n3551 GND.n1900 19.3944
R6201 GND.n3551 GND.n3550 19.3944
R6202 GND.n3861 GND.n3860 19.3944
R6203 GND.n3860 GND.n1531 19.3944
R6204 GND.n3853 GND.n1531 19.3944
R6205 GND.n3847 GND.n3846 19.3944
R6206 GND.n3846 GND.n3845 19.3944
R6207 GND.n3845 GND.n3844 19.3944
R6208 GND.n3844 GND.n3842 19.3944
R6209 GND.n3842 GND.n3839 19.3944
R6210 GND.n3839 GND.n3838 19.3944
R6211 GND.n3838 GND.n3835 19.3944
R6212 GND.n3835 GND.n3834 19.3944
R6213 GND.n3834 GND.n3831 19.3944
R6214 GND.n3831 GND.n3830 19.3944
R6215 GND.n3830 GND.n3827 19.3944
R6216 GND.n3827 GND.n3826 19.3944
R6217 GND.n3826 GND.n1527 19.3944
R6218 GND.n3865 GND.n1527 19.3944
R6219 GND.n2163 GND.n2162 19.3944
R6220 GND.n3391 GND.n2162 19.3944
R6221 GND.n3391 GND.n3390 19.3944
R6222 GND.n3390 GND.n3389 19.3944
R6223 GND.n3389 GND.n2168 19.3944
R6224 GND.n3379 GND.n23 19.3944
R6225 GND.n2187 GND.n23 19.3944
R6226 GND.n5498 GND.n16 19.3944
R6227 GND.n2231 GND.n17 19.3944
R6228 GND.n5495 GND.n25 19.3944
R6229 GND.n5495 GND.n26 19.3944
R6230 GND.n5485 GND.n26 19.3944
R6231 GND.n5485 GND.n5484 19.3944
R6232 GND.n5484 GND.n5483 19.3944
R6233 GND.n5483 GND.n49 19.3944
R6234 GND.n4200 GND.n4199 19.3944
R6235 GND.n4199 GND.n4198 19.3944
R6236 GND.n4198 GND.n1146 19.3944
R6237 GND.n4192 GND.n1146 19.3944
R6238 GND.n4192 GND.n4191 19.3944
R6239 GND.n4191 GND.n4190 19.3944
R6240 GND.n4190 GND.n1154 19.3944
R6241 GND.n4184 GND.n1154 19.3944
R6242 GND.n4184 GND.n4183 19.3944
R6243 GND.n4183 GND.n4182 19.3944
R6244 GND.n4182 GND.n1162 19.3944
R6245 GND.n4176 GND.n1162 19.3944
R6246 GND.n4176 GND.n4175 19.3944
R6247 GND.n4175 GND.n4174 19.3944
R6248 GND.n4174 GND.n1170 19.3944
R6249 GND.n4168 GND.n1170 19.3944
R6250 GND.n4168 GND.n4167 19.3944
R6251 GND.n4167 GND.n4166 19.3944
R6252 GND.n4166 GND.n1178 19.3944
R6253 GND.n4160 GND.n1178 19.3944
R6254 GND.n4160 GND.n4159 19.3944
R6255 GND.n4159 GND.n4158 19.3944
R6256 GND.n4158 GND.n1186 19.3944
R6257 GND.n4152 GND.n1186 19.3944
R6258 GND.n4152 GND.n4151 19.3944
R6259 GND.n4151 GND.n4150 19.3944
R6260 GND.n4150 GND.n1194 19.3944
R6261 GND.n4144 GND.n1194 19.3944
R6262 GND.n4144 GND.n4143 19.3944
R6263 GND.n4143 GND.n4142 19.3944
R6264 GND.n4142 GND.n1202 19.3944
R6265 GND.n4136 GND.n1202 19.3944
R6266 GND.n4136 GND.n4135 19.3944
R6267 GND.n4135 GND.n4134 19.3944
R6268 GND.n4134 GND.n1210 19.3944
R6269 GND.n4128 GND.n1210 19.3944
R6270 GND.n4128 GND.n4127 19.3944
R6271 GND.n4127 GND.n4126 19.3944
R6272 GND.n4126 GND.n1218 19.3944
R6273 GND.n4120 GND.n1218 19.3944
R6274 GND.n4120 GND.n4119 19.3944
R6275 GND.n4119 GND.n4118 19.3944
R6276 GND.n4118 GND.n1226 19.3944
R6277 GND.n4112 GND.n1226 19.3944
R6278 GND.n4112 GND.n4111 19.3944
R6279 GND.n4111 GND.n4110 19.3944
R6280 GND.n4110 GND.n1234 19.3944
R6281 GND.n4104 GND.n1234 19.3944
R6282 GND.n4104 GND.n4103 19.3944
R6283 GND.n4103 GND.n4102 19.3944
R6284 GND.n4102 GND.n1242 19.3944
R6285 GND.n4096 GND.n1242 19.3944
R6286 GND.n4096 GND.n4095 19.3944
R6287 GND.n4095 GND.n4094 19.3944
R6288 GND.n4094 GND.n1250 19.3944
R6289 GND.n4088 GND.n1250 19.3944
R6290 GND.n4088 GND.n4087 19.3944
R6291 GND.n4087 GND.n4086 19.3944
R6292 GND.n4086 GND.n1258 19.3944
R6293 GND.n4080 GND.n1258 19.3944
R6294 GND.n4080 GND.n4079 19.3944
R6295 GND.n4079 GND.n4078 19.3944
R6296 GND.n4078 GND.n1266 19.3944
R6297 GND.n4072 GND.n1266 19.3944
R6298 GND.n4072 GND.n4071 19.3944
R6299 GND.n4071 GND.n4070 19.3944
R6300 GND.n4070 GND.n1274 19.3944
R6301 GND.n4064 GND.n1274 19.3944
R6302 GND.n4064 GND.n4063 19.3944
R6303 GND.n4063 GND.n4062 19.3944
R6304 GND.n4062 GND.n1282 19.3944
R6305 GND.n4056 GND.n1282 19.3944
R6306 GND.n4056 GND.n4055 19.3944
R6307 GND.n4055 GND.n4054 19.3944
R6308 GND.n4054 GND.n1290 19.3944
R6309 GND.n4048 GND.n1290 19.3944
R6310 GND.n4048 GND.n4047 19.3944
R6311 GND.n4047 GND.n4046 19.3944
R6312 GND.n4046 GND.n1298 19.3944
R6313 GND.n4040 GND.n1298 19.3944
R6314 GND.n4040 GND.n4039 19.3944
R6315 GND.n4039 GND.n4038 19.3944
R6316 GND.n4038 GND.n1306 19.3944
R6317 GND.n4032 GND.n1306 19.3944
R6318 GND.n4032 GND.n4031 19.3944
R6319 GND.n4031 GND.n4030 19.3944
R6320 GND.n4030 GND.n1314 19.3944
R6321 GND.n4024 GND.n1314 19.3944
R6322 GND.n4024 GND.n4023 19.3944
R6323 GND.n4023 GND.n4022 19.3944
R6324 GND.n4022 GND.n1322 19.3944
R6325 GND.n4016 GND.n1322 19.3944
R6326 GND.n4016 GND.n4015 19.3944
R6327 GND.n4015 GND.n4014 19.3944
R6328 GND.n4014 GND.n1330 19.3944
R6329 GND.n4008 GND.n1330 19.3944
R6330 GND.n4008 GND.n4007 19.3944
R6331 GND.n4007 GND.n4006 19.3944
R6332 GND.n4006 GND.n1338 19.3944
R6333 GND.n4000 GND.n1338 19.3944
R6334 GND.n4000 GND.n3999 19.3944
R6335 GND.n3999 GND.n3998 19.3944
R6336 GND.n3998 GND.n1346 19.3944
R6337 GND.n3992 GND.n1346 19.3944
R6338 GND.n3992 GND.n3991 19.3944
R6339 GND.n3991 GND.n3990 19.3944
R6340 GND.n3990 GND.n1354 19.3944
R6341 GND.n2440 GND.n1354 19.3944
R6342 GND.n2515 GND.n2440 19.3944
R6343 GND.n2515 GND.n2514 19.3944
R6344 GND.n2514 GND.n2513 19.3944
R6345 GND.n2509 GND.n2446 19.3944
R6346 GND.n2505 GND.n2451 19.3944
R6347 GND.n2503 GND.n2502 19.3944
R6348 GND.n2499 GND.n2498 19.3944
R6349 GND.n2495 GND.n2494 19.3944
R6350 GND.n2494 GND.n2493 19.3944
R6351 GND.n2493 GND.n2455 19.3944
R6352 GND.n2489 GND.n2455 19.3944
R6353 GND.n2489 GND.n2488 19.3944
R6354 GND.n2488 GND.n2487 19.3944
R6355 GND.n2487 GND.n2461 19.3944
R6356 GND.n2481 GND.n2461 19.3944
R6357 GND.n2481 GND.n2480 19.3944
R6358 GND.n2480 GND.n2479 19.3944
R6359 GND.n2479 GND.n2467 19.3944
R6360 GND.n2471 GND.n2467 19.3944
R6361 GND.n2471 GND.n1565 19.3944
R6362 GND.n3802 GND.n1565 19.3944
R6363 GND.n3802 GND.n3801 19.3944
R6364 GND.n3801 GND.n3800 19.3944
R6365 GND.n3800 GND.n1569 19.3944
R6366 GND.n2882 GND.n1569 19.3944
R6367 GND.n2885 GND.n2882 19.3944
R6368 GND.n2885 GND.n2879 19.3944
R6369 GND.n2890 GND.n2879 19.3944
R6370 GND.n2890 GND.n1657 19.3944
R6371 GND.n3703 GND.n1657 19.3944
R6372 GND.n3703 GND.n3702 19.3944
R6373 GND.n3702 GND.n3701 19.3944
R6374 GND.n3701 GND.n1661 19.3944
R6375 GND.n1690 GND.n1661 19.3944
R6376 GND.n1690 GND.n1687 19.3944
R6377 GND.n3682 GND.n1687 19.3944
R6378 GND.n3682 GND.n3681 19.3944
R6379 GND.n3681 GND.n3680 19.3944
R6380 GND.n3680 GND.n1696 19.3944
R6381 GND.n3668 GND.n1696 19.3944
R6382 GND.n3668 GND.n3667 19.3944
R6383 GND.n3667 GND.n3666 19.3944
R6384 GND.n3666 GND.n1714 19.3944
R6385 GND.n3654 GND.n1714 19.3944
R6386 GND.n3654 GND.n3653 19.3944
R6387 GND.n3653 GND.n3652 19.3944
R6388 GND.n3652 GND.n1731 19.3944
R6389 GND.n3640 GND.n1731 19.3944
R6390 GND.n3640 GND.n3639 19.3944
R6391 GND.n3639 GND.n3638 19.3944
R6392 GND.n3638 GND.n1749 19.3944
R6393 GND.n3626 GND.n1749 19.3944
R6394 GND.n3626 GND.n3625 19.3944
R6395 GND.n3625 GND.n3624 19.3944
R6396 GND.n3624 GND.n1766 19.3944
R6397 GND.n3612 GND.n1766 19.3944
R6398 GND.n3612 GND.n3611 19.3944
R6399 GND.n3611 GND.n3610 19.3944
R6400 GND.n3610 GND.n1784 19.3944
R6401 GND.n1812 GND.n1784 19.3944
R6402 GND.n1812 GND.n1809 19.3944
R6403 GND.n3591 GND.n1809 19.3944
R6404 GND.n3591 GND.n3590 19.3944
R6405 GND.n3590 GND.n3589 19.3944
R6406 GND.n3589 GND.n1818 19.3944
R6407 GND.n1864 GND.n1818 19.3944
R6408 GND.n3572 GND.n1864 19.3944
R6409 GND.n3572 GND.n3571 19.3944
R6410 GND.n3571 GND.n3570 19.3944
R6411 GND.n3570 GND.n1870 19.3944
R6412 GND.n1887 GND.n1870 19.3944
R6413 GND.n3558 GND.n1887 19.3944
R6414 GND.n3558 GND.n3557 19.3944
R6415 GND.n3557 GND.n3556 19.3944
R6416 GND.n3556 GND.n1893 19.3944
R6417 GND.n3506 GND.n1893 19.3944
R6418 GND.n3506 GND.n3505 19.3944
R6419 GND.n3505 GND.n3504 19.3944
R6420 GND.n3504 GND.n1944 19.3944
R6421 GND.n2199 GND.n1944 19.3944
R6422 GND.n2203 GND.n2199 19.3944
R6423 GND.n2203 GND.n2198 19.3944
R6424 GND.n2207 GND.n2198 19.3944
R6425 GND.n2207 GND.n2196 19.3944
R6426 GND.n2212 GND.n2196 19.3944
R6427 GND.n2212 GND.n2194 19.3944
R6428 GND.n2216 GND.n2194 19.3944
R6429 GND.n3374 GND.n2218 19.3944
R6430 GND.n3372 GND.n3371 19.3944
R6431 GND.n3359 GND.n3341 19.3944
R6432 GND.n3357 GND.n3356 19.3944
R6433 GND.n3353 GND.n3352 19.3944
R6434 GND.n3352 GND.n3351 19.3944
R6435 GND.n3351 GND.n3348 19.3944
R6436 GND.n3348 GND.n64 19.3944
R6437 GND.n5471 GND.n64 19.3944
R6438 GND.n5471 GND.n5470 19.3944
R6439 GND.n5470 GND.n5469 19.3944
R6440 GND.n5469 GND.n68 19.3944
R6441 GND.n5463 GND.n68 19.3944
R6442 GND.n5463 GND.n5462 19.3944
R6443 GND.n5462 GND.n5461 19.3944
R6444 GND.n5461 GND.n265 19.3944
R6445 GND.n5455 GND.n265 19.3944
R6446 GND.n5455 GND.n5454 19.3944
R6447 GND.n5454 GND.n5453 19.3944
R6448 GND.n5453 GND.n273 19.3944
R6449 GND.n5447 GND.n273 19.3944
R6450 GND.n5447 GND.n5446 19.3944
R6451 GND.n5446 GND.n5445 19.3944
R6452 GND.n5445 GND.n281 19.3944
R6453 GND.n5439 GND.n281 19.3944
R6454 GND.n5439 GND.n5438 19.3944
R6455 GND.n5438 GND.n5437 19.3944
R6456 GND.n5437 GND.n289 19.3944
R6457 GND.n5431 GND.n289 19.3944
R6458 GND.n5431 GND.n5430 19.3944
R6459 GND.n5430 GND.n5429 19.3944
R6460 GND.n5429 GND.n297 19.3944
R6461 GND.n5423 GND.n297 19.3944
R6462 GND.n5423 GND.n5422 19.3944
R6463 GND.n5422 GND.n5421 19.3944
R6464 GND.n5421 GND.n305 19.3944
R6465 GND.n5415 GND.n305 19.3944
R6466 GND.n5415 GND.n5414 19.3944
R6467 GND.n5414 GND.n5413 19.3944
R6468 GND.n5413 GND.n313 19.3944
R6469 GND.n5407 GND.n313 19.3944
R6470 GND.n5407 GND.n5406 19.3944
R6471 GND.n5406 GND.n5405 19.3944
R6472 GND.n5405 GND.n321 19.3944
R6473 GND.n5399 GND.n321 19.3944
R6474 GND.n5399 GND.n5398 19.3944
R6475 GND.n5398 GND.n5397 19.3944
R6476 GND.n5397 GND.n329 19.3944
R6477 GND.n5391 GND.n329 19.3944
R6478 GND.n5391 GND.n5390 19.3944
R6479 GND.n5390 GND.n5389 19.3944
R6480 GND.n5389 GND.n337 19.3944
R6481 GND.n5383 GND.n337 19.3944
R6482 GND.n5383 GND.n5382 19.3944
R6483 GND.n5382 GND.n5381 19.3944
R6484 GND.n5381 GND.n345 19.3944
R6485 GND.n5375 GND.n345 19.3944
R6486 GND.n5375 GND.n5374 19.3944
R6487 GND.n5374 GND.n5373 19.3944
R6488 GND.n5373 GND.n353 19.3944
R6489 GND.n5367 GND.n353 19.3944
R6490 GND.n5367 GND.n5366 19.3944
R6491 GND.n5366 GND.n5365 19.3944
R6492 GND.n5365 GND.n361 19.3944
R6493 GND.n5359 GND.n361 19.3944
R6494 GND.n5359 GND.n5358 19.3944
R6495 GND.n5358 GND.n5357 19.3944
R6496 GND.n5357 GND.n369 19.3944
R6497 GND.n5351 GND.n369 19.3944
R6498 GND.n5351 GND.n5350 19.3944
R6499 GND.n5350 GND.n5349 19.3944
R6500 GND.n5349 GND.n377 19.3944
R6501 GND.n5343 GND.n377 19.3944
R6502 GND.n5343 GND.n5342 19.3944
R6503 GND.n5342 GND.n5341 19.3944
R6504 GND.n5341 GND.n385 19.3944
R6505 GND.n5335 GND.n385 19.3944
R6506 GND.n5335 GND.n5334 19.3944
R6507 GND.n5334 GND.n5333 19.3944
R6508 GND.n5333 GND.n393 19.3944
R6509 GND.n5327 GND.n393 19.3944
R6510 GND.n5327 GND.n5326 19.3944
R6511 GND.n5326 GND.n5325 19.3944
R6512 GND.n5325 GND.n401 19.3944
R6513 GND.n5319 GND.n401 19.3944
R6514 GND.n5319 GND.n5318 19.3944
R6515 GND.n5318 GND.n5317 19.3944
R6516 GND.n5317 GND.n409 19.3944
R6517 GND.n5311 GND.n409 19.3944
R6518 GND.n5311 GND.n5310 19.3944
R6519 GND.n5310 GND.n5309 19.3944
R6520 GND.n5309 GND.n417 19.3944
R6521 GND.n5303 GND.n417 19.3944
R6522 GND.n5303 GND.n5302 19.3944
R6523 GND.n5302 GND.n5301 19.3944
R6524 GND.n5301 GND.n425 19.3944
R6525 GND.n5295 GND.n425 19.3944
R6526 GND.n5295 GND.n5294 19.3944
R6527 GND.n5294 GND.n5293 19.3944
R6528 GND.n5293 GND.n433 19.3944
R6529 GND.n5287 GND.n433 19.3944
R6530 GND.n5287 GND.n5286 19.3944
R6531 GND.n5286 GND.n5285 19.3944
R6532 GND.n5285 GND.n441 19.3944
R6533 GND.n5279 GND.n441 19.3944
R6534 GND.n5279 GND.n5278 19.3944
R6535 GND.n5278 GND.n5277 19.3944
R6536 GND.n5277 GND.n449 19.3944
R6537 GND.n5271 GND.n449 19.3944
R6538 GND.n5271 GND.n5270 19.3944
R6539 GND.n5270 GND.n5269 19.3944
R6540 GND.n5269 GND.n457 19.3944
R6541 GND.n5263 GND.n457 19.3944
R6542 GND.n5263 GND.n5262 19.3944
R6543 GND.n5262 GND.n5261 19.3944
R6544 GND.n2596 GND.n2595 19.3944
R6545 GND.n2601 GND.n2596 19.3944
R6546 GND.n2601 GND.n2592 19.3944
R6547 GND.n2605 GND.n2592 19.3944
R6548 GND.n2605 GND.n2590 19.3944
R6549 GND.n2611 GND.n2590 19.3944
R6550 GND.n2611 GND.n2588 19.3944
R6551 GND.n2615 GND.n2588 19.3944
R6552 GND.n2615 GND.n2583 19.3944
R6553 GND.n2621 GND.n2583 19.3944
R6554 GND.n2625 GND.n2581 19.3944
R6555 GND.n2625 GND.n2579 19.3944
R6556 GND.n2631 GND.n2579 19.3944
R6557 GND.n2631 GND.n2577 19.3944
R6558 GND.n2635 GND.n2577 19.3944
R6559 GND.n2635 GND.n2575 19.3944
R6560 GND.n2641 GND.n2575 19.3944
R6561 GND.n2641 GND.n2573 19.3944
R6562 GND.n2646 GND.n2573 19.3944
R6563 GND.n2646 GND.n2571 19.3944
R6564 GND.n2652 GND.n2571 19.3944
R6565 GND.n2653 GND.n2652 19.3944
R6566 GND.n2656 GND.n2565 19.3944
R6567 GND.n2662 GND.n2565 19.3944
R6568 GND.n2662 GND.n2563 19.3944
R6569 GND.n2666 GND.n2563 19.3944
R6570 GND.n2666 GND.n2561 19.3944
R6571 GND.n2672 GND.n2561 19.3944
R6572 GND.n2672 GND.n2559 19.3944
R6573 GND.n2676 GND.n2559 19.3944
R6574 GND.n2676 GND.n2557 19.3944
R6575 GND.n2682 GND.n2557 19.3944
R6576 GND.n2682 GND.n2555 19.3944
R6577 GND.n2694 GND.n2553 19.3944
R6578 GND.n2694 GND.n2551 19.3944
R6579 GND.n2698 GND.n2551 19.3944
R6580 GND.n2698 GND.n2549 19.3944
R6581 GND.n2704 GND.n2549 19.3944
R6582 GND.n2704 GND.n2547 19.3944
R6583 GND.n2708 GND.n2547 19.3944
R6584 GND.n2708 GND.n2545 19.3944
R6585 GND.n2714 GND.n2545 19.3944
R6586 GND.n2714 GND.n2543 19.3944
R6587 GND.n2718 GND.n2543 19.3944
R6588 GND.n3985 GND.n3984 19.3944
R6589 GND.n3984 GND.n3983 19.3944
R6590 GND.n3983 GND.n1366 19.3944
R6591 GND.n2431 GND.n1366 19.3944
R6592 GND.n2778 GND.n2431 19.3944
R6593 GND.n2783 GND.n2780 19.3944
R6594 GND.n2783 GND.n2782 19.3944
R6595 GND.n2803 GND.n2408 19.3944
R6596 GND.n2808 GND.n2805 19.3944
R6597 GND.n2806 GND.n2388 19.3944
R6598 GND.n2830 GND.n2388 19.3944
R6599 GND.n2830 GND.n2386 19.3944
R6600 GND.n2834 GND.n2386 19.3944
R6601 GND.n2834 GND.n1418 19.3944
R6602 GND.n3948 GND.n1418 19.3944
R6603 GND.n4312 GND.n4311 19.3944
R6604 GND.n4311 GND.n4310 19.3944
R6605 GND.n4310 GND.n1034 19.3944
R6606 GND.n4304 GND.n1034 19.3944
R6607 GND.n4304 GND.n4303 19.3944
R6608 GND.n4303 GND.n4302 19.3944
R6609 GND.n4302 GND.n1042 19.3944
R6610 GND.n4296 GND.n1042 19.3944
R6611 GND.n4296 GND.n4295 19.3944
R6612 GND.n4295 GND.n4294 19.3944
R6613 GND.n4294 GND.n1050 19.3944
R6614 GND.n4288 GND.n1050 19.3944
R6615 GND.n4288 GND.n4287 19.3944
R6616 GND.n4287 GND.n4286 19.3944
R6617 GND.n4286 GND.n1058 19.3944
R6618 GND.n4280 GND.n1058 19.3944
R6619 GND.n4280 GND.n4279 19.3944
R6620 GND.n4279 GND.n4278 19.3944
R6621 GND.n4278 GND.n1066 19.3944
R6622 GND.n4272 GND.n1066 19.3944
R6623 GND.n4272 GND.n4271 19.3944
R6624 GND.n4271 GND.n4270 19.3944
R6625 GND.n4270 GND.n1074 19.3944
R6626 GND.n4264 GND.n1074 19.3944
R6627 GND.n4264 GND.n4263 19.3944
R6628 GND.n4263 GND.n4262 19.3944
R6629 GND.n4262 GND.n1082 19.3944
R6630 GND.n4256 GND.n1082 19.3944
R6631 GND.n4256 GND.n4255 19.3944
R6632 GND.n4255 GND.n4254 19.3944
R6633 GND.n4254 GND.n1090 19.3944
R6634 GND.n4248 GND.n1090 19.3944
R6635 GND.n4248 GND.n4247 19.3944
R6636 GND.n4247 GND.n4246 19.3944
R6637 GND.n4246 GND.n1098 19.3944
R6638 GND.n4240 GND.n1098 19.3944
R6639 GND.n4240 GND.n4239 19.3944
R6640 GND.n4239 GND.n4238 19.3944
R6641 GND.n4238 GND.n1106 19.3944
R6642 GND.n4232 GND.n1106 19.3944
R6643 GND.n4232 GND.n4231 19.3944
R6644 GND.n4231 GND.n4230 19.3944
R6645 GND.n4230 GND.n1114 19.3944
R6646 GND.n4224 GND.n1114 19.3944
R6647 GND.n4224 GND.n4223 19.3944
R6648 GND.n4223 GND.n4222 19.3944
R6649 GND.n4222 GND.n1122 19.3944
R6650 GND.n4216 GND.n1122 19.3944
R6651 GND.n4216 GND.n4215 19.3944
R6652 GND.n4215 GND.n4214 19.3944
R6653 GND.n4214 GND.n1130 19.3944
R6654 GND.n4208 GND.n1130 19.3944
R6655 GND.n4208 GND.n4207 19.3944
R6656 GND.n4207 GND.n4206 19.3944
R6657 GND.n4206 GND.n1138 19.3944
R6658 GND.n2731 GND.n2537 19.3944
R6659 GND.n2731 GND.n2535 19.3944
R6660 GND.n2737 GND.n2535 19.3944
R6661 GND.n2737 GND.n2533 19.3944
R6662 GND.n2741 GND.n2533 19.3944
R6663 GND.n2741 GND.n2531 19.3944
R6664 GND.n2747 GND.n2531 19.3944
R6665 GND.n2747 GND.n2529 19.3944
R6666 GND.n2751 GND.n2529 19.3944
R6667 GND.n2751 GND.n2527 19.3944
R6668 GND.n2763 GND.n2759 19.3944
R6669 GND.n2764 GND.n2763 19.3944
R6670 GND.n2764 GND.n2520 19.3944
R6671 GND.n2769 GND.n2520 19.3944
R6672 GND.n2769 GND.n2521 19.3944
R6673 GND.n2521 GND.n2420 19.3944
R6674 GND.n2787 GND.n2420 19.3944
R6675 GND.n2787 GND.n2417 19.3944
R6676 GND.n2793 GND.n2417 19.3944
R6677 GND.n2793 GND.n2418 19.3944
R6678 GND.n2418 GND.n2399 19.3944
R6679 GND.n2812 GND.n2399 19.3944
R6680 GND.n2812 GND.n2396 19.3944
R6681 GND.n2822 GND.n2396 19.3944
R6682 GND.n2822 GND.n2397 19.3944
R6683 GND.n2818 GND.n2397 19.3944
R6684 GND.n2818 GND.n2379 19.3944
R6685 GND.n2841 GND.n2379 19.3944
R6686 GND.n2842 GND.n2841 19.3944
R6687 GND.n3914 GND.n1452 18.6187
R6688 GND.n3457 GND.n3456 18.6187
R6689 GND.n2795 GND.t130 18.343
R6690 GND.n2476 GND.n2475 18.343
R6691 GND.n2475 GND.n2474 18.343
R6692 GND.n2474 GND.n2473 18.343
R6693 GND.n2473 GND.n1560 18.343
R6694 GND.n3805 GND.n1560 18.343
R6695 GND.n3805 GND.n3804 18.343
R6696 GND.n3804 GND.n1562 18.343
R6697 GND.n1572 GND.n1571 18.343
R6698 GND.n3798 GND.n1572 18.343
R6699 GND.n3798 GND.n3797 18.343
R6700 GND.n3797 GND.n1574 18.343
R6701 GND.n2870 GND.n1574 18.343
R6702 GND.n2870 GND.n1585 18.343
R6703 GND.n3791 GND.n1585 18.343
R6704 GND.n2351 GND.n1605 18.343
R6705 GND.t70 GND.n2892 18.343
R6706 GND.n3706 GND.n3705 18.343
R6707 GND.n3691 GND.n1673 18.343
R6708 GND.n3685 GND.n3684 18.343
R6709 GND.n3678 GND.n1698 18.343
R6710 GND.n2979 GND.n1706 18.343
R6711 GND.n3031 GND.n3030 18.343
R6712 GND.n3062 GND.n2310 18.343
R6713 GND.n3010 GND.n1735 18.343
R6714 GND.n3010 GND.n1741 18.343
R6715 GND.n2303 GND.n2302 18.343
R6716 GND.n2285 GND.n2284 18.343
R6717 GND.n2990 GND.n1770 18.343
R6718 GND.n3614 GND.n1778 18.343
R6719 GND.n3608 GND.n3607 18.343
R6720 GND.n3601 GND.t104 18.343
R6721 GND.n3593 GND.n1806 18.343
R6722 GND.n3587 GND.n1820 18.343
R6723 GND.n3587 GND.n1822 18.343
R6724 GND.n3159 GND.n1829 18.343
R6725 GND.n3574 GND.n1861 18.343
R6726 GND.n2009 GND.n1861 18.343
R6727 GND.n3568 GND.n1872 18.343
R6728 GND.n3568 GND.n3567 18.343
R6729 GND.n3567 GND.n1874 18.343
R6730 GND.n3187 GND.n1874 18.343
R6731 GND.n3187 GND.n1883 18.343
R6732 GND.n3561 GND.n1883 18.343
R6733 GND.n3561 GND.n3560 18.343
R6734 GND.n3195 GND.n3194 18.343
R6735 GND.n3194 GND.n1895 18.343
R6736 GND.n3554 GND.n1895 18.343
R6737 GND.n3554 GND.n3553 18.343
R6738 GND.n3553 GND.n1897 18.343
R6739 GND.n3509 GND.n1897 18.343
R6740 GND.n3509 GND.n3508 18.343
R6741 GND.n5500 GND.t1 18.343
R6742 GND.n1632 GND.n1631 18.2581
R6743 GND.n1856 GND.n1855 18.2581
R6744 GND.n1621 GND.n1620 17.9571
R6745 GND.n1853 GND.n1852 17.9571
R6746 GND.t16 GND.n2383 17.6093
R6747 GND.n2975 GND.n2974 17.6093
R6748 GND.n3671 GND.n3670 17.6093
R6749 GND.n3622 GND.n3621 17.6093
R6750 GND.n2274 GND.n2273 17.6093
R6751 GND.t32 GND.n2158 17.6093
R6752 GND.n3891 GND.n3890 17.2611
R6753 GND.n3432 GND.n3431 17.2611
R6754 GND.n182 GND.n181 17.2611
R6755 GND.n2688 GND.n2555 17.2611
R6756 GND.n3712 GND.n1643 16.8756
R6757 GND.n3698 GND.n1664 16.8756
R6758 GND.n3019 GND.n3016 16.8756
R6759 GND.n3072 GND.n2301 16.8756
R6760 GND.n3181 GND.n3160 16.8756
R6761 GND.n3664 GND.n1716 16.1419
R6762 GND.n3628 GND.n1760 16.1419
R6763 GND.n2267 GND.n1788 16.1419
R6764 GND.n2816 GND.t16 15.4082
R6765 GND.n2341 GND.n2340 15.4082
R6766 GND.n3048 GND.n2318 15.4082
R6767 GND.n2317 GND.t4 15.4082
R6768 GND.n2292 GND.t5 15.4082
R6769 GND.n3083 GND.n2293 15.4082
R6770 GND.n3142 GND.n3141 15.4082
R6771 GND.n3239 GND.t32 15.4082
R6772 GND.n3872 GND.n3871 14.9338
R6773 GND.n3408 GND.n2141 14.9338
R6774 GND.n157 GND.n154 14.9338
R6775 GND.n2718 GND.n2541 14.9338
R6776 GND.t130 GND.n2410 14.6745
R6777 GND.n3692 GND.n1670 14.6745
R6778 GND.n3657 GND.n3656 14.6745
R6779 GND.n3636 GND.n3635 14.6745
R6780 GND.n3600 GND.n1799 14.6745
R6781 GND.n3369 GND.t1 14.6745
R6782 GND.n3787 GND.n1634 14.6737
R6783 GND.n2066 GND.n1858 14.6737
R6784 GND.n3035 GND.n3034 13.9408
R6785 GND.n3100 GND.n2283 13.9408
R6786 GND.n1839 GND.n1838 13.5524
R6787 GND.n2911 GND.n2898 13.2071
R6788 GND.n2951 GND.n2346 13.2071
R6789 GND.n3650 GND.n1733 13.2071
R6790 GND.n3642 GND.n1743 13.2071
R6791 GND.n3130 GND.n3129 13.2071
R6792 GND.n3581 GND.n1828 13.2071
R6793 GND.n1633 GND.n1609 13.1884
R6794 GND.n1628 GND.n1627 13.1884
R6795 GND.n1627 GND.n1626 13.1884
R6796 GND.n1626 GND.n1612 13.1884
R6797 GND.n1622 GND.n1612 13.1884
R6798 GND.n1841 GND.n1840 13.1884
R6799 GND.n1841 GND.n1836 13.1884
R6800 GND.n1845 GND.n1836 13.1884
R6801 GND.n1846 GND.n1845 13.1884
R6802 GND.n3791 GND.n3790 12.8403
R6803 GND.n2351 GND.t9 12.4734
R6804 GND.n2903 GND.t122 12.4734
R6805 GND.n3677 GND.n1700 12.4734
R6806 GND.n2980 GND.n1700 12.4734
R6807 GND.n2991 GND.n1776 12.4734
R6808 GND.n3615 GND.n1776 12.4734
R6809 GND.n2517 GND.t12 11.7397
R6810 GND.n2904 GND.n2346 11.7397
R6811 GND.n2950 GND.t49 11.7397
R6812 GND.n3650 GND.n3649 11.7397
R6813 GND.n3643 GND.n3642 11.7397
R6814 GND.n3129 GND.t85 11.7397
R6815 GND.t52 GND.n44 11.7397
R6816 GND.n1857 GND.n1834 11.6369
R6817 GND.n3871 GND.n3870 11.055
R6818 GND.n3404 GND.n2141 11.055
R6819 GND.n154 GND.n149 11.055
R6820 GND.n2723 GND.n2541 11.055
R6821 GND.t23 GND.n1682 11.006
R6822 GND.n2973 GND.n2337 11.006
R6823 GND.n3035 GND.n1708 11.006
R6824 GND.n3100 GND.n1768 11.006
R6825 GND.n3120 GND.n3111 11.006
R6826 GND.n3594 GND.t43 11.006
R6827 GND.n2022 GND.n2005 10.6151
R6828 GND.n2025 GND.n2022 10.6151
R6829 GND.n2026 GND.n2025 10.6151
R6830 GND.n2030 GND.n2029 10.6151
R6831 GND.n2033 GND.n2030 10.6151
R6832 GND.n2034 GND.n2033 10.6151
R6833 GND.n2037 GND.n2034 10.6151
R6834 GND.n2038 GND.n2037 10.6151
R6835 GND.n2041 GND.n2038 10.6151
R6836 GND.n2042 GND.n2041 10.6151
R6837 GND.n2045 GND.n2042 10.6151
R6838 GND.n2046 GND.n2045 10.6151
R6839 GND.n2049 GND.n2046 10.6151
R6840 GND.n2051 GND.n2049 10.6151
R6841 GND.n2052 GND.n2051 10.6151
R6842 GND.n2054 GND.n2052 10.6151
R6843 GND.n3715 GND.n1639 10.6151
R6844 GND.n2896 GND.n1639 10.6151
R6845 GND.n2896 GND.n2895 10.6151
R6846 GND.n2895 GND.n2894 10.6151
R6847 GND.n2894 GND.n2344 10.6151
R6848 GND.n2953 GND.n2344 10.6151
R6849 GND.n2954 GND.n2953 10.6151
R6850 GND.n2957 GND.n2954 10.6151
R6851 GND.n2958 GND.n2957 10.6151
R6852 GND.n2959 GND.n2958 10.6151
R6853 GND.n2963 GND.n2959 10.6151
R6854 GND.n2963 GND.n2962 10.6151
R6855 GND.n2962 GND.n2961 10.6151
R6856 GND.n2961 GND.n2335 10.6151
R6857 GND.n2977 GND.n2335 10.6151
R6858 GND.n2978 GND.n2977 10.6151
R6859 GND.n2982 GND.n2978 10.6151
R6860 GND.n2983 GND.n2982 10.6151
R6861 GND.n2984 GND.n2983 10.6151
R6862 GND.n3028 GND.n2984 10.6151
R6863 GND.n3028 GND.n3027 10.6151
R6864 GND.n3027 GND.n3026 10.6151
R6865 GND.n3026 GND.n3025 10.6151
R6866 GND.n3025 GND.n3023 10.6151
R6867 GND.n3023 GND.n3022 10.6151
R6868 GND.n3022 GND.n2985 10.6151
R6869 GND.n3014 GND.n2985 10.6151
R6870 GND.n3014 GND.n3013 10.6151
R6871 GND.n3013 GND.n3012 10.6151
R6872 GND.n3012 GND.n3009 10.6151
R6873 GND.n3009 GND.n3008 10.6151
R6874 GND.n3008 GND.n2986 10.6151
R6875 GND.n3004 GND.n2986 10.6151
R6876 GND.n3004 GND.n3003 10.6151
R6877 GND.n3003 GND.n3002 10.6151
R6878 GND.n3002 GND.n3000 10.6151
R6879 GND.n3000 GND.n2999 10.6151
R6880 GND.n2999 GND.n2987 10.6151
R6881 GND.n2995 GND.n2987 10.6151
R6882 GND.n2995 GND.n2994 10.6151
R6883 GND.n2994 GND.n2993 10.6151
R6884 GND.n2993 GND.n2989 10.6151
R6885 GND.n2989 GND.n2988 10.6151
R6886 GND.n2988 GND.n2272 10.6151
R6887 GND.n2272 GND.n2270 10.6151
R6888 GND.n3124 GND.n2270 10.6151
R6889 GND.n3125 GND.n3124 10.6151
R6890 GND.n3139 GND.n3125 10.6151
R6891 GND.n3139 GND.n3138 10.6151
R6892 GND.n3138 GND.n3137 10.6151
R6893 GND.n3137 GND.n3133 10.6151
R6894 GND.n3133 GND.n3132 10.6151
R6895 GND.n3132 GND.n1825 10.6151
R6896 GND.n3585 GND.n1825 10.6151
R6897 GND.n3585 GND.n3584 10.6151
R6898 GND.n3584 GND.n3583 10.6151
R6899 GND.n3583 GND.n1826 10.6151
R6900 GND.n2053 GND.n1826 10.6151
R6901 GND.n3751 GND.n3748 10.6151
R6902 GND.n3748 GND.n3747 10.6151
R6903 GND.n3747 GND.n3744 10.6151
R6904 GND.n3742 GND.n3739 10.6151
R6905 GND.n3739 GND.n3738 10.6151
R6906 GND.n3738 GND.n3735 10.6151
R6907 GND.n3735 GND.n3734 10.6151
R6908 GND.n3734 GND.n3731 10.6151
R6909 GND.n3731 GND.n3730 10.6151
R6910 GND.n3730 GND.n3727 10.6151
R6911 GND.n3727 GND.n3726 10.6151
R6912 GND.n3726 GND.n3723 10.6151
R6913 GND.n3723 GND.n3722 10.6151
R6914 GND.n3722 GND.n3719 10.6151
R6915 GND.n3719 GND.n3718 10.6151
R6916 GND.n3718 GND.n3716 10.6151
R6917 GND.n3787 GND.n3786 10.6151
R6918 GND.n3786 GND.n3785 10.6151
R6919 GND.n3785 GND.n3784 10.6151
R6920 GND.n3784 GND.n3782 10.6151
R6921 GND.n3782 GND.n3779 10.6151
R6922 GND.n3779 GND.n3778 10.6151
R6923 GND.n3778 GND.n3775 10.6151
R6924 GND.n3775 GND.n3774 10.6151
R6925 GND.n3774 GND.n3771 10.6151
R6926 GND.n3771 GND.n3770 10.6151
R6927 GND.n3770 GND.n3767 10.6151
R6928 GND.n3767 GND.n3766 10.6151
R6929 GND.n3766 GND.n3763 10.6151
R6930 GND.n3761 GND.n3758 10.6151
R6931 GND.n3758 GND.n3757 10.6151
R6932 GND.n3757 GND.n3754 10.6151
R6933 GND.n2067 GND.n2066 10.6151
R6934 GND.n2099 GND.n2067 10.6151
R6935 GND.n2099 GND.n2098 10.6151
R6936 GND.n2098 GND.n2097 10.6151
R6937 GND.n2097 GND.n2094 10.6151
R6938 GND.n2094 GND.n2093 10.6151
R6939 GND.n2093 GND.n2090 10.6151
R6940 GND.n2090 GND.n2089 10.6151
R6941 GND.n2089 GND.n2086 10.6151
R6942 GND.n2086 GND.n2085 10.6151
R6943 GND.n2085 GND.n2082 10.6151
R6944 GND.n2082 GND.n2081 10.6151
R6945 GND.n2081 GND.n2078 10.6151
R6946 GND.n2076 GND.n2073 10.6151
R6947 GND.n2073 GND.n2072 10.6151
R6948 GND.n2072 GND.n2006 10.6151
R6949 GND.n2902 GND.n2901 10.6151
R6950 GND.n2909 GND.n2902 10.6151
R6951 GND.n2909 GND.n2908 10.6151
R6952 GND.n2908 GND.n2907 10.6151
R6953 GND.n2907 GND.n2906 10.6151
R6954 GND.n2906 GND.n1667 10.6151
R6955 GND.n3696 GND.n1667 10.6151
R6956 GND.n3696 GND.n3695 10.6151
R6957 GND.n3695 GND.n3694 10.6151
R6958 GND.n3694 GND.n1668 10.6151
R6959 GND.n2339 GND.n1668 10.6151
R6960 GND.n2969 GND.n2339 10.6151
R6961 GND.n2970 GND.n2969 10.6151
R6962 GND.n2971 GND.n2970 10.6151
R6963 GND.n2971 GND.n1703 10.6151
R6964 GND.n3675 GND.n1703 10.6151
R6965 GND.n3675 GND.n3674 10.6151
R6966 GND.n3674 GND.n3673 10.6151
R6967 GND.n3673 GND.n1704 10.6151
R6968 GND.n3032 GND.n1704 10.6151
R6969 GND.n3032 GND.n1720 10.6151
R6970 GND.n3661 GND.n1720 10.6151
R6971 GND.n3661 GND.n3660 10.6151
R6972 GND.n3660 GND.n3659 10.6151
R6973 GND.n3659 GND.n1721 10.6151
R6974 GND.n3017 GND.n1721 10.6151
R6975 GND.n3017 GND.n1738 10.6151
R6976 GND.n3647 GND.n1738 10.6151
R6977 GND.n3647 GND.n3646 10.6151
R6978 GND.n3646 GND.n3645 10.6151
R6979 GND.n3645 GND.n1739 10.6151
R6980 GND.n2299 GND.n1739 10.6151
R6981 GND.n2299 GND.n1756 10.6151
R6982 GND.n3633 GND.n1756 10.6151
R6983 GND.n3633 GND.n3632 10.6151
R6984 GND.n3632 GND.n3631 10.6151
R6985 GND.n3631 GND.n1757 10.6151
R6986 GND.n2281 GND.n1757 10.6151
R6987 GND.n2281 GND.n1773 10.6151
R6988 GND.n3619 GND.n1773 10.6151
R6989 GND.n3619 GND.n3618 10.6151
R6990 GND.n3618 GND.n3617 10.6151
R6991 GND.n3617 GND.n1774 10.6151
R6992 GND.n3118 GND.n1774 10.6151
R6993 GND.n3118 GND.n3117 10.6151
R6994 GND.n3117 GND.n3116 10.6151
R6995 GND.n3116 GND.n3113 10.6151
R6996 GND.n3113 GND.n1802 10.6151
R6997 GND.n3598 GND.n1802 10.6151
R6998 GND.n3598 GND.n3597 10.6151
R6999 GND.n3597 GND.n3596 10.6151
R7000 GND.n3596 GND.n1803 10.6151
R7001 GND.n3127 GND.n1803 10.6151
R7002 GND.n3127 GND.n3126 10.6151
R7003 GND.n3126 GND.n1833 10.6151
R7004 GND.n3579 GND.n1833 10.6151
R7005 GND.n3579 GND.n3578 10.6151
R7006 GND.n3578 GND.n3577 10.6151
R7007 GND.n1571 GND.t39 10.2723
R7008 GND.n3713 GND.n1641 10.2723
R7009 GND.n3656 GND.n1725 10.2723
R7010 GND.n3636 GND.n1751 10.2723
R7011 GND.n3575 GND.n3574 10.2723
R7012 GND.n3560 GND.t88 10.2723
R7013 GND.n2966 GND.n2340 9.5386
R7014 GND.n3142 GND.n2268 9.5386
R7015 GND.n2029 GND.n2021 9.36635
R7016 GND.n3743 GND.n3742 9.36635
R7017 GND.n3763 GND.n3762 9.36635
R7018 GND.n2078 GND.n2077 9.36635
R7019 GND.n1027 GND.n1026 9.3005
R7020 GND.n4319 GND.n4318 9.3005
R7021 GND.n4320 GND.n1025 9.3005
R7022 GND.n4322 GND.n4321 9.3005
R7023 GND.n1021 GND.n1020 9.3005
R7024 GND.n4329 GND.n4328 9.3005
R7025 GND.n4330 GND.n1019 9.3005
R7026 GND.n4332 GND.n4331 9.3005
R7027 GND.n1015 GND.n1014 9.3005
R7028 GND.n4339 GND.n4338 9.3005
R7029 GND.n4340 GND.n1013 9.3005
R7030 GND.n4342 GND.n4341 9.3005
R7031 GND.n1009 GND.n1008 9.3005
R7032 GND.n4349 GND.n4348 9.3005
R7033 GND.n4350 GND.n1007 9.3005
R7034 GND.n4352 GND.n4351 9.3005
R7035 GND.n1003 GND.n1002 9.3005
R7036 GND.n4359 GND.n4358 9.3005
R7037 GND.n4360 GND.n1001 9.3005
R7038 GND.n4362 GND.n4361 9.3005
R7039 GND.n997 GND.n996 9.3005
R7040 GND.n4369 GND.n4368 9.3005
R7041 GND.n4370 GND.n995 9.3005
R7042 GND.n4372 GND.n4371 9.3005
R7043 GND.n991 GND.n990 9.3005
R7044 GND.n4379 GND.n4378 9.3005
R7045 GND.n4380 GND.n989 9.3005
R7046 GND.n4382 GND.n4381 9.3005
R7047 GND.n985 GND.n984 9.3005
R7048 GND.n4389 GND.n4388 9.3005
R7049 GND.n4390 GND.n983 9.3005
R7050 GND.n4392 GND.n4391 9.3005
R7051 GND.n979 GND.n978 9.3005
R7052 GND.n4399 GND.n4398 9.3005
R7053 GND.n4400 GND.n977 9.3005
R7054 GND.n4402 GND.n4401 9.3005
R7055 GND.n973 GND.n972 9.3005
R7056 GND.n4409 GND.n4408 9.3005
R7057 GND.n4410 GND.n971 9.3005
R7058 GND.n4412 GND.n4411 9.3005
R7059 GND.n967 GND.n966 9.3005
R7060 GND.n4419 GND.n4418 9.3005
R7061 GND.n4420 GND.n965 9.3005
R7062 GND.n4422 GND.n4421 9.3005
R7063 GND.n961 GND.n960 9.3005
R7064 GND.n4429 GND.n4428 9.3005
R7065 GND.n4430 GND.n959 9.3005
R7066 GND.n4432 GND.n4431 9.3005
R7067 GND.n955 GND.n954 9.3005
R7068 GND.n4439 GND.n4438 9.3005
R7069 GND.n4440 GND.n953 9.3005
R7070 GND.n4442 GND.n4441 9.3005
R7071 GND.n949 GND.n948 9.3005
R7072 GND.n4449 GND.n4448 9.3005
R7073 GND.n4450 GND.n947 9.3005
R7074 GND.n4452 GND.n4451 9.3005
R7075 GND.n943 GND.n942 9.3005
R7076 GND.n4459 GND.n4458 9.3005
R7077 GND.n4460 GND.n941 9.3005
R7078 GND.n4462 GND.n4461 9.3005
R7079 GND.n937 GND.n936 9.3005
R7080 GND.n4469 GND.n4468 9.3005
R7081 GND.n4470 GND.n935 9.3005
R7082 GND.n4472 GND.n4471 9.3005
R7083 GND.n931 GND.n930 9.3005
R7084 GND.n4479 GND.n4478 9.3005
R7085 GND.n4480 GND.n929 9.3005
R7086 GND.n4482 GND.n4481 9.3005
R7087 GND.n925 GND.n924 9.3005
R7088 GND.n4489 GND.n4488 9.3005
R7089 GND.n4490 GND.n923 9.3005
R7090 GND.n4492 GND.n4491 9.3005
R7091 GND.n919 GND.n918 9.3005
R7092 GND.n4499 GND.n4498 9.3005
R7093 GND.n4500 GND.n917 9.3005
R7094 GND.n4502 GND.n4501 9.3005
R7095 GND.n913 GND.n912 9.3005
R7096 GND.n4509 GND.n4508 9.3005
R7097 GND.n4510 GND.n911 9.3005
R7098 GND.n4512 GND.n4511 9.3005
R7099 GND.n907 GND.n906 9.3005
R7100 GND.n4519 GND.n4518 9.3005
R7101 GND.n4520 GND.n905 9.3005
R7102 GND.n4522 GND.n4521 9.3005
R7103 GND.n901 GND.n900 9.3005
R7104 GND.n4529 GND.n4528 9.3005
R7105 GND.n4530 GND.n899 9.3005
R7106 GND.n4532 GND.n4531 9.3005
R7107 GND.n895 GND.n894 9.3005
R7108 GND.n4539 GND.n4538 9.3005
R7109 GND.n4540 GND.n893 9.3005
R7110 GND.n4542 GND.n4541 9.3005
R7111 GND.n889 GND.n888 9.3005
R7112 GND.n4549 GND.n4548 9.3005
R7113 GND.n4550 GND.n887 9.3005
R7114 GND.n4552 GND.n4551 9.3005
R7115 GND.n883 GND.n882 9.3005
R7116 GND.n4559 GND.n4558 9.3005
R7117 GND.n4560 GND.n881 9.3005
R7118 GND.n4562 GND.n4561 9.3005
R7119 GND.n877 GND.n876 9.3005
R7120 GND.n4569 GND.n4568 9.3005
R7121 GND.n4570 GND.n875 9.3005
R7122 GND.n4572 GND.n4571 9.3005
R7123 GND.n871 GND.n870 9.3005
R7124 GND.n4579 GND.n4578 9.3005
R7125 GND.n4580 GND.n869 9.3005
R7126 GND.n4582 GND.n4581 9.3005
R7127 GND.n865 GND.n864 9.3005
R7128 GND.n4589 GND.n4588 9.3005
R7129 GND.n4590 GND.n863 9.3005
R7130 GND.n4592 GND.n4591 9.3005
R7131 GND.n859 GND.n858 9.3005
R7132 GND.n4599 GND.n4598 9.3005
R7133 GND.n4600 GND.n857 9.3005
R7134 GND.n4602 GND.n4601 9.3005
R7135 GND.n853 GND.n852 9.3005
R7136 GND.n4609 GND.n4608 9.3005
R7137 GND.n4610 GND.n851 9.3005
R7138 GND.n4612 GND.n4611 9.3005
R7139 GND.n847 GND.n846 9.3005
R7140 GND.n4619 GND.n4618 9.3005
R7141 GND.n4620 GND.n845 9.3005
R7142 GND.n4622 GND.n4621 9.3005
R7143 GND.n841 GND.n840 9.3005
R7144 GND.n4629 GND.n4628 9.3005
R7145 GND.n4630 GND.n839 9.3005
R7146 GND.n4632 GND.n4631 9.3005
R7147 GND.n835 GND.n834 9.3005
R7148 GND.n4639 GND.n4638 9.3005
R7149 GND.n4640 GND.n833 9.3005
R7150 GND.n4642 GND.n4641 9.3005
R7151 GND.n829 GND.n828 9.3005
R7152 GND.n4649 GND.n4648 9.3005
R7153 GND.n4650 GND.n827 9.3005
R7154 GND.n4652 GND.n4651 9.3005
R7155 GND.n823 GND.n822 9.3005
R7156 GND.n4659 GND.n4658 9.3005
R7157 GND.n4660 GND.n821 9.3005
R7158 GND.n4662 GND.n4661 9.3005
R7159 GND.n817 GND.n816 9.3005
R7160 GND.n4669 GND.n4668 9.3005
R7161 GND.n4670 GND.n815 9.3005
R7162 GND.n4672 GND.n4671 9.3005
R7163 GND.n811 GND.n810 9.3005
R7164 GND.n4679 GND.n4678 9.3005
R7165 GND.n4680 GND.n809 9.3005
R7166 GND.n4682 GND.n4681 9.3005
R7167 GND.n805 GND.n804 9.3005
R7168 GND.n4689 GND.n4688 9.3005
R7169 GND.n4690 GND.n803 9.3005
R7170 GND.n4692 GND.n4691 9.3005
R7171 GND.n799 GND.n798 9.3005
R7172 GND.n4699 GND.n4698 9.3005
R7173 GND.n4700 GND.n797 9.3005
R7174 GND.n4702 GND.n4701 9.3005
R7175 GND.n793 GND.n792 9.3005
R7176 GND.n4709 GND.n4708 9.3005
R7177 GND.n4710 GND.n791 9.3005
R7178 GND.n4712 GND.n4711 9.3005
R7179 GND.n787 GND.n786 9.3005
R7180 GND.n4719 GND.n4718 9.3005
R7181 GND.n4720 GND.n785 9.3005
R7182 GND.n4722 GND.n4721 9.3005
R7183 GND.n781 GND.n780 9.3005
R7184 GND.n4729 GND.n4728 9.3005
R7185 GND.n4730 GND.n779 9.3005
R7186 GND.n4732 GND.n4731 9.3005
R7187 GND.n775 GND.n774 9.3005
R7188 GND.n4739 GND.n4738 9.3005
R7189 GND.n4740 GND.n773 9.3005
R7190 GND.n4742 GND.n4741 9.3005
R7191 GND.n769 GND.n768 9.3005
R7192 GND.n4749 GND.n4748 9.3005
R7193 GND.n4750 GND.n767 9.3005
R7194 GND.n4752 GND.n4751 9.3005
R7195 GND.n763 GND.n762 9.3005
R7196 GND.n4759 GND.n4758 9.3005
R7197 GND.n4760 GND.n761 9.3005
R7198 GND.n4762 GND.n4761 9.3005
R7199 GND.n757 GND.n756 9.3005
R7200 GND.n4769 GND.n4768 9.3005
R7201 GND.n4770 GND.n755 9.3005
R7202 GND.n4772 GND.n4771 9.3005
R7203 GND.n751 GND.n750 9.3005
R7204 GND.n4779 GND.n4778 9.3005
R7205 GND.n4780 GND.n749 9.3005
R7206 GND.n4782 GND.n4781 9.3005
R7207 GND.n745 GND.n744 9.3005
R7208 GND.n4789 GND.n4788 9.3005
R7209 GND.n4790 GND.n743 9.3005
R7210 GND.n4792 GND.n4791 9.3005
R7211 GND.n739 GND.n738 9.3005
R7212 GND.n4799 GND.n4798 9.3005
R7213 GND.n4800 GND.n737 9.3005
R7214 GND.n4802 GND.n4801 9.3005
R7215 GND.n733 GND.n732 9.3005
R7216 GND.n4809 GND.n4808 9.3005
R7217 GND.n4810 GND.n731 9.3005
R7218 GND.n4812 GND.n4811 9.3005
R7219 GND.n727 GND.n726 9.3005
R7220 GND.n4819 GND.n4818 9.3005
R7221 GND.n4820 GND.n725 9.3005
R7222 GND.n4822 GND.n4821 9.3005
R7223 GND.n721 GND.n720 9.3005
R7224 GND.n4829 GND.n4828 9.3005
R7225 GND.n4830 GND.n719 9.3005
R7226 GND.n4832 GND.n4831 9.3005
R7227 GND.n715 GND.n714 9.3005
R7228 GND.n4839 GND.n4838 9.3005
R7229 GND.n4840 GND.n713 9.3005
R7230 GND.n4842 GND.n4841 9.3005
R7231 GND.n709 GND.n708 9.3005
R7232 GND.n4849 GND.n4848 9.3005
R7233 GND.n4850 GND.n707 9.3005
R7234 GND.n4852 GND.n4851 9.3005
R7235 GND.n703 GND.n702 9.3005
R7236 GND.n4859 GND.n4858 9.3005
R7237 GND.n4860 GND.n701 9.3005
R7238 GND.n4862 GND.n4861 9.3005
R7239 GND.n697 GND.n696 9.3005
R7240 GND.n4869 GND.n4868 9.3005
R7241 GND.n4870 GND.n695 9.3005
R7242 GND.n4872 GND.n4871 9.3005
R7243 GND.n691 GND.n690 9.3005
R7244 GND.n4879 GND.n4878 9.3005
R7245 GND.n4880 GND.n689 9.3005
R7246 GND.n4882 GND.n4881 9.3005
R7247 GND.n685 GND.n684 9.3005
R7248 GND.n4889 GND.n4888 9.3005
R7249 GND.n4890 GND.n683 9.3005
R7250 GND.n4892 GND.n4891 9.3005
R7251 GND.n679 GND.n678 9.3005
R7252 GND.n4899 GND.n4898 9.3005
R7253 GND.n4900 GND.n677 9.3005
R7254 GND.n4902 GND.n4901 9.3005
R7255 GND.n673 GND.n672 9.3005
R7256 GND.n4909 GND.n4908 9.3005
R7257 GND.n4910 GND.n671 9.3005
R7258 GND.n4912 GND.n4911 9.3005
R7259 GND.n667 GND.n666 9.3005
R7260 GND.n4919 GND.n4918 9.3005
R7261 GND.n4920 GND.n665 9.3005
R7262 GND.n4922 GND.n4921 9.3005
R7263 GND.n661 GND.n660 9.3005
R7264 GND.n4929 GND.n4928 9.3005
R7265 GND.n4930 GND.n659 9.3005
R7266 GND.n4932 GND.n4931 9.3005
R7267 GND.n655 GND.n654 9.3005
R7268 GND.n4939 GND.n4938 9.3005
R7269 GND.n4940 GND.n653 9.3005
R7270 GND.n4942 GND.n4941 9.3005
R7271 GND.n649 GND.n648 9.3005
R7272 GND.n4949 GND.n4948 9.3005
R7273 GND.n4950 GND.n647 9.3005
R7274 GND.n4952 GND.n4951 9.3005
R7275 GND.n643 GND.n642 9.3005
R7276 GND.n4959 GND.n4958 9.3005
R7277 GND.n4960 GND.n641 9.3005
R7278 GND.n4962 GND.n4961 9.3005
R7279 GND.n637 GND.n636 9.3005
R7280 GND.n4969 GND.n4968 9.3005
R7281 GND.n4970 GND.n635 9.3005
R7282 GND.n4972 GND.n4971 9.3005
R7283 GND.n631 GND.n630 9.3005
R7284 GND.n4979 GND.n4978 9.3005
R7285 GND.n4980 GND.n629 9.3005
R7286 GND.n4982 GND.n4981 9.3005
R7287 GND.n625 GND.n624 9.3005
R7288 GND.n4989 GND.n4988 9.3005
R7289 GND.n4990 GND.n623 9.3005
R7290 GND.n4992 GND.n4991 9.3005
R7291 GND.n619 GND.n618 9.3005
R7292 GND.n4999 GND.n4998 9.3005
R7293 GND.n5000 GND.n617 9.3005
R7294 GND.n5002 GND.n5001 9.3005
R7295 GND.n613 GND.n612 9.3005
R7296 GND.n5009 GND.n5008 9.3005
R7297 GND.n5010 GND.n611 9.3005
R7298 GND.n5012 GND.n5011 9.3005
R7299 GND.n607 GND.n606 9.3005
R7300 GND.n5019 GND.n5018 9.3005
R7301 GND.n5020 GND.n605 9.3005
R7302 GND.n5022 GND.n5021 9.3005
R7303 GND.n601 GND.n600 9.3005
R7304 GND.n5029 GND.n5028 9.3005
R7305 GND.n5030 GND.n599 9.3005
R7306 GND.n5032 GND.n5031 9.3005
R7307 GND.n595 GND.n594 9.3005
R7308 GND.n5039 GND.n5038 9.3005
R7309 GND.n5040 GND.n593 9.3005
R7310 GND.n5042 GND.n5041 9.3005
R7311 GND.n589 GND.n588 9.3005
R7312 GND.n5049 GND.n5048 9.3005
R7313 GND.n5050 GND.n587 9.3005
R7314 GND.n5052 GND.n5051 9.3005
R7315 GND.n583 GND.n582 9.3005
R7316 GND.n5059 GND.n5058 9.3005
R7317 GND.n5060 GND.n581 9.3005
R7318 GND.n5062 GND.n5061 9.3005
R7319 GND.n577 GND.n576 9.3005
R7320 GND.n5069 GND.n5068 9.3005
R7321 GND.n5070 GND.n575 9.3005
R7322 GND.n5072 GND.n5071 9.3005
R7323 GND.n571 GND.n570 9.3005
R7324 GND.n5079 GND.n5078 9.3005
R7325 GND.n5080 GND.n569 9.3005
R7326 GND.n5082 GND.n5081 9.3005
R7327 GND.n565 GND.n564 9.3005
R7328 GND.n5089 GND.n5088 9.3005
R7329 GND.n5090 GND.n563 9.3005
R7330 GND.n5092 GND.n5091 9.3005
R7331 GND.n559 GND.n558 9.3005
R7332 GND.n5099 GND.n5098 9.3005
R7333 GND.n5100 GND.n557 9.3005
R7334 GND.n5102 GND.n5101 9.3005
R7335 GND.n553 GND.n552 9.3005
R7336 GND.n5109 GND.n5108 9.3005
R7337 GND.n5110 GND.n551 9.3005
R7338 GND.n5113 GND.n5111 9.3005
R7339 GND.n5112 GND.n547 9.3005
R7340 GND.n5121 GND.n546 9.3005
R7341 GND.n5123 GND.n5122 9.3005
R7342 GND.n542 GND.n541 9.3005
R7343 GND.n5130 GND.n5129 9.3005
R7344 GND.n5131 GND.n540 9.3005
R7345 GND.n5133 GND.n5132 9.3005
R7346 GND.n536 GND.n535 9.3005
R7347 GND.n5140 GND.n5139 9.3005
R7348 GND.n5141 GND.n534 9.3005
R7349 GND.n5143 GND.n5142 9.3005
R7350 GND.n530 GND.n529 9.3005
R7351 GND.n5150 GND.n5149 9.3005
R7352 GND.n5151 GND.n528 9.3005
R7353 GND.n5153 GND.n5152 9.3005
R7354 GND.n524 GND.n523 9.3005
R7355 GND.n5160 GND.n5159 9.3005
R7356 GND.n5161 GND.n522 9.3005
R7357 GND.n5163 GND.n5162 9.3005
R7358 GND.n518 GND.n517 9.3005
R7359 GND.n5170 GND.n5169 9.3005
R7360 GND.n5171 GND.n516 9.3005
R7361 GND.n5173 GND.n5172 9.3005
R7362 GND.n512 GND.n511 9.3005
R7363 GND.n5180 GND.n5179 9.3005
R7364 GND.n5181 GND.n510 9.3005
R7365 GND.n5183 GND.n5182 9.3005
R7366 GND.n506 GND.n505 9.3005
R7367 GND.n5190 GND.n5189 9.3005
R7368 GND.n5191 GND.n504 9.3005
R7369 GND.n5193 GND.n5192 9.3005
R7370 GND.n500 GND.n499 9.3005
R7371 GND.n5200 GND.n5199 9.3005
R7372 GND.n5201 GND.n498 9.3005
R7373 GND.n5203 GND.n5202 9.3005
R7374 GND.n494 GND.n493 9.3005
R7375 GND.n5210 GND.n5209 9.3005
R7376 GND.n5211 GND.n492 9.3005
R7377 GND.n5213 GND.n5212 9.3005
R7378 GND.n488 GND.n487 9.3005
R7379 GND.n5220 GND.n5219 9.3005
R7380 GND.n5221 GND.n486 9.3005
R7381 GND.n5223 GND.n5222 9.3005
R7382 GND.n482 GND.n481 9.3005
R7383 GND.n5230 GND.n5229 9.3005
R7384 GND.n5231 GND.n480 9.3005
R7385 GND.n5233 GND.n5232 9.3005
R7386 GND.n476 GND.n475 9.3005
R7387 GND.n5240 GND.n5239 9.3005
R7388 GND.n5241 GND.n474 9.3005
R7389 GND.n5243 GND.n5242 9.3005
R7390 GND.n470 GND.n469 9.3005
R7391 GND.n5250 GND.n5249 9.3005
R7392 GND.n5251 GND.n468 9.3005
R7393 GND.n5255 GND.n5252 9.3005
R7394 GND.n5254 GND.n5253 9.3005
R7395 GND.n5120 GND.n5119 9.3005
R7396 GND.n2861 GND.n2860 9.3005
R7397 GND.n2862 GND.n2356 9.3005
R7398 GND.n2866 GND.n2865 9.3005
R7399 GND.n2867 GND.n2355 9.3005
R7400 GND.n2869 GND.n2868 9.3005
R7401 GND.n2872 GND.n2354 9.3005
R7402 GND.n2874 GND.n2873 9.3005
R7403 GND.n2875 GND.n2353 9.3005
R7404 GND.n2877 GND.n2876 9.3005
R7405 GND.n2913 GND.n2350 9.3005
R7406 GND.n2915 GND.n2914 9.3005
R7407 GND.n2916 GND.n2349 9.3005
R7408 GND.n2943 GND.n2917 9.3005
R7409 GND.n2942 GND.n2918 9.3005
R7410 GND.n2941 GND.n2919 9.3005
R7411 GND.n2940 GND.n2920 9.3005
R7412 GND.n2938 GND.n2921 9.3005
R7413 GND.n2937 GND.n2922 9.3005
R7414 GND.n2925 GND.n2923 9.3005
R7415 GND.n2933 GND.n2926 9.3005
R7416 GND.n2932 GND.n2927 9.3005
R7417 GND.n2931 GND.n2928 9.3005
R7418 GND.n2930 GND.n2929 9.3005
R7419 GND.n2315 GND.n2314 9.3005
R7420 GND.n3052 GND.n3051 9.3005
R7421 GND.n3053 GND.n2313 9.3005
R7422 GND.n3060 GND.n3054 9.3005
R7423 GND.n3059 GND.n3055 9.3005
R7424 GND.n3058 GND.n3056 9.3005
R7425 GND.n2297 GND.n2296 9.3005
R7426 GND.n3075 GND.n3074 9.3005
R7427 GND.n3076 GND.n2295 9.3005
R7428 GND.n3081 GND.n3077 9.3005
R7429 GND.n3080 GND.n3079 9.3005
R7430 GND.n3078 GND.n2280 9.3005
R7431 GND.n2278 GND.n2277 9.3005
R7432 GND.n3105 GND.n3104 9.3005
R7433 GND.n3106 GND.n2276 9.3005
R7434 GND.n3109 GND.n3108 9.3005
R7435 GND.n3107 GND.n2266 9.3005
R7436 GND.n3144 GND.n2265 9.3005
R7437 GND.n3146 GND.n3145 9.3005
R7438 GND.n3147 GND.n2264 9.3005
R7439 GND.n3149 GND.n3148 9.3005
R7440 GND.n2262 GND.n2261 9.3005
R7441 GND.n3154 GND.n3153 9.3005
R7442 GND.n3155 GND.n2260 9.3005
R7443 GND.n3158 GND.n3157 9.3005
R7444 GND.n3156 GND.n2257 9.3005
R7445 GND.n3185 GND.n2258 9.3005
R7446 GND.n3186 GND.n2256 9.3005
R7447 GND.n3190 GND.n3189 9.3005
R7448 GND.n3191 GND.n2255 9.3005
R7449 GND.n3193 GND.n3192 9.3005
R7450 GND.n3198 GND.n2254 9.3005
R7451 GND.n3200 GND.n3199 9.3005
R7452 GND.n3201 GND.n1938 9.3005
R7453 GND.n2859 GND.n2357 9.3005
R7454 GND.n1527 GND.n1525 9.3005
R7455 GND.n3826 GND.n3823 9.3005
R7456 GND.n3827 GND.n3822 9.3005
R7457 GND.n3830 GND.n3821 9.3005
R7458 GND.n3831 GND.n3820 9.3005
R7459 GND.n3834 GND.n3819 9.3005
R7460 GND.n3835 GND.n3818 9.3005
R7461 GND.n3838 GND.n3817 9.3005
R7462 GND.n3839 GND.n3816 9.3005
R7463 GND.n3842 GND.n3815 9.3005
R7464 GND.n3844 GND.n3814 9.3005
R7465 GND.n3845 GND.n3813 9.3005
R7466 GND.n3846 GND.n3812 9.3005
R7467 GND.n3847 GND.n3811 9.3005
R7468 GND.n3808 GND.n1555 9.3005
R7469 GND.n3807 GND.n1557 9.3005
R7470 GND.n1578 GND.n1558 9.3005
R7471 GND.n1579 GND.n1577 9.3005
R7472 GND.n3795 GND.n1580 9.3005
R7473 GND.n3794 GND.n1581 9.3005
R7474 GND.n3793 GND.n1582 9.3005
R7475 GND.n1645 GND.n1583 9.3005
R7476 GND.n3710 GND.n1646 9.3005
R7477 GND.n3709 GND.n1647 9.3005
R7478 GND.n3708 GND.n1648 9.3005
R7479 GND.n2945 GND.n1649 9.3005
R7480 GND.n2948 GND.n2947 9.3005
R7481 GND.n2946 GND.n1676 9.3005
R7482 GND.n3689 GND.n1677 9.3005
R7483 GND.n3688 GND.n1678 9.3005
R7484 GND.n3687 GND.n1679 9.3005
R7485 GND.n2326 GND.n1680 9.3005
R7486 GND.n2327 GND.n2325 9.3005
R7487 GND.n2329 GND.n2328 9.3005
R7488 GND.n2323 GND.n2322 9.3005
R7489 GND.n3038 GND.n3037 9.3005
R7490 GND.n3039 GND.n2321 9.3005
R7491 GND.n3046 GND.n3040 9.3005
R7492 GND.n3045 GND.n3041 9.3005
R7493 GND.n3044 GND.n3043 9.3005
R7494 GND.n3042 GND.n2309 9.3005
R7495 GND.n2307 GND.n2306 9.3005
R7496 GND.n3067 GND.n3066 9.3005
R7497 GND.n3068 GND.n2305 9.3005
R7498 GND.n3070 GND.n3069 9.3005
R7499 GND.n2290 GND.n2289 9.3005
R7500 GND.n3086 GND.n3085 9.3005
R7501 GND.n3087 GND.n2288 9.3005
R7502 GND.n3098 GND.n3088 9.3005
R7503 GND.n3097 GND.n3089 9.3005
R7504 GND.n3096 GND.n3090 9.3005
R7505 GND.n3093 GND.n3092 9.3005
R7506 GND.n3091 GND.n1791 9.3005
R7507 GND.n3605 GND.n1792 9.3005
R7508 GND.n3604 GND.n1793 9.3005
R7509 GND.n3603 GND.n1794 9.3005
R7510 GND.n3166 GND.n1795 9.3005
R7511 GND.n3168 GND.n3167 9.3005
R7512 GND.n3165 GND.n3164 9.3005
R7513 GND.n3173 GND.n3172 9.3005
R7514 GND.n3174 GND.n3163 9.3005
R7515 GND.n3179 GND.n3175 9.3005
R7516 GND.n3178 GND.n3177 9.3005
R7517 GND.n3176 GND.n1877 9.3005
R7518 GND.n3565 GND.n1878 9.3005
R7519 GND.n3564 GND.n1879 9.3005
R7520 GND.n3563 GND.n1880 9.3005
R7521 GND.n1901 GND.n1881 9.3005
R7522 GND.n1902 GND.n1900 9.3005
R7523 GND.n3551 GND.n1903 9.3005
R7524 GND.n3550 GND.n3549 9.3005
R7525 GND.n3810 GND.n3809 9.3005
R7526 GND.n1905 GND.n1904 9.3005
R7527 GND.n3542 GND.n1918 9.3005
R7528 GND.n3541 GND.n1919 9.3005
R7529 GND.n3540 GND.n1920 9.3005
R7530 GND.n3537 GND.n1921 9.3005
R7531 GND.n3536 GND.n1922 9.3005
R7532 GND.n3533 GND.n1923 9.3005
R7533 GND.n3532 GND.n1924 9.3005
R7534 GND.n3529 GND.n1925 9.3005
R7535 GND.n3528 GND.n1926 9.3005
R7536 GND.n3525 GND.n1927 9.3005
R7537 GND.n3524 GND.n1928 9.3005
R7538 GND.n3521 GND.n1929 9.3005
R7539 GND.n3548 GND.n3547 9.3005
R7540 GND.n3217 GND.n3216 9.3005
R7541 GND.n3214 GND.n2253 9.3005
R7542 GND.n3213 GND.n3212 9.3005
R7543 GND.n3209 GND.n3206 9.3005
R7544 GND.n3205 GND.n3204 9.3005
R7545 GND.n3203 GND.n3202 9.3005
R7546 GND.n3520 GND.n1930 9.3005
R7547 GND.n3517 GND.n1934 9.3005
R7548 GND.n3516 GND.n1935 9.3005
R7549 GND.n3513 GND.n1936 9.3005
R7550 GND.n3512 GND.n1937 9.3005
R7551 GND.n3230 GND.n2248 9.3005
R7552 GND.n3227 GND.n3226 9.3005
R7553 GND.n3225 GND.n2251 9.3005
R7554 GND.n3224 GND.n3223 9.3005
R7555 GND.n3220 GND.n2252 9.3005
R7556 GND.n3234 GND.n3233 9.3005
R7557 GND.n3237 GND.n3236 9.3005
R7558 GND.n3238 GND.n2244 9.3005
R7559 GND.n3242 GND.n3241 9.3005
R7560 GND.n3243 GND.n2243 9.3005
R7561 GND.n3252 GND.n3244 9.3005
R7562 GND.n3251 GND.n3245 9.3005
R7563 GND.n3250 GND.n3246 9.3005
R7564 GND.n3249 GND.n3247 9.3005
R7565 GND.n7 GND.n5 9.3005
R7566 GND.n3235 GND.n2245 9.3005
R7567 GND.n5503 GND.n5502 9.3005
R7568 GND.n8 GND.n6 9.3005
R7569 GND.n2237 GND.n2236 9.3005
R7570 GND.n3336 GND.n2238 9.3005
R7571 GND.n3335 GND.n2239 9.3005
R7572 GND.n3334 GND.n2240 9.3005
R7573 GND.n3273 GND.n2241 9.3005
R7574 GND.n3324 GND.n3274 9.3005
R7575 GND.n3323 GND.n3275 9.3005
R7576 GND.n3322 GND.n3321 9.3005
R7577 GND.n3293 GND.n3292 9.3005
R7578 GND.n3287 GND.n3286 9.3005
R7579 GND.n3300 GND.n3299 9.3005
R7580 GND.n3301 GND.n3285 9.3005
R7581 GND.n3303 GND.n3302 9.3005
R7582 GND.n3283 GND.n3282 9.3005
R7583 GND.n3311 GND.n3310 9.3005
R7584 GND.n3312 GND.n3281 9.3005
R7585 GND.n3314 GND.n3313 9.3005
R7586 GND.n3315 GND.n3276 9.3005
R7587 GND.n3320 GND.n3319 9.3005
R7588 GND.n3291 GND.n3290 9.3005
R7589 GND.n255 GND.n254 9.3005
R7590 GND.n253 GND.n98 9.3005
R7591 GND.n252 GND.n251 9.3005
R7592 GND.n248 GND.n99 9.3005
R7593 GND.n245 GND.n100 9.3005
R7594 GND.n244 GND.n101 9.3005
R7595 GND.n241 GND.n102 9.3005
R7596 GND.n240 GND.n103 9.3005
R7597 GND.n237 GND.n104 9.3005
R7598 GND.n236 GND.n105 9.3005
R7599 GND.n233 GND.n109 9.3005
R7600 GND.n232 GND.n110 9.3005
R7601 GND.n229 GND.n111 9.3005
R7602 GND.n228 GND.n112 9.3005
R7603 GND.n225 GND.n113 9.3005
R7604 GND.n224 GND.n114 9.3005
R7605 GND.n221 GND.n115 9.3005
R7606 GND.n220 GND.n116 9.3005
R7607 GND.n217 GND.n117 9.3005
R7608 GND.n216 GND.n118 9.3005
R7609 GND.n213 GND.n119 9.3005
R7610 GND.n212 GND.n120 9.3005
R7611 GND.n209 GND.n121 9.3005
R7612 GND.n205 GND.n122 9.3005
R7613 GND.n202 GND.n123 9.3005
R7614 GND.n201 GND.n124 9.3005
R7615 GND.n198 GND.n125 9.3005
R7616 GND.n197 GND.n126 9.3005
R7617 GND.n194 GND.n127 9.3005
R7618 GND.n193 GND.n128 9.3005
R7619 GND.n190 GND.n129 9.3005
R7620 GND.n189 GND.n130 9.3005
R7621 GND.n186 GND.n131 9.3005
R7622 GND.n185 GND.n132 9.3005
R7623 GND.n182 GND.n133 9.3005
R7624 GND.n181 GND.n180 9.3005
R7625 GND.n179 GND.n134 9.3005
R7626 GND.n178 GND.n177 9.3005
R7627 GND.n174 GND.n139 9.3005
R7628 GND.n173 GND.n140 9.3005
R7629 GND.n170 GND.n141 9.3005
R7630 GND.n169 GND.n142 9.3005
R7631 GND.n166 GND.n143 9.3005
R7632 GND.n165 GND.n144 9.3005
R7633 GND.n162 GND.n145 9.3005
R7634 GND.n161 GND.n146 9.3005
R7635 GND.n158 GND.n147 9.3005
R7636 GND.n157 GND.n148 9.3005
R7637 GND.n154 GND.n153 9.3005
R7638 GND.n152 GND.n149 9.3005
R7639 GND.n256 GND.n97 9.3005
R7640 GND.n3398 GND.n3397 9.3005
R7641 GND.n2153 GND.n2152 9.3005
R7642 GND.n2177 GND.n2176 9.3005
R7643 GND.n3385 GND.n2178 9.3005
R7644 GND.n3384 GND.n2179 9.3005
R7645 GND.n3383 GND.n2180 9.3005
R7646 GND.n3259 GND.n2181 9.3005
R7647 GND.n3260 GND.n2224 9.3005
R7648 GND.n3366 GND.n2225 9.3005
R7649 GND.n3365 GND.n2226 9.3005
R7650 GND.n3364 GND.n2227 9.3005
R7651 GND.n3268 GND.n2228 9.3005
R7652 GND.n3269 GND.n35 9.3005
R7653 GND.n5491 GND.n36 9.3005
R7654 GND.n5490 GND.n37 9.3005
R7655 GND.n5489 GND.n38 9.3005
R7656 GND.n3272 GND.n39 9.3005
R7657 GND.n5479 GND.n56 9.3005
R7658 GND.n5478 GND.n5477 9.3005
R7659 GND.n3399 GND.n2151 9.3005
R7660 GND.n3397 GND.n3396 9.3005
R7661 GND.n3395 GND.n2153 9.3005
R7662 GND.n2177 GND.n2154 9.3005
R7663 GND.n2242 GND.n2178 9.3005
R7664 GND.n3256 GND.n2179 9.3005
R7665 GND.n3257 GND.n2180 9.3005
R7666 GND.n3259 GND.n3258 9.3005
R7667 GND.n3262 GND.n3260 9.3005
R7668 GND.n3263 GND.n2225 9.3005
R7669 GND.n3264 GND.n2226 9.3005
R7670 GND.n3265 GND.n2227 9.3005
R7671 GND.n3268 GND.n3267 9.3005
R7672 GND.n3270 GND.n3269 9.3005
R7673 GND.n3271 GND.n36 9.3005
R7674 GND.n3330 GND.n37 9.3005
R7675 GND.n3329 GND.n38 9.3005
R7676 GND.n3328 GND.n3272 9.3005
R7677 GND.n58 GND.n56 9.3005
R7678 GND.n5477 GND.n5476 9.3005
R7679 GND.n2151 GND.n2145 9.3005
R7680 GND.n3408 GND.n3407 9.3005
R7681 GND.n3409 GND.n2136 9.3005
R7682 GND.n3412 GND.n2135 9.3005
R7683 GND.n3413 GND.n2134 9.3005
R7684 GND.n3416 GND.n2133 9.3005
R7685 GND.n3417 GND.n2132 9.3005
R7686 GND.n3420 GND.n2131 9.3005
R7687 GND.n3421 GND.n2130 9.3005
R7688 GND.n3424 GND.n2129 9.3005
R7689 GND.n3425 GND.n2128 9.3005
R7690 GND.n3428 GND.n2127 9.3005
R7691 GND.n3430 GND.n2126 9.3005
R7692 GND.n3432 GND.n2121 9.3005
R7693 GND.n3435 GND.n2120 9.3005
R7694 GND.n3436 GND.n2119 9.3005
R7695 GND.n3439 GND.n2118 9.3005
R7696 GND.n3440 GND.n2117 9.3005
R7697 GND.n3443 GND.n2116 9.3005
R7698 GND.n3444 GND.n2115 9.3005
R7699 GND.n3447 GND.n2114 9.3005
R7700 GND.n3448 GND.n2113 9.3005
R7701 GND.n3451 GND.n2112 9.3005
R7702 GND.n3452 GND.n2111 9.3005
R7703 GND.n3455 GND.n2110 9.3005
R7704 GND.n3457 GND.n2004 9.3005
R7705 GND.n3460 GND.n2003 9.3005
R7706 GND.n3461 GND.n2002 9.3005
R7707 GND.n3464 GND.n2001 9.3005
R7708 GND.n3465 GND.n2000 9.3005
R7709 GND.n3468 GND.n1999 9.3005
R7710 GND.n3469 GND.n1998 9.3005
R7711 GND.n3472 GND.n1997 9.3005
R7712 GND.n3473 GND.n1996 9.3005
R7713 GND.n3476 GND.n1995 9.3005
R7714 GND.n3477 GND.n1994 9.3005
R7715 GND.n3480 GND.n1990 9.3005
R7716 GND.n3481 GND.n1989 9.3005
R7717 GND.n3484 GND.n1988 9.3005
R7718 GND.n3485 GND.n1987 9.3005
R7719 GND.n3488 GND.n1986 9.3005
R7720 GND.n3489 GND.n1985 9.3005
R7721 GND.n3492 GND.n1984 9.3005
R7722 GND.n3494 GND.n1983 9.3005
R7723 GND.n3495 GND.n1982 9.3005
R7724 GND.n3496 GND.n1981 9.3005
R7725 GND.n3497 GND.n1980 9.3005
R7726 GND.n3431 GND.n2123 9.3005
R7727 GND.n3406 GND.n2141 9.3005
R7728 GND.n3405 GND.n3404 9.3005
R7729 GND.n2165 GND.n2162 9.3005
R7730 GND.n3391 GND.n2166 9.3005
R7731 GND.n3390 GND.n2167 9.3005
R7732 GND.n3389 GND.n19 9.3005
R7733 GND.n26 GND.n18 9.3005
R7734 GND.n5485 GND.n46 9.3005
R7735 GND.n5484 GND.n47 9.3005
R7736 GND.n5483 GND.n48 9.3005
R7737 GND.n96 GND.n49 9.3005
R7738 GND.n2164 GND.n2163 9.3005
R7739 GND.n5496 GND.n23 9.3005
R7740 GND.n5496 GND.n5495 9.3005
R7741 GND.n2494 GND.n2447 9.3005
R7742 GND.n2493 GND.n2454 9.3005
R7743 GND.n2457 GND.n2455 9.3005
R7744 GND.n2489 GND.n2458 9.3005
R7745 GND.n2488 GND.n2459 9.3005
R7746 GND.n2487 GND.n2460 9.3005
R7747 GND.n2463 GND.n2461 9.3005
R7748 GND.n2481 GND.n2464 9.3005
R7749 GND.n2480 GND.n2465 9.3005
R7750 GND.n2479 GND.n2466 9.3005
R7751 GND.n2468 GND.n2467 9.3005
R7752 GND.n2471 GND.n2470 9.3005
R7753 GND.n2469 GND.n1565 9.3005
R7754 GND.n3802 GND.n1566 9.3005
R7755 GND.n3801 GND.n1567 9.3005
R7756 GND.n3800 GND.n1568 9.3005
R7757 GND.n2880 GND.n1569 9.3005
R7758 GND.n2882 GND.n2881 9.3005
R7759 GND.n2886 GND.n2885 9.3005
R7760 GND.n2887 GND.n2879 9.3005
R7761 GND.n2890 GND.n2889 9.3005
R7762 GND.n2888 GND.n1657 9.3005
R7763 GND.n3703 GND.n1658 9.3005
R7764 GND.n3702 GND.n1659 9.3005
R7765 GND.n3701 GND.n1660 9.3005
R7766 GND.n1688 GND.n1661 9.3005
R7767 GND.n1691 GND.n1690 9.3005
R7768 GND.n1692 GND.n1687 9.3005
R7769 GND.n3682 GND.n1693 9.3005
R7770 GND.n3681 GND.n1694 9.3005
R7771 GND.n3680 GND.n1695 9.3005
R7772 GND.n1710 GND.n1696 9.3005
R7773 GND.n3668 GND.n1711 9.3005
R7774 GND.n3667 GND.n1712 9.3005
R7775 GND.n3666 GND.n1713 9.3005
R7776 GND.n1727 GND.n1714 9.3005
R7777 GND.n3654 GND.n1728 9.3005
R7778 GND.n3653 GND.n1729 9.3005
R7779 GND.n3652 GND.n1730 9.3005
R7780 GND.n1745 GND.n1731 9.3005
R7781 GND.n3640 GND.n1746 9.3005
R7782 GND.n3639 GND.n1747 9.3005
R7783 GND.n3638 GND.n1748 9.3005
R7784 GND.n1762 GND.n1749 9.3005
R7785 GND.n3626 GND.n1763 9.3005
R7786 GND.n3625 GND.n1764 9.3005
R7787 GND.n3624 GND.n1765 9.3005
R7788 GND.n1780 GND.n1766 9.3005
R7789 GND.n3612 GND.n1781 9.3005
R7790 GND.n3611 GND.n1782 9.3005
R7791 GND.n3610 GND.n1783 9.3005
R7792 GND.n1810 GND.n1784 9.3005
R7793 GND.n1813 GND.n1812 9.3005
R7794 GND.n1814 GND.n1809 9.3005
R7795 GND.n3591 GND.n1815 9.3005
R7796 GND.n3590 GND.n1816 9.3005
R7797 GND.n3589 GND.n1817 9.3005
R7798 GND.n1865 GND.n1818 9.3005
R7799 GND.n1866 GND.n1864 9.3005
R7800 GND.n3572 GND.n1867 9.3005
R7801 GND.n3571 GND.n1868 9.3005
R7802 GND.n3570 GND.n1869 9.3005
R7803 GND.n1888 GND.n1870 9.3005
R7804 GND.n1889 GND.n1887 9.3005
R7805 GND.n3558 GND.n1890 9.3005
R7806 GND.n3557 GND.n1891 9.3005
R7807 GND.n3556 GND.n1892 9.3005
R7808 GND.n1940 GND.n1893 9.3005
R7809 GND.n3506 GND.n1941 9.3005
R7810 GND.n3505 GND.n1942 9.3005
R7811 GND.n3504 GND.n1943 9.3005
R7812 GND.n2200 GND.n1944 9.3005
R7813 GND.n2201 GND.n2199 9.3005
R7814 GND.n2203 GND.n2202 9.3005
R7815 GND.n2198 GND.n2197 9.3005
R7816 GND.n2208 GND.n2207 9.3005
R7817 GND.n2209 GND.n2196 9.3005
R7818 GND.n2212 GND.n2211 9.3005
R7819 GND.n2210 GND.n2194 9.3005
R7820 GND.n3352 GND.n3344 9.3005
R7821 GND.n3351 GND.n3345 9.3005
R7822 GND.n3348 GND.n3347 9.3005
R7823 GND.n3346 GND.n64 9.3005
R7824 GND.n5471 GND.n65 9.3005
R7825 GND.n5470 GND.n66 9.3005
R7826 GND.n5469 GND.n67 9.3005
R7827 GND.n261 GND.n68 9.3005
R7828 GND.n5463 GND.n262 9.3005
R7829 GND.n5462 GND.n263 9.3005
R7830 GND.n5461 GND.n264 9.3005
R7831 GND.n269 GND.n265 9.3005
R7832 GND.n5455 GND.n270 9.3005
R7833 GND.n5454 GND.n271 9.3005
R7834 GND.n5453 GND.n272 9.3005
R7835 GND.n277 GND.n273 9.3005
R7836 GND.n5447 GND.n278 9.3005
R7837 GND.n5446 GND.n279 9.3005
R7838 GND.n5445 GND.n280 9.3005
R7839 GND.n285 GND.n281 9.3005
R7840 GND.n5439 GND.n286 9.3005
R7841 GND.n5438 GND.n287 9.3005
R7842 GND.n5437 GND.n288 9.3005
R7843 GND.n293 GND.n289 9.3005
R7844 GND.n5431 GND.n294 9.3005
R7845 GND.n5430 GND.n295 9.3005
R7846 GND.n5429 GND.n296 9.3005
R7847 GND.n301 GND.n297 9.3005
R7848 GND.n5423 GND.n302 9.3005
R7849 GND.n5422 GND.n303 9.3005
R7850 GND.n5421 GND.n304 9.3005
R7851 GND.n309 GND.n305 9.3005
R7852 GND.n5415 GND.n310 9.3005
R7853 GND.n5414 GND.n311 9.3005
R7854 GND.n5413 GND.n312 9.3005
R7855 GND.n317 GND.n313 9.3005
R7856 GND.n5407 GND.n318 9.3005
R7857 GND.n5406 GND.n319 9.3005
R7858 GND.n5405 GND.n320 9.3005
R7859 GND.n325 GND.n321 9.3005
R7860 GND.n5399 GND.n326 9.3005
R7861 GND.n5398 GND.n327 9.3005
R7862 GND.n5397 GND.n328 9.3005
R7863 GND.n333 GND.n329 9.3005
R7864 GND.n5391 GND.n334 9.3005
R7865 GND.n5390 GND.n335 9.3005
R7866 GND.n5389 GND.n336 9.3005
R7867 GND.n341 GND.n337 9.3005
R7868 GND.n5383 GND.n342 9.3005
R7869 GND.n5382 GND.n343 9.3005
R7870 GND.n5381 GND.n344 9.3005
R7871 GND.n349 GND.n345 9.3005
R7872 GND.n5375 GND.n350 9.3005
R7873 GND.n5374 GND.n351 9.3005
R7874 GND.n5373 GND.n352 9.3005
R7875 GND.n357 GND.n353 9.3005
R7876 GND.n5367 GND.n358 9.3005
R7877 GND.n5366 GND.n359 9.3005
R7878 GND.n5365 GND.n360 9.3005
R7879 GND.n365 GND.n361 9.3005
R7880 GND.n5359 GND.n366 9.3005
R7881 GND.n5358 GND.n367 9.3005
R7882 GND.n5357 GND.n368 9.3005
R7883 GND.n373 GND.n369 9.3005
R7884 GND.n5351 GND.n374 9.3005
R7885 GND.n5350 GND.n375 9.3005
R7886 GND.n5349 GND.n376 9.3005
R7887 GND.n381 GND.n377 9.3005
R7888 GND.n5343 GND.n382 9.3005
R7889 GND.n5342 GND.n383 9.3005
R7890 GND.n5341 GND.n384 9.3005
R7891 GND.n389 GND.n385 9.3005
R7892 GND.n5335 GND.n390 9.3005
R7893 GND.n5334 GND.n391 9.3005
R7894 GND.n5333 GND.n392 9.3005
R7895 GND.n397 GND.n393 9.3005
R7896 GND.n5327 GND.n398 9.3005
R7897 GND.n5326 GND.n399 9.3005
R7898 GND.n5325 GND.n400 9.3005
R7899 GND.n405 GND.n401 9.3005
R7900 GND.n5319 GND.n406 9.3005
R7901 GND.n5318 GND.n407 9.3005
R7902 GND.n5317 GND.n408 9.3005
R7903 GND.n413 GND.n409 9.3005
R7904 GND.n5311 GND.n414 9.3005
R7905 GND.n5310 GND.n415 9.3005
R7906 GND.n5309 GND.n416 9.3005
R7907 GND.n421 GND.n417 9.3005
R7908 GND.n5303 GND.n422 9.3005
R7909 GND.n5302 GND.n423 9.3005
R7910 GND.n5301 GND.n424 9.3005
R7911 GND.n429 GND.n425 9.3005
R7912 GND.n5295 GND.n430 9.3005
R7913 GND.n5294 GND.n431 9.3005
R7914 GND.n5293 GND.n432 9.3005
R7915 GND.n437 GND.n433 9.3005
R7916 GND.n5287 GND.n438 9.3005
R7917 GND.n5286 GND.n439 9.3005
R7918 GND.n5285 GND.n440 9.3005
R7919 GND.n445 GND.n441 9.3005
R7920 GND.n5279 GND.n446 9.3005
R7921 GND.n5278 GND.n447 9.3005
R7922 GND.n5277 GND.n448 9.3005
R7923 GND.n453 GND.n449 9.3005
R7924 GND.n5271 GND.n454 9.3005
R7925 GND.n5270 GND.n455 9.3005
R7926 GND.n5269 GND.n456 9.3005
R7927 GND.n461 GND.n457 9.3005
R7928 GND.n5263 GND.n462 9.3005
R7929 GND.n5262 GND.n463 9.3005
R7930 GND.n5261 GND.n464 9.3005
R7931 GND.n2718 GND.n2717 9.3005
R7932 GND.n2716 GND.n2543 9.3005
R7933 GND.n2715 GND.n2714 9.3005
R7934 GND.n2545 GND.n2544 9.3005
R7935 GND.n2708 GND.n2707 9.3005
R7936 GND.n2706 GND.n2547 9.3005
R7937 GND.n2705 GND.n2704 9.3005
R7938 GND.n2549 GND.n2548 9.3005
R7939 GND.n2698 GND.n2697 9.3005
R7940 GND.n2696 GND.n2551 9.3005
R7941 GND.n2695 GND.n2694 9.3005
R7942 GND.n2553 GND.n2552 9.3005
R7943 GND.n2684 GND.n2555 9.3005
R7944 GND.n2683 GND.n2682 9.3005
R7945 GND.n2557 GND.n2556 9.3005
R7946 GND.n2676 GND.n2675 9.3005
R7947 GND.n2674 GND.n2559 9.3005
R7948 GND.n2673 GND.n2672 9.3005
R7949 GND.n2561 GND.n2560 9.3005
R7950 GND.n2666 GND.n2665 9.3005
R7951 GND.n2664 GND.n2563 9.3005
R7952 GND.n2663 GND.n2662 9.3005
R7953 GND.n2565 GND.n2564 9.3005
R7954 GND.n2656 GND.n2655 9.3005
R7955 GND.n2652 GND.n2570 9.3005
R7956 GND.n2644 GND.n2571 9.3005
R7957 GND.n2646 GND.n2645 9.3005
R7958 GND.n2643 GND.n2573 9.3005
R7959 GND.n2642 GND.n2641 9.3005
R7960 GND.n2575 GND.n2574 9.3005
R7961 GND.n2635 GND.n2634 9.3005
R7962 GND.n2633 GND.n2577 9.3005
R7963 GND.n2632 GND.n2631 9.3005
R7964 GND.n2579 GND.n2578 9.3005
R7965 GND.n2625 GND.n2624 9.3005
R7966 GND.n2623 GND.n2581 9.3005
R7967 GND.n2622 GND.n2621 9.3005
R7968 GND.n2583 GND.n2582 9.3005
R7969 GND.n2615 GND.n2614 9.3005
R7970 GND.n2613 GND.n2588 9.3005
R7971 GND.n2612 GND.n2611 9.3005
R7972 GND.n2590 GND.n2589 9.3005
R7973 GND.n2605 GND.n2604 9.3005
R7974 GND.n2603 GND.n2592 9.3005
R7975 GND.n2602 GND.n2601 9.3005
R7976 GND.n2596 GND.n2593 9.3005
R7977 GND.n2595 GND.n2594 9.3005
R7978 GND.n2654 GND.n2653 9.3005
R7979 GND.n2688 GND.n2685 9.3005
R7980 GND.n2541 GND.n2538 9.3005
R7981 GND.n2724 GND.n2723 9.3005
R7982 GND.n3984 GND.n1364 9.3005
R7983 GND.n3983 GND.n1365 9.3005
R7984 GND.n2429 GND.n1366 9.3005
R7985 GND.n2431 GND.n2430 9.3005
R7986 GND.n2831 GND.n2830 9.3005
R7987 GND.n2832 GND.n2386 9.3005
R7988 GND.n2834 GND.n2833 9.3005
R7989 GND.n1419 GND.n1418 9.3005
R7990 GND.n3948 GND.n3947 9.3005
R7991 GND.n3985 GND.n1363 9.3005
R7992 GND.n2783 GND.n2387 9.3005
R7993 GND.n2388 GND.n2387 9.3005
R7994 GND.n4199 GND.n1144 9.3005
R7995 GND.n4198 GND.n1145 9.3005
R7996 GND.n1150 GND.n1146 9.3005
R7997 GND.n4192 GND.n1151 9.3005
R7998 GND.n4191 GND.n1152 9.3005
R7999 GND.n4190 GND.n1153 9.3005
R8000 GND.n1158 GND.n1154 9.3005
R8001 GND.n4184 GND.n1159 9.3005
R8002 GND.n4183 GND.n1160 9.3005
R8003 GND.n4182 GND.n1161 9.3005
R8004 GND.n1166 GND.n1162 9.3005
R8005 GND.n4176 GND.n1167 9.3005
R8006 GND.n4175 GND.n1168 9.3005
R8007 GND.n4174 GND.n1169 9.3005
R8008 GND.n1174 GND.n1170 9.3005
R8009 GND.n4168 GND.n1175 9.3005
R8010 GND.n4167 GND.n1176 9.3005
R8011 GND.n4166 GND.n1177 9.3005
R8012 GND.n1182 GND.n1178 9.3005
R8013 GND.n4160 GND.n1183 9.3005
R8014 GND.n4159 GND.n1184 9.3005
R8015 GND.n4158 GND.n1185 9.3005
R8016 GND.n1190 GND.n1186 9.3005
R8017 GND.n4152 GND.n1191 9.3005
R8018 GND.n4151 GND.n1192 9.3005
R8019 GND.n4150 GND.n1193 9.3005
R8020 GND.n1198 GND.n1194 9.3005
R8021 GND.n4144 GND.n1199 9.3005
R8022 GND.n4143 GND.n1200 9.3005
R8023 GND.n4142 GND.n1201 9.3005
R8024 GND.n1206 GND.n1202 9.3005
R8025 GND.n4136 GND.n1207 9.3005
R8026 GND.n4135 GND.n1208 9.3005
R8027 GND.n4134 GND.n1209 9.3005
R8028 GND.n1214 GND.n1210 9.3005
R8029 GND.n4128 GND.n1215 9.3005
R8030 GND.n4127 GND.n1216 9.3005
R8031 GND.n4126 GND.n1217 9.3005
R8032 GND.n1222 GND.n1218 9.3005
R8033 GND.n4120 GND.n1223 9.3005
R8034 GND.n4119 GND.n1224 9.3005
R8035 GND.n4118 GND.n1225 9.3005
R8036 GND.n1230 GND.n1226 9.3005
R8037 GND.n4112 GND.n1231 9.3005
R8038 GND.n4111 GND.n1232 9.3005
R8039 GND.n4110 GND.n1233 9.3005
R8040 GND.n1238 GND.n1234 9.3005
R8041 GND.n4104 GND.n1239 9.3005
R8042 GND.n4103 GND.n1240 9.3005
R8043 GND.n4102 GND.n1241 9.3005
R8044 GND.n1246 GND.n1242 9.3005
R8045 GND.n4096 GND.n1247 9.3005
R8046 GND.n4095 GND.n1248 9.3005
R8047 GND.n4094 GND.n1249 9.3005
R8048 GND.n1254 GND.n1250 9.3005
R8049 GND.n4088 GND.n1255 9.3005
R8050 GND.n4087 GND.n1256 9.3005
R8051 GND.n4086 GND.n1257 9.3005
R8052 GND.n1262 GND.n1258 9.3005
R8053 GND.n4080 GND.n1263 9.3005
R8054 GND.n4079 GND.n1264 9.3005
R8055 GND.n4078 GND.n1265 9.3005
R8056 GND.n1270 GND.n1266 9.3005
R8057 GND.n4072 GND.n1271 9.3005
R8058 GND.n4071 GND.n1272 9.3005
R8059 GND.n4070 GND.n1273 9.3005
R8060 GND.n1278 GND.n1274 9.3005
R8061 GND.n4064 GND.n1279 9.3005
R8062 GND.n4063 GND.n1280 9.3005
R8063 GND.n4062 GND.n1281 9.3005
R8064 GND.n1286 GND.n1282 9.3005
R8065 GND.n4056 GND.n1287 9.3005
R8066 GND.n4055 GND.n1288 9.3005
R8067 GND.n4054 GND.n1289 9.3005
R8068 GND.n1294 GND.n1290 9.3005
R8069 GND.n4048 GND.n1295 9.3005
R8070 GND.n4047 GND.n1296 9.3005
R8071 GND.n4046 GND.n1297 9.3005
R8072 GND.n1302 GND.n1298 9.3005
R8073 GND.n4040 GND.n1303 9.3005
R8074 GND.n4039 GND.n1304 9.3005
R8075 GND.n4038 GND.n1305 9.3005
R8076 GND.n1310 GND.n1306 9.3005
R8077 GND.n4032 GND.n1311 9.3005
R8078 GND.n4031 GND.n1312 9.3005
R8079 GND.n4030 GND.n1313 9.3005
R8080 GND.n1318 GND.n1314 9.3005
R8081 GND.n4024 GND.n1319 9.3005
R8082 GND.n4023 GND.n1320 9.3005
R8083 GND.n4022 GND.n1321 9.3005
R8084 GND.n1326 GND.n1322 9.3005
R8085 GND.n4016 GND.n1327 9.3005
R8086 GND.n4015 GND.n1328 9.3005
R8087 GND.n4014 GND.n1329 9.3005
R8088 GND.n1334 GND.n1330 9.3005
R8089 GND.n4008 GND.n1335 9.3005
R8090 GND.n4007 GND.n1336 9.3005
R8091 GND.n4006 GND.n1337 9.3005
R8092 GND.n1342 GND.n1338 9.3005
R8093 GND.n4000 GND.n1343 9.3005
R8094 GND.n3999 GND.n1344 9.3005
R8095 GND.n3998 GND.n1345 9.3005
R8096 GND.n1350 GND.n1346 9.3005
R8097 GND.n3992 GND.n1351 9.3005
R8098 GND.n3991 GND.n1352 9.3005
R8099 GND.n3990 GND.n1353 9.3005
R8100 GND.n2441 GND.n1354 9.3005
R8101 GND.n2442 GND.n2440 9.3005
R8102 GND.n2515 GND.n2443 9.3005
R8103 GND.n2514 GND.n2444 9.3005
R8104 GND.n4200 GND.n1143 9.3005
R8105 GND.n4206 GND.n1137 9.3005
R8106 GND.n4207 GND.n1136 9.3005
R8107 GND.n4208 GND.n1135 9.3005
R8108 GND.n1134 GND.n1130 9.3005
R8109 GND.n4214 GND.n1129 9.3005
R8110 GND.n4215 GND.n1128 9.3005
R8111 GND.n4216 GND.n1127 9.3005
R8112 GND.n1126 GND.n1122 9.3005
R8113 GND.n4222 GND.n1121 9.3005
R8114 GND.n4223 GND.n1120 9.3005
R8115 GND.n4224 GND.n1119 9.3005
R8116 GND.n1118 GND.n1114 9.3005
R8117 GND.n4230 GND.n1113 9.3005
R8118 GND.n4231 GND.n1112 9.3005
R8119 GND.n4232 GND.n1111 9.3005
R8120 GND.n1110 GND.n1106 9.3005
R8121 GND.n4238 GND.n1105 9.3005
R8122 GND.n4239 GND.n1104 9.3005
R8123 GND.n4240 GND.n1103 9.3005
R8124 GND.n1102 GND.n1098 9.3005
R8125 GND.n4246 GND.n1097 9.3005
R8126 GND.n4247 GND.n1096 9.3005
R8127 GND.n4248 GND.n1095 9.3005
R8128 GND.n1094 GND.n1090 9.3005
R8129 GND.n4254 GND.n1089 9.3005
R8130 GND.n4255 GND.n1088 9.3005
R8131 GND.n4256 GND.n1087 9.3005
R8132 GND.n1086 GND.n1082 9.3005
R8133 GND.n4262 GND.n1081 9.3005
R8134 GND.n4263 GND.n1080 9.3005
R8135 GND.n4264 GND.n1079 9.3005
R8136 GND.n1078 GND.n1074 9.3005
R8137 GND.n4270 GND.n1073 9.3005
R8138 GND.n4271 GND.n1072 9.3005
R8139 GND.n4272 GND.n1071 9.3005
R8140 GND.n1070 GND.n1066 9.3005
R8141 GND.n4278 GND.n1065 9.3005
R8142 GND.n4279 GND.n1064 9.3005
R8143 GND.n4280 GND.n1063 9.3005
R8144 GND.n1062 GND.n1058 9.3005
R8145 GND.n4286 GND.n1057 9.3005
R8146 GND.n4287 GND.n1056 9.3005
R8147 GND.n4288 GND.n1055 9.3005
R8148 GND.n1054 GND.n1050 9.3005
R8149 GND.n4294 GND.n1049 9.3005
R8150 GND.n4295 GND.n1048 9.3005
R8151 GND.n4296 GND.n1047 9.3005
R8152 GND.n1046 GND.n1042 9.3005
R8153 GND.n4302 GND.n1041 9.3005
R8154 GND.n4303 GND.n1040 9.3005
R8155 GND.n4304 GND.n1039 9.3005
R8156 GND.n1038 GND.n1034 9.3005
R8157 GND.n4310 GND.n1033 9.3005
R8158 GND.n4311 GND.n1032 9.3005
R8159 GND.n4312 GND.n1031 9.3005
R8160 GND.n1142 GND.n1138 9.3005
R8161 GND.n2790 GND.n2418 9.3005
R8162 GND.n2399 GND.n2398 9.3005
R8163 GND.n2813 GND.n2812 9.3005
R8164 GND.n2814 GND.n2396 9.3005
R8165 GND.n2822 GND.n2821 9.3005
R8166 GND.n2820 GND.n2397 9.3005
R8167 GND.n2819 GND.n2818 9.3005
R8168 GND.n2815 GND.n2379 9.3005
R8169 GND.n2841 GND.n2378 9.3005
R8170 GND.n2843 GND.n2842 9.3005
R8171 GND.n2855 GND.n2360 9.3005
R8172 GND.n2854 GND.n2853 9.3005
R8173 GND.n2852 GND.n2370 9.3005
R8174 GND.n2851 GND.n2850 9.3005
R8175 GND.n2849 GND.n2371 9.3005
R8176 GND.n2847 GND.n2844 9.3005
R8177 GND.n3858 GND.n3857 9.3005
R8178 GND.n3856 GND.n3855 9.3005
R8179 GND.n1540 GND.n1539 9.3005
R8180 GND.n2361 GND.n2359 9.3005
R8181 GND.n2857 GND.n2856 9.3005
R8182 GND.n1534 GND.n1532 9.3005
R8183 GND.n1533 GND.n1531 9.3005
R8184 GND.n3860 GND.n3859 9.3005
R8185 GND.n3861 GND.n1526 9.3005
R8186 GND.n3866 GND.n3865 9.3005
R8187 GND.n3854 GND.n3853 9.3005
R8188 GND.n3914 GND.n1449 9.3005
R8189 GND.n3915 GND.n1446 9.3005
R8190 GND.n3917 GND.n3916 9.3005
R8191 GND.n3918 GND.n1445 9.3005
R8192 GND.n3920 GND.n3919 9.3005
R8193 GND.n3921 GND.n1441 9.3005
R8194 GND.n3923 GND.n3922 9.3005
R8195 GND.n3924 GND.n1440 9.3005
R8196 GND.n3926 GND.n3925 9.3005
R8197 GND.n3927 GND.n1436 9.3005
R8198 GND.n3929 GND.n3928 9.3005
R8199 GND.n3931 GND.n3930 9.3005
R8200 GND.n3932 GND.n1429 9.3005
R8201 GND.n3934 GND.n3933 9.3005
R8202 GND.n3935 GND.n1428 9.3005
R8203 GND.n3937 GND.n3936 9.3005
R8204 GND.n3938 GND.n1424 9.3005
R8205 GND.n3940 GND.n3939 9.3005
R8206 GND.n3941 GND.n1423 9.3005
R8207 GND.n3943 GND.n3942 9.3005
R8208 GND.n3944 GND.n1420 9.3005
R8209 GND.n3946 GND.n3945 9.3005
R8210 GND.n3908 GND.n3907 9.3005
R8211 GND.n3906 GND.n1469 9.3005
R8212 GND.n3905 GND.n3904 9.3005
R8213 GND.n3903 GND.n1471 9.3005
R8214 GND.n3902 GND.n3901 9.3005
R8215 GND.n3900 GND.n1477 9.3005
R8216 GND.n3899 GND.n3898 9.3005
R8217 GND.n3897 GND.n1478 9.3005
R8218 GND.n3896 GND.n3895 9.3005
R8219 GND.n3894 GND.n1485 9.3005
R8220 GND.n3893 GND.n3892 9.3005
R8221 GND.n3891 GND.n1486 9.3005
R8222 GND.n3890 GND.n1493 9.3005
R8223 GND.n3889 GND.n3888 9.3005
R8224 GND.n3887 GND.n1497 9.3005
R8225 GND.n3886 GND.n3885 9.3005
R8226 GND.n3884 GND.n1498 9.3005
R8227 GND.n3883 GND.n3882 9.3005
R8228 GND.n3881 GND.n1505 9.3005
R8229 GND.n3880 GND.n3879 9.3005
R8230 GND.n3878 GND.n1506 9.3005
R8231 GND.n3877 GND.n3876 9.3005
R8232 GND.n3875 GND.n1513 9.3005
R8233 GND.n3874 GND.n3873 9.3005
R8234 GND.n3872 GND.n1514 9.3005
R8235 GND.n3871 GND.n1522 9.3005
R8236 GND.n3870 GND.n3869 9.3005
R8237 GND.n1375 GND.n1373 9.3005
R8238 GND.n3979 GND.n3978 9.3005
R8239 GND.n1376 GND.n1374 9.3005
R8240 GND.n3974 GND.n1381 9.3005
R8241 GND.n3973 GND.n1382 9.3005
R8242 GND.n3972 GND.n1383 9.3005
R8243 GND.n2424 GND.n1384 9.3005
R8244 GND.n3968 GND.n1389 9.3005
R8245 GND.n3967 GND.n1390 9.3005
R8246 GND.n3966 GND.n1391 9.3005
R8247 GND.n2797 GND.n1392 9.3005
R8248 GND.n3962 GND.n1397 9.3005
R8249 GND.n3961 GND.n1398 9.3005
R8250 GND.n3960 GND.n1399 9.3005
R8251 GND.n2826 GND.n1400 9.3005
R8252 GND.n3956 GND.n1405 9.3005
R8253 GND.n3955 GND.n1406 9.3005
R8254 GND.n3954 GND.n1407 9.3005
R8255 GND.n1414 GND.n1408 9.3005
R8256 GND.n2727 GND.n2725 9.3005
R8257 GND.n1377 GND.n1375 9.3005
R8258 GND.n3978 GND.n3977 9.3005
R8259 GND.n3976 GND.n1376 9.3005
R8260 GND.n3975 GND.n3974 9.3005
R8261 GND.n3973 GND.n1380 9.3005
R8262 GND.n3972 GND.n3971 9.3005
R8263 GND.n3970 GND.n1384 9.3005
R8264 GND.n3969 GND.n3968 9.3005
R8265 GND.n3967 GND.n1388 9.3005
R8266 GND.n3966 GND.n3965 9.3005
R8267 GND.n3964 GND.n1392 9.3005
R8268 GND.n3963 GND.n3962 9.3005
R8269 GND.n3961 GND.n1396 9.3005
R8270 GND.n3960 GND.n3959 9.3005
R8271 GND.n3958 GND.n1400 9.3005
R8272 GND.n3957 GND.n3956 9.3005
R8273 GND.n3955 GND.n1404 9.3005
R8274 GND.n3954 GND.n3953 9.3005
R8275 GND.n3952 GND.n1408 9.3005
R8276 GND.n2727 GND.n2726 9.3005
R8277 GND.n2527 GND.n2523 9.3005
R8278 GND.n2751 GND.n2750 9.3005
R8279 GND.n2749 GND.n2529 9.3005
R8280 GND.n2748 GND.n2747 9.3005
R8281 GND.n2531 GND.n2530 9.3005
R8282 GND.n2741 GND.n2740 9.3005
R8283 GND.n2739 GND.n2533 9.3005
R8284 GND.n2738 GND.n2737 9.3005
R8285 GND.n2535 GND.n2534 9.3005
R8286 GND.n2731 GND.n2730 9.3005
R8287 GND.n2729 GND.n2537 9.3005
R8288 GND.n2757 GND.n2756 9.3005
R8289 GND.n2763 GND.n2522 9.3005
R8290 GND.n2765 GND.n2764 9.3005
R8291 GND.n2766 GND.n2520 9.3005
R8292 GND.n2769 GND.n2768 9.3005
R8293 GND.n2767 GND.n2521 9.3005
R8294 GND.n2420 GND.n2419 9.3005
R8295 GND.n2788 GND.n2787 9.3005
R8296 GND.n2789 GND.n2417 9.3005
R8297 GND.n2793 GND.n2792 9.3005
R8298 GND.n2759 GND.n2758 9.3005
R8299 GND.n2966 GND.n2965 8.8049
R8300 GND.n2337 GND.t136 8.8049
R8301 GND.n3664 GND.n3663 8.8049
R8302 GND.n3629 GND.n3628 8.8049
R8303 GND.n3111 GND.t134 8.8049
R8304 GND.n2268 GND.n2267 8.8049
R8305 GND.n3890 GND.n3889 8.72777
R8306 GND.n3431 GND.n3430 8.72777
R8307 GND.n181 GND.n134 8.72777
R8308 GND.n2688 GND.n2553 8.72777
R8309 GND.t39 GND.n1562 8.0712
R8310 GND.n3713 GND.n3712 8.0712
R8311 GND.t3 GND.n1651 8.0712
R8312 GND.n2955 GND.n1664 8.0712
R8313 GND.n3016 GND.n1725 8.0712
R8314 GND.n3072 GND.n1751 8.0712
R8315 GND.n3135 GND.n3134 8.0712
R8316 GND.n1830 GND.t0 8.0712
R8317 GND.n3195 GND.t88 8.0712
R8318 GND.n2955 GND.t63 7.70435
R8319 GND.n3135 GND.t56 7.70435
R8320 GND.n2974 GND.n2973 7.3375
R8321 GND.n3670 GND.n1708 7.3375
R8322 GND.n3622 GND.n1768 7.3375
R8323 GND.n3120 GND.n2274 7.3375
R8324 GND.t36 GND.n1872 7.3375
R8325 GND.n3048 GND.t133 6.97065
R8326 GND.n3083 GND.t7 6.97065
R8327 GND.n3706 GND.n1651 6.6038
R8328 GND.n2904 GND.n2903 6.6038
R8329 GND.n3699 GND.t49 6.6038
R8330 GND.n3649 GND.n1735 6.6038
R8331 GND.n3643 GND.n1741 6.6038
R8332 GND.t85 GND.n1820 6.6038
R8333 GND.n1830 GND.n1822 6.6038
R8334 GND.n208 GND.n205 6.4005
R8335 GND.n2656 GND.n2569 6.4005
R8336 GND.n3520 GND.n1933 6.20656
R8337 GND.n3865 GND.n3864 6.20656
R8338 GND.n2848 GND.n2847 6.01262
R8339 GND.n3319 GND.n3279 6.01262
R8340 GND.n3233 GND.n3231 6.01262
R8341 GND.n2756 GND.n2526 6.01262
R8342 GND.t9 GND.n1641 5.8701
R8343 GND.n3705 GND.t122 5.8701
R8344 GND.n3678 GND.n3677 5.8701
R8345 GND.n2980 GND.n2979 5.8701
R8346 GND.n2991 GND.n2990 5.8701
R8347 GND.n3615 GND.n3614 5.8701
R8348 GND.n3134 GND.t43 5.8701
R8349 GND.n3790 GND.n1605 5.50325
R8350 GND.n2102 GND.n2009 5.50325
R8351 GND.n2102 GND.t36 5.50325
R8352 GND.t70 GND.n2911 5.1364
R8353 GND.n2951 GND.n2950 5.1364
R8354 GND.n2965 GND.t23 5.1364
R8355 GND.t136 GND.n1684 5.1364
R8356 GND.n3062 GND.n1733 5.1364
R8357 GND.n2303 GND.n1743 5.1364
R8358 GND.t134 GND.n1786 5.1364
R8359 GND.n3130 GND.n1806 5.1364
R8360 GND.n3581 GND.n1829 5.1364
R8361 GND.n3181 GND.t92 5.1364
R8362 GND.n3994 GND.n1348 4.76955
R8363 GND.n5467 GND.n258 4.76955
R8364 GND.n2168 GND.n24 4.74817
R8365 GND.n22 GND.n16 4.74817
R8366 GND.n5497 GND.n17 4.74817
R8367 GND.n25 GND.n21 4.74817
R8368 GND.n3379 GND.n24 4.74817
R8369 GND.n2187 GND.n22 4.74817
R8370 GND.n5498 GND.n5497 4.74817
R8371 GND.n2231 GND.n21 4.74817
R8372 GND.n2513 GND.n2512 4.74817
R8373 GND.n2510 GND.n2451 4.74817
R8374 GND.n2503 GND.n2450 4.74817
R8375 GND.n2499 GND.n2449 4.74817
R8376 GND.n2495 GND.n2448 4.74817
R8377 GND.n2218 GND.n2217 4.74817
R8378 GND.n3373 GND.n3372 4.74817
R8379 GND.n3341 GND.n2219 4.74817
R8380 GND.n3358 GND.n3357 4.74817
R8381 GND.n3353 GND.n3342 4.74817
R8382 GND.n2217 GND.n2216 4.74817
R8383 GND.n3374 GND.n3373 4.74817
R8384 GND.n3371 GND.n2219 4.74817
R8385 GND.n3359 GND.n3358 4.74817
R8386 GND.n3356 GND.n3342 4.74817
R8387 GND.n2779 GND.n2778 4.74817
R8388 GND.n2781 GND.n2408 4.74817
R8389 GND.n2805 GND.n2804 4.74817
R8390 GND.n2807 GND.n2806 4.74817
R8391 GND.n2780 GND.n2779 4.74817
R8392 GND.n2782 GND.n2781 4.74817
R8393 GND.n2804 GND.n2803 4.74817
R8394 GND.n2808 GND.n2807 4.74817
R8395 GND.n2512 GND.n2446 4.74817
R8396 GND.n2510 GND.n2509 4.74817
R8397 GND.n2505 GND.n2450 4.74817
R8398 GND.n2502 GND.n2449 4.74817
R8399 GND.n2498 GND.n2448 4.74817
R8400 GND.n5509 GND.n5504 4.62047
R8401 GND.n2791 GND.n4 4.62047
R8402 GND.n3456 GND.n2107 4.6132
R8403 GND.n1470 GND.n1452 4.6132
R8404 GND.n3684 GND.n1684 4.4027
R8405 GND.n3034 GND.n3031 4.4027
R8406 GND.n2284 GND.n2283 4.4027
R8407 GND.n3608 GND.n1786 4.4027
R8408 GND.n3928 GND.n1435 4.07323
R8409 GND.n3477 GND.n1993 4.07323
R8410 GND.n233 GND.n108 4.07323
R8411 GND.n2586 GND.n2581 4.07323
R8412 GND.n3 GND.n2 3.8023
R8413 GND.n5508 GND.n5507 3.8023
R8414 GND.n3988 GND.n3987 3.669
R8415 GND.n2761 GND.n1359 3.669
R8416 GND.n3981 GND.n1368 3.669
R8417 GND.n2518 GND.n2517 3.669
R8418 GND.n2771 GND.n2437 3.669
R8419 GND.n2776 GND.n2433 3.669
R8420 GND.n2773 GND.n2436 3.669
R8421 GND.n2785 GND.n2422 3.669
R8422 GND.n2427 GND.n2423 3.669
R8423 GND.n2795 GND.n2414 3.669
R8424 GND.n2801 GND.n2410 3.669
R8425 GND.n2798 GND.n2412 3.669
R8426 GND.n2810 GND.n2401 3.669
R8427 GND.n2406 GND.n2402 3.669
R8428 GND.n2824 GND.n2394 3.669
R8429 GND.n2828 GND.n2390 3.669
R8430 GND.n2816 GND.n2392 3.669
R8431 GND.n2836 GND.n2383 3.669
R8432 GND.n2839 GND.n2381 3.669
R8433 GND.n3950 GND.n1411 3.669
R8434 GND.n2898 GND.t3 3.669
R8435 GND.n3657 GND.n1723 3.669
R8436 GND.n3635 GND.n1753 3.669
R8437 GND.n3601 GND.n3600 3.669
R8438 GND.n3401 GND.n2148 3.669
R8439 GND.n2246 GND.n2156 3.669
R8440 GND.n3393 GND.n2158 3.669
R8441 GND.n3239 GND.n2170 3.669
R8442 GND.n3387 GND.n2173 3.669
R8443 GND.n3254 GND.n2183 3.669
R8444 GND.n3381 GND.n2186 3.669
R8445 GND.n3377 GND.n3376 3.669
R8446 GND.n2221 GND.n2191 3.669
R8447 GND.n3369 GND.n3368 3.669
R8448 GND.n5500 GND.n12 3.669
R8449 GND.n3362 GND.n3361 3.669
R8450 GND.n3339 GND.n2233 3.669
R8451 GND.n3338 GND.n29 3.669
R8452 GND.n5493 GND.n32 3.669
R8453 GND.n3332 GND.n41 3.669
R8454 GND.n5487 GND.n44 3.669
R8455 GND.n3326 GND.n51 3.669
R8456 GND.n5481 GND.n54 3.669
R8457 GND.n5474 GND.n5473 3.669
R8458 GND.n4 GND.n3 3.13796
R8459 GND.n5509 GND.n5508 3.13796
R8460 GND.n3692 GND.t107 2.9353
R8461 GND.n2341 GND.n1673 2.9353
R8462 GND.n2318 GND.n2317 2.9353
R8463 GND.t4 GND.n1723 2.9353
R8464 GND.t5 GND.n1753 2.9353
R8465 GND.n2293 GND.n2292 2.9353
R8466 GND.n3141 GND.t104 2.9353
R8467 GND.t0 GND.t67 2.9353
R8468 GND.n3575 GND.t92 2.9353
R8469 GND.n1 GND.n0 2.71602
R8470 GND.n2 GND.n1 2.71602
R8471 GND.n5506 GND.n5505 2.71602
R8472 GND.n5507 GND.n5506 2.71602
R8473 GND.n2484 GND.n1467 2.56845
R8474 GND.t63 GND.n1670 2.56845
R8475 GND.n3663 GND.t133 2.56845
R8476 GND.n3629 GND.t7 2.56845
R8477 GND.t56 GND.n1799 2.56845
R8478 GND.n3500 GND.n1976 2.56845
R8479 GND.n3931 GND.n1435 2.52171
R8480 GND.n3480 GND.n1993 2.52171
R8481 GND.n236 GND.n108 2.52171
R8482 GND.n2621 GND.n2586 2.52171
R8483 GND GND.n4 2.36659
R8484 GND.n5496 GND.n24 2.27742
R8485 GND.n5496 GND.n22 2.27742
R8486 GND.n5497 GND.n5496 2.27742
R8487 GND.n5496 GND.n21 2.27742
R8488 GND.n2217 GND.n20 2.27742
R8489 GND.n3373 GND.n20 2.27742
R8490 GND.n2219 GND.n20 2.27742
R8491 GND.n3358 GND.n20 2.27742
R8492 GND.n3342 GND.n20 2.27742
R8493 GND.n2779 GND.n2387 2.27742
R8494 GND.n2781 GND.n2387 2.27742
R8495 GND.n2804 GND.n2387 2.27742
R8496 GND.n2807 GND.n2387 2.27742
R8497 GND.n2512 GND.n2511 2.27742
R8498 GND.n2511 GND.n2510 2.27742
R8499 GND.n2511 GND.n2450 2.27742
R8500 GND.n2511 GND.n2449 2.27742
R8501 GND.n2511 GND.n2448 2.27742
R8502 GND.n3850 GND.n1551 2.2016
R8503 GND.n3685 GND.n1682 2.2016
R8504 GND.n3030 GND.n1716 2.2016
R8505 GND.n2285 GND.n1760 2.2016
R8506 GND.n3607 GND.n1788 2.2016
R8507 GND.n3545 GND.n1907 2.2016
R8508 GND GND.n5509 2.19715
R8509 GND.n1629 GND.n1611 2.19141
R8510 GND.n1624 GND.n1623 2.19141
R8511 GND.n1842 GND.n1837 2.19141
R8512 GND.n1844 GND.n1835 2.19141
R8513 GND.n1852 GND.n1834 1.55202
R8514 GND.n2892 GND.n1643 1.4679
R8515 GND.n3699 GND.n3698 1.4679
R8516 GND.n3019 GND.n2310 1.4679
R8517 GND.n2302 GND.n2301 1.4679
R8518 GND.n3594 GND.n3593 1.4679
R8519 GND.n3160 GND.n3159 1.4679
R8520 GND.n2026 GND.n2021 1.24928
R8521 GND.n3744 GND.n3743 1.24928
R8522 GND.n3762 GND.n3761 1.24928
R8523 GND.n2077 GND.n2076 1.24928
R8524 GND.n3908 GND.n1452 0.776258
R8525 GND.n3456 GND.n3455 0.776258
R8526 GND.t107 GND.n3691 0.7342
R8527 GND.n2975 GND.n1698 0.7342
R8528 GND.n3671 GND.n1706 0.7342
R8529 GND.n3621 GND.n1770 0.7342
R8530 GND.n2273 GND.n1778 0.7342
R8531 GND.t67 GND.n1828 0.7342
R8532 GND.n2849 GND.n2848 0.582318
R8533 GND.n3315 GND.n3279 0.582318
R8534 GND.n3231 GND.n3230 0.582318
R8535 GND.n2527 GND.n2526 0.582318
R8536 GND.n3321 GND.n3320 0.544707
R8537 GND.n2758 GND.n2757 0.544707
R8538 GND.n97 GND.n96 0.529463
R8539 GND.n2164 GND.n1980 0.529463
R8540 GND.n3947 GND.n3946 0.529463
R8541 GND.n2594 GND.n1363 0.529463
R8542 GND.n3811 GND.n3810 0.456293
R8543 GND.n3549 GND.n3548 0.456293
R8544 GND.n1031 GND.n1026 0.445622
R8545 GND.n5120 GND.n547 0.445622
R8546 GND.n5253 GND.n464 0.445622
R8547 GND.n1143 GND.n1142 0.445622
R8548 GND.n3517 GND.n1933 0.388379
R8549 GND.n3864 GND.n3861 0.388379
R8550 GND.n5496 GND.n20 0.388125
R8551 GND.n2511 GND.n2387 0.388125
R8552 GND.n3235 GND.n3234 0.370491
R8553 GND.n2844 GND.n2843 0.370491
R8554 GND.n2105 GND.n2005 0.312695
R8555 GND.n3753 GND.n3751 0.312695
R8556 GND.n3754 GND.n3753 0.312695
R8557 GND.n2105 GND.n2006 0.312695
R8558 GND.n3291 GND.n57 0.306902
R8559 GND.n2729 GND.n2728 0.306902
R8560 GND.n152 GND.n57 0.291659
R8561 GND.n3405 GND.n2143 0.291659
R8562 GND.n2728 GND.n2724 0.291659
R8563 GND.n3869 GND.n3868 0.291659
R8564 GND.n2107 GND.n2004 0.229039
R8565 GND.n2110 GND.n2107 0.229039
R8566 GND.n1470 GND.n1449 0.229039
R8567 GND.n3907 GND.n1470 0.229039
R8568 GND.n209 GND.n208 0.194439
R8569 GND.n2653 GND.n2569 0.194439
R8570 GND.n2859 GND.n2858 0.175805
R8571 GND.n3215 GND.n3201 0.175805
R8572 GND.n4319 GND.n1026 0.152939
R8573 GND.n4320 GND.n4319 0.152939
R8574 GND.n4321 GND.n4320 0.152939
R8575 GND.n4321 GND.n1020 0.152939
R8576 GND.n4329 GND.n1020 0.152939
R8577 GND.n4330 GND.n4329 0.152939
R8578 GND.n4331 GND.n4330 0.152939
R8579 GND.n4331 GND.n1014 0.152939
R8580 GND.n4339 GND.n1014 0.152939
R8581 GND.n4340 GND.n4339 0.152939
R8582 GND.n4341 GND.n4340 0.152939
R8583 GND.n4341 GND.n1008 0.152939
R8584 GND.n4349 GND.n1008 0.152939
R8585 GND.n4350 GND.n4349 0.152939
R8586 GND.n4351 GND.n4350 0.152939
R8587 GND.n4351 GND.n1002 0.152939
R8588 GND.n4359 GND.n1002 0.152939
R8589 GND.n4360 GND.n4359 0.152939
R8590 GND.n4361 GND.n4360 0.152939
R8591 GND.n4361 GND.n996 0.152939
R8592 GND.n4369 GND.n996 0.152939
R8593 GND.n4370 GND.n4369 0.152939
R8594 GND.n4371 GND.n4370 0.152939
R8595 GND.n4371 GND.n990 0.152939
R8596 GND.n4379 GND.n990 0.152939
R8597 GND.n4380 GND.n4379 0.152939
R8598 GND.n4381 GND.n4380 0.152939
R8599 GND.n4381 GND.n984 0.152939
R8600 GND.n4389 GND.n984 0.152939
R8601 GND.n4390 GND.n4389 0.152939
R8602 GND.n4391 GND.n4390 0.152939
R8603 GND.n4391 GND.n978 0.152939
R8604 GND.n4399 GND.n978 0.152939
R8605 GND.n4400 GND.n4399 0.152939
R8606 GND.n4401 GND.n4400 0.152939
R8607 GND.n4401 GND.n972 0.152939
R8608 GND.n4409 GND.n972 0.152939
R8609 GND.n4410 GND.n4409 0.152939
R8610 GND.n4411 GND.n4410 0.152939
R8611 GND.n4411 GND.n966 0.152939
R8612 GND.n4419 GND.n966 0.152939
R8613 GND.n4420 GND.n4419 0.152939
R8614 GND.n4421 GND.n4420 0.152939
R8615 GND.n4421 GND.n960 0.152939
R8616 GND.n4429 GND.n960 0.152939
R8617 GND.n4430 GND.n4429 0.152939
R8618 GND.n4431 GND.n4430 0.152939
R8619 GND.n4431 GND.n954 0.152939
R8620 GND.n4439 GND.n954 0.152939
R8621 GND.n4440 GND.n4439 0.152939
R8622 GND.n4441 GND.n4440 0.152939
R8623 GND.n4441 GND.n948 0.152939
R8624 GND.n4449 GND.n948 0.152939
R8625 GND.n4450 GND.n4449 0.152939
R8626 GND.n4451 GND.n4450 0.152939
R8627 GND.n4451 GND.n942 0.152939
R8628 GND.n4459 GND.n942 0.152939
R8629 GND.n4460 GND.n4459 0.152939
R8630 GND.n4461 GND.n4460 0.152939
R8631 GND.n4461 GND.n936 0.152939
R8632 GND.n4469 GND.n936 0.152939
R8633 GND.n4470 GND.n4469 0.152939
R8634 GND.n4471 GND.n4470 0.152939
R8635 GND.n4471 GND.n930 0.152939
R8636 GND.n4479 GND.n930 0.152939
R8637 GND.n4480 GND.n4479 0.152939
R8638 GND.n4481 GND.n4480 0.152939
R8639 GND.n4481 GND.n924 0.152939
R8640 GND.n4489 GND.n924 0.152939
R8641 GND.n4490 GND.n4489 0.152939
R8642 GND.n4491 GND.n4490 0.152939
R8643 GND.n4491 GND.n918 0.152939
R8644 GND.n4499 GND.n918 0.152939
R8645 GND.n4500 GND.n4499 0.152939
R8646 GND.n4501 GND.n4500 0.152939
R8647 GND.n4501 GND.n912 0.152939
R8648 GND.n4509 GND.n912 0.152939
R8649 GND.n4510 GND.n4509 0.152939
R8650 GND.n4511 GND.n4510 0.152939
R8651 GND.n4511 GND.n906 0.152939
R8652 GND.n4519 GND.n906 0.152939
R8653 GND.n4520 GND.n4519 0.152939
R8654 GND.n4521 GND.n4520 0.152939
R8655 GND.n4521 GND.n900 0.152939
R8656 GND.n4529 GND.n900 0.152939
R8657 GND.n4530 GND.n4529 0.152939
R8658 GND.n4531 GND.n4530 0.152939
R8659 GND.n4531 GND.n894 0.152939
R8660 GND.n4539 GND.n894 0.152939
R8661 GND.n4540 GND.n4539 0.152939
R8662 GND.n4541 GND.n4540 0.152939
R8663 GND.n4541 GND.n888 0.152939
R8664 GND.n4549 GND.n888 0.152939
R8665 GND.n4550 GND.n4549 0.152939
R8666 GND.n4551 GND.n4550 0.152939
R8667 GND.n4551 GND.n882 0.152939
R8668 GND.n4559 GND.n882 0.152939
R8669 GND.n4560 GND.n4559 0.152939
R8670 GND.n4561 GND.n4560 0.152939
R8671 GND.n4561 GND.n876 0.152939
R8672 GND.n4569 GND.n876 0.152939
R8673 GND.n4570 GND.n4569 0.152939
R8674 GND.n4571 GND.n4570 0.152939
R8675 GND.n4571 GND.n870 0.152939
R8676 GND.n4579 GND.n870 0.152939
R8677 GND.n4580 GND.n4579 0.152939
R8678 GND.n4581 GND.n4580 0.152939
R8679 GND.n4581 GND.n864 0.152939
R8680 GND.n4589 GND.n864 0.152939
R8681 GND.n4590 GND.n4589 0.152939
R8682 GND.n4591 GND.n4590 0.152939
R8683 GND.n4591 GND.n858 0.152939
R8684 GND.n4599 GND.n858 0.152939
R8685 GND.n4600 GND.n4599 0.152939
R8686 GND.n4601 GND.n4600 0.152939
R8687 GND.n4601 GND.n852 0.152939
R8688 GND.n4609 GND.n852 0.152939
R8689 GND.n4610 GND.n4609 0.152939
R8690 GND.n4611 GND.n4610 0.152939
R8691 GND.n4611 GND.n846 0.152939
R8692 GND.n4619 GND.n846 0.152939
R8693 GND.n4620 GND.n4619 0.152939
R8694 GND.n4621 GND.n4620 0.152939
R8695 GND.n4621 GND.n840 0.152939
R8696 GND.n4629 GND.n840 0.152939
R8697 GND.n4630 GND.n4629 0.152939
R8698 GND.n4631 GND.n4630 0.152939
R8699 GND.n4631 GND.n834 0.152939
R8700 GND.n4639 GND.n834 0.152939
R8701 GND.n4640 GND.n4639 0.152939
R8702 GND.n4641 GND.n4640 0.152939
R8703 GND.n4641 GND.n828 0.152939
R8704 GND.n4649 GND.n828 0.152939
R8705 GND.n4650 GND.n4649 0.152939
R8706 GND.n4651 GND.n4650 0.152939
R8707 GND.n4651 GND.n822 0.152939
R8708 GND.n4659 GND.n822 0.152939
R8709 GND.n4660 GND.n4659 0.152939
R8710 GND.n4661 GND.n4660 0.152939
R8711 GND.n4661 GND.n816 0.152939
R8712 GND.n4669 GND.n816 0.152939
R8713 GND.n4670 GND.n4669 0.152939
R8714 GND.n4671 GND.n4670 0.152939
R8715 GND.n4671 GND.n810 0.152939
R8716 GND.n4679 GND.n810 0.152939
R8717 GND.n4680 GND.n4679 0.152939
R8718 GND.n4681 GND.n4680 0.152939
R8719 GND.n4681 GND.n804 0.152939
R8720 GND.n4689 GND.n804 0.152939
R8721 GND.n4690 GND.n4689 0.152939
R8722 GND.n4691 GND.n4690 0.152939
R8723 GND.n4691 GND.n798 0.152939
R8724 GND.n4699 GND.n798 0.152939
R8725 GND.n4700 GND.n4699 0.152939
R8726 GND.n4701 GND.n4700 0.152939
R8727 GND.n4701 GND.n792 0.152939
R8728 GND.n4709 GND.n792 0.152939
R8729 GND.n4710 GND.n4709 0.152939
R8730 GND.n4711 GND.n4710 0.152939
R8731 GND.n4711 GND.n786 0.152939
R8732 GND.n4719 GND.n786 0.152939
R8733 GND.n4720 GND.n4719 0.152939
R8734 GND.n4721 GND.n4720 0.152939
R8735 GND.n4721 GND.n780 0.152939
R8736 GND.n4729 GND.n780 0.152939
R8737 GND.n4730 GND.n4729 0.152939
R8738 GND.n4731 GND.n4730 0.152939
R8739 GND.n4731 GND.n774 0.152939
R8740 GND.n4739 GND.n774 0.152939
R8741 GND.n4740 GND.n4739 0.152939
R8742 GND.n4741 GND.n4740 0.152939
R8743 GND.n4741 GND.n768 0.152939
R8744 GND.n4749 GND.n768 0.152939
R8745 GND.n4750 GND.n4749 0.152939
R8746 GND.n4751 GND.n4750 0.152939
R8747 GND.n4751 GND.n762 0.152939
R8748 GND.n4759 GND.n762 0.152939
R8749 GND.n4760 GND.n4759 0.152939
R8750 GND.n4761 GND.n4760 0.152939
R8751 GND.n4761 GND.n756 0.152939
R8752 GND.n4769 GND.n756 0.152939
R8753 GND.n4770 GND.n4769 0.152939
R8754 GND.n4771 GND.n4770 0.152939
R8755 GND.n4771 GND.n750 0.152939
R8756 GND.n4779 GND.n750 0.152939
R8757 GND.n4780 GND.n4779 0.152939
R8758 GND.n4781 GND.n4780 0.152939
R8759 GND.n4781 GND.n744 0.152939
R8760 GND.n4789 GND.n744 0.152939
R8761 GND.n4790 GND.n4789 0.152939
R8762 GND.n4791 GND.n4790 0.152939
R8763 GND.n4791 GND.n738 0.152939
R8764 GND.n4799 GND.n738 0.152939
R8765 GND.n4800 GND.n4799 0.152939
R8766 GND.n4801 GND.n4800 0.152939
R8767 GND.n4801 GND.n732 0.152939
R8768 GND.n4809 GND.n732 0.152939
R8769 GND.n4810 GND.n4809 0.152939
R8770 GND.n4811 GND.n4810 0.152939
R8771 GND.n4811 GND.n726 0.152939
R8772 GND.n4819 GND.n726 0.152939
R8773 GND.n4820 GND.n4819 0.152939
R8774 GND.n4821 GND.n4820 0.152939
R8775 GND.n4821 GND.n720 0.152939
R8776 GND.n4829 GND.n720 0.152939
R8777 GND.n4830 GND.n4829 0.152939
R8778 GND.n4831 GND.n4830 0.152939
R8779 GND.n4831 GND.n714 0.152939
R8780 GND.n4839 GND.n714 0.152939
R8781 GND.n4840 GND.n4839 0.152939
R8782 GND.n4841 GND.n4840 0.152939
R8783 GND.n4841 GND.n708 0.152939
R8784 GND.n4849 GND.n708 0.152939
R8785 GND.n4850 GND.n4849 0.152939
R8786 GND.n4851 GND.n4850 0.152939
R8787 GND.n4851 GND.n702 0.152939
R8788 GND.n4859 GND.n702 0.152939
R8789 GND.n4860 GND.n4859 0.152939
R8790 GND.n4861 GND.n4860 0.152939
R8791 GND.n4861 GND.n696 0.152939
R8792 GND.n4869 GND.n696 0.152939
R8793 GND.n4870 GND.n4869 0.152939
R8794 GND.n4871 GND.n4870 0.152939
R8795 GND.n4871 GND.n690 0.152939
R8796 GND.n4879 GND.n690 0.152939
R8797 GND.n4880 GND.n4879 0.152939
R8798 GND.n4881 GND.n4880 0.152939
R8799 GND.n4881 GND.n684 0.152939
R8800 GND.n4889 GND.n684 0.152939
R8801 GND.n4890 GND.n4889 0.152939
R8802 GND.n4891 GND.n4890 0.152939
R8803 GND.n4891 GND.n678 0.152939
R8804 GND.n4899 GND.n678 0.152939
R8805 GND.n4900 GND.n4899 0.152939
R8806 GND.n4901 GND.n4900 0.152939
R8807 GND.n4901 GND.n672 0.152939
R8808 GND.n4909 GND.n672 0.152939
R8809 GND.n4910 GND.n4909 0.152939
R8810 GND.n4911 GND.n4910 0.152939
R8811 GND.n4911 GND.n666 0.152939
R8812 GND.n4919 GND.n666 0.152939
R8813 GND.n4920 GND.n4919 0.152939
R8814 GND.n4921 GND.n4920 0.152939
R8815 GND.n4921 GND.n660 0.152939
R8816 GND.n4929 GND.n660 0.152939
R8817 GND.n4930 GND.n4929 0.152939
R8818 GND.n4931 GND.n4930 0.152939
R8819 GND.n4931 GND.n654 0.152939
R8820 GND.n4939 GND.n654 0.152939
R8821 GND.n4940 GND.n4939 0.152939
R8822 GND.n4941 GND.n4940 0.152939
R8823 GND.n4941 GND.n648 0.152939
R8824 GND.n4949 GND.n648 0.152939
R8825 GND.n4950 GND.n4949 0.152939
R8826 GND.n4951 GND.n4950 0.152939
R8827 GND.n4951 GND.n642 0.152939
R8828 GND.n4959 GND.n642 0.152939
R8829 GND.n4960 GND.n4959 0.152939
R8830 GND.n4961 GND.n4960 0.152939
R8831 GND.n4961 GND.n636 0.152939
R8832 GND.n4969 GND.n636 0.152939
R8833 GND.n4970 GND.n4969 0.152939
R8834 GND.n4971 GND.n4970 0.152939
R8835 GND.n4971 GND.n630 0.152939
R8836 GND.n4979 GND.n630 0.152939
R8837 GND.n4980 GND.n4979 0.152939
R8838 GND.n4981 GND.n4980 0.152939
R8839 GND.n4981 GND.n624 0.152939
R8840 GND.n4989 GND.n624 0.152939
R8841 GND.n4990 GND.n4989 0.152939
R8842 GND.n4991 GND.n4990 0.152939
R8843 GND.n4991 GND.n618 0.152939
R8844 GND.n4999 GND.n618 0.152939
R8845 GND.n5000 GND.n4999 0.152939
R8846 GND.n5001 GND.n5000 0.152939
R8847 GND.n5001 GND.n612 0.152939
R8848 GND.n5009 GND.n612 0.152939
R8849 GND.n5010 GND.n5009 0.152939
R8850 GND.n5011 GND.n5010 0.152939
R8851 GND.n5011 GND.n606 0.152939
R8852 GND.n5019 GND.n606 0.152939
R8853 GND.n5020 GND.n5019 0.152939
R8854 GND.n5021 GND.n5020 0.152939
R8855 GND.n5021 GND.n600 0.152939
R8856 GND.n5029 GND.n600 0.152939
R8857 GND.n5030 GND.n5029 0.152939
R8858 GND.n5031 GND.n5030 0.152939
R8859 GND.n5031 GND.n594 0.152939
R8860 GND.n5039 GND.n594 0.152939
R8861 GND.n5040 GND.n5039 0.152939
R8862 GND.n5041 GND.n5040 0.152939
R8863 GND.n5041 GND.n588 0.152939
R8864 GND.n5049 GND.n588 0.152939
R8865 GND.n5050 GND.n5049 0.152939
R8866 GND.n5051 GND.n5050 0.152939
R8867 GND.n5051 GND.n582 0.152939
R8868 GND.n5059 GND.n582 0.152939
R8869 GND.n5060 GND.n5059 0.152939
R8870 GND.n5061 GND.n5060 0.152939
R8871 GND.n5061 GND.n576 0.152939
R8872 GND.n5069 GND.n576 0.152939
R8873 GND.n5070 GND.n5069 0.152939
R8874 GND.n5071 GND.n5070 0.152939
R8875 GND.n5071 GND.n570 0.152939
R8876 GND.n5079 GND.n570 0.152939
R8877 GND.n5080 GND.n5079 0.152939
R8878 GND.n5081 GND.n5080 0.152939
R8879 GND.n5081 GND.n564 0.152939
R8880 GND.n5089 GND.n564 0.152939
R8881 GND.n5090 GND.n5089 0.152939
R8882 GND.n5091 GND.n5090 0.152939
R8883 GND.n5091 GND.n558 0.152939
R8884 GND.n5099 GND.n558 0.152939
R8885 GND.n5100 GND.n5099 0.152939
R8886 GND.n5101 GND.n5100 0.152939
R8887 GND.n5101 GND.n552 0.152939
R8888 GND.n5109 GND.n552 0.152939
R8889 GND.n5110 GND.n5109 0.152939
R8890 GND.n5111 GND.n5110 0.152939
R8891 GND.n5111 GND.n547 0.152939
R8892 GND.n5121 GND.n5120 0.152939
R8893 GND.n5122 GND.n5121 0.152939
R8894 GND.n5122 GND.n541 0.152939
R8895 GND.n5130 GND.n541 0.152939
R8896 GND.n5131 GND.n5130 0.152939
R8897 GND.n5132 GND.n5131 0.152939
R8898 GND.n5132 GND.n535 0.152939
R8899 GND.n5140 GND.n535 0.152939
R8900 GND.n5141 GND.n5140 0.152939
R8901 GND.n5142 GND.n5141 0.152939
R8902 GND.n5142 GND.n529 0.152939
R8903 GND.n5150 GND.n529 0.152939
R8904 GND.n5151 GND.n5150 0.152939
R8905 GND.n5152 GND.n5151 0.152939
R8906 GND.n5152 GND.n523 0.152939
R8907 GND.n5160 GND.n523 0.152939
R8908 GND.n5161 GND.n5160 0.152939
R8909 GND.n5162 GND.n5161 0.152939
R8910 GND.n5162 GND.n517 0.152939
R8911 GND.n5170 GND.n517 0.152939
R8912 GND.n5171 GND.n5170 0.152939
R8913 GND.n5172 GND.n5171 0.152939
R8914 GND.n5172 GND.n511 0.152939
R8915 GND.n5180 GND.n511 0.152939
R8916 GND.n5181 GND.n5180 0.152939
R8917 GND.n5182 GND.n5181 0.152939
R8918 GND.n5182 GND.n505 0.152939
R8919 GND.n5190 GND.n505 0.152939
R8920 GND.n5191 GND.n5190 0.152939
R8921 GND.n5192 GND.n5191 0.152939
R8922 GND.n5192 GND.n499 0.152939
R8923 GND.n5200 GND.n499 0.152939
R8924 GND.n5201 GND.n5200 0.152939
R8925 GND.n5202 GND.n5201 0.152939
R8926 GND.n5202 GND.n493 0.152939
R8927 GND.n5210 GND.n493 0.152939
R8928 GND.n5211 GND.n5210 0.152939
R8929 GND.n5212 GND.n5211 0.152939
R8930 GND.n5212 GND.n487 0.152939
R8931 GND.n5220 GND.n487 0.152939
R8932 GND.n5221 GND.n5220 0.152939
R8933 GND.n5222 GND.n5221 0.152939
R8934 GND.n5222 GND.n481 0.152939
R8935 GND.n5230 GND.n481 0.152939
R8936 GND.n5231 GND.n5230 0.152939
R8937 GND.n5232 GND.n5231 0.152939
R8938 GND.n5232 GND.n475 0.152939
R8939 GND.n5240 GND.n475 0.152939
R8940 GND.n5241 GND.n5240 0.152939
R8941 GND.n5242 GND.n5241 0.152939
R8942 GND.n5242 GND.n469 0.152939
R8943 GND.n5250 GND.n469 0.152939
R8944 GND.n5251 GND.n5250 0.152939
R8945 GND.n5252 GND.n5251 0.152939
R8946 GND.n5253 GND.n5252 0.152939
R8947 GND.n3345 GND.n3344 0.152939
R8948 GND.n3347 GND.n3345 0.152939
R8949 GND.n3347 GND.n3346 0.152939
R8950 GND.n3346 GND.n65 0.152939
R8951 GND.n66 GND.n65 0.152939
R8952 GND.n67 GND.n66 0.152939
R8953 GND.n261 GND.n67 0.152939
R8954 GND.n262 GND.n261 0.152939
R8955 GND.n263 GND.n262 0.152939
R8956 GND.n264 GND.n263 0.152939
R8957 GND.n269 GND.n264 0.152939
R8958 GND.n270 GND.n269 0.152939
R8959 GND.n271 GND.n270 0.152939
R8960 GND.n272 GND.n271 0.152939
R8961 GND.n277 GND.n272 0.152939
R8962 GND.n278 GND.n277 0.152939
R8963 GND.n279 GND.n278 0.152939
R8964 GND.n280 GND.n279 0.152939
R8965 GND.n285 GND.n280 0.152939
R8966 GND.n286 GND.n285 0.152939
R8967 GND.n287 GND.n286 0.152939
R8968 GND.n288 GND.n287 0.152939
R8969 GND.n293 GND.n288 0.152939
R8970 GND.n294 GND.n293 0.152939
R8971 GND.n295 GND.n294 0.152939
R8972 GND.n296 GND.n295 0.152939
R8973 GND.n301 GND.n296 0.152939
R8974 GND.n302 GND.n301 0.152939
R8975 GND.n303 GND.n302 0.152939
R8976 GND.n304 GND.n303 0.152939
R8977 GND.n309 GND.n304 0.152939
R8978 GND.n310 GND.n309 0.152939
R8979 GND.n311 GND.n310 0.152939
R8980 GND.n312 GND.n311 0.152939
R8981 GND.n317 GND.n312 0.152939
R8982 GND.n318 GND.n317 0.152939
R8983 GND.n319 GND.n318 0.152939
R8984 GND.n320 GND.n319 0.152939
R8985 GND.n325 GND.n320 0.152939
R8986 GND.n326 GND.n325 0.152939
R8987 GND.n327 GND.n326 0.152939
R8988 GND.n328 GND.n327 0.152939
R8989 GND.n333 GND.n328 0.152939
R8990 GND.n334 GND.n333 0.152939
R8991 GND.n335 GND.n334 0.152939
R8992 GND.n336 GND.n335 0.152939
R8993 GND.n341 GND.n336 0.152939
R8994 GND.n342 GND.n341 0.152939
R8995 GND.n343 GND.n342 0.152939
R8996 GND.n344 GND.n343 0.152939
R8997 GND.n349 GND.n344 0.152939
R8998 GND.n350 GND.n349 0.152939
R8999 GND.n351 GND.n350 0.152939
R9000 GND.n352 GND.n351 0.152939
R9001 GND.n357 GND.n352 0.152939
R9002 GND.n358 GND.n357 0.152939
R9003 GND.n359 GND.n358 0.152939
R9004 GND.n360 GND.n359 0.152939
R9005 GND.n365 GND.n360 0.152939
R9006 GND.n366 GND.n365 0.152939
R9007 GND.n367 GND.n366 0.152939
R9008 GND.n368 GND.n367 0.152939
R9009 GND.n373 GND.n368 0.152939
R9010 GND.n374 GND.n373 0.152939
R9011 GND.n375 GND.n374 0.152939
R9012 GND.n376 GND.n375 0.152939
R9013 GND.n381 GND.n376 0.152939
R9014 GND.n382 GND.n381 0.152939
R9015 GND.n383 GND.n382 0.152939
R9016 GND.n384 GND.n383 0.152939
R9017 GND.n389 GND.n384 0.152939
R9018 GND.n390 GND.n389 0.152939
R9019 GND.n391 GND.n390 0.152939
R9020 GND.n392 GND.n391 0.152939
R9021 GND.n397 GND.n392 0.152939
R9022 GND.n398 GND.n397 0.152939
R9023 GND.n399 GND.n398 0.152939
R9024 GND.n400 GND.n399 0.152939
R9025 GND.n405 GND.n400 0.152939
R9026 GND.n406 GND.n405 0.152939
R9027 GND.n407 GND.n406 0.152939
R9028 GND.n408 GND.n407 0.152939
R9029 GND.n413 GND.n408 0.152939
R9030 GND.n414 GND.n413 0.152939
R9031 GND.n415 GND.n414 0.152939
R9032 GND.n416 GND.n415 0.152939
R9033 GND.n421 GND.n416 0.152939
R9034 GND.n422 GND.n421 0.152939
R9035 GND.n423 GND.n422 0.152939
R9036 GND.n424 GND.n423 0.152939
R9037 GND.n429 GND.n424 0.152939
R9038 GND.n430 GND.n429 0.152939
R9039 GND.n431 GND.n430 0.152939
R9040 GND.n432 GND.n431 0.152939
R9041 GND.n437 GND.n432 0.152939
R9042 GND.n438 GND.n437 0.152939
R9043 GND.n439 GND.n438 0.152939
R9044 GND.n440 GND.n439 0.152939
R9045 GND.n445 GND.n440 0.152939
R9046 GND.n446 GND.n445 0.152939
R9047 GND.n447 GND.n446 0.152939
R9048 GND.n448 GND.n447 0.152939
R9049 GND.n453 GND.n448 0.152939
R9050 GND.n454 GND.n453 0.152939
R9051 GND.n455 GND.n454 0.152939
R9052 GND.n456 GND.n455 0.152939
R9053 GND.n461 GND.n456 0.152939
R9054 GND.n462 GND.n461 0.152939
R9055 GND.n463 GND.n462 0.152939
R9056 GND.n464 GND.n463 0.152939
R9057 GND.n46 GND.n18 0.152939
R9058 GND.n47 GND.n46 0.152939
R9059 GND.n48 GND.n47 0.152939
R9060 GND.n96 GND.n48 0.152939
R9061 GND.n2860 GND.n2859 0.152939
R9062 GND.n2860 GND.n2356 0.152939
R9063 GND.n2866 GND.n2356 0.152939
R9064 GND.n2867 GND.n2866 0.152939
R9065 GND.n2868 GND.n2867 0.152939
R9066 GND.n2868 GND.n2354 0.152939
R9067 GND.n2874 GND.n2354 0.152939
R9068 GND.n2875 GND.n2874 0.152939
R9069 GND.n2876 GND.n2875 0.152939
R9070 GND.n2876 GND.n2350 0.152939
R9071 GND.n2915 GND.n2350 0.152939
R9072 GND.n2916 GND.n2915 0.152939
R9073 GND.n2917 GND.n2916 0.152939
R9074 GND.n2918 GND.n2917 0.152939
R9075 GND.n2919 GND.n2918 0.152939
R9076 GND.n2920 GND.n2919 0.152939
R9077 GND.n2921 GND.n2920 0.152939
R9078 GND.n2922 GND.n2921 0.152939
R9079 GND.n2925 GND.n2922 0.152939
R9080 GND.n2926 GND.n2925 0.152939
R9081 GND.n2927 GND.n2926 0.152939
R9082 GND.n2928 GND.n2927 0.152939
R9083 GND.n2929 GND.n2928 0.152939
R9084 GND.n2929 GND.n2314 0.152939
R9085 GND.n3052 GND.n2314 0.152939
R9086 GND.n3053 GND.n3052 0.152939
R9087 GND.n3054 GND.n3053 0.152939
R9088 GND.n3055 GND.n3054 0.152939
R9089 GND.n3056 GND.n3055 0.152939
R9090 GND.n3056 GND.n2296 0.152939
R9091 GND.n3075 GND.n2296 0.152939
R9092 GND.n3076 GND.n3075 0.152939
R9093 GND.n3077 GND.n3076 0.152939
R9094 GND.n3079 GND.n3077 0.152939
R9095 GND.n3079 GND.n3078 0.152939
R9096 GND.n3078 GND.n2277 0.152939
R9097 GND.n3105 GND.n2277 0.152939
R9098 GND.n3106 GND.n3105 0.152939
R9099 GND.n3108 GND.n3106 0.152939
R9100 GND.n3108 GND.n3107 0.152939
R9101 GND.n3107 GND.n2265 0.152939
R9102 GND.n3146 GND.n2265 0.152939
R9103 GND.n3147 GND.n3146 0.152939
R9104 GND.n3148 GND.n3147 0.152939
R9105 GND.n3148 GND.n2261 0.152939
R9106 GND.n3154 GND.n2261 0.152939
R9107 GND.n3155 GND.n3154 0.152939
R9108 GND.n3157 GND.n3155 0.152939
R9109 GND.n3157 GND.n3156 0.152939
R9110 GND.n3156 GND.n2258 0.152939
R9111 GND.n2258 GND.n2256 0.152939
R9112 GND.n3190 GND.n2256 0.152939
R9113 GND.n3191 GND.n3190 0.152939
R9114 GND.n3192 GND.n3191 0.152939
R9115 GND.n3192 GND.n2254 0.152939
R9116 GND.n3200 GND.n2254 0.152939
R9117 GND.n3201 GND.n3200 0.152939
R9118 GND.n3812 GND.n3811 0.152939
R9119 GND.n3813 GND.n3812 0.152939
R9120 GND.n3814 GND.n3813 0.152939
R9121 GND.n3815 GND.n3814 0.152939
R9122 GND.n3816 GND.n3815 0.152939
R9123 GND.n3817 GND.n3816 0.152939
R9124 GND.n3818 GND.n3817 0.152939
R9125 GND.n3819 GND.n3818 0.152939
R9126 GND.n3820 GND.n3819 0.152939
R9127 GND.n3821 GND.n3820 0.152939
R9128 GND.n3822 GND.n3821 0.152939
R9129 GND.n3823 GND.n3822 0.152939
R9130 GND.n3823 GND.n1525 0.152939
R9131 GND.n3810 GND.n1555 0.152939
R9132 GND.n1557 GND.n1555 0.152939
R9133 GND.n1578 GND.n1557 0.152939
R9134 GND.n1579 GND.n1578 0.152939
R9135 GND.n1580 GND.n1579 0.152939
R9136 GND.n1581 GND.n1580 0.152939
R9137 GND.n1582 GND.n1581 0.152939
R9138 GND.n1645 GND.n1582 0.152939
R9139 GND.n1646 GND.n1645 0.152939
R9140 GND.n1647 GND.n1646 0.152939
R9141 GND.n1648 GND.n1647 0.152939
R9142 GND.n2945 GND.n1648 0.152939
R9143 GND.n2947 GND.n2945 0.152939
R9144 GND.n2947 GND.n2946 0.152939
R9145 GND.n2946 GND.n1677 0.152939
R9146 GND.n1678 GND.n1677 0.152939
R9147 GND.n1679 GND.n1678 0.152939
R9148 GND.n2326 GND.n1679 0.152939
R9149 GND.n2327 GND.n2326 0.152939
R9150 GND.n2328 GND.n2327 0.152939
R9151 GND.n2328 GND.n2322 0.152939
R9152 GND.n3038 GND.n2322 0.152939
R9153 GND.n3039 GND.n3038 0.152939
R9154 GND.n3040 GND.n3039 0.152939
R9155 GND.n3041 GND.n3040 0.152939
R9156 GND.n3043 GND.n3041 0.152939
R9157 GND.n3043 GND.n3042 0.152939
R9158 GND.n3042 GND.n2306 0.152939
R9159 GND.n3067 GND.n2306 0.152939
R9160 GND.n3068 GND.n3067 0.152939
R9161 GND.n3069 GND.n3068 0.152939
R9162 GND.n3069 GND.n2289 0.152939
R9163 GND.n3086 GND.n2289 0.152939
R9164 GND.n3087 GND.n3086 0.152939
R9165 GND.n3088 GND.n3087 0.152939
R9166 GND.n3089 GND.n3088 0.152939
R9167 GND.n3090 GND.n3089 0.152939
R9168 GND.n3092 GND.n3090 0.152939
R9169 GND.n3092 GND.n3091 0.152939
R9170 GND.n3091 GND.n1792 0.152939
R9171 GND.n1793 GND.n1792 0.152939
R9172 GND.n1794 GND.n1793 0.152939
R9173 GND.n3166 GND.n1794 0.152939
R9174 GND.n3167 GND.n3166 0.152939
R9175 GND.n3167 GND.n3164 0.152939
R9176 GND.n3173 GND.n3164 0.152939
R9177 GND.n3174 GND.n3173 0.152939
R9178 GND.n3175 GND.n3174 0.152939
R9179 GND.n3177 GND.n3175 0.152939
R9180 GND.n3177 GND.n3176 0.152939
R9181 GND.n3176 GND.n1878 0.152939
R9182 GND.n1879 GND.n1878 0.152939
R9183 GND.n1880 GND.n1879 0.152939
R9184 GND.n1901 GND.n1880 0.152939
R9185 GND.n1902 GND.n1901 0.152939
R9186 GND.n1903 GND.n1902 0.152939
R9187 GND.n3549 GND.n1903 0.152939
R9188 GND.n3548 GND.n1904 0.152939
R9189 GND.n1918 GND.n1904 0.152939
R9190 GND.n1919 GND.n1918 0.152939
R9191 GND.n1920 GND.n1919 0.152939
R9192 GND.n1921 GND.n1920 0.152939
R9193 GND.n1922 GND.n1921 0.152939
R9194 GND.n1923 GND.n1922 0.152939
R9195 GND.n1924 GND.n1923 0.152939
R9196 GND.n1925 GND.n1924 0.152939
R9197 GND.n1926 GND.n1925 0.152939
R9198 GND.n1927 GND.n1926 0.152939
R9199 GND.n1928 GND.n1927 0.152939
R9200 GND.n1929 GND.n1928 0.152939
R9201 GND.n3236 GND.n3235 0.152939
R9202 GND.n3236 GND.n2244 0.152939
R9203 GND.n3242 GND.n2244 0.152939
R9204 GND.n3243 GND.n3242 0.152939
R9205 GND.n3244 GND.n3243 0.152939
R9206 GND.n3245 GND.n3244 0.152939
R9207 GND.n3246 GND.n3245 0.152939
R9208 GND.n3247 GND.n3246 0.152939
R9209 GND.n3247 GND.n5 0.152939
R9210 GND.n5503 GND.n6 0.152939
R9211 GND.n2237 GND.n6 0.152939
R9212 GND.n2238 GND.n2237 0.152939
R9213 GND.n2239 GND.n2238 0.152939
R9214 GND.n2240 GND.n2239 0.152939
R9215 GND.n3273 GND.n2240 0.152939
R9216 GND.n3274 GND.n3273 0.152939
R9217 GND.n3275 GND.n3274 0.152939
R9218 GND.n3321 GND.n3275 0.152939
R9219 GND.n3292 GND.n3291 0.152939
R9220 GND.n3292 GND.n3286 0.152939
R9221 GND.n3300 GND.n3286 0.152939
R9222 GND.n3301 GND.n3300 0.152939
R9223 GND.n3302 GND.n3301 0.152939
R9224 GND.n3302 GND.n3282 0.152939
R9225 GND.n3311 GND.n3282 0.152939
R9226 GND.n3312 GND.n3311 0.152939
R9227 GND.n3313 GND.n3312 0.152939
R9228 GND.n3313 GND.n3276 0.152939
R9229 GND.n3320 GND.n3276 0.152939
R9230 GND.n254 GND.n97 0.152939
R9231 GND.n254 GND.n253 0.152939
R9232 GND.n253 GND.n252 0.152939
R9233 GND.n252 GND.n99 0.152939
R9234 GND.n100 GND.n99 0.152939
R9235 GND.n101 GND.n100 0.152939
R9236 GND.n102 GND.n101 0.152939
R9237 GND.n103 GND.n102 0.152939
R9238 GND.n104 GND.n103 0.152939
R9239 GND.n105 GND.n104 0.152939
R9240 GND.n109 GND.n105 0.152939
R9241 GND.n110 GND.n109 0.152939
R9242 GND.n111 GND.n110 0.152939
R9243 GND.n112 GND.n111 0.152939
R9244 GND.n113 GND.n112 0.152939
R9245 GND.n114 GND.n113 0.152939
R9246 GND.n115 GND.n114 0.152939
R9247 GND.n116 GND.n115 0.152939
R9248 GND.n117 GND.n116 0.152939
R9249 GND.n118 GND.n117 0.152939
R9250 GND.n119 GND.n118 0.152939
R9251 GND.n120 GND.n119 0.152939
R9252 GND.n121 GND.n120 0.152939
R9253 GND.n122 GND.n121 0.152939
R9254 GND.n123 GND.n122 0.152939
R9255 GND.n124 GND.n123 0.152939
R9256 GND.n125 GND.n124 0.152939
R9257 GND.n126 GND.n125 0.152939
R9258 GND.n127 GND.n126 0.152939
R9259 GND.n128 GND.n127 0.152939
R9260 GND.n129 GND.n128 0.152939
R9261 GND.n130 GND.n129 0.152939
R9262 GND.n131 GND.n130 0.152939
R9263 GND.n132 GND.n131 0.152939
R9264 GND.n133 GND.n132 0.152939
R9265 GND.n180 GND.n133 0.152939
R9266 GND.n180 GND.n179 0.152939
R9267 GND.n179 GND.n178 0.152939
R9268 GND.n178 GND.n139 0.152939
R9269 GND.n140 GND.n139 0.152939
R9270 GND.n141 GND.n140 0.152939
R9271 GND.n142 GND.n141 0.152939
R9272 GND.n143 GND.n142 0.152939
R9273 GND.n144 GND.n143 0.152939
R9274 GND.n145 GND.n144 0.152939
R9275 GND.n146 GND.n145 0.152939
R9276 GND.n147 GND.n146 0.152939
R9277 GND.n148 GND.n147 0.152939
R9278 GND.n153 GND.n148 0.152939
R9279 GND.n153 GND.n152 0.152939
R9280 GND.n1981 GND.n1980 0.152939
R9281 GND.n1982 GND.n1981 0.152939
R9282 GND.n1983 GND.n1982 0.152939
R9283 GND.n1984 GND.n1983 0.152939
R9284 GND.n1985 GND.n1984 0.152939
R9285 GND.n1986 GND.n1985 0.152939
R9286 GND.n1987 GND.n1986 0.152939
R9287 GND.n1988 GND.n1987 0.152939
R9288 GND.n1989 GND.n1988 0.152939
R9289 GND.n1990 GND.n1989 0.152939
R9290 GND.n1994 GND.n1990 0.152939
R9291 GND.n1995 GND.n1994 0.152939
R9292 GND.n1996 GND.n1995 0.152939
R9293 GND.n1997 GND.n1996 0.152939
R9294 GND.n1998 GND.n1997 0.152939
R9295 GND.n1999 GND.n1998 0.152939
R9296 GND.n2000 GND.n1999 0.152939
R9297 GND.n2001 GND.n2000 0.152939
R9298 GND.n2002 GND.n2001 0.152939
R9299 GND.n2003 GND.n2002 0.152939
R9300 GND.n2004 GND.n2003 0.152939
R9301 GND.n2111 GND.n2110 0.152939
R9302 GND.n2112 GND.n2111 0.152939
R9303 GND.n2113 GND.n2112 0.152939
R9304 GND.n2114 GND.n2113 0.152939
R9305 GND.n2115 GND.n2114 0.152939
R9306 GND.n2116 GND.n2115 0.152939
R9307 GND.n2117 GND.n2116 0.152939
R9308 GND.n2118 GND.n2117 0.152939
R9309 GND.n2119 GND.n2118 0.152939
R9310 GND.n2120 GND.n2119 0.152939
R9311 GND.n2121 GND.n2120 0.152939
R9312 GND.n2123 GND.n2121 0.152939
R9313 GND.n2126 GND.n2123 0.152939
R9314 GND.n2127 GND.n2126 0.152939
R9315 GND.n2128 GND.n2127 0.152939
R9316 GND.n2129 GND.n2128 0.152939
R9317 GND.n2130 GND.n2129 0.152939
R9318 GND.n2131 GND.n2130 0.152939
R9319 GND.n2132 GND.n2131 0.152939
R9320 GND.n2133 GND.n2132 0.152939
R9321 GND.n2134 GND.n2133 0.152939
R9322 GND.n2135 GND.n2134 0.152939
R9323 GND.n2136 GND.n2135 0.152939
R9324 GND.n3407 GND.n2136 0.152939
R9325 GND.n3407 GND.n3406 0.152939
R9326 GND.n3406 GND.n3405 0.152939
R9327 GND.n2165 GND.n2164 0.152939
R9328 GND.n2166 GND.n2165 0.152939
R9329 GND.n2167 GND.n2166 0.152939
R9330 GND.n2167 GND.n19 0.152939
R9331 GND.n2454 GND.n2447 0.152939
R9332 GND.n2457 GND.n2454 0.152939
R9333 GND.n2458 GND.n2457 0.152939
R9334 GND.n2459 GND.n2458 0.152939
R9335 GND.n2460 GND.n2459 0.152939
R9336 GND.n2463 GND.n2460 0.152939
R9337 GND.n2464 GND.n2463 0.152939
R9338 GND.n2465 GND.n2464 0.152939
R9339 GND.n2466 GND.n2465 0.152939
R9340 GND.n2468 GND.n2466 0.152939
R9341 GND.n2470 GND.n2468 0.152939
R9342 GND.n2470 GND.n2469 0.152939
R9343 GND.n2469 GND.n1566 0.152939
R9344 GND.n1567 GND.n1566 0.152939
R9345 GND.n1568 GND.n1567 0.152939
R9346 GND.n2880 GND.n1568 0.152939
R9347 GND.n2881 GND.n2880 0.152939
R9348 GND.n2886 GND.n2881 0.152939
R9349 GND.n2887 GND.n2886 0.152939
R9350 GND.n2889 GND.n2887 0.152939
R9351 GND.n2889 GND.n2888 0.152939
R9352 GND.n2888 GND.n1658 0.152939
R9353 GND.n1659 GND.n1658 0.152939
R9354 GND.n1660 GND.n1659 0.152939
R9355 GND.n1688 GND.n1660 0.152939
R9356 GND.n1691 GND.n1688 0.152939
R9357 GND.n1692 GND.n1691 0.152939
R9358 GND.n1693 GND.n1692 0.152939
R9359 GND.n1694 GND.n1693 0.152939
R9360 GND.n1695 GND.n1694 0.152939
R9361 GND.n1710 GND.n1695 0.152939
R9362 GND.n1711 GND.n1710 0.152939
R9363 GND.n1712 GND.n1711 0.152939
R9364 GND.n1713 GND.n1712 0.152939
R9365 GND.n1727 GND.n1713 0.152939
R9366 GND.n1728 GND.n1727 0.152939
R9367 GND.n1729 GND.n1728 0.152939
R9368 GND.n1730 GND.n1729 0.152939
R9369 GND.n1745 GND.n1730 0.152939
R9370 GND.n1746 GND.n1745 0.152939
R9371 GND.n1747 GND.n1746 0.152939
R9372 GND.n1748 GND.n1747 0.152939
R9373 GND.n1762 GND.n1748 0.152939
R9374 GND.n1763 GND.n1762 0.152939
R9375 GND.n1764 GND.n1763 0.152939
R9376 GND.n1765 GND.n1764 0.152939
R9377 GND.n1780 GND.n1765 0.152939
R9378 GND.n1781 GND.n1780 0.152939
R9379 GND.n1782 GND.n1781 0.152939
R9380 GND.n1783 GND.n1782 0.152939
R9381 GND.n1810 GND.n1783 0.152939
R9382 GND.n1813 GND.n1810 0.152939
R9383 GND.n1814 GND.n1813 0.152939
R9384 GND.n1815 GND.n1814 0.152939
R9385 GND.n1816 GND.n1815 0.152939
R9386 GND.n1817 GND.n1816 0.152939
R9387 GND.n1865 GND.n1817 0.152939
R9388 GND.n1866 GND.n1865 0.152939
R9389 GND.n1867 GND.n1866 0.152939
R9390 GND.n1868 GND.n1867 0.152939
R9391 GND.n1869 GND.n1868 0.152939
R9392 GND.n1888 GND.n1869 0.152939
R9393 GND.n1889 GND.n1888 0.152939
R9394 GND.n1890 GND.n1889 0.152939
R9395 GND.n1891 GND.n1890 0.152939
R9396 GND.n1892 GND.n1891 0.152939
R9397 GND.n1940 GND.n1892 0.152939
R9398 GND.n1941 GND.n1940 0.152939
R9399 GND.n1942 GND.n1941 0.152939
R9400 GND.n1943 GND.n1942 0.152939
R9401 GND.n2200 GND.n1943 0.152939
R9402 GND.n2201 GND.n2200 0.152939
R9403 GND.n2202 GND.n2201 0.152939
R9404 GND.n2202 GND.n2197 0.152939
R9405 GND.n2208 GND.n2197 0.152939
R9406 GND.n2209 GND.n2208 0.152939
R9407 GND.n2211 GND.n2209 0.152939
R9408 GND.n2211 GND.n2210 0.152939
R9409 GND.n2832 GND.n2831 0.152939
R9410 GND.n2833 GND.n2832 0.152939
R9411 GND.n2833 GND.n1419 0.152939
R9412 GND.n3947 GND.n1419 0.152939
R9413 GND.n2594 GND.n2593 0.152939
R9414 GND.n2602 GND.n2593 0.152939
R9415 GND.n2603 GND.n2602 0.152939
R9416 GND.n2604 GND.n2603 0.152939
R9417 GND.n2604 GND.n2589 0.152939
R9418 GND.n2612 GND.n2589 0.152939
R9419 GND.n2613 GND.n2612 0.152939
R9420 GND.n2614 GND.n2613 0.152939
R9421 GND.n2614 GND.n2582 0.152939
R9422 GND.n2622 GND.n2582 0.152939
R9423 GND.n2623 GND.n2622 0.152939
R9424 GND.n2624 GND.n2623 0.152939
R9425 GND.n2624 GND.n2578 0.152939
R9426 GND.n2632 GND.n2578 0.152939
R9427 GND.n2633 GND.n2632 0.152939
R9428 GND.n2634 GND.n2633 0.152939
R9429 GND.n2634 GND.n2574 0.152939
R9430 GND.n2642 GND.n2574 0.152939
R9431 GND.n2643 GND.n2642 0.152939
R9432 GND.n2645 GND.n2643 0.152939
R9433 GND.n2645 GND.n2644 0.152939
R9434 GND.n2644 GND.n2570 0.152939
R9435 GND.n2654 GND.n2570 0.152939
R9436 GND.n2655 GND.n2654 0.152939
R9437 GND.n2655 GND.n2564 0.152939
R9438 GND.n2663 GND.n2564 0.152939
R9439 GND.n2664 GND.n2663 0.152939
R9440 GND.n2665 GND.n2664 0.152939
R9441 GND.n2665 GND.n2560 0.152939
R9442 GND.n2673 GND.n2560 0.152939
R9443 GND.n2674 GND.n2673 0.152939
R9444 GND.n2675 GND.n2674 0.152939
R9445 GND.n2675 GND.n2556 0.152939
R9446 GND.n2683 GND.n2556 0.152939
R9447 GND.n2684 GND.n2683 0.152939
R9448 GND.n2685 GND.n2684 0.152939
R9449 GND.n2685 GND.n2552 0.152939
R9450 GND.n2695 GND.n2552 0.152939
R9451 GND.n2696 GND.n2695 0.152939
R9452 GND.n2697 GND.n2696 0.152939
R9453 GND.n2697 GND.n2548 0.152939
R9454 GND.n2705 GND.n2548 0.152939
R9455 GND.n2706 GND.n2705 0.152939
R9456 GND.n2707 GND.n2706 0.152939
R9457 GND.n2707 GND.n2544 0.152939
R9458 GND.n2715 GND.n2544 0.152939
R9459 GND.n2716 GND.n2715 0.152939
R9460 GND.n2717 GND.n2716 0.152939
R9461 GND.n2717 GND.n2538 0.152939
R9462 GND.n2724 GND.n2538 0.152939
R9463 GND.n1364 GND.n1363 0.152939
R9464 GND.n1365 GND.n1364 0.152939
R9465 GND.n2429 GND.n1365 0.152939
R9466 GND.n2430 GND.n2429 0.152939
R9467 GND.n1144 GND.n1143 0.152939
R9468 GND.n1145 GND.n1144 0.152939
R9469 GND.n1150 GND.n1145 0.152939
R9470 GND.n1151 GND.n1150 0.152939
R9471 GND.n1152 GND.n1151 0.152939
R9472 GND.n1153 GND.n1152 0.152939
R9473 GND.n1158 GND.n1153 0.152939
R9474 GND.n1159 GND.n1158 0.152939
R9475 GND.n1160 GND.n1159 0.152939
R9476 GND.n1161 GND.n1160 0.152939
R9477 GND.n1166 GND.n1161 0.152939
R9478 GND.n1167 GND.n1166 0.152939
R9479 GND.n1168 GND.n1167 0.152939
R9480 GND.n1169 GND.n1168 0.152939
R9481 GND.n1174 GND.n1169 0.152939
R9482 GND.n1175 GND.n1174 0.152939
R9483 GND.n1176 GND.n1175 0.152939
R9484 GND.n1177 GND.n1176 0.152939
R9485 GND.n1182 GND.n1177 0.152939
R9486 GND.n1183 GND.n1182 0.152939
R9487 GND.n1184 GND.n1183 0.152939
R9488 GND.n1185 GND.n1184 0.152939
R9489 GND.n1190 GND.n1185 0.152939
R9490 GND.n1191 GND.n1190 0.152939
R9491 GND.n1192 GND.n1191 0.152939
R9492 GND.n1193 GND.n1192 0.152939
R9493 GND.n1198 GND.n1193 0.152939
R9494 GND.n1199 GND.n1198 0.152939
R9495 GND.n1200 GND.n1199 0.152939
R9496 GND.n1201 GND.n1200 0.152939
R9497 GND.n1206 GND.n1201 0.152939
R9498 GND.n1207 GND.n1206 0.152939
R9499 GND.n1208 GND.n1207 0.152939
R9500 GND.n1209 GND.n1208 0.152939
R9501 GND.n1214 GND.n1209 0.152939
R9502 GND.n1215 GND.n1214 0.152939
R9503 GND.n1216 GND.n1215 0.152939
R9504 GND.n1217 GND.n1216 0.152939
R9505 GND.n1222 GND.n1217 0.152939
R9506 GND.n1223 GND.n1222 0.152939
R9507 GND.n1224 GND.n1223 0.152939
R9508 GND.n1225 GND.n1224 0.152939
R9509 GND.n1230 GND.n1225 0.152939
R9510 GND.n1231 GND.n1230 0.152939
R9511 GND.n1232 GND.n1231 0.152939
R9512 GND.n1233 GND.n1232 0.152939
R9513 GND.n1238 GND.n1233 0.152939
R9514 GND.n1239 GND.n1238 0.152939
R9515 GND.n1240 GND.n1239 0.152939
R9516 GND.n1241 GND.n1240 0.152939
R9517 GND.n1246 GND.n1241 0.152939
R9518 GND.n1247 GND.n1246 0.152939
R9519 GND.n1248 GND.n1247 0.152939
R9520 GND.n1249 GND.n1248 0.152939
R9521 GND.n1254 GND.n1249 0.152939
R9522 GND.n1255 GND.n1254 0.152939
R9523 GND.n1256 GND.n1255 0.152939
R9524 GND.n1257 GND.n1256 0.152939
R9525 GND.n1262 GND.n1257 0.152939
R9526 GND.n1263 GND.n1262 0.152939
R9527 GND.n1264 GND.n1263 0.152939
R9528 GND.n1265 GND.n1264 0.152939
R9529 GND.n1270 GND.n1265 0.152939
R9530 GND.n1271 GND.n1270 0.152939
R9531 GND.n1272 GND.n1271 0.152939
R9532 GND.n1273 GND.n1272 0.152939
R9533 GND.n1278 GND.n1273 0.152939
R9534 GND.n1279 GND.n1278 0.152939
R9535 GND.n1280 GND.n1279 0.152939
R9536 GND.n1281 GND.n1280 0.152939
R9537 GND.n1286 GND.n1281 0.152939
R9538 GND.n1287 GND.n1286 0.152939
R9539 GND.n1288 GND.n1287 0.152939
R9540 GND.n1289 GND.n1288 0.152939
R9541 GND.n1294 GND.n1289 0.152939
R9542 GND.n1295 GND.n1294 0.152939
R9543 GND.n1296 GND.n1295 0.152939
R9544 GND.n1297 GND.n1296 0.152939
R9545 GND.n1302 GND.n1297 0.152939
R9546 GND.n1303 GND.n1302 0.152939
R9547 GND.n1304 GND.n1303 0.152939
R9548 GND.n1305 GND.n1304 0.152939
R9549 GND.n1310 GND.n1305 0.152939
R9550 GND.n1311 GND.n1310 0.152939
R9551 GND.n1312 GND.n1311 0.152939
R9552 GND.n1313 GND.n1312 0.152939
R9553 GND.n1318 GND.n1313 0.152939
R9554 GND.n1319 GND.n1318 0.152939
R9555 GND.n1320 GND.n1319 0.152939
R9556 GND.n1321 GND.n1320 0.152939
R9557 GND.n1326 GND.n1321 0.152939
R9558 GND.n1327 GND.n1326 0.152939
R9559 GND.n1328 GND.n1327 0.152939
R9560 GND.n1329 GND.n1328 0.152939
R9561 GND.n1334 GND.n1329 0.152939
R9562 GND.n1335 GND.n1334 0.152939
R9563 GND.n1336 GND.n1335 0.152939
R9564 GND.n1337 GND.n1336 0.152939
R9565 GND.n1342 GND.n1337 0.152939
R9566 GND.n1343 GND.n1342 0.152939
R9567 GND.n1344 GND.n1343 0.152939
R9568 GND.n1345 GND.n1344 0.152939
R9569 GND.n1350 GND.n1345 0.152939
R9570 GND.n1351 GND.n1350 0.152939
R9571 GND.n1352 GND.n1351 0.152939
R9572 GND.n1353 GND.n1352 0.152939
R9573 GND.n2441 GND.n1353 0.152939
R9574 GND.n2442 GND.n2441 0.152939
R9575 GND.n2443 GND.n2442 0.152939
R9576 GND.n2444 GND.n2443 0.152939
R9577 GND.n1032 GND.n1031 0.152939
R9578 GND.n1033 GND.n1032 0.152939
R9579 GND.n1038 GND.n1033 0.152939
R9580 GND.n1039 GND.n1038 0.152939
R9581 GND.n1040 GND.n1039 0.152939
R9582 GND.n1041 GND.n1040 0.152939
R9583 GND.n1046 GND.n1041 0.152939
R9584 GND.n1047 GND.n1046 0.152939
R9585 GND.n1048 GND.n1047 0.152939
R9586 GND.n1049 GND.n1048 0.152939
R9587 GND.n1054 GND.n1049 0.152939
R9588 GND.n1055 GND.n1054 0.152939
R9589 GND.n1056 GND.n1055 0.152939
R9590 GND.n1057 GND.n1056 0.152939
R9591 GND.n1062 GND.n1057 0.152939
R9592 GND.n1063 GND.n1062 0.152939
R9593 GND.n1064 GND.n1063 0.152939
R9594 GND.n1065 GND.n1064 0.152939
R9595 GND.n1070 GND.n1065 0.152939
R9596 GND.n1071 GND.n1070 0.152939
R9597 GND.n1072 GND.n1071 0.152939
R9598 GND.n1073 GND.n1072 0.152939
R9599 GND.n1078 GND.n1073 0.152939
R9600 GND.n1079 GND.n1078 0.152939
R9601 GND.n1080 GND.n1079 0.152939
R9602 GND.n1081 GND.n1080 0.152939
R9603 GND.n1086 GND.n1081 0.152939
R9604 GND.n1087 GND.n1086 0.152939
R9605 GND.n1088 GND.n1087 0.152939
R9606 GND.n1089 GND.n1088 0.152939
R9607 GND.n1094 GND.n1089 0.152939
R9608 GND.n1095 GND.n1094 0.152939
R9609 GND.n1096 GND.n1095 0.152939
R9610 GND.n1097 GND.n1096 0.152939
R9611 GND.n1102 GND.n1097 0.152939
R9612 GND.n1103 GND.n1102 0.152939
R9613 GND.n1104 GND.n1103 0.152939
R9614 GND.n1105 GND.n1104 0.152939
R9615 GND.n1110 GND.n1105 0.152939
R9616 GND.n1111 GND.n1110 0.152939
R9617 GND.n1112 GND.n1111 0.152939
R9618 GND.n1113 GND.n1112 0.152939
R9619 GND.n1118 GND.n1113 0.152939
R9620 GND.n1119 GND.n1118 0.152939
R9621 GND.n1120 GND.n1119 0.152939
R9622 GND.n1121 GND.n1120 0.152939
R9623 GND.n1126 GND.n1121 0.152939
R9624 GND.n1127 GND.n1126 0.152939
R9625 GND.n1128 GND.n1127 0.152939
R9626 GND.n1129 GND.n1128 0.152939
R9627 GND.n1134 GND.n1129 0.152939
R9628 GND.n1135 GND.n1134 0.152939
R9629 GND.n1136 GND.n1135 0.152939
R9630 GND.n1137 GND.n1136 0.152939
R9631 GND.n1142 GND.n1137 0.152939
R9632 GND.n2790 GND.n2398 0.152939
R9633 GND.n2813 GND.n2398 0.152939
R9634 GND.n2814 GND.n2813 0.152939
R9635 GND.n2821 GND.n2814 0.152939
R9636 GND.n2821 GND.n2820 0.152939
R9637 GND.n2820 GND.n2819 0.152939
R9638 GND.n2819 GND.n2815 0.152939
R9639 GND.n2815 GND.n2378 0.152939
R9640 GND.n2843 GND.n2378 0.152939
R9641 GND.n3946 GND.n1420 0.152939
R9642 GND.n3942 GND.n1420 0.152939
R9643 GND.n3942 GND.n3941 0.152939
R9644 GND.n3941 GND.n3940 0.152939
R9645 GND.n3940 GND.n1424 0.152939
R9646 GND.n3936 GND.n1424 0.152939
R9647 GND.n3936 GND.n3935 0.152939
R9648 GND.n3935 GND.n3934 0.152939
R9649 GND.n3934 GND.n1429 0.152939
R9650 GND.n3930 GND.n1429 0.152939
R9651 GND.n3930 GND.n3929 0.152939
R9652 GND.n3929 GND.n1436 0.152939
R9653 GND.n3925 GND.n1436 0.152939
R9654 GND.n3925 GND.n3924 0.152939
R9655 GND.n3924 GND.n3923 0.152939
R9656 GND.n3923 GND.n1441 0.152939
R9657 GND.n3919 GND.n1441 0.152939
R9658 GND.n3919 GND.n3918 0.152939
R9659 GND.n3918 GND.n3917 0.152939
R9660 GND.n3917 GND.n1446 0.152939
R9661 GND.n1449 GND.n1446 0.152939
R9662 GND.n3907 GND.n3906 0.152939
R9663 GND.n3906 GND.n3905 0.152939
R9664 GND.n3905 GND.n1471 0.152939
R9665 GND.n3901 GND.n1471 0.152939
R9666 GND.n3901 GND.n3900 0.152939
R9667 GND.n3900 GND.n3899 0.152939
R9668 GND.n3899 GND.n1478 0.152939
R9669 GND.n3895 GND.n1478 0.152939
R9670 GND.n3895 GND.n3894 0.152939
R9671 GND.n3894 GND.n3893 0.152939
R9672 GND.n3893 GND.n1486 0.152939
R9673 GND.n1493 GND.n1486 0.152939
R9674 GND.n3888 GND.n1493 0.152939
R9675 GND.n3888 GND.n3887 0.152939
R9676 GND.n3887 GND.n3886 0.152939
R9677 GND.n3886 GND.n1498 0.152939
R9678 GND.n3882 GND.n1498 0.152939
R9679 GND.n3882 GND.n3881 0.152939
R9680 GND.n3881 GND.n3880 0.152939
R9681 GND.n3880 GND.n1506 0.152939
R9682 GND.n3876 GND.n1506 0.152939
R9683 GND.n3876 GND.n3875 0.152939
R9684 GND.n3875 GND.n3874 0.152939
R9685 GND.n3874 GND.n1514 0.152939
R9686 GND.n1522 GND.n1514 0.152939
R9687 GND.n3869 GND.n1522 0.152939
R9688 GND.n2730 GND.n2729 0.152939
R9689 GND.n2730 GND.n2534 0.152939
R9690 GND.n2738 GND.n2534 0.152939
R9691 GND.n2739 GND.n2738 0.152939
R9692 GND.n2740 GND.n2739 0.152939
R9693 GND.n2740 GND.n2530 0.152939
R9694 GND.n2748 GND.n2530 0.152939
R9695 GND.n2749 GND.n2748 0.152939
R9696 GND.n2750 GND.n2749 0.152939
R9697 GND.n2750 GND.n2523 0.152939
R9698 GND.n2757 GND.n2523 0.152939
R9699 GND.n2758 GND.n2522 0.152939
R9700 GND.n2765 GND.n2522 0.152939
R9701 GND.n2766 GND.n2765 0.152939
R9702 GND.n2768 GND.n2766 0.152939
R9703 GND.n2768 GND.n2767 0.152939
R9704 GND.n2767 GND.n2419 0.152939
R9705 GND.n2788 GND.n2419 0.152939
R9706 GND.n2789 GND.n2788 0.152939
R9707 GND.n2792 GND.n2789 0.152939
R9708 GND.n3344 GND.n20 0.0919634
R9709 GND.n2511 GND.n2444 0.0919634
R9710 GND.n5496 GND.n18 0.0767195
R9711 GND.n5496 GND.n19 0.0767195
R9712 GND.n2831 GND.n2387 0.0767195
R9713 GND.n2430 GND.n2387 0.0767195
R9714 GND.n5504 GND.n5 0.0695946
R9715 GND.n5504 GND.n5503 0.0695946
R9716 GND.n2791 GND.n2790 0.0695946
R9717 GND.n2792 GND.n2791 0.0695946
R9718 GND.n3867 GND.n1525 0.063
R9719 GND.n2142 GND.n1929 0.063
R9720 GND.n2143 GND.n2142 0.063
R9721 GND.n3868 GND.n3867 0.063
R9722 GND.n2511 GND.n2447 0.0614756
R9723 GND.n2210 GND.n20 0.0614756
R9724 GND.n2151 GND.n2143 0.0534891
R9725 GND.n5477 GND.n57 0.0534891
R9726 GND.n2728 GND.n2727 0.0534891
R9727 GND.n3868 GND.n1408 0.0534891
R9728 GND.n3224 GND.n2252 0.044054
R9729 GND.n3225 GND.n3224 0.044054
R9730 GND.n3226 GND.n3225 0.044054
R9731 GND.n3226 GND.n2248 0.044054
R9732 GND.n3234 GND.n2248 0.044054
R9733 GND.n2853 GND.n2360 0.044054
R9734 GND.n2853 GND.n2852 0.044054
R9735 GND.n2852 GND.n2851 0.044054
R9736 GND.n2851 GND.n2371 0.044054
R9737 GND.n2844 GND.n2371 0.044054
R9738 GND.n3216 GND.n2252 0.0417311
R9739 GND.n2857 GND.n2360 0.0417311
R9740 GND.n3397 GND.n2151 0.0344674
R9741 GND.n3397 GND.n2153 0.0344674
R9742 GND.n2177 GND.n2153 0.0344674
R9743 GND.n2178 GND.n2177 0.0344674
R9744 GND.n2179 GND.n2178 0.0344674
R9745 GND.n2180 GND.n2179 0.0344674
R9746 GND.n3259 GND.n2180 0.0344674
R9747 GND.n3260 GND.n3259 0.0344674
R9748 GND.n3260 GND.n2225 0.0344674
R9749 GND.n2226 GND.n2225 0.0344674
R9750 GND.n2227 GND.n2226 0.0344674
R9751 GND.n3268 GND.n2227 0.0344674
R9752 GND.n3269 GND.n3268 0.0344674
R9753 GND.n3269 GND.n36 0.0344674
R9754 GND.n37 GND.n36 0.0344674
R9755 GND.n38 GND.n37 0.0344674
R9756 GND.n3272 GND.n38 0.0344674
R9757 GND.n3272 GND.n56 0.0344674
R9758 GND.n5477 GND.n56 0.0344674
R9759 GND.n2727 GND.n1375 0.0344674
R9760 GND.n3978 GND.n1375 0.0344674
R9761 GND.n3978 GND.n1376 0.0344674
R9762 GND.n3974 GND.n1376 0.0344674
R9763 GND.n3974 GND.n3973 0.0344674
R9764 GND.n3973 GND.n3972 0.0344674
R9765 GND.n3972 GND.n1384 0.0344674
R9766 GND.n3968 GND.n1384 0.0344674
R9767 GND.n3968 GND.n3967 0.0344674
R9768 GND.n3967 GND.n3966 0.0344674
R9769 GND.n3966 GND.n1392 0.0344674
R9770 GND.n3962 GND.n1392 0.0344674
R9771 GND.n3962 GND.n3961 0.0344674
R9772 GND.n3961 GND.n3960 0.0344674
R9773 GND.n3960 GND.n1400 0.0344674
R9774 GND.n3956 GND.n1400 0.0344674
R9775 GND.n3956 GND.n3955 0.0344674
R9776 GND.n3955 GND.n3954 0.0344674
R9777 GND.n3954 GND.n1408 0.0344674
R9778 GND.n1934 GND.n1930 0.0343753
R9779 GND.n3214 GND.n3213 0.0343753
R9780 GND.n3866 GND.n1526 0.0343753
R9781 GND.n2359 GND.n1540 0.0343753
R9782 GND.n3202 GND.n1935 0.0340366
R9783 GND.n3204 GND.n1936 0.0340366
R9784 GND.n3206 GND.n1937 0.0340366
R9785 GND.n3859 GND.n1532 0.0340366
R9786 GND.n3858 GND.n1533 0.0340366
R9787 GND.n3855 GND.n3854 0.0340366
R9788 GND.n3215 GND.n3214 0.0286165
R9789 GND.n2858 GND.n2359 0.0286165
R9790 GND.n2142 GND.n1930 0.0204865
R9791 GND.n3867 GND.n3866 0.0204865
R9792 GND.n3216 GND.n3215 0.00625881
R9793 GND.n2858 GND.n2857 0.00625881
R9794 GND.n3202 GND.n1934 0.000838753
R9795 GND.n3204 GND.n1935 0.000838753
R9796 GND.n3206 GND.n1936 0.000838753
R9797 GND.n3213 GND.n1937 0.000838753
R9798 GND.n1532 GND.n1526 0.000838753
R9799 GND.n3859 GND.n3858 0.000838753
R9800 GND.n3855 GND.n1533 0.000838753
R9801 GND.n3854 GND.n1540 0.000838753
R9802 a_n14320_7092.n24 a_n14320_7092.t7 120.427
R9803 a_n14320_7092.n15 a_n14320_7092.t6 113.434
R9804 a_n14320_7092.n14 a_n14320_7092.t5 110.305
R9805 a_n14320_7092.n14 a_n14320_7092.t3 107.061
R9806 a_n14320_7092.n14 a_n14320_7092.t2 103.931
R9807 a_n14320_7092.n15 a_n14320_7092.t1 103.931
R9808 a_n14320_7092.t0 a_n14320_7092.n15 103.931
R9809 a_n14320_7092.n24 a_n14320_7092.t4 88.2359
R9810 a_n14320_7092.n5 a_n14320_7092.t21 44.664
R9811 a_n14320_7092.n4 a_n14320_7092.t39 44.664
R9812 a_n14320_7092.n4 a_n14320_7092.t16 44.664
R9813 a_n14320_7092.n4 a_n14320_7092.t28 44.664
R9814 a_n14320_7092.n11 a_n14320_7092.t46 44.664
R9815 a_n14320_7092.n23 a_n14320_7092.t38 46.6563
R9816 a_n14320_7092.n17 a_n14320_7092.t15 46.6561
R9817 a_n14320_7092.n18 a_n14320_7092.t32 46.6561
R9818 a_n14320_7092.n19 a_n14320_7092.t9 46.6561
R9819 a_n14320_7092.n20 a_n14320_7092.t22 46.6561
R9820 a_n14320_7092.n6 a_n14320_7092.n16 1.80487
R9821 a_n14320_7092.n6 a_n14320_7092.n17 2.05575
R9822 a_n14320_7092.n1 a_n14320_7092.n18 2.05575
R9823 a_n14320_7092.n1 a_n14320_7092.n19 2.05575
R9824 a_n14320_7092.n1 a_n14320_7092.n20 2.05575
R9825 a_n14320_7092.n22 a_n14320_7092.n23 2.05575
R9826 a_n14320_7092.n22 a_n14320_7092.n21 1.80487
R9827 a_n14320_7092.n13 a_n14320_7092.n24 12.4106
R9828 a_n14320_7092.n25 a_n14320_7092.n13 11.4887
R9829 a_n14320_7092.n16 a_n14320_7092.t8 45.0831
R9830 a_n14320_7092.n16 a_n14320_7092.t35 42.079
R9831 a_n14320_7092.n17 a_n14320_7092.t40 41.9024
R9832 a_n14320_7092.n0 a_n14320_7092.t24 45.0831
R9833 a_n14320_7092.n0 a_n14320_7092.t14 42.079
R9834 a_n14320_7092.n18 a_n14320_7092.t19 41.9024
R9835 a_n14320_7092.n2 a_n14320_7092.t42 45.0831
R9836 a_n14320_7092.n2 a_n14320_7092.t29 42.079
R9837 a_n14320_7092.n19 a_n14320_7092.t34 41.9024
R9838 a_n14320_7092.n3 a_n14320_7092.t17 45.0831
R9839 a_n14320_7092.n3 a_n14320_7092.t37 42.079
R9840 a_n14320_7092.n20 a_n14320_7092.t36 41.9024
R9841 a_n14320_7092.n23 a_n14320_7092.t12 41.9024
R9842 a_n14320_7092.n21 a_n14320_7092.t13 42.079
R9843 a_n14320_7092.n21 a_n14320_7092.t31 45.0831
R9844 a_n14320_7092.n7 a_n14320_7092.t47 45.224
R9845 a_n14320_7092.n7 a_n14320_7092.t30 41.7162
R9846 a_n14320_7092.n5 a_n14320_7092.t11 44.8812
R9847 a_n14320_7092.n8 a_n14320_7092.t23 45.224
R9848 a_n14320_7092.n8 a_n14320_7092.t10 41.7162
R9849 a_n14320_7092.n4 a_n14320_7092.t26 44.8812
R9850 a_n14320_7092.n9 a_n14320_7092.t41 45.224
R9851 a_n14320_7092.n9 a_n14320_7092.t25 41.7162
R9852 a_n14320_7092.n4 a_n14320_7092.t44 44.8812
R9853 a_n14320_7092.n10 a_n14320_7092.t43 45.224
R9854 a_n14320_7092.n10 a_n14320_7092.t18 41.7162
R9855 a_n14320_7092.n4 a_n14320_7092.t27 44.8812
R9856 a_n14320_7092.n12 a_n14320_7092.t20 45.224
R9857 a_n14320_7092.n12 a_n14320_7092.t33 41.7162
R9858 a_n14320_7092.n11 a_n14320_7092.t45 44.8812
R9859 a_n14320_7092.n5 a_n14320_7092.n7 2.54617
R9860 a_n14320_7092.n11 a_n14320_7092.n12 2.54617
R9861 a_n14320_7092.n25 a_n14320_7092.n14 46.0782
R9862 a_n14320_7092.n15 a_n14320_7092.n25 38.9319
R9863 a_n14320_7092.n1 a_n14320_7092.n6 10.6887
R9864 a_n14320_7092.n4 a_n14320_7092.n5 10.6887
R9865 a_n14320_7092.n13 a_n14320_7092.n1 9.91667
R9866 a_n14320_7092.n4 a_n14320_7092.n10 7.98439
R9867 a_n14320_7092.n4 a_n14320_7092.n9 7.98439
R9868 a_n14320_7092.n4 a_n14320_7092.n8 7.98439
R9869 a_n14320_7092.n1 a_n14320_7092.n3 7.24309
R9870 a_n14320_7092.n1 a_n14320_7092.n2 7.24309
R9871 a_n14320_7092.n1 a_n14320_7092.n0 7.24309
R9872 a_n14320_7092.n1 a_n14320_7092.n22 7.18872
R9873 a_n14320_7092.n4 a_n14320_7092.n11 7.18872
R9874 a_n14320_7092.n13 a_n14320_7092.n4 6.65362
R9875 VOUT.n47 VOUT.n45 157.475
R9876 VOUT.n43 VOUT.n41 157.475
R9877 VOUT.n39 VOUT.n37 157.475
R9878 VOUT.n35 VOUT.n33 157.475
R9879 VOUT.n32 VOUT.n30 157.475
R9880 VOUT.n17 VOUT.n15 157.475
R9881 VOUT.n13 VOUT.n11 157.475
R9882 VOUT.n9 VOUT.n7 157.475
R9883 VOUT.n5 VOUT.n3 157.475
R9884 VOUT.n2 VOUT.n0 157.475
R9885 VOUT.n43 VOUT.n42 152.69
R9886 VOUT.n39 VOUT.n38 152.69
R9887 VOUT.n35 VOUT.n34 152.69
R9888 VOUT.n32 VOUT.n31 152.69
R9889 VOUT.n17 VOUT.n16 152.69
R9890 VOUT.n13 VOUT.n12 152.69
R9891 VOUT.n9 VOUT.n8 152.69
R9892 VOUT.n5 VOUT.n4 152.69
R9893 VOUT.n2 VOUT.n1 152.69
R9894 VOUT.n47 VOUT.n46 152.69
R9895 VOUT.n50 VOUT.t45 85.2228
R9896 VOUT.n54 VOUT.t1 84.2012
R9897 VOUT.n52 VOUT.t3 82.5072
R9898 VOUT.n51 VOUT.t0 82.5072
R9899 VOUT.n50 VOUT.t47 82.5072
R9900 VOUT.n56 VOUT.t46 81.4857
R9901 VOUT.n55 VOUT.t44 81.4857
R9902 VOUT.n54 VOUT.t2 81.4857
R9903 VOUT.n46 VOUT.t33 13.2678
R9904 VOUT.n46 VOUT.t24 13.2678
R9905 VOUT.n45 VOUT.t18 13.2678
R9906 VOUT.n45 VOUT.t9 13.2678
R9907 VOUT.n42 VOUT.t30 13.2678
R9908 VOUT.n42 VOUT.t28 13.2678
R9909 VOUT.n41 VOUT.t14 13.2678
R9910 VOUT.n41 VOUT.t29 13.2678
R9911 VOUT.n38 VOUT.t43 13.2678
R9912 VOUT.n38 VOUT.t4 13.2678
R9913 VOUT.n37 VOUT.t39 13.2678
R9914 VOUT.n37 VOUT.t11 13.2678
R9915 VOUT.n34 VOUT.t22 13.2678
R9916 VOUT.n34 VOUT.t17 13.2678
R9917 VOUT.n33 VOUT.t26 13.2678
R9918 VOUT.n33 VOUT.t8 13.2678
R9919 VOUT.n31 VOUT.t19 13.2678
R9920 VOUT.n31 VOUT.t7 13.2678
R9921 VOUT.n30 VOUT.t5 13.2678
R9922 VOUT.n30 VOUT.t42 13.2678
R9923 VOUT.n15 VOUT.t16 13.2678
R9924 VOUT.n15 VOUT.t6 13.2678
R9925 VOUT.n16 VOUT.t25 13.2678
R9926 VOUT.n16 VOUT.t21 13.2678
R9927 VOUT.n11 VOUT.t13 13.2678
R9928 VOUT.n11 VOUT.t36 13.2678
R9929 VOUT.n12 VOUT.t12 13.2678
R9930 VOUT.n12 VOUT.t32 13.2678
R9931 VOUT.n7 VOUT.t38 13.2678
R9932 VOUT.n7 VOUT.t31 13.2678
R9933 VOUT.n8 VOUT.t15 13.2678
R9934 VOUT.n8 VOUT.t40 13.2678
R9935 VOUT.n3 VOUT.t35 13.2678
R9936 VOUT.n3 VOUT.t37 13.2678
R9937 VOUT.n4 VOUT.t23 13.2678
R9938 VOUT.n4 VOUT.t27 13.2678
R9939 VOUT.n0 VOUT.t10 13.2678
R9940 VOUT.n0 VOUT.t34 13.2678
R9941 VOUT.n1 VOUT.t20 13.2678
R9942 VOUT.n1 VOUT.t41 13.2678
R9943 VOUT.n53 VOUT.n49 10.0047
R9944 VOUT.n36 VOUT.n32 9.76774
R9945 VOUT.n6 VOUT.n2 9.76774
R9946 VOUT.n48 VOUT.n47 7.7936
R9947 VOUT.n44 VOUT.n43 7.7936
R9948 VOUT.n40 VOUT.n39 7.7936
R9949 VOUT.n36 VOUT.n35 7.7936
R9950 VOUT.n18 VOUT.n17 7.7936
R9951 VOUT.n14 VOUT.n13 7.7936
R9952 VOUT.n10 VOUT.n9 7.7936
R9953 VOUT.n6 VOUT.n5 7.7936
R9954 VOUT.n49 VOUT.n48 6.31567
R9955 VOUT.n19 VOUT.n18 6.31567
R9956 VOUT.n53 VOUT.n52 5.58291
R9957 VOUT.n57 VOUT.n56 5.58291
R9958 VOUT.n58 VOUT.n57 5.25635
R9959 VOUT.n58 VOUT.n19 4.72936
R9960 VOUT.n49 VOUT.n19 4.67105
R9961 VOUT.n29 VOUT 3.41035
R9962 VOUT.n51 VOUT.n50 2.71602
R9963 VOUT.n52 VOUT.n51 2.71602
R9964 VOUT.n55 VOUT.n54 2.71602
R9965 VOUT.n56 VOUT.n55 2.71602
R9966 VOUT.n40 VOUT.n36 1.97464
R9967 VOUT.n44 VOUT.n40 1.97464
R9968 VOUT.n48 VOUT.n44 1.97464
R9969 VOUT.n10 VOUT.n6 1.97464
R9970 VOUT.n14 VOUT.n10 1.97464
R9971 VOUT.n18 VOUT.n14 1.97464
R9972 VOUT.n57 VOUT.n53 1.56341
R9973 VOUT.n29 VOUT.n28 0.343116
R9974 VOUT.n58 VOUT.n29 0.332085
R9975 VOUT.n22 VOUT.n21 0.0947519
R9976 VOUT.n27 VOUT.n26 0.0947519
R9977 VOUT.n24 VOUT.n23 0.0947519
R9978 VOUT.n21 VOUT.t50 0.056164
R9979 VOUT.n23 VOUT.t48 0.056164
R9980 VOUT.n27 VOUT.t52 0.056164
R9981 VOUT.n22 VOUT.t53 0.0555192
R9982 VOUT.n24 VOUT.t51 0.0555192
R9983 VOUT.n26 VOUT.t49 0.0555192
R9984 VOUT.n21 VOUT.n20 0.0480384
R9985 VOUT.n25 VOUT.n22 0.0466438
R9986 VOUT.n26 VOUT.n25 0.0466438
R9987 VOUT.n28 VOUT.n20 0.0391444
R9988 VOUT VOUT.n58 0.0099
R9989 VOUT.n23 VOUT.n20 0.00939398
R9990 VOUT.n28 VOUT.n27 0.00939398
R9991 VOUT.n25 VOUT.n24 0.00799933
R9992 VDD.n138 VDD.n132 756.745
R9993 VDD.n125 VDD.n119 756.745
R9994 VDD.n112 VDD.n106 756.745
R9995 VDD.n99 VDD.n93 756.745
R9996 VDD.n86 VDD.n80 756.745
R9997 VDD.n73 VDD.n67 756.745
R9998 VDD.n60 VDD.n54 756.745
R9999 VDD.n47 VDD.n41 756.745
R10000 VDD.n35 VDD.n29 756.745
R10001 VDD.n22 VDD.n16 756.745
R10002 VDD.n1731 VDD.n1725 756.745
R10003 VDD.n1744 VDD.n1738 756.745
R10004 VDD.n1705 VDD.n1699 756.745
R10005 VDD.n1718 VDD.n1712 756.745
R10006 VDD.n1679 VDD.n1673 756.745
R10007 VDD.n1692 VDD.n1686 756.745
R10008 VDD.n1653 VDD.n1647 756.745
R10009 VDD.n1666 VDD.n1660 756.745
R10010 VDD.n1628 VDD.n1622 756.745
R10011 VDD.n1641 VDD.n1635 756.745
R10012 VDD.n139 VDD.n138 585
R10013 VDD.n137 VDD.n136 585
R10014 VDD.n126 VDD.n125 585
R10015 VDD.n124 VDD.n123 585
R10016 VDD.n113 VDD.n112 585
R10017 VDD.n111 VDD.n110 585
R10018 VDD.n100 VDD.n99 585
R10019 VDD.n98 VDD.n97 585
R10020 VDD.n87 VDD.n86 585
R10021 VDD.n85 VDD.n84 585
R10022 VDD.n74 VDD.n73 585
R10023 VDD.n72 VDD.n71 585
R10024 VDD.n61 VDD.n60 585
R10025 VDD.n59 VDD.n58 585
R10026 VDD.n48 VDD.n47 585
R10027 VDD.n46 VDD.n45 585
R10028 VDD.n36 VDD.n35 585
R10029 VDD.n34 VDD.n33 585
R10030 VDD.n23 VDD.n22 585
R10031 VDD.n21 VDD.n20 585
R10032 VDD.n1732 VDD.n1731 585
R10033 VDD.n1730 VDD.n1729 585
R10034 VDD.n1745 VDD.n1744 585
R10035 VDD.n1743 VDD.n1742 585
R10036 VDD.n1706 VDD.n1705 585
R10037 VDD.n1704 VDD.n1703 585
R10038 VDD.n1719 VDD.n1718 585
R10039 VDD.n1717 VDD.n1716 585
R10040 VDD.n1680 VDD.n1679 585
R10041 VDD.n1678 VDD.n1677 585
R10042 VDD.n1693 VDD.n1692 585
R10043 VDD.n1691 VDD.n1690 585
R10044 VDD.n1654 VDD.n1653 585
R10045 VDD.n1652 VDD.n1651 585
R10046 VDD.n1667 VDD.n1666 585
R10047 VDD.n1665 VDD.n1664 585
R10048 VDD.n1629 VDD.n1628 585
R10049 VDD.n1627 VDD.n1626 585
R10050 VDD.n1642 VDD.n1641 585
R10051 VDD.n1640 VDD.n1639 585
R10052 VDD.n3877 VDD.n243 510.733
R10053 VDD.n3788 VDD.n3787 510.733
R10054 VDD.n3579 VDD.n449 510.733
R10055 VDD.n3581 VDD.n447 510.733
R10056 VDD.n2211 VDD.n1100 510.733
R10057 VDD.n2213 VDD.n1092 510.733
R10058 VDD.n1481 VDD.n1309 510.733
R10059 VDD.n1478 VDD.n1307 510.733
R10060 VDD.n135 VDD.t142 355.474
R10061 VDD.n122 VDD.t151 355.474
R10062 VDD.n109 VDD.t160 355.474
R10063 VDD.n96 VDD.t165 355.474
R10064 VDD.n83 VDD.t173 355.474
R10065 VDD.n70 VDD.t136 355.474
R10066 VDD.n57 VDD.t150 355.474
R10067 VDD.n44 VDD.t158 355.474
R10068 VDD.n32 VDD.t167 355.474
R10069 VDD.n19 VDD.t174 355.474
R10070 VDD.n1728 VDD.t132 355.474
R10071 VDD.n1741 VDD.t130 355.474
R10072 VDD.n1702 VDD.t155 355.474
R10073 VDD.n1715 VDD.t154 355.474
R10074 VDD.n1676 VDD.t133 355.474
R10075 VDD.n1689 VDD.t166 355.474
R10076 VDD.n1650 VDD.t156 355.474
R10077 VDD.n1663 VDD.t140 355.474
R10078 VDD.n1625 VDD.t171 355.474
R10079 VDD.n1638 VDD.t161 355.474
R10080 VDD.n1312 VDD.t57 330.918
R10081 VDD.n1414 VDD.t108 330.918
R10082 VDD.n1371 VDD.t70 330.918
R10083 VDD.n1447 VDD.t79 330.918
R10084 VDD.n1464 VDD.t54 330.918
R10085 VDD.n2218 VDD.t110 330.918
R10086 VDD.n1954 VDD.t66 330.918
R10087 VDD.n1993 VDD.t120 330.918
R10088 VDD.n1917 VDD.t43 330.918
R10089 VDD.n2029 VDD.t98 330.918
R10090 VDD.n3790 VDD.t39 330.918
R10091 VDD.n308 VDD.t85 330.918
R10092 VDD.n3826 VDD.t59 330.918
R10093 VDD.n275 VDD.t46 330.918
R10094 VDD.n259 VDD.t101 330.918
R10095 VDD.n482 VDD.t36 330.918
R10096 VDD.n3521 VDD.t105 330.918
R10097 VDD.n3550 VDD.t50 330.918
R10098 VDD.n3455 VDD.t96 330.918
R10099 VDD.n451 VDD.t76 330.918
R10100 VDD.n3101 VDD.n774 298.538
R10101 VDD.n3422 VDD.n514 298.538
R10102 VDD.n3432 VDD.n506 298.538
R10103 VDD.n2833 VDD.n2745 298.538
R10104 VDD.n2691 VDD.n809 298.538
R10105 VDD.n2649 VDD.n2648 298.538
R10106 VDD.n1071 VDD.n1057 298.538
R10107 VDD.n2396 VDD.n1059 298.538
R10108 VDD.n3388 VDD.n3387 298.538
R10109 VDD.n3347 VDD.n3346 298.538
R10110 VDD.n3054 VDD.n2746 298.538
R10111 VDD.n3099 VDD.n2747 298.538
R10112 VDD.n2742 VDD.n798 298.538
R10113 VDD.n2698 VDD.n797 298.538
R10114 VDD.n2389 VDD.n1058 298.538
R10115 VDD.n2398 VDD.n1056 298.538
R10116 VDD.n1083 VDD.t116 246.15
R10117 VDD.n801 VDD.t71 246.15
R10118 VDD.n2053 VDD.t80 246.15
R10119 VDD.n811 VDD.t61 246.15
R10120 VDD.n2758 VDD.t87 246.15
R10121 VDD.n501 VDD.t122 246.15
R10122 VDD.n2826 VDD.t91 246.15
R10123 VDD.n537 VDD.t112 246.15
R10124 VDD.n1313 VDD.t56 223.281
R10125 VDD.n1415 VDD.t107 223.281
R10126 VDD.n1372 VDD.t69 223.281
R10127 VDD.n1448 VDD.t78 223.281
R10128 VDD.n1465 VDD.t53 223.281
R10129 VDD.n2219 VDD.t111 223.281
R10130 VDD.n1955 VDD.t67 223.281
R10131 VDD.n1994 VDD.t121 223.281
R10132 VDD.n1918 VDD.t44 223.281
R10133 VDD.n2030 VDD.t99 223.281
R10134 VDD.n3791 VDD.t40 223.281
R10135 VDD.n309 VDD.t86 223.281
R10136 VDD.n3827 VDD.t60 223.281
R10137 VDD.n276 VDD.t47 223.281
R10138 VDD.n260 VDD.t102 223.281
R10139 VDD.n483 VDD.t35 223.281
R10140 VDD.n3522 VDD.t104 223.281
R10141 VDD.n3551 VDD.t49 223.281
R10142 VDD.n3456 VDD.t95 223.281
R10143 VDD.n452 VDD.t75 223.281
R10144 VDD.n1312 VDD.t55 210.389
R10145 VDD.n1414 VDD.t106 210.389
R10146 VDD.n1371 VDD.t68 210.389
R10147 VDD.n1447 VDD.t77 210.389
R10148 VDD.n1464 VDD.t51 210.389
R10149 VDD.n2218 VDD.t109 210.389
R10150 VDD.n1954 VDD.t65 210.389
R10151 VDD.n1993 VDD.t119 210.389
R10152 VDD.n1917 VDD.t41 210.389
R10153 VDD.n2029 VDD.t97 210.389
R10154 VDD.n3790 VDD.t37 210.389
R10155 VDD.n308 VDD.t84 210.389
R10156 VDD.n3826 VDD.t58 210.389
R10157 VDD.n275 VDD.t45 210.389
R10158 VDD.n259 VDD.t100 210.389
R10159 VDD.n482 VDD.t33 210.389
R10160 VDD.n3521 VDD.t103 210.389
R10161 VDD.n3550 VDD.t48 210.389
R10162 VDD.n3455 VDD.t94 210.389
R10163 VDD.n451 VDD.t74 210.389
R10164 VDD.n1098 VDD.t26 209.835
R10165 VDD.t25 VDD.n448 209.835
R10166 VDD.n1083 VDD.t118 191.381
R10167 VDD.n801 VDD.t72 191.381
R10168 VDD.n2053 VDD.t83 191.381
R10169 VDD.n811 VDD.t63 191.381
R10170 VDD.n2758 VDD.t90 191.381
R10171 VDD.n501 VDD.t123 191.381
R10172 VDD.n2826 VDD.t93 191.381
R10173 VDD.n537 VDD.t114 191.381
R10174 VDD.n3389 VDD.n3388 185
R10175 VDD.n3388 VDD.n511 185
R10176 VDD.n3390 VDD.n512 185
R10177 VDD.n3427 VDD.n512 185
R10178 VDD.n3391 VDD.n521 185
R10179 VDD.n521 VDD.n509 185
R10180 VDD.n3393 VDD.n3392 185
R10181 VDD.n3394 VDD.n3393 185
R10182 VDD.n522 VDD.n520 185
R10183 VDD.n520 VDD.n517 185
R10184 VDD.n3326 VDD.n543 185
R10185 VDD.n3336 VDD.n543 185
R10186 VDD.n3327 VDD.n551 185
R10187 VDD.n551 VDD.n541 185
R10188 VDD.n3329 VDD.n3328 185
R10189 VDD.n3330 VDD.n3329 185
R10190 VDD.n3325 VDD.n550 185
R10191 VDD.n550 VDD.n547 185
R10192 VDD.n3324 VDD.n3323 185
R10193 VDD.n3323 VDD.n3322 185
R10194 VDD.n553 VDD.n552 185
R10195 VDD.n562 VDD.n553 185
R10196 VDD.n3315 VDD.n3314 185
R10197 VDD.n3316 VDD.n3315 185
R10198 VDD.n3313 VDD.n563 185
R10199 VDD.n563 VDD.n559 185
R10200 VDD.n3312 VDD.n3311 185
R10201 VDD.n3311 VDD.n3310 185
R10202 VDD.n565 VDD.n564 185
R10203 VDD.n566 VDD.n565 185
R10204 VDD.n3303 VDD.n3302 185
R10205 VDD.n3304 VDD.n3303 185
R10206 VDD.n3301 VDD.n575 185
R10207 VDD.n575 VDD.n572 185
R10208 VDD.n3300 VDD.n3299 185
R10209 VDD.n3299 VDD.n3298 185
R10210 VDD.n577 VDD.n576 185
R10211 VDD.n578 VDD.n577 185
R10212 VDD.n3291 VDD.n3290 185
R10213 VDD.n3292 VDD.n3291 185
R10214 VDD.n3289 VDD.n586 185
R10215 VDD.n2956 VDD.n586 185
R10216 VDD.n3288 VDD.n3287 185
R10217 VDD.n3287 VDD.n3286 185
R10218 VDD.n588 VDD.n587 185
R10219 VDD.n589 VDD.n588 185
R10220 VDD.n3279 VDD.n3278 185
R10221 VDD.n3280 VDD.n3279 185
R10222 VDD.n3277 VDD.n598 185
R10223 VDD.n598 VDD.n595 185
R10224 VDD.n3276 VDD.n3275 185
R10225 VDD.n3275 VDD.n3274 185
R10226 VDD.n600 VDD.n599 185
R10227 VDD.n601 VDD.n600 185
R10228 VDD.n3267 VDD.n3266 185
R10229 VDD.n3268 VDD.n3267 185
R10230 VDD.n3265 VDD.n610 185
R10231 VDD.n610 VDD.n607 185
R10232 VDD.n3264 VDD.n3263 185
R10233 VDD.n3263 VDD.n3262 185
R10234 VDD.n612 VDD.n611 185
R10235 VDD.n613 VDD.n612 185
R10236 VDD.n3255 VDD.n3254 185
R10237 VDD.n3256 VDD.n3255 185
R10238 VDD.n3253 VDD.n622 185
R10239 VDD.n622 VDD.n619 185
R10240 VDD.n3252 VDD.n3251 185
R10241 VDD.n3251 VDD.n3250 185
R10242 VDD.n624 VDD.n623 185
R10243 VDD.n625 VDD.n624 185
R10244 VDD.n3243 VDD.n3242 185
R10245 VDD.n3244 VDD.n3243 185
R10246 VDD.n3241 VDD.n634 185
R10247 VDD.n634 VDD.n631 185
R10248 VDD.n3240 VDD.n3239 185
R10249 VDD.n3239 VDD.n3238 185
R10250 VDD.n636 VDD.n635 185
R10251 VDD.n637 VDD.n636 185
R10252 VDD.n3231 VDD.n3230 185
R10253 VDD.n3232 VDD.n3231 185
R10254 VDD.n3229 VDD.n646 185
R10255 VDD.n646 VDD.n643 185
R10256 VDD.n3228 VDD.n3227 185
R10257 VDD.n3227 VDD.n3226 185
R10258 VDD.n648 VDD.n647 185
R10259 VDD.n657 VDD.n648 185
R10260 VDD.n3219 VDD.n3218 185
R10261 VDD.n3220 VDD.n3219 185
R10262 VDD.n3217 VDD.n658 185
R10263 VDD.n658 VDD.n654 185
R10264 VDD.n3216 VDD.n3215 185
R10265 VDD.n3215 VDD.n3214 185
R10266 VDD.n660 VDD.n659 185
R10267 VDD.n661 VDD.n660 185
R10268 VDD.n3207 VDD.n3206 185
R10269 VDD.n3208 VDD.n3207 185
R10270 VDD.n3205 VDD.n670 185
R10271 VDD.n670 VDD.n667 185
R10272 VDD.n3204 VDD.n3203 185
R10273 VDD.n3203 VDD.n3202 185
R10274 VDD.n672 VDD.n671 185
R10275 VDD.n673 VDD.n672 185
R10276 VDD.n3195 VDD.n3194 185
R10277 VDD.n3196 VDD.n3195 185
R10278 VDD.n3193 VDD.n682 185
R10279 VDD.n682 VDD.n679 185
R10280 VDD.n3192 VDD.n3191 185
R10281 VDD.n3191 VDD.n3190 185
R10282 VDD.n684 VDD.n683 185
R10283 VDD.n685 VDD.n684 185
R10284 VDD.n3183 VDD.n3182 185
R10285 VDD.n3184 VDD.n3183 185
R10286 VDD.n3181 VDD.n694 185
R10287 VDD.n694 VDD.n691 185
R10288 VDD.n3180 VDD.n3179 185
R10289 VDD.n3179 VDD.n3178 185
R10290 VDD.n696 VDD.n695 185
R10291 VDD.n705 VDD.n696 185
R10292 VDD.n3171 VDD.n3170 185
R10293 VDD.n3172 VDD.n3171 185
R10294 VDD.n3169 VDD.n706 185
R10295 VDD.n706 VDD.n702 185
R10296 VDD.n3168 VDD.n3167 185
R10297 VDD.n3167 VDD.n3166 185
R10298 VDD.n708 VDD.n707 185
R10299 VDD.n709 VDD.n708 185
R10300 VDD.n3159 VDD.n3158 185
R10301 VDD.n3160 VDD.n3159 185
R10302 VDD.n3157 VDD.n718 185
R10303 VDD.n718 VDD.n715 185
R10304 VDD.n3156 VDD.n3155 185
R10305 VDD.n3155 VDD.n3154 185
R10306 VDD.n720 VDD.n719 185
R10307 VDD.n721 VDD.n720 185
R10308 VDD.n3147 VDD.n3146 185
R10309 VDD.n3148 VDD.n3147 185
R10310 VDD.n3145 VDD.n730 185
R10311 VDD.n730 VDD.n727 185
R10312 VDD.n3144 VDD.n3143 185
R10313 VDD.n3143 VDD.n3142 185
R10314 VDD.n732 VDD.n731 185
R10315 VDD.n733 VDD.n732 185
R10316 VDD.n3135 VDD.n3134 185
R10317 VDD.n3136 VDD.n3135 185
R10318 VDD.n3133 VDD.n742 185
R10319 VDD.n742 VDD.n739 185
R10320 VDD.n3132 VDD.n3131 185
R10321 VDD.n3131 VDD.n3130 185
R10322 VDD.n744 VDD.n743 185
R10323 VDD.n745 VDD.n744 185
R10324 VDD.n3123 VDD.n3122 185
R10325 VDD.n3124 VDD.n3123 185
R10326 VDD.n3121 VDD.n754 185
R10327 VDD.n754 VDD.n751 185
R10328 VDD.n3120 VDD.n3119 185
R10329 VDD.n3119 VDD.n3118 185
R10330 VDD.n756 VDD.n755 185
R10331 VDD.n757 VDD.n756 185
R10332 VDD.n3111 VDD.n3110 185
R10333 VDD.n3112 VDD.n3111 185
R10334 VDD.n3109 VDD.n766 185
R10335 VDD.n766 VDD.n763 185
R10336 VDD.n3108 VDD.n3107 185
R10337 VDD.n3107 VDD.n3106 185
R10338 VDD.n768 VDD.n767 185
R10339 VDD.n769 VDD.n768 185
R10340 VDD.n3099 VDD.n3098 185
R10341 VDD.n3100 VDD.n3099 185
R10342 VDD.n3097 VDD.n2747 185
R10343 VDD.n3096 VDD.n3095 185
R10344 VDD.n3093 VDD.n2748 185
R10345 VDD.n3091 VDD.n3090 185
R10346 VDD.n3089 VDD.n2749 185
R10347 VDD.n3088 VDD.n3087 185
R10348 VDD.n3085 VDD.n2750 185
R10349 VDD.n3083 VDD.n3082 185
R10350 VDD.n3081 VDD.n2751 185
R10351 VDD.n3080 VDD.n3079 185
R10352 VDD.n3077 VDD.n2752 185
R10353 VDD.n3075 VDD.n3074 185
R10354 VDD.n3073 VDD.n2753 185
R10355 VDD.n3072 VDD.n3071 185
R10356 VDD.n3069 VDD.n2754 185
R10357 VDD.n3067 VDD.n3066 185
R10358 VDD.n3065 VDD.n2755 185
R10359 VDD.n3064 VDD.n3063 185
R10360 VDD.n3061 VDD.n2756 185
R10361 VDD.n3059 VDD.n3058 185
R10362 VDD.n3056 VDD.n2757 185
R10363 VDD.n3055 VDD.n3054 185
R10364 VDD.n3348 VDD.n3347 185
R10365 VDD.n3349 VDD.n536 185
R10366 VDD.n3352 VDD.n3351 185
R10367 VDD.n3354 VDD.n534 185
R10368 VDD.n3356 VDD.n3355 185
R10369 VDD.n3357 VDD.n533 185
R10370 VDD.n3359 VDD.n3358 185
R10371 VDD.n3361 VDD.n531 185
R10372 VDD.n3363 VDD.n3362 185
R10373 VDD.n3364 VDD.n530 185
R10374 VDD.n3366 VDD.n3365 185
R10375 VDD.n3369 VDD.n3368 185
R10376 VDD.n3371 VDD.n3370 185
R10377 VDD.n3373 VDD.n528 185
R10378 VDD.n3375 VDD.n3374 185
R10379 VDD.n3376 VDD.n527 185
R10380 VDD.n3378 VDD.n3377 185
R10381 VDD.n3380 VDD.n525 185
R10382 VDD.n3382 VDD.n3381 185
R10383 VDD.n3383 VDD.n524 185
R10384 VDD.n3385 VDD.n3384 185
R10385 VDD.n3387 VDD.n523 185
R10386 VDD.n3346 VDD.n3344 185
R10387 VDD.n3346 VDD.n511 185
R10388 VDD.n3343 VDD.n510 185
R10389 VDD.n3427 VDD.n510 185
R10390 VDD.n3342 VDD.n3341 185
R10391 VDD.n3341 VDD.n509 185
R10392 VDD.n3340 VDD.n519 185
R10393 VDD.n3394 VDD.n519 185
R10394 VDD.n3339 VDD.n3338 185
R10395 VDD.n3338 VDD.n517 185
R10396 VDD.n3337 VDD.n539 185
R10397 VDD.n3337 VDD.n3336 185
R10398 VDD.n2760 VDD.n540 185
R10399 VDD.n541 VDD.n540 185
R10400 VDD.n2761 VDD.n549 185
R10401 VDD.n3330 VDD.n549 185
R10402 VDD.n2763 VDD.n2762 185
R10403 VDD.n2762 VDD.n547 185
R10404 VDD.n2764 VDD.n555 185
R10405 VDD.n3322 VDD.n555 185
R10406 VDD.n2766 VDD.n2765 185
R10407 VDD.n2765 VDD.n562 185
R10408 VDD.n2767 VDD.n561 185
R10409 VDD.n3316 VDD.n561 185
R10410 VDD.n2769 VDD.n2768 185
R10411 VDD.n2768 VDD.n559 185
R10412 VDD.n2770 VDD.n568 185
R10413 VDD.n3310 VDD.n568 185
R10414 VDD.n2772 VDD.n2771 185
R10415 VDD.n2771 VDD.n566 185
R10416 VDD.n2773 VDD.n574 185
R10417 VDD.n3304 VDD.n574 185
R10418 VDD.n2775 VDD.n2774 185
R10419 VDD.n2774 VDD.n572 185
R10420 VDD.n2776 VDD.n580 185
R10421 VDD.n3298 VDD.n580 185
R10422 VDD.n2778 VDD.n2777 185
R10423 VDD.n2777 VDD.n578 185
R10424 VDD.n2779 VDD.n585 185
R10425 VDD.n3292 VDD.n585 185
R10426 VDD.n2958 VDD.n2957 185
R10427 VDD.n2957 VDD.n2956 185
R10428 VDD.n2959 VDD.n591 185
R10429 VDD.n3286 VDD.n591 185
R10430 VDD.n2961 VDD.n2960 185
R10431 VDD.n2960 VDD.n589 185
R10432 VDD.n2962 VDD.n597 185
R10433 VDD.n3280 VDD.n597 185
R10434 VDD.n2964 VDD.n2963 185
R10435 VDD.n2963 VDD.n595 185
R10436 VDD.n2965 VDD.n603 185
R10437 VDD.n3274 VDD.n603 185
R10438 VDD.n2967 VDD.n2966 185
R10439 VDD.n2966 VDD.n601 185
R10440 VDD.n2968 VDD.n609 185
R10441 VDD.n3268 VDD.n609 185
R10442 VDD.n2970 VDD.n2969 185
R10443 VDD.n2969 VDD.n607 185
R10444 VDD.n2971 VDD.n615 185
R10445 VDD.n3262 VDD.n615 185
R10446 VDD.n2973 VDD.n2972 185
R10447 VDD.n2972 VDD.n613 185
R10448 VDD.n2974 VDD.n621 185
R10449 VDD.n3256 VDD.n621 185
R10450 VDD.n2976 VDD.n2975 185
R10451 VDD.n2975 VDD.n619 185
R10452 VDD.n2977 VDD.n627 185
R10453 VDD.n3250 VDD.n627 185
R10454 VDD.n2979 VDD.n2978 185
R10455 VDD.n2978 VDD.n625 185
R10456 VDD.n2980 VDD.n633 185
R10457 VDD.n3244 VDD.n633 185
R10458 VDD.n2982 VDD.n2981 185
R10459 VDD.n2981 VDD.n631 185
R10460 VDD.n2983 VDD.n639 185
R10461 VDD.n3238 VDD.n639 185
R10462 VDD.n2985 VDD.n2984 185
R10463 VDD.n2984 VDD.n637 185
R10464 VDD.n2986 VDD.n645 185
R10465 VDD.n3232 VDD.n645 185
R10466 VDD.n2988 VDD.n2987 185
R10467 VDD.n2987 VDD.n643 185
R10468 VDD.n2989 VDD.n650 185
R10469 VDD.n3226 VDD.n650 185
R10470 VDD.n2991 VDD.n2990 185
R10471 VDD.n2990 VDD.n657 185
R10472 VDD.n2992 VDD.n656 185
R10473 VDD.n3220 VDD.n656 185
R10474 VDD.n2994 VDD.n2993 185
R10475 VDD.n2993 VDD.n654 185
R10476 VDD.n2995 VDD.n663 185
R10477 VDD.n3214 VDD.n663 185
R10478 VDD.n2997 VDD.n2996 185
R10479 VDD.n2996 VDD.n661 185
R10480 VDD.n2998 VDD.n669 185
R10481 VDD.n3208 VDD.n669 185
R10482 VDD.n3000 VDD.n2999 185
R10483 VDD.n2999 VDD.n667 185
R10484 VDD.n3001 VDD.n675 185
R10485 VDD.n3202 VDD.n675 185
R10486 VDD.n3003 VDD.n3002 185
R10487 VDD.n3002 VDD.n673 185
R10488 VDD.n3004 VDD.n681 185
R10489 VDD.n3196 VDD.n681 185
R10490 VDD.n3006 VDD.n3005 185
R10491 VDD.n3005 VDD.n679 185
R10492 VDD.n3007 VDD.n687 185
R10493 VDD.n3190 VDD.n687 185
R10494 VDD.n3009 VDD.n3008 185
R10495 VDD.n3008 VDD.n685 185
R10496 VDD.n3010 VDD.n693 185
R10497 VDD.n3184 VDD.n693 185
R10498 VDD.n3012 VDD.n3011 185
R10499 VDD.n3011 VDD.n691 185
R10500 VDD.n3013 VDD.n698 185
R10501 VDD.n3178 VDD.n698 185
R10502 VDD.n3015 VDD.n3014 185
R10503 VDD.n3014 VDD.n705 185
R10504 VDD.n3016 VDD.n704 185
R10505 VDD.n3172 VDD.n704 185
R10506 VDD.n3018 VDD.n3017 185
R10507 VDD.n3017 VDD.n702 185
R10508 VDD.n3019 VDD.n711 185
R10509 VDD.n3166 VDD.n711 185
R10510 VDD.n3021 VDD.n3020 185
R10511 VDD.n3020 VDD.n709 185
R10512 VDD.n3022 VDD.n717 185
R10513 VDD.n3160 VDD.n717 185
R10514 VDD.n3024 VDD.n3023 185
R10515 VDD.n3023 VDD.n715 185
R10516 VDD.n3025 VDD.n723 185
R10517 VDD.n3154 VDD.n723 185
R10518 VDD.n3027 VDD.n3026 185
R10519 VDD.n3026 VDD.n721 185
R10520 VDD.n3028 VDD.n729 185
R10521 VDD.n3148 VDD.n729 185
R10522 VDD.n3030 VDD.n3029 185
R10523 VDD.n3029 VDD.n727 185
R10524 VDD.n3031 VDD.n735 185
R10525 VDD.n3142 VDD.n735 185
R10526 VDD.n3033 VDD.n3032 185
R10527 VDD.n3032 VDD.n733 185
R10528 VDD.n3034 VDD.n741 185
R10529 VDD.n3136 VDD.n741 185
R10530 VDD.n3036 VDD.n3035 185
R10531 VDD.n3035 VDD.n739 185
R10532 VDD.n3037 VDD.n747 185
R10533 VDD.n3130 VDD.n747 185
R10534 VDD.n3039 VDD.n3038 185
R10535 VDD.n3038 VDD.n745 185
R10536 VDD.n3040 VDD.n753 185
R10537 VDD.n3124 VDD.n753 185
R10538 VDD.n3042 VDD.n3041 185
R10539 VDD.n3041 VDD.n751 185
R10540 VDD.n3043 VDD.n759 185
R10541 VDD.n3118 VDD.n759 185
R10542 VDD.n3045 VDD.n3044 185
R10543 VDD.n3044 VDD.n757 185
R10544 VDD.n3046 VDD.n765 185
R10545 VDD.n3112 VDD.n765 185
R10546 VDD.n3048 VDD.n3047 185
R10547 VDD.n3047 VDD.n763 185
R10548 VDD.n3049 VDD.n771 185
R10549 VDD.n3106 VDD.n771 185
R10550 VDD.n3051 VDD.n3050 185
R10551 VDD.n3050 VDD.n769 185
R10552 VDD.n3052 VDD.n2746 185
R10553 VDD.n3100 VDD.n2746 185
R10554 VDD.n2211 VDD.n2210 185
R10555 VDD.n2212 VDD.n2211 185
R10556 VDD.n1101 VDD.n1099 185
R10557 VDD.n1099 VDD.n1096 185
R10558 VDD.n1894 VDD.n1893 185
R10559 VDD.n1893 VDD.n1892 185
R10560 VDD.n1104 VDD.n1103 185
R10561 VDD.n1105 VDD.n1104 185
R10562 VDD.n1883 VDD.n1882 185
R10563 VDD.n1884 VDD.n1883 185
R10564 VDD.n1113 VDD.n1112 185
R10565 VDD.n1112 VDD.n1111 185
R10566 VDD.n1878 VDD.n1877 185
R10567 VDD.n1877 VDD.n1876 185
R10568 VDD.n1116 VDD.n1115 185
R10569 VDD.n1117 VDD.n1116 185
R10570 VDD.n1867 VDD.n1866 185
R10571 VDD.n1868 VDD.n1867 185
R10572 VDD.n1125 VDD.n1124 185
R10573 VDD.n1124 VDD.n1123 185
R10574 VDD.n1862 VDD.n1861 185
R10575 VDD.n1861 VDD.n1860 185
R10576 VDD.n1128 VDD.n1127 185
R10577 VDD.n1129 VDD.n1128 185
R10578 VDD.n1851 VDD.n1850 185
R10579 VDD.n1852 VDD.n1851 185
R10580 VDD.n1137 VDD.n1136 185
R10581 VDD.n1136 VDD.n1135 185
R10582 VDD.n1846 VDD.n1845 185
R10583 VDD.n1845 VDD.n1844 185
R10584 VDD.n1140 VDD.n1139 185
R10585 VDD.n1141 VDD.n1140 185
R10586 VDD.n1835 VDD.n1834 185
R10587 VDD.n1836 VDD.n1835 185
R10588 VDD.n1149 VDD.n1148 185
R10589 VDD.n1148 VDD.n1147 185
R10590 VDD.n1830 VDD.n1829 185
R10591 VDD.n1829 VDD.n1828 185
R10592 VDD.n1152 VDD.n1151 185
R10593 VDD.n1159 VDD.n1152 185
R10594 VDD.n1819 VDD.n1818 185
R10595 VDD.n1820 VDD.n1819 185
R10596 VDD.n1161 VDD.n1160 185
R10597 VDD.n1160 VDD.n1158 185
R10598 VDD.n1814 VDD.n1813 185
R10599 VDD.n1813 VDD.n1812 185
R10600 VDD.n1164 VDD.n1163 185
R10601 VDD.n1165 VDD.n1164 185
R10602 VDD.n1803 VDD.n1802 185
R10603 VDD.n1804 VDD.n1803 185
R10604 VDD.n1173 VDD.n1172 185
R10605 VDD.n1172 VDD.n1171 185
R10606 VDD.n1798 VDD.n1797 185
R10607 VDD.n1797 VDD.n1796 185
R10608 VDD.n1176 VDD.n1175 185
R10609 VDD.n1177 VDD.n1176 185
R10610 VDD.n1787 VDD.n1786 185
R10611 VDD.n1788 VDD.n1787 185
R10612 VDD.n1185 VDD.n1184 185
R10613 VDD.n1184 VDD.n1183 185
R10614 VDD.n1782 VDD.n1781 185
R10615 VDD.n1781 VDD.n1780 185
R10616 VDD.n1188 VDD.n1187 185
R10617 VDD.n1189 VDD.n1188 185
R10618 VDD.n1771 VDD.n1770 185
R10619 VDD.n1772 VDD.n1771 185
R10620 VDD.n1197 VDD.n1196 185
R10621 VDD.n1196 VDD.n1195 185
R10622 VDD.n1766 VDD.n1765 185
R10623 VDD.n1765 VDD.n1764 185
R10624 VDD.n1200 VDD.n1199 185
R10625 VDD.n1201 VDD.n1200 185
R10626 VDD.n1755 VDD.n1754 185
R10627 VDD.n1756 VDD.n1755 185
R10628 VDD.n1209 VDD.n1208 185
R10629 VDD.n1208 VDD.n1207 185
R10630 VDD.n1619 VDD.n1618 185
R10631 VDD.n1618 VDD.n1617 185
R10632 VDD.n1212 VDD.n1211 185
R10633 VDD.n1213 VDD.n1212 185
R10634 VDD.n1608 VDD.n1607 185
R10635 VDD.n1609 VDD.n1608 185
R10636 VDD.n1221 VDD.n1220 185
R10637 VDD.n1220 VDD.n1219 185
R10638 VDD.n1603 VDD.n1602 185
R10639 VDD.n1602 VDD.n1601 185
R10640 VDD.n1224 VDD.n1223 185
R10641 VDD.n1225 VDD.n1224 185
R10642 VDD.n1592 VDD.n1591 185
R10643 VDD.n1593 VDD.n1592 185
R10644 VDD.n1233 VDD.n1232 185
R10645 VDD.n1232 VDD.n1231 185
R10646 VDD.n1587 VDD.n1586 185
R10647 VDD.n1586 VDD.n1585 185
R10648 VDD.n1236 VDD.n1235 185
R10649 VDD.n1237 VDD.n1236 185
R10650 VDD.n1576 VDD.n1575 185
R10651 VDD.n1577 VDD.n1576 185
R10652 VDD.n1245 VDD.n1244 185
R10653 VDD.n1244 VDD.n1243 185
R10654 VDD.n1571 VDD.n1570 185
R10655 VDD.n1570 VDD.n1569 185
R10656 VDD.n1248 VDD.n1247 185
R10657 VDD.n1249 VDD.n1248 185
R10658 VDD.n1560 VDD.n1559 185
R10659 VDD.n1561 VDD.n1560 185
R10660 VDD.n1256 VDD.n1255 185
R10661 VDD.n1552 VDD.n1255 185
R10662 VDD.n1555 VDD.n1554 185
R10663 VDD.n1554 VDD.n1553 185
R10664 VDD.n1259 VDD.n1258 185
R10665 VDD.n1260 VDD.n1259 185
R10666 VDD.n1543 VDD.n1542 185
R10667 VDD.n1544 VDD.n1543 185
R10668 VDD.n1268 VDD.n1267 185
R10669 VDD.n1267 VDD.n1266 185
R10670 VDD.n1538 VDD.n1537 185
R10671 VDD.n1537 VDD.n1536 185
R10672 VDD.n1271 VDD.n1270 185
R10673 VDD.n1272 VDD.n1271 185
R10674 VDD.n1527 VDD.n1526 185
R10675 VDD.n1528 VDD.n1527 185
R10676 VDD.n1280 VDD.n1279 185
R10677 VDD.n1279 VDD.n1278 185
R10678 VDD.n1522 VDD.n1521 185
R10679 VDD.n1521 VDD.n1520 185
R10680 VDD.n1283 VDD.n1282 185
R10681 VDD.n1284 VDD.n1283 185
R10682 VDD.n1511 VDD.n1510 185
R10683 VDD.n1512 VDD.n1511 185
R10684 VDD.n1292 VDD.n1291 185
R10685 VDD.n1291 VDD.n1290 185
R10686 VDD.n1506 VDD.n1505 185
R10687 VDD.n1505 VDD.n1504 185
R10688 VDD.n1295 VDD.n1294 185
R10689 VDD.n1296 VDD.n1295 185
R10690 VDD.n1495 VDD.n1494 185
R10691 VDD.n1496 VDD.n1495 185
R10692 VDD.n1304 VDD.n1303 185
R10693 VDD.n1303 VDD.n1302 185
R10694 VDD.n1490 VDD.n1489 185
R10695 VDD.n1489 VDD.n1488 185
R10696 VDD.n1307 VDD.n1306 185
R10697 VDD.n1308 VDD.n1307 185
R10698 VDD.n1478 VDD.n1477 185
R10699 VDD.n1476 VDD.n1338 185
R10700 VDD.n1340 VDD.n1337 185
R10701 VDD.n1480 VDD.n1337 185
R10702 VDD.n1472 VDD.n1342 185
R10703 VDD.n1471 VDD.n1343 185
R10704 VDD.n1470 VDD.n1344 185
R10705 VDD.n1462 VDD.n1345 185
R10706 VDD.n1466 VDD.n1463 185
R10707 VDD.n1461 VDD.n1347 185
R10708 VDD.n1460 VDD.n1348 185
R10709 VDD.n1351 VDD.n1349 185
R10710 VDD.n1456 VDD.n1352 185
R10711 VDD.n1455 VDD.n1353 185
R10712 VDD.n1454 VDD.n1354 185
R10713 VDD.n1357 VDD.n1355 185
R10714 VDD.n1450 VDD.n1358 185
R10715 VDD.n1449 VDD.n1446 185
R10716 VDD.n1445 VDD.n1444 185
R10717 VDD.n1361 VDD.n1359 185
R10718 VDD.n1440 VDD.n1362 185
R10719 VDD.n1439 VDD.n1363 185
R10720 VDD.n1438 VDD.n1364 185
R10721 VDD.n1367 VDD.n1365 185
R10722 VDD.n1434 VDD.n1368 185
R10723 VDD.n1433 VDD.n1369 185
R10724 VDD.n1432 VDD.n1370 185
R10725 VDD.n1429 VDD.n1375 185
R10726 VDD.n1428 VDD.n1376 185
R10727 VDD.n1427 VDD.n1377 185
R10728 VDD.n1379 VDD.n1378 185
R10729 VDD.n1423 VDD.n1381 185
R10730 VDD.n1422 VDD.n1382 185
R10731 VDD.n1421 VDD.n1383 185
R10732 VDD.n1385 VDD.n1384 185
R10733 VDD.n1417 VDD.n1387 185
R10734 VDD.n1416 VDD.n1413 185
R10735 VDD.n1412 VDD.n1388 185
R10736 VDD.n1390 VDD.n1389 185
R10737 VDD.n1408 VDD.n1392 185
R10738 VDD.n1407 VDD.n1393 185
R10739 VDD.n1406 VDD.n1394 185
R10740 VDD.n1396 VDD.n1395 185
R10741 VDD.n1402 VDD.n1398 185
R10742 VDD.n1401 VDD.n1399 185
R10743 VDD.n1400 VDD.n1315 185
R10744 VDD.n1482 VDD.n1481 185
R10745 VDD.n1481 VDD.n1480 185
R10746 VDD.n2217 VDD.n1092 185
R10747 VDD.n2221 VDD.n1091 185
R10748 VDD.n2222 VDD.n1090 185
R10749 VDD.n1963 VDD.n1089 185
R10750 VDD.n1965 VDD.n1964 185
R10751 VDD.n1967 VDD.n1961 185
R10752 VDD.n1969 VDD.n1968 185
R10753 VDD.n1971 VDD.n1958 185
R10754 VDD.n1973 VDD.n1972 185
R10755 VDD.n1959 VDD.n1953 185
R10756 VDD.n1977 VDD.n1957 185
R10757 VDD.n1978 VDD.n1949 185
R10758 VDD.n1980 VDD.n1979 185
R10759 VDD.n1982 VDD.n1947 185
R10760 VDD.n1984 VDD.n1983 185
R10761 VDD.n1985 VDD.n1942 185
R10762 VDD.n1987 VDD.n1986 185
R10763 VDD.n1989 VDD.n1940 185
R10764 VDD.n1991 VDD.n1990 185
R10765 VDD.n1992 VDD.n1935 185
R10766 VDD.n1997 VDD.n1996 185
R10767 VDD.n1999 VDD.n1933 185
R10768 VDD.n2001 VDD.n2000 185
R10769 VDD.n2002 VDD.n1928 185
R10770 VDD.n2004 VDD.n2003 185
R10771 VDD.n2006 VDD.n1926 185
R10772 VDD.n2008 VDD.n2007 185
R10773 VDD.n2009 VDD.n1921 185
R10774 VDD.n2011 VDD.n2010 185
R10775 VDD.n2013 VDD.n1919 185
R10776 VDD.n2015 VDD.n2014 185
R10777 VDD.n2016 VDD.n1912 185
R10778 VDD.n2018 VDD.n2017 185
R10779 VDD.n2020 VDD.n1911 185
R10780 VDD.n2021 VDD.n1908 185
R10781 VDD.n2024 VDD.n2023 185
R10782 VDD.n1910 VDD.n1906 185
R10783 VDD.n2028 VDD.n1905 185
R10784 VDD.n2032 VDD.n2031 185
R10785 VDD.n2034 VDD.n1903 185
R10786 VDD.n2036 VDD.n2035 185
R10787 VDD.n1901 VDD.n1900 185
R10788 VDD.n2202 VDD.n2201 185
R10789 VDD.n2204 VDD.n1898 185
R10790 VDD.n2206 VDD.n2205 185
R10791 VDD.n2207 VDD.n1100 185
R10792 VDD.n2214 VDD.n2213 185
R10793 VDD.n2213 VDD.n2212 185
R10794 VDD.n1095 VDD.n1094 185
R10795 VDD.n1096 VDD.n1095 185
R10796 VDD.n1891 VDD.n1890 185
R10797 VDD.n1892 VDD.n1891 185
R10798 VDD.n1107 VDD.n1106 185
R10799 VDD.n1106 VDD.n1105 185
R10800 VDD.n1886 VDD.n1885 185
R10801 VDD.n1885 VDD.n1884 185
R10802 VDD.n1110 VDD.n1109 185
R10803 VDD.n1111 VDD.n1110 185
R10804 VDD.n1875 VDD.n1874 185
R10805 VDD.n1876 VDD.n1875 185
R10806 VDD.n1119 VDD.n1118 185
R10807 VDD.n1118 VDD.n1117 185
R10808 VDD.n1870 VDD.n1869 185
R10809 VDD.n1869 VDD.n1868 185
R10810 VDD.n1122 VDD.n1121 185
R10811 VDD.n1123 VDD.n1122 185
R10812 VDD.n1859 VDD.n1858 185
R10813 VDD.n1860 VDD.n1859 185
R10814 VDD.n1131 VDD.n1130 185
R10815 VDD.n1130 VDD.n1129 185
R10816 VDD.n1854 VDD.n1853 185
R10817 VDD.n1853 VDD.n1852 185
R10818 VDD.n1134 VDD.n1133 185
R10819 VDD.n1135 VDD.n1134 185
R10820 VDD.n1843 VDD.n1842 185
R10821 VDD.n1844 VDD.n1843 185
R10822 VDD.n1143 VDD.n1142 185
R10823 VDD.n1142 VDD.n1141 185
R10824 VDD.n1838 VDD.n1837 185
R10825 VDD.n1837 VDD.n1836 185
R10826 VDD.n1146 VDD.n1145 185
R10827 VDD.n1147 VDD.n1146 185
R10828 VDD.n1827 VDD.n1826 185
R10829 VDD.n1828 VDD.n1827 185
R10830 VDD.n1154 VDD.n1153 185
R10831 VDD.n1159 VDD.n1153 185
R10832 VDD.n1822 VDD.n1821 185
R10833 VDD.n1821 VDD.n1820 185
R10834 VDD.n1157 VDD.n1156 185
R10835 VDD.n1158 VDD.n1157 185
R10836 VDD.n1811 VDD.n1810 185
R10837 VDD.n1812 VDD.n1811 185
R10838 VDD.n1167 VDD.n1166 185
R10839 VDD.n1166 VDD.n1165 185
R10840 VDD.n1806 VDD.n1805 185
R10841 VDD.n1805 VDD.n1804 185
R10842 VDD.n1170 VDD.n1169 185
R10843 VDD.n1171 VDD.n1170 185
R10844 VDD.n1795 VDD.n1794 185
R10845 VDD.n1796 VDD.n1795 185
R10846 VDD.n1179 VDD.n1178 185
R10847 VDD.n1178 VDD.n1177 185
R10848 VDD.n1790 VDD.n1789 185
R10849 VDD.n1789 VDD.n1788 185
R10850 VDD.n1182 VDD.n1181 185
R10851 VDD.n1183 VDD.n1182 185
R10852 VDD.n1779 VDD.n1778 185
R10853 VDD.n1780 VDD.n1779 185
R10854 VDD.n1191 VDD.n1190 185
R10855 VDD.n1190 VDD.n1189 185
R10856 VDD.n1774 VDD.n1773 185
R10857 VDD.n1773 VDD.n1772 185
R10858 VDD.n1194 VDD.n1193 185
R10859 VDD.n1195 VDD.n1194 185
R10860 VDD.n1763 VDD.n1762 185
R10861 VDD.n1764 VDD.n1763 185
R10862 VDD.n1203 VDD.n1202 185
R10863 VDD.n1202 VDD.n1201 185
R10864 VDD.n1758 VDD.n1757 185
R10865 VDD.n1757 VDD.n1756 185
R10866 VDD.n1206 VDD.n1205 185
R10867 VDD.n1207 VDD.n1206 185
R10868 VDD.n1616 VDD.n1615 185
R10869 VDD.n1617 VDD.n1616 185
R10870 VDD.n1215 VDD.n1214 185
R10871 VDD.n1214 VDD.n1213 185
R10872 VDD.n1611 VDD.n1610 185
R10873 VDD.n1610 VDD.n1609 185
R10874 VDD.n1218 VDD.n1217 185
R10875 VDD.n1219 VDD.n1218 185
R10876 VDD.n1600 VDD.n1599 185
R10877 VDD.n1601 VDD.n1600 185
R10878 VDD.n1227 VDD.n1226 185
R10879 VDD.n1226 VDD.n1225 185
R10880 VDD.n1595 VDD.n1594 185
R10881 VDD.n1594 VDD.n1593 185
R10882 VDD.n1230 VDD.n1229 185
R10883 VDD.n1231 VDD.n1230 185
R10884 VDD.n1584 VDD.n1583 185
R10885 VDD.n1585 VDD.n1584 185
R10886 VDD.n1239 VDD.n1238 185
R10887 VDD.n1238 VDD.n1237 185
R10888 VDD.n1579 VDD.n1578 185
R10889 VDD.n1578 VDD.n1577 185
R10890 VDD.n1242 VDD.n1241 185
R10891 VDD.n1243 VDD.n1242 185
R10892 VDD.n1568 VDD.n1567 185
R10893 VDD.n1569 VDD.n1568 185
R10894 VDD.n1251 VDD.n1250 185
R10895 VDD.n1250 VDD.n1249 185
R10896 VDD.n1563 VDD.n1562 185
R10897 VDD.n1562 VDD.n1561 185
R10898 VDD.n1254 VDD.n1253 185
R10899 VDD.n1552 VDD.n1254 185
R10900 VDD.n1551 VDD.n1550 185
R10901 VDD.n1553 VDD.n1551 185
R10902 VDD.n1262 VDD.n1261 185
R10903 VDD.n1261 VDD.n1260 185
R10904 VDD.n1546 VDD.n1545 185
R10905 VDD.n1545 VDD.n1544 185
R10906 VDD.n1265 VDD.n1264 185
R10907 VDD.n1266 VDD.n1265 185
R10908 VDD.n1535 VDD.n1534 185
R10909 VDD.n1536 VDD.n1535 185
R10910 VDD.n1274 VDD.n1273 185
R10911 VDD.n1273 VDD.n1272 185
R10912 VDD.n1530 VDD.n1529 185
R10913 VDD.n1529 VDD.n1528 185
R10914 VDD.n1277 VDD.n1276 185
R10915 VDD.n1278 VDD.n1277 185
R10916 VDD.n1519 VDD.n1518 185
R10917 VDD.n1520 VDD.n1519 185
R10918 VDD.n1286 VDD.n1285 185
R10919 VDD.n1285 VDD.n1284 185
R10920 VDD.n1514 VDD.n1513 185
R10921 VDD.n1513 VDD.n1512 185
R10922 VDD.n1289 VDD.n1288 185
R10923 VDD.n1290 VDD.n1289 185
R10924 VDD.n1503 VDD.n1502 185
R10925 VDD.n1504 VDD.n1503 185
R10926 VDD.n1298 VDD.n1297 185
R10927 VDD.n1297 VDD.n1296 185
R10928 VDD.n1498 VDD.n1497 185
R10929 VDD.n1497 VDD.n1496 185
R10930 VDD.n1301 VDD.n1300 185
R10931 VDD.n1302 VDD.n1301 185
R10932 VDD.n1487 VDD.n1486 185
R10933 VDD.n1488 VDD.n1487 185
R10934 VDD.n1310 VDD.n1309 185
R10935 VDD.n1309 VDD.n1308 185
R10936 VDD.n2693 VDD.n809 185
R10937 VDD.n809 VDD.n775 185
R10938 VDD.n2695 VDD.n2694 185
R10939 VDD.n2696 VDD.n2695 185
R10940 VDD.n810 VDD.n808 185
R10941 VDD.n808 VDD.n805 185
R10942 VDD.n2641 VDD.n2640 185
R10943 VDD.n2642 VDD.n2641 185
R10944 VDD.n2639 VDD.n819 185
R10945 VDD.n819 VDD.n816 185
R10946 VDD.n2638 VDD.n2637 185
R10947 VDD.n2637 VDD.n2636 185
R10948 VDD.n821 VDD.n820 185
R10949 VDD.n822 VDD.n821 185
R10950 VDD.n2624 VDD.n2623 185
R10951 VDD.n2625 VDD.n2624 185
R10952 VDD.n2622 VDD.n832 185
R10953 VDD.n832 VDD.n829 185
R10954 VDD.n2621 VDD.n2620 185
R10955 VDD.n2620 VDD.n2619 185
R10956 VDD.n834 VDD.n833 185
R10957 VDD.n835 VDD.n834 185
R10958 VDD.n2612 VDD.n2611 185
R10959 VDD.n2613 VDD.n2612 185
R10960 VDD.n2610 VDD.n844 185
R10961 VDD.n844 VDD.n841 185
R10962 VDD.n2609 VDD.n2608 185
R10963 VDD.n2608 VDD.n2607 185
R10964 VDD.n846 VDD.n845 185
R10965 VDD.n847 VDD.n846 185
R10966 VDD.n2600 VDD.n2599 185
R10967 VDD.n2601 VDD.n2600 185
R10968 VDD.n2598 VDD.n856 185
R10969 VDD.n856 VDD.n853 185
R10970 VDD.n2597 VDD.n2596 185
R10971 VDD.n2596 VDD.n2595 185
R10972 VDD.n858 VDD.n857 185
R10973 VDD.n859 VDD.n858 185
R10974 VDD.n2588 VDD.n2587 185
R10975 VDD.n2589 VDD.n2588 185
R10976 VDD.n2586 VDD.n868 185
R10977 VDD.n868 VDD.n865 185
R10978 VDD.n2585 VDD.n2584 185
R10979 VDD.n2584 VDD.n2583 185
R10980 VDD.n870 VDD.n869 185
R10981 VDD.n871 VDD.n870 185
R10982 VDD.n2576 VDD.n2575 185
R10983 VDD.n2577 VDD.n2576 185
R10984 VDD.n2574 VDD.n880 185
R10985 VDD.n880 VDD.n877 185
R10986 VDD.n2573 VDD.n2572 185
R10987 VDD.n2572 VDD.n2571 185
R10988 VDD.n882 VDD.n881 185
R10989 VDD.n891 VDD.n882 185
R10990 VDD.n2564 VDD.n2563 185
R10991 VDD.n2565 VDD.n2564 185
R10992 VDD.n2562 VDD.n892 185
R10993 VDD.n892 VDD.n888 185
R10994 VDD.n2561 VDD.n2560 185
R10995 VDD.n2560 VDD.n2559 185
R10996 VDD.n894 VDD.n893 185
R10997 VDD.n895 VDD.n894 185
R10998 VDD.n2552 VDD.n2551 185
R10999 VDD.n2553 VDD.n2552 185
R11000 VDD.n2550 VDD.n904 185
R11001 VDD.n904 VDD.n901 185
R11002 VDD.n2549 VDD.n2548 185
R11003 VDD.n2548 VDD.n2547 185
R11004 VDD.n906 VDD.n905 185
R11005 VDD.n907 VDD.n906 185
R11006 VDD.n2540 VDD.n2539 185
R11007 VDD.n2541 VDD.n2540 185
R11008 VDD.n2538 VDD.n916 185
R11009 VDD.n916 VDD.n913 185
R11010 VDD.n2537 VDD.n2536 185
R11011 VDD.n2536 VDD.n2535 185
R11012 VDD.n918 VDD.n917 185
R11013 VDD.n919 VDD.n918 185
R11014 VDD.n2528 VDD.n2527 185
R11015 VDD.n2529 VDD.n2528 185
R11016 VDD.n2526 VDD.n928 185
R11017 VDD.n928 VDD.n925 185
R11018 VDD.n2525 VDD.n2524 185
R11019 VDD.n2524 VDD.n2523 185
R11020 VDD.n930 VDD.n929 185
R11021 VDD.n939 VDD.n930 185
R11022 VDD.n2516 VDD.n2515 185
R11023 VDD.n2517 VDD.n2516 185
R11024 VDD.n2514 VDD.n940 185
R11025 VDD.n940 VDD.n936 185
R11026 VDD.n2513 VDD.n2512 185
R11027 VDD.n2512 VDD.n2511 185
R11028 VDD.n942 VDD.n941 185
R11029 VDD.n943 VDD.n942 185
R11030 VDD.n2504 VDD.n2503 185
R11031 VDD.n2505 VDD.n2504 185
R11032 VDD.n2502 VDD.n952 185
R11033 VDD.n952 VDD.n949 185
R11034 VDD.n2501 VDD.n2500 185
R11035 VDD.n2500 VDD.n2499 185
R11036 VDD.n954 VDD.n953 185
R11037 VDD.n955 VDD.n954 185
R11038 VDD.n2492 VDD.n2491 185
R11039 VDD.n2493 VDD.n2492 185
R11040 VDD.n2490 VDD.n964 185
R11041 VDD.n964 VDD.n961 185
R11042 VDD.n2489 VDD.n2488 185
R11043 VDD.n2488 VDD.n2487 185
R11044 VDD.n966 VDD.n965 185
R11045 VDD.n967 VDD.n966 185
R11046 VDD.n2480 VDD.n2479 185
R11047 VDD.n2481 VDD.n2480 185
R11048 VDD.n2478 VDD.n976 185
R11049 VDD.n976 VDD.n973 185
R11050 VDD.n2477 VDD.n2476 185
R11051 VDD.n2476 VDD.n2475 185
R11052 VDD.n978 VDD.n977 185
R11053 VDD.n979 VDD.n978 185
R11054 VDD.n2468 VDD.n2467 185
R11055 VDD.n2469 VDD.n2468 185
R11056 VDD.n2466 VDD.n988 185
R11057 VDD.n988 VDD.n985 185
R11058 VDD.n2465 VDD.n2464 185
R11059 VDD.n2464 VDD.n2463 185
R11060 VDD.n990 VDD.n989 185
R11061 VDD.n991 VDD.n990 185
R11062 VDD.n2456 VDD.n2455 185
R11063 VDD.n2457 VDD.n2456 185
R11064 VDD.n2454 VDD.n999 185
R11065 VDD.n1005 VDD.n999 185
R11066 VDD.n2453 VDD.n2452 185
R11067 VDD.n2452 VDD.n2451 185
R11068 VDD.n1001 VDD.n1000 185
R11069 VDD.n1002 VDD.n1001 185
R11070 VDD.n2444 VDD.n2443 185
R11071 VDD.n2445 VDD.n2444 185
R11072 VDD.n2442 VDD.n1012 185
R11073 VDD.n1012 VDD.n1009 185
R11074 VDD.n2441 VDD.n2440 185
R11075 VDD.n2440 VDD.n2439 185
R11076 VDD.n1014 VDD.n1013 185
R11077 VDD.n1015 VDD.n1014 185
R11078 VDD.n2432 VDD.n2431 185
R11079 VDD.n2433 VDD.n2432 185
R11080 VDD.n2430 VDD.n1024 185
R11081 VDD.n1024 VDD.n1021 185
R11082 VDD.n2429 VDD.n2428 185
R11083 VDD.n2428 VDD.n2427 185
R11084 VDD.n1026 VDD.n1025 185
R11085 VDD.n1035 VDD.n1026 185
R11086 VDD.n2420 VDD.n2419 185
R11087 VDD.n2421 VDD.n2420 185
R11088 VDD.n2418 VDD.n1036 185
R11089 VDD.n1036 VDD.n1032 185
R11090 VDD.n2417 VDD.n2416 185
R11091 VDD.n2416 VDD.n2415 185
R11092 VDD.n1038 VDD.n1037 185
R11093 VDD.n1039 VDD.n1038 185
R11094 VDD.n2408 VDD.n2407 185
R11095 VDD.n2409 VDD.n2408 185
R11096 VDD.n2406 VDD.n1048 185
R11097 VDD.n1048 VDD.n1045 185
R11098 VDD.n2405 VDD.n2404 185
R11099 VDD.n2404 VDD.n2403 185
R11100 VDD.n1050 VDD.n1049 185
R11101 VDD.n1051 VDD.n1050 185
R11102 VDD.n2396 VDD.n2395 185
R11103 VDD.n2397 VDD.n2396 185
R11104 VDD.n2394 VDD.n1059 185
R11105 VDD.n2393 VDD.n2392 185
R11106 VDD.n1061 VDD.n1060 185
R11107 VDD.n2390 VDD.n1061 185
R11108 VDD.n2039 VDD.n2038 185
R11109 VDD.n2041 VDD.n2040 185
R11110 VDD.n2043 VDD.n2042 185
R11111 VDD.n2045 VDD.n2044 185
R11112 VDD.n2047 VDD.n2046 185
R11113 VDD.n2049 VDD.n2048 185
R11114 VDD.n2051 VDD.n2050 185
R11115 VDD.n2194 VDD.n2052 185
R11116 VDD.n2196 VDD.n2195 185
R11117 VDD.n2193 VDD.n2192 185
R11118 VDD.n2191 VDD.n2190 185
R11119 VDD.n2189 VDD.n2188 185
R11120 VDD.n2187 VDD.n2186 185
R11121 VDD.n2185 VDD.n2184 185
R11122 VDD.n2183 VDD.n2182 185
R11123 VDD.n2181 VDD.n2180 185
R11124 VDD.n2179 VDD.n2178 185
R11125 VDD.n2176 VDD.n2175 185
R11126 VDD.n2174 VDD.n1071 185
R11127 VDD.n2390 VDD.n1071 185
R11128 VDD.n2650 VDD.n2649 185
R11129 VDD.n2652 VDD.n2651 185
R11130 VDD.n2654 VDD.n2653 185
R11131 VDD.n2656 VDD.n2655 185
R11132 VDD.n2658 VDD.n2657 185
R11133 VDD.n2660 VDD.n2659 185
R11134 VDD.n2662 VDD.n2661 185
R11135 VDD.n2664 VDD.n2663 185
R11136 VDD.n2666 VDD.n2665 185
R11137 VDD.n2668 VDD.n2667 185
R11138 VDD.n2670 VDD.n2669 185
R11139 VDD.n2672 VDD.n2671 185
R11140 VDD.n2674 VDD.n2673 185
R11141 VDD.n2676 VDD.n2675 185
R11142 VDD.n2678 VDD.n2677 185
R11143 VDD.n2680 VDD.n2679 185
R11144 VDD.n2682 VDD.n2681 185
R11145 VDD.n2684 VDD.n2683 185
R11146 VDD.n2686 VDD.n2685 185
R11147 VDD.n2688 VDD.n2687 185
R11148 VDD.n2690 VDD.n2689 185
R11149 VDD.n2692 VDD.n2691 185
R11150 VDD.n2648 VDD.n2647 185
R11151 VDD.n2648 VDD.n775 185
R11152 VDD.n2646 VDD.n806 185
R11153 VDD.n2696 VDD.n806 185
R11154 VDD.n2645 VDD.n2644 185
R11155 VDD.n2644 VDD.n805 185
R11156 VDD.n2643 VDD.n814 185
R11157 VDD.n2643 VDD.n2642 185
R11158 VDD.n2055 VDD.n815 185
R11159 VDD.n816 VDD.n815 185
R11160 VDD.n2056 VDD.n823 185
R11161 VDD.n2636 VDD.n823 185
R11162 VDD.n2058 VDD.n2057 185
R11163 VDD.n2057 VDD.n822 185
R11164 VDD.n2059 VDD.n830 185
R11165 VDD.n2625 VDD.n830 185
R11166 VDD.n2061 VDD.n2060 185
R11167 VDD.n2060 VDD.n829 185
R11168 VDD.n2062 VDD.n836 185
R11169 VDD.n2619 VDD.n836 185
R11170 VDD.n2064 VDD.n2063 185
R11171 VDD.n2063 VDD.n835 185
R11172 VDD.n2065 VDD.n842 185
R11173 VDD.n2613 VDD.n842 185
R11174 VDD.n2067 VDD.n2066 185
R11175 VDD.n2066 VDD.n841 185
R11176 VDD.n2068 VDD.n848 185
R11177 VDD.n2607 VDD.n848 185
R11178 VDD.n2070 VDD.n2069 185
R11179 VDD.n2069 VDD.n847 185
R11180 VDD.n2071 VDD.n854 185
R11181 VDD.n2601 VDD.n854 185
R11182 VDD.n2073 VDD.n2072 185
R11183 VDD.n2072 VDD.n853 185
R11184 VDD.n2074 VDD.n860 185
R11185 VDD.n2595 VDD.n860 185
R11186 VDD.n2076 VDD.n2075 185
R11187 VDD.n2075 VDD.n859 185
R11188 VDD.n2077 VDD.n866 185
R11189 VDD.n2589 VDD.n866 185
R11190 VDD.n2079 VDD.n2078 185
R11191 VDD.n2078 VDD.n865 185
R11192 VDD.n2080 VDD.n872 185
R11193 VDD.n2583 VDD.n872 185
R11194 VDD.n2082 VDD.n2081 185
R11195 VDD.n2081 VDD.n871 185
R11196 VDD.n2083 VDD.n878 185
R11197 VDD.n2577 VDD.n878 185
R11198 VDD.n2085 VDD.n2084 185
R11199 VDD.n2084 VDD.n877 185
R11200 VDD.n2086 VDD.n883 185
R11201 VDD.n2571 VDD.n883 185
R11202 VDD.n2088 VDD.n2087 185
R11203 VDD.n2087 VDD.n891 185
R11204 VDD.n2089 VDD.n889 185
R11205 VDD.n2565 VDD.n889 185
R11206 VDD.n2091 VDD.n2090 185
R11207 VDD.n2090 VDD.n888 185
R11208 VDD.n2092 VDD.n896 185
R11209 VDD.n2559 VDD.n896 185
R11210 VDD.n2094 VDD.n2093 185
R11211 VDD.n2093 VDD.n895 185
R11212 VDD.n2095 VDD.n902 185
R11213 VDD.n2553 VDD.n902 185
R11214 VDD.n2097 VDD.n2096 185
R11215 VDD.n2096 VDD.n901 185
R11216 VDD.n2098 VDD.n908 185
R11217 VDD.n2547 VDD.n908 185
R11218 VDD.n2100 VDD.n2099 185
R11219 VDD.n2099 VDD.n907 185
R11220 VDD.n2101 VDD.n914 185
R11221 VDD.n2541 VDD.n914 185
R11222 VDD.n2103 VDD.n2102 185
R11223 VDD.n2102 VDD.n913 185
R11224 VDD.n2104 VDD.n920 185
R11225 VDD.n2535 VDD.n920 185
R11226 VDD.n2106 VDD.n2105 185
R11227 VDD.n2105 VDD.n919 185
R11228 VDD.n2107 VDD.n926 185
R11229 VDD.n2529 VDD.n926 185
R11230 VDD.n2109 VDD.n2108 185
R11231 VDD.n2108 VDD.n925 185
R11232 VDD.n2110 VDD.n931 185
R11233 VDD.n2523 VDD.n931 185
R11234 VDD.n2112 VDD.n2111 185
R11235 VDD.n2111 VDD.n939 185
R11236 VDD.n2113 VDD.n937 185
R11237 VDD.n2517 VDD.n937 185
R11238 VDD.n2115 VDD.n2114 185
R11239 VDD.n2114 VDD.n936 185
R11240 VDD.n2116 VDD.n944 185
R11241 VDD.n2511 VDD.n944 185
R11242 VDD.n2118 VDD.n2117 185
R11243 VDD.n2117 VDD.n943 185
R11244 VDD.n2119 VDD.n950 185
R11245 VDD.n2505 VDD.n950 185
R11246 VDD.n2121 VDD.n2120 185
R11247 VDD.n2120 VDD.n949 185
R11248 VDD.n2122 VDD.n956 185
R11249 VDD.n2499 VDD.n956 185
R11250 VDD.n2124 VDD.n2123 185
R11251 VDD.n2123 VDD.n955 185
R11252 VDD.n2125 VDD.n962 185
R11253 VDD.n2493 VDD.n962 185
R11254 VDD.n2127 VDD.n2126 185
R11255 VDD.n2126 VDD.n961 185
R11256 VDD.n2128 VDD.n968 185
R11257 VDD.n2487 VDD.n968 185
R11258 VDD.n2130 VDD.n2129 185
R11259 VDD.n2129 VDD.n967 185
R11260 VDD.n2131 VDD.n974 185
R11261 VDD.n2481 VDD.n974 185
R11262 VDD.n2133 VDD.n2132 185
R11263 VDD.n2132 VDD.n973 185
R11264 VDD.n2134 VDD.n980 185
R11265 VDD.n2475 VDD.n980 185
R11266 VDD.n2136 VDD.n2135 185
R11267 VDD.n2135 VDD.n979 185
R11268 VDD.n2137 VDD.n986 185
R11269 VDD.n2469 VDD.n986 185
R11270 VDD.n2139 VDD.n2138 185
R11271 VDD.n2138 VDD.n985 185
R11272 VDD.n2140 VDD.n992 185
R11273 VDD.n2463 VDD.n992 185
R11274 VDD.n2142 VDD.n2141 185
R11275 VDD.n2141 VDD.n991 185
R11276 VDD.n2143 VDD.n997 185
R11277 VDD.n2457 VDD.n997 185
R11278 VDD.n2145 VDD.n2144 185
R11279 VDD.n2144 VDD.n1005 185
R11280 VDD.n2146 VDD.n1003 185
R11281 VDD.n2451 VDD.n1003 185
R11282 VDD.n2148 VDD.n2147 185
R11283 VDD.n2147 VDD.n1002 185
R11284 VDD.n2149 VDD.n1010 185
R11285 VDD.n2445 VDD.n1010 185
R11286 VDD.n2151 VDD.n2150 185
R11287 VDD.n2150 VDD.n1009 185
R11288 VDD.n2152 VDD.n1016 185
R11289 VDD.n2439 VDD.n1016 185
R11290 VDD.n2154 VDD.n2153 185
R11291 VDD.n2153 VDD.n1015 185
R11292 VDD.n2155 VDD.n1022 185
R11293 VDD.n2433 VDD.n1022 185
R11294 VDD.n2157 VDD.n2156 185
R11295 VDD.n2156 VDD.n1021 185
R11296 VDD.n2158 VDD.n1027 185
R11297 VDD.n2427 VDD.n1027 185
R11298 VDD.n2160 VDD.n2159 185
R11299 VDD.n2159 VDD.n1035 185
R11300 VDD.n2161 VDD.n1033 185
R11301 VDD.n2421 VDD.n1033 185
R11302 VDD.n2163 VDD.n2162 185
R11303 VDD.n2162 VDD.n1032 185
R11304 VDD.n2164 VDD.n1040 185
R11305 VDD.n2415 VDD.n1040 185
R11306 VDD.n2166 VDD.n2165 185
R11307 VDD.n2165 VDD.n1039 185
R11308 VDD.n2167 VDD.n1046 185
R11309 VDD.n2409 VDD.n1046 185
R11310 VDD.n2169 VDD.n2168 185
R11311 VDD.n2168 VDD.n1045 185
R11312 VDD.n2170 VDD.n1052 185
R11313 VDD.n2403 VDD.n1052 185
R11314 VDD.n2172 VDD.n2171 185
R11315 VDD.n2171 VDD.n1051 185
R11316 VDD.n2173 VDD.n1057 185
R11317 VDD.n2397 VDD.n1057 185
R11318 VDD.n3881 VDD.n243 185
R11319 VDD.n243 VDD.n242 185
R11320 VDD.n3883 VDD.n3882 185
R11321 VDD.n3884 VDD.n3883 185
R11322 VDD.n238 VDD.n237 185
R11323 VDD.n3885 VDD.n238 185
R11324 VDD.n3888 VDD.n3887 185
R11325 VDD.n3887 VDD.n3886 185
R11326 VDD.n3889 VDD.n232 185
R11327 VDD.n232 VDD.n231 185
R11328 VDD.n3891 VDD.n3890 185
R11329 VDD.n3892 VDD.n3891 185
R11330 VDD.n227 VDD.n226 185
R11331 VDD.n3893 VDD.n227 185
R11332 VDD.n3896 VDD.n3895 185
R11333 VDD.n3895 VDD.n3894 185
R11334 VDD.n3897 VDD.n221 185
R11335 VDD.n221 VDD.n220 185
R11336 VDD.n3899 VDD.n3898 185
R11337 VDD.n3900 VDD.n3899 185
R11338 VDD.n216 VDD.n215 185
R11339 VDD.n3901 VDD.n216 185
R11340 VDD.n3904 VDD.n3903 185
R11341 VDD.n3903 VDD.n3902 185
R11342 VDD.n3905 VDD.n210 185
R11343 VDD.n210 VDD.n209 185
R11344 VDD.n3907 VDD.n3906 185
R11345 VDD.n3908 VDD.n3907 185
R11346 VDD.n205 VDD.n204 185
R11347 VDD.n3909 VDD.n205 185
R11348 VDD.n3912 VDD.n3911 185
R11349 VDD.n3911 VDD.n3910 185
R11350 VDD.n3913 VDD.n199 185
R11351 VDD.n199 VDD.n198 185
R11352 VDD.n3915 VDD.n3914 185
R11353 VDD.n3916 VDD.n3915 185
R11354 VDD.n194 VDD.n193 185
R11355 VDD.n3917 VDD.n194 185
R11356 VDD.n3920 VDD.n3919 185
R11357 VDD.n3919 VDD.n3918 185
R11358 VDD.n3921 VDD.n188 185
R11359 VDD.n188 VDD.n187 185
R11360 VDD.n3923 VDD.n3922 185
R11361 VDD.n3924 VDD.n3923 185
R11362 VDD.n183 VDD.n182 185
R11363 VDD.n3925 VDD.n183 185
R11364 VDD.n3928 VDD.n3927 185
R11365 VDD.n3927 VDD.n3926 185
R11366 VDD.n3929 VDD.n177 185
R11367 VDD.n177 VDD.n176 185
R11368 VDD.n3931 VDD.n3930 185
R11369 VDD.n3932 VDD.n3931 185
R11370 VDD.n172 VDD.n171 185
R11371 VDD.n3933 VDD.n172 185
R11372 VDD.n3936 VDD.n3935 185
R11373 VDD.n3935 VDD.n3934 185
R11374 VDD.n3937 VDD.n166 185
R11375 VDD.n166 VDD.n165 185
R11376 VDD.n3939 VDD.n3938 185
R11377 VDD.n3940 VDD.n3939 185
R11378 VDD.n161 VDD.n160 185
R11379 VDD.n3941 VDD.n161 185
R11380 VDD.n3944 VDD.n3943 185
R11381 VDD.n3943 VDD.n3942 185
R11382 VDD.n3945 VDD.n156 185
R11383 VDD.n156 VDD.n155 185
R11384 VDD.n3947 VDD.n3946 185
R11385 VDD.n3948 VDD.n3947 185
R11386 VDD.n150 VDD.n148 185
R11387 VDD.n3949 VDD.n150 185
R11388 VDD.n3952 VDD.n3951 185
R11389 VDD.n3951 VDD.n3950 185
R11390 VDD.n149 VDD.n147 185
R11391 VDD.n151 VDD.n149 185
R11392 VDD.n3720 VDD.n3719 185
R11393 VDD.n3721 VDD.n3720 185
R11394 VDD.n351 VDD.n350 185
R11395 VDD.n350 VDD.n349 185
R11396 VDD.n3715 VDD.n3714 185
R11397 VDD.n3714 VDD.n3713 185
R11398 VDD.n354 VDD.n353 185
R11399 VDD.n355 VDD.n354 185
R11400 VDD.n3701 VDD.n3700 185
R11401 VDD.n3702 VDD.n3701 185
R11402 VDD.n362 VDD.n361 185
R11403 VDD.n3693 VDD.n361 185
R11404 VDD.n3696 VDD.n3695 185
R11405 VDD.n3695 VDD.n3694 185
R11406 VDD.n365 VDD.n364 185
R11407 VDD.n366 VDD.n365 185
R11408 VDD.n3684 VDD.n3683 185
R11409 VDD.n3685 VDD.n3684 185
R11410 VDD.n374 VDD.n373 185
R11411 VDD.n373 VDD.n372 185
R11412 VDD.n3679 VDD.n3678 185
R11413 VDD.n3678 VDD.n3677 185
R11414 VDD.n377 VDD.n376 185
R11415 VDD.n378 VDD.n377 185
R11416 VDD.n3668 VDD.n3667 185
R11417 VDD.n3669 VDD.n3668 185
R11418 VDD.n386 VDD.n385 185
R11419 VDD.n385 VDD.n384 185
R11420 VDD.n3663 VDD.n3662 185
R11421 VDD.n3662 VDD.n3661 185
R11422 VDD.n389 VDD.n388 185
R11423 VDD.n390 VDD.n389 185
R11424 VDD.n3652 VDD.n3651 185
R11425 VDD.n3653 VDD.n3652 185
R11426 VDD.n398 VDD.n397 185
R11427 VDD.n397 VDD.n396 185
R11428 VDD.n3647 VDD.n3646 185
R11429 VDD.n3646 VDD.n3645 185
R11430 VDD.n401 VDD.n400 185
R11431 VDD.n402 VDD.n401 185
R11432 VDD.n3636 VDD.n3635 185
R11433 VDD.n3637 VDD.n3636 185
R11434 VDD.n410 VDD.n409 185
R11435 VDD.n409 VDD.n408 185
R11436 VDD.n3631 VDD.n3630 185
R11437 VDD.n3630 VDD.n3629 185
R11438 VDD.n413 VDD.n412 185
R11439 VDD.n414 VDD.n413 185
R11440 VDD.n3620 VDD.n3619 185
R11441 VDD.n3621 VDD.n3620 185
R11442 VDD.n422 VDD.n421 185
R11443 VDD.n421 VDD.n420 185
R11444 VDD.n3615 VDD.n3614 185
R11445 VDD.n3614 VDD.n3613 185
R11446 VDD.n425 VDD.n424 185
R11447 VDD.n426 VDD.n425 185
R11448 VDD.n3604 VDD.n3603 185
R11449 VDD.n3605 VDD.n3604 185
R11450 VDD.n433 VDD.n432 185
R11451 VDD.n3596 VDD.n432 185
R11452 VDD.n3599 VDD.n3598 185
R11453 VDD.n3598 VDD.n3597 185
R11454 VDD.n436 VDD.n435 185
R11455 VDD.n437 VDD.n436 185
R11456 VDD.n3587 VDD.n3586 185
R11457 VDD.n3588 VDD.n3587 185
R11458 VDD.n445 VDD.n444 185
R11459 VDD.n444 VDD.n443 185
R11460 VDD.n3582 VDD.n3581 185
R11461 VDD.n3581 VDD.n3580 185
R11462 VDD.n3460 VDD.n447 185
R11463 VDD.n3465 VDD.n3463 185
R11464 VDD.n3466 VDD.n3459 185
R11465 VDD.n3466 VDD.n448 185
R11466 VDD.n3469 VDD.n3468 185
R11467 VDD.n3471 VDD.n3458 185
R11468 VDD.n3473 VDD.n3472 185
R11469 VDD.n3476 VDD.n3475 185
R11470 VDD.n3477 VDD.n3454 185
R11471 VDD.n492 VDD.n491 185
R11472 VDD.n3482 VDD.n3481 185
R11473 VDD.n3484 VDD.n490 185
R11474 VDD.n3487 VDD.n3486 185
R11475 VDD.n488 VDD.n487 185
R11476 VDD.n3492 VDD.n3491 185
R11477 VDD.n3494 VDD.n486 185
R11478 VDD.n3497 VDD.n3496 185
R11479 VDD.n484 VDD.n481 185
R11480 VDD.n3502 VDD.n3501 185
R11481 VDD.n3504 VDD.n480 185
R11482 VDD.n3507 VDD.n3506 185
R11483 VDD.n478 VDD.n477 185
R11484 VDD.n3512 VDD.n3511 185
R11485 VDD.n3514 VDD.n476 185
R11486 VDD.n3517 VDD.n3516 185
R11487 VDD.n474 VDD.n473 185
R11488 VDD.n3525 VDD.n3524 185
R11489 VDD.n3527 VDD.n472 185
R11490 VDD.n3530 VDD.n3529 185
R11491 VDD.n470 VDD.n469 185
R11492 VDD.n3535 VDD.n3534 185
R11493 VDD.n3537 VDD.n468 185
R11494 VDD.n3540 VDD.n3539 185
R11495 VDD.n466 VDD.n465 185
R11496 VDD.n3545 VDD.n3544 185
R11497 VDD.n3547 VDD.n464 185
R11498 VDD.n3552 VDD.n3549 185
R11499 VDD.n462 VDD.n461 185
R11500 VDD.n3557 VDD.n3556 185
R11501 VDD.n3559 VDD.n460 185
R11502 VDD.n3562 VDD.n3561 185
R11503 VDD.n456 VDD.n455 185
R11504 VDD.n3567 VDD.n3566 185
R11505 VDD.n3569 VDD.n454 185
R11506 VDD.n3570 VDD.n453 185
R11507 VDD.n3573 VDD.n3572 185
R11508 VDD.n3575 VDD.n449 185
R11509 VDD.n449 VDD.n448 185
R11510 VDD.n3789 VDD.n3788 185
R11511 VDD.n3793 VDD.n322 185
R11512 VDD.n3795 VDD.n3794 185
R11513 VDD.n3797 VDD.n320 185
R11514 VDD.n3799 VDD.n3798 185
R11515 VDD.n3800 VDD.n316 185
R11516 VDD.n3802 VDD.n3801 185
R11517 VDD.n3804 VDD.n313 185
R11518 VDD.n3806 VDD.n3805 185
R11519 VDD.n314 VDD.n307 185
R11520 VDD.n3810 VDD.n311 185
R11521 VDD.n3811 VDD.n303 185
R11522 VDD.n3813 VDD.n3812 185
R11523 VDD.n3815 VDD.n301 185
R11524 VDD.n3817 VDD.n3816 185
R11525 VDD.n3818 VDD.n296 185
R11526 VDD.n3820 VDD.n3819 185
R11527 VDD.n3822 VDD.n294 185
R11528 VDD.n3824 VDD.n3823 185
R11529 VDD.n3825 VDD.n289 185
R11530 VDD.n3830 VDD.n3829 185
R11531 VDD.n3832 VDD.n287 185
R11532 VDD.n3834 VDD.n3833 185
R11533 VDD.n3835 VDD.n282 185
R11534 VDD.n3837 VDD.n3836 185
R11535 VDD.n3839 VDD.n281 185
R11536 VDD.n3840 VDD.n278 185
R11537 VDD.n3843 VDD.n3842 185
R11538 VDD.n280 VDD.n274 185
R11539 VDD.n3847 VDD.n271 185
R11540 VDD.n3849 VDD.n3848 185
R11541 VDD.n3851 VDD.n269 185
R11542 VDD.n3853 VDD.n3852 185
R11543 VDD.n3854 VDD.n265 185
R11544 VDD.n3856 VDD.n3855 185
R11545 VDD.n3858 VDD.n263 185
R11546 VDD.n3860 VDD.n3859 185
R11547 VDD.n258 VDD.n257 185
R11548 VDD.n3865 VDD.n3864 185
R11549 VDD.n3867 VDD.n255 185
R11550 VDD.n3869 VDD.n3868 185
R11551 VDD.n3870 VDD.n250 185
R11552 VDD.n3872 VDD.n3871 185
R11553 VDD.n3874 VDD.n249 185
R11554 VDD.n3875 VDD.n247 185
R11555 VDD.n3878 VDD.n3877 185
R11556 VDD.n3787 VDD.n3786 185
R11557 VDD.n3787 VDD.n242 185
R11558 VDD.n328 VDD.n241 185
R11559 VDD.n3884 VDD.n241 185
R11560 VDD.n3782 VDD.n240 185
R11561 VDD.n3885 VDD.n240 185
R11562 VDD.n3781 VDD.n239 185
R11563 VDD.n3886 VDD.n239 185
R11564 VDD.n3780 VDD.n3779 185
R11565 VDD.n3779 VDD.n231 185
R11566 VDD.n330 VDD.n230 185
R11567 VDD.n3892 VDD.n230 185
R11568 VDD.n3775 VDD.n229 185
R11569 VDD.n3893 VDD.n229 185
R11570 VDD.n3774 VDD.n228 185
R11571 VDD.n3894 VDD.n228 185
R11572 VDD.n3773 VDD.n3772 185
R11573 VDD.n3772 VDD.n220 185
R11574 VDD.n332 VDD.n219 185
R11575 VDD.n3900 VDD.n219 185
R11576 VDD.n3768 VDD.n218 185
R11577 VDD.n3901 VDD.n218 185
R11578 VDD.n3767 VDD.n217 185
R11579 VDD.n3902 VDD.n217 185
R11580 VDD.n3766 VDD.n3765 185
R11581 VDD.n3765 VDD.n209 185
R11582 VDD.n334 VDD.n208 185
R11583 VDD.n3908 VDD.n208 185
R11584 VDD.n3761 VDD.n207 185
R11585 VDD.n3909 VDD.n207 185
R11586 VDD.n3760 VDD.n206 185
R11587 VDD.n3910 VDD.n206 185
R11588 VDD.n3759 VDD.n3758 185
R11589 VDD.n3758 VDD.n198 185
R11590 VDD.n336 VDD.n197 185
R11591 VDD.n3916 VDD.n197 185
R11592 VDD.n3754 VDD.n196 185
R11593 VDD.n3917 VDD.n196 185
R11594 VDD.n3753 VDD.n195 185
R11595 VDD.n3918 VDD.n195 185
R11596 VDD.n3752 VDD.n3751 185
R11597 VDD.n3751 VDD.n187 185
R11598 VDD.n338 VDD.n186 185
R11599 VDD.n3924 VDD.n186 185
R11600 VDD.n3747 VDD.n185 185
R11601 VDD.n3925 VDD.n185 185
R11602 VDD.n3746 VDD.n184 185
R11603 VDD.n3926 VDD.n184 185
R11604 VDD.n3745 VDD.n3744 185
R11605 VDD.n3744 VDD.n176 185
R11606 VDD.n340 VDD.n175 185
R11607 VDD.n3932 VDD.n175 185
R11608 VDD.n3740 VDD.n174 185
R11609 VDD.n3933 VDD.n174 185
R11610 VDD.n3739 VDD.n173 185
R11611 VDD.n3934 VDD.n173 185
R11612 VDD.n3738 VDD.n3737 185
R11613 VDD.n3737 VDD.n165 185
R11614 VDD.n342 VDD.n164 185
R11615 VDD.n3940 VDD.n164 185
R11616 VDD.n3733 VDD.n163 185
R11617 VDD.n3941 VDD.n163 185
R11618 VDD.n3732 VDD.n162 185
R11619 VDD.n3942 VDD.n162 185
R11620 VDD.n3731 VDD.n3730 185
R11621 VDD.n3730 VDD.n155 185
R11622 VDD.n344 VDD.n154 185
R11623 VDD.n3948 VDD.n154 185
R11624 VDD.n3726 VDD.n153 185
R11625 VDD.n3949 VDD.n153 185
R11626 VDD.n3725 VDD.n152 185
R11627 VDD.n3950 VDD.n152 185
R11628 VDD.n3724 VDD.n3723 185
R11629 VDD.n3723 VDD.n151 185
R11630 VDD.n3722 VDD.n346 185
R11631 VDD.n3722 VDD.n3721 185
R11632 VDD.n3710 VDD.n348 185
R11633 VDD.n349 VDD.n348 185
R11634 VDD.n3712 VDD.n3711 185
R11635 VDD.n3713 VDD.n3712 185
R11636 VDD.n357 VDD.n356 185
R11637 VDD.n356 VDD.n355 185
R11638 VDD.n3704 VDD.n3703 185
R11639 VDD.n3703 VDD.n3702 185
R11640 VDD.n360 VDD.n359 185
R11641 VDD.n3693 VDD.n360 185
R11642 VDD.n3692 VDD.n3691 185
R11643 VDD.n3694 VDD.n3692 185
R11644 VDD.n368 VDD.n367 185
R11645 VDD.n367 VDD.n366 185
R11646 VDD.n3687 VDD.n3686 185
R11647 VDD.n3686 VDD.n3685 185
R11648 VDD.n371 VDD.n370 185
R11649 VDD.n372 VDD.n371 185
R11650 VDD.n3676 VDD.n3675 185
R11651 VDD.n3677 VDD.n3676 185
R11652 VDD.n380 VDD.n379 185
R11653 VDD.n379 VDD.n378 185
R11654 VDD.n3671 VDD.n3670 185
R11655 VDD.n3670 VDD.n3669 185
R11656 VDD.n383 VDD.n382 185
R11657 VDD.n384 VDD.n383 185
R11658 VDD.n3660 VDD.n3659 185
R11659 VDD.n3661 VDD.n3660 185
R11660 VDD.n392 VDD.n391 185
R11661 VDD.n391 VDD.n390 185
R11662 VDD.n3655 VDD.n3654 185
R11663 VDD.n3654 VDD.n3653 185
R11664 VDD.n395 VDD.n394 185
R11665 VDD.n396 VDD.n395 185
R11666 VDD.n3644 VDD.n3643 185
R11667 VDD.n3645 VDD.n3644 185
R11668 VDD.n404 VDD.n403 185
R11669 VDD.n403 VDD.n402 185
R11670 VDD.n3639 VDD.n3638 185
R11671 VDD.n3638 VDD.n3637 185
R11672 VDD.n407 VDD.n406 185
R11673 VDD.n408 VDD.n407 185
R11674 VDD.n3628 VDD.n3627 185
R11675 VDD.n3629 VDD.n3628 185
R11676 VDD.n416 VDD.n415 185
R11677 VDD.n415 VDD.n414 185
R11678 VDD.n3623 VDD.n3622 185
R11679 VDD.n3622 VDD.n3621 185
R11680 VDD.n419 VDD.n418 185
R11681 VDD.n420 VDD.n419 185
R11682 VDD.n3612 VDD.n3611 185
R11683 VDD.n3613 VDD.n3612 185
R11684 VDD.n428 VDD.n427 185
R11685 VDD.n427 VDD.n426 185
R11686 VDD.n3607 VDD.n3606 185
R11687 VDD.n3606 VDD.n3605 185
R11688 VDD.n431 VDD.n430 185
R11689 VDD.n3596 VDD.n431 185
R11690 VDD.n3595 VDD.n3594 185
R11691 VDD.n3597 VDD.n3595 185
R11692 VDD.n439 VDD.n438 185
R11693 VDD.n438 VDD.n437 185
R11694 VDD.n3590 VDD.n3589 185
R11695 VDD.n3589 VDD.n3588 185
R11696 VDD.n442 VDD.n441 185
R11697 VDD.n443 VDD.n442 185
R11698 VDD.n3579 VDD.n3578 185
R11699 VDD.n3580 VDD.n3579 185
R11700 VDD.n774 VDD.n773 185
R11701 VDD.n2792 VDD.n2791 185
R11702 VDD.n2793 VDD.n2789 185
R11703 VDD.n2789 VDD.n2744 185
R11704 VDD.n2795 VDD.n2794 185
R11705 VDD.n2797 VDD.n2788 185
R11706 VDD.n2800 VDD.n2799 185
R11707 VDD.n2801 VDD.n2787 185
R11708 VDD.n2803 VDD.n2802 185
R11709 VDD.n2805 VDD.n2786 185
R11710 VDD.n2808 VDD.n2807 185
R11711 VDD.n2809 VDD.n2785 185
R11712 VDD.n2811 VDD.n2810 185
R11713 VDD.n2813 VDD.n2784 185
R11714 VDD.n2816 VDD.n2815 185
R11715 VDD.n2817 VDD.n2783 185
R11716 VDD.n2819 VDD.n2818 185
R11717 VDD.n2821 VDD.n2782 185
R11718 VDD.n2824 VDD.n2823 185
R11719 VDD.n2825 VDD.n2781 185
R11720 VDD.n2830 VDD.n2829 185
R11721 VDD.n2832 VDD.n2780 185
R11722 VDD.n2834 VDD.n2833 185
R11723 VDD.n2833 VDD.n2744 185
R11724 VDD.n3432 VDD.n3431 185
R11725 VDD.n3434 VDD.n505 185
R11726 VDD.n3436 VDD.n3435 185
R11727 VDD.n3437 VDD.n500 185
R11728 VDD.n3439 VDD.n3438 185
R11729 VDD.n3441 VDD.n498 185
R11730 VDD.n3443 VDD.n3442 185
R11731 VDD.n3444 VDD.n497 185
R11732 VDD.n3446 VDD.n3445 185
R11733 VDD.n3448 VDD.n494 185
R11734 VDD.n3450 VDD.n3449 185
R11735 VDD.n3405 VDD.n493 185
R11736 VDD.n3407 VDD.n3406 185
R11737 VDD.n3408 VDD.n3403 185
R11738 VDD.n3410 VDD.n3409 185
R11739 VDD.n3412 VDD.n3401 185
R11740 VDD.n3414 VDD.n3413 185
R11741 VDD.n3415 VDD.n3400 185
R11742 VDD.n3417 VDD.n3416 185
R11743 VDD.n3419 VDD.n3399 185
R11744 VDD.n3420 VDD.n3398 185
R11745 VDD.n3423 VDD.n3422 185
R11746 VDD.n3430 VDD.n506 185
R11747 VDD.n511 VDD.n506 185
R11748 VDD.n3429 VDD.n3428 185
R11749 VDD.n3428 VDD.n3427 185
R11750 VDD.n508 VDD.n507 185
R11751 VDD.n509 VDD.n508 185
R11752 VDD.n2929 VDD.n518 185
R11753 VDD.n3394 VDD.n518 185
R11754 VDD.n2931 VDD.n2930 185
R11755 VDD.n2930 VDD.n517 185
R11756 VDD.n2932 VDD.n542 185
R11757 VDD.n3336 VDD.n542 185
R11758 VDD.n2934 VDD.n2933 185
R11759 VDD.n2933 VDD.n541 185
R11760 VDD.n2935 VDD.n548 185
R11761 VDD.n3330 VDD.n548 185
R11762 VDD.n2937 VDD.n2936 185
R11763 VDD.n2936 VDD.n547 185
R11764 VDD.n2938 VDD.n554 185
R11765 VDD.n3322 VDD.n554 185
R11766 VDD.n2940 VDD.n2939 185
R11767 VDD.n2939 VDD.n562 185
R11768 VDD.n2941 VDD.n560 185
R11769 VDD.n3316 VDD.n560 185
R11770 VDD.n2943 VDD.n2942 185
R11771 VDD.n2942 VDD.n559 185
R11772 VDD.n2944 VDD.n567 185
R11773 VDD.n3310 VDD.n567 185
R11774 VDD.n2946 VDD.n2945 185
R11775 VDD.n2945 VDD.n566 185
R11776 VDD.n2947 VDD.n573 185
R11777 VDD.n3304 VDD.n573 185
R11778 VDD.n2949 VDD.n2948 185
R11779 VDD.n2948 VDD.n572 185
R11780 VDD.n2950 VDD.n579 185
R11781 VDD.n3298 VDD.n579 185
R11782 VDD.n2952 VDD.n2951 185
R11783 VDD.n2951 VDD.n578 185
R11784 VDD.n2953 VDD.n584 185
R11785 VDD.n3292 VDD.n584 185
R11786 VDD.n2955 VDD.n2954 185
R11787 VDD.n2956 VDD.n2955 185
R11788 VDD.n2928 VDD.n590 185
R11789 VDD.n3286 VDD.n590 185
R11790 VDD.n2927 VDD.n2926 185
R11791 VDD.n2926 VDD.n589 185
R11792 VDD.n2925 VDD.n596 185
R11793 VDD.n3280 VDD.n596 185
R11794 VDD.n2924 VDD.n2923 185
R11795 VDD.n2923 VDD.n595 185
R11796 VDD.n2922 VDD.n602 185
R11797 VDD.n3274 VDD.n602 185
R11798 VDD.n2921 VDD.n2920 185
R11799 VDD.n2920 VDD.n601 185
R11800 VDD.n2919 VDD.n608 185
R11801 VDD.n3268 VDD.n608 185
R11802 VDD.n2918 VDD.n2917 185
R11803 VDD.n2917 VDD.n607 185
R11804 VDD.n2916 VDD.n614 185
R11805 VDD.n3262 VDD.n614 185
R11806 VDD.n2915 VDD.n2914 185
R11807 VDD.n2914 VDD.n613 185
R11808 VDD.n2913 VDD.n620 185
R11809 VDD.n3256 VDD.n620 185
R11810 VDD.n2912 VDD.n2911 185
R11811 VDD.n2911 VDD.n619 185
R11812 VDD.n2910 VDD.n626 185
R11813 VDD.n3250 VDD.n626 185
R11814 VDD.n2909 VDD.n2908 185
R11815 VDD.n2908 VDD.n625 185
R11816 VDD.n2907 VDD.n632 185
R11817 VDD.n3244 VDD.n632 185
R11818 VDD.n2906 VDD.n2905 185
R11819 VDD.n2905 VDD.n631 185
R11820 VDD.n2904 VDD.n638 185
R11821 VDD.n3238 VDD.n638 185
R11822 VDD.n2903 VDD.n2902 185
R11823 VDD.n2902 VDD.n637 185
R11824 VDD.n2901 VDD.n644 185
R11825 VDD.n3232 VDD.n644 185
R11826 VDD.n2900 VDD.n2899 185
R11827 VDD.n2899 VDD.n643 185
R11828 VDD.n2898 VDD.n649 185
R11829 VDD.n3226 VDD.n649 185
R11830 VDD.n2897 VDD.n2896 185
R11831 VDD.n2896 VDD.n657 185
R11832 VDD.n2895 VDD.n655 185
R11833 VDD.n3220 VDD.n655 185
R11834 VDD.n2894 VDD.n2893 185
R11835 VDD.n2893 VDD.n654 185
R11836 VDD.n2892 VDD.n662 185
R11837 VDD.n3214 VDD.n662 185
R11838 VDD.n2891 VDD.n2890 185
R11839 VDD.n2890 VDD.n661 185
R11840 VDD.n2889 VDD.n668 185
R11841 VDD.n3208 VDD.n668 185
R11842 VDD.n2888 VDD.n2887 185
R11843 VDD.n2887 VDD.n667 185
R11844 VDD.n2886 VDD.n674 185
R11845 VDD.n3202 VDD.n674 185
R11846 VDD.n2885 VDD.n2884 185
R11847 VDD.n2884 VDD.n673 185
R11848 VDD.n2883 VDD.n680 185
R11849 VDD.n3196 VDD.n680 185
R11850 VDD.n2882 VDD.n2881 185
R11851 VDD.n2881 VDD.n679 185
R11852 VDD.n2880 VDD.n686 185
R11853 VDD.n3190 VDD.n686 185
R11854 VDD.n2879 VDD.n2878 185
R11855 VDD.n2878 VDD.n685 185
R11856 VDD.n2877 VDD.n692 185
R11857 VDD.n3184 VDD.n692 185
R11858 VDD.n2876 VDD.n2875 185
R11859 VDD.n2875 VDD.n691 185
R11860 VDD.n2874 VDD.n697 185
R11861 VDD.n3178 VDD.n697 185
R11862 VDD.n2873 VDD.n2872 185
R11863 VDD.n2872 VDD.n705 185
R11864 VDD.n2871 VDD.n703 185
R11865 VDD.n3172 VDD.n703 185
R11866 VDD.n2870 VDD.n2869 185
R11867 VDD.n2869 VDD.n702 185
R11868 VDD.n2868 VDD.n710 185
R11869 VDD.n3166 VDD.n710 185
R11870 VDD.n2867 VDD.n2866 185
R11871 VDD.n2866 VDD.n709 185
R11872 VDD.n2865 VDD.n716 185
R11873 VDD.n3160 VDD.n716 185
R11874 VDD.n2864 VDD.n2863 185
R11875 VDD.n2863 VDD.n715 185
R11876 VDD.n2862 VDD.n722 185
R11877 VDD.n3154 VDD.n722 185
R11878 VDD.n2861 VDD.n2860 185
R11879 VDD.n2860 VDD.n721 185
R11880 VDD.n2859 VDD.n728 185
R11881 VDD.n3148 VDD.n728 185
R11882 VDD.n2858 VDD.n2857 185
R11883 VDD.n2857 VDD.n727 185
R11884 VDD.n2856 VDD.n734 185
R11885 VDD.n3142 VDD.n734 185
R11886 VDD.n2855 VDD.n2854 185
R11887 VDD.n2854 VDD.n733 185
R11888 VDD.n2853 VDD.n740 185
R11889 VDD.n3136 VDD.n740 185
R11890 VDD.n2852 VDD.n2851 185
R11891 VDD.n2851 VDD.n739 185
R11892 VDD.n2850 VDD.n746 185
R11893 VDD.n3130 VDD.n746 185
R11894 VDD.n2849 VDD.n2848 185
R11895 VDD.n2848 VDD.n745 185
R11896 VDD.n2847 VDD.n752 185
R11897 VDD.n3124 VDD.n752 185
R11898 VDD.n2846 VDD.n2845 185
R11899 VDD.n2845 VDD.n751 185
R11900 VDD.n2844 VDD.n758 185
R11901 VDD.n3118 VDD.n758 185
R11902 VDD.n2843 VDD.n2842 185
R11903 VDD.n2842 VDD.n757 185
R11904 VDD.n2841 VDD.n764 185
R11905 VDD.n3112 VDD.n764 185
R11906 VDD.n2840 VDD.n2839 185
R11907 VDD.n2839 VDD.n763 185
R11908 VDD.n2838 VDD.n770 185
R11909 VDD.n3106 VDD.n770 185
R11910 VDD.n2837 VDD.n2836 185
R11911 VDD.n2836 VDD.n769 185
R11912 VDD.n2835 VDD.n2745 185
R11913 VDD.n3100 VDD.n2745 185
R11914 VDD.n3102 VDD.n3101 185
R11915 VDD.n3101 VDD.n3100 185
R11916 VDD.n3103 VDD.n772 185
R11917 VDD.n772 VDD.n769 185
R11918 VDD.n3105 VDD.n3104 185
R11919 VDD.n3106 VDD.n3105 185
R11920 VDD.n762 VDD.n761 185
R11921 VDD.n763 VDD.n762 185
R11922 VDD.n3114 VDD.n3113 185
R11923 VDD.n3113 VDD.n3112 185
R11924 VDD.n3115 VDD.n760 185
R11925 VDD.n760 VDD.n757 185
R11926 VDD.n3117 VDD.n3116 185
R11927 VDD.n3118 VDD.n3117 185
R11928 VDD.n750 VDD.n749 185
R11929 VDD.n751 VDD.n750 185
R11930 VDD.n3126 VDD.n3125 185
R11931 VDD.n3125 VDD.n3124 185
R11932 VDD.n3127 VDD.n748 185
R11933 VDD.n748 VDD.n745 185
R11934 VDD.n3129 VDD.n3128 185
R11935 VDD.n3130 VDD.n3129 185
R11936 VDD.n738 VDD.n737 185
R11937 VDD.n739 VDD.n738 185
R11938 VDD.n3138 VDD.n3137 185
R11939 VDD.n3137 VDD.n3136 185
R11940 VDD.n3139 VDD.n736 185
R11941 VDD.n736 VDD.n733 185
R11942 VDD.n3141 VDD.n3140 185
R11943 VDD.n3142 VDD.n3141 185
R11944 VDD.n726 VDD.n725 185
R11945 VDD.n727 VDD.n726 185
R11946 VDD.n3150 VDD.n3149 185
R11947 VDD.n3149 VDD.n3148 185
R11948 VDD.n3151 VDD.n724 185
R11949 VDD.n724 VDD.n721 185
R11950 VDD.n3153 VDD.n3152 185
R11951 VDD.n3154 VDD.n3153 185
R11952 VDD.n714 VDD.n713 185
R11953 VDD.n715 VDD.n714 185
R11954 VDD.n3162 VDD.n3161 185
R11955 VDD.n3161 VDD.n3160 185
R11956 VDD.n3163 VDD.n712 185
R11957 VDD.n712 VDD.n709 185
R11958 VDD.n3165 VDD.n3164 185
R11959 VDD.n3166 VDD.n3165 185
R11960 VDD.n701 VDD.n700 185
R11961 VDD.n702 VDD.n701 185
R11962 VDD.n3174 VDD.n3173 185
R11963 VDD.n3173 VDD.n3172 185
R11964 VDD.n3175 VDD.n699 185
R11965 VDD.n705 VDD.n699 185
R11966 VDD.n3177 VDD.n3176 185
R11967 VDD.n3178 VDD.n3177 185
R11968 VDD.n690 VDD.n689 185
R11969 VDD.n691 VDD.n690 185
R11970 VDD.n3186 VDD.n3185 185
R11971 VDD.n3185 VDD.n3184 185
R11972 VDD.n3187 VDD.n688 185
R11973 VDD.n688 VDD.n685 185
R11974 VDD.n3189 VDD.n3188 185
R11975 VDD.n3190 VDD.n3189 185
R11976 VDD.n678 VDD.n677 185
R11977 VDD.n679 VDD.n678 185
R11978 VDD.n3198 VDD.n3197 185
R11979 VDD.n3197 VDD.n3196 185
R11980 VDD.n3199 VDD.n676 185
R11981 VDD.n676 VDD.n673 185
R11982 VDD.n3201 VDD.n3200 185
R11983 VDD.n3202 VDD.n3201 185
R11984 VDD.n666 VDD.n665 185
R11985 VDD.n667 VDD.n666 185
R11986 VDD.n3210 VDD.n3209 185
R11987 VDD.n3209 VDD.n3208 185
R11988 VDD.n3211 VDD.n664 185
R11989 VDD.n664 VDD.n661 185
R11990 VDD.n3213 VDD.n3212 185
R11991 VDD.n3214 VDD.n3213 185
R11992 VDD.n653 VDD.n652 185
R11993 VDD.n654 VDD.n653 185
R11994 VDD.n3222 VDD.n3221 185
R11995 VDD.n3221 VDD.n3220 185
R11996 VDD.n3223 VDD.n651 185
R11997 VDD.n657 VDD.n651 185
R11998 VDD.n3225 VDD.n3224 185
R11999 VDD.n3226 VDD.n3225 185
R12000 VDD.n642 VDD.n641 185
R12001 VDD.n643 VDD.n642 185
R12002 VDD.n3234 VDD.n3233 185
R12003 VDD.n3233 VDD.n3232 185
R12004 VDD.n3235 VDD.n640 185
R12005 VDD.n640 VDD.n637 185
R12006 VDD.n3237 VDD.n3236 185
R12007 VDD.n3238 VDD.n3237 185
R12008 VDD.n630 VDD.n629 185
R12009 VDD.n631 VDD.n630 185
R12010 VDD.n3246 VDD.n3245 185
R12011 VDD.n3245 VDD.n3244 185
R12012 VDD.n3247 VDD.n628 185
R12013 VDD.n628 VDD.n625 185
R12014 VDD.n3249 VDD.n3248 185
R12015 VDD.n3250 VDD.n3249 185
R12016 VDD.n618 VDD.n617 185
R12017 VDD.n619 VDD.n618 185
R12018 VDD.n3258 VDD.n3257 185
R12019 VDD.n3257 VDD.n3256 185
R12020 VDD.n3259 VDD.n616 185
R12021 VDD.n616 VDD.n613 185
R12022 VDD.n3261 VDD.n3260 185
R12023 VDD.n3262 VDD.n3261 185
R12024 VDD.n606 VDD.n605 185
R12025 VDD.n607 VDD.n606 185
R12026 VDD.n3270 VDD.n3269 185
R12027 VDD.n3269 VDD.n3268 185
R12028 VDD.n3271 VDD.n604 185
R12029 VDD.n604 VDD.n601 185
R12030 VDD.n3273 VDD.n3272 185
R12031 VDD.n3274 VDD.n3273 185
R12032 VDD.n594 VDD.n593 185
R12033 VDD.n595 VDD.n594 185
R12034 VDD.n3282 VDD.n3281 185
R12035 VDD.n3281 VDD.n3280 185
R12036 VDD.n3283 VDD.n592 185
R12037 VDD.n592 VDD.n589 185
R12038 VDD.n3285 VDD.n3284 185
R12039 VDD.n3286 VDD.n3285 185
R12040 VDD.n583 VDD.n582 185
R12041 VDD.n2956 VDD.n583 185
R12042 VDD.n3294 VDD.n3293 185
R12043 VDD.n3293 VDD.n3292 185
R12044 VDD.n3295 VDD.n581 185
R12045 VDD.n581 VDD.n578 185
R12046 VDD.n3297 VDD.n3296 185
R12047 VDD.n3298 VDD.n3297 185
R12048 VDD.n571 VDD.n570 185
R12049 VDD.n572 VDD.n571 185
R12050 VDD.n3306 VDD.n3305 185
R12051 VDD.n3305 VDD.n3304 185
R12052 VDD.n3307 VDD.n569 185
R12053 VDD.n569 VDD.n566 185
R12054 VDD.n3309 VDD.n3308 185
R12055 VDD.n3310 VDD.n3309 185
R12056 VDD.n558 VDD.n557 185
R12057 VDD.n559 VDD.n558 185
R12058 VDD.n3318 VDD.n3317 185
R12059 VDD.n3317 VDD.n3316 185
R12060 VDD.n3319 VDD.n556 185
R12061 VDD.n562 VDD.n556 185
R12062 VDD.n3321 VDD.n3320 185
R12063 VDD.n3322 VDD.n3321 185
R12064 VDD.n546 VDD.n545 185
R12065 VDD.n547 VDD.n546 185
R12066 VDD.n3332 VDD.n3331 185
R12067 VDD.n3331 VDD.n3330 185
R12068 VDD.n3333 VDD.n544 185
R12069 VDD.n544 VDD.n541 185
R12070 VDD.n3335 VDD.n3334 185
R12071 VDD.n3336 VDD.n3335 185
R12072 VDD.n516 VDD.n515 185
R12073 VDD.n517 VDD.n516 185
R12074 VDD.n3396 VDD.n3395 185
R12075 VDD.n3395 VDD.n3394 185
R12076 VDD.n3397 VDD.n513 185
R12077 VDD.n513 VDD.n509 185
R12078 VDD.n3426 VDD.n3425 185
R12079 VDD.n3427 VDD.n3426 185
R12080 VDD.n3424 VDD.n514 185
R12081 VDD.n514 VDD.n511 185
R12082 VDD.n800 VDD.n798 185
R12083 VDD.n798 VDD.n775 185
R12084 VDD.n2629 VDD.n807 185
R12085 VDD.n2696 VDD.n807 185
R12086 VDD.n2631 VDD.n2630 185
R12087 VDD.n2630 VDD.n805 185
R12088 VDD.n2632 VDD.n818 185
R12089 VDD.n2642 VDD.n818 185
R12090 VDD.n2633 VDD.n826 185
R12091 VDD.n826 VDD.n816 185
R12092 VDD.n2635 VDD.n2634 185
R12093 VDD.n2636 VDD.n2635 185
R12094 VDD.n2628 VDD.n825 185
R12095 VDD.n825 VDD.n822 185
R12096 VDD.n2627 VDD.n2626 185
R12097 VDD.n2626 VDD.n2625 185
R12098 VDD.n828 VDD.n827 185
R12099 VDD.n829 VDD.n828 185
R12100 VDD.n2618 VDD.n2617 185
R12101 VDD.n2619 VDD.n2618 185
R12102 VDD.n2616 VDD.n838 185
R12103 VDD.n838 VDD.n835 185
R12104 VDD.n2615 VDD.n2614 185
R12105 VDD.n2614 VDD.n2613 185
R12106 VDD.n840 VDD.n839 185
R12107 VDD.n841 VDD.n840 185
R12108 VDD.n2606 VDD.n2605 185
R12109 VDD.n2607 VDD.n2606 185
R12110 VDD.n2604 VDD.n850 185
R12111 VDD.n850 VDD.n847 185
R12112 VDD.n2603 VDD.n2602 185
R12113 VDD.n2602 VDD.n2601 185
R12114 VDD.n852 VDD.n851 185
R12115 VDD.n853 VDD.n852 185
R12116 VDD.n2594 VDD.n2593 185
R12117 VDD.n2595 VDD.n2594 185
R12118 VDD.n2592 VDD.n862 185
R12119 VDD.n862 VDD.n859 185
R12120 VDD.n2591 VDD.n2590 185
R12121 VDD.n2590 VDD.n2589 185
R12122 VDD.n864 VDD.n863 185
R12123 VDD.n865 VDD.n864 185
R12124 VDD.n2582 VDD.n2581 185
R12125 VDD.n2583 VDD.n2582 185
R12126 VDD.n2580 VDD.n874 185
R12127 VDD.n874 VDD.n871 185
R12128 VDD.n2579 VDD.n2578 185
R12129 VDD.n2578 VDD.n2577 185
R12130 VDD.n876 VDD.n875 185
R12131 VDD.n877 VDD.n876 185
R12132 VDD.n2570 VDD.n2569 185
R12133 VDD.n2571 VDD.n2570 185
R12134 VDD.n2568 VDD.n885 185
R12135 VDD.n891 VDD.n885 185
R12136 VDD.n2567 VDD.n2566 185
R12137 VDD.n2566 VDD.n2565 185
R12138 VDD.n887 VDD.n886 185
R12139 VDD.n888 VDD.n887 185
R12140 VDD.n2558 VDD.n2557 185
R12141 VDD.n2559 VDD.n2558 185
R12142 VDD.n2556 VDD.n898 185
R12143 VDD.n898 VDD.n895 185
R12144 VDD.n2555 VDD.n2554 185
R12145 VDD.n2554 VDD.n2553 185
R12146 VDD.n900 VDD.n899 185
R12147 VDD.n901 VDD.n900 185
R12148 VDD.n2546 VDD.n2545 185
R12149 VDD.n2547 VDD.n2546 185
R12150 VDD.n2544 VDD.n910 185
R12151 VDD.n910 VDD.n907 185
R12152 VDD.n2543 VDD.n2542 185
R12153 VDD.n2542 VDD.n2541 185
R12154 VDD.n912 VDD.n911 185
R12155 VDD.n913 VDD.n912 185
R12156 VDD.n2534 VDD.n2533 185
R12157 VDD.n2535 VDD.n2534 185
R12158 VDD.n2532 VDD.n922 185
R12159 VDD.n922 VDD.n919 185
R12160 VDD.n2531 VDD.n2530 185
R12161 VDD.n2530 VDD.n2529 185
R12162 VDD.n924 VDD.n923 185
R12163 VDD.n925 VDD.n924 185
R12164 VDD.n2522 VDD.n2521 185
R12165 VDD.n2523 VDD.n2522 185
R12166 VDD.n2520 VDD.n933 185
R12167 VDD.n939 VDD.n933 185
R12168 VDD.n2519 VDD.n2518 185
R12169 VDD.n2518 VDD.n2517 185
R12170 VDD.n935 VDD.n934 185
R12171 VDD.n936 VDD.n935 185
R12172 VDD.n2510 VDD.n2509 185
R12173 VDD.n2511 VDD.n2510 185
R12174 VDD.n2508 VDD.n946 185
R12175 VDD.n946 VDD.n943 185
R12176 VDD.n2507 VDD.n2506 185
R12177 VDD.n2506 VDD.n2505 185
R12178 VDD.n948 VDD.n947 185
R12179 VDD.n949 VDD.n948 185
R12180 VDD.n2498 VDD.n2497 185
R12181 VDD.n2499 VDD.n2498 185
R12182 VDD.n2496 VDD.n958 185
R12183 VDD.n958 VDD.n955 185
R12184 VDD.n2495 VDD.n2494 185
R12185 VDD.n2494 VDD.n2493 185
R12186 VDD.n960 VDD.n959 185
R12187 VDD.n961 VDD.n960 185
R12188 VDD.n2486 VDD.n2485 185
R12189 VDD.n2487 VDD.n2486 185
R12190 VDD.n2484 VDD.n970 185
R12191 VDD.n970 VDD.n967 185
R12192 VDD.n2483 VDD.n2482 185
R12193 VDD.n2482 VDD.n2481 185
R12194 VDD.n972 VDD.n971 185
R12195 VDD.n973 VDD.n972 185
R12196 VDD.n2474 VDD.n2473 185
R12197 VDD.n2475 VDD.n2474 185
R12198 VDD.n2472 VDD.n982 185
R12199 VDD.n982 VDD.n979 185
R12200 VDD.n2471 VDD.n2470 185
R12201 VDD.n2470 VDD.n2469 185
R12202 VDD.n984 VDD.n983 185
R12203 VDD.n985 VDD.n984 185
R12204 VDD.n2462 VDD.n2461 185
R12205 VDD.n2463 VDD.n2462 185
R12206 VDD.n2460 VDD.n994 185
R12207 VDD.n994 VDD.n991 185
R12208 VDD.n2459 VDD.n2458 185
R12209 VDD.n2458 VDD.n2457 185
R12210 VDD.n996 VDD.n995 185
R12211 VDD.n1005 VDD.n996 185
R12212 VDD.n2450 VDD.n2449 185
R12213 VDD.n2451 VDD.n2450 185
R12214 VDD.n2448 VDD.n1006 185
R12215 VDD.n1006 VDD.n1002 185
R12216 VDD.n2447 VDD.n2446 185
R12217 VDD.n2446 VDD.n2445 185
R12218 VDD.n1008 VDD.n1007 185
R12219 VDD.n1009 VDD.n1008 185
R12220 VDD.n2438 VDD.n2437 185
R12221 VDD.n2439 VDD.n2438 185
R12222 VDD.n2436 VDD.n1018 185
R12223 VDD.n1018 VDD.n1015 185
R12224 VDD.n2435 VDD.n2434 185
R12225 VDD.n2434 VDD.n2433 185
R12226 VDD.n1020 VDD.n1019 185
R12227 VDD.n1021 VDD.n1020 185
R12228 VDD.n2426 VDD.n2425 185
R12229 VDD.n2427 VDD.n2426 185
R12230 VDD.n2424 VDD.n1029 185
R12231 VDD.n1035 VDD.n1029 185
R12232 VDD.n2423 VDD.n2422 185
R12233 VDD.n2422 VDD.n2421 185
R12234 VDD.n1031 VDD.n1030 185
R12235 VDD.n1032 VDD.n1031 185
R12236 VDD.n2414 VDD.n2413 185
R12237 VDD.n2415 VDD.n2414 185
R12238 VDD.n2412 VDD.n1042 185
R12239 VDD.n1042 VDD.n1039 185
R12240 VDD.n2411 VDD.n2410 185
R12241 VDD.n2410 VDD.n2409 185
R12242 VDD.n1044 VDD.n1043 185
R12243 VDD.n1045 VDD.n1044 185
R12244 VDD.n2402 VDD.n2401 185
R12245 VDD.n2403 VDD.n2402 185
R12246 VDD.n2400 VDD.n1054 185
R12247 VDD.n1054 VDD.n1051 185
R12248 VDD.n2399 VDD.n2398 185
R12249 VDD.n2398 VDD.n2397 185
R12250 VDD.n2700 VDD.n797 185
R12251 VDD.n2743 VDD.n797 185
R12252 VDD.n2702 VDD.n2701 185
R12253 VDD.n2705 VDD.n2704 185
R12254 VDD.n2707 VDD.n2706 185
R12255 VDD.n2709 VDD.n2708 185
R12256 VDD.n2711 VDD.n2710 185
R12257 VDD.n2713 VDD.n2712 185
R12258 VDD.n2715 VDD.n2714 185
R12259 VDD.n2717 VDD.n2716 185
R12260 VDD.n2719 VDD.n2718 185
R12261 VDD.n2721 VDD.n2720 185
R12262 VDD.n2723 VDD.n2722 185
R12263 VDD.n2725 VDD.n2724 185
R12264 VDD.n2727 VDD.n2726 185
R12265 VDD.n2729 VDD.n2728 185
R12266 VDD.n2731 VDD.n2730 185
R12267 VDD.n2733 VDD.n2732 185
R12268 VDD.n2735 VDD.n2734 185
R12269 VDD.n2737 VDD.n2736 185
R12270 VDD.n2739 VDD.n2738 185
R12271 VDD.n2740 VDD.n799 185
R12272 VDD.n2742 VDD.n2741 185
R12273 VDD.n2743 VDD.n2742 185
R12274 VDD.n2699 VDD.n2698 185
R12275 VDD.n2698 VDD.n775 185
R12276 VDD.n2697 VDD.n803 185
R12277 VDD.n2697 VDD.n2696 185
R12278 VDD.n2266 VDD.n804 185
R12279 VDD.n805 VDD.n804 185
R12280 VDD.n2267 VDD.n817 185
R12281 VDD.n2642 VDD.n817 185
R12282 VDD.n2269 VDD.n2268 185
R12283 VDD.n2268 VDD.n816 185
R12284 VDD.n2270 VDD.n824 185
R12285 VDD.n2636 VDD.n824 185
R12286 VDD.n2272 VDD.n2271 185
R12287 VDD.n2271 VDD.n822 185
R12288 VDD.n2273 VDD.n831 185
R12289 VDD.n2625 VDD.n831 185
R12290 VDD.n2275 VDD.n2274 185
R12291 VDD.n2274 VDD.n829 185
R12292 VDD.n2276 VDD.n837 185
R12293 VDD.n2619 VDD.n837 185
R12294 VDD.n2278 VDD.n2277 185
R12295 VDD.n2277 VDD.n835 185
R12296 VDD.n2279 VDD.n843 185
R12297 VDD.n2613 VDD.n843 185
R12298 VDD.n2281 VDD.n2280 185
R12299 VDD.n2280 VDD.n841 185
R12300 VDD.n2282 VDD.n849 185
R12301 VDD.n2607 VDD.n849 185
R12302 VDD.n2284 VDD.n2283 185
R12303 VDD.n2283 VDD.n847 185
R12304 VDD.n2285 VDD.n855 185
R12305 VDD.n2601 VDD.n855 185
R12306 VDD.n2287 VDD.n2286 185
R12307 VDD.n2286 VDD.n853 185
R12308 VDD.n2288 VDD.n861 185
R12309 VDD.n2595 VDD.n861 185
R12310 VDD.n2290 VDD.n2289 185
R12311 VDD.n2289 VDD.n859 185
R12312 VDD.n2291 VDD.n867 185
R12313 VDD.n2589 VDD.n867 185
R12314 VDD.n2293 VDD.n2292 185
R12315 VDD.n2292 VDD.n865 185
R12316 VDD.n2294 VDD.n873 185
R12317 VDD.n2583 VDD.n873 185
R12318 VDD.n2296 VDD.n2295 185
R12319 VDD.n2295 VDD.n871 185
R12320 VDD.n2297 VDD.n879 185
R12321 VDD.n2577 VDD.n879 185
R12322 VDD.n2299 VDD.n2298 185
R12323 VDD.n2298 VDD.n877 185
R12324 VDD.n2300 VDD.n884 185
R12325 VDD.n2571 VDD.n884 185
R12326 VDD.n2302 VDD.n2301 185
R12327 VDD.n2301 VDD.n891 185
R12328 VDD.n2303 VDD.n890 185
R12329 VDD.n2565 VDD.n890 185
R12330 VDD.n2305 VDD.n2304 185
R12331 VDD.n2304 VDD.n888 185
R12332 VDD.n2306 VDD.n897 185
R12333 VDD.n2559 VDD.n897 185
R12334 VDD.n2308 VDD.n2307 185
R12335 VDD.n2307 VDD.n895 185
R12336 VDD.n2309 VDD.n903 185
R12337 VDD.n2553 VDD.n903 185
R12338 VDD.n2311 VDD.n2310 185
R12339 VDD.n2310 VDD.n901 185
R12340 VDD.n2312 VDD.n909 185
R12341 VDD.n2547 VDD.n909 185
R12342 VDD.n2314 VDD.n2313 185
R12343 VDD.n2313 VDD.n907 185
R12344 VDD.n2315 VDD.n915 185
R12345 VDD.n2541 VDD.n915 185
R12346 VDD.n2317 VDD.n2316 185
R12347 VDD.n2316 VDD.n913 185
R12348 VDD.n2318 VDD.n921 185
R12349 VDD.n2535 VDD.n921 185
R12350 VDD.n2320 VDD.n2319 185
R12351 VDD.n2319 VDD.n919 185
R12352 VDD.n2321 VDD.n927 185
R12353 VDD.n2529 VDD.n927 185
R12354 VDD.n2323 VDD.n2322 185
R12355 VDD.n2322 VDD.n925 185
R12356 VDD.n2324 VDD.n932 185
R12357 VDD.n2523 VDD.n932 185
R12358 VDD.n2326 VDD.n2325 185
R12359 VDD.n2325 VDD.n939 185
R12360 VDD.n2327 VDD.n938 185
R12361 VDD.n2517 VDD.n938 185
R12362 VDD.n2329 VDD.n2328 185
R12363 VDD.n2328 VDD.n936 185
R12364 VDD.n2330 VDD.n945 185
R12365 VDD.n2511 VDD.n945 185
R12366 VDD.n2332 VDD.n2331 185
R12367 VDD.n2331 VDD.n943 185
R12368 VDD.n2333 VDD.n951 185
R12369 VDD.n2505 VDD.n951 185
R12370 VDD.n2335 VDD.n2334 185
R12371 VDD.n2334 VDD.n949 185
R12372 VDD.n2336 VDD.n957 185
R12373 VDD.n2499 VDD.n957 185
R12374 VDD.n2338 VDD.n2337 185
R12375 VDD.n2337 VDD.n955 185
R12376 VDD.n2339 VDD.n963 185
R12377 VDD.n2493 VDD.n963 185
R12378 VDD.n2341 VDD.n2340 185
R12379 VDD.n2340 VDD.n961 185
R12380 VDD.n2342 VDD.n969 185
R12381 VDD.n2487 VDD.n969 185
R12382 VDD.n2344 VDD.n2343 185
R12383 VDD.n2343 VDD.n967 185
R12384 VDD.n2345 VDD.n975 185
R12385 VDD.n2481 VDD.n975 185
R12386 VDD.n2347 VDD.n2346 185
R12387 VDD.n2346 VDD.n973 185
R12388 VDD.n2348 VDD.n981 185
R12389 VDD.n2475 VDD.n981 185
R12390 VDD.n2350 VDD.n2349 185
R12391 VDD.n2349 VDD.n979 185
R12392 VDD.n2351 VDD.n987 185
R12393 VDD.n2469 VDD.n987 185
R12394 VDD.n2353 VDD.n2352 185
R12395 VDD.n2352 VDD.n985 185
R12396 VDD.n2354 VDD.n993 185
R12397 VDD.n2463 VDD.n993 185
R12398 VDD.n2356 VDD.n2355 185
R12399 VDD.n2355 VDD.n991 185
R12400 VDD.n2357 VDD.n998 185
R12401 VDD.n2457 VDD.n998 185
R12402 VDD.n2359 VDD.n2358 185
R12403 VDD.n2358 VDD.n1005 185
R12404 VDD.n2360 VDD.n1004 185
R12405 VDD.n2451 VDD.n1004 185
R12406 VDD.n2362 VDD.n2361 185
R12407 VDD.n2361 VDD.n1002 185
R12408 VDD.n2363 VDD.n1011 185
R12409 VDD.n2445 VDD.n1011 185
R12410 VDD.n2365 VDD.n2364 185
R12411 VDD.n2364 VDD.n1009 185
R12412 VDD.n2366 VDD.n1017 185
R12413 VDD.n2439 VDD.n1017 185
R12414 VDD.n2368 VDD.n2367 185
R12415 VDD.n2367 VDD.n1015 185
R12416 VDD.n2369 VDD.n1023 185
R12417 VDD.n2433 VDD.n1023 185
R12418 VDD.n2371 VDD.n2370 185
R12419 VDD.n2370 VDD.n1021 185
R12420 VDD.n2372 VDD.n1028 185
R12421 VDD.n2427 VDD.n1028 185
R12422 VDD.n2374 VDD.n2373 185
R12423 VDD.n2373 VDD.n1035 185
R12424 VDD.n2375 VDD.n1034 185
R12425 VDD.n2421 VDD.n1034 185
R12426 VDD.n2377 VDD.n2376 185
R12427 VDD.n2376 VDD.n1032 185
R12428 VDD.n2378 VDD.n1041 185
R12429 VDD.n2415 VDD.n1041 185
R12430 VDD.n2380 VDD.n2379 185
R12431 VDD.n2379 VDD.n1039 185
R12432 VDD.n2381 VDD.n1047 185
R12433 VDD.n2409 VDD.n1047 185
R12434 VDD.n2383 VDD.n2382 185
R12435 VDD.n2382 VDD.n1045 185
R12436 VDD.n2384 VDD.n1053 185
R12437 VDD.n2403 VDD.n1053 185
R12438 VDD.n2386 VDD.n2385 185
R12439 VDD.n2385 VDD.n1051 185
R12440 VDD.n2387 VDD.n1058 185
R12441 VDD.n2397 VDD.n1058 185
R12442 VDD.n1056 VDD.n1055 185
R12443 VDD.n2390 VDD.n1056 185
R12444 VDD.n2227 VDD.n2226 185
R12445 VDD.n2229 VDD.n2228 185
R12446 VDD.n2231 VDD.n2230 185
R12447 VDD.n2233 VDD.n2232 185
R12448 VDD.n2235 VDD.n2234 185
R12449 VDD.n2237 VDD.n2236 185
R12450 VDD.n2239 VDD.n2238 185
R12451 VDD.n2241 VDD.n2240 185
R12452 VDD.n2243 VDD.n2242 185
R12453 VDD.n2245 VDD.n2244 185
R12454 VDD.n2247 VDD.n2246 185
R12455 VDD.n2249 VDD.n2248 185
R12456 VDD.n2251 VDD.n2250 185
R12457 VDD.n2253 VDD.n2252 185
R12458 VDD.n2255 VDD.n2254 185
R12459 VDD.n2257 VDD.n2256 185
R12460 VDD.n2259 VDD.n2258 185
R12461 VDD.n2261 VDD.n2260 185
R12462 VDD.n2263 VDD.n2262 185
R12463 VDD.n2265 VDD.n1082 185
R12464 VDD.n2389 VDD.n2388 185
R12465 VDD.n2390 VDD.n2389 185
R12466 VDD.n138 VDD.n137 171.744
R12467 VDD.n125 VDD.n124 171.744
R12468 VDD.n112 VDD.n111 171.744
R12469 VDD.n99 VDD.n98 171.744
R12470 VDD.n86 VDD.n85 171.744
R12471 VDD.n73 VDD.n72 171.744
R12472 VDD.n60 VDD.n59 171.744
R12473 VDD.n47 VDD.n46 171.744
R12474 VDD.n35 VDD.n34 171.744
R12475 VDD.n22 VDD.n21 171.744
R12476 VDD.n1731 VDD.n1730 171.744
R12477 VDD.n1744 VDD.n1743 171.744
R12478 VDD.n1705 VDD.n1704 171.744
R12479 VDD.n1718 VDD.n1717 171.744
R12480 VDD.n1679 VDD.n1678 171.744
R12481 VDD.n1692 VDD.n1691 171.744
R12482 VDD.n1653 VDD.n1652 171.744
R12483 VDD.n1666 VDD.n1665 171.744
R12484 VDD.n1628 VDD.n1627 171.744
R12485 VDD.n1641 VDD.n1640 171.744
R12486 VDD.n2390 VDD.t26 158.333
R12487 VDD.n496 VDD.t25 158.333
R12488 VDD.n3875 VDD.n3874 146.341
R12489 VDD.n3872 VDD.n250 146.341
R12490 VDD.n3868 VDD.n3867 146.341
R12491 VDD.n3865 VDD.n257 146.341
R12492 VDD.n3859 VDD.n3858 146.341
R12493 VDD.n3856 VDD.n265 146.341
R12494 VDD.n3852 VDD.n3851 146.341
R12495 VDD.n3849 VDD.n271 146.341
R12496 VDD.n3842 VDD.n280 146.341
R12497 VDD.n3840 VDD.n3839 146.341
R12498 VDD.n3837 VDD.n282 146.341
R12499 VDD.n3833 VDD.n3832 146.341
R12500 VDD.n3830 VDD.n289 146.341
R12501 VDD.n3823 VDD.n3822 146.341
R12502 VDD.n3820 VDD.n296 146.341
R12503 VDD.n3816 VDD.n3815 146.341
R12504 VDD.n3813 VDD.n303 146.341
R12505 VDD.n314 VDD.n311 146.341
R12506 VDD.n3805 VDD.n3804 146.341
R12507 VDD.n3802 VDD.n316 146.341
R12508 VDD.n3798 VDD.n3797 146.341
R12509 VDD.n3795 VDD.n322 146.341
R12510 VDD.n3579 VDD.n442 146.341
R12511 VDD.n3589 VDD.n442 146.341
R12512 VDD.n3589 VDD.n438 146.341
R12513 VDD.n3595 VDD.n438 146.341
R12514 VDD.n3595 VDD.n431 146.341
R12515 VDD.n3606 VDD.n431 146.341
R12516 VDD.n3606 VDD.n427 146.341
R12517 VDD.n3612 VDD.n427 146.341
R12518 VDD.n3612 VDD.n419 146.341
R12519 VDD.n3622 VDD.n419 146.341
R12520 VDD.n3622 VDD.n415 146.341
R12521 VDD.n3628 VDD.n415 146.341
R12522 VDD.n3628 VDD.n407 146.341
R12523 VDD.n3638 VDD.n407 146.341
R12524 VDD.n3638 VDD.n403 146.341
R12525 VDD.n3644 VDD.n403 146.341
R12526 VDD.n3644 VDD.n395 146.341
R12527 VDD.n3654 VDD.n395 146.341
R12528 VDD.n3654 VDD.n391 146.341
R12529 VDD.n3660 VDD.n391 146.341
R12530 VDD.n3660 VDD.n383 146.341
R12531 VDD.n3670 VDD.n383 146.341
R12532 VDD.n3670 VDD.n379 146.341
R12533 VDD.n3676 VDD.n379 146.341
R12534 VDD.n3676 VDD.n371 146.341
R12535 VDD.n3686 VDD.n371 146.341
R12536 VDD.n3686 VDD.n367 146.341
R12537 VDD.n3692 VDD.n367 146.341
R12538 VDD.n3692 VDD.n360 146.341
R12539 VDD.n3703 VDD.n360 146.341
R12540 VDD.n3703 VDD.n356 146.341
R12541 VDD.n3712 VDD.n356 146.341
R12542 VDD.n3712 VDD.n348 146.341
R12543 VDD.n3722 VDD.n348 146.341
R12544 VDD.n3723 VDD.n3722 146.341
R12545 VDD.n3723 VDD.n152 146.341
R12546 VDD.n153 VDD.n152 146.341
R12547 VDD.n154 VDD.n153 146.341
R12548 VDD.n3730 VDD.n154 146.341
R12549 VDD.n3730 VDD.n162 146.341
R12550 VDD.n163 VDD.n162 146.341
R12551 VDD.n164 VDD.n163 146.341
R12552 VDD.n3737 VDD.n164 146.341
R12553 VDD.n3737 VDD.n173 146.341
R12554 VDD.n174 VDD.n173 146.341
R12555 VDD.n175 VDD.n174 146.341
R12556 VDD.n3744 VDD.n175 146.341
R12557 VDD.n3744 VDD.n184 146.341
R12558 VDD.n185 VDD.n184 146.341
R12559 VDD.n186 VDD.n185 146.341
R12560 VDD.n3751 VDD.n186 146.341
R12561 VDD.n3751 VDD.n195 146.341
R12562 VDD.n196 VDD.n195 146.341
R12563 VDD.n197 VDD.n196 146.341
R12564 VDD.n3758 VDD.n197 146.341
R12565 VDD.n3758 VDD.n206 146.341
R12566 VDD.n207 VDD.n206 146.341
R12567 VDD.n208 VDD.n207 146.341
R12568 VDD.n3765 VDD.n208 146.341
R12569 VDD.n3765 VDD.n217 146.341
R12570 VDD.n218 VDD.n217 146.341
R12571 VDD.n219 VDD.n218 146.341
R12572 VDD.n3772 VDD.n219 146.341
R12573 VDD.n3772 VDD.n228 146.341
R12574 VDD.n229 VDD.n228 146.341
R12575 VDD.n230 VDD.n229 146.341
R12576 VDD.n3779 VDD.n230 146.341
R12577 VDD.n3779 VDD.n239 146.341
R12578 VDD.n240 VDD.n239 146.341
R12579 VDD.n241 VDD.n240 146.341
R12580 VDD.n3787 VDD.n241 146.341
R12581 VDD.n3466 VDD.n3465 146.341
R12582 VDD.n3468 VDD.n3466 146.341
R12583 VDD.n3473 VDD.n3458 146.341
R12584 VDD.n3475 VDD.n3454 146.341
R12585 VDD.n3482 VDD.n491 146.341
R12586 VDD.n3486 VDD.n3484 146.341
R12587 VDD.n3492 VDD.n487 146.341
R12588 VDD.n3496 VDD.n3494 146.341
R12589 VDD.n3502 VDD.n481 146.341
R12590 VDD.n3506 VDD.n3504 146.341
R12591 VDD.n3512 VDD.n477 146.341
R12592 VDD.n3516 VDD.n3514 146.341
R12593 VDD.n3525 VDD.n473 146.341
R12594 VDD.n3529 VDD.n3527 146.341
R12595 VDD.n3535 VDD.n469 146.341
R12596 VDD.n3539 VDD.n3537 146.341
R12597 VDD.n3545 VDD.n465 146.341
R12598 VDD.n3549 VDD.n3547 146.341
R12599 VDD.n3557 VDD.n461 146.341
R12600 VDD.n3561 VDD.n3559 146.341
R12601 VDD.n3567 VDD.n455 146.341
R12602 VDD.n3570 VDD.n3569 146.341
R12603 VDD.n3572 VDD.n449 146.341
R12604 VDD.n3581 VDD.n444 146.341
R12605 VDD.n3587 VDD.n444 146.341
R12606 VDD.n3587 VDD.n436 146.341
R12607 VDD.n3598 VDD.n436 146.341
R12608 VDD.n3598 VDD.n432 146.341
R12609 VDD.n3604 VDD.n432 146.341
R12610 VDD.n3604 VDD.n425 146.341
R12611 VDD.n3614 VDD.n425 146.341
R12612 VDD.n3614 VDD.n421 146.341
R12613 VDD.n3620 VDD.n421 146.341
R12614 VDD.n3620 VDD.n413 146.341
R12615 VDD.n3630 VDD.n413 146.341
R12616 VDD.n3630 VDD.n409 146.341
R12617 VDD.n3636 VDD.n409 146.341
R12618 VDD.n3636 VDD.n401 146.341
R12619 VDD.n3646 VDD.n401 146.341
R12620 VDD.n3646 VDD.n397 146.341
R12621 VDD.n3652 VDD.n397 146.341
R12622 VDD.n3652 VDD.n389 146.341
R12623 VDD.n3662 VDD.n389 146.341
R12624 VDD.n3662 VDD.n385 146.341
R12625 VDD.n3668 VDD.n385 146.341
R12626 VDD.n3668 VDD.n377 146.341
R12627 VDD.n3678 VDD.n377 146.341
R12628 VDD.n3678 VDD.n373 146.341
R12629 VDD.n3684 VDD.n373 146.341
R12630 VDD.n3684 VDD.n365 146.341
R12631 VDD.n3695 VDD.n365 146.341
R12632 VDD.n3695 VDD.n361 146.341
R12633 VDD.n3701 VDD.n361 146.341
R12634 VDD.n3701 VDD.n354 146.341
R12635 VDD.n3714 VDD.n354 146.341
R12636 VDD.n3714 VDD.n350 146.341
R12637 VDD.n3720 VDD.n350 146.341
R12638 VDD.n3720 VDD.n149 146.341
R12639 VDD.n3951 VDD.n149 146.341
R12640 VDD.n3951 VDD.n150 146.341
R12641 VDD.n3947 VDD.n150 146.341
R12642 VDD.n3947 VDD.n156 146.341
R12643 VDD.n3943 VDD.n156 146.341
R12644 VDD.n3943 VDD.n161 146.341
R12645 VDD.n3939 VDD.n161 146.341
R12646 VDD.n3939 VDD.n166 146.341
R12647 VDD.n3935 VDD.n166 146.341
R12648 VDD.n3935 VDD.n172 146.341
R12649 VDD.n3931 VDD.n172 146.341
R12650 VDD.n3931 VDD.n177 146.341
R12651 VDD.n3927 VDD.n177 146.341
R12652 VDD.n3927 VDD.n183 146.341
R12653 VDD.n3923 VDD.n183 146.341
R12654 VDD.n3923 VDD.n188 146.341
R12655 VDD.n3919 VDD.n188 146.341
R12656 VDD.n3919 VDD.n194 146.341
R12657 VDD.n3915 VDD.n194 146.341
R12658 VDD.n3915 VDD.n199 146.341
R12659 VDD.n3911 VDD.n199 146.341
R12660 VDD.n3911 VDD.n205 146.341
R12661 VDD.n3907 VDD.n205 146.341
R12662 VDD.n3907 VDD.n210 146.341
R12663 VDD.n3903 VDD.n210 146.341
R12664 VDD.n3903 VDD.n216 146.341
R12665 VDD.n3899 VDD.n216 146.341
R12666 VDD.n3899 VDD.n221 146.341
R12667 VDD.n3895 VDD.n221 146.341
R12668 VDD.n3895 VDD.n227 146.341
R12669 VDD.n3891 VDD.n227 146.341
R12670 VDD.n3891 VDD.n232 146.341
R12671 VDD.n3887 VDD.n232 146.341
R12672 VDD.n3887 VDD.n238 146.341
R12673 VDD.n3883 VDD.n238 146.341
R12674 VDD.n3883 VDD.n243 146.341
R12675 VDD.n2205 VDD.n2204 146.341
R12676 VDD.n2202 VDD.n1900 146.341
R12677 VDD.n2035 VDD.n2034 146.341
R12678 VDD.n2032 VDD.n1905 146.341
R12679 VDD.n2023 VDD.n1910 146.341
R12680 VDD.n2021 VDD.n2020 146.341
R12681 VDD.n2018 VDD.n1912 146.341
R12682 VDD.n2014 VDD.n2013 146.341
R12683 VDD.n2011 VDD.n1921 146.341
R12684 VDD.n2007 VDD.n2006 146.341
R12685 VDD.n2004 VDD.n1928 146.341
R12686 VDD.n2000 VDD.n1999 146.341
R12687 VDD.n1997 VDD.n1935 146.341
R12688 VDD.n1990 VDD.n1989 146.341
R12689 VDD.n1987 VDD.n1942 146.341
R12690 VDD.n1983 VDD.n1982 146.341
R12691 VDD.n1980 VDD.n1949 146.341
R12692 VDD.n1959 VDD.n1957 146.341
R12693 VDD.n1972 VDD.n1971 146.341
R12694 VDD.n1969 VDD.n1967 146.341
R12695 VDD.n1965 VDD.n1963 146.341
R12696 VDD.n1091 VDD.n1090 146.341
R12697 VDD.n1487 VDD.n1309 146.341
R12698 VDD.n1487 VDD.n1301 146.341
R12699 VDD.n1497 VDD.n1301 146.341
R12700 VDD.n1497 VDD.n1297 146.341
R12701 VDD.n1503 VDD.n1297 146.341
R12702 VDD.n1503 VDD.n1289 146.341
R12703 VDD.n1513 VDD.n1289 146.341
R12704 VDD.n1513 VDD.n1285 146.341
R12705 VDD.n1519 VDD.n1285 146.341
R12706 VDD.n1519 VDD.n1277 146.341
R12707 VDD.n1529 VDD.n1277 146.341
R12708 VDD.n1529 VDD.n1273 146.341
R12709 VDD.n1535 VDD.n1273 146.341
R12710 VDD.n1535 VDD.n1265 146.341
R12711 VDD.n1545 VDD.n1265 146.341
R12712 VDD.n1545 VDD.n1261 146.341
R12713 VDD.n1551 VDD.n1261 146.341
R12714 VDD.n1551 VDD.n1254 146.341
R12715 VDD.n1562 VDD.n1254 146.341
R12716 VDD.n1562 VDD.n1250 146.341
R12717 VDD.n1568 VDD.n1250 146.341
R12718 VDD.n1568 VDD.n1242 146.341
R12719 VDD.n1578 VDD.n1242 146.341
R12720 VDD.n1578 VDD.n1238 146.341
R12721 VDD.n1584 VDD.n1238 146.341
R12722 VDD.n1584 VDD.n1230 146.341
R12723 VDD.n1594 VDD.n1230 146.341
R12724 VDD.n1594 VDD.n1226 146.341
R12725 VDD.n1600 VDD.n1226 146.341
R12726 VDD.n1600 VDD.n1218 146.341
R12727 VDD.n1610 VDD.n1218 146.341
R12728 VDD.n1610 VDD.n1214 146.341
R12729 VDD.n1616 VDD.n1214 146.341
R12730 VDD.n1616 VDD.n1206 146.341
R12731 VDD.n1757 VDD.n1206 146.341
R12732 VDD.n1757 VDD.n1202 146.341
R12733 VDD.n1763 VDD.n1202 146.341
R12734 VDD.n1763 VDD.n1194 146.341
R12735 VDD.n1773 VDD.n1194 146.341
R12736 VDD.n1773 VDD.n1190 146.341
R12737 VDD.n1779 VDD.n1190 146.341
R12738 VDD.n1779 VDD.n1182 146.341
R12739 VDD.n1789 VDD.n1182 146.341
R12740 VDD.n1789 VDD.n1178 146.341
R12741 VDD.n1795 VDD.n1178 146.341
R12742 VDD.n1795 VDD.n1170 146.341
R12743 VDD.n1805 VDD.n1170 146.341
R12744 VDD.n1805 VDD.n1166 146.341
R12745 VDD.n1811 VDD.n1166 146.341
R12746 VDD.n1811 VDD.n1157 146.341
R12747 VDD.n1821 VDD.n1157 146.341
R12748 VDD.n1821 VDD.n1153 146.341
R12749 VDD.n1827 VDD.n1153 146.341
R12750 VDD.n1827 VDD.n1146 146.341
R12751 VDD.n1837 VDD.n1146 146.341
R12752 VDD.n1837 VDD.n1142 146.341
R12753 VDD.n1843 VDD.n1142 146.341
R12754 VDD.n1843 VDD.n1134 146.341
R12755 VDD.n1853 VDD.n1134 146.341
R12756 VDD.n1853 VDD.n1130 146.341
R12757 VDD.n1859 VDD.n1130 146.341
R12758 VDD.n1859 VDD.n1122 146.341
R12759 VDD.n1869 VDD.n1122 146.341
R12760 VDD.n1869 VDD.n1118 146.341
R12761 VDD.n1875 VDD.n1118 146.341
R12762 VDD.n1875 VDD.n1110 146.341
R12763 VDD.n1885 VDD.n1110 146.341
R12764 VDD.n1885 VDD.n1106 146.341
R12765 VDD.n1891 VDD.n1106 146.341
R12766 VDD.n1891 VDD.n1095 146.341
R12767 VDD.n2213 VDD.n1095 146.341
R12768 VDD.n1338 VDD.n1337 146.341
R12769 VDD.n1342 VDD.n1337 146.341
R12770 VDD.n1344 VDD.n1343 146.341
R12771 VDD.n1463 VDD.n1462 146.341
R12772 VDD.n1348 VDD.n1347 146.341
R12773 VDD.n1352 VDD.n1351 146.341
R12774 VDD.n1354 VDD.n1353 146.341
R12775 VDD.n1358 VDD.n1357 146.341
R12776 VDD.n1446 VDD.n1445 146.341
R12777 VDD.n1362 VDD.n1361 146.341
R12778 VDD.n1364 VDD.n1363 146.341
R12779 VDD.n1368 VDD.n1367 146.341
R12780 VDD.n1370 VDD.n1369 146.341
R12781 VDD.n1376 VDD.n1375 146.341
R12782 VDD.n1378 VDD.n1377 146.341
R12783 VDD.n1382 VDD.n1381 146.341
R12784 VDD.n1384 VDD.n1383 146.341
R12785 VDD.n1413 VDD.n1387 146.341
R12786 VDD.n1389 VDD.n1388 146.341
R12787 VDD.n1393 VDD.n1392 146.341
R12788 VDD.n1395 VDD.n1394 146.341
R12789 VDD.n1399 VDD.n1398 146.341
R12790 VDD.n1481 VDD.n1315 146.341
R12791 VDD.n1489 VDD.n1307 146.341
R12792 VDD.n1489 VDD.n1303 146.341
R12793 VDD.n1495 VDD.n1303 146.341
R12794 VDD.n1495 VDD.n1295 146.341
R12795 VDD.n1505 VDD.n1295 146.341
R12796 VDD.n1505 VDD.n1291 146.341
R12797 VDD.n1511 VDD.n1291 146.341
R12798 VDD.n1511 VDD.n1283 146.341
R12799 VDD.n1521 VDD.n1283 146.341
R12800 VDD.n1521 VDD.n1279 146.341
R12801 VDD.n1527 VDD.n1279 146.341
R12802 VDD.n1527 VDD.n1271 146.341
R12803 VDD.n1537 VDD.n1271 146.341
R12804 VDD.n1537 VDD.n1267 146.341
R12805 VDD.n1543 VDD.n1267 146.341
R12806 VDD.n1543 VDD.n1259 146.341
R12807 VDD.n1554 VDD.n1259 146.341
R12808 VDD.n1554 VDD.n1255 146.341
R12809 VDD.n1560 VDD.n1255 146.341
R12810 VDD.n1560 VDD.n1248 146.341
R12811 VDD.n1570 VDD.n1248 146.341
R12812 VDD.n1570 VDD.n1244 146.341
R12813 VDD.n1576 VDD.n1244 146.341
R12814 VDD.n1576 VDD.n1236 146.341
R12815 VDD.n1586 VDD.n1236 146.341
R12816 VDD.n1586 VDD.n1232 146.341
R12817 VDD.n1592 VDD.n1232 146.341
R12818 VDD.n1592 VDD.n1224 146.341
R12819 VDD.n1602 VDD.n1224 146.341
R12820 VDD.n1602 VDD.n1220 146.341
R12821 VDD.n1608 VDD.n1220 146.341
R12822 VDD.n1608 VDD.n1212 146.341
R12823 VDD.n1618 VDD.n1212 146.341
R12824 VDD.n1618 VDD.n1208 146.341
R12825 VDD.n1755 VDD.n1208 146.341
R12826 VDD.n1755 VDD.n1200 146.341
R12827 VDD.n1765 VDD.n1200 146.341
R12828 VDD.n1765 VDD.n1196 146.341
R12829 VDD.n1771 VDD.n1196 146.341
R12830 VDD.n1771 VDD.n1188 146.341
R12831 VDD.n1781 VDD.n1188 146.341
R12832 VDD.n1781 VDD.n1184 146.341
R12833 VDD.n1787 VDD.n1184 146.341
R12834 VDD.n1787 VDD.n1176 146.341
R12835 VDD.n1797 VDD.n1176 146.341
R12836 VDD.n1797 VDD.n1172 146.341
R12837 VDD.n1803 VDD.n1172 146.341
R12838 VDD.n1803 VDD.n1164 146.341
R12839 VDD.n1813 VDD.n1164 146.341
R12840 VDD.n1813 VDD.n1160 146.341
R12841 VDD.n1819 VDD.n1160 146.341
R12842 VDD.n1819 VDD.n1152 146.341
R12843 VDD.n1829 VDD.n1152 146.341
R12844 VDD.n1829 VDD.n1148 146.341
R12845 VDD.n1835 VDD.n1148 146.341
R12846 VDD.n1835 VDD.n1140 146.341
R12847 VDD.n1845 VDD.n1140 146.341
R12848 VDD.n1845 VDD.n1136 146.341
R12849 VDD.n1851 VDD.n1136 146.341
R12850 VDD.n1851 VDD.n1128 146.341
R12851 VDD.n1861 VDD.n1128 146.341
R12852 VDD.n1861 VDD.n1124 146.341
R12853 VDD.n1867 VDD.n1124 146.341
R12854 VDD.n1867 VDD.n1116 146.341
R12855 VDD.n1877 VDD.n1116 146.341
R12856 VDD.n1877 VDD.n1112 146.341
R12857 VDD.n1883 VDD.n1112 146.341
R12858 VDD.n1883 VDD.n1104 146.341
R12859 VDD.n1893 VDD.n1104 146.341
R12860 VDD.n1893 VDD.n1099 146.341
R12861 VDD.n2211 VDD.n1099 146.341
R12862 VDD.n131 VDD.n130 136.012
R12863 VDD.n105 VDD.n104 136.012
R12864 VDD.n79 VDD.n78 136.012
R12865 VDD.n53 VDD.n52 136.012
R12866 VDD.n28 VDD.n27 136.012
R12867 VDD.n1737 VDD.n1736 136.012
R12868 VDD.n1711 VDD.n1710 136.012
R12869 VDD.n1685 VDD.n1684 136.012
R12870 VDD.n1659 VDD.n1658 136.012
R12871 VDD.n1634 VDD.n1633 136.012
R12872 VDD.n2744 VDD.n2743 126.32
R12873 VDD.n1084 VDD.t117 120.981
R12874 VDD.n802 VDD.t73 120.981
R12875 VDD.n2054 VDD.t82 120.981
R12876 VDD.n812 VDD.t64 120.981
R12877 VDD.n2759 VDD.t89 120.981
R12878 VDD.n502 VDD.t124 120.981
R12879 VDD.n2827 VDD.t92 120.981
R12880 VDD.n538 VDD.t115 120.981
R12881 VDD.n1313 VDD.n1312 107.636
R12882 VDD.n1415 VDD.n1414 107.636
R12883 VDD.n1372 VDD.n1371 107.636
R12884 VDD.n1448 VDD.n1447 107.636
R12885 VDD.n1465 VDD.n1464 107.636
R12886 VDD.n2219 VDD.n2218 107.636
R12887 VDD.n1955 VDD.n1954 107.636
R12888 VDD.n1994 VDD.n1993 107.636
R12889 VDD.n1918 VDD.n1917 107.636
R12890 VDD.n2030 VDD.n2029 107.636
R12891 VDD.n3791 VDD.n3790 107.636
R12892 VDD.n309 VDD.n308 107.636
R12893 VDD.n3827 VDD.n3826 107.636
R12894 VDD.n276 VDD.n275 107.636
R12895 VDD.n260 VDD.n259 107.636
R12896 VDD.n483 VDD.n482 107.636
R12897 VDD.n3522 VDD.n3521 107.636
R12898 VDD.n3551 VDD.n3550 107.636
R12899 VDD.n3456 VDD.n3455 107.636
R12900 VDD.n452 VDD.n451 107.636
R12901 VDD.n9 VDD.n7 107.061
R12902 VDD.n2 VDD.n0 107.061
R12903 VDD.n9 VDD.n8 103.931
R12904 VDD.n11 VDD.n10 103.931
R12905 VDD.n13 VDD.n12 103.931
R12906 VDD.n6 VDD.n5 103.931
R12907 VDD.n4 VDD.n3 103.931
R12908 VDD.n2 VDD.n1 103.931
R12909 VDD.n3101 VDD.n772 99.5127
R12910 VDD.n3105 VDD.n772 99.5127
R12911 VDD.n3105 VDD.n762 99.5127
R12912 VDD.n3113 VDD.n762 99.5127
R12913 VDD.n3113 VDD.n760 99.5127
R12914 VDD.n3117 VDD.n760 99.5127
R12915 VDD.n3117 VDD.n750 99.5127
R12916 VDD.n3125 VDD.n750 99.5127
R12917 VDD.n3125 VDD.n748 99.5127
R12918 VDD.n3129 VDD.n748 99.5127
R12919 VDD.n3129 VDD.n738 99.5127
R12920 VDD.n3137 VDD.n738 99.5127
R12921 VDD.n3137 VDD.n736 99.5127
R12922 VDD.n3141 VDD.n736 99.5127
R12923 VDD.n3141 VDD.n726 99.5127
R12924 VDD.n3149 VDD.n726 99.5127
R12925 VDD.n3149 VDD.n724 99.5127
R12926 VDD.n3153 VDD.n724 99.5127
R12927 VDD.n3153 VDD.n714 99.5127
R12928 VDD.n3161 VDD.n714 99.5127
R12929 VDD.n3161 VDD.n712 99.5127
R12930 VDD.n3165 VDD.n712 99.5127
R12931 VDD.n3165 VDD.n701 99.5127
R12932 VDD.n3173 VDD.n701 99.5127
R12933 VDD.n3173 VDD.n699 99.5127
R12934 VDD.n3177 VDD.n699 99.5127
R12935 VDD.n3177 VDD.n690 99.5127
R12936 VDD.n3185 VDD.n690 99.5127
R12937 VDD.n3185 VDD.n688 99.5127
R12938 VDD.n3189 VDD.n688 99.5127
R12939 VDD.n3189 VDD.n678 99.5127
R12940 VDD.n3197 VDD.n678 99.5127
R12941 VDD.n3197 VDD.n676 99.5127
R12942 VDD.n3201 VDD.n676 99.5127
R12943 VDD.n3201 VDD.n666 99.5127
R12944 VDD.n3209 VDD.n666 99.5127
R12945 VDD.n3209 VDD.n664 99.5127
R12946 VDD.n3213 VDD.n664 99.5127
R12947 VDD.n3213 VDD.n653 99.5127
R12948 VDD.n3221 VDD.n653 99.5127
R12949 VDD.n3221 VDD.n651 99.5127
R12950 VDD.n3225 VDD.n651 99.5127
R12951 VDD.n3225 VDD.n642 99.5127
R12952 VDD.n3233 VDD.n642 99.5127
R12953 VDD.n3233 VDD.n640 99.5127
R12954 VDD.n3237 VDD.n640 99.5127
R12955 VDD.n3237 VDD.n630 99.5127
R12956 VDD.n3245 VDD.n630 99.5127
R12957 VDD.n3245 VDD.n628 99.5127
R12958 VDD.n3249 VDD.n628 99.5127
R12959 VDD.n3249 VDD.n618 99.5127
R12960 VDD.n3257 VDD.n618 99.5127
R12961 VDD.n3257 VDD.n616 99.5127
R12962 VDD.n3261 VDD.n616 99.5127
R12963 VDD.n3261 VDD.n606 99.5127
R12964 VDD.n3269 VDD.n606 99.5127
R12965 VDD.n3269 VDD.n604 99.5127
R12966 VDD.n3273 VDD.n604 99.5127
R12967 VDD.n3273 VDD.n594 99.5127
R12968 VDD.n3281 VDD.n594 99.5127
R12969 VDD.n3281 VDD.n592 99.5127
R12970 VDD.n3285 VDD.n592 99.5127
R12971 VDD.n3285 VDD.n583 99.5127
R12972 VDD.n3293 VDD.n583 99.5127
R12973 VDD.n3293 VDD.n581 99.5127
R12974 VDD.n3297 VDD.n581 99.5127
R12975 VDD.n3297 VDD.n571 99.5127
R12976 VDD.n3305 VDD.n571 99.5127
R12977 VDD.n3305 VDD.n569 99.5127
R12978 VDD.n3309 VDD.n569 99.5127
R12979 VDD.n3309 VDD.n558 99.5127
R12980 VDD.n3317 VDD.n558 99.5127
R12981 VDD.n3317 VDD.n556 99.5127
R12982 VDD.n3321 VDD.n556 99.5127
R12983 VDD.n3321 VDD.n546 99.5127
R12984 VDD.n3331 VDD.n546 99.5127
R12985 VDD.n3331 VDD.n544 99.5127
R12986 VDD.n3335 VDD.n544 99.5127
R12987 VDD.n3335 VDD.n516 99.5127
R12988 VDD.n3395 VDD.n516 99.5127
R12989 VDD.n3395 VDD.n513 99.5127
R12990 VDD.n3426 VDD.n513 99.5127
R12991 VDD.n3426 VDD.n514 99.5127
R12992 VDD.n3420 VDD.n3419 99.5127
R12993 VDD.n3417 VDD.n3400 99.5127
R12994 VDD.n3413 VDD.n3412 99.5127
R12995 VDD.n3410 VDD.n3403 99.5127
R12996 VDD.n3406 VDD.n3405 99.5127
R12997 VDD.n3449 VDD.n3448 99.5127
R12998 VDD.n3446 VDD.n497 99.5127
R12999 VDD.n3442 VDD.n3441 99.5127
R13000 VDD.n3439 VDD.n500 99.5127
R13001 VDD.n3435 VDD.n3434 99.5127
R13002 VDD.n2836 VDD.n2745 99.5127
R13003 VDD.n2836 VDD.n770 99.5127
R13004 VDD.n2839 VDD.n770 99.5127
R13005 VDD.n2839 VDD.n764 99.5127
R13006 VDD.n2842 VDD.n764 99.5127
R13007 VDD.n2842 VDD.n758 99.5127
R13008 VDD.n2845 VDD.n758 99.5127
R13009 VDD.n2845 VDD.n752 99.5127
R13010 VDD.n2848 VDD.n752 99.5127
R13011 VDD.n2848 VDD.n746 99.5127
R13012 VDD.n2851 VDD.n746 99.5127
R13013 VDD.n2851 VDD.n740 99.5127
R13014 VDD.n2854 VDD.n740 99.5127
R13015 VDD.n2854 VDD.n734 99.5127
R13016 VDD.n2857 VDD.n734 99.5127
R13017 VDD.n2857 VDD.n728 99.5127
R13018 VDD.n2860 VDD.n728 99.5127
R13019 VDD.n2860 VDD.n722 99.5127
R13020 VDD.n2863 VDD.n722 99.5127
R13021 VDD.n2863 VDD.n716 99.5127
R13022 VDD.n2866 VDD.n716 99.5127
R13023 VDD.n2866 VDD.n710 99.5127
R13024 VDD.n2869 VDD.n710 99.5127
R13025 VDD.n2869 VDD.n703 99.5127
R13026 VDD.n2872 VDD.n703 99.5127
R13027 VDD.n2872 VDD.n697 99.5127
R13028 VDD.n2875 VDD.n697 99.5127
R13029 VDD.n2875 VDD.n692 99.5127
R13030 VDD.n2878 VDD.n692 99.5127
R13031 VDD.n2878 VDD.n686 99.5127
R13032 VDD.n2881 VDD.n686 99.5127
R13033 VDD.n2881 VDD.n680 99.5127
R13034 VDD.n2884 VDD.n680 99.5127
R13035 VDD.n2884 VDD.n674 99.5127
R13036 VDD.n2887 VDD.n674 99.5127
R13037 VDD.n2887 VDD.n668 99.5127
R13038 VDD.n2890 VDD.n668 99.5127
R13039 VDD.n2890 VDD.n662 99.5127
R13040 VDD.n2893 VDD.n662 99.5127
R13041 VDD.n2893 VDD.n655 99.5127
R13042 VDD.n2896 VDD.n655 99.5127
R13043 VDD.n2896 VDD.n649 99.5127
R13044 VDD.n2899 VDD.n649 99.5127
R13045 VDD.n2899 VDD.n644 99.5127
R13046 VDD.n2902 VDD.n644 99.5127
R13047 VDD.n2902 VDD.n638 99.5127
R13048 VDD.n2905 VDD.n638 99.5127
R13049 VDD.n2905 VDD.n632 99.5127
R13050 VDD.n2908 VDD.n632 99.5127
R13051 VDD.n2908 VDD.n626 99.5127
R13052 VDD.n2911 VDD.n626 99.5127
R13053 VDD.n2911 VDD.n620 99.5127
R13054 VDD.n2914 VDD.n620 99.5127
R13055 VDD.n2914 VDD.n614 99.5127
R13056 VDD.n2917 VDD.n614 99.5127
R13057 VDD.n2917 VDD.n608 99.5127
R13058 VDD.n2920 VDD.n608 99.5127
R13059 VDD.n2920 VDD.n602 99.5127
R13060 VDD.n2923 VDD.n602 99.5127
R13061 VDD.n2923 VDD.n596 99.5127
R13062 VDD.n2926 VDD.n596 99.5127
R13063 VDD.n2926 VDD.n590 99.5127
R13064 VDD.n2955 VDD.n590 99.5127
R13065 VDD.n2955 VDD.n584 99.5127
R13066 VDD.n2951 VDD.n584 99.5127
R13067 VDD.n2951 VDD.n579 99.5127
R13068 VDD.n2948 VDD.n579 99.5127
R13069 VDD.n2948 VDD.n573 99.5127
R13070 VDD.n2945 VDD.n573 99.5127
R13071 VDD.n2945 VDD.n567 99.5127
R13072 VDD.n2942 VDD.n567 99.5127
R13073 VDD.n2942 VDD.n560 99.5127
R13074 VDD.n2939 VDD.n560 99.5127
R13075 VDD.n2939 VDD.n554 99.5127
R13076 VDD.n2936 VDD.n554 99.5127
R13077 VDD.n2936 VDD.n548 99.5127
R13078 VDD.n2933 VDD.n548 99.5127
R13079 VDD.n2933 VDD.n542 99.5127
R13080 VDD.n2930 VDD.n542 99.5127
R13081 VDD.n2930 VDD.n518 99.5127
R13082 VDD.n518 VDD.n508 99.5127
R13083 VDD.n3428 VDD.n508 99.5127
R13084 VDD.n3428 VDD.n506 99.5127
R13085 VDD.n2791 VDD.n2789 99.5127
R13086 VDD.n2795 VDD.n2789 99.5127
R13087 VDD.n2799 VDD.n2797 99.5127
R13088 VDD.n2803 VDD.n2787 99.5127
R13089 VDD.n2807 VDD.n2805 99.5127
R13090 VDD.n2811 VDD.n2785 99.5127
R13091 VDD.n2815 VDD.n2813 99.5127
R13092 VDD.n2819 VDD.n2783 99.5127
R13093 VDD.n2823 VDD.n2821 99.5127
R13094 VDD.n2830 VDD.n2781 99.5127
R13095 VDD.n2833 VDD.n2832 99.5127
R13096 VDD.n2689 VDD.n2688 99.5127
R13097 VDD.n2685 VDD.n2684 99.5127
R13098 VDD.n2681 VDD.n2680 99.5127
R13099 VDD.n2677 VDD.n2676 99.5127
R13100 VDD.n2673 VDD.n2672 99.5127
R13101 VDD.n2669 VDD.n2668 99.5127
R13102 VDD.n2665 VDD.n2664 99.5127
R13103 VDD.n2661 VDD.n2660 99.5127
R13104 VDD.n2657 VDD.n2656 99.5127
R13105 VDD.n2653 VDD.n2652 99.5127
R13106 VDD.n2171 VDD.n1057 99.5127
R13107 VDD.n2171 VDD.n1052 99.5127
R13108 VDD.n2168 VDD.n1052 99.5127
R13109 VDD.n2168 VDD.n1046 99.5127
R13110 VDD.n2165 VDD.n1046 99.5127
R13111 VDD.n2165 VDD.n1040 99.5127
R13112 VDD.n2162 VDD.n1040 99.5127
R13113 VDD.n2162 VDD.n1033 99.5127
R13114 VDD.n2159 VDD.n1033 99.5127
R13115 VDD.n2159 VDD.n1027 99.5127
R13116 VDD.n2156 VDD.n1027 99.5127
R13117 VDD.n2156 VDD.n1022 99.5127
R13118 VDD.n2153 VDD.n1022 99.5127
R13119 VDD.n2153 VDD.n1016 99.5127
R13120 VDD.n2150 VDD.n1016 99.5127
R13121 VDD.n2150 VDD.n1010 99.5127
R13122 VDD.n2147 VDD.n1010 99.5127
R13123 VDD.n2147 VDD.n1003 99.5127
R13124 VDD.n2144 VDD.n1003 99.5127
R13125 VDD.n2144 VDD.n997 99.5127
R13126 VDD.n2141 VDD.n997 99.5127
R13127 VDD.n2141 VDD.n992 99.5127
R13128 VDD.n2138 VDD.n992 99.5127
R13129 VDD.n2138 VDD.n986 99.5127
R13130 VDD.n2135 VDD.n986 99.5127
R13131 VDD.n2135 VDD.n980 99.5127
R13132 VDD.n2132 VDD.n980 99.5127
R13133 VDD.n2132 VDD.n974 99.5127
R13134 VDD.n2129 VDD.n974 99.5127
R13135 VDD.n2129 VDD.n968 99.5127
R13136 VDD.n2126 VDD.n968 99.5127
R13137 VDD.n2126 VDD.n962 99.5127
R13138 VDD.n2123 VDD.n962 99.5127
R13139 VDD.n2123 VDD.n956 99.5127
R13140 VDD.n2120 VDD.n956 99.5127
R13141 VDD.n2120 VDD.n950 99.5127
R13142 VDD.n2117 VDD.n950 99.5127
R13143 VDD.n2117 VDD.n944 99.5127
R13144 VDD.n2114 VDD.n944 99.5127
R13145 VDD.n2114 VDD.n937 99.5127
R13146 VDD.n2111 VDD.n937 99.5127
R13147 VDD.n2111 VDD.n931 99.5127
R13148 VDD.n2108 VDD.n931 99.5127
R13149 VDD.n2108 VDD.n926 99.5127
R13150 VDD.n2105 VDD.n926 99.5127
R13151 VDD.n2105 VDD.n920 99.5127
R13152 VDD.n2102 VDD.n920 99.5127
R13153 VDD.n2102 VDD.n914 99.5127
R13154 VDD.n2099 VDD.n914 99.5127
R13155 VDD.n2099 VDD.n908 99.5127
R13156 VDD.n2096 VDD.n908 99.5127
R13157 VDD.n2096 VDD.n902 99.5127
R13158 VDD.n2093 VDD.n902 99.5127
R13159 VDD.n2093 VDD.n896 99.5127
R13160 VDD.n2090 VDD.n896 99.5127
R13161 VDD.n2090 VDD.n889 99.5127
R13162 VDD.n2087 VDD.n889 99.5127
R13163 VDD.n2087 VDD.n883 99.5127
R13164 VDD.n2084 VDD.n883 99.5127
R13165 VDD.n2084 VDD.n878 99.5127
R13166 VDD.n2081 VDD.n878 99.5127
R13167 VDD.n2081 VDD.n872 99.5127
R13168 VDD.n2078 VDD.n872 99.5127
R13169 VDD.n2078 VDD.n866 99.5127
R13170 VDD.n2075 VDD.n866 99.5127
R13171 VDD.n2075 VDD.n860 99.5127
R13172 VDD.n2072 VDD.n860 99.5127
R13173 VDD.n2072 VDD.n854 99.5127
R13174 VDD.n2069 VDD.n854 99.5127
R13175 VDD.n2069 VDD.n848 99.5127
R13176 VDD.n2066 VDD.n848 99.5127
R13177 VDD.n2066 VDD.n842 99.5127
R13178 VDD.n2063 VDD.n842 99.5127
R13179 VDD.n2063 VDD.n836 99.5127
R13180 VDD.n2060 VDD.n836 99.5127
R13181 VDD.n2060 VDD.n830 99.5127
R13182 VDD.n2057 VDD.n830 99.5127
R13183 VDD.n2057 VDD.n823 99.5127
R13184 VDD.n823 VDD.n815 99.5127
R13185 VDD.n2643 VDD.n815 99.5127
R13186 VDD.n2644 VDD.n2643 99.5127
R13187 VDD.n2644 VDD.n806 99.5127
R13188 VDD.n2648 VDD.n806 99.5127
R13189 VDD.n2392 VDD.n1061 99.5127
R13190 VDD.n2038 VDD.n1061 99.5127
R13191 VDD.n2042 VDD.n2041 99.5127
R13192 VDD.n2046 VDD.n2045 99.5127
R13193 VDD.n2050 VDD.n2049 99.5127
R13194 VDD.n2195 VDD.n2194 99.5127
R13195 VDD.n2192 VDD.n2191 99.5127
R13196 VDD.n2188 VDD.n2187 99.5127
R13197 VDD.n2184 VDD.n2183 99.5127
R13198 VDD.n2180 VDD.n2179 99.5127
R13199 VDD.n2175 VDD.n1071 99.5127
R13200 VDD.n2396 VDD.n1050 99.5127
R13201 VDD.n2404 VDD.n1050 99.5127
R13202 VDD.n2404 VDD.n1048 99.5127
R13203 VDD.n2408 VDD.n1048 99.5127
R13204 VDD.n2408 VDD.n1038 99.5127
R13205 VDD.n2416 VDD.n1038 99.5127
R13206 VDD.n2416 VDD.n1036 99.5127
R13207 VDD.n2420 VDD.n1036 99.5127
R13208 VDD.n2420 VDD.n1026 99.5127
R13209 VDD.n2428 VDD.n1026 99.5127
R13210 VDD.n2428 VDD.n1024 99.5127
R13211 VDD.n2432 VDD.n1024 99.5127
R13212 VDD.n2432 VDD.n1014 99.5127
R13213 VDD.n2440 VDD.n1014 99.5127
R13214 VDD.n2440 VDD.n1012 99.5127
R13215 VDD.n2444 VDD.n1012 99.5127
R13216 VDD.n2444 VDD.n1001 99.5127
R13217 VDD.n2452 VDD.n1001 99.5127
R13218 VDD.n2452 VDD.n999 99.5127
R13219 VDD.n2456 VDD.n999 99.5127
R13220 VDD.n2456 VDD.n990 99.5127
R13221 VDD.n2464 VDD.n990 99.5127
R13222 VDD.n2464 VDD.n988 99.5127
R13223 VDD.n2468 VDD.n988 99.5127
R13224 VDD.n2468 VDD.n978 99.5127
R13225 VDD.n2476 VDD.n978 99.5127
R13226 VDD.n2476 VDD.n976 99.5127
R13227 VDD.n2480 VDD.n976 99.5127
R13228 VDD.n2480 VDD.n966 99.5127
R13229 VDD.n2488 VDD.n966 99.5127
R13230 VDD.n2488 VDD.n964 99.5127
R13231 VDD.n2492 VDD.n964 99.5127
R13232 VDD.n2492 VDD.n954 99.5127
R13233 VDD.n2500 VDD.n954 99.5127
R13234 VDD.n2500 VDD.n952 99.5127
R13235 VDD.n2504 VDD.n952 99.5127
R13236 VDD.n2504 VDD.n942 99.5127
R13237 VDD.n2512 VDD.n942 99.5127
R13238 VDD.n2512 VDD.n940 99.5127
R13239 VDD.n2516 VDD.n940 99.5127
R13240 VDD.n2516 VDD.n930 99.5127
R13241 VDD.n2524 VDD.n930 99.5127
R13242 VDD.n2524 VDD.n928 99.5127
R13243 VDD.n2528 VDD.n928 99.5127
R13244 VDD.n2528 VDD.n918 99.5127
R13245 VDD.n2536 VDD.n918 99.5127
R13246 VDD.n2536 VDD.n916 99.5127
R13247 VDD.n2540 VDD.n916 99.5127
R13248 VDD.n2540 VDD.n906 99.5127
R13249 VDD.n2548 VDD.n906 99.5127
R13250 VDD.n2548 VDD.n904 99.5127
R13251 VDD.n2552 VDD.n904 99.5127
R13252 VDD.n2552 VDD.n894 99.5127
R13253 VDD.n2560 VDD.n894 99.5127
R13254 VDD.n2560 VDD.n892 99.5127
R13255 VDD.n2564 VDD.n892 99.5127
R13256 VDD.n2564 VDD.n882 99.5127
R13257 VDD.n2572 VDD.n882 99.5127
R13258 VDD.n2572 VDD.n880 99.5127
R13259 VDD.n2576 VDD.n880 99.5127
R13260 VDD.n2576 VDD.n870 99.5127
R13261 VDD.n2584 VDD.n870 99.5127
R13262 VDD.n2584 VDD.n868 99.5127
R13263 VDD.n2588 VDD.n868 99.5127
R13264 VDD.n2588 VDD.n858 99.5127
R13265 VDD.n2596 VDD.n858 99.5127
R13266 VDD.n2596 VDD.n856 99.5127
R13267 VDD.n2600 VDD.n856 99.5127
R13268 VDD.n2600 VDD.n846 99.5127
R13269 VDD.n2608 VDD.n846 99.5127
R13270 VDD.n2608 VDD.n844 99.5127
R13271 VDD.n2612 VDD.n844 99.5127
R13272 VDD.n2612 VDD.n834 99.5127
R13273 VDD.n2620 VDD.n834 99.5127
R13274 VDD.n2620 VDD.n832 99.5127
R13275 VDD.n2624 VDD.n832 99.5127
R13276 VDD.n2624 VDD.n821 99.5127
R13277 VDD.n2637 VDD.n821 99.5127
R13278 VDD.n2637 VDD.n819 99.5127
R13279 VDD.n2641 VDD.n819 99.5127
R13280 VDD.n2641 VDD.n808 99.5127
R13281 VDD.n2695 VDD.n808 99.5127
R13282 VDD.n2695 VDD.n809 99.5127
R13283 VDD.n3385 VDD.n524 99.5127
R13284 VDD.n3381 VDD.n3380 99.5127
R13285 VDD.n3378 VDD.n527 99.5127
R13286 VDD.n3374 VDD.n3373 99.5127
R13287 VDD.n3371 VDD.n3368 99.5127
R13288 VDD.n3366 VDD.n530 99.5127
R13289 VDD.n3362 VDD.n3361 99.5127
R13290 VDD.n3359 VDD.n533 99.5127
R13291 VDD.n3355 VDD.n3354 99.5127
R13292 VDD.n3352 VDD.n536 99.5127
R13293 VDD.n3050 VDD.n2746 99.5127
R13294 VDD.n3050 VDD.n771 99.5127
R13295 VDD.n3047 VDD.n771 99.5127
R13296 VDD.n3047 VDD.n765 99.5127
R13297 VDD.n3044 VDD.n765 99.5127
R13298 VDD.n3044 VDD.n759 99.5127
R13299 VDD.n3041 VDD.n759 99.5127
R13300 VDD.n3041 VDD.n753 99.5127
R13301 VDD.n3038 VDD.n753 99.5127
R13302 VDD.n3038 VDD.n747 99.5127
R13303 VDD.n3035 VDD.n747 99.5127
R13304 VDD.n3035 VDD.n741 99.5127
R13305 VDD.n3032 VDD.n741 99.5127
R13306 VDD.n3032 VDD.n735 99.5127
R13307 VDD.n3029 VDD.n735 99.5127
R13308 VDD.n3029 VDD.n729 99.5127
R13309 VDD.n3026 VDD.n729 99.5127
R13310 VDD.n3026 VDD.n723 99.5127
R13311 VDD.n3023 VDD.n723 99.5127
R13312 VDD.n3023 VDD.n717 99.5127
R13313 VDD.n3020 VDD.n717 99.5127
R13314 VDD.n3020 VDD.n711 99.5127
R13315 VDD.n3017 VDD.n711 99.5127
R13316 VDD.n3017 VDD.n704 99.5127
R13317 VDD.n3014 VDD.n704 99.5127
R13318 VDD.n3014 VDD.n698 99.5127
R13319 VDD.n3011 VDD.n698 99.5127
R13320 VDD.n3011 VDD.n693 99.5127
R13321 VDD.n3008 VDD.n693 99.5127
R13322 VDD.n3008 VDD.n687 99.5127
R13323 VDD.n3005 VDD.n687 99.5127
R13324 VDD.n3005 VDD.n681 99.5127
R13325 VDD.n3002 VDD.n681 99.5127
R13326 VDD.n3002 VDD.n675 99.5127
R13327 VDD.n2999 VDD.n675 99.5127
R13328 VDD.n2999 VDD.n669 99.5127
R13329 VDD.n2996 VDD.n669 99.5127
R13330 VDD.n2996 VDD.n663 99.5127
R13331 VDD.n2993 VDD.n663 99.5127
R13332 VDD.n2993 VDD.n656 99.5127
R13333 VDD.n2990 VDD.n656 99.5127
R13334 VDD.n2990 VDD.n650 99.5127
R13335 VDD.n2987 VDD.n650 99.5127
R13336 VDD.n2987 VDD.n645 99.5127
R13337 VDD.n2984 VDD.n645 99.5127
R13338 VDD.n2984 VDD.n639 99.5127
R13339 VDD.n2981 VDD.n639 99.5127
R13340 VDD.n2981 VDD.n633 99.5127
R13341 VDD.n2978 VDD.n633 99.5127
R13342 VDD.n2978 VDD.n627 99.5127
R13343 VDD.n2975 VDD.n627 99.5127
R13344 VDD.n2975 VDD.n621 99.5127
R13345 VDD.n2972 VDD.n621 99.5127
R13346 VDD.n2972 VDD.n615 99.5127
R13347 VDD.n2969 VDD.n615 99.5127
R13348 VDD.n2969 VDD.n609 99.5127
R13349 VDD.n2966 VDD.n609 99.5127
R13350 VDD.n2966 VDD.n603 99.5127
R13351 VDD.n2963 VDD.n603 99.5127
R13352 VDD.n2963 VDD.n597 99.5127
R13353 VDD.n2960 VDD.n597 99.5127
R13354 VDD.n2960 VDD.n591 99.5127
R13355 VDD.n2957 VDD.n591 99.5127
R13356 VDD.n2957 VDD.n585 99.5127
R13357 VDD.n2777 VDD.n585 99.5127
R13358 VDD.n2777 VDD.n580 99.5127
R13359 VDD.n2774 VDD.n580 99.5127
R13360 VDD.n2774 VDD.n574 99.5127
R13361 VDD.n2771 VDD.n574 99.5127
R13362 VDD.n2771 VDD.n568 99.5127
R13363 VDD.n2768 VDD.n568 99.5127
R13364 VDD.n2768 VDD.n561 99.5127
R13365 VDD.n2765 VDD.n561 99.5127
R13366 VDD.n2765 VDD.n555 99.5127
R13367 VDD.n2762 VDD.n555 99.5127
R13368 VDD.n2762 VDD.n549 99.5127
R13369 VDD.n549 VDD.n540 99.5127
R13370 VDD.n3337 VDD.n540 99.5127
R13371 VDD.n3338 VDD.n3337 99.5127
R13372 VDD.n3338 VDD.n519 99.5127
R13373 VDD.n3341 VDD.n519 99.5127
R13374 VDD.n3341 VDD.n510 99.5127
R13375 VDD.n3346 VDD.n510 99.5127
R13376 VDD.n3095 VDD.n3093 99.5127
R13377 VDD.n3091 VDD.n2749 99.5127
R13378 VDD.n3087 VDD.n3085 99.5127
R13379 VDD.n3083 VDD.n2751 99.5127
R13380 VDD.n3079 VDD.n3077 99.5127
R13381 VDD.n3075 VDD.n2753 99.5127
R13382 VDD.n3071 VDD.n3069 99.5127
R13383 VDD.n3067 VDD.n2755 99.5127
R13384 VDD.n3063 VDD.n3061 99.5127
R13385 VDD.n3059 VDD.n2757 99.5127
R13386 VDD.n3099 VDD.n768 99.5127
R13387 VDD.n3107 VDD.n768 99.5127
R13388 VDD.n3107 VDD.n766 99.5127
R13389 VDD.n3111 VDD.n766 99.5127
R13390 VDD.n3111 VDD.n756 99.5127
R13391 VDD.n3119 VDD.n756 99.5127
R13392 VDD.n3119 VDD.n754 99.5127
R13393 VDD.n3123 VDD.n754 99.5127
R13394 VDD.n3123 VDD.n744 99.5127
R13395 VDD.n3131 VDD.n744 99.5127
R13396 VDD.n3131 VDD.n742 99.5127
R13397 VDD.n3135 VDD.n742 99.5127
R13398 VDD.n3135 VDD.n732 99.5127
R13399 VDD.n3143 VDD.n732 99.5127
R13400 VDD.n3143 VDD.n730 99.5127
R13401 VDD.n3147 VDD.n730 99.5127
R13402 VDD.n3147 VDD.n720 99.5127
R13403 VDD.n3155 VDD.n720 99.5127
R13404 VDD.n3155 VDD.n718 99.5127
R13405 VDD.n3159 VDD.n718 99.5127
R13406 VDD.n3159 VDD.n708 99.5127
R13407 VDD.n3167 VDD.n708 99.5127
R13408 VDD.n3167 VDD.n706 99.5127
R13409 VDD.n3171 VDD.n706 99.5127
R13410 VDD.n3171 VDD.n696 99.5127
R13411 VDD.n3179 VDD.n696 99.5127
R13412 VDD.n3179 VDD.n694 99.5127
R13413 VDD.n3183 VDD.n694 99.5127
R13414 VDD.n3183 VDD.n684 99.5127
R13415 VDD.n3191 VDD.n684 99.5127
R13416 VDD.n3191 VDD.n682 99.5127
R13417 VDD.n3195 VDD.n682 99.5127
R13418 VDD.n3195 VDD.n672 99.5127
R13419 VDD.n3203 VDD.n672 99.5127
R13420 VDD.n3203 VDD.n670 99.5127
R13421 VDD.n3207 VDD.n670 99.5127
R13422 VDD.n3207 VDD.n660 99.5127
R13423 VDD.n3215 VDD.n660 99.5127
R13424 VDD.n3215 VDD.n658 99.5127
R13425 VDD.n3219 VDD.n658 99.5127
R13426 VDD.n3219 VDD.n648 99.5127
R13427 VDD.n3227 VDD.n648 99.5127
R13428 VDD.n3227 VDD.n646 99.5127
R13429 VDD.n3231 VDD.n646 99.5127
R13430 VDD.n3231 VDD.n636 99.5127
R13431 VDD.n3239 VDD.n636 99.5127
R13432 VDD.n3239 VDD.n634 99.5127
R13433 VDD.n3243 VDD.n634 99.5127
R13434 VDD.n3243 VDD.n624 99.5127
R13435 VDD.n3251 VDD.n624 99.5127
R13436 VDD.n3251 VDD.n622 99.5127
R13437 VDD.n3255 VDD.n622 99.5127
R13438 VDD.n3255 VDD.n612 99.5127
R13439 VDD.n3263 VDD.n612 99.5127
R13440 VDD.n3263 VDD.n610 99.5127
R13441 VDD.n3267 VDD.n610 99.5127
R13442 VDD.n3267 VDD.n600 99.5127
R13443 VDD.n3275 VDD.n600 99.5127
R13444 VDD.n3275 VDD.n598 99.5127
R13445 VDD.n3279 VDD.n598 99.5127
R13446 VDD.n3279 VDD.n588 99.5127
R13447 VDD.n3287 VDD.n588 99.5127
R13448 VDD.n3287 VDD.n586 99.5127
R13449 VDD.n3291 VDD.n586 99.5127
R13450 VDD.n3291 VDD.n577 99.5127
R13451 VDD.n3299 VDD.n577 99.5127
R13452 VDD.n3299 VDD.n575 99.5127
R13453 VDD.n3303 VDD.n575 99.5127
R13454 VDD.n3303 VDD.n565 99.5127
R13455 VDD.n3311 VDD.n565 99.5127
R13456 VDD.n3311 VDD.n563 99.5127
R13457 VDD.n3315 VDD.n563 99.5127
R13458 VDD.n3315 VDD.n553 99.5127
R13459 VDD.n3323 VDD.n553 99.5127
R13460 VDD.n3323 VDD.n550 99.5127
R13461 VDD.n3329 VDD.n550 99.5127
R13462 VDD.n3329 VDD.n551 99.5127
R13463 VDD.n551 VDD.n543 99.5127
R13464 VDD.n543 VDD.n520 99.5127
R13465 VDD.n3393 VDD.n520 99.5127
R13466 VDD.n3393 VDD.n521 99.5127
R13467 VDD.n521 VDD.n512 99.5127
R13468 VDD.n3388 VDD.n512 99.5127
R13469 VDD.n2742 VDD.n799 99.5127
R13470 VDD.n2738 VDD.n2737 99.5127
R13471 VDD.n2734 VDD.n2733 99.5127
R13472 VDD.n2730 VDD.n2729 99.5127
R13473 VDD.n2726 VDD.n2725 99.5127
R13474 VDD.n2722 VDD.n2721 99.5127
R13475 VDD.n2718 VDD.n2717 99.5127
R13476 VDD.n2714 VDD.n2713 99.5127
R13477 VDD.n2710 VDD.n2709 99.5127
R13478 VDD.n2706 VDD.n2705 99.5127
R13479 VDD.n2701 VDD.n797 99.5127
R13480 VDD.n2385 VDD.n1058 99.5127
R13481 VDD.n2385 VDD.n1053 99.5127
R13482 VDD.n2382 VDD.n1053 99.5127
R13483 VDD.n2382 VDD.n1047 99.5127
R13484 VDD.n2379 VDD.n1047 99.5127
R13485 VDD.n2379 VDD.n1041 99.5127
R13486 VDD.n2376 VDD.n1041 99.5127
R13487 VDD.n2376 VDD.n1034 99.5127
R13488 VDD.n2373 VDD.n1034 99.5127
R13489 VDD.n2373 VDD.n1028 99.5127
R13490 VDD.n2370 VDD.n1028 99.5127
R13491 VDD.n2370 VDD.n1023 99.5127
R13492 VDD.n2367 VDD.n1023 99.5127
R13493 VDD.n2367 VDD.n1017 99.5127
R13494 VDD.n2364 VDD.n1017 99.5127
R13495 VDD.n2364 VDD.n1011 99.5127
R13496 VDD.n2361 VDD.n1011 99.5127
R13497 VDD.n2361 VDD.n1004 99.5127
R13498 VDD.n2358 VDD.n1004 99.5127
R13499 VDD.n2358 VDD.n998 99.5127
R13500 VDD.n2355 VDD.n998 99.5127
R13501 VDD.n2355 VDD.n993 99.5127
R13502 VDD.n2352 VDD.n993 99.5127
R13503 VDD.n2352 VDD.n987 99.5127
R13504 VDD.n2349 VDD.n987 99.5127
R13505 VDD.n2349 VDD.n981 99.5127
R13506 VDD.n2346 VDD.n981 99.5127
R13507 VDD.n2346 VDD.n975 99.5127
R13508 VDD.n2343 VDD.n975 99.5127
R13509 VDD.n2343 VDD.n969 99.5127
R13510 VDD.n2340 VDD.n969 99.5127
R13511 VDD.n2340 VDD.n963 99.5127
R13512 VDD.n2337 VDD.n963 99.5127
R13513 VDD.n2337 VDD.n957 99.5127
R13514 VDD.n2334 VDD.n957 99.5127
R13515 VDD.n2334 VDD.n951 99.5127
R13516 VDD.n2331 VDD.n951 99.5127
R13517 VDD.n2331 VDD.n945 99.5127
R13518 VDD.n2328 VDD.n945 99.5127
R13519 VDD.n2328 VDD.n938 99.5127
R13520 VDD.n2325 VDD.n938 99.5127
R13521 VDD.n2325 VDD.n932 99.5127
R13522 VDD.n2322 VDD.n932 99.5127
R13523 VDD.n2322 VDD.n927 99.5127
R13524 VDD.n2319 VDD.n927 99.5127
R13525 VDD.n2319 VDD.n921 99.5127
R13526 VDD.n2316 VDD.n921 99.5127
R13527 VDD.n2316 VDD.n915 99.5127
R13528 VDD.n2313 VDD.n915 99.5127
R13529 VDD.n2313 VDD.n909 99.5127
R13530 VDD.n2310 VDD.n909 99.5127
R13531 VDD.n2310 VDD.n903 99.5127
R13532 VDD.n2307 VDD.n903 99.5127
R13533 VDD.n2307 VDD.n897 99.5127
R13534 VDD.n2304 VDD.n897 99.5127
R13535 VDD.n2304 VDD.n890 99.5127
R13536 VDD.n2301 VDD.n890 99.5127
R13537 VDD.n2301 VDD.n884 99.5127
R13538 VDD.n2298 VDD.n884 99.5127
R13539 VDD.n2298 VDD.n879 99.5127
R13540 VDD.n2295 VDD.n879 99.5127
R13541 VDD.n2295 VDD.n873 99.5127
R13542 VDD.n2292 VDD.n873 99.5127
R13543 VDD.n2292 VDD.n867 99.5127
R13544 VDD.n2289 VDD.n867 99.5127
R13545 VDD.n2289 VDD.n861 99.5127
R13546 VDD.n2286 VDD.n861 99.5127
R13547 VDD.n2286 VDD.n855 99.5127
R13548 VDD.n2283 VDD.n855 99.5127
R13549 VDD.n2283 VDD.n849 99.5127
R13550 VDD.n2280 VDD.n849 99.5127
R13551 VDD.n2280 VDD.n843 99.5127
R13552 VDD.n2277 VDD.n843 99.5127
R13553 VDD.n2277 VDD.n837 99.5127
R13554 VDD.n2274 VDD.n837 99.5127
R13555 VDD.n2274 VDD.n831 99.5127
R13556 VDD.n2271 VDD.n831 99.5127
R13557 VDD.n2271 VDD.n824 99.5127
R13558 VDD.n2268 VDD.n824 99.5127
R13559 VDD.n2268 VDD.n817 99.5127
R13560 VDD.n817 VDD.n804 99.5127
R13561 VDD.n2697 VDD.n804 99.5127
R13562 VDD.n2698 VDD.n2697 99.5127
R13563 VDD.n2226 VDD.n1056 99.5127
R13564 VDD.n2230 VDD.n2229 99.5127
R13565 VDD.n2234 VDD.n2233 99.5127
R13566 VDD.n2238 VDD.n2237 99.5127
R13567 VDD.n2242 VDD.n2241 99.5127
R13568 VDD.n2246 VDD.n2245 99.5127
R13569 VDD.n2250 VDD.n2249 99.5127
R13570 VDD.n2254 VDD.n2253 99.5127
R13571 VDD.n2258 VDD.n2257 99.5127
R13572 VDD.n2262 VDD.n2261 99.5127
R13573 VDD.n2389 VDD.n1082 99.5127
R13574 VDD.n2398 VDD.n1054 99.5127
R13575 VDD.n2402 VDD.n1054 99.5127
R13576 VDD.n2402 VDD.n1044 99.5127
R13577 VDD.n2410 VDD.n1044 99.5127
R13578 VDD.n2410 VDD.n1042 99.5127
R13579 VDD.n2414 VDD.n1042 99.5127
R13580 VDD.n2414 VDD.n1031 99.5127
R13581 VDD.n2422 VDD.n1031 99.5127
R13582 VDD.n2422 VDD.n1029 99.5127
R13583 VDD.n2426 VDD.n1029 99.5127
R13584 VDD.n2426 VDD.n1020 99.5127
R13585 VDD.n2434 VDD.n1020 99.5127
R13586 VDD.n2434 VDD.n1018 99.5127
R13587 VDD.n2438 VDD.n1018 99.5127
R13588 VDD.n2438 VDD.n1008 99.5127
R13589 VDD.n2446 VDD.n1008 99.5127
R13590 VDD.n2446 VDD.n1006 99.5127
R13591 VDD.n2450 VDD.n1006 99.5127
R13592 VDD.n2450 VDD.n996 99.5127
R13593 VDD.n2458 VDD.n996 99.5127
R13594 VDD.n2458 VDD.n994 99.5127
R13595 VDD.n2462 VDD.n994 99.5127
R13596 VDD.n2462 VDD.n984 99.5127
R13597 VDD.n2470 VDD.n984 99.5127
R13598 VDD.n2470 VDD.n982 99.5127
R13599 VDD.n2474 VDD.n982 99.5127
R13600 VDD.n2474 VDD.n972 99.5127
R13601 VDD.n2482 VDD.n972 99.5127
R13602 VDD.n2482 VDD.n970 99.5127
R13603 VDD.n2486 VDD.n970 99.5127
R13604 VDD.n2486 VDD.n960 99.5127
R13605 VDD.n2494 VDD.n960 99.5127
R13606 VDD.n2494 VDD.n958 99.5127
R13607 VDD.n2498 VDD.n958 99.5127
R13608 VDD.n2498 VDD.n948 99.5127
R13609 VDD.n2506 VDD.n948 99.5127
R13610 VDD.n2506 VDD.n946 99.5127
R13611 VDD.n2510 VDD.n946 99.5127
R13612 VDD.n2510 VDD.n935 99.5127
R13613 VDD.n2518 VDD.n935 99.5127
R13614 VDD.n2518 VDD.n933 99.5127
R13615 VDD.n2522 VDD.n933 99.5127
R13616 VDD.n2522 VDD.n924 99.5127
R13617 VDD.n2530 VDD.n924 99.5127
R13618 VDD.n2530 VDD.n922 99.5127
R13619 VDD.n2534 VDD.n922 99.5127
R13620 VDD.n2534 VDD.n912 99.5127
R13621 VDD.n2542 VDD.n912 99.5127
R13622 VDD.n2542 VDD.n910 99.5127
R13623 VDD.n2546 VDD.n910 99.5127
R13624 VDD.n2546 VDD.n900 99.5127
R13625 VDD.n2554 VDD.n900 99.5127
R13626 VDD.n2554 VDD.n898 99.5127
R13627 VDD.n2558 VDD.n898 99.5127
R13628 VDD.n2558 VDD.n887 99.5127
R13629 VDD.n2566 VDD.n887 99.5127
R13630 VDD.n2566 VDD.n885 99.5127
R13631 VDD.n2570 VDD.n885 99.5127
R13632 VDD.n2570 VDD.n876 99.5127
R13633 VDD.n2578 VDD.n876 99.5127
R13634 VDD.n2578 VDD.n874 99.5127
R13635 VDD.n2582 VDD.n874 99.5127
R13636 VDD.n2582 VDD.n864 99.5127
R13637 VDD.n2590 VDD.n864 99.5127
R13638 VDD.n2590 VDD.n862 99.5127
R13639 VDD.n2594 VDD.n862 99.5127
R13640 VDD.n2594 VDD.n852 99.5127
R13641 VDD.n2602 VDD.n852 99.5127
R13642 VDD.n2602 VDD.n850 99.5127
R13643 VDD.n2606 VDD.n850 99.5127
R13644 VDD.n2606 VDD.n840 99.5127
R13645 VDD.n2614 VDD.n840 99.5127
R13646 VDD.n2614 VDD.n838 99.5127
R13647 VDD.n2618 VDD.n838 99.5127
R13648 VDD.n2618 VDD.n828 99.5127
R13649 VDD.n2626 VDD.n828 99.5127
R13650 VDD.n2626 VDD.n825 99.5127
R13651 VDD.n2635 VDD.n825 99.5127
R13652 VDD.n2635 VDD.n826 99.5127
R13653 VDD.n826 VDD.n818 99.5127
R13654 VDD.n2630 VDD.n818 99.5127
R13655 VDD.n2630 VDD.n807 99.5127
R13656 VDD.n807 VDD.n798 99.5127
R13657 VDD.n137 VDD.t142 85.8723
R13658 VDD.n124 VDD.t151 85.8723
R13659 VDD.n111 VDD.t160 85.8723
R13660 VDD.n98 VDD.t165 85.8723
R13661 VDD.n85 VDD.t173 85.8723
R13662 VDD.n72 VDD.t136 85.8723
R13663 VDD.n59 VDD.t150 85.8723
R13664 VDD.n46 VDD.t158 85.8723
R13665 VDD.n34 VDD.t167 85.8723
R13666 VDD.n21 VDD.t174 85.8723
R13667 VDD.n1730 VDD.t132 85.8723
R13668 VDD.n1743 VDD.t130 85.8723
R13669 VDD.n1704 VDD.t155 85.8723
R13670 VDD.n1717 VDD.t154 85.8723
R13671 VDD.n1678 VDD.t133 85.8723
R13672 VDD.n1691 VDD.t166 85.8723
R13673 VDD.n1652 VDD.t156 85.8723
R13674 VDD.n1665 VDD.t140 85.8723
R13675 VDD.n1627 VDD.t171 85.8723
R13676 VDD.n1640 VDD.t161 85.8723
R13677 VDD.n3094 VDD.n2744 72.8958
R13678 VDD.n3092 VDD.n2744 72.8958
R13679 VDD.n3086 VDD.n2744 72.8958
R13680 VDD.n3084 VDD.n2744 72.8958
R13681 VDD.n3078 VDD.n2744 72.8958
R13682 VDD.n3076 VDD.n2744 72.8958
R13683 VDD.n3070 VDD.n2744 72.8958
R13684 VDD.n3068 VDD.n2744 72.8958
R13685 VDD.n3062 VDD.n2744 72.8958
R13686 VDD.n3060 VDD.n2744 72.8958
R13687 VDD.n3053 VDD.n2744 72.8958
R13688 VDD.n3345 VDD.n496 72.8958
R13689 VDD.n3353 VDD.n496 72.8958
R13690 VDD.n535 VDD.n496 72.8958
R13691 VDD.n3360 VDD.n496 72.8958
R13692 VDD.n532 VDD.n496 72.8958
R13693 VDD.n3367 VDD.n496 72.8958
R13694 VDD.n3372 VDD.n496 72.8958
R13695 VDD.n529 VDD.n496 72.8958
R13696 VDD.n3379 VDD.n496 72.8958
R13697 VDD.n526 VDD.n496 72.8958
R13698 VDD.n3386 VDD.n496 72.8958
R13699 VDD.n2391 VDD.n2390 72.8958
R13700 VDD.n2390 VDD.n1062 72.8958
R13701 VDD.n2390 VDD.n1063 72.8958
R13702 VDD.n2390 VDD.n1064 72.8958
R13703 VDD.n2390 VDD.n1065 72.8958
R13704 VDD.n2390 VDD.n1066 72.8958
R13705 VDD.n2390 VDD.n1067 72.8958
R13706 VDD.n2390 VDD.n1068 72.8958
R13707 VDD.n2390 VDD.n1069 72.8958
R13708 VDD.n2390 VDD.n1070 72.8958
R13709 VDD.n2743 VDD.n786 72.8958
R13710 VDD.n2743 VDD.n785 72.8958
R13711 VDD.n2743 VDD.n784 72.8958
R13712 VDD.n2743 VDD.n783 72.8958
R13713 VDD.n2743 VDD.n782 72.8958
R13714 VDD.n2743 VDD.n781 72.8958
R13715 VDD.n2743 VDD.n780 72.8958
R13716 VDD.n2743 VDD.n779 72.8958
R13717 VDD.n2743 VDD.n778 72.8958
R13718 VDD.n2743 VDD.n777 72.8958
R13719 VDD.n2743 VDD.n776 72.8958
R13720 VDD.n2790 VDD.n2744 72.8958
R13721 VDD.n2796 VDD.n2744 72.8958
R13722 VDD.n2798 VDD.n2744 72.8958
R13723 VDD.n2804 VDD.n2744 72.8958
R13724 VDD.n2806 VDD.n2744 72.8958
R13725 VDD.n2812 VDD.n2744 72.8958
R13726 VDD.n2814 VDD.n2744 72.8958
R13727 VDD.n2820 VDD.n2744 72.8958
R13728 VDD.n2822 VDD.n2744 72.8958
R13729 VDD.n2831 VDD.n2744 72.8958
R13730 VDD.n3433 VDD.n496 72.8958
R13731 VDD.n504 VDD.n496 72.8958
R13732 VDD.n3440 VDD.n496 72.8958
R13733 VDD.n499 VDD.n496 72.8958
R13734 VDD.n3447 VDD.n496 72.8958
R13735 VDD.n496 VDD.n495 72.8958
R13736 VDD.n3404 VDD.n496 72.8958
R13737 VDD.n3411 VDD.n496 72.8958
R13738 VDD.n3402 VDD.n496 72.8958
R13739 VDD.n3418 VDD.n496 72.8958
R13740 VDD.n3421 VDD.n496 72.8958
R13741 VDD.n2743 VDD.n796 72.8958
R13742 VDD.n2743 VDD.n795 72.8958
R13743 VDD.n2743 VDD.n794 72.8958
R13744 VDD.n2743 VDD.n793 72.8958
R13745 VDD.n2743 VDD.n792 72.8958
R13746 VDD.n2743 VDD.n791 72.8958
R13747 VDD.n2743 VDD.n790 72.8958
R13748 VDD.n2743 VDD.n789 72.8958
R13749 VDD.n2743 VDD.n788 72.8958
R13750 VDD.n2743 VDD.n787 72.8958
R13751 VDD.n2390 VDD.n1072 72.8958
R13752 VDD.n2390 VDD.n1073 72.8958
R13753 VDD.n2390 VDD.n1074 72.8958
R13754 VDD.n2390 VDD.n1075 72.8958
R13755 VDD.n2390 VDD.n1076 72.8958
R13756 VDD.n2390 VDD.n1077 72.8958
R13757 VDD.n2390 VDD.n1078 72.8958
R13758 VDD.n2390 VDD.n1079 72.8958
R13759 VDD.n2390 VDD.n1080 72.8958
R13760 VDD.n2390 VDD.n1081 72.8958
R13761 VDD.n1084 VDD.n1083 70.4005
R13762 VDD.n802 VDD.n801 70.4005
R13763 VDD.n2054 VDD.n2053 70.4005
R13764 VDD.n812 VDD.n811 70.4005
R13765 VDD.n2759 VDD.n2758 70.4005
R13766 VDD.n502 VDD.n501 70.4005
R13767 VDD.n2827 VDD.n2826 70.4005
R13768 VDD.n538 VDD.n537 70.4005
R13769 VDD.n1480 VDD.n1479 66.2847
R13770 VDD.n1480 VDD.n1316 66.2847
R13771 VDD.n1480 VDD.n1317 66.2847
R13772 VDD.n1480 VDD.n1318 66.2847
R13773 VDD.n1480 VDD.n1319 66.2847
R13774 VDD.n1480 VDD.n1320 66.2847
R13775 VDD.n1480 VDD.n1321 66.2847
R13776 VDD.n1480 VDD.n1322 66.2847
R13777 VDD.n1480 VDD.n1323 66.2847
R13778 VDD.n1480 VDD.n1324 66.2847
R13779 VDD.n1480 VDD.n1325 66.2847
R13780 VDD.n1480 VDD.n1326 66.2847
R13781 VDD.n1480 VDD.n1327 66.2847
R13782 VDD.n1480 VDD.n1328 66.2847
R13783 VDD.n1480 VDD.n1329 66.2847
R13784 VDD.n1480 VDD.n1330 66.2847
R13785 VDD.n1480 VDD.n1331 66.2847
R13786 VDD.n1480 VDD.n1332 66.2847
R13787 VDD.n1480 VDD.n1333 66.2847
R13788 VDD.n1480 VDD.n1334 66.2847
R13789 VDD.n1480 VDD.n1335 66.2847
R13790 VDD.n1480 VDD.n1336 66.2847
R13791 VDD.n1098 VDD.n1097 66.2847
R13792 VDD.n1962 VDD.n1098 66.2847
R13793 VDD.n1966 VDD.n1098 66.2847
R13794 VDD.n1970 VDD.n1098 66.2847
R13795 VDD.n1960 VDD.n1098 66.2847
R13796 VDD.n1956 VDD.n1098 66.2847
R13797 VDD.n1981 VDD.n1098 66.2847
R13798 VDD.n1948 VDD.n1098 66.2847
R13799 VDD.n1988 VDD.n1098 66.2847
R13800 VDD.n1941 VDD.n1098 66.2847
R13801 VDD.n1998 VDD.n1098 66.2847
R13802 VDD.n1934 VDD.n1098 66.2847
R13803 VDD.n2005 VDD.n1098 66.2847
R13804 VDD.n1927 VDD.n1098 66.2847
R13805 VDD.n2012 VDD.n1098 66.2847
R13806 VDD.n1920 VDD.n1098 66.2847
R13807 VDD.n2019 VDD.n1098 66.2847
R13808 VDD.n2022 VDD.n1098 66.2847
R13809 VDD.n1909 VDD.n1098 66.2847
R13810 VDD.n2033 VDD.n1098 66.2847
R13811 VDD.n1904 VDD.n1098 66.2847
R13812 VDD.n2203 VDD.n1098 66.2847
R13813 VDD.n1899 VDD.n1098 66.2847
R13814 VDD.n3464 VDD.n448 66.2847
R13815 VDD.n3467 VDD.n448 66.2847
R13816 VDD.n3474 VDD.n448 66.2847
R13817 VDD.n3453 VDD.n448 66.2847
R13818 VDD.n3483 VDD.n448 66.2847
R13819 VDD.n3485 VDD.n448 66.2847
R13820 VDD.n3493 VDD.n448 66.2847
R13821 VDD.n3495 VDD.n448 66.2847
R13822 VDD.n3503 VDD.n448 66.2847
R13823 VDD.n3505 VDD.n448 66.2847
R13824 VDD.n3513 VDD.n448 66.2847
R13825 VDD.n3515 VDD.n448 66.2847
R13826 VDD.n3526 VDD.n448 66.2847
R13827 VDD.n3528 VDD.n448 66.2847
R13828 VDD.n3536 VDD.n448 66.2847
R13829 VDD.n3538 VDD.n448 66.2847
R13830 VDD.n3546 VDD.n448 66.2847
R13831 VDD.n3548 VDD.n448 66.2847
R13832 VDD.n3558 VDD.n448 66.2847
R13833 VDD.n3560 VDD.n448 66.2847
R13834 VDD.n3568 VDD.n448 66.2847
R13835 VDD.n3571 VDD.n448 66.2847
R13836 VDD.n327 VDD.n248 66.2847
R13837 VDD.n3796 VDD.n248 66.2847
R13838 VDD.n321 VDD.n248 66.2847
R13839 VDD.n3803 VDD.n248 66.2847
R13840 VDD.n315 VDD.n248 66.2847
R13841 VDD.n310 VDD.n248 66.2847
R13842 VDD.n3814 VDD.n248 66.2847
R13843 VDD.n302 VDD.n248 66.2847
R13844 VDD.n3821 VDD.n248 66.2847
R13845 VDD.n295 VDD.n248 66.2847
R13846 VDD.n3831 VDD.n248 66.2847
R13847 VDD.n288 VDD.n248 66.2847
R13848 VDD.n3838 VDD.n248 66.2847
R13849 VDD.n3841 VDD.n248 66.2847
R13850 VDD.n279 VDD.n248 66.2847
R13851 VDD.n3850 VDD.n248 66.2847
R13852 VDD.n270 VDD.n248 66.2847
R13853 VDD.n3857 VDD.n248 66.2847
R13854 VDD.n264 VDD.n248 66.2847
R13855 VDD.n3866 VDD.n248 66.2847
R13856 VDD.n256 VDD.n248 66.2847
R13857 VDD.n3873 VDD.n248 66.2847
R13858 VDD.n3876 VDD.n248 66.2847
R13859 VDD.n3876 VDD.n3875 52.4337
R13860 VDD.n3873 VDD.n3872 52.4337
R13861 VDD.n3868 VDD.n256 52.4337
R13862 VDD.n3866 VDD.n3865 52.4337
R13863 VDD.n3859 VDD.n264 52.4337
R13864 VDD.n3857 VDD.n3856 52.4337
R13865 VDD.n3852 VDD.n270 52.4337
R13866 VDD.n3850 VDD.n3849 52.4337
R13867 VDD.n280 VDD.n279 52.4337
R13868 VDD.n3841 VDD.n3840 52.4337
R13869 VDD.n3838 VDD.n3837 52.4337
R13870 VDD.n3833 VDD.n288 52.4337
R13871 VDD.n3831 VDD.n3830 52.4337
R13872 VDD.n3823 VDD.n295 52.4337
R13873 VDD.n3821 VDD.n3820 52.4337
R13874 VDD.n3816 VDD.n302 52.4337
R13875 VDD.n3814 VDD.n3813 52.4337
R13876 VDD.n311 VDD.n310 52.4337
R13877 VDD.n3805 VDD.n315 52.4337
R13878 VDD.n3803 VDD.n3802 52.4337
R13879 VDD.n3798 VDD.n321 52.4337
R13880 VDD.n3796 VDD.n3795 52.4337
R13881 VDD.n3788 VDD.n327 52.4337
R13882 VDD.n3464 VDD.n447 52.4337
R13883 VDD.n3468 VDD.n3467 52.4337
R13884 VDD.n3474 VDD.n3473 52.4337
R13885 VDD.n3454 VDD.n3453 52.4337
R13886 VDD.n3483 VDD.n3482 52.4337
R13887 VDD.n3486 VDD.n3485 52.4337
R13888 VDD.n3493 VDD.n3492 52.4337
R13889 VDD.n3496 VDD.n3495 52.4337
R13890 VDD.n3503 VDD.n3502 52.4337
R13891 VDD.n3506 VDD.n3505 52.4337
R13892 VDD.n3513 VDD.n3512 52.4337
R13893 VDD.n3516 VDD.n3515 52.4337
R13894 VDD.n3526 VDD.n3525 52.4337
R13895 VDD.n3529 VDD.n3528 52.4337
R13896 VDD.n3536 VDD.n3535 52.4337
R13897 VDD.n3539 VDD.n3538 52.4337
R13898 VDD.n3546 VDD.n3545 52.4337
R13899 VDD.n3549 VDD.n3548 52.4337
R13900 VDD.n3558 VDD.n3557 52.4337
R13901 VDD.n3561 VDD.n3560 52.4337
R13902 VDD.n3568 VDD.n3567 52.4337
R13903 VDD.n3571 VDD.n3570 52.4337
R13904 VDD.n2205 VDD.n1899 52.4337
R13905 VDD.n2203 VDD.n2202 52.4337
R13906 VDD.n2035 VDD.n1904 52.4337
R13907 VDD.n2033 VDD.n2032 52.4337
R13908 VDD.n1910 VDD.n1909 52.4337
R13909 VDD.n2022 VDD.n2021 52.4337
R13910 VDD.n2019 VDD.n2018 52.4337
R13911 VDD.n2014 VDD.n1920 52.4337
R13912 VDD.n2012 VDD.n2011 52.4337
R13913 VDD.n2007 VDD.n1927 52.4337
R13914 VDD.n2005 VDD.n2004 52.4337
R13915 VDD.n2000 VDD.n1934 52.4337
R13916 VDD.n1998 VDD.n1997 52.4337
R13917 VDD.n1990 VDD.n1941 52.4337
R13918 VDD.n1988 VDD.n1987 52.4337
R13919 VDD.n1983 VDD.n1948 52.4337
R13920 VDD.n1981 VDD.n1980 52.4337
R13921 VDD.n1957 VDD.n1956 52.4337
R13922 VDD.n1972 VDD.n1960 52.4337
R13923 VDD.n1970 VDD.n1969 52.4337
R13924 VDD.n1966 VDD.n1965 52.4337
R13925 VDD.n1962 VDD.n1090 52.4337
R13926 VDD.n1097 VDD.n1092 52.4337
R13927 VDD.n1479 VDD.n1478 52.4337
R13928 VDD.n1342 VDD.n1316 52.4337
R13929 VDD.n1344 VDD.n1317 52.4337
R13930 VDD.n1463 VDD.n1318 52.4337
R13931 VDD.n1348 VDD.n1319 52.4337
R13932 VDD.n1352 VDD.n1320 52.4337
R13933 VDD.n1354 VDD.n1321 52.4337
R13934 VDD.n1358 VDD.n1322 52.4337
R13935 VDD.n1445 VDD.n1323 52.4337
R13936 VDD.n1362 VDD.n1324 52.4337
R13937 VDD.n1364 VDD.n1325 52.4337
R13938 VDD.n1368 VDD.n1326 52.4337
R13939 VDD.n1370 VDD.n1327 52.4337
R13940 VDD.n1376 VDD.n1328 52.4337
R13941 VDD.n1378 VDD.n1329 52.4337
R13942 VDD.n1382 VDD.n1330 52.4337
R13943 VDD.n1384 VDD.n1331 52.4337
R13944 VDD.n1413 VDD.n1332 52.4337
R13945 VDD.n1389 VDD.n1333 52.4337
R13946 VDD.n1393 VDD.n1334 52.4337
R13947 VDD.n1395 VDD.n1335 52.4337
R13948 VDD.n1399 VDD.n1336 52.4337
R13949 VDD.n1479 VDD.n1338 52.4337
R13950 VDD.n1343 VDD.n1316 52.4337
R13951 VDD.n1462 VDD.n1317 52.4337
R13952 VDD.n1347 VDD.n1318 52.4337
R13953 VDD.n1351 VDD.n1319 52.4337
R13954 VDD.n1353 VDD.n1320 52.4337
R13955 VDD.n1357 VDD.n1321 52.4337
R13956 VDD.n1446 VDD.n1322 52.4337
R13957 VDD.n1361 VDD.n1323 52.4337
R13958 VDD.n1363 VDD.n1324 52.4337
R13959 VDD.n1367 VDD.n1325 52.4337
R13960 VDD.n1369 VDD.n1326 52.4337
R13961 VDD.n1375 VDD.n1327 52.4337
R13962 VDD.n1377 VDD.n1328 52.4337
R13963 VDD.n1381 VDD.n1329 52.4337
R13964 VDD.n1383 VDD.n1330 52.4337
R13965 VDD.n1387 VDD.n1331 52.4337
R13966 VDD.n1388 VDD.n1332 52.4337
R13967 VDD.n1392 VDD.n1333 52.4337
R13968 VDD.n1394 VDD.n1334 52.4337
R13969 VDD.n1398 VDD.n1335 52.4337
R13970 VDD.n1336 VDD.n1315 52.4337
R13971 VDD.n1097 VDD.n1091 52.4337
R13972 VDD.n1963 VDD.n1962 52.4337
R13973 VDD.n1967 VDD.n1966 52.4337
R13974 VDD.n1971 VDD.n1970 52.4337
R13975 VDD.n1960 VDD.n1959 52.4337
R13976 VDD.n1956 VDD.n1949 52.4337
R13977 VDD.n1982 VDD.n1981 52.4337
R13978 VDD.n1948 VDD.n1942 52.4337
R13979 VDD.n1989 VDD.n1988 52.4337
R13980 VDD.n1941 VDD.n1935 52.4337
R13981 VDD.n1999 VDD.n1998 52.4337
R13982 VDD.n1934 VDD.n1928 52.4337
R13983 VDD.n2006 VDD.n2005 52.4337
R13984 VDD.n1927 VDD.n1921 52.4337
R13985 VDD.n2013 VDD.n2012 52.4337
R13986 VDD.n1920 VDD.n1912 52.4337
R13987 VDD.n2020 VDD.n2019 52.4337
R13988 VDD.n2023 VDD.n2022 52.4337
R13989 VDD.n1909 VDD.n1905 52.4337
R13990 VDD.n2034 VDD.n2033 52.4337
R13991 VDD.n1904 VDD.n1900 52.4337
R13992 VDD.n2204 VDD.n2203 52.4337
R13993 VDD.n1899 VDD.n1100 52.4337
R13994 VDD.n3465 VDD.n3464 52.4337
R13995 VDD.n3467 VDD.n3458 52.4337
R13996 VDD.n3475 VDD.n3474 52.4337
R13997 VDD.n3453 VDD.n491 52.4337
R13998 VDD.n3484 VDD.n3483 52.4337
R13999 VDD.n3485 VDD.n487 52.4337
R14000 VDD.n3494 VDD.n3493 52.4337
R14001 VDD.n3495 VDD.n481 52.4337
R14002 VDD.n3504 VDD.n3503 52.4337
R14003 VDD.n3505 VDD.n477 52.4337
R14004 VDD.n3514 VDD.n3513 52.4337
R14005 VDD.n3515 VDD.n473 52.4337
R14006 VDD.n3527 VDD.n3526 52.4337
R14007 VDD.n3528 VDD.n469 52.4337
R14008 VDD.n3537 VDD.n3536 52.4337
R14009 VDD.n3538 VDD.n465 52.4337
R14010 VDD.n3547 VDD.n3546 52.4337
R14011 VDD.n3548 VDD.n461 52.4337
R14012 VDD.n3559 VDD.n3558 52.4337
R14013 VDD.n3560 VDD.n455 52.4337
R14014 VDD.n3569 VDD.n3568 52.4337
R14015 VDD.n3572 VDD.n3571 52.4337
R14016 VDD.n327 VDD.n322 52.4337
R14017 VDD.n3797 VDD.n3796 52.4337
R14018 VDD.n321 VDD.n316 52.4337
R14019 VDD.n3804 VDD.n3803 52.4337
R14020 VDD.n315 VDD.n314 52.4337
R14021 VDD.n310 VDD.n303 52.4337
R14022 VDD.n3815 VDD.n3814 52.4337
R14023 VDD.n302 VDD.n296 52.4337
R14024 VDD.n3822 VDD.n3821 52.4337
R14025 VDD.n295 VDD.n289 52.4337
R14026 VDD.n3832 VDD.n3831 52.4337
R14027 VDD.n288 VDD.n282 52.4337
R14028 VDD.n3839 VDD.n3838 52.4337
R14029 VDD.n3842 VDD.n3841 52.4337
R14030 VDD.n279 VDD.n271 52.4337
R14031 VDD.n3851 VDD.n3850 52.4337
R14032 VDD.n270 VDD.n265 52.4337
R14033 VDD.n3858 VDD.n3857 52.4337
R14034 VDD.n264 VDD.n257 52.4337
R14035 VDD.n3867 VDD.n3866 52.4337
R14036 VDD.n256 VDD.n250 52.4337
R14037 VDD.n3874 VDD.n3873 52.4337
R14038 VDD.n3877 VDD.n3876 52.4337
R14039 VDD.n3421 VDD.n3420 39.2114
R14040 VDD.n3418 VDD.n3417 39.2114
R14041 VDD.n3413 VDD.n3402 39.2114
R14042 VDD.n3411 VDD.n3410 39.2114
R14043 VDD.n3406 VDD.n3404 39.2114
R14044 VDD.n3449 VDD.n495 39.2114
R14045 VDD.n3447 VDD.n3446 39.2114
R14046 VDD.n3442 VDD.n499 39.2114
R14047 VDD.n3440 VDD.n3439 39.2114
R14048 VDD.n3435 VDD.n504 39.2114
R14049 VDD.n3433 VDD.n3432 39.2114
R14050 VDD.n2790 VDD.n774 39.2114
R14051 VDD.n2796 VDD.n2795 39.2114
R14052 VDD.n2799 VDD.n2798 39.2114
R14053 VDD.n2804 VDD.n2803 39.2114
R14054 VDD.n2807 VDD.n2806 39.2114
R14055 VDD.n2812 VDD.n2811 39.2114
R14056 VDD.n2815 VDD.n2814 39.2114
R14057 VDD.n2820 VDD.n2819 39.2114
R14058 VDD.n2823 VDD.n2822 39.2114
R14059 VDD.n2831 VDD.n2830 39.2114
R14060 VDD.n2689 VDD.n776 39.2114
R14061 VDD.n2685 VDD.n777 39.2114
R14062 VDD.n2681 VDD.n778 39.2114
R14063 VDD.n2677 VDD.n779 39.2114
R14064 VDD.n2673 VDD.n780 39.2114
R14065 VDD.n2669 VDD.n781 39.2114
R14066 VDD.n2665 VDD.n782 39.2114
R14067 VDD.n2661 VDD.n783 39.2114
R14068 VDD.n2657 VDD.n784 39.2114
R14069 VDD.n2653 VDD.n785 39.2114
R14070 VDD.n2649 VDD.n786 39.2114
R14071 VDD.n2391 VDD.n1059 39.2114
R14072 VDD.n2038 VDD.n1062 39.2114
R14073 VDD.n2042 VDD.n1063 39.2114
R14074 VDD.n2046 VDD.n1064 39.2114
R14075 VDD.n2050 VDD.n1065 39.2114
R14076 VDD.n2195 VDD.n1066 39.2114
R14077 VDD.n2191 VDD.n1067 39.2114
R14078 VDD.n2187 VDD.n1068 39.2114
R14079 VDD.n2183 VDD.n1069 39.2114
R14080 VDD.n2179 VDD.n1070 39.2114
R14081 VDD.n3386 VDD.n3385 39.2114
R14082 VDD.n3381 VDD.n526 39.2114
R14083 VDD.n3379 VDD.n3378 39.2114
R14084 VDD.n3374 VDD.n529 39.2114
R14085 VDD.n3372 VDD.n3371 39.2114
R14086 VDD.n3367 VDD.n3366 39.2114
R14087 VDD.n3362 VDD.n532 39.2114
R14088 VDD.n3360 VDD.n3359 39.2114
R14089 VDD.n3355 VDD.n535 39.2114
R14090 VDD.n3353 VDD.n3352 39.2114
R14091 VDD.n3347 VDD.n3345 39.2114
R14092 VDD.n3094 VDD.n2747 39.2114
R14093 VDD.n3093 VDD.n3092 39.2114
R14094 VDD.n3086 VDD.n2749 39.2114
R14095 VDD.n3085 VDD.n3084 39.2114
R14096 VDD.n3078 VDD.n2751 39.2114
R14097 VDD.n3077 VDD.n3076 39.2114
R14098 VDD.n3070 VDD.n2753 39.2114
R14099 VDD.n3069 VDD.n3068 39.2114
R14100 VDD.n3062 VDD.n2755 39.2114
R14101 VDD.n3061 VDD.n3060 39.2114
R14102 VDD.n3053 VDD.n2757 39.2114
R14103 VDD.n3095 VDD.n3094 39.2114
R14104 VDD.n3092 VDD.n3091 39.2114
R14105 VDD.n3087 VDD.n3086 39.2114
R14106 VDD.n3084 VDD.n3083 39.2114
R14107 VDD.n3079 VDD.n3078 39.2114
R14108 VDD.n3076 VDD.n3075 39.2114
R14109 VDD.n3071 VDD.n3070 39.2114
R14110 VDD.n3068 VDD.n3067 39.2114
R14111 VDD.n3063 VDD.n3062 39.2114
R14112 VDD.n3060 VDD.n3059 39.2114
R14113 VDD.n3054 VDD.n3053 39.2114
R14114 VDD.n3345 VDD.n536 39.2114
R14115 VDD.n3354 VDD.n3353 39.2114
R14116 VDD.n535 VDD.n533 39.2114
R14117 VDD.n3361 VDD.n3360 39.2114
R14118 VDD.n532 VDD.n530 39.2114
R14119 VDD.n3368 VDD.n3367 39.2114
R14120 VDD.n3373 VDD.n3372 39.2114
R14121 VDD.n529 VDD.n527 39.2114
R14122 VDD.n3380 VDD.n3379 39.2114
R14123 VDD.n526 VDD.n524 39.2114
R14124 VDD.n3387 VDD.n3386 39.2114
R14125 VDD.n2392 VDD.n2391 39.2114
R14126 VDD.n2041 VDD.n1062 39.2114
R14127 VDD.n2045 VDD.n1063 39.2114
R14128 VDD.n2049 VDD.n1064 39.2114
R14129 VDD.n2194 VDD.n1065 39.2114
R14130 VDD.n2192 VDD.n1066 39.2114
R14131 VDD.n2188 VDD.n1067 39.2114
R14132 VDD.n2184 VDD.n1068 39.2114
R14133 VDD.n2180 VDD.n1069 39.2114
R14134 VDD.n2175 VDD.n1070 39.2114
R14135 VDD.n2652 VDD.n786 39.2114
R14136 VDD.n2656 VDD.n785 39.2114
R14137 VDD.n2660 VDD.n784 39.2114
R14138 VDD.n2664 VDD.n783 39.2114
R14139 VDD.n2668 VDD.n782 39.2114
R14140 VDD.n2672 VDD.n781 39.2114
R14141 VDD.n2676 VDD.n780 39.2114
R14142 VDD.n2680 VDD.n779 39.2114
R14143 VDD.n2684 VDD.n778 39.2114
R14144 VDD.n2688 VDD.n777 39.2114
R14145 VDD.n2691 VDD.n776 39.2114
R14146 VDD.n2791 VDD.n2790 39.2114
R14147 VDD.n2797 VDD.n2796 39.2114
R14148 VDD.n2798 VDD.n2787 39.2114
R14149 VDD.n2805 VDD.n2804 39.2114
R14150 VDD.n2806 VDD.n2785 39.2114
R14151 VDD.n2813 VDD.n2812 39.2114
R14152 VDD.n2814 VDD.n2783 39.2114
R14153 VDD.n2821 VDD.n2820 39.2114
R14154 VDD.n2822 VDD.n2781 39.2114
R14155 VDD.n2832 VDD.n2831 39.2114
R14156 VDD.n3434 VDD.n3433 39.2114
R14157 VDD.n504 VDD.n500 39.2114
R14158 VDD.n3441 VDD.n3440 39.2114
R14159 VDD.n499 VDD.n497 39.2114
R14160 VDD.n3448 VDD.n3447 39.2114
R14161 VDD.n3405 VDD.n495 39.2114
R14162 VDD.n3404 VDD.n3403 39.2114
R14163 VDD.n3412 VDD.n3411 39.2114
R14164 VDD.n3402 VDD.n3400 39.2114
R14165 VDD.n3419 VDD.n3418 39.2114
R14166 VDD.n3422 VDD.n3421 39.2114
R14167 VDD.n799 VDD.n787 39.2114
R14168 VDD.n2737 VDD.n788 39.2114
R14169 VDD.n2733 VDD.n789 39.2114
R14170 VDD.n2729 VDD.n790 39.2114
R14171 VDD.n2725 VDD.n791 39.2114
R14172 VDD.n2721 VDD.n792 39.2114
R14173 VDD.n2717 VDD.n793 39.2114
R14174 VDD.n2713 VDD.n794 39.2114
R14175 VDD.n2709 VDD.n795 39.2114
R14176 VDD.n2705 VDD.n796 39.2114
R14177 VDD.n2226 VDD.n1072 39.2114
R14178 VDD.n2230 VDD.n1073 39.2114
R14179 VDD.n2234 VDD.n1074 39.2114
R14180 VDD.n2238 VDD.n1075 39.2114
R14181 VDD.n2242 VDD.n1076 39.2114
R14182 VDD.n2246 VDD.n1077 39.2114
R14183 VDD.n2250 VDD.n1078 39.2114
R14184 VDD.n2254 VDD.n1079 39.2114
R14185 VDD.n2258 VDD.n1080 39.2114
R14186 VDD.n2262 VDD.n1081 39.2114
R14187 VDD.n2701 VDD.n796 39.2114
R14188 VDD.n2706 VDD.n795 39.2114
R14189 VDD.n2710 VDD.n794 39.2114
R14190 VDD.n2714 VDD.n793 39.2114
R14191 VDD.n2718 VDD.n792 39.2114
R14192 VDD.n2722 VDD.n791 39.2114
R14193 VDD.n2726 VDD.n790 39.2114
R14194 VDD.n2730 VDD.n789 39.2114
R14195 VDD.n2734 VDD.n788 39.2114
R14196 VDD.n2738 VDD.n787 39.2114
R14197 VDD.n2229 VDD.n1072 39.2114
R14198 VDD.n2233 VDD.n1073 39.2114
R14199 VDD.n2237 VDD.n1074 39.2114
R14200 VDD.n2241 VDD.n1075 39.2114
R14201 VDD.n2245 VDD.n1076 39.2114
R14202 VDD.n2249 VDD.n1077 39.2114
R14203 VDD.n2253 VDD.n1078 39.2114
R14204 VDD.n2257 VDD.n1079 39.2114
R14205 VDD.n2261 VDD.n1080 39.2114
R14206 VDD.n1082 VDD.n1081 39.2114
R14207 VDD.n131 VDD.n129 37.9395
R14208 VDD.n105 VDD.n103 37.9395
R14209 VDD.n79 VDD.n77 37.9395
R14210 VDD.n53 VDD.n51 37.9395
R14211 VDD.n28 VDD.n26 37.9395
R14212 VDD.n1737 VDD.n1735 37.9395
R14213 VDD.n1711 VDD.n1709 37.9395
R14214 VDD.n1685 VDD.n1683 37.9395
R14215 VDD.n1659 VDD.n1657 37.9395
R14216 VDD.n1634 VDD.n1632 37.9395
R14217 VDD.n1314 VDD.n1313 37.2369
R14218 VDD.n1416 VDD.n1415 37.2369
R14219 VDD.n1373 VDD.n1372 37.2369
R14220 VDD.n1449 VDD.n1448 37.2369
R14221 VDD.n1466 VDD.n1465 37.2369
R14222 VDD.n2220 VDD.n2219 37.2369
R14223 VDD.n1977 VDD.n1955 37.2369
R14224 VDD.n1995 VDD.n1994 37.2369
R14225 VDD.n1919 VDD.n1918 37.2369
R14226 VDD.n2031 VDD.n2030 37.2369
R14227 VDD.n3792 VDD.n3791 37.2369
R14228 VDD.n3810 VDD.n309 37.2369
R14229 VDD.n3828 VDD.n3827 37.2369
R14230 VDD.n3847 VDD.n276 37.2369
R14231 VDD.n3864 VDD.n260 37.2369
R14232 VDD.n484 VDD.n483 37.2369
R14233 VDD.n3523 VDD.n3522 37.2369
R14234 VDD.n3552 VDD.n3551 37.2369
R14235 VDD.n3477 VDD.n3456 37.2369
R14236 VDD.n3574 VDD.n452 37.2369
R14237 VDD.n143 VDD.n142 33.155
R14238 VDD.n117 VDD.n116 33.155
R14239 VDD.n91 VDD.n90 33.155
R14240 VDD.n65 VDD.n64 33.155
R14241 VDD.n40 VDD.n39 33.155
R14242 VDD.n1749 VDD.n1748 33.155
R14243 VDD.n1723 VDD.n1722 33.155
R14244 VDD.n1697 VDD.n1696 33.155
R14245 VDD.n1671 VDD.n1670 33.155
R14246 VDD.n1646 VDD.n1645 33.155
R14247 VDD.n1480 VDD.n1308 33.0591
R14248 VDD.n2212 VDD.n1098 33.0591
R14249 VDD.n3580 VDD.n448 33.0591
R14250 VDD.n248 VDD.n242 33.0591
R14251 VDD.n2395 VDD.n2394 31.8444
R14252 VDD.n2693 VDD.n2692 31.8444
R14253 VDD.n2650 VDD.n2647 31.8444
R14254 VDD.n2174 VDD.n2173 31.8444
R14255 VDD.n2835 VDD.n2834 31.8444
R14256 VDD.n3431 VDD.n3430 31.8444
R14257 VDD.n3102 VDD.n773 31.8444
R14258 VDD.n3424 VDD.n3423 31.8444
R14259 VDD.n3389 VDD.n523 31.8444
R14260 VDD.n3348 VDD.n3344 31.8444
R14261 VDD.n3055 VDD.n3052 31.8444
R14262 VDD.n3098 VDD.n3097 31.8444
R14263 VDD.n2399 VDD.n1055 31.8444
R14264 VDD.n2741 VDD.n800 31.8444
R14265 VDD.n2700 VDD.n2699 31.8444
R14266 VDD.n2388 VDD.n2387 31.8444
R14267 VDD.n2264 VDD.n1084 30.449
R14268 VDD.n2703 VDD.n802 30.449
R14269 VDD.n2177 VDD.n2054 30.449
R14270 VDD.n813 VDD.n812 30.449
R14271 VDD.n3057 VDD.n2759 30.449
R14272 VDD.n503 VDD.n502 30.449
R14273 VDD.n2828 VDD.n2827 30.449
R14274 VDD.n3350 VDD.n538 30.449
R14275 VDD.n2743 VDD.n775 23.4895
R14276 VDD.n3100 VDD.n2744 23.4895
R14277 VDD.n1486 VDD.n1310 19.3944
R14278 VDD.n1486 VDD.n1300 19.3944
R14279 VDD.n1498 VDD.n1300 19.3944
R14280 VDD.n1498 VDD.n1298 19.3944
R14281 VDD.n1502 VDD.n1298 19.3944
R14282 VDD.n1502 VDD.n1288 19.3944
R14283 VDD.n1514 VDD.n1288 19.3944
R14284 VDD.n1514 VDD.n1286 19.3944
R14285 VDD.n1518 VDD.n1286 19.3944
R14286 VDD.n1518 VDD.n1276 19.3944
R14287 VDD.n1530 VDD.n1276 19.3944
R14288 VDD.n1530 VDD.n1274 19.3944
R14289 VDD.n1534 VDD.n1274 19.3944
R14290 VDD.n1534 VDD.n1264 19.3944
R14291 VDD.n1546 VDD.n1264 19.3944
R14292 VDD.n1546 VDD.n1262 19.3944
R14293 VDD.n1550 VDD.n1262 19.3944
R14294 VDD.n1550 VDD.n1253 19.3944
R14295 VDD.n1563 VDD.n1253 19.3944
R14296 VDD.n1563 VDD.n1251 19.3944
R14297 VDD.n1567 VDD.n1251 19.3944
R14298 VDD.n1567 VDD.n1241 19.3944
R14299 VDD.n1579 VDD.n1241 19.3944
R14300 VDD.n1579 VDD.n1239 19.3944
R14301 VDD.n1583 VDD.n1239 19.3944
R14302 VDD.n1583 VDD.n1229 19.3944
R14303 VDD.n1595 VDD.n1229 19.3944
R14304 VDD.n1595 VDD.n1227 19.3944
R14305 VDD.n1599 VDD.n1227 19.3944
R14306 VDD.n1599 VDD.n1217 19.3944
R14307 VDD.n1611 VDD.n1217 19.3944
R14308 VDD.n1611 VDD.n1215 19.3944
R14309 VDD.n1615 VDD.n1215 19.3944
R14310 VDD.n1615 VDD.n1205 19.3944
R14311 VDD.n1758 VDD.n1205 19.3944
R14312 VDD.n1758 VDD.n1203 19.3944
R14313 VDD.n1762 VDD.n1203 19.3944
R14314 VDD.n1762 VDD.n1193 19.3944
R14315 VDD.n1774 VDD.n1193 19.3944
R14316 VDD.n1774 VDD.n1191 19.3944
R14317 VDD.n1778 VDD.n1191 19.3944
R14318 VDD.n1778 VDD.n1181 19.3944
R14319 VDD.n1790 VDD.n1181 19.3944
R14320 VDD.n1790 VDD.n1179 19.3944
R14321 VDD.n1794 VDD.n1179 19.3944
R14322 VDD.n1794 VDD.n1169 19.3944
R14323 VDD.n1806 VDD.n1169 19.3944
R14324 VDD.n1806 VDD.n1167 19.3944
R14325 VDD.n1810 VDD.n1167 19.3944
R14326 VDD.n1810 VDD.n1156 19.3944
R14327 VDD.n1822 VDD.n1156 19.3944
R14328 VDD.n1822 VDD.n1154 19.3944
R14329 VDD.n1826 VDD.n1154 19.3944
R14330 VDD.n1826 VDD.n1145 19.3944
R14331 VDD.n1838 VDD.n1145 19.3944
R14332 VDD.n1838 VDD.n1143 19.3944
R14333 VDD.n1842 VDD.n1143 19.3944
R14334 VDD.n1842 VDD.n1133 19.3944
R14335 VDD.n1854 VDD.n1133 19.3944
R14336 VDD.n1854 VDD.n1131 19.3944
R14337 VDD.n1858 VDD.n1131 19.3944
R14338 VDD.n1858 VDD.n1121 19.3944
R14339 VDD.n1870 VDD.n1121 19.3944
R14340 VDD.n1870 VDD.n1119 19.3944
R14341 VDD.n1874 VDD.n1119 19.3944
R14342 VDD.n1874 VDD.n1109 19.3944
R14343 VDD.n1886 VDD.n1109 19.3944
R14344 VDD.n1886 VDD.n1107 19.3944
R14345 VDD.n1890 VDD.n1107 19.3944
R14346 VDD.n1890 VDD.n1094 19.3944
R14347 VDD.n2214 VDD.n1094 19.3944
R14348 VDD.n1412 VDD.n1390 19.3944
R14349 VDD.n1408 VDD.n1390 19.3944
R14350 VDD.n1408 VDD.n1407 19.3944
R14351 VDD.n1407 VDD.n1406 19.3944
R14352 VDD.n1406 VDD.n1396 19.3944
R14353 VDD.n1402 VDD.n1396 19.3944
R14354 VDD.n1402 VDD.n1401 19.3944
R14355 VDD.n1401 VDD.n1400 19.3944
R14356 VDD.n1429 VDD.n1428 19.3944
R14357 VDD.n1428 VDD.n1427 19.3944
R14358 VDD.n1427 VDD.n1379 19.3944
R14359 VDD.n1423 VDD.n1379 19.3944
R14360 VDD.n1423 VDD.n1422 19.3944
R14361 VDD.n1422 VDD.n1421 19.3944
R14362 VDD.n1421 VDD.n1385 19.3944
R14363 VDD.n1417 VDD.n1385 19.3944
R14364 VDD.n1444 VDD.n1359 19.3944
R14365 VDD.n1440 VDD.n1359 19.3944
R14366 VDD.n1440 VDD.n1439 19.3944
R14367 VDD.n1439 VDD.n1438 19.3944
R14368 VDD.n1438 VDD.n1365 19.3944
R14369 VDD.n1434 VDD.n1365 19.3944
R14370 VDD.n1434 VDD.n1433 19.3944
R14371 VDD.n1433 VDD.n1432 19.3944
R14372 VDD.n1461 VDD.n1460 19.3944
R14373 VDD.n1460 VDD.n1349 19.3944
R14374 VDD.n1456 VDD.n1349 19.3944
R14375 VDD.n1456 VDD.n1455 19.3944
R14376 VDD.n1455 VDD.n1454 19.3944
R14377 VDD.n1454 VDD.n1355 19.3944
R14378 VDD.n1450 VDD.n1355 19.3944
R14379 VDD.n1477 VDD.n1476 19.3944
R14380 VDD.n1476 VDD.n1340 19.3944
R14381 VDD.n1472 VDD.n1340 19.3944
R14382 VDD.n1472 VDD.n1471 19.3944
R14383 VDD.n1471 VDD.n1470 19.3944
R14384 VDD.n1470 VDD.n1345 19.3944
R14385 VDD.n1973 VDD.n1953 19.3944
R14386 VDD.n1973 VDD.n1958 19.3944
R14387 VDD.n1968 VDD.n1958 19.3944
R14388 VDD.n1964 VDD.n1961 19.3944
R14389 VDD.n2222 VDD.n1089 19.3944
R14390 VDD.n2222 VDD.n2221 19.3944
R14391 VDD.n1992 VDD.n1991 19.3944
R14392 VDD.n1991 VDD.n1940 19.3944
R14393 VDD.n1986 VDD.n1940 19.3944
R14394 VDD.n1986 VDD.n1985 19.3944
R14395 VDD.n1985 VDD.n1984 19.3944
R14396 VDD.n1984 VDD.n1947 19.3944
R14397 VDD.n1979 VDD.n1947 19.3944
R14398 VDD.n1979 VDD.n1978 19.3944
R14399 VDD.n2010 VDD.n2009 19.3944
R14400 VDD.n2009 VDD.n2008 19.3944
R14401 VDD.n2008 VDD.n1926 19.3944
R14402 VDD.n2003 VDD.n1926 19.3944
R14403 VDD.n2003 VDD.n2002 19.3944
R14404 VDD.n2002 VDD.n2001 19.3944
R14405 VDD.n2001 VDD.n1933 19.3944
R14406 VDD.n1996 VDD.n1933 19.3944
R14407 VDD.n2028 VDD.n1906 19.3944
R14408 VDD.n2024 VDD.n1906 19.3944
R14409 VDD.n2024 VDD.n1908 19.3944
R14410 VDD.n1911 VDD.n1908 19.3944
R14411 VDD.n2017 VDD.n1911 19.3944
R14412 VDD.n2017 VDD.n2016 19.3944
R14413 VDD.n2016 VDD.n2015 19.3944
R14414 VDD.n2207 VDD.n2206 19.3944
R14415 VDD.n2206 VDD.n1898 19.3944
R14416 VDD.n2201 VDD.n1898 19.3944
R14417 VDD.n2036 VDD.n1901 19.3944
R14418 VDD.n1490 VDD.n1306 19.3944
R14419 VDD.n1490 VDD.n1304 19.3944
R14420 VDD.n1494 VDD.n1304 19.3944
R14421 VDD.n1494 VDD.n1294 19.3944
R14422 VDD.n1506 VDD.n1294 19.3944
R14423 VDD.n1506 VDD.n1292 19.3944
R14424 VDD.n1510 VDD.n1292 19.3944
R14425 VDD.n1510 VDD.n1282 19.3944
R14426 VDD.n1522 VDD.n1282 19.3944
R14427 VDD.n1522 VDD.n1280 19.3944
R14428 VDD.n1526 VDD.n1280 19.3944
R14429 VDD.n1526 VDD.n1270 19.3944
R14430 VDD.n1538 VDD.n1270 19.3944
R14431 VDD.n1538 VDD.n1268 19.3944
R14432 VDD.n1542 VDD.n1268 19.3944
R14433 VDD.n1542 VDD.n1258 19.3944
R14434 VDD.n1555 VDD.n1258 19.3944
R14435 VDD.n1555 VDD.n1256 19.3944
R14436 VDD.n1559 VDD.n1256 19.3944
R14437 VDD.n1559 VDD.n1247 19.3944
R14438 VDD.n1571 VDD.n1247 19.3944
R14439 VDD.n1571 VDD.n1245 19.3944
R14440 VDD.n1575 VDD.n1245 19.3944
R14441 VDD.n1575 VDD.n1235 19.3944
R14442 VDD.n1587 VDD.n1235 19.3944
R14443 VDD.n1587 VDD.n1233 19.3944
R14444 VDD.n1591 VDD.n1233 19.3944
R14445 VDD.n1591 VDD.n1223 19.3944
R14446 VDD.n1603 VDD.n1223 19.3944
R14447 VDD.n1603 VDD.n1221 19.3944
R14448 VDD.n1607 VDD.n1221 19.3944
R14449 VDD.n1607 VDD.n1211 19.3944
R14450 VDD.n1619 VDD.n1211 19.3944
R14451 VDD.n1619 VDD.n1209 19.3944
R14452 VDD.n1754 VDD.n1209 19.3944
R14453 VDD.n1754 VDD.n1199 19.3944
R14454 VDD.n1766 VDD.n1199 19.3944
R14455 VDD.n1766 VDD.n1197 19.3944
R14456 VDD.n1770 VDD.n1197 19.3944
R14457 VDD.n1770 VDD.n1187 19.3944
R14458 VDD.n1782 VDD.n1187 19.3944
R14459 VDD.n1782 VDD.n1185 19.3944
R14460 VDD.n1786 VDD.n1185 19.3944
R14461 VDD.n1786 VDD.n1175 19.3944
R14462 VDD.n1798 VDD.n1175 19.3944
R14463 VDD.n1798 VDD.n1173 19.3944
R14464 VDD.n1802 VDD.n1173 19.3944
R14465 VDD.n1802 VDD.n1163 19.3944
R14466 VDD.n1814 VDD.n1163 19.3944
R14467 VDD.n1814 VDD.n1161 19.3944
R14468 VDD.n1818 VDD.n1161 19.3944
R14469 VDD.n1818 VDD.n1151 19.3944
R14470 VDD.n1830 VDD.n1151 19.3944
R14471 VDD.n1830 VDD.n1149 19.3944
R14472 VDD.n1834 VDD.n1149 19.3944
R14473 VDD.n1834 VDD.n1139 19.3944
R14474 VDD.n1846 VDD.n1139 19.3944
R14475 VDD.n1846 VDD.n1137 19.3944
R14476 VDD.n1850 VDD.n1137 19.3944
R14477 VDD.n1850 VDD.n1127 19.3944
R14478 VDD.n1862 VDD.n1127 19.3944
R14479 VDD.n1862 VDD.n1125 19.3944
R14480 VDD.n1866 VDD.n1125 19.3944
R14481 VDD.n1866 VDD.n1115 19.3944
R14482 VDD.n1878 VDD.n1115 19.3944
R14483 VDD.n1878 VDD.n1113 19.3944
R14484 VDD.n1882 VDD.n1113 19.3944
R14485 VDD.n1882 VDD.n1103 19.3944
R14486 VDD.n1894 VDD.n1103 19.3944
R14487 VDD.n1894 VDD.n1101 19.3944
R14488 VDD.n2210 VDD.n1101 19.3944
R14489 VDD.n3578 VDD.n441 19.3944
R14490 VDD.n3590 VDD.n441 19.3944
R14491 VDD.n3590 VDD.n439 19.3944
R14492 VDD.n3594 VDD.n439 19.3944
R14493 VDD.n3594 VDD.n430 19.3944
R14494 VDD.n3607 VDD.n430 19.3944
R14495 VDD.n3607 VDD.n428 19.3944
R14496 VDD.n3611 VDD.n428 19.3944
R14497 VDD.n3611 VDD.n418 19.3944
R14498 VDD.n3623 VDD.n418 19.3944
R14499 VDD.n3623 VDD.n416 19.3944
R14500 VDD.n3627 VDD.n416 19.3944
R14501 VDD.n3627 VDD.n406 19.3944
R14502 VDD.n3639 VDD.n406 19.3944
R14503 VDD.n3639 VDD.n404 19.3944
R14504 VDD.n3643 VDD.n404 19.3944
R14505 VDD.n3643 VDD.n394 19.3944
R14506 VDD.n3655 VDD.n394 19.3944
R14507 VDD.n3655 VDD.n392 19.3944
R14508 VDD.n3659 VDD.n392 19.3944
R14509 VDD.n3659 VDD.n382 19.3944
R14510 VDD.n3671 VDD.n382 19.3944
R14511 VDD.n3671 VDD.n380 19.3944
R14512 VDD.n3675 VDD.n380 19.3944
R14513 VDD.n3675 VDD.n370 19.3944
R14514 VDD.n3687 VDD.n370 19.3944
R14515 VDD.n3687 VDD.n368 19.3944
R14516 VDD.n3691 VDD.n368 19.3944
R14517 VDD.n3691 VDD.n359 19.3944
R14518 VDD.n3704 VDD.n359 19.3944
R14519 VDD.n3704 VDD.n357 19.3944
R14520 VDD.n3711 VDD.n357 19.3944
R14521 VDD.n3711 VDD.n3710 19.3944
R14522 VDD.n3710 VDD.n346 19.3944
R14523 VDD.n3724 VDD.n346 19.3944
R14524 VDD.n3725 VDD.n3724 19.3944
R14525 VDD.n3726 VDD.n3725 19.3944
R14526 VDD.n3726 VDD.n344 19.3944
R14527 VDD.n3731 VDD.n344 19.3944
R14528 VDD.n3732 VDD.n3731 19.3944
R14529 VDD.n3733 VDD.n3732 19.3944
R14530 VDD.n3733 VDD.n342 19.3944
R14531 VDD.n3738 VDD.n342 19.3944
R14532 VDD.n3739 VDD.n3738 19.3944
R14533 VDD.n3740 VDD.n3739 19.3944
R14534 VDD.n3740 VDD.n340 19.3944
R14535 VDD.n3745 VDD.n340 19.3944
R14536 VDD.n3746 VDD.n3745 19.3944
R14537 VDD.n3747 VDD.n3746 19.3944
R14538 VDD.n3747 VDD.n338 19.3944
R14539 VDD.n3752 VDD.n338 19.3944
R14540 VDD.n3753 VDD.n3752 19.3944
R14541 VDD.n3754 VDD.n3753 19.3944
R14542 VDD.n3754 VDD.n336 19.3944
R14543 VDD.n3759 VDD.n336 19.3944
R14544 VDD.n3760 VDD.n3759 19.3944
R14545 VDD.n3761 VDD.n3760 19.3944
R14546 VDD.n3761 VDD.n334 19.3944
R14547 VDD.n3766 VDD.n334 19.3944
R14548 VDD.n3767 VDD.n3766 19.3944
R14549 VDD.n3768 VDD.n3767 19.3944
R14550 VDD.n3768 VDD.n332 19.3944
R14551 VDD.n3773 VDD.n332 19.3944
R14552 VDD.n3774 VDD.n3773 19.3944
R14553 VDD.n3775 VDD.n3774 19.3944
R14554 VDD.n3775 VDD.n330 19.3944
R14555 VDD.n3780 VDD.n330 19.3944
R14556 VDD.n3781 VDD.n3780 19.3944
R14557 VDD.n3782 VDD.n3781 19.3944
R14558 VDD.n3782 VDD.n328 19.3944
R14559 VDD.n3786 VDD.n328 19.3944
R14560 VDD.n3806 VDD.n307 19.3944
R14561 VDD.n3806 VDD.n313 19.3944
R14562 VDD.n3801 VDD.n313 19.3944
R14563 VDD.n3801 VDD.n3800 19.3944
R14564 VDD.n3800 VDD.n3799 19.3944
R14565 VDD.n3799 VDD.n320 19.3944
R14566 VDD.n3794 VDD.n320 19.3944
R14567 VDD.n3794 VDD.n3793 19.3944
R14568 VDD.n3825 VDD.n3824 19.3944
R14569 VDD.n3824 VDD.n294 19.3944
R14570 VDD.n3819 VDD.n294 19.3944
R14571 VDD.n3819 VDD.n3818 19.3944
R14572 VDD.n3818 VDD.n3817 19.3944
R14573 VDD.n3817 VDD.n301 19.3944
R14574 VDD.n3812 VDD.n301 19.3944
R14575 VDD.n3812 VDD.n3811 19.3944
R14576 VDD.n3843 VDD.n274 19.3944
R14577 VDD.n3843 VDD.n278 19.3944
R14578 VDD.n281 VDD.n278 19.3944
R14579 VDD.n3836 VDD.n281 19.3944
R14580 VDD.n3836 VDD.n3835 19.3944
R14581 VDD.n3835 VDD.n3834 19.3944
R14582 VDD.n3834 VDD.n287 19.3944
R14583 VDD.n3829 VDD.n287 19.3944
R14584 VDD.n3860 VDD.n258 19.3944
R14585 VDD.n3860 VDD.n263 19.3944
R14586 VDD.n3855 VDD.n263 19.3944
R14587 VDD.n3855 VDD.n3854 19.3944
R14588 VDD.n3854 VDD.n3853 19.3944
R14589 VDD.n3853 VDD.n269 19.3944
R14590 VDD.n3848 VDD.n269 19.3944
R14591 VDD.n3878 VDD.n247 19.3944
R14592 VDD.n249 VDD.n247 19.3944
R14593 VDD.n3871 VDD.n249 19.3944
R14594 VDD.n3871 VDD.n3870 19.3944
R14595 VDD.n3870 VDD.n3869 19.3944
R14596 VDD.n3869 VDD.n255 19.3944
R14597 VDD.n3582 VDD.n445 19.3944
R14598 VDD.n3586 VDD.n445 19.3944
R14599 VDD.n3586 VDD.n435 19.3944
R14600 VDD.n3599 VDD.n435 19.3944
R14601 VDD.n3599 VDD.n433 19.3944
R14602 VDD.n3603 VDD.n433 19.3944
R14603 VDD.n3603 VDD.n424 19.3944
R14604 VDD.n3615 VDD.n424 19.3944
R14605 VDD.n3615 VDD.n422 19.3944
R14606 VDD.n3619 VDD.n422 19.3944
R14607 VDD.n3619 VDD.n412 19.3944
R14608 VDD.n3631 VDD.n412 19.3944
R14609 VDD.n3631 VDD.n410 19.3944
R14610 VDD.n3635 VDD.n410 19.3944
R14611 VDD.n3635 VDD.n400 19.3944
R14612 VDD.n3647 VDD.n400 19.3944
R14613 VDD.n3647 VDD.n398 19.3944
R14614 VDD.n3651 VDD.n398 19.3944
R14615 VDD.n3651 VDD.n388 19.3944
R14616 VDD.n3663 VDD.n388 19.3944
R14617 VDD.n3663 VDD.n386 19.3944
R14618 VDD.n3667 VDD.n386 19.3944
R14619 VDD.n3667 VDD.n376 19.3944
R14620 VDD.n3679 VDD.n376 19.3944
R14621 VDD.n3679 VDD.n374 19.3944
R14622 VDD.n3683 VDD.n374 19.3944
R14623 VDD.n3683 VDD.n364 19.3944
R14624 VDD.n3696 VDD.n364 19.3944
R14625 VDD.n3696 VDD.n362 19.3944
R14626 VDD.n3700 VDD.n362 19.3944
R14627 VDD.n3700 VDD.n353 19.3944
R14628 VDD.n3715 VDD.n353 19.3944
R14629 VDD.n3715 VDD.n351 19.3944
R14630 VDD.n3719 VDD.n351 19.3944
R14631 VDD.n3719 VDD.n147 19.3944
R14632 VDD.n3952 VDD.n147 19.3944
R14633 VDD.n3952 VDD.n148 19.3944
R14634 VDD.n3946 VDD.n148 19.3944
R14635 VDD.n3946 VDD.n3945 19.3944
R14636 VDD.n3945 VDD.n3944 19.3944
R14637 VDD.n3944 VDD.n160 19.3944
R14638 VDD.n3938 VDD.n160 19.3944
R14639 VDD.n3938 VDD.n3937 19.3944
R14640 VDD.n3937 VDD.n3936 19.3944
R14641 VDD.n3936 VDD.n171 19.3944
R14642 VDD.n3930 VDD.n171 19.3944
R14643 VDD.n3930 VDD.n3929 19.3944
R14644 VDD.n3929 VDD.n3928 19.3944
R14645 VDD.n3928 VDD.n182 19.3944
R14646 VDD.n3922 VDD.n182 19.3944
R14647 VDD.n3922 VDD.n3921 19.3944
R14648 VDD.n3921 VDD.n3920 19.3944
R14649 VDD.n3920 VDD.n193 19.3944
R14650 VDD.n3914 VDD.n193 19.3944
R14651 VDD.n3914 VDD.n3913 19.3944
R14652 VDD.n3913 VDD.n3912 19.3944
R14653 VDD.n3912 VDD.n204 19.3944
R14654 VDD.n3906 VDD.n204 19.3944
R14655 VDD.n3906 VDD.n3905 19.3944
R14656 VDD.n3905 VDD.n3904 19.3944
R14657 VDD.n3904 VDD.n215 19.3944
R14658 VDD.n3898 VDD.n215 19.3944
R14659 VDD.n3898 VDD.n3897 19.3944
R14660 VDD.n3897 VDD.n3896 19.3944
R14661 VDD.n3896 VDD.n226 19.3944
R14662 VDD.n3890 VDD.n226 19.3944
R14663 VDD.n3890 VDD.n3889 19.3944
R14664 VDD.n3889 VDD.n3888 19.3944
R14665 VDD.n3888 VDD.n237 19.3944
R14666 VDD.n3882 VDD.n237 19.3944
R14667 VDD.n3882 VDD.n3881 19.3944
R14668 VDD.n3481 VDD.n492 19.3944
R14669 VDD.n3481 VDD.n490 19.3944
R14670 VDD.n3487 VDD.n490 19.3944
R14671 VDD.n3487 VDD.n488 19.3944
R14672 VDD.n3491 VDD.n488 19.3944
R14673 VDD.n3491 VDD.n486 19.3944
R14674 VDD.n3497 VDD.n486 19.3944
R14675 VDD.n3501 VDD.n480 19.3944
R14676 VDD.n3507 VDD.n480 19.3944
R14677 VDD.n3507 VDD.n478 19.3944
R14678 VDD.n3511 VDD.n478 19.3944
R14679 VDD.n3511 VDD.n476 19.3944
R14680 VDD.n3517 VDD.n476 19.3944
R14681 VDD.n3517 VDD.n474 19.3944
R14682 VDD.n3524 VDD.n474 19.3944
R14683 VDD.n3530 VDD.n472 19.3944
R14684 VDD.n3530 VDD.n470 19.3944
R14685 VDD.n3534 VDD.n470 19.3944
R14686 VDD.n3534 VDD.n468 19.3944
R14687 VDD.n3540 VDD.n468 19.3944
R14688 VDD.n3540 VDD.n466 19.3944
R14689 VDD.n3544 VDD.n466 19.3944
R14690 VDD.n3544 VDD.n464 19.3944
R14691 VDD.n3463 VDD.n3460 19.3944
R14692 VDD.n3463 VDD.n3459 19.3944
R14693 VDD.n3469 VDD.n3459 19.3944
R14694 VDD.n3472 VDD.n3471 19.3944
R14695 VDD.n3556 VDD.n462 19.3944
R14696 VDD.n3556 VDD.n460 19.3944
R14697 VDD.n3562 VDD.n460 19.3944
R14698 VDD.n3566 VDD.n456 19.3944
R14699 VDD.n454 VDD.n453 19.3944
R14700 VDD.n3573 VDD.n453 19.3944
R14701 VDD.n1466 VDD.n1461 19.2005
R14702 VDD.n2031 VDD.n2028 19.2005
R14703 VDD.n3864 VDD.n258 19.2005
R14704 VDD.n3477 VDD.n492 19.2005
R14705 VDD.n2397 VDD.t182 17.5738
R14706 VDD.n511 VDD.t0 17.5738
R14707 VDD.n1488 VDD.n1308 17.3998
R14708 VDD.n1488 VDD.n1302 17.3998
R14709 VDD.n1496 VDD.n1302 17.3998
R14710 VDD.n1496 VDD.n1296 17.3998
R14711 VDD.n1504 VDD.n1296 17.3998
R14712 VDD.n1512 VDD.n1290 17.3998
R14713 VDD.n1512 VDD.n1284 17.3998
R14714 VDD.n1520 VDD.n1284 17.3998
R14715 VDD.n1520 VDD.n1278 17.3998
R14716 VDD.n1528 VDD.n1278 17.3998
R14717 VDD.n1528 VDD.n1272 17.3998
R14718 VDD.n1536 VDD.n1272 17.3998
R14719 VDD.n1536 VDD.n1266 17.3998
R14720 VDD.n1544 VDD.n1266 17.3998
R14721 VDD.n1544 VDD.n1260 17.3998
R14722 VDD.n1553 VDD.n1260 17.3998
R14723 VDD.n1553 VDD.n1552 17.3998
R14724 VDD.n1561 VDD.n1249 17.3998
R14725 VDD.n1569 VDD.n1249 17.3998
R14726 VDD.n1569 VDD.n1243 17.3998
R14727 VDD.n1577 VDD.n1243 17.3998
R14728 VDD.n1577 VDD.n1237 17.3998
R14729 VDD.n1585 VDD.n1237 17.3998
R14730 VDD.n1585 VDD.n1231 17.3998
R14731 VDD.n1593 VDD.n1231 17.3998
R14732 VDD.n1593 VDD.n1225 17.3998
R14733 VDD.n1601 VDD.n1225 17.3998
R14734 VDD.n1609 VDD.n1219 17.3998
R14735 VDD.n1609 VDD.n1213 17.3998
R14736 VDD.n1617 VDD.n1213 17.3998
R14737 VDD.n1617 VDD.n1207 17.3998
R14738 VDD.n1756 VDD.n1207 17.3998
R14739 VDD.n1756 VDD.n1201 17.3998
R14740 VDD.n1764 VDD.n1201 17.3998
R14741 VDD.n1764 VDD.n1195 17.3998
R14742 VDD.n1772 VDD.n1195 17.3998
R14743 VDD.n1772 VDD.n1189 17.3998
R14744 VDD.n1780 VDD.n1189 17.3998
R14745 VDD.n1788 VDD.n1183 17.3998
R14746 VDD.n1788 VDD.n1177 17.3998
R14747 VDD.n1796 VDD.n1177 17.3998
R14748 VDD.n1796 VDD.n1171 17.3998
R14749 VDD.n1804 VDD.n1171 17.3998
R14750 VDD.n1804 VDD.n1165 17.3998
R14751 VDD.n1812 VDD.n1165 17.3998
R14752 VDD.n1812 VDD.n1158 17.3998
R14753 VDD.n1820 VDD.n1158 17.3998
R14754 VDD.n1820 VDD.n1159 17.3998
R14755 VDD.n1828 VDD.n1147 17.3998
R14756 VDD.n1836 VDD.n1147 17.3998
R14757 VDD.n1836 VDD.n1141 17.3998
R14758 VDD.n1844 VDD.n1141 17.3998
R14759 VDD.n1844 VDD.n1135 17.3998
R14760 VDD.n1852 VDD.n1135 17.3998
R14761 VDD.n1852 VDD.n1129 17.3998
R14762 VDD.n1860 VDD.n1129 17.3998
R14763 VDD.n1860 VDD.n1123 17.3998
R14764 VDD.n1868 VDD.n1123 17.3998
R14765 VDD.n1868 VDD.n1117 17.3998
R14766 VDD.n1876 VDD.n1117 17.3998
R14767 VDD.n1884 VDD.n1111 17.3998
R14768 VDD.n1884 VDD.n1105 17.3998
R14769 VDD.n1892 VDD.n1105 17.3998
R14770 VDD.n1892 VDD.n1096 17.3998
R14771 VDD.n2212 VDD.n1096 17.3998
R14772 VDD.n3580 VDD.n443 17.3998
R14773 VDD.n3588 VDD.n443 17.3998
R14774 VDD.n3588 VDD.n437 17.3998
R14775 VDD.n3597 VDD.n437 17.3998
R14776 VDD.n3597 VDD.n3596 17.3998
R14777 VDD.n3605 VDD.n426 17.3998
R14778 VDD.n3613 VDD.n426 17.3998
R14779 VDD.n3613 VDD.n420 17.3998
R14780 VDD.n3621 VDD.n420 17.3998
R14781 VDD.n3621 VDD.n414 17.3998
R14782 VDD.n3629 VDD.n414 17.3998
R14783 VDD.n3629 VDD.n408 17.3998
R14784 VDD.n3637 VDD.n408 17.3998
R14785 VDD.n3637 VDD.n402 17.3998
R14786 VDD.n3645 VDD.n402 17.3998
R14787 VDD.n3645 VDD.n396 17.3998
R14788 VDD.n3653 VDD.n396 17.3998
R14789 VDD.n3661 VDD.n390 17.3998
R14790 VDD.n3661 VDD.n384 17.3998
R14791 VDD.n3669 VDD.n384 17.3998
R14792 VDD.n3669 VDD.n378 17.3998
R14793 VDD.n3677 VDD.n378 17.3998
R14794 VDD.n3677 VDD.n372 17.3998
R14795 VDD.n3685 VDD.n372 17.3998
R14796 VDD.n3685 VDD.n366 17.3998
R14797 VDD.n3694 VDD.n366 17.3998
R14798 VDD.n3694 VDD.n3693 17.3998
R14799 VDD.n3702 VDD.n355 17.3998
R14800 VDD.n3713 VDD.n355 17.3998
R14801 VDD.n3713 VDD.n349 17.3998
R14802 VDD.n3721 VDD.n349 17.3998
R14803 VDD.n3721 VDD.n151 17.3998
R14804 VDD.n3950 VDD.n151 17.3998
R14805 VDD.n3950 VDD.n3949 17.3998
R14806 VDD.n3949 VDD.n3948 17.3998
R14807 VDD.n3948 VDD.n155 17.3998
R14808 VDD.n3942 VDD.n155 17.3998
R14809 VDD.n3942 VDD.n3941 17.3998
R14810 VDD.n3940 VDD.n165 17.3998
R14811 VDD.n3934 VDD.n165 17.3998
R14812 VDD.n3934 VDD.n3933 17.3998
R14813 VDD.n3933 VDD.n3932 17.3998
R14814 VDD.n3932 VDD.n176 17.3998
R14815 VDD.n3926 VDD.n176 17.3998
R14816 VDD.n3926 VDD.n3925 17.3998
R14817 VDD.n3925 VDD.n3924 17.3998
R14818 VDD.n3924 VDD.n187 17.3998
R14819 VDD.n3918 VDD.n187 17.3998
R14820 VDD.n3917 VDD.n3916 17.3998
R14821 VDD.n3916 VDD.n198 17.3998
R14822 VDD.n3910 VDD.n198 17.3998
R14823 VDD.n3910 VDD.n3909 17.3998
R14824 VDD.n3909 VDD.n3908 17.3998
R14825 VDD.n3908 VDD.n209 17.3998
R14826 VDD.n3902 VDD.n209 17.3998
R14827 VDD.n3902 VDD.n3901 17.3998
R14828 VDD.n3901 VDD.n3900 17.3998
R14829 VDD.n3900 VDD.n220 17.3998
R14830 VDD.n3894 VDD.n220 17.3998
R14831 VDD.n3894 VDD.n3893 17.3998
R14832 VDD.n3892 VDD.n231 17.3998
R14833 VDD.n3886 VDD.n231 17.3998
R14834 VDD.n3886 VDD.n3885 17.3998
R14835 VDD.n3885 VDD.n3884 17.3998
R14836 VDD.n3884 VDD.n242 17.3998
R14837 VDD.n1601 VDD.t127 16.5298
R14838 VDD.t148 VDD.n1183 16.5298
R14839 VDD.n3693 VDD.t143 16.5298
R14840 VDD.t138 VDD.n3940 16.5298
R14841 VDD.n136 VDD.n135 15.8418
R14842 VDD.n123 VDD.n122 15.8418
R14843 VDD.n110 VDD.n109 15.8418
R14844 VDD.n97 VDD.n96 15.8418
R14845 VDD.n84 VDD.n83 15.8418
R14846 VDD.n71 VDD.n70 15.8418
R14847 VDD.n58 VDD.n57 15.8418
R14848 VDD.n45 VDD.n44 15.8418
R14849 VDD.n33 VDD.n32 15.8418
R14850 VDD.n20 VDD.n19 15.8418
R14851 VDD.n1729 VDD.n1728 15.8418
R14852 VDD.n1742 VDD.n1741 15.8418
R14853 VDD.n1703 VDD.n1702 15.8418
R14854 VDD.n1716 VDD.n1715 15.8418
R14855 VDD.n1677 VDD.n1676 15.8418
R14856 VDD.n1690 VDD.n1689 15.8418
R14857 VDD.n1651 VDD.n1650 15.8418
R14858 VDD.n1664 VDD.n1663 15.8418
R14859 VDD.n1626 VDD.n1625 15.8418
R14860 VDD.n1639 VDD.n1638 15.8418
R14861 VDD.n1450 VDD.n1449 15.3217
R14862 VDD.n2015 VDD.n1919 15.3217
R14863 VDD.n3848 VDD.n3847 15.3217
R14864 VDD.n3497 VDD.n484 15.3217
R14865 VDD.n1552 VDD.t129 14.7899
R14866 VDD.n1828 VDD.t131 14.7899
R14867 VDD.n3653 VDD.t135 14.7899
R14868 VDD.t141 VDD.n3917 14.7899
R14869 VDD.n130 VDD.t169 13.2678
R14870 VDD.n130 VDD.t170 13.2678
R14871 VDD.n104 VDD.t144 13.2678
R14872 VDD.n104 VDD.t145 13.2678
R14873 VDD.n78 VDD.t153 13.2678
R14874 VDD.n78 VDD.t147 13.2678
R14875 VDD.n52 VDD.t168 13.2678
R14876 VDD.n52 VDD.t163 13.2678
R14877 VDD.n27 VDD.t146 13.2678
R14878 VDD.n27 VDD.t139 13.2678
R14879 VDD.n1736 VDD.t162 13.2678
R14880 VDD.n1736 VDD.t149 13.2678
R14881 VDD.n1710 VDD.t134 13.2678
R14882 VDD.n1710 VDD.t164 13.2678
R14883 VDD.n1684 VDD.t137 13.2678
R14884 VDD.n1684 VDD.t157 13.2678
R14885 VDD.n1658 VDD.t159 13.2678
R14886 VDD.n1658 VDD.t172 13.2678
R14887 VDD.n1633 VDD.t128 13.2678
R14888 VDD.n1633 VDD.t152 13.2678
R14889 VDD.n1416 VDD.n1412 12.9944
R14890 VDD.n1417 VDD.n1416 12.9944
R14891 VDD.n1977 VDD.n1953 12.9944
R14892 VDD.n1978 VDD.n1977 12.9944
R14893 VDD.n3810 VDD.n307 12.9944
R14894 VDD.n3811 VDD.n3810 12.9944
R14895 VDD.n3552 VDD.n464 12.9944
R14896 VDD.n3552 VDD.n462 12.9944
R14897 VDD.n139 VDD.n134 12.8005
R14898 VDD.n126 VDD.n121 12.8005
R14899 VDD.n113 VDD.n108 12.8005
R14900 VDD.n100 VDD.n95 12.8005
R14901 VDD.n87 VDD.n82 12.8005
R14902 VDD.n74 VDD.n69 12.8005
R14903 VDD.n61 VDD.n56 12.8005
R14904 VDD.n48 VDD.n43 12.8005
R14905 VDD.n36 VDD.n31 12.8005
R14906 VDD.n23 VDD.n18 12.8005
R14907 VDD.n1732 VDD.n1727 12.8005
R14908 VDD.n1745 VDD.n1740 12.8005
R14909 VDD.n1706 VDD.n1701 12.8005
R14910 VDD.n1719 VDD.n1714 12.8005
R14911 VDD.n1680 VDD.n1675 12.8005
R14912 VDD.n1693 VDD.n1688 12.8005
R14913 VDD.n1654 VDD.n1649 12.8005
R14914 VDD.n1667 VDD.n1662 12.8005
R14915 VDD.n1629 VDD.n1624 12.8005
R14916 VDD.n1642 VDD.n1637 12.8005
R14917 VDD.n140 VDD.n132 12.0247
R14918 VDD.n127 VDD.n119 12.0247
R14919 VDD.n114 VDD.n106 12.0247
R14920 VDD.n101 VDD.n93 12.0247
R14921 VDD.n88 VDD.n80 12.0247
R14922 VDD.n75 VDD.n67 12.0247
R14923 VDD.n62 VDD.n54 12.0247
R14924 VDD.n49 VDD.n41 12.0247
R14925 VDD.n37 VDD.n29 12.0247
R14926 VDD.n24 VDD.n16 12.0247
R14927 VDD.n1733 VDD.n1725 12.0247
R14928 VDD.n1746 VDD.n1738 12.0247
R14929 VDD.n1707 VDD.n1699 12.0247
R14930 VDD.n1720 VDD.n1712 12.0247
R14931 VDD.n1681 VDD.n1673 12.0247
R14932 VDD.n1694 VDD.n1686 12.0247
R14933 VDD.n1655 VDD.n1647 12.0247
R14934 VDD.n1668 VDD.n1660 12.0247
R14935 VDD.n1630 VDD.n1622 12.0247
R14936 VDD.n1643 VDD.n1635 12.0247
R14937 VDD.n2397 VDD.n1051 11.832
R14938 VDD.n2403 VDD.n1051 11.832
R14939 VDD.n2403 VDD.n1045 11.832
R14940 VDD.n2409 VDD.n1045 11.832
R14941 VDD.n2409 VDD.n1039 11.832
R14942 VDD.n2415 VDD.n1039 11.832
R14943 VDD.n2421 VDD.n1032 11.832
R14944 VDD.n2421 VDD.n1035 11.832
R14945 VDD.n2427 VDD.n1021 11.832
R14946 VDD.n2433 VDD.n1021 11.832
R14947 VDD.n2433 VDD.n1015 11.832
R14948 VDD.n2439 VDD.n1015 11.832
R14949 VDD.n2439 VDD.n1009 11.832
R14950 VDD.n2445 VDD.n1009 11.832
R14951 VDD.n2445 VDD.n1002 11.832
R14952 VDD.n2451 VDD.n1002 11.832
R14953 VDD.n2451 VDD.n1005 11.832
R14954 VDD.n2463 VDD.n991 11.832
R14955 VDD.n2463 VDD.n985 11.832
R14956 VDD.n2469 VDD.n985 11.832
R14957 VDD.n2469 VDD.n979 11.832
R14958 VDD.n2475 VDD.n979 11.832
R14959 VDD.n2475 VDD.n973 11.832
R14960 VDD.n2481 VDD.n973 11.832
R14961 VDD.n2481 VDD.n967 11.832
R14962 VDD.n2487 VDD.n967 11.832
R14963 VDD.n2493 VDD.n961 11.832
R14964 VDD.n2493 VDD.n955 11.832
R14965 VDD.n2499 VDD.n955 11.832
R14966 VDD.n2499 VDD.n949 11.832
R14967 VDD.n2505 VDD.n949 11.832
R14968 VDD.n2505 VDD.n943 11.832
R14969 VDD.n2511 VDD.n943 11.832
R14970 VDD.n2511 VDD.n936 11.832
R14971 VDD.n2517 VDD.n936 11.832
R14972 VDD.n2517 VDD.n939 11.832
R14973 VDD.n2523 VDD.n925 11.832
R14974 VDD.n2529 VDD.n925 11.832
R14975 VDD.n2529 VDD.n919 11.832
R14976 VDD.n2535 VDD.n919 11.832
R14977 VDD.n2541 VDD.n913 11.832
R14978 VDD.n2541 VDD.n907 11.832
R14979 VDD.n2547 VDD.n907 11.832
R14980 VDD.n2547 VDD.n901 11.832
R14981 VDD.n2553 VDD.n901 11.832
R14982 VDD.n2559 VDD.n895 11.832
R14983 VDD.n2559 VDD.n888 11.832
R14984 VDD.n2565 VDD.n888 11.832
R14985 VDD.n2565 VDD.n891 11.832
R14986 VDD.n2571 VDD.n877 11.832
R14987 VDD.n2577 VDD.n877 11.832
R14988 VDD.n2577 VDD.n871 11.832
R14989 VDD.n2583 VDD.n871 11.832
R14990 VDD.n2589 VDD.n865 11.832
R14991 VDD.n2589 VDD.n859 11.832
R14992 VDD.n2595 VDD.n859 11.832
R14993 VDD.n2595 VDD.n853 11.832
R14994 VDD.n2601 VDD.n853 11.832
R14995 VDD.n2607 VDD.n847 11.832
R14996 VDD.n2607 VDD.n841 11.832
R14997 VDD.n2613 VDD.n841 11.832
R14998 VDD.n2613 VDD.n835 11.832
R14999 VDD.n2619 VDD.n835 11.832
R15000 VDD.n2619 VDD.n829 11.832
R15001 VDD.n2625 VDD.n829 11.832
R15002 VDD.n2636 VDD.n822 11.832
R15003 VDD.n2642 VDD.n816 11.832
R15004 VDD.n2642 VDD.n805 11.832
R15005 VDD.n2696 VDD.n805 11.832
R15006 VDD.n2696 VDD.n775 11.832
R15007 VDD.n3100 VDD.n769 11.832
R15008 VDD.n3106 VDD.n769 11.832
R15009 VDD.n3106 VDD.n763 11.832
R15010 VDD.n3112 VDD.n763 11.832
R15011 VDD.n3118 VDD.n757 11.832
R15012 VDD.n3124 VDD.n751 11.832
R15013 VDD.n3124 VDD.n745 11.832
R15014 VDD.n3130 VDD.n745 11.832
R15015 VDD.n3130 VDD.n739 11.832
R15016 VDD.n3136 VDD.n739 11.832
R15017 VDD.n3136 VDD.n733 11.832
R15018 VDD.n3142 VDD.n733 11.832
R15019 VDD.n3148 VDD.n727 11.832
R15020 VDD.n3148 VDD.n721 11.832
R15021 VDD.n3154 VDD.n721 11.832
R15022 VDD.n3154 VDD.n715 11.832
R15023 VDD.n3160 VDD.n715 11.832
R15024 VDD.n3166 VDD.n709 11.832
R15025 VDD.n3166 VDD.n702 11.832
R15026 VDD.n3172 VDD.n702 11.832
R15027 VDD.n3172 VDD.n705 11.832
R15028 VDD.n3178 VDD.n691 11.832
R15029 VDD.n3184 VDD.n691 11.832
R15030 VDD.n3184 VDD.n685 11.832
R15031 VDD.n3190 VDD.n685 11.832
R15032 VDD.n3196 VDD.n679 11.832
R15033 VDD.n3196 VDD.n673 11.832
R15034 VDD.n3202 VDD.n673 11.832
R15035 VDD.n3202 VDD.n667 11.832
R15036 VDD.n3208 VDD.n667 11.832
R15037 VDD.n3214 VDD.n661 11.832
R15038 VDD.n3214 VDD.n654 11.832
R15039 VDD.n3220 VDD.n654 11.832
R15040 VDD.n3220 VDD.n657 11.832
R15041 VDD.n3226 VDD.n643 11.832
R15042 VDD.n3232 VDD.n643 11.832
R15043 VDD.n3232 VDD.n637 11.832
R15044 VDD.n3238 VDD.n637 11.832
R15045 VDD.n3238 VDD.n631 11.832
R15046 VDD.n3244 VDD.n631 11.832
R15047 VDD.n3244 VDD.n625 11.832
R15048 VDD.n3250 VDD.n625 11.832
R15049 VDD.n3250 VDD.n619 11.832
R15050 VDD.n3256 VDD.n619 11.832
R15051 VDD.n3262 VDD.n613 11.832
R15052 VDD.n3262 VDD.n607 11.832
R15053 VDD.n3268 VDD.n607 11.832
R15054 VDD.n3268 VDD.n601 11.832
R15055 VDD.n3274 VDD.n601 11.832
R15056 VDD.n3274 VDD.n595 11.832
R15057 VDD.n3280 VDD.n595 11.832
R15058 VDD.n3280 VDD.n589 11.832
R15059 VDD.n3286 VDD.n589 11.832
R15060 VDD.n3292 VDD.n578 11.832
R15061 VDD.n3298 VDD.n578 11.832
R15062 VDD.n3298 VDD.n572 11.832
R15063 VDD.n3304 VDD.n572 11.832
R15064 VDD.n3304 VDD.n566 11.832
R15065 VDD.n3310 VDD.n566 11.832
R15066 VDD.n3310 VDD.n559 11.832
R15067 VDD.n3316 VDD.n559 11.832
R15068 VDD.n3316 VDD.n562 11.832
R15069 VDD.n3322 VDD.n547 11.832
R15070 VDD.n3330 VDD.n547 11.832
R15071 VDD.n3336 VDD.n541 11.832
R15072 VDD.n3336 VDD.n517 11.832
R15073 VDD.n3394 VDD.n517 11.832
R15074 VDD.n3394 VDD.n509 11.832
R15075 VDD.n3427 VDD.n509 11.832
R15076 VDD.n3427 VDD.n511 11.832
R15077 VDD.t2 VDD.n847 10.962
R15078 VDD.n3142 VDD.t29 10.962
R15079 VDD.n1449 VDD.n1444 10.6672
R15080 VDD.n2010 VDD.n1919 10.6672
R15081 VDD.n3847 VDD.n274 10.6672
R15082 VDD.n3501 VDD.n484 10.6672
R15083 VDD.n2395 VDD.n1049 10.6151
R15084 VDD.n2405 VDD.n1049 10.6151
R15085 VDD.n2406 VDD.n2405 10.6151
R15086 VDD.n2407 VDD.n2406 10.6151
R15087 VDD.n2407 VDD.n1037 10.6151
R15088 VDD.n2417 VDD.n1037 10.6151
R15089 VDD.n2418 VDD.n2417 10.6151
R15090 VDD.n2419 VDD.n2418 10.6151
R15091 VDD.n2419 VDD.n1025 10.6151
R15092 VDD.n2429 VDD.n1025 10.6151
R15093 VDD.n2430 VDD.n2429 10.6151
R15094 VDD.n2431 VDD.n2430 10.6151
R15095 VDD.n2431 VDD.n1013 10.6151
R15096 VDD.n2441 VDD.n1013 10.6151
R15097 VDD.n2442 VDD.n2441 10.6151
R15098 VDD.n2443 VDD.n2442 10.6151
R15099 VDD.n2443 VDD.n1000 10.6151
R15100 VDD.n2453 VDD.n1000 10.6151
R15101 VDD.n2454 VDD.n2453 10.6151
R15102 VDD.n2455 VDD.n2454 10.6151
R15103 VDD.n2455 VDD.n989 10.6151
R15104 VDD.n2465 VDD.n989 10.6151
R15105 VDD.n2466 VDD.n2465 10.6151
R15106 VDD.n2467 VDD.n2466 10.6151
R15107 VDD.n2467 VDD.n977 10.6151
R15108 VDD.n2477 VDD.n977 10.6151
R15109 VDD.n2478 VDD.n2477 10.6151
R15110 VDD.n2479 VDD.n2478 10.6151
R15111 VDD.n2479 VDD.n965 10.6151
R15112 VDD.n2489 VDD.n965 10.6151
R15113 VDD.n2490 VDD.n2489 10.6151
R15114 VDD.n2491 VDD.n2490 10.6151
R15115 VDD.n2491 VDD.n953 10.6151
R15116 VDD.n2501 VDD.n953 10.6151
R15117 VDD.n2502 VDD.n2501 10.6151
R15118 VDD.n2503 VDD.n2502 10.6151
R15119 VDD.n2503 VDD.n941 10.6151
R15120 VDD.n2513 VDD.n941 10.6151
R15121 VDD.n2514 VDD.n2513 10.6151
R15122 VDD.n2515 VDD.n2514 10.6151
R15123 VDD.n2515 VDD.n929 10.6151
R15124 VDD.n2525 VDD.n929 10.6151
R15125 VDD.n2526 VDD.n2525 10.6151
R15126 VDD.n2527 VDD.n2526 10.6151
R15127 VDD.n2527 VDD.n917 10.6151
R15128 VDD.n2537 VDD.n917 10.6151
R15129 VDD.n2538 VDD.n2537 10.6151
R15130 VDD.n2539 VDD.n2538 10.6151
R15131 VDD.n2539 VDD.n905 10.6151
R15132 VDD.n2549 VDD.n905 10.6151
R15133 VDD.n2550 VDD.n2549 10.6151
R15134 VDD.n2551 VDD.n2550 10.6151
R15135 VDD.n2551 VDD.n893 10.6151
R15136 VDD.n2561 VDD.n893 10.6151
R15137 VDD.n2562 VDD.n2561 10.6151
R15138 VDD.n2563 VDD.n2562 10.6151
R15139 VDD.n2563 VDD.n881 10.6151
R15140 VDD.n2573 VDD.n881 10.6151
R15141 VDD.n2574 VDD.n2573 10.6151
R15142 VDD.n2575 VDD.n2574 10.6151
R15143 VDD.n2575 VDD.n869 10.6151
R15144 VDD.n2585 VDD.n869 10.6151
R15145 VDD.n2586 VDD.n2585 10.6151
R15146 VDD.n2587 VDD.n2586 10.6151
R15147 VDD.n2587 VDD.n857 10.6151
R15148 VDD.n2597 VDD.n857 10.6151
R15149 VDD.n2598 VDD.n2597 10.6151
R15150 VDD.n2599 VDD.n2598 10.6151
R15151 VDD.n2599 VDD.n845 10.6151
R15152 VDD.n2609 VDD.n845 10.6151
R15153 VDD.n2610 VDD.n2609 10.6151
R15154 VDD.n2611 VDD.n2610 10.6151
R15155 VDD.n2611 VDD.n833 10.6151
R15156 VDD.n2621 VDD.n833 10.6151
R15157 VDD.n2622 VDD.n2621 10.6151
R15158 VDD.n2623 VDD.n2622 10.6151
R15159 VDD.n2623 VDD.n820 10.6151
R15160 VDD.n2638 VDD.n820 10.6151
R15161 VDD.n2639 VDD.n2638 10.6151
R15162 VDD.n2640 VDD.n2639 10.6151
R15163 VDD.n2640 VDD.n810 10.6151
R15164 VDD.n2694 VDD.n810 10.6151
R15165 VDD.n2694 VDD.n2693 10.6151
R15166 VDD.n2692 VDD.n2690 10.6151
R15167 VDD.n2690 VDD.n2687 10.6151
R15168 VDD.n2687 VDD.n2686 10.6151
R15169 VDD.n2686 VDD.n2683 10.6151
R15170 VDD.n2683 VDD.n2682 10.6151
R15171 VDD.n2682 VDD.n2679 10.6151
R15172 VDD.n2679 VDD.n2678 10.6151
R15173 VDD.n2678 VDD.n2675 10.6151
R15174 VDD.n2675 VDD.n2674 10.6151
R15175 VDD.n2674 VDD.n2671 10.6151
R15176 VDD.n2671 VDD.n2670 10.6151
R15177 VDD.n2670 VDD.n2667 10.6151
R15178 VDD.n2667 VDD.n2666 10.6151
R15179 VDD.n2666 VDD.n2663 10.6151
R15180 VDD.n2663 VDD.n2662 10.6151
R15181 VDD.n2662 VDD.n2659 10.6151
R15182 VDD.n2659 VDD.n2658 10.6151
R15183 VDD.n2658 VDD.n2655 10.6151
R15184 VDD.n2655 VDD.n2654 10.6151
R15185 VDD.n2651 VDD.n2650 10.6151
R15186 VDD.n2173 VDD.n2172 10.6151
R15187 VDD.n2172 VDD.n2170 10.6151
R15188 VDD.n2170 VDD.n2169 10.6151
R15189 VDD.n2169 VDD.n2167 10.6151
R15190 VDD.n2167 VDD.n2166 10.6151
R15191 VDD.n2166 VDD.n2164 10.6151
R15192 VDD.n2164 VDD.n2163 10.6151
R15193 VDD.n2163 VDD.n2161 10.6151
R15194 VDD.n2161 VDD.n2160 10.6151
R15195 VDD.n2160 VDD.n2158 10.6151
R15196 VDD.n2158 VDD.n2157 10.6151
R15197 VDD.n2157 VDD.n2155 10.6151
R15198 VDD.n2155 VDD.n2154 10.6151
R15199 VDD.n2154 VDD.n2152 10.6151
R15200 VDD.n2152 VDD.n2151 10.6151
R15201 VDD.n2151 VDD.n2149 10.6151
R15202 VDD.n2149 VDD.n2148 10.6151
R15203 VDD.n2148 VDD.n2146 10.6151
R15204 VDD.n2146 VDD.n2145 10.6151
R15205 VDD.n2145 VDD.n2143 10.6151
R15206 VDD.n2143 VDD.n2142 10.6151
R15207 VDD.n2142 VDD.n2140 10.6151
R15208 VDD.n2140 VDD.n2139 10.6151
R15209 VDD.n2139 VDD.n2137 10.6151
R15210 VDD.n2137 VDD.n2136 10.6151
R15211 VDD.n2136 VDD.n2134 10.6151
R15212 VDD.n2134 VDD.n2133 10.6151
R15213 VDD.n2133 VDD.n2131 10.6151
R15214 VDD.n2131 VDD.n2130 10.6151
R15215 VDD.n2130 VDD.n2128 10.6151
R15216 VDD.n2128 VDD.n2127 10.6151
R15217 VDD.n2127 VDD.n2125 10.6151
R15218 VDD.n2125 VDD.n2124 10.6151
R15219 VDD.n2124 VDD.n2122 10.6151
R15220 VDD.n2122 VDD.n2121 10.6151
R15221 VDD.n2121 VDD.n2119 10.6151
R15222 VDD.n2119 VDD.n2118 10.6151
R15223 VDD.n2118 VDD.n2116 10.6151
R15224 VDD.n2116 VDD.n2115 10.6151
R15225 VDD.n2115 VDD.n2113 10.6151
R15226 VDD.n2113 VDD.n2112 10.6151
R15227 VDD.n2112 VDD.n2110 10.6151
R15228 VDD.n2110 VDD.n2109 10.6151
R15229 VDD.n2109 VDD.n2107 10.6151
R15230 VDD.n2107 VDD.n2106 10.6151
R15231 VDD.n2106 VDD.n2104 10.6151
R15232 VDD.n2104 VDD.n2103 10.6151
R15233 VDD.n2103 VDD.n2101 10.6151
R15234 VDD.n2101 VDD.n2100 10.6151
R15235 VDD.n2100 VDD.n2098 10.6151
R15236 VDD.n2098 VDD.n2097 10.6151
R15237 VDD.n2097 VDD.n2095 10.6151
R15238 VDD.n2095 VDD.n2094 10.6151
R15239 VDD.n2094 VDD.n2092 10.6151
R15240 VDD.n2092 VDD.n2091 10.6151
R15241 VDD.n2091 VDD.n2089 10.6151
R15242 VDD.n2089 VDD.n2088 10.6151
R15243 VDD.n2088 VDD.n2086 10.6151
R15244 VDD.n2086 VDD.n2085 10.6151
R15245 VDD.n2085 VDD.n2083 10.6151
R15246 VDD.n2083 VDD.n2082 10.6151
R15247 VDD.n2082 VDD.n2080 10.6151
R15248 VDD.n2080 VDD.n2079 10.6151
R15249 VDD.n2079 VDD.n2077 10.6151
R15250 VDD.n2077 VDD.n2076 10.6151
R15251 VDD.n2076 VDD.n2074 10.6151
R15252 VDD.n2074 VDD.n2073 10.6151
R15253 VDD.n2073 VDD.n2071 10.6151
R15254 VDD.n2071 VDD.n2070 10.6151
R15255 VDD.n2070 VDD.n2068 10.6151
R15256 VDD.n2068 VDD.n2067 10.6151
R15257 VDD.n2067 VDD.n2065 10.6151
R15258 VDD.n2065 VDD.n2064 10.6151
R15259 VDD.n2064 VDD.n2062 10.6151
R15260 VDD.n2062 VDD.n2061 10.6151
R15261 VDD.n2061 VDD.n2059 10.6151
R15262 VDD.n2059 VDD.n2058 10.6151
R15263 VDD.n2058 VDD.n2056 10.6151
R15264 VDD.n2056 VDD.n2055 10.6151
R15265 VDD.n2055 VDD.n814 10.6151
R15266 VDD.n2645 VDD.n814 10.6151
R15267 VDD.n2646 VDD.n2645 10.6151
R15268 VDD.n2647 VDD.n2646 10.6151
R15269 VDD.n2394 VDD.n2393 10.6151
R15270 VDD.n2393 VDD.n1060 10.6151
R15271 VDD.n2039 VDD.n1060 10.6151
R15272 VDD.n2040 VDD.n2039 10.6151
R15273 VDD.n2043 VDD.n2040 10.6151
R15274 VDD.n2044 VDD.n2043 10.6151
R15275 VDD.n2047 VDD.n2044 10.6151
R15276 VDD.n2048 VDD.n2047 10.6151
R15277 VDD.n2051 VDD.n2048 10.6151
R15278 VDD.n2052 VDD.n2051 10.6151
R15279 VDD.n2196 VDD.n2193 10.6151
R15280 VDD.n2193 VDD.n2190 10.6151
R15281 VDD.n2190 VDD.n2189 10.6151
R15282 VDD.n2189 VDD.n2186 10.6151
R15283 VDD.n2186 VDD.n2185 10.6151
R15284 VDD.n2185 VDD.n2182 10.6151
R15285 VDD.n2182 VDD.n2181 10.6151
R15286 VDD.n2181 VDD.n2178 10.6151
R15287 VDD.n2176 VDD.n2174 10.6151
R15288 VDD.n2837 VDD.n2835 10.6151
R15289 VDD.n2838 VDD.n2837 10.6151
R15290 VDD.n2840 VDD.n2838 10.6151
R15291 VDD.n2841 VDD.n2840 10.6151
R15292 VDD.n2843 VDD.n2841 10.6151
R15293 VDD.n2844 VDD.n2843 10.6151
R15294 VDD.n2846 VDD.n2844 10.6151
R15295 VDD.n2847 VDD.n2846 10.6151
R15296 VDD.n2849 VDD.n2847 10.6151
R15297 VDD.n2850 VDD.n2849 10.6151
R15298 VDD.n2852 VDD.n2850 10.6151
R15299 VDD.n2853 VDD.n2852 10.6151
R15300 VDD.n2855 VDD.n2853 10.6151
R15301 VDD.n2856 VDD.n2855 10.6151
R15302 VDD.n2858 VDD.n2856 10.6151
R15303 VDD.n2859 VDD.n2858 10.6151
R15304 VDD.n2861 VDD.n2859 10.6151
R15305 VDD.n2862 VDD.n2861 10.6151
R15306 VDD.n2864 VDD.n2862 10.6151
R15307 VDD.n2865 VDD.n2864 10.6151
R15308 VDD.n2867 VDD.n2865 10.6151
R15309 VDD.n2868 VDD.n2867 10.6151
R15310 VDD.n2870 VDD.n2868 10.6151
R15311 VDD.n2871 VDD.n2870 10.6151
R15312 VDD.n2873 VDD.n2871 10.6151
R15313 VDD.n2874 VDD.n2873 10.6151
R15314 VDD.n2876 VDD.n2874 10.6151
R15315 VDD.n2877 VDD.n2876 10.6151
R15316 VDD.n2879 VDD.n2877 10.6151
R15317 VDD.n2880 VDD.n2879 10.6151
R15318 VDD.n2882 VDD.n2880 10.6151
R15319 VDD.n2883 VDD.n2882 10.6151
R15320 VDD.n2885 VDD.n2883 10.6151
R15321 VDD.n2886 VDD.n2885 10.6151
R15322 VDD.n2888 VDD.n2886 10.6151
R15323 VDD.n2889 VDD.n2888 10.6151
R15324 VDD.n2891 VDD.n2889 10.6151
R15325 VDD.n2892 VDD.n2891 10.6151
R15326 VDD.n2894 VDD.n2892 10.6151
R15327 VDD.n2895 VDD.n2894 10.6151
R15328 VDD.n2897 VDD.n2895 10.6151
R15329 VDD.n2898 VDD.n2897 10.6151
R15330 VDD.n2900 VDD.n2898 10.6151
R15331 VDD.n2901 VDD.n2900 10.6151
R15332 VDD.n2903 VDD.n2901 10.6151
R15333 VDD.n2904 VDD.n2903 10.6151
R15334 VDD.n2906 VDD.n2904 10.6151
R15335 VDD.n2907 VDD.n2906 10.6151
R15336 VDD.n2909 VDD.n2907 10.6151
R15337 VDD.n2910 VDD.n2909 10.6151
R15338 VDD.n2912 VDD.n2910 10.6151
R15339 VDD.n2913 VDD.n2912 10.6151
R15340 VDD.n2915 VDD.n2913 10.6151
R15341 VDD.n2916 VDD.n2915 10.6151
R15342 VDD.n2918 VDD.n2916 10.6151
R15343 VDD.n2919 VDD.n2918 10.6151
R15344 VDD.n2921 VDD.n2919 10.6151
R15345 VDD.n2922 VDD.n2921 10.6151
R15346 VDD.n2924 VDD.n2922 10.6151
R15347 VDD.n2925 VDD.n2924 10.6151
R15348 VDD.n2927 VDD.n2925 10.6151
R15349 VDD.n2928 VDD.n2927 10.6151
R15350 VDD.n2954 VDD.n2928 10.6151
R15351 VDD.n2954 VDD.n2953 10.6151
R15352 VDD.n2953 VDD.n2952 10.6151
R15353 VDD.n2952 VDD.n2950 10.6151
R15354 VDD.n2950 VDD.n2949 10.6151
R15355 VDD.n2949 VDD.n2947 10.6151
R15356 VDD.n2947 VDD.n2946 10.6151
R15357 VDD.n2946 VDD.n2944 10.6151
R15358 VDD.n2944 VDD.n2943 10.6151
R15359 VDD.n2943 VDD.n2941 10.6151
R15360 VDD.n2941 VDD.n2940 10.6151
R15361 VDD.n2940 VDD.n2938 10.6151
R15362 VDD.n2938 VDD.n2937 10.6151
R15363 VDD.n2937 VDD.n2935 10.6151
R15364 VDD.n2935 VDD.n2934 10.6151
R15365 VDD.n2934 VDD.n2932 10.6151
R15366 VDD.n2932 VDD.n2931 10.6151
R15367 VDD.n2931 VDD.n2929 10.6151
R15368 VDD.n2929 VDD.n507 10.6151
R15369 VDD.n3429 VDD.n507 10.6151
R15370 VDD.n3430 VDD.n3429 10.6151
R15371 VDD.n2792 VDD.n773 10.6151
R15372 VDD.n2793 VDD.n2792 10.6151
R15373 VDD.n2794 VDD.n2793 10.6151
R15374 VDD.n2794 VDD.n2788 10.6151
R15375 VDD.n2800 VDD.n2788 10.6151
R15376 VDD.n2801 VDD.n2800 10.6151
R15377 VDD.n2802 VDD.n2801 10.6151
R15378 VDD.n2802 VDD.n2786 10.6151
R15379 VDD.n2808 VDD.n2786 10.6151
R15380 VDD.n2809 VDD.n2808 10.6151
R15381 VDD.n2810 VDD.n2809 10.6151
R15382 VDD.n2810 VDD.n2784 10.6151
R15383 VDD.n2816 VDD.n2784 10.6151
R15384 VDD.n2817 VDD.n2816 10.6151
R15385 VDD.n2818 VDD.n2817 10.6151
R15386 VDD.n2818 VDD.n2782 10.6151
R15387 VDD.n2824 VDD.n2782 10.6151
R15388 VDD.n2825 VDD.n2824 10.6151
R15389 VDD.n2829 VDD.n2825 10.6151
R15390 VDD.n2834 VDD.n2780 10.6151
R15391 VDD.n3103 VDD.n3102 10.6151
R15392 VDD.n3104 VDD.n3103 10.6151
R15393 VDD.n3104 VDD.n761 10.6151
R15394 VDD.n3114 VDD.n761 10.6151
R15395 VDD.n3115 VDD.n3114 10.6151
R15396 VDD.n3116 VDD.n3115 10.6151
R15397 VDD.n3116 VDD.n749 10.6151
R15398 VDD.n3126 VDD.n749 10.6151
R15399 VDD.n3127 VDD.n3126 10.6151
R15400 VDD.n3128 VDD.n3127 10.6151
R15401 VDD.n3128 VDD.n737 10.6151
R15402 VDD.n3138 VDD.n737 10.6151
R15403 VDD.n3139 VDD.n3138 10.6151
R15404 VDD.n3140 VDD.n3139 10.6151
R15405 VDD.n3140 VDD.n725 10.6151
R15406 VDD.n3150 VDD.n725 10.6151
R15407 VDD.n3151 VDD.n3150 10.6151
R15408 VDD.n3152 VDD.n3151 10.6151
R15409 VDD.n3152 VDD.n713 10.6151
R15410 VDD.n3162 VDD.n713 10.6151
R15411 VDD.n3163 VDD.n3162 10.6151
R15412 VDD.n3164 VDD.n3163 10.6151
R15413 VDD.n3164 VDD.n700 10.6151
R15414 VDD.n3174 VDD.n700 10.6151
R15415 VDD.n3175 VDD.n3174 10.6151
R15416 VDD.n3176 VDD.n3175 10.6151
R15417 VDD.n3176 VDD.n689 10.6151
R15418 VDD.n3186 VDD.n689 10.6151
R15419 VDD.n3187 VDD.n3186 10.6151
R15420 VDD.n3188 VDD.n3187 10.6151
R15421 VDD.n3188 VDD.n677 10.6151
R15422 VDD.n3198 VDD.n677 10.6151
R15423 VDD.n3199 VDD.n3198 10.6151
R15424 VDD.n3200 VDD.n3199 10.6151
R15425 VDD.n3200 VDD.n665 10.6151
R15426 VDD.n3210 VDD.n665 10.6151
R15427 VDD.n3211 VDD.n3210 10.6151
R15428 VDD.n3212 VDD.n3211 10.6151
R15429 VDD.n3212 VDD.n652 10.6151
R15430 VDD.n3222 VDD.n652 10.6151
R15431 VDD.n3223 VDD.n3222 10.6151
R15432 VDD.n3224 VDD.n3223 10.6151
R15433 VDD.n3224 VDD.n641 10.6151
R15434 VDD.n3234 VDD.n641 10.6151
R15435 VDD.n3235 VDD.n3234 10.6151
R15436 VDD.n3236 VDD.n3235 10.6151
R15437 VDD.n3236 VDD.n629 10.6151
R15438 VDD.n3246 VDD.n629 10.6151
R15439 VDD.n3247 VDD.n3246 10.6151
R15440 VDD.n3248 VDD.n3247 10.6151
R15441 VDD.n3248 VDD.n617 10.6151
R15442 VDD.n3258 VDD.n617 10.6151
R15443 VDD.n3259 VDD.n3258 10.6151
R15444 VDD.n3260 VDD.n3259 10.6151
R15445 VDD.n3260 VDD.n605 10.6151
R15446 VDD.n3270 VDD.n605 10.6151
R15447 VDD.n3271 VDD.n3270 10.6151
R15448 VDD.n3272 VDD.n3271 10.6151
R15449 VDD.n3272 VDD.n593 10.6151
R15450 VDD.n3282 VDD.n593 10.6151
R15451 VDD.n3283 VDD.n3282 10.6151
R15452 VDD.n3284 VDD.n3283 10.6151
R15453 VDD.n3284 VDD.n582 10.6151
R15454 VDD.n3294 VDD.n582 10.6151
R15455 VDD.n3295 VDD.n3294 10.6151
R15456 VDD.n3296 VDD.n3295 10.6151
R15457 VDD.n3296 VDD.n570 10.6151
R15458 VDD.n3306 VDD.n570 10.6151
R15459 VDD.n3307 VDD.n3306 10.6151
R15460 VDD.n3308 VDD.n3307 10.6151
R15461 VDD.n3308 VDD.n557 10.6151
R15462 VDD.n3318 VDD.n557 10.6151
R15463 VDD.n3319 VDD.n3318 10.6151
R15464 VDD.n3320 VDD.n3319 10.6151
R15465 VDD.n3320 VDD.n545 10.6151
R15466 VDD.n3332 VDD.n545 10.6151
R15467 VDD.n3333 VDD.n3332 10.6151
R15468 VDD.n3334 VDD.n3333 10.6151
R15469 VDD.n3334 VDD.n515 10.6151
R15470 VDD.n3396 VDD.n515 10.6151
R15471 VDD.n3397 VDD.n3396 10.6151
R15472 VDD.n3425 VDD.n3397 10.6151
R15473 VDD.n3425 VDD.n3424 10.6151
R15474 VDD.n3423 VDD.n3398 10.6151
R15475 VDD.n3399 VDD.n3398 10.6151
R15476 VDD.n3416 VDD.n3399 10.6151
R15477 VDD.n3416 VDD.n3415 10.6151
R15478 VDD.n3415 VDD.n3414 10.6151
R15479 VDD.n3414 VDD.n3401 10.6151
R15480 VDD.n3409 VDD.n3401 10.6151
R15481 VDD.n3409 VDD.n3408 10.6151
R15482 VDD.n3408 VDD.n3407 10.6151
R15483 VDD.n3407 VDD.n493 10.6151
R15484 VDD.n3450 VDD.n494 10.6151
R15485 VDD.n3445 VDD.n494 10.6151
R15486 VDD.n3445 VDD.n3444 10.6151
R15487 VDD.n3444 VDD.n3443 10.6151
R15488 VDD.n3443 VDD.n498 10.6151
R15489 VDD.n3438 VDD.n498 10.6151
R15490 VDD.n3438 VDD.n3437 10.6151
R15491 VDD.n3437 VDD.n3436 10.6151
R15492 VDD.n3431 VDD.n505 10.6151
R15493 VDD.n3384 VDD.n523 10.6151
R15494 VDD.n3384 VDD.n3383 10.6151
R15495 VDD.n3383 VDD.n3382 10.6151
R15496 VDD.n3382 VDD.n525 10.6151
R15497 VDD.n3377 VDD.n525 10.6151
R15498 VDD.n3377 VDD.n3376 10.6151
R15499 VDD.n3376 VDD.n3375 10.6151
R15500 VDD.n3375 VDD.n528 10.6151
R15501 VDD.n3370 VDD.n528 10.6151
R15502 VDD.n3370 VDD.n3369 10.6151
R15503 VDD.n3365 VDD.n3364 10.6151
R15504 VDD.n3364 VDD.n3363 10.6151
R15505 VDD.n3363 VDD.n531 10.6151
R15506 VDD.n3358 VDD.n531 10.6151
R15507 VDD.n3358 VDD.n3357 10.6151
R15508 VDD.n3357 VDD.n3356 10.6151
R15509 VDD.n3356 VDD.n534 10.6151
R15510 VDD.n3351 VDD.n534 10.6151
R15511 VDD.n3349 VDD.n3348 10.6151
R15512 VDD.n3052 VDD.n3051 10.6151
R15513 VDD.n3051 VDD.n3049 10.6151
R15514 VDD.n3049 VDD.n3048 10.6151
R15515 VDD.n3048 VDD.n3046 10.6151
R15516 VDD.n3046 VDD.n3045 10.6151
R15517 VDD.n3045 VDD.n3043 10.6151
R15518 VDD.n3043 VDD.n3042 10.6151
R15519 VDD.n3042 VDD.n3040 10.6151
R15520 VDD.n3040 VDD.n3039 10.6151
R15521 VDD.n3039 VDD.n3037 10.6151
R15522 VDD.n3037 VDD.n3036 10.6151
R15523 VDD.n3036 VDD.n3034 10.6151
R15524 VDD.n3034 VDD.n3033 10.6151
R15525 VDD.n3033 VDD.n3031 10.6151
R15526 VDD.n3031 VDD.n3030 10.6151
R15527 VDD.n3030 VDD.n3028 10.6151
R15528 VDD.n3028 VDD.n3027 10.6151
R15529 VDD.n3027 VDD.n3025 10.6151
R15530 VDD.n3025 VDD.n3024 10.6151
R15531 VDD.n3024 VDD.n3022 10.6151
R15532 VDD.n3022 VDD.n3021 10.6151
R15533 VDD.n3021 VDD.n3019 10.6151
R15534 VDD.n3019 VDD.n3018 10.6151
R15535 VDD.n3018 VDD.n3016 10.6151
R15536 VDD.n3016 VDD.n3015 10.6151
R15537 VDD.n3015 VDD.n3013 10.6151
R15538 VDD.n3013 VDD.n3012 10.6151
R15539 VDD.n3012 VDD.n3010 10.6151
R15540 VDD.n3010 VDD.n3009 10.6151
R15541 VDD.n3009 VDD.n3007 10.6151
R15542 VDD.n3007 VDD.n3006 10.6151
R15543 VDD.n3006 VDD.n3004 10.6151
R15544 VDD.n3004 VDD.n3003 10.6151
R15545 VDD.n3003 VDD.n3001 10.6151
R15546 VDD.n3001 VDD.n3000 10.6151
R15547 VDD.n3000 VDD.n2998 10.6151
R15548 VDD.n2998 VDD.n2997 10.6151
R15549 VDD.n2997 VDD.n2995 10.6151
R15550 VDD.n2995 VDD.n2994 10.6151
R15551 VDD.n2994 VDD.n2992 10.6151
R15552 VDD.n2992 VDD.n2991 10.6151
R15553 VDD.n2991 VDD.n2989 10.6151
R15554 VDD.n2989 VDD.n2988 10.6151
R15555 VDD.n2988 VDD.n2986 10.6151
R15556 VDD.n2986 VDD.n2985 10.6151
R15557 VDD.n2985 VDD.n2983 10.6151
R15558 VDD.n2983 VDD.n2982 10.6151
R15559 VDD.n2982 VDD.n2980 10.6151
R15560 VDD.n2980 VDD.n2979 10.6151
R15561 VDD.n2979 VDD.n2977 10.6151
R15562 VDD.n2977 VDD.n2976 10.6151
R15563 VDD.n2976 VDD.n2974 10.6151
R15564 VDD.n2974 VDD.n2973 10.6151
R15565 VDD.n2973 VDD.n2971 10.6151
R15566 VDD.n2971 VDD.n2970 10.6151
R15567 VDD.n2970 VDD.n2968 10.6151
R15568 VDD.n2968 VDD.n2967 10.6151
R15569 VDD.n2967 VDD.n2965 10.6151
R15570 VDD.n2965 VDD.n2964 10.6151
R15571 VDD.n2964 VDD.n2962 10.6151
R15572 VDD.n2962 VDD.n2961 10.6151
R15573 VDD.n2961 VDD.n2959 10.6151
R15574 VDD.n2959 VDD.n2958 10.6151
R15575 VDD.n2958 VDD.n2779 10.6151
R15576 VDD.n2779 VDD.n2778 10.6151
R15577 VDD.n2778 VDD.n2776 10.6151
R15578 VDD.n2776 VDD.n2775 10.6151
R15579 VDD.n2775 VDD.n2773 10.6151
R15580 VDD.n2773 VDD.n2772 10.6151
R15581 VDD.n2772 VDD.n2770 10.6151
R15582 VDD.n2770 VDD.n2769 10.6151
R15583 VDD.n2769 VDD.n2767 10.6151
R15584 VDD.n2767 VDD.n2766 10.6151
R15585 VDD.n2766 VDD.n2764 10.6151
R15586 VDD.n2764 VDD.n2763 10.6151
R15587 VDD.n2763 VDD.n2761 10.6151
R15588 VDD.n2761 VDD.n2760 10.6151
R15589 VDD.n2760 VDD.n539 10.6151
R15590 VDD.n3339 VDD.n539 10.6151
R15591 VDD.n3340 VDD.n3339 10.6151
R15592 VDD.n3342 VDD.n3340 10.6151
R15593 VDD.n3343 VDD.n3342 10.6151
R15594 VDD.n3344 VDD.n3343 10.6151
R15595 VDD.n3097 VDD.n3096 10.6151
R15596 VDD.n3096 VDD.n2748 10.6151
R15597 VDD.n3090 VDD.n2748 10.6151
R15598 VDD.n3090 VDD.n3089 10.6151
R15599 VDD.n3089 VDD.n3088 10.6151
R15600 VDD.n3088 VDD.n2750 10.6151
R15601 VDD.n3082 VDD.n2750 10.6151
R15602 VDD.n3082 VDD.n3081 10.6151
R15603 VDD.n3081 VDD.n3080 10.6151
R15604 VDD.n3080 VDD.n2752 10.6151
R15605 VDD.n3074 VDD.n2752 10.6151
R15606 VDD.n3074 VDD.n3073 10.6151
R15607 VDD.n3073 VDD.n3072 10.6151
R15608 VDD.n3072 VDD.n2754 10.6151
R15609 VDD.n3066 VDD.n2754 10.6151
R15610 VDD.n3066 VDD.n3065 10.6151
R15611 VDD.n3065 VDD.n3064 10.6151
R15612 VDD.n3064 VDD.n2756 10.6151
R15613 VDD.n3058 VDD.n2756 10.6151
R15614 VDD.n3056 VDD.n3055 10.6151
R15615 VDD.n3098 VDD.n767 10.6151
R15616 VDD.n3108 VDD.n767 10.6151
R15617 VDD.n3109 VDD.n3108 10.6151
R15618 VDD.n3110 VDD.n3109 10.6151
R15619 VDD.n3110 VDD.n755 10.6151
R15620 VDD.n3120 VDD.n755 10.6151
R15621 VDD.n3121 VDD.n3120 10.6151
R15622 VDD.n3122 VDD.n3121 10.6151
R15623 VDD.n3122 VDD.n743 10.6151
R15624 VDD.n3132 VDD.n743 10.6151
R15625 VDD.n3133 VDD.n3132 10.6151
R15626 VDD.n3134 VDD.n3133 10.6151
R15627 VDD.n3134 VDD.n731 10.6151
R15628 VDD.n3144 VDD.n731 10.6151
R15629 VDD.n3145 VDD.n3144 10.6151
R15630 VDD.n3146 VDD.n3145 10.6151
R15631 VDD.n3146 VDD.n719 10.6151
R15632 VDD.n3156 VDD.n719 10.6151
R15633 VDD.n3157 VDD.n3156 10.6151
R15634 VDD.n3158 VDD.n3157 10.6151
R15635 VDD.n3158 VDD.n707 10.6151
R15636 VDD.n3168 VDD.n707 10.6151
R15637 VDD.n3169 VDD.n3168 10.6151
R15638 VDD.n3170 VDD.n3169 10.6151
R15639 VDD.n3170 VDD.n695 10.6151
R15640 VDD.n3180 VDD.n695 10.6151
R15641 VDD.n3181 VDD.n3180 10.6151
R15642 VDD.n3182 VDD.n3181 10.6151
R15643 VDD.n3182 VDD.n683 10.6151
R15644 VDD.n3192 VDD.n683 10.6151
R15645 VDD.n3193 VDD.n3192 10.6151
R15646 VDD.n3194 VDD.n3193 10.6151
R15647 VDD.n3194 VDD.n671 10.6151
R15648 VDD.n3204 VDD.n671 10.6151
R15649 VDD.n3205 VDD.n3204 10.6151
R15650 VDD.n3206 VDD.n3205 10.6151
R15651 VDD.n3206 VDD.n659 10.6151
R15652 VDD.n3216 VDD.n659 10.6151
R15653 VDD.n3217 VDD.n3216 10.6151
R15654 VDD.n3218 VDD.n3217 10.6151
R15655 VDD.n3218 VDD.n647 10.6151
R15656 VDD.n3228 VDD.n647 10.6151
R15657 VDD.n3229 VDD.n3228 10.6151
R15658 VDD.n3230 VDD.n3229 10.6151
R15659 VDD.n3230 VDD.n635 10.6151
R15660 VDD.n3240 VDD.n635 10.6151
R15661 VDD.n3241 VDD.n3240 10.6151
R15662 VDD.n3242 VDD.n3241 10.6151
R15663 VDD.n3242 VDD.n623 10.6151
R15664 VDD.n3252 VDD.n623 10.6151
R15665 VDD.n3253 VDD.n3252 10.6151
R15666 VDD.n3254 VDD.n3253 10.6151
R15667 VDD.n3254 VDD.n611 10.6151
R15668 VDD.n3264 VDD.n611 10.6151
R15669 VDD.n3265 VDD.n3264 10.6151
R15670 VDD.n3266 VDD.n3265 10.6151
R15671 VDD.n3266 VDD.n599 10.6151
R15672 VDD.n3276 VDD.n599 10.6151
R15673 VDD.n3277 VDD.n3276 10.6151
R15674 VDD.n3278 VDD.n3277 10.6151
R15675 VDD.n3278 VDD.n587 10.6151
R15676 VDD.n3288 VDD.n587 10.6151
R15677 VDD.n3289 VDD.n3288 10.6151
R15678 VDD.n3290 VDD.n3289 10.6151
R15679 VDD.n3290 VDD.n576 10.6151
R15680 VDD.n3300 VDD.n576 10.6151
R15681 VDD.n3301 VDD.n3300 10.6151
R15682 VDD.n3302 VDD.n3301 10.6151
R15683 VDD.n3302 VDD.n564 10.6151
R15684 VDD.n3312 VDD.n564 10.6151
R15685 VDD.n3313 VDD.n3312 10.6151
R15686 VDD.n3314 VDD.n3313 10.6151
R15687 VDD.n3314 VDD.n552 10.6151
R15688 VDD.n3324 VDD.n552 10.6151
R15689 VDD.n3325 VDD.n3324 10.6151
R15690 VDD.n3328 VDD.n3325 10.6151
R15691 VDD.n3328 VDD.n3327 10.6151
R15692 VDD.n3327 VDD.n3326 10.6151
R15693 VDD.n3326 VDD.n522 10.6151
R15694 VDD.n3392 VDD.n522 10.6151
R15695 VDD.n3392 VDD.n3391 10.6151
R15696 VDD.n3391 VDD.n3390 10.6151
R15697 VDD.n3390 VDD.n3389 10.6151
R15698 VDD.n2400 VDD.n2399 10.6151
R15699 VDD.n2401 VDD.n2400 10.6151
R15700 VDD.n2401 VDD.n1043 10.6151
R15701 VDD.n2411 VDD.n1043 10.6151
R15702 VDD.n2412 VDD.n2411 10.6151
R15703 VDD.n2413 VDD.n2412 10.6151
R15704 VDD.n2413 VDD.n1030 10.6151
R15705 VDD.n2423 VDD.n1030 10.6151
R15706 VDD.n2424 VDD.n2423 10.6151
R15707 VDD.n2425 VDD.n2424 10.6151
R15708 VDD.n2425 VDD.n1019 10.6151
R15709 VDD.n2435 VDD.n1019 10.6151
R15710 VDD.n2436 VDD.n2435 10.6151
R15711 VDD.n2437 VDD.n2436 10.6151
R15712 VDD.n2437 VDD.n1007 10.6151
R15713 VDD.n2447 VDD.n1007 10.6151
R15714 VDD.n2448 VDD.n2447 10.6151
R15715 VDD.n2449 VDD.n2448 10.6151
R15716 VDD.n2449 VDD.n995 10.6151
R15717 VDD.n2459 VDD.n995 10.6151
R15718 VDD.n2460 VDD.n2459 10.6151
R15719 VDD.n2461 VDD.n2460 10.6151
R15720 VDD.n2461 VDD.n983 10.6151
R15721 VDD.n2471 VDD.n983 10.6151
R15722 VDD.n2472 VDD.n2471 10.6151
R15723 VDD.n2473 VDD.n2472 10.6151
R15724 VDD.n2473 VDD.n971 10.6151
R15725 VDD.n2483 VDD.n971 10.6151
R15726 VDD.n2484 VDD.n2483 10.6151
R15727 VDD.n2485 VDD.n2484 10.6151
R15728 VDD.n2485 VDD.n959 10.6151
R15729 VDD.n2495 VDD.n959 10.6151
R15730 VDD.n2496 VDD.n2495 10.6151
R15731 VDD.n2497 VDD.n2496 10.6151
R15732 VDD.n2497 VDD.n947 10.6151
R15733 VDD.n2507 VDD.n947 10.6151
R15734 VDD.n2508 VDD.n2507 10.6151
R15735 VDD.n2509 VDD.n2508 10.6151
R15736 VDD.n2509 VDD.n934 10.6151
R15737 VDD.n2519 VDD.n934 10.6151
R15738 VDD.n2520 VDD.n2519 10.6151
R15739 VDD.n2521 VDD.n2520 10.6151
R15740 VDD.n2521 VDD.n923 10.6151
R15741 VDD.n2531 VDD.n923 10.6151
R15742 VDD.n2532 VDD.n2531 10.6151
R15743 VDD.n2533 VDD.n2532 10.6151
R15744 VDD.n2533 VDD.n911 10.6151
R15745 VDD.n2543 VDD.n911 10.6151
R15746 VDD.n2544 VDD.n2543 10.6151
R15747 VDD.n2545 VDD.n2544 10.6151
R15748 VDD.n2545 VDD.n899 10.6151
R15749 VDD.n2555 VDD.n899 10.6151
R15750 VDD.n2556 VDD.n2555 10.6151
R15751 VDD.n2557 VDD.n2556 10.6151
R15752 VDD.n2557 VDD.n886 10.6151
R15753 VDD.n2567 VDD.n886 10.6151
R15754 VDD.n2568 VDD.n2567 10.6151
R15755 VDD.n2569 VDD.n2568 10.6151
R15756 VDD.n2569 VDD.n875 10.6151
R15757 VDD.n2579 VDD.n875 10.6151
R15758 VDD.n2580 VDD.n2579 10.6151
R15759 VDD.n2581 VDD.n2580 10.6151
R15760 VDD.n2581 VDD.n863 10.6151
R15761 VDD.n2591 VDD.n863 10.6151
R15762 VDD.n2592 VDD.n2591 10.6151
R15763 VDD.n2593 VDD.n2592 10.6151
R15764 VDD.n2593 VDD.n851 10.6151
R15765 VDD.n2603 VDD.n851 10.6151
R15766 VDD.n2604 VDD.n2603 10.6151
R15767 VDD.n2605 VDD.n2604 10.6151
R15768 VDD.n2605 VDD.n839 10.6151
R15769 VDD.n2615 VDD.n839 10.6151
R15770 VDD.n2616 VDD.n2615 10.6151
R15771 VDD.n2617 VDD.n2616 10.6151
R15772 VDD.n2617 VDD.n827 10.6151
R15773 VDD.n2627 VDD.n827 10.6151
R15774 VDD.n2628 VDD.n2627 10.6151
R15775 VDD.n2634 VDD.n2628 10.6151
R15776 VDD.n2634 VDD.n2633 10.6151
R15777 VDD.n2633 VDD.n2632 10.6151
R15778 VDD.n2632 VDD.n2631 10.6151
R15779 VDD.n2631 VDD.n2629 10.6151
R15780 VDD.n2629 VDD.n800 10.6151
R15781 VDD.n2741 VDD.n2740 10.6151
R15782 VDD.n2740 VDD.n2739 10.6151
R15783 VDD.n2739 VDD.n2736 10.6151
R15784 VDD.n2736 VDD.n2735 10.6151
R15785 VDD.n2735 VDD.n2732 10.6151
R15786 VDD.n2732 VDD.n2731 10.6151
R15787 VDD.n2731 VDD.n2728 10.6151
R15788 VDD.n2728 VDD.n2727 10.6151
R15789 VDD.n2727 VDD.n2724 10.6151
R15790 VDD.n2724 VDD.n2723 10.6151
R15791 VDD.n2723 VDD.n2720 10.6151
R15792 VDD.n2720 VDD.n2719 10.6151
R15793 VDD.n2719 VDD.n2716 10.6151
R15794 VDD.n2716 VDD.n2715 10.6151
R15795 VDD.n2715 VDD.n2712 10.6151
R15796 VDD.n2712 VDD.n2711 10.6151
R15797 VDD.n2711 VDD.n2708 10.6151
R15798 VDD.n2708 VDD.n2707 10.6151
R15799 VDD.n2707 VDD.n2704 10.6151
R15800 VDD.n2702 VDD.n2700 10.6151
R15801 VDD.n2387 VDD.n2386 10.6151
R15802 VDD.n2386 VDD.n2384 10.6151
R15803 VDD.n2384 VDD.n2383 10.6151
R15804 VDD.n2383 VDD.n2381 10.6151
R15805 VDD.n2381 VDD.n2380 10.6151
R15806 VDD.n2380 VDD.n2378 10.6151
R15807 VDD.n2378 VDD.n2377 10.6151
R15808 VDD.n2377 VDD.n2375 10.6151
R15809 VDD.n2375 VDD.n2374 10.6151
R15810 VDD.n2374 VDD.n2372 10.6151
R15811 VDD.n2372 VDD.n2371 10.6151
R15812 VDD.n2371 VDD.n2369 10.6151
R15813 VDD.n2369 VDD.n2368 10.6151
R15814 VDD.n2368 VDD.n2366 10.6151
R15815 VDD.n2366 VDD.n2365 10.6151
R15816 VDD.n2365 VDD.n2363 10.6151
R15817 VDD.n2363 VDD.n2362 10.6151
R15818 VDD.n2362 VDD.n2360 10.6151
R15819 VDD.n2360 VDD.n2359 10.6151
R15820 VDD.n2359 VDD.n2357 10.6151
R15821 VDD.n2357 VDD.n2356 10.6151
R15822 VDD.n2356 VDD.n2354 10.6151
R15823 VDD.n2354 VDD.n2353 10.6151
R15824 VDD.n2353 VDD.n2351 10.6151
R15825 VDD.n2351 VDD.n2350 10.6151
R15826 VDD.n2350 VDD.n2348 10.6151
R15827 VDD.n2348 VDD.n2347 10.6151
R15828 VDD.n2347 VDD.n2345 10.6151
R15829 VDD.n2345 VDD.n2344 10.6151
R15830 VDD.n2344 VDD.n2342 10.6151
R15831 VDD.n2342 VDD.n2341 10.6151
R15832 VDD.n2341 VDD.n2339 10.6151
R15833 VDD.n2339 VDD.n2338 10.6151
R15834 VDD.n2338 VDD.n2336 10.6151
R15835 VDD.n2336 VDD.n2335 10.6151
R15836 VDD.n2335 VDD.n2333 10.6151
R15837 VDD.n2333 VDD.n2332 10.6151
R15838 VDD.n2332 VDD.n2330 10.6151
R15839 VDD.n2330 VDD.n2329 10.6151
R15840 VDD.n2329 VDD.n2327 10.6151
R15841 VDD.n2327 VDD.n2326 10.6151
R15842 VDD.n2326 VDD.n2324 10.6151
R15843 VDD.n2324 VDD.n2323 10.6151
R15844 VDD.n2323 VDD.n2321 10.6151
R15845 VDD.n2321 VDD.n2320 10.6151
R15846 VDD.n2320 VDD.n2318 10.6151
R15847 VDD.n2318 VDD.n2317 10.6151
R15848 VDD.n2317 VDD.n2315 10.6151
R15849 VDD.n2315 VDD.n2314 10.6151
R15850 VDD.n2314 VDD.n2312 10.6151
R15851 VDD.n2312 VDD.n2311 10.6151
R15852 VDD.n2311 VDD.n2309 10.6151
R15853 VDD.n2309 VDD.n2308 10.6151
R15854 VDD.n2308 VDD.n2306 10.6151
R15855 VDD.n2306 VDD.n2305 10.6151
R15856 VDD.n2305 VDD.n2303 10.6151
R15857 VDD.n2303 VDD.n2302 10.6151
R15858 VDD.n2302 VDD.n2300 10.6151
R15859 VDD.n2300 VDD.n2299 10.6151
R15860 VDD.n2299 VDD.n2297 10.6151
R15861 VDD.n2297 VDD.n2296 10.6151
R15862 VDD.n2296 VDD.n2294 10.6151
R15863 VDD.n2294 VDD.n2293 10.6151
R15864 VDD.n2293 VDD.n2291 10.6151
R15865 VDD.n2291 VDD.n2290 10.6151
R15866 VDD.n2290 VDD.n2288 10.6151
R15867 VDD.n2288 VDD.n2287 10.6151
R15868 VDD.n2287 VDD.n2285 10.6151
R15869 VDD.n2285 VDD.n2284 10.6151
R15870 VDD.n2284 VDD.n2282 10.6151
R15871 VDD.n2282 VDD.n2281 10.6151
R15872 VDD.n2281 VDD.n2279 10.6151
R15873 VDD.n2279 VDD.n2278 10.6151
R15874 VDD.n2278 VDD.n2276 10.6151
R15875 VDD.n2276 VDD.n2275 10.6151
R15876 VDD.n2275 VDD.n2273 10.6151
R15877 VDD.n2273 VDD.n2272 10.6151
R15878 VDD.n2272 VDD.n2270 10.6151
R15879 VDD.n2270 VDD.n2269 10.6151
R15880 VDD.n2269 VDD.n2267 10.6151
R15881 VDD.n2267 VDD.n2266 10.6151
R15882 VDD.n2266 VDD.n803 10.6151
R15883 VDD.n2699 VDD.n803 10.6151
R15884 VDD.n2227 VDD.n1055 10.6151
R15885 VDD.n2228 VDD.n2227 10.6151
R15886 VDD.n2231 VDD.n2228 10.6151
R15887 VDD.n2232 VDD.n2231 10.6151
R15888 VDD.n2235 VDD.n2232 10.6151
R15889 VDD.n2236 VDD.n2235 10.6151
R15890 VDD.n2239 VDD.n2236 10.6151
R15891 VDD.n2240 VDD.n2239 10.6151
R15892 VDD.n2243 VDD.n2240 10.6151
R15893 VDD.n2244 VDD.n2243 10.6151
R15894 VDD.n2248 VDD.n2247 10.6151
R15895 VDD.n2251 VDD.n2248 10.6151
R15896 VDD.n2252 VDD.n2251 10.6151
R15897 VDD.n2255 VDD.n2252 10.6151
R15898 VDD.n2256 VDD.n2255 10.6151
R15899 VDD.n2259 VDD.n2256 10.6151
R15900 VDD.n2260 VDD.n2259 10.6151
R15901 VDD.n2263 VDD.n2260 10.6151
R15902 VDD.n2388 VDD.n2265 10.6151
R15903 VDD.n1005 VDD.t21 10.2661
R15904 VDD.n3292 VDD.t7 10.2661
R15905 VDD.t20 VDD.n991 10.0921
R15906 VDD.n2583 VDD.t18 10.0921
R15907 VDD.t177 VDD.n709 10.0921
R15908 VDD.n3286 VDD.t4 10.0921
R15909 VDD.n2199 VDD.n2197 9.94894
R15910 VDD.n3452 VDD.n3451 9.94894
R15911 VDD.n3564 VDD.n459 9.94894
R15912 VDD.n2225 VDD.n2224 9.94894
R15913 VDD.n1504 VDD.t52 9.91808
R15914 VDD.t42 VDD.n1111 9.91808
R15915 VDD.n3596 VDD.t34 9.91808
R15916 VDD.t38 VDD.n3892 9.91808
R15917 VDD.t6 VDD.n895 9.74409
R15918 VDD.n3190 VDD.t19 9.74409
R15919 VDD.n2427 VDD.t175 9.5701
R15920 VDD.n562 VDD.t31 9.5701
R15921 VDD.n142 VDD.n141 9.45567
R15922 VDD.n129 VDD.n128 9.45567
R15923 VDD.n116 VDD.n115 9.45567
R15924 VDD.n103 VDD.n102 9.45567
R15925 VDD.n90 VDD.n89 9.45567
R15926 VDD.n77 VDD.n76 9.45567
R15927 VDD.n64 VDD.n63 9.45567
R15928 VDD.n51 VDD.n50 9.45567
R15929 VDD.n39 VDD.n38 9.45567
R15930 VDD.n26 VDD.n25 9.45567
R15931 VDD.n1735 VDD.n1734 9.45567
R15932 VDD.n1748 VDD.n1747 9.45567
R15933 VDD.n1709 VDD.n1708 9.45567
R15934 VDD.n1722 VDD.n1721 9.45567
R15935 VDD.n1683 VDD.n1682 9.45567
R15936 VDD.n1696 VDD.n1695 9.45567
R15937 VDD.n1657 VDD.n1656 9.45567
R15938 VDD.n1670 VDD.n1669 9.45567
R15939 VDD.n1632 VDD.n1631 9.45567
R15940 VDD.n1645 VDD.n1644 9.45567
R15941 VDD.n2028 VDD.n2027 9.3005
R15942 VDD.n2026 VDD.n1906 9.3005
R15943 VDD.n2025 VDD.n2024 9.3005
R15944 VDD.n1908 VDD.n1907 9.3005
R15945 VDD.n1913 VDD.n1911 9.3005
R15946 VDD.n2017 VDD.n1914 9.3005
R15947 VDD.n2016 VDD.n1915 9.3005
R15948 VDD.n2015 VDD.n1916 9.3005
R15949 VDD.n1922 VDD.n1919 9.3005
R15950 VDD.n2010 VDD.n1923 9.3005
R15951 VDD.n2009 VDD.n1924 9.3005
R15952 VDD.n2008 VDD.n1925 9.3005
R15953 VDD.n1929 VDD.n1926 9.3005
R15954 VDD.n2003 VDD.n1930 9.3005
R15955 VDD.n2002 VDD.n1931 9.3005
R15956 VDD.n2001 VDD.n1932 9.3005
R15957 VDD.n1936 VDD.n1933 9.3005
R15958 VDD.n1996 VDD.n1937 9.3005
R15959 VDD.n1992 VDD.n1938 9.3005
R15960 VDD.n1991 VDD.n1939 9.3005
R15961 VDD.n1943 VDD.n1940 9.3005
R15962 VDD.n1986 VDD.n1944 9.3005
R15963 VDD.n1985 VDD.n1945 9.3005
R15964 VDD.n1984 VDD.n1946 9.3005
R15965 VDD.n1950 VDD.n1947 9.3005
R15966 VDD.n1979 VDD.n1951 9.3005
R15967 VDD.n1978 VDD.n1952 9.3005
R15968 VDD.n1977 VDD.n1976 9.3005
R15969 VDD.n1975 VDD.n1953 9.3005
R15970 VDD.n1974 VDD.n1973 9.3005
R15971 VDD.n1958 VDD.n1085 9.3005
R15972 VDD.n2031 VDD.n1902 9.3005
R15973 VDD.n2206 VDD.n1897 9.3005
R15974 VDD.n2198 VDD.n1898 9.3005
R15975 VDD.n2208 VDD.n2207 9.3005
R15976 VDD.n1199 VDD.n1198 9.3005
R15977 VDD.n1767 VDD.n1766 9.3005
R15978 VDD.n1768 VDD.n1197 9.3005
R15979 VDD.n1770 VDD.n1769 9.3005
R15980 VDD.n1187 VDD.n1186 9.3005
R15981 VDD.n1783 VDD.n1782 9.3005
R15982 VDD.n1784 VDD.n1185 9.3005
R15983 VDD.n1786 VDD.n1785 9.3005
R15984 VDD.n1175 VDD.n1174 9.3005
R15985 VDD.n1799 VDD.n1798 9.3005
R15986 VDD.n1800 VDD.n1173 9.3005
R15987 VDD.n1802 VDD.n1801 9.3005
R15988 VDD.n1163 VDD.n1162 9.3005
R15989 VDD.n1815 VDD.n1814 9.3005
R15990 VDD.n1816 VDD.n1161 9.3005
R15991 VDD.n1818 VDD.n1817 9.3005
R15992 VDD.n1151 VDD.n1150 9.3005
R15993 VDD.n1831 VDD.n1830 9.3005
R15994 VDD.n1832 VDD.n1149 9.3005
R15995 VDD.n1834 VDD.n1833 9.3005
R15996 VDD.n1139 VDD.n1138 9.3005
R15997 VDD.n1847 VDD.n1846 9.3005
R15998 VDD.n1848 VDD.n1137 9.3005
R15999 VDD.n1850 VDD.n1849 9.3005
R16000 VDD.n1127 VDD.n1126 9.3005
R16001 VDD.n1863 VDD.n1862 9.3005
R16002 VDD.n1864 VDD.n1125 9.3005
R16003 VDD.n1866 VDD.n1865 9.3005
R16004 VDD.n1115 VDD.n1114 9.3005
R16005 VDD.n1879 VDD.n1878 9.3005
R16006 VDD.n1880 VDD.n1113 9.3005
R16007 VDD.n1882 VDD.n1881 9.3005
R16008 VDD.n1103 VDD.n1102 9.3005
R16009 VDD.n1895 VDD.n1894 9.3005
R16010 VDD.n1896 VDD.n1101 9.3005
R16011 VDD.n2210 VDD.n2209 9.3005
R16012 VDD.n141 VDD.n140 9.3005
R16013 VDD.n134 VDD.n133 9.3005
R16014 VDD.n128 VDD.n127 9.3005
R16015 VDD.n121 VDD.n120 9.3005
R16016 VDD.n115 VDD.n114 9.3005
R16017 VDD.n108 VDD.n107 9.3005
R16018 VDD.n102 VDD.n101 9.3005
R16019 VDD.n95 VDD.n94 9.3005
R16020 VDD.n89 VDD.n88 9.3005
R16021 VDD.n82 VDD.n81 9.3005
R16022 VDD.n76 VDD.n75 9.3005
R16023 VDD.n69 VDD.n68 9.3005
R16024 VDD.n63 VDD.n62 9.3005
R16025 VDD.n56 VDD.n55 9.3005
R16026 VDD.n50 VDD.n49 9.3005
R16027 VDD.n43 VDD.n42 9.3005
R16028 VDD.n38 VDD.n37 9.3005
R16029 VDD.n31 VDD.n30 9.3005
R16030 VDD.n25 VDD.n24 9.3005
R16031 VDD.n18 VDD.n17 9.3005
R16032 VDD.n3553 VDD.n3552 9.3005
R16033 VDD.n464 VDD.n463 9.3005
R16034 VDD.n3544 VDD.n3543 9.3005
R16035 VDD.n3542 VDD.n466 9.3005
R16036 VDD.n3541 VDD.n3540 9.3005
R16037 VDD.n468 VDD.n467 9.3005
R16038 VDD.n3534 VDD.n3533 9.3005
R16039 VDD.n3532 VDD.n470 9.3005
R16040 VDD.n3531 VDD.n3530 9.3005
R16041 VDD.n472 VDD.n471 9.3005
R16042 VDD.n3524 VDD.n3520 9.3005
R16043 VDD.n3519 VDD.n474 9.3005
R16044 VDD.n3518 VDD.n3517 9.3005
R16045 VDD.n476 VDD.n475 9.3005
R16046 VDD.n3511 VDD.n3510 9.3005
R16047 VDD.n3509 VDD.n478 9.3005
R16048 VDD.n3508 VDD.n3507 9.3005
R16049 VDD.n480 VDD.n479 9.3005
R16050 VDD.n3501 VDD.n3500 9.3005
R16051 VDD.n3498 VDD.n3497 9.3005
R16052 VDD.n486 VDD.n485 9.3005
R16053 VDD.n3491 VDD.n3490 9.3005
R16054 VDD.n3489 VDD.n488 9.3005
R16055 VDD.n3488 VDD.n3487 9.3005
R16056 VDD.n490 VDD.n489 9.3005
R16057 VDD.n3481 VDD.n3480 9.3005
R16058 VDD.n3479 VDD.n492 9.3005
R16059 VDD.n3499 VDD.n484 9.3005
R16060 VDD.n3478 VDD.n3477 9.3005
R16061 VDD.n3461 VDD.n3459 9.3005
R16062 VDD.n3463 VDD.n3462 9.3005
R16063 VDD.n3460 VDD.n446 9.3005
R16064 VDD.n3584 VDD.n445 9.3005
R16065 VDD.n3586 VDD.n3585 9.3005
R16066 VDD.n435 VDD.n434 9.3005
R16067 VDD.n3600 VDD.n3599 9.3005
R16068 VDD.n3601 VDD.n433 9.3005
R16069 VDD.n3603 VDD.n3602 9.3005
R16070 VDD.n424 VDD.n423 9.3005
R16071 VDD.n3616 VDD.n3615 9.3005
R16072 VDD.n3617 VDD.n422 9.3005
R16073 VDD.n3619 VDD.n3618 9.3005
R16074 VDD.n412 VDD.n411 9.3005
R16075 VDD.n3632 VDD.n3631 9.3005
R16076 VDD.n3633 VDD.n410 9.3005
R16077 VDD.n3635 VDD.n3634 9.3005
R16078 VDD.n400 VDD.n399 9.3005
R16079 VDD.n3648 VDD.n3647 9.3005
R16080 VDD.n3649 VDD.n398 9.3005
R16081 VDD.n3651 VDD.n3650 9.3005
R16082 VDD.n388 VDD.n387 9.3005
R16083 VDD.n3664 VDD.n3663 9.3005
R16084 VDD.n3665 VDD.n386 9.3005
R16085 VDD.n3667 VDD.n3666 9.3005
R16086 VDD.n376 VDD.n375 9.3005
R16087 VDD.n3680 VDD.n3679 9.3005
R16088 VDD.n3681 VDD.n374 9.3005
R16089 VDD.n3683 VDD.n3682 9.3005
R16090 VDD.n364 VDD.n363 9.3005
R16091 VDD.n3697 VDD.n3696 9.3005
R16092 VDD.n3698 VDD.n362 9.3005
R16093 VDD.n3700 VDD.n3699 9.3005
R16094 VDD.n353 VDD.n352 9.3005
R16095 VDD.n3716 VDD.n3715 9.3005
R16096 VDD.n3717 VDD.n351 9.3005
R16097 VDD.n3719 VDD.n3718 9.3005
R16098 VDD.n147 VDD.n145 9.3005
R16099 VDD.n3583 VDD.n3582 9.3005
R16100 VDD.n3953 VDD.n3952 9.3005
R16101 VDD.n148 VDD.n146 9.3005
R16102 VDD.n3946 VDD.n157 9.3005
R16103 VDD.n3945 VDD.n158 9.3005
R16104 VDD.n3944 VDD.n159 9.3005
R16105 VDD.n167 VDD.n160 9.3005
R16106 VDD.n3938 VDD.n168 9.3005
R16107 VDD.n3937 VDD.n169 9.3005
R16108 VDD.n3936 VDD.n170 9.3005
R16109 VDD.n178 VDD.n171 9.3005
R16110 VDD.n3930 VDD.n179 9.3005
R16111 VDD.n3929 VDD.n180 9.3005
R16112 VDD.n3928 VDD.n181 9.3005
R16113 VDD.n189 VDD.n182 9.3005
R16114 VDD.n3922 VDD.n190 9.3005
R16115 VDD.n3921 VDD.n191 9.3005
R16116 VDD.n3920 VDD.n192 9.3005
R16117 VDD.n200 VDD.n193 9.3005
R16118 VDD.n3914 VDD.n201 9.3005
R16119 VDD.n3913 VDD.n202 9.3005
R16120 VDD.n3912 VDD.n203 9.3005
R16121 VDD.n211 VDD.n204 9.3005
R16122 VDD.n3906 VDD.n212 9.3005
R16123 VDD.n3905 VDD.n213 9.3005
R16124 VDD.n3904 VDD.n214 9.3005
R16125 VDD.n222 VDD.n215 9.3005
R16126 VDD.n3898 VDD.n223 9.3005
R16127 VDD.n3897 VDD.n224 9.3005
R16128 VDD.n3896 VDD.n225 9.3005
R16129 VDD.n233 VDD.n226 9.3005
R16130 VDD.n3890 VDD.n234 9.3005
R16131 VDD.n3889 VDD.n235 9.3005
R16132 VDD.n3888 VDD.n236 9.3005
R16133 VDD.n244 VDD.n237 9.3005
R16134 VDD.n3882 VDD.n245 9.3005
R16135 VDD.n3881 VDD.n3880 9.3005
R16136 VDD.n247 VDD.n246 9.3005
R16137 VDD.n251 VDD.n249 9.3005
R16138 VDD.n3871 VDD.n252 9.3005
R16139 VDD.n3870 VDD.n253 9.3005
R16140 VDD.n3869 VDD.n254 9.3005
R16141 VDD.n261 VDD.n255 9.3005
R16142 VDD.n3864 VDD.n3863 9.3005
R16143 VDD.n3862 VDD.n258 9.3005
R16144 VDD.n3861 VDD.n3860 9.3005
R16145 VDD.n263 VDD.n262 9.3005
R16146 VDD.n3855 VDD.n266 9.3005
R16147 VDD.n3854 VDD.n267 9.3005
R16148 VDD.n3853 VDD.n268 9.3005
R16149 VDD.n272 VDD.n269 9.3005
R16150 VDD.n3848 VDD.n273 9.3005
R16151 VDD.n3847 VDD.n3846 9.3005
R16152 VDD.n3845 VDD.n274 9.3005
R16153 VDD.n3844 VDD.n3843 9.3005
R16154 VDD.n278 VDD.n277 9.3005
R16155 VDD.n283 VDD.n281 9.3005
R16156 VDD.n3836 VDD.n284 9.3005
R16157 VDD.n3835 VDD.n285 9.3005
R16158 VDD.n3834 VDD.n286 9.3005
R16159 VDD.n290 VDD.n287 9.3005
R16160 VDD.n3829 VDD.n291 9.3005
R16161 VDD.n3825 VDD.n292 9.3005
R16162 VDD.n3824 VDD.n293 9.3005
R16163 VDD.n297 VDD.n294 9.3005
R16164 VDD.n3819 VDD.n298 9.3005
R16165 VDD.n3818 VDD.n299 9.3005
R16166 VDD.n3817 VDD.n300 9.3005
R16167 VDD.n304 VDD.n301 9.3005
R16168 VDD.n3812 VDD.n305 9.3005
R16169 VDD.n3811 VDD.n306 9.3005
R16170 VDD.n3810 VDD.n3809 9.3005
R16171 VDD.n3808 VDD.n307 9.3005
R16172 VDD.n3807 VDD.n3806 9.3005
R16173 VDD.n313 VDD.n312 9.3005
R16174 VDD.n3801 VDD.n317 9.3005
R16175 VDD.n3800 VDD.n318 9.3005
R16176 VDD.n3799 VDD.n319 9.3005
R16177 VDD.n323 VDD.n320 9.3005
R16178 VDD.n3794 VDD.n324 9.3005
R16179 VDD.n3793 VDD.n325 9.3005
R16180 VDD.n3789 VDD.n326 9.3005
R16181 VDD.n3879 VDD.n3878 9.3005
R16182 VDD.n441 VDD.n440 9.3005
R16183 VDD.n3591 VDD.n3590 9.3005
R16184 VDD.n3592 VDD.n439 9.3005
R16185 VDD.n3594 VDD.n3593 9.3005
R16186 VDD.n430 VDD.n429 9.3005
R16187 VDD.n3608 VDD.n3607 9.3005
R16188 VDD.n3609 VDD.n428 9.3005
R16189 VDD.n3611 VDD.n3610 9.3005
R16190 VDD.n418 VDD.n417 9.3005
R16191 VDD.n3624 VDD.n3623 9.3005
R16192 VDD.n3625 VDD.n416 9.3005
R16193 VDD.n3627 VDD.n3626 9.3005
R16194 VDD.n406 VDD.n405 9.3005
R16195 VDD.n3640 VDD.n3639 9.3005
R16196 VDD.n3641 VDD.n404 9.3005
R16197 VDD.n3643 VDD.n3642 9.3005
R16198 VDD.n394 VDD.n393 9.3005
R16199 VDD.n3656 VDD.n3655 9.3005
R16200 VDD.n3657 VDD.n392 9.3005
R16201 VDD.n3659 VDD.n3658 9.3005
R16202 VDD.n382 VDD.n381 9.3005
R16203 VDD.n3672 VDD.n3671 9.3005
R16204 VDD.n3673 VDD.n380 9.3005
R16205 VDD.n3675 VDD.n3674 9.3005
R16206 VDD.n370 VDD.n369 9.3005
R16207 VDD.n3688 VDD.n3687 9.3005
R16208 VDD.n3689 VDD.n368 9.3005
R16209 VDD.n3691 VDD.n3690 9.3005
R16210 VDD.n359 VDD.n358 9.3005
R16211 VDD.n3705 VDD.n3704 9.3005
R16212 VDD.n3706 VDD.n357 9.3005
R16213 VDD.n3711 VDD.n3707 9.3005
R16214 VDD.n3710 VDD.n3709 9.3005
R16215 VDD.n3708 VDD.n346 9.3005
R16216 VDD.n3724 VDD.n347 9.3005
R16217 VDD.n3725 VDD.n345 9.3005
R16218 VDD.n3727 VDD.n3726 9.3005
R16219 VDD.n3728 VDD.n344 9.3005
R16220 VDD.n3731 VDD.n3729 9.3005
R16221 VDD.n3732 VDD.n343 9.3005
R16222 VDD.n3734 VDD.n3733 9.3005
R16223 VDD.n3735 VDD.n342 9.3005
R16224 VDD.n3738 VDD.n3736 9.3005
R16225 VDD.n3739 VDD.n341 9.3005
R16226 VDD.n3741 VDD.n3740 9.3005
R16227 VDD.n3742 VDD.n340 9.3005
R16228 VDD.n3745 VDD.n3743 9.3005
R16229 VDD.n3746 VDD.n339 9.3005
R16230 VDD.n3748 VDD.n3747 9.3005
R16231 VDD.n3749 VDD.n338 9.3005
R16232 VDD.n3752 VDD.n3750 9.3005
R16233 VDD.n3753 VDD.n337 9.3005
R16234 VDD.n3755 VDD.n3754 9.3005
R16235 VDD.n3756 VDD.n336 9.3005
R16236 VDD.n3759 VDD.n3757 9.3005
R16237 VDD.n3760 VDD.n335 9.3005
R16238 VDD.n3762 VDD.n3761 9.3005
R16239 VDD.n3763 VDD.n334 9.3005
R16240 VDD.n3766 VDD.n3764 9.3005
R16241 VDD.n3767 VDD.n333 9.3005
R16242 VDD.n3769 VDD.n3768 9.3005
R16243 VDD.n3770 VDD.n332 9.3005
R16244 VDD.n3773 VDD.n3771 9.3005
R16245 VDD.n3774 VDD.n331 9.3005
R16246 VDD.n3776 VDD.n3775 9.3005
R16247 VDD.n3777 VDD.n330 9.3005
R16248 VDD.n3780 VDD.n3778 9.3005
R16249 VDD.n3781 VDD.n329 9.3005
R16250 VDD.n3783 VDD.n3782 9.3005
R16251 VDD.n3784 VDD.n328 9.3005
R16252 VDD.n3786 VDD.n3785 9.3005
R16253 VDD.n3578 VDD.n3577 9.3005
R16254 VDD.n3576 VDD.n3575 9.3005
R16255 VDD.n3573 VDD.n450 9.3005
R16256 VDD.n458 VDD.n453 9.3005
R16257 VDD.n460 VDD.n457 9.3005
R16258 VDD.n3556 VDD.n3555 9.3005
R16259 VDD.n3554 VDD.n462 9.3005
R16260 VDD.n2223 VDD.n2222 9.3005
R16261 VDD.n2221 VDD.n1088 9.3005
R16262 VDD.n2217 VDD.n2216 9.3005
R16263 VDD.n1486 VDD.n1485 9.3005
R16264 VDD.n1300 VDD.n1299 9.3005
R16265 VDD.n1499 VDD.n1498 9.3005
R16266 VDD.n1500 VDD.n1298 9.3005
R16267 VDD.n1502 VDD.n1501 9.3005
R16268 VDD.n1288 VDD.n1287 9.3005
R16269 VDD.n1515 VDD.n1514 9.3005
R16270 VDD.n1516 VDD.n1286 9.3005
R16271 VDD.n1518 VDD.n1517 9.3005
R16272 VDD.n1276 VDD.n1275 9.3005
R16273 VDD.n1531 VDD.n1530 9.3005
R16274 VDD.n1532 VDD.n1274 9.3005
R16275 VDD.n1534 VDD.n1533 9.3005
R16276 VDD.n1264 VDD.n1263 9.3005
R16277 VDD.n1547 VDD.n1546 9.3005
R16278 VDD.n1548 VDD.n1262 9.3005
R16279 VDD.n1550 VDD.n1549 9.3005
R16280 VDD.n1253 VDD.n1252 9.3005
R16281 VDD.n1564 VDD.n1563 9.3005
R16282 VDD.n1565 VDD.n1251 9.3005
R16283 VDD.n1567 VDD.n1566 9.3005
R16284 VDD.n1241 VDD.n1240 9.3005
R16285 VDD.n1580 VDD.n1579 9.3005
R16286 VDD.n1581 VDD.n1239 9.3005
R16287 VDD.n1583 VDD.n1582 9.3005
R16288 VDD.n1229 VDD.n1228 9.3005
R16289 VDD.n1596 VDD.n1595 9.3005
R16290 VDD.n1597 VDD.n1227 9.3005
R16291 VDD.n1599 VDD.n1598 9.3005
R16292 VDD.n1217 VDD.n1216 9.3005
R16293 VDD.n1612 VDD.n1611 9.3005
R16294 VDD.n1613 VDD.n1215 9.3005
R16295 VDD.n1615 VDD.n1614 9.3005
R16296 VDD.n1205 VDD.n1204 9.3005
R16297 VDD.n1759 VDD.n1758 9.3005
R16298 VDD.n1760 VDD.n1203 9.3005
R16299 VDD.n1762 VDD.n1761 9.3005
R16300 VDD.n1193 VDD.n1192 9.3005
R16301 VDD.n1775 VDD.n1774 9.3005
R16302 VDD.n1776 VDD.n1191 9.3005
R16303 VDD.n1778 VDD.n1777 9.3005
R16304 VDD.n1181 VDD.n1180 9.3005
R16305 VDD.n1791 VDD.n1790 9.3005
R16306 VDD.n1792 VDD.n1179 9.3005
R16307 VDD.n1794 VDD.n1793 9.3005
R16308 VDD.n1169 VDD.n1168 9.3005
R16309 VDD.n1807 VDD.n1806 9.3005
R16310 VDD.n1808 VDD.n1167 9.3005
R16311 VDD.n1810 VDD.n1809 9.3005
R16312 VDD.n1156 VDD.n1155 9.3005
R16313 VDD.n1823 VDD.n1822 9.3005
R16314 VDD.n1824 VDD.n1154 9.3005
R16315 VDD.n1826 VDD.n1825 9.3005
R16316 VDD.n1145 VDD.n1144 9.3005
R16317 VDD.n1839 VDD.n1838 9.3005
R16318 VDD.n1840 VDD.n1143 9.3005
R16319 VDD.n1842 VDD.n1841 9.3005
R16320 VDD.n1133 VDD.n1132 9.3005
R16321 VDD.n1855 VDD.n1854 9.3005
R16322 VDD.n1856 VDD.n1131 9.3005
R16323 VDD.n1858 VDD.n1857 9.3005
R16324 VDD.n1121 VDD.n1120 9.3005
R16325 VDD.n1871 VDD.n1870 9.3005
R16326 VDD.n1872 VDD.n1119 9.3005
R16327 VDD.n1874 VDD.n1873 9.3005
R16328 VDD.n1109 VDD.n1108 9.3005
R16329 VDD.n1887 VDD.n1886 9.3005
R16330 VDD.n1888 VDD.n1107 9.3005
R16331 VDD.n1890 VDD.n1889 9.3005
R16332 VDD.n1094 VDD.n1093 9.3005
R16333 VDD.n2215 VDD.n2214 9.3005
R16334 VDD.n1484 VDD.n1310 9.3005
R16335 VDD.n1400 VDD.n1311 9.3005
R16336 VDD.n1401 VDD.n1397 9.3005
R16337 VDD.n1403 VDD.n1402 9.3005
R16338 VDD.n1404 VDD.n1396 9.3005
R16339 VDD.n1406 VDD.n1405 9.3005
R16340 VDD.n1407 VDD.n1391 9.3005
R16341 VDD.n1409 VDD.n1408 9.3005
R16342 VDD.n1410 VDD.n1390 9.3005
R16343 VDD.n1412 VDD.n1411 9.3005
R16344 VDD.n1416 VDD.n1386 9.3005
R16345 VDD.n1418 VDD.n1417 9.3005
R16346 VDD.n1419 VDD.n1385 9.3005
R16347 VDD.n1421 VDD.n1420 9.3005
R16348 VDD.n1422 VDD.n1380 9.3005
R16349 VDD.n1424 VDD.n1423 9.3005
R16350 VDD.n1425 VDD.n1379 9.3005
R16351 VDD.n1427 VDD.n1426 9.3005
R16352 VDD.n1428 VDD.n1374 9.3005
R16353 VDD.n1430 VDD.n1429 9.3005
R16354 VDD.n1432 VDD.n1431 9.3005
R16355 VDD.n1433 VDD.n1366 9.3005
R16356 VDD.n1435 VDD.n1434 9.3005
R16357 VDD.n1436 VDD.n1365 9.3005
R16358 VDD.n1438 VDD.n1437 9.3005
R16359 VDD.n1439 VDD.n1360 9.3005
R16360 VDD.n1441 VDD.n1440 9.3005
R16361 VDD.n1442 VDD.n1359 9.3005
R16362 VDD.n1444 VDD.n1443 9.3005
R16363 VDD.n1451 VDD.n1450 9.3005
R16364 VDD.n1452 VDD.n1355 9.3005
R16365 VDD.n1454 VDD.n1453 9.3005
R16366 VDD.n1455 VDD.n1350 9.3005
R16367 VDD.n1457 VDD.n1456 9.3005
R16368 VDD.n1458 VDD.n1349 9.3005
R16369 VDD.n1460 VDD.n1459 9.3005
R16370 VDD.n1461 VDD.n1346 9.3005
R16371 VDD.n1467 VDD.n1466 9.3005
R16372 VDD.n1468 VDD.n1345 9.3005
R16373 VDD.n1470 VDD.n1469 9.3005
R16374 VDD.n1471 VDD.n1341 9.3005
R16375 VDD.n1473 VDD.n1472 9.3005
R16376 VDD.n1474 VDD.n1340 9.3005
R16377 VDD.n1476 VDD.n1475 9.3005
R16378 VDD.n1477 VDD.n1339 9.3005
R16379 VDD.n1449 VDD.n1356 9.3005
R16380 VDD.n1483 VDD.n1482 9.3005
R16381 VDD.n1491 VDD.n1490 9.3005
R16382 VDD.n1492 VDD.n1304 9.3005
R16383 VDD.n1494 VDD.n1493 9.3005
R16384 VDD.n1294 VDD.n1293 9.3005
R16385 VDD.n1507 VDD.n1506 9.3005
R16386 VDD.n1508 VDD.n1292 9.3005
R16387 VDD.n1510 VDD.n1509 9.3005
R16388 VDD.n1282 VDD.n1281 9.3005
R16389 VDD.n1523 VDD.n1522 9.3005
R16390 VDD.n1524 VDD.n1280 9.3005
R16391 VDD.n1526 VDD.n1525 9.3005
R16392 VDD.n1270 VDD.n1269 9.3005
R16393 VDD.n1539 VDD.n1538 9.3005
R16394 VDD.n1540 VDD.n1268 9.3005
R16395 VDD.n1542 VDD.n1541 9.3005
R16396 VDD.n1258 VDD.n1257 9.3005
R16397 VDD.n1556 VDD.n1555 9.3005
R16398 VDD.n1557 VDD.n1256 9.3005
R16399 VDD.n1559 VDD.n1558 9.3005
R16400 VDD.n1247 VDD.n1246 9.3005
R16401 VDD.n1572 VDD.n1571 9.3005
R16402 VDD.n1573 VDD.n1245 9.3005
R16403 VDD.n1575 VDD.n1574 9.3005
R16404 VDD.n1235 VDD.n1234 9.3005
R16405 VDD.n1588 VDD.n1587 9.3005
R16406 VDD.n1589 VDD.n1233 9.3005
R16407 VDD.n1591 VDD.n1590 9.3005
R16408 VDD.n1223 VDD.n1222 9.3005
R16409 VDD.n1604 VDD.n1603 9.3005
R16410 VDD.n1605 VDD.n1221 9.3005
R16411 VDD.n1607 VDD.n1606 9.3005
R16412 VDD.n1211 VDD.n1210 9.3005
R16413 VDD.n1620 VDD.n1619 9.3005
R16414 VDD.n1621 VDD.n1209 9.3005
R16415 VDD.n1754 VDD.n1753 9.3005
R16416 VDD.n1306 VDD.n1305 9.3005
R16417 VDD.n1734 VDD.n1733 9.3005
R16418 VDD.n1727 VDD.n1726 9.3005
R16419 VDD.n1747 VDD.n1746 9.3005
R16420 VDD.n1740 VDD.n1739 9.3005
R16421 VDD.n1708 VDD.n1707 9.3005
R16422 VDD.n1701 VDD.n1700 9.3005
R16423 VDD.n1721 VDD.n1720 9.3005
R16424 VDD.n1714 VDD.n1713 9.3005
R16425 VDD.n1682 VDD.n1681 9.3005
R16426 VDD.n1675 VDD.n1674 9.3005
R16427 VDD.n1695 VDD.n1694 9.3005
R16428 VDD.n1688 VDD.n1687 9.3005
R16429 VDD.n1656 VDD.n1655 9.3005
R16430 VDD.n1649 VDD.n1648 9.3005
R16431 VDD.n1669 VDD.n1668 9.3005
R16432 VDD.n1662 VDD.n1661 9.3005
R16433 VDD.n1631 VDD.n1630 9.3005
R16434 VDD.n1624 VDD.n1623 9.3005
R16435 VDD.n1644 VDD.n1643 9.3005
R16436 VDD.n1637 VDD.n1636 9.3005
R16437 VDD.n2636 VDD.t16 8.87413
R16438 VDD.t125 VDD.n757 8.87413
R16439 VDD.t81 VDD.n1032 8.70013
R16440 VDD.n2625 VDD.t62 8.70013
R16441 VDD.t88 VDD.n751 8.70013
R16442 VDD.n3330 VDD.t113 8.70013
R16443 VDD.n2535 VDD.t10 8.52614
R16444 VDD.t180 VDD.n661 8.52614
R16445 VDD.n2651 VDD.n813 8.27367
R16446 VDD.n2177 VDD.n2176 8.27367
R16447 VDD.n2828 VDD.n2780 8.27367
R16448 VDD.n505 VDD.n503 8.27367
R16449 VDD.n3350 VDD.n3349 8.27367
R16450 VDD.n3057 VDD.n3056 8.27367
R16451 VDD.n2703 VDD.n2702 8.27367
R16452 VDD.n2265 VDD.n2264 8.27367
R16453 VDD.n15 VDD.n14 8.2594
R16454 VDD.n3955 VDD.n3954 8.09137
R16455 VDD.n1752 VDD.n1751 8.09137
R16456 VDD.t52 VDD.n1290 7.48219
R16457 VDD.n1876 VDD.t42 7.48219
R16458 VDD.n3605 VDD.t34 7.48219
R16459 VDD.n3893 VDD.t38 7.48219
R16460 VDD.n2571 VDD.t23 7.1342
R16461 VDD.n705 VDD.t27 7.1342
R16462 VDD.n66 VDD.n40 6.85826
R16463 VDD.n1672 VDD.n1646 6.85826
R16464 VDD.n1466 VDD.n1345 6.78838
R16465 VDD.n2031 VDD.n1903 6.78838
R16466 VDD.n3864 VDD.n255 6.78838
R16467 VDD.n3477 VDD.n3476 6.78838
R16468 VDD.n2487 VDD.t178 6.43823
R16469 VDD.t14 VDD.n613 6.43823
R16470 VDD.n7 VDD.t32 6.37403
R16471 VDD.n7 VDD.t1 6.37403
R16472 VDD.n8 VDD.t15 6.37403
R16473 VDD.n8 VDD.t8 6.37403
R16474 VDD.n10 VDD.t28 6.37403
R16475 VDD.n10 VDD.t181 6.37403
R16476 VDD.n12 VDD.t126 6.37403
R16477 VDD.n12 VDD.t30 6.37403
R16478 VDD.n5 VDD.t3 6.37403
R16479 VDD.n5 VDD.t17 6.37403
R16480 VDD.n3 VDD.t11 6.37403
R16481 VDD.n3 VDD.t24 6.37403
R16482 VDD.n1 VDD.t22 6.37403
R16483 VDD.n1 VDD.t179 6.37403
R16484 VDD.n0 VDD.t183 6.37403
R16485 VDD.n0 VDD.t176 6.37403
R16486 VDD.n2390 VDD.t182 5.91625
R16487 VDD.n939 VDD.t13 5.91625
R16488 VDD.n2523 VDD.t13 5.91625
R16489 VDD.n657 VDD.t5 5.91625
R16490 VDD.n3226 VDD.t5 5.91625
R16491 VDD.t0 VDD.n496 5.91625
R16492 VDD.n3955 VDD.n144 5.39442
R16493 VDD.n1751 VDD.n1750 5.39442
R16494 VDD.n2197 VDD.n2052 5.30782
R16495 VDD.n2197 VDD.n2196 5.30782
R16496 VDD.n3451 VDD.n493 5.30782
R16497 VDD.n3451 VDD.n3450 5.30782
R16498 VDD.n3369 VDD.n459 5.30782
R16499 VDD.n3365 VDD.n459 5.30782
R16500 VDD.n2244 VDD.n2225 5.30782
R16501 VDD.n2247 VDD.n2225 5.30782
R16502 VDD.n144 VDD.n143 4.88412
R16503 VDD.n118 VDD.n117 4.88412
R16504 VDD.n92 VDD.n91 4.88412
R16505 VDD.n66 VDD.n65 4.88412
R16506 VDD.n1750 VDD.n1749 4.88412
R16507 VDD.n1724 VDD.n1723 4.88412
R16508 VDD.n1698 VDD.n1697 4.88412
R16509 VDD.n1672 VDD.n1671 4.88412
R16510 VDD.n143 VDD.n131 4.78498
R16511 VDD.n117 VDD.n105 4.78498
R16512 VDD.n91 VDD.n79 4.78498
R16513 VDD.n65 VDD.n53 4.78498
R16514 VDD.n40 VDD.n28 4.78498
R16515 VDD.n1749 VDD.n1737 4.78498
R16516 VDD.n1723 VDD.n1711 4.78498
R16517 VDD.n1697 VDD.n1685 4.78498
R16518 VDD.n1671 VDD.n1659 4.78498
R16519 VDD.n1646 VDD.n1634 4.78498
R16520 VDD.n1968 VDD.n1086 4.74817
R16521 VDD.n1964 VDD.n1087 4.74817
R16522 VDD.n2201 VDD.n2200 4.74817
R16523 VDD.n2037 VDD.n1903 4.74817
R16524 VDD.n2200 VDD.n1901 4.74817
R16525 VDD.n2037 VDD.n2036 4.74817
R16526 VDD.n3470 VDD.n3469 4.74817
R16527 VDD.n3476 VDD.n3457 4.74817
R16528 VDD.n3472 VDD.n3457 4.74817
R16529 VDD.n3471 VDD.n3470 4.74817
R16530 VDD.n3563 VDD.n456 4.74817
R16531 VDD.n3565 VDD.n454 4.74817
R16532 VDD.n3566 VDD.n3565 4.74817
R16533 VDD.n3563 VDD.n3562 4.74817
R16534 VDD.n1961 VDD.n1086 4.74817
R16535 VDD.n1089 VDD.n1087 4.74817
R16536 VDD.n891 VDD.t23 4.6983
R16537 VDD.n3178 VDD.t27 4.6983
R16538 VDD.n1482 VDD.n1314 4.46111
R16539 VDD.n1432 VDD.n1373 4.46111
R16540 VDD.n2220 VDD.n2217 4.46111
R16541 VDD.n1996 VDD.n1995 4.46111
R16542 VDD.n3792 VDD.n3789 4.46111
R16543 VDD.n3829 VDD.n3828 4.46111
R16544 VDD.n3524 VDD.n3523 4.46111
R16545 VDD.n3575 VDD.n3574 4.46111
R16546 VDD.n135 VDD.n133 4.29255
R16547 VDD.n122 VDD.n120 4.29255
R16548 VDD.n109 VDD.n107 4.29255
R16549 VDD.n96 VDD.n94 4.29255
R16550 VDD.n83 VDD.n81 4.29255
R16551 VDD.n70 VDD.n68 4.29255
R16552 VDD.n57 VDD.n55 4.29255
R16553 VDD.n44 VDD.n42 4.29255
R16554 VDD.n32 VDD.n30 4.29255
R16555 VDD.n19 VDD.n17 4.29255
R16556 VDD.n1728 VDD.n1726 4.29255
R16557 VDD.n1741 VDD.n1739 4.29255
R16558 VDD.n1702 VDD.n1700 4.29255
R16559 VDD.n1715 VDD.n1713 4.29255
R16560 VDD.n1676 VDD.n1674 4.29255
R16561 VDD.n1689 VDD.n1687 4.29255
R16562 VDD.n1650 VDD.n1648 4.29255
R16563 VDD.n1663 VDD.n1661 4.29255
R16564 VDD.n1625 VDD.n1623 4.29255
R16565 VDD.n1638 VDD.n1636 4.29255
R16566 VDD.n11 VDD.n9 3.93584
R16567 VDD.n4 VDD.n2 3.93584
R16568 VDD.t178 VDD.t9 3.30636
R16569 VDD.t10 VDD.n913 3.30636
R16570 VDD.n3208 VDD.t180 3.30636
R16571 VDD.t12 VDD.t14 3.30636
R16572 VDD.n2415 VDD.t81 3.13237
R16573 VDD.t62 VDD.n822 3.13237
R16574 VDD.n3118 VDD.t88 3.13237
R16575 VDD.t113 VDD.n541 3.13237
R16576 VDD.n13 VDD.n11 3.12981
R16577 VDD.n6 VDD.n4 3.12981
R16578 VDD.t16 VDD.n816 2.95838
R16579 VDD.n3112 VDD.t125 2.95838
R16580 VDD.n1561 VDD.t129 2.61039
R16581 VDD.n1159 VDD.t131 2.61039
R16582 VDD.t135 VDD.n390 2.61039
R16583 VDD.n3918 VDD.t141 2.61039
R16584 VDD.n14 VDD.n13 2.43301
R16585 VDD.n14 VDD.n6 2.43301
R16586 VDD.n2654 VDD.n813 2.34196
R16587 VDD.n2178 VDD.n2177 2.34196
R16588 VDD.n2829 VDD.n2828 2.34196
R16589 VDD.n3436 VDD.n503 2.34196
R16590 VDD.n3351 VDD.n3350 2.34196
R16591 VDD.n3058 VDD.n3057 2.34196
R16592 VDD.n2704 VDD.n2703 2.34196
R16593 VDD.n2264 VDD.n2263 2.34196
R16594 VDD.n2200 VDD.n2199 2.27742
R16595 VDD.n2199 VDD.n2037 2.27742
R16596 VDD.n3457 VDD.n3452 2.27742
R16597 VDD.n3470 VDD.n3452 2.27742
R16598 VDD.n3565 VDD.n3564 2.27742
R16599 VDD.n3564 VDD.n3563 2.27742
R16600 VDD.n2224 VDD.n1086 2.27742
R16601 VDD.n2224 VDD.n1087 2.27742
R16602 VDD.n1035 VDD.t175 2.2624
R16603 VDD.n3322 VDD.t31 2.2624
R16604 VDD.n1400 VDD.n1314 2.13383
R16605 VDD.n1429 VDD.n1373 2.13383
R16606 VDD.n2221 VDD.n2220 2.13383
R16607 VDD.n1995 VDD.n1992 2.13383
R16608 VDD.n3793 VDD.n3792 2.13383
R16609 VDD.n3828 VDD.n3825 2.13383
R16610 VDD.n3523 VDD.n472 2.13383
R16611 VDD.n3574 VDD.n3573 2.13383
R16612 VDD.t9 VDD.n961 2.08841
R16613 VDD.n2553 VDD.t6 2.08841
R16614 VDD.t19 VDD.n679 2.08841
R16615 VDD.n3256 VDD.t12 2.08841
R16616 VDD.n92 VDD.n66 1.97464
R16617 VDD.n118 VDD.n92 1.97464
R16618 VDD.n144 VDD.n118 1.97464
R16619 VDD.n1698 VDD.n1672 1.97464
R16620 VDD.n1724 VDD.n1698 1.97464
R16621 VDD.n1750 VDD.n1724 1.97464
R16622 VDD.n142 VDD.n132 1.93989
R16623 VDD.n129 VDD.n119 1.93989
R16624 VDD.n116 VDD.n106 1.93989
R16625 VDD.n103 VDD.n93 1.93989
R16626 VDD.n90 VDD.n80 1.93989
R16627 VDD.n77 VDD.n67 1.93989
R16628 VDD.n64 VDD.n54 1.93989
R16629 VDD.n51 VDD.n41 1.93989
R16630 VDD.n39 VDD.n29 1.93989
R16631 VDD.n26 VDD.n16 1.93989
R16632 VDD.n1735 VDD.n1725 1.93989
R16633 VDD.n1748 VDD.n1738 1.93989
R16634 VDD.n1709 VDD.n1699 1.93989
R16635 VDD.n1722 VDD.n1712 1.93989
R16636 VDD.n1683 VDD.n1673 1.93989
R16637 VDD.n1696 VDD.n1686 1.93989
R16638 VDD.n1657 VDD.n1647 1.93989
R16639 VDD.n1670 VDD.n1660 1.93989
R16640 VDD.n1632 VDD.n1622 1.93989
R16641 VDD.n1645 VDD.n1635 1.93989
R16642 VDD.n1751 VDD.n15 1.86217
R16643 VDD VDD.n3955 1.85434
R16644 VDD.n2457 VDD.t20 1.74043
R16645 VDD.t18 VDD.n865 1.74043
R16646 VDD.n3160 VDD.t177 1.74043
R16647 VDD.n2956 VDD.t4 1.74043
R16648 VDD.n2457 VDD.t21 1.56643
R16649 VDD.n2956 VDD.t7 1.56643
R16650 VDD.n140 VDD.n139 1.16414
R16651 VDD.n127 VDD.n126 1.16414
R16652 VDD.n114 VDD.n113 1.16414
R16653 VDD.n101 VDD.n100 1.16414
R16654 VDD.n88 VDD.n87 1.16414
R16655 VDD.n75 VDD.n74 1.16414
R16656 VDD.n62 VDD.n61 1.16414
R16657 VDD.n49 VDD.n48 1.16414
R16658 VDD.n37 VDD.n36 1.16414
R16659 VDD.n24 VDD.n23 1.16414
R16660 VDD.n1733 VDD.n1732 1.16414
R16661 VDD.n1746 VDD.n1745 1.16414
R16662 VDD.n1707 VDD.n1706 1.16414
R16663 VDD.n1720 VDD.n1719 1.16414
R16664 VDD.n1681 VDD.n1680 1.16414
R16665 VDD.n1694 VDD.n1693 1.16414
R16666 VDD.n1655 VDD.n1654 1.16414
R16667 VDD.n1668 VDD.n1667 1.16414
R16668 VDD.n1630 VDD.n1629 1.16414
R16669 VDD.n1643 VDD.n1642 1.16414
R16670 VDD.t127 VDD.n1219 0.870463
R16671 VDD.n1780 VDD.t148 0.870463
R16672 VDD.n2601 VDD.t2 0.870463
R16673 VDD.t29 VDD.n727 0.870463
R16674 VDD.n3702 VDD.t143 0.870463
R16675 VDD.n3941 VDD.t138 0.870463
R16676 VDD.n2209 VDD.n2208 0.532512
R16677 VDD.n3583 VDD.n446 0.532512
R16678 VDD.n3880 VDD.n3879 0.532512
R16679 VDD.n3785 VDD.n326 0.532512
R16680 VDD.n3577 VDD.n3576 0.532512
R16681 VDD.n2216 VDD.n2215 0.532512
R16682 VDD.n1484 VDD.n1483 0.532512
R16683 VDD.n1339 VDD.n1305 0.532512
R16684 VDD.n136 VDD.n134 0.388379
R16685 VDD.n123 VDD.n121 0.388379
R16686 VDD.n110 VDD.n108 0.388379
R16687 VDD.n97 VDD.n95 0.388379
R16688 VDD.n84 VDD.n82 0.388379
R16689 VDD.n71 VDD.n69 0.388379
R16690 VDD.n58 VDD.n56 0.388379
R16691 VDD.n45 VDD.n43 0.388379
R16692 VDD.n33 VDD.n31 0.388379
R16693 VDD.n20 VDD.n18 0.388379
R16694 VDD.n1729 VDD.n1727 0.388379
R16695 VDD.n1742 VDD.n1740 0.388379
R16696 VDD.n1703 VDD.n1701 0.388379
R16697 VDD.n1716 VDD.n1714 0.388379
R16698 VDD.n1677 VDD.n1675 0.388379
R16699 VDD.n1690 VDD.n1688 0.388379
R16700 VDD.n1651 VDD.n1649 0.388379
R16701 VDD.n1664 VDD.n1662 0.388379
R16702 VDD.n1626 VDD.n1624 0.388379
R16703 VDD.n1639 VDD.n1637 0.388379
R16704 VDD.n141 VDD.n133 0.155672
R16705 VDD.n128 VDD.n120 0.155672
R16706 VDD.n115 VDD.n107 0.155672
R16707 VDD.n102 VDD.n94 0.155672
R16708 VDD.n89 VDD.n81 0.155672
R16709 VDD.n76 VDD.n68 0.155672
R16710 VDD.n63 VDD.n55 0.155672
R16711 VDD.n50 VDD.n42 0.155672
R16712 VDD.n38 VDD.n30 0.155672
R16713 VDD.n25 VDD.n17 0.155672
R16714 VDD.n1734 VDD.n1726 0.155672
R16715 VDD.n1747 VDD.n1739 0.155672
R16716 VDD.n1708 VDD.n1700 0.155672
R16717 VDD.n1721 VDD.n1713 0.155672
R16718 VDD.n1682 VDD.n1674 0.155672
R16719 VDD.n1695 VDD.n1687 0.155672
R16720 VDD.n1656 VDD.n1648 0.155672
R16721 VDD.n1669 VDD.n1661 0.155672
R16722 VDD.n1631 VDD.n1623 0.155672
R16723 VDD.n1644 VDD.n1636 0.155672
R16724 VDD.n2027 VDD.n1902 0.152939
R16725 VDD.n2027 VDD.n2026 0.152939
R16726 VDD.n2026 VDD.n2025 0.152939
R16727 VDD.n2025 VDD.n1907 0.152939
R16728 VDD.n1913 VDD.n1907 0.152939
R16729 VDD.n1914 VDD.n1913 0.152939
R16730 VDD.n1915 VDD.n1914 0.152939
R16731 VDD.n1916 VDD.n1915 0.152939
R16732 VDD.n1922 VDD.n1916 0.152939
R16733 VDD.n1923 VDD.n1922 0.152939
R16734 VDD.n1924 VDD.n1923 0.152939
R16735 VDD.n1925 VDD.n1924 0.152939
R16736 VDD.n1929 VDD.n1925 0.152939
R16737 VDD.n1930 VDD.n1929 0.152939
R16738 VDD.n1931 VDD.n1930 0.152939
R16739 VDD.n1932 VDD.n1931 0.152939
R16740 VDD.n1936 VDD.n1932 0.152939
R16741 VDD.n1937 VDD.n1936 0.152939
R16742 VDD.n1938 VDD.n1937 0.152939
R16743 VDD.n1939 VDD.n1938 0.152939
R16744 VDD.n1943 VDD.n1939 0.152939
R16745 VDD.n1944 VDD.n1943 0.152939
R16746 VDD.n1945 VDD.n1944 0.152939
R16747 VDD.n1946 VDD.n1945 0.152939
R16748 VDD.n1950 VDD.n1946 0.152939
R16749 VDD.n1951 VDD.n1950 0.152939
R16750 VDD.n1952 VDD.n1951 0.152939
R16751 VDD.n1976 VDD.n1952 0.152939
R16752 VDD.n1976 VDD.n1975 0.152939
R16753 VDD.n1975 VDD.n1974 0.152939
R16754 VDD.n1974 VDD.n1085 0.152939
R16755 VDD.n2208 VDD.n1897 0.152939
R16756 VDD.n2198 VDD.n1897 0.152939
R16757 VDD.n1767 VDD.n1198 0.152939
R16758 VDD.n1768 VDD.n1767 0.152939
R16759 VDD.n1769 VDD.n1768 0.152939
R16760 VDD.n1769 VDD.n1186 0.152939
R16761 VDD.n1783 VDD.n1186 0.152939
R16762 VDD.n1784 VDD.n1783 0.152939
R16763 VDD.n1785 VDD.n1784 0.152939
R16764 VDD.n1785 VDD.n1174 0.152939
R16765 VDD.n1799 VDD.n1174 0.152939
R16766 VDD.n1800 VDD.n1799 0.152939
R16767 VDD.n1801 VDD.n1800 0.152939
R16768 VDD.n1801 VDD.n1162 0.152939
R16769 VDD.n1815 VDD.n1162 0.152939
R16770 VDD.n1816 VDD.n1815 0.152939
R16771 VDD.n1817 VDD.n1816 0.152939
R16772 VDD.n1817 VDD.n1150 0.152939
R16773 VDD.n1831 VDD.n1150 0.152939
R16774 VDD.n1832 VDD.n1831 0.152939
R16775 VDD.n1833 VDD.n1832 0.152939
R16776 VDD.n1833 VDD.n1138 0.152939
R16777 VDD.n1847 VDD.n1138 0.152939
R16778 VDD.n1848 VDD.n1847 0.152939
R16779 VDD.n1849 VDD.n1848 0.152939
R16780 VDD.n1849 VDD.n1126 0.152939
R16781 VDD.n1863 VDD.n1126 0.152939
R16782 VDD.n1864 VDD.n1863 0.152939
R16783 VDD.n1865 VDD.n1864 0.152939
R16784 VDD.n1865 VDD.n1114 0.152939
R16785 VDD.n1879 VDD.n1114 0.152939
R16786 VDD.n1880 VDD.n1879 0.152939
R16787 VDD.n1881 VDD.n1880 0.152939
R16788 VDD.n1881 VDD.n1102 0.152939
R16789 VDD.n1895 VDD.n1102 0.152939
R16790 VDD.n1896 VDD.n1895 0.152939
R16791 VDD.n2209 VDD.n1896 0.152939
R16792 VDD.n3479 VDD.n3478 0.152939
R16793 VDD.n3480 VDD.n3479 0.152939
R16794 VDD.n3480 VDD.n489 0.152939
R16795 VDD.n3488 VDD.n489 0.152939
R16796 VDD.n3489 VDD.n3488 0.152939
R16797 VDD.n3490 VDD.n3489 0.152939
R16798 VDD.n3490 VDD.n485 0.152939
R16799 VDD.n3498 VDD.n485 0.152939
R16800 VDD.n3499 VDD.n3498 0.152939
R16801 VDD.n3500 VDD.n3499 0.152939
R16802 VDD.n3500 VDD.n479 0.152939
R16803 VDD.n3508 VDD.n479 0.152939
R16804 VDD.n3509 VDD.n3508 0.152939
R16805 VDD.n3510 VDD.n3509 0.152939
R16806 VDD.n3510 VDD.n475 0.152939
R16807 VDD.n3518 VDD.n475 0.152939
R16808 VDD.n3519 VDD.n3518 0.152939
R16809 VDD.n3520 VDD.n3519 0.152939
R16810 VDD.n3520 VDD.n471 0.152939
R16811 VDD.n3531 VDD.n471 0.152939
R16812 VDD.n3532 VDD.n3531 0.152939
R16813 VDD.n3533 VDD.n3532 0.152939
R16814 VDD.n3533 VDD.n467 0.152939
R16815 VDD.n3541 VDD.n467 0.152939
R16816 VDD.n3542 VDD.n3541 0.152939
R16817 VDD.n3543 VDD.n3542 0.152939
R16818 VDD.n3543 VDD.n463 0.152939
R16819 VDD.n3553 VDD.n463 0.152939
R16820 VDD.n3554 VDD.n3553 0.152939
R16821 VDD.n3555 VDD.n3554 0.152939
R16822 VDD.n3555 VDD.n457 0.152939
R16823 VDD.n3462 VDD.n446 0.152939
R16824 VDD.n3462 VDD.n3461 0.152939
R16825 VDD.n3584 VDD.n3583 0.152939
R16826 VDD.n3585 VDD.n3584 0.152939
R16827 VDD.n3585 VDD.n434 0.152939
R16828 VDD.n3600 VDD.n434 0.152939
R16829 VDD.n3601 VDD.n3600 0.152939
R16830 VDD.n3602 VDD.n3601 0.152939
R16831 VDD.n3602 VDD.n423 0.152939
R16832 VDD.n3616 VDD.n423 0.152939
R16833 VDD.n3617 VDD.n3616 0.152939
R16834 VDD.n3618 VDD.n3617 0.152939
R16835 VDD.n3618 VDD.n411 0.152939
R16836 VDD.n3632 VDD.n411 0.152939
R16837 VDD.n3633 VDD.n3632 0.152939
R16838 VDD.n3634 VDD.n3633 0.152939
R16839 VDD.n3634 VDD.n399 0.152939
R16840 VDD.n3648 VDD.n399 0.152939
R16841 VDD.n3649 VDD.n3648 0.152939
R16842 VDD.n3650 VDD.n3649 0.152939
R16843 VDD.n3650 VDD.n387 0.152939
R16844 VDD.n3664 VDD.n387 0.152939
R16845 VDD.n3665 VDD.n3664 0.152939
R16846 VDD.n3666 VDD.n3665 0.152939
R16847 VDD.n3666 VDD.n375 0.152939
R16848 VDD.n3680 VDD.n375 0.152939
R16849 VDD.n3681 VDD.n3680 0.152939
R16850 VDD.n3682 VDD.n3681 0.152939
R16851 VDD.n3682 VDD.n363 0.152939
R16852 VDD.n3697 VDD.n363 0.152939
R16853 VDD.n3698 VDD.n3697 0.152939
R16854 VDD.n3699 VDD.n3698 0.152939
R16855 VDD.n3699 VDD.n352 0.152939
R16856 VDD.n3716 VDD.n352 0.152939
R16857 VDD.n3717 VDD.n3716 0.152939
R16858 VDD.n3718 VDD.n3717 0.152939
R16859 VDD.n3718 VDD.n145 0.152939
R16860 VDD.n3953 VDD.n146 0.152939
R16861 VDD.n157 VDD.n146 0.152939
R16862 VDD.n158 VDD.n157 0.152939
R16863 VDD.n159 VDD.n158 0.152939
R16864 VDD.n167 VDD.n159 0.152939
R16865 VDD.n168 VDD.n167 0.152939
R16866 VDD.n169 VDD.n168 0.152939
R16867 VDD.n170 VDD.n169 0.152939
R16868 VDD.n178 VDD.n170 0.152939
R16869 VDD.n179 VDD.n178 0.152939
R16870 VDD.n180 VDD.n179 0.152939
R16871 VDD.n181 VDD.n180 0.152939
R16872 VDD.n189 VDD.n181 0.152939
R16873 VDD.n190 VDD.n189 0.152939
R16874 VDD.n191 VDD.n190 0.152939
R16875 VDD.n192 VDD.n191 0.152939
R16876 VDD.n200 VDD.n192 0.152939
R16877 VDD.n201 VDD.n200 0.152939
R16878 VDD.n202 VDD.n201 0.152939
R16879 VDD.n203 VDD.n202 0.152939
R16880 VDD.n211 VDD.n203 0.152939
R16881 VDD.n212 VDD.n211 0.152939
R16882 VDD.n213 VDD.n212 0.152939
R16883 VDD.n214 VDD.n213 0.152939
R16884 VDD.n222 VDD.n214 0.152939
R16885 VDD.n223 VDD.n222 0.152939
R16886 VDD.n224 VDD.n223 0.152939
R16887 VDD.n225 VDD.n224 0.152939
R16888 VDD.n233 VDD.n225 0.152939
R16889 VDD.n234 VDD.n233 0.152939
R16890 VDD.n235 VDD.n234 0.152939
R16891 VDD.n236 VDD.n235 0.152939
R16892 VDD.n244 VDD.n236 0.152939
R16893 VDD.n245 VDD.n244 0.152939
R16894 VDD.n3880 VDD.n245 0.152939
R16895 VDD.n3879 VDD.n246 0.152939
R16896 VDD.n251 VDD.n246 0.152939
R16897 VDD.n252 VDD.n251 0.152939
R16898 VDD.n253 VDD.n252 0.152939
R16899 VDD.n254 VDD.n253 0.152939
R16900 VDD.n261 VDD.n254 0.152939
R16901 VDD.n3863 VDD.n261 0.152939
R16902 VDD.n3863 VDD.n3862 0.152939
R16903 VDD.n3862 VDD.n3861 0.152939
R16904 VDD.n3861 VDD.n262 0.152939
R16905 VDD.n266 VDD.n262 0.152939
R16906 VDD.n267 VDD.n266 0.152939
R16907 VDD.n268 VDD.n267 0.152939
R16908 VDD.n272 VDD.n268 0.152939
R16909 VDD.n273 VDD.n272 0.152939
R16910 VDD.n3846 VDD.n273 0.152939
R16911 VDD.n3846 VDD.n3845 0.152939
R16912 VDD.n3845 VDD.n3844 0.152939
R16913 VDD.n3844 VDD.n277 0.152939
R16914 VDD.n283 VDD.n277 0.152939
R16915 VDD.n284 VDD.n283 0.152939
R16916 VDD.n285 VDD.n284 0.152939
R16917 VDD.n286 VDD.n285 0.152939
R16918 VDD.n290 VDD.n286 0.152939
R16919 VDD.n291 VDD.n290 0.152939
R16920 VDD.n292 VDD.n291 0.152939
R16921 VDD.n293 VDD.n292 0.152939
R16922 VDD.n297 VDD.n293 0.152939
R16923 VDD.n298 VDD.n297 0.152939
R16924 VDD.n299 VDD.n298 0.152939
R16925 VDD.n300 VDD.n299 0.152939
R16926 VDD.n304 VDD.n300 0.152939
R16927 VDD.n305 VDD.n304 0.152939
R16928 VDD.n306 VDD.n305 0.152939
R16929 VDD.n3809 VDD.n306 0.152939
R16930 VDD.n3809 VDD.n3808 0.152939
R16931 VDD.n3808 VDD.n3807 0.152939
R16932 VDD.n3807 VDD.n312 0.152939
R16933 VDD.n317 VDD.n312 0.152939
R16934 VDD.n318 VDD.n317 0.152939
R16935 VDD.n319 VDD.n318 0.152939
R16936 VDD.n323 VDD.n319 0.152939
R16937 VDD.n324 VDD.n323 0.152939
R16938 VDD.n325 VDD.n324 0.152939
R16939 VDD.n326 VDD.n325 0.152939
R16940 VDD.n3577 VDD.n440 0.152939
R16941 VDD.n3591 VDD.n440 0.152939
R16942 VDD.n3592 VDD.n3591 0.152939
R16943 VDD.n3593 VDD.n3592 0.152939
R16944 VDD.n3593 VDD.n429 0.152939
R16945 VDD.n3608 VDD.n429 0.152939
R16946 VDD.n3609 VDD.n3608 0.152939
R16947 VDD.n3610 VDD.n3609 0.152939
R16948 VDD.n3610 VDD.n417 0.152939
R16949 VDD.n3624 VDD.n417 0.152939
R16950 VDD.n3625 VDD.n3624 0.152939
R16951 VDD.n3626 VDD.n3625 0.152939
R16952 VDD.n3626 VDD.n405 0.152939
R16953 VDD.n3640 VDD.n405 0.152939
R16954 VDD.n3641 VDD.n3640 0.152939
R16955 VDD.n3642 VDD.n3641 0.152939
R16956 VDD.n3642 VDD.n393 0.152939
R16957 VDD.n3656 VDD.n393 0.152939
R16958 VDD.n3657 VDD.n3656 0.152939
R16959 VDD.n3658 VDD.n3657 0.152939
R16960 VDD.n3658 VDD.n381 0.152939
R16961 VDD.n3672 VDD.n381 0.152939
R16962 VDD.n3673 VDD.n3672 0.152939
R16963 VDD.n3674 VDD.n3673 0.152939
R16964 VDD.n3674 VDD.n369 0.152939
R16965 VDD.n3688 VDD.n369 0.152939
R16966 VDD.n3689 VDD.n3688 0.152939
R16967 VDD.n3690 VDD.n3689 0.152939
R16968 VDD.n3690 VDD.n358 0.152939
R16969 VDD.n3705 VDD.n358 0.152939
R16970 VDD.n3706 VDD.n3705 0.152939
R16971 VDD.n3707 VDD.n3706 0.152939
R16972 VDD.n3709 VDD.n3707 0.152939
R16973 VDD.n3709 VDD.n3708 0.152939
R16974 VDD.n3708 VDD.n347 0.152939
R16975 VDD.n347 VDD.n345 0.152939
R16976 VDD.n3727 VDD.n345 0.152939
R16977 VDD.n3728 VDD.n3727 0.152939
R16978 VDD.n3729 VDD.n3728 0.152939
R16979 VDD.n3729 VDD.n343 0.152939
R16980 VDD.n3734 VDD.n343 0.152939
R16981 VDD.n3735 VDD.n3734 0.152939
R16982 VDD.n3736 VDD.n3735 0.152939
R16983 VDD.n3736 VDD.n341 0.152939
R16984 VDD.n3741 VDD.n341 0.152939
R16985 VDD.n3742 VDD.n3741 0.152939
R16986 VDD.n3743 VDD.n3742 0.152939
R16987 VDD.n3743 VDD.n339 0.152939
R16988 VDD.n3748 VDD.n339 0.152939
R16989 VDD.n3749 VDD.n3748 0.152939
R16990 VDD.n3750 VDD.n3749 0.152939
R16991 VDD.n3750 VDD.n337 0.152939
R16992 VDD.n3755 VDD.n337 0.152939
R16993 VDD.n3756 VDD.n3755 0.152939
R16994 VDD.n3757 VDD.n3756 0.152939
R16995 VDD.n3757 VDD.n335 0.152939
R16996 VDD.n3762 VDD.n335 0.152939
R16997 VDD.n3763 VDD.n3762 0.152939
R16998 VDD.n3764 VDD.n3763 0.152939
R16999 VDD.n3764 VDD.n333 0.152939
R17000 VDD.n3769 VDD.n333 0.152939
R17001 VDD.n3770 VDD.n3769 0.152939
R17002 VDD.n3771 VDD.n3770 0.152939
R17003 VDD.n3771 VDD.n331 0.152939
R17004 VDD.n3776 VDD.n331 0.152939
R17005 VDD.n3777 VDD.n3776 0.152939
R17006 VDD.n3778 VDD.n3777 0.152939
R17007 VDD.n3778 VDD.n329 0.152939
R17008 VDD.n3783 VDD.n329 0.152939
R17009 VDD.n3784 VDD.n3783 0.152939
R17010 VDD.n3785 VDD.n3784 0.152939
R17011 VDD.n458 VDD.n450 0.152939
R17012 VDD.n3576 VDD.n450 0.152939
R17013 VDD.n2223 VDD.n1088 0.152939
R17014 VDD.n2216 VDD.n1088 0.152939
R17015 VDD.n1485 VDD.n1484 0.152939
R17016 VDD.n1485 VDD.n1299 0.152939
R17017 VDD.n1499 VDD.n1299 0.152939
R17018 VDD.n1500 VDD.n1499 0.152939
R17019 VDD.n1501 VDD.n1500 0.152939
R17020 VDD.n1501 VDD.n1287 0.152939
R17021 VDD.n1515 VDD.n1287 0.152939
R17022 VDD.n1516 VDD.n1515 0.152939
R17023 VDD.n1517 VDD.n1516 0.152939
R17024 VDD.n1517 VDD.n1275 0.152939
R17025 VDD.n1531 VDD.n1275 0.152939
R17026 VDD.n1532 VDD.n1531 0.152939
R17027 VDD.n1533 VDD.n1532 0.152939
R17028 VDD.n1533 VDD.n1263 0.152939
R17029 VDD.n1547 VDD.n1263 0.152939
R17030 VDD.n1548 VDD.n1547 0.152939
R17031 VDD.n1549 VDD.n1548 0.152939
R17032 VDD.n1549 VDD.n1252 0.152939
R17033 VDD.n1564 VDD.n1252 0.152939
R17034 VDD.n1565 VDD.n1564 0.152939
R17035 VDD.n1566 VDD.n1565 0.152939
R17036 VDD.n1566 VDD.n1240 0.152939
R17037 VDD.n1580 VDD.n1240 0.152939
R17038 VDD.n1581 VDD.n1580 0.152939
R17039 VDD.n1582 VDD.n1581 0.152939
R17040 VDD.n1582 VDD.n1228 0.152939
R17041 VDD.n1596 VDD.n1228 0.152939
R17042 VDD.n1597 VDD.n1596 0.152939
R17043 VDD.n1598 VDD.n1597 0.152939
R17044 VDD.n1598 VDD.n1216 0.152939
R17045 VDD.n1612 VDD.n1216 0.152939
R17046 VDD.n1613 VDD.n1612 0.152939
R17047 VDD.n1614 VDD.n1613 0.152939
R17048 VDD.n1614 VDD.n1204 0.152939
R17049 VDD.n1759 VDD.n1204 0.152939
R17050 VDD.n1760 VDD.n1759 0.152939
R17051 VDD.n1761 VDD.n1760 0.152939
R17052 VDD.n1761 VDD.n1192 0.152939
R17053 VDD.n1775 VDD.n1192 0.152939
R17054 VDD.n1776 VDD.n1775 0.152939
R17055 VDD.n1777 VDD.n1776 0.152939
R17056 VDD.n1777 VDD.n1180 0.152939
R17057 VDD.n1791 VDD.n1180 0.152939
R17058 VDD.n1792 VDD.n1791 0.152939
R17059 VDD.n1793 VDD.n1792 0.152939
R17060 VDD.n1793 VDD.n1168 0.152939
R17061 VDD.n1807 VDD.n1168 0.152939
R17062 VDD.n1808 VDD.n1807 0.152939
R17063 VDD.n1809 VDD.n1808 0.152939
R17064 VDD.n1809 VDD.n1155 0.152939
R17065 VDD.n1823 VDD.n1155 0.152939
R17066 VDD.n1824 VDD.n1823 0.152939
R17067 VDD.n1825 VDD.n1824 0.152939
R17068 VDD.n1825 VDD.n1144 0.152939
R17069 VDD.n1839 VDD.n1144 0.152939
R17070 VDD.n1840 VDD.n1839 0.152939
R17071 VDD.n1841 VDD.n1840 0.152939
R17072 VDD.n1841 VDD.n1132 0.152939
R17073 VDD.n1855 VDD.n1132 0.152939
R17074 VDD.n1856 VDD.n1855 0.152939
R17075 VDD.n1857 VDD.n1856 0.152939
R17076 VDD.n1857 VDD.n1120 0.152939
R17077 VDD.n1871 VDD.n1120 0.152939
R17078 VDD.n1872 VDD.n1871 0.152939
R17079 VDD.n1873 VDD.n1872 0.152939
R17080 VDD.n1873 VDD.n1108 0.152939
R17081 VDD.n1887 VDD.n1108 0.152939
R17082 VDD.n1888 VDD.n1887 0.152939
R17083 VDD.n1889 VDD.n1888 0.152939
R17084 VDD.n1889 VDD.n1093 0.152939
R17085 VDD.n2215 VDD.n1093 0.152939
R17086 VDD.n1475 VDD.n1339 0.152939
R17087 VDD.n1475 VDD.n1474 0.152939
R17088 VDD.n1474 VDD.n1473 0.152939
R17089 VDD.n1473 VDD.n1341 0.152939
R17090 VDD.n1469 VDD.n1341 0.152939
R17091 VDD.n1469 VDD.n1468 0.152939
R17092 VDD.n1468 VDD.n1467 0.152939
R17093 VDD.n1467 VDD.n1346 0.152939
R17094 VDD.n1459 VDD.n1346 0.152939
R17095 VDD.n1459 VDD.n1458 0.152939
R17096 VDD.n1458 VDD.n1457 0.152939
R17097 VDD.n1457 VDD.n1350 0.152939
R17098 VDD.n1453 VDD.n1350 0.152939
R17099 VDD.n1453 VDD.n1452 0.152939
R17100 VDD.n1452 VDD.n1451 0.152939
R17101 VDD.n1451 VDD.n1356 0.152939
R17102 VDD.n1443 VDD.n1356 0.152939
R17103 VDD.n1443 VDD.n1442 0.152939
R17104 VDD.n1442 VDD.n1441 0.152939
R17105 VDD.n1441 VDD.n1360 0.152939
R17106 VDD.n1437 VDD.n1360 0.152939
R17107 VDD.n1437 VDD.n1436 0.152939
R17108 VDD.n1436 VDD.n1435 0.152939
R17109 VDD.n1435 VDD.n1366 0.152939
R17110 VDD.n1431 VDD.n1366 0.152939
R17111 VDD.n1431 VDD.n1430 0.152939
R17112 VDD.n1430 VDD.n1374 0.152939
R17113 VDD.n1426 VDD.n1374 0.152939
R17114 VDD.n1426 VDD.n1425 0.152939
R17115 VDD.n1425 VDD.n1424 0.152939
R17116 VDD.n1424 VDD.n1380 0.152939
R17117 VDD.n1420 VDD.n1380 0.152939
R17118 VDD.n1420 VDD.n1419 0.152939
R17119 VDD.n1419 VDD.n1418 0.152939
R17120 VDD.n1418 VDD.n1386 0.152939
R17121 VDD.n1411 VDD.n1386 0.152939
R17122 VDD.n1411 VDD.n1410 0.152939
R17123 VDD.n1410 VDD.n1409 0.152939
R17124 VDD.n1409 VDD.n1391 0.152939
R17125 VDD.n1405 VDD.n1391 0.152939
R17126 VDD.n1405 VDD.n1404 0.152939
R17127 VDD.n1404 VDD.n1403 0.152939
R17128 VDD.n1403 VDD.n1397 0.152939
R17129 VDD.n1397 VDD.n1311 0.152939
R17130 VDD.n1483 VDD.n1311 0.152939
R17131 VDD.n1491 VDD.n1305 0.152939
R17132 VDD.n1492 VDD.n1491 0.152939
R17133 VDD.n1493 VDD.n1492 0.152939
R17134 VDD.n1493 VDD.n1293 0.152939
R17135 VDD.n1507 VDD.n1293 0.152939
R17136 VDD.n1508 VDD.n1507 0.152939
R17137 VDD.n1509 VDD.n1508 0.152939
R17138 VDD.n1509 VDD.n1281 0.152939
R17139 VDD.n1523 VDD.n1281 0.152939
R17140 VDD.n1524 VDD.n1523 0.152939
R17141 VDD.n1525 VDD.n1524 0.152939
R17142 VDD.n1525 VDD.n1269 0.152939
R17143 VDD.n1539 VDD.n1269 0.152939
R17144 VDD.n1540 VDD.n1539 0.152939
R17145 VDD.n1541 VDD.n1540 0.152939
R17146 VDD.n1541 VDD.n1257 0.152939
R17147 VDD.n1556 VDD.n1257 0.152939
R17148 VDD.n1557 VDD.n1556 0.152939
R17149 VDD.n1558 VDD.n1557 0.152939
R17150 VDD.n1558 VDD.n1246 0.152939
R17151 VDD.n1572 VDD.n1246 0.152939
R17152 VDD.n1573 VDD.n1572 0.152939
R17153 VDD.n1574 VDD.n1573 0.152939
R17154 VDD.n1574 VDD.n1234 0.152939
R17155 VDD.n1588 VDD.n1234 0.152939
R17156 VDD.n1589 VDD.n1588 0.152939
R17157 VDD.n1590 VDD.n1589 0.152939
R17158 VDD.n1590 VDD.n1222 0.152939
R17159 VDD.n1604 VDD.n1222 0.152939
R17160 VDD.n1605 VDD.n1604 0.152939
R17161 VDD.n1606 VDD.n1605 0.152939
R17162 VDD.n1606 VDD.n1210 0.152939
R17163 VDD.n1620 VDD.n1210 0.152939
R17164 VDD.n1621 VDD.n1620 0.152939
R17165 VDD.n1753 VDD.n1621 0.152939
R17166 VDD.n2199 VDD.n2198 0.128549
R17167 VDD.n3461 VDD.n3452 0.128549
R17168 VDD.n3564 VDD.n458 0.128549
R17169 VDD.n2224 VDD.n2223 0.128549
R17170 VDD.n1752 VDD.n1198 0.0695946
R17171 VDD.n3954 VDD.n145 0.0695946
R17172 VDD.n3954 VDD.n3953 0.0695946
R17173 VDD.n1753 VDD.n1752 0.0695946
R17174 VDD.n2199 VDD.n1902 0.0248902
R17175 VDD.n2224 VDD.n1085 0.0248902
R17176 VDD.n3478 VDD.n3452 0.0248902
R17177 VDD.n3564 VDD.n457 0.0248902
R17178 VDD VDD.n15 0.00833333
R17179 a_n6573_8708.n4 a_n6573_8708.n3 7.01317
R17180 a_n6573_8708.n17 a_n6573_8708.n3 4.70034
R17181 a_n6573_8708.n6 a_n6573_8708.n5 7.01317
R17182 a_n6573_8708.n16 a_n6573_8708.n5 4.70034
R17183 a_n6573_8708.n11 a_n6573_8708.n0 4.70026
R17184 a_n6573_8708.n20 a_n6573_8708.n0 4.70026
R17185 a_n6573_8708.n19 a_n6573_8708.n0 4.70026
R17186 a_n6573_8708.n18 a_n6573_8708.n0 4.70026
R17187 a_n6573_8708.n8 a_n6573_8708.n7 7.01317
R17188 a_n6573_8708.n15 a_n6573_8708.n7 4.70034
R17189 a_n6573_8708.n10 a_n6573_8708.n9 7.01317
R17190 a_n6573_8708.n9 a_n6573_8708.n14 4.70034
R17191 a_n6573_8708.n58 a_n6573_8708.t1 119.138
R17192 a_n6573_8708.t3 a_n6573_8708.n13 96.7557
R17193 a_n6573_8708.n12 a_n6573_8708.t7 93.6263
R17194 a_n6573_8708.n12 a_n6573_8708.t19 90.3822
R17195 a_n6573_8708.n58 a_n6573_8708.t0 87.4995
R17196 a_n6573_8708.n13 a_n6573_8708.t9 87.2529
R17197 a_n6573_8708.n13 a_n6573_8708.t5 87.2529
R17198 a_n6573_8708.n12 a_n6573_8708.t17 87.2529
R17199 a_n6573_8708.n0 a_n6573_8708.n33 3.92153
R17200 a_n6573_8708.n0 a_n6573_8708.n1 3.92152
R17201 a_n6573_8708.n0 a_n6573_8708.n31 3.92153
R17202 a_n6573_8708.n7 a_n6573_8708.n27 3.74957
R17203 a_n6573_8708.n5 a_n6573_8708.n25 3.74957
R17204 a_n6573_8708.n3 a_n6573_8708.n23 3.74957
R17205 a_n6573_8708.n39 a_n6573_8708.n10 72.3794
R17206 a_n6573_8708.n42 a_n6573_8708.n8 72.3794
R17207 a_n6573_8708.n37 a_n6573_8708.n6 72.3794
R17208 a_n6573_8708.n36 a_n6573_8708.n4 72.3794
R17209 a_n6573_8708.n39 a_n6573_8708.t8 37.246
R17210 a_n6573_8708.n29 a_n6573_8708.t4 69.3436
R17211 a_n6573_8708.n38 a_n6573_8708.t14 37.246
R17212 a_n6573_8708.n40 a_n6573_8708.t20 37.246
R17213 a_n6573_8708.n30 a_n6573_8708.t2 69.3438
R17214 a_n6573_8708.n42 a_n6573_8708.t23 37.246
R17215 a_n6573_8708.n27 a_n6573_8708.t30 69.3436
R17216 a_n6573_8708.n41 a_n6573_8708.t34 37.246
R17217 a_n6573_8708.n43 a_n6573_8708.t41 37.246
R17218 a_n6573_8708.n28 a_n6573_8708.t29 69.3438
R17219 a_n6573_8708.n37 a_n6573_8708.t16 37.246
R17220 a_n6573_8708.n25 a_n6573_8708.t18 69.3436
R17221 a_n6573_8708.n45 a_n6573_8708.t10 37.246
R17222 a_n6573_8708.n44 a_n6573_8708.t12 37.246
R17223 a_n6573_8708.n26 a_n6573_8708.t6 69.3438
R17224 a_n6573_8708.n36 a_n6573_8708.t33 37.246
R17225 a_n6573_8708.n23 a_n6573_8708.t35 69.3436
R17226 a_n6573_8708.n47 a_n6573_8708.t43 37.246
R17227 a_n6573_8708.n46 a_n6573_8708.t40 37.246
R17228 a_n6573_8708.n24 a_n6573_8708.t46 69.3438
R17229 a_n6573_8708.n2 a_n6573_8708.t36 68.7679
R17230 a_n6573_8708.n56 a_n6573_8708.t24 37.246
R17231 a_n6573_8708.n49 a_n6573_8708.t28 37.246
R17232 a_n6573_8708.n34 a_n6573_8708.t22 68.7676
R17233 a_n6573_8708.n21 a_n6573_8708.t26 68.7679
R17234 a_n6573_8708.n55 a_n6573_8708.t38 37.246
R17235 a_n6573_8708.n50 a_n6573_8708.t25 37.246
R17236 a_n6573_8708.n33 a_n6573_8708.t45 68.7676
R17237 a_n6573_8708.n1 a_n6573_8708.t37 68.7679
R17238 a_n6573_8708.n54 a_n6573_8708.t42 37.246
R17239 a_n6573_8708.n51 a_n6573_8708.t44 37.246
R17240 a_n6573_8708.n32 a_n6573_8708.t31 68.7676
R17241 a_n6573_8708.n22 a_n6573_8708.t39 68.7679
R17242 a_n6573_8708.n53 a_n6573_8708.t32 37.246
R17243 a_n6573_8708.n52 a_n6573_8708.t47 37.246
R17244 a_n6573_8708.n31 a_n6573_8708.t27 68.7676
R17245 a_n6573_8708.n9 a_n6573_8708.n58 24.7041
R17246 a_n6573_8708.n29 a_n6573_8708.n38 68.505
R17247 a_n6573_8708.n14 a_n6573_8708.n39 48.5071
R17248 a_n6573_8708.n10 a_n6573_8708.n40 52.7921
R17249 a_n6573_8708.n27 a_n6573_8708.n41 68.505
R17250 a_n6573_8708.n41 a_n6573_8708.n15 54.9002
R17251 a_n6573_8708.n15 a_n6573_8708.n42 48.5071
R17252 a_n6573_8708.n8 a_n6573_8708.n43 52.7921
R17253 a_n6573_8708.n45 a_n6573_8708.n25 68.505
R17254 a_n6573_8708.n45 a_n6573_8708.n16 54.9002
R17255 a_n6573_8708.n16 a_n6573_8708.n37 48.5071
R17256 a_n6573_8708.n44 a_n6573_8708.n6 52.7921
R17257 a_n6573_8708.n47 a_n6573_8708.n23 68.505
R17258 a_n6573_8708.n47 a_n6573_8708.n17 54.9002
R17259 a_n6573_8708.n17 a_n6573_8708.n36 48.5071
R17260 a_n6573_8708.n46 a_n6573_8708.n4 52.7921
R17261 a_n6573_8708.n56 a_n6573_8708.n2 71.7742
R17262 a_n6573_8708.n18 a_n6573_8708.n56 51.7038
R17263 a_n6573_8708.n55 a_n6573_8708.n21 71.7742
R17264 a_n6573_8708.n19 a_n6573_8708.n55 51.7038
R17265 a_n6573_8708.n51 a_n6573_8708.n20 51.7034
R17266 a_n6573_8708.n52 a_n6573_8708.n11 51.7034
R17267 a_n6573_8708.n34 a_n6573_8708.n49 71.7745
R17268 a_n6573_8708.n33 a_n6573_8708.n50 71.7745
R17269 a_n6573_8708.n1 a_n6573_8708.n54 71.7742
R17270 a_n6573_8708.n32 a_n6573_8708.n51 71.7745
R17271 a_n6573_8708.n22 a_n6573_8708.n53 71.7742
R17272 a_n6573_8708.n31 a_n6573_8708.n52 71.7745
R17273 a_n6573_8708.n30 a_n6573_8708.n40 68.5052
R17274 a_n6573_8708.n28 a_n6573_8708.n43 68.5052
R17275 a_n6573_8708.n26 a_n6573_8708.n44 68.5052
R17276 a_n6573_8708.n24 a_n6573_8708.n46 68.5052
R17277 a_n6573_8708.n7 a_n6573_8708.n57 12.983
R17278 a_n6573_8708.n3 a_n6573_8708.n35 12.9678
R17279 a_n6573_8708.n35 a_n6573_8708.n9 11.9546
R17280 a_n6573_8708.n48 a_n6573_8708.n5 9.64965
R17281 a_n6573_8708.n57 a_n6573_8708.n0 6.83904
R17282 a_n6573_8708.n5 a_n6573_8708.n3 6.56773
R17283 a_n6573_8708.n14 a_n6573_8708.n38 54.9002
R17284 a_n6573_8708.t9 a_n6573_8708.t21 6.37403
R17285 a_n6573_8708.t5 a_n6573_8708.t15 6.37403
R17286 a_n6573_8708.t17 a_n6573_8708.t13 6.37403
R17287 a_n6573_8708.t19 a_n6573_8708.t11 6.37403
R17288 a_n6573_8708.n9 a_n6573_8708.n7 4.15343
R17289 a_n6573_8708.n57 a_n6573_8708.n48 3.31868
R17290 a_n6573_8708.n18 a_n6573_8708.n49 51.7034
R17291 a_n6573_8708.n19 a_n6573_8708.n50 51.7034
R17292 a_n6573_8708.n54 a_n6573_8708.n20 51.7038
R17293 a_n6573_8708.n53 a_n6573_8708.n11 51.7038
R17294 a_n6573_8708.n48 a_n6573_8708.n12 15.2899
R17295 a_n6573_8708.n13 a_n6573_8708.n35 14.5522
R17296 a_n6573_8708.n0 a_n6573_8708.n32 10.1331
R17297 a_n6573_8708.n2 a_n6573_8708.n0 10.1331
R17298 a_n6573_8708.n7 a_n6573_8708.n28 9.76123
R17299 a_n6573_8708.n5 a_n6573_8708.n26 9.76123
R17300 a_n6573_8708.n3 a_n6573_8708.n24 9.76123
R17301 a_n6573_8708.n9 a_n6573_8708.n30 9.13177
R17302 a_n6573_8708.n0 a_n6573_8708.n22 8.60751
R17303 a_n6573_8708.n21 a_n6573_8708.n0 8.40372
R17304 a_n6573_8708.n0 a_n6573_8708.n35 7.86745
R17305 a_n6573_8708.n9 a_n6573_8708.n29 6.75544
R17306 a_n6573_8708.n0 a_n6573_8708.n34 6.54862
R17307 a_n6651_8904.n1 a_n6651_8904.t12 113.434
R17308 a_n6651_8904.n3 a_n6651_8904.t13 111.385
R17309 a_n6651_8904.n1 a_n6651_8904.n0 103.931
R17310 a_n6651_8904.n5 a_n6651_8904.n4 103.931
R17311 a_n6651_8904.n3 a_n6651_8904.n2 103.931
R17312 a_n6651_8904.n15 a_n6651_8904.n14 103.931
R17313 a_n6651_8904.n7 a_n6651_8904.t4 96.7557
R17314 a_n6651_8904.n12 a_n6651_8904.t7 93.6264
R17315 a_n6651_8904.n9 a_n6651_8904.t2 93.6264
R17316 a_n6651_8904.n8 a_n6651_8904.t0 93.6264
R17317 a_n6651_8904.n11 a_n6651_8904.n10 87.2529
R17318 a_n6651_8904.n7 a_n6651_8904.n6 87.2529
R17319 a_n6651_8904.n13 a_n6651_8904.n5 28.0067
R17320 a_n6651_8904.n14 a_n6651_8904.n13 15.2087
R17321 a_n6651_8904.n13 a_n6651_8904.n12 7.04576
R17322 a_n6651_8904.n0 a_n6651_8904.t9 6.37403
R17323 a_n6651_8904.n0 a_n6651_8904.t11 6.37403
R17324 a_n6651_8904.n10 a_n6651_8904.t6 6.37403
R17325 a_n6651_8904.n10 a_n6651_8904.t3 6.37403
R17326 a_n6651_8904.n6 a_n6651_8904.t1 6.37403
R17327 a_n6651_8904.n6 a_n6651_8904.t5 6.37403
R17328 a_n6651_8904.n4 a_n6651_8904.t8 6.37403
R17329 a_n6651_8904.n4 a_n6651_8904.t17 6.37403
R17330 a_n6651_8904.n2 a_n6651_8904.t10 6.37403
R17331 a_n6651_8904.n2 a_n6651_8904.t15 6.37403
R17332 a_n6651_8904.t16 a_n6651_8904.n15 6.37403
R17333 a_n6651_8904.n15 a_n6651_8904.t14 6.37403
R17334 a_n6651_8904.n8 a_n6651_8904.n7 3.12981
R17335 a_n6651_8904.n11 a_n6651_8904.n9 3.12981
R17336 a_n6651_8904.n12 a_n6651_8904.n11 3.12981
R17337 a_n6651_8904.n14 a_n6651_8904.n1 3.12981
R17338 a_n6651_8904.n5 a_n6651_8904.n3 1.08086
R17339 a_n6651_8904.n9 a_n6651_8904.n8 0.806535
R17340 a_n5180_7124.n6 a_n5180_7124.t7 96.7557
R17341 a_n5180_7124.t17 a_n5180_7124.n16 96.7557
R17342 a_n5180_7124.n1 a_n5180_7124.t9 96.7556
R17343 a_n5180_7124.n7 a_n5180_7124.t5 93.6264
R17344 a_n5180_7124.n8 a_n5180_7124.t8 93.6264
R17345 a_n5180_7124.n11 a_n5180_7124.t4 93.6264
R17346 a_n5180_7124.n16 a_n5180_7124.n15 87.2529
R17347 a_n5180_7124.n14 a_n5180_7124.n13 87.2529
R17348 a_n5180_7124.n1 a_n5180_7124.n0 87.2529
R17349 a_n5180_7124.n3 a_n5180_7124.n2 87.2529
R17350 a_n5180_7124.n6 a_n5180_7124.n5 87.2529
R17351 a_n5180_7124.n10 a_n5180_7124.n9 87.2529
R17352 a_n5180_7124.n14 a_n5180_7124.n12 38.4152
R17353 a_n5180_7124.n4 a_n5180_7124.n3 11.7807
R17354 a_n5180_7124.n4 a_n5180_7124.t0 9.86523
R17355 a_n5180_7124.n12 a_n5180_7124.n11 7.04576
R17356 a_n5180_7124.n15 a_n5180_7124.t18 6.37403
R17357 a_n5180_7124.n15 a_n5180_7124.t11 6.37403
R17358 a_n5180_7124.n13 a_n5180_7124.t16 6.37403
R17359 a_n5180_7124.n13 a_n5180_7124.t14 6.37403
R17360 a_n5180_7124.n0 a_n5180_7124.t15 6.37403
R17361 a_n5180_7124.n0 a_n5180_7124.t12 6.37403
R17362 a_n5180_7124.n2 a_n5180_7124.t13 6.37403
R17363 a_n5180_7124.n2 a_n5180_7124.t10 6.37403
R17364 a_n5180_7124.n5 a_n5180_7124.t3 6.37403
R17365 a_n5180_7124.n5 a_n5180_7124.t2 6.37403
R17366 a_n5180_7124.n9 a_n5180_7124.t6 6.37403
R17367 a_n5180_7124.n9 a_n5180_7124.t1 6.37403
R17368 a_n5180_7124.n12 a_n5180_7124.n4 3.31868
R17369 a_n5180_7124.n3 a_n5180_7124.n1 3.12981
R17370 a_n5180_7124.n11 a_n5180_7124.n10 3.12981
R17371 a_n5180_7124.n10 a_n5180_7124.n8 3.12981
R17372 a_n5180_7124.n7 a_n5180_7124.n6 3.12981
R17373 a_n5180_7124.n16 a_n5180_7124.n14 3.12981
R17374 a_n5180_7124.n8 a_n5180_7124.n7 0.806535
R17375 VN.n2 VN.t1 243.97
R17376 VN.n5 VN.t0 243.255
R17377 VN.n2 VN.n1 223.454
R17378 VN.n4 VN.n3 223.454
R17379 VN.n0 VN.t7 86.9589
R17380 VN.n0 VN.t6 70.3441
R17381 VN.n1 VN.t2 19.8005
R17382 VN.n1 VN.t4 19.8005
R17383 VN.n3 VN.t3 19.8005
R17384 VN.n3 VN.t5 19.8005
R17385 VN VN.n6 16.5269
R17386 VN.n6 VN.n5 5.04791
R17387 VN.n6 VN.n0 1.188
R17388 VN.n5 VN.n4 0.716017
R17389 VN.n4 VN.n2 0.716017
R17390 DIFFPAIR_BIAS.n14 DIFFPAIR_BIAS.n0 289.615
R17391 DIFFPAIR_BIAS.n33 DIFFPAIR_BIAS.n19 289.615
R17392 DIFFPAIR_BIAS.n53 DIFFPAIR_BIAS.n39 289.615
R17393 DIFFPAIR_BIAS.n15 DIFFPAIR_BIAS.n14 185
R17394 DIFFPAIR_BIAS.n13 DIFFPAIR_BIAS.n12 185
R17395 DIFFPAIR_BIAS.n4 DIFFPAIR_BIAS.n3 185
R17396 DIFFPAIR_BIAS.n7 DIFFPAIR_BIAS.n6 185
R17397 DIFFPAIR_BIAS.n34 DIFFPAIR_BIAS.n33 185
R17398 DIFFPAIR_BIAS.n32 DIFFPAIR_BIAS.n31 185
R17399 DIFFPAIR_BIAS.n23 DIFFPAIR_BIAS.n22 185
R17400 DIFFPAIR_BIAS.n26 DIFFPAIR_BIAS.n25 185
R17401 DIFFPAIR_BIAS.n54 DIFFPAIR_BIAS.n53 185
R17402 DIFFPAIR_BIAS.n52 DIFFPAIR_BIAS.n51 185
R17403 DIFFPAIR_BIAS.n43 DIFFPAIR_BIAS.n42 185
R17404 DIFFPAIR_BIAS.n46 DIFFPAIR_BIAS.n45 185
R17405 DIFFPAIR_BIAS.t3 DIFFPAIR_BIAS.n5 147.888
R17406 DIFFPAIR_BIAS.t5 DIFFPAIR_BIAS.n24 147.888
R17407 DIFFPAIR_BIAS.t1 DIFFPAIR_BIAS.n44 147.888
R17408 DIFFPAIR_BIAS.n64 DIFFPAIR_BIAS.t6 142.5
R17409 DIFFPAIR_BIAS.n63 DIFFPAIR_BIAS.t7 141.083
R17410 DIFFPAIR_BIAS.n62 DIFFPAIR_BIAS.t8 141.083
R17411 DIFFPAIR_BIAS.n14 DIFFPAIR_BIAS.n13 104.615
R17412 DIFFPAIR_BIAS.n13 DIFFPAIR_BIAS.n3 104.615
R17413 DIFFPAIR_BIAS.n6 DIFFPAIR_BIAS.n3 104.615
R17414 DIFFPAIR_BIAS.n33 DIFFPAIR_BIAS.n32 104.615
R17415 DIFFPAIR_BIAS.n32 DIFFPAIR_BIAS.n22 104.615
R17416 DIFFPAIR_BIAS.n25 DIFFPAIR_BIAS.n22 104.615
R17417 DIFFPAIR_BIAS.n53 DIFFPAIR_BIAS.n52 104.615
R17418 DIFFPAIR_BIAS.n52 DIFFPAIR_BIAS.n42 104.615
R17419 DIFFPAIR_BIAS.n45 DIFFPAIR_BIAS.n42 104.615
R17420 DIFFPAIR_BIAS.n59 DIFFPAIR_BIAS.t2 102.475
R17421 DIFFPAIR_BIAS.n59 DIFFPAIR_BIAS.t4 100.391
R17422 DIFFPAIR_BIAS.n60 DIFFPAIR_BIAS.t0 100.391
R17423 DIFFPAIR_BIAS.n38 DIFFPAIR_BIAS.n18 74.4516
R17424 DIFFPAIR_BIAS.n38 DIFFPAIR_BIAS.n37 72.3702
R17425 DIFFPAIR_BIAS.n58 DIFFPAIR_BIAS.n57 72.3702
R17426 DIFFPAIR_BIAS.n6 DIFFPAIR_BIAS.t3 52.3082
R17427 DIFFPAIR_BIAS.n25 DIFFPAIR_BIAS.t5 52.3082
R17428 DIFFPAIR_BIAS.n45 DIFFPAIR_BIAS.t1 52.3082
R17429 DIFFPAIR_BIAS.n7 DIFFPAIR_BIAS.n5 15.6496
R17430 DIFFPAIR_BIAS.n26 DIFFPAIR_BIAS.n24 15.6496
R17431 DIFFPAIR_BIAS.n46 DIFFPAIR_BIAS.n44 15.6496
R17432 DIFFPAIR_BIAS.n8 DIFFPAIR_BIAS.n4 12.8005
R17433 DIFFPAIR_BIAS.n27 DIFFPAIR_BIAS.n23 12.8005
R17434 DIFFPAIR_BIAS.n47 DIFFPAIR_BIAS.n43 12.8005
R17435 DIFFPAIR_BIAS.n12 DIFFPAIR_BIAS.n11 12.0247
R17436 DIFFPAIR_BIAS.n31 DIFFPAIR_BIAS.n30 12.0247
R17437 DIFFPAIR_BIAS.n51 DIFFPAIR_BIAS.n50 12.0247
R17438 DIFFPAIR_BIAS.n15 DIFFPAIR_BIAS.n2 11.249
R17439 DIFFPAIR_BIAS.n34 DIFFPAIR_BIAS.n21 11.249
R17440 DIFFPAIR_BIAS.n54 DIFFPAIR_BIAS.n41 11.249
R17441 DIFFPAIR_BIAS.n16 DIFFPAIR_BIAS.n0 10.4732
R17442 DIFFPAIR_BIAS.n35 DIFFPAIR_BIAS.n19 10.4732
R17443 DIFFPAIR_BIAS.n55 DIFFPAIR_BIAS.n39 10.4732
R17444 DIFFPAIR_BIAS.n18 DIFFPAIR_BIAS.n17 9.45567
R17445 DIFFPAIR_BIAS.n37 DIFFPAIR_BIAS.n36 9.45567
R17446 DIFFPAIR_BIAS.n57 DIFFPAIR_BIAS.n56 9.45567
R17447 DIFFPAIR_BIAS.n17 DIFFPAIR_BIAS.n16 9.3005
R17448 DIFFPAIR_BIAS.n2 DIFFPAIR_BIAS.n1 9.3005
R17449 DIFFPAIR_BIAS.n11 DIFFPAIR_BIAS.n10 9.3005
R17450 DIFFPAIR_BIAS.n9 DIFFPAIR_BIAS.n8 9.3005
R17451 DIFFPAIR_BIAS.n36 DIFFPAIR_BIAS.n35 9.3005
R17452 DIFFPAIR_BIAS.n21 DIFFPAIR_BIAS.n20 9.3005
R17453 DIFFPAIR_BIAS.n30 DIFFPAIR_BIAS.n29 9.3005
R17454 DIFFPAIR_BIAS.n28 DIFFPAIR_BIAS.n27 9.3005
R17455 DIFFPAIR_BIAS.n56 DIFFPAIR_BIAS.n55 9.3005
R17456 DIFFPAIR_BIAS.n41 DIFFPAIR_BIAS.n40 9.3005
R17457 DIFFPAIR_BIAS.n50 DIFFPAIR_BIAS.n49 9.3005
R17458 DIFFPAIR_BIAS.n48 DIFFPAIR_BIAS.n47 9.3005
R17459 DIFFPAIR_BIAS.n61 DIFFPAIR_BIAS.n60 5.3272
R17460 DIFFPAIR_BIAS.n61 DIFFPAIR_BIAS.n58 5.13582
R17461 DIFFPAIR_BIAS.n9 DIFFPAIR_BIAS.n5 4.40546
R17462 DIFFPAIR_BIAS.n28 DIFFPAIR_BIAS.n24 4.40546
R17463 DIFFPAIR_BIAS.n48 DIFFPAIR_BIAS.n44 4.40546
R17464 DIFFPAIR_BIAS.n62 DIFFPAIR_BIAS.n61 4.32378
R17465 DIFFPAIR_BIAS.n18 DIFFPAIR_BIAS.n0 3.49141
R17466 DIFFPAIR_BIAS.n37 DIFFPAIR_BIAS.n19 3.49141
R17467 DIFFPAIR_BIAS.n57 DIFFPAIR_BIAS.n39 3.49141
R17468 DIFFPAIR_BIAS.n16 DIFFPAIR_BIAS.n15 2.71565
R17469 DIFFPAIR_BIAS.n35 DIFFPAIR_BIAS.n34 2.71565
R17470 DIFFPAIR_BIAS.n55 DIFFPAIR_BIAS.n54 2.71565
R17471 DIFFPAIR_BIAS.n60 DIFFPAIR_BIAS.n59 2.08358
R17472 DIFFPAIR_BIAS.n63 DIFFPAIR_BIAS.n62 2.08355
R17473 DIFFPAIR_BIAS.n58 DIFFPAIR_BIAS.n38 2.0819
R17474 DIFFPAIR_BIAS.n12 DIFFPAIR_BIAS.n2 1.93989
R17475 DIFFPAIR_BIAS.n31 DIFFPAIR_BIAS.n21 1.93989
R17476 DIFFPAIR_BIAS.n51 DIFFPAIR_BIAS.n41 1.93989
R17477 DIFFPAIR_BIAS DIFFPAIR_BIAS.n64 1.19612
R17478 DIFFPAIR_BIAS.n11 DIFFPAIR_BIAS.n4 1.16414
R17479 DIFFPAIR_BIAS.n30 DIFFPAIR_BIAS.n23 1.16414
R17480 DIFFPAIR_BIAS.n50 DIFFPAIR_BIAS.n43 1.16414
R17481 DIFFPAIR_BIAS.n8 DIFFPAIR_BIAS.n7 0.388379
R17482 DIFFPAIR_BIAS.n27 DIFFPAIR_BIAS.n26 0.388379
R17483 DIFFPAIR_BIAS.n47 DIFFPAIR_BIAS.n46 0.388379
R17484 DIFFPAIR_BIAS.n64 DIFFPAIR_BIAS.n63 0.376161
R17485 DIFFPAIR_BIAS.n17 DIFFPAIR_BIAS.n1 0.155672
R17486 DIFFPAIR_BIAS.n10 DIFFPAIR_BIAS.n1 0.155672
R17487 DIFFPAIR_BIAS.n10 DIFFPAIR_BIAS.n9 0.155672
R17488 DIFFPAIR_BIAS.n36 DIFFPAIR_BIAS.n20 0.155672
R17489 DIFFPAIR_BIAS.n29 DIFFPAIR_BIAS.n20 0.155672
R17490 DIFFPAIR_BIAS.n29 DIFFPAIR_BIAS.n28 0.155672
R17491 DIFFPAIR_BIAS.n56 DIFFPAIR_BIAS.n40 0.155672
R17492 DIFFPAIR_BIAS.n49 DIFFPAIR_BIAS.n40 0.155672
R17493 DIFFPAIR_BIAS.n49 DIFFPAIR_BIAS.n48 0.155672
R17494 a_n1379_n2440.n25 a_n1379_n2440.n1 215.069
R17495 a_n1379_n2440.n22 a_n1379_n2440.n3 215.069
R17496 a_n1379_n2440.n5 a_n1379_n2440.n29 215.069
R17497 a_n1379_n2440.n0 a_n1379_n2440.n1 7.91264
R17498 a_n1379_n2440.n25 a_n1379_n2440.n7 185
R17499 a_n1379_n2440.n17 a_n1379_n2440.n16 185
R17500 a_n1379_n2440.n12 a_n1379_n2440.n24 187.962
R17501 a_n1379_n2440.n2 a_n1379_n2440.n3 7.91264
R17502 a_n1379_n2440.n22 a_n1379_n2440.n9 185
R17503 a_n1379_n2440.n19 a_n1379_n2440.n18 185
R17504 a_n1379_n2440.n13 a_n1379_n2440.n21 187.962
R17505 a_n1379_n2440.n4 a_n1379_n2440.n5 7.91264
R17506 a_n1379_n2440.n29 a_n1379_n2440.n11 185
R17507 a_n1379_n2440.n10 a_n1379_n2440.n30 185
R17508 a_n1379_n2440.n15 a_n1379_n2440.n20 187.962
R17509 a_n1379_n2440.n27 a_n1379_n2440.n23 115.178
R17510 a_n1379_n2440.n28 a_n1379_n2440.n27 115.178
R17511 a_n1379_n2440.n27 a_n1379_n2440.n26 113.097
R17512 a_n1379_n2440.n25 a_n1379_n2440.n16 104.615
R17513 a_n1379_n2440.n24 a_n1379_n2440.n16 104.615
R17514 a_n1379_n2440.n22 a_n1379_n2440.n18 104.615
R17515 a_n1379_n2440.n21 a_n1379_n2440.n18 104.615
R17516 a_n1379_n2440.n30 a_n1379_n2440.n29 104.615
R17517 a_n1379_n2440.n30 a_n1379_n2440.n20 104.615
R17518 a_n1379_n2440.n24 a_n1379_n2440.t2 52.3082
R17519 a_n1379_n2440.n21 a_n1379_n2440.t1 52.3082
R17520 a_n1379_n2440.t0 a_n1379_n2440.n20 52.3082
R17521 a_n1379_n2440.n12 a_n1379_n2440.n17 4.42678
R17522 a_n1379_n2440.n13 a_n1379_n2440.n19 4.42678
R17523 a_n1379_n2440.n15 a_n1379_n2440.n10 4.42678
R17524 a_n1379_n2440.n7 a_n1379_n2440.n17 12.0247
R17525 a_n1379_n2440.n9 a_n1379_n2440.n19 12.0247
R17526 a_n1379_n2440.n11 a_n1379_n2440.n10 12.0247
R17527 a_n1379_n2440.n26 a_n1379_n2440.n6 9.45567
R17528 a_n1379_n2440.n23 a_n1379_n2440.n8 9.45567
R17529 a_n1379_n2440.n14 a_n1379_n2440.n28 9.45567
R17530 a_n1379_n2440.n6 a_n1379_n2440.t2 150.207
R17531 a_n1379_n2440.n8 a_n1379_n2440.t1 150.207
R17532 a_n1379_n2440.t0 a_n1379_n2440.n14 150.207
R17533 a_n1379_n2440.n6 a_n1379_n2440.n0 3.91495
R17534 a_n1379_n2440.n8 a_n1379_n2440.n2 3.91495
R17535 a_n1379_n2440.n14 a_n1379_n2440.n4 3.91495
R17536 a_n1379_n2440.n11 a_n1379_n2440.n4 3.6652
R17537 a_n1379_n2440.n9 a_n1379_n2440.n2 3.6652
R17538 a_n1379_n2440.n7 a_n1379_n2440.n0 3.6652
R17539 a_n1379_n2440.n14 a_n1379_n2440.n15 2.42091
R17540 a_n1379_n2440.n13 a_n1379_n2440.n8 2.42091
R17541 a_n1379_n2440.n12 a_n1379_n2440.n6 2.42091
R17542 a_n1379_n2440.n26 a_n1379_n2440.n1 9.74451
R17543 a_n1379_n2440.n23 a_n1379_n2440.n3 9.74451
R17544 a_n1379_n2440.n5 a_n1379_n2440.n28 9.74451
R17545 a_n874_n120.n24 a_n874_n120.n19 289.615
R17546 a_n874_n120.n35 a_n874_n120.n30 289.615
R17547 a_n874_n120.n44 a_n874_n120.n17 289.615
R17548 a_n874_n120.n25 a_n874_n120.n24 185
R17549 a_n874_n120.n23 a_n874_n120.n22 185
R17550 a_n874_n120.n3 a_n874_n120.n2 185
R17551 a_n874_n120.n11 a_n874_n120.n21 185
R17552 a_n874_n120.n36 a_n874_n120.n35 185
R17553 a_n874_n120.n34 a_n874_n120.n33 185
R17554 a_n874_n120.n5 a_n874_n120.n4 185
R17555 a_n874_n120.n13 a_n874_n120.n32 185
R17556 a_n874_n120.n18 a_n874_n120.n17 185
R17557 a_n874_n120.n48 a_n874_n120.n47 185
R17558 a_n874_n120.n6 a_n874_n120.n49 185
R17559 a_n874_n120.n15 a_n874_n120.n14 185
R17560 a_n874_n120.n1 a_n874_n120.n38 140.831
R17561 a_n874_n120.n0 a_n874_n120.n27 140.637
R17562 a_n874_n120.n43 a_n874_n120.n42 140.637
R17563 a_n874_n120.n24 a_n874_n120.n23 104.615
R17564 a_n874_n120.n23 a_n874_n120.n2 104.615
R17565 a_n874_n120.n21 a_n874_n120.n2 104.615
R17566 a_n874_n120.n35 a_n874_n120.n34 104.615
R17567 a_n874_n120.n34 a_n874_n120.n4 104.615
R17568 a_n874_n120.n32 a_n874_n120.n4 104.615
R17569 a_n874_n120.n48 a_n874_n120.n17 104.615
R17570 a_n874_n120.n49 a_n874_n120.n48 104.615
R17571 a_n874_n120.n49 a_n874_n120.n14 104.615
R17572 a_n874_n120.n29 a_n874_n120.t0 70.8207
R17573 a_n874_n120.n40 a_n874_n120.t1 70.8205
R17574 a_n874_n120.n39 a_n874_n120.t6 70.8205
R17575 a_n874_n120.n28 a_n874_n120.t5 70.8205
R17576 a_n874_n120.n21 a_n874_n120.t3 52.3082
R17577 a_n874_n120.n32 a_n874_n120.t2 52.3082
R17578 a_n874_n120.t4 a_n874_n120.n14 52.3082
R17579 a_n874_n120.n11 a_n874_n120.n10 5.0984
R17580 a_n874_n120.n13 a_n874_n120.n12 5.0984
R17581 a_n874_n120.n16 a_n874_n120.n15 5.0984
R17582 a_n874_n120.n11 a_n874_n120.n3 12.8005
R17583 a_n874_n120.n13 a_n874_n120.n5 12.8005
R17584 a_n874_n120.n15 a_n874_n120.n6 12.8005
R17585 a_n874_n120.n1 a_n874_n120.n29 12.1055
R17586 a_n874_n120.n22 a_n874_n120.n3 12.0247
R17587 a_n874_n120.n33 a_n874_n120.n5 12.0247
R17588 a_n874_n120.n47 a_n874_n120.n6 12.0247
R17589 a_n874_n120.n25 a_n874_n120.n20 11.249
R17590 a_n874_n120.n36 a_n874_n120.n31 11.249
R17591 a_n874_n120.n46 a_n874_n120.n18 11.249
R17592 a_n874_n120.n41 a_n874_n120.n28 10.5538
R17593 a_n874_n120.n26 a_n874_n120.n19 10.4732
R17594 a_n874_n120.n37 a_n874_n120.n30 10.4732
R17595 a_n874_n120.n45 a_n874_n120.n44 10.4732
R17596 a_n874_n120.n27 a_n874_n120.n9 9.45567
R17597 a_n874_n120.n38 a_n874_n120.n8 9.45567
R17598 a_n874_n120.n7 a_n874_n120.n43 9.45567
R17599 a_n874_n120.n9 a_n874_n120.n26 9.3005
R17600 a_n874_n120.n20 a_n874_n120.n9 9.3005
R17601 a_n874_n120.n8 a_n874_n120.n37 9.3005
R17602 a_n874_n120.n31 a_n874_n120.n8 9.3005
R17603 a_n874_n120.n7 a_n874_n120.n45 9.3005
R17604 a_n874_n120.n46 a_n874_n120.n7 9.3005
R17605 a_n874_n120.n39 a_n874_n120.n1 8.36688
R17606 a_n874_n120.n41 a_n874_n120.n40 6.81516
R17607 a_n874_n120.n10 a_n874_n120.t3 150.207
R17608 a_n874_n120.n12 a_n874_n120.t2 150.207
R17609 a_n874_n120.t4 a_n874_n120.n16 150.207
R17610 a_n874_n120.n7 a_n874_n120.n6 10.4641
R17611 a_n874_n120.n5 a_n874_n120.n8 10.4641
R17612 a_n874_n120.n3 a_n874_n120.n9 10.4641
R17613 a_n874_n120.n1 a_n874_n120.n0 3.51169
R17614 a_n874_n120.n27 a_n874_n120.n19 3.49141
R17615 a_n874_n120.n38 a_n874_n120.n30 3.49141
R17616 a_n874_n120.n44 a_n874_n120.n43 3.49141
R17617 a_n874_n120.n42 a_n874_n120.n41 3.2268
R17618 a_n874_n120.n26 a_n874_n120.n25 2.71565
R17619 a_n874_n120.n37 a_n874_n120.n36 2.71565
R17620 a_n874_n120.n45 a_n874_n120.n18 2.71565
R17621 a_n874_n120.n42 a_n874_n120.n0 2.0819
R17622 a_n874_n120.n29 a_n874_n120.n28 2.02205
R17623 a_n874_n120.n40 a_n874_n120.n39 2.02205
R17624 a_n874_n120.n22 a_n874_n120.n20 1.93989
R17625 a_n874_n120.n33 a_n874_n120.n31 1.93989
R17626 a_n874_n120.n47 a_n874_n120.n46 1.93989
R17627 a_n874_n120.n9 a_n874_n120.n10 1.90135
R17628 a_n874_n120.n8 a_n874_n120.n12 1.90135
R17629 a_n874_n120.n16 a_n874_n120.n7 1.90135
R17630 CS_BIAS.n5 CS_BIAS.t0 120.767
R17631 CS_BIAS.n0 CS_BIAS.t2 120.287
R17632 CS_BIAS.n4 CS_BIAS.t9 113.302
R17633 CS_BIAS.n9 CS_BIAS.t5 113.302
R17634 CS_BIAS.n8 CS_BIAS.t8 113.302
R17635 CS_BIAS.n7 CS_BIAS.t10 113.302
R17636 CS_BIAS.n3 CS_BIAS.t7 113.3
R17637 CS_BIAS.n2 CS_BIAS.t4 113.3
R17638 CS_BIAS.n1 CS_BIAS.t6 108.188
R17639 CS_BIAS.n6 CS_BIAS.t11 108.188
R17640 CS_BIAS.n5 CS_BIAS.t1 76.5654
R17641 CS_BIAS.n0 CS_BIAS.t3 76.0848
R17642 CS_BIAS.n1 CS_BIAS.n0 10.0382
R17643 CS_BIAS.n6 CS_BIAS.n5 9.55757
R17644 CS_BIAS.n10 CS_BIAS.n4 7.85594
R17645 CS_BIAS.n2 CS_BIAS.n1 7.50554
R17646 CS_BIAS.n7 CS_BIAS.n6 7.50554
R17647 CS_BIAS.n10 CS_BIAS.n9 6.54308
R17648 CS_BIAS CS_BIAS.n10 4.90972
R17649 CS_BIAS.n3 CS_BIAS.n2 2.40202
R17650 CS_BIAS.n4 CS_BIAS.n3 2.40202
R17651 CS_BIAS.n8 CS_BIAS.n7 2.40202
R17652 CS_BIAS.n9 CS_BIAS.n8 2.40202
R17653 VP.n2 VP.t5 243.97
R17654 VP.n5 VP.t0 243.255
R17655 VP.n4 VP.n3 223.454
R17656 VP.n2 VP.n1 223.454
R17657 VP.n0 VP.t7 87.1736
R17658 VP.n0 VP.t6 70.5612
R17659 VP.n3 VP.t2 19.8005
R17660 VP.n3 VP.t4 19.8005
R17661 VP.n1 VP.t1 19.8005
R17662 VP.n1 VP.t3 19.8005
R17663 VP VP.n6 14.1384
R17664 VP.n6 VP.n5 4.80222
R17665 VP.n6 VP.n0 0.972091
R17666 VP.n4 VP.n2 0.716017
R17667 VP.n5 VP.n4 0.716017
R17668 a_n2095_n2440.n22 a_n2095_n2440.n17 289.615
R17669 a_n2095_n2440.n31 a_n2095_n2440.n26 289.615
R17670 a_n2095_n2440.n37 a_n2095_n2440.n15 289.615
R17671 a_n2095_n2440.n23 a_n2095_n2440.n22 185
R17672 a_n2095_n2440.n21 a_n2095_n2440.n20 185
R17673 a_n2095_n2440.n1 a_n2095_n2440.n0 185
R17674 a_n2095_n2440.n9 a_n2095_n2440.n19 185
R17675 a_n2095_n2440.n32 a_n2095_n2440.n31 185
R17676 a_n2095_n2440.n30 a_n2095_n2440.n29 185
R17677 a_n2095_n2440.n3 a_n2095_n2440.n2 185
R17678 a_n2095_n2440.n11 a_n2095_n2440.n28 185
R17679 a_n2095_n2440.n16 a_n2095_n2440.n15 185
R17680 a_n2095_n2440.n41 a_n2095_n2440.n40 185
R17681 a_n2095_n2440.n4 a_n2095_n2440.n42 185
R17682 a_n2095_n2440.n13 a_n2095_n2440.n12 185
R17683 a_n2095_n2440.n22 a_n2095_n2440.n21 104.615
R17684 a_n2095_n2440.n21 a_n2095_n2440.n0 104.615
R17685 a_n2095_n2440.n19 a_n2095_n2440.n0 104.615
R17686 a_n2095_n2440.n31 a_n2095_n2440.n30 104.615
R17687 a_n2095_n2440.n30 a_n2095_n2440.n2 104.615
R17688 a_n2095_n2440.n28 a_n2095_n2440.n2 104.615
R17689 a_n2095_n2440.n41 a_n2095_n2440.n15 104.615
R17690 a_n2095_n2440.n42 a_n2095_n2440.n41 104.615
R17691 a_n2095_n2440.n42 a_n2095_n2440.n12 104.615
R17692 a_n2095_n2440.n19 a_n2095_n2440.t2 52.3082
R17693 a_n2095_n2440.n28 a_n2095_n2440.t0 52.3082
R17694 a_n2095_n2440.t1 a_n2095_n2440.n12 52.3082
R17695 a_n2095_n2440.n35 a_n2095_n2440.n25 46.9122
R17696 a_n2095_n2440.n36 a_n2095_n2440.n35 46.9122
R17697 a_n2095_n2440.n35 a_n2095_n2440.n34 44.8308
R17698 a_n2095_n2440.n9 a_n2095_n2440.n8 5.0984
R17699 a_n2095_n2440.n11 a_n2095_n2440.n10 5.0984
R17700 a_n2095_n2440.n14 a_n2095_n2440.n13 5.0984
R17701 a_n2095_n2440.n9 a_n2095_n2440.n1 12.8005
R17702 a_n2095_n2440.n11 a_n2095_n2440.n3 12.8005
R17703 a_n2095_n2440.n13 a_n2095_n2440.n4 12.8005
R17704 a_n2095_n2440.n20 a_n2095_n2440.n1 12.0247
R17705 a_n2095_n2440.n29 a_n2095_n2440.n3 12.0247
R17706 a_n2095_n2440.n40 a_n2095_n2440.n4 12.0247
R17707 a_n2095_n2440.n23 a_n2095_n2440.n18 11.249
R17708 a_n2095_n2440.n32 a_n2095_n2440.n27 11.249
R17709 a_n2095_n2440.n39 a_n2095_n2440.n16 11.249
R17710 a_n2095_n2440.n24 a_n2095_n2440.n17 10.4732
R17711 a_n2095_n2440.n33 a_n2095_n2440.n26 10.4732
R17712 a_n2095_n2440.n38 a_n2095_n2440.n37 10.4732
R17713 a_n2095_n2440.n25 a_n2095_n2440.n7 9.45567
R17714 a_n2095_n2440.n34 a_n2095_n2440.n6 9.45567
R17715 a_n2095_n2440.n5 a_n2095_n2440.n36 9.45567
R17716 a_n2095_n2440.n7 a_n2095_n2440.n24 9.3005
R17717 a_n2095_n2440.n18 a_n2095_n2440.n7 9.3005
R17718 a_n2095_n2440.n6 a_n2095_n2440.n33 9.3005
R17719 a_n2095_n2440.n27 a_n2095_n2440.n6 9.3005
R17720 a_n2095_n2440.n5 a_n2095_n2440.n38 9.3005
R17721 a_n2095_n2440.n39 a_n2095_n2440.n5 9.3005
R17722 a_n2095_n2440.n8 a_n2095_n2440.t2 150.207
R17723 a_n2095_n2440.n10 a_n2095_n2440.t0 150.207
R17724 a_n2095_n2440.t1 a_n2095_n2440.n14 150.207
R17725 a_n2095_n2440.n5 a_n2095_n2440.n4 10.4641
R17726 a_n2095_n2440.n3 a_n2095_n2440.n6 10.4641
R17727 a_n2095_n2440.n1 a_n2095_n2440.n7 10.4641
R17728 a_n2095_n2440.n25 a_n2095_n2440.n17 3.49141
R17729 a_n2095_n2440.n34 a_n2095_n2440.n26 3.49141
R17730 a_n2095_n2440.n37 a_n2095_n2440.n36 3.49141
R17731 a_n2095_n2440.n24 a_n2095_n2440.n23 2.71565
R17732 a_n2095_n2440.n33 a_n2095_n2440.n32 2.71565
R17733 a_n2095_n2440.n38 a_n2095_n2440.n16 2.71565
R17734 a_n2095_n2440.n20 a_n2095_n2440.n18 1.93989
R17735 a_n2095_n2440.n29 a_n2095_n2440.n27 1.93989
R17736 a_n2095_n2440.n40 a_n2095_n2440.n39 1.93989
R17737 a_n2095_n2440.n7 a_n2095_n2440.n8 1.90135
R17738 a_n2095_n2440.n6 a_n2095_n2440.n10 1.90135
R17739 a_n2095_n2440.n14 a_n2095_n2440.n5 1.90135
C0 VOUT VN 0.936043f
C1 CS_BIAS VP 0.278854f
C2 CS_BIAS VN 0.249318f
C3 CS_BIAS DIFFPAIR_BIAS 0.013021f
C4 VP VN 9.63485f
C5 VP DIFFPAIR_BIAS 0.005394f
C6 a_6779_8904# VDD 1.3156f
C7 VN DIFFPAIR_BIAS 0.005394f
C8 VDD VOUT 50.181896f
C9 a_n7595_8904# VDD 1.31611f
C10 VOUT CS_BIAS 10.709901f
C11 VDD VN 0.1064f
C12 VOUT VP 4.4733f
C13 DIFFPAIR_BIAS GND 17.311876f
C14 VN GND 26.13329f
C15 VP GND 25.75918f
C16 CS_BIAS GND 43.45151f
C17 VOUT GND 55.761627f
C18 VDD GND 0.534119p
C19 a_6779_8904# GND 0.421883f
C20 a_n7595_8904# GND 0.421883f
C21 a_n2095_n2440.n0 GND 0.021523f
C22 a_n2095_n2440.n1 GND 0.018748f
C23 a_n2095_n2440.n2 GND 0.021523f
C24 a_n2095_n2440.n3 GND 0.018748f
C25 a_n2095_n2440.n4 GND 0.018748f
C26 a_n2095_n2440.n5 GND 0.320373f
C27 a_n2095_n2440.n6 GND 0.320373f
C28 a_n2095_n2440.n7 GND 0.320373f
C29 a_n2095_n2440.n8 GND 0.064401f
C30 a_n2095_n2440.n9 GND 0.021774f
C31 a_n2095_n2440.n10 GND 0.064401f
C32 a_n2095_n2440.n11 GND 0.021774f
C33 a_n2095_n2440.n12 GND 0.016143f
C34 a_n2095_n2440.n13 GND 0.021774f
C35 a_n2095_n2440.n14 GND 0.064401f
C36 a_n2095_n2440.n15 GND 0.046999f
C37 a_n2095_n2440.n16 GND 0.009642f
C38 a_n2095_n2440.n17 GND 0.024048f
C39 a_n2095_n2440.n18 GND 0.009106f
C40 a_n2095_n2440.t2 GND 0.036806f
C41 a_n2095_n2440.n19 GND 0.016143f
C42 a_n2095_n2440.n20 GND 0.009642f
C43 a_n2095_n2440.n21 GND 0.021523f
C44 a_n2095_n2440.n22 GND 0.046999f
C45 a_n2095_n2440.n23 GND 0.009642f
C46 a_n2095_n2440.n24 GND 0.009106f
C47 a_n2095_n2440.n25 GND 0.097997f
C48 a_n2095_n2440.n26 GND 0.024048f
C49 a_n2095_n2440.n27 GND 0.009106f
C50 a_n2095_n2440.t0 GND 0.036806f
C51 a_n2095_n2440.n28 GND 0.016143f
C52 a_n2095_n2440.n29 GND 0.009642f
C53 a_n2095_n2440.n30 GND 0.021523f
C54 a_n2095_n2440.n31 GND 0.046999f
C55 a_n2095_n2440.n32 GND 0.009642f
C56 a_n2095_n2440.n33 GND 0.009106f
C57 a_n2095_n2440.n34 GND 0.074597f
C58 a_n2095_n2440.n35 GND 1.92666f
C59 a_n2095_n2440.n36 GND 0.111251f
C60 a_n2095_n2440.n37 GND 0.024048f
C61 a_n2095_n2440.n38 GND 0.009106f
C62 a_n2095_n2440.n39 GND 0.009106f
C63 a_n2095_n2440.n40 GND 0.009642f
C64 a_n2095_n2440.n41 GND 0.021523f
C65 a_n2095_n2440.n42 GND 0.021523f
C66 a_n2095_n2440.t1 GND 0.036806f
C67 VP.t6 GND 0.683107f
C68 VP.t7 GND 0.842103f
C69 VP.n0 GND 1.57534f
C70 VP.t5 GND 0.031656f
C71 VP.t1 GND 0.005653f
C72 VP.t3 GND 0.005653f
C73 VP.n1 GND 0.018334f
C74 VP.n2 GND 0.142326f
C75 VP.t2 GND 0.005653f
C76 VP.t4 GND 0.005653f
C77 VP.n3 GND 0.018334f
C78 VP.n4 GND 0.076922f
C79 VP.t0 GND 0.031464f
C80 VP.n5 GND 0.085384f
C81 VP.n6 GND 2.15124f
C82 CS_BIAS.t6 GND 0.199495f
C83 CS_BIAS.t2 GND 0.210241f
C84 CS_BIAS.t3 GND 0.085935f
C85 CS_BIAS.n0 GND 0.197676f
C86 CS_BIAS.n1 GND 0.135063f
C87 CS_BIAS.t4 GND 0.203212f
C88 CS_BIAS.n2 GND 0.154633f
C89 CS_BIAS.t7 GND 0.203212f
C90 CS_BIAS.n3 GND 0.133868f
C91 CS_BIAS.t9 GND 0.203213f
C92 CS_BIAS.n4 GND 0.330364f
C93 CS_BIAS.t11 GND 0.199495f
C94 CS_BIAS.t1 GND 0.086127f
C95 CS_BIAS.t0 GND 0.210775f
C96 CS_BIAS.n5 GND 0.214947f
C97 CS_BIAS.n6 GND 0.133146f
C98 CS_BIAS.t10 GND 0.203213f
C99 CS_BIAS.n7 GND 0.154633f
C100 CS_BIAS.t8 GND 0.203213f
C101 CS_BIAS.n8 GND 0.133867f
C102 CS_BIAS.t5 GND 0.203213f
C103 CS_BIAS.n9 GND 0.188043f
C104 CS_BIAS.n10 GND 3.8132f
C105 a_n874_n120.n0 GND 0.552481f
C106 a_n874_n120.n1 GND 1.18466f
C107 a_n874_n120.n2 GND 0.0202f
C108 a_n874_n120.n3 GND 0.017595f
C109 a_n874_n120.n4 GND 0.0202f
C110 a_n874_n120.n5 GND 0.017595f
C111 a_n874_n120.n6 GND 0.017595f
C112 a_n874_n120.n7 GND 0.300671f
C113 a_n874_n120.n8 GND 0.300671f
C114 a_n874_n120.n9 GND 0.300671f
C115 a_n874_n120.n10 GND 0.060441f
C116 a_n874_n120.n11 GND 0.020435f
C117 a_n874_n120.n12 GND 0.060441f
C118 a_n874_n120.n13 GND 0.020435f
C119 a_n874_n120.n14 GND 0.01515f
C120 a_n874_n120.n15 GND 0.020435f
C121 a_n874_n120.n16 GND 0.060441f
C122 a_n874_n120.n17 GND 0.044109f
C123 a_n874_n120.n18 GND 0.009049f
C124 a_n874_n120.n19 GND 0.022569f
C125 a_n874_n120.n20 GND 0.008546f
C126 a_n874_n120.t3 GND 0.034543f
C127 a_n874_n120.n21 GND 0.01515f
C128 a_n874_n120.n22 GND 0.009049f
C129 a_n874_n120.n23 GND 0.0202f
C130 a_n874_n120.n24 GND 0.044109f
C131 a_n874_n120.n25 GND 0.009049f
C132 a_n874_n120.n26 GND 0.008546f
C133 a_n874_n120.n27 GND 0.09424f
C134 a_n874_n120.t5 GND 0.285561f
C135 a_n874_n120.n28 GND 0.57598f
C136 a_n874_n120.t0 GND 0.285562f
C137 a_n874_n120.n29 GND 0.683926f
C138 a_n874_n120.n30 GND 0.022569f
C139 a_n874_n120.n31 GND 0.008546f
C140 a_n874_n120.t2 GND 0.034543f
C141 a_n874_n120.n32 GND 0.01515f
C142 a_n874_n120.n33 GND 0.009049f
C143 a_n874_n120.n34 GND 0.0202f
C144 a_n874_n120.n35 GND 0.044109f
C145 a_n874_n120.n36 GND 0.009049f
C146 a_n874_n120.n37 GND 0.008546f
C147 a_n874_n120.n38 GND 0.094429f
C148 a_n874_n120.t6 GND 0.285561f
C149 a_n874_n120.n39 GND 0.573366f
C150 a_n874_n120.t1 GND 0.285561f
C151 a_n874_n120.n40 GND 0.468275f
C152 a_n874_n120.n41 GND 0.770056f
C153 a_n874_n120.n42 GND 0.692793f
C154 a_n874_n120.n43 GND 0.09424f
C155 a_n874_n120.n44 GND 0.022569f
C156 a_n874_n120.n45 GND 0.008546f
C157 a_n874_n120.n46 GND 0.008546f
C158 a_n874_n120.n47 GND 0.009049f
C159 a_n874_n120.n48 GND 0.0202f
C160 a_n874_n120.n49 GND 0.0202f
C161 a_n874_n120.t4 GND 0.034543f
C162 a_n1379_n2440.n0 GND 0.01362f
C163 a_n1379_n2440.n1 GND 0.058654f
C164 a_n1379_n2440.n2 GND 0.01362f
C165 a_n1379_n2440.n3 GND 0.058654f
C166 a_n1379_n2440.n4 GND 0.01362f
C167 a_n1379_n2440.n5 GND 0.058654f
C168 a_n1379_n2440.n6 GND 0.553698f
C169 a_n1379_n2440.n7 GND 0.026979f
C170 a_n1379_n2440.n8 GND 0.553698f
C171 a_n1379_n2440.n9 GND 0.026979f
C172 a_n1379_n2440.n10 GND 0.026979f
C173 a_n1379_n2440.n11 GND 0.026979f
C174 a_n1379_n2440.n12 GND 0.03084f
C175 a_n1379_n2440.n13 GND 0.03084f
C176 a_n1379_n2440.n14 GND 0.553698f
C177 a_n1379_n2440.n15 GND 0.03084f
C178 a_n1379_n2440.n16 GND 0.030973f
C179 a_n1379_n2440.n17 GND 0.026979f
C180 a_n1379_n2440.n18 GND 0.030973f
C181 a_n1379_n2440.n19 GND 0.026979f
C182 a_n1379_n2440.t2 GND 0.052965f
C183 a_n1379_n2440.t1 GND 0.052965f
C184 a_n1379_n2440.n20 GND 0.023723f
C185 a_n1379_n2440.n21 GND 0.023723f
C186 a_n1379_n2440.n22 GND 0.065707f
C187 a_n1379_n2440.n23 GND 0.160087f
C188 a_n1379_n2440.n24 GND 0.023723f
C189 a_n1379_n2440.n25 GND 0.065707f
C190 a_n1379_n2440.n26 GND 0.145387f
C191 a_n1379_n2440.n27 GND 2.7768f
C192 a_n1379_n2440.n28 GND 0.165314f
C193 a_n1379_n2440.n29 GND 0.065707f
C194 a_n1379_n2440.n30 GND 0.030973f
C195 a_n1379_n2440.t0 GND 0.052965f
C196 DIFFPAIR_BIAS.t6 GND 0.48964f
C197 DIFFPAIR_BIAS.n0 GND 0.006835f
C198 DIFFPAIR_BIAS.n1 GND 0.004816f
C199 DIFFPAIR_BIAS.n2 GND 0.002588f
C200 DIFFPAIR_BIAS.n3 GND 0.006117f
C201 DIFFPAIR_BIAS.n4 GND 0.00274f
C202 DIFFPAIR_BIAS.n5 GND 0.01859f
C203 DIFFPAIR_BIAS.t3 GND 0.010174f
C204 DIFFPAIR_BIAS.n6 GND 0.004588f
C205 DIFFPAIR_BIAS.n7 GND 0.0036f
C206 DIFFPAIR_BIAS.n8 GND 0.002588f
C207 DIFFPAIR_BIAS.n9 GND 0.069367f
C208 DIFFPAIR_BIAS.n10 GND 0.004816f
C209 DIFFPAIR_BIAS.n11 GND 0.002588f
C210 DIFFPAIR_BIAS.n12 GND 0.00274f
C211 DIFFPAIR_BIAS.n13 GND 0.006117f
C212 DIFFPAIR_BIAS.n14 GND 0.013358f
C213 DIFFPAIR_BIAS.n15 GND 0.00274f
C214 DIFFPAIR_BIAS.n16 GND 0.002588f
C215 DIFFPAIR_BIAS.n17 GND 0.012054f
C216 DIFFPAIR_BIAS.n18 GND 0.02474f
C217 DIFFPAIR_BIAS.n19 GND 0.006835f
C218 DIFFPAIR_BIAS.n20 GND 0.004816f
C219 DIFFPAIR_BIAS.n21 GND 0.002588f
C220 DIFFPAIR_BIAS.n22 GND 0.006117f
C221 DIFFPAIR_BIAS.n23 GND 0.00274f
C222 DIFFPAIR_BIAS.n24 GND 0.01859f
C223 DIFFPAIR_BIAS.t5 GND 0.010174f
C224 DIFFPAIR_BIAS.n25 GND 0.004588f
C225 DIFFPAIR_BIAS.n26 GND 0.0036f
C226 DIFFPAIR_BIAS.n27 GND 0.002588f
C227 DIFFPAIR_BIAS.n28 GND 0.069367f
C228 DIFFPAIR_BIAS.n29 GND 0.004816f
C229 DIFFPAIR_BIAS.n30 GND 0.002588f
C230 DIFFPAIR_BIAS.n31 GND 0.00274f
C231 DIFFPAIR_BIAS.n32 GND 0.006117f
C232 DIFFPAIR_BIAS.n33 GND 0.013358f
C233 DIFFPAIR_BIAS.n34 GND 0.00274f
C234 DIFFPAIR_BIAS.n35 GND 0.002588f
C235 DIFFPAIR_BIAS.n36 GND 0.012054f
C236 DIFFPAIR_BIAS.n37 GND 0.020131f
C237 DIFFPAIR_BIAS.n38 GND 0.341263f
C238 DIFFPAIR_BIAS.n39 GND 0.006835f
C239 DIFFPAIR_BIAS.n40 GND 0.004816f
C240 DIFFPAIR_BIAS.n41 GND 0.002588f
C241 DIFFPAIR_BIAS.n42 GND 0.006117f
C242 DIFFPAIR_BIAS.n43 GND 0.00274f
C243 DIFFPAIR_BIAS.n44 GND 0.01859f
C244 DIFFPAIR_BIAS.t1 GND 0.010174f
C245 DIFFPAIR_BIAS.n45 GND 0.004588f
C246 DIFFPAIR_BIAS.n46 GND 0.0036f
C247 DIFFPAIR_BIAS.n47 GND 0.002588f
C248 DIFFPAIR_BIAS.n48 GND 0.069367f
C249 DIFFPAIR_BIAS.n49 GND 0.004816f
C250 DIFFPAIR_BIAS.n50 GND 0.002588f
C251 DIFFPAIR_BIAS.n51 GND 0.00274f
C252 DIFFPAIR_BIAS.n52 GND 0.006117f
C253 DIFFPAIR_BIAS.n53 GND 0.013358f
C254 DIFFPAIR_BIAS.n54 GND 0.00274f
C255 DIFFPAIR_BIAS.n55 GND 0.002588f
C256 DIFFPAIR_BIAS.n56 GND 0.012054f
C257 DIFFPAIR_BIAS.n57 GND 0.020131f
C258 DIFFPAIR_BIAS.n58 GND 0.210199f
C259 DIFFPAIR_BIAS.t0 GND 0.465411f
C260 DIFFPAIR_BIAS.t4 GND 0.465411f
C261 DIFFPAIR_BIAS.t2 GND 0.470993f
C262 DIFFPAIR_BIAS.n59 GND 0.592093f
C263 DIFFPAIR_BIAS.n60 GND 0.359809f
C264 DIFFPAIR_BIAS.n61 GND 0.638789f
C265 DIFFPAIR_BIAS.t8 GND 0.48644f
C266 DIFFPAIR_BIAS.n62 GND 0.308929f
C267 DIFFPAIR_BIAS.t7 GND 0.48644f
C268 DIFFPAIR_BIAS.n63 GND 0.256841f
C269 DIFFPAIR_BIAS.n64 GND 0.624648f
C270 VN.t6 GND 0.37593f
C271 VN.t7 GND 0.462728f
C272 VN.n0 GND 0.861663f
C273 VN.t1 GND 0.017469f
C274 VN.t2 GND 0.00312f
C275 VN.t4 GND 0.00312f
C276 VN.n1 GND 0.010117f
C277 VN.n2 GND 0.07854f
C278 VN.t3 GND 0.00312f
C279 VN.t5 GND 0.00312f
C280 VN.n3 GND 0.010117f
C281 VN.n4 GND 0.042448f
C282 VN.t0 GND 0.017363f
C283 VN.n5 GND 0.052607f
C284 VN.n6 GND 1.63875f
C285 a_n5180_7124.t0 GND 66.4765f
C286 a_n5180_7124.t9 GND 0.406554f
C287 a_n5180_7124.t15 GND 0.050277f
C288 a_n5180_7124.t12 GND 0.050277f
C289 a_n5180_7124.n0 GND 0.282746f
C290 a_n5180_7124.n1 GND 0.816569f
C291 a_n5180_7124.t13 GND 0.050277f
C292 a_n5180_7124.t10 GND 0.050277f
C293 a_n5180_7124.n2 GND 0.282746f
C294 a_n5180_7124.n3 GND 0.747192f
C295 a_n5180_7124.n4 GND 3.43031f
C296 a_n5180_7124.t7 GND 0.406556f
C297 a_n5180_7124.t3 GND 0.050277f
C298 a_n5180_7124.t2 GND 0.050277f
C299 a_n5180_7124.n5 GND 0.282746f
C300 a_n5180_7124.n6 GND 0.816567f
C301 a_n5180_7124.t5 GND 0.394705f
C302 a_n5180_7124.n7 GND 0.393781f
C303 a_n5180_7124.t8 GND 0.394705f
C304 a_n5180_7124.n8 GND 0.393781f
C305 a_n5180_7124.t6 GND 0.050277f
C306 a_n5180_7124.t1 GND 0.050277f
C307 a_n5180_7124.n9 GND 0.282746f
C308 a_n5180_7124.n10 GND 0.462012f
C309 a_n5180_7124.t4 GND 0.394705f
C310 a_n5180_7124.n11 GND 0.539973f
C311 a_n5180_7124.n12 GND 1.4006f
C312 a_n5180_7124.t16 GND 0.050277f
C313 a_n5180_7124.t14 GND 0.050277f
C314 a_n5180_7124.n13 GND 0.282746f
C315 a_n5180_7124.n14 GND 1.30254f
C316 a_n5180_7124.t18 GND 0.050277f
C317 a_n5180_7124.t11 GND 0.050277f
C318 a_n5180_7124.n15 GND 0.282746f
C319 a_n5180_7124.n16 GND 0.816567f
C320 a_n5180_7124.t17 GND 0.406556f
C321 a_n6651_8904.t14 GND 0.138098f
C322 a_n6651_8904.t12 GND 1.21425f
C323 a_n6651_8904.t9 GND 0.138098f
C324 a_n6651_8904.t11 GND 0.138098f
C325 a_n6651_8904.n0 GND 0.875822f
C326 a_n6651_8904.n1 GND 2.13934f
C327 a_n6651_8904.t13 GND 1.20388f
C328 a_n6651_8904.t10 GND 0.138098f
C329 a_n6651_8904.t15 GND 0.138098f
C330 a_n6651_8904.n2 GND 0.875822f
C331 a_n6651_8904.n3 GND 4.14175f
C332 a_n6651_8904.t8 GND 0.138098f
C333 a_n6651_8904.t17 GND 0.138098f
C334 a_n6651_8904.n4 GND 0.875822f
C335 a_n6651_8904.n5 GND 5.36779f
C336 a_n6651_8904.t4 GND 1.11671f
C337 a_n6651_8904.t1 GND 0.138098f
C338 a_n6651_8904.t5 GND 0.138098f
C339 a_n6651_8904.n6 GND 0.776637f
C340 a_n6651_8904.n7 GND 2.24292f
C341 a_n6651_8904.t0 GND 1.08416f
C342 a_n6651_8904.n8 GND 1.08162f
C343 a_n6651_8904.t2 GND 1.08416f
C344 a_n6651_8904.n9 GND 1.08162f
C345 a_n6651_8904.t6 GND 0.138098f
C346 a_n6651_8904.t3 GND 0.138098f
C347 a_n6651_8904.n10 GND 0.776637f
C348 a_n6651_8904.n11 GND 1.26904f
C349 a_n6651_8904.t7 GND 1.08416f
C350 a_n6651_8904.n12 GND 1.48318f
C351 a_n6651_8904.n13 GND 3.95893f
C352 a_n6651_8904.n14 GND 2.23275f
C353 a_n6651_8904.n15 GND 0.875823f
C354 a_n6651_8904.t16 GND 0.138098f
C355 a_n6573_8708.n0 GND 4.96384f
C356 a_n6573_8708.n1 GND 0.593848f
C357 a_n6573_8708.n2 GND 0.593848f
C358 a_n6573_8708.n3 GND 2.06371f
C359 a_n6573_8708.n4 GND 0.183109f
C360 a_n6573_8708.n5 GND 1.9762f
C361 a_n6573_8708.n6 GND 0.183109f
C362 a_n6573_8708.n7 GND 1.93211f
C363 a_n6573_8708.n8 GND 0.183109f
C364 a_n6573_8708.n9 GND 3.92556f
C365 a_n6573_8708.n10 GND 0.183109f
C366 a_n6573_8708.n11 GND 0.176649f
C367 a_n6573_8708.n12 GND 1.69623f
C368 a_n6573_8708.n13 GND 1.59579f
C369 a_n6573_8708.n14 GND 0.176077f
C370 a_n6573_8708.n15 GND 0.176077f
C371 a_n6573_8708.n16 GND 0.176077f
C372 a_n6573_8708.n17 GND 0.176077f
C373 a_n6573_8708.n18 GND 0.176649f
C374 a_n6573_8708.n19 GND 0.176649f
C375 a_n6573_8708.n20 GND 0.176649f
C376 a_n6573_8708.n21 GND 0.593848f
C377 a_n6573_8708.n22 GND 0.593848f
C378 a_n6573_8708.n23 GND 0.591781f
C379 a_n6573_8708.n24 GND 0.59178f
C380 a_n6573_8708.n25 GND 0.591781f
C381 a_n6573_8708.n26 GND 0.59178f
C382 a_n6573_8708.n27 GND 0.591781f
C383 a_n6573_8708.n28 GND 0.59178f
C384 a_n6573_8708.n29 GND 0.591781f
C385 a_n6573_8708.n30 GND 0.59178f
C386 a_n6573_8708.n31 GND 0.59385f
C387 a_n6573_8708.n32 GND 0.59385f
C388 a_n6573_8708.n33 GND 0.59385f
C389 a_n6573_8708.n34 GND 0.59385f
C390 a_n6573_8708.n35 GND 1.1333f
C391 a_n6573_8708.n36 GND 0.761173f
C392 a_n6573_8708.n37 GND 0.761173f
C393 a_n6573_8708.t4 GND 1.81172f
C394 a_n6573_8708.t14 GND 1.45379f
C395 a_n6573_8708.n38 GND 0.764358f
C396 a_n6573_8708.t8 GND 1.45379f
C397 a_n6573_8708.n39 GND 0.761173f
C398 a_n6573_8708.t20 GND 1.45379f
C399 a_n6573_8708.n40 GND 0.757326f
C400 a_n6573_8708.t2 GND 1.81172f
C401 a_n6573_8708.t30 GND 1.81172f
C402 a_n6573_8708.t34 GND 1.45379f
C403 a_n6573_8708.n41 GND 0.764358f
C404 a_n6573_8708.t23 GND 1.45379f
C405 a_n6573_8708.n42 GND 0.761173f
C406 a_n6573_8708.t41 GND 1.45379f
C407 a_n6573_8708.n43 GND 0.757326f
C408 a_n6573_8708.t29 GND 1.81172f
C409 a_n6573_8708.t19 GND 0.360109f
C410 a_n6573_8708.t11 GND 0.051848f
C411 a_n6573_8708.t17 GND 0.343433f
C412 a_n6573_8708.t13 GND 0.051848f
C413 a_n6573_8708.t7 GND 0.407041f
C414 a_n6573_8708.t6 GND 1.81172f
C415 a_n6573_8708.t12 GND 1.45379f
C416 a_n6573_8708.n44 GND 0.757326f
C417 a_n6573_8708.t16 GND 1.45379f
C418 a_n6573_8708.t10 GND 1.45379f
C419 a_n6573_8708.n45 GND 0.764358f
C420 a_n6573_8708.t18 GND 1.81172f
C421 a_n6573_8708.t46 GND 1.81172f
C422 a_n6573_8708.t40 GND 1.45379f
C423 a_n6573_8708.n46 GND 0.757326f
C424 a_n6573_8708.t33 GND 1.45379f
C425 a_n6573_8708.t43 GND 1.45379f
C426 a_n6573_8708.n47 GND 0.764358f
C427 a_n6573_8708.t35 GND 1.81172f
C428 a_n6573_8708.n48 GND 0.678708f
C429 a_n6573_8708.t22 GND 1.80668f
C430 a_n6573_8708.t28 GND 1.45379f
C431 a_n6573_8708.n49 GND 0.765601f
C432 a_n6573_8708.t36 GND 1.80668f
C433 a_n6573_8708.t45 GND 1.80668f
C434 a_n6573_8708.t25 GND 1.45379f
C435 a_n6573_8708.n50 GND 0.765601f
C436 a_n6573_8708.t26 GND 1.80668f
C437 a_n6573_8708.t31 GND 1.80668f
C438 a_n6573_8708.t44 GND 1.45379f
C439 a_n6573_8708.n51 GND 0.765601f
C440 a_n6573_8708.t37 GND 1.80668f
C441 a_n6573_8708.t27 GND 1.80668f
C442 a_n6573_8708.t47 GND 1.45379f
C443 a_n6573_8708.n52 GND 0.765601f
C444 a_n6573_8708.t39 GND 1.80668f
C445 a_n6573_8708.t32 GND 1.45379f
C446 a_n6573_8708.n53 GND 0.765602f
C447 a_n6573_8708.t42 GND 1.45379f
C448 a_n6573_8708.n54 GND 0.765602f
C449 a_n6573_8708.t38 GND 1.45379f
C450 a_n6573_8708.n55 GND 0.765602f
C451 a_n6573_8708.t24 GND 1.45379f
C452 a_n6573_8708.n56 GND 0.765602f
C453 a_n6573_8708.n57 GND 0.661709f
C454 a_n6573_8708.t1 GND 0.429046f
C455 a_n6573_8708.t0 GND 0.257506f
C456 a_n6573_8708.n58 GND 3.0547f
C457 a_n6573_8708.t5 GND 0.343433f
C458 a_n6573_8708.t15 GND 0.051848f
C459 a_n6573_8708.t9 GND 0.343433f
C460 a_n6573_8708.t21 GND 0.051848f
C461 a_n6573_8708.t3 GND 0.419265f
C462 VDD.t183 GND 0.016423f
C463 VDD.t176 GND 0.016423f
C464 VDD.n0 GND 0.108433f
C465 VDD.t22 GND 0.016423f
C466 VDD.t179 GND 0.016423f
C467 VDD.n1 GND 0.104157f
C468 VDD.n2 GND 0.297274f
C469 VDD.t11 GND 0.016423f
C470 VDD.t24 GND 0.016423f
C471 VDD.n3 GND 0.104157f
C472 VDD.n4 GND 0.155247f
C473 VDD.t3 GND 0.016423f
C474 VDD.t17 GND 0.016423f
C475 VDD.n5 GND 0.104157f
C476 VDD.n6 GND 0.135548f
C477 VDD.t32 GND 0.016423f
C478 VDD.t1 GND 0.016423f
C479 VDD.n7 GND 0.108433f
C480 VDD.t15 GND 0.016423f
C481 VDD.t8 GND 0.016423f
C482 VDD.n8 GND 0.104157f
C483 VDD.n9 GND 0.297274f
C484 VDD.t28 GND 0.016423f
C485 VDD.t181 GND 0.016423f
C486 VDD.n10 GND 0.104157f
C487 VDD.n11 GND 0.155247f
C488 VDD.t126 GND 0.016423f
C489 VDD.t30 GND 0.016423f
C490 VDD.n12 GND 0.104157f
C491 VDD.n13 GND 0.135548f
C492 VDD.n14 GND 0.092609f
C493 VDD.n15 GND 2.67329f
C494 VDD.n16 GND 0.004201f
C495 VDD.n17 GND 0.028145f
C496 VDD.n18 GND 0.00219f
C497 VDD.t174 GND 0.011388f
C498 VDD.n19 GND 0.013332f
C499 VDD.n20 GND 0.003052f
C500 VDD.n21 GND 0.003882f
C501 VDD.n22 GND 0.011589f
C502 VDD.n23 GND 0.002319f
C503 VDD.n24 GND 0.00219f
C504 VDD.n25 GND 0.009698f
C505 VDD.n26 GND 0.014383f
C506 VDD.t146 GND 0.00789f
C507 VDD.t139 GND 0.00789f
C508 VDD.n27 GND 0.032694f
C509 VDD.n28 GND 0.23237f
C510 VDD.n29 GND 0.004201f
C511 VDD.n30 GND 0.028145f
C512 VDD.n31 GND 0.00219f
C513 VDD.t167 GND 0.011388f
C514 VDD.n32 GND 0.013332f
C515 VDD.n33 GND 0.003052f
C516 VDD.n34 GND 0.003882f
C517 VDD.n35 GND 0.011589f
C518 VDD.n36 GND 0.002319f
C519 VDD.n37 GND 0.00219f
C520 VDD.n38 GND 0.009698f
C521 VDD.n39 GND 0.005795f
C522 VDD.n40 GND 0.090594f
C523 VDD.n41 GND 0.004201f
C524 VDD.n42 GND 0.028145f
C525 VDD.n43 GND 0.00219f
C526 VDD.t158 GND 0.011388f
C527 VDD.n44 GND 0.013332f
C528 VDD.n45 GND 0.003052f
C529 VDD.n46 GND 0.003882f
C530 VDD.n47 GND 0.011589f
C531 VDD.n48 GND 0.002319f
C532 VDD.n49 GND 0.00219f
C533 VDD.n50 GND 0.009698f
C534 VDD.n51 GND 0.014383f
C535 VDD.t168 GND 0.00789f
C536 VDD.t163 GND 0.00789f
C537 VDD.n52 GND 0.032694f
C538 VDD.n53 GND 0.23237f
C539 VDD.n54 GND 0.004201f
C540 VDD.n55 GND 0.028145f
C541 VDD.n56 GND 0.00219f
C542 VDD.t150 GND 0.011388f
C543 VDD.n57 GND 0.013332f
C544 VDD.n58 GND 0.003052f
C545 VDD.n59 GND 0.003882f
C546 VDD.n60 GND 0.011589f
C547 VDD.n61 GND 0.002319f
C548 VDD.n62 GND 0.00219f
C549 VDD.n63 GND 0.009698f
C550 VDD.n64 GND 0.005795f
C551 VDD.n65 GND 0.081291f
C552 VDD.n66 GND 0.079615f
C553 VDD.n67 GND 0.004201f
C554 VDD.n68 GND 0.028145f
C555 VDD.n69 GND 0.00219f
C556 VDD.t136 GND 0.011388f
C557 VDD.n70 GND 0.013332f
C558 VDD.n71 GND 0.003052f
C559 VDD.n72 GND 0.003882f
C560 VDD.n73 GND 0.011589f
C561 VDD.n74 GND 0.002319f
C562 VDD.n75 GND 0.00219f
C563 VDD.n76 GND 0.009698f
C564 VDD.n77 GND 0.014383f
C565 VDD.t153 GND 0.00789f
C566 VDD.t147 GND 0.00789f
C567 VDD.n78 GND 0.032694f
C568 VDD.n79 GND 0.23237f
C569 VDD.n80 GND 0.004201f
C570 VDD.n81 GND 0.028145f
C571 VDD.n82 GND 0.00219f
C572 VDD.t173 GND 0.011388f
C573 VDD.n83 GND 0.013332f
C574 VDD.n84 GND 0.003052f
C575 VDD.n85 GND 0.003882f
C576 VDD.n86 GND 0.011589f
C577 VDD.n87 GND 0.002319f
C578 VDD.n88 GND 0.00219f
C579 VDD.n89 GND 0.009698f
C580 VDD.n90 GND 0.005795f
C581 VDD.n91 GND 0.081291f
C582 VDD.n92 GND 0.0566f
C583 VDD.n93 GND 0.004201f
C584 VDD.n94 GND 0.028145f
C585 VDD.n95 GND 0.00219f
C586 VDD.t165 GND 0.011388f
C587 VDD.n96 GND 0.013332f
C588 VDD.n97 GND 0.003052f
C589 VDD.n98 GND 0.003882f
C590 VDD.n99 GND 0.011589f
C591 VDD.n100 GND 0.002319f
C592 VDD.n101 GND 0.00219f
C593 VDD.n102 GND 0.009698f
C594 VDD.n103 GND 0.014383f
C595 VDD.t144 GND 0.00789f
C596 VDD.t145 GND 0.00789f
C597 VDD.n104 GND 0.032694f
C598 VDD.n105 GND 0.23237f
C599 VDD.n106 GND 0.004201f
C600 VDD.n107 GND 0.028145f
C601 VDD.n108 GND 0.00219f
C602 VDD.t160 GND 0.011388f
C603 VDD.n109 GND 0.013332f
C604 VDD.n110 GND 0.003052f
C605 VDD.n111 GND 0.003882f
C606 VDD.n112 GND 0.011589f
C607 VDD.n113 GND 0.002319f
C608 VDD.n114 GND 0.00219f
C609 VDD.n115 GND 0.009698f
C610 VDD.n116 GND 0.005795f
C611 VDD.n117 GND 0.081291f
C612 VDD.n118 GND 0.0566f
C613 VDD.n119 GND 0.004201f
C614 VDD.n120 GND 0.028145f
C615 VDD.n121 GND 0.00219f
C616 VDD.t151 GND 0.011388f
C617 VDD.n122 GND 0.013332f
C618 VDD.n123 GND 0.003052f
C619 VDD.n124 GND 0.003882f
C620 VDD.n125 GND 0.011589f
C621 VDD.n126 GND 0.002319f
C622 VDD.n127 GND 0.00219f
C623 VDD.n128 GND 0.009698f
C624 VDD.n129 GND 0.014383f
C625 VDD.t169 GND 0.00789f
C626 VDD.t170 GND 0.00789f
C627 VDD.n130 GND 0.032694f
C628 VDD.n131 GND 0.23237f
C629 VDD.n132 GND 0.004201f
C630 VDD.n133 GND 0.028145f
C631 VDD.n134 GND 0.00219f
C632 VDD.t142 GND 0.011388f
C633 VDD.n135 GND 0.013332f
C634 VDD.n136 GND 0.003052f
C635 VDD.n137 GND 0.003882f
C636 VDD.n138 GND 0.011589f
C637 VDD.n139 GND 0.002319f
C638 VDD.n140 GND 0.00219f
C639 VDD.n141 GND 0.009698f
C640 VDD.n142 GND 0.005795f
C641 VDD.n143 GND 0.081291f
C642 VDD.n144 GND 0.152614f
C643 VDD.n145 GND 0.00615f
C644 VDD.n146 GND 0.008002f
C645 VDD.n147 GND 0.00644f
C646 VDD.n148 GND 0.00644f
C647 VDD.n149 GND 0.008002f
C648 VDD.n150 GND 0.008002f
C649 VDD.n151 GND 0.532804f
C650 VDD.n152 GND 0.008002f
C651 VDD.n153 GND 0.008002f
C652 VDD.n154 GND 0.008002f
C653 VDD.n155 GND 0.532804f
C654 VDD.n156 GND 0.008002f
C655 VDD.n157 GND 0.008002f
C656 VDD.n158 GND 0.008002f
C657 VDD.n159 GND 0.008002f
C658 VDD.n160 GND 0.00644f
C659 VDD.n161 GND 0.008002f
C660 VDD.n162 GND 0.008002f
C661 VDD.n163 GND 0.008002f
C662 VDD.n164 GND 0.008002f
C663 VDD.n165 GND 0.532804f
C664 VDD.n166 GND 0.008002f
C665 VDD.n167 GND 0.008002f
C666 VDD.n168 GND 0.008002f
C667 VDD.n169 GND 0.008002f
C668 VDD.n170 GND 0.008002f
C669 VDD.n171 GND 0.00644f
C670 VDD.n172 GND 0.008002f
C671 VDD.n173 GND 0.008002f
C672 VDD.n174 GND 0.008002f
C673 VDD.n175 GND 0.008002f
C674 VDD.n176 GND 0.532804f
C675 VDD.n177 GND 0.008002f
C676 VDD.n178 GND 0.008002f
C677 VDD.n179 GND 0.008002f
C678 VDD.n180 GND 0.008002f
C679 VDD.n181 GND 0.008002f
C680 VDD.n182 GND 0.00644f
C681 VDD.n183 GND 0.008002f
C682 VDD.n184 GND 0.008002f
C683 VDD.n185 GND 0.008002f
C684 VDD.n186 GND 0.008002f
C685 VDD.n187 GND 0.532804f
C686 VDD.n188 GND 0.008002f
C687 VDD.n189 GND 0.008002f
C688 VDD.n190 GND 0.008002f
C689 VDD.n191 GND 0.008002f
C690 VDD.n192 GND 0.008002f
C691 VDD.n193 GND 0.00644f
C692 VDD.n194 GND 0.008002f
C693 VDD.n195 GND 0.008002f
C694 VDD.n196 GND 0.008002f
C695 VDD.n197 GND 0.008002f
C696 VDD.n198 GND 0.532804f
C697 VDD.n199 GND 0.008002f
C698 VDD.n200 GND 0.008002f
C699 VDD.n201 GND 0.008002f
C700 VDD.n202 GND 0.008002f
C701 VDD.n203 GND 0.008002f
C702 VDD.n204 GND 0.00644f
C703 VDD.n205 GND 0.008002f
C704 VDD.n206 GND 0.008002f
C705 VDD.n207 GND 0.008002f
C706 VDD.n208 GND 0.008002f
C707 VDD.n209 GND 0.532804f
C708 VDD.n210 GND 0.008002f
C709 VDD.n211 GND 0.008002f
C710 VDD.n212 GND 0.008002f
C711 VDD.n213 GND 0.008002f
C712 VDD.n214 GND 0.008002f
C713 VDD.n215 GND 0.00644f
C714 VDD.n216 GND 0.008002f
C715 VDD.n217 GND 0.008002f
C716 VDD.n218 GND 0.008002f
C717 VDD.n219 GND 0.008002f
C718 VDD.n220 GND 0.532804f
C719 VDD.n221 GND 0.008002f
C720 VDD.n222 GND 0.008002f
C721 VDD.n223 GND 0.008002f
C722 VDD.n224 GND 0.008002f
C723 VDD.n225 GND 0.008002f
C724 VDD.n226 GND 0.00644f
C725 VDD.n227 GND 0.008002f
C726 VDD.n228 GND 0.008002f
C727 VDD.n229 GND 0.008002f
C728 VDD.n230 GND 0.008002f
C729 VDD.n231 GND 0.532804f
C730 VDD.n232 GND 0.008002f
C731 VDD.n233 GND 0.008002f
C732 VDD.n234 GND 0.008002f
C733 VDD.n235 GND 0.008002f
C734 VDD.n236 GND 0.008002f
C735 VDD.n237 GND 0.00644f
C736 VDD.n238 GND 0.008002f
C737 VDD.n239 GND 0.008002f
C738 VDD.n240 GND 0.008002f
C739 VDD.n241 GND 0.008002f
C740 VDD.n242 GND 0.772565f
C741 VDD.n243 GND 0.019459f
C742 VDD.n244 GND 0.008002f
C743 VDD.n245 GND 0.008002f
C744 VDD.n246 GND 0.008002f
C745 VDD.n247 GND 0.00644f
C746 VDD.n248 GND 1.24676f
C747 VDD.n249 GND 0.00644f
C748 VDD.n250 GND 0.008002f
C749 VDD.n251 GND 0.008002f
C750 VDD.n252 GND 0.008002f
C751 VDD.n253 GND 0.008002f
C752 VDD.n254 GND 0.008002f
C753 VDD.n255 GND 0.004347f
C754 VDD.n257 GND 0.008002f
C755 VDD.n258 GND 0.006408f
C756 VDD.t102 GND 0.029464f
C757 VDD.t101 GND 0.049829f
C758 VDD.t100 GND 0.498044f
C759 VDD.n259 GND 0.083391f
C760 VDD.n260 GND 0.066666f
C761 VDD.n261 GND 0.008002f
C762 VDD.n262 GND 0.008002f
C763 VDD.n263 GND 0.00644f
C764 VDD.n265 GND 0.008002f
C765 VDD.n266 GND 0.008002f
C766 VDD.n267 GND 0.008002f
C767 VDD.n268 GND 0.008002f
C768 VDD.n269 GND 0.00644f
C769 VDD.n271 GND 0.008002f
C770 VDD.n272 GND 0.008002f
C771 VDD.n273 GND 0.008002f
C772 VDD.n274 GND 0.004991f
C773 VDD.t47 GND 0.029464f
C774 VDD.t46 GND 0.049829f
C775 VDD.t45 GND 0.498044f
C776 VDD.n275 GND 0.083391f
C777 VDD.n276 GND 0.066666f
C778 VDD.n277 GND 0.008002f
C779 VDD.n278 GND 0.00644f
C780 VDD.n280 GND 0.008002f
C781 VDD.n281 GND 0.00644f
C782 VDD.n282 GND 0.008002f
C783 VDD.n283 GND 0.008002f
C784 VDD.n284 GND 0.008002f
C785 VDD.n285 GND 0.008002f
C786 VDD.n286 GND 0.008002f
C787 VDD.n287 GND 0.00644f
C788 VDD.n289 GND 0.008002f
C789 VDD.n290 GND 0.008002f
C790 VDD.n291 GND 0.008002f
C791 VDD.n292 GND 0.008002f
C792 VDD.n293 GND 0.008002f
C793 VDD.n294 GND 0.00644f
C794 VDD.n296 GND 0.008002f
C795 VDD.n297 GND 0.008002f
C796 VDD.n298 GND 0.008002f
C797 VDD.n299 GND 0.008002f
C798 VDD.n300 GND 0.008002f
C799 VDD.n301 GND 0.00644f
C800 VDD.n303 GND 0.008002f
C801 VDD.n304 GND 0.008002f
C802 VDD.n305 GND 0.008002f
C803 VDD.n306 GND 0.008002f
C804 VDD.n307 GND 0.005378f
C805 VDD.t86 GND 0.029464f
C806 VDD.t85 GND 0.049829f
C807 VDD.t84 GND 0.498044f
C808 VDD.n308 GND 0.083391f
C809 VDD.n309 GND 0.066666f
C810 VDD.n311 GND 0.008002f
C811 VDD.n312 GND 0.008002f
C812 VDD.n313 GND 0.00644f
C813 VDD.n314 GND 0.008002f
C814 VDD.n316 GND 0.008002f
C815 VDD.n317 GND 0.008002f
C816 VDD.n318 GND 0.008002f
C817 VDD.n319 GND 0.008002f
C818 VDD.n320 GND 0.00644f
C819 VDD.n322 GND 0.008002f
C820 VDD.n323 GND 0.008002f
C821 VDD.n324 GND 0.008002f
C822 VDD.n325 GND 0.008002f
C823 VDD.n326 GND 0.01975f
C824 VDD.n328 GND 0.00644f
C825 VDD.n329 GND 0.008002f
C826 VDD.n330 GND 0.00644f
C827 VDD.n331 GND 0.008002f
C828 VDD.n332 GND 0.00644f
C829 VDD.n333 GND 0.008002f
C830 VDD.n334 GND 0.00644f
C831 VDD.n335 GND 0.008002f
C832 VDD.n336 GND 0.00644f
C833 VDD.n337 GND 0.008002f
C834 VDD.n338 GND 0.00644f
C835 VDD.n339 GND 0.008002f
C836 VDD.n340 GND 0.00644f
C837 VDD.n341 GND 0.008002f
C838 VDD.n342 GND 0.00644f
C839 VDD.n343 GND 0.008002f
C840 VDD.n344 GND 0.00644f
C841 VDD.n345 GND 0.008002f
C842 VDD.n346 GND 0.00644f
C843 VDD.n347 GND 0.008002f
C844 VDD.n348 GND 0.008002f
C845 VDD.n349 GND 0.532804f
C846 VDD.n350 GND 0.008002f
C847 VDD.n351 GND 0.00644f
C848 VDD.n352 GND 0.008002f
C849 VDD.n353 GND 0.00644f
C850 VDD.n354 GND 0.008002f
C851 VDD.n355 GND 0.532804f
C852 VDD.n356 GND 0.008002f
C853 VDD.n357 GND 0.00644f
C854 VDD.n358 GND 0.008002f
C855 VDD.n359 GND 0.00644f
C856 VDD.n360 GND 0.008002f
C857 VDD.t143 GND 0.266402f
C858 VDD.n361 GND 0.008002f
C859 VDD.n362 GND 0.00644f
C860 VDD.n363 GND 0.008002f
C861 VDD.n364 GND 0.00644f
C862 VDD.n365 GND 0.008002f
C863 VDD.n366 GND 0.532804f
C864 VDD.n367 GND 0.008002f
C865 VDD.n368 GND 0.00644f
C866 VDD.n369 GND 0.008002f
C867 VDD.n370 GND 0.00644f
C868 VDD.n371 GND 0.008002f
C869 VDD.n372 GND 0.532804f
C870 VDD.n373 GND 0.008002f
C871 VDD.n374 GND 0.00644f
C872 VDD.n375 GND 0.008002f
C873 VDD.n376 GND 0.00644f
C874 VDD.n377 GND 0.008002f
C875 VDD.n378 GND 0.532804f
C876 VDD.n379 GND 0.008002f
C877 VDD.n380 GND 0.00644f
C878 VDD.n381 GND 0.008002f
C879 VDD.n382 GND 0.00644f
C880 VDD.n383 GND 0.008002f
C881 VDD.n384 GND 0.532804f
C882 VDD.n385 GND 0.008002f
C883 VDD.n386 GND 0.00644f
C884 VDD.n387 GND 0.008002f
C885 VDD.n388 GND 0.00644f
C886 VDD.n389 GND 0.008002f
C887 VDD.n390 GND 0.306362f
C888 VDD.n391 GND 0.008002f
C889 VDD.n392 GND 0.00644f
C890 VDD.n393 GND 0.008002f
C891 VDD.n394 GND 0.00644f
C892 VDD.n395 GND 0.008002f
C893 VDD.n396 GND 0.532804f
C894 VDD.t135 GND 0.266402f
C895 VDD.n397 GND 0.008002f
C896 VDD.n398 GND 0.00644f
C897 VDD.n399 GND 0.008002f
C898 VDD.n400 GND 0.00644f
C899 VDD.n401 GND 0.008002f
C900 VDD.n402 GND 0.532804f
C901 VDD.n403 GND 0.008002f
C902 VDD.n404 GND 0.00644f
C903 VDD.n405 GND 0.008002f
C904 VDD.n406 GND 0.00644f
C905 VDD.n407 GND 0.008002f
C906 VDD.n408 GND 0.532804f
C907 VDD.n409 GND 0.008002f
C908 VDD.n410 GND 0.00644f
C909 VDD.n411 GND 0.008002f
C910 VDD.n412 GND 0.00644f
C911 VDD.n413 GND 0.008002f
C912 VDD.n414 GND 0.532804f
C913 VDD.n415 GND 0.008002f
C914 VDD.n416 GND 0.00644f
C915 VDD.n417 GND 0.008002f
C916 VDD.n418 GND 0.00644f
C917 VDD.n419 GND 0.008002f
C918 VDD.n420 GND 0.532804f
C919 VDD.n421 GND 0.008002f
C920 VDD.n422 GND 0.00644f
C921 VDD.n423 GND 0.008002f
C922 VDD.n424 GND 0.00644f
C923 VDD.n425 GND 0.008002f
C924 VDD.n426 GND 0.532804f
C925 VDD.n427 GND 0.008002f
C926 VDD.n428 GND 0.00644f
C927 VDD.n429 GND 0.008002f
C928 VDD.n430 GND 0.00644f
C929 VDD.n431 GND 0.008002f
C930 VDD.t34 GND 0.266402f
C931 VDD.n432 GND 0.008002f
C932 VDD.n433 GND 0.00644f
C933 VDD.n434 GND 0.008002f
C934 VDD.n435 GND 0.00644f
C935 VDD.n436 GND 0.008002f
C936 VDD.n437 GND 0.532804f
C937 VDD.n438 GND 0.008002f
C938 VDD.n439 GND 0.00644f
C939 VDD.n440 GND 0.008002f
C940 VDD.n441 GND 0.00644f
C941 VDD.n442 GND 0.008002f
C942 VDD.n443 GND 0.532804f
C943 VDD.n444 GND 0.008002f
C944 VDD.n445 GND 0.00644f
C945 VDD.n446 GND 0.01975f
C946 VDD.n447 GND 0.01975f
C947 VDD.n448 GND 3.71897f
C948 VDD.n449 GND 0.01975f
C949 VDD.n450 GND 0.008002f
C950 VDD.t75 GND 0.029464f
C951 VDD.t76 GND 0.049829f
C952 VDD.t74 GND 0.498044f
C953 VDD.n451 GND 0.083391f
C954 VDD.n452 GND 0.066666f
C955 VDD.n453 GND 0.00644f
C956 VDD.n454 GND 0.00644f
C957 VDD.n455 GND 0.008002f
C958 VDD.n456 GND 0.00644f
C959 VDD.n457 GND 0.004641f
C960 VDD.n458 GND 0.007362f
C961 VDD.n459 GND 0.027582f
C962 VDD.n460 GND 0.00644f
C963 VDD.n461 GND 0.008002f
C964 VDD.n462 GND 0.005378f
C965 VDD.n463 GND 0.008002f
C966 VDD.n464 GND 0.005378f
C967 VDD.n465 GND 0.008002f
C968 VDD.n466 GND 0.00644f
C969 VDD.n467 GND 0.008002f
C970 VDD.n468 GND 0.00644f
C971 VDD.n469 GND 0.008002f
C972 VDD.n470 GND 0.00644f
C973 VDD.n471 GND 0.008002f
C974 VDD.n472 GND 0.003574f
C975 VDD.n473 GND 0.008002f
C976 VDD.n474 GND 0.00644f
C977 VDD.n475 GND 0.008002f
C978 VDD.n476 GND 0.00644f
C979 VDD.n477 GND 0.008002f
C980 VDD.n478 GND 0.00644f
C981 VDD.n479 GND 0.008002f
C982 VDD.n480 GND 0.00644f
C983 VDD.n481 GND 0.008002f
C984 VDD.t35 GND 0.029464f
C985 VDD.t36 GND 0.049829f
C986 VDD.t33 GND 0.498044f
C987 VDD.n482 GND 0.083391f
C988 VDD.n483 GND 0.066666f
C989 VDD.n484 GND 0.013139f
C990 VDD.n485 GND 0.008002f
C991 VDD.n486 GND 0.00644f
C992 VDD.n487 GND 0.008002f
C993 VDD.n488 GND 0.00644f
C994 VDD.n489 GND 0.008002f
C995 VDD.n490 GND 0.00644f
C996 VDD.n491 GND 0.008002f
C997 VDD.n492 GND 0.006408f
C998 VDD.n493 GND 0.004081f
C999 VDD.n494 GND 0.005441f
C1000 VDD.t25 GND 5.63706f
C1001 VDD.n496 GND 2.51483f
C1002 VDD.n497 GND 0.005441f
C1003 VDD.n498 GND 0.005441f
C1004 VDD.n500 GND 0.005441f
C1005 VDD.t124 GND 0.111051f
C1006 VDD.t123 GND 0.129192f
C1007 VDD.t122 GND 0.629305f
C1008 VDD.n501 GND 0.086428f
C1009 VDD.n502 GND 0.052244f
C1010 VDD.n503 GND 0.007776f
C1011 VDD.n505 GND 0.004841f
C1012 VDD.n506 GND 0.011992f
C1013 VDD.n507 GND 0.005441f
C1014 VDD.n508 GND 0.005441f
C1015 VDD.n509 GND 0.362306f
C1016 VDD.n510 GND 0.005441f
C1017 VDD.t0 GND 0.359642f
C1018 VDD.n511 GND 0.450219f
C1019 VDD.n512 GND 0.005441f
C1020 VDD.n513 GND 0.005441f
C1021 VDD.n514 GND 0.011992f
C1022 VDD.n515 GND 0.005441f
C1023 VDD.n516 GND 0.005441f
C1024 VDD.n517 GND 0.362306f
C1025 VDD.n518 GND 0.005441f
C1026 VDD.n519 GND 0.005441f
C1027 VDD.n520 GND 0.005441f
C1028 VDD.n521 GND 0.005441f
C1029 VDD.n522 GND 0.005441f
C1030 VDD.n523 GND 0.013054f
C1031 VDD.n524 GND 0.005441f
C1032 VDD.n525 GND 0.005441f
C1033 VDD.n527 GND 0.005441f
C1034 VDD.n528 GND 0.005441f
C1035 VDD.n530 GND 0.005441f
C1036 VDD.n531 GND 0.005441f
C1037 VDD.n533 GND 0.005441f
C1038 VDD.n534 GND 0.005441f
C1039 VDD.n536 GND 0.005441f
C1040 VDD.t115 GND 0.111051f
C1041 VDD.t114 GND 0.129192f
C1042 VDD.t112 GND 0.629305f
C1043 VDD.n537 GND 0.086428f
C1044 VDD.n538 GND 0.052244f
C1045 VDD.n539 GND 0.005441f
C1046 VDD.n540 GND 0.005441f
C1047 VDD.n541 GND 0.229106f
C1048 VDD.n542 GND 0.005441f
C1049 VDD.n543 GND 0.005441f
C1050 VDD.n544 GND 0.005441f
C1051 VDD.n545 GND 0.005441f
C1052 VDD.n546 GND 0.005441f
C1053 VDD.n547 GND 0.362306f
C1054 VDD.n548 GND 0.005441f
C1055 VDD.n549 GND 0.005441f
C1056 VDD.t113 GND 0.181153f
C1057 VDD.n550 GND 0.005441f
C1058 VDD.n551 GND 0.005441f
C1059 VDD.n552 GND 0.005441f
C1060 VDD.n553 GND 0.005441f
C1061 VDD.t31 GND 0.181153f
C1062 VDD.n554 GND 0.005441f
C1063 VDD.n555 GND 0.005441f
C1064 VDD.n556 GND 0.005441f
C1065 VDD.n557 GND 0.005441f
C1066 VDD.n558 GND 0.005441f
C1067 VDD.n559 GND 0.362306f
C1068 VDD.n560 GND 0.005441f
C1069 VDD.n561 GND 0.005441f
C1070 VDD.n562 GND 0.327674f
C1071 VDD.n563 GND 0.005441f
C1072 VDD.n564 GND 0.005441f
C1073 VDD.n565 GND 0.005441f
C1074 VDD.n566 GND 0.362306f
C1075 VDD.n567 GND 0.005441f
C1076 VDD.n568 GND 0.005441f
C1077 VDD.n569 GND 0.005441f
C1078 VDD.n570 GND 0.005441f
C1079 VDD.n571 GND 0.005441f
C1080 VDD.n572 GND 0.362306f
C1081 VDD.n573 GND 0.005441f
C1082 VDD.n574 GND 0.005441f
C1083 VDD.n575 GND 0.005441f
C1084 VDD.n576 GND 0.005441f
C1085 VDD.n577 GND 0.005441f
C1086 VDD.n578 GND 0.362306f
C1087 VDD.n579 GND 0.005441f
C1088 VDD.n580 GND 0.005441f
C1089 VDD.n581 GND 0.005441f
C1090 VDD.n582 GND 0.005441f
C1091 VDD.n583 GND 0.005441f
C1092 VDD.t7 GND 0.181153f
C1093 VDD.n584 GND 0.005441f
C1094 VDD.n585 GND 0.005441f
C1095 VDD.n586 GND 0.005441f
C1096 VDD.n587 GND 0.005441f
C1097 VDD.n588 GND 0.005441f
C1098 VDD.n589 GND 0.362306f
C1099 VDD.n590 GND 0.005441f
C1100 VDD.n591 GND 0.005441f
C1101 VDD.t4 GND 0.181153f
C1102 VDD.n592 GND 0.005441f
C1103 VDD.n593 GND 0.005441f
C1104 VDD.n594 GND 0.005441f
C1105 VDD.n595 GND 0.362306f
C1106 VDD.n596 GND 0.005441f
C1107 VDD.n597 GND 0.005441f
C1108 VDD.n598 GND 0.005441f
C1109 VDD.n599 GND 0.005441f
C1110 VDD.n600 GND 0.005441f
C1111 VDD.n601 GND 0.362306f
C1112 VDD.n602 GND 0.005441f
C1113 VDD.n603 GND 0.005441f
C1114 VDD.n604 GND 0.005441f
C1115 VDD.n605 GND 0.005441f
C1116 VDD.n606 GND 0.005441f
C1117 VDD.n607 GND 0.362306f
C1118 VDD.n608 GND 0.005441f
C1119 VDD.n609 GND 0.005441f
C1120 VDD.n610 GND 0.005441f
C1121 VDD.n611 GND 0.005441f
C1122 VDD.n612 GND 0.005441f
C1123 VDD.n613 GND 0.279722f
C1124 VDD.n614 GND 0.005441f
C1125 VDD.n615 GND 0.005441f
C1126 VDD.n616 GND 0.005441f
C1127 VDD.n617 GND 0.005441f
C1128 VDD.n618 GND 0.005441f
C1129 VDD.n619 GND 0.362306f
C1130 VDD.n620 GND 0.005441f
C1131 VDD.n621 GND 0.005441f
C1132 VDD.t14 GND 0.149185f
C1133 VDD.t12 GND 0.082585f
C1134 VDD.n622 GND 0.005441f
C1135 VDD.n623 GND 0.005441f
C1136 VDD.n624 GND 0.005441f
C1137 VDD.n625 GND 0.362306f
C1138 VDD.n626 GND 0.005441f
C1139 VDD.n627 GND 0.005441f
C1140 VDD.n628 GND 0.005441f
C1141 VDD.n629 GND 0.005441f
C1142 VDD.n630 GND 0.005441f
C1143 VDD.n631 GND 0.362306f
C1144 VDD.n632 GND 0.005441f
C1145 VDD.n633 GND 0.005441f
C1146 VDD.n634 GND 0.005441f
C1147 VDD.n635 GND 0.005441f
C1148 VDD.n636 GND 0.005441f
C1149 VDD.n637 GND 0.362306f
C1150 VDD.n638 GND 0.005441f
C1151 VDD.n639 GND 0.005441f
C1152 VDD.n640 GND 0.005441f
C1153 VDD.n641 GND 0.005441f
C1154 VDD.n642 GND 0.005441f
C1155 VDD.n643 GND 0.362306f
C1156 VDD.n644 GND 0.005441f
C1157 VDD.n645 GND 0.005441f
C1158 VDD.n646 GND 0.005441f
C1159 VDD.n647 GND 0.005441f
C1160 VDD.n648 GND 0.005441f
C1161 VDD.t5 GND 0.181153f
C1162 VDD.n649 GND 0.005441f
C1163 VDD.n650 GND 0.005441f
C1164 VDD.n651 GND 0.005441f
C1165 VDD.n652 GND 0.005441f
C1166 VDD.n653 GND 0.005441f
C1167 VDD.n654 GND 0.362306f
C1168 VDD.n655 GND 0.005441f
C1169 VDD.n656 GND 0.005441f
C1170 VDD.n657 GND 0.27173f
C1171 VDD.n658 GND 0.005441f
C1172 VDD.n659 GND 0.005441f
C1173 VDD.n660 GND 0.005441f
C1174 VDD.n661 GND 0.31169f
C1175 VDD.n662 GND 0.005441f
C1176 VDD.n663 GND 0.005441f
C1177 VDD.n664 GND 0.005441f
C1178 VDD.n665 GND 0.005441f
C1179 VDD.n666 GND 0.005441f
C1180 VDD.n667 GND 0.362306f
C1181 VDD.n668 GND 0.005441f
C1182 VDD.n669 GND 0.005441f
C1183 VDD.t180 GND 0.181153f
C1184 VDD.n670 GND 0.005441f
C1185 VDD.n671 GND 0.005441f
C1186 VDD.n672 GND 0.005441f
C1187 VDD.n673 GND 0.362306f
C1188 VDD.n674 GND 0.005441f
C1189 VDD.n675 GND 0.005441f
C1190 VDD.n676 GND 0.005441f
C1191 VDD.n677 GND 0.005441f
C1192 VDD.n678 GND 0.005441f
C1193 VDD.n679 GND 0.213121f
C1194 VDD.n680 GND 0.005441f
C1195 VDD.n681 GND 0.005441f
C1196 VDD.n682 GND 0.005441f
C1197 VDD.n683 GND 0.005441f
C1198 VDD.n684 GND 0.005441f
C1199 VDD.n685 GND 0.362306f
C1200 VDD.n686 GND 0.005441f
C1201 VDD.n687 GND 0.005441f
C1202 VDD.t19 GND 0.181153f
C1203 VDD.n688 GND 0.005441f
C1204 VDD.n689 GND 0.005441f
C1205 VDD.n690 GND 0.005441f
C1206 VDD.n691 GND 0.362306f
C1207 VDD.n692 GND 0.005441f
C1208 VDD.n693 GND 0.005441f
C1209 VDD.n694 GND 0.005441f
C1210 VDD.n695 GND 0.005441f
C1211 VDD.n696 GND 0.005441f
C1212 VDD.t27 GND 0.181153f
C1213 VDD.n697 GND 0.005441f
C1214 VDD.n698 GND 0.005441f
C1215 VDD.n699 GND 0.005441f
C1216 VDD.n700 GND 0.005441f
C1217 VDD.n701 GND 0.005441f
C1218 VDD.n702 GND 0.362306f
C1219 VDD.n703 GND 0.005441f
C1220 VDD.n704 GND 0.005441f
C1221 VDD.n705 GND 0.290378f
C1222 VDD.n706 GND 0.005441f
C1223 VDD.n707 GND 0.005441f
C1224 VDD.n708 GND 0.005441f
C1225 VDD.n709 GND 0.335666f
C1226 VDD.n710 GND 0.005441f
C1227 VDD.n711 GND 0.005441f
C1228 VDD.n712 GND 0.005441f
C1229 VDD.n713 GND 0.005441f
C1230 VDD.n714 GND 0.005441f
C1231 VDD.n715 GND 0.362306f
C1232 VDD.n716 GND 0.005441f
C1233 VDD.n717 GND 0.005441f
C1234 VDD.t177 GND 0.181153f
C1235 VDD.n718 GND 0.005441f
C1236 VDD.n719 GND 0.005441f
C1237 VDD.n720 GND 0.005441f
C1238 VDD.n721 GND 0.362306f
C1239 VDD.n722 GND 0.005441f
C1240 VDD.n723 GND 0.005441f
C1241 VDD.n724 GND 0.005441f
C1242 VDD.n725 GND 0.005441f
C1243 VDD.n726 GND 0.005441f
C1244 VDD.n727 GND 0.194473f
C1245 VDD.n728 GND 0.005441f
C1246 VDD.n729 GND 0.005441f
C1247 VDD.n730 GND 0.005441f
C1248 VDD.n731 GND 0.005441f
C1249 VDD.n732 GND 0.005441f
C1250 VDD.n733 GND 0.362306f
C1251 VDD.n734 GND 0.005441f
C1252 VDD.n735 GND 0.005441f
C1253 VDD.t29 GND 0.181153f
C1254 VDD.n736 GND 0.005441f
C1255 VDD.n737 GND 0.005441f
C1256 VDD.n738 GND 0.005441f
C1257 VDD.n739 GND 0.362306f
C1258 VDD.n740 GND 0.005441f
C1259 VDD.n741 GND 0.005441f
C1260 VDD.n742 GND 0.005441f
C1261 VDD.n743 GND 0.005441f
C1262 VDD.n744 GND 0.005441f
C1263 VDD.n745 GND 0.362306f
C1264 VDD.n746 GND 0.005441f
C1265 VDD.n747 GND 0.005441f
C1266 VDD.n748 GND 0.005441f
C1267 VDD.n749 GND 0.005441f
C1268 VDD.n750 GND 0.005441f
C1269 VDD.n751 GND 0.314354f
C1270 VDD.n752 GND 0.005441f
C1271 VDD.n753 GND 0.005441f
C1272 VDD.n754 GND 0.005441f
C1273 VDD.n755 GND 0.005441f
C1274 VDD.n756 GND 0.005441f
C1275 VDD.n757 GND 0.317018f
C1276 VDD.n758 GND 0.005441f
C1277 VDD.n759 GND 0.005441f
C1278 VDD.t88 GND 0.181153f
C1279 VDD.n760 GND 0.005441f
C1280 VDD.n761 GND 0.005441f
C1281 VDD.n762 GND 0.005441f
C1282 VDD.n763 GND 0.362306f
C1283 VDD.n764 GND 0.005441f
C1284 VDD.n765 GND 0.005441f
C1285 VDD.t125 GND 0.181153f
C1286 VDD.n766 GND 0.005441f
C1287 VDD.n767 GND 0.005441f
C1288 VDD.n768 GND 0.005441f
C1289 VDD.n769 GND 0.362306f
C1290 VDD.n770 GND 0.005441f
C1291 VDD.n771 GND 0.005441f
C1292 VDD.n772 GND 0.005441f
C1293 VDD.n773 GND 0.013054f
C1294 VDD.n774 GND 0.013054f
C1295 VDD.n775 GND 0.540796f
C1296 VDD.n797 GND 0.013054f
C1297 VDD.n798 GND 0.011992f
C1298 VDD.n799 GND 0.005441f
C1299 VDD.n800 GND 0.011992f
C1300 VDD.t73 GND 0.111051f
C1301 VDD.t72 GND 0.129192f
C1302 VDD.t71 GND 0.629305f
C1303 VDD.n801 GND 0.086428f
C1304 VDD.n802 GND 0.052244f
C1305 VDD.n803 GND 0.005441f
C1306 VDD.n804 GND 0.005441f
C1307 VDD.n805 GND 0.362306f
C1308 VDD.n806 GND 0.005441f
C1309 VDD.n807 GND 0.005441f
C1310 VDD.n808 GND 0.005441f
C1311 VDD.n809 GND 0.011992f
C1312 VDD.n810 GND 0.005441f
C1313 VDD.t64 GND 0.111051f
C1314 VDD.t63 GND 0.129192f
C1315 VDD.t61 GND 0.629305f
C1316 VDD.n811 GND 0.086428f
C1317 VDD.n812 GND 0.052244f
C1318 VDD.n813 GND 0.007776f
C1319 VDD.n814 GND 0.005441f
C1320 VDD.n815 GND 0.005441f
C1321 VDD.n816 GND 0.226442f
C1322 VDD.n817 GND 0.005441f
C1323 VDD.n818 GND 0.005441f
C1324 VDD.n819 GND 0.005441f
C1325 VDD.n820 GND 0.005441f
C1326 VDD.n821 GND 0.005441f
C1327 VDD.n822 GND 0.229106f
C1328 VDD.n823 GND 0.005441f
C1329 VDD.n824 GND 0.005441f
C1330 VDD.t16 GND 0.181153f
C1331 VDD.n825 GND 0.005441f
C1332 VDD.n826 GND 0.005441f
C1333 VDD.n827 GND 0.005441f
C1334 VDD.n828 GND 0.005441f
C1335 VDD.n829 GND 0.362306f
C1336 VDD.n830 GND 0.005441f
C1337 VDD.n831 GND 0.005441f
C1338 VDD.t62 GND 0.181153f
C1339 VDD.n832 GND 0.005441f
C1340 VDD.n833 GND 0.005441f
C1341 VDD.n834 GND 0.005441f
C1342 VDD.n835 GND 0.362306f
C1343 VDD.n836 GND 0.005441f
C1344 VDD.n837 GND 0.005441f
C1345 VDD.n838 GND 0.005441f
C1346 VDD.n839 GND 0.005441f
C1347 VDD.n840 GND 0.005441f
C1348 VDD.n841 GND 0.362306f
C1349 VDD.n842 GND 0.005441f
C1350 VDD.n843 GND 0.005441f
C1351 VDD.n844 GND 0.005441f
C1352 VDD.n845 GND 0.005441f
C1353 VDD.n846 GND 0.005441f
C1354 VDD.n847 GND 0.348986f
C1355 VDD.n848 GND 0.005441f
C1356 VDD.n849 GND 0.005441f
C1357 VDD.n850 GND 0.005441f
C1358 VDD.n851 GND 0.005441f
C1359 VDD.n852 GND 0.005441f
C1360 VDD.n853 GND 0.362306f
C1361 VDD.n854 GND 0.005441f
C1362 VDD.n855 GND 0.005441f
C1363 VDD.t2 GND 0.181153f
C1364 VDD.n856 GND 0.005441f
C1365 VDD.n857 GND 0.005441f
C1366 VDD.n858 GND 0.005441f
C1367 VDD.n859 GND 0.362306f
C1368 VDD.n860 GND 0.005441f
C1369 VDD.n861 GND 0.005441f
C1370 VDD.n862 GND 0.005441f
C1371 VDD.n863 GND 0.005441f
C1372 VDD.n864 GND 0.005441f
C1373 VDD.n865 GND 0.207793f
C1374 VDD.n866 GND 0.005441f
C1375 VDD.n867 GND 0.005441f
C1376 VDD.n868 GND 0.005441f
C1377 VDD.n869 GND 0.005441f
C1378 VDD.n870 GND 0.005441f
C1379 VDD.n871 GND 0.362306f
C1380 VDD.n872 GND 0.005441f
C1381 VDD.n873 GND 0.005441f
C1382 VDD.t18 GND 0.181153f
C1383 VDD.n874 GND 0.005441f
C1384 VDD.n875 GND 0.005441f
C1385 VDD.n876 GND 0.005441f
C1386 VDD.n877 GND 0.362306f
C1387 VDD.n878 GND 0.005441f
C1388 VDD.n879 GND 0.005441f
C1389 VDD.n880 GND 0.005441f
C1390 VDD.n881 GND 0.005441f
C1391 VDD.n882 GND 0.005441f
C1392 VDD.t23 GND 0.181153f
C1393 VDD.n883 GND 0.005441f
C1394 VDD.n884 GND 0.005441f
C1395 VDD.n885 GND 0.005441f
C1396 VDD.n886 GND 0.005441f
C1397 VDD.n887 GND 0.005441f
C1398 VDD.n888 GND 0.362306f
C1399 VDD.n889 GND 0.005441f
C1400 VDD.n890 GND 0.005441f
C1401 VDD.n891 GND 0.253082f
C1402 VDD.n892 GND 0.005441f
C1403 VDD.n893 GND 0.005441f
C1404 VDD.n894 GND 0.005441f
C1405 VDD.n895 GND 0.330338f
C1406 VDD.n896 GND 0.005441f
C1407 VDD.n897 GND 0.005441f
C1408 VDD.n898 GND 0.005441f
C1409 VDD.n899 GND 0.005441f
C1410 VDD.n900 GND 0.005441f
C1411 VDD.n901 GND 0.362306f
C1412 VDD.n902 GND 0.005441f
C1413 VDD.n903 GND 0.005441f
C1414 VDD.t6 GND 0.181153f
C1415 VDD.n904 GND 0.005441f
C1416 VDD.n905 GND 0.005441f
C1417 VDD.n906 GND 0.005441f
C1418 VDD.n907 GND 0.362306f
C1419 VDD.n908 GND 0.005441f
C1420 VDD.n909 GND 0.005441f
C1421 VDD.n910 GND 0.005441f
C1422 VDD.n911 GND 0.005441f
C1423 VDD.n912 GND 0.005441f
C1424 VDD.n913 GND 0.23177f
C1425 VDD.n914 GND 0.005441f
C1426 VDD.n915 GND 0.005441f
C1427 VDD.n916 GND 0.005441f
C1428 VDD.n917 GND 0.005441f
C1429 VDD.n918 GND 0.005441f
C1430 VDD.n919 GND 0.362306f
C1431 VDD.n920 GND 0.005441f
C1432 VDD.n921 GND 0.005441f
C1433 VDD.t10 GND 0.181153f
C1434 VDD.n922 GND 0.005441f
C1435 VDD.n923 GND 0.005441f
C1436 VDD.n924 GND 0.005441f
C1437 VDD.n925 GND 0.362306f
C1438 VDD.n926 GND 0.005441f
C1439 VDD.n927 GND 0.005441f
C1440 VDD.n928 GND 0.005441f
C1441 VDD.n929 GND 0.005441f
C1442 VDD.n930 GND 0.005441f
C1443 VDD.t13 GND 0.181153f
C1444 VDD.n931 GND 0.005441f
C1445 VDD.n932 GND 0.005441f
C1446 VDD.n933 GND 0.005441f
C1447 VDD.n934 GND 0.005441f
C1448 VDD.n935 GND 0.005441f
C1449 VDD.n936 GND 0.362306f
C1450 VDD.n937 GND 0.005441f
C1451 VDD.n938 GND 0.005441f
C1452 VDD.n939 GND 0.27173f
C1453 VDD.n940 GND 0.005441f
C1454 VDD.n941 GND 0.005441f
C1455 VDD.n942 GND 0.005441f
C1456 VDD.n943 GND 0.362306f
C1457 VDD.n944 GND 0.005441f
C1458 VDD.n945 GND 0.005441f
C1459 VDD.n946 GND 0.005441f
C1460 VDD.n947 GND 0.005441f
C1461 VDD.n948 GND 0.005441f
C1462 VDD.n949 GND 0.362306f
C1463 VDD.n950 GND 0.005441f
C1464 VDD.n951 GND 0.005441f
C1465 VDD.n952 GND 0.005441f
C1466 VDD.n953 GND 0.005441f
C1467 VDD.n954 GND 0.005441f
C1468 VDD.n955 GND 0.362306f
C1469 VDD.n956 GND 0.005441f
C1470 VDD.n957 GND 0.005441f
C1471 VDD.n958 GND 0.005441f
C1472 VDD.n959 GND 0.005441f
C1473 VDD.n960 GND 0.005441f
C1474 VDD.n961 GND 0.213121f
C1475 VDD.n962 GND 0.005441f
C1476 VDD.n963 GND 0.005441f
C1477 VDD.n964 GND 0.005441f
C1478 VDD.n965 GND 0.005441f
C1479 VDD.n966 GND 0.005441f
C1480 VDD.n967 GND 0.362306f
C1481 VDD.n968 GND 0.005441f
C1482 VDD.n969 GND 0.005441f
C1483 VDD.t9 GND 0.082585f
C1484 VDD.t178 GND 0.149185f
C1485 VDD.n970 GND 0.005441f
C1486 VDD.n971 GND 0.005441f
C1487 VDD.n972 GND 0.005441f
C1488 VDD.n973 GND 0.362306f
C1489 VDD.n974 GND 0.005441f
C1490 VDD.n975 GND 0.005441f
C1491 VDD.n976 GND 0.005441f
C1492 VDD.n977 GND 0.005441f
C1493 VDD.n978 GND 0.005441f
C1494 VDD.n979 GND 0.362306f
C1495 VDD.n980 GND 0.005441f
C1496 VDD.n981 GND 0.005441f
C1497 VDD.n982 GND 0.005441f
C1498 VDD.n983 GND 0.005441f
C1499 VDD.n984 GND 0.005441f
C1500 VDD.n985 GND 0.362306f
C1501 VDD.n986 GND 0.005441f
C1502 VDD.n987 GND 0.005441f
C1503 VDD.n988 GND 0.005441f
C1504 VDD.n989 GND 0.005441f
C1505 VDD.n990 GND 0.005441f
C1506 VDD.n991 GND 0.335666f
C1507 VDD.n992 GND 0.005441f
C1508 VDD.n993 GND 0.005441f
C1509 VDD.n994 GND 0.005441f
C1510 VDD.n995 GND 0.005441f
C1511 VDD.n996 GND 0.005441f
C1512 VDD.t21 GND 0.181153f
C1513 VDD.n997 GND 0.005441f
C1514 VDD.n998 GND 0.005441f
C1515 VDD.t20 GND 0.181153f
C1516 VDD.n999 GND 0.005441f
C1517 VDD.n1000 GND 0.005441f
C1518 VDD.n1001 GND 0.005441f
C1519 VDD.n1002 GND 0.362306f
C1520 VDD.n1003 GND 0.005441f
C1521 VDD.n1004 GND 0.005441f
C1522 VDD.n1005 GND 0.33833f
C1523 VDD.n1006 GND 0.005441f
C1524 VDD.n1007 GND 0.005441f
C1525 VDD.n1008 GND 0.005441f
C1526 VDD.n1009 GND 0.362306f
C1527 VDD.n1010 GND 0.005441f
C1528 VDD.n1011 GND 0.005441f
C1529 VDD.n1012 GND 0.005441f
C1530 VDD.n1013 GND 0.005441f
C1531 VDD.n1014 GND 0.005441f
C1532 VDD.n1015 GND 0.362306f
C1533 VDD.n1016 GND 0.005441f
C1534 VDD.n1017 GND 0.005441f
C1535 VDD.n1018 GND 0.005441f
C1536 VDD.n1019 GND 0.005441f
C1537 VDD.n1020 GND 0.005441f
C1538 VDD.n1021 GND 0.362306f
C1539 VDD.n1022 GND 0.005441f
C1540 VDD.n1023 GND 0.005441f
C1541 VDD.n1024 GND 0.005441f
C1542 VDD.n1025 GND 0.005441f
C1543 VDD.n1026 GND 0.005441f
C1544 VDD.t175 GND 0.181153f
C1545 VDD.n1027 GND 0.005441f
C1546 VDD.n1028 GND 0.005441f
C1547 VDD.n1029 GND 0.005441f
C1548 VDD.n1030 GND 0.005441f
C1549 VDD.n1031 GND 0.005441f
C1550 VDD.n1032 GND 0.314354f
C1551 VDD.n1033 GND 0.005441f
C1552 VDD.n1034 GND 0.005441f
C1553 VDD.n1035 GND 0.215785f
C1554 VDD.n1036 GND 0.005441f
C1555 VDD.n1037 GND 0.005441f
C1556 VDD.n1038 GND 0.005441f
C1557 VDD.n1039 GND 0.362306f
C1558 VDD.n1040 GND 0.005441f
C1559 VDD.n1041 GND 0.005441f
C1560 VDD.t81 GND 0.181153f
C1561 VDD.n1042 GND 0.005441f
C1562 VDD.n1043 GND 0.005441f
C1563 VDD.n1044 GND 0.005441f
C1564 VDD.n1045 GND 0.362306f
C1565 VDD.n1046 GND 0.005441f
C1566 VDD.n1047 GND 0.005441f
C1567 VDD.n1048 GND 0.005441f
C1568 VDD.n1049 GND 0.005441f
C1569 VDD.n1050 GND 0.005441f
C1570 VDD.n1051 GND 0.362306f
C1571 VDD.n1052 GND 0.005441f
C1572 VDD.n1053 GND 0.005441f
C1573 VDD.n1054 GND 0.005441f
C1574 VDD.n1055 GND 0.013054f
C1575 VDD.n1056 GND 0.013054f
C1576 VDD.t182 GND 0.359642f
C1577 VDD.n1057 GND 0.011992f
C1578 VDD.n1058 GND 0.011992f
C1579 VDD.n1059 GND 0.013054f
C1580 VDD.n1060 GND 0.005441f
C1581 VDD.n1061 GND 0.005441f
C1582 VDD.t26 GND 5.63706f
C1583 VDD.n1071 GND 0.013054f
C1584 VDD.n1082 GND 0.005441f
C1585 VDD.t117 GND 0.111051f
C1586 VDD.t118 GND 0.129192f
C1587 VDD.t116 GND 0.629305f
C1588 VDD.n1083 GND 0.086428f
C1589 VDD.n1084 GND 0.052244f
C1590 VDD.n1085 GND 0.004641f
C1591 VDD.n1088 GND 0.008002f
C1592 VDD.n1089 GND 0.00644f
C1593 VDD.n1090 GND 0.008002f
C1594 VDD.n1091 GND 0.008002f
C1595 VDD.n1092 GND 0.01975f
C1596 VDD.n1093 GND 0.008002f
C1597 VDD.n1094 GND 0.00644f
C1598 VDD.n1095 GND 0.008002f
C1599 VDD.n1096 GND 0.532804f
C1600 VDD.n1098 GND 3.71897f
C1601 VDD.n1099 GND 0.008002f
C1602 VDD.n1100 GND 0.01975f
C1603 VDD.n1101 GND 0.00644f
C1604 VDD.n1102 GND 0.008002f
C1605 VDD.n1103 GND 0.00644f
C1606 VDD.n1104 GND 0.008002f
C1607 VDD.n1105 GND 0.532804f
C1608 VDD.n1106 GND 0.008002f
C1609 VDD.n1107 GND 0.00644f
C1610 VDD.n1108 GND 0.008002f
C1611 VDD.n1109 GND 0.00644f
C1612 VDD.n1110 GND 0.008002f
C1613 VDD.n1111 GND 0.418251f
C1614 VDD.n1112 GND 0.008002f
C1615 VDD.n1113 GND 0.00644f
C1616 VDD.n1114 GND 0.008002f
C1617 VDD.n1115 GND 0.00644f
C1618 VDD.n1116 GND 0.008002f
C1619 VDD.n1117 GND 0.532804f
C1620 VDD.n1118 GND 0.008002f
C1621 VDD.n1119 GND 0.00644f
C1622 VDD.n1120 GND 0.008002f
C1623 VDD.n1121 GND 0.00644f
C1624 VDD.n1122 GND 0.008002f
C1625 VDD.n1123 GND 0.532804f
C1626 VDD.n1124 GND 0.008002f
C1627 VDD.n1125 GND 0.00644f
C1628 VDD.n1126 GND 0.008002f
C1629 VDD.n1127 GND 0.00644f
C1630 VDD.n1128 GND 0.008002f
C1631 VDD.n1129 GND 0.532804f
C1632 VDD.n1130 GND 0.008002f
C1633 VDD.n1131 GND 0.00644f
C1634 VDD.n1132 GND 0.008002f
C1635 VDD.n1133 GND 0.00644f
C1636 VDD.n1134 GND 0.008002f
C1637 VDD.n1135 GND 0.532804f
C1638 VDD.n1136 GND 0.008002f
C1639 VDD.n1137 GND 0.00644f
C1640 VDD.n1138 GND 0.008002f
C1641 VDD.n1139 GND 0.00644f
C1642 VDD.n1140 GND 0.008002f
C1643 VDD.n1141 GND 0.532804f
C1644 VDD.n1142 GND 0.008002f
C1645 VDD.n1143 GND 0.00644f
C1646 VDD.n1144 GND 0.008002f
C1647 VDD.n1145 GND 0.00644f
C1648 VDD.n1146 GND 0.008002f
C1649 VDD.n1147 GND 0.532804f
C1650 VDD.n1148 GND 0.008002f
C1651 VDD.n1149 GND 0.00644f
C1652 VDD.n1150 GND 0.008002f
C1653 VDD.n1151 GND 0.00644f
C1654 VDD.n1152 GND 0.008002f
C1655 VDD.t131 GND 0.266402f
C1656 VDD.n1153 GND 0.008002f
C1657 VDD.n1154 GND 0.00644f
C1658 VDD.n1155 GND 0.008002f
C1659 VDD.n1156 GND 0.00644f
C1660 VDD.n1157 GND 0.008002f
C1661 VDD.n1158 GND 0.532804f
C1662 VDD.n1159 GND 0.306362f
C1663 VDD.n1160 GND 0.008002f
C1664 VDD.n1161 GND 0.00644f
C1665 VDD.n1162 GND 0.008002f
C1666 VDD.n1163 GND 0.00644f
C1667 VDD.n1164 GND 0.008002f
C1668 VDD.n1165 GND 0.532804f
C1669 VDD.n1166 GND 0.008002f
C1670 VDD.n1167 GND 0.00644f
C1671 VDD.n1168 GND 0.008002f
C1672 VDD.n1169 GND 0.00644f
C1673 VDD.n1170 GND 0.008002f
C1674 VDD.n1171 GND 0.532804f
C1675 VDD.n1172 GND 0.008002f
C1676 VDD.n1173 GND 0.00644f
C1677 VDD.n1174 GND 0.008002f
C1678 VDD.n1175 GND 0.00644f
C1679 VDD.n1176 GND 0.008002f
C1680 VDD.n1177 GND 0.532804f
C1681 VDD.n1178 GND 0.008002f
C1682 VDD.n1179 GND 0.00644f
C1683 VDD.n1180 GND 0.008002f
C1684 VDD.n1181 GND 0.00644f
C1685 VDD.n1182 GND 0.008002f
C1686 VDD.n1183 GND 0.519484f
C1687 VDD.n1184 GND 0.008002f
C1688 VDD.n1185 GND 0.00644f
C1689 VDD.n1186 GND 0.008002f
C1690 VDD.n1187 GND 0.00644f
C1691 VDD.n1188 GND 0.008002f
C1692 VDD.n1189 GND 0.532804f
C1693 VDD.n1190 GND 0.008002f
C1694 VDD.n1191 GND 0.00644f
C1695 VDD.n1192 GND 0.008002f
C1696 VDD.n1193 GND 0.00644f
C1697 VDD.n1194 GND 0.008002f
C1698 VDD.n1195 GND 0.532804f
C1699 VDD.n1196 GND 0.008002f
C1700 VDD.n1197 GND 0.00644f
C1701 VDD.n1198 GND 0.00615f
C1702 VDD.n1199 GND 0.00644f
C1703 VDD.n1200 GND 0.008002f
C1704 VDD.n1201 GND 0.532804f
C1705 VDD.n1202 GND 0.008002f
C1706 VDD.n1203 GND 0.00644f
C1707 VDD.n1204 GND 0.008002f
C1708 VDD.n1205 GND 0.00644f
C1709 VDD.n1206 GND 0.008002f
C1710 VDD.n1207 GND 0.532804f
C1711 VDD.n1208 GND 0.008002f
C1712 VDD.n1209 GND 0.00644f
C1713 VDD.n1210 GND 0.008002f
C1714 VDD.n1211 GND 0.00644f
C1715 VDD.n1212 GND 0.008002f
C1716 VDD.n1213 GND 0.532804f
C1717 VDD.n1214 GND 0.008002f
C1718 VDD.n1215 GND 0.00644f
C1719 VDD.n1216 GND 0.008002f
C1720 VDD.n1217 GND 0.00644f
C1721 VDD.n1218 GND 0.008002f
C1722 VDD.n1219 GND 0.279722f
C1723 VDD.n1220 GND 0.008002f
C1724 VDD.n1221 GND 0.00644f
C1725 VDD.n1222 GND 0.008002f
C1726 VDD.n1223 GND 0.00644f
C1727 VDD.n1224 GND 0.008002f
C1728 VDD.n1225 GND 0.532804f
C1729 VDD.n1226 GND 0.008002f
C1730 VDD.n1227 GND 0.00644f
C1731 VDD.n1228 GND 0.008002f
C1732 VDD.n1229 GND 0.00644f
C1733 VDD.n1230 GND 0.008002f
C1734 VDD.n1231 GND 0.532804f
C1735 VDD.n1232 GND 0.008002f
C1736 VDD.n1233 GND 0.00644f
C1737 VDD.n1234 GND 0.008002f
C1738 VDD.n1235 GND 0.00644f
C1739 VDD.n1236 GND 0.008002f
C1740 VDD.n1237 GND 0.532804f
C1741 VDD.n1238 GND 0.008002f
C1742 VDD.n1239 GND 0.00644f
C1743 VDD.n1240 GND 0.008002f
C1744 VDD.n1241 GND 0.00644f
C1745 VDD.n1242 GND 0.008002f
C1746 VDD.n1243 GND 0.532804f
C1747 VDD.n1244 GND 0.008002f
C1748 VDD.n1245 GND 0.00644f
C1749 VDD.n1246 GND 0.008002f
C1750 VDD.n1247 GND 0.00644f
C1751 VDD.n1248 GND 0.008002f
C1752 VDD.n1249 GND 0.532804f
C1753 VDD.n1250 GND 0.008002f
C1754 VDD.n1251 GND 0.00644f
C1755 VDD.n1252 GND 0.008002f
C1756 VDD.n1253 GND 0.00644f
C1757 VDD.n1254 GND 0.008002f
C1758 VDD.t129 GND 0.266402f
C1759 VDD.n1255 GND 0.008002f
C1760 VDD.n1256 GND 0.00644f
C1761 VDD.n1257 GND 0.008002f
C1762 VDD.n1258 GND 0.00644f
C1763 VDD.n1259 GND 0.008002f
C1764 VDD.n1260 GND 0.532804f
C1765 VDD.n1261 GND 0.008002f
C1766 VDD.n1262 GND 0.00644f
C1767 VDD.n1263 GND 0.008002f
C1768 VDD.n1264 GND 0.00644f
C1769 VDD.n1265 GND 0.008002f
C1770 VDD.n1266 GND 0.532804f
C1771 VDD.n1267 GND 0.008002f
C1772 VDD.n1268 GND 0.00644f
C1773 VDD.n1269 GND 0.008002f
C1774 VDD.n1270 GND 0.00644f
C1775 VDD.n1271 GND 0.008002f
C1776 VDD.n1272 GND 0.532804f
C1777 VDD.n1273 GND 0.008002f
C1778 VDD.n1274 GND 0.00644f
C1779 VDD.n1275 GND 0.008002f
C1780 VDD.n1276 GND 0.00644f
C1781 VDD.n1277 GND 0.008002f
C1782 VDD.n1278 GND 0.532804f
C1783 VDD.n1279 GND 0.008002f
C1784 VDD.n1280 GND 0.00644f
C1785 VDD.n1281 GND 0.008002f
C1786 VDD.n1282 GND 0.00644f
C1787 VDD.n1283 GND 0.008002f
C1788 VDD.n1284 GND 0.532804f
C1789 VDD.n1285 GND 0.008002f
C1790 VDD.n1286 GND 0.00644f
C1791 VDD.n1287 GND 0.008002f
C1792 VDD.n1288 GND 0.00644f
C1793 VDD.n1289 GND 0.008002f
C1794 VDD.n1290 GND 0.380955f
C1795 VDD.n1291 GND 0.008002f
C1796 VDD.n1292 GND 0.00644f
C1797 VDD.n1293 GND 0.008002f
C1798 VDD.n1294 GND 0.00644f
C1799 VDD.n1295 GND 0.008002f
C1800 VDD.n1296 GND 0.532804f
C1801 VDD.n1297 GND 0.008002f
C1802 VDD.n1298 GND 0.00644f
C1803 VDD.n1299 GND 0.008002f
C1804 VDD.n1300 GND 0.00644f
C1805 VDD.n1301 GND 0.008002f
C1806 VDD.n1302 GND 0.532804f
C1807 VDD.n1303 GND 0.008002f
C1808 VDD.n1304 GND 0.00644f
C1809 VDD.n1305 GND 0.019459f
C1810 VDD.n1306 GND 0.005346f
C1811 VDD.n1307 GND 0.019459f
C1812 VDD.n1308 GND 0.772565f
C1813 VDD.n1309 GND 0.019459f
C1814 VDD.n1310 GND 0.005346f
C1815 VDD.n1311 GND 0.008002f
C1816 VDD.t56 GND 0.029464f
C1817 VDD.t57 GND 0.049829f
C1818 VDD.t55 GND 0.498044f
C1819 VDD.n1312 GND 0.083391f
C1820 VDD.n1313 GND 0.066666f
C1821 VDD.n1314 GND 0.009918f
C1822 VDD.n1315 GND 0.008002f
C1823 VDD.n1337 GND 0.008002f
C1824 VDD.n1338 GND 0.008002f
C1825 VDD.n1339 GND 0.01975f
C1826 VDD.n1340 GND 0.00644f
C1827 VDD.n1341 GND 0.008002f
C1828 VDD.n1342 GND 0.008002f
C1829 VDD.n1343 GND 0.008002f
C1830 VDD.n1344 GND 0.008002f
C1831 VDD.n1345 GND 0.004347f
C1832 VDD.n1346 GND 0.008002f
C1833 VDD.n1347 GND 0.008002f
C1834 VDD.n1348 GND 0.008002f
C1835 VDD.n1349 GND 0.00644f
C1836 VDD.n1350 GND 0.008002f
C1837 VDD.n1351 GND 0.008002f
C1838 VDD.n1352 GND 0.008002f
C1839 VDD.n1353 GND 0.008002f
C1840 VDD.n1354 GND 0.008002f
C1841 VDD.n1355 GND 0.00644f
C1842 VDD.n1356 GND 0.008002f
C1843 VDD.n1357 GND 0.008002f
C1844 VDD.n1358 GND 0.008002f
C1845 VDD.n1359 GND 0.00644f
C1846 VDD.n1360 GND 0.008002f
C1847 VDD.n1361 GND 0.008002f
C1848 VDD.n1362 GND 0.008002f
C1849 VDD.n1363 GND 0.008002f
C1850 VDD.n1364 GND 0.008002f
C1851 VDD.n1365 GND 0.00644f
C1852 VDD.n1366 GND 0.008002f
C1853 VDD.n1367 GND 0.008002f
C1854 VDD.n1368 GND 0.008002f
C1855 VDD.n1369 GND 0.008002f
C1856 VDD.n1370 GND 0.008002f
C1857 VDD.t69 GND 0.029464f
C1858 VDD.t70 GND 0.049829f
C1859 VDD.t68 GND 0.498044f
C1860 VDD.n1371 GND 0.083391f
C1861 VDD.n1372 GND 0.066666f
C1862 VDD.n1373 GND 0.009918f
C1863 VDD.n1374 GND 0.008002f
C1864 VDD.n1375 GND 0.008002f
C1865 VDD.n1376 GND 0.008002f
C1866 VDD.n1377 GND 0.008002f
C1867 VDD.n1378 GND 0.008002f
C1868 VDD.n1379 GND 0.00644f
C1869 VDD.n1380 GND 0.008002f
C1870 VDD.n1381 GND 0.008002f
C1871 VDD.n1382 GND 0.008002f
C1872 VDD.n1383 GND 0.008002f
C1873 VDD.n1384 GND 0.008002f
C1874 VDD.n1385 GND 0.00644f
C1875 VDD.n1386 GND 0.008002f
C1876 VDD.n1387 GND 0.008002f
C1877 VDD.n1388 GND 0.008002f
C1878 VDD.n1389 GND 0.008002f
C1879 VDD.n1390 GND 0.00644f
C1880 VDD.n1391 GND 0.008002f
C1881 VDD.n1392 GND 0.008002f
C1882 VDD.n1393 GND 0.008002f
C1883 VDD.n1394 GND 0.008002f
C1884 VDD.n1395 GND 0.008002f
C1885 VDD.n1396 GND 0.00644f
C1886 VDD.n1397 GND 0.008002f
C1887 VDD.n1398 GND 0.008002f
C1888 VDD.n1399 GND 0.008002f
C1889 VDD.n1400 GND 0.003574f
C1890 VDD.n1401 GND 0.00644f
C1891 VDD.n1402 GND 0.00644f
C1892 VDD.n1403 GND 0.008002f
C1893 VDD.n1404 GND 0.008002f
C1894 VDD.n1405 GND 0.008002f
C1895 VDD.n1406 GND 0.00644f
C1896 VDD.n1407 GND 0.00644f
C1897 VDD.n1408 GND 0.00644f
C1898 VDD.n1409 GND 0.008002f
C1899 VDD.n1410 GND 0.008002f
C1900 VDD.n1411 GND 0.008002f
C1901 VDD.n1412 GND 0.005378f
C1902 VDD.n1413 GND 0.008002f
C1903 VDD.t107 GND 0.029464f
C1904 VDD.t108 GND 0.049829f
C1905 VDD.t106 GND 0.498044f
C1906 VDD.n1414 GND 0.083391f
C1907 VDD.n1415 GND 0.066666f
C1908 VDD.n1416 GND 0.013139f
C1909 VDD.n1417 GND 0.005378f
C1910 VDD.n1418 GND 0.008002f
C1911 VDD.n1419 GND 0.008002f
C1912 VDD.n1420 GND 0.008002f
C1913 VDD.n1421 GND 0.00644f
C1914 VDD.n1422 GND 0.00644f
C1915 VDD.n1423 GND 0.00644f
C1916 VDD.n1424 GND 0.008002f
C1917 VDD.n1425 GND 0.008002f
C1918 VDD.n1426 GND 0.008002f
C1919 VDD.n1427 GND 0.00644f
C1920 VDD.n1428 GND 0.00644f
C1921 VDD.n1429 GND 0.003574f
C1922 VDD.n1430 GND 0.008002f
C1923 VDD.n1431 GND 0.008002f
C1924 VDD.n1432 GND 0.003961f
C1925 VDD.n1433 GND 0.00644f
C1926 VDD.n1434 GND 0.00644f
C1927 VDD.n1435 GND 0.008002f
C1928 VDD.n1436 GND 0.008002f
C1929 VDD.n1437 GND 0.008002f
C1930 VDD.n1438 GND 0.00644f
C1931 VDD.n1439 GND 0.00644f
C1932 VDD.n1440 GND 0.00644f
C1933 VDD.n1441 GND 0.008002f
C1934 VDD.n1442 GND 0.008002f
C1935 VDD.n1443 GND 0.008002f
C1936 VDD.n1444 GND 0.004991f
C1937 VDD.n1445 GND 0.008002f
C1938 VDD.n1446 GND 0.008002f
C1939 VDD.t78 GND 0.029464f
C1940 VDD.t79 GND 0.049829f
C1941 VDD.t77 GND 0.498044f
C1942 VDD.n1447 GND 0.083391f
C1943 VDD.n1448 GND 0.066666f
C1944 VDD.n1449 GND 0.013139f
C1945 VDD.n1450 GND 0.005764f
C1946 VDD.n1451 GND 0.008002f
C1947 VDD.n1452 GND 0.008002f
C1948 VDD.n1453 GND 0.008002f
C1949 VDD.n1454 GND 0.00644f
C1950 VDD.n1455 GND 0.00644f
C1951 VDD.n1456 GND 0.00644f
C1952 VDD.n1457 GND 0.008002f
C1953 VDD.n1458 GND 0.008002f
C1954 VDD.n1459 GND 0.008002f
C1955 VDD.n1460 GND 0.00644f
C1956 VDD.n1461 GND 0.006408f
C1957 VDD.n1462 GND 0.008002f
C1958 VDD.n1463 GND 0.008002f
C1959 VDD.t53 GND 0.029464f
C1960 VDD.t54 GND 0.049829f
C1961 VDD.t51 GND 0.498044f
C1962 VDD.n1464 GND 0.083391f
C1963 VDD.n1465 GND 0.066666f
C1964 VDD.n1466 GND 0.013139f
C1965 VDD.n1467 GND 0.008002f
C1966 VDD.n1468 GND 0.008002f
C1967 VDD.n1469 GND 0.008002f
C1968 VDD.n1470 GND 0.00644f
C1969 VDD.n1471 GND 0.00644f
C1970 VDD.n1472 GND 0.00644f
C1971 VDD.n1473 GND 0.008002f
C1972 VDD.n1474 GND 0.008002f
C1973 VDD.n1475 GND 0.008002f
C1974 VDD.n1476 GND 0.00644f
C1975 VDD.n1477 GND 0.005346f
C1976 VDD.n1478 GND 0.01975f
C1977 VDD.n1480 GND 1.24676f
C1978 VDD.n1481 GND 0.01975f
C1979 VDD.n1482 GND 0.002866f
C1980 VDD.n1483 GND 0.01975f
C1981 VDD.n1484 GND 0.019459f
C1982 VDD.n1485 GND 0.008002f
C1983 VDD.n1486 GND 0.00644f
C1984 VDD.n1487 GND 0.008002f
C1985 VDD.n1488 GND 0.532804f
C1986 VDD.n1489 GND 0.008002f
C1987 VDD.n1490 GND 0.00644f
C1988 VDD.n1491 GND 0.008002f
C1989 VDD.n1492 GND 0.008002f
C1990 VDD.n1493 GND 0.008002f
C1991 VDD.n1494 GND 0.00644f
C1992 VDD.n1495 GND 0.008002f
C1993 VDD.n1496 GND 0.532804f
C1994 VDD.n1497 GND 0.008002f
C1995 VDD.n1498 GND 0.00644f
C1996 VDD.n1499 GND 0.008002f
C1997 VDD.n1500 GND 0.008002f
C1998 VDD.n1501 GND 0.008002f
C1999 VDD.n1502 GND 0.00644f
C2000 VDD.n1503 GND 0.008002f
C2001 VDD.t52 GND 0.266402f
C2002 VDD.n1504 GND 0.418251f
C2003 VDD.n1505 GND 0.008002f
C2004 VDD.n1506 GND 0.00644f
C2005 VDD.n1507 GND 0.008002f
C2006 VDD.n1508 GND 0.008002f
C2007 VDD.n1509 GND 0.008002f
C2008 VDD.n1510 GND 0.00644f
C2009 VDD.n1511 GND 0.008002f
C2010 VDD.n1512 GND 0.532804f
C2011 VDD.n1513 GND 0.008002f
C2012 VDD.n1514 GND 0.00644f
C2013 VDD.n1515 GND 0.008002f
C2014 VDD.n1516 GND 0.008002f
C2015 VDD.n1517 GND 0.008002f
C2016 VDD.n1518 GND 0.00644f
C2017 VDD.n1519 GND 0.008002f
C2018 VDD.n1520 GND 0.532804f
C2019 VDD.n1521 GND 0.008002f
C2020 VDD.n1522 GND 0.00644f
C2021 VDD.n1523 GND 0.008002f
C2022 VDD.n1524 GND 0.008002f
C2023 VDD.n1525 GND 0.008002f
C2024 VDD.n1526 GND 0.00644f
C2025 VDD.n1527 GND 0.008002f
C2026 VDD.n1528 GND 0.532804f
C2027 VDD.n1529 GND 0.008002f
C2028 VDD.n1530 GND 0.00644f
C2029 VDD.n1531 GND 0.008002f
C2030 VDD.n1532 GND 0.008002f
C2031 VDD.n1533 GND 0.008002f
C2032 VDD.n1534 GND 0.00644f
C2033 VDD.n1535 GND 0.008002f
C2034 VDD.n1536 GND 0.532804f
C2035 VDD.n1537 GND 0.008002f
C2036 VDD.n1538 GND 0.00644f
C2037 VDD.n1539 GND 0.008002f
C2038 VDD.n1540 GND 0.008002f
C2039 VDD.n1541 GND 0.008002f
C2040 VDD.n1542 GND 0.00644f
C2041 VDD.n1543 GND 0.008002f
C2042 VDD.n1544 GND 0.532804f
C2043 VDD.n1545 GND 0.008002f
C2044 VDD.n1546 GND 0.00644f
C2045 VDD.n1547 GND 0.008002f
C2046 VDD.n1548 GND 0.008002f
C2047 VDD.n1549 GND 0.008002f
C2048 VDD.n1550 GND 0.00644f
C2049 VDD.n1551 GND 0.008002f
C2050 VDD.n1552 GND 0.492843f
C2051 VDD.n1553 GND 0.532804f
C2052 VDD.n1554 GND 0.008002f
C2053 VDD.n1555 GND 0.00644f
C2054 VDD.n1556 GND 0.008002f
C2055 VDD.n1557 GND 0.008002f
C2056 VDD.n1558 GND 0.008002f
C2057 VDD.n1559 GND 0.00644f
C2058 VDD.n1560 GND 0.008002f
C2059 VDD.n1561 GND 0.306362f
C2060 VDD.n1562 GND 0.008002f
C2061 VDD.n1563 GND 0.00644f
C2062 VDD.n1564 GND 0.008002f
C2063 VDD.n1565 GND 0.008002f
C2064 VDD.n1566 GND 0.008002f
C2065 VDD.n1567 GND 0.00644f
C2066 VDD.n1568 GND 0.008002f
C2067 VDD.n1569 GND 0.532804f
C2068 VDD.n1570 GND 0.008002f
C2069 VDD.n1571 GND 0.00644f
C2070 VDD.n1572 GND 0.008002f
C2071 VDD.n1573 GND 0.008002f
C2072 VDD.n1574 GND 0.008002f
C2073 VDD.n1575 GND 0.00644f
C2074 VDD.n1576 GND 0.008002f
C2075 VDD.n1577 GND 0.532804f
C2076 VDD.n1578 GND 0.008002f
C2077 VDD.n1579 GND 0.00644f
C2078 VDD.n1580 GND 0.008002f
C2079 VDD.n1581 GND 0.008002f
C2080 VDD.n1582 GND 0.008002f
C2081 VDD.n1583 GND 0.00644f
C2082 VDD.n1584 GND 0.008002f
C2083 VDD.n1585 GND 0.532804f
C2084 VDD.n1586 GND 0.008002f
C2085 VDD.n1587 GND 0.00644f
C2086 VDD.n1588 GND 0.008002f
C2087 VDD.n1589 GND 0.008002f
C2088 VDD.n1590 GND 0.008002f
C2089 VDD.n1591 GND 0.00644f
C2090 VDD.n1592 GND 0.008002f
C2091 VDD.n1593 GND 0.532804f
C2092 VDD.n1594 GND 0.008002f
C2093 VDD.n1595 GND 0.00644f
C2094 VDD.n1596 GND 0.008002f
C2095 VDD.n1597 GND 0.008002f
C2096 VDD.n1598 GND 0.008002f
C2097 VDD.n1599 GND 0.00644f
C2098 VDD.n1600 GND 0.008002f
C2099 VDD.t127 GND 0.266402f
C2100 VDD.n1601 GND 0.519484f
C2101 VDD.n1602 GND 0.008002f
C2102 VDD.n1603 GND 0.00644f
C2103 VDD.n1604 GND 0.008002f
C2104 VDD.n1605 GND 0.008002f
C2105 VDD.n1606 GND 0.008002f
C2106 VDD.n1607 GND 0.00644f
C2107 VDD.n1608 GND 0.008002f
C2108 VDD.n1609 GND 0.532804f
C2109 VDD.n1610 GND 0.008002f
C2110 VDD.n1611 GND 0.00644f
C2111 VDD.n1612 GND 0.008002f
C2112 VDD.n1613 GND 0.008002f
C2113 VDD.n1614 GND 0.008002f
C2114 VDD.n1615 GND 0.00644f
C2115 VDD.n1616 GND 0.008002f
C2116 VDD.n1617 GND 0.532804f
C2117 VDD.n1618 GND 0.008002f
C2118 VDD.n1619 GND 0.00644f
C2119 VDD.n1620 GND 0.008002f
C2120 VDD.n1621 GND 0.008002f
C2121 VDD.n1622 GND 0.004201f
C2122 VDD.n1623 GND 0.028145f
C2123 VDD.n1624 GND 0.00219f
C2124 VDD.t171 GND 0.011388f
C2125 VDD.n1625 GND 0.013332f
C2126 VDD.n1626 GND 0.003052f
C2127 VDD.n1627 GND 0.003882f
C2128 VDD.n1628 GND 0.011589f
C2129 VDD.n1629 GND 0.002319f
C2130 VDD.n1630 GND 0.00219f
C2131 VDD.n1631 GND 0.009698f
C2132 VDD.n1632 GND 0.014383f
C2133 VDD.t128 GND 0.00789f
C2134 VDD.t152 GND 0.00789f
C2135 VDD.n1633 GND 0.032694f
C2136 VDD.n1634 GND 0.23237f
C2137 VDD.n1635 GND 0.004201f
C2138 VDD.n1636 GND 0.028145f
C2139 VDD.n1637 GND 0.00219f
C2140 VDD.t161 GND 0.011388f
C2141 VDD.n1638 GND 0.013332f
C2142 VDD.n1639 GND 0.003052f
C2143 VDD.n1640 GND 0.003882f
C2144 VDD.n1641 GND 0.011589f
C2145 VDD.n1642 GND 0.002319f
C2146 VDD.n1643 GND 0.00219f
C2147 VDD.n1644 GND 0.009698f
C2148 VDD.n1645 GND 0.005795f
C2149 VDD.n1646 GND 0.090594f
C2150 VDD.n1647 GND 0.004201f
C2151 VDD.n1648 GND 0.028145f
C2152 VDD.n1649 GND 0.00219f
C2153 VDD.t156 GND 0.011388f
C2154 VDD.n1650 GND 0.013332f
C2155 VDD.n1651 GND 0.003052f
C2156 VDD.n1652 GND 0.003882f
C2157 VDD.n1653 GND 0.011589f
C2158 VDD.n1654 GND 0.002319f
C2159 VDD.n1655 GND 0.00219f
C2160 VDD.n1656 GND 0.009698f
C2161 VDD.n1657 GND 0.014383f
C2162 VDD.t159 GND 0.00789f
C2163 VDD.t172 GND 0.00789f
C2164 VDD.n1658 GND 0.032694f
C2165 VDD.n1659 GND 0.23237f
C2166 VDD.n1660 GND 0.004201f
C2167 VDD.n1661 GND 0.028145f
C2168 VDD.n1662 GND 0.00219f
C2169 VDD.t140 GND 0.011388f
C2170 VDD.n1663 GND 0.013332f
C2171 VDD.n1664 GND 0.003052f
C2172 VDD.n1665 GND 0.003882f
C2173 VDD.n1666 GND 0.011589f
C2174 VDD.n1667 GND 0.002319f
C2175 VDD.n1668 GND 0.00219f
C2176 VDD.n1669 GND 0.009698f
C2177 VDD.n1670 GND 0.005795f
C2178 VDD.n1671 GND 0.081291f
C2179 VDD.n1672 GND 0.079615f
C2180 VDD.n1673 GND 0.004201f
C2181 VDD.n1674 GND 0.028145f
C2182 VDD.n1675 GND 0.00219f
C2183 VDD.t133 GND 0.011388f
C2184 VDD.n1676 GND 0.013332f
C2185 VDD.n1677 GND 0.003052f
C2186 VDD.n1678 GND 0.003882f
C2187 VDD.n1679 GND 0.011589f
C2188 VDD.n1680 GND 0.002319f
C2189 VDD.n1681 GND 0.00219f
C2190 VDD.n1682 GND 0.009698f
C2191 VDD.n1683 GND 0.014383f
C2192 VDD.t137 GND 0.00789f
C2193 VDD.t157 GND 0.00789f
C2194 VDD.n1684 GND 0.032694f
C2195 VDD.n1685 GND 0.23237f
C2196 VDD.n1686 GND 0.004201f
C2197 VDD.n1687 GND 0.028145f
C2198 VDD.n1688 GND 0.00219f
C2199 VDD.t166 GND 0.011388f
C2200 VDD.n1689 GND 0.013332f
C2201 VDD.n1690 GND 0.003052f
C2202 VDD.n1691 GND 0.003882f
C2203 VDD.n1692 GND 0.011589f
C2204 VDD.n1693 GND 0.002319f
C2205 VDD.n1694 GND 0.00219f
C2206 VDD.n1695 GND 0.009698f
C2207 VDD.n1696 GND 0.005795f
C2208 VDD.n1697 GND 0.081291f
C2209 VDD.n1698 GND 0.0566f
C2210 VDD.n1699 GND 0.004201f
C2211 VDD.n1700 GND 0.028145f
C2212 VDD.n1701 GND 0.00219f
C2213 VDD.t155 GND 0.011388f
C2214 VDD.n1702 GND 0.013332f
C2215 VDD.n1703 GND 0.003052f
C2216 VDD.n1704 GND 0.003882f
C2217 VDD.n1705 GND 0.011589f
C2218 VDD.n1706 GND 0.002319f
C2219 VDD.n1707 GND 0.00219f
C2220 VDD.n1708 GND 0.009698f
C2221 VDD.n1709 GND 0.014383f
C2222 VDD.t134 GND 0.00789f
C2223 VDD.t164 GND 0.00789f
C2224 VDD.n1710 GND 0.032694f
C2225 VDD.n1711 GND 0.23237f
C2226 VDD.n1712 GND 0.004201f
C2227 VDD.n1713 GND 0.028145f
C2228 VDD.n1714 GND 0.00219f
C2229 VDD.t154 GND 0.011388f
C2230 VDD.n1715 GND 0.013332f
C2231 VDD.n1716 GND 0.003052f
C2232 VDD.n1717 GND 0.003882f
C2233 VDD.n1718 GND 0.011589f
C2234 VDD.n1719 GND 0.002319f
C2235 VDD.n1720 GND 0.00219f
C2236 VDD.n1721 GND 0.009698f
C2237 VDD.n1722 GND 0.005795f
C2238 VDD.n1723 GND 0.081291f
C2239 VDD.n1724 GND 0.0566f
C2240 VDD.n1725 GND 0.004201f
C2241 VDD.n1726 GND 0.028145f
C2242 VDD.n1727 GND 0.00219f
C2243 VDD.t132 GND 0.011388f
C2244 VDD.n1728 GND 0.013332f
C2245 VDD.n1729 GND 0.003052f
C2246 VDD.n1730 GND 0.003882f
C2247 VDD.n1731 GND 0.011589f
C2248 VDD.n1732 GND 0.002319f
C2249 VDD.n1733 GND 0.00219f
C2250 VDD.n1734 GND 0.009698f
C2251 VDD.n1735 GND 0.014383f
C2252 VDD.t162 GND 0.00789f
C2253 VDD.t149 GND 0.00789f
C2254 VDD.n1736 GND 0.032694f
C2255 VDD.n1737 GND 0.23237f
C2256 VDD.n1738 GND 0.004201f
C2257 VDD.n1739 GND 0.028145f
C2258 VDD.n1740 GND 0.00219f
C2259 VDD.t130 GND 0.011388f
C2260 VDD.n1741 GND 0.013332f
C2261 VDD.n1742 GND 0.003052f
C2262 VDD.n1743 GND 0.003882f
C2263 VDD.n1744 GND 0.011589f
C2264 VDD.n1745 GND 0.002319f
C2265 VDD.n1746 GND 0.00219f
C2266 VDD.n1747 GND 0.009698f
C2267 VDD.n1748 GND 0.005795f
C2268 VDD.n1749 GND 0.081291f
C2269 VDD.n1750 GND 0.152614f
C2270 VDD.n1751 GND 2.7637f
C2271 VDD.n1752 GND 0.232322f
C2272 VDD.n1753 GND 0.00615f
C2273 VDD.n1754 GND 0.00644f
C2274 VDD.n1755 GND 0.008002f
C2275 VDD.n1756 GND 0.532804f
C2276 VDD.n1757 GND 0.008002f
C2277 VDD.n1758 GND 0.00644f
C2278 VDD.n1759 GND 0.008002f
C2279 VDD.n1760 GND 0.008002f
C2280 VDD.n1761 GND 0.008002f
C2281 VDD.n1762 GND 0.00644f
C2282 VDD.n1763 GND 0.008002f
C2283 VDD.n1764 GND 0.532804f
C2284 VDD.n1765 GND 0.008002f
C2285 VDD.n1766 GND 0.00644f
C2286 VDD.n1767 GND 0.008002f
C2287 VDD.n1768 GND 0.008002f
C2288 VDD.n1769 GND 0.008002f
C2289 VDD.n1770 GND 0.00644f
C2290 VDD.n1771 GND 0.008002f
C2291 VDD.n1772 GND 0.532804f
C2292 VDD.n1773 GND 0.008002f
C2293 VDD.n1774 GND 0.00644f
C2294 VDD.n1775 GND 0.008002f
C2295 VDD.n1776 GND 0.008002f
C2296 VDD.n1777 GND 0.008002f
C2297 VDD.n1778 GND 0.00644f
C2298 VDD.n1779 GND 0.008002f
C2299 VDD.t148 GND 0.266402f
C2300 VDD.n1780 GND 0.279722f
C2301 VDD.n1781 GND 0.008002f
C2302 VDD.n1782 GND 0.00644f
C2303 VDD.n1783 GND 0.008002f
C2304 VDD.n1784 GND 0.008002f
C2305 VDD.n1785 GND 0.008002f
C2306 VDD.n1786 GND 0.00644f
C2307 VDD.n1787 GND 0.008002f
C2308 VDD.n1788 GND 0.532804f
C2309 VDD.n1789 GND 0.008002f
C2310 VDD.n1790 GND 0.00644f
C2311 VDD.n1791 GND 0.008002f
C2312 VDD.n1792 GND 0.008002f
C2313 VDD.n1793 GND 0.008002f
C2314 VDD.n1794 GND 0.00644f
C2315 VDD.n1795 GND 0.008002f
C2316 VDD.n1796 GND 0.532804f
C2317 VDD.n1797 GND 0.008002f
C2318 VDD.n1798 GND 0.00644f
C2319 VDD.n1799 GND 0.008002f
C2320 VDD.n1800 GND 0.008002f
C2321 VDD.n1801 GND 0.008002f
C2322 VDD.n1802 GND 0.00644f
C2323 VDD.n1803 GND 0.008002f
C2324 VDD.n1804 GND 0.532804f
C2325 VDD.n1805 GND 0.008002f
C2326 VDD.n1806 GND 0.00644f
C2327 VDD.n1807 GND 0.008002f
C2328 VDD.n1808 GND 0.008002f
C2329 VDD.n1809 GND 0.008002f
C2330 VDD.n1810 GND 0.00644f
C2331 VDD.n1811 GND 0.008002f
C2332 VDD.n1812 GND 0.532804f
C2333 VDD.n1813 GND 0.008002f
C2334 VDD.n1814 GND 0.00644f
C2335 VDD.n1815 GND 0.008002f
C2336 VDD.n1816 GND 0.008002f
C2337 VDD.n1817 GND 0.008002f
C2338 VDD.n1818 GND 0.00644f
C2339 VDD.n1819 GND 0.008002f
C2340 VDD.n1820 GND 0.532804f
C2341 VDD.n1821 GND 0.008002f
C2342 VDD.n1822 GND 0.00644f
C2343 VDD.n1823 GND 0.008002f
C2344 VDD.n1824 GND 0.008002f
C2345 VDD.n1825 GND 0.008002f
C2346 VDD.n1826 GND 0.00644f
C2347 VDD.n1827 GND 0.008002f
C2348 VDD.n1828 GND 0.492843f
C2349 VDD.n1829 GND 0.008002f
C2350 VDD.n1830 GND 0.00644f
C2351 VDD.n1831 GND 0.008002f
C2352 VDD.n1832 GND 0.008002f
C2353 VDD.n1833 GND 0.008002f
C2354 VDD.n1834 GND 0.00644f
C2355 VDD.n1835 GND 0.008002f
C2356 VDD.n1836 GND 0.532804f
C2357 VDD.n1837 GND 0.008002f
C2358 VDD.n1838 GND 0.00644f
C2359 VDD.n1839 GND 0.008002f
C2360 VDD.n1840 GND 0.008002f
C2361 VDD.n1841 GND 0.008002f
C2362 VDD.n1842 GND 0.00644f
C2363 VDD.n1843 GND 0.008002f
C2364 VDD.n1844 GND 0.532804f
C2365 VDD.n1845 GND 0.008002f
C2366 VDD.n1846 GND 0.00644f
C2367 VDD.n1847 GND 0.008002f
C2368 VDD.n1848 GND 0.008002f
C2369 VDD.n1849 GND 0.008002f
C2370 VDD.n1850 GND 0.00644f
C2371 VDD.n1851 GND 0.008002f
C2372 VDD.n1852 GND 0.532804f
C2373 VDD.n1853 GND 0.008002f
C2374 VDD.n1854 GND 0.00644f
C2375 VDD.n1855 GND 0.008002f
C2376 VDD.n1856 GND 0.008002f
C2377 VDD.n1857 GND 0.008002f
C2378 VDD.n1858 GND 0.00644f
C2379 VDD.n1859 GND 0.008002f
C2380 VDD.n1860 GND 0.532804f
C2381 VDD.n1861 GND 0.008002f
C2382 VDD.n1862 GND 0.00644f
C2383 VDD.n1863 GND 0.008002f
C2384 VDD.n1864 GND 0.008002f
C2385 VDD.n1865 GND 0.008002f
C2386 VDD.n1866 GND 0.00644f
C2387 VDD.n1867 GND 0.008002f
C2388 VDD.n1868 GND 0.532804f
C2389 VDD.n1869 GND 0.008002f
C2390 VDD.n1870 GND 0.00644f
C2391 VDD.n1871 GND 0.008002f
C2392 VDD.n1872 GND 0.008002f
C2393 VDD.n1873 GND 0.008002f
C2394 VDD.n1874 GND 0.00644f
C2395 VDD.n1875 GND 0.008002f
C2396 VDD.t42 GND 0.266402f
C2397 VDD.n1876 GND 0.380955f
C2398 VDD.n1877 GND 0.008002f
C2399 VDD.n1878 GND 0.00644f
C2400 VDD.n1879 GND 0.008002f
C2401 VDD.n1880 GND 0.008002f
C2402 VDD.n1881 GND 0.008002f
C2403 VDD.n1882 GND 0.00644f
C2404 VDD.n1883 GND 0.008002f
C2405 VDD.n1884 GND 0.532804f
C2406 VDD.n1885 GND 0.008002f
C2407 VDD.n1886 GND 0.00644f
C2408 VDD.n1887 GND 0.008002f
C2409 VDD.n1888 GND 0.008002f
C2410 VDD.n1889 GND 0.008002f
C2411 VDD.n1890 GND 0.00644f
C2412 VDD.n1891 GND 0.008002f
C2413 VDD.n1892 GND 0.532804f
C2414 VDD.n1893 GND 0.008002f
C2415 VDD.n1894 GND 0.00644f
C2416 VDD.n1895 GND 0.008002f
C2417 VDD.n1896 GND 0.008002f
C2418 VDD.n1897 GND 0.008002f
C2419 VDD.n1898 GND 0.00644f
C2420 VDD.n1900 GND 0.008002f
C2421 VDD.n1901 GND 0.00644f
C2422 VDD.n1902 GND 0.004641f
C2423 VDD.n1903 GND 0.004347f
C2424 VDD.n1905 GND 0.008002f
C2425 VDD.n1906 GND 0.00644f
C2426 VDD.n1907 GND 0.008002f
C2427 VDD.n1908 GND 0.00644f
C2428 VDD.n1910 GND 0.008002f
C2429 VDD.n1911 GND 0.00644f
C2430 VDD.n1912 GND 0.008002f
C2431 VDD.n1913 GND 0.008002f
C2432 VDD.n1914 GND 0.008002f
C2433 VDD.n1915 GND 0.008002f
C2434 VDD.n1916 GND 0.008002f
C2435 VDD.t44 GND 0.029464f
C2436 VDD.t43 GND 0.049829f
C2437 VDD.t41 GND 0.498044f
C2438 VDD.n1917 GND 0.083391f
C2439 VDD.n1918 GND 0.066666f
C2440 VDD.n1919 GND 0.013139f
C2441 VDD.n1921 GND 0.008002f
C2442 VDD.n1922 GND 0.008002f
C2443 VDD.n1923 GND 0.008002f
C2444 VDD.n1924 GND 0.008002f
C2445 VDD.n1925 GND 0.008002f
C2446 VDD.n1926 GND 0.00644f
C2447 VDD.n1928 GND 0.008002f
C2448 VDD.n1929 GND 0.008002f
C2449 VDD.n1930 GND 0.008002f
C2450 VDD.n1931 GND 0.008002f
C2451 VDD.n1932 GND 0.008002f
C2452 VDD.n1933 GND 0.00644f
C2453 VDD.n1935 GND 0.008002f
C2454 VDD.n1936 GND 0.008002f
C2455 VDD.n1937 GND 0.008002f
C2456 VDD.n1938 GND 0.008002f
C2457 VDD.n1939 GND 0.008002f
C2458 VDD.n1940 GND 0.00644f
C2459 VDD.n1942 GND 0.008002f
C2460 VDD.n1943 GND 0.008002f
C2461 VDD.n1944 GND 0.008002f
C2462 VDD.n1945 GND 0.008002f
C2463 VDD.n1946 GND 0.008002f
C2464 VDD.n1947 GND 0.00644f
C2465 VDD.n1949 GND 0.008002f
C2466 VDD.n1950 GND 0.008002f
C2467 VDD.n1951 GND 0.008002f
C2468 VDD.n1952 GND 0.008002f
C2469 VDD.n1953 GND 0.005378f
C2470 VDD.t67 GND 0.029464f
C2471 VDD.t66 GND 0.049829f
C2472 VDD.t65 GND 0.498044f
C2473 VDD.n1954 GND 0.083391f
C2474 VDD.n1955 GND 0.066666f
C2475 VDD.n1957 GND 0.008002f
C2476 VDD.n1958 GND 0.00644f
C2477 VDD.n1959 GND 0.008002f
C2478 VDD.n1961 GND 0.00644f
C2479 VDD.n1963 GND 0.008002f
C2480 VDD.n1964 GND 0.00644f
C2481 VDD.n1965 GND 0.008002f
C2482 VDD.n1967 GND 0.008002f
C2483 VDD.n1968 GND 0.00644f
C2484 VDD.n1969 GND 0.008002f
C2485 VDD.n1971 GND 0.008002f
C2486 VDD.n1972 GND 0.008002f
C2487 VDD.n1973 GND 0.00644f
C2488 VDD.n1974 GND 0.008002f
C2489 VDD.n1975 GND 0.008002f
C2490 VDD.n1976 GND 0.008002f
C2491 VDD.n1977 GND 0.013139f
C2492 VDD.n1978 GND 0.005378f
C2493 VDD.n1979 GND 0.00644f
C2494 VDD.n1980 GND 0.008002f
C2495 VDD.n1982 GND 0.008002f
C2496 VDD.n1983 GND 0.008002f
C2497 VDD.n1984 GND 0.00644f
C2498 VDD.n1985 GND 0.00644f
C2499 VDD.n1986 GND 0.00644f
C2500 VDD.n1987 GND 0.008002f
C2501 VDD.n1989 GND 0.008002f
C2502 VDD.n1990 GND 0.008002f
C2503 VDD.n1991 GND 0.00644f
C2504 VDD.n1992 GND 0.003574f
C2505 VDD.t121 GND 0.029464f
C2506 VDD.t120 GND 0.049829f
C2507 VDD.t119 GND 0.498044f
C2508 VDD.n1993 GND 0.083391f
C2509 VDD.n1994 GND 0.066666f
C2510 VDD.n1995 GND 0.009918f
C2511 VDD.n1996 GND 0.003961f
C2512 VDD.n1997 GND 0.008002f
C2513 VDD.n1999 GND 0.008002f
C2514 VDD.n2000 GND 0.008002f
C2515 VDD.n2001 GND 0.00644f
C2516 VDD.n2002 GND 0.00644f
C2517 VDD.n2003 GND 0.00644f
C2518 VDD.n2004 GND 0.008002f
C2519 VDD.n2006 GND 0.008002f
C2520 VDD.n2007 GND 0.008002f
C2521 VDD.n2008 GND 0.00644f
C2522 VDD.n2009 GND 0.00644f
C2523 VDD.n2010 GND 0.004991f
C2524 VDD.n2011 GND 0.008002f
C2525 VDD.n2013 GND 0.008002f
C2526 VDD.n2014 GND 0.008002f
C2527 VDD.n2015 GND 0.005764f
C2528 VDD.n2016 GND 0.00644f
C2529 VDD.n2017 GND 0.00644f
C2530 VDD.n2018 GND 0.008002f
C2531 VDD.n2020 GND 0.008002f
C2532 VDD.n2021 GND 0.008002f
C2533 VDD.n2023 GND 0.008002f
C2534 VDD.n2024 GND 0.00644f
C2535 VDD.n2025 GND 0.008002f
C2536 VDD.n2026 GND 0.008002f
C2537 VDD.n2027 GND 0.008002f
C2538 VDD.n2028 GND 0.006408f
C2539 VDD.t99 GND 0.029464f
C2540 VDD.t98 GND 0.049829f
C2541 VDD.t97 GND 0.498044f
C2542 VDD.n2029 GND 0.083391f
C2543 VDD.n2030 GND 0.066666f
C2544 VDD.n2031 GND 0.013139f
C2545 VDD.n2032 GND 0.008002f
C2546 VDD.n2034 GND 0.008002f
C2547 VDD.n2035 GND 0.008002f
C2548 VDD.n2036 GND 0.00644f
C2549 VDD.n2038 GND 0.005441f
C2550 VDD.n2039 GND 0.005441f
C2551 VDD.n2040 GND 0.005441f
C2552 VDD.n2041 GND 0.005441f
C2553 VDD.n2042 GND 0.005441f
C2554 VDD.n2043 GND 0.005441f
C2555 VDD.n2044 GND 0.005441f
C2556 VDD.n2045 GND 0.005441f
C2557 VDD.n2046 GND 0.005441f
C2558 VDD.n2047 GND 0.005441f
C2559 VDD.n2048 GND 0.005441f
C2560 VDD.n2049 GND 0.005441f
C2561 VDD.n2050 GND 0.005441f
C2562 VDD.n2051 GND 0.005441f
C2563 VDD.n2052 GND 0.004081f
C2564 VDD.t82 GND 0.111051f
C2565 VDD.t83 GND 0.129192f
C2566 VDD.t80 GND 0.629305f
C2567 VDD.n2053 GND 0.086428f
C2568 VDD.n2054 GND 0.052244f
C2569 VDD.n2055 GND 0.005441f
C2570 VDD.n2056 GND 0.005441f
C2571 VDD.n2057 GND 0.005441f
C2572 VDD.n2058 GND 0.005441f
C2573 VDD.n2059 GND 0.005441f
C2574 VDD.n2060 GND 0.005441f
C2575 VDD.n2061 GND 0.005441f
C2576 VDD.n2062 GND 0.005441f
C2577 VDD.n2063 GND 0.005441f
C2578 VDD.n2064 GND 0.005441f
C2579 VDD.n2065 GND 0.005441f
C2580 VDD.n2066 GND 0.005441f
C2581 VDD.n2067 GND 0.005441f
C2582 VDD.n2068 GND 0.005441f
C2583 VDD.n2069 GND 0.005441f
C2584 VDD.n2070 GND 0.005441f
C2585 VDD.n2071 GND 0.005441f
C2586 VDD.n2072 GND 0.005441f
C2587 VDD.n2073 GND 0.005441f
C2588 VDD.n2074 GND 0.005441f
C2589 VDD.n2075 GND 0.005441f
C2590 VDD.n2076 GND 0.005441f
C2591 VDD.n2077 GND 0.005441f
C2592 VDD.n2078 GND 0.005441f
C2593 VDD.n2079 GND 0.005441f
C2594 VDD.n2080 GND 0.005441f
C2595 VDD.n2081 GND 0.005441f
C2596 VDD.n2082 GND 0.005441f
C2597 VDD.n2083 GND 0.005441f
C2598 VDD.n2084 GND 0.005441f
C2599 VDD.n2085 GND 0.005441f
C2600 VDD.n2086 GND 0.005441f
C2601 VDD.n2087 GND 0.005441f
C2602 VDD.n2088 GND 0.005441f
C2603 VDD.n2089 GND 0.005441f
C2604 VDD.n2090 GND 0.005441f
C2605 VDD.n2091 GND 0.005441f
C2606 VDD.n2092 GND 0.005441f
C2607 VDD.n2093 GND 0.005441f
C2608 VDD.n2094 GND 0.005441f
C2609 VDD.n2095 GND 0.005441f
C2610 VDD.n2096 GND 0.005441f
C2611 VDD.n2097 GND 0.005441f
C2612 VDD.n2098 GND 0.005441f
C2613 VDD.n2099 GND 0.005441f
C2614 VDD.n2100 GND 0.005441f
C2615 VDD.n2101 GND 0.005441f
C2616 VDD.n2102 GND 0.005441f
C2617 VDD.n2103 GND 0.005441f
C2618 VDD.n2104 GND 0.005441f
C2619 VDD.n2105 GND 0.005441f
C2620 VDD.n2106 GND 0.005441f
C2621 VDD.n2107 GND 0.005441f
C2622 VDD.n2108 GND 0.005441f
C2623 VDD.n2109 GND 0.005441f
C2624 VDD.n2110 GND 0.005441f
C2625 VDD.n2111 GND 0.005441f
C2626 VDD.n2112 GND 0.005441f
C2627 VDD.n2113 GND 0.005441f
C2628 VDD.n2114 GND 0.005441f
C2629 VDD.n2115 GND 0.005441f
C2630 VDD.n2116 GND 0.005441f
C2631 VDD.n2117 GND 0.005441f
C2632 VDD.n2118 GND 0.005441f
C2633 VDD.n2119 GND 0.005441f
C2634 VDD.n2120 GND 0.005441f
C2635 VDD.n2121 GND 0.005441f
C2636 VDD.n2122 GND 0.005441f
C2637 VDD.n2123 GND 0.005441f
C2638 VDD.n2124 GND 0.005441f
C2639 VDD.n2125 GND 0.005441f
C2640 VDD.n2126 GND 0.005441f
C2641 VDD.n2127 GND 0.005441f
C2642 VDD.n2128 GND 0.005441f
C2643 VDD.n2129 GND 0.005441f
C2644 VDD.n2130 GND 0.005441f
C2645 VDD.n2131 GND 0.005441f
C2646 VDD.n2132 GND 0.005441f
C2647 VDD.n2133 GND 0.005441f
C2648 VDD.n2134 GND 0.005441f
C2649 VDD.n2135 GND 0.005441f
C2650 VDD.n2136 GND 0.005441f
C2651 VDD.n2137 GND 0.005441f
C2652 VDD.n2138 GND 0.005441f
C2653 VDD.n2139 GND 0.005441f
C2654 VDD.n2140 GND 0.005441f
C2655 VDD.n2141 GND 0.005441f
C2656 VDD.n2142 GND 0.005441f
C2657 VDD.n2143 GND 0.005441f
C2658 VDD.n2144 GND 0.005441f
C2659 VDD.n2145 GND 0.005441f
C2660 VDD.n2146 GND 0.005441f
C2661 VDD.n2147 GND 0.005441f
C2662 VDD.n2148 GND 0.005441f
C2663 VDD.n2149 GND 0.005441f
C2664 VDD.n2150 GND 0.005441f
C2665 VDD.n2151 GND 0.005441f
C2666 VDD.n2152 GND 0.005441f
C2667 VDD.n2153 GND 0.005441f
C2668 VDD.n2154 GND 0.005441f
C2669 VDD.n2155 GND 0.005441f
C2670 VDD.n2156 GND 0.005441f
C2671 VDD.n2157 GND 0.005441f
C2672 VDD.n2158 GND 0.005441f
C2673 VDD.n2159 GND 0.005441f
C2674 VDD.n2160 GND 0.005441f
C2675 VDD.n2161 GND 0.005441f
C2676 VDD.n2162 GND 0.005441f
C2677 VDD.n2163 GND 0.005441f
C2678 VDD.n2164 GND 0.005441f
C2679 VDD.n2165 GND 0.005441f
C2680 VDD.n2166 GND 0.005441f
C2681 VDD.n2167 GND 0.005441f
C2682 VDD.n2168 GND 0.005441f
C2683 VDD.n2169 GND 0.005441f
C2684 VDD.n2170 GND 0.005441f
C2685 VDD.n2171 GND 0.005441f
C2686 VDD.n2172 GND 0.005441f
C2687 VDD.n2173 GND 0.011992f
C2688 VDD.n2174 GND 0.013054f
C2689 VDD.n2175 GND 0.005441f
C2690 VDD.n2176 GND 0.004841f
C2691 VDD.n2177 GND 0.007776f
C2692 VDD.n2178 GND 0.003321f
C2693 VDD.n2179 GND 0.005441f
C2694 VDD.n2180 GND 0.005441f
C2695 VDD.n2181 GND 0.005441f
C2696 VDD.n2182 GND 0.005441f
C2697 VDD.n2183 GND 0.005441f
C2698 VDD.n2184 GND 0.005441f
C2699 VDD.n2185 GND 0.005441f
C2700 VDD.n2186 GND 0.005441f
C2701 VDD.n2187 GND 0.005441f
C2702 VDD.n2188 GND 0.005441f
C2703 VDD.n2189 GND 0.005441f
C2704 VDD.n2190 GND 0.005441f
C2705 VDD.n2191 GND 0.005441f
C2706 VDD.n2192 GND 0.005441f
C2707 VDD.n2193 GND 0.005441f
C2708 VDD.n2194 GND 0.005441f
C2709 VDD.n2195 GND 0.005441f
C2710 VDD.n2196 GND 0.004081f
C2711 VDD.n2197 GND 0.030651f
C2712 VDD.n2198 GND 0.007362f
C2713 VDD.n2199 GND 0.802014f
C2714 VDD.n2201 GND 0.00644f
C2715 VDD.n2202 GND 0.008002f
C2716 VDD.n2204 GND 0.008002f
C2717 VDD.n2205 GND 0.008002f
C2718 VDD.n2206 GND 0.00644f
C2719 VDD.n2207 GND 0.005346f
C2720 VDD.n2208 GND 0.01975f
C2721 VDD.n2209 GND 0.019459f
C2722 VDD.n2210 GND 0.005346f
C2723 VDD.n2211 GND 0.019459f
C2724 VDD.n2212 GND 0.772565f
C2725 VDD.n2213 GND 0.019459f
C2726 VDD.n2214 GND 0.005346f
C2727 VDD.n2215 GND 0.019459f
C2728 VDD.n2216 GND 0.01975f
C2729 VDD.n2217 GND 0.002866f
C2730 VDD.t111 GND 0.029464f
C2731 VDD.t110 GND 0.049829f
C2732 VDD.t109 GND 0.498044f
C2733 VDD.n2218 GND 0.083391f
C2734 VDD.n2219 GND 0.066666f
C2735 VDD.n2220 GND 0.009918f
C2736 VDD.n2221 GND 0.003574f
C2737 VDD.n2222 GND 0.00644f
C2738 VDD.n2223 GND 0.007362f
C2739 VDD.n2224 GND 0.802014f
C2740 VDD.n2225 GND 0.030651f
C2741 VDD.n2226 GND 0.005441f
C2742 VDD.n2227 GND 0.005441f
C2743 VDD.n2228 GND 0.005441f
C2744 VDD.n2229 GND 0.005441f
C2745 VDD.n2230 GND 0.005441f
C2746 VDD.n2231 GND 0.005441f
C2747 VDD.n2232 GND 0.005441f
C2748 VDD.n2233 GND 0.005441f
C2749 VDD.n2234 GND 0.005441f
C2750 VDD.n2235 GND 0.005441f
C2751 VDD.n2236 GND 0.005441f
C2752 VDD.n2237 GND 0.005441f
C2753 VDD.n2238 GND 0.005441f
C2754 VDD.n2239 GND 0.005441f
C2755 VDD.n2240 GND 0.005441f
C2756 VDD.n2241 GND 0.005441f
C2757 VDD.n2242 GND 0.005441f
C2758 VDD.n2243 GND 0.005441f
C2759 VDD.n2244 GND 0.004081f
C2760 VDD.n2245 GND 0.005441f
C2761 VDD.n2246 GND 0.005441f
C2762 VDD.n2247 GND 0.004081f
C2763 VDD.n2248 GND 0.005441f
C2764 VDD.n2249 GND 0.005441f
C2765 VDD.n2250 GND 0.005441f
C2766 VDD.n2251 GND 0.005441f
C2767 VDD.n2252 GND 0.005441f
C2768 VDD.n2253 GND 0.005441f
C2769 VDD.n2254 GND 0.005441f
C2770 VDD.n2255 GND 0.005441f
C2771 VDD.n2256 GND 0.005441f
C2772 VDD.n2257 GND 0.005441f
C2773 VDD.n2258 GND 0.005441f
C2774 VDD.n2259 GND 0.005441f
C2775 VDD.n2260 GND 0.005441f
C2776 VDD.n2261 GND 0.005441f
C2777 VDD.n2262 GND 0.005441f
C2778 VDD.n2263 GND 0.003321f
C2779 VDD.n2264 GND 0.007776f
C2780 VDD.n2265 GND 0.004841f
C2781 VDD.n2266 GND 0.005441f
C2782 VDD.n2267 GND 0.005441f
C2783 VDD.n2268 GND 0.005441f
C2784 VDD.n2269 GND 0.005441f
C2785 VDD.n2270 GND 0.005441f
C2786 VDD.n2271 GND 0.005441f
C2787 VDD.n2272 GND 0.005441f
C2788 VDD.n2273 GND 0.005441f
C2789 VDD.n2274 GND 0.005441f
C2790 VDD.n2275 GND 0.005441f
C2791 VDD.n2276 GND 0.005441f
C2792 VDD.n2277 GND 0.005441f
C2793 VDD.n2278 GND 0.005441f
C2794 VDD.n2279 GND 0.005441f
C2795 VDD.n2280 GND 0.005441f
C2796 VDD.n2281 GND 0.005441f
C2797 VDD.n2282 GND 0.005441f
C2798 VDD.n2283 GND 0.005441f
C2799 VDD.n2284 GND 0.005441f
C2800 VDD.n2285 GND 0.005441f
C2801 VDD.n2286 GND 0.005441f
C2802 VDD.n2287 GND 0.005441f
C2803 VDD.n2288 GND 0.005441f
C2804 VDD.n2289 GND 0.005441f
C2805 VDD.n2290 GND 0.005441f
C2806 VDD.n2291 GND 0.005441f
C2807 VDD.n2292 GND 0.005441f
C2808 VDD.n2293 GND 0.005441f
C2809 VDD.n2294 GND 0.005441f
C2810 VDD.n2295 GND 0.005441f
C2811 VDD.n2296 GND 0.005441f
C2812 VDD.n2297 GND 0.005441f
C2813 VDD.n2298 GND 0.005441f
C2814 VDD.n2299 GND 0.005441f
C2815 VDD.n2300 GND 0.005441f
C2816 VDD.n2301 GND 0.005441f
C2817 VDD.n2302 GND 0.005441f
C2818 VDD.n2303 GND 0.005441f
C2819 VDD.n2304 GND 0.005441f
C2820 VDD.n2305 GND 0.005441f
C2821 VDD.n2306 GND 0.005441f
C2822 VDD.n2307 GND 0.005441f
C2823 VDD.n2308 GND 0.005441f
C2824 VDD.n2309 GND 0.005441f
C2825 VDD.n2310 GND 0.005441f
C2826 VDD.n2311 GND 0.005441f
C2827 VDD.n2312 GND 0.005441f
C2828 VDD.n2313 GND 0.005441f
C2829 VDD.n2314 GND 0.005441f
C2830 VDD.n2315 GND 0.005441f
C2831 VDD.n2316 GND 0.005441f
C2832 VDD.n2317 GND 0.005441f
C2833 VDD.n2318 GND 0.005441f
C2834 VDD.n2319 GND 0.005441f
C2835 VDD.n2320 GND 0.005441f
C2836 VDD.n2321 GND 0.005441f
C2837 VDD.n2322 GND 0.005441f
C2838 VDD.n2323 GND 0.005441f
C2839 VDD.n2324 GND 0.005441f
C2840 VDD.n2325 GND 0.005441f
C2841 VDD.n2326 GND 0.005441f
C2842 VDD.n2327 GND 0.005441f
C2843 VDD.n2328 GND 0.005441f
C2844 VDD.n2329 GND 0.005441f
C2845 VDD.n2330 GND 0.005441f
C2846 VDD.n2331 GND 0.005441f
C2847 VDD.n2332 GND 0.005441f
C2848 VDD.n2333 GND 0.005441f
C2849 VDD.n2334 GND 0.005441f
C2850 VDD.n2335 GND 0.005441f
C2851 VDD.n2336 GND 0.005441f
C2852 VDD.n2337 GND 0.005441f
C2853 VDD.n2338 GND 0.005441f
C2854 VDD.n2339 GND 0.005441f
C2855 VDD.n2340 GND 0.005441f
C2856 VDD.n2341 GND 0.005441f
C2857 VDD.n2342 GND 0.005441f
C2858 VDD.n2343 GND 0.005441f
C2859 VDD.n2344 GND 0.005441f
C2860 VDD.n2345 GND 0.005441f
C2861 VDD.n2346 GND 0.005441f
C2862 VDD.n2347 GND 0.005441f
C2863 VDD.n2348 GND 0.005441f
C2864 VDD.n2349 GND 0.005441f
C2865 VDD.n2350 GND 0.005441f
C2866 VDD.n2351 GND 0.005441f
C2867 VDD.n2352 GND 0.005441f
C2868 VDD.n2353 GND 0.005441f
C2869 VDD.n2354 GND 0.005441f
C2870 VDD.n2355 GND 0.005441f
C2871 VDD.n2356 GND 0.005441f
C2872 VDD.n2357 GND 0.005441f
C2873 VDD.n2358 GND 0.005441f
C2874 VDD.n2359 GND 0.005441f
C2875 VDD.n2360 GND 0.005441f
C2876 VDD.n2361 GND 0.005441f
C2877 VDD.n2362 GND 0.005441f
C2878 VDD.n2363 GND 0.005441f
C2879 VDD.n2364 GND 0.005441f
C2880 VDD.n2365 GND 0.005441f
C2881 VDD.n2366 GND 0.005441f
C2882 VDD.n2367 GND 0.005441f
C2883 VDD.n2368 GND 0.005441f
C2884 VDD.n2369 GND 0.005441f
C2885 VDD.n2370 GND 0.005441f
C2886 VDD.n2371 GND 0.005441f
C2887 VDD.n2372 GND 0.005441f
C2888 VDD.n2373 GND 0.005441f
C2889 VDD.n2374 GND 0.005441f
C2890 VDD.n2375 GND 0.005441f
C2891 VDD.n2376 GND 0.005441f
C2892 VDD.n2377 GND 0.005441f
C2893 VDD.n2378 GND 0.005441f
C2894 VDD.n2379 GND 0.005441f
C2895 VDD.n2380 GND 0.005441f
C2896 VDD.n2381 GND 0.005441f
C2897 VDD.n2382 GND 0.005441f
C2898 VDD.n2383 GND 0.005441f
C2899 VDD.n2384 GND 0.005441f
C2900 VDD.n2385 GND 0.005441f
C2901 VDD.n2386 GND 0.005441f
C2902 VDD.n2387 GND 0.011992f
C2903 VDD.n2388 GND 0.013054f
C2904 VDD.n2389 GND 0.013054f
C2905 VDD.n2390 GND 2.51483f
C2906 VDD.n2392 GND 0.005441f
C2907 VDD.n2393 GND 0.005441f
C2908 VDD.n2394 GND 0.013054f
C2909 VDD.n2395 GND 0.011992f
C2910 VDD.n2396 GND 0.011992f
C2911 VDD.n2397 GND 0.450219f
C2912 VDD.n2398 GND 0.011992f
C2913 VDD.n2399 GND 0.011992f
C2914 VDD.n2400 GND 0.005441f
C2915 VDD.n2401 GND 0.005441f
C2916 VDD.n2402 GND 0.005441f
C2917 VDD.n2403 GND 0.362306f
C2918 VDD.n2404 GND 0.005441f
C2919 VDD.n2405 GND 0.005441f
C2920 VDD.n2406 GND 0.005441f
C2921 VDD.n2407 GND 0.005441f
C2922 VDD.n2408 GND 0.005441f
C2923 VDD.n2409 GND 0.362306f
C2924 VDD.n2410 GND 0.005441f
C2925 VDD.n2411 GND 0.005441f
C2926 VDD.n2412 GND 0.005441f
C2927 VDD.n2413 GND 0.005441f
C2928 VDD.n2414 GND 0.005441f
C2929 VDD.n2415 GND 0.229106f
C2930 VDD.n2416 GND 0.005441f
C2931 VDD.n2417 GND 0.005441f
C2932 VDD.n2418 GND 0.005441f
C2933 VDD.n2419 GND 0.005441f
C2934 VDD.n2420 GND 0.005441f
C2935 VDD.n2421 GND 0.362306f
C2936 VDD.n2422 GND 0.005441f
C2937 VDD.n2423 GND 0.005441f
C2938 VDD.n2424 GND 0.005441f
C2939 VDD.n2425 GND 0.005441f
C2940 VDD.n2426 GND 0.005441f
C2941 VDD.n2427 GND 0.327674f
C2942 VDD.n2428 GND 0.005441f
C2943 VDD.n2429 GND 0.005441f
C2944 VDD.n2430 GND 0.005441f
C2945 VDD.n2431 GND 0.005441f
C2946 VDD.n2432 GND 0.005441f
C2947 VDD.n2433 GND 0.362306f
C2948 VDD.n2434 GND 0.005441f
C2949 VDD.n2435 GND 0.005441f
C2950 VDD.n2436 GND 0.005441f
C2951 VDD.n2437 GND 0.005441f
C2952 VDD.n2438 GND 0.005441f
C2953 VDD.n2439 GND 0.362306f
C2954 VDD.n2440 GND 0.005441f
C2955 VDD.n2441 GND 0.005441f
C2956 VDD.n2442 GND 0.005441f
C2957 VDD.n2443 GND 0.005441f
C2958 VDD.n2444 GND 0.005441f
C2959 VDD.n2445 GND 0.362306f
C2960 VDD.n2446 GND 0.005441f
C2961 VDD.n2447 GND 0.005441f
C2962 VDD.n2448 GND 0.005441f
C2963 VDD.n2449 GND 0.005441f
C2964 VDD.n2450 GND 0.005441f
C2965 VDD.n2451 GND 0.362306f
C2966 VDD.n2452 GND 0.005441f
C2967 VDD.n2453 GND 0.005441f
C2968 VDD.n2454 GND 0.005441f
C2969 VDD.n2455 GND 0.005441f
C2970 VDD.n2456 GND 0.005441f
C2971 VDD.n2457 GND 0.050616f
C2972 VDD.n2458 GND 0.005441f
C2973 VDD.n2459 GND 0.005441f
C2974 VDD.n2460 GND 0.005441f
C2975 VDD.n2461 GND 0.005441f
C2976 VDD.n2462 GND 0.005441f
C2977 VDD.n2463 GND 0.362306f
C2978 VDD.n2464 GND 0.005441f
C2979 VDD.n2465 GND 0.005441f
C2980 VDD.n2466 GND 0.005441f
C2981 VDD.n2467 GND 0.005441f
C2982 VDD.n2468 GND 0.005441f
C2983 VDD.n2469 GND 0.362306f
C2984 VDD.n2470 GND 0.005441f
C2985 VDD.n2471 GND 0.005441f
C2986 VDD.n2472 GND 0.005441f
C2987 VDD.n2473 GND 0.005441f
C2988 VDD.n2474 GND 0.005441f
C2989 VDD.n2475 GND 0.362306f
C2990 VDD.n2476 GND 0.005441f
C2991 VDD.n2477 GND 0.005441f
C2992 VDD.n2478 GND 0.005441f
C2993 VDD.n2479 GND 0.005441f
C2994 VDD.n2480 GND 0.005441f
C2995 VDD.n2481 GND 0.362306f
C2996 VDD.n2482 GND 0.005441f
C2997 VDD.n2483 GND 0.005441f
C2998 VDD.n2484 GND 0.005441f
C2999 VDD.n2485 GND 0.005441f
C3000 VDD.n2486 GND 0.005441f
C3001 VDD.n2487 GND 0.279722f
C3002 VDD.n2488 GND 0.005441f
C3003 VDD.n2489 GND 0.005441f
C3004 VDD.n2490 GND 0.005441f
C3005 VDD.n2491 GND 0.005441f
C3006 VDD.n2492 GND 0.005441f
C3007 VDD.n2493 GND 0.362306f
C3008 VDD.n2494 GND 0.005441f
C3009 VDD.n2495 GND 0.005441f
C3010 VDD.n2496 GND 0.005441f
C3011 VDD.n2497 GND 0.005441f
C3012 VDD.n2498 GND 0.005441f
C3013 VDD.n2499 GND 0.362306f
C3014 VDD.n2500 GND 0.005441f
C3015 VDD.n2501 GND 0.005441f
C3016 VDD.n2502 GND 0.005441f
C3017 VDD.n2503 GND 0.005441f
C3018 VDD.n2504 GND 0.005441f
C3019 VDD.n2505 GND 0.362306f
C3020 VDD.n2506 GND 0.005441f
C3021 VDD.n2507 GND 0.005441f
C3022 VDD.n2508 GND 0.005441f
C3023 VDD.n2509 GND 0.005441f
C3024 VDD.n2510 GND 0.005441f
C3025 VDD.n2511 GND 0.362306f
C3026 VDD.n2512 GND 0.005441f
C3027 VDD.n2513 GND 0.005441f
C3028 VDD.n2514 GND 0.005441f
C3029 VDD.n2515 GND 0.005441f
C3030 VDD.n2516 GND 0.005441f
C3031 VDD.n2517 GND 0.362306f
C3032 VDD.n2518 GND 0.005441f
C3033 VDD.n2519 GND 0.005441f
C3034 VDD.n2520 GND 0.005441f
C3035 VDD.n2521 GND 0.005441f
C3036 VDD.n2522 GND 0.005441f
C3037 VDD.n2523 GND 0.27173f
C3038 VDD.n2524 GND 0.005441f
C3039 VDD.n2525 GND 0.005441f
C3040 VDD.n2526 GND 0.005441f
C3041 VDD.n2527 GND 0.005441f
C3042 VDD.n2528 GND 0.005441f
C3043 VDD.n2529 GND 0.362306f
C3044 VDD.n2530 GND 0.005441f
C3045 VDD.n2531 GND 0.005441f
C3046 VDD.n2532 GND 0.005441f
C3047 VDD.n2533 GND 0.005441f
C3048 VDD.n2534 GND 0.005441f
C3049 VDD.n2535 GND 0.31169f
C3050 VDD.n2536 GND 0.005441f
C3051 VDD.n2537 GND 0.005441f
C3052 VDD.n2538 GND 0.005441f
C3053 VDD.n2539 GND 0.005441f
C3054 VDD.n2540 GND 0.005441f
C3055 VDD.n2541 GND 0.362306f
C3056 VDD.n2542 GND 0.005441f
C3057 VDD.n2543 GND 0.005441f
C3058 VDD.n2544 GND 0.005441f
C3059 VDD.n2545 GND 0.005441f
C3060 VDD.n2546 GND 0.005441f
C3061 VDD.n2547 GND 0.362306f
C3062 VDD.n2548 GND 0.005441f
C3063 VDD.n2549 GND 0.005441f
C3064 VDD.n2550 GND 0.005441f
C3065 VDD.n2551 GND 0.005441f
C3066 VDD.n2552 GND 0.005441f
C3067 VDD.n2553 GND 0.213121f
C3068 VDD.n2554 GND 0.005441f
C3069 VDD.n2555 GND 0.005441f
C3070 VDD.n2556 GND 0.005441f
C3071 VDD.n2557 GND 0.005441f
C3072 VDD.n2558 GND 0.005441f
C3073 VDD.n2559 GND 0.362306f
C3074 VDD.n2560 GND 0.005441f
C3075 VDD.n2561 GND 0.005441f
C3076 VDD.n2562 GND 0.005441f
C3077 VDD.n2563 GND 0.005441f
C3078 VDD.n2564 GND 0.005441f
C3079 VDD.n2565 GND 0.362306f
C3080 VDD.n2566 GND 0.005441f
C3081 VDD.n2567 GND 0.005441f
C3082 VDD.n2568 GND 0.005441f
C3083 VDD.n2569 GND 0.005441f
C3084 VDD.n2570 GND 0.005441f
C3085 VDD.n2571 GND 0.290378f
C3086 VDD.n2572 GND 0.005441f
C3087 VDD.n2573 GND 0.005441f
C3088 VDD.n2574 GND 0.005441f
C3089 VDD.n2575 GND 0.005441f
C3090 VDD.n2576 GND 0.005441f
C3091 VDD.n2577 GND 0.362306f
C3092 VDD.n2578 GND 0.005441f
C3093 VDD.n2579 GND 0.005441f
C3094 VDD.n2580 GND 0.005441f
C3095 VDD.n2581 GND 0.005441f
C3096 VDD.n2582 GND 0.005441f
C3097 VDD.n2583 GND 0.335666f
C3098 VDD.n2584 GND 0.005441f
C3099 VDD.n2585 GND 0.005441f
C3100 VDD.n2586 GND 0.005441f
C3101 VDD.n2587 GND 0.005441f
C3102 VDD.n2588 GND 0.005441f
C3103 VDD.n2589 GND 0.362306f
C3104 VDD.n2590 GND 0.005441f
C3105 VDD.n2591 GND 0.005441f
C3106 VDD.n2592 GND 0.005441f
C3107 VDD.n2593 GND 0.005441f
C3108 VDD.n2594 GND 0.005441f
C3109 VDD.n2595 GND 0.362306f
C3110 VDD.n2596 GND 0.005441f
C3111 VDD.n2597 GND 0.005441f
C3112 VDD.n2598 GND 0.005441f
C3113 VDD.n2599 GND 0.005441f
C3114 VDD.n2600 GND 0.005441f
C3115 VDD.n2601 GND 0.194473f
C3116 VDD.n2602 GND 0.005441f
C3117 VDD.n2603 GND 0.005441f
C3118 VDD.n2604 GND 0.005441f
C3119 VDD.n2605 GND 0.005441f
C3120 VDD.n2606 GND 0.005441f
C3121 VDD.n2607 GND 0.362306f
C3122 VDD.n2608 GND 0.005441f
C3123 VDD.n2609 GND 0.005441f
C3124 VDD.n2610 GND 0.005441f
C3125 VDD.n2611 GND 0.005441f
C3126 VDD.n2612 GND 0.005441f
C3127 VDD.n2613 GND 0.362306f
C3128 VDD.n2614 GND 0.005441f
C3129 VDD.n2615 GND 0.005441f
C3130 VDD.n2616 GND 0.005441f
C3131 VDD.n2617 GND 0.005441f
C3132 VDD.n2618 GND 0.005441f
C3133 VDD.n2619 GND 0.362306f
C3134 VDD.n2620 GND 0.005441f
C3135 VDD.n2621 GND 0.005441f
C3136 VDD.n2622 GND 0.005441f
C3137 VDD.n2623 GND 0.005441f
C3138 VDD.n2624 GND 0.005441f
C3139 VDD.n2625 GND 0.314354f
C3140 VDD.n2626 GND 0.005441f
C3141 VDD.n2627 GND 0.005441f
C3142 VDD.n2628 GND 0.005441f
C3143 VDD.n2629 GND 0.005441f
C3144 VDD.n2630 GND 0.005441f
C3145 VDD.n2631 GND 0.005441f
C3146 VDD.n2632 GND 0.005441f
C3147 VDD.n2633 GND 0.005441f
C3148 VDD.n2634 GND 0.005441f
C3149 VDD.n2635 GND 0.005441f
C3150 VDD.n2636 GND 0.317018f
C3151 VDD.n2637 GND 0.005441f
C3152 VDD.n2638 GND 0.005441f
C3153 VDD.n2639 GND 0.005441f
C3154 VDD.n2640 GND 0.005441f
C3155 VDD.n2641 GND 0.005441f
C3156 VDD.n2642 GND 0.362306f
C3157 VDD.n2643 GND 0.005441f
C3158 VDD.n2644 GND 0.005441f
C3159 VDD.n2645 GND 0.005441f
C3160 VDD.n2646 GND 0.005441f
C3161 VDD.n2647 GND 0.012652f
C3162 VDD.n2648 GND 0.011992f
C3163 VDD.n2649 GND 0.013054f
C3164 VDD.n2650 GND 0.012394f
C3165 VDD.n2651 GND 0.004841f
C3166 VDD.n2652 GND 0.005441f
C3167 VDD.n2653 GND 0.005441f
C3168 VDD.n2654 GND 0.003321f
C3169 VDD.n2655 GND 0.005441f
C3170 VDD.n2656 GND 0.005441f
C3171 VDD.n2657 GND 0.005441f
C3172 VDD.n2658 GND 0.005441f
C3173 VDD.n2659 GND 0.005441f
C3174 VDD.n2660 GND 0.005441f
C3175 VDD.n2661 GND 0.005441f
C3176 VDD.n2662 GND 0.005441f
C3177 VDD.n2663 GND 0.005441f
C3178 VDD.n2664 GND 0.005441f
C3179 VDD.n2665 GND 0.005441f
C3180 VDD.n2666 GND 0.005441f
C3181 VDD.n2667 GND 0.005441f
C3182 VDD.n2668 GND 0.005441f
C3183 VDD.n2669 GND 0.005441f
C3184 VDD.n2670 GND 0.005441f
C3185 VDD.n2671 GND 0.005441f
C3186 VDD.n2672 GND 0.005441f
C3187 VDD.n2673 GND 0.005441f
C3188 VDD.n2674 GND 0.005441f
C3189 VDD.n2675 GND 0.005441f
C3190 VDD.n2676 GND 0.005441f
C3191 VDD.n2677 GND 0.005441f
C3192 VDD.n2678 GND 0.005441f
C3193 VDD.n2679 GND 0.005441f
C3194 VDD.n2680 GND 0.005441f
C3195 VDD.n2681 GND 0.005441f
C3196 VDD.n2682 GND 0.005441f
C3197 VDD.n2683 GND 0.005441f
C3198 VDD.n2684 GND 0.005441f
C3199 VDD.n2685 GND 0.005441f
C3200 VDD.n2686 GND 0.005441f
C3201 VDD.n2687 GND 0.005441f
C3202 VDD.n2688 GND 0.005441f
C3203 VDD.n2689 GND 0.005441f
C3204 VDD.n2690 GND 0.005441f
C3205 VDD.n2691 GND 0.013054f
C3206 VDD.n2692 GND 0.013054f
C3207 VDD.n2693 GND 0.011992f
C3208 VDD.n2694 GND 0.005441f
C3209 VDD.n2695 GND 0.005441f
C3210 VDD.n2696 GND 0.362306f
C3211 VDD.n2697 GND 0.005441f
C3212 VDD.n2698 GND 0.011992f
C3213 VDD.n2699 GND 0.012652f
C3214 VDD.n2700 GND 0.012394f
C3215 VDD.n2701 GND 0.005441f
C3216 VDD.n2702 GND 0.004841f
C3217 VDD.n2703 GND 0.007776f
C3218 VDD.n2704 GND 0.003321f
C3219 VDD.n2705 GND 0.005441f
C3220 VDD.n2706 GND 0.005441f
C3221 VDD.n2707 GND 0.005441f
C3222 VDD.n2708 GND 0.005441f
C3223 VDD.n2709 GND 0.005441f
C3224 VDD.n2710 GND 0.005441f
C3225 VDD.n2711 GND 0.005441f
C3226 VDD.n2712 GND 0.005441f
C3227 VDD.n2713 GND 0.005441f
C3228 VDD.n2714 GND 0.005441f
C3229 VDD.n2715 GND 0.005441f
C3230 VDD.n2716 GND 0.005441f
C3231 VDD.n2717 GND 0.005441f
C3232 VDD.n2718 GND 0.005441f
C3233 VDD.n2719 GND 0.005441f
C3234 VDD.n2720 GND 0.005441f
C3235 VDD.n2721 GND 0.005441f
C3236 VDD.n2722 GND 0.005441f
C3237 VDD.n2723 GND 0.005441f
C3238 VDD.n2724 GND 0.005441f
C3239 VDD.n2725 GND 0.005441f
C3240 VDD.n2726 GND 0.005441f
C3241 VDD.n2727 GND 0.005441f
C3242 VDD.n2728 GND 0.005441f
C3243 VDD.n2729 GND 0.005441f
C3244 VDD.n2730 GND 0.005441f
C3245 VDD.n2731 GND 0.005441f
C3246 VDD.n2732 GND 0.005441f
C3247 VDD.n2733 GND 0.005441f
C3248 VDD.n2734 GND 0.005441f
C3249 VDD.n2735 GND 0.005441f
C3250 VDD.n2736 GND 0.005441f
C3251 VDD.n2737 GND 0.005441f
C3252 VDD.n2738 GND 0.005441f
C3253 VDD.n2739 GND 0.005441f
C3254 VDD.n2740 GND 0.005441f
C3255 VDD.n2741 GND 0.013054f
C3256 VDD.n2742 GND 0.013054f
C3257 VDD.n2743 GND 2.29372f
C3258 VDD.n2744 GND 2.29372f
C3259 VDD.n2745 GND 0.011992f
C3260 VDD.n2746 GND 0.011992f
C3261 VDD.n2747 GND 0.013054f
C3262 VDD.n2748 GND 0.005441f
C3263 VDD.n2749 GND 0.005441f
C3264 VDD.n2750 GND 0.005441f
C3265 VDD.n2751 GND 0.005441f
C3266 VDD.n2752 GND 0.005441f
C3267 VDD.n2753 GND 0.005441f
C3268 VDD.n2754 GND 0.005441f
C3269 VDD.n2755 GND 0.005441f
C3270 VDD.n2756 GND 0.005441f
C3271 VDD.n2757 GND 0.005441f
C3272 VDD.t89 GND 0.111051f
C3273 VDD.t90 GND 0.129192f
C3274 VDD.t87 GND 0.629305f
C3275 VDD.n2758 GND 0.086428f
C3276 VDD.n2759 GND 0.052244f
C3277 VDD.n2760 GND 0.005441f
C3278 VDD.n2761 GND 0.005441f
C3279 VDD.n2762 GND 0.005441f
C3280 VDD.n2763 GND 0.005441f
C3281 VDD.n2764 GND 0.005441f
C3282 VDD.n2765 GND 0.005441f
C3283 VDD.n2766 GND 0.005441f
C3284 VDD.n2767 GND 0.005441f
C3285 VDD.n2768 GND 0.005441f
C3286 VDD.n2769 GND 0.005441f
C3287 VDD.n2770 GND 0.005441f
C3288 VDD.n2771 GND 0.005441f
C3289 VDD.n2772 GND 0.005441f
C3290 VDD.n2773 GND 0.005441f
C3291 VDD.n2774 GND 0.005441f
C3292 VDD.n2775 GND 0.005441f
C3293 VDD.n2776 GND 0.005441f
C3294 VDD.n2777 GND 0.005441f
C3295 VDD.n2778 GND 0.005441f
C3296 VDD.n2779 GND 0.005441f
C3297 VDD.n2780 GND 0.004841f
C3298 VDD.n2781 GND 0.005441f
C3299 VDD.n2782 GND 0.005441f
C3300 VDD.n2783 GND 0.005441f
C3301 VDD.n2784 GND 0.005441f
C3302 VDD.n2785 GND 0.005441f
C3303 VDD.n2786 GND 0.005441f
C3304 VDD.n2787 GND 0.005441f
C3305 VDD.n2788 GND 0.005441f
C3306 VDD.n2789 GND 0.005441f
C3307 VDD.n2791 GND 0.005441f
C3308 VDD.n2792 GND 0.005441f
C3309 VDD.n2793 GND 0.005441f
C3310 VDD.n2794 GND 0.005441f
C3311 VDD.n2795 GND 0.005441f
C3312 VDD.n2797 GND 0.005441f
C3313 VDD.n2799 GND 0.005441f
C3314 VDD.n2800 GND 0.005441f
C3315 VDD.n2801 GND 0.005441f
C3316 VDD.n2802 GND 0.005441f
C3317 VDD.n2803 GND 0.005441f
C3318 VDD.n2805 GND 0.005441f
C3319 VDD.n2807 GND 0.005441f
C3320 VDD.n2808 GND 0.005441f
C3321 VDD.n2809 GND 0.005441f
C3322 VDD.n2810 GND 0.005441f
C3323 VDD.n2811 GND 0.005441f
C3324 VDD.n2813 GND 0.005441f
C3325 VDD.n2815 GND 0.005441f
C3326 VDD.n2816 GND 0.005441f
C3327 VDD.n2817 GND 0.005441f
C3328 VDD.n2818 GND 0.005441f
C3329 VDD.n2819 GND 0.005441f
C3330 VDD.n2821 GND 0.005441f
C3331 VDD.n2823 GND 0.005441f
C3332 VDD.n2824 GND 0.005441f
C3333 VDD.n2825 GND 0.005441f
C3334 VDD.t92 GND 0.111051f
C3335 VDD.t93 GND 0.129192f
C3336 VDD.t91 GND 0.629305f
C3337 VDD.n2826 GND 0.086428f
C3338 VDD.n2827 GND 0.052244f
C3339 VDD.n2828 GND 0.007776f
C3340 VDD.n2829 GND 0.003321f
C3341 VDD.n2830 GND 0.005441f
C3342 VDD.n2832 GND 0.005441f
C3343 VDD.n2833 GND 0.013054f
C3344 VDD.n2834 GND 0.013054f
C3345 VDD.n2835 GND 0.011992f
C3346 VDD.n2836 GND 0.005441f
C3347 VDD.n2837 GND 0.005441f
C3348 VDD.n2838 GND 0.005441f
C3349 VDD.n2839 GND 0.005441f
C3350 VDD.n2840 GND 0.005441f
C3351 VDD.n2841 GND 0.005441f
C3352 VDD.n2842 GND 0.005441f
C3353 VDD.n2843 GND 0.005441f
C3354 VDD.n2844 GND 0.005441f
C3355 VDD.n2845 GND 0.005441f
C3356 VDD.n2846 GND 0.005441f
C3357 VDD.n2847 GND 0.005441f
C3358 VDD.n2848 GND 0.005441f
C3359 VDD.n2849 GND 0.005441f
C3360 VDD.n2850 GND 0.005441f
C3361 VDD.n2851 GND 0.005441f
C3362 VDD.n2852 GND 0.005441f
C3363 VDD.n2853 GND 0.005441f
C3364 VDD.n2854 GND 0.005441f
C3365 VDD.n2855 GND 0.005441f
C3366 VDD.n2856 GND 0.005441f
C3367 VDD.n2857 GND 0.005441f
C3368 VDD.n2858 GND 0.005441f
C3369 VDD.n2859 GND 0.005441f
C3370 VDD.n2860 GND 0.005441f
C3371 VDD.n2861 GND 0.005441f
C3372 VDD.n2862 GND 0.005441f
C3373 VDD.n2863 GND 0.005441f
C3374 VDD.n2864 GND 0.005441f
C3375 VDD.n2865 GND 0.005441f
C3376 VDD.n2866 GND 0.005441f
C3377 VDD.n2867 GND 0.005441f
C3378 VDD.n2868 GND 0.005441f
C3379 VDD.n2869 GND 0.005441f
C3380 VDD.n2870 GND 0.005441f
C3381 VDD.n2871 GND 0.005441f
C3382 VDD.n2872 GND 0.005441f
C3383 VDD.n2873 GND 0.005441f
C3384 VDD.n2874 GND 0.005441f
C3385 VDD.n2875 GND 0.005441f
C3386 VDD.n2876 GND 0.005441f
C3387 VDD.n2877 GND 0.005441f
C3388 VDD.n2878 GND 0.005441f
C3389 VDD.n2879 GND 0.005441f
C3390 VDD.n2880 GND 0.005441f
C3391 VDD.n2881 GND 0.005441f
C3392 VDD.n2882 GND 0.005441f
C3393 VDD.n2883 GND 0.005441f
C3394 VDD.n2884 GND 0.005441f
C3395 VDD.n2885 GND 0.005441f
C3396 VDD.n2886 GND 0.005441f
C3397 VDD.n2887 GND 0.005441f
C3398 VDD.n2888 GND 0.005441f
C3399 VDD.n2889 GND 0.005441f
C3400 VDD.n2890 GND 0.005441f
C3401 VDD.n2891 GND 0.005441f
C3402 VDD.n2892 GND 0.005441f
C3403 VDD.n2893 GND 0.005441f
C3404 VDD.n2894 GND 0.005441f
C3405 VDD.n2895 GND 0.005441f
C3406 VDD.n2896 GND 0.005441f
C3407 VDD.n2897 GND 0.005441f
C3408 VDD.n2898 GND 0.005441f
C3409 VDD.n2899 GND 0.005441f
C3410 VDD.n2900 GND 0.005441f
C3411 VDD.n2901 GND 0.005441f
C3412 VDD.n2902 GND 0.005441f
C3413 VDD.n2903 GND 0.005441f
C3414 VDD.n2904 GND 0.005441f
C3415 VDD.n2905 GND 0.005441f
C3416 VDD.n2906 GND 0.005441f
C3417 VDD.n2907 GND 0.005441f
C3418 VDD.n2908 GND 0.005441f
C3419 VDD.n2909 GND 0.005441f
C3420 VDD.n2910 GND 0.005441f
C3421 VDD.n2911 GND 0.005441f
C3422 VDD.n2912 GND 0.005441f
C3423 VDD.n2913 GND 0.005441f
C3424 VDD.n2914 GND 0.005441f
C3425 VDD.n2915 GND 0.005441f
C3426 VDD.n2916 GND 0.005441f
C3427 VDD.n2917 GND 0.005441f
C3428 VDD.n2918 GND 0.005441f
C3429 VDD.n2919 GND 0.005441f
C3430 VDD.n2920 GND 0.005441f
C3431 VDD.n2921 GND 0.005441f
C3432 VDD.n2922 GND 0.005441f
C3433 VDD.n2923 GND 0.005441f
C3434 VDD.n2924 GND 0.005441f
C3435 VDD.n2925 GND 0.005441f
C3436 VDD.n2926 GND 0.005441f
C3437 VDD.n2927 GND 0.005441f
C3438 VDD.n2928 GND 0.005441f
C3439 VDD.n2929 GND 0.005441f
C3440 VDD.n2930 GND 0.005441f
C3441 VDD.n2931 GND 0.005441f
C3442 VDD.n2932 GND 0.005441f
C3443 VDD.n2933 GND 0.005441f
C3444 VDD.n2934 GND 0.005441f
C3445 VDD.n2935 GND 0.005441f
C3446 VDD.n2936 GND 0.005441f
C3447 VDD.n2937 GND 0.005441f
C3448 VDD.n2938 GND 0.005441f
C3449 VDD.n2939 GND 0.005441f
C3450 VDD.n2940 GND 0.005441f
C3451 VDD.n2941 GND 0.005441f
C3452 VDD.n2942 GND 0.005441f
C3453 VDD.n2943 GND 0.005441f
C3454 VDD.n2944 GND 0.005441f
C3455 VDD.n2945 GND 0.005441f
C3456 VDD.n2946 GND 0.005441f
C3457 VDD.n2947 GND 0.005441f
C3458 VDD.n2948 GND 0.005441f
C3459 VDD.n2949 GND 0.005441f
C3460 VDD.n2950 GND 0.005441f
C3461 VDD.n2951 GND 0.005441f
C3462 VDD.n2952 GND 0.005441f
C3463 VDD.n2953 GND 0.005441f
C3464 VDD.n2954 GND 0.005441f
C3465 VDD.n2955 GND 0.005441f
C3466 VDD.n2956 GND 0.050616f
C3467 VDD.n2957 GND 0.005441f
C3468 VDD.n2958 GND 0.005441f
C3469 VDD.n2959 GND 0.005441f
C3470 VDD.n2960 GND 0.005441f
C3471 VDD.n2961 GND 0.005441f
C3472 VDD.n2962 GND 0.005441f
C3473 VDD.n2963 GND 0.005441f
C3474 VDD.n2964 GND 0.005441f
C3475 VDD.n2965 GND 0.005441f
C3476 VDD.n2966 GND 0.005441f
C3477 VDD.n2967 GND 0.005441f
C3478 VDD.n2968 GND 0.005441f
C3479 VDD.n2969 GND 0.005441f
C3480 VDD.n2970 GND 0.005441f
C3481 VDD.n2971 GND 0.005441f
C3482 VDD.n2972 GND 0.005441f
C3483 VDD.n2973 GND 0.005441f
C3484 VDD.n2974 GND 0.005441f
C3485 VDD.n2975 GND 0.005441f
C3486 VDD.n2976 GND 0.005441f
C3487 VDD.n2977 GND 0.005441f
C3488 VDD.n2978 GND 0.005441f
C3489 VDD.n2979 GND 0.005441f
C3490 VDD.n2980 GND 0.005441f
C3491 VDD.n2981 GND 0.005441f
C3492 VDD.n2982 GND 0.005441f
C3493 VDD.n2983 GND 0.005441f
C3494 VDD.n2984 GND 0.005441f
C3495 VDD.n2985 GND 0.005441f
C3496 VDD.n2986 GND 0.005441f
C3497 VDD.n2987 GND 0.005441f
C3498 VDD.n2988 GND 0.005441f
C3499 VDD.n2989 GND 0.005441f
C3500 VDD.n2990 GND 0.005441f
C3501 VDD.n2991 GND 0.005441f
C3502 VDD.n2992 GND 0.005441f
C3503 VDD.n2993 GND 0.005441f
C3504 VDD.n2994 GND 0.005441f
C3505 VDD.n2995 GND 0.005441f
C3506 VDD.n2996 GND 0.005441f
C3507 VDD.n2997 GND 0.005441f
C3508 VDD.n2998 GND 0.005441f
C3509 VDD.n2999 GND 0.005441f
C3510 VDD.n3000 GND 0.005441f
C3511 VDD.n3001 GND 0.005441f
C3512 VDD.n3002 GND 0.005441f
C3513 VDD.n3003 GND 0.005441f
C3514 VDD.n3004 GND 0.005441f
C3515 VDD.n3005 GND 0.005441f
C3516 VDD.n3006 GND 0.005441f
C3517 VDD.n3007 GND 0.005441f
C3518 VDD.n3008 GND 0.005441f
C3519 VDD.n3009 GND 0.005441f
C3520 VDD.n3010 GND 0.005441f
C3521 VDD.n3011 GND 0.005441f
C3522 VDD.n3012 GND 0.005441f
C3523 VDD.n3013 GND 0.005441f
C3524 VDD.n3014 GND 0.005441f
C3525 VDD.n3015 GND 0.005441f
C3526 VDD.n3016 GND 0.005441f
C3527 VDD.n3017 GND 0.005441f
C3528 VDD.n3018 GND 0.005441f
C3529 VDD.n3019 GND 0.005441f
C3530 VDD.n3020 GND 0.005441f
C3531 VDD.n3021 GND 0.005441f
C3532 VDD.n3022 GND 0.005441f
C3533 VDD.n3023 GND 0.005441f
C3534 VDD.n3024 GND 0.005441f
C3535 VDD.n3025 GND 0.005441f
C3536 VDD.n3026 GND 0.005441f
C3537 VDD.n3027 GND 0.005441f
C3538 VDD.n3028 GND 0.005441f
C3539 VDD.n3029 GND 0.005441f
C3540 VDD.n3030 GND 0.005441f
C3541 VDD.n3031 GND 0.005441f
C3542 VDD.n3032 GND 0.005441f
C3543 VDD.n3033 GND 0.005441f
C3544 VDD.n3034 GND 0.005441f
C3545 VDD.n3035 GND 0.005441f
C3546 VDD.n3036 GND 0.005441f
C3547 VDD.n3037 GND 0.005441f
C3548 VDD.n3038 GND 0.005441f
C3549 VDD.n3039 GND 0.005441f
C3550 VDD.n3040 GND 0.005441f
C3551 VDD.n3041 GND 0.005441f
C3552 VDD.n3042 GND 0.005441f
C3553 VDD.n3043 GND 0.005441f
C3554 VDD.n3044 GND 0.005441f
C3555 VDD.n3045 GND 0.005441f
C3556 VDD.n3046 GND 0.005441f
C3557 VDD.n3047 GND 0.005441f
C3558 VDD.n3048 GND 0.005441f
C3559 VDD.n3049 GND 0.005441f
C3560 VDD.n3050 GND 0.005441f
C3561 VDD.n3051 GND 0.005441f
C3562 VDD.n3052 GND 0.011992f
C3563 VDD.n3054 GND 0.013054f
C3564 VDD.n3055 GND 0.013054f
C3565 VDD.n3056 GND 0.004841f
C3566 VDD.n3057 GND 0.007776f
C3567 VDD.n3058 GND 0.003321f
C3568 VDD.n3059 GND 0.005441f
C3569 VDD.n3061 GND 0.005441f
C3570 VDD.n3063 GND 0.005441f
C3571 VDD.n3064 GND 0.005441f
C3572 VDD.n3065 GND 0.005441f
C3573 VDD.n3066 GND 0.005441f
C3574 VDD.n3067 GND 0.005441f
C3575 VDD.n3069 GND 0.005441f
C3576 VDD.n3071 GND 0.005441f
C3577 VDD.n3072 GND 0.005441f
C3578 VDD.n3073 GND 0.005441f
C3579 VDD.n3074 GND 0.005441f
C3580 VDD.n3075 GND 0.005441f
C3581 VDD.n3077 GND 0.005441f
C3582 VDD.n3079 GND 0.005441f
C3583 VDD.n3080 GND 0.005441f
C3584 VDD.n3081 GND 0.005441f
C3585 VDD.n3082 GND 0.005441f
C3586 VDD.n3083 GND 0.005441f
C3587 VDD.n3085 GND 0.005441f
C3588 VDD.n3087 GND 0.005441f
C3589 VDD.n3088 GND 0.005441f
C3590 VDD.n3089 GND 0.005441f
C3591 VDD.n3090 GND 0.005441f
C3592 VDD.n3091 GND 0.005441f
C3593 VDD.n3093 GND 0.005441f
C3594 VDD.n3095 GND 0.005441f
C3595 VDD.n3096 GND 0.005441f
C3596 VDD.n3097 GND 0.013054f
C3597 VDD.n3098 GND 0.011992f
C3598 VDD.n3099 GND 0.011992f
C3599 VDD.n3100 GND 0.540796f
C3600 VDD.n3101 GND 0.011992f
C3601 VDD.n3102 GND 0.011992f
C3602 VDD.n3103 GND 0.005441f
C3603 VDD.n3104 GND 0.005441f
C3604 VDD.n3105 GND 0.005441f
C3605 VDD.n3106 GND 0.362306f
C3606 VDD.n3107 GND 0.005441f
C3607 VDD.n3108 GND 0.005441f
C3608 VDD.n3109 GND 0.005441f
C3609 VDD.n3110 GND 0.005441f
C3610 VDD.n3111 GND 0.005441f
C3611 VDD.n3112 GND 0.226442f
C3612 VDD.n3113 GND 0.005441f
C3613 VDD.n3114 GND 0.005441f
C3614 VDD.n3115 GND 0.005441f
C3615 VDD.n3116 GND 0.005441f
C3616 VDD.n3117 GND 0.005441f
C3617 VDD.n3118 GND 0.229106f
C3618 VDD.n3119 GND 0.005441f
C3619 VDD.n3120 GND 0.005441f
C3620 VDD.n3121 GND 0.005441f
C3621 VDD.n3122 GND 0.005441f
C3622 VDD.n3123 GND 0.005441f
C3623 VDD.n3124 GND 0.362306f
C3624 VDD.n3125 GND 0.005441f
C3625 VDD.n3126 GND 0.005441f
C3626 VDD.n3127 GND 0.005441f
C3627 VDD.n3128 GND 0.005441f
C3628 VDD.n3129 GND 0.005441f
C3629 VDD.n3130 GND 0.362306f
C3630 VDD.n3131 GND 0.005441f
C3631 VDD.n3132 GND 0.005441f
C3632 VDD.n3133 GND 0.005441f
C3633 VDD.n3134 GND 0.005441f
C3634 VDD.n3135 GND 0.005441f
C3635 VDD.n3136 GND 0.362306f
C3636 VDD.n3137 GND 0.005441f
C3637 VDD.n3138 GND 0.005441f
C3638 VDD.n3139 GND 0.005441f
C3639 VDD.n3140 GND 0.005441f
C3640 VDD.n3141 GND 0.005441f
C3641 VDD.n3142 GND 0.348986f
C3642 VDD.n3143 GND 0.005441f
C3643 VDD.n3144 GND 0.005441f
C3644 VDD.n3145 GND 0.005441f
C3645 VDD.n3146 GND 0.005441f
C3646 VDD.n3147 GND 0.005441f
C3647 VDD.n3148 GND 0.362306f
C3648 VDD.n3149 GND 0.005441f
C3649 VDD.n3150 GND 0.005441f
C3650 VDD.n3151 GND 0.005441f
C3651 VDD.n3152 GND 0.005441f
C3652 VDD.n3153 GND 0.005441f
C3653 VDD.n3154 GND 0.362306f
C3654 VDD.n3155 GND 0.005441f
C3655 VDD.n3156 GND 0.005441f
C3656 VDD.n3157 GND 0.005441f
C3657 VDD.n3158 GND 0.005441f
C3658 VDD.n3159 GND 0.005441f
C3659 VDD.n3160 GND 0.207793f
C3660 VDD.n3161 GND 0.005441f
C3661 VDD.n3162 GND 0.005441f
C3662 VDD.n3163 GND 0.005441f
C3663 VDD.n3164 GND 0.005441f
C3664 VDD.n3165 GND 0.005441f
C3665 VDD.n3166 GND 0.362306f
C3666 VDD.n3167 GND 0.005441f
C3667 VDD.n3168 GND 0.005441f
C3668 VDD.n3169 GND 0.005441f
C3669 VDD.n3170 GND 0.005441f
C3670 VDD.n3171 GND 0.005441f
C3671 VDD.n3172 GND 0.362306f
C3672 VDD.n3173 GND 0.005441f
C3673 VDD.n3174 GND 0.005441f
C3674 VDD.n3175 GND 0.005441f
C3675 VDD.n3176 GND 0.005441f
C3676 VDD.n3177 GND 0.005441f
C3677 VDD.n3178 GND 0.253082f
C3678 VDD.n3179 GND 0.005441f
C3679 VDD.n3180 GND 0.005441f
C3680 VDD.n3181 GND 0.005441f
C3681 VDD.n3182 GND 0.005441f
C3682 VDD.n3183 GND 0.005441f
C3683 VDD.n3184 GND 0.362306f
C3684 VDD.n3185 GND 0.005441f
C3685 VDD.n3186 GND 0.005441f
C3686 VDD.n3187 GND 0.005441f
C3687 VDD.n3188 GND 0.005441f
C3688 VDD.n3189 GND 0.005441f
C3689 VDD.n3190 GND 0.330338f
C3690 VDD.n3191 GND 0.005441f
C3691 VDD.n3192 GND 0.005441f
C3692 VDD.n3193 GND 0.005441f
C3693 VDD.n3194 GND 0.005441f
C3694 VDD.n3195 GND 0.005441f
C3695 VDD.n3196 GND 0.362306f
C3696 VDD.n3197 GND 0.005441f
C3697 VDD.n3198 GND 0.005441f
C3698 VDD.n3199 GND 0.005441f
C3699 VDD.n3200 GND 0.005441f
C3700 VDD.n3201 GND 0.005441f
C3701 VDD.n3202 GND 0.362306f
C3702 VDD.n3203 GND 0.005441f
C3703 VDD.n3204 GND 0.005441f
C3704 VDD.n3205 GND 0.005441f
C3705 VDD.n3206 GND 0.005441f
C3706 VDD.n3207 GND 0.005441f
C3707 VDD.n3208 GND 0.23177f
C3708 VDD.n3209 GND 0.005441f
C3709 VDD.n3210 GND 0.005441f
C3710 VDD.n3211 GND 0.005441f
C3711 VDD.n3212 GND 0.005441f
C3712 VDD.n3213 GND 0.005441f
C3713 VDD.n3214 GND 0.362306f
C3714 VDD.n3215 GND 0.005441f
C3715 VDD.n3216 GND 0.005441f
C3716 VDD.n3217 GND 0.005441f
C3717 VDD.n3218 GND 0.005441f
C3718 VDD.n3219 GND 0.005441f
C3719 VDD.n3220 GND 0.362306f
C3720 VDD.n3221 GND 0.005441f
C3721 VDD.n3222 GND 0.005441f
C3722 VDD.n3223 GND 0.005441f
C3723 VDD.n3224 GND 0.005441f
C3724 VDD.n3225 GND 0.005441f
C3725 VDD.n3226 GND 0.27173f
C3726 VDD.n3227 GND 0.005441f
C3727 VDD.n3228 GND 0.005441f
C3728 VDD.n3229 GND 0.005441f
C3729 VDD.n3230 GND 0.005441f
C3730 VDD.n3231 GND 0.005441f
C3731 VDD.n3232 GND 0.362306f
C3732 VDD.n3233 GND 0.005441f
C3733 VDD.n3234 GND 0.005441f
C3734 VDD.n3235 GND 0.005441f
C3735 VDD.n3236 GND 0.005441f
C3736 VDD.n3237 GND 0.005441f
C3737 VDD.n3238 GND 0.362306f
C3738 VDD.n3239 GND 0.005441f
C3739 VDD.n3240 GND 0.005441f
C3740 VDD.n3241 GND 0.005441f
C3741 VDD.n3242 GND 0.005441f
C3742 VDD.n3243 GND 0.005441f
C3743 VDD.n3244 GND 0.362306f
C3744 VDD.n3245 GND 0.005441f
C3745 VDD.n3246 GND 0.005441f
C3746 VDD.n3247 GND 0.005441f
C3747 VDD.n3248 GND 0.005441f
C3748 VDD.n3249 GND 0.005441f
C3749 VDD.n3250 GND 0.362306f
C3750 VDD.n3251 GND 0.005441f
C3751 VDD.n3252 GND 0.005441f
C3752 VDD.n3253 GND 0.005441f
C3753 VDD.n3254 GND 0.005441f
C3754 VDD.n3255 GND 0.005441f
C3755 VDD.n3256 GND 0.213121f
C3756 VDD.n3257 GND 0.005441f
C3757 VDD.n3258 GND 0.005441f
C3758 VDD.n3259 GND 0.005441f
C3759 VDD.n3260 GND 0.005441f
C3760 VDD.n3261 GND 0.005441f
C3761 VDD.n3262 GND 0.362306f
C3762 VDD.n3263 GND 0.005441f
C3763 VDD.n3264 GND 0.005441f
C3764 VDD.n3265 GND 0.005441f
C3765 VDD.n3266 GND 0.005441f
C3766 VDD.n3267 GND 0.005441f
C3767 VDD.n3268 GND 0.362306f
C3768 VDD.n3269 GND 0.005441f
C3769 VDD.n3270 GND 0.005441f
C3770 VDD.n3271 GND 0.005441f
C3771 VDD.n3272 GND 0.005441f
C3772 VDD.n3273 GND 0.005441f
C3773 VDD.n3274 GND 0.362306f
C3774 VDD.n3275 GND 0.005441f
C3775 VDD.n3276 GND 0.005441f
C3776 VDD.n3277 GND 0.005441f
C3777 VDD.n3278 GND 0.005441f
C3778 VDD.n3279 GND 0.005441f
C3779 VDD.n3280 GND 0.362306f
C3780 VDD.n3281 GND 0.005441f
C3781 VDD.n3282 GND 0.005441f
C3782 VDD.n3283 GND 0.005441f
C3783 VDD.n3284 GND 0.005441f
C3784 VDD.n3285 GND 0.005441f
C3785 VDD.n3286 GND 0.335666f
C3786 VDD.n3287 GND 0.005441f
C3787 VDD.n3288 GND 0.005441f
C3788 VDD.n3289 GND 0.005441f
C3789 VDD.n3290 GND 0.005441f
C3790 VDD.n3291 GND 0.005441f
C3791 VDD.n3292 GND 0.33833f
C3792 VDD.n3293 GND 0.005441f
C3793 VDD.n3294 GND 0.005441f
C3794 VDD.n3295 GND 0.005441f
C3795 VDD.n3296 GND 0.005441f
C3796 VDD.n3297 GND 0.005441f
C3797 VDD.n3298 GND 0.362306f
C3798 VDD.n3299 GND 0.005441f
C3799 VDD.n3300 GND 0.005441f
C3800 VDD.n3301 GND 0.005441f
C3801 VDD.n3302 GND 0.005441f
C3802 VDD.n3303 GND 0.005441f
C3803 VDD.n3304 GND 0.362306f
C3804 VDD.n3305 GND 0.005441f
C3805 VDD.n3306 GND 0.005441f
C3806 VDD.n3307 GND 0.005441f
C3807 VDD.n3308 GND 0.005441f
C3808 VDD.n3309 GND 0.005441f
C3809 VDD.n3310 GND 0.362306f
C3810 VDD.n3311 GND 0.005441f
C3811 VDD.n3312 GND 0.005441f
C3812 VDD.n3313 GND 0.005441f
C3813 VDD.n3314 GND 0.005441f
C3814 VDD.n3315 GND 0.005441f
C3815 VDD.n3316 GND 0.362306f
C3816 VDD.n3317 GND 0.005441f
C3817 VDD.n3318 GND 0.005441f
C3818 VDD.n3319 GND 0.005441f
C3819 VDD.n3320 GND 0.005441f
C3820 VDD.n3321 GND 0.005441f
C3821 VDD.n3322 GND 0.215785f
C3822 VDD.n3323 GND 0.005441f
C3823 VDD.n3324 GND 0.005441f
C3824 VDD.n3325 GND 0.005441f
C3825 VDD.n3326 GND 0.005441f
C3826 VDD.n3327 GND 0.005441f
C3827 VDD.n3328 GND 0.005441f
C3828 VDD.n3329 GND 0.005441f
C3829 VDD.n3330 GND 0.314354f
C3830 VDD.n3331 GND 0.005441f
C3831 VDD.n3332 GND 0.005441f
C3832 VDD.n3333 GND 0.005441f
C3833 VDD.n3334 GND 0.005441f
C3834 VDD.n3335 GND 0.005441f
C3835 VDD.n3336 GND 0.362306f
C3836 VDD.n3337 GND 0.005441f
C3837 VDD.n3338 GND 0.005441f
C3838 VDD.n3339 GND 0.005441f
C3839 VDD.n3340 GND 0.005441f
C3840 VDD.n3341 GND 0.005441f
C3841 VDD.n3342 GND 0.005441f
C3842 VDD.n3343 GND 0.005441f
C3843 VDD.n3344 GND 0.012652f
C3844 VDD.n3346 GND 0.011992f
C3845 VDD.n3347 GND 0.013054f
C3846 VDD.n3348 GND 0.012394f
C3847 VDD.n3349 GND 0.004841f
C3848 VDD.n3350 GND 0.007776f
C3849 VDD.n3351 GND 0.003321f
C3850 VDD.n3352 GND 0.005441f
C3851 VDD.n3354 GND 0.005441f
C3852 VDD.n3355 GND 0.005441f
C3853 VDD.n3356 GND 0.005441f
C3854 VDD.n3357 GND 0.005441f
C3855 VDD.n3358 GND 0.005441f
C3856 VDD.n3359 GND 0.005441f
C3857 VDD.n3361 GND 0.005441f
C3858 VDD.n3362 GND 0.005441f
C3859 VDD.n3363 GND 0.005441f
C3860 VDD.n3364 GND 0.005441f
C3861 VDD.n3365 GND 0.004081f
C3862 VDD.n3366 GND 0.005441f
C3863 VDD.n3368 GND 0.005441f
C3864 VDD.n3369 GND 0.004081f
C3865 VDD.n3370 GND 0.005441f
C3866 VDD.n3371 GND 0.005441f
C3867 VDD.n3373 GND 0.005441f
C3868 VDD.n3374 GND 0.005441f
C3869 VDD.n3375 GND 0.005441f
C3870 VDD.n3376 GND 0.005441f
C3871 VDD.n3377 GND 0.005441f
C3872 VDD.n3378 GND 0.005441f
C3873 VDD.n3380 GND 0.005441f
C3874 VDD.n3381 GND 0.005441f
C3875 VDD.n3382 GND 0.005441f
C3876 VDD.n3383 GND 0.005441f
C3877 VDD.n3384 GND 0.005441f
C3878 VDD.n3385 GND 0.005441f
C3879 VDD.n3387 GND 0.013054f
C3880 VDD.n3388 GND 0.011992f
C3881 VDD.n3389 GND 0.011992f
C3882 VDD.n3390 GND 0.005441f
C3883 VDD.n3391 GND 0.005441f
C3884 VDD.n3392 GND 0.005441f
C3885 VDD.n3393 GND 0.005441f
C3886 VDD.n3394 GND 0.362306f
C3887 VDD.n3395 GND 0.005441f
C3888 VDD.n3396 GND 0.005441f
C3889 VDD.n3397 GND 0.005441f
C3890 VDD.n3398 GND 0.005441f
C3891 VDD.n3399 GND 0.005441f
C3892 VDD.n3400 GND 0.005441f
C3893 VDD.n3401 GND 0.005441f
C3894 VDD.n3403 GND 0.005441f
C3895 VDD.n3405 GND 0.005441f
C3896 VDD.n3406 GND 0.005441f
C3897 VDD.n3407 GND 0.005441f
C3898 VDD.n3408 GND 0.005441f
C3899 VDD.n3409 GND 0.005441f
C3900 VDD.n3410 GND 0.005441f
C3901 VDD.n3412 GND 0.005441f
C3902 VDD.n3413 GND 0.005441f
C3903 VDD.n3414 GND 0.005441f
C3904 VDD.n3415 GND 0.005441f
C3905 VDD.n3416 GND 0.005441f
C3906 VDD.n3417 GND 0.005441f
C3907 VDD.n3419 GND 0.005441f
C3908 VDD.n3420 GND 0.005441f
C3909 VDD.n3422 GND 0.013054f
C3910 VDD.n3423 GND 0.013054f
C3911 VDD.n3424 GND 0.011992f
C3912 VDD.n3425 GND 0.005441f
C3913 VDD.n3426 GND 0.005441f
C3914 VDD.n3427 GND 0.362306f
C3915 VDD.n3428 GND 0.005441f
C3916 VDD.n3429 GND 0.005441f
C3917 VDD.n3430 GND 0.012652f
C3918 VDD.n3431 GND 0.012394f
C3919 VDD.n3432 GND 0.013054f
C3920 VDD.n3434 GND 0.005441f
C3921 VDD.n3435 GND 0.005441f
C3922 VDD.n3436 GND 0.003321f
C3923 VDD.n3437 GND 0.005441f
C3924 VDD.n3438 GND 0.005441f
C3925 VDD.n3439 GND 0.005441f
C3926 VDD.n3441 GND 0.005441f
C3927 VDD.n3442 GND 0.005441f
C3928 VDD.n3443 GND 0.005441f
C3929 VDD.n3444 GND 0.005441f
C3930 VDD.n3445 GND 0.005441f
C3931 VDD.n3446 GND 0.005441f
C3932 VDD.n3448 GND 0.005441f
C3933 VDD.n3449 GND 0.005441f
C3934 VDD.n3450 GND 0.004081f
C3935 VDD.n3451 GND 0.027582f
C3936 VDD.n3452 GND 0.805083f
C3937 VDD.n3454 GND 0.008002f
C3938 VDD.t95 GND 0.029464f
C3939 VDD.t96 GND 0.049829f
C3940 VDD.t94 GND 0.498044f
C3941 VDD.n3455 GND 0.083391f
C3942 VDD.n3456 GND 0.066666f
C3943 VDD.n3458 GND 0.008002f
C3944 VDD.n3459 GND 0.00644f
C3945 VDD.n3460 GND 0.005346f
C3946 VDD.n3461 GND 0.007362f
C3947 VDD.n3462 GND 0.008002f
C3948 VDD.n3463 GND 0.00644f
C3949 VDD.n3465 GND 0.008002f
C3950 VDD.n3466 GND 0.008002f
C3951 VDD.n3468 GND 0.008002f
C3952 VDD.n3469 GND 0.00644f
C3953 VDD.n3471 GND 0.00644f
C3954 VDD.n3472 GND 0.00644f
C3955 VDD.n3473 GND 0.008002f
C3956 VDD.n3475 GND 0.008002f
C3957 VDD.n3476 GND 0.004347f
C3958 VDD.n3477 GND 0.013139f
C3959 VDD.n3478 GND 0.004641f
C3960 VDD.n3479 GND 0.008002f
C3961 VDD.n3480 GND 0.008002f
C3962 VDD.n3481 GND 0.00644f
C3963 VDD.n3482 GND 0.008002f
C3964 VDD.n3484 GND 0.008002f
C3965 VDD.n3486 GND 0.008002f
C3966 VDD.n3487 GND 0.00644f
C3967 VDD.n3488 GND 0.008002f
C3968 VDD.n3489 GND 0.008002f
C3969 VDD.n3490 GND 0.008002f
C3970 VDD.n3491 GND 0.00644f
C3971 VDD.n3492 GND 0.008002f
C3972 VDD.n3494 GND 0.008002f
C3973 VDD.n3496 GND 0.008002f
C3974 VDD.n3497 GND 0.005764f
C3975 VDD.n3498 GND 0.008002f
C3976 VDD.n3499 GND 0.008002f
C3977 VDD.n3500 GND 0.008002f
C3978 VDD.n3501 GND 0.004991f
C3979 VDD.n3502 GND 0.008002f
C3980 VDD.n3504 GND 0.008002f
C3981 VDD.n3506 GND 0.008002f
C3982 VDD.n3507 GND 0.00644f
C3983 VDD.n3508 GND 0.008002f
C3984 VDD.n3509 GND 0.008002f
C3985 VDD.n3510 GND 0.008002f
C3986 VDD.n3511 GND 0.00644f
C3987 VDD.n3512 GND 0.008002f
C3988 VDD.n3514 GND 0.008002f
C3989 VDD.n3516 GND 0.008002f
C3990 VDD.n3517 GND 0.00644f
C3991 VDD.n3518 GND 0.008002f
C3992 VDD.n3519 GND 0.008002f
C3993 VDD.n3520 GND 0.008002f
C3994 VDD.t104 GND 0.029464f
C3995 VDD.t105 GND 0.049829f
C3996 VDD.t103 GND 0.498044f
C3997 VDD.n3521 GND 0.083391f
C3998 VDD.n3522 GND 0.066666f
C3999 VDD.n3523 GND 0.009918f
C4000 VDD.n3524 GND 0.003961f
C4001 VDD.n3525 GND 0.008002f
C4002 VDD.n3527 GND 0.008002f
C4003 VDD.n3529 GND 0.008002f
C4004 VDD.n3530 GND 0.00644f
C4005 VDD.n3531 GND 0.008002f
C4006 VDD.n3532 GND 0.008002f
C4007 VDD.n3533 GND 0.008002f
C4008 VDD.n3534 GND 0.00644f
C4009 VDD.n3535 GND 0.008002f
C4010 VDD.n3537 GND 0.008002f
C4011 VDD.n3539 GND 0.008002f
C4012 VDD.n3540 GND 0.00644f
C4013 VDD.n3541 GND 0.008002f
C4014 VDD.n3542 GND 0.008002f
C4015 VDD.n3543 GND 0.008002f
C4016 VDD.n3544 GND 0.00644f
C4017 VDD.n3545 GND 0.008002f
C4018 VDD.n3547 GND 0.008002f
C4019 VDD.n3549 GND 0.008002f
C4020 VDD.t49 GND 0.029464f
C4021 VDD.t50 GND 0.049829f
C4022 VDD.t48 GND 0.498044f
C4023 VDD.n3550 GND 0.083391f
C4024 VDD.n3551 GND 0.066666f
C4025 VDD.n3552 GND 0.013139f
C4026 VDD.n3553 GND 0.008002f
C4027 VDD.n3554 GND 0.008002f
C4028 VDD.n3555 GND 0.008002f
C4029 VDD.n3556 GND 0.00644f
C4030 VDD.n3557 GND 0.008002f
C4031 VDD.n3559 GND 0.008002f
C4032 VDD.n3561 GND 0.008002f
C4033 VDD.n3562 GND 0.00644f
C4034 VDD.n3564 GND 0.805083f
C4035 VDD.n3566 GND 0.00644f
C4036 VDD.n3567 GND 0.008002f
C4037 VDD.n3569 GND 0.008002f
C4038 VDD.n3570 GND 0.008002f
C4039 VDD.n3572 GND 0.008002f
C4040 VDD.n3573 GND 0.003574f
C4041 VDD.n3574 GND 0.009918f
C4042 VDD.n3575 GND 0.002866f
C4043 VDD.n3576 GND 0.01975f
C4044 VDD.n3577 GND 0.019459f
C4045 VDD.n3578 GND 0.005346f
C4046 VDD.n3579 GND 0.019459f
C4047 VDD.n3580 GND 0.772565f
C4048 VDD.n3581 GND 0.019459f
C4049 VDD.n3582 GND 0.005346f
C4050 VDD.n3583 GND 0.019459f
C4051 VDD.n3584 GND 0.008002f
C4052 VDD.n3585 GND 0.008002f
C4053 VDD.n3586 GND 0.00644f
C4054 VDD.n3587 GND 0.008002f
C4055 VDD.n3588 GND 0.532804f
C4056 VDD.n3589 GND 0.008002f
C4057 VDD.n3590 GND 0.00644f
C4058 VDD.n3591 GND 0.008002f
C4059 VDD.n3592 GND 0.008002f
C4060 VDD.n3593 GND 0.008002f
C4061 VDD.n3594 GND 0.00644f
C4062 VDD.n3595 GND 0.008002f
C4063 VDD.n3596 GND 0.418251f
C4064 VDD.n3597 GND 0.532804f
C4065 VDD.n3598 GND 0.008002f
C4066 VDD.n3599 GND 0.00644f
C4067 VDD.n3600 GND 0.008002f
C4068 VDD.n3601 GND 0.008002f
C4069 VDD.n3602 GND 0.008002f
C4070 VDD.n3603 GND 0.00644f
C4071 VDD.n3604 GND 0.008002f
C4072 VDD.n3605 GND 0.380955f
C4073 VDD.n3606 GND 0.008002f
C4074 VDD.n3607 GND 0.00644f
C4075 VDD.n3608 GND 0.008002f
C4076 VDD.n3609 GND 0.008002f
C4077 VDD.n3610 GND 0.008002f
C4078 VDD.n3611 GND 0.00644f
C4079 VDD.n3612 GND 0.008002f
C4080 VDD.n3613 GND 0.532804f
C4081 VDD.n3614 GND 0.008002f
C4082 VDD.n3615 GND 0.00644f
C4083 VDD.n3616 GND 0.008002f
C4084 VDD.n3617 GND 0.008002f
C4085 VDD.n3618 GND 0.008002f
C4086 VDD.n3619 GND 0.00644f
C4087 VDD.n3620 GND 0.008002f
C4088 VDD.n3621 GND 0.532804f
C4089 VDD.n3622 GND 0.008002f
C4090 VDD.n3623 GND 0.00644f
C4091 VDD.n3624 GND 0.008002f
C4092 VDD.n3625 GND 0.008002f
C4093 VDD.n3626 GND 0.008002f
C4094 VDD.n3627 GND 0.00644f
C4095 VDD.n3628 GND 0.008002f
C4096 VDD.n3629 GND 0.532804f
C4097 VDD.n3630 GND 0.008002f
C4098 VDD.n3631 GND 0.00644f
C4099 VDD.n3632 GND 0.008002f
C4100 VDD.n3633 GND 0.008002f
C4101 VDD.n3634 GND 0.008002f
C4102 VDD.n3635 GND 0.00644f
C4103 VDD.n3636 GND 0.008002f
C4104 VDD.n3637 GND 0.532804f
C4105 VDD.n3638 GND 0.008002f
C4106 VDD.n3639 GND 0.00644f
C4107 VDD.n3640 GND 0.008002f
C4108 VDD.n3641 GND 0.008002f
C4109 VDD.n3642 GND 0.008002f
C4110 VDD.n3643 GND 0.00644f
C4111 VDD.n3644 GND 0.008002f
C4112 VDD.n3645 GND 0.532804f
C4113 VDD.n3646 GND 0.008002f
C4114 VDD.n3647 GND 0.00644f
C4115 VDD.n3648 GND 0.008002f
C4116 VDD.n3649 GND 0.008002f
C4117 VDD.n3650 GND 0.008002f
C4118 VDD.n3651 GND 0.00644f
C4119 VDD.n3652 GND 0.008002f
C4120 VDD.n3653 GND 0.492843f
C4121 VDD.n3654 GND 0.008002f
C4122 VDD.n3655 GND 0.00644f
C4123 VDD.n3656 GND 0.008002f
C4124 VDD.n3657 GND 0.008002f
C4125 VDD.n3658 GND 0.008002f
C4126 VDD.n3659 GND 0.00644f
C4127 VDD.n3660 GND 0.008002f
C4128 VDD.n3661 GND 0.532804f
C4129 VDD.n3662 GND 0.008002f
C4130 VDD.n3663 GND 0.00644f
C4131 VDD.n3664 GND 0.008002f
C4132 VDD.n3665 GND 0.008002f
C4133 VDD.n3666 GND 0.008002f
C4134 VDD.n3667 GND 0.00644f
C4135 VDD.n3668 GND 0.008002f
C4136 VDD.n3669 GND 0.532804f
C4137 VDD.n3670 GND 0.008002f
C4138 VDD.n3671 GND 0.00644f
C4139 VDD.n3672 GND 0.008002f
C4140 VDD.n3673 GND 0.008002f
C4141 VDD.n3674 GND 0.008002f
C4142 VDD.n3675 GND 0.00644f
C4143 VDD.n3676 GND 0.008002f
C4144 VDD.n3677 GND 0.532804f
C4145 VDD.n3678 GND 0.008002f
C4146 VDD.n3679 GND 0.00644f
C4147 VDD.n3680 GND 0.008002f
C4148 VDD.n3681 GND 0.008002f
C4149 VDD.n3682 GND 0.008002f
C4150 VDD.n3683 GND 0.00644f
C4151 VDD.n3684 GND 0.008002f
C4152 VDD.n3685 GND 0.532804f
C4153 VDD.n3686 GND 0.008002f
C4154 VDD.n3687 GND 0.00644f
C4155 VDD.n3688 GND 0.008002f
C4156 VDD.n3689 GND 0.008002f
C4157 VDD.n3690 GND 0.008002f
C4158 VDD.n3691 GND 0.00644f
C4159 VDD.n3692 GND 0.008002f
C4160 VDD.n3693 GND 0.519484f
C4161 VDD.n3694 GND 0.532804f
C4162 VDD.n3695 GND 0.008002f
C4163 VDD.n3696 GND 0.00644f
C4164 VDD.n3697 GND 0.008002f
C4165 VDD.n3698 GND 0.008002f
C4166 VDD.n3699 GND 0.008002f
C4167 VDD.n3700 GND 0.00644f
C4168 VDD.n3701 GND 0.008002f
C4169 VDD.n3702 GND 0.279722f
C4170 VDD.n3703 GND 0.008002f
C4171 VDD.n3704 GND 0.00644f
C4172 VDD.n3705 GND 0.008002f
C4173 VDD.n3706 GND 0.008002f
C4174 VDD.n3707 GND 0.008002f
C4175 VDD.n3708 GND 0.008002f
C4176 VDD.n3709 GND 0.008002f
C4177 VDD.n3710 GND 0.00644f
C4178 VDD.n3711 GND 0.00644f
C4179 VDD.n3712 GND 0.008002f
C4180 VDD.n3713 GND 0.532804f
C4181 VDD.n3714 GND 0.008002f
C4182 VDD.n3715 GND 0.00644f
C4183 VDD.n3716 GND 0.008002f
C4184 VDD.n3717 GND 0.008002f
C4185 VDD.n3718 GND 0.008002f
C4186 VDD.n3719 GND 0.00644f
C4187 VDD.n3720 GND 0.008002f
C4188 VDD.n3721 GND 0.532804f
C4189 VDD.n3722 GND 0.008002f
C4190 VDD.n3723 GND 0.008002f
C4191 VDD.n3724 GND 0.00644f
C4192 VDD.n3725 GND 0.00644f
C4193 VDD.n3726 GND 0.00644f
C4194 VDD.n3727 GND 0.008002f
C4195 VDD.n3728 GND 0.008002f
C4196 VDD.n3729 GND 0.008002f
C4197 VDD.n3730 GND 0.008002f
C4198 VDD.n3731 GND 0.00644f
C4199 VDD.n3732 GND 0.00644f
C4200 VDD.n3733 GND 0.00644f
C4201 VDD.n3734 GND 0.008002f
C4202 VDD.n3735 GND 0.008002f
C4203 VDD.n3736 GND 0.008002f
C4204 VDD.n3737 GND 0.008002f
C4205 VDD.n3738 GND 0.00644f
C4206 VDD.n3739 GND 0.00644f
C4207 VDD.n3740 GND 0.00644f
C4208 VDD.n3741 GND 0.008002f
C4209 VDD.n3742 GND 0.008002f
C4210 VDD.n3743 GND 0.008002f
C4211 VDD.n3744 GND 0.008002f
C4212 VDD.n3745 GND 0.00644f
C4213 VDD.n3746 GND 0.00644f
C4214 VDD.n3747 GND 0.00644f
C4215 VDD.n3748 GND 0.008002f
C4216 VDD.n3749 GND 0.008002f
C4217 VDD.n3750 GND 0.008002f
C4218 VDD.n3751 GND 0.008002f
C4219 VDD.n3752 GND 0.00644f
C4220 VDD.n3753 GND 0.00644f
C4221 VDD.n3754 GND 0.00644f
C4222 VDD.n3755 GND 0.008002f
C4223 VDD.n3756 GND 0.008002f
C4224 VDD.n3757 GND 0.008002f
C4225 VDD.n3758 GND 0.008002f
C4226 VDD.n3759 GND 0.00644f
C4227 VDD.n3760 GND 0.00644f
C4228 VDD.n3761 GND 0.00644f
C4229 VDD.n3762 GND 0.008002f
C4230 VDD.n3763 GND 0.008002f
C4231 VDD.n3764 GND 0.008002f
C4232 VDD.n3765 GND 0.008002f
C4233 VDD.n3766 GND 0.00644f
C4234 VDD.n3767 GND 0.00644f
C4235 VDD.n3768 GND 0.00644f
C4236 VDD.n3769 GND 0.008002f
C4237 VDD.n3770 GND 0.008002f
C4238 VDD.n3771 GND 0.008002f
C4239 VDD.n3772 GND 0.008002f
C4240 VDD.n3773 GND 0.00644f
C4241 VDD.n3774 GND 0.00644f
C4242 VDD.n3775 GND 0.00644f
C4243 VDD.n3776 GND 0.008002f
C4244 VDD.n3777 GND 0.008002f
C4245 VDD.n3778 GND 0.008002f
C4246 VDD.n3779 GND 0.008002f
C4247 VDD.n3780 GND 0.00644f
C4248 VDD.n3781 GND 0.00644f
C4249 VDD.n3782 GND 0.00644f
C4250 VDD.n3783 GND 0.008002f
C4251 VDD.n3784 GND 0.008002f
C4252 VDD.n3785 GND 0.019459f
C4253 VDD.n3786 GND 0.005346f
C4254 VDD.n3787 GND 0.019459f
C4255 VDD.n3788 GND 0.01975f
C4256 VDD.n3789 GND 0.002866f
C4257 VDD.t40 GND 0.029464f
C4258 VDD.t39 GND 0.049829f
C4259 VDD.t37 GND 0.498044f
C4260 VDD.n3790 GND 0.083391f
C4261 VDD.n3791 GND 0.066666f
C4262 VDD.n3792 GND 0.009918f
C4263 VDD.n3793 GND 0.003574f
C4264 VDD.n3794 GND 0.00644f
C4265 VDD.n3795 GND 0.008002f
C4266 VDD.n3797 GND 0.008002f
C4267 VDD.n3798 GND 0.008002f
C4268 VDD.n3799 GND 0.00644f
C4269 VDD.n3800 GND 0.00644f
C4270 VDD.n3801 GND 0.00644f
C4271 VDD.n3802 GND 0.008002f
C4272 VDD.n3804 GND 0.008002f
C4273 VDD.n3805 GND 0.008002f
C4274 VDD.n3806 GND 0.00644f
C4275 VDD.n3807 GND 0.008002f
C4276 VDD.n3808 GND 0.008002f
C4277 VDD.n3809 GND 0.008002f
C4278 VDD.n3810 GND 0.013139f
C4279 VDD.n3811 GND 0.005378f
C4280 VDD.n3812 GND 0.00644f
C4281 VDD.n3813 GND 0.008002f
C4282 VDD.n3815 GND 0.008002f
C4283 VDD.n3816 GND 0.008002f
C4284 VDD.n3817 GND 0.00644f
C4285 VDD.n3818 GND 0.00644f
C4286 VDD.n3819 GND 0.00644f
C4287 VDD.n3820 GND 0.008002f
C4288 VDD.n3822 GND 0.008002f
C4289 VDD.n3823 GND 0.008002f
C4290 VDD.n3824 GND 0.00644f
C4291 VDD.n3825 GND 0.003574f
C4292 VDD.t60 GND 0.029464f
C4293 VDD.t59 GND 0.049829f
C4294 VDD.t58 GND 0.498044f
C4295 VDD.n3826 GND 0.083391f
C4296 VDD.n3827 GND 0.066666f
C4297 VDD.n3828 GND 0.009918f
C4298 VDD.n3829 GND 0.003961f
C4299 VDD.n3830 GND 0.008002f
C4300 VDD.n3832 GND 0.008002f
C4301 VDD.n3833 GND 0.008002f
C4302 VDD.n3834 GND 0.00644f
C4303 VDD.n3835 GND 0.00644f
C4304 VDD.n3836 GND 0.00644f
C4305 VDD.n3837 GND 0.008002f
C4306 VDD.n3839 GND 0.008002f
C4307 VDD.n3840 GND 0.008002f
C4308 VDD.n3842 GND 0.008002f
C4309 VDD.n3843 GND 0.00644f
C4310 VDD.n3844 GND 0.008002f
C4311 VDD.n3845 GND 0.008002f
C4312 VDD.n3846 GND 0.008002f
C4313 VDD.n3847 GND 0.013139f
C4314 VDD.n3848 GND 0.005764f
C4315 VDD.n3849 GND 0.008002f
C4316 VDD.n3851 GND 0.008002f
C4317 VDD.n3852 GND 0.008002f
C4318 VDD.n3853 GND 0.00644f
C4319 VDD.n3854 GND 0.00644f
C4320 VDD.n3855 GND 0.00644f
C4321 VDD.n3856 GND 0.008002f
C4322 VDD.n3858 GND 0.008002f
C4323 VDD.n3859 GND 0.008002f
C4324 VDD.n3860 GND 0.00644f
C4325 VDD.n3861 GND 0.008002f
C4326 VDD.n3862 GND 0.008002f
C4327 VDD.n3863 GND 0.008002f
C4328 VDD.n3864 GND 0.013139f
C4329 VDD.n3865 GND 0.008002f
C4330 VDD.n3867 GND 0.008002f
C4331 VDD.n3868 GND 0.008002f
C4332 VDD.n3869 GND 0.00644f
C4333 VDD.n3870 GND 0.00644f
C4334 VDD.n3871 GND 0.00644f
C4335 VDD.n3872 GND 0.008002f
C4336 VDD.n3874 GND 0.008002f
C4337 VDD.n3875 GND 0.008002f
C4338 VDD.n3877 GND 0.01975f
C4339 VDD.n3878 GND 0.005346f
C4340 VDD.n3879 GND 0.01975f
C4341 VDD.n3880 GND 0.019459f
C4342 VDD.n3881 GND 0.005346f
C4343 VDD.n3882 GND 0.00644f
C4344 VDD.n3883 GND 0.008002f
C4345 VDD.n3884 GND 0.532804f
C4346 VDD.n3885 GND 0.532804f
C4347 VDD.n3886 GND 0.532804f
C4348 VDD.n3887 GND 0.008002f
C4349 VDD.n3888 GND 0.00644f
C4350 VDD.n3889 GND 0.00644f
C4351 VDD.n3890 GND 0.00644f
C4352 VDD.n3891 GND 0.008002f
C4353 VDD.n3892 GND 0.418251f
C4354 VDD.t38 GND 0.266402f
C4355 VDD.n3893 GND 0.380955f
C4356 VDD.n3894 GND 0.532804f
C4357 VDD.n3895 GND 0.008002f
C4358 VDD.n3896 GND 0.00644f
C4359 VDD.n3897 GND 0.00644f
C4360 VDD.n3898 GND 0.00644f
C4361 VDD.n3899 GND 0.008002f
C4362 VDD.n3900 GND 0.532804f
C4363 VDD.n3901 GND 0.532804f
C4364 VDD.n3902 GND 0.532804f
C4365 VDD.n3903 GND 0.008002f
C4366 VDD.n3904 GND 0.00644f
C4367 VDD.n3905 GND 0.00644f
C4368 VDD.n3906 GND 0.00644f
C4369 VDD.n3907 GND 0.008002f
C4370 VDD.n3908 GND 0.532804f
C4371 VDD.n3909 GND 0.532804f
C4372 VDD.n3910 GND 0.532804f
C4373 VDD.n3911 GND 0.008002f
C4374 VDD.n3912 GND 0.00644f
C4375 VDD.n3913 GND 0.00644f
C4376 VDD.n3914 GND 0.00644f
C4377 VDD.n3915 GND 0.008002f
C4378 VDD.n3916 GND 0.532804f
C4379 VDD.n3917 GND 0.492843f
C4380 VDD.t141 GND 0.266402f
C4381 VDD.n3918 GND 0.306362f
C4382 VDD.n3919 GND 0.008002f
C4383 VDD.n3920 GND 0.00644f
C4384 VDD.n3921 GND 0.00644f
C4385 VDD.n3922 GND 0.00644f
C4386 VDD.n3923 GND 0.008002f
C4387 VDD.n3924 GND 0.532804f
C4388 VDD.n3925 GND 0.532804f
C4389 VDD.n3926 GND 0.532804f
C4390 VDD.n3927 GND 0.008002f
C4391 VDD.n3928 GND 0.00644f
C4392 VDD.n3929 GND 0.00644f
C4393 VDD.n3930 GND 0.00644f
C4394 VDD.n3931 GND 0.008002f
C4395 VDD.n3932 GND 0.532804f
C4396 VDD.n3933 GND 0.532804f
C4397 VDD.n3934 GND 0.532804f
C4398 VDD.n3935 GND 0.008002f
C4399 VDD.n3936 GND 0.00644f
C4400 VDD.n3937 GND 0.00644f
C4401 VDD.n3938 GND 0.00644f
C4402 VDD.n3939 GND 0.008002f
C4403 VDD.n3940 GND 0.519484f
C4404 VDD.t138 GND 0.266402f
C4405 VDD.n3941 GND 0.279722f
C4406 VDD.n3942 GND 0.532804f
C4407 VDD.n3943 GND 0.008002f
C4408 VDD.n3944 GND 0.00644f
C4409 VDD.n3945 GND 0.00644f
C4410 VDD.n3946 GND 0.00644f
C4411 VDD.n3947 GND 0.008002f
C4412 VDD.n3948 GND 0.532804f
C4413 VDD.n3949 GND 0.532804f
C4414 VDD.n3950 GND 0.532804f
C4415 VDD.n3951 GND 0.008002f
C4416 VDD.n3952 GND 0.00644f
C4417 VDD.n3953 GND 0.00615f
C4418 VDD.n3954 GND 0.232322f
C4419 VDD.n3955 GND 2.75555f
C4420 VOUT.t10 GND 0.014762f
C4421 VOUT.t34 GND 0.014762f
C4422 VOUT.n0 GND 0.081709f
C4423 VOUT.t20 GND 0.014762f
C4424 VOUT.t41 GND 0.014762f
C4425 VOUT.n1 GND 0.071797f
C4426 VOUT.n2 GND 0.675338f
C4427 VOUT.t35 GND 0.014762f
C4428 VOUT.t37 GND 0.014762f
C4429 VOUT.n3 GND 0.081709f
C4430 VOUT.t23 GND 0.014762f
C4431 VOUT.t27 GND 0.014762f
C4432 VOUT.n4 GND 0.071797f
C4433 VOUT.n5 GND 0.655627f
C4434 VOUT.n6 GND 0.220762f
C4435 VOUT.t38 GND 0.014762f
C4436 VOUT.t31 GND 0.014762f
C4437 VOUT.n7 GND 0.081709f
C4438 VOUT.t15 GND 0.014762f
C4439 VOUT.t40 GND 0.014762f
C4440 VOUT.n8 GND 0.071797f
C4441 VOUT.n9 GND 0.655627f
C4442 VOUT.n10 GND 0.142952f
C4443 VOUT.t13 GND 0.014762f
C4444 VOUT.t36 GND 0.014762f
C4445 VOUT.n11 GND 0.081709f
C4446 VOUT.t12 GND 0.014762f
C4447 VOUT.t32 GND 0.014762f
C4448 VOUT.n12 GND 0.071797f
C4449 VOUT.n13 GND 0.655627f
C4450 VOUT.n14 GND 0.142952f
C4451 VOUT.t16 GND 0.014762f
C4452 VOUT.t6 GND 0.014762f
C4453 VOUT.n15 GND 0.081709f
C4454 VOUT.t25 GND 0.014762f
C4455 VOUT.t21 GND 0.014762f
C4456 VOUT.n16 GND 0.071797f
C4457 VOUT.n17 GND 0.655627f
C4458 VOUT.n18 GND 0.291818f
C4459 VOUT.n19 GND 10.0367f
C4460 VOUT.n20 GND 3.90827f
C4461 VOUT.t52 GND 5.47823f
C4462 VOUT.t49 GND 5.50791f
C4463 VOUT.t53 GND 5.50791f
C4464 VOUT.t50 GND 5.47823f
C4465 VOUT.n21 GND 4.77574f
C4466 VOUT.n22 GND 4.64154f
C4467 VOUT.t48 GND 5.47823f
C4468 VOUT.n23 GND 2.16601f
C4469 VOUT.t51 GND 5.50791f
C4470 VOUT.n24 GND 1.81765f
C4471 VOUT.n25 GND 4.56518f
C4472 VOUT.n26 GND 4.64154f
C4473 VOUT.n27 GND 2.16601f
C4474 VOUT.n28 GND 5.40835f
C4475 VOUT.n29 GND 2.14691f
C4476 VOUT.t5 GND 0.014762f
C4477 VOUT.t42 GND 0.014762f
C4478 VOUT.n30 GND 0.081709f
C4479 VOUT.t19 GND 0.014762f
C4480 VOUT.t7 GND 0.014762f
C4481 VOUT.n31 GND 0.071797f
C4482 VOUT.n32 GND 0.675338f
C4483 VOUT.t26 GND 0.014762f
C4484 VOUT.t8 GND 0.014762f
C4485 VOUT.n33 GND 0.081709f
C4486 VOUT.t22 GND 0.014762f
C4487 VOUT.t17 GND 0.014762f
C4488 VOUT.n34 GND 0.071797f
C4489 VOUT.n35 GND 0.655627f
C4490 VOUT.n36 GND 0.220762f
C4491 VOUT.t39 GND 0.014762f
C4492 VOUT.t11 GND 0.014762f
C4493 VOUT.n37 GND 0.081709f
C4494 VOUT.t43 GND 0.014762f
C4495 VOUT.t4 GND 0.014762f
C4496 VOUT.n38 GND 0.071797f
C4497 VOUT.n39 GND 0.655627f
C4498 VOUT.n40 GND 0.142952f
C4499 VOUT.t14 GND 0.014762f
C4500 VOUT.t29 GND 0.014762f
C4501 VOUT.n41 GND 0.081709f
C4502 VOUT.t30 GND 0.014762f
C4503 VOUT.t28 GND 0.014762f
C4504 VOUT.n42 GND 0.071797f
C4505 VOUT.n43 GND 0.655627f
C4506 VOUT.n44 GND 0.142952f
C4507 VOUT.t18 GND 0.014762f
C4508 VOUT.t9 GND 0.014762f
C4509 VOUT.n45 GND 0.081709f
C4510 VOUT.t33 GND 0.014762f
C4511 VOUT.t24 GND 0.014762f
C4512 VOUT.n46 GND 0.071797f
C4513 VOUT.n47 GND 0.655628f
C4514 VOUT.n48 GND 0.291818f
C4515 VOUT.n49 GND 13.753901f
C4516 VOUT.t45 GND 0.273165f
C4517 VOUT.t47 GND 0.2653f
C4518 VOUT.n50 GND 0.549443f
C4519 VOUT.t0 GND 0.2653f
C4520 VOUT.n51 GND 0.310478f
C4521 VOUT.t3 GND 0.2653f
C4522 VOUT.n52 GND 0.428665f
C4523 VOUT.n53 GND 11.526f
C4524 VOUT.t1 GND 0.27217f
C4525 VOUT.t2 GND 0.264173f
C4526 VOUT.n54 GND 0.551565f
C4527 VOUT.t44 GND 0.264173f
C4528 VOUT.n55 GND 0.311604f
C4529 VOUT.t46 GND 0.264173f
C4530 VOUT.n56 GND 0.429792f
C4531 VOUT.n57 GND 8.18925f
C4532 VOUT.n58 GND 7.17279f
C4533 a_n14320_7092.t1 GND 0.466615f
C4534 a_n14320_7092.t3 GND 0.48118f
C4535 a_n14320_7092.t2 GND 0.466615f
C4536 a_n14320_7092.t0 GND 0.466616f
C4537 a_n14320_7092.n0 GND 0.765191f
C4538 a_n14320_7092.n1 GND 8.42933f
C4539 a_n14320_7092.n2 GND 0.765191f
C4540 a_n14320_7092.n3 GND 0.765191f
C4541 a_n14320_7092.n4 GND 11.7635f
C4542 a_n14320_7092.n5 GND 3.06192f
C4543 a_n14320_7092.n6 GND 2.01559f
C4544 a_n14320_7092.n7 GND 0.756636f
C4545 a_n14320_7092.n8 GND 0.756636f
C4546 a_n14320_7092.n9 GND 0.756636f
C4547 a_n14320_7092.n10 GND 0.756636f
C4548 a_n14320_7092.n11 GND 3.09638f
C4549 a_n14320_7092.n12 GND 0.756636f
C4550 a_n14320_7092.n13 GND 20.634f
C4551 a_n14320_7092.n14 GND 2.95842f
C4552 a_n14320_7092.n15 GND 2.40563f
C4553 a_n14320_7092.n16 GND 0.765191f
C4554 a_n14320_7092.n17 GND 1.03323f
C4555 a_n14320_7092.n18 GND 1.03323f
C4556 a_n14320_7092.n19 GND 1.03323f
C4557 a_n14320_7092.n20 GND 1.03323f
C4558 a_n14320_7092.n21 GND 0.765191f
C4559 a_n14320_7092.n22 GND 2.05005f
C4560 a_n14320_7092.n23 GND 1.03323f
C4561 a_n14320_7092.t6 GND 0.491821f
C4562 a_n14320_7092.t5 GND 0.481216f
C4563 a_n14320_7092.t4 GND 0.279165f
C4564 a_n14320_7092.t7 GND 0.482019f
C4565 a_n14320_7092.n24 GND 1.92126f
C4566 a_n14320_7092.t45 GND 1.67229f
C4567 a_n14320_7092.t33 GND 1.6417f
C4568 a_n14320_7092.t20 GND 1.67751f
C4569 a_n14320_7092.t46 GND 1.68439f
C4570 a_n14320_7092.t27 GND 1.67229f
C4571 a_n14320_7092.t18 GND 1.6417f
C4572 a_n14320_7092.t43 GND 1.67751f
C4573 a_n14320_7092.t28 GND 1.68439f
C4574 a_n14320_7092.t44 GND 1.67229f
C4575 a_n14320_7092.t25 GND 1.6417f
C4576 a_n14320_7092.t41 GND 1.67751f
C4577 a_n14320_7092.t16 GND 1.68439f
C4578 a_n14320_7092.t26 GND 1.67229f
C4579 a_n14320_7092.t10 GND 1.6417f
C4580 a_n14320_7092.t23 GND 1.67751f
C4581 a_n14320_7092.t39 GND 1.68439f
C4582 a_n14320_7092.t11 GND 1.67229f
C4583 a_n14320_7092.t30 GND 1.6417f
C4584 a_n14320_7092.t47 GND 1.67751f
C4585 a_n14320_7092.t21 GND 1.68439f
C4586 a_n14320_7092.t31 GND 1.67845f
C4587 a_n14320_7092.t13 GND 1.64076f
C4588 a_n14320_7092.t12 GND 1.63961f
C4589 a_n14320_7092.t38 GND 1.7216f
C4590 a_n14320_7092.t17 GND 1.67845f
C4591 a_n14320_7092.t37 GND 1.64076f
C4592 a_n14320_7092.t36 GND 1.63961f
C4593 a_n14320_7092.t22 GND 1.7216f
C4594 a_n14320_7092.t42 GND 1.67845f
C4595 a_n14320_7092.t29 GND 1.64076f
C4596 a_n14320_7092.t34 GND 1.63961f
C4597 a_n14320_7092.t9 GND 1.7216f
C4598 a_n14320_7092.t24 GND 1.67845f
C4599 a_n14320_7092.t14 GND 1.64076f
C4600 a_n14320_7092.t19 GND 1.63961f
C4601 a_n14320_7092.t32 GND 1.7216f
C4602 a_n14320_7092.t8 GND 1.67845f
C4603 a_n14320_7092.t35 GND 1.64076f
C4604 a_n14320_7092.t40 GND 1.63961f
C4605 a_n14320_7092.t15 GND 1.7216f
C4606 a_n14320_7092.n25 GND 3.49186f
.ends

