* NGSPICE file created from diff_pair_sample_1321.ext - technology: sky130A

.subckt diff_pair_sample_1321 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t7 VN.t0 VTAIL.t9 w_n4100_n1956# sky130_fd_pr__pfet_01v8 ad=0.8151 pd=5.27 as=0.8151 ps=5.27 w=4.94 l=2.8
X1 B.t11 B.t9 B.t10 w_n4100_n1956# sky130_fd_pr__pfet_01v8 ad=1.9266 pd=10.66 as=0 ps=0 w=4.94 l=2.8
X2 VTAIL.t14 VN.t1 VDD2.t6 w_n4100_n1956# sky130_fd_pr__pfet_01v8 ad=0.8151 pd=5.27 as=0.8151 ps=5.27 w=4.94 l=2.8
X3 VDD1.t7 VP.t0 VTAIL.t1 w_n4100_n1956# sky130_fd_pr__pfet_01v8 ad=0.8151 pd=5.27 as=0.8151 ps=5.27 w=4.94 l=2.8
X4 VTAIL.t11 VN.t2 VDD2.t5 w_n4100_n1956# sky130_fd_pr__pfet_01v8 ad=1.9266 pd=10.66 as=0.8151 ps=5.27 w=4.94 l=2.8
X5 VTAIL.t15 VN.t3 VDD2.t4 w_n4100_n1956# sky130_fd_pr__pfet_01v8 ad=0.8151 pd=5.27 as=0.8151 ps=5.27 w=4.94 l=2.8
X6 VDD2.t3 VN.t4 VTAIL.t13 w_n4100_n1956# sky130_fd_pr__pfet_01v8 ad=0.8151 pd=5.27 as=1.9266 ps=10.66 w=4.94 l=2.8
X7 VDD2.t2 VN.t5 VTAIL.t12 w_n4100_n1956# sky130_fd_pr__pfet_01v8 ad=0.8151 pd=5.27 as=1.9266 ps=10.66 w=4.94 l=2.8
X8 VDD2.t1 VN.t6 VTAIL.t10 w_n4100_n1956# sky130_fd_pr__pfet_01v8 ad=0.8151 pd=5.27 as=0.8151 ps=5.27 w=4.94 l=2.8
X9 VDD1.t6 VP.t1 VTAIL.t2 w_n4100_n1956# sky130_fd_pr__pfet_01v8 ad=0.8151 pd=5.27 as=1.9266 ps=10.66 w=4.94 l=2.8
X10 B.t8 B.t6 B.t7 w_n4100_n1956# sky130_fd_pr__pfet_01v8 ad=1.9266 pd=10.66 as=0 ps=0 w=4.94 l=2.8
X11 VDD1.t5 VP.t2 VTAIL.t3 w_n4100_n1956# sky130_fd_pr__pfet_01v8 ad=0.8151 pd=5.27 as=0.8151 ps=5.27 w=4.94 l=2.8
X12 VTAIL.t4 VP.t3 VDD1.t4 w_n4100_n1956# sky130_fd_pr__pfet_01v8 ad=1.9266 pd=10.66 as=0.8151 ps=5.27 w=4.94 l=2.8
X13 VDD1.t3 VP.t4 VTAIL.t5 w_n4100_n1956# sky130_fd_pr__pfet_01v8 ad=0.8151 pd=5.27 as=1.9266 ps=10.66 w=4.94 l=2.8
X14 VTAIL.t6 VP.t5 VDD1.t2 w_n4100_n1956# sky130_fd_pr__pfet_01v8 ad=1.9266 pd=10.66 as=0.8151 ps=5.27 w=4.94 l=2.8
X15 B.t5 B.t3 B.t4 w_n4100_n1956# sky130_fd_pr__pfet_01v8 ad=1.9266 pd=10.66 as=0 ps=0 w=4.94 l=2.8
X16 VTAIL.t8 VN.t7 VDD2.t0 w_n4100_n1956# sky130_fd_pr__pfet_01v8 ad=1.9266 pd=10.66 as=0.8151 ps=5.27 w=4.94 l=2.8
X17 VTAIL.t0 VP.t6 VDD1.t1 w_n4100_n1956# sky130_fd_pr__pfet_01v8 ad=0.8151 pd=5.27 as=0.8151 ps=5.27 w=4.94 l=2.8
X18 B.t2 B.t0 B.t1 w_n4100_n1956# sky130_fd_pr__pfet_01v8 ad=1.9266 pd=10.66 as=0 ps=0 w=4.94 l=2.8
X19 VTAIL.t7 VP.t7 VDD1.t0 w_n4100_n1956# sky130_fd_pr__pfet_01v8 ad=0.8151 pd=5.27 as=0.8151 ps=5.27 w=4.94 l=2.8
R0 VN.n56 VN.n55 161.3
R1 VN.n54 VN.n30 161.3
R2 VN.n53 VN.n52 161.3
R3 VN.n51 VN.n31 161.3
R4 VN.n50 VN.n49 161.3
R5 VN.n48 VN.n32 161.3
R6 VN.n46 VN.n45 161.3
R7 VN.n44 VN.n33 161.3
R8 VN.n43 VN.n42 161.3
R9 VN.n41 VN.n34 161.3
R10 VN.n40 VN.n39 161.3
R11 VN.n38 VN.n35 161.3
R12 VN.n27 VN.n26 161.3
R13 VN.n25 VN.n1 161.3
R14 VN.n24 VN.n23 161.3
R15 VN.n22 VN.n2 161.3
R16 VN.n21 VN.n20 161.3
R17 VN.n19 VN.n3 161.3
R18 VN.n17 VN.n16 161.3
R19 VN.n15 VN.n4 161.3
R20 VN.n14 VN.n13 161.3
R21 VN.n12 VN.n5 161.3
R22 VN.n11 VN.n10 161.3
R23 VN.n9 VN.n6 161.3
R24 VN.n37 VN.t4 74.4816
R25 VN.n8 VN.t2 74.4816
R26 VN.n28 VN.n0 68.3588
R27 VN.n57 VN.n29 68.3588
R28 VN.n8 VN.n7 58.3801
R29 VN.n37 VN.n36 58.3801
R30 VN.n13 VN.n12 56.5617
R31 VN.n42 VN.n41 56.5617
R32 VN.n24 VN.n2 52.2023
R33 VN.n53 VN.n31 52.2023
R34 VN VN.n57 46.7481
R35 VN.n7 VN.t6 42.5198
R36 VN.n18 VN.t3 42.5198
R37 VN.n0 VN.t5 42.5198
R38 VN.n36 VN.t1 42.5198
R39 VN.n47 VN.t0 42.5198
R40 VN.n29 VN.t7 42.5198
R41 VN.n25 VN.n24 28.9518
R42 VN.n54 VN.n53 28.9518
R43 VN.n11 VN.n6 24.5923
R44 VN.n12 VN.n11 24.5923
R45 VN.n13 VN.n4 24.5923
R46 VN.n17 VN.n4 24.5923
R47 VN.n20 VN.n19 24.5923
R48 VN.n20 VN.n2 24.5923
R49 VN.n26 VN.n25 24.5923
R50 VN.n41 VN.n40 24.5923
R51 VN.n40 VN.n35 24.5923
R52 VN.n49 VN.n31 24.5923
R53 VN.n49 VN.n48 24.5923
R54 VN.n46 VN.n33 24.5923
R55 VN.n42 VN.n33 24.5923
R56 VN.n55 VN.n54 24.5923
R57 VN.n26 VN.n0 21.8872
R58 VN.n55 VN.n29 21.8872
R59 VN.n7 VN.n6 15.4934
R60 VN.n18 VN.n17 15.4934
R61 VN.n36 VN.n35 15.4934
R62 VN.n47 VN.n46 15.4934
R63 VN.n19 VN.n18 9.09948
R64 VN.n48 VN.n47 9.09948
R65 VN.n38 VN.n37 5.39044
R66 VN.n9 VN.n8 5.39044
R67 VN.n57 VN.n56 0.354861
R68 VN.n28 VN.n27 0.354861
R69 VN VN.n28 0.267071
R70 VN.n56 VN.n30 0.189894
R71 VN.n52 VN.n30 0.189894
R72 VN.n52 VN.n51 0.189894
R73 VN.n51 VN.n50 0.189894
R74 VN.n50 VN.n32 0.189894
R75 VN.n45 VN.n32 0.189894
R76 VN.n45 VN.n44 0.189894
R77 VN.n44 VN.n43 0.189894
R78 VN.n43 VN.n34 0.189894
R79 VN.n39 VN.n34 0.189894
R80 VN.n39 VN.n38 0.189894
R81 VN.n10 VN.n9 0.189894
R82 VN.n10 VN.n5 0.189894
R83 VN.n14 VN.n5 0.189894
R84 VN.n15 VN.n14 0.189894
R85 VN.n16 VN.n15 0.189894
R86 VN.n16 VN.n3 0.189894
R87 VN.n21 VN.n3 0.189894
R88 VN.n22 VN.n21 0.189894
R89 VN.n23 VN.n22 0.189894
R90 VN.n23 VN.n1 0.189894
R91 VN.n27 VN.n1 0.189894
R92 VTAIL.n11 VTAIL.t4 90.7298
R93 VTAIL.n10 VTAIL.t13 90.7298
R94 VTAIL.n7 VTAIL.t8 90.7298
R95 VTAIL.n15 VTAIL.t12 90.7297
R96 VTAIL.n2 VTAIL.t11 90.7297
R97 VTAIL.n3 VTAIL.t5 90.7297
R98 VTAIL.n6 VTAIL.t6 90.7297
R99 VTAIL.n14 VTAIL.t2 90.7297
R100 VTAIL.n13 VTAIL.n12 84.1499
R101 VTAIL.n9 VTAIL.n8 84.1499
R102 VTAIL.n1 VTAIL.n0 84.1496
R103 VTAIL.n5 VTAIL.n4 84.1496
R104 VTAIL.n15 VTAIL.n14 19.3238
R105 VTAIL.n7 VTAIL.n6 19.3238
R106 VTAIL.n0 VTAIL.t10 6.58046
R107 VTAIL.n0 VTAIL.t15 6.58046
R108 VTAIL.n4 VTAIL.t3 6.58046
R109 VTAIL.n4 VTAIL.t0 6.58046
R110 VTAIL.n12 VTAIL.t1 6.58046
R111 VTAIL.n12 VTAIL.t7 6.58046
R112 VTAIL.n8 VTAIL.t9 6.58046
R113 VTAIL.n8 VTAIL.t14 6.58046
R114 VTAIL.n9 VTAIL.n7 2.69878
R115 VTAIL.n10 VTAIL.n9 2.69878
R116 VTAIL.n13 VTAIL.n11 2.69878
R117 VTAIL.n14 VTAIL.n13 2.69878
R118 VTAIL.n6 VTAIL.n5 2.69878
R119 VTAIL.n5 VTAIL.n3 2.69878
R120 VTAIL.n2 VTAIL.n1 2.69878
R121 VTAIL VTAIL.n15 2.64059
R122 VTAIL.n11 VTAIL.n10 0.470328
R123 VTAIL.n3 VTAIL.n2 0.470328
R124 VTAIL VTAIL.n1 0.0586897
R125 VDD2.n2 VDD2.n1 102.123
R126 VDD2.n2 VDD2.n0 102.123
R127 VDD2 VDD2.n5 102.12
R128 VDD2.n4 VDD2.n3 100.829
R129 VDD2.n4 VDD2.n2 40.1162
R130 VDD2.n5 VDD2.t6 6.58046
R131 VDD2.n5 VDD2.t3 6.58046
R132 VDD2.n3 VDD2.t0 6.58046
R133 VDD2.n3 VDD2.t7 6.58046
R134 VDD2.n1 VDD2.t4 6.58046
R135 VDD2.n1 VDD2.t2 6.58046
R136 VDD2.n0 VDD2.t5 6.58046
R137 VDD2.n0 VDD2.t1 6.58046
R138 VDD2 VDD2.n4 1.40783
R139 B.n492 B.n491 585
R140 B.n493 B.n58 585
R141 B.n495 B.n494 585
R142 B.n496 B.n57 585
R143 B.n498 B.n497 585
R144 B.n499 B.n56 585
R145 B.n501 B.n500 585
R146 B.n502 B.n55 585
R147 B.n504 B.n503 585
R148 B.n505 B.n54 585
R149 B.n507 B.n506 585
R150 B.n508 B.n53 585
R151 B.n510 B.n509 585
R152 B.n511 B.n52 585
R153 B.n513 B.n512 585
R154 B.n514 B.n51 585
R155 B.n516 B.n515 585
R156 B.n517 B.n50 585
R157 B.n519 B.n518 585
R158 B.n520 B.n49 585
R159 B.n522 B.n521 585
R160 B.n524 B.n523 585
R161 B.n525 B.n45 585
R162 B.n527 B.n526 585
R163 B.n528 B.n44 585
R164 B.n530 B.n529 585
R165 B.n531 B.n43 585
R166 B.n533 B.n532 585
R167 B.n534 B.n42 585
R168 B.n536 B.n535 585
R169 B.n538 B.n39 585
R170 B.n540 B.n539 585
R171 B.n541 B.n38 585
R172 B.n543 B.n542 585
R173 B.n544 B.n37 585
R174 B.n546 B.n545 585
R175 B.n547 B.n36 585
R176 B.n549 B.n548 585
R177 B.n550 B.n35 585
R178 B.n552 B.n551 585
R179 B.n553 B.n34 585
R180 B.n555 B.n554 585
R181 B.n556 B.n33 585
R182 B.n558 B.n557 585
R183 B.n559 B.n32 585
R184 B.n561 B.n560 585
R185 B.n562 B.n31 585
R186 B.n564 B.n563 585
R187 B.n565 B.n30 585
R188 B.n567 B.n566 585
R189 B.n568 B.n29 585
R190 B.n490 B.n59 585
R191 B.n489 B.n488 585
R192 B.n487 B.n60 585
R193 B.n486 B.n485 585
R194 B.n484 B.n61 585
R195 B.n483 B.n482 585
R196 B.n481 B.n62 585
R197 B.n480 B.n479 585
R198 B.n478 B.n63 585
R199 B.n477 B.n476 585
R200 B.n475 B.n64 585
R201 B.n474 B.n473 585
R202 B.n472 B.n65 585
R203 B.n471 B.n470 585
R204 B.n469 B.n66 585
R205 B.n468 B.n467 585
R206 B.n466 B.n67 585
R207 B.n465 B.n464 585
R208 B.n463 B.n68 585
R209 B.n462 B.n461 585
R210 B.n460 B.n69 585
R211 B.n459 B.n458 585
R212 B.n457 B.n70 585
R213 B.n456 B.n455 585
R214 B.n454 B.n71 585
R215 B.n453 B.n452 585
R216 B.n451 B.n72 585
R217 B.n450 B.n449 585
R218 B.n448 B.n73 585
R219 B.n447 B.n446 585
R220 B.n445 B.n74 585
R221 B.n444 B.n443 585
R222 B.n442 B.n75 585
R223 B.n441 B.n440 585
R224 B.n439 B.n76 585
R225 B.n438 B.n437 585
R226 B.n436 B.n77 585
R227 B.n435 B.n434 585
R228 B.n433 B.n78 585
R229 B.n432 B.n431 585
R230 B.n430 B.n79 585
R231 B.n429 B.n428 585
R232 B.n427 B.n80 585
R233 B.n426 B.n425 585
R234 B.n424 B.n81 585
R235 B.n423 B.n422 585
R236 B.n421 B.n82 585
R237 B.n420 B.n419 585
R238 B.n418 B.n83 585
R239 B.n417 B.n416 585
R240 B.n415 B.n84 585
R241 B.n414 B.n413 585
R242 B.n412 B.n85 585
R243 B.n411 B.n410 585
R244 B.n409 B.n86 585
R245 B.n408 B.n407 585
R246 B.n406 B.n87 585
R247 B.n405 B.n404 585
R248 B.n403 B.n88 585
R249 B.n402 B.n401 585
R250 B.n400 B.n89 585
R251 B.n399 B.n398 585
R252 B.n397 B.n90 585
R253 B.n396 B.n395 585
R254 B.n394 B.n91 585
R255 B.n393 B.n392 585
R256 B.n391 B.n92 585
R257 B.n390 B.n389 585
R258 B.n388 B.n93 585
R259 B.n387 B.n386 585
R260 B.n385 B.n94 585
R261 B.n384 B.n383 585
R262 B.n382 B.n95 585
R263 B.n381 B.n380 585
R264 B.n379 B.n96 585
R265 B.n378 B.n377 585
R266 B.n376 B.n97 585
R267 B.n375 B.n374 585
R268 B.n373 B.n98 585
R269 B.n372 B.n371 585
R270 B.n370 B.n99 585
R271 B.n369 B.n368 585
R272 B.n367 B.n100 585
R273 B.n366 B.n365 585
R274 B.n364 B.n101 585
R275 B.n363 B.n362 585
R276 B.n361 B.n102 585
R277 B.n360 B.n359 585
R278 B.n358 B.n103 585
R279 B.n357 B.n356 585
R280 B.n355 B.n104 585
R281 B.n354 B.n353 585
R282 B.n352 B.n105 585
R283 B.n351 B.n350 585
R284 B.n349 B.n106 585
R285 B.n348 B.n347 585
R286 B.n346 B.n107 585
R287 B.n345 B.n344 585
R288 B.n343 B.n108 585
R289 B.n342 B.n341 585
R290 B.n340 B.n109 585
R291 B.n339 B.n338 585
R292 B.n337 B.n110 585
R293 B.n336 B.n335 585
R294 B.n334 B.n111 585
R295 B.n333 B.n332 585
R296 B.n331 B.n112 585
R297 B.n330 B.n329 585
R298 B.n328 B.n113 585
R299 B.n250 B.n143 585
R300 B.n252 B.n251 585
R301 B.n253 B.n142 585
R302 B.n255 B.n254 585
R303 B.n256 B.n141 585
R304 B.n258 B.n257 585
R305 B.n259 B.n140 585
R306 B.n261 B.n260 585
R307 B.n262 B.n139 585
R308 B.n264 B.n263 585
R309 B.n265 B.n138 585
R310 B.n267 B.n266 585
R311 B.n268 B.n137 585
R312 B.n270 B.n269 585
R313 B.n271 B.n136 585
R314 B.n273 B.n272 585
R315 B.n274 B.n135 585
R316 B.n276 B.n275 585
R317 B.n277 B.n134 585
R318 B.n279 B.n278 585
R319 B.n280 B.n131 585
R320 B.n283 B.n282 585
R321 B.n284 B.n130 585
R322 B.n286 B.n285 585
R323 B.n287 B.n129 585
R324 B.n289 B.n288 585
R325 B.n290 B.n128 585
R326 B.n292 B.n291 585
R327 B.n293 B.n127 585
R328 B.n295 B.n294 585
R329 B.n297 B.n296 585
R330 B.n298 B.n123 585
R331 B.n300 B.n299 585
R332 B.n301 B.n122 585
R333 B.n303 B.n302 585
R334 B.n304 B.n121 585
R335 B.n306 B.n305 585
R336 B.n307 B.n120 585
R337 B.n309 B.n308 585
R338 B.n310 B.n119 585
R339 B.n312 B.n311 585
R340 B.n313 B.n118 585
R341 B.n315 B.n314 585
R342 B.n316 B.n117 585
R343 B.n318 B.n317 585
R344 B.n319 B.n116 585
R345 B.n321 B.n320 585
R346 B.n322 B.n115 585
R347 B.n324 B.n323 585
R348 B.n325 B.n114 585
R349 B.n327 B.n326 585
R350 B.n249 B.n248 585
R351 B.n247 B.n144 585
R352 B.n246 B.n245 585
R353 B.n244 B.n145 585
R354 B.n243 B.n242 585
R355 B.n241 B.n146 585
R356 B.n240 B.n239 585
R357 B.n238 B.n147 585
R358 B.n237 B.n236 585
R359 B.n235 B.n148 585
R360 B.n234 B.n233 585
R361 B.n232 B.n149 585
R362 B.n231 B.n230 585
R363 B.n229 B.n150 585
R364 B.n228 B.n227 585
R365 B.n226 B.n151 585
R366 B.n225 B.n224 585
R367 B.n223 B.n152 585
R368 B.n222 B.n221 585
R369 B.n220 B.n153 585
R370 B.n219 B.n218 585
R371 B.n217 B.n154 585
R372 B.n216 B.n215 585
R373 B.n214 B.n155 585
R374 B.n213 B.n212 585
R375 B.n211 B.n156 585
R376 B.n210 B.n209 585
R377 B.n208 B.n157 585
R378 B.n207 B.n206 585
R379 B.n205 B.n158 585
R380 B.n204 B.n203 585
R381 B.n202 B.n159 585
R382 B.n201 B.n200 585
R383 B.n199 B.n160 585
R384 B.n198 B.n197 585
R385 B.n196 B.n161 585
R386 B.n195 B.n194 585
R387 B.n193 B.n162 585
R388 B.n192 B.n191 585
R389 B.n190 B.n163 585
R390 B.n189 B.n188 585
R391 B.n187 B.n164 585
R392 B.n186 B.n185 585
R393 B.n184 B.n165 585
R394 B.n183 B.n182 585
R395 B.n181 B.n166 585
R396 B.n180 B.n179 585
R397 B.n178 B.n167 585
R398 B.n177 B.n176 585
R399 B.n175 B.n168 585
R400 B.n174 B.n173 585
R401 B.n172 B.n169 585
R402 B.n171 B.n170 585
R403 B.n2 B.n0 585
R404 B.n649 B.n1 585
R405 B.n648 B.n647 585
R406 B.n646 B.n3 585
R407 B.n645 B.n644 585
R408 B.n643 B.n4 585
R409 B.n642 B.n641 585
R410 B.n640 B.n5 585
R411 B.n639 B.n638 585
R412 B.n637 B.n6 585
R413 B.n636 B.n635 585
R414 B.n634 B.n7 585
R415 B.n633 B.n632 585
R416 B.n631 B.n8 585
R417 B.n630 B.n629 585
R418 B.n628 B.n9 585
R419 B.n627 B.n626 585
R420 B.n625 B.n10 585
R421 B.n624 B.n623 585
R422 B.n622 B.n11 585
R423 B.n621 B.n620 585
R424 B.n619 B.n12 585
R425 B.n618 B.n617 585
R426 B.n616 B.n13 585
R427 B.n615 B.n614 585
R428 B.n613 B.n14 585
R429 B.n612 B.n611 585
R430 B.n610 B.n15 585
R431 B.n609 B.n608 585
R432 B.n607 B.n16 585
R433 B.n606 B.n605 585
R434 B.n604 B.n17 585
R435 B.n603 B.n602 585
R436 B.n601 B.n18 585
R437 B.n600 B.n599 585
R438 B.n598 B.n19 585
R439 B.n597 B.n596 585
R440 B.n595 B.n20 585
R441 B.n594 B.n593 585
R442 B.n592 B.n21 585
R443 B.n591 B.n590 585
R444 B.n589 B.n22 585
R445 B.n588 B.n587 585
R446 B.n586 B.n23 585
R447 B.n585 B.n584 585
R448 B.n583 B.n24 585
R449 B.n582 B.n581 585
R450 B.n580 B.n25 585
R451 B.n579 B.n578 585
R452 B.n577 B.n26 585
R453 B.n576 B.n575 585
R454 B.n574 B.n27 585
R455 B.n573 B.n572 585
R456 B.n571 B.n28 585
R457 B.n570 B.n569 585
R458 B.n651 B.n650 585
R459 B.n248 B.n143 545.355
R460 B.n570 B.n29 545.355
R461 B.n326 B.n113 545.355
R462 B.n492 B.n59 545.355
R463 B.n124 B.t0 250.85
R464 B.n132 B.t9 250.85
R465 B.n40 B.t3 250.85
R466 B.n46 B.t6 250.85
R467 B.n124 B.t2 178.792
R468 B.n46 B.t7 178.792
R469 B.n132 B.t11 178.787
R470 B.n40 B.t4 178.787
R471 B.n248 B.n247 163.367
R472 B.n247 B.n246 163.367
R473 B.n246 B.n145 163.367
R474 B.n242 B.n145 163.367
R475 B.n242 B.n241 163.367
R476 B.n241 B.n240 163.367
R477 B.n240 B.n147 163.367
R478 B.n236 B.n147 163.367
R479 B.n236 B.n235 163.367
R480 B.n235 B.n234 163.367
R481 B.n234 B.n149 163.367
R482 B.n230 B.n149 163.367
R483 B.n230 B.n229 163.367
R484 B.n229 B.n228 163.367
R485 B.n228 B.n151 163.367
R486 B.n224 B.n151 163.367
R487 B.n224 B.n223 163.367
R488 B.n223 B.n222 163.367
R489 B.n222 B.n153 163.367
R490 B.n218 B.n153 163.367
R491 B.n218 B.n217 163.367
R492 B.n217 B.n216 163.367
R493 B.n216 B.n155 163.367
R494 B.n212 B.n155 163.367
R495 B.n212 B.n211 163.367
R496 B.n211 B.n210 163.367
R497 B.n210 B.n157 163.367
R498 B.n206 B.n157 163.367
R499 B.n206 B.n205 163.367
R500 B.n205 B.n204 163.367
R501 B.n204 B.n159 163.367
R502 B.n200 B.n159 163.367
R503 B.n200 B.n199 163.367
R504 B.n199 B.n198 163.367
R505 B.n198 B.n161 163.367
R506 B.n194 B.n161 163.367
R507 B.n194 B.n193 163.367
R508 B.n193 B.n192 163.367
R509 B.n192 B.n163 163.367
R510 B.n188 B.n163 163.367
R511 B.n188 B.n187 163.367
R512 B.n187 B.n186 163.367
R513 B.n186 B.n165 163.367
R514 B.n182 B.n165 163.367
R515 B.n182 B.n181 163.367
R516 B.n181 B.n180 163.367
R517 B.n180 B.n167 163.367
R518 B.n176 B.n167 163.367
R519 B.n176 B.n175 163.367
R520 B.n175 B.n174 163.367
R521 B.n174 B.n169 163.367
R522 B.n170 B.n169 163.367
R523 B.n170 B.n2 163.367
R524 B.n650 B.n2 163.367
R525 B.n650 B.n649 163.367
R526 B.n649 B.n648 163.367
R527 B.n648 B.n3 163.367
R528 B.n644 B.n3 163.367
R529 B.n644 B.n643 163.367
R530 B.n643 B.n642 163.367
R531 B.n642 B.n5 163.367
R532 B.n638 B.n5 163.367
R533 B.n638 B.n637 163.367
R534 B.n637 B.n636 163.367
R535 B.n636 B.n7 163.367
R536 B.n632 B.n7 163.367
R537 B.n632 B.n631 163.367
R538 B.n631 B.n630 163.367
R539 B.n630 B.n9 163.367
R540 B.n626 B.n9 163.367
R541 B.n626 B.n625 163.367
R542 B.n625 B.n624 163.367
R543 B.n624 B.n11 163.367
R544 B.n620 B.n11 163.367
R545 B.n620 B.n619 163.367
R546 B.n619 B.n618 163.367
R547 B.n618 B.n13 163.367
R548 B.n614 B.n13 163.367
R549 B.n614 B.n613 163.367
R550 B.n613 B.n612 163.367
R551 B.n612 B.n15 163.367
R552 B.n608 B.n15 163.367
R553 B.n608 B.n607 163.367
R554 B.n607 B.n606 163.367
R555 B.n606 B.n17 163.367
R556 B.n602 B.n17 163.367
R557 B.n602 B.n601 163.367
R558 B.n601 B.n600 163.367
R559 B.n600 B.n19 163.367
R560 B.n596 B.n19 163.367
R561 B.n596 B.n595 163.367
R562 B.n595 B.n594 163.367
R563 B.n594 B.n21 163.367
R564 B.n590 B.n21 163.367
R565 B.n590 B.n589 163.367
R566 B.n589 B.n588 163.367
R567 B.n588 B.n23 163.367
R568 B.n584 B.n23 163.367
R569 B.n584 B.n583 163.367
R570 B.n583 B.n582 163.367
R571 B.n582 B.n25 163.367
R572 B.n578 B.n25 163.367
R573 B.n578 B.n577 163.367
R574 B.n577 B.n576 163.367
R575 B.n576 B.n27 163.367
R576 B.n572 B.n27 163.367
R577 B.n572 B.n571 163.367
R578 B.n571 B.n570 163.367
R579 B.n252 B.n143 163.367
R580 B.n253 B.n252 163.367
R581 B.n254 B.n253 163.367
R582 B.n254 B.n141 163.367
R583 B.n258 B.n141 163.367
R584 B.n259 B.n258 163.367
R585 B.n260 B.n259 163.367
R586 B.n260 B.n139 163.367
R587 B.n264 B.n139 163.367
R588 B.n265 B.n264 163.367
R589 B.n266 B.n265 163.367
R590 B.n266 B.n137 163.367
R591 B.n270 B.n137 163.367
R592 B.n271 B.n270 163.367
R593 B.n272 B.n271 163.367
R594 B.n272 B.n135 163.367
R595 B.n276 B.n135 163.367
R596 B.n277 B.n276 163.367
R597 B.n278 B.n277 163.367
R598 B.n278 B.n131 163.367
R599 B.n283 B.n131 163.367
R600 B.n284 B.n283 163.367
R601 B.n285 B.n284 163.367
R602 B.n285 B.n129 163.367
R603 B.n289 B.n129 163.367
R604 B.n290 B.n289 163.367
R605 B.n291 B.n290 163.367
R606 B.n291 B.n127 163.367
R607 B.n295 B.n127 163.367
R608 B.n296 B.n295 163.367
R609 B.n296 B.n123 163.367
R610 B.n300 B.n123 163.367
R611 B.n301 B.n300 163.367
R612 B.n302 B.n301 163.367
R613 B.n302 B.n121 163.367
R614 B.n306 B.n121 163.367
R615 B.n307 B.n306 163.367
R616 B.n308 B.n307 163.367
R617 B.n308 B.n119 163.367
R618 B.n312 B.n119 163.367
R619 B.n313 B.n312 163.367
R620 B.n314 B.n313 163.367
R621 B.n314 B.n117 163.367
R622 B.n318 B.n117 163.367
R623 B.n319 B.n318 163.367
R624 B.n320 B.n319 163.367
R625 B.n320 B.n115 163.367
R626 B.n324 B.n115 163.367
R627 B.n325 B.n324 163.367
R628 B.n326 B.n325 163.367
R629 B.n330 B.n113 163.367
R630 B.n331 B.n330 163.367
R631 B.n332 B.n331 163.367
R632 B.n332 B.n111 163.367
R633 B.n336 B.n111 163.367
R634 B.n337 B.n336 163.367
R635 B.n338 B.n337 163.367
R636 B.n338 B.n109 163.367
R637 B.n342 B.n109 163.367
R638 B.n343 B.n342 163.367
R639 B.n344 B.n343 163.367
R640 B.n344 B.n107 163.367
R641 B.n348 B.n107 163.367
R642 B.n349 B.n348 163.367
R643 B.n350 B.n349 163.367
R644 B.n350 B.n105 163.367
R645 B.n354 B.n105 163.367
R646 B.n355 B.n354 163.367
R647 B.n356 B.n355 163.367
R648 B.n356 B.n103 163.367
R649 B.n360 B.n103 163.367
R650 B.n361 B.n360 163.367
R651 B.n362 B.n361 163.367
R652 B.n362 B.n101 163.367
R653 B.n366 B.n101 163.367
R654 B.n367 B.n366 163.367
R655 B.n368 B.n367 163.367
R656 B.n368 B.n99 163.367
R657 B.n372 B.n99 163.367
R658 B.n373 B.n372 163.367
R659 B.n374 B.n373 163.367
R660 B.n374 B.n97 163.367
R661 B.n378 B.n97 163.367
R662 B.n379 B.n378 163.367
R663 B.n380 B.n379 163.367
R664 B.n380 B.n95 163.367
R665 B.n384 B.n95 163.367
R666 B.n385 B.n384 163.367
R667 B.n386 B.n385 163.367
R668 B.n386 B.n93 163.367
R669 B.n390 B.n93 163.367
R670 B.n391 B.n390 163.367
R671 B.n392 B.n391 163.367
R672 B.n392 B.n91 163.367
R673 B.n396 B.n91 163.367
R674 B.n397 B.n396 163.367
R675 B.n398 B.n397 163.367
R676 B.n398 B.n89 163.367
R677 B.n402 B.n89 163.367
R678 B.n403 B.n402 163.367
R679 B.n404 B.n403 163.367
R680 B.n404 B.n87 163.367
R681 B.n408 B.n87 163.367
R682 B.n409 B.n408 163.367
R683 B.n410 B.n409 163.367
R684 B.n410 B.n85 163.367
R685 B.n414 B.n85 163.367
R686 B.n415 B.n414 163.367
R687 B.n416 B.n415 163.367
R688 B.n416 B.n83 163.367
R689 B.n420 B.n83 163.367
R690 B.n421 B.n420 163.367
R691 B.n422 B.n421 163.367
R692 B.n422 B.n81 163.367
R693 B.n426 B.n81 163.367
R694 B.n427 B.n426 163.367
R695 B.n428 B.n427 163.367
R696 B.n428 B.n79 163.367
R697 B.n432 B.n79 163.367
R698 B.n433 B.n432 163.367
R699 B.n434 B.n433 163.367
R700 B.n434 B.n77 163.367
R701 B.n438 B.n77 163.367
R702 B.n439 B.n438 163.367
R703 B.n440 B.n439 163.367
R704 B.n440 B.n75 163.367
R705 B.n444 B.n75 163.367
R706 B.n445 B.n444 163.367
R707 B.n446 B.n445 163.367
R708 B.n446 B.n73 163.367
R709 B.n450 B.n73 163.367
R710 B.n451 B.n450 163.367
R711 B.n452 B.n451 163.367
R712 B.n452 B.n71 163.367
R713 B.n456 B.n71 163.367
R714 B.n457 B.n456 163.367
R715 B.n458 B.n457 163.367
R716 B.n458 B.n69 163.367
R717 B.n462 B.n69 163.367
R718 B.n463 B.n462 163.367
R719 B.n464 B.n463 163.367
R720 B.n464 B.n67 163.367
R721 B.n468 B.n67 163.367
R722 B.n469 B.n468 163.367
R723 B.n470 B.n469 163.367
R724 B.n470 B.n65 163.367
R725 B.n474 B.n65 163.367
R726 B.n475 B.n474 163.367
R727 B.n476 B.n475 163.367
R728 B.n476 B.n63 163.367
R729 B.n480 B.n63 163.367
R730 B.n481 B.n480 163.367
R731 B.n482 B.n481 163.367
R732 B.n482 B.n61 163.367
R733 B.n486 B.n61 163.367
R734 B.n487 B.n486 163.367
R735 B.n488 B.n487 163.367
R736 B.n488 B.n59 163.367
R737 B.n566 B.n29 163.367
R738 B.n566 B.n565 163.367
R739 B.n565 B.n564 163.367
R740 B.n564 B.n31 163.367
R741 B.n560 B.n31 163.367
R742 B.n560 B.n559 163.367
R743 B.n559 B.n558 163.367
R744 B.n558 B.n33 163.367
R745 B.n554 B.n33 163.367
R746 B.n554 B.n553 163.367
R747 B.n553 B.n552 163.367
R748 B.n552 B.n35 163.367
R749 B.n548 B.n35 163.367
R750 B.n548 B.n547 163.367
R751 B.n547 B.n546 163.367
R752 B.n546 B.n37 163.367
R753 B.n542 B.n37 163.367
R754 B.n542 B.n541 163.367
R755 B.n541 B.n540 163.367
R756 B.n540 B.n39 163.367
R757 B.n535 B.n39 163.367
R758 B.n535 B.n534 163.367
R759 B.n534 B.n533 163.367
R760 B.n533 B.n43 163.367
R761 B.n529 B.n43 163.367
R762 B.n529 B.n528 163.367
R763 B.n528 B.n527 163.367
R764 B.n527 B.n45 163.367
R765 B.n523 B.n45 163.367
R766 B.n523 B.n522 163.367
R767 B.n522 B.n49 163.367
R768 B.n518 B.n49 163.367
R769 B.n518 B.n517 163.367
R770 B.n517 B.n516 163.367
R771 B.n516 B.n51 163.367
R772 B.n512 B.n51 163.367
R773 B.n512 B.n511 163.367
R774 B.n511 B.n510 163.367
R775 B.n510 B.n53 163.367
R776 B.n506 B.n53 163.367
R777 B.n506 B.n505 163.367
R778 B.n505 B.n504 163.367
R779 B.n504 B.n55 163.367
R780 B.n500 B.n55 163.367
R781 B.n500 B.n499 163.367
R782 B.n499 B.n498 163.367
R783 B.n498 B.n57 163.367
R784 B.n494 B.n57 163.367
R785 B.n494 B.n493 163.367
R786 B.n493 B.n492 163.367
R787 B.n125 B.t1 118.09
R788 B.n47 B.t8 118.09
R789 B.n133 B.t10 118.085
R790 B.n41 B.t5 118.085
R791 B.n125 B.n124 60.7035
R792 B.n133 B.n132 60.7035
R793 B.n41 B.n40 60.7035
R794 B.n47 B.n46 60.7035
R795 B.n126 B.n125 59.5399
R796 B.n281 B.n133 59.5399
R797 B.n537 B.n41 59.5399
R798 B.n48 B.n47 59.5399
R799 B.n569 B.n568 35.4346
R800 B.n328 B.n327 35.4346
R801 B.n250 B.n249 35.4346
R802 B.n491 B.n490 35.4346
R803 B B.n651 18.0485
R804 B.n568 B.n567 10.6151
R805 B.n567 B.n30 10.6151
R806 B.n563 B.n30 10.6151
R807 B.n563 B.n562 10.6151
R808 B.n562 B.n561 10.6151
R809 B.n561 B.n32 10.6151
R810 B.n557 B.n32 10.6151
R811 B.n557 B.n556 10.6151
R812 B.n556 B.n555 10.6151
R813 B.n555 B.n34 10.6151
R814 B.n551 B.n34 10.6151
R815 B.n551 B.n550 10.6151
R816 B.n550 B.n549 10.6151
R817 B.n549 B.n36 10.6151
R818 B.n545 B.n36 10.6151
R819 B.n545 B.n544 10.6151
R820 B.n544 B.n543 10.6151
R821 B.n543 B.n38 10.6151
R822 B.n539 B.n38 10.6151
R823 B.n539 B.n538 10.6151
R824 B.n536 B.n42 10.6151
R825 B.n532 B.n42 10.6151
R826 B.n532 B.n531 10.6151
R827 B.n531 B.n530 10.6151
R828 B.n530 B.n44 10.6151
R829 B.n526 B.n44 10.6151
R830 B.n526 B.n525 10.6151
R831 B.n525 B.n524 10.6151
R832 B.n521 B.n520 10.6151
R833 B.n520 B.n519 10.6151
R834 B.n519 B.n50 10.6151
R835 B.n515 B.n50 10.6151
R836 B.n515 B.n514 10.6151
R837 B.n514 B.n513 10.6151
R838 B.n513 B.n52 10.6151
R839 B.n509 B.n52 10.6151
R840 B.n509 B.n508 10.6151
R841 B.n508 B.n507 10.6151
R842 B.n507 B.n54 10.6151
R843 B.n503 B.n54 10.6151
R844 B.n503 B.n502 10.6151
R845 B.n502 B.n501 10.6151
R846 B.n501 B.n56 10.6151
R847 B.n497 B.n56 10.6151
R848 B.n497 B.n496 10.6151
R849 B.n496 B.n495 10.6151
R850 B.n495 B.n58 10.6151
R851 B.n491 B.n58 10.6151
R852 B.n329 B.n328 10.6151
R853 B.n329 B.n112 10.6151
R854 B.n333 B.n112 10.6151
R855 B.n334 B.n333 10.6151
R856 B.n335 B.n334 10.6151
R857 B.n335 B.n110 10.6151
R858 B.n339 B.n110 10.6151
R859 B.n340 B.n339 10.6151
R860 B.n341 B.n340 10.6151
R861 B.n341 B.n108 10.6151
R862 B.n345 B.n108 10.6151
R863 B.n346 B.n345 10.6151
R864 B.n347 B.n346 10.6151
R865 B.n347 B.n106 10.6151
R866 B.n351 B.n106 10.6151
R867 B.n352 B.n351 10.6151
R868 B.n353 B.n352 10.6151
R869 B.n353 B.n104 10.6151
R870 B.n357 B.n104 10.6151
R871 B.n358 B.n357 10.6151
R872 B.n359 B.n358 10.6151
R873 B.n359 B.n102 10.6151
R874 B.n363 B.n102 10.6151
R875 B.n364 B.n363 10.6151
R876 B.n365 B.n364 10.6151
R877 B.n365 B.n100 10.6151
R878 B.n369 B.n100 10.6151
R879 B.n370 B.n369 10.6151
R880 B.n371 B.n370 10.6151
R881 B.n371 B.n98 10.6151
R882 B.n375 B.n98 10.6151
R883 B.n376 B.n375 10.6151
R884 B.n377 B.n376 10.6151
R885 B.n377 B.n96 10.6151
R886 B.n381 B.n96 10.6151
R887 B.n382 B.n381 10.6151
R888 B.n383 B.n382 10.6151
R889 B.n383 B.n94 10.6151
R890 B.n387 B.n94 10.6151
R891 B.n388 B.n387 10.6151
R892 B.n389 B.n388 10.6151
R893 B.n389 B.n92 10.6151
R894 B.n393 B.n92 10.6151
R895 B.n394 B.n393 10.6151
R896 B.n395 B.n394 10.6151
R897 B.n395 B.n90 10.6151
R898 B.n399 B.n90 10.6151
R899 B.n400 B.n399 10.6151
R900 B.n401 B.n400 10.6151
R901 B.n401 B.n88 10.6151
R902 B.n405 B.n88 10.6151
R903 B.n406 B.n405 10.6151
R904 B.n407 B.n406 10.6151
R905 B.n407 B.n86 10.6151
R906 B.n411 B.n86 10.6151
R907 B.n412 B.n411 10.6151
R908 B.n413 B.n412 10.6151
R909 B.n413 B.n84 10.6151
R910 B.n417 B.n84 10.6151
R911 B.n418 B.n417 10.6151
R912 B.n419 B.n418 10.6151
R913 B.n419 B.n82 10.6151
R914 B.n423 B.n82 10.6151
R915 B.n424 B.n423 10.6151
R916 B.n425 B.n424 10.6151
R917 B.n425 B.n80 10.6151
R918 B.n429 B.n80 10.6151
R919 B.n430 B.n429 10.6151
R920 B.n431 B.n430 10.6151
R921 B.n431 B.n78 10.6151
R922 B.n435 B.n78 10.6151
R923 B.n436 B.n435 10.6151
R924 B.n437 B.n436 10.6151
R925 B.n437 B.n76 10.6151
R926 B.n441 B.n76 10.6151
R927 B.n442 B.n441 10.6151
R928 B.n443 B.n442 10.6151
R929 B.n443 B.n74 10.6151
R930 B.n447 B.n74 10.6151
R931 B.n448 B.n447 10.6151
R932 B.n449 B.n448 10.6151
R933 B.n449 B.n72 10.6151
R934 B.n453 B.n72 10.6151
R935 B.n454 B.n453 10.6151
R936 B.n455 B.n454 10.6151
R937 B.n455 B.n70 10.6151
R938 B.n459 B.n70 10.6151
R939 B.n460 B.n459 10.6151
R940 B.n461 B.n460 10.6151
R941 B.n461 B.n68 10.6151
R942 B.n465 B.n68 10.6151
R943 B.n466 B.n465 10.6151
R944 B.n467 B.n466 10.6151
R945 B.n467 B.n66 10.6151
R946 B.n471 B.n66 10.6151
R947 B.n472 B.n471 10.6151
R948 B.n473 B.n472 10.6151
R949 B.n473 B.n64 10.6151
R950 B.n477 B.n64 10.6151
R951 B.n478 B.n477 10.6151
R952 B.n479 B.n478 10.6151
R953 B.n479 B.n62 10.6151
R954 B.n483 B.n62 10.6151
R955 B.n484 B.n483 10.6151
R956 B.n485 B.n484 10.6151
R957 B.n485 B.n60 10.6151
R958 B.n489 B.n60 10.6151
R959 B.n490 B.n489 10.6151
R960 B.n251 B.n250 10.6151
R961 B.n251 B.n142 10.6151
R962 B.n255 B.n142 10.6151
R963 B.n256 B.n255 10.6151
R964 B.n257 B.n256 10.6151
R965 B.n257 B.n140 10.6151
R966 B.n261 B.n140 10.6151
R967 B.n262 B.n261 10.6151
R968 B.n263 B.n262 10.6151
R969 B.n263 B.n138 10.6151
R970 B.n267 B.n138 10.6151
R971 B.n268 B.n267 10.6151
R972 B.n269 B.n268 10.6151
R973 B.n269 B.n136 10.6151
R974 B.n273 B.n136 10.6151
R975 B.n274 B.n273 10.6151
R976 B.n275 B.n274 10.6151
R977 B.n275 B.n134 10.6151
R978 B.n279 B.n134 10.6151
R979 B.n280 B.n279 10.6151
R980 B.n282 B.n130 10.6151
R981 B.n286 B.n130 10.6151
R982 B.n287 B.n286 10.6151
R983 B.n288 B.n287 10.6151
R984 B.n288 B.n128 10.6151
R985 B.n292 B.n128 10.6151
R986 B.n293 B.n292 10.6151
R987 B.n294 B.n293 10.6151
R988 B.n298 B.n297 10.6151
R989 B.n299 B.n298 10.6151
R990 B.n299 B.n122 10.6151
R991 B.n303 B.n122 10.6151
R992 B.n304 B.n303 10.6151
R993 B.n305 B.n304 10.6151
R994 B.n305 B.n120 10.6151
R995 B.n309 B.n120 10.6151
R996 B.n310 B.n309 10.6151
R997 B.n311 B.n310 10.6151
R998 B.n311 B.n118 10.6151
R999 B.n315 B.n118 10.6151
R1000 B.n316 B.n315 10.6151
R1001 B.n317 B.n316 10.6151
R1002 B.n317 B.n116 10.6151
R1003 B.n321 B.n116 10.6151
R1004 B.n322 B.n321 10.6151
R1005 B.n323 B.n322 10.6151
R1006 B.n323 B.n114 10.6151
R1007 B.n327 B.n114 10.6151
R1008 B.n249 B.n144 10.6151
R1009 B.n245 B.n144 10.6151
R1010 B.n245 B.n244 10.6151
R1011 B.n244 B.n243 10.6151
R1012 B.n243 B.n146 10.6151
R1013 B.n239 B.n146 10.6151
R1014 B.n239 B.n238 10.6151
R1015 B.n238 B.n237 10.6151
R1016 B.n237 B.n148 10.6151
R1017 B.n233 B.n148 10.6151
R1018 B.n233 B.n232 10.6151
R1019 B.n232 B.n231 10.6151
R1020 B.n231 B.n150 10.6151
R1021 B.n227 B.n150 10.6151
R1022 B.n227 B.n226 10.6151
R1023 B.n226 B.n225 10.6151
R1024 B.n225 B.n152 10.6151
R1025 B.n221 B.n152 10.6151
R1026 B.n221 B.n220 10.6151
R1027 B.n220 B.n219 10.6151
R1028 B.n219 B.n154 10.6151
R1029 B.n215 B.n154 10.6151
R1030 B.n215 B.n214 10.6151
R1031 B.n214 B.n213 10.6151
R1032 B.n213 B.n156 10.6151
R1033 B.n209 B.n156 10.6151
R1034 B.n209 B.n208 10.6151
R1035 B.n208 B.n207 10.6151
R1036 B.n207 B.n158 10.6151
R1037 B.n203 B.n158 10.6151
R1038 B.n203 B.n202 10.6151
R1039 B.n202 B.n201 10.6151
R1040 B.n201 B.n160 10.6151
R1041 B.n197 B.n160 10.6151
R1042 B.n197 B.n196 10.6151
R1043 B.n196 B.n195 10.6151
R1044 B.n195 B.n162 10.6151
R1045 B.n191 B.n162 10.6151
R1046 B.n191 B.n190 10.6151
R1047 B.n190 B.n189 10.6151
R1048 B.n189 B.n164 10.6151
R1049 B.n185 B.n164 10.6151
R1050 B.n185 B.n184 10.6151
R1051 B.n184 B.n183 10.6151
R1052 B.n183 B.n166 10.6151
R1053 B.n179 B.n166 10.6151
R1054 B.n179 B.n178 10.6151
R1055 B.n178 B.n177 10.6151
R1056 B.n177 B.n168 10.6151
R1057 B.n173 B.n168 10.6151
R1058 B.n173 B.n172 10.6151
R1059 B.n172 B.n171 10.6151
R1060 B.n171 B.n0 10.6151
R1061 B.n647 B.n1 10.6151
R1062 B.n647 B.n646 10.6151
R1063 B.n646 B.n645 10.6151
R1064 B.n645 B.n4 10.6151
R1065 B.n641 B.n4 10.6151
R1066 B.n641 B.n640 10.6151
R1067 B.n640 B.n639 10.6151
R1068 B.n639 B.n6 10.6151
R1069 B.n635 B.n6 10.6151
R1070 B.n635 B.n634 10.6151
R1071 B.n634 B.n633 10.6151
R1072 B.n633 B.n8 10.6151
R1073 B.n629 B.n8 10.6151
R1074 B.n629 B.n628 10.6151
R1075 B.n628 B.n627 10.6151
R1076 B.n627 B.n10 10.6151
R1077 B.n623 B.n10 10.6151
R1078 B.n623 B.n622 10.6151
R1079 B.n622 B.n621 10.6151
R1080 B.n621 B.n12 10.6151
R1081 B.n617 B.n12 10.6151
R1082 B.n617 B.n616 10.6151
R1083 B.n616 B.n615 10.6151
R1084 B.n615 B.n14 10.6151
R1085 B.n611 B.n14 10.6151
R1086 B.n611 B.n610 10.6151
R1087 B.n610 B.n609 10.6151
R1088 B.n609 B.n16 10.6151
R1089 B.n605 B.n16 10.6151
R1090 B.n605 B.n604 10.6151
R1091 B.n604 B.n603 10.6151
R1092 B.n603 B.n18 10.6151
R1093 B.n599 B.n18 10.6151
R1094 B.n599 B.n598 10.6151
R1095 B.n598 B.n597 10.6151
R1096 B.n597 B.n20 10.6151
R1097 B.n593 B.n20 10.6151
R1098 B.n593 B.n592 10.6151
R1099 B.n592 B.n591 10.6151
R1100 B.n591 B.n22 10.6151
R1101 B.n587 B.n22 10.6151
R1102 B.n587 B.n586 10.6151
R1103 B.n586 B.n585 10.6151
R1104 B.n585 B.n24 10.6151
R1105 B.n581 B.n24 10.6151
R1106 B.n581 B.n580 10.6151
R1107 B.n580 B.n579 10.6151
R1108 B.n579 B.n26 10.6151
R1109 B.n575 B.n26 10.6151
R1110 B.n575 B.n574 10.6151
R1111 B.n574 B.n573 10.6151
R1112 B.n573 B.n28 10.6151
R1113 B.n569 B.n28 10.6151
R1114 B.n537 B.n536 6.5566
R1115 B.n524 B.n48 6.5566
R1116 B.n282 B.n281 6.5566
R1117 B.n294 B.n126 6.5566
R1118 B.n538 B.n537 4.05904
R1119 B.n521 B.n48 4.05904
R1120 B.n281 B.n280 4.05904
R1121 B.n297 B.n126 4.05904
R1122 B.n651 B.n0 2.81026
R1123 B.n651 B.n1 2.81026
R1124 VP.n19 VP.n16 161.3
R1125 VP.n21 VP.n20 161.3
R1126 VP.n22 VP.n15 161.3
R1127 VP.n24 VP.n23 161.3
R1128 VP.n25 VP.n14 161.3
R1129 VP.n27 VP.n26 161.3
R1130 VP.n29 VP.n13 161.3
R1131 VP.n31 VP.n30 161.3
R1132 VP.n32 VP.n12 161.3
R1133 VP.n34 VP.n33 161.3
R1134 VP.n35 VP.n11 161.3
R1135 VP.n37 VP.n36 161.3
R1136 VP.n69 VP.n68 161.3
R1137 VP.n67 VP.n1 161.3
R1138 VP.n66 VP.n65 161.3
R1139 VP.n64 VP.n2 161.3
R1140 VP.n63 VP.n62 161.3
R1141 VP.n61 VP.n3 161.3
R1142 VP.n59 VP.n58 161.3
R1143 VP.n57 VP.n4 161.3
R1144 VP.n56 VP.n55 161.3
R1145 VP.n54 VP.n5 161.3
R1146 VP.n53 VP.n52 161.3
R1147 VP.n51 VP.n6 161.3
R1148 VP.n50 VP.n49 161.3
R1149 VP.n47 VP.n7 161.3
R1150 VP.n46 VP.n45 161.3
R1151 VP.n44 VP.n8 161.3
R1152 VP.n43 VP.n42 161.3
R1153 VP.n41 VP.n9 161.3
R1154 VP.n18 VP.t3 74.4814
R1155 VP.n40 VP.n39 68.3588
R1156 VP.n70 VP.n0 68.3588
R1157 VP.n38 VP.n10 68.3588
R1158 VP.n18 VP.n17 58.3802
R1159 VP.n55 VP.n54 56.5617
R1160 VP.n23 VP.n22 56.5617
R1161 VP.n46 VP.n8 52.2023
R1162 VP.n66 VP.n2 52.2023
R1163 VP.n34 VP.n12 52.2023
R1164 VP.n39 VP.n38 46.5829
R1165 VP.n40 VP.t5 42.5198
R1166 VP.n48 VP.t2 42.5198
R1167 VP.n60 VP.t6 42.5198
R1168 VP.n0 VP.t4 42.5198
R1169 VP.n10 VP.t1 42.5198
R1170 VP.n28 VP.t7 42.5198
R1171 VP.n17 VP.t0 42.5198
R1172 VP.n42 VP.n8 28.9518
R1173 VP.n67 VP.n66 28.9518
R1174 VP.n35 VP.n34 28.9518
R1175 VP.n42 VP.n41 24.5923
R1176 VP.n47 VP.n46 24.5923
R1177 VP.n49 VP.n47 24.5923
R1178 VP.n53 VP.n6 24.5923
R1179 VP.n54 VP.n53 24.5923
R1180 VP.n55 VP.n4 24.5923
R1181 VP.n59 VP.n4 24.5923
R1182 VP.n62 VP.n61 24.5923
R1183 VP.n62 VP.n2 24.5923
R1184 VP.n68 VP.n67 24.5923
R1185 VP.n36 VP.n35 24.5923
R1186 VP.n23 VP.n14 24.5923
R1187 VP.n27 VP.n14 24.5923
R1188 VP.n30 VP.n29 24.5923
R1189 VP.n30 VP.n12 24.5923
R1190 VP.n21 VP.n16 24.5923
R1191 VP.n22 VP.n21 24.5923
R1192 VP.n41 VP.n40 21.8872
R1193 VP.n68 VP.n0 21.8872
R1194 VP.n36 VP.n10 21.8872
R1195 VP.n48 VP.n6 15.4934
R1196 VP.n60 VP.n59 15.4934
R1197 VP.n28 VP.n27 15.4934
R1198 VP.n17 VP.n16 15.4934
R1199 VP.n49 VP.n48 9.09948
R1200 VP.n61 VP.n60 9.09948
R1201 VP.n29 VP.n28 9.09948
R1202 VP.n19 VP.n18 5.3904
R1203 VP.n38 VP.n37 0.354861
R1204 VP.n39 VP.n9 0.354861
R1205 VP.n70 VP.n69 0.354861
R1206 VP VP.n70 0.267071
R1207 VP.n20 VP.n19 0.189894
R1208 VP.n20 VP.n15 0.189894
R1209 VP.n24 VP.n15 0.189894
R1210 VP.n25 VP.n24 0.189894
R1211 VP.n26 VP.n25 0.189894
R1212 VP.n26 VP.n13 0.189894
R1213 VP.n31 VP.n13 0.189894
R1214 VP.n32 VP.n31 0.189894
R1215 VP.n33 VP.n32 0.189894
R1216 VP.n33 VP.n11 0.189894
R1217 VP.n37 VP.n11 0.189894
R1218 VP.n43 VP.n9 0.189894
R1219 VP.n44 VP.n43 0.189894
R1220 VP.n45 VP.n44 0.189894
R1221 VP.n45 VP.n7 0.189894
R1222 VP.n50 VP.n7 0.189894
R1223 VP.n51 VP.n50 0.189894
R1224 VP.n52 VP.n51 0.189894
R1225 VP.n52 VP.n5 0.189894
R1226 VP.n56 VP.n5 0.189894
R1227 VP.n57 VP.n56 0.189894
R1228 VP.n58 VP.n57 0.189894
R1229 VP.n58 VP.n3 0.189894
R1230 VP.n63 VP.n3 0.189894
R1231 VP.n64 VP.n63 0.189894
R1232 VP.n65 VP.n64 0.189894
R1233 VP.n65 VP.n1 0.189894
R1234 VP.n69 VP.n1 0.189894
R1235 VDD1 VDD1.n0 102.237
R1236 VDD1.n3 VDD1.n2 102.123
R1237 VDD1.n3 VDD1.n1 102.123
R1238 VDD1.n5 VDD1.n4 100.829
R1239 VDD1.n5 VDD1.n3 40.6992
R1240 VDD1.n4 VDD1.t0 6.58046
R1241 VDD1.n4 VDD1.t6 6.58046
R1242 VDD1.n0 VDD1.t4 6.58046
R1243 VDD1.n0 VDD1.t7 6.58046
R1244 VDD1.n2 VDD1.t1 6.58046
R1245 VDD1.n2 VDD1.t3 6.58046
R1246 VDD1.n1 VDD1.t2 6.58046
R1247 VDD1.n1 VDD1.t5 6.58046
R1248 VDD1 VDD1.n5 1.29145
C0 B VTAIL 2.70599f
C1 VDD2 VP 0.545538f
C2 VN VP 6.59775f
C3 VDD2 VDD1 1.88109f
C4 VP B 2.12353f
C5 VDD1 VN 0.152358f
C6 VDD1 B 1.51939f
C7 VP VTAIL 4.89131f
C8 VDD2 w_n4100_n1956# 1.95176f
C9 VDD1 VTAIL 5.84378f
C10 w_n4100_n1956# VN 8.27799f
C11 w_n4100_n1956# B 8.456281f
C12 w_n4100_n1956# VTAIL 2.64306f
C13 VDD1 VP 4.28688f
C14 w_n4100_n1956# VP 8.81076f
C15 VDD2 VN 3.89967f
C16 VDD2 B 1.62182f
C17 w_n4100_n1956# VDD1 1.82896f
C18 VN B 1.2293f
C19 VDD2 VTAIL 5.89953f
C20 VN VTAIL 4.8772f
C21 VDD2 VSUBS 1.577552f
C22 VDD1 VSUBS 2.275379f
C23 VTAIL VSUBS 0.687588f
C24 VN VSUBS 6.75085f
C25 VP VSUBS 3.290928f
C26 B VSUBS 4.36209f
C27 w_n4100_n1956# VSUBS 0.100516p
C28 VDD1.t4 VSUBS 0.096373f
C29 VDD1.t7 VSUBS 0.096373f
C30 VDD1.n0 VSUBS 0.613127f
C31 VDD1.t2 VSUBS 0.096373f
C32 VDD1.t5 VSUBS 0.096373f
C33 VDD1.n1 VSUBS 0.612233f
C34 VDD1.t1 VSUBS 0.096373f
C35 VDD1.t3 VSUBS 0.096373f
C36 VDD1.n2 VSUBS 0.612233f
C37 VDD1.n3 VSUBS 3.3236f
C38 VDD1.t0 VSUBS 0.096373f
C39 VDD1.t6 VSUBS 0.096373f
C40 VDD1.n4 VSUBS 0.603308f
C41 VDD1.n5 VSUBS 2.64664f
C42 VP.t4 VSUBS 1.55342f
C43 VP.n0 VSUBS 0.758475f
C44 VP.n1 VSUBS 0.042974f
C45 VP.n2 VSUBS 0.076778f
C46 VP.n3 VSUBS 0.042974f
C47 VP.t6 VSUBS 1.55342f
C48 VP.n4 VSUBS 0.079691f
C49 VP.n5 VSUBS 0.042974f
C50 VP.n6 VSUBS 0.065135f
C51 VP.n7 VSUBS 0.042974f
C52 VP.n8 VSUBS 0.043303f
C53 VP.n9 VSUBS 0.069348f
C54 VP.t5 VSUBS 1.55342f
C55 VP.t1 VSUBS 1.55342f
C56 VP.n10 VSUBS 0.758475f
C57 VP.n11 VSUBS 0.042974f
C58 VP.n12 VSUBS 0.076778f
C59 VP.n13 VSUBS 0.042974f
C60 VP.t7 VSUBS 1.55342f
C61 VP.n14 VSUBS 0.079691f
C62 VP.n15 VSUBS 0.042974f
C63 VP.n16 VSUBS 0.065135f
C64 VP.t3 VSUBS 1.92745f
C65 VP.t0 VSUBS 1.55342f
C66 VP.n17 VSUBS 0.730637f
C67 VP.n18 VSUBS 0.699679f
C68 VP.n19 VSUBS 0.453256f
C69 VP.n20 VSUBS 0.042974f
C70 VP.n21 VSUBS 0.079691f
C71 VP.n22 VSUBS 0.062469f
C72 VP.n23 VSUBS 0.062469f
C73 VP.n24 VSUBS 0.042974f
C74 VP.n25 VSUBS 0.042974f
C75 VP.n26 VSUBS 0.042974f
C76 VP.n27 VSUBS 0.065135f
C77 VP.n28 VSUBS 0.594616f
C78 VP.n29 VSUBS 0.054906f
C79 VP.n30 VSUBS 0.079691f
C80 VP.n31 VSUBS 0.042974f
C81 VP.n32 VSUBS 0.042974f
C82 VP.n33 VSUBS 0.042974f
C83 VP.n34 VSUBS 0.043303f
C84 VP.n35 VSUBS 0.084549f
C85 VP.n36 VSUBS 0.075363f
C86 VP.n37 VSUBS 0.069348f
C87 VP.n38 VSUBS 2.18073f
C88 VP.n39 VSUBS 2.21399f
C89 VP.n40 VSUBS 0.758475f
C90 VP.n41 VSUBS 0.075363f
C91 VP.n42 VSUBS 0.084549f
C92 VP.n43 VSUBS 0.042974f
C93 VP.n44 VSUBS 0.042974f
C94 VP.n45 VSUBS 0.042974f
C95 VP.n46 VSUBS 0.076778f
C96 VP.n47 VSUBS 0.079691f
C97 VP.t2 VSUBS 1.55342f
C98 VP.n48 VSUBS 0.594616f
C99 VP.n49 VSUBS 0.054906f
C100 VP.n50 VSUBS 0.042974f
C101 VP.n51 VSUBS 0.042974f
C102 VP.n52 VSUBS 0.042974f
C103 VP.n53 VSUBS 0.079691f
C104 VP.n54 VSUBS 0.062469f
C105 VP.n55 VSUBS 0.062469f
C106 VP.n56 VSUBS 0.042974f
C107 VP.n57 VSUBS 0.042974f
C108 VP.n58 VSUBS 0.042974f
C109 VP.n59 VSUBS 0.065135f
C110 VP.n60 VSUBS 0.594616f
C111 VP.n61 VSUBS 0.054906f
C112 VP.n62 VSUBS 0.079691f
C113 VP.n63 VSUBS 0.042974f
C114 VP.n64 VSUBS 0.042974f
C115 VP.n65 VSUBS 0.042974f
C116 VP.n66 VSUBS 0.043303f
C117 VP.n67 VSUBS 0.084549f
C118 VP.n68 VSUBS 0.075363f
C119 VP.n69 VSUBS 0.069348f
C120 VP.n70 VSUBS 0.083224f
C121 B.n0 VSUBS 0.006372f
C122 B.n1 VSUBS 0.006372f
C123 B.n2 VSUBS 0.010076f
C124 B.n3 VSUBS 0.010076f
C125 B.n4 VSUBS 0.010076f
C126 B.n5 VSUBS 0.010076f
C127 B.n6 VSUBS 0.010076f
C128 B.n7 VSUBS 0.010076f
C129 B.n8 VSUBS 0.010076f
C130 B.n9 VSUBS 0.010076f
C131 B.n10 VSUBS 0.010076f
C132 B.n11 VSUBS 0.010076f
C133 B.n12 VSUBS 0.010076f
C134 B.n13 VSUBS 0.010076f
C135 B.n14 VSUBS 0.010076f
C136 B.n15 VSUBS 0.010076f
C137 B.n16 VSUBS 0.010076f
C138 B.n17 VSUBS 0.010076f
C139 B.n18 VSUBS 0.010076f
C140 B.n19 VSUBS 0.010076f
C141 B.n20 VSUBS 0.010076f
C142 B.n21 VSUBS 0.010076f
C143 B.n22 VSUBS 0.010076f
C144 B.n23 VSUBS 0.010076f
C145 B.n24 VSUBS 0.010076f
C146 B.n25 VSUBS 0.010076f
C147 B.n26 VSUBS 0.010076f
C148 B.n27 VSUBS 0.010076f
C149 B.n28 VSUBS 0.010076f
C150 B.n29 VSUBS 0.025416f
C151 B.n30 VSUBS 0.010076f
C152 B.n31 VSUBS 0.010076f
C153 B.n32 VSUBS 0.010076f
C154 B.n33 VSUBS 0.010076f
C155 B.n34 VSUBS 0.010076f
C156 B.n35 VSUBS 0.010076f
C157 B.n36 VSUBS 0.010076f
C158 B.n37 VSUBS 0.010076f
C159 B.n38 VSUBS 0.010076f
C160 B.n39 VSUBS 0.010076f
C161 B.t5 VSUBS 0.197938f
C162 B.t4 VSUBS 0.227722f
C163 B.t3 VSUBS 0.952851f
C164 B.n40 VSUBS 0.150104f
C165 B.n41 VSUBS 0.102093f
C166 B.n42 VSUBS 0.010076f
C167 B.n43 VSUBS 0.010076f
C168 B.n44 VSUBS 0.010076f
C169 B.n45 VSUBS 0.010076f
C170 B.t8 VSUBS 0.197938f
C171 B.t7 VSUBS 0.227721f
C172 B.t6 VSUBS 0.952851f
C173 B.n46 VSUBS 0.150105f
C174 B.n47 VSUBS 0.102093f
C175 B.n48 VSUBS 0.023346f
C176 B.n49 VSUBS 0.010076f
C177 B.n50 VSUBS 0.010076f
C178 B.n51 VSUBS 0.010076f
C179 B.n52 VSUBS 0.010076f
C180 B.n53 VSUBS 0.010076f
C181 B.n54 VSUBS 0.010076f
C182 B.n55 VSUBS 0.010076f
C183 B.n56 VSUBS 0.010076f
C184 B.n57 VSUBS 0.010076f
C185 B.n58 VSUBS 0.010076f
C186 B.n59 VSUBS 0.024372f
C187 B.n60 VSUBS 0.010076f
C188 B.n61 VSUBS 0.010076f
C189 B.n62 VSUBS 0.010076f
C190 B.n63 VSUBS 0.010076f
C191 B.n64 VSUBS 0.010076f
C192 B.n65 VSUBS 0.010076f
C193 B.n66 VSUBS 0.010076f
C194 B.n67 VSUBS 0.010076f
C195 B.n68 VSUBS 0.010076f
C196 B.n69 VSUBS 0.010076f
C197 B.n70 VSUBS 0.010076f
C198 B.n71 VSUBS 0.010076f
C199 B.n72 VSUBS 0.010076f
C200 B.n73 VSUBS 0.010076f
C201 B.n74 VSUBS 0.010076f
C202 B.n75 VSUBS 0.010076f
C203 B.n76 VSUBS 0.010076f
C204 B.n77 VSUBS 0.010076f
C205 B.n78 VSUBS 0.010076f
C206 B.n79 VSUBS 0.010076f
C207 B.n80 VSUBS 0.010076f
C208 B.n81 VSUBS 0.010076f
C209 B.n82 VSUBS 0.010076f
C210 B.n83 VSUBS 0.010076f
C211 B.n84 VSUBS 0.010076f
C212 B.n85 VSUBS 0.010076f
C213 B.n86 VSUBS 0.010076f
C214 B.n87 VSUBS 0.010076f
C215 B.n88 VSUBS 0.010076f
C216 B.n89 VSUBS 0.010076f
C217 B.n90 VSUBS 0.010076f
C218 B.n91 VSUBS 0.010076f
C219 B.n92 VSUBS 0.010076f
C220 B.n93 VSUBS 0.010076f
C221 B.n94 VSUBS 0.010076f
C222 B.n95 VSUBS 0.010076f
C223 B.n96 VSUBS 0.010076f
C224 B.n97 VSUBS 0.010076f
C225 B.n98 VSUBS 0.010076f
C226 B.n99 VSUBS 0.010076f
C227 B.n100 VSUBS 0.010076f
C228 B.n101 VSUBS 0.010076f
C229 B.n102 VSUBS 0.010076f
C230 B.n103 VSUBS 0.010076f
C231 B.n104 VSUBS 0.010076f
C232 B.n105 VSUBS 0.010076f
C233 B.n106 VSUBS 0.010076f
C234 B.n107 VSUBS 0.010076f
C235 B.n108 VSUBS 0.010076f
C236 B.n109 VSUBS 0.010076f
C237 B.n110 VSUBS 0.010076f
C238 B.n111 VSUBS 0.010076f
C239 B.n112 VSUBS 0.010076f
C240 B.n113 VSUBS 0.024372f
C241 B.n114 VSUBS 0.010076f
C242 B.n115 VSUBS 0.010076f
C243 B.n116 VSUBS 0.010076f
C244 B.n117 VSUBS 0.010076f
C245 B.n118 VSUBS 0.010076f
C246 B.n119 VSUBS 0.010076f
C247 B.n120 VSUBS 0.010076f
C248 B.n121 VSUBS 0.010076f
C249 B.n122 VSUBS 0.010076f
C250 B.n123 VSUBS 0.010076f
C251 B.t1 VSUBS 0.197938f
C252 B.t2 VSUBS 0.227721f
C253 B.t0 VSUBS 0.952851f
C254 B.n124 VSUBS 0.150105f
C255 B.n125 VSUBS 0.102093f
C256 B.n126 VSUBS 0.023346f
C257 B.n127 VSUBS 0.010076f
C258 B.n128 VSUBS 0.010076f
C259 B.n129 VSUBS 0.010076f
C260 B.n130 VSUBS 0.010076f
C261 B.n131 VSUBS 0.010076f
C262 B.t10 VSUBS 0.197938f
C263 B.t11 VSUBS 0.227722f
C264 B.t9 VSUBS 0.952851f
C265 B.n132 VSUBS 0.150104f
C266 B.n133 VSUBS 0.102093f
C267 B.n134 VSUBS 0.010076f
C268 B.n135 VSUBS 0.010076f
C269 B.n136 VSUBS 0.010076f
C270 B.n137 VSUBS 0.010076f
C271 B.n138 VSUBS 0.010076f
C272 B.n139 VSUBS 0.010076f
C273 B.n140 VSUBS 0.010076f
C274 B.n141 VSUBS 0.010076f
C275 B.n142 VSUBS 0.010076f
C276 B.n143 VSUBS 0.025416f
C277 B.n144 VSUBS 0.010076f
C278 B.n145 VSUBS 0.010076f
C279 B.n146 VSUBS 0.010076f
C280 B.n147 VSUBS 0.010076f
C281 B.n148 VSUBS 0.010076f
C282 B.n149 VSUBS 0.010076f
C283 B.n150 VSUBS 0.010076f
C284 B.n151 VSUBS 0.010076f
C285 B.n152 VSUBS 0.010076f
C286 B.n153 VSUBS 0.010076f
C287 B.n154 VSUBS 0.010076f
C288 B.n155 VSUBS 0.010076f
C289 B.n156 VSUBS 0.010076f
C290 B.n157 VSUBS 0.010076f
C291 B.n158 VSUBS 0.010076f
C292 B.n159 VSUBS 0.010076f
C293 B.n160 VSUBS 0.010076f
C294 B.n161 VSUBS 0.010076f
C295 B.n162 VSUBS 0.010076f
C296 B.n163 VSUBS 0.010076f
C297 B.n164 VSUBS 0.010076f
C298 B.n165 VSUBS 0.010076f
C299 B.n166 VSUBS 0.010076f
C300 B.n167 VSUBS 0.010076f
C301 B.n168 VSUBS 0.010076f
C302 B.n169 VSUBS 0.010076f
C303 B.n170 VSUBS 0.010076f
C304 B.n171 VSUBS 0.010076f
C305 B.n172 VSUBS 0.010076f
C306 B.n173 VSUBS 0.010076f
C307 B.n174 VSUBS 0.010076f
C308 B.n175 VSUBS 0.010076f
C309 B.n176 VSUBS 0.010076f
C310 B.n177 VSUBS 0.010076f
C311 B.n178 VSUBS 0.010076f
C312 B.n179 VSUBS 0.010076f
C313 B.n180 VSUBS 0.010076f
C314 B.n181 VSUBS 0.010076f
C315 B.n182 VSUBS 0.010076f
C316 B.n183 VSUBS 0.010076f
C317 B.n184 VSUBS 0.010076f
C318 B.n185 VSUBS 0.010076f
C319 B.n186 VSUBS 0.010076f
C320 B.n187 VSUBS 0.010076f
C321 B.n188 VSUBS 0.010076f
C322 B.n189 VSUBS 0.010076f
C323 B.n190 VSUBS 0.010076f
C324 B.n191 VSUBS 0.010076f
C325 B.n192 VSUBS 0.010076f
C326 B.n193 VSUBS 0.010076f
C327 B.n194 VSUBS 0.010076f
C328 B.n195 VSUBS 0.010076f
C329 B.n196 VSUBS 0.010076f
C330 B.n197 VSUBS 0.010076f
C331 B.n198 VSUBS 0.010076f
C332 B.n199 VSUBS 0.010076f
C333 B.n200 VSUBS 0.010076f
C334 B.n201 VSUBS 0.010076f
C335 B.n202 VSUBS 0.010076f
C336 B.n203 VSUBS 0.010076f
C337 B.n204 VSUBS 0.010076f
C338 B.n205 VSUBS 0.010076f
C339 B.n206 VSUBS 0.010076f
C340 B.n207 VSUBS 0.010076f
C341 B.n208 VSUBS 0.010076f
C342 B.n209 VSUBS 0.010076f
C343 B.n210 VSUBS 0.010076f
C344 B.n211 VSUBS 0.010076f
C345 B.n212 VSUBS 0.010076f
C346 B.n213 VSUBS 0.010076f
C347 B.n214 VSUBS 0.010076f
C348 B.n215 VSUBS 0.010076f
C349 B.n216 VSUBS 0.010076f
C350 B.n217 VSUBS 0.010076f
C351 B.n218 VSUBS 0.010076f
C352 B.n219 VSUBS 0.010076f
C353 B.n220 VSUBS 0.010076f
C354 B.n221 VSUBS 0.010076f
C355 B.n222 VSUBS 0.010076f
C356 B.n223 VSUBS 0.010076f
C357 B.n224 VSUBS 0.010076f
C358 B.n225 VSUBS 0.010076f
C359 B.n226 VSUBS 0.010076f
C360 B.n227 VSUBS 0.010076f
C361 B.n228 VSUBS 0.010076f
C362 B.n229 VSUBS 0.010076f
C363 B.n230 VSUBS 0.010076f
C364 B.n231 VSUBS 0.010076f
C365 B.n232 VSUBS 0.010076f
C366 B.n233 VSUBS 0.010076f
C367 B.n234 VSUBS 0.010076f
C368 B.n235 VSUBS 0.010076f
C369 B.n236 VSUBS 0.010076f
C370 B.n237 VSUBS 0.010076f
C371 B.n238 VSUBS 0.010076f
C372 B.n239 VSUBS 0.010076f
C373 B.n240 VSUBS 0.010076f
C374 B.n241 VSUBS 0.010076f
C375 B.n242 VSUBS 0.010076f
C376 B.n243 VSUBS 0.010076f
C377 B.n244 VSUBS 0.010076f
C378 B.n245 VSUBS 0.010076f
C379 B.n246 VSUBS 0.010076f
C380 B.n247 VSUBS 0.010076f
C381 B.n248 VSUBS 0.024372f
C382 B.n249 VSUBS 0.024372f
C383 B.n250 VSUBS 0.025416f
C384 B.n251 VSUBS 0.010076f
C385 B.n252 VSUBS 0.010076f
C386 B.n253 VSUBS 0.010076f
C387 B.n254 VSUBS 0.010076f
C388 B.n255 VSUBS 0.010076f
C389 B.n256 VSUBS 0.010076f
C390 B.n257 VSUBS 0.010076f
C391 B.n258 VSUBS 0.010076f
C392 B.n259 VSUBS 0.010076f
C393 B.n260 VSUBS 0.010076f
C394 B.n261 VSUBS 0.010076f
C395 B.n262 VSUBS 0.010076f
C396 B.n263 VSUBS 0.010076f
C397 B.n264 VSUBS 0.010076f
C398 B.n265 VSUBS 0.010076f
C399 B.n266 VSUBS 0.010076f
C400 B.n267 VSUBS 0.010076f
C401 B.n268 VSUBS 0.010076f
C402 B.n269 VSUBS 0.010076f
C403 B.n270 VSUBS 0.010076f
C404 B.n271 VSUBS 0.010076f
C405 B.n272 VSUBS 0.010076f
C406 B.n273 VSUBS 0.010076f
C407 B.n274 VSUBS 0.010076f
C408 B.n275 VSUBS 0.010076f
C409 B.n276 VSUBS 0.010076f
C410 B.n277 VSUBS 0.010076f
C411 B.n278 VSUBS 0.010076f
C412 B.n279 VSUBS 0.010076f
C413 B.n280 VSUBS 0.006964f
C414 B.n281 VSUBS 0.023346f
C415 B.n282 VSUBS 0.00815f
C416 B.n283 VSUBS 0.010076f
C417 B.n284 VSUBS 0.010076f
C418 B.n285 VSUBS 0.010076f
C419 B.n286 VSUBS 0.010076f
C420 B.n287 VSUBS 0.010076f
C421 B.n288 VSUBS 0.010076f
C422 B.n289 VSUBS 0.010076f
C423 B.n290 VSUBS 0.010076f
C424 B.n291 VSUBS 0.010076f
C425 B.n292 VSUBS 0.010076f
C426 B.n293 VSUBS 0.010076f
C427 B.n294 VSUBS 0.00815f
C428 B.n295 VSUBS 0.010076f
C429 B.n296 VSUBS 0.010076f
C430 B.n297 VSUBS 0.006964f
C431 B.n298 VSUBS 0.010076f
C432 B.n299 VSUBS 0.010076f
C433 B.n300 VSUBS 0.010076f
C434 B.n301 VSUBS 0.010076f
C435 B.n302 VSUBS 0.010076f
C436 B.n303 VSUBS 0.010076f
C437 B.n304 VSUBS 0.010076f
C438 B.n305 VSUBS 0.010076f
C439 B.n306 VSUBS 0.010076f
C440 B.n307 VSUBS 0.010076f
C441 B.n308 VSUBS 0.010076f
C442 B.n309 VSUBS 0.010076f
C443 B.n310 VSUBS 0.010076f
C444 B.n311 VSUBS 0.010076f
C445 B.n312 VSUBS 0.010076f
C446 B.n313 VSUBS 0.010076f
C447 B.n314 VSUBS 0.010076f
C448 B.n315 VSUBS 0.010076f
C449 B.n316 VSUBS 0.010076f
C450 B.n317 VSUBS 0.010076f
C451 B.n318 VSUBS 0.010076f
C452 B.n319 VSUBS 0.010076f
C453 B.n320 VSUBS 0.010076f
C454 B.n321 VSUBS 0.010076f
C455 B.n322 VSUBS 0.010076f
C456 B.n323 VSUBS 0.010076f
C457 B.n324 VSUBS 0.010076f
C458 B.n325 VSUBS 0.010076f
C459 B.n326 VSUBS 0.025416f
C460 B.n327 VSUBS 0.025416f
C461 B.n328 VSUBS 0.024372f
C462 B.n329 VSUBS 0.010076f
C463 B.n330 VSUBS 0.010076f
C464 B.n331 VSUBS 0.010076f
C465 B.n332 VSUBS 0.010076f
C466 B.n333 VSUBS 0.010076f
C467 B.n334 VSUBS 0.010076f
C468 B.n335 VSUBS 0.010076f
C469 B.n336 VSUBS 0.010076f
C470 B.n337 VSUBS 0.010076f
C471 B.n338 VSUBS 0.010076f
C472 B.n339 VSUBS 0.010076f
C473 B.n340 VSUBS 0.010076f
C474 B.n341 VSUBS 0.010076f
C475 B.n342 VSUBS 0.010076f
C476 B.n343 VSUBS 0.010076f
C477 B.n344 VSUBS 0.010076f
C478 B.n345 VSUBS 0.010076f
C479 B.n346 VSUBS 0.010076f
C480 B.n347 VSUBS 0.010076f
C481 B.n348 VSUBS 0.010076f
C482 B.n349 VSUBS 0.010076f
C483 B.n350 VSUBS 0.010076f
C484 B.n351 VSUBS 0.010076f
C485 B.n352 VSUBS 0.010076f
C486 B.n353 VSUBS 0.010076f
C487 B.n354 VSUBS 0.010076f
C488 B.n355 VSUBS 0.010076f
C489 B.n356 VSUBS 0.010076f
C490 B.n357 VSUBS 0.010076f
C491 B.n358 VSUBS 0.010076f
C492 B.n359 VSUBS 0.010076f
C493 B.n360 VSUBS 0.010076f
C494 B.n361 VSUBS 0.010076f
C495 B.n362 VSUBS 0.010076f
C496 B.n363 VSUBS 0.010076f
C497 B.n364 VSUBS 0.010076f
C498 B.n365 VSUBS 0.010076f
C499 B.n366 VSUBS 0.010076f
C500 B.n367 VSUBS 0.010076f
C501 B.n368 VSUBS 0.010076f
C502 B.n369 VSUBS 0.010076f
C503 B.n370 VSUBS 0.010076f
C504 B.n371 VSUBS 0.010076f
C505 B.n372 VSUBS 0.010076f
C506 B.n373 VSUBS 0.010076f
C507 B.n374 VSUBS 0.010076f
C508 B.n375 VSUBS 0.010076f
C509 B.n376 VSUBS 0.010076f
C510 B.n377 VSUBS 0.010076f
C511 B.n378 VSUBS 0.010076f
C512 B.n379 VSUBS 0.010076f
C513 B.n380 VSUBS 0.010076f
C514 B.n381 VSUBS 0.010076f
C515 B.n382 VSUBS 0.010076f
C516 B.n383 VSUBS 0.010076f
C517 B.n384 VSUBS 0.010076f
C518 B.n385 VSUBS 0.010076f
C519 B.n386 VSUBS 0.010076f
C520 B.n387 VSUBS 0.010076f
C521 B.n388 VSUBS 0.010076f
C522 B.n389 VSUBS 0.010076f
C523 B.n390 VSUBS 0.010076f
C524 B.n391 VSUBS 0.010076f
C525 B.n392 VSUBS 0.010076f
C526 B.n393 VSUBS 0.010076f
C527 B.n394 VSUBS 0.010076f
C528 B.n395 VSUBS 0.010076f
C529 B.n396 VSUBS 0.010076f
C530 B.n397 VSUBS 0.010076f
C531 B.n398 VSUBS 0.010076f
C532 B.n399 VSUBS 0.010076f
C533 B.n400 VSUBS 0.010076f
C534 B.n401 VSUBS 0.010076f
C535 B.n402 VSUBS 0.010076f
C536 B.n403 VSUBS 0.010076f
C537 B.n404 VSUBS 0.010076f
C538 B.n405 VSUBS 0.010076f
C539 B.n406 VSUBS 0.010076f
C540 B.n407 VSUBS 0.010076f
C541 B.n408 VSUBS 0.010076f
C542 B.n409 VSUBS 0.010076f
C543 B.n410 VSUBS 0.010076f
C544 B.n411 VSUBS 0.010076f
C545 B.n412 VSUBS 0.010076f
C546 B.n413 VSUBS 0.010076f
C547 B.n414 VSUBS 0.010076f
C548 B.n415 VSUBS 0.010076f
C549 B.n416 VSUBS 0.010076f
C550 B.n417 VSUBS 0.010076f
C551 B.n418 VSUBS 0.010076f
C552 B.n419 VSUBS 0.010076f
C553 B.n420 VSUBS 0.010076f
C554 B.n421 VSUBS 0.010076f
C555 B.n422 VSUBS 0.010076f
C556 B.n423 VSUBS 0.010076f
C557 B.n424 VSUBS 0.010076f
C558 B.n425 VSUBS 0.010076f
C559 B.n426 VSUBS 0.010076f
C560 B.n427 VSUBS 0.010076f
C561 B.n428 VSUBS 0.010076f
C562 B.n429 VSUBS 0.010076f
C563 B.n430 VSUBS 0.010076f
C564 B.n431 VSUBS 0.010076f
C565 B.n432 VSUBS 0.010076f
C566 B.n433 VSUBS 0.010076f
C567 B.n434 VSUBS 0.010076f
C568 B.n435 VSUBS 0.010076f
C569 B.n436 VSUBS 0.010076f
C570 B.n437 VSUBS 0.010076f
C571 B.n438 VSUBS 0.010076f
C572 B.n439 VSUBS 0.010076f
C573 B.n440 VSUBS 0.010076f
C574 B.n441 VSUBS 0.010076f
C575 B.n442 VSUBS 0.010076f
C576 B.n443 VSUBS 0.010076f
C577 B.n444 VSUBS 0.010076f
C578 B.n445 VSUBS 0.010076f
C579 B.n446 VSUBS 0.010076f
C580 B.n447 VSUBS 0.010076f
C581 B.n448 VSUBS 0.010076f
C582 B.n449 VSUBS 0.010076f
C583 B.n450 VSUBS 0.010076f
C584 B.n451 VSUBS 0.010076f
C585 B.n452 VSUBS 0.010076f
C586 B.n453 VSUBS 0.010076f
C587 B.n454 VSUBS 0.010076f
C588 B.n455 VSUBS 0.010076f
C589 B.n456 VSUBS 0.010076f
C590 B.n457 VSUBS 0.010076f
C591 B.n458 VSUBS 0.010076f
C592 B.n459 VSUBS 0.010076f
C593 B.n460 VSUBS 0.010076f
C594 B.n461 VSUBS 0.010076f
C595 B.n462 VSUBS 0.010076f
C596 B.n463 VSUBS 0.010076f
C597 B.n464 VSUBS 0.010076f
C598 B.n465 VSUBS 0.010076f
C599 B.n466 VSUBS 0.010076f
C600 B.n467 VSUBS 0.010076f
C601 B.n468 VSUBS 0.010076f
C602 B.n469 VSUBS 0.010076f
C603 B.n470 VSUBS 0.010076f
C604 B.n471 VSUBS 0.010076f
C605 B.n472 VSUBS 0.010076f
C606 B.n473 VSUBS 0.010076f
C607 B.n474 VSUBS 0.010076f
C608 B.n475 VSUBS 0.010076f
C609 B.n476 VSUBS 0.010076f
C610 B.n477 VSUBS 0.010076f
C611 B.n478 VSUBS 0.010076f
C612 B.n479 VSUBS 0.010076f
C613 B.n480 VSUBS 0.010076f
C614 B.n481 VSUBS 0.010076f
C615 B.n482 VSUBS 0.010076f
C616 B.n483 VSUBS 0.010076f
C617 B.n484 VSUBS 0.010076f
C618 B.n485 VSUBS 0.010076f
C619 B.n486 VSUBS 0.010076f
C620 B.n487 VSUBS 0.010076f
C621 B.n488 VSUBS 0.010076f
C622 B.n489 VSUBS 0.010076f
C623 B.n490 VSUBS 0.02547f
C624 B.n491 VSUBS 0.024319f
C625 B.n492 VSUBS 0.025416f
C626 B.n493 VSUBS 0.010076f
C627 B.n494 VSUBS 0.010076f
C628 B.n495 VSUBS 0.010076f
C629 B.n496 VSUBS 0.010076f
C630 B.n497 VSUBS 0.010076f
C631 B.n498 VSUBS 0.010076f
C632 B.n499 VSUBS 0.010076f
C633 B.n500 VSUBS 0.010076f
C634 B.n501 VSUBS 0.010076f
C635 B.n502 VSUBS 0.010076f
C636 B.n503 VSUBS 0.010076f
C637 B.n504 VSUBS 0.010076f
C638 B.n505 VSUBS 0.010076f
C639 B.n506 VSUBS 0.010076f
C640 B.n507 VSUBS 0.010076f
C641 B.n508 VSUBS 0.010076f
C642 B.n509 VSUBS 0.010076f
C643 B.n510 VSUBS 0.010076f
C644 B.n511 VSUBS 0.010076f
C645 B.n512 VSUBS 0.010076f
C646 B.n513 VSUBS 0.010076f
C647 B.n514 VSUBS 0.010076f
C648 B.n515 VSUBS 0.010076f
C649 B.n516 VSUBS 0.010076f
C650 B.n517 VSUBS 0.010076f
C651 B.n518 VSUBS 0.010076f
C652 B.n519 VSUBS 0.010076f
C653 B.n520 VSUBS 0.010076f
C654 B.n521 VSUBS 0.006964f
C655 B.n522 VSUBS 0.010076f
C656 B.n523 VSUBS 0.010076f
C657 B.n524 VSUBS 0.00815f
C658 B.n525 VSUBS 0.010076f
C659 B.n526 VSUBS 0.010076f
C660 B.n527 VSUBS 0.010076f
C661 B.n528 VSUBS 0.010076f
C662 B.n529 VSUBS 0.010076f
C663 B.n530 VSUBS 0.010076f
C664 B.n531 VSUBS 0.010076f
C665 B.n532 VSUBS 0.010076f
C666 B.n533 VSUBS 0.010076f
C667 B.n534 VSUBS 0.010076f
C668 B.n535 VSUBS 0.010076f
C669 B.n536 VSUBS 0.00815f
C670 B.n537 VSUBS 0.023346f
C671 B.n538 VSUBS 0.006964f
C672 B.n539 VSUBS 0.010076f
C673 B.n540 VSUBS 0.010076f
C674 B.n541 VSUBS 0.010076f
C675 B.n542 VSUBS 0.010076f
C676 B.n543 VSUBS 0.010076f
C677 B.n544 VSUBS 0.010076f
C678 B.n545 VSUBS 0.010076f
C679 B.n546 VSUBS 0.010076f
C680 B.n547 VSUBS 0.010076f
C681 B.n548 VSUBS 0.010076f
C682 B.n549 VSUBS 0.010076f
C683 B.n550 VSUBS 0.010076f
C684 B.n551 VSUBS 0.010076f
C685 B.n552 VSUBS 0.010076f
C686 B.n553 VSUBS 0.010076f
C687 B.n554 VSUBS 0.010076f
C688 B.n555 VSUBS 0.010076f
C689 B.n556 VSUBS 0.010076f
C690 B.n557 VSUBS 0.010076f
C691 B.n558 VSUBS 0.010076f
C692 B.n559 VSUBS 0.010076f
C693 B.n560 VSUBS 0.010076f
C694 B.n561 VSUBS 0.010076f
C695 B.n562 VSUBS 0.010076f
C696 B.n563 VSUBS 0.010076f
C697 B.n564 VSUBS 0.010076f
C698 B.n565 VSUBS 0.010076f
C699 B.n566 VSUBS 0.010076f
C700 B.n567 VSUBS 0.010076f
C701 B.n568 VSUBS 0.025416f
C702 B.n569 VSUBS 0.024372f
C703 B.n570 VSUBS 0.024372f
C704 B.n571 VSUBS 0.010076f
C705 B.n572 VSUBS 0.010076f
C706 B.n573 VSUBS 0.010076f
C707 B.n574 VSUBS 0.010076f
C708 B.n575 VSUBS 0.010076f
C709 B.n576 VSUBS 0.010076f
C710 B.n577 VSUBS 0.010076f
C711 B.n578 VSUBS 0.010076f
C712 B.n579 VSUBS 0.010076f
C713 B.n580 VSUBS 0.010076f
C714 B.n581 VSUBS 0.010076f
C715 B.n582 VSUBS 0.010076f
C716 B.n583 VSUBS 0.010076f
C717 B.n584 VSUBS 0.010076f
C718 B.n585 VSUBS 0.010076f
C719 B.n586 VSUBS 0.010076f
C720 B.n587 VSUBS 0.010076f
C721 B.n588 VSUBS 0.010076f
C722 B.n589 VSUBS 0.010076f
C723 B.n590 VSUBS 0.010076f
C724 B.n591 VSUBS 0.010076f
C725 B.n592 VSUBS 0.010076f
C726 B.n593 VSUBS 0.010076f
C727 B.n594 VSUBS 0.010076f
C728 B.n595 VSUBS 0.010076f
C729 B.n596 VSUBS 0.010076f
C730 B.n597 VSUBS 0.010076f
C731 B.n598 VSUBS 0.010076f
C732 B.n599 VSUBS 0.010076f
C733 B.n600 VSUBS 0.010076f
C734 B.n601 VSUBS 0.010076f
C735 B.n602 VSUBS 0.010076f
C736 B.n603 VSUBS 0.010076f
C737 B.n604 VSUBS 0.010076f
C738 B.n605 VSUBS 0.010076f
C739 B.n606 VSUBS 0.010076f
C740 B.n607 VSUBS 0.010076f
C741 B.n608 VSUBS 0.010076f
C742 B.n609 VSUBS 0.010076f
C743 B.n610 VSUBS 0.010076f
C744 B.n611 VSUBS 0.010076f
C745 B.n612 VSUBS 0.010076f
C746 B.n613 VSUBS 0.010076f
C747 B.n614 VSUBS 0.010076f
C748 B.n615 VSUBS 0.010076f
C749 B.n616 VSUBS 0.010076f
C750 B.n617 VSUBS 0.010076f
C751 B.n618 VSUBS 0.010076f
C752 B.n619 VSUBS 0.010076f
C753 B.n620 VSUBS 0.010076f
C754 B.n621 VSUBS 0.010076f
C755 B.n622 VSUBS 0.010076f
C756 B.n623 VSUBS 0.010076f
C757 B.n624 VSUBS 0.010076f
C758 B.n625 VSUBS 0.010076f
C759 B.n626 VSUBS 0.010076f
C760 B.n627 VSUBS 0.010076f
C761 B.n628 VSUBS 0.010076f
C762 B.n629 VSUBS 0.010076f
C763 B.n630 VSUBS 0.010076f
C764 B.n631 VSUBS 0.010076f
C765 B.n632 VSUBS 0.010076f
C766 B.n633 VSUBS 0.010076f
C767 B.n634 VSUBS 0.010076f
C768 B.n635 VSUBS 0.010076f
C769 B.n636 VSUBS 0.010076f
C770 B.n637 VSUBS 0.010076f
C771 B.n638 VSUBS 0.010076f
C772 B.n639 VSUBS 0.010076f
C773 B.n640 VSUBS 0.010076f
C774 B.n641 VSUBS 0.010076f
C775 B.n642 VSUBS 0.010076f
C776 B.n643 VSUBS 0.010076f
C777 B.n644 VSUBS 0.010076f
C778 B.n645 VSUBS 0.010076f
C779 B.n646 VSUBS 0.010076f
C780 B.n647 VSUBS 0.010076f
C781 B.n648 VSUBS 0.010076f
C782 B.n649 VSUBS 0.010076f
C783 B.n650 VSUBS 0.010076f
C784 B.n651 VSUBS 0.022816f
C785 VDD2.t5 VSUBS 0.094363f
C786 VDD2.t1 VSUBS 0.094363f
C787 VDD2.n0 VSUBS 0.59946f
C788 VDD2.t4 VSUBS 0.094363f
C789 VDD2.t2 VSUBS 0.094363f
C790 VDD2.n1 VSUBS 0.59946f
C791 VDD2.n2 VSUBS 3.20383f
C792 VDD2.t0 VSUBS 0.094363f
C793 VDD2.t7 VSUBS 0.094363f
C794 VDD2.n3 VSUBS 0.590724f
C795 VDD2.n4 VSUBS 2.56163f
C796 VDD2.t6 VSUBS 0.094363f
C797 VDD2.t3 VSUBS 0.094363f
C798 VDD2.n5 VSUBS 0.599432f
C799 VTAIL.t10 VSUBS 0.120874f
C800 VTAIL.t15 VSUBS 0.120874f
C801 VTAIL.n0 VSUBS 0.664255f
C802 VTAIL.n1 VSUBS 0.797599f
C803 VTAIL.t11 VSUBS 0.930595f
C804 VTAIL.n2 VSUBS 0.901985f
C805 VTAIL.t5 VSUBS 0.930595f
C806 VTAIL.n3 VSUBS 0.901985f
C807 VTAIL.t3 VSUBS 0.120874f
C808 VTAIL.t0 VSUBS 0.120874f
C809 VTAIL.n4 VSUBS 0.664255f
C810 VTAIL.n5 VSUBS 1.06101f
C811 VTAIL.t6 VSUBS 0.930595f
C812 VTAIL.n6 VSUBS 1.96982f
C813 VTAIL.t8 VSUBS 0.9306f
C814 VTAIL.n7 VSUBS 1.96981f
C815 VTAIL.t9 VSUBS 0.120874f
C816 VTAIL.t14 VSUBS 0.120874f
C817 VTAIL.n8 VSUBS 0.664259f
C818 VTAIL.n9 VSUBS 1.061f
C819 VTAIL.t13 VSUBS 0.9306f
C820 VTAIL.n10 VSUBS 0.90198f
C821 VTAIL.t4 VSUBS 0.9306f
C822 VTAIL.n11 VSUBS 0.90198f
C823 VTAIL.t1 VSUBS 0.120874f
C824 VTAIL.t7 VSUBS 0.120874f
C825 VTAIL.n12 VSUBS 0.664259f
C826 VTAIL.n13 VSUBS 1.061f
C827 VTAIL.t2 VSUBS 0.930595f
C828 VTAIL.n14 VSUBS 1.96982f
C829 VTAIL.t12 VSUBS 0.930595f
C830 VTAIL.n15 VSUBS 1.96401f
C831 VN.t5 VSUBS 1.37577f
C832 VN.n0 VSUBS 0.671733f
C833 VN.n1 VSUBS 0.038059f
C834 VN.n2 VSUBS 0.067997f
C835 VN.n3 VSUBS 0.038059f
C836 VN.t3 VSUBS 1.37577f
C837 VN.n4 VSUBS 0.070577f
C838 VN.n5 VSUBS 0.038059f
C839 VN.n6 VSUBS 0.057686f
C840 VN.t6 VSUBS 1.37577f
C841 VN.n7 VSUBS 0.647079f
C842 VN.t2 VSUBS 1.70702f
C843 VN.n8 VSUBS 0.61966f
C844 VN.n9 VSUBS 0.401419f
C845 VN.n10 VSUBS 0.038059f
C846 VN.n11 VSUBS 0.070577f
C847 VN.n12 VSUBS 0.055325f
C848 VN.n13 VSUBS 0.055325f
C849 VN.n14 VSUBS 0.038059f
C850 VN.n15 VSUBS 0.038059f
C851 VN.n16 VSUBS 0.038059f
C852 VN.n17 VSUBS 0.057686f
C853 VN.n18 VSUBS 0.526614f
C854 VN.n19 VSUBS 0.048627f
C855 VN.n20 VSUBS 0.070577f
C856 VN.n21 VSUBS 0.038059f
C857 VN.n22 VSUBS 0.038059f
C858 VN.n23 VSUBS 0.038059f
C859 VN.n24 VSUBS 0.03835f
C860 VN.n25 VSUBS 0.074879f
C861 VN.n26 VSUBS 0.066745f
C862 VN.n27 VSUBS 0.061417f
C863 VN.n28 VSUBS 0.073706f
C864 VN.t7 VSUBS 1.37577f
C865 VN.n29 VSUBS 0.671733f
C866 VN.n30 VSUBS 0.038059f
C867 VN.n31 VSUBS 0.067997f
C868 VN.n32 VSUBS 0.038059f
C869 VN.t0 VSUBS 1.37577f
C870 VN.n33 VSUBS 0.070577f
C871 VN.n34 VSUBS 0.038059f
C872 VN.n35 VSUBS 0.057686f
C873 VN.t4 VSUBS 1.70702f
C874 VN.t1 VSUBS 1.37577f
C875 VN.n36 VSUBS 0.647079f
C876 VN.n37 VSUBS 0.61966f
C877 VN.n38 VSUBS 0.401419f
C878 VN.n39 VSUBS 0.038059f
C879 VN.n40 VSUBS 0.070577f
C880 VN.n41 VSUBS 0.055325f
C881 VN.n42 VSUBS 0.055325f
C882 VN.n43 VSUBS 0.038059f
C883 VN.n44 VSUBS 0.038059f
C884 VN.n45 VSUBS 0.038059f
C885 VN.n46 VSUBS 0.057686f
C886 VN.n47 VSUBS 0.526614f
C887 VN.n48 VSUBS 0.048627f
C888 VN.n49 VSUBS 0.070577f
C889 VN.n50 VSUBS 0.038059f
C890 VN.n51 VSUBS 0.038059f
C891 VN.n52 VSUBS 0.038059f
C892 VN.n53 VSUBS 0.03835f
C893 VN.n54 VSUBS 0.074879f
C894 VN.n55 VSUBS 0.066745f
C895 VN.n56 VSUBS 0.061417f
C896 VN.n57 VSUBS 1.94731f
.ends

