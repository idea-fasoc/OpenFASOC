* NGSPICE file created from diff_pair_sample_0214.ext - technology: sky130A

.subckt diff_pair_sample_0214 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t7 w_n2114_n1078# sky130_fd_pr__pfet_01v8 ad=0.2145 pd=1.88 as=0.09075 ps=0.88 w=0.55 l=1.1
X1 B.t11 B.t9 B.t10 w_n2114_n1078# sky130_fd_pr__pfet_01v8 ad=0.2145 pd=1.88 as=0 ps=0 w=0.55 l=1.1
X2 VTAIL.t5 VN.t0 VDD2.t5 w_n2114_n1078# sky130_fd_pr__pfet_01v8 ad=0.09075 pd=0.88 as=0.09075 ps=0.88 w=0.55 l=1.1
X3 VDD2.t4 VN.t1 VTAIL.t0 w_n2114_n1078# sky130_fd_pr__pfet_01v8 ad=0.09075 pd=0.88 as=0.2145 ps=1.88 w=0.55 l=1.1
X4 VDD1.t4 VP.t1 VTAIL.t11 w_n2114_n1078# sky130_fd_pr__pfet_01v8 ad=0.09075 pd=0.88 as=0.2145 ps=1.88 w=0.55 l=1.1
X5 VDD2.t3 VN.t2 VTAIL.t1 w_n2114_n1078# sky130_fd_pr__pfet_01v8 ad=0.2145 pd=1.88 as=0.09075 ps=0.88 w=0.55 l=1.1
X6 VDD1.t3 VP.t2 VTAIL.t6 w_n2114_n1078# sky130_fd_pr__pfet_01v8 ad=0.2145 pd=1.88 as=0.09075 ps=0.88 w=0.55 l=1.1
X7 VDD2.t2 VN.t3 VTAIL.t2 w_n2114_n1078# sky130_fd_pr__pfet_01v8 ad=0.09075 pd=0.88 as=0.2145 ps=1.88 w=0.55 l=1.1
X8 VTAIL.t10 VP.t3 VDD1.t2 w_n2114_n1078# sky130_fd_pr__pfet_01v8 ad=0.09075 pd=0.88 as=0.09075 ps=0.88 w=0.55 l=1.1
X9 VTAIL.t3 VN.t4 VDD2.t1 w_n2114_n1078# sky130_fd_pr__pfet_01v8 ad=0.09075 pd=0.88 as=0.09075 ps=0.88 w=0.55 l=1.1
X10 VDD1.t1 VP.t4 VTAIL.t9 w_n2114_n1078# sky130_fd_pr__pfet_01v8 ad=0.09075 pd=0.88 as=0.2145 ps=1.88 w=0.55 l=1.1
X11 B.t8 B.t6 B.t7 w_n2114_n1078# sky130_fd_pr__pfet_01v8 ad=0.2145 pd=1.88 as=0 ps=0 w=0.55 l=1.1
X12 VDD2.t0 VN.t5 VTAIL.t4 w_n2114_n1078# sky130_fd_pr__pfet_01v8 ad=0.2145 pd=1.88 as=0.09075 ps=0.88 w=0.55 l=1.1
X13 B.t5 B.t3 B.t4 w_n2114_n1078# sky130_fd_pr__pfet_01v8 ad=0.2145 pd=1.88 as=0 ps=0 w=0.55 l=1.1
X14 VTAIL.t8 VP.t5 VDD1.t0 w_n2114_n1078# sky130_fd_pr__pfet_01v8 ad=0.09075 pd=0.88 as=0.09075 ps=0.88 w=0.55 l=1.1
X15 B.t2 B.t0 B.t1 w_n2114_n1078# sky130_fd_pr__pfet_01v8 ad=0.2145 pd=1.88 as=0 ps=0 w=0.55 l=1.1
R0 VP.n5 VP.n2 161.3
R1 VP.n13 VP.n0 161.3
R2 VP.n12 VP.n11 161.3
R3 VP.n10 VP.n1 161.3
R4 VP.n7 VP.n6 80.6037
R5 VP.n15 VP.n14 80.6037
R6 VP.n9 VP.n8 80.6037
R7 VP.n3 VP.t2 71.0394
R8 VP.n8 VP.n1 50.6472
R9 VP.n14 VP.n13 50.6472
R10 VP.n6 VP.n5 50.6472
R11 VP.n8 VP.t0 47.9814
R12 VP.n14 VP.t1 47.9814
R13 VP.n6 VP.t4 47.9814
R14 VP.n9 VP.n7 34.3082
R15 VP.n4 VP.n3 32.6873
R16 VP.n3 VP.n2 28.1202
R17 VP.n12 VP.n1 24.4675
R18 VP.n13 VP.n12 24.4675
R19 VP.n5 VP.n4 24.4675
R20 VP.n12 VP.t3 12.0505
R21 VP.n4 VP.t5 12.0505
R22 VP.n7 VP.n2 0.285035
R23 VP.n10 VP.n9 0.285035
R24 VP.n15 VP.n0 0.285035
R25 VP.n11 VP.n10 0.189894
R26 VP.n11 VP.n0 0.189894
R27 VP VP.n15 0.146778
R28 VTAIL.n11 VTAIL.t0 675.316
R29 VTAIL.n2 VTAIL.t11 675.316
R30 VTAIL.n10 VTAIL.t9 675.316
R31 VTAIL.n7 VTAIL.t2 675.316
R32 VTAIL.n1 VTAIL.n0 616.216
R33 VTAIL.n4 VTAIL.n3 616.216
R34 VTAIL.n9 VTAIL.n8 616.216
R35 VTAIL.n6 VTAIL.n5 616.216
R36 VTAIL.n0 VTAIL.t1 59.1005
R37 VTAIL.n0 VTAIL.t3 59.1005
R38 VTAIL.n3 VTAIL.t7 59.1005
R39 VTAIL.n3 VTAIL.t10 59.1005
R40 VTAIL.n8 VTAIL.t6 59.1005
R41 VTAIL.n8 VTAIL.t8 59.1005
R42 VTAIL.n5 VTAIL.t4 59.1005
R43 VTAIL.n5 VTAIL.t5 59.1005
R44 VTAIL.n6 VTAIL.n4 15.3065
R45 VTAIL.n11 VTAIL.n10 14.0738
R46 VTAIL.n7 VTAIL.n6 1.23326
R47 VTAIL.n10 VTAIL.n9 1.23326
R48 VTAIL.n4 VTAIL.n2 1.23326
R49 VTAIL.n9 VTAIL.n7 1.08671
R50 VTAIL.n2 VTAIL.n1 1.08671
R51 VTAIL VTAIL.n11 0.866879
R52 VTAIL VTAIL.n1 0.366879
R53 VDD1 VDD1.t3 692.977
R54 VDD1.n1 VDD1.t5 692.864
R55 VDD1.n1 VDD1.n0 633.148
R56 VDD1.n3 VDD1.n2 632.894
R57 VDD1.n2 VDD1.t0 59.1005
R58 VDD1.n2 VDD1.t1 59.1005
R59 VDD1.n0 VDD1.t2 59.1005
R60 VDD1.n0 VDD1.t4 59.1005
R61 VDD1.n3 VDD1.n1 29.3953
R62 VDD1 VDD1.n3 0.2505
R63 B.n145 B.t5 692.197
R64 B.n67 B.t11 692.197
R65 B.n20 B.t7 692.197
R66 B.n27 B.t1 692.197
R67 B.n146 B.t4 664.465
R68 B.n68 B.t10 664.465
R69 B.n21 B.t8 664.465
R70 B.n28 B.t2 664.465
R71 B.n239 B.n238 585
R72 B.n240 B.n31 585
R73 B.n242 B.n241 585
R74 B.n243 B.n30 585
R75 B.n245 B.n244 585
R76 B.n246 B.n29 585
R77 B.n248 B.n247 585
R78 B.n249 B.n26 585
R79 B.n252 B.n251 585
R80 B.n253 B.n25 585
R81 B.n255 B.n254 585
R82 B.n256 B.n24 585
R83 B.n258 B.n257 585
R84 B.n259 B.n23 585
R85 B.n261 B.n260 585
R86 B.n262 B.n19 585
R87 B.n264 B.n263 585
R88 B.n265 B.n18 585
R89 B.n267 B.n266 585
R90 B.n268 B.n17 585
R91 B.n270 B.n269 585
R92 B.n271 B.n16 585
R93 B.n273 B.n272 585
R94 B.n274 B.n15 585
R95 B.n276 B.n275 585
R96 B.n237 B.n32 585
R97 B.n236 B.n235 585
R98 B.n234 B.n33 585
R99 B.n233 B.n232 585
R100 B.n231 B.n34 585
R101 B.n230 B.n229 585
R102 B.n228 B.n35 585
R103 B.n227 B.n226 585
R104 B.n225 B.n36 585
R105 B.n224 B.n223 585
R106 B.n222 B.n37 585
R107 B.n221 B.n220 585
R108 B.n219 B.n38 585
R109 B.n218 B.n217 585
R110 B.n216 B.n39 585
R111 B.n215 B.n214 585
R112 B.n213 B.n40 585
R113 B.n212 B.n211 585
R114 B.n210 B.n41 585
R115 B.n209 B.n208 585
R116 B.n207 B.n42 585
R117 B.n206 B.n205 585
R118 B.n204 B.n43 585
R119 B.n203 B.n202 585
R120 B.n201 B.n44 585
R121 B.n200 B.n199 585
R122 B.n198 B.n45 585
R123 B.n197 B.n196 585
R124 B.n195 B.n46 585
R125 B.n194 B.n193 585
R126 B.n192 B.n47 585
R127 B.n191 B.n190 585
R128 B.n189 B.n48 585
R129 B.n188 B.n187 585
R130 B.n186 B.n49 585
R131 B.n185 B.n184 585
R132 B.n183 B.n50 585
R133 B.n182 B.n181 585
R134 B.n180 B.n51 585
R135 B.n179 B.n178 585
R136 B.n177 B.n52 585
R137 B.n176 B.n175 585
R138 B.n174 B.n53 585
R139 B.n173 B.n172 585
R140 B.n171 B.n54 585
R141 B.n170 B.n169 585
R142 B.n168 B.n55 585
R143 B.n167 B.n166 585
R144 B.n165 B.n56 585
R145 B.n164 B.n163 585
R146 B.n162 B.n57 585
R147 B.n121 B.n120 585
R148 B.n122 B.n71 585
R149 B.n124 B.n123 585
R150 B.n125 B.n70 585
R151 B.n127 B.n126 585
R152 B.n128 B.n69 585
R153 B.n130 B.n129 585
R154 B.n131 B.n66 585
R155 B.n134 B.n133 585
R156 B.n135 B.n65 585
R157 B.n137 B.n136 585
R158 B.n138 B.n64 585
R159 B.n140 B.n139 585
R160 B.n141 B.n63 585
R161 B.n143 B.n142 585
R162 B.n144 B.n62 585
R163 B.n149 B.n148 585
R164 B.n150 B.n61 585
R165 B.n152 B.n151 585
R166 B.n153 B.n60 585
R167 B.n155 B.n154 585
R168 B.n156 B.n59 585
R169 B.n158 B.n157 585
R170 B.n159 B.n58 585
R171 B.n161 B.n160 585
R172 B.n119 B.n72 585
R173 B.n118 B.n117 585
R174 B.n116 B.n73 585
R175 B.n115 B.n114 585
R176 B.n113 B.n74 585
R177 B.n112 B.n111 585
R178 B.n110 B.n75 585
R179 B.n109 B.n108 585
R180 B.n107 B.n76 585
R181 B.n106 B.n105 585
R182 B.n104 B.n77 585
R183 B.n103 B.n102 585
R184 B.n101 B.n78 585
R185 B.n100 B.n99 585
R186 B.n98 B.n79 585
R187 B.n97 B.n96 585
R188 B.n95 B.n80 585
R189 B.n94 B.n93 585
R190 B.n92 B.n81 585
R191 B.n91 B.n90 585
R192 B.n89 B.n82 585
R193 B.n88 B.n87 585
R194 B.n86 B.n83 585
R195 B.n85 B.n84 585
R196 B.n2 B.n0 585
R197 B.n313 B.n1 585
R198 B.n312 B.n311 585
R199 B.n310 B.n3 585
R200 B.n309 B.n308 585
R201 B.n307 B.n4 585
R202 B.n306 B.n305 585
R203 B.n304 B.n5 585
R204 B.n303 B.n302 585
R205 B.n301 B.n6 585
R206 B.n300 B.n299 585
R207 B.n298 B.n7 585
R208 B.n297 B.n296 585
R209 B.n295 B.n8 585
R210 B.n294 B.n293 585
R211 B.n292 B.n9 585
R212 B.n291 B.n290 585
R213 B.n289 B.n10 585
R214 B.n288 B.n287 585
R215 B.n286 B.n11 585
R216 B.n285 B.n284 585
R217 B.n283 B.n12 585
R218 B.n282 B.n281 585
R219 B.n280 B.n13 585
R220 B.n279 B.n278 585
R221 B.n277 B.n14 585
R222 B.n315 B.n314 585
R223 B.n121 B.n72 526.135
R224 B.n277 B.n276 526.135
R225 B.n162 B.n161 526.135
R226 B.n239 B.n32 526.135
R227 B.n145 B.t3 206.263
R228 B.n67 B.t9 206.263
R229 B.n20 B.t6 206.263
R230 B.n27 B.t0 206.263
R231 B.n117 B.n72 163.367
R232 B.n117 B.n116 163.367
R233 B.n116 B.n115 163.367
R234 B.n115 B.n74 163.367
R235 B.n111 B.n74 163.367
R236 B.n111 B.n110 163.367
R237 B.n110 B.n109 163.367
R238 B.n109 B.n76 163.367
R239 B.n105 B.n76 163.367
R240 B.n105 B.n104 163.367
R241 B.n104 B.n103 163.367
R242 B.n103 B.n78 163.367
R243 B.n99 B.n78 163.367
R244 B.n99 B.n98 163.367
R245 B.n98 B.n97 163.367
R246 B.n97 B.n80 163.367
R247 B.n93 B.n80 163.367
R248 B.n93 B.n92 163.367
R249 B.n92 B.n91 163.367
R250 B.n91 B.n82 163.367
R251 B.n87 B.n82 163.367
R252 B.n87 B.n86 163.367
R253 B.n86 B.n85 163.367
R254 B.n85 B.n2 163.367
R255 B.n314 B.n2 163.367
R256 B.n314 B.n313 163.367
R257 B.n313 B.n312 163.367
R258 B.n312 B.n3 163.367
R259 B.n308 B.n3 163.367
R260 B.n308 B.n307 163.367
R261 B.n307 B.n306 163.367
R262 B.n306 B.n5 163.367
R263 B.n302 B.n5 163.367
R264 B.n302 B.n301 163.367
R265 B.n301 B.n300 163.367
R266 B.n300 B.n7 163.367
R267 B.n296 B.n7 163.367
R268 B.n296 B.n295 163.367
R269 B.n295 B.n294 163.367
R270 B.n294 B.n9 163.367
R271 B.n290 B.n9 163.367
R272 B.n290 B.n289 163.367
R273 B.n289 B.n288 163.367
R274 B.n288 B.n11 163.367
R275 B.n284 B.n11 163.367
R276 B.n284 B.n283 163.367
R277 B.n283 B.n282 163.367
R278 B.n282 B.n13 163.367
R279 B.n278 B.n13 163.367
R280 B.n278 B.n277 163.367
R281 B.n122 B.n121 163.367
R282 B.n123 B.n122 163.367
R283 B.n123 B.n70 163.367
R284 B.n127 B.n70 163.367
R285 B.n128 B.n127 163.367
R286 B.n129 B.n128 163.367
R287 B.n129 B.n66 163.367
R288 B.n134 B.n66 163.367
R289 B.n135 B.n134 163.367
R290 B.n136 B.n135 163.367
R291 B.n136 B.n64 163.367
R292 B.n140 B.n64 163.367
R293 B.n141 B.n140 163.367
R294 B.n142 B.n141 163.367
R295 B.n142 B.n62 163.367
R296 B.n149 B.n62 163.367
R297 B.n150 B.n149 163.367
R298 B.n151 B.n150 163.367
R299 B.n151 B.n60 163.367
R300 B.n155 B.n60 163.367
R301 B.n156 B.n155 163.367
R302 B.n157 B.n156 163.367
R303 B.n157 B.n58 163.367
R304 B.n161 B.n58 163.367
R305 B.n163 B.n162 163.367
R306 B.n163 B.n56 163.367
R307 B.n167 B.n56 163.367
R308 B.n168 B.n167 163.367
R309 B.n169 B.n168 163.367
R310 B.n169 B.n54 163.367
R311 B.n173 B.n54 163.367
R312 B.n174 B.n173 163.367
R313 B.n175 B.n174 163.367
R314 B.n175 B.n52 163.367
R315 B.n179 B.n52 163.367
R316 B.n180 B.n179 163.367
R317 B.n181 B.n180 163.367
R318 B.n181 B.n50 163.367
R319 B.n185 B.n50 163.367
R320 B.n186 B.n185 163.367
R321 B.n187 B.n186 163.367
R322 B.n187 B.n48 163.367
R323 B.n191 B.n48 163.367
R324 B.n192 B.n191 163.367
R325 B.n193 B.n192 163.367
R326 B.n193 B.n46 163.367
R327 B.n197 B.n46 163.367
R328 B.n198 B.n197 163.367
R329 B.n199 B.n198 163.367
R330 B.n199 B.n44 163.367
R331 B.n203 B.n44 163.367
R332 B.n204 B.n203 163.367
R333 B.n205 B.n204 163.367
R334 B.n205 B.n42 163.367
R335 B.n209 B.n42 163.367
R336 B.n210 B.n209 163.367
R337 B.n211 B.n210 163.367
R338 B.n211 B.n40 163.367
R339 B.n215 B.n40 163.367
R340 B.n216 B.n215 163.367
R341 B.n217 B.n216 163.367
R342 B.n217 B.n38 163.367
R343 B.n221 B.n38 163.367
R344 B.n222 B.n221 163.367
R345 B.n223 B.n222 163.367
R346 B.n223 B.n36 163.367
R347 B.n227 B.n36 163.367
R348 B.n228 B.n227 163.367
R349 B.n229 B.n228 163.367
R350 B.n229 B.n34 163.367
R351 B.n233 B.n34 163.367
R352 B.n234 B.n233 163.367
R353 B.n235 B.n234 163.367
R354 B.n235 B.n32 163.367
R355 B.n276 B.n15 163.367
R356 B.n272 B.n15 163.367
R357 B.n272 B.n271 163.367
R358 B.n271 B.n270 163.367
R359 B.n270 B.n17 163.367
R360 B.n266 B.n17 163.367
R361 B.n266 B.n265 163.367
R362 B.n265 B.n264 163.367
R363 B.n264 B.n19 163.367
R364 B.n260 B.n19 163.367
R365 B.n260 B.n259 163.367
R366 B.n259 B.n258 163.367
R367 B.n258 B.n24 163.367
R368 B.n254 B.n24 163.367
R369 B.n254 B.n253 163.367
R370 B.n253 B.n252 163.367
R371 B.n252 B.n26 163.367
R372 B.n247 B.n26 163.367
R373 B.n247 B.n246 163.367
R374 B.n246 B.n245 163.367
R375 B.n245 B.n30 163.367
R376 B.n241 B.n30 163.367
R377 B.n241 B.n240 163.367
R378 B.n240 B.n239 163.367
R379 B.n147 B.n146 59.5399
R380 B.n132 B.n68 59.5399
R381 B.n22 B.n21 59.5399
R382 B.n250 B.n28 59.5399
R383 B.n275 B.n14 34.1859
R384 B.n238 B.n237 34.1859
R385 B.n160 B.n57 34.1859
R386 B.n120 B.n119 34.1859
R387 B.n146 B.n145 27.7338
R388 B.n68 B.n67 27.7338
R389 B.n21 B.n20 27.7338
R390 B.n28 B.n27 27.7338
R391 B B.n315 18.0485
R392 B.n275 B.n274 10.6151
R393 B.n274 B.n273 10.6151
R394 B.n273 B.n16 10.6151
R395 B.n269 B.n16 10.6151
R396 B.n269 B.n268 10.6151
R397 B.n268 B.n267 10.6151
R398 B.n267 B.n18 10.6151
R399 B.n263 B.n262 10.6151
R400 B.n262 B.n261 10.6151
R401 B.n261 B.n23 10.6151
R402 B.n257 B.n23 10.6151
R403 B.n257 B.n256 10.6151
R404 B.n256 B.n255 10.6151
R405 B.n255 B.n25 10.6151
R406 B.n251 B.n25 10.6151
R407 B.n249 B.n248 10.6151
R408 B.n248 B.n29 10.6151
R409 B.n244 B.n29 10.6151
R410 B.n244 B.n243 10.6151
R411 B.n243 B.n242 10.6151
R412 B.n242 B.n31 10.6151
R413 B.n238 B.n31 10.6151
R414 B.n164 B.n57 10.6151
R415 B.n165 B.n164 10.6151
R416 B.n166 B.n165 10.6151
R417 B.n166 B.n55 10.6151
R418 B.n170 B.n55 10.6151
R419 B.n171 B.n170 10.6151
R420 B.n172 B.n171 10.6151
R421 B.n172 B.n53 10.6151
R422 B.n176 B.n53 10.6151
R423 B.n177 B.n176 10.6151
R424 B.n178 B.n177 10.6151
R425 B.n178 B.n51 10.6151
R426 B.n182 B.n51 10.6151
R427 B.n183 B.n182 10.6151
R428 B.n184 B.n183 10.6151
R429 B.n184 B.n49 10.6151
R430 B.n188 B.n49 10.6151
R431 B.n189 B.n188 10.6151
R432 B.n190 B.n189 10.6151
R433 B.n190 B.n47 10.6151
R434 B.n194 B.n47 10.6151
R435 B.n195 B.n194 10.6151
R436 B.n196 B.n195 10.6151
R437 B.n196 B.n45 10.6151
R438 B.n200 B.n45 10.6151
R439 B.n201 B.n200 10.6151
R440 B.n202 B.n201 10.6151
R441 B.n202 B.n43 10.6151
R442 B.n206 B.n43 10.6151
R443 B.n207 B.n206 10.6151
R444 B.n208 B.n207 10.6151
R445 B.n208 B.n41 10.6151
R446 B.n212 B.n41 10.6151
R447 B.n213 B.n212 10.6151
R448 B.n214 B.n213 10.6151
R449 B.n214 B.n39 10.6151
R450 B.n218 B.n39 10.6151
R451 B.n219 B.n218 10.6151
R452 B.n220 B.n219 10.6151
R453 B.n220 B.n37 10.6151
R454 B.n224 B.n37 10.6151
R455 B.n225 B.n224 10.6151
R456 B.n226 B.n225 10.6151
R457 B.n226 B.n35 10.6151
R458 B.n230 B.n35 10.6151
R459 B.n231 B.n230 10.6151
R460 B.n232 B.n231 10.6151
R461 B.n232 B.n33 10.6151
R462 B.n236 B.n33 10.6151
R463 B.n237 B.n236 10.6151
R464 B.n120 B.n71 10.6151
R465 B.n124 B.n71 10.6151
R466 B.n125 B.n124 10.6151
R467 B.n126 B.n125 10.6151
R468 B.n126 B.n69 10.6151
R469 B.n130 B.n69 10.6151
R470 B.n131 B.n130 10.6151
R471 B.n133 B.n65 10.6151
R472 B.n137 B.n65 10.6151
R473 B.n138 B.n137 10.6151
R474 B.n139 B.n138 10.6151
R475 B.n139 B.n63 10.6151
R476 B.n143 B.n63 10.6151
R477 B.n144 B.n143 10.6151
R478 B.n148 B.n144 10.6151
R479 B.n152 B.n61 10.6151
R480 B.n153 B.n152 10.6151
R481 B.n154 B.n153 10.6151
R482 B.n154 B.n59 10.6151
R483 B.n158 B.n59 10.6151
R484 B.n159 B.n158 10.6151
R485 B.n160 B.n159 10.6151
R486 B.n119 B.n118 10.6151
R487 B.n118 B.n73 10.6151
R488 B.n114 B.n73 10.6151
R489 B.n114 B.n113 10.6151
R490 B.n113 B.n112 10.6151
R491 B.n112 B.n75 10.6151
R492 B.n108 B.n75 10.6151
R493 B.n108 B.n107 10.6151
R494 B.n107 B.n106 10.6151
R495 B.n106 B.n77 10.6151
R496 B.n102 B.n77 10.6151
R497 B.n102 B.n101 10.6151
R498 B.n101 B.n100 10.6151
R499 B.n100 B.n79 10.6151
R500 B.n96 B.n79 10.6151
R501 B.n96 B.n95 10.6151
R502 B.n95 B.n94 10.6151
R503 B.n94 B.n81 10.6151
R504 B.n90 B.n81 10.6151
R505 B.n90 B.n89 10.6151
R506 B.n89 B.n88 10.6151
R507 B.n88 B.n83 10.6151
R508 B.n84 B.n83 10.6151
R509 B.n84 B.n0 10.6151
R510 B.n311 B.n1 10.6151
R511 B.n311 B.n310 10.6151
R512 B.n310 B.n309 10.6151
R513 B.n309 B.n4 10.6151
R514 B.n305 B.n4 10.6151
R515 B.n305 B.n304 10.6151
R516 B.n304 B.n303 10.6151
R517 B.n303 B.n6 10.6151
R518 B.n299 B.n6 10.6151
R519 B.n299 B.n298 10.6151
R520 B.n298 B.n297 10.6151
R521 B.n297 B.n8 10.6151
R522 B.n293 B.n8 10.6151
R523 B.n293 B.n292 10.6151
R524 B.n292 B.n291 10.6151
R525 B.n291 B.n10 10.6151
R526 B.n287 B.n10 10.6151
R527 B.n287 B.n286 10.6151
R528 B.n286 B.n285 10.6151
R529 B.n285 B.n12 10.6151
R530 B.n281 B.n12 10.6151
R531 B.n281 B.n280 10.6151
R532 B.n280 B.n279 10.6151
R533 B.n279 B.n14 10.6151
R534 B.n263 B.n22 6.5566
R535 B.n251 B.n250 6.5566
R536 B.n133 B.n132 6.5566
R537 B.n148 B.n147 6.5566
R538 B.n22 B.n18 4.05904
R539 B.n250 B.n249 4.05904
R540 B.n132 B.n131 4.05904
R541 B.n147 B.n61 4.05904
R542 B.n315 B.n0 2.81026
R543 B.n315 B.n1 2.81026
R544 VN.n9 VN.n6 161.3
R545 VN.n3 VN.n0 161.3
R546 VN.n11 VN.n10 80.6037
R547 VN.n5 VN.n4 80.6037
R548 VN.n1 VN.t2 71.0394
R549 VN.n7 VN.t3 71.0394
R550 VN.n4 VN.n3 50.6472
R551 VN.n10 VN.n9 50.6472
R552 VN.n4 VN.t1 47.9814
R553 VN.n10 VN.t5 47.9814
R554 VN VN.n11 34.5938
R555 VN.n2 VN.n1 32.6873
R556 VN.n8 VN.n7 32.6873
R557 VN.n7 VN.n6 28.1202
R558 VN.n1 VN.n0 28.1202
R559 VN.n3 VN.n2 24.4675
R560 VN.n9 VN.n8 24.4675
R561 VN.n2 VN.t4 12.0505
R562 VN.n8 VN.t0 12.0505
R563 VN.n11 VN.n6 0.285035
R564 VN.n5 VN.n0 0.285035
R565 VN VN.n5 0.146778
R566 VDD2.n1 VDD2.t3 692.864
R567 VDD2.n2 VDD2.t0 691.995
R568 VDD2.n1 VDD2.n0 633.148
R569 VDD2 VDD2.n3 633.144
R570 VDD2.n3 VDD2.t5 59.1005
R571 VDD2.n3 VDD2.t2 59.1005
R572 VDD2.n0 VDD2.t1 59.1005
R573 VDD2.n0 VDD2.t4 59.1005
R574 VDD2.n2 VDD2.n1 28.1959
R575 VDD2 VDD2.n2 0.983259
C0 VTAIL B 0.667824f
C1 VDD2 VP 0.340117f
C2 VDD1 VP 0.75982f
C3 VTAIL VP 1.0999f
C4 VN w_n2114_n1078# 3.37586f
C5 VN B 0.671562f
C6 w_n2114_n1078# B 4.40126f
C7 VDD2 VDD1 0.855366f
C8 VN VP 3.35732f
C9 VTAIL VDD2 2.51212f
C10 VP w_n2114_n1078# 3.63556f
C11 VTAIL VDD1 2.46889f
C12 VP B 1.11178f
C13 VN VDD2 0.579462f
C14 VDD2 w_n2114_n1078# 1.11246f
C15 VN VDD1 0.157318f
C16 VDD1 w_n2114_n1078# 1.0771f
C17 VTAIL VN 1.08578f
C18 VDD2 B 0.861436f
C19 VTAIL w_n2114_n1078# 1.07625f
C20 VDD1 B 0.822604f
C21 VDD2 VSUBS 0.615344f
C22 VDD1 VSUBS 0.886627f
C23 VTAIL VSUBS 0.315306f
C24 VN VSUBS 3.9748f
C25 VP VSUBS 1.267046f
C26 B VSUBS 2.071203f
C27 w_n2114_n1078# VSUBS 29.553698f
C28 VDD2.t3 VSUBS 0.041845f
C29 VDD2.t1 VSUBS 0.00904f
C30 VDD2.t4 VSUBS 0.00904f
C31 VDD2.n0 VSUBS 0.020147f
C32 VDD2.n1 VSUBS 1.04729f
C33 VDD2.t0 VSUBS 0.041687f
C34 VDD2.n2 VSUBS 1.0471f
C35 VDD2.t5 VSUBS 0.00904f
C36 VDD2.t2 VSUBS 0.00904f
C37 VDD2.n3 VSUBS 0.020146f
C38 VN.n0 VSUBS 0.359363f
C39 VN.t4 VSUBS 0.043104f
C40 VN.t2 VSUBS 0.224072f
C41 VN.n1 VSUBS 0.176756f
C42 VN.n2 VSUBS 0.202022f
C43 VN.n3 VSUBS 0.08498f
C44 VN.t1 VSUBS 0.151858f
C45 VN.n4 VSUBS 0.206073f
C46 VN.n5 VSUBS 0.060439f
C47 VN.n6 VSUBS 0.359363f
C48 VN.t0 VSUBS 0.043104f
C49 VN.t3 VSUBS 0.224072f
C50 VN.n7 VSUBS 0.176756f
C51 VN.n8 VSUBS 0.202022f
C52 VN.n9 VSUBS 0.08498f
C53 VN.t5 VSUBS 0.151858f
C54 VN.n10 VSUBS 0.206073f
C55 VN.n11 VSUBS 1.91024f
C56 B.n0 VSUBS 0.006854f
C57 B.n1 VSUBS 0.006854f
C58 B.n2 VSUBS 0.010838f
C59 B.n3 VSUBS 0.010838f
C60 B.n4 VSUBS 0.010838f
C61 B.n5 VSUBS 0.010838f
C62 B.n6 VSUBS 0.010838f
C63 B.n7 VSUBS 0.010838f
C64 B.n8 VSUBS 0.010838f
C65 B.n9 VSUBS 0.010838f
C66 B.n10 VSUBS 0.010838f
C67 B.n11 VSUBS 0.010838f
C68 B.n12 VSUBS 0.010838f
C69 B.n13 VSUBS 0.010838f
C70 B.n14 VSUBS 0.025856f
C71 B.n15 VSUBS 0.010838f
C72 B.n16 VSUBS 0.010838f
C73 B.n17 VSUBS 0.010838f
C74 B.n18 VSUBS 0.007491f
C75 B.n19 VSUBS 0.010838f
C76 B.t8 VSUBS 0.01593f
C77 B.t7 VSUBS 0.01732f
C78 B.t6 VSUBS 0.051755f
C79 B.n20 VSUBS 0.055386f
C80 B.n21 VSUBS 0.050138f
C81 B.n22 VSUBS 0.025111f
C82 B.n23 VSUBS 0.010838f
C83 B.n24 VSUBS 0.010838f
C84 B.n25 VSUBS 0.010838f
C85 B.n26 VSUBS 0.010838f
C86 B.t2 VSUBS 0.01593f
C87 B.t1 VSUBS 0.01732f
C88 B.t0 VSUBS 0.051755f
C89 B.n27 VSUBS 0.055386f
C90 B.n28 VSUBS 0.050138f
C91 B.n29 VSUBS 0.010838f
C92 B.n30 VSUBS 0.010838f
C93 B.n31 VSUBS 0.010838f
C94 B.n32 VSUBS 0.025856f
C95 B.n33 VSUBS 0.010838f
C96 B.n34 VSUBS 0.010838f
C97 B.n35 VSUBS 0.010838f
C98 B.n36 VSUBS 0.010838f
C99 B.n37 VSUBS 0.010838f
C100 B.n38 VSUBS 0.010838f
C101 B.n39 VSUBS 0.010838f
C102 B.n40 VSUBS 0.010838f
C103 B.n41 VSUBS 0.010838f
C104 B.n42 VSUBS 0.010838f
C105 B.n43 VSUBS 0.010838f
C106 B.n44 VSUBS 0.010838f
C107 B.n45 VSUBS 0.010838f
C108 B.n46 VSUBS 0.010838f
C109 B.n47 VSUBS 0.010838f
C110 B.n48 VSUBS 0.010838f
C111 B.n49 VSUBS 0.010838f
C112 B.n50 VSUBS 0.010838f
C113 B.n51 VSUBS 0.010838f
C114 B.n52 VSUBS 0.010838f
C115 B.n53 VSUBS 0.010838f
C116 B.n54 VSUBS 0.010838f
C117 B.n55 VSUBS 0.010838f
C118 B.n56 VSUBS 0.010838f
C119 B.n57 VSUBS 0.025856f
C120 B.n58 VSUBS 0.010838f
C121 B.n59 VSUBS 0.010838f
C122 B.n60 VSUBS 0.010838f
C123 B.n61 VSUBS 0.007491f
C124 B.n62 VSUBS 0.010838f
C125 B.n63 VSUBS 0.010838f
C126 B.n64 VSUBS 0.010838f
C127 B.n65 VSUBS 0.010838f
C128 B.n66 VSUBS 0.010838f
C129 B.t10 VSUBS 0.01593f
C130 B.t11 VSUBS 0.01732f
C131 B.t9 VSUBS 0.051755f
C132 B.n67 VSUBS 0.055386f
C133 B.n68 VSUBS 0.050138f
C134 B.n69 VSUBS 0.010838f
C135 B.n70 VSUBS 0.010838f
C136 B.n71 VSUBS 0.010838f
C137 B.n72 VSUBS 0.025856f
C138 B.n73 VSUBS 0.010838f
C139 B.n74 VSUBS 0.010838f
C140 B.n75 VSUBS 0.010838f
C141 B.n76 VSUBS 0.010838f
C142 B.n77 VSUBS 0.010838f
C143 B.n78 VSUBS 0.010838f
C144 B.n79 VSUBS 0.010838f
C145 B.n80 VSUBS 0.010838f
C146 B.n81 VSUBS 0.010838f
C147 B.n82 VSUBS 0.010838f
C148 B.n83 VSUBS 0.010838f
C149 B.n84 VSUBS 0.010838f
C150 B.n85 VSUBS 0.010838f
C151 B.n86 VSUBS 0.010838f
C152 B.n87 VSUBS 0.010838f
C153 B.n88 VSUBS 0.010838f
C154 B.n89 VSUBS 0.010838f
C155 B.n90 VSUBS 0.010838f
C156 B.n91 VSUBS 0.010838f
C157 B.n92 VSUBS 0.010838f
C158 B.n93 VSUBS 0.010838f
C159 B.n94 VSUBS 0.010838f
C160 B.n95 VSUBS 0.010838f
C161 B.n96 VSUBS 0.010838f
C162 B.n97 VSUBS 0.010838f
C163 B.n98 VSUBS 0.010838f
C164 B.n99 VSUBS 0.010838f
C165 B.n100 VSUBS 0.010838f
C166 B.n101 VSUBS 0.010838f
C167 B.n102 VSUBS 0.010838f
C168 B.n103 VSUBS 0.010838f
C169 B.n104 VSUBS 0.010838f
C170 B.n105 VSUBS 0.010838f
C171 B.n106 VSUBS 0.010838f
C172 B.n107 VSUBS 0.010838f
C173 B.n108 VSUBS 0.010838f
C174 B.n109 VSUBS 0.010838f
C175 B.n110 VSUBS 0.010838f
C176 B.n111 VSUBS 0.010838f
C177 B.n112 VSUBS 0.010838f
C178 B.n113 VSUBS 0.010838f
C179 B.n114 VSUBS 0.010838f
C180 B.n115 VSUBS 0.010838f
C181 B.n116 VSUBS 0.010838f
C182 B.n117 VSUBS 0.010838f
C183 B.n118 VSUBS 0.010838f
C184 B.n119 VSUBS 0.025856f
C185 B.n120 VSUBS 0.026423f
C186 B.n121 VSUBS 0.026423f
C187 B.n122 VSUBS 0.010838f
C188 B.n123 VSUBS 0.010838f
C189 B.n124 VSUBS 0.010838f
C190 B.n125 VSUBS 0.010838f
C191 B.n126 VSUBS 0.010838f
C192 B.n127 VSUBS 0.010838f
C193 B.n128 VSUBS 0.010838f
C194 B.n129 VSUBS 0.010838f
C195 B.n130 VSUBS 0.010838f
C196 B.n131 VSUBS 0.007491f
C197 B.n132 VSUBS 0.025111f
C198 B.n133 VSUBS 0.008766f
C199 B.n134 VSUBS 0.010838f
C200 B.n135 VSUBS 0.010838f
C201 B.n136 VSUBS 0.010838f
C202 B.n137 VSUBS 0.010838f
C203 B.n138 VSUBS 0.010838f
C204 B.n139 VSUBS 0.010838f
C205 B.n140 VSUBS 0.010838f
C206 B.n141 VSUBS 0.010838f
C207 B.n142 VSUBS 0.010838f
C208 B.n143 VSUBS 0.010838f
C209 B.n144 VSUBS 0.010838f
C210 B.t4 VSUBS 0.01593f
C211 B.t5 VSUBS 0.01732f
C212 B.t3 VSUBS 0.051755f
C213 B.n145 VSUBS 0.055386f
C214 B.n146 VSUBS 0.050138f
C215 B.n147 VSUBS 0.025111f
C216 B.n148 VSUBS 0.008766f
C217 B.n149 VSUBS 0.010838f
C218 B.n150 VSUBS 0.010838f
C219 B.n151 VSUBS 0.010838f
C220 B.n152 VSUBS 0.010838f
C221 B.n153 VSUBS 0.010838f
C222 B.n154 VSUBS 0.010838f
C223 B.n155 VSUBS 0.010838f
C224 B.n156 VSUBS 0.010838f
C225 B.n157 VSUBS 0.010838f
C226 B.n158 VSUBS 0.010838f
C227 B.n159 VSUBS 0.010838f
C228 B.n160 VSUBS 0.026423f
C229 B.n161 VSUBS 0.026423f
C230 B.n162 VSUBS 0.025856f
C231 B.n163 VSUBS 0.010838f
C232 B.n164 VSUBS 0.010838f
C233 B.n165 VSUBS 0.010838f
C234 B.n166 VSUBS 0.010838f
C235 B.n167 VSUBS 0.010838f
C236 B.n168 VSUBS 0.010838f
C237 B.n169 VSUBS 0.010838f
C238 B.n170 VSUBS 0.010838f
C239 B.n171 VSUBS 0.010838f
C240 B.n172 VSUBS 0.010838f
C241 B.n173 VSUBS 0.010838f
C242 B.n174 VSUBS 0.010838f
C243 B.n175 VSUBS 0.010838f
C244 B.n176 VSUBS 0.010838f
C245 B.n177 VSUBS 0.010838f
C246 B.n178 VSUBS 0.010838f
C247 B.n179 VSUBS 0.010838f
C248 B.n180 VSUBS 0.010838f
C249 B.n181 VSUBS 0.010838f
C250 B.n182 VSUBS 0.010838f
C251 B.n183 VSUBS 0.010838f
C252 B.n184 VSUBS 0.010838f
C253 B.n185 VSUBS 0.010838f
C254 B.n186 VSUBS 0.010838f
C255 B.n187 VSUBS 0.010838f
C256 B.n188 VSUBS 0.010838f
C257 B.n189 VSUBS 0.010838f
C258 B.n190 VSUBS 0.010838f
C259 B.n191 VSUBS 0.010838f
C260 B.n192 VSUBS 0.010838f
C261 B.n193 VSUBS 0.010838f
C262 B.n194 VSUBS 0.010838f
C263 B.n195 VSUBS 0.010838f
C264 B.n196 VSUBS 0.010838f
C265 B.n197 VSUBS 0.010838f
C266 B.n198 VSUBS 0.010838f
C267 B.n199 VSUBS 0.010838f
C268 B.n200 VSUBS 0.010838f
C269 B.n201 VSUBS 0.010838f
C270 B.n202 VSUBS 0.010838f
C271 B.n203 VSUBS 0.010838f
C272 B.n204 VSUBS 0.010838f
C273 B.n205 VSUBS 0.010838f
C274 B.n206 VSUBS 0.010838f
C275 B.n207 VSUBS 0.010838f
C276 B.n208 VSUBS 0.010838f
C277 B.n209 VSUBS 0.010838f
C278 B.n210 VSUBS 0.010838f
C279 B.n211 VSUBS 0.010838f
C280 B.n212 VSUBS 0.010838f
C281 B.n213 VSUBS 0.010838f
C282 B.n214 VSUBS 0.010838f
C283 B.n215 VSUBS 0.010838f
C284 B.n216 VSUBS 0.010838f
C285 B.n217 VSUBS 0.010838f
C286 B.n218 VSUBS 0.010838f
C287 B.n219 VSUBS 0.010838f
C288 B.n220 VSUBS 0.010838f
C289 B.n221 VSUBS 0.010838f
C290 B.n222 VSUBS 0.010838f
C291 B.n223 VSUBS 0.010838f
C292 B.n224 VSUBS 0.010838f
C293 B.n225 VSUBS 0.010838f
C294 B.n226 VSUBS 0.010838f
C295 B.n227 VSUBS 0.010838f
C296 B.n228 VSUBS 0.010838f
C297 B.n229 VSUBS 0.010838f
C298 B.n230 VSUBS 0.010838f
C299 B.n231 VSUBS 0.010838f
C300 B.n232 VSUBS 0.010838f
C301 B.n233 VSUBS 0.010838f
C302 B.n234 VSUBS 0.010838f
C303 B.n235 VSUBS 0.010838f
C304 B.n236 VSUBS 0.010838f
C305 B.n237 VSUBS 0.02708f
C306 B.n238 VSUBS 0.0252f
C307 B.n239 VSUBS 0.026423f
C308 B.n240 VSUBS 0.010838f
C309 B.n241 VSUBS 0.010838f
C310 B.n242 VSUBS 0.010838f
C311 B.n243 VSUBS 0.010838f
C312 B.n244 VSUBS 0.010838f
C313 B.n245 VSUBS 0.010838f
C314 B.n246 VSUBS 0.010838f
C315 B.n247 VSUBS 0.010838f
C316 B.n248 VSUBS 0.010838f
C317 B.n249 VSUBS 0.007491f
C318 B.n250 VSUBS 0.025111f
C319 B.n251 VSUBS 0.008766f
C320 B.n252 VSUBS 0.010838f
C321 B.n253 VSUBS 0.010838f
C322 B.n254 VSUBS 0.010838f
C323 B.n255 VSUBS 0.010838f
C324 B.n256 VSUBS 0.010838f
C325 B.n257 VSUBS 0.010838f
C326 B.n258 VSUBS 0.010838f
C327 B.n259 VSUBS 0.010838f
C328 B.n260 VSUBS 0.010838f
C329 B.n261 VSUBS 0.010838f
C330 B.n262 VSUBS 0.010838f
C331 B.n263 VSUBS 0.008766f
C332 B.n264 VSUBS 0.010838f
C333 B.n265 VSUBS 0.010838f
C334 B.n266 VSUBS 0.010838f
C335 B.n267 VSUBS 0.010838f
C336 B.n268 VSUBS 0.010838f
C337 B.n269 VSUBS 0.010838f
C338 B.n270 VSUBS 0.010838f
C339 B.n271 VSUBS 0.010838f
C340 B.n272 VSUBS 0.010838f
C341 B.n273 VSUBS 0.010838f
C342 B.n274 VSUBS 0.010838f
C343 B.n275 VSUBS 0.026423f
C344 B.n276 VSUBS 0.026423f
C345 B.n277 VSUBS 0.025856f
C346 B.n278 VSUBS 0.010838f
C347 B.n279 VSUBS 0.010838f
C348 B.n280 VSUBS 0.010838f
C349 B.n281 VSUBS 0.010838f
C350 B.n282 VSUBS 0.010838f
C351 B.n283 VSUBS 0.010838f
C352 B.n284 VSUBS 0.010838f
C353 B.n285 VSUBS 0.010838f
C354 B.n286 VSUBS 0.010838f
C355 B.n287 VSUBS 0.010838f
C356 B.n288 VSUBS 0.010838f
C357 B.n289 VSUBS 0.010838f
C358 B.n290 VSUBS 0.010838f
C359 B.n291 VSUBS 0.010838f
C360 B.n292 VSUBS 0.010838f
C361 B.n293 VSUBS 0.010838f
C362 B.n294 VSUBS 0.010838f
C363 B.n295 VSUBS 0.010838f
C364 B.n296 VSUBS 0.010838f
C365 B.n297 VSUBS 0.010838f
C366 B.n298 VSUBS 0.010838f
C367 B.n299 VSUBS 0.010838f
C368 B.n300 VSUBS 0.010838f
C369 B.n301 VSUBS 0.010838f
C370 B.n302 VSUBS 0.010838f
C371 B.n303 VSUBS 0.010838f
C372 B.n304 VSUBS 0.010838f
C373 B.n305 VSUBS 0.010838f
C374 B.n306 VSUBS 0.010838f
C375 B.n307 VSUBS 0.010838f
C376 B.n308 VSUBS 0.010838f
C377 B.n309 VSUBS 0.010838f
C378 B.n310 VSUBS 0.010838f
C379 B.n311 VSUBS 0.010838f
C380 B.n312 VSUBS 0.010838f
C381 B.n313 VSUBS 0.010838f
C382 B.n314 VSUBS 0.010838f
C383 B.n315 VSUBS 0.024542f
C384 VDD1.t3 VSUBS 0.040627f
C385 VDD1.t5 VSUBS 0.040597f
C386 VDD1.t2 VSUBS 0.008771f
C387 VDD1.t4 VSUBS 0.008771f
C388 VDD1.n0 VSUBS 0.019547f
C389 VDD1.n1 VSUBS 1.07932f
C390 VDD1.t0 VSUBS 0.008771f
C391 VDD1.t1 VSUBS 0.008771f
C392 VDD1.n2 VSUBS 0.019483f
C393 VDD1.n3 VSUBS 1.05673f
C394 VTAIL.t1 VSUBS 0.013895f
C395 VTAIL.t3 VSUBS 0.013895f
C396 VTAIL.n0 VSUBS 0.02873f
C397 VTAIL.n1 VSUBS 0.193327f
C398 VTAIL.t11 VSUBS 0.06201f
C399 VTAIL.n2 VSUBS 0.287191f
C400 VTAIL.t7 VSUBS 0.013895f
C401 VTAIL.t10 VSUBS 0.013895f
C402 VTAIL.n3 VSUBS 0.02873f
C403 VTAIL.n4 VSUBS 0.907775f
C404 VTAIL.t4 VSUBS 0.013895f
C405 VTAIL.t5 VSUBS 0.013895f
C406 VTAIL.n5 VSUBS 0.02873f
C407 VTAIL.n6 VSUBS 0.907775f
C408 VTAIL.t2 VSUBS 0.06201f
C409 VTAIL.n7 VSUBS 0.287191f
C410 VTAIL.t6 VSUBS 0.013895f
C411 VTAIL.t8 VSUBS 0.013895f
C412 VTAIL.n8 VSUBS 0.02873f
C413 VTAIL.n9 VSUBS 0.282576f
C414 VTAIL.t9 VSUBS 0.06201f
C415 VTAIL.n10 VSUBS 0.785399f
C416 VTAIL.t0 VSUBS 0.06201f
C417 VTAIL.n11 VSUBS 0.747657f
C418 VP.n0 VSUBS 0.089844f
C419 VP.t3 VSUBS 0.044972f
C420 VP.n1 VSUBS 0.088662f
C421 VP.n2 VSUBS 0.374934f
C422 VP.t4 VSUBS 0.158438f
C423 VP.t5 VSUBS 0.044972f
C424 VP.t2 VSUBS 0.233781f
C425 VP.n3 VSUBS 0.184415f
C426 VP.n4 VSUBS 0.210776f
C427 VP.n5 VSUBS 0.088662f
C428 VP.n6 VSUBS 0.215003f
C429 VP.n7 VSUBS 1.95374f
C430 VP.t0 VSUBS 0.158438f
C431 VP.n8 VSUBS 0.215003f
C432 VP.n9 VSUBS 2.02429f
C433 VP.n10 VSUBS 0.089844f
C434 VP.n11 VSUBS 0.067331f
C435 VP.n12 VSUBS 0.16354f
C436 VP.n13 VSUBS 0.088662f
C437 VP.t1 VSUBS 0.158438f
C438 VP.n14 VSUBS 0.215003f
C439 VP.n15 VSUBS 0.063058f
.ends

