* NGSPICE file created from diff_pair_sample_1485.ext - technology: sky130A

.subckt diff_pair_sample_1485 VTAIL VN VP B VDD2 VDD1
X0 B.t23 B.t21 B.t22 B.t11 sky130_fd_pr__nfet_01v8 ad=2.3361 pd=12.76 as=0 ps=0 w=5.99 l=0.59
X1 B.t20 B.t18 B.t19 B.t15 sky130_fd_pr__nfet_01v8 ad=2.3361 pd=12.76 as=0 ps=0 w=5.99 l=0.59
X2 VTAIL.t17 VP.t0 VDD1.t1 B.t5 sky130_fd_pr__nfet_01v8 ad=0.98835 pd=6.32 as=0.98835 ps=6.32 w=5.99 l=0.59
X3 VTAIL.t2 VN.t0 VDD2.t9 B.t1 sky130_fd_pr__nfet_01v8 ad=0.98835 pd=6.32 as=0.98835 ps=6.32 w=5.99 l=0.59
X4 VTAIL.t1 VN.t1 VDD2.t8 B.t5 sky130_fd_pr__nfet_01v8 ad=0.98835 pd=6.32 as=0.98835 ps=6.32 w=5.99 l=0.59
X5 VTAIL.t3 VN.t2 VDD2.t7 B.t0 sky130_fd_pr__nfet_01v8 ad=0.98835 pd=6.32 as=0.98835 ps=6.32 w=5.99 l=0.59
X6 VTAIL.t5 VN.t3 VDD2.t6 B.t4 sky130_fd_pr__nfet_01v8 ad=0.98835 pd=6.32 as=0.98835 ps=6.32 w=5.99 l=0.59
X7 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=2.3361 pd=12.76 as=0 ps=0 w=5.99 l=0.59
X8 VDD2.t5 VN.t4 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=0.98835 pd=6.32 as=0.98835 ps=6.32 w=5.99 l=0.59
X9 VDD1.t2 VP.t1 VTAIL.t16 B.t3 sky130_fd_pr__nfet_01v8 ad=2.3361 pd=12.76 as=0.98835 ps=6.32 w=5.99 l=0.59
X10 VDD2.t4 VN.t5 VTAIL.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=2.3361 pd=12.76 as=0.98835 ps=6.32 w=5.99 l=0.59
X11 VDD1.t3 VP.t2 VTAIL.t15 B.t8 sky130_fd_pr__nfet_01v8 ad=0.98835 pd=6.32 as=2.3361 ps=12.76 w=5.99 l=0.59
X12 VTAIL.t14 VP.t3 VDD1.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=0.98835 pd=6.32 as=0.98835 ps=6.32 w=5.99 l=0.59
X13 VDD1.t5 VP.t4 VTAIL.t13 B.t7 sky130_fd_pr__nfet_01v8 ad=0.98835 pd=6.32 as=0.98835 ps=6.32 w=5.99 l=0.59
X14 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=2.3361 pd=12.76 as=0 ps=0 w=5.99 l=0.59
X15 VDD2.t3 VN.t6 VTAIL.t18 B.t9 sky130_fd_pr__nfet_01v8 ad=0.98835 pd=6.32 as=2.3361 ps=12.76 w=5.99 l=0.59
X16 VDD1.t6 VP.t5 VTAIL.t12 B.t6 sky130_fd_pr__nfet_01v8 ad=2.3361 pd=12.76 as=0.98835 ps=6.32 w=5.99 l=0.59
X17 VDD1.t8 VP.t6 VTAIL.t11 B.t2 sky130_fd_pr__nfet_01v8 ad=0.98835 pd=6.32 as=0.98835 ps=6.32 w=5.99 l=0.59
X18 VDD2.t2 VN.t7 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=2.3361 pd=12.76 as=0.98835 ps=6.32 w=5.99 l=0.59
X19 VDD1.t7 VP.t7 VTAIL.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=0.98835 pd=6.32 as=2.3361 ps=12.76 w=5.99 l=0.59
X20 VDD2.t1 VN.t8 VTAIL.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=0.98835 pd=6.32 as=0.98835 ps=6.32 w=5.99 l=0.59
X21 VTAIL.t9 VP.t8 VDD1.t9 B.t0 sky130_fd_pr__nfet_01v8 ad=0.98835 pd=6.32 as=0.98835 ps=6.32 w=5.99 l=0.59
X22 VTAIL.t8 VP.t9 VDD1.t0 B.t4 sky130_fd_pr__nfet_01v8 ad=0.98835 pd=6.32 as=0.98835 ps=6.32 w=5.99 l=0.59
X23 VDD2.t0 VN.t9 VTAIL.t19 B.t8 sky130_fd_pr__nfet_01v8 ad=0.98835 pd=6.32 as=2.3361 ps=12.76 w=5.99 l=0.59
R0 B.n493 B.n492 585
R1 B.n494 B.n493 585
R2 B.n192 B.n77 585
R3 B.n191 B.n190 585
R4 B.n189 B.n188 585
R5 B.n187 B.n186 585
R6 B.n185 B.n184 585
R7 B.n183 B.n182 585
R8 B.n181 B.n180 585
R9 B.n179 B.n178 585
R10 B.n177 B.n176 585
R11 B.n175 B.n174 585
R12 B.n173 B.n172 585
R13 B.n171 B.n170 585
R14 B.n169 B.n168 585
R15 B.n167 B.n166 585
R16 B.n165 B.n164 585
R17 B.n163 B.n162 585
R18 B.n161 B.n160 585
R19 B.n159 B.n158 585
R20 B.n157 B.n156 585
R21 B.n155 B.n154 585
R22 B.n153 B.n152 585
R23 B.n151 B.n150 585
R24 B.n149 B.n148 585
R25 B.n146 B.n145 585
R26 B.n144 B.n143 585
R27 B.n142 B.n141 585
R28 B.n140 B.n139 585
R29 B.n138 B.n137 585
R30 B.n136 B.n135 585
R31 B.n134 B.n133 585
R32 B.n132 B.n131 585
R33 B.n130 B.n129 585
R34 B.n128 B.n127 585
R35 B.n126 B.n125 585
R36 B.n124 B.n123 585
R37 B.n122 B.n121 585
R38 B.n120 B.n119 585
R39 B.n118 B.n117 585
R40 B.n116 B.n115 585
R41 B.n114 B.n113 585
R42 B.n112 B.n111 585
R43 B.n110 B.n109 585
R44 B.n108 B.n107 585
R45 B.n106 B.n105 585
R46 B.n104 B.n103 585
R47 B.n102 B.n101 585
R48 B.n100 B.n99 585
R49 B.n98 B.n97 585
R50 B.n96 B.n95 585
R51 B.n94 B.n93 585
R52 B.n92 B.n91 585
R53 B.n90 B.n89 585
R54 B.n88 B.n87 585
R55 B.n86 B.n85 585
R56 B.n84 B.n83 585
R57 B.n47 B.n46 585
R58 B.n491 B.n48 585
R59 B.n495 B.n48 585
R60 B.n490 B.n489 585
R61 B.n489 B.n44 585
R62 B.n488 B.n43 585
R63 B.n501 B.n43 585
R64 B.n487 B.n42 585
R65 B.n502 B.n42 585
R66 B.n486 B.n41 585
R67 B.n503 B.n41 585
R68 B.n485 B.n484 585
R69 B.n484 B.n37 585
R70 B.n483 B.n36 585
R71 B.n509 B.n36 585
R72 B.n482 B.n35 585
R73 B.n510 B.n35 585
R74 B.n481 B.n34 585
R75 B.n511 B.n34 585
R76 B.n480 B.n479 585
R77 B.n479 B.n30 585
R78 B.n478 B.n29 585
R79 B.n517 B.n29 585
R80 B.n477 B.n28 585
R81 B.n518 B.n28 585
R82 B.n476 B.n27 585
R83 B.n519 B.n27 585
R84 B.n475 B.n474 585
R85 B.n474 B.n26 585
R86 B.n473 B.n22 585
R87 B.n525 B.n22 585
R88 B.n472 B.n21 585
R89 B.n526 B.n21 585
R90 B.n471 B.n20 585
R91 B.n527 B.n20 585
R92 B.n470 B.n469 585
R93 B.n469 B.n16 585
R94 B.n468 B.n15 585
R95 B.n533 B.n15 585
R96 B.n467 B.n14 585
R97 B.n534 B.n14 585
R98 B.n466 B.n13 585
R99 B.n535 B.n13 585
R100 B.n465 B.n464 585
R101 B.n464 B.n12 585
R102 B.n463 B.n462 585
R103 B.n463 B.n8 585
R104 B.n461 B.n7 585
R105 B.n542 B.n7 585
R106 B.n460 B.n6 585
R107 B.n543 B.n6 585
R108 B.n459 B.n5 585
R109 B.n544 B.n5 585
R110 B.n458 B.n457 585
R111 B.n457 B.n4 585
R112 B.n456 B.n193 585
R113 B.n456 B.n455 585
R114 B.n445 B.n194 585
R115 B.n448 B.n194 585
R116 B.n447 B.n446 585
R117 B.n449 B.n447 585
R118 B.n444 B.n199 585
R119 B.n199 B.n198 585
R120 B.n443 B.n442 585
R121 B.n442 B.n441 585
R122 B.n201 B.n200 585
R123 B.n202 B.n201 585
R124 B.n434 B.n433 585
R125 B.n435 B.n434 585
R126 B.n432 B.n207 585
R127 B.n207 B.n206 585
R128 B.n431 B.n430 585
R129 B.n430 B.n429 585
R130 B.n209 B.n208 585
R131 B.n422 B.n209 585
R132 B.n421 B.n420 585
R133 B.n423 B.n421 585
R134 B.n419 B.n214 585
R135 B.n214 B.n213 585
R136 B.n418 B.n417 585
R137 B.n417 B.n416 585
R138 B.n216 B.n215 585
R139 B.n217 B.n216 585
R140 B.n409 B.n408 585
R141 B.n410 B.n409 585
R142 B.n407 B.n222 585
R143 B.n222 B.n221 585
R144 B.n406 B.n405 585
R145 B.n405 B.n404 585
R146 B.n224 B.n223 585
R147 B.n225 B.n224 585
R148 B.n397 B.n396 585
R149 B.n398 B.n397 585
R150 B.n395 B.n230 585
R151 B.n230 B.n229 585
R152 B.n394 B.n393 585
R153 B.n393 B.n392 585
R154 B.n232 B.n231 585
R155 B.n233 B.n232 585
R156 B.n385 B.n384 585
R157 B.n386 B.n385 585
R158 B.n236 B.n235 585
R159 B.n272 B.n270 585
R160 B.n273 B.n269 585
R161 B.n273 B.n237 585
R162 B.n276 B.n275 585
R163 B.n277 B.n268 585
R164 B.n279 B.n278 585
R165 B.n281 B.n267 585
R166 B.n284 B.n283 585
R167 B.n285 B.n266 585
R168 B.n287 B.n286 585
R169 B.n289 B.n265 585
R170 B.n292 B.n291 585
R171 B.n293 B.n264 585
R172 B.n295 B.n294 585
R173 B.n297 B.n263 585
R174 B.n300 B.n299 585
R175 B.n301 B.n262 585
R176 B.n303 B.n302 585
R177 B.n305 B.n261 585
R178 B.n308 B.n307 585
R179 B.n309 B.n260 585
R180 B.n311 B.n310 585
R181 B.n313 B.n259 585
R182 B.n316 B.n315 585
R183 B.n318 B.n256 585
R184 B.n320 B.n319 585
R185 B.n322 B.n255 585
R186 B.n325 B.n324 585
R187 B.n326 B.n254 585
R188 B.n328 B.n327 585
R189 B.n330 B.n253 585
R190 B.n333 B.n332 585
R191 B.n334 B.n250 585
R192 B.n337 B.n336 585
R193 B.n339 B.n249 585
R194 B.n342 B.n341 585
R195 B.n343 B.n248 585
R196 B.n345 B.n344 585
R197 B.n347 B.n247 585
R198 B.n350 B.n349 585
R199 B.n351 B.n246 585
R200 B.n353 B.n352 585
R201 B.n355 B.n245 585
R202 B.n358 B.n357 585
R203 B.n359 B.n244 585
R204 B.n361 B.n360 585
R205 B.n363 B.n243 585
R206 B.n366 B.n365 585
R207 B.n367 B.n242 585
R208 B.n369 B.n368 585
R209 B.n371 B.n241 585
R210 B.n374 B.n373 585
R211 B.n375 B.n240 585
R212 B.n377 B.n376 585
R213 B.n379 B.n239 585
R214 B.n382 B.n381 585
R215 B.n383 B.n238 585
R216 B.n388 B.n387 585
R217 B.n387 B.n386 585
R218 B.n389 B.n234 585
R219 B.n234 B.n233 585
R220 B.n391 B.n390 585
R221 B.n392 B.n391 585
R222 B.n228 B.n227 585
R223 B.n229 B.n228 585
R224 B.n400 B.n399 585
R225 B.n399 B.n398 585
R226 B.n401 B.n226 585
R227 B.n226 B.n225 585
R228 B.n403 B.n402 585
R229 B.n404 B.n403 585
R230 B.n220 B.n219 585
R231 B.n221 B.n220 585
R232 B.n412 B.n411 585
R233 B.n411 B.n410 585
R234 B.n413 B.n218 585
R235 B.n218 B.n217 585
R236 B.n415 B.n414 585
R237 B.n416 B.n415 585
R238 B.n212 B.n211 585
R239 B.n213 B.n212 585
R240 B.n425 B.n424 585
R241 B.n424 B.n423 585
R242 B.n426 B.n210 585
R243 B.n422 B.n210 585
R244 B.n428 B.n427 585
R245 B.n429 B.n428 585
R246 B.n205 B.n204 585
R247 B.n206 B.n205 585
R248 B.n437 B.n436 585
R249 B.n436 B.n435 585
R250 B.n438 B.n203 585
R251 B.n203 B.n202 585
R252 B.n440 B.n439 585
R253 B.n441 B.n440 585
R254 B.n197 B.n196 585
R255 B.n198 B.n197 585
R256 B.n451 B.n450 585
R257 B.n450 B.n449 585
R258 B.n452 B.n195 585
R259 B.n448 B.n195 585
R260 B.n454 B.n453 585
R261 B.n455 B.n454 585
R262 B.n3 B.n0 585
R263 B.n4 B.n3 585
R264 B.n541 B.n1 585
R265 B.n542 B.n541 585
R266 B.n540 B.n539 585
R267 B.n540 B.n8 585
R268 B.n538 B.n9 585
R269 B.n12 B.n9 585
R270 B.n537 B.n536 585
R271 B.n536 B.n535 585
R272 B.n11 B.n10 585
R273 B.n534 B.n11 585
R274 B.n532 B.n531 585
R275 B.n533 B.n532 585
R276 B.n530 B.n17 585
R277 B.n17 B.n16 585
R278 B.n529 B.n528 585
R279 B.n528 B.n527 585
R280 B.n19 B.n18 585
R281 B.n526 B.n19 585
R282 B.n524 B.n523 585
R283 B.n525 B.n524 585
R284 B.n522 B.n23 585
R285 B.n26 B.n23 585
R286 B.n521 B.n520 585
R287 B.n520 B.n519 585
R288 B.n25 B.n24 585
R289 B.n518 B.n25 585
R290 B.n516 B.n515 585
R291 B.n517 B.n516 585
R292 B.n514 B.n31 585
R293 B.n31 B.n30 585
R294 B.n513 B.n512 585
R295 B.n512 B.n511 585
R296 B.n33 B.n32 585
R297 B.n510 B.n33 585
R298 B.n508 B.n507 585
R299 B.n509 B.n508 585
R300 B.n506 B.n38 585
R301 B.n38 B.n37 585
R302 B.n505 B.n504 585
R303 B.n504 B.n503 585
R304 B.n40 B.n39 585
R305 B.n502 B.n40 585
R306 B.n500 B.n499 585
R307 B.n501 B.n500 585
R308 B.n498 B.n45 585
R309 B.n45 B.n44 585
R310 B.n497 B.n496 585
R311 B.n496 B.n495 585
R312 B.n545 B.n544 585
R313 B.n543 B.n2 585
R314 B.n496 B.n47 511.721
R315 B.n493 B.n48 511.721
R316 B.n385 B.n238 511.721
R317 B.n387 B.n236 511.721
R318 B.n80 B.t10 449.247
R319 B.n78 B.t21 449.247
R320 B.n251 B.t14 449.247
R321 B.n257 B.t18 449.247
R322 B.n494 B.n76 256.663
R323 B.n494 B.n75 256.663
R324 B.n494 B.n74 256.663
R325 B.n494 B.n73 256.663
R326 B.n494 B.n72 256.663
R327 B.n494 B.n71 256.663
R328 B.n494 B.n70 256.663
R329 B.n494 B.n69 256.663
R330 B.n494 B.n68 256.663
R331 B.n494 B.n67 256.663
R332 B.n494 B.n66 256.663
R333 B.n494 B.n65 256.663
R334 B.n494 B.n64 256.663
R335 B.n494 B.n63 256.663
R336 B.n494 B.n62 256.663
R337 B.n494 B.n61 256.663
R338 B.n494 B.n60 256.663
R339 B.n494 B.n59 256.663
R340 B.n494 B.n58 256.663
R341 B.n494 B.n57 256.663
R342 B.n494 B.n56 256.663
R343 B.n494 B.n55 256.663
R344 B.n494 B.n54 256.663
R345 B.n494 B.n53 256.663
R346 B.n494 B.n52 256.663
R347 B.n494 B.n51 256.663
R348 B.n494 B.n50 256.663
R349 B.n494 B.n49 256.663
R350 B.n271 B.n237 256.663
R351 B.n274 B.n237 256.663
R352 B.n280 B.n237 256.663
R353 B.n282 B.n237 256.663
R354 B.n288 B.n237 256.663
R355 B.n290 B.n237 256.663
R356 B.n296 B.n237 256.663
R357 B.n298 B.n237 256.663
R358 B.n304 B.n237 256.663
R359 B.n306 B.n237 256.663
R360 B.n312 B.n237 256.663
R361 B.n314 B.n237 256.663
R362 B.n321 B.n237 256.663
R363 B.n323 B.n237 256.663
R364 B.n329 B.n237 256.663
R365 B.n331 B.n237 256.663
R366 B.n338 B.n237 256.663
R367 B.n340 B.n237 256.663
R368 B.n346 B.n237 256.663
R369 B.n348 B.n237 256.663
R370 B.n354 B.n237 256.663
R371 B.n356 B.n237 256.663
R372 B.n362 B.n237 256.663
R373 B.n364 B.n237 256.663
R374 B.n370 B.n237 256.663
R375 B.n372 B.n237 256.663
R376 B.n378 B.n237 256.663
R377 B.n380 B.n237 256.663
R378 B.n547 B.n546 256.663
R379 B.n78 B.t22 196.636
R380 B.n251 B.t17 196.636
R381 B.n80 B.t12 196.636
R382 B.n257 B.t20 196.636
R383 B.n79 B.t23 178.792
R384 B.n252 B.t16 178.792
R385 B.n81 B.t13 178.792
R386 B.n258 B.t19 178.792
R387 B.n85 B.n84 163.367
R388 B.n89 B.n88 163.367
R389 B.n93 B.n92 163.367
R390 B.n97 B.n96 163.367
R391 B.n101 B.n100 163.367
R392 B.n105 B.n104 163.367
R393 B.n109 B.n108 163.367
R394 B.n113 B.n112 163.367
R395 B.n117 B.n116 163.367
R396 B.n121 B.n120 163.367
R397 B.n125 B.n124 163.367
R398 B.n129 B.n128 163.367
R399 B.n133 B.n132 163.367
R400 B.n137 B.n136 163.367
R401 B.n141 B.n140 163.367
R402 B.n145 B.n144 163.367
R403 B.n150 B.n149 163.367
R404 B.n154 B.n153 163.367
R405 B.n158 B.n157 163.367
R406 B.n162 B.n161 163.367
R407 B.n166 B.n165 163.367
R408 B.n170 B.n169 163.367
R409 B.n174 B.n173 163.367
R410 B.n178 B.n177 163.367
R411 B.n182 B.n181 163.367
R412 B.n186 B.n185 163.367
R413 B.n190 B.n189 163.367
R414 B.n493 B.n77 163.367
R415 B.n385 B.n232 163.367
R416 B.n393 B.n232 163.367
R417 B.n393 B.n230 163.367
R418 B.n397 B.n230 163.367
R419 B.n397 B.n224 163.367
R420 B.n405 B.n224 163.367
R421 B.n405 B.n222 163.367
R422 B.n409 B.n222 163.367
R423 B.n409 B.n216 163.367
R424 B.n417 B.n216 163.367
R425 B.n417 B.n214 163.367
R426 B.n421 B.n214 163.367
R427 B.n421 B.n209 163.367
R428 B.n430 B.n209 163.367
R429 B.n430 B.n207 163.367
R430 B.n434 B.n207 163.367
R431 B.n434 B.n201 163.367
R432 B.n442 B.n201 163.367
R433 B.n442 B.n199 163.367
R434 B.n447 B.n199 163.367
R435 B.n447 B.n194 163.367
R436 B.n456 B.n194 163.367
R437 B.n457 B.n456 163.367
R438 B.n457 B.n5 163.367
R439 B.n6 B.n5 163.367
R440 B.n7 B.n6 163.367
R441 B.n463 B.n7 163.367
R442 B.n464 B.n463 163.367
R443 B.n464 B.n13 163.367
R444 B.n14 B.n13 163.367
R445 B.n15 B.n14 163.367
R446 B.n469 B.n15 163.367
R447 B.n469 B.n20 163.367
R448 B.n21 B.n20 163.367
R449 B.n22 B.n21 163.367
R450 B.n474 B.n22 163.367
R451 B.n474 B.n27 163.367
R452 B.n28 B.n27 163.367
R453 B.n29 B.n28 163.367
R454 B.n479 B.n29 163.367
R455 B.n479 B.n34 163.367
R456 B.n35 B.n34 163.367
R457 B.n36 B.n35 163.367
R458 B.n484 B.n36 163.367
R459 B.n484 B.n41 163.367
R460 B.n42 B.n41 163.367
R461 B.n43 B.n42 163.367
R462 B.n489 B.n43 163.367
R463 B.n489 B.n48 163.367
R464 B.n273 B.n272 163.367
R465 B.n275 B.n273 163.367
R466 B.n279 B.n268 163.367
R467 B.n283 B.n281 163.367
R468 B.n287 B.n266 163.367
R469 B.n291 B.n289 163.367
R470 B.n295 B.n264 163.367
R471 B.n299 B.n297 163.367
R472 B.n303 B.n262 163.367
R473 B.n307 B.n305 163.367
R474 B.n311 B.n260 163.367
R475 B.n315 B.n313 163.367
R476 B.n320 B.n256 163.367
R477 B.n324 B.n322 163.367
R478 B.n328 B.n254 163.367
R479 B.n332 B.n330 163.367
R480 B.n337 B.n250 163.367
R481 B.n341 B.n339 163.367
R482 B.n345 B.n248 163.367
R483 B.n349 B.n347 163.367
R484 B.n353 B.n246 163.367
R485 B.n357 B.n355 163.367
R486 B.n361 B.n244 163.367
R487 B.n365 B.n363 163.367
R488 B.n369 B.n242 163.367
R489 B.n373 B.n371 163.367
R490 B.n377 B.n240 163.367
R491 B.n381 B.n379 163.367
R492 B.n387 B.n234 163.367
R493 B.n391 B.n234 163.367
R494 B.n391 B.n228 163.367
R495 B.n399 B.n228 163.367
R496 B.n399 B.n226 163.367
R497 B.n403 B.n226 163.367
R498 B.n403 B.n220 163.367
R499 B.n411 B.n220 163.367
R500 B.n411 B.n218 163.367
R501 B.n415 B.n218 163.367
R502 B.n415 B.n212 163.367
R503 B.n424 B.n212 163.367
R504 B.n424 B.n210 163.367
R505 B.n428 B.n210 163.367
R506 B.n428 B.n205 163.367
R507 B.n436 B.n205 163.367
R508 B.n436 B.n203 163.367
R509 B.n440 B.n203 163.367
R510 B.n440 B.n197 163.367
R511 B.n450 B.n197 163.367
R512 B.n450 B.n195 163.367
R513 B.n454 B.n195 163.367
R514 B.n454 B.n3 163.367
R515 B.n545 B.n3 163.367
R516 B.n541 B.n2 163.367
R517 B.n541 B.n540 163.367
R518 B.n540 B.n9 163.367
R519 B.n536 B.n9 163.367
R520 B.n536 B.n11 163.367
R521 B.n532 B.n11 163.367
R522 B.n532 B.n17 163.367
R523 B.n528 B.n17 163.367
R524 B.n528 B.n19 163.367
R525 B.n524 B.n19 163.367
R526 B.n524 B.n23 163.367
R527 B.n520 B.n23 163.367
R528 B.n520 B.n25 163.367
R529 B.n516 B.n25 163.367
R530 B.n516 B.n31 163.367
R531 B.n512 B.n31 163.367
R532 B.n512 B.n33 163.367
R533 B.n508 B.n33 163.367
R534 B.n508 B.n38 163.367
R535 B.n504 B.n38 163.367
R536 B.n504 B.n40 163.367
R537 B.n500 B.n40 163.367
R538 B.n500 B.n45 163.367
R539 B.n496 B.n45 163.367
R540 B.n386 B.n237 110.343
R541 B.n495 B.n494 110.343
R542 B.n49 B.n47 71.676
R543 B.n85 B.n50 71.676
R544 B.n89 B.n51 71.676
R545 B.n93 B.n52 71.676
R546 B.n97 B.n53 71.676
R547 B.n101 B.n54 71.676
R548 B.n105 B.n55 71.676
R549 B.n109 B.n56 71.676
R550 B.n113 B.n57 71.676
R551 B.n117 B.n58 71.676
R552 B.n121 B.n59 71.676
R553 B.n125 B.n60 71.676
R554 B.n129 B.n61 71.676
R555 B.n133 B.n62 71.676
R556 B.n137 B.n63 71.676
R557 B.n141 B.n64 71.676
R558 B.n145 B.n65 71.676
R559 B.n150 B.n66 71.676
R560 B.n154 B.n67 71.676
R561 B.n158 B.n68 71.676
R562 B.n162 B.n69 71.676
R563 B.n166 B.n70 71.676
R564 B.n170 B.n71 71.676
R565 B.n174 B.n72 71.676
R566 B.n178 B.n73 71.676
R567 B.n182 B.n74 71.676
R568 B.n186 B.n75 71.676
R569 B.n190 B.n76 71.676
R570 B.n77 B.n76 71.676
R571 B.n189 B.n75 71.676
R572 B.n185 B.n74 71.676
R573 B.n181 B.n73 71.676
R574 B.n177 B.n72 71.676
R575 B.n173 B.n71 71.676
R576 B.n169 B.n70 71.676
R577 B.n165 B.n69 71.676
R578 B.n161 B.n68 71.676
R579 B.n157 B.n67 71.676
R580 B.n153 B.n66 71.676
R581 B.n149 B.n65 71.676
R582 B.n144 B.n64 71.676
R583 B.n140 B.n63 71.676
R584 B.n136 B.n62 71.676
R585 B.n132 B.n61 71.676
R586 B.n128 B.n60 71.676
R587 B.n124 B.n59 71.676
R588 B.n120 B.n58 71.676
R589 B.n116 B.n57 71.676
R590 B.n112 B.n56 71.676
R591 B.n108 B.n55 71.676
R592 B.n104 B.n54 71.676
R593 B.n100 B.n53 71.676
R594 B.n96 B.n52 71.676
R595 B.n92 B.n51 71.676
R596 B.n88 B.n50 71.676
R597 B.n84 B.n49 71.676
R598 B.n271 B.n236 71.676
R599 B.n275 B.n274 71.676
R600 B.n280 B.n279 71.676
R601 B.n283 B.n282 71.676
R602 B.n288 B.n287 71.676
R603 B.n291 B.n290 71.676
R604 B.n296 B.n295 71.676
R605 B.n299 B.n298 71.676
R606 B.n304 B.n303 71.676
R607 B.n307 B.n306 71.676
R608 B.n312 B.n311 71.676
R609 B.n315 B.n314 71.676
R610 B.n321 B.n320 71.676
R611 B.n324 B.n323 71.676
R612 B.n329 B.n328 71.676
R613 B.n332 B.n331 71.676
R614 B.n338 B.n337 71.676
R615 B.n341 B.n340 71.676
R616 B.n346 B.n345 71.676
R617 B.n349 B.n348 71.676
R618 B.n354 B.n353 71.676
R619 B.n357 B.n356 71.676
R620 B.n362 B.n361 71.676
R621 B.n365 B.n364 71.676
R622 B.n370 B.n369 71.676
R623 B.n373 B.n372 71.676
R624 B.n378 B.n377 71.676
R625 B.n381 B.n380 71.676
R626 B.n272 B.n271 71.676
R627 B.n274 B.n268 71.676
R628 B.n281 B.n280 71.676
R629 B.n282 B.n266 71.676
R630 B.n289 B.n288 71.676
R631 B.n290 B.n264 71.676
R632 B.n297 B.n296 71.676
R633 B.n298 B.n262 71.676
R634 B.n305 B.n304 71.676
R635 B.n306 B.n260 71.676
R636 B.n313 B.n312 71.676
R637 B.n314 B.n256 71.676
R638 B.n322 B.n321 71.676
R639 B.n323 B.n254 71.676
R640 B.n330 B.n329 71.676
R641 B.n331 B.n250 71.676
R642 B.n339 B.n338 71.676
R643 B.n340 B.n248 71.676
R644 B.n347 B.n346 71.676
R645 B.n348 B.n246 71.676
R646 B.n355 B.n354 71.676
R647 B.n356 B.n244 71.676
R648 B.n363 B.n362 71.676
R649 B.n364 B.n242 71.676
R650 B.n371 B.n370 71.676
R651 B.n372 B.n240 71.676
R652 B.n379 B.n378 71.676
R653 B.n380 B.n238 71.676
R654 B.n546 B.n545 71.676
R655 B.n546 B.n2 71.676
R656 B.n386 B.n233 66.4009
R657 B.n392 B.n233 66.4009
R658 B.n392 B.n229 66.4009
R659 B.n398 B.n229 66.4009
R660 B.n404 B.n225 66.4009
R661 B.n404 B.n221 66.4009
R662 B.n410 B.n221 66.4009
R663 B.n410 B.n217 66.4009
R664 B.n416 B.n217 66.4009
R665 B.n423 B.n213 66.4009
R666 B.n423 B.n422 66.4009
R667 B.n429 B.n206 66.4009
R668 B.n435 B.n206 66.4009
R669 B.n441 B.n202 66.4009
R670 B.n449 B.n198 66.4009
R671 B.n449 B.n448 66.4009
R672 B.n455 B.n4 66.4009
R673 B.n544 B.n4 66.4009
R674 B.n544 B.n543 66.4009
R675 B.n543 B.n542 66.4009
R676 B.n542 B.n8 66.4009
R677 B.n535 B.n12 66.4009
R678 B.n535 B.n534 66.4009
R679 B.n533 B.n16 66.4009
R680 B.n527 B.n526 66.4009
R681 B.n526 B.n525 66.4009
R682 B.n519 B.n26 66.4009
R683 B.n519 B.n518 66.4009
R684 B.n517 B.n30 66.4009
R685 B.n511 B.n30 66.4009
R686 B.n511 B.n510 66.4009
R687 B.n510 B.n509 66.4009
R688 B.n509 B.n37 66.4009
R689 B.n503 B.n502 66.4009
R690 B.n502 B.n501 66.4009
R691 B.n501 B.n44 66.4009
R692 B.n495 B.n44 66.4009
R693 B.n82 B.n81 59.5399
R694 B.n147 B.n79 59.5399
R695 B.n335 B.n252 59.5399
R696 B.n317 B.n258 59.5399
R697 B.t2 B.n202 57.6126
R698 B.t7 B.n16 57.6126
R699 B.n441 B.t0 55.6596
R700 B.t4 B.n533 55.6596
R701 B.n398 B.t15 53.7067
R702 B.n503 B.t11 53.7067
R703 B.n416 B.t6 47.8478
R704 B.t8 B.n517 47.8478
R705 B.n429 B.t1 38.0831
R706 B.n525 B.t5 38.0831
R707 B.n448 B.t9 36.1301
R708 B.n12 B.t3 36.1301
R709 B.n388 B.n235 33.2493
R710 B.n384 B.n383 33.2493
R711 B.n492 B.n491 33.2493
R712 B.n497 B.n46 33.2493
R713 B.n455 B.t9 30.2713
R714 B.t3 B.n8 30.2713
R715 B.n422 B.t1 28.3183
R716 B.n26 B.t5 28.3183
R717 B.t6 B.n213 18.5535
R718 B.n518 B.t8 18.5535
R719 B B.n547 18.0485
R720 B.n81 B.n80 17.8429
R721 B.n79 B.n78 17.8429
R722 B.n252 B.n251 17.8429
R723 B.n258 B.n257 17.8429
R724 B.t15 B.n225 12.6947
R725 B.t11 B.n37 12.6947
R726 B.t0 B.n198 10.7417
R727 B.n534 B.t4 10.7417
R728 B.n389 B.n388 10.6151
R729 B.n390 B.n389 10.6151
R730 B.n390 B.n227 10.6151
R731 B.n400 B.n227 10.6151
R732 B.n401 B.n400 10.6151
R733 B.n402 B.n401 10.6151
R734 B.n402 B.n219 10.6151
R735 B.n412 B.n219 10.6151
R736 B.n413 B.n412 10.6151
R737 B.n414 B.n413 10.6151
R738 B.n414 B.n211 10.6151
R739 B.n425 B.n211 10.6151
R740 B.n426 B.n425 10.6151
R741 B.n427 B.n426 10.6151
R742 B.n427 B.n204 10.6151
R743 B.n437 B.n204 10.6151
R744 B.n438 B.n437 10.6151
R745 B.n439 B.n438 10.6151
R746 B.n439 B.n196 10.6151
R747 B.n451 B.n196 10.6151
R748 B.n452 B.n451 10.6151
R749 B.n453 B.n452 10.6151
R750 B.n453 B.n0 10.6151
R751 B.n270 B.n235 10.6151
R752 B.n270 B.n269 10.6151
R753 B.n276 B.n269 10.6151
R754 B.n277 B.n276 10.6151
R755 B.n278 B.n277 10.6151
R756 B.n278 B.n267 10.6151
R757 B.n284 B.n267 10.6151
R758 B.n285 B.n284 10.6151
R759 B.n286 B.n285 10.6151
R760 B.n286 B.n265 10.6151
R761 B.n292 B.n265 10.6151
R762 B.n293 B.n292 10.6151
R763 B.n294 B.n293 10.6151
R764 B.n294 B.n263 10.6151
R765 B.n300 B.n263 10.6151
R766 B.n301 B.n300 10.6151
R767 B.n302 B.n301 10.6151
R768 B.n302 B.n261 10.6151
R769 B.n308 B.n261 10.6151
R770 B.n309 B.n308 10.6151
R771 B.n310 B.n309 10.6151
R772 B.n310 B.n259 10.6151
R773 B.n316 B.n259 10.6151
R774 B.n319 B.n318 10.6151
R775 B.n319 B.n255 10.6151
R776 B.n325 B.n255 10.6151
R777 B.n326 B.n325 10.6151
R778 B.n327 B.n326 10.6151
R779 B.n327 B.n253 10.6151
R780 B.n333 B.n253 10.6151
R781 B.n334 B.n333 10.6151
R782 B.n336 B.n249 10.6151
R783 B.n342 B.n249 10.6151
R784 B.n343 B.n342 10.6151
R785 B.n344 B.n343 10.6151
R786 B.n344 B.n247 10.6151
R787 B.n350 B.n247 10.6151
R788 B.n351 B.n350 10.6151
R789 B.n352 B.n351 10.6151
R790 B.n352 B.n245 10.6151
R791 B.n358 B.n245 10.6151
R792 B.n359 B.n358 10.6151
R793 B.n360 B.n359 10.6151
R794 B.n360 B.n243 10.6151
R795 B.n366 B.n243 10.6151
R796 B.n367 B.n366 10.6151
R797 B.n368 B.n367 10.6151
R798 B.n368 B.n241 10.6151
R799 B.n374 B.n241 10.6151
R800 B.n375 B.n374 10.6151
R801 B.n376 B.n375 10.6151
R802 B.n376 B.n239 10.6151
R803 B.n382 B.n239 10.6151
R804 B.n383 B.n382 10.6151
R805 B.n384 B.n231 10.6151
R806 B.n394 B.n231 10.6151
R807 B.n395 B.n394 10.6151
R808 B.n396 B.n395 10.6151
R809 B.n396 B.n223 10.6151
R810 B.n406 B.n223 10.6151
R811 B.n407 B.n406 10.6151
R812 B.n408 B.n407 10.6151
R813 B.n408 B.n215 10.6151
R814 B.n418 B.n215 10.6151
R815 B.n419 B.n418 10.6151
R816 B.n420 B.n419 10.6151
R817 B.n420 B.n208 10.6151
R818 B.n431 B.n208 10.6151
R819 B.n432 B.n431 10.6151
R820 B.n433 B.n432 10.6151
R821 B.n433 B.n200 10.6151
R822 B.n443 B.n200 10.6151
R823 B.n444 B.n443 10.6151
R824 B.n446 B.n444 10.6151
R825 B.n446 B.n445 10.6151
R826 B.n445 B.n193 10.6151
R827 B.n458 B.n193 10.6151
R828 B.n459 B.n458 10.6151
R829 B.n460 B.n459 10.6151
R830 B.n461 B.n460 10.6151
R831 B.n462 B.n461 10.6151
R832 B.n465 B.n462 10.6151
R833 B.n466 B.n465 10.6151
R834 B.n467 B.n466 10.6151
R835 B.n468 B.n467 10.6151
R836 B.n470 B.n468 10.6151
R837 B.n471 B.n470 10.6151
R838 B.n472 B.n471 10.6151
R839 B.n473 B.n472 10.6151
R840 B.n475 B.n473 10.6151
R841 B.n476 B.n475 10.6151
R842 B.n477 B.n476 10.6151
R843 B.n478 B.n477 10.6151
R844 B.n480 B.n478 10.6151
R845 B.n481 B.n480 10.6151
R846 B.n482 B.n481 10.6151
R847 B.n483 B.n482 10.6151
R848 B.n485 B.n483 10.6151
R849 B.n486 B.n485 10.6151
R850 B.n487 B.n486 10.6151
R851 B.n488 B.n487 10.6151
R852 B.n490 B.n488 10.6151
R853 B.n491 B.n490 10.6151
R854 B.n539 B.n1 10.6151
R855 B.n539 B.n538 10.6151
R856 B.n538 B.n537 10.6151
R857 B.n537 B.n10 10.6151
R858 B.n531 B.n10 10.6151
R859 B.n531 B.n530 10.6151
R860 B.n530 B.n529 10.6151
R861 B.n529 B.n18 10.6151
R862 B.n523 B.n18 10.6151
R863 B.n523 B.n522 10.6151
R864 B.n522 B.n521 10.6151
R865 B.n521 B.n24 10.6151
R866 B.n515 B.n24 10.6151
R867 B.n515 B.n514 10.6151
R868 B.n514 B.n513 10.6151
R869 B.n513 B.n32 10.6151
R870 B.n507 B.n32 10.6151
R871 B.n507 B.n506 10.6151
R872 B.n506 B.n505 10.6151
R873 B.n505 B.n39 10.6151
R874 B.n499 B.n39 10.6151
R875 B.n499 B.n498 10.6151
R876 B.n498 B.n497 10.6151
R877 B.n83 B.n46 10.6151
R878 B.n86 B.n83 10.6151
R879 B.n87 B.n86 10.6151
R880 B.n90 B.n87 10.6151
R881 B.n91 B.n90 10.6151
R882 B.n94 B.n91 10.6151
R883 B.n95 B.n94 10.6151
R884 B.n98 B.n95 10.6151
R885 B.n99 B.n98 10.6151
R886 B.n102 B.n99 10.6151
R887 B.n103 B.n102 10.6151
R888 B.n106 B.n103 10.6151
R889 B.n107 B.n106 10.6151
R890 B.n110 B.n107 10.6151
R891 B.n111 B.n110 10.6151
R892 B.n114 B.n111 10.6151
R893 B.n115 B.n114 10.6151
R894 B.n118 B.n115 10.6151
R895 B.n119 B.n118 10.6151
R896 B.n122 B.n119 10.6151
R897 B.n123 B.n122 10.6151
R898 B.n126 B.n123 10.6151
R899 B.n127 B.n126 10.6151
R900 B.n131 B.n130 10.6151
R901 B.n134 B.n131 10.6151
R902 B.n135 B.n134 10.6151
R903 B.n138 B.n135 10.6151
R904 B.n139 B.n138 10.6151
R905 B.n142 B.n139 10.6151
R906 B.n143 B.n142 10.6151
R907 B.n146 B.n143 10.6151
R908 B.n151 B.n148 10.6151
R909 B.n152 B.n151 10.6151
R910 B.n155 B.n152 10.6151
R911 B.n156 B.n155 10.6151
R912 B.n159 B.n156 10.6151
R913 B.n160 B.n159 10.6151
R914 B.n163 B.n160 10.6151
R915 B.n164 B.n163 10.6151
R916 B.n167 B.n164 10.6151
R917 B.n168 B.n167 10.6151
R918 B.n171 B.n168 10.6151
R919 B.n172 B.n171 10.6151
R920 B.n175 B.n172 10.6151
R921 B.n176 B.n175 10.6151
R922 B.n179 B.n176 10.6151
R923 B.n180 B.n179 10.6151
R924 B.n183 B.n180 10.6151
R925 B.n184 B.n183 10.6151
R926 B.n187 B.n184 10.6151
R927 B.n188 B.n187 10.6151
R928 B.n191 B.n188 10.6151
R929 B.n192 B.n191 10.6151
R930 B.n492 B.n192 10.6151
R931 B.n435 B.t2 8.78878
R932 B.n527 B.t7 8.78878
R933 B.n547 B.n0 8.11757
R934 B.n547 B.n1 8.11757
R935 B.n318 B.n317 6.5566
R936 B.n335 B.n334 6.5566
R937 B.n130 B.n82 6.5566
R938 B.n147 B.n146 6.5566
R939 B.n317 B.n316 4.05904
R940 B.n336 B.n335 4.05904
R941 B.n127 B.n82 4.05904
R942 B.n148 B.n147 4.05904
R943 VP.n6 VP.t1 337.387
R944 VP.n14 VP.t5 311.666
R945 VP.n16 VP.t3 311.666
R946 VP.n1 VP.t6 311.666
R947 VP.n20 VP.t8 311.666
R948 VP.n22 VP.t7 311.666
R949 VP.n11 VP.t2 311.666
R950 VP.n9 VP.t0 311.666
R951 VP.n8 VP.t4 311.666
R952 VP.n7 VP.t9 311.666
R953 VP.n23 VP.n22 161.3
R954 VP.n9 VP.n4 161.3
R955 VP.n10 VP.n3 161.3
R956 VP.n12 VP.n11 161.3
R957 VP.n21 VP.n0 161.3
R958 VP.n20 VP.n19 161.3
R959 VP.n17 VP.n16 161.3
R960 VP.n15 VP.n2 161.3
R961 VP.n14 VP.n13 161.3
R962 VP.n8 VP.n5 80.6037
R963 VP.n18 VP.n1 80.6037
R964 VP.n16 VP.n1 48.2005
R965 VP.n20 VP.n1 48.2005
R966 VP.n9 VP.n8 48.2005
R967 VP.n8 VP.n7 48.2005
R968 VP.n6 VP.n5 45.1242
R969 VP.n15 VP.n14 43.0884
R970 VP.n22 VP.n21 43.0884
R971 VP.n11 VP.n10 43.0884
R972 VP.n13 VP.n12 37.6293
R973 VP.n7 VP.n6 15.1442
R974 VP.n16 VP.n15 5.11262
R975 VP.n21 VP.n20 5.11262
R976 VP.n10 VP.n9 5.11262
R977 VP.n5 VP.n4 0.285035
R978 VP.n18 VP.n17 0.285035
R979 VP.n19 VP.n18 0.285035
R980 VP.n4 VP.n3 0.189894
R981 VP.n12 VP.n3 0.189894
R982 VP.n13 VP.n2 0.189894
R983 VP.n17 VP.n2 0.189894
R984 VP.n19 VP.n0 0.189894
R985 VP.n23 VP.n0 0.189894
R986 VP VP.n23 0.0516364
R987 VDD1.n26 VDD1.n0 289.615
R988 VDD1.n59 VDD1.n33 289.615
R989 VDD1.n27 VDD1.n26 185
R990 VDD1.n25 VDD1.n24 185
R991 VDD1.n4 VDD1.n3 185
R992 VDD1.n19 VDD1.n18 185
R993 VDD1.n17 VDD1.n16 185
R994 VDD1.n8 VDD1.n7 185
R995 VDD1.n11 VDD1.n10 185
R996 VDD1.n44 VDD1.n43 185
R997 VDD1.n41 VDD1.n40 185
R998 VDD1.n50 VDD1.n49 185
R999 VDD1.n52 VDD1.n51 185
R1000 VDD1.n37 VDD1.n36 185
R1001 VDD1.n58 VDD1.n57 185
R1002 VDD1.n60 VDD1.n59 185
R1003 VDD1.t2 VDD1.n9 147.661
R1004 VDD1.t6 VDD1.n42 147.661
R1005 VDD1.n26 VDD1.n25 104.615
R1006 VDD1.n25 VDD1.n3 104.615
R1007 VDD1.n18 VDD1.n3 104.615
R1008 VDD1.n18 VDD1.n17 104.615
R1009 VDD1.n17 VDD1.n7 104.615
R1010 VDD1.n10 VDD1.n7 104.615
R1011 VDD1.n43 VDD1.n40 104.615
R1012 VDD1.n50 VDD1.n40 104.615
R1013 VDD1.n51 VDD1.n50 104.615
R1014 VDD1.n51 VDD1.n36 104.615
R1015 VDD1.n58 VDD1.n36 104.615
R1016 VDD1.n59 VDD1.n58 104.615
R1017 VDD1.n67 VDD1.n66 67.5362
R1018 VDD1.n32 VDD1.n31 66.9969
R1019 VDD1.n69 VDD1.n68 66.9967
R1020 VDD1.n65 VDD1.n64 66.9967
R1021 VDD1.n10 VDD1.t2 52.3082
R1022 VDD1.n43 VDD1.t6 52.3082
R1023 VDD1.n32 VDD1.n30 49.4633
R1024 VDD1.n65 VDD1.n63 49.4633
R1025 VDD1.n69 VDD1.n67 33.6259
R1026 VDD1.n11 VDD1.n9 15.6674
R1027 VDD1.n44 VDD1.n42 15.6674
R1028 VDD1.n12 VDD1.n8 12.8005
R1029 VDD1.n45 VDD1.n41 12.8005
R1030 VDD1.n16 VDD1.n15 12.0247
R1031 VDD1.n49 VDD1.n48 12.0247
R1032 VDD1.n19 VDD1.n6 11.249
R1033 VDD1.n52 VDD1.n39 11.249
R1034 VDD1.n20 VDD1.n4 10.4732
R1035 VDD1.n53 VDD1.n37 10.4732
R1036 VDD1.n24 VDD1.n23 9.69747
R1037 VDD1.n57 VDD1.n56 9.69747
R1038 VDD1.n30 VDD1.n29 9.45567
R1039 VDD1.n63 VDD1.n62 9.45567
R1040 VDD1.n29 VDD1.n28 9.3005
R1041 VDD1.n2 VDD1.n1 9.3005
R1042 VDD1.n23 VDD1.n22 9.3005
R1043 VDD1.n21 VDD1.n20 9.3005
R1044 VDD1.n6 VDD1.n5 9.3005
R1045 VDD1.n15 VDD1.n14 9.3005
R1046 VDD1.n13 VDD1.n12 9.3005
R1047 VDD1.n62 VDD1.n61 9.3005
R1048 VDD1.n35 VDD1.n34 9.3005
R1049 VDD1.n56 VDD1.n55 9.3005
R1050 VDD1.n54 VDD1.n53 9.3005
R1051 VDD1.n39 VDD1.n38 9.3005
R1052 VDD1.n48 VDD1.n47 9.3005
R1053 VDD1.n46 VDD1.n45 9.3005
R1054 VDD1.n27 VDD1.n2 8.92171
R1055 VDD1.n60 VDD1.n35 8.92171
R1056 VDD1.n28 VDD1.n0 8.14595
R1057 VDD1.n61 VDD1.n33 8.14595
R1058 VDD1.n30 VDD1.n0 5.81868
R1059 VDD1.n63 VDD1.n33 5.81868
R1060 VDD1.n28 VDD1.n27 5.04292
R1061 VDD1.n61 VDD1.n60 5.04292
R1062 VDD1.n13 VDD1.n9 4.38594
R1063 VDD1.n46 VDD1.n42 4.38594
R1064 VDD1.n24 VDD1.n2 4.26717
R1065 VDD1.n57 VDD1.n35 4.26717
R1066 VDD1.n23 VDD1.n4 3.49141
R1067 VDD1.n56 VDD1.n37 3.49141
R1068 VDD1.n68 VDD1.t1 3.30601
R1069 VDD1.n68 VDD1.t3 3.30601
R1070 VDD1.n31 VDD1.t0 3.30601
R1071 VDD1.n31 VDD1.t5 3.30601
R1072 VDD1.n66 VDD1.t9 3.30601
R1073 VDD1.n66 VDD1.t7 3.30601
R1074 VDD1.n64 VDD1.t4 3.30601
R1075 VDD1.n64 VDD1.t8 3.30601
R1076 VDD1.n20 VDD1.n19 2.71565
R1077 VDD1.n53 VDD1.n52 2.71565
R1078 VDD1.n16 VDD1.n6 1.93989
R1079 VDD1.n49 VDD1.n39 1.93989
R1080 VDD1.n15 VDD1.n8 1.16414
R1081 VDD1.n48 VDD1.n41 1.16414
R1082 VDD1 VDD1.n69 0.537138
R1083 VDD1.n12 VDD1.n11 0.388379
R1084 VDD1.n45 VDD1.n44 0.388379
R1085 VDD1 VDD1.n32 0.256966
R1086 VDD1.n29 VDD1.n1 0.155672
R1087 VDD1.n22 VDD1.n1 0.155672
R1088 VDD1.n22 VDD1.n21 0.155672
R1089 VDD1.n21 VDD1.n5 0.155672
R1090 VDD1.n14 VDD1.n5 0.155672
R1091 VDD1.n14 VDD1.n13 0.155672
R1092 VDD1.n47 VDD1.n46 0.155672
R1093 VDD1.n47 VDD1.n38 0.155672
R1094 VDD1.n54 VDD1.n38 0.155672
R1095 VDD1.n55 VDD1.n54 0.155672
R1096 VDD1.n55 VDD1.n34 0.155672
R1097 VDD1.n62 VDD1.n34 0.155672
R1098 VDD1.n67 VDD1.n65 0.14343
R1099 VTAIL.n136 VTAIL.n110 289.615
R1100 VTAIL.n28 VTAIL.n2 289.615
R1101 VTAIL.n104 VTAIL.n78 289.615
R1102 VTAIL.n68 VTAIL.n42 289.615
R1103 VTAIL.n121 VTAIL.n120 185
R1104 VTAIL.n118 VTAIL.n117 185
R1105 VTAIL.n127 VTAIL.n126 185
R1106 VTAIL.n129 VTAIL.n128 185
R1107 VTAIL.n114 VTAIL.n113 185
R1108 VTAIL.n135 VTAIL.n134 185
R1109 VTAIL.n137 VTAIL.n136 185
R1110 VTAIL.n13 VTAIL.n12 185
R1111 VTAIL.n10 VTAIL.n9 185
R1112 VTAIL.n19 VTAIL.n18 185
R1113 VTAIL.n21 VTAIL.n20 185
R1114 VTAIL.n6 VTAIL.n5 185
R1115 VTAIL.n27 VTAIL.n26 185
R1116 VTAIL.n29 VTAIL.n28 185
R1117 VTAIL.n105 VTAIL.n104 185
R1118 VTAIL.n103 VTAIL.n102 185
R1119 VTAIL.n82 VTAIL.n81 185
R1120 VTAIL.n97 VTAIL.n96 185
R1121 VTAIL.n95 VTAIL.n94 185
R1122 VTAIL.n86 VTAIL.n85 185
R1123 VTAIL.n89 VTAIL.n88 185
R1124 VTAIL.n69 VTAIL.n68 185
R1125 VTAIL.n67 VTAIL.n66 185
R1126 VTAIL.n46 VTAIL.n45 185
R1127 VTAIL.n61 VTAIL.n60 185
R1128 VTAIL.n59 VTAIL.n58 185
R1129 VTAIL.n50 VTAIL.n49 185
R1130 VTAIL.n53 VTAIL.n52 185
R1131 VTAIL.t19 VTAIL.n119 147.661
R1132 VTAIL.t10 VTAIL.n11 147.661
R1133 VTAIL.t15 VTAIL.n87 147.661
R1134 VTAIL.t18 VTAIL.n51 147.661
R1135 VTAIL.n120 VTAIL.n117 104.615
R1136 VTAIL.n127 VTAIL.n117 104.615
R1137 VTAIL.n128 VTAIL.n127 104.615
R1138 VTAIL.n128 VTAIL.n113 104.615
R1139 VTAIL.n135 VTAIL.n113 104.615
R1140 VTAIL.n136 VTAIL.n135 104.615
R1141 VTAIL.n12 VTAIL.n9 104.615
R1142 VTAIL.n19 VTAIL.n9 104.615
R1143 VTAIL.n20 VTAIL.n19 104.615
R1144 VTAIL.n20 VTAIL.n5 104.615
R1145 VTAIL.n27 VTAIL.n5 104.615
R1146 VTAIL.n28 VTAIL.n27 104.615
R1147 VTAIL.n104 VTAIL.n103 104.615
R1148 VTAIL.n103 VTAIL.n81 104.615
R1149 VTAIL.n96 VTAIL.n81 104.615
R1150 VTAIL.n96 VTAIL.n95 104.615
R1151 VTAIL.n95 VTAIL.n85 104.615
R1152 VTAIL.n88 VTAIL.n85 104.615
R1153 VTAIL.n68 VTAIL.n67 104.615
R1154 VTAIL.n67 VTAIL.n45 104.615
R1155 VTAIL.n60 VTAIL.n45 104.615
R1156 VTAIL.n60 VTAIL.n59 104.615
R1157 VTAIL.n59 VTAIL.n49 104.615
R1158 VTAIL.n52 VTAIL.n49 104.615
R1159 VTAIL.n120 VTAIL.t19 52.3082
R1160 VTAIL.n12 VTAIL.t10 52.3082
R1161 VTAIL.n88 VTAIL.t15 52.3082
R1162 VTAIL.n52 VTAIL.t18 52.3082
R1163 VTAIL.n77 VTAIL.n76 50.3181
R1164 VTAIL.n75 VTAIL.n74 50.3181
R1165 VTAIL.n41 VTAIL.n40 50.3181
R1166 VTAIL.n39 VTAIL.n38 50.3181
R1167 VTAIL.n143 VTAIL.n142 50.3179
R1168 VTAIL.n1 VTAIL.n0 50.3179
R1169 VTAIL.n35 VTAIL.n34 50.3179
R1170 VTAIL.n37 VTAIL.n36 50.3179
R1171 VTAIL.n141 VTAIL.n140 31.9914
R1172 VTAIL.n33 VTAIL.n32 31.9914
R1173 VTAIL.n109 VTAIL.n108 31.9914
R1174 VTAIL.n73 VTAIL.n72 31.9914
R1175 VTAIL.n39 VTAIL.n37 19.1169
R1176 VTAIL.n141 VTAIL.n109 18.3238
R1177 VTAIL.n121 VTAIL.n119 15.6674
R1178 VTAIL.n13 VTAIL.n11 15.6674
R1179 VTAIL.n89 VTAIL.n87 15.6674
R1180 VTAIL.n53 VTAIL.n51 15.6674
R1181 VTAIL.n122 VTAIL.n118 12.8005
R1182 VTAIL.n14 VTAIL.n10 12.8005
R1183 VTAIL.n90 VTAIL.n86 12.8005
R1184 VTAIL.n54 VTAIL.n50 12.8005
R1185 VTAIL.n126 VTAIL.n125 12.0247
R1186 VTAIL.n18 VTAIL.n17 12.0247
R1187 VTAIL.n94 VTAIL.n93 12.0247
R1188 VTAIL.n58 VTAIL.n57 12.0247
R1189 VTAIL.n129 VTAIL.n116 11.249
R1190 VTAIL.n21 VTAIL.n8 11.249
R1191 VTAIL.n97 VTAIL.n84 11.249
R1192 VTAIL.n61 VTAIL.n48 11.249
R1193 VTAIL.n130 VTAIL.n114 10.4732
R1194 VTAIL.n22 VTAIL.n6 10.4732
R1195 VTAIL.n98 VTAIL.n82 10.4732
R1196 VTAIL.n62 VTAIL.n46 10.4732
R1197 VTAIL.n134 VTAIL.n133 9.69747
R1198 VTAIL.n26 VTAIL.n25 9.69747
R1199 VTAIL.n102 VTAIL.n101 9.69747
R1200 VTAIL.n66 VTAIL.n65 9.69747
R1201 VTAIL.n140 VTAIL.n139 9.45567
R1202 VTAIL.n32 VTAIL.n31 9.45567
R1203 VTAIL.n108 VTAIL.n107 9.45567
R1204 VTAIL.n72 VTAIL.n71 9.45567
R1205 VTAIL.n139 VTAIL.n138 9.3005
R1206 VTAIL.n112 VTAIL.n111 9.3005
R1207 VTAIL.n133 VTAIL.n132 9.3005
R1208 VTAIL.n131 VTAIL.n130 9.3005
R1209 VTAIL.n116 VTAIL.n115 9.3005
R1210 VTAIL.n125 VTAIL.n124 9.3005
R1211 VTAIL.n123 VTAIL.n122 9.3005
R1212 VTAIL.n31 VTAIL.n30 9.3005
R1213 VTAIL.n4 VTAIL.n3 9.3005
R1214 VTAIL.n25 VTAIL.n24 9.3005
R1215 VTAIL.n23 VTAIL.n22 9.3005
R1216 VTAIL.n8 VTAIL.n7 9.3005
R1217 VTAIL.n17 VTAIL.n16 9.3005
R1218 VTAIL.n15 VTAIL.n14 9.3005
R1219 VTAIL.n107 VTAIL.n106 9.3005
R1220 VTAIL.n80 VTAIL.n79 9.3005
R1221 VTAIL.n101 VTAIL.n100 9.3005
R1222 VTAIL.n99 VTAIL.n98 9.3005
R1223 VTAIL.n84 VTAIL.n83 9.3005
R1224 VTAIL.n93 VTAIL.n92 9.3005
R1225 VTAIL.n91 VTAIL.n90 9.3005
R1226 VTAIL.n71 VTAIL.n70 9.3005
R1227 VTAIL.n44 VTAIL.n43 9.3005
R1228 VTAIL.n65 VTAIL.n64 9.3005
R1229 VTAIL.n63 VTAIL.n62 9.3005
R1230 VTAIL.n48 VTAIL.n47 9.3005
R1231 VTAIL.n57 VTAIL.n56 9.3005
R1232 VTAIL.n55 VTAIL.n54 9.3005
R1233 VTAIL.n137 VTAIL.n112 8.92171
R1234 VTAIL.n29 VTAIL.n4 8.92171
R1235 VTAIL.n105 VTAIL.n80 8.92171
R1236 VTAIL.n69 VTAIL.n44 8.92171
R1237 VTAIL.n138 VTAIL.n110 8.14595
R1238 VTAIL.n30 VTAIL.n2 8.14595
R1239 VTAIL.n106 VTAIL.n78 8.14595
R1240 VTAIL.n70 VTAIL.n42 8.14595
R1241 VTAIL.n140 VTAIL.n110 5.81868
R1242 VTAIL.n32 VTAIL.n2 5.81868
R1243 VTAIL.n108 VTAIL.n78 5.81868
R1244 VTAIL.n72 VTAIL.n42 5.81868
R1245 VTAIL.n138 VTAIL.n137 5.04292
R1246 VTAIL.n30 VTAIL.n29 5.04292
R1247 VTAIL.n106 VTAIL.n105 5.04292
R1248 VTAIL.n70 VTAIL.n69 5.04292
R1249 VTAIL.n123 VTAIL.n119 4.38594
R1250 VTAIL.n15 VTAIL.n11 4.38594
R1251 VTAIL.n91 VTAIL.n87 4.38594
R1252 VTAIL.n55 VTAIL.n51 4.38594
R1253 VTAIL.n134 VTAIL.n112 4.26717
R1254 VTAIL.n26 VTAIL.n4 4.26717
R1255 VTAIL.n102 VTAIL.n80 4.26717
R1256 VTAIL.n66 VTAIL.n44 4.26717
R1257 VTAIL.n133 VTAIL.n114 3.49141
R1258 VTAIL.n25 VTAIL.n6 3.49141
R1259 VTAIL.n101 VTAIL.n82 3.49141
R1260 VTAIL.n65 VTAIL.n46 3.49141
R1261 VTAIL.n142 VTAIL.t7 3.30601
R1262 VTAIL.n142 VTAIL.t1 3.30601
R1263 VTAIL.n0 VTAIL.t4 3.30601
R1264 VTAIL.n0 VTAIL.t5 3.30601
R1265 VTAIL.n34 VTAIL.t11 3.30601
R1266 VTAIL.n34 VTAIL.t9 3.30601
R1267 VTAIL.n36 VTAIL.t12 3.30601
R1268 VTAIL.n36 VTAIL.t14 3.30601
R1269 VTAIL.n76 VTAIL.t13 3.30601
R1270 VTAIL.n76 VTAIL.t17 3.30601
R1271 VTAIL.n74 VTAIL.t16 3.30601
R1272 VTAIL.n74 VTAIL.t8 3.30601
R1273 VTAIL.n40 VTAIL.t0 3.30601
R1274 VTAIL.n40 VTAIL.t3 3.30601
R1275 VTAIL.n38 VTAIL.t6 3.30601
R1276 VTAIL.n38 VTAIL.t2 3.30601
R1277 VTAIL.n130 VTAIL.n129 2.71565
R1278 VTAIL.n22 VTAIL.n21 2.71565
R1279 VTAIL.n98 VTAIL.n97 2.71565
R1280 VTAIL.n62 VTAIL.n61 2.71565
R1281 VTAIL.n126 VTAIL.n116 1.93989
R1282 VTAIL.n18 VTAIL.n8 1.93989
R1283 VTAIL.n94 VTAIL.n84 1.93989
R1284 VTAIL.n58 VTAIL.n48 1.93989
R1285 VTAIL.n125 VTAIL.n118 1.16414
R1286 VTAIL.n17 VTAIL.n10 1.16414
R1287 VTAIL.n93 VTAIL.n86 1.16414
R1288 VTAIL.n57 VTAIL.n50 1.16414
R1289 VTAIL.n75 VTAIL.n73 0.866879
R1290 VTAIL.n33 VTAIL.n1 0.866879
R1291 VTAIL.n41 VTAIL.n39 0.793603
R1292 VTAIL.n73 VTAIL.n41 0.793603
R1293 VTAIL.n77 VTAIL.n75 0.793603
R1294 VTAIL.n109 VTAIL.n77 0.793603
R1295 VTAIL.n37 VTAIL.n35 0.793603
R1296 VTAIL.n35 VTAIL.n33 0.793603
R1297 VTAIL.n143 VTAIL.n141 0.793603
R1298 VTAIL VTAIL.n1 0.653517
R1299 VTAIL.n122 VTAIL.n121 0.388379
R1300 VTAIL.n14 VTAIL.n13 0.388379
R1301 VTAIL.n90 VTAIL.n89 0.388379
R1302 VTAIL.n54 VTAIL.n53 0.388379
R1303 VTAIL.n124 VTAIL.n123 0.155672
R1304 VTAIL.n124 VTAIL.n115 0.155672
R1305 VTAIL.n131 VTAIL.n115 0.155672
R1306 VTAIL.n132 VTAIL.n131 0.155672
R1307 VTAIL.n132 VTAIL.n111 0.155672
R1308 VTAIL.n139 VTAIL.n111 0.155672
R1309 VTAIL.n16 VTAIL.n15 0.155672
R1310 VTAIL.n16 VTAIL.n7 0.155672
R1311 VTAIL.n23 VTAIL.n7 0.155672
R1312 VTAIL.n24 VTAIL.n23 0.155672
R1313 VTAIL.n24 VTAIL.n3 0.155672
R1314 VTAIL.n31 VTAIL.n3 0.155672
R1315 VTAIL.n107 VTAIL.n79 0.155672
R1316 VTAIL.n100 VTAIL.n79 0.155672
R1317 VTAIL.n100 VTAIL.n99 0.155672
R1318 VTAIL.n99 VTAIL.n83 0.155672
R1319 VTAIL.n92 VTAIL.n83 0.155672
R1320 VTAIL.n92 VTAIL.n91 0.155672
R1321 VTAIL.n71 VTAIL.n43 0.155672
R1322 VTAIL.n64 VTAIL.n43 0.155672
R1323 VTAIL.n64 VTAIL.n63 0.155672
R1324 VTAIL.n63 VTAIL.n47 0.155672
R1325 VTAIL.n56 VTAIL.n47 0.155672
R1326 VTAIL.n56 VTAIL.n55 0.155672
R1327 VTAIL VTAIL.n143 0.140586
R1328 VN.n3 VN.t5 337.387
R1329 VN.n13 VN.t6 337.387
R1330 VN.n2 VN.t3 311.666
R1331 VN.n1 VN.t4 311.666
R1332 VN.n6 VN.t1 311.666
R1333 VN.n8 VN.t9 311.666
R1334 VN.n12 VN.t2 311.666
R1335 VN.n11 VN.t8 311.666
R1336 VN.n16 VN.t0 311.666
R1337 VN.n18 VN.t7 311.666
R1338 VN.n9 VN.n8 161.3
R1339 VN.n19 VN.n18 161.3
R1340 VN.n17 VN.n10 161.3
R1341 VN.n16 VN.n15 161.3
R1342 VN.n7 VN.n0 161.3
R1343 VN.n6 VN.n5 161.3
R1344 VN.n14 VN.n11 80.6037
R1345 VN.n4 VN.n1 80.6037
R1346 VN.n2 VN.n1 48.2005
R1347 VN.n6 VN.n1 48.2005
R1348 VN.n12 VN.n11 48.2005
R1349 VN.n16 VN.n11 48.2005
R1350 VN.n14 VN.n13 45.1242
R1351 VN.n4 VN.n3 45.1242
R1352 VN.n8 VN.n7 43.0884
R1353 VN.n18 VN.n17 43.0884
R1354 VN VN.n19 38.01
R1355 VN.n3 VN.n2 15.1442
R1356 VN.n13 VN.n12 15.1442
R1357 VN.n7 VN.n6 5.11262
R1358 VN.n17 VN.n16 5.11262
R1359 VN.n15 VN.n14 0.285035
R1360 VN.n5 VN.n4 0.285035
R1361 VN.n19 VN.n10 0.189894
R1362 VN.n15 VN.n10 0.189894
R1363 VN.n5 VN.n0 0.189894
R1364 VN.n9 VN.n0 0.189894
R1365 VN VN.n9 0.0516364
R1366 VDD2.n61 VDD2.n35 289.615
R1367 VDD2.n26 VDD2.n0 289.615
R1368 VDD2.n62 VDD2.n61 185
R1369 VDD2.n60 VDD2.n59 185
R1370 VDD2.n39 VDD2.n38 185
R1371 VDD2.n54 VDD2.n53 185
R1372 VDD2.n52 VDD2.n51 185
R1373 VDD2.n43 VDD2.n42 185
R1374 VDD2.n46 VDD2.n45 185
R1375 VDD2.n11 VDD2.n10 185
R1376 VDD2.n8 VDD2.n7 185
R1377 VDD2.n17 VDD2.n16 185
R1378 VDD2.n19 VDD2.n18 185
R1379 VDD2.n4 VDD2.n3 185
R1380 VDD2.n25 VDD2.n24 185
R1381 VDD2.n27 VDD2.n26 185
R1382 VDD2.t2 VDD2.n44 147.661
R1383 VDD2.t4 VDD2.n9 147.661
R1384 VDD2.n61 VDD2.n60 104.615
R1385 VDD2.n60 VDD2.n38 104.615
R1386 VDD2.n53 VDD2.n38 104.615
R1387 VDD2.n53 VDD2.n52 104.615
R1388 VDD2.n52 VDD2.n42 104.615
R1389 VDD2.n45 VDD2.n42 104.615
R1390 VDD2.n10 VDD2.n7 104.615
R1391 VDD2.n17 VDD2.n7 104.615
R1392 VDD2.n18 VDD2.n17 104.615
R1393 VDD2.n18 VDD2.n3 104.615
R1394 VDD2.n25 VDD2.n3 104.615
R1395 VDD2.n26 VDD2.n25 104.615
R1396 VDD2.n34 VDD2.n33 67.5362
R1397 VDD2 VDD2.n69 67.5334
R1398 VDD2.n68 VDD2.n67 66.9969
R1399 VDD2.n32 VDD2.n31 66.9967
R1400 VDD2.n45 VDD2.t2 52.3082
R1401 VDD2.n10 VDD2.t4 52.3082
R1402 VDD2.n32 VDD2.n30 49.4633
R1403 VDD2.n66 VDD2.n65 48.6702
R1404 VDD2.n66 VDD2.n34 32.6463
R1405 VDD2.n46 VDD2.n44 15.6674
R1406 VDD2.n11 VDD2.n9 15.6674
R1407 VDD2.n47 VDD2.n43 12.8005
R1408 VDD2.n12 VDD2.n8 12.8005
R1409 VDD2.n51 VDD2.n50 12.0247
R1410 VDD2.n16 VDD2.n15 12.0247
R1411 VDD2.n54 VDD2.n41 11.249
R1412 VDD2.n19 VDD2.n6 11.249
R1413 VDD2.n55 VDD2.n39 10.4732
R1414 VDD2.n20 VDD2.n4 10.4732
R1415 VDD2.n59 VDD2.n58 9.69747
R1416 VDD2.n24 VDD2.n23 9.69747
R1417 VDD2.n65 VDD2.n64 9.45567
R1418 VDD2.n30 VDD2.n29 9.45567
R1419 VDD2.n64 VDD2.n63 9.3005
R1420 VDD2.n37 VDD2.n36 9.3005
R1421 VDD2.n58 VDD2.n57 9.3005
R1422 VDD2.n56 VDD2.n55 9.3005
R1423 VDD2.n41 VDD2.n40 9.3005
R1424 VDD2.n50 VDD2.n49 9.3005
R1425 VDD2.n48 VDD2.n47 9.3005
R1426 VDD2.n29 VDD2.n28 9.3005
R1427 VDD2.n2 VDD2.n1 9.3005
R1428 VDD2.n23 VDD2.n22 9.3005
R1429 VDD2.n21 VDD2.n20 9.3005
R1430 VDD2.n6 VDD2.n5 9.3005
R1431 VDD2.n15 VDD2.n14 9.3005
R1432 VDD2.n13 VDD2.n12 9.3005
R1433 VDD2.n62 VDD2.n37 8.92171
R1434 VDD2.n27 VDD2.n2 8.92171
R1435 VDD2.n63 VDD2.n35 8.14595
R1436 VDD2.n28 VDD2.n0 8.14595
R1437 VDD2.n65 VDD2.n35 5.81868
R1438 VDD2.n30 VDD2.n0 5.81868
R1439 VDD2.n63 VDD2.n62 5.04292
R1440 VDD2.n28 VDD2.n27 5.04292
R1441 VDD2.n48 VDD2.n44 4.38594
R1442 VDD2.n13 VDD2.n9 4.38594
R1443 VDD2.n59 VDD2.n37 4.26717
R1444 VDD2.n24 VDD2.n2 4.26717
R1445 VDD2.n58 VDD2.n39 3.49141
R1446 VDD2.n23 VDD2.n4 3.49141
R1447 VDD2.n69 VDD2.t7 3.30601
R1448 VDD2.n69 VDD2.t3 3.30601
R1449 VDD2.n67 VDD2.t9 3.30601
R1450 VDD2.n67 VDD2.t1 3.30601
R1451 VDD2.n33 VDD2.t8 3.30601
R1452 VDD2.n33 VDD2.t0 3.30601
R1453 VDD2.n31 VDD2.t6 3.30601
R1454 VDD2.n31 VDD2.t5 3.30601
R1455 VDD2.n55 VDD2.n54 2.71565
R1456 VDD2.n20 VDD2.n19 2.71565
R1457 VDD2.n51 VDD2.n41 1.93989
R1458 VDD2.n16 VDD2.n6 1.93989
R1459 VDD2.n50 VDD2.n43 1.16414
R1460 VDD2.n15 VDD2.n8 1.16414
R1461 VDD2.n68 VDD2.n66 0.793603
R1462 VDD2.n47 VDD2.n46 0.388379
R1463 VDD2.n12 VDD2.n11 0.388379
R1464 VDD2 VDD2.n68 0.256966
R1465 VDD2.n64 VDD2.n36 0.155672
R1466 VDD2.n57 VDD2.n36 0.155672
R1467 VDD2.n57 VDD2.n56 0.155672
R1468 VDD2.n56 VDD2.n40 0.155672
R1469 VDD2.n49 VDD2.n40 0.155672
R1470 VDD2.n49 VDD2.n48 0.155672
R1471 VDD2.n14 VDD2.n13 0.155672
R1472 VDD2.n14 VDD2.n5 0.155672
R1473 VDD2.n21 VDD2.n5 0.155672
R1474 VDD2.n22 VDD2.n21 0.155672
R1475 VDD2.n22 VDD2.n1 0.155672
R1476 VDD2.n29 VDD2.n1 0.155672
R1477 VDD2.n34 VDD2.n32 0.14343
C0 VTAIL VP 3.34062f
C1 VTAIL VDD1 8.85452f
C2 VN VDD2 3.24924f
C3 VDD2 VP 0.3267f
C4 VN VP 4.32369f
C5 VDD2 VDD1 0.90257f
C6 VN VDD1 0.148821f
C7 VDD1 VP 3.42446f
C8 VDD2 VTAIL 8.891081f
C9 VN VTAIL 3.32624f
C10 VDD2 B 3.774201f
C11 VDD1 B 3.691777f
C12 VTAIL B 4.103954f
C13 VN B 8.18143f
C14 VP B 6.482685f
C15 VDD2.n0 B 0.035176f
C16 VDD2.n1 B 0.025146f
C17 VDD2.n2 B 0.013513f
C18 VDD2.n3 B 0.031939f
C19 VDD2.n4 B 0.014307f
C20 VDD2.n5 B 0.025146f
C21 VDD2.n6 B 0.013513f
C22 VDD2.n7 B 0.031939f
C23 VDD2.n8 B 0.014307f
C24 VDD2.n9 B 0.107539f
C25 VDD2.t4 B 0.052052f
C26 VDD2.n10 B 0.023954f
C27 VDD2.n11 B 0.018866f
C28 VDD2.n12 B 0.013513f
C29 VDD2.n13 B 0.59719f
C30 VDD2.n14 B 0.025146f
C31 VDD2.n15 B 0.013513f
C32 VDD2.n16 B 0.014307f
C33 VDD2.n17 B 0.031939f
C34 VDD2.n18 B 0.031939f
C35 VDD2.n19 B 0.014307f
C36 VDD2.n20 B 0.013513f
C37 VDD2.n21 B 0.025146f
C38 VDD2.n22 B 0.025146f
C39 VDD2.n23 B 0.013513f
C40 VDD2.n24 B 0.014307f
C41 VDD2.n25 B 0.031939f
C42 VDD2.n26 B 0.068842f
C43 VDD2.n27 B 0.014307f
C44 VDD2.n28 B 0.013513f
C45 VDD2.n29 B 0.057781f
C46 VDD2.n30 B 0.057648f
C47 VDD2.t6 B 0.11903f
C48 VDD2.t5 B 0.11903f
C49 VDD2.n31 B 0.992438f
C50 VDD2.n32 B 0.39474f
C51 VDD2.t8 B 0.11903f
C52 VDD2.t0 B 0.11903f
C53 VDD2.n33 B 0.995021f
C54 VDD2.n34 B 1.49326f
C55 VDD2.n35 B 0.035176f
C56 VDD2.n36 B 0.025146f
C57 VDD2.n37 B 0.013513f
C58 VDD2.n38 B 0.031939f
C59 VDD2.n39 B 0.014307f
C60 VDD2.n40 B 0.025146f
C61 VDD2.n41 B 0.013513f
C62 VDD2.n42 B 0.031939f
C63 VDD2.n43 B 0.014307f
C64 VDD2.n44 B 0.107539f
C65 VDD2.t2 B 0.052052f
C66 VDD2.n45 B 0.023954f
C67 VDD2.n46 B 0.018866f
C68 VDD2.n47 B 0.013513f
C69 VDD2.n48 B 0.59719f
C70 VDD2.n49 B 0.025146f
C71 VDD2.n50 B 0.013513f
C72 VDD2.n51 B 0.014307f
C73 VDD2.n52 B 0.031939f
C74 VDD2.n53 B 0.031939f
C75 VDD2.n54 B 0.014307f
C76 VDD2.n55 B 0.013513f
C77 VDD2.n56 B 0.025146f
C78 VDD2.n57 B 0.025146f
C79 VDD2.n58 B 0.013513f
C80 VDD2.n59 B 0.014307f
C81 VDD2.n60 B 0.031939f
C82 VDD2.n61 B 0.068842f
C83 VDD2.n62 B 0.014307f
C84 VDD2.n63 B 0.013513f
C85 VDD2.n64 B 0.057781f
C86 VDD2.n65 B 0.055844f
C87 VDD2.n66 B 1.64397f
C88 VDD2.t9 B 0.11903f
C89 VDD2.t1 B 0.11903f
C90 VDD2.n67 B 0.992443f
C91 VDD2.n68 B 0.289173f
C92 VDD2.t7 B 0.11903f
C93 VDD2.t3 B 0.11903f
C94 VDD2.n69 B 0.994997f
C95 VN.n0 B 0.045606f
C96 VN.t4 B 0.467778f
C97 VN.n1 B 0.229074f
C98 VN.t5 B 0.484431f
C99 VN.t3 B 0.467778f
C100 VN.n2 B 0.227864f
C101 VN.n3 B 0.204612f
C102 VN.n4 B 0.219043f
C103 VN.n5 B 0.060856f
C104 VN.t1 B 0.467778f
C105 VN.n6 B 0.219709f
C106 VN.n7 B 0.010349f
C107 VN.t9 B 0.467778f
C108 VN.n8 B 0.217741f
C109 VN.n9 B 0.035343f
C110 VN.n10 B 0.045606f
C111 VN.t8 B 0.467778f
C112 VN.n11 B 0.229074f
C113 VN.t0 B 0.467778f
C114 VN.t6 B 0.484431f
C115 VN.t2 B 0.467778f
C116 VN.n12 B 0.227864f
C117 VN.n13 B 0.204612f
C118 VN.n14 B 0.219043f
C119 VN.n15 B 0.060856f
C120 VN.n16 B 0.219709f
C121 VN.n17 B 0.010349f
C122 VN.t7 B 0.467778f
C123 VN.n18 B 0.217741f
C124 VN.n19 B 1.58592f
C125 VTAIL.t4 B 0.132701f
C126 VTAIL.t5 B 0.132701f
C127 VTAIL.n0 B 1.03276f
C128 VTAIL.n1 B 0.400394f
C129 VTAIL.n2 B 0.039216f
C130 VTAIL.n3 B 0.028035f
C131 VTAIL.n4 B 0.015064f
C132 VTAIL.n5 B 0.035607f
C133 VTAIL.n6 B 0.015951f
C134 VTAIL.n7 B 0.028035f
C135 VTAIL.n8 B 0.015064f
C136 VTAIL.n9 B 0.035607f
C137 VTAIL.n10 B 0.015951f
C138 VTAIL.n11 B 0.11989f
C139 VTAIL.t10 B 0.05803f
C140 VTAIL.n12 B 0.026705f
C141 VTAIL.n13 B 0.021033f
C142 VTAIL.n14 B 0.015064f
C143 VTAIL.n15 B 0.665781f
C144 VTAIL.n16 B 0.028035f
C145 VTAIL.n17 B 0.015064f
C146 VTAIL.n18 B 0.015951f
C147 VTAIL.n19 B 0.035607f
C148 VTAIL.n20 B 0.035607f
C149 VTAIL.n21 B 0.015951f
C150 VTAIL.n22 B 0.015064f
C151 VTAIL.n23 B 0.028035f
C152 VTAIL.n24 B 0.028035f
C153 VTAIL.n25 B 0.015064f
C154 VTAIL.n26 B 0.015951f
C155 VTAIL.n27 B 0.035607f
C156 VTAIL.n28 B 0.076749f
C157 VTAIL.n29 B 0.015951f
C158 VTAIL.n30 B 0.015064f
C159 VTAIL.n31 B 0.064418f
C160 VTAIL.n32 B 0.042898f
C161 VTAIL.n33 B 0.173634f
C162 VTAIL.t11 B 0.132701f
C163 VTAIL.t9 B 0.132701f
C164 VTAIL.n34 B 1.03276f
C165 VTAIL.n35 B 0.40643f
C166 VTAIL.t12 B 0.132701f
C167 VTAIL.t14 B 0.132701f
C168 VTAIL.n36 B 1.03276f
C169 VTAIL.n37 B 1.32535f
C170 VTAIL.t6 B 0.132701f
C171 VTAIL.t2 B 0.132701f
C172 VTAIL.n38 B 1.03277f
C173 VTAIL.n39 B 1.32535f
C174 VTAIL.t0 B 0.132701f
C175 VTAIL.t3 B 0.132701f
C176 VTAIL.n40 B 1.03277f
C177 VTAIL.n41 B 0.406422f
C178 VTAIL.n42 B 0.039216f
C179 VTAIL.n43 B 0.028035f
C180 VTAIL.n44 B 0.015064f
C181 VTAIL.n45 B 0.035607f
C182 VTAIL.n46 B 0.015951f
C183 VTAIL.n47 B 0.028035f
C184 VTAIL.n48 B 0.015064f
C185 VTAIL.n49 B 0.035607f
C186 VTAIL.n50 B 0.015951f
C187 VTAIL.n51 B 0.11989f
C188 VTAIL.t18 B 0.05803f
C189 VTAIL.n52 B 0.026705f
C190 VTAIL.n53 B 0.021033f
C191 VTAIL.n54 B 0.015064f
C192 VTAIL.n55 B 0.665781f
C193 VTAIL.n56 B 0.028035f
C194 VTAIL.n57 B 0.015064f
C195 VTAIL.n58 B 0.015951f
C196 VTAIL.n59 B 0.035607f
C197 VTAIL.n60 B 0.035607f
C198 VTAIL.n61 B 0.015951f
C199 VTAIL.n62 B 0.015064f
C200 VTAIL.n63 B 0.028035f
C201 VTAIL.n64 B 0.028035f
C202 VTAIL.n65 B 0.015064f
C203 VTAIL.n66 B 0.015951f
C204 VTAIL.n67 B 0.035607f
C205 VTAIL.n68 B 0.076749f
C206 VTAIL.n69 B 0.015951f
C207 VTAIL.n70 B 0.015064f
C208 VTAIL.n71 B 0.064418f
C209 VTAIL.n72 B 0.042898f
C210 VTAIL.n73 B 0.173634f
C211 VTAIL.t16 B 0.132701f
C212 VTAIL.t8 B 0.132701f
C213 VTAIL.n74 B 1.03277f
C214 VTAIL.n75 B 0.413042f
C215 VTAIL.t13 B 0.132701f
C216 VTAIL.t17 B 0.132701f
C217 VTAIL.n76 B 1.03277f
C218 VTAIL.n77 B 0.406422f
C219 VTAIL.n78 B 0.039216f
C220 VTAIL.n79 B 0.028035f
C221 VTAIL.n80 B 0.015064f
C222 VTAIL.n81 B 0.035607f
C223 VTAIL.n82 B 0.015951f
C224 VTAIL.n83 B 0.028035f
C225 VTAIL.n84 B 0.015064f
C226 VTAIL.n85 B 0.035607f
C227 VTAIL.n86 B 0.015951f
C228 VTAIL.n87 B 0.11989f
C229 VTAIL.t15 B 0.05803f
C230 VTAIL.n88 B 0.026705f
C231 VTAIL.n89 B 0.021033f
C232 VTAIL.n90 B 0.015064f
C233 VTAIL.n91 B 0.665781f
C234 VTAIL.n92 B 0.028035f
C235 VTAIL.n93 B 0.015064f
C236 VTAIL.n94 B 0.015951f
C237 VTAIL.n95 B 0.035607f
C238 VTAIL.n96 B 0.035607f
C239 VTAIL.n97 B 0.015951f
C240 VTAIL.n98 B 0.015064f
C241 VTAIL.n99 B 0.028035f
C242 VTAIL.n100 B 0.028035f
C243 VTAIL.n101 B 0.015064f
C244 VTAIL.n102 B 0.015951f
C245 VTAIL.n103 B 0.035607f
C246 VTAIL.n104 B 0.076749f
C247 VTAIL.n105 B 0.015951f
C248 VTAIL.n106 B 0.015064f
C249 VTAIL.n107 B 0.064418f
C250 VTAIL.n108 B 0.042898f
C251 VTAIL.n109 B 1.0143f
C252 VTAIL.n110 B 0.039216f
C253 VTAIL.n111 B 0.028035f
C254 VTAIL.n112 B 0.015064f
C255 VTAIL.n113 B 0.035607f
C256 VTAIL.n114 B 0.015951f
C257 VTAIL.n115 B 0.028035f
C258 VTAIL.n116 B 0.015064f
C259 VTAIL.n117 B 0.035607f
C260 VTAIL.n118 B 0.015951f
C261 VTAIL.n119 B 0.11989f
C262 VTAIL.t19 B 0.05803f
C263 VTAIL.n120 B 0.026705f
C264 VTAIL.n121 B 0.021033f
C265 VTAIL.n122 B 0.015064f
C266 VTAIL.n123 B 0.665781f
C267 VTAIL.n124 B 0.028035f
C268 VTAIL.n125 B 0.015064f
C269 VTAIL.n126 B 0.015951f
C270 VTAIL.n127 B 0.035607f
C271 VTAIL.n128 B 0.035607f
C272 VTAIL.n129 B 0.015951f
C273 VTAIL.n130 B 0.015064f
C274 VTAIL.n131 B 0.028035f
C275 VTAIL.n132 B 0.028035f
C276 VTAIL.n133 B 0.015064f
C277 VTAIL.n134 B 0.015951f
C278 VTAIL.n135 B 0.035607f
C279 VTAIL.n136 B 0.076749f
C280 VTAIL.n137 B 0.015951f
C281 VTAIL.n138 B 0.015064f
C282 VTAIL.n139 B 0.064418f
C283 VTAIL.n140 B 0.042898f
C284 VTAIL.n141 B 1.0143f
C285 VTAIL.t7 B 0.132701f
C286 VTAIL.t1 B 0.132701f
C287 VTAIL.n142 B 1.03276f
C288 VTAIL.n143 B 0.34744f
C289 VDD1.n0 B 0.035485f
C290 VDD1.n1 B 0.025367f
C291 VDD1.n2 B 0.013631f
C292 VDD1.n3 B 0.032219f
C293 VDD1.n4 B 0.014433f
C294 VDD1.n5 B 0.025367f
C295 VDD1.n6 B 0.013631f
C296 VDD1.n7 B 0.032219f
C297 VDD1.n8 B 0.014433f
C298 VDD1.n9 B 0.108484f
C299 VDD1.t2 B 0.052509f
C300 VDD1.n10 B 0.024164f
C301 VDD1.n11 B 0.019032f
C302 VDD1.n12 B 0.013631f
C303 VDD1.n13 B 0.602437f
C304 VDD1.n14 B 0.025367f
C305 VDD1.n15 B 0.013631f
C306 VDD1.n16 B 0.014433f
C307 VDD1.n17 B 0.032219f
C308 VDD1.n18 B 0.032219f
C309 VDD1.n19 B 0.014433f
C310 VDD1.n20 B 0.013631f
C311 VDD1.n21 B 0.025367f
C312 VDD1.n22 B 0.025367f
C313 VDD1.n23 B 0.013631f
C314 VDD1.n24 B 0.014433f
C315 VDD1.n25 B 0.032219f
C316 VDD1.n26 B 0.069447f
C317 VDD1.n27 B 0.014433f
C318 VDD1.n28 B 0.013631f
C319 VDD1.n29 B 0.058289f
C320 VDD1.n30 B 0.058154f
C321 VDD1.t0 B 0.120075f
C322 VDD1.t5 B 0.120075f
C323 VDD1.n31 B 1.00116f
C324 VDD1.n32 B 0.403369f
C325 VDD1.n33 B 0.035485f
C326 VDD1.n34 B 0.025367f
C327 VDD1.n35 B 0.013631f
C328 VDD1.n36 B 0.032219f
C329 VDD1.n37 B 0.014433f
C330 VDD1.n38 B 0.025367f
C331 VDD1.n39 B 0.013631f
C332 VDD1.n40 B 0.032219f
C333 VDD1.n41 B 0.014433f
C334 VDD1.n42 B 0.108484f
C335 VDD1.t6 B 0.052509f
C336 VDD1.n43 B 0.024164f
C337 VDD1.n44 B 0.019032f
C338 VDD1.n45 B 0.013631f
C339 VDD1.n46 B 0.602437f
C340 VDD1.n47 B 0.025367f
C341 VDD1.n48 B 0.013631f
C342 VDD1.n49 B 0.014433f
C343 VDD1.n50 B 0.032219f
C344 VDD1.n51 B 0.032219f
C345 VDD1.n52 B 0.014433f
C346 VDD1.n53 B 0.013631f
C347 VDD1.n54 B 0.025367f
C348 VDD1.n55 B 0.025367f
C349 VDD1.n56 B 0.013631f
C350 VDD1.n57 B 0.014433f
C351 VDD1.n58 B 0.032219f
C352 VDD1.n59 B 0.069447f
C353 VDD1.n60 B 0.014433f
C354 VDD1.n61 B 0.013631f
C355 VDD1.n62 B 0.058289f
C356 VDD1.n63 B 0.058154f
C357 VDD1.t4 B 0.120075f
C358 VDD1.t8 B 0.120075f
C359 VDD1.n64 B 1.00116f
C360 VDD1.n65 B 0.398208f
C361 VDD1.t9 B 0.120075f
C362 VDD1.t7 B 0.120075f
C363 VDD1.n66 B 1.00376f
C364 VDD1.n67 B 1.57967f
C365 VDD1.t1 B 0.120075f
C366 VDD1.t3 B 0.120075f
C367 VDD1.n68 B 1.00116f
C368 VDD1.n69 B 1.89018f
C369 VP.n0 B 0.046728f
C370 VP.t6 B 0.479286f
C371 VP.n1 B 0.23471f
C372 VP.n2 B 0.046728f
C373 VP.n3 B 0.046728f
C374 VP.t2 B 0.479286f
C375 VP.t0 B 0.479286f
C376 VP.n4 B 0.062353f
C377 VP.t4 B 0.479286f
C378 VP.n5 B 0.224432f
C379 VP.t9 B 0.479286f
C380 VP.t1 B 0.496349f
C381 VP.n6 B 0.209645f
C382 VP.n7 B 0.233469f
C383 VP.n8 B 0.23471f
C384 VP.n9 B 0.225114f
C385 VP.n10 B 0.010603f
C386 VP.n11 B 0.223098f
C387 VP.n12 B 1.59404f
C388 VP.n13 B 1.63868f
C389 VP.t5 B 0.479286f
C390 VP.n14 B 0.223098f
C391 VP.n15 B 0.010603f
C392 VP.t3 B 0.479286f
C393 VP.n16 B 0.225114f
C394 VP.n17 B 0.062353f
C395 VP.n18 B 0.062207f
C396 VP.n19 B 0.062353f
C397 VP.t8 B 0.479286f
C398 VP.n20 B 0.225114f
C399 VP.n21 B 0.010603f
C400 VP.t7 B 0.479286f
C401 VP.n22 B 0.223098f
C402 VP.n23 B 0.036212f
.ends

