* NGSPICE file created from diff_pair_sample_0556.ext - technology: sky130A

.subckt diff_pair_sample_0556 VTAIL VN VP B VDD2 VDD1
X0 B.t19 B.t17 B.t18 B.t14 sky130_fd_pr__nfet_01v8 ad=7.5153 pd=39.32 as=0 ps=0 w=19.27 l=0.41
X1 VDD2.t5 VN.t0 VTAIL.t8 B.t1 sky130_fd_pr__nfet_01v8 ad=7.5153 pd=39.32 as=3.17955 ps=19.6 w=19.27 l=0.41
X2 VDD1.t5 VP.t0 VTAIL.t0 B.t4 sky130_fd_pr__nfet_01v8 ad=7.5153 pd=39.32 as=3.17955 ps=19.6 w=19.27 l=0.41
X3 B.t16 B.t13 B.t15 B.t14 sky130_fd_pr__nfet_01v8 ad=7.5153 pd=39.32 as=0 ps=0 w=19.27 l=0.41
X4 VTAIL.t5 VP.t1 VDD1.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=3.17955 pd=19.6 as=3.17955 ps=19.6 w=19.27 l=0.41
X5 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=7.5153 pd=39.32 as=0 ps=0 w=19.27 l=0.41
X6 VDD1.t3 VP.t2 VTAIL.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=3.17955 pd=19.6 as=7.5153 ps=39.32 w=19.27 l=0.41
X7 VDD1.t2 VP.t3 VTAIL.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=3.17955 pd=19.6 as=7.5153 ps=39.32 w=19.27 l=0.41
X8 VDD2.t4 VN.t1 VTAIL.t9 B.t4 sky130_fd_pr__nfet_01v8 ad=7.5153 pd=39.32 as=3.17955 ps=19.6 w=19.27 l=0.41
X9 VDD2.t3 VN.t2 VTAIL.t10 B.t3 sky130_fd_pr__nfet_01v8 ad=3.17955 pd=19.6 as=7.5153 ps=39.32 w=19.27 l=0.41
X10 VTAIL.t6 VN.t3 VDD2.t2 B.t5 sky130_fd_pr__nfet_01v8 ad=3.17955 pd=19.6 as=3.17955 ps=19.6 w=19.27 l=0.41
X11 VDD1.t1 VP.t4 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=7.5153 pd=39.32 as=3.17955 ps=19.6 w=19.27 l=0.41
X12 VDD2.t1 VN.t4 VTAIL.t11 B.t2 sky130_fd_pr__nfet_01v8 ad=3.17955 pd=19.6 as=7.5153 ps=39.32 w=19.27 l=0.41
X13 VTAIL.t2 VP.t5 VDD1.t0 B.t5 sky130_fd_pr__nfet_01v8 ad=3.17955 pd=19.6 as=3.17955 ps=19.6 w=19.27 l=0.41
X14 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=7.5153 pd=39.32 as=0 ps=0 w=19.27 l=0.41
X15 VTAIL.t7 VN.t5 VDD2.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=3.17955 pd=19.6 as=3.17955 ps=19.6 w=19.27 l=0.41
R0 B.n482 B.t10 1341.75
R1 B.n479 B.t6 1341.75
R2 B.n105 B.t13 1341.75
R3 B.n103 B.t17 1341.75
R4 B.n829 B.n828 585
R5 B.n377 B.n102 585
R6 B.n376 B.n375 585
R7 B.n374 B.n373 585
R8 B.n372 B.n371 585
R9 B.n370 B.n369 585
R10 B.n368 B.n367 585
R11 B.n366 B.n365 585
R12 B.n364 B.n363 585
R13 B.n362 B.n361 585
R14 B.n360 B.n359 585
R15 B.n358 B.n357 585
R16 B.n356 B.n355 585
R17 B.n354 B.n353 585
R18 B.n352 B.n351 585
R19 B.n350 B.n349 585
R20 B.n348 B.n347 585
R21 B.n346 B.n345 585
R22 B.n344 B.n343 585
R23 B.n342 B.n341 585
R24 B.n340 B.n339 585
R25 B.n338 B.n337 585
R26 B.n336 B.n335 585
R27 B.n334 B.n333 585
R28 B.n332 B.n331 585
R29 B.n330 B.n329 585
R30 B.n328 B.n327 585
R31 B.n326 B.n325 585
R32 B.n324 B.n323 585
R33 B.n322 B.n321 585
R34 B.n320 B.n319 585
R35 B.n318 B.n317 585
R36 B.n316 B.n315 585
R37 B.n314 B.n313 585
R38 B.n312 B.n311 585
R39 B.n310 B.n309 585
R40 B.n308 B.n307 585
R41 B.n306 B.n305 585
R42 B.n304 B.n303 585
R43 B.n302 B.n301 585
R44 B.n300 B.n299 585
R45 B.n298 B.n297 585
R46 B.n296 B.n295 585
R47 B.n294 B.n293 585
R48 B.n292 B.n291 585
R49 B.n290 B.n289 585
R50 B.n288 B.n287 585
R51 B.n286 B.n285 585
R52 B.n284 B.n283 585
R53 B.n282 B.n281 585
R54 B.n280 B.n279 585
R55 B.n278 B.n277 585
R56 B.n276 B.n275 585
R57 B.n274 B.n273 585
R58 B.n272 B.n271 585
R59 B.n270 B.n269 585
R60 B.n268 B.n267 585
R61 B.n266 B.n265 585
R62 B.n264 B.n263 585
R63 B.n262 B.n261 585
R64 B.n260 B.n259 585
R65 B.n258 B.n257 585
R66 B.n256 B.n255 585
R67 B.n253 B.n252 585
R68 B.n251 B.n250 585
R69 B.n249 B.n248 585
R70 B.n247 B.n246 585
R71 B.n245 B.n244 585
R72 B.n243 B.n242 585
R73 B.n241 B.n240 585
R74 B.n239 B.n238 585
R75 B.n237 B.n236 585
R76 B.n235 B.n234 585
R77 B.n232 B.n231 585
R78 B.n230 B.n229 585
R79 B.n228 B.n227 585
R80 B.n226 B.n225 585
R81 B.n224 B.n223 585
R82 B.n222 B.n221 585
R83 B.n220 B.n219 585
R84 B.n218 B.n217 585
R85 B.n216 B.n215 585
R86 B.n214 B.n213 585
R87 B.n212 B.n211 585
R88 B.n210 B.n209 585
R89 B.n208 B.n207 585
R90 B.n206 B.n205 585
R91 B.n204 B.n203 585
R92 B.n202 B.n201 585
R93 B.n200 B.n199 585
R94 B.n198 B.n197 585
R95 B.n196 B.n195 585
R96 B.n194 B.n193 585
R97 B.n192 B.n191 585
R98 B.n190 B.n189 585
R99 B.n188 B.n187 585
R100 B.n186 B.n185 585
R101 B.n184 B.n183 585
R102 B.n182 B.n181 585
R103 B.n180 B.n179 585
R104 B.n178 B.n177 585
R105 B.n176 B.n175 585
R106 B.n174 B.n173 585
R107 B.n172 B.n171 585
R108 B.n170 B.n169 585
R109 B.n168 B.n167 585
R110 B.n166 B.n165 585
R111 B.n164 B.n163 585
R112 B.n162 B.n161 585
R113 B.n160 B.n159 585
R114 B.n158 B.n157 585
R115 B.n156 B.n155 585
R116 B.n154 B.n153 585
R117 B.n152 B.n151 585
R118 B.n150 B.n149 585
R119 B.n148 B.n147 585
R120 B.n146 B.n145 585
R121 B.n144 B.n143 585
R122 B.n142 B.n141 585
R123 B.n140 B.n139 585
R124 B.n138 B.n137 585
R125 B.n136 B.n135 585
R126 B.n134 B.n133 585
R127 B.n132 B.n131 585
R128 B.n130 B.n129 585
R129 B.n128 B.n127 585
R130 B.n126 B.n125 585
R131 B.n124 B.n123 585
R132 B.n122 B.n121 585
R133 B.n120 B.n119 585
R134 B.n118 B.n117 585
R135 B.n116 B.n115 585
R136 B.n114 B.n113 585
R137 B.n112 B.n111 585
R138 B.n110 B.n109 585
R139 B.n108 B.n107 585
R140 B.n827 B.n34 585
R141 B.n832 B.n34 585
R142 B.n826 B.n33 585
R143 B.n833 B.n33 585
R144 B.n825 B.n824 585
R145 B.n824 B.n29 585
R146 B.n823 B.n28 585
R147 B.n839 B.n28 585
R148 B.n822 B.n27 585
R149 B.n840 B.n27 585
R150 B.n821 B.n26 585
R151 B.n841 B.n26 585
R152 B.n820 B.n819 585
R153 B.n819 B.n22 585
R154 B.n818 B.n21 585
R155 B.n847 B.n21 585
R156 B.n817 B.n20 585
R157 B.n848 B.n20 585
R158 B.n816 B.n19 585
R159 B.n849 B.n19 585
R160 B.n815 B.n814 585
R161 B.n814 B.n15 585
R162 B.n813 B.n14 585
R163 B.n855 B.n14 585
R164 B.n812 B.n13 585
R165 B.n856 B.n13 585
R166 B.n811 B.n12 585
R167 B.n857 B.n12 585
R168 B.n810 B.n809 585
R169 B.n809 B.n11 585
R170 B.n808 B.n7 585
R171 B.n863 B.n7 585
R172 B.n807 B.n6 585
R173 B.n864 B.n6 585
R174 B.n806 B.n5 585
R175 B.n865 B.n5 585
R176 B.n805 B.n804 585
R177 B.n804 B.n4 585
R178 B.n803 B.n378 585
R179 B.n803 B.n802 585
R180 B.n792 B.n379 585
R181 B.n795 B.n379 585
R182 B.n794 B.n793 585
R183 B.n796 B.n794 585
R184 B.n791 B.n383 585
R185 B.n387 B.n383 585
R186 B.n790 B.n789 585
R187 B.n789 B.n788 585
R188 B.n385 B.n384 585
R189 B.n386 B.n385 585
R190 B.n781 B.n780 585
R191 B.n782 B.n781 585
R192 B.n779 B.n392 585
R193 B.n392 B.n391 585
R194 B.n778 B.n777 585
R195 B.n777 B.n776 585
R196 B.n394 B.n393 585
R197 B.n395 B.n394 585
R198 B.n769 B.n768 585
R199 B.n770 B.n769 585
R200 B.n767 B.n399 585
R201 B.n403 B.n399 585
R202 B.n766 B.n765 585
R203 B.n765 B.n764 585
R204 B.n401 B.n400 585
R205 B.n402 B.n401 585
R206 B.n757 B.n756 585
R207 B.n758 B.n757 585
R208 B.n755 B.n408 585
R209 B.n408 B.n407 585
R210 B.n750 B.n749 585
R211 B.n748 B.n478 585
R212 B.n747 B.n477 585
R213 B.n752 B.n477 585
R214 B.n746 B.n745 585
R215 B.n744 B.n743 585
R216 B.n742 B.n741 585
R217 B.n740 B.n739 585
R218 B.n738 B.n737 585
R219 B.n736 B.n735 585
R220 B.n734 B.n733 585
R221 B.n732 B.n731 585
R222 B.n730 B.n729 585
R223 B.n728 B.n727 585
R224 B.n726 B.n725 585
R225 B.n724 B.n723 585
R226 B.n722 B.n721 585
R227 B.n720 B.n719 585
R228 B.n718 B.n717 585
R229 B.n716 B.n715 585
R230 B.n714 B.n713 585
R231 B.n712 B.n711 585
R232 B.n710 B.n709 585
R233 B.n708 B.n707 585
R234 B.n706 B.n705 585
R235 B.n704 B.n703 585
R236 B.n702 B.n701 585
R237 B.n700 B.n699 585
R238 B.n698 B.n697 585
R239 B.n696 B.n695 585
R240 B.n694 B.n693 585
R241 B.n692 B.n691 585
R242 B.n690 B.n689 585
R243 B.n688 B.n687 585
R244 B.n686 B.n685 585
R245 B.n684 B.n683 585
R246 B.n682 B.n681 585
R247 B.n680 B.n679 585
R248 B.n678 B.n677 585
R249 B.n676 B.n675 585
R250 B.n674 B.n673 585
R251 B.n672 B.n671 585
R252 B.n670 B.n669 585
R253 B.n668 B.n667 585
R254 B.n666 B.n665 585
R255 B.n664 B.n663 585
R256 B.n662 B.n661 585
R257 B.n660 B.n659 585
R258 B.n658 B.n657 585
R259 B.n656 B.n655 585
R260 B.n654 B.n653 585
R261 B.n652 B.n651 585
R262 B.n650 B.n649 585
R263 B.n648 B.n647 585
R264 B.n646 B.n645 585
R265 B.n644 B.n643 585
R266 B.n642 B.n641 585
R267 B.n640 B.n639 585
R268 B.n638 B.n637 585
R269 B.n636 B.n635 585
R270 B.n634 B.n633 585
R271 B.n632 B.n631 585
R272 B.n630 B.n629 585
R273 B.n628 B.n627 585
R274 B.n626 B.n625 585
R275 B.n624 B.n623 585
R276 B.n622 B.n621 585
R277 B.n620 B.n619 585
R278 B.n618 B.n617 585
R279 B.n616 B.n615 585
R280 B.n614 B.n613 585
R281 B.n612 B.n611 585
R282 B.n610 B.n609 585
R283 B.n608 B.n607 585
R284 B.n606 B.n605 585
R285 B.n604 B.n603 585
R286 B.n602 B.n601 585
R287 B.n600 B.n599 585
R288 B.n598 B.n597 585
R289 B.n596 B.n595 585
R290 B.n594 B.n593 585
R291 B.n592 B.n591 585
R292 B.n590 B.n589 585
R293 B.n588 B.n587 585
R294 B.n586 B.n585 585
R295 B.n584 B.n583 585
R296 B.n582 B.n581 585
R297 B.n580 B.n579 585
R298 B.n578 B.n577 585
R299 B.n576 B.n575 585
R300 B.n574 B.n573 585
R301 B.n572 B.n571 585
R302 B.n570 B.n569 585
R303 B.n568 B.n567 585
R304 B.n566 B.n565 585
R305 B.n564 B.n563 585
R306 B.n562 B.n561 585
R307 B.n560 B.n559 585
R308 B.n558 B.n557 585
R309 B.n556 B.n555 585
R310 B.n554 B.n553 585
R311 B.n552 B.n551 585
R312 B.n550 B.n549 585
R313 B.n548 B.n547 585
R314 B.n546 B.n545 585
R315 B.n544 B.n543 585
R316 B.n542 B.n541 585
R317 B.n540 B.n539 585
R318 B.n538 B.n537 585
R319 B.n536 B.n535 585
R320 B.n534 B.n533 585
R321 B.n532 B.n531 585
R322 B.n530 B.n529 585
R323 B.n528 B.n527 585
R324 B.n526 B.n525 585
R325 B.n524 B.n523 585
R326 B.n522 B.n521 585
R327 B.n520 B.n519 585
R328 B.n518 B.n517 585
R329 B.n516 B.n515 585
R330 B.n514 B.n513 585
R331 B.n512 B.n511 585
R332 B.n510 B.n509 585
R333 B.n508 B.n507 585
R334 B.n506 B.n505 585
R335 B.n504 B.n503 585
R336 B.n502 B.n501 585
R337 B.n500 B.n499 585
R338 B.n498 B.n497 585
R339 B.n496 B.n495 585
R340 B.n494 B.n493 585
R341 B.n492 B.n491 585
R342 B.n490 B.n489 585
R343 B.n488 B.n487 585
R344 B.n486 B.n485 585
R345 B.n410 B.n409 585
R346 B.n754 B.n753 585
R347 B.n753 B.n752 585
R348 B.n406 B.n405 585
R349 B.n407 B.n406 585
R350 B.n760 B.n759 585
R351 B.n759 B.n758 585
R352 B.n761 B.n404 585
R353 B.n404 B.n402 585
R354 B.n763 B.n762 585
R355 B.n764 B.n763 585
R356 B.n398 B.n397 585
R357 B.n403 B.n398 585
R358 B.n772 B.n771 585
R359 B.n771 B.n770 585
R360 B.n773 B.n396 585
R361 B.n396 B.n395 585
R362 B.n775 B.n774 585
R363 B.n776 B.n775 585
R364 B.n390 B.n389 585
R365 B.n391 B.n390 585
R366 B.n784 B.n783 585
R367 B.n783 B.n782 585
R368 B.n785 B.n388 585
R369 B.n388 B.n386 585
R370 B.n787 B.n786 585
R371 B.n788 B.n787 585
R372 B.n382 B.n381 585
R373 B.n387 B.n382 585
R374 B.n798 B.n797 585
R375 B.n797 B.n796 585
R376 B.n799 B.n380 585
R377 B.n795 B.n380 585
R378 B.n801 B.n800 585
R379 B.n802 B.n801 585
R380 B.n2 B.n0 585
R381 B.n4 B.n2 585
R382 B.n3 B.n1 585
R383 B.n864 B.n3 585
R384 B.n862 B.n861 585
R385 B.n863 B.n862 585
R386 B.n860 B.n8 585
R387 B.n11 B.n8 585
R388 B.n859 B.n858 585
R389 B.n858 B.n857 585
R390 B.n10 B.n9 585
R391 B.n856 B.n10 585
R392 B.n854 B.n853 585
R393 B.n855 B.n854 585
R394 B.n852 B.n16 585
R395 B.n16 B.n15 585
R396 B.n851 B.n850 585
R397 B.n850 B.n849 585
R398 B.n18 B.n17 585
R399 B.n848 B.n18 585
R400 B.n846 B.n845 585
R401 B.n847 B.n846 585
R402 B.n844 B.n23 585
R403 B.n23 B.n22 585
R404 B.n843 B.n842 585
R405 B.n842 B.n841 585
R406 B.n25 B.n24 585
R407 B.n840 B.n25 585
R408 B.n838 B.n837 585
R409 B.n839 B.n838 585
R410 B.n836 B.n30 585
R411 B.n30 B.n29 585
R412 B.n835 B.n834 585
R413 B.n834 B.n833 585
R414 B.n32 B.n31 585
R415 B.n832 B.n32 585
R416 B.n867 B.n866 585
R417 B.n866 B.n865 585
R418 B.n750 B.n406 434.841
R419 B.n107 B.n32 434.841
R420 B.n753 B.n408 434.841
R421 B.n829 B.n34 434.841
R422 B.n831 B.n830 256.663
R423 B.n831 B.n101 256.663
R424 B.n831 B.n100 256.663
R425 B.n831 B.n99 256.663
R426 B.n831 B.n98 256.663
R427 B.n831 B.n97 256.663
R428 B.n831 B.n96 256.663
R429 B.n831 B.n95 256.663
R430 B.n831 B.n94 256.663
R431 B.n831 B.n93 256.663
R432 B.n831 B.n92 256.663
R433 B.n831 B.n91 256.663
R434 B.n831 B.n90 256.663
R435 B.n831 B.n89 256.663
R436 B.n831 B.n88 256.663
R437 B.n831 B.n87 256.663
R438 B.n831 B.n86 256.663
R439 B.n831 B.n85 256.663
R440 B.n831 B.n84 256.663
R441 B.n831 B.n83 256.663
R442 B.n831 B.n82 256.663
R443 B.n831 B.n81 256.663
R444 B.n831 B.n80 256.663
R445 B.n831 B.n79 256.663
R446 B.n831 B.n78 256.663
R447 B.n831 B.n77 256.663
R448 B.n831 B.n76 256.663
R449 B.n831 B.n75 256.663
R450 B.n831 B.n74 256.663
R451 B.n831 B.n73 256.663
R452 B.n831 B.n72 256.663
R453 B.n831 B.n71 256.663
R454 B.n831 B.n70 256.663
R455 B.n831 B.n69 256.663
R456 B.n831 B.n68 256.663
R457 B.n831 B.n67 256.663
R458 B.n831 B.n66 256.663
R459 B.n831 B.n65 256.663
R460 B.n831 B.n64 256.663
R461 B.n831 B.n63 256.663
R462 B.n831 B.n62 256.663
R463 B.n831 B.n61 256.663
R464 B.n831 B.n60 256.663
R465 B.n831 B.n59 256.663
R466 B.n831 B.n58 256.663
R467 B.n831 B.n57 256.663
R468 B.n831 B.n56 256.663
R469 B.n831 B.n55 256.663
R470 B.n831 B.n54 256.663
R471 B.n831 B.n53 256.663
R472 B.n831 B.n52 256.663
R473 B.n831 B.n51 256.663
R474 B.n831 B.n50 256.663
R475 B.n831 B.n49 256.663
R476 B.n831 B.n48 256.663
R477 B.n831 B.n47 256.663
R478 B.n831 B.n46 256.663
R479 B.n831 B.n45 256.663
R480 B.n831 B.n44 256.663
R481 B.n831 B.n43 256.663
R482 B.n831 B.n42 256.663
R483 B.n831 B.n41 256.663
R484 B.n831 B.n40 256.663
R485 B.n831 B.n39 256.663
R486 B.n831 B.n38 256.663
R487 B.n831 B.n37 256.663
R488 B.n831 B.n36 256.663
R489 B.n831 B.n35 256.663
R490 B.n752 B.n751 256.663
R491 B.n752 B.n411 256.663
R492 B.n752 B.n412 256.663
R493 B.n752 B.n413 256.663
R494 B.n752 B.n414 256.663
R495 B.n752 B.n415 256.663
R496 B.n752 B.n416 256.663
R497 B.n752 B.n417 256.663
R498 B.n752 B.n418 256.663
R499 B.n752 B.n419 256.663
R500 B.n752 B.n420 256.663
R501 B.n752 B.n421 256.663
R502 B.n752 B.n422 256.663
R503 B.n752 B.n423 256.663
R504 B.n752 B.n424 256.663
R505 B.n752 B.n425 256.663
R506 B.n752 B.n426 256.663
R507 B.n752 B.n427 256.663
R508 B.n752 B.n428 256.663
R509 B.n752 B.n429 256.663
R510 B.n752 B.n430 256.663
R511 B.n752 B.n431 256.663
R512 B.n752 B.n432 256.663
R513 B.n752 B.n433 256.663
R514 B.n752 B.n434 256.663
R515 B.n752 B.n435 256.663
R516 B.n752 B.n436 256.663
R517 B.n752 B.n437 256.663
R518 B.n752 B.n438 256.663
R519 B.n752 B.n439 256.663
R520 B.n752 B.n440 256.663
R521 B.n752 B.n441 256.663
R522 B.n752 B.n442 256.663
R523 B.n752 B.n443 256.663
R524 B.n752 B.n444 256.663
R525 B.n752 B.n445 256.663
R526 B.n752 B.n446 256.663
R527 B.n752 B.n447 256.663
R528 B.n752 B.n448 256.663
R529 B.n752 B.n449 256.663
R530 B.n752 B.n450 256.663
R531 B.n752 B.n451 256.663
R532 B.n752 B.n452 256.663
R533 B.n752 B.n453 256.663
R534 B.n752 B.n454 256.663
R535 B.n752 B.n455 256.663
R536 B.n752 B.n456 256.663
R537 B.n752 B.n457 256.663
R538 B.n752 B.n458 256.663
R539 B.n752 B.n459 256.663
R540 B.n752 B.n460 256.663
R541 B.n752 B.n461 256.663
R542 B.n752 B.n462 256.663
R543 B.n752 B.n463 256.663
R544 B.n752 B.n464 256.663
R545 B.n752 B.n465 256.663
R546 B.n752 B.n466 256.663
R547 B.n752 B.n467 256.663
R548 B.n752 B.n468 256.663
R549 B.n752 B.n469 256.663
R550 B.n752 B.n470 256.663
R551 B.n752 B.n471 256.663
R552 B.n752 B.n472 256.663
R553 B.n752 B.n473 256.663
R554 B.n752 B.n474 256.663
R555 B.n752 B.n475 256.663
R556 B.n752 B.n476 256.663
R557 B.n759 B.n406 163.367
R558 B.n759 B.n404 163.367
R559 B.n763 B.n404 163.367
R560 B.n763 B.n398 163.367
R561 B.n771 B.n398 163.367
R562 B.n771 B.n396 163.367
R563 B.n775 B.n396 163.367
R564 B.n775 B.n390 163.367
R565 B.n783 B.n390 163.367
R566 B.n783 B.n388 163.367
R567 B.n787 B.n388 163.367
R568 B.n787 B.n382 163.367
R569 B.n797 B.n382 163.367
R570 B.n797 B.n380 163.367
R571 B.n801 B.n380 163.367
R572 B.n801 B.n2 163.367
R573 B.n866 B.n2 163.367
R574 B.n866 B.n3 163.367
R575 B.n862 B.n3 163.367
R576 B.n862 B.n8 163.367
R577 B.n858 B.n8 163.367
R578 B.n858 B.n10 163.367
R579 B.n854 B.n10 163.367
R580 B.n854 B.n16 163.367
R581 B.n850 B.n16 163.367
R582 B.n850 B.n18 163.367
R583 B.n846 B.n18 163.367
R584 B.n846 B.n23 163.367
R585 B.n842 B.n23 163.367
R586 B.n842 B.n25 163.367
R587 B.n838 B.n25 163.367
R588 B.n838 B.n30 163.367
R589 B.n834 B.n30 163.367
R590 B.n834 B.n32 163.367
R591 B.n478 B.n477 163.367
R592 B.n745 B.n477 163.367
R593 B.n743 B.n742 163.367
R594 B.n739 B.n738 163.367
R595 B.n735 B.n734 163.367
R596 B.n731 B.n730 163.367
R597 B.n727 B.n726 163.367
R598 B.n723 B.n722 163.367
R599 B.n719 B.n718 163.367
R600 B.n715 B.n714 163.367
R601 B.n711 B.n710 163.367
R602 B.n707 B.n706 163.367
R603 B.n703 B.n702 163.367
R604 B.n699 B.n698 163.367
R605 B.n695 B.n694 163.367
R606 B.n691 B.n690 163.367
R607 B.n687 B.n686 163.367
R608 B.n683 B.n682 163.367
R609 B.n679 B.n678 163.367
R610 B.n675 B.n674 163.367
R611 B.n671 B.n670 163.367
R612 B.n667 B.n666 163.367
R613 B.n663 B.n662 163.367
R614 B.n659 B.n658 163.367
R615 B.n655 B.n654 163.367
R616 B.n651 B.n650 163.367
R617 B.n647 B.n646 163.367
R618 B.n643 B.n642 163.367
R619 B.n639 B.n638 163.367
R620 B.n635 B.n634 163.367
R621 B.n631 B.n630 163.367
R622 B.n627 B.n626 163.367
R623 B.n623 B.n622 163.367
R624 B.n619 B.n618 163.367
R625 B.n615 B.n614 163.367
R626 B.n611 B.n610 163.367
R627 B.n607 B.n606 163.367
R628 B.n603 B.n602 163.367
R629 B.n599 B.n598 163.367
R630 B.n595 B.n594 163.367
R631 B.n591 B.n590 163.367
R632 B.n587 B.n586 163.367
R633 B.n583 B.n582 163.367
R634 B.n579 B.n578 163.367
R635 B.n575 B.n574 163.367
R636 B.n571 B.n570 163.367
R637 B.n567 B.n566 163.367
R638 B.n563 B.n562 163.367
R639 B.n559 B.n558 163.367
R640 B.n555 B.n554 163.367
R641 B.n551 B.n550 163.367
R642 B.n547 B.n546 163.367
R643 B.n543 B.n542 163.367
R644 B.n539 B.n538 163.367
R645 B.n535 B.n534 163.367
R646 B.n531 B.n530 163.367
R647 B.n527 B.n526 163.367
R648 B.n523 B.n522 163.367
R649 B.n519 B.n518 163.367
R650 B.n515 B.n514 163.367
R651 B.n511 B.n510 163.367
R652 B.n507 B.n506 163.367
R653 B.n503 B.n502 163.367
R654 B.n499 B.n498 163.367
R655 B.n495 B.n494 163.367
R656 B.n491 B.n490 163.367
R657 B.n487 B.n486 163.367
R658 B.n753 B.n410 163.367
R659 B.n757 B.n408 163.367
R660 B.n757 B.n401 163.367
R661 B.n765 B.n401 163.367
R662 B.n765 B.n399 163.367
R663 B.n769 B.n399 163.367
R664 B.n769 B.n394 163.367
R665 B.n777 B.n394 163.367
R666 B.n777 B.n392 163.367
R667 B.n781 B.n392 163.367
R668 B.n781 B.n385 163.367
R669 B.n789 B.n385 163.367
R670 B.n789 B.n383 163.367
R671 B.n794 B.n383 163.367
R672 B.n794 B.n379 163.367
R673 B.n803 B.n379 163.367
R674 B.n804 B.n803 163.367
R675 B.n804 B.n5 163.367
R676 B.n6 B.n5 163.367
R677 B.n7 B.n6 163.367
R678 B.n809 B.n7 163.367
R679 B.n809 B.n12 163.367
R680 B.n13 B.n12 163.367
R681 B.n14 B.n13 163.367
R682 B.n814 B.n14 163.367
R683 B.n814 B.n19 163.367
R684 B.n20 B.n19 163.367
R685 B.n21 B.n20 163.367
R686 B.n819 B.n21 163.367
R687 B.n819 B.n26 163.367
R688 B.n27 B.n26 163.367
R689 B.n28 B.n27 163.367
R690 B.n824 B.n28 163.367
R691 B.n824 B.n33 163.367
R692 B.n34 B.n33 163.367
R693 B.n111 B.n110 163.367
R694 B.n115 B.n114 163.367
R695 B.n119 B.n118 163.367
R696 B.n123 B.n122 163.367
R697 B.n127 B.n126 163.367
R698 B.n131 B.n130 163.367
R699 B.n135 B.n134 163.367
R700 B.n139 B.n138 163.367
R701 B.n143 B.n142 163.367
R702 B.n147 B.n146 163.367
R703 B.n151 B.n150 163.367
R704 B.n155 B.n154 163.367
R705 B.n159 B.n158 163.367
R706 B.n163 B.n162 163.367
R707 B.n167 B.n166 163.367
R708 B.n171 B.n170 163.367
R709 B.n175 B.n174 163.367
R710 B.n179 B.n178 163.367
R711 B.n183 B.n182 163.367
R712 B.n187 B.n186 163.367
R713 B.n191 B.n190 163.367
R714 B.n195 B.n194 163.367
R715 B.n199 B.n198 163.367
R716 B.n203 B.n202 163.367
R717 B.n207 B.n206 163.367
R718 B.n211 B.n210 163.367
R719 B.n215 B.n214 163.367
R720 B.n219 B.n218 163.367
R721 B.n223 B.n222 163.367
R722 B.n227 B.n226 163.367
R723 B.n231 B.n230 163.367
R724 B.n236 B.n235 163.367
R725 B.n240 B.n239 163.367
R726 B.n244 B.n243 163.367
R727 B.n248 B.n247 163.367
R728 B.n252 B.n251 163.367
R729 B.n257 B.n256 163.367
R730 B.n261 B.n260 163.367
R731 B.n265 B.n264 163.367
R732 B.n269 B.n268 163.367
R733 B.n273 B.n272 163.367
R734 B.n277 B.n276 163.367
R735 B.n281 B.n280 163.367
R736 B.n285 B.n284 163.367
R737 B.n289 B.n288 163.367
R738 B.n293 B.n292 163.367
R739 B.n297 B.n296 163.367
R740 B.n301 B.n300 163.367
R741 B.n305 B.n304 163.367
R742 B.n309 B.n308 163.367
R743 B.n313 B.n312 163.367
R744 B.n317 B.n316 163.367
R745 B.n321 B.n320 163.367
R746 B.n325 B.n324 163.367
R747 B.n329 B.n328 163.367
R748 B.n333 B.n332 163.367
R749 B.n337 B.n336 163.367
R750 B.n341 B.n340 163.367
R751 B.n345 B.n344 163.367
R752 B.n349 B.n348 163.367
R753 B.n353 B.n352 163.367
R754 B.n357 B.n356 163.367
R755 B.n361 B.n360 163.367
R756 B.n365 B.n364 163.367
R757 B.n369 B.n368 163.367
R758 B.n373 B.n372 163.367
R759 B.n375 B.n102 163.367
R760 B.n482 B.t12 85.99
R761 B.n103 B.t18 85.99
R762 B.n479 B.t9 85.9643
R763 B.n105 B.t15 85.9643
R764 B.n751 B.n750 71.676
R765 B.n745 B.n411 71.676
R766 B.n742 B.n412 71.676
R767 B.n738 B.n413 71.676
R768 B.n734 B.n414 71.676
R769 B.n730 B.n415 71.676
R770 B.n726 B.n416 71.676
R771 B.n722 B.n417 71.676
R772 B.n718 B.n418 71.676
R773 B.n714 B.n419 71.676
R774 B.n710 B.n420 71.676
R775 B.n706 B.n421 71.676
R776 B.n702 B.n422 71.676
R777 B.n698 B.n423 71.676
R778 B.n694 B.n424 71.676
R779 B.n690 B.n425 71.676
R780 B.n686 B.n426 71.676
R781 B.n682 B.n427 71.676
R782 B.n678 B.n428 71.676
R783 B.n674 B.n429 71.676
R784 B.n670 B.n430 71.676
R785 B.n666 B.n431 71.676
R786 B.n662 B.n432 71.676
R787 B.n658 B.n433 71.676
R788 B.n654 B.n434 71.676
R789 B.n650 B.n435 71.676
R790 B.n646 B.n436 71.676
R791 B.n642 B.n437 71.676
R792 B.n638 B.n438 71.676
R793 B.n634 B.n439 71.676
R794 B.n630 B.n440 71.676
R795 B.n626 B.n441 71.676
R796 B.n622 B.n442 71.676
R797 B.n618 B.n443 71.676
R798 B.n614 B.n444 71.676
R799 B.n610 B.n445 71.676
R800 B.n606 B.n446 71.676
R801 B.n602 B.n447 71.676
R802 B.n598 B.n448 71.676
R803 B.n594 B.n449 71.676
R804 B.n590 B.n450 71.676
R805 B.n586 B.n451 71.676
R806 B.n582 B.n452 71.676
R807 B.n578 B.n453 71.676
R808 B.n574 B.n454 71.676
R809 B.n570 B.n455 71.676
R810 B.n566 B.n456 71.676
R811 B.n562 B.n457 71.676
R812 B.n558 B.n458 71.676
R813 B.n554 B.n459 71.676
R814 B.n550 B.n460 71.676
R815 B.n546 B.n461 71.676
R816 B.n542 B.n462 71.676
R817 B.n538 B.n463 71.676
R818 B.n534 B.n464 71.676
R819 B.n530 B.n465 71.676
R820 B.n526 B.n466 71.676
R821 B.n522 B.n467 71.676
R822 B.n518 B.n468 71.676
R823 B.n514 B.n469 71.676
R824 B.n510 B.n470 71.676
R825 B.n506 B.n471 71.676
R826 B.n502 B.n472 71.676
R827 B.n498 B.n473 71.676
R828 B.n494 B.n474 71.676
R829 B.n490 B.n475 71.676
R830 B.n486 B.n476 71.676
R831 B.n107 B.n35 71.676
R832 B.n111 B.n36 71.676
R833 B.n115 B.n37 71.676
R834 B.n119 B.n38 71.676
R835 B.n123 B.n39 71.676
R836 B.n127 B.n40 71.676
R837 B.n131 B.n41 71.676
R838 B.n135 B.n42 71.676
R839 B.n139 B.n43 71.676
R840 B.n143 B.n44 71.676
R841 B.n147 B.n45 71.676
R842 B.n151 B.n46 71.676
R843 B.n155 B.n47 71.676
R844 B.n159 B.n48 71.676
R845 B.n163 B.n49 71.676
R846 B.n167 B.n50 71.676
R847 B.n171 B.n51 71.676
R848 B.n175 B.n52 71.676
R849 B.n179 B.n53 71.676
R850 B.n183 B.n54 71.676
R851 B.n187 B.n55 71.676
R852 B.n191 B.n56 71.676
R853 B.n195 B.n57 71.676
R854 B.n199 B.n58 71.676
R855 B.n203 B.n59 71.676
R856 B.n207 B.n60 71.676
R857 B.n211 B.n61 71.676
R858 B.n215 B.n62 71.676
R859 B.n219 B.n63 71.676
R860 B.n223 B.n64 71.676
R861 B.n227 B.n65 71.676
R862 B.n231 B.n66 71.676
R863 B.n236 B.n67 71.676
R864 B.n240 B.n68 71.676
R865 B.n244 B.n69 71.676
R866 B.n248 B.n70 71.676
R867 B.n252 B.n71 71.676
R868 B.n257 B.n72 71.676
R869 B.n261 B.n73 71.676
R870 B.n265 B.n74 71.676
R871 B.n269 B.n75 71.676
R872 B.n273 B.n76 71.676
R873 B.n277 B.n77 71.676
R874 B.n281 B.n78 71.676
R875 B.n285 B.n79 71.676
R876 B.n289 B.n80 71.676
R877 B.n293 B.n81 71.676
R878 B.n297 B.n82 71.676
R879 B.n301 B.n83 71.676
R880 B.n305 B.n84 71.676
R881 B.n309 B.n85 71.676
R882 B.n313 B.n86 71.676
R883 B.n317 B.n87 71.676
R884 B.n321 B.n88 71.676
R885 B.n325 B.n89 71.676
R886 B.n329 B.n90 71.676
R887 B.n333 B.n91 71.676
R888 B.n337 B.n92 71.676
R889 B.n341 B.n93 71.676
R890 B.n345 B.n94 71.676
R891 B.n349 B.n95 71.676
R892 B.n353 B.n96 71.676
R893 B.n357 B.n97 71.676
R894 B.n361 B.n98 71.676
R895 B.n365 B.n99 71.676
R896 B.n369 B.n100 71.676
R897 B.n373 B.n101 71.676
R898 B.n830 B.n102 71.676
R899 B.n830 B.n829 71.676
R900 B.n375 B.n101 71.676
R901 B.n372 B.n100 71.676
R902 B.n368 B.n99 71.676
R903 B.n364 B.n98 71.676
R904 B.n360 B.n97 71.676
R905 B.n356 B.n96 71.676
R906 B.n352 B.n95 71.676
R907 B.n348 B.n94 71.676
R908 B.n344 B.n93 71.676
R909 B.n340 B.n92 71.676
R910 B.n336 B.n91 71.676
R911 B.n332 B.n90 71.676
R912 B.n328 B.n89 71.676
R913 B.n324 B.n88 71.676
R914 B.n320 B.n87 71.676
R915 B.n316 B.n86 71.676
R916 B.n312 B.n85 71.676
R917 B.n308 B.n84 71.676
R918 B.n304 B.n83 71.676
R919 B.n300 B.n82 71.676
R920 B.n296 B.n81 71.676
R921 B.n292 B.n80 71.676
R922 B.n288 B.n79 71.676
R923 B.n284 B.n78 71.676
R924 B.n280 B.n77 71.676
R925 B.n276 B.n76 71.676
R926 B.n272 B.n75 71.676
R927 B.n268 B.n74 71.676
R928 B.n264 B.n73 71.676
R929 B.n260 B.n72 71.676
R930 B.n256 B.n71 71.676
R931 B.n251 B.n70 71.676
R932 B.n247 B.n69 71.676
R933 B.n243 B.n68 71.676
R934 B.n239 B.n67 71.676
R935 B.n235 B.n66 71.676
R936 B.n230 B.n65 71.676
R937 B.n226 B.n64 71.676
R938 B.n222 B.n63 71.676
R939 B.n218 B.n62 71.676
R940 B.n214 B.n61 71.676
R941 B.n210 B.n60 71.676
R942 B.n206 B.n59 71.676
R943 B.n202 B.n58 71.676
R944 B.n198 B.n57 71.676
R945 B.n194 B.n56 71.676
R946 B.n190 B.n55 71.676
R947 B.n186 B.n54 71.676
R948 B.n182 B.n53 71.676
R949 B.n178 B.n52 71.676
R950 B.n174 B.n51 71.676
R951 B.n170 B.n50 71.676
R952 B.n166 B.n49 71.676
R953 B.n162 B.n48 71.676
R954 B.n158 B.n47 71.676
R955 B.n154 B.n46 71.676
R956 B.n150 B.n45 71.676
R957 B.n146 B.n44 71.676
R958 B.n142 B.n43 71.676
R959 B.n138 B.n42 71.676
R960 B.n134 B.n41 71.676
R961 B.n130 B.n40 71.676
R962 B.n126 B.n39 71.676
R963 B.n122 B.n38 71.676
R964 B.n118 B.n37 71.676
R965 B.n114 B.n36 71.676
R966 B.n110 B.n35 71.676
R967 B.n751 B.n478 71.676
R968 B.n743 B.n411 71.676
R969 B.n739 B.n412 71.676
R970 B.n735 B.n413 71.676
R971 B.n731 B.n414 71.676
R972 B.n727 B.n415 71.676
R973 B.n723 B.n416 71.676
R974 B.n719 B.n417 71.676
R975 B.n715 B.n418 71.676
R976 B.n711 B.n419 71.676
R977 B.n707 B.n420 71.676
R978 B.n703 B.n421 71.676
R979 B.n699 B.n422 71.676
R980 B.n695 B.n423 71.676
R981 B.n691 B.n424 71.676
R982 B.n687 B.n425 71.676
R983 B.n683 B.n426 71.676
R984 B.n679 B.n427 71.676
R985 B.n675 B.n428 71.676
R986 B.n671 B.n429 71.676
R987 B.n667 B.n430 71.676
R988 B.n663 B.n431 71.676
R989 B.n659 B.n432 71.676
R990 B.n655 B.n433 71.676
R991 B.n651 B.n434 71.676
R992 B.n647 B.n435 71.676
R993 B.n643 B.n436 71.676
R994 B.n639 B.n437 71.676
R995 B.n635 B.n438 71.676
R996 B.n631 B.n439 71.676
R997 B.n627 B.n440 71.676
R998 B.n623 B.n441 71.676
R999 B.n619 B.n442 71.676
R1000 B.n615 B.n443 71.676
R1001 B.n611 B.n444 71.676
R1002 B.n607 B.n445 71.676
R1003 B.n603 B.n446 71.676
R1004 B.n599 B.n447 71.676
R1005 B.n595 B.n448 71.676
R1006 B.n591 B.n449 71.676
R1007 B.n587 B.n450 71.676
R1008 B.n583 B.n451 71.676
R1009 B.n579 B.n452 71.676
R1010 B.n575 B.n453 71.676
R1011 B.n571 B.n454 71.676
R1012 B.n567 B.n455 71.676
R1013 B.n563 B.n456 71.676
R1014 B.n559 B.n457 71.676
R1015 B.n555 B.n458 71.676
R1016 B.n551 B.n459 71.676
R1017 B.n547 B.n460 71.676
R1018 B.n543 B.n461 71.676
R1019 B.n539 B.n462 71.676
R1020 B.n535 B.n463 71.676
R1021 B.n531 B.n464 71.676
R1022 B.n527 B.n465 71.676
R1023 B.n523 B.n466 71.676
R1024 B.n519 B.n467 71.676
R1025 B.n515 B.n468 71.676
R1026 B.n511 B.n469 71.676
R1027 B.n507 B.n470 71.676
R1028 B.n503 B.n471 71.676
R1029 B.n499 B.n472 71.676
R1030 B.n495 B.n473 71.676
R1031 B.n491 B.n474 71.676
R1032 B.n487 B.n475 71.676
R1033 B.n476 B.n410 71.676
R1034 B.n483 B.t11 71.6385
R1035 B.n104 B.t19 71.6385
R1036 B.n480 B.t8 71.6128
R1037 B.n106 B.t16 71.6128
R1038 B.n484 B.n483 59.5399
R1039 B.n481 B.n480 59.5399
R1040 B.n233 B.n106 59.5399
R1041 B.n254 B.n104 59.5399
R1042 B.n752 B.n407 49.7459
R1043 B.n832 B.n831 49.7459
R1044 B.n758 B.n407 30.4751
R1045 B.n758 B.n402 30.4751
R1046 B.n764 B.n402 30.4751
R1047 B.n764 B.n403 30.4751
R1048 B.n770 B.n395 30.4751
R1049 B.n776 B.n395 30.4751
R1050 B.n776 B.n391 30.4751
R1051 B.n782 B.n391 30.4751
R1052 B.n788 B.n386 30.4751
R1053 B.n788 B.n387 30.4751
R1054 B.n796 B.n795 30.4751
R1055 B.n802 B.n4 30.4751
R1056 B.n865 B.n4 30.4751
R1057 B.n865 B.n864 30.4751
R1058 B.n864 B.n863 30.4751
R1059 B.n857 B.n11 30.4751
R1060 B.n856 B.n855 30.4751
R1061 B.n855 B.n15 30.4751
R1062 B.n849 B.n848 30.4751
R1063 B.n848 B.n847 30.4751
R1064 B.n847 B.n22 30.4751
R1065 B.n841 B.n22 30.4751
R1066 B.n840 B.n839 30.4751
R1067 B.n839 B.n29 30.4751
R1068 B.n833 B.n29 30.4751
R1069 B.n833 B.n832 30.4751
R1070 B.n782 B.t1 29.1307
R1071 B.n849 B.t2 29.1307
R1072 B.n108 B.n31 28.2542
R1073 B.n828 B.n827 28.2542
R1074 B.n755 B.n754 28.2542
R1075 B.n749 B.n405 28.2542
R1076 B.n796 B.t5 26.4417
R1077 B.n857 B.t0 26.4417
R1078 B.n802 B.t3 21.0639
R1079 B.n863 B.t4 21.0639
R1080 B B.n867 18.0485
R1081 B.n403 B.t7 17.4786
R1082 B.t14 B.n840 17.4786
R1083 B.n483 B.n482 14.352
R1084 B.n480 B.n479 14.352
R1085 B.n106 B.n105 14.352
R1086 B.n104 B.n103 14.352
R1087 B.n770 B.t7 12.997
R1088 B.n841 B.t14 12.997
R1089 B.n109 B.n108 10.6151
R1090 B.n112 B.n109 10.6151
R1091 B.n113 B.n112 10.6151
R1092 B.n116 B.n113 10.6151
R1093 B.n117 B.n116 10.6151
R1094 B.n120 B.n117 10.6151
R1095 B.n121 B.n120 10.6151
R1096 B.n124 B.n121 10.6151
R1097 B.n125 B.n124 10.6151
R1098 B.n128 B.n125 10.6151
R1099 B.n129 B.n128 10.6151
R1100 B.n132 B.n129 10.6151
R1101 B.n133 B.n132 10.6151
R1102 B.n136 B.n133 10.6151
R1103 B.n137 B.n136 10.6151
R1104 B.n140 B.n137 10.6151
R1105 B.n141 B.n140 10.6151
R1106 B.n144 B.n141 10.6151
R1107 B.n145 B.n144 10.6151
R1108 B.n148 B.n145 10.6151
R1109 B.n149 B.n148 10.6151
R1110 B.n152 B.n149 10.6151
R1111 B.n153 B.n152 10.6151
R1112 B.n156 B.n153 10.6151
R1113 B.n157 B.n156 10.6151
R1114 B.n160 B.n157 10.6151
R1115 B.n161 B.n160 10.6151
R1116 B.n164 B.n161 10.6151
R1117 B.n165 B.n164 10.6151
R1118 B.n168 B.n165 10.6151
R1119 B.n169 B.n168 10.6151
R1120 B.n172 B.n169 10.6151
R1121 B.n173 B.n172 10.6151
R1122 B.n176 B.n173 10.6151
R1123 B.n177 B.n176 10.6151
R1124 B.n180 B.n177 10.6151
R1125 B.n181 B.n180 10.6151
R1126 B.n184 B.n181 10.6151
R1127 B.n185 B.n184 10.6151
R1128 B.n188 B.n185 10.6151
R1129 B.n189 B.n188 10.6151
R1130 B.n192 B.n189 10.6151
R1131 B.n193 B.n192 10.6151
R1132 B.n196 B.n193 10.6151
R1133 B.n197 B.n196 10.6151
R1134 B.n200 B.n197 10.6151
R1135 B.n201 B.n200 10.6151
R1136 B.n204 B.n201 10.6151
R1137 B.n205 B.n204 10.6151
R1138 B.n208 B.n205 10.6151
R1139 B.n209 B.n208 10.6151
R1140 B.n212 B.n209 10.6151
R1141 B.n213 B.n212 10.6151
R1142 B.n216 B.n213 10.6151
R1143 B.n217 B.n216 10.6151
R1144 B.n220 B.n217 10.6151
R1145 B.n221 B.n220 10.6151
R1146 B.n224 B.n221 10.6151
R1147 B.n225 B.n224 10.6151
R1148 B.n228 B.n225 10.6151
R1149 B.n229 B.n228 10.6151
R1150 B.n232 B.n229 10.6151
R1151 B.n237 B.n234 10.6151
R1152 B.n238 B.n237 10.6151
R1153 B.n241 B.n238 10.6151
R1154 B.n242 B.n241 10.6151
R1155 B.n245 B.n242 10.6151
R1156 B.n246 B.n245 10.6151
R1157 B.n249 B.n246 10.6151
R1158 B.n250 B.n249 10.6151
R1159 B.n253 B.n250 10.6151
R1160 B.n258 B.n255 10.6151
R1161 B.n259 B.n258 10.6151
R1162 B.n262 B.n259 10.6151
R1163 B.n263 B.n262 10.6151
R1164 B.n266 B.n263 10.6151
R1165 B.n267 B.n266 10.6151
R1166 B.n270 B.n267 10.6151
R1167 B.n271 B.n270 10.6151
R1168 B.n274 B.n271 10.6151
R1169 B.n275 B.n274 10.6151
R1170 B.n278 B.n275 10.6151
R1171 B.n279 B.n278 10.6151
R1172 B.n282 B.n279 10.6151
R1173 B.n283 B.n282 10.6151
R1174 B.n286 B.n283 10.6151
R1175 B.n287 B.n286 10.6151
R1176 B.n290 B.n287 10.6151
R1177 B.n291 B.n290 10.6151
R1178 B.n294 B.n291 10.6151
R1179 B.n295 B.n294 10.6151
R1180 B.n298 B.n295 10.6151
R1181 B.n299 B.n298 10.6151
R1182 B.n302 B.n299 10.6151
R1183 B.n303 B.n302 10.6151
R1184 B.n306 B.n303 10.6151
R1185 B.n307 B.n306 10.6151
R1186 B.n310 B.n307 10.6151
R1187 B.n311 B.n310 10.6151
R1188 B.n314 B.n311 10.6151
R1189 B.n315 B.n314 10.6151
R1190 B.n318 B.n315 10.6151
R1191 B.n319 B.n318 10.6151
R1192 B.n322 B.n319 10.6151
R1193 B.n323 B.n322 10.6151
R1194 B.n326 B.n323 10.6151
R1195 B.n327 B.n326 10.6151
R1196 B.n330 B.n327 10.6151
R1197 B.n331 B.n330 10.6151
R1198 B.n334 B.n331 10.6151
R1199 B.n335 B.n334 10.6151
R1200 B.n338 B.n335 10.6151
R1201 B.n339 B.n338 10.6151
R1202 B.n342 B.n339 10.6151
R1203 B.n343 B.n342 10.6151
R1204 B.n346 B.n343 10.6151
R1205 B.n347 B.n346 10.6151
R1206 B.n350 B.n347 10.6151
R1207 B.n351 B.n350 10.6151
R1208 B.n354 B.n351 10.6151
R1209 B.n355 B.n354 10.6151
R1210 B.n358 B.n355 10.6151
R1211 B.n359 B.n358 10.6151
R1212 B.n362 B.n359 10.6151
R1213 B.n363 B.n362 10.6151
R1214 B.n366 B.n363 10.6151
R1215 B.n367 B.n366 10.6151
R1216 B.n370 B.n367 10.6151
R1217 B.n371 B.n370 10.6151
R1218 B.n374 B.n371 10.6151
R1219 B.n376 B.n374 10.6151
R1220 B.n377 B.n376 10.6151
R1221 B.n828 B.n377 10.6151
R1222 B.n756 B.n755 10.6151
R1223 B.n756 B.n400 10.6151
R1224 B.n766 B.n400 10.6151
R1225 B.n767 B.n766 10.6151
R1226 B.n768 B.n767 10.6151
R1227 B.n768 B.n393 10.6151
R1228 B.n778 B.n393 10.6151
R1229 B.n779 B.n778 10.6151
R1230 B.n780 B.n779 10.6151
R1231 B.n780 B.n384 10.6151
R1232 B.n790 B.n384 10.6151
R1233 B.n791 B.n790 10.6151
R1234 B.n793 B.n791 10.6151
R1235 B.n793 B.n792 10.6151
R1236 B.n792 B.n378 10.6151
R1237 B.n805 B.n378 10.6151
R1238 B.n806 B.n805 10.6151
R1239 B.n807 B.n806 10.6151
R1240 B.n808 B.n807 10.6151
R1241 B.n810 B.n808 10.6151
R1242 B.n811 B.n810 10.6151
R1243 B.n812 B.n811 10.6151
R1244 B.n813 B.n812 10.6151
R1245 B.n815 B.n813 10.6151
R1246 B.n816 B.n815 10.6151
R1247 B.n817 B.n816 10.6151
R1248 B.n818 B.n817 10.6151
R1249 B.n820 B.n818 10.6151
R1250 B.n821 B.n820 10.6151
R1251 B.n822 B.n821 10.6151
R1252 B.n823 B.n822 10.6151
R1253 B.n825 B.n823 10.6151
R1254 B.n826 B.n825 10.6151
R1255 B.n827 B.n826 10.6151
R1256 B.n749 B.n748 10.6151
R1257 B.n748 B.n747 10.6151
R1258 B.n747 B.n746 10.6151
R1259 B.n746 B.n744 10.6151
R1260 B.n744 B.n741 10.6151
R1261 B.n741 B.n740 10.6151
R1262 B.n740 B.n737 10.6151
R1263 B.n737 B.n736 10.6151
R1264 B.n736 B.n733 10.6151
R1265 B.n733 B.n732 10.6151
R1266 B.n732 B.n729 10.6151
R1267 B.n729 B.n728 10.6151
R1268 B.n728 B.n725 10.6151
R1269 B.n725 B.n724 10.6151
R1270 B.n724 B.n721 10.6151
R1271 B.n721 B.n720 10.6151
R1272 B.n720 B.n717 10.6151
R1273 B.n717 B.n716 10.6151
R1274 B.n716 B.n713 10.6151
R1275 B.n713 B.n712 10.6151
R1276 B.n712 B.n709 10.6151
R1277 B.n709 B.n708 10.6151
R1278 B.n708 B.n705 10.6151
R1279 B.n705 B.n704 10.6151
R1280 B.n704 B.n701 10.6151
R1281 B.n701 B.n700 10.6151
R1282 B.n700 B.n697 10.6151
R1283 B.n697 B.n696 10.6151
R1284 B.n696 B.n693 10.6151
R1285 B.n693 B.n692 10.6151
R1286 B.n692 B.n689 10.6151
R1287 B.n689 B.n688 10.6151
R1288 B.n688 B.n685 10.6151
R1289 B.n685 B.n684 10.6151
R1290 B.n684 B.n681 10.6151
R1291 B.n681 B.n680 10.6151
R1292 B.n680 B.n677 10.6151
R1293 B.n677 B.n676 10.6151
R1294 B.n676 B.n673 10.6151
R1295 B.n673 B.n672 10.6151
R1296 B.n672 B.n669 10.6151
R1297 B.n669 B.n668 10.6151
R1298 B.n668 B.n665 10.6151
R1299 B.n665 B.n664 10.6151
R1300 B.n664 B.n661 10.6151
R1301 B.n661 B.n660 10.6151
R1302 B.n660 B.n657 10.6151
R1303 B.n657 B.n656 10.6151
R1304 B.n656 B.n653 10.6151
R1305 B.n653 B.n652 10.6151
R1306 B.n652 B.n649 10.6151
R1307 B.n649 B.n648 10.6151
R1308 B.n648 B.n645 10.6151
R1309 B.n645 B.n644 10.6151
R1310 B.n644 B.n641 10.6151
R1311 B.n641 B.n640 10.6151
R1312 B.n640 B.n637 10.6151
R1313 B.n637 B.n636 10.6151
R1314 B.n636 B.n633 10.6151
R1315 B.n633 B.n632 10.6151
R1316 B.n632 B.n629 10.6151
R1317 B.n629 B.n628 10.6151
R1318 B.n625 B.n624 10.6151
R1319 B.n624 B.n621 10.6151
R1320 B.n621 B.n620 10.6151
R1321 B.n620 B.n617 10.6151
R1322 B.n617 B.n616 10.6151
R1323 B.n616 B.n613 10.6151
R1324 B.n613 B.n612 10.6151
R1325 B.n612 B.n609 10.6151
R1326 B.n609 B.n608 10.6151
R1327 B.n605 B.n604 10.6151
R1328 B.n604 B.n601 10.6151
R1329 B.n601 B.n600 10.6151
R1330 B.n600 B.n597 10.6151
R1331 B.n597 B.n596 10.6151
R1332 B.n596 B.n593 10.6151
R1333 B.n593 B.n592 10.6151
R1334 B.n592 B.n589 10.6151
R1335 B.n589 B.n588 10.6151
R1336 B.n588 B.n585 10.6151
R1337 B.n585 B.n584 10.6151
R1338 B.n584 B.n581 10.6151
R1339 B.n581 B.n580 10.6151
R1340 B.n580 B.n577 10.6151
R1341 B.n577 B.n576 10.6151
R1342 B.n576 B.n573 10.6151
R1343 B.n573 B.n572 10.6151
R1344 B.n572 B.n569 10.6151
R1345 B.n569 B.n568 10.6151
R1346 B.n568 B.n565 10.6151
R1347 B.n565 B.n564 10.6151
R1348 B.n564 B.n561 10.6151
R1349 B.n561 B.n560 10.6151
R1350 B.n560 B.n557 10.6151
R1351 B.n557 B.n556 10.6151
R1352 B.n556 B.n553 10.6151
R1353 B.n553 B.n552 10.6151
R1354 B.n552 B.n549 10.6151
R1355 B.n549 B.n548 10.6151
R1356 B.n548 B.n545 10.6151
R1357 B.n545 B.n544 10.6151
R1358 B.n544 B.n541 10.6151
R1359 B.n541 B.n540 10.6151
R1360 B.n540 B.n537 10.6151
R1361 B.n537 B.n536 10.6151
R1362 B.n536 B.n533 10.6151
R1363 B.n533 B.n532 10.6151
R1364 B.n532 B.n529 10.6151
R1365 B.n529 B.n528 10.6151
R1366 B.n528 B.n525 10.6151
R1367 B.n525 B.n524 10.6151
R1368 B.n524 B.n521 10.6151
R1369 B.n521 B.n520 10.6151
R1370 B.n520 B.n517 10.6151
R1371 B.n517 B.n516 10.6151
R1372 B.n516 B.n513 10.6151
R1373 B.n513 B.n512 10.6151
R1374 B.n512 B.n509 10.6151
R1375 B.n509 B.n508 10.6151
R1376 B.n508 B.n505 10.6151
R1377 B.n505 B.n504 10.6151
R1378 B.n504 B.n501 10.6151
R1379 B.n501 B.n500 10.6151
R1380 B.n500 B.n497 10.6151
R1381 B.n497 B.n496 10.6151
R1382 B.n496 B.n493 10.6151
R1383 B.n493 B.n492 10.6151
R1384 B.n492 B.n489 10.6151
R1385 B.n489 B.n488 10.6151
R1386 B.n488 B.n485 10.6151
R1387 B.n485 B.n409 10.6151
R1388 B.n754 B.n409 10.6151
R1389 B.n760 B.n405 10.6151
R1390 B.n761 B.n760 10.6151
R1391 B.n762 B.n761 10.6151
R1392 B.n762 B.n397 10.6151
R1393 B.n772 B.n397 10.6151
R1394 B.n773 B.n772 10.6151
R1395 B.n774 B.n773 10.6151
R1396 B.n774 B.n389 10.6151
R1397 B.n784 B.n389 10.6151
R1398 B.n785 B.n784 10.6151
R1399 B.n786 B.n785 10.6151
R1400 B.n786 B.n381 10.6151
R1401 B.n798 B.n381 10.6151
R1402 B.n799 B.n798 10.6151
R1403 B.n800 B.n799 10.6151
R1404 B.n800 B.n0 10.6151
R1405 B.n861 B.n1 10.6151
R1406 B.n861 B.n860 10.6151
R1407 B.n860 B.n859 10.6151
R1408 B.n859 B.n9 10.6151
R1409 B.n853 B.n9 10.6151
R1410 B.n853 B.n852 10.6151
R1411 B.n852 B.n851 10.6151
R1412 B.n851 B.n17 10.6151
R1413 B.n845 B.n17 10.6151
R1414 B.n845 B.n844 10.6151
R1415 B.n844 B.n843 10.6151
R1416 B.n843 B.n24 10.6151
R1417 B.n837 B.n24 10.6151
R1418 B.n837 B.n836 10.6151
R1419 B.n836 B.n835 10.6151
R1420 B.n835 B.n31 10.6151
R1421 B.n795 B.t3 9.41179
R1422 B.n11 B.t4 9.41179
R1423 B.n233 B.n232 9.36635
R1424 B.n255 B.n254 9.36635
R1425 B.n628 B.n481 9.36635
R1426 B.n605 B.n484 9.36635
R1427 B.n387 B.t5 4.03391
R1428 B.t0 B.n856 4.03391
R1429 B.n867 B.n0 2.81026
R1430 B.n867 B.n1 2.81026
R1431 B.t1 B.n386 1.34497
R1432 B.t2 B.n15 1.34497
R1433 B.n234 B.n233 1.24928
R1434 B.n254 B.n253 1.24928
R1435 B.n625 B.n481 1.24928
R1436 B.n608 B.n484 1.24928
R1437 VN.n0 VN.t1 1253.23
R1438 VN.n4 VN.t2 1253.23
R1439 VN.n2 VN.t4 1234.21
R1440 VN.n6 VN.t0 1234.21
R1441 VN.n1 VN.t5 1229.1
R1442 VN.n5 VN.t3 1229.1
R1443 VN.n3 VN.n2 161.3
R1444 VN.n7 VN.n6 161.3
R1445 VN.n7 VN.n4 71.3843
R1446 VN.n3 VN.n0 71.3843
R1447 VN VN.n7 46.0403
R1448 VN.n2 VN.n1 43.0884
R1449 VN.n6 VN.n5 43.0884
R1450 VN.n5 VN.n4 18.9966
R1451 VN.n1 VN.n0 18.9966
R1452 VN VN.n3 0.0516364
R1453 VTAIL.n7 VTAIL.t10 43.9902
R1454 VTAIL.n11 VTAIL.t11 43.9899
R1455 VTAIL.n2 VTAIL.t1 43.9899
R1456 VTAIL.n10 VTAIL.t4 43.9899
R1457 VTAIL.n9 VTAIL.n8 42.9627
R1458 VTAIL.n6 VTAIL.n5 42.9627
R1459 VTAIL.n1 VTAIL.n0 42.9626
R1460 VTAIL.n4 VTAIL.n3 42.9626
R1461 VTAIL.n6 VTAIL.n4 30.2548
R1462 VTAIL.n11 VTAIL.n10 29.6169
R1463 VTAIL.n0 VTAIL.t9 1.028
R1464 VTAIL.n0 VTAIL.t7 1.028
R1465 VTAIL.n3 VTAIL.t3 1.028
R1466 VTAIL.n3 VTAIL.t2 1.028
R1467 VTAIL.n8 VTAIL.t0 1.028
R1468 VTAIL.n8 VTAIL.t5 1.028
R1469 VTAIL.n5 VTAIL.t8 1.028
R1470 VTAIL.n5 VTAIL.t6 1.028
R1471 VTAIL.n9 VTAIL.n7 0.789293
R1472 VTAIL.n2 VTAIL.n1 0.789293
R1473 VTAIL.n7 VTAIL.n6 0.638431
R1474 VTAIL.n10 VTAIL.n9 0.638431
R1475 VTAIL.n4 VTAIL.n2 0.638431
R1476 VTAIL VTAIL.n11 0.420759
R1477 VTAIL VTAIL.n1 0.218172
R1478 VDD2.n1 VDD2.t4 61.0918
R1479 VDD2.n2 VDD2.t5 60.6689
R1480 VDD2.n1 VDD2.n0 59.7455
R1481 VDD2 VDD2.n3 59.7426
R1482 VDD2.n2 VDD2.n1 42.4006
R1483 VDD2.n3 VDD2.t2 1.028
R1484 VDD2.n3 VDD2.t3 1.028
R1485 VDD2.n0 VDD2.t0 1.028
R1486 VDD2.n0 VDD2.t1 1.028
R1487 VDD2 VDD2.n2 0.537138
R1488 VP.n1 VP.t0 1253.23
R1489 VP.n8 VP.t3 1234.21
R1490 VP.n6 VP.t4 1234.21
R1491 VP.n3 VP.t2 1234.21
R1492 VP.n7 VP.t5 1229.1
R1493 VP.n2 VP.t1 1229.1
R1494 VP.n9 VP.n8 161.3
R1495 VP.n4 VP.n3 161.3
R1496 VP.n7 VP.n0 161.3
R1497 VP.n6 VP.n5 161.3
R1498 VP.n4 VP.n1 71.3843
R1499 VP.n5 VP.n4 45.6596
R1500 VP.n7 VP.n6 43.0884
R1501 VP.n8 VP.n7 43.0884
R1502 VP.n3 VP.n2 43.0884
R1503 VP.n2 VP.n1 18.9966
R1504 VP.n5 VP.n0 0.189894
R1505 VP.n9 VP.n0 0.189894
R1506 VP VP.n9 0.0516364
R1507 VDD1 VDD1.t5 61.2056
R1508 VDD1.n1 VDD1.t1 61.0918
R1509 VDD1.n1 VDD1.n0 59.7455
R1510 VDD1.n3 VDD1.n2 59.6413
R1511 VDD1.n3 VDD1.n1 43.3026
R1512 VDD1.n2 VDD1.t4 1.028
R1513 VDD1.n2 VDD1.t3 1.028
R1514 VDD1.n0 VDD1.t0 1.028
R1515 VDD1.n0 VDD1.t2 1.028
R1516 VDD1 VDD1.n3 0.101793
C0 VTAIL VN 4.31972f
C1 VN VDD2 5.0321f
C2 VP VN 6.14418f
C3 VDD1 VN 0.147729f
C4 VTAIL VDD2 18.7309f
C5 VP VTAIL 4.3348f
C6 VP VDD2 0.274429f
C7 VDD1 VTAIL 18.7049f
C8 VDD1 VDD2 0.610498f
C9 VP VDD1 5.15098f
C10 VDD2 B 5.585059f
C11 VDD1 B 5.800718f
C12 VTAIL B 8.680893f
C13 VN B 8.0356f
C14 VP B 5.379718f
C15 VDD1.t5 B 4.62537f
C16 VDD1.t1 B 4.62467f
C17 VDD1.t0 B 0.395999f
C18 VDD1.t2 B 0.395999f
C19 VDD1.n0 B 3.61567f
C20 VDD1.n1 B 2.59319f
C21 VDD1.t4 B 0.395999f
C22 VDD1.t3 B 0.395999f
C23 VDD1.n2 B 3.61513f
C24 VDD1.n3 B 2.84429f
C25 VP.n0 B 0.054649f
C26 VP.t4 B 1.22527f
C27 VP.t0 B 1.2323f
C28 VP.n1 B 0.456553f
C29 VP.t1 B 1.2234f
C30 VP.n2 B 0.472635f
C31 VP.t2 B 1.22527f
C32 VP.n3 B 0.463179f
C33 VP.n4 B 2.70515f
C34 VP.n5 B 2.62614f
C35 VP.n6 B 0.463179f
C36 VP.t5 B 1.2234f
C37 VP.n7 B 0.472635f
C38 VP.t3 B 1.22527f
C39 VP.n8 B 0.463179f
C40 VP.n9 B 0.042351f
C41 VDD2.t4 B 4.60448f
C42 VDD2.t0 B 0.39427f
C43 VDD2.t1 B 0.39427f
C44 VDD2.n0 B 3.59988f
C45 VDD2.n1 B 2.50761f
C46 VDD2.t5 B 4.60214f
C47 VDD2.n2 B 2.86607f
C48 VDD2.t2 B 0.39427f
C49 VDD2.t3 B 0.39427f
C50 VDD2.n3 B 3.59983f
C51 VTAIL.t9 B 0.397102f
C52 VTAIL.t7 B 0.397102f
C53 VTAIL.n0 B 3.54188f
C54 VTAIL.n1 B 0.352091f
C55 VTAIL.t1 B 4.52612f
C56 VTAIL.n2 B 0.48617f
C57 VTAIL.t3 B 0.397102f
C58 VTAIL.t2 B 0.397102f
C59 VTAIL.n3 B 3.54188f
C60 VTAIL.n4 B 2.17844f
C61 VTAIL.t8 B 0.397102f
C62 VTAIL.t6 B 0.397102f
C63 VTAIL.n5 B 3.54187f
C64 VTAIL.n6 B 2.17845f
C65 VTAIL.t10 B 4.52612f
C66 VTAIL.n7 B 0.486164f
C67 VTAIL.t0 B 0.397102f
C68 VTAIL.t5 B 0.397102f
C69 VTAIL.n8 B 3.54187f
C70 VTAIL.n9 B 0.387413f
C71 VTAIL.t4 B 4.52612f
C72 VTAIL.n10 B 2.2236f
C73 VTAIL.t11 B 4.52612f
C74 VTAIL.n11 B 2.20531f
C75 VN.t1 B 1.21054f
C76 VN.n0 B 0.448491f
C77 VN.t5 B 1.20179f
C78 VN.n1 B 0.464289f
C79 VN.t4 B 1.20363f
C80 VN.n2 B 0.455f
C81 VN.n3 B 0.161481f
C82 VN.t2 B 1.21054f
C83 VN.n4 B 0.448491f
C84 VN.t0 B 1.20363f
C85 VN.t3 B 1.20179f
C86 VN.n5 B 0.464289f
C87 VN.n6 B 0.455f
C88 VN.n7 B 2.69246f
.ends

