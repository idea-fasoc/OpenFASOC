* NGSPICE file created from diff_pair_sample_0006.ext - technology: sky130A

.subckt diff_pair_sample_0006 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=7.215 pd=37.78 as=0 ps=0 w=18.5 l=3.53
X1 B.t12 B.t10 B.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=7.215 pd=37.78 as=0 ps=0 w=18.5 l=3.53
X2 VDD1.t1 VP.t0 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=7.215 pd=37.78 as=7.215 ps=37.78 w=18.5 l=3.53
X3 VDD2.t1 VN.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=7.215 pd=37.78 as=7.215 ps=37.78 w=18.5 l=3.53
X4 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=7.215 pd=37.78 as=0 ps=0 w=18.5 l=3.53
X5 VDD2.t0 VN.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=7.215 pd=37.78 as=7.215 ps=37.78 w=18.5 l=3.53
X6 VDD1.t0 VP.t1 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=7.215 pd=37.78 as=7.215 ps=37.78 w=18.5 l=3.53
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=7.215 pd=37.78 as=0 ps=0 w=18.5 l=3.53
R0 B.n914 B.n913 585
R1 B.n915 B.n914 585
R2 B.n387 B.n125 585
R3 B.n386 B.n385 585
R4 B.n384 B.n383 585
R5 B.n382 B.n381 585
R6 B.n380 B.n379 585
R7 B.n378 B.n377 585
R8 B.n376 B.n375 585
R9 B.n374 B.n373 585
R10 B.n372 B.n371 585
R11 B.n370 B.n369 585
R12 B.n368 B.n367 585
R13 B.n366 B.n365 585
R14 B.n364 B.n363 585
R15 B.n362 B.n361 585
R16 B.n360 B.n359 585
R17 B.n358 B.n357 585
R18 B.n356 B.n355 585
R19 B.n354 B.n353 585
R20 B.n352 B.n351 585
R21 B.n350 B.n349 585
R22 B.n348 B.n347 585
R23 B.n346 B.n345 585
R24 B.n344 B.n343 585
R25 B.n342 B.n341 585
R26 B.n340 B.n339 585
R27 B.n338 B.n337 585
R28 B.n336 B.n335 585
R29 B.n334 B.n333 585
R30 B.n332 B.n331 585
R31 B.n330 B.n329 585
R32 B.n328 B.n327 585
R33 B.n326 B.n325 585
R34 B.n324 B.n323 585
R35 B.n322 B.n321 585
R36 B.n320 B.n319 585
R37 B.n318 B.n317 585
R38 B.n316 B.n315 585
R39 B.n314 B.n313 585
R40 B.n312 B.n311 585
R41 B.n310 B.n309 585
R42 B.n308 B.n307 585
R43 B.n306 B.n305 585
R44 B.n304 B.n303 585
R45 B.n302 B.n301 585
R46 B.n300 B.n299 585
R47 B.n298 B.n297 585
R48 B.n296 B.n295 585
R49 B.n294 B.n293 585
R50 B.n292 B.n291 585
R51 B.n290 B.n289 585
R52 B.n288 B.n287 585
R53 B.n286 B.n285 585
R54 B.n284 B.n283 585
R55 B.n282 B.n281 585
R56 B.n280 B.n279 585
R57 B.n278 B.n277 585
R58 B.n276 B.n275 585
R59 B.n274 B.n273 585
R60 B.n272 B.n271 585
R61 B.n270 B.n269 585
R62 B.n268 B.n267 585
R63 B.n266 B.n265 585
R64 B.n264 B.n263 585
R65 B.n262 B.n261 585
R66 B.n260 B.n259 585
R67 B.n258 B.n257 585
R68 B.n256 B.n255 585
R69 B.n254 B.n253 585
R70 B.n252 B.n251 585
R71 B.n249 B.n248 585
R72 B.n247 B.n246 585
R73 B.n245 B.n244 585
R74 B.n243 B.n242 585
R75 B.n241 B.n240 585
R76 B.n239 B.n238 585
R77 B.n237 B.n236 585
R78 B.n235 B.n234 585
R79 B.n233 B.n232 585
R80 B.n231 B.n230 585
R81 B.n229 B.n228 585
R82 B.n227 B.n226 585
R83 B.n225 B.n224 585
R84 B.n223 B.n222 585
R85 B.n221 B.n220 585
R86 B.n219 B.n218 585
R87 B.n217 B.n216 585
R88 B.n215 B.n214 585
R89 B.n213 B.n212 585
R90 B.n211 B.n210 585
R91 B.n209 B.n208 585
R92 B.n207 B.n206 585
R93 B.n205 B.n204 585
R94 B.n203 B.n202 585
R95 B.n201 B.n200 585
R96 B.n199 B.n198 585
R97 B.n197 B.n196 585
R98 B.n195 B.n194 585
R99 B.n193 B.n192 585
R100 B.n191 B.n190 585
R101 B.n189 B.n188 585
R102 B.n187 B.n186 585
R103 B.n185 B.n184 585
R104 B.n183 B.n182 585
R105 B.n181 B.n180 585
R106 B.n179 B.n178 585
R107 B.n177 B.n176 585
R108 B.n175 B.n174 585
R109 B.n173 B.n172 585
R110 B.n171 B.n170 585
R111 B.n169 B.n168 585
R112 B.n167 B.n166 585
R113 B.n165 B.n164 585
R114 B.n163 B.n162 585
R115 B.n161 B.n160 585
R116 B.n159 B.n158 585
R117 B.n157 B.n156 585
R118 B.n155 B.n154 585
R119 B.n153 B.n152 585
R120 B.n151 B.n150 585
R121 B.n149 B.n148 585
R122 B.n147 B.n146 585
R123 B.n145 B.n144 585
R124 B.n143 B.n142 585
R125 B.n141 B.n140 585
R126 B.n139 B.n138 585
R127 B.n137 B.n136 585
R128 B.n135 B.n134 585
R129 B.n133 B.n132 585
R130 B.n60 B.n59 585
R131 B.n918 B.n917 585
R132 B.n912 B.n126 585
R133 B.n126 B.n57 585
R134 B.n911 B.n56 585
R135 B.n922 B.n56 585
R136 B.n910 B.n55 585
R137 B.n923 B.n55 585
R138 B.n909 B.n54 585
R139 B.n924 B.n54 585
R140 B.n908 B.n907 585
R141 B.n907 B.n50 585
R142 B.n906 B.n49 585
R143 B.n930 B.n49 585
R144 B.n905 B.n48 585
R145 B.n931 B.n48 585
R146 B.n904 B.n47 585
R147 B.n932 B.n47 585
R148 B.n903 B.n902 585
R149 B.n902 B.n43 585
R150 B.n901 B.n42 585
R151 B.n938 B.n42 585
R152 B.n900 B.n41 585
R153 B.n939 B.n41 585
R154 B.n899 B.n40 585
R155 B.n940 B.n40 585
R156 B.n898 B.n897 585
R157 B.n897 B.n36 585
R158 B.n896 B.n35 585
R159 B.n946 B.n35 585
R160 B.n895 B.n34 585
R161 B.n947 B.n34 585
R162 B.n894 B.n33 585
R163 B.n948 B.n33 585
R164 B.n893 B.n892 585
R165 B.n892 B.n29 585
R166 B.n891 B.n28 585
R167 B.n954 B.n28 585
R168 B.n890 B.n27 585
R169 B.n955 B.n27 585
R170 B.n889 B.n26 585
R171 B.n956 B.n26 585
R172 B.n888 B.n887 585
R173 B.n887 B.n22 585
R174 B.n886 B.n21 585
R175 B.n962 B.n21 585
R176 B.n885 B.n20 585
R177 B.n963 B.n20 585
R178 B.n884 B.n19 585
R179 B.n964 B.n19 585
R180 B.n883 B.n882 585
R181 B.n882 B.n15 585
R182 B.n881 B.n14 585
R183 B.n970 B.n14 585
R184 B.n880 B.n13 585
R185 B.n971 B.n13 585
R186 B.n879 B.n12 585
R187 B.n972 B.n12 585
R188 B.n878 B.n877 585
R189 B.n877 B.n8 585
R190 B.n876 B.n7 585
R191 B.n978 B.n7 585
R192 B.n875 B.n6 585
R193 B.n979 B.n6 585
R194 B.n874 B.n5 585
R195 B.n980 B.n5 585
R196 B.n873 B.n872 585
R197 B.n872 B.n4 585
R198 B.n871 B.n388 585
R199 B.n871 B.n870 585
R200 B.n861 B.n389 585
R201 B.n390 B.n389 585
R202 B.n863 B.n862 585
R203 B.n864 B.n863 585
R204 B.n860 B.n395 585
R205 B.n395 B.n394 585
R206 B.n859 B.n858 585
R207 B.n858 B.n857 585
R208 B.n397 B.n396 585
R209 B.n398 B.n397 585
R210 B.n850 B.n849 585
R211 B.n851 B.n850 585
R212 B.n848 B.n403 585
R213 B.n403 B.n402 585
R214 B.n847 B.n846 585
R215 B.n846 B.n845 585
R216 B.n405 B.n404 585
R217 B.n406 B.n405 585
R218 B.n838 B.n837 585
R219 B.n839 B.n838 585
R220 B.n836 B.n411 585
R221 B.n411 B.n410 585
R222 B.n835 B.n834 585
R223 B.n834 B.n833 585
R224 B.n413 B.n412 585
R225 B.n414 B.n413 585
R226 B.n826 B.n825 585
R227 B.n827 B.n826 585
R228 B.n824 B.n419 585
R229 B.n419 B.n418 585
R230 B.n823 B.n822 585
R231 B.n822 B.n821 585
R232 B.n421 B.n420 585
R233 B.n422 B.n421 585
R234 B.n814 B.n813 585
R235 B.n815 B.n814 585
R236 B.n812 B.n427 585
R237 B.n427 B.n426 585
R238 B.n811 B.n810 585
R239 B.n810 B.n809 585
R240 B.n429 B.n428 585
R241 B.n430 B.n429 585
R242 B.n802 B.n801 585
R243 B.n803 B.n802 585
R244 B.n800 B.n435 585
R245 B.n435 B.n434 585
R246 B.n799 B.n798 585
R247 B.n798 B.n797 585
R248 B.n437 B.n436 585
R249 B.n438 B.n437 585
R250 B.n790 B.n789 585
R251 B.n791 B.n790 585
R252 B.n788 B.n443 585
R253 B.n443 B.n442 585
R254 B.n787 B.n786 585
R255 B.n786 B.n785 585
R256 B.n445 B.n444 585
R257 B.n446 B.n445 585
R258 B.n781 B.n780 585
R259 B.n449 B.n448 585
R260 B.n777 B.n776 585
R261 B.n778 B.n777 585
R262 B.n775 B.n514 585
R263 B.n774 B.n773 585
R264 B.n772 B.n771 585
R265 B.n770 B.n769 585
R266 B.n768 B.n767 585
R267 B.n766 B.n765 585
R268 B.n764 B.n763 585
R269 B.n762 B.n761 585
R270 B.n760 B.n759 585
R271 B.n758 B.n757 585
R272 B.n756 B.n755 585
R273 B.n754 B.n753 585
R274 B.n752 B.n751 585
R275 B.n750 B.n749 585
R276 B.n748 B.n747 585
R277 B.n746 B.n745 585
R278 B.n744 B.n743 585
R279 B.n742 B.n741 585
R280 B.n740 B.n739 585
R281 B.n738 B.n737 585
R282 B.n736 B.n735 585
R283 B.n734 B.n733 585
R284 B.n732 B.n731 585
R285 B.n730 B.n729 585
R286 B.n728 B.n727 585
R287 B.n726 B.n725 585
R288 B.n724 B.n723 585
R289 B.n722 B.n721 585
R290 B.n720 B.n719 585
R291 B.n718 B.n717 585
R292 B.n716 B.n715 585
R293 B.n714 B.n713 585
R294 B.n712 B.n711 585
R295 B.n710 B.n709 585
R296 B.n708 B.n707 585
R297 B.n706 B.n705 585
R298 B.n704 B.n703 585
R299 B.n702 B.n701 585
R300 B.n700 B.n699 585
R301 B.n698 B.n697 585
R302 B.n696 B.n695 585
R303 B.n694 B.n693 585
R304 B.n692 B.n691 585
R305 B.n690 B.n689 585
R306 B.n688 B.n687 585
R307 B.n686 B.n685 585
R308 B.n684 B.n683 585
R309 B.n682 B.n681 585
R310 B.n680 B.n679 585
R311 B.n678 B.n677 585
R312 B.n676 B.n675 585
R313 B.n674 B.n673 585
R314 B.n672 B.n671 585
R315 B.n670 B.n669 585
R316 B.n668 B.n667 585
R317 B.n666 B.n665 585
R318 B.n664 B.n663 585
R319 B.n662 B.n661 585
R320 B.n660 B.n659 585
R321 B.n658 B.n657 585
R322 B.n656 B.n655 585
R323 B.n654 B.n653 585
R324 B.n652 B.n651 585
R325 B.n650 B.n649 585
R326 B.n648 B.n647 585
R327 B.n646 B.n645 585
R328 B.n644 B.n643 585
R329 B.n641 B.n640 585
R330 B.n639 B.n638 585
R331 B.n637 B.n636 585
R332 B.n635 B.n634 585
R333 B.n633 B.n632 585
R334 B.n631 B.n630 585
R335 B.n629 B.n628 585
R336 B.n627 B.n626 585
R337 B.n625 B.n624 585
R338 B.n623 B.n622 585
R339 B.n621 B.n620 585
R340 B.n619 B.n618 585
R341 B.n617 B.n616 585
R342 B.n615 B.n614 585
R343 B.n613 B.n612 585
R344 B.n611 B.n610 585
R345 B.n609 B.n608 585
R346 B.n607 B.n606 585
R347 B.n605 B.n604 585
R348 B.n603 B.n602 585
R349 B.n601 B.n600 585
R350 B.n599 B.n598 585
R351 B.n597 B.n596 585
R352 B.n595 B.n594 585
R353 B.n593 B.n592 585
R354 B.n591 B.n590 585
R355 B.n589 B.n588 585
R356 B.n587 B.n586 585
R357 B.n585 B.n584 585
R358 B.n583 B.n582 585
R359 B.n581 B.n580 585
R360 B.n579 B.n578 585
R361 B.n577 B.n576 585
R362 B.n575 B.n574 585
R363 B.n573 B.n572 585
R364 B.n571 B.n570 585
R365 B.n569 B.n568 585
R366 B.n567 B.n566 585
R367 B.n565 B.n564 585
R368 B.n563 B.n562 585
R369 B.n561 B.n560 585
R370 B.n559 B.n558 585
R371 B.n557 B.n556 585
R372 B.n555 B.n554 585
R373 B.n553 B.n552 585
R374 B.n551 B.n550 585
R375 B.n549 B.n548 585
R376 B.n547 B.n546 585
R377 B.n545 B.n544 585
R378 B.n543 B.n542 585
R379 B.n541 B.n540 585
R380 B.n539 B.n538 585
R381 B.n537 B.n536 585
R382 B.n535 B.n534 585
R383 B.n533 B.n532 585
R384 B.n531 B.n530 585
R385 B.n529 B.n528 585
R386 B.n527 B.n526 585
R387 B.n525 B.n524 585
R388 B.n523 B.n522 585
R389 B.n521 B.n520 585
R390 B.n782 B.n447 585
R391 B.n447 B.n446 585
R392 B.n784 B.n783 585
R393 B.n785 B.n784 585
R394 B.n441 B.n440 585
R395 B.n442 B.n441 585
R396 B.n793 B.n792 585
R397 B.n792 B.n791 585
R398 B.n794 B.n439 585
R399 B.n439 B.n438 585
R400 B.n796 B.n795 585
R401 B.n797 B.n796 585
R402 B.n433 B.n432 585
R403 B.n434 B.n433 585
R404 B.n805 B.n804 585
R405 B.n804 B.n803 585
R406 B.n806 B.n431 585
R407 B.n431 B.n430 585
R408 B.n808 B.n807 585
R409 B.n809 B.n808 585
R410 B.n425 B.n424 585
R411 B.n426 B.n425 585
R412 B.n817 B.n816 585
R413 B.n816 B.n815 585
R414 B.n818 B.n423 585
R415 B.n423 B.n422 585
R416 B.n820 B.n819 585
R417 B.n821 B.n820 585
R418 B.n417 B.n416 585
R419 B.n418 B.n417 585
R420 B.n829 B.n828 585
R421 B.n828 B.n827 585
R422 B.n830 B.n415 585
R423 B.n415 B.n414 585
R424 B.n832 B.n831 585
R425 B.n833 B.n832 585
R426 B.n409 B.n408 585
R427 B.n410 B.n409 585
R428 B.n841 B.n840 585
R429 B.n840 B.n839 585
R430 B.n842 B.n407 585
R431 B.n407 B.n406 585
R432 B.n844 B.n843 585
R433 B.n845 B.n844 585
R434 B.n401 B.n400 585
R435 B.n402 B.n401 585
R436 B.n853 B.n852 585
R437 B.n852 B.n851 585
R438 B.n854 B.n399 585
R439 B.n399 B.n398 585
R440 B.n856 B.n855 585
R441 B.n857 B.n856 585
R442 B.n393 B.n392 585
R443 B.n394 B.n393 585
R444 B.n866 B.n865 585
R445 B.n865 B.n864 585
R446 B.n867 B.n391 585
R447 B.n391 B.n390 585
R448 B.n869 B.n868 585
R449 B.n870 B.n869 585
R450 B.n2 B.n0 585
R451 B.n4 B.n2 585
R452 B.n3 B.n1 585
R453 B.n979 B.n3 585
R454 B.n977 B.n976 585
R455 B.n978 B.n977 585
R456 B.n975 B.n9 585
R457 B.n9 B.n8 585
R458 B.n974 B.n973 585
R459 B.n973 B.n972 585
R460 B.n11 B.n10 585
R461 B.n971 B.n11 585
R462 B.n969 B.n968 585
R463 B.n970 B.n969 585
R464 B.n967 B.n16 585
R465 B.n16 B.n15 585
R466 B.n966 B.n965 585
R467 B.n965 B.n964 585
R468 B.n18 B.n17 585
R469 B.n963 B.n18 585
R470 B.n961 B.n960 585
R471 B.n962 B.n961 585
R472 B.n959 B.n23 585
R473 B.n23 B.n22 585
R474 B.n958 B.n957 585
R475 B.n957 B.n956 585
R476 B.n25 B.n24 585
R477 B.n955 B.n25 585
R478 B.n953 B.n952 585
R479 B.n954 B.n953 585
R480 B.n951 B.n30 585
R481 B.n30 B.n29 585
R482 B.n950 B.n949 585
R483 B.n949 B.n948 585
R484 B.n32 B.n31 585
R485 B.n947 B.n32 585
R486 B.n945 B.n944 585
R487 B.n946 B.n945 585
R488 B.n943 B.n37 585
R489 B.n37 B.n36 585
R490 B.n942 B.n941 585
R491 B.n941 B.n940 585
R492 B.n39 B.n38 585
R493 B.n939 B.n39 585
R494 B.n937 B.n936 585
R495 B.n938 B.n937 585
R496 B.n935 B.n44 585
R497 B.n44 B.n43 585
R498 B.n934 B.n933 585
R499 B.n933 B.n932 585
R500 B.n46 B.n45 585
R501 B.n931 B.n46 585
R502 B.n929 B.n928 585
R503 B.n930 B.n929 585
R504 B.n927 B.n51 585
R505 B.n51 B.n50 585
R506 B.n926 B.n925 585
R507 B.n925 B.n924 585
R508 B.n53 B.n52 585
R509 B.n923 B.n53 585
R510 B.n921 B.n920 585
R511 B.n922 B.n921 585
R512 B.n919 B.n58 585
R513 B.n58 B.n57 585
R514 B.n982 B.n981 585
R515 B.n981 B.n980 585
R516 B.n780 B.n447 473.281
R517 B.n917 B.n58 473.281
R518 B.n520 B.n445 473.281
R519 B.n914 B.n126 473.281
R520 B.n518 B.t10 335.423
R521 B.n515 B.t2 335.423
R522 B.n130 B.t6 335.423
R523 B.n127 B.t13 335.423
R524 B.n915 B.n124 256.663
R525 B.n915 B.n123 256.663
R526 B.n915 B.n122 256.663
R527 B.n915 B.n121 256.663
R528 B.n915 B.n120 256.663
R529 B.n915 B.n119 256.663
R530 B.n915 B.n118 256.663
R531 B.n915 B.n117 256.663
R532 B.n915 B.n116 256.663
R533 B.n915 B.n115 256.663
R534 B.n915 B.n114 256.663
R535 B.n915 B.n113 256.663
R536 B.n915 B.n112 256.663
R537 B.n915 B.n111 256.663
R538 B.n915 B.n110 256.663
R539 B.n915 B.n109 256.663
R540 B.n915 B.n108 256.663
R541 B.n915 B.n107 256.663
R542 B.n915 B.n106 256.663
R543 B.n915 B.n105 256.663
R544 B.n915 B.n104 256.663
R545 B.n915 B.n103 256.663
R546 B.n915 B.n102 256.663
R547 B.n915 B.n101 256.663
R548 B.n915 B.n100 256.663
R549 B.n915 B.n99 256.663
R550 B.n915 B.n98 256.663
R551 B.n915 B.n97 256.663
R552 B.n915 B.n96 256.663
R553 B.n915 B.n95 256.663
R554 B.n915 B.n94 256.663
R555 B.n915 B.n93 256.663
R556 B.n915 B.n92 256.663
R557 B.n915 B.n91 256.663
R558 B.n915 B.n90 256.663
R559 B.n915 B.n89 256.663
R560 B.n915 B.n88 256.663
R561 B.n915 B.n87 256.663
R562 B.n915 B.n86 256.663
R563 B.n915 B.n85 256.663
R564 B.n915 B.n84 256.663
R565 B.n915 B.n83 256.663
R566 B.n915 B.n82 256.663
R567 B.n915 B.n81 256.663
R568 B.n915 B.n80 256.663
R569 B.n915 B.n79 256.663
R570 B.n915 B.n78 256.663
R571 B.n915 B.n77 256.663
R572 B.n915 B.n76 256.663
R573 B.n915 B.n75 256.663
R574 B.n915 B.n74 256.663
R575 B.n915 B.n73 256.663
R576 B.n915 B.n72 256.663
R577 B.n915 B.n71 256.663
R578 B.n915 B.n70 256.663
R579 B.n915 B.n69 256.663
R580 B.n915 B.n68 256.663
R581 B.n915 B.n67 256.663
R582 B.n915 B.n66 256.663
R583 B.n915 B.n65 256.663
R584 B.n915 B.n64 256.663
R585 B.n915 B.n63 256.663
R586 B.n915 B.n62 256.663
R587 B.n915 B.n61 256.663
R588 B.n916 B.n915 256.663
R589 B.n779 B.n778 256.663
R590 B.n778 B.n450 256.663
R591 B.n778 B.n451 256.663
R592 B.n778 B.n452 256.663
R593 B.n778 B.n453 256.663
R594 B.n778 B.n454 256.663
R595 B.n778 B.n455 256.663
R596 B.n778 B.n456 256.663
R597 B.n778 B.n457 256.663
R598 B.n778 B.n458 256.663
R599 B.n778 B.n459 256.663
R600 B.n778 B.n460 256.663
R601 B.n778 B.n461 256.663
R602 B.n778 B.n462 256.663
R603 B.n778 B.n463 256.663
R604 B.n778 B.n464 256.663
R605 B.n778 B.n465 256.663
R606 B.n778 B.n466 256.663
R607 B.n778 B.n467 256.663
R608 B.n778 B.n468 256.663
R609 B.n778 B.n469 256.663
R610 B.n778 B.n470 256.663
R611 B.n778 B.n471 256.663
R612 B.n778 B.n472 256.663
R613 B.n778 B.n473 256.663
R614 B.n778 B.n474 256.663
R615 B.n778 B.n475 256.663
R616 B.n778 B.n476 256.663
R617 B.n778 B.n477 256.663
R618 B.n778 B.n478 256.663
R619 B.n778 B.n479 256.663
R620 B.n778 B.n480 256.663
R621 B.n778 B.n481 256.663
R622 B.n778 B.n482 256.663
R623 B.n778 B.n483 256.663
R624 B.n778 B.n484 256.663
R625 B.n778 B.n485 256.663
R626 B.n778 B.n486 256.663
R627 B.n778 B.n487 256.663
R628 B.n778 B.n488 256.663
R629 B.n778 B.n489 256.663
R630 B.n778 B.n490 256.663
R631 B.n778 B.n491 256.663
R632 B.n778 B.n492 256.663
R633 B.n778 B.n493 256.663
R634 B.n778 B.n494 256.663
R635 B.n778 B.n495 256.663
R636 B.n778 B.n496 256.663
R637 B.n778 B.n497 256.663
R638 B.n778 B.n498 256.663
R639 B.n778 B.n499 256.663
R640 B.n778 B.n500 256.663
R641 B.n778 B.n501 256.663
R642 B.n778 B.n502 256.663
R643 B.n778 B.n503 256.663
R644 B.n778 B.n504 256.663
R645 B.n778 B.n505 256.663
R646 B.n778 B.n506 256.663
R647 B.n778 B.n507 256.663
R648 B.n778 B.n508 256.663
R649 B.n778 B.n509 256.663
R650 B.n778 B.n510 256.663
R651 B.n778 B.n511 256.663
R652 B.n778 B.n512 256.663
R653 B.n778 B.n513 256.663
R654 B.n784 B.n447 163.367
R655 B.n784 B.n441 163.367
R656 B.n792 B.n441 163.367
R657 B.n792 B.n439 163.367
R658 B.n796 B.n439 163.367
R659 B.n796 B.n433 163.367
R660 B.n804 B.n433 163.367
R661 B.n804 B.n431 163.367
R662 B.n808 B.n431 163.367
R663 B.n808 B.n425 163.367
R664 B.n816 B.n425 163.367
R665 B.n816 B.n423 163.367
R666 B.n820 B.n423 163.367
R667 B.n820 B.n417 163.367
R668 B.n828 B.n417 163.367
R669 B.n828 B.n415 163.367
R670 B.n832 B.n415 163.367
R671 B.n832 B.n409 163.367
R672 B.n840 B.n409 163.367
R673 B.n840 B.n407 163.367
R674 B.n844 B.n407 163.367
R675 B.n844 B.n401 163.367
R676 B.n852 B.n401 163.367
R677 B.n852 B.n399 163.367
R678 B.n856 B.n399 163.367
R679 B.n856 B.n393 163.367
R680 B.n865 B.n393 163.367
R681 B.n865 B.n391 163.367
R682 B.n869 B.n391 163.367
R683 B.n869 B.n2 163.367
R684 B.n981 B.n2 163.367
R685 B.n981 B.n3 163.367
R686 B.n977 B.n3 163.367
R687 B.n977 B.n9 163.367
R688 B.n973 B.n9 163.367
R689 B.n973 B.n11 163.367
R690 B.n969 B.n11 163.367
R691 B.n969 B.n16 163.367
R692 B.n965 B.n16 163.367
R693 B.n965 B.n18 163.367
R694 B.n961 B.n18 163.367
R695 B.n961 B.n23 163.367
R696 B.n957 B.n23 163.367
R697 B.n957 B.n25 163.367
R698 B.n953 B.n25 163.367
R699 B.n953 B.n30 163.367
R700 B.n949 B.n30 163.367
R701 B.n949 B.n32 163.367
R702 B.n945 B.n32 163.367
R703 B.n945 B.n37 163.367
R704 B.n941 B.n37 163.367
R705 B.n941 B.n39 163.367
R706 B.n937 B.n39 163.367
R707 B.n937 B.n44 163.367
R708 B.n933 B.n44 163.367
R709 B.n933 B.n46 163.367
R710 B.n929 B.n46 163.367
R711 B.n929 B.n51 163.367
R712 B.n925 B.n51 163.367
R713 B.n925 B.n53 163.367
R714 B.n921 B.n53 163.367
R715 B.n921 B.n58 163.367
R716 B.n777 B.n449 163.367
R717 B.n777 B.n514 163.367
R718 B.n773 B.n772 163.367
R719 B.n769 B.n768 163.367
R720 B.n765 B.n764 163.367
R721 B.n761 B.n760 163.367
R722 B.n757 B.n756 163.367
R723 B.n753 B.n752 163.367
R724 B.n749 B.n748 163.367
R725 B.n745 B.n744 163.367
R726 B.n741 B.n740 163.367
R727 B.n737 B.n736 163.367
R728 B.n733 B.n732 163.367
R729 B.n729 B.n728 163.367
R730 B.n725 B.n724 163.367
R731 B.n721 B.n720 163.367
R732 B.n717 B.n716 163.367
R733 B.n713 B.n712 163.367
R734 B.n709 B.n708 163.367
R735 B.n705 B.n704 163.367
R736 B.n701 B.n700 163.367
R737 B.n697 B.n696 163.367
R738 B.n693 B.n692 163.367
R739 B.n689 B.n688 163.367
R740 B.n685 B.n684 163.367
R741 B.n681 B.n680 163.367
R742 B.n677 B.n676 163.367
R743 B.n673 B.n672 163.367
R744 B.n669 B.n668 163.367
R745 B.n665 B.n664 163.367
R746 B.n661 B.n660 163.367
R747 B.n657 B.n656 163.367
R748 B.n653 B.n652 163.367
R749 B.n649 B.n648 163.367
R750 B.n645 B.n644 163.367
R751 B.n640 B.n639 163.367
R752 B.n636 B.n635 163.367
R753 B.n632 B.n631 163.367
R754 B.n628 B.n627 163.367
R755 B.n624 B.n623 163.367
R756 B.n620 B.n619 163.367
R757 B.n616 B.n615 163.367
R758 B.n612 B.n611 163.367
R759 B.n608 B.n607 163.367
R760 B.n604 B.n603 163.367
R761 B.n600 B.n599 163.367
R762 B.n596 B.n595 163.367
R763 B.n592 B.n591 163.367
R764 B.n588 B.n587 163.367
R765 B.n584 B.n583 163.367
R766 B.n580 B.n579 163.367
R767 B.n576 B.n575 163.367
R768 B.n572 B.n571 163.367
R769 B.n568 B.n567 163.367
R770 B.n564 B.n563 163.367
R771 B.n560 B.n559 163.367
R772 B.n556 B.n555 163.367
R773 B.n552 B.n551 163.367
R774 B.n548 B.n547 163.367
R775 B.n544 B.n543 163.367
R776 B.n540 B.n539 163.367
R777 B.n536 B.n535 163.367
R778 B.n532 B.n531 163.367
R779 B.n528 B.n527 163.367
R780 B.n524 B.n523 163.367
R781 B.n786 B.n445 163.367
R782 B.n786 B.n443 163.367
R783 B.n790 B.n443 163.367
R784 B.n790 B.n437 163.367
R785 B.n798 B.n437 163.367
R786 B.n798 B.n435 163.367
R787 B.n802 B.n435 163.367
R788 B.n802 B.n429 163.367
R789 B.n810 B.n429 163.367
R790 B.n810 B.n427 163.367
R791 B.n814 B.n427 163.367
R792 B.n814 B.n421 163.367
R793 B.n822 B.n421 163.367
R794 B.n822 B.n419 163.367
R795 B.n826 B.n419 163.367
R796 B.n826 B.n413 163.367
R797 B.n834 B.n413 163.367
R798 B.n834 B.n411 163.367
R799 B.n838 B.n411 163.367
R800 B.n838 B.n405 163.367
R801 B.n846 B.n405 163.367
R802 B.n846 B.n403 163.367
R803 B.n850 B.n403 163.367
R804 B.n850 B.n397 163.367
R805 B.n858 B.n397 163.367
R806 B.n858 B.n395 163.367
R807 B.n863 B.n395 163.367
R808 B.n863 B.n389 163.367
R809 B.n871 B.n389 163.367
R810 B.n872 B.n871 163.367
R811 B.n872 B.n5 163.367
R812 B.n6 B.n5 163.367
R813 B.n7 B.n6 163.367
R814 B.n877 B.n7 163.367
R815 B.n877 B.n12 163.367
R816 B.n13 B.n12 163.367
R817 B.n14 B.n13 163.367
R818 B.n882 B.n14 163.367
R819 B.n882 B.n19 163.367
R820 B.n20 B.n19 163.367
R821 B.n21 B.n20 163.367
R822 B.n887 B.n21 163.367
R823 B.n887 B.n26 163.367
R824 B.n27 B.n26 163.367
R825 B.n28 B.n27 163.367
R826 B.n892 B.n28 163.367
R827 B.n892 B.n33 163.367
R828 B.n34 B.n33 163.367
R829 B.n35 B.n34 163.367
R830 B.n897 B.n35 163.367
R831 B.n897 B.n40 163.367
R832 B.n41 B.n40 163.367
R833 B.n42 B.n41 163.367
R834 B.n902 B.n42 163.367
R835 B.n902 B.n47 163.367
R836 B.n48 B.n47 163.367
R837 B.n49 B.n48 163.367
R838 B.n907 B.n49 163.367
R839 B.n907 B.n54 163.367
R840 B.n55 B.n54 163.367
R841 B.n56 B.n55 163.367
R842 B.n126 B.n56 163.367
R843 B.n132 B.n60 163.367
R844 B.n136 B.n135 163.367
R845 B.n140 B.n139 163.367
R846 B.n144 B.n143 163.367
R847 B.n148 B.n147 163.367
R848 B.n152 B.n151 163.367
R849 B.n156 B.n155 163.367
R850 B.n160 B.n159 163.367
R851 B.n164 B.n163 163.367
R852 B.n168 B.n167 163.367
R853 B.n172 B.n171 163.367
R854 B.n176 B.n175 163.367
R855 B.n180 B.n179 163.367
R856 B.n184 B.n183 163.367
R857 B.n188 B.n187 163.367
R858 B.n192 B.n191 163.367
R859 B.n196 B.n195 163.367
R860 B.n200 B.n199 163.367
R861 B.n204 B.n203 163.367
R862 B.n208 B.n207 163.367
R863 B.n212 B.n211 163.367
R864 B.n216 B.n215 163.367
R865 B.n220 B.n219 163.367
R866 B.n224 B.n223 163.367
R867 B.n228 B.n227 163.367
R868 B.n232 B.n231 163.367
R869 B.n236 B.n235 163.367
R870 B.n240 B.n239 163.367
R871 B.n244 B.n243 163.367
R872 B.n248 B.n247 163.367
R873 B.n253 B.n252 163.367
R874 B.n257 B.n256 163.367
R875 B.n261 B.n260 163.367
R876 B.n265 B.n264 163.367
R877 B.n269 B.n268 163.367
R878 B.n273 B.n272 163.367
R879 B.n277 B.n276 163.367
R880 B.n281 B.n280 163.367
R881 B.n285 B.n284 163.367
R882 B.n289 B.n288 163.367
R883 B.n293 B.n292 163.367
R884 B.n297 B.n296 163.367
R885 B.n301 B.n300 163.367
R886 B.n305 B.n304 163.367
R887 B.n309 B.n308 163.367
R888 B.n313 B.n312 163.367
R889 B.n317 B.n316 163.367
R890 B.n321 B.n320 163.367
R891 B.n325 B.n324 163.367
R892 B.n329 B.n328 163.367
R893 B.n333 B.n332 163.367
R894 B.n337 B.n336 163.367
R895 B.n341 B.n340 163.367
R896 B.n345 B.n344 163.367
R897 B.n349 B.n348 163.367
R898 B.n353 B.n352 163.367
R899 B.n357 B.n356 163.367
R900 B.n361 B.n360 163.367
R901 B.n365 B.n364 163.367
R902 B.n369 B.n368 163.367
R903 B.n373 B.n372 163.367
R904 B.n377 B.n376 163.367
R905 B.n381 B.n380 163.367
R906 B.n385 B.n384 163.367
R907 B.n914 B.n125 163.367
R908 B.n518 B.t12 144.796
R909 B.n127 B.t14 144.796
R910 B.n515 B.t5 144.77
R911 B.n130 B.t8 144.77
R912 B.n519 B.n518 74.8611
R913 B.n516 B.n515 74.8611
R914 B.n131 B.n130 74.8611
R915 B.n128 B.n127 74.8611
R916 B.n780 B.n779 71.676
R917 B.n514 B.n450 71.676
R918 B.n772 B.n451 71.676
R919 B.n768 B.n452 71.676
R920 B.n764 B.n453 71.676
R921 B.n760 B.n454 71.676
R922 B.n756 B.n455 71.676
R923 B.n752 B.n456 71.676
R924 B.n748 B.n457 71.676
R925 B.n744 B.n458 71.676
R926 B.n740 B.n459 71.676
R927 B.n736 B.n460 71.676
R928 B.n732 B.n461 71.676
R929 B.n728 B.n462 71.676
R930 B.n724 B.n463 71.676
R931 B.n720 B.n464 71.676
R932 B.n716 B.n465 71.676
R933 B.n712 B.n466 71.676
R934 B.n708 B.n467 71.676
R935 B.n704 B.n468 71.676
R936 B.n700 B.n469 71.676
R937 B.n696 B.n470 71.676
R938 B.n692 B.n471 71.676
R939 B.n688 B.n472 71.676
R940 B.n684 B.n473 71.676
R941 B.n680 B.n474 71.676
R942 B.n676 B.n475 71.676
R943 B.n672 B.n476 71.676
R944 B.n668 B.n477 71.676
R945 B.n664 B.n478 71.676
R946 B.n660 B.n479 71.676
R947 B.n656 B.n480 71.676
R948 B.n652 B.n481 71.676
R949 B.n648 B.n482 71.676
R950 B.n644 B.n483 71.676
R951 B.n639 B.n484 71.676
R952 B.n635 B.n485 71.676
R953 B.n631 B.n486 71.676
R954 B.n627 B.n487 71.676
R955 B.n623 B.n488 71.676
R956 B.n619 B.n489 71.676
R957 B.n615 B.n490 71.676
R958 B.n611 B.n491 71.676
R959 B.n607 B.n492 71.676
R960 B.n603 B.n493 71.676
R961 B.n599 B.n494 71.676
R962 B.n595 B.n495 71.676
R963 B.n591 B.n496 71.676
R964 B.n587 B.n497 71.676
R965 B.n583 B.n498 71.676
R966 B.n579 B.n499 71.676
R967 B.n575 B.n500 71.676
R968 B.n571 B.n501 71.676
R969 B.n567 B.n502 71.676
R970 B.n563 B.n503 71.676
R971 B.n559 B.n504 71.676
R972 B.n555 B.n505 71.676
R973 B.n551 B.n506 71.676
R974 B.n547 B.n507 71.676
R975 B.n543 B.n508 71.676
R976 B.n539 B.n509 71.676
R977 B.n535 B.n510 71.676
R978 B.n531 B.n511 71.676
R979 B.n527 B.n512 71.676
R980 B.n523 B.n513 71.676
R981 B.n917 B.n916 71.676
R982 B.n132 B.n61 71.676
R983 B.n136 B.n62 71.676
R984 B.n140 B.n63 71.676
R985 B.n144 B.n64 71.676
R986 B.n148 B.n65 71.676
R987 B.n152 B.n66 71.676
R988 B.n156 B.n67 71.676
R989 B.n160 B.n68 71.676
R990 B.n164 B.n69 71.676
R991 B.n168 B.n70 71.676
R992 B.n172 B.n71 71.676
R993 B.n176 B.n72 71.676
R994 B.n180 B.n73 71.676
R995 B.n184 B.n74 71.676
R996 B.n188 B.n75 71.676
R997 B.n192 B.n76 71.676
R998 B.n196 B.n77 71.676
R999 B.n200 B.n78 71.676
R1000 B.n204 B.n79 71.676
R1001 B.n208 B.n80 71.676
R1002 B.n212 B.n81 71.676
R1003 B.n216 B.n82 71.676
R1004 B.n220 B.n83 71.676
R1005 B.n224 B.n84 71.676
R1006 B.n228 B.n85 71.676
R1007 B.n232 B.n86 71.676
R1008 B.n236 B.n87 71.676
R1009 B.n240 B.n88 71.676
R1010 B.n244 B.n89 71.676
R1011 B.n248 B.n90 71.676
R1012 B.n253 B.n91 71.676
R1013 B.n257 B.n92 71.676
R1014 B.n261 B.n93 71.676
R1015 B.n265 B.n94 71.676
R1016 B.n269 B.n95 71.676
R1017 B.n273 B.n96 71.676
R1018 B.n277 B.n97 71.676
R1019 B.n281 B.n98 71.676
R1020 B.n285 B.n99 71.676
R1021 B.n289 B.n100 71.676
R1022 B.n293 B.n101 71.676
R1023 B.n297 B.n102 71.676
R1024 B.n301 B.n103 71.676
R1025 B.n305 B.n104 71.676
R1026 B.n309 B.n105 71.676
R1027 B.n313 B.n106 71.676
R1028 B.n317 B.n107 71.676
R1029 B.n321 B.n108 71.676
R1030 B.n325 B.n109 71.676
R1031 B.n329 B.n110 71.676
R1032 B.n333 B.n111 71.676
R1033 B.n337 B.n112 71.676
R1034 B.n341 B.n113 71.676
R1035 B.n345 B.n114 71.676
R1036 B.n349 B.n115 71.676
R1037 B.n353 B.n116 71.676
R1038 B.n357 B.n117 71.676
R1039 B.n361 B.n118 71.676
R1040 B.n365 B.n119 71.676
R1041 B.n369 B.n120 71.676
R1042 B.n373 B.n121 71.676
R1043 B.n377 B.n122 71.676
R1044 B.n381 B.n123 71.676
R1045 B.n385 B.n124 71.676
R1046 B.n125 B.n124 71.676
R1047 B.n384 B.n123 71.676
R1048 B.n380 B.n122 71.676
R1049 B.n376 B.n121 71.676
R1050 B.n372 B.n120 71.676
R1051 B.n368 B.n119 71.676
R1052 B.n364 B.n118 71.676
R1053 B.n360 B.n117 71.676
R1054 B.n356 B.n116 71.676
R1055 B.n352 B.n115 71.676
R1056 B.n348 B.n114 71.676
R1057 B.n344 B.n113 71.676
R1058 B.n340 B.n112 71.676
R1059 B.n336 B.n111 71.676
R1060 B.n332 B.n110 71.676
R1061 B.n328 B.n109 71.676
R1062 B.n324 B.n108 71.676
R1063 B.n320 B.n107 71.676
R1064 B.n316 B.n106 71.676
R1065 B.n312 B.n105 71.676
R1066 B.n308 B.n104 71.676
R1067 B.n304 B.n103 71.676
R1068 B.n300 B.n102 71.676
R1069 B.n296 B.n101 71.676
R1070 B.n292 B.n100 71.676
R1071 B.n288 B.n99 71.676
R1072 B.n284 B.n98 71.676
R1073 B.n280 B.n97 71.676
R1074 B.n276 B.n96 71.676
R1075 B.n272 B.n95 71.676
R1076 B.n268 B.n94 71.676
R1077 B.n264 B.n93 71.676
R1078 B.n260 B.n92 71.676
R1079 B.n256 B.n91 71.676
R1080 B.n252 B.n90 71.676
R1081 B.n247 B.n89 71.676
R1082 B.n243 B.n88 71.676
R1083 B.n239 B.n87 71.676
R1084 B.n235 B.n86 71.676
R1085 B.n231 B.n85 71.676
R1086 B.n227 B.n84 71.676
R1087 B.n223 B.n83 71.676
R1088 B.n219 B.n82 71.676
R1089 B.n215 B.n81 71.676
R1090 B.n211 B.n80 71.676
R1091 B.n207 B.n79 71.676
R1092 B.n203 B.n78 71.676
R1093 B.n199 B.n77 71.676
R1094 B.n195 B.n76 71.676
R1095 B.n191 B.n75 71.676
R1096 B.n187 B.n74 71.676
R1097 B.n183 B.n73 71.676
R1098 B.n179 B.n72 71.676
R1099 B.n175 B.n71 71.676
R1100 B.n171 B.n70 71.676
R1101 B.n167 B.n69 71.676
R1102 B.n163 B.n68 71.676
R1103 B.n159 B.n67 71.676
R1104 B.n155 B.n66 71.676
R1105 B.n151 B.n65 71.676
R1106 B.n147 B.n64 71.676
R1107 B.n143 B.n63 71.676
R1108 B.n139 B.n62 71.676
R1109 B.n135 B.n61 71.676
R1110 B.n916 B.n60 71.676
R1111 B.n779 B.n449 71.676
R1112 B.n773 B.n450 71.676
R1113 B.n769 B.n451 71.676
R1114 B.n765 B.n452 71.676
R1115 B.n761 B.n453 71.676
R1116 B.n757 B.n454 71.676
R1117 B.n753 B.n455 71.676
R1118 B.n749 B.n456 71.676
R1119 B.n745 B.n457 71.676
R1120 B.n741 B.n458 71.676
R1121 B.n737 B.n459 71.676
R1122 B.n733 B.n460 71.676
R1123 B.n729 B.n461 71.676
R1124 B.n725 B.n462 71.676
R1125 B.n721 B.n463 71.676
R1126 B.n717 B.n464 71.676
R1127 B.n713 B.n465 71.676
R1128 B.n709 B.n466 71.676
R1129 B.n705 B.n467 71.676
R1130 B.n701 B.n468 71.676
R1131 B.n697 B.n469 71.676
R1132 B.n693 B.n470 71.676
R1133 B.n689 B.n471 71.676
R1134 B.n685 B.n472 71.676
R1135 B.n681 B.n473 71.676
R1136 B.n677 B.n474 71.676
R1137 B.n673 B.n475 71.676
R1138 B.n669 B.n476 71.676
R1139 B.n665 B.n477 71.676
R1140 B.n661 B.n478 71.676
R1141 B.n657 B.n479 71.676
R1142 B.n653 B.n480 71.676
R1143 B.n649 B.n481 71.676
R1144 B.n645 B.n482 71.676
R1145 B.n640 B.n483 71.676
R1146 B.n636 B.n484 71.676
R1147 B.n632 B.n485 71.676
R1148 B.n628 B.n486 71.676
R1149 B.n624 B.n487 71.676
R1150 B.n620 B.n488 71.676
R1151 B.n616 B.n489 71.676
R1152 B.n612 B.n490 71.676
R1153 B.n608 B.n491 71.676
R1154 B.n604 B.n492 71.676
R1155 B.n600 B.n493 71.676
R1156 B.n596 B.n494 71.676
R1157 B.n592 B.n495 71.676
R1158 B.n588 B.n496 71.676
R1159 B.n584 B.n497 71.676
R1160 B.n580 B.n498 71.676
R1161 B.n576 B.n499 71.676
R1162 B.n572 B.n500 71.676
R1163 B.n568 B.n501 71.676
R1164 B.n564 B.n502 71.676
R1165 B.n560 B.n503 71.676
R1166 B.n556 B.n504 71.676
R1167 B.n552 B.n505 71.676
R1168 B.n548 B.n506 71.676
R1169 B.n544 B.n507 71.676
R1170 B.n540 B.n508 71.676
R1171 B.n536 B.n509 71.676
R1172 B.n532 B.n510 71.676
R1173 B.n528 B.n511 71.676
R1174 B.n524 B.n512 71.676
R1175 B.n520 B.n513 71.676
R1176 B.n519 B.t11 69.9348
R1177 B.n128 B.t15 69.9348
R1178 B.n516 B.t4 69.9101
R1179 B.n131 B.t9 69.9101
R1180 B.n642 B.n519 59.5399
R1181 B.n517 B.n516 59.5399
R1182 B.n250 B.n131 59.5399
R1183 B.n129 B.n128 59.5399
R1184 B.n778 B.n446 51.357
R1185 B.n915 B.n57 51.357
R1186 B.n785 B.n446 31.4621
R1187 B.n785 B.n442 31.4621
R1188 B.n791 B.n442 31.4621
R1189 B.n791 B.n438 31.4621
R1190 B.n797 B.n438 31.4621
R1191 B.n797 B.n434 31.4621
R1192 B.n803 B.n434 31.4621
R1193 B.n803 B.n430 31.4621
R1194 B.n809 B.n430 31.4621
R1195 B.n815 B.n426 31.4621
R1196 B.n815 B.n422 31.4621
R1197 B.n821 B.n422 31.4621
R1198 B.n821 B.n418 31.4621
R1199 B.n827 B.n418 31.4621
R1200 B.n827 B.n414 31.4621
R1201 B.n833 B.n414 31.4621
R1202 B.n833 B.n410 31.4621
R1203 B.n839 B.n410 31.4621
R1204 B.n839 B.n406 31.4621
R1205 B.n845 B.n406 31.4621
R1206 B.n845 B.n402 31.4621
R1207 B.n851 B.n402 31.4621
R1208 B.n857 B.n398 31.4621
R1209 B.n857 B.n394 31.4621
R1210 B.n864 B.n394 31.4621
R1211 B.n864 B.n390 31.4621
R1212 B.n870 B.n390 31.4621
R1213 B.n870 B.n4 31.4621
R1214 B.n980 B.n4 31.4621
R1215 B.n980 B.n979 31.4621
R1216 B.n979 B.n978 31.4621
R1217 B.n978 B.n8 31.4621
R1218 B.n972 B.n8 31.4621
R1219 B.n972 B.n971 31.4621
R1220 B.n971 B.n970 31.4621
R1221 B.n970 B.n15 31.4621
R1222 B.n964 B.n963 31.4621
R1223 B.n963 B.n962 31.4621
R1224 B.n962 B.n22 31.4621
R1225 B.n956 B.n22 31.4621
R1226 B.n956 B.n955 31.4621
R1227 B.n955 B.n954 31.4621
R1228 B.n954 B.n29 31.4621
R1229 B.n948 B.n29 31.4621
R1230 B.n948 B.n947 31.4621
R1231 B.n947 B.n946 31.4621
R1232 B.n946 B.n36 31.4621
R1233 B.n940 B.n36 31.4621
R1234 B.n940 B.n939 31.4621
R1235 B.n938 B.n43 31.4621
R1236 B.n932 B.n43 31.4621
R1237 B.n932 B.n931 31.4621
R1238 B.n931 B.n930 31.4621
R1239 B.n930 B.n50 31.4621
R1240 B.n924 B.n50 31.4621
R1241 B.n924 B.n923 31.4621
R1242 B.n923 B.n922 31.4621
R1243 B.n922 B.n57 31.4621
R1244 B.n919 B.n918 30.7517
R1245 B.n521 B.n444 30.7517
R1246 B.n782 B.n781 30.7517
R1247 B.n913 B.n912 30.7517
R1248 B.t3 B.n426 26.3727
R1249 B.n939 B.t7 26.3727
R1250 B.n851 B.t1 22.6714
R1251 B.n964 B.t0 22.6714
R1252 B B.n982 18.0485
R1253 B.n918 B.n59 10.6151
R1254 B.n133 B.n59 10.6151
R1255 B.n134 B.n133 10.6151
R1256 B.n137 B.n134 10.6151
R1257 B.n138 B.n137 10.6151
R1258 B.n141 B.n138 10.6151
R1259 B.n142 B.n141 10.6151
R1260 B.n145 B.n142 10.6151
R1261 B.n146 B.n145 10.6151
R1262 B.n149 B.n146 10.6151
R1263 B.n150 B.n149 10.6151
R1264 B.n153 B.n150 10.6151
R1265 B.n154 B.n153 10.6151
R1266 B.n157 B.n154 10.6151
R1267 B.n158 B.n157 10.6151
R1268 B.n161 B.n158 10.6151
R1269 B.n162 B.n161 10.6151
R1270 B.n165 B.n162 10.6151
R1271 B.n166 B.n165 10.6151
R1272 B.n169 B.n166 10.6151
R1273 B.n170 B.n169 10.6151
R1274 B.n173 B.n170 10.6151
R1275 B.n174 B.n173 10.6151
R1276 B.n177 B.n174 10.6151
R1277 B.n178 B.n177 10.6151
R1278 B.n181 B.n178 10.6151
R1279 B.n182 B.n181 10.6151
R1280 B.n185 B.n182 10.6151
R1281 B.n186 B.n185 10.6151
R1282 B.n189 B.n186 10.6151
R1283 B.n190 B.n189 10.6151
R1284 B.n193 B.n190 10.6151
R1285 B.n194 B.n193 10.6151
R1286 B.n197 B.n194 10.6151
R1287 B.n198 B.n197 10.6151
R1288 B.n201 B.n198 10.6151
R1289 B.n202 B.n201 10.6151
R1290 B.n205 B.n202 10.6151
R1291 B.n206 B.n205 10.6151
R1292 B.n209 B.n206 10.6151
R1293 B.n210 B.n209 10.6151
R1294 B.n213 B.n210 10.6151
R1295 B.n214 B.n213 10.6151
R1296 B.n217 B.n214 10.6151
R1297 B.n218 B.n217 10.6151
R1298 B.n221 B.n218 10.6151
R1299 B.n222 B.n221 10.6151
R1300 B.n225 B.n222 10.6151
R1301 B.n226 B.n225 10.6151
R1302 B.n229 B.n226 10.6151
R1303 B.n230 B.n229 10.6151
R1304 B.n233 B.n230 10.6151
R1305 B.n234 B.n233 10.6151
R1306 B.n237 B.n234 10.6151
R1307 B.n238 B.n237 10.6151
R1308 B.n241 B.n238 10.6151
R1309 B.n242 B.n241 10.6151
R1310 B.n245 B.n242 10.6151
R1311 B.n246 B.n245 10.6151
R1312 B.n249 B.n246 10.6151
R1313 B.n254 B.n251 10.6151
R1314 B.n255 B.n254 10.6151
R1315 B.n258 B.n255 10.6151
R1316 B.n259 B.n258 10.6151
R1317 B.n262 B.n259 10.6151
R1318 B.n263 B.n262 10.6151
R1319 B.n266 B.n263 10.6151
R1320 B.n267 B.n266 10.6151
R1321 B.n271 B.n270 10.6151
R1322 B.n274 B.n271 10.6151
R1323 B.n275 B.n274 10.6151
R1324 B.n278 B.n275 10.6151
R1325 B.n279 B.n278 10.6151
R1326 B.n282 B.n279 10.6151
R1327 B.n283 B.n282 10.6151
R1328 B.n286 B.n283 10.6151
R1329 B.n287 B.n286 10.6151
R1330 B.n290 B.n287 10.6151
R1331 B.n291 B.n290 10.6151
R1332 B.n294 B.n291 10.6151
R1333 B.n295 B.n294 10.6151
R1334 B.n298 B.n295 10.6151
R1335 B.n299 B.n298 10.6151
R1336 B.n302 B.n299 10.6151
R1337 B.n303 B.n302 10.6151
R1338 B.n306 B.n303 10.6151
R1339 B.n307 B.n306 10.6151
R1340 B.n310 B.n307 10.6151
R1341 B.n311 B.n310 10.6151
R1342 B.n314 B.n311 10.6151
R1343 B.n315 B.n314 10.6151
R1344 B.n318 B.n315 10.6151
R1345 B.n319 B.n318 10.6151
R1346 B.n322 B.n319 10.6151
R1347 B.n323 B.n322 10.6151
R1348 B.n326 B.n323 10.6151
R1349 B.n327 B.n326 10.6151
R1350 B.n330 B.n327 10.6151
R1351 B.n331 B.n330 10.6151
R1352 B.n334 B.n331 10.6151
R1353 B.n335 B.n334 10.6151
R1354 B.n338 B.n335 10.6151
R1355 B.n339 B.n338 10.6151
R1356 B.n342 B.n339 10.6151
R1357 B.n343 B.n342 10.6151
R1358 B.n346 B.n343 10.6151
R1359 B.n347 B.n346 10.6151
R1360 B.n350 B.n347 10.6151
R1361 B.n351 B.n350 10.6151
R1362 B.n354 B.n351 10.6151
R1363 B.n355 B.n354 10.6151
R1364 B.n358 B.n355 10.6151
R1365 B.n359 B.n358 10.6151
R1366 B.n362 B.n359 10.6151
R1367 B.n363 B.n362 10.6151
R1368 B.n366 B.n363 10.6151
R1369 B.n367 B.n366 10.6151
R1370 B.n370 B.n367 10.6151
R1371 B.n371 B.n370 10.6151
R1372 B.n374 B.n371 10.6151
R1373 B.n375 B.n374 10.6151
R1374 B.n378 B.n375 10.6151
R1375 B.n379 B.n378 10.6151
R1376 B.n382 B.n379 10.6151
R1377 B.n383 B.n382 10.6151
R1378 B.n386 B.n383 10.6151
R1379 B.n387 B.n386 10.6151
R1380 B.n913 B.n387 10.6151
R1381 B.n787 B.n444 10.6151
R1382 B.n788 B.n787 10.6151
R1383 B.n789 B.n788 10.6151
R1384 B.n789 B.n436 10.6151
R1385 B.n799 B.n436 10.6151
R1386 B.n800 B.n799 10.6151
R1387 B.n801 B.n800 10.6151
R1388 B.n801 B.n428 10.6151
R1389 B.n811 B.n428 10.6151
R1390 B.n812 B.n811 10.6151
R1391 B.n813 B.n812 10.6151
R1392 B.n813 B.n420 10.6151
R1393 B.n823 B.n420 10.6151
R1394 B.n824 B.n823 10.6151
R1395 B.n825 B.n824 10.6151
R1396 B.n825 B.n412 10.6151
R1397 B.n835 B.n412 10.6151
R1398 B.n836 B.n835 10.6151
R1399 B.n837 B.n836 10.6151
R1400 B.n837 B.n404 10.6151
R1401 B.n847 B.n404 10.6151
R1402 B.n848 B.n847 10.6151
R1403 B.n849 B.n848 10.6151
R1404 B.n849 B.n396 10.6151
R1405 B.n859 B.n396 10.6151
R1406 B.n860 B.n859 10.6151
R1407 B.n862 B.n860 10.6151
R1408 B.n862 B.n861 10.6151
R1409 B.n861 B.n388 10.6151
R1410 B.n873 B.n388 10.6151
R1411 B.n874 B.n873 10.6151
R1412 B.n875 B.n874 10.6151
R1413 B.n876 B.n875 10.6151
R1414 B.n878 B.n876 10.6151
R1415 B.n879 B.n878 10.6151
R1416 B.n880 B.n879 10.6151
R1417 B.n881 B.n880 10.6151
R1418 B.n883 B.n881 10.6151
R1419 B.n884 B.n883 10.6151
R1420 B.n885 B.n884 10.6151
R1421 B.n886 B.n885 10.6151
R1422 B.n888 B.n886 10.6151
R1423 B.n889 B.n888 10.6151
R1424 B.n890 B.n889 10.6151
R1425 B.n891 B.n890 10.6151
R1426 B.n893 B.n891 10.6151
R1427 B.n894 B.n893 10.6151
R1428 B.n895 B.n894 10.6151
R1429 B.n896 B.n895 10.6151
R1430 B.n898 B.n896 10.6151
R1431 B.n899 B.n898 10.6151
R1432 B.n900 B.n899 10.6151
R1433 B.n901 B.n900 10.6151
R1434 B.n903 B.n901 10.6151
R1435 B.n904 B.n903 10.6151
R1436 B.n905 B.n904 10.6151
R1437 B.n906 B.n905 10.6151
R1438 B.n908 B.n906 10.6151
R1439 B.n909 B.n908 10.6151
R1440 B.n910 B.n909 10.6151
R1441 B.n911 B.n910 10.6151
R1442 B.n912 B.n911 10.6151
R1443 B.n781 B.n448 10.6151
R1444 B.n776 B.n448 10.6151
R1445 B.n776 B.n775 10.6151
R1446 B.n775 B.n774 10.6151
R1447 B.n774 B.n771 10.6151
R1448 B.n771 B.n770 10.6151
R1449 B.n770 B.n767 10.6151
R1450 B.n767 B.n766 10.6151
R1451 B.n766 B.n763 10.6151
R1452 B.n763 B.n762 10.6151
R1453 B.n762 B.n759 10.6151
R1454 B.n759 B.n758 10.6151
R1455 B.n758 B.n755 10.6151
R1456 B.n755 B.n754 10.6151
R1457 B.n754 B.n751 10.6151
R1458 B.n751 B.n750 10.6151
R1459 B.n750 B.n747 10.6151
R1460 B.n747 B.n746 10.6151
R1461 B.n746 B.n743 10.6151
R1462 B.n743 B.n742 10.6151
R1463 B.n742 B.n739 10.6151
R1464 B.n739 B.n738 10.6151
R1465 B.n738 B.n735 10.6151
R1466 B.n735 B.n734 10.6151
R1467 B.n734 B.n731 10.6151
R1468 B.n731 B.n730 10.6151
R1469 B.n730 B.n727 10.6151
R1470 B.n727 B.n726 10.6151
R1471 B.n726 B.n723 10.6151
R1472 B.n723 B.n722 10.6151
R1473 B.n722 B.n719 10.6151
R1474 B.n719 B.n718 10.6151
R1475 B.n718 B.n715 10.6151
R1476 B.n715 B.n714 10.6151
R1477 B.n714 B.n711 10.6151
R1478 B.n711 B.n710 10.6151
R1479 B.n710 B.n707 10.6151
R1480 B.n707 B.n706 10.6151
R1481 B.n706 B.n703 10.6151
R1482 B.n703 B.n702 10.6151
R1483 B.n702 B.n699 10.6151
R1484 B.n699 B.n698 10.6151
R1485 B.n698 B.n695 10.6151
R1486 B.n695 B.n694 10.6151
R1487 B.n694 B.n691 10.6151
R1488 B.n691 B.n690 10.6151
R1489 B.n690 B.n687 10.6151
R1490 B.n687 B.n686 10.6151
R1491 B.n686 B.n683 10.6151
R1492 B.n683 B.n682 10.6151
R1493 B.n682 B.n679 10.6151
R1494 B.n679 B.n678 10.6151
R1495 B.n678 B.n675 10.6151
R1496 B.n675 B.n674 10.6151
R1497 B.n674 B.n671 10.6151
R1498 B.n671 B.n670 10.6151
R1499 B.n670 B.n667 10.6151
R1500 B.n667 B.n666 10.6151
R1501 B.n666 B.n663 10.6151
R1502 B.n663 B.n662 10.6151
R1503 B.n659 B.n658 10.6151
R1504 B.n658 B.n655 10.6151
R1505 B.n655 B.n654 10.6151
R1506 B.n654 B.n651 10.6151
R1507 B.n651 B.n650 10.6151
R1508 B.n650 B.n647 10.6151
R1509 B.n647 B.n646 10.6151
R1510 B.n646 B.n643 10.6151
R1511 B.n641 B.n638 10.6151
R1512 B.n638 B.n637 10.6151
R1513 B.n637 B.n634 10.6151
R1514 B.n634 B.n633 10.6151
R1515 B.n633 B.n630 10.6151
R1516 B.n630 B.n629 10.6151
R1517 B.n629 B.n626 10.6151
R1518 B.n626 B.n625 10.6151
R1519 B.n625 B.n622 10.6151
R1520 B.n622 B.n621 10.6151
R1521 B.n621 B.n618 10.6151
R1522 B.n618 B.n617 10.6151
R1523 B.n617 B.n614 10.6151
R1524 B.n614 B.n613 10.6151
R1525 B.n613 B.n610 10.6151
R1526 B.n610 B.n609 10.6151
R1527 B.n609 B.n606 10.6151
R1528 B.n606 B.n605 10.6151
R1529 B.n605 B.n602 10.6151
R1530 B.n602 B.n601 10.6151
R1531 B.n601 B.n598 10.6151
R1532 B.n598 B.n597 10.6151
R1533 B.n597 B.n594 10.6151
R1534 B.n594 B.n593 10.6151
R1535 B.n593 B.n590 10.6151
R1536 B.n590 B.n589 10.6151
R1537 B.n589 B.n586 10.6151
R1538 B.n586 B.n585 10.6151
R1539 B.n585 B.n582 10.6151
R1540 B.n582 B.n581 10.6151
R1541 B.n581 B.n578 10.6151
R1542 B.n578 B.n577 10.6151
R1543 B.n577 B.n574 10.6151
R1544 B.n574 B.n573 10.6151
R1545 B.n573 B.n570 10.6151
R1546 B.n570 B.n569 10.6151
R1547 B.n569 B.n566 10.6151
R1548 B.n566 B.n565 10.6151
R1549 B.n565 B.n562 10.6151
R1550 B.n562 B.n561 10.6151
R1551 B.n561 B.n558 10.6151
R1552 B.n558 B.n557 10.6151
R1553 B.n557 B.n554 10.6151
R1554 B.n554 B.n553 10.6151
R1555 B.n553 B.n550 10.6151
R1556 B.n550 B.n549 10.6151
R1557 B.n549 B.n546 10.6151
R1558 B.n546 B.n545 10.6151
R1559 B.n545 B.n542 10.6151
R1560 B.n542 B.n541 10.6151
R1561 B.n541 B.n538 10.6151
R1562 B.n538 B.n537 10.6151
R1563 B.n537 B.n534 10.6151
R1564 B.n534 B.n533 10.6151
R1565 B.n533 B.n530 10.6151
R1566 B.n530 B.n529 10.6151
R1567 B.n529 B.n526 10.6151
R1568 B.n526 B.n525 10.6151
R1569 B.n525 B.n522 10.6151
R1570 B.n522 B.n521 10.6151
R1571 B.n783 B.n782 10.6151
R1572 B.n783 B.n440 10.6151
R1573 B.n793 B.n440 10.6151
R1574 B.n794 B.n793 10.6151
R1575 B.n795 B.n794 10.6151
R1576 B.n795 B.n432 10.6151
R1577 B.n805 B.n432 10.6151
R1578 B.n806 B.n805 10.6151
R1579 B.n807 B.n806 10.6151
R1580 B.n807 B.n424 10.6151
R1581 B.n817 B.n424 10.6151
R1582 B.n818 B.n817 10.6151
R1583 B.n819 B.n818 10.6151
R1584 B.n819 B.n416 10.6151
R1585 B.n829 B.n416 10.6151
R1586 B.n830 B.n829 10.6151
R1587 B.n831 B.n830 10.6151
R1588 B.n831 B.n408 10.6151
R1589 B.n841 B.n408 10.6151
R1590 B.n842 B.n841 10.6151
R1591 B.n843 B.n842 10.6151
R1592 B.n843 B.n400 10.6151
R1593 B.n853 B.n400 10.6151
R1594 B.n854 B.n853 10.6151
R1595 B.n855 B.n854 10.6151
R1596 B.n855 B.n392 10.6151
R1597 B.n866 B.n392 10.6151
R1598 B.n867 B.n866 10.6151
R1599 B.n868 B.n867 10.6151
R1600 B.n868 B.n0 10.6151
R1601 B.n976 B.n1 10.6151
R1602 B.n976 B.n975 10.6151
R1603 B.n975 B.n974 10.6151
R1604 B.n974 B.n10 10.6151
R1605 B.n968 B.n10 10.6151
R1606 B.n968 B.n967 10.6151
R1607 B.n967 B.n966 10.6151
R1608 B.n966 B.n17 10.6151
R1609 B.n960 B.n17 10.6151
R1610 B.n960 B.n959 10.6151
R1611 B.n959 B.n958 10.6151
R1612 B.n958 B.n24 10.6151
R1613 B.n952 B.n24 10.6151
R1614 B.n952 B.n951 10.6151
R1615 B.n951 B.n950 10.6151
R1616 B.n950 B.n31 10.6151
R1617 B.n944 B.n31 10.6151
R1618 B.n944 B.n943 10.6151
R1619 B.n943 B.n942 10.6151
R1620 B.n942 B.n38 10.6151
R1621 B.n936 B.n38 10.6151
R1622 B.n936 B.n935 10.6151
R1623 B.n935 B.n934 10.6151
R1624 B.n934 B.n45 10.6151
R1625 B.n928 B.n45 10.6151
R1626 B.n928 B.n927 10.6151
R1627 B.n927 B.n926 10.6151
R1628 B.n926 B.n52 10.6151
R1629 B.n920 B.n52 10.6151
R1630 B.n920 B.n919 10.6151
R1631 B.t1 B.n398 8.79125
R1632 B.t0 B.n15 8.79125
R1633 B.n251 B.n250 6.5566
R1634 B.n267 B.n129 6.5566
R1635 B.n659 B.n517 6.5566
R1636 B.n643 B.n642 6.5566
R1637 B.n809 B.t3 5.08988
R1638 B.t7 B.n938 5.08988
R1639 B.n250 B.n249 4.05904
R1640 B.n270 B.n129 4.05904
R1641 B.n662 B.n517 4.05904
R1642 B.n642 B.n641 4.05904
R1643 B.n982 B.n0 2.81026
R1644 B.n982 B.n1 2.81026
R1645 VP.n0 VP.t0 217.196
R1646 VP.n0 VP.t1 165.149
R1647 VP VP.n0 0.526373
R1648 VTAIL.n1 VTAIL.t1 43.0861
R1649 VTAIL.n3 VTAIL.t0 43.086
R1650 VTAIL.n0 VTAIL.t2 43.086
R1651 VTAIL.n2 VTAIL.t3 43.086
R1652 VTAIL.n1 VTAIL.n0 34.9703
R1653 VTAIL.n3 VTAIL.n2 31.6427
R1654 VTAIL.n2 VTAIL.n1 2.13412
R1655 VTAIL VTAIL.n0 1.36041
R1656 VTAIL VTAIL.n3 0.774207
R1657 VDD1 VDD1.t0 107.385
R1658 VDD1 VDD1.t1 60.6549
R1659 VN VN.t0 217.103
R1660 VN VN.t1 165.675
R1661 VDD2.n0 VDD2.t0 106.028
R1662 VDD2.n0 VDD2.t1 59.7648
R1663 VDD2 VDD2.n0 0.890586
C0 VDD1 VP 4.54888f
C1 VN VTAIL 3.74648f
C2 VN VDD2 4.32792f
C3 VTAIL VDD2 6.9392f
C4 VN VP 7.090549f
C5 VTAIL VP 3.76077f
C6 VN VDD1 0.148883f
C7 VTAIL VDD1 6.88266f
C8 VP VDD2 0.372881f
C9 VDD1 VDD2 0.776924f
C10 VDD2 B 5.932191f
C11 VDD1 B 9.69981f
C12 VTAIL B 10.478756f
C13 VN B 13.07365f
C14 VP B 7.982452f
C15 VDD2.t0 B 4.17576f
C16 VDD2.t1 B 3.38452f
C17 VDD2.n0 B 3.47556f
C18 VN.t1 B 4.68644f
C19 VN.t0 B 5.36279f
C20 VDD1.t1 B 3.42681f
C21 VDD1.t0 B 4.27078f
C22 VTAIL.t2 B 3.29597f
C23 VTAIL.n0 B 2.08599f
C24 VTAIL.t1 B 3.29599f
C25 VTAIL.n1 B 2.13549f
C26 VTAIL.t3 B 3.29597f
C27 VTAIL.n2 B 1.92254f
C28 VTAIL.t0 B 3.29597f
C29 VTAIL.n3 B 1.8355f
C30 VP.t0 B 5.48189f
C31 VP.t1 B 4.78551f
C32 VP.n0 B 5.04067f
.ends

