* NGSPICE file created from diff_pair_sample_0587.ext - technology: sky130A

.subckt diff_pair_sample_0587 VTAIL VN VP B VDD2 VDD1
X0 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=5.6043 pd=29.52 as=0 ps=0 w=14.37 l=1.97
X1 VDD2.t3 VN.t0 VTAIL.t7 B.t0 sky130_fd_pr__nfet_01v8 ad=2.37105 pd=14.7 as=5.6043 ps=29.52 w=14.37 l=1.97
X2 VTAIL.t5 VN.t1 VDD2.t2 B.t17 sky130_fd_pr__nfet_01v8 ad=5.6043 pd=29.52 as=2.37105 ps=14.7 w=14.37 l=1.97
X3 VTAIL.t1 VP.t0 VDD1.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=5.6043 pd=29.52 as=2.37105 ps=14.7 w=14.37 l=1.97
X4 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=5.6043 pd=29.52 as=0 ps=0 w=14.37 l=1.97
X5 VTAIL.t3 VP.t1 VDD1.t2 B.t17 sky130_fd_pr__nfet_01v8 ad=5.6043 pd=29.52 as=2.37105 ps=14.7 w=14.37 l=1.97
X6 B.t9 B.t7 B.t8 B.t4 sky130_fd_pr__nfet_01v8 ad=5.6043 pd=29.52 as=0 ps=0 w=14.37 l=1.97
X7 B.t6 B.t3 B.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=5.6043 pd=29.52 as=0 ps=0 w=14.37 l=1.97
X8 VDD1.t1 VP.t2 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=2.37105 pd=14.7 as=5.6043 ps=29.52 w=14.37 l=1.97
X9 VDD2.t1 VN.t2 VTAIL.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=2.37105 pd=14.7 as=5.6043 ps=29.52 w=14.37 l=1.97
X10 VTAIL.t4 VN.t3 VDD2.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=5.6043 pd=29.52 as=2.37105 ps=14.7 w=14.37 l=1.97
X11 VDD1.t0 VP.t3 VTAIL.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=2.37105 pd=14.7 as=5.6043 ps=29.52 w=14.37 l=1.97
R0 B.n775 B.n774 585
R1 B.n776 B.n775 585
R2 B.n324 B.n109 585
R3 B.n323 B.n322 585
R4 B.n321 B.n320 585
R5 B.n319 B.n318 585
R6 B.n317 B.n316 585
R7 B.n315 B.n314 585
R8 B.n313 B.n312 585
R9 B.n311 B.n310 585
R10 B.n309 B.n308 585
R11 B.n307 B.n306 585
R12 B.n305 B.n304 585
R13 B.n303 B.n302 585
R14 B.n301 B.n300 585
R15 B.n299 B.n298 585
R16 B.n297 B.n296 585
R17 B.n295 B.n294 585
R18 B.n293 B.n292 585
R19 B.n291 B.n290 585
R20 B.n289 B.n288 585
R21 B.n287 B.n286 585
R22 B.n285 B.n284 585
R23 B.n283 B.n282 585
R24 B.n281 B.n280 585
R25 B.n279 B.n278 585
R26 B.n277 B.n276 585
R27 B.n275 B.n274 585
R28 B.n273 B.n272 585
R29 B.n271 B.n270 585
R30 B.n269 B.n268 585
R31 B.n267 B.n266 585
R32 B.n265 B.n264 585
R33 B.n263 B.n262 585
R34 B.n261 B.n260 585
R35 B.n259 B.n258 585
R36 B.n257 B.n256 585
R37 B.n255 B.n254 585
R38 B.n253 B.n252 585
R39 B.n251 B.n250 585
R40 B.n249 B.n248 585
R41 B.n247 B.n246 585
R42 B.n245 B.n244 585
R43 B.n243 B.n242 585
R44 B.n241 B.n240 585
R45 B.n239 B.n238 585
R46 B.n237 B.n236 585
R47 B.n235 B.n234 585
R48 B.n233 B.n232 585
R49 B.n231 B.n230 585
R50 B.n229 B.n228 585
R51 B.n227 B.n226 585
R52 B.n225 B.n224 585
R53 B.n223 B.n222 585
R54 B.n221 B.n220 585
R55 B.n219 B.n218 585
R56 B.n217 B.n216 585
R57 B.n215 B.n214 585
R58 B.n213 B.n212 585
R59 B.n210 B.n209 585
R60 B.n208 B.n207 585
R61 B.n206 B.n205 585
R62 B.n204 B.n203 585
R63 B.n202 B.n201 585
R64 B.n200 B.n199 585
R65 B.n198 B.n197 585
R66 B.n196 B.n195 585
R67 B.n194 B.n193 585
R68 B.n192 B.n191 585
R69 B.n190 B.n189 585
R70 B.n188 B.n187 585
R71 B.n186 B.n185 585
R72 B.n184 B.n183 585
R73 B.n182 B.n181 585
R74 B.n180 B.n179 585
R75 B.n178 B.n177 585
R76 B.n176 B.n175 585
R77 B.n174 B.n173 585
R78 B.n172 B.n171 585
R79 B.n170 B.n169 585
R80 B.n168 B.n167 585
R81 B.n166 B.n165 585
R82 B.n164 B.n163 585
R83 B.n162 B.n161 585
R84 B.n160 B.n159 585
R85 B.n158 B.n157 585
R86 B.n156 B.n155 585
R87 B.n154 B.n153 585
R88 B.n152 B.n151 585
R89 B.n150 B.n149 585
R90 B.n148 B.n147 585
R91 B.n146 B.n145 585
R92 B.n144 B.n143 585
R93 B.n142 B.n141 585
R94 B.n140 B.n139 585
R95 B.n138 B.n137 585
R96 B.n136 B.n135 585
R97 B.n134 B.n133 585
R98 B.n132 B.n131 585
R99 B.n130 B.n129 585
R100 B.n128 B.n127 585
R101 B.n126 B.n125 585
R102 B.n124 B.n123 585
R103 B.n122 B.n121 585
R104 B.n120 B.n119 585
R105 B.n118 B.n117 585
R106 B.n116 B.n115 585
R107 B.n54 B.n53 585
R108 B.n773 B.n55 585
R109 B.n777 B.n55 585
R110 B.n772 B.n771 585
R111 B.n771 B.n51 585
R112 B.n770 B.n50 585
R113 B.n783 B.n50 585
R114 B.n769 B.n49 585
R115 B.n784 B.n49 585
R116 B.n768 B.n48 585
R117 B.n785 B.n48 585
R118 B.n767 B.n766 585
R119 B.n766 B.n44 585
R120 B.n765 B.n43 585
R121 B.n791 B.n43 585
R122 B.n764 B.n42 585
R123 B.n792 B.n42 585
R124 B.n763 B.n41 585
R125 B.n793 B.n41 585
R126 B.n762 B.n761 585
R127 B.n761 B.n37 585
R128 B.n760 B.n36 585
R129 B.n799 B.n36 585
R130 B.n759 B.n35 585
R131 B.n800 B.n35 585
R132 B.n758 B.n34 585
R133 B.n801 B.n34 585
R134 B.n757 B.n756 585
R135 B.n756 B.n30 585
R136 B.n755 B.n29 585
R137 B.n807 B.n29 585
R138 B.n754 B.n28 585
R139 B.n808 B.n28 585
R140 B.n753 B.n27 585
R141 B.n809 B.n27 585
R142 B.n752 B.n751 585
R143 B.n751 B.n23 585
R144 B.n750 B.n22 585
R145 B.n815 B.n22 585
R146 B.n749 B.n21 585
R147 B.n816 B.n21 585
R148 B.n748 B.n20 585
R149 B.n817 B.n20 585
R150 B.n747 B.n746 585
R151 B.n746 B.n16 585
R152 B.n745 B.n15 585
R153 B.n823 B.n15 585
R154 B.n744 B.n14 585
R155 B.n824 B.n14 585
R156 B.n743 B.n13 585
R157 B.n825 B.n13 585
R158 B.n742 B.n741 585
R159 B.n741 B.n12 585
R160 B.n740 B.n739 585
R161 B.n740 B.n8 585
R162 B.n738 B.n7 585
R163 B.n832 B.n7 585
R164 B.n737 B.n6 585
R165 B.n833 B.n6 585
R166 B.n736 B.n5 585
R167 B.n834 B.n5 585
R168 B.n735 B.n734 585
R169 B.n734 B.n4 585
R170 B.n733 B.n325 585
R171 B.n733 B.n732 585
R172 B.n723 B.n326 585
R173 B.n327 B.n326 585
R174 B.n725 B.n724 585
R175 B.n726 B.n725 585
R176 B.n722 B.n331 585
R177 B.n335 B.n331 585
R178 B.n721 B.n720 585
R179 B.n720 B.n719 585
R180 B.n333 B.n332 585
R181 B.n334 B.n333 585
R182 B.n712 B.n711 585
R183 B.n713 B.n712 585
R184 B.n710 B.n340 585
R185 B.n340 B.n339 585
R186 B.n709 B.n708 585
R187 B.n708 B.n707 585
R188 B.n342 B.n341 585
R189 B.n343 B.n342 585
R190 B.n700 B.n699 585
R191 B.n701 B.n700 585
R192 B.n698 B.n348 585
R193 B.n348 B.n347 585
R194 B.n697 B.n696 585
R195 B.n696 B.n695 585
R196 B.n350 B.n349 585
R197 B.n351 B.n350 585
R198 B.n688 B.n687 585
R199 B.n689 B.n688 585
R200 B.n686 B.n356 585
R201 B.n356 B.n355 585
R202 B.n685 B.n684 585
R203 B.n684 B.n683 585
R204 B.n358 B.n357 585
R205 B.n359 B.n358 585
R206 B.n676 B.n675 585
R207 B.n677 B.n676 585
R208 B.n674 B.n364 585
R209 B.n364 B.n363 585
R210 B.n673 B.n672 585
R211 B.n672 B.n671 585
R212 B.n366 B.n365 585
R213 B.n367 B.n366 585
R214 B.n664 B.n663 585
R215 B.n665 B.n664 585
R216 B.n662 B.n372 585
R217 B.n372 B.n371 585
R218 B.n661 B.n660 585
R219 B.n660 B.n659 585
R220 B.n374 B.n373 585
R221 B.n375 B.n374 585
R222 B.n652 B.n651 585
R223 B.n653 B.n652 585
R224 B.n378 B.n377 585
R225 B.n440 B.n439 585
R226 B.n441 B.n437 585
R227 B.n437 B.n379 585
R228 B.n443 B.n442 585
R229 B.n445 B.n436 585
R230 B.n448 B.n447 585
R231 B.n449 B.n435 585
R232 B.n451 B.n450 585
R233 B.n453 B.n434 585
R234 B.n456 B.n455 585
R235 B.n457 B.n433 585
R236 B.n459 B.n458 585
R237 B.n461 B.n432 585
R238 B.n464 B.n463 585
R239 B.n465 B.n431 585
R240 B.n467 B.n466 585
R241 B.n469 B.n430 585
R242 B.n472 B.n471 585
R243 B.n473 B.n429 585
R244 B.n475 B.n474 585
R245 B.n477 B.n428 585
R246 B.n480 B.n479 585
R247 B.n481 B.n427 585
R248 B.n483 B.n482 585
R249 B.n485 B.n426 585
R250 B.n488 B.n487 585
R251 B.n489 B.n425 585
R252 B.n491 B.n490 585
R253 B.n493 B.n424 585
R254 B.n496 B.n495 585
R255 B.n497 B.n423 585
R256 B.n499 B.n498 585
R257 B.n501 B.n422 585
R258 B.n504 B.n503 585
R259 B.n505 B.n421 585
R260 B.n507 B.n506 585
R261 B.n509 B.n420 585
R262 B.n512 B.n511 585
R263 B.n513 B.n419 585
R264 B.n515 B.n514 585
R265 B.n517 B.n418 585
R266 B.n520 B.n519 585
R267 B.n521 B.n417 585
R268 B.n523 B.n522 585
R269 B.n525 B.n416 585
R270 B.n528 B.n527 585
R271 B.n529 B.n415 585
R272 B.n531 B.n530 585
R273 B.n533 B.n414 585
R274 B.n536 B.n535 585
R275 B.n537 B.n410 585
R276 B.n539 B.n538 585
R277 B.n541 B.n409 585
R278 B.n544 B.n543 585
R279 B.n545 B.n408 585
R280 B.n547 B.n546 585
R281 B.n549 B.n407 585
R282 B.n552 B.n551 585
R283 B.n554 B.n404 585
R284 B.n556 B.n555 585
R285 B.n558 B.n403 585
R286 B.n561 B.n560 585
R287 B.n562 B.n402 585
R288 B.n564 B.n563 585
R289 B.n566 B.n401 585
R290 B.n569 B.n568 585
R291 B.n570 B.n400 585
R292 B.n572 B.n571 585
R293 B.n574 B.n399 585
R294 B.n577 B.n576 585
R295 B.n578 B.n398 585
R296 B.n580 B.n579 585
R297 B.n582 B.n397 585
R298 B.n585 B.n584 585
R299 B.n586 B.n396 585
R300 B.n588 B.n587 585
R301 B.n590 B.n395 585
R302 B.n593 B.n592 585
R303 B.n594 B.n394 585
R304 B.n596 B.n595 585
R305 B.n598 B.n393 585
R306 B.n601 B.n600 585
R307 B.n602 B.n392 585
R308 B.n604 B.n603 585
R309 B.n606 B.n391 585
R310 B.n609 B.n608 585
R311 B.n610 B.n390 585
R312 B.n612 B.n611 585
R313 B.n614 B.n389 585
R314 B.n617 B.n616 585
R315 B.n618 B.n388 585
R316 B.n620 B.n619 585
R317 B.n622 B.n387 585
R318 B.n625 B.n624 585
R319 B.n626 B.n386 585
R320 B.n628 B.n627 585
R321 B.n630 B.n385 585
R322 B.n633 B.n632 585
R323 B.n634 B.n384 585
R324 B.n636 B.n635 585
R325 B.n638 B.n383 585
R326 B.n641 B.n640 585
R327 B.n642 B.n382 585
R328 B.n644 B.n643 585
R329 B.n646 B.n381 585
R330 B.n649 B.n648 585
R331 B.n650 B.n380 585
R332 B.n655 B.n654 585
R333 B.n654 B.n653 585
R334 B.n656 B.n376 585
R335 B.n376 B.n375 585
R336 B.n658 B.n657 585
R337 B.n659 B.n658 585
R338 B.n370 B.n369 585
R339 B.n371 B.n370 585
R340 B.n667 B.n666 585
R341 B.n666 B.n665 585
R342 B.n668 B.n368 585
R343 B.n368 B.n367 585
R344 B.n670 B.n669 585
R345 B.n671 B.n670 585
R346 B.n362 B.n361 585
R347 B.n363 B.n362 585
R348 B.n679 B.n678 585
R349 B.n678 B.n677 585
R350 B.n680 B.n360 585
R351 B.n360 B.n359 585
R352 B.n682 B.n681 585
R353 B.n683 B.n682 585
R354 B.n354 B.n353 585
R355 B.n355 B.n354 585
R356 B.n691 B.n690 585
R357 B.n690 B.n689 585
R358 B.n692 B.n352 585
R359 B.n352 B.n351 585
R360 B.n694 B.n693 585
R361 B.n695 B.n694 585
R362 B.n346 B.n345 585
R363 B.n347 B.n346 585
R364 B.n703 B.n702 585
R365 B.n702 B.n701 585
R366 B.n704 B.n344 585
R367 B.n344 B.n343 585
R368 B.n706 B.n705 585
R369 B.n707 B.n706 585
R370 B.n338 B.n337 585
R371 B.n339 B.n338 585
R372 B.n715 B.n714 585
R373 B.n714 B.n713 585
R374 B.n716 B.n336 585
R375 B.n336 B.n334 585
R376 B.n718 B.n717 585
R377 B.n719 B.n718 585
R378 B.n330 B.n329 585
R379 B.n335 B.n330 585
R380 B.n728 B.n727 585
R381 B.n727 B.n726 585
R382 B.n729 B.n328 585
R383 B.n328 B.n327 585
R384 B.n731 B.n730 585
R385 B.n732 B.n731 585
R386 B.n3 B.n0 585
R387 B.n4 B.n3 585
R388 B.n831 B.n1 585
R389 B.n832 B.n831 585
R390 B.n830 B.n829 585
R391 B.n830 B.n8 585
R392 B.n828 B.n9 585
R393 B.n12 B.n9 585
R394 B.n827 B.n826 585
R395 B.n826 B.n825 585
R396 B.n11 B.n10 585
R397 B.n824 B.n11 585
R398 B.n822 B.n821 585
R399 B.n823 B.n822 585
R400 B.n820 B.n17 585
R401 B.n17 B.n16 585
R402 B.n819 B.n818 585
R403 B.n818 B.n817 585
R404 B.n19 B.n18 585
R405 B.n816 B.n19 585
R406 B.n814 B.n813 585
R407 B.n815 B.n814 585
R408 B.n812 B.n24 585
R409 B.n24 B.n23 585
R410 B.n811 B.n810 585
R411 B.n810 B.n809 585
R412 B.n26 B.n25 585
R413 B.n808 B.n26 585
R414 B.n806 B.n805 585
R415 B.n807 B.n806 585
R416 B.n804 B.n31 585
R417 B.n31 B.n30 585
R418 B.n803 B.n802 585
R419 B.n802 B.n801 585
R420 B.n33 B.n32 585
R421 B.n800 B.n33 585
R422 B.n798 B.n797 585
R423 B.n799 B.n798 585
R424 B.n796 B.n38 585
R425 B.n38 B.n37 585
R426 B.n795 B.n794 585
R427 B.n794 B.n793 585
R428 B.n40 B.n39 585
R429 B.n792 B.n40 585
R430 B.n790 B.n789 585
R431 B.n791 B.n790 585
R432 B.n788 B.n45 585
R433 B.n45 B.n44 585
R434 B.n787 B.n786 585
R435 B.n786 B.n785 585
R436 B.n47 B.n46 585
R437 B.n784 B.n47 585
R438 B.n782 B.n781 585
R439 B.n783 B.n782 585
R440 B.n780 B.n52 585
R441 B.n52 B.n51 585
R442 B.n779 B.n778 585
R443 B.n778 B.n777 585
R444 B.n835 B.n834 585
R445 B.n833 B.n2 585
R446 B.n778 B.n54 463.671
R447 B.n775 B.n55 463.671
R448 B.n652 B.n380 463.671
R449 B.n654 B.n378 463.671
R450 B.n113 B.t3 382.642
R451 B.n110 B.t7 382.642
R452 B.n405 B.t10 382.642
R453 B.n411 B.t14 382.642
R454 B.n776 B.n108 256.663
R455 B.n776 B.n107 256.663
R456 B.n776 B.n106 256.663
R457 B.n776 B.n105 256.663
R458 B.n776 B.n104 256.663
R459 B.n776 B.n103 256.663
R460 B.n776 B.n102 256.663
R461 B.n776 B.n101 256.663
R462 B.n776 B.n100 256.663
R463 B.n776 B.n99 256.663
R464 B.n776 B.n98 256.663
R465 B.n776 B.n97 256.663
R466 B.n776 B.n96 256.663
R467 B.n776 B.n95 256.663
R468 B.n776 B.n94 256.663
R469 B.n776 B.n93 256.663
R470 B.n776 B.n92 256.663
R471 B.n776 B.n91 256.663
R472 B.n776 B.n90 256.663
R473 B.n776 B.n89 256.663
R474 B.n776 B.n88 256.663
R475 B.n776 B.n87 256.663
R476 B.n776 B.n86 256.663
R477 B.n776 B.n85 256.663
R478 B.n776 B.n84 256.663
R479 B.n776 B.n83 256.663
R480 B.n776 B.n82 256.663
R481 B.n776 B.n81 256.663
R482 B.n776 B.n80 256.663
R483 B.n776 B.n79 256.663
R484 B.n776 B.n78 256.663
R485 B.n776 B.n77 256.663
R486 B.n776 B.n76 256.663
R487 B.n776 B.n75 256.663
R488 B.n776 B.n74 256.663
R489 B.n776 B.n73 256.663
R490 B.n776 B.n72 256.663
R491 B.n776 B.n71 256.663
R492 B.n776 B.n70 256.663
R493 B.n776 B.n69 256.663
R494 B.n776 B.n68 256.663
R495 B.n776 B.n67 256.663
R496 B.n776 B.n66 256.663
R497 B.n776 B.n65 256.663
R498 B.n776 B.n64 256.663
R499 B.n776 B.n63 256.663
R500 B.n776 B.n62 256.663
R501 B.n776 B.n61 256.663
R502 B.n776 B.n60 256.663
R503 B.n776 B.n59 256.663
R504 B.n776 B.n58 256.663
R505 B.n776 B.n57 256.663
R506 B.n776 B.n56 256.663
R507 B.n438 B.n379 256.663
R508 B.n444 B.n379 256.663
R509 B.n446 B.n379 256.663
R510 B.n452 B.n379 256.663
R511 B.n454 B.n379 256.663
R512 B.n460 B.n379 256.663
R513 B.n462 B.n379 256.663
R514 B.n468 B.n379 256.663
R515 B.n470 B.n379 256.663
R516 B.n476 B.n379 256.663
R517 B.n478 B.n379 256.663
R518 B.n484 B.n379 256.663
R519 B.n486 B.n379 256.663
R520 B.n492 B.n379 256.663
R521 B.n494 B.n379 256.663
R522 B.n500 B.n379 256.663
R523 B.n502 B.n379 256.663
R524 B.n508 B.n379 256.663
R525 B.n510 B.n379 256.663
R526 B.n516 B.n379 256.663
R527 B.n518 B.n379 256.663
R528 B.n524 B.n379 256.663
R529 B.n526 B.n379 256.663
R530 B.n532 B.n379 256.663
R531 B.n534 B.n379 256.663
R532 B.n540 B.n379 256.663
R533 B.n542 B.n379 256.663
R534 B.n548 B.n379 256.663
R535 B.n550 B.n379 256.663
R536 B.n557 B.n379 256.663
R537 B.n559 B.n379 256.663
R538 B.n565 B.n379 256.663
R539 B.n567 B.n379 256.663
R540 B.n573 B.n379 256.663
R541 B.n575 B.n379 256.663
R542 B.n581 B.n379 256.663
R543 B.n583 B.n379 256.663
R544 B.n589 B.n379 256.663
R545 B.n591 B.n379 256.663
R546 B.n597 B.n379 256.663
R547 B.n599 B.n379 256.663
R548 B.n605 B.n379 256.663
R549 B.n607 B.n379 256.663
R550 B.n613 B.n379 256.663
R551 B.n615 B.n379 256.663
R552 B.n621 B.n379 256.663
R553 B.n623 B.n379 256.663
R554 B.n629 B.n379 256.663
R555 B.n631 B.n379 256.663
R556 B.n637 B.n379 256.663
R557 B.n639 B.n379 256.663
R558 B.n645 B.n379 256.663
R559 B.n647 B.n379 256.663
R560 B.n837 B.n836 256.663
R561 B.n117 B.n116 163.367
R562 B.n121 B.n120 163.367
R563 B.n125 B.n124 163.367
R564 B.n129 B.n128 163.367
R565 B.n133 B.n132 163.367
R566 B.n137 B.n136 163.367
R567 B.n141 B.n140 163.367
R568 B.n145 B.n144 163.367
R569 B.n149 B.n148 163.367
R570 B.n153 B.n152 163.367
R571 B.n157 B.n156 163.367
R572 B.n161 B.n160 163.367
R573 B.n165 B.n164 163.367
R574 B.n169 B.n168 163.367
R575 B.n173 B.n172 163.367
R576 B.n177 B.n176 163.367
R577 B.n181 B.n180 163.367
R578 B.n185 B.n184 163.367
R579 B.n189 B.n188 163.367
R580 B.n193 B.n192 163.367
R581 B.n197 B.n196 163.367
R582 B.n201 B.n200 163.367
R583 B.n205 B.n204 163.367
R584 B.n209 B.n208 163.367
R585 B.n214 B.n213 163.367
R586 B.n218 B.n217 163.367
R587 B.n222 B.n221 163.367
R588 B.n226 B.n225 163.367
R589 B.n230 B.n229 163.367
R590 B.n234 B.n233 163.367
R591 B.n238 B.n237 163.367
R592 B.n242 B.n241 163.367
R593 B.n246 B.n245 163.367
R594 B.n250 B.n249 163.367
R595 B.n254 B.n253 163.367
R596 B.n258 B.n257 163.367
R597 B.n262 B.n261 163.367
R598 B.n266 B.n265 163.367
R599 B.n270 B.n269 163.367
R600 B.n274 B.n273 163.367
R601 B.n278 B.n277 163.367
R602 B.n282 B.n281 163.367
R603 B.n286 B.n285 163.367
R604 B.n290 B.n289 163.367
R605 B.n294 B.n293 163.367
R606 B.n298 B.n297 163.367
R607 B.n302 B.n301 163.367
R608 B.n306 B.n305 163.367
R609 B.n310 B.n309 163.367
R610 B.n314 B.n313 163.367
R611 B.n318 B.n317 163.367
R612 B.n322 B.n321 163.367
R613 B.n775 B.n109 163.367
R614 B.n652 B.n374 163.367
R615 B.n660 B.n374 163.367
R616 B.n660 B.n372 163.367
R617 B.n664 B.n372 163.367
R618 B.n664 B.n366 163.367
R619 B.n672 B.n366 163.367
R620 B.n672 B.n364 163.367
R621 B.n676 B.n364 163.367
R622 B.n676 B.n358 163.367
R623 B.n684 B.n358 163.367
R624 B.n684 B.n356 163.367
R625 B.n688 B.n356 163.367
R626 B.n688 B.n350 163.367
R627 B.n696 B.n350 163.367
R628 B.n696 B.n348 163.367
R629 B.n700 B.n348 163.367
R630 B.n700 B.n342 163.367
R631 B.n708 B.n342 163.367
R632 B.n708 B.n340 163.367
R633 B.n712 B.n340 163.367
R634 B.n712 B.n333 163.367
R635 B.n720 B.n333 163.367
R636 B.n720 B.n331 163.367
R637 B.n725 B.n331 163.367
R638 B.n725 B.n326 163.367
R639 B.n733 B.n326 163.367
R640 B.n734 B.n733 163.367
R641 B.n734 B.n5 163.367
R642 B.n6 B.n5 163.367
R643 B.n7 B.n6 163.367
R644 B.n740 B.n7 163.367
R645 B.n741 B.n740 163.367
R646 B.n741 B.n13 163.367
R647 B.n14 B.n13 163.367
R648 B.n15 B.n14 163.367
R649 B.n746 B.n15 163.367
R650 B.n746 B.n20 163.367
R651 B.n21 B.n20 163.367
R652 B.n22 B.n21 163.367
R653 B.n751 B.n22 163.367
R654 B.n751 B.n27 163.367
R655 B.n28 B.n27 163.367
R656 B.n29 B.n28 163.367
R657 B.n756 B.n29 163.367
R658 B.n756 B.n34 163.367
R659 B.n35 B.n34 163.367
R660 B.n36 B.n35 163.367
R661 B.n761 B.n36 163.367
R662 B.n761 B.n41 163.367
R663 B.n42 B.n41 163.367
R664 B.n43 B.n42 163.367
R665 B.n766 B.n43 163.367
R666 B.n766 B.n48 163.367
R667 B.n49 B.n48 163.367
R668 B.n50 B.n49 163.367
R669 B.n771 B.n50 163.367
R670 B.n771 B.n55 163.367
R671 B.n439 B.n437 163.367
R672 B.n443 B.n437 163.367
R673 B.n447 B.n445 163.367
R674 B.n451 B.n435 163.367
R675 B.n455 B.n453 163.367
R676 B.n459 B.n433 163.367
R677 B.n463 B.n461 163.367
R678 B.n467 B.n431 163.367
R679 B.n471 B.n469 163.367
R680 B.n475 B.n429 163.367
R681 B.n479 B.n477 163.367
R682 B.n483 B.n427 163.367
R683 B.n487 B.n485 163.367
R684 B.n491 B.n425 163.367
R685 B.n495 B.n493 163.367
R686 B.n499 B.n423 163.367
R687 B.n503 B.n501 163.367
R688 B.n507 B.n421 163.367
R689 B.n511 B.n509 163.367
R690 B.n515 B.n419 163.367
R691 B.n519 B.n517 163.367
R692 B.n523 B.n417 163.367
R693 B.n527 B.n525 163.367
R694 B.n531 B.n415 163.367
R695 B.n535 B.n533 163.367
R696 B.n539 B.n410 163.367
R697 B.n543 B.n541 163.367
R698 B.n547 B.n408 163.367
R699 B.n551 B.n549 163.367
R700 B.n556 B.n404 163.367
R701 B.n560 B.n558 163.367
R702 B.n564 B.n402 163.367
R703 B.n568 B.n566 163.367
R704 B.n572 B.n400 163.367
R705 B.n576 B.n574 163.367
R706 B.n580 B.n398 163.367
R707 B.n584 B.n582 163.367
R708 B.n588 B.n396 163.367
R709 B.n592 B.n590 163.367
R710 B.n596 B.n394 163.367
R711 B.n600 B.n598 163.367
R712 B.n604 B.n392 163.367
R713 B.n608 B.n606 163.367
R714 B.n612 B.n390 163.367
R715 B.n616 B.n614 163.367
R716 B.n620 B.n388 163.367
R717 B.n624 B.n622 163.367
R718 B.n628 B.n386 163.367
R719 B.n632 B.n630 163.367
R720 B.n636 B.n384 163.367
R721 B.n640 B.n638 163.367
R722 B.n644 B.n382 163.367
R723 B.n648 B.n646 163.367
R724 B.n654 B.n376 163.367
R725 B.n658 B.n376 163.367
R726 B.n658 B.n370 163.367
R727 B.n666 B.n370 163.367
R728 B.n666 B.n368 163.367
R729 B.n670 B.n368 163.367
R730 B.n670 B.n362 163.367
R731 B.n678 B.n362 163.367
R732 B.n678 B.n360 163.367
R733 B.n682 B.n360 163.367
R734 B.n682 B.n354 163.367
R735 B.n690 B.n354 163.367
R736 B.n690 B.n352 163.367
R737 B.n694 B.n352 163.367
R738 B.n694 B.n346 163.367
R739 B.n702 B.n346 163.367
R740 B.n702 B.n344 163.367
R741 B.n706 B.n344 163.367
R742 B.n706 B.n338 163.367
R743 B.n714 B.n338 163.367
R744 B.n714 B.n336 163.367
R745 B.n718 B.n336 163.367
R746 B.n718 B.n330 163.367
R747 B.n727 B.n330 163.367
R748 B.n727 B.n328 163.367
R749 B.n731 B.n328 163.367
R750 B.n731 B.n3 163.367
R751 B.n835 B.n3 163.367
R752 B.n831 B.n2 163.367
R753 B.n831 B.n830 163.367
R754 B.n830 B.n9 163.367
R755 B.n826 B.n9 163.367
R756 B.n826 B.n11 163.367
R757 B.n822 B.n11 163.367
R758 B.n822 B.n17 163.367
R759 B.n818 B.n17 163.367
R760 B.n818 B.n19 163.367
R761 B.n814 B.n19 163.367
R762 B.n814 B.n24 163.367
R763 B.n810 B.n24 163.367
R764 B.n810 B.n26 163.367
R765 B.n806 B.n26 163.367
R766 B.n806 B.n31 163.367
R767 B.n802 B.n31 163.367
R768 B.n802 B.n33 163.367
R769 B.n798 B.n33 163.367
R770 B.n798 B.n38 163.367
R771 B.n794 B.n38 163.367
R772 B.n794 B.n40 163.367
R773 B.n790 B.n40 163.367
R774 B.n790 B.n45 163.367
R775 B.n786 B.n45 163.367
R776 B.n786 B.n47 163.367
R777 B.n782 B.n47 163.367
R778 B.n782 B.n52 163.367
R779 B.n778 B.n52 163.367
R780 B.n110 B.t8 113.873
R781 B.n405 B.t13 113.873
R782 B.n113 B.t5 113.855
R783 B.n411 B.t16 113.855
R784 B.n56 B.n54 71.676
R785 B.n117 B.n57 71.676
R786 B.n121 B.n58 71.676
R787 B.n125 B.n59 71.676
R788 B.n129 B.n60 71.676
R789 B.n133 B.n61 71.676
R790 B.n137 B.n62 71.676
R791 B.n141 B.n63 71.676
R792 B.n145 B.n64 71.676
R793 B.n149 B.n65 71.676
R794 B.n153 B.n66 71.676
R795 B.n157 B.n67 71.676
R796 B.n161 B.n68 71.676
R797 B.n165 B.n69 71.676
R798 B.n169 B.n70 71.676
R799 B.n173 B.n71 71.676
R800 B.n177 B.n72 71.676
R801 B.n181 B.n73 71.676
R802 B.n185 B.n74 71.676
R803 B.n189 B.n75 71.676
R804 B.n193 B.n76 71.676
R805 B.n197 B.n77 71.676
R806 B.n201 B.n78 71.676
R807 B.n205 B.n79 71.676
R808 B.n209 B.n80 71.676
R809 B.n214 B.n81 71.676
R810 B.n218 B.n82 71.676
R811 B.n222 B.n83 71.676
R812 B.n226 B.n84 71.676
R813 B.n230 B.n85 71.676
R814 B.n234 B.n86 71.676
R815 B.n238 B.n87 71.676
R816 B.n242 B.n88 71.676
R817 B.n246 B.n89 71.676
R818 B.n250 B.n90 71.676
R819 B.n254 B.n91 71.676
R820 B.n258 B.n92 71.676
R821 B.n262 B.n93 71.676
R822 B.n266 B.n94 71.676
R823 B.n270 B.n95 71.676
R824 B.n274 B.n96 71.676
R825 B.n278 B.n97 71.676
R826 B.n282 B.n98 71.676
R827 B.n286 B.n99 71.676
R828 B.n290 B.n100 71.676
R829 B.n294 B.n101 71.676
R830 B.n298 B.n102 71.676
R831 B.n302 B.n103 71.676
R832 B.n306 B.n104 71.676
R833 B.n310 B.n105 71.676
R834 B.n314 B.n106 71.676
R835 B.n318 B.n107 71.676
R836 B.n322 B.n108 71.676
R837 B.n109 B.n108 71.676
R838 B.n321 B.n107 71.676
R839 B.n317 B.n106 71.676
R840 B.n313 B.n105 71.676
R841 B.n309 B.n104 71.676
R842 B.n305 B.n103 71.676
R843 B.n301 B.n102 71.676
R844 B.n297 B.n101 71.676
R845 B.n293 B.n100 71.676
R846 B.n289 B.n99 71.676
R847 B.n285 B.n98 71.676
R848 B.n281 B.n97 71.676
R849 B.n277 B.n96 71.676
R850 B.n273 B.n95 71.676
R851 B.n269 B.n94 71.676
R852 B.n265 B.n93 71.676
R853 B.n261 B.n92 71.676
R854 B.n257 B.n91 71.676
R855 B.n253 B.n90 71.676
R856 B.n249 B.n89 71.676
R857 B.n245 B.n88 71.676
R858 B.n241 B.n87 71.676
R859 B.n237 B.n86 71.676
R860 B.n233 B.n85 71.676
R861 B.n229 B.n84 71.676
R862 B.n225 B.n83 71.676
R863 B.n221 B.n82 71.676
R864 B.n217 B.n81 71.676
R865 B.n213 B.n80 71.676
R866 B.n208 B.n79 71.676
R867 B.n204 B.n78 71.676
R868 B.n200 B.n77 71.676
R869 B.n196 B.n76 71.676
R870 B.n192 B.n75 71.676
R871 B.n188 B.n74 71.676
R872 B.n184 B.n73 71.676
R873 B.n180 B.n72 71.676
R874 B.n176 B.n71 71.676
R875 B.n172 B.n70 71.676
R876 B.n168 B.n69 71.676
R877 B.n164 B.n68 71.676
R878 B.n160 B.n67 71.676
R879 B.n156 B.n66 71.676
R880 B.n152 B.n65 71.676
R881 B.n148 B.n64 71.676
R882 B.n144 B.n63 71.676
R883 B.n140 B.n62 71.676
R884 B.n136 B.n61 71.676
R885 B.n132 B.n60 71.676
R886 B.n128 B.n59 71.676
R887 B.n124 B.n58 71.676
R888 B.n120 B.n57 71.676
R889 B.n116 B.n56 71.676
R890 B.n438 B.n378 71.676
R891 B.n444 B.n443 71.676
R892 B.n447 B.n446 71.676
R893 B.n452 B.n451 71.676
R894 B.n455 B.n454 71.676
R895 B.n460 B.n459 71.676
R896 B.n463 B.n462 71.676
R897 B.n468 B.n467 71.676
R898 B.n471 B.n470 71.676
R899 B.n476 B.n475 71.676
R900 B.n479 B.n478 71.676
R901 B.n484 B.n483 71.676
R902 B.n487 B.n486 71.676
R903 B.n492 B.n491 71.676
R904 B.n495 B.n494 71.676
R905 B.n500 B.n499 71.676
R906 B.n503 B.n502 71.676
R907 B.n508 B.n507 71.676
R908 B.n511 B.n510 71.676
R909 B.n516 B.n515 71.676
R910 B.n519 B.n518 71.676
R911 B.n524 B.n523 71.676
R912 B.n527 B.n526 71.676
R913 B.n532 B.n531 71.676
R914 B.n535 B.n534 71.676
R915 B.n540 B.n539 71.676
R916 B.n543 B.n542 71.676
R917 B.n548 B.n547 71.676
R918 B.n551 B.n550 71.676
R919 B.n557 B.n556 71.676
R920 B.n560 B.n559 71.676
R921 B.n565 B.n564 71.676
R922 B.n568 B.n567 71.676
R923 B.n573 B.n572 71.676
R924 B.n576 B.n575 71.676
R925 B.n581 B.n580 71.676
R926 B.n584 B.n583 71.676
R927 B.n589 B.n588 71.676
R928 B.n592 B.n591 71.676
R929 B.n597 B.n596 71.676
R930 B.n600 B.n599 71.676
R931 B.n605 B.n604 71.676
R932 B.n608 B.n607 71.676
R933 B.n613 B.n612 71.676
R934 B.n616 B.n615 71.676
R935 B.n621 B.n620 71.676
R936 B.n624 B.n623 71.676
R937 B.n629 B.n628 71.676
R938 B.n632 B.n631 71.676
R939 B.n637 B.n636 71.676
R940 B.n640 B.n639 71.676
R941 B.n645 B.n644 71.676
R942 B.n648 B.n647 71.676
R943 B.n439 B.n438 71.676
R944 B.n445 B.n444 71.676
R945 B.n446 B.n435 71.676
R946 B.n453 B.n452 71.676
R947 B.n454 B.n433 71.676
R948 B.n461 B.n460 71.676
R949 B.n462 B.n431 71.676
R950 B.n469 B.n468 71.676
R951 B.n470 B.n429 71.676
R952 B.n477 B.n476 71.676
R953 B.n478 B.n427 71.676
R954 B.n485 B.n484 71.676
R955 B.n486 B.n425 71.676
R956 B.n493 B.n492 71.676
R957 B.n494 B.n423 71.676
R958 B.n501 B.n500 71.676
R959 B.n502 B.n421 71.676
R960 B.n509 B.n508 71.676
R961 B.n510 B.n419 71.676
R962 B.n517 B.n516 71.676
R963 B.n518 B.n417 71.676
R964 B.n525 B.n524 71.676
R965 B.n526 B.n415 71.676
R966 B.n533 B.n532 71.676
R967 B.n534 B.n410 71.676
R968 B.n541 B.n540 71.676
R969 B.n542 B.n408 71.676
R970 B.n549 B.n548 71.676
R971 B.n550 B.n404 71.676
R972 B.n558 B.n557 71.676
R973 B.n559 B.n402 71.676
R974 B.n566 B.n565 71.676
R975 B.n567 B.n400 71.676
R976 B.n574 B.n573 71.676
R977 B.n575 B.n398 71.676
R978 B.n582 B.n581 71.676
R979 B.n583 B.n396 71.676
R980 B.n590 B.n589 71.676
R981 B.n591 B.n394 71.676
R982 B.n598 B.n597 71.676
R983 B.n599 B.n392 71.676
R984 B.n606 B.n605 71.676
R985 B.n607 B.n390 71.676
R986 B.n614 B.n613 71.676
R987 B.n615 B.n388 71.676
R988 B.n622 B.n621 71.676
R989 B.n623 B.n386 71.676
R990 B.n630 B.n629 71.676
R991 B.n631 B.n384 71.676
R992 B.n638 B.n637 71.676
R993 B.n639 B.n382 71.676
R994 B.n646 B.n645 71.676
R995 B.n647 B.n380 71.676
R996 B.n836 B.n835 71.676
R997 B.n836 B.n2 71.676
R998 B.n111 B.t9 69.2667
R999 B.n406 B.t12 69.2667
R1000 B.n114 B.t6 69.248
R1001 B.n412 B.t15 69.248
R1002 B.n653 B.n379 65.5133
R1003 B.n777 B.n776 65.5133
R1004 B.n211 B.n114 59.5399
R1005 B.n112 B.n111 59.5399
R1006 B.n553 B.n406 59.5399
R1007 B.n413 B.n412 59.5399
R1008 B.n114 B.n113 44.6066
R1009 B.n111 B.n110 44.6066
R1010 B.n406 B.n405 44.6066
R1011 B.n412 B.n411 44.6066
R1012 B.n653 B.n375 38.0763
R1013 B.n659 B.n375 38.0763
R1014 B.n659 B.n371 38.0763
R1015 B.n665 B.n371 38.0763
R1016 B.n665 B.n367 38.0763
R1017 B.n671 B.n367 38.0763
R1018 B.n677 B.n363 38.0763
R1019 B.n677 B.n359 38.0763
R1020 B.n683 B.n359 38.0763
R1021 B.n683 B.n355 38.0763
R1022 B.n689 B.n355 38.0763
R1023 B.n689 B.n351 38.0763
R1024 B.n695 B.n351 38.0763
R1025 B.n695 B.n347 38.0763
R1026 B.n701 B.n347 38.0763
R1027 B.n707 B.n343 38.0763
R1028 B.n707 B.n339 38.0763
R1029 B.n713 B.n339 38.0763
R1030 B.n713 B.n334 38.0763
R1031 B.n719 B.n334 38.0763
R1032 B.n719 B.n335 38.0763
R1033 B.n726 B.n327 38.0763
R1034 B.n732 B.n327 38.0763
R1035 B.n732 B.n4 38.0763
R1036 B.n834 B.n4 38.0763
R1037 B.n834 B.n833 38.0763
R1038 B.n833 B.n832 38.0763
R1039 B.n832 B.n8 38.0763
R1040 B.n12 B.n8 38.0763
R1041 B.n825 B.n12 38.0763
R1042 B.n824 B.n823 38.0763
R1043 B.n823 B.n16 38.0763
R1044 B.n817 B.n16 38.0763
R1045 B.n817 B.n816 38.0763
R1046 B.n816 B.n815 38.0763
R1047 B.n815 B.n23 38.0763
R1048 B.n809 B.n808 38.0763
R1049 B.n808 B.n807 38.0763
R1050 B.n807 B.n30 38.0763
R1051 B.n801 B.n30 38.0763
R1052 B.n801 B.n800 38.0763
R1053 B.n800 B.n799 38.0763
R1054 B.n799 B.n37 38.0763
R1055 B.n793 B.n37 38.0763
R1056 B.n793 B.n792 38.0763
R1057 B.n791 B.n44 38.0763
R1058 B.n785 B.n44 38.0763
R1059 B.n785 B.n784 38.0763
R1060 B.n784 B.n783 38.0763
R1061 B.n783 B.n51 38.0763
R1062 B.n777 B.n51 38.0763
R1063 B.n655 B.n377 30.1273
R1064 B.n651 B.n650 30.1273
R1065 B.n774 B.n773 30.1273
R1066 B.n779 B.n53 30.1273
R1067 B.n671 B.t11 29.6773
R1068 B.t4 B.n791 29.6773
R1069 B.n701 B.t17 28.5574
R1070 B.n809 B.t0 28.5574
R1071 B.n335 B.t2 19.5984
R1072 B.t1 B.n824 19.5984
R1073 B.n726 B.t2 18.4785
R1074 B.n825 B.t1 18.4785
R1075 B B.n837 18.0485
R1076 B.n656 B.n655 10.6151
R1077 B.n657 B.n656 10.6151
R1078 B.n657 B.n369 10.6151
R1079 B.n667 B.n369 10.6151
R1080 B.n668 B.n667 10.6151
R1081 B.n669 B.n668 10.6151
R1082 B.n669 B.n361 10.6151
R1083 B.n679 B.n361 10.6151
R1084 B.n680 B.n679 10.6151
R1085 B.n681 B.n680 10.6151
R1086 B.n681 B.n353 10.6151
R1087 B.n691 B.n353 10.6151
R1088 B.n692 B.n691 10.6151
R1089 B.n693 B.n692 10.6151
R1090 B.n693 B.n345 10.6151
R1091 B.n703 B.n345 10.6151
R1092 B.n704 B.n703 10.6151
R1093 B.n705 B.n704 10.6151
R1094 B.n705 B.n337 10.6151
R1095 B.n715 B.n337 10.6151
R1096 B.n716 B.n715 10.6151
R1097 B.n717 B.n716 10.6151
R1098 B.n717 B.n329 10.6151
R1099 B.n728 B.n329 10.6151
R1100 B.n729 B.n728 10.6151
R1101 B.n730 B.n729 10.6151
R1102 B.n730 B.n0 10.6151
R1103 B.n440 B.n377 10.6151
R1104 B.n441 B.n440 10.6151
R1105 B.n442 B.n441 10.6151
R1106 B.n442 B.n436 10.6151
R1107 B.n448 B.n436 10.6151
R1108 B.n449 B.n448 10.6151
R1109 B.n450 B.n449 10.6151
R1110 B.n450 B.n434 10.6151
R1111 B.n456 B.n434 10.6151
R1112 B.n457 B.n456 10.6151
R1113 B.n458 B.n457 10.6151
R1114 B.n458 B.n432 10.6151
R1115 B.n464 B.n432 10.6151
R1116 B.n465 B.n464 10.6151
R1117 B.n466 B.n465 10.6151
R1118 B.n466 B.n430 10.6151
R1119 B.n472 B.n430 10.6151
R1120 B.n473 B.n472 10.6151
R1121 B.n474 B.n473 10.6151
R1122 B.n474 B.n428 10.6151
R1123 B.n480 B.n428 10.6151
R1124 B.n481 B.n480 10.6151
R1125 B.n482 B.n481 10.6151
R1126 B.n482 B.n426 10.6151
R1127 B.n488 B.n426 10.6151
R1128 B.n489 B.n488 10.6151
R1129 B.n490 B.n489 10.6151
R1130 B.n490 B.n424 10.6151
R1131 B.n496 B.n424 10.6151
R1132 B.n497 B.n496 10.6151
R1133 B.n498 B.n497 10.6151
R1134 B.n498 B.n422 10.6151
R1135 B.n504 B.n422 10.6151
R1136 B.n505 B.n504 10.6151
R1137 B.n506 B.n505 10.6151
R1138 B.n506 B.n420 10.6151
R1139 B.n512 B.n420 10.6151
R1140 B.n513 B.n512 10.6151
R1141 B.n514 B.n513 10.6151
R1142 B.n514 B.n418 10.6151
R1143 B.n520 B.n418 10.6151
R1144 B.n521 B.n520 10.6151
R1145 B.n522 B.n521 10.6151
R1146 B.n522 B.n416 10.6151
R1147 B.n528 B.n416 10.6151
R1148 B.n529 B.n528 10.6151
R1149 B.n530 B.n529 10.6151
R1150 B.n530 B.n414 10.6151
R1151 B.n537 B.n536 10.6151
R1152 B.n538 B.n537 10.6151
R1153 B.n538 B.n409 10.6151
R1154 B.n544 B.n409 10.6151
R1155 B.n545 B.n544 10.6151
R1156 B.n546 B.n545 10.6151
R1157 B.n546 B.n407 10.6151
R1158 B.n552 B.n407 10.6151
R1159 B.n555 B.n554 10.6151
R1160 B.n555 B.n403 10.6151
R1161 B.n561 B.n403 10.6151
R1162 B.n562 B.n561 10.6151
R1163 B.n563 B.n562 10.6151
R1164 B.n563 B.n401 10.6151
R1165 B.n569 B.n401 10.6151
R1166 B.n570 B.n569 10.6151
R1167 B.n571 B.n570 10.6151
R1168 B.n571 B.n399 10.6151
R1169 B.n577 B.n399 10.6151
R1170 B.n578 B.n577 10.6151
R1171 B.n579 B.n578 10.6151
R1172 B.n579 B.n397 10.6151
R1173 B.n585 B.n397 10.6151
R1174 B.n586 B.n585 10.6151
R1175 B.n587 B.n586 10.6151
R1176 B.n587 B.n395 10.6151
R1177 B.n593 B.n395 10.6151
R1178 B.n594 B.n593 10.6151
R1179 B.n595 B.n594 10.6151
R1180 B.n595 B.n393 10.6151
R1181 B.n601 B.n393 10.6151
R1182 B.n602 B.n601 10.6151
R1183 B.n603 B.n602 10.6151
R1184 B.n603 B.n391 10.6151
R1185 B.n609 B.n391 10.6151
R1186 B.n610 B.n609 10.6151
R1187 B.n611 B.n610 10.6151
R1188 B.n611 B.n389 10.6151
R1189 B.n617 B.n389 10.6151
R1190 B.n618 B.n617 10.6151
R1191 B.n619 B.n618 10.6151
R1192 B.n619 B.n387 10.6151
R1193 B.n625 B.n387 10.6151
R1194 B.n626 B.n625 10.6151
R1195 B.n627 B.n626 10.6151
R1196 B.n627 B.n385 10.6151
R1197 B.n633 B.n385 10.6151
R1198 B.n634 B.n633 10.6151
R1199 B.n635 B.n634 10.6151
R1200 B.n635 B.n383 10.6151
R1201 B.n641 B.n383 10.6151
R1202 B.n642 B.n641 10.6151
R1203 B.n643 B.n642 10.6151
R1204 B.n643 B.n381 10.6151
R1205 B.n649 B.n381 10.6151
R1206 B.n650 B.n649 10.6151
R1207 B.n651 B.n373 10.6151
R1208 B.n661 B.n373 10.6151
R1209 B.n662 B.n661 10.6151
R1210 B.n663 B.n662 10.6151
R1211 B.n663 B.n365 10.6151
R1212 B.n673 B.n365 10.6151
R1213 B.n674 B.n673 10.6151
R1214 B.n675 B.n674 10.6151
R1215 B.n675 B.n357 10.6151
R1216 B.n685 B.n357 10.6151
R1217 B.n686 B.n685 10.6151
R1218 B.n687 B.n686 10.6151
R1219 B.n687 B.n349 10.6151
R1220 B.n697 B.n349 10.6151
R1221 B.n698 B.n697 10.6151
R1222 B.n699 B.n698 10.6151
R1223 B.n699 B.n341 10.6151
R1224 B.n709 B.n341 10.6151
R1225 B.n710 B.n709 10.6151
R1226 B.n711 B.n710 10.6151
R1227 B.n711 B.n332 10.6151
R1228 B.n721 B.n332 10.6151
R1229 B.n722 B.n721 10.6151
R1230 B.n724 B.n722 10.6151
R1231 B.n724 B.n723 10.6151
R1232 B.n723 B.n325 10.6151
R1233 B.n735 B.n325 10.6151
R1234 B.n736 B.n735 10.6151
R1235 B.n737 B.n736 10.6151
R1236 B.n738 B.n737 10.6151
R1237 B.n739 B.n738 10.6151
R1238 B.n742 B.n739 10.6151
R1239 B.n743 B.n742 10.6151
R1240 B.n744 B.n743 10.6151
R1241 B.n745 B.n744 10.6151
R1242 B.n747 B.n745 10.6151
R1243 B.n748 B.n747 10.6151
R1244 B.n749 B.n748 10.6151
R1245 B.n750 B.n749 10.6151
R1246 B.n752 B.n750 10.6151
R1247 B.n753 B.n752 10.6151
R1248 B.n754 B.n753 10.6151
R1249 B.n755 B.n754 10.6151
R1250 B.n757 B.n755 10.6151
R1251 B.n758 B.n757 10.6151
R1252 B.n759 B.n758 10.6151
R1253 B.n760 B.n759 10.6151
R1254 B.n762 B.n760 10.6151
R1255 B.n763 B.n762 10.6151
R1256 B.n764 B.n763 10.6151
R1257 B.n765 B.n764 10.6151
R1258 B.n767 B.n765 10.6151
R1259 B.n768 B.n767 10.6151
R1260 B.n769 B.n768 10.6151
R1261 B.n770 B.n769 10.6151
R1262 B.n772 B.n770 10.6151
R1263 B.n773 B.n772 10.6151
R1264 B.n829 B.n1 10.6151
R1265 B.n829 B.n828 10.6151
R1266 B.n828 B.n827 10.6151
R1267 B.n827 B.n10 10.6151
R1268 B.n821 B.n10 10.6151
R1269 B.n821 B.n820 10.6151
R1270 B.n820 B.n819 10.6151
R1271 B.n819 B.n18 10.6151
R1272 B.n813 B.n18 10.6151
R1273 B.n813 B.n812 10.6151
R1274 B.n812 B.n811 10.6151
R1275 B.n811 B.n25 10.6151
R1276 B.n805 B.n25 10.6151
R1277 B.n805 B.n804 10.6151
R1278 B.n804 B.n803 10.6151
R1279 B.n803 B.n32 10.6151
R1280 B.n797 B.n32 10.6151
R1281 B.n797 B.n796 10.6151
R1282 B.n796 B.n795 10.6151
R1283 B.n795 B.n39 10.6151
R1284 B.n789 B.n39 10.6151
R1285 B.n789 B.n788 10.6151
R1286 B.n788 B.n787 10.6151
R1287 B.n787 B.n46 10.6151
R1288 B.n781 B.n46 10.6151
R1289 B.n781 B.n780 10.6151
R1290 B.n780 B.n779 10.6151
R1291 B.n115 B.n53 10.6151
R1292 B.n118 B.n115 10.6151
R1293 B.n119 B.n118 10.6151
R1294 B.n122 B.n119 10.6151
R1295 B.n123 B.n122 10.6151
R1296 B.n126 B.n123 10.6151
R1297 B.n127 B.n126 10.6151
R1298 B.n130 B.n127 10.6151
R1299 B.n131 B.n130 10.6151
R1300 B.n134 B.n131 10.6151
R1301 B.n135 B.n134 10.6151
R1302 B.n138 B.n135 10.6151
R1303 B.n139 B.n138 10.6151
R1304 B.n142 B.n139 10.6151
R1305 B.n143 B.n142 10.6151
R1306 B.n146 B.n143 10.6151
R1307 B.n147 B.n146 10.6151
R1308 B.n150 B.n147 10.6151
R1309 B.n151 B.n150 10.6151
R1310 B.n154 B.n151 10.6151
R1311 B.n155 B.n154 10.6151
R1312 B.n158 B.n155 10.6151
R1313 B.n159 B.n158 10.6151
R1314 B.n162 B.n159 10.6151
R1315 B.n163 B.n162 10.6151
R1316 B.n166 B.n163 10.6151
R1317 B.n167 B.n166 10.6151
R1318 B.n170 B.n167 10.6151
R1319 B.n171 B.n170 10.6151
R1320 B.n174 B.n171 10.6151
R1321 B.n175 B.n174 10.6151
R1322 B.n178 B.n175 10.6151
R1323 B.n179 B.n178 10.6151
R1324 B.n182 B.n179 10.6151
R1325 B.n183 B.n182 10.6151
R1326 B.n186 B.n183 10.6151
R1327 B.n187 B.n186 10.6151
R1328 B.n190 B.n187 10.6151
R1329 B.n191 B.n190 10.6151
R1330 B.n194 B.n191 10.6151
R1331 B.n195 B.n194 10.6151
R1332 B.n198 B.n195 10.6151
R1333 B.n199 B.n198 10.6151
R1334 B.n202 B.n199 10.6151
R1335 B.n203 B.n202 10.6151
R1336 B.n206 B.n203 10.6151
R1337 B.n207 B.n206 10.6151
R1338 B.n210 B.n207 10.6151
R1339 B.n215 B.n212 10.6151
R1340 B.n216 B.n215 10.6151
R1341 B.n219 B.n216 10.6151
R1342 B.n220 B.n219 10.6151
R1343 B.n223 B.n220 10.6151
R1344 B.n224 B.n223 10.6151
R1345 B.n227 B.n224 10.6151
R1346 B.n228 B.n227 10.6151
R1347 B.n232 B.n231 10.6151
R1348 B.n235 B.n232 10.6151
R1349 B.n236 B.n235 10.6151
R1350 B.n239 B.n236 10.6151
R1351 B.n240 B.n239 10.6151
R1352 B.n243 B.n240 10.6151
R1353 B.n244 B.n243 10.6151
R1354 B.n247 B.n244 10.6151
R1355 B.n248 B.n247 10.6151
R1356 B.n251 B.n248 10.6151
R1357 B.n252 B.n251 10.6151
R1358 B.n255 B.n252 10.6151
R1359 B.n256 B.n255 10.6151
R1360 B.n259 B.n256 10.6151
R1361 B.n260 B.n259 10.6151
R1362 B.n263 B.n260 10.6151
R1363 B.n264 B.n263 10.6151
R1364 B.n267 B.n264 10.6151
R1365 B.n268 B.n267 10.6151
R1366 B.n271 B.n268 10.6151
R1367 B.n272 B.n271 10.6151
R1368 B.n275 B.n272 10.6151
R1369 B.n276 B.n275 10.6151
R1370 B.n279 B.n276 10.6151
R1371 B.n280 B.n279 10.6151
R1372 B.n283 B.n280 10.6151
R1373 B.n284 B.n283 10.6151
R1374 B.n287 B.n284 10.6151
R1375 B.n288 B.n287 10.6151
R1376 B.n291 B.n288 10.6151
R1377 B.n292 B.n291 10.6151
R1378 B.n295 B.n292 10.6151
R1379 B.n296 B.n295 10.6151
R1380 B.n299 B.n296 10.6151
R1381 B.n300 B.n299 10.6151
R1382 B.n303 B.n300 10.6151
R1383 B.n304 B.n303 10.6151
R1384 B.n307 B.n304 10.6151
R1385 B.n308 B.n307 10.6151
R1386 B.n311 B.n308 10.6151
R1387 B.n312 B.n311 10.6151
R1388 B.n315 B.n312 10.6151
R1389 B.n316 B.n315 10.6151
R1390 B.n319 B.n316 10.6151
R1391 B.n320 B.n319 10.6151
R1392 B.n323 B.n320 10.6151
R1393 B.n324 B.n323 10.6151
R1394 B.n774 B.n324 10.6151
R1395 B.t17 B.n343 9.51946
R1396 B.t0 B.n23 9.51946
R1397 B.t11 B.n363 8.39958
R1398 B.n792 B.t4 8.39958
R1399 B.n837 B.n0 8.11757
R1400 B.n837 B.n1 8.11757
R1401 B.n536 B.n413 6.5566
R1402 B.n553 B.n552 6.5566
R1403 B.n212 B.n211 6.5566
R1404 B.n228 B.n112 6.5566
R1405 B.n414 B.n413 4.05904
R1406 B.n554 B.n553 4.05904
R1407 B.n211 B.n210 4.05904
R1408 B.n231 B.n112 4.05904
R1409 VN.n0 VN.t3 211.214
R1410 VN.n1 VN.t2 211.214
R1411 VN.n0 VN.t0 210.686
R1412 VN.n1 VN.t1 210.686
R1413 VN VN.n1 53.7892
R1414 VN VN.n0 7.39144
R1415 VTAIL.n5 VTAIL.t1 47.4104
R1416 VTAIL.n4 VTAIL.t6 47.4104
R1417 VTAIL.n3 VTAIL.t5 47.4104
R1418 VTAIL.n7 VTAIL.t7 47.4103
R1419 VTAIL.n0 VTAIL.t4 47.4103
R1420 VTAIL.n1 VTAIL.t0 47.4103
R1421 VTAIL.n2 VTAIL.t3 47.4103
R1422 VTAIL.n6 VTAIL.t2 47.4103
R1423 VTAIL.n7 VTAIL.n6 26.7376
R1424 VTAIL.n3 VTAIL.n2 26.7376
R1425 VTAIL.n4 VTAIL.n3 1.98326
R1426 VTAIL.n6 VTAIL.n5 1.98326
R1427 VTAIL.n2 VTAIL.n1 1.98326
R1428 VTAIL VTAIL.n0 1.05007
R1429 VTAIL VTAIL.n7 0.93369
R1430 VTAIL.n5 VTAIL.n4 0.470328
R1431 VTAIL.n1 VTAIL.n0 0.470328
R1432 VDD2.n2 VDD2.n0 104.763
R1433 VDD2.n2 VDD2.n1 62.7112
R1434 VDD2.n1 VDD2.t2 1.37837
R1435 VDD2.n1 VDD2.t1 1.37837
R1436 VDD2.n0 VDD2.t0 1.37837
R1437 VDD2.n0 VDD2.t3 1.37837
R1438 VDD2 VDD2.n2 0.0586897
R1439 VP.n2 VP.t0 211.214
R1440 VP.n2 VP.t2 210.686
R1441 VP.n4 VP.t1 175.796
R1442 VP.n11 VP.t3 175.796
R1443 VP.n10 VP.n0 161.3
R1444 VP.n9 VP.n8 161.3
R1445 VP.n7 VP.n1 161.3
R1446 VP.n6 VP.n5 161.3
R1447 VP.n4 VP.n3 91.1828
R1448 VP.n12 VP.n11 91.1828
R1449 VP.n9 VP.n1 56.5193
R1450 VP.n3 VP.n2 53.5103
R1451 VP.n5 VP.n1 24.4675
R1452 VP.n10 VP.n9 24.4675
R1453 VP.n5 VP.n4 19.5741
R1454 VP.n11 VP.n10 19.5741
R1455 VP.n6 VP.n3 0.278367
R1456 VP.n12 VP.n0 0.278367
R1457 VP.n7 VP.n6 0.189894
R1458 VP.n8 VP.n7 0.189894
R1459 VP.n8 VP.n0 0.189894
R1460 VP VP.n12 0.153454
R1461 VDD1 VDD1.n1 105.287
R1462 VDD1 VDD1.n0 62.7694
R1463 VDD1.n0 VDD1.t3 1.37837
R1464 VDD1.n0 VDD1.t1 1.37837
R1465 VDD1.n1 VDD1.t2 1.37837
R1466 VDD1.n1 VDD1.t0 1.37837
C0 VDD2 VN 5.3122f
C1 VDD2 VTAIL 6.06604f
C2 VP VDD1 5.51741f
C3 VTAIL VN 5.04137f
C4 VDD2 VDD1 0.876286f
C5 VP VDD2 0.354343f
C6 VDD1 VTAIL 6.01605f
C7 VDD1 VN 0.148556f
C8 VP VN 6.17811f
C9 VP VTAIL 5.05548f
C10 VDD2 B 3.596326f
C11 VDD1 B 7.75201f
C12 VTAIL B 11.112899f
C13 VN B 9.77728f
C14 VP B 7.765774f
C15 VDD1.t3 B 0.302472f
C16 VDD1.t1 B 0.302472f
C17 VDD1.n0 B 2.7309f
C18 VDD1.t2 B 0.302472f
C19 VDD1.t0 B 0.302472f
C20 VDD1.n1 B 3.46886f
C21 VP.n0 B 0.03977f
C22 VP.t3 B 2.33762f
C23 VP.n1 B 0.044035f
C24 VP.t2 B 2.49986f
C25 VP.t0 B 2.50233f
C26 VP.n2 B 3.15829f
C27 VP.n3 B 1.73239f
C28 VP.t1 B 2.33762f
C29 VP.n4 B 0.916168f
C30 VP.n5 B 0.050669f
C31 VP.n6 B 0.03977f
C32 VP.n7 B 0.030165f
C33 VP.n8 B 0.030165f
C34 VP.n9 B 0.044035f
C35 VP.n10 B 0.050669f
C36 VP.n11 B 0.916168f
C37 VP.n12 B 0.036655f
C38 VDD2.t0 B 0.302429f
C39 VDD2.t3 B 0.302429f
C40 VDD2.n0 B 3.44163f
C41 VDD2.t2 B 0.302429f
C42 VDD2.t1 B 0.302429f
C43 VDD2.n1 B 2.73014f
C44 VDD2.n2 B 3.84263f
C45 VTAIL.t4 B 1.9902f
C46 VTAIL.n0 B 0.280896f
C47 VTAIL.t0 B 1.9902f
C48 VTAIL.n1 B 0.32796f
C49 VTAIL.t3 B 1.9902f
C50 VTAIL.n2 B 1.24164f
C51 VTAIL.t5 B 1.99021f
C52 VTAIL.n3 B 1.24163f
C53 VTAIL.t6 B 1.99021f
C54 VTAIL.n4 B 0.327946f
C55 VTAIL.t1 B 1.99021f
C56 VTAIL.n5 B 0.327946f
C57 VTAIL.t2 B 1.9902f
C58 VTAIL.n6 B 1.24164f
C59 VTAIL.t7 B 1.9902f
C60 VTAIL.n7 B 1.18871f
C61 VN.t3 B 2.45146f
C62 VN.t0 B 2.44904f
C63 VN.n0 B 1.67223f
C64 VN.t2 B 2.45146f
C65 VN.t1 B 2.44904f
C66 VN.n1 B 3.10916f
.ends

