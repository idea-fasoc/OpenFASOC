* NGSPICE file created from diff_pair_sample_1157.ext - technology: sky130A

.subckt diff_pair_sample_1157 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=6.8172 pd=35.74 as=6.8172 ps=35.74 w=17.48 l=0.92
X1 B.t15 B.t13 B.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=6.8172 pd=35.74 as=0 ps=0 w=17.48 l=0.92
X2 B.t12 B.t10 B.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=6.8172 pd=35.74 as=0 ps=0 w=17.48 l=0.92
X3 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=6.8172 pd=35.74 as=0 ps=0 w=17.48 l=0.92
X4 VDD1.t1 VP.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=6.8172 pd=35.74 as=6.8172 ps=35.74 w=17.48 l=0.92
X5 VDD1.t0 VP.t1 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=6.8172 pd=35.74 as=6.8172 ps=35.74 w=17.48 l=0.92
X6 VDD2.t0 VN.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=6.8172 pd=35.74 as=6.8172 ps=35.74 w=17.48 l=0.92
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=6.8172 pd=35.74 as=0 ps=0 w=17.48 l=0.92
R0 VN VN.t0 706.648
R1 VN VN.t1 661.951
R2 VTAIL.n386 VTAIL.n294 289.615
R3 VTAIL.n92 VTAIL.n0 289.615
R4 VTAIL.n288 VTAIL.n196 289.615
R5 VTAIL.n190 VTAIL.n98 289.615
R6 VTAIL.n327 VTAIL.n326 185
R7 VTAIL.n329 VTAIL.n328 185
R8 VTAIL.n322 VTAIL.n321 185
R9 VTAIL.n335 VTAIL.n334 185
R10 VTAIL.n337 VTAIL.n336 185
R11 VTAIL.n318 VTAIL.n317 185
R12 VTAIL.n343 VTAIL.n342 185
R13 VTAIL.n345 VTAIL.n344 185
R14 VTAIL.n314 VTAIL.n313 185
R15 VTAIL.n351 VTAIL.n350 185
R16 VTAIL.n353 VTAIL.n352 185
R17 VTAIL.n310 VTAIL.n309 185
R18 VTAIL.n359 VTAIL.n358 185
R19 VTAIL.n361 VTAIL.n360 185
R20 VTAIL.n306 VTAIL.n305 185
R21 VTAIL.n368 VTAIL.n367 185
R22 VTAIL.n369 VTAIL.n304 185
R23 VTAIL.n371 VTAIL.n370 185
R24 VTAIL.n302 VTAIL.n301 185
R25 VTAIL.n377 VTAIL.n376 185
R26 VTAIL.n379 VTAIL.n378 185
R27 VTAIL.n298 VTAIL.n297 185
R28 VTAIL.n385 VTAIL.n384 185
R29 VTAIL.n387 VTAIL.n386 185
R30 VTAIL.n33 VTAIL.n32 185
R31 VTAIL.n35 VTAIL.n34 185
R32 VTAIL.n28 VTAIL.n27 185
R33 VTAIL.n41 VTAIL.n40 185
R34 VTAIL.n43 VTAIL.n42 185
R35 VTAIL.n24 VTAIL.n23 185
R36 VTAIL.n49 VTAIL.n48 185
R37 VTAIL.n51 VTAIL.n50 185
R38 VTAIL.n20 VTAIL.n19 185
R39 VTAIL.n57 VTAIL.n56 185
R40 VTAIL.n59 VTAIL.n58 185
R41 VTAIL.n16 VTAIL.n15 185
R42 VTAIL.n65 VTAIL.n64 185
R43 VTAIL.n67 VTAIL.n66 185
R44 VTAIL.n12 VTAIL.n11 185
R45 VTAIL.n74 VTAIL.n73 185
R46 VTAIL.n75 VTAIL.n10 185
R47 VTAIL.n77 VTAIL.n76 185
R48 VTAIL.n8 VTAIL.n7 185
R49 VTAIL.n83 VTAIL.n82 185
R50 VTAIL.n85 VTAIL.n84 185
R51 VTAIL.n4 VTAIL.n3 185
R52 VTAIL.n91 VTAIL.n90 185
R53 VTAIL.n93 VTAIL.n92 185
R54 VTAIL.n289 VTAIL.n288 185
R55 VTAIL.n287 VTAIL.n286 185
R56 VTAIL.n200 VTAIL.n199 185
R57 VTAIL.n281 VTAIL.n280 185
R58 VTAIL.n279 VTAIL.n278 185
R59 VTAIL.n204 VTAIL.n203 185
R60 VTAIL.n208 VTAIL.n206 185
R61 VTAIL.n273 VTAIL.n272 185
R62 VTAIL.n271 VTAIL.n270 185
R63 VTAIL.n210 VTAIL.n209 185
R64 VTAIL.n265 VTAIL.n264 185
R65 VTAIL.n263 VTAIL.n262 185
R66 VTAIL.n214 VTAIL.n213 185
R67 VTAIL.n257 VTAIL.n256 185
R68 VTAIL.n255 VTAIL.n254 185
R69 VTAIL.n218 VTAIL.n217 185
R70 VTAIL.n249 VTAIL.n248 185
R71 VTAIL.n247 VTAIL.n246 185
R72 VTAIL.n222 VTAIL.n221 185
R73 VTAIL.n241 VTAIL.n240 185
R74 VTAIL.n239 VTAIL.n238 185
R75 VTAIL.n226 VTAIL.n225 185
R76 VTAIL.n233 VTAIL.n232 185
R77 VTAIL.n231 VTAIL.n230 185
R78 VTAIL.n191 VTAIL.n190 185
R79 VTAIL.n189 VTAIL.n188 185
R80 VTAIL.n102 VTAIL.n101 185
R81 VTAIL.n183 VTAIL.n182 185
R82 VTAIL.n181 VTAIL.n180 185
R83 VTAIL.n106 VTAIL.n105 185
R84 VTAIL.n110 VTAIL.n108 185
R85 VTAIL.n175 VTAIL.n174 185
R86 VTAIL.n173 VTAIL.n172 185
R87 VTAIL.n112 VTAIL.n111 185
R88 VTAIL.n167 VTAIL.n166 185
R89 VTAIL.n165 VTAIL.n164 185
R90 VTAIL.n116 VTAIL.n115 185
R91 VTAIL.n159 VTAIL.n158 185
R92 VTAIL.n157 VTAIL.n156 185
R93 VTAIL.n120 VTAIL.n119 185
R94 VTAIL.n151 VTAIL.n150 185
R95 VTAIL.n149 VTAIL.n148 185
R96 VTAIL.n124 VTAIL.n123 185
R97 VTAIL.n143 VTAIL.n142 185
R98 VTAIL.n141 VTAIL.n140 185
R99 VTAIL.n128 VTAIL.n127 185
R100 VTAIL.n135 VTAIL.n134 185
R101 VTAIL.n133 VTAIL.n132 185
R102 VTAIL.n325 VTAIL.t1 147.659
R103 VTAIL.n31 VTAIL.t0 147.659
R104 VTAIL.n229 VTAIL.t3 147.659
R105 VTAIL.n131 VTAIL.t2 147.659
R106 VTAIL.n328 VTAIL.n327 104.615
R107 VTAIL.n328 VTAIL.n321 104.615
R108 VTAIL.n335 VTAIL.n321 104.615
R109 VTAIL.n336 VTAIL.n335 104.615
R110 VTAIL.n336 VTAIL.n317 104.615
R111 VTAIL.n343 VTAIL.n317 104.615
R112 VTAIL.n344 VTAIL.n343 104.615
R113 VTAIL.n344 VTAIL.n313 104.615
R114 VTAIL.n351 VTAIL.n313 104.615
R115 VTAIL.n352 VTAIL.n351 104.615
R116 VTAIL.n352 VTAIL.n309 104.615
R117 VTAIL.n359 VTAIL.n309 104.615
R118 VTAIL.n360 VTAIL.n359 104.615
R119 VTAIL.n360 VTAIL.n305 104.615
R120 VTAIL.n368 VTAIL.n305 104.615
R121 VTAIL.n369 VTAIL.n368 104.615
R122 VTAIL.n370 VTAIL.n369 104.615
R123 VTAIL.n370 VTAIL.n301 104.615
R124 VTAIL.n377 VTAIL.n301 104.615
R125 VTAIL.n378 VTAIL.n377 104.615
R126 VTAIL.n378 VTAIL.n297 104.615
R127 VTAIL.n385 VTAIL.n297 104.615
R128 VTAIL.n386 VTAIL.n385 104.615
R129 VTAIL.n34 VTAIL.n33 104.615
R130 VTAIL.n34 VTAIL.n27 104.615
R131 VTAIL.n41 VTAIL.n27 104.615
R132 VTAIL.n42 VTAIL.n41 104.615
R133 VTAIL.n42 VTAIL.n23 104.615
R134 VTAIL.n49 VTAIL.n23 104.615
R135 VTAIL.n50 VTAIL.n49 104.615
R136 VTAIL.n50 VTAIL.n19 104.615
R137 VTAIL.n57 VTAIL.n19 104.615
R138 VTAIL.n58 VTAIL.n57 104.615
R139 VTAIL.n58 VTAIL.n15 104.615
R140 VTAIL.n65 VTAIL.n15 104.615
R141 VTAIL.n66 VTAIL.n65 104.615
R142 VTAIL.n66 VTAIL.n11 104.615
R143 VTAIL.n74 VTAIL.n11 104.615
R144 VTAIL.n75 VTAIL.n74 104.615
R145 VTAIL.n76 VTAIL.n75 104.615
R146 VTAIL.n76 VTAIL.n7 104.615
R147 VTAIL.n83 VTAIL.n7 104.615
R148 VTAIL.n84 VTAIL.n83 104.615
R149 VTAIL.n84 VTAIL.n3 104.615
R150 VTAIL.n91 VTAIL.n3 104.615
R151 VTAIL.n92 VTAIL.n91 104.615
R152 VTAIL.n288 VTAIL.n287 104.615
R153 VTAIL.n287 VTAIL.n199 104.615
R154 VTAIL.n280 VTAIL.n199 104.615
R155 VTAIL.n280 VTAIL.n279 104.615
R156 VTAIL.n279 VTAIL.n203 104.615
R157 VTAIL.n208 VTAIL.n203 104.615
R158 VTAIL.n272 VTAIL.n208 104.615
R159 VTAIL.n272 VTAIL.n271 104.615
R160 VTAIL.n271 VTAIL.n209 104.615
R161 VTAIL.n264 VTAIL.n209 104.615
R162 VTAIL.n264 VTAIL.n263 104.615
R163 VTAIL.n263 VTAIL.n213 104.615
R164 VTAIL.n256 VTAIL.n213 104.615
R165 VTAIL.n256 VTAIL.n255 104.615
R166 VTAIL.n255 VTAIL.n217 104.615
R167 VTAIL.n248 VTAIL.n217 104.615
R168 VTAIL.n248 VTAIL.n247 104.615
R169 VTAIL.n247 VTAIL.n221 104.615
R170 VTAIL.n240 VTAIL.n221 104.615
R171 VTAIL.n240 VTAIL.n239 104.615
R172 VTAIL.n239 VTAIL.n225 104.615
R173 VTAIL.n232 VTAIL.n225 104.615
R174 VTAIL.n232 VTAIL.n231 104.615
R175 VTAIL.n190 VTAIL.n189 104.615
R176 VTAIL.n189 VTAIL.n101 104.615
R177 VTAIL.n182 VTAIL.n101 104.615
R178 VTAIL.n182 VTAIL.n181 104.615
R179 VTAIL.n181 VTAIL.n105 104.615
R180 VTAIL.n110 VTAIL.n105 104.615
R181 VTAIL.n174 VTAIL.n110 104.615
R182 VTAIL.n174 VTAIL.n173 104.615
R183 VTAIL.n173 VTAIL.n111 104.615
R184 VTAIL.n166 VTAIL.n111 104.615
R185 VTAIL.n166 VTAIL.n165 104.615
R186 VTAIL.n165 VTAIL.n115 104.615
R187 VTAIL.n158 VTAIL.n115 104.615
R188 VTAIL.n158 VTAIL.n157 104.615
R189 VTAIL.n157 VTAIL.n119 104.615
R190 VTAIL.n150 VTAIL.n119 104.615
R191 VTAIL.n150 VTAIL.n149 104.615
R192 VTAIL.n149 VTAIL.n123 104.615
R193 VTAIL.n142 VTAIL.n123 104.615
R194 VTAIL.n142 VTAIL.n141 104.615
R195 VTAIL.n141 VTAIL.n127 104.615
R196 VTAIL.n134 VTAIL.n127 104.615
R197 VTAIL.n134 VTAIL.n133 104.615
R198 VTAIL.n327 VTAIL.t1 52.3082
R199 VTAIL.n33 VTAIL.t0 52.3082
R200 VTAIL.n231 VTAIL.t3 52.3082
R201 VTAIL.n133 VTAIL.t2 52.3082
R202 VTAIL.n391 VTAIL.n390 31.4096
R203 VTAIL.n97 VTAIL.n96 31.4096
R204 VTAIL.n293 VTAIL.n292 31.4096
R205 VTAIL.n195 VTAIL.n194 31.4096
R206 VTAIL.n195 VTAIL.n97 29.6083
R207 VTAIL.n391 VTAIL.n293 28.5307
R208 VTAIL.n326 VTAIL.n325 15.6677
R209 VTAIL.n32 VTAIL.n31 15.6677
R210 VTAIL.n230 VTAIL.n229 15.6677
R211 VTAIL.n132 VTAIL.n131 15.6677
R212 VTAIL.n371 VTAIL.n302 13.1884
R213 VTAIL.n77 VTAIL.n8 13.1884
R214 VTAIL.n206 VTAIL.n204 13.1884
R215 VTAIL.n108 VTAIL.n106 13.1884
R216 VTAIL.n329 VTAIL.n324 12.8005
R217 VTAIL.n372 VTAIL.n304 12.8005
R218 VTAIL.n376 VTAIL.n375 12.8005
R219 VTAIL.n35 VTAIL.n30 12.8005
R220 VTAIL.n78 VTAIL.n10 12.8005
R221 VTAIL.n82 VTAIL.n81 12.8005
R222 VTAIL.n278 VTAIL.n277 12.8005
R223 VTAIL.n274 VTAIL.n273 12.8005
R224 VTAIL.n233 VTAIL.n228 12.8005
R225 VTAIL.n180 VTAIL.n179 12.8005
R226 VTAIL.n176 VTAIL.n175 12.8005
R227 VTAIL.n135 VTAIL.n130 12.8005
R228 VTAIL.n330 VTAIL.n322 12.0247
R229 VTAIL.n367 VTAIL.n366 12.0247
R230 VTAIL.n379 VTAIL.n300 12.0247
R231 VTAIL.n36 VTAIL.n28 12.0247
R232 VTAIL.n73 VTAIL.n72 12.0247
R233 VTAIL.n85 VTAIL.n6 12.0247
R234 VTAIL.n281 VTAIL.n202 12.0247
R235 VTAIL.n270 VTAIL.n207 12.0247
R236 VTAIL.n234 VTAIL.n226 12.0247
R237 VTAIL.n183 VTAIL.n104 12.0247
R238 VTAIL.n172 VTAIL.n109 12.0247
R239 VTAIL.n136 VTAIL.n128 12.0247
R240 VTAIL.n334 VTAIL.n333 11.249
R241 VTAIL.n365 VTAIL.n306 11.249
R242 VTAIL.n380 VTAIL.n298 11.249
R243 VTAIL.n40 VTAIL.n39 11.249
R244 VTAIL.n71 VTAIL.n12 11.249
R245 VTAIL.n86 VTAIL.n4 11.249
R246 VTAIL.n282 VTAIL.n200 11.249
R247 VTAIL.n269 VTAIL.n210 11.249
R248 VTAIL.n238 VTAIL.n237 11.249
R249 VTAIL.n184 VTAIL.n102 11.249
R250 VTAIL.n171 VTAIL.n112 11.249
R251 VTAIL.n140 VTAIL.n139 11.249
R252 VTAIL.n337 VTAIL.n320 10.4732
R253 VTAIL.n362 VTAIL.n361 10.4732
R254 VTAIL.n384 VTAIL.n383 10.4732
R255 VTAIL.n43 VTAIL.n26 10.4732
R256 VTAIL.n68 VTAIL.n67 10.4732
R257 VTAIL.n90 VTAIL.n89 10.4732
R258 VTAIL.n286 VTAIL.n285 10.4732
R259 VTAIL.n266 VTAIL.n265 10.4732
R260 VTAIL.n241 VTAIL.n224 10.4732
R261 VTAIL.n188 VTAIL.n187 10.4732
R262 VTAIL.n168 VTAIL.n167 10.4732
R263 VTAIL.n143 VTAIL.n126 10.4732
R264 VTAIL.n338 VTAIL.n318 9.69747
R265 VTAIL.n358 VTAIL.n308 9.69747
R266 VTAIL.n387 VTAIL.n296 9.69747
R267 VTAIL.n44 VTAIL.n24 9.69747
R268 VTAIL.n64 VTAIL.n14 9.69747
R269 VTAIL.n93 VTAIL.n2 9.69747
R270 VTAIL.n289 VTAIL.n198 9.69747
R271 VTAIL.n262 VTAIL.n212 9.69747
R272 VTAIL.n242 VTAIL.n222 9.69747
R273 VTAIL.n191 VTAIL.n100 9.69747
R274 VTAIL.n164 VTAIL.n114 9.69747
R275 VTAIL.n144 VTAIL.n124 9.69747
R276 VTAIL.n390 VTAIL.n389 9.45567
R277 VTAIL.n96 VTAIL.n95 9.45567
R278 VTAIL.n292 VTAIL.n291 9.45567
R279 VTAIL.n194 VTAIL.n193 9.45567
R280 VTAIL.n389 VTAIL.n388 9.3005
R281 VTAIL.n296 VTAIL.n295 9.3005
R282 VTAIL.n383 VTAIL.n382 9.3005
R283 VTAIL.n381 VTAIL.n380 9.3005
R284 VTAIL.n300 VTAIL.n299 9.3005
R285 VTAIL.n375 VTAIL.n374 9.3005
R286 VTAIL.n347 VTAIL.n346 9.3005
R287 VTAIL.n316 VTAIL.n315 9.3005
R288 VTAIL.n341 VTAIL.n340 9.3005
R289 VTAIL.n339 VTAIL.n338 9.3005
R290 VTAIL.n320 VTAIL.n319 9.3005
R291 VTAIL.n333 VTAIL.n332 9.3005
R292 VTAIL.n331 VTAIL.n330 9.3005
R293 VTAIL.n324 VTAIL.n323 9.3005
R294 VTAIL.n349 VTAIL.n348 9.3005
R295 VTAIL.n312 VTAIL.n311 9.3005
R296 VTAIL.n355 VTAIL.n354 9.3005
R297 VTAIL.n357 VTAIL.n356 9.3005
R298 VTAIL.n308 VTAIL.n307 9.3005
R299 VTAIL.n363 VTAIL.n362 9.3005
R300 VTAIL.n365 VTAIL.n364 9.3005
R301 VTAIL.n366 VTAIL.n303 9.3005
R302 VTAIL.n373 VTAIL.n372 9.3005
R303 VTAIL.n95 VTAIL.n94 9.3005
R304 VTAIL.n2 VTAIL.n1 9.3005
R305 VTAIL.n89 VTAIL.n88 9.3005
R306 VTAIL.n87 VTAIL.n86 9.3005
R307 VTAIL.n6 VTAIL.n5 9.3005
R308 VTAIL.n81 VTAIL.n80 9.3005
R309 VTAIL.n53 VTAIL.n52 9.3005
R310 VTAIL.n22 VTAIL.n21 9.3005
R311 VTAIL.n47 VTAIL.n46 9.3005
R312 VTAIL.n45 VTAIL.n44 9.3005
R313 VTAIL.n26 VTAIL.n25 9.3005
R314 VTAIL.n39 VTAIL.n38 9.3005
R315 VTAIL.n37 VTAIL.n36 9.3005
R316 VTAIL.n30 VTAIL.n29 9.3005
R317 VTAIL.n55 VTAIL.n54 9.3005
R318 VTAIL.n18 VTAIL.n17 9.3005
R319 VTAIL.n61 VTAIL.n60 9.3005
R320 VTAIL.n63 VTAIL.n62 9.3005
R321 VTAIL.n14 VTAIL.n13 9.3005
R322 VTAIL.n69 VTAIL.n68 9.3005
R323 VTAIL.n71 VTAIL.n70 9.3005
R324 VTAIL.n72 VTAIL.n9 9.3005
R325 VTAIL.n79 VTAIL.n78 9.3005
R326 VTAIL.n216 VTAIL.n215 9.3005
R327 VTAIL.n259 VTAIL.n258 9.3005
R328 VTAIL.n261 VTAIL.n260 9.3005
R329 VTAIL.n212 VTAIL.n211 9.3005
R330 VTAIL.n267 VTAIL.n266 9.3005
R331 VTAIL.n269 VTAIL.n268 9.3005
R332 VTAIL.n207 VTAIL.n205 9.3005
R333 VTAIL.n275 VTAIL.n274 9.3005
R334 VTAIL.n291 VTAIL.n290 9.3005
R335 VTAIL.n198 VTAIL.n197 9.3005
R336 VTAIL.n285 VTAIL.n284 9.3005
R337 VTAIL.n283 VTAIL.n282 9.3005
R338 VTAIL.n202 VTAIL.n201 9.3005
R339 VTAIL.n277 VTAIL.n276 9.3005
R340 VTAIL.n253 VTAIL.n252 9.3005
R341 VTAIL.n251 VTAIL.n250 9.3005
R342 VTAIL.n220 VTAIL.n219 9.3005
R343 VTAIL.n245 VTAIL.n244 9.3005
R344 VTAIL.n243 VTAIL.n242 9.3005
R345 VTAIL.n224 VTAIL.n223 9.3005
R346 VTAIL.n237 VTAIL.n236 9.3005
R347 VTAIL.n235 VTAIL.n234 9.3005
R348 VTAIL.n228 VTAIL.n227 9.3005
R349 VTAIL.n118 VTAIL.n117 9.3005
R350 VTAIL.n161 VTAIL.n160 9.3005
R351 VTAIL.n163 VTAIL.n162 9.3005
R352 VTAIL.n114 VTAIL.n113 9.3005
R353 VTAIL.n169 VTAIL.n168 9.3005
R354 VTAIL.n171 VTAIL.n170 9.3005
R355 VTAIL.n109 VTAIL.n107 9.3005
R356 VTAIL.n177 VTAIL.n176 9.3005
R357 VTAIL.n193 VTAIL.n192 9.3005
R358 VTAIL.n100 VTAIL.n99 9.3005
R359 VTAIL.n187 VTAIL.n186 9.3005
R360 VTAIL.n185 VTAIL.n184 9.3005
R361 VTAIL.n104 VTAIL.n103 9.3005
R362 VTAIL.n179 VTAIL.n178 9.3005
R363 VTAIL.n155 VTAIL.n154 9.3005
R364 VTAIL.n153 VTAIL.n152 9.3005
R365 VTAIL.n122 VTAIL.n121 9.3005
R366 VTAIL.n147 VTAIL.n146 9.3005
R367 VTAIL.n145 VTAIL.n144 9.3005
R368 VTAIL.n126 VTAIL.n125 9.3005
R369 VTAIL.n139 VTAIL.n138 9.3005
R370 VTAIL.n137 VTAIL.n136 9.3005
R371 VTAIL.n130 VTAIL.n129 9.3005
R372 VTAIL.n342 VTAIL.n341 8.92171
R373 VTAIL.n357 VTAIL.n310 8.92171
R374 VTAIL.n388 VTAIL.n294 8.92171
R375 VTAIL.n48 VTAIL.n47 8.92171
R376 VTAIL.n63 VTAIL.n16 8.92171
R377 VTAIL.n94 VTAIL.n0 8.92171
R378 VTAIL.n290 VTAIL.n196 8.92171
R379 VTAIL.n261 VTAIL.n214 8.92171
R380 VTAIL.n246 VTAIL.n245 8.92171
R381 VTAIL.n192 VTAIL.n98 8.92171
R382 VTAIL.n163 VTAIL.n116 8.92171
R383 VTAIL.n148 VTAIL.n147 8.92171
R384 VTAIL.n345 VTAIL.n316 8.14595
R385 VTAIL.n354 VTAIL.n353 8.14595
R386 VTAIL.n51 VTAIL.n22 8.14595
R387 VTAIL.n60 VTAIL.n59 8.14595
R388 VTAIL.n258 VTAIL.n257 8.14595
R389 VTAIL.n249 VTAIL.n220 8.14595
R390 VTAIL.n160 VTAIL.n159 8.14595
R391 VTAIL.n151 VTAIL.n122 8.14595
R392 VTAIL.n346 VTAIL.n314 7.3702
R393 VTAIL.n350 VTAIL.n312 7.3702
R394 VTAIL.n52 VTAIL.n20 7.3702
R395 VTAIL.n56 VTAIL.n18 7.3702
R396 VTAIL.n254 VTAIL.n216 7.3702
R397 VTAIL.n250 VTAIL.n218 7.3702
R398 VTAIL.n156 VTAIL.n118 7.3702
R399 VTAIL.n152 VTAIL.n120 7.3702
R400 VTAIL.n349 VTAIL.n314 6.59444
R401 VTAIL.n350 VTAIL.n349 6.59444
R402 VTAIL.n55 VTAIL.n20 6.59444
R403 VTAIL.n56 VTAIL.n55 6.59444
R404 VTAIL.n254 VTAIL.n253 6.59444
R405 VTAIL.n253 VTAIL.n218 6.59444
R406 VTAIL.n156 VTAIL.n155 6.59444
R407 VTAIL.n155 VTAIL.n120 6.59444
R408 VTAIL.n346 VTAIL.n345 5.81868
R409 VTAIL.n353 VTAIL.n312 5.81868
R410 VTAIL.n52 VTAIL.n51 5.81868
R411 VTAIL.n59 VTAIL.n18 5.81868
R412 VTAIL.n257 VTAIL.n216 5.81868
R413 VTAIL.n250 VTAIL.n249 5.81868
R414 VTAIL.n159 VTAIL.n118 5.81868
R415 VTAIL.n152 VTAIL.n151 5.81868
R416 VTAIL.n342 VTAIL.n316 5.04292
R417 VTAIL.n354 VTAIL.n310 5.04292
R418 VTAIL.n390 VTAIL.n294 5.04292
R419 VTAIL.n48 VTAIL.n22 5.04292
R420 VTAIL.n60 VTAIL.n16 5.04292
R421 VTAIL.n96 VTAIL.n0 5.04292
R422 VTAIL.n292 VTAIL.n196 5.04292
R423 VTAIL.n258 VTAIL.n214 5.04292
R424 VTAIL.n246 VTAIL.n220 5.04292
R425 VTAIL.n194 VTAIL.n98 5.04292
R426 VTAIL.n160 VTAIL.n116 5.04292
R427 VTAIL.n148 VTAIL.n122 5.04292
R428 VTAIL.n325 VTAIL.n323 4.38563
R429 VTAIL.n31 VTAIL.n29 4.38563
R430 VTAIL.n229 VTAIL.n227 4.38563
R431 VTAIL.n131 VTAIL.n129 4.38563
R432 VTAIL.n341 VTAIL.n318 4.26717
R433 VTAIL.n358 VTAIL.n357 4.26717
R434 VTAIL.n388 VTAIL.n387 4.26717
R435 VTAIL.n47 VTAIL.n24 4.26717
R436 VTAIL.n64 VTAIL.n63 4.26717
R437 VTAIL.n94 VTAIL.n93 4.26717
R438 VTAIL.n290 VTAIL.n289 4.26717
R439 VTAIL.n262 VTAIL.n261 4.26717
R440 VTAIL.n245 VTAIL.n222 4.26717
R441 VTAIL.n192 VTAIL.n191 4.26717
R442 VTAIL.n164 VTAIL.n163 4.26717
R443 VTAIL.n147 VTAIL.n124 4.26717
R444 VTAIL.n338 VTAIL.n337 3.49141
R445 VTAIL.n361 VTAIL.n308 3.49141
R446 VTAIL.n384 VTAIL.n296 3.49141
R447 VTAIL.n44 VTAIL.n43 3.49141
R448 VTAIL.n67 VTAIL.n14 3.49141
R449 VTAIL.n90 VTAIL.n2 3.49141
R450 VTAIL.n286 VTAIL.n198 3.49141
R451 VTAIL.n265 VTAIL.n212 3.49141
R452 VTAIL.n242 VTAIL.n241 3.49141
R453 VTAIL.n188 VTAIL.n100 3.49141
R454 VTAIL.n167 VTAIL.n114 3.49141
R455 VTAIL.n144 VTAIL.n143 3.49141
R456 VTAIL.n334 VTAIL.n320 2.71565
R457 VTAIL.n362 VTAIL.n306 2.71565
R458 VTAIL.n383 VTAIL.n298 2.71565
R459 VTAIL.n40 VTAIL.n26 2.71565
R460 VTAIL.n68 VTAIL.n12 2.71565
R461 VTAIL.n89 VTAIL.n4 2.71565
R462 VTAIL.n285 VTAIL.n200 2.71565
R463 VTAIL.n266 VTAIL.n210 2.71565
R464 VTAIL.n238 VTAIL.n224 2.71565
R465 VTAIL.n187 VTAIL.n102 2.71565
R466 VTAIL.n168 VTAIL.n112 2.71565
R467 VTAIL.n140 VTAIL.n126 2.71565
R468 VTAIL.n333 VTAIL.n322 1.93989
R469 VTAIL.n367 VTAIL.n365 1.93989
R470 VTAIL.n380 VTAIL.n379 1.93989
R471 VTAIL.n39 VTAIL.n28 1.93989
R472 VTAIL.n73 VTAIL.n71 1.93989
R473 VTAIL.n86 VTAIL.n85 1.93989
R474 VTAIL.n282 VTAIL.n281 1.93989
R475 VTAIL.n270 VTAIL.n269 1.93989
R476 VTAIL.n237 VTAIL.n226 1.93989
R477 VTAIL.n184 VTAIL.n183 1.93989
R478 VTAIL.n172 VTAIL.n171 1.93989
R479 VTAIL.n139 VTAIL.n128 1.93989
R480 VTAIL.n330 VTAIL.n329 1.16414
R481 VTAIL.n366 VTAIL.n304 1.16414
R482 VTAIL.n376 VTAIL.n300 1.16414
R483 VTAIL.n36 VTAIL.n35 1.16414
R484 VTAIL.n72 VTAIL.n10 1.16414
R485 VTAIL.n82 VTAIL.n6 1.16414
R486 VTAIL.n278 VTAIL.n202 1.16414
R487 VTAIL.n273 VTAIL.n207 1.16414
R488 VTAIL.n234 VTAIL.n233 1.16414
R489 VTAIL.n180 VTAIL.n104 1.16414
R490 VTAIL.n175 VTAIL.n109 1.16414
R491 VTAIL.n136 VTAIL.n135 1.16414
R492 VTAIL.n293 VTAIL.n195 1.00912
R493 VTAIL VTAIL.n97 0.797914
R494 VTAIL.n326 VTAIL.n324 0.388379
R495 VTAIL.n372 VTAIL.n371 0.388379
R496 VTAIL.n375 VTAIL.n302 0.388379
R497 VTAIL.n32 VTAIL.n30 0.388379
R498 VTAIL.n78 VTAIL.n77 0.388379
R499 VTAIL.n81 VTAIL.n8 0.388379
R500 VTAIL.n277 VTAIL.n204 0.388379
R501 VTAIL.n274 VTAIL.n206 0.388379
R502 VTAIL.n230 VTAIL.n228 0.388379
R503 VTAIL.n179 VTAIL.n106 0.388379
R504 VTAIL.n176 VTAIL.n108 0.388379
R505 VTAIL.n132 VTAIL.n130 0.388379
R506 VTAIL VTAIL.n391 0.211707
R507 VTAIL.n331 VTAIL.n323 0.155672
R508 VTAIL.n332 VTAIL.n331 0.155672
R509 VTAIL.n332 VTAIL.n319 0.155672
R510 VTAIL.n339 VTAIL.n319 0.155672
R511 VTAIL.n340 VTAIL.n339 0.155672
R512 VTAIL.n340 VTAIL.n315 0.155672
R513 VTAIL.n347 VTAIL.n315 0.155672
R514 VTAIL.n348 VTAIL.n347 0.155672
R515 VTAIL.n348 VTAIL.n311 0.155672
R516 VTAIL.n355 VTAIL.n311 0.155672
R517 VTAIL.n356 VTAIL.n355 0.155672
R518 VTAIL.n356 VTAIL.n307 0.155672
R519 VTAIL.n363 VTAIL.n307 0.155672
R520 VTAIL.n364 VTAIL.n363 0.155672
R521 VTAIL.n364 VTAIL.n303 0.155672
R522 VTAIL.n373 VTAIL.n303 0.155672
R523 VTAIL.n374 VTAIL.n373 0.155672
R524 VTAIL.n374 VTAIL.n299 0.155672
R525 VTAIL.n381 VTAIL.n299 0.155672
R526 VTAIL.n382 VTAIL.n381 0.155672
R527 VTAIL.n382 VTAIL.n295 0.155672
R528 VTAIL.n389 VTAIL.n295 0.155672
R529 VTAIL.n37 VTAIL.n29 0.155672
R530 VTAIL.n38 VTAIL.n37 0.155672
R531 VTAIL.n38 VTAIL.n25 0.155672
R532 VTAIL.n45 VTAIL.n25 0.155672
R533 VTAIL.n46 VTAIL.n45 0.155672
R534 VTAIL.n46 VTAIL.n21 0.155672
R535 VTAIL.n53 VTAIL.n21 0.155672
R536 VTAIL.n54 VTAIL.n53 0.155672
R537 VTAIL.n54 VTAIL.n17 0.155672
R538 VTAIL.n61 VTAIL.n17 0.155672
R539 VTAIL.n62 VTAIL.n61 0.155672
R540 VTAIL.n62 VTAIL.n13 0.155672
R541 VTAIL.n69 VTAIL.n13 0.155672
R542 VTAIL.n70 VTAIL.n69 0.155672
R543 VTAIL.n70 VTAIL.n9 0.155672
R544 VTAIL.n79 VTAIL.n9 0.155672
R545 VTAIL.n80 VTAIL.n79 0.155672
R546 VTAIL.n80 VTAIL.n5 0.155672
R547 VTAIL.n87 VTAIL.n5 0.155672
R548 VTAIL.n88 VTAIL.n87 0.155672
R549 VTAIL.n88 VTAIL.n1 0.155672
R550 VTAIL.n95 VTAIL.n1 0.155672
R551 VTAIL.n291 VTAIL.n197 0.155672
R552 VTAIL.n284 VTAIL.n197 0.155672
R553 VTAIL.n284 VTAIL.n283 0.155672
R554 VTAIL.n283 VTAIL.n201 0.155672
R555 VTAIL.n276 VTAIL.n201 0.155672
R556 VTAIL.n276 VTAIL.n275 0.155672
R557 VTAIL.n275 VTAIL.n205 0.155672
R558 VTAIL.n268 VTAIL.n205 0.155672
R559 VTAIL.n268 VTAIL.n267 0.155672
R560 VTAIL.n267 VTAIL.n211 0.155672
R561 VTAIL.n260 VTAIL.n211 0.155672
R562 VTAIL.n260 VTAIL.n259 0.155672
R563 VTAIL.n259 VTAIL.n215 0.155672
R564 VTAIL.n252 VTAIL.n215 0.155672
R565 VTAIL.n252 VTAIL.n251 0.155672
R566 VTAIL.n251 VTAIL.n219 0.155672
R567 VTAIL.n244 VTAIL.n219 0.155672
R568 VTAIL.n244 VTAIL.n243 0.155672
R569 VTAIL.n243 VTAIL.n223 0.155672
R570 VTAIL.n236 VTAIL.n223 0.155672
R571 VTAIL.n236 VTAIL.n235 0.155672
R572 VTAIL.n235 VTAIL.n227 0.155672
R573 VTAIL.n193 VTAIL.n99 0.155672
R574 VTAIL.n186 VTAIL.n99 0.155672
R575 VTAIL.n186 VTAIL.n185 0.155672
R576 VTAIL.n185 VTAIL.n103 0.155672
R577 VTAIL.n178 VTAIL.n103 0.155672
R578 VTAIL.n178 VTAIL.n177 0.155672
R579 VTAIL.n177 VTAIL.n107 0.155672
R580 VTAIL.n170 VTAIL.n107 0.155672
R581 VTAIL.n170 VTAIL.n169 0.155672
R582 VTAIL.n169 VTAIL.n113 0.155672
R583 VTAIL.n162 VTAIL.n113 0.155672
R584 VTAIL.n162 VTAIL.n161 0.155672
R585 VTAIL.n161 VTAIL.n117 0.155672
R586 VTAIL.n154 VTAIL.n117 0.155672
R587 VTAIL.n154 VTAIL.n153 0.155672
R588 VTAIL.n153 VTAIL.n121 0.155672
R589 VTAIL.n146 VTAIL.n121 0.155672
R590 VTAIL.n146 VTAIL.n145 0.155672
R591 VTAIL.n145 VTAIL.n125 0.155672
R592 VTAIL.n138 VTAIL.n125 0.155672
R593 VTAIL.n138 VTAIL.n137 0.155672
R594 VTAIL.n137 VTAIL.n129 0.155672
R595 VDD2.n189 VDD2.n97 289.615
R596 VDD2.n92 VDD2.n0 289.615
R597 VDD2.n190 VDD2.n189 185
R598 VDD2.n188 VDD2.n187 185
R599 VDD2.n101 VDD2.n100 185
R600 VDD2.n182 VDD2.n181 185
R601 VDD2.n180 VDD2.n179 185
R602 VDD2.n105 VDD2.n104 185
R603 VDD2.n109 VDD2.n107 185
R604 VDD2.n174 VDD2.n173 185
R605 VDD2.n172 VDD2.n171 185
R606 VDD2.n111 VDD2.n110 185
R607 VDD2.n166 VDD2.n165 185
R608 VDD2.n164 VDD2.n163 185
R609 VDD2.n115 VDD2.n114 185
R610 VDD2.n158 VDD2.n157 185
R611 VDD2.n156 VDD2.n155 185
R612 VDD2.n119 VDD2.n118 185
R613 VDD2.n150 VDD2.n149 185
R614 VDD2.n148 VDD2.n147 185
R615 VDD2.n123 VDD2.n122 185
R616 VDD2.n142 VDD2.n141 185
R617 VDD2.n140 VDD2.n139 185
R618 VDD2.n127 VDD2.n126 185
R619 VDD2.n134 VDD2.n133 185
R620 VDD2.n132 VDD2.n131 185
R621 VDD2.n33 VDD2.n32 185
R622 VDD2.n35 VDD2.n34 185
R623 VDD2.n28 VDD2.n27 185
R624 VDD2.n41 VDD2.n40 185
R625 VDD2.n43 VDD2.n42 185
R626 VDD2.n24 VDD2.n23 185
R627 VDD2.n49 VDD2.n48 185
R628 VDD2.n51 VDD2.n50 185
R629 VDD2.n20 VDD2.n19 185
R630 VDD2.n57 VDD2.n56 185
R631 VDD2.n59 VDD2.n58 185
R632 VDD2.n16 VDD2.n15 185
R633 VDD2.n65 VDD2.n64 185
R634 VDD2.n67 VDD2.n66 185
R635 VDD2.n12 VDD2.n11 185
R636 VDD2.n74 VDD2.n73 185
R637 VDD2.n75 VDD2.n10 185
R638 VDD2.n77 VDD2.n76 185
R639 VDD2.n8 VDD2.n7 185
R640 VDD2.n83 VDD2.n82 185
R641 VDD2.n85 VDD2.n84 185
R642 VDD2.n4 VDD2.n3 185
R643 VDD2.n91 VDD2.n90 185
R644 VDD2.n93 VDD2.n92 185
R645 VDD2.n130 VDD2.t1 147.659
R646 VDD2.n31 VDD2.t0 147.659
R647 VDD2.n189 VDD2.n188 104.615
R648 VDD2.n188 VDD2.n100 104.615
R649 VDD2.n181 VDD2.n100 104.615
R650 VDD2.n181 VDD2.n180 104.615
R651 VDD2.n180 VDD2.n104 104.615
R652 VDD2.n109 VDD2.n104 104.615
R653 VDD2.n173 VDD2.n109 104.615
R654 VDD2.n173 VDD2.n172 104.615
R655 VDD2.n172 VDD2.n110 104.615
R656 VDD2.n165 VDD2.n110 104.615
R657 VDD2.n165 VDD2.n164 104.615
R658 VDD2.n164 VDD2.n114 104.615
R659 VDD2.n157 VDD2.n114 104.615
R660 VDD2.n157 VDD2.n156 104.615
R661 VDD2.n156 VDD2.n118 104.615
R662 VDD2.n149 VDD2.n118 104.615
R663 VDD2.n149 VDD2.n148 104.615
R664 VDD2.n148 VDD2.n122 104.615
R665 VDD2.n141 VDD2.n122 104.615
R666 VDD2.n141 VDD2.n140 104.615
R667 VDD2.n140 VDD2.n126 104.615
R668 VDD2.n133 VDD2.n126 104.615
R669 VDD2.n133 VDD2.n132 104.615
R670 VDD2.n34 VDD2.n33 104.615
R671 VDD2.n34 VDD2.n27 104.615
R672 VDD2.n41 VDD2.n27 104.615
R673 VDD2.n42 VDD2.n41 104.615
R674 VDD2.n42 VDD2.n23 104.615
R675 VDD2.n49 VDD2.n23 104.615
R676 VDD2.n50 VDD2.n49 104.615
R677 VDD2.n50 VDD2.n19 104.615
R678 VDD2.n57 VDD2.n19 104.615
R679 VDD2.n58 VDD2.n57 104.615
R680 VDD2.n58 VDD2.n15 104.615
R681 VDD2.n65 VDD2.n15 104.615
R682 VDD2.n66 VDD2.n65 104.615
R683 VDD2.n66 VDD2.n11 104.615
R684 VDD2.n74 VDD2.n11 104.615
R685 VDD2.n75 VDD2.n74 104.615
R686 VDD2.n76 VDD2.n75 104.615
R687 VDD2.n76 VDD2.n7 104.615
R688 VDD2.n83 VDD2.n7 104.615
R689 VDD2.n84 VDD2.n83 104.615
R690 VDD2.n84 VDD2.n3 104.615
R691 VDD2.n91 VDD2.n3 104.615
R692 VDD2.n92 VDD2.n91 104.615
R693 VDD2.n194 VDD2.n96 88.9892
R694 VDD2.n132 VDD2.t1 52.3082
R695 VDD2.n33 VDD2.t0 52.3082
R696 VDD2.n194 VDD2.n193 48.0884
R697 VDD2.n131 VDD2.n130 15.6677
R698 VDD2.n32 VDD2.n31 15.6677
R699 VDD2.n107 VDD2.n105 13.1884
R700 VDD2.n77 VDD2.n8 13.1884
R701 VDD2.n179 VDD2.n178 12.8005
R702 VDD2.n175 VDD2.n174 12.8005
R703 VDD2.n134 VDD2.n129 12.8005
R704 VDD2.n35 VDD2.n30 12.8005
R705 VDD2.n78 VDD2.n10 12.8005
R706 VDD2.n82 VDD2.n81 12.8005
R707 VDD2.n182 VDD2.n103 12.0247
R708 VDD2.n171 VDD2.n108 12.0247
R709 VDD2.n135 VDD2.n127 12.0247
R710 VDD2.n36 VDD2.n28 12.0247
R711 VDD2.n73 VDD2.n72 12.0247
R712 VDD2.n85 VDD2.n6 12.0247
R713 VDD2.n183 VDD2.n101 11.249
R714 VDD2.n170 VDD2.n111 11.249
R715 VDD2.n139 VDD2.n138 11.249
R716 VDD2.n40 VDD2.n39 11.249
R717 VDD2.n71 VDD2.n12 11.249
R718 VDD2.n86 VDD2.n4 11.249
R719 VDD2.n187 VDD2.n186 10.4732
R720 VDD2.n167 VDD2.n166 10.4732
R721 VDD2.n142 VDD2.n125 10.4732
R722 VDD2.n43 VDD2.n26 10.4732
R723 VDD2.n68 VDD2.n67 10.4732
R724 VDD2.n90 VDD2.n89 10.4732
R725 VDD2.n190 VDD2.n99 9.69747
R726 VDD2.n163 VDD2.n113 9.69747
R727 VDD2.n143 VDD2.n123 9.69747
R728 VDD2.n44 VDD2.n24 9.69747
R729 VDD2.n64 VDD2.n14 9.69747
R730 VDD2.n93 VDD2.n2 9.69747
R731 VDD2.n193 VDD2.n192 9.45567
R732 VDD2.n96 VDD2.n95 9.45567
R733 VDD2.n117 VDD2.n116 9.3005
R734 VDD2.n160 VDD2.n159 9.3005
R735 VDD2.n162 VDD2.n161 9.3005
R736 VDD2.n113 VDD2.n112 9.3005
R737 VDD2.n168 VDD2.n167 9.3005
R738 VDD2.n170 VDD2.n169 9.3005
R739 VDD2.n108 VDD2.n106 9.3005
R740 VDD2.n176 VDD2.n175 9.3005
R741 VDD2.n192 VDD2.n191 9.3005
R742 VDD2.n99 VDD2.n98 9.3005
R743 VDD2.n186 VDD2.n185 9.3005
R744 VDD2.n184 VDD2.n183 9.3005
R745 VDD2.n103 VDD2.n102 9.3005
R746 VDD2.n178 VDD2.n177 9.3005
R747 VDD2.n154 VDD2.n153 9.3005
R748 VDD2.n152 VDD2.n151 9.3005
R749 VDD2.n121 VDD2.n120 9.3005
R750 VDD2.n146 VDD2.n145 9.3005
R751 VDD2.n144 VDD2.n143 9.3005
R752 VDD2.n125 VDD2.n124 9.3005
R753 VDD2.n138 VDD2.n137 9.3005
R754 VDD2.n136 VDD2.n135 9.3005
R755 VDD2.n129 VDD2.n128 9.3005
R756 VDD2.n95 VDD2.n94 9.3005
R757 VDD2.n2 VDD2.n1 9.3005
R758 VDD2.n89 VDD2.n88 9.3005
R759 VDD2.n87 VDD2.n86 9.3005
R760 VDD2.n6 VDD2.n5 9.3005
R761 VDD2.n81 VDD2.n80 9.3005
R762 VDD2.n53 VDD2.n52 9.3005
R763 VDD2.n22 VDD2.n21 9.3005
R764 VDD2.n47 VDD2.n46 9.3005
R765 VDD2.n45 VDD2.n44 9.3005
R766 VDD2.n26 VDD2.n25 9.3005
R767 VDD2.n39 VDD2.n38 9.3005
R768 VDD2.n37 VDD2.n36 9.3005
R769 VDD2.n30 VDD2.n29 9.3005
R770 VDD2.n55 VDD2.n54 9.3005
R771 VDD2.n18 VDD2.n17 9.3005
R772 VDD2.n61 VDD2.n60 9.3005
R773 VDD2.n63 VDD2.n62 9.3005
R774 VDD2.n14 VDD2.n13 9.3005
R775 VDD2.n69 VDD2.n68 9.3005
R776 VDD2.n71 VDD2.n70 9.3005
R777 VDD2.n72 VDD2.n9 9.3005
R778 VDD2.n79 VDD2.n78 9.3005
R779 VDD2.n191 VDD2.n97 8.92171
R780 VDD2.n162 VDD2.n115 8.92171
R781 VDD2.n147 VDD2.n146 8.92171
R782 VDD2.n48 VDD2.n47 8.92171
R783 VDD2.n63 VDD2.n16 8.92171
R784 VDD2.n94 VDD2.n0 8.92171
R785 VDD2.n159 VDD2.n158 8.14595
R786 VDD2.n150 VDD2.n121 8.14595
R787 VDD2.n51 VDD2.n22 8.14595
R788 VDD2.n60 VDD2.n59 8.14595
R789 VDD2.n155 VDD2.n117 7.3702
R790 VDD2.n151 VDD2.n119 7.3702
R791 VDD2.n52 VDD2.n20 7.3702
R792 VDD2.n56 VDD2.n18 7.3702
R793 VDD2.n155 VDD2.n154 6.59444
R794 VDD2.n154 VDD2.n119 6.59444
R795 VDD2.n55 VDD2.n20 6.59444
R796 VDD2.n56 VDD2.n55 6.59444
R797 VDD2.n158 VDD2.n117 5.81868
R798 VDD2.n151 VDD2.n150 5.81868
R799 VDD2.n52 VDD2.n51 5.81868
R800 VDD2.n59 VDD2.n18 5.81868
R801 VDD2.n193 VDD2.n97 5.04292
R802 VDD2.n159 VDD2.n115 5.04292
R803 VDD2.n147 VDD2.n121 5.04292
R804 VDD2.n48 VDD2.n22 5.04292
R805 VDD2.n60 VDD2.n16 5.04292
R806 VDD2.n96 VDD2.n0 5.04292
R807 VDD2.n130 VDD2.n128 4.38563
R808 VDD2.n31 VDD2.n29 4.38563
R809 VDD2.n191 VDD2.n190 4.26717
R810 VDD2.n163 VDD2.n162 4.26717
R811 VDD2.n146 VDD2.n123 4.26717
R812 VDD2.n47 VDD2.n24 4.26717
R813 VDD2.n64 VDD2.n63 4.26717
R814 VDD2.n94 VDD2.n93 4.26717
R815 VDD2.n187 VDD2.n99 3.49141
R816 VDD2.n166 VDD2.n113 3.49141
R817 VDD2.n143 VDD2.n142 3.49141
R818 VDD2.n44 VDD2.n43 3.49141
R819 VDD2.n67 VDD2.n14 3.49141
R820 VDD2.n90 VDD2.n2 3.49141
R821 VDD2.n186 VDD2.n101 2.71565
R822 VDD2.n167 VDD2.n111 2.71565
R823 VDD2.n139 VDD2.n125 2.71565
R824 VDD2.n40 VDD2.n26 2.71565
R825 VDD2.n68 VDD2.n12 2.71565
R826 VDD2.n89 VDD2.n4 2.71565
R827 VDD2.n183 VDD2.n182 1.93989
R828 VDD2.n171 VDD2.n170 1.93989
R829 VDD2.n138 VDD2.n127 1.93989
R830 VDD2.n39 VDD2.n28 1.93989
R831 VDD2.n73 VDD2.n71 1.93989
R832 VDD2.n86 VDD2.n85 1.93989
R833 VDD2.n179 VDD2.n103 1.16414
R834 VDD2.n174 VDD2.n108 1.16414
R835 VDD2.n135 VDD2.n134 1.16414
R836 VDD2.n36 VDD2.n35 1.16414
R837 VDD2.n72 VDD2.n10 1.16414
R838 VDD2.n82 VDD2.n6 1.16414
R839 VDD2.n178 VDD2.n105 0.388379
R840 VDD2.n175 VDD2.n107 0.388379
R841 VDD2.n131 VDD2.n129 0.388379
R842 VDD2.n32 VDD2.n30 0.388379
R843 VDD2.n78 VDD2.n77 0.388379
R844 VDD2.n81 VDD2.n8 0.388379
R845 VDD2 VDD2.n194 0.328086
R846 VDD2.n192 VDD2.n98 0.155672
R847 VDD2.n185 VDD2.n98 0.155672
R848 VDD2.n185 VDD2.n184 0.155672
R849 VDD2.n184 VDD2.n102 0.155672
R850 VDD2.n177 VDD2.n102 0.155672
R851 VDD2.n177 VDD2.n176 0.155672
R852 VDD2.n176 VDD2.n106 0.155672
R853 VDD2.n169 VDD2.n106 0.155672
R854 VDD2.n169 VDD2.n168 0.155672
R855 VDD2.n168 VDD2.n112 0.155672
R856 VDD2.n161 VDD2.n112 0.155672
R857 VDD2.n161 VDD2.n160 0.155672
R858 VDD2.n160 VDD2.n116 0.155672
R859 VDD2.n153 VDD2.n116 0.155672
R860 VDD2.n153 VDD2.n152 0.155672
R861 VDD2.n152 VDD2.n120 0.155672
R862 VDD2.n145 VDD2.n120 0.155672
R863 VDD2.n145 VDD2.n144 0.155672
R864 VDD2.n144 VDD2.n124 0.155672
R865 VDD2.n137 VDD2.n124 0.155672
R866 VDD2.n137 VDD2.n136 0.155672
R867 VDD2.n136 VDD2.n128 0.155672
R868 VDD2.n37 VDD2.n29 0.155672
R869 VDD2.n38 VDD2.n37 0.155672
R870 VDD2.n38 VDD2.n25 0.155672
R871 VDD2.n45 VDD2.n25 0.155672
R872 VDD2.n46 VDD2.n45 0.155672
R873 VDD2.n46 VDD2.n21 0.155672
R874 VDD2.n53 VDD2.n21 0.155672
R875 VDD2.n54 VDD2.n53 0.155672
R876 VDD2.n54 VDD2.n17 0.155672
R877 VDD2.n61 VDD2.n17 0.155672
R878 VDD2.n62 VDD2.n61 0.155672
R879 VDD2.n62 VDD2.n13 0.155672
R880 VDD2.n69 VDD2.n13 0.155672
R881 VDD2.n70 VDD2.n69 0.155672
R882 VDD2.n70 VDD2.n9 0.155672
R883 VDD2.n79 VDD2.n9 0.155672
R884 VDD2.n80 VDD2.n79 0.155672
R885 VDD2.n80 VDD2.n5 0.155672
R886 VDD2.n87 VDD2.n5 0.155672
R887 VDD2.n88 VDD2.n87 0.155672
R888 VDD2.n88 VDD2.n1 0.155672
R889 VDD2.n95 VDD2.n1 0.155672
R890 B.n99 B.t13 660.25
R891 B.n97 B.t6 660.25
R892 B.n439 B.t10 660.25
R893 B.n437 B.t2 660.25
R894 B.n759 B.n758 585
R895 B.n760 B.n759 585
R896 B.n345 B.n95 585
R897 B.n344 B.n343 585
R898 B.n342 B.n341 585
R899 B.n340 B.n339 585
R900 B.n338 B.n337 585
R901 B.n336 B.n335 585
R902 B.n334 B.n333 585
R903 B.n332 B.n331 585
R904 B.n330 B.n329 585
R905 B.n328 B.n327 585
R906 B.n326 B.n325 585
R907 B.n324 B.n323 585
R908 B.n322 B.n321 585
R909 B.n320 B.n319 585
R910 B.n318 B.n317 585
R911 B.n316 B.n315 585
R912 B.n314 B.n313 585
R913 B.n312 B.n311 585
R914 B.n310 B.n309 585
R915 B.n308 B.n307 585
R916 B.n306 B.n305 585
R917 B.n304 B.n303 585
R918 B.n302 B.n301 585
R919 B.n300 B.n299 585
R920 B.n298 B.n297 585
R921 B.n296 B.n295 585
R922 B.n294 B.n293 585
R923 B.n292 B.n291 585
R924 B.n290 B.n289 585
R925 B.n288 B.n287 585
R926 B.n286 B.n285 585
R927 B.n284 B.n283 585
R928 B.n282 B.n281 585
R929 B.n280 B.n279 585
R930 B.n278 B.n277 585
R931 B.n276 B.n275 585
R932 B.n274 B.n273 585
R933 B.n272 B.n271 585
R934 B.n270 B.n269 585
R935 B.n268 B.n267 585
R936 B.n266 B.n265 585
R937 B.n264 B.n263 585
R938 B.n262 B.n261 585
R939 B.n260 B.n259 585
R940 B.n258 B.n257 585
R941 B.n256 B.n255 585
R942 B.n254 B.n253 585
R943 B.n252 B.n251 585
R944 B.n250 B.n249 585
R945 B.n248 B.n247 585
R946 B.n246 B.n245 585
R947 B.n244 B.n243 585
R948 B.n242 B.n241 585
R949 B.n240 B.n239 585
R950 B.n238 B.n237 585
R951 B.n236 B.n235 585
R952 B.n234 B.n233 585
R953 B.n231 B.n230 585
R954 B.n229 B.n228 585
R955 B.n227 B.n226 585
R956 B.n225 B.n224 585
R957 B.n223 B.n222 585
R958 B.n221 B.n220 585
R959 B.n219 B.n218 585
R960 B.n217 B.n216 585
R961 B.n215 B.n214 585
R962 B.n213 B.n212 585
R963 B.n211 B.n210 585
R964 B.n209 B.n208 585
R965 B.n207 B.n206 585
R966 B.n205 B.n204 585
R967 B.n203 B.n202 585
R968 B.n201 B.n200 585
R969 B.n199 B.n198 585
R970 B.n197 B.n196 585
R971 B.n195 B.n194 585
R972 B.n193 B.n192 585
R973 B.n191 B.n190 585
R974 B.n189 B.n188 585
R975 B.n187 B.n186 585
R976 B.n185 B.n184 585
R977 B.n183 B.n182 585
R978 B.n181 B.n180 585
R979 B.n179 B.n178 585
R980 B.n177 B.n176 585
R981 B.n175 B.n174 585
R982 B.n173 B.n172 585
R983 B.n171 B.n170 585
R984 B.n169 B.n168 585
R985 B.n167 B.n166 585
R986 B.n165 B.n164 585
R987 B.n163 B.n162 585
R988 B.n161 B.n160 585
R989 B.n159 B.n158 585
R990 B.n157 B.n156 585
R991 B.n155 B.n154 585
R992 B.n153 B.n152 585
R993 B.n151 B.n150 585
R994 B.n149 B.n148 585
R995 B.n147 B.n146 585
R996 B.n145 B.n144 585
R997 B.n143 B.n142 585
R998 B.n141 B.n140 585
R999 B.n139 B.n138 585
R1000 B.n137 B.n136 585
R1001 B.n135 B.n134 585
R1002 B.n133 B.n132 585
R1003 B.n131 B.n130 585
R1004 B.n129 B.n128 585
R1005 B.n127 B.n126 585
R1006 B.n125 B.n124 585
R1007 B.n123 B.n122 585
R1008 B.n121 B.n120 585
R1009 B.n119 B.n118 585
R1010 B.n117 B.n116 585
R1011 B.n115 B.n114 585
R1012 B.n113 B.n112 585
R1013 B.n111 B.n110 585
R1014 B.n109 B.n108 585
R1015 B.n107 B.n106 585
R1016 B.n105 B.n104 585
R1017 B.n103 B.n102 585
R1018 B.n33 B.n32 585
R1019 B.n763 B.n762 585
R1020 B.n757 B.n96 585
R1021 B.n96 B.n30 585
R1022 B.n756 B.n29 585
R1023 B.n767 B.n29 585
R1024 B.n755 B.n28 585
R1025 B.n768 B.n28 585
R1026 B.n754 B.n27 585
R1027 B.n769 B.n27 585
R1028 B.n753 B.n752 585
R1029 B.n752 B.n23 585
R1030 B.n751 B.n22 585
R1031 B.n775 B.n22 585
R1032 B.n750 B.n21 585
R1033 B.n776 B.n21 585
R1034 B.n749 B.n20 585
R1035 B.n777 B.n20 585
R1036 B.n748 B.n747 585
R1037 B.n747 B.n16 585
R1038 B.n746 B.n15 585
R1039 B.n783 B.n15 585
R1040 B.n745 B.n14 585
R1041 B.n784 B.n14 585
R1042 B.n744 B.n13 585
R1043 B.n785 B.n13 585
R1044 B.n743 B.n742 585
R1045 B.n742 B.n12 585
R1046 B.n741 B.n740 585
R1047 B.n741 B.n8 585
R1048 B.n739 B.n7 585
R1049 B.n792 B.n7 585
R1050 B.n738 B.n6 585
R1051 B.n793 B.n6 585
R1052 B.n737 B.n5 585
R1053 B.n794 B.n5 585
R1054 B.n736 B.n735 585
R1055 B.n735 B.n4 585
R1056 B.n734 B.n346 585
R1057 B.n734 B.n733 585
R1058 B.n723 B.n347 585
R1059 B.n726 B.n347 585
R1060 B.n725 B.n724 585
R1061 B.n727 B.n725 585
R1062 B.n722 B.n352 585
R1063 B.n352 B.n351 585
R1064 B.n721 B.n720 585
R1065 B.n720 B.n719 585
R1066 B.n354 B.n353 585
R1067 B.n355 B.n354 585
R1068 B.n712 B.n711 585
R1069 B.n713 B.n712 585
R1070 B.n710 B.n360 585
R1071 B.n360 B.n359 585
R1072 B.n709 B.n708 585
R1073 B.n708 B.n707 585
R1074 B.n362 B.n361 585
R1075 B.n363 B.n362 585
R1076 B.n700 B.n699 585
R1077 B.n701 B.n700 585
R1078 B.n698 B.n368 585
R1079 B.n368 B.n367 585
R1080 B.n697 B.n696 585
R1081 B.n696 B.n695 585
R1082 B.n370 B.n369 585
R1083 B.n371 B.n370 585
R1084 B.n691 B.n690 585
R1085 B.n374 B.n373 585
R1086 B.n687 B.n686 585
R1087 B.n688 B.n687 585
R1088 B.n685 B.n436 585
R1089 B.n684 B.n683 585
R1090 B.n682 B.n681 585
R1091 B.n680 B.n679 585
R1092 B.n678 B.n677 585
R1093 B.n676 B.n675 585
R1094 B.n674 B.n673 585
R1095 B.n672 B.n671 585
R1096 B.n670 B.n669 585
R1097 B.n668 B.n667 585
R1098 B.n666 B.n665 585
R1099 B.n664 B.n663 585
R1100 B.n662 B.n661 585
R1101 B.n660 B.n659 585
R1102 B.n658 B.n657 585
R1103 B.n656 B.n655 585
R1104 B.n654 B.n653 585
R1105 B.n652 B.n651 585
R1106 B.n650 B.n649 585
R1107 B.n648 B.n647 585
R1108 B.n646 B.n645 585
R1109 B.n644 B.n643 585
R1110 B.n642 B.n641 585
R1111 B.n640 B.n639 585
R1112 B.n638 B.n637 585
R1113 B.n636 B.n635 585
R1114 B.n634 B.n633 585
R1115 B.n632 B.n631 585
R1116 B.n630 B.n629 585
R1117 B.n628 B.n627 585
R1118 B.n626 B.n625 585
R1119 B.n624 B.n623 585
R1120 B.n622 B.n621 585
R1121 B.n620 B.n619 585
R1122 B.n618 B.n617 585
R1123 B.n616 B.n615 585
R1124 B.n614 B.n613 585
R1125 B.n612 B.n611 585
R1126 B.n610 B.n609 585
R1127 B.n608 B.n607 585
R1128 B.n606 B.n605 585
R1129 B.n604 B.n603 585
R1130 B.n602 B.n601 585
R1131 B.n600 B.n599 585
R1132 B.n598 B.n597 585
R1133 B.n596 B.n595 585
R1134 B.n594 B.n593 585
R1135 B.n592 B.n591 585
R1136 B.n590 B.n589 585
R1137 B.n588 B.n587 585
R1138 B.n586 B.n585 585
R1139 B.n584 B.n583 585
R1140 B.n582 B.n581 585
R1141 B.n580 B.n579 585
R1142 B.n578 B.n577 585
R1143 B.n575 B.n574 585
R1144 B.n573 B.n572 585
R1145 B.n571 B.n570 585
R1146 B.n569 B.n568 585
R1147 B.n567 B.n566 585
R1148 B.n565 B.n564 585
R1149 B.n563 B.n562 585
R1150 B.n561 B.n560 585
R1151 B.n559 B.n558 585
R1152 B.n557 B.n556 585
R1153 B.n555 B.n554 585
R1154 B.n553 B.n552 585
R1155 B.n551 B.n550 585
R1156 B.n549 B.n548 585
R1157 B.n547 B.n546 585
R1158 B.n545 B.n544 585
R1159 B.n543 B.n542 585
R1160 B.n541 B.n540 585
R1161 B.n539 B.n538 585
R1162 B.n537 B.n536 585
R1163 B.n535 B.n534 585
R1164 B.n533 B.n532 585
R1165 B.n531 B.n530 585
R1166 B.n529 B.n528 585
R1167 B.n527 B.n526 585
R1168 B.n525 B.n524 585
R1169 B.n523 B.n522 585
R1170 B.n521 B.n520 585
R1171 B.n519 B.n518 585
R1172 B.n517 B.n516 585
R1173 B.n515 B.n514 585
R1174 B.n513 B.n512 585
R1175 B.n511 B.n510 585
R1176 B.n509 B.n508 585
R1177 B.n507 B.n506 585
R1178 B.n505 B.n504 585
R1179 B.n503 B.n502 585
R1180 B.n501 B.n500 585
R1181 B.n499 B.n498 585
R1182 B.n497 B.n496 585
R1183 B.n495 B.n494 585
R1184 B.n493 B.n492 585
R1185 B.n491 B.n490 585
R1186 B.n489 B.n488 585
R1187 B.n487 B.n486 585
R1188 B.n485 B.n484 585
R1189 B.n483 B.n482 585
R1190 B.n481 B.n480 585
R1191 B.n479 B.n478 585
R1192 B.n477 B.n476 585
R1193 B.n475 B.n474 585
R1194 B.n473 B.n472 585
R1195 B.n471 B.n470 585
R1196 B.n469 B.n468 585
R1197 B.n467 B.n466 585
R1198 B.n465 B.n464 585
R1199 B.n463 B.n462 585
R1200 B.n461 B.n460 585
R1201 B.n459 B.n458 585
R1202 B.n457 B.n456 585
R1203 B.n455 B.n454 585
R1204 B.n453 B.n452 585
R1205 B.n451 B.n450 585
R1206 B.n449 B.n448 585
R1207 B.n447 B.n446 585
R1208 B.n445 B.n444 585
R1209 B.n443 B.n442 585
R1210 B.n692 B.n372 585
R1211 B.n372 B.n371 585
R1212 B.n694 B.n693 585
R1213 B.n695 B.n694 585
R1214 B.n366 B.n365 585
R1215 B.n367 B.n366 585
R1216 B.n703 B.n702 585
R1217 B.n702 B.n701 585
R1218 B.n704 B.n364 585
R1219 B.n364 B.n363 585
R1220 B.n706 B.n705 585
R1221 B.n707 B.n706 585
R1222 B.n358 B.n357 585
R1223 B.n359 B.n358 585
R1224 B.n715 B.n714 585
R1225 B.n714 B.n713 585
R1226 B.n716 B.n356 585
R1227 B.n356 B.n355 585
R1228 B.n718 B.n717 585
R1229 B.n719 B.n718 585
R1230 B.n350 B.n349 585
R1231 B.n351 B.n350 585
R1232 B.n729 B.n728 585
R1233 B.n728 B.n727 585
R1234 B.n730 B.n348 585
R1235 B.n726 B.n348 585
R1236 B.n732 B.n731 585
R1237 B.n733 B.n732 585
R1238 B.n3 B.n0 585
R1239 B.n4 B.n3 585
R1240 B.n791 B.n1 585
R1241 B.n792 B.n791 585
R1242 B.n790 B.n789 585
R1243 B.n790 B.n8 585
R1244 B.n788 B.n9 585
R1245 B.n12 B.n9 585
R1246 B.n787 B.n786 585
R1247 B.n786 B.n785 585
R1248 B.n11 B.n10 585
R1249 B.n784 B.n11 585
R1250 B.n782 B.n781 585
R1251 B.n783 B.n782 585
R1252 B.n780 B.n17 585
R1253 B.n17 B.n16 585
R1254 B.n779 B.n778 585
R1255 B.n778 B.n777 585
R1256 B.n19 B.n18 585
R1257 B.n776 B.n19 585
R1258 B.n774 B.n773 585
R1259 B.n775 B.n774 585
R1260 B.n772 B.n24 585
R1261 B.n24 B.n23 585
R1262 B.n771 B.n770 585
R1263 B.n770 B.n769 585
R1264 B.n26 B.n25 585
R1265 B.n768 B.n26 585
R1266 B.n766 B.n765 585
R1267 B.n767 B.n766 585
R1268 B.n764 B.n31 585
R1269 B.n31 B.n30 585
R1270 B.n795 B.n794 585
R1271 B.n793 B.n2 585
R1272 B.n762 B.n31 506.916
R1273 B.n759 B.n96 506.916
R1274 B.n442 B.n370 506.916
R1275 B.n690 B.n372 506.916
R1276 B.n97 B.t8 400.726
R1277 B.n439 B.t12 400.726
R1278 B.n99 B.t14 400.726
R1279 B.n437 B.t5 400.726
R1280 B.n98 B.t9 376.483
R1281 B.n440 B.t11 376.483
R1282 B.n100 B.t15 376.483
R1283 B.n438 B.t4 376.483
R1284 B.n760 B.n94 256.663
R1285 B.n760 B.n93 256.663
R1286 B.n760 B.n92 256.663
R1287 B.n760 B.n91 256.663
R1288 B.n760 B.n90 256.663
R1289 B.n760 B.n89 256.663
R1290 B.n760 B.n88 256.663
R1291 B.n760 B.n87 256.663
R1292 B.n760 B.n86 256.663
R1293 B.n760 B.n85 256.663
R1294 B.n760 B.n84 256.663
R1295 B.n760 B.n83 256.663
R1296 B.n760 B.n82 256.663
R1297 B.n760 B.n81 256.663
R1298 B.n760 B.n80 256.663
R1299 B.n760 B.n79 256.663
R1300 B.n760 B.n78 256.663
R1301 B.n760 B.n77 256.663
R1302 B.n760 B.n76 256.663
R1303 B.n760 B.n75 256.663
R1304 B.n760 B.n74 256.663
R1305 B.n760 B.n73 256.663
R1306 B.n760 B.n72 256.663
R1307 B.n760 B.n71 256.663
R1308 B.n760 B.n70 256.663
R1309 B.n760 B.n69 256.663
R1310 B.n760 B.n68 256.663
R1311 B.n760 B.n67 256.663
R1312 B.n760 B.n66 256.663
R1313 B.n760 B.n65 256.663
R1314 B.n760 B.n64 256.663
R1315 B.n760 B.n63 256.663
R1316 B.n760 B.n62 256.663
R1317 B.n760 B.n61 256.663
R1318 B.n760 B.n60 256.663
R1319 B.n760 B.n59 256.663
R1320 B.n760 B.n58 256.663
R1321 B.n760 B.n57 256.663
R1322 B.n760 B.n56 256.663
R1323 B.n760 B.n55 256.663
R1324 B.n760 B.n54 256.663
R1325 B.n760 B.n53 256.663
R1326 B.n760 B.n52 256.663
R1327 B.n760 B.n51 256.663
R1328 B.n760 B.n50 256.663
R1329 B.n760 B.n49 256.663
R1330 B.n760 B.n48 256.663
R1331 B.n760 B.n47 256.663
R1332 B.n760 B.n46 256.663
R1333 B.n760 B.n45 256.663
R1334 B.n760 B.n44 256.663
R1335 B.n760 B.n43 256.663
R1336 B.n760 B.n42 256.663
R1337 B.n760 B.n41 256.663
R1338 B.n760 B.n40 256.663
R1339 B.n760 B.n39 256.663
R1340 B.n760 B.n38 256.663
R1341 B.n760 B.n37 256.663
R1342 B.n760 B.n36 256.663
R1343 B.n760 B.n35 256.663
R1344 B.n760 B.n34 256.663
R1345 B.n761 B.n760 256.663
R1346 B.n689 B.n688 256.663
R1347 B.n688 B.n375 256.663
R1348 B.n688 B.n376 256.663
R1349 B.n688 B.n377 256.663
R1350 B.n688 B.n378 256.663
R1351 B.n688 B.n379 256.663
R1352 B.n688 B.n380 256.663
R1353 B.n688 B.n381 256.663
R1354 B.n688 B.n382 256.663
R1355 B.n688 B.n383 256.663
R1356 B.n688 B.n384 256.663
R1357 B.n688 B.n385 256.663
R1358 B.n688 B.n386 256.663
R1359 B.n688 B.n387 256.663
R1360 B.n688 B.n388 256.663
R1361 B.n688 B.n389 256.663
R1362 B.n688 B.n390 256.663
R1363 B.n688 B.n391 256.663
R1364 B.n688 B.n392 256.663
R1365 B.n688 B.n393 256.663
R1366 B.n688 B.n394 256.663
R1367 B.n688 B.n395 256.663
R1368 B.n688 B.n396 256.663
R1369 B.n688 B.n397 256.663
R1370 B.n688 B.n398 256.663
R1371 B.n688 B.n399 256.663
R1372 B.n688 B.n400 256.663
R1373 B.n688 B.n401 256.663
R1374 B.n688 B.n402 256.663
R1375 B.n688 B.n403 256.663
R1376 B.n688 B.n404 256.663
R1377 B.n688 B.n405 256.663
R1378 B.n688 B.n406 256.663
R1379 B.n688 B.n407 256.663
R1380 B.n688 B.n408 256.663
R1381 B.n688 B.n409 256.663
R1382 B.n688 B.n410 256.663
R1383 B.n688 B.n411 256.663
R1384 B.n688 B.n412 256.663
R1385 B.n688 B.n413 256.663
R1386 B.n688 B.n414 256.663
R1387 B.n688 B.n415 256.663
R1388 B.n688 B.n416 256.663
R1389 B.n688 B.n417 256.663
R1390 B.n688 B.n418 256.663
R1391 B.n688 B.n419 256.663
R1392 B.n688 B.n420 256.663
R1393 B.n688 B.n421 256.663
R1394 B.n688 B.n422 256.663
R1395 B.n688 B.n423 256.663
R1396 B.n688 B.n424 256.663
R1397 B.n688 B.n425 256.663
R1398 B.n688 B.n426 256.663
R1399 B.n688 B.n427 256.663
R1400 B.n688 B.n428 256.663
R1401 B.n688 B.n429 256.663
R1402 B.n688 B.n430 256.663
R1403 B.n688 B.n431 256.663
R1404 B.n688 B.n432 256.663
R1405 B.n688 B.n433 256.663
R1406 B.n688 B.n434 256.663
R1407 B.n688 B.n435 256.663
R1408 B.n797 B.n796 256.663
R1409 B.n102 B.n33 163.367
R1410 B.n106 B.n105 163.367
R1411 B.n110 B.n109 163.367
R1412 B.n114 B.n113 163.367
R1413 B.n118 B.n117 163.367
R1414 B.n122 B.n121 163.367
R1415 B.n126 B.n125 163.367
R1416 B.n130 B.n129 163.367
R1417 B.n134 B.n133 163.367
R1418 B.n138 B.n137 163.367
R1419 B.n142 B.n141 163.367
R1420 B.n146 B.n145 163.367
R1421 B.n150 B.n149 163.367
R1422 B.n154 B.n153 163.367
R1423 B.n158 B.n157 163.367
R1424 B.n162 B.n161 163.367
R1425 B.n166 B.n165 163.367
R1426 B.n170 B.n169 163.367
R1427 B.n174 B.n173 163.367
R1428 B.n178 B.n177 163.367
R1429 B.n182 B.n181 163.367
R1430 B.n186 B.n185 163.367
R1431 B.n190 B.n189 163.367
R1432 B.n194 B.n193 163.367
R1433 B.n198 B.n197 163.367
R1434 B.n202 B.n201 163.367
R1435 B.n206 B.n205 163.367
R1436 B.n210 B.n209 163.367
R1437 B.n214 B.n213 163.367
R1438 B.n218 B.n217 163.367
R1439 B.n222 B.n221 163.367
R1440 B.n226 B.n225 163.367
R1441 B.n230 B.n229 163.367
R1442 B.n235 B.n234 163.367
R1443 B.n239 B.n238 163.367
R1444 B.n243 B.n242 163.367
R1445 B.n247 B.n246 163.367
R1446 B.n251 B.n250 163.367
R1447 B.n255 B.n254 163.367
R1448 B.n259 B.n258 163.367
R1449 B.n263 B.n262 163.367
R1450 B.n267 B.n266 163.367
R1451 B.n271 B.n270 163.367
R1452 B.n275 B.n274 163.367
R1453 B.n279 B.n278 163.367
R1454 B.n283 B.n282 163.367
R1455 B.n287 B.n286 163.367
R1456 B.n291 B.n290 163.367
R1457 B.n295 B.n294 163.367
R1458 B.n299 B.n298 163.367
R1459 B.n303 B.n302 163.367
R1460 B.n307 B.n306 163.367
R1461 B.n311 B.n310 163.367
R1462 B.n315 B.n314 163.367
R1463 B.n319 B.n318 163.367
R1464 B.n323 B.n322 163.367
R1465 B.n327 B.n326 163.367
R1466 B.n331 B.n330 163.367
R1467 B.n335 B.n334 163.367
R1468 B.n339 B.n338 163.367
R1469 B.n343 B.n342 163.367
R1470 B.n759 B.n95 163.367
R1471 B.n696 B.n370 163.367
R1472 B.n696 B.n368 163.367
R1473 B.n700 B.n368 163.367
R1474 B.n700 B.n362 163.367
R1475 B.n708 B.n362 163.367
R1476 B.n708 B.n360 163.367
R1477 B.n712 B.n360 163.367
R1478 B.n712 B.n354 163.367
R1479 B.n720 B.n354 163.367
R1480 B.n720 B.n352 163.367
R1481 B.n725 B.n352 163.367
R1482 B.n725 B.n347 163.367
R1483 B.n734 B.n347 163.367
R1484 B.n735 B.n734 163.367
R1485 B.n735 B.n5 163.367
R1486 B.n6 B.n5 163.367
R1487 B.n7 B.n6 163.367
R1488 B.n741 B.n7 163.367
R1489 B.n742 B.n741 163.367
R1490 B.n742 B.n13 163.367
R1491 B.n14 B.n13 163.367
R1492 B.n15 B.n14 163.367
R1493 B.n747 B.n15 163.367
R1494 B.n747 B.n20 163.367
R1495 B.n21 B.n20 163.367
R1496 B.n22 B.n21 163.367
R1497 B.n752 B.n22 163.367
R1498 B.n752 B.n27 163.367
R1499 B.n28 B.n27 163.367
R1500 B.n29 B.n28 163.367
R1501 B.n96 B.n29 163.367
R1502 B.n687 B.n374 163.367
R1503 B.n687 B.n436 163.367
R1504 B.n683 B.n682 163.367
R1505 B.n679 B.n678 163.367
R1506 B.n675 B.n674 163.367
R1507 B.n671 B.n670 163.367
R1508 B.n667 B.n666 163.367
R1509 B.n663 B.n662 163.367
R1510 B.n659 B.n658 163.367
R1511 B.n655 B.n654 163.367
R1512 B.n651 B.n650 163.367
R1513 B.n647 B.n646 163.367
R1514 B.n643 B.n642 163.367
R1515 B.n639 B.n638 163.367
R1516 B.n635 B.n634 163.367
R1517 B.n631 B.n630 163.367
R1518 B.n627 B.n626 163.367
R1519 B.n623 B.n622 163.367
R1520 B.n619 B.n618 163.367
R1521 B.n615 B.n614 163.367
R1522 B.n611 B.n610 163.367
R1523 B.n607 B.n606 163.367
R1524 B.n603 B.n602 163.367
R1525 B.n599 B.n598 163.367
R1526 B.n595 B.n594 163.367
R1527 B.n591 B.n590 163.367
R1528 B.n587 B.n586 163.367
R1529 B.n583 B.n582 163.367
R1530 B.n579 B.n578 163.367
R1531 B.n574 B.n573 163.367
R1532 B.n570 B.n569 163.367
R1533 B.n566 B.n565 163.367
R1534 B.n562 B.n561 163.367
R1535 B.n558 B.n557 163.367
R1536 B.n554 B.n553 163.367
R1537 B.n550 B.n549 163.367
R1538 B.n546 B.n545 163.367
R1539 B.n542 B.n541 163.367
R1540 B.n538 B.n537 163.367
R1541 B.n534 B.n533 163.367
R1542 B.n530 B.n529 163.367
R1543 B.n526 B.n525 163.367
R1544 B.n522 B.n521 163.367
R1545 B.n518 B.n517 163.367
R1546 B.n514 B.n513 163.367
R1547 B.n510 B.n509 163.367
R1548 B.n506 B.n505 163.367
R1549 B.n502 B.n501 163.367
R1550 B.n498 B.n497 163.367
R1551 B.n494 B.n493 163.367
R1552 B.n490 B.n489 163.367
R1553 B.n486 B.n485 163.367
R1554 B.n482 B.n481 163.367
R1555 B.n478 B.n477 163.367
R1556 B.n474 B.n473 163.367
R1557 B.n470 B.n469 163.367
R1558 B.n466 B.n465 163.367
R1559 B.n462 B.n461 163.367
R1560 B.n458 B.n457 163.367
R1561 B.n454 B.n453 163.367
R1562 B.n450 B.n449 163.367
R1563 B.n446 B.n445 163.367
R1564 B.n694 B.n372 163.367
R1565 B.n694 B.n366 163.367
R1566 B.n702 B.n366 163.367
R1567 B.n702 B.n364 163.367
R1568 B.n706 B.n364 163.367
R1569 B.n706 B.n358 163.367
R1570 B.n714 B.n358 163.367
R1571 B.n714 B.n356 163.367
R1572 B.n718 B.n356 163.367
R1573 B.n718 B.n350 163.367
R1574 B.n728 B.n350 163.367
R1575 B.n728 B.n348 163.367
R1576 B.n732 B.n348 163.367
R1577 B.n732 B.n3 163.367
R1578 B.n795 B.n3 163.367
R1579 B.n791 B.n2 163.367
R1580 B.n791 B.n790 163.367
R1581 B.n790 B.n9 163.367
R1582 B.n786 B.n9 163.367
R1583 B.n786 B.n11 163.367
R1584 B.n782 B.n11 163.367
R1585 B.n782 B.n17 163.367
R1586 B.n778 B.n17 163.367
R1587 B.n778 B.n19 163.367
R1588 B.n774 B.n19 163.367
R1589 B.n774 B.n24 163.367
R1590 B.n770 B.n24 163.367
R1591 B.n770 B.n26 163.367
R1592 B.n766 B.n26 163.367
R1593 B.n766 B.n31 163.367
R1594 B.n762 B.n761 71.676
R1595 B.n102 B.n34 71.676
R1596 B.n106 B.n35 71.676
R1597 B.n110 B.n36 71.676
R1598 B.n114 B.n37 71.676
R1599 B.n118 B.n38 71.676
R1600 B.n122 B.n39 71.676
R1601 B.n126 B.n40 71.676
R1602 B.n130 B.n41 71.676
R1603 B.n134 B.n42 71.676
R1604 B.n138 B.n43 71.676
R1605 B.n142 B.n44 71.676
R1606 B.n146 B.n45 71.676
R1607 B.n150 B.n46 71.676
R1608 B.n154 B.n47 71.676
R1609 B.n158 B.n48 71.676
R1610 B.n162 B.n49 71.676
R1611 B.n166 B.n50 71.676
R1612 B.n170 B.n51 71.676
R1613 B.n174 B.n52 71.676
R1614 B.n178 B.n53 71.676
R1615 B.n182 B.n54 71.676
R1616 B.n186 B.n55 71.676
R1617 B.n190 B.n56 71.676
R1618 B.n194 B.n57 71.676
R1619 B.n198 B.n58 71.676
R1620 B.n202 B.n59 71.676
R1621 B.n206 B.n60 71.676
R1622 B.n210 B.n61 71.676
R1623 B.n214 B.n62 71.676
R1624 B.n218 B.n63 71.676
R1625 B.n222 B.n64 71.676
R1626 B.n226 B.n65 71.676
R1627 B.n230 B.n66 71.676
R1628 B.n235 B.n67 71.676
R1629 B.n239 B.n68 71.676
R1630 B.n243 B.n69 71.676
R1631 B.n247 B.n70 71.676
R1632 B.n251 B.n71 71.676
R1633 B.n255 B.n72 71.676
R1634 B.n259 B.n73 71.676
R1635 B.n263 B.n74 71.676
R1636 B.n267 B.n75 71.676
R1637 B.n271 B.n76 71.676
R1638 B.n275 B.n77 71.676
R1639 B.n279 B.n78 71.676
R1640 B.n283 B.n79 71.676
R1641 B.n287 B.n80 71.676
R1642 B.n291 B.n81 71.676
R1643 B.n295 B.n82 71.676
R1644 B.n299 B.n83 71.676
R1645 B.n303 B.n84 71.676
R1646 B.n307 B.n85 71.676
R1647 B.n311 B.n86 71.676
R1648 B.n315 B.n87 71.676
R1649 B.n319 B.n88 71.676
R1650 B.n323 B.n89 71.676
R1651 B.n327 B.n90 71.676
R1652 B.n331 B.n91 71.676
R1653 B.n335 B.n92 71.676
R1654 B.n339 B.n93 71.676
R1655 B.n343 B.n94 71.676
R1656 B.n95 B.n94 71.676
R1657 B.n342 B.n93 71.676
R1658 B.n338 B.n92 71.676
R1659 B.n334 B.n91 71.676
R1660 B.n330 B.n90 71.676
R1661 B.n326 B.n89 71.676
R1662 B.n322 B.n88 71.676
R1663 B.n318 B.n87 71.676
R1664 B.n314 B.n86 71.676
R1665 B.n310 B.n85 71.676
R1666 B.n306 B.n84 71.676
R1667 B.n302 B.n83 71.676
R1668 B.n298 B.n82 71.676
R1669 B.n294 B.n81 71.676
R1670 B.n290 B.n80 71.676
R1671 B.n286 B.n79 71.676
R1672 B.n282 B.n78 71.676
R1673 B.n278 B.n77 71.676
R1674 B.n274 B.n76 71.676
R1675 B.n270 B.n75 71.676
R1676 B.n266 B.n74 71.676
R1677 B.n262 B.n73 71.676
R1678 B.n258 B.n72 71.676
R1679 B.n254 B.n71 71.676
R1680 B.n250 B.n70 71.676
R1681 B.n246 B.n69 71.676
R1682 B.n242 B.n68 71.676
R1683 B.n238 B.n67 71.676
R1684 B.n234 B.n66 71.676
R1685 B.n229 B.n65 71.676
R1686 B.n225 B.n64 71.676
R1687 B.n221 B.n63 71.676
R1688 B.n217 B.n62 71.676
R1689 B.n213 B.n61 71.676
R1690 B.n209 B.n60 71.676
R1691 B.n205 B.n59 71.676
R1692 B.n201 B.n58 71.676
R1693 B.n197 B.n57 71.676
R1694 B.n193 B.n56 71.676
R1695 B.n189 B.n55 71.676
R1696 B.n185 B.n54 71.676
R1697 B.n181 B.n53 71.676
R1698 B.n177 B.n52 71.676
R1699 B.n173 B.n51 71.676
R1700 B.n169 B.n50 71.676
R1701 B.n165 B.n49 71.676
R1702 B.n161 B.n48 71.676
R1703 B.n157 B.n47 71.676
R1704 B.n153 B.n46 71.676
R1705 B.n149 B.n45 71.676
R1706 B.n145 B.n44 71.676
R1707 B.n141 B.n43 71.676
R1708 B.n137 B.n42 71.676
R1709 B.n133 B.n41 71.676
R1710 B.n129 B.n40 71.676
R1711 B.n125 B.n39 71.676
R1712 B.n121 B.n38 71.676
R1713 B.n117 B.n37 71.676
R1714 B.n113 B.n36 71.676
R1715 B.n109 B.n35 71.676
R1716 B.n105 B.n34 71.676
R1717 B.n761 B.n33 71.676
R1718 B.n690 B.n689 71.676
R1719 B.n436 B.n375 71.676
R1720 B.n682 B.n376 71.676
R1721 B.n678 B.n377 71.676
R1722 B.n674 B.n378 71.676
R1723 B.n670 B.n379 71.676
R1724 B.n666 B.n380 71.676
R1725 B.n662 B.n381 71.676
R1726 B.n658 B.n382 71.676
R1727 B.n654 B.n383 71.676
R1728 B.n650 B.n384 71.676
R1729 B.n646 B.n385 71.676
R1730 B.n642 B.n386 71.676
R1731 B.n638 B.n387 71.676
R1732 B.n634 B.n388 71.676
R1733 B.n630 B.n389 71.676
R1734 B.n626 B.n390 71.676
R1735 B.n622 B.n391 71.676
R1736 B.n618 B.n392 71.676
R1737 B.n614 B.n393 71.676
R1738 B.n610 B.n394 71.676
R1739 B.n606 B.n395 71.676
R1740 B.n602 B.n396 71.676
R1741 B.n598 B.n397 71.676
R1742 B.n594 B.n398 71.676
R1743 B.n590 B.n399 71.676
R1744 B.n586 B.n400 71.676
R1745 B.n582 B.n401 71.676
R1746 B.n578 B.n402 71.676
R1747 B.n573 B.n403 71.676
R1748 B.n569 B.n404 71.676
R1749 B.n565 B.n405 71.676
R1750 B.n561 B.n406 71.676
R1751 B.n557 B.n407 71.676
R1752 B.n553 B.n408 71.676
R1753 B.n549 B.n409 71.676
R1754 B.n545 B.n410 71.676
R1755 B.n541 B.n411 71.676
R1756 B.n537 B.n412 71.676
R1757 B.n533 B.n413 71.676
R1758 B.n529 B.n414 71.676
R1759 B.n525 B.n415 71.676
R1760 B.n521 B.n416 71.676
R1761 B.n517 B.n417 71.676
R1762 B.n513 B.n418 71.676
R1763 B.n509 B.n419 71.676
R1764 B.n505 B.n420 71.676
R1765 B.n501 B.n421 71.676
R1766 B.n497 B.n422 71.676
R1767 B.n493 B.n423 71.676
R1768 B.n489 B.n424 71.676
R1769 B.n485 B.n425 71.676
R1770 B.n481 B.n426 71.676
R1771 B.n477 B.n427 71.676
R1772 B.n473 B.n428 71.676
R1773 B.n469 B.n429 71.676
R1774 B.n465 B.n430 71.676
R1775 B.n461 B.n431 71.676
R1776 B.n457 B.n432 71.676
R1777 B.n453 B.n433 71.676
R1778 B.n449 B.n434 71.676
R1779 B.n445 B.n435 71.676
R1780 B.n689 B.n374 71.676
R1781 B.n683 B.n375 71.676
R1782 B.n679 B.n376 71.676
R1783 B.n675 B.n377 71.676
R1784 B.n671 B.n378 71.676
R1785 B.n667 B.n379 71.676
R1786 B.n663 B.n380 71.676
R1787 B.n659 B.n381 71.676
R1788 B.n655 B.n382 71.676
R1789 B.n651 B.n383 71.676
R1790 B.n647 B.n384 71.676
R1791 B.n643 B.n385 71.676
R1792 B.n639 B.n386 71.676
R1793 B.n635 B.n387 71.676
R1794 B.n631 B.n388 71.676
R1795 B.n627 B.n389 71.676
R1796 B.n623 B.n390 71.676
R1797 B.n619 B.n391 71.676
R1798 B.n615 B.n392 71.676
R1799 B.n611 B.n393 71.676
R1800 B.n607 B.n394 71.676
R1801 B.n603 B.n395 71.676
R1802 B.n599 B.n396 71.676
R1803 B.n595 B.n397 71.676
R1804 B.n591 B.n398 71.676
R1805 B.n587 B.n399 71.676
R1806 B.n583 B.n400 71.676
R1807 B.n579 B.n401 71.676
R1808 B.n574 B.n402 71.676
R1809 B.n570 B.n403 71.676
R1810 B.n566 B.n404 71.676
R1811 B.n562 B.n405 71.676
R1812 B.n558 B.n406 71.676
R1813 B.n554 B.n407 71.676
R1814 B.n550 B.n408 71.676
R1815 B.n546 B.n409 71.676
R1816 B.n542 B.n410 71.676
R1817 B.n538 B.n411 71.676
R1818 B.n534 B.n412 71.676
R1819 B.n530 B.n413 71.676
R1820 B.n526 B.n414 71.676
R1821 B.n522 B.n415 71.676
R1822 B.n518 B.n416 71.676
R1823 B.n514 B.n417 71.676
R1824 B.n510 B.n418 71.676
R1825 B.n506 B.n419 71.676
R1826 B.n502 B.n420 71.676
R1827 B.n498 B.n421 71.676
R1828 B.n494 B.n422 71.676
R1829 B.n490 B.n423 71.676
R1830 B.n486 B.n424 71.676
R1831 B.n482 B.n425 71.676
R1832 B.n478 B.n426 71.676
R1833 B.n474 B.n427 71.676
R1834 B.n470 B.n428 71.676
R1835 B.n466 B.n429 71.676
R1836 B.n462 B.n430 71.676
R1837 B.n458 B.n431 71.676
R1838 B.n454 B.n432 71.676
R1839 B.n450 B.n433 71.676
R1840 B.n446 B.n434 71.676
R1841 B.n442 B.n435 71.676
R1842 B.n796 B.n795 71.676
R1843 B.n796 B.n2 71.676
R1844 B.n101 B.n100 59.5399
R1845 B.n232 B.n98 59.5399
R1846 B.n441 B.n440 59.5399
R1847 B.n576 B.n438 59.5399
R1848 B.n688 B.n371 58.4418
R1849 B.n760 B.n30 58.4418
R1850 B.n692 B.n691 32.9371
R1851 B.n443 B.n369 32.9371
R1852 B.n758 B.n757 32.9371
R1853 B.n764 B.n763 32.9371
R1854 B.n695 B.n371 32.8435
R1855 B.n695 B.n367 32.8435
R1856 B.n701 B.n367 32.8435
R1857 B.n701 B.n363 32.8435
R1858 B.n707 B.n363 32.8435
R1859 B.n713 B.n359 32.8435
R1860 B.n713 B.n355 32.8435
R1861 B.n719 B.n355 32.8435
R1862 B.n719 B.n351 32.8435
R1863 B.n727 B.n351 32.8435
R1864 B.n727 B.n726 32.8435
R1865 B.n733 B.n4 32.8435
R1866 B.n794 B.n4 32.8435
R1867 B.n794 B.n793 32.8435
R1868 B.n793 B.n792 32.8435
R1869 B.n792 B.n8 32.8435
R1870 B.n785 B.n12 32.8435
R1871 B.n785 B.n784 32.8435
R1872 B.n784 B.n783 32.8435
R1873 B.n783 B.n16 32.8435
R1874 B.n777 B.n16 32.8435
R1875 B.n777 B.n776 32.8435
R1876 B.n775 B.n23 32.8435
R1877 B.n769 B.n23 32.8435
R1878 B.n769 B.n768 32.8435
R1879 B.n768 B.n767 32.8435
R1880 B.n767 B.n30 32.8435
R1881 B.n733 B.t0 30.9116
R1882 B.t1 B.n8 30.9116
R1883 B.t3 B.n359 27.0477
R1884 B.n776 B.t7 27.0477
R1885 B.n100 B.n99 24.2429
R1886 B.n98 B.n97 24.2429
R1887 B.n440 B.n439 24.2429
R1888 B.n438 B.n437 24.2429
R1889 B B.n797 18.0485
R1890 B.n693 B.n692 10.6151
R1891 B.n693 B.n365 10.6151
R1892 B.n703 B.n365 10.6151
R1893 B.n704 B.n703 10.6151
R1894 B.n705 B.n704 10.6151
R1895 B.n705 B.n357 10.6151
R1896 B.n715 B.n357 10.6151
R1897 B.n716 B.n715 10.6151
R1898 B.n717 B.n716 10.6151
R1899 B.n717 B.n349 10.6151
R1900 B.n729 B.n349 10.6151
R1901 B.n730 B.n729 10.6151
R1902 B.n731 B.n730 10.6151
R1903 B.n731 B.n0 10.6151
R1904 B.n691 B.n373 10.6151
R1905 B.n686 B.n373 10.6151
R1906 B.n686 B.n685 10.6151
R1907 B.n685 B.n684 10.6151
R1908 B.n684 B.n681 10.6151
R1909 B.n681 B.n680 10.6151
R1910 B.n680 B.n677 10.6151
R1911 B.n677 B.n676 10.6151
R1912 B.n676 B.n673 10.6151
R1913 B.n673 B.n672 10.6151
R1914 B.n672 B.n669 10.6151
R1915 B.n669 B.n668 10.6151
R1916 B.n668 B.n665 10.6151
R1917 B.n665 B.n664 10.6151
R1918 B.n664 B.n661 10.6151
R1919 B.n661 B.n660 10.6151
R1920 B.n660 B.n657 10.6151
R1921 B.n657 B.n656 10.6151
R1922 B.n656 B.n653 10.6151
R1923 B.n653 B.n652 10.6151
R1924 B.n652 B.n649 10.6151
R1925 B.n649 B.n648 10.6151
R1926 B.n648 B.n645 10.6151
R1927 B.n645 B.n644 10.6151
R1928 B.n644 B.n641 10.6151
R1929 B.n641 B.n640 10.6151
R1930 B.n640 B.n637 10.6151
R1931 B.n637 B.n636 10.6151
R1932 B.n636 B.n633 10.6151
R1933 B.n633 B.n632 10.6151
R1934 B.n632 B.n629 10.6151
R1935 B.n629 B.n628 10.6151
R1936 B.n628 B.n625 10.6151
R1937 B.n625 B.n624 10.6151
R1938 B.n624 B.n621 10.6151
R1939 B.n621 B.n620 10.6151
R1940 B.n620 B.n617 10.6151
R1941 B.n617 B.n616 10.6151
R1942 B.n616 B.n613 10.6151
R1943 B.n613 B.n612 10.6151
R1944 B.n612 B.n609 10.6151
R1945 B.n609 B.n608 10.6151
R1946 B.n608 B.n605 10.6151
R1947 B.n605 B.n604 10.6151
R1948 B.n604 B.n601 10.6151
R1949 B.n601 B.n600 10.6151
R1950 B.n600 B.n597 10.6151
R1951 B.n597 B.n596 10.6151
R1952 B.n596 B.n593 10.6151
R1953 B.n593 B.n592 10.6151
R1954 B.n592 B.n589 10.6151
R1955 B.n589 B.n588 10.6151
R1956 B.n588 B.n585 10.6151
R1957 B.n585 B.n584 10.6151
R1958 B.n584 B.n581 10.6151
R1959 B.n581 B.n580 10.6151
R1960 B.n580 B.n577 10.6151
R1961 B.n575 B.n572 10.6151
R1962 B.n572 B.n571 10.6151
R1963 B.n571 B.n568 10.6151
R1964 B.n568 B.n567 10.6151
R1965 B.n567 B.n564 10.6151
R1966 B.n564 B.n563 10.6151
R1967 B.n563 B.n560 10.6151
R1968 B.n560 B.n559 10.6151
R1969 B.n556 B.n555 10.6151
R1970 B.n555 B.n552 10.6151
R1971 B.n552 B.n551 10.6151
R1972 B.n551 B.n548 10.6151
R1973 B.n548 B.n547 10.6151
R1974 B.n547 B.n544 10.6151
R1975 B.n544 B.n543 10.6151
R1976 B.n543 B.n540 10.6151
R1977 B.n540 B.n539 10.6151
R1978 B.n539 B.n536 10.6151
R1979 B.n536 B.n535 10.6151
R1980 B.n535 B.n532 10.6151
R1981 B.n532 B.n531 10.6151
R1982 B.n531 B.n528 10.6151
R1983 B.n528 B.n527 10.6151
R1984 B.n527 B.n524 10.6151
R1985 B.n524 B.n523 10.6151
R1986 B.n523 B.n520 10.6151
R1987 B.n520 B.n519 10.6151
R1988 B.n519 B.n516 10.6151
R1989 B.n516 B.n515 10.6151
R1990 B.n515 B.n512 10.6151
R1991 B.n512 B.n511 10.6151
R1992 B.n511 B.n508 10.6151
R1993 B.n508 B.n507 10.6151
R1994 B.n507 B.n504 10.6151
R1995 B.n504 B.n503 10.6151
R1996 B.n503 B.n500 10.6151
R1997 B.n500 B.n499 10.6151
R1998 B.n499 B.n496 10.6151
R1999 B.n496 B.n495 10.6151
R2000 B.n495 B.n492 10.6151
R2001 B.n492 B.n491 10.6151
R2002 B.n491 B.n488 10.6151
R2003 B.n488 B.n487 10.6151
R2004 B.n487 B.n484 10.6151
R2005 B.n484 B.n483 10.6151
R2006 B.n483 B.n480 10.6151
R2007 B.n480 B.n479 10.6151
R2008 B.n479 B.n476 10.6151
R2009 B.n476 B.n475 10.6151
R2010 B.n475 B.n472 10.6151
R2011 B.n472 B.n471 10.6151
R2012 B.n471 B.n468 10.6151
R2013 B.n468 B.n467 10.6151
R2014 B.n467 B.n464 10.6151
R2015 B.n464 B.n463 10.6151
R2016 B.n463 B.n460 10.6151
R2017 B.n460 B.n459 10.6151
R2018 B.n459 B.n456 10.6151
R2019 B.n456 B.n455 10.6151
R2020 B.n455 B.n452 10.6151
R2021 B.n452 B.n451 10.6151
R2022 B.n451 B.n448 10.6151
R2023 B.n448 B.n447 10.6151
R2024 B.n447 B.n444 10.6151
R2025 B.n444 B.n443 10.6151
R2026 B.n697 B.n369 10.6151
R2027 B.n698 B.n697 10.6151
R2028 B.n699 B.n698 10.6151
R2029 B.n699 B.n361 10.6151
R2030 B.n709 B.n361 10.6151
R2031 B.n710 B.n709 10.6151
R2032 B.n711 B.n710 10.6151
R2033 B.n711 B.n353 10.6151
R2034 B.n721 B.n353 10.6151
R2035 B.n722 B.n721 10.6151
R2036 B.n724 B.n722 10.6151
R2037 B.n724 B.n723 10.6151
R2038 B.n723 B.n346 10.6151
R2039 B.n736 B.n346 10.6151
R2040 B.n737 B.n736 10.6151
R2041 B.n738 B.n737 10.6151
R2042 B.n739 B.n738 10.6151
R2043 B.n740 B.n739 10.6151
R2044 B.n743 B.n740 10.6151
R2045 B.n744 B.n743 10.6151
R2046 B.n745 B.n744 10.6151
R2047 B.n746 B.n745 10.6151
R2048 B.n748 B.n746 10.6151
R2049 B.n749 B.n748 10.6151
R2050 B.n750 B.n749 10.6151
R2051 B.n751 B.n750 10.6151
R2052 B.n753 B.n751 10.6151
R2053 B.n754 B.n753 10.6151
R2054 B.n755 B.n754 10.6151
R2055 B.n756 B.n755 10.6151
R2056 B.n757 B.n756 10.6151
R2057 B.n789 B.n1 10.6151
R2058 B.n789 B.n788 10.6151
R2059 B.n788 B.n787 10.6151
R2060 B.n787 B.n10 10.6151
R2061 B.n781 B.n10 10.6151
R2062 B.n781 B.n780 10.6151
R2063 B.n780 B.n779 10.6151
R2064 B.n779 B.n18 10.6151
R2065 B.n773 B.n18 10.6151
R2066 B.n773 B.n772 10.6151
R2067 B.n772 B.n771 10.6151
R2068 B.n771 B.n25 10.6151
R2069 B.n765 B.n25 10.6151
R2070 B.n765 B.n764 10.6151
R2071 B.n763 B.n32 10.6151
R2072 B.n103 B.n32 10.6151
R2073 B.n104 B.n103 10.6151
R2074 B.n107 B.n104 10.6151
R2075 B.n108 B.n107 10.6151
R2076 B.n111 B.n108 10.6151
R2077 B.n112 B.n111 10.6151
R2078 B.n115 B.n112 10.6151
R2079 B.n116 B.n115 10.6151
R2080 B.n119 B.n116 10.6151
R2081 B.n120 B.n119 10.6151
R2082 B.n123 B.n120 10.6151
R2083 B.n124 B.n123 10.6151
R2084 B.n127 B.n124 10.6151
R2085 B.n128 B.n127 10.6151
R2086 B.n131 B.n128 10.6151
R2087 B.n132 B.n131 10.6151
R2088 B.n135 B.n132 10.6151
R2089 B.n136 B.n135 10.6151
R2090 B.n139 B.n136 10.6151
R2091 B.n140 B.n139 10.6151
R2092 B.n143 B.n140 10.6151
R2093 B.n144 B.n143 10.6151
R2094 B.n147 B.n144 10.6151
R2095 B.n148 B.n147 10.6151
R2096 B.n151 B.n148 10.6151
R2097 B.n152 B.n151 10.6151
R2098 B.n155 B.n152 10.6151
R2099 B.n156 B.n155 10.6151
R2100 B.n159 B.n156 10.6151
R2101 B.n160 B.n159 10.6151
R2102 B.n163 B.n160 10.6151
R2103 B.n164 B.n163 10.6151
R2104 B.n167 B.n164 10.6151
R2105 B.n168 B.n167 10.6151
R2106 B.n171 B.n168 10.6151
R2107 B.n172 B.n171 10.6151
R2108 B.n175 B.n172 10.6151
R2109 B.n176 B.n175 10.6151
R2110 B.n179 B.n176 10.6151
R2111 B.n180 B.n179 10.6151
R2112 B.n183 B.n180 10.6151
R2113 B.n184 B.n183 10.6151
R2114 B.n187 B.n184 10.6151
R2115 B.n188 B.n187 10.6151
R2116 B.n191 B.n188 10.6151
R2117 B.n192 B.n191 10.6151
R2118 B.n195 B.n192 10.6151
R2119 B.n196 B.n195 10.6151
R2120 B.n199 B.n196 10.6151
R2121 B.n200 B.n199 10.6151
R2122 B.n203 B.n200 10.6151
R2123 B.n204 B.n203 10.6151
R2124 B.n207 B.n204 10.6151
R2125 B.n208 B.n207 10.6151
R2126 B.n211 B.n208 10.6151
R2127 B.n212 B.n211 10.6151
R2128 B.n216 B.n215 10.6151
R2129 B.n219 B.n216 10.6151
R2130 B.n220 B.n219 10.6151
R2131 B.n223 B.n220 10.6151
R2132 B.n224 B.n223 10.6151
R2133 B.n227 B.n224 10.6151
R2134 B.n228 B.n227 10.6151
R2135 B.n231 B.n228 10.6151
R2136 B.n236 B.n233 10.6151
R2137 B.n237 B.n236 10.6151
R2138 B.n240 B.n237 10.6151
R2139 B.n241 B.n240 10.6151
R2140 B.n244 B.n241 10.6151
R2141 B.n245 B.n244 10.6151
R2142 B.n248 B.n245 10.6151
R2143 B.n249 B.n248 10.6151
R2144 B.n252 B.n249 10.6151
R2145 B.n253 B.n252 10.6151
R2146 B.n256 B.n253 10.6151
R2147 B.n257 B.n256 10.6151
R2148 B.n260 B.n257 10.6151
R2149 B.n261 B.n260 10.6151
R2150 B.n264 B.n261 10.6151
R2151 B.n265 B.n264 10.6151
R2152 B.n268 B.n265 10.6151
R2153 B.n269 B.n268 10.6151
R2154 B.n272 B.n269 10.6151
R2155 B.n273 B.n272 10.6151
R2156 B.n276 B.n273 10.6151
R2157 B.n277 B.n276 10.6151
R2158 B.n280 B.n277 10.6151
R2159 B.n281 B.n280 10.6151
R2160 B.n284 B.n281 10.6151
R2161 B.n285 B.n284 10.6151
R2162 B.n288 B.n285 10.6151
R2163 B.n289 B.n288 10.6151
R2164 B.n292 B.n289 10.6151
R2165 B.n293 B.n292 10.6151
R2166 B.n296 B.n293 10.6151
R2167 B.n297 B.n296 10.6151
R2168 B.n300 B.n297 10.6151
R2169 B.n301 B.n300 10.6151
R2170 B.n304 B.n301 10.6151
R2171 B.n305 B.n304 10.6151
R2172 B.n308 B.n305 10.6151
R2173 B.n309 B.n308 10.6151
R2174 B.n312 B.n309 10.6151
R2175 B.n313 B.n312 10.6151
R2176 B.n316 B.n313 10.6151
R2177 B.n317 B.n316 10.6151
R2178 B.n320 B.n317 10.6151
R2179 B.n321 B.n320 10.6151
R2180 B.n324 B.n321 10.6151
R2181 B.n325 B.n324 10.6151
R2182 B.n328 B.n325 10.6151
R2183 B.n329 B.n328 10.6151
R2184 B.n332 B.n329 10.6151
R2185 B.n333 B.n332 10.6151
R2186 B.n336 B.n333 10.6151
R2187 B.n337 B.n336 10.6151
R2188 B.n340 B.n337 10.6151
R2189 B.n341 B.n340 10.6151
R2190 B.n344 B.n341 10.6151
R2191 B.n345 B.n344 10.6151
R2192 B.n758 B.n345 10.6151
R2193 B.n797 B.n0 8.11757
R2194 B.n797 B.n1 8.11757
R2195 B.n576 B.n575 7.18099
R2196 B.n559 B.n441 7.18099
R2197 B.n215 B.n101 7.18099
R2198 B.n232 B.n231 7.18099
R2199 B.n707 B.t3 5.79633
R2200 B.t7 B.n775 5.79633
R2201 B.n577 B.n576 3.43465
R2202 B.n556 B.n441 3.43465
R2203 B.n212 B.n101 3.43465
R2204 B.n233 B.n232 3.43465
R2205 B.n726 B.t0 1.93244
R2206 B.n12 B.t1 1.93244
R2207 VP.n0 VP.t1 706.266
R2208 VP.n0 VP.t0 661.899
R2209 VP VP.n0 0.0516364
R2210 VDD1.n92 VDD1.n0 289.615
R2211 VDD1.n189 VDD1.n97 289.615
R2212 VDD1.n93 VDD1.n92 185
R2213 VDD1.n91 VDD1.n90 185
R2214 VDD1.n4 VDD1.n3 185
R2215 VDD1.n85 VDD1.n84 185
R2216 VDD1.n83 VDD1.n82 185
R2217 VDD1.n8 VDD1.n7 185
R2218 VDD1.n12 VDD1.n10 185
R2219 VDD1.n77 VDD1.n76 185
R2220 VDD1.n75 VDD1.n74 185
R2221 VDD1.n14 VDD1.n13 185
R2222 VDD1.n69 VDD1.n68 185
R2223 VDD1.n67 VDD1.n66 185
R2224 VDD1.n18 VDD1.n17 185
R2225 VDD1.n61 VDD1.n60 185
R2226 VDD1.n59 VDD1.n58 185
R2227 VDD1.n22 VDD1.n21 185
R2228 VDD1.n53 VDD1.n52 185
R2229 VDD1.n51 VDD1.n50 185
R2230 VDD1.n26 VDD1.n25 185
R2231 VDD1.n45 VDD1.n44 185
R2232 VDD1.n43 VDD1.n42 185
R2233 VDD1.n30 VDD1.n29 185
R2234 VDD1.n37 VDD1.n36 185
R2235 VDD1.n35 VDD1.n34 185
R2236 VDD1.n130 VDD1.n129 185
R2237 VDD1.n132 VDD1.n131 185
R2238 VDD1.n125 VDD1.n124 185
R2239 VDD1.n138 VDD1.n137 185
R2240 VDD1.n140 VDD1.n139 185
R2241 VDD1.n121 VDD1.n120 185
R2242 VDD1.n146 VDD1.n145 185
R2243 VDD1.n148 VDD1.n147 185
R2244 VDD1.n117 VDD1.n116 185
R2245 VDD1.n154 VDD1.n153 185
R2246 VDD1.n156 VDD1.n155 185
R2247 VDD1.n113 VDD1.n112 185
R2248 VDD1.n162 VDD1.n161 185
R2249 VDD1.n164 VDD1.n163 185
R2250 VDD1.n109 VDD1.n108 185
R2251 VDD1.n171 VDD1.n170 185
R2252 VDD1.n172 VDD1.n107 185
R2253 VDD1.n174 VDD1.n173 185
R2254 VDD1.n105 VDD1.n104 185
R2255 VDD1.n180 VDD1.n179 185
R2256 VDD1.n182 VDD1.n181 185
R2257 VDD1.n101 VDD1.n100 185
R2258 VDD1.n188 VDD1.n187 185
R2259 VDD1.n190 VDD1.n189 185
R2260 VDD1.n33 VDD1.t0 147.659
R2261 VDD1.n128 VDD1.t1 147.659
R2262 VDD1.n92 VDD1.n91 104.615
R2263 VDD1.n91 VDD1.n3 104.615
R2264 VDD1.n84 VDD1.n3 104.615
R2265 VDD1.n84 VDD1.n83 104.615
R2266 VDD1.n83 VDD1.n7 104.615
R2267 VDD1.n12 VDD1.n7 104.615
R2268 VDD1.n76 VDD1.n12 104.615
R2269 VDD1.n76 VDD1.n75 104.615
R2270 VDD1.n75 VDD1.n13 104.615
R2271 VDD1.n68 VDD1.n13 104.615
R2272 VDD1.n68 VDD1.n67 104.615
R2273 VDD1.n67 VDD1.n17 104.615
R2274 VDD1.n60 VDD1.n17 104.615
R2275 VDD1.n60 VDD1.n59 104.615
R2276 VDD1.n59 VDD1.n21 104.615
R2277 VDD1.n52 VDD1.n21 104.615
R2278 VDD1.n52 VDD1.n51 104.615
R2279 VDD1.n51 VDD1.n25 104.615
R2280 VDD1.n44 VDD1.n25 104.615
R2281 VDD1.n44 VDD1.n43 104.615
R2282 VDD1.n43 VDD1.n29 104.615
R2283 VDD1.n36 VDD1.n29 104.615
R2284 VDD1.n36 VDD1.n35 104.615
R2285 VDD1.n131 VDD1.n130 104.615
R2286 VDD1.n131 VDD1.n124 104.615
R2287 VDD1.n138 VDD1.n124 104.615
R2288 VDD1.n139 VDD1.n138 104.615
R2289 VDD1.n139 VDD1.n120 104.615
R2290 VDD1.n146 VDD1.n120 104.615
R2291 VDD1.n147 VDD1.n146 104.615
R2292 VDD1.n147 VDD1.n116 104.615
R2293 VDD1.n154 VDD1.n116 104.615
R2294 VDD1.n155 VDD1.n154 104.615
R2295 VDD1.n155 VDD1.n112 104.615
R2296 VDD1.n162 VDD1.n112 104.615
R2297 VDD1.n163 VDD1.n162 104.615
R2298 VDD1.n163 VDD1.n108 104.615
R2299 VDD1.n171 VDD1.n108 104.615
R2300 VDD1.n172 VDD1.n171 104.615
R2301 VDD1.n173 VDD1.n172 104.615
R2302 VDD1.n173 VDD1.n104 104.615
R2303 VDD1.n180 VDD1.n104 104.615
R2304 VDD1.n181 VDD1.n180 104.615
R2305 VDD1.n181 VDD1.n100 104.615
R2306 VDD1.n188 VDD1.n100 104.615
R2307 VDD1.n189 VDD1.n188 104.615
R2308 VDD1 VDD1.n193 89.7834
R2309 VDD1.n35 VDD1.t0 52.3082
R2310 VDD1.n130 VDD1.t1 52.3082
R2311 VDD1 VDD1.n96 48.416
R2312 VDD1.n34 VDD1.n33 15.6677
R2313 VDD1.n129 VDD1.n128 15.6677
R2314 VDD1.n10 VDD1.n8 13.1884
R2315 VDD1.n174 VDD1.n105 13.1884
R2316 VDD1.n82 VDD1.n81 12.8005
R2317 VDD1.n78 VDD1.n77 12.8005
R2318 VDD1.n37 VDD1.n32 12.8005
R2319 VDD1.n132 VDD1.n127 12.8005
R2320 VDD1.n175 VDD1.n107 12.8005
R2321 VDD1.n179 VDD1.n178 12.8005
R2322 VDD1.n85 VDD1.n6 12.0247
R2323 VDD1.n74 VDD1.n11 12.0247
R2324 VDD1.n38 VDD1.n30 12.0247
R2325 VDD1.n133 VDD1.n125 12.0247
R2326 VDD1.n170 VDD1.n169 12.0247
R2327 VDD1.n182 VDD1.n103 12.0247
R2328 VDD1.n86 VDD1.n4 11.249
R2329 VDD1.n73 VDD1.n14 11.249
R2330 VDD1.n42 VDD1.n41 11.249
R2331 VDD1.n137 VDD1.n136 11.249
R2332 VDD1.n168 VDD1.n109 11.249
R2333 VDD1.n183 VDD1.n101 11.249
R2334 VDD1.n90 VDD1.n89 10.4732
R2335 VDD1.n70 VDD1.n69 10.4732
R2336 VDD1.n45 VDD1.n28 10.4732
R2337 VDD1.n140 VDD1.n123 10.4732
R2338 VDD1.n165 VDD1.n164 10.4732
R2339 VDD1.n187 VDD1.n186 10.4732
R2340 VDD1.n93 VDD1.n2 9.69747
R2341 VDD1.n66 VDD1.n16 9.69747
R2342 VDD1.n46 VDD1.n26 9.69747
R2343 VDD1.n141 VDD1.n121 9.69747
R2344 VDD1.n161 VDD1.n111 9.69747
R2345 VDD1.n190 VDD1.n99 9.69747
R2346 VDD1.n96 VDD1.n95 9.45567
R2347 VDD1.n193 VDD1.n192 9.45567
R2348 VDD1.n20 VDD1.n19 9.3005
R2349 VDD1.n63 VDD1.n62 9.3005
R2350 VDD1.n65 VDD1.n64 9.3005
R2351 VDD1.n16 VDD1.n15 9.3005
R2352 VDD1.n71 VDD1.n70 9.3005
R2353 VDD1.n73 VDD1.n72 9.3005
R2354 VDD1.n11 VDD1.n9 9.3005
R2355 VDD1.n79 VDD1.n78 9.3005
R2356 VDD1.n95 VDD1.n94 9.3005
R2357 VDD1.n2 VDD1.n1 9.3005
R2358 VDD1.n89 VDD1.n88 9.3005
R2359 VDD1.n87 VDD1.n86 9.3005
R2360 VDD1.n6 VDD1.n5 9.3005
R2361 VDD1.n81 VDD1.n80 9.3005
R2362 VDD1.n57 VDD1.n56 9.3005
R2363 VDD1.n55 VDD1.n54 9.3005
R2364 VDD1.n24 VDD1.n23 9.3005
R2365 VDD1.n49 VDD1.n48 9.3005
R2366 VDD1.n47 VDD1.n46 9.3005
R2367 VDD1.n28 VDD1.n27 9.3005
R2368 VDD1.n41 VDD1.n40 9.3005
R2369 VDD1.n39 VDD1.n38 9.3005
R2370 VDD1.n32 VDD1.n31 9.3005
R2371 VDD1.n192 VDD1.n191 9.3005
R2372 VDD1.n99 VDD1.n98 9.3005
R2373 VDD1.n186 VDD1.n185 9.3005
R2374 VDD1.n184 VDD1.n183 9.3005
R2375 VDD1.n103 VDD1.n102 9.3005
R2376 VDD1.n178 VDD1.n177 9.3005
R2377 VDD1.n150 VDD1.n149 9.3005
R2378 VDD1.n119 VDD1.n118 9.3005
R2379 VDD1.n144 VDD1.n143 9.3005
R2380 VDD1.n142 VDD1.n141 9.3005
R2381 VDD1.n123 VDD1.n122 9.3005
R2382 VDD1.n136 VDD1.n135 9.3005
R2383 VDD1.n134 VDD1.n133 9.3005
R2384 VDD1.n127 VDD1.n126 9.3005
R2385 VDD1.n152 VDD1.n151 9.3005
R2386 VDD1.n115 VDD1.n114 9.3005
R2387 VDD1.n158 VDD1.n157 9.3005
R2388 VDD1.n160 VDD1.n159 9.3005
R2389 VDD1.n111 VDD1.n110 9.3005
R2390 VDD1.n166 VDD1.n165 9.3005
R2391 VDD1.n168 VDD1.n167 9.3005
R2392 VDD1.n169 VDD1.n106 9.3005
R2393 VDD1.n176 VDD1.n175 9.3005
R2394 VDD1.n94 VDD1.n0 8.92171
R2395 VDD1.n65 VDD1.n18 8.92171
R2396 VDD1.n50 VDD1.n49 8.92171
R2397 VDD1.n145 VDD1.n144 8.92171
R2398 VDD1.n160 VDD1.n113 8.92171
R2399 VDD1.n191 VDD1.n97 8.92171
R2400 VDD1.n62 VDD1.n61 8.14595
R2401 VDD1.n53 VDD1.n24 8.14595
R2402 VDD1.n148 VDD1.n119 8.14595
R2403 VDD1.n157 VDD1.n156 8.14595
R2404 VDD1.n58 VDD1.n20 7.3702
R2405 VDD1.n54 VDD1.n22 7.3702
R2406 VDD1.n149 VDD1.n117 7.3702
R2407 VDD1.n153 VDD1.n115 7.3702
R2408 VDD1.n58 VDD1.n57 6.59444
R2409 VDD1.n57 VDD1.n22 6.59444
R2410 VDD1.n152 VDD1.n117 6.59444
R2411 VDD1.n153 VDD1.n152 6.59444
R2412 VDD1.n61 VDD1.n20 5.81868
R2413 VDD1.n54 VDD1.n53 5.81868
R2414 VDD1.n149 VDD1.n148 5.81868
R2415 VDD1.n156 VDD1.n115 5.81868
R2416 VDD1.n96 VDD1.n0 5.04292
R2417 VDD1.n62 VDD1.n18 5.04292
R2418 VDD1.n50 VDD1.n24 5.04292
R2419 VDD1.n145 VDD1.n119 5.04292
R2420 VDD1.n157 VDD1.n113 5.04292
R2421 VDD1.n193 VDD1.n97 5.04292
R2422 VDD1.n33 VDD1.n31 4.38563
R2423 VDD1.n128 VDD1.n126 4.38563
R2424 VDD1.n94 VDD1.n93 4.26717
R2425 VDD1.n66 VDD1.n65 4.26717
R2426 VDD1.n49 VDD1.n26 4.26717
R2427 VDD1.n144 VDD1.n121 4.26717
R2428 VDD1.n161 VDD1.n160 4.26717
R2429 VDD1.n191 VDD1.n190 4.26717
R2430 VDD1.n90 VDD1.n2 3.49141
R2431 VDD1.n69 VDD1.n16 3.49141
R2432 VDD1.n46 VDD1.n45 3.49141
R2433 VDD1.n141 VDD1.n140 3.49141
R2434 VDD1.n164 VDD1.n111 3.49141
R2435 VDD1.n187 VDD1.n99 3.49141
R2436 VDD1.n89 VDD1.n4 2.71565
R2437 VDD1.n70 VDD1.n14 2.71565
R2438 VDD1.n42 VDD1.n28 2.71565
R2439 VDD1.n137 VDD1.n123 2.71565
R2440 VDD1.n165 VDD1.n109 2.71565
R2441 VDD1.n186 VDD1.n101 2.71565
R2442 VDD1.n86 VDD1.n85 1.93989
R2443 VDD1.n74 VDD1.n73 1.93989
R2444 VDD1.n41 VDD1.n30 1.93989
R2445 VDD1.n136 VDD1.n125 1.93989
R2446 VDD1.n170 VDD1.n168 1.93989
R2447 VDD1.n183 VDD1.n182 1.93989
R2448 VDD1.n82 VDD1.n6 1.16414
R2449 VDD1.n77 VDD1.n11 1.16414
R2450 VDD1.n38 VDD1.n37 1.16414
R2451 VDD1.n133 VDD1.n132 1.16414
R2452 VDD1.n169 VDD1.n107 1.16414
R2453 VDD1.n179 VDD1.n103 1.16414
R2454 VDD1.n81 VDD1.n8 0.388379
R2455 VDD1.n78 VDD1.n10 0.388379
R2456 VDD1.n34 VDD1.n32 0.388379
R2457 VDD1.n129 VDD1.n127 0.388379
R2458 VDD1.n175 VDD1.n174 0.388379
R2459 VDD1.n178 VDD1.n105 0.388379
R2460 VDD1.n95 VDD1.n1 0.155672
R2461 VDD1.n88 VDD1.n1 0.155672
R2462 VDD1.n88 VDD1.n87 0.155672
R2463 VDD1.n87 VDD1.n5 0.155672
R2464 VDD1.n80 VDD1.n5 0.155672
R2465 VDD1.n80 VDD1.n79 0.155672
R2466 VDD1.n79 VDD1.n9 0.155672
R2467 VDD1.n72 VDD1.n9 0.155672
R2468 VDD1.n72 VDD1.n71 0.155672
R2469 VDD1.n71 VDD1.n15 0.155672
R2470 VDD1.n64 VDD1.n15 0.155672
R2471 VDD1.n64 VDD1.n63 0.155672
R2472 VDD1.n63 VDD1.n19 0.155672
R2473 VDD1.n56 VDD1.n19 0.155672
R2474 VDD1.n56 VDD1.n55 0.155672
R2475 VDD1.n55 VDD1.n23 0.155672
R2476 VDD1.n48 VDD1.n23 0.155672
R2477 VDD1.n48 VDD1.n47 0.155672
R2478 VDD1.n47 VDD1.n27 0.155672
R2479 VDD1.n40 VDD1.n27 0.155672
R2480 VDD1.n40 VDD1.n39 0.155672
R2481 VDD1.n39 VDD1.n31 0.155672
R2482 VDD1.n134 VDD1.n126 0.155672
R2483 VDD1.n135 VDD1.n134 0.155672
R2484 VDD1.n135 VDD1.n122 0.155672
R2485 VDD1.n142 VDD1.n122 0.155672
R2486 VDD1.n143 VDD1.n142 0.155672
R2487 VDD1.n143 VDD1.n118 0.155672
R2488 VDD1.n150 VDD1.n118 0.155672
R2489 VDD1.n151 VDD1.n150 0.155672
R2490 VDD1.n151 VDD1.n114 0.155672
R2491 VDD1.n158 VDD1.n114 0.155672
R2492 VDD1.n159 VDD1.n158 0.155672
R2493 VDD1.n159 VDD1.n110 0.155672
R2494 VDD1.n166 VDD1.n110 0.155672
R2495 VDD1.n167 VDD1.n166 0.155672
R2496 VDD1.n167 VDD1.n106 0.155672
R2497 VDD1.n176 VDD1.n106 0.155672
R2498 VDD1.n177 VDD1.n176 0.155672
R2499 VDD1.n177 VDD1.n102 0.155672
R2500 VDD1.n184 VDD1.n102 0.155672
R2501 VDD1.n185 VDD1.n184 0.155672
R2502 VDD1.n185 VDD1.n98 0.155672
R2503 VDD1.n192 VDD1.n98 0.155672
C0 VP VTAIL 2.36777f
C1 VP VN 5.673759f
C2 VDD1 VDD2 0.485244f
C3 VDD1 VTAIL 7.2295f
C4 VDD2 VTAIL 7.262919f
C5 VDD1 VN 0.149022f
C6 VDD2 VN 3.06554f
C7 VDD1 VP 3.17602f
C8 VDD2 VP 0.26524f
C9 VN VTAIL 2.35303f
C10 VDD2 B 4.823386f
C11 VDD1 B 7.688019f
C12 VTAIL B 8.604833f
C13 VN B 10.64818f
C14 VP B 4.670987f
C15 VDD1.n0 B 0.02761f
C16 VDD1.n1 B 0.020428f
C17 VDD1.n2 B 0.010977f
C18 VDD1.n3 B 0.025945f
C19 VDD1.n4 B 0.011623f
C20 VDD1.n5 B 0.020428f
C21 VDD1.n6 B 0.010977f
C22 VDD1.n7 B 0.025945f
C23 VDD1.n8 B 0.0113f
C24 VDD1.n9 B 0.020428f
C25 VDD1.n10 B 0.0113f
C26 VDD1.n11 B 0.010977f
C27 VDD1.n12 B 0.025945f
C28 VDD1.n13 B 0.025945f
C29 VDD1.n14 B 0.011623f
C30 VDD1.n15 B 0.020428f
C31 VDD1.n16 B 0.010977f
C32 VDD1.n17 B 0.025945f
C33 VDD1.n18 B 0.011623f
C34 VDD1.n19 B 0.020428f
C35 VDD1.n20 B 0.010977f
C36 VDD1.n21 B 0.025945f
C37 VDD1.n22 B 0.011623f
C38 VDD1.n23 B 0.020428f
C39 VDD1.n24 B 0.010977f
C40 VDD1.n25 B 0.025945f
C41 VDD1.n26 B 0.011623f
C42 VDD1.n27 B 0.020428f
C43 VDD1.n28 B 0.010977f
C44 VDD1.n29 B 0.025945f
C45 VDD1.n30 B 0.011623f
C46 VDD1.n31 B 1.56123f
C47 VDD1.n32 B 0.010977f
C48 VDD1.t0 B 0.042955f
C49 VDD1.n33 B 0.145936f
C50 VDD1.n34 B 0.015327f
C51 VDD1.n35 B 0.019459f
C52 VDD1.n36 B 0.025945f
C53 VDD1.n37 B 0.011623f
C54 VDD1.n38 B 0.010977f
C55 VDD1.n39 B 0.020428f
C56 VDD1.n40 B 0.020428f
C57 VDD1.n41 B 0.010977f
C58 VDD1.n42 B 0.011623f
C59 VDD1.n43 B 0.025945f
C60 VDD1.n44 B 0.025945f
C61 VDD1.n45 B 0.011623f
C62 VDD1.n46 B 0.010977f
C63 VDD1.n47 B 0.020428f
C64 VDD1.n48 B 0.020428f
C65 VDD1.n49 B 0.010977f
C66 VDD1.n50 B 0.011623f
C67 VDD1.n51 B 0.025945f
C68 VDD1.n52 B 0.025945f
C69 VDD1.n53 B 0.011623f
C70 VDD1.n54 B 0.010977f
C71 VDD1.n55 B 0.020428f
C72 VDD1.n56 B 0.020428f
C73 VDD1.n57 B 0.010977f
C74 VDD1.n58 B 0.011623f
C75 VDD1.n59 B 0.025945f
C76 VDD1.n60 B 0.025945f
C77 VDD1.n61 B 0.011623f
C78 VDD1.n62 B 0.010977f
C79 VDD1.n63 B 0.020428f
C80 VDD1.n64 B 0.020428f
C81 VDD1.n65 B 0.010977f
C82 VDD1.n66 B 0.011623f
C83 VDD1.n67 B 0.025945f
C84 VDD1.n68 B 0.025945f
C85 VDD1.n69 B 0.011623f
C86 VDD1.n70 B 0.010977f
C87 VDD1.n71 B 0.020428f
C88 VDD1.n72 B 0.020428f
C89 VDD1.n73 B 0.010977f
C90 VDD1.n74 B 0.011623f
C91 VDD1.n75 B 0.025945f
C92 VDD1.n76 B 0.025945f
C93 VDD1.n77 B 0.011623f
C94 VDD1.n78 B 0.010977f
C95 VDD1.n79 B 0.020428f
C96 VDD1.n80 B 0.020428f
C97 VDD1.n81 B 0.010977f
C98 VDD1.n82 B 0.011623f
C99 VDD1.n83 B 0.025945f
C100 VDD1.n84 B 0.025945f
C101 VDD1.n85 B 0.011623f
C102 VDD1.n86 B 0.010977f
C103 VDD1.n87 B 0.020428f
C104 VDD1.n88 B 0.020428f
C105 VDD1.n89 B 0.010977f
C106 VDD1.n90 B 0.011623f
C107 VDD1.n91 B 0.025945f
C108 VDD1.n92 B 0.054218f
C109 VDD1.n93 B 0.011623f
C110 VDD1.n94 B 0.010977f
C111 VDD1.n95 B 0.046101f
C112 VDD1.n96 B 0.044624f
C113 VDD1.n97 B 0.02761f
C114 VDD1.n98 B 0.020428f
C115 VDD1.n99 B 0.010977f
C116 VDD1.n100 B 0.025945f
C117 VDD1.n101 B 0.011623f
C118 VDD1.n102 B 0.020428f
C119 VDD1.n103 B 0.010977f
C120 VDD1.n104 B 0.025945f
C121 VDD1.n105 B 0.0113f
C122 VDD1.n106 B 0.020428f
C123 VDD1.n107 B 0.011623f
C124 VDD1.n108 B 0.025945f
C125 VDD1.n109 B 0.011623f
C126 VDD1.n110 B 0.020428f
C127 VDD1.n111 B 0.010977f
C128 VDD1.n112 B 0.025945f
C129 VDD1.n113 B 0.011623f
C130 VDD1.n114 B 0.020428f
C131 VDD1.n115 B 0.010977f
C132 VDD1.n116 B 0.025945f
C133 VDD1.n117 B 0.011623f
C134 VDD1.n118 B 0.020428f
C135 VDD1.n119 B 0.010977f
C136 VDD1.n120 B 0.025945f
C137 VDD1.n121 B 0.011623f
C138 VDD1.n122 B 0.020428f
C139 VDD1.n123 B 0.010977f
C140 VDD1.n124 B 0.025945f
C141 VDD1.n125 B 0.011623f
C142 VDD1.n126 B 1.56123f
C143 VDD1.n127 B 0.010977f
C144 VDD1.t1 B 0.042955f
C145 VDD1.n128 B 0.145936f
C146 VDD1.n129 B 0.015327f
C147 VDD1.n130 B 0.019459f
C148 VDD1.n131 B 0.025945f
C149 VDD1.n132 B 0.011623f
C150 VDD1.n133 B 0.010977f
C151 VDD1.n134 B 0.020428f
C152 VDD1.n135 B 0.020428f
C153 VDD1.n136 B 0.010977f
C154 VDD1.n137 B 0.011623f
C155 VDD1.n138 B 0.025945f
C156 VDD1.n139 B 0.025945f
C157 VDD1.n140 B 0.011623f
C158 VDD1.n141 B 0.010977f
C159 VDD1.n142 B 0.020428f
C160 VDD1.n143 B 0.020428f
C161 VDD1.n144 B 0.010977f
C162 VDD1.n145 B 0.011623f
C163 VDD1.n146 B 0.025945f
C164 VDD1.n147 B 0.025945f
C165 VDD1.n148 B 0.011623f
C166 VDD1.n149 B 0.010977f
C167 VDD1.n150 B 0.020428f
C168 VDD1.n151 B 0.020428f
C169 VDD1.n152 B 0.010977f
C170 VDD1.n153 B 0.011623f
C171 VDD1.n154 B 0.025945f
C172 VDD1.n155 B 0.025945f
C173 VDD1.n156 B 0.011623f
C174 VDD1.n157 B 0.010977f
C175 VDD1.n158 B 0.020428f
C176 VDD1.n159 B 0.020428f
C177 VDD1.n160 B 0.010977f
C178 VDD1.n161 B 0.011623f
C179 VDD1.n162 B 0.025945f
C180 VDD1.n163 B 0.025945f
C181 VDD1.n164 B 0.011623f
C182 VDD1.n165 B 0.010977f
C183 VDD1.n166 B 0.020428f
C184 VDD1.n167 B 0.020428f
C185 VDD1.n168 B 0.010977f
C186 VDD1.n169 B 0.010977f
C187 VDD1.n170 B 0.011623f
C188 VDD1.n171 B 0.025945f
C189 VDD1.n172 B 0.025945f
C190 VDD1.n173 B 0.025945f
C191 VDD1.n174 B 0.0113f
C192 VDD1.n175 B 0.010977f
C193 VDD1.n176 B 0.020428f
C194 VDD1.n177 B 0.020428f
C195 VDD1.n178 B 0.010977f
C196 VDD1.n179 B 0.011623f
C197 VDD1.n180 B 0.025945f
C198 VDD1.n181 B 0.025945f
C199 VDD1.n182 B 0.011623f
C200 VDD1.n183 B 0.010977f
C201 VDD1.n184 B 0.020428f
C202 VDD1.n185 B 0.020428f
C203 VDD1.n186 B 0.010977f
C204 VDD1.n187 B 0.011623f
C205 VDD1.n188 B 0.025945f
C206 VDD1.n189 B 0.054218f
C207 VDD1.n190 B 0.011623f
C208 VDD1.n191 B 0.010977f
C209 VDD1.n192 B 0.046101f
C210 VDD1.n193 B 0.707413f
C211 VP.t1 B 2.7831f
C212 VP.t0 B 2.59236f
C213 VP.n0 B 5.89932f
C214 VDD2.n0 B 0.027812f
C215 VDD2.n1 B 0.020577f
C216 VDD2.n2 B 0.011057f
C217 VDD2.n3 B 0.026135f
C218 VDD2.n4 B 0.011708f
C219 VDD2.n5 B 0.020577f
C220 VDD2.n6 B 0.011057f
C221 VDD2.n7 B 0.026135f
C222 VDD2.n8 B 0.011382f
C223 VDD2.n9 B 0.020577f
C224 VDD2.n10 B 0.011708f
C225 VDD2.n11 B 0.026135f
C226 VDD2.n12 B 0.011708f
C227 VDD2.n13 B 0.020577f
C228 VDD2.n14 B 0.011057f
C229 VDD2.n15 B 0.026135f
C230 VDD2.n16 B 0.011708f
C231 VDD2.n17 B 0.020577f
C232 VDD2.n18 B 0.011057f
C233 VDD2.n19 B 0.026135f
C234 VDD2.n20 B 0.011708f
C235 VDD2.n21 B 0.020577f
C236 VDD2.n22 B 0.011057f
C237 VDD2.n23 B 0.026135f
C238 VDD2.n24 B 0.011708f
C239 VDD2.n25 B 0.020577f
C240 VDD2.n26 B 0.011057f
C241 VDD2.n27 B 0.026135f
C242 VDD2.n28 B 0.011708f
C243 VDD2.n29 B 1.57264f
C244 VDD2.n30 B 0.011057f
C245 VDD2.t0 B 0.043269f
C246 VDD2.n31 B 0.147002f
C247 VDD2.n32 B 0.015439f
C248 VDD2.n33 B 0.019601f
C249 VDD2.n34 B 0.026135f
C250 VDD2.n35 B 0.011708f
C251 VDD2.n36 B 0.011057f
C252 VDD2.n37 B 0.020577f
C253 VDD2.n38 B 0.020577f
C254 VDD2.n39 B 0.011057f
C255 VDD2.n40 B 0.011708f
C256 VDD2.n41 B 0.026135f
C257 VDD2.n42 B 0.026135f
C258 VDD2.n43 B 0.011708f
C259 VDD2.n44 B 0.011057f
C260 VDD2.n45 B 0.020577f
C261 VDD2.n46 B 0.020577f
C262 VDD2.n47 B 0.011057f
C263 VDD2.n48 B 0.011708f
C264 VDD2.n49 B 0.026135f
C265 VDD2.n50 B 0.026135f
C266 VDD2.n51 B 0.011708f
C267 VDD2.n52 B 0.011057f
C268 VDD2.n53 B 0.020577f
C269 VDD2.n54 B 0.020577f
C270 VDD2.n55 B 0.011057f
C271 VDD2.n56 B 0.011708f
C272 VDD2.n57 B 0.026135f
C273 VDD2.n58 B 0.026135f
C274 VDD2.n59 B 0.011708f
C275 VDD2.n60 B 0.011057f
C276 VDD2.n61 B 0.020577f
C277 VDD2.n62 B 0.020577f
C278 VDD2.n63 B 0.011057f
C279 VDD2.n64 B 0.011708f
C280 VDD2.n65 B 0.026135f
C281 VDD2.n66 B 0.026135f
C282 VDD2.n67 B 0.011708f
C283 VDD2.n68 B 0.011057f
C284 VDD2.n69 B 0.020577f
C285 VDD2.n70 B 0.020577f
C286 VDD2.n71 B 0.011057f
C287 VDD2.n72 B 0.011057f
C288 VDD2.n73 B 0.011708f
C289 VDD2.n74 B 0.026135f
C290 VDD2.n75 B 0.026135f
C291 VDD2.n76 B 0.026135f
C292 VDD2.n77 B 0.011382f
C293 VDD2.n78 B 0.011057f
C294 VDD2.n79 B 0.020577f
C295 VDD2.n80 B 0.020577f
C296 VDD2.n81 B 0.011057f
C297 VDD2.n82 B 0.011708f
C298 VDD2.n83 B 0.026135f
C299 VDD2.n84 B 0.026135f
C300 VDD2.n85 B 0.011708f
C301 VDD2.n86 B 0.011057f
C302 VDD2.n87 B 0.020577f
C303 VDD2.n88 B 0.020577f
C304 VDD2.n89 B 0.011057f
C305 VDD2.n90 B 0.011708f
C306 VDD2.n91 B 0.026135f
C307 VDD2.n92 B 0.054614f
C308 VDD2.n93 B 0.011708f
C309 VDD2.n94 B 0.011057f
C310 VDD2.n95 B 0.046438f
C311 VDD2.n96 B 0.680992f
C312 VDD2.n97 B 0.027812f
C313 VDD2.n98 B 0.020577f
C314 VDD2.n99 B 0.011057f
C315 VDD2.n100 B 0.026135f
C316 VDD2.n101 B 0.011708f
C317 VDD2.n102 B 0.020577f
C318 VDD2.n103 B 0.011057f
C319 VDD2.n104 B 0.026135f
C320 VDD2.n105 B 0.011382f
C321 VDD2.n106 B 0.020577f
C322 VDD2.n107 B 0.011382f
C323 VDD2.n108 B 0.011057f
C324 VDD2.n109 B 0.026135f
C325 VDD2.n110 B 0.026135f
C326 VDD2.n111 B 0.011708f
C327 VDD2.n112 B 0.020577f
C328 VDD2.n113 B 0.011057f
C329 VDD2.n114 B 0.026135f
C330 VDD2.n115 B 0.011708f
C331 VDD2.n116 B 0.020577f
C332 VDD2.n117 B 0.011057f
C333 VDD2.n118 B 0.026135f
C334 VDD2.n119 B 0.011708f
C335 VDD2.n120 B 0.020577f
C336 VDD2.n121 B 0.011057f
C337 VDD2.n122 B 0.026135f
C338 VDD2.n123 B 0.011708f
C339 VDD2.n124 B 0.020577f
C340 VDD2.n125 B 0.011057f
C341 VDD2.n126 B 0.026135f
C342 VDD2.n127 B 0.011708f
C343 VDD2.n128 B 1.57264f
C344 VDD2.n129 B 0.011057f
C345 VDD2.t1 B 0.043269f
C346 VDD2.n130 B 0.147002f
C347 VDD2.n131 B 0.015439f
C348 VDD2.n132 B 0.019601f
C349 VDD2.n133 B 0.026135f
C350 VDD2.n134 B 0.011708f
C351 VDD2.n135 B 0.011057f
C352 VDD2.n136 B 0.020577f
C353 VDD2.n137 B 0.020577f
C354 VDD2.n138 B 0.011057f
C355 VDD2.n139 B 0.011708f
C356 VDD2.n140 B 0.026135f
C357 VDD2.n141 B 0.026135f
C358 VDD2.n142 B 0.011708f
C359 VDD2.n143 B 0.011057f
C360 VDD2.n144 B 0.020577f
C361 VDD2.n145 B 0.020577f
C362 VDD2.n146 B 0.011057f
C363 VDD2.n147 B 0.011708f
C364 VDD2.n148 B 0.026135f
C365 VDD2.n149 B 0.026135f
C366 VDD2.n150 B 0.011708f
C367 VDD2.n151 B 0.011057f
C368 VDD2.n152 B 0.020577f
C369 VDD2.n153 B 0.020577f
C370 VDD2.n154 B 0.011057f
C371 VDD2.n155 B 0.011708f
C372 VDD2.n156 B 0.026135f
C373 VDD2.n157 B 0.026135f
C374 VDD2.n158 B 0.011708f
C375 VDD2.n159 B 0.011057f
C376 VDD2.n160 B 0.020577f
C377 VDD2.n161 B 0.020577f
C378 VDD2.n162 B 0.011057f
C379 VDD2.n163 B 0.011708f
C380 VDD2.n164 B 0.026135f
C381 VDD2.n165 B 0.026135f
C382 VDD2.n166 B 0.011708f
C383 VDD2.n167 B 0.011057f
C384 VDD2.n168 B 0.020577f
C385 VDD2.n169 B 0.020577f
C386 VDD2.n170 B 0.011057f
C387 VDD2.n171 B 0.011708f
C388 VDD2.n172 B 0.026135f
C389 VDD2.n173 B 0.026135f
C390 VDD2.n174 B 0.011708f
C391 VDD2.n175 B 0.011057f
C392 VDD2.n176 B 0.020577f
C393 VDD2.n177 B 0.020577f
C394 VDD2.n178 B 0.011057f
C395 VDD2.n179 B 0.011708f
C396 VDD2.n180 B 0.026135f
C397 VDD2.n181 B 0.026135f
C398 VDD2.n182 B 0.011708f
C399 VDD2.n183 B 0.011057f
C400 VDD2.n184 B 0.020577f
C401 VDD2.n185 B 0.020577f
C402 VDD2.n186 B 0.011057f
C403 VDD2.n187 B 0.011708f
C404 VDD2.n188 B 0.026135f
C405 VDD2.n189 B 0.054614f
C406 VDD2.n190 B 0.011708f
C407 VDD2.n191 B 0.011057f
C408 VDD2.n192 B 0.046438f
C409 VDD2.n193 B 0.044539f
C410 VDD2.n194 B 2.70276f
C411 VTAIL.n0 B 0.027066f
C412 VTAIL.n1 B 0.020025f
C413 VTAIL.n2 B 0.010761f
C414 VTAIL.n3 B 0.025434f
C415 VTAIL.n4 B 0.011394f
C416 VTAIL.n5 B 0.020025f
C417 VTAIL.n6 B 0.010761f
C418 VTAIL.n7 B 0.025434f
C419 VTAIL.n8 B 0.011077f
C420 VTAIL.n9 B 0.020025f
C421 VTAIL.n10 B 0.011394f
C422 VTAIL.n11 B 0.025434f
C423 VTAIL.n12 B 0.011394f
C424 VTAIL.n13 B 0.020025f
C425 VTAIL.n14 B 0.010761f
C426 VTAIL.n15 B 0.025434f
C427 VTAIL.n16 B 0.011394f
C428 VTAIL.n17 B 0.020025f
C429 VTAIL.n18 B 0.010761f
C430 VTAIL.n19 B 0.025434f
C431 VTAIL.n20 B 0.011394f
C432 VTAIL.n21 B 0.020025f
C433 VTAIL.n22 B 0.010761f
C434 VTAIL.n23 B 0.025434f
C435 VTAIL.n24 B 0.011394f
C436 VTAIL.n25 B 0.020025f
C437 VTAIL.n26 B 0.010761f
C438 VTAIL.n27 B 0.025434f
C439 VTAIL.n28 B 0.011394f
C440 VTAIL.n29 B 1.53047f
C441 VTAIL.n30 B 0.010761f
C442 VTAIL.t0 B 0.042109f
C443 VTAIL.n31 B 0.14306f
C444 VTAIL.n32 B 0.015025f
C445 VTAIL.n33 B 0.019076f
C446 VTAIL.n34 B 0.025434f
C447 VTAIL.n35 B 0.011394f
C448 VTAIL.n36 B 0.010761f
C449 VTAIL.n37 B 0.020025f
C450 VTAIL.n38 B 0.020025f
C451 VTAIL.n39 B 0.010761f
C452 VTAIL.n40 B 0.011394f
C453 VTAIL.n41 B 0.025434f
C454 VTAIL.n42 B 0.025434f
C455 VTAIL.n43 B 0.011394f
C456 VTAIL.n44 B 0.010761f
C457 VTAIL.n45 B 0.020025f
C458 VTAIL.n46 B 0.020025f
C459 VTAIL.n47 B 0.010761f
C460 VTAIL.n48 B 0.011394f
C461 VTAIL.n49 B 0.025434f
C462 VTAIL.n50 B 0.025434f
C463 VTAIL.n51 B 0.011394f
C464 VTAIL.n52 B 0.010761f
C465 VTAIL.n53 B 0.020025f
C466 VTAIL.n54 B 0.020025f
C467 VTAIL.n55 B 0.010761f
C468 VTAIL.n56 B 0.011394f
C469 VTAIL.n57 B 0.025434f
C470 VTAIL.n58 B 0.025434f
C471 VTAIL.n59 B 0.011394f
C472 VTAIL.n60 B 0.010761f
C473 VTAIL.n61 B 0.020025f
C474 VTAIL.n62 B 0.020025f
C475 VTAIL.n63 B 0.010761f
C476 VTAIL.n64 B 0.011394f
C477 VTAIL.n65 B 0.025434f
C478 VTAIL.n66 B 0.025434f
C479 VTAIL.n67 B 0.011394f
C480 VTAIL.n68 B 0.010761f
C481 VTAIL.n69 B 0.020025f
C482 VTAIL.n70 B 0.020025f
C483 VTAIL.n71 B 0.010761f
C484 VTAIL.n72 B 0.010761f
C485 VTAIL.n73 B 0.011394f
C486 VTAIL.n74 B 0.025434f
C487 VTAIL.n75 B 0.025434f
C488 VTAIL.n76 B 0.025434f
C489 VTAIL.n77 B 0.011077f
C490 VTAIL.n78 B 0.010761f
C491 VTAIL.n79 B 0.020025f
C492 VTAIL.n80 B 0.020025f
C493 VTAIL.n81 B 0.010761f
C494 VTAIL.n82 B 0.011394f
C495 VTAIL.n83 B 0.025434f
C496 VTAIL.n84 B 0.025434f
C497 VTAIL.n85 B 0.011394f
C498 VTAIL.n86 B 0.010761f
C499 VTAIL.n87 B 0.020025f
C500 VTAIL.n88 B 0.020025f
C501 VTAIL.n89 B 0.010761f
C502 VTAIL.n90 B 0.011394f
C503 VTAIL.n91 B 0.025434f
C504 VTAIL.n92 B 0.05315f
C505 VTAIL.n93 B 0.011394f
C506 VTAIL.n94 B 0.010761f
C507 VTAIL.n95 B 0.045193f
C508 VTAIL.n96 B 0.029509f
C509 VTAIL.n97 B 1.45247f
C510 VTAIL.n98 B 0.027066f
C511 VTAIL.n99 B 0.020025f
C512 VTAIL.n100 B 0.010761f
C513 VTAIL.n101 B 0.025434f
C514 VTAIL.n102 B 0.011394f
C515 VTAIL.n103 B 0.020025f
C516 VTAIL.n104 B 0.010761f
C517 VTAIL.n105 B 0.025434f
C518 VTAIL.n106 B 0.011077f
C519 VTAIL.n107 B 0.020025f
C520 VTAIL.n108 B 0.011077f
C521 VTAIL.n109 B 0.010761f
C522 VTAIL.n110 B 0.025434f
C523 VTAIL.n111 B 0.025434f
C524 VTAIL.n112 B 0.011394f
C525 VTAIL.n113 B 0.020025f
C526 VTAIL.n114 B 0.010761f
C527 VTAIL.n115 B 0.025434f
C528 VTAIL.n116 B 0.011394f
C529 VTAIL.n117 B 0.020025f
C530 VTAIL.n118 B 0.010761f
C531 VTAIL.n119 B 0.025434f
C532 VTAIL.n120 B 0.011394f
C533 VTAIL.n121 B 0.020025f
C534 VTAIL.n122 B 0.010761f
C535 VTAIL.n123 B 0.025434f
C536 VTAIL.n124 B 0.011394f
C537 VTAIL.n125 B 0.020025f
C538 VTAIL.n126 B 0.010761f
C539 VTAIL.n127 B 0.025434f
C540 VTAIL.n128 B 0.011394f
C541 VTAIL.n129 B 1.53047f
C542 VTAIL.n130 B 0.010761f
C543 VTAIL.t2 B 0.042109f
C544 VTAIL.n131 B 0.14306f
C545 VTAIL.n132 B 0.015025f
C546 VTAIL.n133 B 0.019076f
C547 VTAIL.n134 B 0.025434f
C548 VTAIL.n135 B 0.011394f
C549 VTAIL.n136 B 0.010761f
C550 VTAIL.n137 B 0.020025f
C551 VTAIL.n138 B 0.020025f
C552 VTAIL.n139 B 0.010761f
C553 VTAIL.n140 B 0.011394f
C554 VTAIL.n141 B 0.025434f
C555 VTAIL.n142 B 0.025434f
C556 VTAIL.n143 B 0.011394f
C557 VTAIL.n144 B 0.010761f
C558 VTAIL.n145 B 0.020025f
C559 VTAIL.n146 B 0.020025f
C560 VTAIL.n147 B 0.010761f
C561 VTAIL.n148 B 0.011394f
C562 VTAIL.n149 B 0.025434f
C563 VTAIL.n150 B 0.025434f
C564 VTAIL.n151 B 0.011394f
C565 VTAIL.n152 B 0.010761f
C566 VTAIL.n153 B 0.020025f
C567 VTAIL.n154 B 0.020025f
C568 VTAIL.n155 B 0.010761f
C569 VTAIL.n156 B 0.011394f
C570 VTAIL.n157 B 0.025434f
C571 VTAIL.n158 B 0.025434f
C572 VTAIL.n159 B 0.011394f
C573 VTAIL.n160 B 0.010761f
C574 VTAIL.n161 B 0.020025f
C575 VTAIL.n162 B 0.020025f
C576 VTAIL.n163 B 0.010761f
C577 VTAIL.n164 B 0.011394f
C578 VTAIL.n165 B 0.025434f
C579 VTAIL.n166 B 0.025434f
C580 VTAIL.n167 B 0.011394f
C581 VTAIL.n168 B 0.010761f
C582 VTAIL.n169 B 0.020025f
C583 VTAIL.n170 B 0.020025f
C584 VTAIL.n171 B 0.010761f
C585 VTAIL.n172 B 0.011394f
C586 VTAIL.n173 B 0.025434f
C587 VTAIL.n174 B 0.025434f
C588 VTAIL.n175 B 0.011394f
C589 VTAIL.n176 B 0.010761f
C590 VTAIL.n177 B 0.020025f
C591 VTAIL.n178 B 0.020025f
C592 VTAIL.n179 B 0.010761f
C593 VTAIL.n180 B 0.011394f
C594 VTAIL.n181 B 0.025434f
C595 VTAIL.n182 B 0.025434f
C596 VTAIL.n183 B 0.011394f
C597 VTAIL.n184 B 0.010761f
C598 VTAIL.n185 B 0.020025f
C599 VTAIL.n186 B 0.020025f
C600 VTAIL.n187 B 0.010761f
C601 VTAIL.n188 B 0.011394f
C602 VTAIL.n189 B 0.025434f
C603 VTAIL.n190 B 0.05315f
C604 VTAIL.n191 B 0.011394f
C605 VTAIL.n192 B 0.010761f
C606 VTAIL.n193 B 0.045193f
C607 VTAIL.n194 B 0.029509f
C608 VTAIL.n195 B 1.4661f
C609 VTAIL.n196 B 0.027066f
C610 VTAIL.n197 B 0.020025f
C611 VTAIL.n198 B 0.010761f
C612 VTAIL.n199 B 0.025434f
C613 VTAIL.n200 B 0.011394f
C614 VTAIL.n201 B 0.020025f
C615 VTAIL.n202 B 0.010761f
C616 VTAIL.n203 B 0.025434f
C617 VTAIL.n204 B 0.011077f
C618 VTAIL.n205 B 0.020025f
C619 VTAIL.n206 B 0.011077f
C620 VTAIL.n207 B 0.010761f
C621 VTAIL.n208 B 0.025434f
C622 VTAIL.n209 B 0.025434f
C623 VTAIL.n210 B 0.011394f
C624 VTAIL.n211 B 0.020025f
C625 VTAIL.n212 B 0.010761f
C626 VTAIL.n213 B 0.025434f
C627 VTAIL.n214 B 0.011394f
C628 VTAIL.n215 B 0.020025f
C629 VTAIL.n216 B 0.010761f
C630 VTAIL.n217 B 0.025434f
C631 VTAIL.n218 B 0.011394f
C632 VTAIL.n219 B 0.020025f
C633 VTAIL.n220 B 0.010761f
C634 VTAIL.n221 B 0.025434f
C635 VTAIL.n222 B 0.011394f
C636 VTAIL.n223 B 0.020025f
C637 VTAIL.n224 B 0.010761f
C638 VTAIL.n225 B 0.025434f
C639 VTAIL.n226 B 0.011394f
C640 VTAIL.n227 B 1.53047f
C641 VTAIL.n228 B 0.010761f
C642 VTAIL.t3 B 0.042109f
C643 VTAIL.n229 B 0.14306f
C644 VTAIL.n230 B 0.015025f
C645 VTAIL.n231 B 0.019076f
C646 VTAIL.n232 B 0.025434f
C647 VTAIL.n233 B 0.011394f
C648 VTAIL.n234 B 0.010761f
C649 VTAIL.n235 B 0.020025f
C650 VTAIL.n236 B 0.020025f
C651 VTAIL.n237 B 0.010761f
C652 VTAIL.n238 B 0.011394f
C653 VTAIL.n239 B 0.025434f
C654 VTAIL.n240 B 0.025434f
C655 VTAIL.n241 B 0.011394f
C656 VTAIL.n242 B 0.010761f
C657 VTAIL.n243 B 0.020025f
C658 VTAIL.n244 B 0.020025f
C659 VTAIL.n245 B 0.010761f
C660 VTAIL.n246 B 0.011394f
C661 VTAIL.n247 B 0.025434f
C662 VTAIL.n248 B 0.025434f
C663 VTAIL.n249 B 0.011394f
C664 VTAIL.n250 B 0.010761f
C665 VTAIL.n251 B 0.020025f
C666 VTAIL.n252 B 0.020025f
C667 VTAIL.n253 B 0.010761f
C668 VTAIL.n254 B 0.011394f
C669 VTAIL.n255 B 0.025434f
C670 VTAIL.n256 B 0.025434f
C671 VTAIL.n257 B 0.011394f
C672 VTAIL.n258 B 0.010761f
C673 VTAIL.n259 B 0.020025f
C674 VTAIL.n260 B 0.020025f
C675 VTAIL.n261 B 0.010761f
C676 VTAIL.n262 B 0.011394f
C677 VTAIL.n263 B 0.025434f
C678 VTAIL.n264 B 0.025434f
C679 VTAIL.n265 B 0.011394f
C680 VTAIL.n266 B 0.010761f
C681 VTAIL.n267 B 0.020025f
C682 VTAIL.n268 B 0.020025f
C683 VTAIL.n269 B 0.010761f
C684 VTAIL.n270 B 0.011394f
C685 VTAIL.n271 B 0.025434f
C686 VTAIL.n272 B 0.025434f
C687 VTAIL.n273 B 0.011394f
C688 VTAIL.n274 B 0.010761f
C689 VTAIL.n275 B 0.020025f
C690 VTAIL.n276 B 0.020025f
C691 VTAIL.n277 B 0.010761f
C692 VTAIL.n278 B 0.011394f
C693 VTAIL.n279 B 0.025434f
C694 VTAIL.n280 B 0.025434f
C695 VTAIL.n281 B 0.011394f
C696 VTAIL.n282 B 0.010761f
C697 VTAIL.n283 B 0.020025f
C698 VTAIL.n284 B 0.020025f
C699 VTAIL.n285 B 0.010761f
C700 VTAIL.n286 B 0.011394f
C701 VTAIL.n287 B 0.025434f
C702 VTAIL.n288 B 0.05315f
C703 VTAIL.n289 B 0.011394f
C704 VTAIL.n290 B 0.010761f
C705 VTAIL.n291 B 0.045193f
C706 VTAIL.n292 B 0.029509f
C707 VTAIL.n293 B 1.39657f
C708 VTAIL.n294 B 0.027066f
C709 VTAIL.n295 B 0.020025f
C710 VTAIL.n296 B 0.010761f
C711 VTAIL.n297 B 0.025434f
C712 VTAIL.n298 B 0.011394f
C713 VTAIL.n299 B 0.020025f
C714 VTAIL.n300 B 0.010761f
C715 VTAIL.n301 B 0.025434f
C716 VTAIL.n302 B 0.011077f
C717 VTAIL.n303 B 0.020025f
C718 VTAIL.n304 B 0.011394f
C719 VTAIL.n305 B 0.025434f
C720 VTAIL.n306 B 0.011394f
C721 VTAIL.n307 B 0.020025f
C722 VTAIL.n308 B 0.010761f
C723 VTAIL.n309 B 0.025434f
C724 VTAIL.n310 B 0.011394f
C725 VTAIL.n311 B 0.020025f
C726 VTAIL.n312 B 0.010761f
C727 VTAIL.n313 B 0.025434f
C728 VTAIL.n314 B 0.011394f
C729 VTAIL.n315 B 0.020025f
C730 VTAIL.n316 B 0.010761f
C731 VTAIL.n317 B 0.025434f
C732 VTAIL.n318 B 0.011394f
C733 VTAIL.n319 B 0.020025f
C734 VTAIL.n320 B 0.010761f
C735 VTAIL.n321 B 0.025434f
C736 VTAIL.n322 B 0.011394f
C737 VTAIL.n323 B 1.53047f
C738 VTAIL.n324 B 0.010761f
C739 VTAIL.t1 B 0.042109f
C740 VTAIL.n325 B 0.14306f
C741 VTAIL.n326 B 0.015025f
C742 VTAIL.n327 B 0.019076f
C743 VTAIL.n328 B 0.025434f
C744 VTAIL.n329 B 0.011394f
C745 VTAIL.n330 B 0.010761f
C746 VTAIL.n331 B 0.020025f
C747 VTAIL.n332 B 0.020025f
C748 VTAIL.n333 B 0.010761f
C749 VTAIL.n334 B 0.011394f
C750 VTAIL.n335 B 0.025434f
C751 VTAIL.n336 B 0.025434f
C752 VTAIL.n337 B 0.011394f
C753 VTAIL.n338 B 0.010761f
C754 VTAIL.n339 B 0.020025f
C755 VTAIL.n340 B 0.020025f
C756 VTAIL.n341 B 0.010761f
C757 VTAIL.n342 B 0.011394f
C758 VTAIL.n343 B 0.025434f
C759 VTAIL.n344 B 0.025434f
C760 VTAIL.n345 B 0.011394f
C761 VTAIL.n346 B 0.010761f
C762 VTAIL.n347 B 0.020025f
C763 VTAIL.n348 B 0.020025f
C764 VTAIL.n349 B 0.010761f
C765 VTAIL.n350 B 0.011394f
C766 VTAIL.n351 B 0.025434f
C767 VTAIL.n352 B 0.025434f
C768 VTAIL.n353 B 0.011394f
C769 VTAIL.n354 B 0.010761f
C770 VTAIL.n355 B 0.020025f
C771 VTAIL.n356 B 0.020025f
C772 VTAIL.n357 B 0.010761f
C773 VTAIL.n358 B 0.011394f
C774 VTAIL.n359 B 0.025434f
C775 VTAIL.n360 B 0.025434f
C776 VTAIL.n361 B 0.011394f
C777 VTAIL.n362 B 0.010761f
C778 VTAIL.n363 B 0.020025f
C779 VTAIL.n364 B 0.020025f
C780 VTAIL.n365 B 0.010761f
C781 VTAIL.n366 B 0.010761f
C782 VTAIL.n367 B 0.011394f
C783 VTAIL.n368 B 0.025434f
C784 VTAIL.n369 B 0.025434f
C785 VTAIL.n370 B 0.025434f
C786 VTAIL.n371 B 0.011077f
C787 VTAIL.n372 B 0.010761f
C788 VTAIL.n373 B 0.020025f
C789 VTAIL.n374 B 0.020025f
C790 VTAIL.n375 B 0.010761f
C791 VTAIL.n376 B 0.011394f
C792 VTAIL.n377 B 0.025434f
C793 VTAIL.n378 B 0.025434f
C794 VTAIL.n379 B 0.011394f
C795 VTAIL.n380 B 0.010761f
C796 VTAIL.n381 B 0.020025f
C797 VTAIL.n382 B 0.020025f
C798 VTAIL.n383 B 0.010761f
C799 VTAIL.n384 B 0.011394f
C800 VTAIL.n385 B 0.025434f
C801 VTAIL.n386 B 0.05315f
C802 VTAIL.n387 B 0.011394f
C803 VTAIL.n388 B 0.010761f
C804 VTAIL.n389 B 0.045193f
C805 VTAIL.n390 B 0.029509f
C806 VTAIL.n391 B 1.34511f
C807 VN.t1 B 2.55293f
C808 VN.t0 B 2.74434f
.ends

