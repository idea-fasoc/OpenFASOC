* NGSPICE file created from diff_pair_sample_0519.ext - technology: sky130A

.subckt diff_pair_sample_0519 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t9 VN.t0 VTAIL.t10 w_n4066_n4000# sky130_fd_pr__pfet_01v8 ad=2.5014 pd=15.49 as=2.5014 ps=15.49 w=15.16 l=2.25
X1 VDD2.t8 VN.t1 VTAIL.t11 w_n4066_n4000# sky130_fd_pr__pfet_01v8 ad=5.9124 pd=31.1 as=2.5014 ps=15.49 w=15.16 l=2.25
X2 B.t11 B.t9 B.t10 w_n4066_n4000# sky130_fd_pr__pfet_01v8 ad=5.9124 pd=31.1 as=0 ps=0 w=15.16 l=2.25
X3 B.t8 B.t6 B.t7 w_n4066_n4000# sky130_fd_pr__pfet_01v8 ad=5.9124 pd=31.1 as=0 ps=0 w=15.16 l=2.25
X4 VDD2.t7 VN.t2 VTAIL.t12 w_n4066_n4000# sky130_fd_pr__pfet_01v8 ad=2.5014 pd=15.49 as=2.5014 ps=15.49 w=15.16 l=2.25
X5 VTAIL.t5 VP.t0 VDD1.t9 w_n4066_n4000# sky130_fd_pr__pfet_01v8 ad=2.5014 pd=15.49 as=2.5014 ps=15.49 w=15.16 l=2.25
X6 VTAIL.t4 VP.t1 VDD1.t8 w_n4066_n4000# sky130_fd_pr__pfet_01v8 ad=2.5014 pd=15.49 as=2.5014 ps=15.49 w=15.16 l=2.25
X7 VTAIL.t13 VN.t3 VDD2.t6 w_n4066_n4000# sky130_fd_pr__pfet_01v8 ad=2.5014 pd=15.49 as=2.5014 ps=15.49 w=15.16 l=2.25
X8 VDD1.t7 VP.t2 VTAIL.t16 w_n4066_n4000# sky130_fd_pr__pfet_01v8 ad=2.5014 pd=15.49 as=5.9124 ps=31.1 w=15.16 l=2.25
X9 VDD2.t5 VN.t4 VTAIL.t15 w_n4066_n4000# sky130_fd_pr__pfet_01v8 ad=2.5014 pd=15.49 as=5.9124 ps=31.1 w=15.16 l=2.25
X10 B.t5 B.t3 B.t4 w_n4066_n4000# sky130_fd_pr__pfet_01v8 ad=5.9124 pd=31.1 as=0 ps=0 w=15.16 l=2.25
X11 B.t2 B.t0 B.t1 w_n4066_n4000# sky130_fd_pr__pfet_01v8 ad=5.9124 pd=31.1 as=0 ps=0 w=15.16 l=2.25
X12 VTAIL.t14 VN.t5 VDD2.t4 w_n4066_n4000# sky130_fd_pr__pfet_01v8 ad=2.5014 pd=15.49 as=2.5014 ps=15.49 w=15.16 l=2.25
X13 VDD1.t6 VP.t3 VTAIL.t3 w_n4066_n4000# sky130_fd_pr__pfet_01v8 ad=2.5014 pd=15.49 as=2.5014 ps=15.49 w=15.16 l=2.25
X14 VTAIL.t0 VP.t4 VDD1.t5 w_n4066_n4000# sky130_fd_pr__pfet_01v8 ad=2.5014 pd=15.49 as=2.5014 ps=15.49 w=15.16 l=2.25
X15 VDD2.t3 VN.t6 VTAIL.t9 w_n4066_n4000# sky130_fd_pr__pfet_01v8 ad=5.9124 pd=31.1 as=2.5014 ps=15.49 w=15.16 l=2.25
X16 VTAIL.t6 VN.t7 VDD2.t2 w_n4066_n4000# sky130_fd_pr__pfet_01v8 ad=2.5014 pd=15.49 as=2.5014 ps=15.49 w=15.16 l=2.25
X17 VDD2.t1 VN.t8 VTAIL.t7 w_n4066_n4000# sky130_fd_pr__pfet_01v8 ad=2.5014 pd=15.49 as=5.9124 ps=31.1 w=15.16 l=2.25
X18 VDD1.t4 VP.t5 VTAIL.t2 w_n4066_n4000# sky130_fd_pr__pfet_01v8 ad=5.9124 pd=31.1 as=2.5014 ps=15.49 w=15.16 l=2.25
X19 VTAIL.t1 VP.t6 VDD1.t3 w_n4066_n4000# sky130_fd_pr__pfet_01v8 ad=2.5014 pd=15.49 as=2.5014 ps=15.49 w=15.16 l=2.25
X20 VTAIL.t8 VN.t9 VDD2.t0 w_n4066_n4000# sky130_fd_pr__pfet_01v8 ad=2.5014 pd=15.49 as=2.5014 ps=15.49 w=15.16 l=2.25
X21 VDD1.t2 VP.t7 VTAIL.t17 w_n4066_n4000# sky130_fd_pr__pfet_01v8 ad=2.5014 pd=15.49 as=2.5014 ps=15.49 w=15.16 l=2.25
X22 VDD1.t1 VP.t8 VTAIL.t19 w_n4066_n4000# sky130_fd_pr__pfet_01v8 ad=5.9124 pd=31.1 as=2.5014 ps=15.49 w=15.16 l=2.25
X23 VDD1.t0 VP.t9 VTAIL.t18 w_n4066_n4000# sky130_fd_pr__pfet_01v8 ad=2.5014 pd=15.49 as=5.9124 ps=31.1 w=15.16 l=2.25
R0 VN.n8 VN.t1 196.519
R1 VN.n44 VN.t4 196.519
R2 VN.n9 VN.t9 162.381
R3 VN.n5 VN.t2 162.381
R4 VN.n26 VN.t5 162.381
R5 VN.n34 VN.t8 162.381
R6 VN.n45 VN.t7 162.381
R7 VN.n41 VN.t0 162.381
R8 VN.n62 VN.t3 162.381
R9 VN.n70 VN.t6 162.381
R10 VN.n69 VN.n36 161.3
R11 VN.n68 VN.n67 161.3
R12 VN.n66 VN.n37 161.3
R13 VN.n65 VN.n64 161.3
R14 VN.n63 VN.n38 161.3
R15 VN.n61 VN.n60 161.3
R16 VN.n59 VN.n39 161.3
R17 VN.n58 VN.n57 161.3
R18 VN.n56 VN.n40 161.3
R19 VN.n55 VN.n54 161.3
R20 VN.n53 VN.n52 161.3
R21 VN.n51 VN.n42 161.3
R22 VN.n50 VN.n49 161.3
R23 VN.n48 VN.n43 161.3
R24 VN.n47 VN.n46 161.3
R25 VN.n33 VN.n0 161.3
R26 VN.n32 VN.n31 161.3
R27 VN.n30 VN.n1 161.3
R28 VN.n29 VN.n28 161.3
R29 VN.n27 VN.n2 161.3
R30 VN.n25 VN.n24 161.3
R31 VN.n23 VN.n3 161.3
R32 VN.n22 VN.n21 161.3
R33 VN.n20 VN.n4 161.3
R34 VN.n19 VN.n18 161.3
R35 VN.n17 VN.n16 161.3
R36 VN.n15 VN.n6 161.3
R37 VN.n14 VN.n13 161.3
R38 VN.n12 VN.n7 161.3
R39 VN.n11 VN.n10 161.3
R40 VN.n35 VN.n34 90.7429
R41 VN.n71 VN.n70 90.7429
R42 VN.n9 VN.n8 55.0386
R43 VN.n45 VN.n44 55.0386
R44 VN VN.n71 53.9755
R45 VN.n32 VN.n1 52.2023
R46 VN.n68 VN.n37 52.2023
R47 VN.n14 VN.n7 44.4521
R48 VN.n21 VN.n3 44.4521
R49 VN.n50 VN.n43 44.4521
R50 VN.n57 VN.n39 44.4521
R51 VN.n15 VN.n14 36.702
R52 VN.n21 VN.n20 36.702
R53 VN.n51 VN.n50 36.702
R54 VN.n57 VN.n56 36.702
R55 VN.n28 VN.n1 28.9518
R56 VN.n64 VN.n37 28.9518
R57 VN.n10 VN.n7 24.5923
R58 VN.n16 VN.n15 24.5923
R59 VN.n20 VN.n19 24.5923
R60 VN.n25 VN.n3 24.5923
R61 VN.n28 VN.n27 24.5923
R62 VN.n33 VN.n32 24.5923
R63 VN.n46 VN.n43 24.5923
R64 VN.n56 VN.n55 24.5923
R65 VN.n52 VN.n51 24.5923
R66 VN.n64 VN.n63 24.5923
R67 VN.n61 VN.n39 24.5923
R68 VN.n69 VN.n68 24.5923
R69 VN.n34 VN.n33 20.1658
R70 VN.n70 VN.n69 20.1658
R71 VN.n10 VN.n9 16.2311
R72 VN.n26 VN.n25 16.2311
R73 VN.n46 VN.n45 16.2311
R74 VN.n62 VN.n61 16.2311
R75 VN.n16 VN.n5 12.2964
R76 VN.n19 VN.n5 12.2964
R77 VN.n55 VN.n41 12.2964
R78 VN.n52 VN.n41 12.2964
R79 VN.n47 VN.n44 8.94118
R80 VN.n11 VN.n8 8.94118
R81 VN.n27 VN.n26 8.36172
R82 VN.n63 VN.n62 8.36172
R83 VN.n71 VN.n36 0.278335
R84 VN.n35 VN.n0 0.278335
R85 VN.n67 VN.n36 0.189894
R86 VN.n67 VN.n66 0.189894
R87 VN.n66 VN.n65 0.189894
R88 VN.n65 VN.n38 0.189894
R89 VN.n60 VN.n38 0.189894
R90 VN.n60 VN.n59 0.189894
R91 VN.n59 VN.n58 0.189894
R92 VN.n58 VN.n40 0.189894
R93 VN.n54 VN.n40 0.189894
R94 VN.n54 VN.n53 0.189894
R95 VN.n53 VN.n42 0.189894
R96 VN.n49 VN.n42 0.189894
R97 VN.n49 VN.n48 0.189894
R98 VN.n48 VN.n47 0.189894
R99 VN.n12 VN.n11 0.189894
R100 VN.n13 VN.n12 0.189894
R101 VN.n13 VN.n6 0.189894
R102 VN.n17 VN.n6 0.189894
R103 VN.n18 VN.n17 0.189894
R104 VN.n18 VN.n4 0.189894
R105 VN.n22 VN.n4 0.189894
R106 VN.n23 VN.n22 0.189894
R107 VN.n24 VN.n23 0.189894
R108 VN.n24 VN.n2 0.189894
R109 VN.n29 VN.n2 0.189894
R110 VN.n30 VN.n29 0.189894
R111 VN.n31 VN.n30 0.189894
R112 VN.n31 VN.n0 0.189894
R113 VN VN.n35 0.153485
R114 VTAIL.n11 VTAIL.t15 59.0735
R115 VTAIL.n17 VTAIL.t7 59.0733
R116 VTAIL.n2 VTAIL.t16 59.0733
R117 VTAIL.n16 VTAIL.t18 59.0733
R118 VTAIL.n15 VTAIL.n14 56.9294
R119 VTAIL.n13 VTAIL.n12 56.9294
R120 VTAIL.n10 VTAIL.n9 56.9294
R121 VTAIL.n8 VTAIL.n7 56.9294
R122 VTAIL.n19 VTAIL.n18 56.9291
R123 VTAIL.n1 VTAIL.n0 56.9291
R124 VTAIL.n4 VTAIL.n3 56.9291
R125 VTAIL.n6 VTAIL.n5 56.9291
R126 VTAIL.n8 VTAIL.n6 29.8841
R127 VTAIL.n17 VTAIL.n16 27.66
R128 VTAIL.n10 VTAIL.n8 2.22464
R129 VTAIL.n11 VTAIL.n10 2.22464
R130 VTAIL.n15 VTAIL.n13 2.22464
R131 VTAIL.n16 VTAIL.n15 2.22464
R132 VTAIL.n6 VTAIL.n4 2.22464
R133 VTAIL.n4 VTAIL.n2 2.22464
R134 VTAIL.n19 VTAIL.n17 2.22464
R135 VTAIL.n18 VTAIL.t12 2.14463
R136 VTAIL.n18 VTAIL.t14 2.14463
R137 VTAIL.n0 VTAIL.t11 2.14463
R138 VTAIL.n0 VTAIL.t8 2.14463
R139 VTAIL.n3 VTAIL.t17 2.14463
R140 VTAIL.n3 VTAIL.t1 2.14463
R141 VTAIL.n5 VTAIL.t19 2.14463
R142 VTAIL.n5 VTAIL.t5 2.14463
R143 VTAIL.n14 VTAIL.t3 2.14463
R144 VTAIL.n14 VTAIL.t0 2.14463
R145 VTAIL.n12 VTAIL.t2 2.14463
R146 VTAIL.n12 VTAIL.t4 2.14463
R147 VTAIL.n9 VTAIL.t10 2.14463
R148 VTAIL.n9 VTAIL.t6 2.14463
R149 VTAIL.n7 VTAIL.t9 2.14463
R150 VTAIL.n7 VTAIL.t13 2.14463
R151 VTAIL VTAIL.n1 1.72679
R152 VTAIL.n13 VTAIL.n11 1.5824
R153 VTAIL.n2 VTAIL.n1 1.5824
R154 VTAIL VTAIL.n19 0.498345
R155 VDD2.n1 VDD2.t8 77.9762
R156 VDD2.n4 VDD2.t3 75.7523
R157 VDD2.n3 VDD2.n2 75.2207
R158 VDD2 VDD2.n7 75.2179
R159 VDD2.n6 VDD2.n5 73.6082
R160 VDD2.n1 VDD2.n0 73.6079
R161 VDD2.n4 VDD2.n3 47.3489
R162 VDD2.n6 VDD2.n4 2.22464
R163 VDD2.n7 VDD2.t2 2.14463
R164 VDD2.n7 VDD2.t5 2.14463
R165 VDD2.n5 VDD2.t6 2.14463
R166 VDD2.n5 VDD2.t9 2.14463
R167 VDD2.n2 VDD2.t4 2.14463
R168 VDD2.n2 VDD2.t1 2.14463
R169 VDD2.n0 VDD2.t0 2.14463
R170 VDD2.n0 VDD2.t7 2.14463
R171 VDD2 VDD2.n6 0.614724
R172 VDD2.n3 VDD2.n1 0.501188
R173 B.n474 B.n473 585
R174 B.n472 B.n143 585
R175 B.n471 B.n470 585
R176 B.n469 B.n144 585
R177 B.n468 B.n467 585
R178 B.n466 B.n145 585
R179 B.n465 B.n464 585
R180 B.n463 B.n146 585
R181 B.n462 B.n461 585
R182 B.n460 B.n147 585
R183 B.n459 B.n458 585
R184 B.n457 B.n148 585
R185 B.n456 B.n455 585
R186 B.n454 B.n149 585
R187 B.n453 B.n452 585
R188 B.n451 B.n150 585
R189 B.n450 B.n449 585
R190 B.n448 B.n151 585
R191 B.n447 B.n446 585
R192 B.n445 B.n152 585
R193 B.n444 B.n443 585
R194 B.n442 B.n153 585
R195 B.n441 B.n440 585
R196 B.n439 B.n154 585
R197 B.n438 B.n437 585
R198 B.n436 B.n155 585
R199 B.n435 B.n434 585
R200 B.n433 B.n156 585
R201 B.n432 B.n431 585
R202 B.n430 B.n157 585
R203 B.n429 B.n428 585
R204 B.n427 B.n158 585
R205 B.n426 B.n425 585
R206 B.n424 B.n159 585
R207 B.n423 B.n422 585
R208 B.n421 B.n160 585
R209 B.n420 B.n419 585
R210 B.n418 B.n161 585
R211 B.n417 B.n416 585
R212 B.n415 B.n162 585
R213 B.n414 B.n413 585
R214 B.n412 B.n163 585
R215 B.n411 B.n410 585
R216 B.n409 B.n164 585
R217 B.n408 B.n407 585
R218 B.n406 B.n165 585
R219 B.n405 B.n404 585
R220 B.n403 B.n166 585
R221 B.n402 B.n401 585
R222 B.n400 B.n167 585
R223 B.n399 B.n398 585
R224 B.n397 B.n396 585
R225 B.n395 B.n171 585
R226 B.n394 B.n393 585
R227 B.n392 B.n172 585
R228 B.n391 B.n390 585
R229 B.n389 B.n173 585
R230 B.n388 B.n387 585
R231 B.n386 B.n174 585
R232 B.n385 B.n384 585
R233 B.n382 B.n175 585
R234 B.n381 B.n380 585
R235 B.n379 B.n178 585
R236 B.n378 B.n377 585
R237 B.n376 B.n179 585
R238 B.n375 B.n374 585
R239 B.n373 B.n180 585
R240 B.n372 B.n371 585
R241 B.n370 B.n181 585
R242 B.n369 B.n368 585
R243 B.n367 B.n182 585
R244 B.n366 B.n365 585
R245 B.n364 B.n183 585
R246 B.n363 B.n362 585
R247 B.n361 B.n184 585
R248 B.n360 B.n359 585
R249 B.n358 B.n185 585
R250 B.n357 B.n356 585
R251 B.n355 B.n186 585
R252 B.n354 B.n353 585
R253 B.n352 B.n187 585
R254 B.n351 B.n350 585
R255 B.n349 B.n188 585
R256 B.n348 B.n347 585
R257 B.n346 B.n189 585
R258 B.n345 B.n344 585
R259 B.n343 B.n190 585
R260 B.n342 B.n341 585
R261 B.n340 B.n191 585
R262 B.n339 B.n338 585
R263 B.n337 B.n192 585
R264 B.n336 B.n335 585
R265 B.n334 B.n193 585
R266 B.n333 B.n332 585
R267 B.n331 B.n194 585
R268 B.n330 B.n329 585
R269 B.n328 B.n195 585
R270 B.n327 B.n326 585
R271 B.n325 B.n196 585
R272 B.n324 B.n323 585
R273 B.n322 B.n197 585
R274 B.n321 B.n320 585
R275 B.n319 B.n198 585
R276 B.n318 B.n317 585
R277 B.n316 B.n199 585
R278 B.n315 B.n314 585
R279 B.n313 B.n200 585
R280 B.n312 B.n311 585
R281 B.n310 B.n201 585
R282 B.n309 B.n308 585
R283 B.n307 B.n202 585
R284 B.n475 B.n142 585
R285 B.n477 B.n476 585
R286 B.n478 B.n141 585
R287 B.n480 B.n479 585
R288 B.n481 B.n140 585
R289 B.n483 B.n482 585
R290 B.n484 B.n139 585
R291 B.n486 B.n485 585
R292 B.n487 B.n138 585
R293 B.n489 B.n488 585
R294 B.n490 B.n137 585
R295 B.n492 B.n491 585
R296 B.n493 B.n136 585
R297 B.n495 B.n494 585
R298 B.n496 B.n135 585
R299 B.n498 B.n497 585
R300 B.n499 B.n134 585
R301 B.n501 B.n500 585
R302 B.n502 B.n133 585
R303 B.n504 B.n503 585
R304 B.n505 B.n132 585
R305 B.n507 B.n506 585
R306 B.n508 B.n131 585
R307 B.n510 B.n509 585
R308 B.n511 B.n130 585
R309 B.n513 B.n512 585
R310 B.n514 B.n129 585
R311 B.n516 B.n515 585
R312 B.n517 B.n128 585
R313 B.n519 B.n518 585
R314 B.n520 B.n127 585
R315 B.n522 B.n521 585
R316 B.n523 B.n126 585
R317 B.n525 B.n524 585
R318 B.n526 B.n125 585
R319 B.n528 B.n527 585
R320 B.n529 B.n124 585
R321 B.n531 B.n530 585
R322 B.n532 B.n123 585
R323 B.n534 B.n533 585
R324 B.n535 B.n122 585
R325 B.n537 B.n536 585
R326 B.n538 B.n121 585
R327 B.n540 B.n539 585
R328 B.n541 B.n120 585
R329 B.n543 B.n542 585
R330 B.n544 B.n119 585
R331 B.n546 B.n545 585
R332 B.n547 B.n118 585
R333 B.n549 B.n548 585
R334 B.n550 B.n117 585
R335 B.n552 B.n551 585
R336 B.n553 B.n116 585
R337 B.n555 B.n554 585
R338 B.n556 B.n115 585
R339 B.n558 B.n557 585
R340 B.n559 B.n114 585
R341 B.n561 B.n560 585
R342 B.n562 B.n113 585
R343 B.n564 B.n563 585
R344 B.n565 B.n112 585
R345 B.n567 B.n566 585
R346 B.n568 B.n111 585
R347 B.n570 B.n569 585
R348 B.n571 B.n110 585
R349 B.n573 B.n572 585
R350 B.n574 B.n109 585
R351 B.n576 B.n575 585
R352 B.n577 B.n108 585
R353 B.n579 B.n578 585
R354 B.n580 B.n107 585
R355 B.n582 B.n581 585
R356 B.n583 B.n106 585
R357 B.n585 B.n584 585
R358 B.n586 B.n105 585
R359 B.n588 B.n587 585
R360 B.n589 B.n104 585
R361 B.n591 B.n590 585
R362 B.n592 B.n103 585
R363 B.n594 B.n593 585
R364 B.n595 B.n102 585
R365 B.n597 B.n596 585
R366 B.n598 B.n101 585
R367 B.n600 B.n599 585
R368 B.n601 B.n100 585
R369 B.n603 B.n602 585
R370 B.n604 B.n99 585
R371 B.n606 B.n605 585
R372 B.n607 B.n98 585
R373 B.n609 B.n608 585
R374 B.n610 B.n97 585
R375 B.n612 B.n611 585
R376 B.n613 B.n96 585
R377 B.n615 B.n614 585
R378 B.n616 B.n95 585
R379 B.n618 B.n617 585
R380 B.n619 B.n94 585
R381 B.n621 B.n620 585
R382 B.n622 B.n93 585
R383 B.n624 B.n623 585
R384 B.n625 B.n92 585
R385 B.n627 B.n626 585
R386 B.n628 B.n91 585
R387 B.n630 B.n629 585
R388 B.n631 B.n90 585
R389 B.n633 B.n632 585
R390 B.n634 B.n89 585
R391 B.n636 B.n635 585
R392 B.n804 B.n803 585
R393 B.n802 B.n29 585
R394 B.n801 B.n800 585
R395 B.n799 B.n30 585
R396 B.n798 B.n797 585
R397 B.n796 B.n31 585
R398 B.n795 B.n794 585
R399 B.n793 B.n32 585
R400 B.n792 B.n791 585
R401 B.n790 B.n33 585
R402 B.n789 B.n788 585
R403 B.n787 B.n34 585
R404 B.n786 B.n785 585
R405 B.n784 B.n35 585
R406 B.n783 B.n782 585
R407 B.n781 B.n36 585
R408 B.n780 B.n779 585
R409 B.n778 B.n37 585
R410 B.n777 B.n776 585
R411 B.n775 B.n38 585
R412 B.n774 B.n773 585
R413 B.n772 B.n39 585
R414 B.n771 B.n770 585
R415 B.n769 B.n40 585
R416 B.n768 B.n767 585
R417 B.n766 B.n41 585
R418 B.n765 B.n764 585
R419 B.n763 B.n42 585
R420 B.n762 B.n761 585
R421 B.n760 B.n43 585
R422 B.n759 B.n758 585
R423 B.n757 B.n44 585
R424 B.n756 B.n755 585
R425 B.n754 B.n45 585
R426 B.n753 B.n752 585
R427 B.n751 B.n46 585
R428 B.n750 B.n749 585
R429 B.n748 B.n47 585
R430 B.n747 B.n746 585
R431 B.n745 B.n48 585
R432 B.n744 B.n743 585
R433 B.n742 B.n49 585
R434 B.n741 B.n740 585
R435 B.n739 B.n50 585
R436 B.n738 B.n737 585
R437 B.n736 B.n51 585
R438 B.n735 B.n734 585
R439 B.n733 B.n52 585
R440 B.n732 B.n731 585
R441 B.n730 B.n53 585
R442 B.n729 B.n728 585
R443 B.n727 B.n726 585
R444 B.n725 B.n57 585
R445 B.n724 B.n723 585
R446 B.n722 B.n58 585
R447 B.n721 B.n720 585
R448 B.n719 B.n59 585
R449 B.n718 B.n717 585
R450 B.n716 B.n60 585
R451 B.n715 B.n714 585
R452 B.n712 B.n61 585
R453 B.n711 B.n710 585
R454 B.n709 B.n64 585
R455 B.n708 B.n707 585
R456 B.n706 B.n65 585
R457 B.n705 B.n704 585
R458 B.n703 B.n66 585
R459 B.n702 B.n701 585
R460 B.n700 B.n67 585
R461 B.n699 B.n698 585
R462 B.n697 B.n68 585
R463 B.n696 B.n695 585
R464 B.n694 B.n69 585
R465 B.n693 B.n692 585
R466 B.n691 B.n70 585
R467 B.n690 B.n689 585
R468 B.n688 B.n71 585
R469 B.n687 B.n686 585
R470 B.n685 B.n72 585
R471 B.n684 B.n683 585
R472 B.n682 B.n73 585
R473 B.n681 B.n680 585
R474 B.n679 B.n74 585
R475 B.n678 B.n677 585
R476 B.n676 B.n75 585
R477 B.n675 B.n674 585
R478 B.n673 B.n76 585
R479 B.n672 B.n671 585
R480 B.n670 B.n77 585
R481 B.n669 B.n668 585
R482 B.n667 B.n78 585
R483 B.n666 B.n665 585
R484 B.n664 B.n79 585
R485 B.n663 B.n662 585
R486 B.n661 B.n80 585
R487 B.n660 B.n659 585
R488 B.n658 B.n81 585
R489 B.n657 B.n656 585
R490 B.n655 B.n82 585
R491 B.n654 B.n653 585
R492 B.n652 B.n83 585
R493 B.n651 B.n650 585
R494 B.n649 B.n84 585
R495 B.n648 B.n647 585
R496 B.n646 B.n85 585
R497 B.n645 B.n644 585
R498 B.n643 B.n86 585
R499 B.n642 B.n641 585
R500 B.n640 B.n87 585
R501 B.n639 B.n638 585
R502 B.n637 B.n88 585
R503 B.n805 B.n28 585
R504 B.n807 B.n806 585
R505 B.n808 B.n27 585
R506 B.n810 B.n809 585
R507 B.n811 B.n26 585
R508 B.n813 B.n812 585
R509 B.n814 B.n25 585
R510 B.n816 B.n815 585
R511 B.n817 B.n24 585
R512 B.n819 B.n818 585
R513 B.n820 B.n23 585
R514 B.n822 B.n821 585
R515 B.n823 B.n22 585
R516 B.n825 B.n824 585
R517 B.n826 B.n21 585
R518 B.n828 B.n827 585
R519 B.n829 B.n20 585
R520 B.n831 B.n830 585
R521 B.n832 B.n19 585
R522 B.n834 B.n833 585
R523 B.n835 B.n18 585
R524 B.n837 B.n836 585
R525 B.n838 B.n17 585
R526 B.n840 B.n839 585
R527 B.n841 B.n16 585
R528 B.n843 B.n842 585
R529 B.n844 B.n15 585
R530 B.n846 B.n845 585
R531 B.n847 B.n14 585
R532 B.n849 B.n848 585
R533 B.n850 B.n13 585
R534 B.n852 B.n851 585
R535 B.n853 B.n12 585
R536 B.n855 B.n854 585
R537 B.n856 B.n11 585
R538 B.n858 B.n857 585
R539 B.n859 B.n10 585
R540 B.n861 B.n860 585
R541 B.n862 B.n9 585
R542 B.n864 B.n863 585
R543 B.n865 B.n8 585
R544 B.n867 B.n866 585
R545 B.n868 B.n7 585
R546 B.n870 B.n869 585
R547 B.n871 B.n6 585
R548 B.n873 B.n872 585
R549 B.n874 B.n5 585
R550 B.n876 B.n875 585
R551 B.n877 B.n4 585
R552 B.n879 B.n878 585
R553 B.n880 B.n3 585
R554 B.n882 B.n881 585
R555 B.n883 B.n0 585
R556 B.n2 B.n1 585
R557 B.n229 B.n228 585
R558 B.n231 B.n230 585
R559 B.n232 B.n227 585
R560 B.n234 B.n233 585
R561 B.n235 B.n226 585
R562 B.n237 B.n236 585
R563 B.n238 B.n225 585
R564 B.n240 B.n239 585
R565 B.n241 B.n224 585
R566 B.n243 B.n242 585
R567 B.n244 B.n223 585
R568 B.n246 B.n245 585
R569 B.n247 B.n222 585
R570 B.n249 B.n248 585
R571 B.n250 B.n221 585
R572 B.n252 B.n251 585
R573 B.n253 B.n220 585
R574 B.n255 B.n254 585
R575 B.n256 B.n219 585
R576 B.n258 B.n257 585
R577 B.n259 B.n218 585
R578 B.n261 B.n260 585
R579 B.n262 B.n217 585
R580 B.n264 B.n263 585
R581 B.n265 B.n216 585
R582 B.n267 B.n266 585
R583 B.n268 B.n215 585
R584 B.n270 B.n269 585
R585 B.n271 B.n214 585
R586 B.n273 B.n272 585
R587 B.n274 B.n213 585
R588 B.n276 B.n275 585
R589 B.n277 B.n212 585
R590 B.n279 B.n278 585
R591 B.n280 B.n211 585
R592 B.n282 B.n281 585
R593 B.n283 B.n210 585
R594 B.n285 B.n284 585
R595 B.n286 B.n209 585
R596 B.n288 B.n287 585
R597 B.n289 B.n208 585
R598 B.n291 B.n290 585
R599 B.n292 B.n207 585
R600 B.n294 B.n293 585
R601 B.n295 B.n206 585
R602 B.n297 B.n296 585
R603 B.n298 B.n205 585
R604 B.n300 B.n299 585
R605 B.n301 B.n204 585
R606 B.n303 B.n302 585
R607 B.n304 B.n203 585
R608 B.n306 B.n305 585
R609 B.n307 B.n306 554.963
R610 B.n475 B.n474 554.963
R611 B.n637 B.n636 554.963
R612 B.n805 B.n804 554.963
R613 B.n176 B.t0 369.83
R614 B.n168 B.t9 369.83
R615 B.n62 B.t6 369.83
R616 B.n54 B.t3 369.83
R617 B.n885 B.n884 256.663
R618 B.n884 B.n883 235.042
R619 B.n884 B.n2 235.042
R620 B.n308 B.n307 163.367
R621 B.n308 B.n201 163.367
R622 B.n312 B.n201 163.367
R623 B.n313 B.n312 163.367
R624 B.n314 B.n313 163.367
R625 B.n314 B.n199 163.367
R626 B.n318 B.n199 163.367
R627 B.n319 B.n318 163.367
R628 B.n320 B.n319 163.367
R629 B.n320 B.n197 163.367
R630 B.n324 B.n197 163.367
R631 B.n325 B.n324 163.367
R632 B.n326 B.n325 163.367
R633 B.n326 B.n195 163.367
R634 B.n330 B.n195 163.367
R635 B.n331 B.n330 163.367
R636 B.n332 B.n331 163.367
R637 B.n332 B.n193 163.367
R638 B.n336 B.n193 163.367
R639 B.n337 B.n336 163.367
R640 B.n338 B.n337 163.367
R641 B.n338 B.n191 163.367
R642 B.n342 B.n191 163.367
R643 B.n343 B.n342 163.367
R644 B.n344 B.n343 163.367
R645 B.n344 B.n189 163.367
R646 B.n348 B.n189 163.367
R647 B.n349 B.n348 163.367
R648 B.n350 B.n349 163.367
R649 B.n350 B.n187 163.367
R650 B.n354 B.n187 163.367
R651 B.n355 B.n354 163.367
R652 B.n356 B.n355 163.367
R653 B.n356 B.n185 163.367
R654 B.n360 B.n185 163.367
R655 B.n361 B.n360 163.367
R656 B.n362 B.n361 163.367
R657 B.n362 B.n183 163.367
R658 B.n366 B.n183 163.367
R659 B.n367 B.n366 163.367
R660 B.n368 B.n367 163.367
R661 B.n368 B.n181 163.367
R662 B.n372 B.n181 163.367
R663 B.n373 B.n372 163.367
R664 B.n374 B.n373 163.367
R665 B.n374 B.n179 163.367
R666 B.n378 B.n179 163.367
R667 B.n379 B.n378 163.367
R668 B.n380 B.n379 163.367
R669 B.n380 B.n175 163.367
R670 B.n385 B.n175 163.367
R671 B.n386 B.n385 163.367
R672 B.n387 B.n386 163.367
R673 B.n387 B.n173 163.367
R674 B.n391 B.n173 163.367
R675 B.n392 B.n391 163.367
R676 B.n393 B.n392 163.367
R677 B.n393 B.n171 163.367
R678 B.n397 B.n171 163.367
R679 B.n398 B.n397 163.367
R680 B.n398 B.n167 163.367
R681 B.n402 B.n167 163.367
R682 B.n403 B.n402 163.367
R683 B.n404 B.n403 163.367
R684 B.n404 B.n165 163.367
R685 B.n408 B.n165 163.367
R686 B.n409 B.n408 163.367
R687 B.n410 B.n409 163.367
R688 B.n410 B.n163 163.367
R689 B.n414 B.n163 163.367
R690 B.n415 B.n414 163.367
R691 B.n416 B.n415 163.367
R692 B.n416 B.n161 163.367
R693 B.n420 B.n161 163.367
R694 B.n421 B.n420 163.367
R695 B.n422 B.n421 163.367
R696 B.n422 B.n159 163.367
R697 B.n426 B.n159 163.367
R698 B.n427 B.n426 163.367
R699 B.n428 B.n427 163.367
R700 B.n428 B.n157 163.367
R701 B.n432 B.n157 163.367
R702 B.n433 B.n432 163.367
R703 B.n434 B.n433 163.367
R704 B.n434 B.n155 163.367
R705 B.n438 B.n155 163.367
R706 B.n439 B.n438 163.367
R707 B.n440 B.n439 163.367
R708 B.n440 B.n153 163.367
R709 B.n444 B.n153 163.367
R710 B.n445 B.n444 163.367
R711 B.n446 B.n445 163.367
R712 B.n446 B.n151 163.367
R713 B.n450 B.n151 163.367
R714 B.n451 B.n450 163.367
R715 B.n452 B.n451 163.367
R716 B.n452 B.n149 163.367
R717 B.n456 B.n149 163.367
R718 B.n457 B.n456 163.367
R719 B.n458 B.n457 163.367
R720 B.n458 B.n147 163.367
R721 B.n462 B.n147 163.367
R722 B.n463 B.n462 163.367
R723 B.n464 B.n463 163.367
R724 B.n464 B.n145 163.367
R725 B.n468 B.n145 163.367
R726 B.n469 B.n468 163.367
R727 B.n470 B.n469 163.367
R728 B.n470 B.n143 163.367
R729 B.n474 B.n143 163.367
R730 B.n636 B.n89 163.367
R731 B.n632 B.n89 163.367
R732 B.n632 B.n631 163.367
R733 B.n631 B.n630 163.367
R734 B.n630 B.n91 163.367
R735 B.n626 B.n91 163.367
R736 B.n626 B.n625 163.367
R737 B.n625 B.n624 163.367
R738 B.n624 B.n93 163.367
R739 B.n620 B.n93 163.367
R740 B.n620 B.n619 163.367
R741 B.n619 B.n618 163.367
R742 B.n618 B.n95 163.367
R743 B.n614 B.n95 163.367
R744 B.n614 B.n613 163.367
R745 B.n613 B.n612 163.367
R746 B.n612 B.n97 163.367
R747 B.n608 B.n97 163.367
R748 B.n608 B.n607 163.367
R749 B.n607 B.n606 163.367
R750 B.n606 B.n99 163.367
R751 B.n602 B.n99 163.367
R752 B.n602 B.n601 163.367
R753 B.n601 B.n600 163.367
R754 B.n600 B.n101 163.367
R755 B.n596 B.n101 163.367
R756 B.n596 B.n595 163.367
R757 B.n595 B.n594 163.367
R758 B.n594 B.n103 163.367
R759 B.n590 B.n103 163.367
R760 B.n590 B.n589 163.367
R761 B.n589 B.n588 163.367
R762 B.n588 B.n105 163.367
R763 B.n584 B.n105 163.367
R764 B.n584 B.n583 163.367
R765 B.n583 B.n582 163.367
R766 B.n582 B.n107 163.367
R767 B.n578 B.n107 163.367
R768 B.n578 B.n577 163.367
R769 B.n577 B.n576 163.367
R770 B.n576 B.n109 163.367
R771 B.n572 B.n109 163.367
R772 B.n572 B.n571 163.367
R773 B.n571 B.n570 163.367
R774 B.n570 B.n111 163.367
R775 B.n566 B.n111 163.367
R776 B.n566 B.n565 163.367
R777 B.n565 B.n564 163.367
R778 B.n564 B.n113 163.367
R779 B.n560 B.n113 163.367
R780 B.n560 B.n559 163.367
R781 B.n559 B.n558 163.367
R782 B.n558 B.n115 163.367
R783 B.n554 B.n115 163.367
R784 B.n554 B.n553 163.367
R785 B.n553 B.n552 163.367
R786 B.n552 B.n117 163.367
R787 B.n548 B.n117 163.367
R788 B.n548 B.n547 163.367
R789 B.n547 B.n546 163.367
R790 B.n546 B.n119 163.367
R791 B.n542 B.n119 163.367
R792 B.n542 B.n541 163.367
R793 B.n541 B.n540 163.367
R794 B.n540 B.n121 163.367
R795 B.n536 B.n121 163.367
R796 B.n536 B.n535 163.367
R797 B.n535 B.n534 163.367
R798 B.n534 B.n123 163.367
R799 B.n530 B.n123 163.367
R800 B.n530 B.n529 163.367
R801 B.n529 B.n528 163.367
R802 B.n528 B.n125 163.367
R803 B.n524 B.n125 163.367
R804 B.n524 B.n523 163.367
R805 B.n523 B.n522 163.367
R806 B.n522 B.n127 163.367
R807 B.n518 B.n127 163.367
R808 B.n518 B.n517 163.367
R809 B.n517 B.n516 163.367
R810 B.n516 B.n129 163.367
R811 B.n512 B.n129 163.367
R812 B.n512 B.n511 163.367
R813 B.n511 B.n510 163.367
R814 B.n510 B.n131 163.367
R815 B.n506 B.n131 163.367
R816 B.n506 B.n505 163.367
R817 B.n505 B.n504 163.367
R818 B.n504 B.n133 163.367
R819 B.n500 B.n133 163.367
R820 B.n500 B.n499 163.367
R821 B.n499 B.n498 163.367
R822 B.n498 B.n135 163.367
R823 B.n494 B.n135 163.367
R824 B.n494 B.n493 163.367
R825 B.n493 B.n492 163.367
R826 B.n492 B.n137 163.367
R827 B.n488 B.n137 163.367
R828 B.n488 B.n487 163.367
R829 B.n487 B.n486 163.367
R830 B.n486 B.n139 163.367
R831 B.n482 B.n139 163.367
R832 B.n482 B.n481 163.367
R833 B.n481 B.n480 163.367
R834 B.n480 B.n141 163.367
R835 B.n476 B.n141 163.367
R836 B.n476 B.n475 163.367
R837 B.n804 B.n29 163.367
R838 B.n800 B.n29 163.367
R839 B.n800 B.n799 163.367
R840 B.n799 B.n798 163.367
R841 B.n798 B.n31 163.367
R842 B.n794 B.n31 163.367
R843 B.n794 B.n793 163.367
R844 B.n793 B.n792 163.367
R845 B.n792 B.n33 163.367
R846 B.n788 B.n33 163.367
R847 B.n788 B.n787 163.367
R848 B.n787 B.n786 163.367
R849 B.n786 B.n35 163.367
R850 B.n782 B.n35 163.367
R851 B.n782 B.n781 163.367
R852 B.n781 B.n780 163.367
R853 B.n780 B.n37 163.367
R854 B.n776 B.n37 163.367
R855 B.n776 B.n775 163.367
R856 B.n775 B.n774 163.367
R857 B.n774 B.n39 163.367
R858 B.n770 B.n39 163.367
R859 B.n770 B.n769 163.367
R860 B.n769 B.n768 163.367
R861 B.n768 B.n41 163.367
R862 B.n764 B.n41 163.367
R863 B.n764 B.n763 163.367
R864 B.n763 B.n762 163.367
R865 B.n762 B.n43 163.367
R866 B.n758 B.n43 163.367
R867 B.n758 B.n757 163.367
R868 B.n757 B.n756 163.367
R869 B.n756 B.n45 163.367
R870 B.n752 B.n45 163.367
R871 B.n752 B.n751 163.367
R872 B.n751 B.n750 163.367
R873 B.n750 B.n47 163.367
R874 B.n746 B.n47 163.367
R875 B.n746 B.n745 163.367
R876 B.n745 B.n744 163.367
R877 B.n744 B.n49 163.367
R878 B.n740 B.n49 163.367
R879 B.n740 B.n739 163.367
R880 B.n739 B.n738 163.367
R881 B.n738 B.n51 163.367
R882 B.n734 B.n51 163.367
R883 B.n734 B.n733 163.367
R884 B.n733 B.n732 163.367
R885 B.n732 B.n53 163.367
R886 B.n728 B.n53 163.367
R887 B.n728 B.n727 163.367
R888 B.n727 B.n57 163.367
R889 B.n723 B.n57 163.367
R890 B.n723 B.n722 163.367
R891 B.n722 B.n721 163.367
R892 B.n721 B.n59 163.367
R893 B.n717 B.n59 163.367
R894 B.n717 B.n716 163.367
R895 B.n716 B.n715 163.367
R896 B.n715 B.n61 163.367
R897 B.n710 B.n61 163.367
R898 B.n710 B.n709 163.367
R899 B.n709 B.n708 163.367
R900 B.n708 B.n65 163.367
R901 B.n704 B.n65 163.367
R902 B.n704 B.n703 163.367
R903 B.n703 B.n702 163.367
R904 B.n702 B.n67 163.367
R905 B.n698 B.n67 163.367
R906 B.n698 B.n697 163.367
R907 B.n697 B.n696 163.367
R908 B.n696 B.n69 163.367
R909 B.n692 B.n69 163.367
R910 B.n692 B.n691 163.367
R911 B.n691 B.n690 163.367
R912 B.n690 B.n71 163.367
R913 B.n686 B.n71 163.367
R914 B.n686 B.n685 163.367
R915 B.n685 B.n684 163.367
R916 B.n684 B.n73 163.367
R917 B.n680 B.n73 163.367
R918 B.n680 B.n679 163.367
R919 B.n679 B.n678 163.367
R920 B.n678 B.n75 163.367
R921 B.n674 B.n75 163.367
R922 B.n674 B.n673 163.367
R923 B.n673 B.n672 163.367
R924 B.n672 B.n77 163.367
R925 B.n668 B.n77 163.367
R926 B.n668 B.n667 163.367
R927 B.n667 B.n666 163.367
R928 B.n666 B.n79 163.367
R929 B.n662 B.n79 163.367
R930 B.n662 B.n661 163.367
R931 B.n661 B.n660 163.367
R932 B.n660 B.n81 163.367
R933 B.n656 B.n81 163.367
R934 B.n656 B.n655 163.367
R935 B.n655 B.n654 163.367
R936 B.n654 B.n83 163.367
R937 B.n650 B.n83 163.367
R938 B.n650 B.n649 163.367
R939 B.n649 B.n648 163.367
R940 B.n648 B.n85 163.367
R941 B.n644 B.n85 163.367
R942 B.n644 B.n643 163.367
R943 B.n643 B.n642 163.367
R944 B.n642 B.n87 163.367
R945 B.n638 B.n87 163.367
R946 B.n638 B.n637 163.367
R947 B.n806 B.n805 163.367
R948 B.n806 B.n27 163.367
R949 B.n810 B.n27 163.367
R950 B.n811 B.n810 163.367
R951 B.n812 B.n811 163.367
R952 B.n812 B.n25 163.367
R953 B.n816 B.n25 163.367
R954 B.n817 B.n816 163.367
R955 B.n818 B.n817 163.367
R956 B.n818 B.n23 163.367
R957 B.n822 B.n23 163.367
R958 B.n823 B.n822 163.367
R959 B.n824 B.n823 163.367
R960 B.n824 B.n21 163.367
R961 B.n828 B.n21 163.367
R962 B.n829 B.n828 163.367
R963 B.n830 B.n829 163.367
R964 B.n830 B.n19 163.367
R965 B.n834 B.n19 163.367
R966 B.n835 B.n834 163.367
R967 B.n836 B.n835 163.367
R968 B.n836 B.n17 163.367
R969 B.n840 B.n17 163.367
R970 B.n841 B.n840 163.367
R971 B.n842 B.n841 163.367
R972 B.n842 B.n15 163.367
R973 B.n846 B.n15 163.367
R974 B.n847 B.n846 163.367
R975 B.n848 B.n847 163.367
R976 B.n848 B.n13 163.367
R977 B.n852 B.n13 163.367
R978 B.n853 B.n852 163.367
R979 B.n854 B.n853 163.367
R980 B.n854 B.n11 163.367
R981 B.n858 B.n11 163.367
R982 B.n859 B.n858 163.367
R983 B.n860 B.n859 163.367
R984 B.n860 B.n9 163.367
R985 B.n864 B.n9 163.367
R986 B.n865 B.n864 163.367
R987 B.n866 B.n865 163.367
R988 B.n866 B.n7 163.367
R989 B.n870 B.n7 163.367
R990 B.n871 B.n870 163.367
R991 B.n872 B.n871 163.367
R992 B.n872 B.n5 163.367
R993 B.n876 B.n5 163.367
R994 B.n877 B.n876 163.367
R995 B.n878 B.n877 163.367
R996 B.n878 B.n3 163.367
R997 B.n882 B.n3 163.367
R998 B.n883 B.n882 163.367
R999 B.n229 B.n2 163.367
R1000 B.n230 B.n229 163.367
R1001 B.n230 B.n227 163.367
R1002 B.n234 B.n227 163.367
R1003 B.n235 B.n234 163.367
R1004 B.n236 B.n235 163.367
R1005 B.n236 B.n225 163.367
R1006 B.n240 B.n225 163.367
R1007 B.n241 B.n240 163.367
R1008 B.n242 B.n241 163.367
R1009 B.n242 B.n223 163.367
R1010 B.n246 B.n223 163.367
R1011 B.n247 B.n246 163.367
R1012 B.n248 B.n247 163.367
R1013 B.n248 B.n221 163.367
R1014 B.n252 B.n221 163.367
R1015 B.n253 B.n252 163.367
R1016 B.n254 B.n253 163.367
R1017 B.n254 B.n219 163.367
R1018 B.n258 B.n219 163.367
R1019 B.n259 B.n258 163.367
R1020 B.n260 B.n259 163.367
R1021 B.n260 B.n217 163.367
R1022 B.n264 B.n217 163.367
R1023 B.n265 B.n264 163.367
R1024 B.n266 B.n265 163.367
R1025 B.n266 B.n215 163.367
R1026 B.n270 B.n215 163.367
R1027 B.n271 B.n270 163.367
R1028 B.n272 B.n271 163.367
R1029 B.n272 B.n213 163.367
R1030 B.n276 B.n213 163.367
R1031 B.n277 B.n276 163.367
R1032 B.n278 B.n277 163.367
R1033 B.n278 B.n211 163.367
R1034 B.n282 B.n211 163.367
R1035 B.n283 B.n282 163.367
R1036 B.n284 B.n283 163.367
R1037 B.n284 B.n209 163.367
R1038 B.n288 B.n209 163.367
R1039 B.n289 B.n288 163.367
R1040 B.n290 B.n289 163.367
R1041 B.n290 B.n207 163.367
R1042 B.n294 B.n207 163.367
R1043 B.n295 B.n294 163.367
R1044 B.n296 B.n295 163.367
R1045 B.n296 B.n205 163.367
R1046 B.n300 B.n205 163.367
R1047 B.n301 B.n300 163.367
R1048 B.n302 B.n301 163.367
R1049 B.n302 B.n203 163.367
R1050 B.n306 B.n203 163.367
R1051 B.n168 B.t10 160.453
R1052 B.n62 B.t8 160.453
R1053 B.n176 B.t1 160.435
R1054 B.n54 B.t5 160.435
R1055 B.n169 B.t11 110.418
R1056 B.n63 B.t7 110.418
R1057 B.n177 B.t2 110.398
R1058 B.n55 B.t4 110.398
R1059 B.n383 B.n177 59.5399
R1060 B.n170 B.n169 59.5399
R1061 B.n713 B.n63 59.5399
R1062 B.n56 B.n55 59.5399
R1063 B.n177 B.n176 50.0369
R1064 B.n169 B.n168 50.0369
R1065 B.n63 B.n62 50.0369
R1066 B.n55 B.n54 50.0369
R1067 B.n803 B.n28 36.059
R1068 B.n635 B.n88 36.059
R1069 B.n305 B.n202 36.059
R1070 B.n473 B.n142 36.059
R1071 B B.n885 18.0485
R1072 B.n807 B.n28 10.6151
R1073 B.n808 B.n807 10.6151
R1074 B.n809 B.n808 10.6151
R1075 B.n809 B.n26 10.6151
R1076 B.n813 B.n26 10.6151
R1077 B.n814 B.n813 10.6151
R1078 B.n815 B.n814 10.6151
R1079 B.n815 B.n24 10.6151
R1080 B.n819 B.n24 10.6151
R1081 B.n820 B.n819 10.6151
R1082 B.n821 B.n820 10.6151
R1083 B.n821 B.n22 10.6151
R1084 B.n825 B.n22 10.6151
R1085 B.n826 B.n825 10.6151
R1086 B.n827 B.n826 10.6151
R1087 B.n827 B.n20 10.6151
R1088 B.n831 B.n20 10.6151
R1089 B.n832 B.n831 10.6151
R1090 B.n833 B.n832 10.6151
R1091 B.n833 B.n18 10.6151
R1092 B.n837 B.n18 10.6151
R1093 B.n838 B.n837 10.6151
R1094 B.n839 B.n838 10.6151
R1095 B.n839 B.n16 10.6151
R1096 B.n843 B.n16 10.6151
R1097 B.n844 B.n843 10.6151
R1098 B.n845 B.n844 10.6151
R1099 B.n845 B.n14 10.6151
R1100 B.n849 B.n14 10.6151
R1101 B.n850 B.n849 10.6151
R1102 B.n851 B.n850 10.6151
R1103 B.n851 B.n12 10.6151
R1104 B.n855 B.n12 10.6151
R1105 B.n856 B.n855 10.6151
R1106 B.n857 B.n856 10.6151
R1107 B.n857 B.n10 10.6151
R1108 B.n861 B.n10 10.6151
R1109 B.n862 B.n861 10.6151
R1110 B.n863 B.n862 10.6151
R1111 B.n863 B.n8 10.6151
R1112 B.n867 B.n8 10.6151
R1113 B.n868 B.n867 10.6151
R1114 B.n869 B.n868 10.6151
R1115 B.n869 B.n6 10.6151
R1116 B.n873 B.n6 10.6151
R1117 B.n874 B.n873 10.6151
R1118 B.n875 B.n874 10.6151
R1119 B.n875 B.n4 10.6151
R1120 B.n879 B.n4 10.6151
R1121 B.n880 B.n879 10.6151
R1122 B.n881 B.n880 10.6151
R1123 B.n881 B.n0 10.6151
R1124 B.n803 B.n802 10.6151
R1125 B.n802 B.n801 10.6151
R1126 B.n801 B.n30 10.6151
R1127 B.n797 B.n30 10.6151
R1128 B.n797 B.n796 10.6151
R1129 B.n796 B.n795 10.6151
R1130 B.n795 B.n32 10.6151
R1131 B.n791 B.n32 10.6151
R1132 B.n791 B.n790 10.6151
R1133 B.n790 B.n789 10.6151
R1134 B.n789 B.n34 10.6151
R1135 B.n785 B.n34 10.6151
R1136 B.n785 B.n784 10.6151
R1137 B.n784 B.n783 10.6151
R1138 B.n783 B.n36 10.6151
R1139 B.n779 B.n36 10.6151
R1140 B.n779 B.n778 10.6151
R1141 B.n778 B.n777 10.6151
R1142 B.n777 B.n38 10.6151
R1143 B.n773 B.n38 10.6151
R1144 B.n773 B.n772 10.6151
R1145 B.n772 B.n771 10.6151
R1146 B.n771 B.n40 10.6151
R1147 B.n767 B.n40 10.6151
R1148 B.n767 B.n766 10.6151
R1149 B.n766 B.n765 10.6151
R1150 B.n765 B.n42 10.6151
R1151 B.n761 B.n42 10.6151
R1152 B.n761 B.n760 10.6151
R1153 B.n760 B.n759 10.6151
R1154 B.n759 B.n44 10.6151
R1155 B.n755 B.n44 10.6151
R1156 B.n755 B.n754 10.6151
R1157 B.n754 B.n753 10.6151
R1158 B.n753 B.n46 10.6151
R1159 B.n749 B.n46 10.6151
R1160 B.n749 B.n748 10.6151
R1161 B.n748 B.n747 10.6151
R1162 B.n747 B.n48 10.6151
R1163 B.n743 B.n48 10.6151
R1164 B.n743 B.n742 10.6151
R1165 B.n742 B.n741 10.6151
R1166 B.n741 B.n50 10.6151
R1167 B.n737 B.n50 10.6151
R1168 B.n737 B.n736 10.6151
R1169 B.n736 B.n735 10.6151
R1170 B.n735 B.n52 10.6151
R1171 B.n731 B.n52 10.6151
R1172 B.n731 B.n730 10.6151
R1173 B.n730 B.n729 10.6151
R1174 B.n726 B.n725 10.6151
R1175 B.n725 B.n724 10.6151
R1176 B.n724 B.n58 10.6151
R1177 B.n720 B.n58 10.6151
R1178 B.n720 B.n719 10.6151
R1179 B.n719 B.n718 10.6151
R1180 B.n718 B.n60 10.6151
R1181 B.n714 B.n60 10.6151
R1182 B.n712 B.n711 10.6151
R1183 B.n711 B.n64 10.6151
R1184 B.n707 B.n64 10.6151
R1185 B.n707 B.n706 10.6151
R1186 B.n706 B.n705 10.6151
R1187 B.n705 B.n66 10.6151
R1188 B.n701 B.n66 10.6151
R1189 B.n701 B.n700 10.6151
R1190 B.n700 B.n699 10.6151
R1191 B.n699 B.n68 10.6151
R1192 B.n695 B.n68 10.6151
R1193 B.n695 B.n694 10.6151
R1194 B.n694 B.n693 10.6151
R1195 B.n693 B.n70 10.6151
R1196 B.n689 B.n70 10.6151
R1197 B.n689 B.n688 10.6151
R1198 B.n688 B.n687 10.6151
R1199 B.n687 B.n72 10.6151
R1200 B.n683 B.n72 10.6151
R1201 B.n683 B.n682 10.6151
R1202 B.n682 B.n681 10.6151
R1203 B.n681 B.n74 10.6151
R1204 B.n677 B.n74 10.6151
R1205 B.n677 B.n676 10.6151
R1206 B.n676 B.n675 10.6151
R1207 B.n675 B.n76 10.6151
R1208 B.n671 B.n76 10.6151
R1209 B.n671 B.n670 10.6151
R1210 B.n670 B.n669 10.6151
R1211 B.n669 B.n78 10.6151
R1212 B.n665 B.n78 10.6151
R1213 B.n665 B.n664 10.6151
R1214 B.n664 B.n663 10.6151
R1215 B.n663 B.n80 10.6151
R1216 B.n659 B.n80 10.6151
R1217 B.n659 B.n658 10.6151
R1218 B.n658 B.n657 10.6151
R1219 B.n657 B.n82 10.6151
R1220 B.n653 B.n82 10.6151
R1221 B.n653 B.n652 10.6151
R1222 B.n652 B.n651 10.6151
R1223 B.n651 B.n84 10.6151
R1224 B.n647 B.n84 10.6151
R1225 B.n647 B.n646 10.6151
R1226 B.n646 B.n645 10.6151
R1227 B.n645 B.n86 10.6151
R1228 B.n641 B.n86 10.6151
R1229 B.n641 B.n640 10.6151
R1230 B.n640 B.n639 10.6151
R1231 B.n639 B.n88 10.6151
R1232 B.n635 B.n634 10.6151
R1233 B.n634 B.n633 10.6151
R1234 B.n633 B.n90 10.6151
R1235 B.n629 B.n90 10.6151
R1236 B.n629 B.n628 10.6151
R1237 B.n628 B.n627 10.6151
R1238 B.n627 B.n92 10.6151
R1239 B.n623 B.n92 10.6151
R1240 B.n623 B.n622 10.6151
R1241 B.n622 B.n621 10.6151
R1242 B.n621 B.n94 10.6151
R1243 B.n617 B.n94 10.6151
R1244 B.n617 B.n616 10.6151
R1245 B.n616 B.n615 10.6151
R1246 B.n615 B.n96 10.6151
R1247 B.n611 B.n96 10.6151
R1248 B.n611 B.n610 10.6151
R1249 B.n610 B.n609 10.6151
R1250 B.n609 B.n98 10.6151
R1251 B.n605 B.n98 10.6151
R1252 B.n605 B.n604 10.6151
R1253 B.n604 B.n603 10.6151
R1254 B.n603 B.n100 10.6151
R1255 B.n599 B.n100 10.6151
R1256 B.n599 B.n598 10.6151
R1257 B.n598 B.n597 10.6151
R1258 B.n597 B.n102 10.6151
R1259 B.n593 B.n102 10.6151
R1260 B.n593 B.n592 10.6151
R1261 B.n592 B.n591 10.6151
R1262 B.n591 B.n104 10.6151
R1263 B.n587 B.n104 10.6151
R1264 B.n587 B.n586 10.6151
R1265 B.n586 B.n585 10.6151
R1266 B.n585 B.n106 10.6151
R1267 B.n581 B.n106 10.6151
R1268 B.n581 B.n580 10.6151
R1269 B.n580 B.n579 10.6151
R1270 B.n579 B.n108 10.6151
R1271 B.n575 B.n108 10.6151
R1272 B.n575 B.n574 10.6151
R1273 B.n574 B.n573 10.6151
R1274 B.n573 B.n110 10.6151
R1275 B.n569 B.n110 10.6151
R1276 B.n569 B.n568 10.6151
R1277 B.n568 B.n567 10.6151
R1278 B.n567 B.n112 10.6151
R1279 B.n563 B.n112 10.6151
R1280 B.n563 B.n562 10.6151
R1281 B.n562 B.n561 10.6151
R1282 B.n561 B.n114 10.6151
R1283 B.n557 B.n114 10.6151
R1284 B.n557 B.n556 10.6151
R1285 B.n556 B.n555 10.6151
R1286 B.n555 B.n116 10.6151
R1287 B.n551 B.n116 10.6151
R1288 B.n551 B.n550 10.6151
R1289 B.n550 B.n549 10.6151
R1290 B.n549 B.n118 10.6151
R1291 B.n545 B.n118 10.6151
R1292 B.n545 B.n544 10.6151
R1293 B.n544 B.n543 10.6151
R1294 B.n543 B.n120 10.6151
R1295 B.n539 B.n120 10.6151
R1296 B.n539 B.n538 10.6151
R1297 B.n538 B.n537 10.6151
R1298 B.n537 B.n122 10.6151
R1299 B.n533 B.n122 10.6151
R1300 B.n533 B.n532 10.6151
R1301 B.n532 B.n531 10.6151
R1302 B.n531 B.n124 10.6151
R1303 B.n527 B.n124 10.6151
R1304 B.n527 B.n526 10.6151
R1305 B.n526 B.n525 10.6151
R1306 B.n525 B.n126 10.6151
R1307 B.n521 B.n126 10.6151
R1308 B.n521 B.n520 10.6151
R1309 B.n520 B.n519 10.6151
R1310 B.n519 B.n128 10.6151
R1311 B.n515 B.n128 10.6151
R1312 B.n515 B.n514 10.6151
R1313 B.n514 B.n513 10.6151
R1314 B.n513 B.n130 10.6151
R1315 B.n509 B.n130 10.6151
R1316 B.n509 B.n508 10.6151
R1317 B.n508 B.n507 10.6151
R1318 B.n507 B.n132 10.6151
R1319 B.n503 B.n132 10.6151
R1320 B.n503 B.n502 10.6151
R1321 B.n502 B.n501 10.6151
R1322 B.n501 B.n134 10.6151
R1323 B.n497 B.n134 10.6151
R1324 B.n497 B.n496 10.6151
R1325 B.n496 B.n495 10.6151
R1326 B.n495 B.n136 10.6151
R1327 B.n491 B.n136 10.6151
R1328 B.n491 B.n490 10.6151
R1329 B.n490 B.n489 10.6151
R1330 B.n489 B.n138 10.6151
R1331 B.n485 B.n138 10.6151
R1332 B.n485 B.n484 10.6151
R1333 B.n484 B.n483 10.6151
R1334 B.n483 B.n140 10.6151
R1335 B.n479 B.n140 10.6151
R1336 B.n479 B.n478 10.6151
R1337 B.n478 B.n477 10.6151
R1338 B.n477 B.n142 10.6151
R1339 B.n228 B.n1 10.6151
R1340 B.n231 B.n228 10.6151
R1341 B.n232 B.n231 10.6151
R1342 B.n233 B.n232 10.6151
R1343 B.n233 B.n226 10.6151
R1344 B.n237 B.n226 10.6151
R1345 B.n238 B.n237 10.6151
R1346 B.n239 B.n238 10.6151
R1347 B.n239 B.n224 10.6151
R1348 B.n243 B.n224 10.6151
R1349 B.n244 B.n243 10.6151
R1350 B.n245 B.n244 10.6151
R1351 B.n245 B.n222 10.6151
R1352 B.n249 B.n222 10.6151
R1353 B.n250 B.n249 10.6151
R1354 B.n251 B.n250 10.6151
R1355 B.n251 B.n220 10.6151
R1356 B.n255 B.n220 10.6151
R1357 B.n256 B.n255 10.6151
R1358 B.n257 B.n256 10.6151
R1359 B.n257 B.n218 10.6151
R1360 B.n261 B.n218 10.6151
R1361 B.n262 B.n261 10.6151
R1362 B.n263 B.n262 10.6151
R1363 B.n263 B.n216 10.6151
R1364 B.n267 B.n216 10.6151
R1365 B.n268 B.n267 10.6151
R1366 B.n269 B.n268 10.6151
R1367 B.n269 B.n214 10.6151
R1368 B.n273 B.n214 10.6151
R1369 B.n274 B.n273 10.6151
R1370 B.n275 B.n274 10.6151
R1371 B.n275 B.n212 10.6151
R1372 B.n279 B.n212 10.6151
R1373 B.n280 B.n279 10.6151
R1374 B.n281 B.n280 10.6151
R1375 B.n281 B.n210 10.6151
R1376 B.n285 B.n210 10.6151
R1377 B.n286 B.n285 10.6151
R1378 B.n287 B.n286 10.6151
R1379 B.n287 B.n208 10.6151
R1380 B.n291 B.n208 10.6151
R1381 B.n292 B.n291 10.6151
R1382 B.n293 B.n292 10.6151
R1383 B.n293 B.n206 10.6151
R1384 B.n297 B.n206 10.6151
R1385 B.n298 B.n297 10.6151
R1386 B.n299 B.n298 10.6151
R1387 B.n299 B.n204 10.6151
R1388 B.n303 B.n204 10.6151
R1389 B.n304 B.n303 10.6151
R1390 B.n305 B.n304 10.6151
R1391 B.n309 B.n202 10.6151
R1392 B.n310 B.n309 10.6151
R1393 B.n311 B.n310 10.6151
R1394 B.n311 B.n200 10.6151
R1395 B.n315 B.n200 10.6151
R1396 B.n316 B.n315 10.6151
R1397 B.n317 B.n316 10.6151
R1398 B.n317 B.n198 10.6151
R1399 B.n321 B.n198 10.6151
R1400 B.n322 B.n321 10.6151
R1401 B.n323 B.n322 10.6151
R1402 B.n323 B.n196 10.6151
R1403 B.n327 B.n196 10.6151
R1404 B.n328 B.n327 10.6151
R1405 B.n329 B.n328 10.6151
R1406 B.n329 B.n194 10.6151
R1407 B.n333 B.n194 10.6151
R1408 B.n334 B.n333 10.6151
R1409 B.n335 B.n334 10.6151
R1410 B.n335 B.n192 10.6151
R1411 B.n339 B.n192 10.6151
R1412 B.n340 B.n339 10.6151
R1413 B.n341 B.n340 10.6151
R1414 B.n341 B.n190 10.6151
R1415 B.n345 B.n190 10.6151
R1416 B.n346 B.n345 10.6151
R1417 B.n347 B.n346 10.6151
R1418 B.n347 B.n188 10.6151
R1419 B.n351 B.n188 10.6151
R1420 B.n352 B.n351 10.6151
R1421 B.n353 B.n352 10.6151
R1422 B.n353 B.n186 10.6151
R1423 B.n357 B.n186 10.6151
R1424 B.n358 B.n357 10.6151
R1425 B.n359 B.n358 10.6151
R1426 B.n359 B.n184 10.6151
R1427 B.n363 B.n184 10.6151
R1428 B.n364 B.n363 10.6151
R1429 B.n365 B.n364 10.6151
R1430 B.n365 B.n182 10.6151
R1431 B.n369 B.n182 10.6151
R1432 B.n370 B.n369 10.6151
R1433 B.n371 B.n370 10.6151
R1434 B.n371 B.n180 10.6151
R1435 B.n375 B.n180 10.6151
R1436 B.n376 B.n375 10.6151
R1437 B.n377 B.n376 10.6151
R1438 B.n377 B.n178 10.6151
R1439 B.n381 B.n178 10.6151
R1440 B.n382 B.n381 10.6151
R1441 B.n384 B.n174 10.6151
R1442 B.n388 B.n174 10.6151
R1443 B.n389 B.n388 10.6151
R1444 B.n390 B.n389 10.6151
R1445 B.n390 B.n172 10.6151
R1446 B.n394 B.n172 10.6151
R1447 B.n395 B.n394 10.6151
R1448 B.n396 B.n395 10.6151
R1449 B.n400 B.n399 10.6151
R1450 B.n401 B.n400 10.6151
R1451 B.n401 B.n166 10.6151
R1452 B.n405 B.n166 10.6151
R1453 B.n406 B.n405 10.6151
R1454 B.n407 B.n406 10.6151
R1455 B.n407 B.n164 10.6151
R1456 B.n411 B.n164 10.6151
R1457 B.n412 B.n411 10.6151
R1458 B.n413 B.n412 10.6151
R1459 B.n413 B.n162 10.6151
R1460 B.n417 B.n162 10.6151
R1461 B.n418 B.n417 10.6151
R1462 B.n419 B.n418 10.6151
R1463 B.n419 B.n160 10.6151
R1464 B.n423 B.n160 10.6151
R1465 B.n424 B.n423 10.6151
R1466 B.n425 B.n424 10.6151
R1467 B.n425 B.n158 10.6151
R1468 B.n429 B.n158 10.6151
R1469 B.n430 B.n429 10.6151
R1470 B.n431 B.n430 10.6151
R1471 B.n431 B.n156 10.6151
R1472 B.n435 B.n156 10.6151
R1473 B.n436 B.n435 10.6151
R1474 B.n437 B.n436 10.6151
R1475 B.n437 B.n154 10.6151
R1476 B.n441 B.n154 10.6151
R1477 B.n442 B.n441 10.6151
R1478 B.n443 B.n442 10.6151
R1479 B.n443 B.n152 10.6151
R1480 B.n447 B.n152 10.6151
R1481 B.n448 B.n447 10.6151
R1482 B.n449 B.n448 10.6151
R1483 B.n449 B.n150 10.6151
R1484 B.n453 B.n150 10.6151
R1485 B.n454 B.n453 10.6151
R1486 B.n455 B.n454 10.6151
R1487 B.n455 B.n148 10.6151
R1488 B.n459 B.n148 10.6151
R1489 B.n460 B.n459 10.6151
R1490 B.n461 B.n460 10.6151
R1491 B.n461 B.n146 10.6151
R1492 B.n465 B.n146 10.6151
R1493 B.n466 B.n465 10.6151
R1494 B.n467 B.n466 10.6151
R1495 B.n467 B.n144 10.6151
R1496 B.n471 B.n144 10.6151
R1497 B.n472 B.n471 10.6151
R1498 B.n473 B.n472 10.6151
R1499 B.n885 B.n0 8.11757
R1500 B.n885 B.n1 8.11757
R1501 B.n726 B.n56 6.5566
R1502 B.n714 B.n713 6.5566
R1503 B.n384 B.n383 6.5566
R1504 B.n396 B.n170 6.5566
R1505 B.n729 B.n56 4.05904
R1506 B.n713 B.n712 4.05904
R1507 B.n383 B.n382 4.05904
R1508 B.n399 B.n170 4.05904
R1509 VP.n19 VP.t5 196.519
R1510 VP.n48 VP.t8 162.381
R1511 VP.n56 VP.t0 162.381
R1512 VP.n5 VP.t7 162.381
R1513 VP.n73 VP.t6 162.381
R1514 VP.n81 VP.t2 162.381
R1515 VP.n45 VP.t9 162.381
R1516 VP.n37 VP.t4 162.381
R1517 VP.n16 VP.t3 162.381
R1518 VP.n20 VP.t1 162.381
R1519 VP.n22 VP.n21 161.3
R1520 VP.n23 VP.n18 161.3
R1521 VP.n25 VP.n24 161.3
R1522 VP.n26 VP.n17 161.3
R1523 VP.n28 VP.n27 161.3
R1524 VP.n30 VP.n29 161.3
R1525 VP.n31 VP.n15 161.3
R1526 VP.n33 VP.n32 161.3
R1527 VP.n34 VP.n14 161.3
R1528 VP.n36 VP.n35 161.3
R1529 VP.n38 VP.n13 161.3
R1530 VP.n40 VP.n39 161.3
R1531 VP.n41 VP.n12 161.3
R1532 VP.n43 VP.n42 161.3
R1533 VP.n44 VP.n11 161.3
R1534 VP.n80 VP.n0 161.3
R1535 VP.n79 VP.n78 161.3
R1536 VP.n77 VP.n1 161.3
R1537 VP.n76 VP.n75 161.3
R1538 VP.n74 VP.n2 161.3
R1539 VP.n72 VP.n71 161.3
R1540 VP.n70 VP.n3 161.3
R1541 VP.n69 VP.n68 161.3
R1542 VP.n67 VP.n4 161.3
R1543 VP.n66 VP.n65 161.3
R1544 VP.n64 VP.n63 161.3
R1545 VP.n62 VP.n6 161.3
R1546 VP.n61 VP.n60 161.3
R1547 VP.n59 VP.n7 161.3
R1548 VP.n58 VP.n57 161.3
R1549 VP.n55 VP.n8 161.3
R1550 VP.n54 VP.n53 161.3
R1551 VP.n52 VP.n9 161.3
R1552 VP.n51 VP.n50 161.3
R1553 VP.n49 VP.n10 161.3
R1554 VP.n48 VP.n47 90.7429
R1555 VP.n82 VP.n81 90.7429
R1556 VP.n46 VP.n45 90.7429
R1557 VP.n20 VP.n19 55.0386
R1558 VP.n47 VP.n46 53.6966
R1559 VP.n50 VP.n9 52.2023
R1560 VP.n79 VP.n1 52.2023
R1561 VP.n43 VP.n12 52.2023
R1562 VP.n61 VP.n7 44.4521
R1563 VP.n68 VP.n3 44.4521
R1564 VP.n32 VP.n14 44.4521
R1565 VP.n25 VP.n18 44.4521
R1566 VP.n62 VP.n61 36.702
R1567 VP.n68 VP.n67 36.702
R1568 VP.n32 VP.n31 36.702
R1569 VP.n26 VP.n25 36.702
R1570 VP.n54 VP.n9 28.9518
R1571 VP.n75 VP.n1 28.9518
R1572 VP.n39 VP.n12 28.9518
R1573 VP.n50 VP.n49 24.5923
R1574 VP.n55 VP.n54 24.5923
R1575 VP.n57 VP.n7 24.5923
R1576 VP.n63 VP.n62 24.5923
R1577 VP.n67 VP.n66 24.5923
R1578 VP.n72 VP.n3 24.5923
R1579 VP.n75 VP.n74 24.5923
R1580 VP.n80 VP.n79 24.5923
R1581 VP.n44 VP.n43 24.5923
R1582 VP.n36 VP.n14 24.5923
R1583 VP.n39 VP.n38 24.5923
R1584 VP.n27 VP.n26 24.5923
R1585 VP.n31 VP.n30 24.5923
R1586 VP.n21 VP.n18 24.5923
R1587 VP.n49 VP.n48 20.1658
R1588 VP.n81 VP.n80 20.1658
R1589 VP.n45 VP.n44 20.1658
R1590 VP.n57 VP.n56 16.2311
R1591 VP.n73 VP.n72 16.2311
R1592 VP.n37 VP.n36 16.2311
R1593 VP.n21 VP.n20 16.2311
R1594 VP.n63 VP.n5 12.2964
R1595 VP.n66 VP.n5 12.2964
R1596 VP.n27 VP.n16 12.2964
R1597 VP.n30 VP.n16 12.2964
R1598 VP.n22 VP.n19 8.94118
R1599 VP.n56 VP.n55 8.36172
R1600 VP.n74 VP.n73 8.36172
R1601 VP.n38 VP.n37 8.36172
R1602 VP.n46 VP.n11 0.278335
R1603 VP.n47 VP.n10 0.278335
R1604 VP.n82 VP.n0 0.278335
R1605 VP.n23 VP.n22 0.189894
R1606 VP.n24 VP.n23 0.189894
R1607 VP.n24 VP.n17 0.189894
R1608 VP.n28 VP.n17 0.189894
R1609 VP.n29 VP.n28 0.189894
R1610 VP.n29 VP.n15 0.189894
R1611 VP.n33 VP.n15 0.189894
R1612 VP.n34 VP.n33 0.189894
R1613 VP.n35 VP.n34 0.189894
R1614 VP.n35 VP.n13 0.189894
R1615 VP.n40 VP.n13 0.189894
R1616 VP.n41 VP.n40 0.189894
R1617 VP.n42 VP.n41 0.189894
R1618 VP.n42 VP.n11 0.189894
R1619 VP.n51 VP.n10 0.189894
R1620 VP.n52 VP.n51 0.189894
R1621 VP.n53 VP.n52 0.189894
R1622 VP.n53 VP.n8 0.189894
R1623 VP.n58 VP.n8 0.189894
R1624 VP.n59 VP.n58 0.189894
R1625 VP.n60 VP.n59 0.189894
R1626 VP.n60 VP.n6 0.189894
R1627 VP.n64 VP.n6 0.189894
R1628 VP.n65 VP.n64 0.189894
R1629 VP.n65 VP.n4 0.189894
R1630 VP.n69 VP.n4 0.189894
R1631 VP.n70 VP.n69 0.189894
R1632 VP.n71 VP.n70 0.189894
R1633 VP.n71 VP.n2 0.189894
R1634 VP.n76 VP.n2 0.189894
R1635 VP.n77 VP.n76 0.189894
R1636 VP.n78 VP.n77 0.189894
R1637 VP.n78 VP.n0 0.189894
R1638 VP VP.n82 0.153485
R1639 VDD1.n1 VDD1.t4 77.9765
R1640 VDD1.n3 VDD1.t1 77.9762
R1641 VDD1.n5 VDD1.n4 75.2207
R1642 VDD1.n1 VDD1.n0 73.6082
R1643 VDD1.n7 VDD1.n6 73.608
R1644 VDD1.n3 VDD1.n2 73.6079
R1645 VDD1.n7 VDD1.n5 49.044
R1646 VDD1.n6 VDD1.t5 2.14463
R1647 VDD1.n6 VDD1.t0 2.14463
R1648 VDD1.n0 VDD1.t8 2.14463
R1649 VDD1.n0 VDD1.t6 2.14463
R1650 VDD1.n4 VDD1.t3 2.14463
R1651 VDD1.n4 VDD1.t7 2.14463
R1652 VDD1.n2 VDD1.t9 2.14463
R1653 VDD1.n2 VDD1.t2 2.14463
R1654 VDD1 VDD1.n7 1.61041
R1655 VDD1 VDD1.n1 0.614724
R1656 VDD1.n5 VDD1.n3 0.501188
C0 w_n4066_n4000# VDD1 2.87417f
C1 VP B 2.12135f
C2 VTAIL VDD1 11.944099f
C3 VDD2 VDD1 1.94593f
C4 VN VDD1 0.152728f
C5 w_n4066_n4000# VTAIL 3.60615f
C6 w_n4066_n4000# VDD2 2.99961f
C7 B VDD1 2.5908f
C8 VN w_n4066_n4000# 8.63469f
C9 VP VDD1 13.3205f
C10 VTAIL VDD2 11.991401f
C11 VN VTAIL 13.297f
C12 VN VDD2 12.938299f
C13 B w_n4066_n4000# 10.8444f
C14 VP w_n4066_n4000# 9.16298f
C15 B VTAIL 4.27006f
C16 B VDD2 2.69508f
C17 VP VTAIL 13.3114f
C18 VP VDD2 0.539393f
C19 B VN 1.23493f
C20 VP VN 8.45898f
C21 VDD2 VSUBS 2.04279f
C22 VDD1 VSUBS 1.889177f
C23 VTAIL VSUBS 1.324479f
C24 VN VSUBS 7.23544f
C25 VP VSUBS 3.912f
C26 B VSUBS 5.198293f
C27 w_n4066_n4000# VSUBS 0.199413p
C28 VDD1.t4 VSUBS 3.45553f
C29 VDD1.t8 VSUBS 0.323485f
C30 VDD1.t6 VSUBS 0.323485f
C31 VDD1.n0 VSUBS 2.64103f
C32 VDD1.n1 VSUBS 1.53046f
C33 VDD1.t1 VSUBS 3.45553f
C34 VDD1.t9 VSUBS 0.323485f
C35 VDD1.t2 VSUBS 0.323485f
C36 VDD1.n2 VSUBS 2.64103f
C37 VDD1.n3 VSUBS 1.52184f
C38 VDD1.t3 VSUBS 0.323485f
C39 VDD1.t7 VSUBS 0.323485f
C40 VDD1.n4 VSUBS 2.65927f
C41 VDD1.n5 VSUBS 3.55891f
C42 VDD1.t5 VSUBS 0.323485f
C43 VDD1.t0 VSUBS 0.323485f
C44 VDD1.n6 VSUBS 2.64102f
C45 VDD1.n7 VSUBS 3.814f
C46 VP.n0 VSUBS 0.040568f
C47 VP.t2 VSUBS 2.87692f
C48 VP.n1 VSUBS 0.031008f
C49 VP.n2 VSUBS 0.030772f
C50 VP.t6 VSUBS 2.87692f
C51 VP.n3 VSUBS 0.05933f
C52 VP.n4 VSUBS 0.030772f
C53 VP.t7 VSUBS 2.87692f
C54 VP.n5 VSUBS 1.00871f
C55 VP.n6 VSUBS 0.030772f
C56 VP.n7 VSUBS 0.05933f
C57 VP.n8 VSUBS 0.030772f
C58 VP.t0 VSUBS 2.87692f
C59 VP.n9 VSUBS 0.031008f
C60 VP.n10 VSUBS 0.040568f
C61 VP.t8 VSUBS 2.87692f
C62 VP.n11 VSUBS 0.040568f
C63 VP.t9 VSUBS 2.87692f
C64 VP.n12 VSUBS 0.031008f
C65 VP.n13 VSUBS 0.030772f
C66 VP.t4 VSUBS 2.87692f
C67 VP.n14 VSUBS 0.05933f
C68 VP.n15 VSUBS 0.030772f
C69 VP.t3 VSUBS 2.87692f
C70 VP.n16 VSUBS 1.00871f
C71 VP.n17 VSUBS 0.030772f
C72 VP.n18 VSUBS 0.05933f
C73 VP.t5 VSUBS 3.08238f
C74 VP.n19 VSUBS 1.0731f
C75 VP.t1 VSUBS 2.87692f
C76 VP.n20 VSUBS 1.09289f
C77 VP.n21 VSUBS 0.047486f
C78 VP.n22 VSUBS 0.263097f
C79 VP.n23 VSUBS 0.030772f
C80 VP.n24 VSUBS 0.030772f
C81 VP.n25 VSUBS 0.025487f
C82 VP.n26 VSUBS 0.061712f
C83 VP.n27 VSUBS 0.042979f
C84 VP.n28 VSUBS 0.030772f
C85 VP.n29 VSUBS 0.030772f
C86 VP.n30 VSUBS 0.042979f
C87 VP.n31 VSUBS 0.061712f
C88 VP.n32 VSUBS 0.025487f
C89 VP.n33 VSUBS 0.030772f
C90 VP.n34 VSUBS 0.030772f
C91 VP.n35 VSUBS 0.030772f
C92 VP.n36 VSUBS 0.047486f
C93 VP.n37 VSUBS 1.00871f
C94 VP.n38 VSUBS 0.038472f
C95 VP.n39 VSUBS 0.060543f
C96 VP.n40 VSUBS 0.030772f
C97 VP.n41 VSUBS 0.030772f
C98 VP.n42 VSUBS 0.030772f
C99 VP.n43 VSUBS 0.054979f
C100 VP.n44 VSUBS 0.051994f
C101 VP.n45 VSUBS 1.11462f
C102 VP.n46 VSUBS 1.88689f
C103 VP.n47 VSUBS 1.90755f
C104 VP.n48 VSUBS 1.11462f
C105 VP.n49 VSUBS 0.051994f
C106 VP.n50 VSUBS 0.054979f
C107 VP.n51 VSUBS 0.030772f
C108 VP.n52 VSUBS 0.030772f
C109 VP.n53 VSUBS 0.030772f
C110 VP.n54 VSUBS 0.060543f
C111 VP.n55 VSUBS 0.038472f
C112 VP.n56 VSUBS 1.00871f
C113 VP.n57 VSUBS 0.047486f
C114 VP.n58 VSUBS 0.030772f
C115 VP.n59 VSUBS 0.030772f
C116 VP.n60 VSUBS 0.030772f
C117 VP.n61 VSUBS 0.025487f
C118 VP.n62 VSUBS 0.061712f
C119 VP.n63 VSUBS 0.042979f
C120 VP.n64 VSUBS 0.030772f
C121 VP.n65 VSUBS 0.030772f
C122 VP.n66 VSUBS 0.042979f
C123 VP.n67 VSUBS 0.061712f
C124 VP.n68 VSUBS 0.025487f
C125 VP.n69 VSUBS 0.030772f
C126 VP.n70 VSUBS 0.030772f
C127 VP.n71 VSUBS 0.030772f
C128 VP.n72 VSUBS 0.047486f
C129 VP.n73 VSUBS 1.00871f
C130 VP.n74 VSUBS 0.038472f
C131 VP.n75 VSUBS 0.060543f
C132 VP.n76 VSUBS 0.030772f
C133 VP.n77 VSUBS 0.030772f
C134 VP.n78 VSUBS 0.030772f
C135 VP.n79 VSUBS 0.054979f
C136 VP.n80 VSUBS 0.051994f
C137 VP.n81 VSUBS 1.11462f
C138 VP.n82 VSUBS 0.038323f
C139 B.n0 VSUBS 0.007769f
C140 B.n1 VSUBS 0.007769f
C141 B.n2 VSUBS 0.01149f
C142 B.n3 VSUBS 0.008805f
C143 B.n4 VSUBS 0.008805f
C144 B.n5 VSUBS 0.008805f
C145 B.n6 VSUBS 0.008805f
C146 B.n7 VSUBS 0.008805f
C147 B.n8 VSUBS 0.008805f
C148 B.n9 VSUBS 0.008805f
C149 B.n10 VSUBS 0.008805f
C150 B.n11 VSUBS 0.008805f
C151 B.n12 VSUBS 0.008805f
C152 B.n13 VSUBS 0.008805f
C153 B.n14 VSUBS 0.008805f
C154 B.n15 VSUBS 0.008805f
C155 B.n16 VSUBS 0.008805f
C156 B.n17 VSUBS 0.008805f
C157 B.n18 VSUBS 0.008805f
C158 B.n19 VSUBS 0.008805f
C159 B.n20 VSUBS 0.008805f
C160 B.n21 VSUBS 0.008805f
C161 B.n22 VSUBS 0.008805f
C162 B.n23 VSUBS 0.008805f
C163 B.n24 VSUBS 0.008805f
C164 B.n25 VSUBS 0.008805f
C165 B.n26 VSUBS 0.008805f
C166 B.n27 VSUBS 0.008805f
C167 B.n28 VSUBS 0.02161f
C168 B.n29 VSUBS 0.008805f
C169 B.n30 VSUBS 0.008805f
C170 B.n31 VSUBS 0.008805f
C171 B.n32 VSUBS 0.008805f
C172 B.n33 VSUBS 0.008805f
C173 B.n34 VSUBS 0.008805f
C174 B.n35 VSUBS 0.008805f
C175 B.n36 VSUBS 0.008805f
C176 B.n37 VSUBS 0.008805f
C177 B.n38 VSUBS 0.008805f
C178 B.n39 VSUBS 0.008805f
C179 B.n40 VSUBS 0.008805f
C180 B.n41 VSUBS 0.008805f
C181 B.n42 VSUBS 0.008805f
C182 B.n43 VSUBS 0.008805f
C183 B.n44 VSUBS 0.008805f
C184 B.n45 VSUBS 0.008805f
C185 B.n46 VSUBS 0.008805f
C186 B.n47 VSUBS 0.008805f
C187 B.n48 VSUBS 0.008805f
C188 B.n49 VSUBS 0.008805f
C189 B.n50 VSUBS 0.008805f
C190 B.n51 VSUBS 0.008805f
C191 B.n52 VSUBS 0.008805f
C192 B.n53 VSUBS 0.008805f
C193 B.t4 VSUBS 0.635387f
C194 B.t5 VSUBS 0.659138f
C195 B.t3 VSUBS 1.90489f
C196 B.n54 VSUBS 0.335796f
C197 B.n55 VSUBS 0.088712f
C198 B.n56 VSUBS 0.0204f
C199 B.n57 VSUBS 0.008805f
C200 B.n58 VSUBS 0.008805f
C201 B.n59 VSUBS 0.008805f
C202 B.n60 VSUBS 0.008805f
C203 B.n61 VSUBS 0.008805f
C204 B.t7 VSUBS 0.635369f
C205 B.t8 VSUBS 0.659122f
C206 B.t6 VSUBS 1.90489f
C207 B.n62 VSUBS 0.335812f
C208 B.n63 VSUBS 0.08873f
C209 B.n64 VSUBS 0.008805f
C210 B.n65 VSUBS 0.008805f
C211 B.n66 VSUBS 0.008805f
C212 B.n67 VSUBS 0.008805f
C213 B.n68 VSUBS 0.008805f
C214 B.n69 VSUBS 0.008805f
C215 B.n70 VSUBS 0.008805f
C216 B.n71 VSUBS 0.008805f
C217 B.n72 VSUBS 0.008805f
C218 B.n73 VSUBS 0.008805f
C219 B.n74 VSUBS 0.008805f
C220 B.n75 VSUBS 0.008805f
C221 B.n76 VSUBS 0.008805f
C222 B.n77 VSUBS 0.008805f
C223 B.n78 VSUBS 0.008805f
C224 B.n79 VSUBS 0.008805f
C225 B.n80 VSUBS 0.008805f
C226 B.n81 VSUBS 0.008805f
C227 B.n82 VSUBS 0.008805f
C228 B.n83 VSUBS 0.008805f
C229 B.n84 VSUBS 0.008805f
C230 B.n85 VSUBS 0.008805f
C231 B.n86 VSUBS 0.008805f
C232 B.n87 VSUBS 0.008805f
C233 B.n88 VSUBS 0.022415f
C234 B.n89 VSUBS 0.008805f
C235 B.n90 VSUBS 0.008805f
C236 B.n91 VSUBS 0.008805f
C237 B.n92 VSUBS 0.008805f
C238 B.n93 VSUBS 0.008805f
C239 B.n94 VSUBS 0.008805f
C240 B.n95 VSUBS 0.008805f
C241 B.n96 VSUBS 0.008805f
C242 B.n97 VSUBS 0.008805f
C243 B.n98 VSUBS 0.008805f
C244 B.n99 VSUBS 0.008805f
C245 B.n100 VSUBS 0.008805f
C246 B.n101 VSUBS 0.008805f
C247 B.n102 VSUBS 0.008805f
C248 B.n103 VSUBS 0.008805f
C249 B.n104 VSUBS 0.008805f
C250 B.n105 VSUBS 0.008805f
C251 B.n106 VSUBS 0.008805f
C252 B.n107 VSUBS 0.008805f
C253 B.n108 VSUBS 0.008805f
C254 B.n109 VSUBS 0.008805f
C255 B.n110 VSUBS 0.008805f
C256 B.n111 VSUBS 0.008805f
C257 B.n112 VSUBS 0.008805f
C258 B.n113 VSUBS 0.008805f
C259 B.n114 VSUBS 0.008805f
C260 B.n115 VSUBS 0.008805f
C261 B.n116 VSUBS 0.008805f
C262 B.n117 VSUBS 0.008805f
C263 B.n118 VSUBS 0.008805f
C264 B.n119 VSUBS 0.008805f
C265 B.n120 VSUBS 0.008805f
C266 B.n121 VSUBS 0.008805f
C267 B.n122 VSUBS 0.008805f
C268 B.n123 VSUBS 0.008805f
C269 B.n124 VSUBS 0.008805f
C270 B.n125 VSUBS 0.008805f
C271 B.n126 VSUBS 0.008805f
C272 B.n127 VSUBS 0.008805f
C273 B.n128 VSUBS 0.008805f
C274 B.n129 VSUBS 0.008805f
C275 B.n130 VSUBS 0.008805f
C276 B.n131 VSUBS 0.008805f
C277 B.n132 VSUBS 0.008805f
C278 B.n133 VSUBS 0.008805f
C279 B.n134 VSUBS 0.008805f
C280 B.n135 VSUBS 0.008805f
C281 B.n136 VSUBS 0.008805f
C282 B.n137 VSUBS 0.008805f
C283 B.n138 VSUBS 0.008805f
C284 B.n139 VSUBS 0.008805f
C285 B.n140 VSUBS 0.008805f
C286 B.n141 VSUBS 0.008805f
C287 B.n142 VSUBS 0.022553f
C288 B.n143 VSUBS 0.008805f
C289 B.n144 VSUBS 0.008805f
C290 B.n145 VSUBS 0.008805f
C291 B.n146 VSUBS 0.008805f
C292 B.n147 VSUBS 0.008805f
C293 B.n148 VSUBS 0.008805f
C294 B.n149 VSUBS 0.008805f
C295 B.n150 VSUBS 0.008805f
C296 B.n151 VSUBS 0.008805f
C297 B.n152 VSUBS 0.008805f
C298 B.n153 VSUBS 0.008805f
C299 B.n154 VSUBS 0.008805f
C300 B.n155 VSUBS 0.008805f
C301 B.n156 VSUBS 0.008805f
C302 B.n157 VSUBS 0.008805f
C303 B.n158 VSUBS 0.008805f
C304 B.n159 VSUBS 0.008805f
C305 B.n160 VSUBS 0.008805f
C306 B.n161 VSUBS 0.008805f
C307 B.n162 VSUBS 0.008805f
C308 B.n163 VSUBS 0.008805f
C309 B.n164 VSUBS 0.008805f
C310 B.n165 VSUBS 0.008805f
C311 B.n166 VSUBS 0.008805f
C312 B.n167 VSUBS 0.008805f
C313 B.t11 VSUBS 0.635369f
C314 B.t10 VSUBS 0.659122f
C315 B.t9 VSUBS 1.90489f
C316 B.n168 VSUBS 0.335812f
C317 B.n169 VSUBS 0.08873f
C318 B.n170 VSUBS 0.0204f
C319 B.n171 VSUBS 0.008805f
C320 B.n172 VSUBS 0.008805f
C321 B.n173 VSUBS 0.008805f
C322 B.n174 VSUBS 0.008805f
C323 B.n175 VSUBS 0.008805f
C324 B.t2 VSUBS 0.635387f
C325 B.t1 VSUBS 0.659138f
C326 B.t0 VSUBS 1.90489f
C327 B.n176 VSUBS 0.335796f
C328 B.n177 VSUBS 0.088712f
C329 B.n178 VSUBS 0.008805f
C330 B.n179 VSUBS 0.008805f
C331 B.n180 VSUBS 0.008805f
C332 B.n181 VSUBS 0.008805f
C333 B.n182 VSUBS 0.008805f
C334 B.n183 VSUBS 0.008805f
C335 B.n184 VSUBS 0.008805f
C336 B.n185 VSUBS 0.008805f
C337 B.n186 VSUBS 0.008805f
C338 B.n187 VSUBS 0.008805f
C339 B.n188 VSUBS 0.008805f
C340 B.n189 VSUBS 0.008805f
C341 B.n190 VSUBS 0.008805f
C342 B.n191 VSUBS 0.008805f
C343 B.n192 VSUBS 0.008805f
C344 B.n193 VSUBS 0.008805f
C345 B.n194 VSUBS 0.008805f
C346 B.n195 VSUBS 0.008805f
C347 B.n196 VSUBS 0.008805f
C348 B.n197 VSUBS 0.008805f
C349 B.n198 VSUBS 0.008805f
C350 B.n199 VSUBS 0.008805f
C351 B.n200 VSUBS 0.008805f
C352 B.n201 VSUBS 0.008805f
C353 B.n202 VSUBS 0.022415f
C354 B.n203 VSUBS 0.008805f
C355 B.n204 VSUBS 0.008805f
C356 B.n205 VSUBS 0.008805f
C357 B.n206 VSUBS 0.008805f
C358 B.n207 VSUBS 0.008805f
C359 B.n208 VSUBS 0.008805f
C360 B.n209 VSUBS 0.008805f
C361 B.n210 VSUBS 0.008805f
C362 B.n211 VSUBS 0.008805f
C363 B.n212 VSUBS 0.008805f
C364 B.n213 VSUBS 0.008805f
C365 B.n214 VSUBS 0.008805f
C366 B.n215 VSUBS 0.008805f
C367 B.n216 VSUBS 0.008805f
C368 B.n217 VSUBS 0.008805f
C369 B.n218 VSUBS 0.008805f
C370 B.n219 VSUBS 0.008805f
C371 B.n220 VSUBS 0.008805f
C372 B.n221 VSUBS 0.008805f
C373 B.n222 VSUBS 0.008805f
C374 B.n223 VSUBS 0.008805f
C375 B.n224 VSUBS 0.008805f
C376 B.n225 VSUBS 0.008805f
C377 B.n226 VSUBS 0.008805f
C378 B.n227 VSUBS 0.008805f
C379 B.n228 VSUBS 0.008805f
C380 B.n229 VSUBS 0.008805f
C381 B.n230 VSUBS 0.008805f
C382 B.n231 VSUBS 0.008805f
C383 B.n232 VSUBS 0.008805f
C384 B.n233 VSUBS 0.008805f
C385 B.n234 VSUBS 0.008805f
C386 B.n235 VSUBS 0.008805f
C387 B.n236 VSUBS 0.008805f
C388 B.n237 VSUBS 0.008805f
C389 B.n238 VSUBS 0.008805f
C390 B.n239 VSUBS 0.008805f
C391 B.n240 VSUBS 0.008805f
C392 B.n241 VSUBS 0.008805f
C393 B.n242 VSUBS 0.008805f
C394 B.n243 VSUBS 0.008805f
C395 B.n244 VSUBS 0.008805f
C396 B.n245 VSUBS 0.008805f
C397 B.n246 VSUBS 0.008805f
C398 B.n247 VSUBS 0.008805f
C399 B.n248 VSUBS 0.008805f
C400 B.n249 VSUBS 0.008805f
C401 B.n250 VSUBS 0.008805f
C402 B.n251 VSUBS 0.008805f
C403 B.n252 VSUBS 0.008805f
C404 B.n253 VSUBS 0.008805f
C405 B.n254 VSUBS 0.008805f
C406 B.n255 VSUBS 0.008805f
C407 B.n256 VSUBS 0.008805f
C408 B.n257 VSUBS 0.008805f
C409 B.n258 VSUBS 0.008805f
C410 B.n259 VSUBS 0.008805f
C411 B.n260 VSUBS 0.008805f
C412 B.n261 VSUBS 0.008805f
C413 B.n262 VSUBS 0.008805f
C414 B.n263 VSUBS 0.008805f
C415 B.n264 VSUBS 0.008805f
C416 B.n265 VSUBS 0.008805f
C417 B.n266 VSUBS 0.008805f
C418 B.n267 VSUBS 0.008805f
C419 B.n268 VSUBS 0.008805f
C420 B.n269 VSUBS 0.008805f
C421 B.n270 VSUBS 0.008805f
C422 B.n271 VSUBS 0.008805f
C423 B.n272 VSUBS 0.008805f
C424 B.n273 VSUBS 0.008805f
C425 B.n274 VSUBS 0.008805f
C426 B.n275 VSUBS 0.008805f
C427 B.n276 VSUBS 0.008805f
C428 B.n277 VSUBS 0.008805f
C429 B.n278 VSUBS 0.008805f
C430 B.n279 VSUBS 0.008805f
C431 B.n280 VSUBS 0.008805f
C432 B.n281 VSUBS 0.008805f
C433 B.n282 VSUBS 0.008805f
C434 B.n283 VSUBS 0.008805f
C435 B.n284 VSUBS 0.008805f
C436 B.n285 VSUBS 0.008805f
C437 B.n286 VSUBS 0.008805f
C438 B.n287 VSUBS 0.008805f
C439 B.n288 VSUBS 0.008805f
C440 B.n289 VSUBS 0.008805f
C441 B.n290 VSUBS 0.008805f
C442 B.n291 VSUBS 0.008805f
C443 B.n292 VSUBS 0.008805f
C444 B.n293 VSUBS 0.008805f
C445 B.n294 VSUBS 0.008805f
C446 B.n295 VSUBS 0.008805f
C447 B.n296 VSUBS 0.008805f
C448 B.n297 VSUBS 0.008805f
C449 B.n298 VSUBS 0.008805f
C450 B.n299 VSUBS 0.008805f
C451 B.n300 VSUBS 0.008805f
C452 B.n301 VSUBS 0.008805f
C453 B.n302 VSUBS 0.008805f
C454 B.n303 VSUBS 0.008805f
C455 B.n304 VSUBS 0.008805f
C456 B.n305 VSUBS 0.02161f
C457 B.n306 VSUBS 0.02161f
C458 B.n307 VSUBS 0.022415f
C459 B.n308 VSUBS 0.008805f
C460 B.n309 VSUBS 0.008805f
C461 B.n310 VSUBS 0.008805f
C462 B.n311 VSUBS 0.008805f
C463 B.n312 VSUBS 0.008805f
C464 B.n313 VSUBS 0.008805f
C465 B.n314 VSUBS 0.008805f
C466 B.n315 VSUBS 0.008805f
C467 B.n316 VSUBS 0.008805f
C468 B.n317 VSUBS 0.008805f
C469 B.n318 VSUBS 0.008805f
C470 B.n319 VSUBS 0.008805f
C471 B.n320 VSUBS 0.008805f
C472 B.n321 VSUBS 0.008805f
C473 B.n322 VSUBS 0.008805f
C474 B.n323 VSUBS 0.008805f
C475 B.n324 VSUBS 0.008805f
C476 B.n325 VSUBS 0.008805f
C477 B.n326 VSUBS 0.008805f
C478 B.n327 VSUBS 0.008805f
C479 B.n328 VSUBS 0.008805f
C480 B.n329 VSUBS 0.008805f
C481 B.n330 VSUBS 0.008805f
C482 B.n331 VSUBS 0.008805f
C483 B.n332 VSUBS 0.008805f
C484 B.n333 VSUBS 0.008805f
C485 B.n334 VSUBS 0.008805f
C486 B.n335 VSUBS 0.008805f
C487 B.n336 VSUBS 0.008805f
C488 B.n337 VSUBS 0.008805f
C489 B.n338 VSUBS 0.008805f
C490 B.n339 VSUBS 0.008805f
C491 B.n340 VSUBS 0.008805f
C492 B.n341 VSUBS 0.008805f
C493 B.n342 VSUBS 0.008805f
C494 B.n343 VSUBS 0.008805f
C495 B.n344 VSUBS 0.008805f
C496 B.n345 VSUBS 0.008805f
C497 B.n346 VSUBS 0.008805f
C498 B.n347 VSUBS 0.008805f
C499 B.n348 VSUBS 0.008805f
C500 B.n349 VSUBS 0.008805f
C501 B.n350 VSUBS 0.008805f
C502 B.n351 VSUBS 0.008805f
C503 B.n352 VSUBS 0.008805f
C504 B.n353 VSUBS 0.008805f
C505 B.n354 VSUBS 0.008805f
C506 B.n355 VSUBS 0.008805f
C507 B.n356 VSUBS 0.008805f
C508 B.n357 VSUBS 0.008805f
C509 B.n358 VSUBS 0.008805f
C510 B.n359 VSUBS 0.008805f
C511 B.n360 VSUBS 0.008805f
C512 B.n361 VSUBS 0.008805f
C513 B.n362 VSUBS 0.008805f
C514 B.n363 VSUBS 0.008805f
C515 B.n364 VSUBS 0.008805f
C516 B.n365 VSUBS 0.008805f
C517 B.n366 VSUBS 0.008805f
C518 B.n367 VSUBS 0.008805f
C519 B.n368 VSUBS 0.008805f
C520 B.n369 VSUBS 0.008805f
C521 B.n370 VSUBS 0.008805f
C522 B.n371 VSUBS 0.008805f
C523 B.n372 VSUBS 0.008805f
C524 B.n373 VSUBS 0.008805f
C525 B.n374 VSUBS 0.008805f
C526 B.n375 VSUBS 0.008805f
C527 B.n376 VSUBS 0.008805f
C528 B.n377 VSUBS 0.008805f
C529 B.n378 VSUBS 0.008805f
C530 B.n379 VSUBS 0.008805f
C531 B.n380 VSUBS 0.008805f
C532 B.n381 VSUBS 0.008805f
C533 B.n382 VSUBS 0.006086f
C534 B.n383 VSUBS 0.0204f
C535 B.n384 VSUBS 0.007122f
C536 B.n385 VSUBS 0.008805f
C537 B.n386 VSUBS 0.008805f
C538 B.n387 VSUBS 0.008805f
C539 B.n388 VSUBS 0.008805f
C540 B.n389 VSUBS 0.008805f
C541 B.n390 VSUBS 0.008805f
C542 B.n391 VSUBS 0.008805f
C543 B.n392 VSUBS 0.008805f
C544 B.n393 VSUBS 0.008805f
C545 B.n394 VSUBS 0.008805f
C546 B.n395 VSUBS 0.008805f
C547 B.n396 VSUBS 0.007122f
C548 B.n397 VSUBS 0.008805f
C549 B.n398 VSUBS 0.008805f
C550 B.n399 VSUBS 0.006086f
C551 B.n400 VSUBS 0.008805f
C552 B.n401 VSUBS 0.008805f
C553 B.n402 VSUBS 0.008805f
C554 B.n403 VSUBS 0.008805f
C555 B.n404 VSUBS 0.008805f
C556 B.n405 VSUBS 0.008805f
C557 B.n406 VSUBS 0.008805f
C558 B.n407 VSUBS 0.008805f
C559 B.n408 VSUBS 0.008805f
C560 B.n409 VSUBS 0.008805f
C561 B.n410 VSUBS 0.008805f
C562 B.n411 VSUBS 0.008805f
C563 B.n412 VSUBS 0.008805f
C564 B.n413 VSUBS 0.008805f
C565 B.n414 VSUBS 0.008805f
C566 B.n415 VSUBS 0.008805f
C567 B.n416 VSUBS 0.008805f
C568 B.n417 VSUBS 0.008805f
C569 B.n418 VSUBS 0.008805f
C570 B.n419 VSUBS 0.008805f
C571 B.n420 VSUBS 0.008805f
C572 B.n421 VSUBS 0.008805f
C573 B.n422 VSUBS 0.008805f
C574 B.n423 VSUBS 0.008805f
C575 B.n424 VSUBS 0.008805f
C576 B.n425 VSUBS 0.008805f
C577 B.n426 VSUBS 0.008805f
C578 B.n427 VSUBS 0.008805f
C579 B.n428 VSUBS 0.008805f
C580 B.n429 VSUBS 0.008805f
C581 B.n430 VSUBS 0.008805f
C582 B.n431 VSUBS 0.008805f
C583 B.n432 VSUBS 0.008805f
C584 B.n433 VSUBS 0.008805f
C585 B.n434 VSUBS 0.008805f
C586 B.n435 VSUBS 0.008805f
C587 B.n436 VSUBS 0.008805f
C588 B.n437 VSUBS 0.008805f
C589 B.n438 VSUBS 0.008805f
C590 B.n439 VSUBS 0.008805f
C591 B.n440 VSUBS 0.008805f
C592 B.n441 VSUBS 0.008805f
C593 B.n442 VSUBS 0.008805f
C594 B.n443 VSUBS 0.008805f
C595 B.n444 VSUBS 0.008805f
C596 B.n445 VSUBS 0.008805f
C597 B.n446 VSUBS 0.008805f
C598 B.n447 VSUBS 0.008805f
C599 B.n448 VSUBS 0.008805f
C600 B.n449 VSUBS 0.008805f
C601 B.n450 VSUBS 0.008805f
C602 B.n451 VSUBS 0.008805f
C603 B.n452 VSUBS 0.008805f
C604 B.n453 VSUBS 0.008805f
C605 B.n454 VSUBS 0.008805f
C606 B.n455 VSUBS 0.008805f
C607 B.n456 VSUBS 0.008805f
C608 B.n457 VSUBS 0.008805f
C609 B.n458 VSUBS 0.008805f
C610 B.n459 VSUBS 0.008805f
C611 B.n460 VSUBS 0.008805f
C612 B.n461 VSUBS 0.008805f
C613 B.n462 VSUBS 0.008805f
C614 B.n463 VSUBS 0.008805f
C615 B.n464 VSUBS 0.008805f
C616 B.n465 VSUBS 0.008805f
C617 B.n466 VSUBS 0.008805f
C618 B.n467 VSUBS 0.008805f
C619 B.n468 VSUBS 0.008805f
C620 B.n469 VSUBS 0.008805f
C621 B.n470 VSUBS 0.008805f
C622 B.n471 VSUBS 0.008805f
C623 B.n472 VSUBS 0.008805f
C624 B.n473 VSUBS 0.021473f
C625 B.n474 VSUBS 0.022415f
C626 B.n475 VSUBS 0.02161f
C627 B.n476 VSUBS 0.008805f
C628 B.n477 VSUBS 0.008805f
C629 B.n478 VSUBS 0.008805f
C630 B.n479 VSUBS 0.008805f
C631 B.n480 VSUBS 0.008805f
C632 B.n481 VSUBS 0.008805f
C633 B.n482 VSUBS 0.008805f
C634 B.n483 VSUBS 0.008805f
C635 B.n484 VSUBS 0.008805f
C636 B.n485 VSUBS 0.008805f
C637 B.n486 VSUBS 0.008805f
C638 B.n487 VSUBS 0.008805f
C639 B.n488 VSUBS 0.008805f
C640 B.n489 VSUBS 0.008805f
C641 B.n490 VSUBS 0.008805f
C642 B.n491 VSUBS 0.008805f
C643 B.n492 VSUBS 0.008805f
C644 B.n493 VSUBS 0.008805f
C645 B.n494 VSUBS 0.008805f
C646 B.n495 VSUBS 0.008805f
C647 B.n496 VSUBS 0.008805f
C648 B.n497 VSUBS 0.008805f
C649 B.n498 VSUBS 0.008805f
C650 B.n499 VSUBS 0.008805f
C651 B.n500 VSUBS 0.008805f
C652 B.n501 VSUBS 0.008805f
C653 B.n502 VSUBS 0.008805f
C654 B.n503 VSUBS 0.008805f
C655 B.n504 VSUBS 0.008805f
C656 B.n505 VSUBS 0.008805f
C657 B.n506 VSUBS 0.008805f
C658 B.n507 VSUBS 0.008805f
C659 B.n508 VSUBS 0.008805f
C660 B.n509 VSUBS 0.008805f
C661 B.n510 VSUBS 0.008805f
C662 B.n511 VSUBS 0.008805f
C663 B.n512 VSUBS 0.008805f
C664 B.n513 VSUBS 0.008805f
C665 B.n514 VSUBS 0.008805f
C666 B.n515 VSUBS 0.008805f
C667 B.n516 VSUBS 0.008805f
C668 B.n517 VSUBS 0.008805f
C669 B.n518 VSUBS 0.008805f
C670 B.n519 VSUBS 0.008805f
C671 B.n520 VSUBS 0.008805f
C672 B.n521 VSUBS 0.008805f
C673 B.n522 VSUBS 0.008805f
C674 B.n523 VSUBS 0.008805f
C675 B.n524 VSUBS 0.008805f
C676 B.n525 VSUBS 0.008805f
C677 B.n526 VSUBS 0.008805f
C678 B.n527 VSUBS 0.008805f
C679 B.n528 VSUBS 0.008805f
C680 B.n529 VSUBS 0.008805f
C681 B.n530 VSUBS 0.008805f
C682 B.n531 VSUBS 0.008805f
C683 B.n532 VSUBS 0.008805f
C684 B.n533 VSUBS 0.008805f
C685 B.n534 VSUBS 0.008805f
C686 B.n535 VSUBS 0.008805f
C687 B.n536 VSUBS 0.008805f
C688 B.n537 VSUBS 0.008805f
C689 B.n538 VSUBS 0.008805f
C690 B.n539 VSUBS 0.008805f
C691 B.n540 VSUBS 0.008805f
C692 B.n541 VSUBS 0.008805f
C693 B.n542 VSUBS 0.008805f
C694 B.n543 VSUBS 0.008805f
C695 B.n544 VSUBS 0.008805f
C696 B.n545 VSUBS 0.008805f
C697 B.n546 VSUBS 0.008805f
C698 B.n547 VSUBS 0.008805f
C699 B.n548 VSUBS 0.008805f
C700 B.n549 VSUBS 0.008805f
C701 B.n550 VSUBS 0.008805f
C702 B.n551 VSUBS 0.008805f
C703 B.n552 VSUBS 0.008805f
C704 B.n553 VSUBS 0.008805f
C705 B.n554 VSUBS 0.008805f
C706 B.n555 VSUBS 0.008805f
C707 B.n556 VSUBS 0.008805f
C708 B.n557 VSUBS 0.008805f
C709 B.n558 VSUBS 0.008805f
C710 B.n559 VSUBS 0.008805f
C711 B.n560 VSUBS 0.008805f
C712 B.n561 VSUBS 0.008805f
C713 B.n562 VSUBS 0.008805f
C714 B.n563 VSUBS 0.008805f
C715 B.n564 VSUBS 0.008805f
C716 B.n565 VSUBS 0.008805f
C717 B.n566 VSUBS 0.008805f
C718 B.n567 VSUBS 0.008805f
C719 B.n568 VSUBS 0.008805f
C720 B.n569 VSUBS 0.008805f
C721 B.n570 VSUBS 0.008805f
C722 B.n571 VSUBS 0.008805f
C723 B.n572 VSUBS 0.008805f
C724 B.n573 VSUBS 0.008805f
C725 B.n574 VSUBS 0.008805f
C726 B.n575 VSUBS 0.008805f
C727 B.n576 VSUBS 0.008805f
C728 B.n577 VSUBS 0.008805f
C729 B.n578 VSUBS 0.008805f
C730 B.n579 VSUBS 0.008805f
C731 B.n580 VSUBS 0.008805f
C732 B.n581 VSUBS 0.008805f
C733 B.n582 VSUBS 0.008805f
C734 B.n583 VSUBS 0.008805f
C735 B.n584 VSUBS 0.008805f
C736 B.n585 VSUBS 0.008805f
C737 B.n586 VSUBS 0.008805f
C738 B.n587 VSUBS 0.008805f
C739 B.n588 VSUBS 0.008805f
C740 B.n589 VSUBS 0.008805f
C741 B.n590 VSUBS 0.008805f
C742 B.n591 VSUBS 0.008805f
C743 B.n592 VSUBS 0.008805f
C744 B.n593 VSUBS 0.008805f
C745 B.n594 VSUBS 0.008805f
C746 B.n595 VSUBS 0.008805f
C747 B.n596 VSUBS 0.008805f
C748 B.n597 VSUBS 0.008805f
C749 B.n598 VSUBS 0.008805f
C750 B.n599 VSUBS 0.008805f
C751 B.n600 VSUBS 0.008805f
C752 B.n601 VSUBS 0.008805f
C753 B.n602 VSUBS 0.008805f
C754 B.n603 VSUBS 0.008805f
C755 B.n604 VSUBS 0.008805f
C756 B.n605 VSUBS 0.008805f
C757 B.n606 VSUBS 0.008805f
C758 B.n607 VSUBS 0.008805f
C759 B.n608 VSUBS 0.008805f
C760 B.n609 VSUBS 0.008805f
C761 B.n610 VSUBS 0.008805f
C762 B.n611 VSUBS 0.008805f
C763 B.n612 VSUBS 0.008805f
C764 B.n613 VSUBS 0.008805f
C765 B.n614 VSUBS 0.008805f
C766 B.n615 VSUBS 0.008805f
C767 B.n616 VSUBS 0.008805f
C768 B.n617 VSUBS 0.008805f
C769 B.n618 VSUBS 0.008805f
C770 B.n619 VSUBS 0.008805f
C771 B.n620 VSUBS 0.008805f
C772 B.n621 VSUBS 0.008805f
C773 B.n622 VSUBS 0.008805f
C774 B.n623 VSUBS 0.008805f
C775 B.n624 VSUBS 0.008805f
C776 B.n625 VSUBS 0.008805f
C777 B.n626 VSUBS 0.008805f
C778 B.n627 VSUBS 0.008805f
C779 B.n628 VSUBS 0.008805f
C780 B.n629 VSUBS 0.008805f
C781 B.n630 VSUBS 0.008805f
C782 B.n631 VSUBS 0.008805f
C783 B.n632 VSUBS 0.008805f
C784 B.n633 VSUBS 0.008805f
C785 B.n634 VSUBS 0.008805f
C786 B.n635 VSUBS 0.02161f
C787 B.n636 VSUBS 0.02161f
C788 B.n637 VSUBS 0.022415f
C789 B.n638 VSUBS 0.008805f
C790 B.n639 VSUBS 0.008805f
C791 B.n640 VSUBS 0.008805f
C792 B.n641 VSUBS 0.008805f
C793 B.n642 VSUBS 0.008805f
C794 B.n643 VSUBS 0.008805f
C795 B.n644 VSUBS 0.008805f
C796 B.n645 VSUBS 0.008805f
C797 B.n646 VSUBS 0.008805f
C798 B.n647 VSUBS 0.008805f
C799 B.n648 VSUBS 0.008805f
C800 B.n649 VSUBS 0.008805f
C801 B.n650 VSUBS 0.008805f
C802 B.n651 VSUBS 0.008805f
C803 B.n652 VSUBS 0.008805f
C804 B.n653 VSUBS 0.008805f
C805 B.n654 VSUBS 0.008805f
C806 B.n655 VSUBS 0.008805f
C807 B.n656 VSUBS 0.008805f
C808 B.n657 VSUBS 0.008805f
C809 B.n658 VSUBS 0.008805f
C810 B.n659 VSUBS 0.008805f
C811 B.n660 VSUBS 0.008805f
C812 B.n661 VSUBS 0.008805f
C813 B.n662 VSUBS 0.008805f
C814 B.n663 VSUBS 0.008805f
C815 B.n664 VSUBS 0.008805f
C816 B.n665 VSUBS 0.008805f
C817 B.n666 VSUBS 0.008805f
C818 B.n667 VSUBS 0.008805f
C819 B.n668 VSUBS 0.008805f
C820 B.n669 VSUBS 0.008805f
C821 B.n670 VSUBS 0.008805f
C822 B.n671 VSUBS 0.008805f
C823 B.n672 VSUBS 0.008805f
C824 B.n673 VSUBS 0.008805f
C825 B.n674 VSUBS 0.008805f
C826 B.n675 VSUBS 0.008805f
C827 B.n676 VSUBS 0.008805f
C828 B.n677 VSUBS 0.008805f
C829 B.n678 VSUBS 0.008805f
C830 B.n679 VSUBS 0.008805f
C831 B.n680 VSUBS 0.008805f
C832 B.n681 VSUBS 0.008805f
C833 B.n682 VSUBS 0.008805f
C834 B.n683 VSUBS 0.008805f
C835 B.n684 VSUBS 0.008805f
C836 B.n685 VSUBS 0.008805f
C837 B.n686 VSUBS 0.008805f
C838 B.n687 VSUBS 0.008805f
C839 B.n688 VSUBS 0.008805f
C840 B.n689 VSUBS 0.008805f
C841 B.n690 VSUBS 0.008805f
C842 B.n691 VSUBS 0.008805f
C843 B.n692 VSUBS 0.008805f
C844 B.n693 VSUBS 0.008805f
C845 B.n694 VSUBS 0.008805f
C846 B.n695 VSUBS 0.008805f
C847 B.n696 VSUBS 0.008805f
C848 B.n697 VSUBS 0.008805f
C849 B.n698 VSUBS 0.008805f
C850 B.n699 VSUBS 0.008805f
C851 B.n700 VSUBS 0.008805f
C852 B.n701 VSUBS 0.008805f
C853 B.n702 VSUBS 0.008805f
C854 B.n703 VSUBS 0.008805f
C855 B.n704 VSUBS 0.008805f
C856 B.n705 VSUBS 0.008805f
C857 B.n706 VSUBS 0.008805f
C858 B.n707 VSUBS 0.008805f
C859 B.n708 VSUBS 0.008805f
C860 B.n709 VSUBS 0.008805f
C861 B.n710 VSUBS 0.008805f
C862 B.n711 VSUBS 0.008805f
C863 B.n712 VSUBS 0.006086f
C864 B.n713 VSUBS 0.0204f
C865 B.n714 VSUBS 0.007122f
C866 B.n715 VSUBS 0.008805f
C867 B.n716 VSUBS 0.008805f
C868 B.n717 VSUBS 0.008805f
C869 B.n718 VSUBS 0.008805f
C870 B.n719 VSUBS 0.008805f
C871 B.n720 VSUBS 0.008805f
C872 B.n721 VSUBS 0.008805f
C873 B.n722 VSUBS 0.008805f
C874 B.n723 VSUBS 0.008805f
C875 B.n724 VSUBS 0.008805f
C876 B.n725 VSUBS 0.008805f
C877 B.n726 VSUBS 0.007122f
C878 B.n727 VSUBS 0.008805f
C879 B.n728 VSUBS 0.008805f
C880 B.n729 VSUBS 0.006086f
C881 B.n730 VSUBS 0.008805f
C882 B.n731 VSUBS 0.008805f
C883 B.n732 VSUBS 0.008805f
C884 B.n733 VSUBS 0.008805f
C885 B.n734 VSUBS 0.008805f
C886 B.n735 VSUBS 0.008805f
C887 B.n736 VSUBS 0.008805f
C888 B.n737 VSUBS 0.008805f
C889 B.n738 VSUBS 0.008805f
C890 B.n739 VSUBS 0.008805f
C891 B.n740 VSUBS 0.008805f
C892 B.n741 VSUBS 0.008805f
C893 B.n742 VSUBS 0.008805f
C894 B.n743 VSUBS 0.008805f
C895 B.n744 VSUBS 0.008805f
C896 B.n745 VSUBS 0.008805f
C897 B.n746 VSUBS 0.008805f
C898 B.n747 VSUBS 0.008805f
C899 B.n748 VSUBS 0.008805f
C900 B.n749 VSUBS 0.008805f
C901 B.n750 VSUBS 0.008805f
C902 B.n751 VSUBS 0.008805f
C903 B.n752 VSUBS 0.008805f
C904 B.n753 VSUBS 0.008805f
C905 B.n754 VSUBS 0.008805f
C906 B.n755 VSUBS 0.008805f
C907 B.n756 VSUBS 0.008805f
C908 B.n757 VSUBS 0.008805f
C909 B.n758 VSUBS 0.008805f
C910 B.n759 VSUBS 0.008805f
C911 B.n760 VSUBS 0.008805f
C912 B.n761 VSUBS 0.008805f
C913 B.n762 VSUBS 0.008805f
C914 B.n763 VSUBS 0.008805f
C915 B.n764 VSUBS 0.008805f
C916 B.n765 VSUBS 0.008805f
C917 B.n766 VSUBS 0.008805f
C918 B.n767 VSUBS 0.008805f
C919 B.n768 VSUBS 0.008805f
C920 B.n769 VSUBS 0.008805f
C921 B.n770 VSUBS 0.008805f
C922 B.n771 VSUBS 0.008805f
C923 B.n772 VSUBS 0.008805f
C924 B.n773 VSUBS 0.008805f
C925 B.n774 VSUBS 0.008805f
C926 B.n775 VSUBS 0.008805f
C927 B.n776 VSUBS 0.008805f
C928 B.n777 VSUBS 0.008805f
C929 B.n778 VSUBS 0.008805f
C930 B.n779 VSUBS 0.008805f
C931 B.n780 VSUBS 0.008805f
C932 B.n781 VSUBS 0.008805f
C933 B.n782 VSUBS 0.008805f
C934 B.n783 VSUBS 0.008805f
C935 B.n784 VSUBS 0.008805f
C936 B.n785 VSUBS 0.008805f
C937 B.n786 VSUBS 0.008805f
C938 B.n787 VSUBS 0.008805f
C939 B.n788 VSUBS 0.008805f
C940 B.n789 VSUBS 0.008805f
C941 B.n790 VSUBS 0.008805f
C942 B.n791 VSUBS 0.008805f
C943 B.n792 VSUBS 0.008805f
C944 B.n793 VSUBS 0.008805f
C945 B.n794 VSUBS 0.008805f
C946 B.n795 VSUBS 0.008805f
C947 B.n796 VSUBS 0.008805f
C948 B.n797 VSUBS 0.008805f
C949 B.n798 VSUBS 0.008805f
C950 B.n799 VSUBS 0.008805f
C951 B.n800 VSUBS 0.008805f
C952 B.n801 VSUBS 0.008805f
C953 B.n802 VSUBS 0.008805f
C954 B.n803 VSUBS 0.022415f
C955 B.n804 VSUBS 0.022415f
C956 B.n805 VSUBS 0.02161f
C957 B.n806 VSUBS 0.008805f
C958 B.n807 VSUBS 0.008805f
C959 B.n808 VSUBS 0.008805f
C960 B.n809 VSUBS 0.008805f
C961 B.n810 VSUBS 0.008805f
C962 B.n811 VSUBS 0.008805f
C963 B.n812 VSUBS 0.008805f
C964 B.n813 VSUBS 0.008805f
C965 B.n814 VSUBS 0.008805f
C966 B.n815 VSUBS 0.008805f
C967 B.n816 VSUBS 0.008805f
C968 B.n817 VSUBS 0.008805f
C969 B.n818 VSUBS 0.008805f
C970 B.n819 VSUBS 0.008805f
C971 B.n820 VSUBS 0.008805f
C972 B.n821 VSUBS 0.008805f
C973 B.n822 VSUBS 0.008805f
C974 B.n823 VSUBS 0.008805f
C975 B.n824 VSUBS 0.008805f
C976 B.n825 VSUBS 0.008805f
C977 B.n826 VSUBS 0.008805f
C978 B.n827 VSUBS 0.008805f
C979 B.n828 VSUBS 0.008805f
C980 B.n829 VSUBS 0.008805f
C981 B.n830 VSUBS 0.008805f
C982 B.n831 VSUBS 0.008805f
C983 B.n832 VSUBS 0.008805f
C984 B.n833 VSUBS 0.008805f
C985 B.n834 VSUBS 0.008805f
C986 B.n835 VSUBS 0.008805f
C987 B.n836 VSUBS 0.008805f
C988 B.n837 VSUBS 0.008805f
C989 B.n838 VSUBS 0.008805f
C990 B.n839 VSUBS 0.008805f
C991 B.n840 VSUBS 0.008805f
C992 B.n841 VSUBS 0.008805f
C993 B.n842 VSUBS 0.008805f
C994 B.n843 VSUBS 0.008805f
C995 B.n844 VSUBS 0.008805f
C996 B.n845 VSUBS 0.008805f
C997 B.n846 VSUBS 0.008805f
C998 B.n847 VSUBS 0.008805f
C999 B.n848 VSUBS 0.008805f
C1000 B.n849 VSUBS 0.008805f
C1001 B.n850 VSUBS 0.008805f
C1002 B.n851 VSUBS 0.008805f
C1003 B.n852 VSUBS 0.008805f
C1004 B.n853 VSUBS 0.008805f
C1005 B.n854 VSUBS 0.008805f
C1006 B.n855 VSUBS 0.008805f
C1007 B.n856 VSUBS 0.008805f
C1008 B.n857 VSUBS 0.008805f
C1009 B.n858 VSUBS 0.008805f
C1010 B.n859 VSUBS 0.008805f
C1011 B.n860 VSUBS 0.008805f
C1012 B.n861 VSUBS 0.008805f
C1013 B.n862 VSUBS 0.008805f
C1014 B.n863 VSUBS 0.008805f
C1015 B.n864 VSUBS 0.008805f
C1016 B.n865 VSUBS 0.008805f
C1017 B.n866 VSUBS 0.008805f
C1018 B.n867 VSUBS 0.008805f
C1019 B.n868 VSUBS 0.008805f
C1020 B.n869 VSUBS 0.008805f
C1021 B.n870 VSUBS 0.008805f
C1022 B.n871 VSUBS 0.008805f
C1023 B.n872 VSUBS 0.008805f
C1024 B.n873 VSUBS 0.008805f
C1025 B.n874 VSUBS 0.008805f
C1026 B.n875 VSUBS 0.008805f
C1027 B.n876 VSUBS 0.008805f
C1028 B.n877 VSUBS 0.008805f
C1029 B.n878 VSUBS 0.008805f
C1030 B.n879 VSUBS 0.008805f
C1031 B.n880 VSUBS 0.008805f
C1032 B.n881 VSUBS 0.008805f
C1033 B.n882 VSUBS 0.008805f
C1034 B.n883 VSUBS 0.01149f
C1035 B.n884 VSUBS 0.01224f
C1036 B.n885 VSUBS 0.02434f
C1037 VDD2.t8 VSUBS 3.4555f
C1038 VDD2.t0 VSUBS 0.323482f
C1039 VDD2.t7 VSUBS 0.323482f
C1040 VDD2.n0 VSUBS 2.641f
C1041 VDD2.n1 VSUBS 1.52182f
C1042 VDD2.t4 VSUBS 0.323482f
C1043 VDD2.t1 VSUBS 0.323482f
C1044 VDD2.n2 VSUBS 2.65924f
C1045 VDD2.n3 VSUBS 3.43184f
C1046 VDD2.t3 VSUBS 3.43266f
C1047 VDD2.n4 VSUBS 3.79176f
C1048 VDD2.t6 VSUBS 0.323482f
C1049 VDD2.t9 VSUBS 0.323482f
C1050 VDD2.n5 VSUBS 2.64101f
C1051 VDD2.n6 VSUBS 0.75264f
C1052 VDD2.t2 VSUBS 0.323482f
C1053 VDD2.t5 VSUBS 0.323482f
C1054 VDD2.n7 VSUBS 2.65919f
C1055 VTAIL.t11 VSUBS 0.332314f
C1056 VTAIL.t8 VSUBS 0.332314f
C1057 VTAIL.n0 VSUBS 2.56246f
C1058 VTAIL.n1 VSUBS 0.928136f
C1059 VTAIL.t16 VSUBS 3.35493f
C1060 VTAIL.n2 VSUBS 1.08648f
C1061 VTAIL.t17 VSUBS 0.332314f
C1062 VTAIL.t1 VSUBS 0.332314f
C1063 VTAIL.n3 VSUBS 2.56246f
C1064 VTAIL.n4 VSUBS 1.03004f
C1065 VTAIL.t19 VSUBS 0.332314f
C1066 VTAIL.t5 VSUBS 0.332314f
C1067 VTAIL.n5 VSUBS 2.56246f
C1068 VTAIL.n6 VSUBS 2.77378f
C1069 VTAIL.t9 VSUBS 0.332314f
C1070 VTAIL.t13 VSUBS 0.332314f
C1071 VTAIL.n7 VSUBS 2.56246f
C1072 VTAIL.n8 VSUBS 2.77378f
C1073 VTAIL.t10 VSUBS 0.332314f
C1074 VTAIL.t6 VSUBS 0.332314f
C1075 VTAIL.n9 VSUBS 2.56246f
C1076 VTAIL.n10 VSUBS 1.03004f
C1077 VTAIL.t15 VSUBS 3.35493f
C1078 VTAIL.n11 VSUBS 1.08647f
C1079 VTAIL.t2 VSUBS 0.332314f
C1080 VTAIL.t4 VSUBS 0.332314f
C1081 VTAIL.n12 VSUBS 2.56246f
C1082 VTAIL.n13 VSUBS 0.97263f
C1083 VTAIL.t3 VSUBS 0.332314f
C1084 VTAIL.t0 VSUBS 0.332314f
C1085 VTAIL.n14 VSUBS 2.56246f
C1086 VTAIL.n15 VSUBS 1.03004f
C1087 VTAIL.t18 VSUBS 3.35493f
C1088 VTAIL.n16 VSUBS 2.68882f
C1089 VTAIL.t7 VSUBS 3.35493f
C1090 VTAIL.n17 VSUBS 2.68882f
C1091 VTAIL.t12 VSUBS 0.332314f
C1092 VTAIL.t14 VSUBS 0.332314f
C1093 VTAIL.n18 VSUBS 2.56246f
C1094 VTAIL.n19 VSUBS 0.87574f
C1095 VN.n0 VSUBS 0.037822f
C1096 VN.t8 VSUBS 2.68221f
C1097 VN.n1 VSUBS 0.028909f
C1098 VN.n2 VSUBS 0.02869f
C1099 VN.t5 VSUBS 2.68221f
C1100 VN.n3 VSUBS 0.055315f
C1101 VN.n4 VSUBS 0.02869f
C1102 VN.t2 VSUBS 2.68221f
C1103 VN.n5 VSUBS 0.940437f
C1104 VN.n6 VSUBS 0.02869f
C1105 VN.n7 VSUBS 0.055315f
C1106 VN.t1 VSUBS 2.87377f
C1107 VN.n8 VSUBS 1.00047f
C1108 VN.t9 VSUBS 2.68221f
C1109 VN.n9 VSUBS 1.01892f
C1110 VN.n10 VSUBS 0.044273f
C1111 VN.n11 VSUBS 0.245291f
C1112 VN.n12 VSUBS 0.02869f
C1113 VN.n13 VSUBS 0.02869f
C1114 VN.n14 VSUBS 0.023762f
C1115 VN.n15 VSUBS 0.057535f
C1116 VN.n16 VSUBS 0.04007f
C1117 VN.n17 VSUBS 0.02869f
C1118 VN.n18 VSUBS 0.02869f
C1119 VN.n19 VSUBS 0.04007f
C1120 VN.n20 VSUBS 0.057535f
C1121 VN.n21 VSUBS 0.023762f
C1122 VN.n22 VSUBS 0.02869f
C1123 VN.n23 VSUBS 0.02869f
C1124 VN.n24 VSUBS 0.02869f
C1125 VN.n25 VSUBS 0.044273f
C1126 VN.n26 VSUBS 0.940437f
C1127 VN.n27 VSUBS 0.035868f
C1128 VN.n28 VSUBS 0.056446f
C1129 VN.n29 VSUBS 0.02869f
C1130 VN.n30 VSUBS 0.02869f
C1131 VN.n31 VSUBS 0.02869f
C1132 VN.n32 VSUBS 0.051258f
C1133 VN.n33 VSUBS 0.048475f
C1134 VN.n34 VSUBS 1.03918f
C1135 VN.n35 VSUBS 0.035729f
C1136 VN.n36 VSUBS 0.037822f
C1137 VN.t6 VSUBS 2.68221f
C1138 VN.n37 VSUBS 0.028909f
C1139 VN.n38 VSUBS 0.02869f
C1140 VN.t3 VSUBS 2.68221f
C1141 VN.n39 VSUBS 0.055315f
C1142 VN.n40 VSUBS 0.02869f
C1143 VN.t0 VSUBS 2.68221f
C1144 VN.n41 VSUBS 0.940437f
C1145 VN.n42 VSUBS 0.02869f
C1146 VN.n43 VSUBS 0.055315f
C1147 VN.t4 VSUBS 2.87377f
C1148 VN.n44 VSUBS 1.00047f
C1149 VN.t7 VSUBS 2.68221f
C1150 VN.n45 VSUBS 1.01892f
C1151 VN.n46 VSUBS 0.044273f
C1152 VN.n47 VSUBS 0.245291f
C1153 VN.n48 VSUBS 0.02869f
C1154 VN.n49 VSUBS 0.02869f
C1155 VN.n50 VSUBS 0.023762f
C1156 VN.n51 VSUBS 0.057535f
C1157 VN.n52 VSUBS 0.04007f
C1158 VN.n53 VSUBS 0.02869f
C1159 VN.n54 VSUBS 0.02869f
C1160 VN.n55 VSUBS 0.04007f
C1161 VN.n56 VSUBS 0.057535f
C1162 VN.n57 VSUBS 0.023762f
C1163 VN.n58 VSUBS 0.02869f
C1164 VN.n59 VSUBS 0.02869f
C1165 VN.n60 VSUBS 0.02869f
C1166 VN.n61 VSUBS 0.044273f
C1167 VN.n62 VSUBS 0.940437f
C1168 VN.n63 VSUBS 0.035868f
C1169 VN.n64 VSUBS 0.056446f
C1170 VN.n65 VSUBS 0.02869f
C1171 VN.n66 VSUBS 0.02869f
C1172 VN.n67 VSUBS 0.02869f
C1173 VN.n68 VSUBS 0.051258f
C1174 VN.n69 VSUBS 0.048475f
C1175 VN.n70 VSUBS 1.03918f
C1176 VN.n71 VSUBS 1.77443f
.ends

