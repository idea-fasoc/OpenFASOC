* NGSPICE file created from diff_pair_sample_1537.ext - technology: sky130A

.subckt diff_pair_sample_1537 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t15 B.t1 sky130_fd_pr__nfet_01v8 ad=0.6468 pd=4.25 as=1.5288 ps=8.62 w=3.92 l=1.8
X1 B.t23 B.t21 B.t22 B.t11 sky130_fd_pr__nfet_01v8 ad=1.5288 pd=8.62 as=0 ps=0 w=3.92 l=1.8
X2 VDD2.t9 VN.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.6468 pd=4.25 as=1.5288 ps=8.62 w=3.92 l=1.8
X3 VDD1.t8 VP.t1 VTAIL.t17 B.t6 sky130_fd_pr__nfet_01v8 ad=1.5288 pd=8.62 as=0.6468 ps=4.25 w=3.92 l=1.8
X4 VTAIL.t7 VN.t1 VDD2.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=0.6468 pd=4.25 as=0.6468 ps=4.25 w=3.92 l=1.8
X5 VTAIL.t11 VP.t2 VDD1.t7 B.t8 sky130_fd_pr__nfet_01v8 ad=0.6468 pd=4.25 as=0.6468 ps=4.25 w=3.92 l=1.8
X6 VDD1.t6 VP.t3 VTAIL.t14 B.t2 sky130_fd_pr__nfet_01v8 ad=1.5288 pd=8.62 as=0.6468 ps=4.25 w=3.92 l=1.8
X7 VDD2.t7 VN.t2 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.6468 pd=4.25 as=0.6468 ps=4.25 w=3.92 l=1.8
X8 VDD2.t6 VN.t3 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=1.5288 pd=8.62 as=0.6468 ps=4.25 w=3.92 l=1.8
X9 B.t20 B.t18 B.t19 B.t15 sky130_fd_pr__nfet_01v8 ad=1.5288 pd=8.62 as=0 ps=0 w=3.92 l=1.8
X10 VDD2.t5 VN.t4 VTAIL.t9 B.t9 sky130_fd_pr__nfet_01v8 ad=0.6468 pd=4.25 as=0.6468 ps=4.25 w=3.92 l=1.8
X11 VTAIL.t12 VP.t4 VDD1.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=0.6468 pd=4.25 as=0.6468 ps=4.25 w=3.92 l=1.8
X12 VDD1.t4 VP.t5 VTAIL.t10 B.t3 sky130_fd_pr__nfet_01v8 ad=0.6468 pd=4.25 as=0.6468 ps=4.25 w=3.92 l=1.8
X13 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=1.5288 pd=8.62 as=0 ps=0 w=3.92 l=1.8
X14 VDD1.t3 VP.t6 VTAIL.t13 B.t0 sky130_fd_pr__nfet_01v8 ad=0.6468 pd=4.25 as=1.5288 ps=8.62 w=3.92 l=1.8
X15 VDD2.t4 VN.t5 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.6468 pd=4.25 as=1.5288 ps=8.62 w=3.92 l=1.8
X16 VTAIL.t16 VP.t7 VDD1.t2 B.t7 sky130_fd_pr__nfet_01v8 ad=0.6468 pd=4.25 as=0.6468 ps=4.25 w=3.92 l=1.8
X17 VTAIL.t8 VN.t6 VDD2.t3 B.t8 sky130_fd_pr__nfet_01v8 ad=0.6468 pd=4.25 as=0.6468 ps=4.25 w=3.92 l=1.8
X18 VTAIL.t18 VP.t8 VDD1.t1 B.t5 sky130_fd_pr__nfet_01v8 ad=0.6468 pd=4.25 as=0.6468 ps=4.25 w=3.92 l=1.8
X19 VDD2.t2 VN.t7 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.5288 pd=8.62 as=0.6468 ps=4.25 w=3.92 l=1.8
X20 VDD1.t0 VP.t9 VTAIL.t19 B.t9 sky130_fd_pr__nfet_01v8 ad=0.6468 pd=4.25 as=0.6468 ps=4.25 w=3.92 l=1.8
X21 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=1.5288 pd=8.62 as=0 ps=0 w=3.92 l=1.8
X22 VTAIL.t4 VN.t8 VDD2.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=0.6468 pd=4.25 as=0.6468 ps=4.25 w=3.92 l=1.8
X23 VTAIL.t5 VN.t9 VDD2.t0 B.t5 sky130_fd_pr__nfet_01v8 ad=0.6468 pd=4.25 as=0.6468 ps=4.25 w=3.92 l=1.8
R0 VP.n42 VP.n9 185.4
R1 VP.n74 VP.n73 185.4
R2 VP.n41 VP.n40 185.4
R3 VP.n19 VP.n16 161.3
R4 VP.n21 VP.n20 161.3
R5 VP.n22 VP.n15 161.3
R6 VP.n24 VP.n23 161.3
R7 VP.n26 VP.n14 161.3
R8 VP.n28 VP.n27 161.3
R9 VP.n29 VP.n13 161.3
R10 VP.n31 VP.n30 161.3
R11 VP.n33 VP.n12 161.3
R12 VP.n35 VP.n34 161.3
R13 VP.n36 VP.n11 161.3
R14 VP.n38 VP.n37 161.3
R15 VP.n39 VP.n10 161.3
R16 VP.n72 VP.n0 161.3
R17 VP.n71 VP.n70 161.3
R18 VP.n69 VP.n1 161.3
R19 VP.n68 VP.n67 161.3
R20 VP.n66 VP.n2 161.3
R21 VP.n64 VP.n63 161.3
R22 VP.n62 VP.n3 161.3
R23 VP.n61 VP.n60 161.3
R24 VP.n59 VP.n4 161.3
R25 VP.n57 VP.n56 161.3
R26 VP.n55 VP.n5 161.3
R27 VP.n54 VP.n53 161.3
R28 VP.n52 VP.n6 161.3
R29 VP.n50 VP.n49 161.3
R30 VP.n48 VP.n7 161.3
R31 VP.n47 VP.n46 161.3
R32 VP.n45 VP.n8 161.3
R33 VP.n44 VP.n43 161.3
R34 VP.n17 VP.t3 84.766
R35 VP.n53 VP.n5 56.5617
R36 VP.n60 VP.n3 56.5617
R37 VP.n27 VP.n13 56.5617
R38 VP.n20 VP.n15 56.5617
R39 VP.n9 VP.t1 52.4849
R40 VP.n51 VP.t8 52.4849
R41 VP.n58 VP.t5 52.4849
R42 VP.n65 VP.t4 52.4849
R43 VP.n73 VP.t0 52.4849
R44 VP.n40 VP.t6 52.4849
R45 VP.n32 VP.t2 52.4849
R46 VP.n25 VP.t9 52.4849
R47 VP.n18 VP.t7 52.4849
R48 VP.n18 VP.n17 51.1748
R49 VP.n46 VP.n7 45.9053
R50 VP.n67 VP.n1 45.9053
R51 VP.n34 VP.n11 45.9053
R52 VP.n42 VP.n41 42.4967
R53 VP.n46 VP.n45 35.2488
R54 VP.n71 VP.n1 35.2488
R55 VP.n38 VP.n11 35.2488
R56 VP.n45 VP.n44 24.5923
R57 VP.n50 VP.n7 24.5923
R58 VP.n53 VP.n52 24.5923
R59 VP.n57 VP.n5 24.5923
R60 VP.n60 VP.n59 24.5923
R61 VP.n64 VP.n3 24.5923
R62 VP.n67 VP.n66 24.5923
R63 VP.n72 VP.n71 24.5923
R64 VP.n39 VP.n38 24.5923
R65 VP.n31 VP.n13 24.5923
R66 VP.n34 VP.n33 24.5923
R67 VP.n24 VP.n15 24.5923
R68 VP.n27 VP.n26 24.5923
R69 VP.n20 VP.n19 24.5923
R70 VP.n52 VP.n51 18.6903
R71 VP.n65 VP.n64 18.6903
R72 VP.n32 VP.n31 18.6903
R73 VP.n19 VP.n18 18.6903
R74 VP.n17 VP.n16 12.512
R75 VP.n58 VP.n57 12.2964
R76 VP.n59 VP.n58 12.2964
R77 VP.n25 VP.n24 12.2964
R78 VP.n26 VP.n25 12.2964
R79 VP.n51 VP.n50 5.90254
R80 VP.n66 VP.n65 5.90254
R81 VP.n33 VP.n32 5.90254
R82 VP.n44 VP.n9 0.492337
R83 VP.n73 VP.n72 0.492337
R84 VP.n40 VP.n39 0.492337
R85 VP.n21 VP.n16 0.189894
R86 VP.n22 VP.n21 0.189894
R87 VP.n23 VP.n22 0.189894
R88 VP.n23 VP.n14 0.189894
R89 VP.n28 VP.n14 0.189894
R90 VP.n29 VP.n28 0.189894
R91 VP.n30 VP.n29 0.189894
R92 VP.n30 VP.n12 0.189894
R93 VP.n35 VP.n12 0.189894
R94 VP.n36 VP.n35 0.189894
R95 VP.n37 VP.n36 0.189894
R96 VP.n37 VP.n10 0.189894
R97 VP.n41 VP.n10 0.189894
R98 VP.n43 VP.n42 0.189894
R99 VP.n43 VP.n8 0.189894
R100 VP.n47 VP.n8 0.189894
R101 VP.n48 VP.n47 0.189894
R102 VP.n49 VP.n48 0.189894
R103 VP.n49 VP.n6 0.189894
R104 VP.n54 VP.n6 0.189894
R105 VP.n55 VP.n54 0.189894
R106 VP.n56 VP.n55 0.189894
R107 VP.n56 VP.n4 0.189894
R108 VP.n61 VP.n4 0.189894
R109 VP.n62 VP.n61 0.189894
R110 VP.n63 VP.n62 0.189894
R111 VP.n63 VP.n2 0.189894
R112 VP.n68 VP.n2 0.189894
R113 VP.n69 VP.n68 0.189894
R114 VP.n70 VP.n69 0.189894
R115 VP.n70 VP.n0 0.189894
R116 VP.n74 VP.n0 0.189894
R117 VP VP.n74 0.0516364
R118 VTAIL.n88 VTAIL.n74 289.615
R119 VTAIL.n16 VTAIL.n2 289.615
R120 VTAIL.n68 VTAIL.n54 289.615
R121 VTAIL.n44 VTAIL.n30 289.615
R122 VTAIL.n81 VTAIL.n80 185
R123 VTAIL.n78 VTAIL.n77 185
R124 VTAIL.n87 VTAIL.n86 185
R125 VTAIL.n89 VTAIL.n88 185
R126 VTAIL.n9 VTAIL.n8 185
R127 VTAIL.n6 VTAIL.n5 185
R128 VTAIL.n15 VTAIL.n14 185
R129 VTAIL.n17 VTAIL.n16 185
R130 VTAIL.n69 VTAIL.n68 185
R131 VTAIL.n67 VTAIL.n66 185
R132 VTAIL.n58 VTAIL.n57 185
R133 VTAIL.n61 VTAIL.n60 185
R134 VTAIL.n45 VTAIL.n44 185
R135 VTAIL.n43 VTAIL.n42 185
R136 VTAIL.n34 VTAIL.n33 185
R137 VTAIL.n37 VTAIL.n36 185
R138 VTAIL.t0 VTAIL.n79 147.888
R139 VTAIL.t15 VTAIL.n7 147.888
R140 VTAIL.t13 VTAIL.n59 147.888
R141 VTAIL.t1 VTAIL.n35 147.888
R142 VTAIL.n80 VTAIL.n77 104.615
R143 VTAIL.n87 VTAIL.n77 104.615
R144 VTAIL.n88 VTAIL.n87 104.615
R145 VTAIL.n8 VTAIL.n5 104.615
R146 VTAIL.n15 VTAIL.n5 104.615
R147 VTAIL.n16 VTAIL.n15 104.615
R148 VTAIL.n68 VTAIL.n67 104.615
R149 VTAIL.n67 VTAIL.n57 104.615
R150 VTAIL.n60 VTAIL.n57 104.615
R151 VTAIL.n44 VTAIL.n43 104.615
R152 VTAIL.n43 VTAIL.n33 104.615
R153 VTAIL.n36 VTAIL.n33 104.615
R154 VTAIL.n53 VTAIL.n52 58.3368
R155 VTAIL.n51 VTAIL.n50 58.3368
R156 VTAIL.n29 VTAIL.n28 58.3368
R157 VTAIL.n27 VTAIL.n26 58.3368
R158 VTAIL.n95 VTAIL.n94 58.3367
R159 VTAIL.n1 VTAIL.n0 58.3367
R160 VTAIL.n23 VTAIL.n22 58.3367
R161 VTAIL.n25 VTAIL.n24 58.3367
R162 VTAIL.n80 VTAIL.t0 52.3082
R163 VTAIL.n8 VTAIL.t15 52.3082
R164 VTAIL.n60 VTAIL.t13 52.3082
R165 VTAIL.n36 VTAIL.t1 52.3082
R166 VTAIL.n93 VTAIL.n92 33.7369
R167 VTAIL.n21 VTAIL.n20 33.7369
R168 VTAIL.n73 VTAIL.n72 33.7369
R169 VTAIL.n49 VTAIL.n48 33.7369
R170 VTAIL.n27 VTAIL.n25 19.4186
R171 VTAIL.n93 VTAIL.n73 17.5824
R172 VTAIL.n81 VTAIL.n79 15.6496
R173 VTAIL.n9 VTAIL.n7 15.6496
R174 VTAIL.n61 VTAIL.n59 15.6496
R175 VTAIL.n37 VTAIL.n35 15.6496
R176 VTAIL.n82 VTAIL.n78 12.8005
R177 VTAIL.n10 VTAIL.n6 12.8005
R178 VTAIL.n62 VTAIL.n58 12.8005
R179 VTAIL.n38 VTAIL.n34 12.8005
R180 VTAIL.n86 VTAIL.n85 12.0247
R181 VTAIL.n14 VTAIL.n13 12.0247
R182 VTAIL.n66 VTAIL.n65 12.0247
R183 VTAIL.n42 VTAIL.n41 12.0247
R184 VTAIL.n89 VTAIL.n76 11.249
R185 VTAIL.n17 VTAIL.n4 11.249
R186 VTAIL.n69 VTAIL.n56 11.249
R187 VTAIL.n45 VTAIL.n32 11.249
R188 VTAIL.n90 VTAIL.n74 10.4732
R189 VTAIL.n18 VTAIL.n2 10.4732
R190 VTAIL.n70 VTAIL.n54 10.4732
R191 VTAIL.n46 VTAIL.n30 10.4732
R192 VTAIL.n92 VTAIL.n91 9.45567
R193 VTAIL.n20 VTAIL.n19 9.45567
R194 VTAIL.n72 VTAIL.n71 9.45567
R195 VTAIL.n48 VTAIL.n47 9.45567
R196 VTAIL.n91 VTAIL.n90 9.3005
R197 VTAIL.n76 VTAIL.n75 9.3005
R198 VTAIL.n85 VTAIL.n84 9.3005
R199 VTAIL.n83 VTAIL.n82 9.3005
R200 VTAIL.n19 VTAIL.n18 9.3005
R201 VTAIL.n4 VTAIL.n3 9.3005
R202 VTAIL.n13 VTAIL.n12 9.3005
R203 VTAIL.n11 VTAIL.n10 9.3005
R204 VTAIL.n71 VTAIL.n70 9.3005
R205 VTAIL.n56 VTAIL.n55 9.3005
R206 VTAIL.n65 VTAIL.n64 9.3005
R207 VTAIL.n63 VTAIL.n62 9.3005
R208 VTAIL.n47 VTAIL.n46 9.3005
R209 VTAIL.n32 VTAIL.n31 9.3005
R210 VTAIL.n41 VTAIL.n40 9.3005
R211 VTAIL.n39 VTAIL.n38 9.3005
R212 VTAIL.n94 VTAIL.t9 5.05152
R213 VTAIL.n94 VTAIL.t8 5.05152
R214 VTAIL.n0 VTAIL.t2 5.05152
R215 VTAIL.n0 VTAIL.t7 5.05152
R216 VTAIL.n22 VTAIL.t10 5.05152
R217 VTAIL.n22 VTAIL.t12 5.05152
R218 VTAIL.n24 VTAIL.t17 5.05152
R219 VTAIL.n24 VTAIL.t18 5.05152
R220 VTAIL.n52 VTAIL.t19 5.05152
R221 VTAIL.n52 VTAIL.t11 5.05152
R222 VTAIL.n50 VTAIL.t14 5.05152
R223 VTAIL.n50 VTAIL.t16 5.05152
R224 VTAIL.n28 VTAIL.t3 5.05152
R225 VTAIL.n28 VTAIL.t4 5.05152
R226 VTAIL.n26 VTAIL.t6 5.05152
R227 VTAIL.n26 VTAIL.t5 5.05152
R228 VTAIL.n83 VTAIL.n79 4.40546
R229 VTAIL.n11 VTAIL.n7 4.40546
R230 VTAIL.n63 VTAIL.n59 4.40546
R231 VTAIL.n39 VTAIL.n35 4.40546
R232 VTAIL.n92 VTAIL.n74 3.49141
R233 VTAIL.n20 VTAIL.n2 3.49141
R234 VTAIL.n72 VTAIL.n54 3.49141
R235 VTAIL.n48 VTAIL.n30 3.49141
R236 VTAIL.n90 VTAIL.n89 2.71565
R237 VTAIL.n18 VTAIL.n17 2.71565
R238 VTAIL.n70 VTAIL.n69 2.71565
R239 VTAIL.n46 VTAIL.n45 2.71565
R240 VTAIL.n86 VTAIL.n76 1.93989
R241 VTAIL.n14 VTAIL.n4 1.93989
R242 VTAIL.n66 VTAIL.n56 1.93989
R243 VTAIL.n42 VTAIL.n32 1.93989
R244 VTAIL.n29 VTAIL.n27 1.83671
R245 VTAIL.n49 VTAIL.n29 1.83671
R246 VTAIL.n53 VTAIL.n51 1.83671
R247 VTAIL.n73 VTAIL.n53 1.83671
R248 VTAIL.n25 VTAIL.n23 1.83671
R249 VTAIL.n23 VTAIL.n21 1.83671
R250 VTAIL.n95 VTAIL.n93 1.83671
R251 VTAIL VTAIL.n1 1.43584
R252 VTAIL.n51 VTAIL.n49 1.38843
R253 VTAIL.n21 VTAIL.n1 1.38843
R254 VTAIL.n85 VTAIL.n78 1.16414
R255 VTAIL.n13 VTAIL.n6 1.16414
R256 VTAIL.n65 VTAIL.n58 1.16414
R257 VTAIL.n41 VTAIL.n34 1.16414
R258 VTAIL VTAIL.n95 0.401362
R259 VTAIL.n82 VTAIL.n81 0.388379
R260 VTAIL.n10 VTAIL.n9 0.388379
R261 VTAIL.n62 VTAIL.n61 0.388379
R262 VTAIL.n38 VTAIL.n37 0.388379
R263 VTAIL.n84 VTAIL.n83 0.155672
R264 VTAIL.n84 VTAIL.n75 0.155672
R265 VTAIL.n91 VTAIL.n75 0.155672
R266 VTAIL.n12 VTAIL.n11 0.155672
R267 VTAIL.n12 VTAIL.n3 0.155672
R268 VTAIL.n19 VTAIL.n3 0.155672
R269 VTAIL.n71 VTAIL.n55 0.155672
R270 VTAIL.n64 VTAIL.n55 0.155672
R271 VTAIL.n64 VTAIL.n63 0.155672
R272 VTAIL.n47 VTAIL.n31 0.155672
R273 VTAIL.n40 VTAIL.n31 0.155672
R274 VTAIL.n40 VTAIL.n39 0.155672
R275 VDD1.n14 VDD1.n0 289.615
R276 VDD1.n35 VDD1.n21 289.615
R277 VDD1.n15 VDD1.n14 185
R278 VDD1.n13 VDD1.n12 185
R279 VDD1.n4 VDD1.n3 185
R280 VDD1.n7 VDD1.n6 185
R281 VDD1.n28 VDD1.n27 185
R282 VDD1.n25 VDD1.n24 185
R283 VDD1.n34 VDD1.n33 185
R284 VDD1.n36 VDD1.n35 185
R285 VDD1.t6 VDD1.n5 147.888
R286 VDD1.t8 VDD1.n26 147.888
R287 VDD1.n14 VDD1.n13 104.615
R288 VDD1.n13 VDD1.n3 104.615
R289 VDD1.n6 VDD1.n3 104.615
R290 VDD1.n27 VDD1.n24 104.615
R291 VDD1.n34 VDD1.n24 104.615
R292 VDD1.n35 VDD1.n34 104.615
R293 VDD1.n43 VDD1.n42 76.3373
R294 VDD1.n20 VDD1.n19 75.0156
R295 VDD1.n45 VDD1.n44 75.0155
R296 VDD1.n41 VDD1.n40 75.0155
R297 VDD1.n6 VDD1.t6 52.3082
R298 VDD1.n27 VDD1.t8 52.3082
R299 VDD1.n20 VDD1.n18 52.2519
R300 VDD1.n41 VDD1.n39 52.2519
R301 VDD1.n45 VDD1.n43 37.3177
R302 VDD1.n7 VDD1.n5 15.6496
R303 VDD1.n28 VDD1.n26 15.6496
R304 VDD1.n8 VDD1.n4 12.8005
R305 VDD1.n29 VDD1.n25 12.8005
R306 VDD1.n12 VDD1.n11 12.0247
R307 VDD1.n33 VDD1.n32 12.0247
R308 VDD1.n15 VDD1.n2 11.249
R309 VDD1.n36 VDD1.n23 11.249
R310 VDD1.n16 VDD1.n0 10.4732
R311 VDD1.n37 VDD1.n21 10.4732
R312 VDD1.n18 VDD1.n17 9.45567
R313 VDD1.n39 VDD1.n38 9.45567
R314 VDD1.n17 VDD1.n16 9.3005
R315 VDD1.n2 VDD1.n1 9.3005
R316 VDD1.n11 VDD1.n10 9.3005
R317 VDD1.n9 VDD1.n8 9.3005
R318 VDD1.n38 VDD1.n37 9.3005
R319 VDD1.n23 VDD1.n22 9.3005
R320 VDD1.n32 VDD1.n31 9.3005
R321 VDD1.n30 VDD1.n29 9.3005
R322 VDD1.n44 VDD1.t7 5.05152
R323 VDD1.n44 VDD1.t3 5.05152
R324 VDD1.n19 VDD1.t2 5.05152
R325 VDD1.n19 VDD1.t0 5.05152
R326 VDD1.n42 VDD1.t5 5.05152
R327 VDD1.n42 VDD1.t9 5.05152
R328 VDD1.n40 VDD1.t1 5.05152
R329 VDD1.n40 VDD1.t4 5.05152
R330 VDD1.n9 VDD1.n5 4.40546
R331 VDD1.n30 VDD1.n26 4.40546
R332 VDD1.n18 VDD1.n0 3.49141
R333 VDD1.n39 VDD1.n21 3.49141
R334 VDD1.n16 VDD1.n15 2.71565
R335 VDD1.n37 VDD1.n36 2.71565
R336 VDD1.n12 VDD1.n2 1.93989
R337 VDD1.n33 VDD1.n23 1.93989
R338 VDD1 VDD1.n45 1.31947
R339 VDD1.n11 VDD1.n4 1.16414
R340 VDD1.n32 VDD1.n25 1.16414
R341 VDD1 VDD1.n20 0.517741
R342 VDD1.n43 VDD1.n41 0.404206
R343 VDD1.n8 VDD1.n7 0.388379
R344 VDD1.n29 VDD1.n28 0.388379
R345 VDD1.n17 VDD1.n1 0.155672
R346 VDD1.n10 VDD1.n1 0.155672
R347 VDD1.n10 VDD1.n9 0.155672
R348 VDD1.n31 VDD1.n30 0.155672
R349 VDD1.n31 VDD1.n22 0.155672
R350 VDD1.n38 VDD1.n22 0.155672
R351 B.n602 B.n601 585
R352 B.n603 B.n602 585
R353 B.n200 B.n107 585
R354 B.n199 B.n198 585
R355 B.n197 B.n196 585
R356 B.n195 B.n194 585
R357 B.n193 B.n192 585
R358 B.n191 B.n190 585
R359 B.n189 B.n188 585
R360 B.n187 B.n186 585
R361 B.n185 B.n184 585
R362 B.n183 B.n182 585
R363 B.n181 B.n180 585
R364 B.n179 B.n178 585
R365 B.n177 B.n176 585
R366 B.n175 B.n174 585
R367 B.n173 B.n172 585
R368 B.n171 B.n170 585
R369 B.n169 B.n168 585
R370 B.n166 B.n165 585
R371 B.n164 B.n163 585
R372 B.n162 B.n161 585
R373 B.n160 B.n159 585
R374 B.n158 B.n157 585
R375 B.n156 B.n155 585
R376 B.n154 B.n153 585
R377 B.n152 B.n151 585
R378 B.n150 B.n149 585
R379 B.n148 B.n147 585
R380 B.n146 B.n145 585
R381 B.n144 B.n143 585
R382 B.n142 B.n141 585
R383 B.n140 B.n139 585
R384 B.n138 B.n137 585
R385 B.n136 B.n135 585
R386 B.n134 B.n133 585
R387 B.n132 B.n131 585
R388 B.n130 B.n129 585
R389 B.n128 B.n127 585
R390 B.n126 B.n125 585
R391 B.n124 B.n123 585
R392 B.n122 B.n121 585
R393 B.n120 B.n119 585
R394 B.n118 B.n117 585
R395 B.n116 B.n115 585
R396 B.n114 B.n113 585
R397 B.n600 B.n84 585
R398 B.n604 B.n84 585
R399 B.n599 B.n83 585
R400 B.n605 B.n83 585
R401 B.n598 B.n597 585
R402 B.n597 B.n79 585
R403 B.n596 B.n78 585
R404 B.n611 B.n78 585
R405 B.n595 B.n77 585
R406 B.n612 B.n77 585
R407 B.n594 B.n76 585
R408 B.n613 B.n76 585
R409 B.n593 B.n592 585
R410 B.n592 B.n75 585
R411 B.n591 B.n71 585
R412 B.n619 B.n71 585
R413 B.n590 B.n70 585
R414 B.n620 B.n70 585
R415 B.n589 B.n69 585
R416 B.n621 B.n69 585
R417 B.n588 B.n587 585
R418 B.n587 B.n65 585
R419 B.n586 B.n64 585
R420 B.n627 B.n64 585
R421 B.n585 B.n63 585
R422 B.n628 B.n63 585
R423 B.n584 B.n62 585
R424 B.n629 B.n62 585
R425 B.n583 B.n582 585
R426 B.n582 B.n58 585
R427 B.n581 B.n57 585
R428 B.n635 B.n57 585
R429 B.n580 B.n56 585
R430 B.n636 B.n56 585
R431 B.n579 B.n55 585
R432 B.n637 B.n55 585
R433 B.n578 B.n577 585
R434 B.n577 B.n51 585
R435 B.n576 B.n50 585
R436 B.n643 B.n50 585
R437 B.n575 B.n49 585
R438 B.n644 B.n49 585
R439 B.n574 B.n48 585
R440 B.n645 B.n48 585
R441 B.n573 B.n572 585
R442 B.n572 B.n44 585
R443 B.n571 B.n43 585
R444 B.n651 B.n43 585
R445 B.n570 B.n42 585
R446 B.n652 B.n42 585
R447 B.n569 B.n41 585
R448 B.n653 B.n41 585
R449 B.n568 B.n567 585
R450 B.n567 B.n37 585
R451 B.n566 B.n36 585
R452 B.n659 B.n36 585
R453 B.n565 B.n35 585
R454 B.n660 B.n35 585
R455 B.n564 B.n34 585
R456 B.n661 B.n34 585
R457 B.n563 B.n562 585
R458 B.n562 B.n30 585
R459 B.n561 B.n29 585
R460 B.n667 B.n29 585
R461 B.n560 B.n28 585
R462 B.n668 B.n28 585
R463 B.n559 B.n27 585
R464 B.n669 B.n27 585
R465 B.n558 B.n557 585
R466 B.n557 B.n26 585
R467 B.n556 B.n22 585
R468 B.n675 B.n22 585
R469 B.n555 B.n21 585
R470 B.n676 B.n21 585
R471 B.n554 B.n20 585
R472 B.n677 B.n20 585
R473 B.n553 B.n552 585
R474 B.n552 B.n16 585
R475 B.n551 B.n15 585
R476 B.n683 B.n15 585
R477 B.n550 B.n14 585
R478 B.n684 B.n14 585
R479 B.n549 B.n13 585
R480 B.n685 B.n13 585
R481 B.n548 B.n547 585
R482 B.n547 B.n12 585
R483 B.n546 B.n545 585
R484 B.n546 B.n8 585
R485 B.n544 B.n7 585
R486 B.n692 B.n7 585
R487 B.n543 B.n6 585
R488 B.n693 B.n6 585
R489 B.n542 B.n5 585
R490 B.n694 B.n5 585
R491 B.n541 B.n540 585
R492 B.n540 B.n4 585
R493 B.n539 B.n201 585
R494 B.n539 B.n538 585
R495 B.n529 B.n202 585
R496 B.n203 B.n202 585
R497 B.n531 B.n530 585
R498 B.n532 B.n531 585
R499 B.n528 B.n207 585
R500 B.n211 B.n207 585
R501 B.n527 B.n526 585
R502 B.n526 B.n525 585
R503 B.n209 B.n208 585
R504 B.n210 B.n209 585
R505 B.n518 B.n517 585
R506 B.n519 B.n518 585
R507 B.n516 B.n216 585
R508 B.n216 B.n215 585
R509 B.n515 B.n514 585
R510 B.n514 B.n513 585
R511 B.n218 B.n217 585
R512 B.n506 B.n218 585
R513 B.n505 B.n504 585
R514 B.n507 B.n505 585
R515 B.n503 B.n223 585
R516 B.n223 B.n222 585
R517 B.n502 B.n501 585
R518 B.n501 B.n500 585
R519 B.n225 B.n224 585
R520 B.n226 B.n225 585
R521 B.n493 B.n492 585
R522 B.n494 B.n493 585
R523 B.n491 B.n230 585
R524 B.n234 B.n230 585
R525 B.n490 B.n489 585
R526 B.n489 B.n488 585
R527 B.n232 B.n231 585
R528 B.n233 B.n232 585
R529 B.n481 B.n480 585
R530 B.n482 B.n481 585
R531 B.n479 B.n239 585
R532 B.n239 B.n238 585
R533 B.n478 B.n477 585
R534 B.n477 B.n476 585
R535 B.n241 B.n240 585
R536 B.n242 B.n241 585
R537 B.n469 B.n468 585
R538 B.n470 B.n469 585
R539 B.n467 B.n247 585
R540 B.n247 B.n246 585
R541 B.n466 B.n465 585
R542 B.n465 B.n464 585
R543 B.n249 B.n248 585
R544 B.n250 B.n249 585
R545 B.n457 B.n456 585
R546 B.n458 B.n457 585
R547 B.n455 B.n255 585
R548 B.n255 B.n254 585
R549 B.n454 B.n453 585
R550 B.n453 B.n452 585
R551 B.n257 B.n256 585
R552 B.n258 B.n257 585
R553 B.n445 B.n444 585
R554 B.n446 B.n445 585
R555 B.n443 B.n263 585
R556 B.n263 B.n262 585
R557 B.n442 B.n441 585
R558 B.n441 B.n440 585
R559 B.n265 B.n264 585
R560 B.n266 B.n265 585
R561 B.n433 B.n432 585
R562 B.n434 B.n433 585
R563 B.n431 B.n271 585
R564 B.n271 B.n270 585
R565 B.n430 B.n429 585
R566 B.n429 B.n428 585
R567 B.n273 B.n272 585
R568 B.n421 B.n273 585
R569 B.n420 B.n419 585
R570 B.n422 B.n420 585
R571 B.n418 B.n278 585
R572 B.n278 B.n277 585
R573 B.n417 B.n416 585
R574 B.n416 B.n415 585
R575 B.n280 B.n279 585
R576 B.n281 B.n280 585
R577 B.n408 B.n407 585
R578 B.n409 B.n408 585
R579 B.n406 B.n286 585
R580 B.n286 B.n285 585
R581 B.n400 B.n399 585
R582 B.n398 B.n310 585
R583 B.n397 B.n309 585
R584 B.n402 B.n309 585
R585 B.n396 B.n395 585
R586 B.n394 B.n393 585
R587 B.n392 B.n391 585
R588 B.n390 B.n389 585
R589 B.n388 B.n387 585
R590 B.n386 B.n385 585
R591 B.n384 B.n383 585
R592 B.n382 B.n381 585
R593 B.n380 B.n379 585
R594 B.n378 B.n377 585
R595 B.n376 B.n375 585
R596 B.n374 B.n373 585
R597 B.n372 B.n371 585
R598 B.n370 B.n369 585
R599 B.n368 B.n367 585
R600 B.n365 B.n364 585
R601 B.n363 B.n362 585
R602 B.n361 B.n360 585
R603 B.n359 B.n358 585
R604 B.n357 B.n356 585
R605 B.n355 B.n354 585
R606 B.n353 B.n352 585
R607 B.n351 B.n350 585
R608 B.n349 B.n348 585
R609 B.n347 B.n346 585
R610 B.n345 B.n344 585
R611 B.n343 B.n342 585
R612 B.n341 B.n340 585
R613 B.n339 B.n338 585
R614 B.n337 B.n336 585
R615 B.n335 B.n334 585
R616 B.n333 B.n332 585
R617 B.n331 B.n330 585
R618 B.n329 B.n328 585
R619 B.n327 B.n326 585
R620 B.n325 B.n324 585
R621 B.n323 B.n322 585
R622 B.n321 B.n320 585
R623 B.n319 B.n318 585
R624 B.n317 B.n316 585
R625 B.n288 B.n287 585
R626 B.n405 B.n404 585
R627 B.n284 B.n283 585
R628 B.n285 B.n284 585
R629 B.n411 B.n410 585
R630 B.n410 B.n409 585
R631 B.n412 B.n282 585
R632 B.n282 B.n281 585
R633 B.n414 B.n413 585
R634 B.n415 B.n414 585
R635 B.n276 B.n275 585
R636 B.n277 B.n276 585
R637 B.n424 B.n423 585
R638 B.n423 B.n422 585
R639 B.n425 B.n274 585
R640 B.n421 B.n274 585
R641 B.n427 B.n426 585
R642 B.n428 B.n427 585
R643 B.n269 B.n268 585
R644 B.n270 B.n269 585
R645 B.n436 B.n435 585
R646 B.n435 B.n434 585
R647 B.n437 B.n267 585
R648 B.n267 B.n266 585
R649 B.n439 B.n438 585
R650 B.n440 B.n439 585
R651 B.n261 B.n260 585
R652 B.n262 B.n261 585
R653 B.n448 B.n447 585
R654 B.n447 B.n446 585
R655 B.n449 B.n259 585
R656 B.n259 B.n258 585
R657 B.n451 B.n450 585
R658 B.n452 B.n451 585
R659 B.n253 B.n252 585
R660 B.n254 B.n253 585
R661 B.n460 B.n459 585
R662 B.n459 B.n458 585
R663 B.n461 B.n251 585
R664 B.n251 B.n250 585
R665 B.n463 B.n462 585
R666 B.n464 B.n463 585
R667 B.n245 B.n244 585
R668 B.n246 B.n245 585
R669 B.n472 B.n471 585
R670 B.n471 B.n470 585
R671 B.n473 B.n243 585
R672 B.n243 B.n242 585
R673 B.n475 B.n474 585
R674 B.n476 B.n475 585
R675 B.n237 B.n236 585
R676 B.n238 B.n237 585
R677 B.n484 B.n483 585
R678 B.n483 B.n482 585
R679 B.n485 B.n235 585
R680 B.n235 B.n233 585
R681 B.n487 B.n486 585
R682 B.n488 B.n487 585
R683 B.n229 B.n228 585
R684 B.n234 B.n229 585
R685 B.n496 B.n495 585
R686 B.n495 B.n494 585
R687 B.n497 B.n227 585
R688 B.n227 B.n226 585
R689 B.n499 B.n498 585
R690 B.n500 B.n499 585
R691 B.n221 B.n220 585
R692 B.n222 B.n221 585
R693 B.n509 B.n508 585
R694 B.n508 B.n507 585
R695 B.n510 B.n219 585
R696 B.n506 B.n219 585
R697 B.n512 B.n511 585
R698 B.n513 B.n512 585
R699 B.n214 B.n213 585
R700 B.n215 B.n214 585
R701 B.n521 B.n520 585
R702 B.n520 B.n519 585
R703 B.n522 B.n212 585
R704 B.n212 B.n210 585
R705 B.n524 B.n523 585
R706 B.n525 B.n524 585
R707 B.n206 B.n205 585
R708 B.n211 B.n206 585
R709 B.n534 B.n533 585
R710 B.n533 B.n532 585
R711 B.n535 B.n204 585
R712 B.n204 B.n203 585
R713 B.n537 B.n536 585
R714 B.n538 B.n537 585
R715 B.n3 B.n0 585
R716 B.n4 B.n3 585
R717 B.n691 B.n1 585
R718 B.n692 B.n691 585
R719 B.n690 B.n689 585
R720 B.n690 B.n8 585
R721 B.n688 B.n9 585
R722 B.n12 B.n9 585
R723 B.n687 B.n686 585
R724 B.n686 B.n685 585
R725 B.n11 B.n10 585
R726 B.n684 B.n11 585
R727 B.n682 B.n681 585
R728 B.n683 B.n682 585
R729 B.n680 B.n17 585
R730 B.n17 B.n16 585
R731 B.n679 B.n678 585
R732 B.n678 B.n677 585
R733 B.n19 B.n18 585
R734 B.n676 B.n19 585
R735 B.n674 B.n673 585
R736 B.n675 B.n674 585
R737 B.n672 B.n23 585
R738 B.n26 B.n23 585
R739 B.n671 B.n670 585
R740 B.n670 B.n669 585
R741 B.n25 B.n24 585
R742 B.n668 B.n25 585
R743 B.n666 B.n665 585
R744 B.n667 B.n666 585
R745 B.n664 B.n31 585
R746 B.n31 B.n30 585
R747 B.n663 B.n662 585
R748 B.n662 B.n661 585
R749 B.n33 B.n32 585
R750 B.n660 B.n33 585
R751 B.n658 B.n657 585
R752 B.n659 B.n658 585
R753 B.n656 B.n38 585
R754 B.n38 B.n37 585
R755 B.n655 B.n654 585
R756 B.n654 B.n653 585
R757 B.n40 B.n39 585
R758 B.n652 B.n40 585
R759 B.n650 B.n649 585
R760 B.n651 B.n650 585
R761 B.n648 B.n45 585
R762 B.n45 B.n44 585
R763 B.n647 B.n646 585
R764 B.n646 B.n645 585
R765 B.n47 B.n46 585
R766 B.n644 B.n47 585
R767 B.n642 B.n641 585
R768 B.n643 B.n642 585
R769 B.n640 B.n52 585
R770 B.n52 B.n51 585
R771 B.n639 B.n638 585
R772 B.n638 B.n637 585
R773 B.n54 B.n53 585
R774 B.n636 B.n54 585
R775 B.n634 B.n633 585
R776 B.n635 B.n634 585
R777 B.n632 B.n59 585
R778 B.n59 B.n58 585
R779 B.n631 B.n630 585
R780 B.n630 B.n629 585
R781 B.n61 B.n60 585
R782 B.n628 B.n61 585
R783 B.n626 B.n625 585
R784 B.n627 B.n626 585
R785 B.n624 B.n66 585
R786 B.n66 B.n65 585
R787 B.n623 B.n622 585
R788 B.n622 B.n621 585
R789 B.n68 B.n67 585
R790 B.n620 B.n68 585
R791 B.n618 B.n617 585
R792 B.n619 B.n618 585
R793 B.n616 B.n72 585
R794 B.n75 B.n72 585
R795 B.n615 B.n614 585
R796 B.n614 B.n613 585
R797 B.n74 B.n73 585
R798 B.n612 B.n74 585
R799 B.n610 B.n609 585
R800 B.n611 B.n610 585
R801 B.n608 B.n80 585
R802 B.n80 B.n79 585
R803 B.n607 B.n606 585
R804 B.n606 B.n605 585
R805 B.n82 B.n81 585
R806 B.n604 B.n82 585
R807 B.n695 B.n694 585
R808 B.n693 B.n2 585
R809 B.n113 B.n82 554.963
R810 B.n602 B.n84 554.963
R811 B.n404 B.n286 554.963
R812 B.n400 B.n284 554.963
R813 B.n110 B.t14 258.89
R814 B.n108 B.t18 258.89
R815 B.n313 B.t21 258.89
R816 B.n311 B.t10 258.89
R817 B.n603 B.n106 256.663
R818 B.n603 B.n105 256.663
R819 B.n603 B.n104 256.663
R820 B.n603 B.n103 256.663
R821 B.n603 B.n102 256.663
R822 B.n603 B.n101 256.663
R823 B.n603 B.n100 256.663
R824 B.n603 B.n99 256.663
R825 B.n603 B.n98 256.663
R826 B.n603 B.n97 256.663
R827 B.n603 B.n96 256.663
R828 B.n603 B.n95 256.663
R829 B.n603 B.n94 256.663
R830 B.n603 B.n93 256.663
R831 B.n603 B.n92 256.663
R832 B.n603 B.n91 256.663
R833 B.n603 B.n90 256.663
R834 B.n603 B.n89 256.663
R835 B.n603 B.n88 256.663
R836 B.n603 B.n87 256.663
R837 B.n603 B.n86 256.663
R838 B.n603 B.n85 256.663
R839 B.n402 B.n401 256.663
R840 B.n402 B.n289 256.663
R841 B.n402 B.n290 256.663
R842 B.n402 B.n291 256.663
R843 B.n402 B.n292 256.663
R844 B.n402 B.n293 256.663
R845 B.n402 B.n294 256.663
R846 B.n402 B.n295 256.663
R847 B.n402 B.n296 256.663
R848 B.n402 B.n297 256.663
R849 B.n402 B.n298 256.663
R850 B.n402 B.n299 256.663
R851 B.n402 B.n300 256.663
R852 B.n402 B.n301 256.663
R853 B.n402 B.n302 256.663
R854 B.n402 B.n303 256.663
R855 B.n402 B.n304 256.663
R856 B.n402 B.n305 256.663
R857 B.n402 B.n306 256.663
R858 B.n402 B.n307 256.663
R859 B.n402 B.n308 256.663
R860 B.n403 B.n402 256.663
R861 B.n697 B.n696 256.663
R862 B.n108 B.t19 185.018
R863 B.n313 B.t23 185.018
R864 B.n110 B.t16 185.018
R865 B.n311 B.t13 185.018
R866 B.n402 B.n285 163.893
R867 B.n604 B.n603 163.893
R868 B.n117 B.n116 163.367
R869 B.n121 B.n120 163.367
R870 B.n125 B.n124 163.367
R871 B.n129 B.n128 163.367
R872 B.n133 B.n132 163.367
R873 B.n137 B.n136 163.367
R874 B.n141 B.n140 163.367
R875 B.n145 B.n144 163.367
R876 B.n149 B.n148 163.367
R877 B.n153 B.n152 163.367
R878 B.n157 B.n156 163.367
R879 B.n161 B.n160 163.367
R880 B.n165 B.n164 163.367
R881 B.n170 B.n169 163.367
R882 B.n174 B.n173 163.367
R883 B.n178 B.n177 163.367
R884 B.n182 B.n181 163.367
R885 B.n186 B.n185 163.367
R886 B.n190 B.n189 163.367
R887 B.n194 B.n193 163.367
R888 B.n198 B.n197 163.367
R889 B.n602 B.n107 163.367
R890 B.n408 B.n286 163.367
R891 B.n408 B.n280 163.367
R892 B.n416 B.n280 163.367
R893 B.n416 B.n278 163.367
R894 B.n420 B.n278 163.367
R895 B.n420 B.n273 163.367
R896 B.n429 B.n273 163.367
R897 B.n429 B.n271 163.367
R898 B.n433 B.n271 163.367
R899 B.n433 B.n265 163.367
R900 B.n441 B.n265 163.367
R901 B.n441 B.n263 163.367
R902 B.n445 B.n263 163.367
R903 B.n445 B.n257 163.367
R904 B.n453 B.n257 163.367
R905 B.n453 B.n255 163.367
R906 B.n457 B.n255 163.367
R907 B.n457 B.n249 163.367
R908 B.n465 B.n249 163.367
R909 B.n465 B.n247 163.367
R910 B.n469 B.n247 163.367
R911 B.n469 B.n241 163.367
R912 B.n477 B.n241 163.367
R913 B.n477 B.n239 163.367
R914 B.n481 B.n239 163.367
R915 B.n481 B.n232 163.367
R916 B.n489 B.n232 163.367
R917 B.n489 B.n230 163.367
R918 B.n493 B.n230 163.367
R919 B.n493 B.n225 163.367
R920 B.n501 B.n225 163.367
R921 B.n501 B.n223 163.367
R922 B.n505 B.n223 163.367
R923 B.n505 B.n218 163.367
R924 B.n514 B.n218 163.367
R925 B.n514 B.n216 163.367
R926 B.n518 B.n216 163.367
R927 B.n518 B.n209 163.367
R928 B.n526 B.n209 163.367
R929 B.n526 B.n207 163.367
R930 B.n531 B.n207 163.367
R931 B.n531 B.n202 163.367
R932 B.n539 B.n202 163.367
R933 B.n540 B.n539 163.367
R934 B.n540 B.n5 163.367
R935 B.n6 B.n5 163.367
R936 B.n7 B.n6 163.367
R937 B.n546 B.n7 163.367
R938 B.n547 B.n546 163.367
R939 B.n547 B.n13 163.367
R940 B.n14 B.n13 163.367
R941 B.n15 B.n14 163.367
R942 B.n552 B.n15 163.367
R943 B.n552 B.n20 163.367
R944 B.n21 B.n20 163.367
R945 B.n22 B.n21 163.367
R946 B.n557 B.n22 163.367
R947 B.n557 B.n27 163.367
R948 B.n28 B.n27 163.367
R949 B.n29 B.n28 163.367
R950 B.n562 B.n29 163.367
R951 B.n562 B.n34 163.367
R952 B.n35 B.n34 163.367
R953 B.n36 B.n35 163.367
R954 B.n567 B.n36 163.367
R955 B.n567 B.n41 163.367
R956 B.n42 B.n41 163.367
R957 B.n43 B.n42 163.367
R958 B.n572 B.n43 163.367
R959 B.n572 B.n48 163.367
R960 B.n49 B.n48 163.367
R961 B.n50 B.n49 163.367
R962 B.n577 B.n50 163.367
R963 B.n577 B.n55 163.367
R964 B.n56 B.n55 163.367
R965 B.n57 B.n56 163.367
R966 B.n582 B.n57 163.367
R967 B.n582 B.n62 163.367
R968 B.n63 B.n62 163.367
R969 B.n64 B.n63 163.367
R970 B.n587 B.n64 163.367
R971 B.n587 B.n69 163.367
R972 B.n70 B.n69 163.367
R973 B.n71 B.n70 163.367
R974 B.n592 B.n71 163.367
R975 B.n592 B.n76 163.367
R976 B.n77 B.n76 163.367
R977 B.n78 B.n77 163.367
R978 B.n597 B.n78 163.367
R979 B.n597 B.n83 163.367
R980 B.n84 B.n83 163.367
R981 B.n310 B.n309 163.367
R982 B.n395 B.n309 163.367
R983 B.n393 B.n392 163.367
R984 B.n389 B.n388 163.367
R985 B.n385 B.n384 163.367
R986 B.n381 B.n380 163.367
R987 B.n377 B.n376 163.367
R988 B.n373 B.n372 163.367
R989 B.n369 B.n368 163.367
R990 B.n364 B.n363 163.367
R991 B.n360 B.n359 163.367
R992 B.n356 B.n355 163.367
R993 B.n352 B.n351 163.367
R994 B.n348 B.n347 163.367
R995 B.n344 B.n343 163.367
R996 B.n340 B.n339 163.367
R997 B.n336 B.n335 163.367
R998 B.n332 B.n331 163.367
R999 B.n328 B.n327 163.367
R1000 B.n324 B.n323 163.367
R1001 B.n320 B.n319 163.367
R1002 B.n316 B.n288 163.367
R1003 B.n410 B.n284 163.367
R1004 B.n410 B.n282 163.367
R1005 B.n414 B.n282 163.367
R1006 B.n414 B.n276 163.367
R1007 B.n423 B.n276 163.367
R1008 B.n423 B.n274 163.367
R1009 B.n427 B.n274 163.367
R1010 B.n427 B.n269 163.367
R1011 B.n435 B.n269 163.367
R1012 B.n435 B.n267 163.367
R1013 B.n439 B.n267 163.367
R1014 B.n439 B.n261 163.367
R1015 B.n447 B.n261 163.367
R1016 B.n447 B.n259 163.367
R1017 B.n451 B.n259 163.367
R1018 B.n451 B.n253 163.367
R1019 B.n459 B.n253 163.367
R1020 B.n459 B.n251 163.367
R1021 B.n463 B.n251 163.367
R1022 B.n463 B.n245 163.367
R1023 B.n471 B.n245 163.367
R1024 B.n471 B.n243 163.367
R1025 B.n475 B.n243 163.367
R1026 B.n475 B.n237 163.367
R1027 B.n483 B.n237 163.367
R1028 B.n483 B.n235 163.367
R1029 B.n487 B.n235 163.367
R1030 B.n487 B.n229 163.367
R1031 B.n495 B.n229 163.367
R1032 B.n495 B.n227 163.367
R1033 B.n499 B.n227 163.367
R1034 B.n499 B.n221 163.367
R1035 B.n508 B.n221 163.367
R1036 B.n508 B.n219 163.367
R1037 B.n512 B.n219 163.367
R1038 B.n512 B.n214 163.367
R1039 B.n520 B.n214 163.367
R1040 B.n520 B.n212 163.367
R1041 B.n524 B.n212 163.367
R1042 B.n524 B.n206 163.367
R1043 B.n533 B.n206 163.367
R1044 B.n533 B.n204 163.367
R1045 B.n537 B.n204 163.367
R1046 B.n537 B.n3 163.367
R1047 B.n695 B.n3 163.367
R1048 B.n691 B.n2 163.367
R1049 B.n691 B.n690 163.367
R1050 B.n690 B.n9 163.367
R1051 B.n686 B.n9 163.367
R1052 B.n686 B.n11 163.367
R1053 B.n682 B.n11 163.367
R1054 B.n682 B.n17 163.367
R1055 B.n678 B.n17 163.367
R1056 B.n678 B.n19 163.367
R1057 B.n674 B.n19 163.367
R1058 B.n674 B.n23 163.367
R1059 B.n670 B.n23 163.367
R1060 B.n670 B.n25 163.367
R1061 B.n666 B.n25 163.367
R1062 B.n666 B.n31 163.367
R1063 B.n662 B.n31 163.367
R1064 B.n662 B.n33 163.367
R1065 B.n658 B.n33 163.367
R1066 B.n658 B.n38 163.367
R1067 B.n654 B.n38 163.367
R1068 B.n654 B.n40 163.367
R1069 B.n650 B.n40 163.367
R1070 B.n650 B.n45 163.367
R1071 B.n646 B.n45 163.367
R1072 B.n646 B.n47 163.367
R1073 B.n642 B.n47 163.367
R1074 B.n642 B.n52 163.367
R1075 B.n638 B.n52 163.367
R1076 B.n638 B.n54 163.367
R1077 B.n634 B.n54 163.367
R1078 B.n634 B.n59 163.367
R1079 B.n630 B.n59 163.367
R1080 B.n630 B.n61 163.367
R1081 B.n626 B.n61 163.367
R1082 B.n626 B.n66 163.367
R1083 B.n622 B.n66 163.367
R1084 B.n622 B.n68 163.367
R1085 B.n618 B.n68 163.367
R1086 B.n618 B.n72 163.367
R1087 B.n614 B.n72 163.367
R1088 B.n614 B.n74 163.367
R1089 B.n610 B.n74 163.367
R1090 B.n610 B.n80 163.367
R1091 B.n606 B.n80 163.367
R1092 B.n606 B.n82 163.367
R1093 B.n109 B.t20 143.708
R1094 B.n314 B.t22 143.708
R1095 B.n111 B.t17 143.708
R1096 B.n312 B.t12 143.708
R1097 B.n409 B.n285 81.3491
R1098 B.n409 B.n281 81.3491
R1099 B.n415 B.n281 81.3491
R1100 B.n415 B.n277 81.3491
R1101 B.n422 B.n277 81.3491
R1102 B.n422 B.n421 81.3491
R1103 B.n428 B.n270 81.3491
R1104 B.n434 B.n270 81.3491
R1105 B.n434 B.n266 81.3491
R1106 B.n440 B.n266 81.3491
R1107 B.n440 B.n262 81.3491
R1108 B.n446 B.n262 81.3491
R1109 B.n446 B.n258 81.3491
R1110 B.n452 B.n258 81.3491
R1111 B.n458 B.n254 81.3491
R1112 B.n458 B.n250 81.3491
R1113 B.n464 B.n250 81.3491
R1114 B.n464 B.n246 81.3491
R1115 B.n470 B.n246 81.3491
R1116 B.n476 B.n242 81.3491
R1117 B.n476 B.n238 81.3491
R1118 B.n482 B.n238 81.3491
R1119 B.n482 B.n233 81.3491
R1120 B.n488 B.n233 81.3491
R1121 B.n488 B.n234 81.3491
R1122 B.n494 B.n226 81.3491
R1123 B.n500 B.n226 81.3491
R1124 B.n500 B.n222 81.3491
R1125 B.n507 B.n222 81.3491
R1126 B.n507 B.n506 81.3491
R1127 B.n513 B.n215 81.3491
R1128 B.n519 B.n215 81.3491
R1129 B.n519 B.n210 81.3491
R1130 B.n525 B.n210 81.3491
R1131 B.n525 B.n211 81.3491
R1132 B.n532 B.n203 81.3491
R1133 B.n538 B.n203 81.3491
R1134 B.n538 B.n4 81.3491
R1135 B.n694 B.n4 81.3491
R1136 B.n694 B.n693 81.3491
R1137 B.n693 B.n692 81.3491
R1138 B.n692 B.n8 81.3491
R1139 B.n12 B.n8 81.3491
R1140 B.n685 B.n12 81.3491
R1141 B.n684 B.n683 81.3491
R1142 B.n683 B.n16 81.3491
R1143 B.n677 B.n16 81.3491
R1144 B.n677 B.n676 81.3491
R1145 B.n676 B.n675 81.3491
R1146 B.n669 B.n26 81.3491
R1147 B.n669 B.n668 81.3491
R1148 B.n668 B.n667 81.3491
R1149 B.n667 B.n30 81.3491
R1150 B.n661 B.n30 81.3491
R1151 B.n660 B.n659 81.3491
R1152 B.n659 B.n37 81.3491
R1153 B.n653 B.n37 81.3491
R1154 B.n653 B.n652 81.3491
R1155 B.n652 B.n651 81.3491
R1156 B.n651 B.n44 81.3491
R1157 B.n645 B.n644 81.3491
R1158 B.n644 B.n643 81.3491
R1159 B.n643 B.n51 81.3491
R1160 B.n637 B.n51 81.3491
R1161 B.n637 B.n636 81.3491
R1162 B.n635 B.n58 81.3491
R1163 B.n629 B.n58 81.3491
R1164 B.n629 B.n628 81.3491
R1165 B.n628 B.n627 81.3491
R1166 B.n627 B.n65 81.3491
R1167 B.n621 B.n65 81.3491
R1168 B.n621 B.n620 81.3491
R1169 B.n620 B.n619 81.3491
R1170 B.n613 B.n75 81.3491
R1171 B.n613 B.n612 81.3491
R1172 B.n612 B.n611 81.3491
R1173 B.n611 B.n79 81.3491
R1174 B.n605 B.n79 81.3491
R1175 B.n605 B.n604 81.3491
R1176 B.n470 B.t5 78.9565
R1177 B.n645 B.t8 78.9565
R1178 B.n113 B.n85 71.676
R1179 B.n117 B.n86 71.676
R1180 B.n121 B.n87 71.676
R1181 B.n125 B.n88 71.676
R1182 B.n129 B.n89 71.676
R1183 B.n133 B.n90 71.676
R1184 B.n137 B.n91 71.676
R1185 B.n141 B.n92 71.676
R1186 B.n145 B.n93 71.676
R1187 B.n149 B.n94 71.676
R1188 B.n153 B.n95 71.676
R1189 B.n157 B.n96 71.676
R1190 B.n161 B.n97 71.676
R1191 B.n165 B.n98 71.676
R1192 B.n170 B.n99 71.676
R1193 B.n174 B.n100 71.676
R1194 B.n178 B.n101 71.676
R1195 B.n182 B.n102 71.676
R1196 B.n186 B.n103 71.676
R1197 B.n190 B.n104 71.676
R1198 B.n194 B.n105 71.676
R1199 B.n198 B.n106 71.676
R1200 B.n107 B.n106 71.676
R1201 B.n197 B.n105 71.676
R1202 B.n193 B.n104 71.676
R1203 B.n189 B.n103 71.676
R1204 B.n185 B.n102 71.676
R1205 B.n181 B.n101 71.676
R1206 B.n177 B.n100 71.676
R1207 B.n173 B.n99 71.676
R1208 B.n169 B.n98 71.676
R1209 B.n164 B.n97 71.676
R1210 B.n160 B.n96 71.676
R1211 B.n156 B.n95 71.676
R1212 B.n152 B.n94 71.676
R1213 B.n148 B.n93 71.676
R1214 B.n144 B.n92 71.676
R1215 B.n140 B.n91 71.676
R1216 B.n136 B.n90 71.676
R1217 B.n132 B.n89 71.676
R1218 B.n128 B.n88 71.676
R1219 B.n124 B.n87 71.676
R1220 B.n120 B.n86 71.676
R1221 B.n116 B.n85 71.676
R1222 B.n401 B.n400 71.676
R1223 B.n395 B.n289 71.676
R1224 B.n392 B.n290 71.676
R1225 B.n388 B.n291 71.676
R1226 B.n384 B.n292 71.676
R1227 B.n380 B.n293 71.676
R1228 B.n376 B.n294 71.676
R1229 B.n372 B.n295 71.676
R1230 B.n368 B.n296 71.676
R1231 B.n363 B.n297 71.676
R1232 B.n359 B.n298 71.676
R1233 B.n355 B.n299 71.676
R1234 B.n351 B.n300 71.676
R1235 B.n347 B.n301 71.676
R1236 B.n343 B.n302 71.676
R1237 B.n339 B.n303 71.676
R1238 B.n335 B.n304 71.676
R1239 B.n331 B.n305 71.676
R1240 B.n327 B.n306 71.676
R1241 B.n323 B.n307 71.676
R1242 B.n319 B.n308 71.676
R1243 B.n403 B.n288 71.676
R1244 B.n401 B.n310 71.676
R1245 B.n393 B.n289 71.676
R1246 B.n389 B.n290 71.676
R1247 B.n385 B.n291 71.676
R1248 B.n381 B.n292 71.676
R1249 B.n377 B.n293 71.676
R1250 B.n373 B.n294 71.676
R1251 B.n369 B.n295 71.676
R1252 B.n364 B.n296 71.676
R1253 B.n360 B.n297 71.676
R1254 B.n356 B.n298 71.676
R1255 B.n352 B.n299 71.676
R1256 B.n348 B.n300 71.676
R1257 B.n344 B.n301 71.676
R1258 B.n340 B.n302 71.676
R1259 B.n336 B.n303 71.676
R1260 B.n332 B.n304 71.676
R1261 B.n328 B.n305 71.676
R1262 B.n324 B.n306 71.676
R1263 B.n320 B.n307 71.676
R1264 B.n316 B.n308 71.676
R1265 B.n404 B.n403 71.676
R1266 B.n696 B.n695 71.676
R1267 B.n696 B.n2 71.676
R1268 B.n428 B.t11 62.2082
R1269 B.n494 B.t3 62.2082
R1270 B.n211 B.t1 62.2082
R1271 B.t2 B.n684 62.2082
R1272 B.n661 B.t9 62.2082
R1273 B.n619 B.t15 62.2082
R1274 B.n112 B.n111 59.5399
R1275 B.n167 B.n109 59.5399
R1276 B.n315 B.n314 59.5399
R1277 B.n366 B.n312 59.5399
R1278 B.n452 B.t6 57.423
R1279 B.t0 B.n635 57.423
R1280 B.n111 B.n110 41.3096
R1281 B.n109 B.n108 41.3096
R1282 B.n314 B.n313 41.3096
R1283 B.n312 B.n311 41.3096
R1284 B.n506 B.t4 40.6748
R1285 B.n513 B.t4 40.6748
R1286 B.n675 B.t7 40.6748
R1287 B.n26 B.t7 40.6748
R1288 B.n399 B.n283 36.059
R1289 B.n406 B.n405 36.059
R1290 B.n601 B.n600 36.059
R1291 B.n114 B.n81 36.059
R1292 B.t6 B.n254 23.9265
R1293 B.n636 B.t0 23.9265
R1294 B.n421 B.t11 19.1413
R1295 B.n234 B.t3 19.1413
R1296 B.n532 B.t1 19.1413
R1297 B.n685 B.t2 19.1413
R1298 B.t9 B.n660 19.1413
R1299 B.n75 B.t15 19.1413
R1300 B B.n697 18.0485
R1301 B.n411 B.n283 10.6151
R1302 B.n412 B.n411 10.6151
R1303 B.n413 B.n412 10.6151
R1304 B.n413 B.n275 10.6151
R1305 B.n424 B.n275 10.6151
R1306 B.n425 B.n424 10.6151
R1307 B.n426 B.n425 10.6151
R1308 B.n426 B.n268 10.6151
R1309 B.n436 B.n268 10.6151
R1310 B.n437 B.n436 10.6151
R1311 B.n438 B.n437 10.6151
R1312 B.n438 B.n260 10.6151
R1313 B.n448 B.n260 10.6151
R1314 B.n449 B.n448 10.6151
R1315 B.n450 B.n449 10.6151
R1316 B.n450 B.n252 10.6151
R1317 B.n460 B.n252 10.6151
R1318 B.n461 B.n460 10.6151
R1319 B.n462 B.n461 10.6151
R1320 B.n462 B.n244 10.6151
R1321 B.n472 B.n244 10.6151
R1322 B.n473 B.n472 10.6151
R1323 B.n474 B.n473 10.6151
R1324 B.n474 B.n236 10.6151
R1325 B.n484 B.n236 10.6151
R1326 B.n485 B.n484 10.6151
R1327 B.n486 B.n485 10.6151
R1328 B.n486 B.n228 10.6151
R1329 B.n496 B.n228 10.6151
R1330 B.n497 B.n496 10.6151
R1331 B.n498 B.n497 10.6151
R1332 B.n498 B.n220 10.6151
R1333 B.n509 B.n220 10.6151
R1334 B.n510 B.n509 10.6151
R1335 B.n511 B.n510 10.6151
R1336 B.n511 B.n213 10.6151
R1337 B.n521 B.n213 10.6151
R1338 B.n522 B.n521 10.6151
R1339 B.n523 B.n522 10.6151
R1340 B.n523 B.n205 10.6151
R1341 B.n534 B.n205 10.6151
R1342 B.n535 B.n534 10.6151
R1343 B.n536 B.n535 10.6151
R1344 B.n536 B.n0 10.6151
R1345 B.n399 B.n398 10.6151
R1346 B.n398 B.n397 10.6151
R1347 B.n397 B.n396 10.6151
R1348 B.n396 B.n394 10.6151
R1349 B.n394 B.n391 10.6151
R1350 B.n391 B.n390 10.6151
R1351 B.n390 B.n387 10.6151
R1352 B.n387 B.n386 10.6151
R1353 B.n386 B.n383 10.6151
R1354 B.n383 B.n382 10.6151
R1355 B.n382 B.n379 10.6151
R1356 B.n379 B.n378 10.6151
R1357 B.n378 B.n375 10.6151
R1358 B.n375 B.n374 10.6151
R1359 B.n374 B.n371 10.6151
R1360 B.n371 B.n370 10.6151
R1361 B.n370 B.n367 10.6151
R1362 B.n365 B.n362 10.6151
R1363 B.n362 B.n361 10.6151
R1364 B.n361 B.n358 10.6151
R1365 B.n358 B.n357 10.6151
R1366 B.n357 B.n354 10.6151
R1367 B.n354 B.n353 10.6151
R1368 B.n353 B.n350 10.6151
R1369 B.n350 B.n349 10.6151
R1370 B.n346 B.n345 10.6151
R1371 B.n345 B.n342 10.6151
R1372 B.n342 B.n341 10.6151
R1373 B.n341 B.n338 10.6151
R1374 B.n338 B.n337 10.6151
R1375 B.n337 B.n334 10.6151
R1376 B.n334 B.n333 10.6151
R1377 B.n333 B.n330 10.6151
R1378 B.n330 B.n329 10.6151
R1379 B.n329 B.n326 10.6151
R1380 B.n326 B.n325 10.6151
R1381 B.n325 B.n322 10.6151
R1382 B.n322 B.n321 10.6151
R1383 B.n321 B.n318 10.6151
R1384 B.n318 B.n317 10.6151
R1385 B.n317 B.n287 10.6151
R1386 B.n405 B.n287 10.6151
R1387 B.n407 B.n406 10.6151
R1388 B.n407 B.n279 10.6151
R1389 B.n417 B.n279 10.6151
R1390 B.n418 B.n417 10.6151
R1391 B.n419 B.n418 10.6151
R1392 B.n419 B.n272 10.6151
R1393 B.n430 B.n272 10.6151
R1394 B.n431 B.n430 10.6151
R1395 B.n432 B.n431 10.6151
R1396 B.n432 B.n264 10.6151
R1397 B.n442 B.n264 10.6151
R1398 B.n443 B.n442 10.6151
R1399 B.n444 B.n443 10.6151
R1400 B.n444 B.n256 10.6151
R1401 B.n454 B.n256 10.6151
R1402 B.n455 B.n454 10.6151
R1403 B.n456 B.n455 10.6151
R1404 B.n456 B.n248 10.6151
R1405 B.n466 B.n248 10.6151
R1406 B.n467 B.n466 10.6151
R1407 B.n468 B.n467 10.6151
R1408 B.n468 B.n240 10.6151
R1409 B.n478 B.n240 10.6151
R1410 B.n479 B.n478 10.6151
R1411 B.n480 B.n479 10.6151
R1412 B.n480 B.n231 10.6151
R1413 B.n490 B.n231 10.6151
R1414 B.n491 B.n490 10.6151
R1415 B.n492 B.n491 10.6151
R1416 B.n492 B.n224 10.6151
R1417 B.n502 B.n224 10.6151
R1418 B.n503 B.n502 10.6151
R1419 B.n504 B.n503 10.6151
R1420 B.n504 B.n217 10.6151
R1421 B.n515 B.n217 10.6151
R1422 B.n516 B.n515 10.6151
R1423 B.n517 B.n516 10.6151
R1424 B.n517 B.n208 10.6151
R1425 B.n527 B.n208 10.6151
R1426 B.n528 B.n527 10.6151
R1427 B.n530 B.n528 10.6151
R1428 B.n530 B.n529 10.6151
R1429 B.n529 B.n201 10.6151
R1430 B.n541 B.n201 10.6151
R1431 B.n542 B.n541 10.6151
R1432 B.n543 B.n542 10.6151
R1433 B.n544 B.n543 10.6151
R1434 B.n545 B.n544 10.6151
R1435 B.n548 B.n545 10.6151
R1436 B.n549 B.n548 10.6151
R1437 B.n550 B.n549 10.6151
R1438 B.n551 B.n550 10.6151
R1439 B.n553 B.n551 10.6151
R1440 B.n554 B.n553 10.6151
R1441 B.n555 B.n554 10.6151
R1442 B.n556 B.n555 10.6151
R1443 B.n558 B.n556 10.6151
R1444 B.n559 B.n558 10.6151
R1445 B.n560 B.n559 10.6151
R1446 B.n561 B.n560 10.6151
R1447 B.n563 B.n561 10.6151
R1448 B.n564 B.n563 10.6151
R1449 B.n565 B.n564 10.6151
R1450 B.n566 B.n565 10.6151
R1451 B.n568 B.n566 10.6151
R1452 B.n569 B.n568 10.6151
R1453 B.n570 B.n569 10.6151
R1454 B.n571 B.n570 10.6151
R1455 B.n573 B.n571 10.6151
R1456 B.n574 B.n573 10.6151
R1457 B.n575 B.n574 10.6151
R1458 B.n576 B.n575 10.6151
R1459 B.n578 B.n576 10.6151
R1460 B.n579 B.n578 10.6151
R1461 B.n580 B.n579 10.6151
R1462 B.n581 B.n580 10.6151
R1463 B.n583 B.n581 10.6151
R1464 B.n584 B.n583 10.6151
R1465 B.n585 B.n584 10.6151
R1466 B.n586 B.n585 10.6151
R1467 B.n588 B.n586 10.6151
R1468 B.n589 B.n588 10.6151
R1469 B.n590 B.n589 10.6151
R1470 B.n591 B.n590 10.6151
R1471 B.n593 B.n591 10.6151
R1472 B.n594 B.n593 10.6151
R1473 B.n595 B.n594 10.6151
R1474 B.n596 B.n595 10.6151
R1475 B.n598 B.n596 10.6151
R1476 B.n599 B.n598 10.6151
R1477 B.n600 B.n599 10.6151
R1478 B.n689 B.n1 10.6151
R1479 B.n689 B.n688 10.6151
R1480 B.n688 B.n687 10.6151
R1481 B.n687 B.n10 10.6151
R1482 B.n681 B.n10 10.6151
R1483 B.n681 B.n680 10.6151
R1484 B.n680 B.n679 10.6151
R1485 B.n679 B.n18 10.6151
R1486 B.n673 B.n18 10.6151
R1487 B.n673 B.n672 10.6151
R1488 B.n672 B.n671 10.6151
R1489 B.n671 B.n24 10.6151
R1490 B.n665 B.n24 10.6151
R1491 B.n665 B.n664 10.6151
R1492 B.n664 B.n663 10.6151
R1493 B.n663 B.n32 10.6151
R1494 B.n657 B.n32 10.6151
R1495 B.n657 B.n656 10.6151
R1496 B.n656 B.n655 10.6151
R1497 B.n655 B.n39 10.6151
R1498 B.n649 B.n39 10.6151
R1499 B.n649 B.n648 10.6151
R1500 B.n648 B.n647 10.6151
R1501 B.n647 B.n46 10.6151
R1502 B.n641 B.n46 10.6151
R1503 B.n641 B.n640 10.6151
R1504 B.n640 B.n639 10.6151
R1505 B.n639 B.n53 10.6151
R1506 B.n633 B.n53 10.6151
R1507 B.n633 B.n632 10.6151
R1508 B.n632 B.n631 10.6151
R1509 B.n631 B.n60 10.6151
R1510 B.n625 B.n60 10.6151
R1511 B.n625 B.n624 10.6151
R1512 B.n624 B.n623 10.6151
R1513 B.n623 B.n67 10.6151
R1514 B.n617 B.n67 10.6151
R1515 B.n617 B.n616 10.6151
R1516 B.n616 B.n615 10.6151
R1517 B.n615 B.n73 10.6151
R1518 B.n609 B.n73 10.6151
R1519 B.n609 B.n608 10.6151
R1520 B.n608 B.n607 10.6151
R1521 B.n607 B.n81 10.6151
R1522 B.n115 B.n114 10.6151
R1523 B.n118 B.n115 10.6151
R1524 B.n119 B.n118 10.6151
R1525 B.n122 B.n119 10.6151
R1526 B.n123 B.n122 10.6151
R1527 B.n126 B.n123 10.6151
R1528 B.n127 B.n126 10.6151
R1529 B.n130 B.n127 10.6151
R1530 B.n131 B.n130 10.6151
R1531 B.n134 B.n131 10.6151
R1532 B.n135 B.n134 10.6151
R1533 B.n138 B.n135 10.6151
R1534 B.n139 B.n138 10.6151
R1535 B.n142 B.n139 10.6151
R1536 B.n143 B.n142 10.6151
R1537 B.n146 B.n143 10.6151
R1538 B.n147 B.n146 10.6151
R1539 B.n151 B.n150 10.6151
R1540 B.n154 B.n151 10.6151
R1541 B.n155 B.n154 10.6151
R1542 B.n158 B.n155 10.6151
R1543 B.n159 B.n158 10.6151
R1544 B.n162 B.n159 10.6151
R1545 B.n163 B.n162 10.6151
R1546 B.n166 B.n163 10.6151
R1547 B.n171 B.n168 10.6151
R1548 B.n172 B.n171 10.6151
R1549 B.n175 B.n172 10.6151
R1550 B.n176 B.n175 10.6151
R1551 B.n179 B.n176 10.6151
R1552 B.n180 B.n179 10.6151
R1553 B.n183 B.n180 10.6151
R1554 B.n184 B.n183 10.6151
R1555 B.n187 B.n184 10.6151
R1556 B.n188 B.n187 10.6151
R1557 B.n191 B.n188 10.6151
R1558 B.n192 B.n191 10.6151
R1559 B.n195 B.n192 10.6151
R1560 B.n196 B.n195 10.6151
R1561 B.n199 B.n196 10.6151
R1562 B.n200 B.n199 10.6151
R1563 B.n601 B.n200 10.6151
R1564 B.n697 B.n0 8.11757
R1565 B.n697 B.n1 8.11757
R1566 B.n366 B.n365 6.5566
R1567 B.n349 B.n315 6.5566
R1568 B.n150 B.n112 6.5566
R1569 B.n167 B.n166 6.5566
R1570 B.n367 B.n366 4.05904
R1571 B.n346 B.n315 4.05904
R1572 B.n147 B.n112 4.05904
R1573 B.n168 B.n167 4.05904
R1574 B.t5 B.n242 2.3931
R1575 B.t8 B.n44 2.3931
R1576 VN.n31 VN.n30 185.4
R1577 VN.n63 VN.n62 185.4
R1578 VN.n61 VN.n32 161.3
R1579 VN.n60 VN.n59 161.3
R1580 VN.n58 VN.n33 161.3
R1581 VN.n57 VN.n56 161.3
R1582 VN.n55 VN.n34 161.3
R1583 VN.n53 VN.n52 161.3
R1584 VN.n51 VN.n35 161.3
R1585 VN.n50 VN.n49 161.3
R1586 VN.n48 VN.n36 161.3
R1587 VN.n46 VN.n45 161.3
R1588 VN.n44 VN.n37 161.3
R1589 VN.n43 VN.n42 161.3
R1590 VN.n41 VN.n38 161.3
R1591 VN.n29 VN.n0 161.3
R1592 VN.n28 VN.n27 161.3
R1593 VN.n26 VN.n1 161.3
R1594 VN.n25 VN.n24 161.3
R1595 VN.n23 VN.n2 161.3
R1596 VN.n21 VN.n20 161.3
R1597 VN.n19 VN.n3 161.3
R1598 VN.n18 VN.n17 161.3
R1599 VN.n16 VN.n4 161.3
R1600 VN.n14 VN.n13 161.3
R1601 VN.n12 VN.n5 161.3
R1602 VN.n11 VN.n10 161.3
R1603 VN.n9 VN.n6 161.3
R1604 VN.n7 VN.t7 84.766
R1605 VN.n39 VN.t5 84.766
R1606 VN.n10 VN.n5 56.5617
R1607 VN.n17 VN.n3 56.5617
R1608 VN.n42 VN.n37 56.5617
R1609 VN.n49 VN.n35 56.5617
R1610 VN.n8 VN.t1 52.4849
R1611 VN.n15 VN.t4 52.4849
R1612 VN.n22 VN.t6 52.4849
R1613 VN.n30 VN.t0 52.4849
R1614 VN.n40 VN.t8 52.4849
R1615 VN.n47 VN.t2 52.4849
R1616 VN.n54 VN.t9 52.4849
R1617 VN.n62 VN.t3 52.4849
R1618 VN.n8 VN.n7 51.1748
R1619 VN.n40 VN.n39 51.1748
R1620 VN.n24 VN.n1 45.9053
R1621 VN.n56 VN.n33 45.9053
R1622 VN VN.n63 42.8774
R1623 VN.n28 VN.n1 35.2488
R1624 VN.n60 VN.n33 35.2488
R1625 VN.n10 VN.n9 24.5923
R1626 VN.n14 VN.n5 24.5923
R1627 VN.n17 VN.n16 24.5923
R1628 VN.n21 VN.n3 24.5923
R1629 VN.n24 VN.n23 24.5923
R1630 VN.n29 VN.n28 24.5923
R1631 VN.n42 VN.n41 24.5923
R1632 VN.n49 VN.n48 24.5923
R1633 VN.n46 VN.n37 24.5923
R1634 VN.n56 VN.n55 24.5923
R1635 VN.n53 VN.n35 24.5923
R1636 VN.n61 VN.n60 24.5923
R1637 VN.n9 VN.n8 18.6903
R1638 VN.n22 VN.n21 18.6903
R1639 VN.n41 VN.n40 18.6903
R1640 VN.n54 VN.n53 18.6903
R1641 VN.n39 VN.n38 12.512
R1642 VN.n7 VN.n6 12.512
R1643 VN.n15 VN.n14 12.2964
R1644 VN.n16 VN.n15 12.2964
R1645 VN.n48 VN.n47 12.2964
R1646 VN.n47 VN.n46 12.2964
R1647 VN.n23 VN.n22 5.90254
R1648 VN.n55 VN.n54 5.90254
R1649 VN.n30 VN.n29 0.492337
R1650 VN.n62 VN.n61 0.492337
R1651 VN.n63 VN.n32 0.189894
R1652 VN.n59 VN.n32 0.189894
R1653 VN.n59 VN.n58 0.189894
R1654 VN.n58 VN.n57 0.189894
R1655 VN.n57 VN.n34 0.189894
R1656 VN.n52 VN.n34 0.189894
R1657 VN.n52 VN.n51 0.189894
R1658 VN.n51 VN.n50 0.189894
R1659 VN.n50 VN.n36 0.189894
R1660 VN.n45 VN.n36 0.189894
R1661 VN.n45 VN.n44 0.189894
R1662 VN.n44 VN.n43 0.189894
R1663 VN.n43 VN.n38 0.189894
R1664 VN.n11 VN.n6 0.189894
R1665 VN.n12 VN.n11 0.189894
R1666 VN.n13 VN.n12 0.189894
R1667 VN.n13 VN.n4 0.189894
R1668 VN.n18 VN.n4 0.189894
R1669 VN.n19 VN.n18 0.189894
R1670 VN.n20 VN.n19 0.189894
R1671 VN.n20 VN.n2 0.189894
R1672 VN.n25 VN.n2 0.189894
R1673 VN.n26 VN.n25 0.189894
R1674 VN.n27 VN.n26 0.189894
R1675 VN.n27 VN.n0 0.189894
R1676 VN.n31 VN.n0 0.189894
R1677 VN VN.n31 0.0516364
R1678 VDD2.n37 VDD2.n23 289.615
R1679 VDD2.n14 VDD2.n0 289.615
R1680 VDD2.n38 VDD2.n37 185
R1681 VDD2.n36 VDD2.n35 185
R1682 VDD2.n27 VDD2.n26 185
R1683 VDD2.n30 VDD2.n29 185
R1684 VDD2.n7 VDD2.n6 185
R1685 VDD2.n4 VDD2.n3 185
R1686 VDD2.n13 VDD2.n12 185
R1687 VDD2.n15 VDD2.n14 185
R1688 VDD2.t6 VDD2.n28 147.888
R1689 VDD2.t2 VDD2.n5 147.888
R1690 VDD2.n37 VDD2.n36 104.615
R1691 VDD2.n36 VDD2.n26 104.615
R1692 VDD2.n29 VDD2.n26 104.615
R1693 VDD2.n6 VDD2.n3 104.615
R1694 VDD2.n13 VDD2.n3 104.615
R1695 VDD2.n14 VDD2.n13 104.615
R1696 VDD2.n22 VDD2.n21 76.3373
R1697 VDD2 VDD2.n45 76.3345
R1698 VDD2.n44 VDD2.n43 75.0156
R1699 VDD2.n20 VDD2.n19 75.0155
R1700 VDD2.n29 VDD2.t6 52.3082
R1701 VDD2.n6 VDD2.t2 52.3082
R1702 VDD2.n20 VDD2.n18 52.2519
R1703 VDD2.n42 VDD2.n41 50.4157
R1704 VDD2.n42 VDD2.n22 35.8166
R1705 VDD2.n30 VDD2.n28 15.6496
R1706 VDD2.n7 VDD2.n5 15.6496
R1707 VDD2.n31 VDD2.n27 12.8005
R1708 VDD2.n8 VDD2.n4 12.8005
R1709 VDD2.n35 VDD2.n34 12.0247
R1710 VDD2.n12 VDD2.n11 12.0247
R1711 VDD2.n38 VDD2.n25 11.249
R1712 VDD2.n15 VDD2.n2 11.249
R1713 VDD2.n39 VDD2.n23 10.4732
R1714 VDD2.n16 VDD2.n0 10.4732
R1715 VDD2.n41 VDD2.n40 9.45567
R1716 VDD2.n18 VDD2.n17 9.45567
R1717 VDD2.n40 VDD2.n39 9.3005
R1718 VDD2.n25 VDD2.n24 9.3005
R1719 VDD2.n34 VDD2.n33 9.3005
R1720 VDD2.n32 VDD2.n31 9.3005
R1721 VDD2.n17 VDD2.n16 9.3005
R1722 VDD2.n2 VDD2.n1 9.3005
R1723 VDD2.n11 VDD2.n10 9.3005
R1724 VDD2.n9 VDD2.n8 9.3005
R1725 VDD2.n45 VDD2.t1 5.05152
R1726 VDD2.n45 VDD2.t4 5.05152
R1727 VDD2.n43 VDD2.t0 5.05152
R1728 VDD2.n43 VDD2.t7 5.05152
R1729 VDD2.n21 VDD2.t3 5.05152
R1730 VDD2.n21 VDD2.t9 5.05152
R1731 VDD2.n19 VDD2.t8 5.05152
R1732 VDD2.n19 VDD2.t5 5.05152
R1733 VDD2.n32 VDD2.n28 4.40546
R1734 VDD2.n9 VDD2.n5 4.40546
R1735 VDD2.n41 VDD2.n23 3.49141
R1736 VDD2.n18 VDD2.n0 3.49141
R1737 VDD2.n39 VDD2.n38 2.71565
R1738 VDD2.n16 VDD2.n15 2.71565
R1739 VDD2.n35 VDD2.n25 1.93989
R1740 VDD2.n12 VDD2.n2 1.93989
R1741 VDD2.n44 VDD2.n42 1.83671
R1742 VDD2.n34 VDD2.n27 1.16414
R1743 VDD2.n11 VDD2.n4 1.16414
R1744 VDD2 VDD2.n44 0.517741
R1745 VDD2.n22 VDD2.n20 0.404206
R1746 VDD2.n31 VDD2.n30 0.388379
R1747 VDD2.n8 VDD2.n7 0.388379
R1748 VDD2.n40 VDD2.n24 0.155672
R1749 VDD2.n33 VDD2.n24 0.155672
R1750 VDD2.n33 VDD2.n32 0.155672
R1751 VDD2.n10 VDD2.n9 0.155672
R1752 VDD2.n10 VDD2.n1 0.155672
R1753 VDD2.n17 VDD2.n1 0.155672
C0 VDD1 VN 0.156178f
C1 VTAIL VP 4.36427f
C2 VDD1 VDD2 1.65236f
C3 VTAIL VN 4.35007f
C4 VN VP 5.72448f
C5 VTAIL VDD2 6.09916f
C6 VP VDD2 0.485973f
C7 VTAIL VDD1 6.05208f
C8 VN VDD2 3.52658f
C9 VDD1 VP 3.85355f
C10 VDD2 B 4.81408f
C11 VDD1 B 4.797912f
C12 VTAIL B 4.078586f
C13 VN B 13.524149f
C14 VP B 12.038127f
C15 VDD2.n0 B 0.031524f
C16 VDD2.n1 B 0.022867f
C17 VDD2.n2 B 0.012288f
C18 VDD2.n3 B 0.029043f
C19 VDD2.n4 B 0.01301f
C20 VDD2.n5 B 0.087626f
C21 VDD2.t2 B 0.048154f
C22 VDD2.n6 B 0.021782f
C23 VDD2.n7 B 0.017094f
C24 VDD2.n8 B 0.012288f
C25 VDD2.n9 B 0.323491f
C26 VDD2.n10 B 0.022867f
C27 VDD2.n11 B 0.012288f
C28 VDD2.n12 B 0.01301f
C29 VDD2.n13 B 0.029043f
C30 VDD2.n14 B 0.061782f
C31 VDD2.n15 B 0.01301f
C32 VDD2.n16 B 0.012288f
C33 VDD2.n17 B 0.055354f
C34 VDD2.n18 B 0.056655f
C35 VDD2.t8 B 0.070834f
C36 VDD2.t5 B 0.070834f
C37 VDD2.n19 B 0.554704f
C38 VDD2.n20 B 0.518228f
C39 VDD2.t3 B 0.070834f
C40 VDD2.t9 B 0.070834f
C41 VDD2.n21 B 0.561973f
C42 VDD2.n22 B 1.82206f
C43 VDD2.n23 B 0.031524f
C44 VDD2.n24 B 0.022867f
C45 VDD2.n25 B 0.012288f
C46 VDD2.n26 B 0.029043f
C47 VDD2.n27 B 0.01301f
C48 VDD2.n28 B 0.087626f
C49 VDD2.t6 B 0.048154f
C50 VDD2.n29 B 0.021782f
C51 VDD2.n30 B 0.017094f
C52 VDD2.n31 B 0.012288f
C53 VDD2.n32 B 0.323491f
C54 VDD2.n33 B 0.022867f
C55 VDD2.n34 B 0.012288f
C56 VDD2.n35 B 0.01301f
C57 VDD2.n36 B 0.029043f
C58 VDD2.n37 B 0.061782f
C59 VDD2.n38 B 0.01301f
C60 VDD2.n39 B 0.012288f
C61 VDD2.n40 B 0.055354f
C62 VDD2.n41 B 0.050303f
C63 VDD2.n42 B 1.77706f
C64 VDD2.t0 B 0.070834f
C65 VDD2.t7 B 0.070834f
C66 VDD2.n43 B 0.554707f
C67 VDD2.n44 B 0.350874f
C68 VDD2.t1 B 0.070834f
C69 VDD2.t4 B 0.070834f
C70 VDD2.n45 B 0.561947f
C71 VN.n0 B 0.030785f
C72 VN.t0 B 0.556982f
C73 VN.n1 B 0.026072f
C74 VN.n2 B 0.030785f
C75 VN.t6 B 0.556982f
C76 VN.n3 B 0.039214f
C77 VN.n4 B 0.030785f
C78 VN.t4 B 0.556982f
C79 VN.n5 B 0.050287f
C80 VN.n6 B 0.225168f
C81 VN.t1 B 0.556982f
C82 VN.t7 B 0.699863f
C83 VN.n7 B 0.295349f
C84 VN.n8 B 0.306651f
C85 VN.n9 B 0.050324f
C86 VN.n10 B 0.039214f
C87 VN.n11 B 0.030785f
C88 VN.n12 B 0.030785f
C89 VN.n13 B 0.030785f
C90 VN.n14 B 0.042996f
C91 VN.n15 B 0.231098f
C92 VN.n16 B 0.042996f
C93 VN.n17 B 0.050287f
C94 VN.n18 B 0.030785f
C95 VN.n19 B 0.030785f
C96 VN.n20 B 0.030785f
C97 VN.n21 B 0.050324f
C98 VN.n22 B 0.231098f
C99 VN.n23 B 0.035669f
C100 VN.n24 B 0.058658f
C101 VN.n25 B 0.030785f
C102 VN.n26 B 0.030785f
C103 VN.n27 B 0.030785f
C104 VN.n28 B 0.061859f
C105 VN.n29 B 0.029469f
C106 VN.n30 B 0.295967f
C107 VN.n31 B 0.033549f
C108 VN.n32 B 0.030785f
C109 VN.t3 B 0.556982f
C110 VN.n33 B 0.026072f
C111 VN.n34 B 0.030785f
C112 VN.t9 B 0.556982f
C113 VN.n35 B 0.039214f
C114 VN.n36 B 0.030785f
C115 VN.t2 B 0.556982f
C116 VN.n37 B 0.050287f
C117 VN.n38 B 0.225168f
C118 VN.t8 B 0.556982f
C119 VN.t5 B 0.699863f
C120 VN.n39 B 0.295349f
C121 VN.n40 B 0.306651f
C122 VN.n41 B 0.050324f
C123 VN.n42 B 0.039214f
C124 VN.n43 B 0.030785f
C125 VN.n44 B 0.030785f
C126 VN.n45 B 0.030785f
C127 VN.n46 B 0.042996f
C128 VN.n47 B 0.231098f
C129 VN.n48 B 0.042996f
C130 VN.n49 B 0.050287f
C131 VN.n50 B 0.030785f
C132 VN.n51 B 0.030785f
C133 VN.n52 B 0.030785f
C134 VN.n53 B 0.050324f
C135 VN.n54 B 0.231098f
C136 VN.n55 B 0.035669f
C137 VN.n56 B 0.058658f
C138 VN.n57 B 0.030785f
C139 VN.n58 B 0.030785f
C140 VN.n59 B 0.030785f
C141 VN.n60 B 0.061859f
C142 VN.n61 B 0.029469f
C143 VN.n62 B 0.295967f
C144 VN.n63 B 1.32559f
C145 VDD1.n0 B 0.032551f
C146 VDD1.n1 B 0.023612f
C147 VDD1.n2 B 0.012688f
C148 VDD1.n3 B 0.029989f
C149 VDD1.n4 B 0.013434f
C150 VDD1.n5 B 0.09048f
C151 VDD1.t6 B 0.049723f
C152 VDD1.n6 B 0.022492f
C153 VDD1.n7 B 0.017651f
C154 VDD1.n8 B 0.012688f
C155 VDD1.n9 B 0.334031f
C156 VDD1.n10 B 0.023612f
C157 VDD1.n11 B 0.012688f
C158 VDD1.n12 B 0.013434f
C159 VDD1.n13 B 0.029989f
C160 VDD1.n14 B 0.063795f
C161 VDD1.n15 B 0.013434f
C162 VDD1.n16 B 0.012688f
C163 VDD1.n17 B 0.057157f
C164 VDD1.n18 B 0.058501f
C165 VDD1.t2 B 0.073142f
C166 VDD1.t0 B 0.073142f
C167 VDD1.n19 B 0.572781f
C168 VDD1.n20 B 0.542393f
C169 VDD1.n21 B 0.032551f
C170 VDD1.n22 B 0.023612f
C171 VDD1.n23 B 0.012688f
C172 VDD1.n24 B 0.029989f
C173 VDD1.n25 B 0.013434f
C174 VDD1.n26 B 0.09048f
C175 VDD1.t8 B 0.049723f
C176 VDD1.n27 B 0.022492f
C177 VDD1.n28 B 0.017651f
C178 VDD1.n29 B 0.012688f
C179 VDD1.n30 B 0.334031f
C180 VDD1.n31 B 0.023612f
C181 VDD1.n32 B 0.012688f
C182 VDD1.n33 B 0.013434f
C183 VDD1.n34 B 0.029989f
C184 VDD1.n35 B 0.063795f
C185 VDD1.n36 B 0.013434f
C186 VDD1.n37 B 0.012688f
C187 VDD1.n38 B 0.057157f
C188 VDD1.n39 B 0.058501f
C189 VDD1.t1 B 0.073142f
C190 VDD1.t4 B 0.073142f
C191 VDD1.n40 B 0.572778f
C192 VDD1.n41 B 0.535113f
C193 VDD1.t5 B 0.073142f
C194 VDD1.t9 B 0.073142f
C195 VDD1.n42 B 0.580283f
C196 VDD1.n43 B 1.97408f
C197 VDD1.t7 B 0.073142f
C198 VDD1.t3 B 0.073142f
C199 VDD1.n44 B 0.572778f
C200 VDD1.n45 B 2.07569f
C201 VTAIL.t2 B 0.0933f
C202 VTAIL.t7 B 0.0933f
C203 VTAIL.n0 B 0.66545f
C204 VTAIL.n1 B 0.532022f
C205 VTAIL.n2 B 0.041522f
C206 VTAIL.n3 B 0.030119f
C207 VTAIL.n4 B 0.016185f
C208 VTAIL.n5 B 0.038255f
C209 VTAIL.n6 B 0.017137f
C210 VTAIL.n7 B 0.115418f
C211 VTAIL.t15 B 0.063427f
C212 VTAIL.n8 B 0.028691f
C213 VTAIL.n9 B 0.022515f
C214 VTAIL.n10 B 0.016185f
C215 VTAIL.n11 B 0.426095f
C216 VTAIL.n12 B 0.030119f
C217 VTAIL.n13 B 0.016185f
C218 VTAIL.n14 B 0.017137f
C219 VTAIL.n15 B 0.038255f
C220 VTAIL.n16 B 0.081378f
C221 VTAIL.n17 B 0.017137f
C222 VTAIL.n18 B 0.016185f
C223 VTAIL.n19 B 0.072911f
C224 VTAIL.n20 B 0.045486f
C225 VTAIL.n21 B 0.34049f
C226 VTAIL.t10 B 0.0933f
C227 VTAIL.t12 B 0.0933f
C228 VTAIL.n22 B 0.66545f
C229 VTAIL.n23 B 0.614432f
C230 VTAIL.t17 B 0.0933f
C231 VTAIL.t18 B 0.0933f
C232 VTAIL.n24 B 0.66545f
C233 VTAIL.n25 B 1.52974f
C234 VTAIL.t6 B 0.0933f
C235 VTAIL.t5 B 0.0933f
C236 VTAIL.n26 B 0.665454f
C237 VTAIL.n27 B 1.52973f
C238 VTAIL.t3 B 0.0933f
C239 VTAIL.t4 B 0.0933f
C240 VTAIL.n28 B 0.665454f
C241 VTAIL.n29 B 0.614428f
C242 VTAIL.n30 B 0.041522f
C243 VTAIL.n31 B 0.030119f
C244 VTAIL.n32 B 0.016185f
C245 VTAIL.n33 B 0.038255f
C246 VTAIL.n34 B 0.017137f
C247 VTAIL.n35 B 0.115418f
C248 VTAIL.t1 B 0.063427f
C249 VTAIL.n36 B 0.028691f
C250 VTAIL.n37 B 0.022515f
C251 VTAIL.n38 B 0.016185f
C252 VTAIL.n39 B 0.426095f
C253 VTAIL.n40 B 0.030119f
C254 VTAIL.n41 B 0.016185f
C255 VTAIL.n42 B 0.017137f
C256 VTAIL.n43 B 0.038255f
C257 VTAIL.n44 B 0.081378f
C258 VTAIL.n45 B 0.017137f
C259 VTAIL.n46 B 0.016185f
C260 VTAIL.n47 B 0.072911f
C261 VTAIL.n48 B 0.045486f
C262 VTAIL.n49 B 0.34049f
C263 VTAIL.t14 B 0.0933f
C264 VTAIL.t16 B 0.0933f
C265 VTAIL.n50 B 0.665454f
C266 VTAIL.n51 B 0.570922f
C267 VTAIL.t19 B 0.0933f
C268 VTAIL.t11 B 0.0933f
C269 VTAIL.n52 B 0.665454f
C270 VTAIL.n53 B 0.614428f
C271 VTAIL.n54 B 0.041522f
C272 VTAIL.n55 B 0.030119f
C273 VTAIL.n56 B 0.016185f
C274 VTAIL.n57 B 0.038255f
C275 VTAIL.n58 B 0.017137f
C276 VTAIL.n59 B 0.115418f
C277 VTAIL.t13 B 0.063427f
C278 VTAIL.n60 B 0.028691f
C279 VTAIL.n61 B 0.022515f
C280 VTAIL.n62 B 0.016185f
C281 VTAIL.n63 B 0.426095f
C282 VTAIL.n64 B 0.030119f
C283 VTAIL.n65 B 0.016185f
C284 VTAIL.n66 B 0.017137f
C285 VTAIL.n67 B 0.038255f
C286 VTAIL.n68 B 0.081378f
C287 VTAIL.n69 B 0.017137f
C288 VTAIL.n70 B 0.016185f
C289 VTAIL.n71 B 0.072911f
C290 VTAIL.n72 B 0.045486f
C291 VTAIL.n73 B 1.1211f
C292 VTAIL.n74 B 0.041522f
C293 VTAIL.n75 B 0.030119f
C294 VTAIL.n76 B 0.016185f
C295 VTAIL.n77 B 0.038255f
C296 VTAIL.n78 B 0.017137f
C297 VTAIL.n79 B 0.115418f
C298 VTAIL.t0 B 0.063427f
C299 VTAIL.n80 B 0.028691f
C300 VTAIL.n81 B 0.022515f
C301 VTAIL.n82 B 0.016185f
C302 VTAIL.n83 B 0.426095f
C303 VTAIL.n84 B 0.030119f
C304 VTAIL.n85 B 0.016185f
C305 VTAIL.n86 B 0.017137f
C306 VTAIL.n87 B 0.038255f
C307 VTAIL.n88 B 0.081378f
C308 VTAIL.n89 B 0.017137f
C309 VTAIL.n90 B 0.016185f
C310 VTAIL.n91 B 0.072911f
C311 VTAIL.n92 B 0.045486f
C312 VTAIL.n93 B 1.1211f
C313 VTAIL.t9 B 0.0933f
C314 VTAIL.t8 B 0.0933f
C315 VTAIL.n94 B 0.66545f
C316 VTAIL.n95 B 0.47513f
C317 VP.n0 B 0.031791f
C318 VP.t0 B 0.575194f
C319 VP.n1 B 0.026924f
C320 VP.n2 B 0.031791f
C321 VP.t4 B 0.575194f
C322 VP.n3 B 0.040496f
C323 VP.n4 B 0.031791f
C324 VP.t5 B 0.575194f
C325 VP.n5 B 0.051931f
C326 VP.n6 B 0.031791f
C327 VP.t8 B 0.575194f
C328 VP.n7 B 0.060576f
C329 VP.n8 B 0.031791f
C330 VP.t1 B 0.575194f
C331 VP.n9 B 0.305644f
C332 VP.n10 B 0.031791f
C333 VP.t6 B 0.575194f
C334 VP.n11 B 0.026924f
C335 VP.n12 B 0.031791f
C336 VP.t2 B 0.575194f
C337 VP.n13 B 0.040496f
C338 VP.n14 B 0.031791f
C339 VP.t9 B 0.575194f
C340 VP.n15 B 0.051931f
C341 VP.n16 B 0.23253f
C342 VP.t7 B 0.575194f
C343 VP.t3 B 0.722747f
C344 VP.n17 B 0.305006f
C345 VP.n18 B 0.316678f
C346 VP.n19 B 0.051969f
C347 VP.n20 B 0.040496f
C348 VP.n21 B 0.031791f
C349 VP.n22 B 0.031791f
C350 VP.n23 B 0.031791f
C351 VP.n24 B 0.044402f
C352 VP.n25 B 0.238654f
C353 VP.n26 B 0.044402f
C354 VP.n27 B 0.051931f
C355 VP.n28 B 0.031791f
C356 VP.n29 B 0.031791f
C357 VP.n30 B 0.031791f
C358 VP.n31 B 0.051969f
C359 VP.n32 B 0.238654f
C360 VP.n33 B 0.036835f
C361 VP.n34 B 0.060576f
C362 VP.n35 B 0.031791f
C363 VP.n36 B 0.031791f
C364 VP.n37 B 0.031791f
C365 VP.n38 B 0.063882f
C366 VP.n39 B 0.030432f
C367 VP.n40 B 0.305644f
C368 VP.n41 B 1.34808f
C369 VP.n42 B 1.37505f
C370 VP.n43 B 0.031791f
C371 VP.n44 B 0.030432f
C372 VP.n45 B 0.063882f
C373 VP.n46 B 0.026924f
C374 VP.n47 B 0.031791f
C375 VP.n48 B 0.031791f
C376 VP.n49 B 0.031791f
C377 VP.n50 B 0.036835f
C378 VP.n51 B 0.238654f
C379 VP.n52 B 0.051969f
C380 VP.n53 B 0.040496f
C381 VP.n54 B 0.031791f
C382 VP.n55 B 0.031791f
C383 VP.n56 B 0.031791f
C384 VP.n57 B 0.044402f
C385 VP.n58 B 0.238654f
C386 VP.n59 B 0.044402f
C387 VP.n60 B 0.051931f
C388 VP.n61 B 0.031791f
C389 VP.n62 B 0.031791f
C390 VP.n63 B 0.031791f
C391 VP.n64 B 0.051969f
C392 VP.n65 B 0.238654f
C393 VP.n66 B 0.036835f
C394 VP.n67 B 0.060576f
C395 VP.n68 B 0.031791f
C396 VP.n69 B 0.031791f
C397 VP.n70 B 0.031791f
C398 VP.n71 B 0.063882f
C399 VP.n72 B 0.030432f
C400 VP.n73 B 0.305644f
C401 VP.n74 B 0.034646f
.ends

