* NGSPICE file created from diff_pair_sample_1734.ext - technology: sky130A

.subckt diff_pair_sample_1734 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n3010_n3812# sky130_fd_pr__pfet_01v8 ad=5.5458 pd=29.22 as=0 ps=0 w=14.22 l=1.71
X1 VTAIL.t14 VP.t0 VDD1.t2 w_n3010_n3812# sky130_fd_pr__pfet_01v8 ad=2.3463 pd=14.55 as=2.3463 ps=14.55 w=14.22 l=1.71
X2 VDD2.t7 VN.t0 VTAIL.t1 w_n3010_n3812# sky130_fd_pr__pfet_01v8 ad=2.3463 pd=14.55 as=2.3463 ps=14.55 w=14.22 l=1.71
X3 VTAIL.t6 VN.t1 VDD2.t6 w_n3010_n3812# sky130_fd_pr__pfet_01v8 ad=5.5458 pd=29.22 as=2.3463 ps=14.55 w=14.22 l=1.71
X4 VTAIL.t4 VN.t2 VDD2.t5 w_n3010_n3812# sky130_fd_pr__pfet_01v8 ad=5.5458 pd=29.22 as=2.3463 ps=14.55 w=14.22 l=1.71
X5 VTAIL.t5 VN.t3 VDD2.t4 w_n3010_n3812# sky130_fd_pr__pfet_01v8 ad=2.3463 pd=14.55 as=2.3463 ps=14.55 w=14.22 l=1.71
X6 VDD2.t3 VN.t4 VTAIL.t3 w_n3010_n3812# sky130_fd_pr__pfet_01v8 ad=2.3463 pd=14.55 as=5.5458 ps=29.22 w=14.22 l=1.71
X7 B.t8 B.t6 B.t7 w_n3010_n3812# sky130_fd_pr__pfet_01v8 ad=5.5458 pd=29.22 as=0 ps=0 w=14.22 l=1.71
X8 VDD1.t3 VP.t1 VTAIL.t13 w_n3010_n3812# sky130_fd_pr__pfet_01v8 ad=2.3463 pd=14.55 as=5.5458 ps=29.22 w=14.22 l=1.71
X9 VTAIL.t15 VN.t5 VDD2.t2 w_n3010_n3812# sky130_fd_pr__pfet_01v8 ad=2.3463 pd=14.55 as=2.3463 ps=14.55 w=14.22 l=1.71
X10 B.t5 B.t3 B.t4 w_n3010_n3812# sky130_fd_pr__pfet_01v8 ad=5.5458 pd=29.22 as=0 ps=0 w=14.22 l=1.71
X11 VDD2.t1 VN.t6 VTAIL.t2 w_n3010_n3812# sky130_fd_pr__pfet_01v8 ad=2.3463 pd=14.55 as=5.5458 ps=29.22 w=14.22 l=1.71
X12 VDD1.t6 VP.t2 VTAIL.t12 w_n3010_n3812# sky130_fd_pr__pfet_01v8 ad=2.3463 pd=14.55 as=5.5458 ps=29.22 w=14.22 l=1.71
X13 VTAIL.t11 VP.t3 VDD1.t0 w_n3010_n3812# sky130_fd_pr__pfet_01v8 ad=2.3463 pd=14.55 as=2.3463 ps=14.55 w=14.22 l=1.71
X14 VTAIL.t10 VP.t4 VDD1.t1 w_n3010_n3812# sky130_fd_pr__pfet_01v8 ad=5.5458 pd=29.22 as=2.3463 ps=14.55 w=14.22 l=1.71
X15 VTAIL.t9 VP.t5 VDD1.t7 w_n3010_n3812# sky130_fd_pr__pfet_01v8 ad=5.5458 pd=29.22 as=2.3463 ps=14.55 w=14.22 l=1.71
X16 VDD2.t0 VN.t7 VTAIL.t0 w_n3010_n3812# sky130_fd_pr__pfet_01v8 ad=2.3463 pd=14.55 as=2.3463 ps=14.55 w=14.22 l=1.71
X17 B.t2 B.t0 B.t1 w_n3010_n3812# sky130_fd_pr__pfet_01v8 ad=5.5458 pd=29.22 as=0 ps=0 w=14.22 l=1.71
X18 VDD1.t4 VP.t6 VTAIL.t8 w_n3010_n3812# sky130_fd_pr__pfet_01v8 ad=2.3463 pd=14.55 as=2.3463 ps=14.55 w=14.22 l=1.71
X19 VDD1.t5 VP.t7 VTAIL.t7 w_n3010_n3812# sky130_fd_pr__pfet_01v8 ad=2.3463 pd=14.55 as=2.3463 ps=14.55 w=14.22 l=1.71
R0 B.n525 B.n78 585
R1 B.n527 B.n526 585
R2 B.n528 B.n77 585
R3 B.n530 B.n529 585
R4 B.n531 B.n76 585
R5 B.n533 B.n532 585
R6 B.n534 B.n75 585
R7 B.n536 B.n535 585
R8 B.n537 B.n74 585
R9 B.n539 B.n538 585
R10 B.n540 B.n73 585
R11 B.n542 B.n541 585
R12 B.n543 B.n72 585
R13 B.n545 B.n544 585
R14 B.n546 B.n71 585
R15 B.n548 B.n547 585
R16 B.n549 B.n70 585
R17 B.n551 B.n550 585
R18 B.n552 B.n69 585
R19 B.n554 B.n553 585
R20 B.n555 B.n68 585
R21 B.n557 B.n556 585
R22 B.n558 B.n67 585
R23 B.n560 B.n559 585
R24 B.n561 B.n66 585
R25 B.n563 B.n562 585
R26 B.n564 B.n65 585
R27 B.n566 B.n565 585
R28 B.n567 B.n64 585
R29 B.n569 B.n568 585
R30 B.n570 B.n63 585
R31 B.n572 B.n571 585
R32 B.n573 B.n62 585
R33 B.n575 B.n574 585
R34 B.n576 B.n61 585
R35 B.n578 B.n577 585
R36 B.n579 B.n60 585
R37 B.n581 B.n580 585
R38 B.n582 B.n59 585
R39 B.n584 B.n583 585
R40 B.n585 B.n58 585
R41 B.n587 B.n586 585
R42 B.n588 B.n57 585
R43 B.n590 B.n589 585
R44 B.n591 B.n56 585
R45 B.n593 B.n592 585
R46 B.n594 B.n55 585
R47 B.n596 B.n595 585
R48 B.n598 B.n597 585
R49 B.n599 B.n51 585
R50 B.n601 B.n600 585
R51 B.n602 B.n50 585
R52 B.n604 B.n603 585
R53 B.n605 B.n49 585
R54 B.n607 B.n606 585
R55 B.n608 B.n48 585
R56 B.n610 B.n609 585
R57 B.n611 B.n45 585
R58 B.n614 B.n613 585
R59 B.n615 B.n44 585
R60 B.n617 B.n616 585
R61 B.n618 B.n43 585
R62 B.n620 B.n619 585
R63 B.n621 B.n42 585
R64 B.n623 B.n622 585
R65 B.n624 B.n41 585
R66 B.n626 B.n625 585
R67 B.n627 B.n40 585
R68 B.n629 B.n628 585
R69 B.n630 B.n39 585
R70 B.n632 B.n631 585
R71 B.n633 B.n38 585
R72 B.n635 B.n634 585
R73 B.n636 B.n37 585
R74 B.n638 B.n637 585
R75 B.n639 B.n36 585
R76 B.n641 B.n640 585
R77 B.n642 B.n35 585
R78 B.n644 B.n643 585
R79 B.n645 B.n34 585
R80 B.n647 B.n646 585
R81 B.n648 B.n33 585
R82 B.n650 B.n649 585
R83 B.n651 B.n32 585
R84 B.n653 B.n652 585
R85 B.n654 B.n31 585
R86 B.n656 B.n655 585
R87 B.n657 B.n30 585
R88 B.n659 B.n658 585
R89 B.n660 B.n29 585
R90 B.n662 B.n661 585
R91 B.n663 B.n28 585
R92 B.n665 B.n664 585
R93 B.n666 B.n27 585
R94 B.n668 B.n667 585
R95 B.n669 B.n26 585
R96 B.n671 B.n670 585
R97 B.n672 B.n25 585
R98 B.n674 B.n673 585
R99 B.n675 B.n24 585
R100 B.n677 B.n676 585
R101 B.n678 B.n23 585
R102 B.n680 B.n679 585
R103 B.n681 B.n22 585
R104 B.n683 B.n682 585
R105 B.n684 B.n21 585
R106 B.n524 B.n523 585
R107 B.n522 B.n79 585
R108 B.n521 B.n520 585
R109 B.n519 B.n80 585
R110 B.n518 B.n517 585
R111 B.n516 B.n81 585
R112 B.n515 B.n514 585
R113 B.n513 B.n82 585
R114 B.n512 B.n511 585
R115 B.n510 B.n83 585
R116 B.n509 B.n508 585
R117 B.n507 B.n84 585
R118 B.n506 B.n505 585
R119 B.n504 B.n85 585
R120 B.n503 B.n502 585
R121 B.n501 B.n86 585
R122 B.n500 B.n499 585
R123 B.n498 B.n87 585
R124 B.n497 B.n496 585
R125 B.n495 B.n88 585
R126 B.n494 B.n493 585
R127 B.n492 B.n89 585
R128 B.n491 B.n490 585
R129 B.n489 B.n90 585
R130 B.n488 B.n487 585
R131 B.n486 B.n91 585
R132 B.n485 B.n484 585
R133 B.n483 B.n92 585
R134 B.n482 B.n481 585
R135 B.n480 B.n93 585
R136 B.n479 B.n478 585
R137 B.n477 B.n94 585
R138 B.n476 B.n475 585
R139 B.n474 B.n95 585
R140 B.n473 B.n472 585
R141 B.n471 B.n96 585
R142 B.n470 B.n469 585
R143 B.n468 B.n97 585
R144 B.n467 B.n466 585
R145 B.n465 B.n98 585
R146 B.n464 B.n463 585
R147 B.n462 B.n99 585
R148 B.n461 B.n460 585
R149 B.n459 B.n100 585
R150 B.n458 B.n457 585
R151 B.n456 B.n101 585
R152 B.n455 B.n454 585
R153 B.n453 B.n102 585
R154 B.n452 B.n451 585
R155 B.n450 B.n103 585
R156 B.n449 B.n448 585
R157 B.n447 B.n104 585
R158 B.n446 B.n445 585
R159 B.n444 B.n105 585
R160 B.n443 B.n442 585
R161 B.n441 B.n106 585
R162 B.n440 B.n439 585
R163 B.n438 B.n107 585
R164 B.n437 B.n436 585
R165 B.n435 B.n108 585
R166 B.n434 B.n433 585
R167 B.n432 B.n109 585
R168 B.n431 B.n430 585
R169 B.n429 B.n110 585
R170 B.n428 B.n427 585
R171 B.n426 B.n111 585
R172 B.n425 B.n424 585
R173 B.n423 B.n112 585
R174 B.n422 B.n421 585
R175 B.n420 B.n113 585
R176 B.n419 B.n418 585
R177 B.n417 B.n114 585
R178 B.n416 B.n415 585
R179 B.n414 B.n115 585
R180 B.n413 B.n412 585
R181 B.n411 B.n116 585
R182 B.n410 B.n409 585
R183 B.n249 B.n174 585
R184 B.n251 B.n250 585
R185 B.n252 B.n173 585
R186 B.n254 B.n253 585
R187 B.n255 B.n172 585
R188 B.n257 B.n256 585
R189 B.n258 B.n171 585
R190 B.n260 B.n259 585
R191 B.n261 B.n170 585
R192 B.n263 B.n262 585
R193 B.n264 B.n169 585
R194 B.n266 B.n265 585
R195 B.n267 B.n168 585
R196 B.n269 B.n268 585
R197 B.n270 B.n167 585
R198 B.n272 B.n271 585
R199 B.n273 B.n166 585
R200 B.n275 B.n274 585
R201 B.n276 B.n165 585
R202 B.n278 B.n277 585
R203 B.n279 B.n164 585
R204 B.n281 B.n280 585
R205 B.n282 B.n163 585
R206 B.n284 B.n283 585
R207 B.n285 B.n162 585
R208 B.n287 B.n286 585
R209 B.n288 B.n161 585
R210 B.n290 B.n289 585
R211 B.n291 B.n160 585
R212 B.n293 B.n292 585
R213 B.n294 B.n159 585
R214 B.n296 B.n295 585
R215 B.n297 B.n158 585
R216 B.n299 B.n298 585
R217 B.n300 B.n157 585
R218 B.n302 B.n301 585
R219 B.n303 B.n156 585
R220 B.n305 B.n304 585
R221 B.n306 B.n155 585
R222 B.n308 B.n307 585
R223 B.n309 B.n154 585
R224 B.n311 B.n310 585
R225 B.n312 B.n153 585
R226 B.n314 B.n313 585
R227 B.n315 B.n152 585
R228 B.n317 B.n316 585
R229 B.n318 B.n151 585
R230 B.n320 B.n319 585
R231 B.n322 B.n321 585
R232 B.n323 B.n147 585
R233 B.n325 B.n324 585
R234 B.n326 B.n146 585
R235 B.n328 B.n327 585
R236 B.n329 B.n145 585
R237 B.n331 B.n330 585
R238 B.n332 B.n144 585
R239 B.n334 B.n333 585
R240 B.n335 B.n141 585
R241 B.n338 B.n337 585
R242 B.n339 B.n140 585
R243 B.n341 B.n340 585
R244 B.n342 B.n139 585
R245 B.n344 B.n343 585
R246 B.n345 B.n138 585
R247 B.n347 B.n346 585
R248 B.n348 B.n137 585
R249 B.n350 B.n349 585
R250 B.n351 B.n136 585
R251 B.n353 B.n352 585
R252 B.n354 B.n135 585
R253 B.n356 B.n355 585
R254 B.n357 B.n134 585
R255 B.n359 B.n358 585
R256 B.n360 B.n133 585
R257 B.n362 B.n361 585
R258 B.n363 B.n132 585
R259 B.n365 B.n364 585
R260 B.n366 B.n131 585
R261 B.n368 B.n367 585
R262 B.n369 B.n130 585
R263 B.n371 B.n370 585
R264 B.n372 B.n129 585
R265 B.n374 B.n373 585
R266 B.n375 B.n128 585
R267 B.n377 B.n376 585
R268 B.n378 B.n127 585
R269 B.n380 B.n379 585
R270 B.n381 B.n126 585
R271 B.n383 B.n382 585
R272 B.n384 B.n125 585
R273 B.n386 B.n385 585
R274 B.n387 B.n124 585
R275 B.n389 B.n388 585
R276 B.n390 B.n123 585
R277 B.n392 B.n391 585
R278 B.n393 B.n122 585
R279 B.n395 B.n394 585
R280 B.n396 B.n121 585
R281 B.n398 B.n397 585
R282 B.n399 B.n120 585
R283 B.n401 B.n400 585
R284 B.n402 B.n119 585
R285 B.n404 B.n403 585
R286 B.n405 B.n118 585
R287 B.n407 B.n406 585
R288 B.n408 B.n117 585
R289 B.n248 B.n247 585
R290 B.n246 B.n175 585
R291 B.n245 B.n244 585
R292 B.n243 B.n176 585
R293 B.n242 B.n241 585
R294 B.n240 B.n177 585
R295 B.n239 B.n238 585
R296 B.n237 B.n178 585
R297 B.n236 B.n235 585
R298 B.n234 B.n179 585
R299 B.n233 B.n232 585
R300 B.n231 B.n180 585
R301 B.n230 B.n229 585
R302 B.n228 B.n181 585
R303 B.n227 B.n226 585
R304 B.n225 B.n182 585
R305 B.n224 B.n223 585
R306 B.n222 B.n183 585
R307 B.n221 B.n220 585
R308 B.n219 B.n184 585
R309 B.n218 B.n217 585
R310 B.n216 B.n185 585
R311 B.n215 B.n214 585
R312 B.n213 B.n186 585
R313 B.n212 B.n211 585
R314 B.n210 B.n187 585
R315 B.n209 B.n208 585
R316 B.n207 B.n188 585
R317 B.n206 B.n205 585
R318 B.n204 B.n189 585
R319 B.n203 B.n202 585
R320 B.n201 B.n190 585
R321 B.n200 B.n199 585
R322 B.n198 B.n191 585
R323 B.n197 B.n196 585
R324 B.n195 B.n192 585
R325 B.n194 B.n193 585
R326 B.n2 B.n0 585
R327 B.n741 B.n1 585
R328 B.n740 B.n739 585
R329 B.n738 B.n3 585
R330 B.n737 B.n736 585
R331 B.n735 B.n4 585
R332 B.n734 B.n733 585
R333 B.n732 B.n5 585
R334 B.n731 B.n730 585
R335 B.n729 B.n6 585
R336 B.n728 B.n727 585
R337 B.n726 B.n7 585
R338 B.n725 B.n724 585
R339 B.n723 B.n8 585
R340 B.n722 B.n721 585
R341 B.n720 B.n9 585
R342 B.n719 B.n718 585
R343 B.n717 B.n10 585
R344 B.n716 B.n715 585
R345 B.n714 B.n11 585
R346 B.n713 B.n712 585
R347 B.n711 B.n12 585
R348 B.n710 B.n709 585
R349 B.n708 B.n13 585
R350 B.n707 B.n706 585
R351 B.n705 B.n14 585
R352 B.n704 B.n703 585
R353 B.n702 B.n15 585
R354 B.n701 B.n700 585
R355 B.n699 B.n16 585
R356 B.n698 B.n697 585
R357 B.n696 B.n17 585
R358 B.n695 B.n694 585
R359 B.n693 B.n18 585
R360 B.n692 B.n691 585
R361 B.n690 B.n19 585
R362 B.n689 B.n688 585
R363 B.n687 B.n20 585
R364 B.n686 B.n685 585
R365 B.n743 B.n742 585
R366 B.n249 B.n248 506.916
R367 B.n686 B.n21 506.916
R368 B.n410 B.n117 506.916
R369 B.n525 B.n524 506.916
R370 B.n142 B.t5 455.327
R371 B.n52 B.t7 455.327
R372 B.n148 B.t2 455.327
R373 B.n46 B.t10 455.327
R374 B.n143 B.t4 415.764
R375 B.n53 B.t8 415.764
R376 B.n149 B.t1 415.764
R377 B.n47 B.t11 415.764
R378 B.n142 B.t3 406.555
R379 B.n148 B.t0 406.555
R380 B.n46 B.t9 406.555
R381 B.n52 B.t6 406.555
R382 B.n248 B.n175 163.367
R383 B.n244 B.n175 163.367
R384 B.n244 B.n243 163.367
R385 B.n243 B.n242 163.367
R386 B.n242 B.n177 163.367
R387 B.n238 B.n177 163.367
R388 B.n238 B.n237 163.367
R389 B.n237 B.n236 163.367
R390 B.n236 B.n179 163.367
R391 B.n232 B.n179 163.367
R392 B.n232 B.n231 163.367
R393 B.n231 B.n230 163.367
R394 B.n230 B.n181 163.367
R395 B.n226 B.n181 163.367
R396 B.n226 B.n225 163.367
R397 B.n225 B.n224 163.367
R398 B.n224 B.n183 163.367
R399 B.n220 B.n183 163.367
R400 B.n220 B.n219 163.367
R401 B.n219 B.n218 163.367
R402 B.n218 B.n185 163.367
R403 B.n214 B.n185 163.367
R404 B.n214 B.n213 163.367
R405 B.n213 B.n212 163.367
R406 B.n212 B.n187 163.367
R407 B.n208 B.n187 163.367
R408 B.n208 B.n207 163.367
R409 B.n207 B.n206 163.367
R410 B.n206 B.n189 163.367
R411 B.n202 B.n189 163.367
R412 B.n202 B.n201 163.367
R413 B.n201 B.n200 163.367
R414 B.n200 B.n191 163.367
R415 B.n196 B.n191 163.367
R416 B.n196 B.n195 163.367
R417 B.n195 B.n194 163.367
R418 B.n194 B.n2 163.367
R419 B.n742 B.n2 163.367
R420 B.n742 B.n741 163.367
R421 B.n741 B.n740 163.367
R422 B.n740 B.n3 163.367
R423 B.n736 B.n3 163.367
R424 B.n736 B.n735 163.367
R425 B.n735 B.n734 163.367
R426 B.n734 B.n5 163.367
R427 B.n730 B.n5 163.367
R428 B.n730 B.n729 163.367
R429 B.n729 B.n728 163.367
R430 B.n728 B.n7 163.367
R431 B.n724 B.n7 163.367
R432 B.n724 B.n723 163.367
R433 B.n723 B.n722 163.367
R434 B.n722 B.n9 163.367
R435 B.n718 B.n9 163.367
R436 B.n718 B.n717 163.367
R437 B.n717 B.n716 163.367
R438 B.n716 B.n11 163.367
R439 B.n712 B.n11 163.367
R440 B.n712 B.n711 163.367
R441 B.n711 B.n710 163.367
R442 B.n710 B.n13 163.367
R443 B.n706 B.n13 163.367
R444 B.n706 B.n705 163.367
R445 B.n705 B.n704 163.367
R446 B.n704 B.n15 163.367
R447 B.n700 B.n15 163.367
R448 B.n700 B.n699 163.367
R449 B.n699 B.n698 163.367
R450 B.n698 B.n17 163.367
R451 B.n694 B.n17 163.367
R452 B.n694 B.n693 163.367
R453 B.n693 B.n692 163.367
R454 B.n692 B.n19 163.367
R455 B.n688 B.n19 163.367
R456 B.n688 B.n687 163.367
R457 B.n687 B.n686 163.367
R458 B.n250 B.n249 163.367
R459 B.n250 B.n173 163.367
R460 B.n254 B.n173 163.367
R461 B.n255 B.n254 163.367
R462 B.n256 B.n255 163.367
R463 B.n256 B.n171 163.367
R464 B.n260 B.n171 163.367
R465 B.n261 B.n260 163.367
R466 B.n262 B.n261 163.367
R467 B.n262 B.n169 163.367
R468 B.n266 B.n169 163.367
R469 B.n267 B.n266 163.367
R470 B.n268 B.n267 163.367
R471 B.n268 B.n167 163.367
R472 B.n272 B.n167 163.367
R473 B.n273 B.n272 163.367
R474 B.n274 B.n273 163.367
R475 B.n274 B.n165 163.367
R476 B.n278 B.n165 163.367
R477 B.n279 B.n278 163.367
R478 B.n280 B.n279 163.367
R479 B.n280 B.n163 163.367
R480 B.n284 B.n163 163.367
R481 B.n285 B.n284 163.367
R482 B.n286 B.n285 163.367
R483 B.n286 B.n161 163.367
R484 B.n290 B.n161 163.367
R485 B.n291 B.n290 163.367
R486 B.n292 B.n291 163.367
R487 B.n292 B.n159 163.367
R488 B.n296 B.n159 163.367
R489 B.n297 B.n296 163.367
R490 B.n298 B.n297 163.367
R491 B.n298 B.n157 163.367
R492 B.n302 B.n157 163.367
R493 B.n303 B.n302 163.367
R494 B.n304 B.n303 163.367
R495 B.n304 B.n155 163.367
R496 B.n308 B.n155 163.367
R497 B.n309 B.n308 163.367
R498 B.n310 B.n309 163.367
R499 B.n310 B.n153 163.367
R500 B.n314 B.n153 163.367
R501 B.n315 B.n314 163.367
R502 B.n316 B.n315 163.367
R503 B.n316 B.n151 163.367
R504 B.n320 B.n151 163.367
R505 B.n321 B.n320 163.367
R506 B.n321 B.n147 163.367
R507 B.n325 B.n147 163.367
R508 B.n326 B.n325 163.367
R509 B.n327 B.n326 163.367
R510 B.n327 B.n145 163.367
R511 B.n331 B.n145 163.367
R512 B.n332 B.n331 163.367
R513 B.n333 B.n332 163.367
R514 B.n333 B.n141 163.367
R515 B.n338 B.n141 163.367
R516 B.n339 B.n338 163.367
R517 B.n340 B.n339 163.367
R518 B.n340 B.n139 163.367
R519 B.n344 B.n139 163.367
R520 B.n345 B.n344 163.367
R521 B.n346 B.n345 163.367
R522 B.n346 B.n137 163.367
R523 B.n350 B.n137 163.367
R524 B.n351 B.n350 163.367
R525 B.n352 B.n351 163.367
R526 B.n352 B.n135 163.367
R527 B.n356 B.n135 163.367
R528 B.n357 B.n356 163.367
R529 B.n358 B.n357 163.367
R530 B.n358 B.n133 163.367
R531 B.n362 B.n133 163.367
R532 B.n363 B.n362 163.367
R533 B.n364 B.n363 163.367
R534 B.n364 B.n131 163.367
R535 B.n368 B.n131 163.367
R536 B.n369 B.n368 163.367
R537 B.n370 B.n369 163.367
R538 B.n370 B.n129 163.367
R539 B.n374 B.n129 163.367
R540 B.n375 B.n374 163.367
R541 B.n376 B.n375 163.367
R542 B.n376 B.n127 163.367
R543 B.n380 B.n127 163.367
R544 B.n381 B.n380 163.367
R545 B.n382 B.n381 163.367
R546 B.n382 B.n125 163.367
R547 B.n386 B.n125 163.367
R548 B.n387 B.n386 163.367
R549 B.n388 B.n387 163.367
R550 B.n388 B.n123 163.367
R551 B.n392 B.n123 163.367
R552 B.n393 B.n392 163.367
R553 B.n394 B.n393 163.367
R554 B.n394 B.n121 163.367
R555 B.n398 B.n121 163.367
R556 B.n399 B.n398 163.367
R557 B.n400 B.n399 163.367
R558 B.n400 B.n119 163.367
R559 B.n404 B.n119 163.367
R560 B.n405 B.n404 163.367
R561 B.n406 B.n405 163.367
R562 B.n406 B.n117 163.367
R563 B.n411 B.n410 163.367
R564 B.n412 B.n411 163.367
R565 B.n412 B.n115 163.367
R566 B.n416 B.n115 163.367
R567 B.n417 B.n416 163.367
R568 B.n418 B.n417 163.367
R569 B.n418 B.n113 163.367
R570 B.n422 B.n113 163.367
R571 B.n423 B.n422 163.367
R572 B.n424 B.n423 163.367
R573 B.n424 B.n111 163.367
R574 B.n428 B.n111 163.367
R575 B.n429 B.n428 163.367
R576 B.n430 B.n429 163.367
R577 B.n430 B.n109 163.367
R578 B.n434 B.n109 163.367
R579 B.n435 B.n434 163.367
R580 B.n436 B.n435 163.367
R581 B.n436 B.n107 163.367
R582 B.n440 B.n107 163.367
R583 B.n441 B.n440 163.367
R584 B.n442 B.n441 163.367
R585 B.n442 B.n105 163.367
R586 B.n446 B.n105 163.367
R587 B.n447 B.n446 163.367
R588 B.n448 B.n447 163.367
R589 B.n448 B.n103 163.367
R590 B.n452 B.n103 163.367
R591 B.n453 B.n452 163.367
R592 B.n454 B.n453 163.367
R593 B.n454 B.n101 163.367
R594 B.n458 B.n101 163.367
R595 B.n459 B.n458 163.367
R596 B.n460 B.n459 163.367
R597 B.n460 B.n99 163.367
R598 B.n464 B.n99 163.367
R599 B.n465 B.n464 163.367
R600 B.n466 B.n465 163.367
R601 B.n466 B.n97 163.367
R602 B.n470 B.n97 163.367
R603 B.n471 B.n470 163.367
R604 B.n472 B.n471 163.367
R605 B.n472 B.n95 163.367
R606 B.n476 B.n95 163.367
R607 B.n477 B.n476 163.367
R608 B.n478 B.n477 163.367
R609 B.n478 B.n93 163.367
R610 B.n482 B.n93 163.367
R611 B.n483 B.n482 163.367
R612 B.n484 B.n483 163.367
R613 B.n484 B.n91 163.367
R614 B.n488 B.n91 163.367
R615 B.n489 B.n488 163.367
R616 B.n490 B.n489 163.367
R617 B.n490 B.n89 163.367
R618 B.n494 B.n89 163.367
R619 B.n495 B.n494 163.367
R620 B.n496 B.n495 163.367
R621 B.n496 B.n87 163.367
R622 B.n500 B.n87 163.367
R623 B.n501 B.n500 163.367
R624 B.n502 B.n501 163.367
R625 B.n502 B.n85 163.367
R626 B.n506 B.n85 163.367
R627 B.n507 B.n506 163.367
R628 B.n508 B.n507 163.367
R629 B.n508 B.n83 163.367
R630 B.n512 B.n83 163.367
R631 B.n513 B.n512 163.367
R632 B.n514 B.n513 163.367
R633 B.n514 B.n81 163.367
R634 B.n518 B.n81 163.367
R635 B.n519 B.n518 163.367
R636 B.n520 B.n519 163.367
R637 B.n520 B.n79 163.367
R638 B.n524 B.n79 163.367
R639 B.n682 B.n21 163.367
R640 B.n682 B.n681 163.367
R641 B.n681 B.n680 163.367
R642 B.n680 B.n23 163.367
R643 B.n676 B.n23 163.367
R644 B.n676 B.n675 163.367
R645 B.n675 B.n674 163.367
R646 B.n674 B.n25 163.367
R647 B.n670 B.n25 163.367
R648 B.n670 B.n669 163.367
R649 B.n669 B.n668 163.367
R650 B.n668 B.n27 163.367
R651 B.n664 B.n27 163.367
R652 B.n664 B.n663 163.367
R653 B.n663 B.n662 163.367
R654 B.n662 B.n29 163.367
R655 B.n658 B.n29 163.367
R656 B.n658 B.n657 163.367
R657 B.n657 B.n656 163.367
R658 B.n656 B.n31 163.367
R659 B.n652 B.n31 163.367
R660 B.n652 B.n651 163.367
R661 B.n651 B.n650 163.367
R662 B.n650 B.n33 163.367
R663 B.n646 B.n33 163.367
R664 B.n646 B.n645 163.367
R665 B.n645 B.n644 163.367
R666 B.n644 B.n35 163.367
R667 B.n640 B.n35 163.367
R668 B.n640 B.n639 163.367
R669 B.n639 B.n638 163.367
R670 B.n638 B.n37 163.367
R671 B.n634 B.n37 163.367
R672 B.n634 B.n633 163.367
R673 B.n633 B.n632 163.367
R674 B.n632 B.n39 163.367
R675 B.n628 B.n39 163.367
R676 B.n628 B.n627 163.367
R677 B.n627 B.n626 163.367
R678 B.n626 B.n41 163.367
R679 B.n622 B.n41 163.367
R680 B.n622 B.n621 163.367
R681 B.n621 B.n620 163.367
R682 B.n620 B.n43 163.367
R683 B.n616 B.n43 163.367
R684 B.n616 B.n615 163.367
R685 B.n615 B.n614 163.367
R686 B.n614 B.n45 163.367
R687 B.n609 B.n45 163.367
R688 B.n609 B.n608 163.367
R689 B.n608 B.n607 163.367
R690 B.n607 B.n49 163.367
R691 B.n603 B.n49 163.367
R692 B.n603 B.n602 163.367
R693 B.n602 B.n601 163.367
R694 B.n601 B.n51 163.367
R695 B.n597 B.n51 163.367
R696 B.n597 B.n596 163.367
R697 B.n596 B.n55 163.367
R698 B.n592 B.n55 163.367
R699 B.n592 B.n591 163.367
R700 B.n591 B.n590 163.367
R701 B.n590 B.n57 163.367
R702 B.n586 B.n57 163.367
R703 B.n586 B.n585 163.367
R704 B.n585 B.n584 163.367
R705 B.n584 B.n59 163.367
R706 B.n580 B.n59 163.367
R707 B.n580 B.n579 163.367
R708 B.n579 B.n578 163.367
R709 B.n578 B.n61 163.367
R710 B.n574 B.n61 163.367
R711 B.n574 B.n573 163.367
R712 B.n573 B.n572 163.367
R713 B.n572 B.n63 163.367
R714 B.n568 B.n63 163.367
R715 B.n568 B.n567 163.367
R716 B.n567 B.n566 163.367
R717 B.n566 B.n65 163.367
R718 B.n562 B.n65 163.367
R719 B.n562 B.n561 163.367
R720 B.n561 B.n560 163.367
R721 B.n560 B.n67 163.367
R722 B.n556 B.n67 163.367
R723 B.n556 B.n555 163.367
R724 B.n555 B.n554 163.367
R725 B.n554 B.n69 163.367
R726 B.n550 B.n69 163.367
R727 B.n550 B.n549 163.367
R728 B.n549 B.n548 163.367
R729 B.n548 B.n71 163.367
R730 B.n544 B.n71 163.367
R731 B.n544 B.n543 163.367
R732 B.n543 B.n542 163.367
R733 B.n542 B.n73 163.367
R734 B.n538 B.n73 163.367
R735 B.n538 B.n537 163.367
R736 B.n537 B.n536 163.367
R737 B.n536 B.n75 163.367
R738 B.n532 B.n75 163.367
R739 B.n532 B.n531 163.367
R740 B.n531 B.n530 163.367
R741 B.n530 B.n77 163.367
R742 B.n526 B.n77 163.367
R743 B.n526 B.n525 163.367
R744 B.n336 B.n143 59.5399
R745 B.n150 B.n149 59.5399
R746 B.n612 B.n47 59.5399
R747 B.n54 B.n53 59.5399
R748 B.n143 B.n142 39.5641
R749 B.n149 B.n148 39.5641
R750 B.n47 B.n46 39.5641
R751 B.n53 B.n52 39.5641
R752 B.n685 B.n684 32.9371
R753 B.n523 B.n78 32.9371
R754 B.n409 B.n408 32.9371
R755 B.n247 B.n174 32.9371
R756 B B.n743 18.0485
R757 B.n684 B.n683 10.6151
R758 B.n683 B.n22 10.6151
R759 B.n679 B.n22 10.6151
R760 B.n679 B.n678 10.6151
R761 B.n678 B.n677 10.6151
R762 B.n677 B.n24 10.6151
R763 B.n673 B.n24 10.6151
R764 B.n673 B.n672 10.6151
R765 B.n672 B.n671 10.6151
R766 B.n671 B.n26 10.6151
R767 B.n667 B.n26 10.6151
R768 B.n667 B.n666 10.6151
R769 B.n666 B.n665 10.6151
R770 B.n665 B.n28 10.6151
R771 B.n661 B.n28 10.6151
R772 B.n661 B.n660 10.6151
R773 B.n660 B.n659 10.6151
R774 B.n659 B.n30 10.6151
R775 B.n655 B.n30 10.6151
R776 B.n655 B.n654 10.6151
R777 B.n654 B.n653 10.6151
R778 B.n653 B.n32 10.6151
R779 B.n649 B.n32 10.6151
R780 B.n649 B.n648 10.6151
R781 B.n648 B.n647 10.6151
R782 B.n647 B.n34 10.6151
R783 B.n643 B.n34 10.6151
R784 B.n643 B.n642 10.6151
R785 B.n642 B.n641 10.6151
R786 B.n641 B.n36 10.6151
R787 B.n637 B.n36 10.6151
R788 B.n637 B.n636 10.6151
R789 B.n636 B.n635 10.6151
R790 B.n635 B.n38 10.6151
R791 B.n631 B.n38 10.6151
R792 B.n631 B.n630 10.6151
R793 B.n630 B.n629 10.6151
R794 B.n629 B.n40 10.6151
R795 B.n625 B.n40 10.6151
R796 B.n625 B.n624 10.6151
R797 B.n624 B.n623 10.6151
R798 B.n623 B.n42 10.6151
R799 B.n619 B.n42 10.6151
R800 B.n619 B.n618 10.6151
R801 B.n618 B.n617 10.6151
R802 B.n617 B.n44 10.6151
R803 B.n613 B.n44 10.6151
R804 B.n611 B.n610 10.6151
R805 B.n610 B.n48 10.6151
R806 B.n606 B.n48 10.6151
R807 B.n606 B.n605 10.6151
R808 B.n605 B.n604 10.6151
R809 B.n604 B.n50 10.6151
R810 B.n600 B.n50 10.6151
R811 B.n600 B.n599 10.6151
R812 B.n599 B.n598 10.6151
R813 B.n595 B.n594 10.6151
R814 B.n594 B.n593 10.6151
R815 B.n593 B.n56 10.6151
R816 B.n589 B.n56 10.6151
R817 B.n589 B.n588 10.6151
R818 B.n588 B.n587 10.6151
R819 B.n587 B.n58 10.6151
R820 B.n583 B.n58 10.6151
R821 B.n583 B.n582 10.6151
R822 B.n582 B.n581 10.6151
R823 B.n581 B.n60 10.6151
R824 B.n577 B.n60 10.6151
R825 B.n577 B.n576 10.6151
R826 B.n576 B.n575 10.6151
R827 B.n575 B.n62 10.6151
R828 B.n571 B.n62 10.6151
R829 B.n571 B.n570 10.6151
R830 B.n570 B.n569 10.6151
R831 B.n569 B.n64 10.6151
R832 B.n565 B.n64 10.6151
R833 B.n565 B.n564 10.6151
R834 B.n564 B.n563 10.6151
R835 B.n563 B.n66 10.6151
R836 B.n559 B.n66 10.6151
R837 B.n559 B.n558 10.6151
R838 B.n558 B.n557 10.6151
R839 B.n557 B.n68 10.6151
R840 B.n553 B.n68 10.6151
R841 B.n553 B.n552 10.6151
R842 B.n552 B.n551 10.6151
R843 B.n551 B.n70 10.6151
R844 B.n547 B.n70 10.6151
R845 B.n547 B.n546 10.6151
R846 B.n546 B.n545 10.6151
R847 B.n545 B.n72 10.6151
R848 B.n541 B.n72 10.6151
R849 B.n541 B.n540 10.6151
R850 B.n540 B.n539 10.6151
R851 B.n539 B.n74 10.6151
R852 B.n535 B.n74 10.6151
R853 B.n535 B.n534 10.6151
R854 B.n534 B.n533 10.6151
R855 B.n533 B.n76 10.6151
R856 B.n529 B.n76 10.6151
R857 B.n529 B.n528 10.6151
R858 B.n528 B.n527 10.6151
R859 B.n527 B.n78 10.6151
R860 B.n409 B.n116 10.6151
R861 B.n413 B.n116 10.6151
R862 B.n414 B.n413 10.6151
R863 B.n415 B.n414 10.6151
R864 B.n415 B.n114 10.6151
R865 B.n419 B.n114 10.6151
R866 B.n420 B.n419 10.6151
R867 B.n421 B.n420 10.6151
R868 B.n421 B.n112 10.6151
R869 B.n425 B.n112 10.6151
R870 B.n426 B.n425 10.6151
R871 B.n427 B.n426 10.6151
R872 B.n427 B.n110 10.6151
R873 B.n431 B.n110 10.6151
R874 B.n432 B.n431 10.6151
R875 B.n433 B.n432 10.6151
R876 B.n433 B.n108 10.6151
R877 B.n437 B.n108 10.6151
R878 B.n438 B.n437 10.6151
R879 B.n439 B.n438 10.6151
R880 B.n439 B.n106 10.6151
R881 B.n443 B.n106 10.6151
R882 B.n444 B.n443 10.6151
R883 B.n445 B.n444 10.6151
R884 B.n445 B.n104 10.6151
R885 B.n449 B.n104 10.6151
R886 B.n450 B.n449 10.6151
R887 B.n451 B.n450 10.6151
R888 B.n451 B.n102 10.6151
R889 B.n455 B.n102 10.6151
R890 B.n456 B.n455 10.6151
R891 B.n457 B.n456 10.6151
R892 B.n457 B.n100 10.6151
R893 B.n461 B.n100 10.6151
R894 B.n462 B.n461 10.6151
R895 B.n463 B.n462 10.6151
R896 B.n463 B.n98 10.6151
R897 B.n467 B.n98 10.6151
R898 B.n468 B.n467 10.6151
R899 B.n469 B.n468 10.6151
R900 B.n469 B.n96 10.6151
R901 B.n473 B.n96 10.6151
R902 B.n474 B.n473 10.6151
R903 B.n475 B.n474 10.6151
R904 B.n475 B.n94 10.6151
R905 B.n479 B.n94 10.6151
R906 B.n480 B.n479 10.6151
R907 B.n481 B.n480 10.6151
R908 B.n481 B.n92 10.6151
R909 B.n485 B.n92 10.6151
R910 B.n486 B.n485 10.6151
R911 B.n487 B.n486 10.6151
R912 B.n487 B.n90 10.6151
R913 B.n491 B.n90 10.6151
R914 B.n492 B.n491 10.6151
R915 B.n493 B.n492 10.6151
R916 B.n493 B.n88 10.6151
R917 B.n497 B.n88 10.6151
R918 B.n498 B.n497 10.6151
R919 B.n499 B.n498 10.6151
R920 B.n499 B.n86 10.6151
R921 B.n503 B.n86 10.6151
R922 B.n504 B.n503 10.6151
R923 B.n505 B.n504 10.6151
R924 B.n505 B.n84 10.6151
R925 B.n509 B.n84 10.6151
R926 B.n510 B.n509 10.6151
R927 B.n511 B.n510 10.6151
R928 B.n511 B.n82 10.6151
R929 B.n515 B.n82 10.6151
R930 B.n516 B.n515 10.6151
R931 B.n517 B.n516 10.6151
R932 B.n517 B.n80 10.6151
R933 B.n521 B.n80 10.6151
R934 B.n522 B.n521 10.6151
R935 B.n523 B.n522 10.6151
R936 B.n251 B.n174 10.6151
R937 B.n252 B.n251 10.6151
R938 B.n253 B.n252 10.6151
R939 B.n253 B.n172 10.6151
R940 B.n257 B.n172 10.6151
R941 B.n258 B.n257 10.6151
R942 B.n259 B.n258 10.6151
R943 B.n259 B.n170 10.6151
R944 B.n263 B.n170 10.6151
R945 B.n264 B.n263 10.6151
R946 B.n265 B.n264 10.6151
R947 B.n265 B.n168 10.6151
R948 B.n269 B.n168 10.6151
R949 B.n270 B.n269 10.6151
R950 B.n271 B.n270 10.6151
R951 B.n271 B.n166 10.6151
R952 B.n275 B.n166 10.6151
R953 B.n276 B.n275 10.6151
R954 B.n277 B.n276 10.6151
R955 B.n277 B.n164 10.6151
R956 B.n281 B.n164 10.6151
R957 B.n282 B.n281 10.6151
R958 B.n283 B.n282 10.6151
R959 B.n283 B.n162 10.6151
R960 B.n287 B.n162 10.6151
R961 B.n288 B.n287 10.6151
R962 B.n289 B.n288 10.6151
R963 B.n289 B.n160 10.6151
R964 B.n293 B.n160 10.6151
R965 B.n294 B.n293 10.6151
R966 B.n295 B.n294 10.6151
R967 B.n295 B.n158 10.6151
R968 B.n299 B.n158 10.6151
R969 B.n300 B.n299 10.6151
R970 B.n301 B.n300 10.6151
R971 B.n301 B.n156 10.6151
R972 B.n305 B.n156 10.6151
R973 B.n306 B.n305 10.6151
R974 B.n307 B.n306 10.6151
R975 B.n307 B.n154 10.6151
R976 B.n311 B.n154 10.6151
R977 B.n312 B.n311 10.6151
R978 B.n313 B.n312 10.6151
R979 B.n313 B.n152 10.6151
R980 B.n317 B.n152 10.6151
R981 B.n318 B.n317 10.6151
R982 B.n319 B.n318 10.6151
R983 B.n323 B.n322 10.6151
R984 B.n324 B.n323 10.6151
R985 B.n324 B.n146 10.6151
R986 B.n328 B.n146 10.6151
R987 B.n329 B.n328 10.6151
R988 B.n330 B.n329 10.6151
R989 B.n330 B.n144 10.6151
R990 B.n334 B.n144 10.6151
R991 B.n335 B.n334 10.6151
R992 B.n337 B.n140 10.6151
R993 B.n341 B.n140 10.6151
R994 B.n342 B.n341 10.6151
R995 B.n343 B.n342 10.6151
R996 B.n343 B.n138 10.6151
R997 B.n347 B.n138 10.6151
R998 B.n348 B.n347 10.6151
R999 B.n349 B.n348 10.6151
R1000 B.n349 B.n136 10.6151
R1001 B.n353 B.n136 10.6151
R1002 B.n354 B.n353 10.6151
R1003 B.n355 B.n354 10.6151
R1004 B.n355 B.n134 10.6151
R1005 B.n359 B.n134 10.6151
R1006 B.n360 B.n359 10.6151
R1007 B.n361 B.n360 10.6151
R1008 B.n361 B.n132 10.6151
R1009 B.n365 B.n132 10.6151
R1010 B.n366 B.n365 10.6151
R1011 B.n367 B.n366 10.6151
R1012 B.n367 B.n130 10.6151
R1013 B.n371 B.n130 10.6151
R1014 B.n372 B.n371 10.6151
R1015 B.n373 B.n372 10.6151
R1016 B.n373 B.n128 10.6151
R1017 B.n377 B.n128 10.6151
R1018 B.n378 B.n377 10.6151
R1019 B.n379 B.n378 10.6151
R1020 B.n379 B.n126 10.6151
R1021 B.n383 B.n126 10.6151
R1022 B.n384 B.n383 10.6151
R1023 B.n385 B.n384 10.6151
R1024 B.n385 B.n124 10.6151
R1025 B.n389 B.n124 10.6151
R1026 B.n390 B.n389 10.6151
R1027 B.n391 B.n390 10.6151
R1028 B.n391 B.n122 10.6151
R1029 B.n395 B.n122 10.6151
R1030 B.n396 B.n395 10.6151
R1031 B.n397 B.n396 10.6151
R1032 B.n397 B.n120 10.6151
R1033 B.n401 B.n120 10.6151
R1034 B.n402 B.n401 10.6151
R1035 B.n403 B.n402 10.6151
R1036 B.n403 B.n118 10.6151
R1037 B.n407 B.n118 10.6151
R1038 B.n408 B.n407 10.6151
R1039 B.n247 B.n246 10.6151
R1040 B.n246 B.n245 10.6151
R1041 B.n245 B.n176 10.6151
R1042 B.n241 B.n176 10.6151
R1043 B.n241 B.n240 10.6151
R1044 B.n240 B.n239 10.6151
R1045 B.n239 B.n178 10.6151
R1046 B.n235 B.n178 10.6151
R1047 B.n235 B.n234 10.6151
R1048 B.n234 B.n233 10.6151
R1049 B.n233 B.n180 10.6151
R1050 B.n229 B.n180 10.6151
R1051 B.n229 B.n228 10.6151
R1052 B.n228 B.n227 10.6151
R1053 B.n227 B.n182 10.6151
R1054 B.n223 B.n182 10.6151
R1055 B.n223 B.n222 10.6151
R1056 B.n222 B.n221 10.6151
R1057 B.n221 B.n184 10.6151
R1058 B.n217 B.n184 10.6151
R1059 B.n217 B.n216 10.6151
R1060 B.n216 B.n215 10.6151
R1061 B.n215 B.n186 10.6151
R1062 B.n211 B.n186 10.6151
R1063 B.n211 B.n210 10.6151
R1064 B.n210 B.n209 10.6151
R1065 B.n209 B.n188 10.6151
R1066 B.n205 B.n188 10.6151
R1067 B.n205 B.n204 10.6151
R1068 B.n204 B.n203 10.6151
R1069 B.n203 B.n190 10.6151
R1070 B.n199 B.n190 10.6151
R1071 B.n199 B.n198 10.6151
R1072 B.n198 B.n197 10.6151
R1073 B.n197 B.n192 10.6151
R1074 B.n193 B.n192 10.6151
R1075 B.n193 B.n0 10.6151
R1076 B.n739 B.n1 10.6151
R1077 B.n739 B.n738 10.6151
R1078 B.n738 B.n737 10.6151
R1079 B.n737 B.n4 10.6151
R1080 B.n733 B.n4 10.6151
R1081 B.n733 B.n732 10.6151
R1082 B.n732 B.n731 10.6151
R1083 B.n731 B.n6 10.6151
R1084 B.n727 B.n6 10.6151
R1085 B.n727 B.n726 10.6151
R1086 B.n726 B.n725 10.6151
R1087 B.n725 B.n8 10.6151
R1088 B.n721 B.n8 10.6151
R1089 B.n721 B.n720 10.6151
R1090 B.n720 B.n719 10.6151
R1091 B.n719 B.n10 10.6151
R1092 B.n715 B.n10 10.6151
R1093 B.n715 B.n714 10.6151
R1094 B.n714 B.n713 10.6151
R1095 B.n713 B.n12 10.6151
R1096 B.n709 B.n12 10.6151
R1097 B.n709 B.n708 10.6151
R1098 B.n708 B.n707 10.6151
R1099 B.n707 B.n14 10.6151
R1100 B.n703 B.n14 10.6151
R1101 B.n703 B.n702 10.6151
R1102 B.n702 B.n701 10.6151
R1103 B.n701 B.n16 10.6151
R1104 B.n697 B.n16 10.6151
R1105 B.n697 B.n696 10.6151
R1106 B.n696 B.n695 10.6151
R1107 B.n695 B.n18 10.6151
R1108 B.n691 B.n18 10.6151
R1109 B.n691 B.n690 10.6151
R1110 B.n690 B.n689 10.6151
R1111 B.n689 B.n20 10.6151
R1112 B.n685 B.n20 10.6151
R1113 B.n613 B.n612 9.36635
R1114 B.n595 B.n54 9.36635
R1115 B.n319 B.n150 9.36635
R1116 B.n337 B.n336 9.36635
R1117 B.n743 B.n0 2.81026
R1118 B.n743 B.n1 2.81026
R1119 B.n612 B.n611 1.24928
R1120 B.n598 B.n54 1.24928
R1121 B.n322 B.n150 1.24928
R1122 B.n336 B.n335 1.24928
R1123 VP.n12 VP.t5 229.371
R1124 VP.n31 VP.t4 200.411
R1125 VP.n38 VP.t6 200.411
R1126 VP.n46 VP.t3 200.411
R1127 VP.n53 VP.t2 200.411
R1128 VP.n28 VP.t1 200.411
R1129 VP.n21 VP.t0 200.411
R1130 VP.n13 VP.t7 200.411
R1131 VP.n31 VP.n30 182.722
R1132 VP.n54 VP.n53 182.722
R1133 VP.n29 VP.n28 182.722
R1134 VP.n14 VP.n11 161.3
R1135 VP.n16 VP.n15 161.3
R1136 VP.n17 VP.n10 161.3
R1137 VP.n19 VP.n18 161.3
R1138 VP.n20 VP.n9 161.3
R1139 VP.n23 VP.n22 161.3
R1140 VP.n24 VP.n8 161.3
R1141 VP.n26 VP.n25 161.3
R1142 VP.n27 VP.n7 161.3
R1143 VP.n52 VP.n0 161.3
R1144 VP.n51 VP.n50 161.3
R1145 VP.n49 VP.n1 161.3
R1146 VP.n48 VP.n47 161.3
R1147 VP.n45 VP.n2 161.3
R1148 VP.n44 VP.n43 161.3
R1149 VP.n42 VP.n3 161.3
R1150 VP.n41 VP.n40 161.3
R1151 VP.n39 VP.n4 161.3
R1152 VP.n37 VP.n36 161.3
R1153 VP.n35 VP.n5 161.3
R1154 VP.n34 VP.n33 161.3
R1155 VP.n32 VP.n6 161.3
R1156 VP.n13 VP.n12 67.3788
R1157 VP.n30 VP.n29 48.2808
R1158 VP.n33 VP.n5 44.3055
R1159 VP.n51 VP.n1 44.3055
R1160 VP.n26 VP.n8 44.3055
R1161 VP.n40 VP.n3 40.4106
R1162 VP.n44 VP.n3 40.4106
R1163 VP.n19 VP.n10 40.4106
R1164 VP.n15 VP.n10 40.4106
R1165 VP.n37 VP.n5 36.5157
R1166 VP.n47 VP.n1 36.5157
R1167 VP.n22 VP.n8 36.5157
R1168 VP.n33 VP.n32 24.3439
R1169 VP.n40 VP.n39 24.3439
R1170 VP.n45 VP.n44 24.3439
R1171 VP.n52 VP.n51 24.3439
R1172 VP.n27 VP.n26 24.3439
R1173 VP.n20 VP.n19 24.3439
R1174 VP.n15 VP.n14 24.3439
R1175 VP.n38 VP.n37 23.3702
R1176 VP.n47 VP.n46 23.3702
R1177 VP.n22 VP.n21 23.3702
R1178 VP.n12 VP.n11 18.7354
R1179 VP.n32 VP.n31 2.92171
R1180 VP.n53 VP.n52 2.92171
R1181 VP.n28 VP.n27 2.92171
R1182 VP.n39 VP.n38 0.974237
R1183 VP.n46 VP.n45 0.974237
R1184 VP.n21 VP.n20 0.974237
R1185 VP.n14 VP.n13 0.974237
R1186 VP.n16 VP.n11 0.189894
R1187 VP.n17 VP.n16 0.189894
R1188 VP.n18 VP.n17 0.189894
R1189 VP.n18 VP.n9 0.189894
R1190 VP.n23 VP.n9 0.189894
R1191 VP.n24 VP.n23 0.189894
R1192 VP.n25 VP.n24 0.189894
R1193 VP.n25 VP.n7 0.189894
R1194 VP.n29 VP.n7 0.189894
R1195 VP.n30 VP.n6 0.189894
R1196 VP.n34 VP.n6 0.189894
R1197 VP.n35 VP.n34 0.189894
R1198 VP.n36 VP.n35 0.189894
R1199 VP.n36 VP.n4 0.189894
R1200 VP.n41 VP.n4 0.189894
R1201 VP.n42 VP.n41 0.189894
R1202 VP.n43 VP.n42 0.189894
R1203 VP.n43 VP.n2 0.189894
R1204 VP.n48 VP.n2 0.189894
R1205 VP.n49 VP.n48 0.189894
R1206 VP.n50 VP.n49 0.189894
R1207 VP.n50 VP.n0 0.189894
R1208 VP.n54 VP.n0 0.189894
R1209 VP VP.n54 0.0516364
R1210 VDD1 VDD1.n0 71.4068
R1211 VDD1.n3 VDD1.n2 71.2933
R1212 VDD1.n3 VDD1.n1 71.2933
R1213 VDD1.n5 VDD1.n4 70.4693
R1214 VDD1.n5 VDD1.n3 44.4707
R1215 VDD1.n4 VDD1.t2 2.28637
R1216 VDD1.n4 VDD1.t3 2.28637
R1217 VDD1.n0 VDD1.t7 2.28637
R1218 VDD1.n0 VDD1.t5 2.28637
R1219 VDD1.n2 VDD1.t0 2.28637
R1220 VDD1.n2 VDD1.t6 2.28637
R1221 VDD1.n1 VDD1.t1 2.28637
R1222 VDD1.n1 VDD1.t4 2.28637
R1223 VDD1 VDD1.n5 0.821621
R1224 VTAIL.n626 VTAIL.n554 756.745
R1225 VTAIL.n74 VTAIL.n2 756.745
R1226 VTAIL.n152 VTAIL.n80 756.745
R1227 VTAIL.n232 VTAIL.n160 756.745
R1228 VTAIL.n548 VTAIL.n476 756.745
R1229 VTAIL.n468 VTAIL.n396 756.745
R1230 VTAIL.n390 VTAIL.n318 756.745
R1231 VTAIL.n310 VTAIL.n238 756.745
R1232 VTAIL.n578 VTAIL.n577 585
R1233 VTAIL.n583 VTAIL.n582 585
R1234 VTAIL.n585 VTAIL.n584 585
R1235 VTAIL.n574 VTAIL.n573 585
R1236 VTAIL.n591 VTAIL.n590 585
R1237 VTAIL.n593 VTAIL.n592 585
R1238 VTAIL.n570 VTAIL.n569 585
R1239 VTAIL.n600 VTAIL.n599 585
R1240 VTAIL.n601 VTAIL.n568 585
R1241 VTAIL.n603 VTAIL.n602 585
R1242 VTAIL.n566 VTAIL.n565 585
R1243 VTAIL.n609 VTAIL.n608 585
R1244 VTAIL.n611 VTAIL.n610 585
R1245 VTAIL.n562 VTAIL.n561 585
R1246 VTAIL.n617 VTAIL.n616 585
R1247 VTAIL.n619 VTAIL.n618 585
R1248 VTAIL.n558 VTAIL.n557 585
R1249 VTAIL.n625 VTAIL.n624 585
R1250 VTAIL.n627 VTAIL.n626 585
R1251 VTAIL.n26 VTAIL.n25 585
R1252 VTAIL.n31 VTAIL.n30 585
R1253 VTAIL.n33 VTAIL.n32 585
R1254 VTAIL.n22 VTAIL.n21 585
R1255 VTAIL.n39 VTAIL.n38 585
R1256 VTAIL.n41 VTAIL.n40 585
R1257 VTAIL.n18 VTAIL.n17 585
R1258 VTAIL.n48 VTAIL.n47 585
R1259 VTAIL.n49 VTAIL.n16 585
R1260 VTAIL.n51 VTAIL.n50 585
R1261 VTAIL.n14 VTAIL.n13 585
R1262 VTAIL.n57 VTAIL.n56 585
R1263 VTAIL.n59 VTAIL.n58 585
R1264 VTAIL.n10 VTAIL.n9 585
R1265 VTAIL.n65 VTAIL.n64 585
R1266 VTAIL.n67 VTAIL.n66 585
R1267 VTAIL.n6 VTAIL.n5 585
R1268 VTAIL.n73 VTAIL.n72 585
R1269 VTAIL.n75 VTAIL.n74 585
R1270 VTAIL.n104 VTAIL.n103 585
R1271 VTAIL.n109 VTAIL.n108 585
R1272 VTAIL.n111 VTAIL.n110 585
R1273 VTAIL.n100 VTAIL.n99 585
R1274 VTAIL.n117 VTAIL.n116 585
R1275 VTAIL.n119 VTAIL.n118 585
R1276 VTAIL.n96 VTAIL.n95 585
R1277 VTAIL.n126 VTAIL.n125 585
R1278 VTAIL.n127 VTAIL.n94 585
R1279 VTAIL.n129 VTAIL.n128 585
R1280 VTAIL.n92 VTAIL.n91 585
R1281 VTAIL.n135 VTAIL.n134 585
R1282 VTAIL.n137 VTAIL.n136 585
R1283 VTAIL.n88 VTAIL.n87 585
R1284 VTAIL.n143 VTAIL.n142 585
R1285 VTAIL.n145 VTAIL.n144 585
R1286 VTAIL.n84 VTAIL.n83 585
R1287 VTAIL.n151 VTAIL.n150 585
R1288 VTAIL.n153 VTAIL.n152 585
R1289 VTAIL.n184 VTAIL.n183 585
R1290 VTAIL.n189 VTAIL.n188 585
R1291 VTAIL.n191 VTAIL.n190 585
R1292 VTAIL.n180 VTAIL.n179 585
R1293 VTAIL.n197 VTAIL.n196 585
R1294 VTAIL.n199 VTAIL.n198 585
R1295 VTAIL.n176 VTAIL.n175 585
R1296 VTAIL.n206 VTAIL.n205 585
R1297 VTAIL.n207 VTAIL.n174 585
R1298 VTAIL.n209 VTAIL.n208 585
R1299 VTAIL.n172 VTAIL.n171 585
R1300 VTAIL.n215 VTAIL.n214 585
R1301 VTAIL.n217 VTAIL.n216 585
R1302 VTAIL.n168 VTAIL.n167 585
R1303 VTAIL.n223 VTAIL.n222 585
R1304 VTAIL.n225 VTAIL.n224 585
R1305 VTAIL.n164 VTAIL.n163 585
R1306 VTAIL.n231 VTAIL.n230 585
R1307 VTAIL.n233 VTAIL.n232 585
R1308 VTAIL.n549 VTAIL.n548 585
R1309 VTAIL.n547 VTAIL.n546 585
R1310 VTAIL.n480 VTAIL.n479 585
R1311 VTAIL.n541 VTAIL.n540 585
R1312 VTAIL.n539 VTAIL.n538 585
R1313 VTAIL.n484 VTAIL.n483 585
R1314 VTAIL.n533 VTAIL.n532 585
R1315 VTAIL.n531 VTAIL.n530 585
R1316 VTAIL.n488 VTAIL.n487 585
R1317 VTAIL.n525 VTAIL.n524 585
R1318 VTAIL.n523 VTAIL.n490 585
R1319 VTAIL.n522 VTAIL.n521 585
R1320 VTAIL.n493 VTAIL.n491 585
R1321 VTAIL.n516 VTAIL.n515 585
R1322 VTAIL.n514 VTAIL.n513 585
R1323 VTAIL.n497 VTAIL.n496 585
R1324 VTAIL.n508 VTAIL.n507 585
R1325 VTAIL.n506 VTAIL.n505 585
R1326 VTAIL.n501 VTAIL.n500 585
R1327 VTAIL.n469 VTAIL.n468 585
R1328 VTAIL.n467 VTAIL.n466 585
R1329 VTAIL.n400 VTAIL.n399 585
R1330 VTAIL.n461 VTAIL.n460 585
R1331 VTAIL.n459 VTAIL.n458 585
R1332 VTAIL.n404 VTAIL.n403 585
R1333 VTAIL.n453 VTAIL.n452 585
R1334 VTAIL.n451 VTAIL.n450 585
R1335 VTAIL.n408 VTAIL.n407 585
R1336 VTAIL.n445 VTAIL.n444 585
R1337 VTAIL.n443 VTAIL.n410 585
R1338 VTAIL.n442 VTAIL.n441 585
R1339 VTAIL.n413 VTAIL.n411 585
R1340 VTAIL.n436 VTAIL.n435 585
R1341 VTAIL.n434 VTAIL.n433 585
R1342 VTAIL.n417 VTAIL.n416 585
R1343 VTAIL.n428 VTAIL.n427 585
R1344 VTAIL.n426 VTAIL.n425 585
R1345 VTAIL.n421 VTAIL.n420 585
R1346 VTAIL.n391 VTAIL.n390 585
R1347 VTAIL.n389 VTAIL.n388 585
R1348 VTAIL.n322 VTAIL.n321 585
R1349 VTAIL.n383 VTAIL.n382 585
R1350 VTAIL.n381 VTAIL.n380 585
R1351 VTAIL.n326 VTAIL.n325 585
R1352 VTAIL.n375 VTAIL.n374 585
R1353 VTAIL.n373 VTAIL.n372 585
R1354 VTAIL.n330 VTAIL.n329 585
R1355 VTAIL.n367 VTAIL.n366 585
R1356 VTAIL.n365 VTAIL.n332 585
R1357 VTAIL.n364 VTAIL.n363 585
R1358 VTAIL.n335 VTAIL.n333 585
R1359 VTAIL.n358 VTAIL.n357 585
R1360 VTAIL.n356 VTAIL.n355 585
R1361 VTAIL.n339 VTAIL.n338 585
R1362 VTAIL.n350 VTAIL.n349 585
R1363 VTAIL.n348 VTAIL.n347 585
R1364 VTAIL.n343 VTAIL.n342 585
R1365 VTAIL.n311 VTAIL.n310 585
R1366 VTAIL.n309 VTAIL.n308 585
R1367 VTAIL.n242 VTAIL.n241 585
R1368 VTAIL.n303 VTAIL.n302 585
R1369 VTAIL.n301 VTAIL.n300 585
R1370 VTAIL.n246 VTAIL.n245 585
R1371 VTAIL.n295 VTAIL.n294 585
R1372 VTAIL.n293 VTAIL.n292 585
R1373 VTAIL.n250 VTAIL.n249 585
R1374 VTAIL.n287 VTAIL.n286 585
R1375 VTAIL.n285 VTAIL.n252 585
R1376 VTAIL.n284 VTAIL.n283 585
R1377 VTAIL.n255 VTAIL.n253 585
R1378 VTAIL.n278 VTAIL.n277 585
R1379 VTAIL.n276 VTAIL.n275 585
R1380 VTAIL.n259 VTAIL.n258 585
R1381 VTAIL.n270 VTAIL.n269 585
R1382 VTAIL.n268 VTAIL.n267 585
R1383 VTAIL.n263 VTAIL.n262 585
R1384 VTAIL.n579 VTAIL.t2 329.036
R1385 VTAIL.n27 VTAIL.t6 329.036
R1386 VTAIL.n105 VTAIL.t12 329.036
R1387 VTAIL.n185 VTAIL.t10 329.036
R1388 VTAIL.n422 VTAIL.t9 329.036
R1389 VTAIL.n344 VTAIL.t3 329.036
R1390 VTAIL.n264 VTAIL.t4 329.036
R1391 VTAIL.n502 VTAIL.t13 329.036
R1392 VTAIL.n583 VTAIL.n577 171.744
R1393 VTAIL.n584 VTAIL.n583 171.744
R1394 VTAIL.n584 VTAIL.n573 171.744
R1395 VTAIL.n591 VTAIL.n573 171.744
R1396 VTAIL.n592 VTAIL.n591 171.744
R1397 VTAIL.n592 VTAIL.n569 171.744
R1398 VTAIL.n600 VTAIL.n569 171.744
R1399 VTAIL.n601 VTAIL.n600 171.744
R1400 VTAIL.n602 VTAIL.n601 171.744
R1401 VTAIL.n602 VTAIL.n565 171.744
R1402 VTAIL.n609 VTAIL.n565 171.744
R1403 VTAIL.n610 VTAIL.n609 171.744
R1404 VTAIL.n610 VTAIL.n561 171.744
R1405 VTAIL.n617 VTAIL.n561 171.744
R1406 VTAIL.n618 VTAIL.n617 171.744
R1407 VTAIL.n618 VTAIL.n557 171.744
R1408 VTAIL.n625 VTAIL.n557 171.744
R1409 VTAIL.n626 VTAIL.n625 171.744
R1410 VTAIL.n31 VTAIL.n25 171.744
R1411 VTAIL.n32 VTAIL.n31 171.744
R1412 VTAIL.n32 VTAIL.n21 171.744
R1413 VTAIL.n39 VTAIL.n21 171.744
R1414 VTAIL.n40 VTAIL.n39 171.744
R1415 VTAIL.n40 VTAIL.n17 171.744
R1416 VTAIL.n48 VTAIL.n17 171.744
R1417 VTAIL.n49 VTAIL.n48 171.744
R1418 VTAIL.n50 VTAIL.n49 171.744
R1419 VTAIL.n50 VTAIL.n13 171.744
R1420 VTAIL.n57 VTAIL.n13 171.744
R1421 VTAIL.n58 VTAIL.n57 171.744
R1422 VTAIL.n58 VTAIL.n9 171.744
R1423 VTAIL.n65 VTAIL.n9 171.744
R1424 VTAIL.n66 VTAIL.n65 171.744
R1425 VTAIL.n66 VTAIL.n5 171.744
R1426 VTAIL.n73 VTAIL.n5 171.744
R1427 VTAIL.n74 VTAIL.n73 171.744
R1428 VTAIL.n109 VTAIL.n103 171.744
R1429 VTAIL.n110 VTAIL.n109 171.744
R1430 VTAIL.n110 VTAIL.n99 171.744
R1431 VTAIL.n117 VTAIL.n99 171.744
R1432 VTAIL.n118 VTAIL.n117 171.744
R1433 VTAIL.n118 VTAIL.n95 171.744
R1434 VTAIL.n126 VTAIL.n95 171.744
R1435 VTAIL.n127 VTAIL.n126 171.744
R1436 VTAIL.n128 VTAIL.n127 171.744
R1437 VTAIL.n128 VTAIL.n91 171.744
R1438 VTAIL.n135 VTAIL.n91 171.744
R1439 VTAIL.n136 VTAIL.n135 171.744
R1440 VTAIL.n136 VTAIL.n87 171.744
R1441 VTAIL.n143 VTAIL.n87 171.744
R1442 VTAIL.n144 VTAIL.n143 171.744
R1443 VTAIL.n144 VTAIL.n83 171.744
R1444 VTAIL.n151 VTAIL.n83 171.744
R1445 VTAIL.n152 VTAIL.n151 171.744
R1446 VTAIL.n189 VTAIL.n183 171.744
R1447 VTAIL.n190 VTAIL.n189 171.744
R1448 VTAIL.n190 VTAIL.n179 171.744
R1449 VTAIL.n197 VTAIL.n179 171.744
R1450 VTAIL.n198 VTAIL.n197 171.744
R1451 VTAIL.n198 VTAIL.n175 171.744
R1452 VTAIL.n206 VTAIL.n175 171.744
R1453 VTAIL.n207 VTAIL.n206 171.744
R1454 VTAIL.n208 VTAIL.n207 171.744
R1455 VTAIL.n208 VTAIL.n171 171.744
R1456 VTAIL.n215 VTAIL.n171 171.744
R1457 VTAIL.n216 VTAIL.n215 171.744
R1458 VTAIL.n216 VTAIL.n167 171.744
R1459 VTAIL.n223 VTAIL.n167 171.744
R1460 VTAIL.n224 VTAIL.n223 171.744
R1461 VTAIL.n224 VTAIL.n163 171.744
R1462 VTAIL.n231 VTAIL.n163 171.744
R1463 VTAIL.n232 VTAIL.n231 171.744
R1464 VTAIL.n548 VTAIL.n547 171.744
R1465 VTAIL.n547 VTAIL.n479 171.744
R1466 VTAIL.n540 VTAIL.n479 171.744
R1467 VTAIL.n540 VTAIL.n539 171.744
R1468 VTAIL.n539 VTAIL.n483 171.744
R1469 VTAIL.n532 VTAIL.n483 171.744
R1470 VTAIL.n532 VTAIL.n531 171.744
R1471 VTAIL.n531 VTAIL.n487 171.744
R1472 VTAIL.n524 VTAIL.n487 171.744
R1473 VTAIL.n524 VTAIL.n523 171.744
R1474 VTAIL.n523 VTAIL.n522 171.744
R1475 VTAIL.n522 VTAIL.n491 171.744
R1476 VTAIL.n515 VTAIL.n491 171.744
R1477 VTAIL.n515 VTAIL.n514 171.744
R1478 VTAIL.n514 VTAIL.n496 171.744
R1479 VTAIL.n507 VTAIL.n496 171.744
R1480 VTAIL.n507 VTAIL.n506 171.744
R1481 VTAIL.n506 VTAIL.n500 171.744
R1482 VTAIL.n468 VTAIL.n467 171.744
R1483 VTAIL.n467 VTAIL.n399 171.744
R1484 VTAIL.n460 VTAIL.n399 171.744
R1485 VTAIL.n460 VTAIL.n459 171.744
R1486 VTAIL.n459 VTAIL.n403 171.744
R1487 VTAIL.n452 VTAIL.n403 171.744
R1488 VTAIL.n452 VTAIL.n451 171.744
R1489 VTAIL.n451 VTAIL.n407 171.744
R1490 VTAIL.n444 VTAIL.n407 171.744
R1491 VTAIL.n444 VTAIL.n443 171.744
R1492 VTAIL.n443 VTAIL.n442 171.744
R1493 VTAIL.n442 VTAIL.n411 171.744
R1494 VTAIL.n435 VTAIL.n411 171.744
R1495 VTAIL.n435 VTAIL.n434 171.744
R1496 VTAIL.n434 VTAIL.n416 171.744
R1497 VTAIL.n427 VTAIL.n416 171.744
R1498 VTAIL.n427 VTAIL.n426 171.744
R1499 VTAIL.n426 VTAIL.n420 171.744
R1500 VTAIL.n390 VTAIL.n389 171.744
R1501 VTAIL.n389 VTAIL.n321 171.744
R1502 VTAIL.n382 VTAIL.n321 171.744
R1503 VTAIL.n382 VTAIL.n381 171.744
R1504 VTAIL.n381 VTAIL.n325 171.744
R1505 VTAIL.n374 VTAIL.n325 171.744
R1506 VTAIL.n374 VTAIL.n373 171.744
R1507 VTAIL.n373 VTAIL.n329 171.744
R1508 VTAIL.n366 VTAIL.n329 171.744
R1509 VTAIL.n366 VTAIL.n365 171.744
R1510 VTAIL.n365 VTAIL.n364 171.744
R1511 VTAIL.n364 VTAIL.n333 171.744
R1512 VTAIL.n357 VTAIL.n333 171.744
R1513 VTAIL.n357 VTAIL.n356 171.744
R1514 VTAIL.n356 VTAIL.n338 171.744
R1515 VTAIL.n349 VTAIL.n338 171.744
R1516 VTAIL.n349 VTAIL.n348 171.744
R1517 VTAIL.n348 VTAIL.n342 171.744
R1518 VTAIL.n310 VTAIL.n309 171.744
R1519 VTAIL.n309 VTAIL.n241 171.744
R1520 VTAIL.n302 VTAIL.n241 171.744
R1521 VTAIL.n302 VTAIL.n301 171.744
R1522 VTAIL.n301 VTAIL.n245 171.744
R1523 VTAIL.n294 VTAIL.n245 171.744
R1524 VTAIL.n294 VTAIL.n293 171.744
R1525 VTAIL.n293 VTAIL.n249 171.744
R1526 VTAIL.n286 VTAIL.n249 171.744
R1527 VTAIL.n286 VTAIL.n285 171.744
R1528 VTAIL.n285 VTAIL.n284 171.744
R1529 VTAIL.n284 VTAIL.n253 171.744
R1530 VTAIL.n277 VTAIL.n253 171.744
R1531 VTAIL.n277 VTAIL.n276 171.744
R1532 VTAIL.n276 VTAIL.n258 171.744
R1533 VTAIL.n269 VTAIL.n258 171.744
R1534 VTAIL.n269 VTAIL.n268 171.744
R1535 VTAIL.n268 VTAIL.n262 171.744
R1536 VTAIL.t2 VTAIL.n577 85.8723
R1537 VTAIL.t6 VTAIL.n25 85.8723
R1538 VTAIL.t12 VTAIL.n103 85.8723
R1539 VTAIL.t10 VTAIL.n183 85.8723
R1540 VTAIL.t13 VTAIL.n500 85.8723
R1541 VTAIL.t9 VTAIL.n420 85.8723
R1542 VTAIL.t3 VTAIL.n342 85.8723
R1543 VTAIL.t4 VTAIL.n262 85.8723
R1544 VTAIL.n1 VTAIL.n0 53.7905
R1545 VTAIL.n159 VTAIL.n158 53.7905
R1546 VTAIL.n475 VTAIL.n474 53.7905
R1547 VTAIL.n317 VTAIL.n316 53.7905
R1548 VTAIL.n631 VTAIL.n630 31.0217
R1549 VTAIL.n79 VTAIL.n78 31.0217
R1550 VTAIL.n157 VTAIL.n156 31.0217
R1551 VTAIL.n237 VTAIL.n236 31.0217
R1552 VTAIL.n553 VTAIL.n552 31.0217
R1553 VTAIL.n473 VTAIL.n472 31.0217
R1554 VTAIL.n395 VTAIL.n394 31.0217
R1555 VTAIL.n315 VTAIL.n314 31.0217
R1556 VTAIL.n631 VTAIL.n553 26.3841
R1557 VTAIL.n315 VTAIL.n237 26.3841
R1558 VTAIL.n603 VTAIL.n568 13.1884
R1559 VTAIL.n51 VTAIL.n16 13.1884
R1560 VTAIL.n129 VTAIL.n94 13.1884
R1561 VTAIL.n209 VTAIL.n174 13.1884
R1562 VTAIL.n525 VTAIL.n490 13.1884
R1563 VTAIL.n445 VTAIL.n410 13.1884
R1564 VTAIL.n367 VTAIL.n332 13.1884
R1565 VTAIL.n287 VTAIL.n252 13.1884
R1566 VTAIL.n599 VTAIL.n598 12.8005
R1567 VTAIL.n604 VTAIL.n566 12.8005
R1568 VTAIL.n47 VTAIL.n46 12.8005
R1569 VTAIL.n52 VTAIL.n14 12.8005
R1570 VTAIL.n125 VTAIL.n124 12.8005
R1571 VTAIL.n130 VTAIL.n92 12.8005
R1572 VTAIL.n205 VTAIL.n204 12.8005
R1573 VTAIL.n210 VTAIL.n172 12.8005
R1574 VTAIL.n526 VTAIL.n488 12.8005
R1575 VTAIL.n521 VTAIL.n492 12.8005
R1576 VTAIL.n446 VTAIL.n408 12.8005
R1577 VTAIL.n441 VTAIL.n412 12.8005
R1578 VTAIL.n368 VTAIL.n330 12.8005
R1579 VTAIL.n363 VTAIL.n334 12.8005
R1580 VTAIL.n288 VTAIL.n250 12.8005
R1581 VTAIL.n283 VTAIL.n254 12.8005
R1582 VTAIL.n597 VTAIL.n570 12.0247
R1583 VTAIL.n608 VTAIL.n607 12.0247
R1584 VTAIL.n45 VTAIL.n18 12.0247
R1585 VTAIL.n56 VTAIL.n55 12.0247
R1586 VTAIL.n123 VTAIL.n96 12.0247
R1587 VTAIL.n134 VTAIL.n133 12.0247
R1588 VTAIL.n203 VTAIL.n176 12.0247
R1589 VTAIL.n214 VTAIL.n213 12.0247
R1590 VTAIL.n530 VTAIL.n529 12.0247
R1591 VTAIL.n520 VTAIL.n493 12.0247
R1592 VTAIL.n450 VTAIL.n449 12.0247
R1593 VTAIL.n440 VTAIL.n413 12.0247
R1594 VTAIL.n372 VTAIL.n371 12.0247
R1595 VTAIL.n362 VTAIL.n335 12.0247
R1596 VTAIL.n292 VTAIL.n291 12.0247
R1597 VTAIL.n282 VTAIL.n255 12.0247
R1598 VTAIL.n594 VTAIL.n593 11.249
R1599 VTAIL.n611 VTAIL.n564 11.249
R1600 VTAIL.n42 VTAIL.n41 11.249
R1601 VTAIL.n59 VTAIL.n12 11.249
R1602 VTAIL.n120 VTAIL.n119 11.249
R1603 VTAIL.n137 VTAIL.n90 11.249
R1604 VTAIL.n200 VTAIL.n199 11.249
R1605 VTAIL.n217 VTAIL.n170 11.249
R1606 VTAIL.n533 VTAIL.n486 11.249
R1607 VTAIL.n517 VTAIL.n516 11.249
R1608 VTAIL.n453 VTAIL.n406 11.249
R1609 VTAIL.n437 VTAIL.n436 11.249
R1610 VTAIL.n375 VTAIL.n328 11.249
R1611 VTAIL.n359 VTAIL.n358 11.249
R1612 VTAIL.n295 VTAIL.n248 11.249
R1613 VTAIL.n279 VTAIL.n278 11.249
R1614 VTAIL.n579 VTAIL.n578 10.7239
R1615 VTAIL.n27 VTAIL.n26 10.7239
R1616 VTAIL.n105 VTAIL.n104 10.7239
R1617 VTAIL.n185 VTAIL.n184 10.7239
R1618 VTAIL.n502 VTAIL.n501 10.7239
R1619 VTAIL.n422 VTAIL.n421 10.7239
R1620 VTAIL.n344 VTAIL.n343 10.7239
R1621 VTAIL.n264 VTAIL.n263 10.7239
R1622 VTAIL.n590 VTAIL.n572 10.4732
R1623 VTAIL.n612 VTAIL.n562 10.4732
R1624 VTAIL.n38 VTAIL.n20 10.4732
R1625 VTAIL.n60 VTAIL.n10 10.4732
R1626 VTAIL.n116 VTAIL.n98 10.4732
R1627 VTAIL.n138 VTAIL.n88 10.4732
R1628 VTAIL.n196 VTAIL.n178 10.4732
R1629 VTAIL.n218 VTAIL.n168 10.4732
R1630 VTAIL.n534 VTAIL.n484 10.4732
R1631 VTAIL.n513 VTAIL.n495 10.4732
R1632 VTAIL.n454 VTAIL.n404 10.4732
R1633 VTAIL.n433 VTAIL.n415 10.4732
R1634 VTAIL.n376 VTAIL.n326 10.4732
R1635 VTAIL.n355 VTAIL.n337 10.4732
R1636 VTAIL.n296 VTAIL.n246 10.4732
R1637 VTAIL.n275 VTAIL.n257 10.4732
R1638 VTAIL.n589 VTAIL.n574 9.69747
R1639 VTAIL.n616 VTAIL.n615 9.69747
R1640 VTAIL.n37 VTAIL.n22 9.69747
R1641 VTAIL.n64 VTAIL.n63 9.69747
R1642 VTAIL.n115 VTAIL.n100 9.69747
R1643 VTAIL.n142 VTAIL.n141 9.69747
R1644 VTAIL.n195 VTAIL.n180 9.69747
R1645 VTAIL.n222 VTAIL.n221 9.69747
R1646 VTAIL.n538 VTAIL.n537 9.69747
R1647 VTAIL.n512 VTAIL.n497 9.69747
R1648 VTAIL.n458 VTAIL.n457 9.69747
R1649 VTAIL.n432 VTAIL.n417 9.69747
R1650 VTAIL.n380 VTAIL.n379 9.69747
R1651 VTAIL.n354 VTAIL.n339 9.69747
R1652 VTAIL.n300 VTAIL.n299 9.69747
R1653 VTAIL.n274 VTAIL.n259 9.69747
R1654 VTAIL.n630 VTAIL.n629 9.45567
R1655 VTAIL.n78 VTAIL.n77 9.45567
R1656 VTAIL.n156 VTAIL.n155 9.45567
R1657 VTAIL.n236 VTAIL.n235 9.45567
R1658 VTAIL.n552 VTAIL.n551 9.45567
R1659 VTAIL.n472 VTAIL.n471 9.45567
R1660 VTAIL.n394 VTAIL.n393 9.45567
R1661 VTAIL.n314 VTAIL.n313 9.45567
R1662 VTAIL.n556 VTAIL.n555 9.3005
R1663 VTAIL.n629 VTAIL.n628 9.3005
R1664 VTAIL.n621 VTAIL.n620 9.3005
R1665 VTAIL.n560 VTAIL.n559 9.3005
R1666 VTAIL.n615 VTAIL.n614 9.3005
R1667 VTAIL.n613 VTAIL.n612 9.3005
R1668 VTAIL.n564 VTAIL.n563 9.3005
R1669 VTAIL.n607 VTAIL.n606 9.3005
R1670 VTAIL.n605 VTAIL.n604 9.3005
R1671 VTAIL.n581 VTAIL.n580 9.3005
R1672 VTAIL.n576 VTAIL.n575 9.3005
R1673 VTAIL.n587 VTAIL.n586 9.3005
R1674 VTAIL.n589 VTAIL.n588 9.3005
R1675 VTAIL.n572 VTAIL.n571 9.3005
R1676 VTAIL.n595 VTAIL.n594 9.3005
R1677 VTAIL.n597 VTAIL.n596 9.3005
R1678 VTAIL.n598 VTAIL.n567 9.3005
R1679 VTAIL.n623 VTAIL.n622 9.3005
R1680 VTAIL.n4 VTAIL.n3 9.3005
R1681 VTAIL.n77 VTAIL.n76 9.3005
R1682 VTAIL.n69 VTAIL.n68 9.3005
R1683 VTAIL.n8 VTAIL.n7 9.3005
R1684 VTAIL.n63 VTAIL.n62 9.3005
R1685 VTAIL.n61 VTAIL.n60 9.3005
R1686 VTAIL.n12 VTAIL.n11 9.3005
R1687 VTAIL.n55 VTAIL.n54 9.3005
R1688 VTAIL.n53 VTAIL.n52 9.3005
R1689 VTAIL.n29 VTAIL.n28 9.3005
R1690 VTAIL.n24 VTAIL.n23 9.3005
R1691 VTAIL.n35 VTAIL.n34 9.3005
R1692 VTAIL.n37 VTAIL.n36 9.3005
R1693 VTAIL.n20 VTAIL.n19 9.3005
R1694 VTAIL.n43 VTAIL.n42 9.3005
R1695 VTAIL.n45 VTAIL.n44 9.3005
R1696 VTAIL.n46 VTAIL.n15 9.3005
R1697 VTAIL.n71 VTAIL.n70 9.3005
R1698 VTAIL.n82 VTAIL.n81 9.3005
R1699 VTAIL.n155 VTAIL.n154 9.3005
R1700 VTAIL.n147 VTAIL.n146 9.3005
R1701 VTAIL.n86 VTAIL.n85 9.3005
R1702 VTAIL.n141 VTAIL.n140 9.3005
R1703 VTAIL.n139 VTAIL.n138 9.3005
R1704 VTAIL.n90 VTAIL.n89 9.3005
R1705 VTAIL.n133 VTAIL.n132 9.3005
R1706 VTAIL.n131 VTAIL.n130 9.3005
R1707 VTAIL.n107 VTAIL.n106 9.3005
R1708 VTAIL.n102 VTAIL.n101 9.3005
R1709 VTAIL.n113 VTAIL.n112 9.3005
R1710 VTAIL.n115 VTAIL.n114 9.3005
R1711 VTAIL.n98 VTAIL.n97 9.3005
R1712 VTAIL.n121 VTAIL.n120 9.3005
R1713 VTAIL.n123 VTAIL.n122 9.3005
R1714 VTAIL.n124 VTAIL.n93 9.3005
R1715 VTAIL.n149 VTAIL.n148 9.3005
R1716 VTAIL.n162 VTAIL.n161 9.3005
R1717 VTAIL.n235 VTAIL.n234 9.3005
R1718 VTAIL.n227 VTAIL.n226 9.3005
R1719 VTAIL.n166 VTAIL.n165 9.3005
R1720 VTAIL.n221 VTAIL.n220 9.3005
R1721 VTAIL.n219 VTAIL.n218 9.3005
R1722 VTAIL.n170 VTAIL.n169 9.3005
R1723 VTAIL.n213 VTAIL.n212 9.3005
R1724 VTAIL.n211 VTAIL.n210 9.3005
R1725 VTAIL.n187 VTAIL.n186 9.3005
R1726 VTAIL.n182 VTAIL.n181 9.3005
R1727 VTAIL.n193 VTAIL.n192 9.3005
R1728 VTAIL.n195 VTAIL.n194 9.3005
R1729 VTAIL.n178 VTAIL.n177 9.3005
R1730 VTAIL.n201 VTAIL.n200 9.3005
R1731 VTAIL.n203 VTAIL.n202 9.3005
R1732 VTAIL.n204 VTAIL.n173 9.3005
R1733 VTAIL.n229 VTAIL.n228 9.3005
R1734 VTAIL.n478 VTAIL.n477 9.3005
R1735 VTAIL.n545 VTAIL.n544 9.3005
R1736 VTAIL.n543 VTAIL.n542 9.3005
R1737 VTAIL.n482 VTAIL.n481 9.3005
R1738 VTAIL.n537 VTAIL.n536 9.3005
R1739 VTAIL.n535 VTAIL.n534 9.3005
R1740 VTAIL.n486 VTAIL.n485 9.3005
R1741 VTAIL.n529 VTAIL.n528 9.3005
R1742 VTAIL.n527 VTAIL.n526 9.3005
R1743 VTAIL.n492 VTAIL.n489 9.3005
R1744 VTAIL.n520 VTAIL.n519 9.3005
R1745 VTAIL.n518 VTAIL.n517 9.3005
R1746 VTAIL.n495 VTAIL.n494 9.3005
R1747 VTAIL.n512 VTAIL.n511 9.3005
R1748 VTAIL.n510 VTAIL.n509 9.3005
R1749 VTAIL.n499 VTAIL.n498 9.3005
R1750 VTAIL.n504 VTAIL.n503 9.3005
R1751 VTAIL.n551 VTAIL.n550 9.3005
R1752 VTAIL.n424 VTAIL.n423 9.3005
R1753 VTAIL.n419 VTAIL.n418 9.3005
R1754 VTAIL.n430 VTAIL.n429 9.3005
R1755 VTAIL.n432 VTAIL.n431 9.3005
R1756 VTAIL.n415 VTAIL.n414 9.3005
R1757 VTAIL.n438 VTAIL.n437 9.3005
R1758 VTAIL.n440 VTAIL.n439 9.3005
R1759 VTAIL.n412 VTAIL.n409 9.3005
R1760 VTAIL.n471 VTAIL.n470 9.3005
R1761 VTAIL.n398 VTAIL.n397 9.3005
R1762 VTAIL.n465 VTAIL.n464 9.3005
R1763 VTAIL.n463 VTAIL.n462 9.3005
R1764 VTAIL.n402 VTAIL.n401 9.3005
R1765 VTAIL.n457 VTAIL.n456 9.3005
R1766 VTAIL.n455 VTAIL.n454 9.3005
R1767 VTAIL.n406 VTAIL.n405 9.3005
R1768 VTAIL.n449 VTAIL.n448 9.3005
R1769 VTAIL.n447 VTAIL.n446 9.3005
R1770 VTAIL.n346 VTAIL.n345 9.3005
R1771 VTAIL.n341 VTAIL.n340 9.3005
R1772 VTAIL.n352 VTAIL.n351 9.3005
R1773 VTAIL.n354 VTAIL.n353 9.3005
R1774 VTAIL.n337 VTAIL.n336 9.3005
R1775 VTAIL.n360 VTAIL.n359 9.3005
R1776 VTAIL.n362 VTAIL.n361 9.3005
R1777 VTAIL.n334 VTAIL.n331 9.3005
R1778 VTAIL.n393 VTAIL.n392 9.3005
R1779 VTAIL.n320 VTAIL.n319 9.3005
R1780 VTAIL.n387 VTAIL.n386 9.3005
R1781 VTAIL.n385 VTAIL.n384 9.3005
R1782 VTAIL.n324 VTAIL.n323 9.3005
R1783 VTAIL.n379 VTAIL.n378 9.3005
R1784 VTAIL.n377 VTAIL.n376 9.3005
R1785 VTAIL.n328 VTAIL.n327 9.3005
R1786 VTAIL.n371 VTAIL.n370 9.3005
R1787 VTAIL.n369 VTAIL.n368 9.3005
R1788 VTAIL.n266 VTAIL.n265 9.3005
R1789 VTAIL.n261 VTAIL.n260 9.3005
R1790 VTAIL.n272 VTAIL.n271 9.3005
R1791 VTAIL.n274 VTAIL.n273 9.3005
R1792 VTAIL.n257 VTAIL.n256 9.3005
R1793 VTAIL.n280 VTAIL.n279 9.3005
R1794 VTAIL.n282 VTAIL.n281 9.3005
R1795 VTAIL.n254 VTAIL.n251 9.3005
R1796 VTAIL.n313 VTAIL.n312 9.3005
R1797 VTAIL.n240 VTAIL.n239 9.3005
R1798 VTAIL.n307 VTAIL.n306 9.3005
R1799 VTAIL.n305 VTAIL.n304 9.3005
R1800 VTAIL.n244 VTAIL.n243 9.3005
R1801 VTAIL.n299 VTAIL.n298 9.3005
R1802 VTAIL.n297 VTAIL.n296 9.3005
R1803 VTAIL.n248 VTAIL.n247 9.3005
R1804 VTAIL.n291 VTAIL.n290 9.3005
R1805 VTAIL.n289 VTAIL.n288 9.3005
R1806 VTAIL.n586 VTAIL.n585 8.92171
R1807 VTAIL.n619 VTAIL.n560 8.92171
R1808 VTAIL.n34 VTAIL.n33 8.92171
R1809 VTAIL.n67 VTAIL.n8 8.92171
R1810 VTAIL.n112 VTAIL.n111 8.92171
R1811 VTAIL.n145 VTAIL.n86 8.92171
R1812 VTAIL.n192 VTAIL.n191 8.92171
R1813 VTAIL.n225 VTAIL.n166 8.92171
R1814 VTAIL.n541 VTAIL.n482 8.92171
R1815 VTAIL.n509 VTAIL.n508 8.92171
R1816 VTAIL.n461 VTAIL.n402 8.92171
R1817 VTAIL.n429 VTAIL.n428 8.92171
R1818 VTAIL.n383 VTAIL.n324 8.92171
R1819 VTAIL.n351 VTAIL.n350 8.92171
R1820 VTAIL.n303 VTAIL.n244 8.92171
R1821 VTAIL.n271 VTAIL.n270 8.92171
R1822 VTAIL.n582 VTAIL.n576 8.14595
R1823 VTAIL.n620 VTAIL.n558 8.14595
R1824 VTAIL.n630 VTAIL.n554 8.14595
R1825 VTAIL.n30 VTAIL.n24 8.14595
R1826 VTAIL.n68 VTAIL.n6 8.14595
R1827 VTAIL.n78 VTAIL.n2 8.14595
R1828 VTAIL.n108 VTAIL.n102 8.14595
R1829 VTAIL.n146 VTAIL.n84 8.14595
R1830 VTAIL.n156 VTAIL.n80 8.14595
R1831 VTAIL.n188 VTAIL.n182 8.14595
R1832 VTAIL.n226 VTAIL.n164 8.14595
R1833 VTAIL.n236 VTAIL.n160 8.14595
R1834 VTAIL.n552 VTAIL.n476 8.14595
R1835 VTAIL.n542 VTAIL.n480 8.14595
R1836 VTAIL.n505 VTAIL.n499 8.14595
R1837 VTAIL.n472 VTAIL.n396 8.14595
R1838 VTAIL.n462 VTAIL.n400 8.14595
R1839 VTAIL.n425 VTAIL.n419 8.14595
R1840 VTAIL.n394 VTAIL.n318 8.14595
R1841 VTAIL.n384 VTAIL.n322 8.14595
R1842 VTAIL.n347 VTAIL.n341 8.14595
R1843 VTAIL.n314 VTAIL.n238 8.14595
R1844 VTAIL.n304 VTAIL.n242 8.14595
R1845 VTAIL.n267 VTAIL.n261 8.14595
R1846 VTAIL.n581 VTAIL.n578 7.3702
R1847 VTAIL.n624 VTAIL.n623 7.3702
R1848 VTAIL.n628 VTAIL.n627 7.3702
R1849 VTAIL.n29 VTAIL.n26 7.3702
R1850 VTAIL.n72 VTAIL.n71 7.3702
R1851 VTAIL.n76 VTAIL.n75 7.3702
R1852 VTAIL.n107 VTAIL.n104 7.3702
R1853 VTAIL.n150 VTAIL.n149 7.3702
R1854 VTAIL.n154 VTAIL.n153 7.3702
R1855 VTAIL.n187 VTAIL.n184 7.3702
R1856 VTAIL.n230 VTAIL.n229 7.3702
R1857 VTAIL.n234 VTAIL.n233 7.3702
R1858 VTAIL.n550 VTAIL.n549 7.3702
R1859 VTAIL.n546 VTAIL.n545 7.3702
R1860 VTAIL.n504 VTAIL.n501 7.3702
R1861 VTAIL.n470 VTAIL.n469 7.3702
R1862 VTAIL.n466 VTAIL.n465 7.3702
R1863 VTAIL.n424 VTAIL.n421 7.3702
R1864 VTAIL.n392 VTAIL.n391 7.3702
R1865 VTAIL.n388 VTAIL.n387 7.3702
R1866 VTAIL.n346 VTAIL.n343 7.3702
R1867 VTAIL.n312 VTAIL.n311 7.3702
R1868 VTAIL.n308 VTAIL.n307 7.3702
R1869 VTAIL.n266 VTAIL.n263 7.3702
R1870 VTAIL.n624 VTAIL.n556 6.59444
R1871 VTAIL.n627 VTAIL.n556 6.59444
R1872 VTAIL.n72 VTAIL.n4 6.59444
R1873 VTAIL.n75 VTAIL.n4 6.59444
R1874 VTAIL.n150 VTAIL.n82 6.59444
R1875 VTAIL.n153 VTAIL.n82 6.59444
R1876 VTAIL.n230 VTAIL.n162 6.59444
R1877 VTAIL.n233 VTAIL.n162 6.59444
R1878 VTAIL.n549 VTAIL.n478 6.59444
R1879 VTAIL.n546 VTAIL.n478 6.59444
R1880 VTAIL.n469 VTAIL.n398 6.59444
R1881 VTAIL.n466 VTAIL.n398 6.59444
R1882 VTAIL.n391 VTAIL.n320 6.59444
R1883 VTAIL.n388 VTAIL.n320 6.59444
R1884 VTAIL.n311 VTAIL.n240 6.59444
R1885 VTAIL.n308 VTAIL.n240 6.59444
R1886 VTAIL.n582 VTAIL.n581 5.81868
R1887 VTAIL.n623 VTAIL.n558 5.81868
R1888 VTAIL.n628 VTAIL.n554 5.81868
R1889 VTAIL.n30 VTAIL.n29 5.81868
R1890 VTAIL.n71 VTAIL.n6 5.81868
R1891 VTAIL.n76 VTAIL.n2 5.81868
R1892 VTAIL.n108 VTAIL.n107 5.81868
R1893 VTAIL.n149 VTAIL.n84 5.81868
R1894 VTAIL.n154 VTAIL.n80 5.81868
R1895 VTAIL.n188 VTAIL.n187 5.81868
R1896 VTAIL.n229 VTAIL.n164 5.81868
R1897 VTAIL.n234 VTAIL.n160 5.81868
R1898 VTAIL.n550 VTAIL.n476 5.81868
R1899 VTAIL.n545 VTAIL.n480 5.81868
R1900 VTAIL.n505 VTAIL.n504 5.81868
R1901 VTAIL.n470 VTAIL.n396 5.81868
R1902 VTAIL.n465 VTAIL.n400 5.81868
R1903 VTAIL.n425 VTAIL.n424 5.81868
R1904 VTAIL.n392 VTAIL.n318 5.81868
R1905 VTAIL.n387 VTAIL.n322 5.81868
R1906 VTAIL.n347 VTAIL.n346 5.81868
R1907 VTAIL.n312 VTAIL.n238 5.81868
R1908 VTAIL.n307 VTAIL.n242 5.81868
R1909 VTAIL.n267 VTAIL.n266 5.81868
R1910 VTAIL.n585 VTAIL.n576 5.04292
R1911 VTAIL.n620 VTAIL.n619 5.04292
R1912 VTAIL.n33 VTAIL.n24 5.04292
R1913 VTAIL.n68 VTAIL.n67 5.04292
R1914 VTAIL.n111 VTAIL.n102 5.04292
R1915 VTAIL.n146 VTAIL.n145 5.04292
R1916 VTAIL.n191 VTAIL.n182 5.04292
R1917 VTAIL.n226 VTAIL.n225 5.04292
R1918 VTAIL.n542 VTAIL.n541 5.04292
R1919 VTAIL.n508 VTAIL.n499 5.04292
R1920 VTAIL.n462 VTAIL.n461 5.04292
R1921 VTAIL.n428 VTAIL.n419 5.04292
R1922 VTAIL.n384 VTAIL.n383 5.04292
R1923 VTAIL.n350 VTAIL.n341 5.04292
R1924 VTAIL.n304 VTAIL.n303 5.04292
R1925 VTAIL.n270 VTAIL.n261 5.04292
R1926 VTAIL.n586 VTAIL.n574 4.26717
R1927 VTAIL.n616 VTAIL.n560 4.26717
R1928 VTAIL.n34 VTAIL.n22 4.26717
R1929 VTAIL.n64 VTAIL.n8 4.26717
R1930 VTAIL.n112 VTAIL.n100 4.26717
R1931 VTAIL.n142 VTAIL.n86 4.26717
R1932 VTAIL.n192 VTAIL.n180 4.26717
R1933 VTAIL.n222 VTAIL.n166 4.26717
R1934 VTAIL.n538 VTAIL.n482 4.26717
R1935 VTAIL.n509 VTAIL.n497 4.26717
R1936 VTAIL.n458 VTAIL.n402 4.26717
R1937 VTAIL.n429 VTAIL.n417 4.26717
R1938 VTAIL.n380 VTAIL.n324 4.26717
R1939 VTAIL.n351 VTAIL.n339 4.26717
R1940 VTAIL.n300 VTAIL.n244 4.26717
R1941 VTAIL.n271 VTAIL.n259 4.26717
R1942 VTAIL.n590 VTAIL.n589 3.49141
R1943 VTAIL.n615 VTAIL.n562 3.49141
R1944 VTAIL.n38 VTAIL.n37 3.49141
R1945 VTAIL.n63 VTAIL.n10 3.49141
R1946 VTAIL.n116 VTAIL.n115 3.49141
R1947 VTAIL.n141 VTAIL.n88 3.49141
R1948 VTAIL.n196 VTAIL.n195 3.49141
R1949 VTAIL.n221 VTAIL.n168 3.49141
R1950 VTAIL.n537 VTAIL.n484 3.49141
R1951 VTAIL.n513 VTAIL.n512 3.49141
R1952 VTAIL.n457 VTAIL.n404 3.49141
R1953 VTAIL.n433 VTAIL.n432 3.49141
R1954 VTAIL.n379 VTAIL.n326 3.49141
R1955 VTAIL.n355 VTAIL.n354 3.49141
R1956 VTAIL.n299 VTAIL.n246 3.49141
R1957 VTAIL.n275 VTAIL.n274 3.49141
R1958 VTAIL.n593 VTAIL.n572 2.71565
R1959 VTAIL.n612 VTAIL.n611 2.71565
R1960 VTAIL.n41 VTAIL.n20 2.71565
R1961 VTAIL.n60 VTAIL.n59 2.71565
R1962 VTAIL.n119 VTAIL.n98 2.71565
R1963 VTAIL.n138 VTAIL.n137 2.71565
R1964 VTAIL.n199 VTAIL.n178 2.71565
R1965 VTAIL.n218 VTAIL.n217 2.71565
R1966 VTAIL.n534 VTAIL.n533 2.71565
R1967 VTAIL.n516 VTAIL.n495 2.71565
R1968 VTAIL.n454 VTAIL.n453 2.71565
R1969 VTAIL.n436 VTAIL.n415 2.71565
R1970 VTAIL.n376 VTAIL.n375 2.71565
R1971 VTAIL.n358 VTAIL.n337 2.71565
R1972 VTAIL.n296 VTAIL.n295 2.71565
R1973 VTAIL.n278 VTAIL.n257 2.71565
R1974 VTAIL.n503 VTAIL.n502 2.41282
R1975 VTAIL.n423 VTAIL.n422 2.41282
R1976 VTAIL.n345 VTAIL.n344 2.41282
R1977 VTAIL.n265 VTAIL.n264 2.41282
R1978 VTAIL.n580 VTAIL.n579 2.41282
R1979 VTAIL.n28 VTAIL.n27 2.41282
R1980 VTAIL.n106 VTAIL.n105 2.41282
R1981 VTAIL.n186 VTAIL.n185 2.41282
R1982 VTAIL.n0 VTAIL.t1 2.28637
R1983 VTAIL.n0 VTAIL.t5 2.28637
R1984 VTAIL.n158 VTAIL.t8 2.28637
R1985 VTAIL.n158 VTAIL.t11 2.28637
R1986 VTAIL.n474 VTAIL.t7 2.28637
R1987 VTAIL.n474 VTAIL.t14 2.28637
R1988 VTAIL.n316 VTAIL.t0 2.28637
R1989 VTAIL.n316 VTAIL.t15 2.28637
R1990 VTAIL.n594 VTAIL.n570 1.93989
R1991 VTAIL.n608 VTAIL.n564 1.93989
R1992 VTAIL.n42 VTAIL.n18 1.93989
R1993 VTAIL.n56 VTAIL.n12 1.93989
R1994 VTAIL.n120 VTAIL.n96 1.93989
R1995 VTAIL.n134 VTAIL.n90 1.93989
R1996 VTAIL.n200 VTAIL.n176 1.93989
R1997 VTAIL.n214 VTAIL.n170 1.93989
R1998 VTAIL.n530 VTAIL.n486 1.93989
R1999 VTAIL.n517 VTAIL.n493 1.93989
R2000 VTAIL.n450 VTAIL.n406 1.93989
R2001 VTAIL.n437 VTAIL.n413 1.93989
R2002 VTAIL.n372 VTAIL.n328 1.93989
R2003 VTAIL.n359 VTAIL.n335 1.93989
R2004 VTAIL.n292 VTAIL.n248 1.93989
R2005 VTAIL.n279 VTAIL.n255 1.93989
R2006 VTAIL.n317 VTAIL.n315 1.75912
R2007 VTAIL.n395 VTAIL.n317 1.75912
R2008 VTAIL.n475 VTAIL.n473 1.75912
R2009 VTAIL.n553 VTAIL.n475 1.75912
R2010 VTAIL.n237 VTAIL.n159 1.75912
R2011 VTAIL.n159 VTAIL.n157 1.75912
R2012 VTAIL.n79 VTAIL.n1 1.75912
R2013 VTAIL VTAIL.n631 1.70093
R2014 VTAIL.n599 VTAIL.n597 1.16414
R2015 VTAIL.n607 VTAIL.n566 1.16414
R2016 VTAIL.n47 VTAIL.n45 1.16414
R2017 VTAIL.n55 VTAIL.n14 1.16414
R2018 VTAIL.n125 VTAIL.n123 1.16414
R2019 VTAIL.n133 VTAIL.n92 1.16414
R2020 VTAIL.n205 VTAIL.n203 1.16414
R2021 VTAIL.n213 VTAIL.n172 1.16414
R2022 VTAIL.n529 VTAIL.n488 1.16414
R2023 VTAIL.n521 VTAIL.n520 1.16414
R2024 VTAIL.n449 VTAIL.n408 1.16414
R2025 VTAIL.n441 VTAIL.n440 1.16414
R2026 VTAIL.n371 VTAIL.n330 1.16414
R2027 VTAIL.n363 VTAIL.n362 1.16414
R2028 VTAIL.n291 VTAIL.n250 1.16414
R2029 VTAIL.n283 VTAIL.n282 1.16414
R2030 VTAIL.n473 VTAIL.n395 0.470328
R2031 VTAIL.n157 VTAIL.n79 0.470328
R2032 VTAIL.n598 VTAIL.n568 0.388379
R2033 VTAIL.n604 VTAIL.n603 0.388379
R2034 VTAIL.n46 VTAIL.n16 0.388379
R2035 VTAIL.n52 VTAIL.n51 0.388379
R2036 VTAIL.n124 VTAIL.n94 0.388379
R2037 VTAIL.n130 VTAIL.n129 0.388379
R2038 VTAIL.n204 VTAIL.n174 0.388379
R2039 VTAIL.n210 VTAIL.n209 0.388379
R2040 VTAIL.n526 VTAIL.n525 0.388379
R2041 VTAIL.n492 VTAIL.n490 0.388379
R2042 VTAIL.n446 VTAIL.n445 0.388379
R2043 VTAIL.n412 VTAIL.n410 0.388379
R2044 VTAIL.n368 VTAIL.n367 0.388379
R2045 VTAIL.n334 VTAIL.n332 0.388379
R2046 VTAIL.n288 VTAIL.n287 0.388379
R2047 VTAIL.n254 VTAIL.n252 0.388379
R2048 VTAIL.n580 VTAIL.n575 0.155672
R2049 VTAIL.n587 VTAIL.n575 0.155672
R2050 VTAIL.n588 VTAIL.n587 0.155672
R2051 VTAIL.n588 VTAIL.n571 0.155672
R2052 VTAIL.n595 VTAIL.n571 0.155672
R2053 VTAIL.n596 VTAIL.n595 0.155672
R2054 VTAIL.n596 VTAIL.n567 0.155672
R2055 VTAIL.n605 VTAIL.n567 0.155672
R2056 VTAIL.n606 VTAIL.n605 0.155672
R2057 VTAIL.n606 VTAIL.n563 0.155672
R2058 VTAIL.n613 VTAIL.n563 0.155672
R2059 VTAIL.n614 VTAIL.n613 0.155672
R2060 VTAIL.n614 VTAIL.n559 0.155672
R2061 VTAIL.n621 VTAIL.n559 0.155672
R2062 VTAIL.n622 VTAIL.n621 0.155672
R2063 VTAIL.n622 VTAIL.n555 0.155672
R2064 VTAIL.n629 VTAIL.n555 0.155672
R2065 VTAIL.n28 VTAIL.n23 0.155672
R2066 VTAIL.n35 VTAIL.n23 0.155672
R2067 VTAIL.n36 VTAIL.n35 0.155672
R2068 VTAIL.n36 VTAIL.n19 0.155672
R2069 VTAIL.n43 VTAIL.n19 0.155672
R2070 VTAIL.n44 VTAIL.n43 0.155672
R2071 VTAIL.n44 VTAIL.n15 0.155672
R2072 VTAIL.n53 VTAIL.n15 0.155672
R2073 VTAIL.n54 VTAIL.n53 0.155672
R2074 VTAIL.n54 VTAIL.n11 0.155672
R2075 VTAIL.n61 VTAIL.n11 0.155672
R2076 VTAIL.n62 VTAIL.n61 0.155672
R2077 VTAIL.n62 VTAIL.n7 0.155672
R2078 VTAIL.n69 VTAIL.n7 0.155672
R2079 VTAIL.n70 VTAIL.n69 0.155672
R2080 VTAIL.n70 VTAIL.n3 0.155672
R2081 VTAIL.n77 VTAIL.n3 0.155672
R2082 VTAIL.n106 VTAIL.n101 0.155672
R2083 VTAIL.n113 VTAIL.n101 0.155672
R2084 VTAIL.n114 VTAIL.n113 0.155672
R2085 VTAIL.n114 VTAIL.n97 0.155672
R2086 VTAIL.n121 VTAIL.n97 0.155672
R2087 VTAIL.n122 VTAIL.n121 0.155672
R2088 VTAIL.n122 VTAIL.n93 0.155672
R2089 VTAIL.n131 VTAIL.n93 0.155672
R2090 VTAIL.n132 VTAIL.n131 0.155672
R2091 VTAIL.n132 VTAIL.n89 0.155672
R2092 VTAIL.n139 VTAIL.n89 0.155672
R2093 VTAIL.n140 VTAIL.n139 0.155672
R2094 VTAIL.n140 VTAIL.n85 0.155672
R2095 VTAIL.n147 VTAIL.n85 0.155672
R2096 VTAIL.n148 VTAIL.n147 0.155672
R2097 VTAIL.n148 VTAIL.n81 0.155672
R2098 VTAIL.n155 VTAIL.n81 0.155672
R2099 VTAIL.n186 VTAIL.n181 0.155672
R2100 VTAIL.n193 VTAIL.n181 0.155672
R2101 VTAIL.n194 VTAIL.n193 0.155672
R2102 VTAIL.n194 VTAIL.n177 0.155672
R2103 VTAIL.n201 VTAIL.n177 0.155672
R2104 VTAIL.n202 VTAIL.n201 0.155672
R2105 VTAIL.n202 VTAIL.n173 0.155672
R2106 VTAIL.n211 VTAIL.n173 0.155672
R2107 VTAIL.n212 VTAIL.n211 0.155672
R2108 VTAIL.n212 VTAIL.n169 0.155672
R2109 VTAIL.n219 VTAIL.n169 0.155672
R2110 VTAIL.n220 VTAIL.n219 0.155672
R2111 VTAIL.n220 VTAIL.n165 0.155672
R2112 VTAIL.n227 VTAIL.n165 0.155672
R2113 VTAIL.n228 VTAIL.n227 0.155672
R2114 VTAIL.n228 VTAIL.n161 0.155672
R2115 VTAIL.n235 VTAIL.n161 0.155672
R2116 VTAIL.n551 VTAIL.n477 0.155672
R2117 VTAIL.n544 VTAIL.n477 0.155672
R2118 VTAIL.n544 VTAIL.n543 0.155672
R2119 VTAIL.n543 VTAIL.n481 0.155672
R2120 VTAIL.n536 VTAIL.n481 0.155672
R2121 VTAIL.n536 VTAIL.n535 0.155672
R2122 VTAIL.n535 VTAIL.n485 0.155672
R2123 VTAIL.n528 VTAIL.n485 0.155672
R2124 VTAIL.n528 VTAIL.n527 0.155672
R2125 VTAIL.n527 VTAIL.n489 0.155672
R2126 VTAIL.n519 VTAIL.n489 0.155672
R2127 VTAIL.n519 VTAIL.n518 0.155672
R2128 VTAIL.n518 VTAIL.n494 0.155672
R2129 VTAIL.n511 VTAIL.n494 0.155672
R2130 VTAIL.n511 VTAIL.n510 0.155672
R2131 VTAIL.n510 VTAIL.n498 0.155672
R2132 VTAIL.n503 VTAIL.n498 0.155672
R2133 VTAIL.n471 VTAIL.n397 0.155672
R2134 VTAIL.n464 VTAIL.n397 0.155672
R2135 VTAIL.n464 VTAIL.n463 0.155672
R2136 VTAIL.n463 VTAIL.n401 0.155672
R2137 VTAIL.n456 VTAIL.n401 0.155672
R2138 VTAIL.n456 VTAIL.n455 0.155672
R2139 VTAIL.n455 VTAIL.n405 0.155672
R2140 VTAIL.n448 VTAIL.n405 0.155672
R2141 VTAIL.n448 VTAIL.n447 0.155672
R2142 VTAIL.n447 VTAIL.n409 0.155672
R2143 VTAIL.n439 VTAIL.n409 0.155672
R2144 VTAIL.n439 VTAIL.n438 0.155672
R2145 VTAIL.n438 VTAIL.n414 0.155672
R2146 VTAIL.n431 VTAIL.n414 0.155672
R2147 VTAIL.n431 VTAIL.n430 0.155672
R2148 VTAIL.n430 VTAIL.n418 0.155672
R2149 VTAIL.n423 VTAIL.n418 0.155672
R2150 VTAIL.n393 VTAIL.n319 0.155672
R2151 VTAIL.n386 VTAIL.n319 0.155672
R2152 VTAIL.n386 VTAIL.n385 0.155672
R2153 VTAIL.n385 VTAIL.n323 0.155672
R2154 VTAIL.n378 VTAIL.n323 0.155672
R2155 VTAIL.n378 VTAIL.n377 0.155672
R2156 VTAIL.n377 VTAIL.n327 0.155672
R2157 VTAIL.n370 VTAIL.n327 0.155672
R2158 VTAIL.n370 VTAIL.n369 0.155672
R2159 VTAIL.n369 VTAIL.n331 0.155672
R2160 VTAIL.n361 VTAIL.n331 0.155672
R2161 VTAIL.n361 VTAIL.n360 0.155672
R2162 VTAIL.n360 VTAIL.n336 0.155672
R2163 VTAIL.n353 VTAIL.n336 0.155672
R2164 VTAIL.n353 VTAIL.n352 0.155672
R2165 VTAIL.n352 VTAIL.n340 0.155672
R2166 VTAIL.n345 VTAIL.n340 0.155672
R2167 VTAIL.n313 VTAIL.n239 0.155672
R2168 VTAIL.n306 VTAIL.n239 0.155672
R2169 VTAIL.n306 VTAIL.n305 0.155672
R2170 VTAIL.n305 VTAIL.n243 0.155672
R2171 VTAIL.n298 VTAIL.n243 0.155672
R2172 VTAIL.n298 VTAIL.n297 0.155672
R2173 VTAIL.n297 VTAIL.n247 0.155672
R2174 VTAIL.n290 VTAIL.n247 0.155672
R2175 VTAIL.n290 VTAIL.n289 0.155672
R2176 VTAIL.n289 VTAIL.n251 0.155672
R2177 VTAIL.n281 VTAIL.n251 0.155672
R2178 VTAIL.n281 VTAIL.n280 0.155672
R2179 VTAIL.n280 VTAIL.n256 0.155672
R2180 VTAIL.n273 VTAIL.n256 0.155672
R2181 VTAIL.n273 VTAIL.n272 0.155672
R2182 VTAIL.n272 VTAIL.n260 0.155672
R2183 VTAIL.n265 VTAIL.n260 0.155672
R2184 VTAIL VTAIL.n1 0.0586897
R2185 VN.n5 VN.t1 229.371
R2186 VN.n28 VN.t4 229.371
R2187 VN.n6 VN.t0 200.411
R2188 VN.n14 VN.t3 200.411
R2189 VN.n21 VN.t6 200.411
R2190 VN.n29 VN.t5 200.411
R2191 VN.n37 VN.t7 200.411
R2192 VN.n44 VN.t2 200.411
R2193 VN.n22 VN.n21 182.722
R2194 VN.n45 VN.n44 182.722
R2195 VN.n43 VN.n23 161.3
R2196 VN.n42 VN.n41 161.3
R2197 VN.n40 VN.n24 161.3
R2198 VN.n39 VN.n38 161.3
R2199 VN.n36 VN.n25 161.3
R2200 VN.n35 VN.n34 161.3
R2201 VN.n33 VN.n26 161.3
R2202 VN.n32 VN.n31 161.3
R2203 VN.n30 VN.n27 161.3
R2204 VN.n20 VN.n0 161.3
R2205 VN.n19 VN.n18 161.3
R2206 VN.n17 VN.n1 161.3
R2207 VN.n16 VN.n15 161.3
R2208 VN.n13 VN.n2 161.3
R2209 VN.n12 VN.n11 161.3
R2210 VN.n10 VN.n3 161.3
R2211 VN.n9 VN.n8 161.3
R2212 VN.n7 VN.n4 161.3
R2213 VN.n6 VN.n5 67.3788
R2214 VN.n29 VN.n28 67.3788
R2215 VN VN.n45 48.6615
R2216 VN.n19 VN.n1 44.3055
R2217 VN.n42 VN.n24 44.3055
R2218 VN.n8 VN.n3 40.4106
R2219 VN.n12 VN.n3 40.4106
R2220 VN.n31 VN.n26 40.4106
R2221 VN.n35 VN.n26 40.4106
R2222 VN.n15 VN.n1 36.5157
R2223 VN.n38 VN.n24 36.5157
R2224 VN.n8 VN.n7 24.3439
R2225 VN.n13 VN.n12 24.3439
R2226 VN.n20 VN.n19 24.3439
R2227 VN.n31 VN.n30 24.3439
R2228 VN.n36 VN.n35 24.3439
R2229 VN.n43 VN.n42 24.3439
R2230 VN.n15 VN.n14 23.3702
R2231 VN.n38 VN.n37 23.3702
R2232 VN.n28 VN.n27 18.7354
R2233 VN.n5 VN.n4 18.7354
R2234 VN.n21 VN.n20 2.92171
R2235 VN.n44 VN.n43 2.92171
R2236 VN.n7 VN.n6 0.974237
R2237 VN.n14 VN.n13 0.974237
R2238 VN.n30 VN.n29 0.974237
R2239 VN.n37 VN.n36 0.974237
R2240 VN.n45 VN.n23 0.189894
R2241 VN.n41 VN.n23 0.189894
R2242 VN.n41 VN.n40 0.189894
R2243 VN.n40 VN.n39 0.189894
R2244 VN.n39 VN.n25 0.189894
R2245 VN.n34 VN.n25 0.189894
R2246 VN.n34 VN.n33 0.189894
R2247 VN.n33 VN.n32 0.189894
R2248 VN.n32 VN.n27 0.189894
R2249 VN.n9 VN.n4 0.189894
R2250 VN.n10 VN.n9 0.189894
R2251 VN.n11 VN.n10 0.189894
R2252 VN.n11 VN.n2 0.189894
R2253 VN.n16 VN.n2 0.189894
R2254 VN.n17 VN.n16 0.189894
R2255 VN.n18 VN.n17 0.189894
R2256 VN.n18 VN.n0 0.189894
R2257 VN.n22 VN.n0 0.189894
R2258 VN VN.n22 0.0516364
R2259 VDD2.n2 VDD2.n1 71.2933
R2260 VDD2.n2 VDD2.n0 71.2933
R2261 VDD2 VDD2.n5 71.2905
R2262 VDD2.n4 VDD2.n3 70.4693
R2263 VDD2.n4 VDD2.n2 43.8877
R2264 VDD2.n5 VDD2.t2 2.28637
R2265 VDD2.n5 VDD2.t3 2.28637
R2266 VDD2.n3 VDD2.t5 2.28637
R2267 VDD2.n3 VDD2.t0 2.28637
R2268 VDD2.n1 VDD2.t4 2.28637
R2269 VDD2.n1 VDD2.t1 2.28637
R2270 VDD2.n0 VDD2.t6 2.28637
R2271 VDD2.n0 VDD2.t7 2.28637
R2272 VDD2 VDD2.n4 0.938
C0 VDD2 w_n3010_n3812# 1.79422f
C1 VTAIL w_n3010_n3812# 4.67371f
C2 VP VN 6.99104f
C3 VDD1 VDD2 1.31171f
C4 VTAIL VDD1 9.20996f
C5 VN w_n3010_n3812# 5.93482f
C6 VTAIL VDD2 9.25841f
C7 VN VDD1 0.149401f
C8 VN VDD2 9.251151f
C9 VN VTAIL 9.263339f
C10 B VP 1.687f
C11 B w_n3010_n3812# 9.37482f
C12 VP w_n3010_n3812# 6.32296f
C13 B VDD1 1.4385f
C14 B VDD2 1.50652f
C15 VP VDD1 9.52505f
C16 B VTAIL 5.21031f
C17 VP VDD2 0.424247f
C18 VP VTAIL 9.27744f
C19 VDD1 w_n3010_n3812# 1.71685f
C20 B VN 1.04109f
C21 VDD2 VSUBS 1.644096f
C22 VDD1 VSUBS 2.126377f
C23 VTAIL VSUBS 1.253682f
C24 VN VSUBS 5.73335f
C25 VP VSUBS 2.739221f
C26 B VSUBS 4.196338f
C27 w_n3010_n3812# VSUBS 0.140832p
C28 VDD2.t6 VSUBS 0.280057f
C29 VDD2.t7 VSUBS 0.280057f
C30 VDD2.n0 VSUBS 2.24817f
C31 VDD2.t4 VSUBS 0.280057f
C32 VDD2.t1 VSUBS 0.280057f
C33 VDD2.n1 VSUBS 2.24817f
C34 VDD2.n2 VSUBS 3.45115f
C35 VDD2.t5 VSUBS 0.280057f
C36 VDD2.t0 VSUBS 0.280057f
C37 VDD2.n3 VSUBS 2.24001f
C38 VDD2.n4 VSUBS 3.08541f
C39 VDD2.t2 VSUBS 0.280057f
C40 VDD2.t3 VSUBS 0.280057f
C41 VDD2.n5 VSUBS 2.24814f
C42 VN.n0 VSUBS 0.034941f
C43 VN.t6 VSUBS 2.32524f
C44 VN.n1 VSUBS 0.029005f
C45 VN.n2 VSUBS 0.034941f
C46 VN.t3 VSUBS 2.32524f
C47 VN.n3 VSUBS 0.028275f
C48 VN.n4 VSUBS 0.222879f
C49 VN.t0 VSUBS 2.32524f
C50 VN.t1 VSUBS 2.44833f
C51 VN.n5 VSUBS 0.92281f
C52 VN.n6 VSUBS 0.886498f
C53 VN.n7 VSUBS 0.034426f
C54 VN.n8 VSUBS 0.069816f
C55 VN.n9 VSUBS 0.034941f
C56 VN.n10 VSUBS 0.034941f
C57 VN.n11 VSUBS 0.034941f
C58 VN.n12 VSUBS 0.069816f
C59 VN.n13 VSUBS 0.034426f
C60 VN.n14 VSUBS 0.825999f
C61 VN.n15 VSUBS 0.06954f
C62 VN.n16 VSUBS 0.034941f
C63 VN.n17 VSUBS 0.034941f
C64 VN.n18 VSUBS 0.034941f
C65 VN.n19 VSUBS 0.068068f
C66 VN.n20 VSUBS 0.037011f
C67 VN.n21 VSUBS 0.899177f
C68 VN.n22 VSUBS 0.036796f
C69 VN.n23 VSUBS 0.034941f
C70 VN.t2 VSUBS 2.32524f
C71 VN.n24 VSUBS 0.029005f
C72 VN.n25 VSUBS 0.034941f
C73 VN.t7 VSUBS 2.32524f
C74 VN.n26 VSUBS 0.028275f
C75 VN.n27 VSUBS 0.222879f
C76 VN.t5 VSUBS 2.32524f
C77 VN.t4 VSUBS 2.44833f
C78 VN.n28 VSUBS 0.92281f
C79 VN.n29 VSUBS 0.886498f
C80 VN.n30 VSUBS 0.034426f
C81 VN.n31 VSUBS 0.069816f
C82 VN.n32 VSUBS 0.034941f
C83 VN.n33 VSUBS 0.034941f
C84 VN.n34 VSUBS 0.034941f
C85 VN.n35 VSUBS 0.069816f
C86 VN.n36 VSUBS 0.034426f
C87 VN.n37 VSUBS 0.825999f
C88 VN.n38 VSUBS 0.06954f
C89 VN.n39 VSUBS 0.034941f
C90 VN.n40 VSUBS 0.034941f
C91 VN.n41 VSUBS 0.034941f
C92 VN.n42 VSUBS 0.068068f
C93 VN.n43 VSUBS 0.037011f
C94 VN.n44 VSUBS 0.899177f
C95 VN.n45 VSUBS 1.83391f
C96 VTAIL.t1 VSUBS 0.2689f
C97 VTAIL.t5 VSUBS 0.2689f
C98 VTAIL.n0 VSUBS 2.00683f
C99 VTAIL.n1 VSUBS 0.720244f
C100 VTAIL.n2 VSUBS 0.026802f
C101 VTAIL.n3 VSUBS 0.02393f
C102 VTAIL.n4 VSUBS 0.012859f
C103 VTAIL.n5 VSUBS 0.030394f
C104 VTAIL.n6 VSUBS 0.013615f
C105 VTAIL.n7 VSUBS 0.02393f
C106 VTAIL.n8 VSUBS 0.012859f
C107 VTAIL.n9 VSUBS 0.030394f
C108 VTAIL.n10 VSUBS 0.013615f
C109 VTAIL.n11 VSUBS 0.02393f
C110 VTAIL.n12 VSUBS 0.012859f
C111 VTAIL.n13 VSUBS 0.030394f
C112 VTAIL.n14 VSUBS 0.013615f
C113 VTAIL.n15 VSUBS 0.02393f
C114 VTAIL.n16 VSUBS 0.013237f
C115 VTAIL.n17 VSUBS 0.030394f
C116 VTAIL.n18 VSUBS 0.013615f
C117 VTAIL.n19 VSUBS 0.02393f
C118 VTAIL.n20 VSUBS 0.012859f
C119 VTAIL.n21 VSUBS 0.030394f
C120 VTAIL.n22 VSUBS 0.013615f
C121 VTAIL.n23 VSUBS 0.02393f
C122 VTAIL.n24 VSUBS 0.012859f
C123 VTAIL.n25 VSUBS 0.022795f
C124 VTAIL.n26 VSUBS 0.022864f
C125 VTAIL.t6 VSUBS 0.065671f
C126 VTAIL.n27 VSUBS 0.212478f
C127 VTAIL.n28 VSUBS 1.40852f
C128 VTAIL.n29 VSUBS 0.012859f
C129 VTAIL.n30 VSUBS 0.013615f
C130 VTAIL.n31 VSUBS 0.030394f
C131 VTAIL.n32 VSUBS 0.030394f
C132 VTAIL.n33 VSUBS 0.013615f
C133 VTAIL.n34 VSUBS 0.012859f
C134 VTAIL.n35 VSUBS 0.02393f
C135 VTAIL.n36 VSUBS 0.02393f
C136 VTAIL.n37 VSUBS 0.012859f
C137 VTAIL.n38 VSUBS 0.013615f
C138 VTAIL.n39 VSUBS 0.030394f
C139 VTAIL.n40 VSUBS 0.030394f
C140 VTAIL.n41 VSUBS 0.013615f
C141 VTAIL.n42 VSUBS 0.012859f
C142 VTAIL.n43 VSUBS 0.02393f
C143 VTAIL.n44 VSUBS 0.02393f
C144 VTAIL.n45 VSUBS 0.012859f
C145 VTAIL.n46 VSUBS 0.012859f
C146 VTAIL.n47 VSUBS 0.013615f
C147 VTAIL.n48 VSUBS 0.030394f
C148 VTAIL.n49 VSUBS 0.030394f
C149 VTAIL.n50 VSUBS 0.030394f
C150 VTAIL.n51 VSUBS 0.013237f
C151 VTAIL.n52 VSUBS 0.012859f
C152 VTAIL.n53 VSUBS 0.02393f
C153 VTAIL.n54 VSUBS 0.02393f
C154 VTAIL.n55 VSUBS 0.012859f
C155 VTAIL.n56 VSUBS 0.013615f
C156 VTAIL.n57 VSUBS 0.030394f
C157 VTAIL.n58 VSUBS 0.030394f
C158 VTAIL.n59 VSUBS 0.013615f
C159 VTAIL.n60 VSUBS 0.012859f
C160 VTAIL.n61 VSUBS 0.02393f
C161 VTAIL.n62 VSUBS 0.02393f
C162 VTAIL.n63 VSUBS 0.012859f
C163 VTAIL.n64 VSUBS 0.013615f
C164 VTAIL.n65 VSUBS 0.030394f
C165 VTAIL.n66 VSUBS 0.030394f
C166 VTAIL.n67 VSUBS 0.013615f
C167 VTAIL.n68 VSUBS 0.012859f
C168 VTAIL.n69 VSUBS 0.02393f
C169 VTAIL.n70 VSUBS 0.02393f
C170 VTAIL.n71 VSUBS 0.012859f
C171 VTAIL.n72 VSUBS 0.013615f
C172 VTAIL.n73 VSUBS 0.030394f
C173 VTAIL.n74 VSUBS 0.075312f
C174 VTAIL.n75 VSUBS 0.013615f
C175 VTAIL.n76 VSUBS 0.012859f
C176 VTAIL.n77 VSUBS 0.053351f
C177 VTAIL.n78 VSUBS 0.037889f
C178 VTAIL.n79 VSUBS 0.19116f
C179 VTAIL.n80 VSUBS 0.026802f
C180 VTAIL.n81 VSUBS 0.02393f
C181 VTAIL.n82 VSUBS 0.012859f
C182 VTAIL.n83 VSUBS 0.030394f
C183 VTAIL.n84 VSUBS 0.013615f
C184 VTAIL.n85 VSUBS 0.02393f
C185 VTAIL.n86 VSUBS 0.012859f
C186 VTAIL.n87 VSUBS 0.030394f
C187 VTAIL.n88 VSUBS 0.013615f
C188 VTAIL.n89 VSUBS 0.02393f
C189 VTAIL.n90 VSUBS 0.012859f
C190 VTAIL.n91 VSUBS 0.030394f
C191 VTAIL.n92 VSUBS 0.013615f
C192 VTAIL.n93 VSUBS 0.02393f
C193 VTAIL.n94 VSUBS 0.013237f
C194 VTAIL.n95 VSUBS 0.030394f
C195 VTAIL.n96 VSUBS 0.013615f
C196 VTAIL.n97 VSUBS 0.02393f
C197 VTAIL.n98 VSUBS 0.012859f
C198 VTAIL.n99 VSUBS 0.030394f
C199 VTAIL.n100 VSUBS 0.013615f
C200 VTAIL.n101 VSUBS 0.02393f
C201 VTAIL.n102 VSUBS 0.012859f
C202 VTAIL.n103 VSUBS 0.022795f
C203 VTAIL.n104 VSUBS 0.022864f
C204 VTAIL.t12 VSUBS 0.065671f
C205 VTAIL.n105 VSUBS 0.212478f
C206 VTAIL.n106 VSUBS 1.40852f
C207 VTAIL.n107 VSUBS 0.012859f
C208 VTAIL.n108 VSUBS 0.013615f
C209 VTAIL.n109 VSUBS 0.030394f
C210 VTAIL.n110 VSUBS 0.030394f
C211 VTAIL.n111 VSUBS 0.013615f
C212 VTAIL.n112 VSUBS 0.012859f
C213 VTAIL.n113 VSUBS 0.02393f
C214 VTAIL.n114 VSUBS 0.02393f
C215 VTAIL.n115 VSUBS 0.012859f
C216 VTAIL.n116 VSUBS 0.013615f
C217 VTAIL.n117 VSUBS 0.030394f
C218 VTAIL.n118 VSUBS 0.030394f
C219 VTAIL.n119 VSUBS 0.013615f
C220 VTAIL.n120 VSUBS 0.012859f
C221 VTAIL.n121 VSUBS 0.02393f
C222 VTAIL.n122 VSUBS 0.02393f
C223 VTAIL.n123 VSUBS 0.012859f
C224 VTAIL.n124 VSUBS 0.012859f
C225 VTAIL.n125 VSUBS 0.013615f
C226 VTAIL.n126 VSUBS 0.030394f
C227 VTAIL.n127 VSUBS 0.030394f
C228 VTAIL.n128 VSUBS 0.030394f
C229 VTAIL.n129 VSUBS 0.013237f
C230 VTAIL.n130 VSUBS 0.012859f
C231 VTAIL.n131 VSUBS 0.02393f
C232 VTAIL.n132 VSUBS 0.02393f
C233 VTAIL.n133 VSUBS 0.012859f
C234 VTAIL.n134 VSUBS 0.013615f
C235 VTAIL.n135 VSUBS 0.030394f
C236 VTAIL.n136 VSUBS 0.030394f
C237 VTAIL.n137 VSUBS 0.013615f
C238 VTAIL.n138 VSUBS 0.012859f
C239 VTAIL.n139 VSUBS 0.02393f
C240 VTAIL.n140 VSUBS 0.02393f
C241 VTAIL.n141 VSUBS 0.012859f
C242 VTAIL.n142 VSUBS 0.013615f
C243 VTAIL.n143 VSUBS 0.030394f
C244 VTAIL.n144 VSUBS 0.030394f
C245 VTAIL.n145 VSUBS 0.013615f
C246 VTAIL.n146 VSUBS 0.012859f
C247 VTAIL.n147 VSUBS 0.02393f
C248 VTAIL.n148 VSUBS 0.02393f
C249 VTAIL.n149 VSUBS 0.012859f
C250 VTAIL.n150 VSUBS 0.013615f
C251 VTAIL.n151 VSUBS 0.030394f
C252 VTAIL.n152 VSUBS 0.075312f
C253 VTAIL.n153 VSUBS 0.013615f
C254 VTAIL.n154 VSUBS 0.012859f
C255 VTAIL.n155 VSUBS 0.053351f
C256 VTAIL.n156 VSUBS 0.037889f
C257 VTAIL.n157 VSUBS 0.19116f
C258 VTAIL.t8 VSUBS 0.2689f
C259 VTAIL.t11 VSUBS 0.2689f
C260 VTAIL.n158 VSUBS 2.00683f
C261 VTAIL.n159 VSUBS 0.851359f
C262 VTAIL.n160 VSUBS 0.026802f
C263 VTAIL.n161 VSUBS 0.02393f
C264 VTAIL.n162 VSUBS 0.012859f
C265 VTAIL.n163 VSUBS 0.030394f
C266 VTAIL.n164 VSUBS 0.013615f
C267 VTAIL.n165 VSUBS 0.02393f
C268 VTAIL.n166 VSUBS 0.012859f
C269 VTAIL.n167 VSUBS 0.030394f
C270 VTAIL.n168 VSUBS 0.013615f
C271 VTAIL.n169 VSUBS 0.02393f
C272 VTAIL.n170 VSUBS 0.012859f
C273 VTAIL.n171 VSUBS 0.030394f
C274 VTAIL.n172 VSUBS 0.013615f
C275 VTAIL.n173 VSUBS 0.02393f
C276 VTAIL.n174 VSUBS 0.013237f
C277 VTAIL.n175 VSUBS 0.030394f
C278 VTAIL.n176 VSUBS 0.013615f
C279 VTAIL.n177 VSUBS 0.02393f
C280 VTAIL.n178 VSUBS 0.012859f
C281 VTAIL.n179 VSUBS 0.030394f
C282 VTAIL.n180 VSUBS 0.013615f
C283 VTAIL.n181 VSUBS 0.02393f
C284 VTAIL.n182 VSUBS 0.012859f
C285 VTAIL.n183 VSUBS 0.022795f
C286 VTAIL.n184 VSUBS 0.022864f
C287 VTAIL.t10 VSUBS 0.065671f
C288 VTAIL.n185 VSUBS 0.212478f
C289 VTAIL.n186 VSUBS 1.40852f
C290 VTAIL.n187 VSUBS 0.012859f
C291 VTAIL.n188 VSUBS 0.013615f
C292 VTAIL.n189 VSUBS 0.030394f
C293 VTAIL.n190 VSUBS 0.030394f
C294 VTAIL.n191 VSUBS 0.013615f
C295 VTAIL.n192 VSUBS 0.012859f
C296 VTAIL.n193 VSUBS 0.02393f
C297 VTAIL.n194 VSUBS 0.02393f
C298 VTAIL.n195 VSUBS 0.012859f
C299 VTAIL.n196 VSUBS 0.013615f
C300 VTAIL.n197 VSUBS 0.030394f
C301 VTAIL.n198 VSUBS 0.030394f
C302 VTAIL.n199 VSUBS 0.013615f
C303 VTAIL.n200 VSUBS 0.012859f
C304 VTAIL.n201 VSUBS 0.02393f
C305 VTAIL.n202 VSUBS 0.02393f
C306 VTAIL.n203 VSUBS 0.012859f
C307 VTAIL.n204 VSUBS 0.012859f
C308 VTAIL.n205 VSUBS 0.013615f
C309 VTAIL.n206 VSUBS 0.030394f
C310 VTAIL.n207 VSUBS 0.030394f
C311 VTAIL.n208 VSUBS 0.030394f
C312 VTAIL.n209 VSUBS 0.013237f
C313 VTAIL.n210 VSUBS 0.012859f
C314 VTAIL.n211 VSUBS 0.02393f
C315 VTAIL.n212 VSUBS 0.02393f
C316 VTAIL.n213 VSUBS 0.012859f
C317 VTAIL.n214 VSUBS 0.013615f
C318 VTAIL.n215 VSUBS 0.030394f
C319 VTAIL.n216 VSUBS 0.030394f
C320 VTAIL.n217 VSUBS 0.013615f
C321 VTAIL.n218 VSUBS 0.012859f
C322 VTAIL.n219 VSUBS 0.02393f
C323 VTAIL.n220 VSUBS 0.02393f
C324 VTAIL.n221 VSUBS 0.012859f
C325 VTAIL.n222 VSUBS 0.013615f
C326 VTAIL.n223 VSUBS 0.030394f
C327 VTAIL.n224 VSUBS 0.030394f
C328 VTAIL.n225 VSUBS 0.013615f
C329 VTAIL.n226 VSUBS 0.012859f
C330 VTAIL.n227 VSUBS 0.02393f
C331 VTAIL.n228 VSUBS 0.02393f
C332 VTAIL.n229 VSUBS 0.012859f
C333 VTAIL.n230 VSUBS 0.013615f
C334 VTAIL.n231 VSUBS 0.030394f
C335 VTAIL.n232 VSUBS 0.075312f
C336 VTAIL.n233 VSUBS 0.013615f
C337 VTAIL.n234 VSUBS 0.012859f
C338 VTAIL.n235 VSUBS 0.053351f
C339 VTAIL.n236 VSUBS 0.037889f
C340 VTAIL.n237 VSUBS 1.56081f
C341 VTAIL.n238 VSUBS 0.026802f
C342 VTAIL.n239 VSUBS 0.02393f
C343 VTAIL.n240 VSUBS 0.012859f
C344 VTAIL.n241 VSUBS 0.030394f
C345 VTAIL.n242 VSUBS 0.013615f
C346 VTAIL.n243 VSUBS 0.02393f
C347 VTAIL.n244 VSUBS 0.012859f
C348 VTAIL.n245 VSUBS 0.030394f
C349 VTAIL.n246 VSUBS 0.013615f
C350 VTAIL.n247 VSUBS 0.02393f
C351 VTAIL.n248 VSUBS 0.012859f
C352 VTAIL.n249 VSUBS 0.030394f
C353 VTAIL.n250 VSUBS 0.013615f
C354 VTAIL.n251 VSUBS 0.02393f
C355 VTAIL.n252 VSUBS 0.013237f
C356 VTAIL.n253 VSUBS 0.030394f
C357 VTAIL.n254 VSUBS 0.012859f
C358 VTAIL.n255 VSUBS 0.013615f
C359 VTAIL.n256 VSUBS 0.02393f
C360 VTAIL.n257 VSUBS 0.012859f
C361 VTAIL.n258 VSUBS 0.030394f
C362 VTAIL.n259 VSUBS 0.013615f
C363 VTAIL.n260 VSUBS 0.02393f
C364 VTAIL.n261 VSUBS 0.012859f
C365 VTAIL.n262 VSUBS 0.022795f
C366 VTAIL.n263 VSUBS 0.022864f
C367 VTAIL.t4 VSUBS 0.065671f
C368 VTAIL.n264 VSUBS 0.212478f
C369 VTAIL.n265 VSUBS 1.40852f
C370 VTAIL.n266 VSUBS 0.012859f
C371 VTAIL.n267 VSUBS 0.013615f
C372 VTAIL.n268 VSUBS 0.030394f
C373 VTAIL.n269 VSUBS 0.030394f
C374 VTAIL.n270 VSUBS 0.013615f
C375 VTAIL.n271 VSUBS 0.012859f
C376 VTAIL.n272 VSUBS 0.02393f
C377 VTAIL.n273 VSUBS 0.02393f
C378 VTAIL.n274 VSUBS 0.012859f
C379 VTAIL.n275 VSUBS 0.013615f
C380 VTAIL.n276 VSUBS 0.030394f
C381 VTAIL.n277 VSUBS 0.030394f
C382 VTAIL.n278 VSUBS 0.013615f
C383 VTAIL.n279 VSUBS 0.012859f
C384 VTAIL.n280 VSUBS 0.02393f
C385 VTAIL.n281 VSUBS 0.02393f
C386 VTAIL.n282 VSUBS 0.012859f
C387 VTAIL.n283 VSUBS 0.013615f
C388 VTAIL.n284 VSUBS 0.030394f
C389 VTAIL.n285 VSUBS 0.030394f
C390 VTAIL.n286 VSUBS 0.030394f
C391 VTAIL.n287 VSUBS 0.013237f
C392 VTAIL.n288 VSUBS 0.012859f
C393 VTAIL.n289 VSUBS 0.02393f
C394 VTAIL.n290 VSUBS 0.02393f
C395 VTAIL.n291 VSUBS 0.012859f
C396 VTAIL.n292 VSUBS 0.013615f
C397 VTAIL.n293 VSUBS 0.030394f
C398 VTAIL.n294 VSUBS 0.030394f
C399 VTAIL.n295 VSUBS 0.013615f
C400 VTAIL.n296 VSUBS 0.012859f
C401 VTAIL.n297 VSUBS 0.02393f
C402 VTAIL.n298 VSUBS 0.02393f
C403 VTAIL.n299 VSUBS 0.012859f
C404 VTAIL.n300 VSUBS 0.013615f
C405 VTAIL.n301 VSUBS 0.030394f
C406 VTAIL.n302 VSUBS 0.030394f
C407 VTAIL.n303 VSUBS 0.013615f
C408 VTAIL.n304 VSUBS 0.012859f
C409 VTAIL.n305 VSUBS 0.02393f
C410 VTAIL.n306 VSUBS 0.02393f
C411 VTAIL.n307 VSUBS 0.012859f
C412 VTAIL.n308 VSUBS 0.013615f
C413 VTAIL.n309 VSUBS 0.030394f
C414 VTAIL.n310 VSUBS 0.075312f
C415 VTAIL.n311 VSUBS 0.013615f
C416 VTAIL.n312 VSUBS 0.012859f
C417 VTAIL.n313 VSUBS 0.053351f
C418 VTAIL.n314 VSUBS 0.037889f
C419 VTAIL.n315 VSUBS 1.56081f
C420 VTAIL.t0 VSUBS 0.2689f
C421 VTAIL.t15 VSUBS 0.2689f
C422 VTAIL.n316 VSUBS 2.00684f
C423 VTAIL.n317 VSUBS 0.851349f
C424 VTAIL.n318 VSUBS 0.026802f
C425 VTAIL.n319 VSUBS 0.02393f
C426 VTAIL.n320 VSUBS 0.012859f
C427 VTAIL.n321 VSUBS 0.030394f
C428 VTAIL.n322 VSUBS 0.013615f
C429 VTAIL.n323 VSUBS 0.02393f
C430 VTAIL.n324 VSUBS 0.012859f
C431 VTAIL.n325 VSUBS 0.030394f
C432 VTAIL.n326 VSUBS 0.013615f
C433 VTAIL.n327 VSUBS 0.02393f
C434 VTAIL.n328 VSUBS 0.012859f
C435 VTAIL.n329 VSUBS 0.030394f
C436 VTAIL.n330 VSUBS 0.013615f
C437 VTAIL.n331 VSUBS 0.02393f
C438 VTAIL.n332 VSUBS 0.013237f
C439 VTAIL.n333 VSUBS 0.030394f
C440 VTAIL.n334 VSUBS 0.012859f
C441 VTAIL.n335 VSUBS 0.013615f
C442 VTAIL.n336 VSUBS 0.02393f
C443 VTAIL.n337 VSUBS 0.012859f
C444 VTAIL.n338 VSUBS 0.030394f
C445 VTAIL.n339 VSUBS 0.013615f
C446 VTAIL.n340 VSUBS 0.02393f
C447 VTAIL.n341 VSUBS 0.012859f
C448 VTAIL.n342 VSUBS 0.022795f
C449 VTAIL.n343 VSUBS 0.022864f
C450 VTAIL.t3 VSUBS 0.065671f
C451 VTAIL.n344 VSUBS 0.212478f
C452 VTAIL.n345 VSUBS 1.40852f
C453 VTAIL.n346 VSUBS 0.012859f
C454 VTAIL.n347 VSUBS 0.013615f
C455 VTAIL.n348 VSUBS 0.030394f
C456 VTAIL.n349 VSUBS 0.030394f
C457 VTAIL.n350 VSUBS 0.013615f
C458 VTAIL.n351 VSUBS 0.012859f
C459 VTAIL.n352 VSUBS 0.02393f
C460 VTAIL.n353 VSUBS 0.02393f
C461 VTAIL.n354 VSUBS 0.012859f
C462 VTAIL.n355 VSUBS 0.013615f
C463 VTAIL.n356 VSUBS 0.030394f
C464 VTAIL.n357 VSUBS 0.030394f
C465 VTAIL.n358 VSUBS 0.013615f
C466 VTAIL.n359 VSUBS 0.012859f
C467 VTAIL.n360 VSUBS 0.02393f
C468 VTAIL.n361 VSUBS 0.02393f
C469 VTAIL.n362 VSUBS 0.012859f
C470 VTAIL.n363 VSUBS 0.013615f
C471 VTAIL.n364 VSUBS 0.030394f
C472 VTAIL.n365 VSUBS 0.030394f
C473 VTAIL.n366 VSUBS 0.030394f
C474 VTAIL.n367 VSUBS 0.013237f
C475 VTAIL.n368 VSUBS 0.012859f
C476 VTAIL.n369 VSUBS 0.02393f
C477 VTAIL.n370 VSUBS 0.02393f
C478 VTAIL.n371 VSUBS 0.012859f
C479 VTAIL.n372 VSUBS 0.013615f
C480 VTAIL.n373 VSUBS 0.030394f
C481 VTAIL.n374 VSUBS 0.030394f
C482 VTAIL.n375 VSUBS 0.013615f
C483 VTAIL.n376 VSUBS 0.012859f
C484 VTAIL.n377 VSUBS 0.02393f
C485 VTAIL.n378 VSUBS 0.02393f
C486 VTAIL.n379 VSUBS 0.012859f
C487 VTAIL.n380 VSUBS 0.013615f
C488 VTAIL.n381 VSUBS 0.030394f
C489 VTAIL.n382 VSUBS 0.030394f
C490 VTAIL.n383 VSUBS 0.013615f
C491 VTAIL.n384 VSUBS 0.012859f
C492 VTAIL.n385 VSUBS 0.02393f
C493 VTAIL.n386 VSUBS 0.02393f
C494 VTAIL.n387 VSUBS 0.012859f
C495 VTAIL.n388 VSUBS 0.013615f
C496 VTAIL.n389 VSUBS 0.030394f
C497 VTAIL.n390 VSUBS 0.075312f
C498 VTAIL.n391 VSUBS 0.013615f
C499 VTAIL.n392 VSUBS 0.012859f
C500 VTAIL.n393 VSUBS 0.053351f
C501 VTAIL.n394 VSUBS 0.037889f
C502 VTAIL.n395 VSUBS 0.19116f
C503 VTAIL.n396 VSUBS 0.026802f
C504 VTAIL.n397 VSUBS 0.02393f
C505 VTAIL.n398 VSUBS 0.012859f
C506 VTAIL.n399 VSUBS 0.030394f
C507 VTAIL.n400 VSUBS 0.013615f
C508 VTAIL.n401 VSUBS 0.02393f
C509 VTAIL.n402 VSUBS 0.012859f
C510 VTAIL.n403 VSUBS 0.030394f
C511 VTAIL.n404 VSUBS 0.013615f
C512 VTAIL.n405 VSUBS 0.02393f
C513 VTAIL.n406 VSUBS 0.012859f
C514 VTAIL.n407 VSUBS 0.030394f
C515 VTAIL.n408 VSUBS 0.013615f
C516 VTAIL.n409 VSUBS 0.02393f
C517 VTAIL.n410 VSUBS 0.013237f
C518 VTAIL.n411 VSUBS 0.030394f
C519 VTAIL.n412 VSUBS 0.012859f
C520 VTAIL.n413 VSUBS 0.013615f
C521 VTAIL.n414 VSUBS 0.02393f
C522 VTAIL.n415 VSUBS 0.012859f
C523 VTAIL.n416 VSUBS 0.030394f
C524 VTAIL.n417 VSUBS 0.013615f
C525 VTAIL.n418 VSUBS 0.02393f
C526 VTAIL.n419 VSUBS 0.012859f
C527 VTAIL.n420 VSUBS 0.022795f
C528 VTAIL.n421 VSUBS 0.022864f
C529 VTAIL.t9 VSUBS 0.065671f
C530 VTAIL.n422 VSUBS 0.212478f
C531 VTAIL.n423 VSUBS 1.40852f
C532 VTAIL.n424 VSUBS 0.012859f
C533 VTAIL.n425 VSUBS 0.013615f
C534 VTAIL.n426 VSUBS 0.030394f
C535 VTAIL.n427 VSUBS 0.030394f
C536 VTAIL.n428 VSUBS 0.013615f
C537 VTAIL.n429 VSUBS 0.012859f
C538 VTAIL.n430 VSUBS 0.02393f
C539 VTAIL.n431 VSUBS 0.02393f
C540 VTAIL.n432 VSUBS 0.012859f
C541 VTAIL.n433 VSUBS 0.013615f
C542 VTAIL.n434 VSUBS 0.030394f
C543 VTAIL.n435 VSUBS 0.030394f
C544 VTAIL.n436 VSUBS 0.013615f
C545 VTAIL.n437 VSUBS 0.012859f
C546 VTAIL.n438 VSUBS 0.02393f
C547 VTAIL.n439 VSUBS 0.02393f
C548 VTAIL.n440 VSUBS 0.012859f
C549 VTAIL.n441 VSUBS 0.013615f
C550 VTAIL.n442 VSUBS 0.030394f
C551 VTAIL.n443 VSUBS 0.030394f
C552 VTAIL.n444 VSUBS 0.030394f
C553 VTAIL.n445 VSUBS 0.013237f
C554 VTAIL.n446 VSUBS 0.012859f
C555 VTAIL.n447 VSUBS 0.02393f
C556 VTAIL.n448 VSUBS 0.02393f
C557 VTAIL.n449 VSUBS 0.012859f
C558 VTAIL.n450 VSUBS 0.013615f
C559 VTAIL.n451 VSUBS 0.030394f
C560 VTAIL.n452 VSUBS 0.030394f
C561 VTAIL.n453 VSUBS 0.013615f
C562 VTAIL.n454 VSUBS 0.012859f
C563 VTAIL.n455 VSUBS 0.02393f
C564 VTAIL.n456 VSUBS 0.02393f
C565 VTAIL.n457 VSUBS 0.012859f
C566 VTAIL.n458 VSUBS 0.013615f
C567 VTAIL.n459 VSUBS 0.030394f
C568 VTAIL.n460 VSUBS 0.030394f
C569 VTAIL.n461 VSUBS 0.013615f
C570 VTAIL.n462 VSUBS 0.012859f
C571 VTAIL.n463 VSUBS 0.02393f
C572 VTAIL.n464 VSUBS 0.02393f
C573 VTAIL.n465 VSUBS 0.012859f
C574 VTAIL.n466 VSUBS 0.013615f
C575 VTAIL.n467 VSUBS 0.030394f
C576 VTAIL.n468 VSUBS 0.075312f
C577 VTAIL.n469 VSUBS 0.013615f
C578 VTAIL.n470 VSUBS 0.012859f
C579 VTAIL.n471 VSUBS 0.053351f
C580 VTAIL.n472 VSUBS 0.037889f
C581 VTAIL.n473 VSUBS 0.19116f
C582 VTAIL.t7 VSUBS 0.2689f
C583 VTAIL.t14 VSUBS 0.2689f
C584 VTAIL.n474 VSUBS 2.00684f
C585 VTAIL.n475 VSUBS 0.851349f
C586 VTAIL.n476 VSUBS 0.026802f
C587 VTAIL.n477 VSUBS 0.02393f
C588 VTAIL.n478 VSUBS 0.012859f
C589 VTAIL.n479 VSUBS 0.030394f
C590 VTAIL.n480 VSUBS 0.013615f
C591 VTAIL.n481 VSUBS 0.02393f
C592 VTAIL.n482 VSUBS 0.012859f
C593 VTAIL.n483 VSUBS 0.030394f
C594 VTAIL.n484 VSUBS 0.013615f
C595 VTAIL.n485 VSUBS 0.02393f
C596 VTAIL.n486 VSUBS 0.012859f
C597 VTAIL.n487 VSUBS 0.030394f
C598 VTAIL.n488 VSUBS 0.013615f
C599 VTAIL.n489 VSUBS 0.02393f
C600 VTAIL.n490 VSUBS 0.013237f
C601 VTAIL.n491 VSUBS 0.030394f
C602 VTAIL.n492 VSUBS 0.012859f
C603 VTAIL.n493 VSUBS 0.013615f
C604 VTAIL.n494 VSUBS 0.02393f
C605 VTAIL.n495 VSUBS 0.012859f
C606 VTAIL.n496 VSUBS 0.030394f
C607 VTAIL.n497 VSUBS 0.013615f
C608 VTAIL.n498 VSUBS 0.02393f
C609 VTAIL.n499 VSUBS 0.012859f
C610 VTAIL.n500 VSUBS 0.022795f
C611 VTAIL.n501 VSUBS 0.022864f
C612 VTAIL.t13 VSUBS 0.065671f
C613 VTAIL.n502 VSUBS 0.212478f
C614 VTAIL.n503 VSUBS 1.40852f
C615 VTAIL.n504 VSUBS 0.012859f
C616 VTAIL.n505 VSUBS 0.013615f
C617 VTAIL.n506 VSUBS 0.030394f
C618 VTAIL.n507 VSUBS 0.030394f
C619 VTAIL.n508 VSUBS 0.013615f
C620 VTAIL.n509 VSUBS 0.012859f
C621 VTAIL.n510 VSUBS 0.02393f
C622 VTAIL.n511 VSUBS 0.02393f
C623 VTAIL.n512 VSUBS 0.012859f
C624 VTAIL.n513 VSUBS 0.013615f
C625 VTAIL.n514 VSUBS 0.030394f
C626 VTAIL.n515 VSUBS 0.030394f
C627 VTAIL.n516 VSUBS 0.013615f
C628 VTAIL.n517 VSUBS 0.012859f
C629 VTAIL.n518 VSUBS 0.02393f
C630 VTAIL.n519 VSUBS 0.02393f
C631 VTAIL.n520 VSUBS 0.012859f
C632 VTAIL.n521 VSUBS 0.013615f
C633 VTAIL.n522 VSUBS 0.030394f
C634 VTAIL.n523 VSUBS 0.030394f
C635 VTAIL.n524 VSUBS 0.030394f
C636 VTAIL.n525 VSUBS 0.013237f
C637 VTAIL.n526 VSUBS 0.012859f
C638 VTAIL.n527 VSUBS 0.02393f
C639 VTAIL.n528 VSUBS 0.02393f
C640 VTAIL.n529 VSUBS 0.012859f
C641 VTAIL.n530 VSUBS 0.013615f
C642 VTAIL.n531 VSUBS 0.030394f
C643 VTAIL.n532 VSUBS 0.030394f
C644 VTAIL.n533 VSUBS 0.013615f
C645 VTAIL.n534 VSUBS 0.012859f
C646 VTAIL.n535 VSUBS 0.02393f
C647 VTAIL.n536 VSUBS 0.02393f
C648 VTAIL.n537 VSUBS 0.012859f
C649 VTAIL.n538 VSUBS 0.013615f
C650 VTAIL.n539 VSUBS 0.030394f
C651 VTAIL.n540 VSUBS 0.030394f
C652 VTAIL.n541 VSUBS 0.013615f
C653 VTAIL.n542 VSUBS 0.012859f
C654 VTAIL.n543 VSUBS 0.02393f
C655 VTAIL.n544 VSUBS 0.02393f
C656 VTAIL.n545 VSUBS 0.012859f
C657 VTAIL.n546 VSUBS 0.013615f
C658 VTAIL.n547 VSUBS 0.030394f
C659 VTAIL.n548 VSUBS 0.075312f
C660 VTAIL.n549 VSUBS 0.013615f
C661 VTAIL.n550 VSUBS 0.012859f
C662 VTAIL.n551 VSUBS 0.053351f
C663 VTAIL.n552 VSUBS 0.037889f
C664 VTAIL.n553 VSUBS 1.56081f
C665 VTAIL.n554 VSUBS 0.026802f
C666 VTAIL.n555 VSUBS 0.02393f
C667 VTAIL.n556 VSUBS 0.012859f
C668 VTAIL.n557 VSUBS 0.030394f
C669 VTAIL.n558 VSUBS 0.013615f
C670 VTAIL.n559 VSUBS 0.02393f
C671 VTAIL.n560 VSUBS 0.012859f
C672 VTAIL.n561 VSUBS 0.030394f
C673 VTAIL.n562 VSUBS 0.013615f
C674 VTAIL.n563 VSUBS 0.02393f
C675 VTAIL.n564 VSUBS 0.012859f
C676 VTAIL.n565 VSUBS 0.030394f
C677 VTAIL.n566 VSUBS 0.013615f
C678 VTAIL.n567 VSUBS 0.02393f
C679 VTAIL.n568 VSUBS 0.013237f
C680 VTAIL.n569 VSUBS 0.030394f
C681 VTAIL.n570 VSUBS 0.013615f
C682 VTAIL.n571 VSUBS 0.02393f
C683 VTAIL.n572 VSUBS 0.012859f
C684 VTAIL.n573 VSUBS 0.030394f
C685 VTAIL.n574 VSUBS 0.013615f
C686 VTAIL.n575 VSUBS 0.02393f
C687 VTAIL.n576 VSUBS 0.012859f
C688 VTAIL.n577 VSUBS 0.022795f
C689 VTAIL.n578 VSUBS 0.022864f
C690 VTAIL.t2 VSUBS 0.065671f
C691 VTAIL.n579 VSUBS 0.212478f
C692 VTAIL.n580 VSUBS 1.40852f
C693 VTAIL.n581 VSUBS 0.012859f
C694 VTAIL.n582 VSUBS 0.013615f
C695 VTAIL.n583 VSUBS 0.030394f
C696 VTAIL.n584 VSUBS 0.030394f
C697 VTAIL.n585 VSUBS 0.013615f
C698 VTAIL.n586 VSUBS 0.012859f
C699 VTAIL.n587 VSUBS 0.02393f
C700 VTAIL.n588 VSUBS 0.02393f
C701 VTAIL.n589 VSUBS 0.012859f
C702 VTAIL.n590 VSUBS 0.013615f
C703 VTAIL.n591 VSUBS 0.030394f
C704 VTAIL.n592 VSUBS 0.030394f
C705 VTAIL.n593 VSUBS 0.013615f
C706 VTAIL.n594 VSUBS 0.012859f
C707 VTAIL.n595 VSUBS 0.02393f
C708 VTAIL.n596 VSUBS 0.02393f
C709 VTAIL.n597 VSUBS 0.012859f
C710 VTAIL.n598 VSUBS 0.012859f
C711 VTAIL.n599 VSUBS 0.013615f
C712 VTAIL.n600 VSUBS 0.030394f
C713 VTAIL.n601 VSUBS 0.030394f
C714 VTAIL.n602 VSUBS 0.030394f
C715 VTAIL.n603 VSUBS 0.013237f
C716 VTAIL.n604 VSUBS 0.012859f
C717 VTAIL.n605 VSUBS 0.02393f
C718 VTAIL.n606 VSUBS 0.02393f
C719 VTAIL.n607 VSUBS 0.012859f
C720 VTAIL.n608 VSUBS 0.013615f
C721 VTAIL.n609 VSUBS 0.030394f
C722 VTAIL.n610 VSUBS 0.030394f
C723 VTAIL.n611 VSUBS 0.013615f
C724 VTAIL.n612 VSUBS 0.012859f
C725 VTAIL.n613 VSUBS 0.02393f
C726 VTAIL.n614 VSUBS 0.02393f
C727 VTAIL.n615 VSUBS 0.012859f
C728 VTAIL.n616 VSUBS 0.013615f
C729 VTAIL.n617 VSUBS 0.030394f
C730 VTAIL.n618 VSUBS 0.030394f
C731 VTAIL.n619 VSUBS 0.013615f
C732 VTAIL.n620 VSUBS 0.012859f
C733 VTAIL.n621 VSUBS 0.02393f
C734 VTAIL.n622 VSUBS 0.02393f
C735 VTAIL.n623 VSUBS 0.012859f
C736 VTAIL.n624 VSUBS 0.013615f
C737 VTAIL.n625 VSUBS 0.030394f
C738 VTAIL.n626 VSUBS 0.075312f
C739 VTAIL.n627 VSUBS 0.013615f
C740 VTAIL.n628 VSUBS 0.012859f
C741 VTAIL.n629 VSUBS 0.053351f
C742 VTAIL.n630 VSUBS 0.037889f
C743 VTAIL.n631 VSUBS 1.55633f
C744 VDD1.t7 VSUBS 0.280176f
C745 VDD1.t5 VSUBS 0.280176f
C746 VDD1.n0 VSUBS 2.25035f
C747 VDD1.t1 VSUBS 0.280176f
C748 VDD1.t4 VSUBS 0.280176f
C749 VDD1.n1 VSUBS 2.24912f
C750 VDD1.t0 VSUBS 0.280176f
C751 VDD1.t6 VSUBS 0.280176f
C752 VDD1.n2 VSUBS 2.24912f
C753 VDD1.n3 VSUBS 3.50499f
C754 VDD1.t2 VSUBS 0.280176f
C755 VDD1.t3 VSUBS 0.280176f
C756 VDD1.n4 VSUBS 2.24096f
C757 VDD1.n5 VSUBS 3.11709f
C758 VP.n0 VSUBS 0.035662f
C759 VP.t2 VSUBS 2.37323f
C760 VP.n1 VSUBS 0.029604f
C761 VP.n2 VSUBS 0.035662f
C762 VP.t3 VSUBS 2.37323f
C763 VP.n3 VSUBS 0.028858f
C764 VP.n4 VSUBS 0.035662f
C765 VP.t6 VSUBS 2.37323f
C766 VP.n5 VSUBS 0.029604f
C767 VP.n6 VSUBS 0.035662f
C768 VP.t4 VSUBS 2.37323f
C769 VP.n7 VSUBS 0.035662f
C770 VP.t1 VSUBS 2.37323f
C771 VP.n8 VSUBS 0.029604f
C772 VP.n9 VSUBS 0.035662f
C773 VP.t0 VSUBS 2.37323f
C774 VP.n10 VSUBS 0.028858f
C775 VP.n11 VSUBS 0.227479f
C776 VP.t7 VSUBS 2.37323f
C777 VP.t5 VSUBS 2.49886f
C778 VP.n12 VSUBS 0.941855f
C779 VP.n13 VSUBS 0.904795f
C780 VP.n14 VSUBS 0.035137f
C781 VP.n15 VSUBS 0.071256f
C782 VP.n16 VSUBS 0.035662f
C783 VP.n17 VSUBS 0.035662f
C784 VP.n18 VSUBS 0.035662f
C785 VP.n19 VSUBS 0.071256f
C786 VP.n20 VSUBS 0.035137f
C787 VP.n21 VSUBS 0.843046f
C788 VP.n22 VSUBS 0.070976f
C789 VP.n23 VSUBS 0.035662f
C790 VP.n24 VSUBS 0.035662f
C791 VP.n25 VSUBS 0.035662f
C792 VP.n26 VSUBS 0.069473f
C793 VP.n27 VSUBS 0.037775f
C794 VP.n28 VSUBS 0.917735f
C795 VP.n29 VSUBS 1.84853f
C796 VP.n30 VSUBS 1.87501f
C797 VP.n31 VSUBS 0.917735f
C798 VP.n32 VSUBS 0.037775f
C799 VP.n33 VSUBS 0.069473f
C800 VP.n34 VSUBS 0.035662f
C801 VP.n35 VSUBS 0.035662f
C802 VP.n36 VSUBS 0.035662f
C803 VP.n37 VSUBS 0.070976f
C804 VP.n38 VSUBS 0.843046f
C805 VP.n39 VSUBS 0.035137f
C806 VP.n40 VSUBS 0.071256f
C807 VP.n41 VSUBS 0.035662f
C808 VP.n42 VSUBS 0.035662f
C809 VP.n43 VSUBS 0.035662f
C810 VP.n44 VSUBS 0.071256f
C811 VP.n45 VSUBS 0.035137f
C812 VP.n46 VSUBS 0.843046f
C813 VP.n47 VSUBS 0.070976f
C814 VP.n48 VSUBS 0.035662f
C815 VP.n49 VSUBS 0.035662f
C816 VP.n50 VSUBS 0.035662f
C817 VP.n51 VSUBS 0.069473f
C818 VP.n52 VSUBS 0.037775f
C819 VP.n53 VSUBS 0.917735f
C820 VP.n54 VSUBS 0.037556f
C821 B.n0 VSUBS 0.00443f
C822 B.n1 VSUBS 0.00443f
C823 B.n2 VSUBS 0.007006f
C824 B.n3 VSUBS 0.007006f
C825 B.n4 VSUBS 0.007006f
C826 B.n5 VSUBS 0.007006f
C827 B.n6 VSUBS 0.007006f
C828 B.n7 VSUBS 0.007006f
C829 B.n8 VSUBS 0.007006f
C830 B.n9 VSUBS 0.007006f
C831 B.n10 VSUBS 0.007006f
C832 B.n11 VSUBS 0.007006f
C833 B.n12 VSUBS 0.007006f
C834 B.n13 VSUBS 0.007006f
C835 B.n14 VSUBS 0.007006f
C836 B.n15 VSUBS 0.007006f
C837 B.n16 VSUBS 0.007006f
C838 B.n17 VSUBS 0.007006f
C839 B.n18 VSUBS 0.007006f
C840 B.n19 VSUBS 0.007006f
C841 B.n20 VSUBS 0.007006f
C842 B.n21 VSUBS 0.016994f
C843 B.n22 VSUBS 0.007006f
C844 B.n23 VSUBS 0.007006f
C845 B.n24 VSUBS 0.007006f
C846 B.n25 VSUBS 0.007006f
C847 B.n26 VSUBS 0.007006f
C848 B.n27 VSUBS 0.007006f
C849 B.n28 VSUBS 0.007006f
C850 B.n29 VSUBS 0.007006f
C851 B.n30 VSUBS 0.007006f
C852 B.n31 VSUBS 0.007006f
C853 B.n32 VSUBS 0.007006f
C854 B.n33 VSUBS 0.007006f
C855 B.n34 VSUBS 0.007006f
C856 B.n35 VSUBS 0.007006f
C857 B.n36 VSUBS 0.007006f
C858 B.n37 VSUBS 0.007006f
C859 B.n38 VSUBS 0.007006f
C860 B.n39 VSUBS 0.007006f
C861 B.n40 VSUBS 0.007006f
C862 B.n41 VSUBS 0.007006f
C863 B.n42 VSUBS 0.007006f
C864 B.n43 VSUBS 0.007006f
C865 B.n44 VSUBS 0.007006f
C866 B.n45 VSUBS 0.007006f
C867 B.t11 VSUBS 0.261847f
C868 B.t10 VSUBS 0.285137f
C869 B.t9 VSUBS 1.06271f
C870 B.n46 VSUBS 0.426459f
C871 B.n47 VSUBS 0.278026f
C872 B.n48 VSUBS 0.007006f
C873 B.n49 VSUBS 0.007006f
C874 B.n50 VSUBS 0.007006f
C875 B.n51 VSUBS 0.007006f
C876 B.t8 VSUBS 0.26185f
C877 B.t7 VSUBS 0.28514f
C878 B.t6 VSUBS 1.06271f
C879 B.n52 VSUBS 0.426456f
C880 B.n53 VSUBS 0.278023f
C881 B.n54 VSUBS 0.016231f
C882 B.n55 VSUBS 0.007006f
C883 B.n56 VSUBS 0.007006f
C884 B.n57 VSUBS 0.007006f
C885 B.n58 VSUBS 0.007006f
C886 B.n59 VSUBS 0.007006f
C887 B.n60 VSUBS 0.007006f
C888 B.n61 VSUBS 0.007006f
C889 B.n62 VSUBS 0.007006f
C890 B.n63 VSUBS 0.007006f
C891 B.n64 VSUBS 0.007006f
C892 B.n65 VSUBS 0.007006f
C893 B.n66 VSUBS 0.007006f
C894 B.n67 VSUBS 0.007006f
C895 B.n68 VSUBS 0.007006f
C896 B.n69 VSUBS 0.007006f
C897 B.n70 VSUBS 0.007006f
C898 B.n71 VSUBS 0.007006f
C899 B.n72 VSUBS 0.007006f
C900 B.n73 VSUBS 0.007006f
C901 B.n74 VSUBS 0.007006f
C902 B.n75 VSUBS 0.007006f
C903 B.n76 VSUBS 0.007006f
C904 B.n77 VSUBS 0.007006f
C905 B.n78 VSUBS 0.016174f
C906 B.n79 VSUBS 0.007006f
C907 B.n80 VSUBS 0.007006f
C908 B.n81 VSUBS 0.007006f
C909 B.n82 VSUBS 0.007006f
C910 B.n83 VSUBS 0.007006f
C911 B.n84 VSUBS 0.007006f
C912 B.n85 VSUBS 0.007006f
C913 B.n86 VSUBS 0.007006f
C914 B.n87 VSUBS 0.007006f
C915 B.n88 VSUBS 0.007006f
C916 B.n89 VSUBS 0.007006f
C917 B.n90 VSUBS 0.007006f
C918 B.n91 VSUBS 0.007006f
C919 B.n92 VSUBS 0.007006f
C920 B.n93 VSUBS 0.007006f
C921 B.n94 VSUBS 0.007006f
C922 B.n95 VSUBS 0.007006f
C923 B.n96 VSUBS 0.007006f
C924 B.n97 VSUBS 0.007006f
C925 B.n98 VSUBS 0.007006f
C926 B.n99 VSUBS 0.007006f
C927 B.n100 VSUBS 0.007006f
C928 B.n101 VSUBS 0.007006f
C929 B.n102 VSUBS 0.007006f
C930 B.n103 VSUBS 0.007006f
C931 B.n104 VSUBS 0.007006f
C932 B.n105 VSUBS 0.007006f
C933 B.n106 VSUBS 0.007006f
C934 B.n107 VSUBS 0.007006f
C935 B.n108 VSUBS 0.007006f
C936 B.n109 VSUBS 0.007006f
C937 B.n110 VSUBS 0.007006f
C938 B.n111 VSUBS 0.007006f
C939 B.n112 VSUBS 0.007006f
C940 B.n113 VSUBS 0.007006f
C941 B.n114 VSUBS 0.007006f
C942 B.n115 VSUBS 0.007006f
C943 B.n116 VSUBS 0.007006f
C944 B.n117 VSUBS 0.016994f
C945 B.n118 VSUBS 0.007006f
C946 B.n119 VSUBS 0.007006f
C947 B.n120 VSUBS 0.007006f
C948 B.n121 VSUBS 0.007006f
C949 B.n122 VSUBS 0.007006f
C950 B.n123 VSUBS 0.007006f
C951 B.n124 VSUBS 0.007006f
C952 B.n125 VSUBS 0.007006f
C953 B.n126 VSUBS 0.007006f
C954 B.n127 VSUBS 0.007006f
C955 B.n128 VSUBS 0.007006f
C956 B.n129 VSUBS 0.007006f
C957 B.n130 VSUBS 0.007006f
C958 B.n131 VSUBS 0.007006f
C959 B.n132 VSUBS 0.007006f
C960 B.n133 VSUBS 0.007006f
C961 B.n134 VSUBS 0.007006f
C962 B.n135 VSUBS 0.007006f
C963 B.n136 VSUBS 0.007006f
C964 B.n137 VSUBS 0.007006f
C965 B.n138 VSUBS 0.007006f
C966 B.n139 VSUBS 0.007006f
C967 B.n140 VSUBS 0.007006f
C968 B.n141 VSUBS 0.007006f
C969 B.t4 VSUBS 0.26185f
C970 B.t5 VSUBS 0.28514f
C971 B.t3 VSUBS 1.06271f
C972 B.n142 VSUBS 0.426456f
C973 B.n143 VSUBS 0.278023f
C974 B.n144 VSUBS 0.007006f
C975 B.n145 VSUBS 0.007006f
C976 B.n146 VSUBS 0.007006f
C977 B.n147 VSUBS 0.007006f
C978 B.t1 VSUBS 0.261847f
C979 B.t2 VSUBS 0.285137f
C980 B.t0 VSUBS 1.06271f
C981 B.n148 VSUBS 0.426459f
C982 B.n149 VSUBS 0.278026f
C983 B.n150 VSUBS 0.016231f
C984 B.n151 VSUBS 0.007006f
C985 B.n152 VSUBS 0.007006f
C986 B.n153 VSUBS 0.007006f
C987 B.n154 VSUBS 0.007006f
C988 B.n155 VSUBS 0.007006f
C989 B.n156 VSUBS 0.007006f
C990 B.n157 VSUBS 0.007006f
C991 B.n158 VSUBS 0.007006f
C992 B.n159 VSUBS 0.007006f
C993 B.n160 VSUBS 0.007006f
C994 B.n161 VSUBS 0.007006f
C995 B.n162 VSUBS 0.007006f
C996 B.n163 VSUBS 0.007006f
C997 B.n164 VSUBS 0.007006f
C998 B.n165 VSUBS 0.007006f
C999 B.n166 VSUBS 0.007006f
C1000 B.n167 VSUBS 0.007006f
C1001 B.n168 VSUBS 0.007006f
C1002 B.n169 VSUBS 0.007006f
C1003 B.n170 VSUBS 0.007006f
C1004 B.n171 VSUBS 0.007006f
C1005 B.n172 VSUBS 0.007006f
C1006 B.n173 VSUBS 0.007006f
C1007 B.n174 VSUBS 0.016994f
C1008 B.n175 VSUBS 0.007006f
C1009 B.n176 VSUBS 0.007006f
C1010 B.n177 VSUBS 0.007006f
C1011 B.n178 VSUBS 0.007006f
C1012 B.n179 VSUBS 0.007006f
C1013 B.n180 VSUBS 0.007006f
C1014 B.n181 VSUBS 0.007006f
C1015 B.n182 VSUBS 0.007006f
C1016 B.n183 VSUBS 0.007006f
C1017 B.n184 VSUBS 0.007006f
C1018 B.n185 VSUBS 0.007006f
C1019 B.n186 VSUBS 0.007006f
C1020 B.n187 VSUBS 0.007006f
C1021 B.n188 VSUBS 0.007006f
C1022 B.n189 VSUBS 0.007006f
C1023 B.n190 VSUBS 0.007006f
C1024 B.n191 VSUBS 0.007006f
C1025 B.n192 VSUBS 0.007006f
C1026 B.n193 VSUBS 0.007006f
C1027 B.n194 VSUBS 0.007006f
C1028 B.n195 VSUBS 0.007006f
C1029 B.n196 VSUBS 0.007006f
C1030 B.n197 VSUBS 0.007006f
C1031 B.n198 VSUBS 0.007006f
C1032 B.n199 VSUBS 0.007006f
C1033 B.n200 VSUBS 0.007006f
C1034 B.n201 VSUBS 0.007006f
C1035 B.n202 VSUBS 0.007006f
C1036 B.n203 VSUBS 0.007006f
C1037 B.n204 VSUBS 0.007006f
C1038 B.n205 VSUBS 0.007006f
C1039 B.n206 VSUBS 0.007006f
C1040 B.n207 VSUBS 0.007006f
C1041 B.n208 VSUBS 0.007006f
C1042 B.n209 VSUBS 0.007006f
C1043 B.n210 VSUBS 0.007006f
C1044 B.n211 VSUBS 0.007006f
C1045 B.n212 VSUBS 0.007006f
C1046 B.n213 VSUBS 0.007006f
C1047 B.n214 VSUBS 0.007006f
C1048 B.n215 VSUBS 0.007006f
C1049 B.n216 VSUBS 0.007006f
C1050 B.n217 VSUBS 0.007006f
C1051 B.n218 VSUBS 0.007006f
C1052 B.n219 VSUBS 0.007006f
C1053 B.n220 VSUBS 0.007006f
C1054 B.n221 VSUBS 0.007006f
C1055 B.n222 VSUBS 0.007006f
C1056 B.n223 VSUBS 0.007006f
C1057 B.n224 VSUBS 0.007006f
C1058 B.n225 VSUBS 0.007006f
C1059 B.n226 VSUBS 0.007006f
C1060 B.n227 VSUBS 0.007006f
C1061 B.n228 VSUBS 0.007006f
C1062 B.n229 VSUBS 0.007006f
C1063 B.n230 VSUBS 0.007006f
C1064 B.n231 VSUBS 0.007006f
C1065 B.n232 VSUBS 0.007006f
C1066 B.n233 VSUBS 0.007006f
C1067 B.n234 VSUBS 0.007006f
C1068 B.n235 VSUBS 0.007006f
C1069 B.n236 VSUBS 0.007006f
C1070 B.n237 VSUBS 0.007006f
C1071 B.n238 VSUBS 0.007006f
C1072 B.n239 VSUBS 0.007006f
C1073 B.n240 VSUBS 0.007006f
C1074 B.n241 VSUBS 0.007006f
C1075 B.n242 VSUBS 0.007006f
C1076 B.n243 VSUBS 0.007006f
C1077 B.n244 VSUBS 0.007006f
C1078 B.n245 VSUBS 0.007006f
C1079 B.n246 VSUBS 0.007006f
C1080 B.n247 VSUBS 0.015973f
C1081 B.n248 VSUBS 0.015973f
C1082 B.n249 VSUBS 0.016994f
C1083 B.n250 VSUBS 0.007006f
C1084 B.n251 VSUBS 0.007006f
C1085 B.n252 VSUBS 0.007006f
C1086 B.n253 VSUBS 0.007006f
C1087 B.n254 VSUBS 0.007006f
C1088 B.n255 VSUBS 0.007006f
C1089 B.n256 VSUBS 0.007006f
C1090 B.n257 VSUBS 0.007006f
C1091 B.n258 VSUBS 0.007006f
C1092 B.n259 VSUBS 0.007006f
C1093 B.n260 VSUBS 0.007006f
C1094 B.n261 VSUBS 0.007006f
C1095 B.n262 VSUBS 0.007006f
C1096 B.n263 VSUBS 0.007006f
C1097 B.n264 VSUBS 0.007006f
C1098 B.n265 VSUBS 0.007006f
C1099 B.n266 VSUBS 0.007006f
C1100 B.n267 VSUBS 0.007006f
C1101 B.n268 VSUBS 0.007006f
C1102 B.n269 VSUBS 0.007006f
C1103 B.n270 VSUBS 0.007006f
C1104 B.n271 VSUBS 0.007006f
C1105 B.n272 VSUBS 0.007006f
C1106 B.n273 VSUBS 0.007006f
C1107 B.n274 VSUBS 0.007006f
C1108 B.n275 VSUBS 0.007006f
C1109 B.n276 VSUBS 0.007006f
C1110 B.n277 VSUBS 0.007006f
C1111 B.n278 VSUBS 0.007006f
C1112 B.n279 VSUBS 0.007006f
C1113 B.n280 VSUBS 0.007006f
C1114 B.n281 VSUBS 0.007006f
C1115 B.n282 VSUBS 0.007006f
C1116 B.n283 VSUBS 0.007006f
C1117 B.n284 VSUBS 0.007006f
C1118 B.n285 VSUBS 0.007006f
C1119 B.n286 VSUBS 0.007006f
C1120 B.n287 VSUBS 0.007006f
C1121 B.n288 VSUBS 0.007006f
C1122 B.n289 VSUBS 0.007006f
C1123 B.n290 VSUBS 0.007006f
C1124 B.n291 VSUBS 0.007006f
C1125 B.n292 VSUBS 0.007006f
C1126 B.n293 VSUBS 0.007006f
C1127 B.n294 VSUBS 0.007006f
C1128 B.n295 VSUBS 0.007006f
C1129 B.n296 VSUBS 0.007006f
C1130 B.n297 VSUBS 0.007006f
C1131 B.n298 VSUBS 0.007006f
C1132 B.n299 VSUBS 0.007006f
C1133 B.n300 VSUBS 0.007006f
C1134 B.n301 VSUBS 0.007006f
C1135 B.n302 VSUBS 0.007006f
C1136 B.n303 VSUBS 0.007006f
C1137 B.n304 VSUBS 0.007006f
C1138 B.n305 VSUBS 0.007006f
C1139 B.n306 VSUBS 0.007006f
C1140 B.n307 VSUBS 0.007006f
C1141 B.n308 VSUBS 0.007006f
C1142 B.n309 VSUBS 0.007006f
C1143 B.n310 VSUBS 0.007006f
C1144 B.n311 VSUBS 0.007006f
C1145 B.n312 VSUBS 0.007006f
C1146 B.n313 VSUBS 0.007006f
C1147 B.n314 VSUBS 0.007006f
C1148 B.n315 VSUBS 0.007006f
C1149 B.n316 VSUBS 0.007006f
C1150 B.n317 VSUBS 0.007006f
C1151 B.n318 VSUBS 0.007006f
C1152 B.n319 VSUBS 0.006594f
C1153 B.n320 VSUBS 0.007006f
C1154 B.n321 VSUBS 0.007006f
C1155 B.n322 VSUBS 0.003915f
C1156 B.n323 VSUBS 0.007006f
C1157 B.n324 VSUBS 0.007006f
C1158 B.n325 VSUBS 0.007006f
C1159 B.n326 VSUBS 0.007006f
C1160 B.n327 VSUBS 0.007006f
C1161 B.n328 VSUBS 0.007006f
C1162 B.n329 VSUBS 0.007006f
C1163 B.n330 VSUBS 0.007006f
C1164 B.n331 VSUBS 0.007006f
C1165 B.n332 VSUBS 0.007006f
C1166 B.n333 VSUBS 0.007006f
C1167 B.n334 VSUBS 0.007006f
C1168 B.n335 VSUBS 0.003915f
C1169 B.n336 VSUBS 0.016231f
C1170 B.n337 VSUBS 0.006594f
C1171 B.n338 VSUBS 0.007006f
C1172 B.n339 VSUBS 0.007006f
C1173 B.n340 VSUBS 0.007006f
C1174 B.n341 VSUBS 0.007006f
C1175 B.n342 VSUBS 0.007006f
C1176 B.n343 VSUBS 0.007006f
C1177 B.n344 VSUBS 0.007006f
C1178 B.n345 VSUBS 0.007006f
C1179 B.n346 VSUBS 0.007006f
C1180 B.n347 VSUBS 0.007006f
C1181 B.n348 VSUBS 0.007006f
C1182 B.n349 VSUBS 0.007006f
C1183 B.n350 VSUBS 0.007006f
C1184 B.n351 VSUBS 0.007006f
C1185 B.n352 VSUBS 0.007006f
C1186 B.n353 VSUBS 0.007006f
C1187 B.n354 VSUBS 0.007006f
C1188 B.n355 VSUBS 0.007006f
C1189 B.n356 VSUBS 0.007006f
C1190 B.n357 VSUBS 0.007006f
C1191 B.n358 VSUBS 0.007006f
C1192 B.n359 VSUBS 0.007006f
C1193 B.n360 VSUBS 0.007006f
C1194 B.n361 VSUBS 0.007006f
C1195 B.n362 VSUBS 0.007006f
C1196 B.n363 VSUBS 0.007006f
C1197 B.n364 VSUBS 0.007006f
C1198 B.n365 VSUBS 0.007006f
C1199 B.n366 VSUBS 0.007006f
C1200 B.n367 VSUBS 0.007006f
C1201 B.n368 VSUBS 0.007006f
C1202 B.n369 VSUBS 0.007006f
C1203 B.n370 VSUBS 0.007006f
C1204 B.n371 VSUBS 0.007006f
C1205 B.n372 VSUBS 0.007006f
C1206 B.n373 VSUBS 0.007006f
C1207 B.n374 VSUBS 0.007006f
C1208 B.n375 VSUBS 0.007006f
C1209 B.n376 VSUBS 0.007006f
C1210 B.n377 VSUBS 0.007006f
C1211 B.n378 VSUBS 0.007006f
C1212 B.n379 VSUBS 0.007006f
C1213 B.n380 VSUBS 0.007006f
C1214 B.n381 VSUBS 0.007006f
C1215 B.n382 VSUBS 0.007006f
C1216 B.n383 VSUBS 0.007006f
C1217 B.n384 VSUBS 0.007006f
C1218 B.n385 VSUBS 0.007006f
C1219 B.n386 VSUBS 0.007006f
C1220 B.n387 VSUBS 0.007006f
C1221 B.n388 VSUBS 0.007006f
C1222 B.n389 VSUBS 0.007006f
C1223 B.n390 VSUBS 0.007006f
C1224 B.n391 VSUBS 0.007006f
C1225 B.n392 VSUBS 0.007006f
C1226 B.n393 VSUBS 0.007006f
C1227 B.n394 VSUBS 0.007006f
C1228 B.n395 VSUBS 0.007006f
C1229 B.n396 VSUBS 0.007006f
C1230 B.n397 VSUBS 0.007006f
C1231 B.n398 VSUBS 0.007006f
C1232 B.n399 VSUBS 0.007006f
C1233 B.n400 VSUBS 0.007006f
C1234 B.n401 VSUBS 0.007006f
C1235 B.n402 VSUBS 0.007006f
C1236 B.n403 VSUBS 0.007006f
C1237 B.n404 VSUBS 0.007006f
C1238 B.n405 VSUBS 0.007006f
C1239 B.n406 VSUBS 0.007006f
C1240 B.n407 VSUBS 0.007006f
C1241 B.n408 VSUBS 0.016994f
C1242 B.n409 VSUBS 0.015973f
C1243 B.n410 VSUBS 0.015973f
C1244 B.n411 VSUBS 0.007006f
C1245 B.n412 VSUBS 0.007006f
C1246 B.n413 VSUBS 0.007006f
C1247 B.n414 VSUBS 0.007006f
C1248 B.n415 VSUBS 0.007006f
C1249 B.n416 VSUBS 0.007006f
C1250 B.n417 VSUBS 0.007006f
C1251 B.n418 VSUBS 0.007006f
C1252 B.n419 VSUBS 0.007006f
C1253 B.n420 VSUBS 0.007006f
C1254 B.n421 VSUBS 0.007006f
C1255 B.n422 VSUBS 0.007006f
C1256 B.n423 VSUBS 0.007006f
C1257 B.n424 VSUBS 0.007006f
C1258 B.n425 VSUBS 0.007006f
C1259 B.n426 VSUBS 0.007006f
C1260 B.n427 VSUBS 0.007006f
C1261 B.n428 VSUBS 0.007006f
C1262 B.n429 VSUBS 0.007006f
C1263 B.n430 VSUBS 0.007006f
C1264 B.n431 VSUBS 0.007006f
C1265 B.n432 VSUBS 0.007006f
C1266 B.n433 VSUBS 0.007006f
C1267 B.n434 VSUBS 0.007006f
C1268 B.n435 VSUBS 0.007006f
C1269 B.n436 VSUBS 0.007006f
C1270 B.n437 VSUBS 0.007006f
C1271 B.n438 VSUBS 0.007006f
C1272 B.n439 VSUBS 0.007006f
C1273 B.n440 VSUBS 0.007006f
C1274 B.n441 VSUBS 0.007006f
C1275 B.n442 VSUBS 0.007006f
C1276 B.n443 VSUBS 0.007006f
C1277 B.n444 VSUBS 0.007006f
C1278 B.n445 VSUBS 0.007006f
C1279 B.n446 VSUBS 0.007006f
C1280 B.n447 VSUBS 0.007006f
C1281 B.n448 VSUBS 0.007006f
C1282 B.n449 VSUBS 0.007006f
C1283 B.n450 VSUBS 0.007006f
C1284 B.n451 VSUBS 0.007006f
C1285 B.n452 VSUBS 0.007006f
C1286 B.n453 VSUBS 0.007006f
C1287 B.n454 VSUBS 0.007006f
C1288 B.n455 VSUBS 0.007006f
C1289 B.n456 VSUBS 0.007006f
C1290 B.n457 VSUBS 0.007006f
C1291 B.n458 VSUBS 0.007006f
C1292 B.n459 VSUBS 0.007006f
C1293 B.n460 VSUBS 0.007006f
C1294 B.n461 VSUBS 0.007006f
C1295 B.n462 VSUBS 0.007006f
C1296 B.n463 VSUBS 0.007006f
C1297 B.n464 VSUBS 0.007006f
C1298 B.n465 VSUBS 0.007006f
C1299 B.n466 VSUBS 0.007006f
C1300 B.n467 VSUBS 0.007006f
C1301 B.n468 VSUBS 0.007006f
C1302 B.n469 VSUBS 0.007006f
C1303 B.n470 VSUBS 0.007006f
C1304 B.n471 VSUBS 0.007006f
C1305 B.n472 VSUBS 0.007006f
C1306 B.n473 VSUBS 0.007006f
C1307 B.n474 VSUBS 0.007006f
C1308 B.n475 VSUBS 0.007006f
C1309 B.n476 VSUBS 0.007006f
C1310 B.n477 VSUBS 0.007006f
C1311 B.n478 VSUBS 0.007006f
C1312 B.n479 VSUBS 0.007006f
C1313 B.n480 VSUBS 0.007006f
C1314 B.n481 VSUBS 0.007006f
C1315 B.n482 VSUBS 0.007006f
C1316 B.n483 VSUBS 0.007006f
C1317 B.n484 VSUBS 0.007006f
C1318 B.n485 VSUBS 0.007006f
C1319 B.n486 VSUBS 0.007006f
C1320 B.n487 VSUBS 0.007006f
C1321 B.n488 VSUBS 0.007006f
C1322 B.n489 VSUBS 0.007006f
C1323 B.n490 VSUBS 0.007006f
C1324 B.n491 VSUBS 0.007006f
C1325 B.n492 VSUBS 0.007006f
C1326 B.n493 VSUBS 0.007006f
C1327 B.n494 VSUBS 0.007006f
C1328 B.n495 VSUBS 0.007006f
C1329 B.n496 VSUBS 0.007006f
C1330 B.n497 VSUBS 0.007006f
C1331 B.n498 VSUBS 0.007006f
C1332 B.n499 VSUBS 0.007006f
C1333 B.n500 VSUBS 0.007006f
C1334 B.n501 VSUBS 0.007006f
C1335 B.n502 VSUBS 0.007006f
C1336 B.n503 VSUBS 0.007006f
C1337 B.n504 VSUBS 0.007006f
C1338 B.n505 VSUBS 0.007006f
C1339 B.n506 VSUBS 0.007006f
C1340 B.n507 VSUBS 0.007006f
C1341 B.n508 VSUBS 0.007006f
C1342 B.n509 VSUBS 0.007006f
C1343 B.n510 VSUBS 0.007006f
C1344 B.n511 VSUBS 0.007006f
C1345 B.n512 VSUBS 0.007006f
C1346 B.n513 VSUBS 0.007006f
C1347 B.n514 VSUBS 0.007006f
C1348 B.n515 VSUBS 0.007006f
C1349 B.n516 VSUBS 0.007006f
C1350 B.n517 VSUBS 0.007006f
C1351 B.n518 VSUBS 0.007006f
C1352 B.n519 VSUBS 0.007006f
C1353 B.n520 VSUBS 0.007006f
C1354 B.n521 VSUBS 0.007006f
C1355 B.n522 VSUBS 0.007006f
C1356 B.n523 VSUBS 0.016794f
C1357 B.n524 VSUBS 0.015973f
C1358 B.n525 VSUBS 0.016994f
C1359 B.n526 VSUBS 0.007006f
C1360 B.n527 VSUBS 0.007006f
C1361 B.n528 VSUBS 0.007006f
C1362 B.n529 VSUBS 0.007006f
C1363 B.n530 VSUBS 0.007006f
C1364 B.n531 VSUBS 0.007006f
C1365 B.n532 VSUBS 0.007006f
C1366 B.n533 VSUBS 0.007006f
C1367 B.n534 VSUBS 0.007006f
C1368 B.n535 VSUBS 0.007006f
C1369 B.n536 VSUBS 0.007006f
C1370 B.n537 VSUBS 0.007006f
C1371 B.n538 VSUBS 0.007006f
C1372 B.n539 VSUBS 0.007006f
C1373 B.n540 VSUBS 0.007006f
C1374 B.n541 VSUBS 0.007006f
C1375 B.n542 VSUBS 0.007006f
C1376 B.n543 VSUBS 0.007006f
C1377 B.n544 VSUBS 0.007006f
C1378 B.n545 VSUBS 0.007006f
C1379 B.n546 VSUBS 0.007006f
C1380 B.n547 VSUBS 0.007006f
C1381 B.n548 VSUBS 0.007006f
C1382 B.n549 VSUBS 0.007006f
C1383 B.n550 VSUBS 0.007006f
C1384 B.n551 VSUBS 0.007006f
C1385 B.n552 VSUBS 0.007006f
C1386 B.n553 VSUBS 0.007006f
C1387 B.n554 VSUBS 0.007006f
C1388 B.n555 VSUBS 0.007006f
C1389 B.n556 VSUBS 0.007006f
C1390 B.n557 VSUBS 0.007006f
C1391 B.n558 VSUBS 0.007006f
C1392 B.n559 VSUBS 0.007006f
C1393 B.n560 VSUBS 0.007006f
C1394 B.n561 VSUBS 0.007006f
C1395 B.n562 VSUBS 0.007006f
C1396 B.n563 VSUBS 0.007006f
C1397 B.n564 VSUBS 0.007006f
C1398 B.n565 VSUBS 0.007006f
C1399 B.n566 VSUBS 0.007006f
C1400 B.n567 VSUBS 0.007006f
C1401 B.n568 VSUBS 0.007006f
C1402 B.n569 VSUBS 0.007006f
C1403 B.n570 VSUBS 0.007006f
C1404 B.n571 VSUBS 0.007006f
C1405 B.n572 VSUBS 0.007006f
C1406 B.n573 VSUBS 0.007006f
C1407 B.n574 VSUBS 0.007006f
C1408 B.n575 VSUBS 0.007006f
C1409 B.n576 VSUBS 0.007006f
C1410 B.n577 VSUBS 0.007006f
C1411 B.n578 VSUBS 0.007006f
C1412 B.n579 VSUBS 0.007006f
C1413 B.n580 VSUBS 0.007006f
C1414 B.n581 VSUBS 0.007006f
C1415 B.n582 VSUBS 0.007006f
C1416 B.n583 VSUBS 0.007006f
C1417 B.n584 VSUBS 0.007006f
C1418 B.n585 VSUBS 0.007006f
C1419 B.n586 VSUBS 0.007006f
C1420 B.n587 VSUBS 0.007006f
C1421 B.n588 VSUBS 0.007006f
C1422 B.n589 VSUBS 0.007006f
C1423 B.n590 VSUBS 0.007006f
C1424 B.n591 VSUBS 0.007006f
C1425 B.n592 VSUBS 0.007006f
C1426 B.n593 VSUBS 0.007006f
C1427 B.n594 VSUBS 0.007006f
C1428 B.n595 VSUBS 0.006594f
C1429 B.n596 VSUBS 0.007006f
C1430 B.n597 VSUBS 0.007006f
C1431 B.n598 VSUBS 0.003915f
C1432 B.n599 VSUBS 0.007006f
C1433 B.n600 VSUBS 0.007006f
C1434 B.n601 VSUBS 0.007006f
C1435 B.n602 VSUBS 0.007006f
C1436 B.n603 VSUBS 0.007006f
C1437 B.n604 VSUBS 0.007006f
C1438 B.n605 VSUBS 0.007006f
C1439 B.n606 VSUBS 0.007006f
C1440 B.n607 VSUBS 0.007006f
C1441 B.n608 VSUBS 0.007006f
C1442 B.n609 VSUBS 0.007006f
C1443 B.n610 VSUBS 0.007006f
C1444 B.n611 VSUBS 0.003915f
C1445 B.n612 VSUBS 0.016231f
C1446 B.n613 VSUBS 0.006594f
C1447 B.n614 VSUBS 0.007006f
C1448 B.n615 VSUBS 0.007006f
C1449 B.n616 VSUBS 0.007006f
C1450 B.n617 VSUBS 0.007006f
C1451 B.n618 VSUBS 0.007006f
C1452 B.n619 VSUBS 0.007006f
C1453 B.n620 VSUBS 0.007006f
C1454 B.n621 VSUBS 0.007006f
C1455 B.n622 VSUBS 0.007006f
C1456 B.n623 VSUBS 0.007006f
C1457 B.n624 VSUBS 0.007006f
C1458 B.n625 VSUBS 0.007006f
C1459 B.n626 VSUBS 0.007006f
C1460 B.n627 VSUBS 0.007006f
C1461 B.n628 VSUBS 0.007006f
C1462 B.n629 VSUBS 0.007006f
C1463 B.n630 VSUBS 0.007006f
C1464 B.n631 VSUBS 0.007006f
C1465 B.n632 VSUBS 0.007006f
C1466 B.n633 VSUBS 0.007006f
C1467 B.n634 VSUBS 0.007006f
C1468 B.n635 VSUBS 0.007006f
C1469 B.n636 VSUBS 0.007006f
C1470 B.n637 VSUBS 0.007006f
C1471 B.n638 VSUBS 0.007006f
C1472 B.n639 VSUBS 0.007006f
C1473 B.n640 VSUBS 0.007006f
C1474 B.n641 VSUBS 0.007006f
C1475 B.n642 VSUBS 0.007006f
C1476 B.n643 VSUBS 0.007006f
C1477 B.n644 VSUBS 0.007006f
C1478 B.n645 VSUBS 0.007006f
C1479 B.n646 VSUBS 0.007006f
C1480 B.n647 VSUBS 0.007006f
C1481 B.n648 VSUBS 0.007006f
C1482 B.n649 VSUBS 0.007006f
C1483 B.n650 VSUBS 0.007006f
C1484 B.n651 VSUBS 0.007006f
C1485 B.n652 VSUBS 0.007006f
C1486 B.n653 VSUBS 0.007006f
C1487 B.n654 VSUBS 0.007006f
C1488 B.n655 VSUBS 0.007006f
C1489 B.n656 VSUBS 0.007006f
C1490 B.n657 VSUBS 0.007006f
C1491 B.n658 VSUBS 0.007006f
C1492 B.n659 VSUBS 0.007006f
C1493 B.n660 VSUBS 0.007006f
C1494 B.n661 VSUBS 0.007006f
C1495 B.n662 VSUBS 0.007006f
C1496 B.n663 VSUBS 0.007006f
C1497 B.n664 VSUBS 0.007006f
C1498 B.n665 VSUBS 0.007006f
C1499 B.n666 VSUBS 0.007006f
C1500 B.n667 VSUBS 0.007006f
C1501 B.n668 VSUBS 0.007006f
C1502 B.n669 VSUBS 0.007006f
C1503 B.n670 VSUBS 0.007006f
C1504 B.n671 VSUBS 0.007006f
C1505 B.n672 VSUBS 0.007006f
C1506 B.n673 VSUBS 0.007006f
C1507 B.n674 VSUBS 0.007006f
C1508 B.n675 VSUBS 0.007006f
C1509 B.n676 VSUBS 0.007006f
C1510 B.n677 VSUBS 0.007006f
C1511 B.n678 VSUBS 0.007006f
C1512 B.n679 VSUBS 0.007006f
C1513 B.n680 VSUBS 0.007006f
C1514 B.n681 VSUBS 0.007006f
C1515 B.n682 VSUBS 0.007006f
C1516 B.n683 VSUBS 0.007006f
C1517 B.n684 VSUBS 0.016994f
C1518 B.n685 VSUBS 0.015973f
C1519 B.n686 VSUBS 0.015973f
C1520 B.n687 VSUBS 0.007006f
C1521 B.n688 VSUBS 0.007006f
C1522 B.n689 VSUBS 0.007006f
C1523 B.n690 VSUBS 0.007006f
C1524 B.n691 VSUBS 0.007006f
C1525 B.n692 VSUBS 0.007006f
C1526 B.n693 VSUBS 0.007006f
C1527 B.n694 VSUBS 0.007006f
C1528 B.n695 VSUBS 0.007006f
C1529 B.n696 VSUBS 0.007006f
C1530 B.n697 VSUBS 0.007006f
C1531 B.n698 VSUBS 0.007006f
C1532 B.n699 VSUBS 0.007006f
C1533 B.n700 VSUBS 0.007006f
C1534 B.n701 VSUBS 0.007006f
C1535 B.n702 VSUBS 0.007006f
C1536 B.n703 VSUBS 0.007006f
C1537 B.n704 VSUBS 0.007006f
C1538 B.n705 VSUBS 0.007006f
C1539 B.n706 VSUBS 0.007006f
C1540 B.n707 VSUBS 0.007006f
C1541 B.n708 VSUBS 0.007006f
C1542 B.n709 VSUBS 0.007006f
C1543 B.n710 VSUBS 0.007006f
C1544 B.n711 VSUBS 0.007006f
C1545 B.n712 VSUBS 0.007006f
C1546 B.n713 VSUBS 0.007006f
C1547 B.n714 VSUBS 0.007006f
C1548 B.n715 VSUBS 0.007006f
C1549 B.n716 VSUBS 0.007006f
C1550 B.n717 VSUBS 0.007006f
C1551 B.n718 VSUBS 0.007006f
C1552 B.n719 VSUBS 0.007006f
C1553 B.n720 VSUBS 0.007006f
C1554 B.n721 VSUBS 0.007006f
C1555 B.n722 VSUBS 0.007006f
C1556 B.n723 VSUBS 0.007006f
C1557 B.n724 VSUBS 0.007006f
C1558 B.n725 VSUBS 0.007006f
C1559 B.n726 VSUBS 0.007006f
C1560 B.n727 VSUBS 0.007006f
C1561 B.n728 VSUBS 0.007006f
C1562 B.n729 VSUBS 0.007006f
C1563 B.n730 VSUBS 0.007006f
C1564 B.n731 VSUBS 0.007006f
C1565 B.n732 VSUBS 0.007006f
C1566 B.n733 VSUBS 0.007006f
C1567 B.n734 VSUBS 0.007006f
C1568 B.n735 VSUBS 0.007006f
C1569 B.n736 VSUBS 0.007006f
C1570 B.n737 VSUBS 0.007006f
C1571 B.n738 VSUBS 0.007006f
C1572 B.n739 VSUBS 0.007006f
C1573 B.n740 VSUBS 0.007006f
C1574 B.n741 VSUBS 0.007006f
C1575 B.n742 VSUBS 0.007006f
C1576 B.n743 VSUBS 0.015863f
.ends

