* NGSPICE file created from diff_pair_sample_0991.ext - technology: sky130A

.subckt diff_pair_sample_0991 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t11 VP.t0 VDD1.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=3.14325 pd=19.38 as=3.14325 ps=19.38 w=19.05 l=2.18
X1 VDD2.t5 VN.t0 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=3.14325 pd=19.38 as=7.4295 ps=38.88 w=19.05 l=2.18
X2 VDD1.t0 VP.t1 VTAIL.t10 B.t3 sky130_fd_pr__nfet_01v8 ad=3.14325 pd=19.38 as=7.4295 ps=38.88 w=19.05 l=2.18
X3 VDD1.t5 VP.t2 VTAIL.t9 B.t2 sky130_fd_pr__nfet_01v8 ad=3.14325 pd=19.38 as=7.4295 ps=38.88 w=19.05 l=2.18
X4 B.t19 B.t17 B.t18 B.t14 sky130_fd_pr__nfet_01v8 ad=7.4295 pd=38.88 as=0 ps=0 w=19.05 l=2.18
X5 VTAIL.t8 VP.t3 VDD1.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=3.14325 pd=19.38 as=3.14325 ps=19.38 w=19.05 l=2.18
X6 VDD2.t4 VN.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=7.4295 pd=38.88 as=3.14325 ps=19.38 w=19.05 l=2.18
X7 VTAIL.t4 VN.t2 VDD2.t3 B.t4 sky130_fd_pr__nfet_01v8 ad=3.14325 pd=19.38 as=3.14325 ps=19.38 w=19.05 l=2.18
X8 VTAIL.t0 VN.t3 VDD2.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=3.14325 pd=19.38 as=3.14325 ps=19.38 w=19.05 l=2.18
X9 VDD2.t1 VN.t4 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=7.4295 pd=38.88 as=3.14325 ps=19.38 w=19.05 l=2.18
X10 VDD1.t3 VP.t4 VTAIL.t7 B.t5 sky130_fd_pr__nfet_01v8 ad=7.4295 pd=38.88 as=3.14325 ps=19.38 w=19.05 l=2.18
X11 B.t16 B.t13 B.t15 B.t14 sky130_fd_pr__nfet_01v8 ad=7.4295 pd=38.88 as=0 ps=0 w=19.05 l=2.18
X12 VDD2.t0 VN.t5 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=3.14325 pd=19.38 as=7.4295 ps=38.88 w=19.05 l=2.18
X13 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=7.4295 pd=38.88 as=0 ps=0 w=19.05 l=2.18
X14 VDD1.t2 VP.t5 VTAIL.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=7.4295 pd=38.88 as=3.14325 ps=19.38 w=19.05 l=2.18
X15 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=7.4295 pd=38.88 as=0 ps=0 w=19.05 l=2.18
R0 VP.n9 VP.t4 242.743
R1 VP.n5 VP.t5 210.6
R2 VP.n29 VP.t0 210.6
R3 VP.n37 VP.t1 210.6
R4 VP.n18 VP.t2 210.6
R5 VP.n10 VP.t3 210.6
R6 VP.n11 VP.n8 161.3
R7 VP.n13 VP.n12 161.3
R8 VP.n14 VP.n7 161.3
R9 VP.n16 VP.n15 161.3
R10 VP.n17 VP.n6 161.3
R11 VP.n36 VP.n0 161.3
R12 VP.n35 VP.n34 161.3
R13 VP.n33 VP.n1 161.3
R14 VP.n32 VP.n31 161.3
R15 VP.n30 VP.n2 161.3
R16 VP.n28 VP.n27 161.3
R17 VP.n26 VP.n3 161.3
R18 VP.n25 VP.n24 161.3
R19 VP.n23 VP.n4 161.3
R20 VP.n22 VP.n21 161.3
R21 VP.n20 VP.n5 98.0336
R22 VP.n38 VP.n37 98.0336
R23 VP.n19 VP.n18 98.0336
R24 VP.n10 VP.n9 59.258
R25 VP.n20 VP.n19 52.3291
R26 VP.n24 VP.n23 40.979
R27 VP.n35 VP.n1 40.979
R28 VP.n16 VP.n7 40.979
R29 VP.n24 VP.n3 40.0078
R30 VP.n31 VP.n1 40.0078
R31 VP.n12 VP.n7 40.0078
R32 VP.n23 VP.n22 24.4675
R33 VP.n28 VP.n3 24.4675
R34 VP.n31 VP.n30 24.4675
R35 VP.n36 VP.n35 24.4675
R36 VP.n17 VP.n16 24.4675
R37 VP.n12 VP.n11 24.4675
R38 VP.n22 VP.n5 12.7233
R39 VP.n37 VP.n36 12.7233
R40 VP.n18 VP.n17 12.7233
R41 VP.n29 VP.n28 12.234
R42 VP.n30 VP.n29 12.234
R43 VP.n11 VP.n10 12.234
R44 VP.n9 VP.n8 9.6787
R45 VP.n19 VP.n6 0.278367
R46 VP.n21 VP.n20 0.278367
R47 VP.n38 VP.n0 0.278367
R48 VP.n13 VP.n8 0.189894
R49 VP.n14 VP.n13 0.189894
R50 VP.n15 VP.n14 0.189894
R51 VP.n15 VP.n6 0.189894
R52 VP.n21 VP.n4 0.189894
R53 VP.n25 VP.n4 0.189894
R54 VP.n26 VP.n25 0.189894
R55 VP.n27 VP.n26 0.189894
R56 VP.n27 VP.n2 0.189894
R57 VP.n32 VP.n2 0.189894
R58 VP.n33 VP.n32 0.189894
R59 VP.n34 VP.n33 0.189894
R60 VP.n34 VP.n0 0.189894
R61 VP VP.n38 0.153454
R62 VDD1 VDD1.t3 64.6654
R63 VDD1.n1 VDD1.t2 64.5517
R64 VDD1.n1 VDD1.n0 62.4294
R65 VDD1.n3 VDD1.n2 61.9448
R66 VDD1.n3 VDD1.n1 48.8349
R67 VDD1.n2 VDD1.t4 1.03987
R68 VDD1.n2 VDD1.t5 1.03987
R69 VDD1.n0 VDD1.t1 1.03987
R70 VDD1.n0 VDD1.t0 1.03987
R71 VDD1 VDD1.n3 0.483259
R72 VTAIL.n7 VTAIL.t3 46.3055
R73 VTAIL.n11 VTAIL.t2 46.3054
R74 VTAIL.n2 VTAIL.t10 46.3054
R75 VTAIL.n10 VTAIL.t9 46.3054
R76 VTAIL.n9 VTAIL.n8 45.2662
R77 VTAIL.n6 VTAIL.n5 45.2662
R78 VTAIL.n1 VTAIL.n0 45.265
R79 VTAIL.n4 VTAIL.n3 45.265
R80 VTAIL.n6 VTAIL.n4 33.1169
R81 VTAIL.n11 VTAIL.n10 30.9531
R82 VTAIL.n7 VTAIL.n6 2.16429
R83 VTAIL.n10 VTAIL.n9 2.16429
R84 VTAIL.n4 VTAIL.n2 2.16429
R85 VTAIL VTAIL.n11 1.56516
R86 VTAIL.n9 VTAIL.n7 1.55222
R87 VTAIL.n2 VTAIL.n1 1.55222
R88 VTAIL.n0 VTAIL.t5 1.03987
R89 VTAIL.n0 VTAIL.t4 1.03987
R90 VTAIL.n3 VTAIL.t6 1.03987
R91 VTAIL.n3 VTAIL.t11 1.03987
R92 VTAIL.n8 VTAIL.t7 1.03987
R93 VTAIL.n8 VTAIL.t8 1.03987
R94 VTAIL.n5 VTAIL.t1 1.03987
R95 VTAIL.n5 VTAIL.t0 1.03987
R96 VTAIL VTAIL.n1 0.599638
R97 B.n982 B.n981 585
R98 B.n408 B.n137 585
R99 B.n407 B.n406 585
R100 B.n405 B.n404 585
R101 B.n403 B.n402 585
R102 B.n401 B.n400 585
R103 B.n399 B.n398 585
R104 B.n397 B.n396 585
R105 B.n395 B.n394 585
R106 B.n393 B.n392 585
R107 B.n391 B.n390 585
R108 B.n389 B.n388 585
R109 B.n387 B.n386 585
R110 B.n385 B.n384 585
R111 B.n383 B.n382 585
R112 B.n381 B.n380 585
R113 B.n379 B.n378 585
R114 B.n377 B.n376 585
R115 B.n375 B.n374 585
R116 B.n373 B.n372 585
R117 B.n371 B.n370 585
R118 B.n369 B.n368 585
R119 B.n367 B.n366 585
R120 B.n365 B.n364 585
R121 B.n363 B.n362 585
R122 B.n361 B.n360 585
R123 B.n359 B.n358 585
R124 B.n357 B.n356 585
R125 B.n355 B.n354 585
R126 B.n353 B.n352 585
R127 B.n351 B.n350 585
R128 B.n349 B.n348 585
R129 B.n347 B.n346 585
R130 B.n345 B.n344 585
R131 B.n343 B.n342 585
R132 B.n341 B.n340 585
R133 B.n339 B.n338 585
R134 B.n337 B.n336 585
R135 B.n335 B.n334 585
R136 B.n333 B.n332 585
R137 B.n331 B.n330 585
R138 B.n329 B.n328 585
R139 B.n327 B.n326 585
R140 B.n325 B.n324 585
R141 B.n323 B.n322 585
R142 B.n321 B.n320 585
R143 B.n319 B.n318 585
R144 B.n317 B.n316 585
R145 B.n315 B.n314 585
R146 B.n313 B.n312 585
R147 B.n311 B.n310 585
R148 B.n309 B.n308 585
R149 B.n307 B.n306 585
R150 B.n305 B.n304 585
R151 B.n303 B.n302 585
R152 B.n301 B.n300 585
R153 B.n299 B.n298 585
R154 B.n297 B.n296 585
R155 B.n295 B.n294 585
R156 B.n293 B.n292 585
R157 B.n291 B.n290 585
R158 B.n289 B.n288 585
R159 B.n287 B.n286 585
R160 B.n285 B.n284 585
R161 B.n283 B.n282 585
R162 B.n281 B.n280 585
R163 B.n279 B.n278 585
R164 B.n277 B.n276 585
R165 B.n275 B.n274 585
R166 B.n273 B.n272 585
R167 B.n271 B.n270 585
R168 B.n269 B.n268 585
R169 B.n267 B.n266 585
R170 B.n265 B.n264 585
R171 B.n263 B.n262 585
R172 B.n261 B.n260 585
R173 B.n259 B.n258 585
R174 B.n257 B.n256 585
R175 B.n255 B.n254 585
R176 B.n253 B.n252 585
R177 B.n251 B.n250 585
R178 B.n249 B.n248 585
R179 B.n247 B.n246 585
R180 B.n245 B.n244 585
R181 B.n243 B.n242 585
R182 B.n241 B.n240 585
R183 B.n239 B.n238 585
R184 B.n237 B.n236 585
R185 B.n235 B.n234 585
R186 B.n233 B.n232 585
R187 B.n231 B.n230 585
R188 B.n229 B.n228 585
R189 B.n227 B.n226 585
R190 B.n225 B.n224 585
R191 B.n223 B.n222 585
R192 B.n221 B.n220 585
R193 B.n219 B.n218 585
R194 B.n217 B.n216 585
R195 B.n215 B.n214 585
R196 B.n213 B.n212 585
R197 B.n211 B.n210 585
R198 B.n209 B.n208 585
R199 B.n207 B.n206 585
R200 B.n205 B.n204 585
R201 B.n203 B.n202 585
R202 B.n201 B.n200 585
R203 B.n199 B.n198 585
R204 B.n197 B.n196 585
R205 B.n195 B.n194 585
R206 B.n193 B.n192 585
R207 B.n191 B.n190 585
R208 B.n189 B.n188 585
R209 B.n187 B.n186 585
R210 B.n185 B.n184 585
R211 B.n183 B.n182 585
R212 B.n181 B.n180 585
R213 B.n179 B.n178 585
R214 B.n177 B.n176 585
R215 B.n175 B.n174 585
R216 B.n173 B.n172 585
R217 B.n171 B.n170 585
R218 B.n169 B.n168 585
R219 B.n167 B.n166 585
R220 B.n165 B.n164 585
R221 B.n163 B.n162 585
R222 B.n161 B.n160 585
R223 B.n159 B.n158 585
R224 B.n157 B.n156 585
R225 B.n155 B.n154 585
R226 B.n153 B.n152 585
R227 B.n151 B.n150 585
R228 B.n149 B.n148 585
R229 B.n147 B.n146 585
R230 B.n145 B.n144 585
R231 B.n980 B.n70 585
R232 B.n985 B.n70 585
R233 B.n979 B.n69 585
R234 B.n986 B.n69 585
R235 B.n978 B.n977 585
R236 B.n977 B.n65 585
R237 B.n976 B.n64 585
R238 B.n992 B.n64 585
R239 B.n975 B.n63 585
R240 B.n993 B.n63 585
R241 B.n974 B.n62 585
R242 B.n994 B.n62 585
R243 B.n973 B.n972 585
R244 B.n972 B.n61 585
R245 B.n971 B.n57 585
R246 B.n1000 B.n57 585
R247 B.n970 B.n56 585
R248 B.n1001 B.n56 585
R249 B.n969 B.n55 585
R250 B.n1002 B.n55 585
R251 B.n968 B.n967 585
R252 B.n967 B.n51 585
R253 B.n966 B.n50 585
R254 B.n1008 B.n50 585
R255 B.n965 B.n49 585
R256 B.n1009 B.n49 585
R257 B.n964 B.n48 585
R258 B.n1010 B.n48 585
R259 B.n963 B.n962 585
R260 B.n962 B.n44 585
R261 B.n961 B.n43 585
R262 B.n1016 B.n43 585
R263 B.n960 B.n42 585
R264 B.n1017 B.n42 585
R265 B.n959 B.n41 585
R266 B.n1018 B.n41 585
R267 B.n958 B.n957 585
R268 B.n957 B.n37 585
R269 B.n956 B.n36 585
R270 B.n1024 B.n36 585
R271 B.n955 B.n35 585
R272 B.n1025 B.n35 585
R273 B.n954 B.n34 585
R274 B.n1026 B.n34 585
R275 B.n953 B.n952 585
R276 B.n952 B.n30 585
R277 B.n951 B.n29 585
R278 B.n1032 B.n29 585
R279 B.n950 B.n28 585
R280 B.n1033 B.n28 585
R281 B.n949 B.n27 585
R282 B.n1034 B.n27 585
R283 B.n948 B.n947 585
R284 B.n947 B.n23 585
R285 B.n946 B.n22 585
R286 B.n1040 B.n22 585
R287 B.n945 B.n21 585
R288 B.n1041 B.n21 585
R289 B.n944 B.n20 585
R290 B.n1042 B.n20 585
R291 B.n943 B.n942 585
R292 B.n942 B.n16 585
R293 B.n941 B.n15 585
R294 B.n1048 B.n15 585
R295 B.n940 B.n14 585
R296 B.n1049 B.n14 585
R297 B.n939 B.n13 585
R298 B.n1050 B.n13 585
R299 B.n938 B.n937 585
R300 B.n937 B.n12 585
R301 B.n936 B.n935 585
R302 B.n936 B.n8 585
R303 B.n934 B.n7 585
R304 B.n1057 B.n7 585
R305 B.n933 B.n6 585
R306 B.n1058 B.n6 585
R307 B.n932 B.n5 585
R308 B.n1059 B.n5 585
R309 B.n931 B.n930 585
R310 B.n930 B.n4 585
R311 B.n929 B.n409 585
R312 B.n929 B.n928 585
R313 B.n919 B.n410 585
R314 B.n411 B.n410 585
R315 B.n921 B.n920 585
R316 B.n922 B.n921 585
R317 B.n918 B.n415 585
R318 B.n419 B.n415 585
R319 B.n917 B.n916 585
R320 B.n916 B.n915 585
R321 B.n417 B.n416 585
R322 B.n418 B.n417 585
R323 B.n908 B.n907 585
R324 B.n909 B.n908 585
R325 B.n906 B.n424 585
R326 B.n424 B.n423 585
R327 B.n905 B.n904 585
R328 B.n904 B.n903 585
R329 B.n426 B.n425 585
R330 B.n427 B.n426 585
R331 B.n896 B.n895 585
R332 B.n897 B.n896 585
R333 B.n894 B.n431 585
R334 B.n435 B.n431 585
R335 B.n893 B.n892 585
R336 B.n892 B.n891 585
R337 B.n433 B.n432 585
R338 B.n434 B.n433 585
R339 B.n884 B.n883 585
R340 B.n885 B.n884 585
R341 B.n882 B.n440 585
R342 B.n440 B.n439 585
R343 B.n881 B.n880 585
R344 B.n880 B.n879 585
R345 B.n442 B.n441 585
R346 B.n443 B.n442 585
R347 B.n872 B.n871 585
R348 B.n873 B.n872 585
R349 B.n870 B.n448 585
R350 B.n448 B.n447 585
R351 B.n869 B.n868 585
R352 B.n868 B.n867 585
R353 B.n450 B.n449 585
R354 B.n451 B.n450 585
R355 B.n860 B.n859 585
R356 B.n861 B.n860 585
R357 B.n858 B.n456 585
R358 B.n456 B.n455 585
R359 B.n857 B.n856 585
R360 B.n856 B.n855 585
R361 B.n458 B.n457 585
R362 B.n459 B.n458 585
R363 B.n848 B.n847 585
R364 B.n849 B.n848 585
R365 B.n846 B.n464 585
R366 B.n464 B.n463 585
R367 B.n845 B.n844 585
R368 B.n844 B.n843 585
R369 B.n466 B.n465 585
R370 B.n836 B.n466 585
R371 B.n835 B.n834 585
R372 B.n837 B.n835 585
R373 B.n833 B.n471 585
R374 B.n471 B.n470 585
R375 B.n832 B.n831 585
R376 B.n831 B.n830 585
R377 B.n473 B.n472 585
R378 B.n474 B.n473 585
R379 B.n823 B.n822 585
R380 B.n824 B.n823 585
R381 B.n821 B.n479 585
R382 B.n479 B.n478 585
R383 B.n816 B.n815 585
R384 B.n814 B.n548 585
R385 B.n813 B.n547 585
R386 B.n818 B.n547 585
R387 B.n812 B.n811 585
R388 B.n810 B.n809 585
R389 B.n808 B.n807 585
R390 B.n806 B.n805 585
R391 B.n804 B.n803 585
R392 B.n802 B.n801 585
R393 B.n800 B.n799 585
R394 B.n798 B.n797 585
R395 B.n796 B.n795 585
R396 B.n794 B.n793 585
R397 B.n792 B.n791 585
R398 B.n790 B.n789 585
R399 B.n788 B.n787 585
R400 B.n786 B.n785 585
R401 B.n784 B.n783 585
R402 B.n782 B.n781 585
R403 B.n780 B.n779 585
R404 B.n778 B.n777 585
R405 B.n776 B.n775 585
R406 B.n774 B.n773 585
R407 B.n772 B.n771 585
R408 B.n770 B.n769 585
R409 B.n768 B.n767 585
R410 B.n766 B.n765 585
R411 B.n764 B.n763 585
R412 B.n762 B.n761 585
R413 B.n760 B.n759 585
R414 B.n758 B.n757 585
R415 B.n756 B.n755 585
R416 B.n754 B.n753 585
R417 B.n752 B.n751 585
R418 B.n750 B.n749 585
R419 B.n748 B.n747 585
R420 B.n746 B.n745 585
R421 B.n744 B.n743 585
R422 B.n742 B.n741 585
R423 B.n740 B.n739 585
R424 B.n738 B.n737 585
R425 B.n736 B.n735 585
R426 B.n734 B.n733 585
R427 B.n732 B.n731 585
R428 B.n730 B.n729 585
R429 B.n728 B.n727 585
R430 B.n726 B.n725 585
R431 B.n724 B.n723 585
R432 B.n722 B.n721 585
R433 B.n720 B.n719 585
R434 B.n718 B.n717 585
R435 B.n716 B.n715 585
R436 B.n714 B.n713 585
R437 B.n712 B.n711 585
R438 B.n710 B.n709 585
R439 B.n708 B.n707 585
R440 B.n706 B.n705 585
R441 B.n704 B.n703 585
R442 B.n702 B.n701 585
R443 B.n700 B.n699 585
R444 B.n698 B.n697 585
R445 B.n696 B.n695 585
R446 B.n693 B.n692 585
R447 B.n691 B.n690 585
R448 B.n689 B.n688 585
R449 B.n687 B.n686 585
R450 B.n685 B.n684 585
R451 B.n683 B.n682 585
R452 B.n681 B.n680 585
R453 B.n679 B.n678 585
R454 B.n677 B.n676 585
R455 B.n675 B.n674 585
R456 B.n672 B.n671 585
R457 B.n670 B.n669 585
R458 B.n668 B.n667 585
R459 B.n666 B.n665 585
R460 B.n664 B.n663 585
R461 B.n662 B.n661 585
R462 B.n660 B.n659 585
R463 B.n658 B.n657 585
R464 B.n656 B.n655 585
R465 B.n654 B.n653 585
R466 B.n652 B.n651 585
R467 B.n650 B.n649 585
R468 B.n648 B.n647 585
R469 B.n646 B.n645 585
R470 B.n644 B.n643 585
R471 B.n642 B.n641 585
R472 B.n640 B.n639 585
R473 B.n638 B.n637 585
R474 B.n636 B.n635 585
R475 B.n634 B.n633 585
R476 B.n632 B.n631 585
R477 B.n630 B.n629 585
R478 B.n628 B.n627 585
R479 B.n626 B.n625 585
R480 B.n624 B.n623 585
R481 B.n622 B.n621 585
R482 B.n620 B.n619 585
R483 B.n618 B.n617 585
R484 B.n616 B.n615 585
R485 B.n614 B.n613 585
R486 B.n612 B.n611 585
R487 B.n610 B.n609 585
R488 B.n608 B.n607 585
R489 B.n606 B.n605 585
R490 B.n604 B.n603 585
R491 B.n602 B.n601 585
R492 B.n600 B.n599 585
R493 B.n598 B.n597 585
R494 B.n596 B.n595 585
R495 B.n594 B.n593 585
R496 B.n592 B.n591 585
R497 B.n590 B.n589 585
R498 B.n588 B.n587 585
R499 B.n586 B.n585 585
R500 B.n584 B.n583 585
R501 B.n582 B.n581 585
R502 B.n580 B.n579 585
R503 B.n578 B.n577 585
R504 B.n576 B.n575 585
R505 B.n574 B.n573 585
R506 B.n572 B.n571 585
R507 B.n570 B.n569 585
R508 B.n568 B.n567 585
R509 B.n566 B.n565 585
R510 B.n564 B.n563 585
R511 B.n562 B.n561 585
R512 B.n560 B.n559 585
R513 B.n558 B.n557 585
R514 B.n556 B.n555 585
R515 B.n554 B.n553 585
R516 B.n481 B.n480 585
R517 B.n820 B.n819 585
R518 B.n819 B.n818 585
R519 B.n477 B.n476 585
R520 B.n478 B.n477 585
R521 B.n826 B.n825 585
R522 B.n825 B.n824 585
R523 B.n827 B.n475 585
R524 B.n475 B.n474 585
R525 B.n829 B.n828 585
R526 B.n830 B.n829 585
R527 B.n469 B.n468 585
R528 B.n470 B.n469 585
R529 B.n839 B.n838 585
R530 B.n838 B.n837 585
R531 B.n840 B.n467 585
R532 B.n836 B.n467 585
R533 B.n842 B.n841 585
R534 B.n843 B.n842 585
R535 B.n462 B.n461 585
R536 B.n463 B.n462 585
R537 B.n851 B.n850 585
R538 B.n850 B.n849 585
R539 B.n852 B.n460 585
R540 B.n460 B.n459 585
R541 B.n854 B.n853 585
R542 B.n855 B.n854 585
R543 B.n454 B.n453 585
R544 B.n455 B.n454 585
R545 B.n863 B.n862 585
R546 B.n862 B.n861 585
R547 B.n864 B.n452 585
R548 B.n452 B.n451 585
R549 B.n866 B.n865 585
R550 B.n867 B.n866 585
R551 B.n446 B.n445 585
R552 B.n447 B.n446 585
R553 B.n875 B.n874 585
R554 B.n874 B.n873 585
R555 B.n876 B.n444 585
R556 B.n444 B.n443 585
R557 B.n878 B.n877 585
R558 B.n879 B.n878 585
R559 B.n438 B.n437 585
R560 B.n439 B.n438 585
R561 B.n887 B.n886 585
R562 B.n886 B.n885 585
R563 B.n888 B.n436 585
R564 B.n436 B.n434 585
R565 B.n890 B.n889 585
R566 B.n891 B.n890 585
R567 B.n430 B.n429 585
R568 B.n435 B.n430 585
R569 B.n899 B.n898 585
R570 B.n898 B.n897 585
R571 B.n900 B.n428 585
R572 B.n428 B.n427 585
R573 B.n902 B.n901 585
R574 B.n903 B.n902 585
R575 B.n422 B.n421 585
R576 B.n423 B.n422 585
R577 B.n911 B.n910 585
R578 B.n910 B.n909 585
R579 B.n912 B.n420 585
R580 B.n420 B.n418 585
R581 B.n914 B.n913 585
R582 B.n915 B.n914 585
R583 B.n414 B.n413 585
R584 B.n419 B.n414 585
R585 B.n924 B.n923 585
R586 B.n923 B.n922 585
R587 B.n925 B.n412 585
R588 B.n412 B.n411 585
R589 B.n927 B.n926 585
R590 B.n928 B.n927 585
R591 B.n3 B.n0 585
R592 B.n4 B.n3 585
R593 B.n1056 B.n1 585
R594 B.n1057 B.n1056 585
R595 B.n1055 B.n1054 585
R596 B.n1055 B.n8 585
R597 B.n1053 B.n9 585
R598 B.n12 B.n9 585
R599 B.n1052 B.n1051 585
R600 B.n1051 B.n1050 585
R601 B.n11 B.n10 585
R602 B.n1049 B.n11 585
R603 B.n1047 B.n1046 585
R604 B.n1048 B.n1047 585
R605 B.n1045 B.n17 585
R606 B.n17 B.n16 585
R607 B.n1044 B.n1043 585
R608 B.n1043 B.n1042 585
R609 B.n19 B.n18 585
R610 B.n1041 B.n19 585
R611 B.n1039 B.n1038 585
R612 B.n1040 B.n1039 585
R613 B.n1037 B.n24 585
R614 B.n24 B.n23 585
R615 B.n1036 B.n1035 585
R616 B.n1035 B.n1034 585
R617 B.n26 B.n25 585
R618 B.n1033 B.n26 585
R619 B.n1031 B.n1030 585
R620 B.n1032 B.n1031 585
R621 B.n1029 B.n31 585
R622 B.n31 B.n30 585
R623 B.n1028 B.n1027 585
R624 B.n1027 B.n1026 585
R625 B.n33 B.n32 585
R626 B.n1025 B.n33 585
R627 B.n1023 B.n1022 585
R628 B.n1024 B.n1023 585
R629 B.n1021 B.n38 585
R630 B.n38 B.n37 585
R631 B.n1020 B.n1019 585
R632 B.n1019 B.n1018 585
R633 B.n40 B.n39 585
R634 B.n1017 B.n40 585
R635 B.n1015 B.n1014 585
R636 B.n1016 B.n1015 585
R637 B.n1013 B.n45 585
R638 B.n45 B.n44 585
R639 B.n1012 B.n1011 585
R640 B.n1011 B.n1010 585
R641 B.n47 B.n46 585
R642 B.n1009 B.n47 585
R643 B.n1007 B.n1006 585
R644 B.n1008 B.n1007 585
R645 B.n1005 B.n52 585
R646 B.n52 B.n51 585
R647 B.n1004 B.n1003 585
R648 B.n1003 B.n1002 585
R649 B.n54 B.n53 585
R650 B.n1001 B.n54 585
R651 B.n999 B.n998 585
R652 B.n1000 B.n999 585
R653 B.n997 B.n58 585
R654 B.n61 B.n58 585
R655 B.n996 B.n995 585
R656 B.n995 B.n994 585
R657 B.n60 B.n59 585
R658 B.n993 B.n60 585
R659 B.n991 B.n990 585
R660 B.n992 B.n991 585
R661 B.n989 B.n66 585
R662 B.n66 B.n65 585
R663 B.n988 B.n987 585
R664 B.n987 B.n986 585
R665 B.n68 B.n67 585
R666 B.n985 B.n68 585
R667 B.n1060 B.n1059 585
R668 B.n1058 B.n2 585
R669 B.n144 B.n68 545.355
R670 B.n982 B.n70 545.355
R671 B.n819 B.n479 545.355
R672 B.n816 B.n477 545.355
R673 B.n141 B.t13 417.909
R674 B.n138 B.t17 417.909
R675 B.n551 B.t10 417.909
R676 B.n549 B.t6 417.909
R677 B.n984 B.n983 256.663
R678 B.n984 B.n136 256.663
R679 B.n984 B.n135 256.663
R680 B.n984 B.n134 256.663
R681 B.n984 B.n133 256.663
R682 B.n984 B.n132 256.663
R683 B.n984 B.n131 256.663
R684 B.n984 B.n130 256.663
R685 B.n984 B.n129 256.663
R686 B.n984 B.n128 256.663
R687 B.n984 B.n127 256.663
R688 B.n984 B.n126 256.663
R689 B.n984 B.n125 256.663
R690 B.n984 B.n124 256.663
R691 B.n984 B.n123 256.663
R692 B.n984 B.n122 256.663
R693 B.n984 B.n121 256.663
R694 B.n984 B.n120 256.663
R695 B.n984 B.n119 256.663
R696 B.n984 B.n118 256.663
R697 B.n984 B.n117 256.663
R698 B.n984 B.n116 256.663
R699 B.n984 B.n115 256.663
R700 B.n984 B.n114 256.663
R701 B.n984 B.n113 256.663
R702 B.n984 B.n112 256.663
R703 B.n984 B.n111 256.663
R704 B.n984 B.n110 256.663
R705 B.n984 B.n109 256.663
R706 B.n984 B.n108 256.663
R707 B.n984 B.n107 256.663
R708 B.n984 B.n106 256.663
R709 B.n984 B.n105 256.663
R710 B.n984 B.n104 256.663
R711 B.n984 B.n103 256.663
R712 B.n984 B.n102 256.663
R713 B.n984 B.n101 256.663
R714 B.n984 B.n100 256.663
R715 B.n984 B.n99 256.663
R716 B.n984 B.n98 256.663
R717 B.n984 B.n97 256.663
R718 B.n984 B.n96 256.663
R719 B.n984 B.n95 256.663
R720 B.n984 B.n94 256.663
R721 B.n984 B.n93 256.663
R722 B.n984 B.n92 256.663
R723 B.n984 B.n91 256.663
R724 B.n984 B.n90 256.663
R725 B.n984 B.n89 256.663
R726 B.n984 B.n88 256.663
R727 B.n984 B.n87 256.663
R728 B.n984 B.n86 256.663
R729 B.n984 B.n85 256.663
R730 B.n984 B.n84 256.663
R731 B.n984 B.n83 256.663
R732 B.n984 B.n82 256.663
R733 B.n984 B.n81 256.663
R734 B.n984 B.n80 256.663
R735 B.n984 B.n79 256.663
R736 B.n984 B.n78 256.663
R737 B.n984 B.n77 256.663
R738 B.n984 B.n76 256.663
R739 B.n984 B.n75 256.663
R740 B.n984 B.n74 256.663
R741 B.n984 B.n73 256.663
R742 B.n984 B.n72 256.663
R743 B.n984 B.n71 256.663
R744 B.n818 B.n817 256.663
R745 B.n818 B.n482 256.663
R746 B.n818 B.n483 256.663
R747 B.n818 B.n484 256.663
R748 B.n818 B.n485 256.663
R749 B.n818 B.n486 256.663
R750 B.n818 B.n487 256.663
R751 B.n818 B.n488 256.663
R752 B.n818 B.n489 256.663
R753 B.n818 B.n490 256.663
R754 B.n818 B.n491 256.663
R755 B.n818 B.n492 256.663
R756 B.n818 B.n493 256.663
R757 B.n818 B.n494 256.663
R758 B.n818 B.n495 256.663
R759 B.n818 B.n496 256.663
R760 B.n818 B.n497 256.663
R761 B.n818 B.n498 256.663
R762 B.n818 B.n499 256.663
R763 B.n818 B.n500 256.663
R764 B.n818 B.n501 256.663
R765 B.n818 B.n502 256.663
R766 B.n818 B.n503 256.663
R767 B.n818 B.n504 256.663
R768 B.n818 B.n505 256.663
R769 B.n818 B.n506 256.663
R770 B.n818 B.n507 256.663
R771 B.n818 B.n508 256.663
R772 B.n818 B.n509 256.663
R773 B.n818 B.n510 256.663
R774 B.n818 B.n511 256.663
R775 B.n818 B.n512 256.663
R776 B.n818 B.n513 256.663
R777 B.n818 B.n514 256.663
R778 B.n818 B.n515 256.663
R779 B.n818 B.n516 256.663
R780 B.n818 B.n517 256.663
R781 B.n818 B.n518 256.663
R782 B.n818 B.n519 256.663
R783 B.n818 B.n520 256.663
R784 B.n818 B.n521 256.663
R785 B.n818 B.n522 256.663
R786 B.n818 B.n523 256.663
R787 B.n818 B.n524 256.663
R788 B.n818 B.n525 256.663
R789 B.n818 B.n526 256.663
R790 B.n818 B.n527 256.663
R791 B.n818 B.n528 256.663
R792 B.n818 B.n529 256.663
R793 B.n818 B.n530 256.663
R794 B.n818 B.n531 256.663
R795 B.n818 B.n532 256.663
R796 B.n818 B.n533 256.663
R797 B.n818 B.n534 256.663
R798 B.n818 B.n535 256.663
R799 B.n818 B.n536 256.663
R800 B.n818 B.n537 256.663
R801 B.n818 B.n538 256.663
R802 B.n818 B.n539 256.663
R803 B.n818 B.n540 256.663
R804 B.n818 B.n541 256.663
R805 B.n818 B.n542 256.663
R806 B.n818 B.n543 256.663
R807 B.n818 B.n544 256.663
R808 B.n818 B.n545 256.663
R809 B.n818 B.n546 256.663
R810 B.n1062 B.n1061 256.663
R811 B.n148 B.n147 163.367
R812 B.n152 B.n151 163.367
R813 B.n156 B.n155 163.367
R814 B.n160 B.n159 163.367
R815 B.n164 B.n163 163.367
R816 B.n168 B.n167 163.367
R817 B.n172 B.n171 163.367
R818 B.n176 B.n175 163.367
R819 B.n180 B.n179 163.367
R820 B.n184 B.n183 163.367
R821 B.n188 B.n187 163.367
R822 B.n192 B.n191 163.367
R823 B.n196 B.n195 163.367
R824 B.n200 B.n199 163.367
R825 B.n204 B.n203 163.367
R826 B.n208 B.n207 163.367
R827 B.n212 B.n211 163.367
R828 B.n216 B.n215 163.367
R829 B.n220 B.n219 163.367
R830 B.n224 B.n223 163.367
R831 B.n228 B.n227 163.367
R832 B.n232 B.n231 163.367
R833 B.n236 B.n235 163.367
R834 B.n240 B.n239 163.367
R835 B.n244 B.n243 163.367
R836 B.n248 B.n247 163.367
R837 B.n252 B.n251 163.367
R838 B.n256 B.n255 163.367
R839 B.n260 B.n259 163.367
R840 B.n264 B.n263 163.367
R841 B.n268 B.n267 163.367
R842 B.n272 B.n271 163.367
R843 B.n276 B.n275 163.367
R844 B.n280 B.n279 163.367
R845 B.n284 B.n283 163.367
R846 B.n288 B.n287 163.367
R847 B.n292 B.n291 163.367
R848 B.n296 B.n295 163.367
R849 B.n300 B.n299 163.367
R850 B.n304 B.n303 163.367
R851 B.n308 B.n307 163.367
R852 B.n312 B.n311 163.367
R853 B.n316 B.n315 163.367
R854 B.n320 B.n319 163.367
R855 B.n324 B.n323 163.367
R856 B.n328 B.n327 163.367
R857 B.n332 B.n331 163.367
R858 B.n336 B.n335 163.367
R859 B.n340 B.n339 163.367
R860 B.n344 B.n343 163.367
R861 B.n348 B.n347 163.367
R862 B.n352 B.n351 163.367
R863 B.n356 B.n355 163.367
R864 B.n360 B.n359 163.367
R865 B.n364 B.n363 163.367
R866 B.n368 B.n367 163.367
R867 B.n372 B.n371 163.367
R868 B.n376 B.n375 163.367
R869 B.n380 B.n379 163.367
R870 B.n384 B.n383 163.367
R871 B.n388 B.n387 163.367
R872 B.n392 B.n391 163.367
R873 B.n396 B.n395 163.367
R874 B.n400 B.n399 163.367
R875 B.n404 B.n403 163.367
R876 B.n406 B.n137 163.367
R877 B.n823 B.n479 163.367
R878 B.n823 B.n473 163.367
R879 B.n831 B.n473 163.367
R880 B.n831 B.n471 163.367
R881 B.n835 B.n471 163.367
R882 B.n835 B.n466 163.367
R883 B.n844 B.n466 163.367
R884 B.n844 B.n464 163.367
R885 B.n848 B.n464 163.367
R886 B.n848 B.n458 163.367
R887 B.n856 B.n458 163.367
R888 B.n856 B.n456 163.367
R889 B.n860 B.n456 163.367
R890 B.n860 B.n450 163.367
R891 B.n868 B.n450 163.367
R892 B.n868 B.n448 163.367
R893 B.n872 B.n448 163.367
R894 B.n872 B.n442 163.367
R895 B.n880 B.n442 163.367
R896 B.n880 B.n440 163.367
R897 B.n884 B.n440 163.367
R898 B.n884 B.n433 163.367
R899 B.n892 B.n433 163.367
R900 B.n892 B.n431 163.367
R901 B.n896 B.n431 163.367
R902 B.n896 B.n426 163.367
R903 B.n904 B.n426 163.367
R904 B.n904 B.n424 163.367
R905 B.n908 B.n424 163.367
R906 B.n908 B.n417 163.367
R907 B.n916 B.n417 163.367
R908 B.n916 B.n415 163.367
R909 B.n921 B.n415 163.367
R910 B.n921 B.n410 163.367
R911 B.n929 B.n410 163.367
R912 B.n930 B.n929 163.367
R913 B.n930 B.n5 163.367
R914 B.n6 B.n5 163.367
R915 B.n7 B.n6 163.367
R916 B.n936 B.n7 163.367
R917 B.n937 B.n936 163.367
R918 B.n937 B.n13 163.367
R919 B.n14 B.n13 163.367
R920 B.n15 B.n14 163.367
R921 B.n942 B.n15 163.367
R922 B.n942 B.n20 163.367
R923 B.n21 B.n20 163.367
R924 B.n22 B.n21 163.367
R925 B.n947 B.n22 163.367
R926 B.n947 B.n27 163.367
R927 B.n28 B.n27 163.367
R928 B.n29 B.n28 163.367
R929 B.n952 B.n29 163.367
R930 B.n952 B.n34 163.367
R931 B.n35 B.n34 163.367
R932 B.n36 B.n35 163.367
R933 B.n957 B.n36 163.367
R934 B.n957 B.n41 163.367
R935 B.n42 B.n41 163.367
R936 B.n43 B.n42 163.367
R937 B.n962 B.n43 163.367
R938 B.n962 B.n48 163.367
R939 B.n49 B.n48 163.367
R940 B.n50 B.n49 163.367
R941 B.n967 B.n50 163.367
R942 B.n967 B.n55 163.367
R943 B.n56 B.n55 163.367
R944 B.n57 B.n56 163.367
R945 B.n972 B.n57 163.367
R946 B.n972 B.n62 163.367
R947 B.n63 B.n62 163.367
R948 B.n64 B.n63 163.367
R949 B.n977 B.n64 163.367
R950 B.n977 B.n69 163.367
R951 B.n70 B.n69 163.367
R952 B.n548 B.n547 163.367
R953 B.n811 B.n547 163.367
R954 B.n809 B.n808 163.367
R955 B.n805 B.n804 163.367
R956 B.n801 B.n800 163.367
R957 B.n797 B.n796 163.367
R958 B.n793 B.n792 163.367
R959 B.n789 B.n788 163.367
R960 B.n785 B.n784 163.367
R961 B.n781 B.n780 163.367
R962 B.n777 B.n776 163.367
R963 B.n773 B.n772 163.367
R964 B.n769 B.n768 163.367
R965 B.n765 B.n764 163.367
R966 B.n761 B.n760 163.367
R967 B.n757 B.n756 163.367
R968 B.n753 B.n752 163.367
R969 B.n749 B.n748 163.367
R970 B.n745 B.n744 163.367
R971 B.n741 B.n740 163.367
R972 B.n737 B.n736 163.367
R973 B.n733 B.n732 163.367
R974 B.n729 B.n728 163.367
R975 B.n725 B.n724 163.367
R976 B.n721 B.n720 163.367
R977 B.n717 B.n716 163.367
R978 B.n713 B.n712 163.367
R979 B.n709 B.n708 163.367
R980 B.n705 B.n704 163.367
R981 B.n701 B.n700 163.367
R982 B.n697 B.n696 163.367
R983 B.n692 B.n691 163.367
R984 B.n688 B.n687 163.367
R985 B.n684 B.n683 163.367
R986 B.n680 B.n679 163.367
R987 B.n676 B.n675 163.367
R988 B.n671 B.n670 163.367
R989 B.n667 B.n666 163.367
R990 B.n663 B.n662 163.367
R991 B.n659 B.n658 163.367
R992 B.n655 B.n654 163.367
R993 B.n651 B.n650 163.367
R994 B.n647 B.n646 163.367
R995 B.n643 B.n642 163.367
R996 B.n639 B.n638 163.367
R997 B.n635 B.n634 163.367
R998 B.n631 B.n630 163.367
R999 B.n627 B.n626 163.367
R1000 B.n623 B.n622 163.367
R1001 B.n619 B.n618 163.367
R1002 B.n615 B.n614 163.367
R1003 B.n611 B.n610 163.367
R1004 B.n607 B.n606 163.367
R1005 B.n603 B.n602 163.367
R1006 B.n599 B.n598 163.367
R1007 B.n595 B.n594 163.367
R1008 B.n591 B.n590 163.367
R1009 B.n587 B.n586 163.367
R1010 B.n583 B.n582 163.367
R1011 B.n579 B.n578 163.367
R1012 B.n575 B.n574 163.367
R1013 B.n571 B.n570 163.367
R1014 B.n567 B.n566 163.367
R1015 B.n563 B.n562 163.367
R1016 B.n559 B.n558 163.367
R1017 B.n555 B.n554 163.367
R1018 B.n819 B.n481 163.367
R1019 B.n825 B.n477 163.367
R1020 B.n825 B.n475 163.367
R1021 B.n829 B.n475 163.367
R1022 B.n829 B.n469 163.367
R1023 B.n838 B.n469 163.367
R1024 B.n838 B.n467 163.367
R1025 B.n842 B.n467 163.367
R1026 B.n842 B.n462 163.367
R1027 B.n850 B.n462 163.367
R1028 B.n850 B.n460 163.367
R1029 B.n854 B.n460 163.367
R1030 B.n854 B.n454 163.367
R1031 B.n862 B.n454 163.367
R1032 B.n862 B.n452 163.367
R1033 B.n866 B.n452 163.367
R1034 B.n866 B.n446 163.367
R1035 B.n874 B.n446 163.367
R1036 B.n874 B.n444 163.367
R1037 B.n878 B.n444 163.367
R1038 B.n878 B.n438 163.367
R1039 B.n886 B.n438 163.367
R1040 B.n886 B.n436 163.367
R1041 B.n890 B.n436 163.367
R1042 B.n890 B.n430 163.367
R1043 B.n898 B.n430 163.367
R1044 B.n898 B.n428 163.367
R1045 B.n902 B.n428 163.367
R1046 B.n902 B.n422 163.367
R1047 B.n910 B.n422 163.367
R1048 B.n910 B.n420 163.367
R1049 B.n914 B.n420 163.367
R1050 B.n914 B.n414 163.367
R1051 B.n923 B.n414 163.367
R1052 B.n923 B.n412 163.367
R1053 B.n927 B.n412 163.367
R1054 B.n927 B.n3 163.367
R1055 B.n1060 B.n3 163.367
R1056 B.n1056 B.n2 163.367
R1057 B.n1056 B.n1055 163.367
R1058 B.n1055 B.n9 163.367
R1059 B.n1051 B.n9 163.367
R1060 B.n1051 B.n11 163.367
R1061 B.n1047 B.n11 163.367
R1062 B.n1047 B.n17 163.367
R1063 B.n1043 B.n17 163.367
R1064 B.n1043 B.n19 163.367
R1065 B.n1039 B.n19 163.367
R1066 B.n1039 B.n24 163.367
R1067 B.n1035 B.n24 163.367
R1068 B.n1035 B.n26 163.367
R1069 B.n1031 B.n26 163.367
R1070 B.n1031 B.n31 163.367
R1071 B.n1027 B.n31 163.367
R1072 B.n1027 B.n33 163.367
R1073 B.n1023 B.n33 163.367
R1074 B.n1023 B.n38 163.367
R1075 B.n1019 B.n38 163.367
R1076 B.n1019 B.n40 163.367
R1077 B.n1015 B.n40 163.367
R1078 B.n1015 B.n45 163.367
R1079 B.n1011 B.n45 163.367
R1080 B.n1011 B.n47 163.367
R1081 B.n1007 B.n47 163.367
R1082 B.n1007 B.n52 163.367
R1083 B.n1003 B.n52 163.367
R1084 B.n1003 B.n54 163.367
R1085 B.n999 B.n54 163.367
R1086 B.n999 B.n58 163.367
R1087 B.n995 B.n58 163.367
R1088 B.n995 B.n60 163.367
R1089 B.n991 B.n60 163.367
R1090 B.n991 B.n66 163.367
R1091 B.n987 B.n66 163.367
R1092 B.n987 B.n68 163.367
R1093 B.n138 B.t18 116.062
R1094 B.n551 B.t12 116.062
R1095 B.n141 B.t15 116.037
R1096 B.n549 B.t9 116.037
R1097 B.n144 B.n71 71.676
R1098 B.n148 B.n72 71.676
R1099 B.n152 B.n73 71.676
R1100 B.n156 B.n74 71.676
R1101 B.n160 B.n75 71.676
R1102 B.n164 B.n76 71.676
R1103 B.n168 B.n77 71.676
R1104 B.n172 B.n78 71.676
R1105 B.n176 B.n79 71.676
R1106 B.n180 B.n80 71.676
R1107 B.n184 B.n81 71.676
R1108 B.n188 B.n82 71.676
R1109 B.n192 B.n83 71.676
R1110 B.n196 B.n84 71.676
R1111 B.n200 B.n85 71.676
R1112 B.n204 B.n86 71.676
R1113 B.n208 B.n87 71.676
R1114 B.n212 B.n88 71.676
R1115 B.n216 B.n89 71.676
R1116 B.n220 B.n90 71.676
R1117 B.n224 B.n91 71.676
R1118 B.n228 B.n92 71.676
R1119 B.n232 B.n93 71.676
R1120 B.n236 B.n94 71.676
R1121 B.n240 B.n95 71.676
R1122 B.n244 B.n96 71.676
R1123 B.n248 B.n97 71.676
R1124 B.n252 B.n98 71.676
R1125 B.n256 B.n99 71.676
R1126 B.n260 B.n100 71.676
R1127 B.n264 B.n101 71.676
R1128 B.n268 B.n102 71.676
R1129 B.n272 B.n103 71.676
R1130 B.n276 B.n104 71.676
R1131 B.n280 B.n105 71.676
R1132 B.n284 B.n106 71.676
R1133 B.n288 B.n107 71.676
R1134 B.n292 B.n108 71.676
R1135 B.n296 B.n109 71.676
R1136 B.n300 B.n110 71.676
R1137 B.n304 B.n111 71.676
R1138 B.n308 B.n112 71.676
R1139 B.n312 B.n113 71.676
R1140 B.n316 B.n114 71.676
R1141 B.n320 B.n115 71.676
R1142 B.n324 B.n116 71.676
R1143 B.n328 B.n117 71.676
R1144 B.n332 B.n118 71.676
R1145 B.n336 B.n119 71.676
R1146 B.n340 B.n120 71.676
R1147 B.n344 B.n121 71.676
R1148 B.n348 B.n122 71.676
R1149 B.n352 B.n123 71.676
R1150 B.n356 B.n124 71.676
R1151 B.n360 B.n125 71.676
R1152 B.n364 B.n126 71.676
R1153 B.n368 B.n127 71.676
R1154 B.n372 B.n128 71.676
R1155 B.n376 B.n129 71.676
R1156 B.n380 B.n130 71.676
R1157 B.n384 B.n131 71.676
R1158 B.n388 B.n132 71.676
R1159 B.n392 B.n133 71.676
R1160 B.n396 B.n134 71.676
R1161 B.n400 B.n135 71.676
R1162 B.n404 B.n136 71.676
R1163 B.n983 B.n137 71.676
R1164 B.n983 B.n982 71.676
R1165 B.n406 B.n136 71.676
R1166 B.n403 B.n135 71.676
R1167 B.n399 B.n134 71.676
R1168 B.n395 B.n133 71.676
R1169 B.n391 B.n132 71.676
R1170 B.n387 B.n131 71.676
R1171 B.n383 B.n130 71.676
R1172 B.n379 B.n129 71.676
R1173 B.n375 B.n128 71.676
R1174 B.n371 B.n127 71.676
R1175 B.n367 B.n126 71.676
R1176 B.n363 B.n125 71.676
R1177 B.n359 B.n124 71.676
R1178 B.n355 B.n123 71.676
R1179 B.n351 B.n122 71.676
R1180 B.n347 B.n121 71.676
R1181 B.n343 B.n120 71.676
R1182 B.n339 B.n119 71.676
R1183 B.n335 B.n118 71.676
R1184 B.n331 B.n117 71.676
R1185 B.n327 B.n116 71.676
R1186 B.n323 B.n115 71.676
R1187 B.n319 B.n114 71.676
R1188 B.n315 B.n113 71.676
R1189 B.n311 B.n112 71.676
R1190 B.n307 B.n111 71.676
R1191 B.n303 B.n110 71.676
R1192 B.n299 B.n109 71.676
R1193 B.n295 B.n108 71.676
R1194 B.n291 B.n107 71.676
R1195 B.n287 B.n106 71.676
R1196 B.n283 B.n105 71.676
R1197 B.n279 B.n104 71.676
R1198 B.n275 B.n103 71.676
R1199 B.n271 B.n102 71.676
R1200 B.n267 B.n101 71.676
R1201 B.n263 B.n100 71.676
R1202 B.n259 B.n99 71.676
R1203 B.n255 B.n98 71.676
R1204 B.n251 B.n97 71.676
R1205 B.n247 B.n96 71.676
R1206 B.n243 B.n95 71.676
R1207 B.n239 B.n94 71.676
R1208 B.n235 B.n93 71.676
R1209 B.n231 B.n92 71.676
R1210 B.n227 B.n91 71.676
R1211 B.n223 B.n90 71.676
R1212 B.n219 B.n89 71.676
R1213 B.n215 B.n88 71.676
R1214 B.n211 B.n87 71.676
R1215 B.n207 B.n86 71.676
R1216 B.n203 B.n85 71.676
R1217 B.n199 B.n84 71.676
R1218 B.n195 B.n83 71.676
R1219 B.n191 B.n82 71.676
R1220 B.n187 B.n81 71.676
R1221 B.n183 B.n80 71.676
R1222 B.n179 B.n79 71.676
R1223 B.n175 B.n78 71.676
R1224 B.n171 B.n77 71.676
R1225 B.n167 B.n76 71.676
R1226 B.n163 B.n75 71.676
R1227 B.n159 B.n74 71.676
R1228 B.n155 B.n73 71.676
R1229 B.n151 B.n72 71.676
R1230 B.n147 B.n71 71.676
R1231 B.n817 B.n816 71.676
R1232 B.n811 B.n482 71.676
R1233 B.n808 B.n483 71.676
R1234 B.n804 B.n484 71.676
R1235 B.n800 B.n485 71.676
R1236 B.n796 B.n486 71.676
R1237 B.n792 B.n487 71.676
R1238 B.n788 B.n488 71.676
R1239 B.n784 B.n489 71.676
R1240 B.n780 B.n490 71.676
R1241 B.n776 B.n491 71.676
R1242 B.n772 B.n492 71.676
R1243 B.n768 B.n493 71.676
R1244 B.n764 B.n494 71.676
R1245 B.n760 B.n495 71.676
R1246 B.n756 B.n496 71.676
R1247 B.n752 B.n497 71.676
R1248 B.n748 B.n498 71.676
R1249 B.n744 B.n499 71.676
R1250 B.n740 B.n500 71.676
R1251 B.n736 B.n501 71.676
R1252 B.n732 B.n502 71.676
R1253 B.n728 B.n503 71.676
R1254 B.n724 B.n504 71.676
R1255 B.n720 B.n505 71.676
R1256 B.n716 B.n506 71.676
R1257 B.n712 B.n507 71.676
R1258 B.n708 B.n508 71.676
R1259 B.n704 B.n509 71.676
R1260 B.n700 B.n510 71.676
R1261 B.n696 B.n511 71.676
R1262 B.n691 B.n512 71.676
R1263 B.n687 B.n513 71.676
R1264 B.n683 B.n514 71.676
R1265 B.n679 B.n515 71.676
R1266 B.n675 B.n516 71.676
R1267 B.n670 B.n517 71.676
R1268 B.n666 B.n518 71.676
R1269 B.n662 B.n519 71.676
R1270 B.n658 B.n520 71.676
R1271 B.n654 B.n521 71.676
R1272 B.n650 B.n522 71.676
R1273 B.n646 B.n523 71.676
R1274 B.n642 B.n524 71.676
R1275 B.n638 B.n525 71.676
R1276 B.n634 B.n526 71.676
R1277 B.n630 B.n527 71.676
R1278 B.n626 B.n528 71.676
R1279 B.n622 B.n529 71.676
R1280 B.n618 B.n530 71.676
R1281 B.n614 B.n531 71.676
R1282 B.n610 B.n532 71.676
R1283 B.n606 B.n533 71.676
R1284 B.n602 B.n534 71.676
R1285 B.n598 B.n535 71.676
R1286 B.n594 B.n536 71.676
R1287 B.n590 B.n537 71.676
R1288 B.n586 B.n538 71.676
R1289 B.n582 B.n539 71.676
R1290 B.n578 B.n540 71.676
R1291 B.n574 B.n541 71.676
R1292 B.n570 B.n542 71.676
R1293 B.n566 B.n543 71.676
R1294 B.n562 B.n544 71.676
R1295 B.n558 B.n545 71.676
R1296 B.n554 B.n546 71.676
R1297 B.n817 B.n548 71.676
R1298 B.n809 B.n482 71.676
R1299 B.n805 B.n483 71.676
R1300 B.n801 B.n484 71.676
R1301 B.n797 B.n485 71.676
R1302 B.n793 B.n486 71.676
R1303 B.n789 B.n487 71.676
R1304 B.n785 B.n488 71.676
R1305 B.n781 B.n489 71.676
R1306 B.n777 B.n490 71.676
R1307 B.n773 B.n491 71.676
R1308 B.n769 B.n492 71.676
R1309 B.n765 B.n493 71.676
R1310 B.n761 B.n494 71.676
R1311 B.n757 B.n495 71.676
R1312 B.n753 B.n496 71.676
R1313 B.n749 B.n497 71.676
R1314 B.n745 B.n498 71.676
R1315 B.n741 B.n499 71.676
R1316 B.n737 B.n500 71.676
R1317 B.n733 B.n501 71.676
R1318 B.n729 B.n502 71.676
R1319 B.n725 B.n503 71.676
R1320 B.n721 B.n504 71.676
R1321 B.n717 B.n505 71.676
R1322 B.n713 B.n506 71.676
R1323 B.n709 B.n507 71.676
R1324 B.n705 B.n508 71.676
R1325 B.n701 B.n509 71.676
R1326 B.n697 B.n510 71.676
R1327 B.n692 B.n511 71.676
R1328 B.n688 B.n512 71.676
R1329 B.n684 B.n513 71.676
R1330 B.n680 B.n514 71.676
R1331 B.n676 B.n515 71.676
R1332 B.n671 B.n516 71.676
R1333 B.n667 B.n517 71.676
R1334 B.n663 B.n518 71.676
R1335 B.n659 B.n519 71.676
R1336 B.n655 B.n520 71.676
R1337 B.n651 B.n521 71.676
R1338 B.n647 B.n522 71.676
R1339 B.n643 B.n523 71.676
R1340 B.n639 B.n524 71.676
R1341 B.n635 B.n525 71.676
R1342 B.n631 B.n526 71.676
R1343 B.n627 B.n527 71.676
R1344 B.n623 B.n528 71.676
R1345 B.n619 B.n529 71.676
R1346 B.n615 B.n530 71.676
R1347 B.n611 B.n531 71.676
R1348 B.n607 B.n532 71.676
R1349 B.n603 B.n533 71.676
R1350 B.n599 B.n534 71.676
R1351 B.n595 B.n535 71.676
R1352 B.n591 B.n536 71.676
R1353 B.n587 B.n537 71.676
R1354 B.n583 B.n538 71.676
R1355 B.n579 B.n539 71.676
R1356 B.n575 B.n540 71.676
R1357 B.n571 B.n541 71.676
R1358 B.n567 B.n542 71.676
R1359 B.n563 B.n543 71.676
R1360 B.n559 B.n544 71.676
R1361 B.n555 B.n545 71.676
R1362 B.n546 B.n481 71.676
R1363 B.n1061 B.n1060 71.676
R1364 B.n1061 B.n2 71.676
R1365 B.n139 B.t19 67.3837
R1366 B.n552 B.t11 67.3837
R1367 B.n142 B.t16 67.358
R1368 B.n550 B.t8 67.358
R1369 B.n818 B.n478 60.1444
R1370 B.n985 B.n984 60.1444
R1371 B.n143 B.n142 59.5399
R1372 B.n140 B.n139 59.5399
R1373 B.n673 B.n552 59.5399
R1374 B.n694 B.n550 59.5399
R1375 B.n142 B.n141 48.6793
R1376 B.n139 B.n138 48.6793
R1377 B.n552 B.n551 48.6793
R1378 B.n550 B.n549 48.6793
R1379 B.n815 B.n476 35.4346
R1380 B.n821 B.n820 35.4346
R1381 B.n145 B.n67 35.4346
R1382 B.n981 B.n980 35.4346
R1383 B.n824 B.n478 30.7508
R1384 B.n824 B.n474 30.7508
R1385 B.n830 B.n474 30.7508
R1386 B.n830 B.n470 30.7508
R1387 B.n837 B.n470 30.7508
R1388 B.n837 B.n836 30.7508
R1389 B.n843 B.n463 30.7508
R1390 B.n849 B.n463 30.7508
R1391 B.n849 B.n459 30.7508
R1392 B.n855 B.n459 30.7508
R1393 B.n855 B.n455 30.7508
R1394 B.n861 B.n455 30.7508
R1395 B.n861 B.n451 30.7508
R1396 B.n867 B.n451 30.7508
R1397 B.n867 B.n447 30.7508
R1398 B.n873 B.n447 30.7508
R1399 B.n879 B.n443 30.7508
R1400 B.n879 B.n439 30.7508
R1401 B.n885 B.n439 30.7508
R1402 B.n885 B.n434 30.7508
R1403 B.n891 B.n434 30.7508
R1404 B.n891 B.n435 30.7508
R1405 B.n897 B.n427 30.7508
R1406 B.n903 B.n427 30.7508
R1407 B.n903 B.n423 30.7508
R1408 B.n909 B.n423 30.7508
R1409 B.n909 B.n418 30.7508
R1410 B.n915 B.n418 30.7508
R1411 B.n915 B.n419 30.7508
R1412 B.n922 B.n411 30.7508
R1413 B.n928 B.n411 30.7508
R1414 B.n928 B.n4 30.7508
R1415 B.n1059 B.n4 30.7508
R1416 B.n1059 B.n1058 30.7508
R1417 B.n1058 B.n1057 30.7508
R1418 B.n1057 B.n8 30.7508
R1419 B.n12 B.n8 30.7508
R1420 B.n1050 B.n12 30.7508
R1421 B.n1049 B.n1048 30.7508
R1422 B.n1048 B.n16 30.7508
R1423 B.n1042 B.n16 30.7508
R1424 B.n1042 B.n1041 30.7508
R1425 B.n1041 B.n1040 30.7508
R1426 B.n1040 B.n23 30.7508
R1427 B.n1034 B.n23 30.7508
R1428 B.n1033 B.n1032 30.7508
R1429 B.n1032 B.n30 30.7508
R1430 B.n1026 B.n30 30.7508
R1431 B.n1026 B.n1025 30.7508
R1432 B.n1025 B.n1024 30.7508
R1433 B.n1024 B.n37 30.7508
R1434 B.n1018 B.n1017 30.7508
R1435 B.n1017 B.n1016 30.7508
R1436 B.n1016 B.n44 30.7508
R1437 B.n1010 B.n44 30.7508
R1438 B.n1010 B.n1009 30.7508
R1439 B.n1009 B.n1008 30.7508
R1440 B.n1008 B.n51 30.7508
R1441 B.n1002 B.n51 30.7508
R1442 B.n1002 B.n1001 30.7508
R1443 B.n1001 B.n1000 30.7508
R1444 B.n994 B.n61 30.7508
R1445 B.n994 B.n993 30.7508
R1446 B.n993 B.n992 30.7508
R1447 B.n992 B.n65 30.7508
R1448 B.n986 B.n65 30.7508
R1449 B.n986 B.n985 30.7508
R1450 B.n836 B.t7 26.2287
R1451 B.n61 B.t14 26.2287
R1452 B.n435 B.t0 25.3242
R1453 B.t4 B.n1033 25.3242
R1454 B.n922 B.t3 24.4198
R1455 B.n1050 B.t5 24.4198
R1456 B B.n1062 18.0485
R1457 B.t1 B.n443 17.1845
R1458 B.t2 B.n37 17.1845
R1459 B.n873 B.t1 13.5668
R1460 B.n1018 B.t2 13.5668
R1461 B.n826 B.n476 10.6151
R1462 B.n827 B.n826 10.6151
R1463 B.n828 B.n827 10.6151
R1464 B.n828 B.n468 10.6151
R1465 B.n839 B.n468 10.6151
R1466 B.n840 B.n839 10.6151
R1467 B.n841 B.n840 10.6151
R1468 B.n841 B.n461 10.6151
R1469 B.n851 B.n461 10.6151
R1470 B.n852 B.n851 10.6151
R1471 B.n853 B.n852 10.6151
R1472 B.n853 B.n453 10.6151
R1473 B.n863 B.n453 10.6151
R1474 B.n864 B.n863 10.6151
R1475 B.n865 B.n864 10.6151
R1476 B.n865 B.n445 10.6151
R1477 B.n875 B.n445 10.6151
R1478 B.n876 B.n875 10.6151
R1479 B.n877 B.n876 10.6151
R1480 B.n877 B.n437 10.6151
R1481 B.n887 B.n437 10.6151
R1482 B.n888 B.n887 10.6151
R1483 B.n889 B.n888 10.6151
R1484 B.n889 B.n429 10.6151
R1485 B.n899 B.n429 10.6151
R1486 B.n900 B.n899 10.6151
R1487 B.n901 B.n900 10.6151
R1488 B.n901 B.n421 10.6151
R1489 B.n911 B.n421 10.6151
R1490 B.n912 B.n911 10.6151
R1491 B.n913 B.n912 10.6151
R1492 B.n913 B.n413 10.6151
R1493 B.n924 B.n413 10.6151
R1494 B.n925 B.n924 10.6151
R1495 B.n926 B.n925 10.6151
R1496 B.n926 B.n0 10.6151
R1497 B.n815 B.n814 10.6151
R1498 B.n814 B.n813 10.6151
R1499 B.n813 B.n812 10.6151
R1500 B.n812 B.n810 10.6151
R1501 B.n810 B.n807 10.6151
R1502 B.n807 B.n806 10.6151
R1503 B.n806 B.n803 10.6151
R1504 B.n803 B.n802 10.6151
R1505 B.n802 B.n799 10.6151
R1506 B.n799 B.n798 10.6151
R1507 B.n798 B.n795 10.6151
R1508 B.n795 B.n794 10.6151
R1509 B.n794 B.n791 10.6151
R1510 B.n791 B.n790 10.6151
R1511 B.n790 B.n787 10.6151
R1512 B.n787 B.n786 10.6151
R1513 B.n786 B.n783 10.6151
R1514 B.n783 B.n782 10.6151
R1515 B.n782 B.n779 10.6151
R1516 B.n779 B.n778 10.6151
R1517 B.n778 B.n775 10.6151
R1518 B.n775 B.n774 10.6151
R1519 B.n774 B.n771 10.6151
R1520 B.n771 B.n770 10.6151
R1521 B.n770 B.n767 10.6151
R1522 B.n767 B.n766 10.6151
R1523 B.n766 B.n763 10.6151
R1524 B.n763 B.n762 10.6151
R1525 B.n762 B.n759 10.6151
R1526 B.n759 B.n758 10.6151
R1527 B.n758 B.n755 10.6151
R1528 B.n755 B.n754 10.6151
R1529 B.n754 B.n751 10.6151
R1530 B.n751 B.n750 10.6151
R1531 B.n750 B.n747 10.6151
R1532 B.n747 B.n746 10.6151
R1533 B.n746 B.n743 10.6151
R1534 B.n743 B.n742 10.6151
R1535 B.n742 B.n739 10.6151
R1536 B.n739 B.n738 10.6151
R1537 B.n738 B.n735 10.6151
R1538 B.n735 B.n734 10.6151
R1539 B.n734 B.n731 10.6151
R1540 B.n731 B.n730 10.6151
R1541 B.n730 B.n727 10.6151
R1542 B.n727 B.n726 10.6151
R1543 B.n726 B.n723 10.6151
R1544 B.n723 B.n722 10.6151
R1545 B.n722 B.n719 10.6151
R1546 B.n719 B.n718 10.6151
R1547 B.n718 B.n715 10.6151
R1548 B.n715 B.n714 10.6151
R1549 B.n714 B.n711 10.6151
R1550 B.n711 B.n710 10.6151
R1551 B.n710 B.n707 10.6151
R1552 B.n707 B.n706 10.6151
R1553 B.n706 B.n703 10.6151
R1554 B.n703 B.n702 10.6151
R1555 B.n702 B.n699 10.6151
R1556 B.n699 B.n698 10.6151
R1557 B.n698 B.n695 10.6151
R1558 B.n693 B.n690 10.6151
R1559 B.n690 B.n689 10.6151
R1560 B.n689 B.n686 10.6151
R1561 B.n686 B.n685 10.6151
R1562 B.n685 B.n682 10.6151
R1563 B.n682 B.n681 10.6151
R1564 B.n681 B.n678 10.6151
R1565 B.n678 B.n677 10.6151
R1566 B.n677 B.n674 10.6151
R1567 B.n672 B.n669 10.6151
R1568 B.n669 B.n668 10.6151
R1569 B.n668 B.n665 10.6151
R1570 B.n665 B.n664 10.6151
R1571 B.n664 B.n661 10.6151
R1572 B.n661 B.n660 10.6151
R1573 B.n660 B.n657 10.6151
R1574 B.n657 B.n656 10.6151
R1575 B.n656 B.n653 10.6151
R1576 B.n653 B.n652 10.6151
R1577 B.n652 B.n649 10.6151
R1578 B.n649 B.n648 10.6151
R1579 B.n648 B.n645 10.6151
R1580 B.n645 B.n644 10.6151
R1581 B.n644 B.n641 10.6151
R1582 B.n641 B.n640 10.6151
R1583 B.n640 B.n637 10.6151
R1584 B.n637 B.n636 10.6151
R1585 B.n636 B.n633 10.6151
R1586 B.n633 B.n632 10.6151
R1587 B.n632 B.n629 10.6151
R1588 B.n629 B.n628 10.6151
R1589 B.n628 B.n625 10.6151
R1590 B.n625 B.n624 10.6151
R1591 B.n624 B.n621 10.6151
R1592 B.n621 B.n620 10.6151
R1593 B.n620 B.n617 10.6151
R1594 B.n617 B.n616 10.6151
R1595 B.n616 B.n613 10.6151
R1596 B.n613 B.n612 10.6151
R1597 B.n612 B.n609 10.6151
R1598 B.n609 B.n608 10.6151
R1599 B.n608 B.n605 10.6151
R1600 B.n605 B.n604 10.6151
R1601 B.n604 B.n601 10.6151
R1602 B.n601 B.n600 10.6151
R1603 B.n600 B.n597 10.6151
R1604 B.n597 B.n596 10.6151
R1605 B.n596 B.n593 10.6151
R1606 B.n593 B.n592 10.6151
R1607 B.n592 B.n589 10.6151
R1608 B.n589 B.n588 10.6151
R1609 B.n588 B.n585 10.6151
R1610 B.n585 B.n584 10.6151
R1611 B.n584 B.n581 10.6151
R1612 B.n581 B.n580 10.6151
R1613 B.n580 B.n577 10.6151
R1614 B.n577 B.n576 10.6151
R1615 B.n576 B.n573 10.6151
R1616 B.n573 B.n572 10.6151
R1617 B.n572 B.n569 10.6151
R1618 B.n569 B.n568 10.6151
R1619 B.n568 B.n565 10.6151
R1620 B.n565 B.n564 10.6151
R1621 B.n564 B.n561 10.6151
R1622 B.n561 B.n560 10.6151
R1623 B.n560 B.n557 10.6151
R1624 B.n557 B.n556 10.6151
R1625 B.n556 B.n553 10.6151
R1626 B.n553 B.n480 10.6151
R1627 B.n820 B.n480 10.6151
R1628 B.n822 B.n821 10.6151
R1629 B.n822 B.n472 10.6151
R1630 B.n832 B.n472 10.6151
R1631 B.n833 B.n832 10.6151
R1632 B.n834 B.n833 10.6151
R1633 B.n834 B.n465 10.6151
R1634 B.n845 B.n465 10.6151
R1635 B.n846 B.n845 10.6151
R1636 B.n847 B.n846 10.6151
R1637 B.n847 B.n457 10.6151
R1638 B.n857 B.n457 10.6151
R1639 B.n858 B.n857 10.6151
R1640 B.n859 B.n858 10.6151
R1641 B.n859 B.n449 10.6151
R1642 B.n869 B.n449 10.6151
R1643 B.n870 B.n869 10.6151
R1644 B.n871 B.n870 10.6151
R1645 B.n871 B.n441 10.6151
R1646 B.n881 B.n441 10.6151
R1647 B.n882 B.n881 10.6151
R1648 B.n883 B.n882 10.6151
R1649 B.n883 B.n432 10.6151
R1650 B.n893 B.n432 10.6151
R1651 B.n894 B.n893 10.6151
R1652 B.n895 B.n894 10.6151
R1653 B.n895 B.n425 10.6151
R1654 B.n905 B.n425 10.6151
R1655 B.n906 B.n905 10.6151
R1656 B.n907 B.n906 10.6151
R1657 B.n907 B.n416 10.6151
R1658 B.n917 B.n416 10.6151
R1659 B.n918 B.n917 10.6151
R1660 B.n920 B.n918 10.6151
R1661 B.n920 B.n919 10.6151
R1662 B.n919 B.n409 10.6151
R1663 B.n931 B.n409 10.6151
R1664 B.n932 B.n931 10.6151
R1665 B.n933 B.n932 10.6151
R1666 B.n934 B.n933 10.6151
R1667 B.n935 B.n934 10.6151
R1668 B.n938 B.n935 10.6151
R1669 B.n939 B.n938 10.6151
R1670 B.n940 B.n939 10.6151
R1671 B.n941 B.n940 10.6151
R1672 B.n943 B.n941 10.6151
R1673 B.n944 B.n943 10.6151
R1674 B.n945 B.n944 10.6151
R1675 B.n946 B.n945 10.6151
R1676 B.n948 B.n946 10.6151
R1677 B.n949 B.n948 10.6151
R1678 B.n950 B.n949 10.6151
R1679 B.n951 B.n950 10.6151
R1680 B.n953 B.n951 10.6151
R1681 B.n954 B.n953 10.6151
R1682 B.n955 B.n954 10.6151
R1683 B.n956 B.n955 10.6151
R1684 B.n958 B.n956 10.6151
R1685 B.n959 B.n958 10.6151
R1686 B.n960 B.n959 10.6151
R1687 B.n961 B.n960 10.6151
R1688 B.n963 B.n961 10.6151
R1689 B.n964 B.n963 10.6151
R1690 B.n965 B.n964 10.6151
R1691 B.n966 B.n965 10.6151
R1692 B.n968 B.n966 10.6151
R1693 B.n969 B.n968 10.6151
R1694 B.n970 B.n969 10.6151
R1695 B.n971 B.n970 10.6151
R1696 B.n973 B.n971 10.6151
R1697 B.n974 B.n973 10.6151
R1698 B.n975 B.n974 10.6151
R1699 B.n976 B.n975 10.6151
R1700 B.n978 B.n976 10.6151
R1701 B.n979 B.n978 10.6151
R1702 B.n980 B.n979 10.6151
R1703 B.n1054 B.n1 10.6151
R1704 B.n1054 B.n1053 10.6151
R1705 B.n1053 B.n1052 10.6151
R1706 B.n1052 B.n10 10.6151
R1707 B.n1046 B.n10 10.6151
R1708 B.n1046 B.n1045 10.6151
R1709 B.n1045 B.n1044 10.6151
R1710 B.n1044 B.n18 10.6151
R1711 B.n1038 B.n18 10.6151
R1712 B.n1038 B.n1037 10.6151
R1713 B.n1037 B.n1036 10.6151
R1714 B.n1036 B.n25 10.6151
R1715 B.n1030 B.n25 10.6151
R1716 B.n1030 B.n1029 10.6151
R1717 B.n1029 B.n1028 10.6151
R1718 B.n1028 B.n32 10.6151
R1719 B.n1022 B.n32 10.6151
R1720 B.n1022 B.n1021 10.6151
R1721 B.n1021 B.n1020 10.6151
R1722 B.n1020 B.n39 10.6151
R1723 B.n1014 B.n39 10.6151
R1724 B.n1014 B.n1013 10.6151
R1725 B.n1013 B.n1012 10.6151
R1726 B.n1012 B.n46 10.6151
R1727 B.n1006 B.n46 10.6151
R1728 B.n1006 B.n1005 10.6151
R1729 B.n1005 B.n1004 10.6151
R1730 B.n1004 B.n53 10.6151
R1731 B.n998 B.n53 10.6151
R1732 B.n998 B.n997 10.6151
R1733 B.n997 B.n996 10.6151
R1734 B.n996 B.n59 10.6151
R1735 B.n990 B.n59 10.6151
R1736 B.n990 B.n989 10.6151
R1737 B.n989 B.n988 10.6151
R1738 B.n988 B.n67 10.6151
R1739 B.n146 B.n145 10.6151
R1740 B.n149 B.n146 10.6151
R1741 B.n150 B.n149 10.6151
R1742 B.n153 B.n150 10.6151
R1743 B.n154 B.n153 10.6151
R1744 B.n157 B.n154 10.6151
R1745 B.n158 B.n157 10.6151
R1746 B.n161 B.n158 10.6151
R1747 B.n162 B.n161 10.6151
R1748 B.n165 B.n162 10.6151
R1749 B.n166 B.n165 10.6151
R1750 B.n169 B.n166 10.6151
R1751 B.n170 B.n169 10.6151
R1752 B.n173 B.n170 10.6151
R1753 B.n174 B.n173 10.6151
R1754 B.n177 B.n174 10.6151
R1755 B.n178 B.n177 10.6151
R1756 B.n181 B.n178 10.6151
R1757 B.n182 B.n181 10.6151
R1758 B.n185 B.n182 10.6151
R1759 B.n186 B.n185 10.6151
R1760 B.n189 B.n186 10.6151
R1761 B.n190 B.n189 10.6151
R1762 B.n193 B.n190 10.6151
R1763 B.n194 B.n193 10.6151
R1764 B.n197 B.n194 10.6151
R1765 B.n198 B.n197 10.6151
R1766 B.n201 B.n198 10.6151
R1767 B.n202 B.n201 10.6151
R1768 B.n205 B.n202 10.6151
R1769 B.n206 B.n205 10.6151
R1770 B.n209 B.n206 10.6151
R1771 B.n210 B.n209 10.6151
R1772 B.n213 B.n210 10.6151
R1773 B.n214 B.n213 10.6151
R1774 B.n217 B.n214 10.6151
R1775 B.n218 B.n217 10.6151
R1776 B.n221 B.n218 10.6151
R1777 B.n222 B.n221 10.6151
R1778 B.n225 B.n222 10.6151
R1779 B.n226 B.n225 10.6151
R1780 B.n229 B.n226 10.6151
R1781 B.n230 B.n229 10.6151
R1782 B.n233 B.n230 10.6151
R1783 B.n234 B.n233 10.6151
R1784 B.n237 B.n234 10.6151
R1785 B.n238 B.n237 10.6151
R1786 B.n241 B.n238 10.6151
R1787 B.n242 B.n241 10.6151
R1788 B.n245 B.n242 10.6151
R1789 B.n246 B.n245 10.6151
R1790 B.n249 B.n246 10.6151
R1791 B.n250 B.n249 10.6151
R1792 B.n253 B.n250 10.6151
R1793 B.n254 B.n253 10.6151
R1794 B.n257 B.n254 10.6151
R1795 B.n258 B.n257 10.6151
R1796 B.n261 B.n258 10.6151
R1797 B.n262 B.n261 10.6151
R1798 B.n265 B.n262 10.6151
R1799 B.n266 B.n265 10.6151
R1800 B.n270 B.n269 10.6151
R1801 B.n273 B.n270 10.6151
R1802 B.n274 B.n273 10.6151
R1803 B.n277 B.n274 10.6151
R1804 B.n278 B.n277 10.6151
R1805 B.n281 B.n278 10.6151
R1806 B.n282 B.n281 10.6151
R1807 B.n285 B.n282 10.6151
R1808 B.n286 B.n285 10.6151
R1809 B.n290 B.n289 10.6151
R1810 B.n293 B.n290 10.6151
R1811 B.n294 B.n293 10.6151
R1812 B.n297 B.n294 10.6151
R1813 B.n298 B.n297 10.6151
R1814 B.n301 B.n298 10.6151
R1815 B.n302 B.n301 10.6151
R1816 B.n305 B.n302 10.6151
R1817 B.n306 B.n305 10.6151
R1818 B.n309 B.n306 10.6151
R1819 B.n310 B.n309 10.6151
R1820 B.n313 B.n310 10.6151
R1821 B.n314 B.n313 10.6151
R1822 B.n317 B.n314 10.6151
R1823 B.n318 B.n317 10.6151
R1824 B.n321 B.n318 10.6151
R1825 B.n322 B.n321 10.6151
R1826 B.n325 B.n322 10.6151
R1827 B.n326 B.n325 10.6151
R1828 B.n329 B.n326 10.6151
R1829 B.n330 B.n329 10.6151
R1830 B.n333 B.n330 10.6151
R1831 B.n334 B.n333 10.6151
R1832 B.n337 B.n334 10.6151
R1833 B.n338 B.n337 10.6151
R1834 B.n341 B.n338 10.6151
R1835 B.n342 B.n341 10.6151
R1836 B.n345 B.n342 10.6151
R1837 B.n346 B.n345 10.6151
R1838 B.n349 B.n346 10.6151
R1839 B.n350 B.n349 10.6151
R1840 B.n353 B.n350 10.6151
R1841 B.n354 B.n353 10.6151
R1842 B.n357 B.n354 10.6151
R1843 B.n358 B.n357 10.6151
R1844 B.n361 B.n358 10.6151
R1845 B.n362 B.n361 10.6151
R1846 B.n365 B.n362 10.6151
R1847 B.n366 B.n365 10.6151
R1848 B.n369 B.n366 10.6151
R1849 B.n370 B.n369 10.6151
R1850 B.n373 B.n370 10.6151
R1851 B.n374 B.n373 10.6151
R1852 B.n377 B.n374 10.6151
R1853 B.n378 B.n377 10.6151
R1854 B.n381 B.n378 10.6151
R1855 B.n382 B.n381 10.6151
R1856 B.n385 B.n382 10.6151
R1857 B.n386 B.n385 10.6151
R1858 B.n389 B.n386 10.6151
R1859 B.n390 B.n389 10.6151
R1860 B.n393 B.n390 10.6151
R1861 B.n394 B.n393 10.6151
R1862 B.n397 B.n394 10.6151
R1863 B.n398 B.n397 10.6151
R1864 B.n401 B.n398 10.6151
R1865 B.n402 B.n401 10.6151
R1866 B.n405 B.n402 10.6151
R1867 B.n407 B.n405 10.6151
R1868 B.n408 B.n407 10.6151
R1869 B.n981 B.n408 10.6151
R1870 B.n695 B.n694 9.36635
R1871 B.n673 B.n672 9.36635
R1872 B.n266 B.n143 9.36635
R1873 B.n289 B.n140 9.36635
R1874 B.n1062 B.n0 8.11757
R1875 B.n1062 B.n1 8.11757
R1876 B.n419 B.t3 6.33144
R1877 B.t5 B.n1049 6.33144
R1878 B.n897 B.t0 5.42702
R1879 B.n1034 B.t4 5.42702
R1880 B.n843 B.t7 4.5226
R1881 B.n1000 B.t14 4.5226
R1882 B.n694 B.n693 1.24928
R1883 B.n674 B.n673 1.24928
R1884 B.n269 B.n143 1.24928
R1885 B.n286 B.n140 1.24928
R1886 VN.n3 VN.t4 242.743
R1887 VN.n17 VN.t5 242.743
R1888 VN.n4 VN.t2 210.6
R1889 VN.n12 VN.t0 210.6
R1890 VN.n18 VN.t3 210.6
R1891 VN.n26 VN.t1 210.6
R1892 VN.n25 VN.n14 161.3
R1893 VN.n24 VN.n23 161.3
R1894 VN.n22 VN.n15 161.3
R1895 VN.n21 VN.n20 161.3
R1896 VN.n19 VN.n16 161.3
R1897 VN.n11 VN.n0 161.3
R1898 VN.n10 VN.n9 161.3
R1899 VN.n8 VN.n1 161.3
R1900 VN.n7 VN.n6 161.3
R1901 VN.n5 VN.n2 161.3
R1902 VN.n13 VN.n12 98.0336
R1903 VN.n27 VN.n26 98.0336
R1904 VN.n4 VN.n3 59.258
R1905 VN.n18 VN.n17 59.258
R1906 VN VN.n27 52.608
R1907 VN.n10 VN.n1 40.979
R1908 VN.n24 VN.n15 40.979
R1909 VN.n6 VN.n1 40.0078
R1910 VN.n20 VN.n15 40.0078
R1911 VN.n6 VN.n5 24.4675
R1912 VN.n11 VN.n10 24.4675
R1913 VN.n20 VN.n19 24.4675
R1914 VN.n25 VN.n24 24.4675
R1915 VN.n12 VN.n11 12.7233
R1916 VN.n26 VN.n25 12.7233
R1917 VN.n5 VN.n4 12.234
R1918 VN.n19 VN.n18 12.234
R1919 VN.n17 VN.n16 9.6787
R1920 VN.n3 VN.n2 9.6787
R1921 VN.n27 VN.n14 0.278367
R1922 VN.n13 VN.n0 0.278367
R1923 VN.n23 VN.n14 0.189894
R1924 VN.n23 VN.n22 0.189894
R1925 VN.n22 VN.n21 0.189894
R1926 VN.n21 VN.n16 0.189894
R1927 VN.n7 VN.n2 0.189894
R1928 VN.n8 VN.n7 0.189894
R1929 VN.n9 VN.n8 0.189894
R1930 VN.n9 VN.n0 0.189894
R1931 VN VN.n13 0.153454
R1932 VDD2.n1 VDD2.t1 64.5517
R1933 VDD2.n2 VDD2.t4 62.9843
R1934 VDD2.n1 VDD2.n0 62.4294
R1935 VDD2 VDD2.n3 62.4276
R1936 VDD2.n2 VDD2.n1 47.17
R1937 VDD2 VDD2.n2 1.68153
R1938 VDD2.n3 VDD2.t2 1.03987
R1939 VDD2.n3 VDD2.t0 1.03987
R1940 VDD2.n0 VDD2.t3 1.03987
R1941 VDD2.n0 VDD2.t5 1.03987
C0 VDD2 VP 0.423157f
C1 VDD1 VTAIL 10.445299f
C2 VN VTAIL 9.83629f
C3 VDD2 VTAIL 10.4908f
C4 VDD1 VN 0.149949f
C5 VTAIL VP 9.850739f
C6 VDD2 VDD1 1.2429f
C7 VDD2 VN 10.079401f
C8 VDD1 VP 10.3479f
C9 VN VP 7.82773f
C10 VDD2 B 6.918177f
C11 VDD1 B 7.218508f
C12 VTAIL B 10.316821f
C13 VN B 12.328091f
C14 VP B 10.73079f
C15 VDD2.t1 B 3.7581f
C16 VDD2.t3 B 0.320583f
C17 VDD2.t5 B 0.320583f
C18 VDD2.n0 B 2.93577f
C19 VDD2.n1 B 2.69105f
C20 VDD2.t4 B 3.74973f
C21 VDD2.n2 B 2.73977f
C22 VDD2.t2 B 0.320583f
C23 VDD2.t0 B 0.320583f
C24 VDD2.n3 B 2.93573f
C25 VN.n0 B 0.032803f
C26 VN.t0 B 2.84507f
C27 VN.n1 B 0.020123f
C28 VN.n2 B 0.211205f
C29 VN.t2 B 2.84507f
C30 VN.t4 B 2.99335f
C31 VN.n3 B 1.04626f
C32 VN.n4 B 1.05198f
C33 VN.n5 B 0.034925f
C34 VN.n6 B 0.049573f
C35 VN.n7 B 0.024881f
C36 VN.n8 B 0.024881f
C37 VN.n9 B 0.024881f
C38 VN.n10 B 0.049324f
C39 VN.n11 B 0.035383f
C40 VN.n12 B 1.06092f
C41 VN.n13 B 0.035756f
C42 VN.n14 B 0.032803f
C43 VN.t1 B 2.84507f
C44 VN.n15 B 0.020123f
C45 VN.n16 B 0.211205f
C46 VN.t3 B 2.84507f
C47 VN.t5 B 2.99335f
C48 VN.n17 B 1.04626f
C49 VN.n18 B 1.05198f
C50 VN.n19 B 0.034925f
C51 VN.n20 B 0.049573f
C52 VN.n21 B 0.024881f
C53 VN.n22 B 0.024881f
C54 VN.n23 B 0.024881f
C55 VN.n24 B 0.049324f
C56 VN.n25 B 0.035383f
C57 VN.n26 B 1.06092f
C58 VN.n27 B 1.48663f
C59 VTAIL.t5 B 0.335141f
C60 VTAIL.t4 B 0.335141f
C61 VTAIL.n0 B 3.00158f
C62 VTAIL.n1 B 0.368027f
C63 VTAIL.t10 B 3.83522f
C64 VTAIL.n2 B 0.560651f
C65 VTAIL.t6 B 0.335141f
C66 VTAIL.t11 B 0.335141f
C67 VTAIL.n3 B 3.00158f
C68 VTAIL.n4 B 2.15988f
C69 VTAIL.t1 B 0.335141f
C70 VTAIL.t0 B 0.335141f
C71 VTAIL.n5 B 3.00159f
C72 VTAIL.n6 B 2.15988f
C73 VTAIL.t3 B 3.83524f
C74 VTAIL.n7 B 0.560623f
C75 VTAIL.t7 B 0.335141f
C76 VTAIL.t8 B 0.335141f
C77 VTAIL.n8 B 3.00159f
C78 VTAIL.n9 B 0.48026f
C79 VTAIL.t9 B 3.83522f
C80 VTAIL.n10 B 2.08505f
C81 VTAIL.t2 B 3.83522f
C82 VTAIL.n11 B 2.04207f
C83 VDD1.t3 B 3.76279f
C84 VDD1.t2 B 3.76198f
C85 VDD1.t1 B 0.320914f
C86 VDD1.t0 B 0.320914f
C87 VDD1.n0 B 2.9388f
C88 VDD1.n1 B 2.7939f
C89 VDD1.t4 B 0.320914f
C90 VDD1.t5 B 0.320914f
C91 VDD1.n2 B 2.93596f
C92 VDD1.n3 B 2.73002f
C93 VP.n0 B 0.0332f
C94 VP.t1 B 2.87952f
C95 VP.n1 B 0.020367f
C96 VP.n2 B 0.025182f
C97 VP.t0 B 2.87952f
C98 VP.n3 B 0.050173f
C99 VP.n4 B 0.025182f
C100 VP.t5 B 2.87952f
C101 VP.n5 B 1.07376f
C102 VP.n6 B 0.0332f
C103 VP.t2 B 2.87952f
C104 VP.n7 B 0.020367f
C105 VP.n8 B 0.213762f
C106 VP.t3 B 2.87952f
C107 VP.t4 B 3.02959f
C108 VP.n9 B 1.05893f
C109 VP.n10 B 1.06472f
C110 VP.n11 B 0.035348f
C111 VP.n12 B 0.050173f
C112 VP.n13 B 0.025182f
C113 VP.n14 B 0.025182f
C114 VP.n15 B 0.025182f
C115 VP.n16 B 0.049921f
C116 VP.n17 B 0.035811f
C117 VP.n18 B 1.07376f
C118 VP.n19 B 1.49119f
C119 VP.n20 B 1.50849f
C120 VP.n21 B 0.0332f
C121 VP.n22 B 0.035811f
C122 VP.n23 B 0.049921f
C123 VP.n24 B 0.020367f
C124 VP.n25 B 0.025182f
C125 VP.n26 B 0.025182f
C126 VP.n27 B 0.025182f
C127 VP.n28 B 0.035348f
C128 VP.n29 B 1.0001f
C129 VP.n30 B 0.035348f
C130 VP.n31 B 0.050173f
C131 VP.n32 B 0.025182f
C132 VP.n33 B 0.025182f
C133 VP.n34 B 0.025182f
C134 VP.n35 B 0.049921f
C135 VP.n36 B 0.035811f
C136 VP.n37 B 1.07376f
C137 VP.n38 B 0.036188f
.ends

