* NGSPICE file created from opamp_sample_0002.ext - technology: sky130A

.subckt opamp_sample_0002 GND VOUT VDD VN VP CS_BIAS DIFFPAIR_BIAS
X0 VDD.t194 a_n7677_8299.t20 VOUT.t54 VDD.t127 sky130_fd_pr__pfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X1 a_n2686_8422.t19 a_n2686_12778.t32 a_n7677_8299.t1 VDD.t4 sky130_fd_pr__pfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X2 VOUT.t53 a_n7677_8299.t21 VDD.t193 VDD.t137 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X3 GND.t158 GND.t156 GND.t157 GND.t79 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X4 CS_BIAS.t31 CS_BIAS.t30 GND.t41 GND.t40 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X5 GND.t165 CS_BIAS.t32 VOUT.t24 GND.t0 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=2
X6 a_n2686_8422.t7 a_n2686_12778.t33 VDD.t29 VDD.t28 sky130_fd_pr__pfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=1
X7 GND.t155 GND.t153 GND.t154 GND.t103 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X8 VOUT.t10 CS_BIAS.t33 GND.t50 GND.t42 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X9 VDD.t192 a_n7677_8299.t22 VOUT.t52 VDD.t154 sky130_fd_pr__pfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X10 GND.t163 CS_BIAS.t34 VOUT.t22 GND.t48 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X11 GND.t152 GND.t150 GND.t151 GND.t79 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X12 VDD.t114 VDD.t112 VDD.t113 VDD.t71 sky130_fd_pr__pfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X13 GND.t149 GND.t147 VN.t4 GND.t148 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X14 GND.t146 GND.t144 GND.t145 GND.t75 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X15 a_n2511_10556.t11 a_n2686_12778.t19 a_n2686_12778.t20 VDD.t8 sky130_fd_pr__pfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X16 a_n7677_8299.t19 a_n2686_12778.t34 a_n2686_8422.t18 VDD.t36 sky130_fd_pr__pfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X17 VDD.t111 VDD.t109 VDD.t110 VDD.t87 sky130_fd_pr__pfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=1
X18 GND.t64 CS_BIAS.t28 CS_BIAS.t29 GND.t9 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X19 VDD.t191 a_n7677_8299.t23 VOUT.t61 VDD.t119 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X20 VDD.t190 a_n7677_8299.t24 VOUT.t60 VDD.t143 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X21 VOUT.t19 CS_BIAS.t35 GND.t66 GND.t28 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X22 VOUT.t59 a_n7677_8299.t25 VDD.t189 VDD.t156 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X23 VDD.t188 a_n7677_8299.t26 VOUT.t58 VDD.t160 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X24 a_n7677_8299.t0 VN.t5 a_n1455_n3928.t15 GND.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X25 GND.t143 GND.t141 VP.t4 GND.t142 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X26 GND.t170 CS_BIAS.t26 CS_BIAS.t27 GND.t2 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X27 VDD.t187 a_n7677_8299.t27 VOUT.t76 VDD.t158 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X28 GND.t59 CS_BIAS.t36 VOUT.t16 GND.t32 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X29 GND.t10 CS_BIAS.t37 VOUT.t2 GND.t9 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X30 VOUT.t75 a_n7677_8299.t28 VDD.t186 VDD.t156 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X31 VOUT.t92 a_n2686_8422.t20 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X32 VDD.t108 VDD.t106 VDD.t107 VDD.t63 sky130_fd_pr__pfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X33 a_n7677_8299.t5 a_n2686_12778.t35 a_n2686_8422.t17 VDD.t7 sky130_fd_pr__pfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=1
X34 VDD.t105 VDD.t102 VDD.t104 VDD.t103 sky130_fd_pr__pfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=1
X35 GND.t58 CS_BIAS.t38 VOUT.t15 GND.t57 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=2
X36 VDD.t196 a_n2686_12778.t36 a_n2511_10556.t19 VDD.t195 sky130_fd_pr__pfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=1
X37 VDD.t185 a_n7677_8299.t29 VOUT.t74 VDD.t135 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X38 GND.t140 GND.t138 GND.t139 GND.t83 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X39 VOUT.t73 a_n7677_8299.t30 VDD.t184 VDD.t145 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X40 a_n2686_8422.t16 a_n2686_12778.t37 a_n7677_8299.t10 VDD.t33 sky130_fd_pr__pfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=1
X41 a_n1455_n3928.t6 DIFFPAIR_BIAS.t8 GND.t35 GND.t34 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=2
X42 CS_BIAS.t25 CS_BIAS.t24 GND.t47 GND.t46 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X43 a_n2511_10556.t10 a_n2686_12778.t25 a_n2686_12778.t26 VDD.t36 sky130_fd_pr__pfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X44 GND.t137 GND.t135 GND.t136 GND.t75 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X45 VDD.t183 a_n7677_8299.t31 VOUT.t49 VDD.t149 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X46 DIFFPAIR_BIAS.t7 DIFFPAIR_BIAS.t6 GND.t174 GND.t173 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=2
X47 GND.t134 GND.t131 GND.t133 GND.t132 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=2
X48 VDD.t10 a_n2686_12778.t38 a_n2511_10556.t18 VDD.t9 sky130_fd_pr__pfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X49 VDD.t17 a_n2686_12778.t39 a_n2686_8422.t6 VDD.t16 sky130_fd_pr__pfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=1
X50 a_n7677_8299.t6 a_n2686_12778.t40 a_n2686_8422.t15 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=1
X51 GND.t130 GND.t128 GND.t129 GND.t90 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X52 GND.t127 GND.t124 GND.t126 GND.t125 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=2
X53 GND.t53 CS_BIAS.t39 VOUT.t12 GND.t0 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=2
X54 a_n1455_n3928.t0 VP.t5 a_n2686_12778.t0 GND.t13 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X55 GND.t123 GND.t121 GND.t122 GND.t103 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X56 VN.t3 GND.t118 GND.t120 GND.t119 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X57 DIFFPAIR_BIAS.t5 DIFFPAIR_BIAS.t4 GND.t12 GND.t11 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=2
X58 VOUT.t48 a_n7677_8299.t32 VDD.t182 VDD.t125 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X59 GND.t117 GND.t115 VP.t3 GND.t116 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X60 a_n2686_8422.t14 a_n2686_12778.t41 a_n7677_8299.t16 VDD.t197 sky130_fd_pr__pfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X61 VDD.t35 a_n2686_12778.t42 a_n2686_8422.t5 VDD.t34 sky130_fd_pr__pfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=1
X62 VOUT.t47 a_n7677_8299.t33 VDD.t181 VDD.t139 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X63 CS_BIAS.t23 CS_BIAS.t22 GND.t178 GND.t61 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X64 a_n1455_n3928.t2 DIFFPAIR_BIAS.t9 GND.t17 GND.t16 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=2
X65 VDD.t101 VDD.t99 VDD.t100 VDD.t44 sky130_fd_pr__pfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X66 a_n2686_8422.t13 a_n2686_12778.t43 a_n7677_8299.t11 VDD.t1 sky130_fd_pr__pfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X67 VDD.t180 a_n7677_8299.t34 VOUT.t46 VDD.t141 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X68 VDD.t179 a_n7677_8299.t35 VOUT.t80 VDD.t141 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X69 a_n1455_n3928.t14 VN.t6 a_n7677_8299.t15 GND.t21 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X70 a_n2686_12778.t5 VP.t6 a_n1455_n3928.t17 GND.t27 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X71 VDD.t199 a_n2686_12778.t44 a_n2511_10556.t17 VDD.t198 sky130_fd_pr__pfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=1
X72 a_n2511_10556.t16 a_n2686_12778.t45 VDD.t6 VDD.t5 sky130_fd_pr__pfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=1
X73 VDD.t98 VDD.t96 VDD.t97 VDD.t67 sky130_fd_pr__pfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=1
X74 GND.t114 GND.t112 VP.t2 GND.t113 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X75 VOUT.t79 a_n7677_8299.t36 VDD.t178 VDD.t137 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X76 VOUT.t78 a_n7677_8299.t37 VDD.t177 VDD.t132 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X77 VOUT.t88 CS_BIAS.t40 GND.t172 GND.t40 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X78 GND.t44 CS_BIAS.t41 VOUT.t9 GND.t9 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X79 GND.t33 CS_BIAS.t42 VOUT.t7 GND.t32 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X80 a_n7677_8299.t12 VN.t7 a_n1455_n3928.t13 GND.t63 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X81 VOUT.t90 CS_BIAS.t43 GND.t177 GND.t38 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=2
X82 a_n2686_12778.t1 VP.t7 a_n1455_n3928.t3 GND.t20 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X83 a_n1455_n3928.t12 VN.t8 a_n7677_8299.t13 GND.t60 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X84 VOUT.t77 a_n7677_8299.t38 VDD.t176 VDD.t130 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X85 a_n7677_8299.t17 a_n2686_12778.t46 a_n2686_8422.t12 VDD.t8 sky130_fd_pr__pfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X86 VN.t2 GND.t109 GND.t111 GND.t110 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X87 GND.t49 CS_BIAS.t20 CS_BIAS.t21 GND.t48 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X88 VOUT.t45 a_n7677_8299.t39 VDD.t175 VDD.t115 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X89 GND.t108 GND.t106 GND.t107 GND.t68 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X90 VDD.t174 a_n7677_8299.t40 VOUT.t44 VDD.t127 sky130_fd_pr__pfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X91 VDD.t95 VDD.t93 VDD.t94 VDD.t52 sky130_fd_pr__pfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=1
X92 a_n2511_10556.t9 a_n2686_12778.t11 a_n2686_12778.t12 VDD.t7 sky130_fd_pr__pfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=1
X93 VOUT.t11 CS_BIAS.t44 GND.t51 GND.t46 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X94 VDD.t173 a_n7677_8299.t41 VOUT.t43 VDD.t123 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X95 a_n1455_n3928.t19 VP.t8 a_n2686_12778.t31 GND.t52 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X96 VOUT.t21 CS_BIAS.t45 GND.t161 GND.t160 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X97 a_n2686_12778.t22 a_n2686_12778.t21 a_n2511_10556.t8 VDD.t33 sky130_fd_pr__pfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=1
X98 VDD.t31 a_n2686_12778.t47 a_n2686_8422.t4 VDD.t30 sky130_fd_pr__pfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X99 VOUT.t42 a_n7677_8299.t42 VDD.t172 VDD.t121 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X100 VOUT.t31 a_n7677_8299.t43 VDD.t171 VDD.t117 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X101 a_n2686_12778.t16 a_n2686_12778.t15 a_n2511_10556.t7 VDD.t25 sky130_fd_pr__pfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=1
X102 GND.t171 CS_BIAS.t18 CS_BIAS.t19 GND.t57 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=2
X103 GND.t105 GND.t102 GND.t104 GND.t103 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X104 a_n7677_8299.t18 a_n2686_12778.t48 a_n2686_8422.t11 VDD.t32 sky130_fd_pr__pfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X105 GND.t5 CS_BIAS.t46 VOUT.t1 GND.t4 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X106 VOUT.t30 a_n7677_8299.t44 VDD.t170 VDD.t115 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X107 VDD.t169 a_n7677_8299.t45 VOUT.t29 VDD.t158 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X108 a_n2686_8422.t10 a_n2686_12778.t49 a_n7677_8299.t7 VDD.t25 sky130_fd_pr__pfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=1
X109 CS_BIAS.t17 CS_BIAS.t16 GND.t168 GND.t38 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=2
X110 VDD.t92 VDD.t90 VDD.t91 VDD.t40 sky130_fd_pr__pfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X111 VOUT.t93 a_n2686_8422.t20 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X112 CS_BIAS.t15 CS_BIAS.t14 GND.t56 GND.t24 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=2
X113 VDD.t168 a_n7677_8299.t46 VOUT.t28 VDD.t149 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X114 GND.t101 GND.t99 GND.t100 GND.t83 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X115 VDD.t21 a_n2686_12778.t50 a_n2686_8422.t3 VDD.t20 sky130_fd_pr__pfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X116 GND.t1 CS_BIAS.t12 CS_BIAS.t13 GND.t0 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=2
X117 VDD.t89 VDD.t86 VDD.t88 VDD.t87 sky130_fd_pr__pfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=1
X118 a_n2511_10556.t6 a_n2686_12778.t27 a_n2686_12778.t28 VDD.t22 sky130_fd_pr__pfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X119 a_n2686_8422.t2 a_n2686_12778.t51 VDD.t3 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X120 VOUT.t26 CS_BIAS.t47 GND.t167 GND.t40 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X121 VDD.t167 a_n7677_8299.t47 VOUT.t68 VDD.t154 sky130_fd_pr__pfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X122 a_n2511_10556.t15 a_n2686_12778.t52 VDD.t12 VDD.t11 sky130_fd_pr__pfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X123 GND.t162 CS_BIAS.t10 CS_BIAS.t11 GND.t4 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X124 GND.t98 GND.t96 VN.t1 GND.t97 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X125 CS_BIAS.t9 CS_BIAS.t8 GND.t43 GND.t42 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X126 DIFFPAIR_BIAS.t3 DIFFPAIR_BIAS.t2 GND.t19 GND.t18 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=2
X127 VOUT.t8 CS_BIAS.t48 GND.t39 GND.t38 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=2
X128 a_n2511_10556.t14 a_n2686_12778.t53 VDD.t38 VDD.t37 sky130_fd_pr__pfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=1
X129 VP.t1 GND.t93 GND.t95 GND.t94 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X130 a_n7677_8299.t9 a_n2686_12778.t54 a_n2686_8422.t9 VDD.t22 sky130_fd_pr__pfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X131 VOUT.t67 a_n7677_8299.t48 VDD.t166 VDD.t139 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X132 VDD.t85 VDD.t83 VDD.t84 VDD.t71 sky130_fd_pr__pfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X133 VDD.t165 a_n7677_8299.t49 VOUT.t66 VDD.t119 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X134 GND.t45 CS_BIAS.t6 CS_BIAS.t7 GND.t32 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X135 VOUT.t65 a_n7677_8299.t50 VDD.t164 VDD.t117 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X136 VOUT.t17 CS_BIAS.t49 GND.t62 GND.t61 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X137 VDD.t163 a_n7677_8299.t51 VOUT.t87 VDD.t160 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X138 VDD.t162 a_n7677_8299.t52 VOUT.t86 VDD.t143 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X139 a_n2686_12778.t10 a_n2686_12778.t9 a_n2511_10556.t5 VDD.t13 sky130_fd_pr__pfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X140 GND.t164 CS_BIAS.t50 VOUT.t23 GND.t2 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X141 VDD.t161 a_n7677_8299.t53 VOUT.t85 VDD.t160 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X142 VOUT.t18 CS_BIAS.t51 GND.t65 GND.t46 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X143 VOUT.t27 CS_BIAS.t52 GND.t169 GND.t160 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X144 VDD.t82 VDD.t80 VDD.t81 VDD.t59 sky130_fd_pr__pfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=1
X145 VOUT.t94 a_n2686_8422.t20 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X146 VDD.t27 a_n2686_12778.t55 a_n2511_10556.t13 VDD.t26 sky130_fd_pr__pfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X147 VOUT.t95 a_n2686_8422.t20 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X148 GND.t54 CS_BIAS.t53 VOUT.t13 GND.t7 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X149 VDD.t79 VDD.t77 VDD.t78 VDD.t40 sky130_fd_pr__pfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X150 VDD.t159 a_n7677_8299.t54 VOUT.t84 VDD.t158 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X151 VDD.t76 VDD.t74 VDD.t75 VDD.t63 sky130_fd_pr__pfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X152 GND.t92 GND.t89 GND.t91 GND.t90 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X153 VOUT.t83 a_n7677_8299.t55 VDD.t157 VDD.t156 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X154 GND.t8 CS_BIAS.t4 CS_BIAS.t5 GND.t7 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X155 a_n1455_n3928.t7 DIFFPAIR_BIAS.t10 GND.t37 GND.t36 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=2
X156 VOUT.t14 CS_BIAS.t54 GND.t55 GND.t24 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=2
X157 GND.t31 CS_BIAS.t55 VOUT.t6 GND.t4 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X158 a_n2511_10556.t12 a_n2686_12778.t56 VDD.t15 VDD.t14 sky130_fd_pr__pfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X159 VDD.t155 a_n7677_8299.t56 VOUT.t64 VDD.t154 sky130_fd_pr__pfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X160 CS_BIAS.t3 CS_BIAS.t2 GND.t176 GND.t160 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X161 VDD.t153 a_n7677_8299.t57 VOUT.t63 VDD.t135 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X162 a_n1455_n3928.t11 VN.t9 a_n7677_8299.t14 GND.t13 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X163 VOUT.t62 a_n7677_8299.t58 VDD.t152 VDD.t145 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X164 a_n2686_12778.t3 VP.t9 a_n1455_n3928.t5 GND.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X165 VOUT.t57 a_n7677_8299.t59 VDD.t151 VDD.t130 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X166 GND.t88 GND.t86 VN.t0 GND.t87 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X167 GND.t85 GND.t82 GND.t84 GND.t83 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X168 VDD.t73 VDD.t70 VDD.t72 VDD.t71 sky130_fd_pr__pfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X169 VDD.t150 a_n7677_8299.t60 VOUT.t56 VDD.t149 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X170 VDD.t69 VDD.t66 VDD.t68 VDD.t67 sky130_fd_pr__pfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=1
X171 VOUT.t96 a_n2686_8422.t20 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X172 VDD.t65 VDD.t62 VDD.t64 VDD.t63 sky130_fd_pr__pfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X173 VOUT.t55 a_n7677_8299.t61 VDD.t148 VDD.t121 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X174 a_n2511_10556.t4 a_n2686_12778.t23 a_n2686_12778.t24 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=1
X175 CS_BIAS.t1 CS_BIAS.t0 GND.t30 GND.t28 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X176 a_n7677_8299.t3 VN.t10 a_n1455_n3928.t10 GND.t27 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X177 VDD.t61 VDD.t58 VDD.t60 VDD.t59 sky130_fd_pr__pfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=1
X178 VOUT.t36 a_n7677_8299.t62 VDD.t147 VDD.t125 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X179 VOUT.t35 a_n7677_8299.t63 VDD.t146 VDD.t145 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X180 VDD.t144 a_n7677_8299.t64 VOUT.t34 VDD.t143 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X181 VOUT.t25 CS_BIAS.t56 GND.t166 GND.t61 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X182 a_n2686_12778.t6 VP.t10 a_n1455_n3928.t18 GND.t63 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X183 VDD.t57 VDD.t55 VDD.t56 VDD.t44 sky130_fd_pr__pfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X184 VDD.t142 a_n7677_8299.t65 VOUT.t33 VDD.t141 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X185 a_n2511_10556.t3 a_n2686_12778.t29 a_n2686_12778.t30 VDD.t32 sky130_fd_pr__pfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X186 a_n1455_n3928.t16 VP.t11 a_n2686_12778.t4 GND.t60 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X187 GND.t3 CS_BIAS.t57 VOUT.t0 GND.t2 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X188 VOUT.t32 a_n7677_8299.t66 VDD.t140 VDD.t139 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X189 a_n2686_8422.t8 a_n2686_12778.t57 a_n7677_8299.t4 VDD.t13 sky130_fd_pr__pfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X190 VOUT.t51 a_n7677_8299.t67 VDD.t138 VDD.t137 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X191 a_n1455_n3928.t1 DIFFPAIR_BIAS.t11 GND.t15 GND.t14 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=2
X192 VDD.t136 a_n7677_8299.t68 VOUT.t50 VDD.t135 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X193 GND.t26 CS_BIAS.t58 VOUT.t4 GND.t7 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X194 a_n2686_12778.t14 a_n2686_12778.t13 a_n2511_10556.t2 VDD.t197 sky130_fd_pr__pfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X195 VOUT.t72 a_n7677_8299.t69 VDD.t134 VDD.t132 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X196 VOUT.t97 a_n2686_8422.t20 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X197 VOUT.t71 a_n7677_8299.t70 VDD.t133 VDD.t132 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X198 VOUT.t91 CS_BIAS.t59 GND.t179 GND.t42 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X199 VOUT.t3 CS_BIAS.t60 GND.t25 GND.t24 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=2
X200 VOUT.t39 a_n7677_8299.t71 VDD.t131 VDD.t130 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X201 GND.t175 CS_BIAS.t61 VOUT.t89 GND.t48 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X202 GND.t81 GND.t78 GND.t80 GND.t79 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X203 VDD.t129 a_n7677_8299.t72 VOUT.t38 VDD.t123 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X204 a_n1455_n3928.t4 VP.t12 a_n2686_12778.t2 GND.t21 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X205 VDD.t54 VDD.t51 VDD.t53 VDD.t52 sky130_fd_pr__pfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=1
X206 VDD.t50 VDD.t47 VDD.t49 VDD.t48 sky130_fd_pr__pfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=1
X207 GND.t77 GND.t74 GND.t76 GND.t75 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X208 a_n2686_8422.t1 a_n2686_12778.t58 VDD.t19 VDD.t18 sky130_fd_pr__pfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=1
X209 VDD.t128 a_n7677_8299.t73 VOUT.t37 VDD.t127 sky130_fd_pr__pfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X210 VOUT.t70 a_n7677_8299.t74 VDD.t126 VDD.t125 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X211 DIFFPAIR_BIAS.t1 DIFFPAIR_BIAS.t0 GND.t23 GND.t22 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=2
X212 VOUT.t5 CS_BIAS.t62 GND.t29 GND.t28 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X213 a_n7677_8299.t2 VN.t11 a_n1455_n3928.t9 GND.t20 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X214 VDD.t124 a_n7677_8299.t75 VOUT.t69 VDD.t123 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X215 VOUT.t41 a_n7677_8299.t76 VDD.t122 VDD.t121 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X216 a_n2686_8422.t0 a_n2686_12778.t59 VDD.t24 VDD.t23 sky130_fd_pr__pfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X217 VDD.t120 a_n7677_8299.t77 VOUT.t40 VDD.t119 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X218 VDD.t46 VDD.t43 VDD.t45 VDD.t44 sky130_fd_pr__pfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X219 VOUT.t82 a_n7677_8299.t78 VDD.t118 VDD.t117 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X220 VP.t0 GND.t71 GND.t73 GND.t72 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X221 VOUT.t81 a_n7677_8299.t79 VDD.t116 VDD.t115 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X222 GND.t70 GND.t67 GND.t69 GND.t68 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X223 GND.t159 CS_BIAS.t63 VOUT.t20 GND.t57 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=2
X224 a_n2686_12778.t8 a_n2686_12778.t7 a_n2511_10556.t1 VDD.t4 sky130_fd_pr__pfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X225 a_n1455_n3928.t8 VN.t12 a_n7677_8299.t8 GND.t52 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X226 a_n2686_12778.t18 a_n2686_12778.t17 a_n2511_10556.t0 VDD.t1 sky130_fd_pr__pfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X227 VDD.t42 VDD.t39 VDD.t41 VDD.t40 sky130_fd_pr__pfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
R0 a_n7677_8299.n172 a_n7677_8299.t63 223.136
R1 a_n7677_8299.n160 a_n7677_8299.t30 223.136
R2 a_n7677_8299.n149 a_n7677_8299.t58 223.136
R3 a_n7677_8299.n133 a_n7677_8299.t20 223.136
R4 a_n7677_8299.n118 a_n7677_8299.t73 223.136
R5 a_n7677_8299.n104 a_n7677_8299.t40 223.136
R6 a_n7677_8299.n11 a_n7677_8299.t56 223.097
R7 a_n7677_8299.n10 a_n7677_8299.t47 223.097
R8 a_n7677_8299.n9 a_n7677_8299.t22 223.097
R9 a_n7677_8299.n142 a_n7677_8299.t74 207.983
R10 a_n7677_8299.n127 a_n7677_8299.t32 207.983
R11 a_n7677_8299.n113 a_n7677_8299.t62 207.983
R12 a_n7677_8299.n178 a_n7677_8299.t50 168.701
R13 a_n7677_8299.n177 a_n7677_8299.t64 168.701
R14 a_n7677_8299.n168 a_n7677_8299.t48 168.701
R15 a_n7677_8299.n174 a_n7677_8299.t46 168.701
R16 a_n7677_8299.n173 a_n7677_8299.t59 168.701
R17 a_n7677_8299.n169 a_n7677_8299.t72 168.701
R18 a_n7677_8299.n170 a_n7677_8299.t39 168.701
R19 a_n7677_8299.n171 a_n7677_8299.t51 168.701
R20 a_n7677_8299.n166 a_n7677_8299.t43 168.701
R21 a_n7677_8299.n165 a_n7677_8299.t24 168.701
R22 a_n7677_8299.n156 a_n7677_8299.t33 168.701
R23 a_n7677_8299.n162 a_n7677_8299.t31 168.701
R24 a_n7677_8299.n161 a_n7677_8299.t71 168.701
R25 a_n7677_8299.n157 a_n7677_8299.t41 168.701
R26 a_n7677_8299.n158 a_n7677_8299.t79 168.701
R27 a_n7677_8299.n159 a_n7677_8299.t53 168.701
R28 a_n7677_8299.n155 a_n7677_8299.t78 168.701
R29 a_n7677_8299.n154 a_n7677_8299.t52 168.701
R30 a_n7677_8299.n145 a_n7677_8299.t66 168.701
R31 a_n7677_8299.n153 a_n7677_8299.t60 168.701
R32 a_n7677_8299.n152 a_n7677_8299.t38 168.701
R33 a_n7677_8299.n146 a_n7677_8299.t75 168.701
R34 a_n7677_8299.n147 a_n7677_8299.t44 168.701
R35 a_n7677_8299.n148 a_n7677_8299.t26 168.701
R36 a_n7677_8299.n132 a_n7677_8299.t69 168.701
R37 a_n7677_8299.n131 a_n7677_8299.t35 168.701
R38 a_n7677_8299.n130 a_n7677_8299.t25 168.701
R39 a_n7677_8299.n136 a_n7677_8299.t77 168.701
R40 a_n7677_8299.n137 a_n7677_8299.t61 168.701
R41 a_n7677_8299.n23 a_n7677_8299.t45 168.701
R42 a_n7677_8299.n139 a_n7677_8299.t21 168.701
R43 a_n7677_8299.n140 a_n7677_8299.t68 168.701
R44 a_n7677_8299.n117 a_n7677_8299.t37 168.701
R45 a_n7677_8299.n116 a_n7677_8299.t65 168.701
R46 a_n7677_8299.n115 a_n7677_8299.t28 168.701
R47 a_n7677_8299.n121 a_n7677_8299.t49 168.701
R48 a_n7677_8299.n122 a_n7677_8299.t76 168.701
R49 a_n7677_8299.n25 a_n7677_8299.t27 168.701
R50 a_n7677_8299.n124 a_n7677_8299.t67 168.701
R51 a_n7677_8299.n125 a_n7677_8299.t29 168.701
R52 a_n7677_8299.n103 a_n7677_8299.t70 168.701
R53 a_n7677_8299.n102 a_n7677_8299.t34 168.701
R54 a_n7677_8299.n101 a_n7677_8299.t55 168.701
R55 a_n7677_8299.n107 a_n7677_8299.t23 168.701
R56 a_n7677_8299.n108 a_n7677_8299.t42 168.701
R57 a_n7677_8299.n27 a_n7677_8299.t54 168.701
R58 a_n7677_8299.n110 a_n7677_8299.t36 168.701
R59 a_n7677_8299.n111 a_n7677_8299.t57 168.701
R60 a_n7677_8299.n19 a_n7677_8299.n0 39.6376
R61 a_n7677_8299.n5 a_n7677_8299.n0 39.7274
R62 a_n7677_8299.n29 a_n7677_8299.n0 68.6201
R63 a_n7677_8299.n20 a_n7677_8299.n0 39.6373
R64 a_n7677_8299.n175 a_n7677_8299.n0 161.3
R65 a_n7677_8299.n1 a_n7677_8299.n176 161.3
R66 a_n7677_8299.n21 a_n7677_8299.n1 39.7274
R67 a_n7677_8299.n22 a_n7677_8299.n1 39.6376
R68 a_n7677_8299.n15 a_n7677_8299.n2 39.6376
R69 a_n7677_8299.n6 a_n7677_8299.n2 39.7274
R70 a_n7677_8299.n30 a_n7677_8299.n2 68.6201
R71 a_n7677_8299.n16 a_n7677_8299.n2 39.6373
R72 a_n7677_8299.n163 a_n7677_8299.n2 161.3
R73 a_n7677_8299.n3 a_n7677_8299.n164 161.3
R74 a_n7677_8299.n17 a_n7677_8299.n3 39.7274
R75 a_n7677_8299.n18 a_n7677_8299.n3 39.6376
R76 a_n7677_8299.n35 a_n7677_8299.n33 71.8318
R77 a_n7677_8299.n34 a_n7677_8299.n150 161.3
R78 a_n7677_8299.n151 a_n7677_8299.n34 161.3
R79 a_n7677_8299.n32 a_n7677_8299.n7 74.8341
R80 a_n7677_8299.n31 a_n7677_8299.n4 68.6201
R81 a_n7677_8299.n12 a_n7677_8299.n4 39.6373
R82 a_n7677_8299.n4 a_n7677_8299.n8 68.6201
R83 a_n7677_8299.n13 a_n7677_8299.n4 39.7274
R84 a_n7677_8299.n14 a_n7677_8299.n4 39.6376
R85 a_n7677_8299.n141 a_n7677_8299.n53 161.3
R86 a_n7677_8299.n50 a_n7677_8299.n53 161.3
R87 a_n7677_8299.n52 a_n7677_8299.n51 71.4497
R88 a_n7677_8299.n49 a_n7677_8299.n48 68.7078
R89 a_n7677_8299.n24 a_n7677_8299.n23 11.426
R90 a_n7677_8299.n47 a_n7677_8299.n24 74.9385
R91 a_n7677_8299.n138 a_n7677_8299.n46 161.3
R92 a_n7677_8299.n43 a_n7677_8299.n46 161.3
R93 a_n7677_8299.n45 a_n7677_8299.n44 71.6402
R94 a_n7677_8299.n42 a_n7677_8299.n41 68.6201
R95 a_n7677_8299.n38 a_n7677_8299.n40 74.8341
R96 a_n7677_8299.n135 a_n7677_8299.n39 161.3
R97 a_n7677_8299.n39 a_n7677_8299.n134 161.3
R98 a_n7677_8299.n37 a_n7677_8299.n36 71.8318
R99 a_n7677_8299.n126 a_n7677_8299.n71 161.3
R100 a_n7677_8299.n68 a_n7677_8299.n71 161.3
R101 a_n7677_8299.n70 a_n7677_8299.n69 71.4497
R102 a_n7677_8299.n67 a_n7677_8299.n66 68.7078
R103 a_n7677_8299.n26 a_n7677_8299.n25 11.426
R104 a_n7677_8299.n65 a_n7677_8299.n26 74.9385
R105 a_n7677_8299.n123 a_n7677_8299.n64 161.3
R106 a_n7677_8299.n61 a_n7677_8299.n64 161.3
R107 a_n7677_8299.n63 a_n7677_8299.n62 71.6402
R108 a_n7677_8299.n60 a_n7677_8299.n59 68.6201
R109 a_n7677_8299.n56 a_n7677_8299.n58 74.8341
R110 a_n7677_8299.n120 a_n7677_8299.n57 161.3
R111 a_n7677_8299.n57 a_n7677_8299.n119 161.3
R112 a_n7677_8299.n55 a_n7677_8299.n54 71.8318
R113 a_n7677_8299.n112 a_n7677_8299.n89 161.3
R114 a_n7677_8299.n86 a_n7677_8299.n89 161.3
R115 a_n7677_8299.n88 a_n7677_8299.n87 71.4497
R116 a_n7677_8299.n85 a_n7677_8299.n84 68.7078
R117 a_n7677_8299.n28 a_n7677_8299.n27 11.426
R118 a_n7677_8299.n83 a_n7677_8299.n28 74.9385
R119 a_n7677_8299.n109 a_n7677_8299.n82 161.3
R120 a_n7677_8299.n79 a_n7677_8299.n82 161.3
R121 a_n7677_8299.n81 a_n7677_8299.n80 71.6402
R122 a_n7677_8299.n78 a_n7677_8299.n77 68.6201
R123 a_n7677_8299.n74 a_n7677_8299.n76 74.8341
R124 a_n7677_8299.n106 a_n7677_8299.n75 161.3
R125 a_n7677_8299.n75 a_n7677_8299.n105 161.3
R126 a_n7677_8299.n73 a_n7677_8299.n72 71.8318
R127 a_n7677_8299.n97 a_n7677_8299.n95 109.74
R128 a_n7677_8299.n92 a_n7677_8299.n90 109.74
R129 a_n7677_8299.n99 a_n7677_8299.n98 109.166
R130 a_n7677_8299.n97 a_n7677_8299.n96 109.166
R131 a_n7677_8299.n92 a_n7677_8299.n91 109.166
R132 a_n7677_8299.n94 a_n7677_8299.n93 109.166
R133 a_n7677_8299.n188 a_n7677_8299.n187 81.2193
R134 a_n7677_8299.n183 a_n7677_8299.n182 81.2191
R135 a_n7677_8299.n187 a_n7677_8299.n186 81.219
R136 a_n7677_8299.n185 a_n7677_8299.n184 80.9324
R137 a_n7677_8299.n1 a_n7677_8299.n11 43.6696
R138 a_n7677_8299.n3 a_n7677_8299.n10 43.6696
R139 a_n7677_8299.n4 a_n7677_8299.n9 43.6696
R140 a_n7677_8299.n143 a_n7677_8299.n142 80.6037
R141 a_n7677_8299.n128 a_n7677_8299.n127 80.6037
R142 a_n7677_8299.n114 a_n7677_8299.n113 80.6037
R143 a_n7677_8299.n176 a_n7677_8299.n175 56.5617
R144 a_n7677_8299.n29 a_n7677_8299.n169 48.4088
R145 a_n7677_8299.n164 a_n7677_8299.n163 56.5617
R146 a_n7677_8299.n30 a_n7677_8299.n157 48.4088
R147 a_n7677_8299.n31 a_n7677_8299.n146 48.4088
R148 a_n7677_8299.n136 a_n7677_8299.n42 40.5394
R149 a_n7677_8299.n24 a_n7677_8299.n138 67.9872
R150 a_n7677_8299.n121 a_n7677_8299.n60 40.5394
R151 a_n7677_8299.n26 a_n7677_8299.n123 67.9872
R152 a_n7677_8299.n107 a_n7677_8299.n78 40.5394
R153 a_n7677_8299.n28 a_n7677_8299.n109 67.9872
R154 a_n7677_8299.n177 a_n7677_8299.n21 51.9316
R155 a_n7677_8299.n165 a_n7677_8299.n17 51.9316
R156 a_n7677_8299.n154 a_n7677_8299.n13 51.9316
R157 a_n7677_8299.n40 a_n7677_8299.n135 67.7116
R158 a_n7677_8299.n139 a_n7677_8299.n49 39.872
R159 a_n7677_8299.n58 a_n7677_8299.n120 67.7116
R160 a_n7677_8299.n124 a_n7677_8299.n67 39.872
R161 a_n7677_8299.n76 a_n7677_8299.n106 67.7116
R162 a_n7677_8299.n110 a_n7677_8299.n85 39.872
R163 a_n7677_8299.n142 a_n7677_8299.n141 55.824
R164 a_n7677_8299.n127 a_n7677_8299.n126 55.824
R165 a_n7677_8299.n113 a_n7677_8299.n112 55.824
R166 a_n7677_8299.n172 a_n7677_8299.n171 47.1841
R167 a_n7677_8299.n160 a_n7677_8299.n159 47.1841
R168 a_n7677_8299.n149 a_n7677_8299.n148 47.1841
R169 a_n7677_8299.n133 a_n7677_8299.n132 47.1841
R170 a_n7677_8299.n118 a_n7677_8299.n117 47.1841
R171 a_n7677_8299.n104 a_n7677_8299.n103 47.1841
R172 a_n7677_8299.n36 a_n7677_8299.n133 43.9713
R173 a_n7677_8299.n54 a_n7677_8299.n118 43.9713
R174 a_n7677_8299.n72 a_n7677_8299.n104 43.9713
R175 a_n7677_8299.n0 a_n7677_8299.n172 43.9713
R176 a_n7677_8299.n2 a_n7677_8299.n160 43.9713
R177 a_n7677_8299.n33 a_n7677_8299.n149 43.9713
R178 a_n7677_8299.n177 a_n7677_8299.n22 41.2665
R179 a_n7677_8299.n165 a_n7677_8299.n18 41.2665
R180 a_n7677_8299.n154 a_n7677_8299.n14 41.2665
R181 a_n7677_8299.n150 a_n7677_8299.n35 59.1846
R182 a_n7677_8299.n134 a_n7677_8299.n37 59.1846
R183 a_n7677_8299.n51 a_n7677_8299.n50 58.0115
R184 a_n7677_8299.n119 a_n7677_8299.n55 59.1846
R185 a_n7677_8299.n69 a_n7677_8299.n68 58.0115
R186 a_n7677_8299.n105 a_n7677_8299.n73 59.1846
R187 a_n7677_8299.n87 a_n7677_8299.n86 58.0115
R188 a_n7677_8299.n173 a_n7677_8299.n20 40.5378
R189 a_n7677_8299.n161 a_n7677_8299.n16 40.5378
R190 a_n7677_8299.n152 a_n7677_8299.n12 40.5378
R191 a_n7677_8299.n44 a_n7677_8299.n43 58.5991
R192 a_n7677_8299.n62 a_n7677_8299.n61 58.5991
R193 a_n7677_8299.n80 a_n7677_8299.n79 58.5991
R194 a_n7677_8299.n19 a_n7677_8299.n171 39.8067
R195 a_n7677_8299.n15 a_n7677_8299.n159 39.8067
R196 a_n7677_8299.n35 a_n7677_8299.n148 25.2628
R197 a_n7677_8299.n187 a_n7677_8299.n185 31.3366
R198 a_n7677_8299.n100 a_n7677_8299.n94 27.4144
R199 a_n7677_8299.n5 a_n7677_8299.n170 51.931
R200 a_n7677_8299.n6 a_n7677_8299.n158 51.931
R201 a_n7677_8299.n32 a_n7677_8299.n151 67.7116
R202 a_n7677_8299.n130 a_n7677_8299.n40 11.8807
R203 a_n7677_8299.n49 a_n7677_8299.n23 48.9635
R204 a_n7677_8299.n115 a_n7677_8299.n58 11.8807
R205 a_n7677_8299.n67 a_n7677_8299.n25 48.9635
R206 a_n7677_8299.n101 a_n7677_8299.n76 11.8807
R207 a_n7677_8299.n85 a_n7677_8299.n27 48.9635
R208 a_n7677_8299.n176 a_n7677_8299.n168 24.3464
R209 a_n7677_8299.n164 a_n7677_8299.n156 24.3464
R210 a_n7677_8299.n8 a_n7677_8299.n145 48.4088
R211 a_n7677_8299.n42 a_n7677_8299.n130 48.4088
R212 a_n7677_8299.n60 a_n7677_8299.n115 48.4088
R213 a_n7677_8299.n78 a_n7677_8299.n101 48.4088
R214 a_n7677_8299.n100 a_n7677_8299.n99 17.7829
R215 a_n7677_8299.n11 a_n7677_8299.n178 47.213
R216 a_n7677_8299.n10 a_n7677_8299.n166 47.213
R217 a_n7677_8299.n9 a_n7677_8299.n155 47.213
R218 a_n7677_8299.n141 a_n7677_8299.n140 16.9689
R219 a_n7677_8299.n126 a_n7677_8299.n125 16.9689
R220 a_n7677_8299.n112 a_n7677_8299.n111 16.9689
R221 a_n7677_8299.n175 a_n7677_8299.n174 16.477
R222 a_n7677_8299.n173 a_n7677_8299.n29 40.5394
R223 a_n7677_8299.n163 a_n7677_8299.n162 16.477
R224 a_n7677_8299.n161 a_n7677_8299.n30 40.5394
R225 a_n7677_8299.n8 a_n7677_8299.n153 40.5394
R226 a_n7677_8299.n152 a_n7677_8299.n31 40.5394
R227 a_n7677_8299.n138 a_n7677_8299.n137 16.477
R228 a_n7677_8299.n123 a_n7677_8299.n122 16.477
R229 a_n7677_8299.n109 a_n7677_8299.n108 16.477
R230 a_n7677_8299.n151 a_n7677_8299.n147 15.9852
R231 a_n7677_8299.n135 a_n7677_8299.n131 15.9852
R232 a_n7677_8299.n120 a_n7677_8299.n116 15.9852
R233 a_n7677_8299.n106 a_n7677_8299.n102 15.9852
R234 a_n7677_8299.n183 a_n7677_8299.n181 12.361
R235 a_n7677_8299.n181 a_n7677_8299.n100 11.4887
R236 a_n7677_8299.n167 a_n7677_8299.n4 8.76042
R237 a_n7677_8299.n129 a_n7677_8299.n114 8.76042
R238 a_n7677_8299.n19 a_n7677_8299.n170 41.266
R239 a_n7677_8299.n15 a_n7677_8299.n158 41.266
R240 a_n7677_8299.n150 a_n7677_8299.n147 8.60764
R241 a_n7677_8299.n134 a_n7677_8299.n131 8.60764
R242 a_n7677_8299.n51 a_n7677_8299.n139 27.0108
R243 a_n7677_8299.n119 a_n7677_8299.n116 8.60764
R244 a_n7677_8299.n69 a_n7677_8299.n124 27.0108
R245 a_n7677_8299.n105 a_n7677_8299.n102 8.60764
R246 a_n7677_8299.n87 a_n7677_8299.n110 27.0108
R247 a_n7677_8299.n174 a_n7677_8299.n20 40.5373
R248 a_n7677_8299.n162 a_n7677_8299.n16 40.5373
R249 a_n7677_8299.n153 a_n7677_8299.n12 40.5373
R250 a_n7677_8299.n44 a_n7677_8299.n136 26.1378
R251 a_n7677_8299.n137 a_n7677_8299.n43 8.11581
R252 a_n7677_8299.n62 a_n7677_8299.n121 26.1378
R253 a_n7677_8299.n122 a_n7677_8299.n61 8.11581
R254 a_n7677_8299.n80 a_n7677_8299.n107 26.1378
R255 a_n7677_8299.n108 a_n7677_8299.n79 8.11581
R256 a_n7677_8299.n178 a_n7677_8299.n22 39.8062
R257 a_n7677_8299.n166 a_n7677_8299.n18 39.8062
R258 a_n7677_8299.n155 a_n7677_8299.n14 39.8062
R259 a_n7677_8299.n37 a_n7677_8299.n132 25.2628
R260 a_n7677_8299.n140 a_n7677_8299.n50 7.62397
R261 a_n7677_8299.n55 a_n7677_8299.n117 25.2628
R262 a_n7677_8299.n125 a_n7677_8299.n68 7.62397
R263 a_n7677_8299.n73 a_n7677_8299.n103 25.2628
R264 a_n7677_8299.n111 a_n7677_8299.n86 7.62397
R265 a_n7677_8299.n180 a_n7677_8299.n144 5.74635
R266 a_n7677_8299.n180 a_n7677_8299.n179 5.5455
R267 a_n7677_8299.n98 a_n7677_8299.t16 5.418
R268 a_n7677_8299.n98 a_n7677_8299.t6 5.418
R269 a_n7677_8299.n96 a_n7677_8299.t11 5.418
R270 a_n7677_8299.n96 a_n7677_8299.t19 5.418
R271 a_n7677_8299.n95 a_n7677_8299.t10 5.418
R272 a_n7677_8299.n95 a_n7677_8299.t17 5.418
R273 a_n7677_8299.n90 a_n7677_8299.t4 5.418
R274 a_n7677_8299.n90 a_n7677_8299.t5 5.418
R275 a_n7677_8299.n91 a_n7677_8299.t1 5.418
R276 a_n7677_8299.n91 a_n7677_8299.t18 5.418
R277 a_n7677_8299.n93 a_n7677_8299.t7 5.418
R278 a_n7677_8299.n93 a_n7677_8299.t9 5.418
R279 a_n7677_8299.n179 a_n7677_8299.n1 5.06913
R280 a_n7677_8299.n167 a_n7677_8299.n3 5.06913
R281 a_n7677_8299.n144 a_n7677_8299.n143 5.06913
R282 a_n7677_8299.n129 a_n7677_8299.n128 5.06913
R283 a_n7677_8299.n179 a_n7677_8299.n167 3.69179
R284 a_n7677_8299.n144 a_n7677_8299.n129 3.69179
R285 a_n7677_8299.n181 a_n7677_8299.n180 3.4105
R286 a_n7677_8299.n186 a_n7677_8299.t14 2.82907
R287 a_n7677_8299.n186 a_n7677_8299.t3 2.82907
R288 a_n7677_8299.n184 a_n7677_8299.t13 2.82907
R289 a_n7677_8299.n184 a_n7677_8299.t12 2.82907
R290 a_n7677_8299.n182 a_n7677_8299.t8 2.82907
R291 a_n7677_8299.n182 a_n7677_8299.t2 2.82907
R292 a_n7677_8299.n188 a_n7677_8299.t15 2.82907
R293 a_n7677_8299.t0 a_n7677_8299.n188 2.82907
R294 a_n7677_8299.n99 a_n7677_8299.n97 0.573776
R295 a_n7677_8299.n94 a_n7677_8299.n92 0.573776
R296 a_n7677_8299.n75 a_n7677_8299.n72 0.568682
R297 a_n7677_8299.n57 a_n7677_8299.n54 0.568682
R298 a_n7677_8299.n39 a_n7677_8299.n36 0.568682
R299 a_n7677_8299.n89 a_n7677_8299.n88 0.379288
R300 a_n7677_8299.n88 a_n7677_8299.n84 0.379288
R301 a_n7677_8299.n84 a_n7677_8299.n83 0.379288
R302 a_n7677_8299.n83 a_n7677_8299.n82 0.379288
R303 a_n7677_8299.n82 a_n7677_8299.n81 0.379288
R304 a_n7677_8299.n81 a_n7677_8299.n77 0.379288
R305 a_n7677_8299.n77 a_n7677_8299.n74 0.379288
R306 a_n7677_8299.n75 a_n7677_8299.n74 0.379288
R307 a_n7677_8299.n71 a_n7677_8299.n70 0.379288
R308 a_n7677_8299.n70 a_n7677_8299.n66 0.379288
R309 a_n7677_8299.n66 a_n7677_8299.n65 0.379288
R310 a_n7677_8299.n65 a_n7677_8299.n64 0.379288
R311 a_n7677_8299.n64 a_n7677_8299.n63 0.379288
R312 a_n7677_8299.n63 a_n7677_8299.n59 0.379288
R313 a_n7677_8299.n59 a_n7677_8299.n56 0.379288
R314 a_n7677_8299.n57 a_n7677_8299.n56 0.379288
R315 a_n7677_8299.n53 a_n7677_8299.n52 0.379288
R316 a_n7677_8299.n52 a_n7677_8299.n48 0.379288
R317 a_n7677_8299.n48 a_n7677_8299.n47 0.379288
R318 a_n7677_8299.n47 a_n7677_8299.n46 0.379288
R319 a_n7677_8299.n46 a_n7677_8299.n45 0.379288
R320 a_n7677_8299.n45 a_n7677_8299.n41 0.379288
R321 a_n7677_8299.n41 a_n7677_8299.n38 0.379288
R322 a_n7677_8299.n39 a_n7677_8299.n38 0.379288
R323 a_n7677_8299.n34 a_n7677_8299.n33 0.379288
R324 a_n7677_8299.n34 a_n7677_8299.n7 0.379288
R325 a_n7677_8299.n185 a_n7677_8299.n183 0.287138
R326 a_n7677_8299.n143 a_n7677_8299.n53 0.285035
R327 a_n7677_8299.n128 a_n7677_8299.n71 0.285035
R328 a_n7677_8299.n114 a_n7677_8299.n89 0.285035
R329 a_n7677_8299.n168 a_n7677_8299.n21 28.5572
R330 a_n7677_8299.n5 a_n7677_8299.n169 28.5577
R331 a_n7677_8299.n156 a_n7677_8299.n17 28.5572
R332 a_n7677_8299.n6 a_n7677_8299.n157 28.5577
R333 a_n7677_8299.n145 a_n7677_8299.n13 28.5572
R334 a_n7677_8299.n32 a_n7677_8299.n146 11.8807
R335 a_n7677_8299.n3 a_n7677_8299.n2 3.88352
R336 a_n7677_8299.n1 a_n7677_8299.n0 3.88352
R337 a_n7677_8299.n4 a_n7677_8299.n7 3.12594
R338 VOUT.n202 VOUT.n200 102.66
R339 VOUT.n192 VOUT.n190 102.66
R340 VOUT.n183 VOUT.n181 102.66
R341 VOUT.n21 VOUT.n19 102.66
R342 VOUT.n11 VOUT.n9 102.66
R343 VOUT.n2 VOUT.n0 102.66
R344 VOUT.n206 VOUT.n205 102.088
R345 VOUT.n204 VOUT.n203 102.088
R346 VOUT.n202 VOUT.n201 102.088
R347 VOUT.n198 VOUT.n197 102.088
R348 VOUT.n196 VOUT.n195 102.088
R349 VOUT.n194 VOUT.n193 102.088
R350 VOUT.n192 VOUT.n191 102.088
R351 VOUT.n189 VOUT.n188 102.088
R352 VOUT.n187 VOUT.n186 102.088
R353 VOUT.n185 VOUT.n184 102.088
R354 VOUT.n183 VOUT.n182 102.088
R355 VOUT.n21 VOUT.n20 102.088
R356 VOUT.n23 VOUT.n22 102.088
R357 VOUT.n25 VOUT.n24 102.088
R358 VOUT.n27 VOUT.n26 102.088
R359 VOUT.n11 VOUT.n10 102.088
R360 VOUT.n13 VOUT.n12 102.088
R361 VOUT.n15 VOUT.n14 102.088
R362 VOUT.n17 VOUT.n16 102.088
R363 VOUT.n2 VOUT.n1 102.088
R364 VOUT.n4 VOUT.n3 102.088
R365 VOUT.n6 VOUT.n5 102.088
R366 VOUT.n8 VOUT.n7 102.088
R367 VOUT.n208 VOUT.n207 102.088
R368 VOUT.n220 VOUT.n218 85.0679
R369 VOUT.n213 VOUT.n211 85.0679
R370 VOUT.n236 VOUT.n234 85.0679
R371 VOUT.n229 VOUT.n227 85.0679
R372 VOUT.n224 VOUT.n223 84.0635
R373 VOUT.n222 VOUT.n221 84.0635
R374 VOUT.n220 VOUT.n219 84.0635
R375 VOUT.n217 VOUT.n216 84.0635
R376 VOUT.n215 VOUT.n214 84.0635
R377 VOUT.n213 VOUT.n212 84.0635
R378 VOUT.n236 VOUT.n235 84.0635
R379 VOUT.n238 VOUT.n237 84.0635
R380 VOUT.n240 VOUT.n239 84.0635
R381 VOUT.n229 VOUT.n228 84.0635
R382 VOUT.n231 VOUT.n230 84.0635
R383 VOUT.n233 VOUT.n232 84.0635
R384 VOUT.n226 VOUT.n210 8.45563
R385 VOUT.n199 VOUT.n189 7.37442
R386 VOUT.n18 VOUT.n8 7.37442
R387 VOUT.n225 VOUT.n217 7.37334
R388 VOUT.n241 VOUT.n233 7.37334
R389 VOUT.n226 VOUT.n225 6.2036
R390 VOUT.n242 VOUT.n241 6.2036
R391 VOUT.n225 VOUT.n224 5.46817
R392 VOUT.n241 VOUT.n240 5.46817
R393 VOUT.n209 VOUT.n208 5.25266
R394 VOUT.n199 VOUT.n198 5.25266
R395 VOUT.n28 VOUT.n27 5.25266
R396 VOUT.n18 VOUT.n17 5.25266
R397 VOUT.n210 VOUT.n209 4.90511
R398 VOUT.n29 VOUT.n28 4.90511
R399 VOUT.n243 VOUT.n29 4.83577
R400 VOUT.n207 VOUT.t58 4.64407
R401 VOUT.n207 VOUT.t62 4.64407
R402 VOUT.n205 VOUT.t69 4.64407
R403 VOUT.n205 VOUT.t30 4.64407
R404 VOUT.n203 VOUT.t56 4.64407
R405 VOUT.n203 VOUT.t77 4.64407
R406 VOUT.n201 VOUT.t86 4.64407
R407 VOUT.n201 VOUT.t32 4.64407
R408 VOUT.n200 VOUT.t52 4.64407
R409 VOUT.n200 VOUT.t82 4.64407
R410 VOUT.n197 VOUT.t85 4.64407
R411 VOUT.n197 VOUT.t73 4.64407
R412 VOUT.n195 VOUT.t43 4.64407
R413 VOUT.n195 VOUT.t81 4.64407
R414 VOUT.n193 VOUT.t49 4.64407
R415 VOUT.n193 VOUT.t39 4.64407
R416 VOUT.n191 VOUT.t60 4.64407
R417 VOUT.n191 VOUT.t47 4.64407
R418 VOUT.n190 VOUT.t68 4.64407
R419 VOUT.n190 VOUT.t31 4.64407
R420 VOUT.n188 VOUT.t87 4.64407
R421 VOUT.n188 VOUT.t35 4.64407
R422 VOUT.n186 VOUT.t38 4.64407
R423 VOUT.n186 VOUT.t45 4.64407
R424 VOUT.n184 VOUT.t28 4.64407
R425 VOUT.n184 VOUT.t57 4.64407
R426 VOUT.n182 VOUT.t34 4.64407
R427 VOUT.n182 VOUT.t67 4.64407
R428 VOUT.n181 VOUT.t64 4.64407
R429 VOUT.n181 VOUT.t65 4.64407
R430 VOUT.n19 VOUT.t63 4.64407
R431 VOUT.n19 VOUT.t36 4.64407
R432 VOUT.n20 VOUT.t84 4.64407
R433 VOUT.n20 VOUT.t79 4.64407
R434 VOUT.n22 VOUT.t61 4.64407
R435 VOUT.n22 VOUT.t42 4.64407
R436 VOUT.n24 VOUT.t46 4.64407
R437 VOUT.n24 VOUT.t83 4.64407
R438 VOUT.n26 VOUT.t44 4.64407
R439 VOUT.n26 VOUT.t71 4.64407
R440 VOUT.n9 VOUT.t74 4.64407
R441 VOUT.n9 VOUT.t48 4.64407
R442 VOUT.n10 VOUT.t76 4.64407
R443 VOUT.n10 VOUT.t51 4.64407
R444 VOUT.n12 VOUT.t66 4.64407
R445 VOUT.n12 VOUT.t41 4.64407
R446 VOUT.n14 VOUT.t33 4.64407
R447 VOUT.n14 VOUT.t75 4.64407
R448 VOUT.n16 VOUT.t37 4.64407
R449 VOUT.n16 VOUT.t78 4.64407
R450 VOUT.n0 VOUT.t50 4.64407
R451 VOUT.n0 VOUT.t70 4.64407
R452 VOUT.n1 VOUT.t29 4.64407
R453 VOUT.n1 VOUT.t53 4.64407
R454 VOUT.n3 VOUT.t40 4.64407
R455 VOUT.n3 VOUT.t55 4.64407
R456 VOUT.n5 VOUT.t80 4.64407
R457 VOUT.n5 VOUT.t59 4.64407
R458 VOUT.n7 VOUT.t54 4.64407
R459 VOUT.n7 VOUT.t72 4.64407
R460 VOUT.n120 VOUT.n73 4.5005
R461 VOUT.n89 VOUT.n73 4.5005
R462 VOUT.n84 VOUT.n68 4.5005
R463 VOUT.n84 VOUT.n70 4.5005
R464 VOUT.n84 VOUT.n67 4.5005
R465 VOUT.n84 VOUT.n71 4.5005
R466 VOUT.n84 VOUT.n66 4.5005
R467 VOUT.n84 VOUT.t97 4.5005
R468 VOUT.n84 VOUT.n65 4.5005
R469 VOUT.n84 VOUT.n72 4.5005
R470 VOUT.n84 VOUT.n73 4.5005
R471 VOUT.n82 VOUT.n68 4.5005
R472 VOUT.n82 VOUT.n70 4.5005
R473 VOUT.n82 VOUT.n67 4.5005
R474 VOUT.n82 VOUT.n71 4.5005
R475 VOUT.n82 VOUT.n66 4.5005
R476 VOUT.n82 VOUT.t97 4.5005
R477 VOUT.n82 VOUT.n65 4.5005
R478 VOUT.n82 VOUT.n72 4.5005
R479 VOUT.n82 VOUT.n73 4.5005
R480 VOUT.n81 VOUT.n68 4.5005
R481 VOUT.n81 VOUT.n70 4.5005
R482 VOUT.n81 VOUT.n67 4.5005
R483 VOUT.n81 VOUT.n71 4.5005
R484 VOUT.n81 VOUT.n66 4.5005
R485 VOUT.n81 VOUT.t97 4.5005
R486 VOUT.n81 VOUT.n65 4.5005
R487 VOUT.n81 VOUT.n72 4.5005
R488 VOUT.n81 VOUT.n73 4.5005
R489 VOUT.n166 VOUT.n68 4.5005
R490 VOUT.n166 VOUT.n70 4.5005
R491 VOUT.n166 VOUT.n67 4.5005
R492 VOUT.n166 VOUT.n71 4.5005
R493 VOUT.n166 VOUT.n66 4.5005
R494 VOUT.n166 VOUT.t97 4.5005
R495 VOUT.n166 VOUT.n65 4.5005
R496 VOUT.n166 VOUT.n72 4.5005
R497 VOUT.n166 VOUT.n73 4.5005
R498 VOUT.n164 VOUT.n68 4.5005
R499 VOUT.n164 VOUT.n70 4.5005
R500 VOUT.n164 VOUT.n67 4.5005
R501 VOUT.n164 VOUT.n71 4.5005
R502 VOUT.n164 VOUT.n66 4.5005
R503 VOUT.n164 VOUT.t97 4.5005
R504 VOUT.n164 VOUT.n65 4.5005
R505 VOUT.n164 VOUT.n72 4.5005
R506 VOUT.n162 VOUT.n68 4.5005
R507 VOUT.n162 VOUT.n70 4.5005
R508 VOUT.n162 VOUT.n67 4.5005
R509 VOUT.n162 VOUT.n71 4.5005
R510 VOUT.n162 VOUT.n66 4.5005
R511 VOUT.n162 VOUT.t97 4.5005
R512 VOUT.n162 VOUT.n65 4.5005
R513 VOUT.n162 VOUT.n72 4.5005
R514 VOUT.n92 VOUT.n68 4.5005
R515 VOUT.n92 VOUT.n70 4.5005
R516 VOUT.n92 VOUT.n67 4.5005
R517 VOUT.n92 VOUT.n71 4.5005
R518 VOUT.n92 VOUT.n66 4.5005
R519 VOUT.n92 VOUT.t97 4.5005
R520 VOUT.n92 VOUT.n65 4.5005
R521 VOUT.n92 VOUT.n72 4.5005
R522 VOUT.n92 VOUT.n73 4.5005
R523 VOUT.n91 VOUT.n68 4.5005
R524 VOUT.n91 VOUT.n70 4.5005
R525 VOUT.n91 VOUT.n67 4.5005
R526 VOUT.n91 VOUT.n71 4.5005
R527 VOUT.n91 VOUT.n66 4.5005
R528 VOUT.n91 VOUT.t97 4.5005
R529 VOUT.n91 VOUT.n65 4.5005
R530 VOUT.n91 VOUT.n72 4.5005
R531 VOUT.n91 VOUT.n73 4.5005
R532 VOUT.n95 VOUT.n68 4.5005
R533 VOUT.n95 VOUT.n70 4.5005
R534 VOUT.n95 VOUT.n67 4.5005
R535 VOUT.n95 VOUT.n71 4.5005
R536 VOUT.n95 VOUT.n66 4.5005
R537 VOUT.n95 VOUT.t97 4.5005
R538 VOUT.n95 VOUT.n65 4.5005
R539 VOUT.n95 VOUT.n72 4.5005
R540 VOUT.n95 VOUT.n73 4.5005
R541 VOUT.n94 VOUT.n68 4.5005
R542 VOUT.n94 VOUT.n70 4.5005
R543 VOUT.n94 VOUT.n67 4.5005
R544 VOUT.n94 VOUT.n71 4.5005
R545 VOUT.n94 VOUT.n66 4.5005
R546 VOUT.n94 VOUT.t97 4.5005
R547 VOUT.n94 VOUT.n65 4.5005
R548 VOUT.n94 VOUT.n72 4.5005
R549 VOUT.n94 VOUT.n73 4.5005
R550 VOUT.n77 VOUT.n68 4.5005
R551 VOUT.n77 VOUT.n70 4.5005
R552 VOUT.n77 VOUT.n67 4.5005
R553 VOUT.n77 VOUT.n71 4.5005
R554 VOUT.n77 VOUT.n66 4.5005
R555 VOUT.n77 VOUT.t97 4.5005
R556 VOUT.n77 VOUT.n65 4.5005
R557 VOUT.n77 VOUT.n72 4.5005
R558 VOUT.n77 VOUT.n73 4.5005
R559 VOUT.n169 VOUT.n68 4.5005
R560 VOUT.n169 VOUT.n70 4.5005
R561 VOUT.n169 VOUT.n67 4.5005
R562 VOUT.n169 VOUT.n71 4.5005
R563 VOUT.n169 VOUT.n66 4.5005
R564 VOUT.n169 VOUT.t97 4.5005
R565 VOUT.n169 VOUT.n65 4.5005
R566 VOUT.n169 VOUT.n72 4.5005
R567 VOUT.n169 VOUT.n73 4.5005
R568 VOUT.n156 VOUT.n127 4.5005
R569 VOUT.n156 VOUT.n133 4.5005
R570 VOUT.n114 VOUT.n103 4.5005
R571 VOUT.n114 VOUT.n105 4.5005
R572 VOUT.n114 VOUT.n102 4.5005
R573 VOUT.n114 VOUT.n106 4.5005
R574 VOUT.n114 VOUT.n101 4.5005
R575 VOUT.n114 VOUT.t94 4.5005
R576 VOUT.n114 VOUT.n100 4.5005
R577 VOUT.n114 VOUT.n107 4.5005
R578 VOUT.n156 VOUT.n114 4.5005
R579 VOUT.n135 VOUT.n103 4.5005
R580 VOUT.n135 VOUT.n105 4.5005
R581 VOUT.n135 VOUT.n102 4.5005
R582 VOUT.n135 VOUT.n106 4.5005
R583 VOUT.n135 VOUT.n101 4.5005
R584 VOUT.n135 VOUT.t94 4.5005
R585 VOUT.n135 VOUT.n100 4.5005
R586 VOUT.n135 VOUT.n107 4.5005
R587 VOUT.n156 VOUT.n135 4.5005
R588 VOUT.n113 VOUT.n103 4.5005
R589 VOUT.n113 VOUT.n105 4.5005
R590 VOUT.n113 VOUT.n102 4.5005
R591 VOUT.n113 VOUT.n106 4.5005
R592 VOUT.n113 VOUT.n101 4.5005
R593 VOUT.n113 VOUT.t94 4.5005
R594 VOUT.n113 VOUT.n100 4.5005
R595 VOUT.n113 VOUT.n107 4.5005
R596 VOUT.n156 VOUT.n113 4.5005
R597 VOUT.n137 VOUT.n103 4.5005
R598 VOUT.n137 VOUT.n105 4.5005
R599 VOUT.n137 VOUT.n102 4.5005
R600 VOUT.n137 VOUT.n106 4.5005
R601 VOUT.n137 VOUT.n101 4.5005
R602 VOUT.n137 VOUT.t94 4.5005
R603 VOUT.n137 VOUT.n100 4.5005
R604 VOUT.n137 VOUT.n107 4.5005
R605 VOUT.n156 VOUT.n137 4.5005
R606 VOUT.n103 VOUT.n98 4.5005
R607 VOUT.n105 VOUT.n98 4.5005
R608 VOUT.n102 VOUT.n98 4.5005
R609 VOUT.n106 VOUT.n98 4.5005
R610 VOUT.n101 VOUT.n98 4.5005
R611 VOUT.t94 VOUT.n98 4.5005
R612 VOUT.n100 VOUT.n98 4.5005
R613 VOUT.n107 VOUT.n98 4.5005
R614 VOUT.n159 VOUT.n103 4.5005
R615 VOUT.n159 VOUT.n105 4.5005
R616 VOUT.n159 VOUT.n102 4.5005
R617 VOUT.n159 VOUT.n106 4.5005
R618 VOUT.n159 VOUT.n101 4.5005
R619 VOUT.n159 VOUT.t94 4.5005
R620 VOUT.n159 VOUT.n100 4.5005
R621 VOUT.n159 VOUT.n107 4.5005
R622 VOUT.n157 VOUT.n103 4.5005
R623 VOUT.n157 VOUT.n105 4.5005
R624 VOUT.n157 VOUT.n102 4.5005
R625 VOUT.n157 VOUT.n106 4.5005
R626 VOUT.n157 VOUT.n101 4.5005
R627 VOUT.n157 VOUT.t94 4.5005
R628 VOUT.n157 VOUT.n100 4.5005
R629 VOUT.n157 VOUT.n107 4.5005
R630 VOUT.n157 VOUT.n156 4.5005
R631 VOUT.n139 VOUT.n103 4.5005
R632 VOUT.n139 VOUT.n105 4.5005
R633 VOUT.n139 VOUT.n102 4.5005
R634 VOUT.n139 VOUT.n106 4.5005
R635 VOUT.n139 VOUT.n101 4.5005
R636 VOUT.n139 VOUT.t94 4.5005
R637 VOUT.n139 VOUT.n100 4.5005
R638 VOUT.n139 VOUT.n107 4.5005
R639 VOUT.n156 VOUT.n139 4.5005
R640 VOUT.n111 VOUT.n103 4.5005
R641 VOUT.n111 VOUT.n105 4.5005
R642 VOUT.n111 VOUT.n102 4.5005
R643 VOUT.n111 VOUT.n106 4.5005
R644 VOUT.n111 VOUT.n101 4.5005
R645 VOUT.n111 VOUT.t94 4.5005
R646 VOUT.n111 VOUT.n100 4.5005
R647 VOUT.n111 VOUT.n107 4.5005
R648 VOUT.n156 VOUT.n111 4.5005
R649 VOUT.n141 VOUT.n103 4.5005
R650 VOUT.n141 VOUT.n105 4.5005
R651 VOUT.n141 VOUT.n102 4.5005
R652 VOUT.n141 VOUT.n106 4.5005
R653 VOUT.n141 VOUT.n101 4.5005
R654 VOUT.n141 VOUT.t94 4.5005
R655 VOUT.n141 VOUT.n100 4.5005
R656 VOUT.n141 VOUT.n107 4.5005
R657 VOUT.n156 VOUT.n141 4.5005
R658 VOUT.n110 VOUT.n103 4.5005
R659 VOUT.n110 VOUT.n105 4.5005
R660 VOUT.n110 VOUT.n102 4.5005
R661 VOUT.n110 VOUT.n106 4.5005
R662 VOUT.n110 VOUT.n101 4.5005
R663 VOUT.n110 VOUT.t94 4.5005
R664 VOUT.n110 VOUT.n100 4.5005
R665 VOUT.n110 VOUT.n107 4.5005
R666 VOUT.n156 VOUT.n110 4.5005
R667 VOUT.n155 VOUT.n103 4.5005
R668 VOUT.n155 VOUT.n105 4.5005
R669 VOUT.n155 VOUT.n102 4.5005
R670 VOUT.n155 VOUT.n106 4.5005
R671 VOUT.n155 VOUT.n101 4.5005
R672 VOUT.n155 VOUT.t94 4.5005
R673 VOUT.n155 VOUT.n100 4.5005
R674 VOUT.n155 VOUT.n107 4.5005
R675 VOUT.n156 VOUT.n155 4.5005
R676 VOUT.n154 VOUT.n39 4.5005
R677 VOUT.n55 VOUT.n39 4.5005
R678 VOUT.n50 VOUT.n34 4.5005
R679 VOUT.n50 VOUT.n36 4.5005
R680 VOUT.n50 VOUT.n33 4.5005
R681 VOUT.n50 VOUT.n37 4.5005
R682 VOUT.n50 VOUT.n32 4.5005
R683 VOUT.n50 VOUT.t95 4.5005
R684 VOUT.n50 VOUT.n31 4.5005
R685 VOUT.n50 VOUT.n38 4.5005
R686 VOUT.n50 VOUT.n39 4.5005
R687 VOUT.n48 VOUT.n34 4.5005
R688 VOUT.n48 VOUT.n36 4.5005
R689 VOUT.n48 VOUT.n33 4.5005
R690 VOUT.n48 VOUT.n37 4.5005
R691 VOUT.n48 VOUT.n32 4.5005
R692 VOUT.n48 VOUT.t95 4.5005
R693 VOUT.n48 VOUT.n31 4.5005
R694 VOUT.n48 VOUT.n38 4.5005
R695 VOUT.n48 VOUT.n39 4.5005
R696 VOUT.n47 VOUT.n34 4.5005
R697 VOUT.n47 VOUT.n36 4.5005
R698 VOUT.n47 VOUT.n33 4.5005
R699 VOUT.n47 VOUT.n37 4.5005
R700 VOUT.n47 VOUT.n32 4.5005
R701 VOUT.n47 VOUT.t95 4.5005
R702 VOUT.n47 VOUT.n31 4.5005
R703 VOUT.n47 VOUT.n38 4.5005
R704 VOUT.n47 VOUT.n39 4.5005
R705 VOUT.n176 VOUT.n34 4.5005
R706 VOUT.n176 VOUT.n36 4.5005
R707 VOUT.n176 VOUT.n33 4.5005
R708 VOUT.n176 VOUT.n37 4.5005
R709 VOUT.n176 VOUT.n32 4.5005
R710 VOUT.n176 VOUT.t95 4.5005
R711 VOUT.n176 VOUT.n31 4.5005
R712 VOUT.n176 VOUT.n38 4.5005
R713 VOUT.n176 VOUT.n39 4.5005
R714 VOUT.n174 VOUT.n34 4.5005
R715 VOUT.n174 VOUT.n36 4.5005
R716 VOUT.n174 VOUT.n33 4.5005
R717 VOUT.n174 VOUT.n37 4.5005
R718 VOUT.n174 VOUT.n32 4.5005
R719 VOUT.n174 VOUT.t95 4.5005
R720 VOUT.n174 VOUT.n31 4.5005
R721 VOUT.n174 VOUT.n38 4.5005
R722 VOUT.n172 VOUT.n34 4.5005
R723 VOUT.n172 VOUT.n36 4.5005
R724 VOUT.n172 VOUT.n33 4.5005
R725 VOUT.n172 VOUT.n37 4.5005
R726 VOUT.n172 VOUT.n32 4.5005
R727 VOUT.n172 VOUT.t95 4.5005
R728 VOUT.n172 VOUT.n31 4.5005
R729 VOUT.n172 VOUT.n38 4.5005
R730 VOUT.n58 VOUT.n34 4.5005
R731 VOUT.n58 VOUT.n36 4.5005
R732 VOUT.n58 VOUT.n33 4.5005
R733 VOUT.n58 VOUT.n37 4.5005
R734 VOUT.n58 VOUT.n32 4.5005
R735 VOUT.n58 VOUT.t95 4.5005
R736 VOUT.n58 VOUT.n31 4.5005
R737 VOUT.n58 VOUT.n38 4.5005
R738 VOUT.n58 VOUT.n39 4.5005
R739 VOUT.n57 VOUT.n34 4.5005
R740 VOUT.n57 VOUT.n36 4.5005
R741 VOUT.n57 VOUT.n33 4.5005
R742 VOUT.n57 VOUT.n37 4.5005
R743 VOUT.n57 VOUT.n32 4.5005
R744 VOUT.n57 VOUT.t95 4.5005
R745 VOUT.n57 VOUT.n31 4.5005
R746 VOUT.n57 VOUT.n38 4.5005
R747 VOUT.n57 VOUT.n39 4.5005
R748 VOUT.n61 VOUT.n34 4.5005
R749 VOUT.n61 VOUT.n36 4.5005
R750 VOUT.n61 VOUT.n33 4.5005
R751 VOUT.n61 VOUT.n37 4.5005
R752 VOUT.n61 VOUT.n32 4.5005
R753 VOUT.n61 VOUT.t95 4.5005
R754 VOUT.n61 VOUT.n31 4.5005
R755 VOUT.n61 VOUT.n38 4.5005
R756 VOUT.n61 VOUT.n39 4.5005
R757 VOUT.n60 VOUT.n34 4.5005
R758 VOUT.n60 VOUT.n36 4.5005
R759 VOUT.n60 VOUT.n33 4.5005
R760 VOUT.n60 VOUT.n37 4.5005
R761 VOUT.n60 VOUT.n32 4.5005
R762 VOUT.n60 VOUT.t95 4.5005
R763 VOUT.n60 VOUT.n31 4.5005
R764 VOUT.n60 VOUT.n38 4.5005
R765 VOUT.n60 VOUT.n39 4.5005
R766 VOUT.n43 VOUT.n34 4.5005
R767 VOUT.n43 VOUT.n36 4.5005
R768 VOUT.n43 VOUT.n33 4.5005
R769 VOUT.n43 VOUT.n37 4.5005
R770 VOUT.n43 VOUT.n32 4.5005
R771 VOUT.n43 VOUT.t95 4.5005
R772 VOUT.n43 VOUT.n31 4.5005
R773 VOUT.n43 VOUT.n38 4.5005
R774 VOUT.n43 VOUT.n39 4.5005
R775 VOUT.n179 VOUT.n34 4.5005
R776 VOUT.n179 VOUT.n36 4.5005
R777 VOUT.n179 VOUT.n33 4.5005
R778 VOUT.n179 VOUT.n37 4.5005
R779 VOUT.n179 VOUT.n32 4.5005
R780 VOUT.n179 VOUT.t95 4.5005
R781 VOUT.n179 VOUT.n31 4.5005
R782 VOUT.n179 VOUT.n38 4.5005
R783 VOUT.n179 VOUT.n39 4.5005
R784 VOUT.n180 VOUT 3.7135
R785 VOUT.n243 VOUT.n242 3.60085
R786 VOUT.n223 VOUT.t0 3.3005
R787 VOUT.n223 VOUT.t3 3.3005
R788 VOUT.n221 VOUT.t22 3.3005
R789 VOUT.n221 VOUT.t19 3.3005
R790 VOUT.n219 VOUT.t6 3.3005
R791 VOUT.n219 VOUT.t27 3.3005
R792 VOUT.n218 VOUT.t15 3.3005
R793 VOUT.n218 VOUT.t18 3.3005
R794 VOUT.n216 VOUT.t23 3.3005
R795 VOUT.n216 VOUT.t14 3.3005
R796 VOUT.n214 VOUT.t89 3.3005
R797 VOUT.n214 VOUT.t5 3.3005
R798 VOUT.n212 VOUT.t1 3.3005
R799 VOUT.n212 VOUT.t21 3.3005
R800 VOUT.n211 VOUT.t20 3.3005
R801 VOUT.n211 VOUT.t11 3.3005
R802 VOUT.n234 VOUT.t9 3.3005
R803 VOUT.n234 VOUT.t8 3.3005
R804 VOUT.n235 VOUT.t7 3.3005
R805 VOUT.n235 VOUT.t10 3.3005
R806 VOUT.n237 VOUT.t4 3.3005
R807 VOUT.n237 VOUT.t25 3.3005
R808 VOUT.n239 VOUT.t12 3.3005
R809 VOUT.n239 VOUT.t26 3.3005
R810 VOUT.n227 VOUT.t2 3.3005
R811 VOUT.n227 VOUT.t90 3.3005
R812 VOUT.n228 VOUT.t16 3.3005
R813 VOUT.n228 VOUT.t91 3.3005
R814 VOUT.n230 VOUT.t13 3.3005
R815 VOUT.n230 VOUT.t17 3.3005
R816 VOUT.n232 VOUT.t24 3.3005
R817 VOUT.n232 VOUT.t88 3.3005
R818 VOUT.n242 VOUT.n226 2.72901
R819 VOUT.n210 VOUT.n29 2.58049
R820 VOUT.n120 VOUT.n118 2.251
R821 VOUT.n120 VOUT.n117 2.251
R822 VOUT.n120 VOUT.n116 2.251
R823 VOUT.n120 VOUT.n115 2.251
R824 VOUT.n89 VOUT.n88 2.251
R825 VOUT.n89 VOUT.n87 2.251
R826 VOUT.n89 VOUT.n86 2.251
R827 VOUT.n89 VOUT.n85 2.251
R828 VOUT.n162 VOUT.n161 2.251
R829 VOUT.n127 VOUT.n125 2.251
R830 VOUT.n127 VOUT.n124 2.251
R831 VOUT.n127 VOUT.n123 2.251
R832 VOUT.n145 VOUT.n127 2.251
R833 VOUT.n133 VOUT.n132 2.251
R834 VOUT.n133 VOUT.n131 2.251
R835 VOUT.n133 VOUT.n130 2.251
R836 VOUT.n133 VOUT.n129 2.251
R837 VOUT.n159 VOUT.n99 2.251
R838 VOUT.n154 VOUT.n152 2.251
R839 VOUT.n154 VOUT.n151 2.251
R840 VOUT.n154 VOUT.n150 2.251
R841 VOUT.n154 VOUT.n149 2.251
R842 VOUT.n55 VOUT.n54 2.251
R843 VOUT.n55 VOUT.n53 2.251
R844 VOUT.n55 VOUT.n52 2.251
R845 VOUT.n55 VOUT.n51 2.251
R846 VOUT.n172 VOUT.n171 2.251
R847 VOUT.n89 VOUT.n69 2.2505
R848 VOUT.n84 VOUT.n69 2.2505
R849 VOUT.n82 VOUT.n69 2.2505
R850 VOUT.n81 VOUT.n69 2.2505
R851 VOUT.n166 VOUT.n69 2.2505
R852 VOUT.n164 VOUT.n69 2.2505
R853 VOUT.n162 VOUT.n69 2.2505
R854 VOUT.n92 VOUT.n69 2.2505
R855 VOUT.n91 VOUT.n69 2.2505
R856 VOUT.n95 VOUT.n69 2.2505
R857 VOUT.n94 VOUT.n69 2.2505
R858 VOUT.n77 VOUT.n69 2.2505
R859 VOUT.n169 VOUT.n69 2.2505
R860 VOUT.n169 VOUT.n168 2.2505
R861 VOUT.n133 VOUT.n104 2.2505
R862 VOUT.n114 VOUT.n104 2.2505
R863 VOUT.n135 VOUT.n104 2.2505
R864 VOUT.n113 VOUT.n104 2.2505
R865 VOUT.n137 VOUT.n104 2.2505
R866 VOUT.n104 VOUT.n98 2.2505
R867 VOUT.n159 VOUT.n104 2.2505
R868 VOUT.n157 VOUT.n104 2.2505
R869 VOUT.n139 VOUT.n104 2.2505
R870 VOUT.n111 VOUT.n104 2.2505
R871 VOUT.n141 VOUT.n104 2.2505
R872 VOUT.n110 VOUT.n104 2.2505
R873 VOUT.n155 VOUT.n104 2.2505
R874 VOUT.n155 VOUT.n108 2.2505
R875 VOUT.n55 VOUT.n35 2.2505
R876 VOUT.n50 VOUT.n35 2.2505
R877 VOUT.n48 VOUT.n35 2.2505
R878 VOUT.n47 VOUT.n35 2.2505
R879 VOUT.n176 VOUT.n35 2.2505
R880 VOUT.n174 VOUT.n35 2.2505
R881 VOUT.n172 VOUT.n35 2.2505
R882 VOUT.n58 VOUT.n35 2.2505
R883 VOUT.n57 VOUT.n35 2.2505
R884 VOUT.n61 VOUT.n35 2.2505
R885 VOUT.n60 VOUT.n35 2.2505
R886 VOUT.n43 VOUT.n35 2.2505
R887 VOUT.n179 VOUT.n35 2.2505
R888 VOUT.n179 VOUT.n178 2.2505
R889 VOUT.n97 VOUT.n90 2.25024
R890 VOUT.n97 VOUT.n83 2.25024
R891 VOUT.n165 VOUT.n97 2.25024
R892 VOUT.n97 VOUT.n93 2.25024
R893 VOUT.n97 VOUT.n96 2.25024
R894 VOUT.n97 VOUT.n64 2.25024
R895 VOUT.n147 VOUT.n144 2.25024
R896 VOUT.n147 VOUT.n143 2.25024
R897 VOUT.n147 VOUT.n142 2.25024
R898 VOUT.n147 VOUT.n109 2.25024
R899 VOUT.n147 VOUT.n146 2.25024
R900 VOUT.n148 VOUT.n147 2.25024
R901 VOUT.n63 VOUT.n56 2.25024
R902 VOUT.n63 VOUT.n49 2.25024
R903 VOUT.n175 VOUT.n63 2.25024
R904 VOUT.n63 VOUT.n59 2.25024
R905 VOUT.n63 VOUT.n62 2.25024
R906 VOUT.n63 VOUT.n30 2.25024
R907 VOUT.n209 VOUT.n199 2.12227
R908 VOUT.n28 VOUT.n18 2.12227
R909 VOUT.n164 VOUT.n74 1.50111
R910 VOUT.n112 VOUT.n98 1.50111
R911 VOUT.n174 VOUT.n40 1.50111
R912 VOUT.n120 VOUT.n119 1.501
R913 VOUT.n127 VOUT.n126 1.501
R914 VOUT.n154 VOUT.n153 1.501
R915 VOUT.n168 VOUT.n79 1.12536
R916 VOUT.n168 VOUT.n80 1.12536
R917 VOUT.n168 VOUT.n167 1.12536
R918 VOUT.n128 VOUT.n108 1.12536
R919 VOUT.n134 VOUT.n108 1.12536
R920 VOUT.n136 VOUT.n108 1.12536
R921 VOUT.n178 VOUT.n45 1.12536
R922 VOUT.n178 VOUT.n46 1.12536
R923 VOUT.n178 VOUT.n177 1.12536
R924 VOUT.n168 VOUT.n75 1.12536
R925 VOUT.n168 VOUT.n76 1.12536
R926 VOUT.n168 VOUT.n78 1.12536
R927 VOUT.n158 VOUT.n108 1.12536
R928 VOUT.n138 VOUT.n108 1.12536
R929 VOUT.n140 VOUT.n108 1.12536
R930 VOUT.n178 VOUT.n41 1.12536
R931 VOUT.n178 VOUT.n42 1.12536
R932 VOUT.n178 VOUT.n44 1.12536
R933 VOUT.n222 VOUT.n220 1.00481
R934 VOUT.n224 VOUT.n222 1.00481
R935 VOUT.n215 VOUT.n213 1.00481
R936 VOUT.n217 VOUT.n215 1.00481
R937 VOUT.n240 VOUT.n238 1.00481
R938 VOUT.n238 VOUT.n236 1.00481
R939 VOUT.n233 VOUT.n231 1.00481
R940 VOUT.n231 VOUT.n229 1.00481
R941 VOUT.n204 VOUT.n202 0.573776
R942 VOUT.n206 VOUT.n204 0.573776
R943 VOUT.n208 VOUT.n206 0.573776
R944 VOUT.n194 VOUT.n192 0.573776
R945 VOUT.n196 VOUT.n194 0.573776
R946 VOUT.n198 VOUT.n196 0.573776
R947 VOUT.n185 VOUT.n183 0.573776
R948 VOUT.n187 VOUT.n185 0.573776
R949 VOUT.n189 VOUT.n187 0.573776
R950 VOUT.n27 VOUT.n25 0.573776
R951 VOUT.n25 VOUT.n23 0.573776
R952 VOUT.n23 VOUT.n21 0.573776
R953 VOUT.n17 VOUT.n15 0.573776
R954 VOUT.n15 VOUT.n13 0.573776
R955 VOUT.n13 VOUT.n11 0.573776
R956 VOUT.n8 VOUT.n6 0.573776
R957 VOUT.n6 VOUT.n4 0.573776
R958 VOUT.n4 VOUT.n2 0.573776
R959 VOUT.n180 VOUT.n179 0.368072
R960 VOUT.n243 VOUT.n180 0.3624
R961 VOUT.n122 VOUT.n121 0.0910737
R962 VOUT.n173 VOUT.n170 0.0723685
R963 VOUT.n127 VOUT.n122 0.0522944
R964 VOUT.n170 VOUT.n169 0.0499135
R965 VOUT.n121 VOUT.n120 0.0499135
R966 VOUT.n155 VOUT.n154 0.0464294
R967 VOUT.n163 VOUT.n160 0.0391444
R968 VOUT.n122 VOUT.t93 0.023435
R969 VOUT.n170 VOUT.t92 0.02262
R970 VOUT.n121 VOUT.t96 0.02262
R971 VOUT VOUT.n243 0.0099
R972 VOUT.n92 VOUT.n75 0.00365111
R973 VOUT.n95 VOUT.n76 0.00365111
R974 VOUT.n78 VOUT.n77 0.00365111
R975 VOUT.n120 VOUT.n79 0.00365111
R976 VOUT.n84 VOUT.n80 0.00365111
R977 VOUT.n167 VOUT.n81 0.00365111
R978 VOUT.n158 VOUT.n157 0.00365111
R979 VOUT.n138 VOUT.n111 0.00365111
R980 VOUT.n140 VOUT.n110 0.00365111
R981 VOUT.n128 VOUT.n127 0.00365111
R982 VOUT.n134 VOUT.n114 0.00365111
R983 VOUT.n136 VOUT.n113 0.00365111
R984 VOUT.n58 VOUT.n41 0.00365111
R985 VOUT.n61 VOUT.n42 0.00365111
R986 VOUT.n44 VOUT.n43 0.00365111
R987 VOUT.n154 VOUT.n45 0.00365111
R988 VOUT.n50 VOUT.n46 0.00365111
R989 VOUT.n177 VOUT.n47 0.00365111
R990 VOUT.n89 VOUT.n79 0.00340054
R991 VOUT.n82 VOUT.n80 0.00340054
R992 VOUT.n167 VOUT.n166 0.00340054
R993 VOUT.n162 VOUT.n75 0.00340054
R994 VOUT.n91 VOUT.n76 0.00340054
R995 VOUT.n94 VOUT.n78 0.00340054
R996 VOUT.n133 VOUT.n128 0.00340054
R997 VOUT.n135 VOUT.n134 0.00340054
R998 VOUT.n137 VOUT.n136 0.00340054
R999 VOUT.n159 VOUT.n158 0.00340054
R1000 VOUT.n139 VOUT.n138 0.00340054
R1001 VOUT.n141 VOUT.n140 0.00340054
R1002 VOUT.n55 VOUT.n45 0.00340054
R1003 VOUT.n48 VOUT.n46 0.00340054
R1004 VOUT.n177 VOUT.n176 0.00340054
R1005 VOUT.n172 VOUT.n41 0.00340054
R1006 VOUT.n57 VOUT.n42 0.00340054
R1007 VOUT.n60 VOUT.n44 0.00340054
R1008 VOUT.n90 VOUT.n84 0.00252698
R1009 VOUT.n83 VOUT.n81 0.00252698
R1010 VOUT.n165 VOUT.n164 0.00252698
R1011 VOUT.n93 VOUT.n91 0.00252698
R1012 VOUT.n96 VOUT.n94 0.00252698
R1013 VOUT.n169 VOUT.n64 0.00252698
R1014 VOUT.n90 VOUT.n89 0.00252698
R1015 VOUT.n83 VOUT.n82 0.00252698
R1016 VOUT.n166 VOUT.n165 0.00252698
R1017 VOUT.n93 VOUT.n92 0.00252698
R1018 VOUT.n96 VOUT.n95 0.00252698
R1019 VOUT.n77 VOUT.n64 0.00252698
R1020 VOUT.n144 VOUT.n114 0.00252698
R1021 VOUT.n143 VOUT.n113 0.00252698
R1022 VOUT.n142 VOUT.n98 0.00252698
R1023 VOUT.n139 VOUT.n109 0.00252698
R1024 VOUT.n146 VOUT.n141 0.00252698
R1025 VOUT.n155 VOUT.n148 0.00252698
R1026 VOUT.n144 VOUT.n133 0.00252698
R1027 VOUT.n143 VOUT.n135 0.00252698
R1028 VOUT.n142 VOUT.n137 0.00252698
R1029 VOUT.n157 VOUT.n109 0.00252698
R1030 VOUT.n146 VOUT.n111 0.00252698
R1031 VOUT.n148 VOUT.n110 0.00252698
R1032 VOUT.n56 VOUT.n50 0.00252698
R1033 VOUT.n49 VOUT.n47 0.00252698
R1034 VOUT.n175 VOUT.n174 0.00252698
R1035 VOUT.n59 VOUT.n57 0.00252698
R1036 VOUT.n62 VOUT.n60 0.00252698
R1037 VOUT.n179 VOUT.n30 0.00252698
R1038 VOUT.n56 VOUT.n55 0.00252698
R1039 VOUT.n49 VOUT.n48 0.00252698
R1040 VOUT.n176 VOUT.n175 0.00252698
R1041 VOUT.n59 VOUT.n58 0.00252698
R1042 VOUT.n62 VOUT.n61 0.00252698
R1043 VOUT.n43 VOUT.n30 0.00252698
R1044 VOUT.n164 VOUT.n163 0.0020275
R1045 VOUT.n163 VOUT.n162 0.0020275
R1046 VOUT.n160 VOUT.n98 0.0020275
R1047 VOUT.n160 VOUT.n159 0.0020275
R1048 VOUT.n174 VOUT.n173 0.0020275
R1049 VOUT.n173 VOUT.n172 0.0020275
R1050 VOUT.n74 VOUT.n73 0.00166668
R1051 VOUT.n156 VOUT.n112 0.00166668
R1052 VOUT.n40 VOUT.n39 0.00166668
R1053 VOUT.n178 VOUT.n40 0.00133328
R1054 VOUT.n112 VOUT.n108 0.00133328
R1055 VOUT.n168 VOUT.n74 0.00133328
R1056 VOUT.n171 VOUT.n63 0.001
R1057 VOUT.n149 VOUT.n63 0.001
R1058 VOUT.n51 VOUT.n31 0.001
R1059 VOUT.n150 VOUT.n31 0.001
R1060 VOUT.n52 VOUT.n32 0.001
R1061 VOUT.n151 VOUT.n32 0.001
R1062 VOUT.n53 VOUT.n33 0.001
R1063 VOUT.n152 VOUT.n33 0.001
R1064 VOUT.n54 VOUT.n34 0.001
R1065 VOUT.n153 VOUT.n34 0.001
R1066 VOUT.n147 VOUT.n99 0.001
R1067 VOUT.n147 VOUT.n145 0.001
R1068 VOUT.n129 VOUT.n100 0.001
R1069 VOUT.n123 VOUT.n100 0.001
R1070 VOUT.n130 VOUT.n101 0.001
R1071 VOUT.n124 VOUT.n101 0.001
R1072 VOUT.n131 VOUT.n102 0.001
R1073 VOUT.n125 VOUT.n102 0.001
R1074 VOUT.n132 VOUT.n103 0.001
R1075 VOUT.n126 VOUT.n103 0.001
R1076 VOUT.n161 VOUT.n97 0.001
R1077 VOUT.n115 VOUT.n97 0.001
R1078 VOUT.n85 VOUT.n65 0.001
R1079 VOUT.n116 VOUT.n65 0.001
R1080 VOUT.n86 VOUT.n66 0.001
R1081 VOUT.n117 VOUT.n66 0.001
R1082 VOUT.n87 VOUT.n67 0.001
R1083 VOUT.n118 VOUT.n67 0.001
R1084 VOUT.n88 VOUT.n68 0.001
R1085 VOUT.n119 VOUT.n68 0.001
R1086 VOUT.n119 VOUT.n69 0.001
R1087 VOUT.n118 VOUT.n70 0.001
R1088 VOUT.n117 VOUT.n71 0.001
R1089 VOUT.n116 VOUT.t97 0.001
R1090 VOUT.n115 VOUT.n72 0.001
R1091 VOUT.n88 VOUT.n70 0.001
R1092 VOUT.n87 VOUT.n71 0.001
R1093 VOUT.n86 VOUT.t97 0.001
R1094 VOUT.n85 VOUT.n72 0.001
R1095 VOUT.n161 VOUT.n73 0.001
R1096 VOUT.n126 VOUT.n104 0.001
R1097 VOUT.n125 VOUT.n105 0.001
R1098 VOUT.n124 VOUT.n106 0.001
R1099 VOUT.n123 VOUT.t94 0.001
R1100 VOUT.n145 VOUT.n107 0.001
R1101 VOUT.n132 VOUT.n105 0.001
R1102 VOUT.n131 VOUT.n106 0.001
R1103 VOUT.n130 VOUT.t94 0.001
R1104 VOUT.n129 VOUT.n107 0.001
R1105 VOUT.n156 VOUT.n99 0.001
R1106 VOUT.n153 VOUT.n35 0.001
R1107 VOUT.n152 VOUT.n36 0.001
R1108 VOUT.n151 VOUT.n37 0.001
R1109 VOUT.n150 VOUT.t95 0.001
R1110 VOUT.n149 VOUT.n38 0.001
R1111 VOUT.n54 VOUT.n36 0.001
R1112 VOUT.n53 VOUT.n37 0.001
R1113 VOUT.n52 VOUT.t95 0.001
R1114 VOUT.n51 VOUT.n38 0.001
R1115 VOUT.n171 VOUT.n39 0.001
R1116 VDD.n2697 VDD.n99 452.195
R1117 VDD.n2590 VDD.n97 452.195
R1118 VDD.n303 VDD.n268 452.195
R1119 VDD.n2483 VDD.n270 452.195
R1120 VDD.n1398 VDD.n716 452.195
R1121 VDD.n1401 VDD.n1400 452.195
R1122 VDD.n887 VDD.n853 452.195
R1123 VDD.n1064 VDD.n855 452.195
R1124 VDD.n969 VDD.t77 371.625
R1125 VDD.n1002 VDD.t90 371.625
R1126 VDD.n1035 VDD.t39 371.625
R1127 VDD.n705 VDD.t43 371.625
R1128 VDD.n1277 VDD.t55 371.625
R1129 VDD.n1242 VDD.t99 371.625
R1130 VDD.n199 VDD.t62 371.625
R1131 VDD.n166 VDD.t74 371.625
R1132 VDD.n131 VDD.t106 371.625
R1133 VDD.n341 VDD.t112 371.625
R1134 VDD.n2450 VDD.t83 371.625
R1135 VDD.n2367 VDD.t70 371.625
R1136 VDD.n689 VDD.t96 347.526
R1137 VDD.n540 VDD.t109 347.526
R1138 VDD.n682 VDD.t66 347.526
R1139 VDD.n550 VDD.t86 347.526
R1140 VDD.n408 VDD.t102 347.526
R1141 VDD.n1887 VDD.t58 347.526
R1142 VDD.n391 VDD.t51 347.526
R1143 VDD.n1893 VDD.t80 347.526
R1144 VDD.n364 VDD.t93 347.526
R1145 VDD.n650 VDD.t47 347.526
R1146 VDD.n2127 VDD.n509 294.147
R1147 VDD.n2331 VDD.n374 294.147
R1148 VDD.n2283 VDD.n371 294.147
R1149 VDD.n1954 VDD.n1871 294.147
R1150 VDD.n1810 VDD.n548 294.147
R1151 VDD.n1759 VDD.n1758 294.147
R1152 VDD.n1584 VDD.n667 294.147
R1153 VDD.n1635 VDD.n669 294.147
R1154 VDD.n2262 VDD.n372 294.147
R1155 VDD.n2334 VDD.n2333 294.147
R1156 VDD.n2073 VDD.n1872 294.147
R1157 VDD.n2125 VDD.n1874 294.147
R1158 VDD.n1868 VDD.n537 294.147
R1159 VDD.n1817 VDD.n536 294.147
R1160 VDD.n1467 VDD.n668 294.147
R1161 VDD.n1637 VDD.n665 294.147
R1162 VDD.n689 VDD.t98 293.986
R1163 VDD.n540 VDD.t110 293.986
R1164 VDD.n682 VDD.t69 293.986
R1165 VDD.n550 VDD.t88 293.986
R1166 VDD.n408 VDD.t104 293.986
R1167 VDD.n408 VDD.t105 293.986
R1168 VDD.n1887 VDD.t61 293.986
R1169 VDD.n391 VDD.t53 293.986
R1170 VDD.n1893 VDD.t82 293.986
R1171 VDD.n364 VDD.t94 293.986
R1172 VDD.n650 VDD.t49 293.986
R1173 VDD.n650 VDD.t50 293.986
R1174 VDD.n690 VDD.t97 268.192
R1175 VDD.n541 VDD.t111 268.192
R1176 VDD.n683 VDD.t68 268.192
R1177 VDD.n551 VDD.t89 268.192
R1178 VDD.n1888 VDD.t60 268.192
R1179 VDD.n392 VDD.t54 268.192
R1180 VDD.n1894 VDD.t81 268.192
R1181 VDD.n365 VDD.t95 268.192
R1182 VDD.n2264 VDD.n372 185
R1183 VDD.n2332 VDD.n372 185
R1184 VDD.n2266 VDD.n2265 185
R1185 VDD.n2265 VDD.n370 185
R1186 VDD.n2267 VDD.n399 185
R1187 VDD.n2277 VDD.n399 185
R1188 VDD.n2268 VDD.n407 185
R1189 VDD.n407 VDD.n397 185
R1190 VDD.n2270 VDD.n2269 185
R1191 VDD.n2271 VDD.n2270 185
R1192 VDD.n2232 VDD.n406 185
R1193 VDD.n406 VDD.n403 185
R1194 VDD.n2230 VDD.n2229 185
R1195 VDD.n2229 VDD.n2228 185
R1196 VDD.n410 VDD.n409 185
R1197 VDD.n411 VDD.n410 185
R1198 VDD.n2221 VDD.n2220 185
R1199 VDD.n2222 VDD.n2221 185
R1200 VDD.n2219 VDD.n420 185
R1201 VDD.n420 VDD.n417 185
R1202 VDD.n2218 VDD.n2217 185
R1203 VDD.n2217 VDD.n2216 185
R1204 VDD.n422 VDD.n421 185
R1205 VDD.n430 VDD.n422 185
R1206 VDD.n2209 VDD.n2208 185
R1207 VDD.n2210 VDD.n2209 185
R1208 VDD.n2207 VDD.n431 185
R1209 VDD.n436 VDD.n431 185
R1210 VDD.n2206 VDD.n2205 185
R1211 VDD.n2205 VDD.n2204 185
R1212 VDD.n433 VDD.n432 185
R1213 VDD.n442 VDD.n433 185
R1214 VDD.n2197 VDD.n2196 185
R1215 VDD.n2198 VDD.n2197 185
R1216 VDD.n2195 VDD.n443 185
R1217 VDD.n448 VDD.n443 185
R1218 VDD.n2194 VDD.n2193 185
R1219 VDD.n2193 VDD.n2192 185
R1220 VDD.n445 VDD.n444 185
R1221 VDD.n454 VDD.n445 185
R1222 VDD.n2185 VDD.n2184 185
R1223 VDD.n2186 VDD.n2185 185
R1224 VDD.n2183 VDD.n455 185
R1225 VDD.n2038 VDD.n455 185
R1226 VDD.n2182 VDD.n2181 185
R1227 VDD.n2181 VDD.n2180 185
R1228 VDD.n457 VDD.n456 185
R1229 VDD.n458 VDD.n457 185
R1230 VDD.n2173 VDD.n2172 185
R1231 VDD.n2174 VDD.n2173 185
R1232 VDD.n2171 VDD.n466 185
R1233 VDD.n2047 VDD.n466 185
R1234 VDD.n2170 VDD.n2169 185
R1235 VDD.n2169 VDD.n2168 185
R1236 VDD.n468 VDD.n467 185
R1237 VDD.n469 VDD.n468 185
R1238 VDD.n2161 VDD.n2160 185
R1239 VDD.n2162 VDD.n2161 185
R1240 VDD.n2159 VDD.n478 185
R1241 VDD.n478 VDD.n475 185
R1242 VDD.n2158 VDD.n2157 185
R1243 VDD.n2157 VDD.n2156 185
R1244 VDD.n480 VDD.n479 185
R1245 VDD.n489 VDD.n480 185
R1246 VDD.n2149 VDD.n2148 185
R1247 VDD.n2150 VDD.n2149 185
R1248 VDD.n2147 VDD.n490 185
R1249 VDD.n490 VDD.n486 185
R1250 VDD.n2146 VDD.n2145 185
R1251 VDD.n2145 VDD.n2144 185
R1252 VDD.n492 VDD.n491 185
R1253 VDD.n500 VDD.n492 185
R1254 VDD.n2137 VDD.n2136 185
R1255 VDD.n2138 VDD.n2137 185
R1256 VDD.n2135 VDD.n501 185
R1257 VDD.n506 VDD.n501 185
R1258 VDD.n2134 VDD.n2133 185
R1259 VDD.n2133 VDD.n2132 185
R1260 VDD.n503 VDD.n502 185
R1261 VDD.n1873 VDD.n503 185
R1262 VDD.n2125 VDD.n2124 185
R1263 VDD.n2126 VDD.n2125 185
R1264 VDD.n2123 VDD.n1874 185
R1265 VDD.n2122 VDD.n2121 185
R1266 VDD.n2119 VDD.n1875 185
R1267 VDD.n2117 VDD.n2116 185
R1268 VDD.n2115 VDD.n1876 185
R1269 VDD.n2114 VDD.n2113 185
R1270 VDD.n2111 VDD.n1877 185
R1271 VDD.n2109 VDD.n2108 185
R1272 VDD.n2107 VDD.n1878 185
R1273 VDD.n2106 VDD.n2105 185
R1274 VDD.n2103 VDD.n1879 185
R1275 VDD.n2101 VDD.n2100 185
R1276 VDD.n2099 VDD.n1880 185
R1277 VDD.n2098 VDD.n2097 185
R1278 VDD.n2095 VDD.n1881 185
R1279 VDD.n2093 VDD.n2092 185
R1280 VDD.n2091 VDD.n1882 185
R1281 VDD.n2090 VDD.n2089 185
R1282 VDD.n2087 VDD.n1883 185
R1283 VDD.n2085 VDD.n2084 185
R1284 VDD.n2083 VDD.n1884 185
R1285 VDD.n2082 VDD.n2081 185
R1286 VDD.n2079 VDD.n1885 185
R1287 VDD.n2077 VDD.n2076 185
R1288 VDD.n2075 VDD.n1886 185
R1289 VDD.n2074 VDD.n2073 185
R1290 VDD.n2335 VDD.n2334 185
R1291 VDD.n2336 VDD.n363 185
R1292 VDD.n2338 VDD.n2337 185
R1293 VDD.n2340 VDD.n361 185
R1294 VDD.n2342 VDD.n2341 185
R1295 VDD.n2343 VDD.n360 185
R1296 VDD.n2345 VDD.n2344 185
R1297 VDD.n2347 VDD.n358 185
R1298 VDD.n2349 VDD.n2348 185
R1299 VDD.n2350 VDD.n357 185
R1300 VDD.n2352 VDD.n2351 185
R1301 VDD.n2354 VDD.n355 185
R1302 VDD.n2356 VDD.n2355 185
R1303 VDD.n2241 VDD.n354 185
R1304 VDD.n2243 VDD.n2242 185
R1305 VDD.n2245 VDD.n2239 185
R1306 VDD.n2247 VDD.n2246 185
R1307 VDD.n2248 VDD.n2238 185
R1308 VDD.n2250 VDD.n2249 185
R1309 VDD.n2252 VDD.n2236 185
R1310 VDD.n2254 VDD.n2253 185
R1311 VDD.n2255 VDD.n2235 185
R1312 VDD.n2257 VDD.n2256 185
R1313 VDD.n2259 VDD.n2234 185
R1314 VDD.n2260 VDD.n2233 185
R1315 VDD.n2263 VDD.n2262 185
R1316 VDD.n2333 VDD.n367 185
R1317 VDD.n2333 VDD.n2332 185
R1318 VDD.n2007 VDD.n369 185
R1319 VDD.n370 VDD.n369 185
R1320 VDD.n2008 VDD.n398 185
R1321 VDD.n2277 VDD.n398 185
R1322 VDD.n2010 VDD.n2009 185
R1323 VDD.n2009 VDD.n397 185
R1324 VDD.n2011 VDD.n405 185
R1325 VDD.n2271 VDD.n405 185
R1326 VDD.n2013 VDD.n2012 185
R1327 VDD.n2012 VDD.n403 185
R1328 VDD.n2014 VDD.n413 185
R1329 VDD.n2228 VDD.n413 185
R1330 VDD.n2016 VDD.n2015 185
R1331 VDD.n2015 VDD.n411 185
R1332 VDD.n2017 VDD.n419 185
R1333 VDD.n2222 VDD.n419 185
R1334 VDD.n2019 VDD.n2018 185
R1335 VDD.n2018 VDD.n417 185
R1336 VDD.n2020 VDD.n424 185
R1337 VDD.n2216 VDD.n424 185
R1338 VDD.n2022 VDD.n2021 185
R1339 VDD.n2021 VDD.n430 185
R1340 VDD.n2023 VDD.n429 185
R1341 VDD.n2210 VDD.n429 185
R1342 VDD.n2025 VDD.n2024 185
R1343 VDD.n2024 VDD.n436 185
R1344 VDD.n2026 VDD.n435 185
R1345 VDD.n2204 VDD.n435 185
R1346 VDD.n2028 VDD.n2027 185
R1347 VDD.n2027 VDD.n442 185
R1348 VDD.n2029 VDD.n441 185
R1349 VDD.n2198 VDD.n441 185
R1350 VDD.n2031 VDD.n2030 185
R1351 VDD.n2030 VDD.n448 185
R1352 VDD.n2032 VDD.n447 185
R1353 VDD.n2192 VDD.n447 185
R1354 VDD.n2034 VDD.n2033 185
R1355 VDD.n2033 VDD.n454 185
R1356 VDD.n2035 VDD.n453 185
R1357 VDD.n2186 VDD.n453 185
R1358 VDD.n2037 VDD.n2036 185
R1359 VDD.n2038 VDD.n2037 185
R1360 VDD.n2006 VDD.n460 185
R1361 VDD.n2180 VDD.n460 185
R1362 VDD.n2005 VDD.n2004 185
R1363 VDD.n2004 VDD.n458 185
R1364 VDD.n1890 VDD.n465 185
R1365 VDD.n2174 VDD.n465 185
R1366 VDD.n2049 VDD.n2048 185
R1367 VDD.n2048 VDD.n2047 185
R1368 VDD.n2050 VDD.n471 185
R1369 VDD.n2168 VDD.n471 185
R1370 VDD.n2052 VDD.n2051 185
R1371 VDD.n2051 VDD.n469 185
R1372 VDD.n2053 VDD.n477 185
R1373 VDD.n2162 VDD.n477 185
R1374 VDD.n2055 VDD.n2054 185
R1375 VDD.n2054 VDD.n475 185
R1376 VDD.n2056 VDD.n482 185
R1377 VDD.n2156 VDD.n482 185
R1378 VDD.n2058 VDD.n2057 185
R1379 VDD.n2057 VDD.n489 185
R1380 VDD.n2059 VDD.n488 185
R1381 VDD.n2150 VDD.n488 185
R1382 VDD.n2061 VDD.n2060 185
R1383 VDD.n2060 VDD.n486 185
R1384 VDD.n2062 VDD.n494 185
R1385 VDD.n2144 VDD.n494 185
R1386 VDD.n2064 VDD.n2063 185
R1387 VDD.n2063 VDD.n500 185
R1388 VDD.n2065 VDD.n499 185
R1389 VDD.n2138 VDD.n499 185
R1390 VDD.n2067 VDD.n2066 185
R1391 VDD.n2066 VDD.n506 185
R1392 VDD.n2068 VDD.n505 185
R1393 VDD.n2132 VDD.n505 185
R1394 VDD.n2070 VDD.n2069 185
R1395 VDD.n2069 VDD.n1873 185
R1396 VDD.n2071 VDD.n1872 185
R1397 VDD.n2126 VDD.n1872 185
R1398 VDD.n1398 VDD.n1397 185
R1399 VDD.n1399 VDD.n1398 185
R1400 VDD.n717 VDD.n715 185
R1401 VDD.n715 VDD.n712 185
R1402 VDD.n1211 VDD.n1210 185
R1403 VDD.n1210 VDD.n1209 185
R1404 VDD.n720 VDD.n719 185
R1405 VDD.n721 VDD.n720 185
R1406 VDD.n1199 VDD.n1198 185
R1407 VDD.n1200 VDD.n1199 185
R1408 VDD.n730 VDD.n729 185
R1409 VDD.n729 VDD.n728 185
R1410 VDD.n1194 VDD.n1193 185
R1411 VDD.n1193 VDD.n1192 185
R1412 VDD.n733 VDD.n732 185
R1413 VDD.n740 VDD.n733 185
R1414 VDD.n1183 VDD.n1182 185
R1415 VDD.n1184 VDD.n1183 185
R1416 VDD.n742 VDD.n741 185
R1417 VDD.n741 VDD.n739 185
R1418 VDD.n1178 VDD.n1177 185
R1419 VDD.n1177 VDD.n1176 185
R1420 VDD.n745 VDD.n744 185
R1421 VDD.n746 VDD.n745 185
R1422 VDD.n1167 VDD.n1166 185
R1423 VDD.n1168 VDD.n1167 185
R1424 VDD.n754 VDD.n753 185
R1425 VDD.n753 VDD.n752 185
R1426 VDD.n1162 VDD.n1161 185
R1427 VDD.n1161 VDD.n1160 185
R1428 VDD.n757 VDD.n756 185
R1429 VDD.n764 VDD.n757 185
R1430 VDD.n1151 VDD.n1150 185
R1431 VDD.n1152 VDD.n1151 185
R1432 VDD.n766 VDD.n765 185
R1433 VDD.n765 VDD.n763 185
R1434 VDD.n1146 VDD.n1145 185
R1435 VDD.n1145 VDD.n1144 185
R1436 VDD.n799 VDD.n798 185
R1437 VDD.n800 VDD.n799 185
R1438 VDD.n1135 VDD.n1134 185
R1439 VDD.n1136 VDD.n1135 185
R1440 VDD.n808 VDD.n807 185
R1441 VDD.n807 VDD.n806 185
R1442 VDD.n1129 VDD.n1128 185
R1443 VDD.n1128 VDD.n1127 185
R1444 VDD.n811 VDD.n810 185
R1445 VDD.n818 VDD.n811 185
R1446 VDD.n1118 VDD.n1117 185
R1447 VDD.n1119 VDD.n1118 185
R1448 VDD.n820 VDD.n819 185
R1449 VDD.n819 VDD.n817 185
R1450 VDD.n1113 VDD.n1112 185
R1451 VDD.n1112 VDD.n1111 185
R1452 VDD.n823 VDD.n822 185
R1453 VDD.n824 VDD.n823 185
R1454 VDD.n1102 VDD.n1101 185
R1455 VDD.n1103 VDD.n1102 185
R1456 VDD.n832 VDD.n831 185
R1457 VDD.n831 VDD.n830 185
R1458 VDD.n1097 VDD.n1096 185
R1459 VDD.n1096 VDD.n1095 185
R1460 VDD.n835 VDD.n834 185
R1461 VDD.n842 VDD.n835 185
R1462 VDD.n1086 VDD.n1085 185
R1463 VDD.n1087 VDD.n1086 185
R1464 VDD.n844 VDD.n843 185
R1465 VDD.n843 VDD.n841 185
R1466 VDD.n1081 VDD.n1080 185
R1467 VDD.n1080 VDD.n1079 185
R1468 VDD.n847 VDD.n846 185
R1469 VDD.n848 VDD.n847 185
R1470 VDD.n1070 VDD.n1069 185
R1471 VDD.n1071 VDD.n1070 185
R1472 VDD.n856 VDD.n855 185
R1473 VDD.n855 VDD.n854 185
R1474 VDD.n1065 VDD.n1064 185
R1475 VDD.n859 VDD.n858 185
R1476 VDD.n1061 VDD.n1060 185
R1477 VDD.n1062 VDD.n1061 185
R1478 VDD.n889 VDD.n888 185
R1479 VDD.n1056 VDD.n891 185
R1480 VDD.n1055 VDD.n892 185
R1481 VDD.n1054 VDD.n893 185
R1482 VDD.n895 VDD.n894 185
R1483 VDD.n1050 VDD.n897 185
R1484 VDD.n1049 VDD.n898 185
R1485 VDD.n1048 VDD.n899 185
R1486 VDD.n901 VDD.n900 185
R1487 VDD.n1044 VDD.n903 185
R1488 VDD.n1043 VDD.n904 185
R1489 VDD.n1042 VDD.n905 185
R1490 VDD.n907 VDD.n906 185
R1491 VDD.n1038 VDD.n909 185
R1492 VDD.n1037 VDD.n1034 185
R1493 VDD.n1033 VDD.n910 185
R1494 VDD.n912 VDD.n911 185
R1495 VDD.n1029 VDD.n914 185
R1496 VDD.n1028 VDD.n915 185
R1497 VDD.n1027 VDD.n916 185
R1498 VDD.n918 VDD.n917 185
R1499 VDD.n1023 VDD.n920 185
R1500 VDD.n1022 VDD.n921 185
R1501 VDD.n1021 VDD.n922 185
R1502 VDD.n924 VDD.n923 185
R1503 VDD.n1017 VDD.n926 185
R1504 VDD.n1016 VDD.n927 185
R1505 VDD.n1015 VDD.n928 185
R1506 VDD.n930 VDD.n929 185
R1507 VDD.n1011 VDD.n932 185
R1508 VDD.n1010 VDD.n933 185
R1509 VDD.n1009 VDD.n934 185
R1510 VDD.n936 VDD.n935 185
R1511 VDD.n1005 VDD.n938 185
R1512 VDD.n1004 VDD.n1001 185
R1513 VDD.n1000 VDD.n939 185
R1514 VDD.n941 VDD.n940 185
R1515 VDD.n996 VDD.n943 185
R1516 VDD.n995 VDD.n944 185
R1517 VDD.n994 VDD.n945 185
R1518 VDD.n947 VDD.n946 185
R1519 VDD.n990 VDD.n949 185
R1520 VDD.n989 VDD.n950 185
R1521 VDD.n988 VDD.n951 185
R1522 VDD.n953 VDD.n952 185
R1523 VDD.n984 VDD.n955 185
R1524 VDD.n983 VDD.n956 185
R1525 VDD.n982 VDD.n957 185
R1526 VDD.n959 VDD.n958 185
R1527 VDD.n978 VDD.n961 185
R1528 VDD.n977 VDD.n962 185
R1529 VDD.n976 VDD.n963 185
R1530 VDD.n965 VDD.n964 185
R1531 VDD.n972 VDD.n967 185
R1532 VDD.n968 VDD.n887 185
R1533 VDD.n1062 VDD.n887 185
R1534 VDD.n1402 VDD.n1401 185
R1535 VDD.n708 VDD.n703 185
R1536 VDD.n1406 VDD.n702 185
R1537 VDD.n1407 VDD.n701 185
R1538 VDD.n1408 VDD.n700 185
R1539 VDD.n1298 VDD.n699 185
R1540 VDD.n1300 VDD.n1299 185
R1541 VDD.n1302 VDD.n1296 185
R1542 VDD.n1304 VDD.n1303 185
R1543 VDD.n1306 VDD.n1294 185
R1544 VDD.n1308 VDD.n1307 185
R1545 VDD.n1309 VDD.n1289 185
R1546 VDD.n1311 VDD.n1310 185
R1547 VDD.n1313 VDD.n1287 185
R1548 VDD.n1315 VDD.n1314 185
R1549 VDD.n1316 VDD.n1283 185
R1550 VDD.n1318 VDD.n1317 185
R1551 VDD.n1320 VDD.n1281 185
R1552 VDD.n1322 VDD.n1321 185
R1553 VDD.n1276 VDD.n1275 185
R1554 VDD.n1327 VDD.n1326 185
R1555 VDD.n1329 VDD.n1273 185
R1556 VDD.n1331 VDD.n1330 185
R1557 VDD.n1332 VDD.n1268 185
R1558 VDD.n1334 VDD.n1333 185
R1559 VDD.n1336 VDD.n1266 185
R1560 VDD.n1338 VDD.n1337 185
R1561 VDD.n1339 VDD.n1261 185
R1562 VDD.n1341 VDD.n1340 185
R1563 VDD.n1343 VDD.n1259 185
R1564 VDD.n1345 VDD.n1344 185
R1565 VDD.n1346 VDD.n1254 185
R1566 VDD.n1348 VDD.n1347 185
R1567 VDD.n1350 VDD.n1252 185
R1568 VDD.n1352 VDD.n1351 185
R1569 VDD.n1353 VDD.n1248 185
R1570 VDD.n1355 VDD.n1354 185
R1571 VDD.n1357 VDD.n1246 185
R1572 VDD.n1359 VDD.n1358 185
R1573 VDD.n1241 VDD.n1240 185
R1574 VDD.n1364 VDD.n1363 185
R1575 VDD.n1366 VDD.n1238 185
R1576 VDD.n1368 VDD.n1367 185
R1577 VDD.n1369 VDD.n1233 185
R1578 VDD.n1371 VDD.n1370 185
R1579 VDD.n1373 VDD.n1231 185
R1580 VDD.n1375 VDD.n1374 185
R1581 VDD.n1376 VDD.n1228 185
R1582 VDD.n1378 VDD.n1377 185
R1583 VDD.n1380 VDD.n1225 185
R1584 VDD.n1382 VDD.n1381 185
R1585 VDD.n1226 VDD.n1223 185
R1586 VDD.n1386 VDD.n1222 185
R1587 VDD.n1387 VDD.n1217 185
R1588 VDD.n1389 VDD.n1388 185
R1589 VDD.n1391 VDD.n1215 185
R1590 VDD.n1393 VDD.n1392 185
R1591 VDD.n1394 VDD.n716 185
R1592 VDD.n1400 VDD.n711 185
R1593 VDD.n1400 VDD.n1399 185
R1594 VDD.n724 VDD.n710 185
R1595 VDD.n712 VDD.n710 185
R1596 VDD.n1208 VDD.n1207 185
R1597 VDD.n1209 VDD.n1208 185
R1598 VDD.n723 VDD.n722 185
R1599 VDD.n722 VDD.n721 185
R1600 VDD.n1202 VDD.n1201 185
R1601 VDD.n1201 VDD.n1200 185
R1602 VDD.n727 VDD.n726 185
R1603 VDD.n728 VDD.n727 185
R1604 VDD.n1191 VDD.n1190 185
R1605 VDD.n1192 VDD.n1191 185
R1606 VDD.n735 VDD.n734 185
R1607 VDD.n740 VDD.n734 185
R1608 VDD.n1186 VDD.n1185 185
R1609 VDD.n1185 VDD.n1184 185
R1610 VDD.n738 VDD.n737 185
R1611 VDD.n739 VDD.n738 185
R1612 VDD.n1175 VDD.n1174 185
R1613 VDD.n1176 VDD.n1175 185
R1614 VDD.n748 VDD.n747 185
R1615 VDD.n747 VDD.n746 185
R1616 VDD.n1170 VDD.n1169 185
R1617 VDD.n1169 VDD.n1168 185
R1618 VDD.n751 VDD.n750 185
R1619 VDD.n752 VDD.n751 185
R1620 VDD.n1159 VDD.n1158 185
R1621 VDD.n1160 VDD.n1159 185
R1622 VDD.n759 VDD.n758 185
R1623 VDD.n764 VDD.n758 185
R1624 VDD.n1154 VDD.n1153 185
R1625 VDD.n1153 VDD.n1152 185
R1626 VDD.n762 VDD.n761 185
R1627 VDD.n763 VDD.n762 185
R1628 VDD.n1143 VDD.n1142 185
R1629 VDD.n1144 VDD.n1143 185
R1630 VDD.n802 VDD.n801 185
R1631 VDD.n801 VDD.n800 185
R1632 VDD.n1138 VDD.n1137 185
R1633 VDD.n1137 VDD.n1136 185
R1634 VDD.n805 VDD.n804 185
R1635 VDD.n806 VDD.n805 185
R1636 VDD.n1126 VDD.n1125 185
R1637 VDD.n1127 VDD.n1126 185
R1638 VDD.n813 VDD.n812 185
R1639 VDD.n818 VDD.n812 185
R1640 VDD.n1121 VDD.n1120 185
R1641 VDD.n1120 VDD.n1119 185
R1642 VDD.n816 VDD.n815 185
R1643 VDD.n817 VDD.n816 185
R1644 VDD.n1110 VDD.n1109 185
R1645 VDD.n1111 VDD.n1110 185
R1646 VDD.n826 VDD.n825 185
R1647 VDD.n825 VDD.n824 185
R1648 VDD.n1105 VDD.n1104 185
R1649 VDD.n1104 VDD.n1103 185
R1650 VDD.n829 VDD.n828 185
R1651 VDD.n830 VDD.n829 185
R1652 VDD.n1094 VDD.n1093 185
R1653 VDD.n1095 VDD.n1094 185
R1654 VDD.n837 VDD.n836 185
R1655 VDD.n842 VDD.n836 185
R1656 VDD.n1089 VDD.n1088 185
R1657 VDD.n1088 VDD.n1087 185
R1658 VDD.n840 VDD.n839 185
R1659 VDD.n841 VDD.n840 185
R1660 VDD.n1078 VDD.n1077 185
R1661 VDD.n1079 VDD.n1078 185
R1662 VDD.n850 VDD.n849 185
R1663 VDD.n849 VDD.n848 185
R1664 VDD.n1073 VDD.n1072 185
R1665 VDD.n1072 VDD.n1071 185
R1666 VDD.n853 VDD.n852 185
R1667 VDD.n854 VDD.n853 185
R1668 VDD.n1812 VDD.n548 185
R1669 VDD.n548 VDD.n510 185
R1670 VDD.n1814 VDD.n1813 185
R1671 VDD.n1815 VDD.n1814 185
R1672 VDD.n549 VDD.n547 185
R1673 VDD.n1753 VDD.n547 185
R1674 VDD.n1743 VDD.n562 185
R1675 VDD.n562 VDD.n554 185
R1676 VDD.n1745 VDD.n1744 185
R1677 VDD.n1746 VDD.n1745 185
R1678 VDD.n1742 VDD.n561 185
R1679 VDD.n561 VDD.n558 185
R1680 VDD.n1741 VDD.n1740 185
R1681 VDD.n1740 VDD.n1739 185
R1682 VDD.n564 VDD.n563 185
R1683 VDD.n565 VDD.n564 185
R1684 VDD.n1732 VDD.n1731 185
R1685 VDD.n1733 VDD.n1732 185
R1686 VDD.n1730 VDD.n574 185
R1687 VDD.n574 VDD.n571 185
R1688 VDD.n1729 VDD.n1728 185
R1689 VDD.n1728 VDD.n1727 185
R1690 VDD.n576 VDD.n575 185
R1691 VDD.n585 VDD.n576 185
R1692 VDD.n1720 VDD.n1719 185
R1693 VDD.n1721 VDD.n1720 185
R1694 VDD.n1718 VDD.n586 185
R1695 VDD.n586 VDD.n582 185
R1696 VDD.n1717 VDD.n1716 185
R1697 VDD.n1716 VDD.n1715 185
R1698 VDD.n588 VDD.n587 185
R1699 VDD.n1540 VDD.n588 185
R1700 VDD.n1708 VDD.n1707 185
R1701 VDD.n1709 VDD.n1708 185
R1702 VDD.n1706 VDD.n597 185
R1703 VDD.n597 VDD.n594 185
R1704 VDD.n1705 VDD.n1704 185
R1705 VDD.n1704 VDD.n1703 185
R1706 VDD.n599 VDD.n598 185
R1707 VDD.n1549 VDD.n599 185
R1708 VDD.n1696 VDD.n1695 185
R1709 VDD.n1697 VDD.n1696 185
R1710 VDD.n1694 VDD.n608 185
R1711 VDD.n608 VDD.n605 185
R1712 VDD.n1693 VDD.n1692 185
R1713 VDD.n1692 VDD.n1691 185
R1714 VDD.n610 VDD.n609 185
R1715 VDD.n611 VDD.n610 185
R1716 VDD.n1684 VDD.n1683 185
R1717 VDD.n1685 VDD.n1684 185
R1718 VDD.n1682 VDD.n620 185
R1719 VDD.n620 VDD.n617 185
R1720 VDD.n1681 VDD.n1680 185
R1721 VDD.n1680 VDD.n1679 185
R1722 VDD.n622 VDD.n621 185
R1723 VDD.n623 VDD.n622 185
R1724 VDD.n1672 VDD.n1671 185
R1725 VDD.n1673 VDD.n1672 185
R1726 VDD.n1670 VDD.n632 185
R1727 VDD.n632 VDD.n629 185
R1728 VDD.n1669 VDD.n1668 185
R1729 VDD.n1668 VDD.n1667 185
R1730 VDD.n634 VDD.n633 185
R1731 VDD.n635 VDD.n634 185
R1732 VDD.n1660 VDD.n1659 185
R1733 VDD.n1661 VDD.n1660 185
R1734 VDD.n1658 VDD.n644 185
R1735 VDD.n644 VDD.n641 185
R1736 VDD.n1657 VDD.n1656 185
R1737 VDD.n1656 VDD.n1655 185
R1738 VDD.n646 VDD.n645 185
R1739 VDD.n655 VDD.n646 185
R1740 VDD.n1647 VDD.n1646 185
R1741 VDD.n1648 VDD.n1647 185
R1742 VDD.n1645 VDD.n656 185
R1743 VDD.n662 VDD.n656 185
R1744 VDD.n1644 VDD.n1643 185
R1745 VDD.n1643 VDD.n1642 185
R1746 VDD.n658 VDD.n657 185
R1747 VDD.n659 VDD.n658 185
R1748 VDD.n1635 VDD.n1634 185
R1749 VDD.n1636 VDD.n1635 185
R1750 VDD.n1633 VDD.n669 185
R1751 VDD.n1632 VDD.n1631 185
R1752 VDD.n1629 VDD.n670 185
R1753 VDD.n1629 VDD.n666 185
R1754 VDD.n1628 VDD.n1627 185
R1755 VDD.n1626 VDD.n1625 185
R1756 VDD.n1624 VDD.n672 185
R1757 VDD.n1622 VDD.n1621 185
R1758 VDD.n1620 VDD.n673 185
R1759 VDD.n1619 VDD.n1618 185
R1760 VDD.n1616 VDD.n674 185
R1761 VDD.n1614 VDD.n1613 185
R1762 VDD.n1612 VDD.n675 185
R1763 VDD.n1611 VDD.n1610 185
R1764 VDD.n1608 VDD.n1607 185
R1765 VDD.n1606 VDD.n1605 185
R1766 VDD.n1604 VDD.n678 185
R1767 VDD.n1602 VDD.n1601 185
R1768 VDD.n1600 VDD.n679 185
R1769 VDD.n1599 VDD.n1598 185
R1770 VDD.n1596 VDD.n680 185
R1771 VDD.n1594 VDD.n1593 185
R1772 VDD.n1592 VDD.n681 185
R1773 VDD.n1591 VDD.n1590 185
R1774 VDD.n1588 VDD.n1587 185
R1775 VDD.n1586 VDD.n1585 185
R1776 VDD.n1584 VDD.n1583 185
R1777 VDD.n1584 VDD.n666 185
R1778 VDD.n1760 VDD.n1759 185
R1779 VDD.n1762 VDD.n1761 185
R1780 VDD.n1764 VDD.n1763 185
R1781 VDD.n1767 VDD.n1766 185
R1782 VDD.n1769 VDD.n1768 185
R1783 VDD.n1771 VDD.n1770 185
R1784 VDD.n1773 VDD.n1772 185
R1785 VDD.n1775 VDD.n1774 185
R1786 VDD.n1777 VDD.n1776 185
R1787 VDD.n1779 VDD.n1778 185
R1788 VDD.n1781 VDD.n1780 185
R1789 VDD.n1783 VDD.n1782 185
R1790 VDD.n1785 VDD.n1784 185
R1791 VDD.n1787 VDD.n1786 185
R1792 VDD.n1789 VDD.n1788 185
R1793 VDD.n1791 VDD.n1790 185
R1794 VDD.n1793 VDD.n1792 185
R1795 VDD.n1795 VDD.n1794 185
R1796 VDD.n1797 VDD.n1796 185
R1797 VDD.n1799 VDD.n1798 185
R1798 VDD.n1801 VDD.n1800 185
R1799 VDD.n1803 VDD.n1802 185
R1800 VDD.n1805 VDD.n1804 185
R1801 VDD.n1807 VDD.n1806 185
R1802 VDD.n1809 VDD.n1808 185
R1803 VDD.n1811 VDD.n1810 185
R1804 VDD.n1758 VDD.n1757 185
R1805 VDD.n1758 VDD.n510 185
R1806 VDD.n1756 VDD.n545 185
R1807 VDD.n1815 VDD.n545 185
R1808 VDD.n1755 VDD.n1754 185
R1809 VDD.n1754 VDD.n1753 185
R1810 VDD.n553 VDD.n552 185
R1811 VDD.n554 VDD.n553 185
R1812 VDD.n1522 VDD.n559 185
R1813 VDD.n1746 VDD.n559 185
R1814 VDD.n1524 VDD.n1523 185
R1815 VDD.n1523 VDD.n558 185
R1816 VDD.n1525 VDD.n566 185
R1817 VDD.n1739 VDD.n566 185
R1818 VDD.n1527 VDD.n1526 185
R1819 VDD.n1526 VDD.n565 185
R1820 VDD.n1528 VDD.n572 185
R1821 VDD.n1733 VDD.n572 185
R1822 VDD.n1530 VDD.n1529 185
R1823 VDD.n1529 VDD.n571 185
R1824 VDD.n1531 VDD.n577 185
R1825 VDD.n1727 VDD.n577 185
R1826 VDD.n1533 VDD.n1532 185
R1827 VDD.n1532 VDD.n585 185
R1828 VDD.n1534 VDD.n583 185
R1829 VDD.n1721 VDD.n583 185
R1830 VDD.n1536 VDD.n1535 185
R1831 VDD.n1535 VDD.n582 185
R1832 VDD.n1537 VDD.n589 185
R1833 VDD.n1715 VDD.n589 185
R1834 VDD.n1539 VDD.n1538 185
R1835 VDD.n1540 VDD.n1539 185
R1836 VDD.n1521 VDD.n595 185
R1837 VDD.n1709 VDD.n595 185
R1838 VDD.n1520 VDD.n1519 185
R1839 VDD.n1519 VDD.n594 185
R1840 VDD.n686 VDD.n600 185
R1841 VDD.n1703 VDD.n600 185
R1842 VDD.n1551 VDD.n1550 185
R1843 VDD.n1550 VDD.n1549 185
R1844 VDD.n1552 VDD.n606 185
R1845 VDD.n1697 VDD.n606 185
R1846 VDD.n1554 VDD.n1553 185
R1847 VDD.n1553 VDD.n605 185
R1848 VDD.n1555 VDD.n612 185
R1849 VDD.n1691 VDD.n612 185
R1850 VDD.n1557 VDD.n1556 185
R1851 VDD.n1556 VDD.n611 185
R1852 VDD.n1558 VDD.n618 185
R1853 VDD.n1685 VDD.n618 185
R1854 VDD.n1560 VDD.n1559 185
R1855 VDD.n1559 VDD.n617 185
R1856 VDD.n1561 VDD.n624 185
R1857 VDD.n1679 VDD.n624 185
R1858 VDD.n1563 VDD.n1562 185
R1859 VDD.n1562 VDD.n623 185
R1860 VDD.n1564 VDD.n630 185
R1861 VDD.n1673 VDD.n630 185
R1862 VDD.n1566 VDD.n1565 185
R1863 VDD.n1565 VDD.n629 185
R1864 VDD.n1567 VDD.n636 185
R1865 VDD.n1667 VDD.n636 185
R1866 VDD.n1569 VDD.n1568 185
R1867 VDD.n1568 VDD.n635 185
R1868 VDD.n1570 VDD.n642 185
R1869 VDD.n1661 VDD.n642 185
R1870 VDD.n1572 VDD.n1571 185
R1871 VDD.n1571 VDD.n641 185
R1872 VDD.n1573 VDD.n647 185
R1873 VDD.n1655 VDD.n647 185
R1874 VDD.n1575 VDD.n1574 185
R1875 VDD.n1574 VDD.n655 185
R1876 VDD.n1576 VDD.n653 185
R1877 VDD.n1648 VDD.n653 185
R1878 VDD.n1578 VDD.n1577 185
R1879 VDD.n1577 VDD.n662 185
R1880 VDD.n1579 VDD.n660 185
R1881 VDD.n1642 VDD.n660 185
R1882 VDD.n1581 VDD.n1580 185
R1883 VDD.n1580 VDD.n659 185
R1884 VDD.n1582 VDD.n667 185
R1885 VDD.n1636 VDD.n667 185
R1886 VDD.n2697 VDD.n2696 185
R1887 VDD.n2698 VDD.n2697 185
R1888 VDD.n94 VDD.n93 185
R1889 VDD.n2699 VDD.n94 185
R1890 VDD.n2702 VDD.n2701 185
R1891 VDD.n2701 VDD.n2700 185
R1892 VDD.n2703 VDD.n88 185
R1893 VDD.n88 VDD.n87 185
R1894 VDD.n2705 VDD.n2704 185
R1895 VDD.n2706 VDD.n2705 185
R1896 VDD.n83 VDD.n82 185
R1897 VDD.n2707 VDD.n83 185
R1898 VDD.n2710 VDD.n2709 185
R1899 VDD.n2709 VDD.n2708 185
R1900 VDD.n2711 VDD.n77 185
R1901 VDD.n77 VDD.n76 185
R1902 VDD.n2713 VDD.n2712 185
R1903 VDD.n2714 VDD.n2713 185
R1904 VDD.n71 VDD.n70 185
R1905 VDD.n2715 VDD.n71 185
R1906 VDD.n2718 VDD.n2717 185
R1907 VDD.n2717 VDD.n2716 185
R1908 VDD.n2719 VDD.n65 185
R1909 VDD.n72 VDD.n65 185
R1910 VDD.n2721 VDD.n2720 185
R1911 VDD.n2722 VDD.n2721 185
R1912 VDD.n61 VDD.n60 185
R1913 VDD.n2723 VDD.n61 185
R1914 VDD.n2726 VDD.n2725 185
R1915 VDD.n2725 VDD.n2724 185
R1916 VDD.n2727 VDD.n56 185
R1917 VDD.n56 VDD.n55 185
R1918 VDD.n2729 VDD.n2728 185
R1919 VDD.n2730 VDD.n2729 185
R1920 VDD.n50 VDD.n48 185
R1921 VDD.n2731 VDD.n50 185
R1922 VDD.n2734 VDD.n2733 185
R1923 VDD.n2733 VDD.n2732 185
R1924 VDD.n49 VDD.n47 185
R1925 VDD.n51 VDD.n49 185
R1926 VDD.n2553 VDD.n2552 185
R1927 VDD.n2554 VDD.n2553 185
R1928 VDD.n223 VDD.n222 185
R1929 VDD.n222 VDD.n221 185
R1930 VDD.n2548 VDD.n2547 185
R1931 VDD.n2547 VDD.n2546 185
R1932 VDD.n226 VDD.n225 185
R1933 VDD.n233 VDD.n226 185
R1934 VDD.n2537 VDD.n2536 185
R1935 VDD.n2538 VDD.n2537 185
R1936 VDD.n235 VDD.n234 185
R1937 VDD.n234 VDD.n232 185
R1938 VDD.n2532 VDD.n2531 185
R1939 VDD.n2531 VDD.n2530 185
R1940 VDD.n238 VDD.n237 185
R1941 VDD.n239 VDD.n238 185
R1942 VDD.n2521 VDD.n2520 185
R1943 VDD.n2522 VDD.n2521 185
R1944 VDD.n247 VDD.n246 185
R1945 VDD.n246 VDD.n245 185
R1946 VDD.n2516 VDD.n2515 185
R1947 VDD.n2515 VDD.n2514 185
R1948 VDD.n250 VDD.n249 185
R1949 VDD.n257 VDD.n250 185
R1950 VDD.n2505 VDD.n2504 185
R1951 VDD.n2506 VDD.n2505 185
R1952 VDD.n259 VDD.n258 185
R1953 VDD.n258 VDD.n256 185
R1954 VDD.n2500 VDD.n2499 185
R1955 VDD.n2499 VDD.n2498 185
R1956 VDD.n262 VDD.n261 185
R1957 VDD.n263 VDD.n262 185
R1958 VDD.n2489 VDD.n2488 185
R1959 VDD.n2490 VDD.n2489 185
R1960 VDD.n271 VDD.n270 185
R1961 VDD.n270 VDD.n269 185
R1962 VDD.n2484 VDD.n2483 185
R1963 VDD.n274 VDD.n273 185
R1964 VDD.n2480 VDD.n2479 185
R1965 VDD.n2481 VDD.n2480 185
R1966 VDD.n2478 VDD.n304 185
R1967 VDD.n2477 VDD.n2476 185
R1968 VDD.n2475 VDD.n2474 185
R1969 VDD.n311 VDD.n308 185
R1970 VDD.n313 VDD.n312 185
R1971 VDD.n2470 VDD.n314 185
R1972 VDD.n2469 VDD.n2468 185
R1973 VDD.n2467 VDD.n2466 185
R1974 VDD.n2465 VDD.n2464 185
R1975 VDD.n2463 VDD.n2462 185
R1976 VDD.n2461 VDD.n2460 185
R1977 VDD.n2459 VDD.n2458 185
R1978 VDD.n2457 VDD.n2456 185
R1979 VDD.n2455 VDD.n2454 185
R1980 VDD.n2453 VDD.n2452 185
R1981 VDD.n2444 VDD.n322 185
R1982 VDD.n2446 VDD.n2445 185
R1983 VDD.n2443 VDD.n2442 185
R1984 VDD.n2441 VDD.n2440 185
R1985 VDD.n2439 VDD.n2438 185
R1986 VDD.n2437 VDD.n2436 185
R1987 VDD.n2435 VDD.n2434 185
R1988 VDD.n2433 VDD.n2432 185
R1989 VDD.n2431 VDD.n2430 185
R1990 VDD.n2429 VDD.n2428 185
R1991 VDD.n2427 VDD.n2426 185
R1992 VDD.n2425 VDD.n2424 185
R1993 VDD.n2423 VDD.n2422 185
R1994 VDD.n2421 VDD.n2420 185
R1995 VDD.n2419 VDD.n2418 185
R1996 VDD.n2417 VDD.n2416 185
R1997 VDD.n2415 VDD.n2414 185
R1998 VDD.n2413 VDD.n2412 185
R1999 VDD.n2411 VDD.n2410 185
R2000 VDD.n2409 VDD.n2408 185
R2001 VDD.n2402 VDD.n340 185
R2002 VDD.n2404 VDD.n2403 185
R2003 VDD.n2401 VDD.n2400 185
R2004 VDD.n2399 VDD.n2398 185
R2005 VDD.n2397 VDD.n2396 185
R2006 VDD.n2395 VDD.n2394 185
R2007 VDD.n2393 VDD.n2392 185
R2008 VDD.n2391 VDD.n2390 185
R2009 VDD.n2389 VDD.n2388 185
R2010 VDD.n2387 VDD.n2386 185
R2011 VDD.n2385 VDD.n2384 185
R2012 VDD.n2383 VDD.n2382 185
R2013 VDD.n2358 VDD.n352 185
R2014 VDD.n2360 VDD.n2359 185
R2015 VDD.n2378 VDD.n2361 185
R2016 VDD.n2377 VDD.n2376 185
R2017 VDD.n2375 VDD.n2374 185
R2018 VDD.n2373 VDD.n2372 185
R2019 VDD.n2371 VDD.n2370 185
R2020 VDD.n2366 VDD.n303 185
R2021 VDD.n2481 VDD.n303 185
R2022 VDD.n2590 VDD.n2589 185
R2023 VDD.n2592 VDD.n197 185
R2024 VDD.n2594 VDD.n2593 185
R2025 VDD.n2595 VDD.n192 185
R2026 VDD.n2597 VDD.n2596 185
R2027 VDD.n2599 VDD.n190 185
R2028 VDD.n2601 VDD.n2600 185
R2029 VDD.n2602 VDD.n185 185
R2030 VDD.n2604 VDD.n2603 185
R2031 VDD.n2606 VDD.n183 185
R2032 VDD.n2608 VDD.n2607 185
R2033 VDD.n2609 VDD.n178 185
R2034 VDD.n2611 VDD.n2610 185
R2035 VDD.n2613 VDD.n176 185
R2036 VDD.n2615 VDD.n2614 185
R2037 VDD.n2616 VDD.n172 185
R2038 VDD.n2618 VDD.n2617 185
R2039 VDD.n2620 VDD.n170 185
R2040 VDD.n2622 VDD.n2621 185
R2041 VDD.n165 VDD.n164 185
R2042 VDD.n2627 VDD.n2626 185
R2043 VDD.n2629 VDD.n162 185
R2044 VDD.n2631 VDD.n2630 185
R2045 VDD.n2632 VDD.n157 185
R2046 VDD.n2634 VDD.n2633 185
R2047 VDD.n2636 VDD.n155 185
R2048 VDD.n2638 VDD.n2637 185
R2049 VDD.n2639 VDD.n150 185
R2050 VDD.n2641 VDD.n2640 185
R2051 VDD.n2643 VDD.n148 185
R2052 VDD.n2645 VDD.n2644 185
R2053 VDD.n2646 VDD.n143 185
R2054 VDD.n2648 VDD.n2647 185
R2055 VDD.n2650 VDD.n141 185
R2056 VDD.n2652 VDD.n2651 185
R2057 VDD.n2653 VDD.n137 185
R2058 VDD.n2655 VDD.n2654 185
R2059 VDD.n2657 VDD.n135 185
R2060 VDD.n2659 VDD.n2658 185
R2061 VDD.n130 VDD.n129 185
R2062 VDD.n2664 VDD.n2663 185
R2063 VDD.n2666 VDD.n127 185
R2064 VDD.n2668 VDD.n2667 185
R2065 VDD.n2669 VDD.n122 185
R2066 VDD.n2671 VDD.n2670 185
R2067 VDD.n2673 VDD.n120 185
R2068 VDD.n2675 VDD.n2674 185
R2069 VDD.n2676 VDD.n115 185
R2070 VDD.n2678 VDD.n2677 185
R2071 VDD.n2680 VDD.n113 185
R2072 VDD.n2682 VDD.n2681 185
R2073 VDD.n2683 VDD.n107 185
R2074 VDD.n2685 VDD.n2684 185
R2075 VDD.n2687 VDD.n106 185
R2076 VDD.n2688 VDD.n105 185
R2077 VDD.n2691 VDD.n2690 185
R2078 VDD.n2692 VDD.n103 185
R2079 VDD.n2693 VDD.n99 185
R2080 VDD.n2586 VDD.n97 185
R2081 VDD.n2698 VDD.n97 185
R2082 VDD.n2585 VDD.n96 185
R2083 VDD.n2699 VDD.n96 185
R2084 VDD.n2584 VDD.n95 185
R2085 VDD.n2700 VDD.n95 185
R2086 VDD.n205 VDD.n204 185
R2087 VDD.n204 VDD.n87 185
R2088 VDD.n2580 VDD.n86 185
R2089 VDD.n2706 VDD.n86 185
R2090 VDD.n2579 VDD.n85 185
R2091 VDD.n2707 VDD.n85 185
R2092 VDD.n2578 VDD.n84 185
R2093 VDD.n2708 VDD.n84 185
R2094 VDD.n208 VDD.n207 185
R2095 VDD.n207 VDD.n76 185
R2096 VDD.n2574 VDD.n75 185
R2097 VDD.n2714 VDD.n75 185
R2098 VDD.n2573 VDD.n74 185
R2099 VDD.n2715 VDD.n74 185
R2100 VDD.n2572 VDD.n73 185
R2101 VDD.n2716 VDD.n73 185
R2102 VDD.n211 VDD.n210 185
R2103 VDD.n210 VDD.n72 185
R2104 VDD.n2568 VDD.n64 185
R2105 VDD.n2722 VDD.n64 185
R2106 VDD.n2567 VDD.n63 185
R2107 VDD.n2723 VDD.n63 185
R2108 VDD.n2566 VDD.n62 185
R2109 VDD.n2724 VDD.n62 185
R2110 VDD.n214 VDD.n213 185
R2111 VDD.n213 VDD.n55 185
R2112 VDD.n2562 VDD.n54 185
R2113 VDD.n2730 VDD.n54 185
R2114 VDD.n2561 VDD.n53 185
R2115 VDD.n2731 VDD.n53 185
R2116 VDD.n2560 VDD.n52 185
R2117 VDD.n2732 VDD.n52 185
R2118 VDD.n220 VDD.n216 185
R2119 VDD.n220 VDD.n51 185
R2120 VDD.n2556 VDD.n2555 185
R2121 VDD.n2555 VDD.n2554 185
R2122 VDD.n219 VDD.n218 185
R2123 VDD.n221 VDD.n219 185
R2124 VDD.n2545 VDD.n2544 185
R2125 VDD.n2546 VDD.n2545 185
R2126 VDD.n228 VDD.n227 185
R2127 VDD.n233 VDD.n227 185
R2128 VDD.n2540 VDD.n2539 185
R2129 VDD.n2539 VDD.n2538 185
R2130 VDD.n231 VDD.n230 185
R2131 VDD.n232 VDD.n231 185
R2132 VDD.n2529 VDD.n2528 185
R2133 VDD.n2530 VDD.n2529 185
R2134 VDD.n241 VDD.n240 185
R2135 VDD.n240 VDD.n239 185
R2136 VDD.n2524 VDD.n2523 185
R2137 VDD.n2523 VDD.n2522 185
R2138 VDD.n244 VDD.n243 185
R2139 VDD.n245 VDD.n244 185
R2140 VDD.n2513 VDD.n2512 185
R2141 VDD.n2514 VDD.n2513 185
R2142 VDD.n252 VDD.n251 185
R2143 VDD.n257 VDD.n251 185
R2144 VDD.n2508 VDD.n2507 185
R2145 VDD.n2507 VDD.n2506 185
R2146 VDD.n255 VDD.n254 185
R2147 VDD.n256 VDD.n255 185
R2148 VDD.n2497 VDD.n2496 185
R2149 VDD.n2498 VDD.n2497 185
R2150 VDD.n265 VDD.n264 185
R2151 VDD.n264 VDD.n263 185
R2152 VDD.n2492 VDD.n2491 185
R2153 VDD.n2491 VDD.n2490 185
R2154 VDD.n268 VDD.n267 185
R2155 VDD.n269 VDD.n268 185
R2156 VDD.n509 VDD.n508 185
R2157 VDD.n1907 VDD.n1906 185
R2158 VDD.n1908 VDD.n1904 185
R2159 VDD.n1904 VDD.n1870 185
R2160 VDD.n1910 VDD.n1909 185
R2161 VDD.n1912 VDD.n1903 185
R2162 VDD.n1915 VDD.n1914 185
R2163 VDD.n1916 VDD.n1902 185
R2164 VDD.n1918 VDD.n1917 185
R2165 VDD.n1920 VDD.n1901 185
R2166 VDD.n1923 VDD.n1922 185
R2167 VDD.n1924 VDD.n1900 185
R2168 VDD.n1926 VDD.n1925 185
R2169 VDD.n1928 VDD.n1899 185
R2170 VDD.n1931 VDD.n1930 185
R2171 VDD.n1932 VDD.n1898 185
R2172 VDD.n1934 VDD.n1933 185
R2173 VDD.n1936 VDD.n1897 185
R2174 VDD.n1939 VDD.n1938 185
R2175 VDD.n1940 VDD.n1896 185
R2176 VDD.n1942 VDD.n1941 185
R2177 VDD.n1944 VDD.n1895 185
R2178 VDD.n1947 VDD.n1946 185
R2179 VDD.n1948 VDD.n1892 185
R2180 VDD.n1951 VDD.n1950 185
R2181 VDD.n1953 VDD.n1891 185
R2182 VDD.n1955 VDD.n1954 185
R2183 VDD.n1954 VDD.n1870 185
R2184 VDD.n2283 VDD.n2282 185
R2185 VDD.n2285 VDD.n393 185
R2186 VDD.n2287 VDD.n2286 185
R2187 VDD.n2289 VDD.n390 185
R2188 VDD.n2291 VDD.n2290 185
R2189 VDD.n2293 VDD.n388 185
R2190 VDD.n2295 VDD.n2294 185
R2191 VDD.n2296 VDD.n387 185
R2192 VDD.n2298 VDD.n2297 185
R2193 VDD.n2300 VDD.n385 185
R2194 VDD.n2302 VDD.n2301 185
R2195 VDD.n2303 VDD.n384 185
R2196 VDD.n2305 VDD.n2304 185
R2197 VDD.n2308 VDD.n2307 185
R2198 VDD.n2310 VDD.n2309 185
R2199 VDD.n2312 VDD.n382 185
R2200 VDD.n2314 VDD.n2313 185
R2201 VDD.n2315 VDD.n381 185
R2202 VDD.n2317 VDD.n2316 185
R2203 VDD.n2319 VDD.n379 185
R2204 VDD.n2321 VDD.n2320 185
R2205 VDD.n2322 VDD.n378 185
R2206 VDD.n2324 VDD.n2323 185
R2207 VDD.n2326 VDD.n376 185
R2208 VDD.n2328 VDD.n2327 185
R2209 VDD.n2329 VDD.n374 185
R2210 VDD.n2281 VDD.n371 185
R2211 VDD.n2332 VDD.n371 185
R2212 VDD.n2280 VDD.n2279 185
R2213 VDD.n2279 VDD.n370 185
R2214 VDD.n2278 VDD.n395 185
R2215 VDD.n2278 VDD.n2277 185
R2216 VDD.n1978 VDD.n396 185
R2217 VDD.n397 VDD.n396 185
R2218 VDD.n1979 VDD.n404 185
R2219 VDD.n2271 VDD.n404 185
R2220 VDD.n1981 VDD.n1980 185
R2221 VDD.n1980 VDD.n403 185
R2222 VDD.n1982 VDD.n412 185
R2223 VDD.n2228 VDD.n412 185
R2224 VDD.n1984 VDD.n1983 185
R2225 VDD.n1983 VDD.n411 185
R2226 VDD.n1985 VDD.n418 185
R2227 VDD.n2222 VDD.n418 185
R2228 VDD.n1987 VDD.n1986 185
R2229 VDD.n1986 VDD.n417 185
R2230 VDD.n1988 VDD.n423 185
R2231 VDD.n2216 VDD.n423 185
R2232 VDD.n1990 VDD.n1989 185
R2233 VDD.n1989 VDD.n430 185
R2234 VDD.n1991 VDD.n428 185
R2235 VDD.n2210 VDD.n428 185
R2236 VDD.n1993 VDD.n1992 185
R2237 VDD.n1992 VDD.n436 185
R2238 VDD.n1994 VDD.n434 185
R2239 VDD.n2204 VDD.n434 185
R2240 VDD.n1996 VDD.n1995 185
R2241 VDD.n1995 VDD.n442 185
R2242 VDD.n1997 VDD.n440 185
R2243 VDD.n2198 VDD.n440 185
R2244 VDD.n1999 VDD.n1998 185
R2245 VDD.n1998 VDD.n448 185
R2246 VDD.n2000 VDD.n446 185
R2247 VDD.n2192 VDD.n446 185
R2248 VDD.n2002 VDD.n2001 185
R2249 VDD.n2001 VDD.n454 185
R2250 VDD.n2003 VDD.n452 185
R2251 VDD.n2186 VDD.n452 185
R2252 VDD.n2040 VDD.n2039 185
R2253 VDD.n2039 VDD.n2038 185
R2254 VDD.n2041 VDD.n459 185
R2255 VDD.n2180 VDD.n459 185
R2256 VDD.n2043 VDD.n2042 185
R2257 VDD.n2042 VDD.n458 185
R2258 VDD.n2044 VDD.n464 185
R2259 VDD.n2174 VDD.n464 185
R2260 VDD.n2046 VDD.n2045 185
R2261 VDD.n2047 VDD.n2046 185
R2262 VDD.n1977 VDD.n470 185
R2263 VDD.n2168 VDD.n470 185
R2264 VDD.n1976 VDD.n1975 185
R2265 VDD.n1975 VDD.n469 185
R2266 VDD.n1974 VDD.n476 185
R2267 VDD.n2162 VDD.n476 185
R2268 VDD.n1973 VDD.n1972 185
R2269 VDD.n1972 VDD.n475 185
R2270 VDD.n1971 VDD.n481 185
R2271 VDD.n2156 VDD.n481 185
R2272 VDD.n1970 VDD.n1969 185
R2273 VDD.n1969 VDD.n489 185
R2274 VDD.n1968 VDD.n487 185
R2275 VDD.n2150 VDD.n487 185
R2276 VDD.n1967 VDD.n1966 185
R2277 VDD.n1966 VDD.n486 185
R2278 VDD.n1965 VDD.n493 185
R2279 VDD.n2144 VDD.n493 185
R2280 VDD.n1964 VDD.n1963 185
R2281 VDD.n1963 VDD.n500 185
R2282 VDD.n1962 VDD.n498 185
R2283 VDD.n2138 VDD.n498 185
R2284 VDD.n1961 VDD.n1960 185
R2285 VDD.n1960 VDD.n506 185
R2286 VDD.n1959 VDD.n504 185
R2287 VDD.n2132 VDD.n504 185
R2288 VDD.n1958 VDD.n1957 185
R2289 VDD.n1957 VDD.n1873 185
R2290 VDD.n1956 VDD.n1871 185
R2291 VDD.n2126 VDD.n1871 185
R2292 VDD.n2128 VDD.n2127 185
R2293 VDD.n2127 VDD.n2126 185
R2294 VDD.n2129 VDD.n507 185
R2295 VDD.n1873 VDD.n507 185
R2296 VDD.n2131 VDD.n2130 185
R2297 VDD.n2132 VDD.n2131 185
R2298 VDD.n497 VDD.n496 185
R2299 VDD.n506 VDD.n497 185
R2300 VDD.n2140 VDD.n2139 185
R2301 VDD.n2139 VDD.n2138 185
R2302 VDD.n2141 VDD.n495 185
R2303 VDD.n500 VDD.n495 185
R2304 VDD.n2143 VDD.n2142 185
R2305 VDD.n2144 VDD.n2143 185
R2306 VDD.n485 VDD.n484 185
R2307 VDD.n486 VDD.n485 185
R2308 VDD.n2152 VDD.n2151 185
R2309 VDD.n2151 VDD.n2150 185
R2310 VDD.n2153 VDD.n483 185
R2311 VDD.n489 VDD.n483 185
R2312 VDD.n2155 VDD.n2154 185
R2313 VDD.n2156 VDD.n2155 185
R2314 VDD.n474 VDD.n473 185
R2315 VDD.n475 VDD.n474 185
R2316 VDD.n2164 VDD.n2163 185
R2317 VDD.n2163 VDD.n2162 185
R2318 VDD.n2165 VDD.n472 185
R2319 VDD.n472 VDD.n469 185
R2320 VDD.n2167 VDD.n2166 185
R2321 VDD.n2168 VDD.n2167 185
R2322 VDD.n463 VDD.n462 185
R2323 VDD.n2047 VDD.n463 185
R2324 VDD.n2176 VDD.n2175 185
R2325 VDD.n2175 VDD.n2174 185
R2326 VDD.n2177 VDD.n461 185
R2327 VDD.n461 VDD.n458 185
R2328 VDD.n2179 VDD.n2178 185
R2329 VDD.n2180 VDD.n2179 185
R2330 VDD.n451 VDD.n450 185
R2331 VDD.n2038 VDD.n451 185
R2332 VDD.n2188 VDD.n2187 185
R2333 VDD.n2187 VDD.n2186 185
R2334 VDD.n2189 VDD.n449 185
R2335 VDD.n454 VDD.n449 185
R2336 VDD.n2191 VDD.n2190 185
R2337 VDD.n2192 VDD.n2191 185
R2338 VDD.n439 VDD.n438 185
R2339 VDD.n448 VDD.n439 185
R2340 VDD.n2200 VDD.n2199 185
R2341 VDD.n2199 VDD.n2198 185
R2342 VDD.n2201 VDD.n437 185
R2343 VDD.n442 VDD.n437 185
R2344 VDD.n2203 VDD.n2202 185
R2345 VDD.n2204 VDD.n2203 185
R2346 VDD.n427 VDD.n426 185
R2347 VDD.n436 VDD.n427 185
R2348 VDD.n2212 VDD.n2211 185
R2349 VDD.n2211 VDD.n2210 185
R2350 VDD.n2213 VDD.n425 185
R2351 VDD.n430 VDD.n425 185
R2352 VDD.n2215 VDD.n2214 185
R2353 VDD.n2216 VDD.n2215 185
R2354 VDD.n416 VDD.n415 185
R2355 VDD.n417 VDD.n416 185
R2356 VDD.n2224 VDD.n2223 185
R2357 VDD.n2223 VDD.n2222 185
R2358 VDD.n2225 VDD.n414 185
R2359 VDD.n414 VDD.n411 185
R2360 VDD.n2227 VDD.n2226 185
R2361 VDD.n2228 VDD.n2227 185
R2362 VDD.n402 VDD.n401 185
R2363 VDD.n403 VDD.n402 185
R2364 VDD.n2273 VDD.n2272 185
R2365 VDD.n2272 VDD.n2271 185
R2366 VDD.n2274 VDD.n400 185
R2367 VDD.n400 VDD.n397 185
R2368 VDD.n2276 VDD.n2275 185
R2369 VDD.n2277 VDD.n2276 185
R2370 VDD.n375 VDD.n373 185
R2371 VDD.n373 VDD.n370 185
R2372 VDD.n2331 VDD.n2330 185
R2373 VDD.n2332 VDD.n2331 185
R2374 VDD.n539 VDD.n537 185
R2375 VDD.n537 VDD.n510 185
R2376 VDD.n1750 VDD.n546 185
R2377 VDD.n1815 VDD.n546 185
R2378 VDD.n1752 VDD.n1751 185
R2379 VDD.n1753 VDD.n1752 185
R2380 VDD.n1749 VDD.n555 185
R2381 VDD.n555 VDD.n554 185
R2382 VDD.n1748 VDD.n1747 185
R2383 VDD.n1747 VDD.n1746 185
R2384 VDD.n557 VDD.n556 185
R2385 VDD.n558 VDD.n557 185
R2386 VDD.n1738 VDD.n1737 185
R2387 VDD.n1739 VDD.n1738 185
R2388 VDD.n1736 VDD.n568 185
R2389 VDD.n568 VDD.n565 185
R2390 VDD.n1735 VDD.n1734 185
R2391 VDD.n1734 VDD.n1733 185
R2392 VDD.n570 VDD.n569 185
R2393 VDD.n571 VDD.n570 185
R2394 VDD.n1726 VDD.n1725 185
R2395 VDD.n1727 VDD.n1726 185
R2396 VDD.n1724 VDD.n579 185
R2397 VDD.n585 VDD.n579 185
R2398 VDD.n1723 VDD.n1722 185
R2399 VDD.n1722 VDD.n1721 185
R2400 VDD.n581 VDD.n580 185
R2401 VDD.n582 VDD.n581 185
R2402 VDD.n1714 VDD.n1713 185
R2403 VDD.n1715 VDD.n1714 185
R2404 VDD.n1712 VDD.n591 185
R2405 VDD.n1540 VDD.n591 185
R2406 VDD.n1711 VDD.n1710 185
R2407 VDD.n1710 VDD.n1709 185
R2408 VDD.n593 VDD.n592 185
R2409 VDD.n594 VDD.n593 185
R2410 VDD.n1702 VDD.n1701 185
R2411 VDD.n1703 VDD.n1702 185
R2412 VDD.n1700 VDD.n602 185
R2413 VDD.n1549 VDD.n602 185
R2414 VDD.n1699 VDD.n1698 185
R2415 VDD.n1698 VDD.n1697 185
R2416 VDD.n604 VDD.n603 185
R2417 VDD.n605 VDD.n604 185
R2418 VDD.n1690 VDD.n1689 185
R2419 VDD.n1691 VDD.n1690 185
R2420 VDD.n1688 VDD.n614 185
R2421 VDD.n614 VDD.n611 185
R2422 VDD.n1687 VDD.n1686 185
R2423 VDD.n1686 VDD.n1685 185
R2424 VDD.n616 VDD.n615 185
R2425 VDD.n617 VDD.n616 185
R2426 VDD.n1678 VDD.n1677 185
R2427 VDD.n1679 VDD.n1678 185
R2428 VDD.n1676 VDD.n626 185
R2429 VDD.n626 VDD.n623 185
R2430 VDD.n1675 VDD.n1674 185
R2431 VDD.n1674 VDD.n1673 185
R2432 VDD.n628 VDD.n627 185
R2433 VDD.n629 VDD.n628 185
R2434 VDD.n1666 VDD.n1665 185
R2435 VDD.n1667 VDD.n1666 185
R2436 VDD.n1664 VDD.n638 185
R2437 VDD.n638 VDD.n635 185
R2438 VDD.n1663 VDD.n1662 185
R2439 VDD.n1662 VDD.n1661 185
R2440 VDD.n640 VDD.n639 185
R2441 VDD.n641 VDD.n640 185
R2442 VDD.n1654 VDD.n1653 185
R2443 VDD.n1655 VDD.n1654 185
R2444 VDD.n1651 VDD.n649 185
R2445 VDD.n655 VDD.n649 185
R2446 VDD.n1650 VDD.n1649 185
R2447 VDD.n1649 VDD.n1648 185
R2448 VDD.n652 VDD.n651 185
R2449 VDD.n662 VDD.n652 185
R2450 VDD.n1641 VDD.n1640 185
R2451 VDD.n1642 VDD.n1641 185
R2452 VDD.n1639 VDD.n663 185
R2453 VDD.n663 VDD.n659 185
R2454 VDD.n1638 VDD.n1637 185
R2455 VDD.n1637 VDD.n1636 185
R2456 VDD.n1819 VDD.n536 185
R2457 VDD.n1869 VDD.n536 185
R2458 VDD.n1821 VDD.n1820 185
R2459 VDD.n1823 VDD.n1822 185
R2460 VDD.n1825 VDD.n1824 185
R2461 VDD.n1827 VDD.n1826 185
R2462 VDD.n1829 VDD.n1828 185
R2463 VDD.n1831 VDD.n1830 185
R2464 VDD.n1833 VDD.n1832 185
R2465 VDD.n1835 VDD.n1834 185
R2466 VDD.n1837 VDD.n1836 185
R2467 VDD.n1839 VDD.n1838 185
R2468 VDD.n1841 VDD.n1840 185
R2469 VDD.n1843 VDD.n1842 185
R2470 VDD.n1845 VDD.n1844 185
R2471 VDD.n1847 VDD.n1846 185
R2472 VDD.n1849 VDD.n1848 185
R2473 VDD.n1851 VDD.n1850 185
R2474 VDD.n1853 VDD.n1852 185
R2475 VDD.n1855 VDD.n1854 185
R2476 VDD.n1857 VDD.n1856 185
R2477 VDD.n1859 VDD.n1858 185
R2478 VDD.n1861 VDD.n1860 185
R2479 VDD.n1863 VDD.n1862 185
R2480 VDD.n1865 VDD.n1864 185
R2481 VDD.n1866 VDD.n538 185
R2482 VDD.n1868 VDD.n1867 185
R2483 VDD.n1869 VDD.n1868 185
R2484 VDD.n1818 VDD.n1817 185
R2485 VDD.n1817 VDD.n510 185
R2486 VDD.n1816 VDD.n543 185
R2487 VDD.n1816 VDD.n1815 185
R2488 VDD.n1500 VDD.n544 185
R2489 VDD.n1753 VDD.n544 185
R2490 VDD.n1502 VDD.n1501 185
R2491 VDD.n1501 VDD.n554 185
R2492 VDD.n1503 VDD.n560 185
R2493 VDD.n1746 VDD.n560 185
R2494 VDD.n1505 VDD.n1504 185
R2495 VDD.n1504 VDD.n558 185
R2496 VDD.n1506 VDD.n567 185
R2497 VDD.n1739 VDD.n567 185
R2498 VDD.n1508 VDD.n1507 185
R2499 VDD.n1507 VDD.n565 185
R2500 VDD.n1509 VDD.n573 185
R2501 VDD.n1733 VDD.n573 185
R2502 VDD.n1511 VDD.n1510 185
R2503 VDD.n1510 VDD.n571 185
R2504 VDD.n1512 VDD.n578 185
R2505 VDD.n1727 VDD.n578 185
R2506 VDD.n1514 VDD.n1513 185
R2507 VDD.n1513 VDD.n585 185
R2508 VDD.n1515 VDD.n584 185
R2509 VDD.n1721 VDD.n584 185
R2510 VDD.n1517 VDD.n1516 185
R2511 VDD.n1516 VDD.n582 185
R2512 VDD.n1518 VDD.n590 185
R2513 VDD.n1715 VDD.n590 185
R2514 VDD.n1542 VDD.n1541 185
R2515 VDD.n1541 VDD.n1540 185
R2516 VDD.n1543 VDD.n596 185
R2517 VDD.n1709 VDD.n596 185
R2518 VDD.n1545 VDD.n1544 185
R2519 VDD.n1544 VDD.n594 185
R2520 VDD.n1546 VDD.n601 185
R2521 VDD.n1703 VDD.n601 185
R2522 VDD.n1548 VDD.n1547 185
R2523 VDD.n1549 VDD.n1548 185
R2524 VDD.n1499 VDD.n607 185
R2525 VDD.n1697 VDD.n607 185
R2526 VDD.n1498 VDD.n1497 185
R2527 VDD.n1497 VDD.n605 185
R2528 VDD.n1496 VDD.n613 185
R2529 VDD.n1691 VDD.n613 185
R2530 VDD.n1495 VDD.n1494 185
R2531 VDD.n1494 VDD.n611 185
R2532 VDD.n1493 VDD.n619 185
R2533 VDD.n1685 VDD.n619 185
R2534 VDD.n1492 VDD.n1491 185
R2535 VDD.n1491 VDD.n617 185
R2536 VDD.n1490 VDD.n625 185
R2537 VDD.n1679 VDD.n625 185
R2538 VDD.n1489 VDD.n1488 185
R2539 VDD.n1488 VDD.n623 185
R2540 VDD.n1487 VDD.n631 185
R2541 VDD.n1673 VDD.n631 185
R2542 VDD.n1486 VDD.n1485 185
R2543 VDD.n1485 VDD.n629 185
R2544 VDD.n1484 VDD.n637 185
R2545 VDD.n1667 VDD.n637 185
R2546 VDD.n1483 VDD.n1482 185
R2547 VDD.n1482 VDD.n635 185
R2548 VDD.n1481 VDD.n643 185
R2549 VDD.n1661 VDD.n643 185
R2550 VDD.n1480 VDD.n1479 185
R2551 VDD.n1479 VDD.n641 185
R2552 VDD.n1478 VDD.n648 185
R2553 VDD.n1655 VDD.n648 185
R2554 VDD.n1477 VDD.n1476 185
R2555 VDD.n1476 VDD.n655 185
R2556 VDD.n1475 VDD.n654 185
R2557 VDD.n1648 VDD.n654 185
R2558 VDD.n1474 VDD.n1473 185
R2559 VDD.n1473 VDD.n662 185
R2560 VDD.n1472 VDD.n661 185
R2561 VDD.n1642 VDD.n661 185
R2562 VDD.n1471 VDD.n1470 185
R2563 VDD.n1470 VDD.n659 185
R2564 VDD.n1469 VDD.n668 185
R2565 VDD.n1636 VDD.n668 185
R2566 VDD.n665 VDD.n664 185
R2567 VDD.n666 VDD.n665 185
R2568 VDD.n1420 VDD.n1419 185
R2569 VDD.n1421 VDD.n1417 185
R2570 VDD.n1423 VDD.n1422 185
R2571 VDD.n1425 VDD.n1416 185
R2572 VDD.n1428 VDD.n1427 185
R2573 VDD.n1429 VDD.n1415 185
R2574 VDD.n1431 VDD.n1430 185
R2575 VDD.n1433 VDD.n1414 185
R2576 VDD.n1436 VDD.n1435 185
R2577 VDD.n1437 VDD.n1413 185
R2578 VDD.n1439 VDD.n1438 185
R2579 VDD.n1441 VDD.n1412 185
R2580 VDD.n1444 VDD.n1443 185
R2581 VDD.n1445 VDD.n694 185
R2582 VDD.n1447 VDD.n1446 185
R2583 VDD.n1449 VDD.n693 185
R2584 VDD.n1452 VDD.n1451 185
R2585 VDD.n1453 VDD.n692 185
R2586 VDD.n1455 VDD.n1454 185
R2587 VDD.n1457 VDD.n691 185
R2588 VDD.n1460 VDD.n1459 185
R2589 VDD.n1461 VDD.n688 185
R2590 VDD.n1464 VDD.n1463 185
R2591 VDD.n1466 VDD.n687 185
R2592 VDD.n1468 VDD.n1467 185
R2593 VDD.n1467 VDD.n666 185
R2594 VDD.n714 VDD.n666 151.596
R2595 VDD.n2481 VDD.n275 151.596
R2596 VDD.n2690 VDD.n103 146.341
R2597 VDD.n2688 VDD.n2687 146.341
R2598 VDD.n2685 VDD.n107 146.341
R2599 VDD.n2681 VDD.n2680 146.341
R2600 VDD.n2678 VDD.n115 146.341
R2601 VDD.n2674 VDD.n2673 146.341
R2602 VDD.n2671 VDD.n122 146.341
R2603 VDD.n2667 VDD.n2666 146.341
R2604 VDD.n2664 VDD.n129 146.341
R2605 VDD.n2658 VDD.n2657 146.341
R2606 VDD.n2655 VDD.n137 146.341
R2607 VDD.n2651 VDD.n2650 146.341
R2608 VDD.n2648 VDD.n143 146.341
R2609 VDD.n2644 VDD.n2643 146.341
R2610 VDD.n2641 VDD.n150 146.341
R2611 VDD.n2637 VDD.n2636 146.341
R2612 VDD.n2634 VDD.n157 146.341
R2613 VDD.n2630 VDD.n2629 146.341
R2614 VDD.n2627 VDD.n164 146.341
R2615 VDD.n2621 VDD.n2620 146.341
R2616 VDD.n2618 VDD.n172 146.341
R2617 VDD.n2614 VDD.n2613 146.341
R2618 VDD.n2611 VDD.n178 146.341
R2619 VDD.n2607 VDD.n2606 146.341
R2620 VDD.n2604 VDD.n185 146.341
R2621 VDD.n2600 VDD.n2599 146.341
R2622 VDD.n2597 VDD.n192 146.341
R2623 VDD.n2593 VDD.n2592 146.341
R2624 VDD.n2491 VDD.n268 146.341
R2625 VDD.n2491 VDD.n264 146.341
R2626 VDD.n2497 VDD.n264 146.341
R2627 VDD.n2497 VDD.n255 146.341
R2628 VDD.n2507 VDD.n255 146.341
R2629 VDD.n2507 VDD.n251 146.341
R2630 VDD.n2513 VDD.n251 146.341
R2631 VDD.n2513 VDD.n244 146.341
R2632 VDD.n2523 VDD.n244 146.341
R2633 VDD.n2523 VDD.n240 146.341
R2634 VDD.n2529 VDD.n240 146.341
R2635 VDD.n2529 VDD.n231 146.341
R2636 VDD.n2539 VDD.n231 146.341
R2637 VDD.n2539 VDD.n227 146.341
R2638 VDD.n2545 VDD.n227 146.341
R2639 VDD.n2545 VDD.n219 146.341
R2640 VDD.n2555 VDD.n219 146.341
R2641 VDD.n2555 VDD.n220 146.341
R2642 VDD.n220 VDD.n52 146.341
R2643 VDD.n53 VDD.n52 146.341
R2644 VDD.n54 VDD.n53 146.341
R2645 VDD.n213 VDD.n54 146.341
R2646 VDD.n213 VDD.n62 146.341
R2647 VDD.n63 VDD.n62 146.341
R2648 VDD.n64 VDD.n63 146.341
R2649 VDD.n210 VDD.n64 146.341
R2650 VDD.n210 VDD.n73 146.341
R2651 VDD.n74 VDD.n73 146.341
R2652 VDD.n75 VDD.n74 146.341
R2653 VDD.n207 VDD.n75 146.341
R2654 VDD.n207 VDD.n84 146.341
R2655 VDD.n85 VDD.n84 146.341
R2656 VDD.n86 VDD.n85 146.341
R2657 VDD.n204 VDD.n86 146.341
R2658 VDD.n204 VDD.n95 146.341
R2659 VDD.n96 VDD.n95 146.341
R2660 VDD.n97 VDD.n96 146.341
R2661 VDD.n2480 VDD.n274 146.341
R2662 VDD.n2480 VDD.n304 146.341
R2663 VDD.n2476 VDD.n2475 146.341
R2664 VDD.n312 VDD.n311 146.341
R2665 VDD.n2468 VDD.n314 146.341
R2666 VDD.n2466 VDD.n2465 146.341
R2667 VDD.n2462 VDD.n2461 146.341
R2668 VDD.n2458 VDD.n2457 146.341
R2669 VDD.n2454 VDD.n2453 146.341
R2670 VDD.n2445 VDD.n2444 146.341
R2671 VDD.n2442 VDD.n2441 146.341
R2672 VDD.n2438 VDD.n2437 146.341
R2673 VDD.n2434 VDD.n2433 146.341
R2674 VDD.n2430 VDD.n2429 146.341
R2675 VDD.n2426 VDD.n2425 146.341
R2676 VDD.n2422 VDD.n2421 146.341
R2677 VDD.n2418 VDD.n2417 146.341
R2678 VDD.n2414 VDD.n2413 146.341
R2679 VDD.n2410 VDD.n2409 146.341
R2680 VDD.n2403 VDD.n2402 146.341
R2681 VDD.n2400 VDD.n2399 146.341
R2682 VDD.n2396 VDD.n2395 146.341
R2683 VDD.n2392 VDD.n2391 146.341
R2684 VDD.n2388 VDD.n2387 146.341
R2685 VDD.n2384 VDD.n2383 146.341
R2686 VDD.n2359 VDD.n2358 146.341
R2687 VDD.n2376 VDD.n2361 146.341
R2688 VDD.n2374 VDD.n2373 146.341
R2689 VDD.n2370 VDD.n303 146.341
R2690 VDD.n2489 VDD.n270 146.341
R2691 VDD.n2489 VDD.n262 146.341
R2692 VDD.n2499 VDD.n262 146.341
R2693 VDD.n2499 VDD.n258 146.341
R2694 VDD.n2505 VDD.n258 146.341
R2695 VDD.n2505 VDD.n250 146.341
R2696 VDD.n2515 VDD.n250 146.341
R2697 VDD.n2515 VDD.n246 146.341
R2698 VDD.n2521 VDD.n246 146.341
R2699 VDD.n2521 VDD.n238 146.341
R2700 VDD.n2531 VDD.n238 146.341
R2701 VDD.n2531 VDD.n234 146.341
R2702 VDD.n2537 VDD.n234 146.341
R2703 VDD.n2537 VDD.n226 146.341
R2704 VDD.n2547 VDD.n226 146.341
R2705 VDD.n2547 VDD.n222 146.341
R2706 VDD.n2553 VDD.n222 146.341
R2707 VDD.n2553 VDD.n49 146.341
R2708 VDD.n2733 VDD.n49 146.341
R2709 VDD.n2733 VDD.n50 146.341
R2710 VDD.n2729 VDD.n50 146.341
R2711 VDD.n2729 VDD.n56 146.341
R2712 VDD.n2725 VDD.n56 146.341
R2713 VDD.n2725 VDD.n61 146.341
R2714 VDD.n2721 VDD.n61 146.341
R2715 VDD.n2721 VDD.n65 146.341
R2716 VDD.n2717 VDD.n65 146.341
R2717 VDD.n2717 VDD.n71 146.341
R2718 VDD.n2713 VDD.n71 146.341
R2719 VDD.n2713 VDD.n77 146.341
R2720 VDD.n2709 VDD.n77 146.341
R2721 VDD.n2709 VDD.n83 146.341
R2722 VDD.n2705 VDD.n83 146.341
R2723 VDD.n2705 VDD.n88 146.341
R2724 VDD.n2701 VDD.n88 146.341
R2725 VDD.n2701 VDD.n94 146.341
R2726 VDD.n2697 VDD.n94 146.341
R2727 VDD.n1392 VDD.n1391 146.341
R2728 VDD.n1389 VDD.n1217 146.341
R2729 VDD.n1226 VDD.n1222 146.341
R2730 VDD.n1381 VDD.n1380 146.341
R2731 VDD.n1378 VDD.n1228 146.341
R2732 VDD.n1374 VDD.n1373 146.341
R2733 VDD.n1371 VDD.n1233 146.341
R2734 VDD.n1367 VDD.n1366 146.341
R2735 VDD.n1364 VDD.n1240 146.341
R2736 VDD.n1358 VDD.n1357 146.341
R2737 VDD.n1355 VDD.n1248 146.341
R2738 VDD.n1351 VDD.n1350 146.341
R2739 VDD.n1348 VDD.n1254 146.341
R2740 VDD.n1344 VDD.n1343 146.341
R2741 VDD.n1341 VDD.n1261 146.341
R2742 VDD.n1337 VDD.n1336 146.341
R2743 VDD.n1334 VDD.n1268 146.341
R2744 VDD.n1330 VDD.n1329 146.341
R2745 VDD.n1327 VDD.n1275 146.341
R2746 VDD.n1321 VDD.n1320 146.341
R2747 VDD.n1318 VDD.n1283 146.341
R2748 VDD.n1314 VDD.n1313 146.341
R2749 VDD.n1311 VDD.n1289 146.341
R2750 VDD.n1307 VDD.n1306 146.341
R2751 VDD.n1304 VDD.n1302 146.341
R2752 VDD.n1300 VDD.n1298 146.341
R2753 VDD.n701 VDD.n700 146.341
R2754 VDD.n708 VDD.n702 146.341
R2755 VDD.n1072 VDD.n853 146.341
R2756 VDD.n1072 VDD.n849 146.341
R2757 VDD.n1078 VDD.n849 146.341
R2758 VDD.n1078 VDD.n840 146.341
R2759 VDD.n1088 VDD.n840 146.341
R2760 VDD.n1088 VDD.n836 146.341
R2761 VDD.n1094 VDD.n836 146.341
R2762 VDD.n1094 VDD.n829 146.341
R2763 VDD.n1104 VDD.n829 146.341
R2764 VDD.n1104 VDD.n825 146.341
R2765 VDD.n1110 VDD.n825 146.341
R2766 VDD.n1110 VDD.n816 146.341
R2767 VDD.n1120 VDD.n816 146.341
R2768 VDD.n1120 VDD.n812 146.341
R2769 VDD.n1126 VDD.n812 146.341
R2770 VDD.n1126 VDD.n805 146.341
R2771 VDD.n1137 VDD.n805 146.341
R2772 VDD.n1137 VDD.n801 146.341
R2773 VDD.n1143 VDD.n801 146.341
R2774 VDD.n1143 VDD.n762 146.341
R2775 VDD.n1153 VDD.n762 146.341
R2776 VDD.n1153 VDD.n758 146.341
R2777 VDD.n1159 VDD.n758 146.341
R2778 VDD.n1159 VDD.n751 146.341
R2779 VDD.n1169 VDD.n751 146.341
R2780 VDD.n1169 VDD.n747 146.341
R2781 VDD.n1175 VDD.n747 146.341
R2782 VDD.n1175 VDD.n738 146.341
R2783 VDD.n1185 VDD.n738 146.341
R2784 VDD.n1185 VDD.n734 146.341
R2785 VDD.n1191 VDD.n734 146.341
R2786 VDD.n1191 VDD.n727 146.341
R2787 VDD.n1201 VDD.n727 146.341
R2788 VDD.n1201 VDD.n722 146.341
R2789 VDD.n1208 VDD.n722 146.341
R2790 VDD.n1208 VDD.n710 146.341
R2791 VDD.n1400 VDD.n710 146.341
R2792 VDD.n1061 VDD.n859 146.341
R2793 VDD.n1061 VDD.n888 146.341
R2794 VDD.n892 VDD.n891 146.341
R2795 VDD.n894 VDD.n893 146.341
R2796 VDD.n898 VDD.n897 146.341
R2797 VDD.n900 VDD.n899 146.341
R2798 VDD.n904 VDD.n903 146.341
R2799 VDD.n906 VDD.n905 146.341
R2800 VDD.n1034 VDD.n909 146.341
R2801 VDD.n911 VDD.n910 146.341
R2802 VDD.n915 VDD.n914 146.341
R2803 VDD.n917 VDD.n916 146.341
R2804 VDD.n921 VDD.n920 146.341
R2805 VDD.n923 VDD.n922 146.341
R2806 VDD.n927 VDD.n926 146.341
R2807 VDD.n929 VDD.n928 146.341
R2808 VDD.n933 VDD.n932 146.341
R2809 VDD.n935 VDD.n934 146.341
R2810 VDD.n1001 VDD.n938 146.341
R2811 VDD.n940 VDD.n939 146.341
R2812 VDD.n944 VDD.n943 146.341
R2813 VDD.n946 VDD.n945 146.341
R2814 VDD.n950 VDD.n949 146.341
R2815 VDD.n952 VDD.n951 146.341
R2816 VDD.n956 VDD.n955 146.341
R2817 VDD.n958 VDD.n957 146.341
R2818 VDD.n962 VDD.n961 146.341
R2819 VDD.n964 VDD.n963 146.341
R2820 VDD.n967 VDD.n887 146.341
R2821 VDD.n1070 VDD.n855 146.341
R2822 VDD.n1070 VDD.n847 146.341
R2823 VDD.n1080 VDD.n847 146.341
R2824 VDD.n1080 VDD.n843 146.341
R2825 VDD.n1086 VDD.n843 146.341
R2826 VDD.n1086 VDD.n835 146.341
R2827 VDD.n1096 VDD.n835 146.341
R2828 VDD.n1096 VDD.n831 146.341
R2829 VDD.n1102 VDD.n831 146.341
R2830 VDD.n1102 VDD.n823 146.341
R2831 VDD.n1112 VDD.n823 146.341
R2832 VDD.n1112 VDD.n819 146.341
R2833 VDD.n1118 VDD.n819 146.341
R2834 VDD.n1118 VDD.n811 146.341
R2835 VDD.n1128 VDD.n811 146.341
R2836 VDD.n1128 VDD.n807 146.341
R2837 VDD.n1135 VDD.n807 146.341
R2838 VDD.n1135 VDD.n799 146.341
R2839 VDD.n1145 VDD.n799 146.341
R2840 VDD.n1145 VDD.n765 146.341
R2841 VDD.n1151 VDD.n765 146.341
R2842 VDD.n1151 VDD.n757 146.341
R2843 VDD.n1161 VDD.n757 146.341
R2844 VDD.n1161 VDD.n753 146.341
R2845 VDD.n1167 VDD.n753 146.341
R2846 VDD.n1167 VDD.n745 146.341
R2847 VDD.n1177 VDD.n745 146.341
R2848 VDD.n1177 VDD.n741 146.341
R2849 VDD.n1183 VDD.n741 146.341
R2850 VDD.n1183 VDD.n733 146.341
R2851 VDD.n1193 VDD.n733 146.341
R2852 VDD.n1193 VDD.n729 146.341
R2853 VDD.n1199 VDD.n729 146.341
R2854 VDD.n1199 VDD.n720 146.341
R2855 VDD.n1210 VDD.n720 146.341
R2856 VDD.n1210 VDD.n715 146.341
R2857 VDD.n1398 VDD.n715 146.341
R2858 VDD.n969 VDD.t79 139.282
R2859 VDD.n1002 VDD.t92 139.282
R2860 VDD.n1035 VDD.t42 139.282
R2861 VDD.n705 VDD.t45 139.282
R2862 VDD.n1277 VDD.t56 139.282
R2863 VDD.n1242 VDD.t100 139.282
R2864 VDD.n199 VDD.t64 139.282
R2865 VDD.n166 VDD.t75 139.282
R2866 VDD.n131 VDD.t107 139.282
R2867 VDD.n341 VDD.t114 139.282
R2868 VDD.n2450 VDD.t85 139.282
R2869 VDD.n2367 VDD.t73 139.282
R2870 VDD.n970 VDD.t78 113.489
R2871 VDD.n1003 VDD.t91 113.489
R2872 VDD.n1036 VDD.t41 113.489
R2873 VDD.n706 VDD.t46 113.489
R2874 VDD.n1278 VDD.t57 113.489
R2875 VDD.n1243 VDD.t101 113.489
R2876 VDD.n200 VDD.t65 113.489
R2877 VDD.n167 VDD.t76 113.489
R2878 VDD.n132 VDD.t108 113.489
R2879 VDD.n342 VDD.t113 113.489
R2880 VDD.n2451 VDD.t84 113.489
R2881 VDD.n2368 VDD.t72 113.489
R2882 VDD.n9 VDD.n7 109.74
R2883 VDD.n2 VDD.n0 109.74
R2884 VDD.n9 VDD.n8 109.166
R2885 VDD.n11 VDD.n10 109.166
R2886 VDD.n13 VDD.n12 109.166
R2887 VDD.n6 VDD.n5 109.166
R2888 VDD.n4 VDD.n3 109.166
R2889 VDD.n2 VDD.n1 109.166
R2890 VDD.n2127 VDD.n507 99.5127
R2891 VDD.n2131 VDD.n507 99.5127
R2892 VDD.n2131 VDD.n497 99.5127
R2893 VDD.n2139 VDD.n497 99.5127
R2894 VDD.n2139 VDD.n495 99.5127
R2895 VDD.n2143 VDD.n495 99.5127
R2896 VDD.n2143 VDD.n485 99.5127
R2897 VDD.n2151 VDD.n485 99.5127
R2898 VDD.n2151 VDD.n483 99.5127
R2899 VDD.n2155 VDD.n483 99.5127
R2900 VDD.n2155 VDD.n474 99.5127
R2901 VDD.n2163 VDD.n474 99.5127
R2902 VDD.n2163 VDD.n472 99.5127
R2903 VDD.n2167 VDD.n472 99.5127
R2904 VDD.n2167 VDD.n463 99.5127
R2905 VDD.n2175 VDD.n463 99.5127
R2906 VDD.n2175 VDD.n461 99.5127
R2907 VDD.n2179 VDD.n461 99.5127
R2908 VDD.n2179 VDD.n451 99.5127
R2909 VDD.n2187 VDD.n451 99.5127
R2910 VDD.n2187 VDD.n449 99.5127
R2911 VDD.n2191 VDD.n449 99.5127
R2912 VDD.n2191 VDD.n439 99.5127
R2913 VDD.n2199 VDD.n439 99.5127
R2914 VDD.n2199 VDD.n437 99.5127
R2915 VDD.n2203 VDD.n437 99.5127
R2916 VDD.n2203 VDD.n427 99.5127
R2917 VDD.n2211 VDD.n427 99.5127
R2918 VDD.n2211 VDD.n425 99.5127
R2919 VDD.n2215 VDD.n425 99.5127
R2920 VDD.n2215 VDD.n416 99.5127
R2921 VDD.n2223 VDD.n416 99.5127
R2922 VDD.n2223 VDD.n414 99.5127
R2923 VDD.n2227 VDD.n414 99.5127
R2924 VDD.n2227 VDD.n402 99.5127
R2925 VDD.n2272 VDD.n402 99.5127
R2926 VDD.n2272 VDD.n400 99.5127
R2927 VDD.n2276 VDD.n400 99.5127
R2928 VDD.n2276 VDD.n373 99.5127
R2929 VDD.n2331 VDD.n373 99.5127
R2930 VDD.n2327 VDD.n2326 99.5127
R2931 VDD.n2324 VDD.n378 99.5127
R2932 VDD.n2320 VDD.n2319 99.5127
R2933 VDD.n2317 VDD.n381 99.5127
R2934 VDD.n2313 VDD.n2312 99.5127
R2935 VDD.n2310 VDD.n2307 99.5127
R2936 VDD.n2305 VDD.n384 99.5127
R2937 VDD.n2301 VDD.n2300 99.5127
R2938 VDD.n2298 VDD.n387 99.5127
R2939 VDD.n2294 VDD.n2293 99.5127
R2940 VDD.n2291 VDD.n390 99.5127
R2941 VDD.n2286 VDD.n2285 99.5127
R2942 VDD.n1957 VDD.n1871 99.5127
R2943 VDD.n1957 VDD.n504 99.5127
R2944 VDD.n1960 VDD.n504 99.5127
R2945 VDD.n1960 VDD.n498 99.5127
R2946 VDD.n1963 VDD.n498 99.5127
R2947 VDD.n1963 VDD.n493 99.5127
R2948 VDD.n1966 VDD.n493 99.5127
R2949 VDD.n1966 VDD.n487 99.5127
R2950 VDD.n1969 VDD.n487 99.5127
R2951 VDD.n1969 VDD.n481 99.5127
R2952 VDD.n1972 VDD.n481 99.5127
R2953 VDD.n1972 VDD.n476 99.5127
R2954 VDD.n1975 VDD.n476 99.5127
R2955 VDD.n1975 VDD.n470 99.5127
R2956 VDD.n2046 VDD.n470 99.5127
R2957 VDD.n2046 VDD.n464 99.5127
R2958 VDD.n2042 VDD.n464 99.5127
R2959 VDD.n2042 VDD.n459 99.5127
R2960 VDD.n2039 VDD.n459 99.5127
R2961 VDD.n2039 VDD.n452 99.5127
R2962 VDD.n2001 VDD.n452 99.5127
R2963 VDD.n2001 VDD.n446 99.5127
R2964 VDD.n1998 VDD.n446 99.5127
R2965 VDD.n1998 VDD.n440 99.5127
R2966 VDD.n1995 VDD.n440 99.5127
R2967 VDD.n1995 VDD.n434 99.5127
R2968 VDD.n1992 VDD.n434 99.5127
R2969 VDD.n1992 VDD.n428 99.5127
R2970 VDD.n1989 VDD.n428 99.5127
R2971 VDD.n1989 VDD.n423 99.5127
R2972 VDD.n1986 VDD.n423 99.5127
R2973 VDD.n1986 VDD.n418 99.5127
R2974 VDD.n1983 VDD.n418 99.5127
R2975 VDD.n1983 VDD.n412 99.5127
R2976 VDD.n1980 VDD.n412 99.5127
R2977 VDD.n1980 VDD.n404 99.5127
R2978 VDD.n404 VDD.n396 99.5127
R2979 VDD.n2278 VDD.n396 99.5127
R2980 VDD.n2279 VDD.n2278 99.5127
R2981 VDD.n2279 VDD.n371 99.5127
R2982 VDD.n1906 VDD.n1904 99.5127
R2983 VDD.n1910 VDD.n1904 99.5127
R2984 VDD.n1914 VDD.n1912 99.5127
R2985 VDD.n1918 VDD.n1902 99.5127
R2986 VDD.n1922 VDD.n1920 99.5127
R2987 VDD.n1926 VDD.n1900 99.5127
R2988 VDD.n1930 VDD.n1928 99.5127
R2989 VDD.n1934 VDD.n1898 99.5127
R2990 VDD.n1938 VDD.n1936 99.5127
R2991 VDD.n1942 VDD.n1896 99.5127
R2992 VDD.n1946 VDD.n1944 99.5127
R2993 VDD.n1951 VDD.n1892 99.5127
R2994 VDD.n1954 VDD.n1953 99.5127
R2995 VDD.n1808 VDD.n1807 99.5127
R2996 VDD.n1804 VDD.n1803 99.5127
R2997 VDD.n1800 VDD.n1799 99.5127
R2998 VDD.n1796 VDD.n1795 99.5127
R2999 VDD.n1792 VDD.n1791 99.5127
R3000 VDD.n1788 VDD.n1787 99.5127
R3001 VDD.n1784 VDD.n1783 99.5127
R3002 VDD.n1780 VDD.n1779 99.5127
R3003 VDD.n1776 VDD.n1775 99.5127
R3004 VDD.n1772 VDD.n1771 99.5127
R3005 VDD.n1768 VDD.n1767 99.5127
R3006 VDD.n1763 VDD.n1762 99.5127
R3007 VDD.n1580 VDD.n667 99.5127
R3008 VDD.n1580 VDD.n660 99.5127
R3009 VDD.n1577 VDD.n660 99.5127
R3010 VDD.n1577 VDD.n653 99.5127
R3011 VDD.n1574 VDD.n653 99.5127
R3012 VDD.n1574 VDD.n647 99.5127
R3013 VDD.n1571 VDD.n647 99.5127
R3014 VDD.n1571 VDD.n642 99.5127
R3015 VDD.n1568 VDD.n642 99.5127
R3016 VDD.n1568 VDD.n636 99.5127
R3017 VDD.n1565 VDD.n636 99.5127
R3018 VDD.n1565 VDD.n630 99.5127
R3019 VDD.n1562 VDD.n630 99.5127
R3020 VDD.n1562 VDD.n624 99.5127
R3021 VDD.n1559 VDD.n624 99.5127
R3022 VDD.n1559 VDD.n618 99.5127
R3023 VDD.n1556 VDD.n618 99.5127
R3024 VDD.n1556 VDD.n612 99.5127
R3025 VDD.n1553 VDD.n612 99.5127
R3026 VDD.n1553 VDD.n606 99.5127
R3027 VDD.n1550 VDD.n606 99.5127
R3028 VDD.n1550 VDD.n600 99.5127
R3029 VDD.n1519 VDD.n600 99.5127
R3030 VDD.n1519 VDD.n595 99.5127
R3031 VDD.n1539 VDD.n595 99.5127
R3032 VDD.n1539 VDD.n589 99.5127
R3033 VDD.n1535 VDD.n589 99.5127
R3034 VDD.n1535 VDD.n583 99.5127
R3035 VDD.n1532 VDD.n583 99.5127
R3036 VDD.n1532 VDD.n577 99.5127
R3037 VDD.n1529 VDD.n577 99.5127
R3038 VDD.n1529 VDD.n572 99.5127
R3039 VDD.n1526 VDD.n572 99.5127
R3040 VDD.n1526 VDD.n566 99.5127
R3041 VDD.n1523 VDD.n566 99.5127
R3042 VDD.n1523 VDD.n559 99.5127
R3043 VDD.n559 VDD.n553 99.5127
R3044 VDD.n1754 VDD.n553 99.5127
R3045 VDD.n1754 VDD.n545 99.5127
R3046 VDD.n1758 VDD.n545 99.5127
R3047 VDD.n1631 VDD.n1629 99.5127
R3048 VDD.n1629 VDD.n1628 99.5127
R3049 VDD.n1625 VDD.n1624 99.5127
R3050 VDD.n1622 VDD.n673 99.5127
R3051 VDD.n1618 VDD.n1616 99.5127
R3052 VDD.n1614 VDD.n675 99.5127
R3053 VDD.n1610 VDD.n1608 99.5127
R3054 VDD.n1605 VDD.n1604 99.5127
R3055 VDD.n1602 VDD.n679 99.5127
R3056 VDD.n1598 VDD.n1596 99.5127
R3057 VDD.n1594 VDD.n681 99.5127
R3058 VDD.n1590 VDD.n1588 99.5127
R3059 VDD.n1585 VDD.n1584 99.5127
R3060 VDD.n1635 VDD.n658 99.5127
R3061 VDD.n1643 VDD.n658 99.5127
R3062 VDD.n1643 VDD.n656 99.5127
R3063 VDD.n1647 VDD.n656 99.5127
R3064 VDD.n1647 VDD.n646 99.5127
R3065 VDD.n1656 VDD.n646 99.5127
R3066 VDD.n1656 VDD.n644 99.5127
R3067 VDD.n1660 VDD.n644 99.5127
R3068 VDD.n1660 VDD.n634 99.5127
R3069 VDD.n1668 VDD.n634 99.5127
R3070 VDD.n1668 VDD.n632 99.5127
R3071 VDD.n1672 VDD.n632 99.5127
R3072 VDD.n1672 VDD.n622 99.5127
R3073 VDD.n1680 VDD.n622 99.5127
R3074 VDD.n1680 VDD.n620 99.5127
R3075 VDD.n1684 VDD.n620 99.5127
R3076 VDD.n1684 VDD.n610 99.5127
R3077 VDD.n1692 VDD.n610 99.5127
R3078 VDD.n1692 VDD.n608 99.5127
R3079 VDD.n1696 VDD.n608 99.5127
R3080 VDD.n1696 VDD.n599 99.5127
R3081 VDD.n1704 VDD.n599 99.5127
R3082 VDD.n1704 VDD.n597 99.5127
R3083 VDD.n1708 VDD.n597 99.5127
R3084 VDD.n1708 VDD.n588 99.5127
R3085 VDD.n1716 VDD.n588 99.5127
R3086 VDD.n1716 VDD.n586 99.5127
R3087 VDD.n1720 VDD.n586 99.5127
R3088 VDD.n1720 VDD.n576 99.5127
R3089 VDD.n1728 VDD.n576 99.5127
R3090 VDD.n1728 VDD.n574 99.5127
R3091 VDD.n1732 VDD.n574 99.5127
R3092 VDD.n1732 VDD.n564 99.5127
R3093 VDD.n1740 VDD.n564 99.5127
R3094 VDD.n1740 VDD.n561 99.5127
R3095 VDD.n1745 VDD.n561 99.5127
R3096 VDD.n1745 VDD.n562 99.5127
R3097 VDD.n562 VDD.n547 99.5127
R3098 VDD.n1814 VDD.n547 99.5127
R3099 VDD.n1814 VDD.n548 99.5127
R3100 VDD.n2260 VDD.n2259 99.5127
R3101 VDD.n2257 VDD.n2235 99.5127
R3102 VDD.n2253 VDD.n2252 99.5127
R3103 VDD.n2250 VDD.n2238 99.5127
R3104 VDD.n2246 VDD.n2245 99.5127
R3105 VDD.n2243 VDD.n2241 99.5127
R3106 VDD.n2355 VDD.n2354 99.5127
R3107 VDD.n2352 VDD.n357 99.5127
R3108 VDD.n2348 VDD.n2347 99.5127
R3109 VDD.n2345 VDD.n360 99.5127
R3110 VDD.n2341 VDD.n2340 99.5127
R3111 VDD.n2338 VDD.n363 99.5127
R3112 VDD.n2069 VDD.n1872 99.5127
R3113 VDD.n2069 VDD.n505 99.5127
R3114 VDD.n2066 VDD.n505 99.5127
R3115 VDD.n2066 VDD.n499 99.5127
R3116 VDD.n2063 VDD.n499 99.5127
R3117 VDD.n2063 VDD.n494 99.5127
R3118 VDD.n2060 VDD.n494 99.5127
R3119 VDD.n2060 VDD.n488 99.5127
R3120 VDD.n2057 VDD.n488 99.5127
R3121 VDD.n2057 VDD.n482 99.5127
R3122 VDD.n2054 VDD.n482 99.5127
R3123 VDD.n2054 VDD.n477 99.5127
R3124 VDD.n2051 VDD.n477 99.5127
R3125 VDD.n2051 VDD.n471 99.5127
R3126 VDD.n2048 VDD.n471 99.5127
R3127 VDD.n2048 VDD.n465 99.5127
R3128 VDD.n2004 VDD.n465 99.5127
R3129 VDD.n2004 VDD.n460 99.5127
R3130 VDD.n2037 VDD.n460 99.5127
R3131 VDD.n2037 VDD.n453 99.5127
R3132 VDD.n2033 VDD.n453 99.5127
R3133 VDD.n2033 VDD.n447 99.5127
R3134 VDD.n2030 VDD.n447 99.5127
R3135 VDD.n2030 VDD.n441 99.5127
R3136 VDD.n2027 VDD.n441 99.5127
R3137 VDD.n2027 VDD.n435 99.5127
R3138 VDD.n2024 VDD.n435 99.5127
R3139 VDD.n2024 VDD.n429 99.5127
R3140 VDD.n2021 VDD.n429 99.5127
R3141 VDD.n2021 VDD.n424 99.5127
R3142 VDD.n2018 VDD.n424 99.5127
R3143 VDD.n2018 VDD.n419 99.5127
R3144 VDD.n2015 VDD.n419 99.5127
R3145 VDD.n2015 VDD.n413 99.5127
R3146 VDD.n2012 VDD.n413 99.5127
R3147 VDD.n2012 VDD.n405 99.5127
R3148 VDD.n2009 VDD.n405 99.5127
R3149 VDD.n2009 VDD.n398 99.5127
R3150 VDD.n398 VDD.n369 99.5127
R3151 VDD.n2333 VDD.n369 99.5127
R3152 VDD.n2121 VDD.n2119 99.5127
R3153 VDD.n2117 VDD.n1876 99.5127
R3154 VDD.n2113 VDD.n2111 99.5127
R3155 VDD.n2109 VDD.n1878 99.5127
R3156 VDD.n2105 VDD.n2103 99.5127
R3157 VDD.n2101 VDD.n1880 99.5127
R3158 VDD.n2097 VDD.n2095 99.5127
R3159 VDD.n2093 VDD.n1882 99.5127
R3160 VDD.n2089 VDD.n2087 99.5127
R3161 VDD.n2085 VDD.n1884 99.5127
R3162 VDD.n2081 VDD.n2079 99.5127
R3163 VDD.n2077 VDD.n1886 99.5127
R3164 VDD.n2125 VDD.n503 99.5127
R3165 VDD.n2133 VDD.n503 99.5127
R3166 VDD.n2133 VDD.n501 99.5127
R3167 VDD.n2137 VDD.n501 99.5127
R3168 VDD.n2137 VDD.n492 99.5127
R3169 VDD.n2145 VDD.n492 99.5127
R3170 VDD.n2145 VDD.n490 99.5127
R3171 VDD.n2149 VDD.n490 99.5127
R3172 VDD.n2149 VDD.n480 99.5127
R3173 VDD.n2157 VDD.n480 99.5127
R3174 VDD.n2157 VDD.n478 99.5127
R3175 VDD.n2161 VDD.n478 99.5127
R3176 VDD.n2161 VDD.n468 99.5127
R3177 VDD.n2169 VDD.n468 99.5127
R3178 VDD.n2169 VDD.n466 99.5127
R3179 VDD.n2173 VDD.n466 99.5127
R3180 VDD.n2173 VDD.n457 99.5127
R3181 VDD.n2181 VDD.n457 99.5127
R3182 VDD.n2181 VDD.n455 99.5127
R3183 VDD.n2185 VDD.n455 99.5127
R3184 VDD.n2185 VDD.n445 99.5127
R3185 VDD.n2193 VDD.n445 99.5127
R3186 VDD.n2193 VDD.n443 99.5127
R3187 VDD.n2197 VDD.n443 99.5127
R3188 VDD.n2197 VDD.n433 99.5127
R3189 VDD.n2205 VDD.n433 99.5127
R3190 VDD.n2205 VDD.n431 99.5127
R3191 VDD.n2209 VDD.n431 99.5127
R3192 VDD.n2209 VDD.n422 99.5127
R3193 VDD.n2217 VDD.n422 99.5127
R3194 VDD.n2217 VDD.n420 99.5127
R3195 VDD.n2221 VDD.n420 99.5127
R3196 VDD.n2221 VDD.n410 99.5127
R3197 VDD.n2229 VDD.n410 99.5127
R3198 VDD.n2229 VDD.n406 99.5127
R3199 VDD.n2270 VDD.n406 99.5127
R3200 VDD.n2270 VDD.n407 99.5127
R3201 VDD.n407 VDD.n399 99.5127
R3202 VDD.n2265 VDD.n399 99.5127
R3203 VDD.n2265 VDD.n372 99.5127
R3204 VDD.n1868 VDD.n538 99.5127
R3205 VDD.n1864 VDD.n1863 99.5127
R3206 VDD.n1860 VDD.n1859 99.5127
R3207 VDD.n1856 VDD.n1855 99.5127
R3208 VDD.n1852 VDD.n1851 99.5127
R3209 VDD.n1848 VDD.n1847 99.5127
R3210 VDD.n1844 VDD.n1843 99.5127
R3211 VDD.n1840 VDD.n1839 99.5127
R3212 VDD.n1836 VDD.n1835 99.5127
R3213 VDD.n1832 VDD.n1831 99.5127
R3214 VDD.n1828 VDD.n1827 99.5127
R3215 VDD.n1824 VDD.n1823 99.5127
R3216 VDD.n1820 VDD.n536 99.5127
R3217 VDD.n1470 VDD.n668 99.5127
R3218 VDD.n1470 VDD.n661 99.5127
R3219 VDD.n1473 VDD.n661 99.5127
R3220 VDD.n1473 VDD.n654 99.5127
R3221 VDD.n1476 VDD.n654 99.5127
R3222 VDD.n1476 VDD.n648 99.5127
R3223 VDD.n1479 VDD.n648 99.5127
R3224 VDD.n1479 VDD.n643 99.5127
R3225 VDD.n1482 VDD.n643 99.5127
R3226 VDD.n1482 VDD.n637 99.5127
R3227 VDD.n1485 VDD.n637 99.5127
R3228 VDD.n1485 VDD.n631 99.5127
R3229 VDD.n1488 VDD.n631 99.5127
R3230 VDD.n1488 VDD.n625 99.5127
R3231 VDD.n1491 VDD.n625 99.5127
R3232 VDD.n1491 VDD.n619 99.5127
R3233 VDD.n1494 VDD.n619 99.5127
R3234 VDD.n1494 VDD.n613 99.5127
R3235 VDD.n1497 VDD.n613 99.5127
R3236 VDD.n1497 VDD.n607 99.5127
R3237 VDD.n1548 VDD.n607 99.5127
R3238 VDD.n1548 VDD.n601 99.5127
R3239 VDD.n1544 VDD.n601 99.5127
R3240 VDD.n1544 VDD.n596 99.5127
R3241 VDD.n1541 VDD.n596 99.5127
R3242 VDD.n1541 VDD.n590 99.5127
R3243 VDD.n1516 VDD.n590 99.5127
R3244 VDD.n1516 VDD.n584 99.5127
R3245 VDD.n1513 VDD.n584 99.5127
R3246 VDD.n1513 VDD.n578 99.5127
R3247 VDD.n1510 VDD.n578 99.5127
R3248 VDD.n1510 VDD.n573 99.5127
R3249 VDD.n1507 VDD.n573 99.5127
R3250 VDD.n1507 VDD.n567 99.5127
R3251 VDD.n1504 VDD.n567 99.5127
R3252 VDD.n1504 VDD.n560 99.5127
R3253 VDD.n1501 VDD.n560 99.5127
R3254 VDD.n1501 VDD.n544 99.5127
R3255 VDD.n1816 VDD.n544 99.5127
R3256 VDD.n1817 VDD.n1816 99.5127
R3257 VDD.n1419 VDD.n665 99.5127
R3258 VDD.n1423 VDD.n1417 99.5127
R3259 VDD.n1427 VDD.n1425 99.5127
R3260 VDD.n1431 VDD.n1415 99.5127
R3261 VDD.n1435 VDD.n1433 99.5127
R3262 VDD.n1439 VDD.n1413 99.5127
R3263 VDD.n1443 VDD.n1441 99.5127
R3264 VDD.n1447 VDD.n694 99.5127
R3265 VDD.n1451 VDD.n1449 99.5127
R3266 VDD.n1455 VDD.n692 99.5127
R3267 VDD.n1459 VDD.n1457 99.5127
R3268 VDD.n1464 VDD.n688 99.5127
R3269 VDD.n1467 VDD.n1466 99.5127
R3270 VDD.n1637 VDD.n663 99.5127
R3271 VDD.n1641 VDD.n663 99.5127
R3272 VDD.n1641 VDD.n652 99.5127
R3273 VDD.n1649 VDD.n652 99.5127
R3274 VDD.n1649 VDD.n649 99.5127
R3275 VDD.n1654 VDD.n649 99.5127
R3276 VDD.n1654 VDD.n640 99.5127
R3277 VDD.n1662 VDD.n640 99.5127
R3278 VDD.n1662 VDD.n638 99.5127
R3279 VDD.n1666 VDD.n638 99.5127
R3280 VDD.n1666 VDD.n628 99.5127
R3281 VDD.n1674 VDD.n628 99.5127
R3282 VDD.n1674 VDD.n626 99.5127
R3283 VDD.n1678 VDD.n626 99.5127
R3284 VDD.n1678 VDD.n616 99.5127
R3285 VDD.n1686 VDD.n616 99.5127
R3286 VDD.n1686 VDD.n614 99.5127
R3287 VDD.n1690 VDD.n614 99.5127
R3288 VDD.n1690 VDD.n604 99.5127
R3289 VDD.n1698 VDD.n604 99.5127
R3290 VDD.n1698 VDD.n602 99.5127
R3291 VDD.n1702 VDD.n602 99.5127
R3292 VDD.n1702 VDD.n593 99.5127
R3293 VDD.n1710 VDD.n593 99.5127
R3294 VDD.n1710 VDD.n591 99.5127
R3295 VDD.n1714 VDD.n591 99.5127
R3296 VDD.n1714 VDD.n581 99.5127
R3297 VDD.n1722 VDD.n581 99.5127
R3298 VDD.n1722 VDD.n579 99.5127
R3299 VDD.n1726 VDD.n579 99.5127
R3300 VDD.n1726 VDD.n570 99.5127
R3301 VDD.n1734 VDD.n570 99.5127
R3302 VDD.n1734 VDD.n568 99.5127
R3303 VDD.n1738 VDD.n568 99.5127
R3304 VDD.n1738 VDD.n557 99.5127
R3305 VDD.n1747 VDD.n557 99.5127
R3306 VDD.n1747 VDD.n555 99.5127
R3307 VDD.n1752 VDD.n555 99.5127
R3308 VDD.n1752 VDD.n546 99.5127
R3309 VDD.n546 VDD.n537 99.5127
R3310 VDD.t5 VDD.t16 94.423
R3311 VDD.n36 VDD.t192 79.3769
R3312 VDD.n26 VDD.t167 79.3769
R3313 VDD.n17 VDD.t155 79.3769
R3314 VDD.n787 VDD.t147 79.3769
R3315 VDD.n777 VDD.t182 79.3769
R3316 VDD.n768 VDD.t126 79.3769
R3317 VDD.n43 VDD.t152 78.8036
R3318 VDD.n33 VDD.t184 78.8036
R3319 VDD.n24 VDD.t146 78.8036
R3320 VDD.n794 VDD.t174 78.8036
R3321 VDD.n784 VDD.t128 78.8036
R3322 VDD.n775 VDD.t194 78.8036
R3323 VDD.n2231 VDD.n408 78.546
R3324 VDD.n1652 VDD.n650 78.546
R3325 VDD.n42 VDD.n41 74.1601
R3326 VDD.n40 VDD.n39 74.1601
R3327 VDD.n38 VDD.n37 74.1601
R3328 VDD.n36 VDD.n35 74.1601
R3329 VDD.n32 VDD.n31 74.1601
R3330 VDD.n30 VDD.n29 74.1601
R3331 VDD.n28 VDD.n27 74.1601
R3332 VDD.n26 VDD.n25 74.1601
R3333 VDD.n23 VDD.n22 74.1601
R3334 VDD.n21 VDD.n20 74.1601
R3335 VDD.n19 VDD.n18 74.1601
R3336 VDD.n17 VDD.n16 74.1601
R3337 VDD.n787 VDD.n786 74.1601
R3338 VDD.n789 VDD.n788 74.1601
R3339 VDD.n791 VDD.n790 74.1601
R3340 VDD.n793 VDD.n792 74.1601
R3341 VDD.n777 VDD.n776 74.1601
R3342 VDD.n779 VDD.n778 74.1601
R3343 VDD.n781 VDD.n780 74.1601
R3344 VDD.n783 VDD.n782 74.1601
R3345 VDD.n768 VDD.n767 74.1601
R3346 VDD.n770 VDD.n769 74.1601
R3347 VDD.n772 VDD.n771 74.1601
R3348 VDD.n774 VDD.n773 74.1601
R3349 VDD.n2120 VDD.n1870 72.8958
R3350 VDD.n2118 VDD.n1870 72.8958
R3351 VDD.n2112 VDD.n1870 72.8958
R3352 VDD.n2110 VDD.n1870 72.8958
R3353 VDD.n2104 VDD.n1870 72.8958
R3354 VDD.n2102 VDD.n1870 72.8958
R3355 VDD.n2096 VDD.n1870 72.8958
R3356 VDD.n2094 VDD.n1870 72.8958
R3357 VDD.n2088 VDD.n1870 72.8958
R3358 VDD.n2086 VDD.n1870 72.8958
R3359 VDD.n2080 VDD.n1870 72.8958
R3360 VDD.n2078 VDD.n1870 72.8958
R3361 VDD.n2072 VDD.n1870 72.8958
R3362 VDD.n368 VDD.n275 72.8958
R3363 VDD.n2339 VDD.n275 72.8958
R3364 VDD.n362 VDD.n275 72.8958
R3365 VDD.n2346 VDD.n275 72.8958
R3366 VDD.n359 VDD.n275 72.8958
R3367 VDD.n2353 VDD.n275 72.8958
R3368 VDD.n356 VDD.n275 72.8958
R3369 VDD.n2244 VDD.n275 72.8958
R3370 VDD.n2240 VDD.n275 72.8958
R3371 VDD.n2251 VDD.n275 72.8958
R3372 VDD.n2237 VDD.n275 72.8958
R3373 VDD.n2258 VDD.n275 72.8958
R3374 VDD.n2261 VDD.n275 72.8958
R3375 VDD.n1630 VDD.n666 72.8958
R3376 VDD.n671 VDD.n666 72.8958
R3377 VDD.n1623 VDD.n666 72.8958
R3378 VDD.n1617 VDD.n666 72.8958
R3379 VDD.n1615 VDD.n666 72.8958
R3380 VDD.n1609 VDD.n666 72.8958
R3381 VDD.n677 VDD.n666 72.8958
R3382 VDD.n1603 VDD.n666 72.8958
R3383 VDD.n1597 VDD.n666 72.8958
R3384 VDD.n1595 VDD.n666 72.8958
R3385 VDD.n1589 VDD.n666 72.8958
R3386 VDD.n685 VDD.n666 72.8958
R3387 VDD.n1869 VDD.n523 72.8958
R3388 VDD.n1869 VDD.n522 72.8958
R3389 VDD.n1869 VDD.n521 72.8958
R3390 VDD.n1869 VDD.n520 72.8958
R3391 VDD.n1869 VDD.n519 72.8958
R3392 VDD.n1869 VDD.n518 72.8958
R3393 VDD.n1869 VDD.n517 72.8958
R3394 VDD.n1869 VDD.n516 72.8958
R3395 VDD.n1869 VDD.n515 72.8958
R3396 VDD.n1869 VDD.n514 72.8958
R3397 VDD.n1869 VDD.n513 72.8958
R3398 VDD.n1869 VDD.n512 72.8958
R3399 VDD.n1869 VDD.n511 72.8958
R3400 VDD.n1905 VDD.n1870 72.8958
R3401 VDD.n1911 VDD.n1870 72.8958
R3402 VDD.n1913 VDD.n1870 72.8958
R3403 VDD.n1919 VDD.n1870 72.8958
R3404 VDD.n1921 VDD.n1870 72.8958
R3405 VDD.n1927 VDD.n1870 72.8958
R3406 VDD.n1929 VDD.n1870 72.8958
R3407 VDD.n1935 VDD.n1870 72.8958
R3408 VDD.n1937 VDD.n1870 72.8958
R3409 VDD.n1943 VDD.n1870 72.8958
R3410 VDD.n1945 VDD.n1870 72.8958
R3411 VDD.n1952 VDD.n1870 72.8958
R3412 VDD.n2284 VDD.n275 72.8958
R3413 VDD.n394 VDD.n275 72.8958
R3414 VDD.n2292 VDD.n275 72.8958
R3415 VDD.n389 VDD.n275 72.8958
R3416 VDD.n2299 VDD.n275 72.8958
R3417 VDD.n386 VDD.n275 72.8958
R3418 VDD.n2306 VDD.n275 72.8958
R3419 VDD.n2311 VDD.n275 72.8958
R3420 VDD.n383 VDD.n275 72.8958
R3421 VDD.n2318 VDD.n275 72.8958
R3422 VDD.n380 VDD.n275 72.8958
R3423 VDD.n2325 VDD.n275 72.8958
R3424 VDD.n377 VDD.n275 72.8958
R3425 VDD.n1869 VDD.n535 72.8958
R3426 VDD.n1869 VDD.n534 72.8958
R3427 VDD.n1869 VDD.n533 72.8958
R3428 VDD.n1869 VDD.n532 72.8958
R3429 VDD.n1869 VDD.n531 72.8958
R3430 VDD.n1869 VDD.n530 72.8958
R3431 VDD.n1869 VDD.n529 72.8958
R3432 VDD.n1869 VDD.n528 72.8958
R3433 VDD.n1869 VDD.n527 72.8958
R3434 VDD.n1869 VDD.n526 72.8958
R3435 VDD.n1869 VDD.n525 72.8958
R3436 VDD.n1869 VDD.n524 72.8958
R3437 VDD.n1418 VDD.n666 72.8958
R3438 VDD.n1424 VDD.n666 72.8958
R3439 VDD.n1426 VDD.n666 72.8958
R3440 VDD.n1432 VDD.n666 72.8958
R3441 VDD.n1434 VDD.n666 72.8958
R3442 VDD.n1440 VDD.n666 72.8958
R3443 VDD.n1442 VDD.n666 72.8958
R3444 VDD.n1448 VDD.n666 72.8958
R3445 VDD.n1450 VDD.n666 72.8958
R3446 VDD.n1456 VDD.n666 72.8958
R3447 VDD.n1458 VDD.n666 72.8958
R3448 VDD.n1465 VDD.n666 72.8958
R3449 VDD.n1063 VDD.n1062 66.2847
R3450 VDD.n1062 VDD.n860 66.2847
R3451 VDD.n1062 VDD.n861 66.2847
R3452 VDD.n1062 VDD.n862 66.2847
R3453 VDD.n1062 VDD.n863 66.2847
R3454 VDD.n1062 VDD.n864 66.2847
R3455 VDD.n1062 VDD.n865 66.2847
R3456 VDD.n1062 VDD.n866 66.2847
R3457 VDD.n1062 VDD.n867 66.2847
R3458 VDD.n1062 VDD.n868 66.2847
R3459 VDD.n1062 VDD.n869 66.2847
R3460 VDD.n1062 VDD.n870 66.2847
R3461 VDD.n1062 VDD.n871 66.2847
R3462 VDD.n1062 VDD.n872 66.2847
R3463 VDD.n1062 VDD.n873 66.2847
R3464 VDD.n1062 VDD.n874 66.2847
R3465 VDD.n1062 VDD.n875 66.2847
R3466 VDD.n1062 VDD.n876 66.2847
R3467 VDD.n1062 VDD.n877 66.2847
R3468 VDD.n1062 VDD.n878 66.2847
R3469 VDD.n1062 VDD.n879 66.2847
R3470 VDD.n1062 VDD.n880 66.2847
R3471 VDD.n1062 VDD.n881 66.2847
R3472 VDD.n1062 VDD.n882 66.2847
R3473 VDD.n1062 VDD.n883 66.2847
R3474 VDD.n1062 VDD.n884 66.2847
R3475 VDD.n1062 VDD.n885 66.2847
R3476 VDD.n1062 VDD.n886 66.2847
R3477 VDD.n714 VDD.n709 66.2847
R3478 VDD.n714 VDD.n713 66.2847
R3479 VDD.n1297 VDD.n714 66.2847
R3480 VDD.n1301 VDD.n714 66.2847
R3481 VDD.n1305 VDD.n714 66.2847
R3482 VDD.n1295 VDD.n714 66.2847
R3483 VDD.n1312 VDD.n714 66.2847
R3484 VDD.n1288 VDD.n714 66.2847
R3485 VDD.n1319 VDD.n714 66.2847
R3486 VDD.n1282 VDD.n714 66.2847
R3487 VDD.n1328 VDD.n714 66.2847
R3488 VDD.n1274 VDD.n714 66.2847
R3489 VDD.n1335 VDD.n714 66.2847
R3490 VDD.n1267 VDD.n714 66.2847
R3491 VDD.n1342 VDD.n714 66.2847
R3492 VDD.n1260 VDD.n714 66.2847
R3493 VDD.n1349 VDD.n714 66.2847
R3494 VDD.n1253 VDD.n714 66.2847
R3495 VDD.n1356 VDD.n714 66.2847
R3496 VDD.n1247 VDD.n714 66.2847
R3497 VDD.n1365 VDD.n714 66.2847
R3498 VDD.n1239 VDD.n714 66.2847
R3499 VDD.n1372 VDD.n714 66.2847
R3500 VDD.n1232 VDD.n714 66.2847
R3501 VDD.n1379 VDD.n714 66.2847
R3502 VDD.n1227 VDD.n714 66.2847
R3503 VDD.n1221 VDD.n714 66.2847
R3504 VDD.n1390 VDD.n714 66.2847
R3505 VDD.n1216 VDD.n714 66.2847
R3506 VDD.n2482 VDD.n2481 66.2847
R3507 VDD.n2481 VDD.n276 66.2847
R3508 VDD.n2481 VDD.n277 66.2847
R3509 VDD.n2481 VDD.n278 66.2847
R3510 VDD.n2481 VDD.n279 66.2847
R3511 VDD.n2481 VDD.n280 66.2847
R3512 VDD.n2481 VDD.n281 66.2847
R3513 VDD.n2481 VDD.n282 66.2847
R3514 VDD.n2481 VDD.n283 66.2847
R3515 VDD.n2481 VDD.n284 66.2847
R3516 VDD.n2481 VDD.n285 66.2847
R3517 VDD.n2481 VDD.n286 66.2847
R3518 VDD.n2481 VDD.n287 66.2847
R3519 VDD.n2481 VDD.n288 66.2847
R3520 VDD.n2481 VDD.n289 66.2847
R3521 VDD.n2481 VDD.n290 66.2847
R3522 VDD.n2481 VDD.n291 66.2847
R3523 VDD.n2481 VDD.n292 66.2847
R3524 VDD.n2481 VDD.n293 66.2847
R3525 VDD.n2481 VDD.n294 66.2847
R3526 VDD.n2481 VDD.n295 66.2847
R3527 VDD.n2481 VDD.n296 66.2847
R3528 VDD.n2481 VDD.n297 66.2847
R3529 VDD.n2481 VDD.n298 66.2847
R3530 VDD.n2481 VDD.n299 66.2847
R3531 VDD.n2481 VDD.n300 66.2847
R3532 VDD.n2481 VDD.n301 66.2847
R3533 VDD.n2481 VDD.n302 66.2847
R3534 VDD.n2591 VDD.n98 66.2847
R3535 VDD.n198 VDD.n98 66.2847
R3536 VDD.n2598 VDD.n98 66.2847
R3537 VDD.n191 VDD.n98 66.2847
R3538 VDD.n2605 VDD.n98 66.2847
R3539 VDD.n184 VDD.n98 66.2847
R3540 VDD.n2612 VDD.n98 66.2847
R3541 VDD.n177 VDD.n98 66.2847
R3542 VDD.n2619 VDD.n98 66.2847
R3543 VDD.n171 VDD.n98 66.2847
R3544 VDD.n2628 VDD.n98 66.2847
R3545 VDD.n163 VDD.n98 66.2847
R3546 VDD.n2635 VDD.n98 66.2847
R3547 VDD.n156 VDD.n98 66.2847
R3548 VDD.n2642 VDD.n98 66.2847
R3549 VDD.n149 VDD.n98 66.2847
R3550 VDD.n2649 VDD.n98 66.2847
R3551 VDD.n142 VDD.n98 66.2847
R3552 VDD.n2656 VDD.n98 66.2847
R3553 VDD.n136 VDD.n98 66.2847
R3554 VDD.n2665 VDD.n98 66.2847
R3555 VDD.n128 VDD.n98 66.2847
R3556 VDD.n2672 VDD.n98 66.2847
R3557 VDD.n121 VDD.n98 66.2847
R3558 VDD.n2679 VDD.n98 66.2847
R3559 VDD.n114 VDD.n98 66.2847
R3560 VDD.n2686 VDD.n98 66.2847
R3561 VDD.n2689 VDD.n98 66.2847
R3562 VDD.n102 VDD.n98 66.2847
R3563 VDD.n103 VDD.n102 52.4337
R3564 VDD.n2689 VDD.n2688 52.4337
R3565 VDD.n2686 VDD.n2685 52.4337
R3566 VDD.n2681 VDD.n114 52.4337
R3567 VDD.n2679 VDD.n2678 52.4337
R3568 VDD.n2674 VDD.n121 52.4337
R3569 VDD.n2672 VDD.n2671 52.4337
R3570 VDD.n2667 VDD.n128 52.4337
R3571 VDD.n2665 VDD.n2664 52.4337
R3572 VDD.n2658 VDD.n136 52.4337
R3573 VDD.n2656 VDD.n2655 52.4337
R3574 VDD.n2651 VDD.n142 52.4337
R3575 VDD.n2649 VDD.n2648 52.4337
R3576 VDD.n2644 VDD.n149 52.4337
R3577 VDD.n2642 VDD.n2641 52.4337
R3578 VDD.n2637 VDD.n156 52.4337
R3579 VDD.n2635 VDD.n2634 52.4337
R3580 VDD.n2630 VDD.n163 52.4337
R3581 VDD.n2628 VDD.n2627 52.4337
R3582 VDD.n2621 VDD.n171 52.4337
R3583 VDD.n2619 VDD.n2618 52.4337
R3584 VDD.n2614 VDD.n177 52.4337
R3585 VDD.n2612 VDD.n2611 52.4337
R3586 VDD.n2607 VDD.n184 52.4337
R3587 VDD.n2605 VDD.n2604 52.4337
R3588 VDD.n2600 VDD.n191 52.4337
R3589 VDD.n2598 VDD.n2597 52.4337
R3590 VDD.n2593 VDD.n198 52.4337
R3591 VDD.n2591 VDD.n2590 52.4337
R3592 VDD.n2483 VDD.n2482 52.4337
R3593 VDD.n304 VDD.n276 52.4337
R3594 VDD.n2475 VDD.n277 52.4337
R3595 VDD.n312 VDD.n278 52.4337
R3596 VDD.n2468 VDD.n279 52.4337
R3597 VDD.n2465 VDD.n280 52.4337
R3598 VDD.n2461 VDD.n281 52.4337
R3599 VDD.n2457 VDD.n282 52.4337
R3600 VDD.n2453 VDD.n283 52.4337
R3601 VDD.n2445 VDD.n284 52.4337
R3602 VDD.n2441 VDD.n285 52.4337
R3603 VDD.n2437 VDD.n286 52.4337
R3604 VDD.n2433 VDD.n287 52.4337
R3605 VDD.n2429 VDD.n288 52.4337
R3606 VDD.n2425 VDD.n289 52.4337
R3607 VDD.n2421 VDD.n290 52.4337
R3608 VDD.n2417 VDD.n291 52.4337
R3609 VDD.n2413 VDD.n292 52.4337
R3610 VDD.n2409 VDD.n293 52.4337
R3611 VDD.n2403 VDD.n294 52.4337
R3612 VDD.n2399 VDD.n295 52.4337
R3613 VDD.n2395 VDD.n296 52.4337
R3614 VDD.n2391 VDD.n297 52.4337
R3615 VDD.n2387 VDD.n298 52.4337
R3616 VDD.n2383 VDD.n299 52.4337
R3617 VDD.n2359 VDD.n300 52.4337
R3618 VDD.n2376 VDD.n301 52.4337
R3619 VDD.n2373 VDD.n302 52.4337
R3620 VDD.n1392 VDD.n1216 52.4337
R3621 VDD.n1390 VDD.n1389 52.4337
R3622 VDD.n1222 VDD.n1221 52.4337
R3623 VDD.n1381 VDD.n1227 52.4337
R3624 VDD.n1379 VDD.n1378 52.4337
R3625 VDD.n1374 VDD.n1232 52.4337
R3626 VDD.n1372 VDD.n1371 52.4337
R3627 VDD.n1367 VDD.n1239 52.4337
R3628 VDD.n1365 VDD.n1364 52.4337
R3629 VDD.n1358 VDD.n1247 52.4337
R3630 VDD.n1356 VDD.n1355 52.4337
R3631 VDD.n1351 VDD.n1253 52.4337
R3632 VDD.n1349 VDD.n1348 52.4337
R3633 VDD.n1344 VDD.n1260 52.4337
R3634 VDD.n1342 VDD.n1341 52.4337
R3635 VDD.n1337 VDD.n1267 52.4337
R3636 VDD.n1335 VDD.n1334 52.4337
R3637 VDD.n1330 VDD.n1274 52.4337
R3638 VDD.n1328 VDD.n1327 52.4337
R3639 VDD.n1321 VDD.n1282 52.4337
R3640 VDD.n1319 VDD.n1318 52.4337
R3641 VDD.n1314 VDD.n1288 52.4337
R3642 VDD.n1312 VDD.n1311 52.4337
R3643 VDD.n1307 VDD.n1295 52.4337
R3644 VDD.n1305 VDD.n1304 52.4337
R3645 VDD.n1301 VDD.n1300 52.4337
R3646 VDD.n1297 VDD.n700 52.4337
R3647 VDD.n713 VDD.n702 52.4337
R3648 VDD.n1401 VDD.n709 52.4337
R3649 VDD.n1064 VDD.n1063 52.4337
R3650 VDD.n888 VDD.n860 52.4337
R3651 VDD.n892 VDD.n861 52.4337
R3652 VDD.n894 VDD.n862 52.4337
R3653 VDD.n898 VDD.n863 52.4337
R3654 VDD.n900 VDD.n864 52.4337
R3655 VDD.n904 VDD.n865 52.4337
R3656 VDD.n906 VDD.n866 52.4337
R3657 VDD.n1034 VDD.n867 52.4337
R3658 VDD.n911 VDD.n868 52.4337
R3659 VDD.n915 VDD.n869 52.4337
R3660 VDD.n917 VDD.n870 52.4337
R3661 VDD.n921 VDD.n871 52.4337
R3662 VDD.n923 VDD.n872 52.4337
R3663 VDD.n927 VDD.n873 52.4337
R3664 VDD.n929 VDD.n874 52.4337
R3665 VDD.n933 VDD.n875 52.4337
R3666 VDD.n935 VDD.n876 52.4337
R3667 VDD.n1001 VDD.n877 52.4337
R3668 VDD.n940 VDD.n878 52.4337
R3669 VDD.n944 VDD.n879 52.4337
R3670 VDD.n946 VDD.n880 52.4337
R3671 VDD.n950 VDD.n881 52.4337
R3672 VDD.n952 VDD.n882 52.4337
R3673 VDD.n956 VDD.n883 52.4337
R3674 VDD.n958 VDD.n884 52.4337
R3675 VDD.n962 VDD.n885 52.4337
R3676 VDD.n964 VDD.n886 52.4337
R3677 VDD.n1063 VDD.n859 52.4337
R3678 VDD.n891 VDD.n860 52.4337
R3679 VDD.n893 VDD.n861 52.4337
R3680 VDD.n897 VDD.n862 52.4337
R3681 VDD.n899 VDD.n863 52.4337
R3682 VDD.n903 VDD.n864 52.4337
R3683 VDD.n905 VDD.n865 52.4337
R3684 VDD.n909 VDD.n866 52.4337
R3685 VDD.n910 VDD.n867 52.4337
R3686 VDD.n914 VDD.n868 52.4337
R3687 VDD.n916 VDD.n869 52.4337
R3688 VDD.n920 VDD.n870 52.4337
R3689 VDD.n922 VDD.n871 52.4337
R3690 VDD.n926 VDD.n872 52.4337
R3691 VDD.n928 VDD.n873 52.4337
R3692 VDD.n932 VDD.n874 52.4337
R3693 VDD.n934 VDD.n875 52.4337
R3694 VDD.n938 VDD.n876 52.4337
R3695 VDD.n939 VDD.n877 52.4337
R3696 VDD.n943 VDD.n878 52.4337
R3697 VDD.n945 VDD.n879 52.4337
R3698 VDD.n949 VDD.n880 52.4337
R3699 VDD.n951 VDD.n881 52.4337
R3700 VDD.n955 VDD.n882 52.4337
R3701 VDD.n957 VDD.n883 52.4337
R3702 VDD.n961 VDD.n884 52.4337
R3703 VDD.n963 VDD.n885 52.4337
R3704 VDD.n967 VDD.n886 52.4337
R3705 VDD.n709 VDD.n708 52.4337
R3706 VDD.n713 VDD.n701 52.4337
R3707 VDD.n1298 VDD.n1297 52.4337
R3708 VDD.n1302 VDD.n1301 52.4337
R3709 VDD.n1306 VDD.n1305 52.4337
R3710 VDD.n1295 VDD.n1289 52.4337
R3711 VDD.n1313 VDD.n1312 52.4337
R3712 VDD.n1288 VDD.n1283 52.4337
R3713 VDD.n1320 VDD.n1319 52.4337
R3714 VDD.n1282 VDD.n1275 52.4337
R3715 VDD.n1329 VDD.n1328 52.4337
R3716 VDD.n1274 VDD.n1268 52.4337
R3717 VDD.n1336 VDD.n1335 52.4337
R3718 VDD.n1267 VDD.n1261 52.4337
R3719 VDD.n1343 VDD.n1342 52.4337
R3720 VDD.n1260 VDD.n1254 52.4337
R3721 VDD.n1350 VDD.n1349 52.4337
R3722 VDD.n1253 VDD.n1248 52.4337
R3723 VDD.n1357 VDD.n1356 52.4337
R3724 VDD.n1247 VDD.n1240 52.4337
R3725 VDD.n1366 VDD.n1365 52.4337
R3726 VDD.n1239 VDD.n1233 52.4337
R3727 VDD.n1373 VDD.n1372 52.4337
R3728 VDD.n1232 VDD.n1228 52.4337
R3729 VDD.n1380 VDD.n1379 52.4337
R3730 VDD.n1227 VDD.n1226 52.4337
R3731 VDD.n1221 VDD.n1217 52.4337
R3732 VDD.n1391 VDD.n1390 52.4337
R3733 VDD.n1216 VDD.n716 52.4337
R3734 VDD.n2482 VDD.n274 52.4337
R3735 VDD.n2476 VDD.n276 52.4337
R3736 VDD.n311 VDD.n277 52.4337
R3737 VDD.n314 VDD.n278 52.4337
R3738 VDD.n2466 VDD.n279 52.4337
R3739 VDD.n2462 VDD.n280 52.4337
R3740 VDD.n2458 VDD.n281 52.4337
R3741 VDD.n2454 VDD.n282 52.4337
R3742 VDD.n2444 VDD.n283 52.4337
R3743 VDD.n2442 VDD.n284 52.4337
R3744 VDD.n2438 VDD.n285 52.4337
R3745 VDD.n2434 VDD.n286 52.4337
R3746 VDD.n2430 VDD.n287 52.4337
R3747 VDD.n2426 VDD.n288 52.4337
R3748 VDD.n2422 VDD.n289 52.4337
R3749 VDD.n2418 VDD.n290 52.4337
R3750 VDD.n2414 VDD.n291 52.4337
R3751 VDD.n2410 VDD.n292 52.4337
R3752 VDD.n2402 VDD.n293 52.4337
R3753 VDD.n2400 VDD.n294 52.4337
R3754 VDD.n2396 VDD.n295 52.4337
R3755 VDD.n2392 VDD.n296 52.4337
R3756 VDD.n2388 VDD.n297 52.4337
R3757 VDD.n2384 VDD.n298 52.4337
R3758 VDD.n2358 VDD.n299 52.4337
R3759 VDD.n2361 VDD.n300 52.4337
R3760 VDD.n2374 VDD.n301 52.4337
R3761 VDD.n2370 VDD.n302 52.4337
R3762 VDD.n2592 VDD.n2591 52.4337
R3763 VDD.n198 VDD.n192 52.4337
R3764 VDD.n2599 VDD.n2598 52.4337
R3765 VDD.n191 VDD.n185 52.4337
R3766 VDD.n2606 VDD.n2605 52.4337
R3767 VDD.n184 VDD.n178 52.4337
R3768 VDD.n2613 VDD.n2612 52.4337
R3769 VDD.n177 VDD.n172 52.4337
R3770 VDD.n2620 VDD.n2619 52.4337
R3771 VDD.n171 VDD.n164 52.4337
R3772 VDD.n2629 VDD.n2628 52.4337
R3773 VDD.n163 VDD.n157 52.4337
R3774 VDD.n2636 VDD.n2635 52.4337
R3775 VDD.n156 VDD.n150 52.4337
R3776 VDD.n2643 VDD.n2642 52.4337
R3777 VDD.n149 VDD.n143 52.4337
R3778 VDD.n2650 VDD.n2649 52.4337
R3779 VDD.n142 VDD.n137 52.4337
R3780 VDD.n2657 VDD.n2656 52.4337
R3781 VDD.n136 VDD.n129 52.4337
R3782 VDD.n2666 VDD.n2665 52.4337
R3783 VDD.n128 VDD.n122 52.4337
R3784 VDD.n2673 VDD.n2672 52.4337
R3785 VDD.n121 VDD.n115 52.4337
R3786 VDD.n2680 VDD.n2679 52.4337
R3787 VDD.n114 VDD.n107 52.4337
R3788 VDD.n2687 VDD.n2686 52.4337
R3789 VDD.n2690 VDD.n2689 52.4337
R3790 VDD.n102 VDD.n99 52.4337
R3791 VDD.n2327 VDD.n377 39.2114
R3792 VDD.n2325 VDD.n2324 39.2114
R3793 VDD.n2320 VDD.n380 39.2114
R3794 VDD.n2318 VDD.n2317 39.2114
R3795 VDD.n2313 VDD.n383 39.2114
R3796 VDD.n2311 VDD.n2310 39.2114
R3797 VDD.n2306 VDD.n2305 39.2114
R3798 VDD.n2301 VDD.n386 39.2114
R3799 VDD.n2299 VDD.n2298 39.2114
R3800 VDD.n2294 VDD.n389 39.2114
R3801 VDD.n2292 VDD.n2291 39.2114
R3802 VDD.n2286 VDD.n394 39.2114
R3803 VDD.n2284 VDD.n2283 39.2114
R3804 VDD.n1905 VDD.n509 39.2114
R3805 VDD.n1911 VDD.n1910 39.2114
R3806 VDD.n1914 VDD.n1913 39.2114
R3807 VDD.n1919 VDD.n1918 39.2114
R3808 VDD.n1922 VDD.n1921 39.2114
R3809 VDD.n1927 VDD.n1926 39.2114
R3810 VDD.n1930 VDD.n1929 39.2114
R3811 VDD.n1935 VDD.n1934 39.2114
R3812 VDD.n1938 VDD.n1937 39.2114
R3813 VDD.n1943 VDD.n1942 39.2114
R3814 VDD.n1946 VDD.n1945 39.2114
R3815 VDD.n1952 VDD.n1951 39.2114
R3816 VDD.n1808 VDD.n511 39.2114
R3817 VDD.n1804 VDD.n512 39.2114
R3818 VDD.n1800 VDD.n513 39.2114
R3819 VDD.n1796 VDD.n514 39.2114
R3820 VDD.n1792 VDD.n515 39.2114
R3821 VDD.n1788 VDD.n516 39.2114
R3822 VDD.n1784 VDD.n517 39.2114
R3823 VDD.n1780 VDD.n518 39.2114
R3824 VDD.n1776 VDD.n519 39.2114
R3825 VDD.n1772 VDD.n520 39.2114
R3826 VDD.n1768 VDD.n521 39.2114
R3827 VDD.n1763 VDD.n522 39.2114
R3828 VDD.n1759 VDD.n523 39.2114
R3829 VDD.n1630 VDD.n669 39.2114
R3830 VDD.n1628 VDD.n671 39.2114
R3831 VDD.n1624 VDD.n1623 39.2114
R3832 VDD.n1617 VDD.n673 39.2114
R3833 VDD.n1616 VDD.n1615 39.2114
R3834 VDD.n1609 VDD.n675 39.2114
R3835 VDD.n1608 VDD.n677 39.2114
R3836 VDD.n1604 VDD.n1603 39.2114
R3837 VDD.n1597 VDD.n679 39.2114
R3838 VDD.n1596 VDD.n1595 39.2114
R3839 VDD.n1589 VDD.n681 39.2114
R3840 VDD.n1588 VDD.n685 39.2114
R3841 VDD.n2261 VDD.n2260 39.2114
R3842 VDD.n2258 VDD.n2257 39.2114
R3843 VDD.n2253 VDD.n2237 39.2114
R3844 VDD.n2251 VDD.n2250 39.2114
R3845 VDD.n2246 VDD.n2240 39.2114
R3846 VDD.n2244 VDD.n2243 39.2114
R3847 VDD.n2355 VDD.n356 39.2114
R3848 VDD.n2353 VDD.n2352 39.2114
R3849 VDD.n2348 VDD.n359 39.2114
R3850 VDD.n2346 VDD.n2345 39.2114
R3851 VDD.n2341 VDD.n362 39.2114
R3852 VDD.n2339 VDD.n2338 39.2114
R3853 VDD.n2334 VDD.n368 39.2114
R3854 VDD.n2120 VDD.n1874 39.2114
R3855 VDD.n2119 VDD.n2118 39.2114
R3856 VDD.n2112 VDD.n1876 39.2114
R3857 VDD.n2111 VDD.n2110 39.2114
R3858 VDD.n2104 VDD.n1878 39.2114
R3859 VDD.n2103 VDD.n2102 39.2114
R3860 VDD.n2096 VDD.n1880 39.2114
R3861 VDD.n2095 VDD.n2094 39.2114
R3862 VDD.n2088 VDD.n1882 39.2114
R3863 VDD.n2087 VDD.n2086 39.2114
R3864 VDD.n2080 VDD.n1884 39.2114
R3865 VDD.n2079 VDD.n2078 39.2114
R3866 VDD.n2072 VDD.n1886 39.2114
R3867 VDD.n2121 VDD.n2120 39.2114
R3868 VDD.n2118 VDD.n2117 39.2114
R3869 VDD.n2113 VDD.n2112 39.2114
R3870 VDD.n2110 VDD.n2109 39.2114
R3871 VDD.n2105 VDD.n2104 39.2114
R3872 VDD.n2102 VDD.n2101 39.2114
R3873 VDD.n2097 VDD.n2096 39.2114
R3874 VDD.n2094 VDD.n2093 39.2114
R3875 VDD.n2089 VDD.n2088 39.2114
R3876 VDD.n2086 VDD.n2085 39.2114
R3877 VDD.n2081 VDD.n2080 39.2114
R3878 VDD.n2078 VDD.n2077 39.2114
R3879 VDD.n2073 VDD.n2072 39.2114
R3880 VDD.n368 VDD.n363 39.2114
R3881 VDD.n2340 VDD.n2339 39.2114
R3882 VDD.n362 VDD.n360 39.2114
R3883 VDD.n2347 VDD.n2346 39.2114
R3884 VDD.n359 VDD.n357 39.2114
R3885 VDD.n2354 VDD.n2353 39.2114
R3886 VDD.n2241 VDD.n356 39.2114
R3887 VDD.n2245 VDD.n2244 39.2114
R3888 VDD.n2240 VDD.n2238 39.2114
R3889 VDD.n2252 VDD.n2251 39.2114
R3890 VDD.n2237 VDD.n2235 39.2114
R3891 VDD.n2259 VDD.n2258 39.2114
R3892 VDD.n2262 VDD.n2261 39.2114
R3893 VDD.n1631 VDD.n1630 39.2114
R3894 VDD.n1625 VDD.n671 39.2114
R3895 VDD.n1623 VDD.n1622 39.2114
R3896 VDD.n1618 VDD.n1617 39.2114
R3897 VDD.n1615 VDD.n1614 39.2114
R3898 VDD.n1610 VDD.n1609 39.2114
R3899 VDD.n1605 VDD.n677 39.2114
R3900 VDD.n1603 VDD.n1602 39.2114
R3901 VDD.n1598 VDD.n1597 39.2114
R3902 VDD.n1595 VDD.n1594 39.2114
R3903 VDD.n1590 VDD.n1589 39.2114
R3904 VDD.n1585 VDD.n685 39.2114
R3905 VDD.n1762 VDD.n523 39.2114
R3906 VDD.n1767 VDD.n522 39.2114
R3907 VDD.n1771 VDD.n521 39.2114
R3908 VDD.n1775 VDD.n520 39.2114
R3909 VDD.n1779 VDD.n519 39.2114
R3910 VDD.n1783 VDD.n518 39.2114
R3911 VDD.n1787 VDD.n517 39.2114
R3912 VDD.n1791 VDD.n516 39.2114
R3913 VDD.n1795 VDD.n515 39.2114
R3914 VDD.n1799 VDD.n514 39.2114
R3915 VDD.n1803 VDD.n513 39.2114
R3916 VDD.n1807 VDD.n512 39.2114
R3917 VDD.n1810 VDD.n511 39.2114
R3918 VDD.n1906 VDD.n1905 39.2114
R3919 VDD.n1912 VDD.n1911 39.2114
R3920 VDD.n1913 VDD.n1902 39.2114
R3921 VDD.n1920 VDD.n1919 39.2114
R3922 VDD.n1921 VDD.n1900 39.2114
R3923 VDD.n1928 VDD.n1927 39.2114
R3924 VDD.n1929 VDD.n1898 39.2114
R3925 VDD.n1936 VDD.n1935 39.2114
R3926 VDD.n1937 VDD.n1896 39.2114
R3927 VDD.n1944 VDD.n1943 39.2114
R3928 VDD.n1945 VDD.n1892 39.2114
R3929 VDD.n1953 VDD.n1952 39.2114
R3930 VDD.n2285 VDD.n2284 39.2114
R3931 VDD.n394 VDD.n390 39.2114
R3932 VDD.n2293 VDD.n2292 39.2114
R3933 VDD.n389 VDD.n387 39.2114
R3934 VDD.n2300 VDD.n2299 39.2114
R3935 VDD.n386 VDD.n384 39.2114
R3936 VDD.n2307 VDD.n2306 39.2114
R3937 VDD.n2312 VDD.n2311 39.2114
R3938 VDD.n383 VDD.n381 39.2114
R3939 VDD.n2319 VDD.n2318 39.2114
R3940 VDD.n380 VDD.n378 39.2114
R3941 VDD.n2326 VDD.n2325 39.2114
R3942 VDD.n377 VDD.n374 39.2114
R3943 VDD.n538 VDD.n524 39.2114
R3944 VDD.n1863 VDD.n525 39.2114
R3945 VDD.n1859 VDD.n526 39.2114
R3946 VDD.n1855 VDD.n527 39.2114
R3947 VDD.n1851 VDD.n528 39.2114
R3948 VDD.n1847 VDD.n529 39.2114
R3949 VDD.n1843 VDD.n530 39.2114
R3950 VDD.n1839 VDD.n531 39.2114
R3951 VDD.n1835 VDD.n532 39.2114
R3952 VDD.n1831 VDD.n533 39.2114
R3953 VDD.n1827 VDD.n534 39.2114
R3954 VDD.n1823 VDD.n535 39.2114
R3955 VDD.n1419 VDD.n1418 39.2114
R3956 VDD.n1424 VDD.n1423 39.2114
R3957 VDD.n1427 VDD.n1426 39.2114
R3958 VDD.n1432 VDD.n1431 39.2114
R3959 VDD.n1435 VDD.n1434 39.2114
R3960 VDD.n1440 VDD.n1439 39.2114
R3961 VDD.n1443 VDD.n1442 39.2114
R3962 VDD.n1448 VDD.n1447 39.2114
R3963 VDD.n1451 VDD.n1450 39.2114
R3964 VDD.n1456 VDD.n1455 39.2114
R3965 VDD.n1459 VDD.n1458 39.2114
R3966 VDD.n1465 VDD.n1464 39.2114
R3967 VDD.n1820 VDD.n535 39.2114
R3968 VDD.n1824 VDD.n534 39.2114
R3969 VDD.n1828 VDD.n533 39.2114
R3970 VDD.n1832 VDD.n532 39.2114
R3971 VDD.n1836 VDD.n531 39.2114
R3972 VDD.n1840 VDD.n530 39.2114
R3973 VDD.n1844 VDD.n529 39.2114
R3974 VDD.n1848 VDD.n528 39.2114
R3975 VDD.n1852 VDD.n527 39.2114
R3976 VDD.n1856 VDD.n526 39.2114
R3977 VDD.n1860 VDD.n525 39.2114
R3978 VDD.n1864 VDD.n524 39.2114
R3979 VDD.n1418 VDD.n1417 39.2114
R3980 VDD.n1425 VDD.n1424 39.2114
R3981 VDD.n1426 VDD.n1415 39.2114
R3982 VDD.n1433 VDD.n1432 39.2114
R3983 VDD.n1434 VDD.n1413 39.2114
R3984 VDD.n1441 VDD.n1440 39.2114
R3985 VDD.n1442 VDD.n694 39.2114
R3986 VDD.n1449 VDD.n1448 39.2114
R3987 VDD.n1450 VDD.n692 39.2114
R3988 VDD.n1457 VDD.n1456 39.2114
R3989 VDD.n1458 VDD.n688 39.2114
R3990 VDD.n1466 VDD.n1465 39.2114
R3991 VDD.n971 VDD.n970 37.4308
R3992 VDD.n1004 VDD.n1003 37.4308
R3993 VDD.n1037 VDD.n1036 37.4308
R3994 VDD.n707 VDD.n706 37.4308
R3995 VDD.n1326 VDD.n1278 37.4308
R3996 VDD.n1363 VDD.n1243 37.4308
R3997 VDD.n201 VDD.n200 37.4308
R3998 VDD.n2626 VDD.n167 37.4308
R3999 VDD.n2663 VDD.n132 37.4308
R4000 VDD.n2408 VDD.n342 37.4308
R4001 VDD.n2452 VDD.n2451 37.4308
R4002 VDD.n2369 VDD.n2368 37.4308
R4003 VDD.n1634 VDD.n1633 31.3761
R4004 VDD.n1812 VDD.n1811 31.3761
R4005 VDD.n1760 VDD.n1757 31.3761
R4006 VDD.n1583 VDD.n1582 31.3761
R4007 VDD.n1956 VDD.n1955 31.3761
R4008 VDD.n2282 VDD.n2281 31.3761
R4009 VDD.n2128 VDD.n508 31.3761
R4010 VDD.n2330 VDD.n2329 31.3761
R4011 VDD.n2264 VDD.n2263 31.3761
R4012 VDD.n2335 VDD.n367 31.3761
R4013 VDD.n2074 VDD.n2071 31.3761
R4014 VDD.n2124 VDD.n2123 31.3761
R4015 VDD.n1638 VDD.n664 31.3761
R4016 VDD.n1867 VDD.n539 31.3761
R4017 VDD.n1819 VDD.n1818 31.3761
R4018 VDD.n1469 VDD.n1468 31.3761
R4019 VDD.n1462 VDD.n690 30.449
R4020 VDD.n542 VDD.n541 30.449
R4021 VDD.n684 VDD.n683 30.449
R4022 VDD.n1765 VDD.n551 30.449
R4023 VDD.n1889 VDD.n1888 30.449
R4024 VDD.n2288 VDD.n392 30.449
R4025 VDD.n1949 VDD.n1894 30.449
R4026 VDD.n366 VDD.n365 30.449
R4027 VDD.n690 VDD.n689 25.7944
R4028 VDD.n541 VDD.n540 25.7944
R4029 VDD.n970 VDD.n969 25.7944
R4030 VDD.n1003 VDD.n1002 25.7944
R4031 VDD.n1036 VDD.n1035 25.7944
R4032 VDD.n706 VDD.n705 25.7944
R4033 VDD.n1278 VDD.n1277 25.7944
R4034 VDD.n1243 VDD.n1242 25.7944
R4035 VDD.n683 VDD.n682 25.7944
R4036 VDD.n551 VDD.n550 25.7944
R4037 VDD.n1888 VDD.n1887 25.7944
R4038 VDD.n200 VDD.n199 25.7944
R4039 VDD.n167 VDD.n166 25.7944
R4040 VDD.n132 VDD.n131 25.7944
R4041 VDD.n342 VDD.n341 25.7944
R4042 VDD.n2451 VDD.n2450 25.7944
R4043 VDD.n392 VDD.n391 25.7944
R4044 VDD.n1894 VDD.n1893 25.7944
R4045 VDD.n2368 VDD.n2367 25.7944
R4046 VDD.n365 VDD.n364 25.7944
R4047 VDD.n1062 VDD.n854 22.6677
R4048 VDD.n1399 VDD.n714 22.6677
R4049 VDD.n2481 VDD.n269 22.6677
R4050 VDD.n2698 VDD.n98 22.6677
R4051 VDD.n1073 VDD.n852 19.3944
R4052 VDD.n1073 VDD.n850 19.3944
R4053 VDD.n1077 VDD.n850 19.3944
R4054 VDD.n1077 VDD.n839 19.3944
R4055 VDD.n1089 VDD.n839 19.3944
R4056 VDD.n1089 VDD.n837 19.3944
R4057 VDD.n1093 VDD.n837 19.3944
R4058 VDD.n1093 VDD.n828 19.3944
R4059 VDD.n1105 VDD.n828 19.3944
R4060 VDD.n1105 VDD.n826 19.3944
R4061 VDD.n1109 VDD.n826 19.3944
R4062 VDD.n1109 VDD.n815 19.3944
R4063 VDD.n1121 VDD.n815 19.3944
R4064 VDD.n1121 VDD.n813 19.3944
R4065 VDD.n1125 VDD.n813 19.3944
R4066 VDD.n1125 VDD.n804 19.3944
R4067 VDD.n1138 VDD.n804 19.3944
R4068 VDD.n1138 VDD.n802 19.3944
R4069 VDD.n1142 VDD.n802 19.3944
R4070 VDD.n1142 VDD.n761 19.3944
R4071 VDD.n1154 VDD.n761 19.3944
R4072 VDD.n1154 VDD.n759 19.3944
R4073 VDD.n1158 VDD.n759 19.3944
R4074 VDD.n1158 VDD.n750 19.3944
R4075 VDD.n1170 VDD.n750 19.3944
R4076 VDD.n1170 VDD.n748 19.3944
R4077 VDD.n1174 VDD.n748 19.3944
R4078 VDD.n1174 VDD.n737 19.3944
R4079 VDD.n1186 VDD.n737 19.3944
R4080 VDD.n1186 VDD.n735 19.3944
R4081 VDD.n1190 VDD.n735 19.3944
R4082 VDD.n1190 VDD.n726 19.3944
R4083 VDD.n1202 VDD.n726 19.3944
R4084 VDD.n1202 VDD.n723 19.3944
R4085 VDD.n1207 VDD.n723 19.3944
R4086 VDD.n1207 VDD.n724 19.3944
R4087 VDD.n724 VDD.n711 19.3944
R4088 VDD.n1000 VDD.n941 19.3944
R4089 VDD.n996 VDD.n941 19.3944
R4090 VDD.n996 VDD.n995 19.3944
R4091 VDD.n995 VDD.n994 19.3944
R4092 VDD.n994 VDD.n947 19.3944
R4093 VDD.n990 VDD.n947 19.3944
R4094 VDD.n990 VDD.n989 19.3944
R4095 VDD.n989 VDD.n988 19.3944
R4096 VDD.n988 VDD.n953 19.3944
R4097 VDD.n984 VDD.n953 19.3944
R4098 VDD.n984 VDD.n983 19.3944
R4099 VDD.n983 VDD.n982 19.3944
R4100 VDD.n982 VDD.n959 19.3944
R4101 VDD.n978 VDD.n959 19.3944
R4102 VDD.n978 VDD.n977 19.3944
R4103 VDD.n977 VDD.n976 19.3944
R4104 VDD.n976 VDD.n965 19.3944
R4105 VDD.n972 VDD.n965 19.3944
R4106 VDD.n1033 VDD.n912 19.3944
R4107 VDD.n1029 VDD.n912 19.3944
R4108 VDD.n1029 VDD.n1028 19.3944
R4109 VDD.n1028 VDD.n1027 19.3944
R4110 VDD.n1027 VDD.n918 19.3944
R4111 VDD.n1023 VDD.n918 19.3944
R4112 VDD.n1023 VDD.n1022 19.3944
R4113 VDD.n1022 VDD.n1021 19.3944
R4114 VDD.n1021 VDD.n924 19.3944
R4115 VDD.n1017 VDD.n924 19.3944
R4116 VDD.n1017 VDD.n1016 19.3944
R4117 VDD.n1016 VDD.n1015 19.3944
R4118 VDD.n1015 VDD.n930 19.3944
R4119 VDD.n1011 VDD.n930 19.3944
R4120 VDD.n1011 VDD.n1010 19.3944
R4121 VDD.n1010 VDD.n1009 19.3944
R4122 VDD.n1009 VDD.n936 19.3944
R4123 VDD.n1005 VDD.n936 19.3944
R4124 VDD.n1065 VDD.n858 19.3944
R4125 VDD.n1060 VDD.n858 19.3944
R4126 VDD.n1060 VDD.n889 19.3944
R4127 VDD.n1056 VDD.n889 19.3944
R4128 VDD.n1056 VDD.n1055 19.3944
R4129 VDD.n1055 VDD.n1054 19.3944
R4130 VDD.n1054 VDD.n895 19.3944
R4131 VDD.n1050 VDD.n895 19.3944
R4132 VDD.n1050 VDD.n1049 19.3944
R4133 VDD.n1049 VDD.n1048 19.3944
R4134 VDD.n1048 VDD.n901 19.3944
R4135 VDD.n1044 VDD.n901 19.3944
R4136 VDD.n1044 VDD.n1043 19.3944
R4137 VDD.n1043 VDD.n1042 19.3944
R4138 VDD.n1042 VDD.n907 19.3944
R4139 VDD.n1038 VDD.n907 19.3944
R4140 VDD.n1322 VDD.n1276 19.3944
R4141 VDD.n1322 VDD.n1281 19.3944
R4142 VDD.n1317 VDD.n1281 19.3944
R4143 VDD.n1317 VDD.n1316 19.3944
R4144 VDD.n1316 VDD.n1315 19.3944
R4145 VDD.n1315 VDD.n1287 19.3944
R4146 VDD.n1310 VDD.n1287 19.3944
R4147 VDD.n1310 VDD.n1309 19.3944
R4148 VDD.n1309 VDD.n1308 19.3944
R4149 VDD.n1308 VDD.n1294 19.3944
R4150 VDD.n1303 VDD.n1294 19.3944
R4151 VDD.n1299 VDD.n1296 19.3944
R4152 VDD.n1408 VDD.n699 19.3944
R4153 VDD.n1408 VDD.n1407 19.3944
R4154 VDD.n1407 VDD.n1406 19.3944
R4155 VDD.n1406 VDD.n703 19.3944
R4156 VDD.n1359 VDD.n1241 19.3944
R4157 VDD.n1359 VDD.n1246 19.3944
R4158 VDD.n1354 VDD.n1246 19.3944
R4159 VDD.n1354 VDD.n1353 19.3944
R4160 VDD.n1353 VDD.n1352 19.3944
R4161 VDD.n1352 VDD.n1252 19.3944
R4162 VDD.n1347 VDD.n1252 19.3944
R4163 VDD.n1347 VDD.n1346 19.3944
R4164 VDD.n1346 VDD.n1345 19.3944
R4165 VDD.n1345 VDD.n1259 19.3944
R4166 VDD.n1340 VDD.n1259 19.3944
R4167 VDD.n1340 VDD.n1339 19.3944
R4168 VDD.n1339 VDD.n1338 19.3944
R4169 VDD.n1338 VDD.n1266 19.3944
R4170 VDD.n1333 VDD.n1266 19.3944
R4171 VDD.n1333 VDD.n1332 19.3944
R4172 VDD.n1332 VDD.n1331 19.3944
R4173 VDD.n1331 VDD.n1273 19.3944
R4174 VDD.n1394 VDD.n1393 19.3944
R4175 VDD.n1393 VDD.n1215 19.3944
R4176 VDD.n1388 VDD.n1215 19.3944
R4177 VDD.n1388 VDD.n1387 19.3944
R4178 VDD.n1387 VDD.n1386 19.3944
R4179 VDD.n1382 VDD.n1223 19.3944
R4180 VDD.n1377 VDD.n1225 19.3944
R4181 VDD.n1377 VDD.n1376 19.3944
R4182 VDD.n1376 VDD.n1375 19.3944
R4183 VDD.n1375 VDD.n1231 19.3944
R4184 VDD.n1370 VDD.n1231 19.3944
R4185 VDD.n1370 VDD.n1369 19.3944
R4186 VDD.n1369 VDD.n1368 19.3944
R4187 VDD.n1368 VDD.n1238 19.3944
R4188 VDD.n1069 VDD.n856 19.3944
R4189 VDD.n1069 VDD.n846 19.3944
R4190 VDD.n1081 VDD.n846 19.3944
R4191 VDD.n1081 VDD.n844 19.3944
R4192 VDD.n1085 VDD.n844 19.3944
R4193 VDD.n1085 VDD.n834 19.3944
R4194 VDD.n1097 VDD.n834 19.3944
R4195 VDD.n1097 VDD.n832 19.3944
R4196 VDD.n1101 VDD.n832 19.3944
R4197 VDD.n1101 VDD.n822 19.3944
R4198 VDD.n1113 VDD.n822 19.3944
R4199 VDD.n1113 VDD.n820 19.3944
R4200 VDD.n1117 VDD.n820 19.3944
R4201 VDD.n1117 VDD.n810 19.3944
R4202 VDD.n1129 VDD.n810 19.3944
R4203 VDD.n1129 VDD.n808 19.3944
R4204 VDD.n1134 VDD.n808 19.3944
R4205 VDD.n1134 VDD.n798 19.3944
R4206 VDD.n1146 VDD.n798 19.3944
R4207 VDD.n1146 VDD.n766 19.3944
R4208 VDD.n1150 VDD.n766 19.3944
R4209 VDD.n1150 VDD.n756 19.3944
R4210 VDD.n1162 VDD.n756 19.3944
R4211 VDD.n1162 VDD.n754 19.3944
R4212 VDD.n1166 VDD.n754 19.3944
R4213 VDD.n1166 VDD.n744 19.3944
R4214 VDD.n1178 VDD.n744 19.3944
R4215 VDD.n1178 VDD.n742 19.3944
R4216 VDD.n1182 VDD.n742 19.3944
R4217 VDD.n1182 VDD.n732 19.3944
R4218 VDD.n1194 VDD.n732 19.3944
R4219 VDD.n1194 VDD.n730 19.3944
R4220 VDD.n1198 VDD.n730 19.3944
R4221 VDD.n1198 VDD.n719 19.3944
R4222 VDD.n1211 VDD.n719 19.3944
R4223 VDD.n1211 VDD.n717 19.3944
R4224 VDD.n1397 VDD.n717 19.3944
R4225 VDD.n2492 VDD.n267 19.3944
R4226 VDD.n2492 VDD.n265 19.3944
R4227 VDD.n2496 VDD.n265 19.3944
R4228 VDD.n2496 VDD.n254 19.3944
R4229 VDD.n2508 VDD.n254 19.3944
R4230 VDD.n2508 VDD.n252 19.3944
R4231 VDD.n2512 VDD.n252 19.3944
R4232 VDD.n2512 VDD.n243 19.3944
R4233 VDD.n2524 VDD.n243 19.3944
R4234 VDD.n2524 VDD.n241 19.3944
R4235 VDD.n2528 VDD.n241 19.3944
R4236 VDD.n2528 VDD.n230 19.3944
R4237 VDD.n2540 VDD.n230 19.3944
R4238 VDD.n2540 VDD.n228 19.3944
R4239 VDD.n2544 VDD.n228 19.3944
R4240 VDD.n2544 VDD.n218 19.3944
R4241 VDD.n2556 VDD.n218 19.3944
R4242 VDD.n2556 VDD.n216 19.3944
R4243 VDD.n2560 VDD.n216 19.3944
R4244 VDD.n2561 VDD.n2560 19.3944
R4245 VDD.n2562 VDD.n2561 19.3944
R4246 VDD.n2562 VDD.n214 19.3944
R4247 VDD.n2566 VDD.n214 19.3944
R4248 VDD.n2567 VDD.n2566 19.3944
R4249 VDD.n2568 VDD.n2567 19.3944
R4250 VDD.n2568 VDD.n211 19.3944
R4251 VDD.n2572 VDD.n211 19.3944
R4252 VDD.n2573 VDD.n2572 19.3944
R4253 VDD.n2574 VDD.n2573 19.3944
R4254 VDD.n2574 VDD.n208 19.3944
R4255 VDD.n2578 VDD.n208 19.3944
R4256 VDD.n2579 VDD.n2578 19.3944
R4257 VDD.n2580 VDD.n2579 19.3944
R4258 VDD.n2580 VDD.n205 19.3944
R4259 VDD.n2584 VDD.n205 19.3944
R4260 VDD.n2585 VDD.n2584 19.3944
R4261 VDD.n2586 VDD.n2585 19.3944
R4262 VDD.n2622 VDD.n165 19.3944
R4263 VDD.n2622 VDD.n170 19.3944
R4264 VDD.n2617 VDD.n170 19.3944
R4265 VDD.n2617 VDD.n2616 19.3944
R4266 VDD.n2616 VDD.n2615 19.3944
R4267 VDD.n2615 VDD.n176 19.3944
R4268 VDD.n2610 VDD.n176 19.3944
R4269 VDD.n2610 VDD.n2609 19.3944
R4270 VDD.n2609 VDD.n2608 19.3944
R4271 VDD.n2608 VDD.n183 19.3944
R4272 VDD.n2603 VDD.n183 19.3944
R4273 VDD.n2603 VDD.n2602 19.3944
R4274 VDD.n2602 VDD.n2601 19.3944
R4275 VDD.n2601 VDD.n190 19.3944
R4276 VDD.n2596 VDD.n190 19.3944
R4277 VDD.n2596 VDD.n2595 19.3944
R4278 VDD.n2595 VDD.n2594 19.3944
R4279 VDD.n2594 VDD.n197 19.3944
R4280 VDD.n2659 VDD.n130 19.3944
R4281 VDD.n2659 VDD.n135 19.3944
R4282 VDD.n2654 VDD.n135 19.3944
R4283 VDD.n2654 VDD.n2653 19.3944
R4284 VDD.n2653 VDD.n2652 19.3944
R4285 VDD.n2652 VDD.n141 19.3944
R4286 VDD.n2647 VDD.n141 19.3944
R4287 VDD.n2647 VDD.n2646 19.3944
R4288 VDD.n2646 VDD.n2645 19.3944
R4289 VDD.n2645 VDD.n148 19.3944
R4290 VDD.n2640 VDD.n148 19.3944
R4291 VDD.n2640 VDD.n2639 19.3944
R4292 VDD.n2639 VDD.n2638 19.3944
R4293 VDD.n2638 VDD.n155 19.3944
R4294 VDD.n2633 VDD.n155 19.3944
R4295 VDD.n2633 VDD.n2632 19.3944
R4296 VDD.n2632 VDD.n2631 19.3944
R4297 VDD.n2631 VDD.n162 19.3944
R4298 VDD.n2693 VDD.n2692 19.3944
R4299 VDD.n2692 VDD.n2691 19.3944
R4300 VDD.n2691 VDD.n105 19.3944
R4301 VDD.n106 VDD.n105 19.3944
R4302 VDD.n2684 VDD.n106 19.3944
R4303 VDD.n2684 VDD.n2683 19.3944
R4304 VDD.n2683 VDD.n2682 19.3944
R4305 VDD.n2682 VDD.n113 19.3944
R4306 VDD.n2677 VDD.n113 19.3944
R4307 VDD.n2677 VDD.n2676 19.3944
R4308 VDD.n2676 VDD.n2675 19.3944
R4309 VDD.n2675 VDD.n120 19.3944
R4310 VDD.n2670 VDD.n120 19.3944
R4311 VDD.n2670 VDD.n2669 19.3944
R4312 VDD.n2669 VDD.n2668 19.3944
R4313 VDD.n2668 VDD.n127 19.3944
R4314 VDD.n2488 VDD.n271 19.3944
R4315 VDD.n2488 VDD.n261 19.3944
R4316 VDD.n2500 VDD.n261 19.3944
R4317 VDD.n2500 VDD.n259 19.3944
R4318 VDD.n2504 VDD.n259 19.3944
R4319 VDD.n2504 VDD.n249 19.3944
R4320 VDD.n2516 VDD.n249 19.3944
R4321 VDD.n2516 VDD.n247 19.3944
R4322 VDD.n2520 VDD.n247 19.3944
R4323 VDD.n2520 VDD.n237 19.3944
R4324 VDD.n2532 VDD.n237 19.3944
R4325 VDD.n2532 VDD.n235 19.3944
R4326 VDD.n2536 VDD.n235 19.3944
R4327 VDD.n2536 VDD.n225 19.3944
R4328 VDD.n2548 VDD.n225 19.3944
R4329 VDD.n2548 VDD.n223 19.3944
R4330 VDD.n2552 VDD.n223 19.3944
R4331 VDD.n2552 VDD.n47 19.3944
R4332 VDD.n2734 VDD.n47 19.3944
R4333 VDD.n2734 VDD.n48 19.3944
R4334 VDD.n2728 VDD.n48 19.3944
R4335 VDD.n2728 VDD.n2727 19.3944
R4336 VDD.n2727 VDD.n2726 19.3944
R4337 VDD.n2726 VDD.n60 19.3944
R4338 VDD.n2720 VDD.n60 19.3944
R4339 VDD.n2720 VDD.n2719 19.3944
R4340 VDD.n2719 VDD.n2718 19.3944
R4341 VDD.n2718 VDD.n70 19.3944
R4342 VDD.n2712 VDD.n70 19.3944
R4343 VDD.n2712 VDD.n2711 19.3944
R4344 VDD.n2711 VDD.n2710 19.3944
R4345 VDD.n2710 VDD.n82 19.3944
R4346 VDD.n2704 VDD.n82 19.3944
R4347 VDD.n2704 VDD.n2703 19.3944
R4348 VDD.n2703 VDD.n2702 19.3944
R4349 VDD.n2702 VDD.n93 19.3944
R4350 VDD.n2696 VDD.n93 19.3944
R4351 VDD.n2446 VDD.n322 19.3944
R4352 VDD.n2446 VDD.n2443 19.3944
R4353 VDD.n2443 VDD.n2440 19.3944
R4354 VDD.n2440 VDD.n2439 19.3944
R4355 VDD.n2439 VDD.n2436 19.3944
R4356 VDD.n2436 VDD.n2435 19.3944
R4357 VDD.n2435 VDD.n2432 19.3944
R4358 VDD.n2432 VDD.n2431 19.3944
R4359 VDD.n2431 VDD.n2428 19.3944
R4360 VDD.n2428 VDD.n2427 19.3944
R4361 VDD.n2427 VDD.n2424 19.3944
R4362 VDD.n2424 VDD.n2423 19.3944
R4363 VDD.n2423 VDD.n2420 19.3944
R4364 VDD.n2420 VDD.n2419 19.3944
R4365 VDD.n2419 VDD.n2416 19.3944
R4366 VDD.n2416 VDD.n2415 19.3944
R4367 VDD.n2415 VDD.n2412 19.3944
R4368 VDD.n2412 VDD.n2411 19.3944
R4369 VDD.n2484 VDD.n273 19.3944
R4370 VDD.n2479 VDD.n273 19.3944
R4371 VDD.n2479 VDD.n2478 19.3944
R4372 VDD.n2478 VDD.n2477 19.3944
R4373 VDD.n2477 VDD.n2474 19.3944
R4374 VDD.n313 VDD.n308 19.3944
R4375 VDD.n2470 VDD.n2469 19.3944
R4376 VDD.n2469 VDD.n2467 19.3944
R4377 VDD.n2467 VDD.n2464 19.3944
R4378 VDD.n2464 VDD.n2463 19.3944
R4379 VDD.n2463 VDD.n2460 19.3944
R4380 VDD.n2460 VDD.n2459 19.3944
R4381 VDD.n2459 VDD.n2456 19.3944
R4382 VDD.n2456 VDD.n2455 19.3944
R4383 VDD.n2404 VDD.n340 19.3944
R4384 VDD.n2404 VDD.n2401 19.3944
R4385 VDD.n2401 VDD.n2398 19.3944
R4386 VDD.n2398 VDD.n2397 19.3944
R4387 VDD.n2397 VDD.n2394 19.3944
R4388 VDD.n2394 VDD.n2393 19.3944
R4389 VDD.n2393 VDD.n2390 19.3944
R4390 VDD.n2390 VDD.n2389 19.3944
R4391 VDD.n2389 VDD.n2386 19.3944
R4392 VDD.n2386 VDD.n2385 19.3944
R4393 VDD.n2385 VDD.n2382 19.3944
R4394 VDD.n2360 VDD.n352 19.3944
R4395 VDD.n2378 VDD.n2377 19.3944
R4396 VDD.n2377 VDD.n2375 19.3944
R4397 VDD.n2375 VDD.n2372 19.3944
R4398 VDD.n2372 VDD.n2371 19.3944
R4399 VDD.n1004 VDD.n1000 19.0066
R4400 VDD.n1326 VDD.n1276 19.0066
R4401 VDD.n2626 VDD.n165 19.0066
R4402 VDD.n2408 VDD.n340 19.0066
R4403 VDD.n1636 VDD.n666 17.3257
R4404 VDD.n1869 VDD.n510 17.3257
R4405 VDD.n2126 VDD.n1870 17.3257
R4406 VDD.n2332 VDD.n275 17.3257
R4407 VDD.n1071 VDD.n854 14.4382
R4408 VDD.n1079 VDD.n848 14.4382
R4409 VDD.n1079 VDD.n841 14.4382
R4410 VDD.n1087 VDD.n841 14.4382
R4411 VDD.n1087 VDD.n842 14.4382
R4412 VDD.n1095 VDD.n830 14.4382
R4413 VDD.n1103 VDD.n830 14.4382
R4414 VDD.n1111 VDD.n824 14.4382
R4415 VDD.n1119 VDD.n817 14.4382
R4416 VDD.n1119 VDD.n818 14.4382
R4417 VDD.n1127 VDD.n806 14.4382
R4418 VDD.n1136 VDD.n806 14.4382
R4419 VDD.n1144 VDD.n800 14.4382
R4420 VDD.n1152 VDD.n763 14.4382
R4421 VDD.n1152 VDD.n764 14.4382
R4422 VDD.n1160 VDD.n752 14.4382
R4423 VDD.n1168 VDD.n752 14.4382
R4424 VDD.n1176 VDD.n746 14.4382
R4425 VDD.n1184 VDD.n739 14.4382
R4426 VDD.n1184 VDD.n740 14.4382
R4427 VDD.n1192 VDD.n728 14.4382
R4428 VDD.n1200 VDD.n728 14.4382
R4429 VDD.n1200 VDD.n721 14.4382
R4430 VDD.n1209 VDD.n721 14.4382
R4431 VDD.n1399 VDD.n712 14.4382
R4432 VDD.n2490 VDD.n269 14.4382
R4433 VDD.n2498 VDD.n263 14.4382
R4434 VDD.n2498 VDD.n256 14.4382
R4435 VDD.n2506 VDD.n256 14.4382
R4436 VDD.n2506 VDD.n257 14.4382
R4437 VDD.n2514 VDD.n245 14.4382
R4438 VDD.n2522 VDD.n245 14.4382
R4439 VDD.n2530 VDD.n239 14.4382
R4440 VDD.n2538 VDD.n232 14.4382
R4441 VDD.n2538 VDD.n233 14.4382
R4442 VDD.n2546 VDD.n221 14.4382
R4443 VDD.n2554 VDD.n221 14.4382
R4444 VDD.n2732 VDD.n51 14.4382
R4445 VDD.n2731 VDD.n2730 14.4382
R4446 VDD.n2730 VDD.n55 14.4382
R4447 VDD.n2724 VDD.n2723 14.4382
R4448 VDD.n2723 VDD.n2722 14.4382
R4449 VDD.n2716 VDD.n72 14.4382
R4450 VDD.n2715 VDD.n2714 14.4382
R4451 VDD.n2714 VDD.n76 14.4382
R4452 VDD.n2708 VDD.n2707 14.4382
R4453 VDD.n2707 VDD.n2706 14.4382
R4454 VDD.n2706 VDD.n87 14.4382
R4455 VDD.n2700 VDD.n87 14.4382
R4456 VDD.n2699 VDD.n2698 14.4382
R4457 VDD.n1037 VDD.n1033 12.9944
R4458 VDD.n1038 VDD.n1037 12.9944
R4459 VDD.n1363 VDD.n1241 12.9944
R4460 VDD.n1363 VDD.n1238 12.9944
R4461 VDD.n2663 VDD.n130 12.9944
R4462 VDD.n2663 VDD.n127 12.9944
R4463 VDD.n2452 VDD.n322 12.9944
R4464 VDD.n2455 VDD.n2452 12.9944
R4465 VDD.n1111 VDD.t141 12.2725
R4466 VDD.t137 VDD.n746 12.2725
R4467 VDD.n2530 VDD.t143 12.2725
R4468 VDD.n72 VDD.t115 12.2725
R4469 VDD.t119 VDD.n800 11.9838
R4470 VDD.n1144 VDD.t121 11.9838
R4471 VDD.t149 VDD.n51 11.9838
R4472 VDD.n2732 VDD.t130 11.9838
R4473 VDD.t132 VDD.n824 11.695
R4474 VDD.n1176 VDD.t135 11.695
R4475 VDD.t117 VDD.n239 11.695
R4476 VDD.n2716 VDD.t160 11.695
R4477 VDD.n1634 VDD.n657 10.6151
R4478 VDD.n1644 VDD.n657 10.6151
R4479 VDD.n1645 VDD.n1644 10.6151
R4480 VDD.n1646 VDD.n1645 10.6151
R4481 VDD.n1646 VDD.n645 10.6151
R4482 VDD.n1657 VDD.n645 10.6151
R4483 VDD.n1658 VDD.n1657 10.6151
R4484 VDD.n1659 VDD.n1658 10.6151
R4485 VDD.n1659 VDD.n633 10.6151
R4486 VDD.n1669 VDD.n633 10.6151
R4487 VDD.n1670 VDD.n1669 10.6151
R4488 VDD.n1671 VDD.n1670 10.6151
R4489 VDD.n1671 VDD.n621 10.6151
R4490 VDD.n1681 VDD.n621 10.6151
R4491 VDD.n1682 VDD.n1681 10.6151
R4492 VDD.n1683 VDD.n1682 10.6151
R4493 VDD.n1683 VDD.n609 10.6151
R4494 VDD.n1693 VDD.n609 10.6151
R4495 VDD.n1694 VDD.n1693 10.6151
R4496 VDD.n1695 VDD.n1694 10.6151
R4497 VDD.n1695 VDD.n598 10.6151
R4498 VDD.n1705 VDD.n598 10.6151
R4499 VDD.n1706 VDD.n1705 10.6151
R4500 VDD.n1707 VDD.n1706 10.6151
R4501 VDD.n1707 VDD.n587 10.6151
R4502 VDD.n1717 VDD.n587 10.6151
R4503 VDD.n1718 VDD.n1717 10.6151
R4504 VDD.n1719 VDD.n1718 10.6151
R4505 VDD.n1719 VDD.n575 10.6151
R4506 VDD.n1729 VDD.n575 10.6151
R4507 VDD.n1730 VDD.n1729 10.6151
R4508 VDD.n1731 VDD.n1730 10.6151
R4509 VDD.n1731 VDD.n563 10.6151
R4510 VDD.n1741 VDD.n563 10.6151
R4511 VDD.n1742 VDD.n1741 10.6151
R4512 VDD.n1744 VDD.n1742 10.6151
R4513 VDD.n1744 VDD.n1743 10.6151
R4514 VDD.n1743 VDD.n549 10.6151
R4515 VDD.n1813 VDD.n549 10.6151
R4516 VDD.n1813 VDD.n1812 10.6151
R4517 VDD.n1811 VDD.n1809 10.6151
R4518 VDD.n1809 VDD.n1806 10.6151
R4519 VDD.n1806 VDD.n1805 10.6151
R4520 VDD.n1805 VDD.n1802 10.6151
R4521 VDD.n1802 VDD.n1801 10.6151
R4522 VDD.n1801 VDD.n1798 10.6151
R4523 VDD.n1798 VDD.n1797 10.6151
R4524 VDD.n1797 VDD.n1794 10.6151
R4525 VDD.n1794 VDD.n1793 10.6151
R4526 VDD.n1793 VDD.n1790 10.6151
R4527 VDD.n1790 VDD.n1789 10.6151
R4528 VDD.n1789 VDD.n1786 10.6151
R4529 VDD.n1786 VDD.n1785 10.6151
R4530 VDD.n1785 VDD.n1782 10.6151
R4531 VDD.n1782 VDD.n1781 10.6151
R4532 VDD.n1781 VDD.n1778 10.6151
R4533 VDD.n1778 VDD.n1777 10.6151
R4534 VDD.n1777 VDD.n1774 10.6151
R4535 VDD.n1774 VDD.n1773 10.6151
R4536 VDD.n1773 VDD.n1770 10.6151
R4537 VDD.n1770 VDD.n1769 10.6151
R4538 VDD.n1769 VDD.n1766 10.6151
R4539 VDD.n1764 VDD.n1761 10.6151
R4540 VDD.n1761 VDD.n1760 10.6151
R4541 VDD.n1582 VDD.n1581 10.6151
R4542 VDD.n1581 VDD.n1579 10.6151
R4543 VDD.n1579 VDD.n1578 10.6151
R4544 VDD.n1578 VDD.n1576 10.6151
R4545 VDD.n1576 VDD.n1575 10.6151
R4546 VDD.n1575 VDD.n1573 10.6151
R4547 VDD.n1573 VDD.n1572 10.6151
R4548 VDD.n1572 VDD.n1570 10.6151
R4549 VDD.n1570 VDD.n1569 10.6151
R4550 VDD.n1569 VDD.n1567 10.6151
R4551 VDD.n1567 VDD.n1566 10.6151
R4552 VDD.n1566 VDD.n1564 10.6151
R4553 VDD.n1564 VDD.n1563 10.6151
R4554 VDD.n1563 VDD.n1561 10.6151
R4555 VDD.n1561 VDD.n1560 10.6151
R4556 VDD.n1560 VDD.n1558 10.6151
R4557 VDD.n1558 VDD.n1557 10.6151
R4558 VDD.n1557 VDD.n1555 10.6151
R4559 VDD.n1555 VDD.n1554 10.6151
R4560 VDD.n1554 VDD.n1552 10.6151
R4561 VDD.n1552 VDD.n1551 10.6151
R4562 VDD.n1551 VDD.n686 10.6151
R4563 VDD.n1520 VDD.n686 10.6151
R4564 VDD.n1521 VDD.n1520 10.6151
R4565 VDD.n1538 VDD.n1521 10.6151
R4566 VDD.n1538 VDD.n1537 10.6151
R4567 VDD.n1537 VDD.n1536 10.6151
R4568 VDD.n1536 VDD.n1534 10.6151
R4569 VDD.n1534 VDD.n1533 10.6151
R4570 VDD.n1533 VDD.n1531 10.6151
R4571 VDD.n1531 VDD.n1530 10.6151
R4572 VDD.n1530 VDD.n1528 10.6151
R4573 VDD.n1528 VDD.n1527 10.6151
R4574 VDD.n1527 VDD.n1525 10.6151
R4575 VDD.n1525 VDD.n1524 10.6151
R4576 VDD.n1524 VDD.n1522 10.6151
R4577 VDD.n1522 VDD.n552 10.6151
R4578 VDD.n1755 VDD.n552 10.6151
R4579 VDD.n1756 VDD.n1755 10.6151
R4580 VDD.n1757 VDD.n1756 10.6151
R4581 VDD.n1633 VDD.n1632 10.6151
R4582 VDD.n1632 VDD.n670 10.6151
R4583 VDD.n1627 VDD.n670 10.6151
R4584 VDD.n1627 VDD.n1626 10.6151
R4585 VDD.n1626 VDD.n672 10.6151
R4586 VDD.n1621 VDD.n672 10.6151
R4587 VDD.n1621 VDD.n1620 10.6151
R4588 VDD.n1620 VDD.n1619 10.6151
R4589 VDD.n1619 VDD.n674 10.6151
R4590 VDD.n1613 VDD.n674 10.6151
R4591 VDD.n1613 VDD.n1612 10.6151
R4592 VDD.n1612 VDD.n1611 10.6151
R4593 VDD.n1607 VDD.n1606 10.6151
R4594 VDD.n1606 VDD.n678 10.6151
R4595 VDD.n1601 VDD.n678 10.6151
R4596 VDD.n1601 VDD.n1600 10.6151
R4597 VDD.n1600 VDD.n1599 10.6151
R4598 VDD.n1599 VDD.n680 10.6151
R4599 VDD.n1593 VDD.n680 10.6151
R4600 VDD.n1593 VDD.n1592 10.6151
R4601 VDD.n1592 VDD.n1591 10.6151
R4602 VDD.n1587 VDD.n1586 10.6151
R4603 VDD.n1586 VDD.n1583 10.6151
R4604 VDD.n1958 VDD.n1956 10.6151
R4605 VDD.n1959 VDD.n1958 10.6151
R4606 VDD.n1961 VDD.n1959 10.6151
R4607 VDD.n1962 VDD.n1961 10.6151
R4608 VDD.n1964 VDD.n1962 10.6151
R4609 VDD.n1965 VDD.n1964 10.6151
R4610 VDD.n1967 VDD.n1965 10.6151
R4611 VDD.n1968 VDD.n1967 10.6151
R4612 VDD.n1970 VDD.n1968 10.6151
R4613 VDD.n1971 VDD.n1970 10.6151
R4614 VDD.n1973 VDD.n1971 10.6151
R4615 VDD.n1974 VDD.n1973 10.6151
R4616 VDD.n1976 VDD.n1974 10.6151
R4617 VDD.n1977 VDD.n1976 10.6151
R4618 VDD.n2045 VDD.n1977 10.6151
R4619 VDD.n2045 VDD.n2044 10.6151
R4620 VDD.n2044 VDD.n2043 10.6151
R4621 VDD.n2043 VDD.n2041 10.6151
R4622 VDD.n2041 VDD.n2040 10.6151
R4623 VDD.n2040 VDD.n2003 10.6151
R4624 VDD.n2003 VDD.n2002 10.6151
R4625 VDD.n2002 VDD.n2000 10.6151
R4626 VDD.n2000 VDD.n1999 10.6151
R4627 VDD.n1999 VDD.n1997 10.6151
R4628 VDD.n1997 VDD.n1996 10.6151
R4629 VDD.n1996 VDD.n1994 10.6151
R4630 VDD.n1994 VDD.n1993 10.6151
R4631 VDD.n1993 VDD.n1991 10.6151
R4632 VDD.n1991 VDD.n1990 10.6151
R4633 VDD.n1990 VDD.n1988 10.6151
R4634 VDD.n1988 VDD.n1987 10.6151
R4635 VDD.n1987 VDD.n1985 10.6151
R4636 VDD.n1985 VDD.n1984 10.6151
R4637 VDD.n1984 VDD.n1982 10.6151
R4638 VDD.n1982 VDD.n1981 10.6151
R4639 VDD.n1981 VDD.n1979 10.6151
R4640 VDD.n1979 VDD.n1978 10.6151
R4641 VDD.n1978 VDD.n395 10.6151
R4642 VDD.n2280 VDD.n395 10.6151
R4643 VDD.n2281 VDD.n2280 10.6151
R4644 VDD.n1907 VDD.n508 10.6151
R4645 VDD.n1908 VDD.n1907 10.6151
R4646 VDD.n1909 VDD.n1908 10.6151
R4647 VDD.n1909 VDD.n1903 10.6151
R4648 VDD.n1915 VDD.n1903 10.6151
R4649 VDD.n1916 VDD.n1915 10.6151
R4650 VDD.n1917 VDD.n1916 10.6151
R4651 VDD.n1917 VDD.n1901 10.6151
R4652 VDD.n1923 VDD.n1901 10.6151
R4653 VDD.n1924 VDD.n1923 10.6151
R4654 VDD.n1925 VDD.n1924 10.6151
R4655 VDD.n1925 VDD.n1899 10.6151
R4656 VDD.n1931 VDD.n1899 10.6151
R4657 VDD.n1932 VDD.n1931 10.6151
R4658 VDD.n1933 VDD.n1932 10.6151
R4659 VDD.n1933 VDD.n1897 10.6151
R4660 VDD.n1939 VDD.n1897 10.6151
R4661 VDD.n1940 VDD.n1939 10.6151
R4662 VDD.n1941 VDD.n1940 10.6151
R4663 VDD.n1941 VDD.n1895 10.6151
R4664 VDD.n1947 VDD.n1895 10.6151
R4665 VDD.n1948 VDD.n1947 10.6151
R4666 VDD.n1950 VDD.n1891 10.6151
R4667 VDD.n1955 VDD.n1891 10.6151
R4668 VDD.n2129 VDD.n2128 10.6151
R4669 VDD.n2130 VDD.n2129 10.6151
R4670 VDD.n2130 VDD.n496 10.6151
R4671 VDD.n2140 VDD.n496 10.6151
R4672 VDD.n2141 VDD.n2140 10.6151
R4673 VDD.n2142 VDD.n2141 10.6151
R4674 VDD.n2142 VDD.n484 10.6151
R4675 VDD.n2152 VDD.n484 10.6151
R4676 VDD.n2153 VDD.n2152 10.6151
R4677 VDD.n2154 VDD.n2153 10.6151
R4678 VDD.n2154 VDD.n473 10.6151
R4679 VDD.n2164 VDD.n473 10.6151
R4680 VDD.n2165 VDD.n2164 10.6151
R4681 VDD.n2166 VDD.n2165 10.6151
R4682 VDD.n2166 VDD.n462 10.6151
R4683 VDD.n2176 VDD.n462 10.6151
R4684 VDD.n2177 VDD.n2176 10.6151
R4685 VDD.n2178 VDD.n2177 10.6151
R4686 VDD.n2178 VDD.n450 10.6151
R4687 VDD.n2188 VDD.n450 10.6151
R4688 VDD.n2189 VDD.n2188 10.6151
R4689 VDD.n2190 VDD.n2189 10.6151
R4690 VDD.n2190 VDD.n438 10.6151
R4691 VDD.n2200 VDD.n438 10.6151
R4692 VDD.n2201 VDD.n2200 10.6151
R4693 VDD.n2202 VDD.n2201 10.6151
R4694 VDD.n2202 VDD.n426 10.6151
R4695 VDD.n2212 VDD.n426 10.6151
R4696 VDD.n2213 VDD.n2212 10.6151
R4697 VDD.n2214 VDD.n2213 10.6151
R4698 VDD.n2214 VDD.n415 10.6151
R4699 VDD.n2224 VDD.n415 10.6151
R4700 VDD.n2225 VDD.n2224 10.6151
R4701 VDD.n2226 VDD.n2225 10.6151
R4702 VDD.n2226 VDD.n401 10.6151
R4703 VDD.n2273 VDD.n401 10.6151
R4704 VDD.n2274 VDD.n2273 10.6151
R4705 VDD.n2275 VDD.n2274 10.6151
R4706 VDD.n2275 VDD.n375 10.6151
R4707 VDD.n2330 VDD.n375 10.6151
R4708 VDD.n2329 VDD.n2328 10.6151
R4709 VDD.n2328 VDD.n376 10.6151
R4710 VDD.n2323 VDD.n376 10.6151
R4711 VDD.n2323 VDD.n2322 10.6151
R4712 VDD.n2322 VDD.n2321 10.6151
R4713 VDD.n2321 VDD.n379 10.6151
R4714 VDD.n2316 VDD.n379 10.6151
R4715 VDD.n2316 VDD.n2315 10.6151
R4716 VDD.n2315 VDD.n2314 10.6151
R4717 VDD.n2314 VDD.n382 10.6151
R4718 VDD.n2309 VDD.n382 10.6151
R4719 VDD.n2309 VDD.n2308 10.6151
R4720 VDD.n2304 VDD.n2303 10.6151
R4721 VDD.n2303 VDD.n2302 10.6151
R4722 VDD.n2302 VDD.n385 10.6151
R4723 VDD.n2297 VDD.n385 10.6151
R4724 VDD.n2297 VDD.n2296 10.6151
R4725 VDD.n2296 VDD.n2295 10.6151
R4726 VDD.n2295 VDD.n388 10.6151
R4727 VDD.n2290 VDD.n388 10.6151
R4728 VDD.n2290 VDD.n2289 10.6151
R4729 VDD.n2287 VDD.n393 10.6151
R4730 VDD.n2282 VDD.n393 10.6151
R4731 VDD.n2263 VDD.n2233 10.6151
R4732 VDD.n2234 VDD.n2233 10.6151
R4733 VDD.n2256 VDD.n2234 10.6151
R4734 VDD.n2256 VDD.n2255 10.6151
R4735 VDD.n2255 VDD.n2254 10.6151
R4736 VDD.n2254 VDD.n2236 10.6151
R4737 VDD.n2249 VDD.n2236 10.6151
R4738 VDD.n2249 VDD.n2248 10.6151
R4739 VDD.n2248 VDD.n2247 10.6151
R4740 VDD.n2247 VDD.n2239 10.6151
R4741 VDD.n2242 VDD.n2239 10.6151
R4742 VDD.n2242 VDD.n354 10.6151
R4743 VDD.n2356 VDD.n355 10.6151
R4744 VDD.n2351 VDD.n355 10.6151
R4745 VDD.n2351 VDD.n2350 10.6151
R4746 VDD.n2350 VDD.n2349 10.6151
R4747 VDD.n2349 VDD.n358 10.6151
R4748 VDD.n2344 VDD.n358 10.6151
R4749 VDD.n2344 VDD.n2343 10.6151
R4750 VDD.n2343 VDD.n2342 10.6151
R4751 VDD.n2342 VDD.n361 10.6151
R4752 VDD.n2337 VDD.n2336 10.6151
R4753 VDD.n2336 VDD.n2335 10.6151
R4754 VDD.n2071 VDD.n2070 10.6151
R4755 VDD.n2070 VDD.n2068 10.6151
R4756 VDD.n2068 VDD.n2067 10.6151
R4757 VDD.n2067 VDD.n2065 10.6151
R4758 VDD.n2065 VDD.n2064 10.6151
R4759 VDD.n2064 VDD.n2062 10.6151
R4760 VDD.n2062 VDD.n2061 10.6151
R4761 VDD.n2061 VDD.n2059 10.6151
R4762 VDD.n2059 VDD.n2058 10.6151
R4763 VDD.n2058 VDD.n2056 10.6151
R4764 VDD.n2056 VDD.n2055 10.6151
R4765 VDD.n2055 VDD.n2053 10.6151
R4766 VDD.n2053 VDD.n2052 10.6151
R4767 VDD.n2052 VDD.n2050 10.6151
R4768 VDD.n2050 VDD.n2049 10.6151
R4769 VDD.n2049 VDD.n1890 10.6151
R4770 VDD.n2005 VDD.n1890 10.6151
R4771 VDD.n2006 VDD.n2005 10.6151
R4772 VDD.n2036 VDD.n2006 10.6151
R4773 VDD.n2036 VDD.n2035 10.6151
R4774 VDD.n2035 VDD.n2034 10.6151
R4775 VDD.n2034 VDD.n2032 10.6151
R4776 VDD.n2032 VDD.n2031 10.6151
R4777 VDD.n2031 VDD.n2029 10.6151
R4778 VDD.n2029 VDD.n2028 10.6151
R4779 VDD.n2028 VDD.n2026 10.6151
R4780 VDD.n2026 VDD.n2025 10.6151
R4781 VDD.n2025 VDD.n2023 10.6151
R4782 VDD.n2023 VDD.n2022 10.6151
R4783 VDD.n2022 VDD.n2020 10.6151
R4784 VDD.n2020 VDD.n2019 10.6151
R4785 VDD.n2019 VDD.n2017 10.6151
R4786 VDD.n2017 VDD.n2016 10.6151
R4787 VDD.n2016 VDD.n2014 10.6151
R4788 VDD.n2014 VDD.n2013 10.6151
R4789 VDD.n2013 VDD.n2011 10.6151
R4790 VDD.n2011 VDD.n2010 10.6151
R4791 VDD.n2010 VDD.n2008 10.6151
R4792 VDD.n2008 VDD.n2007 10.6151
R4793 VDD.n2007 VDD.n367 10.6151
R4794 VDD.n2123 VDD.n2122 10.6151
R4795 VDD.n2122 VDD.n1875 10.6151
R4796 VDD.n2116 VDD.n1875 10.6151
R4797 VDD.n2116 VDD.n2115 10.6151
R4798 VDD.n2115 VDD.n2114 10.6151
R4799 VDD.n2114 VDD.n1877 10.6151
R4800 VDD.n2108 VDD.n1877 10.6151
R4801 VDD.n2108 VDD.n2107 10.6151
R4802 VDD.n2107 VDD.n2106 10.6151
R4803 VDD.n2106 VDD.n1879 10.6151
R4804 VDD.n2100 VDD.n1879 10.6151
R4805 VDD.n2100 VDD.n2099 10.6151
R4806 VDD.n2099 VDD.n2098 10.6151
R4807 VDD.n2098 VDD.n1881 10.6151
R4808 VDD.n2092 VDD.n1881 10.6151
R4809 VDD.n2092 VDD.n2091 10.6151
R4810 VDD.n2091 VDD.n2090 10.6151
R4811 VDD.n2090 VDD.n1883 10.6151
R4812 VDD.n2084 VDD.n1883 10.6151
R4813 VDD.n2084 VDD.n2083 10.6151
R4814 VDD.n2083 VDD.n2082 10.6151
R4815 VDD.n2082 VDD.n1885 10.6151
R4816 VDD.n2076 VDD.n2075 10.6151
R4817 VDD.n2075 VDD.n2074 10.6151
R4818 VDD.n2124 VDD.n502 10.6151
R4819 VDD.n2134 VDD.n502 10.6151
R4820 VDD.n2135 VDD.n2134 10.6151
R4821 VDD.n2136 VDD.n2135 10.6151
R4822 VDD.n2136 VDD.n491 10.6151
R4823 VDD.n2146 VDD.n491 10.6151
R4824 VDD.n2147 VDD.n2146 10.6151
R4825 VDD.n2148 VDD.n2147 10.6151
R4826 VDD.n2148 VDD.n479 10.6151
R4827 VDD.n2158 VDD.n479 10.6151
R4828 VDD.n2159 VDD.n2158 10.6151
R4829 VDD.n2160 VDD.n2159 10.6151
R4830 VDD.n2160 VDD.n467 10.6151
R4831 VDD.n2170 VDD.n467 10.6151
R4832 VDD.n2171 VDD.n2170 10.6151
R4833 VDD.n2172 VDD.n2171 10.6151
R4834 VDD.n2172 VDD.n456 10.6151
R4835 VDD.n2182 VDD.n456 10.6151
R4836 VDD.n2183 VDD.n2182 10.6151
R4837 VDD.n2184 VDD.n2183 10.6151
R4838 VDD.n2184 VDD.n444 10.6151
R4839 VDD.n2194 VDD.n444 10.6151
R4840 VDD.n2195 VDD.n2194 10.6151
R4841 VDD.n2196 VDD.n2195 10.6151
R4842 VDD.n2196 VDD.n432 10.6151
R4843 VDD.n2206 VDD.n432 10.6151
R4844 VDD.n2207 VDD.n2206 10.6151
R4845 VDD.n2208 VDD.n2207 10.6151
R4846 VDD.n2208 VDD.n421 10.6151
R4847 VDD.n2218 VDD.n421 10.6151
R4848 VDD.n2219 VDD.n2218 10.6151
R4849 VDD.n2220 VDD.n2219 10.6151
R4850 VDD.n2220 VDD.n409 10.6151
R4851 VDD.n2230 VDD.n409 10.6151
R4852 VDD.n2269 VDD.n2232 10.6151
R4853 VDD.n2269 VDD.n2268 10.6151
R4854 VDD.n2268 VDD.n2267 10.6151
R4855 VDD.n2267 VDD.n2266 10.6151
R4856 VDD.n2266 VDD.n2264 10.6151
R4857 VDD.n1639 VDD.n1638 10.6151
R4858 VDD.n1640 VDD.n1639 10.6151
R4859 VDD.n1640 VDD.n651 10.6151
R4860 VDD.n1650 VDD.n651 10.6151
R4861 VDD.n1651 VDD.n1650 10.6151
R4862 VDD.n1653 VDD.n639 10.6151
R4863 VDD.n1663 VDD.n639 10.6151
R4864 VDD.n1664 VDD.n1663 10.6151
R4865 VDD.n1665 VDD.n1664 10.6151
R4866 VDD.n1665 VDD.n627 10.6151
R4867 VDD.n1675 VDD.n627 10.6151
R4868 VDD.n1676 VDD.n1675 10.6151
R4869 VDD.n1677 VDD.n1676 10.6151
R4870 VDD.n1677 VDD.n615 10.6151
R4871 VDD.n1687 VDD.n615 10.6151
R4872 VDD.n1688 VDD.n1687 10.6151
R4873 VDD.n1689 VDD.n1688 10.6151
R4874 VDD.n1689 VDD.n603 10.6151
R4875 VDD.n1699 VDD.n603 10.6151
R4876 VDD.n1700 VDD.n1699 10.6151
R4877 VDD.n1701 VDD.n1700 10.6151
R4878 VDD.n1701 VDD.n592 10.6151
R4879 VDD.n1711 VDD.n592 10.6151
R4880 VDD.n1712 VDD.n1711 10.6151
R4881 VDD.n1713 VDD.n1712 10.6151
R4882 VDD.n1713 VDD.n580 10.6151
R4883 VDD.n1723 VDD.n580 10.6151
R4884 VDD.n1724 VDD.n1723 10.6151
R4885 VDD.n1725 VDD.n1724 10.6151
R4886 VDD.n1725 VDD.n569 10.6151
R4887 VDD.n1735 VDD.n569 10.6151
R4888 VDD.n1736 VDD.n1735 10.6151
R4889 VDD.n1737 VDD.n1736 10.6151
R4890 VDD.n1737 VDD.n556 10.6151
R4891 VDD.n1748 VDD.n556 10.6151
R4892 VDD.n1749 VDD.n1748 10.6151
R4893 VDD.n1751 VDD.n1749 10.6151
R4894 VDD.n1751 VDD.n1750 10.6151
R4895 VDD.n1750 VDD.n539 10.6151
R4896 VDD.n1867 VDD.n1866 10.6151
R4897 VDD.n1866 VDD.n1865 10.6151
R4898 VDD.n1865 VDD.n1862 10.6151
R4899 VDD.n1862 VDD.n1861 10.6151
R4900 VDD.n1861 VDD.n1858 10.6151
R4901 VDD.n1858 VDD.n1857 10.6151
R4902 VDD.n1857 VDD.n1854 10.6151
R4903 VDD.n1854 VDD.n1853 10.6151
R4904 VDD.n1853 VDD.n1850 10.6151
R4905 VDD.n1850 VDD.n1849 10.6151
R4906 VDD.n1849 VDD.n1846 10.6151
R4907 VDD.n1846 VDD.n1845 10.6151
R4908 VDD.n1845 VDD.n1842 10.6151
R4909 VDD.n1842 VDD.n1841 10.6151
R4910 VDD.n1841 VDD.n1838 10.6151
R4911 VDD.n1838 VDD.n1837 10.6151
R4912 VDD.n1837 VDD.n1834 10.6151
R4913 VDD.n1834 VDD.n1833 10.6151
R4914 VDD.n1833 VDD.n1830 10.6151
R4915 VDD.n1830 VDD.n1829 10.6151
R4916 VDD.n1829 VDD.n1826 10.6151
R4917 VDD.n1826 VDD.n1825 10.6151
R4918 VDD.n1822 VDD.n1821 10.6151
R4919 VDD.n1821 VDD.n1819 10.6151
R4920 VDD.n1471 VDD.n1469 10.6151
R4921 VDD.n1472 VDD.n1471 10.6151
R4922 VDD.n1474 VDD.n1472 10.6151
R4923 VDD.n1475 VDD.n1474 10.6151
R4924 VDD.n1477 VDD.n1475 10.6151
R4925 VDD.n1478 VDD.n1477 10.6151
R4926 VDD.n1480 VDD.n1478 10.6151
R4927 VDD.n1481 VDD.n1480 10.6151
R4928 VDD.n1483 VDD.n1481 10.6151
R4929 VDD.n1484 VDD.n1483 10.6151
R4930 VDD.n1486 VDD.n1484 10.6151
R4931 VDD.n1487 VDD.n1486 10.6151
R4932 VDD.n1489 VDD.n1487 10.6151
R4933 VDD.n1490 VDD.n1489 10.6151
R4934 VDD.n1492 VDD.n1490 10.6151
R4935 VDD.n1493 VDD.n1492 10.6151
R4936 VDD.n1495 VDD.n1493 10.6151
R4937 VDD.n1496 VDD.n1495 10.6151
R4938 VDD.n1498 VDD.n1496 10.6151
R4939 VDD.n1499 VDD.n1498 10.6151
R4940 VDD.n1547 VDD.n1499 10.6151
R4941 VDD.n1547 VDD.n1546 10.6151
R4942 VDD.n1546 VDD.n1545 10.6151
R4943 VDD.n1545 VDD.n1543 10.6151
R4944 VDD.n1543 VDD.n1542 10.6151
R4945 VDD.n1542 VDD.n1518 10.6151
R4946 VDD.n1518 VDD.n1517 10.6151
R4947 VDD.n1517 VDD.n1515 10.6151
R4948 VDD.n1515 VDD.n1514 10.6151
R4949 VDD.n1514 VDD.n1512 10.6151
R4950 VDD.n1512 VDD.n1511 10.6151
R4951 VDD.n1511 VDD.n1509 10.6151
R4952 VDD.n1509 VDD.n1508 10.6151
R4953 VDD.n1508 VDD.n1506 10.6151
R4954 VDD.n1506 VDD.n1505 10.6151
R4955 VDD.n1505 VDD.n1503 10.6151
R4956 VDD.n1503 VDD.n1502 10.6151
R4957 VDD.n1502 VDD.n1500 10.6151
R4958 VDD.n1500 VDD.n543 10.6151
R4959 VDD.n1818 VDD.n543 10.6151
R4960 VDD.n1420 VDD.n664 10.6151
R4961 VDD.n1421 VDD.n1420 10.6151
R4962 VDD.n1422 VDD.n1421 10.6151
R4963 VDD.n1422 VDD.n1416 10.6151
R4964 VDD.n1428 VDD.n1416 10.6151
R4965 VDD.n1429 VDD.n1428 10.6151
R4966 VDD.n1430 VDD.n1429 10.6151
R4967 VDD.n1430 VDD.n1414 10.6151
R4968 VDD.n1436 VDD.n1414 10.6151
R4969 VDD.n1437 VDD.n1436 10.6151
R4970 VDD.n1438 VDD.n1437 10.6151
R4971 VDD.n1438 VDD.n1412 10.6151
R4972 VDD.n1445 VDD.n1444 10.6151
R4973 VDD.n1446 VDD.n1445 10.6151
R4974 VDD.n1446 VDD.n693 10.6151
R4975 VDD.n1452 VDD.n693 10.6151
R4976 VDD.n1453 VDD.n1452 10.6151
R4977 VDD.n1454 VDD.n1453 10.6151
R4978 VDD.n1454 VDD.n691 10.6151
R4979 VDD.n1460 VDD.n691 10.6151
R4980 VDD.n1461 VDD.n1460 10.6151
R4981 VDD.n1463 VDD.n687 10.6151
R4982 VDD.n1468 VDD.n687 10.6151
R4983 VDD.n1071 VDD.t40 9.96251
R4984 VDD.t44 VDD.n712 9.96251
R4985 VDD.n2490 VDD.t71 9.96251
R4986 VDD.t63 VDD.n2699 9.96251
R4987 VDD.n1636 VDD.n659 9.81813
R4988 VDD.n1642 VDD.n659 9.81813
R4989 VDD.n1642 VDD.n662 9.81813
R4990 VDD.n1648 VDD.n655 9.81813
R4991 VDD.n1655 VDD.n641 9.81813
R4992 VDD.n1661 VDD.n641 9.81813
R4993 VDD.n1661 VDD.n635 9.81813
R4994 VDD.n1667 VDD.n635 9.81813
R4995 VDD.n1673 VDD.n629 9.81813
R4996 VDD.n1679 VDD.n623 9.81813
R4997 VDD.n1685 VDD.n617 9.81813
R4998 VDD.n1691 VDD.n611 9.81813
R4999 VDD.n1697 VDD.n605 9.81813
R5000 VDD.n1703 VDD.n594 9.81813
R5001 VDD.n1709 VDD.n594 9.81813
R5002 VDD.n1715 VDD.n582 9.81813
R5003 VDD.n1721 VDD.n582 9.81813
R5004 VDD.n1721 VDD.n585 9.81813
R5005 VDD.n1733 VDD.n571 9.81813
R5006 VDD.n1733 VDD.n565 9.81813
R5007 VDD.n1739 VDD.n565 9.81813
R5008 VDD.n1746 VDD.n558 9.81813
R5009 VDD.n1753 VDD.n554 9.81813
R5010 VDD.n1815 VDD.n510 9.81813
R5011 VDD.n2126 VDD.n1873 9.81813
R5012 VDD.n2132 VDD.n506 9.81813
R5013 VDD.n2138 VDD.n500 9.81813
R5014 VDD.n2144 VDD.n486 9.81813
R5015 VDD.n2150 VDD.n486 9.81813
R5016 VDD.n2150 VDD.n489 9.81813
R5017 VDD.n2162 VDD.n475 9.81813
R5018 VDD.n2162 VDD.n469 9.81813
R5019 VDD.n2168 VDD.n469 9.81813
R5020 VDD.n2174 VDD.n458 9.81813
R5021 VDD.n2180 VDD.n458 9.81813
R5022 VDD.n2186 VDD.n454 9.81813
R5023 VDD.n2192 VDD.n448 9.81813
R5024 VDD.n2198 VDD.n442 9.81813
R5025 VDD.n2204 VDD.n436 9.81813
R5026 VDD.n2210 VDD.n430 9.81813
R5027 VDD.n2216 VDD.n417 9.81813
R5028 VDD.n2222 VDD.n417 9.81813
R5029 VDD.n2222 VDD.n411 9.81813
R5030 VDD.n2228 VDD.n411 9.81813
R5031 VDD.n2271 VDD.n403 9.81813
R5032 VDD.n2277 VDD.n397 9.81813
R5033 VDD.n2277 VDD.n370 9.81813
R5034 VDD.n2332 VDD.n370 9.81813
R5035 VDD.n1384 VDD.n676 9.61581
R5036 VDD.n2472 VDD.n310 9.61581
R5037 VDD.n2380 VDD.n2357 9.61581
R5038 VDD.n1411 VDD.n1410 9.61581
R5039 VDD.t4 VDD.n605 9.385
R5040 VDD.n1549 VDD.t32 9.385
R5041 VDD.n2038 VDD.t1 9.385
R5042 VDD.n454 VDD.t36 9.385
R5043 VDD.n1361 VDD.n1241 9.3005
R5044 VDD.n1360 VDD.n1359 9.3005
R5045 VDD.n1246 VDD.n1245 9.3005
R5046 VDD.n1354 VDD.n1249 9.3005
R5047 VDD.n1353 VDD.n1250 9.3005
R5048 VDD.n1352 VDD.n1251 9.3005
R5049 VDD.n1255 VDD.n1252 9.3005
R5050 VDD.n1347 VDD.n1256 9.3005
R5051 VDD.n1346 VDD.n1257 9.3005
R5052 VDD.n1345 VDD.n1258 9.3005
R5053 VDD.n1262 VDD.n1259 9.3005
R5054 VDD.n1340 VDD.n1263 9.3005
R5055 VDD.n1339 VDD.n1264 9.3005
R5056 VDD.n1338 VDD.n1265 9.3005
R5057 VDD.n1269 VDD.n1266 9.3005
R5058 VDD.n1333 VDD.n1270 9.3005
R5059 VDD.n1332 VDD.n1271 9.3005
R5060 VDD.n1331 VDD.n1272 9.3005
R5061 VDD.n1279 VDD.n1273 9.3005
R5062 VDD.n1326 VDD.n1325 9.3005
R5063 VDD.n1324 VDD.n1276 9.3005
R5064 VDD.n1323 VDD.n1322 9.3005
R5065 VDD.n1281 VDD.n1280 9.3005
R5066 VDD.n1317 VDD.n1284 9.3005
R5067 VDD.n1316 VDD.n1285 9.3005
R5068 VDD.n1315 VDD.n1286 9.3005
R5069 VDD.n1290 VDD.n1287 9.3005
R5070 VDD.n1310 VDD.n1291 9.3005
R5071 VDD.n1309 VDD.n1292 9.3005
R5072 VDD.n1308 VDD.n1293 9.3005
R5073 VDD.n1294 VDD.n695 9.3005
R5074 VDD.n1363 VDD.n1362 9.3005
R5075 VDD.n1377 VDD.n1224 9.3005
R5076 VDD.n1376 VDD.n1229 9.3005
R5077 VDD.n1375 VDD.n1230 9.3005
R5078 VDD.n1234 VDD.n1231 9.3005
R5079 VDD.n1370 VDD.n1235 9.3005
R5080 VDD.n1369 VDD.n1236 9.3005
R5081 VDD.n1368 VDD.n1237 9.3005
R5082 VDD.n1244 VDD.n1238 9.3005
R5083 VDD.n1393 VDD.n1214 9.3005
R5084 VDD.n1218 VDD.n1215 9.3005
R5085 VDD.n1388 VDD.n1219 9.3005
R5086 VDD.n1387 VDD.n1220 9.3005
R5087 VDD.n1395 VDD.n1394 9.3005
R5088 VDD.n1147 VDD.n1146 9.3005
R5089 VDD.n1148 VDD.n766 9.3005
R5090 VDD.n1150 VDD.n1149 9.3005
R5091 VDD.n756 VDD.n755 9.3005
R5092 VDD.n1163 VDD.n1162 9.3005
R5093 VDD.n1164 VDD.n754 9.3005
R5094 VDD.n1166 VDD.n1165 9.3005
R5095 VDD.n744 VDD.n743 9.3005
R5096 VDD.n1179 VDD.n1178 9.3005
R5097 VDD.n1180 VDD.n742 9.3005
R5098 VDD.n1182 VDD.n1181 9.3005
R5099 VDD.n732 VDD.n731 9.3005
R5100 VDD.n1195 VDD.n1194 9.3005
R5101 VDD.n1196 VDD.n730 9.3005
R5102 VDD.n1198 VDD.n1197 9.3005
R5103 VDD.n719 VDD.n718 9.3005
R5104 VDD.n1212 VDD.n1211 9.3005
R5105 VDD.n1213 VDD.n717 9.3005
R5106 VDD.n1397 VDD.n1396 9.3005
R5107 VDD.n2408 VDD.n2407 9.3005
R5108 VDD.n2411 VDD.n339 9.3005
R5109 VDD.n2412 VDD.n338 9.3005
R5110 VDD.n2415 VDD.n337 9.3005
R5111 VDD.n2416 VDD.n336 9.3005
R5112 VDD.n2419 VDD.n335 9.3005
R5113 VDD.n2420 VDD.n334 9.3005
R5114 VDD.n2423 VDD.n333 9.3005
R5115 VDD.n2424 VDD.n332 9.3005
R5116 VDD.n2427 VDD.n331 9.3005
R5117 VDD.n2428 VDD.n330 9.3005
R5118 VDD.n2431 VDD.n329 9.3005
R5119 VDD.n2432 VDD.n328 9.3005
R5120 VDD.n2435 VDD.n327 9.3005
R5121 VDD.n2436 VDD.n326 9.3005
R5122 VDD.n2439 VDD.n325 9.3005
R5123 VDD.n2440 VDD.n324 9.3005
R5124 VDD.n2443 VDD.n323 9.3005
R5125 VDD.n2447 VDD.n2446 9.3005
R5126 VDD.n2448 VDD.n322 9.3005
R5127 VDD.n2452 VDD.n2449 9.3005
R5128 VDD.n2455 VDD.n321 9.3005
R5129 VDD.n2456 VDD.n320 9.3005
R5130 VDD.n2459 VDD.n319 9.3005
R5131 VDD.n2460 VDD.n318 9.3005
R5132 VDD.n2463 VDD.n317 9.3005
R5133 VDD.n2464 VDD.n316 9.3005
R5134 VDD.n2467 VDD.n315 9.3005
R5135 VDD.n2469 VDD.n309 9.3005
R5136 VDD.n2477 VDD.n307 9.3005
R5137 VDD.n2478 VDD.n306 9.3005
R5138 VDD.n2479 VDD.n305 9.3005
R5139 VDD.n273 VDD.n272 9.3005
R5140 VDD.n2485 VDD.n2484 9.3005
R5141 VDD.n2488 VDD.n2487 9.3005
R5142 VDD.n261 VDD.n260 9.3005
R5143 VDD.n2501 VDD.n2500 9.3005
R5144 VDD.n2502 VDD.n259 9.3005
R5145 VDD.n2504 VDD.n2503 9.3005
R5146 VDD.n249 VDD.n248 9.3005
R5147 VDD.n2517 VDD.n2516 9.3005
R5148 VDD.n2518 VDD.n247 9.3005
R5149 VDD.n2520 VDD.n2519 9.3005
R5150 VDD.n237 VDD.n236 9.3005
R5151 VDD.n2533 VDD.n2532 9.3005
R5152 VDD.n2534 VDD.n235 9.3005
R5153 VDD.n2536 VDD.n2535 9.3005
R5154 VDD.n225 VDD.n224 9.3005
R5155 VDD.n2549 VDD.n2548 9.3005
R5156 VDD.n2550 VDD.n223 9.3005
R5157 VDD.n2552 VDD.n2551 9.3005
R5158 VDD.n47 VDD.n45 9.3005
R5159 VDD.n2486 VDD.n271 9.3005
R5160 VDD.n2735 VDD.n2734 9.3005
R5161 VDD.n48 VDD.n46 9.3005
R5162 VDD.n2728 VDD.n57 9.3005
R5163 VDD.n2727 VDD.n58 9.3005
R5164 VDD.n2726 VDD.n59 9.3005
R5165 VDD.n66 VDD.n60 9.3005
R5166 VDD.n2720 VDD.n67 9.3005
R5167 VDD.n2719 VDD.n68 9.3005
R5168 VDD.n2718 VDD.n69 9.3005
R5169 VDD.n78 VDD.n70 9.3005
R5170 VDD.n2712 VDD.n79 9.3005
R5171 VDD.n2711 VDD.n80 9.3005
R5172 VDD.n2710 VDD.n81 9.3005
R5173 VDD.n89 VDD.n82 9.3005
R5174 VDD.n2704 VDD.n90 9.3005
R5175 VDD.n2703 VDD.n91 9.3005
R5176 VDD.n2702 VDD.n92 9.3005
R5177 VDD.n100 VDD.n93 9.3005
R5178 VDD.n2696 VDD.n2695 9.3005
R5179 VDD.n2692 VDD.n101 9.3005
R5180 VDD.n2691 VDD.n104 9.3005
R5181 VDD.n108 VDD.n105 9.3005
R5182 VDD.n109 VDD.n106 9.3005
R5183 VDD.n2684 VDD.n110 9.3005
R5184 VDD.n2683 VDD.n111 9.3005
R5185 VDD.n2682 VDD.n112 9.3005
R5186 VDD.n116 VDD.n113 9.3005
R5187 VDD.n2677 VDD.n117 9.3005
R5188 VDD.n2676 VDD.n118 9.3005
R5189 VDD.n2675 VDD.n119 9.3005
R5190 VDD.n123 VDD.n120 9.3005
R5191 VDD.n2670 VDD.n124 9.3005
R5192 VDD.n2669 VDD.n125 9.3005
R5193 VDD.n2668 VDD.n126 9.3005
R5194 VDD.n133 VDD.n127 9.3005
R5195 VDD.n2663 VDD.n2662 9.3005
R5196 VDD.n2661 VDD.n130 9.3005
R5197 VDD.n2660 VDD.n2659 9.3005
R5198 VDD.n135 VDD.n134 9.3005
R5199 VDD.n2654 VDD.n138 9.3005
R5200 VDD.n2653 VDD.n139 9.3005
R5201 VDD.n2652 VDD.n140 9.3005
R5202 VDD.n144 VDD.n141 9.3005
R5203 VDD.n2647 VDD.n145 9.3005
R5204 VDD.n2646 VDD.n146 9.3005
R5205 VDD.n2645 VDD.n147 9.3005
R5206 VDD.n151 VDD.n148 9.3005
R5207 VDD.n2640 VDD.n152 9.3005
R5208 VDD.n2639 VDD.n153 9.3005
R5209 VDD.n2638 VDD.n154 9.3005
R5210 VDD.n158 VDD.n155 9.3005
R5211 VDD.n2633 VDD.n159 9.3005
R5212 VDD.n2632 VDD.n160 9.3005
R5213 VDD.n2631 VDD.n161 9.3005
R5214 VDD.n168 VDD.n162 9.3005
R5215 VDD.n2626 VDD.n2625 9.3005
R5216 VDD.n2624 VDD.n165 9.3005
R5217 VDD.n2623 VDD.n2622 9.3005
R5218 VDD.n170 VDD.n169 9.3005
R5219 VDD.n2617 VDD.n173 9.3005
R5220 VDD.n2616 VDD.n174 9.3005
R5221 VDD.n2615 VDD.n175 9.3005
R5222 VDD.n179 VDD.n176 9.3005
R5223 VDD.n2610 VDD.n180 9.3005
R5224 VDD.n2609 VDD.n181 9.3005
R5225 VDD.n2608 VDD.n182 9.3005
R5226 VDD.n186 VDD.n183 9.3005
R5227 VDD.n2603 VDD.n187 9.3005
R5228 VDD.n2602 VDD.n188 9.3005
R5229 VDD.n2601 VDD.n189 9.3005
R5230 VDD.n193 VDD.n190 9.3005
R5231 VDD.n2596 VDD.n194 9.3005
R5232 VDD.n2595 VDD.n195 9.3005
R5233 VDD.n2594 VDD.n196 9.3005
R5234 VDD.n202 VDD.n197 9.3005
R5235 VDD.n2589 VDD.n2588 9.3005
R5236 VDD.n2694 VDD.n2693 9.3005
R5237 VDD.n2493 VDD.n2492 9.3005
R5238 VDD.n2494 VDD.n265 9.3005
R5239 VDD.n2496 VDD.n2495 9.3005
R5240 VDD.n254 VDD.n253 9.3005
R5241 VDD.n2509 VDD.n2508 9.3005
R5242 VDD.n2510 VDD.n252 9.3005
R5243 VDD.n2512 VDD.n2511 9.3005
R5244 VDD.n243 VDD.n242 9.3005
R5245 VDD.n2525 VDD.n2524 9.3005
R5246 VDD.n2526 VDD.n241 9.3005
R5247 VDD.n2528 VDD.n2527 9.3005
R5248 VDD.n230 VDD.n229 9.3005
R5249 VDD.n2541 VDD.n2540 9.3005
R5250 VDD.n2542 VDD.n228 9.3005
R5251 VDD.n2544 VDD.n2543 9.3005
R5252 VDD.n218 VDD.n217 9.3005
R5253 VDD.n2557 VDD.n2556 9.3005
R5254 VDD.n2558 VDD.n216 9.3005
R5255 VDD.n2560 VDD.n2559 9.3005
R5256 VDD.n2561 VDD.n215 9.3005
R5257 VDD.n2563 VDD.n2562 9.3005
R5258 VDD.n2564 VDD.n214 9.3005
R5259 VDD.n2566 VDD.n2565 9.3005
R5260 VDD.n2567 VDD.n212 9.3005
R5261 VDD.n2569 VDD.n2568 9.3005
R5262 VDD.n2570 VDD.n211 9.3005
R5263 VDD.n2572 VDD.n2571 9.3005
R5264 VDD.n2573 VDD.n209 9.3005
R5265 VDD.n2575 VDD.n2574 9.3005
R5266 VDD.n2576 VDD.n208 9.3005
R5267 VDD.n2578 VDD.n2577 9.3005
R5268 VDD.n2579 VDD.n206 9.3005
R5269 VDD.n2581 VDD.n2580 9.3005
R5270 VDD.n2582 VDD.n205 9.3005
R5271 VDD.n2584 VDD.n2583 9.3005
R5272 VDD.n2585 VDD.n203 9.3005
R5273 VDD.n2587 VDD.n2586 9.3005
R5274 VDD.n267 VDD.n266 9.3005
R5275 VDD.n2366 VDD.n2365 9.3005
R5276 VDD.n2371 VDD.n2364 9.3005
R5277 VDD.n2372 VDD.n2363 9.3005
R5278 VDD.n2375 VDD.n2362 9.3005
R5279 VDD.n2377 VDD.n353 9.3005
R5280 VDD.n2385 VDD.n351 9.3005
R5281 VDD.n2386 VDD.n350 9.3005
R5282 VDD.n2389 VDD.n349 9.3005
R5283 VDD.n2390 VDD.n348 9.3005
R5284 VDD.n2393 VDD.n347 9.3005
R5285 VDD.n2394 VDD.n346 9.3005
R5286 VDD.n2397 VDD.n345 9.3005
R5287 VDD.n2398 VDD.n344 9.3005
R5288 VDD.n2401 VDD.n343 9.3005
R5289 VDD.n2405 VDD.n2404 9.3005
R5290 VDD.n2406 VDD.n340 9.3005
R5291 VDD.n1409 VDD.n1408 9.3005
R5292 VDD.n1407 VDD.n698 9.3005
R5293 VDD.n1406 VDD.n1405 9.3005
R5294 VDD.n1404 VDD.n703 9.3005
R5295 VDD.n1403 VDD.n1402 9.3005
R5296 VDD.n1074 VDD.n1073 9.3005
R5297 VDD.n1075 VDD.n850 9.3005
R5298 VDD.n1077 VDD.n1076 9.3005
R5299 VDD.n839 VDD.n838 9.3005
R5300 VDD.n1090 VDD.n1089 9.3005
R5301 VDD.n1091 VDD.n837 9.3005
R5302 VDD.n1093 VDD.n1092 9.3005
R5303 VDD.n828 VDD.n827 9.3005
R5304 VDD.n1106 VDD.n1105 9.3005
R5305 VDD.n1107 VDD.n826 9.3005
R5306 VDD.n1109 VDD.n1108 9.3005
R5307 VDD.n815 VDD.n814 9.3005
R5308 VDD.n1122 VDD.n1121 9.3005
R5309 VDD.n1123 VDD.n813 9.3005
R5310 VDD.n1125 VDD.n1124 9.3005
R5311 VDD.n804 VDD.n803 9.3005
R5312 VDD.n1139 VDD.n1138 9.3005
R5313 VDD.n1140 VDD.n802 9.3005
R5314 VDD.n1142 VDD.n1141 9.3005
R5315 VDD.n761 VDD.n760 9.3005
R5316 VDD.n1155 VDD.n1154 9.3005
R5317 VDD.n1156 VDD.n759 9.3005
R5318 VDD.n1158 VDD.n1157 9.3005
R5319 VDD.n750 VDD.n749 9.3005
R5320 VDD.n1171 VDD.n1170 9.3005
R5321 VDD.n1172 VDD.n748 9.3005
R5322 VDD.n1174 VDD.n1173 9.3005
R5323 VDD.n737 VDD.n736 9.3005
R5324 VDD.n1187 VDD.n1186 9.3005
R5325 VDD.n1188 VDD.n735 9.3005
R5326 VDD.n1190 VDD.n1189 9.3005
R5327 VDD.n726 VDD.n725 9.3005
R5328 VDD.n1203 VDD.n1202 9.3005
R5329 VDD.n1204 VDD.n723 9.3005
R5330 VDD.n1207 VDD.n1206 9.3005
R5331 VDD.n1205 VDD.n724 9.3005
R5332 VDD.n711 VDD.n704 9.3005
R5333 VDD.n852 VDD.n851 9.3005
R5334 VDD.n973 VDD.n972 9.3005
R5335 VDD.n974 VDD.n965 9.3005
R5336 VDD.n976 VDD.n975 9.3005
R5337 VDD.n977 VDD.n960 9.3005
R5338 VDD.n979 VDD.n978 9.3005
R5339 VDD.n980 VDD.n959 9.3005
R5340 VDD.n982 VDD.n981 9.3005
R5341 VDD.n983 VDD.n954 9.3005
R5342 VDD.n985 VDD.n984 9.3005
R5343 VDD.n986 VDD.n953 9.3005
R5344 VDD.n988 VDD.n987 9.3005
R5345 VDD.n989 VDD.n948 9.3005
R5346 VDD.n991 VDD.n990 9.3005
R5347 VDD.n992 VDD.n947 9.3005
R5348 VDD.n994 VDD.n993 9.3005
R5349 VDD.n995 VDD.n942 9.3005
R5350 VDD.n997 VDD.n996 9.3005
R5351 VDD.n998 VDD.n941 9.3005
R5352 VDD.n1000 VDD.n999 9.3005
R5353 VDD.n1004 VDD.n937 9.3005
R5354 VDD.n1006 VDD.n1005 9.3005
R5355 VDD.n1007 VDD.n936 9.3005
R5356 VDD.n1009 VDD.n1008 9.3005
R5357 VDD.n1010 VDD.n931 9.3005
R5358 VDD.n1012 VDD.n1011 9.3005
R5359 VDD.n1013 VDD.n930 9.3005
R5360 VDD.n1015 VDD.n1014 9.3005
R5361 VDD.n1016 VDD.n925 9.3005
R5362 VDD.n1018 VDD.n1017 9.3005
R5363 VDD.n1019 VDD.n924 9.3005
R5364 VDD.n1021 VDD.n1020 9.3005
R5365 VDD.n1022 VDD.n919 9.3005
R5366 VDD.n1024 VDD.n1023 9.3005
R5367 VDD.n1025 VDD.n918 9.3005
R5368 VDD.n1027 VDD.n1026 9.3005
R5369 VDD.n1028 VDD.n913 9.3005
R5370 VDD.n1030 VDD.n1029 9.3005
R5371 VDD.n1031 VDD.n912 9.3005
R5372 VDD.n1033 VDD.n1032 9.3005
R5373 VDD.n1037 VDD.n908 9.3005
R5374 VDD.n1039 VDD.n1038 9.3005
R5375 VDD.n1040 VDD.n907 9.3005
R5376 VDD.n1042 VDD.n1041 9.3005
R5377 VDD.n1043 VDD.n902 9.3005
R5378 VDD.n1045 VDD.n1044 9.3005
R5379 VDD.n1046 VDD.n901 9.3005
R5380 VDD.n1048 VDD.n1047 9.3005
R5381 VDD.n1049 VDD.n896 9.3005
R5382 VDD.n1051 VDD.n1050 9.3005
R5383 VDD.n1052 VDD.n895 9.3005
R5384 VDD.n1054 VDD.n1053 9.3005
R5385 VDD.n1055 VDD.n890 9.3005
R5386 VDD.n1057 VDD.n1056 9.3005
R5387 VDD.n1058 VDD.n889 9.3005
R5388 VDD.n1060 VDD.n1059 9.3005
R5389 VDD.n858 VDD.n857 9.3005
R5390 VDD.n1066 VDD.n1065 9.3005
R5391 VDD.n968 VDD.n966 9.3005
R5392 VDD.n1069 VDD.n1068 9.3005
R5393 VDD.n846 VDD.n845 9.3005
R5394 VDD.n1082 VDD.n1081 9.3005
R5395 VDD.n1083 VDD.n844 9.3005
R5396 VDD.n1085 VDD.n1084 9.3005
R5397 VDD.n834 VDD.n833 9.3005
R5398 VDD.n1098 VDD.n1097 9.3005
R5399 VDD.n1099 VDD.n832 9.3005
R5400 VDD.n1101 VDD.n1100 9.3005
R5401 VDD.n822 VDD.n821 9.3005
R5402 VDD.n1114 VDD.n1113 9.3005
R5403 VDD.n1115 VDD.n820 9.3005
R5404 VDD.n1117 VDD.n1116 9.3005
R5405 VDD.n810 VDD.n809 9.3005
R5406 VDD.n1130 VDD.n1129 9.3005
R5407 VDD.n1131 VDD.n808 9.3005
R5408 VDD.n1134 VDD.n1133 9.3005
R5409 VDD.n1132 VDD.n798 9.3005
R5410 VDD.n1067 VDD.n856 9.3005
R5411 VDD.n1648 VDD.t67 8.80749
R5412 VDD.n1746 VDD.t87 8.80749
R5413 VDD.n2138 VDD.t59 8.80749
R5414 VDD.n2271 VDD.t52 8.80749
R5415 VDD.t22 VDD.n617 8.51874
R5416 VDD.n1540 VDD.t13 8.51874
R5417 VDD.n2047 VDD.t8 8.51874
R5418 VDD.n442 VDD.t197 8.51874
R5419 VDD.n15 VDD.n14 8.32849
R5420 VDD.n2737 VDD.n2736 8.08725
R5421 VDD.n797 VDD.n796 8.08725
R5422 VDD.n1673 VDD.t28 7.79685
R5423 VDD.n2210 VDD.t198 7.79685
R5424 VDD.n842 VDD.t127 7.65248
R5425 VDD.n1192 VDD.t125 7.65248
R5426 VDD.t25 VDD.n629 7.65248
R5427 VDD.n585 VDD.t7 7.65248
R5428 VDD.t33 VDD.n475 7.65248
R5429 VDD.n430 VDD.t0 7.65248
R5430 VDD.n257 VDD.t154 7.65248
R5431 VDD.n2708 VDD.t145 7.65248
R5432 VDD.n818 VDD.t156 7.36372
R5433 VDD.n1160 VDD.t158 7.36372
R5434 VDD.n233 VDD.t139 7.36372
R5435 VDD.n2724 VDD.t123 7.36372
R5436 VDD.n2232 VDD.n2231 7.18099
R5437 VDD.n1652 VDD.n1651 7.18099
R5438 VDD.n1127 VDD.t156 7.07497
R5439 VDD.n764 VDD.t158 7.07497
R5440 VDD.n2546 VDD.t139 7.07497
R5441 VDD.t123 VDD.n55 7.07497
R5442 VDD.n1005 VDD.n1004 6.98232
R5443 VDD.n1326 VDD.n1273 6.98232
R5444 VDD.n2626 VDD.n162 6.98232
R5445 VDD.n2411 VDD.n2408 6.98232
R5446 VDD.n1685 VDD.t20 6.93059
R5447 VDD.n2198 VDD.t14 6.93059
R5448 VDD.n34 VDD.n24 6.82916
R5449 VDD.n785 VDD.n775 6.82916
R5450 VDD.n1095 VDD.t127 6.78621
R5451 VDD.n740 VDD.t125 6.78621
R5452 VDD.n2514 VDD.t154 6.78621
R5453 VDD.t145 VDD.n76 6.78621
R5454 VDD.n655 VDD.t48 6.64184
R5455 VDD.t103 VDD.n403 6.64184
R5456 VDD.n1697 VDD.t23 6.06433
R5457 VDD.n1815 VDD.t2 6.06433
R5458 VDD.n1873 VDD.t26 6.06433
R5459 VDD.n2186 VDD.t9 6.06433
R5460 VDD.n1766 VDD.n1765 5.77611
R5461 VDD.n1591 VDD.n684 5.77611
R5462 VDD.n1949 VDD.n1948 5.77611
R5463 VDD.n2289 VDD.n2288 5.77611
R5464 VDD.n366 VDD.n361 5.77611
R5465 VDD.n1889 VDD.n1885 5.77611
R5466 VDD.n1825 VDD.n542 5.77611
R5467 VDD.n1462 VDD.n1461 5.77611
R5468 VDD.n971 VDD.n968 5.62474
R5469 VDD.n1402 VDD.n707 5.62474
R5470 VDD.n2589 VDD.n201 5.62474
R5471 VDD.n2369 VDD.n2366 5.62474
R5472 VDD.n1727 VDD.t18 5.48682
R5473 VDD.n2156 VDD.t195 5.48682
R5474 VDD.n7 VDD.t15 5.418
R5475 VDD.n7 VDD.t199 5.418
R5476 VDD.n8 VDD.t38 5.418
R5477 VDD.n8 VDD.t10 5.418
R5478 VDD.n10 VDD.t12 5.418
R5479 VDD.n10 VDD.t196 5.418
R5480 VDD.n12 VDD.t6 5.418
R5481 VDD.n12 VDD.t27 5.418
R5482 VDD.n5 VDD.t3 5.418
R5483 VDD.n5 VDD.t17 5.418
R5484 VDD.n3 VDD.t19 5.418
R5485 VDD.n3 VDD.t31 5.418
R5486 VDD.n1 VDD.t24 5.418
R5487 VDD.n1 VDD.t35 5.418
R5488 VDD.n0 VDD.t29 5.418
R5489 VDD.n0 VDD.t21 5.418
R5490 VDD.n1611 VDD.n676 5.30782
R5491 VDD.n1607 VDD.n676 5.30782
R5492 VDD.n2308 VDD.n310 5.30782
R5493 VDD.n2304 VDD.n310 5.30782
R5494 VDD.n2357 VDD.n354 5.30782
R5495 VDD.n2357 VDD.n2356 5.30782
R5496 VDD.n1412 VDD.n1411 5.30782
R5497 VDD.n1444 VDD.n1411 5.30782
R5498 VDD.n1709 VDD.t34 5.19807
R5499 VDD.t30 VDD.n558 5.19807
R5500 VDD.t16 VDD.n1869 5.19807
R5501 VDD.n1870 VDD.t5 5.19807
R5502 VDD.n500 VDD.t11 5.19807
R5503 VDD.n2174 VDD.t37 5.19807
R5504 VDD.n1765 VDD.n1764 4.83952
R5505 VDD.n1587 VDD.n684 4.83952
R5506 VDD.n1950 VDD.n1949 4.83952
R5507 VDD.n2288 VDD.n2287 4.83952
R5508 VDD.n2337 VDD.n366 4.83952
R5509 VDD.n2076 VDD.n1889 4.83952
R5510 VDD.n1822 VDD.n542 4.83952
R5511 VDD.n1463 VDD.n1462 4.83952
R5512 VDD.n1303 VDD.n696 4.74817
R5513 VDD.n1299 VDD.n697 4.74817
R5514 VDD.n1386 VDD.n1385 4.74817
R5515 VDD.n1383 VDD.n1225 4.74817
R5516 VDD.n1385 VDD.n1223 4.74817
R5517 VDD.n1383 VDD.n1382 4.74817
R5518 VDD.n2474 VDD.n2473 4.74817
R5519 VDD.n2471 VDD.n2470 4.74817
R5520 VDD.n2471 VDD.n313 4.74817
R5521 VDD.n2473 VDD.n308 4.74817
R5522 VDD.n2381 VDD.n352 4.74817
R5523 VDD.n2379 VDD.n2378 4.74817
R5524 VDD.n2379 VDD.n2360 4.74817
R5525 VDD.n2382 VDD.n2381 4.74817
R5526 VDD.n1296 VDD.n696 4.74817
R5527 VDD.n699 VDD.n697 4.74817
R5528 VDD.n44 VDD.n43 4.7074
R5529 VDD.n34 VDD.n33 4.7074
R5530 VDD.n795 VDD.n794 4.7074
R5531 VDD.n785 VDD.n784 4.7074
R5532 VDD.n41 VDD.t170 4.64407
R5533 VDD.n41 VDD.t188 4.64407
R5534 VDD.n39 VDD.t176 4.64407
R5535 VDD.n39 VDD.t124 4.64407
R5536 VDD.n37 VDD.t140 4.64407
R5537 VDD.n37 VDD.t150 4.64407
R5538 VDD.n35 VDD.t118 4.64407
R5539 VDD.n35 VDD.t162 4.64407
R5540 VDD.n31 VDD.t116 4.64407
R5541 VDD.n31 VDD.t161 4.64407
R5542 VDD.n29 VDD.t131 4.64407
R5543 VDD.n29 VDD.t173 4.64407
R5544 VDD.n27 VDD.t181 4.64407
R5545 VDD.n27 VDD.t183 4.64407
R5546 VDD.n25 VDD.t171 4.64407
R5547 VDD.n25 VDD.t190 4.64407
R5548 VDD.n22 VDD.t175 4.64407
R5549 VDD.n22 VDD.t163 4.64407
R5550 VDD.n20 VDD.t151 4.64407
R5551 VDD.n20 VDD.t129 4.64407
R5552 VDD.n18 VDD.t166 4.64407
R5553 VDD.n18 VDD.t168 4.64407
R5554 VDD.n16 VDD.t164 4.64407
R5555 VDD.n16 VDD.t144 4.64407
R5556 VDD.n786 VDD.t178 4.64407
R5557 VDD.n786 VDD.t153 4.64407
R5558 VDD.n788 VDD.t172 4.64407
R5559 VDD.n788 VDD.t159 4.64407
R5560 VDD.n790 VDD.t157 4.64407
R5561 VDD.n790 VDD.t191 4.64407
R5562 VDD.n792 VDD.t133 4.64407
R5563 VDD.n792 VDD.t180 4.64407
R5564 VDD.n776 VDD.t138 4.64407
R5565 VDD.n776 VDD.t185 4.64407
R5566 VDD.n778 VDD.t122 4.64407
R5567 VDD.n778 VDD.t187 4.64407
R5568 VDD.n780 VDD.t186 4.64407
R5569 VDD.n780 VDD.t165 4.64407
R5570 VDD.n782 VDD.t177 4.64407
R5571 VDD.n782 VDD.t142 4.64407
R5572 VDD.n767 VDD.t193 4.64407
R5573 VDD.n767 VDD.t136 4.64407
R5574 VDD.n769 VDD.t148 4.64407
R5575 VDD.n769 VDD.t169 4.64407
R5576 VDD.n771 VDD.t189 4.64407
R5577 VDD.n771 VDD.t120 4.64407
R5578 VDD.n773 VDD.t134 4.64407
R5579 VDD.n773 VDD.t179 4.64407
R5580 VDD.n1540 VDD.t34 4.62056
R5581 VDD.n1739 VDD.t30 4.62056
R5582 VDD.n2144 VDD.t11 4.62056
R5583 VDD.n2047 VDD.t37 4.62056
R5584 VDD.n2737 VDD.n44 4.55156
R5585 VDD.n796 VDD.n795 4.55156
R5586 VDD.t40 VDD.n848 4.47618
R5587 VDD.n1209 VDD.t44 4.47618
R5588 VDD.t71 VDD.n263 4.47618
R5589 VDD.n2700 VDD.t63 4.47618
R5590 VDD.t18 VDD.n571 4.33181
R5591 VDD.n489 VDD.t195 4.33181
R5592 VDD.n1549 VDD.t23 3.7543
R5593 VDD.n1753 VDD.t2 3.7543
R5594 VDD.n2132 VDD.t26 3.7543
R5595 VDD.n2038 VDD.t9 3.7543
R5596 VDD.n2231 VDD.n2230 3.43465
R5597 VDD.n1653 VDD.n1652 3.43465
R5598 VDD.n1655 VDD.t48 3.17679
R5599 VDD.n2228 VDD.t103 3.17679
R5600 VDD.t20 VDD.n611 2.88804
R5601 VDD.n448 VDD.t14 2.88804
R5602 VDD.n1103 VDD.t132 2.74366
R5603 VDD.t135 VDD.n739 2.74366
R5604 VDD.n2522 VDD.t117 2.74366
R5605 VDD.t160 VDD.n2715 2.74366
R5606 VDD.n1136 VDD.t119 2.45491
R5607 VDD.t121 VDD.n763 2.45491
R5608 VDD.n2554 VDD.t149 2.45491
R5609 VDD.t130 VDD.n2731 2.45491
R5610 VDD.n1385 VDD.n1384 2.27742
R5611 VDD.n1384 VDD.n1383 2.27742
R5612 VDD.n2472 VDD.n2471 2.27742
R5613 VDD.n2473 VDD.n2472 2.27742
R5614 VDD.n2380 VDD.n2379 2.27742
R5615 VDD.n2381 VDD.n2380 2.27742
R5616 VDD.n1410 VDD.n696 2.27742
R5617 VDD.n1410 VDD.n697 2.27742
R5618 VDD.t141 VDD.n817 2.16615
R5619 VDD.n1168 VDD.t137 2.16615
R5620 VDD.n1667 VDD.t25 2.16615
R5621 VDD.n1727 VDD.t7 2.16615
R5622 VDD.n2156 VDD.t33 2.16615
R5623 VDD.n2216 VDD.t0 2.16615
R5624 VDD.t143 VDD.n232 2.16615
R5625 VDD.n2722 VDD.t115 2.16615
R5626 VDD.n44 VDD.n34 2.12227
R5627 VDD.n795 VDD.n785 2.12227
R5628 VDD.t28 VDD.n623 2.02178
R5629 VDD.n436 VDD.t198 2.02178
R5630 VDD.n1679 VDD.t22 1.29989
R5631 VDD.n1715 VDD.t13 1.29989
R5632 VDD.n2168 VDD.t8 1.29989
R5633 VDD.n2204 VDD.t197 1.29989
R5634 VDD.n662 VDD.t67 1.01114
R5635 VDD.t87 VDD.n554 1.01114
R5636 VDD.n506 VDD.t59 1.01114
R5637 VDD.t52 VDD.n397 1.01114
R5638 VDD.n972 VDD.n971 0.970197
R5639 VDD.n707 VDD.n703 0.970197
R5640 VDD.n201 VDD.n197 0.970197
R5641 VDD.n2371 VDD.n2369 0.970197
R5642 VDD.n796 VDD.n15 0.960867
R5643 VDD VDD.n2737 0.953033
R5644 VDD.n4 VDD.n2 0.728948
R5645 VDD.n11 VDD.n9 0.728948
R5646 VDD.n38 VDD.n36 0.573776
R5647 VDD.n40 VDD.n38 0.573776
R5648 VDD.n42 VDD.n40 0.573776
R5649 VDD.n43 VDD.n42 0.573776
R5650 VDD.n28 VDD.n26 0.573776
R5651 VDD.n30 VDD.n28 0.573776
R5652 VDD.n32 VDD.n30 0.573776
R5653 VDD.n33 VDD.n32 0.573776
R5654 VDD.n19 VDD.n17 0.573776
R5655 VDD.n21 VDD.n19 0.573776
R5656 VDD.n23 VDD.n21 0.573776
R5657 VDD.n24 VDD.n23 0.573776
R5658 VDD.n794 VDD.n793 0.573776
R5659 VDD.n793 VDD.n791 0.573776
R5660 VDD.n791 VDD.n789 0.573776
R5661 VDD.n789 VDD.n787 0.573776
R5662 VDD.n784 VDD.n783 0.573776
R5663 VDD.n783 VDD.n781 0.573776
R5664 VDD.n781 VDD.n779 0.573776
R5665 VDD.n779 VDD.n777 0.573776
R5666 VDD.n775 VDD.n774 0.573776
R5667 VDD.n774 VDD.n772 0.573776
R5668 VDD.n772 VDD.n770 0.573776
R5669 VDD.n770 VDD.n768 0.573776
R5670 VDD.n6 VDD.n4 0.573776
R5671 VDD.n13 VDD.n11 0.573776
R5672 VDD.n14 VDD.n6 0.49619
R5673 VDD.n14 VDD.n13 0.49619
R5674 VDD.n1396 VDD.n1395 0.471537
R5675 VDD.n2486 VDD.n2485 0.471537
R5676 VDD.n2695 VDD.n2694 0.471537
R5677 VDD.n2588 VDD.n2587 0.471537
R5678 VDD.n2365 VDD.n266 0.471537
R5679 VDD.n1403 VDD.n704 0.471537
R5680 VDD.n966 VDD.n851 0.471537
R5681 VDD.n1067 VDD.n1066 0.471537
R5682 VDD.n1691 VDD.t4 0.433631
R5683 VDD.n1703 VDD.t32 0.433631
R5684 VDD.n2180 VDD.t1 0.433631
R5685 VDD.n2192 VDD.t36 0.433631
R5686 VDD.n1229 VDD.n1224 0.152939
R5687 VDD.n1230 VDD.n1229 0.152939
R5688 VDD.n1234 VDD.n1230 0.152939
R5689 VDD.n1235 VDD.n1234 0.152939
R5690 VDD.n1236 VDD.n1235 0.152939
R5691 VDD.n1237 VDD.n1236 0.152939
R5692 VDD.n1244 VDD.n1237 0.152939
R5693 VDD.n1362 VDD.n1244 0.152939
R5694 VDD.n1362 VDD.n1361 0.152939
R5695 VDD.n1361 VDD.n1360 0.152939
R5696 VDD.n1360 VDD.n1245 0.152939
R5697 VDD.n1249 VDD.n1245 0.152939
R5698 VDD.n1250 VDD.n1249 0.152939
R5699 VDD.n1251 VDD.n1250 0.152939
R5700 VDD.n1255 VDD.n1251 0.152939
R5701 VDD.n1256 VDD.n1255 0.152939
R5702 VDD.n1257 VDD.n1256 0.152939
R5703 VDD.n1258 VDD.n1257 0.152939
R5704 VDD.n1262 VDD.n1258 0.152939
R5705 VDD.n1263 VDD.n1262 0.152939
R5706 VDD.n1264 VDD.n1263 0.152939
R5707 VDD.n1265 VDD.n1264 0.152939
R5708 VDD.n1269 VDD.n1265 0.152939
R5709 VDD.n1270 VDD.n1269 0.152939
R5710 VDD.n1271 VDD.n1270 0.152939
R5711 VDD.n1272 VDD.n1271 0.152939
R5712 VDD.n1279 VDD.n1272 0.152939
R5713 VDD.n1325 VDD.n1279 0.152939
R5714 VDD.n1325 VDD.n1324 0.152939
R5715 VDD.n1324 VDD.n1323 0.152939
R5716 VDD.n1323 VDD.n1280 0.152939
R5717 VDD.n1284 VDD.n1280 0.152939
R5718 VDD.n1285 VDD.n1284 0.152939
R5719 VDD.n1286 VDD.n1285 0.152939
R5720 VDD.n1290 VDD.n1286 0.152939
R5721 VDD.n1291 VDD.n1290 0.152939
R5722 VDD.n1292 VDD.n1291 0.152939
R5723 VDD.n1293 VDD.n1292 0.152939
R5724 VDD.n1293 VDD.n695 0.152939
R5725 VDD.n1395 VDD.n1214 0.152939
R5726 VDD.n1218 VDD.n1214 0.152939
R5727 VDD.n1219 VDD.n1218 0.152939
R5728 VDD.n1220 VDD.n1219 0.152939
R5729 VDD.n1148 VDD.n1147 0.152939
R5730 VDD.n1149 VDD.n1148 0.152939
R5731 VDD.n1149 VDD.n755 0.152939
R5732 VDD.n1163 VDD.n755 0.152939
R5733 VDD.n1164 VDD.n1163 0.152939
R5734 VDD.n1165 VDD.n1164 0.152939
R5735 VDD.n1165 VDD.n743 0.152939
R5736 VDD.n1179 VDD.n743 0.152939
R5737 VDD.n1180 VDD.n1179 0.152939
R5738 VDD.n1181 VDD.n1180 0.152939
R5739 VDD.n1181 VDD.n731 0.152939
R5740 VDD.n1195 VDD.n731 0.152939
R5741 VDD.n1196 VDD.n1195 0.152939
R5742 VDD.n1197 VDD.n1196 0.152939
R5743 VDD.n1197 VDD.n718 0.152939
R5744 VDD.n1212 VDD.n718 0.152939
R5745 VDD.n1213 VDD.n1212 0.152939
R5746 VDD.n1396 VDD.n1213 0.152939
R5747 VDD.n315 VDD.n309 0.152939
R5748 VDD.n316 VDD.n315 0.152939
R5749 VDD.n317 VDD.n316 0.152939
R5750 VDD.n318 VDD.n317 0.152939
R5751 VDD.n319 VDD.n318 0.152939
R5752 VDD.n320 VDD.n319 0.152939
R5753 VDD.n321 VDD.n320 0.152939
R5754 VDD.n2449 VDD.n321 0.152939
R5755 VDD.n2449 VDD.n2448 0.152939
R5756 VDD.n2448 VDD.n2447 0.152939
R5757 VDD.n2447 VDD.n323 0.152939
R5758 VDD.n324 VDD.n323 0.152939
R5759 VDD.n325 VDD.n324 0.152939
R5760 VDD.n326 VDD.n325 0.152939
R5761 VDD.n327 VDD.n326 0.152939
R5762 VDD.n328 VDD.n327 0.152939
R5763 VDD.n329 VDD.n328 0.152939
R5764 VDD.n330 VDD.n329 0.152939
R5765 VDD.n331 VDD.n330 0.152939
R5766 VDD.n332 VDD.n331 0.152939
R5767 VDD.n333 VDD.n332 0.152939
R5768 VDD.n334 VDD.n333 0.152939
R5769 VDD.n335 VDD.n334 0.152939
R5770 VDD.n336 VDD.n335 0.152939
R5771 VDD.n337 VDD.n336 0.152939
R5772 VDD.n338 VDD.n337 0.152939
R5773 VDD.n339 VDD.n338 0.152939
R5774 VDD.n2407 VDD.n339 0.152939
R5775 VDD.n2407 VDD.n2406 0.152939
R5776 VDD.n2406 VDD.n2405 0.152939
R5777 VDD.n2405 VDD.n343 0.152939
R5778 VDD.n344 VDD.n343 0.152939
R5779 VDD.n345 VDD.n344 0.152939
R5780 VDD.n346 VDD.n345 0.152939
R5781 VDD.n347 VDD.n346 0.152939
R5782 VDD.n348 VDD.n347 0.152939
R5783 VDD.n349 VDD.n348 0.152939
R5784 VDD.n350 VDD.n349 0.152939
R5785 VDD.n351 VDD.n350 0.152939
R5786 VDD.n2485 VDD.n272 0.152939
R5787 VDD.n305 VDD.n272 0.152939
R5788 VDD.n306 VDD.n305 0.152939
R5789 VDD.n307 VDD.n306 0.152939
R5790 VDD.n2487 VDD.n2486 0.152939
R5791 VDD.n2487 VDD.n260 0.152939
R5792 VDD.n2501 VDD.n260 0.152939
R5793 VDD.n2502 VDD.n2501 0.152939
R5794 VDD.n2503 VDD.n2502 0.152939
R5795 VDD.n2503 VDD.n248 0.152939
R5796 VDD.n2517 VDD.n248 0.152939
R5797 VDD.n2518 VDD.n2517 0.152939
R5798 VDD.n2519 VDD.n2518 0.152939
R5799 VDD.n2519 VDD.n236 0.152939
R5800 VDD.n2533 VDD.n236 0.152939
R5801 VDD.n2534 VDD.n2533 0.152939
R5802 VDD.n2535 VDD.n2534 0.152939
R5803 VDD.n2535 VDD.n224 0.152939
R5804 VDD.n2549 VDD.n224 0.152939
R5805 VDD.n2550 VDD.n2549 0.152939
R5806 VDD.n2551 VDD.n2550 0.152939
R5807 VDD.n2551 VDD.n45 0.152939
R5808 VDD.n2735 VDD.n46 0.152939
R5809 VDD.n57 VDD.n46 0.152939
R5810 VDD.n58 VDD.n57 0.152939
R5811 VDD.n59 VDD.n58 0.152939
R5812 VDD.n66 VDD.n59 0.152939
R5813 VDD.n67 VDD.n66 0.152939
R5814 VDD.n68 VDD.n67 0.152939
R5815 VDD.n69 VDD.n68 0.152939
R5816 VDD.n78 VDD.n69 0.152939
R5817 VDD.n79 VDD.n78 0.152939
R5818 VDD.n80 VDD.n79 0.152939
R5819 VDD.n81 VDD.n80 0.152939
R5820 VDD.n89 VDD.n81 0.152939
R5821 VDD.n90 VDD.n89 0.152939
R5822 VDD.n91 VDD.n90 0.152939
R5823 VDD.n92 VDD.n91 0.152939
R5824 VDD.n100 VDD.n92 0.152939
R5825 VDD.n2695 VDD.n100 0.152939
R5826 VDD.n2694 VDD.n101 0.152939
R5827 VDD.n104 VDD.n101 0.152939
R5828 VDD.n108 VDD.n104 0.152939
R5829 VDD.n109 VDD.n108 0.152939
R5830 VDD.n110 VDD.n109 0.152939
R5831 VDD.n111 VDD.n110 0.152939
R5832 VDD.n112 VDD.n111 0.152939
R5833 VDD.n116 VDD.n112 0.152939
R5834 VDD.n117 VDD.n116 0.152939
R5835 VDD.n118 VDD.n117 0.152939
R5836 VDD.n119 VDD.n118 0.152939
R5837 VDD.n123 VDD.n119 0.152939
R5838 VDD.n124 VDD.n123 0.152939
R5839 VDD.n125 VDD.n124 0.152939
R5840 VDD.n126 VDD.n125 0.152939
R5841 VDD.n133 VDD.n126 0.152939
R5842 VDD.n2662 VDD.n133 0.152939
R5843 VDD.n2662 VDD.n2661 0.152939
R5844 VDD.n2661 VDD.n2660 0.152939
R5845 VDD.n2660 VDD.n134 0.152939
R5846 VDD.n138 VDD.n134 0.152939
R5847 VDD.n139 VDD.n138 0.152939
R5848 VDD.n140 VDD.n139 0.152939
R5849 VDD.n144 VDD.n140 0.152939
R5850 VDD.n145 VDD.n144 0.152939
R5851 VDD.n146 VDD.n145 0.152939
R5852 VDD.n147 VDD.n146 0.152939
R5853 VDD.n151 VDD.n147 0.152939
R5854 VDD.n152 VDD.n151 0.152939
R5855 VDD.n153 VDD.n152 0.152939
R5856 VDD.n154 VDD.n153 0.152939
R5857 VDD.n158 VDD.n154 0.152939
R5858 VDD.n159 VDD.n158 0.152939
R5859 VDD.n160 VDD.n159 0.152939
R5860 VDD.n161 VDD.n160 0.152939
R5861 VDD.n168 VDD.n161 0.152939
R5862 VDD.n2625 VDD.n168 0.152939
R5863 VDD.n2625 VDD.n2624 0.152939
R5864 VDD.n2624 VDD.n2623 0.152939
R5865 VDD.n2623 VDD.n169 0.152939
R5866 VDD.n173 VDD.n169 0.152939
R5867 VDD.n174 VDD.n173 0.152939
R5868 VDD.n175 VDD.n174 0.152939
R5869 VDD.n179 VDD.n175 0.152939
R5870 VDD.n180 VDD.n179 0.152939
R5871 VDD.n181 VDD.n180 0.152939
R5872 VDD.n182 VDD.n181 0.152939
R5873 VDD.n186 VDD.n182 0.152939
R5874 VDD.n187 VDD.n186 0.152939
R5875 VDD.n188 VDD.n187 0.152939
R5876 VDD.n189 VDD.n188 0.152939
R5877 VDD.n193 VDD.n189 0.152939
R5878 VDD.n194 VDD.n193 0.152939
R5879 VDD.n195 VDD.n194 0.152939
R5880 VDD.n196 VDD.n195 0.152939
R5881 VDD.n202 VDD.n196 0.152939
R5882 VDD.n2588 VDD.n202 0.152939
R5883 VDD.n2493 VDD.n266 0.152939
R5884 VDD.n2494 VDD.n2493 0.152939
R5885 VDD.n2495 VDD.n2494 0.152939
R5886 VDD.n2495 VDD.n253 0.152939
R5887 VDD.n2509 VDD.n253 0.152939
R5888 VDD.n2510 VDD.n2509 0.152939
R5889 VDD.n2511 VDD.n2510 0.152939
R5890 VDD.n2511 VDD.n242 0.152939
R5891 VDD.n2525 VDD.n242 0.152939
R5892 VDD.n2526 VDD.n2525 0.152939
R5893 VDD.n2527 VDD.n2526 0.152939
R5894 VDD.n2527 VDD.n229 0.152939
R5895 VDD.n2541 VDD.n229 0.152939
R5896 VDD.n2542 VDD.n2541 0.152939
R5897 VDD.n2543 VDD.n2542 0.152939
R5898 VDD.n2543 VDD.n217 0.152939
R5899 VDD.n2557 VDD.n217 0.152939
R5900 VDD.n2558 VDD.n2557 0.152939
R5901 VDD.n2559 VDD.n2558 0.152939
R5902 VDD.n2559 VDD.n215 0.152939
R5903 VDD.n2563 VDD.n215 0.152939
R5904 VDD.n2564 VDD.n2563 0.152939
R5905 VDD.n2565 VDD.n2564 0.152939
R5906 VDD.n2565 VDD.n212 0.152939
R5907 VDD.n2569 VDD.n212 0.152939
R5908 VDD.n2570 VDD.n2569 0.152939
R5909 VDD.n2571 VDD.n2570 0.152939
R5910 VDD.n2571 VDD.n209 0.152939
R5911 VDD.n2575 VDD.n209 0.152939
R5912 VDD.n2576 VDD.n2575 0.152939
R5913 VDD.n2577 VDD.n2576 0.152939
R5914 VDD.n2577 VDD.n206 0.152939
R5915 VDD.n2581 VDD.n206 0.152939
R5916 VDD.n2582 VDD.n2581 0.152939
R5917 VDD.n2583 VDD.n2582 0.152939
R5918 VDD.n2583 VDD.n203 0.152939
R5919 VDD.n2587 VDD.n203 0.152939
R5920 VDD.n2362 VDD.n353 0.152939
R5921 VDD.n2363 VDD.n2362 0.152939
R5922 VDD.n2364 VDD.n2363 0.152939
R5923 VDD.n2365 VDD.n2364 0.152939
R5924 VDD.n1409 VDD.n698 0.152939
R5925 VDD.n1405 VDD.n698 0.152939
R5926 VDD.n1405 VDD.n1404 0.152939
R5927 VDD.n1404 VDD.n1403 0.152939
R5928 VDD.n1074 VDD.n851 0.152939
R5929 VDD.n1075 VDD.n1074 0.152939
R5930 VDD.n1076 VDD.n1075 0.152939
R5931 VDD.n1076 VDD.n838 0.152939
R5932 VDD.n1090 VDD.n838 0.152939
R5933 VDD.n1091 VDD.n1090 0.152939
R5934 VDD.n1092 VDD.n1091 0.152939
R5935 VDD.n1092 VDD.n827 0.152939
R5936 VDD.n1106 VDD.n827 0.152939
R5937 VDD.n1107 VDD.n1106 0.152939
R5938 VDD.n1108 VDD.n1107 0.152939
R5939 VDD.n1108 VDD.n814 0.152939
R5940 VDD.n1122 VDD.n814 0.152939
R5941 VDD.n1123 VDD.n1122 0.152939
R5942 VDD.n1124 VDD.n1123 0.152939
R5943 VDD.n1124 VDD.n803 0.152939
R5944 VDD.n1139 VDD.n803 0.152939
R5945 VDD.n1140 VDD.n1139 0.152939
R5946 VDD.n1141 VDD.n1140 0.152939
R5947 VDD.n1141 VDD.n760 0.152939
R5948 VDD.n1155 VDD.n760 0.152939
R5949 VDD.n1156 VDD.n1155 0.152939
R5950 VDD.n1157 VDD.n1156 0.152939
R5951 VDD.n1157 VDD.n749 0.152939
R5952 VDD.n1171 VDD.n749 0.152939
R5953 VDD.n1172 VDD.n1171 0.152939
R5954 VDD.n1173 VDD.n1172 0.152939
R5955 VDD.n1173 VDD.n736 0.152939
R5956 VDD.n1187 VDD.n736 0.152939
R5957 VDD.n1188 VDD.n1187 0.152939
R5958 VDD.n1189 VDD.n1188 0.152939
R5959 VDD.n1189 VDD.n725 0.152939
R5960 VDD.n1203 VDD.n725 0.152939
R5961 VDD.n1204 VDD.n1203 0.152939
R5962 VDD.n1206 VDD.n1204 0.152939
R5963 VDD.n1206 VDD.n1205 0.152939
R5964 VDD.n1205 VDD.n704 0.152939
R5965 VDD.n1066 VDD.n857 0.152939
R5966 VDD.n1059 VDD.n857 0.152939
R5967 VDD.n1059 VDD.n1058 0.152939
R5968 VDD.n1058 VDD.n1057 0.152939
R5969 VDD.n1057 VDD.n890 0.152939
R5970 VDD.n1053 VDD.n890 0.152939
R5971 VDD.n1053 VDD.n1052 0.152939
R5972 VDD.n1052 VDD.n1051 0.152939
R5973 VDD.n1051 VDD.n896 0.152939
R5974 VDD.n1047 VDD.n896 0.152939
R5975 VDD.n1047 VDD.n1046 0.152939
R5976 VDD.n1046 VDD.n1045 0.152939
R5977 VDD.n1045 VDD.n902 0.152939
R5978 VDD.n1041 VDD.n902 0.152939
R5979 VDD.n1041 VDD.n1040 0.152939
R5980 VDD.n1040 VDD.n1039 0.152939
R5981 VDD.n1039 VDD.n908 0.152939
R5982 VDD.n1032 VDD.n908 0.152939
R5983 VDD.n1032 VDD.n1031 0.152939
R5984 VDD.n1031 VDD.n1030 0.152939
R5985 VDD.n1030 VDD.n913 0.152939
R5986 VDD.n1026 VDD.n913 0.152939
R5987 VDD.n1026 VDD.n1025 0.152939
R5988 VDD.n1025 VDD.n1024 0.152939
R5989 VDD.n1024 VDD.n919 0.152939
R5990 VDD.n1020 VDD.n919 0.152939
R5991 VDD.n1020 VDD.n1019 0.152939
R5992 VDD.n1019 VDD.n1018 0.152939
R5993 VDD.n1018 VDD.n925 0.152939
R5994 VDD.n1014 VDD.n925 0.152939
R5995 VDD.n1014 VDD.n1013 0.152939
R5996 VDD.n1013 VDD.n1012 0.152939
R5997 VDD.n1012 VDD.n931 0.152939
R5998 VDD.n1008 VDD.n931 0.152939
R5999 VDD.n1008 VDD.n1007 0.152939
R6000 VDD.n1007 VDD.n1006 0.152939
R6001 VDD.n1006 VDD.n937 0.152939
R6002 VDD.n999 VDD.n937 0.152939
R6003 VDD.n999 VDD.n998 0.152939
R6004 VDD.n998 VDD.n997 0.152939
R6005 VDD.n997 VDD.n942 0.152939
R6006 VDD.n993 VDD.n942 0.152939
R6007 VDD.n993 VDD.n992 0.152939
R6008 VDD.n992 VDD.n991 0.152939
R6009 VDD.n991 VDD.n948 0.152939
R6010 VDD.n987 VDD.n948 0.152939
R6011 VDD.n987 VDD.n986 0.152939
R6012 VDD.n986 VDD.n985 0.152939
R6013 VDD.n985 VDD.n954 0.152939
R6014 VDD.n981 VDD.n954 0.152939
R6015 VDD.n981 VDD.n980 0.152939
R6016 VDD.n980 VDD.n979 0.152939
R6017 VDD.n979 VDD.n960 0.152939
R6018 VDD.n975 VDD.n960 0.152939
R6019 VDD.n975 VDD.n974 0.152939
R6020 VDD.n974 VDD.n973 0.152939
R6021 VDD.n973 VDD.n966 0.152939
R6022 VDD.n1068 VDD.n1067 0.152939
R6023 VDD.n1068 VDD.n845 0.152939
R6024 VDD.n1082 VDD.n845 0.152939
R6025 VDD.n1083 VDD.n1082 0.152939
R6026 VDD.n1084 VDD.n1083 0.152939
R6027 VDD.n1084 VDD.n833 0.152939
R6028 VDD.n1098 VDD.n833 0.152939
R6029 VDD.n1099 VDD.n1098 0.152939
R6030 VDD.n1100 VDD.n1099 0.152939
R6031 VDD.n1100 VDD.n821 0.152939
R6032 VDD.n1114 VDD.n821 0.152939
R6033 VDD.n1115 VDD.n1114 0.152939
R6034 VDD.n1116 VDD.n1115 0.152939
R6035 VDD.n1116 VDD.n809 0.152939
R6036 VDD.n1130 VDD.n809 0.152939
R6037 VDD.n1131 VDD.n1130 0.152939
R6038 VDD.n1133 VDD.n1131 0.152939
R6039 VDD.n1133 VDD.n1132 0.152939
R6040 VDD.n1384 VDD.n1220 0.110256
R6041 VDD.n2472 VDD.n307 0.110256
R6042 VDD.n2380 VDD.n353 0.110256
R6043 VDD.n1410 VDD.n1409 0.110256
R6044 VDD.n1147 VDD.n797 0.0695946
R6045 VDD.n2736 VDD.n45 0.0695946
R6046 VDD.n2736 VDD.n2735 0.0695946
R6047 VDD.n1132 VDD.n797 0.0695946
R6048 VDD.n1384 VDD.n1224 0.0431829
R6049 VDD.n1410 VDD.n695 0.0431829
R6050 VDD.n2472 VDD.n309 0.0431829
R6051 VDD.n2380 VDD.n351 0.0431829
R6052 VDD VDD.n15 0.00833333
R6053 a_n2686_12778.n115 a_n2686_12778.n95 756.745
R6054 a_n2686_12778.n86 a_n2686_12778.n66 756.745
R6055 a_n2686_12778.n163 a_n2686_12778.n143 756.745
R6056 a_n2686_12778.n192 a_n2686_12778.n172 756.745
R6057 a_n2686_12778.n116 a_n2686_12778.n115 585
R6058 a_n2686_12778.n114 a_n2686_12778.n113 585
R6059 a_n2686_12778.n98 a_n2686_12778.n97 585
R6060 a_n2686_12778.n110 a_n2686_12778.n109 585
R6061 a_n2686_12778.n108 a_n2686_12778.n107 585
R6062 a_n2686_12778.n101 a_n2686_12778.n100 585
R6063 a_n2686_12778.n104 a_n2686_12778.n103 585
R6064 a_n2686_12778.n87 a_n2686_12778.n86 585
R6065 a_n2686_12778.n85 a_n2686_12778.n84 585
R6066 a_n2686_12778.n69 a_n2686_12778.n68 585
R6067 a_n2686_12778.n81 a_n2686_12778.n80 585
R6068 a_n2686_12778.n79 a_n2686_12778.n78 585
R6069 a_n2686_12778.n72 a_n2686_12778.n71 585
R6070 a_n2686_12778.n75 a_n2686_12778.n74 585
R6071 a_n2686_12778.n164 a_n2686_12778.n163 585
R6072 a_n2686_12778.n162 a_n2686_12778.n161 585
R6073 a_n2686_12778.n146 a_n2686_12778.n145 585
R6074 a_n2686_12778.n158 a_n2686_12778.n157 585
R6075 a_n2686_12778.n156 a_n2686_12778.n155 585
R6076 a_n2686_12778.n149 a_n2686_12778.n148 585
R6077 a_n2686_12778.n152 a_n2686_12778.n151 585
R6078 a_n2686_12778.n193 a_n2686_12778.n192 585
R6079 a_n2686_12778.n191 a_n2686_12778.n190 585
R6080 a_n2686_12778.n175 a_n2686_12778.n174 585
R6081 a_n2686_12778.n187 a_n2686_12778.n186 585
R6082 a_n2686_12778.n185 a_n2686_12778.n184 585
R6083 a_n2686_12778.n178 a_n2686_12778.n177 585
R6084 a_n2686_12778.n181 a_n2686_12778.n180 585
R6085 a_n2686_12778.t24 a_n2686_12778.n102 327.601
R6086 a_n2686_12778.t22 a_n2686_12778.n73 327.601
R6087 a_n2686_12778.t12 a_n2686_12778.n150 327.601
R6088 a_n2686_12778.t16 a_n2686_12778.n179 327.601
R6089 a_n2686_12778.n141 a_n2686_12778.t15 183.883
R6090 a_n2686_12778.n133 a_n2686_12778.t11 183.883
R6091 a_n2686_12778.n225 a_n2686_12778.t53 183.883
R6092 a_n2686_12778.n230 a_n2686_12778.t44 183.883
R6093 a_n2686_12778.n217 a_n2686_12778.t45 183.883
R6094 a_n2686_12778.n222 a_n2686_12778.t36 183.883
R6095 a_n2686_12778.n209 a_n2686_12778.t58 183.883
R6096 a_n2686_12778.n214 a_n2686_12778.t39 183.883
R6097 a_n2686_12778.n201 a_n2686_12778.t33 183.883
R6098 a_n2686_12778.n206 a_n2686_12778.t42 183.883
R6099 a_n2686_12778.n10 a_n2686_12778.t21 206.089
R6100 a_n2686_12778.n8 a_n2686_12778.t49 206.089
R6101 a_n2686_12778.n12 a_n2686_12778.t37 206.089
R6102 a_n2686_12778.n115 a_n2686_12778.n114 171.744
R6103 a_n2686_12778.n114 a_n2686_12778.n97 171.744
R6104 a_n2686_12778.n109 a_n2686_12778.n97 171.744
R6105 a_n2686_12778.n109 a_n2686_12778.n108 171.744
R6106 a_n2686_12778.n108 a_n2686_12778.n100 171.744
R6107 a_n2686_12778.n103 a_n2686_12778.n100 171.744
R6108 a_n2686_12778.n86 a_n2686_12778.n85 171.744
R6109 a_n2686_12778.n85 a_n2686_12778.n68 171.744
R6110 a_n2686_12778.n80 a_n2686_12778.n68 171.744
R6111 a_n2686_12778.n80 a_n2686_12778.n79 171.744
R6112 a_n2686_12778.n79 a_n2686_12778.n71 171.744
R6113 a_n2686_12778.n74 a_n2686_12778.n71 171.744
R6114 a_n2686_12778.n163 a_n2686_12778.n162 171.744
R6115 a_n2686_12778.n162 a_n2686_12778.n145 171.744
R6116 a_n2686_12778.n157 a_n2686_12778.n145 171.744
R6117 a_n2686_12778.n157 a_n2686_12778.n156 171.744
R6118 a_n2686_12778.n156 a_n2686_12778.n148 171.744
R6119 a_n2686_12778.n151 a_n2686_12778.n148 171.744
R6120 a_n2686_12778.n192 a_n2686_12778.n191 171.744
R6121 a_n2686_12778.n191 a_n2686_12778.n174 171.744
R6122 a_n2686_12778.n186 a_n2686_12778.n174 171.744
R6123 a_n2686_12778.n186 a_n2686_12778.n185 171.744
R6124 a_n2686_12778.n185 a_n2686_12778.n177 171.744
R6125 a_n2686_12778.n180 a_n2686_12778.n177 171.744
R6126 a_n2686_12778.n17 a_n2686_12778.n5 68.6201
R6127 a_n2686_12778.n5 a_n2686_12778.n16 71.6402
R6128 a_n2686_12778.n129 a_n2686_12778.n7 161.3
R6129 a_n2686_12778.n7 a_n2686_12778.n15 68.6201
R6130 a_n2686_12778.n19 a_n2686_12778.n3 68.6201
R6131 a_n2686_12778.n3 a_n2686_12778.n18 71.6402
R6132 a_n2686_12778.n126 a_n2686_12778.n9 161.3
R6133 a_n2686_12778.n9 a_n2686_12778.n14 68.6201
R6134 a_n2686_12778.n21 a_n2686_12778.n0 68.6201
R6135 a_n2686_12778.n0 a_n2686_12778.n20 71.6402
R6136 a_n2686_12778.n234 a_n2686_12778.n11 161.3
R6137 a_n2686_12778.n11 a_n2686_12778.n13 68.6201
R6138 a_n2686_12778.n205 a_n2686_12778.n26 161.3
R6139 a_n2686_12778.n22 a_n2686_12778.n26 161.3
R6140 a_n2686_12778.n25 a_n2686_12778.n23 71.6402
R6141 a_n2686_12778.n202 a_n2686_12778.n24 161.3
R6142 a_n2686_12778.n213 a_n2686_12778.n31 161.3
R6143 a_n2686_12778.n27 a_n2686_12778.n31 161.3
R6144 a_n2686_12778.n30 a_n2686_12778.n28 71.6402
R6145 a_n2686_12778.n210 a_n2686_12778.n29 161.3
R6146 a_n2686_12778.n221 a_n2686_12778.n36 161.3
R6147 a_n2686_12778.n32 a_n2686_12778.n36 161.3
R6148 a_n2686_12778.n35 a_n2686_12778.n33 71.6402
R6149 a_n2686_12778.n218 a_n2686_12778.n34 161.3
R6150 a_n2686_12778.n229 a_n2686_12778.n41 161.3
R6151 a_n2686_12778.n37 a_n2686_12778.n41 161.3
R6152 a_n2686_12778.n40 a_n2686_12778.n38 71.6402
R6153 a_n2686_12778.n226 a_n2686_12778.n39 161.3
R6154 a_n2686_12778.n51 a_n2686_12778.n48 74.8341
R6155 a_n2686_12778.n49 a_n2686_12778.n46 68.6201
R6156 a_n2686_12778.n45 a_n2686_12778.n47 71.6402
R6157 a_n2686_12778.n135 a_n2686_12778.n42 161.3
R6158 a_n2686_12778.n137 a_n2686_12778.n42 161.3
R6159 a_n2686_12778.n44 a_n2686_12778.n138 161.3
R6160 a_n2686_12778.n139 a_n2686_12778.n44 161.3
R6161 a_n2686_12778.n140 a_n2686_12778.n43 161.3
R6162 a_n2686_12778.n131 a_n2686_12778.t27 144.601
R6163 a_n2686_12778.n136 a_n2686_12778.t7 144.601
R6164 a_n2686_12778.n134 a_n2686_12778.t29 144.601
R6165 a_n2686_12778.n132 a_n2686_12778.t9 144.601
R6166 a_n2686_12778.n227 a_n2686_12778.t38 144.601
R6167 a_n2686_12778.n228 a_n2686_12778.t56 144.601
R6168 a_n2686_12778.n219 a_n2686_12778.t55 144.601
R6169 a_n2686_12778.n220 a_n2686_12778.t52 144.601
R6170 a_n2686_12778.n211 a_n2686_12778.t47 144.601
R6171 a_n2686_12778.n212 a_n2686_12778.t51 144.601
R6172 a_n2686_12778.n203 a_n2686_12778.t50 144.601
R6173 a_n2686_12778.n204 a_n2686_12778.t59 144.601
R6174 a_n2686_12778.n123 a_n2686_12778.t19 144.601
R6175 a_n2686_12778.n127 a_n2686_12778.t17 144.601
R6176 a_n2686_12778.n125 a_n2686_12778.t25 144.601
R6177 a_n2686_12778.n124 a_n2686_12778.t13 144.601
R6178 a_n2686_12778.n121 a_n2686_12778.t54 144.601
R6179 a_n2686_12778.n130 a_n2686_12778.t32 144.601
R6180 a_n2686_12778.n128 a_n2686_12778.t48 144.601
R6181 a_n2686_12778.n122 a_n2686_12778.t57 144.601
R6182 a_n2686_12778.n64 a_n2686_12778.t46 144.601
R6183 a_n2686_12778.n235 a_n2686_12778.t43 144.601
R6184 a_n2686_12778.n233 a_n2686_12778.t34 144.601
R6185 a_n2686_12778.n65 a_n2686_12778.t41 144.601
R6186 a_n2686_12778.n103 a_n2686_12778.t24 85.8723
R6187 a_n2686_12778.n74 a_n2686_12778.t22 85.8723
R6188 a_n2686_12778.n151 a_n2686_12778.t12 85.8723
R6189 a_n2686_12778.n180 a_n2686_12778.t16 85.8723
R6190 a_n2686_12778.n94 a_n2686_12778.n93 81.2397
R6191 a_n2686_12778.n92 a_n2686_12778.n91 81.2397
R6192 a_n2686_12778.n169 a_n2686_12778.n168 81.2397
R6193 a_n2686_12778.n171 a_n2686_12778.n170 81.2397
R6194 a_n2686_12778.n239 a_n2686_12778.n238 81.219
R6195 a_n2686_12778.n239 a_n2686_12778.n237 81.219
R6196 a_n2686_12778.n243 a_n2686_12778.n242 81.219
R6197 a_n2686_12778.n241 a_n2686_12778.n240 80.9324
R6198 a_n2686_12778.n6 a_n2686_12778.n5 28.1161
R6199 a_n2686_12778.n7 a_n2686_12778.n8 28.1161
R6200 a_n2686_12778.n4 a_n2686_12778.n3 28.1161
R6201 a_n2686_12778.n9 a_n2686_12778.n10 28.1161
R6202 a_n2686_12778.n1 a_n2686_12778.n0 28.1161
R6203 a_n2686_12778.n11 a_n2686_12778.n12 28.1161
R6204 a_n2686_12778.n207 a_n2686_12778.n206 80.6037
R6205 a_n2686_12778.n201 a_n2686_12778.n200 80.6037
R6206 a_n2686_12778.n215 a_n2686_12778.n214 80.6037
R6207 a_n2686_12778.n209 a_n2686_12778.n208 80.6037
R6208 a_n2686_12778.n223 a_n2686_12778.n222 80.6037
R6209 a_n2686_12778.n217 a_n2686_12778.n216 80.6037
R6210 a_n2686_12778.n231 a_n2686_12778.n230 80.6037
R6211 a_n2686_12778.n225 a_n2686_12778.n224 80.6037
R6212 a_n2686_12778.n133 a_n2686_12778.n50 80.6037
R6213 a_n2686_12778.n142 a_n2686_12778.n141 80.6037
R6214 a_n2686_12778.n138 a_n2686_12778.n137 56.5617
R6215 a_n2686_12778.n49 a_n2686_12778.n132 48.4088
R6216 a_n2686_12778.n19 a_n2686_12778.n124 48.4088
R6217 a_n2686_12778.n17 a_n2686_12778.n122 48.4088
R6218 a_n2686_12778.n21 a_n2686_12778.n65 48.4088
R6219 a_n2686_12778.n226 a_n2686_12778.n225 56.3158
R6220 a_n2686_12778.n230 a_n2686_12778.n229 56.3158
R6221 a_n2686_12778.n218 a_n2686_12778.n217 56.3158
R6222 a_n2686_12778.n222 a_n2686_12778.n221 56.3158
R6223 a_n2686_12778.n210 a_n2686_12778.n209 56.3158
R6224 a_n2686_12778.n214 a_n2686_12778.n213 56.3158
R6225 a_n2686_12778.n202 a_n2686_12778.n201 56.3158
R6226 a_n2686_12778.n206 a_n2686_12778.n205 56.3158
R6227 a_n2686_12778.n141 a_n2686_12778.n140 47.4702
R6228 a_n2686_12778.n135 a_n2686_12778.n47 58.5991
R6229 a_n2686_12778.n134 a_n2686_12778.n47 26.1378
R6230 a_n2686_12778.n38 a_n2686_12778.n37 58.5991
R6231 a_n2686_12778.n33 a_n2686_12778.n32 58.5991
R6232 a_n2686_12778.n28 a_n2686_12778.n27 58.5991
R6233 a_n2686_12778.n23 a_n2686_12778.n22 58.5991
R6234 a_n2686_12778.n126 a_n2686_12778.n18 58.5991
R6235 a_n2686_12778.n125 a_n2686_12778.n18 26.1378
R6236 a_n2686_12778.n129 a_n2686_12778.n16 58.5991
R6237 a_n2686_12778.n128 a_n2686_12778.n16 26.1378
R6238 a_n2686_12778.n234 a_n2686_12778.n20 58.5991
R6239 a_n2686_12778.n233 a_n2686_12778.n20 26.1378
R6240 a_n2686_12778.n92 a_n2686_12778.n90 38.3829
R6241 a_n2686_12778.n169 a_n2686_12778.n167 38.3829
R6242 a_n2686_12778.n120 a_n2686_12778.n119 37.8096
R6243 a_n2686_12778.n197 a_n2686_12778.n196 37.8096
R6244 a_n2686_12778.n241 a_n2686_12778.n239 30.598
R6245 a_n2686_12778.n140 a_n2686_12778.n139 25.0767
R6246 a_n2686_12778.n51 a_n2686_12778.n133 59.1045
R6247 a_n2686_12778.n10 a_n2686_12778.n123 32.4972
R6248 a_n2686_12778.n4 a_n2686_12778.t23 206.089
R6249 a_n2686_12778.n8 a_n2686_12778.n121 32.4972
R6250 a_n2686_12778.n6 a_n2686_12778.t35 206.089
R6251 a_n2686_12778.n12 a_n2686_12778.n64 32.4972
R6252 a_n2686_12778.n1 a_n2686_12778.t40 206.089
R6253 a_n2686_12778.n138 a_n2686_12778.n131 24.3464
R6254 a_n2686_12778.n14 a_n2686_12778.n123 48.4088
R6255 a_n2686_12778.n15 a_n2686_12778.n121 48.4088
R6256 a_n2686_12778.n13 a_n2686_12778.n64 48.4088
R6257 a_n2686_12778.n242 a_n2686_12778.n236 23.9181
R6258 a_n2686_12778.n137 a_n2686_12778.n136 16.477
R6259 a_n2686_12778.n134 a_n2686_12778.n49 40.5394
R6260 a_n2686_12778.n227 a_n2686_12778.n226 16.477
R6261 a_n2686_12778.n229 a_n2686_12778.n228 16.477
R6262 a_n2686_12778.n219 a_n2686_12778.n218 16.477
R6263 a_n2686_12778.n221 a_n2686_12778.n220 16.477
R6264 a_n2686_12778.n211 a_n2686_12778.n210 16.477
R6265 a_n2686_12778.n213 a_n2686_12778.n212 16.477
R6266 a_n2686_12778.n203 a_n2686_12778.n202 16.477
R6267 a_n2686_12778.n205 a_n2686_12778.n204 16.477
R6268 a_n2686_12778.n14 a_n2686_12778.n127 40.5394
R6269 a_n2686_12778.n125 a_n2686_12778.n19 40.5394
R6270 a_n2686_12778.n15 a_n2686_12778.n130 40.5394
R6271 a_n2686_12778.n128 a_n2686_12778.n17 40.5394
R6272 a_n2686_12778.n13 a_n2686_12778.n235 40.5394
R6273 a_n2686_12778.n233 a_n2686_12778.n21 40.5394
R6274 a_n2686_12778.n104 a_n2686_12778.n102 16.3865
R6275 a_n2686_12778.n75 a_n2686_12778.n73 16.3865
R6276 a_n2686_12778.n152 a_n2686_12778.n150 16.3865
R6277 a_n2686_12778.n181 a_n2686_12778.n179 16.3865
R6278 a_n2686_12778.n105 a_n2686_12778.n101 12.8005
R6279 a_n2686_12778.n76 a_n2686_12778.n72 12.8005
R6280 a_n2686_12778.n153 a_n2686_12778.n149 12.8005
R6281 a_n2686_12778.n182 a_n2686_12778.n178 12.8005
R6282 a_n2686_12778.n107 a_n2686_12778.n106 12.0247
R6283 a_n2686_12778.n78 a_n2686_12778.n77 12.0247
R6284 a_n2686_12778.n155 a_n2686_12778.n154 12.0247
R6285 a_n2686_12778.n184 a_n2686_12778.n183 12.0247
R6286 a_n2686_12778.n110 a_n2686_12778.n99 11.249
R6287 a_n2686_12778.n81 a_n2686_12778.n70 11.249
R6288 a_n2686_12778.n158 a_n2686_12778.n147 11.249
R6289 a_n2686_12778.n187 a_n2686_12778.n176 11.249
R6290 a_n2686_12778.n199 a_n2686_12778.n7 10.8153
R6291 a_n2686_12778.n0 a_n2686_12778.n232 10.6108
R6292 a_n2686_12778.n111 a_n2686_12778.n98 10.4732
R6293 a_n2686_12778.n82 a_n2686_12778.n69 10.4732
R6294 a_n2686_12778.n159 a_n2686_12778.n146 10.4732
R6295 a_n2686_12778.n188 a_n2686_12778.n175 10.4732
R6296 a_n2686_12778.n113 a_n2686_12778.n112 9.69747
R6297 a_n2686_12778.n84 a_n2686_12778.n83 9.69747
R6298 a_n2686_12778.n161 a_n2686_12778.n160 9.69747
R6299 a_n2686_12778.n190 a_n2686_12778.n189 9.69747
R6300 a_n2686_12778.n119 a_n2686_12778.n118 9.45567
R6301 a_n2686_12778.n90 a_n2686_12778.n89 9.45567
R6302 a_n2686_12778.n167 a_n2686_12778.n166 9.45567
R6303 a_n2686_12778.n196 a_n2686_12778.n195 9.45567
R6304 a_n2686_12778.n198 a_n2686_12778.n142 9.30587
R6305 a_n2686_12778.n118 a_n2686_12778.n117 9.3005
R6306 a_n2686_12778.n96 a_n2686_12778.n53 9.3005
R6307 a_n2686_12778.n112 a_n2686_12778.n53 9.3005
R6308 a_n2686_12778.n52 a_n2686_12778.n111 9.3005
R6309 a_n2686_12778.n99 a_n2686_12778.n52 9.3005
R6310 a_n2686_12778.n106 a_n2686_12778.n54 9.3005
R6311 a_n2686_12778.n54 a_n2686_12778.n105 9.3005
R6312 a_n2686_12778.n89 a_n2686_12778.n88 9.3005
R6313 a_n2686_12778.n67 a_n2686_12778.n56 9.3005
R6314 a_n2686_12778.n83 a_n2686_12778.n56 9.3005
R6315 a_n2686_12778.n55 a_n2686_12778.n82 9.3005
R6316 a_n2686_12778.n70 a_n2686_12778.n55 9.3005
R6317 a_n2686_12778.n77 a_n2686_12778.n57 9.3005
R6318 a_n2686_12778.n57 a_n2686_12778.n76 9.3005
R6319 a_n2686_12778.n166 a_n2686_12778.n165 9.3005
R6320 a_n2686_12778.n144 a_n2686_12778.n59 9.3005
R6321 a_n2686_12778.n160 a_n2686_12778.n59 9.3005
R6322 a_n2686_12778.n58 a_n2686_12778.n159 9.3005
R6323 a_n2686_12778.n147 a_n2686_12778.n58 9.3005
R6324 a_n2686_12778.n154 a_n2686_12778.n60 9.3005
R6325 a_n2686_12778.n60 a_n2686_12778.n153 9.3005
R6326 a_n2686_12778.n195 a_n2686_12778.n194 9.3005
R6327 a_n2686_12778.n173 a_n2686_12778.n62 9.3005
R6328 a_n2686_12778.n189 a_n2686_12778.n62 9.3005
R6329 a_n2686_12778.n61 a_n2686_12778.n188 9.3005
R6330 a_n2686_12778.n176 a_n2686_12778.n61 9.3005
R6331 a_n2686_12778.n183 a_n2686_12778.n63 9.3005
R6332 a_n2686_12778.n63 a_n2686_12778.n182 9.3005
R6333 a_n2686_12778.n116 a_n2686_12778.n96 8.92171
R6334 a_n2686_12778.n87 a_n2686_12778.n67 8.92171
R6335 a_n2686_12778.n164 a_n2686_12778.n144 8.92171
R6336 a_n2686_12778.n193 a_n2686_12778.n173 8.92171
R6337 a_n2686_12778.n2 a_n2686_12778.n120 8.2571
R6338 a_n2686_12778.n117 a_n2686_12778.n95 8.14595
R6339 a_n2686_12778.n88 a_n2686_12778.n66 8.14595
R6340 a_n2686_12778.n165 a_n2686_12778.n143 8.14595
R6341 a_n2686_12778.n194 a_n2686_12778.n172 8.14595
R6342 a_n2686_12778.n136 a_n2686_12778.n135 8.11581
R6343 a_n2686_12778.n38 a_n2686_12778.n227 26.1378
R6344 a_n2686_12778.n228 a_n2686_12778.n37 8.11581
R6345 a_n2686_12778.n33 a_n2686_12778.n219 26.1378
R6346 a_n2686_12778.n220 a_n2686_12778.n32 8.11581
R6347 a_n2686_12778.n28 a_n2686_12778.n211 26.1378
R6348 a_n2686_12778.n212 a_n2686_12778.n27 8.11581
R6349 a_n2686_12778.n23 a_n2686_12778.n203 26.1378
R6350 a_n2686_12778.n204 a_n2686_12778.n22 8.11581
R6351 a_n2686_12778.n127 a_n2686_12778.n126 8.11581
R6352 a_n2686_12778.n130 a_n2686_12778.n129 8.11581
R6353 a_n2686_12778.n235 a_n2686_12778.n234 8.11581
R6354 a_n2686_12778.n232 a_n2686_12778.n231 7.00284
R6355 a_n2686_12778.n200 a_n2686_12778.n199 7.00284
R6356 a_n2686_12778.n3 a_n2686_12778.n2 6.60701
R6357 a_n2686_12778.n119 a_n2686_12778.n95 5.81868
R6358 a_n2686_12778.n90 a_n2686_12778.n66 5.81868
R6359 a_n2686_12778.n167 a_n2686_12778.n143 5.81868
R6360 a_n2686_12778.n196 a_n2686_12778.n172 5.81868
R6361 a_n2686_12778.n198 a_n2686_12778.n197 5.55007
R6362 a_n2686_12778.n93 a_n2686_12778.t26 5.418
R6363 a_n2686_12778.n93 a_n2686_12778.t14 5.418
R6364 a_n2686_12778.n91 a_n2686_12778.t20 5.418
R6365 a_n2686_12778.n91 a_n2686_12778.t18 5.418
R6366 a_n2686_12778.n168 a_n2686_12778.t30 5.418
R6367 a_n2686_12778.n168 a_n2686_12778.t10 5.418
R6368 a_n2686_12778.n170 a_n2686_12778.t28 5.418
R6369 a_n2686_12778.n170 a_n2686_12778.t8 5.418
R6370 a_n2686_12778.n117 a_n2686_12778.n116 5.04292
R6371 a_n2686_12778.n88 a_n2686_12778.n87 5.04292
R6372 a_n2686_12778.n165 a_n2686_12778.n164 5.04292
R6373 a_n2686_12778.n194 a_n2686_12778.n193 5.04292
R6374 a_n2686_12778.n5 a_n2686_12778.n9 4.52033
R6375 a_n2686_12778.n113 a_n2686_12778.n96 4.26717
R6376 a_n2686_12778.n84 a_n2686_12778.n67 4.26717
R6377 a_n2686_12778.n161 a_n2686_12778.n144 4.26717
R6378 a_n2686_12778.n190 a_n2686_12778.n173 4.26717
R6379 a_n2686_12778.n232 a_n2686_12778.n2 4.20883
R6380 a_n2686_12778.n54 a_n2686_12778.n102 3.71286
R6381 a_n2686_12778.n57 a_n2686_12778.n73 3.71286
R6382 a_n2686_12778.n60 a_n2686_12778.n150 3.71286
R6383 a_n2686_12778.n63 a_n2686_12778.n179 3.71286
R6384 a_n2686_12778.n112 a_n2686_12778.n98 3.49141
R6385 a_n2686_12778.n83 a_n2686_12778.n69 3.49141
R6386 a_n2686_12778.n160 a_n2686_12778.n146 3.49141
R6387 a_n2686_12778.n189 a_n2686_12778.n175 3.49141
R6388 a_n2686_12778.n236 a_n2686_12778.n11 3.45549
R6389 a_n2686_12778.n240 a_n2686_12778.t2 2.82907
R6390 a_n2686_12778.n240 a_n2686_12778.t3 2.82907
R6391 a_n2686_12778.n238 a_n2686_12778.t4 2.82907
R6392 a_n2686_12778.n238 a_n2686_12778.t6 2.82907
R6393 a_n2686_12778.n237 a_n2686_12778.t31 2.82907
R6394 a_n2686_12778.n237 a_n2686_12778.t1 2.82907
R6395 a_n2686_12778.t0 a_n2686_12778.n243 2.82907
R6396 a_n2686_12778.n243 a_n2686_12778.t5 2.82907
R6397 a_n2686_12778.n111 a_n2686_12778.n110 2.71565
R6398 a_n2686_12778.n82 a_n2686_12778.n81 2.71565
R6399 a_n2686_12778.n159 a_n2686_12778.n158 2.71565
R6400 a_n2686_12778.n188 a_n2686_12778.n187 2.71565
R6401 a_n2686_12778.n107 a_n2686_12778.n99 1.93989
R6402 a_n2686_12778.n78 a_n2686_12778.n70 1.93989
R6403 a_n2686_12778.n155 a_n2686_12778.n147 1.93989
R6404 a_n2686_12778.n184 a_n2686_12778.n176 1.93989
R6405 a_n2686_12778.n216 a_n2686_12778.n215 1.42563
R6406 a_n2686_12778.n199 a_n2686_12778.n198 1.30542
R6407 a_n2686_12778.n106 a_n2686_12778.n101 1.16414
R6408 a_n2686_12778.n77 a_n2686_12778.n72 1.16414
R6409 a_n2686_12778.n154 a_n2686_12778.n149 1.16414
R6410 a_n2686_12778.n183 a_n2686_12778.n178 1.16414
R6411 a_n2686_12778.n236 a_n2686_12778.n50 1.02746
R6412 a_n2686_12778.n208 a_n2686_12778.n207 0.96351
R6413 a_n2686_12778.n224 a_n2686_12778.n223 0.96351
R6414 a_n2686_12778.n94 a_n2686_12778.n92 0.573776
R6415 a_n2686_12778.n120 a_n2686_12778.n94 0.573776
R6416 a_n2686_12778.n197 a_n2686_12778.n171 0.573776
R6417 a_n2686_12778.n171 a_n2686_12778.n169 0.573776
R6418 a_n2686_12778.n105 a_n2686_12778.n104 0.388379
R6419 a_n2686_12778.n76 a_n2686_12778.n75 0.388379
R6420 a_n2686_12778.n153 a_n2686_12778.n152 0.388379
R6421 a_n2686_12778.n182 a_n2686_12778.n181 0.388379
R6422 a_n2686_12778.n46 a_n2686_12778.n48 0.379288
R6423 a_n2686_12778.n63 a_n2686_12778.n61 0.310845
R6424 a_n2686_12778.n62 a_n2686_12778.n61 0.310845
R6425 a_n2686_12778.n195 a_n2686_12778.n62 0.310845
R6426 a_n2686_12778.n60 a_n2686_12778.n58 0.310845
R6427 a_n2686_12778.n59 a_n2686_12778.n58 0.310845
R6428 a_n2686_12778.n166 a_n2686_12778.n59 0.310845
R6429 a_n2686_12778.n57 a_n2686_12778.n55 0.310845
R6430 a_n2686_12778.n56 a_n2686_12778.n55 0.310845
R6431 a_n2686_12778.n89 a_n2686_12778.n56 0.310845
R6432 a_n2686_12778.n54 a_n2686_12778.n52 0.310845
R6433 a_n2686_12778.n53 a_n2686_12778.n52 0.310845
R6434 a_n2686_12778.n118 a_n2686_12778.n53 0.310845
R6435 a_n2686_12778.n242 a_n2686_12778.n241 0.287138
R6436 a_n2686_12778.n200 a_n2686_12778.n24 0.285035
R6437 a_n2686_12778.n207 a_n2686_12778.n26 0.285035
R6438 a_n2686_12778.n208 a_n2686_12778.n29 0.285035
R6439 a_n2686_12778.n215 a_n2686_12778.n31 0.285035
R6440 a_n2686_12778.n216 a_n2686_12778.n34 0.285035
R6441 a_n2686_12778.n223 a_n2686_12778.n36 0.285035
R6442 a_n2686_12778.n224 a_n2686_12778.n39 0.285035
R6443 a_n2686_12778.n231 a_n2686_12778.n41 0.285035
R6444 a_n2686_12778.n142 a_n2686_12778.n43 0.285035
R6445 a_n2686_12778.n48 a_n2686_12778.n50 0.285035
R6446 a_n2686_12778.n139 a_n2686_12778.n131 0.246418
R6447 a_n2686_12778.n51 a_n2686_12778.n132 11.8807
R6448 a_n2686_12778.n45 a_n2686_12778.n46 0.379288
R6449 a_n2686_12778.n42 a_n2686_12778.n45 0.379288
R6450 a_n2686_12778.n44 a_n2686_12778.n42 0.379288
R6451 a_n2686_12778.n44 a_n2686_12778.n43 0.379288
R6452 a_n2686_12778.n41 a_n2686_12778.n40 0.379288
R6453 a_n2686_12778.n40 a_n2686_12778.n39 0.379288
R6454 a_n2686_12778.n36 a_n2686_12778.n35 0.379288
R6455 a_n2686_12778.n35 a_n2686_12778.n34 0.379288
R6456 a_n2686_12778.n31 a_n2686_12778.n30 0.379288
R6457 a_n2686_12778.n30 a_n2686_12778.n29 0.379288
R6458 a_n2686_12778.n26 a_n2686_12778.n25 0.379288
R6459 a_n2686_12778.n25 a_n2686_12778.n24 0.379288
R6460 a_n2686_12778.n4 a_n2686_12778.n124 32.4972
R6461 a_n2686_12778.n6 a_n2686_12778.n122 32.4972
R6462 a_n2686_12778.n1 a_n2686_12778.n65 32.4972
R6463 a_n2686_12778.n7 a_n2686_12778.n5 2.46351
R6464 a_n2686_12778.n9 a_n2686_12778.n3 2.46351
R6465 a_n2686_12778.n11 a_n2686_12778.n0 2.46351
R6466 a_n2686_8422.n258 a_n2686_8422.n232 756.745
R6467 a_n2686_8422.n226 a_n2686_8422.n200 756.745
R6468 a_n2686_8422.n93 a_n2686_8422.n67 756.745
R6469 a_n2686_8422.n126 a_n2686_8422.n100 756.745
R6470 a_n2686_8422.n158 a_n2686_8422.n132 756.745
R6471 a_n2686_8422.n192 a_n2686_8422.n166 756.745
R6472 a_n2686_8422.n26 a_n2686_8422.n0 756.745
R6473 a_n2686_8422.n61 a_n2686_8422.n35 756.745
R6474 a_n2686_8422.n259 a_n2686_8422.n258 585
R6475 a_n2686_8422.n257 a_n2686_8422.n256 585
R6476 a_n2686_8422.n236 a_n2686_8422.n235 585
R6477 a_n2686_8422.n251 a_n2686_8422.n250 585
R6478 a_n2686_8422.n249 a_n2686_8422.n248 585
R6479 a_n2686_8422.n240 a_n2686_8422.n239 585
R6480 a_n2686_8422.n243 a_n2686_8422.n242 585
R6481 a_n2686_8422.n227 a_n2686_8422.n226 585
R6482 a_n2686_8422.n225 a_n2686_8422.n224 585
R6483 a_n2686_8422.n204 a_n2686_8422.n203 585
R6484 a_n2686_8422.n219 a_n2686_8422.n218 585
R6485 a_n2686_8422.n217 a_n2686_8422.n216 585
R6486 a_n2686_8422.n208 a_n2686_8422.n207 585
R6487 a_n2686_8422.n211 a_n2686_8422.n210 585
R6488 a_n2686_8422.n94 a_n2686_8422.n93 585
R6489 a_n2686_8422.n92 a_n2686_8422.n91 585
R6490 a_n2686_8422.n71 a_n2686_8422.n70 585
R6491 a_n2686_8422.n86 a_n2686_8422.n85 585
R6492 a_n2686_8422.n84 a_n2686_8422.n83 585
R6493 a_n2686_8422.n75 a_n2686_8422.n74 585
R6494 a_n2686_8422.n78 a_n2686_8422.n77 585
R6495 a_n2686_8422.n127 a_n2686_8422.n126 585
R6496 a_n2686_8422.n125 a_n2686_8422.n124 585
R6497 a_n2686_8422.n104 a_n2686_8422.n103 585
R6498 a_n2686_8422.n119 a_n2686_8422.n118 585
R6499 a_n2686_8422.n117 a_n2686_8422.n116 585
R6500 a_n2686_8422.n108 a_n2686_8422.n107 585
R6501 a_n2686_8422.n111 a_n2686_8422.n110 585
R6502 a_n2686_8422.n159 a_n2686_8422.n158 585
R6503 a_n2686_8422.n157 a_n2686_8422.n156 585
R6504 a_n2686_8422.n136 a_n2686_8422.n135 585
R6505 a_n2686_8422.n151 a_n2686_8422.n150 585
R6506 a_n2686_8422.n149 a_n2686_8422.n148 585
R6507 a_n2686_8422.n140 a_n2686_8422.n139 585
R6508 a_n2686_8422.n143 a_n2686_8422.n142 585
R6509 a_n2686_8422.n193 a_n2686_8422.n192 585
R6510 a_n2686_8422.n191 a_n2686_8422.n190 585
R6511 a_n2686_8422.n170 a_n2686_8422.n169 585
R6512 a_n2686_8422.n185 a_n2686_8422.n184 585
R6513 a_n2686_8422.n183 a_n2686_8422.n182 585
R6514 a_n2686_8422.n174 a_n2686_8422.n173 585
R6515 a_n2686_8422.n177 a_n2686_8422.n176 585
R6516 a_n2686_8422.n27 a_n2686_8422.n26 585
R6517 a_n2686_8422.n25 a_n2686_8422.n24 585
R6518 a_n2686_8422.n4 a_n2686_8422.n3 585
R6519 a_n2686_8422.n19 a_n2686_8422.n18 585
R6520 a_n2686_8422.n17 a_n2686_8422.n16 585
R6521 a_n2686_8422.n8 a_n2686_8422.n7 585
R6522 a_n2686_8422.n11 a_n2686_8422.n10 585
R6523 a_n2686_8422.n62 a_n2686_8422.n61 585
R6524 a_n2686_8422.n60 a_n2686_8422.n59 585
R6525 a_n2686_8422.n39 a_n2686_8422.n38 585
R6526 a_n2686_8422.n54 a_n2686_8422.n53 585
R6527 a_n2686_8422.n52 a_n2686_8422.n51 585
R6528 a_n2686_8422.n43 a_n2686_8422.n42 585
R6529 a_n2686_8422.n46 a_n2686_8422.n45 585
R6530 a_n2686_8422.t17 a_n2686_8422.n241 327.601
R6531 a_n2686_8422.t10 a_n2686_8422.n209 327.601
R6532 a_n2686_8422.t6 a_n2686_8422.n76 327.601
R6533 a_n2686_8422.t1 a_n2686_8422.n109 327.601
R6534 a_n2686_8422.t5 a_n2686_8422.n141 327.601
R6535 a_n2686_8422.t7 a_n2686_8422.n175 327.601
R6536 a_n2686_8422.t15 a_n2686_8422.n9 327.601
R6537 a_n2686_8422.t16 a_n2686_8422.n44 327.601
R6538 a_n2686_8422.n258 a_n2686_8422.n257 171.744
R6539 a_n2686_8422.n257 a_n2686_8422.n235 171.744
R6540 a_n2686_8422.n250 a_n2686_8422.n235 171.744
R6541 a_n2686_8422.n250 a_n2686_8422.n249 171.744
R6542 a_n2686_8422.n249 a_n2686_8422.n239 171.744
R6543 a_n2686_8422.n242 a_n2686_8422.n239 171.744
R6544 a_n2686_8422.n226 a_n2686_8422.n225 171.744
R6545 a_n2686_8422.n225 a_n2686_8422.n203 171.744
R6546 a_n2686_8422.n218 a_n2686_8422.n203 171.744
R6547 a_n2686_8422.n218 a_n2686_8422.n217 171.744
R6548 a_n2686_8422.n217 a_n2686_8422.n207 171.744
R6549 a_n2686_8422.n210 a_n2686_8422.n207 171.744
R6550 a_n2686_8422.n93 a_n2686_8422.n92 171.744
R6551 a_n2686_8422.n92 a_n2686_8422.n70 171.744
R6552 a_n2686_8422.n85 a_n2686_8422.n70 171.744
R6553 a_n2686_8422.n85 a_n2686_8422.n84 171.744
R6554 a_n2686_8422.n84 a_n2686_8422.n74 171.744
R6555 a_n2686_8422.n77 a_n2686_8422.n74 171.744
R6556 a_n2686_8422.n126 a_n2686_8422.n125 171.744
R6557 a_n2686_8422.n125 a_n2686_8422.n103 171.744
R6558 a_n2686_8422.n118 a_n2686_8422.n103 171.744
R6559 a_n2686_8422.n118 a_n2686_8422.n117 171.744
R6560 a_n2686_8422.n117 a_n2686_8422.n107 171.744
R6561 a_n2686_8422.n110 a_n2686_8422.n107 171.744
R6562 a_n2686_8422.n158 a_n2686_8422.n157 171.744
R6563 a_n2686_8422.n157 a_n2686_8422.n135 171.744
R6564 a_n2686_8422.n150 a_n2686_8422.n135 171.744
R6565 a_n2686_8422.n150 a_n2686_8422.n149 171.744
R6566 a_n2686_8422.n149 a_n2686_8422.n139 171.744
R6567 a_n2686_8422.n142 a_n2686_8422.n139 171.744
R6568 a_n2686_8422.n192 a_n2686_8422.n191 171.744
R6569 a_n2686_8422.n191 a_n2686_8422.n169 171.744
R6570 a_n2686_8422.n184 a_n2686_8422.n169 171.744
R6571 a_n2686_8422.n184 a_n2686_8422.n183 171.744
R6572 a_n2686_8422.n183 a_n2686_8422.n173 171.744
R6573 a_n2686_8422.n176 a_n2686_8422.n173 171.744
R6574 a_n2686_8422.n26 a_n2686_8422.n25 171.744
R6575 a_n2686_8422.n25 a_n2686_8422.n3 171.744
R6576 a_n2686_8422.n18 a_n2686_8422.n3 171.744
R6577 a_n2686_8422.n18 a_n2686_8422.n17 171.744
R6578 a_n2686_8422.n17 a_n2686_8422.n7 171.744
R6579 a_n2686_8422.n10 a_n2686_8422.n7 171.744
R6580 a_n2686_8422.n61 a_n2686_8422.n60 171.744
R6581 a_n2686_8422.n60 a_n2686_8422.n38 171.744
R6582 a_n2686_8422.n53 a_n2686_8422.n38 171.744
R6583 a_n2686_8422.n53 a_n2686_8422.n52 171.744
R6584 a_n2686_8422.n52 a_n2686_8422.n42 171.744
R6585 a_n2686_8422.n45 a_n2686_8422.n42 171.744
R6586 a_n2686_8422.n242 a_n2686_8422.t17 85.8723
R6587 a_n2686_8422.n210 a_n2686_8422.t10 85.8723
R6588 a_n2686_8422.n77 a_n2686_8422.t6 85.8723
R6589 a_n2686_8422.n110 a_n2686_8422.t1 85.8723
R6590 a_n2686_8422.n142 a_n2686_8422.t5 85.8723
R6591 a_n2686_8422.n176 a_n2686_8422.t7 85.8723
R6592 a_n2686_8422.n10 a_n2686_8422.t15 85.8723
R6593 a_n2686_8422.n45 a_n2686_8422.t16 85.8723
R6594 a_n2686_8422.n264 a_n2686_8422.n263 81.2397
R6595 a_n2686_8422.n99 a_n2686_8422.n98 81.2397
R6596 a_n2686_8422.n165 a_n2686_8422.n164 81.2397
R6597 a_n2686_8422.n32 a_n2686_8422.n31 81.2397
R6598 a_n2686_8422.n34 a_n2686_8422.n33 81.2397
R6599 a_n2686_8422.n266 a_n2686_8422.n265 81.2397
R6600 a_n2686_8422.n264 a_n2686_8422.n262 38.3829
R6601 a_n2686_8422.n99 a_n2686_8422.n97 38.3829
R6602 a_n2686_8422.n32 a_n2686_8422.n30 38.3829
R6603 a_n2686_8422.n231 a_n2686_8422.n230 37.8096
R6604 a_n2686_8422.n131 a_n2686_8422.n130 37.8096
R6605 a_n2686_8422.n163 a_n2686_8422.n162 37.8096
R6606 a_n2686_8422.n197 a_n2686_8422.n196 37.8096
R6607 a_n2686_8422.n66 a_n2686_8422.n65 37.8096
R6608 a_n2686_8422.n198 a_n2686_8422.n66 22.3736
R6609 a_n2686_8422.n243 a_n2686_8422.n241 16.3865
R6610 a_n2686_8422.n211 a_n2686_8422.n209 16.3865
R6611 a_n2686_8422.n78 a_n2686_8422.n76 16.3865
R6612 a_n2686_8422.n111 a_n2686_8422.n109 16.3865
R6613 a_n2686_8422.n143 a_n2686_8422.n141 16.3865
R6614 a_n2686_8422.n177 a_n2686_8422.n175 16.3865
R6615 a_n2686_8422.n11 a_n2686_8422.n9 16.3865
R6616 a_n2686_8422.n46 a_n2686_8422.n44 16.3865
R6617 a_n2686_8422.n244 a_n2686_8422.n240 12.8005
R6618 a_n2686_8422.n212 a_n2686_8422.n208 12.8005
R6619 a_n2686_8422.n79 a_n2686_8422.n75 12.8005
R6620 a_n2686_8422.n112 a_n2686_8422.n108 12.8005
R6621 a_n2686_8422.n144 a_n2686_8422.n140 12.8005
R6622 a_n2686_8422.n178 a_n2686_8422.n174 12.8005
R6623 a_n2686_8422.n12 a_n2686_8422.n8 12.8005
R6624 a_n2686_8422.n47 a_n2686_8422.n43 12.8005
R6625 a_n2686_8422.n248 a_n2686_8422.n247 12.0247
R6626 a_n2686_8422.n216 a_n2686_8422.n215 12.0247
R6627 a_n2686_8422.n83 a_n2686_8422.n82 12.0247
R6628 a_n2686_8422.n116 a_n2686_8422.n115 12.0247
R6629 a_n2686_8422.n148 a_n2686_8422.n147 12.0247
R6630 a_n2686_8422.n182 a_n2686_8422.n181 12.0247
R6631 a_n2686_8422.n16 a_n2686_8422.n15 12.0247
R6632 a_n2686_8422.n51 a_n2686_8422.n50 12.0247
R6633 a_n2686_8422.n251 a_n2686_8422.n238 11.249
R6634 a_n2686_8422.n219 a_n2686_8422.n206 11.249
R6635 a_n2686_8422.n86 a_n2686_8422.n73 11.249
R6636 a_n2686_8422.n119 a_n2686_8422.n106 11.249
R6637 a_n2686_8422.n151 a_n2686_8422.n138 11.249
R6638 a_n2686_8422.n185 a_n2686_8422.n172 11.249
R6639 a_n2686_8422.n19 a_n2686_8422.n6 11.249
R6640 a_n2686_8422.n54 a_n2686_8422.n41 11.249
R6641 a_n2686_8422.n252 a_n2686_8422.n236 10.4732
R6642 a_n2686_8422.n220 a_n2686_8422.n204 10.4732
R6643 a_n2686_8422.n87 a_n2686_8422.n71 10.4732
R6644 a_n2686_8422.n120 a_n2686_8422.n104 10.4732
R6645 a_n2686_8422.n152 a_n2686_8422.n136 10.4732
R6646 a_n2686_8422.n186 a_n2686_8422.n170 10.4732
R6647 a_n2686_8422.n20 a_n2686_8422.n4 10.4732
R6648 a_n2686_8422.n55 a_n2686_8422.n39 10.4732
R6649 a_n2686_8422.n256 a_n2686_8422.n255 9.69747
R6650 a_n2686_8422.n224 a_n2686_8422.n223 9.69747
R6651 a_n2686_8422.n91 a_n2686_8422.n90 9.69747
R6652 a_n2686_8422.n124 a_n2686_8422.n123 9.69747
R6653 a_n2686_8422.n156 a_n2686_8422.n155 9.69747
R6654 a_n2686_8422.n190 a_n2686_8422.n189 9.69747
R6655 a_n2686_8422.n24 a_n2686_8422.n23 9.69747
R6656 a_n2686_8422.n59 a_n2686_8422.n58 9.69747
R6657 a_n2686_8422.n262 a_n2686_8422.n261 9.45567
R6658 a_n2686_8422.n230 a_n2686_8422.n229 9.45567
R6659 a_n2686_8422.n97 a_n2686_8422.n96 9.45567
R6660 a_n2686_8422.n130 a_n2686_8422.n129 9.45567
R6661 a_n2686_8422.n162 a_n2686_8422.n161 9.45567
R6662 a_n2686_8422.n196 a_n2686_8422.n195 9.45567
R6663 a_n2686_8422.n30 a_n2686_8422.n29 9.45567
R6664 a_n2686_8422.n65 a_n2686_8422.n64 9.45567
R6665 a_n2686_8422.n261 a_n2686_8422.n260 9.3005
R6666 a_n2686_8422.n234 a_n2686_8422.n233 9.3005
R6667 a_n2686_8422.n255 a_n2686_8422.n254 9.3005
R6668 a_n2686_8422.n253 a_n2686_8422.n252 9.3005
R6669 a_n2686_8422.n238 a_n2686_8422.n237 9.3005
R6670 a_n2686_8422.n247 a_n2686_8422.n246 9.3005
R6671 a_n2686_8422.n245 a_n2686_8422.n244 9.3005
R6672 a_n2686_8422.n229 a_n2686_8422.n228 9.3005
R6673 a_n2686_8422.n202 a_n2686_8422.n201 9.3005
R6674 a_n2686_8422.n223 a_n2686_8422.n222 9.3005
R6675 a_n2686_8422.n221 a_n2686_8422.n220 9.3005
R6676 a_n2686_8422.n206 a_n2686_8422.n205 9.3005
R6677 a_n2686_8422.n215 a_n2686_8422.n214 9.3005
R6678 a_n2686_8422.n213 a_n2686_8422.n212 9.3005
R6679 a_n2686_8422.n96 a_n2686_8422.n95 9.3005
R6680 a_n2686_8422.n69 a_n2686_8422.n68 9.3005
R6681 a_n2686_8422.n90 a_n2686_8422.n89 9.3005
R6682 a_n2686_8422.n88 a_n2686_8422.n87 9.3005
R6683 a_n2686_8422.n73 a_n2686_8422.n72 9.3005
R6684 a_n2686_8422.n82 a_n2686_8422.n81 9.3005
R6685 a_n2686_8422.n80 a_n2686_8422.n79 9.3005
R6686 a_n2686_8422.n129 a_n2686_8422.n128 9.3005
R6687 a_n2686_8422.n102 a_n2686_8422.n101 9.3005
R6688 a_n2686_8422.n123 a_n2686_8422.n122 9.3005
R6689 a_n2686_8422.n121 a_n2686_8422.n120 9.3005
R6690 a_n2686_8422.n106 a_n2686_8422.n105 9.3005
R6691 a_n2686_8422.n115 a_n2686_8422.n114 9.3005
R6692 a_n2686_8422.n113 a_n2686_8422.n112 9.3005
R6693 a_n2686_8422.n161 a_n2686_8422.n160 9.3005
R6694 a_n2686_8422.n134 a_n2686_8422.n133 9.3005
R6695 a_n2686_8422.n155 a_n2686_8422.n154 9.3005
R6696 a_n2686_8422.n153 a_n2686_8422.n152 9.3005
R6697 a_n2686_8422.n138 a_n2686_8422.n137 9.3005
R6698 a_n2686_8422.n147 a_n2686_8422.n146 9.3005
R6699 a_n2686_8422.n145 a_n2686_8422.n144 9.3005
R6700 a_n2686_8422.n195 a_n2686_8422.n194 9.3005
R6701 a_n2686_8422.n168 a_n2686_8422.n167 9.3005
R6702 a_n2686_8422.n189 a_n2686_8422.n188 9.3005
R6703 a_n2686_8422.n187 a_n2686_8422.n186 9.3005
R6704 a_n2686_8422.n172 a_n2686_8422.n171 9.3005
R6705 a_n2686_8422.n181 a_n2686_8422.n180 9.3005
R6706 a_n2686_8422.n179 a_n2686_8422.n178 9.3005
R6707 a_n2686_8422.n29 a_n2686_8422.n28 9.3005
R6708 a_n2686_8422.n2 a_n2686_8422.n1 9.3005
R6709 a_n2686_8422.n23 a_n2686_8422.n22 9.3005
R6710 a_n2686_8422.n21 a_n2686_8422.n20 9.3005
R6711 a_n2686_8422.n6 a_n2686_8422.n5 9.3005
R6712 a_n2686_8422.n15 a_n2686_8422.n14 9.3005
R6713 a_n2686_8422.n13 a_n2686_8422.n12 9.3005
R6714 a_n2686_8422.n64 a_n2686_8422.n63 9.3005
R6715 a_n2686_8422.n37 a_n2686_8422.n36 9.3005
R6716 a_n2686_8422.n58 a_n2686_8422.n57 9.3005
R6717 a_n2686_8422.n56 a_n2686_8422.n55 9.3005
R6718 a_n2686_8422.n41 a_n2686_8422.n40 9.3005
R6719 a_n2686_8422.n50 a_n2686_8422.n49 9.3005
R6720 a_n2686_8422.n48 a_n2686_8422.n47 9.3005
R6721 a_n2686_8422.n259 a_n2686_8422.n234 8.92171
R6722 a_n2686_8422.n227 a_n2686_8422.n202 8.92171
R6723 a_n2686_8422.n94 a_n2686_8422.n69 8.92171
R6724 a_n2686_8422.n127 a_n2686_8422.n102 8.92171
R6725 a_n2686_8422.n159 a_n2686_8422.n134 8.92171
R6726 a_n2686_8422.n193 a_n2686_8422.n168 8.92171
R6727 a_n2686_8422.n27 a_n2686_8422.n2 8.92171
R6728 a_n2686_8422.n62 a_n2686_8422.n37 8.92171
R6729 a_n2686_8422.n199 a_n2686_8422.t20 8.43517
R6730 a_n2686_8422.n260 a_n2686_8422.n232 8.14595
R6731 a_n2686_8422.n228 a_n2686_8422.n200 8.14595
R6732 a_n2686_8422.n95 a_n2686_8422.n67 8.14595
R6733 a_n2686_8422.n128 a_n2686_8422.n100 8.14595
R6734 a_n2686_8422.n160 a_n2686_8422.n132 8.14595
R6735 a_n2686_8422.n194 a_n2686_8422.n166 8.14595
R6736 a_n2686_8422.n28 a_n2686_8422.n0 8.14595
R6737 a_n2686_8422.n63 a_n2686_8422.n35 8.14595
R6738 a_n2686_8422.n198 a_n2686_8422.n197 5.91753
R6739 a_n2686_8422.n262 a_n2686_8422.n232 5.81868
R6740 a_n2686_8422.n230 a_n2686_8422.n200 5.81868
R6741 a_n2686_8422.n97 a_n2686_8422.n67 5.81868
R6742 a_n2686_8422.n130 a_n2686_8422.n100 5.81868
R6743 a_n2686_8422.n162 a_n2686_8422.n132 5.81868
R6744 a_n2686_8422.n196 a_n2686_8422.n166 5.81868
R6745 a_n2686_8422.n30 a_n2686_8422.n0 5.81868
R6746 a_n2686_8422.n65 a_n2686_8422.n35 5.81868
R6747 a_n2686_8422.n231 a_n2686_8422.n199 5.72895
R6748 a_n2686_8422.n263 a_n2686_8422.t11 5.418
R6749 a_n2686_8422.n263 a_n2686_8422.t8 5.418
R6750 a_n2686_8422.n98 a_n2686_8422.t4 5.418
R6751 a_n2686_8422.n98 a_n2686_8422.t2 5.418
R6752 a_n2686_8422.n164 a_n2686_8422.t3 5.418
R6753 a_n2686_8422.n164 a_n2686_8422.t0 5.418
R6754 a_n2686_8422.n31 a_n2686_8422.t18 5.418
R6755 a_n2686_8422.n31 a_n2686_8422.t14 5.418
R6756 a_n2686_8422.n33 a_n2686_8422.t12 5.418
R6757 a_n2686_8422.n33 a_n2686_8422.t13 5.418
R6758 a_n2686_8422.n266 a_n2686_8422.t9 5.418
R6759 a_n2686_8422.t19 a_n2686_8422.n266 5.418
R6760 a_n2686_8422.n260 a_n2686_8422.n259 5.04292
R6761 a_n2686_8422.n228 a_n2686_8422.n227 5.04292
R6762 a_n2686_8422.n95 a_n2686_8422.n94 5.04292
R6763 a_n2686_8422.n128 a_n2686_8422.n127 5.04292
R6764 a_n2686_8422.n160 a_n2686_8422.n159 5.04292
R6765 a_n2686_8422.n194 a_n2686_8422.n193 5.04292
R6766 a_n2686_8422.n28 a_n2686_8422.n27 5.04292
R6767 a_n2686_8422.n63 a_n2686_8422.n62 5.04292
R6768 a_n2686_8422.n256 a_n2686_8422.n234 4.26717
R6769 a_n2686_8422.n224 a_n2686_8422.n202 4.26717
R6770 a_n2686_8422.n91 a_n2686_8422.n69 4.26717
R6771 a_n2686_8422.n124 a_n2686_8422.n102 4.26717
R6772 a_n2686_8422.n156 a_n2686_8422.n134 4.26717
R6773 a_n2686_8422.n190 a_n2686_8422.n168 4.26717
R6774 a_n2686_8422.n24 a_n2686_8422.n2 4.26717
R6775 a_n2686_8422.n59 a_n2686_8422.n37 4.26717
R6776 a_n2686_8422.n199 a_n2686_8422.n198 4.20883
R6777 a_n2686_8422.n245 a_n2686_8422.n241 3.71286
R6778 a_n2686_8422.n213 a_n2686_8422.n209 3.71286
R6779 a_n2686_8422.n80 a_n2686_8422.n76 3.71286
R6780 a_n2686_8422.n113 a_n2686_8422.n109 3.71286
R6781 a_n2686_8422.n145 a_n2686_8422.n141 3.71286
R6782 a_n2686_8422.n179 a_n2686_8422.n175 3.71286
R6783 a_n2686_8422.n13 a_n2686_8422.n9 3.71286
R6784 a_n2686_8422.n48 a_n2686_8422.n44 3.71286
R6785 a_n2686_8422.n255 a_n2686_8422.n236 3.49141
R6786 a_n2686_8422.n223 a_n2686_8422.n204 3.49141
R6787 a_n2686_8422.n90 a_n2686_8422.n71 3.49141
R6788 a_n2686_8422.n123 a_n2686_8422.n104 3.49141
R6789 a_n2686_8422.n155 a_n2686_8422.n136 3.49141
R6790 a_n2686_8422.n189 a_n2686_8422.n170 3.49141
R6791 a_n2686_8422.n23 a_n2686_8422.n4 3.49141
R6792 a_n2686_8422.n58 a_n2686_8422.n39 3.49141
R6793 a_n2686_8422.n252 a_n2686_8422.n251 2.71565
R6794 a_n2686_8422.n220 a_n2686_8422.n219 2.71565
R6795 a_n2686_8422.n87 a_n2686_8422.n86 2.71565
R6796 a_n2686_8422.n120 a_n2686_8422.n119 2.71565
R6797 a_n2686_8422.n152 a_n2686_8422.n151 2.71565
R6798 a_n2686_8422.n186 a_n2686_8422.n185 2.71565
R6799 a_n2686_8422.n20 a_n2686_8422.n19 2.71565
R6800 a_n2686_8422.n55 a_n2686_8422.n54 2.71565
R6801 a_n2686_8422.n248 a_n2686_8422.n238 1.93989
R6802 a_n2686_8422.n216 a_n2686_8422.n206 1.93989
R6803 a_n2686_8422.n83 a_n2686_8422.n73 1.93989
R6804 a_n2686_8422.n116 a_n2686_8422.n106 1.93989
R6805 a_n2686_8422.n148 a_n2686_8422.n138 1.93989
R6806 a_n2686_8422.n182 a_n2686_8422.n172 1.93989
R6807 a_n2686_8422.n16 a_n2686_8422.n6 1.93989
R6808 a_n2686_8422.n51 a_n2686_8422.n41 1.93989
R6809 a_n2686_8422.n247 a_n2686_8422.n240 1.16414
R6810 a_n2686_8422.n215 a_n2686_8422.n208 1.16414
R6811 a_n2686_8422.n82 a_n2686_8422.n75 1.16414
R6812 a_n2686_8422.n115 a_n2686_8422.n108 1.16414
R6813 a_n2686_8422.n147 a_n2686_8422.n140 1.16414
R6814 a_n2686_8422.n181 a_n2686_8422.n174 1.16414
R6815 a_n2686_8422.n15 a_n2686_8422.n8 1.16414
R6816 a_n2686_8422.n50 a_n2686_8422.n43 1.16414
R6817 a_n2686_8422.n197 a_n2686_8422.n165 0.573776
R6818 a_n2686_8422.n165 a_n2686_8422.n163 0.573776
R6819 a_n2686_8422.n131 a_n2686_8422.n99 0.573776
R6820 a_n2686_8422.n66 a_n2686_8422.n34 0.573776
R6821 a_n2686_8422.n34 a_n2686_8422.n32 0.573776
R6822 a_n2686_8422.n265 a_n2686_8422.n231 0.573776
R6823 a_n2686_8422.n265 a_n2686_8422.n264 0.573776
R6824 a_n2686_8422.n244 a_n2686_8422.n243 0.388379
R6825 a_n2686_8422.n212 a_n2686_8422.n211 0.388379
R6826 a_n2686_8422.n79 a_n2686_8422.n78 0.388379
R6827 a_n2686_8422.n112 a_n2686_8422.n111 0.388379
R6828 a_n2686_8422.n144 a_n2686_8422.n143 0.388379
R6829 a_n2686_8422.n178 a_n2686_8422.n177 0.388379
R6830 a_n2686_8422.n12 a_n2686_8422.n11 0.388379
R6831 a_n2686_8422.n47 a_n2686_8422.n46 0.388379
R6832 a_n2686_8422.n261 a_n2686_8422.n233 0.155672
R6833 a_n2686_8422.n254 a_n2686_8422.n233 0.155672
R6834 a_n2686_8422.n254 a_n2686_8422.n253 0.155672
R6835 a_n2686_8422.n253 a_n2686_8422.n237 0.155672
R6836 a_n2686_8422.n246 a_n2686_8422.n237 0.155672
R6837 a_n2686_8422.n246 a_n2686_8422.n245 0.155672
R6838 a_n2686_8422.n229 a_n2686_8422.n201 0.155672
R6839 a_n2686_8422.n222 a_n2686_8422.n201 0.155672
R6840 a_n2686_8422.n222 a_n2686_8422.n221 0.155672
R6841 a_n2686_8422.n221 a_n2686_8422.n205 0.155672
R6842 a_n2686_8422.n214 a_n2686_8422.n205 0.155672
R6843 a_n2686_8422.n214 a_n2686_8422.n213 0.155672
R6844 a_n2686_8422.n96 a_n2686_8422.n68 0.155672
R6845 a_n2686_8422.n89 a_n2686_8422.n68 0.155672
R6846 a_n2686_8422.n89 a_n2686_8422.n88 0.155672
R6847 a_n2686_8422.n88 a_n2686_8422.n72 0.155672
R6848 a_n2686_8422.n81 a_n2686_8422.n72 0.155672
R6849 a_n2686_8422.n81 a_n2686_8422.n80 0.155672
R6850 a_n2686_8422.n129 a_n2686_8422.n101 0.155672
R6851 a_n2686_8422.n122 a_n2686_8422.n101 0.155672
R6852 a_n2686_8422.n122 a_n2686_8422.n121 0.155672
R6853 a_n2686_8422.n121 a_n2686_8422.n105 0.155672
R6854 a_n2686_8422.n114 a_n2686_8422.n105 0.155672
R6855 a_n2686_8422.n114 a_n2686_8422.n113 0.155672
R6856 a_n2686_8422.n161 a_n2686_8422.n133 0.155672
R6857 a_n2686_8422.n154 a_n2686_8422.n133 0.155672
R6858 a_n2686_8422.n154 a_n2686_8422.n153 0.155672
R6859 a_n2686_8422.n153 a_n2686_8422.n137 0.155672
R6860 a_n2686_8422.n146 a_n2686_8422.n137 0.155672
R6861 a_n2686_8422.n146 a_n2686_8422.n145 0.155672
R6862 a_n2686_8422.n195 a_n2686_8422.n167 0.155672
R6863 a_n2686_8422.n188 a_n2686_8422.n167 0.155672
R6864 a_n2686_8422.n188 a_n2686_8422.n187 0.155672
R6865 a_n2686_8422.n187 a_n2686_8422.n171 0.155672
R6866 a_n2686_8422.n180 a_n2686_8422.n171 0.155672
R6867 a_n2686_8422.n180 a_n2686_8422.n179 0.155672
R6868 a_n2686_8422.n163 a_n2686_8422.n131 0.155672
R6869 a_n2686_8422.n29 a_n2686_8422.n1 0.155672
R6870 a_n2686_8422.n22 a_n2686_8422.n1 0.155672
R6871 a_n2686_8422.n22 a_n2686_8422.n21 0.155672
R6872 a_n2686_8422.n21 a_n2686_8422.n5 0.155672
R6873 a_n2686_8422.n14 a_n2686_8422.n5 0.155672
R6874 a_n2686_8422.n14 a_n2686_8422.n13 0.155672
R6875 a_n2686_8422.n64 a_n2686_8422.n36 0.155672
R6876 a_n2686_8422.n57 a_n2686_8422.n36 0.155672
R6877 a_n2686_8422.n57 a_n2686_8422.n56 0.155672
R6878 a_n2686_8422.n56 a_n2686_8422.n40 0.155672
R6879 a_n2686_8422.n49 a_n2686_8422.n40 0.155672
R6880 a_n2686_8422.n49 a_n2686_8422.n48 0.155672
R6881 GND.n5313 GND.n5312 1759.94
R6882 GND.n4753 GND.n4752 1177.98
R6883 GND.n4253 GND.n1776 766.379
R6884 GND.n3814 GND.n3813 766.379
R6885 GND.n2999 GND.n1401 766.379
R6886 GND.n4536 GND.n1323 766.379
R6887 GND.n1316 GND.n1264 761.573
R6888 GND.n4503 GND.n1262 761.573
R6889 GND.n2577 GND.n1110 761.573
R6890 GND.n2614 GND.n2613 761.573
R6891 GND.n4213 GND.n1852 761.573
R6892 GND.n4216 GND.n1820 761.573
R6893 GND.n5569 GND.n5568 761.573
R6894 GND.n5631 GND.n461 761.573
R6895 GND.n5629 GND.n494 742.355
R6896 GND.n5574 GND.n5573 742.355
R6897 GND.n3644 GND.n1857 742.355
R6898 GND.n3590 GND.n3589 742.355
R6899 GND.n4599 GND.n1266 742.355
R6900 GND.n4601 GND.n1260 742.355
R6901 GND.n4682 GND.n4681 742.355
R6902 GND.n4750 GND.n1114 742.355
R6903 GND.n4883 GND.n954 689.5
R6904 GND.n5314 GND.n700 689.5
R6905 GND.n5481 GND.n5480 689.5
R6906 GND.n2541 GND.n2505 689.5
R6907 GND.n4884 GND.n4883 585
R6908 GND.n4883 GND.n4882 585
R6909 GND.n958 GND.n957 585
R6910 GND.n4881 GND.n958 585
R6911 GND.n4879 GND.n4878 585
R6912 GND.n4880 GND.n4879 585
R6913 GND.n4877 GND.n960 585
R6914 GND.n960 GND.n959 585
R6915 GND.n4876 GND.n4875 585
R6916 GND.n4875 GND.n4874 585
R6917 GND.n965 GND.n964 585
R6918 GND.n4873 GND.n965 585
R6919 GND.n4871 GND.n4870 585
R6920 GND.n4872 GND.n4871 585
R6921 GND.n4869 GND.n967 585
R6922 GND.n967 GND.n966 585
R6923 GND.n4868 GND.n4867 585
R6924 GND.n4867 GND.n4866 585
R6925 GND.n973 GND.n972 585
R6926 GND.n4865 GND.n973 585
R6927 GND.n4863 GND.n4862 585
R6928 GND.n4864 GND.n4863 585
R6929 GND.n4861 GND.n975 585
R6930 GND.n975 GND.n974 585
R6931 GND.n4860 GND.n4859 585
R6932 GND.n4859 GND.n4858 585
R6933 GND.n981 GND.n980 585
R6934 GND.n4857 GND.n981 585
R6935 GND.n4855 GND.n4854 585
R6936 GND.n4856 GND.n4855 585
R6937 GND.n4853 GND.n983 585
R6938 GND.n983 GND.n982 585
R6939 GND.n4852 GND.n4851 585
R6940 GND.n4851 GND.n4850 585
R6941 GND.n989 GND.n988 585
R6942 GND.n4849 GND.n989 585
R6943 GND.n4847 GND.n4846 585
R6944 GND.n4848 GND.n4847 585
R6945 GND.n4845 GND.n991 585
R6946 GND.n991 GND.n990 585
R6947 GND.n4844 GND.n4843 585
R6948 GND.n4843 GND.n4842 585
R6949 GND.n997 GND.n996 585
R6950 GND.n4841 GND.n997 585
R6951 GND.n4839 GND.n4838 585
R6952 GND.n4840 GND.n4839 585
R6953 GND.n4837 GND.n999 585
R6954 GND.n999 GND.n998 585
R6955 GND.n4836 GND.n4835 585
R6956 GND.n4835 GND.n4834 585
R6957 GND.n1005 GND.n1004 585
R6958 GND.n4833 GND.n1005 585
R6959 GND.n4831 GND.n4830 585
R6960 GND.n4832 GND.n4831 585
R6961 GND.n4829 GND.n1007 585
R6962 GND.n1007 GND.n1006 585
R6963 GND.n4828 GND.n4827 585
R6964 GND.n4827 GND.n4826 585
R6965 GND.n1013 GND.n1012 585
R6966 GND.n4825 GND.n1013 585
R6967 GND.n4823 GND.n4822 585
R6968 GND.n4824 GND.n4823 585
R6969 GND.n4821 GND.n1015 585
R6970 GND.n1015 GND.n1014 585
R6971 GND.n4820 GND.n4819 585
R6972 GND.n4819 GND.n4818 585
R6973 GND.n1021 GND.n1020 585
R6974 GND.n4817 GND.n1021 585
R6975 GND.n4815 GND.n4814 585
R6976 GND.n4816 GND.n4815 585
R6977 GND.n4813 GND.n1023 585
R6978 GND.n1023 GND.n1022 585
R6979 GND.n4812 GND.n4811 585
R6980 GND.n4811 GND.n4810 585
R6981 GND.n1029 GND.n1028 585
R6982 GND.n4809 GND.n1029 585
R6983 GND.n4807 GND.n4806 585
R6984 GND.n4808 GND.n4807 585
R6985 GND.n4805 GND.n1031 585
R6986 GND.n1031 GND.n1030 585
R6987 GND.n4804 GND.n4803 585
R6988 GND.n4803 GND.n4802 585
R6989 GND.n1037 GND.n1036 585
R6990 GND.n4801 GND.n1037 585
R6991 GND.n4799 GND.n4798 585
R6992 GND.n4800 GND.n4799 585
R6993 GND.n4797 GND.n1039 585
R6994 GND.n1039 GND.n1038 585
R6995 GND.n4796 GND.n4795 585
R6996 GND.n4795 GND.n4794 585
R6997 GND.n1045 GND.n1044 585
R6998 GND.n4793 GND.n1045 585
R6999 GND.n4791 GND.n4790 585
R7000 GND.n4792 GND.n4791 585
R7001 GND.n4789 GND.n1047 585
R7002 GND.n1047 GND.n1046 585
R7003 GND.n4788 GND.n4787 585
R7004 GND.n4787 GND.n4786 585
R7005 GND.n1053 GND.n1052 585
R7006 GND.n4785 GND.n1053 585
R7007 GND.n4783 GND.n4782 585
R7008 GND.n4784 GND.n4783 585
R7009 GND.n4781 GND.n1055 585
R7010 GND.n1055 GND.n1054 585
R7011 GND.n4780 GND.n4779 585
R7012 GND.n4779 GND.n4778 585
R7013 GND.n1061 GND.n1060 585
R7014 GND.n4777 GND.n1061 585
R7015 GND.n4775 GND.n4774 585
R7016 GND.n4776 GND.n4775 585
R7017 GND.n4773 GND.n1063 585
R7018 GND.n1063 GND.n1062 585
R7019 GND.n4772 GND.n4771 585
R7020 GND.n4771 GND.n4770 585
R7021 GND.n1069 GND.n1068 585
R7022 GND.n4769 GND.n1069 585
R7023 GND.n4767 GND.n4766 585
R7024 GND.n4768 GND.n4767 585
R7025 GND.n4765 GND.n1071 585
R7026 GND.n1071 GND.n1070 585
R7027 GND.n4764 GND.n4763 585
R7028 GND.n4763 GND.n4762 585
R7029 GND.n1077 GND.n1076 585
R7030 GND.n4761 GND.n1077 585
R7031 GND.n4759 GND.n4758 585
R7032 GND.n4760 GND.n4759 585
R7033 GND.n4757 GND.n1079 585
R7034 GND.n1079 GND.n1078 585
R7035 GND.n4756 GND.n4755 585
R7036 GND.n4755 GND.n4754 585
R7037 GND.n1085 GND.n1084 585
R7038 GND.n4753 GND.n1085 585
R7039 GND.n955 GND.n954 585
R7040 GND.n954 GND.n953 585
R7041 GND.n4889 GND.n4888 585
R7042 GND.n4890 GND.n4889 585
R7043 GND.n952 GND.n951 585
R7044 GND.n4891 GND.n952 585
R7045 GND.n4894 GND.n4893 585
R7046 GND.n4893 GND.n4892 585
R7047 GND.n949 GND.n948 585
R7048 GND.n948 GND.n947 585
R7049 GND.n4899 GND.n4898 585
R7050 GND.n4900 GND.n4899 585
R7051 GND.n946 GND.n945 585
R7052 GND.n4901 GND.n946 585
R7053 GND.n4904 GND.n4903 585
R7054 GND.n4903 GND.n4902 585
R7055 GND.n943 GND.n942 585
R7056 GND.n942 GND.n941 585
R7057 GND.n4909 GND.n4908 585
R7058 GND.n4910 GND.n4909 585
R7059 GND.n940 GND.n939 585
R7060 GND.n4911 GND.n940 585
R7061 GND.n4914 GND.n4913 585
R7062 GND.n4913 GND.n4912 585
R7063 GND.n937 GND.n936 585
R7064 GND.n936 GND.n935 585
R7065 GND.n4919 GND.n4918 585
R7066 GND.n4920 GND.n4919 585
R7067 GND.n934 GND.n933 585
R7068 GND.n4921 GND.n934 585
R7069 GND.n4924 GND.n4923 585
R7070 GND.n4923 GND.n4922 585
R7071 GND.n931 GND.n930 585
R7072 GND.n930 GND.n929 585
R7073 GND.n4929 GND.n4928 585
R7074 GND.n4930 GND.n4929 585
R7075 GND.n928 GND.n927 585
R7076 GND.n4931 GND.n928 585
R7077 GND.n4934 GND.n4933 585
R7078 GND.n4933 GND.n4932 585
R7079 GND.n925 GND.n924 585
R7080 GND.n924 GND.n923 585
R7081 GND.n4939 GND.n4938 585
R7082 GND.n4940 GND.n4939 585
R7083 GND.n922 GND.n921 585
R7084 GND.n4941 GND.n922 585
R7085 GND.n4944 GND.n4943 585
R7086 GND.n4943 GND.n4942 585
R7087 GND.n919 GND.n918 585
R7088 GND.n918 GND.n917 585
R7089 GND.n4949 GND.n4948 585
R7090 GND.n4950 GND.n4949 585
R7091 GND.n916 GND.n915 585
R7092 GND.n4951 GND.n916 585
R7093 GND.n4954 GND.n4953 585
R7094 GND.n4953 GND.n4952 585
R7095 GND.n913 GND.n912 585
R7096 GND.n912 GND.n911 585
R7097 GND.n4959 GND.n4958 585
R7098 GND.n4960 GND.n4959 585
R7099 GND.n910 GND.n909 585
R7100 GND.n4961 GND.n910 585
R7101 GND.n4964 GND.n4963 585
R7102 GND.n4963 GND.n4962 585
R7103 GND.n907 GND.n906 585
R7104 GND.n906 GND.n905 585
R7105 GND.n4969 GND.n4968 585
R7106 GND.n4970 GND.n4969 585
R7107 GND.n904 GND.n903 585
R7108 GND.n4971 GND.n904 585
R7109 GND.n4974 GND.n4973 585
R7110 GND.n4973 GND.n4972 585
R7111 GND.n901 GND.n900 585
R7112 GND.n900 GND.n899 585
R7113 GND.n4979 GND.n4978 585
R7114 GND.n4980 GND.n4979 585
R7115 GND.n898 GND.n897 585
R7116 GND.n4981 GND.n898 585
R7117 GND.n4984 GND.n4983 585
R7118 GND.n4983 GND.n4982 585
R7119 GND.n895 GND.n894 585
R7120 GND.n894 GND.n893 585
R7121 GND.n4989 GND.n4988 585
R7122 GND.n4990 GND.n4989 585
R7123 GND.n892 GND.n891 585
R7124 GND.n4991 GND.n892 585
R7125 GND.n4994 GND.n4993 585
R7126 GND.n4993 GND.n4992 585
R7127 GND.n889 GND.n888 585
R7128 GND.n888 GND.n887 585
R7129 GND.n4999 GND.n4998 585
R7130 GND.n5000 GND.n4999 585
R7131 GND.n886 GND.n885 585
R7132 GND.n5001 GND.n886 585
R7133 GND.n5004 GND.n5003 585
R7134 GND.n5003 GND.n5002 585
R7135 GND.n883 GND.n882 585
R7136 GND.n882 GND.n881 585
R7137 GND.n5009 GND.n5008 585
R7138 GND.n5010 GND.n5009 585
R7139 GND.n880 GND.n879 585
R7140 GND.n5011 GND.n880 585
R7141 GND.n5014 GND.n5013 585
R7142 GND.n5013 GND.n5012 585
R7143 GND.n877 GND.n876 585
R7144 GND.n876 GND.n875 585
R7145 GND.n5019 GND.n5018 585
R7146 GND.n5020 GND.n5019 585
R7147 GND.n874 GND.n873 585
R7148 GND.n5021 GND.n874 585
R7149 GND.n5024 GND.n5023 585
R7150 GND.n5023 GND.n5022 585
R7151 GND.n871 GND.n870 585
R7152 GND.n870 GND.n869 585
R7153 GND.n5029 GND.n5028 585
R7154 GND.n5030 GND.n5029 585
R7155 GND.n868 GND.n867 585
R7156 GND.n5031 GND.n868 585
R7157 GND.n5034 GND.n5033 585
R7158 GND.n5033 GND.n5032 585
R7159 GND.n865 GND.n864 585
R7160 GND.n864 GND.n863 585
R7161 GND.n5039 GND.n5038 585
R7162 GND.n5040 GND.n5039 585
R7163 GND.n862 GND.n861 585
R7164 GND.n5041 GND.n862 585
R7165 GND.n5044 GND.n5043 585
R7166 GND.n5043 GND.n5042 585
R7167 GND.n859 GND.n858 585
R7168 GND.n858 GND.n857 585
R7169 GND.n5049 GND.n5048 585
R7170 GND.n5050 GND.n5049 585
R7171 GND.n856 GND.n855 585
R7172 GND.n5051 GND.n856 585
R7173 GND.n5054 GND.n5053 585
R7174 GND.n5053 GND.n5052 585
R7175 GND.n853 GND.n852 585
R7176 GND.n852 GND.n851 585
R7177 GND.n5059 GND.n5058 585
R7178 GND.n5060 GND.n5059 585
R7179 GND.n850 GND.n849 585
R7180 GND.n5061 GND.n850 585
R7181 GND.n5064 GND.n5063 585
R7182 GND.n5063 GND.n5062 585
R7183 GND.n847 GND.n846 585
R7184 GND.n846 GND.n845 585
R7185 GND.n5069 GND.n5068 585
R7186 GND.n5070 GND.n5069 585
R7187 GND.n844 GND.n843 585
R7188 GND.n5071 GND.n844 585
R7189 GND.n5074 GND.n5073 585
R7190 GND.n5073 GND.n5072 585
R7191 GND.n841 GND.n840 585
R7192 GND.n840 GND.n839 585
R7193 GND.n5079 GND.n5078 585
R7194 GND.n5080 GND.n5079 585
R7195 GND.n838 GND.n837 585
R7196 GND.n5081 GND.n838 585
R7197 GND.n5084 GND.n5083 585
R7198 GND.n5083 GND.n5082 585
R7199 GND.n835 GND.n834 585
R7200 GND.n834 GND.n833 585
R7201 GND.n5089 GND.n5088 585
R7202 GND.n5090 GND.n5089 585
R7203 GND.n832 GND.n831 585
R7204 GND.n5091 GND.n832 585
R7205 GND.n5094 GND.n5093 585
R7206 GND.n5093 GND.n5092 585
R7207 GND.n829 GND.n828 585
R7208 GND.n828 GND.n827 585
R7209 GND.n5099 GND.n5098 585
R7210 GND.n5100 GND.n5099 585
R7211 GND.n826 GND.n825 585
R7212 GND.n5101 GND.n826 585
R7213 GND.n5104 GND.n5103 585
R7214 GND.n5103 GND.n5102 585
R7215 GND.n823 GND.n822 585
R7216 GND.n822 GND.n821 585
R7217 GND.n5109 GND.n5108 585
R7218 GND.n5110 GND.n5109 585
R7219 GND.n820 GND.n819 585
R7220 GND.n5111 GND.n820 585
R7221 GND.n5114 GND.n5113 585
R7222 GND.n5113 GND.n5112 585
R7223 GND.n817 GND.n816 585
R7224 GND.n816 GND.n815 585
R7225 GND.n5119 GND.n5118 585
R7226 GND.n5120 GND.n5119 585
R7227 GND.n814 GND.n813 585
R7228 GND.n5121 GND.n814 585
R7229 GND.n5124 GND.n5123 585
R7230 GND.n5123 GND.n5122 585
R7231 GND.n811 GND.n810 585
R7232 GND.n810 GND.n809 585
R7233 GND.n5129 GND.n5128 585
R7234 GND.n5130 GND.n5129 585
R7235 GND.n808 GND.n807 585
R7236 GND.n5131 GND.n808 585
R7237 GND.n5134 GND.n5133 585
R7238 GND.n5133 GND.n5132 585
R7239 GND.n805 GND.n804 585
R7240 GND.n804 GND.n803 585
R7241 GND.n5139 GND.n5138 585
R7242 GND.n5140 GND.n5139 585
R7243 GND.n802 GND.n801 585
R7244 GND.n5141 GND.n802 585
R7245 GND.n5144 GND.n5143 585
R7246 GND.n5143 GND.n5142 585
R7247 GND.n799 GND.n798 585
R7248 GND.n798 GND.n797 585
R7249 GND.n5149 GND.n5148 585
R7250 GND.n5150 GND.n5149 585
R7251 GND.n796 GND.n795 585
R7252 GND.n5151 GND.n796 585
R7253 GND.n5154 GND.n5153 585
R7254 GND.n5153 GND.n5152 585
R7255 GND.n793 GND.n792 585
R7256 GND.n792 GND.n791 585
R7257 GND.n5159 GND.n5158 585
R7258 GND.n5160 GND.n5159 585
R7259 GND.n790 GND.n789 585
R7260 GND.n5161 GND.n790 585
R7261 GND.n5164 GND.n5163 585
R7262 GND.n5163 GND.n5162 585
R7263 GND.n787 GND.n786 585
R7264 GND.n786 GND.n785 585
R7265 GND.n5169 GND.n5168 585
R7266 GND.n5170 GND.n5169 585
R7267 GND.n784 GND.n783 585
R7268 GND.n5171 GND.n784 585
R7269 GND.n5174 GND.n5173 585
R7270 GND.n5173 GND.n5172 585
R7271 GND.n781 GND.n780 585
R7272 GND.n780 GND.n779 585
R7273 GND.n5179 GND.n5178 585
R7274 GND.n5180 GND.n5179 585
R7275 GND.n778 GND.n777 585
R7276 GND.n5181 GND.n778 585
R7277 GND.n5184 GND.n5183 585
R7278 GND.n5183 GND.n5182 585
R7279 GND.n775 GND.n774 585
R7280 GND.n774 GND.n773 585
R7281 GND.n5189 GND.n5188 585
R7282 GND.n5190 GND.n5189 585
R7283 GND.n772 GND.n771 585
R7284 GND.n5191 GND.n772 585
R7285 GND.n5194 GND.n5193 585
R7286 GND.n5193 GND.n5192 585
R7287 GND.n769 GND.n768 585
R7288 GND.n768 GND.n767 585
R7289 GND.n5199 GND.n5198 585
R7290 GND.n5200 GND.n5199 585
R7291 GND.n766 GND.n765 585
R7292 GND.n5201 GND.n766 585
R7293 GND.n5204 GND.n5203 585
R7294 GND.n5203 GND.n5202 585
R7295 GND.n763 GND.n762 585
R7296 GND.n762 GND.n761 585
R7297 GND.n5209 GND.n5208 585
R7298 GND.n5210 GND.n5209 585
R7299 GND.n760 GND.n759 585
R7300 GND.n5211 GND.n760 585
R7301 GND.n5214 GND.n5213 585
R7302 GND.n5213 GND.n5212 585
R7303 GND.n757 GND.n756 585
R7304 GND.n756 GND.n755 585
R7305 GND.n5219 GND.n5218 585
R7306 GND.n5220 GND.n5219 585
R7307 GND.n754 GND.n753 585
R7308 GND.n5221 GND.n754 585
R7309 GND.n5224 GND.n5223 585
R7310 GND.n5223 GND.n5222 585
R7311 GND.n751 GND.n750 585
R7312 GND.n750 GND.n749 585
R7313 GND.n5229 GND.n5228 585
R7314 GND.n5230 GND.n5229 585
R7315 GND.n748 GND.n747 585
R7316 GND.n5231 GND.n748 585
R7317 GND.n5234 GND.n5233 585
R7318 GND.n5233 GND.n5232 585
R7319 GND.n745 GND.n744 585
R7320 GND.n744 GND.n743 585
R7321 GND.n5239 GND.n5238 585
R7322 GND.n5240 GND.n5239 585
R7323 GND.n742 GND.n741 585
R7324 GND.n5241 GND.n742 585
R7325 GND.n5244 GND.n5243 585
R7326 GND.n5243 GND.n5242 585
R7327 GND.n739 GND.n738 585
R7328 GND.n738 GND.n737 585
R7329 GND.n5249 GND.n5248 585
R7330 GND.n5250 GND.n5249 585
R7331 GND.n736 GND.n735 585
R7332 GND.n5251 GND.n736 585
R7333 GND.n5254 GND.n5253 585
R7334 GND.n5253 GND.n5252 585
R7335 GND.n733 GND.n732 585
R7336 GND.n732 GND.n731 585
R7337 GND.n5259 GND.n5258 585
R7338 GND.n5260 GND.n5259 585
R7339 GND.n730 GND.n729 585
R7340 GND.n5261 GND.n730 585
R7341 GND.n5264 GND.n5263 585
R7342 GND.n5263 GND.n5262 585
R7343 GND.n727 GND.n726 585
R7344 GND.n726 GND.n725 585
R7345 GND.n5269 GND.n5268 585
R7346 GND.n5270 GND.n5269 585
R7347 GND.n724 GND.n723 585
R7348 GND.n5271 GND.n724 585
R7349 GND.n5274 GND.n5273 585
R7350 GND.n5273 GND.n5272 585
R7351 GND.n721 GND.n720 585
R7352 GND.n720 GND.n719 585
R7353 GND.n5279 GND.n5278 585
R7354 GND.n5280 GND.n5279 585
R7355 GND.n718 GND.n717 585
R7356 GND.n5281 GND.n718 585
R7357 GND.n5284 GND.n5283 585
R7358 GND.n5283 GND.n5282 585
R7359 GND.n715 GND.n714 585
R7360 GND.n714 GND.n713 585
R7361 GND.n5289 GND.n5288 585
R7362 GND.n5290 GND.n5289 585
R7363 GND.n712 GND.n711 585
R7364 GND.n5291 GND.n712 585
R7365 GND.n5294 GND.n5293 585
R7366 GND.n5293 GND.n5292 585
R7367 GND.n709 GND.n708 585
R7368 GND.n708 GND.n707 585
R7369 GND.n5299 GND.n5298 585
R7370 GND.n5300 GND.n5299 585
R7371 GND.n706 GND.n705 585
R7372 GND.n5301 GND.n706 585
R7373 GND.n5304 GND.n5303 585
R7374 GND.n5303 GND.n5302 585
R7375 GND.n703 GND.n702 585
R7376 GND.n702 GND.n701 585
R7377 GND.n5310 GND.n5309 585
R7378 GND.n5311 GND.n5310 585
R7379 GND.n5308 GND.n700 585
R7380 GND.n5312 GND.n700 585
R7381 GND.n602 GND.n601 585
R7382 GND.n601 GND.n476 585
R7383 GND.n5475 GND.n5474 585
R7384 GND.n5474 GND.n5473 585
R7385 GND.n605 GND.n604 585
R7386 GND.n5472 GND.n605 585
R7387 GND.n5470 GND.n5469 585
R7388 GND.n5471 GND.n5470 585
R7389 GND.n608 GND.n607 585
R7390 GND.n607 GND.n606 585
R7391 GND.n5465 GND.n5464 585
R7392 GND.n5464 GND.n5463 585
R7393 GND.n611 GND.n610 585
R7394 GND.n5462 GND.n611 585
R7395 GND.n5460 GND.n5459 585
R7396 GND.n5461 GND.n5460 585
R7397 GND.n614 GND.n613 585
R7398 GND.n613 GND.n612 585
R7399 GND.n5455 GND.n5454 585
R7400 GND.n5454 GND.n5453 585
R7401 GND.n617 GND.n616 585
R7402 GND.n5452 GND.n617 585
R7403 GND.n5450 GND.n5449 585
R7404 GND.n5451 GND.n5450 585
R7405 GND.n620 GND.n619 585
R7406 GND.n619 GND.n618 585
R7407 GND.n5445 GND.n5444 585
R7408 GND.n5444 GND.n5443 585
R7409 GND.n623 GND.n622 585
R7410 GND.n5442 GND.n623 585
R7411 GND.n5440 GND.n5439 585
R7412 GND.n5441 GND.n5440 585
R7413 GND.n626 GND.n625 585
R7414 GND.n625 GND.n624 585
R7415 GND.n5435 GND.n5434 585
R7416 GND.n5434 GND.n5433 585
R7417 GND.n629 GND.n628 585
R7418 GND.n5432 GND.n629 585
R7419 GND.n5430 GND.n5429 585
R7420 GND.n5431 GND.n5430 585
R7421 GND.n632 GND.n631 585
R7422 GND.n631 GND.n630 585
R7423 GND.n5425 GND.n5424 585
R7424 GND.n5424 GND.n5423 585
R7425 GND.n635 GND.n634 585
R7426 GND.n5422 GND.n635 585
R7427 GND.n5420 GND.n5419 585
R7428 GND.n5421 GND.n5420 585
R7429 GND.n638 GND.n637 585
R7430 GND.n637 GND.n636 585
R7431 GND.n5415 GND.n5414 585
R7432 GND.n5414 GND.n5413 585
R7433 GND.n641 GND.n640 585
R7434 GND.n5412 GND.n641 585
R7435 GND.n5410 GND.n5409 585
R7436 GND.n5411 GND.n5410 585
R7437 GND.n644 GND.n643 585
R7438 GND.n643 GND.n642 585
R7439 GND.n5405 GND.n5404 585
R7440 GND.n5404 GND.n5403 585
R7441 GND.n647 GND.n646 585
R7442 GND.n5402 GND.n647 585
R7443 GND.n5400 GND.n5399 585
R7444 GND.n5401 GND.n5400 585
R7445 GND.n650 GND.n649 585
R7446 GND.n649 GND.n648 585
R7447 GND.n5395 GND.n5394 585
R7448 GND.n5394 GND.n5393 585
R7449 GND.n653 GND.n652 585
R7450 GND.n5392 GND.n653 585
R7451 GND.n5390 GND.n5389 585
R7452 GND.n5391 GND.n5390 585
R7453 GND.n656 GND.n655 585
R7454 GND.n655 GND.n654 585
R7455 GND.n5385 GND.n5384 585
R7456 GND.n5384 GND.n5383 585
R7457 GND.n659 GND.n658 585
R7458 GND.n5382 GND.n659 585
R7459 GND.n5380 GND.n5379 585
R7460 GND.n5381 GND.n5380 585
R7461 GND.n662 GND.n661 585
R7462 GND.n661 GND.n660 585
R7463 GND.n5375 GND.n5374 585
R7464 GND.n5374 GND.n5373 585
R7465 GND.n665 GND.n664 585
R7466 GND.n5372 GND.n665 585
R7467 GND.n5370 GND.n5369 585
R7468 GND.n5371 GND.n5370 585
R7469 GND.n668 GND.n667 585
R7470 GND.n667 GND.n666 585
R7471 GND.n5365 GND.n5364 585
R7472 GND.n5364 GND.n5363 585
R7473 GND.n671 GND.n670 585
R7474 GND.n5362 GND.n671 585
R7475 GND.n5360 GND.n5359 585
R7476 GND.n5361 GND.n5360 585
R7477 GND.n674 GND.n673 585
R7478 GND.n673 GND.n672 585
R7479 GND.n5355 GND.n5354 585
R7480 GND.n5354 GND.n5353 585
R7481 GND.n677 GND.n676 585
R7482 GND.n5352 GND.n677 585
R7483 GND.n5350 GND.n5349 585
R7484 GND.n5351 GND.n5350 585
R7485 GND.n680 GND.n679 585
R7486 GND.n679 GND.n678 585
R7487 GND.n5345 GND.n5344 585
R7488 GND.n5344 GND.n5343 585
R7489 GND.n683 GND.n682 585
R7490 GND.n5342 GND.n683 585
R7491 GND.n5340 GND.n5339 585
R7492 GND.n5341 GND.n5340 585
R7493 GND.n686 GND.n685 585
R7494 GND.n685 GND.n684 585
R7495 GND.n5335 GND.n5334 585
R7496 GND.n5334 GND.n5333 585
R7497 GND.n689 GND.n688 585
R7498 GND.n5332 GND.n689 585
R7499 GND.n5330 GND.n5329 585
R7500 GND.n5331 GND.n5330 585
R7501 GND.n692 GND.n691 585
R7502 GND.n691 GND.n690 585
R7503 GND.n5325 GND.n5324 585
R7504 GND.n5324 GND.n5323 585
R7505 GND.n695 GND.n694 585
R7506 GND.n5322 GND.n695 585
R7507 GND.n5320 GND.n5319 585
R7508 GND.n5321 GND.n5320 585
R7509 GND.n698 GND.n697 585
R7510 GND.n697 GND.n696 585
R7511 GND.n5315 GND.n5314 585
R7512 GND.n5314 GND.n5313 585
R7513 GND.n4206 GND.n1776 585
R7514 GND.n1776 GND.n1760 585
R7515 GND.n1746 GND.n1745 585
R7516 GND.n1748 GND.n1746 585
R7517 GND.n4265 GND.n4264 585
R7518 GND.n4264 GND.n4263 585
R7519 GND.n4266 GND.n1738 585
R7520 GND.n3805 GND.n1738 585
R7521 GND.n4268 GND.n4267 585
R7522 GND.n4269 GND.n4268 585
R7523 GND.n1739 GND.n1737 585
R7524 GND.n1737 GND.n1734 585
R7525 GND.n1719 GND.n1718 585
R7526 GND.n1722 GND.n1719 585
R7527 GND.n4279 GND.n4278 585
R7528 GND.n4278 GND.n4277 585
R7529 GND.n4280 GND.n1711 585
R7530 GND.n2171 GND.n1711 585
R7531 GND.n4282 GND.n4281 585
R7532 GND.n4283 GND.n4282 585
R7533 GND.n1712 GND.n1710 585
R7534 GND.n1710 GND.n1707 585
R7535 GND.n1695 GND.n1694 585
R7536 GND.n1697 GND.n1695 585
R7537 GND.n4293 GND.n4292 585
R7538 GND.n4292 GND.n4291 585
R7539 GND.n4294 GND.n1689 585
R7540 GND.n3757 GND.n1689 585
R7541 GND.n4296 GND.n4295 585
R7542 GND.n4297 GND.n4296 585
R7543 GND.n1677 GND.n1676 585
R7544 GND.n3780 GND.n1677 585
R7545 GND.n4307 GND.n4306 585
R7546 GND.n4306 GND.n4305 585
R7547 GND.n4308 GND.n1666 585
R7548 GND.n3450 GND.n1666 585
R7549 GND.n4310 GND.n4309 585
R7550 GND.n4311 GND.n4310 585
R7551 GND.n1667 GND.n1665 585
R7552 GND.n3441 GND.n1665 585
R7553 GND.n1670 GND.n1669 585
R7554 GND.n1669 GND.n1653 585
R7555 GND.n1642 GND.n1641 585
R7556 GND.n1651 GND.n1642 585
R7557 GND.n4328 GND.n4327 585
R7558 GND.n4327 GND.n4326 585
R7559 GND.n4329 GND.n1631 585
R7560 GND.n3408 GND.n1631 585
R7561 GND.n4331 GND.n4330 585
R7562 GND.n4332 GND.n4331 585
R7563 GND.n1632 GND.n1630 585
R7564 GND.n1630 GND.n1620 585
R7565 GND.n1635 GND.n1634 585
R7566 GND.n1634 GND.n1618 585
R7567 GND.n1602 GND.n1601 585
R7568 GND.n3394 GND.n1602 585
R7569 GND.n4348 GND.n4347 585
R7570 GND.n4347 GND.n4346 585
R7571 GND.n4349 GND.n1588 585
R7572 GND.n2203 GND.n1588 585
R7573 GND.n4351 GND.n4350 585
R7574 GND.n4352 GND.n4351 585
R7575 GND.n1589 GND.n1587 585
R7576 GND.n1587 GND.n1577 585
R7577 GND.n1595 GND.n1594 585
R7578 GND.n1594 GND.n1575 585
R7579 GND.n1593 GND.n1592 585
R7580 GND.n1593 GND.n1561 585
R7581 GND.n1549 GND.n1548 585
R7582 GND.n1559 GND.n1549 585
R7583 GND.n4376 GND.n4375 585
R7584 GND.n4375 GND.n4374 585
R7585 GND.n4377 GND.n1543 585
R7586 GND.n3349 GND.n1543 585
R7587 GND.n4379 GND.n4378 585
R7588 GND.n4380 GND.n4379 585
R7589 GND.n1544 GND.n1542 585
R7590 GND.n3320 GND.n1542 585
R7591 GND.n3285 GND.n3284 585
R7592 GND.n3285 GND.n1532 585
R7593 GND.n3287 GND.n3286 585
R7594 GND.n3286 GND.n1530 585
R7595 GND.n3288 GND.n1524 585
R7596 GND.n4394 GND.n1524 585
R7597 GND.n3290 GND.n3289 585
R7598 GND.n3291 GND.n3290 585
R7599 GND.n2223 GND.n2222 585
R7600 GND.n3256 GND.n2222 585
R7601 GND.n3276 GND.n3275 585
R7602 GND.n3275 GND.n1510 585
R7603 GND.n3274 GND.n2225 585
R7604 GND.n3274 GND.n1504 585
R7605 GND.n3273 GND.n2227 585
R7606 GND.n3273 GND.n3272 585
R7607 GND.n3243 GND.n2226 585
R7608 GND.n2232 GND.n2226 585
R7609 GND.n3244 GND.n3235 585
R7610 GND.n3235 GND.n1492 585
R7611 GND.n3246 GND.n3245 585
R7612 GND.n3247 GND.n3246 585
R7613 GND.n3236 GND.n3234 585
R7614 GND.n3234 GND.n3233 585
R7615 GND.n1471 GND.n1470 585
R7616 GND.n2241 GND.n1471 585
R7617 GND.n4432 GND.n4431 585
R7618 GND.n4431 GND.n4430 585
R7619 GND.n4433 GND.n1463 585
R7620 GND.n3035 GND.n1463 585
R7621 GND.n4435 GND.n4434 585
R7622 GND.n4436 GND.n4435 585
R7623 GND.n1464 GND.n1462 585
R7624 GND.n1462 GND.n1459 585
R7625 GND.n1444 GND.n1443 585
R7626 GND.n1447 GND.n1444 585
R7627 GND.n4446 GND.n4445 585
R7628 GND.n4445 GND.n4444 585
R7629 GND.n4447 GND.n1436 585
R7630 GND.n2269 GND.n1436 585
R7631 GND.n4449 GND.n4448 585
R7632 GND.n4450 GND.n4449 585
R7633 GND.n1437 GND.n1435 585
R7634 GND.n1435 GND.n1432 585
R7635 GND.n1411 GND.n1410 585
R7636 GND.n1414 GND.n1411 585
R7637 GND.n4460 GND.n4459 585
R7638 GND.n4459 GND.n4458 585
R7639 GND.n4461 GND.n1404 585
R7640 GND.n3005 GND.n1404 585
R7641 GND.n4463 GND.n4462 585
R7642 GND.n4464 GND.n4463 585
R7643 GND.n1405 GND.n1323 585
R7644 GND.n4466 GND.n1323 585
R7645 GND.n4537 GND.n4536 585
R7646 GND.n1324 GND.n1322 585
R7647 GND.n4533 GND.n4532 585
R7648 GND.n4534 GND.n4533 585
R7649 GND.n1341 GND.n1340 585
R7650 GND.n4525 GND.n1350 585
R7651 GND.n4524 GND.n1351 585
R7652 GND.n1358 GND.n1352 585
R7653 GND.n4517 GND.n1359 585
R7654 GND.n4516 GND.n1360 585
R7655 GND.n1362 GND.n1361 585
R7656 GND.n4509 GND.n1368 585
R7657 GND.n4508 GND.n1369 585
R7658 GND.n2282 GND.n1370 585
R7659 GND.n2284 GND.n2283 585
R7660 GND.n2963 GND.n2962 585
R7661 GND.n2965 GND.n2964 585
R7662 GND.n2968 GND.n2967 585
R7663 GND.n2966 GND.n2280 585
R7664 GND.n2973 GND.n2972 585
R7665 GND.n2975 GND.n2974 585
R7666 GND.n2978 GND.n2977 585
R7667 GND.n2976 GND.n2278 585
R7668 GND.n2983 GND.n2982 585
R7669 GND.n2985 GND.n2984 585
R7670 GND.n2991 GND.n2987 585
R7671 GND.n2986 GND.n2276 585
R7672 GND.n2996 GND.n2995 585
R7673 GND.n2998 GND.n2997 585
R7674 GND.n3000 GND.n2999 585
R7675 GND.n3815 GND.n3814 585
R7676 GND.n3816 GND.n2164 585
R7677 GND.n2163 GND.n2161 585
R7678 GND.n3820 GND.n2160 585
R7679 GND.n3822 GND.n2157 585
R7680 GND.n3823 GND.n2156 585
R7681 GND.n2155 GND.n2153 585
R7682 GND.n3827 GND.n2152 585
R7683 GND.n3828 GND.n2151 585
R7684 GND.n3829 GND.n2150 585
R7685 GND.n2149 GND.n2147 585
R7686 GND.n3833 GND.n2146 585
R7687 GND.n3834 GND.n2145 585
R7688 GND.n3835 GND.n2144 585
R7689 GND.n2143 GND.n2142 585
R7690 GND.n1818 GND.n1817 585
R7691 GND.n4220 GND.n1816 585
R7692 GND.n4221 GND.n1815 585
R7693 GND.n1814 GND.n1806 585
R7694 GND.n4228 GND.n1805 585
R7695 GND.n4229 GND.n1804 585
R7696 GND.n1798 GND.n1797 585
R7697 GND.n4236 GND.n1796 585
R7698 GND.n4237 GND.n1795 585
R7699 GND.n1794 GND.n1788 585
R7700 GND.n4244 GND.n1787 585
R7701 GND.n4245 GND.n1786 585
R7702 GND.n1778 GND.n1777 585
R7703 GND.n4253 GND.n4252 585
R7704 GND.n4254 GND.n4253 585
R7705 GND.n3813 GND.n3812 585
R7706 GND.n3813 GND.n1760 585
R7707 GND.n2166 GND.n2165 585
R7708 GND.n2165 GND.n1748 585
R7709 GND.n3808 GND.n1747 585
R7710 GND.n4263 GND.n1747 585
R7711 GND.n3807 GND.n3806 585
R7712 GND.n3806 GND.n3805 585
R7713 GND.n3803 GND.n1735 585
R7714 GND.n4269 GND.n1735 585
R7715 GND.n3797 GND.n2168 585
R7716 GND.n3797 GND.n1734 585
R7717 GND.n3799 GND.n3798 585
R7718 GND.n3798 GND.n1722 585
R7719 GND.n3796 GND.n1721 585
R7720 GND.n4277 GND.n1721 585
R7721 GND.n3795 GND.n2172 585
R7722 GND.n2172 GND.n2171 585
R7723 GND.n2170 GND.n1708 585
R7724 GND.n4283 GND.n1708 585
R7725 GND.n3791 GND.n3790 585
R7726 GND.n3790 GND.n1707 585
R7727 GND.n3789 GND.n3788 585
R7728 GND.n3789 GND.n1697 585
R7729 GND.n3787 GND.n1696 585
R7730 GND.n4291 GND.n1696 585
R7731 GND.n3457 GND.n2174 585
R7732 GND.n3757 GND.n3457 585
R7733 GND.n3783 GND.n1688 585
R7734 GND.n4297 GND.n1688 585
R7735 GND.n3782 GND.n3781 585
R7736 GND.n3781 GND.n3780 585
R7737 GND.n2176 GND.n1679 585
R7738 GND.n4305 GND.n1679 585
R7739 GND.n3449 GND.n3448 585
R7740 GND.n3450 GND.n3449 585
R7741 GND.n2182 GND.n1663 585
R7742 GND.n4311 GND.n1663 585
R7743 GND.n3443 GND.n3442 585
R7744 GND.n3442 GND.n3441 585
R7745 GND.n2185 GND.n2184 585
R7746 GND.n2185 GND.n1653 585
R7747 GND.n3402 GND.n3401 585
R7748 GND.n3401 GND.n1651 585
R7749 GND.n2194 GND.n1643 585
R7750 GND.n4326 GND.n1643 585
R7751 GND.n3407 GND.n3406 585
R7752 GND.n3408 GND.n3407 585
R7753 GND.n2193 GND.n1628 585
R7754 GND.n4332 GND.n1628 585
R7755 GND.n3398 GND.n3397 585
R7756 GND.n3397 GND.n1620 585
R7757 GND.n3396 GND.n2196 585
R7758 GND.n3396 GND.n1618 585
R7759 GND.n3395 GND.n2197 585
R7760 GND.n3395 GND.n3394 585
R7761 GND.n3335 GND.n1604 585
R7762 GND.n4346 GND.n1604 585
R7763 GND.n3336 GND.n3332 585
R7764 GND.n3332 GND.n2203 585
R7765 GND.n3337 GND.n1585 585
R7766 GND.n4352 GND.n1585 585
R7767 GND.n3330 GND.n3329 585
R7768 GND.n3329 GND.n1577 585
R7769 GND.n3341 GND.n3328 585
R7770 GND.n3328 GND.n1575 585
R7771 GND.n3342 GND.n3327 585
R7772 GND.n3327 GND.n1561 585
R7773 GND.n3343 GND.n3326 585
R7774 GND.n3326 GND.n1559 585
R7775 GND.n2212 GND.n1551 585
R7776 GND.n4374 GND.n1551 585
R7777 GND.n3348 GND.n3347 585
R7778 GND.n3349 GND.n3348 585
R7779 GND.n2211 GND.n1540 585
R7780 GND.n4380 GND.n1540 585
R7781 GND.n3322 GND.n3321 585
R7782 GND.n3321 GND.n3320 585
R7783 GND.n2215 GND.n2214 585
R7784 GND.n2215 GND.n1532 585
R7785 GND.n3260 GND.n3259 585
R7786 GND.n3259 GND.n1530 585
R7787 GND.n3258 GND.n1522 585
R7788 GND.n4394 GND.n1522 585
R7789 GND.n3264 GND.n2221 585
R7790 GND.n3291 GND.n2221 585
R7791 GND.n3265 GND.n3257 585
R7792 GND.n3257 GND.n3256 585
R7793 GND.n3266 GND.n3254 585
R7794 GND.n3254 GND.n1510 585
R7795 GND.n2236 GND.n2234 585
R7796 GND.n2234 GND.n1504 585
R7797 GND.n3271 GND.n3270 585
R7798 GND.n3272 GND.n3271 585
R7799 GND.n2235 GND.n2233 585
R7800 GND.n2233 GND.n2232 585
R7801 GND.n3250 GND.n3249 585
R7802 GND.n3249 GND.n1492 585
R7803 GND.n3248 GND.n2238 585
R7804 GND.n3248 GND.n3247 585
R7805 GND.n3028 GND.n2239 585
R7806 GND.n3233 GND.n2239 585
R7807 GND.n3029 GND.n3027 585
R7808 GND.n3027 GND.n2241 585
R7809 GND.n2267 GND.n1473 585
R7810 GND.n4430 GND.n1473 585
R7811 GND.n3034 GND.n3033 585
R7812 GND.n3035 GND.n3034 585
R7813 GND.n2266 GND.n1460 585
R7814 GND.n4436 GND.n1460 585
R7815 GND.n3023 GND.n3022 585
R7816 GND.n3022 GND.n1459 585
R7817 GND.n3021 GND.n3020 585
R7818 GND.n3021 GND.n1447 585
R7819 GND.n3019 GND.n1446 585
R7820 GND.n4444 GND.n1446 585
R7821 GND.n2271 GND.n2270 585
R7822 GND.n2270 GND.n2269 585
R7823 GND.n3015 GND.n1433 585
R7824 GND.n4450 GND.n1433 585
R7825 GND.n3014 GND.n3013 585
R7826 GND.n3013 GND.n1432 585
R7827 GND.n3012 GND.n3011 585
R7828 GND.n3012 GND.n1414 585
R7829 GND.n2273 GND.n1413 585
R7830 GND.n4458 GND.n1413 585
R7831 GND.n3007 GND.n3006 585
R7832 GND.n3006 GND.n3005 585
R7833 GND.n3004 GND.n1402 585
R7834 GND.n4464 GND.n1402 585
R7835 GND.n3003 GND.n1401 585
R7836 GND.n4466 GND.n1401 585
R7837 GND.n2952 GND.n1264 585
R7838 GND.n4600 GND.n1264 585
R7839 GND.n2954 GND.n2953 585
R7840 GND.n2955 GND.n2954 585
R7841 GND.n2951 GND.n1255 585
R7842 GND.n2951 GND.n2950 585
R7843 GND.n2290 GND.n1254 585
R7844 GND.n2931 GND.n2290 585
R7845 GND.n2941 GND.n1253 585
R7846 GND.n2942 GND.n2941 585
R7847 GND.n2940 GND.n2300 585
R7848 GND.n2940 GND.n2939 585
R7849 GND.n2299 GND.n1247 585
R7850 GND.n2910 GND.n2299 585
R7851 GND.n2900 GND.n1246 585
R7852 GND.n2900 GND.n2316 585
R7853 GND.n2901 GND.n1245 585
R7854 GND.n2902 GND.n2901 585
R7855 GND.n2899 GND.n2326 585
R7856 GND.n2899 GND.n2898 585
R7857 GND.n2325 GND.n1239 585
R7858 GND.n2765 GND.n2325 585
R7859 GND.n2336 GND.n1238 585
R7860 GND.n2886 GND.n2336 585
R7861 GND.n2873 GND.n1237 585
R7862 GND.n2873 GND.n2872 585
R7863 GND.n2875 GND.n2874 585
R7864 GND.n2876 GND.n2875 585
R7865 GND.n2871 GND.n1231 585
R7866 GND.n2871 GND.n2870 585
R7867 GND.n2346 GND.n1230 585
R7868 GND.n2786 GND.n2346 585
R7869 GND.n2355 GND.n1229 585
R7870 GND.n2861 GND.n2355 585
R7871 GND.n2849 GND.n2847 585
R7872 GND.n2849 GND.n2848 585
R7873 GND.n2850 GND.n1223 585
R7874 GND.n2851 GND.n2850 585
R7875 GND.n2846 GND.n1222 585
R7876 GND.n2846 GND.n2845 585
R7877 GND.n2365 GND.n1221 585
R7878 GND.n2795 GND.n2365 585
R7879 GND.n2376 GND.n2375 585
R7880 GND.n2836 GND.n2376 585
R7881 GND.n2418 GND.n1215 585
R7882 GND.n2746 GND.n2418 585
R7883 GND.n2806 GND.n1214 585
R7884 GND.n2806 GND.n2805 585
R7885 GND.n2807 GND.n1213 585
R7886 GND.n2808 GND.n2807 585
R7887 GND.n2408 GND.n2407 585
R7888 GND.n2813 GND.n2408 585
R7889 GND.n2406 GND.n1207 585
R7890 GND.n2406 GND.n2403 585
R7891 GND.n2393 GND.n1206 585
R7892 GND.n2396 GND.n2393 585
R7893 GND.n2823 GND.n1205 585
R7894 GND.n2823 GND.n2822 585
R7895 GND.n2825 GND.n2824 585
R7896 GND.n2826 GND.n2825 585
R7897 GND.n2392 GND.n1199 585
R7898 GND.n2729 GND.n2392 585
R7899 GND.n2688 GND.n1198 585
R7900 GND.n2688 GND.n2427 585
R7901 GND.n2689 GND.n1197 585
R7902 GND.n2690 GND.n2689 585
R7903 GND.n2438 GND.n2437 585
R7904 GND.n2715 GND.n2438 585
R7905 GND.n2704 GND.n1191 585
R7906 GND.n2704 GND.n2435 585
R7907 GND.n2705 GND.n1190 585
R7908 GND.n2706 GND.n2705 585
R7909 GND.n2703 GND.n1189 585
R7910 GND.n2703 GND.n2702 585
R7911 GND.n2451 GND.n2450 585
R7912 GND.n2463 GND.n2451 585
R7913 GND.n2461 GND.n1183 585
R7914 GND.n2679 GND.n2461 585
R7915 GND.n2667 GND.n1182 585
R7916 GND.n2667 GND.n2666 585
R7917 GND.n2668 GND.n1181 585
R7918 GND.n2669 GND.n2668 585
R7919 GND.n2664 GND.n2473 585
R7920 GND.n2664 GND.n2663 585
R7921 GND.n2472 GND.n1175 585
R7922 GND.n2486 GND.n2472 585
R7923 GND.n2484 GND.n1174 585
R7924 GND.n2654 GND.n2484 585
R7925 GND.n2641 GND.n1173 585
R7926 GND.n2641 GND.n2640 585
R7927 GND.n2643 GND.n2642 585
R7928 GND.n2644 GND.n2643 585
R7929 GND.n2639 GND.n1167 585
R7930 GND.n2639 GND.n2638 585
R7931 GND.n2495 GND.n1166 585
R7932 GND.n2497 GND.n2495 585
R7933 GND.n2543 GND.n1165 585
R7934 GND.n2629 GND.n2543 585
R7935 GND.n2617 GND.n2616 585
R7936 GND.n2617 GND.n2504 585
R7937 GND.n2618 GND.n1159 585
R7938 GND.n2619 GND.n2618 585
R7939 GND.n2615 GND.n1158 585
R7940 GND.n2615 GND.n2552 585
R7941 GND.n2614 GND.n1157 585
R7942 GND.n2614 GND.n1111 585
R7943 GND.n2613 GND.n2612 585
R7944 GND.n2611 GND.n2555 585
R7945 GND.n2557 GND.n2556 585
R7946 GND.n2607 GND.n2559 585
R7947 GND.n2606 GND.n2560 585
R7948 GND.n2605 GND.n2561 585
R7949 GND.n2563 GND.n2562 585
R7950 GND.n2601 GND.n2565 585
R7951 GND.n2600 GND.n2566 585
R7952 GND.n2599 GND.n2567 585
R7953 GND.n2569 GND.n2568 585
R7954 GND.n2595 GND.n2571 585
R7955 GND.n2594 GND.n2572 585
R7956 GND.n2593 GND.n2573 585
R7957 GND.n2575 GND.n2574 585
R7958 GND.n2589 GND.n2586 585
R7959 GND.n2585 GND.n1110 585
R7960 GND.n4752 GND.n1110 585
R7961 GND.n4504 GND.n4503 585
R7962 GND.n4505 GND.n1374 585
R7963 GND.n1389 GND.n1366 585
R7964 GND.n4512 GND.n1365 585
R7965 GND.n4513 GND.n1364 585
R7966 GND.n1387 GND.n1356 585
R7967 GND.n4520 GND.n1355 585
R7968 GND.n4521 GND.n1354 585
R7969 GND.n1384 GND.n1348 585
R7970 GND.n4528 GND.n1347 585
R7971 GND.n4529 GND.n1346 585
R7972 GND.n1382 GND.n1345 585
R7973 GND.n1381 GND.n1380 585
R7974 GND.n1378 GND.n1319 585
R7975 GND.n4541 GND.n1318 585
R7976 GND.n4542 GND.n1317 585
R7977 GND.n4543 GND.n1316 585
R7978 GND.n4501 GND.n1316 585
R7979 GND.n2958 GND.n1262 585
R7980 GND.n4600 GND.n1262 585
R7981 GND.n2957 GND.n2956 585
R7982 GND.n2956 GND.n2955 585
R7983 GND.n2288 GND.n2287 585
R7984 GND.n2950 GND.n2288 585
R7985 GND.n2933 GND.n2932 585
R7986 GND.n2932 GND.n2931 585
R7987 GND.n2304 GND.n2297 585
R7988 GND.n2942 GND.n2297 585
R7989 GND.n2938 GND.n2937 585
R7990 GND.n2939 GND.n2938 585
R7991 GND.n2303 GND.n2302 585
R7992 GND.n2910 GND.n2302 585
R7993 GND.n2892 GND.n2891 585
R7994 GND.n2891 GND.n2316 585
R7995 GND.n2329 GND.n2323 585
R7996 GND.n2902 GND.n2323 585
R7997 GND.n2897 GND.n2896 585
R7998 GND.n2898 GND.n2897 585
R7999 GND.n2328 GND.n2327 585
R8000 GND.n2765 GND.n2327 585
R8001 GND.n2888 GND.n2887 585
R8002 GND.n2887 GND.n2886 585
R8003 GND.n2332 GND.n2331 585
R8004 GND.n2872 GND.n2332 585
R8005 GND.n2349 GND.n2344 585
R8006 GND.n2876 GND.n2344 585
R8007 GND.n2869 GND.n2868 585
R8008 GND.n2870 GND.n2869 585
R8009 GND.n2348 GND.n2347 585
R8010 GND.n2786 GND.n2347 585
R8011 GND.n2863 GND.n2862 585
R8012 GND.n2862 GND.n2861 585
R8013 GND.n2352 GND.n2351 585
R8014 GND.n2848 GND.n2352 585
R8015 GND.n2369 GND.n2363 585
R8016 GND.n2851 GND.n2363 585
R8017 GND.n2844 GND.n2843 585
R8018 GND.n2845 GND.n2844 585
R8019 GND.n2368 GND.n2367 585
R8020 GND.n2795 GND.n2367 585
R8021 GND.n2838 GND.n2837 585
R8022 GND.n2837 GND.n2836 585
R8023 GND.n2372 GND.n2371 585
R8024 GND.n2746 GND.n2372 585
R8025 GND.n2745 GND.n2744 585
R8026 GND.n2805 GND.n2745 585
R8027 GND.n2420 GND.n2416 585
R8028 GND.n2808 GND.n2416 585
R8029 GND.n2740 GND.n2404 585
R8030 GND.n2813 GND.n2404 585
R8031 GND.n2739 GND.n2738 585
R8032 GND.n2738 GND.n2403 585
R8033 GND.n2737 GND.n2736 585
R8034 GND.n2737 GND.n2396 585
R8035 GND.n2422 GND.n2394 585
R8036 GND.n2822 GND.n2394 585
R8037 GND.n2732 GND.n2390 585
R8038 GND.n2826 GND.n2390 585
R8039 GND.n2731 GND.n2730 585
R8040 GND.n2730 GND.n2729 585
R8041 GND.n2425 GND.n2424 585
R8042 GND.n2427 GND.n2425 585
R8043 GND.n2694 GND.n2691 585
R8044 GND.n2691 GND.n2690 585
R8045 GND.n2695 GND.n2436 585
R8046 GND.n2715 GND.n2436 585
R8047 GND.n2696 GND.n2685 585
R8048 GND.n2685 GND.n2435 585
R8049 GND.n2455 GND.n2448 585
R8050 GND.n2706 GND.n2448 585
R8051 GND.n2701 GND.n2700 585
R8052 GND.n2702 GND.n2701 585
R8053 GND.n2454 GND.n2453 585
R8054 GND.n2463 GND.n2453 585
R8055 GND.n2681 GND.n2680 585
R8056 GND.n2680 GND.n2679 585
R8057 GND.n2458 GND.n2457 585
R8058 GND.n2666 GND.n2458 585
R8059 GND.n2477 GND.n2470 585
R8060 GND.n2669 GND.n2470 585
R8061 GND.n2662 GND.n2661 585
R8062 GND.n2663 GND.n2662 585
R8063 GND.n2476 GND.n2475 585
R8064 GND.n2486 GND.n2475 585
R8065 GND.n2656 GND.n2655 585
R8066 GND.n2655 GND.n2654 585
R8067 GND.n2480 GND.n2479 585
R8068 GND.n2640 GND.n2480 585
R8069 GND.n2500 GND.n2493 585
R8070 GND.n2644 GND.n2493 585
R8071 GND.n2637 GND.n2636 585
R8072 GND.n2638 GND.n2637 585
R8073 GND.n2499 GND.n2498 585
R8074 GND.n2498 GND.n2497 585
R8075 GND.n2631 GND.n2630 585
R8076 GND.n2630 GND.n2629 585
R8077 GND.n2503 GND.n2502 585
R8078 GND.n2504 GND.n2503 585
R8079 GND.n2580 GND.n2553 585
R8080 GND.n2619 GND.n2553 585
R8081 GND.n2581 GND.n2578 585
R8082 GND.n2578 GND.n2552 585
R8083 GND.n2582 GND.n2577 585
R8084 GND.n2577 GND.n1111 585
R8085 GND.n4599 GND.n4598 585
R8086 GND.n4600 GND.n4599 585
R8087 GND.n1267 GND.n1265 585
R8088 GND.n2955 GND.n1265 585
R8089 GND.n2949 GND.n2948 585
R8090 GND.n2950 GND.n2949 585
R8091 GND.n2292 GND.n2291 585
R8092 GND.n2931 GND.n2291 585
R8093 GND.n2944 GND.n2943 585
R8094 GND.n2943 GND.n2942 585
R8095 GND.n2295 GND.n2294 585
R8096 GND.n2939 GND.n2295 585
R8097 GND.n2909 GND.n2908 585
R8098 GND.n2910 GND.n2909 585
R8099 GND.n2318 GND.n2317 585
R8100 GND.n2317 GND.n2316 585
R8101 GND.n2904 GND.n2903 585
R8102 GND.n2903 GND.n2902 585
R8103 GND.n2321 GND.n2320 585
R8104 GND.n2898 GND.n2321 585
R8105 GND.n2883 GND.n2338 585
R8106 GND.n2765 GND.n2338 585
R8107 GND.n2885 GND.n2884 585
R8108 GND.n2886 GND.n2885 585
R8109 GND.n2339 GND.n2337 585
R8110 GND.n2872 GND.n2337 585
R8111 GND.n2878 GND.n2877 585
R8112 GND.n2877 GND.n2876 585
R8113 GND.n2342 GND.n2341 585
R8114 GND.n2870 GND.n2342 585
R8115 GND.n2858 GND.n2357 585
R8116 GND.n2786 GND.n2357 585
R8117 GND.n2860 GND.n2859 585
R8118 GND.n2861 GND.n2860 585
R8119 GND.n2358 GND.n2356 585
R8120 GND.n2848 GND.n2356 585
R8121 GND.n2853 GND.n2852 585
R8122 GND.n2852 GND.n2851 585
R8123 GND.n2361 GND.n2360 585
R8124 GND.n2845 GND.n2361 585
R8125 GND.n2833 GND.n2378 585
R8126 GND.n2795 GND.n2378 585
R8127 GND.n2835 GND.n2834 585
R8128 GND.n2836 GND.n2835 585
R8129 GND.n2379 GND.n2377 585
R8130 GND.n2746 GND.n2377 585
R8131 GND.n2414 GND.n2413 585
R8132 GND.n2805 GND.n2413 585
R8133 GND.n2809 GND.n2415 585
R8134 GND.n2809 GND.n2808 585
R8135 GND.n2812 GND.n2811 585
R8136 GND.n2813 GND.n2812 585
R8137 GND.n2810 GND.n2412 585
R8138 GND.n2412 GND.n2403 585
R8139 GND.n2411 GND.n2410 585
R8140 GND.n2411 GND.n2396 585
R8141 GND.n2409 GND.n2388 585
R8142 GND.n2822 GND.n2388 585
R8143 GND.n2828 GND.n2827 585
R8144 GND.n2827 GND.n2826 585
R8145 GND.n2829 GND.n2387 585
R8146 GND.n2729 GND.n2387 585
R8147 GND.n2440 GND.n2386 585
R8148 GND.n2440 GND.n2427 585
R8149 GND.n2712 GND.n2441 585
R8150 GND.n2690 GND.n2441 585
R8151 GND.n2714 GND.n2713 585
R8152 GND.n2715 GND.n2714 585
R8153 GND.n2442 GND.n2439 585
R8154 GND.n2439 GND.n2435 585
R8155 GND.n2708 GND.n2707 585
R8156 GND.n2707 GND.n2706 585
R8157 GND.n2445 GND.n2444 585
R8158 GND.n2702 GND.n2445 585
R8159 GND.n2676 GND.n2464 585
R8160 GND.n2464 GND.n2463 585
R8161 GND.n2678 GND.n2677 585
R8162 GND.n2679 GND.n2678 585
R8163 GND.n2465 GND.n2462 585
R8164 GND.n2666 GND.n2462 585
R8165 GND.n2671 GND.n2670 585
R8166 GND.n2670 GND.n2669 585
R8167 GND.n2468 GND.n2467 585
R8168 GND.n2663 GND.n2468 585
R8169 GND.n2651 GND.n2487 585
R8170 GND.n2487 GND.n2486 585
R8171 GND.n2653 GND.n2652 585
R8172 GND.n2654 GND.n2653 585
R8173 GND.n2488 GND.n2485 585
R8174 GND.n2640 GND.n2485 585
R8175 GND.n2646 GND.n2645 585
R8176 GND.n2645 GND.n2644 585
R8177 GND.n2491 GND.n2490 585
R8178 GND.n2638 GND.n2491 585
R8179 GND.n2626 GND.n2545 585
R8180 GND.n2545 GND.n2497 585
R8181 GND.n2628 GND.n2627 585
R8182 GND.n2629 GND.n2628 585
R8183 GND.n2546 GND.n2544 585
R8184 GND.n2544 GND.n2504 585
R8185 GND.n2621 GND.n2620 585
R8186 GND.n2620 GND.n2619 585
R8187 GND.n2551 GND.n2550 585
R8188 GND.n2552 GND.n2551 585
R8189 GND.n2549 GND.n1114 585
R8190 GND.n1114 GND.n1111 585
R8191 GND.n4750 GND.n4749 585
R8192 GND.n4748 GND.n1113 585
R8193 GND.n4747 GND.n1112 585
R8194 GND.n4752 GND.n1112 585
R8195 GND.n4746 GND.n4745 585
R8196 GND.n4744 GND.n4743 585
R8197 GND.n4742 GND.n4741 585
R8198 GND.n4740 GND.n4739 585
R8199 GND.n4738 GND.n4737 585
R8200 GND.n4736 GND.n4735 585
R8201 GND.n4734 GND.n4733 585
R8202 GND.n4732 GND.n4731 585
R8203 GND.n4730 GND.n4729 585
R8204 GND.n4728 GND.n4727 585
R8205 GND.n4726 GND.n4725 585
R8206 GND.n4724 GND.n4723 585
R8207 GND.n4722 GND.n4721 585
R8208 GND.n4719 GND.n4718 585
R8209 GND.n4717 GND.n4716 585
R8210 GND.n4715 GND.n4714 585
R8211 GND.n4713 GND.n4712 585
R8212 GND.n4711 GND.n4710 585
R8213 GND.n4709 GND.n4708 585
R8214 GND.n4707 GND.n4706 585
R8215 GND.n4705 GND.n4704 585
R8216 GND.n4703 GND.n4702 585
R8217 GND.n4701 GND.n4700 585
R8218 GND.n4699 GND.n4698 585
R8219 GND.n4697 GND.n4696 585
R8220 GND.n4695 GND.n4694 585
R8221 GND.n4693 GND.n4692 585
R8222 GND.n4691 GND.n4690 585
R8223 GND.n4689 GND.n4688 585
R8224 GND.n4687 GND.n1149 585
R8225 GND.n1153 GND.n1150 585
R8226 GND.n4683 GND.n4682 585
R8227 GND.n4546 GND.n1260 585
R8228 GND.n4476 GND.n1314 585
R8229 GND.n4550 GND.n1311 585
R8230 GND.n4551 GND.n1310 585
R8231 GND.n4552 GND.n1309 585
R8232 GND.n4479 GND.n1307 585
R8233 GND.n4556 GND.n1306 585
R8234 GND.n4557 GND.n1305 585
R8235 GND.n4558 GND.n1304 585
R8236 GND.n4482 GND.n1302 585
R8237 GND.n4562 GND.n1301 585
R8238 GND.n4563 GND.n1300 585
R8239 GND.n4564 GND.n1299 585
R8240 GND.n4485 GND.n1297 585
R8241 GND.n4568 GND.n1296 585
R8242 GND.n4569 GND.n1295 585
R8243 GND.n4570 GND.n1294 585
R8244 GND.n4488 GND.n1292 585
R8245 GND.n4574 GND.n1291 585
R8246 GND.n4576 GND.n1285 585
R8247 GND.n4577 GND.n1284 585
R8248 GND.n4492 GND.n1282 585
R8249 GND.n4581 GND.n1281 585
R8250 GND.n4582 GND.n1280 585
R8251 GND.n4583 GND.n1279 585
R8252 GND.n4495 GND.n1277 585
R8253 GND.n4587 GND.n1276 585
R8254 GND.n4588 GND.n1275 585
R8255 GND.n4589 GND.n1274 585
R8256 GND.n4498 GND.n1272 585
R8257 GND.n4593 GND.n1271 585
R8258 GND.n4594 GND.n1270 585
R8259 GND.n4595 GND.n1266 585
R8260 GND.n4501 GND.n1266 585
R8261 GND.n4602 GND.n4601 585
R8262 GND.n4601 GND.n4600 585
R8263 GND.n4603 GND.n1258 585
R8264 GND.n2955 GND.n1258 585
R8265 GND.n4604 GND.n1257 585
R8266 GND.n2950 GND.n1257 585
R8267 GND.n2307 GND.n1252 585
R8268 GND.n2931 GND.n2307 585
R8269 GND.n4608 GND.n1251 585
R8270 GND.n2942 GND.n1251 585
R8271 GND.n4609 GND.n1250 585
R8272 GND.n2939 GND.n1250 585
R8273 GND.n4610 GND.n1249 585
R8274 GND.n2910 GND.n1249 585
R8275 GND.n2315 GND.n1244 585
R8276 GND.n2316 GND.n2315 585
R8277 GND.n4614 GND.n1243 585
R8278 GND.n2902 GND.n1243 585
R8279 GND.n4615 GND.n1242 585
R8280 GND.n2898 GND.n1242 585
R8281 GND.n4616 GND.n1241 585
R8282 GND.n2765 GND.n1241 585
R8283 GND.n2334 GND.n1236 585
R8284 GND.n2886 GND.n2334 585
R8285 GND.n4620 GND.n1235 585
R8286 GND.n2872 GND.n1235 585
R8287 GND.n4621 GND.n1234 585
R8288 GND.n2876 GND.n1234 585
R8289 GND.n4622 GND.n1233 585
R8290 GND.n2870 GND.n1233 585
R8291 GND.n2785 GND.n1228 585
R8292 GND.n2786 GND.n2785 585
R8293 GND.n4626 GND.n1227 585
R8294 GND.n2861 GND.n1227 585
R8295 GND.n4627 GND.n1226 585
R8296 GND.n2848 GND.n1226 585
R8297 GND.n4628 GND.n1225 585
R8298 GND.n2851 GND.n1225 585
R8299 GND.n2366 GND.n1220 585
R8300 GND.n2845 GND.n2366 585
R8301 GND.n4632 GND.n1219 585
R8302 GND.n2795 GND.n1219 585
R8303 GND.n4633 GND.n1218 585
R8304 GND.n2836 GND.n1218 585
R8305 GND.n4634 GND.n1217 585
R8306 GND.n2746 GND.n1217 585
R8307 GND.n2419 GND.n1212 585
R8308 GND.n2805 GND.n2419 585
R8309 GND.n4638 GND.n1211 585
R8310 GND.n2808 GND.n1211 585
R8311 GND.n4639 GND.n1210 585
R8312 GND.n2813 GND.n1210 585
R8313 GND.n4640 GND.n1209 585
R8314 GND.n2403 GND.n1209 585
R8315 GND.n2395 GND.n1204 585
R8316 GND.n2396 GND.n2395 585
R8317 GND.n4644 GND.n1203 585
R8318 GND.n2822 GND.n1203 585
R8319 GND.n4645 GND.n1202 585
R8320 GND.n2826 GND.n1202 585
R8321 GND.n4646 GND.n1201 585
R8322 GND.n2729 GND.n1201 585
R8323 GND.n2426 GND.n1196 585
R8324 GND.n2427 GND.n2426 585
R8325 GND.n4650 GND.n1195 585
R8326 GND.n2690 GND.n1195 585
R8327 GND.n4651 GND.n1194 585
R8328 GND.n2715 GND.n1194 585
R8329 GND.n4652 GND.n1193 585
R8330 GND.n2435 GND.n1193 585
R8331 GND.n2447 GND.n1188 585
R8332 GND.n2706 GND.n2447 585
R8333 GND.n4656 GND.n1187 585
R8334 GND.n2702 GND.n1187 585
R8335 GND.n4657 GND.n1186 585
R8336 GND.n2463 GND.n1186 585
R8337 GND.n4658 GND.n1185 585
R8338 GND.n2679 GND.n1185 585
R8339 GND.n2665 GND.n1180 585
R8340 GND.n2666 GND.n2665 585
R8341 GND.n4662 GND.n1179 585
R8342 GND.n2669 GND.n1179 585
R8343 GND.n4663 GND.n1178 585
R8344 GND.n2663 GND.n1178 585
R8345 GND.n4664 GND.n1177 585
R8346 GND.n2486 GND.n1177 585
R8347 GND.n2482 GND.n1172 585
R8348 GND.n2654 GND.n2482 585
R8349 GND.n4668 GND.n1171 585
R8350 GND.n2640 GND.n1171 585
R8351 GND.n4669 GND.n1170 585
R8352 GND.n2644 GND.n1170 585
R8353 GND.n4670 GND.n1169 585
R8354 GND.n2638 GND.n1169 585
R8355 GND.n2496 GND.n1164 585
R8356 GND.n2497 GND.n2496 585
R8357 GND.n4674 GND.n1163 585
R8358 GND.n2629 GND.n1163 585
R8359 GND.n4675 GND.n1162 585
R8360 GND.n2504 GND.n1162 585
R8361 GND.n4676 GND.n1161 585
R8362 GND.n2619 GND.n1161 585
R8363 GND.n1156 GND.n1155 585
R8364 GND.n2552 GND.n1155 585
R8365 GND.n4681 GND.n4680 585
R8366 GND.n4681 GND.n1111 585
R8367 GND.n5519 GND.n494 585
R8368 GND.n494 GND.n467 585
R8369 GND.n5521 GND.n5520 585
R8370 GND.n5522 GND.n5521 585
R8371 GND.n558 GND.n557 585
R8372 GND.n557 GND.n556 585
R8373 GND.n5515 GND.n5514 585
R8374 GND.n5514 GND.n5513 585
R8375 GND.n561 GND.n560 585
R8376 GND.n562 GND.n561 585
R8377 GND.n5502 GND.n5501 585
R8378 GND.n5503 GND.n5502 585
R8379 GND.n576 GND.n575 585
R8380 GND.n575 GND.n572 585
R8381 GND.n5497 GND.n5496 585
R8382 GND.n5496 GND.n5495 585
R8383 GND.n579 GND.n578 585
R8384 GND.n5487 GND.n579 585
R8385 GND.n4127 GND.n1946 585
R8386 GND.n1946 GND.n594 585
R8387 GND.n4129 GND.n4128 585
R8388 GND.n4130 GND.n4129 585
R8389 GND.n1947 GND.n1945 585
R8390 GND.n1953 GND.n1945 585
R8391 GND.n4122 GND.n4121 585
R8392 GND.n4121 GND.n4120 585
R8393 GND.n1950 GND.n1949 585
R8394 GND.n4117 GND.n1950 585
R8395 GND.n4094 GND.n1969 585
R8396 GND.n1969 GND.n1956 585
R8397 GND.n4096 GND.n4095 585
R8398 GND.n4097 GND.n4096 585
R8399 GND.n1970 GND.n1968 585
R8400 GND.n1968 GND.n1963 585
R8401 GND.n4089 GND.n4088 585
R8402 GND.n4088 GND.n4087 585
R8403 GND.n1973 GND.n1972 585
R8404 GND.n4083 GND.n1973 585
R8405 GND.n4068 GND.n1992 585
R8406 GND.n1992 GND.n1980 585
R8407 GND.n4070 GND.n4069 585
R8408 GND.n4071 GND.n4070 585
R8409 GND.n1993 GND.n1991 585
R8410 GND.n1991 GND.n1988 585
R8411 GND.n4031 GND.n4030 585
R8412 GND.n4032 GND.n4031 585
R8413 GND.n4022 GND.n4021 585
R8414 GND.n4040 GND.n4021 585
R8415 GND.n4044 GND.n4023 585
R8416 GND.n4044 GND.n4043 585
R8417 GND.n4047 GND.n4046 585
R8418 GND.n4048 GND.n4047 585
R8419 GND.n4045 GND.n4020 585
R8420 GND.n4020 GND.n4012 585
R8421 GND.n4019 GND.n4018 585
R8422 GND.n4019 GND.n2011 585
R8423 GND.n4017 GND.n2001 585
R8424 GND.n4057 GND.n2001 585
R8425 GND.n4062 GND.n4061 585
R8426 GND.n4061 GND.n4060 585
R8427 GND.n4063 GND.n2000 585
R8428 GND.n4002 GND.n2000 585
R8429 GND.n2030 GND.n1999 585
R8430 GND.n2030 GND.n2017 585
R8431 GND.n3990 GND.n3989 585
R8432 GND.n3991 GND.n3990 585
R8433 GND.n3988 GND.n2029 585
R8434 GND.n2043 GND.n2029 585
R8435 GND.n2035 GND.n2031 585
R8436 GND.n3978 GND.n2035 585
R8437 GND.n3984 GND.n3983 585
R8438 GND.n3983 GND.n3982 585
R8439 GND.n2034 GND.n2033 585
R8440 GND.n3963 GND.n2034 585
R8441 GND.n3949 GND.n2063 585
R8442 GND.n2063 GND.n2051 585
R8443 GND.n3951 GND.n3950 585
R8444 GND.n3952 GND.n3951 585
R8445 GND.n2064 GND.n2062 585
R8446 GND.n3939 GND.n2062 585
R8447 GND.n3944 GND.n3943 585
R8448 GND.n3943 GND.n3942 585
R8449 GND.n2067 GND.n2066 585
R8450 GND.n3936 GND.n2067 585
R8451 GND.n3924 GND.n2084 585
R8452 GND.n3874 GND.n2084 585
R8453 GND.n3926 GND.n3925 585
R8454 GND.n3927 GND.n3926 585
R8455 GND.n2085 GND.n2083 585
R8456 GND.n3914 GND.n2083 585
R8457 GND.n3919 GND.n3918 585
R8458 GND.n3918 GND.n3917 585
R8459 GND.n2088 GND.n2087 585
R8460 GND.n3912 GND.n2088 585
R8461 GND.n3900 GND.n2107 585
R8462 GND.n2107 GND.n2106 585
R8463 GND.n3902 GND.n3901 585
R8464 GND.n3903 GND.n3902 585
R8465 GND.n2108 GND.n2105 585
R8466 GND.n3890 GND.n2105 585
R8467 GND.n3895 GND.n3894 585
R8468 GND.n3894 GND.n3893 585
R8469 GND.n2111 GND.n2110 585
R8470 GND.n3843 GND.n2111 585
R8471 GND.n3589 GND.n3588 585
R8472 GND.n3589 GND.n2137 585
R8473 GND.n3591 GND.n3590 585
R8474 GND.n3595 GND.n3586 585
R8475 GND.n3597 GND.n3596 585
R8476 GND.n3599 GND.n3598 585
R8477 GND.n3601 GND.n3600 585
R8478 GND.n3605 GND.n3584 585
R8479 GND.n3607 GND.n3606 585
R8480 GND.n3609 GND.n3608 585
R8481 GND.n3611 GND.n3610 585
R8482 GND.n3615 GND.n3582 585
R8483 GND.n3617 GND.n3616 585
R8484 GND.n3619 GND.n3618 585
R8485 GND.n3621 GND.n3620 585
R8486 GND.n3579 GND.n3578 585
R8487 GND.n4214 GND.n1830 585
R8488 GND.n3684 GND.n3683 585
R8489 GND.n3682 GND.n3681 585
R8490 GND.n3680 GND.n3679 585
R8491 GND.n3678 GND.n3677 585
R8492 GND.n3676 GND.n3675 585
R8493 GND.n3674 GND.n3673 585
R8494 GND.n3672 GND.n3671 585
R8495 GND.n3670 GND.n3669 585
R8496 GND.n3668 GND.n3667 585
R8497 GND.n3666 GND.n3665 585
R8498 GND.n3664 GND.n3663 585
R8499 GND.n3662 GND.n3661 585
R8500 GND.n3660 GND.n3659 585
R8501 GND.n3658 GND.n3657 585
R8502 GND.n3656 GND.n3655 585
R8503 GND.n3654 GND.n3653 585
R8504 GND.n3652 GND.n3643 585
R8505 GND.n3649 GND.n3646 585
R8506 GND.n3645 GND.n3644 585
R8507 GND.n5575 GND.n5574 585
R8508 GND.n549 GND.n548 585
R8509 GND.n5579 GND.n545 585
R8510 GND.n5580 GND.n544 585
R8511 GND.n5581 GND.n543 585
R8512 GND.n541 GND.n540 585
R8513 GND.n5585 GND.n539 585
R8514 GND.n5586 GND.n538 585
R8515 GND.n5587 GND.n537 585
R8516 GND.n535 GND.n534 585
R8517 GND.n5591 GND.n533 585
R8518 GND.n5592 GND.n532 585
R8519 GND.n5593 GND.n531 585
R8520 GND.n529 GND.n528 585
R8521 GND.n5597 GND.n527 585
R8522 GND.n5598 GND.n526 585
R8523 GND.n5599 GND.n525 585
R8524 GND.n523 GND.n522 585
R8525 GND.n5603 GND.n521 585
R8526 GND.n5605 GND.n518 585
R8527 GND.n5606 GND.n517 585
R8528 GND.n515 GND.n514 585
R8529 GND.n5610 GND.n513 585
R8530 GND.n5611 GND.n512 585
R8531 GND.n5612 GND.n511 585
R8532 GND.n509 GND.n508 585
R8533 GND.n5616 GND.n507 585
R8534 GND.n5617 GND.n506 585
R8535 GND.n5618 GND.n505 585
R8536 GND.n503 GND.n502 585
R8537 GND.n5622 GND.n501 585
R8538 GND.n5623 GND.n500 585
R8539 GND.n5624 GND.n499 585
R8540 GND.n496 GND.n495 585
R8541 GND.n5629 GND.n5628 585
R8542 GND.n5630 GND.n5629 585
R8543 GND.n5573 GND.n5572 585
R8544 GND.n5573 GND.n467 585
R8545 GND.n552 GND.n551 585
R8546 GND.n5522 GND.n551 585
R8547 GND.n5508 GND.n5507 585
R8548 GND.n5507 GND.n556 585
R8549 GND.n5509 GND.n563 585
R8550 GND.n5513 GND.n563 585
R8551 GND.n5506 GND.n5505 585
R8552 GND.n5505 GND.n562 585
R8553 GND.n5504 GND.n570 585
R8554 GND.n5504 GND.n5503 585
R8555 GND.n5490 GND.n571 585
R8556 GND.n572 GND.n571 585
R8557 GND.n5491 GND.n581 585
R8558 GND.n5495 GND.n581 585
R8559 GND.n5489 GND.n5488 585
R8560 GND.n5488 GND.n5487 585
R8561 GND.n593 GND.n592 585
R8562 GND.n594 GND.n593 585
R8563 GND.n4136 GND.n1939 585
R8564 GND.n4130 GND.n1939 585
R8565 GND.n4137 GND.n1938 585
R8566 GND.n1953 GND.n1938 585
R8567 GND.n4138 GND.n1937 585
R8568 GND.n4120 GND.n1937 585
R8569 GND.n4116 GND.n1932 585
R8570 GND.n4117 GND.n4116 585
R8571 GND.n4142 GND.n1931 585
R8572 GND.n1956 GND.n1931 585
R8573 GND.n4143 GND.n1930 585
R8574 GND.n4097 GND.n1930 585
R8575 GND.n4144 GND.n1929 585
R8576 GND.n1963 GND.n1929 585
R8577 GND.n1975 GND.n1924 585
R8578 GND.n4087 GND.n1975 585
R8579 GND.n4148 GND.n1923 585
R8580 GND.n4083 GND.n1923 585
R8581 GND.n4149 GND.n1922 585
R8582 GND.n1980 GND.n1922 585
R8583 GND.n4150 GND.n1921 585
R8584 GND.n4071 GND.n1921 585
R8585 GND.n1987 GND.n1916 585
R8586 GND.n1988 GND.n1987 585
R8587 GND.n4154 GND.n1915 585
R8588 GND.n4032 GND.n1915 585
R8589 GND.n4155 GND.n1914 585
R8590 GND.n4040 GND.n1914 585
R8591 GND.n4156 GND.n1913 585
R8592 GND.n4043 GND.n1913 585
R8593 GND.n4013 GND.n1908 585
R8594 GND.n4048 GND.n4013 585
R8595 GND.n4160 GND.n1907 585
R8596 GND.n4012 GND.n1907 585
R8597 GND.n4161 GND.n1906 585
R8598 GND.n2011 GND.n1906 585
R8599 GND.n4162 GND.n1905 585
R8600 GND.n4057 GND.n1905 585
R8601 GND.n2003 GND.n1900 585
R8602 GND.n4060 GND.n2003 585
R8603 GND.n4166 GND.n1899 585
R8604 GND.n4002 GND.n1899 585
R8605 GND.n4167 GND.n1898 585
R8606 GND.n2017 GND.n1898 585
R8607 GND.n4168 GND.n1897 585
R8608 GND.n3991 GND.n1897 585
R8609 GND.n2042 GND.n1892 585
R8610 GND.n2043 GND.n2042 585
R8611 GND.n4172 GND.n1891 585
R8612 GND.n3978 GND.n1891 585
R8613 GND.n4173 GND.n1890 585
R8614 GND.n3982 GND.n1890 585
R8615 GND.n4174 GND.n1889 585
R8616 GND.n3963 GND.n1889 585
R8617 GND.n2050 GND.n1884 585
R8618 GND.n2051 GND.n2050 585
R8619 GND.n4178 GND.n1883 585
R8620 GND.n3952 GND.n1883 585
R8621 GND.n4179 GND.n1882 585
R8622 GND.n3939 GND.n1882 585
R8623 GND.n4180 GND.n1881 585
R8624 GND.n3942 GND.n1881 585
R8625 GND.n2073 GND.n1876 585
R8626 GND.n3936 GND.n2073 585
R8627 GND.n4184 GND.n1875 585
R8628 GND.n3874 GND.n1875 585
R8629 GND.n4185 GND.n1874 585
R8630 GND.n3927 GND.n1874 585
R8631 GND.n4186 GND.n1873 585
R8632 GND.n3914 GND.n1873 585
R8633 GND.n2090 GND.n1868 585
R8634 GND.n3917 GND.n2090 585
R8635 GND.n4190 GND.n1867 585
R8636 GND.n3912 GND.n1867 585
R8637 GND.n4191 GND.n1866 585
R8638 GND.n2106 GND.n1866 585
R8639 GND.n4192 GND.n1865 585
R8640 GND.n3903 GND.n1865 585
R8641 GND.n3889 GND.n1860 585
R8642 GND.n3890 GND.n3889 585
R8643 GND.n4196 GND.n1859 585
R8644 GND.n3893 GND.n1859 585
R8645 GND.n4197 GND.n1858 585
R8646 GND.n3843 GND.n1858 585
R8647 GND.n4198 GND.n1857 585
R8648 GND.n2137 GND.n1857 585
R8649 GND.n1685 GND.n1684 585
R8650 GND.n3773 GND.n1685 585
R8651 GND.n4300 GND.n4299 585
R8652 GND.n4299 GND.n4298 585
R8653 GND.n4301 GND.n1682 585
R8654 GND.n3779 GND.n1682 585
R8655 GND.n4303 GND.n4302 585
R8656 GND.n4304 GND.n4303 585
R8657 GND.n1683 GND.n1681 585
R8658 GND.n3451 GND.n1681 585
R8659 GND.n3434 GND.n3433 585
R8660 GND.n3434 GND.n2181 585
R8661 GND.n3436 GND.n3435 585
R8662 GND.n3435 GND.n1664 585
R8663 GND.n3437 GND.n3432 585
R8664 GND.n3432 GND.n1662 585
R8665 GND.n3439 GND.n3438 585
R8666 GND.n3440 GND.n3439 585
R8667 GND.n1650 GND.n1649 585
R8668 GND.n2187 GND.n1650 585
R8669 GND.n4321 GND.n4320 585
R8670 GND.n4320 GND.n4319 585
R8671 GND.n4322 GND.n1647 585
R8672 GND.n3422 GND.n1647 585
R8673 GND.n4324 GND.n4323 585
R8674 GND.n4325 GND.n4324 585
R8675 GND.n1648 GND.n1646 585
R8676 GND.n3418 GND.n1646 585
R8677 GND.n1625 GND.n1624 585
R8678 GND.n2192 GND.n1625 585
R8679 GND.n4334 GND.n4333 585
R8680 GND.n4333 GND.n4332 585
R8681 GND.n4335 GND.n1622 585
R8682 GND.n3372 GND.n1622 585
R8683 GND.n4337 GND.n4336 585
R8684 GND.n4338 GND.n4337 585
R8685 GND.n1623 GND.n1621 585
R8686 GND.n3376 GND.n1621 585
R8687 GND.n3392 GND.n3391 585
R8688 GND.n3393 GND.n3392 585
R8689 GND.n3390 GND.n2201 585
R8690 GND.n2201 GND.n2198 585
R8691 GND.n3389 GND.n3388 585
R8692 GND.n3388 GND.n1603 585
R8693 GND.n3387 GND.n2202 585
R8694 GND.n3387 GND.n3386 585
R8695 GND.n1582 GND.n1581 585
R8696 GND.n2204 GND.n1582 585
R8697 GND.n4355 GND.n4354 585
R8698 GND.n4354 GND.n4353 585
R8699 GND.n4356 GND.n1579 585
R8700 GND.n3366 GND.n1579 585
R8701 GND.n4358 GND.n4357 585
R8702 GND.n4359 GND.n4358 585
R8703 GND.n1580 GND.n1578 585
R8704 GND.n3362 GND.n1578 585
R8705 GND.n1558 GND.n1557 585
R8706 GND.n3360 GND.n1558 585
R8707 GND.n4369 GND.n4368 585
R8708 GND.n4368 GND.n4367 585
R8709 GND.n4370 GND.n1555 585
R8710 GND.n3354 GND.n1555 585
R8711 GND.n4372 GND.n4371 585
R8712 GND.n4373 GND.n4372 585
R8713 GND.n1556 GND.n1554 585
R8714 GND.n3350 GND.n1554 585
R8715 GND.n3315 GND.n3314 585
R8716 GND.n3314 GND.n2210 585
R8717 GND.n3316 GND.n3312 585
R8718 GND.n3312 GND.n1541 585
R8719 GND.n3318 GND.n3317 585
R8720 GND.n3319 GND.n3318 585
R8721 GND.n3313 GND.n3311 585
R8722 GND.n3311 GND.n2216 585
R8723 GND.n1529 GND.n1528 585
R8724 GND.n3304 GND.n1529 585
R8725 GND.n4390 GND.n4389 585
R8726 GND.n4389 GND.n4388 585
R8727 GND.n4391 GND.n1526 585
R8728 GND.n3299 GND.n1526 585
R8729 GND.n4393 GND.n4392 585
R8730 GND.n4394 GND.n4393 585
R8731 GND.n1527 GND.n1525 585
R8732 GND.n1525 GND.n1520 585
R8733 GND.n3293 GND.n3292 585
R8734 GND.n3294 GND.n3293 585
R8735 GND.n1509 GND.n1508 585
R8736 GND.n1512 GND.n1509 585
R8737 GND.n4404 GND.n4403 585
R8738 GND.n4403 GND.n4402 585
R8739 GND.n4405 GND.n1506 585
R8740 GND.n3139 GND.n1506 585
R8741 GND.n4407 GND.n4406 585
R8742 GND.n4408 GND.n4407 585
R8743 GND.n1507 GND.n1505 585
R8744 GND.n1505 GND.n1502 585
R8745 GND.n2229 GND.n2228 585
R8746 GND.n2230 GND.n2229 585
R8747 GND.n1491 GND.n1490 585
R8748 GND.n1494 GND.n1491 585
R8749 GND.n4418 GND.n4417 585
R8750 GND.n4417 GND.n4416 585
R8751 GND.n4419 GND.n1488 585
R8752 GND.n3149 GND.n1488 585
R8753 GND.n4421 GND.n4420 585
R8754 GND.n4422 GND.n4421 585
R8755 GND.n1489 GND.n1487 585
R8756 GND.n1487 GND.n1485 585
R8757 GND.n3230 GND.n3229 585
R8758 GND.n3231 GND.n3230 585
R8759 GND.n3228 GND.n2243 585
R8760 GND.n2243 GND.n1474 585
R8761 GND.n3226 GND.n3225 585
R8762 GND.n2265 GND.n2264 585
R8763 GND.n3222 GND.n3221 585
R8764 GND.n3223 GND.n3222 585
R8765 GND.n3220 GND.n3160 585
R8766 GND.n3219 GND.n3218 585
R8767 GND.n3217 GND.n3216 585
R8768 GND.n3215 GND.n3214 585
R8769 GND.n3213 GND.n3212 585
R8770 GND.n3211 GND.n3210 585
R8771 GND.n3209 GND.n3208 585
R8772 GND.n3207 GND.n3206 585
R8773 GND.n3205 GND.n3204 585
R8774 GND.n3203 GND.n3202 585
R8775 GND.n3201 GND.n3200 585
R8776 GND.n3199 GND.n3198 585
R8777 GND.n3197 GND.n3196 585
R8778 GND.n3195 GND.n3194 585
R8779 GND.n3193 GND.n3192 585
R8780 GND.n3191 GND.n3190 585
R8781 GND.n3189 GND.n3188 585
R8782 GND.n3187 GND.n3186 585
R8783 GND.n3185 GND.n3184 585
R8784 GND.n3183 GND.n3182 585
R8785 GND.n3181 GND.n3180 585
R8786 GND.n3179 GND.n3178 585
R8787 GND.n3177 GND.n3176 585
R8788 GND.n3175 GND.n3174 585
R8789 GND.n3173 GND.n3172 585
R8790 GND.n3171 GND.n3170 585
R8791 GND.n3169 GND.n3168 585
R8792 GND.n3167 GND.n3166 585
R8793 GND.n3165 GND.n3164 585
R8794 GND.n3072 GND.n1290 585
R8795 GND.n3074 GND.n3073 585
R8796 GND.n3076 GND.n3075 585
R8797 GND.n3078 GND.n3077 585
R8798 GND.n3081 GND.n3080 585
R8799 GND.n3083 GND.n3082 585
R8800 GND.n3085 GND.n3084 585
R8801 GND.n3087 GND.n3086 585
R8802 GND.n3089 GND.n3088 585
R8803 GND.n3091 GND.n3090 585
R8804 GND.n3093 GND.n3092 585
R8805 GND.n3095 GND.n3094 585
R8806 GND.n3097 GND.n3096 585
R8807 GND.n3099 GND.n3098 585
R8808 GND.n3101 GND.n3100 585
R8809 GND.n3103 GND.n3102 585
R8810 GND.n3105 GND.n3104 585
R8811 GND.n3107 GND.n3106 585
R8812 GND.n3109 GND.n3108 585
R8813 GND.n3111 GND.n3110 585
R8814 GND.n3113 GND.n3112 585
R8815 GND.n3115 GND.n3114 585
R8816 GND.n3117 GND.n3116 585
R8817 GND.n3119 GND.n3118 585
R8818 GND.n3121 GND.n3120 585
R8819 GND.n3123 GND.n3122 585
R8820 GND.n3125 GND.n3124 585
R8821 GND.n3127 GND.n3126 585
R8822 GND.n3129 GND.n3128 585
R8823 GND.n3131 GND.n3130 585
R8824 GND.n3133 GND.n3132 585
R8825 GND.n3134 GND.n3068 585
R8826 GND.n3158 GND.n3157 585
R8827 GND.n3456 GND.n3455 585
R8828 GND.n3692 GND.n3691 585
R8829 GND.n3694 GND.n3693 585
R8830 GND.n3696 GND.n3695 585
R8831 GND.n3698 GND.n3697 585
R8832 GND.n3700 GND.n3699 585
R8833 GND.n3702 GND.n3701 585
R8834 GND.n3704 GND.n3703 585
R8835 GND.n3706 GND.n3705 585
R8836 GND.n3708 GND.n3707 585
R8837 GND.n3710 GND.n3709 585
R8838 GND.n3712 GND.n3711 585
R8839 GND.n3714 GND.n3713 585
R8840 GND.n3716 GND.n3715 585
R8841 GND.n3718 GND.n3717 585
R8842 GND.n3720 GND.n3719 585
R8843 GND.n3722 GND.n3721 585
R8844 GND.n3724 GND.n3723 585
R8845 GND.n3726 GND.n3725 585
R8846 GND.n3728 GND.n3727 585
R8847 GND.n3730 GND.n3729 585
R8848 GND.n3732 GND.n3731 585
R8849 GND.n3734 GND.n3733 585
R8850 GND.n3736 GND.n3735 585
R8851 GND.n3738 GND.n3737 585
R8852 GND.n3740 GND.n3739 585
R8853 GND.n3742 GND.n3741 585
R8854 GND.n3744 GND.n3743 585
R8855 GND.n3746 GND.n3745 585
R8856 GND.n3749 GND.n3748 585
R8857 GND.n3751 GND.n3750 585
R8858 GND.n3753 GND.n3752 585
R8859 GND.n3755 GND.n3754 585
R8860 GND.n3688 GND.n3687 585
R8861 GND.n3686 GND.n3577 585
R8862 GND.n3576 GND.n3575 585
R8863 GND.n3574 GND.n3573 585
R8864 GND.n3571 GND.n3570 585
R8865 GND.n3569 GND.n3568 585
R8866 GND.n3567 GND.n3566 585
R8867 GND.n3565 GND.n3564 585
R8868 GND.n3563 GND.n3562 585
R8869 GND.n3561 GND.n3560 585
R8870 GND.n3559 GND.n3558 585
R8871 GND.n3557 GND.n3556 585
R8872 GND.n3555 GND.n3554 585
R8873 GND.n3553 GND.n3552 585
R8874 GND.n3551 GND.n3550 585
R8875 GND.n3549 GND.n3548 585
R8876 GND.n3547 GND.n3546 585
R8877 GND.n3545 GND.n3544 585
R8878 GND.n3543 GND.n3542 585
R8879 GND.n3541 GND.n3540 585
R8880 GND.n3539 GND.n3538 585
R8881 GND.n3537 GND.n3536 585
R8882 GND.n3535 GND.n3534 585
R8883 GND.n3533 GND.n3532 585
R8884 GND.n3531 GND.n3530 585
R8885 GND.n3529 GND.n3528 585
R8886 GND.n3527 GND.n3526 585
R8887 GND.n3525 GND.n3524 585
R8888 GND.n3523 GND.n3522 585
R8889 GND.n3521 GND.n3520 585
R8890 GND.n3519 GND.n3518 585
R8891 GND.n3517 GND.n3516 585
R8892 GND.n3515 GND.n3514 585
R8893 GND.n3775 GND.n3774 585
R8894 GND.n3774 GND.n3773 585
R8895 GND.n3776 GND.n1687 585
R8896 GND.n4298 GND.n1687 585
R8897 GND.n3778 GND.n3777 585
R8898 GND.n3779 GND.n3778 585
R8899 GND.n3454 GND.n1680 585
R8900 GND.n4304 GND.n1680 585
R8901 GND.n3453 GND.n3452 585
R8902 GND.n3452 GND.n3451 585
R8903 GND.n2179 GND.n2178 585
R8904 GND.n2181 GND.n2179 585
R8905 GND.n3428 GND.n3427 585
R8906 GND.n3427 GND.n1664 585
R8907 GND.n3429 GND.n2189 585
R8908 GND.n2189 GND.n1662 585
R8909 GND.n3431 GND.n3430 585
R8910 GND.n3440 GND.n3431 585
R8911 GND.n3426 GND.n2188 585
R8912 GND.n2188 GND.n2187 585
R8913 GND.n3425 GND.n1652 585
R8914 GND.n4319 GND.n1652 585
R8915 GND.n3424 GND.n3423 585
R8916 GND.n3423 GND.n3422 585
R8917 GND.n3421 GND.n1644 585
R8918 GND.n4325 GND.n1644 585
R8919 GND.n3420 GND.n3419 585
R8920 GND.n3419 GND.n3418 585
R8921 GND.n2191 GND.n2190 585
R8922 GND.n2192 GND.n2191 585
R8923 GND.n3371 GND.n1627 585
R8924 GND.n4332 GND.n1627 585
R8925 GND.n3374 GND.n3373 585
R8926 GND.n3373 GND.n3372 585
R8927 GND.n3375 GND.n1619 585
R8928 GND.n4338 GND.n1619 585
R8929 GND.n3378 GND.n3377 585
R8930 GND.n3377 GND.n3376 585
R8931 GND.n3379 GND.n2199 585
R8932 GND.n3393 GND.n2199 585
R8933 GND.n3381 GND.n3380 585
R8934 GND.n3380 GND.n2198 585
R8935 GND.n3382 GND.n2206 585
R8936 GND.n2206 GND.n1603 585
R8937 GND.n3384 GND.n3383 585
R8938 GND.n3386 GND.n3384 585
R8939 GND.n3370 GND.n2205 585
R8940 GND.n2205 GND.n2204 585
R8941 GND.n3369 GND.n1584 585
R8942 GND.n4353 GND.n1584 585
R8943 GND.n3368 GND.n3367 585
R8944 GND.n3367 GND.n3366 585
R8945 GND.n3365 GND.n1576 585
R8946 GND.n4359 GND.n1576 585
R8947 GND.n3364 GND.n3363 585
R8948 GND.n3363 GND.n3362 585
R8949 GND.n3359 GND.n3358 585
R8950 GND.n3360 GND.n3359 585
R8951 GND.n3357 GND.n1560 585
R8952 GND.n4367 GND.n1560 585
R8953 GND.n3356 GND.n3355 585
R8954 GND.n3355 GND.n3354 585
R8955 GND.n3353 GND.n1552 585
R8956 GND.n4373 GND.n1552 585
R8957 GND.n3352 GND.n3351 585
R8958 GND.n3351 GND.n3350 585
R8959 GND.n2208 GND.n2207 585
R8960 GND.n2210 GND.n2208 585
R8961 GND.n3308 GND.n2218 585
R8962 GND.n2218 GND.n1541 585
R8963 GND.n3310 GND.n3309 585
R8964 GND.n3319 GND.n3310 585
R8965 GND.n3307 GND.n2217 585
R8966 GND.n2217 GND.n2216 585
R8967 GND.n3306 GND.n3305 585
R8968 GND.n3305 GND.n3304 585
R8969 GND.n3302 GND.n1531 585
R8970 GND.n4388 GND.n1531 585
R8971 GND.n3301 GND.n3300 585
R8972 GND.n3300 GND.n3299 585
R8973 GND.n3298 GND.n1521 585
R8974 GND.n4394 GND.n1521 585
R8975 GND.n3297 GND.n3296 585
R8976 GND.n3296 GND.n1520 585
R8977 GND.n3295 GND.n2219 585
R8978 GND.n3295 GND.n3294 585
R8979 GND.n3136 GND.n2220 585
R8980 GND.n2220 GND.n1512 585
R8981 GND.n3137 GND.n1511 585
R8982 GND.n4402 GND.n1511 585
R8983 GND.n3141 GND.n3140 585
R8984 GND.n3140 GND.n3139 585
R8985 GND.n3142 GND.n1503 585
R8986 GND.n4408 GND.n1503 585
R8987 GND.n3144 GND.n3143 585
R8988 GND.n3144 GND.n1502 585
R8989 GND.n3145 GND.n3135 585
R8990 GND.n3145 GND.n2230 585
R8991 GND.n3147 GND.n3146 585
R8992 GND.n3146 GND.n1494 585
R8993 GND.n3148 GND.n1493 585
R8994 GND.n4416 GND.n1493 585
R8995 GND.n3151 GND.n3150 585
R8996 GND.n3150 GND.n3149 585
R8997 GND.n3152 GND.n1486 585
R8998 GND.n4422 GND.n1486 585
R8999 GND.n3154 GND.n3153 585
R9000 GND.n3153 GND.n1485 585
R9001 GND.n3155 GND.n2242 585
R9002 GND.n3231 GND.n2242 585
R9003 GND.n3156 GND.n3069 585
R9004 GND.n3069 GND.n1474 585
R9005 GND.n2541 GND.n2540 585
R9006 GND.n2542 GND.n2541 585
R9007 GND.n5480 GND.n5479 585
R9008 GND.n5480 GND.n573 585
R9009 GND.n5482 GND.n5481 585
R9010 GND.n5481 GND.n583 585
R9011 GND.n5483 GND.n596 585
R9012 GND.n596 GND.n580 585
R9013 GND.n5485 GND.n5484 585
R9014 GND.n5486 GND.n5485 585
R9015 GND.n597 GND.n595 585
R9016 GND.n1944 GND.n595 585
R9017 GND.n4109 GND.n4108 585
R9018 GND.n4109 GND.n1943 585
R9019 GND.n4111 GND.n4110 585
R9020 GND.n4110 GND.n1954 585
R9021 GND.n4112 GND.n1958 585
R9022 GND.n1958 GND.n1951 585
R9023 GND.n4114 GND.n4113 585
R9024 GND.n4115 GND.n4114 585
R9025 GND.n1959 GND.n1957 585
R9026 GND.n1965 GND.n1957 585
R9027 GND.n4100 GND.n4099 585
R9028 GND.n4099 GND.n4098 585
R9029 GND.n1962 GND.n1961 585
R9030 GND.n1976 GND.n1962 585
R9031 GND.n4079 GND.n1982 585
R9032 GND.n1982 GND.n1974 585
R9033 GND.n4081 GND.n4080 585
R9034 GND.n4082 GND.n4081 585
R9035 GND.n1983 GND.n1981 585
R9036 GND.n1989 GND.n1981 585
R9037 GND.n4074 GND.n4073 585
R9038 GND.n4073 GND.n4072 585
R9039 GND.n1986 GND.n1985 585
R9040 GND.n4029 GND.n1986 585
R9041 GND.n4038 GND.n4037 585
R9042 GND.n4039 GND.n4038 585
R9043 GND.n4035 GND.n4033 585
R9044 GND.n4033 GND.n4027 585
R9045 GND.n4010 GND.n4009 585
R9046 GND.n4014 GND.n4010 585
R9047 GND.n4051 GND.n4050 585
R9048 GND.n4050 GND.n4049 585
R9049 GND.n4053 GND.n2013 585
R9050 GND.n4011 GND.n2013 585
R9051 GND.n4055 GND.n4054 585
R9052 GND.n4056 GND.n4055 585
R9053 GND.n4007 GND.n2012 585
R9054 GND.n2012 GND.n2008 585
R9055 GND.n4006 GND.n4005 585
R9056 GND.n4005 GND.n2002 585
R9057 GND.n4004 GND.n2016 585
R9058 GND.n4004 GND.n4003 585
R9059 GND.n3973 GND.n2015 585
R9060 GND.n2025 GND.n2015 585
R9061 GND.n3974 GND.n2045 585
R9062 GND.n2045 GND.n2024 585
R9063 GND.n3976 GND.n3975 585
R9064 GND.n3977 GND.n3976 585
R9065 GND.n2046 GND.n2044 585
R9066 GND.n2044 GND.n2038 585
R9067 GND.n3967 GND.n3966 585
R9068 GND.n3966 GND.n2036 585
R9069 GND.n3965 GND.n2048 585
R9070 GND.n3965 GND.n3964 585
R9071 GND.n3866 GND.n2049 585
R9072 GND.n2059 GND.n2049 585
R9073 GND.n3868 GND.n3867 585
R9074 GND.n3868 GND.n2058 585
R9075 GND.n3870 GND.n3869 585
R9076 GND.n3869 GND.n2070 585
R9077 GND.n3871 GND.n3859 585
R9078 GND.n3859 GND.n2068 585
R9079 GND.n3873 GND.n3872 585
R9080 GND.n3873 GND.n2072 585
R9081 GND.n3876 GND.n3858 585
R9082 GND.n3876 GND.n3875 585
R9083 GND.n3878 GND.n3877 585
R9084 GND.n3877 GND.n2080 585
R9085 GND.n3879 GND.n3853 585
R9086 GND.n3853 GND.n2092 585
R9087 GND.n3881 GND.n3880 585
R9088 GND.n3881 GND.n2089 585
R9089 GND.n3882 GND.n3852 585
R9090 GND.n3882 GND.n2095 585
R9091 GND.n3884 GND.n3883 585
R9092 GND.n3883 GND.n2103 585
R9093 GND.n3885 GND.n2117 585
R9094 GND.n2117 GND.n2102 585
R9095 GND.n3887 GND.n3886 585
R9096 GND.n3888 GND.n3887 585
R9097 GND.n2118 GND.n2116 585
R9098 GND.n2116 GND.n2112 585
R9099 GND.n3846 GND.n3845 585
R9100 GND.n3845 GND.n3844 585
R9101 GND.n2135 GND.n2120 585
R9102 GND.n2136 GND.n2135 585
R9103 GND.n2134 GND.n2133 585
R9104 GND.n2134 GND.n1851 585
R9105 GND.n2122 GND.n2121 585
R9106 GND.n2121 GND.n1822 585
R9107 GND.n2129 GND.n2128 585
R9108 GND.n2128 GND.n2127 585
R9109 GND.n2126 GND.n2125 585
R9110 GND.n2126 GND.n1761 585
R9111 GND.n1758 GND.n1757 585
R9112 GND.n4255 GND.n1758 585
R9113 GND.n4258 GND.n4257 585
R9114 GND.n4257 GND.n4256 585
R9115 GND.n4259 GND.n1750 585
R9116 GND.n1759 GND.n1750 585
R9117 GND.n4261 GND.n4260 585
R9118 GND.n4262 GND.n4261 585
R9119 GND.n1751 GND.n1749 585
R9120 GND.n3804 GND.n1749 585
R9121 GND.n1732 GND.n1731 585
R9122 GND.n1736 GND.n1732 585
R9123 GND.n4272 GND.n4271 585
R9124 GND.n4271 GND.n4270 585
R9125 GND.n4273 GND.n1724 585
R9126 GND.n1733 GND.n1724 585
R9127 GND.n4275 GND.n4274 585
R9128 GND.n4276 GND.n4275 585
R9129 GND.n1725 GND.n1723 585
R9130 GND.n1723 GND.n1720 585
R9131 GND.n1705 GND.n1704 585
R9132 GND.n1709 GND.n1705 585
R9133 GND.n4286 GND.n4285 585
R9134 GND.n4285 GND.n4284 585
R9135 GND.n4287 GND.n1699 585
R9136 GND.n1706 GND.n1699 585
R9137 GND.n4289 GND.n4288 585
R9138 GND.n4290 GND.n4289 585
R9139 GND.n1700 GND.n1698 585
R9140 GND.n3756 GND.n1698 585
R9141 GND.n3771 GND.n3770 585
R9142 GND.n3772 GND.n3771 585
R9143 GND.n3759 GND.n3758 585
R9144 GND.n3758 GND.n1686 585
R9145 GND.n3765 GND.n3764 585
R9146 GND.n3764 GND.n2177 585
R9147 GND.n3763 GND.n3762 585
R9148 GND.n3763 GND.n1678 585
R9149 GND.n1661 GND.n1660 585
R9150 GND.n2180 GND.n1661 585
R9151 GND.n4314 GND.n4313 585
R9152 GND.n4313 GND.n4312 585
R9153 GND.n4315 GND.n1655 585
R9154 GND.n2186 GND.n1655 585
R9155 GND.n4317 GND.n4316 585
R9156 GND.n4318 GND.n4317 585
R9157 GND.n1656 GND.n1654 585
R9158 GND.n1654 GND.n1645 585
R9159 GND.n3416 GND.n3415 585
R9160 GND.n3417 GND.n3416 585
R9161 GND.n3410 GND.n3409 585
R9162 GND.n3409 GND.n1629 585
R9163 GND.n1617 GND.n1616 585
R9164 GND.n1626 GND.n1617 585
R9165 GND.n4341 GND.n4340 585
R9166 GND.n4340 GND.n4339 585
R9167 GND.n4342 GND.n1606 585
R9168 GND.n2200 GND.n1606 585
R9169 GND.n4344 GND.n4343 585
R9170 GND.n4345 GND.n4344 585
R9171 GND.n1607 GND.n1605 585
R9172 GND.n3385 GND.n1605 585
R9173 GND.n1610 GND.n1609 585
R9174 GND.n1609 GND.n1586 585
R9175 GND.n1574 GND.n1573 585
R9176 GND.n1583 GND.n1574 585
R9177 GND.n4362 GND.n4361 585
R9178 GND.n4361 GND.n4360 585
R9179 GND.n4363 GND.n1563 585
R9180 GND.n3361 GND.n1563 585
R9181 GND.n4365 GND.n4364 585
R9182 GND.n4366 GND.n4365 585
R9183 GND.n1564 GND.n1562 585
R9184 GND.n1562 GND.n1553 585
R9185 GND.n1567 GND.n1566 585
R9186 GND.n1566 GND.n1550 585
R9187 GND.n1539 GND.n1538 585
R9188 GND.n2209 GND.n1539 585
R9189 GND.n4383 GND.n4382 585
R9190 GND.n4382 GND.n4381 585
R9191 GND.n4384 GND.n1533 585
R9192 GND.n3303 GND.n1533 585
R9193 GND.n4386 GND.n4385 585
R9194 GND.n4387 GND.n4386 585
R9195 GND.n1519 GND.n1518 585
R9196 GND.n1523 GND.n1519 585
R9197 GND.n4397 GND.n4396 585
R9198 GND.n4396 GND.n4395 585
R9199 GND.n4398 GND.n1513 585
R9200 GND.n3255 GND.n1513 585
R9201 GND.n4400 GND.n4399 585
R9202 GND.n4401 GND.n4400 585
R9203 GND.n1501 GND.n1500 585
R9204 GND.n3138 GND.n1501 585
R9205 GND.n4411 GND.n4410 585
R9206 GND.n4410 GND.n4409 585
R9207 GND.n4412 GND.n1495 585
R9208 GND.n2231 GND.n1495 585
R9209 GND.n4414 GND.n4413 585
R9210 GND.n4415 GND.n4414 585
R9211 GND.n1484 GND.n1483 585
R9212 GND.n2240 GND.n1484 585
R9213 GND.n4425 GND.n4424 585
R9214 GND.n4424 GND.n4423 585
R9215 GND.n4426 GND.n1476 585
R9216 GND.n3232 GND.n1476 585
R9217 GND.n4428 GND.n4427 585
R9218 GND.n4429 GND.n4428 585
R9219 GND.n1477 GND.n1475 585
R9220 GND.n1475 GND.n1472 585
R9221 GND.n1457 GND.n1456 585
R9222 GND.n1461 GND.n1457 585
R9223 GND.n4439 GND.n4438 585
R9224 GND.n4438 GND.n4437 585
R9225 GND.n4440 GND.n1449 585
R9226 GND.n1458 GND.n1449 585
R9227 GND.n4442 GND.n4441 585
R9228 GND.n4443 GND.n4442 585
R9229 GND.n1450 GND.n1448 585
R9230 GND.n1448 GND.n1445 585
R9231 GND.n1430 GND.n1429 585
R9232 GND.n1434 GND.n1430 585
R9233 GND.n4453 GND.n4452 585
R9234 GND.n4452 GND.n4451 585
R9235 GND.n4454 GND.n1416 585
R9236 GND.n1431 GND.n1416 585
R9237 GND.n4456 GND.n4455 585
R9238 GND.n4457 GND.n4456 585
R9239 GND.n1417 GND.n1415 585
R9240 GND.n1415 GND.n1412 585
R9241 GND.n1423 GND.n1422 585
R9242 GND.n1422 GND.n1403 585
R9243 GND.n1421 GND.n1399 585
R9244 GND.n4465 GND.n1399 585
R9245 GND.n4468 GND.n1400 585
R9246 GND.n4468 GND.n4467 585
R9247 GND.n4469 GND.n1398 585
R9248 GND.n4469 GND.n1339 585
R9249 GND.n4471 GND.n4470 585
R9250 GND.n4470 GND.n1325 585
R9251 GND.n4472 GND.n1393 585
R9252 GND.n1393 GND.n1391 585
R9253 GND.n4474 GND.n4473 585
R9254 GND.n4475 GND.n4474 585
R9255 GND.n1394 GND.n1392 585
R9256 GND.n1392 GND.n1376 585
R9257 GND.n2924 GND.n2923 585
R9258 GND.n2924 GND.n1263 585
R9259 GND.n2926 GND.n2925 585
R9260 GND.n2925 GND.n1261 585
R9261 GND.n2927 GND.n2309 585
R9262 GND.n2309 GND.n2289 585
R9263 GND.n2929 GND.n2928 585
R9264 GND.n2930 GND.n2929 585
R9265 GND.n2310 GND.n2308 585
R9266 GND.n2308 GND.n2298 585
R9267 GND.n2915 GND.n2914 585
R9268 GND.n2914 GND.n2296 585
R9269 GND.n2913 GND.n2312 585
R9270 GND.n2913 GND.n2301 585
R9271 GND.n2912 GND.n2314 585
R9272 GND.n2912 GND.n2911 585
R9273 GND.n2774 GND.n2313 585
R9274 GND.n2324 GND.n2313 585
R9275 GND.n2776 GND.n2775 585
R9276 GND.n2775 GND.n2322 585
R9277 GND.n2777 GND.n2767 585
R9278 GND.n2767 GND.n2766 585
R9279 GND.n2779 GND.n2778 585
R9280 GND.n2779 GND.n2335 585
R9281 GND.n2780 GND.n2764 585
R9282 GND.n2780 GND.n2333 585
R9283 GND.n2782 GND.n2781 585
R9284 GND.n2781 GND.n2345 585
R9285 GND.n2783 GND.n2759 585
R9286 GND.n2759 GND.n2343 585
R9287 GND.n2788 GND.n2784 585
R9288 GND.n2788 GND.n2787 585
R9289 GND.n2789 GND.n2758 585
R9290 GND.n2789 GND.n2354 585
R9291 GND.n2791 GND.n2790 585
R9292 GND.n2790 GND.n2353 585
R9293 GND.n2792 GND.n2753 585
R9294 GND.n2753 GND.n2364 585
R9295 GND.n2794 GND.n2793 585
R9296 GND.n2794 GND.n2362 585
R9297 GND.n2797 GND.n2752 585
R9298 GND.n2797 GND.n2796 585
R9299 GND.n2799 GND.n2798 585
R9300 GND.n2798 GND.n2374 585
R9301 GND.n2800 GND.n2748 585
R9302 GND.n2748 GND.n2373 585
R9303 GND.n2803 GND.n2802 585
R9304 GND.n2804 GND.n2803 585
R9305 GND.n2750 GND.n2747 585
R9306 GND.n2747 GND.n2417 585
R9307 GND.n2401 GND.n2400 585
R9308 GND.n2405 GND.n2401 585
R9309 GND.n2816 GND.n2815 585
R9310 GND.n2815 GND.n2814 585
R9311 GND.n2818 GND.n2398 585
R9312 GND.n2402 GND.n2398 585
R9313 GND.n2820 GND.n2819 585
R9314 GND.n2821 GND.n2820 585
R9315 GND.n2723 GND.n2397 585
R9316 GND.n2397 GND.n2391 585
R9317 GND.n2724 GND.n2429 585
R9318 GND.n2429 GND.n2389 585
R9319 GND.n2727 GND.n2726 585
R9320 GND.n2728 GND.n2727 585
R9321 GND.n2722 GND.n2428 585
R9322 GND.n2687 GND.n2428 585
R9323 GND.n2434 GND.n2430 585
R9324 GND.n2686 GND.n2434 585
R9325 GND.n2718 GND.n2717 585
R9326 GND.n2717 GND.n2716 585
R9327 GND.n2433 GND.n2432 585
R9328 GND.n2449 GND.n2433 585
R9329 GND.n2522 GND.n2521 585
R9330 GND.n2522 GND.n2446 585
R9331 GND.n2524 GND.n2523 585
R9332 GND.n2523 GND.n2452 585
R9333 GND.n2525 GND.n2515 585
R9334 GND.n2515 GND.n2460 585
R9335 GND.n2527 GND.n2526 585
R9336 GND.n2527 GND.n2459 585
R9337 GND.n2528 GND.n2514 585
R9338 GND.n2528 GND.n2471 585
R9339 GND.n2530 GND.n2529 585
R9340 GND.n2529 GND.n2469 585
R9341 GND.n2531 GND.n2509 585
R9342 GND.n2509 GND.n2474 585
R9343 GND.n2533 GND.n2532 585
R9344 GND.n2533 GND.n2483 585
R9345 GND.n2534 GND.n2508 585
R9346 GND.n2534 GND.n2481 585
R9347 GND.n2536 GND.n2535 585
R9348 GND.n2535 GND.n2494 585
R9349 GND.n2537 GND.n2505 585
R9350 GND.n2505 GND.n2492 585
R9351 GND.n4213 GND.n4212 585
R9352 GND.n4214 GND.n4213 585
R9353 GND.n4211 GND.n1853 585
R9354 GND.n4204 GND.n4203 585
R9355 GND.n4202 GND.n1781 585
R9356 GND.n4249 GND.n1782 585
R9357 GND.n4248 GND.n1783 585
R9358 GND.n1843 GND.n1784 585
R9359 GND.n4241 GND.n1790 585
R9360 GND.n4240 GND.n1791 585
R9361 GND.n1846 GND.n1792 585
R9362 GND.n4233 GND.n1800 585
R9363 GND.n4232 GND.n1801 585
R9364 GND.n1848 GND.n1802 585
R9365 GND.n4225 GND.n1808 585
R9366 GND.n4224 GND.n1809 585
R9367 GND.n1821 GND.n1812 585
R9368 GND.n4217 GND.n4216 585
R9369 GND.n5570 GND.n5569 585
R9370 GND.n5569 GND.n467 585
R9371 GND.n5523 GND.n554 585
R9372 GND.n5523 GND.n5522 585
R9373 GND.n567 GND.n555 585
R9374 GND.n556 GND.n555 585
R9375 GND.n5512 GND.n5511 585
R9376 GND.n5513 GND.n5512 585
R9377 GND.n566 GND.n565 585
R9378 GND.n565 GND.n562 585
R9379 GND.n589 GND.n574 585
R9380 GND.n5503 GND.n574 585
R9381 GND.n587 GND.n585 585
R9382 GND.n585 GND.n572 585
R9383 GND.n5494 GND.n5493 585
R9384 GND.n5495 GND.n5494 585
R9385 GND.n586 GND.n584 585
R9386 GND.n5487 GND.n584 585
R9387 GND.n4133 GND.n4132 585
R9388 GND.n4132 GND.n594 585
R9389 GND.n4131 GND.n1940 585
R9390 GND.n4131 GND.n4130 585
R9391 GND.n1942 GND.n1941 585
R9392 GND.n1953 GND.n1942 585
R9393 GND.n4119 GND.n1935 585
R9394 GND.n4120 GND.n4119 585
R9395 GND.n4118 GND.n1934 585
R9396 GND.n4118 GND.n4117 585
R9397 GND.n1955 GND.n1933 585
R9398 GND.n1956 GND.n1955 585
R9399 GND.n1967 GND.n1966 585
R9400 GND.n4097 GND.n1967 585
R9401 GND.n4085 GND.n1927 585
R9402 GND.n4085 GND.n1963 585
R9403 GND.n4086 GND.n1926 585
R9404 GND.n4087 GND.n4086 585
R9405 GND.n4084 GND.n1925 585
R9406 GND.n4084 GND.n4083 585
R9407 GND.n1978 GND.n1977 585
R9408 GND.n1980 GND.n1978 585
R9409 GND.n1990 GND.n1919 585
R9410 GND.n4071 GND.n1990 585
R9411 GND.n4024 GND.n1918 585
R9412 GND.n4024 GND.n1988 585
R9413 GND.n4025 GND.n1917 585
R9414 GND.n4032 GND.n4025 585
R9415 GND.n4041 GND.n4026 585
R9416 GND.n4041 GND.n4040 585
R9417 GND.n4042 GND.n1911 585
R9418 GND.n4043 GND.n4042 585
R9419 GND.n4016 GND.n1910 585
R9420 GND.n4048 GND.n4016 585
R9421 GND.n4015 GND.n1909 585
R9422 GND.n4015 GND.n4012 585
R9423 GND.n2007 GND.n2006 585
R9424 GND.n2011 GND.n2007 585
R9425 GND.n4058 GND.n1903 585
R9426 GND.n4058 GND.n4057 585
R9427 GND.n4059 GND.n1902 585
R9428 GND.n4060 GND.n4059 585
R9429 GND.n2005 GND.n1901 585
R9430 GND.n4002 GND.n2005 585
R9431 GND.n2027 GND.n2026 585
R9432 GND.n2027 GND.n2017 585
R9433 GND.n2028 GND.n1895 585
R9434 GND.n3991 GND.n2028 585
R9435 GND.n2040 GND.n1894 585
R9436 GND.n2043 GND.n2040 585
R9437 GND.n3979 GND.n1893 585
R9438 GND.n3979 GND.n3978 585
R9439 GND.n3981 GND.n3980 585
R9440 GND.n3982 GND.n3981 585
R9441 GND.n2039 GND.n1887 585
R9442 GND.n3963 GND.n2039 585
R9443 GND.n2060 GND.n1886 585
R9444 GND.n2060 GND.n2051 585
R9445 GND.n2061 GND.n1885 585
R9446 GND.n3952 GND.n2061 585
R9447 GND.n3940 GND.n3938 585
R9448 GND.n3940 GND.n3939 585
R9449 GND.n3941 GND.n1879 585
R9450 GND.n3942 GND.n3941 585
R9451 GND.n3937 GND.n1878 585
R9452 GND.n3937 GND.n3936 585
R9453 GND.n2071 GND.n1877 585
R9454 GND.n3874 GND.n2071 585
R9455 GND.n2082 GND.n2081 585
R9456 GND.n3927 GND.n2082 585
R9457 GND.n3915 GND.n1871 585
R9458 GND.n3915 GND.n3914 585
R9459 GND.n3916 GND.n1870 585
R9460 GND.n3917 GND.n3916 585
R9461 GND.n3913 GND.n1869 585
R9462 GND.n3913 GND.n3912 585
R9463 GND.n2094 GND.n2093 585
R9464 GND.n2106 GND.n2094 585
R9465 GND.n2104 GND.n1863 585
R9466 GND.n3903 GND.n2104 585
R9467 GND.n3891 GND.n1862 585
R9468 GND.n3891 GND.n3890 585
R9469 GND.n3892 GND.n1861 585
R9470 GND.n3893 GND.n3892 585
R9471 GND.n2115 GND.n2114 585
R9472 GND.n3843 GND.n2115 585
R9473 GND.n1855 GND.n1852 585
R9474 GND.n2137 GND.n1852 585
R9475 GND.n5632 GND.n5631 585
R9476 GND.n5631 GND.n5630 585
R9477 GND.n466 GND.n465 585
R9478 GND.n5545 GND.n5544 585
R9479 GND.n5543 GND.n5542 585
R9480 GND.n5549 GND.n5541 585
R9481 GND.n5550 GND.n5540 585
R9482 GND.n5551 GND.n5539 585
R9483 GND.n5538 GND.n5536 585
R9484 GND.n5555 GND.n5535 585
R9485 GND.n5556 GND.n5534 585
R9486 GND.n5557 GND.n5533 585
R9487 GND.n5532 GND.n5530 585
R9488 GND.n5561 GND.n5529 585
R9489 GND.n5562 GND.n5528 585
R9490 GND.n5563 GND.n5527 585
R9491 GND.n5526 GND.n5524 585
R9492 GND.n5568 GND.n5567 585
R9493 GND.n5635 GND.n461 585
R9494 GND.n467 GND.n461 585
R9495 GND.n5636 GND.n460 585
R9496 GND.n5522 GND.n460 585
R9497 GND.n5637 GND.n459 585
R9498 GND.n556 GND.n459 585
R9499 GND.n564 GND.n457 585
R9500 GND.n5513 GND.n564 585
R9501 GND.n5641 GND.n456 585
R9502 GND.n562 GND.n456 585
R9503 GND.n5642 GND.n455 585
R9504 GND.n5503 GND.n455 585
R9505 GND.n5643 GND.n454 585
R9506 GND.n572 GND.n454 585
R9507 GND.n582 GND.n452 585
R9508 GND.n5495 GND.n582 585
R9509 GND.n5647 GND.n451 585
R9510 GND.n5487 GND.n451 585
R9511 GND.n5648 GND.n450 585
R9512 GND.n594 GND.n450 585
R9513 GND.n5649 GND.n449 585
R9514 GND.n4130 GND.n449 585
R9515 GND.n1952 GND.n447 585
R9516 GND.n1953 GND.n1952 585
R9517 GND.n5653 GND.n446 585
R9518 GND.n4120 GND.n446 585
R9519 GND.n5654 GND.n445 585
R9520 GND.n4117 GND.n445 585
R9521 GND.n5655 GND.n444 585
R9522 GND.n1956 GND.n444 585
R9523 GND.n1964 GND.n442 585
R9524 GND.n4097 GND.n1964 585
R9525 GND.n5659 GND.n441 585
R9526 GND.n1963 GND.n441 585
R9527 GND.n5660 GND.n440 585
R9528 GND.n4087 GND.n440 585
R9529 GND.n5661 GND.n439 585
R9530 GND.n4083 GND.n439 585
R9531 GND.n1979 GND.n437 585
R9532 GND.n1980 GND.n1979 585
R9533 GND.n5665 GND.n436 585
R9534 GND.n4071 GND.n436 585
R9535 GND.n5666 GND.n435 585
R9536 GND.n1988 GND.n435 585
R9537 GND.n5667 GND.n434 585
R9538 GND.n4032 GND.n434 585
R9539 GND.n4028 GND.n432 585
R9540 GND.n4040 GND.n4028 585
R9541 GND.n5671 GND.n431 585
R9542 GND.n4043 GND.n431 585
R9543 GND.n5672 GND.n430 585
R9544 GND.n4048 GND.n430 585
R9545 GND.n5673 GND.n429 585
R9546 GND.n4012 GND.n429 585
R9547 GND.n2010 GND.n428 585
R9548 GND.n2011 GND.n2010 585
R9549 GND.n3996 GND.n2009 585
R9550 GND.n4057 GND.n2009 585
R9551 GND.n2020 GND.n2004 585
R9552 GND.n4060 GND.n2004 585
R9553 GND.n4001 GND.n4000 585
R9554 GND.n4002 GND.n4001 585
R9555 GND.n2019 GND.n2018 585
R9556 GND.n2018 GND.n2017 585
R9557 GND.n3993 GND.n3992 585
R9558 GND.n3992 GND.n3991 585
R9559 GND.n2023 GND.n2022 585
R9560 GND.n2043 GND.n2023 585
R9561 GND.n3957 GND.n2041 585
R9562 GND.n3978 GND.n2041 585
R9563 GND.n2054 GND.n2037 585
R9564 GND.n3982 GND.n2037 585
R9565 GND.n3962 GND.n3961 585
R9566 GND.n3963 GND.n3962 585
R9567 GND.n2053 GND.n2052 585
R9568 GND.n2052 GND.n2051 585
R9569 GND.n3954 GND.n3953 585
R9570 GND.n3953 GND.n3952 585
R9571 GND.n2057 GND.n2056 585
R9572 GND.n3939 GND.n2057 585
R9573 GND.n2076 GND.n2069 585
R9574 GND.n3942 GND.n2069 585
R9575 GND.n3935 GND.n3934 585
R9576 GND.n3936 GND.n3935 585
R9577 GND.n2075 GND.n2074 585
R9578 GND.n3874 GND.n2074 585
R9579 GND.n3929 GND.n3928 585
R9580 GND.n3928 GND.n3927 585
R9581 GND.n2079 GND.n2078 585
R9582 GND.n3914 GND.n2079 585
R9583 GND.n2098 GND.n2091 585
R9584 GND.n3917 GND.n2091 585
R9585 GND.n3911 GND.n3910 585
R9586 GND.n3912 GND.n3911 585
R9587 GND.n2097 GND.n2096 585
R9588 GND.n2106 GND.n2096 585
R9589 GND.n3905 GND.n3904 585
R9590 GND.n3904 GND.n3903 585
R9591 GND.n2101 GND.n2100 585
R9592 GND.n3890 GND.n2101 585
R9593 GND.n2139 GND.n2113 585
R9594 GND.n3893 GND.n2113 585
R9595 GND.n3842 GND.n3841 585
R9596 GND.n3843 GND.n3842 585
R9597 GND.n2138 GND.n1820 585
R9598 GND.n2137 GND.n1820 585
R9599 GND.n3514 GND.n1685 511.721
R9600 GND.n3774 GND.n3456 511.721
R9601 GND.n3158 GND.n3069 511.721
R9602 GND.n3225 GND.n2243 511.721
R9603 GND.n4882 GND.n953 477.627
R9604 GND.n3070 GND.t89 371.625
R9605 GND.n3689 GND.t106 371.625
R9606 GND.n3161 GND.t128 371.625
R9607 GND.n3492 GND.t67 371.625
R9608 GND.n2158 GND.t131 291.267
R9609 GND.n2988 GND.t124 291.267
R9610 GND.n95 GND.n69 289.615
R9611 GND.n132 GND.n106 289.615
R9612 GND.n164 GND.n138 289.615
R9613 GND.n201 GND.n175 289.615
R9614 GND.n26 GND.n0 289.615
R9615 GND.n63 GND.n37 289.615
R9616 GND.n280 GND.n254 289.615
R9617 GND.n243 GND.n217 289.615
R9618 GND.n349 GND.n323 289.615
R9619 GND.n312 GND.n286 289.615
R9620 GND.n419 GND.n393 289.615
R9621 GND.n382 GND.n356 289.615
R9622 GND.n4890 GND.n953 280.613
R9623 GND.n4891 GND.n4890 280.613
R9624 GND.n4892 GND.n4891 280.613
R9625 GND.n4892 GND.n947 280.613
R9626 GND.n4900 GND.n947 280.613
R9627 GND.n4901 GND.n4900 280.613
R9628 GND.n4902 GND.n4901 280.613
R9629 GND.n4902 GND.n941 280.613
R9630 GND.n4910 GND.n941 280.613
R9631 GND.n4911 GND.n4910 280.613
R9632 GND.n4912 GND.n4911 280.613
R9633 GND.n4912 GND.n935 280.613
R9634 GND.n4920 GND.n935 280.613
R9635 GND.n4921 GND.n4920 280.613
R9636 GND.n4922 GND.n4921 280.613
R9637 GND.n4922 GND.n929 280.613
R9638 GND.n4930 GND.n929 280.613
R9639 GND.n4931 GND.n4930 280.613
R9640 GND.n4932 GND.n4931 280.613
R9641 GND.n4932 GND.n923 280.613
R9642 GND.n4940 GND.n923 280.613
R9643 GND.n4941 GND.n4940 280.613
R9644 GND.n4942 GND.n4941 280.613
R9645 GND.n4942 GND.n917 280.613
R9646 GND.n4950 GND.n917 280.613
R9647 GND.n4951 GND.n4950 280.613
R9648 GND.n4952 GND.n4951 280.613
R9649 GND.n4952 GND.n911 280.613
R9650 GND.n4960 GND.n911 280.613
R9651 GND.n4961 GND.n4960 280.613
R9652 GND.n4962 GND.n4961 280.613
R9653 GND.n4962 GND.n905 280.613
R9654 GND.n4970 GND.n905 280.613
R9655 GND.n4971 GND.n4970 280.613
R9656 GND.n4972 GND.n4971 280.613
R9657 GND.n4972 GND.n899 280.613
R9658 GND.n4980 GND.n899 280.613
R9659 GND.n4981 GND.n4980 280.613
R9660 GND.n4982 GND.n4981 280.613
R9661 GND.n4982 GND.n893 280.613
R9662 GND.n4990 GND.n893 280.613
R9663 GND.n4991 GND.n4990 280.613
R9664 GND.n4992 GND.n4991 280.613
R9665 GND.n4992 GND.n887 280.613
R9666 GND.n5000 GND.n887 280.613
R9667 GND.n5001 GND.n5000 280.613
R9668 GND.n5002 GND.n5001 280.613
R9669 GND.n5002 GND.n881 280.613
R9670 GND.n5010 GND.n881 280.613
R9671 GND.n5011 GND.n5010 280.613
R9672 GND.n5012 GND.n5011 280.613
R9673 GND.n5012 GND.n875 280.613
R9674 GND.n5020 GND.n875 280.613
R9675 GND.n5021 GND.n5020 280.613
R9676 GND.n5022 GND.n5021 280.613
R9677 GND.n5022 GND.n869 280.613
R9678 GND.n5030 GND.n869 280.613
R9679 GND.n5031 GND.n5030 280.613
R9680 GND.n5032 GND.n5031 280.613
R9681 GND.n5032 GND.n863 280.613
R9682 GND.n5040 GND.n863 280.613
R9683 GND.n5041 GND.n5040 280.613
R9684 GND.n5042 GND.n5041 280.613
R9685 GND.n5042 GND.n857 280.613
R9686 GND.n5050 GND.n857 280.613
R9687 GND.n5051 GND.n5050 280.613
R9688 GND.n5052 GND.n5051 280.613
R9689 GND.n5052 GND.n851 280.613
R9690 GND.n5060 GND.n851 280.613
R9691 GND.n5061 GND.n5060 280.613
R9692 GND.n5062 GND.n5061 280.613
R9693 GND.n5062 GND.n845 280.613
R9694 GND.n5070 GND.n845 280.613
R9695 GND.n5071 GND.n5070 280.613
R9696 GND.n5072 GND.n5071 280.613
R9697 GND.n5072 GND.n839 280.613
R9698 GND.n5080 GND.n839 280.613
R9699 GND.n5081 GND.n5080 280.613
R9700 GND.n5082 GND.n5081 280.613
R9701 GND.n5082 GND.n833 280.613
R9702 GND.n5090 GND.n833 280.613
R9703 GND.n5091 GND.n5090 280.613
R9704 GND.n5092 GND.n5091 280.613
R9705 GND.n5092 GND.n827 280.613
R9706 GND.n5100 GND.n827 280.613
R9707 GND.n5101 GND.n5100 280.613
R9708 GND.n5102 GND.n5101 280.613
R9709 GND.n5102 GND.n821 280.613
R9710 GND.n5110 GND.n821 280.613
R9711 GND.n5111 GND.n5110 280.613
R9712 GND.n5112 GND.n5111 280.613
R9713 GND.n5112 GND.n815 280.613
R9714 GND.n5120 GND.n815 280.613
R9715 GND.n5121 GND.n5120 280.613
R9716 GND.n5122 GND.n5121 280.613
R9717 GND.n5122 GND.n809 280.613
R9718 GND.n5130 GND.n809 280.613
R9719 GND.n5131 GND.n5130 280.613
R9720 GND.n5132 GND.n5131 280.613
R9721 GND.n5132 GND.n803 280.613
R9722 GND.n5140 GND.n803 280.613
R9723 GND.n5141 GND.n5140 280.613
R9724 GND.n5142 GND.n5141 280.613
R9725 GND.n5142 GND.n797 280.613
R9726 GND.n5150 GND.n797 280.613
R9727 GND.n5151 GND.n5150 280.613
R9728 GND.n5152 GND.n5151 280.613
R9729 GND.n5152 GND.n791 280.613
R9730 GND.n5160 GND.n791 280.613
R9731 GND.n5161 GND.n5160 280.613
R9732 GND.n5162 GND.n5161 280.613
R9733 GND.n5162 GND.n785 280.613
R9734 GND.n5170 GND.n785 280.613
R9735 GND.n5171 GND.n5170 280.613
R9736 GND.n5172 GND.n5171 280.613
R9737 GND.n5172 GND.n779 280.613
R9738 GND.n5180 GND.n779 280.613
R9739 GND.n5181 GND.n5180 280.613
R9740 GND.n5182 GND.n5181 280.613
R9741 GND.n5182 GND.n773 280.613
R9742 GND.n5190 GND.n773 280.613
R9743 GND.n5191 GND.n5190 280.613
R9744 GND.n5192 GND.n5191 280.613
R9745 GND.n5192 GND.n767 280.613
R9746 GND.n5200 GND.n767 280.613
R9747 GND.n5201 GND.n5200 280.613
R9748 GND.n5202 GND.n5201 280.613
R9749 GND.n5202 GND.n761 280.613
R9750 GND.n5210 GND.n761 280.613
R9751 GND.n5211 GND.n5210 280.613
R9752 GND.n5212 GND.n5211 280.613
R9753 GND.n5212 GND.n755 280.613
R9754 GND.n5220 GND.n755 280.613
R9755 GND.n5221 GND.n5220 280.613
R9756 GND.n5222 GND.n5221 280.613
R9757 GND.n5222 GND.n749 280.613
R9758 GND.n5230 GND.n749 280.613
R9759 GND.n5231 GND.n5230 280.613
R9760 GND.n5232 GND.n5231 280.613
R9761 GND.n5232 GND.n743 280.613
R9762 GND.n5240 GND.n743 280.613
R9763 GND.n5241 GND.n5240 280.613
R9764 GND.n5242 GND.n5241 280.613
R9765 GND.n5242 GND.n737 280.613
R9766 GND.n5250 GND.n737 280.613
R9767 GND.n5251 GND.n5250 280.613
R9768 GND.n5252 GND.n5251 280.613
R9769 GND.n5252 GND.n731 280.613
R9770 GND.n5260 GND.n731 280.613
R9771 GND.n5261 GND.n5260 280.613
R9772 GND.n5262 GND.n5261 280.613
R9773 GND.n5262 GND.n725 280.613
R9774 GND.n5270 GND.n725 280.613
R9775 GND.n5271 GND.n5270 280.613
R9776 GND.n5272 GND.n5271 280.613
R9777 GND.n5272 GND.n719 280.613
R9778 GND.n5280 GND.n719 280.613
R9779 GND.n5281 GND.n5280 280.613
R9780 GND.n5282 GND.n5281 280.613
R9781 GND.n5282 GND.n713 280.613
R9782 GND.n5290 GND.n713 280.613
R9783 GND.n5291 GND.n5290 280.613
R9784 GND.n5292 GND.n5291 280.613
R9785 GND.n5292 GND.n707 280.613
R9786 GND.n5300 GND.n707 280.613
R9787 GND.n5301 GND.n5300 280.613
R9788 GND.n5302 GND.n5301 280.613
R9789 GND.n5302 GND.n701 280.613
R9790 GND.n5311 GND.n701 280.613
R9791 GND.n5312 GND.n5311 280.613
R9792 GND.n463 GND.t156 279.217
R9793 GND.n519 GND.t150 279.217
R9794 GND.n546 GND.t78 279.217
R9795 GND.n1286 GND.t144 279.217
R9796 GND.n1312 GND.t74 279.217
R9797 GND.n1372 GND.t135 279.217
R9798 GND.n2587 GND.t153 279.217
R9799 GND.n3625 GND.t82 279.217
R9800 GND.n3647 GND.t99 279.217
R9801 GND.n1131 GND.t102 279.217
R9802 GND.n1151 GND.t121 279.217
R9803 GND.n1810 GND.t138 279.217
R9804 GND.n2250 GND.t98 260.649
R9805 GND.n3505 GND.t117 260.649
R9806 GND.n3224 GND.n3223 256.663
R9807 GND.n3223 GND.n3036 256.663
R9808 GND.n3223 GND.n3037 256.663
R9809 GND.n3223 GND.n3038 256.663
R9810 GND.n3223 GND.n3039 256.663
R9811 GND.n3223 GND.n3040 256.663
R9812 GND.n3223 GND.n3041 256.663
R9813 GND.n3223 GND.n3042 256.663
R9814 GND.n3223 GND.n3043 256.663
R9815 GND.n3223 GND.n3044 256.663
R9816 GND.n3223 GND.n3045 256.663
R9817 GND.n3223 GND.n3046 256.663
R9818 GND.n3223 GND.n3047 256.663
R9819 GND.n3223 GND.n3048 256.663
R9820 GND.n3223 GND.n3049 256.663
R9821 GND.n3223 GND.n3050 256.663
R9822 GND.n3051 GND.n1290 256.663
R9823 GND.n3223 GND.n3052 256.663
R9824 GND.n3223 GND.n3053 256.663
R9825 GND.n3223 GND.n3054 256.663
R9826 GND.n3223 GND.n3055 256.663
R9827 GND.n3223 GND.n3056 256.663
R9828 GND.n3223 GND.n3057 256.663
R9829 GND.n3223 GND.n3058 256.663
R9830 GND.n3223 GND.n3059 256.663
R9831 GND.n3223 GND.n3060 256.663
R9832 GND.n3223 GND.n3061 256.663
R9833 GND.n3223 GND.n3062 256.663
R9834 GND.n3223 GND.n3063 256.663
R9835 GND.n3223 GND.n3064 256.663
R9836 GND.n3223 GND.n3065 256.663
R9837 GND.n3223 GND.n3066 256.663
R9838 GND.n3223 GND.n3067 256.663
R9839 GND.n3223 GND.n3159 256.663
R9840 GND.n3755 GND.n3475 256.663
R9841 GND.n3755 GND.n3476 256.663
R9842 GND.n3755 GND.n3477 256.663
R9843 GND.n3755 GND.n3478 256.663
R9844 GND.n3755 GND.n3479 256.663
R9845 GND.n3755 GND.n3480 256.663
R9846 GND.n3755 GND.n3481 256.663
R9847 GND.n3755 GND.n3482 256.663
R9848 GND.n3755 GND.n3483 256.663
R9849 GND.n3755 GND.n3484 256.663
R9850 GND.n3755 GND.n3485 256.663
R9851 GND.n3755 GND.n3486 256.663
R9852 GND.n3755 GND.n3487 256.663
R9853 GND.n3755 GND.n3488 256.663
R9854 GND.n3755 GND.n3489 256.663
R9855 GND.n3755 GND.n3490 256.663
R9856 GND.n3688 GND.n3491 256.663
R9857 GND.n3755 GND.n3474 256.663
R9858 GND.n3755 GND.n3473 256.663
R9859 GND.n3755 GND.n3472 256.663
R9860 GND.n3755 GND.n3471 256.663
R9861 GND.n3755 GND.n3470 256.663
R9862 GND.n3755 GND.n3469 256.663
R9863 GND.n3755 GND.n3468 256.663
R9864 GND.n3755 GND.n3467 256.663
R9865 GND.n3755 GND.n3466 256.663
R9866 GND.n3755 GND.n3465 256.663
R9867 GND.n3755 GND.n3464 256.663
R9868 GND.n3755 GND.n3463 256.663
R9869 GND.n3755 GND.n3462 256.663
R9870 GND.n3755 GND.n3461 256.663
R9871 GND.n3755 GND.n3460 256.663
R9872 GND.n3755 GND.n3459 256.663
R9873 GND.n3755 GND.n3458 256.663
R9874 GND.n4535 GND.n4534 242.672
R9875 GND.n4534 GND.n1326 242.672
R9876 GND.n4534 GND.n1327 242.672
R9877 GND.n4534 GND.n1328 242.672
R9878 GND.n4534 GND.n1329 242.672
R9879 GND.n4534 GND.n1330 242.672
R9880 GND.n4534 GND.n1331 242.672
R9881 GND.n4534 GND.n1332 242.672
R9882 GND.n4534 GND.n1333 242.672
R9883 GND.n4534 GND.n1334 242.672
R9884 GND.n4534 GND.n1335 242.672
R9885 GND.n4534 GND.n1336 242.672
R9886 GND.n4534 GND.n1337 242.672
R9887 GND.n4534 GND.n1338 242.672
R9888 GND.n4254 GND.n1762 242.672
R9889 GND.n4254 GND.n1763 242.672
R9890 GND.n4254 GND.n1764 242.672
R9891 GND.n4254 GND.n1765 242.672
R9892 GND.n4254 GND.n1766 242.672
R9893 GND.n4254 GND.n1767 242.672
R9894 GND.n4254 GND.n1768 242.672
R9895 GND.n4254 GND.n1769 242.672
R9896 GND.n4254 GND.n1770 242.672
R9897 GND.n4254 GND.n1771 242.672
R9898 GND.n4254 GND.n1772 242.672
R9899 GND.n4254 GND.n1773 242.672
R9900 GND.n4254 GND.n1774 242.672
R9901 GND.n4254 GND.n1775 242.672
R9902 GND.n4752 GND.n1102 242.672
R9903 GND.n4752 GND.n1103 242.672
R9904 GND.n4752 GND.n1104 242.672
R9905 GND.n4752 GND.n1105 242.672
R9906 GND.n4752 GND.n1106 242.672
R9907 GND.n4752 GND.n1107 242.672
R9908 GND.n4752 GND.n1108 242.672
R9909 GND.n4752 GND.n1109 242.672
R9910 GND.n4502 GND.n4501 242.672
R9911 GND.n4501 GND.n1390 242.672
R9912 GND.n4501 GND.n1388 242.672
R9913 GND.n4501 GND.n1386 242.672
R9914 GND.n4501 GND.n1385 242.672
R9915 GND.n4501 GND.n1383 242.672
R9916 GND.n4501 GND.n1379 242.672
R9917 GND.n4501 GND.n1377 242.672
R9918 GND.n4752 GND.n4751 242.672
R9919 GND.n4752 GND.n1086 242.672
R9920 GND.n4752 GND.n1087 242.672
R9921 GND.n4752 GND.n1088 242.672
R9922 GND.n4752 GND.n1089 242.672
R9923 GND.n4752 GND.n1090 242.672
R9924 GND.n4752 GND.n1091 242.672
R9925 GND.n4752 GND.n1092 242.672
R9926 GND.n4752 GND.n1093 242.672
R9927 GND.n4752 GND.n1094 242.672
R9928 GND.n4752 GND.n1095 242.672
R9929 GND.n4752 GND.n1096 242.672
R9930 GND.n4752 GND.n1097 242.672
R9931 GND.n4752 GND.n1098 242.672
R9932 GND.n4752 GND.n1099 242.672
R9933 GND.n4752 GND.n1100 242.672
R9934 GND.n4752 GND.n1101 242.672
R9935 GND.n4501 GND.n4477 242.672
R9936 GND.n4501 GND.n4478 242.672
R9937 GND.n4501 GND.n4480 242.672
R9938 GND.n4501 GND.n4481 242.672
R9939 GND.n4501 GND.n4483 242.672
R9940 GND.n4501 GND.n4484 242.672
R9941 GND.n4501 GND.n4486 242.672
R9942 GND.n4501 GND.n4487 242.672
R9943 GND.n4501 GND.n4489 242.672
R9944 GND.n4501 GND.n4490 242.672
R9945 GND.n4575 GND.n1289 242.672
R9946 GND.n4501 GND.n4491 242.672
R9947 GND.n4501 GND.n4493 242.672
R9948 GND.n4501 GND.n4494 242.672
R9949 GND.n4501 GND.n4496 242.672
R9950 GND.n4501 GND.n4497 242.672
R9951 GND.n4501 GND.n4499 242.672
R9952 GND.n4501 GND.n4500 242.672
R9953 GND.n4214 GND.n1823 242.672
R9954 GND.n4214 GND.n1824 242.672
R9955 GND.n4214 GND.n1825 242.672
R9956 GND.n4214 GND.n1826 242.672
R9957 GND.n4214 GND.n1827 242.672
R9958 GND.n4214 GND.n1828 242.672
R9959 GND.n4214 GND.n1829 242.672
R9960 GND.n3685 GND.n3580 242.672
R9961 GND.n4214 GND.n1831 242.672
R9962 GND.n4214 GND.n1832 242.672
R9963 GND.n4214 GND.n1833 242.672
R9964 GND.n4214 GND.n1834 242.672
R9965 GND.n4214 GND.n1835 242.672
R9966 GND.n4214 GND.n1836 242.672
R9967 GND.n4214 GND.n1837 242.672
R9968 GND.n4214 GND.n1838 242.672
R9969 GND.n4214 GND.n1839 242.672
R9970 GND.n4214 GND.n1840 242.672
R9971 GND.n5630 GND.n477 242.672
R9972 GND.n5630 GND.n478 242.672
R9973 GND.n5630 GND.n479 242.672
R9974 GND.n5630 GND.n480 242.672
R9975 GND.n5630 GND.n481 242.672
R9976 GND.n5630 GND.n482 242.672
R9977 GND.n5630 GND.n483 242.672
R9978 GND.n5630 GND.n484 242.672
R9979 GND.n5630 GND.n485 242.672
R9980 GND.n5630 GND.n486 242.672
R9981 GND.n5630 GND.n487 242.672
R9982 GND.n5630 GND.n488 242.672
R9983 GND.n5630 GND.n489 242.672
R9984 GND.n5630 GND.n490 242.672
R9985 GND.n5630 GND.n491 242.672
R9986 GND.n5630 GND.n492 242.672
R9987 GND.n5630 GND.n493 242.672
R9988 GND.n4214 GND.n1841 242.672
R9989 GND.n4214 GND.n1842 242.672
R9990 GND.n4214 GND.n1844 242.672
R9991 GND.n4214 GND.n1845 242.672
R9992 GND.n4214 GND.n1847 242.672
R9993 GND.n4214 GND.n1849 242.672
R9994 GND.n4214 GND.n1850 242.672
R9995 GND.n4215 GND.n4214 242.672
R9996 GND.n5630 GND.n475 242.672
R9997 GND.n5630 GND.n474 242.672
R9998 GND.n5630 GND.n473 242.672
R9999 GND.n5630 GND.n472 242.672
R10000 GND.n5630 GND.n471 242.672
R10001 GND.n5630 GND.n470 242.672
R10002 GND.n5630 GND.n469 242.672
R10003 GND.n5630 GND.n468 242.672
R10004 GND.n5629 GND.n495 240.244
R10005 GND.n500 GND.n499 240.244
R10006 GND.n502 GND.n501 240.244
R10007 GND.n506 GND.n505 240.244
R10008 GND.n508 GND.n507 240.244
R10009 GND.n512 GND.n511 240.244
R10010 GND.n514 GND.n513 240.244
R10011 GND.n518 GND.n517 240.244
R10012 GND.n522 GND.n521 240.244
R10013 GND.n526 GND.n525 240.244
R10014 GND.n528 GND.n527 240.244
R10015 GND.n532 GND.n531 240.244
R10016 GND.n534 GND.n533 240.244
R10017 GND.n538 GND.n537 240.244
R10018 GND.n540 GND.n539 240.244
R10019 GND.n544 GND.n543 240.244
R10020 GND.n548 GND.n545 240.244
R10021 GND.n1858 GND.n1857 240.244
R10022 GND.n1859 GND.n1858 240.244
R10023 GND.n3889 GND.n1859 240.244
R10024 GND.n3889 GND.n1865 240.244
R10025 GND.n1866 GND.n1865 240.244
R10026 GND.n1867 GND.n1866 240.244
R10027 GND.n2090 GND.n1867 240.244
R10028 GND.n2090 GND.n1873 240.244
R10029 GND.n1874 GND.n1873 240.244
R10030 GND.n1875 GND.n1874 240.244
R10031 GND.n2073 GND.n1875 240.244
R10032 GND.n2073 GND.n1881 240.244
R10033 GND.n1882 GND.n1881 240.244
R10034 GND.n1883 GND.n1882 240.244
R10035 GND.n2050 GND.n1883 240.244
R10036 GND.n2050 GND.n1889 240.244
R10037 GND.n1890 GND.n1889 240.244
R10038 GND.n1891 GND.n1890 240.244
R10039 GND.n2042 GND.n1891 240.244
R10040 GND.n2042 GND.n1897 240.244
R10041 GND.n1898 GND.n1897 240.244
R10042 GND.n1899 GND.n1898 240.244
R10043 GND.n2003 GND.n1899 240.244
R10044 GND.n2003 GND.n1905 240.244
R10045 GND.n1906 GND.n1905 240.244
R10046 GND.n1907 GND.n1906 240.244
R10047 GND.n4013 GND.n1907 240.244
R10048 GND.n4013 GND.n1913 240.244
R10049 GND.n1914 GND.n1913 240.244
R10050 GND.n1915 GND.n1914 240.244
R10051 GND.n1987 GND.n1915 240.244
R10052 GND.n1987 GND.n1921 240.244
R10053 GND.n1922 GND.n1921 240.244
R10054 GND.n1923 GND.n1922 240.244
R10055 GND.n1975 GND.n1923 240.244
R10056 GND.n1975 GND.n1929 240.244
R10057 GND.n1930 GND.n1929 240.244
R10058 GND.n1931 GND.n1930 240.244
R10059 GND.n4116 GND.n1931 240.244
R10060 GND.n4116 GND.n1937 240.244
R10061 GND.n1938 GND.n1937 240.244
R10062 GND.n1939 GND.n1938 240.244
R10063 GND.n1939 GND.n593 240.244
R10064 GND.n5488 GND.n593 240.244
R10065 GND.n5488 GND.n581 240.244
R10066 GND.n581 GND.n571 240.244
R10067 GND.n5504 GND.n571 240.244
R10068 GND.n5505 GND.n5504 240.244
R10069 GND.n5505 GND.n563 240.244
R10070 GND.n5507 GND.n563 240.244
R10071 GND.n5507 GND.n551 240.244
R10072 GND.n5573 GND.n551 240.244
R10073 GND.n3596 GND.n3595 240.244
R10074 GND.n3600 GND.n3599 240.244
R10075 GND.n3606 GND.n3605 240.244
R10076 GND.n3610 GND.n3609 240.244
R10077 GND.n3616 GND.n3615 240.244
R10078 GND.n3620 GND.n3619 240.244
R10079 GND.n3578 GND.n1830 240.244
R10080 GND.n3683 GND.n3682 240.244
R10081 GND.n3679 GND.n3678 240.244
R10082 GND.n3675 GND.n3674 240.244
R10083 GND.n3671 GND.n3670 240.244
R10084 GND.n3667 GND.n3666 240.244
R10085 GND.n3663 GND.n3662 240.244
R10086 GND.n3659 GND.n3658 240.244
R10087 GND.n3655 GND.n3654 240.244
R10088 GND.n3646 GND.n3643 240.244
R10089 GND.n3589 GND.n2111 240.244
R10090 GND.n3894 GND.n2111 240.244
R10091 GND.n3894 GND.n2105 240.244
R10092 GND.n3902 GND.n2105 240.244
R10093 GND.n3902 GND.n2107 240.244
R10094 GND.n2107 GND.n2088 240.244
R10095 GND.n3918 GND.n2088 240.244
R10096 GND.n3918 GND.n2083 240.244
R10097 GND.n3926 GND.n2083 240.244
R10098 GND.n3926 GND.n2084 240.244
R10099 GND.n2084 GND.n2067 240.244
R10100 GND.n3943 GND.n2067 240.244
R10101 GND.n3943 GND.n2062 240.244
R10102 GND.n3951 GND.n2062 240.244
R10103 GND.n3951 GND.n2063 240.244
R10104 GND.n2063 GND.n2034 240.244
R10105 GND.n3983 GND.n2034 240.244
R10106 GND.n3983 GND.n2035 240.244
R10107 GND.n2035 GND.n2029 240.244
R10108 GND.n3990 GND.n2029 240.244
R10109 GND.n3990 GND.n2030 240.244
R10110 GND.n2030 GND.n2000 240.244
R10111 GND.n4061 GND.n2000 240.244
R10112 GND.n4061 GND.n2001 240.244
R10113 GND.n4019 GND.n2001 240.244
R10114 GND.n4020 GND.n4019 240.244
R10115 GND.n4047 GND.n4020 240.244
R10116 GND.n4047 GND.n4044 240.244
R10117 GND.n4044 GND.n4021 240.244
R10118 GND.n4031 GND.n4021 240.244
R10119 GND.n4031 GND.n1991 240.244
R10120 GND.n4070 GND.n1991 240.244
R10121 GND.n4070 GND.n1992 240.244
R10122 GND.n1992 GND.n1973 240.244
R10123 GND.n4088 GND.n1973 240.244
R10124 GND.n4088 GND.n1968 240.244
R10125 GND.n4096 GND.n1968 240.244
R10126 GND.n4096 GND.n1969 240.244
R10127 GND.n1969 GND.n1950 240.244
R10128 GND.n4121 GND.n1950 240.244
R10129 GND.n4121 GND.n1945 240.244
R10130 GND.n4129 GND.n1945 240.244
R10131 GND.n4129 GND.n1946 240.244
R10132 GND.n1946 GND.n579 240.244
R10133 GND.n5496 GND.n579 240.244
R10134 GND.n5496 GND.n575 240.244
R10135 GND.n5502 GND.n575 240.244
R10136 GND.n5502 GND.n561 240.244
R10137 GND.n5514 GND.n561 240.244
R10138 GND.n5514 GND.n557 240.244
R10139 GND.n5521 GND.n557 240.244
R10140 GND.n5521 GND.n494 240.244
R10141 GND.n1270 GND.n1266 240.244
R10142 GND.n4498 GND.n1271 240.244
R10143 GND.n1275 GND.n1274 240.244
R10144 GND.n4495 GND.n1276 240.244
R10145 GND.n1280 GND.n1279 240.244
R10146 GND.n4492 GND.n1281 240.244
R10147 GND.n1285 GND.n1284 240.244
R10148 GND.n4488 GND.n1291 240.244
R10149 GND.n1295 GND.n1294 240.244
R10150 GND.n4485 GND.n1296 240.244
R10151 GND.n1300 GND.n1299 240.244
R10152 GND.n4482 GND.n1301 240.244
R10153 GND.n1305 GND.n1304 240.244
R10154 GND.n4479 GND.n1306 240.244
R10155 GND.n1310 GND.n1309 240.244
R10156 GND.n4476 GND.n1311 240.244
R10157 GND.n4681 GND.n1155 240.244
R10158 GND.n1161 GND.n1155 240.244
R10159 GND.n1162 GND.n1161 240.244
R10160 GND.n1163 GND.n1162 240.244
R10161 GND.n2496 GND.n1163 240.244
R10162 GND.n2496 GND.n1169 240.244
R10163 GND.n1170 GND.n1169 240.244
R10164 GND.n1171 GND.n1170 240.244
R10165 GND.n2482 GND.n1171 240.244
R10166 GND.n2482 GND.n1177 240.244
R10167 GND.n1178 GND.n1177 240.244
R10168 GND.n1179 GND.n1178 240.244
R10169 GND.n2665 GND.n1179 240.244
R10170 GND.n2665 GND.n1185 240.244
R10171 GND.n1186 GND.n1185 240.244
R10172 GND.n1187 GND.n1186 240.244
R10173 GND.n2447 GND.n1187 240.244
R10174 GND.n2447 GND.n1193 240.244
R10175 GND.n1194 GND.n1193 240.244
R10176 GND.n1195 GND.n1194 240.244
R10177 GND.n2426 GND.n1195 240.244
R10178 GND.n2426 GND.n1201 240.244
R10179 GND.n1202 GND.n1201 240.244
R10180 GND.n1203 GND.n1202 240.244
R10181 GND.n2395 GND.n1203 240.244
R10182 GND.n2395 GND.n1209 240.244
R10183 GND.n1210 GND.n1209 240.244
R10184 GND.n1211 GND.n1210 240.244
R10185 GND.n2419 GND.n1211 240.244
R10186 GND.n2419 GND.n1217 240.244
R10187 GND.n1218 GND.n1217 240.244
R10188 GND.n1219 GND.n1218 240.244
R10189 GND.n2366 GND.n1219 240.244
R10190 GND.n2366 GND.n1225 240.244
R10191 GND.n1226 GND.n1225 240.244
R10192 GND.n1227 GND.n1226 240.244
R10193 GND.n2785 GND.n1227 240.244
R10194 GND.n2785 GND.n1233 240.244
R10195 GND.n1234 GND.n1233 240.244
R10196 GND.n1235 GND.n1234 240.244
R10197 GND.n2334 GND.n1235 240.244
R10198 GND.n2334 GND.n1241 240.244
R10199 GND.n1242 GND.n1241 240.244
R10200 GND.n1243 GND.n1242 240.244
R10201 GND.n2315 GND.n1243 240.244
R10202 GND.n2315 GND.n1249 240.244
R10203 GND.n1250 GND.n1249 240.244
R10204 GND.n1251 GND.n1250 240.244
R10205 GND.n2307 GND.n1251 240.244
R10206 GND.n2307 GND.n1257 240.244
R10207 GND.n1258 GND.n1257 240.244
R10208 GND.n4601 GND.n1258 240.244
R10209 GND.n1113 GND.n1112 240.244
R10210 GND.n4745 GND.n1112 240.244
R10211 GND.n4743 GND.n4742 240.244
R10212 GND.n4739 GND.n4738 240.244
R10213 GND.n4735 GND.n4734 240.244
R10214 GND.n4731 GND.n4730 240.244
R10215 GND.n4727 GND.n4726 240.244
R10216 GND.n4723 GND.n4722 240.244
R10217 GND.n4718 GND.n4717 240.244
R10218 GND.n4714 GND.n4713 240.244
R10219 GND.n4710 GND.n4709 240.244
R10220 GND.n4706 GND.n4705 240.244
R10221 GND.n4702 GND.n4701 240.244
R10222 GND.n4698 GND.n4697 240.244
R10223 GND.n4694 GND.n4693 240.244
R10224 GND.n4690 GND.n4689 240.244
R10225 GND.n1150 GND.n1149 240.244
R10226 GND.n2551 GND.n1114 240.244
R10227 GND.n2620 GND.n2551 240.244
R10228 GND.n2620 GND.n2544 240.244
R10229 GND.n2628 GND.n2544 240.244
R10230 GND.n2628 GND.n2545 240.244
R10231 GND.n2545 GND.n2491 240.244
R10232 GND.n2645 GND.n2491 240.244
R10233 GND.n2645 GND.n2485 240.244
R10234 GND.n2653 GND.n2485 240.244
R10235 GND.n2653 GND.n2487 240.244
R10236 GND.n2487 GND.n2468 240.244
R10237 GND.n2670 GND.n2468 240.244
R10238 GND.n2670 GND.n2462 240.244
R10239 GND.n2678 GND.n2462 240.244
R10240 GND.n2678 GND.n2464 240.244
R10241 GND.n2464 GND.n2445 240.244
R10242 GND.n2707 GND.n2445 240.244
R10243 GND.n2707 GND.n2439 240.244
R10244 GND.n2714 GND.n2439 240.244
R10245 GND.n2714 GND.n2441 240.244
R10246 GND.n2441 GND.n2440 240.244
R10247 GND.n2440 GND.n2387 240.244
R10248 GND.n2827 GND.n2387 240.244
R10249 GND.n2827 GND.n2388 240.244
R10250 GND.n2411 GND.n2388 240.244
R10251 GND.n2412 GND.n2411 240.244
R10252 GND.n2812 GND.n2412 240.244
R10253 GND.n2812 GND.n2809 240.244
R10254 GND.n2809 GND.n2413 240.244
R10255 GND.n2413 GND.n2377 240.244
R10256 GND.n2835 GND.n2377 240.244
R10257 GND.n2835 GND.n2378 240.244
R10258 GND.n2378 GND.n2361 240.244
R10259 GND.n2852 GND.n2361 240.244
R10260 GND.n2852 GND.n2356 240.244
R10261 GND.n2860 GND.n2356 240.244
R10262 GND.n2860 GND.n2357 240.244
R10263 GND.n2357 GND.n2342 240.244
R10264 GND.n2877 GND.n2342 240.244
R10265 GND.n2877 GND.n2337 240.244
R10266 GND.n2885 GND.n2337 240.244
R10267 GND.n2885 GND.n2338 240.244
R10268 GND.n2338 GND.n2321 240.244
R10269 GND.n2903 GND.n2321 240.244
R10270 GND.n2903 GND.n2317 240.244
R10271 GND.n2909 GND.n2317 240.244
R10272 GND.n2909 GND.n2295 240.244
R10273 GND.n2943 GND.n2295 240.244
R10274 GND.n2943 GND.n2291 240.244
R10275 GND.n2949 GND.n2291 240.244
R10276 GND.n2949 GND.n1265 240.244
R10277 GND.n4599 GND.n1265 240.244
R10278 GND.n1317 GND.n1316 240.244
R10279 GND.n1378 GND.n1318 240.244
R10280 GND.n1382 GND.n1381 240.244
R10281 GND.n1347 GND.n1346 240.244
R10282 GND.n1384 GND.n1354 240.244
R10283 GND.n1387 GND.n1355 240.244
R10284 GND.n1365 GND.n1364 240.244
R10285 GND.n1389 GND.n1374 240.244
R10286 GND.n2578 GND.n2577 240.244
R10287 GND.n2578 GND.n2553 240.244
R10288 GND.n2553 GND.n2503 240.244
R10289 GND.n2630 GND.n2503 240.244
R10290 GND.n2630 GND.n2498 240.244
R10291 GND.n2637 GND.n2498 240.244
R10292 GND.n2637 GND.n2493 240.244
R10293 GND.n2493 GND.n2480 240.244
R10294 GND.n2655 GND.n2480 240.244
R10295 GND.n2655 GND.n2475 240.244
R10296 GND.n2662 GND.n2475 240.244
R10297 GND.n2662 GND.n2470 240.244
R10298 GND.n2470 GND.n2458 240.244
R10299 GND.n2680 GND.n2458 240.244
R10300 GND.n2680 GND.n2453 240.244
R10301 GND.n2701 GND.n2453 240.244
R10302 GND.n2701 GND.n2448 240.244
R10303 GND.n2685 GND.n2448 240.244
R10304 GND.n2685 GND.n2436 240.244
R10305 GND.n2691 GND.n2436 240.244
R10306 GND.n2691 GND.n2425 240.244
R10307 GND.n2730 GND.n2425 240.244
R10308 GND.n2730 GND.n2390 240.244
R10309 GND.n2394 GND.n2390 240.244
R10310 GND.n2737 GND.n2394 240.244
R10311 GND.n2738 GND.n2737 240.244
R10312 GND.n2738 GND.n2404 240.244
R10313 GND.n2416 GND.n2404 240.244
R10314 GND.n2745 GND.n2416 240.244
R10315 GND.n2745 GND.n2372 240.244
R10316 GND.n2837 GND.n2372 240.244
R10317 GND.n2837 GND.n2367 240.244
R10318 GND.n2844 GND.n2367 240.244
R10319 GND.n2844 GND.n2363 240.244
R10320 GND.n2363 GND.n2352 240.244
R10321 GND.n2862 GND.n2352 240.244
R10322 GND.n2862 GND.n2347 240.244
R10323 GND.n2869 GND.n2347 240.244
R10324 GND.n2869 GND.n2344 240.244
R10325 GND.n2344 GND.n2332 240.244
R10326 GND.n2887 GND.n2332 240.244
R10327 GND.n2887 GND.n2327 240.244
R10328 GND.n2897 GND.n2327 240.244
R10329 GND.n2897 GND.n2323 240.244
R10330 GND.n2891 GND.n2323 240.244
R10331 GND.n2891 GND.n2302 240.244
R10332 GND.n2938 GND.n2302 240.244
R10333 GND.n2938 GND.n2297 240.244
R10334 GND.n2932 GND.n2297 240.244
R10335 GND.n2932 GND.n2288 240.244
R10336 GND.n2956 GND.n2288 240.244
R10337 GND.n2956 GND.n1262 240.244
R10338 GND.n2556 GND.n2555 240.244
R10339 GND.n2560 GND.n2559 240.244
R10340 GND.n2562 GND.n2561 240.244
R10341 GND.n2566 GND.n2565 240.244
R10342 GND.n2568 GND.n2567 240.244
R10343 GND.n2572 GND.n2571 240.244
R10344 GND.n2574 GND.n2573 240.244
R10345 GND.n2586 GND.n1110 240.244
R10346 GND.n2615 GND.n2614 240.244
R10347 GND.n2618 GND.n2615 240.244
R10348 GND.n2618 GND.n2617 240.244
R10349 GND.n2617 GND.n2543 240.244
R10350 GND.n2543 GND.n2495 240.244
R10351 GND.n2639 GND.n2495 240.244
R10352 GND.n2643 GND.n2639 240.244
R10353 GND.n2643 GND.n2641 240.244
R10354 GND.n2641 GND.n2484 240.244
R10355 GND.n2484 GND.n2472 240.244
R10356 GND.n2664 GND.n2472 240.244
R10357 GND.n2668 GND.n2664 240.244
R10358 GND.n2668 GND.n2667 240.244
R10359 GND.n2667 GND.n2461 240.244
R10360 GND.n2461 GND.n2451 240.244
R10361 GND.n2703 GND.n2451 240.244
R10362 GND.n2705 GND.n2703 240.244
R10363 GND.n2705 GND.n2704 240.244
R10364 GND.n2704 GND.n2438 240.244
R10365 GND.n2689 GND.n2438 240.244
R10366 GND.n2689 GND.n2688 240.244
R10367 GND.n2688 GND.n2392 240.244
R10368 GND.n2825 GND.n2392 240.244
R10369 GND.n2825 GND.n2823 240.244
R10370 GND.n2823 GND.n2393 240.244
R10371 GND.n2406 GND.n2393 240.244
R10372 GND.n2408 GND.n2406 240.244
R10373 GND.n2807 GND.n2408 240.244
R10374 GND.n2807 GND.n2806 240.244
R10375 GND.n2806 GND.n2418 240.244
R10376 GND.n2418 GND.n2376 240.244
R10377 GND.n2376 GND.n2365 240.244
R10378 GND.n2846 GND.n2365 240.244
R10379 GND.n2850 GND.n2846 240.244
R10380 GND.n2850 GND.n2849 240.244
R10381 GND.n2849 GND.n2355 240.244
R10382 GND.n2355 GND.n2346 240.244
R10383 GND.n2871 GND.n2346 240.244
R10384 GND.n2875 GND.n2871 240.244
R10385 GND.n2875 GND.n2873 240.244
R10386 GND.n2873 GND.n2336 240.244
R10387 GND.n2336 GND.n2325 240.244
R10388 GND.n2899 GND.n2325 240.244
R10389 GND.n2901 GND.n2899 240.244
R10390 GND.n2901 GND.n2900 240.244
R10391 GND.n2900 GND.n2299 240.244
R10392 GND.n2940 GND.n2299 240.244
R10393 GND.n2941 GND.n2940 240.244
R10394 GND.n2941 GND.n2290 240.244
R10395 GND.n2951 GND.n2290 240.244
R10396 GND.n2954 GND.n2951 240.244
R10397 GND.n2954 GND.n1264 240.244
R10398 GND.n4253 GND.n1777 240.244
R10399 GND.n1787 GND.n1786 240.244
R10400 GND.n1795 GND.n1794 240.244
R10401 GND.n1797 GND.n1796 240.244
R10402 GND.n1805 GND.n1804 240.244
R10403 GND.n1815 GND.n1814 240.244
R10404 GND.n1817 GND.n1816 240.244
R10405 GND.n2144 GND.n2143 240.244
R10406 GND.n2146 GND.n2145 240.244
R10407 GND.n2150 GND.n2149 240.244
R10408 GND.n2152 GND.n2151 240.244
R10409 GND.n2156 GND.n2155 240.244
R10410 GND.n2160 GND.n2157 240.244
R10411 GND.n2164 GND.n2163 240.244
R10412 GND.n1402 GND.n1401 240.244
R10413 GND.n3006 GND.n1402 240.244
R10414 GND.n3006 GND.n1413 240.244
R10415 GND.n3012 GND.n1413 240.244
R10416 GND.n3013 GND.n3012 240.244
R10417 GND.n3013 GND.n1433 240.244
R10418 GND.n2270 GND.n1433 240.244
R10419 GND.n2270 GND.n1446 240.244
R10420 GND.n3021 GND.n1446 240.244
R10421 GND.n3022 GND.n3021 240.244
R10422 GND.n3022 GND.n1460 240.244
R10423 GND.n3034 GND.n1460 240.244
R10424 GND.n3034 GND.n1473 240.244
R10425 GND.n3027 GND.n1473 240.244
R10426 GND.n3027 GND.n2239 240.244
R10427 GND.n3248 GND.n2239 240.244
R10428 GND.n3249 GND.n3248 240.244
R10429 GND.n3249 GND.n2233 240.244
R10430 GND.n3271 GND.n2233 240.244
R10431 GND.n3271 GND.n2234 240.244
R10432 GND.n3254 GND.n2234 240.244
R10433 GND.n3257 GND.n3254 240.244
R10434 GND.n3257 GND.n2221 240.244
R10435 GND.n2221 GND.n1522 240.244
R10436 GND.n3259 GND.n1522 240.244
R10437 GND.n3259 GND.n2215 240.244
R10438 GND.n3321 GND.n2215 240.244
R10439 GND.n3321 GND.n1540 240.244
R10440 GND.n3348 GND.n1540 240.244
R10441 GND.n3348 GND.n1551 240.244
R10442 GND.n3326 GND.n1551 240.244
R10443 GND.n3327 GND.n3326 240.244
R10444 GND.n3328 GND.n3327 240.244
R10445 GND.n3329 GND.n3328 240.244
R10446 GND.n3329 GND.n1585 240.244
R10447 GND.n3332 GND.n1585 240.244
R10448 GND.n3332 GND.n1604 240.244
R10449 GND.n3395 GND.n1604 240.244
R10450 GND.n3396 GND.n3395 240.244
R10451 GND.n3397 GND.n3396 240.244
R10452 GND.n3397 GND.n1628 240.244
R10453 GND.n3407 GND.n1628 240.244
R10454 GND.n3407 GND.n1643 240.244
R10455 GND.n3401 GND.n1643 240.244
R10456 GND.n3401 GND.n2185 240.244
R10457 GND.n3442 GND.n2185 240.244
R10458 GND.n3442 GND.n1663 240.244
R10459 GND.n3449 GND.n1663 240.244
R10460 GND.n3449 GND.n1679 240.244
R10461 GND.n3781 GND.n1679 240.244
R10462 GND.n3781 GND.n1688 240.244
R10463 GND.n3457 GND.n1688 240.244
R10464 GND.n3457 GND.n1696 240.244
R10465 GND.n3789 GND.n1696 240.244
R10466 GND.n3790 GND.n3789 240.244
R10467 GND.n3790 GND.n1708 240.244
R10468 GND.n2172 GND.n1708 240.244
R10469 GND.n2172 GND.n1721 240.244
R10470 GND.n3798 GND.n1721 240.244
R10471 GND.n3798 GND.n3797 240.244
R10472 GND.n3797 GND.n1735 240.244
R10473 GND.n3806 GND.n1735 240.244
R10474 GND.n3806 GND.n1747 240.244
R10475 GND.n2165 GND.n1747 240.244
R10476 GND.n3813 GND.n2165 240.244
R10477 GND.n4533 GND.n1324 240.244
R10478 GND.n4533 GND.n1340 240.244
R10479 GND.n1351 GND.n1350 240.244
R10480 GND.n1359 GND.n1358 240.244
R10481 GND.n1361 GND.n1360 240.244
R10482 GND.n1369 GND.n1368 240.244
R10483 GND.n2283 GND.n2282 240.244
R10484 GND.n2964 GND.n2963 240.244
R10485 GND.n2967 GND.n2966 240.244
R10486 GND.n2974 GND.n2973 240.244
R10487 GND.n2977 GND.n2976 240.244
R10488 GND.n2984 GND.n2983 240.244
R10489 GND.n2987 GND.n2986 240.244
R10490 GND.n2997 GND.n2996 240.244
R10491 GND.n4463 GND.n1323 240.244
R10492 GND.n4463 GND.n1404 240.244
R10493 GND.n4459 GND.n1404 240.244
R10494 GND.n4459 GND.n1411 240.244
R10495 GND.n1435 GND.n1411 240.244
R10496 GND.n4449 GND.n1435 240.244
R10497 GND.n4449 GND.n1436 240.244
R10498 GND.n4445 GND.n1436 240.244
R10499 GND.n4445 GND.n1444 240.244
R10500 GND.n1462 GND.n1444 240.244
R10501 GND.n4435 GND.n1462 240.244
R10502 GND.n4435 GND.n1463 240.244
R10503 GND.n4431 GND.n1463 240.244
R10504 GND.n4431 GND.n1471 240.244
R10505 GND.n3234 GND.n1471 240.244
R10506 GND.n3246 GND.n3234 240.244
R10507 GND.n3246 GND.n3235 240.244
R10508 GND.n3235 GND.n2226 240.244
R10509 GND.n3273 GND.n2226 240.244
R10510 GND.n3274 GND.n3273 240.244
R10511 GND.n3275 GND.n3274 240.244
R10512 GND.n3275 GND.n2222 240.244
R10513 GND.n3290 GND.n2222 240.244
R10514 GND.n3290 GND.n1524 240.244
R10515 GND.n3286 GND.n1524 240.244
R10516 GND.n3286 GND.n3285 240.244
R10517 GND.n3285 GND.n1542 240.244
R10518 GND.n4379 GND.n1542 240.244
R10519 GND.n4379 GND.n1543 240.244
R10520 GND.n4375 GND.n1543 240.244
R10521 GND.n4375 GND.n1549 240.244
R10522 GND.n1593 GND.n1549 240.244
R10523 GND.n1594 GND.n1593 240.244
R10524 GND.n1594 GND.n1587 240.244
R10525 GND.n4351 GND.n1587 240.244
R10526 GND.n4351 GND.n1588 240.244
R10527 GND.n4347 GND.n1588 240.244
R10528 GND.n4347 GND.n1602 240.244
R10529 GND.n1634 GND.n1602 240.244
R10530 GND.n1634 GND.n1630 240.244
R10531 GND.n4331 GND.n1630 240.244
R10532 GND.n4331 GND.n1631 240.244
R10533 GND.n4327 GND.n1631 240.244
R10534 GND.n4327 GND.n1642 240.244
R10535 GND.n1669 GND.n1642 240.244
R10536 GND.n1669 GND.n1665 240.244
R10537 GND.n4310 GND.n1665 240.244
R10538 GND.n4310 GND.n1666 240.244
R10539 GND.n4306 GND.n1666 240.244
R10540 GND.n4306 GND.n1677 240.244
R10541 GND.n4296 GND.n1677 240.244
R10542 GND.n4296 GND.n1689 240.244
R10543 GND.n4292 GND.n1689 240.244
R10544 GND.n4292 GND.n1695 240.244
R10545 GND.n1710 GND.n1695 240.244
R10546 GND.n4282 GND.n1710 240.244
R10547 GND.n4282 GND.n1711 240.244
R10548 GND.n4278 GND.n1711 240.244
R10549 GND.n4278 GND.n1719 240.244
R10550 GND.n1737 GND.n1719 240.244
R10551 GND.n4268 GND.n1737 240.244
R10552 GND.n4268 GND.n1738 240.244
R10553 GND.n4264 GND.n1738 240.244
R10554 GND.n4264 GND.n1746 240.244
R10555 GND.n1776 GND.n1746 240.244
R10556 GND.n4889 GND.n954 240.244
R10557 GND.n4889 GND.n952 240.244
R10558 GND.n4893 GND.n952 240.244
R10559 GND.n4893 GND.n948 240.244
R10560 GND.n4899 GND.n948 240.244
R10561 GND.n4899 GND.n946 240.244
R10562 GND.n4903 GND.n946 240.244
R10563 GND.n4903 GND.n942 240.244
R10564 GND.n4909 GND.n942 240.244
R10565 GND.n4909 GND.n940 240.244
R10566 GND.n4913 GND.n940 240.244
R10567 GND.n4913 GND.n936 240.244
R10568 GND.n4919 GND.n936 240.244
R10569 GND.n4919 GND.n934 240.244
R10570 GND.n4923 GND.n934 240.244
R10571 GND.n4923 GND.n930 240.244
R10572 GND.n4929 GND.n930 240.244
R10573 GND.n4929 GND.n928 240.244
R10574 GND.n4933 GND.n928 240.244
R10575 GND.n4933 GND.n924 240.244
R10576 GND.n4939 GND.n924 240.244
R10577 GND.n4939 GND.n922 240.244
R10578 GND.n4943 GND.n922 240.244
R10579 GND.n4943 GND.n918 240.244
R10580 GND.n4949 GND.n918 240.244
R10581 GND.n4949 GND.n916 240.244
R10582 GND.n4953 GND.n916 240.244
R10583 GND.n4953 GND.n912 240.244
R10584 GND.n4959 GND.n912 240.244
R10585 GND.n4959 GND.n910 240.244
R10586 GND.n4963 GND.n910 240.244
R10587 GND.n4963 GND.n906 240.244
R10588 GND.n4969 GND.n906 240.244
R10589 GND.n4969 GND.n904 240.244
R10590 GND.n4973 GND.n904 240.244
R10591 GND.n4973 GND.n900 240.244
R10592 GND.n4979 GND.n900 240.244
R10593 GND.n4979 GND.n898 240.244
R10594 GND.n4983 GND.n898 240.244
R10595 GND.n4983 GND.n894 240.244
R10596 GND.n4989 GND.n894 240.244
R10597 GND.n4989 GND.n892 240.244
R10598 GND.n4993 GND.n892 240.244
R10599 GND.n4993 GND.n888 240.244
R10600 GND.n4999 GND.n888 240.244
R10601 GND.n4999 GND.n886 240.244
R10602 GND.n5003 GND.n886 240.244
R10603 GND.n5003 GND.n882 240.244
R10604 GND.n5009 GND.n882 240.244
R10605 GND.n5009 GND.n880 240.244
R10606 GND.n5013 GND.n880 240.244
R10607 GND.n5013 GND.n876 240.244
R10608 GND.n5019 GND.n876 240.244
R10609 GND.n5019 GND.n874 240.244
R10610 GND.n5023 GND.n874 240.244
R10611 GND.n5023 GND.n870 240.244
R10612 GND.n5029 GND.n870 240.244
R10613 GND.n5029 GND.n868 240.244
R10614 GND.n5033 GND.n868 240.244
R10615 GND.n5033 GND.n864 240.244
R10616 GND.n5039 GND.n864 240.244
R10617 GND.n5039 GND.n862 240.244
R10618 GND.n5043 GND.n862 240.244
R10619 GND.n5043 GND.n858 240.244
R10620 GND.n5049 GND.n858 240.244
R10621 GND.n5049 GND.n856 240.244
R10622 GND.n5053 GND.n856 240.244
R10623 GND.n5053 GND.n852 240.244
R10624 GND.n5059 GND.n852 240.244
R10625 GND.n5059 GND.n850 240.244
R10626 GND.n5063 GND.n850 240.244
R10627 GND.n5063 GND.n846 240.244
R10628 GND.n5069 GND.n846 240.244
R10629 GND.n5069 GND.n844 240.244
R10630 GND.n5073 GND.n844 240.244
R10631 GND.n5073 GND.n840 240.244
R10632 GND.n5079 GND.n840 240.244
R10633 GND.n5079 GND.n838 240.244
R10634 GND.n5083 GND.n838 240.244
R10635 GND.n5083 GND.n834 240.244
R10636 GND.n5089 GND.n834 240.244
R10637 GND.n5089 GND.n832 240.244
R10638 GND.n5093 GND.n832 240.244
R10639 GND.n5093 GND.n828 240.244
R10640 GND.n5099 GND.n828 240.244
R10641 GND.n5099 GND.n826 240.244
R10642 GND.n5103 GND.n826 240.244
R10643 GND.n5103 GND.n822 240.244
R10644 GND.n5109 GND.n822 240.244
R10645 GND.n5109 GND.n820 240.244
R10646 GND.n5113 GND.n820 240.244
R10647 GND.n5113 GND.n816 240.244
R10648 GND.n5119 GND.n816 240.244
R10649 GND.n5119 GND.n814 240.244
R10650 GND.n5123 GND.n814 240.244
R10651 GND.n5123 GND.n810 240.244
R10652 GND.n5129 GND.n810 240.244
R10653 GND.n5129 GND.n808 240.244
R10654 GND.n5133 GND.n808 240.244
R10655 GND.n5133 GND.n804 240.244
R10656 GND.n5139 GND.n804 240.244
R10657 GND.n5139 GND.n802 240.244
R10658 GND.n5143 GND.n802 240.244
R10659 GND.n5143 GND.n798 240.244
R10660 GND.n5149 GND.n798 240.244
R10661 GND.n5149 GND.n796 240.244
R10662 GND.n5153 GND.n796 240.244
R10663 GND.n5153 GND.n792 240.244
R10664 GND.n5159 GND.n792 240.244
R10665 GND.n5159 GND.n790 240.244
R10666 GND.n5163 GND.n790 240.244
R10667 GND.n5163 GND.n786 240.244
R10668 GND.n5169 GND.n786 240.244
R10669 GND.n5169 GND.n784 240.244
R10670 GND.n5173 GND.n784 240.244
R10671 GND.n5173 GND.n780 240.244
R10672 GND.n5179 GND.n780 240.244
R10673 GND.n5179 GND.n778 240.244
R10674 GND.n5183 GND.n778 240.244
R10675 GND.n5183 GND.n774 240.244
R10676 GND.n5189 GND.n774 240.244
R10677 GND.n5189 GND.n772 240.244
R10678 GND.n5193 GND.n772 240.244
R10679 GND.n5193 GND.n768 240.244
R10680 GND.n5199 GND.n768 240.244
R10681 GND.n5199 GND.n766 240.244
R10682 GND.n5203 GND.n766 240.244
R10683 GND.n5203 GND.n762 240.244
R10684 GND.n5209 GND.n762 240.244
R10685 GND.n5209 GND.n760 240.244
R10686 GND.n5213 GND.n760 240.244
R10687 GND.n5213 GND.n756 240.244
R10688 GND.n5219 GND.n756 240.244
R10689 GND.n5219 GND.n754 240.244
R10690 GND.n5223 GND.n754 240.244
R10691 GND.n5223 GND.n750 240.244
R10692 GND.n5229 GND.n750 240.244
R10693 GND.n5229 GND.n748 240.244
R10694 GND.n5233 GND.n748 240.244
R10695 GND.n5233 GND.n744 240.244
R10696 GND.n5239 GND.n744 240.244
R10697 GND.n5239 GND.n742 240.244
R10698 GND.n5243 GND.n742 240.244
R10699 GND.n5243 GND.n738 240.244
R10700 GND.n5249 GND.n738 240.244
R10701 GND.n5249 GND.n736 240.244
R10702 GND.n5253 GND.n736 240.244
R10703 GND.n5253 GND.n732 240.244
R10704 GND.n5259 GND.n732 240.244
R10705 GND.n5259 GND.n730 240.244
R10706 GND.n5263 GND.n730 240.244
R10707 GND.n5263 GND.n726 240.244
R10708 GND.n5269 GND.n726 240.244
R10709 GND.n5269 GND.n724 240.244
R10710 GND.n5273 GND.n724 240.244
R10711 GND.n5273 GND.n720 240.244
R10712 GND.n5279 GND.n720 240.244
R10713 GND.n5279 GND.n718 240.244
R10714 GND.n5283 GND.n718 240.244
R10715 GND.n5283 GND.n714 240.244
R10716 GND.n5289 GND.n714 240.244
R10717 GND.n5289 GND.n712 240.244
R10718 GND.n5293 GND.n712 240.244
R10719 GND.n5293 GND.n708 240.244
R10720 GND.n5299 GND.n708 240.244
R10721 GND.n5299 GND.n706 240.244
R10722 GND.n5303 GND.n706 240.244
R10723 GND.n5303 GND.n702 240.244
R10724 GND.n5310 GND.n702 240.244
R10725 GND.n5310 GND.n700 240.244
R10726 GND.n5314 GND.n697 240.244
R10727 GND.n5320 GND.n697 240.244
R10728 GND.n5320 GND.n695 240.244
R10729 GND.n5324 GND.n695 240.244
R10730 GND.n5324 GND.n691 240.244
R10731 GND.n5330 GND.n691 240.244
R10732 GND.n5330 GND.n689 240.244
R10733 GND.n5334 GND.n689 240.244
R10734 GND.n5334 GND.n685 240.244
R10735 GND.n5340 GND.n685 240.244
R10736 GND.n5340 GND.n683 240.244
R10737 GND.n5344 GND.n683 240.244
R10738 GND.n5344 GND.n679 240.244
R10739 GND.n5350 GND.n679 240.244
R10740 GND.n5350 GND.n677 240.244
R10741 GND.n5354 GND.n677 240.244
R10742 GND.n5354 GND.n673 240.244
R10743 GND.n5360 GND.n673 240.244
R10744 GND.n5360 GND.n671 240.244
R10745 GND.n5364 GND.n671 240.244
R10746 GND.n5364 GND.n667 240.244
R10747 GND.n5370 GND.n667 240.244
R10748 GND.n5370 GND.n665 240.244
R10749 GND.n5374 GND.n665 240.244
R10750 GND.n5374 GND.n661 240.244
R10751 GND.n5380 GND.n661 240.244
R10752 GND.n5380 GND.n659 240.244
R10753 GND.n5384 GND.n659 240.244
R10754 GND.n5384 GND.n655 240.244
R10755 GND.n5390 GND.n655 240.244
R10756 GND.n5390 GND.n653 240.244
R10757 GND.n5394 GND.n653 240.244
R10758 GND.n5394 GND.n649 240.244
R10759 GND.n5400 GND.n649 240.244
R10760 GND.n5400 GND.n647 240.244
R10761 GND.n5404 GND.n647 240.244
R10762 GND.n5404 GND.n643 240.244
R10763 GND.n5410 GND.n643 240.244
R10764 GND.n5410 GND.n641 240.244
R10765 GND.n5414 GND.n641 240.244
R10766 GND.n5414 GND.n637 240.244
R10767 GND.n5420 GND.n637 240.244
R10768 GND.n5420 GND.n635 240.244
R10769 GND.n5424 GND.n635 240.244
R10770 GND.n5424 GND.n631 240.244
R10771 GND.n5430 GND.n631 240.244
R10772 GND.n5430 GND.n629 240.244
R10773 GND.n5434 GND.n629 240.244
R10774 GND.n5434 GND.n625 240.244
R10775 GND.n5440 GND.n625 240.244
R10776 GND.n5440 GND.n623 240.244
R10777 GND.n5444 GND.n623 240.244
R10778 GND.n5444 GND.n619 240.244
R10779 GND.n5450 GND.n619 240.244
R10780 GND.n5450 GND.n617 240.244
R10781 GND.n5454 GND.n617 240.244
R10782 GND.n5454 GND.n613 240.244
R10783 GND.n5460 GND.n613 240.244
R10784 GND.n5460 GND.n611 240.244
R10785 GND.n5464 GND.n611 240.244
R10786 GND.n5464 GND.n607 240.244
R10787 GND.n5470 GND.n607 240.244
R10788 GND.n5470 GND.n605 240.244
R10789 GND.n5474 GND.n605 240.244
R10790 GND.n5474 GND.n601 240.244
R10791 GND.n5480 GND.n601 240.244
R10792 GND.n2535 GND.n2505 240.244
R10793 GND.n2535 GND.n2534 240.244
R10794 GND.n2534 GND.n2533 240.244
R10795 GND.n2533 GND.n2509 240.244
R10796 GND.n2529 GND.n2509 240.244
R10797 GND.n2529 GND.n2528 240.244
R10798 GND.n2528 GND.n2527 240.244
R10799 GND.n2527 GND.n2515 240.244
R10800 GND.n2523 GND.n2515 240.244
R10801 GND.n2523 GND.n2522 240.244
R10802 GND.n2522 GND.n2433 240.244
R10803 GND.n2717 GND.n2433 240.244
R10804 GND.n2717 GND.n2434 240.244
R10805 GND.n2434 GND.n2428 240.244
R10806 GND.n2727 GND.n2428 240.244
R10807 GND.n2727 GND.n2429 240.244
R10808 GND.n2429 GND.n2397 240.244
R10809 GND.n2820 GND.n2397 240.244
R10810 GND.n2820 GND.n2398 240.244
R10811 GND.n2815 GND.n2398 240.244
R10812 GND.n2815 GND.n2401 240.244
R10813 GND.n2747 GND.n2401 240.244
R10814 GND.n2803 GND.n2747 240.244
R10815 GND.n2803 GND.n2748 240.244
R10816 GND.n2798 GND.n2748 240.244
R10817 GND.n2798 GND.n2797 240.244
R10818 GND.n2797 GND.n2794 240.244
R10819 GND.n2794 GND.n2753 240.244
R10820 GND.n2790 GND.n2753 240.244
R10821 GND.n2790 GND.n2789 240.244
R10822 GND.n2789 GND.n2788 240.244
R10823 GND.n2788 GND.n2759 240.244
R10824 GND.n2781 GND.n2759 240.244
R10825 GND.n2781 GND.n2780 240.244
R10826 GND.n2780 GND.n2779 240.244
R10827 GND.n2779 GND.n2767 240.244
R10828 GND.n2775 GND.n2767 240.244
R10829 GND.n2775 GND.n2313 240.244
R10830 GND.n2912 GND.n2313 240.244
R10831 GND.n2913 GND.n2912 240.244
R10832 GND.n2914 GND.n2913 240.244
R10833 GND.n2914 GND.n2308 240.244
R10834 GND.n2929 GND.n2308 240.244
R10835 GND.n2929 GND.n2309 240.244
R10836 GND.n2925 GND.n2309 240.244
R10837 GND.n2925 GND.n2924 240.244
R10838 GND.n2924 GND.n1392 240.244
R10839 GND.n4474 GND.n1392 240.244
R10840 GND.n4474 GND.n1393 240.244
R10841 GND.n4470 GND.n1393 240.244
R10842 GND.n4470 GND.n4469 240.244
R10843 GND.n4469 GND.n4468 240.244
R10844 GND.n4468 GND.n1399 240.244
R10845 GND.n1422 GND.n1399 240.244
R10846 GND.n1422 GND.n1415 240.244
R10847 GND.n4456 GND.n1415 240.244
R10848 GND.n4456 GND.n1416 240.244
R10849 GND.n4452 GND.n1416 240.244
R10850 GND.n4452 GND.n1430 240.244
R10851 GND.n1448 GND.n1430 240.244
R10852 GND.n4442 GND.n1448 240.244
R10853 GND.n4442 GND.n1449 240.244
R10854 GND.n4438 GND.n1449 240.244
R10855 GND.n4438 GND.n1457 240.244
R10856 GND.n1475 GND.n1457 240.244
R10857 GND.n4428 GND.n1475 240.244
R10858 GND.n4428 GND.n1476 240.244
R10859 GND.n4424 GND.n1476 240.244
R10860 GND.n4424 GND.n1484 240.244
R10861 GND.n4414 GND.n1484 240.244
R10862 GND.n4414 GND.n1495 240.244
R10863 GND.n4410 GND.n1495 240.244
R10864 GND.n4410 GND.n1501 240.244
R10865 GND.n4400 GND.n1501 240.244
R10866 GND.n4400 GND.n1513 240.244
R10867 GND.n4396 GND.n1513 240.244
R10868 GND.n4396 GND.n1519 240.244
R10869 GND.n4386 GND.n1519 240.244
R10870 GND.n4386 GND.n1533 240.244
R10871 GND.n4382 GND.n1533 240.244
R10872 GND.n4382 GND.n1539 240.244
R10873 GND.n1566 GND.n1539 240.244
R10874 GND.n1566 GND.n1562 240.244
R10875 GND.n4365 GND.n1562 240.244
R10876 GND.n4365 GND.n1563 240.244
R10877 GND.n4361 GND.n1563 240.244
R10878 GND.n4361 GND.n1574 240.244
R10879 GND.n1609 GND.n1574 240.244
R10880 GND.n1609 GND.n1605 240.244
R10881 GND.n4344 GND.n1605 240.244
R10882 GND.n4344 GND.n1606 240.244
R10883 GND.n4340 GND.n1606 240.244
R10884 GND.n4340 GND.n1617 240.244
R10885 GND.n3409 GND.n1617 240.244
R10886 GND.n3416 GND.n3409 240.244
R10887 GND.n3416 GND.n1654 240.244
R10888 GND.n4317 GND.n1654 240.244
R10889 GND.n4317 GND.n1655 240.244
R10890 GND.n4313 GND.n1655 240.244
R10891 GND.n4313 GND.n1661 240.244
R10892 GND.n3763 GND.n1661 240.244
R10893 GND.n3764 GND.n3763 240.244
R10894 GND.n3764 GND.n3758 240.244
R10895 GND.n3771 GND.n3758 240.244
R10896 GND.n3771 GND.n1698 240.244
R10897 GND.n4289 GND.n1698 240.244
R10898 GND.n4289 GND.n1699 240.244
R10899 GND.n4285 GND.n1699 240.244
R10900 GND.n4285 GND.n1705 240.244
R10901 GND.n1723 GND.n1705 240.244
R10902 GND.n4275 GND.n1723 240.244
R10903 GND.n4275 GND.n1724 240.244
R10904 GND.n4271 GND.n1724 240.244
R10905 GND.n4271 GND.n1732 240.244
R10906 GND.n1749 GND.n1732 240.244
R10907 GND.n4261 GND.n1749 240.244
R10908 GND.n4261 GND.n1750 240.244
R10909 GND.n4257 GND.n1750 240.244
R10910 GND.n4257 GND.n1758 240.244
R10911 GND.n2126 GND.n1758 240.244
R10912 GND.n2128 GND.n2126 240.244
R10913 GND.n2128 GND.n2121 240.244
R10914 GND.n2134 GND.n2121 240.244
R10915 GND.n2135 GND.n2134 240.244
R10916 GND.n3845 GND.n2135 240.244
R10917 GND.n3845 GND.n2116 240.244
R10918 GND.n3887 GND.n2116 240.244
R10919 GND.n3887 GND.n2117 240.244
R10920 GND.n3883 GND.n2117 240.244
R10921 GND.n3883 GND.n3882 240.244
R10922 GND.n3882 GND.n3881 240.244
R10923 GND.n3881 GND.n3853 240.244
R10924 GND.n3877 GND.n3853 240.244
R10925 GND.n3877 GND.n3876 240.244
R10926 GND.n3876 GND.n3873 240.244
R10927 GND.n3873 GND.n3859 240.244
R10928 GND.n3869 GND.n3859 240.244
R10929 GND.n3869 GND.n3868 240.244
R10930 GND.n3868 GND.n2049 240.244
R10931 GND.n3965 GND.n2049 240.244
R10932 GND.n3966 GND.n3965 240.244
R10933 GND.n3966 GND.n2044 240.244
R10934 GND.n3976 GND.n2044 240.244
R10935 GND.n3976 GND.n2045 240.244
R10936 GND.n2045 GND.n2015 240.244
R10937 GND.n4004 GND.n2015 240.244
R10938 GND.n4005 GND.n4004 240.244
R10939 GND.n4005 GND.n2012 240.244
R10940 GND.n4055 GND.n2012 240.244
R10941 GND.n4055 GND.n2013 240.244
R10942 GND.n4050 GND.n2013 240.244
R10943 GND.n4050 GND.n4010 240.244
R10944 GND.n4033 GND.n4010 240.244
R10945 GND.n4038 GND.n4033 240.244
R10946 GND.n4038 GND.n1986 240.244
R10947 GND.n4073 GND.n1986 240.244
R10948 GND.n4073 GND.n1981 240.244
R10949 GND.n4081 GND.n1981 240.244
R10950 GND.n4081 GND.n1982 240.244
R10951 GND.n1982 GND.n1962 240.244
R10952 GND.n4099 GND.n1962 240.244
R10953 GND.n4099 GND.n1957 240.244
R10954 GND.n4114 GND.n1957 240.244
R10955 GND.n4114 GND.n1958 240.244
R10956 GND.n4110 GND.n1958 240.244
R10957 GND.n4110 GND.n4109 240.244
R10958 GND.n4109 GND.n595 240.244
R10959 GND.n5485 GND.n595 240.244
R10960 GND.n5485 GND.n596 240.244
R10961 GND.n5481 GND.n596 240.244
R10962 GND.n4883 GND.n958 240.244
R10963 GND.n4879 GND.n958 240.244
R10964 GND.n4879 GND.n960 240.244
R10965 GND.n4875 GND.n960 240.244
R10966 GND.n4875 GND.n965 240.244
R10967 GND.n4871 GND.n965 240.244
R10968 GND.n4871 GND.n967 240.244
R10969 GND.n4867 GND.n967 240.244
R10970 GND.n4867 GND.n973 240.244
R10971 GND.n4863 GND.n973 240.244
R10972 GND.n4863 GND.n975 240.244
R10973 GND.n4859 GND.n975 240.244
R10974 GND.n4859 GND.n981 240.244
R10975 GND.n4855 GND.n981 240.244
R10976 GND.n4855 GND.n983 240.244
R10977 GND.n4851 GND.n983 240.244
R10978 GND.n4851 GND.n989 240.244
R10979 GND.n4847 GND.n989 240.244
R10980 GND.n4847 GND.n991 240.244
R10981 GND.n4843 GND.n991 240.244
R10982 GND.n4843 GND.n997 240.244
R10983 GND.n4839 GND.n997 240.244
R10984 GND.n4839 GND.n999 240.244
R10985 GND.n4835 GND.n999 240.244
R10986 GND.n4835 GND.n1005 240.244
R10987 GND.n4831 GND.n1005 240.244
R10988 GND.n4831 GND.n1007 240.244
R10989 GND.n4827 GND.n1007 240.244
R10990 GND.n4827 GND.n1013 240.244
R10991 GND.n4823 GND.n1013 240.244
R10992 GND.n4823 GND.n1015 240.244
R10993 GND.n4819 GND.n1015 240.244
R10994 GND.n4819 GND.n1021 240.244
R10995 GND.n4815 GND.n1021 240.244
R10996 GND.n4815 GND.n1023 240.244
R10997 GND.n4811 GND.n1023 240.244
R10998 GND.n4811 GND.n1029 240.244
R10999 GND.n4807 GND.n1029 240.244
R11000 GND.n4807 GND.n1031 240.244
R11001 GND.n4803 GND.n1031 240.244
R11002 GND.n4803 GND.n1037 240.244
R11003 GND.n4799 GND.n1037 240.244
R11004 GND.n4799 GND.n1039 240.244
R11005 GND.n4795 GND.n1039 240.244
R11006 GND.n4795 GND.n1045 240.244
R11007 GND.n4791 GND.n1045 240.244
R11008 GND.n4791 GND.n1047 240.244
R11009 GND.n4787 GND.n1047 240.244
R11010 GND.n4787 GND.n1053 240.244
R11011 GND.n4783 GND.n1053 240.244
R11012 GND.n4783 GND.n1055 240.244
R11013 GND.n4779 GND.n1055 240.244
R11014 GND.n4779 GND.n1061 240.244
R11015 GND.n4775 GND.n1061 240.244
R11016 GND.n4775 GND.n1063 240.244
R11017 GND.n4771 GND.n1063 240.244
R11018 GND.n4771 GND.n1069 240.244
R11019 GND.n4767 GND.n1069 240.244
R11020 GND.n4767 GND.n1071 240.244
R11021 GND.n4763 GND.n1071 240.244
R11022 GND.n4763 GND.n1077 240.244
R11023 GND.n4759 GND.n1077 240.244
R11024 GND.n4759 GND.n1079 240.244
R11025 GND.n4755 GND.n1079 240.244
R11026 GND.n4755 GND.n1085 240.244
R11027 GND.n2541 GND.n1085 240.244
R11028 GND.n4213 GND.n1853 240.244
R11029 GND.n4203 GND.n4202 240.244
R11030 GND.n1783 GND.n1782 240.244
R11031 GND.n1843 GND.n1790 240.244
R11032 GND.n1846 GND.n1791 240.244
R11033 GND.n1801 GND.n1800 240.244
R11034 GND.n1848 GND.n1808 240.244
R11035 GND.n1821 GND.n1809 240.244
R11036 GND.n2115 GND.n1852 240.244
R11037 GND.n3892 GND.n2115 240.244
R11038 GND.n3892 GND.n3891 240.244
R11039 GND.n3891 GND.n2104 240.244
R11040 GND.n2104 GND.n2094 240.244
R11041 GND.n3913 GND.n2094 240.244
R11042 GND.n3916 GND.n3913 240.244
R11043 GND.n3916 GND.n3915 240.244
R11044 GND.n3915 GND.n2082 240.244
R11045 GND.n2082 GND.n2071 240.244
R11046 GND.n3937 GND.n2071 240.244
R11047 GND.n3941 GND.n3937 240.244
R11048 GND.n3941 GND.n3940 240.244
R11049 GND.n3940 GND.n2061 240.244
R11050 GND.n2061 GND.n2060 240.244
R11051 GND.n2060 GND.n2039 240.244
R11052 GND.n3981 GND.n2039 240.244
R11053 GND.n3981 GND.n3979 240.244
R11054 GND.n3979 GND.n2040 240.244
R11055 GND.n2040 GND.n2028 240.244
R11056 GND.n2028 GND.n2027 240.244
R11057 GND.n2027 GND.n2005 240.244
R11058 GND.n4059 GND.n2005 240.244
R11059 GND.n4059 GND.n4058 240.244
R11060 GND.n4058 GND.n2007 240.244
R11061 GND.n4015 GND.n2007 240.244
R11062 GND.n4016 GND.n4015 240.244
R11063 GND.n4042 GND.n4016 240.244
R11064 GND.n4042 GND.n4041 240.244
R11065 GND.n4041 GND.n4025 240.244
R11066 GND.n4025 GND.n4024 240.244
R11067 GND.n4024 GND.n1990 240.244
R11068 GND.n1990 GND.n1978 240.244
R11069 GND.n4084 GND.n1978 240.244
R11070 GND.n4086 GND.n4084 240.244
R11071 GND.n4086 GND.n4085 240.244
R11072 GND.n4085 GND.n1967 240.244
R11073 GND.n1967 GND.n1955 240.244
R11074 GND.n4118 GND.n1955 240.244
R11075 GND.n4119 GND.n4118 240.244
R11076 GND.n4119 GND.n1942 240.244
R11077 GND.n4131 GND.n1942 240.244
R11078 GND.n4132 GND.n4131 240.244
R11079 GND.n4132 GND.n584 240.244
R11080 GND.n5494 GND.n584 240.244
R11081 GND.n5494 GND.n585 240.244
R11082 GND.n585 GND.n574 240.244
R11083 GND.n574 GND.n565 240.244
R11084 GND.n5512 GND.n565 240.244
R11085 GND.n5512 GND.n555 240.244
R11086 GND.n5523 GND.n555 240.244
R11087 GND.n5569 GND.n5523 240.244
R11088 GND.n5527 GND.n5526 240.244
R11089 GND.n5529 GND.n5528 240.244
R11090 GND.n5533 GND.n5532 240.244
R11091 GND.n5535 GND.n5534 240.244
R11092 GND.n5539 GND.n5538 240.244
R11093 GND.n5541 GND.n5540 240.244
R11094 GND.n5544 GND.n5543 240.244
R11095 GND.n5631 GND.n466 240.244
R11096 GND.n3842 GND.n1820 240.244
R11097 GND.n3842 GND.n2113 240.244
R11098 GND.n2113 GND.n2101 240.244
R11099 GND.n3904 GND.n2101 240.244
R11100 GND.n3904 GND.n2096 240.244
R11101 GND.n3911 GND.n2096 240.244
R11102 GND.n3911 GND.n2091 240.244
R11103 GND.n2091 GND.n2079 240.244
R11104 GND.n3928 GND.n2079 240.244
R11105 GND.n3928 GND.n2074 240.244
R11106 GND.n3935 GND.n2074 240.244
R11107 GND.n3935 GND.n2069 240.244
R11108 GND.n2069 GND.n2057 240.244
R11109 GND.n3953 GND.n2057 240.244
R11110 GND.n3953 GND.n2052 240.244
R11111 GND.n3962 GND.n2052 240.244
R11112 GND.n3962 GND.n2037 240.244
R11113 GND.n2041 GND.n2037 240.244
R11114 GND.n2041 GND.n2023 240.244
R11115 GND.n3992 GND.n2023 240.244
R11116 GND.n3992 GND.n2018 240.244
R11117 GND.n4001 GND.n2018 240.244
R11118 GND.n4001 GND.n2004 240.244
R11119 GND.n2009 GND.n2004 240.244
R11120 GND.n2010 GND.n2009 240.244
R11121 GND.n2010 GND.n429 240.244
R11122 GND.n430 GND.n429 240.244
R11123 GND.n431 GND.n430 240.244
R11124 GND.n4028 GND.n431 240.244
R11125 GND.n4028 GND.n434 240.244
R11126 GND.n435 GND.n434 240.244
R11127 GND.n436 GND.n435 240.244
R11128 GND.n1979 GND.n436 240.244
R11129 GND.n1979 GND.n439 240.244
R11130 GND.n440 GND.n439 240.244
R11131 GND.n441 GND.n440 240.244
R11132 GND.n1964 GND.n441 240.244
R11133 GND.n1964 GND.n444 240.244
R11134 GND.n445 GND.n444 240.244
R11135 GND.n446 GND.n445 240.244
R11136 GND.n1952 GND.n446 240.244
R11137 GND.n1952 GND.n449 240.244
R11138 GND.n450 GND.n449 240.244
R11139 GND.n451 GND.n450 240.244
R11140 GND.n582 GND.n451 240.244
R11141 GND.n582 GND.n454 240.244
R11142 GND.n455 GND.n454 240.244
R11143 GND.n456 GND.n455 240.244
R11144 GND.n564 GND.n456 240.244
R11145 GND.n564 GND.n459 240.244
R11146 GND.n460 GND.n459 240.244
R11147 GND.n461 GND.n460 240.244
R11148 GND.n2250 GND.n2249 240.132
R11149 GND.n3505 GND.n3504 240.132
R11150 GND.n463 GND.t157 224.174
R11151 GND.n519 GND.t151 224.174
R11152 GND.n546 GND.t80 224.174
R11153 GND.n1286 GND.t145 224.174
R11154 GND.n1312 GND.t76 224.174
R11155 GND.n1372 GND.t136 224.174
R11156 GND.n2587 GND.t155 224.174
R11157 GND.n3625 GND.t85 224.174
R11158 GND.n3647 GND.t101 224.174
R11159 GND.n1131 GND.t105 224.174
R11160 GND.n1151 GND.t123 224.174
R11161 GND.n1810 GND.t140 224.174
R11162 GND.n5630 GND.n476 222.413
R11163 GND.n5313 GND.n696 209.825
R11164 GND.n5321 GND.n696 209.825
R11165 GND.n5322 GND.n5321 209.825
R11166 GND.n5323 GND.n5322 209.825
R11167 GND.n5323 GND.n690 209.825
R11168 GND.n5331 GND.n690 209.825
R11169 GND.n5332 GND.n5331 209.825
R11170 GND.n5333 GND.n5332 209.825
R11171 GND.n5333 GND.n684 209.825
R11172 GND.n5341 GND.n684 209.825
R11173 GND.n5342 GND.n5341 209.825
R11174 GND.n5343 GND.n5342 209.825
R11175 GND.n5343 GND.n678 209.825
R11176 GND.n5351 GND.n678 209.825
R11177 GND.n5352 GND.n5351 209.825
R11178 GND.n5353 GND.n5352 209.825
R11179 GND.n5353 GND.n672 209.825
R11180 GND.n5361 GND.n672 209.825
R11181 GND.n5362 GND.n5361 209.825
R11182 GND.n5363 GND.n5362 209.825
R11183 GND.n5363 GND.n666 209.825
R11184 GND.n5371 GND.n666 209.825
R11185 GND.n5372 GND.n5371 209.825
R11186 GND.n5373 GND.n5372 209.825
R11187 GND.n5373 GND.n660 209.825
R11188 GND.n5381 GND.n660 209.825
R11189 GND.n5382 GND.n5381 209.825
R11190 GND.n5383 GND.n5382 209.825
R11191 GND.n5383 GND.n654 209.825
R11192 GND.n5391 GND.n654 209.825
R11193 GND.n5392 GND.n5391 209.825
R11194 GND.n5393 GND.n5392 209.825
R11195 GND.n5393 GND.n648 209.825
R11196 GND.n5401 GND.n648 209.825
R11197 GND.n5402 GND.n5401 209.825
R11198 GND.n5403 GND.n5402 209.825
R11199 GND.n5403 GND.n642 209.825
R11200 GND.n5411 GND.n642 209.825
R11201 GND.n5412 GND.n5411 209.825
R11202 GND.n5413 GND.n5412 209.825
R11203 GND.n5413 GND.n636 209.825
R11204 GND.n5421 GND.n636 209.825
R11205 GND.n5422 GND.n5421 209.825
R11206 GND.n5423 GND.n5422 209.825
R11207 GND.n5423 GND.n630 209.825
R11208 GND.n5431 GND.n630 209.825
R11209 GND.n5432 GND.n5431 209.825
R11210 GND.n5433 GND.n5432 209.825
R11211 GND.n5433 GND.n624 209.825
R11212 GND.n5441 GND.n624 209.825
R11213 GND.n5442 GND.n5441 209.825
R11214 GND.n5443 GND.n5442 209.825
R11215 GND.n5443 GND.n618 209.825
R11216 GND.n5451 GND.n618 209.825
R11217 GND.n5452 GND.n5451 209.825
R11218 GND.n5453 GND.n5452 209.825
R11219 GND.n5453 GND.n612 209.825
R11220 GND.n5461 GND.n612 209.825
R11221 GND.n5462 GND.n5461 209.825
R11222 GND.n5463 GND.n5462 209.825
R11223 GND.n5463 GND.n606 209.825
R11224 GND.n5471 GND.n606 209.825
R11225 GND.n5472 GND.n5471 209.825
R11226 GND.n5473 GND.n5472 209.825
R11227 GND.n5473 GND.n476 209.825
R11228 GND.n3580 GND.n1831 199.319
R11229 GND.n4491 GND.n1289 199.319
R11230 GND.n4490 GND.n1289 199.319
R11231 GND.n2251 GND.n2248 186.49
R11232 GND.n3506 GND.n3503 186.49
R11233 GND.n96 GND.n95 185
R11234 GND.n94 GND.n93 185
R11235 GND.n73 GND.n72 185
R11236 GND.n88 GND.n87 185
R11237 GND.n86 GND.n85 185
R11238 GND.n77 GND.n76 185
R11239 GND.n80 GND.n79 185
R11240 GND.n133 GND.n132 185
R11241 GND.n131 GND.n130 185
R11242 GND.n110 GND.n109 185
R11243 GND.n125 GND.n124 185
R11244 GND.n123 GND.n122 185
R11245 GND.n114 GND.n113 185
R11246 GND.n117 GND.n116 185
R11247 GND.n165 GND.n164 185
R11248 GND.n163 GND.n162 185
R11249 GND.n142 GND.n141 185
R11250 GND.n157 GND.n156 185
R11251 GND.n155 GND.n154 185
R11252 GND.n146 GND.n145 185
R11253 GND.n149 GND.n148 185
R11254 GND.n202 GND.n201 185
R11255 GND.n200 GND.n199 185
R11256 GND.n179 GND.n178 185
R11257 GND.n194 GND.n193 185
R11258 GND.n192 GND.n191 185
R11259 GND.n183 GND.n182 185
R11260 GND.n186 GND.n185 185
R11261 GND.n27 GND.n26 185
R11262 GND.n25 GND.n24 185
R11263 GND.n4 GND.n3 185
R11264 GND.n19 GND.n18 185
R11265 GND.n17 GND.n16 185
R11266 GND.n8 GND.n7 185
R11267 GND.n11 GND.n10 185
R11268 GND.n64 GND.n63 185
R11269 GND.n62 GND.n61 185
R11270 GND.n41 GND.n40 185
R11271 GND.n56 GND.n55 185
R11272 GND.n54 GND.n53 185
R11273 GND.n45 GND.n44 185
R11274 GND.n48 GND.n47 185
R11275 GND.n281 GND.n280 185
R11276 GND.n279 GND.n278 185
R11277 GND.n258 GND.n257 185
R11278 GND.n273 GND.n272 185
R11279 GND.n271 GND.n270 185
R11280 GND.n262 GND.n261 185
R11281 GND.n265 GND.n264 185
R11282 GND.n244 GND.n243 185
R11283 GND.n242 GND.n241 185
R11284 GND.n221 GND.n220 185
R11285 GND.n236 GND.n235 185
R11286 GND.n234 GND.n233 185
R11287 GND.n225 GND.n224 185
R11288 GND.n228 GND.n227 185
R11289 GND.n350 GND.n349 185
R11290 GND.n348 GND.n347 185
R11291 GND.n327 GND.n326 185
R11292 GND.n342 GND.n341 185
R11293 GND.n340 GND.n339 185
R11294 GND.n331 GND.n330 185
R11295 GND.n334 GND.n333 185
R11296 GND.n313 GND.n312 185
R11297 GND.n311 GND.n310 185
R11298 GND.n290 GND.n289 185
R11299 GND.n305 GND.n304 185
R11300 GND.n303 GND.n302 185
R11301 GND.n294 GND.n293 185
R11302 GND.n297 GND.n296 185
R11303 GND.n420 GND.n419 185
R11304 GND.n418 GND.n417 185
R11305 GND.n397 GND.n396 185
R11306 GND.n412 GND.n411 185
R11307 GND.n410 GND.n409 185
R11308 GND.n401 GND.n400 185
R11309 GND.n404 GND.n403 185
R11310 GND.n383 GND.n382 185
R11311 GND.n381 GND.n380 185
R11312 GND.n360 GND.n359 185
R11313 GND.n375 GND.n374 185
R11314 GND.n373 GND.n372 185
R11315 GND.n364 GND.n363 185
R11316 GND.n367 GND.n366 185
R11317 GND.n464 GND.t158 178.987
R11318 GND.n520 GND.t152 178.987
R11319 GND.n547 GND.t81 178.987
R11320 GND.n1287 GND.t146 178.987
R11321 GND.n1313 GND.t77 178.987
R11322 GND.n1373 GND.t137 178.987
R11323 GND.n2588 GND.t154 178.987
R11324 GND.n3626 GND.t84 178.987
R11325 GND.n3648 GND.t100 178.987
R11326 GND.n1132 GND.t104 178.987
R11327 GND.n1152 GND.t122 178.987
R11328 GND.n1811 GND.t139 178.987
R11329 GND.n210 GND.t15 171.065
R11330 GND.n212 GND.t17 170.103
R11331 GND.n211 GND.t35 170.103
R11332 GND.n210 GND.t37 170.103
R11333 GND.n3518 GND.n3517 163.367
R11334 GND.n3522 GND.n3521 163.367
R11335 GND.n3526 GND.n3525 163.367
R11336 GND.n3530 GND.n3529 163.367
R11337 GND.n3534 GND.n3533 163.367
R11338 GND.n3538 GND.n3537 163.367
R11339 GND.n3542 GND.n3541 163.367
R11340 GND.n3546 GND.n3545 163.367
R11341 GND.n3550 GND.n3549 163.367
R11342 GND.n3554 GND.n3553 163.367
R11343 GND.n3558 GND.n3557 163.367
R11344 GND.n3562 GND.n3561 163.367
R11345 GND.n3566 GND.n3565 163.367
R11346 GND.n3570 GND.n3569 163.367
R11347 GND.n3575 GND.n3574 163.367
R11348 GND.n3687 GND.n3686 163.367
R11349 GND.n3754 GND.n3753 163.367
R11350 GND.n3750 GND.n3749 163.367
R11351 GND.n3745 GND.n3744 163.367
R11352 GND.n3741 GND.n3740 163.367
R11353 GND.n3737 GND.n3736 163.367
R11354 GND.n3733 GND.n3732 163.367
R11355 GND.n3729 GND.n3728 163.367
R11356 GND.n3725 GND.n3724 163.367
R11357 GND.n3721 GND.n3720 163.367
R11358 GND.n3717 GND.n3716 163.367
R11359 GND.n3713 GND.n3712 163.367
R11360 GND.n3709 GND.n3708 163.367
R11361 GND.n3705 GND.n3704 163.367
R11362 GND.n3701 GND.n3700 163.367
R11363 GND.n3697 GND.n3696 163.367
R11364 GND.n3693 GND.n3692 163.367
R11365 GND.n3069 GND.n2242 163.367
R11366 GND.n3153 GND.n2242 163.367
R11367 GND.n3153 GND.n1486 163.367
R11368 GND.n3150 GND.n1486 163.367
R11369 GND.n3150 GND.n1493 163.367
R11370 GND.n3146 GND.n1493 163.367
R11371 GND.n3146 GND.n3145 163.367
R11372 GND.n3145 GND.n3144 163.367
R11373 GND.n3144 GND.n1503 163.367
R11374 GND.n3140 GND.n1503 163.367
R11375 GND.n3140 GND.n1511 163.367
R11376 GND.n2220 GND.n1511 163.367
R11377 GND.n3295 GND.n2220 163.367
R11378 GND.n3296 GND.n3295 163.367
R11379 GND.n3296 GND.n1521 163.367
R11380 GND.n3300 GND.n1521 163.367
R11381 GND.n3300 GND.n1531 163.367
R11382 GND.n3305 GND.n1531 163.367
R11383 GND.n3305 GND.n2217 163.367
R11384 GND.n3310 GND.n2217 163.367
R11385 GND.n3310 GND.n2218 163.367
R11386 GND.n2218 GND.n2208 163.367
R11387 GND.n3351 GND.n2208 163.367
R11388 GND.n3351 GND.n1552 163.367
R11389 GND.n3355 GND.n1552 163.367
R11390 GND.n3355 GND.n1560 163.367
R11391 GND.n3359 GND.n1560 163.367
R11392 GND.n3363 GND.n3359 163.367
R11393 GND.n3363 GND.n1576 163.367
R11394 GND.n3367 GND.n1576 163.367
R11395 GND.n3367 GND.n1584 163.367
R11396 GND.n2205 GND.n1584 163.367
R11397 GND.n3384 GND.n2205 163.367
R11398 GND.n3384 GND.n2206 163.367
R11399 GND.n3380 GND.n2206 163.367
R11400 GND.n3380 GND.n2199 163.367
R11401 GND.n3377 GND.n2199 163.367
R11402 GND.n3377 GND.n1619 163.367
R11403 GND.n3373 GND.n1619 163.367
R11404 GND.n3373 GND.n1627 163.367
R11405 GND.n2191 GND.n1627 163.367
R11406 GND.n3419 GND.n2191 163.367
R11407 GND.n3419 GND.n1644 163.367
R11408 GND.n3423 GND.n1644 163.367
R11409 GND.n3423 GND.n1652 163.367
R11410 GND.n2188 GND.n1652 163.367
R11411 GND.n3431 GND.n2188 163.367
R11412 GND.n3431 GND.n2189 163.367
R11413 GND.n3427 GND.n2189 163.367
R11414 GND.n3427 GND.n2179 163.367
R11415 GND.n3452 GND.n2179 163.367
R11416 GND.n3452 GND.n1680 163.367
R11417 GND.n3778 GND.n1680 163.367
R11418 GND.n3778 GND.n1687 163.367
R11419 GND.n3774 GND.n1687 163.367
R11420 GND.n3222 GND.n2265 163.367
R11421 GND.n3222 GND.n3160 163.367
R11422 GND.n3218 GND.n3217 163.367
R11423 GND.n3214 GND.n3213 163.367
R11424 GND.n3210 GND.n3209 163.367
R11425 GND.n3206 GND.n3205 163.367
R11426 GND.n3202 GND.n3201 163.367
R11427 GND.n3198 GND.n3197 163.367
R11428 GND.n3194 GND.n3193 163.367
R11429 GND.n3190 GND.n3189 163.367
R11430 GND.n3186 GND.n3185 163.367
R11431 GND.n3182 GND.n3181 163.367
R11432 GND.n3178 GND.n3177 163.367
R11433 GND.n3174 GND.n3173 163.367
R11434 GND.n3170 GND.n3169 163.367
R11435 GND.n3166 GND.n3165 163.367
R11436 GND.n3073 GND.n3072 163.367
R11437 GND.n3077 GND.n3076 163.367
R11438 GND.n3082 GND.n3081 163.367
R11439 GND.n3086 GND.n3085 163.367
R11440 GND.n3090 GND.n3089 163.367
R11441 GND.n3094 GND.n3093 163.367
R11442 GND.n3098 GND.n3097 163.367
R11443 GND.n3102 GND.n3101 163.367
R11444 GND.n3106 GND.n3105 163.367
R11445 GND.n3110 GND.n3109 163.367
R11446 GND.n3114 GND.n3113 163.367
R11447 GND.n3118 GND.n3117 163.367
R11448 GND.n3122 GND.n3121 163.367
R11449 GND.n3126 GND.n3125 163.367
R11450 GND.n3130 GND.n3129 163.367
R11451 GND.n3132 GND.n3068 163.367
R11452 GND.n3230 GND.n2243 163.367
R11453 GND.n3230 GND.n1487 163.367
R11454 GND.n4421 GND.n1487 163.367
R11455 GND.n4421 GND.n1488 163.367
R11456 GND.n4417 GND.n1488 163.367
R11457 GND.n4417 GND.n1491 163.367
R11458 GND.n2229 GND.n1491 163.367
R11459 GND.n2229 GND.n1505 163.367
R11460 GND.n4407 GND.n1505 163.367
R11461 GND.n4407 GND.n1506 163.367
R11462 GND.n4403 GND.n1506 163.367
R11463 GND.n4403 GND.n1509 163.367
R11464 GND.n3293 GND.n1509 163.367
R11465 GND.n3293 GND.n1525 163.367
R11466 GND.n4393 GND.n1525 163.367
R11467 GND.n4393 GND.n1526 163.367
R11468 GND.n4389 GND.n1526 163.367
R11469 GND.n4389 GND.n1529 163.367
R11470 GND.n3311 GND.n1529 163.367
R11471 GND.n3318 GND.n3311 163.367
R11472 GND.n3318 GND.n3312 163.367
R11473 GND.n3314 GND.n3312 163.367
R11474 GND.n3314 GND.n1554 163.367
R11475 GND.n4372 GND.n1554 163.367
R11476 GND.n4372 GND.n1555 163.367
R11477 GND.n4368 GND.n1555 163.367
R11478 GND.n4368 GND.n1558 163.367
R11479 GND.n1578 GND.n1558 163.367
R11480 GND.n4358 GND.n1578 163.367
R11481 GND.n4358 GND.n1579 163.367
R11482 GND.n4354 GND.n1579 163.367
R11483 GND.n4354 GND.n1582 163.367
R11484 GND.n3387 GND.n1582 163.367
R11485 GND.n3388 GND.n3387 163.367
R11486 GND.n3388 GND.n2201 163.367
R11487 GND.n3392 GND.n2201 163.367
R11488 GND.n3392 GND.n1621 163.367
R11489 GND.n4337 GND.n1621 163.367
R11490 GND.n4337 GND.n1622 163.367
R11491 GND.n4333 GND.n1622 163.367
R11492 GND.n4333 GND.n1625 163.367
R11493 GND.n1646 GND.n1625 163.367
R11494 GND.n4324 GND.n1646 163.367
R11495 GND.n4324 GND.n1647 163.367
R11496 GND.n4320 GND.n1647 163.367
R11497 GND.n4320 GND.n1650 163.367
R11498 GND.n3439 GND.n1650 163.367
R11499 GND.n3439 GND.n3432 163.367
R11500 GND.n3435 GND.n3432 163.367
R11501 GND.n3435 GND.n3434 163.367
R11502 GND.n3434 GND.n1681 163.367
R11503 GND.n4303 GND.n1681 163.367
R11504 GND.n4303 GND.n1682 163.367
R11505 GND.n4299 GND.n1682 163.367
R11506 GND.n4299 GND.n1685 163.367
R11507 GND.n3512 GND.n3511 156.462
R11508 GND.n2256 GND.n2255 152
R11509 GND.n2257 GND.n2246 152
R11510 GND.n2259 GND.n2258 152
R11511 GND.n2261 GND.n2244 152
R11512 GND.n2263 GND.n2262 152
R11513 GND.n3510 GND.n3494 152
R11514 GND.n3502 GND.n3495 152
R11515 GND.n3501 GND.n3500 152
R11516 GND.n3499 GND.n3496 152
R11517 GND.n3497 GND.t115 150.546
R11518 GND.t39 GND.n78 147.661
R11519 GND.t53 GND.n115 147.661
R11520 GND.t177 GND.n147 147.661
R11521 GND.t165 GND.n184 147.661
R11522 GND.t168 GND.n9 147.661
R11523 GND.t1 GND.n46 147.661
R11524 GND.t25 GND.n263 147.661
R11525 GND.t58 GND.n226 147.661
R11526 GND.t55 GND.n332 147.661
R11527 GND.t159 GND.n295 147.661
R11528 GND.t56 GND.n402 147.661
R11529 GND.t171 GND.n365 147.661
R11530 GND.n3491 GND.n3474 143.351
R11531 GND.n3051 GND.n3050 143.351
R11532 GND.n3052 GND.n3051 143.351
R11533 GND.n2253 GND.t147 130.484
R11534 GND.n2262 GND.t96 126.766
R11535 GND.n2260 GND.t109 126.766
R11536 GND.n2246 GND.t86 126.766
R11537 GND.n2254 GND.t118 126.766
R11538 GND.n3498 GND.t71 126.766
R11539 GND.n3500 GND.t141 126.766
R11540 GND.n3509 GND.t93 126.766
R11541 GND.n3511 GND.t112 126.766
R11542 GND.n2158 GND.t133 118.023
R11543 GND.n2988 GND.t127 118.023
R11544 GND.n4575 GND.n1290 110.912
R11545 GND.n3688 GND.n3685 110.912
R11546 GND.n95 GND.n94 104.615
R11547 GND.n94 GND.n72 104.615
R11548 GND.n87 GND.n72 104.615
R11549 GND.n87 GND.n86 104.615
R11550 GND.n86 GND.n76 104.615
R11551 GND.n79 GND.n76 104.615
R11552 GND.n132 GND.n131 104.615
R11553 GND.n131 GND.n109 104.615
R11554 GND.n124 GND.n109 104.615
R11555 GND.n124 GND.n123 104.615
R11556 GND.n123 GND.n113 104.615
R11557 GND.n116 GND.n113 104.615
R11558 GND.n164 GND.n163 104.615
R11559 GND.n163 GND.n141 104.615
R11560 GND.n156 GND.n141 104.615
R11561 GND.n156 GND.n155 104.615
R11562 GND.n155 GND.n145 104.615
R11563 GND.n148 GND.n145 104.615
R11564 GND.n201 GND.n200 104.615
R11565 GND.n200 GND.n178 104.615
R11566 GND.n193 GND.n178 104.615
R11567 GND.n193 GND.n192 104.615
R11568 GND.n192 GND.n182 104.615
R11569 GND.n185 GND.n182 104.615
R11570 GND.n26 GND.n25 104.615
R11571 GND.n25 GND.n3 104.615
R11572 GND.n18 GND.n3 104.615
R11573 GND.n18 GND.n17 104.615
R11574 GND.n17 GND.n7 104.615
R11575 GND.n10 GND.n7 104.615
R11576 GND.n63 GND.n62 104.615
R11577 GND.n62 GND.n40 104.615
R11578 GND.n55 GND.n40 104.615
R11579 GND.n55 GND.n54 104.615
R11580 GND.n54 GND.n44 104.615
R11581 GND.n47 GND.n44 104.615
R11582 GND.n280 GND.n279 104.615
R11583 GND.n279 GND.n257 104.615
R11584 GND.n272 GND.n257 104.615
R11585 GND.n272 GND.n271 104.615
R11586 GND.n271 GND.n261 104.615
R11587 GND.n264 GND.n261 104.615
R11588 GND.n243 GND.n242 104.615
R11589 GND.n242 GND.n220 104.615
R11590 GND.n235 GND.n220 104.615
R11591 GND.n235 GND.n234 104.615
R11592 GND.n234 GND.n224 104.615
R11593 GND.n227 GND.n224 104.615
R11594 GND.n349 GND.n348 104.615
R11595 GND.n348 GND.n326 104.615
R11596 GND.n341 GND.n326 104.615
R11597 GND.n341 GND.n340 104.615
R11598 GND.n340 GND.n330 104.615
R11599 GND.n333 GND.n330 104.615
R11600 GND.n312 GND.n311 104.615
R11601 GND.n311 GND.n289 104.615
R11602 GND.n304 GND.n289 104.615
R11603 GND.n304 GND.n303 104.615
R11604 GND.n303 GND.n293 104.615
R11605 GND.n296 GND.n293 104.615
R11606 GND.n419 GND.n418 104.615
R11607 GND.n418 GND.n396 104.615
R11608 GND.n411 GND.n396 104.615
R11609 GND.n411 GND.n410 104.615
R11610 GND.n410 GND.n400 104.615
R11611 GND.n403 GND.n400 104.615
R11612 GND.n382 GND.n381 104.615
R11613 GND.n381 GND.n359 104.615
R11614 GND.n374 GND.n359 104.615
R11615 GND.n374 GND.n373 104.615
R11616 GND.n373 GND.n363 104.615
R11617 GND.n366 GND.n363 104.615
R11618 GND.n499 GND.n493 99.6594
R11619 GND.n501 GND.n492 99.6594
R11620 GND.n505 GND.n491 99.6594
R11621 GND.n507 GND.n490 99.6594
R11622 GND.n511 GND.n489 99.6594
R11623 GND.n513 GND.n488 99.6594
R11624 GND.n517 GND.n487 99.6594
R11625 GND.n521 GND.n486 99.6594
R11626 GND.n525 GND.n485 99.6594
R11627 GND.n527 GND.n484 99.6594
R11628 GND.n531 GND.n483 99.6594
R11629 GND.n533 GND.n482 99.6594
R11630 GND.n537 GND.n481 99.6594
R11631 GND.n539 GND.n480 99.6594
R11632 GND.n543 GND.n479 99.6594
R11633 GND.n545 GND.n478 99.6594
R11634 GND.n5574 GND.n477 99.6594
R11635 GND.n3590 GND.n1823 99.6594
R11636 GND.n3596 GND.n1824 99.6594
R11637 GND.n3600 GND.n1825 99.6594
R11638 GND.n3606 GND.n1826 99.6594
R11639 GND.n3610 GND.n1827 99.6594
R11640 GND.n3616 GND.n1828 99.6594
R11641 GND.n3620 GND.n1829 99.6594
R11642 GND.n3580 GND.n1830 99.6594
R11643 GND.n3682 GND.n1832 99.6594
R11644 GND.n3678 GND.n1833 99.6594
R11645 GND.n3674 GND.n1834 99.6594
R11646 GND.n3670 GND.n1835 99.6594
R11647 GND.n3666 GND.n1836 99.6594
R11648 GND.n3662 GND.n1837 99.6594
R11649 GND.n3658 GND.n1838 99.6594
R11650 GND.n3654 GND.n1839 99.6594
R11651 GND.n3646 GND.n1840 99.6594
R11652 GND.n4500 GND.n1271 99.6594
R11653 GND.n4499 GND.n1274 99.6594
R11654 GND.n4497 GND.n1276 99.6594
R11655 GND.n4496 GND.n1279 99.6594
R11656 GND.n4494 GND.n1281 99.6594
R11657 GND.n4493 GND.n1284 99.6594
R11658 GND.n4490 GND.n1291 99.6594
R11659 GND.n4489 GND.n1294 99.6594
R11660 GND.n4487 GND.n1296 99.6594
R11661 GND.n4486 GND.n1299 99.6594
R11662 GND.n4484 GND.n1301 99.6594
R11663 GND.n4483 GND.n1304 99.6594
R11664 GND.n4481 GND.n1306 99.6594
R11665 GND.n4480 GND.n1309 99.6594
R11666 GND.n4478 GND.n1311 99.6594
R11667 GND.n4477 GND.n1260 99.6594
R11668 GND.n4751 GND.n4750 99.6594
R11669 GND.n4745 GND.n1086 99.6594
R11670 GND.n4742 GND.n1087 99.6594
R11671 GND.n4738 GND.n1088 99.6594
R11672 GND.n4734 GND.n1089 99.6594
R11673 GND.n4730 GND.n1090 99.6594
R11674 GND.n4726 GND.n1091 99.6594
R11675 GND.n4722 GND.n1092 99.6594
R11676 GND.n4717 GND.n1093 99.6594
R11677 GND.n4713 GND.n1094 99.6594
R11678 GND.n4709 GND.n1095 99.6594
R11679 GND.n4705 GND.n1096 99.6594
R11680 GND.n4701 GND.n1097 99.6594
R11681 GND.n4697 GND.n1098 99.6594
R11682 GND.n4693 GND.n1099 99.6594
R11683 GND.n4689 GND.n1100 99.6594
R11684 GND.n1150 GND.n1101 99.6594
R11685 GND.n1377 GND.n1318 99.6594
R11686 GND.n1381 GND.n1379 99.6594
R11687 GND.n1383 GND.n1346 99.6594
R11688 GND.n1385 GND.n1384 99.6594
R11689 GND.n1386 GND.n1355 99.6594
R11690 GND.n1388 GND.n1364 99.6594
R11691 GND.n1390 GND.n1389 99.6594
R11692 GND.n4503 GND.n4502 99.6594
R11693 GND.n2613 GND.n1102 99.6594
R11694 GND.n2556 GND.n1103 99.6594
R11695 GND.n2560 GND.n1104 99.6594
R11696 GND.n2562 GND.n1105 99.6594
R11697 GND.n2566 GND.n1106 99.6594
R11698 GND.n2568 GND.n1107 99.6594
R11699 GND.n2572 GND.n1108 99.6594
R11700 GND.n2574 GND.n1109 99.6594
R11701 GND.n1786 GND.n1775 99.6594
R11702 GND.n1794 GND.n1774 99.6594
R11703 GND.n1796 GND.n1773 99.6594
R11704 GND.n1804 GND.n1772 99.6594
R11705 GND.n1814 GND.n1771 99.6594
R11706 GND.n1816 GND.n1770 99.6594
R11707 GND.n2143 GND.n1769 99.6594
R11708 GND.n2145 GND.n1768 99.6594
R11709 GND.n2149 GND.n1767 99.6594
R11710 GND.n2151 GND.n1766 99.6594
R11711 GND.n2155 GND.n1765 99.6594
R11712 GND.n2157 GND.n1764 99.6594
R11713 GND.n2163 GND.n1763 99.6594
R11714 GND.n3814 GND.n1762 99.6594
R11715 GND.n4536 GND.n4535 99.6594
R11716 GND.n1340 GND.n1326 99.6594
R11717 GND.n1351 GND.n1327 99.6594
R11718 GND.n1359 GND.n1328 99.6594
R11719 GND.n1361 GND.n1329 99.6594
R11720 GND.n1369 GND.n1330 99.6594
R11721 GND.n2283 GND.n1331 99.6594
R11722 GND.n2964 GND.n1332 99.6594
R11723 GND.n2966 GND.n1333 99.6594
R11724 GND.n2974 GND.n1334 99.6594
R11725 GND.n2976 GND.n1335 99.6594
R11726 GND.n2984 GND.n1336 99.6594
R11727 GND.n2986 GND.n1337 99.6594
R11728 GND.n2997 GND.n1338 99.6594
R11729 GND.n4535 GND.n1324 99.6594
R11730 GND.n1350 GND.n1326 99.6594
R11731 GND.n1358 GND.n1327 99.6594
R11732 GND.n1360 GND.n1328 99.6594
R11733 GND.n1368 GND.n1329 99.6594
R11734 GND.n2282 GND.n1330 99.6594
R11735 GND.n2963 GND.n1331 99.6594
R11736 GND.n2967 GND.n1332 99.6594
R11737 GND.n2973 GND.n1333 99.6594
R11738 GND.n2977 GND.n1334 99.6594
R11739 GND.n2983 GND.n1335 99.6594
R11740 GND.n2987 GND.n1336 99.6594
R11741 GND.n2996 GND.n1337 99.6594
R11742 GND.n2999 GND.n1338 99.6594
R11743 GND.n2164 GND.n1762 99.6594
R11744 GND.n2160 GND.n1763 99.6594
R11745 GND.n2156 GND.n1764 99.6594
R11746 GND.n2152 GND.n1765 99.6594
R11747 GND.n2150 GND.n1766 99.6594
R11748 GND.n2146 GND.n1767 99.6594
R11749 GND.n2144 GND.n1768 99.6594
R11750 GND.n1817 GND.n1769 99.6594
R11751 GND.n1815 GND.n1770 99.6594
R11752 GND.n1805 GND.n1771 99.6594
R11753 GND.n1797 GND.n1772 99.6594
R11754 GND.n1795 GND.n1773 99.6594
R11755 GND.n1787 GND.n1774 99.6594
R11756 GND.n1777 GND.n1775 99.6594
R11757 GND.n2555 GND.n1102 99.6594
R11758 GND.n2559 GND.n1103 99.6594
R11759 GND.n2561 GND.n1104 99.6594
R11760 GND.n2565 GND.n1105 99.6594
R11761 GND.n2567 GND.n1106 99.6594
R11762 GND.n2571 GND.n1107 99.6594
R11763 GND.n2573 GND.n1108 99.6594
R11764 GND.n2586 GND.n1109 99.6594
R11765 GND.n4502 GND.n1374 99.6594
R11766 GND.n1390 GND.n1365 99.6594
R11767 GND.n1388 GND.n1387 99.6594
R11768 GND.n1386 GND.n1354 99.6594
R11769 GND.n1385 GND.n1347 99.6594
R11770 GND.n1383 GND.n1382 99.6594
R11771 GND.n1379 GND.n1378 99.6594
R11772 GND.n1377 GND.n1317 99.6594
R11773 GND.n4751 GND.n1113 99.6594
R11774 GND.n4743 GND.n1086 99.6594
R11775 GND.n4739 GND.n1087 99.6594
R11776 GND.n4735 GND.n1088 99.6594
R11777 GND.n4731 GND.n1089 99.6594
R11778 GND.n4727 GND.n1090 99.6594
R11779 GND.n4723 GND.n1091 99.6594
R11780 GND.n4718 GND.n1092 99.6594
R11781 GND.n4714 GND.n1093 99.6594
R11782 GND.n4710 GND.n1094 99.6594
R11783 GND.n4706 GND.n1095 99.6594
R11784 GND.n4702 GND.n1096 99.6594
R11785 GND.n4698 GND.n1097 99.6594
R11786 GND.n4694 GND.n1098 99.6594
R11787 GND.n4690 GND.n1099 99.6594
R11788 GND.n1149 GND.n1100 99.6594
R11789 GND.n4682 GND.n1101 99.6594
R11790 GND.n4477 GND.n4476 99.6594
R11791 GND.n4478 GND.n1310 99.6594
R11792 GND.n4480 GND.n4479 99.6594
R11793 GND.n4481 GND.n1305 99.6594
R11794 GND.n4483 GND.n4482 99.6594
R11795 GND.n4484 GND.n1300 99.6594
R11796 GND.n4486 GND.n4485 99.6594
R11797 GND.n4487 GND.n1295 99.6594
R11798 GND.n4489 GND.n4488 99.6594
R11799 GND.n4491 GND.n1285 99.6594
R11800 GND.n4493 GND.n4492 99.6594
R11801 GND.n4494 GND.n1280 99.6594
R11802 GND.n4496 GND.n4495 99.6594
R11803 GND.n4497 GND.n1275 99.6594
R11804 GND.n4499 GND.n4498 99.6594
R11805 GND.n4500 GND.n1270 99.6594
R11806 GND.n3595 GND.n1823 99.6594
R11807 GND.n3599 GND.n1824 99.6594
R11808 GND.n3605 GND.n1825 99.6594
R11809 GND.n3609 GND.n1826 99.6594
R11810 GND.n3615 GND.n1827 99.6594
R11811 GND.n3619 GND.n1828 99.6594
R11812 GND.n3578 GND.n1829 99.6594
R11813 GND.n3683 GND.n1831 99.6594
R11814 GND.n3679 GND.n1832 99.6594
R11815 GND.n3675 GND.n1833 99.6594
R11816 GND.n3671 GND.n1834 99.6594
R11817 GND.n3667 GND.n1835 99.6594
R11818 GND.n3663 GND.n1836 99.6594
R11819 GND.n3659 GND.n1837 99.6594
R11820 GND.n3655 GND.n1838 99.6594
R11821 GND.n3643 GND.n1839 99.6594
R11822 GND.n3644 GND.n1840 99.6594
R11823 GND.n548 GND.n477 99.6594
R11824 GND.n544 GND.n478 99.6594
R11825 GND.n540 GND.n479 99.6594
R11826 GND.n538 GND.n480 99.6594
R11827 GND.n534 GND.n481 99.6594
R11828 GND.n532 GND.n482 99.6594
R11829 GND.n528 GND.n483 99.6594
R11830 GND.n526 GND.n484 99.6594
R11831 GND.n522 GND.n485 99.6594
R11832 GND.n518 GND.n486 99.6594
R11833 GND.n514 GND.n487 99.6594
R11834 GND.n512 GND.n488 99.6594
R11835 GND.n508 GND.n489 99.6594
R11836 GND.n506 GND.n490 99.6594
R11837 GND.n502 GND.n491 99.6594
R11838 GND.n500 GND.n492 99.6594
R11839 GND.n495 GND.n493 99.6594
R11840 GND.n1853 GND.n1841 99.6594
R11841 GND.n4202 GND.n1842 99.6594
R11842 GND.n1844 GND.n1783 99.6594
R11843 GND.n1845 GND.n1790 99.6594
R11844 GND.n1847 GND.n1846 99.6594
R11845 GND.n1849 GND.n1801 99.6594
R11846 GND.n1850 GND.n1808 99.6594
R11847 GND.n4215 GND.n1821 99.6594
R11848 GND.n4203 GND.n1841 99.6594
R11849 GND.n1842 GND.n1782 99.6594
R11850 GND.n1844 GND.n1843 99.6594
R11851 GND.n1845 GND.n1791 99.6594
R11852 GND.n1847 GND.n1800 99.6594
R11853 GND.n1849 GND.n1848 99.6594
R11854 GND.n1850 GND.n1809 99.6594
R11855 GND.n4216 GND.n4215 99.6594
R11856 GND.n5568 GND.n468 99.6594
R11857 GND.n5527 GND.n469 99.6594
R11858 GND.n5529 GND.n470 99.6594
R11859 GND.n5533 GND.n471 99.6594
R11860 GND.n5535 GND.n472 99.6594
R11861 GND.n5539 GND.n473 99.6594
R11862 GND.n5541 GND.n474 99.6594
R11863 GND.n5544 GND.n475 99.6594
R11864 GND.n475 GND.n466 99.6594
R11865 GND.n5543 GND.n474 99.6594
R11866 GND.n5540 GND.n473 99.6594
R11867 GND.n5538 GND.n472 99.6594
R11868 GND.n5534 GND.n471 99.6594
R11869 GND.n5532 GND.n470 99.6594
R11870 GND.n5528 GND.n469 99.6594
R11871 GND.n5526 GND.n468 99.6594
R11872 GND.n3070 GND.t92 98.6378
R11873 GND.n3689 GND.t107 98.6378
R11874 GND.n3161 GND.t130 98.63
R11875 GND.n3492 GND.t69 98.63
R11876 GND.n2253 GND.n2252 81.8399
R11877 GND.n3071 GND.t91 72.8438
R11878 GND.n3690 GND.t108 72.8438
R11879 GND.n2254 GND.n2247 72.8411
R11880 GND.n2260 GND.n2245 72.8411
R11881 GND.n3509 GND.n3508 72.8411
R11882 GND.n3162 GND.t129 72.836
R11883 GND.n3493 GND.t70 72.836
R11884 GND.n2159 GND.t134 72.836
R11885 GND.n2989 GND.t126 72.836
R11886 GND.n3517 GND.n3458 71.676
R11887 GND.n3521 GND.n3459 71.676
R11888 GND.n3525 GND.n3460 71.676
R11889 GND.n3529 GND.n3461 71.676
R11890 GND.n3533 GND.n3462 71.676
R11891 GND.n3537 GND.n3463 71.676
R11892 GND.n3541 GND.n3464 71.676
R11893 GND.n3545 GND.n3465 71.676
R11894 GND.n3549 GND.n3466 71.676
R11895 GND.n3553 GND.n3467 71.676
R11896 GND.n3557 GND.n3468 71.676
R11897 GND.n3561 GND.n3469 71.676
R11898 GND.n3565 GND.n3470 71.676
R11899 GND.n3569 GND.n3471 71.676
R11900 GND.n3574 GND.n3472 71.676
R11901 GND.n3686 GND.n3473 71.676
R11902 GND.n3754 GND.n3491 71.676
R11903 GND.n3750 GND.n3490 71.676
R11904 GND.n3745 GND.n3489 71.676
R11905 GND.n3741 GND.n3488 71.676
R11906 GND.n3737 GND.n3487 71.676
R11907 GND.n3733 GND.n3486 71.676
R11908 GND.n3729 GND.n3485 71.676
R11909 GND.n3725 GND.n3484 71.676
R11910 GND.n3721 GND.n3483 71.676
R11911 GND.n3717 GND.n3482 71.676
R11912 GND.n3713 GND.n3481 71.676
R11913 GND.n3709 GND.n3480 71.676
R11914 GND.n3705 GND.n3479 71.676
R11915 GND.n3701 GND.n3478 71.676
R11916 GND.n3697 GND.n3477 71.676
R11917 GND.n3693 GND.n3476 71.676
R11918 GND.n3475 GND.n3456 71.676
R11919 GND.n3225 GND.n3224 71.676
R11920 GND.n3160 GND.n3036 71.676
R11921 GND.n3217 GND.n3037 71.676
R11922 GND.n3213 GND.n3038 71.676
R11923 GND.n3209 GND.n3039 71.676
R11924 GND.n3205 GND.n3040 71.676
R11925 GND.n3201 GND.n3041 71.676
R11926 GND.n3197 GND.n3042 71.676
R11927 GND.n3193 GND.n3043 71.676
R11928 GND.n3189 GND.n3044 71.676
R11929 GND.n3185 GND.n3045 71.676
R11930 GND.n3181 GND.n3046 71.676
R11931 GND.n3177 GND.n3047 71.676
R11932 GND.n3173 GND.n3048 71.676
R11933 GND.n3169 GND.n3049 71.676
R11934 GND.n3165 GND.n3050 71.676
R11935 GND.n3073 GND.n3053 71.676
R11936 GND.n3077 GND.n3054 71.676
R11937 GND.n3082 GND.n3055 71.676
R11938 GND.n3086 GND.n3056 71.676
R11939 GND.n3090 GND.n3057 71.676
R11940 GND.n3094 GND.n3058 71.676
R11941 GND.n3098 GND.n3059 71.676
R11942 GND.n3102 GND.n3060 71.676
R11943 GND.n3106 GND.n3061 71.676
R11944 GND.n3110 GND.n3062 71.676
R11945 GND.n3114 GND.n3063 71.676
R11946 GND.n3118 GND.n3064 71.676
R11947 GND.n3122 GND.n3065 71.676
R11948 GND.n3126 GND.n3066 71.676
R11949 GND.n3130 GND.n3067 71.676
R11950 GND.n3159 GND.n3068 71.676
R11951 GND.n3224 GND.n2265 71.676
R11952 GND.n3218 GND.n3036 71.676
R11953 GND.n3214 GND.n3037 71.676
R11954 GND.n3210 GND.n3038 71.676
R11955 GND.n3206 GND.n3039 71.676
R11956 GND.n3202 GND.n3040 71.676
R11957 GND.n3198 GND.n3041 71.676
R11958 GND.n3194 GND.n3042 71.676
R11959 GND.n3190 GND.n3043 71.676
R11960 GND.n3186 GND.n3044 71.676
R11961 GND.n3182 GND.n3045 71.676
R11962 GND.n3178 GND.n3046 71.676
R11963 GND.n3174 GND.n3047 71.676
R11964 GND.n3170 GND.n3048 71.676
R11965 GND.n3166 GND.n3049 71.676
R11966 GND.n3072 GND.n3052 71.676
R11967 GND.n3076 GND.n3053 71.676
R11968 GND.n3081 GND.n3054 71.676
R11969 GND.n3085 GND.n3055 71.676
R11970 GND.n3089 GND.n3056 71.676
R11971 GND.n3093 GND.n3057 71.676
R11972 GND.n3097 GND.n3058 71.676
R11973 GND.n3101 GND.n3059 71.676
R11974 GND.n3105 GND.n3060 71.676
R11975 GND.n3109 GND.n3061 71.676
R11976 GND.n3113 GND.n3062 71.676
R11977 GND.n3117 GND.n3063 71.676
R11978 GND.n3121 GND.n3064 71.676
R11979 GND.n3125 GND.n3065 71.676
R11980 GND.n3129 GND.n3066 71.676
R11981 GND.n3132 GND.n3067 71.676
R11982 GND.n3159 GND.n3158 71.676
R11983 GND.n3692 GND.n3475 71.676
R11984 GND.n3696 GND.n3476 71.676
R11985 GND.n3700 GND.n3477 71.676
R11986 GND.n3704 GND.n3478 71.676
R11987 GND.n3708 GND.n3479 71.676
R11988 GND.n3712 GND.n3480 71.676
R11989 GND.n3716 GND.n3481 71.676
R11990 GND.n3720 GND.n3482 71.676
R11991 GND.n3724 GND.n3483 71.676
R11992 GND.n3728 GND.n3484 71.676
R11993 GND.n3732 GND.n3485 71.676
R11994 GND.n3736 GND.n3486 71.676
R11995 GND.n3740 GND.n3487 71.676
R11996 GND.n3744 GND.n3488 71.676
R11997 GND.n3749 GND.n3489 71.676
R11998 GND.n3753 GND.n3490 71.676
R11999 GND.n3687 GND.n3474 71.676
R12000 GND.n3575 GND.n3473 71.676
R12001 GND.n3570 GND.n3472 71.676
R12002 GND.n3566 GND.n3471 71.676
R12003 GND.n3562 GND.n3470 71.676
R12004 GND.n3558 GND.n3469 71.676
R12005 GND.n3554 GND.n3468 71.676
R12006 GND.n3550 GND.n3467 71.676
R12007 GND.n3546 GND.n3466 71.676
R12008 GND.n3542 GND.n3465 71.676
R12009 GND.n3538 GND.n3464 71.676
R12010 GND.n3534 GND.n3463 71.676
R12011 GND.n3530 GND.n3462 71.676
R12012 GND.n3526 GND.n3461 71.676
R12013 GND.n3522 GND.n3460 71.676
R12014 GND.n3518 GND.n3459 71.676
R12015 GND.n3514 GND.n3458 71.676
R12016 GND.n213 GND.t174 69.4414
R12017 GND.n215 GND.t23 68.4792
R12018 GND.n214 GND.t19 68.4792
R12019 GND.n213 GND.t12 68.4792
R12020 GND.n3079 GND.n3071 59.5399
R12021 GND.n3747 GND.n3690 59.5399
R12022 GND.n3163 GND.n3162 59.5399
R12023 GND.n3572 GND.n3493 59.5399
R12024 GND.n3227 GND.n2263 59.1804
R12025 GND.n101 GND.n100 56.1363
R12026 GND.n103 GND.n102 56.1363
R12027 GND.n105 GND.n104 56.1363
R12028 GND.n170 GND.n169 56.1363
R12029 GND.n172 GND.n171 56.1363
R12030 GND.n174 GND.n173 56.1363
R12031 GND.n32 GND.n31 56.1363
R12032 GND.n34 GND.n33 56.1363
R12033 GND.n36 GND.n35 56.1363
R12034 GND.n253 GND.n252 56.1363
R12035 GND.n251 GND.n250 56.1363
R12036 GND.n249 GND.n248 56.1363
R12037 GND.n322 GND.n321 56.1363
R12038 GND.n320 GND.n319 56.1363
R12039 GND.n318 GND.n317 56.1363
R12040 GND.n392 GND.n391 56.1363
R12041 GND.n390 GND.n389 56.1363
R12042 GND.n388 GND.n387 56.1363
R12043 GND.n2251 GND.n2250 54.358
R12044 GND.n3506 GND.n3505 54.358
R12045 GND.n4752 GND.n1111 52.5321
R12046 GND.n5630 GND.n467 52.5321
R12047 GND.n3497 GND.n3496 52.4801
R12048 GND.n79 GND.t39 52.3082
R12049 GND.n116 GND.t53 52.3082
R12050 GND.n148 GND.t177 52.3082
R12051 GND.n185 GND.t165 52.3082
R12052 GND.n10 GND.t168 52.3082
R12053 GND.n47 GND.t1 52.3082
R12054 GND.n264 GND.t25 52.3082
R12055 GND.n227 GND.t58 52.3082
R12056 GND.n333 GND.t55 52.3082
R12057 GND.n296 GND.t159 52.3082
R12058 GND.n403 GND.t56 52.3082
R12059 GND.n366 GND.t171 52.3082
R12060 GND.n4882 GND.n4881 50.3322
R12061 GND.n4881 GND.n4880 50.3322
R12062 GND.n4880 GND.n959 50.3322
R12063 GND.n4874 GND.n959 50.3322
R12064 GND.n4874 GND.n4873 50.3322
R12065 GND.n4873 GND.n4872 50.3322
R12066 GND.n4872 GND.n966 50.3322
R12067 GND.n4866 GND.n966 50.3322
R12068 GND.n4866 GND.n4865 50.3322
R12069 GND.n4865 GND.n4864 50.3322
R12070 GND.n4864 GND.n974 50.3322
R12071 GND.n4858 GND.n974 50.3322
R12072 GND.n4858 GND.n4857 50.3322
R12073 GND.n4857 GND.n4856 50.3322
R12074 GND.n4856 GND.n982 50.3322
R12075 GND.n4850 GND.n982 50.3322
R12076 GND.n4850 GND.n4849 50.3322
R12077 GND.n4849 GND.n4848 50.3322
R12078 GND.n4848 GND.n990 50.3322
R12079 GND.n4842 GND.n990 50.3322
R12080 GND.n4842 GND.n4841 50.3322
R12081 GND.n4841 GND.n4840 50.3322
R12082 GND.n4840 GND.n998 50.3322
R12083 GND.n4834 GND.n998 50.3322
R12084 GND.n4834 GND.n4833 50.3322
R12085 GND.n4833 GND.n4832 50.3322
R12086 GND.n4832 GND.n1006 50.3322
R12087 GND.n4826 GND.n1006 50.3322
R12088 GND.n4826 GND.n4825 50.3322
R12089 GND.n4825 GND.n4824 50.3322
R12090 GND.n4824 GND.n1014 50.3322
R12091 GND.n4818 GND.n1014 50.3322
R12092 GND.n4818 GND.n4817 50.3322
R12093 GND.n4817 GND.n4816 50.3322
R12094 GND.n4816 GND.n1022 50.3322
R12095 GND.n4810 GND.n1022 50.3322
R12096 GND.n4810 GND.n4809 50.3322
R12097 GND.n4809 GND.n4808 50.3322
R12098 GND.n4808 GND.n1030 50.3322
R12099 GND.n4802 GND.n1030 50.3322
R12100 GND.n4802 GND.n4801 50.3322
R12101 GND.n4801 GND.n4800 50.3322
R12102 GND.n4800 GND.n1038 50.3322
R12103 GND.n4794 GND.n1038 50.3322
R12104 GND.n4794 GND.n4793 50.3322
R12105 GND.n4793 GND.n4792 50.3322
R12106 GND.n4792 GND.n1046 50.3322
R12107 GND.n4786 GND.n1046 50.3322
R12108 GND.n4786 GND.n4785 50.3322
R12109 GND.n4785 GND.n4784 50.3322
R12110 GND.n4784 GND.n1054 50.3322
R12111 GND.n4778 GND.n1054 50.3322
R12112 GND.n4778 GND.n4777 50.3322
R12113 GND.n4777 GND.n4776 50.3322
R12114 GND.n4776 GND.n1062 50.3322
R12115 GND.n4770 GND.n1062 50.3322
R12116 GND.n4770 GND.n4769 50.3322
R12117 GND.n4769 GND.n4768 50.3322
R12118 GND.n4768 GND.n1070 50.3322
R12119 GND.n4762 GND.n1070 50.3322
R12120 GND.n4762 GND.n4761 50.3322
R12121 GND.n4761 GND.n4760 50.3322
R12122 GND.n4760 GND.n1078 50.3322
R12123 GND.n4754 GND.n1078 50.3322
R12124 GND.n4754 GND.n4753 50.3322
R12125 GND.n464 GND.n463 45.1884
R12126 GND.n520 GND.n519 45.1884
R12127 GND.n547 GND.n546 45.1884
R12128 GND.n1287 GND.n1286 45.1884
R12129 GND.n1313 GND.n1312 45.1884
R12130 GND.n1373 GND.n1372 45.1884
R12131 GND.n2588 GND.n2587 45.1884
R12132 GND.n2159 GND.n2158 45.1884
R12133 GND.n2989 GND.n2988 45.1884
R12134 GND.n3626 GND.n3625 45.1884
R12135 GND.n3648 GND.n3647 45.1884
R12136 GND.n1132 GND.n1131 45.1884
R12137 GND.n1152 GND.n1151 45.1884
R12138 GND.n1811 GND.n1810 45.1884
R12139 GND.n3513 GND.n3512 44.3322
R12140 GND.n2254 GND.n2253 44.3189
R12141 GND.n465 GND.n464 42.2793
R12142 GND.n5604 GND.n520 42.2793
R12143 GND.n549 GND.n547 42.2793
R12144 GND.n1314 GND.n1313 42.2793
R12145 GND.n4505 GND.n1373 42.2793
R12146 GND.n2589 GND.n2588 42.2793
R12147 GND.n3821 GND.n2159 42.2793
R12148 GND.n2990 GND.n2989 42.2793
R12149 GND.n3649 GND.n3648 42.2793
R12150 GND.n4720 GND.n1132 42.2793
R12151 GND.n1153 GND.n1152 42.2793
R12152 GND.n1812 GND.n1811 42.2793
R12153 GND.n2252 GND.n2251 41.6274
R12154 GND.n3507 GND.n3506 41.6274
R12155 GND.n2261 GND.n2260 40.8975
R12156 GND.n3510 GND.n3509 40.8975
R12157 GND.n101 GND.n99 38.8139
R12158 GND.n170 GND.n168 38.8139
R12159 GND.n32 GND.n30 38.8139
R12160 GND.n249 GND.n247 38.8139
R12161 GND.n318 GND.n316 38.8139
R12162 GND.n388 GND.n386 38.8139
R12163 GND.n137 GND.n136 37.8096
R12164 GND.n206 GND.n205 37.8096
R12165 GND.n68 GND.n67 37.8096
R12166 GND.n285 GND.n284 37.8096
R12167 GND.n354 GND.n353 37.8096
R12168 GND.n424 GND.n423 37.8096
R12169 GND.n4575 GND.n1287 36.9518
R12170 GND.n3685 GND.n3626 36.9518
R12171 GND.n2260 GND.n2259 35.055
R12172 GND.n2255 GND.n2254 35.055
R12173 GND.n3499 GND.n3498 35.055
R12174 GND.n3509 GND.n3495 35.055
R12175 GND.n3775 GND.n3455 33.2493
R12176 GND.n3157 GND.n3156 33.2493
R12177 GND.n2552 GND.n1111 31.6461
R12178 GND.n2619 GND.n2552 31.6461
R12179 GND.n2629 GND.n2504 31.6461
R12180 GND.n2638 GND.n2497 31.6461
R12181 GND.n1376 GND.n1263 31.6461
R12182 GND.n4475 GND.n1391 31.6461
R12183 GND.n1391 GND.n1325 31.6461
R12184 GND.n4467 GND.n1339 31.6461
R12185 GND.n4256 GND.n4255 31.6461
R12186 GND.n2127 GND.n1761 31.6461
R12187 GND.n2127 GND.n1822 31.6461
R12188 GND.n2136 GND.n1851 31.6461
R12189 GND.n5503 GND.n572 31.6461
R12190 GND.n5513 GND.n562 31.6461
R12191 GND.n5522 GND.n556 31.6461
R12192 GND.n5522 GND.n467 31.6461
R12193 GND.n2644 GND.n2492 30.3802
R12194 GND.n2640 GND.n2494 30.3802
R12195 GND.n2654 GND.n2481 30.3802
R12196 GND.n2663 GND.n2474 30.3802
R12197 GND.n2669 GND.n2469 30.3802
R12198 GND.n2666 GND.n2471 30.3802
R12199 GND.n2679 GND.n2459 30.3802
R12200 GND.n2702 GND.n2452 30.3802
R12201 GND.n2706 GND.n2446 30.3802
R12202 GND.n2449 GND.n2435 30.3802
R12203 GND.n2716 GND.n2715 30.3802
R12204 GND.n2690 GND.n2686 30.3802
R12205 GND.n2687 GND.n2427 30.3802
R12206 GND.n2729 GND.n2728 30.3802
R12207 GND.n2826 GND.n2389 30.3802
R12208 GND.n2821 GND.n2396 30.3802
R12209 GND.n2403 GND.n2402 30.3802
R12210 GND.n2814 GND.n2813 30.3802
R12211 GND.n2808 GND.n2405 30.3802
R12212 GND.n2804 GND.n2746 30.3802
R12213 GND.n2836 GND.n2373 30.3802
R12214 GND.n2795 GND.n2374 30.3802
R12215 GND.n2851 GND.n2362 30.3802
R12216 GND.n2848 GND.n2364 30.3802
R12217 GND.n2861 GND.n2353 30.3802
R12218 GND.n2786 GND.n2354 30.3802
R12219 GND.n2876 GND.n2343 30.3802
R12220 GND.n2872 GND.n2345 30.3802
R12221 GND.n2886 GND.n2333 30.3802
R12222 GND.n2765 GND.n2335 30.3802
R12223 GND.n2902 GND.n2322 30.3802
R12224 GND.n2324 GND.n2316 30.3802
R12225 GND.n2911 GND.n2910 30.3802
R12226 GND.n2939 GND.n2301 30.3802
R12227 GND.n2942 GND.n2296 30.3802
R12228 GND.n2931 GND.n2298 30.3802
R12229 GND.n2955 GND.n2289 30.3802
R12230 GND.n4600 GND.n1261 30.3802
R12231 GND.n3844 GND.n2137 30.3802
R12232 GND.n3843 GND.n2112 30.3802
R12233 GND.n3890 GND.n2102 30.3802
R12234 GND.n3903 GND.n2103 30.3802
R12235 GND.n2106 GND.n2095 30.3802
R12236 GND.n3912 GND.n2089 30.3802
R12237 GND.n3917 GND.n2092 30.3802
R12238 GND.n3914 GND.n2080 30.3802
R12239 GND.n3874 GND.n2072 30.3802
R12240 GND.n3936 GND.n2068 30.3802
R12241 GND.n3942 GND.n2070 30.3802
R12242 GND.n3939 GND.n2058 30.3802
R12243 GND.n3964 GND.n2051 30.3802
R12244 GND.n3963 GND.n2036 30.3802
R12245 GND.n3982 GND.n2038 30.3802
R12246 GND.n3978 GND.n3977 30.3802
R12247 GND.n3991 GND.n2025 30.3802
R12248 GND.n4003 GND.n2017 30.3802
R12249 GND.n4002 GND.n2002 30.3802
R12250 GND.n4057 GND.n4056 30.3802
R12251 GND.n4011 GND.n2011 30.3802
R12252 GND.n4049 GND.n4012 30.3802
R12253 GND.n4048 GND.n4014 30.3802
R12254 GND.n4040 GND.n4039 30.3802
R12255 GND.n4032 GND.n4029 30.3802
R12256 GND.n4072 GND.n1988 30.3802
R12257 GND.n4071 GND.n1989 30.3802
R12258 GND.n4082 GND.n1980 30.3802
R12259 GND.n4083 GND.n1974 30.3802
R12260 GND.n4087 GND.n1976 30.3802
R12261 GND.n4098 GND.n1963 30.3802
R12262 GND.n4115 GND.n1956 30.3802
R12263 GND.n4117 GND.n1951 30.3802
R12264 GND.n4120 GND.n1954 30.3802
R12265 GND.n1953 GND.n1943 30.3802
R12266 GND.n5486 GND.n594 30.3802
R12267 GND.n5487 GND.n580 30.3802
R12268 GND.n5495 GND.n583 30.3802
R12269 GND.n2796 GND.t42 30.0638
R12270 GND.t4 GND.n2024 30.0638
R12271 GND.n2619 GND.t103 26.8992
R12272 GND.n2950 GND.t75 26.8992
R12273 GND.n3893 GND.t83 26.8992
R12274 GND.t79 GND.n556 26.8992
R12275 GND.n3071 GND.n3070 25.7944
R12276 GND.n3690 GND.n3689 25.7944
R12277 GND.n3162 GND.n3161 25.7944
R12278 GND.n3493 GND.n3492 25.7944
R12279 GND.n2898 GND.t38 21.8359
R12280 GND.n3927 GND.t57 21.8359
R12281 GND.n2805 GND.t32 21.203
R12282 GND.n4060 GND.t160 21.203
R12283 GND.n3228 GND.n3227 21.0737
R12284 GND.n3513 GND.n1684 21.0737
R12285 GND.t0 GND.n2483 20.5701
R12286 GND.n2463 GND.t40 20.5701
R12287 GND.n4097 GND.t2 20.5701
R12288 GND.t24 GND.n1944 20.5701
R12289 GND.n2542 GND.n2497 19.9372
R12290 GND.t61 GND.n2391 19.9372
R12291 GND.n4027 GND.t48 19.9372
R12292 GND.n5503 GND.n573 19.9372
R12293 GND.n2248 GND.t120 19.8005
R12294 GND.n2248 GND.t149 19.8005
R12295 GND.n2249 GND.t111 19.8005
R12296 GND.n2249 GND.t88 19.8005
R12297 GND.n3503 GND.t95 19.8005
R12298 GND.n3503 GND.t114 19.8005
R12299 GND.n3504 GND.t73 19.8005
R12300 GND.n3504 GND.t143 19.8005
R12301 GND.n4501 GND.n1376 19.6208
R12302 GND.n4214 GND.n1851 19.6208
R12303 GND.n2245 GND.n2244 19.5087
R12304 GND.n2258 GND.n2245 19.5087
R12305 GND.n2256 GND.n2247 19.5087
R12306 GND.n3508 GND.n3502 19.5087
R12307 GND.n5567 GND.n5524 19.3944
R12308 GND.n5563 GND.n5524 19.3944
R12309 GND.n5563 GND.n5562 19.3944
R12310 GND.n5562 GND.n5561 19.3944
R12311 GND.n5561 GND.n5530 19.3944
R12312 GND.n5557 GND.n5530 19.3944
R12313 GND.n5557 GND.n5556 19.3944
R12314 GND.n5556 GND.n5555 19.3944
R12315 GND.n5555 GND.n5536 19.3944
R12316 GND.n5551 GND.n5536 19.3944
R12317 GND.n5551 GND.n5550 19.3944
R12318 GND.n5550 GND.n5549 19.3944
R12319 GND.n5549 GND.n5542 19.3944
R12320 GND.n5545 GND.n5542 19.3944
R12321 GND.n2114 GND.n1855 19.3944
R12322 GND.n2114 GND.n1861 19.3944
R12323 GND.n1862 GND.n1861 19.3944
R12324 GND.n1863 GND.n1862 19.3944
R12325 GND.n2093 GND.n1863 19.3944
R12326 GND.n2093 GND.n1869 19.3944
R12327 GND.n1870 GND.n1869 19.3944
R12328 GND.n1871 GND.n1870 19.3944
R12329 GND.n2081 GND.n1871 19.3944
R12330 GND.n2081 GND.n1877 19.3944
R12331 GND.n1878 GND.n1877 19.3944
R12332 GND.n1879 GND.n1878 19.3944
R12333 GND.n3938 GND.n1879 19.3944
R12334 GND.n3938 GND.n1885 19.3944
R12335 GND.n1886 GND.n1885 19.3944
R12336 GND.n1887 GND.n1886 19.3944
R12337 GND.n3980 GND.n1887 19.3944
R12338 GND.n3980 GND.n1893 19.3944
R12339 GND.n1894 GND.n1893 19.3944
R12340 GND.n1895 GND.n1894 19.3944
R12341 GND.n2026 GND.n1895 19.3944
R12342 GND.n2026 GND.n1901 19.3944
R12343 GND.n1902 GND.n1901 19.3944
R12344 GND.n1903 GND.n1902 19.3944
R12345 GND.n2006 GND.n1903 19.3944
R12346 GND.n2006 GND.n1909 19.3944
R12347 GND.n1910 GND.n1909 19.3944
R12348 GND.n1911 GND.n1910 19.3944
R12349 GND.n4026 GND.n1911 19.3944
R12350 GND.n4026 GND.n1917 19.3944
R12351 GND.n1918 GND.n1917 19.3944
R12352 GND.n1919 GND.n1918 19.3944
R12353 GND.n1977 GND.n1919 19.3944
R12354 GND.n1977 GND.n1925 19.3944
R12355 GND.n1926 GND.n1925 19.3944
R12356 GND.n1927 GND.n1926 19.3944
R12357 GND.n1966 GND.n1927 19.3944
R12358 GND.n1966 GND.n1933 19.3944
R12359 GND.n1934 GND.n1933 19.3944
R12360 GND.n1935 GND.n1934 19.3944
R12361 GND.n1941 GND.n1935 19.3944
R12362 GND.n1941 GND.n1940 19.3944
R12363 GND.n4133 GND.n1940 19.3944
R12364 GND.n4133 GND.n586 19.3944
R12365 GND.n5493 GND.n586 19.3944
R12366 GND.n5493 GND.n587 19.3944
R12367 GND.n589 GND.n587 19.3944
R12368 GND.n589 GND.n566 19.3944
R12369 GND.n5511 GND.n566 19.3944
R12370 GND.n5511 GND.n567 19.3944
R12371 GND.n567 GND.n554 19.3944
R12372 GND.n5570 GND.n554 19.3944
R12373 GND.n4198 GND.n4197 19.3944
R12374 GND.n4197 GND.n4196 19.3944
R12375 GND.n4196 GND.n1860 19.3944
R12376 GND.n4192 GND.n1860 19.3944
R12377 GND.n4192 GND.n4191 19.3944
R12378 GND.n4191 GND.n4190 19.3944
R12379 GND.n4190 GND.n1868 19.3944
R12380 GND.n4186 GND.n1868 19.3944
R12381 GND.n4186 GND.n4185 19.3944
R12382 GND.n4185 GND.n4184 19.3944
R12383 GND.n4184 GND.n1876 19.3944
R12384 GND.n4180 GND.n1876 19.3944
R12385 GND.n4180 GND.n4179 19.3944
R12386 GND.n4179 GND.n4178 19.3944
R12387 GND.n4178 GND.n1884 19.3944
R12388 GND.n4174 GND.n1884 19.3944
R12389 GND.n4174 GND.n4173 19.3944
R12390 GND.n4173 GND.n4172 19.3944
R12391 GND.n4172 GND.n1892 19.3944
R12392 GND.n4168 GND.n1892 19.3944
R12393 GND.n4168 GND.n4167 19.3944
R12394 GND.n4167 GND.n4166 19.3944
R12395 GND.n4166 GND.n1900 19.3944
R12396 GND.n4162 GND.n1900 19.3944
R12397 GND.n4162 GND.n4161 19.3944
R12398 GND.n4161 GND.n4160 19.3944
R12399 GND.n4160 GND.n1908 19.3944
R12400 GND.n4156 GND.n1908 19.3944
R12401 GND.n4156 GND.n4155 19.3944
R12402 GND.n4155 GND.n4154 19.3944
R12403 GND.n4154 GND.n1916 19.3944
R12404 GND.n4150 GND.n1916 19.3944
R12405 GND.n4150 GND.n4149 19.3944
R12406 GND.n4149 GND.n4148 19.3944
R12407 GND.n4148 GND.n1924 19.3944
R12408 GND.n4144 GND.n1924 19.3944
R12409 GND.n4144 GND.n4143 19.3944
R12410 GND.n4143 GND.n4142 19.3944
R12411 GND.n4142 GND.n1932 19.3944
R12412 GND.n4138 GND.n1932 19.3944
R12413 GND.n4138 GND.n4137 19.3944
R12414 GND.n4137 GND.n4136 19.3944
R12415 GND.n4136 GND.n592 19.3944
R12416 GND.n5489 GND.n592 19.3944
R12417 GND.n5491 GND.n5489 19.3944
R12418 GND.n5491 GND.n5490 19.3944
R12419 GND.n5490 GND.n570 19.3944
R12420 GND.n5506 GND.n570 19.3944
R12421 GND.n5509 GND.n5506 19.3944
R12422 GND.n5509 GND.n5508 19.3944
R12423 GND.n5508 GND.n552 19.3944
R12424 GND.n5572 GND.n552 19.3944
R12425 GND.n5628 GND.n496 19.3944
R12426 GND.n5624 GND.n496 19.3944
R12427 GND.n5624 GND.n5623 19.3944
R12428 GND.n5623 GND.n5622 19.3944
R12429 GND.n5622 GND.n503 19.3944
R12430 GND.n5618 GND.n503 19.3944
R12431 GND.n5618 GND.n5617 19.3944
R12432 GND.n5617 GND.n5616 19.3944
R12433 GND.n5616 GND.n509 19.3944
R12434 GND.n5612 GND.n509 19.3944
R12435 GND.n5612 GND.n5611 19.3944
R12436 GND.n5611 GND.n5610 19.3944
R12437 GND.n5610 GND.n515 19.3944
R12438 GND.n5606 GND.n515 19.3944
R12439 GND.n5606 GND.n5605 19.3944
R12440 GND.n5603 GND.n523 19.3944
R12441 GND.n5599 GND.n523 19.3944
R12442 GND.n5599 GND.n5598 19.3944
R12443 GND.n5598 GND.n5597 19.3944
R12444 GND.n5597 GND.n529 19.3944
R12445 GND.n5593 GND.n529 19.3944
R12446 GND.n5593 GND.n5592 19.3944
R12447 GND.n5592 GND.n5591 19.3944
R12448 GND.n5591 GND.n535 19.3944
R12449 GND.n5587 GND.n535 19.3944
R12450 GND.n5587 GND.n5586 19.3944
R12451 GND.n5586 GND.n5585 19.3944
R12452 GND.n5585 GND.n541 19.3944
R12453 GND.n5581 GND.n541 19.3944
R12454 GND.n5581 GND.n5580 19.3944
R12455 GND.n5580 GND.n5579 19.3944
R12456 GND.n4680 GND.n1156 19.3944
R12457 GND.n4676 GND.n1156 19.3944
R12458 GND.n4676 GND.n4675 19.3944
R12459 GND.n4675 GND.n4674 19.3944
R12460 GND.n4674 GND.n1164 19.3944
R12461 GND.n4670 GND.n1164 19.3944
R12462 GND.n4670 GND.n4669 19.3944
R12463 GND.n4669 GND.n4668 19.3944
R12464 GND.n4668 GND.n1172 19.3944
R12465 GND.n4664 GND.n1172 19.3944
R12466 GND.n4664 GND.n4663 19.3944
R12467 GND.n4663 GND.n4662 19.3944
R12468 GND.n4662 GND.n1180 19.3944
R12469 GND.n4658 GND.n1180 19.3944
R12470 GND.n4658 GND.n4657 19.3944
R12471 GND.n4657 GND.n4656 19.3944
R12472 GND.n4656 GND.n1188 19.3944
R12473 GND.n4652 GND.n1188 19.3944
R12474 GND.n4652 GND.n4651 19.3944
R12475 GND.n4651 GND.n4650 19.3944
R12476 GND.n4650 GND.n1196 19.3944
R12477 GND.n4646 GND.n1196 19.3944
R12478 GND.n4646 GND.n4645 19.3944
R12479 GND.n4645 GND.n4644 19.3944
R12480 GND.n4644 GND.n1204 19.3944
R12481 GND.n4640 GND.n1204 19.3944
R12482 GND.n4640 GND.n4639 19.3944
R12483 GND.n4639 GND.n4638 19.3944
R12484 GND.n4638 GND.n1212 19.3944
R12485 GND.n4634 GND.n1212 19.3944
R12486 GND.n4634 GND.n4633 19.3944
R12487 GND.n4633 GND.n4632 19.3944
R12488 GND.n4632 GND.n1220 19.3944
R12489 GND.n4628 GND.n1220 19.3944
R12490 GND.n4628 GND.n4627 19.3944
R12491 GND.n4627 GND.n4626 19.3944
R12492 GND.n4626 GND.n1228 19.3944
R12493 GND.n4622 GND.n1228 19.3944
R12494 GND.n4622 GND.n4621 19.3944
R12495 GND.n4621 GND.n4620 19.3944
R12496 GND.n4620 GND.n1236 19.3944
R12497 GND.n4616 GND.n1236 19.3944
R12498 GND.n4616 GND.n4615 19.3944
R12499 GND.n4615 GND.n4614 19.3944
R12500 GND.n4614 GND.n1244 19.3944
R12501 GND.n4610 GND.n1244 19.3944
R12502 GND.n4610 GND.n4609 19.3944
R12503 GND.n4609 GND.n4608 19.3944
R12504 GND.n4608 GND.n1252 19.3944
R12505 GND.n4604 GND.n1252 19.3944
R12506 GND.n4604 GND.n4603 19.3944
R12507 GND.n4603 GND.n4602 19.3944
R12508 GND.n4595 GND.n4594 19.3944
R12509 GND.n4594 GND.n4593 19.3944
R12510 GND.n4593 GND.n1272 19.3944
R12511 GND.n4589 GND.n1272 19.3944
R12512 GND.n4589 GND.n4588 19.3944
R12513 GND.n4588 GND.n4587 19.3944
R12514 GND.n4587 GND.n1277 19.3944
R12515 GND.n4583 GND.n1277 19.3944
R12516 GND.n4583 GND.n4582 19.3944
R12517 GND.n4582 GND.n4581 19.3944
R12518 GND.n4581 GND.n1282 19.3944
R12519 GND.n4577 GND.n1282 19.3944
R12520 GND.n4577 GND.n4576 19.3944
R12521 GND.n4574 GND.n1292 19.3944
R12522 GND.n4570 GND.n1292 19.3944
R12523 GND.n4570 GND.n4569 19.3944
R12524 GND.n4569 GND.n4568 19.3944
R12525 GND.n4568 GND.n1297 19.3944
R12526 GND.n4564 GND.n1297 19.3944
R12527 GND.n4564 GND.n4563 19.3944
R12528 GND.n4563 GND.n4562 19.3944
R12529 GND.n4562 GND.n1302 19.3944
R12530 GND.n4558 GND.n1302 19.3944
R12531 GND.n4558 GND.n4557 19.3944
R12532 GND.n4557 GND.n4556 19.3944
R12533 GND.n4556 GND.n1307 19.3944
R12534 GND.n4552 GND.n1307 19.3944
R12535 GND.n4552 GND.n4551 19.3944
R12536 GND.n4551 GND.n4550 19.3944
R12537 GND.n2582 GND.n2581 19.3944
R12538 GND.n2581 GND.n2580 19.3944
R12539 GND.n2580 GND.n2502 19.3944
R12540 GND.n2631 GND.n2502 19.3944
R12541 GND.n2631 GND.n2499 19.3944
R12542 GND.n2636 GND.n2499 19.3944
R12543 GND.n2636 GND.n2500 19.3944
R12544 GND.n2500 GND.n2479 19.3944
R12545 GND.n2656 GND.n2479 19.3944
R12546 GND.n2656 GND.n2476 19.3944
R12547 GND.n2661 GND.n2476 19.3944
R12548 GND.n2661 GND.n2477 19.3944
R12549 GND.n2477 GND.n2457 19.3944
R12550 GND.n2681 GND.n2457 19.3944
R12551 GND.n2681 GND.n2454 19.3944
R12552 GND.n2700 GND.n2454 19.3944
R12553 GND.n2700 GND.n2455 19.3944
R12554 GND.n2696 GND.n2455 19.3944
R12555 GND.n2696 GND.n2695 19.3944
R12556 GND.n2695 GND.n2694 19.3944
R12557 GND.n2694 GND.n2424 19.3944
R12558 GND.n2731 GND.n2424 19.3944
R12559 GND.n2732 GND.n2731 19.3944
R12560 GND.n2732 GND.n2422 19.3944
R12561 GND.n2736 GND.n2422 19.3944
R12562 GND.n2739 GND.n2736 19.3944
R12563 GND.n2740 GND.n2739 19.3944
R12564 GND.n2740 GND.n2420 19.3944
R12565 GND.n2744 GND.n2420 19.3944
R12566 GND.n2744 GND.n2371 19.3944
R12567 GND.n2838 GND.n2371 19.3944
R12568 GND.n2838 GND.n2368 19.3944
R12569 GND.n2843 GND.n2368 19.3944
R12570 GND.n2843 GND.n2369 19.3944
R12571 GND.n2369 GND.n2351 19.3944
R12572 GND.n2863 GND.n2351 19.3944
R12573 GND.n2863 GND.n2348 19.3944
R12574 GND.n2868 GND.n2348 19.3944
R12575 GND.n2868 GND.n2349 19.3944
R12576 GND.n2349 GND.n2331 19.3944
R12577 GND.n2888 GND.n2331 19.3944
R12578 GND.n2888 GND.n2328 19.3944
R12579 GND.n2896 GND.n2328 19.3944
R12580 GND.n2896 GND.n2329 19.3944
R12581 GND.n2892 GND.n2329 19.3944
R12582 GND.n2892 GND.n2303 19.3944
R12583 GND.n2937 GND.n2303 19.3944
R12584 GND.n2937 GND.n2304 19.3944
R12585 GND.n2933 GND.n2304 19.3944
R12586 GND.n2933 GND.n2287 19.3944
R12587 GND.n2957 GND.n2287 19.3944
R12588 GND.n2958 GND.n2957 19.3944
R12589 GND.n4543 GND.n4542 19.3944
R12590 GND.n4542 GND.n4541 19.3944
R12591 GND.n4541 GND.n1319 19.3944
R12592 GND.n1380 GND.n1319 19.3944
R12593 GND.n1380 GND.n1345 19.3944
R12594 GND.n4529 GND.n1345 19.3944
R12595 GND.n4529 GND.n4528 19.3944
R12596 GND.n4528 GND.n1348 19.3944
R12597 GND.n4521 GND.n1348 19.3944
R12598 GND.n4521 GND.n4520 19.3944
R12599 GND.n4520 GND.n1356 19.3944
R12600 GND.n4513 GND.n1356 19.3944
R12601 GND.n4513 GND.n4512 19.3944
R12602 GND.n4512 GND.n1366 19.3944
R12603 GND.n2612 GND.n2611 19.3944
R12604 GND.n2611 GND.n2557 19.3944
R12605 GND.n2607 GND.n2557 19.3944
R12606 GND.n2607 GND.n2606 19.3944
R12607 GND.n2606 GND.n2605 19.3944
R12608 GND.n2605 GND.n2563 19.3944
R12609 GND.n2601 GND.n2563 19.3944
R12610 GND.n2601 GND.n2600 19.3944
R12611 GND.n2600 GND.n2599 19.3944
R12612 GND.n2599 GND.n2569 19.3944
R12613 GND.n2595 GND.n2569 19.3944
R12614 GND.n2595 GND.n2594 19.3944
R12615 GND.n2594 GND.n2593 19.3944
R12616 GND.n2593 GND.n2575 19.3944
R12617 GND.n1158 GND.n1157 19.3944
R12618 GND.n1159 GND.n1158 19.3944
R12619 GND.n2616 GND.n1159 19.3944
R12620 GND.n2616 GND.n1165 19.3944
R12621 GND.n1166 GND.n1165 19.3944
R12622 GND.n1167 GND.n1166 19.3944
R12623 GND.n2642 GND.n1167 19.3944
R12624 GND.n2642 GND.n1173 19.3944
R12625 GND.n1174 GND.n1173 19.3944
R12626 GND.n1175 GND.n1174 19.3944
R12627 GND.n2473 GND.n1175 19.3944
R12628 GND.n2473 GND.n1181 19.3944
R12629 GND.n1182 GND.n1181 19.3944
R12630 GND.n1183 GND.n1182 19.3944
R12631 GND.n2450 GND.n1183 19.3944
R12632 GND.n2450 GND.n1189 19.3944
R12633 GND.n1190 GND.n1189 19.3944
R12634 GND.n1191 GND.n1190 19.3944
R12635 GND.n2437 GND.n1191 19.3944
R12636 GND.n2437 GND.n1197 19.3944
R12637 GND.n1198 GND.n1197 19.3944
R12638 GND.n1199 GND.n1198 19.3944
R12639 GND.n2824 GND.n1199 19.3944
R12640 GND.n2824 GND.n1205 19.3944
R12641 GND.n1206 GND.n1205 19.3944
R12642 GND.n1207 GND.n1206 19.3944
R12643 GND.n2407 GND.n1207 19.3944
R12644 GND.n2407 GND.n1213 19.3944
R12645 GND.n1214 GND.n1213 19.3944
R12646 GND.n1215 GND.n1214 19.3944
R12647 GND.n2375 GND.n1215 19.3944
R12648 GND.n2375 GND.n1221 19.3944
R12649 GND.n1222 GND.n1221 19.3944
R12650 GND.n1223 GND.n1222 19.3944
R12651 GND.n2847 GND.n1223 19.3944
R12652 GND.n2847 GND.n1229 19.3944
R12653 GND.n1230 GND.n1229 19.3944
R12654 GND.n1231 GND.n1230 19.3944
R12655 GND.n2874 GND.n1231 19.3944
R12656 GND.n2874 GND.n1237 19.3944
R12657 GND.n1238 GND.n1237 19.3944
R12658 GND.n1239 GND.n1238 19.3944
R12659 GND.n2326 GND.n1239 19.3944
R12660 GND.n2326 GND.n1245 19.3944
R12661 GND.n1246 GND.n1245 19.3944
R12662 GND.n1247 GND.n1246 19.3944
R12663 GND.n2300 GND.n1247 19.3944
R12664 GND.n2300 GND.n1253 19.3944
R12665 GND.n1254 GND.n1253 19.3944
R12666 GND.n1255 GND.n1254 19.3944
R12667 GND.n2953 GND.n1255 19.3944
R12668 GND.n2953 GND.n2952 19.3944
R12669 GND.n3004 GND.n3003 19.3944
R12670 GND.n3007 GND.n3004 19.3944
R12671 GND.n3007 GND.n2273 19.3944
R12672 GND.n3011 GND.n2273 19.3944
R12673 GND.n3014 GND.n3011 19.3944
R12674 GND.n3015 GND.n3014 19.3944
R12675 GND.n3015 GND.n2271 19.3944
R12676 GND.n3019 GND.n2271 19.3944
R12677 GND.n3020 GND.n3019 19.3944
R12678 GND.n3023 GND.n3020 19.3944
R12679 GND.n3023 GND.n2266 19.3944
R12680 GND.n3033 GND.n2266 19.3944
R12681 GND.n3033 GND.n2267 19.3944
R12682 GND.n3029 GND.n2267 19.3944
R12683 GND.n3029 GND.n3028 19.3944
R12684 GND.n3028 GND.n2238 19.3944
R12685 GND.n3250 GND.n2238 19.3944
R12686 GND.n3250 GND.n2235 19.3944
R12687 GND.n3270 GND.n2235 19.3944
R12688 GND.n3270 GND.n2236 19.3944
R12689 GND.n3266 GND.n2236 19.3944
R12690 GND.n3266 GND.n3265 19.3944
R12691 GND.n3265 GND.n3264 19.3944
R12692 GND.n3264 GND.n3258 19.3944
R12693 GND.n3260 GND.n3258 19.3944
R12694 GND.n3260 GND.n2214 19.3944
R12695 GND.n3322 GND.n2214 19.3944
R12696 GND.n3322 GND.n2211 19.3944
R12697 GND.n3347 GND.n2211 19.3944
R12698 GND.n3347 GND.n2212 19.3944
R12699 GND.n3343 GND.n2212 19.3944
R12700 GND.n3343 GND.n3342 19.3944
R12701 GND.n3342 GND.n3341 19.3944
R12702 GND.n3341 GND.n3330 19.3944
R12703 GND.n3337 GND.n3330 19.3944
R12704 GND.n3337 GND.n3336 19.3944
R12705 GND.n3336 GND.n3335 19.3944
R12706 GND.n3335 GND.n2197 19.3944
R12707 GND.n2197 GND.n2196 19.3944
R12708 GND.n3398 GND.n2196 19.3944
R12709 GND.n3398 GND.n2193 19.3944
R12710 GND.n3406 GND.n2193 19.3944
R12711 GND.n3406 GND.n2194 19.3944
R12712 GND.n3402 GND.n2194 19.3944
R12713 GND.n3402 GND.n2184 19.3944
R12714 GND.n3443 GND.n2184 19.3944
R12715 GND.n3443 GND.n2182 19.3944
R12716 GND.n3448 GND.n2182 19.3944
R12717 GND.n3448 GND.n2176 19.3944
R12718 GND.n3782 GND.n2176 19.3944
R12719 GND.n3783 GND.n3782 19.3944
R12720 GND.n3783 GND.n2174 19.3944
R12721 GND.n3787 GND.n2174 19.3944
R12722 GND.n3788 GND.n3787 19.3944
R12723 GND.n3791 GND.n3788 19.3944
R12724 GND.n3791 GND.n2170 19.3944
R12725 GND.n3795 GND.n2170 19.3944
R12726 GND.n3796 GND.n3795 19.3944
R12727 GND.n3799 GND.n3796 19.3944
R12728 GND.n3799 GND.n2168 19.3944
R12729 GND.n3803 GND.n2168 19.3944
R12730 GND.n3807 GND.n3803 19.3944
R12731 GND.n3808 GND.n3807 19.3944
R12732 GND.n3808 GND.n2166 19.3944
R12733 GND.n3812 GND.n2166 19.3944
R12734 GND.n4252 GND.n1778 19.3944
R12735 GND.n4245 GND.n1778 19.3944
R12736 GND.n4245 GND.n4244 19.3944
R12737 GND.n4244 GND.n1788 19.3944
R12738 GND.n4237 GND.n1788 19.3944
R12739 GND.n4237 GND.n4236 19.3944
R12740 GND.n4236 GND.n1798 19.3944
R12741 GND.n4229 GND.n1798 19.3944
R12742 GND.n4229 GND.n4228 19.3944
R12743 GND.n4228 GND.n1806 19.3944
R12744 GND.n4221 GND.n1806 19.3944
R12745 GND.n4221 GND.n4220 19.3944
R12746 GND.n4220 GND.n1818 19.3944
R12747 GND.n2142 GND.n1818 19.3944
R12748 GND.n3835 GND.n2142 19.3944
R12749 GND.n3835 GND.n3834 19.3944
R12750 GND.n3834 GND.n3833 19.3944
R12751 GND.n3833 GND.n2147 19.3944
R12752 GND.n3829 GND.n2147 19.3944
R12753 GND.n3829 GND.n3828 19.3944
R12754 GND.n3828 GND.n3827 19.3944
R12755 GND.n3827 GND.n2153 19.3944
R12756 GND.n3823 GND.n2153 19.3944
R12757 GND.n3823 GND.n3822 19.3944
R12758 GND.n3820 GND.n2161 19.3944
R12759 GND.n3816 GND.n2161 19.3944
R12760 GND.n3816 GND.n3815 19.3944
R12761 GND.n2995 GND.n2276 19.3944
R12762 GND.n2998 GND.n2995 19.3944
R12763 GND.n3000 GND.n2998 19.3944
R12764 GND.n4537 GND.n1322 19.3944
R12765 GND.n4532 GND.n1322 19.3944
R12766 GND.n4532 GND.n1341 19.3944
R12767 GND.n4525 GND.n1341 19.3944
R12768 GND.n4525 GND.n4524 19.3944
R12769 GND.n4524 GND.n1352 19.3944
R12770 GND.n4517 GND.n1352 19.3944
R12771 GND.n4517 GND.n4516 19.3944
R12772 GND.n4516 GND.n1362 19.3944
R12773 GND.n4509 GND.n1362 19.3944
R12774 GND.n4509 GND.n4508 19.3944
R12775 GND.n4508 GND.n1370 19.3944
R12776 GND.n2284 GND.n1370 19.3944
R12777 GND.n2962 GND.n2284 19.3944
R12778 GND.n2965 GND.n2962 19.3944
R12779 GND.n2968 GND.n2965 19.3944
R12780 GND.n2968 GND.n2280 19.3944
R12781 GND.n2972 GND.n2280 19.3944
R12782 GND.n2975 GND.n2972 19.3944
R12783 GND.n2978 GND.n2975 19.3944
R12784 GND.n2978 GND.n2278 19.3944
R12785 GND.n2982 GND.n2278 19.3944
R12786 GND.n2985 GND.n2982 19.3944
R12787 GND.n2991 GND.n2985 19.3944
R12788 GND.n4462 GND.n1405 19.3944
R12789 GND.n4462 GND.n4461 19.3944
R12790 GND.n4461 GND.n4460 19.3944
R12791 GND.n4460 GND.n1410 19.3944
R12792 GND.n1437 GND.n1410 19.3944
R12793 GND.n4448 GND.n1437 19.3944
R12794 GND.n4448 GND.n4447 19.3944
R12795 GND.n4447 GND.n4446 19.3944
R12796 GND.n4446 GND.n1443 19.3944
R12797 GND.n1464 GND.n1443 19.3944
R12798 GND.n4434 GND.n1464 19.3944
R12799 GND.n4434 GND.n4433 19.3944
R12800 GND.n4433 GND.n4432 19.3944
R12801 GND.n4432 GND.n1470 19.3944
R12802 GND.n3236 GND.n1470 19.3944
R12803 GND.n3245 GND.n3236 19.3944
R12804 GND.n3245 GND.n3244 19.3944
R12805 GND.n3244 GND.n3243 19.3944
R12806 GND.n3243 GND.n2227 19.3944
R12807 GND.n2227 GND.n2225 19.3944
R12808 GND.n3276 GND.n2225 19.3944
R12809 GND.n3276 GND.n2223 19.3944
R12810 GND.n3289 GND.n2223 19.3944
R12811 GND.n3289 GND.n3288 19.3944
R12812 GND.n3288 GND.n3287 19.3944
R12813 GND.n3287 GND.n3284 19.3944
R12814 GND.n3284 GND.n1544 19.3944
R12815 GND.n4378 GND.n1544 19.3944
R12816 GND.n4378 GND.n4377 19.3944
R12817 GND.n4377 GND.n4376 19.3944
R12818 GND.n4376 GND.n1548 19.3944
R12819 GND.n1592 GND.n1548 19.3944
R12820 GND.n1595 GND.n1592 19.3944
R12821 GND.n1595 GND.n1589 19.3944
R12822 GND.n4350 GND.n1589 19.3944
R12823 GND.n4350 GND.n4349 19.3944
R12824 GND.n4349 GND.n4348 19.3944
R12825 GND.n4348 GND.n1601 19.3944
R12826 GND.n1635 GND.n1601 19.3944
R12827 GND.n1635 GND.n1632 19.3944
R12828 GND.n4330 GND.n1632 19.3944
R12829 GND.n4330 GND.n4329 19.3944
R12830 GND.n4329 GND.n4328 19.3944
R12831 GND.n4328 GND.n1641 19.3944
R12832 GND.n1670 GND.n1641 19.3944
R12833 GND.n1670 GND.n1667 19.3944
R12834 GND.n4309 GND.n1667 19.3944
R12835 GND.n4309 GND.n4308 19.3944
R12836 GND.n4308 GND.n4307 19.3944
R12837 GND.n4307 GND.n1676 19.3944
R12838 GND.n4295 GND.n1676 19.3944
R12839 GND.n4295 GND.n4294 19.3944
R12840 GND.n4294 GND.n4293 19.3944
R12841 GND.n4293 GND.n1694 19.3944
R12842 GND.n1712 GND.n1694 19.3944
R12843 GND.n4281 GND.n1712 19.3944
R12844 GND.n4281 GND.n4280 19.3944
R12845 GND.n4280 GND.n4279 19.3944
R12846 GND.n4279 GND.n1718 19.3944
R12847 GND.n1739 GND.n1718 19.3944
R12848 GND.n4267 GND.n1739 19.3944
R12849 GND.n4267 GND.n4266 19.3944
R12850 GND.n4266 GND.n4265 19.3944
R12851 GND.n4265 GND.n1745 19.3944
R12852 GND.n4206 GND.n1745 19.3944
R12853 GND.n5315 GND.n698 19.3944
R12854 GND.n5319 GND.n698 19.3944
R12855 GND.n5319 GND.n694 19.3944
R12856 GND.n5325 GND.n694 19.3944
R12857 GND.n5325 GND.n692 19.3944
R12858 GND.n5329 GND.n692 19.3944
R12859 GND.n5329 GND.n688 19.3944
R12860 GND.n5335 GND.n688 19.3944
R12861 GND.n5335 GND.n686 19.3944
R12862 GND.n5339 GND.n686 19.3944
R12863 GND.n5339 GND.n682 19.3944
R12864 GND.n5345 GND.n682 19.3944
R12865 GND.n5345 GND.n680 19.3944
R12866 GND.n5349 GND.n680 19.3944
R12867 GND.n5349 GND.n676 19.3944
R12868 GND.n5355 GND.n676 19.3944
R12869 GND.n5355 GND.n674 19.3944
R12870 GND.n5359 GND.n674 19.3944
R12871 GND.n5359 GND.n670 19.3944
R12872 GND.n5365 GND.n670 19.3944
R12873 GND.n5365 GND.n668 19.3944
R12874 GND.n5369 GND.n668 19.3944
R12875 GND.n5369 GND.n664 19.3944
R12876 GND.n5375 GND.n664 19.3944
R12877 GND.n5375 GND.n662 19.3944
R12878 GND.n5379 GND.n662 19.3944
R12879 GND.n5379 GND.n658 19.3944
R12880 GND.n5385 GND.n658 19.3944
R12881 GND.n5385 GND.n656 19.3944
R12882 GND.n5389 GND.n656 19.3944
R12883 GND.n5389 GND.n652 19.3944
R12884 GND.n5395 GND.n652 19.3944
R12885 GND.n5395 GND.n650 19.3944
R12886 GND.n5399 GND.n650 19.3944
R12887 GND.n5399 GND.n646 19.3944
R12888 GND.n5405 GND.n646 19.3944
R12889 GND.n5405 GND.n644 19.3944
R12890 GND.n5409 GND.n644 19.3944
R12891 GND.n5409 GND.n640 19.3944
R12892 GND.n5415 GND.n640 19.3944
R12893 GND.n5415 GND.n638 19.3944
R12894 GND.n5419 GND.n638 19.3944
R12895 GND.n5419 GND.n634 19.3944
R12896 GND.n5425 GND.n634 19.3944
R12897 GND.n5425 GND.n632 19.3944
R12898 GND.n5429 GND.n632 19.3944
R12899 GND.n5429 GND.n628 19.3944
R12900 GND.n5435 GND.n628 19.3944
R12901 GND.n5435 GND.n626 19.3944
R12902 GND.n5439 GND.n626 19.3944
R12903 GND.n5439 GND.n622 19.3944
R12904 GND.n5445 GND.n622 19.3944
R12905 GND.n5445 GND.n620 19.3944
R12906 GND.n5449 GND.n620 19.3944
R12907 GND.n5449 GND.n616 19.3944
R12908 GND.n5455 GND.n616 19.3944
R12909 GND.n5455 GND.n614 19.3944
R12910 GND.n5459 GND.n614 19.3944
R12911 GND.n5459 GND.n610 19.3944
R12912 GND.n5465 GND.n610 19.3944
R12913 GND.n5465 GND.n608 19.3944
R12914 GND.n5469 GND.n608 19.3944
R12915 GND.n5469 GND.n604 19.3944
R12916 GND.n5475 GND.n604 19.3944
R12917 GND.n5475 GND.n602 19.3944
R12918 GND.n5479 GND.n602 19.3944
R12919 GND.n4888 GND.n955 19.3944
R12920 GND.n4888 GND.n951 19.3944
R12921 GND.n4894 GND.n951 19.3944
R12922 GND.n4894 GND.n949 19.3944
R12923 GND.n4898 GND.n949 19.3944
R12924 GND.n4898 GND.n945 19.3944
R12925 GND.n4904 GND.n945 19.3944
R12926 GND.n4904 GND.n943 19.3944
R12927 GND.n4908 GND.n943 19.3944
R12928 GND.n4908 GND.n939 19.3944
R12929 GND.n4914 GND.n939 19.3944
R12930 GND.n4914 GND.n937 19.3944
R12931 GND.n4918 GND.n937 19.3944
R12932 GND.n4918 GND.n933 19.3944
R12933 GND.n4924 GND.n933 19.3944
R12934 GND.n4924 GND.n931 19.3944
R12935 GND.n4928 GND.n931 19.3944
R12936 GND.n4928 GND.n927 19.3944
R12937 GND.n4934 GND.n927 19.3944
R12938 GND.n4934 GND.n925 19.3944
R12939 GND.n4938 GND.n925 19.3944
R12940 GND.n4938 GND.n921 19.3944
R12941 GND.n4944 GND.n921 19.3944
R12942 GND.n4944 GND.n919 19.3944
R12943 GND.n4948 GND.n919 19.3944
R12944 GND.n4948 GND.n915 19.3944
R12945 GND.n4954 GND.n915 19.3944
R12946 GND.n4954 GND.n913 19.3944
R12947 GND.n4958 GND.n913 19.3944
R12948 GND.n4958 GND.n909 19.3944
R12949 GND.n4964 GND.n909 19.3944
R12950 GND.n4964 GND.n907 19.3944
R12951 GND.n4968 GND.n907 19.3944
R12952 GND.n4968 GND.n903 19.3944
R12953 GND.n4974 GND.n903 19.3944
R12954 GND.n4974 GND.n901 19.3944
R12955 GND.n4978 GND.n901 19.3944
R12956 GND.n4978 GND.n897 19.3944
R12957 GND.n4984 GND.n897 19.3944
R12958 GND.n4984 GND.n895 19.3944
R12959 GND.n4988 GND.n895 19.3944
R12960 GND.n4988 GND.n891 19.3944
R12961 GND.n4994 GND.n891 19.3944
R12962 GND.n4994 GND.n889 19.3944
R12963 GND.n4998 GND.n889 19.3944
R12964 GND.n4998 GND.n885 19.3944
R12965 GND.n5004 GND.n885 19.3944
R12966 GND.n5004 GND.n883 19.3944
R12967 GND.n5008 GND.n883 19.3944
R12968 GND.n5008 GND.n879 19.3944
R12969 GND.n5014 GND.n879 19.3944
R12970 GND.n5014 GND.n877 19.3944
R12971 GND.n5018 GND.n877 19.3944
R12972 GND.n5018 GND.n873 19.3944
R12973 GND.n5024 GND.n873 19.3944
R12974 GND.n5024 GND.n871 19.3944
R12975 GND.n5028 GND.n871 19.3944
R12976 GND.n5028 GND.n867 19.3944
R12977 GND.n5034 GND.n867 19.3944
R12978 GND.n5034 GND.n865 19.3944
R12979 GND.n5038 GND.n865 19.3944
R12980 GND.n5038 GND.n861 19.3944
R12981 GND.n5044 GND.n861 19.3944
R12982 GND.n5044 GND.n859 19.3944
R12983 GND.n5048 GND.n859 19.3944
R12984 GND.n5048 GND.n855 19.3944
R12985 GND.n5054 GND.n855 19.3944
R12986 GND.n5054 GND.n853 19.3944
R12987 GND.n5058 GND.n853 19.3944
R12988 GND.n5058 GND.n849 19.3944
R12989 GND.n5064 GND.n849 19.3944
R12990 GND.n5064 GND.n847 19.3944
R12991 GND.n5068 GND.n847 19.3944
R12992 GND.n5068 GND.n843 19.3944
R12993 GND.n5074 GND.n843 19.3944
R12994 GND.n5074 GND.n841 19.3944
R12995 GND.n5078 GND.n841 19.3944
R12996 GND.n5078 GND.n837 19.3944
R12997 GND.n5084 GND.n837 19.3944
R12998 GND.n5084 GND.n835 19.3944
R12999 GND.n5088 GND.n835 19.3944
R13000 GND.n5088 GND.n831 19.3944
R13001 GND.n5094 GND.n831 19.3944
R13002 GND.n5094 GND.n829 19.3944
R13003 GND.n5098 GND.n829 19.3944
R13004 GND.n5098 GND.n825 19.3944
R13005 GND.n5104 GND.n825 19.3944
R13006 GND.n5104 GND.n823 19.3944
R13007 GND.n5108 GND.n823 19.3944
R13008 GND.n5108 GND.n819 19.3944
R13009 GND.n5114 GND.n819 19.3944
R13010 GND.n5114 GND.n817 19.3944
R13011 GND.n5118 GND.n817 19.3944
R13012 GND.n5118 GND.n813 19.3944
R13013 GND.n5124 GND.n813 19.3944
R13014 GND.n5124 GND.n811 19.3944
R13015 GND.n5128 GND.n811 19.3944
R13016 GND.n5128 GND.n807 19.3944
R13017 GND.n5134 GND.n807 19.3944
R13018 GND.n5134 GND.n805 19.3944
R13019 GND.n5138 GND.n805 19.3944
R13020 GND.n5138 GND.n801 19.3944
R13021 GND.n5144 GND.n801 19.3944
R13022 GND.n5144 GND.n799 19.3944
R13023 GND.n5148 GND.n799 19.3944
R13024 GND.n5148 GND.n795 19.3944
R13025 GND.n5154 GND.n795 19.3944
R13026 GND.n5154 GND.n793 19.3944
R13027 GND.n5158 GND.n793 19.3944
R13028 GND.n5158 GND.n789 19.3944
R13029 GND.n5164 GND.n789 19.3944
R13030 GND.n5164 GND.n787 19.3944
R13031 GND.n5168 GND.n787 19.3944
R13032 GND.n5168 GND.n783 19.3944
R13033 GND.n5174 GND.n783 19.3944
R13034 GND.n5174 GND.n781 19.3944
R13035 GND.n5178 GND.n781 19.3944
R13036 GND.n5178 GND.n777 19.3944
R13037 GND.n5184 GND.n777 19.3944
R13038 GND.n5184 GND.n775 19.3944
R13039 GND.n5188 GND.n775 19.3944
R13040 GND.n5188 GND.n771 19.3944
R13041 GND.n5194 GND.n771 19.3944
R13042 GND.n5194 GND.n769 19.3944
R13043 GND.n5198 GND.n769 19.3944
R13044 GND.n5198 GND.n765 19.3944
R13045 GND.n5204 GND.n765 19.3944
R13046 GND.n5204 GND.n763 19.3944
R13047 GND.n5208 GND.n763 19.3944
R13048 GND.n5208 GND.n759 19.3944
R13049 GND.n5214 GND.n759 19.3944
R13050 GND.n5214 GND.n757 19.3944
R13051 GND.n5218 GND.n757 19.3944
R13052 GND.n5218 GND.n753 19.3944
R13053 GND.n5224 GND.n753 19.3944
R13054 GND.n5224 GND.n751 19.3944
R13055 GND.n5228 GND.n751 19.3944
R13056 GND.n5228 GND.n747 19.3944
R13057 GND.n5234 GND.n747 19.3944
R13058 GND.n5234 GND.n745 19.3944
R13059 GND.n5238 GND.n745 19.3944
R13060 GND.n5238 GND.n741 19.3944
R13061 GND.n5244 GND.n741 19.3944
R13062 GND.n5244 GND.n739 19.3944
R13063 GND.n5248 GND.n739 19.3944
R13064 GND.n5248 GND.n735 19.3944
R13065 GND.n5254 GND.n735 19.3944
R13066 GND.n5254 GND.n733 19.3944
R13067 GND.n5258 GND.n733 19.3944
R13068 GND.n5258 GND.n729 19.3944
R13069 GND.n5264 GND.n729 19.3944
R13070 GND.n5264 GND.n727 19.3944
R13071 GND.n5268 GND.n727 19.3944
R13072 GND.n5268 GND.n723 19.3944
R13073 GND.n5274 GND.n723 19.3944
R13074 GND.n5274 GND.n721 19.3944
R13075 GND.n5278 GND.n721 19.3944
R13076 GND.n5278 GND.n717 19.3944
R13077 GND.n5284 GND.n717 19.3944
R13078 GND.n5284 GND.n715 19.3944
R13079 GND.n5288 GND.n715 19.3944
R13080 GND.n5288 GND.n711 19.3944
R13081 GND.n5294 GND.n711 19.3944
R13082 GND.n5294 GND.n709 19.3944
R13083 GND.n5298 GND.n709 19.3944
R13084 GND.n5298 GND.n705 19.3944
R13085 GND.n5304 GND.n705 19.3944
R13086 GND.n5304 GND.n703 19.3944
R13087 GND.n5309 GND.n703 19.3944
R13088 GND.n5309 GND.n5308 19.3944
R13089 GND.n3591 GND.n3586 19.3944
R13090 GND.n3597 GND.n3586 19.3944
R13091 GND.n3598 GND.n3597 19.3944
R13092 GND.n3601 GND.n3598 19.3944
R13093 GND.n3601 GND.n3584 19.3944
R13094 GND.n3607 GND.n3584 19.3944
R13095 GND.n3608 GND.n3607 19.3944
R13096 GND.n3611 GND.n3608 19.3944
R13097 GND.n3611 GND.n3582 19.3944
R13098 GND.n3617 GND.n3582 19.3944
R13099 GND.n3618 GND.n3617 19.3944
R13100 GND.n3621 GND.n3618 19.3944
R13101 GND.n3621 GND.n3579 19.3944
R13102 GND.n3684 GND.n3681 19.3944
R13103 GND.n3681 GND.n3680 19.3944
R13104 GND.n3680 GND.n3677 19.3944
R13105 GND.n3677 GND.n3676 19.3944
R13106 GND.n3676 GND.n3673 19.3944
R13107 GND.n3673 GND.n3672 19.3944
R13108 GND.n3672 GND.n3669 19.3944
R13109 GND.n3669 GND.n3668 19.3944
R13110 GND.n3668 GND.n3665 19.3944
R13111 GND.n3665 GND.n3664 19.3944
R13112 GND.n3664 GND.n3661 19.3944
R13113 GND.n3661 GND.n3660 19.3944
R13114 GND.n3660 GND.n3657 19.3944
R13115 GND.n3657 GND.n3656 19.3944
R13116 GND.n3656 GND.n3653 19.3944
R13117 GND.n3653 GND.n3652 19.3944
R13118 GND.n3588 GND.n2110 19.3944
R13119 GND.n3895 GND.n2110 19.3944
R13120 GND.n3895 GND.n2108 19.3944
R13121 GND.n3901 GND.n2108 19.3944
R13122 GND.n3901 GND.n3900 19.3944
R13123 GND.n3900 GND.n2087 19.3944
R13124 GND.n3919 GND.n2087 19.3944
R13125 GND.n3919 GND.n2085 19.3944
R13126 GND.n3925 GND.n2085 19.3944
R13127 GND.n3925 GND.n3924 19.3944
R13128 GND.n3924 GND.n2066 19.3944
R13129 GND.n3944 GND.n2066 19.3944
R13130 GND.n3944 GND.n2064 19.3944
R13131 GND.n3950 GND.n2064 19.3944
R13132 GND.n3950 GND.n3949 19.3944
R13133 GND.n3949 GND.n2033 19.3944
R13134 GND.n3984 GND.n2033 19.3944
R13135 GND.n3984 GND.n2031 19.3944
R13136 GND.n3988 GND.n2031 19.3944
R13137 GND.n3989 GND.n3988 19.3944
R13138 GND.n3989 GND.n1999 19.3944
R13139 GND.n4063 GND.n4062 19.3944
R13140 GND.n4018 GND.n4017 19.3944
R13141 GND.n4046 GND.n4045 19.3944
R13142 GND.n4023 GND.n4022 19.3944
R13143 GND.n4030 GND.n1993 19.3944
R13144 GND.n4069 GND.n1993 19.3944
R13145 GND.n4069 GND.n4068 19.3944
R13146 GND.n4068 GND.n1972 19.3944
R13147 GND.n4089 GND.n1972 19.3944
R13148 GND.n4089 GND.n1970 19.3944
R13149 GND.n4095 GND.n1970 19.3944
R13150 GND.n4095 GND.n4094 19.3944
R13151 GND.n4094 GND.n1949 19.3944
R13152 GND.n4122 GND.n1949 19.3944
R13153 GND.n4122 GND.n1947 19.3944
R13154 GND.n4128 GND.n1947 19.3944
R13155 GND.n4128 GND.n4127 19.3944
R13156 GND.n4127 GND.n578 19.3944
R13157 GND.n5497 GND.n578 19.3944
R13158 GND.n5497 GND.n576 19.3944
R13159 GND.n5501 GND.n576 19.3944
R13160 GND.n5501 GND.n560 19.3944
R13161 GND.n5515 GND.n560 19.3944
R13162 GND.n5515 GND.n558 19.3944
R13163 GND.n5520 GND.n558 19.3944
R13164 GND.n5520 GND.n5519 19.3944
R13165 GND.n2537 GND.n2536 19.3944
R13166 GND.n2536 GND.n2508 19.3944
R13167 GND.n2532 GND.n2508 19.3944
R13168 GND.n2532 GND.n2531 19.3944
R13169 GND.n2531 GND.n2530 19.3944
R13170 GND.n2530 GND.n2514 19.3944
R13171 GND.n2526 GND.n2514 19.3944
R13172 GND.n2526 GND.n2525 19.3944
R13173 GND.n2525 GND.n2524 19.3944
R13174 GND.n2524 GND.n2521 19.3944
R13175 GND.n2521 GND.n2432 19.3944
R13176 GND.n2718 GND.n2432 19.3944
R13177 GND.n2718 GND.n2430 19.3944
R13178 GND.n2722 GND.n2430 19.3944
R13179 GND.n2726 GND.n2722 19.3944
R13180 GND.n2724 GND.n2723 19.3944
R13181 GND.n2819 GND.n2818 19.3944
R13182 GND.n2816 GND.n2400 19.3944
R13183 GND.n2802 GND.n2750 19.3944
R13184 GND.n2800 GND.n2799 19.3944
R13185 GND.n2799 GND.n2752 19.3944
R13186 GND.n2793 GND.n2752 19.3944
R13187 GND.n2793 GND.n2792 19.3944
R13188 GND.n2792 GND.n2791 19.3944
R13189 GND.n2791 GND.n2758 19.3944
R13190 GND.n2784 GND.n2758 19.3944
R13191 GND.n2784 GND.n2783 19.3944
R13192 GND.n2783 GND.n2782 19.3944
R13193 GND.n2782 GND.n2764 19.3944
R13194 GND.n2778 GND.n2764 19.3944
R13195 GND.n2778 GND.n2777 19.3944
R13196 GND.n2777 GND.n2776 19.3944
R13197 GND.n2776 GND.n2774 19.3944
R13198 GND.n2774 GND.n2314 19.3944
R13199 GND.n2314 GND.n2312 19.3944
R13200 GND.n2915 GND.n2312 19.3944
R13201 GND.n2915 GND.n2310 19.3944
R13202 GND.n2928 GND.n2310 19.3944
R13203 GND.n2928 GND.n2927 19.3944
R13204 GND.n2927 GND.n2926 19.3944
R13205 GND.n2926 GND.n2923 19.3944
R13206 GND.n2923 GND.n1394 19.3944
R13207 GND.n4473 GND.n1394 19.3944
R13208 GND.n4473 GND.n4472 19.3944
R13209 GND.n4472 GND.n4471 19.3944
R13210 GND.n4471 GND.n1398 19.3944
R13211 GND.n1400 GND.n1398 19.3944
R13212 GND.n1421 GND.n1400 19.3944
R13213 GND.n1423 GND.n1421 19.3944
R13214 GND.n1423 GND.n1417 19.3944
R13215 GND.n4455 GND.n1417 19.3944
R13216 GND.n4455 GND.n4454 19.3944
R13217 GND.n4454 GND.n4453 19.3944
R13218 GND.n4453 GND.n1429 19.3944
R13219 GND.n1450 GND.n1429 19.3944
R13220 GND.n4441 GND.n1450 19.3944
R13221 GND.n4441 GND.n4440 19.3944
R13222 GND.n4440 GND.n4439 19.3944
R13223 GND.n4439 GND.n1456 19.3944
R13224 GND.n1477 GND.n1456 19.3944
R13225 GND.n4427 GND.n1477 19.3944
R13226 GND.n4427 GND.n4426 19.3944
R13227 GND.n4426 GND.n4425 19.3944
R13228 GND.n4425 GND.n1483 19.3944
R13229 GND.n4413 GND.n1483 19.3944
R13230 GND.n4413 GND.n4412 19.3944
R13231 GND.n4412 GND.n4411 19.3944
R13232 GND.n4411 GND.n1500 19.3944
R13233 GND.n4399 GND.n1500 19.3944
R13234 GND.n4399 GND.n4398 19.3944
R13235 GND.n4398 GND.n4397 19.3944
R13236 GND.n4397 GND.n1518 19.3944
R13237 GND.n4385 GND.n1518 19.3944
R13238 GND.n4385 GND.n4384 19.3944
R13239 GND.n4384 GND.n4383 19.3944
R13240 GND.n4383 GND.n1538 19.3944
R13241 GND.n1567 GND.n1538 19.3944
R13242 GND.n1567 GND.n1564 19.3944
R13243 GND.n4364 GND.n1564 19.3944
R13244 GND.n4364 GND.n4363 19.3944
R13245 GND.n4363 GND.n4362 19.3944
R13246 GND.n4362 GND.n1573 19.3944
R13247 GND.n1610 GND.n1573 19.3944
R13248 GND.n1610 GND.n1607 19.3944
R13249 GND.n4343 GND.n1607 19.3944
R13250 GND.n4343 GND.n4342 19.3944
R13251 GND.n4342 GND.n4341 19.3944
R13252 GND.n4341 GND.n1616 19.3944
R13253 GND.n3410 GND.n1616 19.3944
R13254 GND.n3415 GND.n3410 19.3944
R13255 GND.n3415 GND.n1656 19.3944
R13256 GND.n4316 GND.n1656 19.3944
R13257 GND.n4316 GND.n4315 19.3944
R13258 GND.n4315 GND.n4314 19.3944
R13259 GND.n4314 GND.n1660 19.3944
R13260 GND.n3762 GND.n1660 19.3944
R13261 GND.n3765 GND.n3762 19.3944
R13262 GND.n3765 GND.n3759 19.3944
R13263 GND.n3770 GND.n3759 19.3944
R13264 GND.n3770 GND.n1700 19.3944
R13265 GND.n4288 GND.n1700 19.3944
R13266 GND.n4288 GND.n4287 19.3944
R13267 GND.n4287 GND.n4286 19.3944
R13268 GND.n4286 GND.n1704 19.3944
R13269 GND.n1725 GND.n1704 19.3944
R13270 GND.n4274 GND.n1725 19.3944
R13271 GND.n4274 GND.n4273 19.3944
R13272 GND.n4273 GND.n4272 19.3944
R13273 GND.n4272 GND.n1731 19.3944
R13274 GND.n1751 GND.n1731 19.3944
R13275 GND.n4260 GND.n1751 19.3944
R13276 GND.n4260 GND.n4259 19.3944
R13277 GND.n4259 GND.n4258 19.3944
R13278 GND.n4258 GND.n1757 19.3944
R13279 GND.n2125 GND.n1757 19.3944
R13280 GND.n2129 GND.n2125 19.3944
R13281 GND.n2129 GND.n2122 19.3944
R13282 GND.n2133 GND.n2122 19.3944
R13283 GND.n2133 GND.n2120 19.3944
R13284 GND.n3846 GND.n2120 19.3944
R13285 GND.n3846 GND.n2118 19.3944
R13286 GND.n3886 GND.n2118 19.3944
R13287 GND.n3886 GND.n3885 19.3944
R13288 GND.n3885 GND.n3884 19.3944
R13289 GND.n3884 GND.n3852 19.3944
R13290 GND.n3880 GND.n3852 19.3944
R13291 GND.n3880 GND.n3879 19.3944
R13292 GND.n3879 GND.n3878 19.3944
R13293 GND.n3878 GND.n3858 19.3944
R13294 GND.n3872 GND.n3858 19.3944
R13295 GND.n3872 GND.n3871 19.3944
R13296 GND.n3871 GND.n3870 19.3944
R13297 GND.n3870 GND.n3867 19.3944
R13298 GND.n3867 GND.n3866 19.3944
R13299 GND.n3866 GND.n2048 19.3944
R13300 GND.n3967 GND.n2048 19.3944
R13301 GND.n3967 GND.n2046 19.3944
R13302 GND.n3975 GND.n2046 19.3944
R13303 GND.n3975 GND.n3974 19.3944
R13304 GND.n3974 GND.n3973 19.3944
R13305 GND.n3973 GND.n2016 19.3944
R13306 GND.n4007 GND.n4006 19.3944
R13307 GND.n4054 GND.n4053 19.3944
R13308 GND.n4051 GND.n4009 19.3944
R13309 GND.n4037 GND.n4035 19.3944
R13310 GND.n4074 GND.n1985 19.3944
R13311 GND.n4074 GND.n1983 19.3944
R13312 GND.n4080 GND.n1983 19.3944
R13313 GND.n4080 GND.n4079 19.3944
R13314 GND.n4079 GND.n1961 19.3944
R13315 GND.n4100 GND.n1961 19.3944
R13316 GND.n4100 GND.n1959 19.3944
R13317 GND.n4113 GND.n1959 19.3944
R13318 GND.n4113 GND.n4112 19.3944
R13319 GND.n4112 GND.n4111 19.3944
R13320 GND.n4111 GND.n4108 19.3944
R13321 GND.n4108 GND.n597 19.3944
R13322 GND.n5484 GND.n597 19.3944
R13323 GND.n5484 GND.n5483 19.3944
R13324 GND.n5483 GND.n5482 19.3944
R13325 GND.n4749 GND.n4748 19.3944
R13326 GND.n4748 GND.n4747 19.3944
R13327 GND.n4747 GND.n4746 19.3944
R13328 GND.n4746 GND.n4744 19.3944
R13329 GND.n4744 GND.n4741 19.3944
R13330 GND.n4741 GND.n4740 19.3944
R13331 GND.n4740 GND.n4737 19.3944
R13332 GND.n4737 GND.n4736 19.3944
R13333 GND.n4736 GND.n4733 19.3944
R13334 GND.n4733 GND.n4732 19.3944
R13335 GND.n4732 GND.n4729 19.3944
R13336 GND.n4729 GND.n4728 19.3944
R13337 GND.n4728 GND.n4725 19.3944
R13338 GND.n4725 GND.n4724 19.3944
R13339 GND.n4724 GND.n4721 19.3944
R13340 GND.n4719 GND.n4716 19.3944
R13341 GND.n4716 GND.n4715 19.3944
R13342 GND.n4715 GND.n4712 19.3944
R13343 GND.n4712 GND.n4711 19.3944
R13344 GND.n4711 GND.n4708 19.3944
R13345 GND.n4708 GND.n4707 19.3944
R13346 GND.n4707 GND.n4704 19.3944
R13347 GND.n4704 GND.n4703 19.3944
R13348 GND.n4703 GND.n4700 19.3944
R13349 GND.n4700 GND.n4699 19.3944
R13350 GND.n4699 GND.n4696 19.3944
R13351 GND.n4696 GND.n4695 19.3944
R13352 GND.n4695 GND.n4692 19.3944
R13353 GND.n4692 GND.n4691 19.3944
R13354 GND.n4691 GND.n4688 19.3944
R13355 GND.n4688 GND.n4687 19.3944
R13356 GND.n2550 GND.n2549 19.3944
R13357 GND.n2621 GND.n2550 19.3944
R13358 GND.n2621 GND.n2546 19.3944
R13359 GND.n2627 GND.n2546 19.3944
R13360 GND.n2627 GND.n2626 19.3944
R13361 GND.n2626 GND.n2490 19.3944
R13362 GND.n2646 GND.n2490 19.3944
R13363 GND.n2646 GND.n2488 19.3944
R13364 GND.n2652 GND.n2488 19.3944
R13365 GND.n2652 GND.n2651 19.3944
R13366 GND.n2651 GND.n2467 19.3944
R13367 GND.n2671 GND.n2467 19.3944
R13368 GND.n2671 GND.n2465 19.3944
R13369 GND.n2677 GND.n2465 19.3944
R13370 GND.n2677 GND.n2676 19.3944
R13371 GND.n2676 GND.n2444 19.3944
R13372 GND.n2708 GND.n2444 19.3944
R13373 GND.n2708 GND.n2442 19.3944
R13374 GND.n2713 GND.n2442 19.3944
R13375 GND.n2713 GND.n2712 19.3944
R13376 GND.n2712 GND.n2386 19.3944
R13377 GND.n2829 GND.n2828 19.3944
R13378 GND.n2410 GND.n2409 19.3944
R13379 GND.n2811 GND.n2810 19.3944
R13380 GND.n2415 GND.n2414 19.3944
R13381 GND.n2834 GND.n2379 19.3944
R13382 GND.n2834 GND.n2833 19.3944
R13383 GND.n2833 GND.n2360 19.3944
R13384 GND.n2853 GND.n2360 19.3944
R13385 GND.n2853 GND.n2358 19.3944
R13386 GND.n2859 GND.n2358 19.3944
R13387 GND.n2859 GND.n2858 19.3944
R13388 GND.n2858 GND.n2341 19.3944
R13389 GND.n2878 GND.n2341 19.3944
R13390 GND.n2878 GND.n2339 19.3944
R13391 GND.n2884 GND.n2339 19.3944
R13392 GND.n2884 GND.n2883 19.3944
R13393 GND.n2883 GND.n2320 19.3944
R13394 GND.n2904 GND.n2320 19.3944
R13395 GND.n2904 GND.n2318 19.3944
R13396 GND.n2908 GND.n2318 19.3944
R13397 GND.n2908 GND.n2294 19.3944
R13398 GND.n2944 GND.n2294 19.3944
R13399 GND.n2944 GND.n2292 19.3944
R13400 GND.n2948 GND.n2292 19.3944
R13401 GND.n2948 GND.n1267 19.3944
R13402 GND.n4598 GND.n1267 19.3944
R13403 GND.n4884 GND.n957 19.3944
R13404 GND.n4878 GND.n957 19.3944
R13405 GND.n4878 GND.n4877 19.3944
R13406 GND.n4877 GND.n4876 19.3944
R13407 GND.n4876 GND.n964 19.3944
R13408 GND.n4870 GND.n964 19.3944
R13409 GND.n4870 GND.n4869 19.3944
R13410 GND.n4869 GND.n4868 19.3944
R13411 GND.n4868 GND.n972 19.3944
R13412 GND.n4862 GND.n972 19.3944
R13413 GND.n4862 GND.n4861 19.3944
R13414 GND.n4861 GND.n4860 19.3944
R13415 GND.n4860 GND.n980 19.3944
R13416 GND.n4854 GND.n980 19.3944
R13417 GND.n4854 GND.n4853 19.3944
R13418 GND.n4853 GND.n4852 19.3944
R13419 GND.n4852 GND.n988 19.3944
R13420 GND.n4846 GND.n988 19.3944
R13421 GND.n4846 GND.n4845 19.3944
R13422 GND.n4845 GND.n4844 19.3944
R13423 GND.n4844 GND.n996 19.3944
R13424 GND.n4838 GND.n996 19.3944
R13425 GND.n4838 GND.n4837 19.3944
R13426 GND.n4837 GND.n4836 19.3944
R13427 GND.n4836 GND.n1004 19.3944
R13428 GND.n4830 GND.n1004 19.3944
R13429 GND.n4830 GND.n4829 19.3944
R13430 GND.n4829 GND.n4828 19.3944
R13431 GND.n4828 GND.n1012 19.3944
R13432 GND.n4822 GND.n1012 19.3944
R13433 GND.n4822 GND.n4821 19.3944
R13434 GND.n4821 GND.n4820 19.3944
R13435 GND.n4820 GND.n1020 19.3944
R13436 GND.n4814 GND.n1020 19.3944
R13437 GND.n4814 GND.n4813 19.3944
R13438 GND.n4813 GND.n4812 19.3944
R13439 GND.n4812 GND.n1028 19.3944
R13440 GND.n4806 GND.n1028 19.3944
R13441 GND.n4806 GND.n4805 19.3944
R13442 GND.n4805 GND.n4804 19.3944
R13443 GND.n4804 GND.n1036 19.3944
R13444 GND.n4798 GND.n1036 19.3944
R13445 GND.n4798 GND.n4797 19.3944
R13446 GND.n4797 GND.n4796 19.3944
R13447 GND.n4796 GND.n1044 19.3944
R13448 GND.n4790 GND.n1044 19.3944
R13449 GND.n4790 GND.n4789 19.3944
R13450 GND.n4789 GND.n4788 19.3944
R13451 GND.n4788 GND.n1052 19.3944
R13452 GND.n4782 GND.n1052 19.3944
R13453 GND.n4782 GND.n4781 19.3944
R13454 GND.n4781 GND.n4780 19.3944
R13455 GND.n4780 GND.n1060 19.3944
R13456 GND.n4774 GND.n1060 19.3944
R13457 GND.n4774 GND.n4773 19.3944
R13458 GND.n4773 GND.n4772 19.3944
R13459 GND.n4772 GND.n1068 19.3944
R13460 GND.n4766 GND.n1068 19.3944
R13461 GND.n4766 GND.n4765 19.3944
R13462 GND.n4765 GND.n4764 19.3944
R13463 GND.n4764 GND.n1076 19.3944
R13464 GND.n4758 GND.n1076 19.3944
R13465 GND.n4758 GND.n4757 19.3944
R13466 GND.n4757 GND.n4756 19.3944
R13467 GND.n4756 GND.n1084 19.3944
R13468 GND.n2540 GND.n1084 19.3944
R13469 GND.n4212 GND.n4211 19.3944
R13470 GND.n4211 GND.n4204 19.3944
R13471 GND.n4204 GND.n1781 19.3944
R13472 GND.n4249 GND.n1781 19.3944
R13473 GND.n4249 GND.n4248 19.3944
R13474 GND.n4248 GND.n1784 19.3944
R13475 GND.n4241 GND.n1784 19.3944
R13476 GND.n4241 GND.n4240 19.3944
R13477 GND.n4240 GND.n1792 19.3944
R13478 GND.n4233 GND.n1792 19.3944
R13479 GND.n4233 GND.n4232 19.3944
R13480 GND.n4232 GND.n1802 19.3944
R13481 GND.n4225 GND.n1802 19.3944
R13482 GND.n4225 GND.n4224 19.3944
R13483 GND.n3841 GND.n2138 19.3944
R13484 GND.n3841 GND.n2139 19.3944
R13485 GND.n2139 GND.n2100 19.3944
R13486 GND.n3905 GND.n2100 19.3944
R13487 GND.n3905 GND.n2097 19.3944
R13488 GND.n3910 GND.n2097 19.3944
R13489 GND.n3910 GND.n2098 19.3944
R13490 GND.n2098 GND.n2078 19.3944
R13491 GND.n3929 GND.n2078 19.3944
R13492 GND.n3929 GND.n2075 19.3944
R13493 GND.n3934 GND.n2075 19.3944
R13494 GND.n3934 GND.n2076 19.3944
R13495 GND.n2076 GND.n2056 19.3944
R13496 GND.n3954 GND.n2056 19.3944
R13497 GND.n3954 GND.n2053 19.3944
R13498 GND.n3961 GND.n2053 19.3944
R13499 GND.n3961 GND.n2054 19.3944
R13500 GND.n3957 GND.n2054 19.3944
R13501 GND.n3957 GND.n2022 19.3944
R13502 GND.n3993 GND.n2022 19.3944
R13503 GND.n3993 GND.n2019 19.3944
R13504 GND.n4000 GND.n2019 19.3944
R13505 GND.n4000 GND.n2020 19.3944
R13506 GND.n3996 GND.n2020 19.3944
R13507 GND.n3996 GND.n428 19.3944
R13508 GND.n5673 GND.n428 19.3944
R13509 GND.n5673 GND.n5672 19.3944
R13510 GND.n5672 GND.n5671 19.3944
R13511 GND.n5671 GND.n432 19.3944
R13512 GND.n5667 GND.n432 19.3944
R13513 GND.n5667 GND.n5666 19.3944
R13514 GND.n5666 GND.n5665 19.3944
R13515 GND.n5665 GND.n437 19.3944
R13516 GND.n5661 GND.n437 19.3944
R13517 GND.n5661 GND.n5660 19.3944
R13518 GND.n5660 GND.n5659 19.3944
R13519 GND.n5659 GND.n442 19.3944
R13520 GND.n5655 GND.n442 19.3944
R13521 GND.n5655 GND.n5654 19.3944
R13522 GND.n5654 GND.n5653 19.3944
R13523 GND.n5653 GND.n447 19.3944
R13524 GND.n5649 GND.n447 19.3944
R13525 GND.n5649 GND.n5648 19.3944
R13526 GND.n5648 GND.n5647 19.3944
R13527 GND.n5647 GND.n452 19.3944
R13528 GND.n5643 GND.n452 19.3944
R13529 GND.n5643 GND.n5642 19.3944
R13530 GND.n5642 GND.n5641 19.3944
R13531 GND.n5641 GND.n457 19.3944
R13532 GND.n5637 GND.n457 19.3944
R13533 GND.n5637 GND.n5636 19.3944
R13534 GND.n5636 GND.n5635 19.3944
R13535 GND.n2787 GND.t9 19.3043
R13536 GND.t46 GND.n2059 19.3043
R13537 GND.n4576 GND.n4575 18.4247
R13538 GND.n3685 GND.n3579 18.4247
R13539 GND.n5545 GND.n465 18.2308
R13540 GND.n4505 GND.n1366 18.2308
R13541 GND.n2589 GND.n2575 18.2308
R13542 GND.n4224 GND.n1812 18.2308
R13543 GND.n4534 GND.n1339 16.4562
R13544 GND.n4255 GND.n4254 16.4562
R13545 GND.n4467 GND.n4466 15.8233
R13546 GND.n4466 GND.n4465 15.8233
R13547 GND.n4465 GND.n4464 15.8233
R13548 GND.n4464 GND.n1403 15.8233
R13549 GND.n3005 GND.n1403 15.8233
R13550 GND.n4458 GND.n1412 15.8233
R13551 GND.n4458 GND.n4457 15.8233
R13552 GND.n4457 GND.n1414 15.8233
R13553 GND.n1431 GND.n1414 15.8233
R13554 GND.n1432 GND.n1431 15.8233
R13555 GND.n4451 GND.n1432 15.8233
R13556 GND.n4451 GND.n4450 15.8233
R13557 GND.n4450 GND.n1434 15.8233
R13558 GND.n2269 GND.n1434 15.8233
R13559 GND.n2269 GND.n1445 15.8233
R13560 GND.n4444 GND.n1445 15.8233
R13561 GND.n4444 GND.n4443 15.8233
R13562 GND.n4443 GND.n1447 15.8233
R13563 GND.n1459 GND.n1458 15.8233
R13564 GND.n4437 GND.n1459 15.8233
R13565 GND.n4437 GND.n4436 15.8233
R13566 GND.n4436 GND.n1461 15.8233
R13567 GND.n3035 GND.n1461 15.8233
R13568 GND.n4430 GND.n1472 15.8233
R13569 GND.n3233 GND.n3232 15.8233
R13570 GND.n3247 GND.n2240 15.8233
R13571 GND.n4395 GND.n4394 15.8233
R13572 GND.n4394 GND.n1523 15.8233
R13573 GND.n4387 GND.n1532 15.8233
R13574 GND.n4381 GND.n4380 15.8233
R13575 GND.n4374 GND.n1550 15.8233
R13576 GND.n4366 GND.n1561 15.8233
R13577 GND.n4360 GND.n1575 15.8233
R13578 GND.n4352 GND.n1586 15.8233
R13579 GND.n4346 GND.n4345 15.8233
R13580 GND.n4339 GND.n1618 15.8233
R13581 GND.n4332 GND.n1626 15.8233
R13582 GND.n4332 GND.n1629 15.8233
R13583 GND.n4318 GND.n1653 15.8233
R13584 GND.n4312 GND.n4311 15.8233
R13585 GND.n4305 GND.n1678 15.8233
R13586 GND.n3780 GND.n1686 15.8233
R13587 GND.n3772 GND.n3757 15.8233
R13588 GND.n3757 GND.n3756 15.8233
R13589 GND.n4291 GND.n4290 15.8233
R13590 GND.n4290 GND.n1697 15.8233
R13591 GND.n1706 GND.n1697 15.8233
R13592 GND.n1707 GND.n1706 15.8233
R13593 GND.n4284 GND.n1707 15.8233
R13594 GND.n4283 GND.n1709 15.8233
R13595 GND.n2171 GND.n1709 15.8233
R13596 GND.n2171 GND.n1720 15.8233
R13597 GND.n4277 GND.n1720 15.8233
R13598 GND.n4277 GND.n4276 15.8233
R13599 GND.n4276 GND.n1722 15.8233
R13600 GND.n1733 GND.n1722 15.8233
R13601 GND.n1734 GND.n1733 15.8233
R13602 GND.n4270 GND.n1734 15.8233
R13603 GND.n4270 GND.n4269 15.8233
R13604 GND.n4269 GND.n1736 15.8233
R13605 GND.n3805 GND.n1736 15.8233
R13606 GND.n3805 GND.n3804 15.8233
R13607 GND.n4263 GND.n4262 15.8233
R13608 GND.n4262 GND.n1748 15.8233
R13609 GND.n1759 GND.n1748 15.8233
R13610 GND.n1760 GND.n1759 15.8233
R13611 GND.n4256 GND.n1760 15.8233
R13612 GND.n80 GND.n78 15.6674
R13613 GND.n117 GND.n115 15.6674
R13614 GND.n149 GND.n147 15.6674
R13615 GND.n186 GND.n184 15.6674
R13616 GND.n11 GND.n9 15.6674
R13617 GND.n48 GND.n46 15.6674
R13618 GND.n265 GND.n263 15.6674
R13619 GND.n228 GND.n226 15.6674
R13620 GND.n334 GND.n332 15.6674
R13621 GND.n297 GND.n295 15.6674
R13622 GND.n404 GND.n402 15.6674
R13623 GND.n367 GND.n365 15.6674
R13624 GND.n3005 GND.t125 15.5068
R13625 GND.n4263 GND.t132 15.5068
R13626 GND.n4534 GND.n1325 15.1904
R13627 GND.n3231 GND.n2241 15.1904
R13628 GND.n4367 GND.n1559 15.1904
R13629 GND.n4359 GND.n1577 15.1904
R13630 GND.n3451 GND.n3450 15.1904
R13631 GND.n4298 GND.n4297 15.1904
R13632 GND.n4254 GND.n1761 15.1904
R13633 GND.n3498 GND.n3497 15.0827
R13634 GND.n2252 GND.n2247 15.0481
R13635 GND.n3508 GND.n3507 15.0481
R13636 GND.n4401 GND.n1512 14.5575
R13637 GND.n3304 GND.n3303 14.5575
R13638 GND.n3376 GND.n2200 14.5575
R13639 GND.n4325 GND.n1645 14.5575
R13640 GND.n3223 GND.n3035 14.241
R13641 GND.n4430 GND.t97 13.9246
R13642 GND.n3272 GND.n2230 13.9246
R13643 GND.n5579 GND.n549 13.5763
R13644 GND.n4550 GND.n1314 13.5763
R13645 GND.n3652 GND.n3649 13.5763
R13646 GND.n4687 GND.n1153 13.5763
R13647 GND.n2232 GND.t119 13.2916
R13648 GND.n4409 GND.n4408 13.2916
R13649 GND.n3138 GND.t148 13.2916
R13650 GND.n2209 GND.n1541 13.2916
R13651 GND.n3385 GND.n1603 13.2916
R13652 GND.n2187 GND.n2186 13.2916
R13653 GND.n2263 GND.n2244 13.1884
R13654 GND.n2258 GND.n2257 13.1884
R13655 GND.n2257 GND.n2256 13.1884
R13656 GND.n3501 GND.n3496 13.1884
R13657 GND.n3502 GND.n3501 13.1884
R13658 GND.n2259 GND.n2246 13.146
R13659 GND.n2255 GND.n2246 13.146
R13660 GND.n3500 GND.n3499 13.146
R13661 GND.n3500 GND.n3495 13.146
R13662 GND.n81 GND.n77 12.8005
R13663 GND.n118 GND.n114 12.8005
R13664 GND.n150 GND.n146 12.8005
R13665 GND.n187 GND.n183 12.8005
R13666 GND.n12 GND.n8 12.8005
R13667 GND.n49 GND.n45 12.8005
R13668 GND.n266 GND.n262 12.8005
R13669 GND.n229 GND.n225 12.8005
R13670 GND.n335 GND.n331 12.8005
R13671 GND.n298 GND.n294 12.8005
R13672 GND.n405 GND.n401 12.8005
R13673 GND.n368 GND.n364 12.8005
R13674 GND.n3139 GND.n1510 12.6587
R13675 GND.t21 GND.n3255 12.6587
R13676 GND.n3320 GND.n3319 12.6587
R13677 GND.n3394 GND.n2198 12.6587
R13678 GND.n3417 GND.t63 12.6587
R13679 GND.n4319 GND.n1651 12.6587
R13680 GND.n5575 GND.n549 12.4126
R13681 GND.n4546 GND.n1314 12.4126
R13682 GND.n3649 GND.n3645 12.4126
R13683 GND.n4683 GND.n1153 12.4126
R13684 GND.n3227 GND.n3226 12.1761
R13685 GND.n3515 GND.n3513 12.1761
R13686 GND.n4501 GND.n4475 12.0258
R13687 GND.n4415 GND.n1494 12.0258
R13688 GND.n4373 GND.n1553 12.0258
R13689 GND.n4353 GND.n1583 12.0258
R13690 GND.t116 GND.n1662 12.0258
R13691 GND.n2180 GND.n1664 12.0258
R13692 GND.n4214 GND.n1822 12.0258
R13693 GND.n85 GND.n84 12.0247
R13694 GND.n122 GND.n121 12.0247
R13695 GND.n154 GND.n153 12.0247
R13696 GND.n191 GND.n190 12.0247
R13697 GND.n16 GND.n15 12.0247
R13698 GND.n53 GND.n52 12.0247
R13699 GND.n270 GND.n269 12.0247
R13700 GND.n233 GND.n232 12.0247
R13701 GND.n339 GND.n338 12.0247
R13702 GND.n302 GND.n301 12.0247
R13703 GND.n409 GND.n408 12.0247
R13704 GND.n372 GND.n371 12.0247
R13705 GND.n2629 GND.n2542 11.7094
R13706 GND.n573 GND.n562 11.7094
R13707 GND.n3294 GND.n3291 11.3929
R13708 GND.n4388 GND.n1530 11.3929
R13709 GND.n4338 GND.n1620 11.3929
R13710 GND.n3418 GND.n3408 11.3929
R13711 GND.n88 GND.n75 11.249
R13712 GND.n125 GND.n112 11.249
R13713 GND.n157 GND.n144 11.249
R13714 GND.n194 GND.n181 11.249
R13715 GND.n19 GND.n6 11.249
R13716 GND.n56 GND.n43 11.249
R13717 GND.n273 GND.n260 11.249
R13718 GND.n236 GND.n223 11.249
R13719 GND.n342 GND.n329 11.249
R13720 GND.n305 GND.n292 11.249
R13721 GND.n412 GND.n399 11.249
R13722 GND.n375 GND.n362 11.249
R13723 GND.n2870 GND.t9 11.0764
R13724 GND.n3952 GND.t46 11.0764
R13725 GND.n4423 GND.n1485 10.76
R13726 GND.n4423 GND.n4422 10.76
R13727 GND.n3361 GND.n3360 10.76
R13728 GND.n3362 GND.n3361 10.76
R13729 GND.n3779 GND.n2177 10.76
R13730 GND.n3752 GND.n3751 10.6151
R13731 GND.n3751 GND.n3748 10.6151
R13732 GND.n3746 GND.n3743 10.6151
R13733 GND.n3743 GND.n3742 10.6151
R13734 GND.n3742 GND.n3739 10.6151
R13735 GND.n3739 GND.n3738 10.6151
R13736 GND.n3738 GND.n3735 10.6151
R13737 GND.n3735 GND.n3734 10.6151
R13738 GND.n3734 GND.n3731 10.6151
R13739 GND.n3731 GND.n3730 10.6151
R13740 GND.n3730 GND.n3727 10.6151
R13741 GND.n3727 GND.n3726 10.6151
R13742 GND.n3726 GND.n3723 10.6151
R13743 GND.n3723 GND.n3722 10.6151
R13744 GND.n3722 GND.n3719 10.6151
R13745 GND.n3719 GND.n3718 10.6151
R13746 GND.n3718 GND.n3715 10.6151
R13747 GND.n3715 GND.n3714 10.6151
R13748 GND.n3714 GND.n3711 10.6151
R13749 GND.n3711 GND.n3710 10.6151
R13750 GND.n3710 GND.n3707 10.6151
R13751 GND.n3707 GND.n3706 10.6151
R13752 GND.n3706 GND.n3703 10.6151
R13753 GND.n3703 GND.n3702 10.6151
R13754 GND.n3702 GND.n3699 10.6151
R13755 GND.n3699 GND.n3698 10.6151
R13756 GND.n3698 GND.n3695 10.6151
R13757 GND.n3695 GND.n3694 10.6151
R13758 GND.n3694 GND.n3691 10.6151
R13759 GND.n3691 GND.n3455 10.6151
R13760 GND.n3156 GND.n3155 10.6151
R13761 GND.n3155 GND.n3154 10.6151
R13762 GND.n3154 GND.n3152 10.6151
R13763 GND.n3152 GND.n3151 10.6151
R13764 GND.n3151 GND.n3148 10.6151
R13765 GND.n3148 GND.n3147 10.6151
R13766 GND.n3147 GND.n3135 10.6151
R13767 GND.n3143 GND.n3135 10.6151
R13768 GND.n3143 GND.n3142 10.6151
R13769 GND.n3142 GND.n3141 10.6151
R13770 GND.n3141 GND.n3137 10.6151
R13771 GND.n3137 GND.n3136 10.6151
R13772 GND.n3136 GND.n2219 10.6151
R13773 GND.n3297 GND.n2219 10.6151
R13774 GND.n3298 GND.n3297 10.6151
R13775 GND.n3301 GND.n3298 10.6151
R13776 GND.n3302 GND.n3301 10.6151
R13777 GND.n3306 GND.n3302 10.6151
R13778 GND.n3307 GND.n3306 10.6151
R13779 GND.n3309 GND.n3307 10.6151
R13780 GND.n3309 GND.n3308 10.6151
R13781 GND.n3308 GND.n2207 10.6151
R13782 GND.n3352 GND.n2207 10.6151
R13783 GND.n3353 GND.n3352 10.6151
R13784 GND.n3356 GND.n3353 10.6151
R13785 GND.n3357 GND.n3356 10.6151
R13786 GND.n3358 GND.n3357 10.6151
R13787 GND.n3364 GND.n3358 10.6151
R13788 GND.n3365 GND.n3364 10.6151
R13789 GND.n3368 GND.n3365 10.6151
R13790 GND.n3369 GND.n3368 10.6151
R13791 GND.n3370 GND.n3369 10.6151
R13792 GND.n3383 GND.n3370 10.6151
R13793 GND.n3383 GND.n3382 10.6151
R13794 GND.n3382 GND.n3381 10.6151
R13795 GND.n3381 GND.n3379 10.6151
R13796 GND.n3379 GND.n3378 10.6151
R13797 GND.n3378 GND.n3375 10.6151
R13798 GND.n3375 GND.n3374 10.6151
R13799 GND.n3374 GND.n3371 10.6151
R13800 GND.n3371 GND.n2190 10.6151
R13801 GND.n3420 GND.n2190 10.6151
R13802 GND.n3421 GND.n3420 10.6151
R13803 GND.n3424 GND.n3421 10.6151
R13804 GND.n3425 GND.n3424 10.6151
R13805 GND.n3426 GND.n3425 10.6151
R13806 GND.n3430 GND.n3426 10.6151
R13807 GND.n3430 GND.n3429 10.6151
R13808 GND.n3429 GND.n3428 10.6151
R13809 GND.n3428 GND.n2178 10.6151
R13810 GND.n3453 GND.n2178 10.6151
R13811 GND.n3454 GND.n3453 10.6151
R13812 GND.n3777 GND.n3454 10.6151
R13813 GND.n3777 GND.n3776 10.6151
R13814 GND.n3776 GND.n3775 10.6151
R13815 GND.n3075 GND.n3074 10.6151
R13816 GND.n3078 GND.n3075 10.6151
R13817 GND.n3083 GND.n3080 10.6151
R13818 GND.n3084 GND.n3083 10.6151
R13819 GND.n3087 GND.n3084 10.6151
R13820 GND.n3088 GND.n3087 10.6151
R13821 GND.n3091 GND.n3088 10.6151
R13822 GND.n3092 GND.n3091 10.6151
R13823 GND.n3095 GND.n3092 10.6151
R13824 GND.n3096 GND.n3095 10.6151
R13825 GND.n3099 GND.n3096 10.6151
R13826 GND.n3100 GND.n3099 10.6151
R13827 GND.n3103 GND.n3100 10.6151
R13828 GND.n3104 GND.n3103 10.6151
R13829 GND.n3107 GND.n3104 10.6151
R13830 GND.n3108 GND.n3107 10.6151
R13831 GND.n3111 GND.n3108 10.6151
R13832 GND.n3112 GND.n3111 10.6151
R13833 GND.n3115 GND.n3112 10.6151
R13834 GND.n3116 GND.n3115 10.6151
R13835 GND.n3119 GND.n3116 10.6151
R13836 GND.n3120 GND.n3119 10.6151
R13837 GND.n3123 GND.n3120 10.6151
R13838 GND.n3124 GND.n3123 10.6151
R13839 GND.n3127 GND.n3124 10.6151
R13840 GND.n3128 GND.n3127 10.6151
R13841 GND.n3131 GND.n3128 10.6151
R13842 GND.n3133 GND.n3131 10.6151
R13843 GND.n3134 GND.n3133 10.6151
R13844 GND.n3157 GND.n3134 10.6151
R13845 GND.n3226 GND.n2264 10.6151
R13846 GND.n3221 GND.n2264 10.6151
R13847 GND.n3221 GND.n3220 10.6151
R13848 GND.n3220 GND.n3219 10.6151
R13849 GND.n3219 GND.n3216 10.6151
R13850 GND.n3216 GND.n3215 10.6151
R13851 GND.n3215 GND.n3212 10.6151
R13852 GND.n3212 GND.n3211 10.6151
R13853 GND.n3211 GND.n3208 10.6151
R13854 GND.n3208 GND.n3207 10.6151
R13855 GND.n3207 GND.n3204 10.6151
R13856 GND.n3204 GND.n3203 10.6151
R13857 GND.n3203 GND.n3200 10.6151
R13858 GND.n3200 GND.n3199 10.6151
R13859 GND.n3199 GND.n3196 10.6151
R13860 GND.n3196 GND.n3195 10.6151
R13861 GND.n3195 GND.n3192 10.6151
R13862 GND.n3192 GND.n3191 10.6151
R13863 GND.n3191 GND.n3188 10.6151
R13864 GND.n3188 GND.n3187 10.6151
R13865 GND.n3187 GND.n3184 10.6151
R13866 GND.n3184 GND.n3183 10.6151
R13867 GND.n3183 GND.n3180 10.6151
R13868 GND.n3180 GND.n3179 10.6151
R13869 GND.n3179 GND.n3176 10.6151
R13870 GND.n3176 GND.n3175 10.6151
R13871 GND.n3175 GND.n3172 10.6151
R13872 GND.n3172 GND.n3171 10.6151
R13873 GND.n3168 GND.n3167 10.6151
R13874 GND.n3167 GND.n3164 10.6151
R13875 GND.n3516 GND.n3515 10.6151
R13876 GND.n3519 GND.n3516 10.6151
R13877 GND.n3520 GND.n3519 10.6151
R13878 GND.n3523 GND.n3520 10.6151
R13879 GND.n3524 GND.n3523 10.6151
R13880 GND.n3527 GND.n3524 10.6151
R13881 GND.n3528 GND.n3527 10.6151
R13882 GND.n3531 GND.n3528 10.6151
R13883 GND.n3532 GND.n3531 10.6151
R13884 GND.n3535 GND.n3532 10.6151
R13885 GND.n3536 GND.n3535 10.6151
R13886 GND.n3539 GND.n3536 10.6151
R13887 GND.n3540 GND.n3539 10.6151
R13888 GND.n3543 GND.n3540 10.6151
R13889 GND.n3544 GND.n3543 10.6151
R13890 GND.n3547 GND.n3544 10.6151
R13891 GND.n3548 GND.n3547 10.6151
R13892 GND.n3551 GND.n3548 10.6151
R13893 GND.n3552 GND.n3551 10.6151
R13894 GND.n3555 GND.n3552 10.6151
R13895 GND.n3556 GND.n3555 10.6151
R13896 GND.n3559 GND.n3556 10.6151
R13897 GND.n3560 GND.n3559 10.6151
R13898 GND.n3563 GND.n3560 10.6151
R13899 GND.n3564 GND.n3563 10.6151
R13900 GND.n3567 GND.n3564 10.6151
R13901 GND.n3568 GND.n3567 10.6151
R13902 GND.n3571 GND.n3568 10.6151
R13903 GND.n3576 GND.n3573 10.6151
R13904 GND.n3577 GND.n3576 10.6151
R13905 GND.n3229 GND.n3228 10.6151
R13906 GND.n3229 GND.n1489 10.6151
R13907 GND.n4420 GND.n1489 10.6151
R13908 GND.n4420 GND.n4419 10.6151
R13909 GND.n4419 GND.n4418 10.6151
R13910 GND.n4418 GND.n1490 10.6151
R13911 GND.n2228 GND.n1490 10.6151
R13912 GND.n2228 GND.n1507 10.6151
R13913 GND.n4406 GND.n1507 10.6151
R13914 GND.n4406 GND.n4405 10.6151
R13915 GND.n4405 GND.n4404 10.6151
R13916 GND.n4404 GND.n1508 10.6151
R13917 GND.n3292 GND.n1508 10.6151
R13918 GND.n3292 GND.n1527 10.6151
R13919 GND.n4392 GND.n1527 10.6151
R13920 GND.n4392 GND.n4391 10.6151
R13921 GND.n4391 GND.n4390 10.6151
R13922 GND.n4390 GND.n1528 10.6151
R13923 GND.n3313 GND.n1528 10.6151
R13924 GND.n3317 GND.n3313 10.6151
R13925 GND.n3317 GND.n3316 10.6151
R13926 GND.n3316 GND.n3315 10.6151
R13927 GND.n3315 GND.n1556 10.6151
R13928 GND.n4371 GND.n1556 10.6151
R13929 GND.n4371 GND.n4370 10.6151
R13930 GND.n4370 GND.n4369 10.6151
R13931 GND.n4369 GND.n1557 10.6151
R13932 GND.n1580 GND.n1557 10.6151
R13933 GND.n4357 GND.n1580 10.6151
R13934 GND.n4357 GND.n4356 10.6151
R13935 GND.n4356 GND.n4355 10.6151
R13936 GND.n4355 GND.n1581 10.6151
R13937 GND.n2202 GND.n1581 10.6151
R13938 GND.n3389 GND.n2202 10.6151
R13939 GND.n3390 GND.n3389 10.6151
R13940 GND.n3391 GND.n3390 10.6151
R13941 GND.n3391 GND.n1623 10.6151
R13942 GND.n4336 GND.n1623 10.6151
R13943 GND.n4336 GND.n4335 10.6151
R13944 GND.n4335 GND.n4334 10.6151
R13945 GND.n4334 GND.n1624 10.6151
R13946 GND.n1648 GND.n1624 10.6151
R13947 GND.n4323 GND.n1648 10.6151
R13948 GND.n4323 GND.n4322 10.6151
R13949 GND.n4322 GND.n4321 10.6151
R13950 GND.n4321 GND.n1649 10.6151
R13951 GND.n3438 GND.n1649 10.6151
R13952 GND.n3438 GND.n3437 10.6151
R13953 GND.n3437 GND.n3436 10.6151
R13954 GND.n3436 GND.n3433 10.6151
R13955 GND.n3433 GND.n1683 10.6151
R13956 GND.n4302 GND.n1683 10.6151
R13957 GND.n4302 GND.n4301 10.6151
R13958 GND.n4301 GND.n4300 10.6151
R13959 GND.n4300 GND.n1684 10.6151
R13960 GND.n89 GND.n73 10.4732
R13961 GND.n126 GND.n110 10.4732
R13962 GND.n158 GND.n142 10.4732
R13963 GND.n195 GND.n179 10.4732
R13964 GND.n20 GND.n4 10.4732
R13965 GND.n57 GND.n41 10.4732
R13966 GND.n274 GND.n258 10.4732
R13967 GND.n237 GND.n221 10.4732
R13968 GND.n343 GND.n327 10.4732
R13969 GND.n306 GND.n290 10.4732
R13970 GND.n413 GND.n397 10.4732
R13971 GND.n376 GND.n360 10.4732
R13972 GND.n2822 GND.t61 10.4435
R13973 GND.t14 GND.n1447 10.4435
R13974 GND.t22 GND.n4283 10.4435
R13975 GND.n4043 GND.t48 10.4435
R13976 GND.n3291 GND.n1520 10.1271
R13977 GND.n3408 GND.n2192 10.1271
R13978 GND.n2486 GND.t0 9.81063
R13979 GND.t40 GND.n2460 9.81063
R13980 GND.t2 GND.n1965 9.81063
R13981 GND.n4130 GND.t24 9.81063
R13982 GND.n93 GND.n92 9.69747
R13983 GND.n130 GND.n129 9.69747
R13984 GND.n162 GND.n161 9.69747
R13985 GND.n199 GND.n198 9.69747
R13986 GND.n24 GND.n23 9.69747
R13987 GND.n61 GND.n60 9.69747
R13988 GND.n278 GND.n277 9.69747
R13989 GND.n241 GND.n240 9.69747
R13990 GND.n347 GND.n346 9.69747
R13991 GND.n310 GND.n309 9.69747
R13992 GND.n417 GND.n416 9.69747
R13993 GND.n380 GND.n379 9.69747
R13994 GND.n4429 GND.n1474 9.49417
R13995 GND.n3354 GND.n1553 9.49417
R13996 GND.n3366 GND.n1583 9.49417
R13997 GND.n3773 GND.n3772 9.49417
R13998 GND.n4291 GND.t113 9.49417
R13999 GND.n99 GND.n98 9.45567
R14000 GND.n136 GND.n135 9.45567
R14001 GND.n168 GND.n167 9.45567
R14002 GND.n205 GND.n204 9.45567
R14003 GND.n30 GND.n29 9.45567
R14004 GND.n67 GND.n66 9.45567
R14005 GND.n284 GND.n283 9.45567
R14006 GND.n247 GND.n246 9.45567
R14007 GND.n353 GND.n352 9.45567
R14008 GND.n316 GND.n315 9.45567
R14009 GND.n423 GND.n422 9.45567
R14010 GND.n386 GND.n385 9.45567
R14011 GND.n98 GND.n97 9.3005
R14012 GND.n71 GND.n70 9.3005
R14013 GND.n92 GND.n91 9.3005
R14014 GND.n90 GND.n89 9.3005
R14015 GND.n75 GND.n74 9.3005
R14016 GND.n84 GND.n83 9.3005
R14017 GND.n82 GND.n81 9.3005
R14018 GND.n135 GND.n134 9.3005
R14019 GND.n108 GND.n107 9.3005
R14020 GND.n129 GND.n128 9.3005
R14021 GND.n127 GND.n126 9.3005
R14022 GND.n112 GND.n111 9.3005
R14023 GND.n121 GND.n120 9.3005
R14024 GND.n119 GND.n118 9.3005
R14025 GND.n167 GND.n166 9.3005
R14026 GND.n140 GND.n139 9.3005
R14027 GND.n161 GND.n160 9.3005
R14028 GND.n159 GND.n158 9.3005
R14029 GND.n144 GND.n143 9.3005
R14030 GND.n153 GND.n152 9.3005
R14031 GND.n151 GND.n150 9.3005
R14032 GND.n204 GND.n203 9.3005
R14033 GND.n177 GND.n176 9.3005
R14034 GND.n198 GND.n197 9.3005
R14035 GND.n196 GND.n195 9.3005
R14036 GND.n181 GND.n180 9.3005
R14037 GND.n190 GND.n189 9.3005
R14038 GND.n188 GND.n187 9.3005
R14039 GND.n29 GND.n28 9.3005
R14040 GND.n2 GND.n1 9.3005
R14041 GND.n23 GND.n22 9.3005
R14042 GND.n21 GND.n20 9.3005
R14043 GND.n6 GND.n5 9.3005
R14044 GND.n15 GND.n14 9.3005
R14045 GND.n13 GND.n12 9.3005
R14046 GND.n66 GND.n65 9.3005
R14047 GND.n39 GND.n38 9.3005
R14048 GND.n60 GND.n59 9.3005
R14049 GND.n58 GND.n57 9.3005
R14050 GND.n43 GND.n42 9.3005
R14051 GND.n52 GND.n51 9.3005
R14052 GND.n50 GND.n49 9.3005
R14053 GND.n283 GND.n282 9.3005
R14054 GND.n256 GND.n255 9.3005
R14055 GND.n277 GND.n276 9.3005
R14056 GND.n275 GND.n274 9.3005
R14057 GND.n260 GND.n259 9.3005
R14058 GND.n269 GND.n268 9.3005
R14059 GND.n267 GND.n266 9.3005
R14060 GND.n246 GND.n245 9.3005
R14061 GND.n219 GND.n218 9.3005
R14062 GND.n240 GND.n239 9.3005
R14063 GND.n238 GND.n237 9.3005
R14064 GND.n223 GND.n222 9.3005
R14065 GND.n232 GND.n231 9.3005
R14066 GND.n230 GND.n229 9.3005
R14067 GND.n352 GND.n351 9.3005
R14068 GND.n325 GND.n324 9.3005
R14069 GND.n346 GND.n345 9.3005
R14070 GND.n344 GND.n343 9.3005
R14071 GND.n329 GND.n328 9.3005
R14072 GND.n338 GND.n337 9.3005
R14073 GND.n336 GND.n335 9.3005
R14074 GND.n315 GND.n314 9.3005
R14075 GND.n288 GND.n287 9.3005
R14076 GND.n309 GND.n308 9.3005
R14077 GND.n307 GND.n306 9.3005
R14078 GND.n292 GND.n291 9.3005
R14079 GND.n301 GND.n300 9.3005
R14080 GND.n299 GND.n298 9.3005
R14081 GND.n422 GND.n421 9.3005
R14082 GND.n395 GND.n394 9.3005
R14083 GND.n416 GND.n415 9.3005
R14084 GND.n414 GND.n413 9.3005
R14085 GND.n399 GND.n398 9.3005
R14086 GND.n408 GND.n407 9.3005
R14087 GND.n406 GND.n405 9.3005
R14088 GND.n385 GND.n384 9.3005
R14089 GND.n358 GND.n357 9.3005
R14090 GND.n379 GND.n378 9.3005
R14091 GND.n377 GND.n376 9.3005
R14092 GND.n362 GND.n361 9.3005
R14093 GND.n371 GND.n370 9.3005
R14094 GND.n369 GND.n368 9.3005
R14095 GND.n4462 GND.n1407 9.3005
R14096 GND.n4461 GND.n1408 9.3005
R14097 GND.n4460 GND.n1409 9.3005
R14098 GND.n1438 GND.n1410 9.3005
R14099 GND.n1439 GND.n1437 9.3005
R14100 GND.n4448 GND.n1440 9.3005
R14101 GND.n4447 GND.n1441 9.3005
R14102 GND.n4446 GND.n1442 9.3005
R14103 GND.n1465 GND.n1443 9.3005
R14104 GND.n1466 GND.n1464 9.3005
R14105 GND.n4434 GND.n1467 9.3005
R14106 GND.n4433 GND.n1468 9.3005
R14107 GND.n4432 GND.n1469 9.3005
R14108 GND.n3237 GND.n1470 9.3005
R14109 GND.n3238 GND.n3236 9.3005
R14110 GND.n3245 GND.n3239 9.3005
R14111 GND.n3244 GND.n3240 9.3005
R14112 GND.n3243 GND.n3242 9.3005
R14113 GND.n3241 GND.n2227 9.3005
R14114 GND.n2225 GND.n2224 9.3005
R14115 GND.n3277 GND.n3276 9.3005
R14116 GND.n3278 GND.n2223 9.3005
R14117 GND.n3289 GND.n3279 9.3005
R14118 GND.n3288 GND.n3280 9.3005
R14119 GND.n3287 GND.n3281 9.3005
R14120 GND.n3284 GND.n3283 9.3005
R14121 GND.n3282 GND.n1544 9.3005
R14122 GND.n4378 GND.n1545 9.3005
R14123 GND.n4377 GND.n1546 9.3005
R14124 GND.n4376 GND.n1547 9.3005
R14125 GND.n1590 GND.n1548 9.3005
R14126 GND.n1592 GND.n1591 9.3005
R14127 GND.n1596 GND.n1595 9.3005
R14128 GND.n1597 GND.n1589 9.3005
R14129 GND.n4350 GND.n1598 9.3005
R14130 GND.n4349 GND.n1599 9.3005
R14131 GND.n4348 GND.n1600 9.3005
R14132 GND.n1633 GND.n1601 9.3005
R14133 GND.n1636 GND.n1635 9.3005
R14134 GND.n1637 GND.n1632 9.3005
R14135 GND.n4330 GND.n1638 9.3005
R14136 GND.n4329 GND.n1639 9.3005
R14137 GND.n4328 GND.n1640 9.3005
R14138 GND.n1668 GND.n1641 9.3005
R14139 GND.n1671 GND.n1670 9.3005
R14140 GND.n1672 GND.n1667 9.3005
R14141 GND.n4309 GND.n1673 9.3005
R14142 GND.n4308 GND.n1674 9.3005
R14143 GND.n4307 GND.n1675 9.3005
R14144 GND.n1690 GND.n1676 9.3005
R14145 GND.n4295 GND.n1691 9.3005
R14146 GND.n4294 GND.n1692 9.3005
R14147 GND.n4293 GND.n1693 9.3005
R14148 GND.n1713 GND.n1694 9.3005
R14149 GND.n1714 GND.n1712 9.3005
R14150 GND.n4281 GND.n1715 9.3005
R14151 GND.n4280 GND.n1716 9.3005
R14152 GND.n4279 GND.n1717 9.3005
R14153 GND.n1740 GND.n1718 9.3005
R14154 GND.n1741 GND.n1739 9.3005
R14155 GND.n4267 GND.n1742 9.3005
R14156 GND.n4266 GND.n1743 9.3005
R14157 GND.n4265 GND.n1744 9.3005
R14158 GND.n4205 GND.n1745 9.3005
R14159 GND.n4207 GND.n4206 9.3005
R14160 GND.n1406 GND.n1405 9.3005
R14161 GND.n4886 GND.n955 9.3005
R14162 GND.n4888 GND.n4887 9.3005
R14163 GND.n951 GND.n950 9.3005
R14164 GND.n4895 GND.n4894 9.3005
R14165 GND.n4896 GND.n949 9.3005
R14166 GND.n4898 GND.n4897 9.3005
R14167 GND.n945 GND.n944 9.3005
R14168 GND.n4905 GND.n4904 9.3005
R14169 GND.n4906 GND.n943 9.3005
R14170 GND.n4908 GND.n4907 9.3005
R14171 GND.n939 GND.n938 9.3005
R14172 GND.n4915 GND.n4914 9.3005
R14173 GND.n4916 GND.n937 9.3005
R14174 GND.n4918 GND.n4917 9.3005
R14175 GND.n933 GND.n932 9.3005
R14176 GND.n4925 GND.n4924 9.3005
R14177 GND.n4926 GND.n931 9.3005
R14178 GND.n4928 GND.n4927 9.3005
R14179 GND.n927 GND.n926 9.3005
R14180 GND.n4935 GND.n4934 9.3005
R14181 GND.n4936 GND.n925 9.3005
R14182 GND.n4938 GND.n4937 9.3005
R14183 GND.n921 GND.n920 9.3005
R14184 GND.n4945 GND.n4944 9.3005
R14185 GND.n4946 GND.n919 9.3005
R14186 GND.n4948 GND.n4947 9.3005
R14187 GND.n915 GND.n914 9.3005
R14188 GND.n4955 GND.n4954 9.3005
R14189 GND.n4956 GND.n913 9.3005
R14190 GND.n4958 GND.n4957 9.3005
R14191 GND.n909 GND.n908 9.3005
R14192 GND.n4965 GND.n4964 9.3005
R14193 GND.n4966 GND.n907 9.3005
R14194 GND.n4968 GND.n4967 9.3005
R14195 GND.n903 GND.n902 9.3005
R14196 GND.n4975 GND.n4974 9.3005
R14197 GND.n4976 GND.n901 9.3005
R14198 GND.n4978 GND.n4977 9.3005
R14199 GND.n897 GND.n896 9.3005
R14200 GND.n4985 GND.n4984 9.3005
R14201 GND.n4986 GND.n895 9.3005
R14202 GND.n4988 GND.n4987 9.3005
R14203 GND.n891 GND.n890 9.3005
R14204 GND.n4995 GND.n4994 9.3005
R14205 GND.n4996 GND.n889 9.3005
R14206 GND.n4998 GND.n4997 9.3005
R14207 GND.n885 GND.n884 9.3005
R14208 GND.n5005 GND.n5004 9.3005
R14209 GND.n5006 GND.n883 9.3005
R14210 GND.n5008 GND.n5007 9.3005
R14211 GND.n879 GND.n878 9.3005
R14212 GND.n5015 GND.n5014 9.3005
R14213 GND.n5016 GND.n877 9.3005
R14214 GND.n5018 GND.n5017 9.3005
R14215 GND.n873 GND.n872 9.3005
R14216 GND.n5025 GND.n5024 9.3005
R14217 GND.n5026 GND.n871 9.3005
R14218 GND.n5028 GND.n5027 9.3005
R14219 GND.n867 GND.n866 9.3005
R14220 GND.n5035 GND.n5034 9.3005
R14221 GND.n5036 GND.n865 9.3005
R14222 GND.n5038 GND.n5037 9.3005
R14223 GND.n861 GND.n860 9.3005
R14224 GND.n5045 GND.n5044 9.3005
R14225 GND.n5046 GND.n859 9.3005
R14226 GND.n5048 GND.n5047 9.3005
R14227 GND.n855 GND.n854 9.3005
R14228 GND.n5055 GND.n5054 9.3005
R14229 GND.n5056 GND.n853 9.3005
R14230 GND.n5058 GND.n5057 9.3005
R14231 GND.n849 GND.n848 9.3005
R14232 GND.n5065 GND.n5064 9.3005
R14233 GND.n5066 GND.n847 9.3005
R14234 GND.n5068 GND.n5067 9.3005
R14235 GND.n843 GND.n842 9.3005
R14236 GND.n5075 GND.n5074 9.3005
R14237 GND.n5076 GND.n841 9.3005
R14238 GND.n5078 GND.n5077 9.3005
R14239 GND.n837 GND.n836 9.3005
R14240 GND.n5085 GND.n5084 9.3005
R14241 GND.n5086 GND.n835 9.3005
R14242 GND.n5088 GND.n5087 9.3005
R14243 GND.n831 GND.n830 9.3005
R14244 GND.n5095 GND.n5094 9.3005
R14245 GND.n5096 GND.n829 9.3005
R14246 GND.n5098 GND.n5097 9.3005
R14247 GND.n825 GND.n824 9.3005
R14248 GND.n5105 GND.n5104 9.3005
R14249 GND.n5106 GND.n823 9.3005
R14250 GND.n5108 GND.n5107 9.3005
R14251 GND.n819 GND.n818 9.3005
R14252 GND.n5115 GND.n5114 9.3005
R14253 GND.n5116 GND.n817 9.3005
R14254 GND.n5118 GND.n5117 9.3005
R14255 GND.n813 GND.n812 9.3005
R14256 GND.n5125 GND.n5124 9.3005
R14257 GND.n5126 GND.n811 9.3005
R14258 GND.n5128 GND.n5127 9.3005
R14259 GND.n807 GND.n806 9.3005
R14260 GND.n5135 GND.n5134 9.3005
R14261 GND.n5136 GND.n805 9.3005
R14262 GND.n5138 GND.n5137 9.3005
R14263 GND.n801 GND.n800 9.3005
R14264 GND.n5145 GND.n5144 9.3005
R14265 GND.n5146 GND.n799 9.3005
R14266 GND.n5148 GND.n5147 9.3005
R14267 GND.n795 GND.n794 9.3005
R14268 GND.n5155 GND.n5154 9.3005
R14269 GND.n5156 GND.n793 9.3005
R14270 GND.n5158 GND.n5157 9.3005
R14271 GND.n789 GND.n788 9.3005
R14272 GND.n5165 GND.n5164 9.3005
R14273 GND.n5166 GND.n787 9.3005
R14274 GND.n5168 GND.n5167 9.3005
R14275 GND.n783 GND.n782 9.3005
R14276 GND.n5175 GND.n5174 9.3005
R14277 GND.n5176 GND.n781 9.3005
R14278 GND.n5178 GND.n5177 9.3005
R14279 GND.n777 GND.n776 9.3005
R14280 GND.n5185 GND.n5184 9.3005
R14281 GND.n5186 GND.n775 9.3005
R14282 GND.n5188 GND.n5187 9.3005
R14283 GND.n771 GND.n770 9.3005
R14284 GND.n5195 GND.n5194 9.3005
R14285 GND.n5196 GND.n769 9.3005
R14286 GND.n5198 GND.n5197 9.3005
R14287 GND.n765 GND.n764 9.3005
R14288 GND.n5205 GND.n5204 9.3005
R14289 GND.n5206 GND.n763 9.3005
R14290 GND.n5208 GND.n5207 9.3005
R14291 GND.n759 GND.n758 9.3005
R14292 GND.n5215 GND.n5214 9.3005
R14293 GND.n5216 GND.n757 9.3005
R14294 GND.n5218 GND.n5217 9.3005
R14295 GND.n753 GND.n752 9.3005
R14296 GND.n5225 GND.n5224 9.3005
R14297 GND.n5226 GND.n751 9.3005
R14298 GND.n5228 GND.n5227 9.3005
R14299 GND.n747 GND.n746 9.3005
R14300 GND.n5235 GND.n5234 9.3005
R14301 GND.n5236 GND.n745 9.3005
R14302 GND.n5238 GND.n5237 9.3005
R14303 GND.n741 GND.n740 9.3005
R14304 GND.n5245 GND.n5244 9.3005
R14305 GND.n5246 GND.n739 9.3005
R14306 GND.n5248 GND.n5247 9.3005
R14307 GND.n735 GND.n734 9.3005
R14308 GND.n5255 GND.n5254 9.3005
R14309 GND.n5256 GND.n733 9.3005
R14310 GND.n5258 GND.n5257 9.3005
R14311 GND.n729 GND.n728 9.3005
R14312 GND.n5265 GND.n5264 9.3005
R14313 GND.n5266 GND.n727 9.3005
R14314 GND.n5268 GND.n5267 9.3005
R14315 GND.n723 GND.n722 9.3005
R14316 GND.n5275 GND.n5274 9.3005
R14317 GND.n5276 GND.n721 9.3005
R14318 GND.n5278 GND.n5277 9.3005
R14319 GND.n717 GND.n716 9.3005
R14320 GND.n5285 GND.n5284 9.3005
R14321 GND.n5286 GND.n715 9.3005
R14322 GND.n5288 GND.n5287 9.3005
R14323 GND.n711 GND.n710 9.3005
R14324 GND.n5295 GND.n5294 9.3005
R14325 GND.n5296 GND.n709 9.3005
R14326 GND.n5298 GND.n5297 9.3005
R14327 GND.n705 GND.n704 9.3005
R14328 GND.n5305 GND.n5304 9.3005
R14329 GND.n5306 GND.n703 9.3005
R14330 GND.n5309 GND.n5307 9.3005
R14331 GND.n5308 GND.n699 9.3005
R14332 GND.n5317 GND.n698 9.3005
R14333 GND.n5319 GND.n5318 9.3005
R14334 GND.n694 GND.n693 9.3005
R14335 GND.n5326 GND.n5325 9.3005
R14336 GND.n5327 GND.n692 9.3005
R14337 GND.n5329 GND.n5328 9.3005
R14338 GND.n688 GND.n687 9.3005
R14339 GND.n5336 GND.n5335 9.3005
R14340 GND.n5337 GND.n686 9.3005
R14341 GND.n5339 GND.n5338 9.3005
R14342 GND.n682 GND.n681 9.3005
R14343 GND.n5346 GND.n5345 9.3005
R14344 GND.n5347 GND.n680 9.3005
R14345 GND.n5349 GND.n5348 9.3005
R14346 GND.n676 GND.n675 9.3005
R14347 GND.n5356 GND.n5355 9.3005
R14348 GND.n5357 GND.n674 9.3005
R14349 GND.n5359 GND.n5358 9.3005
R14350 GND.n670 GND.n669 9.3005
R14351 GND.n5366 GND.n5365 9.3005
R14352 GND.n5367 GND.n668 9.3005
R14353 GND.n5369 GND.n5368 9.3005
R14354 GND.n664 GND.n663 9.3005
R14355 GND.n5376 GND.n5375 9.3005
R14356 GND.n5377 GND.n662 9.3005
R14357 GND.n5379 GND.n5378 9.3005
R14358 GND.n658 GND.n657 9.3005
R14359 GND.n5386 GND.n5385 9.3005
R14360 GND.n5387 GND.n656 9.3005
R14361 GND.n5389 GND.n5388 9.3005
R14362 GND.n652 GND.n651 9.3005
R14363 GND.n5396 GND.n5395 9.3005
R14364 GND.n5397 GND.n650 9.3005
R14365 GND.n5399 GND.n5398 9.3005
R14366 GND.n646 GND.n645 9.3005
R14367 GND.n5406 GND.n5405 9.3005
R14368 GND.n5407 GND.n644 9.3005
R14369 GND.n5409 GND.n5408 9.3005
R14370 GND.n640 GND.n639 9.3005
R14371 GND.n5416 GND.n5415 9.3005
R14372 GND.n5417 GND.n638 9.3005
R14373 GND.n5419 GND.n5418 9.3005
R14374 GND.n634 GND.n633 9.3005
R14375 GND.n5426 GND.n5425 9.3005
R14376 GND.n5427 GND.n632 9.3005
R14377 GND.n5429 GND.n5428 9.3005
R14378 GND.n628 GND.n627 9.3005
R14379 GND.n5436 GND.n5435 9.3005
R14380 GND.n5437 GND.n626 9.3005
R14381 GND.n5439 GND.n5438 9.3005
R14382 GND.n622 GND.n621 9.3005
R14383 GND.n5446 GND.n5445 9.3005
R14384 GND.n5447 GND.n620 9.3005
R14385 GND.n5449 GND.n5448 9.3005
R14386 GND.n616 GND.n615 9.3005
R14387 GND.n5456 GND.n5455 9.3005
R14388 GND.n5457 GND.n614 9.3005
R14389 GND.n5459 GND.n5458 9.3005
R14390 GND.n610 GND.n609 9.3005
R14391 GND.n5466 GND.n5465 9.3005
R14392 GND.n5467 GND.n608 9.3005
R14393 GND.n5469 GND.n5468 9.3005
R14394 GND.n604 GND.n603 9.3005
R14395 GND.n5476 GND.n5475 9.3005
R14396 GND.n5477 GND.n602 9.3005
R14397 GND.n5479 GND.n5478 9.3005
R14398 GND.n5316 GND.n5315 9.3005
R14399 GND.n3652 GND.n3651 9.3005
R14400 GND.n3653 GND.n3642 9.3005
R14401 GND.n3656 GND.n3641 9.3005
R14402 GND.n3657 GND.n3640 9.3005
R14403 GND.n3660 GND.n3639 9.3005
R14404 GND.n3661 GND.n3638 9.3005
R14405 GND.n3664 GND.n3637 9.3005
R14406 GND.n3665 GND.n3636 9.3005
R14407 GND.n3668 GND.n3635 9.3005
R14408 GND.n3669 GND.n3634 9.3005
R14409 GND.n3672 GND.n3633 9.3005
R14410 GND.n3673 GND.n3632 9.3005
R14411 GND.n3676 GND.n3631 9.3005
R14412 GND.n3677 GND.n3630 9.3005
R14413 GND.n3680 GND.n3629 9.3005
R14414 GND.n3681 GND.n3628 9.3005
R14415 GND.n3684 GND.n3627 9.3005
R14416 GND.n3623 GND.n3579 9.3005
R14417 GND.n3622 GND.n3621 9.3005
R14418 GND.n3618 GND.n3581 9.3005
R14419 GND.n3617 GND.n3614 9.3005
R14420 GND.n3613 GND.n3582 9.3005
R14421 GND.n3612 GND.n3611 9.3005
R14422 GND.n3608 GND.n3583 9.3005
R14423 GND.n3607 GND.n3604 9.3005
R14424 GND.n3603 GND.n3584 9.3005
R14425 GND.n3602 GND.n3601 9.3005
R14426 GND.n3598 GND.n3585 9.3005
R14427 GND.n3597 GND.n3594 9.3005
R14428 GND.n3593 GND.n3586 9.3005
R14429 GND.n3592 GND.n3591 9.3005
R14430 GND.n3650 GND.n3649 9.3005
R14431 GND.n3645 GND.n1854 9.3005
R14432 GND.n2110 GND.n2109 9.3005
R14433 GND.n3896 GND.n3895 9.3005
R14434 GND.n3897 GND.n2108 9.3005
R14435 GND.n3901 GND.n3898 9.3005
R14436 GND.n3900 GND.n3899 9.3005
R14437 GND.n2087 GND.n2086 9.3005
R14438 GND.n3920 GND.n3919 9.3005
R14439 GND.n3921 GND.n2085 9.3005
R14440 GND.n3925 GND.n3922 9.3005
R14441 GND.n3924 GND.n3923 9.3005
R14442 GND.n2066 GND.n2065 9.3005
R14443 GND.n3945 GND.n3944 9.3005
R14444 GND.n3946 GND.n2064 9.3005
R14445 GND.n3950 GND.n3947 9.3005
R14446 GND.n3949 GND.n3948 9.3005
R14447 GND.n2033 GND.n2032 9.3005
R14448 GND.n3985 GND.n3984 9.3005
R14449 GND.n3986 GND.n2031 9.3005
R14450 GND.n3988 GND.n3987 9.3005
R14451 GND.n3989 GND.n1994 9.3005
R14452 GND.n4069 GND.n4066 9.3005
R14453 GND.n4068 GND.n4067 9.3005
R14454 GND.n1972 GND.n1971 9.3005
R14455 GND.n4090 GND.n4089 9.3005
R14456 GND.n4091 GND.n1970 9.3005
R14457 GND.n4095 GND.n4092 9.3005
R14458 GND.n4094 GND.n4093 9.3005
R14459 GND.n1949 GND.n1948 9.3005
R14460 GND.n4123 GND.n4122 9.3005
R14461 GND.n4124 GND.n1947 9.3005
R14462 GND.n4128 GND.n4125 9.3005
R14463 GND.n4127 GND.n4126 9.3005
R14464 GND.n578 GND.n577 9.3005
R14465 GND.n5498 GND.n5497 9.3005
R14466 GND.n5499 GND.n576 9.3005
R14467 GND.n5501 GND.n5500 9.3005
R14468 GND.n560 GND.n559 9.3005
R14469 GND.n5516 GND.n5515 9.3005
R14470 GND.n5517 GND.n558 9.3005
R14471 GND.n5520 GND.n5518 9.3005
R14472 GND.n5519 GND.n497 9.3005
R14473 GND.n3588 GND.n3587 9.3005
R14474 GND.n4065 GND.n1993 9.3005
R14475 GND.n2799 GND.n2751 9.3005
R14476 GND.n2754 GND.n2752 9.3005
R14477 GND.n2793 GND.n2755 9.3005
R14478 GND.n2792 GND.n2756 9.3005
R14479 GND.n2791 GND.n2757 9.3005
R14480 GND.n2760 GND.n2758 9.3005
R14481 GND.n2784 GND.n2761 9.3005
R14482 GND.n2783 GND.n2762 9.3005
R14483 GND.n2782 GND.n2763 9.3005
R14484 GND.n2768 GND.n2764 9.3005
R14485 GND.n2778 GND.n2769 9.3005
R14486 GND.n2777 GND.n2770 9.3005
R14487 GND.n2776 GND.n2771 9.3005
R14488 GND.n2774 GND.n2773 9.3005
R14489 GND.n2772 GND.n2314 9.3005
R14490 GND.n2312 GND.n2311 9.3005
R14491 GND.n2916 GND.n2915 9.3005
R14492 GND.n2917 GND.n2310 9.3005
R14493 GND.n2928 GND.n2918 9.3005
R14494 GND.n2927 GND.n2919 9.3005
R14495 GND.n2926 GND.n2920 9.3005
R14496 GND.n2923 GND.n2922 9.3005
R14497 GND.n2921 GND.n1394 9.3005
R14498 GND.n4473 GND.n1395 9.3005
R14499 GND.n4472 GND.n1396 9.3005
R14500 GND.n4471 GND.n1397 9.3005
R14501 GND.n1418 GND.n1398 9.3005
R14502 GND.n1419 GND.n1400 9.3005
R14503 GND.n1421 GND.n1420 9.3005
R14504 GND.n1424 GND.n1423 9.3005
R14505 GND.n1425 GND.n1417 9.3005
R14506 GND.n4455 GND.n1426 9.3005
R14507 GND.n4454 GND.n1427 9.3005
R14508 GND.n4453 GND.n1428 9.3005
R14509 GND.n1451 GND.n1429 9.3005
R14510 GND.n1452 GND.n1450 9.3005
R14511 GND.n4441 GND.n1453 9.3005
R14512 GND.n4440 GND.n1454 9.3005
R14513 GND.n4439 GND.n1455 9.3005
R14514 GND.n1478 GND.n1456 9.3005
R14515 GND.n1479 GND.n1477 9.3005
R14516 GND.n4427 GND.n1480 9.3005
R14517 GND.n4426 GND.n1481 9.3005
R14518 GND.n4425 GND.n1482 9.3005
R14519 GND.n1496 GND.n1483 9.3005
R14520 GND.n4413 GND.n1497 9.3005
R14521 GND.n4412 GND.n1498 9.3005
R14522 GND.n4411 GND.n1499 9.3005
R14523 GND.n1514 GND.n1500 9.3005
R14524 GND.n4399 GND.n1515 9.3005
R14525 GND.n4398 GND.n1516 9.3005
R14526 GND.n4397 GND.n1517 9.3005
R14527 GND.n1534 GND.n1518 9.3005
R14528 GND.n4385 GND.n1535 9.3005
R14529 GND.n4384 GND.n1536 9.3005
R14530 GND.n4383 GND.n1537 9.3005
R14531 GND.n1565 GND.n1538 9.3005
R14532 GND.n1568 GND.n1567 9.3005
R14533 GND.n1569 GND.n1564 9.3005
R14534 GND.n4364 GND.n1570 9.3005
R14535 GND.n4363 GND.n1571 9.3005
R14536 GND.n4362 GND.n1572 9.3005
R14537 GND.n1608 GND.n1573 9.3005
R14538 GND.n1611 GND.n1610 9.3005
R14539 GND.n1612 GND.n1607 9.3005
R14540 GND.n4343 GND.n1613 9.3005
R14541 GND.n4342 GND.n1614 9.3005
R14542 GND.n4341 GND.n1615 9.3005
R14543 GND.n3411 GND.n1616 9.3005
R14544 GND.n3412 GND.n3410 9.3005
R14545 GND.n3415 GND.n3414 9.3005
R14546 GND.n3413 GND.n1656 9.3005
R14547 GND.n4316 GND.n1657 9.3005
R14548 GND.n4315 GND.n1658 9.3005
R14549 GND.n4314 GND.n1659 9.3005
R14550 GND.n3760 GND.n1660 9.3005
R14551 GND.n3762 GND.n3761 9.3005
R14552 GND.n3766 GND.n3765 9.3005
R14553 GND.n3767 GND.n3759 9.3005
R14554 GND.n3770 GND.n3769 9.3005
R14555 GND.n3768 GND.n1700 9.3005
R14556 GND.n4288 GND.n1701 9.3005
R14557 GND.n4287 GND.n1702 9.3005
R14558 GND.n4286 GND.n1703 9.3005
R14559 GND.n1726 GND.n1704 9.3005
R14560 GND.n1727 GND.n1725 9.3005
R14561 GND.n4274 GND.n1728 9.3005
R14562 GND.n4273 GND.n1729 9.3005
R14563 GND.n4272 GND.n1730 9.3005
R14564 GND.n1752 GND.n1731 9.3005
R14565 GND.n1753 GND.n1751 9.3005
R14566 GND.n4260 GND.n1754 9.3005
R14567 GND.n4259 GND.n1755 9.3005
R14568 GND.n4258 GND.n1756 9.3005
R14569 GND.n2123 GND.n1757 9.3005
R14570 GND.n2125 GND.n2124 9.3005
R14571 GND.n2130 GND.n2129 9.3005
R14572 GND.n2131 GND.n2122 9.3005
R14573 GND.n2133 GND.n2132 9.3005
R14574 GND.n2120 GND.n2119 9.3005
R14575 GND.n3847 GND.n3846 9.3005
R14576 GND.n3848 GND.n2118 9.3005
R14577 GND.n3886 GND.n3849 9.3005
R14578 GND.n3885 GND.n3850 9.3005
R14579 GND.n3884 GND.n3851 9.3005
R14580 GND.n3854 GND.n3852 9.3005
R14581 GND.n3880 GND.n3855 9.3005
R14582 GND.n3879 GND.n3856 9.3005
R14583 GND.n3878 GND.n3857 9.3005
R14584 GND.n3860 GND.n3858 9.3005
R14585 GND.n3872 GND.n3861 9.3005
R14586 GND.n3871 GND.n3862 9.3005
R14587 GND.n3870 GND.n3863 9.3005
R14588 GND.n3867 GND.n3864 9.3005
R14589 GND.n3866 GND.n3865 9.3005
R14590 GND.n2048 GND.n2047 9.3005
R14591 GND.n3968 GND.n3967 9.3005
R14592 GND.n3969 GND.n2046 9.3005
R14593 GND.n3975 GND.n3970 9.3005
R14594 GND.n3974 GND.n3971 9.3005
R14595 GND.n3973 GND.n3972 9.3005
R14596 GND.n4075 GND.n4074 9.3005
R14597 GND.n4076 GND.n1983 9.3005
R14598 GND.n4080 GND.n4077 9.3005
R14599 GND.n4079 GND.n4078 9.3005
R14600 GND.n1961 GND.n1960 9.3005
R14601 GND.n4101 GND.n4100 9.3005
R14602 GND.n4102 GND.n1959 9.3005
R14603 GND.n4113 GND.n4103 9.3005
R14604 GND.n4112 GND.n4104 9.3005
R14605 GND.n4111 GND.n4105 9.3005
R14606 GND.n4108 GND.n4107 9.3005
R14607 GND.n4106 GND.n597 9.3005
R14608 GND.n5484 GND.n598 9.3005
R14609 GND.n5483 GND.n599 9.3005
R14610 GND.n5482 GND.n600 9.3005
R14611 GND.n4687 GND.n4686 9.3005
R14612 GND.n4688 GND.n1148 9.3005
R14613 GND.n4691 GND.n1147 9.3005
R14614 GND.n4692 GND.n1146 9.3005
R14615 GND.n4695 GND.n1145 9.3005
R14616 GND.n4696 GND.n1144 9.3005
R14617 GND.n4699 GND.n1143 9.3005
R14618 GND.n4700 GND.n1142 9.3005
R14619 GND.n4703 GND.n1141 9.3005
R14620 GND.n4704 GND.n1140 9.3005
R14621 GND.n4707 GND.n1139 9.3005
R14622 GND.n4708 GND.n1138 9.3005
R14623 GND.n4711 GND.n1137 9.3005
R14624 GND.n4712 GND.n1136 9.3005
R14625 GND.n4715 GND.n1135 9.3005
R14626 GND.n4716 GND.n1134 9.3005
R14627 GND.n4719 GND.n1133 9.3005
R14628 GND.n4721 GND.n1130 9.3005
R14629 GND.n4724 GND.n1129 9.3005
R14630 GND.n4725 GND.n1128 9.3005
R14631 GND.n4728 GND.n1127 9.3005
R14632 GND.n4729 GND.n1126 9.3005
R14633 GND.n4732 GND.n1125 9.3005
R14634 GND.n4733 GND.n1124 9.3005
R14635 GND.n4736 GND.n1123 9.3005
R14636 GND.n4737 GND.n1122 9.3005
R14637 GND.n4740 GND.n1121 9.3005
R14638 GND.n4741 GND.n1120 9.3005
R14639 GND.n4744 GND.n1119 9.3005
R14640 GND.n4746 GND.n1118 9.3005
R14641 GND.n4747 GND.n1117 9.3005
R14642 GND.n4748 GND.n1116 9.3005
R14643 GND.n4749 GND.n1115 9.3005
R14644 GND.n4685 GND.n1153 9.3005
R14645 GND.n4684 GND.n4683 9.3005
R14646 GND.n2550 GND.n2547 9.3005
R14647 GND.n2622 GND.n2621 9.3005
R14648 GND.n2623 GND.n2546 9.3005
R14649 GND.n2627 GND.n2624 9.3005
R14650 GND.n2626 GND.n2625 9.3005
R14651 GND.n2490 GND.n2489 9.3005
R14652 GND.n2647 GND.n2646 9.3005
R14653 GND.n2648 GND.n2488 9.3005
R14654 GND.n2652 GND.n2649 9.3005
R14655 GND.n2651 GND.n2650 9.3005
R14656 GND.n2467 GND.n2466 9.3005
R14657 GND.n2672 GND.n2671 9.3005
R14658 GND.n2673 GND.n2465 9.3005
R14659 GND.n2677 GND.n2674 9.3005
R14660 GND.n2676 GND.n2675 9.3005
R14661 GND.n2444 GND.n2443 9.3005
R14662 GND.n2709 GND.n2708 9.3005
R14663 GND.n2710 GND.n2442 9.3005
R14664 GND.n2713 GND.n2711 9.3005
R14665 GND.n2712 GND.n2380 9.3005
R14666 GND.n2833 GND.n2832 9.3005
R14667 GND.n2360 GND.n2359 9.3005
R14668 GND.n2854 GND.n2853 9.3005
R14669 GND.n2855 GND.n2358 9.3005
R14670 GND.n2859 GND.n2856 9.3005
R14671 GND.n2858 GND.n2857 9.3005
R14672 GND.n2341 GND.n2340 9.3005
R14673 GND.n2879 GND.n2878 9.3005
R14674 GND.n2880 GND.n2339 9.3005
R14675 GND.n2884 GND.n2881 9.3005
R14676 GND.n2883 GND.n2882 9.3005
R14677 GND.n2320 GND.n2319 9.3005
R14678 GND.n2905 GND.n2904 9.3005
R14679 GND.n2906 GND.n2318 9.3005
R14680 GND.n2908 GND.n2907 9.3005
R14681 GND.n2294 GND.n2293 9.3005
R14682 GND.n2945 GND.n2944 9.3005
R14683 GND.n2946 GND.n2292 9.3005
R14684 GND.n2948 GND.n2947 9.3005
R14685 GND.n1268 GND.n1267 9.3005
R14686 GND.n4598 GND.n4597 9.3005
R14687 GND.n2549 GND.n2548 9.3005
R14688 GND.n2834 GND.n2831 9.3005
R14689 GND.n2536 GND.n2507 9.3005
R14690 GND.n2510 GND.n2508 9.3005
R14691 GND.n2532 GND.n2511 9.3005
R14692 GND.n2531 GND.n2512 9.3005
R14693 GND.n2530 GND.n2513 9.3005
R14694 GND.n2516 GND.n2514 9.3005
R14695 GND.n2526 GND.n2517 9.3005
R14696 GND.n2525 GND.n2518 9.3005
R14697 GND.n2524 GND.n2519 9.3005
R14698 GND.n2521 GND.n2520 9.3005
R14699 GND.n2432 GND.n2431 9.3005
R14700 GND.n2719 GND.n2718 9.3005
R14701 GND.n2720 GND.n2430 9.3005
R14702 GND.n2722 GND.n2721 9.3005
R14703 GND.n2538 GND.n2537 9.3005
R14704 GND.n2506 GND.n1084 9.3005
R14705 GND.n4756 GND.n1083 9.3005
R14706 GND.n4757 GND.n1082 9.3005
R14707 GND.n4758 GND.n1081 9.3005
R14708 GND.n1080 GND.n1076 9.3005
R14709 GND.n4764 GND.n1075 9.3005
R14710 GND.n4765 GND.n1074 9.3005
R14711 GND.n4766 GND.n1073 9.3005
R14712 GND.n1072 GND.n1068 9.3005
R14713 GND.n4772 GND.n1067 9.3005
R14714 GND.n4773 GND.n1066 9.3005
R14715 GND.n4774 GND.n1065 9.3005
R14716 GND.n1064 GND.n1060 9.3005
R14717 GND.n4780 GND.n1059 9.3005
R14718 GND.n4781 GND.n1058 9.3005
R14719 GND.n4782 GND.n1057 9.3005
R14720 GND.n1056 GND.n1052 9.3005
R14721 GND.n4788 GND.n1051 9.3005
R14722 GND.n4789 GND.n1050 9.3005
R14723 GND.n4790 GND.n1049 9.3005
R14724 GND.n1048 GND.n1044 9.3005
R14725 GND.n4796 GND.n1043 9.3005
R14726 GND.n4797 GND.n1042 9.3005
R14727 GND.n4798 GND.n1041 9.3005
R14728 GND.n1040 GND.n1036 9.3005
R14729 GND.n4804 GND.n1035 9.3005
R14730 GND.n4805 GND.n1034 9.3005
R14731 GND.n4806 GND.n1033 9.3005
R14732 GND.n1032 GND.n1028 9.3005
R14733 GND.n4812 GND.n1027 9.3005
R14734 GND.n4813 GND.n1026 9.3005
R14735 GND.n4814 GND.n1025 9.3005
R14736 GND.n1024 GND.n1020 9.3005
R14737 GND.n4820 GND.n1019 9.3005
R14738 GND.n4821 GND.n1018 9.3005
R14739 GND.n4822 GND.n1017 9.3005
R14740 GND.n1016 GND.n1012 9.3005
R14741 GND.n4828 GND.n1011 9.3005
R14742 GND.n4829 GND.n1010 9.3005
R14743 GND.n4830 GND.n1009 9.3005
R14744 GND.n1008 GND.n1004 9.3005
R14745 GND.n4836 GND.n1003 9.3005
R14746 GND.n4837 GND.n1002 9.3005
R14747 GND.n4838 GND.n1001 9.3005
R14748 GND.n1000 GND.n996 9.3005
R14749 GND.n4844 GND.n995 9.3005
R14750 GND.n4845 GND.n994 9.3005
R14751 GND.n4846 GND.n993 9.3005
R14752 GND.n992 GND.n988 9.3005
R14753 GND.n4852 GND.n987 9.3005
R14754 GND.n4853 GND.n986 9.3005
R14755 GND.n4854 GND.n985 9.3005
R14756 GND.n984 GND.n980 9.3005
R14757 GND.n4860 GND.n979 9.3005
R14758 GND.n4861 GND.n978 9.3005
R14759 GND.n4862 GND.n977 9.3005
R14760 GND.n976 GND.n972 9.3005
R14761 GND.n4868 GND.n971 9.3005
R14762 GND.n4869 GND.n970 9.3005
R14763 GND.n4870 GND.n969 9.3005
R14764 GND.n968 GND.n964 9.3005
R14765 GND.n4876 GND.n963 9.3005
R14766 GND.n4877 GND.n962 9.3005
R14767 GND.n4878 GND.n961 9.3005
R14768 GND.n957 GND.n956 9.3005
R14769 GND.n4885 GND.n4884 9.3005
R14770 GND.n2540 GND.n2539 9.3005
R14771 GND.n3841 GND.n3840 9.3005
R14772 GND.n3839 GND.n2139 9.3005
R14773 GND.n2100 GND.n2099 9.3005
R14774 GND.n3906 GND.n3905 9.3005
R14775 GND.n3907 GND.n2097 9.3005
R14776 GND.n3910 GND.n3909 9.3005
R14777 GND.n3908 GND.n2098 9.3005
R14778 GND.n2078 GND.n2077 9.3005
R14779 GND.n3930 GND.n3929 9.3005
R14780 GND.n3931 GND.n2075 9.3005
R14781 GND.n3934 GND.n3933 9.3005
R14782 GND.n3932 GND.n2076 9.3005
R14783 GND.n2056 GND.n2055 9.3005
R14784 GND.n3955 GND.n3954 9.3005
R14785 GND.n3956 GND.n2053 9.3005
R14786 GND.n3961 GND.n3960 9.3005
R14787 GND.n3959 GND.n2054 9.3005
R14788 GND.n3958 GND.n3957 9.3005
R14789 GND.n2022 GND.n2021 9.3005
R14790 GND.n3994 GND.n3993 9.3005
R14791 GND.n3995 GND.n2019 9.3005
R14792 GND.n4000 GND.n3999 9.3005
R14793 GND.n3998 GND.n2020 9.3005
R14794 GND.n3997 GND.n3996 9.3005
R14795 GND.n428 GND.n426 9.3005
R14796 GND.n3838 GND.n2138 9.3005
R14797 GND.n5674 GND.n5673 9.3005
R14798 GND.n5672 GND.n427 9.3005
R14799 GND.n5671 GND.n5670 9.3005
R14800 GND.n5669 GND.n432 9.3005
R14801 GND.n5668 GND.n5667 9.3005
R14802 GND.n5666 GND.n433 9.3005
R14803 GND.n5665 GND.n5664 9.3005
R14804 GND.n5663 GND.n437 9.3005
R14805 GND.n5662 GND.n5661 9.3005
R14806 GND.n5660 GND.n438 9.3005
R14807 GND.n5659 GND.n5658 9.3005
R14808 GND.n5657 GND.n442 9.3005
R14809 GND.n5656 GND.n5655 9.3005
R14810 GND.n5654 GND.n443 9.3005
R14811 GND.n5653 GND.n5652 9.3005
R14812 GND.n5651 GND.n447 9.3005
R14813 GND.n5650 GND.n5649 9.3005
R14814 GND.n5648 GND.n448 9.3005
R14815 GND.n5647 GND.n5646 9.3005
R14816 GND.n5645 GND.n452 9.3005
R14817 GND.n5644 GND.n5643 9.3005
R14818 GND.n5642 GND.n453 9.3005
R14819 GND.n5641 GND.n5640 9.3005
R14820 GND.n5639 GND.n457 9.3005
R14821 GND.n5638 GND.n5637 9.3005
R14822 GND.n5636 GND.n458 9.3005
R14823 GND.n5635 GND.n5634 9.3005
R14824 GND.n5565 GND.n5524 9.3005
R14825 GND.n5564 GND.n5563 9.3005
R14826 GND.n5562 GND.n5525 9.3005
R14827 GND.n5561 GND.n5560 9.3005
R14828 GND.n5559 GND.n5530 9.3005
R14829 GND.n5558 GND.n5557 9.3005
R14830 GND.n5556 GND.n5531 9.3005
R14831 GND.n5555 GND.n5554 9.3005
R14832 GND.n5553 GND.n5536 9.3005
R14833 GND.n5552 GND.n5551 9.3005
R14834 GND.n5550 GND.n5537 9.3005
R14835 GND.n5549 GND.n5548 9.3005
R14836 GND.n5547 GND.n5542 9.3005
R14837 GND.n5546 GND.n5545 9.3005
R14838 GND.n465 GND.n462 9.3005
R14839 GND.n5633 GND.n5632 9.3005
R14840 GND.n5567 GND.n5566 9.3005
R14841 GND.n5626 GND.n496 9.3005
R14842 GND.n5625 GND.n5624 9.3005
R14843 GND.n5623 GND.n498 9.3005
R14844 GND.n5622 GND.n5621 9.3005
R14845 GND.n5620 GND.n503 9.3005
R14846 GND.n5619 GND.n5618 9.3005
R14847 GND.n5617 GND.n504 9.3005
R14848 GND.n5616 GND.n5615 9.3005
R14849 GND.n5614 GND.n509 9.3005
R14850 GND.n5613 GND.n5612 9.3005
R14851 GND.n5611 GND.n510 9.3005
R14852 GND.n5610 GND.n5609 9.3005
R14853 GND.n5608 GND.n515 9.3005
R14854 GND.n5607 GND.n5606 9.3005
R14855 GND.n5605 GND.n516 9.3005
R14856 GND.n5603 GND.n5602 9.3005
R14857 GND.n5601 GND.n523 9.3005
R14858 GND.n5600 GND.n5599 9.3005
R14859 GND.n5598 GND.n524 9.3005
R14860 GND.n5597 GND.n5596 9.3005
R14861 GND.n5595 GND.n529 9.3005
R14862 GND.n5594 GND.n5593 9.3005
R14863 GND.n5592 GND.n530 9.3005
R14864 GND.n5591 GND.n5590 9.3005
R14865 GND.n5589 GND.n535 9.3005
R14866 GND.n5588 GND.n5587 9.3005
R14867 GND.n5586 GND.n536 9.3005
R14868 GND.n5585 GND.n5584 9.3005
R14869 GND.n5583 GND.n541 9.3005
R14870 GND.n5582 GND.n5581 9.3005
R14871 GND.n5580 GND.n542 9.3005
R14872 GND.n5579 GND.n5578 9.3005
R14873 GND.n5577 GND.n549 9.3005
R14874 GND.n5576 GND.n5575 9.3005
R14875 GND.n5628 GND.n5627 9.3005
R14876 GND.n2114 GND.n1856 9.3005
R14877 GND.n4195 GND.n1861 9.3005
R14878 GND.n4194 GND.n1862 9.3005
R14879 GND.n4193 GND.n1863 9.3005
R14880 GND.n2093 GND.n1864 9.3005
R14881 GND.n4189 GND.n1869 9.3005
R14882 GND.n4188 GND.n1870 9.3005
R14883 GND.n4187 GND.n1871 9.3005
R14884 GND.n2081 GND.n1872 9.3005
R14885 GND.n4183 GND.n1877 9.3005
R14886 GND.n4182 GND.n1878 9.3005
R14887 GND.n4181 GND.n1879 9.3005
R14888 GND.n3938 GND.n1880 9.3005
R14889 GND.n4177 GND.n1885 9.3005
R14890 GND.n4176 GND.n1886 9.3005
R14891 GND.n4175 GND.n1887 9.3005
R14892 GND.n3980 GND.n1888 9.3005
R14893 GND.n4171 GND.n1893 9.3005
R14894 GND.n4170 GND.n1894 9.3005
R14895 GND.n4169 GND.n1895 9.3005
R14896 GND.n2026 GND.n1896 9.3005
R14897 GND.n4165 GND.n1901 9.3005
R14898 GND.n4164 GND.n1902 9.3005
R14899 GND.n4163 GND.n1903 9.3005
R14900 GND.n2006 GND.n1904 9.3005
R14901 GND.n4159 GND.n1909 9.3005
R14902 GND.n4158 GND.n1910 9.3005
R14903 GND.n4157 GND.n1911 9.3005
R14904 GND.n4026 GND.n1912 9.3005
R14905 GND.n4153 GND.n1917 9.3005
R14906 GND.n4152 GND.n1918 9.3005
R14907 GND.n4151 GND.n1919 9.3005
R14908 GND.n1977 GND.n1920 9.3005
R14909 GND.n4147 GND.n1925 9.3005
R14910 GND.n4146 GND.n1926 9.3005
R14911 GND.n4145 GND.n1927 9.3005
R14912 GND.n1966 GND.n1928 9.3005
R14913 GND.n4141 GND.n1933 9.3005
R14914 GND.n4140 GND.n1934 9.3005
R14915 GND.n4139 GND.n1935 9.3005
R14916 GND.n1941 GND.n1936 9.3005
R14917 GND.n4135 GND.n1940 9.3005
R14918 GND.n4134 GND.n4133 9.3005
R14919 GND.n588 GND.n586 9.3005
R14920 GND.n5493 GND.n5492 9.3005
R14921 GND.n591 GND.n587 9.3005
R14922 GND.n590 GND.n589 9.3005
R14923 GND.n568 GND.n566 9.3005
R14924 GND.n5511 GND.n5510 9.3005
R14925 GND.n569 GND.n567 9.3005
R14926 GND.n554 GND.n553 9.3005
R14927 GND.n5571 GND.n5570 9.3005
R14928 GND.n4199 GND.n1855 9.3005
R14929 GND.n4197 GND.n1856 9.3005
R14930 GND.n4196 GND.n4195 9.3005
R14931 GND.n4194 GND.n1860 9.3005
R14932 GND.n4193 GND.n4192 9.3005
R14933 GND.n4191 GND.n1864 9.3005
R14934 GND.n4190 GND.n4189 9.3005
R14935 GND.n4188 GND.n1868 9.3005
R14936 GND.n4187 GND.n4186 9.3005
R14937 GND.n4185 GND.n1872 9.3005
R14938 GND.n4184 GND.n4183 9.3005
R14939 GND.n4182 GND.n1876 9.3005
R14940 GND.n4181 GND.n4180 9.3005
R14941 GND.n4179 GND.n1880 9.3005
R14942 GND.n4178 GND.n4177 9.3005
R14943 GND.n4176 GND.n1884 9.3005
R14944 GND.n4175 GND.n4174 9.3005
R14945 GND.n4173 GND.n1888 9.3005
R14946 GND.n4172 GND.n4171 9.3005
R14947 GND.n4170 GND.n1892 9.3005
R14948 GND.n4169 GND.n4168 9.3005
R14949 GND.n4167 GND.n1896 9.3005
R14950 GND.n4166 GND.n4165 9.3005
R14951 GND.n4164 GND.n1900 9.3005
R14952 GND.n4163 GND.n4162 9.3005
R14953 GND.n4161 GND.n1904 9.3005
R14954 GND.n4160 GND.n4159 9.3005
R14955 GND.n4158 GND.n1908 9.3005
R14956 GND.n4157 GND.n4156 9.3005
R14957 GND.n4155 GND.n1912 9.3005
R14958 GND.n4154 GND.n4153 9.3005
R14959 GND.n4152 GND.n1916 9.3005
R14960 GND.n4151 GND.n4150 9.3005
R14961 GND.n4149 GND.n1920 9.3005
R14962 GND.n4148 GND.n4147 9.3005
R14963 GND.n4146 GND.n1924 9.3005
R14964 GND.n4145 GND.n4144 9.3005
R14965 GND.n4143 GND.n1928 9.3005
R14966 GND.n4142 GND.n4141 9.3005
R14967 GND.n4140 GND.n1932 9.3005
R14968 GND.n4139 GND.n4138 9.3005
R14969 GND.n4137 GND.n1936 9.3005
R14970 GND.n4136 GND.n4135 9.3005
R14971 GND.n4134 GND.n592 9.3005
R14972 GND.n5489 GND.n588 9.3005
R14973 GND.n5492 GND.n5491 9.3005
R14974 GND.n5490 GND.n591 9.3005
R14975 GND.n590 GND.n570 9.3005
R14976 GND.n5506 GND.n568 9.3005
R14977 GND.n5510 GND.n5509 9.3005
R14978 GND.n5508 GND.n569 9.3005
R14979 GND.n553 GND.n552 9.3005
R14980 GND.n5572 GND.n5571 9.3005
R14981 GND.n4199 GND.n4198 9.3005
R14982 GND.n4211 GND.n4210 9.3005
R14983 GND.n4212 GND.n4201 9.3005
R14984 GND.n1780 GND.n1778 9.3005
R14985 GND.n4246 GND.n4245 9.3005
R14986 GND.n4244 GND.n4243 9.3005
R14987 GND.n1789 GND.n1788 9.3005
R14988 GND.n4238 GND.n4237 9.3005
R14989 GND.n4236 GND.n4235 9.3005
R14990 GND.n1799 GND.n1798 9.3005
R14991 GND.n4230 GND.n4229 9.3005
R14992 GND.n4228 GND.n4227 9.3005
R14993 GND.n1807 GND.n1806 9.3005
R14994 GND.n4222 GND.n4221 9.3005
R14995 GND.n4220 GND.n4219 9.3005
R14996 GND.n1819 GND.n1818 9.3005
R14997 GND.n2142 GND.n2140 9.3005
R14998 GND.n4252 GND.n4251 9.3005
R14999 GND.n4224 GND.n4223 9.3005
R15000 GND.n4226 GND.n4225 9.3005
R15001 GND.n1803 GND.n1802 9.3005
R15002 GND.n4232 GND.n4231 9.3005
R15003 GND.n4234 GND.n4233 9.3005
R15004 GND.n1793 GND.n1792 9.3005
R15005 GND.n4240 GND.n4239 9.3005
R15006 GND.n4242 GND.n4241 9.3005
R15007 GND.n1785 GND.n1784 9.3005
R15008 GND.n4248 GND.n4247 9.3005
R15009 GND.n4250 GND.n4249 9.3005
R15010 GND.n1781 GND.n1779 9.3005
R15011 GND.n4208 GND.n4204 9.3005
R15012 GND.n1813 GND.n1812 9.3005
R15013 GND.n4218 GND.n4217 9.3005
R15014 GND.n3836 GND.n3835 9.3005
R15015 GND.n3834 GND.n2141 9.3005
R15016 GND.n3833 GND.n3832 9.3005
R15017 GND.n3831 GND.n2147 9.3005
R15018 GND.n3830 GND.n3829 9.3005
R15019 GND.n3828 GND.n2148 9.3005
R15020 GND.n3827 GND.n3826 9.3005
R15021 GND.n3825 GND.n2153 9.3005
R15022 GND.n3824 GND.n3823 9.3005
R15023 GND.n3822 GND.n2154 9.3005
R15024 GND.n3820 GND.n3819 9.3005
R15025 GND.n3818 GND.n2161 9.3005
R15026 GND.n3817 GND.n3816 9.3005
R15027 GND.n3815 GND.n2162 9.3005
R15028 GND.n3004 GND.n2274 9.3005
R15029 GND.n3008 GND.n3007 9.3005
R15030 GND.n3009 GND.n2273 9.3005
R15031 GND.n3011 GND.n3010 9.3005
R15032 GND.n3014 GND.n2272 9.3005
R15033 GND.n3016 GND.n3015 9.3005
R15034 GND.n3017 GND.n2271 9.3005
R15035 GND.n3019 GND.n3018 9.3005
R15036 GND.n3020 GND.n2268 9.3005
R15037 GND.n3024 GND.n3023 9.3005
R15038 GND.n3025 GND.n2266 9.3005
R15039 GND.n3033 GND.n3032 9.3005
R15040 GND.n3031 GND.n2267 9.3005
R15041 GND.n3030 GND.n3029 9.3005
R15042 GND.n3028 GND.n3026 9.3005
R15043 GND.n2238 GND.n2237 9.3005
R15044 GND.n3251 GND.n3250 9.3005
R15045 GND.n3252 GND.n2235 9.3005
R15046 GND.n3270 GND.n3269 9.3005
R15047 GND.n3268 GND.n2236 9.3005
R15048 GND.n3267 GND.n3266 9.3005
R15049 GND.n3265 GND.n3253 9.3005
R15050 GND.n3264 GND.n3263 9.3005
R15051 GND.n3262 GND.n3258 9.3005
R15052 GND.n3261 GND.n3260 9.3005
R15053 GND.n2214 GND.n2213 9.3005
R15054 GND.n3323 GND.n3322 9.3005
R15055 GND.n3324 GND.n2211 9.3005
R15056 GND.n3347 GND.n3346 9.3005
R15057 GND.n3345 GND.n2212 9.3005
R15058 GND.n3344 GND.n3343 9.3005
R15059 GND.n3342 GND.n3325 9.3005
R15060 GND.n3341 GND.n3340 9.3005
R15061 GND.n3339 GND.n3330 9.3005
R15062 GND.n3338 GND.n3337 9.3005
R15063 GND.n3336 GND.n3331 9.3005
R15064 GND.n3335 GND.n3334 9.3005
R15065 GND.n3333 GND.n2197 9.3005
R15066 GND.n2196 GND.n2195 9.3005
R15067 GND.n3399 GND.n3398 9.3005
R15068 GND.n3400 GND.n2193 9.3005
R15069 GND.n3406 GND.n3405 9.3005
R15070 GND.n3404 GND.n2194 9.3005
R15071 GND.n3403 GND.n3402 9.3005
R15072 GND.n2184 GND.n2183 9.3005
R15073 GND.n3444 GND.n3443 9.3005
R15074 GND.n3445 GND.n2182 9.3005
R15075 GND.n3448 GND.n3447 9.3005
R15076 GND.n3446 GND.n2176 9.3005
R15077 GND.n3782 GND.n2175 9.3005
R15078 GND.n3784 GND.n3783 9.3005
R15079 GND.n3785 GND.n2174 9.3005
R15080 GND.n3787 GND.n3786 9.3005
R15081 GND.n3788 GND.n2173 9.3005
R15082 GND.n3792 GND.n3791 9.3005
R15083 GND.n3793 GND.n2170 9.3005
R15084 GND.n3795 GND.n3794 9.3005
R15085 GND.n3796 GND.n2169 9.3005
R15086 GND.n3800 GND.n3799 9.3005
R15087 GND.n3801 GND.n2168 9.3005
R15088 GND.n3803 GND.n3802 9.3005
R15089 GND.n3807 GND.n2167 9.3005
R15090 GND.n3809 GND.n3808 9.3005
R15091 GND.n3810 GND.n2166 9.3005
R15092 GND.n3812 GND.n3811 9.3005
R15093 GND.n3003 GND.n3002 9.3005
R15094 GND.n2998 GND.n2275 9.3005
R15095 GND.n2995 GND.n2994 9.3005
R15096 GND.n2993 GND.n2276 9.3005
R15097 GND.n2992 GND.n2991 9.3005
R15098 GND.n2985 GND.n2277 9.3005
R15099 GND.n2982 GND.n2981 9.3005
R15100 GND.n2980 GND.n2278 9.3005
R15101 GND.n2979 GND.n2978 9.3005
R15102 GND.n2975 GND.n2279 9.3005
R15103 GND.n2972 GND.n2971 9.3005
R15104 GND.n2970 GND.n2280 9.3005
R15105 GND.n2969 GND.n2968 9.3005
R15106 GND.n2965 GND.n2281 9.3005
R15107 GND.n3001 GND.n3000 9.3005
R15108 GND.n2741 GND.n2740 9.3005
R15109 GND.n2742 GND.n2420 9.3005
R15110 GND.n2744 GND.n2743 9.3005
R15111 GND.n2371 GND.n2370 9.3005
R15112 GND.n2839 GND.n2838 9.3005
R15113 GND.n2840 GND.n2368 9.3005
R15114 GND.n2843 GND.n2842 9.3005
R15115 GND.n2841 GND.n2369 9.3005
R15116 GND.n2351 GND.n2350 9.3005
R15117 GND.n2864 GND.n2863 9.3005
R15118 GND.n2865 GND.n2348 9.3005
R15119 GND.n2868 GND.n2867 9.3005
R15120 GND.n2866 GND.n2349 9.3005
R15121 GND.n2331 GND.n2330 9.3005
R15122 GND.n2889 GND.n2888 9.3005
R15123 GND.n2890 GND.n2328 9.3005
R15124 GND.n2896 GND.n2895 9.3005
R15125 GND.n2894 GND.n2329 9.3005
R15126 GND.n2893 GND.n2892 9.3005
R15127 GND.n2305 GND.n2303 9.3005
R15128 GND.n2937 GND.n2936 9.3005
R15129 GND.n2935 GND.n2304 9.3005
R15130 GND.n2934 GND.n2933 9.3005
R15131 GND.n2306 GND.n2287 9.3005
R15132 GND.n2957 GND.n2286 9.3005
R15133 GND.n2959 GND.n2958 9.3005
R15134 GND.n2962 GND.n2961 9.3005
R15135 GND.n2285 GND.n2284 9.3005
R15136 GND.n1371 GND.n1370 9.3005
R15137 GND.n4508 GND.n4507 9.3005
R15138 GND.n4510 GND.n4509 9.3005
R15139 GND.n1363 GND.n1362 9.3005
R15140 GND.n4516 GND.n4515 9.3005
R15141 GND.n4518 GND.n4517 9.3005
R15142 GND.n1353 GND.n1352 9.3005
R15143 GND.n4524 GND.n4523 9.3005
R15144 GND.n4526 GND.n4525 9.3005
R15145 GND.n1344 GND.n1341 9.3005
R15146 GND.n4532 GND.n4531 9.3005
R15147 GND.n1342 GND.n1322 9.3005
R15148 GND.n4538 GND.n4537 9.3005
R15149 GND.n4541 GND.n4540 9.3005
R15150 GND.n4539 GND.n1319 9.3005
R15151 GND.n1380 GND.n1321 9.3005
R15152 GND.n1345 GND.n1343 9.3005
R15153 GND.n4530 GND.n4529 9.3005
R15154 GND.n4528 GND.n4527 9.3005
R15155 GND.n1349 GND.n1348 9.3005
R15156 GND.n4522 GND.n4521 9.3005
R15157 GND.n4520 GND.n4519 9.3005
R15158 GND.n1357 GND.n1356 9.3005
R15159 GND.n4514 GND.n4513 9.3005
R15160 GND.n4512 GND.n4511 9.3005
R15161 GND.n1367 GND.n1366 9.3005
R15162 GND.n4506 GND.n4505 9.3005
R15163 GND.n4504 GND.n1375 9.3005
R15164 GND.n4542 GND.n1315 9.3005
R15165 GND.n4544 GND.n4543 9.3005
R15166 GND.n4576 GND.n1283 9.3005
R15167 GND.n4578 GND.n4577 9.3005
R15168 GND.n4579 GND.n1282 9.3005
R15169 GND.n4581 GND.n4580 9.3005
R15170 GND.n4582 GND.n1278 9.3005
R15171 GND.n4584 GND.n4583 9.3005
R15172 GND.n4585 GND.n1277 9.3005
R15173 GND.n4587 GND.n4586 9.3005
R15174 GND.n4588 GND.n1273 9.3005
R15175 GND.n4590 GND.n4589 9.3005
R15176 GND.n4591 GND.n1272 9.3005
R15177 GND.n4593 GND.n4592 9.3005
R15178 GND.n4594 GND.n1269 9.3005
R15179 GND.n4596 GND.n4595 9.3005
R15180 GND.n4572 GND.n1292 9.3005
R15181 GND.n4571 GND.n4570 9.3005
R15182 GND.n4569 GND.n1293 9.3005
R15183 GND.n4568 GND.n4567 9.3005
R15184 GND.n4566 GND.n1297 9.3005
R15185 GND.n4565 GND.n4564 9.3005
R15186 GND.n4563 GND.n1298 9.3005
R15187 GND.n4562 GND.n4561 9.3005
R15188 GND.n4560 GND.n1302 9.3005
R15189 GND.n4559 GND.n4558 9.3005
R15190 GND.n4557 GND.n1303 9.3005
R15191 GND.n4556 GND.n4555 9.3005
R15192 GND.n4554 GND.n1307 9.3005
R15193 GND.n4553 GND.n4552 9.3005
R15194 GND.n4551 GND.n1308 9.3005
R15195 GND.n4550 GND.n4549 9.3005
R15196 GND.n4548 GND.n1314 9.3005
R15197 GND.n4547 GND.n4546 9.3005
R15198 GND.n4574 GND.n4573 9.3005
R15199 GND.n4678 GND.n1158 9.3005
R15200 GND.n4677 GND.n1159 9.3005
R15201 GND.n2616 GND.n1160 9.3005
R15202 GND.n4673 GND.n1165 9.3005
R15203 GND.n4672 GND.n1166 9.3005
R15204 GND.n4671 GND.n1167 9.3005
R15205 GND.n2642 GND.n1168 9.3005
R15206 GND.n4667 GND.n1173 9.3005
R15207 GND.n4666 GND.n1174 9.3005
R15208 GND.n4665 GND.n1175 9.3005
R15209 GND.n2473 GND.n1176 9.3005
R15210 GND.n4661 GND.n1181 9.3005
R15211 GND.n4660 GND.n1182 9.3005
R15212 GND.n4659 GND.n1183 9.3005
R15213 GND.n2450 GND.n1184 9.3005
R15214 GND.n4655 GND.n1189 9.3005
R15215 GND.n4654 GND.n1190 9.3005
R15216 GND.n4653 GND.n1191 9.3005
R15217 GND.n2437 GND.n1192 9.3005
R15218 GND.n4649 GND.n1197 9.3005
R15219 GND.n4648 GND.n1198 9.3005
R15220 GND.n4647 GND.n1199 9.3005
R15221 GND.n2824 GND.n1200 9.3005
R15222 GND.n4643 GND.n1205 9.3005
R15223 GND.n4642 GND.n1206 9.3005
R15224 GND.n4641 GND.n1207 9.3005
R15225 GND.n2407 GND.n1208 9.3005
R15226 GND.n4637 GND.n1213 9.3005
R15227 GND.n4636 GND.n1214 9.3005
R15228 GND.n4635 GND.n1215 9.3005
R15229 GND.n2375 GND.n1216 9.3005
R15230 GND.n4631 GND.n1221 9.3005
R15231 GND.n4630 GND.n1222 9.3005
R15232 GND.n4629 GND.n1223 9.3005
R15233 GND.n2847 GND.n1224 9.3005
R15234 GND.n4625 GND.n1229 9.3005
R15235 GND.n4624 GND.n1230 9.3005
R15236 GND.n4623 GND.n1231 9.3005
R15237 GND.n2874 GND.n1232 9.3005
R15238 GND.n4619 GND.n1237 9.3005
R15239 GND.n4618 GND.n1238 9.3005
R15240 GND.n4617 GND.n1239 9.3005
R15241 GND.n2326 GND.n1240 9.3005
R15242 GND.n4613 GND.n1245 9.3005
R15243 GND.n4612 GND.n1246 9.3005
R15244 GND.n4611 GND.n1247 9.3005
R15245 GND.n2300 GND.n1248 9.3005
R15246 GND.n4607 GND.n1253 9.3005
R15247 GND.n4606 GND.n1254 9.3005
R15248 GND.n4605 GND.n1255 9.3005
R15249 GND.n2953 GND.n1256 9.3005
R15250 GND.n2952 GND.n1259 9.3005
R15251 GND.n4679 GND.n1157 9.3005
R15252 GND.n4678 GND.n1156 9.3005
R15253 GND.n4677 GND.n4676 9.3005
R15254 GND.n4675 GND.n1160 9.3005
R15255 GND.n4674 GND.n4673 9.3005
R15256 GND.n4672 GND.n1164 9.3005
R15257 GND.n4671 GND.n4670 9.3005
R15258 GND.n4669 GND.n1168 9.3005
R15259 GND.n4668 GND.n4667 9.3005
R15260 GND.n4666 GND.n1172 9.3005
R15261 GND.n4665 GND.n4664 9.3005
R15262 GND.n4663 GND.n1176 9.3005
R15263 GND.n4662 GND.n4661 9.3005
R15264 GND.n4660 GND.n1180 9.3005
R15265 GND.n4659 GND.n4658 9.3005
R15266 GND.n4657 GND.n1184 9.3005
R15267 GND.n4656 GND.n4655 9.3005
R15268 GND.n4654 GND.n1188 9.3005
R15269 GND.n4653 GND.n4652 9.3005
R15270 GND.n4651 GND.n1192 9.3005
R15271 GND.n4650 GND.n4649 9.3005
R15272 GND.n4648 GND.n1196 9.3005
R15273 GND.n4647 GND.n4646 9.3005
R15274 GND.n4645 GND.n1200 9.3005
R15275 GND.n4644 GND.n4643 9.3005
R15276 GND.n4642 GND.n1204 9.3005
R15277 GND.n4641 GND.n4640 9.3005
R15278 GND.n4639 GND.n1208 9.3005
R15279 GND.n4638 GND.n4637 9.3005
R15280 GND.n4636 GND.n1212 9.3005
R15281 GND.n4635 GND.n4634 9.3005
R15282 GND.n4633 GND.n1216 9.3005
R15283 GND.n4632 GND.n4631 9.3005
R15284 GND.n4630 GND.n1220 9.3005
R15285 GND.n4629 GND.n4628 9.3005
R15286 GND.n4627 GND.n1224 9.3005
R15287 GND.n4626 GND.n4625 9.3005
R15288 GND.n4624 GND.n1228 9.3005
R15289 GND.n4623 GND.n4622 9.3005
R15290 GND.n4621 GND.n1232 9.3005
R15291 GND.n4620 GND.n4619 9.3005
R15292 GND.n4618 GND.n1236 9.3005
R15293 GND.n4617 GND.n4616 9.3005
R15294 GND.n4615 GND.n1240 9.3005
R15295 GND.n4614 GND.n4613 9.3005
R15296 GND.n4612 GND.n1244 9.3005
R15297 GND.n4611 GND.n4610 9.3005
R15298 GND.n4609 GND.n1248 9.3005
R15299 GND.n4608 GND.n4607 9.3005
R15300 GND.n4606 GND.n1252 9.3005
R15301 GND.n4605 GND.n4604 9.3005
R15302 GND.n4603 GND.n1256 9.3005
R15303 GND.n4602 GND.n1259 9.3005
R15304 GND.n4680 GND.n4679 9.3005
R15305 GND.n2591 GND.n2575 9.3005
R15306 GND.n2593 GND.n2592 9.3005
R15307 GND.n2594 GND.n2570 9.3005
R15308 GND.n2596 GND.n2595 9.3005
R15309 GND.n2597 GND.n2569 9.3005
R15310 GND.n2599 GND.n2598 9.3005
R15311 GND.n2600 GND.n2564 9.3005
R15312 GND.n2602 GND.n2601 9.3005
R15313 GND.n2603 GND.n2563 9.3005
R15314 GND.n2605 GND.n2604 9.3005
R15315 GND.n2606 GND.n2558 9.3005
R15316 GND.n2608 GND.n2607 9.3005
R15317 GND.n2609 GND.n2557 9.3005
R15318 GND.n2611 GND.n2610 9.3005
R15319 GND.n2612 GND.n2554 9.3005
R15320 GND.n2590 GND.n2589 9.3005
R15321 GND.n2585 GND.n2584 9.3005
R15322 GND.n2581 GND.n2576 9.3005
R15323 GND.n2580 GND.n2579 9.3005
R15324 GND.n2502 GND.n2501 9.3005
R15325 GND.n2632 GND.n2631 9.3005
R15326 GND.n2633 GND.n2499 9.3005
R15327 GND.n2636 GND.n2635 9.3005
R15328 GND.n2634 GND.n2500 9.3005
R15329 GND.n2479 GND.n2478 9.3005
R15330 GND.n2657 GND.n2656 9.3005
R15331 GND.n2658 GND.n2476 9.3005
R15332 GND.n2661 GND.n2660 9.3005
R15333 GND.n2659 GND.n2477 9.3005
R15334 GND.n2457 GND.n2456 9.3005
R15335 GND.n2682 GND.n2681 9.3005
R15336 GND.n2683 GND.n2454 9.3005
R15337 GND.n2700 GND.n2699 9.3005
R15338 GND.n2698 GND.n2455 9.3005
R15339 GND.n2697 GND.n2696 9.3005
R15340 GND.n2695 GND.n2684 9.3005
R15341 GND.n2694 GND.n2693 9.3005
R15342 GND.n2692 GND.n2424 9.3005
R15343 GND.n2731 GND.n2423 9.3005
R15344 GND.n2733 GND.n2732 9.3005
R15345 GND.n2734 GND.n2422 9.3005
R15346 GND.n2736 GND.n2735 9.3005
R15347 GND.n2583 GND.n2582 9.3005
R15348 GND.n2739 GND.n2421 9.3005
R15349 GND.t32 GND.n2417 9.17771
R15350 GND.n2008 GND.t160 9.17771
R15351 GND.n96 GND.n71 8.92171
R15352 GND.n133 GND.n108 8.92171
R15353 GND.n165 GND.n140 8.92171
R15354 GND.n202 GND.n177 8.92171
R15355 GND.n27 GND.n2 8.92171
R15356 GND.n64 GND.n39 8.92171
R15357 GND.n281 GND.n256 8.92171
R15358 GND.n244 GND.n219 8.92171
R15359 GND.n350 GND.n325 8.92171
R15360 GND.n313 GND.n288 8.92171
R15361 GND.n420 GND.n395 8.92171
R15362 GND.n383 GND.n358 8.92171
R15363 GND.n4402 GND.n1510 8.86126
R15364 GND.n3320 GND.n2216 8.86126
R15365 GND.n3394 GND.n3393 8.86126
R15366 GND.n3422 GND.n1651 8.86126
R15367 GND.n3512 GND.n3494 8.72777
R15368 GND.n2766 GND.t38 8.5448
R15369 GND.n3875 GND.t57 8.5448
R15370 GND.n5675 GND.n5674 8.53706
R15371 GND.n2421 GND.n209 8.53706
R15372 GND.n4409 GND.n1502 8.22835
R15373 GND.n2210 GND.n2209 8.22835
R15374 GND.n3386 GND.n3385 8.22835
R15375 GND.n3440 GND.n2186 8.22835
R15376 GND.n97 GND.n69 8.14595
R15377 GND.n134 GND.n106 8.14595
R15378 GND.n166 GND.n138 8.14595
R15379 GND.n203 GND.n175 8.14595
R15380 GND.n28 GND.n0 8.14595
R15381 GND.n65 GND.n37 8.14595
R15382 GND.n282 GND.n254 8.14595
R15383 GND.n245 GND.n217 8.14595
R15384 GND.n351 GND.n323 8.14595
R15385 GND.n314 GND.n286 8.14595
R15386 GND.n421 GND.n393 8.14595
R15387 GND.n384 GND.n356 8.14595
R15388 GND.n3350 GND.t11 7.91189
R15389 GND.n2204 GND.t34 7.91189
R15390 GND.n5632 GND.n465 7.75808
R15391 GND.n4505 GND.n4504 7.75808
R15392 GND.n2589 GND.n2585 7.75808
R15393 GND.n4217 GND.n1812 7.75808
R15394 GND.n3149 GND.t87 7.59544
R15395 GND.t87 GND.n1492 7.59544
R15396 GND.t90 GND.n4415 7.59544
R15397 GND.n3272 GND.n1502 7.59544
R15398 GND.t6 GND.n1530 7.59544
R15399 GND.n3349 GND.n2210 7.59544
R15400 GND.n3386 GND.n2203 7.59544
R15401 GND.t60 GND.n1620 7.59544
R15402 GND.n3441 GND.n3440 7.59544
R15403 GND.n209 GND.n208 7.3623
R15404 GND.n5675 GND.n425 7.3623
R15405 GND.n2262 GND.n2261 7.30353
R15406 GND.n3511 GND.n3510 7.30353
R15407 GND.n4402 GND.n4401 6.96253
R15408 GND.n3303 GND.n2216 6.96253
R15409 GND.n3393 GND.n2200 6.96253
R15410 GND.n3422 GND.n1645 6.96253
R15411 GND.t72 GND.n2180 6.96253
R15412 GND.n4304 GND.t142 6.96253
R15413 GND.n207 GND.n137 6.61257
R15414 GND.n355 GND.n285 6.61257
R15415 GND.n3748 GND.n3747 6.5566
R15416 GND.n3079 GND.n3078 6.5566
R15417 GND.n3168 GND.n3163 6.5566
R15418 GND.n3573 GND.n3572 6.5566
R15419 GND.n2241 GND.n1474 6.32961
R15420 GND.n4416 GND.n1492 6.32961
R15421 GND.n3354 GND.n1559 6.32961
R15422 GND.n3366 GND.n1577 6.32961
R15423 GND.n3450 GND.n2181 6.32961
R15424 GND.n5604 GND.n5603 6.20656
R15425 GND.n4720 GND.n4719 6.20656
R15426 GND.t11 GND.n3349 6.01316
R15427 GND.t34 GND.n2203 6.01316
R15428 GND.n99 GND.n69 5.81868
R15429 GND.n136 GND.n106 5.81868
R15430 GND.n168 GND.n138 5.81868
R15431 GND.n205 GND.n175 5.81868
R15432 GND.n30 GND.n0 5.81868
R15433 GND.n67 GND.n37 5.81868
R15434 GND.n284 GND.n254 5.81868
R15435 GND.n247 GND.n217 5.81868
R15436 GND.n353 GND.n323 5.81868
R15437 GND.n316 GND.n286 5.81868
R15438 GND.n423 GND.n393 5.81868
R15439 GND.n386 GND.n356 5.81868
R15440 GND.n4395 GND.n1520 5.6967
R15441 GND.n3299 GND.n1523 5.6967
R15442 GND.n3372 GND.n1626 5.6967
R15443 GND.n2192 GND.n1629 5.6967
R15444 GND.n3752 GND.n3688 5.62001
R15445 GND.n3074 GND.n1290 5.62001
R15446 GND.n3164 GND.n1290 5.62001
R15447 GND.n3688 GND.n3577 5.62001
R15448 GND.n3821 GND.n3820 5.4308
R15449 GND.n2990 GND.n2276 5.4308
R15450 GND.n1458 GND.t14 5.38025
R15451 GND.n4284 GND.t22 5.38025
R15452 GND.n3360 GND.n1561 5.06379
R15453 GND.n3362 GND.n1575 5.06379
R15454 GND.n3780 GND.n3779 5.06379
R15455 GND.n3773 GND.t94 5.06379
R15456 GND.n97 GND.n96 5.04292
R15457 GND.n134 GND.n133 5.04292
R15458 GND.n166 GND.n165 5.04292
R15459 GND.n203 GND.n202 5.04292
R15460 GND.n28 GND.n27 5.04292
R15461 GND.n65 GND.n64 5.04292
R15462 GND.n282 GND.n281 5.04292
R15463 GND.n245 GND.n244 5.04292
R15464 GND.n351 GND.n350 5.04292
R15465 GND.n314 GND.n313 5.04292
R15466 GND.n421 GND.n420 5.04292
R15467 GND.n384 GND.n383 5.04292
R15468 GND.n208 GND.n68 4.7699
R15469 GND.n425 GND.n424 4.7699
R15470 GND.n4064 GND.n4063 4.74817
R15471 GND.n4017 GND.n1998 4.74817
R15472 GND.n4045 GND.n1997 4.74817
R15473 GND.n4023 GND.n1996 4.74817
R15474 GND.n4030 GND.n1995 4.74817
R15475 GND.n4064 GND.n1999 4.74817
R15476 GND.n4062 GND.n1998 4.74817
R15477 GND.n4018 GND.n1997 4.74817
R15478 GND.n4046 GND.n1996 4.74817
R15479 GND.n4022 GND.n1995 4.74817
R15480 GND.n2726 GND.n2725 4.74817
R15481 GND.n2819 GND.n2399 4.74817
R15482 GND.n2817 GND.n2816 4.74817
R15483 GND.n2750 GND.n2749 4.74817
R15484 GND.n2801 GND.n2800 4.74817
R15485 GND.n4006 GND.n2014 4.74817
R15486 GND.n4054 GND.n4008 4.74817
R15487 GND.n4052 GND.n4051 4.74817
R15488 GND.n4035 GND.n4034 4.74817
R15489 GND.n4036 GND.n1985 4.74817
R15490 GND.n2016 GND.n2014 4.74817
R15491 GND.n4008 GND.n4007 4.74817
R15492 GND.n4053 GND.n4052 4.74817
R15493 GND.n4034 GND.n4009 4.74817
R15494 GND.n4037 GND.n4036 4.74817
R15495 GND.n2830 GND.n2829 4.74817
R15496 GND.n2409 GND.n2385 4.74817
R15497 GND.n2810 GND.n2384 4.74817
R15498 GND.n2415 GND.n2383 4.74817
R15499 GND.n2382 GND.n2379 4.74817
R15500 GND.n2830 GND.n2386 4.74817
R15501 GND.n2828 GND.n2385 4.74817
R15502 GND.n2410 GND.n2384 4.74817
R15503 GND.n2811 GND.n2383 4.74817
R15504 GND.n2414 GND.n2382 4.74817
R15505 GND.n2725 GND.n2724 4.74817
R15506 GND.n2723 GND.n2399 4.74817
R15507 GND.n2818 GND.n2817 4.74817
R15508 GND.n2749 GND.n2400 4.74817
R15509 GND.n2802 GND.n2801 4.74817
R15510 GND.t103 GND.n2504 4.74734
R15511 GND.n3755 GND.t113 4.74734
R15512 GND.n5513 GND.t79 4.74734
R15513 GND.n207 GND.n206 4.7074
R15514 GND.n355 GND.n354 4.7074
R15515 GND.n3685 GND.n3624 4.6132
R15516 GND.n4575 GND.n1288 4.6132
R15517 GND.n3507 GND.n3494 4.46111
R15518 GND.n4388 GND.n4387 4.43088
R15519 GND.n4339 GND.n4338 4.43088
R15520 GND.n82 GND.n78 4.38594
R15521 GND.n119 GND.n115 4.38594
R15522 GND.n151 GND.n147 4.38594
R15523 GND.n188 GND.n184 4.38594
R15524 GND.n13 GND.n9 4.38594
R15525 GND.n50 GND.n46 4.38594
R15526 GND.n267 GND.n263 4.38594
R15527 GND.n230 GND.n226 4.38594
R15528 GND.n336 GND.n332 4.38594
R15529 GND.n299 GND.n295 4.38594
R15530 GND.n406 GND.n402 4.38594
R15531 GND.n369 GND.n365 4.38594
R15532 GND.n93 GND.n71 4.26717
R15533 GND.n130 GND.n108 4.26717
R15534 GND.n162 GND.n140 4.26717
R15535 GND.n199 GND.n177 4.26717
R15536 GND.n24 GND.n2 4.26717
R15537 GND.n61 GND.n39 4.26717
R15538 GND.n278 GND.n256 4.26717
R15539 GND.n241 GND.n219 4.26717
R15540 GND.n347 GND.n325 4.26717
R15541 GND.n310 GND.n288 4.26717
R15542 GND.n417 GND.n395 4.26717
R15543 GND.n380 GND.n358 4.26717
R15544 GND.n216 GND.n212 4.14478
R15545 GND.n3747 GND.n3746 4.05904
R15546 GND.n3080 GND.n3079 4.05904
R15547 GND.n3171 GND.n3163 4.05904
R15548 GND.n3572 GND.n3571 4.05904
R15549 GND.n2232 GND.n1494 3.79797
R15550 GND.n4311 GND.n1664 3.79797
R15551 GND.n2177 GND.t142 3.79797
R15552 GND.n216 GND.n215 3.60163
R15553 GND.n92 GND.n73 3.49141
R15554 GND.n129 GND.n110 3.49141
R15555 GND.n161 GND.n142 3.49141
R15556 GND.n198 GND.n179 3.49141
R15557 GND.n23 GND.n4 3.49141
R15558 GND.n60 GND.n41 3.49141
R15559 GND.n277 GND.n258 3.49141
R15560 GND.n240 GND.n221 3.49141
R15561 GND.n346 GND.n327 3.49141
R15562 GND.n309 GND.n290 3.49141
R15563 GND.n416 GND.n397 3.49141
R15564 GND.n379 GND.n360 3.49141
R15565 GND.n2930 GND.t75 3.48151
R15566 GND.n4422 GND.t173 3.48151
R15567 GND.t16 GND.n4304 3.48151
R15568 GND.n3888 GND.t83 3.48151
R15569 GND.n100 GND.t50 3.3005
R15570 GND.n100 GND.t44 3.3005
R15571 GND.n102 GND.t166 3.3005
R15572 GND.n102 GND.t33 3.3005
R15573 GND.n104 GND.t167 3.3005
R15574 GND.n104 GND.t26 3.3005
R15575 GND.n169 GND.t179 3.3005
R15576 GND.n169 GND.t10 3.3005
R15577 GND.n171 GND.t62 3.3005
R15578 GND.n171 GND.t59 3.3005
R15579 GND.n173 GND.t172 3.3005
R15580 GND.n173 GND.t54 3.3005
R15581 GND.n31 GND.t43 3.3005
R15582 GND.n31 GND.t64 3.3005
R15583 GND.n33 GND.t178 3.3005
R15584 GND.n33 GND.t45 3.3005
R15585 GND.n35 GND.t41 3.3005
R15586 GND.n35 GND.t8 3.3005
R15587 GND.n252 GND.t66 3.3005
R15588 GND.n252 GND.t3 3.3005
R15589 GND.n250 GND.t169 3.3005
R15590 GND.n250 GND.t163 3.3005
R15591 GND.n248 GND.t65 3.3005
R15592 GND.n248 GND.t31 3.3005
R15593 GND.n321 GND.t29 3.3005
R15594 GND.n321 GND.t164 3.3005
R15595 GND.n319 GND.t161 3.3005
R15596 GND.n319 GND.t175 3.3005
R15597 GND.n317 GND.t51 3.3005
R15598 GND.n317 GND.t5 3.3005
R15599 GND.n391 GND.t30 3.3005
R15600 GND.n391 GND.t170 3.3005
R15601 GND.n389 GND.t176 3.3005
R15602 GND.n389 GND.t49 3.3005
R15603 GND.n387 GND.t47 3.3005
R15604 GND.n387 GND.t162 3.3005
R15605 GND.n3233 GND.t110 3.16506
R15606 GND.n3139 GND.n3138 3.16506
R15607 GND.n3256 GND.t21 3.16506
R15608 GND.n4326 GND.t63 3.16506
R15609 GND.n4319 GND.n4318 3.16506
R15610 GND.n89 GND.n88 2.71565
R15611 GND.n126 GND.n125 2.71565
R15612 GND.n158 GND.n157 2.71565
R15613 GND.n195 GND.n194 2.71565
R15614 GND.n20 GND.n19 2.71565
R15615 GND.n57 GND.n56 2.71565
R15616 GND.n274 GND.n273 2.71565
R15617 GND.n237 GND.n236 2.71565
R15618 GND.n343 GND.n342 2.71565
R15619 GND.n306 GND.n305 2.71565
R15620 GND.n413 GND.n412 2.71565
R15621 GND.n376 GND.n375 2.71565
R15622 GND.t119 GND.n2231 2.53215
R15623 GND.n4408 GND.n1504 2.53215
R15624 GND.t148 GND.n1504 2.53215
R15625 GND.n3299 GND.t6 2.53215
R15626 GND.n4381 GND.t13 2.53215
R15627 GND.n4380 GND.n1541 2.53215
R15628 GND.n4374 GND.t27 2.53215
R15629 GND.t52 GND.n4352 2.53215
R15630 GND.n4346 GND.n1603 2.53215
R15631 GND.n4345 GND.t20 2.53215
R15632 GND.n3372 GND.t60 2.53215
R15633 GND.n2187 GND.n1653 2.53215
R15634 GND.n208 GND.n207 2.4477
R15635 GND.n425 GND.n355 2.4477
R15636 GND.n4065 GND.n4064 2.27742
R15637 GND.n4065 GND.n1998 2.27742
R15638 GND.n4065 GND.n1997 2.27742
R15639 GND.n4065 GND.n1996 2.27742
R15640 GND.n4065 GND.n1995 2.27742
R15641 GND.n2014 GND.n1984 2.27742
R15642 GND.n4008 GND.n1984 2.27742
R15643 GND.n4052 GND.n1984 2.27742
R15644 GND.n4034 GND.n1984 2.27742
R15645 GND.n4036 GND.n1984 2.27742
R15646 GND.n2831 GND.n2830 2.27742
R15647 GND.n2831 GND.n2385 2.27742
R15648 GND.n2831 GND.n2384 2.27742
R15649 GND.n2831 GND.n2383 2.27742
R15650 GND.n2831 GND.n2382 2.27742
R15651 GND.n2725 GND.n2381 2.27742
R15652 GND.n2399 GND.n2381 2.27742
R15653 GND.n2817 GND.n2381 2.27742
R15654 GND.n2749 GND.n2381 2.27742
R15655 GND.n2801 GND.n2381 2.27742
R15656 GND.n3255 GND.t36 2.21569
R15657 GND.n3294 GND.t36 2.21569
R15658 GND.n3418 GND.t18 2.21569
R15659 GND.t18 GND.n3417 2.21569
R15660 GND.n85 GND.n75 1.93989
R15661 GND.n122 GND.n112 1.93989
R15662 GND.n154 GND.n144 1.93989
R15663 GND.n191 GND.n181 1.93989
R15664 GND.n16 GND.n6 1.93989
R15665 GND.n53 GND.n43 1.93989
R15666 GND.n270 GND.n260 1.93989
R15667 GND.n233 GND.n223 1.93989
R15668 GND.n339 GND.n329 1.93989
R15669 GND.n302 GND.n292 1.93989
R15670 GND.n409 GND.n399 1.93989
R15671 GND.n372 GND.n362 1.93989
R15672 GND.t97 GND.n4429 1.89923
R15673 GND.t110 GND.n1485 1.89923
R15674 GND.n4416 GND.t90 1.89923
R15675 GND.n2231 GND.n2230 1.89923
R15676 GND.n3350 GND.n1550 1.89923
R15677 GND.n2204 GND.n1586 1.89923
R15678 GND.n3441 GND.t116 1.89923
R15679 GND.n4312 GND.n1662 1.89923
R15680 GND.n2181 GND.t68 1.89923
R15681 GND.n3223 GND.n1472 1.58278
R15682 GND.n3247 GND.t173 1.58278
R15683 GND.n4305 GND.t16 1.58278
R15684 GND.n3756 GND.n3755 1.58278
R15685 GND.n2638 GND.n2492 1.26632
R15686 GND.n2644 GND.n2494 1.26632
R15687 GND.n2640 GND.n2481 1.26632
R15688 GND.n2654 GND.n2483 1.26632
R15689 GND.n2486 GND.n2474 1.26632
R15690 GND.n2663 GND.n2469 1.26632
R15691 GND.n2669 GND.n2471 1.26632
R15692 GND.n2666 GND.n2459 1.26632
R15693 GND.n2679 GND.n2460 1.26632
R15694 GND.n2463 GND.n2452 1.26632
R15695 GND.n2702 GND.n2446 1.26632
R15696 GND.n2706 GND.n2449 1.26632
R15697 GND.n2716 GND.n2435 1.26632
R15698 GND.n2690 GND.n2687 1.26632
R15699 GND.n2728 GND.n2427 1.26632
R15700 GND.n2729 GND.n2389 1.26632
R15701 GND.n2826 GND.n2391 1.26632
R15702 GND.n2822 GND.n2821 1.26632
R15703 GND.n2402 GND.n2396 1.26632
R15704 GND.n2814 GND.n2403 1.26632
R15705 GND.n2813 GND.n2405 1.26632
R15706 GND.n2808 GND.n2417 1.26632
R15707 GND.n2805 GND.n2804 1.26632
R15708 GND.n2746 GND.n2373 1.26632
R15709 GND.n2836 GND.n2374 1.26632
R15710 GND.n2796 GND.n2795 1.26632
R15711 GND.n2845 GND.n2362 1.26632
R15712 GND.n2851 GND.n2364 1.26632
R15713 GND.n2848 GND.n2353 1.26632
R15714 GND.n2861 GND.n2354 1.26632
R15715 GND.n2787 GND.n2786 1.26632
R15716 GND.n2870 GND.n2343 1.26632
R15717 GND.n2876 GND.n2345 1.26632
R15718 GND.n2872 GND.n2333 1.26632
R15719 GND.n2886 GND.n2335 1.26632
R15720 GND.n2766 GND.n2765 1.26632
R15721 GND.n2898 GND.n2322 1.26632
R15722 GND.n2902 GND.n2324 1.26632
R15723 GND.n2911 GND.n2316 1.26632
R15724 GND.n2910 GND.n2301 1.26632
R15725 GND.n2939 GND.n2296 1.26632
R15726 GND.n2942 GND.n2298 1.26632
R15727 GND.n2931 GND.n2930 1.26632
R15728 GND.n2950 GND.n2289 1.26632
R15729 GND.n2955 GND.n1261 1.26632
R15730 GND.n4600 GND.n1263 1.26632
R15731 GND.n3256 GND.n1512 1.26632
R15732 GND.n3304 GND.n1532 1.26632
R15733 GND.t27 GND.n4373 1.26632
R15734 GND.n4353 GND.t52 1.26632
R15735 GND.n3376 GND.n1618 1.26632
R15736 GND.n4326 GND.n4325 1.26632
R15737 GND.n4297 GND.t94 1.26632
R15738 GND.n2137 GND.n2136 1.26632
R15739 GND.n3844 GND.n3843 1.26632
R15740 GND.n3893 GND.n2112 1.26632
R15741 GND.n3890 GND.n3888 1.26632
R15742 GND.n3903 GND.n2102 1.26632
R15743 GND.n2106 GND.n2103 1.26632
R15744 GND.n3912 GND.n2095 1.26632
R15745 GND.n3917 GND.n2089 1.26632
R15746 GND.n3914 GND.n2092 1.26632
R15747 GND.n3927 GND.n2080 1.26632
R15748 GND.n3875 GND.n3874 1.26632
R15749 GND.n3936 GND.n2072 1.26632
R15750 GND.n3942 GND.n2068 1.26632
R15751 GND.n3939 GND.n2070 1.26632
R15752 GND.n3952 GND.n2058 1.26632
R15753 GND.n2059 GND.n2051 1.26632
R15754 GND.n3964 GND.n3963 1.26632
R15755 GND.n3982 GND.n2036 1.26632
R15756 GND.n3978 GND.n2038 1.26632
R15757 GND.n3977 GND.n2043 1.26632
R15758 GND.n3991 GND.n2024 1.26632
R15759 GND.n2025 GND.n2017 1.26632
R15760 GND.n4003 GND.n4002 1.26632
R15761 GND.n4060 GND.n2002 1.26632
R15762 GND.n4057 GND.n2008 1.26632
R15763 GND.n4056 GND.n2011 1.26632
R15764 GND.n4012 GND.n4011 1.26632
R15765 GND.n4049 GND.n4048 1.26632
R15766 GND.n4043 GND.n4014 1.26632
R15767 GND.n4040 GND.n4027 1.26632
R15768 GND.n4039 GND.n4032 1.26632
R15769 GND.n4029 GND.n1988 1.26632
R15770 GND.n4072 GND.n4071 1.26632
R15771 GND.n4083 GND.n4082 1.26632
R15772 GND.n4087 GND.n1974 1.26632
R15773 GND.n1976 GND.n1963 1.26632
R15774 GND.n4098 GND.n4097 1.26632
R15775 GND.n1965 GND.n1956 1.26632
R15776 GND.n4117 GND.n4115 1.26632
R15777 GND.n4120 GND.n1951 1.26632
R15778 GND.n1954 GND.n1953 1.26632
R15779 GND.n4130 GND.n1943 1.26632
R15780 GND.n1944 GND.n594 1.26632
R15781 GND.n5487 GND.n5486 1.26632
R15782 GND.n5495 GND.n580 1.26632
R15783 GND.n583 GND.n572 1.26632
R15784 GND.n84 GND.n77 1.16414
R15785 GND.n121 GND.n114 1.16414
R15786 GND.n153 GND.n146 1.16414
R15787 GND.n190 GND.n183 1.16414
R15788 GND.n15 GND.n8 1.16414
R15789 GND.n52 GND.n45 1.16414
R15790 GND.n269 GND.n262 1.16414
R15791 GND.n232 GND.n225 1.16414
R15792 GND.n338 GND.n331 1.16414
R15793 GND.n301 GND.n294 1.16414
R15794 GND.n408 GND.n401 1.16414
R15795 GND.n371 GND.n364 1.16414
R15796 GND.n3822 GND.n3821 1.16414
R15797 GND.n2991 GND.n2990 1.16414
R15798 GND.n137 GND.n105 1.00481
R15799 GND.n105 GND.n103 1.00481
R15800 GND.n103 GND.n101 1.00481
R15801 GND.n206 GND.n174 1.00481
R15802 GND.n174 GND.n172 1.00481
R15803 GND.n172 GND.n170 1.00481
R15804 GND.n68 GND.n36 1.00481
R15805 GND.n36 GND.n34 1.00481
R15806 GND.n34 GND.n32 1.00481
R15807 GND.n251 GND.n249 1.00481
R15808 GND.n253 GND.n251 1.00481
R15809 GND.n285 GND.n253 1.00481
R15810 GND.n320 GND.n318 1.00481
R15811 GND.n322 GND.n320 1.00481
R15812 GND.n354 GND.n322 1.00481
R15813 GND.n390 GND.n388 1.00481
R15814 GND.n392 GND.n390 1.00481
R15815 GND.n424 GND.n392 1.00481
R15816 GND GND.n209 0.99596
R15817 GND.n4575 GND.n4574 0.970197
R15818 GND.n3685 GND.n3684 0.970197
R15819 GND.n211 GND.n210 0.962709
R15820 GND.n212 GND.n211 0.962709
R15821 GND.n214 GND.n213 0.962709
R15822 GND.n215 GND.n214 0.962709
R15823 GND.n2686 GND.t7 0.949867
R15824 GND.n1989 GND.t28 0.949867
R15825 GND.n3232 GND.n3231 0.633411
R15826 GND.n3149 GND.n2240 0.633411
R15827 GND.n3319 GND.t13 0.633411
R15828 GND.n4367 GND.n4366 0.633411
R15829 GND.n4360 GND.n4359 0.633411
R15830 GND.n2198 GND.t20 0.633411
R15831 GND.t68 GND.t72 0.633411
R15832 GND.n3451 GND.n1678 0.633411
R15833 GND.n4298 GND.n1686 0.633411
R15834 GND.n4065 GND.n1984 0.586625
R15835 GND.n2831 GND.n2381 0.586625
R15836 GND.n5676 GND.n5675 0.57484
R15837 GND.n3811 GND.n2162 0.48678
R15838 GND.n3002 GND.n3001 0.48678
R15839 GND.n5634 GND.n5633 0.483732
R15840 GND.n2584 GND.n2583 0.483732
R15841 GND.n3592 GND.n3587 0.471537
R15842 GND.n2548 GND.n1115 0.471537
R15843 GND.n5627 GND.n497 0.471537
R15844 GND.n4597 GND.n4596 0.471537
R15845 GND.n4886 GND.n4885 0.438
R15846 GND.n5316 GND.n699 0.438
R15847 GND.n5478 GND.n600 0.438
R15848 GND.n2539 GND.n2538 0.438
R15849 GND.n81 GND.n80 0.388379
R15850 GND.n118 GND.n117 0.388379
R15851 GND.n150 GND.n149 0.388379
R15852 GND.n187 GND.n186 0.388379
R15853 GND.n12 GND.n11 0.388379
R15854 GND.n49 GND.n48 0.388379
R15855 GND.n266 GND.n265 0.388379
R15856 GND.n229 GND.n228 0.388379
R15857 GND.n335 GND.n334 0.388379
R15858 GND.n298 GND.n297 0.388379
R15859 GND.n405 GND.n404 0.388379
R15860 GND.n368 GND.n367 0.388379
R15861 GND.n5605 GND.n5604 0.388379
R15862 GND.n4721 GND.n4720 0.388379
R15863 GND.n5676 GND.n216 0.37321
R15864 GND.n2715 GND.t7 0.316956
R15865 GND.n2845 GND.t42 0.316956
R15866 GND.t125 GND.n1412 0.316956
R15867 GND.n3804 GND.t132 0.316956
R15868 GND.n2043 GND.t4 0.316956
R15869 GND.t28 GND.n1980 0.316956
R15870 GND.n5566 GND.n550 0.293183
R15871 GND.n2554 GND.n1154 0.293183
R15872 GND.n4200 GND.n1854 0.280988
R15873 GND.n4684 GND.n1154 0.280988
R15874 GND.n5576 GND.n550 0.280988
R15875 GND.n4547 GND.n4545 0.280988
R15876 GND.n3838 GND.n3837 0.253549
R15877 GND.n2960 GND.n2959 0.253549
R15878 GND.n1406 GND.n1320 0.245927
R15879 GND.n4209 GND.n4207 0.245927
R15880 GND.n3624 GND.n3623 0.229039
R15881 GND.n3627 GND.n3624 0.229039
R15882 GND.n1288 GND.n1283 0.229039
R15883 GND.n4573 GND.n1288 0.229039
R15884 GND GND.n5676 0.213018
R15885 GND.n98 GND.n70 0.155672
R15886 GND.n91 GND.n70 0.155672
R15887 GND.n91 GND.n90 0.155672
R15888 GND.n90 GND.n74 0.155672
R15889 GND.n83 GND.n74 0.155672
R15890 GND.n83 GND.n82 0.155672
R15891 GND.n135 GND.n107 0.155672
R15892 GND.n128 GND.n107 0.155672
R15893 GND.n128 GND.n127 0.155672
R15894 GND.n127 GND.n111 0.155672
R15895 GND.n120 GND.n111 0.155672
R15896 GND.n120 GND.n119 0.155672
R15897 GND.n167 GND.n139 0.155672
R15898 GND.n160 GND.n139 0.155672
R15899 GND.n160 GND.n159 0.155672
R15900 GND.n159 GND.n143 0.155672
R15901 GND.n152 GND.n143 0.155672
R15902 GND.n152 GND.n151 0.155672
R15903 GND.n204 GND.n176 0.155672
R15904 GND.n197 GND.n176 0.155672
R15905 GND.n197 GND.n196 0.155672
R15906 GND.n196 GND.n180 0.155672
R15907 GND.n189 GND.n180 0.155672
R15908 GND.n189 GND.n188 0.155672
R15909 GND.n29 GND.n1 0.155672
R15910 GND.n22 GND.n1 0.155672
R15911 GND.n22 GND.n21 0.155672
R15912 GND.n21 GND.n5 0.155672
R15913 GND.n14 GND.n5 0.155672
R15914 GND.n14 GND.n13 0.155672
R15915 GND.n66 GND.n38 0.155672
R15916 GND.n59 GND.n38 0.155672
R15917 GND.n59 GND.n58 0.155672
R15918 GND.n58 GND.n42 0.155672
R15919 GND.n51 GND.n42 0.155672
R15920 GND.n51 GND.n50 0.155672
R15921 GND.n283 GND.n255 0.155672
R15922 GND.n276 GND.n255 0.155672
R15923 GND.n276 GND.n275 0.155672
R15924 GND.n275 GND.n259 0.155672
R15925 GND.n268 GND.n259 0.155672
R15926 GND.n268 GND.n267 0.155672
R15927 GND.n246 GND.n218 0.155672
R15928 GND.n239 GND.n218 0.155672
R15929 GND.n239 GND.n238 0.155672
R15930 GND.n238 GND.n222 0.155672
R15931 GND.n231 GND.n222 0.155672
R15932 GND.n231 GND.n230 0.155672
R15933 GND.n352 GND.n324 0.155672
R15934 GND.n345 GND.n324 0.155672
R15935 GND.n345 GND.n344 0.155672
R15936 GND.n344 GND.n328 0.155672
R15937 GND.n337 GND.n328 0.155672
R15938 GND.n337 GND.n336 0.155672
R15939 GND.n315 GND.n287 0.155672
R15940 GND.n308 GND.n287 0.155672
R15941 GND.n308 GND.n307 0.155672
R15942 GND.n307 GND.n291 0.155672
R15943 GND.n300 GND.n291 0.155672
R15944 GND.n300 GND.n299 0.155672
R15945 GND.n422 GND.n394 0.155672
R15946 GND.n415 GND.n394 0.155672
R15947 GND.n415 GND.n414 0.155672
R15948 GND.n414 GND.n398 0.155672
R15949 GND.n407 GND.n398 0.155672
R15950 GND.n407 GND.n406 0.155672
R15951 GND.n385 GND.n357 0.155672
R15952 GND.n378 GND.n357 0.155672
R15953 GND.n378 GND.n377 0.155672
R15954 GND.n377 GND.n361 0.155672
R15955 GND.n370 GND.n361 0.155672
R15956 GND.n370 GND.n369 0.155672
R15957 GND.n1407 GND.n1406 0.152939
R15958 GND.n1408 GND.n1407 0.152939
R15959 GND.n1409 GND.n1408 0.152939
R15960 GND.n1438 GND.n1409 0.152939
R15961 GND.n1439 GND.n1438 0.152939
R15962 GND.n1440 GND.n1439 0.152939
R15963 GND.n1441 GND.n1440 0.152939
R15964 GND.n1442 GND.n1441 0.152939
R15965 GND.n1465 GND.n1442 0.152939
R15966 GND.n1466 GND.n1465 0.152939
R15967 GND.n1467 GND.n1466 0.152939
R15968 GND.n1468 GND.n1467 0.152939
R15969 GND.n1469 GND.n1468 0.152939
R15970 GND.n3237 GND.n1469 0.152939
R15971 GND.n3238 GND.n3237 0.152939
R15972 GND.n3239 GND.n3238 0.152939
R15973 GND.n3240 GND.n3239 0.152939
R15974 GND.n3242 GND.n3240 0.152939
R15975 GND.n3242 GND.n3241 0.152939
R15976 GND.n3241 GND.n2224 0.152939
R15977 GND.n3277 GND.n2224 0.152939
R15978 GND.n3278 GND.n3277 0.152939
R15979 GND.n3279 GND.n3278 0.152939
R15980 GND.n3280 GND.n3279 0.152939
R15981 GND.n3281 GND.n3280 0.152939
R15982 GND.n3283 GND.n3281 0.152939
R15983 GND.n3283 GND.n3282 0.152939
R15984 GND.n3282 GND.n1545 0.152939
R15985 GND.n1546 GND.n1545 0.152939
R15986 GND.n1547 GND.n1546 0.152939
R15987 GND.n1590 GND.n1547 0.152939
R15988 GND.n1591 GND.n1590 0.152939
R15989 GND.n1596 GND.n1591 0.152939
R15990 GND.n1597 GND.n1596 0.152939
R15991 GND.n1598 GND.n1597 0.152939
R15992 GND.n1599 GND.n1598 0.152939
R15993 GND.n1600 GND.n1599 0.152939
R15994 GND.n1633 GND.n1600 0.152939
R15995 GND.n1636 GND.n1633 0.152939
R15996 GND.n1637 GND.n1636 0.152939
R15997 GND.n1638 GND.n1637 0.152939
R15998 GND.n1639 GND.n1638 0.152939
R15999 GND.n1640 GND.n1639 0.152939
R16000 GND.n1668 GND.n1640 0.152939
R16001 GND.n1671 GND.n1668 0.152939
R16002 GND.n1672 GND.n1671 0.152939
R16003 GND.n1673 GND.n1672 0.152939
R16004 GND.n1674 GND.n1673 0.152939
R16005 GND.n1675 GND.n1674 0.152939
R16006 GND.n1690 GND.n1675 0.152939
R16007 GND.n1691 GND.n1690 0.152939
R16008 GND.n1692 GND.n1691 0.152939
R16009 GND.n1693 GND.n1692 0.152939
R16010 GND.n1713 GND.n1693 0.152939
R16011 GND.n1714 GND.n1713 0.152939
R16012 GND.n1715 GND.n1714 0.152939
R16013 GND.n1716 GND.n1715 0.152939
R16014 GND.n1717 GND.n1716 0.152939
R16015 GND.n1740 GND.n1717 0.152939
R16016 GND.n1741 GND.n1740 0.152939
R16017 GND.n1742 GND.n1741 0.152939
R16018 GND.n1743 GND.n1742 0.152939
R16019 GND.n1744 GND.n1743 0.152939
R16020 GND.n4205 GND.n1744 0.152939
R16021 GND.n4207 GND.n4205 0.152939
R16022 GND.n4887 GND.n4886 0.152939
R16023 GND.n4887 GND.n950 0.152939
R16024 GND.n4895 GND.n950 0.152939
R16025 GND.n4896 GND.n4895 0.152939
R16026 GND.n4897 GND.n4896 0.152939
R16027 GND.n4897 GND.n944 0.152939
R16028 GND.n4905 GND.n944 0.152939
R16029 GND.n4906 GND.n4905 0.152939
R16030 GND.n4907 GND.n4906 0.152939
R16031 GND.n4907 GND.n938 0.152939
R16032 GND.n4915 GND.n938 0.152939
R16033 GND.n4916 GND.n4915 0.152939
R16034 GND.n4917 GND.n4916 0.152939
R16035 GND.n4917 GND.n932 0.152939
R16036 GND.n4925 GND.n932 0.152939
R16037 GND.n4926 GND.n4925 0.152939
R16038 GND.n4927 GND.n4926 0.152939
R16039 GND.n4927 GND.n926 0.152939
R16040 GND.n4935 GND.n926 0.152939
R16041 GND.n4936 GND.n4935 0.152939
R16042 GND.n4937 GND.n4936 0.152939
R16043 GND.n4937 GND.n920 0.152939
R16044 GND.n4945 GND.n920 0.152939
R16045 GND.n4946 GND.n4945 0.152939
R16046 GND.n4947 GND.n4946 0.152939
R16047 GND.n4947 GND.n914 0.152939
R16048 GND.n4955 GND.n914 0.152939
R16049 GND.n4956 GND.n4955 0.152939
R16050 GND.n4957 GND.n4956 0.152939
R16051 GND.n4957 GND.n908 0.152939
R16052 GND.n4965 GND.n908 0.152939
R16053 GND.n4966 GND.n4965 0.152939
R16054 GND.n4967 GND.n4966 0.152939
R16055 GND.n4967 GND.n902 0.152939
R16056 GND.n4975 GND.n902 0.152939
R16057 GND.n4976 GND.n4975 0.152939
R16058 GND.n4977 GND.n4976 0.152939
R16059 GND.n4977 GND.n896 0.152939
R16060 GND.n4985 GND.n896 0.152939
R16061 GND.n4986 GND.n4985 0.152939
R16062 GND.n4987 GND.n4986 0.152939
R16063 GND.n4987 GND.n890 0.152939
R16064 GND.n4995 GND.n890 0.152939
R16065 GND.n4996 GND.n4995 0.152939
R16066 GND.n4997 GND.n4996 0.152939
R16067 GND.n4997 GND.n884 0.152939
R16068 GND.n5005 GND.n884 0.152939
R16069 GND.n5006 GND.n5005 0.152939
R16070 GND.n5007 GND.n5006 0.152939
R16071 GND.n5007 GND.n878 0.152939
R16072 GND.n5015 GND.n878 0.152939
R16073 GND.n5016 GND.n5015 0.152939
R16074 GND.n5017 GND.n5016 0.152939
R16075 GND.n5017 GND.n872 0.152939
R16076 GND.n5025 GND.n872 0.152939
R16077 GND.n5026 GND.n5025 0.152939
R16078 GND.n5027 GND.n5026 0.152939
R16079 GND.n5027 GND.n866 0.152939
R16080 GND.n5035 GND.n866 0.152939
R16081 GND.n5036 GND.n5035 0.152939
R16082 GND.n5037 GND.n5036 0.152939
R16083 GND.n5037 GND.n860 0.152939
R16084 GND.n5045 GND.n860 0.152939
R16085 GND.n5046 GND.n5045 0.152939
R16086 GND.n5047 GND.n5046 0.152939
R16087 GND.n5047 GND.n854 0.152939
R16088 GND.n5055 GND.n854 0.152939
R16089 GND.n5056 GND.n5055 0.152939
R16090 GND.n5057 GND.n5056 0.152939
R16091 GND.n5057 GND.n848 0.152939
R16092 GND.n5065 GND.n848 0.152939
R16093 GND.n5066 GND.n5065 0.152939
R16094 GND.n5067 GND.n5066 0.152939
R16095 GND.n5067 GND.n842 0.152939
R16096 GND.n5075 GND.n842 0.152939
R16097 GND.n5076 GND.n5075 0.152939
R16098 GND.n5077 GND.n5076 0.152939
R16099 GND.n5077 GND.n836 0.152939
R16100 GND.n5085 GND.n836 0.152939
R16101 GND.n5086 GND.n5085 0.152939
R16102 GND.n5087 GND.n5086 0.152939
R16103 GND.n5087 GND.n830 0.152939
R16104 GND.n5095 GND.n830 0.152939
R16105 GND.n5096 GND.n5095 0.152939
R16106 GND.n5097 GND.n5096 0.152939
R16107 GND.n5097 GND.n824 0.152939
R16108 GND.n5105 GND.n824 0.152939
R16109 GND.n5106 GND.n5105 0.152939
R16110 GND.n5107 GND.n5106 0.152939
R16111 GND.n5107 GND.n818 0.152939
R16112 GND.n5115 GND.n818 0.152939
R16113 GND.n5116 GND.n5115 0.152939
R16114 GND.n5117 GND.n5116 0.152939
R16115 GND.n5117 GND.n812 0.152939
R16116 GND.n5125 GND.n812 0.152939
R16117 GND.n5126 GND.n5125 0.152939
R16118 GND.n5127 GND.n5126 0.152939
R16119 GND.n5127 GND.n806 0.152939
R16120 GND.n5135 GND.n806 0.152939
R16121 GND.n5136 GND.n5135 0.152939
R16122 GND.n5137 GND.n5136 0.152939
R16123 GND.n5137 GND.n800 0.152939
R16124 GND.n5145 GND.n800 0.152939
R16125 GND.n5146 GND.n5145 0.152939
R16126 GND.n5147 GND.n5146 0.152939
R16127 GND.n5147 GND.n794 0.152939
R16128 GND.n5155 GND.n794 0.152939
R16129 GND.n5156 GND.n5155 0.152939
R16130 GND.n5157 GND.n5156 0.152939
R16131 GND.n5157 GND.n788 0.152939
R16132 GND.n5165 GND.n788 0.152939
R16133 GND.n5166 GND.n5165 0.152939
R16134 GND.n5167 GND.n5166 0.152939
R16135 GND.n5167 GND.n782 0.152939
R16136 GND.n5175 GND.n782 0.152939
R16137 GND.n5176 GND.n5175 0.152939
R16138 GND.n5177 GND.n5176 0.152939
R16139 GND.n5177 GND.n776 0.152939
R16140 GND.n5185 GND.n776 0.152939
R16141 GND.n5186 GND.n5185 0.152939
R16142 GND.n5187 GND.n5186 0.152939
R16143 GND.n5187 GND.n770 0.152939
R16144 GND.n5195 GND.n770 0.152939
R16145 GND.n5196 GND.n5195 0.152939
R16146 GND.n5197 GND.n5196 0.152939
R16147 GND.n5197 GND.n764 0.152939
R16148 GND.n5205 GND.n764 0.152939
R16149 GND.n5206 GND.n5205 0.152939
R16150 GND.n5207 GND.n5206 0.152939
R16151 GND.n5207 GND.n758 0.152939
R16152 GND.n5215 GND.n758 0.152939
R16153 GND.n5216 GND.n5215 0.152939
R16154 GND.n5217 GND.n5216 0.152939
R16155 GND.n5217 GND.n752 0.152939
R16156 GND.n5225 GND.n752 0.152939
R16157 GND.n5226 GND.n5225 0.152939
R16158 GND.n5227 GND.n5226 0.152939
R16159 GND.n5227 GND.n746 0.152939
R16160 GND.n5235 GND.n746 0.152939
R16161 GND.n5236 GND.n5235 0.152939
R16162 GND.n5237 GND.n5236 0.152939
R16163 GND.n5237 GND.n740 0.152939
R16164 GND.n5245 GND.n740 0.152939
R16165 GND.n5246 GND.n5245 0.152939
R16166 GND.n5247 GND.n5246 0.152939
R16167 GND.n5247 GND.n734 0.152939
R16168 GND.n5255 GND.n734 0.152939
R16169 GND.n5256 GND.n5255 0.152939
R16170 GND.n5257 GND.n5256 0.152939
R16171 GND.n5257 GND.n728 0.152939
R16172 GND.n5265 GND.n728 0.152939
R16173 GND.n5266 GND.n5265 0.152939
R16174 GND.n5267 GND.n5266 0.152939
R16175 GND.n5267 GND.n722 0.152939
R16176 GND.n5275 GND.n722 0.152939
R16177 GND.n5276 GND.n5275 0.152939
R16178 GND.n5277 GND.n5276 0.152939
R16179 GND.n5277 GND.n716 0.152939
R16180 GND.n5285 GND.n716 0.152939
R16181 GND.n5286 GND.n5285 0.152939
R16182 GND.n5287 GND.n5286 0.152939
R16183 GND.n5287 GND.n710 0.152939
R16184 GND.n5295 GND.n710 0.152939
R16185 GND.n5296 GND.n5295 0.152939
R16186 GND.n5297 GND.n5296 0.152939
R16187 GND.n5297 GND.n704 0.152939
R16188 GND.n5305 GND.n704 0.152939
R16189 GND.n5306 GND.n5305 0.152939
R16190 GND.n5307 GND.n5306 0.152939
R16191 GND.n5307 GND.n699 0.152939
R16192 GND.n5317 GND.n5316 0.152939
R16193 GND.n5318 GND.n5317 0.152939
R16194 GND.n5318 GND.n693 0.152939
R16195 GND.n5326 GND.n693 0.152939
R16196 GND.n5327 GND.n5326 0.152939
R16197 GND.n5328 GND.n5327 0.152939
R16198 GND.n5328 GND.n687 0.152939
R16199 GND.n5336 GND.n687 0.152939
R16200 GND.n5337 GND.n5336 0.152939
R16201 GND.n5338 GND.n5337 0.152939
R16202 GND.n5338 GND.n681 0.152939
R16203 GND.n5346 GND.n681 0.152939
R16204 GND.n5347 GND.n5346 0.152939
R16205 GND.n5348 GND.n5347 0.152939
R16206 GND.n5348 GND.n675 0.152939
R16207 GND.n5356 GND.n675 0.152939
R16208 GND.n5357 GND.n5356 0.152939
R16209 GND.n5358 GND.n5357 0.152939
R16210 GND.n5358 GND.n669 0.152939
R16211 GND.n5366 GND.n669 0.152939
R16212 GND.n5367 GND.n5366 0.152939
R16213 GND.n5368 GND.n5367 0.152939
R16214 GND.n5368 GND.n663 0.152939
R16215 GND.n5376 GND.n663 0.152939
R16216 GND.n5377 GND.n5376 0.152939
R16217 GND.n5378 GND.n5377 0.152939
R16218 GND.n5378 GND.n657 0.152939
R16219 GND.n5386 GND.n657 0.152939
R16220 GND.n5387 GND.n5386 0.152939
R16221 GND.n5388 GND.n5387 0.152939
R16222 GND.n5388 GND.n651 0.152939
R16223 GND.n5396 GND.n651 0.152939
R16224 GND.n5397 GND.n5396 0.152939
R16225 GND.n5398 GND.n5397 0.152939
R16226 GND.n5398 GND.n645 0.152939
R16227 GND.n5406 GND.n645 0.152939
R16228 GND.n5407 GND.n5406 0.152939
R16229 GND.n5408 GND.n5407 0.152939
R16230 GND.n5408 GND.n639 0.152939
R16231 GND.n5416 GND.n639 0.152939
R16232 GND.n5417 GND.n5416 0.152939
R16233 GND.n5418 GND.n5417 0.152939
R16234 GND.n5418 GND.n633 0.152939
R16235 GND.n5426 GND.n633 0.152939
R16236 GND.n5427 GND.n5426 0.152939
R16237 GND.n5428 GND.n5427 0.152939
R16238 GND.n5428 GND.n627 0.152939
R16239 GND.n5436 GND.n627 0.152939
R16240 GND.n5437 GND.n5436 0.152939
R16241 GND.n5438 GND.n5437 0.152939
R16242 GND.n5438 GND.n621 0.152939
R16243 GND.n5446 GND.n621 0.152939
R16244 GND.n5447 GND.n5446 0.152939
R16245 GND.n5448 GND.n5447 0.152939
R16246 GND.n5448 GND.n615 0.152939
R16247 GND.n5456 GND.n615 0.152939
R16248 GND.n5457 GND.n5456 0.152939
R16249 GND.n5458 GND.n5457 0.152939
R16250 GND.n5458 GND.n609 0.152939
R16251 GND.n5466 GND.n609 0.152939
R16252 GND.n5467 GND.n5466 0.152939
R16253 GND.n5468 GND.n5467 0.152939
R16254 GND.n5468 GND.n603 0.152939
R16255 GND.n5476 GND.n603 0.152939
R16256 GND.n5477 GND.n5476 0.152939
R16257 GND.n5478 GND.n5477 0.152939
R16258 GND.n4076 GND.n4075 0.152939
R16259 GND.n4077 GND.n4076 0.152939
R16260 GND.n4078 GND.n4077 0.152939
R16261 GND.n4078 GND.n1960 0.152939
R16262 GND.n4101 GND.n1960 0.152939
R16263 GND.n4102 GND.n4101 0.152939
R16264 GND.n4103 GND.n4102 0.152939
R16265 GND.n4104 GND.n4103 0.152939
R16266 GND.n4105 GND.n4104 0.152939
R16267 GND.n4107 GND.n4105 0.152939
R16268 GND.n4107 GND.n4106 0.152939
R16269 GND.n4106 GND.n598 0.152939
R16270 GND.n599 GND.n598 0.152939
R16271 GND.n600 GND.n599 0.152939
R16272 GND.n4066 GND.n4065 0.152939
R16273 GND.n4067 GND.n4066 0.152939
R16274 GND.n4067 GND.n1971 0.152939
R16275 GND.n4090 GND.n1971 0.152939
R16276 GND.n4091 GND.n4090 0.152939
R16277 GND.n4092 GND.n4091 0.152939
R16278 GND.n4093 GND.n4092 0.152939
R16279 GND.n4093 GND.n1948 0.152939
R16280 GND.n4123 GND.n1948 0.152939
R16281 GND.n4124 GND.n4123 0.152939
R16282 GND.n4125 GND.n4124 0.152939
R16283 GND.n4126 GND.n4125 0.152939
R16284 GND.n4126 GND.n577 0.152939
R16285 GND.n5498 GND.n577 0.152939
R16286 GND.n5499 GND.n5498 0.152939
R16287 GND.n5500 GND.n5499 0.152939
R16288 GND.n5500 GND.n559 0.152939
R16289 GND.n5516 GND.n559 0.152939
R16290 GND.n5517 GND.n5516 0.152939
R16291 GND.n5518 GND.n5517 0.152939
R16292 GND.n5518 GND.n497 0.152939
R16293 GND.n3593 GND.n3592 0.152939
R16294 GND.n3594 GND.n3593 0.152939
R16295 GND.n3594 GND.n3585 0.152939
R16296 GND.n3602 GND.n3585 0.152939
R16297 GND.n3603 GND.n3602 0.152939
R16298 GND.n3604 GND.n3603 0.152939
R16299 GND.n3604 GND.n3583 0.152939
R16300 GND.n3612 GND.n3583 0.152939
R16301 GND.n3613 GND.n3612 0.152939
R16302 GND.n3614 GND.n3613 0.152939
R16303 GND.n3614 GND.n3581 0.152939
R16304 GND.n3622 GND.n3581 0.152939
R16305 GND.n3623 GND.n3622 0.152939
R16306 GND.n3628 GND.n3627 0.152939
R16307 GND.n3629 GND.n3628 0.152939
R16308 GND.n3630 GND.n3629 0.152939
R16309 GND.n3631 GND.n3630 0.152939
R16310 GND.n3632 GND.n3631 0.152939
R16311 GND.n3633 GND.n3632 0.152939
R16312 GND.n3634 GND.n3633 0.152939
R16313 GND.n3635 GND.n3634 0.152939
R16314 GND.n3636 GND.n3635 0.152939
R16315 GND.n3637 GND.n3636 0.152939
R16316 GND.n3638 GND.n3637 0.152939
R16317 GND.n3639 GND.n3638 0.152939
R16318 GND.n3640 GND.n3639 0.152939
R16319 GND.n3641 GND.n3640 0.152939
R16320 GND.n3642 GND.n3641 0.152939
R16321 GND.n3651 GND.n3642 0.152939
R16322 GND.n3651 GND.n3650 0.152939
R16323 GND.n3650 GND.n1854 0.152939
R16324 GND.n3587 GND.n2109 0.152939
R16325 GND.n3896 GND.n2109 0.152939
R16326 GND.n3897 GND.n3896 0.152939
R16327 GND.n3898 GND.n3897 0.152939
R16328 GND.n3899 GND.n3898 0.152939
R16329 GND.n3899 GND.n2086 0.152939
R16330 GND.n3920 GND.n2086 0.152939
R16331 GND.n3921 GND.n3920 0.152939
R16332 GND.n3922 GND.n3921 0.152939
R16333 GND.n3923 GND.n3922 0.152939
R16334 GND.n3923 GND.n2065 0.152939
R16335 GND.n3945 GND.n2065 0.152939
R16336 GND.n3946 GND.n3945 0.152939
R16337 GND.n3947 GND.n3946 0.152939
R16338 GND.n3948 GND.n3947 0.152939
R16339 GND.n3948 GND.n2032 0.152939
R16340 GND.n3985 GND.n2032 0.152939
R16341 GND.n3986 GND.n3985 0.152939
R16342 GND.n3987 GND.n3986 0.152939
R16343 GND.n3987 GND.n1994 0.152939
R16344 GND.n4065 GND.n1994 0.152939
R16345 GND.n2754 GND.n2751 0.152939
R16346 GND.n2755 GND.n2754 0.152939
R16347 GND.n2756 GND.n2755 0.152939
R16348 GND.n2757 GND.n2756 0.152939
R16349 GND.n2760 GND.n2757 0.152939
R16350 GND.n2761 GND.n2760 0.152939
R16351 GND.n2762 GND.n2761 0.152939
R16352 GND.n2763 GND.n2762 0.152939
R16353 GND.n2768 GND.n2763 0.152939
R16354 GND.n2769 GND.n2768 0.152939
R16355 GND.n2770 GND.n2769 0.152939
R16356 GND.n2771 GND.n2770 0.152939
R16357 GND.n2773 GND.n2771 0.152939
R16358 GND.n2773 GND.n2772 0.152939
R16359 GND.n2772 GND.n2311 0.152939
R16360 GND.n2916 GND.n2311 0.152939
R16361 GND.n2917 GND.n2916 0.152939
R16362 GND.n2918 GND.n2917 0.152939
R16363 GND.n2919 GND.n2918 0.152939
R16364 GND.n2920 GND.n2919 0.152939
R16365 GND.n2922 GND.n2920 0.152939
R16366 GND.n2922 GND.n2921 0.152939
R16367 GND.n2921 GND.n1395 0.152939
R16368 GND.n1396 GND.n1395 0.152939
R16369 GND.n1397 GND.n1396 0.152939
R16370 GND.n1418 GND.n1397 0.152939
R16371 GND.n1419 GND.n1418 0.152939
R16372 GND.n1420 GND.n1419 0.152939
R16373 GND.n1424 GND.n1420 0.152939
R16374 GND.n1425 GND.n1424 0.152939
R16375 GND.n1426 GND.n1425 0.152939
R16376 GND.n1427 GND.n1426 0.152939
R16377 GND.n1428 GND.n1427 0.152939
R16378 GND.n1451 GND.n1428 0.152939
R16379 GND.n1452 GND.n1451 0.152939
R16380 GND.n1453 GND.n1452 0.152939
R16381 GND.n1454 GND.n1453 0.152939
R16382 GND.n1455 GND.n1454 0.152939
R16383 GND.n1478 GND.n1455 0.152939
R16384 GND.n1479 GND.n1478 0.152939
R16385 GND.n1480 GND.n1479 0.152939
R16386 GND.n1481 GND.n1480 0.152939
R16387 GND.n1482 GND.n1481 0.152939
R16388 GND.n1496 GND.n1482 0.152939
R16389 GND.n1497 GND.n1496 0.152939
R16390 GND.n1498 GND.n1497 0.152939
R16391 GND.n1499 GND.n1498 0.152939
R16392 GND.n1514 GND.n1499 0.152939
R16393 GND.n1515 GND.n1514 0.152939
R16394 GND.n1516 GND.n1515 0.152939
R16395 GND.n1517 GND.n1516 0.152939
R16396 GND.n1534 GND.n1517 0.152939
R16397 GND.n1535 GND.n1534 0.152939
R16398 GND.n1536 GND.n1535 0.152939
R16399 GND.n1537 GND.n1536 0.152939
R16400 GND.n1565 GND.n1537 0.152939
R16401 GND.n1568 GND.n1565 0.152939
R16402 GND.n1569 GND.n1568 0.152939
R16403 GND.n1570 GND.n1569 0.152939
R16404 GND.n1571 GND.n1570 0.152939
R16405 GND.n1572 GND.n1571 0.152939
R16406 GND.n1608 GND.n1572 0.152939
R16407 GND.n1611 GND.n1608 0.152939
R16408 GND.n1612 GND.n1611 0.152939
R16409 GND.n1613 GND.n1612 0.152939
R16410 GND.n1614 GND.n1613 0.152939
R16411 GND.n1615 GND.n1614 0.152939
R16412 GND.n3411 GND.n1615 0.152939
R16413 GND.n3412 GND.n3411 0.152939
R16414 GND.n3414 GND.n3412 0.152939
R16415 GND.n3414 GND.n3413 0.152939
R16416 GND.n3413 GND.n1657 0.152939
R16417 GND.n1658 GND.n1657 0.152939
R16418 GND.n1659 GND.n1658 0.152939
R16419 GND.n3760 GND.n1659 0.152939
R16420 GND.n3761 GND.n3760 0.152939
R16421 GND.n3766 GND.n3761 0.152939
R16422 GND.n3767 GND.n3766 0.152939
R16423 GND.n3769 GND.n3767 0.152939
R16424 GND.n3769 GND.n3768 0.152939
R16425 GND.n3768 GND.n1701 0.152939
R16426 GND.n1702 GND.n1701 0.152939
R16427 GND.n1703 GND.n1702 0.152939
R16428 GND.n1726 GND.n1703 0.152939
R16429 GND.n1727 GND.n1726 0.152939
R16430 GND.n1728 GND.n1727 0.152939
R16431 GND.n1729 GND.n1728 0.152939
R16432 GND.n1730 GND.n1729 0.152939
R16433 GND.n1752 GND.n1730 0.152939
R16434 GND.n1753 GND.n1752 0.152939
R16435 GND.n1754 GND.n1753 0.152939
R16436 GND.n1755 GND.n1754 0.152939
R16437 GND.n1756 GND.n1755 0.152939
R16438 GND.n2123 GND.n1756 0.152939
R16439 GND.n2124 GND.n2123 0.152939
R16440 GND.n2130 GND.n2124 0.152939
R16441 GND.n2131 GND.n2130 0.152939
R16442 GND.n2132 GND.n2131 0.152939
R16443 GND.n2132 GND.n2119 0.152939
R16444 GND.n3847 GND.n2119 0.152939
R16445 GND.n3848 GND.n3847 0.152939
R16446 GND.n3849 GND.n3848 0.152939
R16447 GND.n3850 GND.n3849 0.152939
R16448 GND.n3851 GND.n3850 0.152939
R16449 GND.n3854 GND.n3851 0.152939
R16450 GND.n3855 GND.n3854 0.152939
R16451 GND.n3856 GND.n3855 0.152939
R16452 GND.n3857 GND.n3856 0.152939
R16453 GND.n3860 GND.n3857 0.152939
R16454 GND.n3861 GND.n3860 0.152939
R16455 GND.n3862 GND.n3861 0.152939
R16456 GND.n3863 GND.n3862 0.152939
R16457 GND.n3864 GND.n3863 0.152939
R16458 GND.n3865 GND.n3864 0.152939
R16459 GND.n3865 GND.n2047 0.152939
R16460 GND.n3968 GND.n2047 0.152939
R16461 GND.n3969 GND.n3968 0.152939
R16462 GND.n3970 GND.n3969 0.152939
R16463 GND.n3971 GND.n3970 0.152939
R16464 GND.n3972 GND.n3971 0.152939
R16465 GND.n2832 GND.n2831 0.152939
R16466 GND.n2832 GND.n2359 0.152939
R16467 GND.n2854 GND.n2359 0.152939
R16468 GND.n2855 GND.n2854 0.152939
R16469 GND.n2856 GND.n2855 0.152939
R16470 GND.n2857 GND.n2856 0.152939
R16471 GND.n2857 GND.n2340 0.152939
R16472 GND.n2879 GND.n2340 0.152939
R16473 GND.n2880 GND.n2879 0.152939
R16474 GND.n2881 GND.n2880 0.152939
R16475 GND.n2882 GND.n2881 0.152939
R16476 GND.n2882 GND.n2319 0.152939
R16477 GND.n2905 GND.n2319 0.152939
R16478 GND.n2906 GND.n2905 0.152939
R16479 GND.n2907 GND.n2906 0.152939
R16480 GND.n2907 GND.n2293 0.152939
R16481 GND.n2945 GND.n2293 0.152939
R16482 GND.n2946 GND.n2945 0.152939
R16483 GND.n2947 GND.n2946 0.152939
R16484 GND.n2947 GND.n1268 0.152939
R16485 GND.n4597 GND.n1268 0.152939
R16486 GND.n1116 GND.n1115 0.152939
R16487 GND.n1117 GND.n1116 0.152939
R16488 GND.n1118 GND.n1117 0.152939
R16489 GND.n1119 GND.n1118 0.152939
R16490 GND.n1120 GND.n1119 0.152939
R16491 GND.n1121 GND.n1120 0.152939
R16492 GND.n1122 GND.n1121 0.152939
R16493 GND.n1123 GND.n1122 0.152939
R16494 GND.n1124 GND.n1123 0.152939
R16495 GND.n1125 GND.n1124 0.152939
R16496 GND.n1126 GND.n1125 0.152939
R16497 GND.n1127 GND.n1126 0.152939
R16498 GND.n1128 GND.n1127 0.152939
R16499 GND.n1129 GND.n1128 0.152939
R16500 GND.n1130 GND.n1129 0.152939
R16501 GND.n1133 GND.n1130 0.152939
R16502 GND.n1134 GND.n1133 0.152939
R16503 GND.n1135 GND.n1134 0.152939
R16504 GND.n1136 GND.n1135 0.152939
R16505 GND.n1137 GND.n1136 0.152939
R16506 GND.n1138 GND.n1137 0.152939
R16507 GND.n1139 GND.n1138 0.152939
R16508 GND.n1140 GND.n1139 0.152939
R16509 GND.n1141 GND.n1140 0.152939
R16510 GND.n1142 GND.n1141 0.152939
R16511 GND.n1143 GND.n1142 0.152939
R16512 GND.n1144 GND.n1143 0.152939
R16513 GND.n1145 GND.n1144 0.152939
R16514 GND.n1146 GND.n1145 0.152939
R16515 GND.n1147 GND.n1146 0.152939
R16516 GND.n1148 GND.n1147 0.152939
R16517 GND.n4686 GND.n1148 0.152939
R16518 GND.n4686 GND.n4685 0.152939
R16519 GND.n4685 GND.n4684 0.152939
R16520 GND.n2548 GND.n2547 0.152939
R16521 GND.n2622 GND.n2547 0.152939
R16522 GND.n2623 GND.n2622 0.152939
R16523 GND.n2624 GND.n2623 0.152939
R16524 GND.n2625 GND.n2624 0.152939
R16525 GND.n2625 GND.n2489 0.152939
R16526 GND.n2647 GND.n2489 0.152939
R16527 GND.n2648 GND.n2647 0.152939
R16528 GND.n2649 GND.n2648 0.152939
R16529 GND.n2650 GND.n2649 0.152939
R16530 GND.n2650 GND.n2466 0.152939
R16531 GND.n2672 GND.n2466 0.152939
R16532 GND.n2673 GND.n2672 0.152939
R16533 GND.n2674 GND.n2673 0.152939
R16534 GND.n2675 GND.n2674 0.152939
R16535 GND.n2675 GND.n2443 0.152939
R16536 GND.n2709 GND.n2443 0.152939
R16537 GND.n2710 GND.n2709 0.152939
R16538 GND.n2711 GND.n2710 0.152939
R16539 GND.n2711 GND.n2380 0.152939
R16540 GND.n2831 GND.n2380 0.152939
R16541 GND.n2538 GND.n2507 0.152939
R16542 GND.n2510 GND.n2507 0.152939
R16543 GND.n2511 GND.n2510 0.152939
R16544 GND.n2512 GND.n2511 0.152939
R16545 GND.n2513 GND.n2512 0.152939
R16546 GND.n2516 GND.n2513 0.152939
R16547 GND.n2517 GND.n2516 0.152939
R16548 GND.n2518 GND.n2517 0.152939
R16549 GND.n2519 GND.n2518 0.152939
R16550 GND.n2520 GND.n2519 0.152939
R16551 GND.n2520 GND.n2431 0.152939
R16552 GND.n2719 GND.n2431 0.152939
R16553 GND.n2720 GND.n2719 0.152939
R16554 GND.n2721 GND.n2720 0.152939
R16555 GND.n4885 GND.n956 0.152939
R16556 GND.n961 GND.n956 0.152939
R16557 GND.n962 GND.n961 0.152939
R16558 GND.n963 GND.n962 0.152939
R16559 GND.n968 GND.n963 0.152939
R16560 GND.n969 GND.n968 0.152939
R16561 GND.n970 GND.n969 0.152939
R16562 GND.n971 GND.n970 0.152939
R16563 GND.n976 GND.n971 0.152939
R16564 GND.n977 GND.n976 0.152939
R16565 GND.n978 GND.n977 0.152939
R16566 GND.n979 GND.n978 0.152939
R16567 GND.n984 GND.n979 0.152939
R16568 GND.n985 GND.n984 0.152939
R16569 GND.n986 GND.n985 0.152939
R16570 GND.n987 GND.n986 0.152939
R16571 GND.n992 GND.n987 0.152939
R16572 GND.n993 GND.n992 0.152939
R16573 GND.n994 GND.n993 0.152939
R16574 GND.n995 GND.n994 0.152939
R16575 GND.n1000 GND.n995 0.152939
R16576 GND.n1001 GND.n1000 0.152939
R16577 GND.n1002 GND.n1001 0.152939
R16578 GND.n1003 GND.n1002 0.152939
R16579 GND.n1008 GND.n1003 0.152939
R16580 GND.n1009 GND.n1008 0.152939
R16581 GND.n1010 GND.n1009 0.152939
R16582 GND.n1011 GND.n1010 0.152939
R16583 GND.n1016 GND.n1011 0.152939
R16584 GND.n1017 GND.n1016 0.152939
R16585 GND.n1018 GND.n1017 0.152939
R16586 GND.n1019 GND.n1018 0.152939
R16587 GND.n1024 GND.n1019 0.152939
R16588 GND.n1025 GND.n1024 0.152939
R16589 GND.n1026 GND.n1025 0.152939
R16590 GND.n1027 GND.n1026 0.152939
R16591 GND.n1032 GND.n1027 0.152939
R16592 GND.n1033 GND.n1032 0.152939
R16593 GND.n1034 GND.n1033 0.152939
R16594 GND.n1035 GND.n1034 0.152939
R16595 GND.n1040 GND.n1035 0.152939
R16596 GND.n1041 GND.n1040 0.152939
R16597 GND.n1042 GND.n1041 0.152939
R16598 GND.n1043 GND.n1042 0.152939
R16599 GND.n1048 GND.n1043 0.152939
R16600 GND.n1049 GND.n1048 0.152939
R16601 GND.n1050 GND.n1049 0.152939
R16602 GND.n1051 GND.n1050 0.152939
R16603 GND.n1056 GND.n1051 0.152939
R16604 GND.n1057 GND.n1056 0.152939
R16605 GND.n1058 GND.n1057 0.152939
R16606 GND.n1059 GND.n1058 0.152939
R16607 GND.n1064 GND.n1059 0.152939
R16608 GND.n1065 GND.n1064 0.152939
R16609 GND.n1066 GND.n1065 0.152939
R16610 GND.n1067 GND.n1066 0.152939
R16611 GND.n1072 GND.n1067 0.152939
R16612 GND.n1073 GND.n1072 0.152939
R16613 GND.n1074 GND.n1073 0.152939
R16614 GND.n1075 GND.n1074 0.152939
R16615 GND.n1080 GND.n1075 0.152939
R16616 GND.n1081 GND.n1080 0.152939
R16617 GND.n1082 GND.n1081 0.152939
R16618 GND.n1083 GND.n1082 0.152939
R16619 GND.n2506 GND.n1083 0.152939
R16620 GND.n2539 GND.n2506 0.152939
R16621 GND.n3840 GND.n3838 0.152939
R16622 GND.n3840 GND.n3839 0.152939
R16623 GND.n3839 GND.n2099 0.152939
R16624 GND.n3906 GND.n2099 0.152939
R16625 GND.n3907 GND.n3906 0.152939
R16626 GND.n3909 GND.n3907 0.152939
R16627 GND.n3909 GND.n3908 0.152939
R16628 GND.n3908 GND.n2077 0.152939
R16629 GND.n3930 GND.n2077 0.152939
R16630 GND.n3931 GND.n3930 0.152939
R16631 GND.n3933 GND.n3931 0.152939
R16632 GND.n3933 GND.n3932 0.152939
R16633 GND.n3932 GND.n2055 0.152939
R16634 GND.n3955 GND.n2055 0.152939
R16635 GND.n3956 GND.n3955 0.152939
R16636 GND.n3960 GND.n3956 0.152939
R16637 GND.n3960 GND.n3959 0.152939
R16638 GND.n3959 GND.n3958 0.152939
R16639 GND.n3958 GND.n2021 0.152939
R16640 GND.n3994 GND.n2021 0.152939
R16641 GND.n3995 GND.n3994 0.152939
R16642 GND.n3999 GND.n3995 0.152939
R16643 GND.n3999 GND.n3998 0.152939
R16644 GND.n3998 GND.n3997 0.152939
R16645 GND.n3997 GND.n426 0.152939
R16646 GND.n5670 GND.n427 0.152939
R16647 GND.n5670 GND.n5669 0.152939
R16648 GND.n5669 GND.n5668 0.152939
R16649 GND.n5668 GND.n433 0.152939
R16650 GND.n5664 GND.n433 0.152939
R16651 GND.n5664 GND.n5663 0.152939
R16652 GND.n5663 GND.n5662 0.152939
R16653 GND.n5662 GND.n438 0.152939
R16654 GND.n5658 GND.n438 0.152939
R16655 GND.n5658 GND.n5657 0.152939
R16656 GND.n5657 GND.n5656 0.152939
R16657 GND.n5656 GND.n443 0.152939
R16658 GND.n5652 GND.n443 0.152939
R16659 GND.n5652 GND.n5651 0.152939
R16660 GND.n5651 GND.n5650 0.152939
R16661 GND.n5650 GND.n448 0.152939
R16662 GND.n5646 GND.n448 0.152939
R16663 GND.n5646 GND.n5645 0.152939
R16664 GND.n5645 GND.n5644 0.152939
R16665 GND.n5644 GND.n453 0.152939
R16666 GND.n5640 GND.n453 0.152939
R16667 GND.n5640 GND.n5639 0.152939
R16668 GND.n5639 GND.n5638 0.152939
R16669 GND.n5638 GND.n458 0.152939
R16670 GND.n5634 GND.n458 0.152939
R16671 GND.n5566 GND.n5565 0.152939
R16672 GND.n5565 GND.n5564 0.152939
R16673 GND.n5564 GND.n5525 0.152939
R16674 GND.n5560 GND.n5525 0.152939
R16675 GND.n5560 GND.n5559 0.152939
R16676 GND.n5559 GND.n5558 0.152939
R16677 GND.n5558 GND.n5531 0.152939
R16678 GND.n5554 GND.n5531 0.152939
R16679 GND.n5554 GND.n5553 0.152939
R16680 GND.n5553 GND.n5552 0.152939
R16681 GND.n5552 GND.n5537 0.152939
R16682 GND.n5548 GND.n5537 0.152939
R16683 GND.n5548 GND.n5547 0.152939
R16684 GND.n5547 GND.n5546 0.152939
R16685 GND.n5546 GND.n462 0.152939
R16686 GND.n5633 GND.n462 0.152939
R16687 GND.n5627 GND.n5626 0.152939
R16688 GND.n5626 GND.n5625 0.152939
R16689 GND.n5625 GND.n498 0.152939
R16690 GND.n5621 GND.n498 0.152939
R16691 GND.n5621 GND.n5620 0.152939
R16692 GND.n5620 GND.n5619 0.152939
R16693 GND.n5619 GND.n504 0.152939
R16694 GND.n5615 GND.n504 0.152939
R16695 GND.n5615 GND.n5614 0.152939
R16696 GND.n5614 GND.n5613 0.152939
R16697 GND.n5613 GND.n510 0.152939
R16698 GND.n5609 GND.n510 0.152939
R16699 GND.n5609 GND.n5608 0.152939
R16700 GND.n5608 GND.n5607 0.152939
R16701 GND.n5607 GND.n516 0.152939
R16702 GND.n5602 GND.n516 0.152939
R16703 GND.n5602 GND.n5601 0.152939
R16704 GND.n5601 GND.n5600 0.152939
R16705 GND.n5600 GND.n524 0.152939
R16706 GND.n5596 GND.n524 0.152939
R16707 GND.n5596 GND.n5595 0.152939
R16708 GND.n5595 GND.n5594 0.152939
R16709 GND.n5594 GND.n530 0.152939
R16710 GND.n5590 GND.n530 0.152939
R16711 GND.n5590 GND.n5589 0.152939
R16712 GND.n5589 GND.n5588 0.152939
R16713 GND.n5588 GND.n536 0.152939
R16714 GND.n5584 GND.n536 0.152939
R16715 GND.n5584 GND.n5583 0.152939
R16716 GND.n5583 GND.n5582 0.152939
R16717 GND.n5582 GND.n542 0.152939
R16718 GND.n5578 GND.n542 0.152939
R16719 GND.n5578 GND.n5577 0.152939
R16720 GND.n5577 GND.n5576 0.152939
R16721 GND.n3836 GND.n2141 0.152939
R16722 GND.n3832 GND.n2141 0.152939
R16723 GND.n3832 GND.n3831 0.152939
R16724 GND.n3831 GND.n3830 0.152939
R16725 GND.n3830 GND.n2148 0.152939
R16726 GND.n3826 GND.n2148 0.152939
R16727 GND.n3826 GND.n3825 0.152939
R16728 GND.n3825 GND.n3824 0.152939
R16729 GND.n3824 GND.n2154 0.152939
R16730 GND.n3819 GND.n2154 0.152939
R16731 GND.n3819 GND.n3818 0.152939
R16732 GND.n3818 GND.n3817 0.152939
R16733 GND.n3817 GND.n2162 0.152939
R16734 GND.n3002 GND.n2274 0.152939
R16735 GND.n3008 GND.n2274 0.152939
R16736 GND.n3009 GND.n3008 0.152939
R16737 GND.n3010 GND.n3009 0.152939
R16738 GND.n3010 GND.n2272 0.152939
R16739 GND.n3016 GND.n2272 0.152939
R16740 GND.n3017 GND.n3016 0.152939
R16741 GND.n3018 GND.n3017 0.152939
R16742 GND.n3018 GND.n2268 0.152939
R16743 GND.n3024 GND.n2268 0.152939
R16744 GND.n3025 GND.n3024 0.152939
R16745 GND.n3032 GND.n3025 0.152939
R16746 GND.n3032 GND.n3031 0.152939
R16747 GND.n3031 GND.n3030 0.152939
R16748 GND.n3030 GND.n3026 0.152939
R16749 GND.n3026 GND.n2237 0.152939
R16750 GND.n3251 GND.n2237 0.152939
R16751 GND.n3252 GND.n3251 0.152939
R16752 GND.n3269 GND.n3252 0.152939
R16753 GND.n3269 GND.n3268 0.152939
R16754 GND.n3268 GND.n3267 0.152939
R16755 GND.n3267 GND.n3253 0.152939
R16756 GND.n3263 GND.n3253 0.152939
R16757 GND.n3263 GND.n3262 0.152939
R16758 GND.n3262 GND.n3261 0.152939
R16759 GND.n3261 GND.n2213 0.152939
R16760 GND.n3323 GND.n2213 0.152939
R16761 GND.n3324 GND.n3323 0.152939
R16762 GND.n3346 GND.n3324 0.152939
R16763 GND.n3346 GND.n3345 0.152939
R16764 GND.n3345 GND.n3344 0.152939
R16765 GND.n3344 GND.n3325 0.152939
R16766 GND.n3340 GND.n3325 0.152939
R16767 GND.n3340 GND.n3339 0.152939
R16768 GND.n3339 GND.n3338 0.152939
R16769 GND.n3338 GND.n3331 0.152939
R16770 GND.n3334 GND.n3331 0.152939
R16771 GND.n3334 GND.n3333 0.152939
R16772 GND.n3333 GND.n2195 0.152939
R16773 GND.n3399 GND.n2195 0.152939
R16774 GND.n3400 GND.n3399 0.152939
R16775 GND.n3405 GND.n3400 0.152939
R16776 GND.n3405 GND.n3404 0.152939
R16777 GND.n3404 GND.n3403 0.152939
R16778 GND.n3403 GND.n2183 0.152939
R16779 GND.n3444 GND.n2183 0.152939
R16780 GND.n3445 GND.n3444 0.152939
R16781 GND.n3447 GND.n3445 0.152939
R16782 GND.n3447 GND.n3446 0.152939
R16783 GND.n3446 GND.n2175 0.152939
R16784 GND.n3784 GND.n2175 0.152939
R16785 GND.n3785 GND.n3784 0.152939
R16786 GND.n3786 GND.n3785 0.152939
R16787 GND.n3786 GND.n2173 0.152939
R16788 GND.n3792 GND.n2173 0.152939
R16789 GND.n3793 GND.n3792 0.152939
R16790 GND.n3794 GND.n3793 0.152939
R16791 GND.n3794 GND.n2169 0.152939
R16792 GND.n3800 GND.n2169 0.152939
R16793 GND.n3801 GND.n3800 0.152939
R16794 GND.n3802 GND.n3801 0.152939
R16795 GND.n3802 GND.n2167 0.152939
R16796 GND.n3809 GND.n2167 0.152939
R16797 GND.n3810 GND.n3809 0.152939
R16798 GND.n3811 GND.n3810 0.152939
R16799 GND.n2969 GND.n2281 0.152939
R16800 GND.n2970 GND.n2969 0.152939
R16801 GND.n2971 GND.n2970 0.152939
R16802 GND.n2971 GND.n2279 0.152939
R16803 GND.n2979 GND.n2279 0.152939
R16804 GND.n2980 GND.n2979 0.152939
R16805 GND.n2981 GND.n2980 0.152939
R16806 GND.n2981 GND.n2277 0.152939
R16807 GND.n2992 GND.n2277 0.152939
R16808 GND.n2993 GND.n2992 0.152939
R16809 GND.n2994 GND.n2993 0.152939
R16810 GND.n2994 GND.n2275 0.152939
R16811 GND.n3001 GND.n2275 0.152939
R16812 GND.n2742 GND.n2741 0.152939
R16813 GND.n2743 GND.n2742 0.152939
R16814 GND.n2743 GND.n2370 0.152939
R16815 GND.n2839 GND.n2370 0.152939
R16816 GND.n2840 GND.n2839 0.152939
R16817 GND.n2842 GND.n2840 0.152939
R16818 GND.n2842 GND.n2841 0.152939
R16819 GND.n2841 GND.n2350 0.152939
R16820 GND.n2864 GND.n2350 0.152939
R16821 GND.n2865 GND.n2864 0.152939
R16822 GND.n2867 GND.n2865 0.152939
R16823 GND.n2867 GND.n2866 0.152939
R16824 GND.n2866 GND.n2330 0.152939
R16825 GND.n2889 GND.n2330 0.152939
R16826 GND.n2890 GND.n2889 0.152939
R16827 GND.n2895 GND.n2890 0.152939
R16828 GND.n2895 GND.n2894 0.152939
R16829 GND.n2894 GND.n2893 0.152939
R16830 GND.n2893 GND.n2305 0.152939
R16831 GND.n2936 GND.n2305 0.152939
R16832 GND.n2936 GND.n2935 0.152939
R16833 GND.n2935 GND.n2934 0.152939
R16834 GND.n2934 GND.n2306 0.152939
R16835 GND.n2306 GND.n2286 0.152939
R16836 GND.n2959 GND.n2286 0.152939
R16837 GND.n4596 GND.n1269 0.152939
R16838 GND.n4592 GND.n1269 0.152939
R16839 GND.n4592 GND.n4591 0.152939
R16840 GND.n4591 GND.n4590 0.152939
R16841 GND.n4590 GND.n1273 0.152939
R16842 GND.n4586 GND.n1273 0.152939
R16843 GND.n4586 GND.n4585 0.152939
R16844 GND.n4585 GND.n4584 0.152939
R16845 GND.n4584 GND.n1278 0.152939
R16846 GND.n4580 GND.n1278 0.152939
R16847 GND.n4580 GND.n4579 0.152939
R16848 GND.n4579 GND.n4578 0.152939
R16849 GND.n4578 GND.n1283 0.152939
R16850 GND.n4573 GND.n4572 0.152939
R16851 GND.n4572 GND.n4571 0.152939
R16852 GND.n4571 GND.n1293 0.152939
R16853 GND.n4567 GND.n1293 0.152939
R16854 GND.n4567 GND.n4566 0.152939
R16855 GND.n4566 GND.n4565 0.152939
R16856 GND.n4565 GND.n1298 0.152939
R16857 GND.n4561 GND.n1298 0.152939
R16858 GND.n4561 GND.n4560 0.152939
R16859 GND.n4560 GND.n4559 0.152939
R16860 GND.n4559 GND.n1303 0.152939
R16861 GND.n4555 GND.n1303 0.152939
R16862 GND.n4555 GND.n4554 0.152939
R16863 GND.n4554 GND.n4553 0.152939
R16864 GND.n4553 GND.n1308 0.152939
R16865 GND.n4549 GND.n1308 0.152939
R16866 GND.n4549 GND.n4548 0.152939
R16867 GND.n4548 GND.n4547 0.152939
R16868 GND.n2610 GND.n2554 0.152939
R16869 GND.n2610 GND.n2609 0.152939
R16870 GND.n2609 GND.n2608 0.152939
R16871 GND.n2608 GND.n2558 0.152939
R16872 GND.n2604 GND.n2558 0.152939
R16873 GND.n2604 GND.n2603 0.152939
R16874 GND.n2603 GND.n2602 0.152939
R16875 GND.n2602 GND.n2564 0.152939
R16876 GND.n2598 GND.n2564 0.152939
R16877 GND.n2598 GND.n2597 0.152939
R16878 GND.n2597 GND.n2596 0.152939
R16879 GND.n2596 GND.n2570 0.152939
R16880 GND.n2592 GND.n2570 0.152939
R16881 GND.n2592 GND.n2591 0.152939
R16882 GND.n2591 GND.n2590 0.152939
R16883 GND.n2590 GND.n2584 0.152939
R16884 GND.n2583 GND.n2576 0.152939
R16885 GND.n2579 GND.n2576 0.152939
R16886 GND.n2579 GND.n2501 0.152939
R16887 GND.n2632 GND.n2501 0.152939
R16888 GND.n2633 GND.n2632 0.152939
R16889 GND.n2635 GND.n2633 0.152939
R16890 GND.n2635 GND.n2634 0.152939
R16891 GND.n2634 GND.n2478 0.152939
R16892 GND.n2657 GND.n2478 0.152939
R16893 GND.n2658 GND.n2657 0.152939
R16894 GND.n2660 GND.n2658 0.152939
R16895 GND.n2660 GND.n2659 0.152939
R16896 GND.n2659 GND.n2456 0.152939
R16897 GND.n2682 GND.n2456 0.152939
R16898 GND.n2683 GND.n2682 0.152939
R16899 GND.n2699 GND.n2683 0.152939
R16900 GND.n2699 GND.n2698 0.152939
R16901 GND.n2698 GND.n2697 0.152939
R16902 GND.n2697 GND.n2684 0.152939
R16903 GND.n2693 GND.n2684 0.152939
R16904 GND.n2693 GND.n2692 0.152939
R16905 GND.n2692 GND.n2423 0.152939
R16906 GND.n2733 GND.n2423 0.152939
R16907 GND.n2734 GND.n2733 0.152939
R16908 GND.n2735 GND.n2734 0.152939
R16909 GND.n4075 GND.n1984 0.146841
R16910 GND.n2721 GND.n2381 0.146841
R16911 GND.n5674 GND.n426 0.145814
R16912 GND.n5674 GND.n427 0.145814
R16913 GND.n2741 GND.n2421 0.145814
R16914 GND.n2735 GND.n2421 0.145814
R16915 GND.n3837 GND.n3836 0.145317
R16916 GND.n2960 GND.n2281 0.145317
R16917 GND.n4201 GND.n4200 0.128997
R16918 GND.n4545 GND.n4544 0.128997
R16919 GND.n4210 GND.n4201 0.0442063
R16920 GND.n4544 GND.n1315 0.0442063
R16921 GND.n4200 GND.n4199 0.0429592
R16922 GND.n5571 GND.n550 0.0429592
R16923 GND.n4679 GND.n1154 0.0429592
R16924 GND.n4545 GND.n1259 0.0429592
R16925 GND.n4210 GND.n4209 0.0349686
R16926 GND.n1320 GND.n1315 0.0349686
R16927 GND.n4199 GND.n1856 0.0344674
R16928 GND.n4195 GND.n1856 0.0344674
R16929 GND.n4195 GND.n4194 0.0344674
R16930 GND.n4194 GND.n4193 0.0344674
R16931 GND.n4193 GND.n1864 0.0344674
R16932 GND.n4189 GND.n1864 0.0344674
R16933 GND.n4189 GND.n4188 0.0344674
R16934 GND.n4188 GND.n4187 0.0344674
R16935 GND.n4187 GND.n1872 0.0344674
R16936 GND.n4183 GND.n1872 0.0344674
R16937 GND.n4183 GND.n4182 0.0344674
R16938 GND.n4182 GND.n4181 0.0344674
R16939 GND.n4181 GND.n1880 0.0344674
R16940 GND.n4177 GND.n1880 0.0344674
R16941 GND.n4177 GND.n4176 0.0344674
R16942 GND.n4176 GND.n4175 0.0344674
R16943 GND.n4175 GND.n1888 0.0344674
R16944 GND.n4171 GND.n1888 0.0344674
R16945 GND.n4171 GND.n4170 0.0344674
R16946 GND.n4170 GND.n4169 0.0344674
R16947 GND.n4169 GND.n1896 0.0344674
R16948 GND.n4165 GND.n1896 0.0344674
R16949 GND.n4165 GND.n4164 0.0344674
R16950 GND.n4164 GND.n4163 0.0344674
R16951 GND.n4163 GND.n1904 0.0344674
R16952 GND.n4159 GND.n1904 0.0344674
R16953 GND.n4159 GND.n4158 0.0344674
R16954 GND.n4158 GND.n4157 0.0344674
R16955 GND.n4157 GND.n1912 0.0344674
R16956 GND.n4153 GND.n1912 0.0344674
R16957 GND.n4153 GND.n4152 0.0344674
R16958 GND.n4152 GND.n4151 0.0344674
R16959 GND.n4151 GND.n1920 0.0344674
R16960 GND.n4147 GND.n1920 0.0344674
R16961 GND.n4147 GND.n4146 0.0344674
R16962 GND.n4146 GND.n4145 0.0344674
R16963 GND.n4145 GND.n1928 0.0344674
R16964 GND.n4141 GND.n1928 0.0344674
R16965 GND.n4141 GND.n4140 0.0344674
R16966 GND.n4140 GND.n4139 0.0344674
R16967 GND.n4139 GND.n1936 0.0344674
R16968 GND.n4135 GND.n1936 0.0344674
R16969 GND.n4135 GND.n4134 0.0344674
R16970 GND.n4134 GND.n588 0.0344674
R16971 GND.n5492 GND.n588 0.0344674
R16972 GND.n5492 GND.n591 0.0344674
R16973 GND.n591 GND.n590 0.0344674
R16974 GND.n590 GND.n568 0.0344674
R16975 GND.n5510 GND.n568 0.0344674
R16976 GND.n5510 GND.n569 0.0344674
R16977 GND.n569 GND.n553 0.0344674
R16978 GND.n5571 GND.n553 0.0344674
R16979 GND.n4208 GND.n1779 0.0344674
R16980 GND.n2140 GND.n1819 0.0344674
R16981 GND.n4540 GND.n4539 0.0344674
R16982 GND.n2961 GND.n2285 0.0344674
R16983 GND.n4679 GND.n4678 0.0344674
R16984 GND.n4678 GND.n4677 0.0344674
R16985 GND.n4677 GND.n1160 0.0344674
R16986 GND.n4673 GND.n1160 0.0344674
R16987 GND.n4673 GND.n4672 0.0344674
R16988 GND.n4672 GND.n4671 0.0344674
R16989 GND.n4671 GND.n1168 0.0344674
R16990 GND.n4667 GND.n1168 0.0344674
R16991 GND.n4667 GND.n4666 0.0344674
R16992 GND.n4666 GND.n4665 0.0344674
R16993 GND.n4665 GND.n1176 0.0344674
R16994 GND.n4661 GND.n1176 0.0344674
R16995 GND.n4661 GND.n4660 0.0344674
R16996 GND.n4660 GND.n4659 0.0344674
R16997 GND.n4659 GND.n1184 0.0344674
R16998 GND.n4655 GND.n1184 0.0344674
R16999 GND.n4655 GND.n4654 0.0344674
R17000 GND.n4654 GND.n4653 0.0344674
R17001 GND.n4653 GND.n1192 0.0344674
R17002 GND.n4649 GND.n1192 0.0344674
R17003 GND.n4649 GND.n4648 0.0344674
R17004 GND.n4648 GND.n4647 0.0344674
R17005 GND.n4647 GND.n1200 0.0344674
R17006 GND.n4643 GND.n1200 0.0344674
R17007 GND.n4643 GND.n4642 0.0344674
R17008 GND.n4642 GND.n4641 0.0344674
R17009 GND.n4641 GND.n1208 0.0344674
R17010 GND.n4637 GND.n1208 0.0344674
R17011 GND.n4637 GND.n4636 0.0344674
R17012 GND.n4636 GND.n4635 0.0344674
R17013 GND.n4635 GND.n1216 0.0344674
R17014 GND.n4631 GND.n1216 0.0344674
R17015 GND.n4631 GND.n4630 0.0344674
R17016 GND.n4630 GND.n4629 0.0344674
R17017 GND.n4629 GND.n1224 0.0344674
R17018 GND.n4625 GND.n1224 0.0344674
R17019 GND.n4625 GND.n4624 0.0344674
R17020 GND.n4624 GND.n4623 0.0344674
R17021 GND.n4623 GND.n1232 0.0344674
R17022 GND.n4619 GND.n1232 0.0344674
R17023 GND.n4619 GND.n4618 0.0344674
R17024 GND.n4618 GND.n4617 0.0344674
R17025 GND.n4617 GND.n1240 0.0344674
R17026 GND.n4613 GND.n1240 0.0344674
R17027 GND.n4613 GND.n4612 0.0344674
R17028 GND.n4612 GND.n4611 0.0344674
R17029 GND.n4611 GND.n1248 0.0344674
R17030 GND.n4607 GND.n1248 0.0344674
R17031 GND.n4607 GND.n4606 0.0344674
R17032 GND.n4606 GND.n4605 0.0344674
R17033 GND.n4605 GND.n1256 0.0344674
R17034 GND.n1259 GND.n1256 0.0344674
R17035 GND.n4251 GND.n4250 0.0188424
R17036 GND.n4247 GND.n1780 0.0188424
R17037 GND.n4246 GND.n1785 0.0188424
R17038 GND.n4243 GND.n4242 0.0188424
R17039 GND.n4239 GND.n1789 0.0188424
R17040 GND.n4238 GND.n1793 0.0188424
R17041 GND.n4235 GND.n4234 0.0188424
R17042 GND.n4231 GND.n1799 0.0188424
R17043 GND.n4230 GND.n1803 0.0188424
R17044 GND.n4227 GND.n4226 0.0188424
R17045 GND.n4223 GND.n1807 0.0188424
R17046 GND.n4222 GND.n1813 0.0188424
R17047 GND.n4219 GND.n4218 0.0188424
R17048 GND.n4538 GND.n1321 0.0188424
R17049 GND.n1343 GND.n1342 0.0188424
R17050 GND.n4531 GND.n4530 0.0188424
R17051 GND.n4527 GND.n1344 0.0188424
R17052 GND.n4526 GND.n1349 0.0188424
R17053 GND.n4523 GND.n4522 0.0188424
R17054 GND.n4519 GND.n1353 0.0188424
R17055 GND.n4518 GND.n1357 0.0188424
R17056 GND.n4515 GND.n4514 0.0188424
R17057 GND.n4511 GND.n1363 0.0188424
R17058 GND.n4510 GND.n1367 0.0188424
R17059 GND.n4507 GND.n4506 0.0188424
R17060 GND.n1375 GND.n1371 0.0188424
R17061 GND.n4251 GND.n1779 0.016125
R17062 GND.n4250 GND.n1780 0.016125
R17063 GND.n4247 GND.n4246 0.016125
R17064 GND.n4243 GND.n1785 0.016125
R17065 GND.n4242 GND.n1789 0.016125
R17066 GND.n4239 GND.n4238 0.016125
R17067 GND.n4235 GND.n1793 0.016125
R17068 GND.n4234 GND.n1799 0.016125
R17069 GND.n4231 GND.n4230 0.016125
R17070 GND.n4227 GND.n1803 0.016125
R17071 GND.n4226 GND.n1807 0.016125
R17072 GND.n4223 GND.n4222 0.016125
R17073 GND.n4219 GND.n1813 0.016125
R17074 GND.n4218 GND.n1819 0.016125
R17075 GND.n4539 GND.n4538 0.016125
R17076 GND.n1342 GND.n1321 0.016125
R17077 GND.n4531 GND.n1343 0.016125
R17078 GND.n4530 GND.n1344 0.016125
R17079 GND.n4527 GND.n4526 0.016125
R17080 GND.n4523 GND.n1349 0.016125
R17081 GND.n4522 GND.n1353 0.016125
R17082 GND.n4519 GND.n4518 0.016125
R17083 GND.n4515 GND.n1357 0.016125
R17084 GND.n4514 GND.n1363 0.016125
R17085 GND.n4511 GND.n4510 0.016125
R17086 GND.n4507 GND.n1367 0.016125
R17087 GND.n4506 GND.n1371 0.016125
R17088 GND.n2285 GND.n1375 0.016125
R17089 GND.n2751 GND.n2381 0.00659756
R17090 GND.n3972 GND.n1984 0.00659756
R17091 GND.n4209 GND.n4208 0.00457609
R17092 GND.n4540 GND.n1320 0.00457609
R17093 GND.n3837 GND.n2140 0.00219837
R17094 GND.n2961 GND.n2960 0.00219837
R17095 CS_BIAS.n201 CS_BIAS.n139 161.3
R17096 CS_BIAS.n200 CS_BIAS.n199 161.3
R17097 CS_BIAS.n198 CS_BIAS.n140 161.3
R17098 CS_BIAS.n197 CS_BIAS.n196 161.3
R17099 CS_BIAS.n194 CS_BIAS.n141 161.3
R17100 CS_BIAS.n193 CS_BIAS.n192 161.3
R17101 CS_BIAS.n191 CS_BIAS.n142 161.3
R17102 CS_BIAS.n190 CS_BIAS.n189 161.3
R17103 CS_BIAS.n188 CS_BIAS.n143 161.3
R17104 CS_BIAS.n186 CS_BIAS.n185 161.3
R17105 CS_BIAS.n184 CS_BIAS.n144 161.3
R17106 CS_BIAS.n183 CS_BIAS.n182 161.3
R17107 CS_BIAS.n181 CS_BIAS.n145 161.3
R17108 CS_BIAS.n180 CS_BIAS.n179 161.3
R17109 CS_BIAS.n178 CS_BIAS.n177 161.3
R17110 CS_BIAS.n176 CS_BIAS.n147 161.3
R17111 CS_BIAS.n175 CS_BIAS.n174 161.3
R17112 CS_BIAS.n173 CS_BIAS.n148 161.3
R17113 CS_BIAS.n172 CS_BIAS.n171 161.3
R17114 CS_BIAS.n170 CS_BIAS.n149 161.3
R17115 CS_BIAS.n169 CS_BIAS.n168 161.3
R17116 CS_BIAS.n167 CS_BIAS.n151 161.3
R17117 CS_BIAS.n166 CS_BIAS.n165 161.3
R17118 CS_BIAS.n163 CS_BIAS.n152 161.3
R17119 CS_BIAS.n162 CS_BIAS.n161 161.3
R17120 CS_BIAS.n160 CS_BIAS.n153 161.3
R17121 CS_BIAS.n159 CS_BIAS.n158 161.3
R17122 CS_BIAS.n157 CS_BIAS.n154 161.3
R17123 CS_BIAS.n28 CS_BIAS.n25 161.3
R17124 CS_BIAS.n30 CS_BIAS.n29 161.3
R17125 CS_BIAS.n31 CS_BIAS.n24 161.3
R17126 CS_BIAS.n33 CS_BIAS.n32 161.3
R17127 CS_BIAS.n34 CS_BIAS.n23 161.3
R17128 CS_BIAS.n37 CS_BIAS.n36 161.3
R17129 CS_BIAS.n38 CS_BIAS.n22 161.3
R17130 CS_BIAS.n40 CS_BIAS.n39 161.3
R17131 CS_BIAS.n41 CS_BIAS.n20 161.3
R17132 CS_BIAS.n43 CS_BIAS.n42 161.3
R17133 CS_BIAS.n44 CS_BIAS.n19 161.3
R17134 CS_BIAS.n46 CS_BIAS.n45 161.3
R17135 CS_BIAS.n47 CS_BIAS.n18 161.3
R17136 CS_BIAS.n49 CS_BIAS.n48 161.3
R17137 CS_BIAS.n51 CS_BIAS.n50 161.3
R17138 CS_BIAS.n52 CS_BIAS.n16 161.3
R17139 CS_BIAS.n54 CS_BIAS.n53 161.3
R17140 CS_BIAS.n55 CS_BIAS.n15 161.3
R17141 CS_BIAS.n57 CS_BIAS.n56 161.3
R17142 CS_BIAS.n59 CS_BIAS.n14 161.3
R17143 CS_BIAS.n61 CS_BIAS.n60 161.3
R17144 CS_BIAS.n62 CS_BIAS.n13 161.3
R17145 CS_BIAS.n64 CS_BIAS.n63 161.3
R17146 CS_BIAS.n65 CS_BIAS.n12 161.3
R17147 CS_BIAS.n68 CS_BIAS.n67 161.3
R17148 CS_BIAS.n69 CS_BIAS.n11 161.3
R17149 CS_BIAS.n71 CS_BIAS.n70 161.3
R17150 CS_BIAS.n72 CS_BIAS.n10 161.3
R17151 CS_BIAS.n92 CS_BIAS.n89 161.3
R17152 CS_BIAS.n94 CS_BIAS.n93 161.3
R17153 CS_BIAS.n95 CS_BIAS.n88 161.3
R17154 CS_BIAS.n97 CS_BIAS.n96 161.3
R17155 CS_BIAS.n98 CS_BIAS.n87 161.3
R17156 CS_BIAS.n101 CS_BIAS.n100 161.3
R17157 CS_BIAS.n102 CS_BIAS.n86 161.3
R17158 CS_BIAS.n104 CS_BIAS.n103 161.3
R17159 CS_BIAS.n105 CS_BIAS.n84 161.3
R17160 CS_BIAS.n107 CS_BIAS.n106 161.3
R17161 CS_BIAS.n108 CS_BIAS.n9 161.3
R17162 CS_BIAS.n110 CS_BIAS.n109 161.3
R17163 CS_BIAS.n111 CS_BIAS.n8 161.3
R17164 CS_BIAS.n113 CS_BIAS.n112 161.3
R17165 CS_BIAS.n115 CS_BIAS.n114 161.3
R17166 CS_BIAS.n116 CS_BIAS.n6 161.3
R17167 CS_BIAS.n118 CS_BIAS.n117 161.3
R17168 CS_BIAS.n119 CS_BIAS.n5 161.3
R17169 CS_BIAS.n121 CS_BIAS.n120 161.3
R17170 CS_BIAS.n123 CS_BIAS.n4 161.3
R17171 CS_BIAS.n125 CS_BIAS.n124 161.3
R17172 CS_BIAS.n126 CS_BIAS.n3 161.3
R17173 CS_BIAS.n128 CS_BIAS.n127 161.3
R17174 CS_BIAS.n129 CS_BIAS.n2 161.3
R17175 CS_BIAS.n132 CS_BIAS.n131 161.3
R17176 CS_BIAS.n133 CS_BIAS.n1 161.3
R17177 CS_BIAS.n135 CS_BIAS.n134 161.3
R17178 CS_BIAS.n136 CS_BIAS.n0 161.3
R17179 CS_BIAS.n406 CS_BIAS.n344 161.3
R17180 CS_BIAS.n405 CS_BIAS.n404 161.3
R17181 CS_BIAS.n403 CS_BIAS.n345 161.3
R17182 CS_BIAS.n402 CS_BIAS.n401 161.3
R17183 CS_BIAS.n399 CS_BIAS.n346 161.3
R17184 CS_BIAS.n398 CS_BIAS.n397 161.3
R17185 CS_BIAS.n396 CS_BIAS.n347 161.3
R17186 CS_BIAS.n395 CS_BIAS.n394 161.3
R17187 CS_BIAS.n393 CS_BIAS.n348 161.3
R17188 CS_BIAS.n391 CS_BIAS.n390 161.3
R17189 CS_BIAS.n389 CS_BIAS.n349 161.3
R17190 CS_BIAS.n388 CS_BIAS.n387 161.3
R17191 CS_BIAS.n386 CS_BIAS.n350 161.3
R17192 CS_BIAS.n385 CS_BIAS.n384 161.3
R17193 CS_BIAS.n383 CS_BIAS.n382 161.3
R17194 CS_BIAS.n381 CS_BIAS.n352 161.3
R17195 CS_BIAS.n380 CS_BIAS.n379 161.3
R17196 CS_BIAS.n378 CS_BIAS.n353 161.3
R17197 CS_BIAS.n377 CS_BIAS.n376 161.3
R17198 CS_BIAS.n374 CS_BIAS.n354 161.3
R17199 CS_BIAS.n373 CS_BIAS.n372 161.3
R17200 CS_BIAS.n371 CS_BIAS.n355 161.3
R17201 CS_BIAS.n370 CS_BIAS.n369 161.3
R17202 CS_BIAS.n367 CS_BIAS.n356 161.3
R17203 CS_BIAS.n366 CS_BIAS.n365 161.3
R17204 CS_BIAS.n364 CS_BIAS.n357 161.3
R17205 CS_BIAS.n363 CS_BIAS.n362 161.3
R17206 CS_BIAS.n361 CS_BIAS.n358 161.3
R17207 CS_BIAS.n305 CS_BIAS.n243 161.3
R17208 CS_BIAS.n304 CS_BIAS.n303 161.3
R17209 CS_BIAS.n302 CS_BIAS.n244 161.3
R17210 CS_BIAS.n301 CS_BIAS.n300 161.3
R17211 CS_BIAS.n298 CS_BIAS.n245 161.3
R17212 CS_BIAS.n297 CS_BIAS.n296 161.3
R17213 CS_BIAS.n295 CS_BIAS.n246 161.3
R17214 CS_BIAS.n294 CS_BIAS.n293 161.3
R17215 CS_BIAS.n292 CS_BIAS.n247 161.3
R17216 CS_BIAS.n290 CS_BIAS.n289 161.3
R17217 CS_BIAS.n288 CS_BIAS.n248 161.3
R17218 CS_BIAS.n287 CS_BIAS.n286 161.3
R17219 CS_BIAS.n285 CS_BIAS.n249 161.3
R17220 CS_BIAS.n284 CS_BIAS.n283 161.3
R17221 CS_BIAS.n282 CS_BIAS.n281 161.3
R17222 CS_BIAS.n280 CS_BIAS.n251 161.3
R17223 CS_BIAS.n279 CS_BIAS.n278 161.3
R17224 CS_BIAS.n277 CS_BIAS.n252 161.3
R17225 CS_BIAS.n276 CS_BIAS.n275 161.3
R17226 CS_BIAS.n273 CS_BIAS.n253 161.3
R17227 CS_BIAS.n272 CS_BIAS.n271 161.3
R17228 CS_BIAS.n270 CS_BIAS.n254 161.3
R17229 CS_BIAS.n269 CS_BIAS.n268 161.3
R17230 CS_BIAS.n266 CS_BIAS.n255 161.3
R17231 CS_BIAS.n265 CS_BIAS.n264 161.3
R17232 CS_BIAS.n263 CS_BIAS.n256 161.3
R17233 CS_BIAS.n262 CS_BIAS.n261 161.3
R17234 CS_BIAS.n260 CS_BIAS.n257 161.3
R17235 CS_BIAS.n315 CS_BIAS.n314 161.3
R17236 CS_BIAS.n239 CS_BIAS.n214 161.3
R17237 CS_BIAS.n238 CS_BIAS.n237 161.3
R17238 CS_BIAS.n235 CS_BIAS.n215 161.3
R17239 CS_BIAS.n234 CS_BIAS.n233 161.3
R17240 CS_BIAS.n232 CS_BIAS.n216 161.3
R17241 CS_BIAS.n231 CS_BIAS.n230 161.3
R17242 CS_BIAS.n228 CS_BIAS.n217 161.3
R17243 CS_BIAS.n227 CS_BIAS.n226 161.3
R17244 CS_BIAS.n225 CS_BIAS.n218 161.3
R17245 CS_BIAS.n224 CS_BIAS.n223 161.3
R17246 CS_BIAS.n222 CS_BIAS.n219 161.3
R17247 CS_BIAS.n341 CS_BIAS.n205 161.3
R17248 CS_BIAS.n340 CS_BIAS.n339 161.3
R17249 CS_BIAS.n338 CS_BIAS.n206 161.3
R17250 CS_BIAS.n337 CS_BIAS.n336 161.3
R17251 CS_BIAS.n334 CS_BIAS.n207 161.3
R17252 CS_BIAS.n333 CS_BIAS.n332 161.3
R17253 CS_BIAS.n331 CS_BIAS.n208 161.3
R17254 CS_BIAS.n330 CS_BIAS.n329 161.3
R17255 CS_BIAS.n328 CS_BIAS.n209 161.3
R17256 CS_BIAS.n326 CS_BIAS.n325 161.3
R17257 CS_BIAS.n324 CS_BIAS.n210 161.3
R17258 CS_BIAS.n323 CS_BIAS.n322 161.3
R17259 CS_BIAS.n321 CS_BIAS.n211 161.3
R17260 CS_BIAS.n320 CS_BIAS.n319 161.3
R17261 CS_BIAS.n318 CS_BIAS.n317 161.3
R17262 CS_BIAS.n316 CS_BIAS.n213 161.3
R17263 CS_BIAS.n155 CS_BIAS.t60 102.697
R17264 CS_BIAS.n359 CS_BIAS.t39 102.697
R17265 CS_BIAS.n258 CS_BIAS.t12 102.697
R17266 CS_BIAS.n220 CS_BIAS.t32 102.697
R17267 CS_BIAS.n26 CS_BIAS.t14 102.697
R17268 CS_BIAS.n90 CS_BIAS.t54 102.697
R17269 CS_BIAS.n203 CS_BIAS.n202 90.9889
R17270 CS_BIAS.n74 CS_BIAS.n73 90.9889
R17271 CS_BIAS.n138 CS_BIAS.n137 90.9889
R17272 CS_BIAS.n408 CS_BIAS.n407 90.9889
R17273 CS_BIAS.n307 CS_BIAS.n306 90.9889
R17274 CS_BIAS.n343 CS_BIAS.n342 90.9889
R17275 CS_BIAS.n81 CS_BIAS.n79 85.0679
R17276 CS_BIAS.n242 CS_BIAS.n240 85.0679
R17277 CS_BIAS.n81 CS_BIAS.n80 84.0635
R17278 CS_BIAS.n78 CS_BIAS.n77 84.0635
R17279 CS_BIAS.n76 CS_BIAS.n75 84.0635
R17280 CS_BIAS.n309 CS_BIAS.n308 84.0635
R17281 CS_BIAS.n311 CS_BIAS.n310 84.0635
R17282 CS_BIAS.n242 CS_BIAS.n241 84.0635
R17283 CS_BIAS.n156 CS_BIAS.t57 72.3005
R17284 CS_BIAS.n164 CS_BIAS.t35 72.3005
R17285 CS_BIAS.n150 CS_BIAS.t34 72.3005
R17286 CS_BIAS.n146 CS_BIAS.t52 72.3005
R17287 CS_BIAS.n187 CS_BIAS.t55 72.3005
R17288 CS_BIAS.n195 CS_BIAS.t51 72.3005
R17289 CS_BIAS.n202 CS_BIAS.t38 72.3005
R17290 CS_BIAS.n73 CS_BIAS.t18 72.3005
R17291 CS_BIAS.n66 CS_BIAS.t24 72.3005
R17292 CS_BIAS.n58 CS_BIAS.t10 72.3005
R17293 CS_BIAS.n17 CS_BIAS.t2 72.3005
R17294 CS_BIAS.n21 CS_BIAS.t20 72.3005
R17295 CS_BIAS.n35 CS_BIAS.t0 72.3005
R17296 CS_BIAS.n27 CS_BIAS.t26 72.3005
R17297 CS_BIAS.n137 CS_BIAS.t63 72.3005
R17298 CS_BIAS.n130 CS_BIAS.t44 72.3005
R17299 CS_BIAS.n122 CS_BIAS.t46 72.3005
R17300 CS_BIAS.n7 CS_BIAS.t45 72.3005
R17301 CS_BIAS.n85 CS_BIAS.t61 72.3005
R17302 CS_BIAS.n99 CS_BIAS.t62 72.3005
R17303 CS_BIAS.n91 CS_BIAS.t50 72.3005
R17304 CS_BIAS.n360 CS_BIAS.t47 72.3005
R17305 CS_BIAS.n368 CS_BIAS.t58 72.3005
R17306 CS_BIAS.n375 CS_BIAS.t56 72.3005
R17307 CS_BIAS.n351 CS_BIAS.t42 72.3005
R17308 CS_BIAS.n392 CS_BIAS.t33 72.3005
R17309 CS_BIAS.n400 CS_BIAS.t41 72.3005
R17310 CS_BIAS.n407 CS_BIAS.t48 72.3005
R17311 CS_BIAS.n259 CS_BIAS.t30 72.3005
R17312 CS_BIAS.n267 CS_BIAS.t4 72.3005
R17313 CS_BIAS.n274 CS_BIAS.t22 72.3005
R17314 CS_BIAS.n250 CS_BIAS.t6 72.3005
R17315 CS_BIAS.n291 CS_BIAS.t8 72.3005
R17316 CS_BIAS.n299 CS_BIAS.t28 72.3005
R17317 CS_BIAS.n306 CS_BIAS.t16 72.3005
R17318 CS_BIAS.n342 CS_BIAS.t43 72.3005
R17319 CS_BIAS.n335 CS_BIAS.t37 72.3005
R17320 CS_BIAS.n327 CS_BIAS.t59 72.3005
R17321 CS_BIAS.n212 CS_BIAS.t36 72.3005
R17322 CS_BIAS.n221 CS_BIAS.t40 72.3005
R17323 CS_BIAS.n229 CS_BIAS.t53 72.3005
R17324 CS_BIAS.n236 CS_BIAS.t49 72.3005
R17325 CS_BIAS.n27 CS_BIAS.n26 66.3065
R17326 CS_BIAS.n91 CS_BIAS.n90 66.3065
R17327 CS_BIAS.n156 CS_BIAS.n155 66.3065
R17328 CS_BIAS.n360 CS_BIAS.n359 66.3065
R17329 CS_BIAS.n259 CS_BIAS.n258 66.3065
R17330 CS_BIAS.n221 CS_BIAS.n220 66.3065
R17331 CS_BIAS.n176 CS_BIAS.n175 56.5617
R17332 CS_BIAS.n200 CS_BIAS.n140 56.5617
R17333 CS_BIAS.n47 CS_BIAS.n46 56.5617
R17334 CS_BIAS.n111 CS_BIAS.n110 56.5617
R17335 CS_BIAS.n381 CS_BIAS.n380 56.5617
R17336 CS_BIAS.n405 CS_BIAS.n345 56.5617
R17337 CS_BIAS.n280 CS_BIAS.n279 56.5617
R17338 CS_BIAS.n304 CS_BIAS.n244 56.5617
R17339 CS_BIAS.n316 CS_BIAS.n315 56.5617
R17340 CS_BIAS.n71 CS_BIAS.n11 56.5617
R17341 CS_BIAS.n135 CS_BIAS.n1 56.5617
R17342 CS_BIAS.n340 CS_BIAS.n206 56.5617
R17343 CS_BIAS.n162 CS_BIAS.n153 49.296
R17344 CS_BIAS.n189 CS_BIAS.n142 49.296
R17345 CS_BIAS.n60 CS_BIAS.n13 49.296
R17346 CS_BIAS.n33 CS_BIAS.n24 49.296
R17347 CS_BIAS.n124 CS_BIAS.n3 49.296
R17348 CS_BIAS.n97 CS_BIAS.n88 49.296
R17349 CS_BIAS.n366 CS_BIAS.n357 49.296
R17350 CS_BIAS.n394 CS_BIAS.n347 49.296
R17351 CS_BIAS.n265 CS_BIAS.n256 49.296
R17352 CS_BIAS.n293 CS_BIAS.n246 49.296
R17353 CS_BIAS.n329 CS_BIAS.n208 49.296
R17354 CS_BIAS.n227 CS_BIAS.n218 49.296
R17355 CS_BIAS.n169 CS_BIAS.n151 48.3272
R17356 CS_BIAS.n182 CS_BIAS.n144 48.3272
R17357 CS_BIAS.n53 CS_BIAS.n15 48.3272
R17358 CS_BIAS.n40 CS_BIAS.n22 48.3272
R17359 CS_BIAS.n117 CS_BIAS.n5 48.3272
R17360 CS_BIAS.n104 CS_BIAS.n86 48.3272
R17361 CS_BIAS.n373 CS_BIAS.n355 48.3272
R17362 CS_BIAS.n387 CS_BIAS.n349 48.3272
R17363 CS_BIAS.n272 CS_BIAS.n254 48.3272
R17364 CS_BIAS.n286 CS_BIAS.n248 48.3272
R17365 CS_BIAS.n322 CS_BIAS.n210 48.3272
R17366 CS_BIAS.n234 CS_BIAS.n216 48.3272
R17367 CS_BIAS.n170 CS_BIAS.n169 32.8269
R17368 CS_BIAS.n182 CS_BIAS.n181 32.8269
R17369 CS_BIAS.n53 CS_BIAS.n52 32.8269
R17370 CS_BIAS.n41 CS_BIAS.n40 32.8269
R17371 CS_BIAS.n117 CS_BIAS.n116 32.8269
R17372 CS_BIAS.n105 CS_BIAS.n104 32.8269
R17373 CS_BIAS.n374 CS_BIAS.n373 32.8269
R17374 CS_BIAS.n387 CS_BIAS.n386 32.8269
R17375 CS_BIAS.n273 CS_BIAS.n272 32.8269
R17376 CS_BIAS.n286 CS_BIAS.n285 32.8269
R17377 CS_BIAS.n322 CS_BIAS.n321 32.8269
R17378 CS_BIAS.n235 CS_BIAS.n234 32.8269
R17379 CS_BIAS.n158 CS_BIAS.n153 31.8581
R17380 CS_BIAS.n193 CS_BIAS.n142 31.8581
R17381 CS_BIAS.n64 CS_BIAS.n13 31.8581
R17382 CS_BIAS.n29 CS_BIAS.n24 31.8581
R17383 CS_BIAS.n128 CS_BIAS.n3 31.8581
R17384 CS_BIAS.n93 CS_BIAS.n88 31.8581
R17385 CS_BIAS.n362 CS_BIAS.n357 31.8581
R17386 CS_BIAS.n398 CS_BIAS.n347 31.8581
R17387 CS_BIAS.n261 CS_BIAS.n256 31.8581
R17388 CS_BIAS.n297 CS_BIAS.n246 31.8581
R17389 CS_BIAS.n333 CS_BIAS.n208 31.8581
R17390 CS_BIAS.n223 CS_BIAS.n218 31.8581
R17391 CS_BIAS.n158 CS_BIAS.n157 24.5923
R17392 CS_BIAS.n165 CS_BIAS.n151 24.5923
R17393 CS_BIAS.n163 CS_BIAS.n162 24.5923
R17394 CS_BIAS.n175 CS_BIAS.n148 24.5923
R17395 CS_BIAS.n171 CS_BIAS.n170 24.5923
R17396 CS_BIAS.n181 CS_BIAS.n180 24.5923
R17397 CS_BIAS.n177 CS_BIAS.n176 24.5923
R17398 CS_BIAS.n189 CS_BIAS.n188 24.5923
R17399 CS_BIAS.n186 CS_BIAS.n144 24.5923
R17400 CS_BIAS.n196 CS_BIAS.n140 24.5923
R17401 CS_BIAS.n194 CS_BIAS.n193 24.5923
R17402 CS_BIAS.n201 CS_BIAS.n200 24.5923
R17403 CS_BIAS.n72 CS_BIAS.n71 24.5923
R17404 CS_BIAS.n67 CS_BIAS.n11 24.5923
R17405 CS_BIAS.n65 CS_BIAS.n64 24.5923
R17406 CS_BIAS.n60 CS_BIAS.n59 24.5923
R17407 CS_BIAS.n57 CS_BIAS.n15 24.5923
R17408 CS_BIAS.n52 CS_BIAS.n51 24.5923
R17409 CS_BIAS.n48 CS_BIAS.n47 24.5923
R17410 CS_BIAS.n46 CS_BIAS.n19 24.5923
R17411 CS_BIAS.n42 CS_BIAS.n41 24.5923
R17412 CS_BIAS.n36 CS_BIAS.n22 24.5923
R17413 CS_BIAS.n34 CS_BIAS.n33 24.5923
R17414 CS_BIAS.n29 CS_BIAS.n28 24.5923
R17415 CS_BIAS.n136 CS_BIAS.n135 24.5923
R17416 CS_BIAS.n131 CS_BIAS.n1 24.5923
R17417 CS_BIAS.n129 CS_BIAS.n128 24.5923
R17418 CS_BIAS.n124 CS_BIAS.n123 24.5923
R17419 CS_BIAS.n121 CS_BIAS.n5 24.5923
R17420 CS_BIAS.n116 CS_BIAS.n115 24.5923
R17421 CS_BIAS.n112 CS_BIAS.n111 24.5923
R17422 CS_BIAS.n110 CS_BIAS.n9 24.5923
R17423 CS_BIAS.n106 CS_BIAS.n105 24.5923
R17424 CS_BIAS.n100 CS_BIAS.n86 24.5923
R17425 CS_BIAS.n98 CS_BIAS.n97 24.5923
R17426 CS_BIAS.n93 CS_BIAS.n92 24.5923
R17427 CS_BIAS.n362 CS_BIAS.n361 24.5923
R17428 CS_BIAS.n367 CS_BIAS.n366 24.5923
R17429 CS_BIAS.n369 CS_BIAS.n355 24.5923
R17430 CS_BIAS.n376 CS_BIAS.n374 24.5923
R17431 CS_BIAS.n380 CS_BIAS.n353 24.5923
R17432 CS_BIAS.n382 CS_BIAS.n381 24.5923
R17433 CS_BIAS.n386 CS_BIAS.n385 24.5923
R17434 CS_BIAS.n391 CS_BIAS.n349 24.5923
R17435 CS_BIAS.n394 CS_BIAS.n393 24.5923
R17436 CS_BIAS.n399 CS_BIAS.n398 24.5923
R17437 CS_BIAS.n401 CS_BIAS.n345 24.5923
R17438 CS_BIAS.n406 CS_BIAS.n405 24.5923
R17439 CS_BIAS.n261 CS_BIAS.n260 24.5923
R17440 CS_BIAS.n266 CS_BIAS.n265 24.5923
R17441 CS_BIAS.n268 CS_BIAS.n254 24.5923
R17442 CS_BIAS.n275 CS_BIAS.n273 24.5923
R17443 CS_BIAS.n279 CS_BIAS.n252 24.5923
R17444 CS_BIAS.n281 CS_BIAS.n280 24.5923
R17445 CS_BIAS.n285 CS_BIAS.n284 24.5923
R17446 CS_BIAS.n290 CS_BIAS.n248 24.5923
R17447 CS_BIAS.n293 CS_BIAS.n292 24.5923
R17448 CS_BIAS.n298 CS_BIAS.n297 24.5923
R17449 CS_BIAS.n300 CS_BIAS.n244 24.5923
R17450 CS_BIAS.n305 CS_BIAS.n304 24.5923
R17451 CS_BIAS.n341 CS_BIAS.n340 24.5923
R17452 CS_BIAS.n334 CS_BIAS.n333 24.5923
R17453 CS_BIAS.n336 CS_BIAS.n206 24.5923
R17454 CS_BIAS.n326 CS_BIAS.n210 24.5923
R17455 CS_BIAS.n329 CS_BIAS.n328 24.5923
R17456 CS_BIAS.n317 CS_BIAS.n316 24.5923
R17457 CS_BIAS.n321 CS_BIAS.n320 24.5923
R17458 CS_BIAS.n223 CS_BIAS.n222 24.5923
R17459 CS_BIAS.n228 CS_BIAS.n227 24.5923
R17460 CS_BIAS.n230 CS_BIAS.n216 24.5923
R17461 CS_BIAS.n237 CS_BIAS.n235 24.5923
R17462 CS_BIAS.n315 CS_BIAS.n214 24.5923
R17463 CS_BIAS.n196 CS_BIAS.n195 20.9036
R17464 CS_BIAS.n67 CS_BIAS.n66 20.9036
R17465 CS_BIAS.n131 CS_BIAS.n130 20.9036
R17466 CS_BIAS.n401 CS_BIAS.n400 20.9036
R17467 CS_BIAS.n300 CS_BIAS.n299 20.9036
R17468 CS_BIAS.n336 CS_BIAS.n335 20.9036
R17469 CS_BIAS.n150 CS_BIAS.n148 20.4117
R17470 CS_BIAS.n177 CS_BIAS.n146 20.4117
R17471 CS_BIAS.n48 CS_BIAS.n17 20.4117
R17472 CS_BIAS.n21 CS_BIAS.n19 20.4117
R17473 CS_BIAS.n112 CS_BIAS.n7 20.4117
R17474 CS_BIAS.n85 CS_BIAS.n9 20.4117
R17475 CS_BIAS.n375 CS_BIAS.n353 20.4117
R17476 CS_BIAS.n382 CS_BIAS.n351 20.4117
R17477 CS_BIAS.n274 CS_BIAS.n252 20.4117
R17478 CS_BIAS.n281 CS_BIAS.n250 20.4117
R17479 CS_BIAS.n317 CS_BIAS.n212 20.4117
R17480 CS_BIAS.n236 CS_BIAS.n214 20.4117
R17481 CS_BIAS.n202 CS_BIAS.n201 19.9199
R17482 CS_BIAS.n73 CS_BIAS.n72 19.9199
R17483 CS_BIAS.n137 CS_BIAS.n136 19.9199
R17484 CS_BIAS.n407 CS_BIAS.n406 19.9199
R17485 CS_BIAS.n306 CS_BIAS.n305 19.9199
R17486 CS_BIAS.n342 CS_BIAS.n341 19.9199
R17487 CS_BIAS.n155 CS_BIAS.n154 13.3071
R17488 CS_BIAS.n359 CS_BIAS.n358 13.3071
R17489 CS_BIAS.n258 CS_BIAS.n257 13.3071
R17490 CS_BIAS.n220 CS_BIAS.n219 13.3071
R17491 CS_BIAS.n26 CS_BIAS.n25 13.3071
R17492 CS_BIAS.n90 CS_BIAS.n89 13.3071
R17493 CS_BIAS.n76 CS_BIAS.n74 13.0832
R17494 CS_BIAS.n309 CS_BIAS.n307 13.0832
R17495 CS_BIAS.n164 CS_BIAS.n163 12.5423
R17496 CS_BIAS.n188 CS_BIAS.n187 12.5423
R17497 CS_BIAS.n59 CS_BIAS.n58 12.5423
R17498 CS_BIAS.n35 CS_BIAS.n34 12.5423
R17499 CS_BIAS.n123 CS_BIAS.n122 12.5423
R17500 CS_BIAS.n99 CS_BIAS.n98 12.5423
R17501 CS_BIAS.n368 CS_BIAS.n367 12.5423
R17502 CS_BIAS.n393 CS_BIAS.n392 12.5423
R17503 CS_BIAS.n267 CS_BIAS.n266 12.5423
R17504 CS_BIAS.n292 CS_BIAS.n291 12.5423
R17505 CS_BIAS.n328 CS_BIAS.n327 12.5423
R17506 CS_BIAS.n229 CS_BIAS.n228 12.5423
R17507 CS_BIAS.n165 CS_BIAS.n164 12.0505
R17508 CS_BIAS.n187 CS_BIAS.n186 12.0505
R17509 CS_BIAS.n58 CS_BIAS.n57 12.0505
R17510 CS_BIAS.n36 CS_BIAS.n35 12.0505
R17511 CS_BIAS.n122 CS_BIAS.n121 12.0505
R17512 CS_BIAS.n100 CS_BIAS.n99 12.0505
R17513 CS_BIAS.n369 CS_BIAS.n368 12.0505
R17514 CS_BIAS.n392 CS_BIAS.n391 12.0505
R17515 CS_BIAS.n268 CS_BIAS.n267 12.0505
R17516 CS_BIAS.n291 CS_BIAS.n290 12.0505
R17517 CS_BIAS.n327 CS_BIAS.n326 12.0505
R17518 CS_BIAS.n230 CS_BIAS.n229 12.0505
R17519 CS_BIAS.n410 CS_BIAS.n204 11.7656
R17520 CS_BIAS.n410 CS_BIAS.n409 10.3158
R17521 CS_BIAS.n83 CS_BIAS.n82 9.50363
R17522 CS_BIAS.n313 CS_BIAS.n312 9.50363
R17523 CS_BIAS.n204 CS_BIAS.n138 8.35614
R17524 CS_BIAS.n409 CS_BIAS.n343 8.35614
R17525 CS_BIAS.n204 CS_BIAS.n203 5.04553
R17526 CS_BIAS.n409 CS_BIAS.n408 5.04553
R17527 CS_BIAS.n171 CS_BIAS.n150 4.18111
R17528 CS_BIAS.n180 CS_BIAS.n146 4.18111
R17529 CS_BIAS.n51 CS_BIAS.n17 4.18111
R17530 CS_BIAS.n42 CS_BIAS.n21 4.18111
R17531 CS_BIAS.n115 CS_BIAS.n7 4.18111
R17532 CS_BIAS.n106 CS_BIAS.n85 4.18111
R17533 CS_BIAS.n376 CS_BIAS.n375 4.18111
R17534 CS_BIAS.n385 CS_BIAS.n351 4.18111
R17535 CS_BIAS.n275 CS_BIAS.n274 4.18111
R17536 CS_BIAS.n284 CS_BIAS.n250 4.18111
R17537 CS_BIAS.n320 CS_BIAS.n212 4.18111
R17538 CS_BIAS.n237 CS_BIAS.n236 4.18111
R17539 CS_BIAS CS_BIAS.n410 3.99076
R17540 CS_BIAS.n157 CS_BIAS.n156 3.68928
R17541 CS_BIAS.n195 CS_BIAS.n194 3.68928
R17542 CS_BIAS.n66 CS_BIAS.n65 3.68928
R17543 CS_BIAS.n28 CS_BIAS.n27 3.68928
R17544 CS_BIAS.n130 CS_BIAS.n129 3.68928
R17545 CS_BIAS.n92 CS_BIAS.n91 3.68928
R17546 CS_BIAS.n361 CS_BIAS.n360 3.68928
R17547 CS_BIAS.n400 CS_BIAS.n399 3.68928
R17548 CS_BIAS.n260 CS_BIAS.n259 3.68928
R17549 CS_BIAS.n299 CS_BIAS.n298 3.68928
R17550 CS_BIAS.n335 CS_BIAS.n334 3.68928
R17551 CS_BIAS.n222 CS_BIAS.n221 3.68928
R17552 CS_BIAS.n79 CS_BIAS.t27 3.3005
R17553 CS_BIAS.n79 CS_BIAS.t15 3.3005
R17554 CS_BIAS.n80 CS_BIAS.t21 3.3005
R17555 CS_BIAS.n80 CS_BIAS.t1 3.3005
R17556 CS_BIAS.n77 CS_BIAS.t11 3.3005
R17557 CS_BIAS.n77 CS_BIAS.t3 3.3005
R17558 CS_BIAS.n75 CS_BIAS.t19 3.3005
R17559 CS_BIAS.n75 CS_BIAS.t25 3.3005
R17560 CS_BIAS.n308 CS_BIAS.t29 3.3005
R17561 CS_BIAS.n308 CS_BIAS.t17 3.3005
R17562 CS_BIAS.n310 CS_BIAS.t7 3.3005
R17563 CS_BIAS.n310 CS_BIAS.t9 3.3005
R17564 CS_BIAS.n241 CS_BIAS.t5 3.3005
R17565 CS_BIAS.n241 CS_BIAS.t23 3.3005
R17566 CS_BIAS.n240 CS_BIAS.t13 3.3005
R17567 CS_BIAS.n240 CS_BIAS.t31 3.3005
R17568 CS_BIAS.n78 CS_BIAS.n76 1.00481
R17569 CS_BIAS.n311 CS_BIAS.n309 1.00481
R17570 CS_BIAS.n82 CS_BIAS.n78 0.502655
R17571 CS_BIAS.n82 CS_BIAS.n81 0.502655
R17572 CS_BIAS.n312 CS_BIAS.n242 0.502655
R17573 CS_BIAS.n312 CS_BIAS.n311 0.502655
R17574 CS_BIAS.n203 CS_BIAS.n139 0.278335
R17575 CS_BIAS.n74 CS_BIAS.n10 0.278335
R17576 CS_BIAS.n138 CS_BIAS.n0 0.278335
R17577 CS_BIAS.n408 CS_BIAS.n344 0.278335
R17578 CS_BIAS.n307 CS_BIAS.n243 0.278335
R17579 CS_BIAS.n343 CS_BIAS.n205 0.278335
R17580 CS_BIAS.n199 CS_BIAS.n139 0.189894
R17581 CS_BIAS.n199 CS_BIAS.n198 0.189894
R17582 CS_BIAS.n198 CS_BIAS.n197 0.189894
R17583 CS_BIAS.n197 CS_BIAS.n141 0.189894
R17584 CS_BIAS.n192 CS_BIAS.n141 0.189894
R17585 CS_BIAS.n192 CS_BIAS.n191 0.189894
R17586 CS_BIAS.n191 CS_BIAS.n190 0.189894
R17587 CS_BIAS.n190 CS_BIAS.n143 0.189894
R17588 CS_BIAS.n185 CS_BIAS.n143 0.189894
R17589 CS_BIAS.n185 CS_BIAS.n184 0.189894
R17590 CS_BIAS.n184 CS_BIAS.n183 0.189894
R17591 CS_BIAS.n183 CS_BIAS.n145 0.189894
R17592 CS_BIAS.n179 CS_BIAS.n145 0.189894
R17593 CS_BIAS.n179 CS_BIAS.n178 0.189894
R17594 CS_BIAS.n178 CS_BIAS.n147 0.189894
R17595 CS_BIAS.n174 CS_BIAS.n147 0.189894
R17596 CS_BIAS.n174 CS_BIAS.n173 0.189894
R17597 CS_BIAS.n173 CS_BIAS.n172 0.189894
R17598 CS_BIAS.n172 CS_BIAS.n149 0.189894
R17599 CS_BIAS.n168 CS_BIAS.n149 0.189894
R17600 CS_BIAS.n168 CS_BIAS.n167 0.189894
R17601 CS_BIAS.n167 CS_BIAS.n166 0.189894
R17602 CS_BIAS.n166 CS_BIAS.n152 0.189894
R17603 CS_BIAS.n161 CS_BIAS.n152 0.189894
R17604 CS_BIAS.n161 CS_BIAS.n160 0.189894
R17605 CS_BIAS.n160 CS_BIAS.n159 0.189894
R17606 CS_BIAS.n159 CS_BIAS.n154 0.189894
R17607 CS_BIAS.n70 CS_BIAS.n10 0.189894
R17608 CS_BIAS.n70 CS_BIAS.n69 0.189894
R17609 CS_BIAS.n69 CS_BIAS.n68 0.189894
R17610 CS_BIAS.n68 CS_BIAS.n12 0.189894
R17611 CS_BIAS.n63 CS_BIAS.n12 0.189894
R17612 CS_BIAS.n63 CS_BIAS.n62 0.189894
R17613 CS_BIAS.n62 CS_BIAS.n61 0.189894
R17614 CS_BIAS.n61 CS_BIAS.n14 0.189894
R17615 CS_BIAS.n56 CS_BIAS.n14 0.189894
R17616 CS_BIAS.n56 CS_BIAS.n55 0.189894
R17617 CS_BIAS.n55 CS_BIAS.n54 0.189894
R17618 CS_BIAS.n54 CS_BIAS.n16 0.189894
R17619 CS_BIAS.n50 CS_BIAS.n16 0.189894
R17620 CS_BIAS.n50 CS_BIAS.n49 0.189894
R17621 CS_BIAS.n49 CS_BIAS.n18 0.189894
R17622 CS_BIAS.n45 CS_BIAS.n18 0.189894
R17623 CS_BIAS.n45 CS_BIAS.n44 0.189894
R17624 CS_BIAS.n44 CS_BIAS.n43 0.189894
R17625 CS_BIAS.n43 CS_BIAS.n20 0.189894
R17626 CS_BIAS.n39 CS_BIAS.n20 0.189894
R17627 CS_BIAS.n39 CS_BIAS.n38 0.189894
R17628 CS_BIAS.n38 CS_BIAS.n37 0.189894
R17629 CS_BIAS.n37 CS_BIAS.n23 0.189894
R17630 CS_BIAS.n32 CS_BIAS.n23 0.189894
R17631 CS_BIAS.n32 CS_BIAS.n31 0.189894
R17632 CS_BIAS.n31 CS_BIAS.n30 0.189894
R17633 CS_BIAS.n30 CS_BIAS.n25 0.189894
R17634 CS_BIAS.n109 CS_BIAS.n108 0.189894
R17635 CS_BIAS.n108 CS_BIAS.n107 0.189894
R17636 CS_BIAS.n107 CS_BIAS.n84 0.189894
R17637 CS_BIAS.n103 CS_BIAS.n84 0.189894
R17638 CS_BIAS.n103 CS_BIAS.n102 0.189894
R17639 CS_BIAS.n102 CS_BIAS.n101 0.189894
R17640 CS_BIAS.n101 CS_BIAS.n87 0.189894
R17641 CS_BIAS.n96 CS_BIAS.n87 0.189894
R17642 CS_BIAS.n96 CS_BIAS.n95 0.189894
R17643 CS_BIAS.n95 CS_BIAS.n94 0.189894
R17644 CS_BIAS.n94 CS_BIAS.n89 0.189894
R17645 CS_BIAS.n134 CS_BIAS.n0 0.189894
R17646 CS_BIAS.n134 CS_BIAS.n133 0.189894
R17647 CS_BIAS.n133 CS_BIAS.n132 0.189894
R17648 CS_BIAS.n132 CS_BIAS.n2 0.189894
R17649 CS_BIAS.n127 CS_BIAS.n2 0.189894
R17650 CS_BIAS.n127 CS_BIAS.n126 0.189894
R17651 CS_BIAS.n126 CS_BIAS.n125 0.189894
R17652 CS_BIAS.n125 CS_BIAS.n4 0.189894
R17653 CS_BIAS.n120 CS_BIAS.n4 0.189894
R17654 CS_BIAS.n120 CS_BIAS.n119 0.189894
R17655 CS_BIAS.n119 CS_BIAS.n118 0.189894
R17656 CS_BIAS.n118 CS_BIAS.n6 0.189894
R17657 CS_BIAS.n114 CS_BIAS.n6 0.189894
R17658 CS_BIAS.n114 CS_BIAS.n113 0.189894
R17659 CS_BIAS.n113 CS_BIAS.n8 0.189894
R17660 CS_BIAS.n363 CS_BIAS.n358 0.189894
R17661 CS_BIAS.n364 CS_BIAS.n363 0.189894
R17662 CS_BIAS.n365 CS_BIAS.n364 0.189894
R17663 CS_BIAS.n365 CS_BIAS.n356 0.189894
R17664 CS_BIAS.n370 CS_BIAS.n356 0.189894
R17665 CS_BIAS.n371 CS_BIAS.n370 0.189894
R17666 CS_BIAS.n372 CS_BIAS.n371 0.189894
R17667 CS_BIAS.n372 CS_BIAS.n354 0.189894
R17668 CS_BIAS.n377 CS_BIAS.n354 0.189894
R17669 CS_BIAS.n378 CS_BIAS.n377 0.189894
R17670 CS_BIAS.n379 CS_BIAS.n378 0.189894
R17671 CS_BIAS.n379 CS_BIAS.n352 0.189894
R17672 CS_BIAS.n383 CS_BIAS.n352 0.189894
R17673 CS_BIAS.n384 CS_BIAS.n383 0.189894
R17674 CS_BIAS.n384 CS_BIAS.n350 0.189894
R17675 CS_BIAS.n388 CS_BIAS.n350 0.189894
R17676 CS_BIAS.n389 CS_BIAS.n388 0.189894
R17677 CS_BIAS.n390 CS_BIAS.n389 0.189894
R17678 CS_BIAS.n390 CS_BIAS.n348 0.189894
R17679 CS_BIAS.n395 CS_BIAS.n348 0.189894
R17680 CS_BIAS.n396 CS_BIAS.n395 0.189894
R17681 CS_BIAS.n397 CS_BIAS.n396 0.189894
R17682 CS_BIAS.n397 CS_BIAS.n346 0.189894
R17683 CS_BIAS.n402 CS_BIAS.n346 0.189894
R17684 CS_BIAS.n403 CS_BIAS.n402 0.189894
R17685 CS_BIAS.n404 CS_BIAS.n403 0.189894
R17686 CS_BIAS.n404 CS_BIAS.n344 0.189894
R17687 CS_BIAS.n262 CS_BIAS.n257 0.189894
R17688 CS_BIAS.n263 CS_BIAS.n262 0.189894
R17689 CS_BIAS.n264 CS_BIAS.n263 0.189894
R17690 CS_BIAS.n264 CS_BIAS.n255 0.189894
R17691 CS_BIAS.n269 CS_BIAS.n255 0.189894
R17692 CS_BIAS.n270 CS_BIAS.n269 0.189894
R17693 CS_BIAS.n271 CS_BIAS.n270 0.189894
R17694 CS_BIAS.n271 CS_BIAS.n253 0.189894
R17695 CS_BIAS.n276 CS_BIAS.n253 0.189894
R17696 CS_BIAS.n277 CS_BIAS.n276 0.189894
R17697 CS_BIAS.n278 CS_BIAS.n277 0.189894
R17698 CS_BIAS.n278 CS_BIAS.n251 0.189894
R17699 CS_BIAS.n282 CS_BIAS.n251 0.189894
R17700 CS_BIAS.n283 CS_BIAS.n282 0.189894
R17701 CS_BIAS.n283 CS_BIAS.n249 0.189894
R17702 CS_BIAS.n287 CS_BIAS.n249 0.189894
R17703 CS_BIAS.n288 CS_BIAS.n287 0.189894
R17704 CS_BIAS.n289 CS_BIAS.n288 0.189894
R17705 CS_BIAS.n289 CS_BIAS.n247 0.189894
R17706 CS_BIAS.n294 CS_BIAS.n247 0.189894
R17707 CS_BIAS.n295 CS_BIAS.n294 0.189894
R17708 CS_BIAS.n296 CS_BIAS.n295 0.189894
R17709 CS_BIAS.n296 CS_BIAS.n245 0.189894
R17710 CS_BIAS.n301 CS_BIAS.n245 0.189894
R17711 CS_BIAS.n302 CS_BIAS.n301 0.189894
R17712 CS_BIAS.n303 CS_BIAS.n302 0.189894
R17713 CS_BIAS.n303 CS_BIAS.n243 0.189894
R17714 CS_BIAS.n224 CS_BIAS.n219 0.189894
R17715 CS_BIAS.n225 CS_BIAS.n224 0.189894
R17716 CS_BIAS.n226 CS_BIAS.n225 0.189894
R17717 CS_BIAS.n226 CS_BIAS.n217 0.189894
R17718 CS_BIAS.n231 CS_BIAS.n217 0.189894
R17719 CS_BIAS.n232 CS_BIAS.n231 0.189894
R17720 CS_BIAS.n233 CS_BIAS.n232 0.189894
R17721 CS_BIAS.n233 CS_BIAS.n215 0.189894
R17722 CS_BIAS.n238 CS_BIAS.n215 0.189894
R17723 CS_BIAS.n239 CS_BIAS.n238 0.189894
R17724 CS_BIAS.n314 CS_BIAS.n239 0.189894
R17725 CS_BIAS.n318 CS_BIAS.n213 0.189894
R17726 CS_BIAS.n319 CS_BIAS.n318 0.189894
R17727 CS_BIAS.n319 CS_BIAS.n211 0.189894
R17728 CS_BIAS.n323 CS_BIAS.n211 0.189894
R17729 CS_BIAS.n324 CS_BIAS.n323 0.189894
R17730 CS_BIAS.n325 CS_BIAS.n324 0.189894
R17731 CS_BIAS.n325 CS_BIAS.n209 0.189894
R17732 CS_BIAS.n330 CS_BIAS.n209 0.189894
R17733 CS_BIAS.n331 CS_BIAS.n330 0.189894
R17734 CS_BIAS.n332 CS_BIAS.n331 0.189894
R17735 CS_BIAS.n332 CS_BIAS.n207 0.189894
R17736 CS_BIAS.n337 CS_BIAS.n207 0.189894
R17737 CS_BIAS.n338 CS_BIAS.n337 0.189894
R17738 CS_BIAS.n339 CS_BIAS.n338 0.189894
R17739 CS_BIAS.n339 CS_BIAS.n205 0.189894
R17740 CS_BIAS.n109 CS_BIAS.n83 0.0762576
R17741 CS_BIAS.n83 CS_BIAS.n8 0.0762576
R17742 CS_BIAS.n314 CS_BIAS.n313 0.0762576
R17743 CS_BIAS.n313 CS_BIAS.n213 0.0762576
R17744 VN.n28 VN.t4 243.97
R17745 VN.n28 VN.n27 223.454
R17746 VN.n30 VN.n29 223.454
R17747 VN.n15 VN.t12 223.244
R17748 VN.n2 VN.t10 223.244
R17749 VN.n24 VN.t7 207.983
R17750 VN.n11 VN.t6 207.983
R17751 VN.n16 VN.t11 168.701
R17752 VN.n22 VN.t8 168.701
R17753 VN.n9 VN.t5 168.701
R17754 VN.n3 VN.t9 168.701
R17755 VN.n23 VN.n13 161.3
R17756 VN.n21 VN.n20 161.3
R17757 VN.n19 VN.n14 161.3
R17758 VN.n18 VN.n17 161.3
R17759 VN.n5 VN.n4 161.3
R17760 VN.n6 VN.n1 161.3
R17761 VN.n8 VN.n7 161.3
R17762 VN.n10 VN.n0 161.3
R17763 VN.n25 VN.n24 80.6037
R17764 VN.n12 VN.n11 80.6037
R17765 VN.n24 VN.n23 56.3158
R17766 VN.n11 VN.n10 56.3158
R17767 VN.n16 VN.n15 46.9082
R17768 VN.n3 VN.n2 46.9082
R17769 VN.n18 VN.n15 43.8991
R17770 VN.n5 VN.n2 43.8991
R17771 VN.n17 VN.n14 40.577
R17772 VN.n21 VN.n14 40.577
R17773 VN.n8 VN.n1 40.577
R17774 VN.n4 VN.n1 40.577
R17775 VN.n26 VN.n25 28.2718
R17776 VN.n27 VN.t0 19.8005
R17777 VN.n27 VN.t3 19.8005
R17778 VN.n29 VN.t1 19.8005
R17779 VN.n29 VN.t2 19.8005
R17780 VN.n23 VN.n22 16.477
R17781 VN.n10 VN.n9 16.477
R17782 VN VN.n31 13.8471
R17783 VN.n26 VN.n12 12.0786
R17784 VN.n17 VN.n16 8.11581
R17785 VN.n22 VN.n21 8.11581
R17786 VN.n9 VN.n8 8.11581
R17787 VN.n4 VN.n3 8.11581
R17788 VN.n31 VN.n30 5.40567
R17789 VN.n31 VN.n26 1.188
R17790 VN.n30 VN.n28 0.716017
R17791 VN.n25 VN.n13 0.285035
R17792 VN.n12 VN.n0 0.285035
R17793 VN.n19 VN.n18 0.189894
R17794 VN.n20 VN.n19 0.189894
R17795 VN.n20 VN.n13 0.189894
R17796 VN.n7 VN.n0 0.189894
R17797 VN.n7 VN.n6 0.189894
R17798 VN.n6 VN.n5 0.189894
R17799 a_n2511_10556.n130 a_n2511_10556.n104 756.745
R17800 a_n2511_10556.n96 a_n2511_10556.n70 756.745
R17801 a_n2511_10556.n64 a_n2511_10556.n38 756.745
R17802 a_n2511_10556.n31 a_n2511_10556.n5 756.745
R17803 a_n2511_10556.n131 a_n2511_10556.n130 585
R17804 a_n2511_10556.n129 a_n2511_10556.n128 585
R17805 a_n2511_10556.n108 a_n2511_10556.n107 585
R17806 a_n2511_10556.n123 a_n2511_10556.n122 585
R17807 a_n2511_10556.n121 a_n2511_10556.n120 585
R17808 a_n2511_10556.n112 a_n2511_10556.n111 585
R17809 a_n2511_10556.n115 a_n2511_10556.n114 585
R17810 a_n2511_10556.n97 a_n2511_10556.n96 585
R17811 a_n2511_10556.n95 a_n2511_10556.n94 585
R17812 a_n2511_10556.n74 a_n2511_10556.n73 585
R17813 a_n2511_10556.n89 a_n2511_10556.n88 585
R17814 a_n2511_10556.n87 a_n2511_10556.n86 585
R17815 a_n2511_10556.n78 a_n2511_10556.n77 585
R17816 a_n2511_10556.n81 a_n2511_10556.n80 585
R17817 a_n2511_10556.n65 a_n2511_10556.n64 585
R17818 a_n2511_10556.n63 a_n2511_10556.n62 585
R17819 a_n2511_10556.n42 a_n2511_10556.n41 585
R17820 a_n2511_10556.n57 a_n2511_10556.n56 585
R17821 a_n2511_10556.n55 a_n2511_10556.n54 585
R17822 a_n2511_10556.n46 a_n2511_10556.n45 585
R17823 a_n2511_10556.n49 a_n2511_10556.n48 585
R17824 a_n2511_10556.n32 a_n2511_10556.n31 585
R17825 a_n2511_10556.n30 a_n2511_10556.n29 585
R17826 a_n2511_10556.n9 a_n2511_10556.n8 585
R17827 a_n2511_10556.n24 a_n2511_10556.n23 585
R17828 a_n2511_10556.n22 a_n2511_10556.n21 585
R17829 a_n2511_10556.n13 a_n2511_10556.n12 585
R17830 a_n2511_10556.n16 a_n2511_10556.n15 585
R17831 a_n2511_10556.t17 a_n2511_10556.n113 327.601
R17832 a_n2511_10556.t14 a_n2511_10556.n79 327.601
R17833 a_n2511_10556.t19 a_n2511_10556.n47 327.601
R17834 a_n2511_10556.t16 a_n2511_10556.n14 327.601
R17835 a_n2511_10556.n130 a_n2511_10556.n129 171.744
R17836 a_n2511_10556.n129 a_n2511_10556.n107 171.744
R17837 a_n2511_10556.n122 a_n2511_10556.n107 171.744
R17838 a_n2511_10556.n122 a_n2511_10556.n121 171.744
R17839 a_n2511_10556.n121 a_n2511_10556.n111 171.744
R17840 a_n2511_10556.n114 a_n2511_10556.n111 171.744
R17841 a_n2511_10556.n96 a_n2511_10556.n95 171.744
R17842 a_n2511_10556.n95 a_n2511_10556.n73 171.744
R17843 a_n2511_10556.n88 a_n2511_10556.n73 171.744
R17844 a_n2511_10556.n88 a_n2511_10556.n87 171.744
R17845 a_n2511_10556.n87 a_n2511_10556.n77 171.744
R17846 a_n2511_10556.n80 a_n2511_10556.n77 171.744
R17847 a_n2511_10556.n64 a_n2511_10556.n63 171.744
R17848 a_n2511_10556.n63 a_n2511_10556.n41 171.744
R17849 a_n2511_10556.n56 a_n2511_10556.n41 171.744
R17850 a_n2511_10556.n56 a_n2511_10556.n55 171.744
R17851 a_n2511_10556.n55 a_n2511_10556.n45 171.744
R17852 a_n2511_10556.n48 a_n2511_10556.n45 171.744
R17853 a_n2511_10556.n31 a_n2511_10556.n30 171.744
R17854 a_n2511_10556.n30 a_n2511_10556.n8 171.744
R17855 a_n2511_10556.n23 a_n2511_10556.n8 171.744
R17856 a_n2511_10556.n23 a_n2511_10556.n22 171.744
R17857 a_n2511_10556.n22 a_n2511_10556.n12 171.744
R17858 a_n2511_10556.n15 a_n2511_10556.n12 171.744
R17859 a_n2511_10556.n141 a_n2511_10556.n140 109.74
R17860 a_n2511_10556.n2 a_n2511_10556.n0 109.401
R17861 a_n2511_10556.n140 a_n2511_10556.n139 109.166
R17862 a_n2511_10556.n4 a_n2511_10556.n3 109.166
R17863 a_n2511_10556.n2 a_n2511_10556.n1 109.166
R17864 a_n2511_10556.n138 a_n2511_10556.n137 109.166
R17865 a_n2511_10556.n114 a_n2511_10556.t17 85.8723
R17866 a_n2511_10556.n80 a_n2511_10556.t14 85.8723
R17867 a_n2511_10556.n48 a_n2511_10556.t19 85.8723
R17868 a_n2511_10556.n15 a_n2511_10556.t16 85.8723
R17869 a_n2511_10556.n103 a_n2511_10556.n102 81.2397
R17870 a_n2511_10556.n37 a_n2511_10556.n36 81.2397
R17871 a_n2511_10556.n37 a_n2511_10556.n35 38.3829
R17872 a_n2511_10556.n135 a_n2511_10556.n134 37.8096
R17873 a_n2511_10556.n101 a_n2511_10556.n100 37.8096
R17874 a_n2511_10556.n69 a_n2511_10556.n68 37.8096
R17875 a_n2511_10556.n115 a_n2511_10556.n113 16.3865
R17876 a_n2511_10556.n81 a_n2511_10556.n79 16.3865
R17877 a_n2511_10556.n49 a_n2511_10556.n47 16.3865
R17878 a_n2511_10556.n16 a_n2511_10556.n14 16.3865
R17879 a_n2511_10556.n136 a_n2511_10556.n4 13.2313
R17880 a_n2511_10556.n116 a_n2511_10556.n112 12.8005
R17881 a_n2511_10556.n82 a_n2511_10556.n78 12.8005
R17882 a_n2511_10556.n50 a_n2511_10556.n46 12.8005
R17883 a_n2511_10556.n17 a_n2511_10556.n13 12.8005
R17884 a_n2511_10556.n120 a_n2511_10556.n119 12.0247
R17885 a_n2511_10556.n86 a_n2511_10556.n85 12.0247
R17886 a_n2511_10556.n54 a_n2511_10556.n53 12.0247
R17887 a_n2511_10556.n21 a_n2511_10556.n20 12.0247
R17888 a_n2511_10556.n123 a_n2511_10556.n110 11.249
R17889 a_n2511_10556.n89 a_n2511_10556.n76 11.249
R17890 a_n2511_10556.n57 a_n2511_10556.n44 11.249
R17891 a_n2511_10556.n24 a_n2511_10556.n11 11.249
R17892 a_n2511_10556.n124 a_n2511_10556.n108 10.4732
R17893 a_n2511_10556.n90 a_n2511_10556.n74 10.4732
R17894 a_n2511_10556.n58 a_n2511_10556.n42 10.4732
R17895 a_n2511_10556.n25 a_n2511_10556.n9 10.4732
R17896 a_n2511_10556.n138 a_n2511_10556.n136 10.4398
R17897 a_n2511_10556.n128 a_n2511_10556.n127 9.69747
R17898 a_n2511_10556.n94 a_n2511_10556.n93 9.69747
R17899 a_n2511_10556.n62 a_n2511_10556.n61 9.69747
R17900 a_n2511_10556.n29 a_n2511_10556.n28 9.69747
R17901 a_n2511_10556.n134 a_n2511_10556.n133 9.45567
R17902 a_n2511_10556.n100 a_n2511_10556.n99 9.45567
R17903 a_n2511_10556.n68 a_n2511_10556.n67 9.45567
R17904 a_n2511_10556.n35 a_n2511_10556.n34 9.45567
R17905 a_n2511_10556.n133 a_n2511_10556.n132 9.3005
R17906 a_n2511_10556.n106 a_n2511_10556.n105 9.3005
R17907 a_n2511_10556.n127 a_n2511_10556.n126 9.3005
R17908 a_n2511_10556.n125 a_n2511_10556.n124 9.3005
R17909 a_n2511_10556.n110 a_n2511_10556.n109 9.3005
R17910 a_n2511_10556.n119 a_n2511_10556.n118 9.3005
R17911 a_n2511_10556.n117 a_n2511_10556.n116 9.3005
R17912 a_n2511_10556.n99 a_n2511_10556.n98 9.3005
R17913 a_n2511_10556.n72 a_n2511_10556.n71 9.3005
R17914 a_n2511_10556.n93 a_n2511_10556.n92 9.3005
R17915 a_n2511_10556.n91 a_n2511_10556.n90 9.3005
R17916 a_n2511_10556.n76 a_n2511_10556.n75 9.3005
R17917 a_n2511_10556.n85 a_n2511_10556.n84 9.3005
R17918 a_n2511_10556.n83 a_n2511_10556.n82 9.3005
R17919 a_n2511_10556.n67 a_n2511_10556.n66 9.3005
R17920 a_n2511_10556.n40 a_n2511_10556.n39 9.3005
R17921 a_n2511_10556.n61 a_n2511_10556.n60 9.3005
R17922 a_n2511_10556.n59 a_n2511_10556.n58 9.3005
R17923 a_n2511_10556.n44 a_n2511_10556.n43 9.3005
R17924 a_n2511_10556.n53 a_n2511_10556.n52 9.3005
R17925 a_n2511_10556.n51 a_n2511_10556.n50 9.3005
R17926 a_n2511_10556.n34 a_n2511_10556.n33 9.3005
R17927 a_n2511_10556.n7 a_n2511_10556.n6 9.3005
R17928 a_n2511_10556.n28 a_n2511_10556.n27 9.3005
R17929 a_n2511_10556.n26 a_n2511_10556.n25 9.3005
R17930 a_n2511_10556.n11 a_n2511_10556.n10 9.3005
R17931 a_n2511_10556.n20 a_n2511_10556.n19 9.3005
R17932 a_n2511_10556.n18 a_n2511_10556.n17 9.3005
R17933 a_n2511_10556.n131 a_n2511_10556.n106 8.92171
R17934 a_n2511_10556.n97 a_n2511_10556.n72 8.92171
R17935 a_n2511_10556.n65 a_n2511_10556.n40 8.92171
R17936 a_n2511_10556.n32 a_n2511_10556.n7 8.92171
R17937 a_n2511_10556.n132 a_n2511_10556.n104 8.14595
R17938 a_n2511_10556.n98 a_n2511_10556.n70 8.14595
R17939 a_n2511_10556.n66 a_n2511_10556.n38 8.14595
R17940 a_n2511_10556.n33 a_n2511_10556.n5 8.14595
R17941 a_n2511_10556.n136 a_n2511_10556.n135 5.91753
R17942 a_n2511_10556.n134 a_n2511_10556.n104 5.81868
R17943 a_n2511_10556.n100 a_n2511_10556.n70 5.81868
R17944 a_n2511_10556.n68 a_n2511_10556.n38 5.81868
R17945 a_n2511_10556.n35 a_n2511_10556.n5 5.81868
R17946 a_n2511_10556.n137 a_n2511_10556.t2 5.418
R17947 a_n2511_10556.n137 a_n2511_10556.t4 5.418
R17948 a_n2511_10556.n139 a_n2511_10556.t0 5.418
R17949 a_n2511_10556.n139 a_n2511_10556.t10 5.418
R17950 a_n2511_10556.n102 a_n2511_10556.t18 5.418
R17951 a_n2511_10556.n102 a_n2511_10556.t12 5.418
R17952 a_n2511_10556.n36 a_n2511_10556.t13 5.418
R17953 a_n2511_10556.n36 a_n2511_10556.t15 5.418
R17954 a_n2511_10556.n3 a_n2511_10556.t5 5.418
R17955 a_n2511_10556.n3 a_n2511_10556.t9 5.418
R17956 a_n2511_10556.n1 a_n2511_10556.t1 5.418
R17957 a_n2511_10556.n1 a_n2511_10556.t3 5.418
R17958 a_n2511_10556.n0 a_n2511_10556.t7 5.418
R17959 a_n2511_10556.n0 a_n2511_10556.t6 5.418
R17960 a_n2511_10556.n141 a_n2511_10556.t8 5.418
R17961 a_n2511_10556.t11 a_n2511_10556.n141 5.418
R17962 a_n2511_10556.n132 a_n2511_10556.n131 5.04292
R17963 a_n2511_10556.n98 a_n2511_10556.n97 5.04292
R17964 a_n2511_10556.n66 a_n2511_10556.n65 5.04292
R17965 a_n2511_10556.n33 a_n2511_10556.n32 5.04292
R17966 a_n2511_10556.n128 a_n2511_10556.n106 4.26717
R17967 a_n2511_10556.n94 a_n2511_10556.n72 4.26717
R17968 a_n2511_10556.n62 a_n2511_10556.n40 4.26717
R17969 a_n2511_10556.n29 a_n2511_10556.n7 4.26717
R17970 a_n2511_10556.n117 a_n2511_10556.n113 3.71286
R17971 a_n2511_10556.n83 a_n2511_10556.n79 3.71286
R17972 a_n2511_10556.n51 a_n2511_10556.n47 3.71286
R17973 a_n2511_10556.n18 a_n2511_10556.n14 3.71286
R17974 a_n2511_10556.n127 a_n2511_10556.n108 3.49141
R17975 a_n2511_10556.n93 a_n2511_10556.n74 3.49141
R17976 a_n2511_10556.n61 a_n2511_10556.n42 3.49141
R17977 a_n2511_10556.n28 a_n2511_10556.n9 3.49141
R17978 a_n2511_10556.n124 a_n2511_10556.n123 2.71565
R17979 a_n2511_10556.n90 a_n2511_10556.n89 2.71565
R17980 a_n2511_10556.n58 a_n2511_10556.n57 2.71565
R17981 a_n2511_10556.n25 a_n2511_10556.n24 2.71565
R17982 a_n2511_10556.n120 a_n2511_10556.n110 1.93989
R17983 a_n2511_10556.n86 a_n2511_10556.n76 1.93989
R17984 a_n2511_10556.n54 a_n2511_10556.n44 1.93989
R17985 a_n2511_10556.n21 a_n2511_10556.n11 1.93989
R17986 a_n2511_10556.n119 a_n2511_10556.n112 1.16414
R17987 a_n2511_10556.n85 a_n2511_10556.n78 1.16414
R17988 a_n2511_10556.n53 a_n2511_10556.n46 1.16414
R17989 a_n2511_10556.n20 a_n2511_10556.n13 1.16414
R17990 a_n2511_10556.n69 a_n2511_10556.n37 0.573776
R17991 a_n2511_10556.n103 a_n2511_10556.n101 0.573776
R17992 a_n2511_10556.n135 a_n2511_10556.n103 0.573776
R17993 a_n2511_10556.n140 a_n2511_10556.n138 0.573776
R17994 a_n2511_10556.n116 a_n2511_10556.n115 0.388379
R17995 a_n2511_10556.n82 a_n2511_10556.n81 0.388379
R17996 a_n2511_10556.n50 a_n2511_10556.n49 0.388379
R17997 a_n2511_10556.n17 a_n2511_10556.n16 0.388379
R17998 a_n2511_10556.n4 a_n2511_10556.n2 0.234655
R17999 a_n2511_10556.n133 a_n2511_10556.n105 0.155672
R18000 a_n2511_10556.n126 a_n2511_10556.n105 0.155672
R18001 a_n2511_10556.n126 a_n2511_10556.n125 0.155672
R18002 a_n2511_10556.n125 a_n2511_10556.n109 0.155672
R18003 a_n2511_10556.n118 a_n2511_10556.n109 0.155672
R18004 a_n2511_10556.n118 a_n2511_10556.n117 0.155672
R18005 a_n2511_10556.n99 a_n2511_10556.n71 0.155672
R18006 a_n2511_10556.n92 a_n2511_10556.n71 0.155672
R18007 a_n2511_10556.n92 a_n2511_10556.n91 0.155672
R18008 a_n2511_10556.n91 a_n2511_10556.n75 0.155672
R18009 a_n2511_10556.n84 a_n2511_10556.n75 0.155672
R18010 a_n2511_10556.n84 a_n2511_10556.n83 0.155672
R18011 a_n2511_10556.n67 a_n2511_10556.n39 0.155672
R18012 a_n2511_10556.n60 a_n2511_10556.n39 0.155672
R18013 a_n2511_10556.n60 a_n2511_10556.n59 0.155672
R18014 a_n2511_10556.n59 a_n2511_10556.n43 0.155672
R18015 a_n2511_10556.n52 a_n2511_10556.n43 0.155672
R18016 a_n2511_10556.n52 a_n2511_10556.n51 0.155672
R18017 a_n2511_10556.n34 a_n2511_10556.n6 0.155672
R18018 a_n2511_10556.n27 a_n2511_10556.n6 0.155672
R18019 a_n2511_10556.n27 a_n2511_10556.n26 0.155672
R18020 a_n2511_10556.n26 a_n2511_10556.n10 0.155672
R18021 a_n2511_10556.n19 a_n2511_10556.n10 0.155672
R18022 a_n2511_10556.n19 a_n2511_10556.n18 0.155672
R18023 a_n2511_10556.n101 a_n2511_10556.n69 0.155672
R18024 a_n1455_n3928.n10 a_n1455_n3928.t1 214.862
R18025 a_n1455_n3928.n13 a_n1455_n3928.t2 214.321
R18026 a_n1455_n3928.n12 a_n1455_n3928.t6 214.321
R18027 a_n1455_n3928.n11 a_n1455_n3928.t7 214.321
R18028 a_n1455_n3928.n4 a_n1455_n3928.t8 55.8337
R18029 a_n1455_n3928.n5 a_n1455_n3928.t17 55.8337
R18030 a_n1455_n3928.n8 a_n1455_n3928.t4 55.8337
R18031 a_n1455_n3928.n1 a_n1455_n3928.t13 55.8335
R18032 a_n1455_n3928.n15 a_n1455_n3928.t18 55.8335
R18033 a_n1455_n3928.n18 a_n1455_n3928.t19 55.8335
R18034 a_n1455_n3928.n19 a_n1455_n3928.t10 55.8335
R18035 a_n1455_n3928.n0 a_n1455_n3928.t14 55.8335
R18036 a_n1455_n3928.n21 a_n1455_n3928.n20 53.0054
R18037 a_n1455_n3928.n3 a_n1455_n3928.n2 53.0052
R18038 a_n1455_n3928.n7 a_n1455_n3928.n6 53.0052
R18039 a_n1455_n3928.n17 a_n1455_n3928.n16 53.0051
R18040 a_n1455_n3928.n9 a_n1455_n3928.n8 12.2632
R18041 a_n1455_n3928.n14 a_n1455_n3928.n1 12.2632
R18042 a_n1455_n3928.n9 a_n1455_n3928.n0 5.18369
R18043 a_n1455_n3928.n15 a_n1455_n3928.n14 5.18369
R18044 a_n1455_n3928.n16 a_n1455_n3928.t3 2.82907
R18045 a_n1455_n3928.n16 a_n1455_n3928.t16 2.82907
R18046 a_n1455_n3928.n2 a_n1455_n3928.t9 2.82907
R18047 a_n1455_n3928.n2 a_n1455_n3928.t12 2.82907
R18048 a_n1455_n3928.n6 a_n1455_n3928.t5 2.82907
R18049 a_n1455_n3928.n6 a_n1455_n3928.t0 2.82907
R18050 a_n1455_n3928.t15 a_n1455_n3928.n21 2.82907
R18051 a_n1455_n3928.n21 a_n1455_n3928.t11 2.82907
R18052 a_n1455_n3928.n14 a_n1455_n3928.n13 2.23674
R18053 a_n1455_n3928.n10 a_n1455_n3928.n9 1.95694
R18054 a_n1455_n3928.n12 a_n1455_n3928.n11 0.962709
R18055 a_n1455_n3928.n13 a_n1455_n3928.n12 0.962709
R18056 a_n1455_n3928.n8 a_n1455_n3928.n7 0.573776
R18057 a_n1455_n3928.n7 a_n1455_n3928.n5 0.573776
R18058 a_n1455_n3928.n4 a_n1455_n3928.n3 0.573776
R18059 a_n1455_n3928.n3 a_n1455_n3928.n1 0.573776
R18060 a_n1455_n3928.n20 a_n1455_n3928.n0 0.573776
R18061 a_n1455_n3928.n20 a_n1455_n3928.n19 0.573776
R18062 a_n1455_n3928.n18 a_n1455_n3928.n17 0.573776
R18063 a_n1455_n3928.n17 a_n1455_n3928.n15 0.573776
R18064 a_n1455_n3928.n11 a_n1455_n3928.n10 0.422738
R18065 a_n1455_n3928.n5 a_n1455_n3928.n4 0.235414
R18066 a_n1455_n3928.n19 a_n1455_n3928.n18 0.235414
R18067 VP.n30 VP.t2 243.255
R18068 VP.n29 VP.n27 224.169
R18069 VP.n29 VP.n28 223.454
R18070 VP.n15 VP.t6 223.244
R18071 VP.n2 VP.t8 223.244
R18072 VP.n24 VP.t12 207.983
R18073 VP.n11 VP.t10 207.983
R18074 VP.n22 VP.t9 168.701
R18075 VP.n16 VP.t5 168.701
R18076 VP.n3 VP.t7 168.701
R18077 VP.n9 VP.t11 168.701
R18078 VP.n18 VP.n17 161.3
R18079 VP.n19 VP.n14 161.3
R18080 VP.n21 VP.n20 161.3
R18081 VP.n23 VP.n13 161.3
R18082 VP.n10 VP.n0 161.3
R18083 VP.n8 VP.n7 161.3
R18084 VP.n6 VP.n1 161.3
R18085 VP.n5 VP.n4 161.3
R18086 VP.n25 VP.n24 80.6037
R18087 VP.n12 VP.n11 80.6037
R18088 VP.n24 VP.n23 56.3158
R18089 VP.n11 VP.n10 56.3158
R18090 VP.n16 VP.n15 46.9082
R18091 VP.n3 VP.n2 46.9082
R18092 VP.n5 VP.n2 43.8991
R18093 VP.n18 VP.n15 43.8991
R18094 VP.n21 VP.n14 40.577
R18095 VP.n17 VP.n14 40.577
R18096 VP.n4 VP.n1 40.577
R18097 VP.n8 VP.n1 40.577
R18098 VP.n26 VP.n25 28.4877
R18099 VP.n28 VP.t4 19.8005
R18100 VP.n28 VP.t1 19.8005
R18101 VP.n27 VP.t3 19.8005
R18102 VP.n27 VP.t0 19.8005
R18103 VP.n23 VP.n22 16.477
R18104 VP.n10 VP.n9 16.477
R18105 VP.n26 VP.n12 12.2945
R18106 VP VP.n31 11.5274
R18107 VP.n22 VP.n21 8.11581
R18108 VP.n17 VP.n16 8.11581
R18109 VP.n4 VP.n3 8.11581
R18110 VP.n9 VP.n8 8.11581
R18111 VP.n31 VP.n30 4.80222
R18112 VP.n31 VP.n26 0.972091
R18113 VP.n30 VP.n29 0.716017
R18114 VP.n25 VP.n13 0.285035
R18115 VP.n12 VP.n0 0.285035
R18116 VP.n20 VP.n13 0.189894
R18117 VP.n20 VP.n19 0.189894
R18118 VP.n19 VP.n18 0.189894
R18119 VP.n6 VP.n5 0.189894
R18120 VP.n7 VP.n6 0.189894
R18121 VP.n7 VP.n0 0.189894
R18122 DIFFPAIR_BIAS.n0 DIFFPAIR_BIAS.t9 190.994
R18123 DIFFPAIR_BIAS.n9 DIFFPAIR_BIAS.t10 189.069
R18124 DIFFPAIR_BIAS.n8 DIFFPAIR_BIAS.t11 189.069
R18125 DIFFPAIR_BIAS.n0 DIFFPAIR_BIAS.t8 189.069
R18126 DIFFPAIR_BIAS.n4 DIFFPAIR_BIAS.t0 144.412
R18127 DIFFPAIR_BIAS.n4 DIFFPAIR_BIAS.t2 142.487
R18128 DIFFPAIR_BIAS.n5 DIFFPAIR_BIAS.t4 142.487
R18129 DIFFPAIR_BIAS.n6 DIFFPAIR_BIAS.t6 142.487
R18130 DIFFPAIR_BIAS.n1 DIFFPAIR_BIAS.t1 113.659
R18131 DIFFPAIR_BIAS.n1 DIFFPAIR_BIAS.t3 112.698
R18132 DIFFPAIR_BIAS.n2 DIFFPAIR_BIAS.t5 112.698
R18133 DIFFPAIR_BIAS.n3 DIFFPAIR_BIAS.t7 112.698
R18134 DIFFPAIR_BIAS.n7 DIFFPAIR_BIAS.n6 5.20947
R18135 DIFFPAIR_BIAS.n7 DIFFPAIR_BIAS.n3 4.45342
R18136 DIFFPAIR_BIAS.n8 DIFFPAIR_BIAS.n7 4.28454
R18137 DIFFPAIR_BIAS.n6 DIFFPAIR_BIAS.n5 1.9266
R18138 DIFFPAIR_BIAS.n5 DIFFPAIR_BIAS.n4 1.9266
R18139 DIFFPAIR_BIAS.n9 DIFFPAIR_BIAS.n8 1.92658
R18140 DIFFPAIR_BIAS.n10 DIFFPAIR_BIAS.n9 1.29913
R18141 DIFFPAIR_BIAS.n3 DIFFPAIR_BIAS.n2 0.962709
R18142 DIFFPAIR_BIAS.n2 DIFFPAIR_BIAS.n1 0.962709
R18143 DIFFPAIR_BIAS DIFFPAIR_BIAS.n10 0.684875
R18144 DIFFPAIR_BIAS.n10 DIFFPAIR_BIAS.n0 0.337251
C0 VDD VN 0.05139f
C1 VOUT VP 2.74686f
C2 VOUT VN 0.804612f
C3 VP VN 8.028561f
C4 VOUT CS_BIAS 23.0378f
C5 VP CS_BIAS 0.306594f
C6 VN CS_BIAS 0.266289f
C7 VP DIFFPAIR_BIAS 2.16e-19
C8 VN DIFFPAIR_BIAS 2.16e-19
C9 CS_BIAS DIFFPAIR_BIAS 0.007973f
C10 VDD VOUT 54.654396f
C11 DIFFPAIR_BIAS GND 34.027576f
C12 CS_BIAS GND 0.111625p
C13 VN GND 26.09265f
C14 VP GND 22.64322f
C15 VOUT GND 62.452892f
C16 VDD GND 0.331217p
C17 DIFFPAIR_BIAS.t8 GND 0.127601f
C18 DIFFPAIR_BIAS.t9 GND 0.128381f
C19 DIFFPAIR_BIAS.n0 GND 0.137143f
C20 DIFFPAIR_BIAS.t1 GND 0.064103f
C21 DIFFPAIR_BIAS.t3 GND 0.06357f
C22 DIFFPAIR_BIAS.n1 GND 0.131903f
C23 DIFFPAIR_BIAS.t5 GND 0.06357f
C24 DIFFPAIR_BIAS.n2 GND 0.069455f
C25 DIFFPAIR_BIAS.t7 GND 0.06357f
C26 DIFFPAIR_BIAS.n3 GND 0.090481f
C27 DIFFPAIR_BIAS.t6 GND 0.120364f
C28 DIFFPAIR_BIAS.t4 GND 0.120364f
C29 DIFFPAIR_BIAS.t2 GND 0.120364f
C30 DIFFPAIR_BIAS.t0 GND 0.121265f
C31 DIFFPAIR_BIAS.n4 GND 0.14338f
C32 DIFFPAIR_BIAS.n5 GND 0.076729f
C33 DIFFPAIR_BIAS.n6 GND 0.08402f
C34 DIFFPAIR_BIAS.n7 GND 0.175839f
C35 DIFFPAIR_BIAS.t11 GND 0.127601f
C36 DIFFPAIR_BIAS.n8 GND 0.070966f
C37 DIFFPAIR_BIAS.t10 GND 0.127601f
C38 DIFFPAIR_BIAS.n9 GND 0.068629f
C39 DIFFPAIR_BIAS.n10 GND 0.04192f
C40 VP.n0 GND 0.037789f
C41 VP.t11 GND 0.529101f
C42 VP.n1 GND 0.022873f
C43 VP.t8 GND 0.589662f
C44 VP.n2 GND 0.251725f
C45 VP.t7 GND 0.529101f
C46 VP.n3 GND 0.236311f
C47 VP.n4 GND 0.038618f
C48 VP.n5 GND 0.121236f
C49 VP.n6 GND 0.02832f
C50 VP.n7 GND 0.02832f
C51 VP.n8 GND 0.038618f
C52 VP.n9 GND 0.211111f
C53 VP.n10 GND 0.038845f
C54 VP.t10 GND 0.572222f
C55 VP.n11 GND 0.254921f
C56 VP.n12 GND 0.351282f
C57 VP.n13 GND 0.037789f
C58 VP.t12 GND 0.572222f
C59 VP.t9 GND 0.529101f
C60 VP.n14 GND 0.022873f
C61 VP.t6 GND 0.589662f
C62 VP.n15 GND 0.251724f
C63 VP.t5 GND 0.529101f
C64 VP.n16 GND 0.236311f
C65 VP.n17 GND 0.038618f
C66 VP.n18 GND 0.121236f
C67 VP.n19 GND 0.02832f
C68 VP.n20 GND 0.02832f
C69 VP.n21 GND 0.038618f
C70 VP.n22 GND 0.211111f
C71 VP.n23 GND 0.038845f
C72 VP.n24 GND 0.254921f
C73 VP.n25 GND 0.769337f
C74 VP.n26 GND 1.15622f
C75 VP.t3 GND 0.00873f
C76 VP.t0 GND 0.00873f
C77 VP.n27 GND 0.028707f
C78 VP.t4 GND 0.00873f
C79 VP.t1 GND 0.00873f
C80 VP.n28 GND 0.028313f
C81 VP.n29 GND 0.241641f
C82 VP.t2 GND 0.048591f
C83 VP.n30 GND 0.131861f
C84 VP.n31 GND 1.77136f
C85 a_n1455_n3928.t14 GND 0.848403f
C86 a_n1455_n3928.n0 GND 0.542321f
C87 a_n1455_n3928.t13 GND 0.848402f
C88 a_n1455_n3928.n1 GND 0.809655f
C89 a_n1455_n3928.t9 GND 0.081631f
C90 a_n1455_n3928.t12 GND 0.081631f
C91 a_n1455_n3928.n2 GND 0.666694f
C92 a_n1455_n3928.n3 GND 0.352373f
C93 a_n1455_n3928.t8 GND 0.848406f
C94 a_n1455_n3928.n4 GND 0.328934f
C95 a_n1455_n3928.t17 GND 0.848406f
C96 a_n1455_n3928.n5 GND 0.328934f
C97 a_n1455_n3928.t5 GND 0.081631f
C98 a_n1455_n3928.t0 GND 0.081631f
C99 a_n1455_n3928.n6 GND 0.666694f
C100 a_n1455_n3928.n7 GND 0.352373f
C101 a_n1455_n3928.t4 GND 0.848406f
C102 a_n1455_n3928.n8 GND 0.809652f
C103 a_n1455_n3928.n9 GND 0.77155f
C104 a_n1455_n3928.t1 GND 1.0552f
C105 a_n1455_n3928.n10 GND 0.948443f
C106 a_n1455_n3928.t7 GND 1.05412f
C107 a_n1455_n3928.n11 GND 0.75976f
C108 a_n1455_n3928.t6 GND 1.05412f
C109 a_n1455_n3928.n12 GND 0.985564f
C110 a_n1455_n3928.t2 GND 1.05412f
C111 a_n1455_n3928.n13 GND 1.3206f
C112 a_n1455_n3928.n14 GND 0.860276f
C113 a_n1455_n3928.t18 GND 0.848403f
C114 a_n1455_n3928.n15 GND 0.542321f
C115 a_n1455_n3928.t3 GND 0.081631f
C116 a_n1455_n3928.t16 GND 0.081631f
C117 a_n1455_n3928.n16 GND 0.666693f
C118 a_n1455_n3928.n17 GND 0.352374f
C119 a_n1455_n3928.t19 GND 0.848403f
C120 a_n1455_n3928.n18 GND 0.328937f
C121 a_n1455_n3928.t10 GND 0.848403f
C122 a_n1455_n3928.n19 GND 0.328937f
C123 a_n1455_n3928.n20 GND 0.352377f
C124 a_n1455_n3928.t11 GND 0.081631f
C125 a_n1455_n3928.n21 GND 0.66669f
C126 a_n1455_n3928.t15 GND 0.081631f
C127 a_n2511_10556.t8 GND 0.115035f
C128 a_n2511_10556.t7 GND 0.115035f
C129 a_n2511_10556.t6 GND 0.115035f
C130 a_n2511_10556.n0 GND 0.830094f
C131 a_n2511_10556.t1 GND 0.115035f
C132 a_n2511_10556.t3 GND 0.115035f
C133 a_n2511_10556.n1 GND 0.827337f
C134 a_n2511_10556.n2 GND 2.52538f
C135 a_n2511_10556.t5 GND 0.115035f
C136 a_n2511_10556.t9 GND 0.115035f
C137 a_n2511_10556.n3 GND 0.827337f
C138 a_n2511_10556.n4 GND 3.96056f
C139 a_n2511_10556.n5 GND 0.026557f
C140 a_n2511_10556.n6 GND 0.024262f
C141 a_n2511_10556.n7 GND 0.013037f
C142 a_n2511_10556.n8 GND 0.030816f
C143 a_n2511_10556.n9 GND 0.013804f
C144 a_n2511_10556.n10 GND 0.024262f
C145 a_n2511_10556.n11 GND 0.013037f
C146 a_n2511_10556.n12 GND 0.030816f
C147 a_n2511_10556.n13 GND 0.013804f
C148 a_n2511_10556.n14 GND 0.107274f
C149 a_n2511_10556.t16 GND 0.066122f
C150 a_n2511_10556.n15 GND 0.023112f
C151 a_n2511_10556.n16 GND 0.019593f
C152 a_n2511_10556.n17 GND 0.013037f
C153 a_n2511_10556.n18 GND 0.556554f
C154 a_n2511_10556.n19 GND 0.024262f
C155 a_n2511_10556.n20 GND 0.013037f
C156 a_n2511_10556.n21 GND 0.013804f
C157 a_n2511_10556.n22 GND 0.030816f
C158 a_n2511_10556.n23 GND 0.030816f
C159 a_n2511_10556.n24 GND 0.013804f
C160 a_n2511_10556.n25 GND 0.013037f
C161 a_n2511_10556.n26 GND 0.024262f
C162 a_n2511_10556.n27 GND 0.024262f
C163 a_n2511_10556.n28 GND 0.013037f
C164 a_n2511_10556.n29 GND 0.013804f
C165 a_n2511_10556.n30 GND 0.030816f
C166 a_n2511_10556.n31 GND 0.074256f
C167 a_n2511_10556.n32 GND 0.013804f
C168 a_n2511_10556.n33 GND 0.013037f
C169 a_n2511_10556.n34 GND 0.056081f
C170 a_n2511_10556.n35 GND 0.046363f
C171 a_n2511_10556.t13 GND 0.115035f
C172 a_n2511_10556.t15 GND 0.115035f
C173 a_n2511_10556.n36 GND 0.708188f
C174 a_n2511_10556.n37 GND 1.00643f
C175 a_n2511_10556.n38 GND 0.026557f
C176 a_n2511_10556.n39 GND 0.024262f
C177 a_n2511_10556.n40 GND 0.013037f
C178 a_n2511_10556.n41 GND 0.030816f
C179 a_n2511_10556.n42 GND 0.013804f
C180 a_n2511_10556.n43 GND 0.024262f
C181 a_n2511_10556.n44 GND 0.013037f
C182 a_n2511_10556.n45 GND 0.030816f
C183 a_n2511_10556.n46 GND 0.013804f
C184 a_n2511_10556.n47 GND 0.107274f
C185 a_n2511_10556.t19 GND 0.066122f
C186 a_n2511_10556.n48 GND 0.023112f
C187 a_n2511_10556.n49 GND 0.019593f
C188 a_n2511_10556.n50 GND 0.013037f
C189 a_n2511_10556.n51 GND 0.556554f
C190 a_n2511_10556.n52 GND 0.024262f
C191 a_n2511_10556.n53 GND 0.013037f
C192 a_n2511_10556.n54 GND 0.013804f
C193 a_n2511_10556.n55 GND 0.030816f
C194 a_n2511_10556.n56 GND 0.030816f
C195 a_n2511_10556.n57 GND 0.013804f
C196 a_n2511_10556.n58 GND 0.013037f
C197 a_n2511_10556.n59 GND 0.024262f
C198 a_n2511_10556.n60 GND 0.024262f
C199 a_n2511_10556.n61 GND 0.013037f
C200 a_n2511_10556.n62 GND 0.013804f
C201 a_n2511_10556.n63 GND 0.030816f
C202 a_n2511_10556.n64 GND 0.074256f
C203 a_n2511_10556.n65 GND 0.013804f
C204 a_n2511_10556.n66 GND 0.013037f
C205 a_n2511_10556.n67 GND 0.056081f
C206 a_n2511_10556.n68 GND 0.043002f
C207 a_n2511_10556.n69 GND 0.25396f
C208 a_n2511_10556.n70 GND 0.026557f
C209 a_n2511_10556.n71 GND 0.024262f
C210 a_n2511_10556.n72 GND 0.013037f
C211 a_n2511_10556.n73 GND 0.030816f
C212 a_n2511_10556.n74 GND 0.013804f
C213 a_n2511_10556.n75 GND 0.024262f
C214 a_n2511_10556.n76 GND 0.013037f
C215 a_n2511_10556.n77 GND 0.030816f
C216 a_n2511_10556.n78 GND 0.013804f
C217 a_n2511_10556.n79 GND 0.107274f
C218 a_n2511_10556.t14 GND 0.066122f
C219 a_n2511_10556.n80 GND 0.023112f
C220 a_n2511_10556.n81 GND 0.019593f
C221 a_n2511_10556.n82 GND 0.013037f
C222 a_n2511_10556.n83 GND 0.556554f
C223 a_n2511_10556.n84 GND 0.024262f
C224 a_n2511_10556.n85 GND 0.013037f
C225 a_n2511_10556.n86 GND 0.013804f
C226 a_n2511_10556.n87 GND 0.030816f
C227 a_n2511_10556.n88 GND 0.030816f
C228 a_n2511_10556.n89 GND 0.013804f
C229 a_n2511_10556.n90 GND 0.013037f
C230 a_n2511_10556.n91 GND 0.024262f
C231 a_n2511_10556.n92 GND 0.024262f
C232 a_n2511_10556.n93 GND 0.013037f
C233 a_n2511_10556.n94 GND 0.013804f
C234 a_n2511_10556.n95 GND 0.030816f
C235 a_n2511_10556.n96 GND 0.074256f
C236 a_n2511_10556.n97 GND 0.013804f
C237 a_n2511_10556.n98 GND 0.013037f
C238 a_n2511_10556.n99 GND 0.056081f
C239 a_n2511_10556.n100 GND 0.043002f
C240 a_n2511_10556.n101 GND 0.25396f
C241 a_n2511_10556.t18 GND 0.115035f
C242 a_n2511_10556.t12 GND 0.115035f
C243 a_n2511_10556.n102 GND 0.708188f
C244 a_n2511_10556.n103 GND 0.78481f
C245 a_n2511_10556.n104 GND 0.026557f
C246 a_n2511_10556.n105 GND 0.024262f
C247 a_n2511_10556.n106 GND 0.013037f
C248 a_n2511_10556.n107 GND 0.030816f
C249 a_n2511_10556.n108 GND 0.013804f
C250 a_n2511_10556.n109 GND 0.024262f
C251 a_n2511_10556.n110 GND 0.013037f
C252 a_n2511_10556.n111 GND 0.030816f
C253 a_n2511_10556.n112 GND 0.013804f
C254 a_n2511_10556.n113 GND 0.107274f
C255 a_n2511_10556.t17 GND 0.066122f
C256 a_n2511_10556.n114 GND 0.023112f
C257 a_n2511_10556.n115 GND 0.019593f
C258 a_n2511_10556.n116 GND 0.013037f
C259 a_n2511_10556.n117 GND 0.556554f
C260 a_n2511_10556.n118 GND 0.024262f
C261 a_n2511_10556.n119 GND 0.013037f
C262 a_n2511_10556.n120 GND 0.013804f
C263 a_n2511_10556.n121 GND 0.030816f
C264 a_n2511_10556.n122 GND 0.030816f
C265 a_n2511_10556.n123 GND 0.013804f
C266 a_n2511_10556.n124 GND 0.013037f
C267 a_n2511_10556.n125 GND 0.024262f
C268 a_n2511_10556.n126 GND 0.024262f
C269 a_n2511_10556.n127 GND 0.013037f
C270 a_n2511_10556.n128 GND 0.013804f
C271 a_n2511_10556.n129 GND 0.030816f
C272 a_n2511_10556.n130 GND 0.074256f
C273 a_n2511_10556.n131 GND 0.013804f
C274 a_n2511_10556.n132 GND 0.013037f
C275 a_n2511_10556.n133 GND 0.056081f
C276 a_n2511_10556.n134 GND 0.043002f
C277 a_n2511_10556.n135 GND 1.00759f
C278 a_n2511_10556.n136 GND 2.19047f
C279 a_n2511_10556.t2 GND 0.115035f
C280 a_n2511_10556.t4 GND 0.115035f
C281 a_n2511_10556.n137 GND 0.827334f
C282 a_n2511_10556.n138 GND 1.64036f
C283 a_n2511_10556.t0 GND 0.115035f
C284 a_n2511_10556.t10 GND 0.115035f
C285 a_n2511_10556.n139 GND 0.827337f
C286 a_n2511_10556.n140 GND 1.45743f
C287 a_n2511_10556.n141 GND 0.831205f
C288 a_n2511_10556.t11 GND 0.115035f
C289 VN.n0 GND 0.026927f
C290 VN.t6 GND 0.407734f
C291 VN.t5 GND 0.377008f
C292 VN.n1 GND 0.016298f
C293 VN.t10 GND 0.420161f
C294 VN.n2 GND 0.179365f
C295 VN.t9 GND 0.377008f
C296 VN.n3 GND 0.168383f
C297 VN.n4 GND 0.027517f
C298 VN.n5 GND 0.086386f
C299 VN.n6 GND 0.020179f
C300 VN.n7 GND 0.020179f
C301 VN.n8 GND 0.027517f
C302 VN.n9 GND 0.150426f
C303 VN.n10 GND 0.027678f
C304 VN.n11 GND 0.181643f
C305 VN.n12 GND 0.245126f
C306 VN.n13 GND 0.026927f
C307 VN.t8 GND 0.377008f
C308 VN.n14 GND 0.016298f
C309 VN.t12 GND 0.420161f
C310 VN.n15 GND 0.179365f
C311 VN.t11 GND 0.377008f
C312 VN.n16 GND 0.168383f
C313 VN.n17 GND 0.027517f
C314 VN.n18 GND 0.086386f
C315 VN.n19 GND 0.020179f
C316 VN.n20 GND 0.020179f
C317 VN.n21 GND 0.027517f
C318 VN.n22 GND 0.150426f
C319 VN.n23 GND 0.027678f
C320 VN.t7 GND 0.407734f
C321 VN.n24 GND 0.181643f
C322 VN.n25 GND 0.540126f
C323 VN.n26 GND 0.815822f
C324 VN.t4 GND 0.034835f
C325 VN.t0 GND 0.006221f
C326 VN.t3 GND 0.006221f
C327 VN.n27 GND 0.020174f
C328 VN.n28 GND 0.156617f
C329 VN.t1 GND 0.006221f
C330 VN.t2 GND 0.006221f
C331 VN.n29 GND 0.020174f
C332 VN.n30 GND 0.11756f
C333 VN.n31 GND 1.9292f
C334 CS_BIAS.n0 GND 0.007636f
C335 CS_BIAS.t63 GND 0.183962f
C336 CS_BIAS.n1 GND 0.008259f
C337 CS_BIAS.n2 GND 0.005792f
C338 CS_BIAS.t44 GND 0.183962f
C339 CS_BIAS.n3 GND 0.005305f
C340 CS_BIAS.n4 GND 0.005792f
C341 CS_BIAS.t46 GND 0.183962f
C342 CS_BIAS.n5 GND 0.010793f
C343 CS_BIAS.n6 GND 0.005792f
C344 CS_BIAS.t45 GND 0.183962f
C345 CS_BIAS.n7 GND 0.07023f
C346 CS_BIAS.n8 GND 0.00506f
C347 CS_BIAS.n9 GND 0.009839f
C348 CS_BIAS.n10 GND 0.007636f
C349 CS_BIAS.t18 GND 0.183962f
C350 CS_BIAS.n11 GND 0.008259f
C351 CS_BIAS.n12 GND 0.005792f
C352 CS_BIAS.t24 GND 0.183962f
C353 CS_BIAS.n13 GND 0.005305f
C354 CS_BIAS.n14 GND 0.005792f
C355 CS_BIAS.t10 GND 0.183962f
C356 CS_BIAS.n15 GND 0.010793f
C357 CS_BIAS.n16 GND 0.005792f
C358 CS_BIAS.t2 GND 0.183962f
C359 CS_BIAS.n17 GND 0.07023f
C360 CS_BIAS.n18 GND 0.005792f
C361 CS_BIAS.n19 GND 0.009839f
C362 CS_BIAS.n20 GND 0.005792f
C363 CS_BIAS.t20 GND 0.183962f
C364 CS_BIAS.n21 GND 0.07023f
C365 CS_BIAS.n22 GND 0.010793f
C366 CS_BIAS.n23 GND 0.005792f
C367 CS_BIAS.t0 GND 0.183962f
C368 CS_BIAS.n24 GND 0.005305f
C369 CS_BIAS.n25 GND 0.043358f
C370 CS_BIAS.t26 GND 0.183962f
C371 CS_BIAS.t14 GND 0.213079f
C372 CS_BIAS.n26 GND 0.084349f
C373 CS_BIAS.n27 GND 0.082279f
C374 CS_BIAS.n28 GND 0.006234f
C375 CS_BIAS.n29 GND 0.011587f
C376 CS_BIAS.n30 GND 0.005792f
C377 CS_BIAS.n31 GND 0.005792f
C378 CS_BIAS.n32 GND 0.005792f
C379 CS_BIAS.n33 GND 0.010688f
C380 CS_BIAS.n34 GND 0.008143f
C381 CS_BIAS.n35 GND 0.07023f
C382 CS_BIAS.n36 GND 0.008037f
C383 CS_BIAS.n37 GND 0.005792f
C384 CS_BIAS.n38 GND 0.005792f
C385 CS_BIAS.n39 GND 0.005792f
C386 CS_BIAS.n40 GND 0.005168f
C387 CS_BIAS.n41 GND 0.011619f
C388 CS_BIAS.n42 GND 0.00634f
C389 CS_BIAS.n43 GND 0.005792f
C390 CS_BIAS.n44 GND 0.005792f
C391 CS_BIAS.n45 GND 0.005792f
C392 CS_BIAS.n46 GND 0.00842f
C393 CS_BIAS.n47 GND 0.00842f
C394 CS_BIAS.n48 GND 0.009839f
C395 CS_BIAS.n49 GND 0.005792f
C396 CS_BIAS.n50 GND 0.005792f
C397 CS_BIAS.n51 GND 0.00634f
C398 CS_BIAS.n52 GND 0.011619f
C399 CS_BIAS.n53 GND 0.005168f
C400 CS_BIAS.n54 GND 0.005792f
C401 CS_BIAS.n55 GND 0.005792f
C402 CS_BIAS.n56 GND 0.005792f
C403 CS_BIAS.n57 GND 0.008037f
C404 CS_BIAS.n58 GND 0.07023f
C405 CS_BIAS.n59 GND 0.008143f
C406 CS_BIAS.n60 GND 0.010688f
C407 CS_BIAS.n61 GND 0.005792f
C408 CS_BIAS.n62 GND 0.005792f
C409 CS_BIAS.n63 GND 0.005792f
C410 CS_BIAS.n64 GND 0.011587f
C411 CS_BIAS.n65 GND 0.006234f
C412 CS_BIAS.n66 GND 0.07023f
C413 CS_BIAS.n67 GND 0.009945f
C414 CS_BIAS.n68 GND 0.005792f
C415 CS_BIAS.n69 GND 0.005792f
C416 CS_BIAS.n70 GND 0.005792f
C417 CS_BIAS.n71 GND 0.00858f
C418 CS_BIAS.n72 GND 0.009733f
C419 CS_BIAS.n73 GND 0.087892f
C420 CS_BIAS.n74 GND 0.058174f
C421 CS_BIAS.t19 GND 0.010713f
C422 CS_BIAS.t25 GND 0.010713f
C423 CS_BIAS.n75 GND 0.093562f
C424 CS_BIAS.n76 GND 0.115968f
C425 CS_BIAS.t11 GND 0.010713f
C426 CS_BIAS.t3 GND 0.010713f
C427 CS_BIAS.n77 GND 0.093562f
C428 CS_BIAS.n78 GND 0.061102f
C429 CS_BIAS.t27 GND 0.010713f
C430 CS_BIAS.t15 GND 0.010713f
C431 CS_BIAS.n79 GND 0.094477f
C432 CS_BIAS.t21 GND 0.010713f
C433 CS_BIAS.t1 GND 0.010713f
C434 CS_BIAS.n80 GND 0.093562f
C435 CS_BIAS.n81 GND 0.137733f
C436 CS_BIAS.n82 GND 0.063874f
C437 CS_BIAS.n83 GND 0.037486f
C438 CS_BIAS.n84 GND 0.005792f
C439 CS_BIAS.t61 GND 0.183962f
C440 CS_BIAS.n85 GND 0.07023f
C441 CS_BIAS.n86 GND 0.010793f
C442 CS_BIAS.n87 GND 0.005792f
C443 CS_BIAS.t62 GND 0.183962f
C444 CS_BIAS.n88 GND 0.005305f
C445 CS_BIAS.n89 GND 0.043358f
C446 CS_BIAS.t50 GND 0.183962f
C447 CS_BIAS.t54 GND 0.213079f
C448 CS_BIAS.n90 GND 0.084349f
C449 CS_BIAS.n91 GND 0.082279f
C450 CS_BIAS.n92 GND 0.006234f
C451 CS_BIAS.n93 GND 0.011587f
C452 CS_BIAS.n94 GND 0.005792f
C453 CS_BIAS.n95 GND 0.005792f
C454 CS_BIAS.n96 GND 0.005792f
C455 CS_BIAS.n97 GND 0.010688f
C456 CS_BIAS.n98 GND 0.008143f
C457 CS_BIAS.n99 GND 0.07023f
C458 CS_BIAS.n100 GND 0.008037f
C459 CS_BIAS.n101 GND 0.005792f
C460 CS_BIAS.n102 GND 0.005792f
C461 CS_BIAS.n103 GND 0.005792f
C462 CS_BIAS.n104 GND 0.005168f
C463 CS_BIAS.n105 GND 0.011619f
C464 CS_BIAS.n106 GND 0.00634f
C465 CS_BIAS.n107 GND 0.005792f
C466 CS_BIAS.n108 GND 0.005792f
C467 CS_BIAS.n109 GND 0.00506f
C468 CS_BIAS.n110 GND 0.00842f
C469 CS_BIAS.n111 GND 0.00842f
C470 CS_BIAS.n112 GND 0.009839f
C471 CS_BIAS.n113 GND 0.005792f
C472 CS_BIAS.n114 GND 0.005792f
C473 CS_BIAS.n115 GND 0.00634f
C474 CS_BIAS.n116 GND 0.011619f
C475 CS_BIAS.n117 GND 0.005168f
C476 CS_BIAS.n118 GND 0.005792f
C477 CS_BIAS.n119 GND 0.005792f
C478 CS_BIAS.n120 GND 0.005792f
C479 CS_BIAS.n121 GND 0.008037f
C480 CS_BIAS.n122 GND 0.07023f
C481 CS_BIAS.n123 GND 0.008143f
C482 CS_BIAS.n124 GND 0.010688f
C483 CS_BIAS.n125 GND 0.005792f
C484 CS_BIAS.n126 GND 0.005792f
C485 CS_BIAS.n127 GND 0.005792f
C486 CS_BIAS.n128 GND 0.011587f
C487 CS_BIAS.n129 GND 0.006234f
C488 CS_BIAS.n130 GND 0.07023f
C489 CS_BIAS.n131 GND 0.009945f
C490 CS_BIAS.n132 GND 0.005792f
C491 CS_BIAS.n133 GND 0.005792f
C492 CS_BIAS.n134 GND 0.005792f
C493 CS_BIAS.n135 GND 0.00858f
C494 CS_BIAS.n136 GND 0.009733f
C495 CS_BIAS.n137 GND 0.087892f
C496 CS_BIAS.n138 GND 0.034855f
C497 CS_BIAS.n139 GND 0.007636f
C498 CS_BIAS.t38 GND 0.183962f
C499 CS_BIAS.n140 GND 0.008259f
C500 CS_BIAS.n141 GND 0.005792f
C501 CS_BIAS.t51 GND 0.183962f
C502 CS_BIAS.n142 GND 0.005305f
C503 CS_BIAS.n143 GND 0.005792f
C504 CS_BIAS.t55 GND 0.183962f
C505 CS_BIAS.n144 GND 0.010793f
C506 CS_BIAS.n145 GND 0.005792f
C507 CS_BIAS.t52 GND 0.183962f
C508 CS_BIAS.n146 GND 0.07023f
C509 CS_BIAS.n147 GND 0.005792f
C510 CS_BIAS.n148 GND 0.009839f
C511 CS_BIAS.n149 GND 0.005792f
C512 CS_BIAS.t34 GND 0.183962f
C513 CS_BIAS.n150 GND 0.07023f
C514 CS_BIAS.n151 GND 0.010793f
C515 CS_BIAS.n152 GND 0.005792f
C516 CS_BIAS.t35 GND 0.183962f
C517 CS_BIAS.n153 GND 0.005305f
C518 CS_BIAS.n154 GND 0.043358f
C519 CS_BIAS.t57 GND 0.183962f
C520 CS_BIAS.t60 GND 0.213079f
C521 CS_BIAS.n155 GND 0.084349f
C522 CS_BIAS.n156 GND 0.082279f
C523 CS_BIAS.n157 GND 0.006234f
C524 CS_BIAS.n158 GND 0.011587f
C525 CS_BIAS.n159 GND 0.005792f
C526 CS_BIAS.n160 GND 0.005792f
C527 CS_BIAS.n161 GND 0.005792f
C528 CS_BIAS.n162 GND 0.010688f
C529 CS_BIAS.n163 GND 0.008143f
C530 CS_BIAS.n164 GND 0.07023f
C531 CS_BIAS.n165 GND 0.008037f
C532 CS_BIAS.n166 GND 0.005792f
C533 CS_BIAS.n167 GND 0.005792f
C534 CS_BIAS.n168 GND 0.005792f
C535 CS_BIAS.n169 GND 0.005168f
C536 CS_BIAS.n170 GND 0.011619f
C537 CS_BIAS.n171 GND 0.00634f
C538 CS_BIAS.n172 GND 0.005792f
C539 CS_BIAS.n173 GND 0.005792f
C540 CS_BIAS.n174 GND 0.005792f
C541 CS_BIAS.n175 GND 0.00842f
C542 CS_BIAS.n176 GND 0.00842f
C543 CS_BIAS.n177 GND 0.009839f
C544 CS_BIAS.n178 GND 0.005792f
C545 CS_BIAS.n179 GND 0.005792f
C546 CS_BIAS.n180 GND 0.00634f
C547 CS_BIAS.n181 GND 0.011619f
C548 CS_BIAS.n182 GND 0.005168f
C549 CS_BIAS.n183 GND 0.005792f
C550 CS_BIAS.n184 GND 0.005792f
C551 CS_BIAS.n185 GND 0.005792f
C552 CS_BIAS.n186 GND 0.008037f
C553 CS_BIAS.n187 GND 0.07023f
C554 CS_BIAS.n188 GND 0.008143f
C555 CS_BIAS.n189 GND 0.010688f
C556 CS_BIAS.n190 GND 0.005792f
C557 CS_BIAS.n191 GND 0.005792f
C558 CS_BIAS.n192 GND 0.005792f
C559 CS_BIAS.n193 GND 0.011587f
C560 CS_BIAS.n194 GND 0.006234f
C561 CS_BIAS.n195 GND 0.07023f
C562 CS_BIAS.n196 GND 0.009945f
C563 CS_BIAS.n197 GND 0.005792f
C564 CS_BIAS.n198 GND 0.005792f
C565 CS_BIAS.n199 GND 0.005792f
C566 CS_BIAS.n200 GND 0.00858f
C567 CS_BIAS.n201 GND 0.009733f
C568 CS_BIAS.n202 GND 0.087892f
C569 CS_BIAS.n203 GND 0.020992f
C570 CS_BIAS.n204 GND 0.262164f
C571 CS_BIAS.n205 GND 0.007636f
C572 CS_BIAS.t43 GND 0.183962f
C573 CS_BIAS.n206 GND 0.008259f
C574 CS_BIAS.n207 GND 0.005792f
C575 CS_BIAS.t37 GND 0.183962f
C576 CS_BIAS.n208 GND 0.005305f
C577 CS_BIAS.n209 GND 0.005792f
C578 CS_BIAS.t59 GND 0.183962f
C579 CS_BIAS.n210 GND 0.010793f
C580 CS_BIAS.n211 GND 0.005792f
C581 CS_BIAS.t36 GND 0.183962f
C582 CS_BIAS.n212 GND 0.07023f
C583 CS_BIAS.n213 GND 0.00506f
C584 CS_BIAS.n214 GND 0.009839f
C585 CS_BIAS.n215 GND 0.005792f
C586 CS_BIAS.n216 GND 0.010793f
C587 CS_BIAS.n217 GND 0.005792f
C588 CS_BIAS.t53 GND 0.183962f
C589 CS_BIAS.n218 GND 0.005305f
C590 CS_BIAS.n219 GND 0.043358f
C591 CS_BIAS.t40 GND 0.183962f
C592 CS_BIAS.t32 GND 0.213079f
C593 CS_BIAS.n220 GND 0.084349f
C594 CS_BIAS.n221 GND 0.082279f
C595 CS_BIAS.n222 GND 0.006234f
C596 CS_BIAS.n223 GND 0.011587f
C597 CS_BIAS.n224 GND 0.005792f
C598 CS_BIAS.n225 GND 0.005792f
C599 CS_BIAS.n226 GND 0.005792f
C600 CS_BIAS.n227 GND 0.010688f
C601 CS_BIAS.n228 GND 0.008143f
C602 CS_BIAS.n229 GND 0.07023f
C603 CS_BIAS.n230 GND 0.008037f
C604 CS_BIAS.n231 GND 0.005792f
C605 CS_BIAS.n232 GND 0.005792f
C606 CS_BIAS.n233 GND 0.005792f
C607 CS_BIAS.n234 GND 0.005168f
C608 CS_BIAS.n235 GND 0.011619f
C609 CS_BIAS.t49 GND 0.183962f
C610 CS_BIAS.n236 GND 0.07023f
C611 CS_BIAS.n237 GND 0.00634f
C612 CS_BIAS.n238 GND 0.005792f
C613 CS_BIAS.n239 GND 0.005792f
C614 CS_BIAS.t13 GND 0.010713f
C615 CS_BIAS.t31 GND 0.010713f
C616 CS_BIAS.n240 GND 0.094477f
C617 CS_BIAS.t5 GND 0.010713f
C618 CS_BIAS.t23 GND 0.010713f
C619 CS_BIAS.n241 GND 0.093562f
C620 CS_BIAS.n242 GND 0.137733f
C621 CS_BIAS.n243 GND 0.007636f
C622 CS_BIAS.t16 GND 0.183962f
C623 CS_BIAS.n244 GND 0.008259f
C624 CS_BIAS.n245 GND 0.005792f
C625 CS_BIAS.t28 GND 0.183962f
C626 CS_BIAS.n246 GND 0.005305f
C627 CS_BIAS.n247 GND 0.005792f
C628 CS_BIAS.t8 GND 0.183962f
C629 CS_BIAS.n248 GND 0.010793f
C630 CS_BIAS.n249 GND 0.005792f
C631 CS_BIAS.t6 GND 0.183962f
C632 CS_BIAS.n250 GND 0.07023f
C633 CS_BIAS.n251 GND 0.005792f
C634 CS_BIAS.n252 GND 0.009839f
C635 CS_BIAS.n253 GND 0.005792f
C636 CS_BIAS.n254 GND 0.010793f
C637 CS_BIAS.n255 GND 0.005792f
C638 CS_BIAS.t4 GND 0.183962f
C639 CS_BIAS.n256 GND 0.005305f
C640 CS_BIAS.n257 GND 0.043358f
C641 CS_BIAS.t30 GND 0.183962f
C642 CS_BIAS.t12 GND 0.213079f
C643 CS_BIAS.n258 GND 0.084349f
C644 CS_BIAS.n259 GND 0.082279f
C645 CS_BIAS.n260 GND 0.006234f
C646 CS_BIAS.n261 GND 0.011587f
C647 CS_BIAS.n262 GND 0.005792f
C648 CS_BIAS.n263 GND 0.005792f
C649 CS_BIAS.n264 GND 0.005792f
C650 CS_BIAS.n265 GND 0.010688f
C651 CS_BIAS.n266 GND 0.008143f
C652 CS_BIAS.n267 GND 0.07023f
C653 CS_BIAS.n268 GND 0.008037f
C654 CS_BIAS.n269 GND 0.005792f
C655 CS_BIAS.n270 GND 0.005792f
C656 CS_BIAS.n271 GND 0.005792f
C657 CS_BIAS.n272 GND 0.005168f
C658 CS_BIAS.n273 GND 0.011619f
C659 CS_BIAS.t22 GND 0.183962f
C660 CS_BIAS.n274 GND 0.07023f
C661 CS_BIAS.n275 GND 0.00634f
C662 CS_BIAS.n276 GND 0.005792f
C663 CS_BIAS.n277 GND 0.005792f
C664 CS_BIAS.n278 GND 0.005792f
C665 CS_BIAS.n279 GND 0.00842f
C666 CS_BIAS.n280 GND 0.00842f
C667 CS_BIAS.n281 GND 0.009839f
C668 CS_BIAS.n282 GND 0.005792f
C669 CS_BIAS.n283 GND 0.005792f
C670 CS_BIAS.n284 GND 0.00634f
C671 CS_BIAS.n285 GND 0.011619f
C672 CS_BIAS.n286 GND 0.005168f
C673 CS_BIAS.n287 GND 0.005792f
C674 CS_BIAS.n288 GND 0.005792f
C675 CS_BIAS.n289 GND 0.005792f
C676 CS_BIAS.n290 GND 0.008037f
C677 CS_BIAS.n291 GND 0.07023f
C678 CS_BIAS.n292 GND 0.008143f
C679 CS_BIAS.n293 GND 0.010688f
C680 CS_BIAS.n294 GND 0.005792f
C681 CS_BIAS.n295 GND 0.005792f
C682 CS_BIAS.n296 GND 0.005792f
C683 CS_BIAS.n297 GND 0.011587f
C684 CS_BIAS.n298 GND 0.006234f
C685 CS_BIAS.n299 GND 0.07023f
C686 CS_BIAS.n300 GND 0.009945f
C687 CS_BIAS.n301 GND 0.005792f
C688 CS_BIAS.n302 GND 0.005792f
C689 CS_BIAS.n303 GND 0.005792f
C690 CS_BIAS.n304 GND 0.00858f
C691 CS_BIAS.n305 GND 0.009733f
C692 CS_BIAS.n306 GND 0.087892f
C693 CS_BIAS.n307 GND 0.058174f
C694 CS_BIAS.t29 GND 0.010713f
C695 CS_BIAS.t17 GND 0.010713f
C696 CS_BIAS.n308 GND 0.093562f
C697 CS_BIAS.n309 GND 0.115968f
C698 CS_BIAS.t7 GND 0.010713f
C699 CS_BIAS.t9 GND 0.010713f
C700 CS_BIAS.n310 GND 0.093562f
C701 CS_BIAS.n311 GND 0.061102f
C702 CS_BIAS.n312 GND 0.063874f
C703 CS_BIAS.n313 GND 0.037486f
C704 CS_BIAS.n314 GND 0.00506f
C705 CS_BIAS.n315 GND 0.00842f
C706 CS_BIAS.n316 GND 0.00842f
C707 CS_BIAS.n317 GND 0.009839f
C708 CS_BIAS.n318 GND 0.005792f
C709 CS_BIAS.n319 GND 0.005792f
C710 CS_BIAS.n320 GND 0.00634f
C711 CS_BIAS.n321 GND 0.011619f
C712 CS_BIAS.n322 GND 0.005168f
C713 CS_BIAS.n323 GND 0.005792f
C714 CS_BIAS.n324 GND 0.005792f
C715 CS_BIAS.n325 GND 0.005792f
C716 CS_BIAS.n326 GND 0.008037f
C717 CS_BIAS.n327 GND 0.07023f
C718 CS_BIAS.n328 GND 0.008143f
C719 CS_BIAS.n329 GND 0.010688f
C720 CS_BIAS.n330 GND 0.005792f
C721 CS_BIAS.n331 GND 0.005792f
C722 CS_BIAS.n332 GND 0.005792f
C723 CS_BIAS.n333 GND 0.011587f
C724 CS_BIAS.n334 GND 0.006234f
C725 CS_BIAS.n335 GND 0.07023f
C726 CS_BIAS.n336 GND 0.009945f
C727 CS_BIAS.n337 GND 0.005792f
C728 CS_BIAS.n338 GND 0.005792f
C729 CS_BIAS.n339 GND 0.005792f
C730 CS_BIAS.n340 GND 0.00858f
C731 CS_BIAS.n341 GND 0.009733f
C732 CS_BIAS.n342 GND 0.087892f
C733 CS_BIAS.n343 GND 0.034855f
C734 CS_BIAS.n344 GND 0.007636f
C735 CS_BIAS.t48 GND 0.183962f
C736 CS_BIAS.n345 GND 0.008259f
C737 CS_BIAS.n346 GND 0.005792f
C738 CS_BIAS.t41 GND 0.183962f
C739 CS_BIAS.n347 GND 0.005305f
C740 CS_BIAS.n348 GND 0.005792f
C741 CS_BIAS.t33 GND 0.183962f
C742 CS_BIAS.n349 GND 0.010793f
C743 CS_BIAS.n350 GND 0.005792f
C744 CS_BIAS.t42 GND 0.183962f
C745 CS_BIAS.n351 GND 0.07023f
C746 CS_BIAS.n352 GND 0.005792f
C747 CS_BIAS.n353 GND 0.009839f
C748 CS_BIAS.n354 GND 0.005792f
C749 CS_BIAS.n355 GND 0.010793f
C750 CS_BIAS.n356 GND 0.005792f
C751 CS_BIAS.t58 GND 0.183962f
C752 CS_BIAS.n357 GND 0.005305f
C753 CS_BIAS.n358 GND 0.043358f
C754 CS_BIAS.t47 GND 0.183962f
C755 CS_BIAS.t39 GND 0.213079f
C756 CS_BIAS.n359 GND 0.084349f
C757 CS_BIAS.n360 GND 0.082279f
C758 CS_BIAS.n361 GND 0.006234f
C759 CS_BIAS.n362 GND 0.011587f
C760 CS_BIAS.n363 GND 0.005792f
C761 CS_BIAS.n364 GND 0.005792f
C762 CS_BIAS.n365 GND 0.005792f
C763 CS_BIAS.n366 GND 0.010688f
C764 CS_BIAS.n367 GND 0.008143f
C765 CS_BIAS.n368 GND 0.07023f
C766 CS_BIAS.n369 GND 0.008037f
C767 CS_BIAS.n370 GND 0.005792f
C768 CS_BIAS.n371 GND 0.005792f
C769 CS_BIAS.n372 GND 0.005792f
C770 CS_BIAS.n373 GND 0.005168f
C771 CS_BIAS.n374 GND 0.011619f
C772 CS_BIAS.t56 GND 0.183962f
C773 CS_BIAS.n375 GND 0.07023f
C774 CS_BIAS.n376 GND 0.00634f
C775 CS_BIAS.n377 GND 0.005792f
C776 CS_BIAS.n378 GND 0.005792f
C777 CS_BIAS.n379 GND 0.005792f
C778 CS_BIAS.n380 GND 0.00842f
C779 CS_BIAS.n381 GND 0.00842f
C780 CS_BIAS.n382 GND 0.009839f
C781 CS_BIAS.n383 GND 0.005792f
C782 CS_BIAS.n384 GND 0.005792f
C783 CS_BIAS.n385 GND 0.00634f
C784 CS_BIAS.n386 GND 0.011619f
C785 CS_BIAS.n387 GND 0.005168f
C786 CS_BIAS.n388 GND 0.005792f
C787 CS_BIAS.n389 GND 0.005792f
C788 CS_BIAS.n390 GND 0.005792f
C789 CS_BIAS.n391 GND 0.008037f
C790 CS_BIAS.n392 GND 0.07023f
C791 CS_BIAS.n393 GND 0.008143f
C792 CS_BIAS.n394 GND 0.010688f
C793 CS_BIAS.n395 GND 0.005792f
C794 CS_BIAS.n396 GND 0.005792f
C795 CS_BIAS.n397 GND 0.005792f
C796 CS_BIAS.n398 GND 0.011587f
C797 CS_BIAS.n399 GND 0.006234f
C798 CS_BIAS.n400 GND 0.07023f
C799 CS_BIAS.n401 GND 0.009945f
C800 CS_BIAS.n402 GND 0.005792f
C801 CS_BIAS.n403 GND 0.005792f
C802 CS_BIAS.n404 GND 0.005792f
C803 CS_BIAS.n405 GND 0.00858f
C804 CS_BIAS.n406 GND 0.009733f
C805 CS_BIAS.n407 GND 0.087892f
C806 CS_BIAS.n408 GND 0.020992f
C807 CS_BIAS.n409 GND 0.157331f
C808 CS_BIAS.n410 GND 2.90828f
C809 a_n2686_8422.t20 GND 98.0738f
C810 a_n2686_8422.t9 GND 0.049091f
C811 a_n2686_8422.n0 GND 0.011333f
C812 a_n2686_8422.n1 GND 0.010354f
C813 a_n2686_8422.n2 GND 0.005564f
C814 a_n2686_8422.n3 GND 0.01315f
C815 a_n2686_8422.n4 GND 0.005891f
C816 a_n2686_8422.n5 GND 0.010354f
C817 a_n2686_8422.n6 GND 0.005564f
C818 a_n2686_8422.n7 GND 0.01315f
C819 a_n2686_8422.n8 GND 0.005891f
C820 a_n2686_8422.n9 GND 0.045779f
C821 a_n2686_8422.t15 GND 0.028217f
C822 a_n2686_8422.n10 GND 0.009863f
C823 a_n2686_8422.n11 GND 0.008361f
C824 a_n2686_8422.n12 GND 0.005564f
C825 a_n2686_8422.n13 GND 0.237506f
C826 a_n2686_8422.n14 GND 0.010354f
C827 a_n2686_8422.n15 GND 0.005564f
C828 a_n2686_8422.n16 GND 0.005891f
C829 a_n2686_8422.n17 GND 0.01315f
C830 a_n2686_8422.n18 GND 0.01315f
C831 a_n2686_8422.n19 GND 0.005891f
C832 a_n2686_8422.n20 GND 0.005564f
C833 a_n2686_8422.n21 GND 0.010354f
C834 a_n2686_8422.n22 GND 0.010354f
C835 a_n2686_8422.n23 GND 0.005564f
C836 a_n2686_8422.n24 GND 0.005891f
C837 a_n2686_8422.n25 GND 0.01315f
C838 a_n2686_8422.n26 GND 0.031688f
C839 a_n2686_8422.n27 GND 0.005891f
C840 a_n2686_8422.n28 GND 0.005564f
C841 a_n2686_8422.n29 GND 0.023932f
C842 a_n2686_8422.n30 GND 0.019785f
C843 a_n2686_8422.t18 GND 0.049091f
C844 a_n2686_8422.t14 GND 0.049091f
C845 a_n2686_8422.n31 GND 0.302215f
C846 a_n2686_8422.n32 GND 0.429488f
C847 a_n2686_8422.t12 GND 0.049091f
C848 a_n2686_8422.t13 GND 0.049091f
C849 a_n2686_8422.n33 GND 0.302215f
C850 a_n2686_8422.n34 GND 0.334913f
C851 a_n2686_8422.n35 GND 0.011333f
C852 a_n2686_8422.n36 GND 0.010354f
C853 a_n2686_8422.n37 GND 0.005564f
C854 a_n2686_8422.n38 GND 0.01315f
C855 a_n2686_8422.n39 GND 0.005891f
C856 a_n2686_8422.n40 GND 0.010354f
C857 a_n2686_8422.n41 GND 0.005564f
C858 a_n2686_8422.n42 GND 0.01315f
C859 a_n2686_8422.n43 GND 0.005891f
C860 a_n2686_8422.n44 GND 0.045779f
C861 a_n2686_8422.t16 GND 0.028217f
C862 a_n2686_8422.n45 GND 0.009863f
C863 a_n2686_8422.n46 GND 0.008361f
C864 a_n2686_8422.n47 GND 0.005564f
C865 a_n2686_8422.n48 GND 0.237506f
C866 a_n2686_8422.n49 GND 0.010354f
C867 a_n2686_8422.n50 GND 0.005564f
C868 a_n2686_8422.n51 GND 0.005891f
C869 a_n2686_8422.n52 GND 0.01315f
C870 a_n2686_8422.n53 GND 0.01315f
C871 a_n2686_8422.n54 GND 0.005891f
C872 a_n2686_8422.n55 GND 0.005564f
C873 a_n2686_8422.n56 GND 0.010354f
C874 a_n2686_8422.n57 GND 0.010354f
C875 a_n2686_8422.n58 GND 0.005564f
C876 a_n2686_8422.n59 GND 0.005891f
C877 a_n2686_8422.n60 GND 0.01315f
C878 a_n2686_8422.n61 GND 0.031688f
C879 a_n2686_8422.n62 GND 0.005891f
C880 a_n2686_8422.n63 GND 0.005564f
C881 a_n2686_8422.n64 GND 0.023932f
C882 a_n2686_8422.n65 GND 0.018351f
C883 a_n2686_8422.n66 GND 0.955844f
C884 a_n2686_8422.n67 GND 0.011333f
C885 a_n2686_8422.n68 GND 0.010354f
C886 a_n2686_8422.n69 GND 0.005564f
C887 a_n2686_8422.n70 GND 0.01315f
C888 a_n2686_8422.n71 GND 0.005891f
C889 a_n2686_8422.n72 GND 0.010354f
C890 a_n2686_8422.n73 GND 0.005564f
C891 a_n2686_8422.n74 GND 0.01315f
C892 a_n2686_8422.n75 GND 0.005891f
C893 a_n2686_8422.n76 GND 0.045779f
C894 a_n2686_8422.t6 GND 0.028217f
C895 a_n2686_8422.n77 GND 0.009863f
C896 a_n2686_8422.n78 GND 0.008361f
C897 a_n2686_8422.n79 GND 0.005564f
C898 a_n2686_8422.n80 GND 0.237506f
C899 a_n2686_8422.n81 GND 0.010354f
C900 a_n2686_8422.n82 GND 0.005564f
C901 a_n2686_8422.n83 GND 0.005891f
C902 a_n2686_8422.n84 GND 0.01315f
C903 a_n2686_8422.n85 GND 0.01315f
C904 a_n2686_8422.n86 GND 0.005891f
C905 a_n2686_8422.n87 GND 0.005564f
C906 a_n2686_8422.n88 GND 0.010354f
C907 a_n2686_8422.n89 GND 0.010354f
C908 a_n2686_8422.n90 GND 0.005564f
C909 a_n2686_8422.n91 GND 0.005891f
C910 a_n2686_8422.n92 GND 0.01315f
C911 a_n2686_8422.n93 GND 0.031688f
C912 a_n2686_8422.n94 GND 0.005891f
C913 a_n2686_8422.n95 GND 0.005564f
C914 a_n2686_8422.n96 GND 0.023932f
C915 a_n2686_8422.n97 GND 0.019785f
C916 a_n2686_8422.t4 GND 0.049091f
C917 a_n2686_8422.t2 GND 0.049091f
C918 a_n2686_8422.n98 GND 0.302215f
C919 a_n2686_8422.n99 GND 0.429488f
C920 a_n2686_8422.n100 GND 0.011333f
C921 a_n2686_8422.n101 GND 0.010354f
C922 a_n2686_8422.n102 GND 0.005564f
C923 a_n2686_8422.n103 GND 0.01315f
C924 a_n2686_8422.n104 GND 0.005891f
C925 a_n2686_8422.n105 GND 0.010354f
C926 a_n2686_8422.n106 GND 0.005564f
C927 a_n2686_8422.n107 GND 0.01315f
C928 a_n2686_8422.n108 GND 0.005891f
C929 a_n2686_8422.n109 GND 0.045779f
C930 a_n2686_8422.t1 GND 0.028217f
C931 a_n2686_8422.n110 GND 0.009863f
C932 a_n2686_8422.n111 GND 0.008361f
C933 a_n2686_8422.n112 GND 0.005564f
C934 a_n2686_8422.n113 GND 0.237506f
C935 a_n2686_8422.n114 GND 0.010354f
C936 a_n2686_8422.n115 GND 0.005564f
C937 a_n2686_8422.n116 GND 0.005891f
C938 a_n2686_8422.n117 GND 0.01315f
C939 a_n2686_8422.n118 GND 0.01315f
C940 a_n2686_8422.n119 GND 0.005891f
C941 a_n2686_8422.n120 GND 0.005564f
C942 a_n2686_8422.n121 GND 0.010354f
C943 a_n2686_8422.n122 GND 0.010354f
C944 a_n2686_8422.n123 GND 0.005564f
C945 a_n2686_8422.n124 GND 0.005891f
C946 a_n2686_8422.n125 GND 0.01315f
C947 a_n2686_8422.n126 GND 0.031688f
C948 a_n2686_8422.n127 GND 0.005891f
C949 a_n2686_8422.n128 GND 0.005564f
C950 a_n2686_8422.n129 GND 0.023932f
C951 a_n2686_8422.n130 GND 0.018351f
C952 a_n2686_8422.n131 GND 0.108376f
C953 a_n2686_8422.n132 GND 0.011333f
C954 a_n2686_8422.n133 GND 0.010354f
C955 a_n2686_8422.n134 GND 0.005564f
C956 a_n2686_8422.n135 GND 0.01315f
C957 a_n2686_8422.n136 GND 0.005891f
C958 a_n2686_8422.n137 GND 0.010354f
C959 a_n2686_8422.n138 GND 0.005564f
C960 a_n2686_8422.n139 GND 0.01315f
C961 a_n2686_8422.n140 GND 0.005891f
C962 a_n2686_8422.n141 GND 0.045779f
C963 a_n2686_8422.t5 GND 0.028217f
C964 a_n2686_8422.n142 GND 0.009863f
C965 a_n2686_8422.n143 GND 0.008361f
C966 a_n2686_8422.n144 GND 0.005564f
C967 a_n2686_8422.n145 GND 0.237506f
C968 a_n2686_8422.n146 GND 0.010354f
C969 a_n2686_8422.n147 GND 0.005564f
C970 a_n2686_8422.n148 GND 0.005891f
C971 a_n2686_8422.n149 GND 0.01315f
C972 a_n2686_8422.n150 GND 0.01315f
C973 a_n2686_8422.n151 GND 0.005891f
C974 a_n2686_8422.n152 GND 0.005564f
C975 a_n2686_8422.n153 GND 0.010354f
C976 a_n2686_8422.n154 GND 0.010354f
C977 a_n2686_8422.n155 GND 0.005564f
C978 a_n2686_8422.n156 GND 0.005891f
C979 a_n2686_8422.n157 GND 0.01315f
C980 a_n2686_8422.n158 GND 0.031688f
C981 a_n2686_8422.n159 GND 0.005891f
C982 a_n2686_8422.n160 GND 0.005564f
C983 a_n2686_8422.n161 GND 0.023932f
C984 a_n2686_8422.n162 GND 0.018351f
C985 a_n2686_8422.n163 GND 0.108376f
C986 a_n2686_8422.t3 GND 0.049091f
C987 a_n2686_8422.t0 GND 0.049091f
C988 a_n2686_8422.n164 GND 0.302215f
C989 a_n2686_8422.n165 GND 0.334913f
C990 a_n2686_8422.n166 GND 0.011333f
C991 a_n2686_8422.n167 GND 0.010354f
C992 a_n2686_8422.n168 GND 0.005564f
C993 a_n2686_8422.n169 GND 0.01315f
C994 a_n2686_8422.n170 GND 0.005891f
C995 a_n2686_8422.n171 GND 0.010354f
C996 a_n2686_8422.n172 GND 0.005564f
C997 a_n2686_8422.n173 GND 0.01315f
C998 a_n2686_8422.n174 GND 0.005891f
C999 a_n2686_8422.n175 GND 0.045779f
C1000 a_n2686_8422.t7 GND 0.028217f
C1001 a_n2686_8422.n176 GND 0.009863f
C1002 a_n2686_8422.n177 GND 0.008361f
C1003 a_n2686_8422.n178 GND 0.005564f
C1004 a_n2686_8422.n179 GND 0.237506f
C1005 a_n2686_8422.n180 GND 0.010354f
C1006 a_n2686_8422.n181 GND 0.005564f
C1007 a_n2686_8422.n182 GND 0.005891f
C1008 a_n2686_8422.n183 GND 0.01315f
C1009 a_n2686_8422.n184 GND 0.01315f
C1010 a_n2686_8422.n185 GND 0.005891f
C1011 a_n2686_8422.n186 GND 0.005564f
C1012 a_n2686_8422.n187 GND 0.010354f
C1013 a_n2686_8422.n188 GND 0.010354f
C1014 a_n2686_8422.n189 GND 0.005564f
C1015 a_n2686_8422.n190 GND 0.005891f
C1016 a_n2686_8422.n191 GND 0.01315f
C1017 a_n2686_8422.n192 GND 0.031688f
C1018 a_n2686_8422.n193 GND 0.005891f
C1019 a_n2686_8422.n194 GND 0.005564f
C1020 a_n2686_8422.n195 GND 0.023932f
C1021 a_n2686_8422.n196 GND 0.018351f
C1022 a_n2686_8422.n197 GND 0.429985f
C1023 a_n2686_8422.n198 GND 1.24148f
C1024 a_n2686_8422.n199 GND 1.43744f
C1025 a_n2686_8422.n200 GND 0.011333f
C1026 a_n2686_8422.n201 GND 0.010354f
C1027 a_n2686_8422.n202 GND 0.005564f
C1028 a_n2686_8422.n203 GND 0.01315f
C1029 a_n2686_8422.n204 GND 0.005891f
C1030 a_n2686_8422.n205 GND 0.010354f
C1031 a_n2686_8422.n206 GND 0.005564f
C1032 a_n2686_8422.n207 GND 0.01315f
C1033 a_n2686_8422.n208 GND 0.005891f
C1034 a_n2686_8422.n209 GND 0.045779f
C1035 a_n2686_8422.t10 GND 0.028217f
C1036 a_n2686_8422.n210 GND 0.009863f
C1037 a_n2686_8422.n211 GND 0.008361f
C1038 a_n2686_8422.n212 GND 0.005564f
C1039 a_n2686_8422.n213 GND 0.237506f
C1040 a_n2686_8422.n214 GND 0.010354f
C1041 a_n2686_8422.n215 GND 0.005564f
C1042 a_n2686_8422.n216 GND 0.005891f
C1043 a_n2686_8422.n217 GND 0.01315f
C1044 a_n2686_8422.n218 GND 0.01315f
C1045 a_n2686_8422.n219 GND 0.005891f
C1046 a_n2686_8422.n220 GND 0.005564f
C1047 a_n2686_8422.n221 GND 0.010354f
C1048 a_n2686_8422.n222 GND 0.010354f
C1049 a_n2686_8422.n223 GND 0.005564f
C1050 a_n2686_8422.n224 GND 0.005891f
C1051 a_n2686_8422.n225 GND 0.01315f
C1052 a_n2686_8422.n226 GND 0.031688f
C1053 a_n2686_8422.n227 GND 0.005891f
C1054 a_n2686_8422.n228 GND 0.005564f
C1055 a_n2686_8422.n229 GND 0.023932f
C1056 a_n2686_8422.n230 GND 0.018351f
C1057 a_n2686_8422.n231 GND 0.390095f
C1058 a_n2686_8422.n232 GND 0.011333f
C1059 a_n2686_8422.n233 GND 0.010354f
C1060 a_n2686_8422.n234 GND 0.005564f
C1061 a_n2686_8422.n235 GND 0.01315f
C1062 a_n2686_8422.n236 GND 0.005891f
C1063 a_n2686_8422.n237 GND 0.010354f
C1064 a_n2686_8422.n238 GND 0.005564f
C1065 a_n2686_8422.n239 GND 0.01315f
C1066 a_n2686_8422.n240 GND 0.005891f
C1067 a_n2686_8422.n241 GND 0.045779f
C1068 a_n2686_8422.t17 GND 0.028217f
C1069 a_n2686_8422.n242 GND 0.009863f
C1070 a_n2686_8422.n243 GND 0.008361f
C1071 a_n2686_8422.n244 GND 0.005564f
C1072 a_n2686_8422.n245 GND 0.237506f
C1073 a_n2686_8422.n246 GND 0.010354f
C1074 a_n2686_8422.n247 GND 0.005564f
C1075 a_n2686_8422.n248 GND 0.005891f
C1076 a_n2686_8422.n249 GND 0.01315f
C1077 a_n2686_8422.n250 GND 0.01315f
C1078 a_n2686_8422.n251 GND 0.005891f
C1079 a_n2686_8422.n252 GND 0.005564f
C1080 a_n2686_8422.n253 GND 0.010354f
C1081 a_n2686_8422.n254 GND 0.010354f
C1082 a_n2686_8422.n255 GND 0.005564f
C1083 a_n2686_8422.n256 GND 0.005891f
C1084 a_n2686_8422.n257 GND 0.01315f
C1085 a_n2686_8422.n258 GND 0.031688f
C1086 a_n2686_8422.n259 GND 0.005891f
C1087 a_n2686_8422.n260 GND 0.005564f
C1088 a_n2686_8422.n261 GND 0.023932f
C1089 a_n2686_8422.n262 GND 0.019785f
C1090 a_n2686_8422.t11 GND 0.049091f
C1091 a_n2686_8422.t8 GND 0.049091f
C1092 a_n2686_8422.n263 GND 0.302215f
C1093 a_n2686_8422.n264 GND 0.429488f
C1094 a_n2686_8422.n265 GND 0.334913f
C1095 a_n2686_8422.n266 GND 0.302215f
C1096 a_n2686_8422.t19 GND 0.049091f
C1097 a_n2686_12778.n0 GND 0.76359f
C1098 a_n2686_12778.n1 GND 0.354832f
C1099 a_n2686_12778.n2 GND 0.760583f
C1100 a_n2686_12778.n3 GND 0.624142f
C1101 a_n2686_12778.n4 GND 0.354832f
C1102 a_n2686_12778.n5 GND 0.682877f
C1103 a_n2686_12778.n6 GND 0.354832f
C1104 a_n2686_12778.n7 GND 0.727612f
C1105 a_n2686_12778.n8 GND 0.354832f
C1106 a_n2686_12778.n9 GND 0.636545f
C1107 a_n2686_12778.n10 GND 0.354832f
C1108 a_n2686_12778.n11 GND 0.555617f
C1109 a_n2686_12778.n12 GND 0.354832f
C1110 a_n2686_12778.n13 GND 0.054355f
C1111 a_n2686_12778.n14 GND 0.054355f
C1112 a_n2686_12778.n15 GND 0.054355f
C1113 a_n2686_12778.n16 GND 0.045529f
C1114 a_n2686_12778.n17 GND 0.054355f
C1115 a_n2686_12778.n18 GND 0.045529f
C1116 a_n2686_12778.n19 GND 0.054355f
C1117 a_n2686_12778.n20 GND 0.045529f
C1118 a_n2686_12778.n21 GND 0.054355f
C1119 a_n2686_12778.n22 GND 0.07469f
C1120 a_n2686_12778.n23 GND 0.045529f
C1121 a_n2686_12778.n24 GND 0.061824f
C1122 a_n2686_12778.n25 GND 0.092664f
C1123 a_n2686_12778.n26 GND 0.108156f
C1124 a_n2686_12778.n27 GND 0.07469f
C1125 a_n2686_12778.n28 GND 0.045529f
C1126 a_n2686_12778.n29 GND 0.061824f
C1127 a_n2686_12778.n30 GND 0.092664f
C1128 a_n2686_12778.n31 GND 0.108156f
C1129 a_n2686_12778.n32 GND 0.07469f
C1130 a_n2686_12778.n33 GND 0.045529f
C1131 a_n2686_12778.n34 GND 0.061824f
C1132 a_n2686_12778.n35 GND 0.092664f
C1133 a_n2686_12778.n36 GND 0.108156f
C1134 a_n2686_12778.n37 GND 0.07469f
C1135 a_n2686_12778.n38 GND 0.045529f
C1136 a_n2686_12778.n39 GND 0.061824f
C1137 a_n2686_12778.n40 GND 0.092664f
C1138 a_n2686_12778.n41 GND 0.108156f
C1139 a_n2686_12778.n42 GND 0.092664f
C1140 a_n2686_12778.n43 GND 0.061824f
C1141 a_n2686_12778.n44 GND 0.092664f
C1142 a_n2686_12778.n45 GND 0.092664f
C1143 a_n2686_12778.n46 GND 0.092664f
C1144 a_n2686_12778.n47 GND 0.045529f
C1145 a_n2686_12778.n48 GND 0.108156f
C1146 a_n2686_12778.n49 GND 0.054355f
C1147 a_n2686_12778.n50 GND 0.123881f
C1148 a_n2686_12778.n51 GND 0.042225f
C1149 a_n2686_12778.n52 GND 0.036148f
C1150 a_n2686_12778.n53 GND 0.036148f
C1151 a_n2686_12778.n54 GND 0.432684f
C1152 a_n2686_12778.n55 GND 0.036148f
C1153 a_n2686_12778.n56 GND 0.036148f
C1154 a_n2686_12778.n57 GND 0.432684f
C1155 a_n2686_12778.n58 GND 0.036148f
C1156 a_n2686_12778.n59 GND 0.036148f
C1157 a_n2686_12778.n60 GND 0.432684f
C1158 a_n2686_12778.n61 GND 0.036148f
C1159 a_n2686_12778.n62 GND 0.036148f
C1160 a_n2686_12778.n63 GND 0.432684f
C1161 a_n2686_12778.t5 GND 0.09998f
C1162 a_n2686_12778.t37 GND 0.847314f
C1163 a_n2686_12778.t46 GND 0.73578f
C1164 a_n2686_12778.n64 GND 0.400864f
C1165 a_n2686_12778.t43 GND 0.73578f
C1166 a_n2686_12778.t34 GND 0.73578f
C1167 a_n2686_12778.t41 GND 0.73578f
C1168 a_n2686_12778.n65 GND 0.400864f
C1169 a_n2686_12778.t40 GND 0.847314f
C1170 a_n2686_12778.n66 GND 0.019784f
C1171 a_n2686_12778.n67 GND 0.009712f
C1172 a_n2686_12778.n68 GND 0.022956f
C1173 a_n2686_12778.n69 GND 0.010284f
C1174 a_n2686_12778.n70 GND 0.009712f
C1175 a_n2686_12778.n71 GND 0.022956f
C1176 a_n2686_12778.n72 GND 0.010284f
C1177 a_n2686_12778.n73 GND 0.079915f
C1178 a_n2686_12778.t22 GND 0.049258f
C1179 a_n2686_12778.n74 GND 0.017217f
C1180 a_n2686_12778.n75 GND 0.014596f
C1181 a_n2686_12778.n76 GND 0.009712f
C1182 a_n2686_12778.n77 GND 0.009712f
C1183 a_n2686_12778.n78 GND 0.010284f
C1184 a_n2686_12778.n79 GND 0.022956f
C1185 a_n2686_12778.n80 GND 0.022956f
C1186 a_n2686_12778.n81 GND 0.010284f
C1187 a_n2686_12778.n82 GND 0.009712f
C1188 a_n2686_12778.n83 GND 0.009712f
C1189 a_n2686_12778.n84 GND 0.010284f
C1190 a_n2686_12778.n85 GND 0.022956f
C1191 a_n2686_12778.n86 GND 0.055317f
C1192 a_n2686_12778.n87 GND 0.010284f
C1193 a_n2686_12778.n88 GND 0.009712f
C1194 a_n2686_12778.n89 GND 0.041778f
C1195 a_n2686_12778.n90 GND 0.034538f
C1196 a_n2686_12778.t20 GND 0.085697f
C1197 a_n2686_12778.t18 GND 0.085697f
C1198 a_n2686_12778.n91 GND 0.527571f
C1199 a_n2686_12778.n92 GND 0.749749f
C1200 a_n2686_12778.t26 GND 0.085697f
C1201 a_n2686_12778.t14 GND 0.085697f
C1202 a_n2686_12778.n93 GND 0.527571f
C1203 a_n2686_12778.n94 GND 0.584651f
C1204 a_n2686_12778.n95 GND 0.019784f
C1205 a_n2686_12778.n96 GND 0.009712f
C1206 a_n2686_12778.n97 GND 0.022956f
C1207 a_n2686_12778.n98 GND 0.010284f
C1208 a_n2686_12778.n99 GND 0.009712f
C1209 a_n2686_12778.n100 GND 0.022956f
C1210 a_n2686_12778.n101 GND 0.010284f
C1211 a_n2686_12778.n102 GND 0.079915f
C1212 a_n2686_12778.t24 GND 0.049258f
C1213 a_n2686_12778.n103 GND 0.017217f
C1214 a_n2686_12778.n104 GND 0.014596f
C1215 a_n2686_12778.n105 GND 0.009712f
C1216 a_n2686_12778.n106 GND 0.009712f
C1217 a_n2686_12778.n107 GND 0.010284f
C1218 a_n2686_12778.n108 GND 0.022956f
C1219 a_n2686_12778.n109 GND 0.022956f
C1220 a_n2686_12778.n110 GND 0.010284f
C1221 a_n2686_12778.n111 GND 0.009712f
C1222 a_n2686_12778.n112 GND 0.009712f
C1223 a_n2686_12778.n113 GND 0.010284f
C1224 a_n2686_12778.n114 GND 0.022956f
C1225 a_n2686_12778.n115 GND 0.055317f
C1226 a_n2686_12778.n116 GND 0.010284f
C1227 a_n2686_12778.n117 GND 0.009712f
C1228 a_n2686_12778.n118 GND 0.041778f
C1229 a_n2686_12778.n119 GND 0.032035f
C1230 a_n2686_12778.n120 GND 0.697509f
C1231 a_n2686_12778.t56 GND 0.73578f
C1232 a_n2686_12778.t38 GND 0.73578f
C1233 a_n2686_12778.t53 GND 0.806329f
C1234 a_n2686_12778.t52 GND 0.73578f
C1235 a_n2686_12778.t55 GND 0.73578f
C1236 a_n2686_12778.t45 GND 0.806329f
C1237 a_n2686_12778.t51 GND 0.73578f
C1238 a_n2686_12778.t47 GND 0.73578f
C1239 a_n2686_12778.t58 GND 0.806329f
C1240 a_n2686_12778.t59 GND 0.73578f
C1241 a_n2686_12778.t50 GND 0.73578f
C1242 a_n2686_12778.t33 GND 0.806329f
C1243 a_n2686_12778.t49 GND 0.847314f
C1244 a_n2686_12778.t54 GND 0.73578f
C1245 a_n2686_12778.n121 GND 0.400864f
C1246 a_n2686_12778.t32 GND 0.73578f
C1247 a_n2686_12778.t48 GND 0.73578f
C1248 a_n2686_12778.t57 GND 0.73578f
C1249 a_n2686_12778.n122 GND 0.400864f
C1250 a_n2686_12778.t35 GND 0.847314f
C1251 a_n2686_12778.t21 GND 0.847314f
C1252 a_n2686_12778.t19 GND 0.73578f
C1253 a_n2686_12778.n123 GND 0.400864f
C1254 a_n2686_12778.t17 GND 0.73578f
C1255 a_n2686_12778.t25 GND 0.73578f
C1256 a_n2686_12778.t13 GND 0.73578f
C1257 a_n2686_12778.n124 GND 0.400864f
C1258 a_n2686_12778.t23 GND 0.847314f
C1259 a_n2686_12778.n125 GND 0.383422f
C1260 a_n2686_12778.n126 GND 0.07469f
C1261 a_n2686_12778.n127 GND 0.339858f
C1262 a_n2686_12778.n128 GND 0.383422f
C1263 a_n2686_12778.n129 GND 0.07469f
C1264 a_n2686_12778.n130 GND 0.339858f
C1265 a_n2686_12778.t15 GND 0.806329f
C1266 a_n2686_12778.t27 GND 0.73578f
C1267 a_n2686_12778.n131 GND 0.302103f
C1268 a_n2686_12778.t7 GND 0.73578f
C1269 a_n2686_12778.t29 GND 0.73578f
C1270 a_n2686_12778.t9 GND 0.73578f
C1271 a_n2686_12778.n132 GND 0.374076f
C1272 a_n2686_12778.t11 GND 0.806329f
C1273 a_n2686_12778.n133 GND 0.380381f
C1274 a_n2686_12778.n134 GND 0.383422f
C1275 a_n2686_12778.n135 GND 0.07469f
C1276 a_n2686_12778.n136 GND 0.302103f
C1277 a_n2686_12778.n137 GND 0.063608f
C1278 a_n2686_12778.n138 GND 0.056671f
C1279 a_n2686_12778.n139 GND 0.04473f
C1280 a_n2686_12778.n140 GND 0.051421f
C1281 a_n2686_12778.n141 GND 0.370259f
C1282 a_n2686_12778.n142 GND 0.409298f
C1283 a_n2686_12778.n143 GND 0.019784f
C1284 a_n2686_12778.n144 GND 0.009712f
C1285 a_n2686_12778.n145 GND 0.022956f
C1286 a_n2686_12778.n146 GND 0.010284f
C1287 a_n2686_12778.n147 GND 0.009712f
C1288 a_n2686_12778.n148 GND 0.022956f
C1289 a_n2686_12778.n149 GND 0.010284f
C1290 a_n2686_12778.n150 GND 0.079915f
C1291 a_n2686_12778.t12 GND 0.049258f
C1292 a_n2686_12778.n151 GND 0.017217f
C1293 a_n2686_12778.n152 GND 0.014596f
C1294 a_n2686_12778.n153 GND 0.009712f
C1295 a_n2686_12778.n154 GND 0.009712f
C1296 a_n2686_12778.n155 GND 0.010284f
C1297 a_n2686_12778.n156 GND 0.022956f
C1298 a_n2686_12778.n157 GND 0.022956f
C1299 a_n2686_12778.n158 GND 0.010284f
C1300 a_n2686_12778.n159 GND 0.009712f
C1301 a_n2686_12778.n160 GND 0.009712f
C1302 a_n2686_12778.n161 GND 0.010284f
C1303 a_n2686_12778.n162 GND 0.022956f
C1304 a_n2686_12778.n163 GND 0.055317f
C1305 a_n2686_12778.n164 GND 0.010284f
C1306 a_n2686_12778.n165 GND 0.009712f
C1307 a_n2686_12778.n166 GND 0.041778f
C1308 a_n2686_12778.n167 GND 0.034538f
C1309 a_n2686_12778.t30 GND 0.085697f
C1310 a_n2686_12778.t10 GND 0.085697f
C1311 a_n2686_12778.n168 GND 0.527571f
C1312 a_n2686_12778.n169 GND 0.749749f
C1313 a_n2686_12778.t28 GND 0.085697f
C1314 a_n2686_12778.t8 GND 0.085697f
C1315 a_n2686_12778.n170 GND 0.527571f
C1316 a_n2686_12778.n171 GND 0.584651f
C1317 a_n2686_12778.n172 GND 0.019784f
C1318 a_n2686_12778.n173 GND 0.009712f
C1319 a_n2686_12778.n174 GND 0.022956f
C1320 a_n2686_12778.n175 GND 0.010284f
C1321 a_n2686_12778.n176 GND 0.009712f
C1322 a_n2686_12778.n177 GND 0.022956f
C1323 a_n2686_12778.n178 GND 0.010284f
C1324 a_n2686_12778.n179 GND 0.079915f
C1325 a_n2686_12778.t16 GND 0.049258f
C1326 a_n2686_12778.n180 GND 0.017217f
C1327 a_n2686_12778.n181 GND 0.014596f
C1328 a_n2686_12778.n182 GND 0.009712f
C1329 a_n2686_12778.n183 GND 0.009712f
C1330 a_n2686_12778.n184 GND 0.010284f
C1331 a_n2686_12778.n185 GND 0.022956f
C1332 a_n2686_12778.n186 GND 0.022956f
C1333 a_n2686_12778.n187 GND 0.010284f
C1334 a_n2686_12778.n188 GND 0.009712f
C1335 a_n2686_12778.n189 GND 0.009712f
C1336 a_n2686_12778.n190 GND 0.010284f
C1337 a_n2686_12778.n191 GND 0.022956f
C1338 a_n2686_12778.n192 GND 0.055317f
C1339 a_n2686_12778.n193 GND 0.010284f
C1340 a_n2686_12778.n194 GND 0.009712f
C1341 a_n2686_12778.n195 GND 0.041778f
C1342 a_n2686_12778.n196 GND 0.032035f
C1343 a_n2686_12778.n197 GND 0.608786f
C1344 a_n2686_12778.n198 GND 0.543706f
C1345 a_n2686_12778.n199 GND 0.726757f
C1346 a_n2686_12778.n200 GND 0.372726f
C1347 a_n2686_12778.n201 GND 0.373777f
C1348 a_n2686_12778.n202 GND 0.063551f
C1349 a_n2686_12778.n203 GND 0.345667f
C1350 a_n2686_12778.n204 GND 0.302103f
C1351 a_n2686_12778.n205 GND 0.063551f
C1352 a_n2686_12778.t42 GND 0.806329f
C1353 a_n2686_12778.n206 GND 0.373777f
C1354 a_n2686_12778.n207 GND 0.121163f
C1355 a_n2686_12778.n208 GND 0.121163f
C1356 a_n2686_12778.n209 GND 0.373777f
C1357 a_n2686_12778.n210 GND 0.063551f
C1358 a_n2686_12778.n211 GND 0.345667f
C1359 a_n2686_12778.n212 GND 0.302103f
C1360 a_n2686_12778.n213 GND 0.063551f
C1361 a_n2686_12778.t39 GND 0.806329f
C1362 a_n2686_12778.n214 GND 0.373777f
C1363 a_n2686_12778.n215 GND 0.156013f
C1364 a_n2686_12778.n216 GND 0.156013f
C1365 a_n2686_12778.n217 GND 0.373777f
C1366 a_n2686_12778.n218 GND 0.063551f
C1367 a_n2686_12778.n219 GND 0.345667f
C1368 a_n2686_12778.n220 GND 0.302103f
C1369 a_n2686_12778.n221 GND 0.063551f
C1370 a_n2686_12778.t36 GND 0.806329f
C1371 a_n2686_12778.n222 GND 0.373777f
C1372 a_n2686_12778.n223 GND 0.121163f
C1373 a_n2686_12778.n224 GND 0.121163f
C1374 a_n2686_12778.n225 GND 0.373777f
C1375 a_n2686_12778.n226 GND 0.063551f
C1376 a_n2686_12778.n227 GND 0.345667f
C1377 a_n2686_12778.n228 GND 0.302103f
C1378 a_n2686_12778.n229 GND 0.063551f
C1379 a_n2686_12778.t44 GND 0.806329f
C1380 a_n2686_12778.n230 GND 0.373777f
C1381 a_n2686_12778.n231 GND 0.372726f
C1382 a_n2686_12778.n232 GND 0.925215f
C1383 a_n2686_12778.n233 GND 0.383422f
C1384 a_n2686_12778.n234 GND 0.07469f
C1385 a_n2686_12778.n235 GND 0.339858f
C1386 a_n2686_12778.n236 GND 2.67653f
C1387 a_n2686_12778.t31 GND 0.09998f
C1388 a_n2686_12778.t1 GND 0.09998f
C1389 a_n2686_12778.n237 GND 0.884701f
C1390 a_n2686_12778.t4 GND 0.09998f
C1391 a_n2686_12778.t6 GND 0.09998f
C1392 a_n2686_12778.n238 GND 0.884701f
C1393 a_n2686_12778.n239 GND 2.22521f
C1394 a_n2686_12778.t2 GND 0.09998f
C1395 a_n2686_12778.t3 GND 0.09998f
C1396 a_n2686_12778.n240 GND 0.883454f
C1397 a_n2686_12778.n241 GND 2.09477f
C1398 a_n2686_12778.n242 GND 2.82663f
C1399 a_n2686_12778.n243 GND 0.884703f
C1400 a_n2686_12778.t0 GND 0.09998f
C1401 VDD.t29 GND 0.021143f
C1402 VDD.t21 GND 0.021143f
C1403 VDD.n0 GND 0.152771f
C1404 VDD.t24 GND 0.021143f
C1405 VDD.t35 GND 0.021143f
C1406 VDD.n1 GND 0.15206f
C1407 VDD.n2 GND 0.276787f
C1408 VDD.t19 GND 0.021143f
C1409 VDD.t31 GND 0.021143f
C1410 VDD.n3 GND 0.15206f
C1411 VDD.n4 GND 0.141412f
C1412 VDD.t3 GND 0.021143f
C1413 VDD.t17 GND 0.021143f
C1414 VDD.n5 GND 0.15206f
C1415 VDD.n6 GND 0.128034f
C1416 VDD.t15 GND 0.021143f
C1417 VDD.t199 GND 0.021143f
C1418 VDD.n7 GND 0.152771f
C1419 VDD.t38 GND 0.021143f
C1420 VDD.t10 GND 0.021143f
C1421 VDD.n8 GND 0.15206f
C1422 VDD.n9 GND 0.276787f
C1423 VDD.t12 GND 0.021143f
C1424 VDD.t196 GND 0.021143f
C1425 VDD.n10 GND 0.15206f
C1426 VDD.n11 GND 0.141412f
C1427 VDD.t6 GND 0.021143f
C1428 VDD.t27 GND 0.021143f
C1429 VDD.n12 GND 0.15206f
C1430 VDD.n13 GND 0.128034f
C1431 VDD.n14 GND 0.084873f
C1432 VDD.n15 GND 2.1359f
C1433 VDD.t155 GND 0.2147f
C1434 VDD.t164 GND 0.024667f
C1435 VDD.t144 GND 0.024667f
C1436 VDD.n16 GND 0.158313f
C1437 VDD.n17 GND 0.280774f
C1438 VDD.t166 GND 0.024667f
C1439 VDD.t168 GND 0.024667f
C1440 VDD.n18 GND 0.158313f
C1441 VDD.n19 GND 0.149623f
C1442 VDD.t151 GND 0.024667f
C1443 VDD.t129 GND 0.024667f
C1444 VDD.n20 GND 0.158313f
C1445 VDD.n21 GND 0.149623f
C1446 VDD.t175 GND 0.024667f
C1447 VDD.t163 GND 0.024667f
C1448 VDD.n22 GND 0.158313f
C1449 VDD.n23 GND 0.149623f
C1450 VDD.t146 GND 0.213746f
C1451 VDD.n24 GND 0.196646f
C1452 VDD.t167 GND 0.2147f
C1453 VDD.t171 GND 0.024667f
C1454 VDD.t190 GND 0.024667f
C1455 VDD.n25 GND 0.158313f
C1456 VDD.n26 GND 0.280774f
C1457 VDD.t181 GND 0.024667f
C1458 VDD.t183 GND 0.024667f
C1459 VDD.n27 GND 0.158313f
C1460 VDD.n28 GND 0.149623f
C1461 VDD.t131 GND 0.024667f
C1462 VDD.t173 GND 0.024667f
C1463 VDD.n29 GND 0.158313f
C1464 VDD.n30 GND 0.149623f
C1465 VDD.t116 GND 0.024667f
C1466 VDD.t161 GND 0.024667f
C1467 VDD.n31 GND 0.158313f
C1468 VDD.n32 GND 0.149623f
C1469 VDD.t184 GND 0.213746f
C1470 VDD.n33 GND 0.156865f
C1471 VDD.n34 GND 0.332902f
C1472 VDD.t192 GND 0.2147f
C1473 VDD.t118 GND 0.024667f
C1474 VDD.t162 GND 0.024667f
C1475 VDD.n35 GND 0.158313f
C1476 VDD.n36 GND 0.280774f
C1477 VDD.t140 GND 0.024667f
C1478 VDD.t150 GND 0.024667f
C1479 VDD.n37 GND 0.158313f
C1480 VDD.n38 GND 0.149623f
C1481 VDD.t176 GND 0.024667f
C1482 VDD.t124 GND 0.024667f
C1483 VDD.n39 GND 0.158313f
C1484 VDD.n40 GND 0.149623f
C1485 VDD.t170 GND 0.024667f
C1486 VDD.t188 GND 0.024667f
C1487 VDD.n41 GND 0.158313f
C1488 VDD.n42 GND 0.149623f
C1489 VDD.t152 GND 0.213746f
C1490 VDD.n43 GND 0.156865f
C1491 VDD.n44 GND 0.30242f
C1492 VDD.n45 GND 0.00673f
C1493 VDD.n46 GND 0.008756f
C1494 VDD.n47 GND 0.007048f
C1495 VDD.n48 GND 0.007048f
C1496 VDD.n49 GND 0.008756f
C1497 VDD.n50 GND 0.008756f
C1498 VDD.n51 GND 0.642906f
C1499 VDD.n52 GND 0.008756f
C1500 VDD.n53 GND 0.008756f
C1501 VDD.n54 GND 0.008756f
C1502 VDD.n55 GND 0.523459f
C1503 VDD.n56 GND 0.008756f
C1504 VDD.n57 GND 0.008756f
C1505 VDD.n58 GND 0.008756f
C1506 VDD.n59 GND 0.008756f
C1507 VDD.n60 GND 0.007048f
C1508 VDD.n61 GND 0.008756f
C1509 VDD.t123 GND 0.351315f
C1510 VDD.n62 GND 0.008756f
C1511 VDD.n63 GND 0.008756f
C1512 VDD.n64 GND 0.008756f
C1513 VDD.t115 GND 0.351315f
C1514 VDD.n65 GND 0.008756f
C1515 VDD.n66 GND 0.008756f
C1516 VDD.n67 GND 0.008756f
C1517 VDD.n68 GND 0.008756f
C1518 VDD.n69 GND 0.008756f
C1519 VDD.n70 GND 0.007048f
C1520 VDD.n71 GND 0.008756f
C1521 VDD.n72 GND 0.649932f
C1522 VDD.n73 GND 0.008756f
C1523 VDD.n74 GND 0.008756f
C1524 VDD.n75 GND 0.008756f
C1525 VDD.n76 GND 0.516432f
C1526 VDD.n77 GND 0.008756f
C1527 VDD.n78 GND 0.008756f
C1528 VDD.n79 GND 0.008756f
C1529 VDD.n80 GND 0.008756f
C1530 VDD.n81 GND 0.008756f
C1531 VDD.n82 GND 0.007048f
C1532 VDD.n83 GND 0.008756f
C1533 VDD.t145 GND 0.351315f
C1534 VDD.n84 GND 0.008756f
C1535 VDD.n85 GND 0.008756f
C1536 VDD.n86 GND 0.008756f
C1537 VDD.n87 GND 0.702629f
C1538 VDD.n88 GND 0.008756f
C1539 VDD.n89 GND 0.008756f
C1540 VDD.n90 GND 0.008756f
C1541 VDD.n91 GND 0.008756f
C1542 VDD.n92 GND 0.008756f
C1543 VDD.n93 GND 0.007048f
C1544 VDD.n94 GND 0.008756f
C1545 VDD.n95 GND 0.008756f
C1546 VDD.n96 GND 0.008756f
C1547 VDD.n97 GND 0.019672f
C1548 VDD.n98 GND 1.52822f
C1549 VDD.n99 GND 0.01973f
C1550 VDD.n100 GND 0.008756f
C1551 VDD.n101 GND 0.008756f
C1552 VDD.n103 GND 0.008756f
C1553 VDD.n104 GND 0.008756f
C1554 VDD.n105 GND 0.007048f
C1555 VDD.n106 GND 0.007048f
C1556 VDD.n107 GND 0.008756f
C1557 VDD.n108 GND 0.008756f
C1558 VDD.n109 GND 0.008756f
C1559 VDD.n110 GND 0.008756f
C1560 VDD.n111 GND 0.008756f
C1561 VDD.n112 GND 0.008756f
C1562 VDD.n113 GND 0.007048f
C1563 VDD.n115 GND 0.008756f
C1564 VDD.n116 GND 0.008756f
C1565 VDD.n117 GND 0.008756f
C1566 VDD.n118 GND 0.008756f
C1567 VDD.n119 GND 0.008756f
C1568 VDD.n120 GND 0.007048f
C1569 VDD.n122 GND 0.008756f
C1570 VDD.n123 GND 0.008756f
C1571 VDD.n124 GND 0.008756f
C1572 VDD.n125 GND 0.008756f
C1573 VDD.n126 GND 0.008756f
C1574 VDD.n127 GND 0.005885f
C1575 VDD.n129 GND 0.008756f
C1576 VDD.n130 GND 0.005885f
C1577 VDD.t108 GND 0.17936f
C1578 VDD.t107 GND 0.187962f
C1579 VDD.t106 GND 0.262044f
C1580 VDD.n131 GND 0.088819f
C1581 VDD.n132 GND 0.050925f
C1582 VDD.n133 GND 0.008756f
C1583 VDD.n134 GND 0.008756f
C1584 VDD.n135 GND 0.007048f
C1585 VDD.n137 GND 0.008756f
C1586 VDD.n138 GND 0.008756f
C1587 VDD.n139 GND 0.008756f
C1588 VDD.n140 GND 0.008756f
C1589 VDD.n141 GND 0.007048f
C1590 VDD.n143 GND 0.008756f
C1591 VDD.n144 GND 0.008756f
C1592 VDD.n145 GND 0.008756f
C1593 VDD.n146 GND 0.008756f
C1594 VDD.n147 GND 0.008756f
C1595 VDD.n148 GND 0.007048f
C1596 VDD.n150 GND 0.008756f
C1597 VDD.n151 GND 0.008756f
C1598 VDD.n152 GND 0.008756f
C1599 VDD.n153 GND 0.008756f
C1600 VDD.n154 GND 0.008756f
C1601 VDD.n155 GND 0.007048f
C1602 VDD.n157 GND 0.008756f
C1603 VDD.n158 GND 0.008756f
C1604 VDD.n159 GND 0.008756f
C1605 VDD.n160 GND 0.008756f
C1606 VDD.n161 GND 0.008756f
C1607 VDD.n162 GND 0.004792f
C1608 VDD.n164 GND 0.008756f
C1609 VDD.n165 GND 0.006977f
C1610 VDD.t76 GND 0.17936f
C1611 VDD.t75 GND 0.187962f
C1612 VDD.t74 GND 0.262044f
C1613 VDD.n166 GND 0.088819f
C1614 VDD.n167 GND 0.050925f
C1615 VDD.n168 GND 0.008756f
C1616 VDD.n169 GND 0.008756f
C1617 VDD.n170 GND 0.007048f
C1618 VDD.n172 GND 0.008756f
C1619 VDD.n173 GND 0.008756f
C1620 VDD.n174 GND 0.008756f
C1621 VDD.n175 GND 0.008756f
C1622 VDD.n176 GND 0.007048f
C1623 VDD.n178 GND 0.008756f
C1624 VDD.n179 GND 0.008756f
C1625 VDD.n180 GND 0.008756f
C1626 VDD.n181 GND 0.008756f
C1627 VDD.n182 GND 0.008756f
C1628 VDD.n183 GND 0.007048f
C1629 VDD.n185 GND 0.008756f
C1630 VDD.n186 GND 0.008756f
C1631 VDD.n187 GND 0.008756f
C1632 VDD.n188 GND 0.008756f
C1633 VDD.n189 GND 0.008756f
C1634 VDD.n190 GND 0.007048f
C1635 VDD.n192 GND 0.008756f
C1636 VDD.n193 GND 0.008756f
C1637 VDD.n194 GND 0.008756f
C1638 VDD.n195 GND 0.008756f
C1639 VDD.n196 GND 0.008756f
C1640 VDD.n197 GND 0.0037f
C1641 VDD.t65 GND 0.17936f
C1642 VDD.t64 GND 0.187962f
C1643 VDD.t62 GND 0.262044f
C1644 VDD.n199 GND 0.088819f
C1645 VDD.n200 GND 0.050925f
C1646 VDD.n201 GND 0.010889f
C1647 VDD.n202 GND 0.008756f
C1648 VDD.n203 GND 0.008756f
C1649 VDD.n204 GND 0.008756f
C1650 VDD.n205 GND 0.007048f
C1651 VDD.n206 GND 0.008756f
C1652 VDD.n207 GND 0.008756f
C1653 VDD.n208 GND 0.007048f
C1654 VDD.n209 GND 0.008756f
C1655 VDD.n210 GND 0.008756f
C1656 VDD.n211 GND 0.007048f
C1657 VDD.n212 GND 0.008756f
C1658 VDD.n213 GND 0.008756f
C1659 VDD.n214 GND 0.007048f
C1660 VDD.n215 GND 0.008756f
C1661 VDD.n216 GND 0.007048f
C1662 VDD.n217 GND 0.008756f
C1663 VDD.n218 GND 0.007048f
C1664 VDD.n219 GND 0.008756f
C1665 VDD.n220 GND 0.008756f
C1666 VDD.n221 GND 0.702629f
C1667 VDD.t149 GND 0.351315f
C1668 VDD.n222 GND 0.008756f
C1669 VDD.n223 GND 0.007048f
C1670 VDD.n224 GND 0.008756f
C1671 VDD.n225 GND 0.007048f
C1672 VDD.n226 GND 0.008756f
C1673 VDD.t139 GND 0.351315f
C1674 VDD.n227 GND 0.008756f
C1675 VDD.n228 GND 0.007048f
C1676 VDD.n229 GND 0.008756f
C1677 VDD.n230 GND 0.007048f
C1678 VDD.n231 GND 0.008756f
C1679 VDD.n232 GND 0.404012f
C1680 VDD.n233 GND 0.530485f
C1681 VDD.n234 GND 0.008756f
C1682 VDD.n235 GND 0.007048f
C1683 VDD.n236 GND 0.008756f
C1684 VDD.n237 GND 0.007048f
C1685 VDD.n238 GND 0.008756f
C1686 VDD.n239 GND 0.635879f
C1687 VDD.n240 GND 0.008756f
C1688 VDD.n241 GND 0.007048f
C1689 VDD.n242 GND 0.008756f
C1690 VDD.n243 GND 0.007048f
C1691 VDD.n244 GND 0.008756f
C1692 VDD.n245 GND 0.702629f
C1693 VDD.t117 GND 0.351315f
C1694 VDD.n246 GND 0.008756f
C1695 VDD.n247 GND 0.007048f
C1696 VDD.n248 GND 0.008756f
C1697 VDD.n249 GND 0.007048f
C1698 VDD.n250 GND 0.008756f
C1699 VDD.t154 GND 0.351315f
C1700 VDD.n251 GND 0.008756f
C1701 VDD.n252 GND 0.007048f
C1702 VDD.n253 GND 0.008756f
C1703 VDD.n254 GND 0.007048f
C1704 VDD.n255 GND 0.008756f
C1705 VDD.n256 GND 0.702629f
C1706 VDD.n257 GND 0.537511f
C1707 VDD.n258 GND 0.008756f
C1708 VDD.n259 GND 0.007048f
C1709 VDD.n260 GND 0.008756f
C1710 VDD.n261 GND 0.007048f
C1711 VDD.n262 GND 0.008756f
C1712 VDD.n263 GND 0.460222f
C1713 VDD.n264 GND 0.008756f
C1714 VDD.n265 GND 0.007048f
C1715 VDD.n266 GND 0.019672f
C1716 VDD.n267 GND 0.00585f
C1717 VDD.n268 GND 0.019672f
C1718 VDD.n269 GND 0.902878f
C1719 VDD.t71 GND 0.351315f
C1720 VDD.n270 GND 0.019672f
C1721 VDD.n271 GND 0.00585f
C1722 VDD.n272 GND 0.008756f
C1723 VDD.n273 GND 0.007048f
C1724 VDD.n274 GND 0.008756f
C1725 VDD.n275 GND 4.11038f
C1726 VDD.n303 GND 0.01973f
C1727 VDD.n304 GND 0.008756f
C1728 VDD.n305 GND 0.008756f
C1729 VDD.n306 GND 0.008756f
C1730 VDD.n307 GND 0.00753f
C1731 VDD.n308 GND 0.007048f
C1732 VDD.n309 GND 0.005604f
C1733 VDD.n310 GND 0.008306f
C1734 VDD.n311 GND 0.008756f
C1735 VDD.n312 GND 0.008756f
C1736 VDD.n313 GND 0.007048f
C1737 VDD.n314 GND 0.008756f
C1738 VDD.n315 GND 0.008756f
C1739 VDD.n316 GND 0.008756f
C1740 VDD.n317 GND 0.008756f
C1741 VDD.n318 GND 0.008756f
C1742 VDD.n319 GND 0.008756f
C1743 VDD.n320 GND 0.008756f
C1744 VDD.n321 GND 0.008756f
C1745 VDD.n322 GND 0.005885f
C1746 VDD.n323 GND 0.008756f
C1747 VDD.n324 GND 0.008756f
C1748 VDD.n325 GND 0.008756f
C1749 VDD.n326 GND 0.008756f
C1750 VDD.n327 GND 0.008756f
C1751 VDD.n328 GND 0.008756f
C1752 VDD.n329 GND 0.008756f
C1753 VDD.n330 GND 0.008756f
C1754 VDD.n331 GND 0.008756f
C1755 VDD.n332 GND 0.008756f
C1756 VDD.n333 GND 0.008756f
C1757 VDD.n334 GND 0.008756f
C1758 VDD.n335 GND 0.008756f
C1759 VDD.n336 GND 0.008756f
C1760 VDD.n337 GND 0.008756f
C1761 VDD.n338 GND 0.008756f
C1762 VDD.n339 GND 0.008756f
C1763 VDD.n340 GND 0.006977f
C1764 VDD.t113 GND 0.17936f
C1765 VDD.t114 GND 0.187962f
C1766 VDD.t112 GND 0.262044f
C1767 VDD.n341 GND 0.088819f
C1768 VDD.n342 GND 0.050925f
C1769 VDD.n343 GND 0.008756f
C1770 VDD.n344 GND 0.008756f
C1771 VDD.n345 GND 0.008756f
C1772 VDD.n346 GND 0.008756f
C1773 VDD.n347 GND 0.008756f
C1774 VDD.n348 GND 0.008756f
C1775 VDD.n349 GND 0.008756f
C1776 VDD.n350 GND 0.008756f
C1777 VDD.n351 GND 0.005604f
C1778 VDD.n352 GND 0.007048f
C1779 VDD.n353 GND 0.00753f
C1780 VDD.n354 GND 0.004466f
C1781 VDD.n355 GND 0.005954f
C1782 VDD.n357 GND 0.005954f
C1783 VDD.n358 GND 0.005954f
C1784 VDD.n360 GND 0.005954f
C1785 VDD.n361 GND 0.004597f
C1786 VDD.n363 GND 0.005954f
C1787 VDD.t95 GND 0.076127f
C1788 VDD.t94 GND 0.086562f
C1789 VDD.t93 GND 0.227136f
C1790 VDD.n364 GND 0.151662f
C1791 VDD.n365 GND 0.122136f
C1792 VDD.n366 GND 0.008509f
C1793 VDD.n367 GND 0.013956f
C1794 VDD.n369 GND 0.005954f
C1795 VDD.n370 GND 0.477788f
C1796 VDD.n371 GND 0.013224f
C1797 VDD.n372 GND 0.013224f
C1798 VDD.n373 GND 0.005954f
C1799 VDD.n374 GND 0.01392f
C1800 VDD.n375 GND 0.005954f
C1801 VDD.n376 GND 0.005954f
C1802 VDD.n378 GND 0.005954f
C1803 VDD.n379 GND 0.005954f
C1804 VDD.n381 GND 0.005954f
C1805 VDD.n382 GND 0.005954f
C1806 VDD.n384 GND 0.005954f
C1807 VDD.n385 GND 0.005954f
C1808 VDD.n387 GND 0.005954f
C1809 VDD.n388 GND 0.005954f
C1810 VDD.n390 GND 0.005954f
C1811 VDD.t54 GND 0.076127f
C1812 VDD.t53 GND 0.086562f
C1813 VDD.t51 GND 0.227136f
C1814 VDD.n391 GND 0.151662f
C1815 VDD.n392 GND 0.122136f
C1816 VDD.n393 GND 0.005954f
C1817 VDD.n395 GND 0.005954f
C1818 VDD.n396 GND 0.005954f
C1819 VDD.n397 GND 0.263486f
C1820 VDD.n398 GND 0.005954f
C1821 VDD.n399 GND 0.005954f
C1822 VDD.n400 GND 0.005954f
C1823 VDD.n401 GND 0.005954f
C1824 VDD.n402 GND 0.005954f
C1825 VDD.n403 GND 0.400499f
C1826 VDD.n404 GND 0.005954f
C1827 VDD.n405 GND 0.005954f
C1828 VDD.t52 GND 0.238894f
C1829 VDD.n406 GND 0.005954f
C1830 VDD.n407 GND 0.005954f
C1831 VDD.t104 GND 0.086562f
C1832 VDD.t102 GND 0.227136f
C1833 VDD.t105 GND 0.086562f
C1834 VDD.n408 GND 0.274428f
C1835 VDD.n409 GND 0.005954f
C1836 VDD.n410 GND 0.005954f
C1837 VDD.n411 GND 0.477788f
C1838 VDD.n412 GND 0.005954f
C1839 VDD.n413 GND 0.005954f
C1840 VDD.t103 GND 0.238894f
C1841 VDD.n414 GND 0.005954f
C1842 VDD.n415 GND 0.005954f
C1843 VDD.n416 GND 0.005954f
C1844 VDD.n417 GND 0.477788f
C1845 VDD.n418 GND 0.005954f
C1846 VDD.n419 GND 0.005954f
C1847 VDD.n420 GND 0.005954f
C1848 VDD.n421 GND 0.005954f
C1849 VDD.n422 GND 0.005954f
C1850 VDD.t0 GND 0.238894f
C1851 VDD.n423 GND 0.005954f
C1852 VDD.n424 GND 0.005954f
C1853 VDD.n425 GND 0.005954f
C1854 VDD.n426 GND 0.005954f
C1855 VDD.n427 GND 0.005954f
C1856 VDD.t198 GND 0.238894f
C1857 VDD.n428 GND 0.005954f
C1858 VDD.n429 GND 0.005954f
C1859 VDD.n430 GND 0.425091f
C1860 VDD.n431 GND 0.005954f
C1861 VDD.n432 GND 0.005954f
C1862 VDD.n433 GND 0.005954f
C1863 VDD.t197 GND 0.238894f
C1864 VDD.n434 GND 0.005954f
C1865 VDD.n435 GND 0.005954f
C1866 VDD.n436 GND 0.288078f
C1867 VDD.n437 GND 0.005954f
C1868 VDD.n438 GND 0.005954f
C1869 VDD.n439 GND 0.005954f
C1870 VDD.t14 GND 0.238894f
C1871 VDD.n440 GND 0.005954f
C1872 VDD.n441 GND 0.005954f
C1873 VDD.n442 GND 0.446169f
C1874 VDD.n443 GND 0.005954f
C1875 VDD.n444 GND 0.005954f
C1876 VDD.n445 GND 0.005954f
C1877 VDD.t36 GND 0.238894f
C1878 VDD.n446 GND 0.005954f
C1879 VDD.n447 GND 0.005954f
C1880 VDD.n448 GND 0.309157f
C1881 VDD.n449 GND 0.005954f
C1882 VDD.n450 GND 0.005954f
C1883 VDD.n451 GND 0.005954f
C1884 VDD.t9 GND 0.238894f
C1885 VDD.n452 GND 0.005954f
C1886 VDD.n453 GND 0.005954f
C1887 VDD.n454 GND 0.467248f
C1888 VDD.n455 GND 0.005954f
C1889 VDD.n456 GND 0.005954f
C1890 VDD.n457 GND 0.005954f
C1891 VDD.n458 GND 0.477788f
C1892 VDD.n459 GND 0.005954f
C1893 VDD.n460 GND 0.005954f
C1894 VDD.t1 GND 0.238894f
C1895 VDD.n461 GND 0.005954f
C1896 VDD.n462 GND 0.005954f
C1897 VDD.n463 GND 0.005954f
C1898 VDD.t37 GND 0.238894f
C1899 VDD.n464 GND 0.005954f
C1900 VDD.n465 GND 0.005954f
C1901 VDD.n466 GND 0.005954f
C1902 VDD.n467 GND 0.005954f
C1903 VDD.n468 GND 0.005954f
C1904 VDD.n469 GND 0.477788f
C1905 VDD.n470 GND 0.005954f
C1906 VDD.n471 GND 0.005954f
C1907 VDD.t8 GND 0.238894f
C1908 VDD.n472 GND 0.005954f
C1909 VDD.n473 GND 0.005954f
C1910 VDD.n474 GND 0.005954f
C1911 VDD.n475 GND 0.425091f
C1912 VDD.n476 GND 0.005954f
C1913 VDD.n477 GND 0.005954f
C1914 VDD.n478 GND 0.005954f
C1915 VDD.n479 GND 0.005954f
C1916 VDD.n480 GND 0.005954f
C1917 VDD.t195 GND 0.238894f
C1918 VDD.n481 GND 0.005954f
C1919 VDD.n482 GND 0.005954f
C1920 VDD.t33 GND 0.238894f
C1921 VDD.n483 GND 0.005954f
C1922 VDD.n484 GND 0.005954f
C1923 VDD.n485 GND 0.005954f
C1924 VDD.n486 GND 0.477788f
C1925 VDD.n487 GND 0.005954f
C1926 VDD.n488 GND 0.005954f
C1927 VDD.n489 GND 0.344288f
C1928 VDD.n490 GND 0.005954f
C1929 VDD.n491 GND 0.005954f
C1930 VDD.n492 GND 0.005954f
C1931 VDD.t11 GND 0.238894f
C1932 VDD.n493 GND 0.005954f
C1933 VDD.n494 GND 0.005954f
C1934 VDD.n495 GND 0.005954f
C1935 VDD.n496 GND 0.005954f
C1936 VDD.n497 GND 0.005954f
C1937 VDD.t59 GND 0.238894f
C1938 VDD.n498 GND 0.005954f
C1939 VDD.n499 GND 0.005954f
C1940 VDD.n500 GND 0.365367f
C1941 VDD.n501 GND 0.005954f
C1942 VDD.n502 GND 0.005954f
C1943 VDD.n503 GND 0.005954f
C1944 VDD.t26 GND 0.238894f
C1945 VDD.n504 GND 0.005954f
C1946 VDD.n505 GND 0.005954f
C1947 VDD.n506 GND 0.263486f
C1948 VDD.n507 GND 0.005954f
C1949 VDD.n508 GND 0.01392f
C1950 VDD.n509 GND 0.01392f
C1951 VDD.n510 GND 0.660471f
C1952 VDD.n536 GND 0.01392f
C1953 VDD.n537 GND 0.013224f
C1954 VDD.n538 GND 0.005954f
C1955 VDD.n539 GND 0.013224f
C1956 VDD.t111 GND 0.076127f
C1957 VDD.t110 GND 0.086562f
C1958 VDD.t109 GND 0.227136f
C1959 VDD.n540 GND 0.151662f
C1960 VDD.n541 GND 0.122136f
C1961 VDD.n542 GND 0.008509f
C1962 VDD.n543 GND 0.005954f
C1963 VDD.n544 GND 0.005954f
C1964 VDD.t2 GND 0.238894f
C1965 VDD.n545 GND 0.005954f
C1966 VDD.n546 GND 0.005954f
C1967 VDD.n547 GND 0.005954f
C1968 VDD.n548 GND 0.013224f
C1969 VDD.n549 GND 0.005954f
C1970 VDD.t89 GND 0.076127f
C1971 VDD.t88 GND 0.086562f
C1972 VDD.t86 GND 0.227136f
C1973 VDD.n550 GND 0.151662f
C1974 VDD.n551 GND 0.122136f
C1975 VDD.n552 GND 0.005954f
C1976 VDD.n553 GND 0.005954f
C1977 VDD.n554 GND 0.263486f
C1978 VDD.n555 GND 0.005954f
C1979 VDD.n556 GND 0.005954f
C1980 VDD.n557 GND 0.005954f
C1981 VDD.n558 GND 0.365367f
C1982 VDD.n559 GND 0.005954f
C1983 VDD.n560 GND 0.005954f
C1984 VDD.t87 GND 0.238894f
C1985 VDD.n561 GND 0.005954f
C1986 VDD.n562 GND 0.005954f
C1987 VDD.n563 GND 0.005954f
C1988 VDD.n564 GND 0.005954f
C1989 VDD.n565 GND 0.477788f
C1990 VDD.n566 GND 0.005954f
C1991 VDD.n567 GND 0.005954f
C1992 VDD.t30 GND 0.238894f
C1993 VDD.n568 GND 0.005954f
C1994 VDD.n569 GND 0.005954f
C1995 VDD.n570 GND 0.005954f
C1996 VDD.n571 GND 0.344288f
C1997 VDD.n572 GND 0.005954f
C1998 VDD.n573 GND 0.005954f
C1999 VDD.n574 GND 0.005954f
C2000 VDD.n575 GND 0.005954f
C2001 VDD.n576 GND 0.005954f
C2002 VDD.t7 GND 0.238894f
C2003 VDD.n577 GND 0.005954f
C2004 VDD.n578 GND 0.005954f
C2005 VDD.t18 GND 0.238894f
C2006 VDD.n579 GND 0.005954f
C2007 VDD.n580 GND 0.005954f
C2008 VDD.n581 GND 0.005954f
C2009 VDD.n582 GND 0.477788f
C2010 VDD.n583 GND 0.005954f
C2011 VDD.n584 GND 0.005954f
C2012 VDD.n585 GND 0.425091f
C2013 VDD.n586 GND 0.005954f
C2014 VDD.n587 GND 0.005954f
C2015 VDD.n588 GND 0.005954f
C2016 VDD.t13 GND 0.238894f
C2017 VDD.n589 GND 0.005954f
C2018 VDD.n590 GND 0.005954f
C2019 VDD.n591 GND 0.005954f
C2020 VDD.n592 GND 0.005954f
C2021 VDD.n593 GND 0.005954f
C2022 VDD.n594 GND 0.477788f
C2023 VDD.n595 GND 0.005954f
C2024 VDD.n596 GND 0.005954f
C2025 VDD.t34 GND 0.238894f
C2026 VDD.n597 GND 0.005954f
C2027 VDD.n598 GND 0.005954f
C2028 VDD.n599 GND 0.005954f
C2029 VDD.t32 GND 0.238894f
C2030 VDD.n600 GND 0.005954f
C2031 VDD.n601 GND 0.005954f
C2032 VDD.n602 GND 0.005954f
C2033 VDD.n603 GND 0.005954f
C2034 VDD.n604 GND 0.005954f
C2035 VDD.n605 GND 0.467248f
C2036 VDD.n606 GND 0.005954f
C2037 VDD.n607 GND 0.005954f
C2038 VDD.t23 GND 0.238894f
C2039 VDD.n608 GND 0.005954f
C2040 VDD.n609 GND 0.005954f
C2041 VDD.n610 GND 0.005954f
C2042 VDD.n611 GND 0.309157f
C2043 VDD.n612 GND 0.005954f
C2044 VDD.n613 GND 0.005954f
C2045 VDD.t4 GND 0.238894f
C2046 VDD.n614 GND 0.005954f
C2047 VDD.n615 GND 0.005954f
C2048 VDD.n616 GND 0.005954f
C2049 VDD.n617 GND 0.446169f
C2050 VDD.n618 GND 0.005954f
C2051 VDD.n619 GND 0.005954f
C2052 VDD.t20 GND 0.238894f
C2053 VDD.n620 GND 0.005954f
C2054 VDD.n621 GND 0.005954f
C2055 VDD.n622 GND 0.005954f
C2056 VDD.n623 GND 0.288078f
C2057 VDD.n624 GND 0.005954f
C2058 VDD.n625 GND 0.005954f
C2059 VDD.t22 GND 0.238894f
C2060 VDD.n626 GND 0.005954f
C2061 VDD.n627 GND 0.005954f
C2062 VDD.n628 GND 0.005954f
C2063 VDD.n629 GND 0.425091f
C2064 VDD.n630 GND 0.005954f
C2065 VDD.n631 GND 0.005954f
C2066 VDD.t28 GND 0.238894f
C2067 VDD.n632 GND 0.005954f
C2068 VDD.n633 GND 0.005954f
C2069 VDD.n634 GND 0.005954f
C2070 VDD.n635 GND 0.477788f
C2071 VDD.n636 GND 0.005954f
C2072 VDD.n637 GND 0.005954f
C2073 VDD.t25 GND 0.238894f
C2074 VDD.n638 GND 0.005954f
C2075 VDD.n639 GND 0.005954f
C2076 VDD.n640 GND 0.005954f
C2077 VDD.n641 GND 0.477788f
C2078 VDD.n642 GND 0.005954f
C2079 VDD.n643 GND 0.005954f
C2080 VDD.n644 GND 0.005954f
C2081 VDD.n645 GND 0.005954f
C2082 VDD.n646 GND 0.005954f
C2083 VDD.t48 GND 0.238894f
C2084 VDD.n647 GND 0.005954f
C2085 VDD.n648 GND 0.005954f
C2086 VDD.n649 GND 0.005954f
C2087 VDD.t49 GND 0.086562f
C2088 VDD.t47 GND 0.227136f
C2089 VDD.t50 GND 0.086562f
C2090 VDD.n650 GND 0.274428f
C2091 VDD.n651 GND 0.005954f
C2092 VDD.n652 GND 0.005954f
C2093 VDD.t67 GND 0.238894f
C2094 VDD.n653 GND 0.005954f
C2095 VDD.n654 GND 0.005954f
C2096 VDD.n655 GND 0.400499f
C2097 VDD.n656 GND 0.005954f
C2098 VDD.n657 GND 0.005954f
C2099 VDD.n658 GND 0.005954f
C2100 VDD.n659 GND 0.477788f
C2101 VDD.n660 GND 0.005954f
C2102 VDD.n661 GND 0.005954f
C2103 VDD.n662 GND 0.263486f
C2104 VDD.n663 GND 0.005954f
C2105 VDD.n664 GND 0.01392f
C2106 VDD.n665 GND 0.01392f
C2107 VDD.n666 GND 4.11038f
C2108 VDD.n667 GND 0.013224f
C2109 VDD.n668 GND 0.013224f
C2110 VDD.n669 GND 0.01392f
C2111 VDD.n670 GND 0.005954f
C2112 VDD.n672 GND 0.005954f
C2113 VDD.n673 GND 0.005954f
C2114 VDD.n674 GND 0.005954f
C2115 VDD.n675 GND 0.005954f
C2116 VDD.n676 GND 0.011781f
C2117 VDD.n678 GND 0.005954f
C2118 VDD.n679 GND 0.005954f
C2119 VDD.n680 GND 0.005954f
C2120 VDD.n681 GND 0.005954f
C2121 VDD.t68 GND 0.076127f
C2122 VDD.t69 GND 0.086562f
C2123 VDD.t66 GND 0.227136f
C2124 VDD.n682 GND 0.151662f
C2125 VDD.n683 GND 0.122136f
C2126 VDD.n684 GND 0.008509f
C2127 VDD.n686 GND 0.005954f
C2128 VDD.n687 GND 0.005954f
C2129 VDD.n688 GND 0.005954f
C2130 VDD.t97 GND 0.076127f
C2131 VDD.t98 GND 0.086562f
C2132 VDD.t96 GND 0.227136f
C2133 VDD.n689 GND 0.151662f
C2134 VDD.n690 GND 0.122136f
C2135 VDD.n691 GND 0.005954f
C2136 VDD.n692 GND 0.005954f
C2137 VDD.n693 GND 0.005954f
C2138 VDD.n694 GND 0.005954f
C2139 VDD.n695 GND 0.005604f
C2140 VDD.n698 GND 0.008756f
C2141 VDD.n699 GND 0.007048f
C2142 VDD.n700 GND 0.008756f
C2143 VDD.n701 GND 0.008756f
C2144 VDD.n702 GND 0.008756f
C2145 VDD.n703 GND 0.0037f
C2146 VDD.n704 GND 0.019672f
C2147 VDD.t46 GND 0.17936f
C2148 VDD.t45 GND 0.187962f
C2149 VDD.t43 GND 0.262044f
C2150 VDD.n705 GND 0.088819f
C2151 VDD.n706 GND 0.050925f
C2152 VDD.n707 GND 0.010889f
C2153 VDD.n708 GND 0.008756f
C2154 VDD.n710 GND 0.008756f
C2155 VDD.n711 GND 0.00585f
C2156 VDD.n712 GND 0.593722f
C2157 VDD.n714 GND 4.24037f
C2158 VDD.n715 GND 0.008756f
C2159 VDD.n716 GND 0.01973f
C2160 VDD.n717 GND 0.007048f
C2161 VDD.n718 GND 0.008756f
C2162 VDD.n719 GND 0.007048f
C2163 VDD.n720 GND 0.008756f
C2164 VDD.n721 GND 0.702629f
C2165 VDD.n722 GND 0.008756f
C2166 VDD.n723 GND 0.007048f
C2167 VDD.n724 GND 0.007048f
C2168 VDD.n725 GND 0.008756f
C2169 VDD.n726 GND 0.007048f
C2170 VDD.n727 GND 0.008756f
C2171 VDD.n728 GND 0.702629f
C2172 VDD.n729 GND 0.008756f
C2173 VDD.n730 GND 0.007048f
C2174 VDD.n731 GND 0.008756f
C2175 VDD.n732 GND 0.007048f
C2176 VDD.n733 GND 0.008756f
C2177 VDD.t125 GND 0.351315f
C2178 VDD.n734 GND 0.008756f
C2179 VDD.n735 GND 0.007048f
C2180 VDD.n736 GND 0.008756f
C2181 VDD.n737 GND 0.007048f
C2182 VDD.n738 GND 0.008756f
C2183 VDD.n739 GND 0.418064f
C2184 VDD.n740 GND 0.516432f
C2185 VDD.n741 GND 0.008756f
C2186 VDD.n742 GND 0.007048f
C2187 VDD.n743 GND 0.008756f
C2188 VDD.n744 GND 0.007048f
C2189 VDD.n745 GND 0.008756f
C2190 VDD.n746 GND 0.649932f
C2191 VDD.n747 GND 0.008756f
C2192 VDD.n748 GND 0.007048f
C2193 VDD.n749 GND 0.008756f
C2194 VDD.n750 GND 0.007048f
C2195 VDD.n751 GND 0.008756f
C2196 VDD.n752 GND 0.702629f
C2197 VDD.t137 GND 0.351315f
C2198 VDD.n753 GND 0.008756f
C2199 VDD.n754 GND 0.007048f
C2200 VDD.n755 GND 0.008756f
C2201 VDD.n756 GND 0.007048f
C2202 VDD.n757 GND 0.008756f
C2203 VDD.t158 GND 0.351315f
C2204 VDD.n758 GND 0.008756f
C2205 VDD.n759 GND 0.007048f
C2206 VDD.n760 GND 0.008756f
C2207 VDD.n761 GND 0.007048f
C2208 VDD.n762 GND 0.008756f
C2209 VDD.n763 GND 0.411038f
C2210 VDD.n764 GND 0.523459f
C2211 VDD.n765 GND 0.008756f
C2212 VDD.n766 GND 0.007048f
C2213 VDD.t126 GND 0.2147f
C2214 VDD.t193 GND 0.024667f
C2215 VDD.t136 GND 0.024667f
C2216 VDD.n767 GND 0.158313f
C2217 VDD.n768 GND 0.280774f
C2218 VDD.t148 GND 0.024667f
C2219 VDD.t169 GND 0.024667f
C2220 VDD.n769 GND 0.158313f
C2221 VDD.n770 GND 0.149623f
C2222 VDD.t189 GND 0.024667f
C2223 VDD.t120 GND 0.024667f
C2224 VDD.n771 GND 0.158313f
C2225 VDD.n772 GND 0.149623f
C2226 VDD.t134 GND 0.024667f
C2227 VDD.t179 GND 0.024667f
C2228 VDD.n773 GND 0.158313f
C2229 VDD.n774 GND 0.149623f
C2230 VDD.t194 GND 0.213746f
C2231 VDD.n775 GND 0.196646f
C2232 VDD.t182 GND 0.2147f
C2233 VDD.t138 GND 0.024667f
C2234 VDD.t185 GND 0.024667f
C2235 VDD.n776 GND 0.158313f
C2236 VDD.n777 GND 0.280774f
C2237 VDD.t122 GND 0.024667f
C2238 VDD.t187 GND 0.024667f
C2239 VDD.n778 GND 0.158313f
C2240 VDD.n779 GND 0.149623f
C2241 VDD.t186 GND 0.024667f
C2242 VDD.t165 GND 0.024667f
C2243 VDD.n780 GND 0.158313f
C2244 VDD.n781 GND 0.149623f
C2245 VDD.t177 GND 0.024667f
C2246 VDD.t142 GND 0.024667f
C2247 VDD.n782 GND 0.158313f
C2248 VDD.n783 GND 0.149623f
C2249 VDD.t128 GND 0.213746f
C2250 VDD.n784 GND 0.156865f
C2251 VDD.n785 GND 0.332902f
C2252 VDD.t147 GND 0.2147f
C2253 VDD.t178 GND 0.024667f
C2254 VDD.t153 GND 0.024667f
C2255 VDD.n786 GND 0.158313f
C2256 VDD.n787 GND 0.280774f
C2257 VDD.t172 GND 0.024667f
C2258 VDD.t159 GND 0.024667f
C2259 VDD.n788 GND 0.158313f
C2260 VDD.n789 GND 0.149623f
C2261 VDD.t157 GND 0.024667f
C2262 VDD.t191 GND 0.024667f
C2263 VDD.n790 GND 0.158313f
C2264 VDD.n791 GND 0.149623f
C2265 VDD.t133 GND 0.024667f
C2266 VDD.t180 GND 0.024667f
C2267 VDD.n792 GND 0.158313f
C2268 VDD.n793 GND 0.149623f
C2269 VDD.t174 GND 0.213746f
C2270 VDD.n794 GND 0.156865f
C2271 VDD.n795 GND 0.30242f
C2272 VDD.n796 GND 1.81635f
C2273 VDD.n797 GND 0.238982f
C2274 VDD.n798 GND 0.007048f
C2275 VDD.n799 GND 0.008756f
C2276 VDD.n800 GND 0.642906f
C2277 VDD.n801 GND 0.008756f
C2278 VDD.n802 GND 0.007048f
C2279 VDD.n803 GND 0.008756f
C2280 VDD.n804 GND 0.007048f
C2281 VDD.n805 GND 0.008756f
C2282 VDD.n806 GND 0.702629f
C2283 VDD.t119 GND 0.351315f
C2284 VDD.n807 GND 0.008756f
C2285 VDD.n808 GND 0.007048f
C2286 VDD.n809 GND 0.008756f
C2287 VDD.n810 GND 0.007048f
C2288 VDD.n811 GND 0.008756f
C2289 VDD.t156 GND 0.351315f
C2290 VDD.n812 GND 0.008756f
C2291 VDD.n813 GND 0.007048f
C2292 VDD.n814 GND 0.008756f
C2293 VDD.n815 GND 0.007048f
C2294 VDD.n816 GND 0.008756f
C2295 VDD.n817 GND 0.404012f
C2296 VDD.n818 GND 0.530485f
C2297 VDD.n819 GND 0.008756f
C2298 VDD.n820 GND 0.007048f
C2299 VDD.n821 GND 0.008756f
C2300 VDD.n822 GND 0.007048f
C2301 VDD.n823 GND 0.008756f
C2302 VDD.n824 GND 0.635879f
C2303 VDD.n825 GND 0.008756f
C2304 VDD.n826 GND 0.007048f
C2305 VDD.n827 GND 0.008756f
C2306 VDD.n828 GND 0.007048f
C2307 VDD.n829 GND 0.008756f
C2308 VDD.n830 GND 0.702629f
C2309 VDD.t132 GND 0.351315f
C2310 VDD.n831 GND 0.008756f
C2311 VDD.n832 GND 0.007048f
C2312 VDD.n833 GND 0.008756f
C2313 VDD.n834 GND 0.007048f
C2314 VDD.n835 GND 0.008756f
C2315 VDD.t127 GND 0.351315f
C2316 VDD.n836 GND 0.008756f
C2317 VDD.n837 GND 0.007048f
C2318 VDD.n838 GND 0.008756f
C2319 VDD.n839 GND 0.007048f
C2320 VDD.n840 GND 0.008756f
C2321 VDD.n841 GND 0.702629f
C2322 VDD.n842 GND 0.537511f
C2323 VDD.n843 GND 0.008756f
C2324 VDD.n844 GND 0.007048f
C2325 VDD.n845 GND 0.008756f
C2326 VDD.n846 GND 0.007048f
C2327 VDD.n847 GND 0.008756f
C2328 VDD.n848 GND 0.460222f
C2329 VDD.n849 GND 0.008756f
C2330 VDD.n850 GND 0.007048f
C2331 VDD.n851 GND 0.019672f
C2332 VDD.n852 GND 0.00585f
C2333 VDD.n853 GND 0.019672f
C2334 VDD.n854 GND 0.902878f
C2335 VDD.t40 GND 0.351315f
C2336 VDD.n855 GND 0.019672f
C2337 VDD.n856 GND 0.00585f
C2338 VDD.n857 GND 0.008756f
C2339 VDD.n858 GND 0.007048f
C2340 VDD.n859 GND 0.008756f
C2341 VDD.n887 GND 0.01973f
C2342 VDD.n888 GND 0.008756f
C2343 VDD.n889 GND 0.007048f
C2344 VDD.n890 GND 0.008756f
C2345 VDD.n891 GND 0.008756f
C2346 VDD.n892 GND 0.008756f
C2347 VDD.n893 GND 0.008756f
C2348 VDD.n894 GND 0.008756f
C2349 VDD.n895 GND 0.007048f
C2350 VDD.n896 GND 0.008756f
C2351 VDD.n897 GND 0.008756f
C2352 VDD.n898 GND 0.008756f
C2353 VDD.n899 GND 0.008756f
C2354 VDD.n900 GND 0.008756f
C2355 VDD.n901 GND 0.007048f
C2356 VDD.n902 GND 0.008756f
C2357 VDD.n903 GND 0.008756f
C2358 VDD.n904 GND 0.008756f
C2359 VDD.n905 GND 0.008756f
C2360 VDD.n906 GND 0.008756f
C2361 VDD.n907 GND 0.007048f
C2362 VDD.n908 GND 0.008756f
C2363 VDD.n909 GND 0.008756f
C2364 VDD.n910 GND 0.008756f
C2365 VDD.n911 GND 0.008756f
C2366 VDD.n912 GND 0.007048f
C2367 VDD.n913 GND 0.008756f
C2368 VDD.n914 GND 0.008756f
C2369 VDD.n915 GND 0.008756f
C2370 VDD.n916 GND 0.008756f
C2371 VDD.n917 GND 0.008756f
C2372 VDD.n918 GND 0.007048f
C2373 VDD.n919 GND 0.008756f
C2374 VDD.n920 GND 0.008756f
C2375 VDD.n921 GND 0.008756f
C2376 VDD.n922 GND 0.008756f
C2377 VDD.n923 GND 0.008756f
C2378 VDD.n924 GND 0.007048f
C2379 VDD.n925 GND 0.008756f
C2380 VDD.n926 GND 0.008756f
C2381 VDD.n927 GND 0.008756f
C2382 VDD.n928 GND 0.008756f
C2383 VDD.n929 GND 0.008756f
C2384 VDD.n930 GND 0.007048f
C2385 VDD.n931 GND 0.008756f
C2386 VDD.n932 GND 0.008756f
C2387 VDD.n933 GND 0.008756f
C2388 VDD.n934 GND 0.008756f
C2389 VDD.n935 GND 0.008756f
C2390 VDD.n936 GND 0.007048f
C2391 VDD.n937 GND 0.008756f
C2392 VDD.n938 GND 0.008756f
C2393 VDD.n939 GND 0.008756f
C2394 VDD.n940 GND 0.008756f
C2395 VDD.n941 GND 0.007048f
C2396 VDD.n942 GND 0.008756f
C2397 VDD.n943 GND 0.008756f
C2398 VDD.n944 GND 0.008756f
C2399 VDD.n945 GND 0.008756f
C2400 VDD.n946 GND 0.008756f
C2401 VDD.n947 GND 0.007048f
C2402 VDD.n948 GND 0.008756f
C2403 VDD.n949 GND 0.008756f
C2404 VDD.n950 GND 0.008756f
C2405 VDD.n951 GND 0.008756f
C2406 VDD.n952 GND 0.008756f
C2407 VDD.n953 GND 0.007048f
C2408 VDD.n954 GND 0.008756f
C2409 VDD.n955 GND 0.008756f
C2410 VDD.n956 GND 0.008756f
C2411 VDD.n957 GND 0.008756f
C2412 VDD.n958 GND 0.008756f
C2413 VDD.n959 GND 0.007048f
C2414 VDD.n960 GND 0.008756f
C2415 VDD.n961 GND 0.008756f
C2416 VDD.n962 GND 0.008756f
C2417 VDD.n963 GND 0.008756f
C2418 VDD.n964 GND 0.008756f
C2419 VDD.n965 GND 0.007048f
C2420 VDD.n966 GND 0.01973f
C2421 VDD.n967 GND 0.008756f
C2422 VDD.n968 GND 0.003348f
C2423 VDD.t78 GND 0.17936f
C2424 VDD.t79 GND 0.187962f
C2425 VDD.t77 GND 0.262044f
C2426 VDD.n969 GND 0.088819f
C2427 VDD.n970 GND 0.050925f
C2428 VDD.n971 GND 0.010889f
C2429 VDD.n972 GND 0.0037f
C2430 VDD.n973 GND 0.008756f
C2431 VDD.n974 GND 0.008756f
C2432 VDD.n975 GND 0.008756f
C2433 VDD.n976 GND 0.007048f
C2434 VDD.n977 GND 0.007048f
C2435 VDD.n978 GND 0.007048f
C2436 VDD.n979 GND 0.008756f
C2437 VDD.n980 GND 0.008756f
C2438 VDD.n981 GND 0.008756f
C2439 VDD.n982 GND 0.007048f
C2440 VDD.n983 GND 0.007048f
C2441 VDD.n984 GND 0.007048f
C2442 VDD.n985 GND 0.008756f
C2443 VDD.n986 GND 0.008756f
C2444 VDD.n987 GND 0.008756f
C2445 VDD.n988 GND 0.007048f
C2446 VDD.n989 GND 0.007048f
C2447 VDD.n990 GND 0.007048f
C2448 VDD.n991 GND 0.008756f
C2449 VDD.n992 GND 0.008756f
C2450 VDD.n993 GND 0.008756f
C2451 VDD.n994 GND 0.007048f
C2452 VDD.n995 GND 0.007048f
C2453 VDD.n996 GND 0.007048f
C2454 VDD.n997 GND 0.008756f
C2455 VDD.n998 GND 0.008756f
C2456 VDD.n999 GND 0.008756f
C2457 VDD.n1000 GND 0.006977f
C2458 VDD.n1001 GND 0.008756f
C2459 VDD.t91 GND 0.17936f
C2460 VDD.t92 GND 0.187962f
C2461 VDD.t90 GND 0.262044f
C2462 VDD.n1002 GND 0.088819f
C2463 VDD.n1003 GND 0.050925f
C2464 VDD.n1004 GND 0.014412f
C2465 VDD.n1005 GND 0.004792f
C2466 VDD.n1006 GND 0.008756f
C2467 VDD.n1007 GND 0.008756f
C2468 VDD.n1008 GND 0.008756f
C2469 VDD.n1009 GND 0.007048f
C2470 VDD.n1010 GND 0.007048f
C2471 VDD.n1011 GND 0.007048f
C2472 VDD.n1012 GND 0.008756f
C2473 VDD.n1013 GND 0.008756f
C2474 VDD.n1014 GND 0.008756f
C2475 VDD.n1015 GND 0.007048f
C2476 VDD.n1016 GND 0.007048f
C2477 VDD.n1017 GND 0.007048f
C2478 VDD.n1018 GND 0.008756f
C2479 VDD.n1019 GND 0.008756f
C2480 VDD.n1020 GND 0.008756f
C2481 VDD.n1021 GND 0.007048f
C2482 VDD.n1022 GND 0.007048f
C2483 VDD.n1023 GND 0.007048f
C2484 VDD.n1024 GND 0.008756f
C2485 VDD.n1025 GND 0.008756f
C2486 VDD.n1026 GND 0.008756f
C2487 VDD.n1027 GND 0.007048f
C2488 VDD.n1028 GND 0.007048f
C2489 VDD.n1029 GND 0.007048f
C2490 VDD.n1030 GND 0.008756f
C2491 VDD.n1031 GND 0.008756f
C2492 VDD.n1032 GND 0.008756f
C2493 VDD.n1033 GND 0.005885f
C2494 VDD.n1034 GND 0.008756f
C2495 VDD.t41 GND 0.17936f
C2496 VDD.t42 GND 0.187962f
C2497 VDD.t39 GND 0.262044f
C2498 VDD.n1035 GND 0.088819f
C2499 VDD.n1036 GND 0.050925f
C2500 VDD.n1037 GND 0.014412f
C2501 VDD.n1038 GND 0.005885f
C2502 VDD.n1039 GND 0.008756f
C2503 VDD.n1040 GND 0.008756f
C2504 VDD.n1041 GND 0.008756f
C2505 VDD.n1042 GND 0.007048f
C2506 VDD.n1043 GND 0.007048f
C2507 VDD.n1044 GND 0.007048f
C2508 VDD.n1045 GND 0.008756f
C2509 VDD.n1046 GND 0.008756f
C2510 VDD.n1047 GND 0.008756f
C2511 VDD.n1048 GND 0.007048f
C2512 VDD.n1049 GND 0.007048f
C2513 VDD.n1050 GND 0.007048f
C2514 VDD.n1051 GND 0.008756f
C2515 VDD.n1052 GND 0.008756f
C2516 VDD.n1053 GND 0.008756f
C2517 VDD.n1054 GND 0.007048f
C2518 VDD.n1055 GND 0.007048f
C2519 VDD.n1056 GND 0.007048f
C2520 VDD.n1057 GND 0.008756f
C2521 VDD.n1058 GND 0.008756f
C2522 VDD.n1059 GND 0.008756f
C2523 VDD.n1060 GND 0.007048f
C2524 VDD.n1061 GND 0.008756f
C2525 VDD.n1062 GND 1.52822f
C2526 VDD.n1064 GND 0.01973f
C2527 VDD.n1065 GND 0.00585f
C2528 VDD.n1066 GND 0.01973f
C2529 VDD.n1067 GND 0.019672f
C2530 VDD.n1068 GND 0.008756f
C2531 VDD.n1069 GND 0.007048f
C2532 VDD.n1070 GND 0.008756f
C2533 VDD.n1071 GND 0.593722f
C2534 VDD.n1072 GND 0.008756f
C2535 VDD.n1073 GND 0.007048f
C2536 VDD.n1074 GND 0.008756f
C2537 VDD.n1075 GND 0.008756f
C2538 VDD.n1076 GND 0.008756f
C2539 VDD.n1077 GND 0.007048f
C2540 VDD.n1078 GND 0.008756f
C2541 VDD.n1079 GND 0.702629f
C2542 VDD.n1080 GND 0.008756f
C2543 VDD.n1081 GND 0.007048f
C2544 VDD.n1082 GND 0.008756f
C2545 VDD.n1083 GND 0.008756f
C2546 VDD.n1084 GND 0.008756f
C2547 VDD.n1085 GND 0.007048f
C2548 VDD.n1086 GND 0.008756f
C2549 VDD.n1087 GND 0.702629f
C2550 VDD.n1088 GND 0.008756f
C2551 VDD.n1089 GND 0.007048f
C2552 VDD.n1090 GND 0.008756f
C2553 VDD.n1091 GND 0.008756f
C2554 VDD.n1092 GND 0.008756f
C2555 VDD.n1093 GND 0.007048f
C2556 VDD.n1094 GND 0.008756f
C2557 VDD.n1095 GND 0.516432f
C2558 VDD.n1096 GND 0.008756f
C2559 VDD.n1097 GND 0.007048f
C2560 VDD.n1098 GND 0.008756f
C2561 VDD.n1099 GND 0.008756f
C2562 VDD.n1100 GND 0.008756f
C2563 VDD.n1101 GND 0.007048f
C2564 VDD.n1102 GND 0.008756f
C2565 VDD.n1103 GND 0.418064f
C2566 VDD.n1104 GND 0.008756f
C2567 VDD.n1105 GND 0.007048f
C2568 VDD.n1106 GND 0.008756f
C2569 VDD.n1107 GND 0.008756f
C2570 VDD.n1108 GND 0.008756f
C2571 VDD.n1109 GND 0.007048f
C2572 VDD.n1110 GND 0.008756f
C2573 VDD.t141 GND 0.351315f
C2574 VDD.n1111 GND 0.649932f
C2575 VDD.n1112 GND 0.008756f
C2576 VDD.n1113 GND 0.007048f
C2577 VDD.n1114 GND 0.008756f
C2578 VDD.n1115 GND 0.008756f
C2579 VDD.n1116 GND 0.008756f
C2580 VDD.n1117 GND 0.007048f
C2581 VDD.n1118 GND 0.008756f
C2582 VDD.n1119 GND 0.702629f
C2583 VDD.n1120 GND 0.008756f
C2584 VDD.n1121 GND 0.007048f
C2585 VDD.n1122 GND 0.008756f
C2586 VDD.n1123 GND 0.008756f
C2587 VDD.n1124 GND 0.008756f
C2588 VDD.n1125 GND 0.007048f
C2589 VDD.n1126 GND 0.008756f
C2590 VDD.n1127 GND 0.523459f
C2591 VDD.n1128 GND 0.008756f
C2592 VDD.n1129 GND 0.007048f
C2593 VDD.n1130 GND 0.008756f
C2594 VDD.n1131 GND 0.008756f
C2595 VDD.n1132 GND 0.00673f
C2596 VDD.n1133 GND 0.008756f
C2597 VDD.n1134 GND 0.007048f
C2598 VDD.n1135 GND 0.008756f
C2599 VDD.n1136 GND 0.411038f
C2600 VDD.n1137 GND 0.008756f
C2601 VDD.n1138 GND 0.007048f
C2602 VDD.n1139 GND 0.008756f
C2603 VDD.n1140 GND 0.008756f
C2604 VDD.n1141 GND 0.008756f
C2605 VDD.n1142 GND 0.007048f
C2606 VDD.n1143 GND 0.008756f
C2607 VDD.t121 GND 0.351315f
C2608 VDD.n1144 GND 0.642906f
C2609 VDD.n1145 GND 0.008756f
C2610 VDD.n1146 GND 0.007048f
C2611 VDD.n1147 GND 0.00673f
C2612 VDD.n1148 GND 0.008756f
C2613 VDD.n1149 GND 0.008756f
C2614 VDD.n1150 GND 0.007048f
C2615 VDD.n1151 GND 0.008756f
C2616 VDD.n1152 GND 0.702629f
C2617 VDD.n1153 GND 0.008756f
C2618 VDD.n1154 GND 0.007048f
C2619 VDD.n1155 GND 0.008756f
C2620 VDD.n1156 GND 0.008756f
C2621 VDD.n1157 GND 0.008756f
C2622 VDD.n1158 GND 0.007048f
C2623 VDD.n1159 GND 0.008756f
C2624 VDD.n1160 GND 0.530485f
C2625 VDD.n1161 GND 0.008756f
C2626 VDD.n1162 GND 0.007048f
C2627 VDD.n1163 GND 0.008756f
C2628 VDD.n1164 GND 0.008756f
C2629 VDD.n1165 GND 0.008756f
C2630 VDD.n1166 GND 0.007048f
C2631 VDD.n1167 GND 0.008756f
C2632 VDD.n1168 GND 0.404012f
C2633 VDD.n1169 GND 0.008756f
C2634 VDD.n1170 GND 0.007048f
C2635 VDD.n1171 GND 0.008756f
C2636 VDD.n1172 GND 0.008756f
C2637 VDD.n1173 GND 0.008756f
C2638 VDD.n1174 GND 0.007048f
C2639 VDD.n1175 GND 0.008756f
C2640 VDD.t135 GND 0.351315f
C2641 VDD.n1176 GND 0.635879f
C2642 VDD.n1177 GND 0.008756f
C2643 VDD.n1178 GND 0.007048f
C2644 VDD.n1179 GND 0.008756f
C2645 VDD.n1180 GND 0.008756f
C2646 VDD.n1181 GND 0.008756f
C2647 VDD.n1182 GND 0.007048f
C2648 VDD.n1183 GND 0.008756f
C2649 VDD.n1184 GND 0.702629f
C2650 VDD.n1185 GND 0.008756f
C2651 VDD.n1186 GND 0.007048f
C2652 VDD.n1187 GND 0.008756f
C2653 VDD.n1188 GND 0.008756f
C2654 VDD.n1189 GND 0.008756f
C2655 VDD.n1190 GND 0.007048f
C2656 VDD.n1191 GND 0.008756f
C2657 VDD.n1192 GND 0.537511f
C2658 VDD.n1193 GND 0.008756f
C2659 VDD.n1194 GND 0.007048f
C2660 VDD.n1195 GND 0.008756f
C2661 VDD.n1196 GND 0.008756f
C2662 VDD.n1197 GND 0.008756f
C2663 VDD.n1198 GND 0.007048f
C2664 VDD.n1199 GND 0.008756f
C2665 VDD.n1200 GND 0.702629f
C2666 VDD.n1201 GND 0.008756f
C2667 VDD.n1202 GND 0.007048f
C2668 VDD.n1203 GND 0.008756f
C2669 VDD.n1204 GND 0.008756f
C2670 VDD.n1205 GND 0.008756f
C2671 VDD.n1206 GND 0.008756f
C2672 VDD.n1207 GND 0.007048f
C2673 VDD.n1208 GND 0.008756f
C2674 VDD.t44 GND 0.351315f
C2675 VDD.n1209 GND 0.460222f
C2676 VDD.n1210 GND 0.008756f
C2677 VDD.n1211 GND 0.007048f
C2678 VDD.n1212 GND 0.008756f
C2679 VDD.n1213 GND 0.008756f
C2680 VDD.n1214 GND 0.008756f
C2681 VDD.n1215 GND 0.007048f
C2682 VDD.n1217 GND 0.008756f
C2683 VDD.n1218 GND 0.008756f
C2684 VDD.n1219 GND 0.008756f
C2685 VDD.n1220 GND 0.00753f
C2686 VDD.n1222 GND 0.008756f
C2687 VDD.n1223 GND 0.007048f
C2688 VDD.n1224 GND 0.005604f
C2689 VDD.n1225 GND 0.007048f
C2690 VDD.n1226 GND 0.008756f
C2691 VDD.n1228 GND 0.008756f
C2692 VDD.n1229 GND 0.008756f
C2693 VDD.n1230 GND 0.008756f
C2694 VDD.n1231 GND 0.007048f
C2695 VDD.n1233 GND 0.008756f
C2696 VDD.n1234 GND 0.008756f
C2697 VDD.n1235 GND 0.008756f
C2698 VDD.n1236 GND 0.008756f
C2699 VDD.n1237 GND 0.008756f
C2700 VDD.n1238 GND 0.005885f
C2701 VDD.n1240 GND 0.008756f
C2702 VDD.n1241 GND 0.005885f
C2703 VDD.t101 GND 0.17936f
C2704 VDD.t100 GND 0.187962f
C2705 VDD.t99 GND 0.262044f
C2706 VDD.n1242 GND 0.088819f
C2707 VDD.n1243 GND 0.050925f
C2708 VDD.n1244 GND 0.008756f
C2709 VDD.n1245 GND 0.008756f
C2710 VDD.n1246 GND 0.007048f
C2711 VDD.n1248 GND 0.008756f
C2712 VDD.n1249 GND 0.008756f
C2713 VDD.n1250 GND 0.008756f
C2714 VDD.n1251 GND 0.008756f
C2715 VDD.n1252 GND 0.007048f
C2716 VDD.n1254 GND 0.008756f
C2717 VDD.n1255 GND 0.008756f
C2718 VDD.n1256 GND 0.008756f
C2719 VDD.n1257 GND 0.008756f
C2720 VDD.n1258 GND 0.008756f
C2721 VDD.n1259 GND 0.007048f
C2722 VDD.n1261 GND 0.008756f
C2723 VDD.n1262 GND 0.008756f
C2724 VDD.n1263 GND 0.008756f
C2725 VDD.n1264 GND 0.008756f
C2726 VDD.n1265 GND 0.008756f
C2727 VDD.n1266 GND 0.007048f
C2728 VDD.n1268 GND 0.008756f
C2729 VDD.n1269 GND 0.008756f
C2730 VDD.n1270 GND 0.008756f
C2731 VDD.n1271 GND 0.008756f
C2732 VDD.n1272 GND 0.008756f
C2733 VDD.n1273 GND 0.004792f
C2734 VDD.n1275 GND 0.008756f
C2735 VDD.n1276 GND 0.006977f
C2736 VDD.t57 GND 0.17936f
C2737 VDD.t56 GND 0.187962f
C2738 VDD.t55 GND 0.262044f
C2739 VDD.n1277 GND 0.088819f
C2740 VDD.n1278 GND 0.050925f
C2741 VDD.n1279 GND 0.008756f
C2742 VDD.n1280 GND 0.008756f
C2743 VDD.n1281 GND 0.007048f
C2744 VDD.n1283 GND 0.008756f
C2745 VDD.n1284 GND 0.008756f
C2746 VDD.n1285 GND 0.008756f
C2747 VDD.n1286 GND 0.008756f
C2748 VDD.n1287 GND 0.007048f
C2749 VDD.n1289 GND 0.008756f
C2750 VDD.n1290 GND 0.008756f
C2751 VDD.n1291 GND 0.008756f
C2752 VDD.n1292 GND 0.008756f
C2753 VDD.n1293 GND 0.008756f
C2754 VDD.n1294 GND 0.007048f
C2755 VDD.n1296 GND 0.007048f
C2756 VDD.n1298 GND 0.008756f
C2757 VDD.n1299 GND 0.007048f
C2758 VDD.n1300 GND 0.008756f
C2759 VDD.n1302 GND 0.008756f
C2760 VDD.n1303 GND 0.007048f
C2761 VDD.n1304 GND 0.008756f
C2762 VDD.n1306 GND 0.008756f
C2763 VDD.n1307 GND 0.008756f
C2764 VDD.n1308 GND 0.007048f
C2765 VDD.n1309 GND 0.007048f
C2766 VDD.n1310 GND 0.007048f
C2767 VDD.n1311 GND 0.008756f
C2768 VDD.n1313 GND 0.008756f
C2769 VDD.n1314 GND 0.008756f
C2770 VDD.n1315 GND 0.007048f
C2771 VDD.n1316 GND 0.007048f
C2772 VDD.n1317 GND 0.007048f
C2773 VDD.n1318 GND 0.008756f
C2774 VDD.n1320 GND 0.008756f
C2775 VDD.n1321 GND 0.008756f
C2776 VDD.n1322 GND 0.007048f
C2777 VDD.n1323 GND 0.008756f
C2778 VDD.n1324 GND 0.008756f
C2779 VDD.n1325 GND 0.008756f
C2780 VDD.n1326 GND 0.014412f
C2781 VDD.n1327 GND 0.008756f
C2782 VDD.n1329 GND 0.008756f
C2783 VDD.n1330 GND 0.008756f
C2784 VDD.n1331 GND 0.007048f
C2785 VDD.n1332 GND 0.007048f
C2786 VDD.n1333 GND 0.007048f
C2787 VDD.n1334 GND 0.008756f
C2788 VDD.n1336 GND 0.008756f
C2789 VDD.n1337 GND 0.008756f
C2790 VDD.n1338 GND 0.007048f
C2791 VDD.n1339 GND 0.007048f
C2792 VDD.n1340 GND 0.007048f
C2793 VDD.n1341 GND 0.008756f
C2794 VDD.n1343 GND 0.008756f
C2795 VDD.n1344 GND 0.008756f
C2796 VDD.n1345 GND 0.007048f
C2797 VDD.n1346 GND 0.007048f
C2798 VDD.n1347 GND 0.007048f
C2799 VDD.n1348 GND 0.008756f
C2800 VDD.n1350 GND 0.008756f
C2801 VDD.n1351 GND 0.008756f
C2802 VDD.n1352 GND 0.007048f
C2803 VDD.n1353 GND 0.007048f
C2804 VDD.n1354 GND 0.007048f
C2805 VDD.n1355 GND 0.008756f
C2806 VDD.n1357 GND 0.008756f
C2807 VDD.n1358 GND 0.008756f
C2808 VDD.n1359 GND 0.007048f
C2809 VDD.n1360 GND 0.008756f
C2810 VDD.n1361 GND 0.008756f
C2811 VDD.n1362 GND 0.008756f
C2812 VDD.n1363 GND 0.014412f
C2813 VDD.n1364 GND 0.008756f
C2814 VDD.n1366 GND 0.008756f
C2815 VDD.n1367 GND 0.008756f
C2816 VDD.n1368 GND 0.007048f
C2817 VDD.n1369 GND 0.007048f
C2818 VDD.n1370 GND 0.007048f
C2819 VDD.n1371 GND 0.008756f
C2820 VDD.n1373 GND 0.008756f
C2821 VDD.n1374 GND 0.008756f
C2822 VDD.n1375 GND 0.007048f
C2823 VDD.n1376 GND 0.007048f
C2824 VDD.n1377 GND 0.007048f
C2825 VDD.n1378 GND 0.008756f
C2826 VDD.n1380 GND 0.008756f
C2827 VDD.n1381 GND 0.008756f
C2828 VDD.n1382 GND 0.007048f
C2829 VDD.n1384 GND 0.444061f
C2830 VDD.n1386 GND 0.007048f
C2831 VDD.n1387 GND 0.007048f
C2832 VDD.n1388 GND 0.007048f
C2833 VDD.n1389 GND 0.008756f
C2834 VDD.n1391 GND 0.008756f
C2835 VDD.n1392 GND 0.008756f
C2836 VDD.n1393 GND 0.007048f
C2837 VDD.n1394 GND 0.00585f
C2838 VDD.n1395 GND 0.01973f
C2839 VDD.n1396 GND 0.019672f
C2840 VDD.n1397 GND 0.00585f
C2841 VDD.n1398 GND 0.019672f
C2842 VDD.n1399 GND 0.902878f
C2843 VDD.n1400 GND 0.019672f
C2844 VDD.n1401 GND 0.01973f
C2845 VDD.n1402 GND 0.003348f
C2846 VDD.n1403 GND 0.01973f
C2847 VDD.n1404 GND 0.008756f
C2848 VDD.n1405 GND 0.008756f
C2849 VDD.n1406 GND 0.007048f
C2850 VDD.n1407 GND 0.007048f
C2851 VDD.n1408 GND 0.007048f
C2852 VDD.n1409 GND 0.00753f
C2853 VDD.n1410 GND 0.444061f
C2854 VDD.n1411 GND 0.011781f
C2855 VDD.n1412 GND 0.004466f
C2856 VDD.n1413 GND 0.005954f
C2857 VDD.n1414 GND 0.005954f
C2858 VDD.n1415 GND 0.005954f
C2859 VDD.n1416 GND 0.005954f
C2860 VDD.n1417 GND 0.005954f
C2861 VDD.n1419 GND 0.005954f
C2862 VDD.n1420 GND 0.005954f
C2863 VDD.n1421 GND 0.005954f
C2864 VDD.n1422 GND 0.005954f
C2865 VDD.n1423 GND 0.005954f
C2866 VDD.n1425 GND 0.005954f
C2867 VDD.n1427 GND 0.005954f
C2868 VDD.n1428 GND 0.005954f
C2869 VDD.n1429 GND 0.005954f
C2870 VDD.n1430 GND 0.005954f
C2871 VDD.n1431 GND 0.005954f
C2872 VDD.n1433 GND 0.005954f
C2873 VDD.n1435 GND 0.005954f
C2874 VDD.n1436 GND 0.005954f
C2875 VDD.n1437 GND 0.005954f
C2876 VDD.n1438 GND 0.005954f
C2877 VDD.n1439 GND 0.005954f
C2878 VDD.n1441 GND 0.005954f
C2879 VDD.n1443 GND 0.005954f
C2880 VDD.n1444 GND 0.004466f
C2881 VDD.n1445 GND 0.005954f
C2882 VDD.n1446 GND 0.005954f
C2883 VDD.n1447 GND 0.005954f
C2884 VDD.n1449 GND 0.005954f
C2885 VDD.n1451 GND 0.005954f
C2886 VDD.n1452 GND 0.005954f
C2887 VDD.n1453 GND 0.005954f
C2888 VDD.n1454 GND 0.005954f
C2889 VDD.n1455 GND 0.005954f
C2890 VDD.n1457 GND 0.005954f
C2891 VDD.n1459 GND 0.005954f
C2892 VDD.n1460 GND 0.005954f
C2893 VDD.n1461 GND 0.004597f
C2894 VDD.n1462 GND 0.008509f
C2895 VDD.n1463 GND 0.004334f
C2896 VDD.n1464 GND 0.005954f
C2897 VDD.n1466 GND 0.005954f
C2898 VDD.n1467 GND 0.01392f
C2899 VDD.n1468 GND 0.01392f
C2900 VDD.n1469 GND 0.013224f
C2901 VDD.n1470 GND 0.005954f
C2902 VDD.n1471 GND 0.005954f
C2903 VDD.n1472 GND 0.005954f
C2904 VDD.n1473 GND 0.005954f
C2905 VDD.n1474 GND 0.005954f
C2906 VDD.n1475 GND 0.005954f
C2907 VDD.n1476 GND 0.005954f
C2908 VDD.n1477 GND 0.005954f
C2909 VDD.n1478 GND 0.005954f
C2910 VDD.n1479 GND 0.005954f
C2911 VDD.n1480 GND 0.005954f
C2912 VDD.n1481 GND 0.005954f
C2913 VDD.n1482 GND 0.005954f
C2914 VDD.n1483 GND 0.005954f
C2915 VDD.n1484 GND 0.005954f
C2916 VDD.n1485 GND 0.005954f
C2917 VDD.n1486 GND 0.005954f
C2918 VDD.n1487 GND 0.005954f
C2919 VDD.n1488 GND 0.005954f
C2920 VDD.n1489 GND 0.005954f
C2921 VDD.n1490 GND 0.005954f
C2922 VDD.n1491 GND 0.005954f
C2923 VDD.n1492 GND 0.005954f
C2924 VDD.n1493 GND 0.005954f
C2925 VDD.n1494 GND 0.005954f
C2926 VDD.n1495 GND 0.005954f
C2927 VDD.n1496 GND 0.005954f
C2928 VDD.n1497 GND 0.005954f
C2929 VDD.n1498 GND 0.005954f
C2930 VDD.n1499 GND 0.005954f
C2931 VDD.n1500 GND 0.005954f
C2932 VDD.n1501 GND 0.005954f
C2933 VDD.n1502 GND 0.005954f
C2934 VDD.n1503 GND 0.005954f
C2935 VDD.n1504 GND 0.005954f
C2936 VDD.n1505 GND 0.005954f
C2937 VDD.n1506 GND 0.005954f
C2938 VDD.n1507 GND 0.005954f
C2939 VDD.n1508 GND 0.005954f
C2940 VDD.n1509 GND 0.005954f
C2941 VDD.n1510 GND 0.005954f
C2942 VDD.n1511 GND 0.005954f
C2943 VDD.n1512 GND 0.005954f
C2944 VDD.n1513 GND 0.005954f
C2945 VDD.n1514 GND 0.005954f
C2946 VDD.n1515 GND 0.005954f
C2947 VDD.n1516 GND 0.005954f
C2948 VDD.n1517 GND 0.005954f
C2949 VDD.n1518 GND 0.005954f
C2950 VDD.n1519 GND 0.005954f
C2951 VDD.n1520 GND 0.005954f
C2952 VDD.n1521 GND 0.005954f
C2953 VDD.n1522 GND 0.005954f
C2954 VDD.n1523 GND 0.005954f
C2955 VDD.n1524 GND 0.005954f
C2956 VDD.n1525 GND 0.005954f
C2957 VDD.n1526 GND 0.005954f
C2958 VDD.n1527 GND 0.005954f
C2959 VDD.n1528 GND 0.005954f
C2960 VDD.n1529 GND 0.005954f
C2961 VDD.n1530 GND 0.005954f
C2962 VDD.n1531 GND 0.005954f
C2963 VDD.n1532 GND 0.005954f
C2964 VDD.n1533 GND 0.005954f
C2965 VDD.n1534 GND 0.005954f
C2966 VDD.n1535 GND 0.005954f
C2967 VDD.n1536 GND 0.005954f
C2968 VDD.n1537 GND 0.005954f
C2969 VDD.n1538 GND 0.005954f
C2970 VDD.n1539 GND 0.005954f
C2971 VDD.n1540 GND 0.319696f
C2972 VDD.n1541 GND 0.005954f
C2973 VDD.n1542 GND 0.005954f
C2974 VDD.n1543 GND 0.005954f
C2975 VDD.n1544 GND 0.005954f
C2976 VDD.n1545 GND 0.005954f
C2977 VDD.n1546 GND 0.005954f
C2978 VDD.n1547 GND 0.005954f
C2979 VDD.n1548 GND 0.005954f
C2980 VDD.n1549 GND 0.319696f
C2981 VDD.n1550 GND 0.005954f
C2982 VDD.n1551 GND 0.005954f
C2983 VDD.n1552 GND 0.005954f
C2984 VDD.n1553 GND 0.005954f
C2985 VDD.n1554 GND 0.005954f
C2986 VDD.n1555 GND 0.005954f
C2987 VDD.n1556 GND 0.005954f
C2988 VDD.n1557 GND 0.005954f
C2989 VDD.n1558 GND 0.005954f
C2990 VDD.n1559 GND 0.005954f
C2991 VDD.n1560 GND 0.005954f
C2992 VDD.n1561 GND 0.005954f
C2993 VDD.n1562 GND 0.005954f
C2994 VDD.n1563 GND 0.005954f
C2995 VDD.n1564 GND 0.005954f
C2996 VDD.n1565 GND 0.005954f
C2997 VDD.n1566 GND 0.005954f
C2998 VDD.n1567 GND 0.005954f
C2999 VDD.n1568 GND 0.005954f
C3000 VDD.n1569 GND 0.005954f
C3001 VDD.n1570 GND 0.005954f
C3002 VDD.n1571 GND 0.005954f
C3003 VDD.n1572 GND 0.005954f
C3004 VDD.n1573 GND 0.005954f
C3005 VDD.n1574 GND 0.005954f
C3006 VDD.n1575 GND 0.005954f
C3007 VDD.n1576 GND 0.005954f
C3008 VDD.n1577 GND 0.005954f
C3009 VDD.n1578 GND 0.005954f
C3010 VDD.n1579 GND 0.005954f
C3011 VDD.n1580 GND 0.005954f
C3012 VDD.n1581 GND 0.005954f
C3013 VDD.n1582 GND 0.013224f
C3014 VDD.n1583 GND 0.01392f
C3015 VDD.n1584 GND 0.01392f
C3016 VDD.n1585 GND 0.005954f
C3017 VDD.n1586 GND 0.005954f
C3018 VDD.n1587 GND 0.004334f
C3019 VDD.n1588 GND 0.005954f
C3020 VDD.n1590 GND 0.005954f
C3021 VDD.n1591 GND 0.004597f
C3022 VDD.n1592 GND 0.005954f
C3023 VDD.n1593 GND 0.005954f
C3024 VDD.n1594 GND 0.005954f
C3025 VDD.n1596 GND 0.005954f
C3026 VDD.n1598 GND 0.005954f
C3027 VDD.n1599 GND 0.005954f
C3028 VDD.n1600 GND 0.005954f
C3029 VDD.n1601 GND 0.005954f
C3030 VDD.n1602 GND 0.005954f
C3031 VDD.n1604 GND 0.005954f
C3032 VDD.n1605 GND 0.005954f
C3033 VDD.n1606 GND 0.005954f
C3034 VDD.n1607 GND 0.004466f
C3035 VDD.n1608 GND 0.005954f
C3036 VDD.n1610 GND 0.005954f
C3037 VDD.n1611 GND 0.004466f
C3038 VDD.n1612 GND 0.005954f
C3039 VDD.n1613 GND 0.005954f
C3040 VDD.n1614 GND 0.005954f
C3041 VDD.n1616 GND 0.005954f
C3042 VDD.n1618 GND 0.005954f
C3043 VDD.n1619 GND 0.005954f
C3044 VDD.n1620 GND 0.005954f
C3045 VDD.n1621 GND 0.005954f
C3046 VDD.n1622 GND 0.005954f
C3047 VDD.n1624 GND 0.005954f
C3048 VDD.n1625 GND 0.005954f
C3049 VDD.n1626 GND 0.005954f
C3050 VDD.n1627 GND 0.005954f
C3051 VDD.n1628 GND 0.005954f
C3052 VDD.n1629 GND 0.005954f
C3053 VDD.n1631 GND 0.005954f
C3054 VDD.n1632 GND 0.005954f
C3055 VDD.n1633 GND 0.01392f
C3056 VDD.n1634 GND 0.013224f
C3057 VDD.n1635 GND 0.013224f
C3058 VDD.n1636 GND 0.660471f
C3059 VDD.n1637 GND 0.013224f
C3060 VDD.n1638 GND 0.013224f
C3061 VDD.n1639 GND 0.005954f
C3062 VDD.n1640 GND 0.005954f
C3063 VDD.n1641 GND 0.005954f
C3064 VDD.n1642 GND 0.477788f
C3065 VDD.n1643 GND 0.005954f
C3066 VDD.n1644 GND 0.005954f
C3067 VDD.n1645 GND 0.005954f
C3068 VDD.n1646 GND 0.005954f
C3069 VDD.n1647 GND 0.005954f
C3070 VDD.n1648 GND 0.453196f
C3071 VDD.n1649 GND 0.005954f
C3072 VDD.n1650 GND 0.005954f
C3073 VDD.n1651 GND 0.004991f
C3074 VDD.n1652 GND 0.017249f
C3075 VDD.n1653 GND 0.00394f
C3076 VDD.n1654 GND 0.005954f
C3077 VDD.n1655 GND 0.316183f
C3078 VDD.n1656 GND 0.005954f
C3079 VDD.n1657 GND 0.005954f
C3080 VDD.n1658 GND 0.005954f
C3081 VDD.n1659 GND 0.005954f
C3082 VDD.n1660 GND 0.005954f
C3083 VDD.n1661 GND 0.477788f
C3084 VDD.n1662 GND 0.005954f
C3085 VDD.n1663 GND 0.005954f
C3086 VDD.n1664 GND 0.005954f
C3087 VDD.n1665 GND 0.005954f
C3088 VDD.n1666 GND 0.005954f
C3089 VDD.n1667 GND 0.291591f
C3090 VDD.n1668 GND 0.005954f
C3091 VDD.n1669 GND 0.005954f
C3092 VDD.n1670 GND 0.005954f
C3093 VDD.n1671 GND 0.005954f
C3094 VDD.n1672 GND 0.005954f
C3095 VDD.n1673 GND 0.428604f
C3096 VDD.n1674 GND 0.005954f
C3097 VDD.n1675 GND 0.005954f
C3098 VDD.n1676 GND 0.005954f
C3099 VDD.n1677 GND 0.005954f
C3100 VDD.n1678 GND 0.005954f
C3101 VDD.n1679 GND 0.270512f
C3102 VDD.n1680 GND 0.005954f
C3103 VDD.n1681 GND 0.005954f
C3104 VDD.n1682 GND 0.005954f
C3105 VDD.n1683 GND 0.005954f
C3106 VDD.n1684 GND 0.005954f
C3107 VDD.n1685 GND 0.407525f
C3108 VDD.n1686 GND 0.005954f
C3109 VDD.n1687 GND 0.005954f
C3110 VDD.n1688 GND 0.005954f
C3111 VDD.n1689 GND 0.005954f
C3112 VDD.n1690 GND 0.005954f
C3113 VDD.n1691 GND 0.249433f
C3114 VDD.n1692 GND 0.005954f
C3115 VDD.n1693 GND 0.005954f
C3116 VDD.n1694 GND 0.005954f
C3117 VDD.n1695 GND 0.005954f
C3118 VDD.n1696 GND 0.005954f
C3119 VDD.n1697 GND 0.386446f
C3120 VDD.n1698 GND 0.005954f
C3121 VDD.n1699 GND 0.005954f
C3122 VDD.n1700 GND 0.005954f
C3123 VDD.n1701 GND 0.005954f
C3124 VDD.n1702 GND 0.005954f
C3125 VDD.n1703 GND 0.249433f
C3126 VDD.n1704 GND 0.005954f
C3127 VDD.n1705 GND 0.005954f
C3128 VDD.n1706 GND 0.005954f
C3129 VDD.n1707 GND 0.005954f
C3130 VDD.n1708 GND 0.005954f
C3131 VDD.n1709 GND 0.365367f
C3132 VDD.n1710 GND 0.005954f
C3133 VDD.n1711 GND 0.005954f
C3134 VDD.n1712 GND 0.005954f
C3135 VDD.n1713 GND 0.005954f
C3136 VDD.n1714 GND 0.005954f
C3137 VDD.n1715 GND 0.270512f
C3138 VDD.n1716 GND 0.005954f
C3139 VDD.n1717 GND 0.005954f
C3140 VDD.n1718 GND 0.005954f
C3141 VDD.n1719 GND 0.005954f
C3142 VDD.n1720 GND 0.005954f
C3143 VDD.n1721 GND 0.477788f
C3144 VDD.n1722 GND 0.005954f
C3145 VDD.n1723 GND 0.005954f
C3146 VDD.n1724 GND 0.005954f
C3147 VDD.n1725 GND 0.005954f
C3148 VDD.n1726 GND 0.005954f
C3149 VDD.n1727 GND 0.186197f
C3150 VDD.n1728 GND 0.005954f
C3151 VDD.n1729 GND 0.005954f
C3152 VDD.n1730 GND 0.005954f
C3153 VDD.n1731 GND 0.005954f
C3154 VDD.n1732 GND 0.005954f
C3155 VDD.n1733 GND 0.477788f
C3156 VDD.n1734 GND 0.005954f
C3157 VDD.n1735 GND 0.005954f
C3158 VDD.n1736 GND 0.005954f
C3159 VDD.n1737 GND 0.005954f
C3160 VDD.n1738 GND 0.005954f
C3161 VDD.n1739 GND 0.351315f
C3162 VDD.n1740 GND 0.005954f
C3163 VDD.n1741 GND 0.005954f
C3164 VDD.n1742 GND 0.005954f
C3165 VDD.n1743 GND 0.005954f
C3166 VDD.n1744 GND 0.005954f
C3167 VDD.n1745 GND 0.005954f
C3168 VDD.n1746 GND 0.453196f
C3169 VDD.n1747 GND 0.005954f
C3170 VDD.n1748 GND 0.005954f
C3171 VDD.n1749 GND 0.005954f
C3172 VDD.n1750 GND 0.005954f
C3173 VDD.n1751 GND 0.005954f
C3174 VDD.n1752 GND 0.005954f
C3175 VDD.n1753 GND 0.330236f
C3176 VDD.n1754 GND 0.005954f
C3177 VDD.n1755 GND 0.005954f
C3178 VDD.n1756 GND 0.005954f
C3179 VDD.n1757 GND 0.013956f
C3180 VDD.n1758 GND 0.013224f
C3181 VDD.n1759 GND 0.01392f
C3182 VDD.n1760 GND 0.013188f
C3183 VDD.n1761 GND 0.005954f
C3184 VDD.n1762 GND 0.005954f
C3185 VDD.n1763 GND 0.005954f
C3186 VDD.n1764 GND 0.004334f
C3187 VDD.n1765 GND 0.008509f
C3188 VDD.n1766 GND 0.004597f
C3189 VDD.n1767 GND 0.005954f
C3190 VDD.n1768 GND 0.005954f
C3191 VDD.n1769 GND 0.005954f
C3192 VDD.n1770 GND 0.005954f
C3193 VDD.n1771 GND 0.005954f
C3194 VDD.n1772 GND 0.005954f
C3195 VDD.n1773 GND 0.005954f
C3196 VDD.n1774 GND 0.005954f
C3197 VDD.n1775 GND 0.005954f
C3198 VDD.n1776 GND 0.005954f
C3199 VDD.n1777 GND 0.005954f
C3200 VDD.n1778 GND 0.005954f
C3201 VDD.n1779 GND 0.005954f
C3202 VDD.n1780 GND 0.005954f
C3203 VDD.n1781 GND 0.005954f
C3204 VDD.n1782 GND 0.005954f
C3205 VDD.n1783 GND 0.005954f
C3206 VDD.n1784 GND 0.005954f
C3207 VDD.n1785 GND 0.005954f
C3208 VDD.n1786 GND 0.005954f
C3209 VDD.n1787 GND 0.005954f
C3210 VDD.n1788 GND 0.005954f
C3211 VDD.n1789 GND 0.005954f
C3212 VDD.n1790 GND 0.005954f
C3213 VDD.n1791 GND 0.005954f
C3214 VDD.n1792 GND 0.005954f
C3215 VDD.n1793 GND 0.005954f
C3216 VDD.n1794 GND 0.005954f
C3217 VDD.n1795 GND 0.005954f
C3218 VDD.n1796 GND 0.005954f
C3219 VDD.n1797 GND 0.005954f
C3220 VDD.n1798 GND 0.005954f
C3221 VDD.n1799 GND 0.005954f
C3222 VDD.n1800 GND 0.005954f
C3223 VDD.n1801 GND 0.005954f
C3224 VDD.n1802 GND 0.005954f
C3225 VDD.n1803 GND 0.005954f
C3226 VDD.n1804 GND 0.005954f
C3227 VDD.n1805 GND 0.005954f
C3228 VDD.n1806 GND 0.005954f
C3229 VDD.n1807 GND 0.005954f
C3230 VDD.n1808 GND 0.005954f
C3231 VDD.n1809 GND 0.005954f
C3232 VDD.n1810 GND 0.01392f
C3233 VDD.n1811 GND 0.01392f
C3234 VDD.n1812 GND 0.013224f
C3235 VDD.n1813 GND 0.005954f
C3236 VDD.n1814 GND 0.005954f
C3237 VDD.n1815 GND 0.386446f
C3238 VDD.n1816 GND 0.005954f
C3239 VDD.n1817 GND 0.013224f
C3240 VDD.n1818 GND 0.013956f
C3241 VDD.n1819 GND 0.013188f
C3242 VDD.n1820 GND 0.005954f
C3243 VDD.n1821 GND 0.005954f
C3244 VDD.n1822 GND 0.004334f
C3245 VDD.n1823 GND 0.005954f
C3246 VDD.n1824 GND 0.005954f
C3247 VDD.n1825 GND 0.004597f
C3248 VDD.n1826 GND 0.005954f
C3249 VDD.n1827 GND 0.005954f
C3250 VDD.n1828 GND 0.005954f
C3251 VDD.n1829 GND 0.005954f
C3252 VDD.n1830 GND 0.005954f
C3253 VDD.n1831 GND 0.005954f
C3254 VDD.n1832 GND 0.005954f
C3255 VDD.n1833 GND 0.005954f
C3256 VDD.n1834 GND 0.005954f
C3257 VDD.n1835 GND 0.005954f
C3258 VDD.n1836 GND 0.005954f
C3259 VDD.n1837 GND 0.005954f
C3260 VDD.n1838 GND 0.005954f
C3261 VDD.n1839 GND 0.005954f
C3262 VDD.n1840 GND 0.005954f
C3263 VDD.n1841 GND 0.005954f
C3264 VDD.n1842 GND 0.005954f
C3265 VDD.n1843 GND 0.005954f
C3266 VDD.n1844 GND 0.005954f
C3267 VDD.n1845 GND 0.005954f
C3268 VDD.n1846 GND 0.005954f
C3269 VDD.n1847 GND 0.005954f
C3270 VDD.n1848 GND 0.005954f
C3271 VDD.n1849 GND 0.005954f
C3272 VDD.n1850 GND 0.005954f
C3273 VDD.n1851 GND 0.005954f
C3274 VDD.n1852 GND 0.005954f
C3275 VDD.n1853 GND 0.005954f
C3276 VDD.n1854 GND 0.005954f
C3277 VDD.n1855 GND 0.005954f
C3278 VDD.n1856 GND 0.005954f
C3279 VDD.n1857 GND 0.005954f
C3280 VDD.n1858 GND 0.005954f
C3281 VDD.n1859 GND 0.005954f
C3282 VDD.n1860 GND 0.005954f
C3283 VDD.n1861 GND 0.005954f
C3284 VDD.n1862 GND 0.005954f
C3285 VDD.n1863 GND 0.005954f
C3286 VDD.n1864 GND 0.005954f
C3287 VDD.n1865 GND 0.005954f
C3288 VDD.n1866 GND 0.005954f
C3289 VDD.n1867 GND 0.01392f
C3290 VDD.n1868 GND 0.01392f
C3291 VDD.n1869 GND 0.548051f
C3292 VDD.t16 GND 2.42407f
C3293 VDD.t5 GND 2.42407f
C3294 VDD.n1870 GND 0.548051f
C3295 VDD.n1871 GND 0.013224f
C3296 VDD.n1872 GND 0.013224f
C3297 VDD.n1873 GND 0.386446f
C3298 VDD.n1874 GND 0.01392f
C3299 VDD.n1875 GND 0.005954f
C3300 VDD.n1876 GND 0.005954f
C3301 VDD.n1877 GND 0.005954f
C3302 VDD.n1878 GND 0.005954f
C3303 VDD.n1879 GND 0.005954f
C3304 VDD.n1880 GND 0.005954f
C3305 VDD.n1881 GND 0.005954f
C3306 VDD.n1882 GND 0.005954f
C3307 VDD.n1883 GND 0.005954f
C3308 VDD.n1884 GND 0.005954f
C3309 VDD.n1885 GND 0.004597f
C3310 VDD.n1886 GND 0.005954f
C3311 VDD.t60 GND 0.076127f
C3312 VDD.t61 GND 0.086562f
C3313 VDD.t58 GND 0.227136f
C3314 VDD.n1887 GND 0.151662f
C3315 VDD.n1888 GND 0.122136f
C3316 VDD.n1889 GND 0.008509f
C3317 VDD.n1890 GND 0.005954f
C3318 VDD.n1891 GND 0.005954f
C3319 VDD.n1892 GND 0.005954f
C3320 VDD.t81 GND 0.076127f
C3321 VDD.t82 GND 0.086562f
C3322 VDD.t80 GND 0.227136f
C3323 VDD.n1893 GND 0.151662f
C3324 VDD.n1894 GND 0.122136f
C3325 VDD.n1895 GND 0.005954f
C3326 VDD.n1896 GND 0.005954f
C3327 VDD.n1897 GND 0.005954f
C3328 VDD.n1898 GND 0.005954f
C3329 VDD.n1899 GND 0.005954f
C3330 VDD.n1900 GND 0.005954f
C3331 VDD.n1901 GND 0.005954f
C3332 VDD.n1902 GND 0.005954f
C3333 VDD.n1903 GND 0.005954f
C3334 VDD.n1904 GND 0.005954f
C3335 VDD.n1906 GND 0.005954f
C3336 VDD.n1907 GND 0.005954f
C3337 VDD.n1908 GND 0.005954f
C3338 VDD.n1909 GND 0.005954f
C3339 VDD.n1910 GND 0.005954f
C3340 VDD.n1912 GND 0.005954f
C3341 VDD.n1914 GND 0.005954f
C3342 VDD.n1915 GND 0.005954f
C3343 VDD.n1916 GND 0.005954f
C3344 VDD.n1917 GND 0.005954f
C3345 VDD.n1918 GND 0.005954f
C3346 VDD.n1920 GND 0.005954f
C3347 VDD.n1922 GND 0.005954f
C3348 VDD.n1923 GND 0.005954f
C3349 VDD.n1924 GND 0.005954f
C3350 VDD.n1925 GND 0.005954f
C3351 VDD.n1926 GND 0.005954f
C3352 VDD.n1928 GND 0.005954f
C3353 VDD.n1930 GND 0.005954f
C3354 VDD.n1931 GND 0.005954f
C3355 VDD.n1932 GND 0.005954f
C3356 VDD.n1933 GND 0.005954f
C3357 VDD.n1934 GND 0.005954f
C3358 VDD.n1936 GND 0.005954f
C3359 VDD.n1938 GND 0.005954f
C3360 VDD.n1939 GND 0.005954f
C3361 VDD.n1940 GND 0.005954f
C3362 VDD.n1941 GND 0.005954f
C3363 VDD.n1942 GND 0.005954f
C3364 VDD.n1944 GND 0.005954f
C3365 VDD.n1946 GND 0.005954f
C3366 VDD.n1947 GND 0.005954f
C3367 VDD.n1948 GND 0.004597f
C3368 VDD.n1949 GND 0.008509f
C3369 VDD.n1950 GND 0.004334f
C3370 VDD.n1951 GND 0.005954f
C3371 VDD.n1953 GND 0.005954f
C3372 VDD.n1954 GND 0.01392f
C3373 VDD.n1955 GND 0.01392f
C3374 VDD.n1956 GND 0.013224f
C3375 VDD.n1957 GND 0.005954f
C3376 VDD.n1958 GND 0.005954f
C3377 VDD.n1959 GND 0.005954f
C3378 VDD.n1960 GND 0.005954f
C3379 VDD.n1961 GND 0.005954f
C3380 VDD.n1962 GND 0.005954f
C3381 VDD.n1963 GND 0.005954f
C3382 VDD.n1964 GND 0.005954f
C3383 VDD.n1965 GND 0.005954f
C3384 VDD.n1966 GND 0.005954f
C3385 VDD.n1967 GND 0.005954f
C3386 VDD.n1968 GND 0.005954f
C3387 VDD.n1969 GND 0.005954f
C3388 VDD.n1970 GND 0.005954f
C3389 VDD.n1971 GND 0.005954f
C3390 VDD.n1972 GND 0.005954f
C3391 VDD.n1973 GND 0.005954f
C3392 VDD.n1974 GND 0.005954f
C3393 VDD.n1975 GND 0.005954f
C3394 VDD.n1976 GND 0.005954f
C3395 VDD.n1977 GND 0.005954f
C3396 VDD.n1978 GND 0.005954f
C3397 VDD.n1979 GND 0.005954f
C3398 VDD.n1980 GND 0.005954f
C3399 VDD.n1981 GND 0.005954f
C3400 VDD.n1982 GND 0.005954f
C3401 VDD.n1983 GND 0.005954f
C3402 VDD.n1984 GND 0.005954f
C3403 VDD.n1985 GND 0.005954f
C3404 VDD.n1986 GND 0.005954f
C3405 VDD.n1987 GND 0.005954f
C3406 VDD.n1988 GND 0.005954f
C3407 VDD.n1989 GND 0.005954f
C3408 VDD.n1990 GND 0.005954f
C3409 VDD.n1991 GND 0.005954f
C3410 VDD.n1992 GND 0.005954f
C3411 VDD.n1993 GND 0.005954f
C3412 VDD.n1994 GND 0.005954f
C3413 VDD.n1995 GND 0.005954f
C3414 VDD.n1996 GND 0.005954f
C3415 VDD.n1997 GND 0.005954f
C3416 VDD.n1998 GND 0.005954f
C3417 VDD.n1999 GND 0.005954f
C3418 VDD.n2000 GND 0.005954f
C3419 VDD.n2001 GND 0.005954f
C3420 VDD.n2002 GND 0.005954f
C3421 VDD.n2003 GND 0.005954f
C3422 VDD.n2004 GND 0.005954f
C3423 VDD.n2005 GND 0.005954f
C3424 VDD.n2006 GND 0.005954f
C3425 VDD.n2007 GND 0.005954f
C3426 VDD.n2008 GND 0.005954f
C3427 VDD.n2009 GND 0.005954f
C3428 VDD.n2010 GND 0.005954f
C3429 VDD.n2011 GND 0.005954f
C3430 VDD.n2012 GND 0.005954f
C3431 VDD.n2013 GND 0.005954f
C3432 VDD.n2014 GND 0.005954f
C3433 VDD.n2015 GND 0.005954f
C3434 VDD.n2016 GND 0.005954f
C3435 VDD.n2017 GND 0.005954f
C3436 VDD.n2018 GND 0.005954f
C3437 VDD.n2019 GND 0.005954f
C3438 VDD.n2020 GND 0.005954f
C3439 VDD.n2021 GND 0.005954f
C3440 VDD.n2022 GND 0.005954f
C3441 VDD.n2023 GND 0.005954f
C3442 VDD.n2024 GND 0.005954f
C3443 VDD.n2025 GND 0.005954f
C3444 VDD.n2026 GND 0.005954f
C3445 VDD.n2027 GND 0.005954f
C3446 VDD.n2028 GND 0.005954f
C3447 VDD.n2029 GND 0.005954f
C3448 VDD.n2030 GND 0.005954f
C3449 VDD.n2031 GND 0.005954f
C3450 VDD.n2032 GND 0.005954f
C3451 VDD.n2033 GND 0.005954f
C3452 VDD.n2034 GND 0.005954f
C3453 VDD.n2035 GND 0.005954f
C3454 VDD.n2036 GND 0.005954f
C3455 VDD.n2037 GND 0.005954f
C3456 VDD.n2038 GND 0.319696f
C3457 VDD.n2039 GND 0.005954f
C3458 VDD.n2040 GND 0.005954f
C3459 VDD.n2041 GND 0.005954f
C3460 VDD.n2042 GND 0.005954f
C3461 VDD.n2043 GND 0.005954f
C3462 VDD.n2044 GND 0.005954f
C3463 VDD.n2045 GND 0.005954f
C3464 VDD.n2046 GND 0.005954f
C3465 VDD.n2047 GND 0.319696f
C3466 VDD.n2048 GND 0.005954f
C3467 VDD.n2049 GND 0.005954f
C3468 VDD.n2050 GND 0.005954f
C3469 VDD.n2051 GND 0.005954f
C3470 VDD.n2052 GND 0.005954f
C3471 VDD.n2053 GND 0.005954f
C3472 VDD.n2054 GND 0.005954f
C3473 VDD.n2055 GND 0.005954f
C3474 VDD.n2056 GND 0.005954f
C3475 VDD.n2057 GND 0.005954f
C3476 VDD.n2058 GND 0.005954f
C3477 VDD.n2059 GND 0.005954f
C3478 VDD.n2060 GND 0.005954f
C3479 VDD.n2061 GND 0.005954f
C3480 VDD.n2062 GND 0.005954f
C3481 VDD.n2063 GND 0.005954f
C3482 VDD.n2064 GND 0.005954f
C3483 VDD.n2065 GND 0.005954f
C3484 VDD.n2066 GND 0.005954f
C3485 VDD.n2067 GND 0.005954f
C3486 VDD.n2068 GND 0.005954f
C3487 VDD.n2069 GND 0.005954f
C3488 VDD.n2070 GND 0.005954f
C3489 VDD.n2071 GND 0.013224f
C3490 VDD.n2073 GND 0.01392f
C3491 VDD.n2074 GND 0.01392f
C3492 VDD.n2075 GND 0.005954f
C3493 VDD.n2076 GND 0.004334f
C3494 VDD.n2077 GND 0.005954f
C3495 VDD.n2079 GND 0.005954f
C3496 VDD.n2081 GND 0.005954f
C3497 VDD.n2082 GND 0.005954f
C3498 VDD.n2083 GND 0.005954f
C3499 VDD.n2084 GND 0.005954f
C3500 VDD.n2085 GND 0.005954f
C3501 VDD.n2087 GND 0.005954f
C3502 VDD.n2089 GND 0.005954f
C3503 VDD.n2090 GND 0.005954f
C3504 VDD.n2091 GND 0.005954f
C3505 VDD.n2092 GND 0.005954f
C3506 VDD.n2093 GND 0.005954f
C3507 VDD.n2095 GND 0.005954f
C3508 VDD.n2097 GND 0.005954f
C3509 VDD.n2098 GND 0.005954f
C3510 VDD.n2099 GND 0.005954f
C3511 VDD.n2100 GND 0.005954f
C3512 VDD.n2101 GND 0.005954f
C3513 VDD.n2103 GND 0.005954f
C3514 VDD.n2105 GND 0.005954f
C3515 VDD.n2106 GND 0.005954f
C3516 VDD.n2107 GND 0.005954f
C3517 VDD.n2108 GND 0.005954f
C3518 VDD.n2109 GND 0.005954f
C3519 VDD.n2111 GND 0.005954f
C3520 VDD.n2113 GND 0.005954f
C3521 VDD.n2114 GND 0.005954f
C3522 VDD.n2115 GND 0.005954f
C3523 VDD.n2116 GND 0.005954f
C3524 VDD.n2117 GND 0.005954f
C3525 VDD.n2119 GND 0.005954f
C3526 VDD.n2121 GND 0.005954f
C3527 VDD.n2122 GND 0.005954f
C3528 VDD.n2123 GND 0.01392f
C3529 VDD.n2124 GND 0.013224f
C3530 VDD.n2125 GND 0.013224f
C3531 VDD.n2126 GND 0.660471f
C3532 VDD.n2127 GND 0.013224f
C3533 VDD.n2128 GND 0.013224f
C3534 VDD.n2129 GND 0.005954f
C3535 VDD.n2130 GND 0.005954f
C3536 VDD.n2131 GND 0.005954f
C3537 VDD.n2132 GND 0.330236f
C3538 VDD.n2133 GND 0.005954f
C3539 VDD.n2134 GND 0.005954f
C3540 VDD.n2135 GND 0.005954f
C3541 VDD.n2136 GND 0.005954f
C3542 VDD.n2137 GND 0.005954f
C3543 VDD.n2138 GND 0.453196f
C3544 VDD.n2139 GND 0.005954f
C3545 VDD.n2140 GND 0.005954f
C3546 VDD.n2141 GND 0.005954f
C3547 VDD.n2142 GND 0.005954f
C3548 VDD.n2143 GND 0.005954f
C3549 VDD.n2144 GND 0.351315f
C3550 VDD.n2145 GND 0.005954f
C3551 VDD.n2146 GND 0.005954f
C3552 VDD.n2147 GND 0.005954f
C3553 VDD.n2148 GND 0.005954f
C3554 VDD.n2149 GND 0.005954f
C3555 VDD.n2150 GND 0.477788f
C3556 VDD.n2151 GND 0.005954f
C3557 VDD.n2152 GND 0.005954f
C3558 VDD.n2153 GND 0.005954f
C3559 VDD.n2154 GND 0.005954f
C3560 VDD.n2155 GND 0.005954f
C3561 VDD.n2156 GND 0.186197f
C3562 VDD.n2157 GND 0.005954f
C3563 VDD.n2158 GND 0.005954f
C3564 VDD.n2159 GND 0.005954f
C3565 VDD.n2160 GND 0.005954f
C3566 VDD.n2161 GND 0.005954f
C3567 VDD.n2162 GND 0.477788f
C3568 VDD.n2163 GND 0.005954f
C3569 VDD.n2164 GND 0.005954f
C3570 VDD.n2165 GND 0.005954f
C3571 VDD.n2166 GND 0.005954f
C3572 VDD.n2167 GND 0.005954f
C3573 VDD.n2168 GND 0.270512f
C3574 VDD.n2169 GND 0.005954f
C3575 VDD.n2170 GND 0.005954f
C3576 VDD.n2171 GND 0.005954f
C3577 VDD.n2172 GND 0.005954f
C3578 VDD.n2173 GND 0.005954f
C3579 VDD.n2174 GND 0.365367f
C3580 VDD.n2175 GND 0.005954f
C3581 VDD.n2176 GND 0.005954f
C3582 VDD.n2177 GND 0.005954f
C3583 VDD.n2178 GND 0.005954f
C3584 VDD.n2179 GND 0.005954f
C3585 VDD.n2180 GND 0.249433f
C3586 VDD.n2181 GND 0.005954f
C3587 VDD.n2182 GND 0.005954f
C3588 VDD.n2183 GND 0.005954f
C3589 VDD.n2184 GND 0.005954f
C3590 VDD.n2185 GND 0.005954f
C3591 VDD.n2186 GND 0.386446f
C3592 VDD.n2187 GND 0.005954f
C3593 VDD.n2188 GND 0.005954f
C3594 VDD.n2189 GND 0.005954f
C3595 VDD.n2190 GND 0.005954f
C3596 VDD.n2191 GND 0.005954f
C3597 VDD.n2192 GND 0.249433f
C3598 VDD.n2193 GND 0.005954f
C3599 VDD.n2194 GND 0.005954f
C3600 VDD.n2195 GND 0.005954f
C3601 VDD.n2196 GND 0.005954f
C3602 VDD.n2197 GND 0.005954f
C3603 VDD.n2198 GND 0.407525f
C3604 VDD.n2199 GND 0.005954f
C3605 VDD.n2200 GND 0.005954f
C3606 VDD.n2201 GND 0.005954f
C3607 VDD.n2202 GND 0.005954f
C3608 VDD.n2203 GND 0.005954f
C3609 VDD.n2204 GND 0.270512f
C3610 VDD.n2205 GND 0.005954f
C3611 VDD.n2206 GND 0.005954f
C3612 VDD.n2207 GND 0.005954f
C3613 VDD.n2208 GND 0.005954f
C3614 VDD.n2209 GND 0.005954f
C3615 VDD.n2210 GND 0.428604f
C3616 VDD.n2211 GND 0.005954f
C3617 VDD.n2212 GND 0.005954f
C3618 VDD.n2213 GND 0.005954f
C3619 VDD.n2214 GND 0.005954f
C3620 VDD.n2215 GND 0.005954f
C3621 VDD.n2216 GND 0.291591f
C3622 VDD.n2217 GND 0.005954f
C3623 VDD.n2218 GND 0.005954f
C3624 VDD.n2219 GND 0.005954f
C3625 VDD.n2220 GND 0.005954f
C3626 VDD.n2221 GND 0.005954f
C3627 VDD.n2222 GND 0.477788f
C3628 VDD.n2223 GND 0.005954f
C3629 VDD.n2224 GND 0.005954f
C3630 VDD.n2225 GND 0.005954f
C3631 VDD.n2226 GND 0.005954f
C3632 VDD.n2227 GND 0.005954f
C3633 VDD.n2228 GND 0.316183f
C3634 VDD.n2229 GND 0.005954f
C3635 VDD.n2230 GND 0.00394f
C3636 VDD.n2231 GND 0.017249f
C3637 VDD.n2232 GND 0.004991f
C3638 VDD.n2233 GND 0.005954f
C3639 VDD.n2234 GND 0.005954f
C3640 VDD.n2235 GND 0.005954f
C3641 VDD.n2236 GND 0.005954f
C3642 VDD.n2238 GND 0.005954f
C3643 VDD.n2239 GND 0.005954f
C3644 VDD.n2241 GND 0.005954f
C3645 VDD.n2242 GND 0.005954f
C3646 VDD.n2243 GND 0.005954f
C3647 VDD.n2245 GND 0.005954f
C3648 VDD.n2246 GND 0.005954f
C3649 VDD.n2247 GND 0.005954f
C3650 VDD.n2248 GND 0.005954f
C3651 VDD.n2249 GND 0.005954f
C3652 VDD.n2250 GND 0.005954f
C3653 VDD.n2252 GND 0.005954f
C3654 VDD.n2253 GND 0.005954f
C3655 VDD.n2254 GND 0.005954f
C3656 VDD.n2255 GND 0.005954f
C3657 VDD.n2256 GND 0.005954f
C3658 VDD.n2257 GND 0.005954f
C3659 VDD.n2259 GND 0.005954f
C3660 VDD.n2260 GND 0.005954f
C3661 VDD.n2262 GND 0.01392f
C3662 VDD.n2263 GND 0.01392f
C3663 VDD.n2264 GND 0.013224f
C3664 VDD.n2265 GND 0.005954f
C3665 VDD.n2266 GND 0.005954f
C3666 VDD.n2267 GND 0.005954f
C3667 VDD.n2268 GND 0.005954f
C3668 VDD.n2269 GND 0.005954f
C3669 VDD.n2270 GND 0.005954f
C3670 VDD.n2271 GND 0.453196f
C3671 VDD.n2272 GND 0.005954f
C3672 VDD.n2273 GND 0.005954f
C3673 VDD.n2274 GND 0.005954f
C3674 VDD.n2275 GND 0.005954f
C3675 VDD.n2276 GND 0.005954f
C3676 VDD.n2277 GND 0.477788f
C3677 VDD.n2278 GND 0.005954f
C3678 VDD.n2279 GND 0.005954f
C3679 VDD.n2280 GND 0.005954f
C3680 VDD.n2281 GND 0.013956f
C3681 VDD.n2282 GND 0.013188f
C3682 VDD.n2283 GND 0.01392f
C3683 VDD.n2285 GND 0.005954f
C3684 VDD.n2286 GND 0.005954f
C3685 VDD.n2287 GND 0.004334f
C3686 VDD.n2288 GND 0.008509f
C3687 VDD.n2289 GND 0.004597f
C3688 VDD.n2290 GND 0.005954f
C3689 VDD.n2291 GND 0.005954f
C3690 VDD.n2293 GND 0.005954f
C3691 VDD.n2294 GND 0.005954f
C3692 VDD.n2295 GND 0.005954f
C3693 VDD.n2296 GND 0.005954f
C3694 VDD.n2297 GND 0.005954f
C3695 VDD.n2298 GND 0.005954f
C3696 VDD.n2300 GND 0.005954f
C3697 VDD.n2301 GND 0.005954f
C3698 VDD.n2302 GND 0.005954f
C3699 VDD.n2303 GND 0.005954f
C3700 VDD.n2304 GND 0.004466f
C3701 VDD.n2305 GND 0.005954f
C3702 VDD.n2307 GND 0.005954f
C3703 VDD.n2308 GND 0.004466f
C3704 VDD.n2309 GND 0.005954f
C3705 VDD.n2310 GND 0.005954f
C3706 VDD.n2312 GND 0.005954f
C3707 VDD.n2313 GND 0.005954f
C3708 VDD.n2314 GND 0.005954f
C3709 VDD.n2315 GND 0.005954f
C3710 VDD.n2316 GND 0.005954f
C3711 VDD.n2317 GND 0.005954f
C3712 VDD.n2319 GND 0.005954f
C3713 VDD.n2320 GND 0.005954f
C3714 VDD.n2321 GND 0.005954f
C3715 VDD.n2322 GND 0.005954f
C3716 VDD.n2323 GND 0.005954f
C3717 VDD.n2324 GND 0.005954f
C3718 VDD.n2326 GND 0.005954f
C3719 VDD.n2327 GND 0.005954f
C3720 VDD.n2328 GND 0.005954f
C3721 VDD.n2329 GND 0.01392f
C3722 VDD.n2330 GND 0.013224f
C3723 VDD.n2331 GND 0.013224f
C3724 VDD.n2332 GND 0.660471f
C3725 VDD.n2333 GND 0.013224f
C3726 VDD.n2334 GND 0.01392f
C3727 VDD.n2335 GND 0.013188f
C3728 VDD.n2336 GND 0.005954f
C3729 VDD.n2337 GND 0.004334f
C3730 VDD.n2338 GND 0.005954f
C3731 VDD.n2340 GND 0.005954f
C3732 VDD.n2341 GND 0.005954f
C3733 VDD.n2342 GND 0.005954f
C3734 VDD.n2343 GND 0.005954f
C3735 VDD.n2344 GND 0.005954f
C3736 VDD.n2345 GND 0.005954f
C3737 VDD.n2347 GND 0.005954f
C3738 VDD.n2348 GND 0.005954f
C3739 VDD.n2349 GND 0.005954f
C3740 VDD.n2350 GND 0.005954f
C3741 VDD.n2351 GND 0.005954f
C3742 VDD.n2352 GND 0.005954f
C3743 VDD.n2354 GND 0.005954f
C3744 VDD.n2355 GND 0.005954f
C3745 VDD.n2356 GND 0.004466f
C3746 VDD.n2357 GND 0.008306f
C3747 VDD.n2358 GND 0.008756f
C3748 VDD.n2359 GND 0.008756f
C3749 VDD.n2360 GND 0.007048f
C3750 VDD.n2361 GND 0.008756f
C3751 VDD.n2362 GND 0.008756f
C3752 VDD.n2363 GND 0.008756f
C3753 VDD.n2364 GND 0.008756f
C3754 VDD.n2365 GND 0.01973f
C3755 VDD.n2366 GND 0.003348f
C3756 VDD.t72 GND 0.17936f
C3757 VDD.t73 GND 0.187962f
C3758 VDD.t70 GND 0.262044f
C3759 VDD.n2367 GND 0.088819f
C3760 VDD.n2368 GND 0.050925f
C3761 VDD.n2369 GND 0.010889f
C3762 VDD.n2370 GND 0.008756f
C3763 VDD.n2371 GND 0.0037f
C3764 VDD.n2372 GND 0.007048f
C3765 VDD.n2373 GND 0.008756f
C3766 VDD.n2374 GND 0.008756f
C3767 VDD.n2375 GND 0.007048f
C3768 VDD.n2376 GND 0.008756f
C3769 VDD.n2377 GND 0.007048f
C3770 VDD.n2378 GND 0.007048f
C3771 VDD.n2380 GND 0.447535f
C3772 VDD.n2382 GND 0.007048f
C3773 VDD.n2383 GND 0.008756f
C3774 VDD.n2384 GND 0.008756f
C3775 VDD.n2385 GND 0.007048f
C3776 VDD.n2386 GND 0.007048f
C3777 VDD.n2387 GND 0.008756f
C3778 VDD.n2388 GND 0.008756f
C3779 VDD.n2389 GND 0.007048f
C3780 VDD.n2390 GND 0.007048f
C3781 VDD.n2391 GND 0.008756f
C3782 VDD.n2392 GND 0.008756f
C3783 VDD.n2393 GND 0.007048f
C3784 VDD.n2394 GND 0.007048f
C3785 VDD.n2395 GND 0.008756f
C3786 VDD.n2396 GND 0.008756f
C3787 VDD.n2397 GND 0.007048f
C3788 VDD.n2398 GND 0.007048f
C3789 VDD.n2399 GND 0.008756f
C3790 VDD.n2400 GND 0.008756f
C3791 VDD.n2401 GND 0.007048f
C3792 VDD.n2402 GND 0.008756f
C3793 VDD.n2403 GND 0.008756f
C3794 VDD.n2404 GND 0.007048f
C3795 VDD.n2405 GND 0.008756f
C3796 VDD.n2406 GND 0.008756f
C3797 VDD.n2407 GND 0.008756f
C3798 VDD.n2408 GND 0.014412f
C3799 VDD.n2409 GND 0.008756f
C3800 VDD.n2410 GND 0.008756f
C3801 VDD.n2411 GND 0.004792f
C3802 VDD.n2412 GND 0.007048f
C3803 VDD.n2413 GND 0.008756f
C3804 VDD.n2414 GND 0.008756f
C3805 VDD.n2415 GND 0.007048f
C3806 VDD.n2416 GND 0.007048f
C3807 VDD.n2417 GND 0.008756f
C3808 VDD.n2418 GND 0.008756f
C3809 VDD.n2419 GND 0.007048f
C3810 VDD.n2420 GND 0.007048f
C3811 VDD.n2421 GND 0.008756f
C3812 VDD.n2422 GND 0.008756f
C3813 VDD.n2423 GND 0.007048f
C3814 VDD.n2424 GND 0.007048f
C3815 VDD.n2425 GND 0.008756f
C3816 VDD.n2426 GND 0.008756f
C3817 VDD.n2427 GND 0.007048f
C3818 VDD.n2428 GND 0.007048f
C3819 VDD.n2429 GND 0.008756f
C3820 VDD.n2430 GND 0.008756f
C3821 VDD.n2431 GND 0.007048f
C3822 VDD.n2432 GND 0.007048f
C3823 VDD.n2433 GND 0.008756f
C3824 VDD.n2434 GND 0.008756f
C3825 VDD.n2435 GND 0.007048f
C3826 VDD.n2436 GND 0.007048f
C3827 VDD.n2437 GND 0.008756f
C3828 VDD.n2438 GND 0.008756f
C3829 VDD.n2439 GND 0.007048f
C3830 VDD.n2440 GND 0.007048f
C3831 VDD.n2441 GND 0.008756f
C3832 VDD.n2442 GND 0.008756f
C3833 VDD.n2443 GND 0.007048f
C3834 VDD.n2444 GND 0.008756f
C3835 VDD.n2445 GND 0.008756f
C3836 VDD.n2446 GND 0.007048f
C3837 VDD.n2447 GND 0.008756f
C3838 VDD.n2448 GND 0.008756f
C3839 VDD.n2449 GND 0.008756f
C3840 VDD.t84 GND 0.17936f
C3841 VDD.t85 GND 0.187962f
C3842 VDD.t83 GND 0.262044f
C3843 VDD.n2450 GND 0.088819f
C3844 VDD.n2451 GND 0.050925f
C3845 VDD.n2452 GND 0.014412f
C3846 VDD.n2453 GND 0.008756f
C3847 VDD.n2454 GND 0.008756f
C3848 VDD.n2455 GND 0.005885f
C3849 VDD.n2456 GND 0.007048f
C3850 VDD.n2457 GND 0.008756f
C3851 VDD.n2458 GND 0.008756f
C3852 VDD.n2459 GND 0.007048f
C3853 VDD.n2460 GND 0.007048f
C3854 VDD.n2461 GND 0.008756f
C3855 VDD.n2462 GND 0.008756f
C3856 VDD.n2463 GND 0.007048f
C3857 VDD.n2464 GND 0.007048f
C3858 VDD.n2465 GND 0.008756f
C3859 VDD.n2466 GND 0.008756f
C3860 VDD.n2467 GND 0.007048f
C3861 VDD.n2468 GND 0.008756f
C3862 VDD.n2469 GND 0.007048f
C3863 VDD.n2470 GND 0.007048f
C3864 VDD.n2472 GND 0.447535f
C3865 VDD.n2474 GND 0.007048f
C3866 VDD.n2475 GND 0.008756f
C3867 VDD.n2476 GND 0.008756f
C3868 VDD.n2477 GND 0.007048f
C3869 VDD.n2478 GND 0.007048f
C3870 VDD.n2479 GND 0.007048f
C3871 VDD.n2480 GND 0.008756f
C3872 VDD.n2481 GND 4.24037f
C3873 VDD.n2483 GND 0.01973f
C3874 VDD.n2484 GND 0.00585f
C3875 VDD.n2485 GND 0.01973f
C3876 VDD.n2486 GND 0.019672f
C3877 VDD.n2487 GND 0.008756f
C3878 VDD.n2488 GND 0.007048f
C3879 VDD.n2489 GND 0.008756f
C3880 VDD.n2490 GND 0.593722f
C3881 VDD.n2491 GND 0.008756f
C3882 VDD.n2492 GND 0.007048f
C3883 VDD.n2493 GND 0.008756f
C3884 VDD.n2494 GND 0.008756f
C3885 VDD.n2495 GND 0.008756f
C3886 VDD.n2496 GND 0.007048f
C3887 VDD.n2497 GND 0.008756f
C3888 VDD.n2498 GND 0.702629f
C3889 VDD.n2499 GND 0.008756f
C3890 VDD.n2500 GND 0.007048f
C3891 VDD.n2501 GND 0.008756f
C3892 VDD.n2502 GND 0.008756f
C3893 VDD.n2503 GND 0.008756f
C3894 VDD.n2504 GND 0.007048f
C3895 VDD.n2505 GND 0.008756f
C3896 VDD.n2506 GND 0.702629f
C3897 VDD.n2507 GND 0.008756f
C3898 VDD.n2508 GND 0.007048f
C3899 VDD.n2509 GND 0.008756f
C3900 VDD.n2510 GND 0.008756f
C3901 VDD.n2511 GND 0.008756f
C3902 VDD.n2512 GND 0.007048f
C3903 VDD.n2513 GND 0.008756f
C3904 VDD.n2514 GND 0.516432f
C3905 VDD.n2515 GND 0.008756f
C3906 VDD.n2516 GND 0.007048f
C3907 VDD.n2517 GND 0.008756f
C3908 VDD.n2518 GND 0.008756f
C3909 VDD.n2519 GND 0.008756f
C3910 VDD.n2520 GND 0.007048f
C3911 VDD.n2521 GND 0.008756f
C3912 VDD.n2522 GND 0.418064f
C3913 VDD.n2523 GND 0.008756f
C3914 VDD.n2524 GND 0.007048f
C3915 VDD.n2525 GND 0.008756f
C3916 VDD.n2526 GND 0.008756f
C3917 VDD.n2527 GND 0.008756f
C3918 VDD.n2528 GND 0.007048f
C3919 VDD.n2529 GND 0.008756f
C3920 VDD.t143 GND 0.351315f
C3921 VDD.n2530 GND 0.649932f
C3922 VDD.n2531 GND 0.008756f
C3923 VDD.n2532 GND 0.007048f
C3924 VDD.n2533 GND 0.008756f
C3925 VDD.n2534 GND 0.008756f
C3926 VDD.n2535 GND 0.008756f
C3927 VDD.n2536 GND 0.007048f
C3928 VDD.n2537 GND 0.008756f
C3929 VDD.n2538 GND 0.702629f
C3930 VDD.n2539 GND 0.008756f
C3931 VDD.n2540 GND 0.007048f
C3932 VDD.n2541 GND 0.008756f
C3933 VDD.n2542 GND 0.008756f
C3934 VDD.n2543 GND 0.008756f
C3935 VDD.n2544 GND 0.007048f
C3936 VDD.n2545 GND 0.008756f
C3937 VDD.n2546 GND 0.523459f
C3938 VDD.n2547 GND 0.008756f
C3939 VDD.n2548 GND 0.007048f
C3940 VDD.n2549 GND 0.008756f
C3941 VDD.n2550 GND 0.008756f
C3942 VDD.n2551 GND 0.008756f
C3943 VDD.n2552 GND 0.007048f
C3944 VDD.n2553 GND 0.008756f
C3945 VDD.n2554 GND 0.411038f
C3946 VDD.n2555 GND 0.008756f
C3947 VDD.n2556 GND 0.007048f
C3948 VDD.n2557 GND 0.008756f
C3949 VDD.n2558 GND 0.008756f
C3950 VDD.n2559 GND 0.008756f
C3951 VDD.n2560 GND 0.007048f
C3952 VDD.n2561 GND 0.007048f
C3953 VDD.n2562 GND 0.007048f
C3954 VDD.n2563 GND 0.008756f
C3955 VDD.n2564 GND 0.008756f
C3956 VDD.n2565 GND 0.008756f
C3957 VDD.n2566 GND 0.007048f
C3958 VDD.n2567 GND 0.007048f
C3959 VDD.n2568 GND 0.007048f
C3960 VDD.n2569 GND 0.008756f
C3961 VDD.n2570 GND 0.008756f
C3962 VDD.n2571 GND 0.008756f
C3963 VDD.n2572 GND 0.007048f
C3964 VDD.n2573 GND 0.007048f
C3965 VDD.n2574 GND 0.007048f
C3966 VDD.n2575 GND 0.008756f
C3967 VDD.n2576 GND 0.008756f
C3968 VDD.n2577 GND 0.008756f
C3969 VDD.n2578 GND 0.007048f
C3970 VDD.n2579 GND 0.007048f
C3971 VDD.n2580 GND 0.007048f
C3972 VDD.n2581 GND 0.008756f
C3973 VDD.n2582 GND 0.008756f
C3974 VDD.n2583 GND 0.008756f
C3975 VDD.n2584 GND 0.007048f
C3976 VDD.n2585 GND 0.007048f
C3977 VDD.n2586 GND 0.00585f
C3978 VDD.n2587 GND 0.019672f
C3979 VDD.n2588 GND 0.01973f
C3980 VDD.n2589 GND 0.003348f
C3981 VDD.n2590 GND 0.01973f
C3982 VDD.n2592 GND 0.008756f
C3983 VDD.n2593 GND 0.008756f
C3984 VDD.n2594 GND 0.007048f
C3985 VDD.n2595 GND 0.007048f
C3986 VDD.n2596 GND 0.007048f
C3987 VDD.n2597 GND 0.008756f
C3988 VDD.n2599 GND 0.008756f
C3989 VDD.n2600 GND 0.008756f
C3990 VDD.n2601 GND 0.007048f
C3991 VDD.n2602 GND 0.007048f
C3992 VDD.n2603 GND 0.007048f
C3993 VDD.n2604 GND 0.008756f
C3994 VDD.n2606 GND 0.008756f
C3995 VDD.n2607 GND 0.008756f
C3996 VDD.n2608 GND 0.007048f
C3997 VDD.n2609 GND 0.007048f
C3998 VDD.n2610 GND 0.007048f
C3999 VDD.n2611 GND 0.008756f
C4000 VDD.n2613 GND 0.008756f
C4001 VDD.n2614 GND 0.008756f
C4002 VDD.n2615 GND 0.007048f
C4003 VDD.n2616 GND 0.007048f
C4004 VDD.n2617 GND 0.007048f
C4005 VDD.n2618 GND 0.008756f
C4006 VDD.n2620 GND 0.008756f
C4007 VDD.n2621 GND 0.008756f
C4008 VDD.n2622 GND 0.007048f
C4009 VDD.n2623 GND 0.008756f
C4010 VDD.n2624 GND 0.008756f
C4011 VDD.n2625 GND 0.008756f
C4012 VDD.n2626 GND 0.014412f
C4013 VDD.n2627 GND 0.008756f
C4014 VDD.n2629 GND 0.008756f
C4015 VDD.n2630 GND 0.008756f
C4016 VDD.n2631 GND 0.007048f
C4017 VDD.n2632 GND 0.007048f
C4018 VDD.n2633 GND 0.007048f
C4019 VDD.n2634 GND 0.008756f
C4020 VDD.n2636 GND 0.008756f
C4021 VDD.n2637 GND 0.008756f
C4022 VDD.n2638 GND 0.007048f
C4023 VDD.n2639 GND 0.007048f
C4024 VDD.n2640 GND 0.007048f
C4025 VDD.n2641 GND 0.008756f
C4026 VDD.n2643 GND 0.008756f
C4027 VDD.n2644 GND 0.008756f
C4028 VDD.n2645 GND 0.007048f
C4029 VDD.n2646 GND 0.007048f
C4030 VDD.n2647 GND 0.007048f
C4031 VDD.n2648 GND 0.008756f
C4032 VDD.n2650 GND 0.008756f
C4033 VDD.n2651 GND 0.008756f
C4034 VDD.n2652 GND 0.007048f
C4035 VDD.n2653 GND 0.007048f
C4036 VDD.n2654 GND 0.007048f
C4037 VDD.n2655 GND 0.008756f
C4038 VDD.n2657 GND 0.008756f
C4039 VDD.n2658 GND 0.008756f
C4040 VDD.n2659 GND 0.007048f
C4041 VDD.n2660 GND 0.008756f
C4042 VDD.n2661 GND 0.008756f
C4043 VDD.n2662 GND 0.008756f
C4044 VDD.n2663 GND 0.014412f
C4045 VDD.n2664 GND 0.008756f
C4046 VDD.n2666 GND 0.008756f
C4047 VDD.n2667 GND 0.008756f
C4048 VDD.n2668 GND 0.007048f
C4049 VDD.n2669 GND 0.007048f
C4050 VDD.n2670 GND 0.007048f
C4051 VDD.n2671 GND 0.008756f
C4052 VDD.n2673 GND 0.008756f
C4053 VDD.n2674 GND 0.008756f
C4054 VDD.n2675 GND 0.007048f
C4055 VDD.n2676 GND 0.007048f
C4056 VDD.n2677 GND 0.007048f
C4057 VDD.n2678 GND 0.008756f
C4058 VDD.n2680 GND 0.008756f
C4059 VDD.n2681 GND 0.008756f
C4060 VDD.n2682 GND 0.007048f
C4061 VDD.n2683 GND 0.007048f
C4062 VDD.n2684 GND 0.007048f
C4063 VDD.n2685 GND 0.008756f
C4064 VDD.n2687 GND 0.008756f
C4065 VDD.n2688 GND 0.008756f
C4066 VDD.n2690 GND 0.008756f
C4067 VDD.n2691 GND 0.007048f
C4068 VDD.n2692 GND 0.007048f
C4069 VDD.n2693 GND 0.00585f
C4070 VDD.n2694 GND 0.01973f
C4071 VDD.n2695 GND 0.019672f
C4072 VDD.n2696 GND 0.00585f
C4073 VDD.n2697 GND 0.019672f
C4074 VDD.n2698 GND 0.902878f
C4075 VDD.n2699 GND 0.593722f
C4076 VDD.t63 GND 0.351315f
C4077 VDD.n2700 GND 0.460222f
C4078 VDD.n2701 GND 0.008756f
C4079 VDD.n2702 GND 0.007048f
C4080 VDD.n2703 GND 0.007048f
C4081 VDD.n2704 GND 0.007048f
C4082 VDD.n2705 GND 0.008756f
C4083 VDD.n2706 GND 0.702629f
C4084 VDD.n2707 GND 0.702629f
C4085 VDD.n2708 GND 0.537511f
C4086 VDD.n2709 GND 0.008756f
C4087 VDD.n2710 GND 0.007048f
C4088 VDD.n2711 GND 0.007048f
C4089 VDD.n2712 GND 0.007048f
C4090 VDD.n2713 GND 0.008756f
C4091 VDD.n2714 GND 0.702629f
C4092 VDD.n2715 GND 0.418064f
C4093 VDD.t160 GND 0.351315f
C4094 VDD.n2716 GND 0.635879f
C4095 VDD.n2717 GND 0.008756f
C4096 VDD.n2718 GND 0.007048f
C4097 VDD.n2719 GND 0.007048f
C4098 VDD.n2720 GND 0.007048f
C4099 VDD.n2721 GND 0.008756f
C4100 VDD.n2722 GND 0.404012f
C4101 VDD.n2723 GND 0.702629f
C4102 VDD.n2724 GND 0.530485f
C4103 VDD.n2725 GND 0.008756f
C4104 VDD.n2726 GND 0.007048f
C4105 VDD.n2727 GND 0.007048f
C4106 VDD.n2728 GND 0.007048f
C4107 VDD.n2729 GND 0.008756f
C4108 VDD.n2730 GND 0.702629f
C4109 VDD.n2731 GND 0.411038f
C4110 VDD.t130 GND 0.351315f
C4111 VDD.n2732 GND 0.642906f
C4112 VDD.n2733 GND 0.008756f
C4113 VDD.n2734 GND 0.007048f
C4114 VDD.n2735 GND 0.00673f
C4115 VDD.n2736 GND 0.238982f
C4116 VDD.n2737 GND 1.80661f
C4117 VOUT.t50 GND 0.039597f
C4118 VOUT.t70 GND 0.039597f
C4119 VOUT.n0 GND 0.295329f
C4120 VOUT.t29 GND 0.039597f
C4121 VOUT.t53 GND 0.039597f
C4122 VOUT.n1 GND 0.294088f
C4123 VOUT.n2 GND 0.437569f
C4124 VOUT.t40 GND 0.039597f
C4125 VOUT.t55 GND 0.039597f
C4126 VOUT.n3 GND 0.294088f
C4127 VOUT.n4 GND 0.216522f
C4128 VOUT.t80 GND 0.039597f
C4129 VOUT.t59 GND 0.039597f
C4130 VOUT.n5 GND 0.294088f
C4131 VOUT.n6 GND 0.216522f
C4132 VOUT.t54 GND 0.039597f
C4133 VOUT.t72 GND 0.039597f
C4134 VOUT.n7 GND 0.294088f
C4135 VOUT.n8 GND 0.361808f
C4136 VOUT.t74 GND 0.039597f
C4137 VOUT.t48 GND 0.039597f
C4138 VOUT.n9 GND 0.295329f
C4139 VOUT.t76 GND 0.039597f
C4140 VOUT.t51 GND 0.039597f
C4141 VOUT.n10 GND 0.294088f
C4142 VOUT.n11 GND 0.437569f
C4143 VOUT.t66 GND 0.039597f
C4144 VOUT.t41 GND 0.039597f
C4145 VOUT.n12 GND 0.294088f
C4146 VOUT.n13 GND 0.216522f
C4147 VOUT.t33 GND 0.039597f
C4148 VOUT.t75 GND 0.039597f
C4149 VOUT.n14 GND 0.294088f
C4150 VOUT.n15 GND 0.216522f
C4151 VOUT.t37 GND 0.039597f
C4152 VOUT.t78 GND 0.039597f
C4153 VOUT.n16 GND 0.294088f
C4154 VOUT.n17 GND 0.299809f
C4155 VOUT.n18 GND 0.556152f
C4156 VOUT.t63 GND 0.039597f
C4157 VOUT.t36 GND 0.039597f
C4158 VOUT.n19 GND 0.295329f
C4159 VOUT.t84 GND 0.039597f
C4160 VOUT.t79 GND 0.039597f
C4161 VOUT.n20 GND 0.294088f
C4162 VOUT.n21 GND 0.437569f
C4163 VOUT.t61 GND 0.039597f
C4164 VOUT.t42 GND 0.039597f
C4165 VOUT.n22 GND 0.294088f
C4166 VOUT.n23 GND 0.216522f
C4167 VOUT.t46 GND 0.039597f
C4168 VOUT.t83 GND 0.039597f
C4169 VOUT.n24 GND 0.294088f
C4170 VOUT.n25 GND 0.216522f
C4171 VOUT.t44 GND 0.039597f
C4172 VOUT.t71 GND 0.039597f
C4173 VOUT.n26 GND 0.294088f
C4174 VOUT.n27 GND 0.299809f
C4175 VOUT.n28 GND 0.540352f
C4176 VOUT.n29 GND 6.05558f
C4177 VOUT.n31 GND 0.641776f
C4178 VOUT.n32 GND 0.481332f
C4179 VOUT.n33 GND 0.641776f
C4180 VOUT.n34 GND 0.641776f
C4181 VOUT.n35 GND 1.72786f
C4182 VOUT.n36 GND 0.641776f
C4183 VOUT.n37 GND 0.641776f
C4184 VOUT.t95 GND 0.80222f
C4185 VOUT.n38 GND 0.641776f
C4186 VOUT.n39 GND 0.641776f
C4187 VOUT.n43 GND 0.641776f
C4188 VOUT.n47 GND 0.641776f
C4189 VOUT.n48 GND 0.641776f
C4190 VOUT.n50 GND 0.641776f
C4191 VOUT.n55 GND 0.641776f
C4192 VOUT.n57 GND 0.641776f
C4193 VOUT.n58 GND 0.641776f
C4194 VOUT.n60 GND 0.641776f
C4195 VOUT.n61 GND 0.641776f
C4196 VOUT.n63 GND 0.641776f
C4197 VOUT.t92 GND 10.724f
C4198 VOUT.n65 GND 0.641776f
C4199 VOUT.n66 GND 0.481332f
C4200 VOUT.n67 GND 0.641776f
C4201 VOUT.n68 GND 0.641776f
C4202 VOUT.n69 GND 1.72786f
C4203 VOUT.n70 GND 0.641776f
C4204 VOUT.n71 GND 0.641776f
C4205 VOUT.t97 GND 0.80222f
C4206 VOUT.n72 GND 0.641776f
C4207 VOUT.n73 GND 0.641776f
C4208 VOUT.n77 GND 0.641776f
C4209 VOUT.n81 GND 0.641776f
C4210 VOUT.n82 GND 0.641776f
C4211 VOUT.n84 GND 0.641776f
C4212 VOUT.n89 GND 0.641776f
C4213 VOUT.n91 GND 0.641776f
C4214 VOUT.n92 GND 0.641776f
C4215 VOUT.n94 GND 0.641776f
C4216 VOUT.n95 GND 0.641776f
C4217 VOUT.n97 GND 0.641776f
C4218 VOUT.n98 GND 0.481332f
C4219 VOUT.n100 GND 0.641776f
C4220 VOUT.n101 GND 0.481332f
C4221 VOUT.n102 GND 0.641776f
C4222 VOUT.n103 GND 0.641776f
C4223 VOUT.n104 GND 1.72786f
C4224 VOUT.n105 GND 0.641776f
C4225 VOUT.n106 GND 0.641776f
C4226 VOUT.t94 GND 0.80222f
C4227 VOUT.n107 GND 0.641776f
C4228 VOUT.n108 GND 1.72786f
C4229 VOUT.n110 GND 0.641776f
C4230 VOUT.n111 GND 0.641776f
C4231 VOUT.n113 GND 0.641776f
C4232 VOUT.n114 GND 0.641776f
C4233 VOUT.t93 GND 10.5492f
C4234 VOUT.t96 GND 10.724f
C4235 VOUT.n120 GND 2.01334f
C4236 VOUT.n121 GND 8.201639f
C4237 VOUT.n122 GND 8.54483f
C4238 VOUT.n127 GND 2.181f
C4239 VOUT.n133 GND 0.641776f
C4240 VOUT.n135 GND 0.641776f
C4241 VOUT.n137 GND 0.641776f
C4242 VOUT.n139 GND 0.641776f
C4243 VOUT.n141 GND 0.641776f
C4244 VOUT.n147 GND 0.641776f
C4245 VOUT.n154 GND 1.17741f
C4246 VOUT.n155 GND 1.17741f
C4247 VOUT.n156 GND 0.641776f
C4248 VOUT.n157 GND 0.641776f
C4249 VOUT.n159 GND 0.481332f
C4250 VOUT.n160 GND 0.412218f
C4251 VOUT.n162 GND 0.481332f
C4252 VOUT.n163 GND 0.412218f
C4253 VOUT.n164 GND 0.481332f
C4254 VOUT.n166 GND 0.641776f
C4255 VOUT.n168 GND 1.72786f
C4256 VOUT.n169 GND 2.01334f
C4257 VOUT.n170 GND 7.5434f
C4258 VOUT.n172 GND 0.481332f
C4259 VOUT.n173 GND 1.2385f
C4260 VOUT.n174 GND 0.481332f
C4261 VOUT.n176 GND 0.641776f
C4262 VOUT.n178 GND 1.72786f
C4263 VOUT.n179 GND 3.2304f
C4264 VOUT.n180 GND 2.16607f
C4265 VOUT.t64 GND 0.039597f
C4266 VOUT.t65 GND 0.039597f
C4267 VOUT.n181 GND 0.295329f
C4268 VOUT.t34 GND 0.039597f
C4269 VOUT.t67 GND 0.039597f
C4270 VOUT.n182 GND 0.294088f
C4271 VOUT.n183 GND 0.437569f
C4272 VOUT.t28 GND 0.039597f
C4273 VOUT.t57 GND 0.039597f
C4274 VOUT.n184 GND 0.294088f
C4275 VOUT.n185 GND 0.216522f
C4276 VOUT.t38 GND 0.039597f
C4277 VOUT.t45 GND 0.039597f
C4278 VOUT.n186 GND 0.294088f
C4279 VOUT.n187 GND 0.216522f
C4280 VOUT.t87 GND 0.039597f
C4281 VOUT.t35 GND 0.039597f
C4282 VOUT.n188 GND 0.294088f
C4283 VOUT.n189 GND 0.361808f
C4284 VOUT.t68 GND 0.039597f
C4285 VOUT.t31 GND 0.039597f
C4286 VOUT.n190 GND 0.295329f
C4287 VOUT.t60 GND 0.039597f
C4288 VOUT.t47 GND 0.039597f
C4289 VOUT.n191 GND 0.294088f
C4290 VOUT.n192 GND 0.437569f
C4291 VOUT.t49 GND 0.039597f
C4292 VOUT.t39 GND 0.039597f
C4293 VOUT.n193 GND 0.294088f
C4294 VOUT.n194 GND 0.216522f
C4295 VOUT.t43 GND 0.039597f
C4296 VOUT.t81 GND 0.039597f
C4297 VOUT.n195 GND 0.294088f
C4298 VOUT.n196 GND 0.216522f
C4299 VOUT.t85 GND 0.039597f
C4300 VOUT.t73 GND 0.039597f
C4301 VOUT.n197 GND 0.294088f
C4302 VOUT.n198 GND 0.299809f
C4303 VOUT.n199 GND 0.556152f
C4304 VOUT.t52 GND 0.039597f
C4305 VOUT.t82 GND 0.039597f
C4306 VOUT.n200 GND 0.295329f
C4307 VOUT.t86 GND 0.039597f
C4308 VOUT.t32 GND 0.039597f
C4309 VOUT.n201 GND 0.294088f
C4310 VOUT.n202 GND 0.437569f
C4311 VOUT.t56 GND 0.039597f
C4312 VOUT.t77 GND 0.039597f
C4313 VOUT.n203 GND 0.294088f
C4314 VOUT.n204 GND 0.216522f
C4315 VOUT.t69 GND 0.039597f
C4316 VOUT.t30 GND 0.039597f
C4317 VOUT.n205 GND 0.294088f
C4318 VOUT.n206 GND 0.216522f
C4319 VOUT.t58 GND 0.039597f
C4320 VOUT.t62 GND 0.039597f
C4321 VOUT.n207 GND 0.294086f
C4322 VOUT.n208 GND 0.29981f
C4323 VOUT.n209 GND 0.540352f
C4324 VOUT.n210 GND 8.69408f
C4325 VOUT.t20 GND 0.03394f
C4326 VOUT.t11 GND 0.03394f
C4327 VOUT.n211 GND 0.299314f
C4328 VOUT.t1 GND 0.03394f
C4329 VOUT.t21 GND 0.03394f
C4330 VOUT.n212 GND 0.296413f
C4331 VOUT.n213 GND 0.482682f
C4332 VOUT.t89 GND 0.03394f
C4333 VOUT.t5 GND 0.03394f
C4334 VOUT.n214 GND 0.296413f
C4335 VOUT.n215 GND 0.239908f
C4336 VOUT.t23 GND 0.03394f
C4337 VOUT.t14 GND 0.03394f
C4338 VOUT.n216 GND 0.296413f
C4339 VOUT.n217 GND 0.369148f
C4340 VOUT.t15 GND 0.03394f
C4341 VOUT.t18 GND 0.03394f
C4342 VOUT.n218 GND 0.299314f
C4343 VOUT.t6 GND 0.03394f
C4344 VOUT.t27 GND 0.03394f
C4345 VOUT.n219 GND 0.296413f
C4346 VOUT.n220 GND 0.482682f
C4347 VOUT.t22 GND 0.03394f
C4348 VOUT.t19 GND 0.03394f
C4349 VOUT.n221 GND 0.296413f
C4350 VOUT.n222 GND 0.239908f
C4351 VOUT.t0 GND 0.03394f
C4352 VOUT.t3 GND 0.03394f
C4353 VOUT.n223 GND 0.296413f
C4354 VOUT.n224 GND 0.317044f
C4355 VOUT.n225 GND 0.820783f
C4356 VOUT.n226 GND 8.86432f
C4357 VOUT.t2 GND 0.03394f
C4358 VOUT.t90 GND 0.03394f
C4359 VOUT.n227 GND 0.299314f
C4360 VOUT.t16 GND 0.03394f
C4361 VOUT.t91 GND 0.03394f
C4362 VOUT.n228 GND 0.296413f
C4363 VOUT.n229 GND 0.482682f
C4364 VOUT.t13 GND 0.03394f
C4365 VOUT.t17 GND 0.03394f
C4366 VOUT.n230 GND 0.296413f
C4367 VOUT.n231 GND 0.239908f
C4368 VOUT.t24 GND 0.03394f
C4369 VOUT.t88 GND 0.03394f
C4370 VOUT.n232 GND 0.296413f
C4371 VOUT.n233 GND 0.369148f
C4372 VOUT.t9 GND 0.03394f
C4373 VOUT.t8 GND 0.03394f
C4374 VOUT.n234 GND 0.299314f
C4375 VOUT.t7 GND 0.03394f
C4376 VOUT.t10 GND 0.03394f
C4377 VOUT.n235 GND 0.296413f
C4378 VOUT.n236 GND 0.482682f
C4379 VOUT.t4 GND 0.03394f
C4380 VOUT.t25 GND 0.03394f
C4381 VOUT.n237 GND 0.296413f
C4382 VOUT.n238 GND 0.239908f
C4383 VOUT.t12 GND 0.03394f
C4384 VOUT.t26 GND 0.03394f
C4385 VOUT.n239 GND 0.296413f
C4386 VOUT.n240 GND 0.317044f
C4387 VOUT.n241 GND 0.820783f
C4388 VOUT.n242 GND 5.33936f
C4389 VOUT.n243 GND 6.29717f
C4390 a_n7677_8299.n0 GND 0.656987f
C4391 a_n7677_8299.n1 GND 0.497097f
C4392 a_n7677_8299.n2 GND 0.656987f
C4393 a_n7677_8299.n3 GND 0.497097f
C4394 a_n7677_8299.n4 GND 0.876082f
C4395 a_n7677_8299.n5 GND 0.038978f
C4396 a_n7677_8299.n6 GND 0.038978f
C4397 a_n7677_8299.n7 GND 0.086056f
C4398 a_n7677_8299.n8 GND 0.050479f
C4399 a_n7677_8299.n9 GND 0.381855f
C4400 a_n7677_8299.n10 GND 0.381855f
C4401 a_n7677_8299.n11 GND 0.381855f
C4402 a_n7677_8299.n12 GND 0.041149f
C4403 a_n7677_8299.n13 GND 0.038977f
C4404 a_n7677_8299.n14 GND 0.041141f
C4405 a_n7677_8299.n15 GND 0.041141f
C4406 a_n7677_8299.n16 GND 0.041149f
C4407 a_n7677_8299.n17 GND 0.038977f
C4408 a_n7677_8299.n18 GND 0.041141f
C4409 a_n7677_8299.n19 GND 0.041141f
C4410 a_n7677_8299.n20 GND 0.041149f
C4411 a_n7677_8299.n21 GND 0.038977f
C4412 a_n7677_8299.n22 GND 0.041141f
C4413 a_n7677_8299.n23 GND 0.387272f
C4414 a_n7677_8299.n24 GND 0.043786f
C4415 a_n7677_8299.n25 GND 0.387272f
C4416 a_n7677_8299.n26 GND 0.043786f
C4417 a_n7677_8299.n27 GND 0.387272f
C4418 a_n7677_8299.n28 GND 0.043786f
C4419 a_n7677_8299.n29 GND 0.050479f
C4420 a_n7677_8299.n30 GND 0.050479f
C4421 a_n7677_8299.n31 GND 0.050479f
C4422 a_n7677_8299.n32 GND 0.043257f
C4423 a_n7677_8299.n33 GND 0.226705f
C4424 a_n7677_8299.n34 GND 0.086056f
C4425 a_n7677_8299.n35 GND 0.042023f
C4426 a_n7677_8299.n36 GND 0.226705f
C4427 a_n7677_8299.n37 GND 0.042023f
C4428 a_n7677_8299.n38 GND 0.086056f
C4429 a_n7677_8299.n39 GND 0.086056f
C4430 a_n7677_8299.n40 GND 0.043257f
C4431 a_n7677_8299.n41 GND 0.086056f
C4432 a_n7677_8299.n42 GND 0.050479f
C4433 a_n7677_8299.n43 GND 0.069364f
C4434 a_n7677_8299.n44 GND 0.042282f
C4435 a_n7677_8299.n45 GND 0.086056f
C4436 a_n7677_8299.n46 GND 0.086056f
C4437 a_n7677_8299.n47 GND 0.086056f
C4438 a_n7677_8299.n48 GND 0.086056f
C4439 a_n7677_8299.n49 GND 0.05002f
C4440 a_n7677_8299.n50 GND 0.069329f
C4441 a_n7677_8299.n51 GND 0.042569f
C4442 a_n7677_8299.n52 GND 0.086056f
C4443 a_n7677_8299.n53 GND 0.100444f
C4444 a_n7677_8299.n54 GND 0.226705f
C4445 a_n7677_8299.n55 GND 0.042023f
C4446 a_n7677_8299.n56 GND 0.086056f
C4447 a_n7677_8299.n57 GND 0.086056f
C4448 a_n7677_8299.n58 GND 0.043257f
C4449 a_n7677_8299.n59 GND 0.086056f
C4450 a_n7677_8299.n60 GND 0.050479f
C4451 a_n7677_8299.n61 GND 0.069364f
C4452 a_n7677_8299.n62 GND 0.042282f
C4453 a_n7677_8299.n63 GND 0.086056f
C4454 a_n7677_8299.n64 GND 0.086056f
C4455 a_n7677_8299.n65 GND 0.086056f
C4456 a_n7677_8299.n66 GND 0.086056f
C4457 a_n7677_8299.n67 GND 0.05002f
C4458 a_n7677_8299.n68 GND 0.069329f
C4459 a_n7677_8299.n69 GND 0.042569f
C4460 a_n7677_8299.n70 GND 0.086056f
C4461 a_n7677_8299.n71 GND 0.100444f
C4462 a_n7677_8299.n72 GND 0.226705f
C4463 a_n7677_8299.n73 GND 0.042023f
C4464 a_n7677_8299.n74 GND 0.086056f
C4465 a_n7677_8299.n75 GND 0.086056f
C4466 a_n7677_8299.n76 GND 0.043257f
C4467 a_n7677_8299.n77 GND 0.086056f
C4468 a_n7677_8299.n78 GND 0.050479f
C4469 a_n7677_8299.n79 GND 0.069364f
C4470 a_n7677_8299.n80 GND 0.042282f
C4471 a_n7677_8299.n81 GND 0.086056f
C4472 a_n7677_8299.n82 GND 0.086056f
C4473 a_n7677_8299.n83 GND 0.086056f
C4474 a_n7677_8299.n84 GND 0.086056f
C4475 a_n7677_8299.n85 GND 0.05002f
C4476 a_n7677_8299.n86 GND 0.069329f
C4477 a_n7677_8299.n87 GND 0.042569f
C4478 a_n7677_8299.n88 GND 0.086056f
C4479 a_n7677_8299.n89 GND 0.100444f
C4480 a_n7677_8299.t15 GND 0.092851f
C4481 a_n7677_8299.t4 GND 0.079586f
C4482 a_n7677_8299.t5 GND 0.079586f
C4483 a_n7677_8299.n90 GND 0.575059f
C4484 a_n7677_8299.t1 GND 0.079586f
C4485 a_n7677_8299.t18 GND 0.079586f
C4486 a_n7677_8299.n91 GND 0.572385f
C4487 a_n7677_8299.n92 GND 1.00831f
C4488 a_n7677_8299.t7 GND 0.079586f
C4489 a_n7677_8299.t9 GND 0.079586f
C4490 a_n7677_8299.n93 GND 0.572385f
C4491 a_n7677_8299.n94 GND 2.25795f
C4492 a_n7677_8299.t10 GND 0.079586f
C4493 a_n7677_8299.t17 GND 0.079586f
C4494 a_n7677_8299.n95 GND 0.575061f
C4495 a_n7677_8299.t11 GND 0.079586f
C4496 a_n7677_8299.t19 GND 0.079586f
C4497 a_n7677_8299.n96 GND 0.572385f
C4498 a_n7677_8299.n97 GND 1.00831f
C4499 a_n7677_8299.t16 GND 0.079586f
C4500 a_n7677_8299.t6 GND 0.079586f
C4501 a_n7677_8299.n98 GND 0.572385f
C4502 a_n7677_8299.n99 GND 1.55752f
C4503 a_n7677_8299.n100 GND 4.83804f
C4504 a_n7677_8299.t57 GND 0.803901f
C4505 a_n7677_8299.t36 GND 0.803901f
C4506 a_n7677_8299.t42 GND 0.803901f
C4507 a_n7677_8299.t23 GND 0.803901f
C4508 a_n7677_8299.t55 GND 0.803901f
C4509 a_n7677_8299.n101 GND 0.387598f
C4510 a_n7677_8299.t34 GND 0.803901f
C4511 a_n7677_8299.n102 GND 0.320757f
C4512 a_n7677_8299.t70 GND 0.803901f
C4513 a_n7677_8299.n103 GND 0.398918f
C4514 a_n7677_8299.t40 GND 0.895722f
C4515 a_n7677_8299.n104 GND 0.382689f
C4516 a_n7677_8299.n105 GND 0.069384f
C4517 a_n7677_8299.n106 GND 0.068166f
C4518 a_n7677_8299.n107 GND 0.396278f
C4519 a_n7677_8299.n108 GND 0.320757f
C4520 a_n7677_8299.n109 GND 0.067918f
C4521 a_n7677_8299.t54 GND 0.803901f
C4522 a_n7677_8299.n110 GND 0.396531f
C4523 a_n7677_8299.n111 GND 0.320757f
C4524 a_n7677_8299.n112 GND 0.058503f
C4525 a_n7677_8299.t62 GND 0.869419f
C4526 a_n7677_8299.n113 GND 0.387049f
C4527 a_n7677_8299.n114 GND 0.2593f
C4528 a_n7677_8299.t29 GND 0.803901f
C4529 a_n7677_8299.t67 GND 0.803901f
C4530 a_n7677_8299.t76 GND 0.803901f
C4531 a_n7677_8299.t49 GND 0.803901f
C4532 a_n7677_8299.t28 GND 0.803901f
C4533 a_n7677_8299.n115 GND 0.387598f
C4534 a_n7677_8299.t65 GND 0.803901f
C4535 a_n7677_8299.n116 GND 0.320757f
C4536 a_n7677_8299.t37 GND 0.803901f
C4537 a_n7677_8299.n117 GND 0.398918f
C4538 a_n7677_8299.t73 GND 0.895722f
C4539 a_n7677_8299.n118 GND 0.382689f
C4540 a_n7677_8299.n119 GND 0.069384f
C4541 a_n7677_8299.n120 GND 0.068166f
C4542 a_n7677_8299.n121 GND 0.396278f
C4543 a_n7677_8299.n122 GND 0.320757f
C4544 a_n7677_8299.n123 GND 0.067918f
C4545 a_n7677_8299.t27 GND 0.803901f
C4546 a_n7677_8299.n124 GND 0.396531f
C4547 a_n7677_8299.n125 GND 0.320757f
C4548 a_n7677_8299.n126 GND 0.058503f
C4549 a_n7677_8299.t32 GND 0.869419f
C4550 a_n7677_8299.n127 GND 0.387049f
C4551 a_n7677_8299.n128 GND 0.138484f
C4552 a_n7677_8299.n129 GND 0.702378f
C4553 a_n7677_8299.t68 GND 0.803901f
C4554 a_n7677_8299.t21 GND 0.803901f
C4555 a_n7677_8299.t61 GND 0.803901f
C4556 a_n7677_8299.t77 GND 0.803901f
C4557 a_n7677_8299.t25 GND 0.803901f
C4558 a_n7677_8299.n130 GND 0.387598f
C4559 a_n7677_8299.t35 GND 0.803901f
C4560 a_n7677_8299.n131 GND 0.320757f
C4561 a_n7677_8299.t69 GND 0.803901f
C4562 a_n7677_8299.n132 GND 0.398918f
C4563 a_n7677_8299.t20 GND 0.895722f
C4564 a_n7677_8299.n133 GND 0.382689f
C4565 a_n7677_8299.n134 GND 0.069384f
C4566 a_n7677_8299.n135 GND 0.068166f
C4567 a_n7677_8299.n136 GND 0.396278f
C4568 a_n7677_8299.n137 GND 0.320757f
C4569 a_n7677_8299.n138 GND 0.067918f
C4570 a_n7677_8299.t45 GND 0.803901f
C4571 a_n7677_8299.n139 GND 0.396531f
C4572 a_n7677_8299.n140 GND 0.320757f
C4573 a_n7677_8299.n141 GND 0.058503f
C4574 a_n7677_8299.t74 GND 0.869419f
C4575 a_n7677_8299.n142 GND 0.387049f
C4576 a_n7677_8299.n143 GND 0.138484f
C4577 a_n7677_8299.n144 GND 1.23574f
C4578 a_n7677_8299.t22 GND 0.895639f
C4579 a_n7677_8299.t78 GND 0.803901f
C4580 a_n7677_8299.t52 GND 0.803901f
C4581 a_n7677_8299.t66 GND 0.803901f
C4582 a_n7677_8299.n145 GND 0.41286f
C4583 a_n7677_8299.t60 GND 0.803901f
C4584 a_n7677_8299.t38 GND 0.803901f
C4585 a_n7677_8299.t75 GND 0.803901f
C4586 a_n7677_8299.n146 GND 0.387598f
C4587 a_n7677_8299.t44 GND 0.803901f
C4588 a_n7677_8299.n147 GND 0.320757f
C4589 a_n7677_8299.t26 GND 0.803901f
C4590 a_n7677_8299.n148 GND 0.398918f
C4591 a_n7677_8299.t58 GND 0.895722f
C4592 a_n7677_8299.n149 GND 0.382689f
C4593 a_n7677_8299.n150 GND 0.069384f
C4594 a_n7677_8299.n151 GND 0.068166f
C4595 a_n7677_8299.n152 GND 0.411298f
C4596 a_n7677_8299.n153 GND 0.411297f
C4597 a_n7677_8299.n154 GND 0.422852f
C4598 a_n7677_8299.n155 GND 0.414285f
C4599 a_n7677_8299.t47 GND 0.895639f
C4600 a_n7677_8299.t43 GND 0.803901f
C4601 a_n7677_8299.t24 GND 0.803901f
C4602 a_n7677_8299.t33 GND 0.803901f
C4603 a_n7677_8299.n156 GND 0.386699f
C4604 a_n7677_8299.t31 GND 0.803901f
C4605 a_n7677_8299.t71 GND 0.803901f
C4606 a_n7677_8299.t41 GND 0.803901f
C4607 a_n7677_8299.n157 GND 0.41286f
C4608 a_n7677_8299.t79 GND 0.803901f
C4609 a_n7677_8299.n158 GND 0.422852f
C4610 a_n7677_8299.t53 GND 0.803901f
C4611 a_n7677_8299.n159 GND 0.414272f
C4612 a_n7677_8299.t30 GND 0.895722f
C4613 a_n7677_8299.n160 GND 0.382689f
C4614 a_n7677_8299.n161 GND 0.411298f
C4615 a_n7677_8299.n162 GND 0.376234f
C4616 a_n7677_8299.n163 GND 0.059073f
C4617 a_n7677_8299.n164 GND 0.052631f
C4618 a_n7677_8299.n165 GND 0.422852f
C4619 a_n7677_8299.n166 GND 0.414285f
C4620 a_n7677_8299.n167 GND 0.702378f
C4621 a_n7677_8299.t56 GND 0.895639f
C4622 a_n7677_8299.t50 GND 0.803901f
C4623 a_n7677_8299.t64 GND 0.803901f
C4624 a_n7677_8299.t48 GND 0.803901f
C4625 a_n7677_8299.n168 GND 0.386699f
C4626 a_n7677_8299.t46 GND 0.803901f
C4627 a_n7677_8299.t59 GND 0.803901f
C4628 a_n7677_8299.t72 GND 0.803901f
C4629 a_n7677_8299.n169 GND 0.41286f
C4630 a_n7677_8299.t39 GND 0.803901f
C4631 a_n7677_8299.n170 GND 0.422852f
C4632 a_n7677_8299.t51 GND 0.803901f
C4633 a_n7677_8299.n171 GND 0.414272f
C4634 a_n7677_8299.t63 GND 0.895722f
C4635 a_n7677_8299.n172 GND 0.382689f
C4636 a_n7677_8299.n173 GND 0.411298f
C4637 a_n7677_8299.n174 GND 0.376234f
C4638 a_n7677_8299.n175 GND 0.059073f
C4639 a_n7677_8299.n176 GND 0.052631f
C4640 a_n7677_8299.n177 GND 0.422852f
C4641 a_n7677_8299.n178 GND 0.414285f
C4642 a_n7677_8299.n179 GND 1.03378f
C4643 a_n7677_8299.n180 GND 11.353001f
C4644 a_n7677_8299.n181 GND 3.69141f
C4645 a_n7677_8299.t8 GND 0.092851f
C4646 a_n7677_8299.t2 GND 0.092851f
C4647 a_n7677_8299.n182 GND 0.821619f
C4648 a_n7677_8299.n183 GND 0.751332f
C4649 a_n7677_8299.t13 GND 0.092851f
C4650 a_n7677_8299.t12 GND 0.092851f
C4651 a_n7677_8299.n184 GND 0.82046f
C4652 a_n7677_8299.n185 GND 1.98942f
C4653 a_n7677_8299.t14 GND 0.092851f
C4654 a_n7677_8299.t3 GND 0.092851f
C4655 a_n7677_8299.n186 GND 0.821619f
C4656 a_n7677_8299.n187 GND 2.10929f
C4657 a_n7677_8299.n188 GND 0.821616f
C4658 a_n7677_8299.t0 GND 0.092851f
.ends

