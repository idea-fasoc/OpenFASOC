* NGSPICE file created from diff_pair_sample_0945.ext - technology: sky130A

.subckt diff_pair_sample_0945 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=3.1239 pd=16.8 as=0 ps=0 w=8.01 l=2.16
X1 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=3.1239 pd=16.8 as=0 ps=0 w=8.01 l=2.16
X2 B.t8 B.t6 B.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=3.1239 pd=16.8 as=0 ps=0 w=8.01 l=2.16
X3 VDD2.t1 VN.t0 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=3.1239 pd=16.8 as=3.1239 ps=16.8 w=8.01 l=2.16
X4 VDD2.t0 VN.t1 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=3.1239 pd=16.8 as=3.1239 ps=16.8 w=8.01 l=2.16
X5 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=3.1239 pd=16.8 as=0 ps=0 w=8.01 l=2.16
X6 VDD1.t1 VP.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=3.1239 pd=16.8 as=3.1239 ps=16.8 w=8.01 l=2.16
X7 VDD1.t0 VP.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=3.1239 pd=16.8 as=3.1239 ps=16.8 w=8.01 l=2.16
R0 B.n401 B.n400 585
R1 B.n401 B.n44 585
R2 B.n404 B.n403 585
R3 B.n405 B.n83 585
R4 B.n407 B.n406 585
R5 B.n409 B.n82 585
R6 B.n412 B.n411 585
R7 B.n413 B.n81 585
R8 B.n415 B.n414 585
R9 B.n417 B.n80 585
R10 B.n420 B.n419 585
R11 B.n421 B.n79 585
R12 B.n423 B.n422 585
R13 B.n425 B.n78 585
R14 B.n428 B.n427 585
R15 B.n429 B.n77 585
R16 B.n431 B.n430 585
R17 B.n433 B.n76 585
R18 B.n436 B.n435 585
R19 B.n437 B.n75 585
R20 B.n439 B.n438 585
R21 B.n441 B.n74 585
R22 B.n444 B.n443 585
R23 B.n445 B.n73 585
R24 B.n447 B.n446 585
R25 B.n449 B.n72 585
R26 B.n452 B.n451 585
R27 B.n453 B.n71 585
R28 B.n455 B.n454 585
R29 B.n457 B.n70 585
R30 B.n460 B.n459 585
R31 B.n462 B.n67 585
R32 B.n464 B.n463 585
R33 B.n466 B.n66 585
R34 B.n469 B.n468 585
R35 B.n470 B.n65 585
R36 B.n472 B.n471 585
R37 B.n474 B.n64 585
R38 B.n476 B.n475 585
R39 B.n478 B.n477 585
R40 B.n481 B.n480 585
R41 B.n482 B.n59 585
R42 B.n484 B.n483 585
R43 B.n486 B.n58 585
R44 B.n489 B.n488 585
R45 B.n490 B.n57 585
R46 B.n492 B.n491 585
R47 B.n494 B.n56 585
R48 B.n497 B.n496 585
R49 B.n498 B.n55 585
R50 B.n500 B.n499 585
R51 B.n502 B.n54 585
R52 B.n505 B.n504 585
R53 B.n506 B.n53 585
R54 B.n508 B.n507 585
R55 B.n510 B.n52 585
R56 B.n513 B.n512 585
R57 B.n514 B.n51 585
R58 B.n516 B.n515 585
R59 B.n518 B.n50 585
R60 B.n521 B.n520 585
R61 B.n522 B.n49 585
R62 B.n524 B.n523 585
R63 B.n526 B.n48 585
R64 B.n529 B.n528 585
R65 B.n530 B.n47 585
R66 B.n532 B.n531 585
R67 B.n534 B.n46 585
R68 B.n537 B.n536 585
R69 B.n538 B.n45 585
R70 B.n399 B.n43 585
R71 B.n541 B.n43 585
R72 B.n398 B.n42 585
R73 B.n542 B.n42 585
R74 B.n397 B.n41 585
R75 B.n543 B.n41 585
R76 B.n396 B.n395 585
R77 B.n395 B.n37 585
R78 B.n394 B.n36 585
R79 B.n549 B.n36 585
R80 B.n393 B.n35 585
R81 B.n550 B.n35 585
R82 B.n392 B.n34 585
R83 B.n551 B.n34 585
R84 B.n391 B.n390 585
R85 B.n390 B.n30 585
R86 B.n389 B.n29 585
R87 B.n557 B.n29 585
R88 B.n388 B.n28 585
R89 B.n558 B.n28 585
R90 B.n387 B.n27 585
R91 B.n559 B.n27 585
R92 B.n386 B.n385 585
R93 B.n385 B.n23 585
R94 B.n384 B.n22 585
R95 B.n565 B.n22 585
R96 B.n383 B.n21 585
R97 B.n566 B.n21 585
R98 B.n382 B.n20 585
R99 B.n567 B.n20 585
R100 B.n381 B.n380 585
R101 B.n380 B.n16 585
R102 B.n379 B.n15 585
R103 B.n573 B.n15 585
R104 B.n378 B.n14 585
R105 B.n574 B.n14 585
R106 B.n377 B.n13 585
R107 B.n575 B.n13 585
R108 B.n376 B.n375 585
R109 B.n375 B.n12 585
R110 B.n374 B.n373 585
R111 B.n374 B.n8 585
R112 B.n372 B.n7 585
R113 B.n582 B.n7 585
R114 B.n371 B.n6 585
R115 B.n583 B.n6 585
R116 B.n370 B.n5 585
R117 B.n584 B.n5 585
R118 B.n369 B.n368 585
R119 B.n368 B.n4 585
R120 B.n367 B.n84 585
R121 B.n367 B.n366 585
R122 B.n357 B.n85 585
R123 B.n86 B.n85 585
R124 B.n359 B.n358 585
R125 B.n360 B.n359 585
R126 B.n356 B.n90 585
R127 B.n94 B.n90 585
R128 B.n355 B.n354 585
R129 B.n354 B.n353 585
R130 B.n92 B.n91 585
R131 B.n93 B.n92 585
R132 B.n346 B.n345 585
R133 B.n347 B.n346 585
R134 B.n344 B.n99 585
R135 B.n99 B.n98 585
R136 B.n343 B.n342 585
R137 B.n342 B.n341 585
R138 B.n101 B.n100 585
R139 B.n102 B.n101 585
R140 B.n334 B.n333 585
R141 B.n335 B.n334 585
R142 B.n332 B.n107 585
R143 B.n107 B.n106 585
R144 B.n331 B.n330 585
R145 B.n330 B.n329 585
R146 B.n109 B.n108 585
R147 B.n110 B.n109 585
R148 B.n322 B.n321 585
R149 B.n323 B.n322 585
R150 B.n320 B.n115 585
R151 B.n115 B.n114 585
R152 B.n319 B.n318 585
R153 B.n318 B.n317 585
R154 B.n117 B.n116 585
R155 B.n118 B.n117 585
R156 B.n310 B.n309 585
R157 B.n311 B.n310 585
R158 B.n308 B.n123 585
R159 B.n123 B.n122 585
R160 B.n307 B.n306 585
R161 B.n306 B.n305 585
R162 B.n302 B.n127 585
R163 B.n301 B.n300 585
R164 B.n298 B.n128 585
R165 B.n298 B.n126 585
R166 B.n297 B.n296 585
R167 B.n295 B.n294 585
R168 B.n293 B.n130 585
R169 B.n291 B.n290 585
R170 B.n289 B.n131 585
R171 B.n288 B.n287 585
R172 B.n285 B.n132 585
R173 B.n283 B.n282 585
R174 B.n281 B.n133 585
R175 B.n280 B.n279 585
R176 B.n277 B.n134 585
R177 B.n275 B.n274 585
R178 B.n273 B.n135 585
R179 B.n272 B.n271 585
R180 B.n269 B.n136 585
R181 B.n267 B.n266 585
R182 B.n265 B.n137 585
R183 B.n264 B.n263 585
R184 B.n261 B.n138 585
R185 B.n259 B.n258 585
R186 B.n257 B.n139 585
R187 B.n256 B.n255 585
R188 B.n253 B.n140 585
R189 B.n251 B.n250 585
R190 B.n249 B.n141 585
R191 B.n248 B.n247 585
R192 B.n245 B.n142 585
R193 B.n243 B.n242 585
R194 B.n241 B.n143 585
R195 B.n240 B.n239 585
R196 B.n237 B.n147 585
R197 B.n235 B.n234 585
R198 B.n233 B.n148 585
R199 B.n232 B.n231 585
R200 B.n229 B.n149 585
R201 B.n227 B.n226 585
R202 B.n224 B.n150 585
R203 B.n223 B.n222 585
R204 B.n220 B.n153 585
R205 B.n218 B.n217 585
R206 B.n216 B.n154 585
R207 B.n215 B.n214 585
R208 B.n212 B.n155 585
R209 B.n210 B.n209 585
R210 B.n208 B.n156 585
R211 B.n207 B.n206 585
R212 B.n204 B.n157 585
R213 B.n202 B.n201 585
R214 B.n200 B.n158 585
R215 B.n199 B.n198 585
R216 B.n196 B.n159 585
R217 B.n194 B.n193 585
R218 B.n192 B.n160 585
R219 B.n191 B.n190 585
R220 B.n188 B.n161 585
R221 B.n186 B.n185 585
R222 B.n184 B.n162 585
R223 B.n183 B.n182 585
R224 B.n180 B.n163 585
R225 B.n178 B.n177 585
R226 B.n176 B.n164 585
R227 B.n175 B.n174 585
R228 B.n172 B.n165 585
R229 B.n170 B.n169 585
R230 B.n168 B.n167 585
R231 B.n125 B.n124 585
R232 B.n304 B.n303 585
R233 B.n305 B.n304 585
R234 B.n121 B.n120 585
R235 B.n122 B.n121 585
R236 B.n313 B.n312 585
R237 B.n312 B.n311 585
R238 B.n314 B.n119 585
R239 B.n119 B.n118 585
R240 B.n316 B.n315 585
R241 B.n317 B.n316 585
R242 B.n113 B.n112 585
R243 B.n114 B.n113 585
R244 B.n325 B.n324 585
R245 B.n324 B.n323 585
R246 B.n326 B.n111 585
R247 B.n111 B.n110 585
R248 B.n328 B.n327 585
R249 B.n329 B.n328 585
R250 B.n105 B.n104 585
R251 B.n106 B.n105 585
R252 B.n337 B.n336 585
R253 B.n336 B.n335 585
R254 B.n338 B.n103 585
R255 B.n103 B.n102 585
R256 B.n340 B.n339 585
R257 B.n341 B.n340 585
R258 B.n97 B.n96 585
R259 B.n98 B.n97 585
R260 B.n349 B.n348 585
R261 B.n348 B.n347 585
R262 B.n350 B.n95 585
R263 B.n95 B.n93 585
R264 B.n352 B.n351 585
R265 B.n353 B.n352 585
R266 B.n89 B.n88 585
R267 B.n94 B.n89 585
R268 B.n362 B.n361 585
R269 B.n361 B.n360 585
R270 B.n363 B.n87 585
R271 B.n87 B.n86 585
R272 B.n365 B.n364 585
R273 B.n366 B.n365 585
R274 B.n3 B.n0 585
R275 B.n4 B.n3 585
R276 B.n581 B.n1 585
R277 B.n582 B.n581 585
R278 B.n580 B.n579 585
R279 B.n580 B.n8 585
R280 B.n578 B.n9 585
R281 B.n12 B.n9 585
R282 B.n577 B.n576 585
R283 B.n576 B.n575 585
R284 B.n11 B.n10 585
R285 B.n574 B.n11 585
R286 B.n572 B.n571 585
R287 B.n573 B.n572 585
R288 B.n570 B.n17 585
R289 B.n17 B.n16 585
R290 B.n569 B.n568 585
R291 B.n568 B.n567 585
R292 B.n19 B.n18 585
R293 B.n566 B.n19 585
R294 B.n564 B.n563 585
R295 B.n565 B.n564 585
R296 B.n562 B.n24 585
R297 B.n24 B.n23 585
R298 B.n561 B.n560 585
R299 B.n560 B.n559 585
R300 B.n26 B.n25 585
R301 B.n558 B.n26 585
R302 B.n556 B.n555 585
R303 B.n557 B.n556 585
R304 B.n554 B.n31 585
R305 B.n31 B.n30 585
R306 B.n553 B.n552 585
R307 B.n552 B.n551 585
R308 B.n33 B.n32 585
R309 B.n550 B.n33 585
R310 B.n548 B.n547 585
R311 B.n549 B.n548 585
R312 B.n546 B.n38 585
R313 B.n38 B.n37 585
R314 B.n545 B.n544 585
R315 B.n544 B.n543 585
R316 B.n40 B.n39 585
R317 B.n542 B.n40 585
R318 B.n540 B.n539 585
R319 B.n541 B.n540 585
R320 B.n585 B.n584 585
R321 B.n583 B.n2 585
R322 B.n540 B.n45 569.379
R323 B.n401 B.n43 569.379
R324 B.n306 B.n125 569.379
R325 B.n304 B.n127 569.379
R326 B.n60 B.t6 296.642
R327 B.n68 B.t2 296.642
R328 B.n151 B.t13 296.642
R329 B.n144 B.t9 296.642
R330 B.n68 B.t4 261.776
R331 B.n151 B.t15 261.776
R332 B.n60 B.t7 261.776
R333 B.n144 B.t12 261.776
R334 B.n402 B.n44 256.663
R335 B.n408 B.n44 256.663
R336 B.n410 B.n44 256.663
R337 B.n416 B.n44 256.663
R338 B.n418 B.n44 256.663
R339 B.n424 B.n44 256.663
R340 B.n426 B.n44 256.663
R341 B.n432 B.n44 256.663
R342 B.n434 B.n44 256.663
R343 B.n440 B.n44 256.663
R344 B.n442 B.n44 256.663
R345 B.n448 B.n44 256.663
R346 B.n450 B.n44 256.663
R347 B.n456 B.n44 256.663
R348 B.n458 B.n44 256.663
R349 B.n465 B.n44 256.663
R350 B.n467 B.n44 256.663
R351 B.n473 B.n44 256.663
R352 B.n63 B.n44 256.663
R353 B.n479 B.n44 256.663
R354 B.n485 B.n44 256.663
R355 B.n487 B.n44 256.663
R356 B.n493 B.n44 256.663
R357 B.n495 B.n44 256.663
R358 B.n501 B.n44 256.663
R359 B.n503 B.n44 256.663
R360 B.n509 B.n44 256.663
R361 B.n511 B.n44 256.663
R362 B.n517 B.n44 256.663
R363 B.n519 B.n44 256.663
R364 B.n525 B.n44 256.663
R365 B.n527 B.n44 256.663
R366 B.n533 B.n44 256.663
R367 B.n535 B.n44 256.663
R368 B.n299 B.n126 256.663
R369 B.n129 B.n126 256.663
R370 B.n292 B.n126 256.663
R371 B.n286 B.n126 256.663
R372 B.n284 B.n126 256.663
R373 B.n278 B.n126 256.663
R374 B.n276 B.n126 256.663
R375 B.n270 B.n126 256.663
R376 B.n268 B.n126 256.663
R377 B.n262 B.n126 256.663
R378 B.n260 B.n126 256.663
R379 B.n254 B.n126 256.663
R380 B.n252 B.n126 256.663
R381 B.n246 B.n126 256.663
R382 B.n244 B.n126 256.663
R383 B.n238 B.n126 256.663
R384 B.n236 B.n126 256.663
R385 B.n230 B.n126 256.663
R386 B.n228 B.n126 256.663
R387 B.n221 B.n126 256.663
R388 B.n219 B.n126 256.663
R389 B.n213 B.n126 256.663
R390 B.n211 B.n126 256.663
R391 B.n205 B.n126 256.663
R392 B.n203 B.n126 256.663
R393 B.n197 B.n126 256.663
R394 B.n195 B.n126 256.663
R395 B.n189 B.n126 256.663
R396 B.n187 B.n126 256.663
R397 B.n181 B.n126 256.663
R398 B.n179 B.n126 256.663
R399 B.n173 B.n126 256.663
R400 B.n171 B.n126 256.663
R401 B.n166 B.n126 256.663
R402 B.n587 B.n586 256.663
R403 B.n69 B.t5 213.486
R404 B.n152 B.t14 213.486
R405 B.n61 B.t8 213.486
R406 B.n145 B.t11 213.486
R407 B.n536 B.n534 163.367
R408 B.n532 B.n47 163.367
R409 B.n528 B.n526 163.367
R410 B.n524 B.n49 163.367
R411 B.n520 B.n518 163.367
R412 B.n516 B.n51 163.367
R413 B.n512 B.n510 163.367
R414 B.n508 B.n53 163.367
R415 B.n504 B.n502 163.367
R416 B.n500 B.n55 163.367
R417 B.n496 B.n494 163.367
R418 B.n492 B.n57 163.367
R419 B.n488 B.n486 163.367
R420 B.n484 B.n59 163.367
R421 B.n480 B.n478 163.367
R422 B.n475 B.n474 163.367
R423 B.n472 B.n65 163.367
R424 B.n468 B.n466 163.367
R425 B.n464 B.n67 163.367
R426 B.n459 B.n457 163.367
R427 B.n455 B.n71 163.367
R428 B.n451 B.n449 163.367
R429 B.n447 B.n73 163.367
R430 B.n443 B.n441 163.367
R431 B.n439 B.n75 163.367
R432 B.n435 B.n433 163.367
R433 B.n431 B.n77 163.367
R434 B.n427 B.n425 163.367
R435 B.n423 B.n79 163.367
R436 B.n419 B.n417 163.367
R437 B.n415 B.n81 163.367
R438 B.n411 B.n409 163.367
R439 B.n407 B.n83 163.367
R440 B.n403 B.n401 163.367
R441 B.n306 B.n123 163.367
R442 B.n310 B.n123 163.367
R443 B.n310 B.n117 163.367
R444 B.n318 B.n117 163.367
R445 B.n318 B.n115 163.367
R446 B.n322 B.n115 163.367
R447 B.n322 B.n109 163.367
R448 B.n330 B.n109 163.367
R449 B.n330 B.n107 163.367
R450 B.n334 B.n107 163.367
R451 B.n334 B.n101 163.367
R452 B.n342 B.n101 163.367
R453 B.n342 B.n99 163.367
R454 B.n346 B.n99 163.367
R455 B.n346 B.n92 163.367
R456 B.n354 B.n92 163.367
R457 B.n354 B.n90 163.367
R458 B.n359 B.n90 163.367
R459 B.n359 B.n85 163.367
R460 B.n367 B.n85 163.367
R461 B.n368 B.n367 163.367
R462 B.n368 B.n5 163.367
R463 B.n6 B.n5 163.367
R464 B.n7 B.n6 163.367
R465 B.n374 B.n7 163.367
R466 B.n375 B.n374 163.367
R467 B.n375 B.n13 163.367
R468 B.n14 B.n13 163.367
R469 B.n15 B.n14 163.367
R470 B.n380 B.n15 163.367
R471 B.n380 B.n20 163.367
R472 B.n21 B.n20 163.367
R473 B.n22 B.n21 163.367
R474 B.n385 B.n22 163.367
R475 B.n385 B.n27 163.367
R476 B.n28 B.n27 163.367
R477 B.n29 B.n28 163.367
R478 B.n390 B.n29 163.367
R479 B.n390 B.n34 163.367
R480 B.n35 B.n34 163.367
R481 B.n36 B.n35 163.367
R482 B.n395 B.n36 163.367
R483 B.n395 B.n41 163.367
R484 B.n42 B.n41 163.367
R485 B.n43 B.n42 163.367
R486 B.n300 B.n298 163.367
R487 B.n298 B.n297 163.367
R488 B.n294 B.n293 163.367
R489 B.n291 B.n131 163.367
R490 B.n287 B.n285 163.367
R491 B.n283 B.n133 163.367
R492 B.n279 B.n277 163.367
R493 B.n275 B.n135 163.367
R494 B.n271 B.n269 163.367
R495 B.n267 B.n137 163.367
R496 B.n263 B.n261 163.367
R497 B.n259 B.n139 163.367
R498 B.n255 B.n253 163.367
R499 B.n251 B.n141 163.367
R500 B.n247 B.n245 163.367
R501 B.n243 B.n143 163.367
R502 B.n239 B.n237 163.367
R503 B.n235 B.n148 163.367
R504 B.n231 B.n229 163.367
R505 B.n227 B.n150 163.367
R506 B.n222 B.n220 163.367
R507 B.n218 B.n154 163.367
R508 B.n214 B.n212 163.367
R509 B.n210 B.n156 163.367
R510 B.n206 B.n204 163.367
R511 B.n202 B.n158 163.367
R512 B.n198 B.n196 163.367
R513 B.n194 B.n160 163.367
R514 B.n190 B.n188 163.367
R515 B.n186 B.n162 163.367
R516 B.n182 B.n180 163.367
R517 B.n178 B.n164 163.367
R518 B.n174 B.n172 163.367
R519 B.n170 B.n167 163.367
R520 B.n304 B.n121 163.367
R521 B.n312 B.n121 163.367
R522 B.n312 B.n119 163.367
R523 B.n316 B.n119 163.367
R524 B.n316 B.n113 163.367
R525 B.n324 B.n113 163.367
R526 B.n324 B.n111 163.367
R527 B.n328 B.n111 163.367
R528 B.n328 B.n105 163.367
R529 B.n336 B.n105 163.367
R530 B.n336 B.n103 163.367
R531 B.n340 B.n103 163.367
R532 B.n340 B.n97 163.367
R533 B.n348 B.n97 163.367
R534 B.n348 B.n95 163.367
R535 B.n352 B.n95 163.367
R536 B.n352 B.n89 163.367
R537 B.n361 B.n89 163.367
R538 B.n361 B.n87 163.367
R539 B.n365 B.n87 163.367
R540 B.n365 B.n3 163.367
R541 B.n585 B.n3 163.367
R542 B.n581 B.n2 163.367
R543 B.n581 B.n580 163.367
R544 B.n580 B.n9 163.367
R545 B.n576 B.n9 163.367
R546 B.n576 B.n11 163.367
R547 B.n572 B.n11 163.367
R548 B.n572 B.n17 163.367
R549 B.n568 B.n17 163.367
R550 B.n568 B.n19 163.367
R551 B.n564 B.n19 163.367
R552 B.n564 B.n24 163.367
R553 B.n560 B.n24 163.367
R554 B.n560 B.n26 163.367
R555 B.n556 B.n26 163.367
R556 B.n556 B.n31 163.367
R557 B.n552 B.n31 163.367
R558 B.n552 B.n33 163.367
R559 B.n548 B.n33 163.367
R560 B.n548 B.n38 163.367
R561 B.n544 B.n38 163.367
R562 B.n544 B.n40 163.367
R563 B.n540 B.n40 163.367
R564 B.n305 B.n126 116.749
R565 B.n541 B.n44 116.749
R566 B.n535 B.n45 71.676
R567 B.n534 B.n533 71.676
R568 B.n527 B.n47 71.676
R569 B.n526 B.n525 71.676
R570 B.n519 B.n49 71.676
R571 B.n518 B.n517 71.676
R572 B.n511 B.n51 71.676
R573 B.n510 B.n509 71.676
R574 B.n503 B.n53 71.676
R575 B.n502 B.n501 71.676
R576 B.n495 B.n55 71.676
R577 B.n494 B.n493 71.676
R578 B.n487 B.n57 71.676
R579 B.n486 B.n485 71.676
R580 B.n479 B.n59 71.676
R581 B.n478 B.n63 71.676
R582 B.n474 B.n473 71.676
R583 B.n467 B.n65 71.676
R584 B.n466 B.n465 71.676
R585 B.n458 B.n67 71.676
R586 B.n457 B.n456 71.676
R587 B.n450 B.n71 71.676
R588 B.n449 B.n448 71.676
R589 B.n442 B.n73 71.676
R590 B.n441 B.n440 71.676
R591 B.n434 B.n75 71.676
R592 B.n433 B.n432 71.676
R593 B.n426 B.n77 71.676
R594 B.n425 B.n424 71.676
R595 B.n418 B.n79 71.676
R596 B.n417 B.n416 71.676
R597 B.n410 B.n81 71.676
R598 B.n409 B.n408 71.676
R599 B.n402 B.n83 71.676
R600 B.n403 B.n402 71.676
R601 B.n408 B.n407 71.676
R602 B.n411 B.n410 71.676
R603 B.n416 B.n415 71.676
R604 B.n419 B.n418 71.676
R605 B.n424 B.n423 71.676
R606 B.n427 B.n426 71.676
R607 B.n432 B.n431 71.676
R608 B.n435 B.n434 71.676
R609 B.n440 B.n439 71.676
R610 B.n443 B.n442 71.676
R611 B.n448 B.n447 71.676
R612 B.n451 B.n450 71.676
R613 B.n456 B.n455 71.676
R614 B.n459 B.n458 71.676
R615 B.n465 B.n464 71.676
R616 B.n468 B.n467 71.676
R617 B.n473 B.n472 71.676
R618 B.n475 B.n63 71.676
R619 B.n480 B.n479 71.676
R620 B.n485 B.n484 71.676
R621 B.n488 B.n487 71.676
R622 B.n493 B.n492 71.676
R623 B.n496 B.n495 71.676
R624 B.n501 B.n500 71.676
R625 B.n504 B.n503 71.676
R626 B.n509 B.n508 71.676
R627 B.n512 B.n511 71.676
R628 B.n517 B.n516 71.676
R629 B.n520 B.n519 71.676
R630 B.n525 B.n524 71.676
R631 B.n528 B.n527 71.676
R632 B.n533 B.n532 71.676
R633 B.n536 B.n535 71.676
R634 B.n299 B.n127 71.676
R635 B.n297 B.n129 71.676
R636 B.n293 B.n292 71.676
R637 B.n286 B.n131 71.676
R638 B.n285 B.n284 71.676
R639 B.n278 B.n133 71.676
R640 B.n277 B.n276 71.676
R641 B.n270 B.n135 71.676
R642 B.n269 B.n268 71.676
R643 B.n262 B.n137 71.676
R644 B.n261 B.n260 71.676
R645 B.n254 B.n139 71.676
R646 B.n253 B.n252 71.676
R647 B.n246 B.n141 71.676
R648 B.n245 B.n244 71.676
R649 B.n238 B.n143 71.676
R650 B.n237 B.n236 71.676
R651 B.n230 B.n148 71.676
R652 B.n229 B.n228 71.676
R653 B.n221 B.n150 71.676
R654 B.n220 B.n219 71.676
R655 B.n213 B.n154 71.676
R656 B.n212 B.n211 71.676
R657 B.n205 B.n156 71.676
R658 B.n204 B.n203 71.676
R659 B.n197 B.n158 71.676
R660 B.n196 B.n195 71.676
R661 B.n189 B.n160 71.676
R662 B.n188 B.n187 71.676
R663 B.n181 B.n162 71.676
R664 B.n180 B.n179 71.676
R665 B.n173 B.n164 71.676
R666 B.n172 B.n171 71.676
R667 B.n167 B.n166 71.676
R668 B.n300 B.n299 71.676
R669 B.n294 B.n129 71.676
R670 B.n292 B.n291 71.676
R671 B.n287 B.n286 71.676
R672 B.n284 B.n283 71.676
R673 B.n279 B.n278 71.676
R674 B.n276 B.n275 71.676
R675 B.n271 B.n270 71.676
R676 B.n268 B.n267 71.676
R677 B.n263 B.n262 71.676
R678 B.n260 B.n259 71.676
R679 B.n255 B.n254 71.676
R680 B.n252 B.n251 71.676
R681 B.n247 B.n246 71.676
R682 B.n244 B.n243 71.676
R683 B.n239 B.n238 71.676
R684 B.n236 B.n235 71.676
R685 B.n231 B.n230 71.676
R686 B.n228 B.n227 71.676
R687 B.n222 B.n221 71.676
R688 B.n219 B.n218 71.676
R689 B.n214 B.n213 71.676
R690 B.n211 B.n210 71.676
R691 B.n206 B.n205 71.676
R692 B.n203 B.n202 71.676
R693 B.n198 B.n197 71.676
R694 B.n195 B.n194 71.676
R695 B.n190 B.n189 71.676
R696 B.n187 B.n186 71.676
R697 B.n182 B.n181 71.676
R698 B.n179 B.n178 71.676
R699 B.n174 B.n173 71.676
R700 B.n171 B.n170 71.676
R701 B.n166 B.n125 71.676
R702 B.n586 B.n585 71.676
R703 B.n586 B.n2 71.676
R704 B.n62 B.n61 59.5399
R705 B.n461 B.n69 59.5399
R706 B.n225 B.n152 59.5399
R707 B.n146 B.n145 59.5399
R708 B.n305 B.n122 56.3046
R709 B.n311 B.n122 56.3046
R710 B.n311 B.n118 56.3046
R711 B.n317 B.n118 56.3046
R712 B.n317 B.n114 56.3046
R713 B.n323 B.n114 56.3046
R714 B.n329 B.n110 56.3046
R715 B.n329 B.n106 56.3046
R716 B.n335 B.n106 56.3046
R717 B.n335 B.n102 56.3046
R718 B.n341 B.n102 56.3046
R719 B.n341 B.n98 56.3046
R720 B.n347 B.n98 56.3046
R721 B.n347 B.n93 56.3046
R722 B.n353 B.n93 56.3046
R723 B.n353 B.n94 56.3046
R724 B.n360 B.n86 56.3046
R725 B.n366 B.n86 56.3046
R726 B.n366 B.n4 56.3046
R727 B.n584 B.n4 56.3046
R728 B.n584 B.n583 56.3046
R729 B.n583 B.n582 56.3046
R730 B.n582 B.n8 56.3046
R731 B.n12 B.n8 56.3046
R732 B.n575 B.n12 56.3046
R733 B.n574 B.n573 56.3046
R734 B.n573 B.n16 56.3046
R735 B.n567 B.n16 56.3046
R736 B.n567 B.n566 56.3046
R737 B.n566 B.n565 56.3046
R738 B.n565 B.n23 56.3046
R739 B.n559 B.n23 56.3046
R740 B.n559 B.n558 56.3046
R741 B.n558 B.n557 56.3046
R742 B.n557 B.n30 56.3046
R743 B.n551 B.n550 56.3046
R744 B.n550 B.n549 56.3046
R745 B.n549 B.n37 56.3046
R746 B.n543 B.n37 56.3046
R747 B.n543 B.n542 56.3046
R748 B.n542 B.n541 56.3046
R749 B.n61 B.n60 48.2914
R750 B.n69 B.n68 48.2914
R751 B.n152 B.n151 48.2914
R752 B.n145 B.n144 48.2914
R753 B.n360 B.t1 43.0566
R754 B.n575 B.t0 43.0566
R755 B.n323 B.t10 39.7446
R756 B.n551 B.t3 39.7446
R757 B.n303 B.n302 36.9956
R758 B.n307 B.n124 36.9956
R759 B.n400 B.n399 36.9956
R760 B.n539 B.n538 36.9956
R761 B B.n587 18.0485
R762 B.t10 B.n110 16.5605
R763 B.t3 B.n30 16.5605
R764 B.n94 B.t1 13.2485
R765 B.t0 B.n574 13.2485
R766 B.n303 B.n120 10.6151
R767 B.n313 B.n120 10.6151
R768 B.n314 B.n313 10.6151
R769 B.n315 B.n314 10.6151
R770 B.n315 B.n112 10.6151
R771 B.n325 B.n112 10.6151
R772 B.n326 B.n325 10.6151
R773 B.n327 B.n326 10.6151
R774 B.n327 B.n104 10.6151
R775 B.n337 B.n104 10.6151
R776 B.n338 B.n337 10.6151
R777 B.n339 B.n338 10.6151
R778 B.n339 B.n96 10.6151
R779 B.n349 B.n96 10.6151
R780 B.n350 B.n349 10.6151
R781 B.n351 B.n350 10.6151
R782 B.n351 B.n88 10.6151
R783 B.n362 B.n88 10.6151
R784 B.n363 B.n362 10.6151
R785 B.n364 B.n363 10.6151
R786 B.n364 B.n0 10.6151
R787 B.n302 B.n301 10.6151
R788 B.n301 B.n128 10.6151
R789 B.n296 B.n128 10.6151
R790 B.n296 B.n295 10.6151
R791 B.n295 B.n130 10.6151
R792 B.n290 B.n130 10.6151
R793 B.n290 B.n289 10.6151
R794 B.n289 B.n288 10.6151
R795 B.n288 B.n132 10.6151
R796 B.n282 B.n132 10.6151
R797 B.n282 B.n281 10.6151
R798 B.n281 B.n280 10.6151
R799 B.n280 B.n134 10.6151
R800 B.n274 B.n134 10.6151
R801 B.n274 B.n273 10.6151
R802 B.n273 B.n272 10.6151
R803 B.n272 B.n136 10.6151
R804 B.n266 B.n136 10.6151
R805 B.n266 B.n265 10.6151
R806 B.n265 B.n264 10.6151
R807 B.n264 B.n138 10.6151
R808 B.n258 B.n138 10.6151
R809 B.n258 B.n257 10.6151
R810 B.n257 B.n256 10.6151
R811 B.n256 B.n140 10.6151
R812 B.n250 B.n140 10.6151
R813 B.n250 B.n249 10.6151
R814 B.n249 B.n248 10.6151
R815 B.n248 B.n142 10.6151
R816 B.n242 B.n241 10.6151
R817 B.n241 B.n240 10.6151
R818 B.n240 B.n147 10.6151
R819 B.n234 B.n147 10.6151
R820 B.n234 B.n233 10.6151
R821 B.n233 B.n232 10.6151
R822 B.n232 B.n149 10.6151
R823 B.n226 B.n149 10.6151
R824 B.n224 B.n223 10.6151
R825 B.n223 B.n153 10.6151
R826 B.n217 B.n153 10.6151
R827 B.n217 B.n216 10.6151
R828 B.n216 B.n215 10.6151
R829 B.n215 B.n155 10.6151
R830 B.n209 B.n155 10.6151
R831 B.n209 B.n208 10.6151
R832 B.n208 B.n207 10.6151
R833 B.n207 B.n157 10.6151
R834 B.n201 B.n157 10.6151
R835 B.n201 B.n200 10.6151
R836 B.n200 B.n199 10.6151
R837 B.n199 B.n159 10.6151
R838 B.n193 B.n159 10.6151
R839 B.n193 B.n192 10.6151
R840 B.n192 B.n191 10.6151
R841 B.n191 B.n161 10.6151
R842 B.n185 B.n161 10.6151
R843 B.n185 B.n184 10.6151
R844 B.n184 B.n183 10.6151
R845 B.n183 B.n163 10.6151
R846 B.n177 B.n163 10.6151
R847 B.n177 B.n176 10.6151
R848 B.n176 B.n175 10.6151
R849 B.n175 B.n165 10.6151
R850 B.n169 B.n165 10.6151
R851 B.n169 B.n168 10.6151
R852 B.n168 B.n124 10.6151
R853 B.n308 B.n307 10.6151
R854 B.n309 B.n308 10.6151
R855 B.n309 B.n116 10.6151
R856 B.n319 B.n116 10.6151
R857 B.n320 B.n319 10.6151
R858 B.n321 B.n320 10.6151
R859 B.n321 B.n108 10.6151
R860 B.n331 B.n108 10.6151
R861 B.n332 B.n331 10.6151
R862 B.n333 B.n332 10.6151
R863 B.n333 B.n100 10.6151
R864 B.n343 B.n100 10.6151
R865 B.n344 B.n343 10.6151
R866 B.n345 B.n344 10.6151
R867 B.n345 B.n91 10.6151
R868 B.n355 B.n91 10.6151
R869 B.n356 B.n355 10.6151
R870 B.n358 B.n356 10.6151
R871 B.n358 B.n357 10.6151
R872 B.n357 B.n84 10.6151
R873 B.n369 B.n84 10.6151
R874 B.n370 B.n369 10.6151
R875 B.n371 B.n370 10.6151
R876 B.n372 B.n371 10.6151
R877 B.n373 B.n372 10.6151
R878 B.n376 B.n373 10.6151
R879 B.n377 B.n376 10.6151
R880 B.n378 B.n377 10.6151
R881 B.n379 B.n378 10.6151
R882 B.n381 B.n379 10.6151
R883 B.n382 B.n381 10.6151
R884 B.n383 B.n382 10.6151
R885 B.n384 B.n383 10.6151
R886 B.n386 B.n384 10.6151
R887 B.n387 B.n386 10.6151
R888 B.n388 B.n387 10.6151
R889 B.n389 B.n388 10.6151
R890 B.n391 B.n389 10.6151
R891 B.n392 B.n391 10.6151
R892 B.n393 B.n392 10.6151
R893 B.n394 B.n393 10.6151
R894 B.n396 B.n394 10.6151
R895 B.n397 B.n396 10.6151
R896 B.n398 B.n397 10.6151
R897 B.n399 B.n398 10.6151
R898 B.n579 B.n1 10.6151
R899 B.n579 B.n578 10.6151
R900 B.n578 B.n577 10.6151
R901 B.n577 B.n10 10.6151
R902 B.n571 B.n10 10.6151
R903 B.n571 B.n570 10.6151
R904 B.n570 B.n569 10.6151
R905 B.n569 B.n18 10.6151
R906 B.n563 B.n18 10.6151
R907 B.n563 B.n562 10.6151
R908 B.n562 B.n561 10.6151
R909 B.n561 B.n25 10.6151
R910 B.n555 B.n25 10.6151
R911 B.n555 B.n554 10.6151
R912 B.n554 B.n553 10.6151
R913 B.n553 B.n32 10.6151
R914 B.n547 B.n32 10.6151
R915 B.n547 B.n546 10.6151
R916 B.n546 B.n545 10.6151
R917 B.n545 B.n39 10.6151
R918 B.n539 B.n39 10.6151
R919 B.n538 B.n537 10.6151
R920 B.n537 B.n46 10.6151
R921 B.n531 B.n46 10.6151
R922 B.n531 B.n530 10.6151
R923 B.n530 B.n529 10.6151
R924 B.n529 B.n48 10.6151
R925 B.n523 B.n48 10.6151
R926 B.n523 B.n522 10.6151
R927 B.n522 B.n521 10.6151
R928 B.n521 B.n50 10.6151
R929 B.n515 B.n50 10.6151
R930 B.n515 B.n514 10.6151
R931 B.n514 B.n513 10.6151
R932 B.n513 B.n52 10.6151
R933 B.n507 B.n52 10.6151
R934 B.n507 B.n506 10.6151
R935 B.n506 B.n505 10.6151
R936 B.n505 B.n54 10.6151
R937 B.n499 B.n54 10.6151
R938 B.n499 B.n498 10.6151
R939 B.n498 B.n497 10.6151
R940 B.n497 B.n56 10.6151
R941 B.n491 B.n56 10.6151
R942 B.n491 B.n490 10.6151
R943 B.n490 B.n489 10.6151
R944 B.n489 B.n58 10.6151
R945 B.n483 B.n58 10.6151
R946 B.n483 B.n482 10.6151
R947 B.n482 B.n481 10.6151
R948 B.n477 B.n476 10.6151
R949 B.n476 B.n64 10.6151
R950 B.n471 B.n64 10.6151
R951 B.n471 B.n470 10.6151
R952 B.n470 B.n469 10.6151
R953 B.n469 B.n66 10.6151
R954 B.n463 B.n66 10.6151
R955 B.n463 B.n462 10.6151
R956 B.n460 B.n70 10.6151
R957 B.n454 B.n70 10.6151
R958 B.n454 B.n453 10.6151
R959 B.n453 B.n452 10.6151
R960 B.n452 B.n72 10.6151
R961 B.n446 B.n72 10.6151
R962 B.n446 B.n445 10.6151
R963 B.n445 B.n444 10.6151
R964 B.n444 B.n74 10.6151
R965 B.n438 B.n74 10.6151
R966 B.n438 B.n437 10.6151
R967 B.n437 B.n436 10.6151
R968 B.n436 B.n76 10.6151
R969 B.n430 B.n76 10.6151
R970 B.n430 B.n429 10.6151
R971 B.n429 B.n428 10.6151
R972 B.n428 B.n78 10.6151
R973 B.n422 B.n78 10.6151
R974 B.n422 B.n421 10.6151
R975 B.n421 B.n420 10.6151
R976 B.n420 B.n80 10.6151
R977 B.n414 B.n80 10.6151
R978 B.n414 B.n413 10.6151
R979 B.n413 B.n412 10.6151
R980 B.n412 B.n82 10.6151
R981 B.n406 B.n82 10.6151
R982 B.n406 B.n405 10.6151
R983 B.n405 B.n404 10.6151
R984 B.n404 B.n400 10.6151
R985 B.n587 B.n0 8.11757
R986 B.n587 B.n1 8.11757
R987 B.n242 B.n146 6.5566
R988 B.n226 B.n225 6.5566
R989 B.n477 B.n62 6.5566
R990 B.n462 B.n461 6.5566
R991 B.n146 B.n142 4.05904
R992 B.n225 B.n224 4.05904
R993 B.n481 B.n62 4.05904
R994 B.n461 B.n460 4.05904
R995 VN VN.t1 179.106
R996 VN VN.t0 138.877
R997 VTAIL.n162 VTAIL.n126 289.615
R998 VTAIL.n36 VTAIL.n0 289.615
R999 VTAIL.n120 VTAIL.n84 289.615
R1000 VTAIL.n78 VTAIL.n42 289.615
R1001 VTAIL.n138 VTAIL.n137 185
R1002 VTAIL.n143 VTAIL.n142 185
R1003 VTAIL.n145 VTAIL.n144 185
R1004 VTAIL.n134 VTAIL.n133 185
R1005 VTAIL.n151 VTAIL.n150 185
R1006 VTAIL.n153 VTAIL.n152 185
R1007 VTAIL.n130 VTAIL.n129 185
R1008 VTAIL.n160 VTAIL.n159 185
R1009 VTAIL.n161 VTAIL.n128 185
R1010 VTAIL.n163 VTAIL.n162 185
R1011 VTAIL.n12 VTAIL.n11 185
R1012 VTAIL.n17 VTAIL.n16 185
R1013 VTAIL.n19 VTAIL.n18 185
R1014 VTAIL.n8 VTAIL.n7 185
R1015 VTAIL.n25 VTAIL.n24 185
R1016 VTAIL.n27 VTAIL.n26 185
R1017 VTAIL.n4 VTAIL.n3 185
R1018 VTAIL.n34 VTAIL.n33 185
R1019 VTAIL.n35 VTAIL.n2 185
R1020 VTAIL.n37 VTAIL.n36 185
R1021 VTAIL.n121 VTAIL.n120 185
R1022 VTAIL.n119 VTAIL.n86 185
R1023 VTAIL.n118 VTAIL.n117 185
R1024 VTAIL.n89 VTAIL.n87 185
R1025 VTAIL.n112 VTAIL.n111 185
R1026 VTAIL.n110 VTAIL.n109 185
R1027 VTAIL.n93 VTAIL.n92 185
R1028 VTAIL.n104 VTAIL.n103 185
R1029 VTAIL.n102 VTAIL.n101 185
R1030 VTAIL.n97 VTAIL.n96 185
R1031 VTAIL.n79 VTAIL.n78 185
R1032 VTAIL.n77 VTAIL.n44 185
R1033 VTAIL.n76 VTAIL.n75 185
R1034 VTAIL.n47 VTAIL.n45 185
R1035 VTAIL.n70 VTAIL.n69 185
R1036 VTAIL.n68 VTAIL.n67 185
R1037 VTAIL.n51 VTAIL.n50 185
R1038 VTAIL.n62 VTAIL.n61 185
R1039 VTAIL.n60 VTAIL.n59 185
R1040 VTAIL.n55 VTAIL.n54 185
R1041 VTAIL.n139 VTAIL.t2 149.524
R1042 VTAIL.n13 VTAIL.t1 149.524
R1043 VTAIL.n98 VTAIL.t0 149.524
R1044 VTAIL.n56 VTAIL.t3 149.524
R1045 VTAIL.n143 VTAIL.n137 104.615
R1046 VTAIL.n144 VTAIL.n143 104.615
R1047 VTAIL.n144 VTAIL.n133 104.615
R1048 VTAIL.n151 VTAIL.n133 104.615
R1049 VTAIL.n152 VTAIL.n151 104.615
R1050 VTAIL.n152 VTAIL.n129 104.615
R1051 VTAIL.n160 VTAIL.n129 104.615
R1052 VTAIL.n161 VTAIL.n160 104.615
R1053 VTAIL.n162 VTAIL.n161 104.615
R1054 VTAIL.n17 VTAIL.n11 104.615
R1055 VTAIL.n18 VTAIL.n17 104.615
R1056 VTAIL.n18 VTAIL.n7 104.615
R1057 VTAIL.n25 VTAIL.n7 104.615
R1058 VTAIL.n26 VTAIL.n25 104.615
R1059 VTAIL.n26 VTAIL.n3 104.615
R1060 VTAIL.n34 VTAIL.n3 104.615
R1061 VTAIL.n35 VTAIL.n34 104.615
R1062 VTAIL.n36 VTAIL.n35 104.615
R1063 VTAIL.n120 VTAIL.n119 104.615
R1064 VTAIL.n119 VTAIL.n118 104.615
R1065 VTAIL.n118 VTAIL.n87 104.615
R1066 VTAIL.n111 VTAIL.n87 104.615
R1067 VTAIL.n111 VTAIL.n110 104.615
R1068 VTAIL.n110 VTAIL.n92 104.615
R1069 VTAIL.n103 VTAIL.n92 104.615
R1070 VTAIL.n103 VTAIL.n102 104.615
R1071 VTAIL.n102 VTAIL.n96 104.615
R1072 VTAIL.n78 VTAIL.n77 104.615
R1073 VTAIL.n77 VTAIL.n76 104.615
R1074 VTAIL.n76 VTAIL.n45 104.615
R1075 VTAIL.n69 VTAIL.n45 104.615
R1076 VTAIL.n69 VTAIL.n68 104.615
R1077 VTAIL.n68 VTAIL.n50 104.615
R1078 VTAIL.n61 VTAIL.n50 104.615
R1079 VTAIL.n61 VTAIL.n60 104.615
R1080 VTAIL.n60 VTAIL.n54 104.615
R1081 VTAIL.t2 VTAIL.n137 52.3082
R1082 VTAIL.t1 VTAIL.n11 52.3082
R1083 VTAIL.t0 VTAIL.n96 52.3082
R1084 VTAIL.t3 VTAIL.n54 52.3082
R1085 VTAIL.n167 VTAIL.n166 36.2581
R1086 VTAIL.n41 VTAIL.n40 36.2581
R1087 VTAIL.n125 VTAIL.n124 36.2581
R1088 VTAIL.n83 VTAIL.n82 36.2581
R1089 VTAIL.n83 VTAIL.n41 23.5652
R1090 VTAIL.n167 VTAIL.n125 21.4186
R1091 VTAIL.n163 VTAIL.n128 13.1884
R1092 VTAIL.n37 VTAIL.n2 13.1884
R1093 VTAIL.n121 VTAIL.n86 13.1884
R1094 VTAIL.n79 VTAIL.n44 13.1884
R1095 VTAIL.n159 VTAIL.n158 12.8005
R1096 VTAIL.n164 VTAIL.n126 12.8005
R1097 VTAIL.n33 VTAIL.n32 12.8005
R1098 VTAIL.n38 VTAIL.n0 12.8005
R1099 VTAIL.n122 VTAIL.n84 12.8005
R1100 VTAIL.n117 VTAIL.n88 12.8005
R1101 VTAIL.n80 VTAIL.n42 12.8005
R1102 VTAIL.n75 VTAIL.n46 12.8005
R1103 VTAIL.n157 VTAIL.n130 12.0247
R1104 VTAIL.n31 VTAIL.n4 12.0247
R1105 VTAIL.n116 VTAIL.n89 12.0247
R1106 VTAIL.n74 VTAIL.n47 12.0247
R1107 VTAIL.n154 VTAIL.n153 11.249
R1108 VTAIL.n28 VTAIL.n27 11.249
R1109 VTAIL.n113 VTAIL.n112 11.249
R1110 VTAIL.n71 VTAIL.n70 11.249
R1111 VTAIL.n150 VTAIL.n132 10.4732
R1112 VTAIL.n24 VTAIL.n6 10.4732
R1113 VTAIL.n109 VTAIL.n91 10.4732
R1114 VTAIL.n67 VTAIL.n49 10.4732
R1115 VTAIL.n139 VTAIL.n138 10.2747
R1116 VTAIL.n13 VTAIL.n12 10.2747
R1117 VTAIL.n98 VTAIL.n97 10.2747
R1118 VTAIL.n56 VTAIL.n55 10.2747
R1119 VTAIL.n149 VTAIL.n134 9.69747
R1120 VTAIL.n23 VTAIL.n8 9.69747
R1121 VTAIL.n108 VTAIL.n93 9.69747
R1122 VTAIL.n66 VTAIL.n51 9.69747
R1123 VTAIL.n166 VTAIL.n165 9.45567
R1124 VTAIL.n40 VTAIL.n39 9.45567
R1125 VTAIL.n124 VTAIL.n123 9.45567
R1126 VTAIL.n82 VTAIL.n81 9.45567
R1127 VTAIL.n165 VTAIL.n164 9.3005
R1128 VTAIL.n141 VTAIL.n140 9.3005
R1129 VTAIL.n136 VTAIL.n135 9.3005
R1130 VTAIL.n147 VTAIL.n146 9.3005
R1131 VTAIL.n149 VTAIL.n148 9.3005
R1132 VTAIL.n132 VTAIL.n131 9.3005
R1133 VTAIL.n155 VTAIL.n154 9.3005
R1134 VTAIL.n157 VTAIL.n156 9.3005
R1135 VTAIL.n158 VTAIL.n127 9.3005
R1136 VTAIL.n39 VTAIL.n38 9.3005
R1137 VTAIL.n15 VTAIL.n14 9.3005
R1138 VTAIL.n10 VTAIL.n9 9.3005
R1139 VTAIL.n21 VTAIL.n20 9.3005
R1140 VTAIL.n23 VTAIL.n22 9.3005
R1141 VTAIL.n6 VTAIL.n5 9.3005
R1142 VTAIL.n29 VTAIL.n28 9.3005
R1143 VTAIL.n31 VTAIL.n30 9.3005
R1144 VTAIL.n32 VTAIL.n1 9.3005
R1145 VTAIL.n100 VTAIL.n99 9.3005
R1146 VTAIL.n95 VTAIL.n94 9.3005
R1147 VTAIL.n106 VTAIL.n105 9.3005
R1148 VTAIL.n108 VTAIL.n107 9.3005
R1149 VTAIL.n91 VTAIL.n90 9.3005
R1150 VTAIL.n114 VTAIL.n113 9.3005
R1151 VTAIL.n116 VTAIL.n115 9.3005
R1152 VTAIL.n88 VTAIL.n85 9.3005
R1153 VTAIL.n123 VTAIL.n122 9.3005
R1154 VTAIL.n58 VTAIL.n57 9.3005
R1155 VTAIL.n53 VTAIL.n52 9.3005
R1156 VTAIL.n64 VTAIL.n63 9.3005
R1157 VTAIL.n66 VTAIL.n65 9.3005
R1158 VTAIL.n49 VTAIL.n48 9.3005
R1159 VTAIL.n72 VTAIL.n71 9.3005
R1160 VTAIL.n74 VTAIL.n73 9.3005
R1161 VTAIL.n46 VTAIL.n43 9.3005
R1162 VTAIL.n81 VTAIL.n80 9.3005
R1163 VTAIL.n146 VTAIL.n145 8.92171
R1164 VTAIL.n20 VTAIL.n19 8.92171
R1165 VTAIL.n105 VTAIL.n104 8.92171
R1166 VTAIL.n63 VTAIL.n62 8.92171
R1167 VTAIL.n142 VTAIL.n136 8.14595
R1168 VTAIL.n16 VTAIL.n10 8.14595
R1169 VTAIL.n101 VTAIL.n95 8.14595
R1170 VTAIL.n59 VTAIL.n53 8.14595
R1171 VTAIL.n141 VTAIL.n138 7.3702
R1172 VTAIL.n15 VTAIL.n12 7.3702
R1173 VTAIL.n100 VTAIL.n97 7.3702
R1174 VTAIL.n58 VTAIL.n55 7.3702
R1175 VTAIL.n142 VTAIL.n141 5.81868
R1176 VTAIL.n16 VTAIL.n15 5.81868
R1177 VTAIL.n101 VTAIL.n100 5.81868
R1178 VTAIL.n59 VTAIL.n58 5.81868
R1179 VTAIL.n145 VTAIL.n136 5.04292
R1180 VTAIL.n19 VTAIL.n10 5.04292
R1181 VTAIL.n104 VTAIL.n95 5.04292
R1182 VTAIL.n62 VTAIL.n53 5.04292
R1183 VTAIL.n146 VTAIL.n134 4.26717
R1184 VTAIL.n20 VTAIL.n8 4.26717
R1185 VTAIL.n105 VTAIL.n93 4.26717
R1186 VTAIL.n63 VTAIL.n51 4.26717
R1187 VTAIL.n150 VTAIL.n149 3.49141
R1188 VTAIL.n24 VTAIL.n23 3.49141
R1189 VTAIL.n109 VTAIL.n108 3.49141
R1190 VTAIL.n67 VTAIL.n66 3.49141
R1191 VTAIL.n140 VTAIL.n139 2.84304
R1192 VTAIL.n14 VTAIL.n13 2.84304
R1193 VTAIL.n99 VTAIL.n98 2.84304
R1194 VTAIL.n57 VTAIL.n56 2.84304
R1195 VTAIL.n153 VTAIL.n132 2.71565
R1196 VTAIL.n27 VTAIL.n6 2.71565
R1197 VTAIL.n112 VTAIL.n91 2.71565
R1198 VTAIL.n70 VTAIL.n49 2.71565
R1199 VTAIL.n154 VTAIL.n130 1.93989
R1200 VTAIL.n28 VTAIL.n4 1.93989
R1201 VTAIL.n113 VTAIL.n89 1.93989
R1202 VTAIL.n71 VTAIL.n47 1.93989
R1203 VTAIL.n125 VTAIL.n83 1.5436
R1204 VTAIL.n159 VTAIL.n157 1.16414
R1205 VTAIL.n166 VTAIL.n126 1.16414
R1206 VTAIL.n33 VTAIL.n31 1.16414
R1207 VTAIL.n40 VTAIL.n0 1.16414
R1208 VTAIL.n124 VTAIL.n84 1.16414
R1209 VTAIL.n117 VTAIL.n116 1.16414
R1210 VTAIL.n82 VTAIL.n42 1.16414
R1211 VTAIL.n75 VTAIL.n74 1.16414
R1212 VTAIL VTAIL.n41 1.06516
R1213 VTAIL VTAIL.n167 0.478948
R1214 VTAIL.n158 VTAIL.n128 0.388379
R1215 VTAIL.n164 VTAIL.n163 0.388379
R1216 VTAIL.n32 VTAIL.n2 0.388379
R1217 VTAIL.n38 VTAIL.n37 0.388379
R1218 VTAIL.n122 VTAIL.n121 0.388379
R1219 VTAIL.n88 VTAIL.n86 0.388379
R1220 VTAIL.n80 VTAIL.n79 0.388379
R1221 VTAIL.n46 VTAIL.n44 0.388379
R1222 VTAIL.n140 VTAIL.n135 0.155672
R1223 VTAIL.n147 VTAIL.n135 0.155672
R1224 VTAIL.n148 VTAIL.n147 0.155672
R1225 VTAIL.n148 VTAIL.n131 0.155672
R1226 VTAIL.n155 VTAIL.n131 0.155672
R1227 VTAIL.n156 VTAIL.n155 0.155672
R1228 VTAIL.n156 VTAIL.n127 0.155672
R1229 VTAIL.n165 VTAIL.n127 0.155672
R1230 VTAIL.n14 VTAIL.n9 0.155672
R1231 VTAIL.n21 VTAIL.n9 0.155672
R1232 VTAIL.n22 VTAIL.n21 0.155672
R1233 VTAIL.n22 VTAIL.n5 0.155672
R1234 VTAIL.n29 VTAIL.n5 0.155672
R1235 VTAIL.n30 VTAIL.n29 0.155672
R1236 VTAIL.n30 VTAIL.n1 0.155672
R1237 VTAIL.n39 VTAIL.n1 0.155672
R1238 VTAIL.n123 VTAIL.n85 0.155672
R1239 VTAIL.n115 VTAIL.n85 0.155672
R1240 VTAIL.n115 VTAIL.n114 0.155672
R1241 VTAIL.n114 VTAIL.n90 0.155672
R1242 VTAIL.n107 VTAIL.n90 0.155672
R1243 VTAIL.n107 VTAIL.n106 0.155672
R1244 VTAIL.n106 VTAIL.n94 0.155672
R1245 VTAIL.n99 VTAIL.n94 0.155672
R1246 VTAIL.n81 VTAIL.n43 0.155672
R1247 VTAIL.n73 VTAIL.n43 0.155672
R1248 VTAIL.n73 VTAIL.n72 0.155672
R1249 VTAIL.n72 VTAIL.n48 0.155672
R1250 VTAIL.n65 VTAIL.n48 0.155672
R1251 VTAIL.n65 VTAIL.n64 0.155672
R1252 VTAIL.n64 VTAIL.n52 0.155672
R1253 VTAIL.n57 VTAIL.n52 0.155672
R1254 VDD2.n77 VDD2.n41 289.615
R1255 VDD2.n36 VDD2.n0 289.615
R1256 VDD2.n78 VDD2.n77 185
R1257 VDD2.n76 VDD2.n43 185
R1258 VDD2.n75 VDD2.n74 185
R1259 VDD2.n46 VDD2.n44 185
R1260 VDD2.n69 VDD2.n68 185
R1261 VDD2.n67 VDD2.n66 185
R1262 VDD2.n50 VDD2.n49 185
R1263 VDD2.n61 VDD2.n60 185
R1264 VDD2.n59 VDD2.n58 185
R1265 VDD2.n54 VDD2.n53 185
R1266 VDD2.n12 VDD2.n11 185
R1267 VDD2.n17 VDD2.n16 185
R1268 VDD2.n19 VDD2.n18 185
R1269 VDD2.n8 VDD2.n7 185
R1270 VDD2.n25 VDD2.n24 185
R1271 VDD2.n27 VDD2.n26 185
R1272 VDD2.n4 VDD2.n3 185
R1273 VDD2.n34 VDD2.n33 185
R1274 VDD2.n35 VDD2.n2 185
R1275 VDD2.n37 VDD2.n36 185
R1276 VDD2.n55 VDD2.t0 149.524
R1277 VDD2.n13 VDD2.t1 149.524
R1278 VDD2.n77 VDD2.n76 104.615
R1279 VDD2.n76 VDD2.n75 104.615
R1280 VDD2.n75 VDD2.n44 104.615
R1281 VDD2.n68 VDD2.n44 104.615
R1282 VDD2.n68 VDD2.n67 104.615
R1283 VDD2.n67 VDD2.n49 104.615
R1284 VDD2.n60 VDD2.n49 104.615
R1285 VDD2.n60 VDD2.n59 104.615
R1286 VDD2.n59 VDD2.n53 104.615
R1287 VDD2.n17 VDD2.n11 104.615
R1288 VDD2.n18 VDD2.n17 104.615
R1289 VDD2.n18 VDD2.n7 104.615
R1290 VDD2.n25 VDD2.n7 104.615
R1291 VDD2.n26 VDD2.n25 104.615
R1292 VDD2.n26 VDD2.n3 104.615
R1293 VDD2.n34 VDD2.n3 104.615
R1294 VDD2.n35 VDD2.n34 104.615
R1295 VDD2.n36 VDD2.n35 104.615
R1296 VDD2.n82 VDD2.n40 87.7946
R1297 VDD2.n82 VDD2.n81 52.9369
R1298 VDD2.t0 VDD2.n53 52.3082
R1299 VDD2.t1 VDD2.n11 52.3082
R1300 VDD2.n78 VDD2.n43 13.1884
R1301 VDD2.n37 VDD2.n2 13.1884
R1302 VDD2.n79 VDD2.n41 12.8005
R1303 VDD2.n74 VDD2.n45 12.8005
R1304 VDD2.n33 VDD2.n32 12.8005
R1305 VDD2.n38 VDD2.n0 12.8005
R1306 VDD2.n73 VDD2.n46 12.0247
R1307 VDD2.n31 VDD2.n4 12.0247
R1308 VDD2.n70 VDD2.n69 11.249
R1309 VDD2.n28 VDD2.n27 11.249
R1310 VDD2.n66 VDD2.n48 10.4732
R1311 VDD2.n24 VDD2.n6 10.4732
R1312 VDD2.n55 VDD2.n54 10.2747
R1313 VDD2.n13 VDD2.n12 10.2747
R1314 VDD2.n65 VDD2.n50 9.69747
R1315 VDD2.n23 VDD2.n8 9.69747
R1316 VDD2.n81 VDD2.n80 9.45567
R1317 VDD2.n40 VDD2.n39 9.45567
R1318 VDD2.n57 VDD2.n56 9.3005
R1319 VDD2.n52 VDD2.n51 9.3005
R1320 VDD2.n63 VDD2.n62 9.3005
R1321 VDD2.n65 VDD2.n64 9.3005
R1322 VDD2.n48 VDD2.n47 9.3005
R1323 VDD2.n71 VDD2.n70 9.3005
R1324 VDD2.n73 VDD2.n72 9.3005
R1325 VDD2.n45 VDD2.n42 9.3005
R1326 VDD2.n80 VDD2.n79 9.3005
R1327 VDD2.n39 VDD2.n38 9.3005
R1328 VDD2.n15 VDD2.n14 9.3005
R1329 VDD2.n10 VDD2.n9 9.3005
R1330 VDD2.n21 VDD2.n20 9.3005
R1331 VDD2.n23 VDD2.n22 9.3005
R1332 VDD2.n6 VDD2.n5 9.3005
R1333 VDD2.n29 VDD2.n28 9.3005
R1334 VDD2.n31 VDD2.n30 9.3005
R1335 VDD2.n32 VDD2.n1 9.3005
R1336 VDD2.n62 VDD2.n61 8.92171
R1337 VDD2.n20 VDD2.n19 8.92171
R1338 VDD2.n58 VDD2.n52 8.14595
R1339 VDD2.n16 VDD2.n10 8.14595
R1340 VDD2.n57 VDD2.n54 7.3702
R1341 VDD2.n15 VDD2.n12 7.3702
R1342 VDD2.n58 VDD2.n57 5.81868
R1343 VDD2.n16 VDD2.n15 5.81868
R1344 VDD2.n61 VDD2.n52 5.04292
R1345 VDD2.n19 VDD2.n10 5.04292
R1346 VDD2.n62 VDD2.n50 4.26717
R1347 VDD2.n20 VDD2.n8 4.26717
R1348 VDD2.n66 VDD2.n65 3.49141
R1349 VDD2.n24 VDD2.n23 3.49141
R1350 VDD2.n56 VDD2.n55 2.84304
R1351 VDD2.n14 VDD2.n13 2.84304
R1352 VDD2.n69 VDD2.n48 2.71565
R1353 VDD2.n27 VDD2.n6 2.71565
R1354 VDD2.n70 VDD2.n46 1.93989
R1355 VDD2.n28 VDD2.n4 1.93989
R1356 VDD2.n81 VDD2.n41 1.16414
R1357 VDD2.n74 VDD2.n73 1.16414
R1358 VDD2.n33 VDD2.n31 1.16414
R1359 VDD2.n40 VDD2.n0 1.16414
R1360 VDD2 VDD2.n82 0.595328
R1361 VDD2.n79 VDD2.n78 0.388379
R1362 VDD2.n45 VDD2.n43 0.388379
R1363 VDD2.n32 VDD2.n2 0.388379
R1364 VDD2.n38 VDD2.n37 0.388379
R1365 VDD2.n80 VDD2.n42 0.155672
R1366 VDD2.n72 VDD2.n42 0.155672
R1367 VDD2.n72 VDD2.n71 0.155672
R1368 VDD2.n71 VDD2.n47 0.155672
R1369 VDD2.n64 VDD2.n47 0.155672
R1370 VDD2.n64 VDD2.n63 0.155672
R1371 VDD2.n63 VDD2.n51 0.155672
R1372 VDD2.n56 VDD2.n51 0.155672
R1373 VDD2.n14 VDD2.n9 0.155672
R1374 VDD2.n21 VDD2.n9 0.155672
R1375 VDD2.n22 VDD2.n21 0.155672
R1376 VDD2.n22 VDD2.n5 0.155672
R1377 VDD2.n29 VDD2.n5 0.155672
R1378 VDD2.n30 VDD2.n29 0.155672
R1379 VDD2.n30 VDD2.n1 0.155672
R1380 VDD2.n39 VDD2.n1 0.155672
R1381 VP.n0 VP.t0 179.008
R1382 VP.n0 VP.t1 138.542
R1383 VP VP.n0 0.336784
R1384 VDD1.n36 VDD1.n0 289.615
R1385 VDD1.n77 VDD1.n41 289.615
R1386 VDD1.n37 VDD1.n36 185
R1387 VDD1.n35 VDD1.n2 185
R1388 VDD1.n34 VDD1.n33 185
R1389 VDD1.n5 VDD1.n3 185
R1390 VDD1.n28 VDD1.n27 185
R1391 VDD1.n26 VDD1.n25 185
R1392 VDD1.n9 VDD1.n8 185
R1393 VDD1.n20 VDD1.n19 185
R1394 VDD1.n18 VDD1.n17 185
R1395 VDD1.n13 VDD1.n12 185
R1396 VDD1.n53 VDD1.n52 185
R1397 VDD1.n58 VDD1.n57 185
R1398 VDD1.n60 VDD1.n59 185
R1399 VDD1.n49 VDD1.n48 185
R1400 VDD1.n66 VDD1.n65 185
R1401 VDD1.n68 VDD1.n67 185
R1402 VDD1.n45 VDD1.n44 185
R1403 VDD1.n75 VDD1.n74 185
R1404 VDD1.n76 VDD1.n43 185
R1405 VDD1.n78 VDD1.n77 185
R1406 VDD1.n14 VDD1.t1 149.524
R1407 VDD1.n54 VDD1.t0 149.524
R1408 VDD1.n36 VDD1.n35 104.615
R1409 VDD1.n35 VDD1.n34 104.615
R1410 VDD1.n34 VDD1.n3 104.615
R1411 VDD1.n27 VDD1.n3 104.615
R1412 VDD1.n27 VDD1.n26 104.615
R1413 VDD1.n26 VDD1.n8 104.615
R1414 VDD1.n19 VDD1.n8 104.615
R1415 VDD1.n19 VDD1.n18 104.615
R1416 VDD1.n18 VDD1.n12 104.615
R1417 VDD1.n58 VDD1.n52 104.615
R1418 VDD1.n59 VDD1.n58 104.615
R1419 VDD1.n59 VDD1.n48 104.615
R1420 VDD1.n66 VDD1.n48 104.615
R1421 VDD1.n67 VDD1.n66 104.615
R1422 VDD1.n67 VDD1.n44 104.615
R1423 VDD1.n75 VDD1.n44 104.615
R1424 VDD1.n76 VDD1.n75 104.615
R1425 VDD1.n77 VDD1.n76 104.615
R1426 VDD1 VDD1.n81 88.856
R1427 VDD1 VDD1.n40 53.5317
R1428 VDD1.t1 VDD1.n12 52.3082
R1429 VDD1.t0 VDD1.n52 52.3082
R1430 VDD1.n37 VDD1.n2 13.1884
R1431 VDD1.n78 VDD1.n43 13.1884
R1432 VDD1.n38 VDD1.n0 12.8005
R1433 VDD1.n33 VDD1.n4 12.8005
R1434 VDD1.n74 VDD1.n73 12.8005
R1435 VDD1.n79 VDD1.n41 12.8005
R1436 VDD1.n32 VDD1.n5 12.0247
R1437 VDD1.n72 VDD1.n45 12.0247
R1438 VDD1.n29 VDD1.n28 11.249
R1439 VDD1.n69 VDD1.n68 11.249
R1440 VDD1.n25 VDD1.n7 10.4732
R1441 VDD1.n65 VDD1.n47 10.4732
R1442 VDD1.n14 VDD1.n13 10.2747
R1443 VDD1.n54 VDD1.n53 10.2747
R1444 VDD1.n24 VDD1.n9 9.69747
R1445 VDD1.n64 VDD1.n49 9.69747
R1446 VDD1.n40 VDD1.n39 9.45567
R1447 VDD1.n81 VDD1.n80 9.45567
R1448 VDD1.n16 VDD1.n15 9.3005
R1449 VDD1.n11 VDD1.n10 9.3005
R1450 VDD1.n22 VDD1.n21 9.3005
R1451 VDD1.n24 VDD1.n23 9.3005
R1452 VDD1.n7 VDD1.n6 9.3005
R1453 VDD1.n30 VDD1.n29 9.3005
R1454 VDD1.n32 VDD1.n31 9.3005
R1455 VDD1.n4 VDD1.n1 9.3005
R1456 VDD1.n39 VDD1.n38 9.3005
R1457 VDD1.n80 VDD1.n79 9.3005
R1458 VDD1.n56 VDD1.n55 9.3005
R1459 VDD1.n51 VDD1.n50 9.3005
R1460 VDD1.n62 VDD1.n61 9.3005
R1461 VDD1.n64 VDD1.n63 9.3005
R1462 VDD1.n47 VDD1.n46 9.3005
R1463 VDD1.n70 VDD1.n69 9.3005
R1464 VDD1.n72 VDD1.n71 9.3005
R1465 VDD1.n73 VDD1.n42 9.3005
R1466 VDD1.n21 VDD1.n20 8.92171
R1467 VDD1.n61 VDD1.n60 8.92171
R1468 VDD1.n17 VDD1.n11 8.14595
R1469 VDD1.n57 VDD1.n51 8.14595
R1470 VDD1.n16 VDD1.n13 7.3702
R1471 VDD1.n56 VDD1.n53 7.3702
R1472 VDD1.n17 VDD1.n16 5.81868
R1473 VDD1.n57 VDD1.n56 5.81868
R1474 VDD1.n20 VDD1.n11 5.04292
R1475 VDD1.n60 VDD1.n51 5.04292
R1476 VDD1.n21 VDD1.n9 4.26717
R1477 VDD1.n61 VDD1.n49 4.26717
R1478 VDD1.n25 VDD1.n24 3.49141
R1479 VDD1.n65 VDD1.n64 3.49141
R1480 VDD1.n15 VDD1.n14 2.84304
R1481 VDD1.n55 VDD1.n54 2.84304
R1482 VDD1.n28 VDD1.n7 2.71565
R1483 VDD1.n68 VDD1.n47 2.71565
R1484 VDD1.n29 VDD1.n5 1.93989
R1485 VDD1.n69 VDD1.n45 1.93989
R1486 VDD1.n40 VDD1.n0 1.16414
R1487 VDD1.n33 VDD1.n32 1.16414
R1488 VDD1.n74 VDD1.n72 1.16414
R1489 VDD1.n81 VDD1.n41 1.16414
R1490 VDD1.n38 VDD1.n37 0.388379
R1491 VDD1.n4 VDD1.n2 0.388379
R1492 VDD1.n73 VDD1.n43 0.388379
R1493 VDD1.n79 VDD1.n78 0.388379
R1494 VDD1.n39 VDD1.n1 0.155672
R1495 VDD1.n31 VDD1.n1 0.155672
R1496 VDD1.n31 VDD1.n30 0.155672
R1497 VDD1.n30 VDD1.n6 0.155672
R1498 VDD1.n23 VDD1.n6 0.155672
R1499 VDD1.n23 VDD1.n22 0.155672
R1500 VDD1.n22 VDD1.n10 0.155672
R1501 VDD1.n15 VDD1.n10 0.155672
R1502 VDD1.n55 VDD1.n50 0.155672
R1503 VDD1.n62 VDD1.n50 0.155672
R1504 VDD1.n63 VDD1.n62 0.155672
R1505 VDD1.n63 VDD1.n46 0.155672
R1506 VDD1.n70 VDD1.n46 0.155672
R1507 VDD1.n71 VDD1.n70 0.155672
R1508 VDD1.n71 VDD1.n42 0.155672
R1509 VDD1.n80 VDD1.n42 0.155672
C0 VN VTAIL 1.68711f
C1 VN VDD2 1.88081f
C2 VDD2 VTAIL 3.98034f
C3 VN VP 4.51381f
C4 VP VTAIL 1.70136f
C5 VN VDD1 0.14792f
C6 VDD2 VP 0.314248f
C7 VDD1 VTAIL 3.93212f
C8 VDD1 VDD2 0.621599f
C9 VDD1 VP 2.04515f
C10 VDD2 B 3.525758f
C11 VDD1 B 5.89965f
C12 VTAIL B 5.525502f
C13 VN B 7.70254f
C14 VP B 5.583113f
C15 VDD1.n0 B 0.028316f
C16 VDD1.n1 B 0.020439f
C17 VDD1.n2 B 0.011306f
C18 VDD1.n3 B 0.02596f
C19 VDD1.n4 B 0.010983f
C20 VDD1.n5 B 0.011629f
C21 VDD1.n6 B 0.020439f
C22 VDD1.n7 B 0.010983f
C23 VDD1.n8 B 0.02596f
C24 VDD1.n9 B 0.011629f
C25 VDD1.n10 B 0.020439f
C26 VDD1.n11 B 0.010983f
C27 VDD1.n12 B 0.01947f
C28 VDD1.n13 B 0.018352f
C29 VDD1.t1 B 0.043423f
C30 VDD1.n14 B 0.116085f
C31 VDD1.n15 B 0.668348f
C32 VDD1.n16 B 0.010983f
C33 VDD1.n17 B 0.011629f
C34 VDD1.n18 B 0.02596f
C35 VDD1.n19 B 0.02596f
C36 VDD1.n20 B 0.011629f
C37 VDD1.n21 B 0.010983f
C38 VDD1.n22 B 0.020439f
C39 VDD1.n23 B 0.020439f
C40 VDD1.n24 B 0.010983f
C41 VDD1.n25 B 0.011629f
C42 VDD1.n26 B 0.02596f
C43 VDD1.n27 B 0.02596f
C44 VDD1.n28 B 0.011629f
C45 VDD1.n29 B 0.010983f
C46 VDD1.n30 B 0.020439f
C47 VDD1.n31 B 0.020439f
C48 VDD1.n32 B 0.010983f
C49 VDD1.n33 B 0.011629f
C50 VDD1.n34 B 0.02596f
C51 VDD1.n35 B 0.02596f
C52 VDD1.n36 B 0.055468f
C53 VDD1.n37 B 0.011306f
C54 VDD1.n38 B 0.010983f
C55 VDD1.n39 B 0.053108f
C56 VDD1.n40 B 0.046115f
C57 VDD1.n41 B 0.028316f
C58 VDD1.n42 B 0.020439f
C59 VDD1.n43 B 0.011306f
C60 VDD1.n44 B 0.02596f
C61 VDD1.n45 B 0.011629f
C62 VDD1.n46 B 0.020439f
C63 VDD1.n47 B 0.010983f
C64 VDD1.n48 B 0.02596f
C65 VDD1.n49 B 0.011629f
C66 VDD1.n50 B 0.020439f
C67 VDD1.n51 B 0.010983f
C68 VDD1.n52 B 0.01947f
C69 VDD1.n53 B 0.018352f
C70 VDD1.t0 B 0.043423f
C71 VDD1.n54 B 0.116085f
C72 VDD1.n55 B 0.668348f
C73 VDD1.n56 B 0.010983f
C74 VDD1.n57 B 0.011629f
C75 VDD1.n58 B 0.02596f
C76 VDD1.n59 B 0.02596f
C77 VDD1.n60 B 0.011629f
C78 VDD1.n61 B 0.010983f
C79 VDD1.n62 B 0.020439f
C80 VDD1.n63 B 0.020439f
C81 VDD1.n64 B 0.010983f
C82 VDD1.n65 B 0.011629f
C83 VDD1.n66 B 0.02596f
C84 VDD1.n67 B 0.02596f
C85 VDD1.n68 B 0.011629f
C86 VDD1.n69 B 0.010983f
C87 VDD1.n70 B 0.020439f
C88 VDD1.n71 B 0.020439f
C89 VDD1.n72 B 0.010983f
C90 VDD1.n73 B 0.010983f
C91 VDD1.n74 B 0.011629f
C92 VDD1.n75 B 0.02596f
C93 VDD1.n76 B 0.02596f
C94 VDD1.n77 B 0.055468f
C95 VDD1.n78 B 0.011306f
C96 VDD1.n79 B 0.010983f
C97 VDD1.n80 B 0.053108f
C98 VDD1.n81 B 0.482298f
C99 VP.t0 B 1.95669f
C100 VP.t1 B 1.58268f
C101 VP.n0 B 2.90294f
C102 VDD2.n0 B 0.019446f
C103 VDD2.n1 B 0.014037f
C104 VDD2.n2 B 0.007765f
C105 VDD2.n3 B 0.017828f
C106 VDD2.n4 B 0.007986f
C107 VDD2.n5 B 0.014037f
C108 VDD2.n6 B 0.007543f
C109 VDD2.n7 B 0.017828f
C110 VDD2.n8 B 0.007986f
C111 VDD2.n9 B 0.014037f
C112 VDD2.n10 B 0.007543f
C113 VDD2.n11 B 0.013371f
C114 VDD2.n12 B 0.012603f
C115 VDD2.t1 B 0.029821f
C116 VDD2.n13 B 0.079722f
C117 VDD2.n14 B 0.45899f
C118 VDD2.n15 B 0.007543f
C119 VDD2.n16 B 0.007986f
C120 VDD2.n17 B 0.017828f
C121 VDD2.n18 B 0.017828f
C122 VDD2.n19 B 0.007986f
C123 VDD2.n20 B 0.007543f
C124 VDD2.n21 B 0.014037f
C125 VDD2.n22 B 0.014037f
C126 VDD2.n23 B 0.007543f
C127 VDD2.n24 B 0.007986f
C128 VDD2.n25 B 0.017828f
C129 VDD2.n26 B 0.017828f
C130 VDD2.n27 B 0.007986f
C131 VDD2.n28 B 0.007543f
C132 VDD2.n29 B 0.014037f
C133 VDD2.n30 B 0.014037f
C134 VDD2.n31 B 0.007543f
C135 VDD2.n32 B 0.007543f
C136 VDD2.n33 B 0.007986f
C137 VDD2.n34 B 0.017828f
C138 VDD2.n35 B 0.017828f
C139 VDD2.n36 B 0.038093f
C140 VDD2.n37 B 0.007765f
C141 VDD2.n38 B 0.007543f
C142 VDD2.n39 B 0.036472f
C143 VDD2.n40 B 0.30861f
C144 VDD2.n41 B 0.019446f
C145 VDD2.n42 B 0.014037f
C146 VDD2.n43 B 0.007765f
C147 VDD2.n44 B 0.017828f
C148 VDD2.n45 B 0.007543f
C149 VDD2.n46 B 0.007986f
C150 VDD2.n47 B 0.014037f
C151 VDD2.n48 B 0.007543f
C152 VDD2.n49 B 0.017828f
C153 VDD2.n50 B 0.007986f
C154 VDD2.n51 B 0.014037f
C155 VDD2.n52 B 0.007543f
C156 VDD2.n53 B 0.013371f
C157 VDD2.n54 B 0.012603f
C158 VDD2.t0 B 0.029821f
C159 VDD2.n55 B 0.079722f
C160 VDD2.n56 B 0.45899f
C161 VDD2.n57 B 0.007543f
C162 VDD2.n58 B 0.007986f
C163 VDD2.n59 B 0.017828f
C164 VDD2.n60 B 0.017828f
C165 VDD2.n61 B 0.007986f
C166 VDD2.n62 B 0.007543f
C167 VDD2.n63 B 0.014037f
C168 VDD2.n64 B 0.014037f
C169 VDD2.n65 B 0.007543f
C170 VDD2.n66 B 0.007986f
C171 VDD2.n67 B 0.017828f
C172 VDD2.n68 B 0.017828f
C173 VDD2.n69 B 0.007986f
C174 VDD2.n70 B 0.007543f
C175 VDD2.n71 B 0.014037f
C176 VDD2.n72 B 0.014037f
C177 VDD2.n73 B 0.007543f
C178 VDD2.n74 B 0.007986f
C179 VDD2.n75 B 0.017828f
C180 VDD2.n76 B 0.017828f
C181 VDD2.n77 B 0.038093f
C182 VDD2.n78 B 0.007765f
C183 VDD2.n79 B 0.007543f
C184 VDD2.n80 B 0.036472f
C185 VDD2.n81 B 0.031045f
C186 VDD2.n82 B 1.44706f
C187 VTAIL.n0 B 0.02107f
C188 VTAIL.n1 B 0.015209f
C189 VTAIL.n2 B 0.008413f
C190 VTAIL.n3 B 0.019317f
C191 VTAIL.n4 B 0.008653f
C192 VTAIL.n5 B 0.015209f
C193 VTAIL.n6 B 0.008173f
C194 VTAIL.n7 B 0.019317f
C195 VTAIL.n8 B 0.008653f
C196 VTAIL.n9 B 0.015209f
C197 VTAIL.n10 B 0.008173f
C198 VTAIL.n11 B 0.014488f
C199 VTAIL.n12 B 0.013656f
C200 VTAIL.t1 B 0.032311f
C201 VTAIL.n13 B 0.086379f
C202 VTAIL.n14 B 0.497318f
C203 VTAIL.n15 B 0.008173f
C204 VTAIL.n16 B 0.008653f
C205 VTAIL.n17 B 0.019317f
C206 VTAIL.n18 B 0.019317f
C207 VTAIL.n19 B 0.008653f
C208 VTAIL.n20 B 0.008173f
C209 VTAIL.n21 B 0.015209f
C210 VTAIL.n22 B 0.015209f
C211 VTAIL.n23 B 0.008173f
C212 VTAIL.n24 B 0.008653f
C213 VTAIL.n25 B 0.019317f
C214 VTAIL.n26 B 0.019317f
C215 VTAIL.n27 B 0.008653f
C216 VTAIL.n28 B 0.008173f
C217 VTAIL.n29 B 0.015209f
C218 VTAIL.n30 B 0.015209f
C219 VTAIL.n31 B 0.008173f
C220 VTAIL.n32 B 0.008173f
C221 VTAIL.n33 B 0.008653f
C222 VTAIL.n34 B 0.019317f
C223 VTAIL.n35 B 0.019317f
C224 VTAIL.n36 B 0.041274f
C225 VTAIL.n37 B 0.008413f
C226 VTAIL.n38 B 0.008173f
C227 VTAIL.n39 B 0.039518f
C228 VTAIL.n40 B 0.023166f
C229 VTAIL.n41 B 0.823019f
C230 VTAIL.n42 B 0.02107f
C231 VTAIL.n43 B 0.015209f
C232 VTAIL.n44 B 0.008413f
C233 VTAIL.n45 B 0.019317f
C234 VTAIL.n46 B 0.008173f
C235 VTAIL.n47 B 0.008653f
C236 VTAIL.n48 B 0.015209f
C237 VTAIL.n49 B 0.008173f
C238 VTAIL.n50 B 0.019317f
C239 VTAIL.n51 B 0.008653f
C240 VTAIL.n52 B 0.015209f
C241 VTAIL.n53 B 0.008173f
C242 VTAIL.n54 B 0.014488f
C243 VTAIL.n55 B 0.013656f
C244 VTAIL.t3 B 0.032311f
C245 VTAIL.n56 B 0.086379f
C246 VTAIL.n57 B 0.497318f
C247 VTAIL.n58 B 0.008173f
C248 VTAIL.n59 B 0.008653f
C249 VTAIL.n60 B 0.019317f
C250 VTAIL.n61 B 0.019317f
C251 VTAIL.n62 B 0.008653f
C252 VTAIL.n63 B 0.008173f
C253 VTAIL.n64 B 0.015209f
C254 VTAIL.n65 B 0.015209f
C255 VTAIL.n66 B 0.008173f
C256 VTAIL.n67 B 0.008653f
C257 VTAIL.n68 B 0.019317f
C258 VTAIL.n69 B 0.019317f
C259 VTAIL.n70 B 0.008653f
C260 VTAIL.n71 B 0.008173f
C261 VTAIL.n72 B 0.015209f
C262 VTAIL.n73 B 0.015209f
C263 VTAIL.n74 B 0.008173f
C264 VTAIL.n75 B 0.008653f
C265 VTAIL.n76 B 0.019317f
C266 VTAIL.n77 B 0.019317f
C267 VTAIL.n78 B 0.041274f
C268 VTAIL.n79 B 0.008413f
C269 VTAIL.n80 B 0.008173f
C270 VTAIL.n81 B 0.039518f
C271 VTAIL.n82 B 0.023166f
C272 VTAIL.n83 B 0.846466f
C273 VTAIL.n84 B 0.02107f
C274 VTAIL.n85 B 0.015209f
C275 VTAIL.n86 B 0.008413f
C276 VTAIL.n87 B 0.019317f
C277 VTAIL.n88 B 0.008173f
C278 VTAIL.n89 B 0.008653f
C279 VTAIL.n90 B 0.015209f
C280 VTAIL.n91 B 0.008173f
C281 VTAIL.n92 B 0.019317f
C282 VTAIL.n93 B 0.008653f
C283 VTAIL.n94 B 0.015209f
C284 VTAIL.n95 B 0.008173f
C285 VTAIL.n96 B 0.014488f
C286 VTAIL.n97 B 0.013656f
C287 VTAIL.t0 B 0.032311f
C288 VTAIL.n98 B 0.086379f
C289 VTAIL.n99 B 0.497318f
C290 VTAIL.n100 B 0.008173f
C291 VTAIL.n101 B 0.008653f
C292 VTAIL.n102 B 0.019317f
C293 VTAIL.n103 B 0.019317f
C294 VTAIL.n104 B 0.008653f
C295 VTAIL.n105 B 0.008173f
C296 VTAIL.n106 B 0.015209f
C297 VTAIL.n107 B 0.015209f
C298 VTAIL.n108 B 0.008173f
C299 VTAIL.n109 B 0.008653f
C300 VTAIL.n110 B 0.019317f
C301 VTAIL.n111 B 0.019317f
C302 VTAIL.n112 B 0.008653f
C303 VTAIL.n113 B 0.008173f
C304 VTAIL.n114 B 0.015209f
C305 VTAIL.n115 B 0.015209f
C306 VTAIL.n116 B 0.008173f
C307 VTAIL.n117 B 0.008653f
C308 VTAIL.n118 B 0.019317f
C309 VTAIL.n119 B 0.019317f
C310 VTAIL.n120 B 0.041274f
C311 VTAIL.n121 B 0.008413f
C312 VTAIL.n122 B 0.008173f
C313 VTAIL.n123 B 0.039518f
C314 VTAIL.n124 B 0.023166f
C315 VTAIL.n125 B 0.741271f
C316 VTAIL.n126 B 0.02107f
C317 VTAIL.n127 B 0.015209f
C318 VTAIL.n128 B 0.008413f
C319 VTAIL.n129 B 0.019317f
C320 VTAIL.n130 B 0.008653f
C321 VTAIL.n131 B 0.015209f
C322 VTAIL.n132 B 0.008173f
C323 VTAIL.n133 B 0.019317f
C324 VTAIL.n134 B 0.008653f
C325 VTAIL.n135 B 0.015209f
C326 VTAIL.n136 B 0.008173f
C327 VTAIL.n137 B 0.014488f
C328 VTAIL.n138 B 0.013656f
C329 VTAIL.t2 B 0.032311f
C330 VTAIL.n139 B 0.086379f
C331 VTAIL.n140 B 0.497318f
C332 VTAIL.n141 B 0.008173f
C333 VTAIL.n142 B 0.008653f
C334 VTAIL.n143 B 0.019317f
C335 VTAIL.n144 B 0.019317f
C336 VTAIL.n145 B 0.008653f
C337 VTAIL.n146 B 0.008173f
C338 VTAIL.n147 B 0.015209f
C339 VTAIL.n148 B 0.015209f
C340 VTAIL.n149 B 0.008173f
C341 VTAIL.n150 B 0.008653f
C342 VTAIL.n151 B 0.019317f
C343 VTAIL.n152 B 0.019317f
C344 VTAIL.n153 B 0.008653f
C345 VTAIL.n154 B 0.008173f
C346 VTAIL.n155 B 0.015209f
C347 VTAIL.n156 B 0.015209f
C348 VTAIL.n157 B 0.008173f
C349 VTAIL.n158 B 0.008173f
C350 VTAIL.n159 B 0.008653f
C351 VTAIL.n160 B 0.019317f
C352 VTAIL.n161 B 0.019317f
C353 VTAIL.n162 B 0.041274f
C354 VTAIL.n163 B 0.008413f
C355 VTAIL.n164 B 0.008173f
C356 VTAIL.n165 B 0.039518f
C357 VTAIL.n166 B 0.023166f
C358 VTAIL.n167 B 0.689096f
C359 VN.t0 B 1.08976f
C360 VN.t1 B 1.34835f
.ends

