* NGSPICE file created from diff_pair_sample_1149.ext - technology: sky130A

.subckt diff_pair_sample_1149 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1768_n2138# sky130_fd_pr__pfet_01v8 ad=2.2815 pd=12.48 as=0 ps=0 w=5.85 l=1
X1 VTAIL.t7 VP.t0 VDD1.t1 w_n1768_n2138# sky130_fd_pr__pfet_01v8 ad=2.2815 pd=12.48 as=0.96525 ps=6.18 w=5.85 l=1
X2 VDD1.t2 VP.t1 VTAIL.t6 w_n1768_n2138# sky130_fd_pr__pfet_01v8 ad=0.96525 pd=6.18 as=2.2815 ps=12.48 w=5.85 l=1
X3 B.t8 B.t6 B.t7 w_n1768_n2138# sky130_fd_pr__pfet_01v8 ad=2.2815 pd=12.48 as=0 ps=0 w=5.85 l=1
X4 VDD2.t3 VN.t0 VTAIL.t1 w_n1768_n2138# sky130_fd_pr__pfet_01v8 ad=0.96525 pd=6.18 as=2.2815 ps=12.48 w=5.85 l=1
X5 VTAIL.t3 VN.t1 VDD2.t2 w_n1768_n2138# sky130_fd_pr__pfet_01v8 ad=2.2815 pd=12.48 as=0.96525 ps=6.18 w=5.85 l=1
X6 B.t5 B.t3 B.t4 w_n1768_n2138# sky130_fd_pr__pfet_01v8 ad=2.2815 pd=12.48 as=0 ps=0 w=5.85 l=1
X7 VDD2.t1 VN.t2 VTAIL.t0 w_n1768_n2138# sky130_fd_pr__pfet_01v8 ad=0.96525 pd=6.18 as=2.2815 ps=12.48 w=5.85 l=1
X8 B.t2 B.t0 B.t1 w_n1768_n2138# sky130_fd_pr__pfet_01v8 ad=2.2815 pd=12.48 as=0 ps=0 w=5.85 l=1
X9 VTAIL.t2 VN.t3 VDD2.t0 w_n1768_n2138# sky130_fd_pr__pfet_01v8 ad=2.2815 pd=12.48 as=0.96525 ps=6.18 w=5.85 l=1
X10 VTAIL.t5 VP.t2 VDD1.t0 w_n1768_n2138# sky130_fd_pr__pfet_01v8 ad=2.2815 pd=12.48 as=0.96525 ps=6.18 w=5.85 l=1
X11 VDD1.t3 VP.t3 VTAIL.t4 w_n1768_n2138# sky130_fd_pr__pfet_01v8 ad=0.96525 pd=6.18 as=2.2815 ps=12.48 w=5.85 l=1
R0 B.n286 B.n285 585
R1 B.n287 B.n44 585
R2 B.n289 B.n288 585
R3 B.n290 B.n43 585
R4 B.n292 B.n291 585
R5 B.n293 B.n42 585
R6 B.n295 B.n294 585
R7 B.n296 B.n41 585
R8 B.n298 B.n297 585
R9 B.n299 B.n40 585
R10 B.n301 B.n300 585
R11 B.n302 B.n39 585
R12 B.n304 B.n303 585
R13 B.n305 B.n38 585
R14 B.n307 B.n306 585
R15 B.n308 B.n37 585
R16 B.n310 B.n309 585
R17 B.n311 B.n36 585
R18 B.n313 B.n312 585
R19 B.n314 B.n35 585
R20 B.n316 B.n315 585
R21 B.n317 B.n34 585
R22 B.n319 B.n318 585
R23 B.n320 B.n31 585
R24 B.n323 B.n322 585
R25 B.n324 B.n30 585
R26 B.n326 B.n325 585
R27 B.n327 B.n29 585
R28 B.n329 B.n328 585
R29 B.n330 B.n28 585
R30 B.n332 B.n331 585
R31 B.n333 B.n27 585
R32 B.n335 B.n334 585
R33 B.n337 B.n336 585
R34 B.n338 B.n23 585
R35 B.n340 B.n339 585
R36 B.n341 B.n22 585
R37 B.n343 B.n342 585
R38 B.n344 B.n21 585
R39 B.n346 B.n345 585
R40 B.n347 B.n20 585
R41 B.n349 B.n348 585
R42 B.n350 B.n19 585
R43 B.n352 B.n351 585
R44 B.n353 B.n18 585
R45 B.n355 B.n354 585
R46 B.n356 B.n17 585
R47 B.n358 B.n357 585
R48 B.n359 B.n16 585
R49 B.n361 B.n360 585
R50 B.n362 B.n15 585
R51 B.n364 B.n363 585
R52 B.n365 B.n14 585
R53 B.n367 B.n366 585
R54 B.n368 B.n13 585
R55 B.n370 B.n369 585
R56 B.n371 B.n12 585
R57 B.n284 B.n45 585
R58 B.n283 B.n282 585
R59 B.n281 B.n46 585
R60 B.n280 B.n279 585
R61 B.n278 B.n47 585
R62 B.n277 B.n276 585
R63 B.n275 B.n48 585
R64 B.n274 B.n273 585
R65 B.n272 B.n49 585
R66 B.n271 B.n270 585
R67 B.n269 B.n50 585
R68 B.n268 B.n267 585
R69 B.n266 B.n51 585
R70 B.n265 B.n264 585
R71 B.n263 B.n52 585
R72 B.n262 B.n261 585
R73 B.n260 B.n53 585
R74 B.n259 B.n258 585
R75 B.n257 B.n54 585
R76 B.n256 B.n255 585
R77 B.n254 B.n55 585
R78 B.n253 B.n252 585
R79 B.n251 B.n56 585
R80 B.n250 B.n249 585
R81 B.n248 B.n57 585
R82 B.n247 B.n246 585
R83 B.n245 B.n58 585
R84 B.n244 B.n243 585
R85 B.n242 B.n59 585
R86 B.n241 B.n240 585
R87 B.n239 B.n60 585
R88 B.n238 B.n237 585
R89 B.n236 B.n61 585
R90 B.n235 B.n234 585
R91 B.n233 B.n62 585
R92 B.n232 B.n231 585
R93 B.n230 B.n63 585
R94 B.n229 B.n228 585
R95 B.n227 B.n64 585
R96 B.n226 B.n225 585
R97 B.n224 B.n65 585
R98 B.n137 B.n98 585
R99 B.n139 B.n138 585
R100 B.n140 B.n97 585
R101 B.n142 B.n141 585
R102 B.n143 B.n96 585
R103 B.n145 B.n144 585
R104 B.n146 B.n95 585
R105 B.n148 B.n147 585
R106 B.n149 B.n94 585
R107 B.n151 B.n150 585
R108 B.n152 B.n93 585
R109 B.n154 B.n153 585
R110 B.n155 B.n92 585
R111 B.n157 B.n156 585
R112 B.n158 B.n91 585
R113 B.n160 B.n159 585
R114 B.n161 B.n90 585
R115 B.n163 B.n162 585
R116 B.n164 B.n89 585
R117 B.n166 B.n165 585
R118 B.n167 B.n88 585
R119 B.n169 B.n168 585
R120 B.n170 B.n87 585
R121 B.n172 B.n171 585
R122 B.n174 B.n173 585
R123 B.n175 B.n83 585
R124 B.n177 B.n176 585
R125 B.n178 B.n82 585
R126 B.n180 B.n179 585
R127 B.n181 B.n81 585
R128 B.n183 B.n182 585
R129 B.n184 B.n80 585
R130 B.n186 B.n185 585
R131 B.n188 B.n77 585
R132 B.n190 B.n189 585
R133 B.n191 B.n76 585
R134 B.n193 B.n192 585
R135 B.n194 B.n75 585
R136 B.n196 B.n195 585
R137 B.n197 B.n74 585
R138 B.n199 B.n198 585
R139 B.n200 B.n73 585
R140 B.n202 B.n201 585
R141 B.n203 B.n72 585
R142 B.n205 B.n204 585
R143 B.n206 B.n71 585
R144 B.n208 B.n207 585
R145 B.n209 B.n70 585
R146 B.n211 B.n210 585
R147 B.n212 B.n69 585
R148 B.n214 B.n213 585
R149 B.n215 B.n68 585
R150 B.n217 B.n216 585
R151 B.n218 B.n67 585
R152 B.n220 B.n219 585
R153 B.n221 B.n66 585
R154 B.n223 B.n222 585
R155 B.n136 B.n135 585
R156 B.n134 B.n99 585
R157 B.n133 B.n132 585
R158 B.n131 B.n100 585
R159 B.n130 B.n129 585
R160 B.n128 B.n101 585
R161 B.n127 B.n126 585
R162 B.n125 B.n102 585
R163 B.n124 B.n123 585
R164 B.n122 B.n103 585
R165 B.n121 B.n120 585
R166 B.n119 B.n104 585
R167 B.n118 B.n117 585
R168 B.n116 B.n105 585
R169 B.n115 B.n114 585
R170 B.n113 B.n106 585
R171 B.n112 B.n111 585
R172 B.n110 B.n107 585
R173 B.n109 B.n108 585
R174 B.n2 B.n0 585
R175 B.n401 B.n1 585
R176 B.n400 B.n399 585
R177 B.n398 B.n3 585
R178 B.n397 B.n396 585
R179 B.n395 B.n4 585
R180 B.n394 B.n393 585
R181 B.n392 B.n5 585
R182 B.n391 B.n390 585
R183 B.n389 B.n6 585
R184 B.n388 B.n387 585
R185 B.n386 B.n7 585
R186 B.n385 B.n384 585
R187 B.n383 B.n8 585
R188 B.n382 B.n381 585
R189 B.n380 B.n9 585
R190 B.n379 B.n378 585
R191 B.n377 B.n10 585
R192 B.n376 B.n375 585
R193 B.n374 B.n11 585
R194 B.n373 B.n372 585
R195 B.n403 B.n402 585
R196 B.n137 B.n136 444.452
R197 B.n372 B.n371 444.452
R198 B.n222 B.n65 444.452
R199 B.n286 B.n45 444.452
R200 B.n78 B.t3 343.911
R201 B.n84 B.t9 343.911
R202 B.n24 B.t6 343.911
R203 B.n32 B.t0 343.911
R204 B.n78 B.t5 291.077
R205 B.n32 B.t1 291.077
R206 B.n84 B.t11 291.077
R207 B.n24 B.t7 291.077
R208 B.n79 B.t4 265.284
R209 B.n33 B.t2 265.284
R210 B.n85 B.t10 265.284
R211 B.n25 B.t8 265.284
R212 B.n136 B.n99 163.367
R213 B.n132 B.n99 163.367
R214 B.n132 B.n131 163.367
R215 B.n131 B.n130 163.367
R216 B.n130 B.n101 163.367
R217 B.n126 B.n101 163.367
R218 B.n126 B.n125 163.367
R219 B.n125 B.n124 163.367
R220 B.n124 B.n103 163.367
R221 B.n120 B.n103 163.367
R222 B.n120 B.n119 163.367
R223 B.n119 B.n118 163.367
R224 B.n118 B.n105 163.367
R225 B.n114 B.n105 163.367
R226 B.n114 B.n113 163.367
R227 B.n113 B.n112 163.367
R228 B.n112 B.n107 163.367
R229 B.n108 B.n107 163.367
R230 B.n108 B.n2 163.367
R231 B.n402 B.n2 163.367
R232 B.n402 B.n401 163.367
R233 B.n401 B.n400 163.367
R234 B.n400 B.n3 163.367
R235 B.n396 B.n3 163.367
R236 B.n396 B.n395 163.367
R237 B.n395 B.n394 163.367
R238 B.n394 B.n5 163.367
R239 B.n390 B.n5 163.367
R240 B.n390 B.n389 163.367
R241 B.n389 B.n388 163.367
R242 B.n388 B.n7 163.367
R243 B.n384 B.n7 163.367
R244 B.n384 B.n383 163.367
R245 B.n383 B.n382 163.367
R246 B.n382 B.n9 163.367
R247 B.n378 B.n9 163.367
R248 B.n378 B.n377 163.367
R249 B.n377 B.n376 163.367
R250 B.n376 B.n11 163.367
R251 B.n372 B.n11 163.367
R252 B.n138 B.n137 163.367
R253 B.n138 B.n97 163.367
R254 B.n142 B.n97 163.367
R255 B.n143 B.n142 163.367
R256 B.n144 B.n143 163.367
R257 B.n144 B.n95 163.367
R258 B.n148 B.n95 163.367
R259 B.n149 B.n148 163.367
R260 B.n150 B.n149 163.367
R261 B.n150 B.n93 163.367
R262 B.n154 B.n93 163.367
R263 B.n155 B.n154 163.367
R264 B.n156 B.n155 163.367
R265 B.n156 B.n91 163.367
R266 B.n160 B.n91 163.367
R267 B.n161 B.n160 163.367
R268 B.n162 B.n161 163.367
R269 B.n162 B.n89 163.367
R270 B.n166 B.n89 163.367
R271 B.n167 B.n166 163.367
R272 B.n168 B.n167 163.367
R273 B.n168 B.n87 163.367
R274 B.n172 B.n87 163.367
R275 B.n173 B.n172 163.367
R276 B.n173 B.n83 163.367
R277 B.n177 B.n83 163.367
R278 B.n178 B.n177 163.367
R279 B.n179 B.n178 163.367
R280 B.n179 B.n81 163.367
R281 B.n183 B.n81 163.367
R282 B.n184 B.n183 163.367
R283 B.n185 B.n184 163.367
R284 B.n185 B.n77 163.367
R285 B.n190 B.n77 163.367
R286 B.n191 B.n190 163.367
R287 B.n192 B.n191 163.367
R288 B.n192 B.n75 163.367
R289 B.n196 B.n75 163.367
R290 B.n197 B.n196 163.367
R291 B.n198 B.n197 163.367
R292 B.n198 B.n73 163.367
R293 B.n202 B.n73 163.367
R294 B.n203 B.n202 163.367
R295 B.n204 B.n203 163.367
R296 B.n204 B.n71 163.367
R297 B.n208 B.n71 163.367
R298 B.n209 B.n208 163.367
R299 B.n210 B.n209 163.367
R300 B.n210 B.n69 163.367
R301 B.n214 B.n69 163.367
R302 B.n215 B.n214 163.367
R303 B.n216 B.n215 163.367
R304 B.n216 B.n67 163.367
R305 B.n220 B.n67 163.367
R306 B.n221 B.n220 163.367
R307 B.n222 B.n221 163.367
R308 B.n226 B.n65 163.367
R309 B.n227 B.n226 163.367
R310 B.n228 B.n227 163.367
R311 B.n228 B.n63 163.367
R312 B.n232 B.n63 163.367
R313 B.n233 B.n232 163.367
R314 B.n234 B.n233 163.367
R315 B.n234 B.n61 163.367
R316 B.n238 B.n61 163.367
R317 B.n239 B.n238 163.367
R318 B.n240 B.n239 163.367
R319 B.n240 B.n59 163.367
R320 B.n244 B.n59 163.367
R321 B.n245 B.n244 163.367
R322 B.n246 B.n245 163.367
R323 B.n246 B.n57 163.367
R324 B.n250 B.n57 163.367
R325 B.n251 B.n250 163.367
R326 B.n252 B.n251 163.367
R327 B.n252 B.n55 163.367
R328 B.n256 B.n55 163.367
R329 B.n257 B.n256 163.367
R330 B.n258 B.n257 163.367
R331 B.n258 B.n53 163.367
R332 B.n262 B.n53 163.367
R333 B.n263 B.n262 163.367
R334 B.n264 B.n263 163.367
R335 B.n264 B.n51 163.367
R336 B.n268 B.n51 163.367
R337 B.n269 B.n268 163.367
R338 B.n270 B.n269 163.367
R339 B.n270 B.n49 163.367
R340 B.n274 B.n49 163.367
R341 B.n275 B.n274 163.367
R342 B.n276 B.n275 163.367
R343 B.n276 B.n47 163.367
R344 B.n280 B.n47 163.367
R345 B.n281 B.n280 163.367
R346 B.n282 B.n281 163.367
R347 B.n282 B.n45 163.367
R348 B.n371 B.n370 163.367
R349 B.n370 B.n13 163.367
R350 B.n366 B.n13 163.367
R351 B.n366 B.n365 163.367
R352 B.n365 B.n364 163.367
R353 B.n364 B.n15 163.367
R354 B.n360 B.n15 163.367
R355 B.n360 B.n359 163.367
R356 B.n359 B.n358 163.367
R357 B.n358 B.n17 163.367
R358 B.n354 B.n17 163.367
R359 B.n354 B.n353 163.367
R360 B.n353 B.n352 163.367
R361 B.n352 B.n19 163.367
R362 B.n348 B.n19 163.367
R363 B.n348 B.n347 163.367
R364 B.n347 B.n346 163.367
R365 B.n346 B.n21 163.367
R366 B.n342 B.n21 163.367
R367 B.n342 B.n341 163.367
R368 B.n341 B.n340 163.367
R369 B.n340 B.n23 163.367
R370 B.n336 B.n23 163.367
R371 B.n336 B.n335 163.367
R372 B.n335 B.n27 163.367
R373 B.n331 B.n27 163.367
R374 B.n331 B.n330 163.367
R375 B.n330 B.n329 163.367
R376 B.n329 B.n29 163.367
R377 B.n325 B.n29 163.367
R378 B.n325 B.n324 163.367
R379 B.n324 B.n323 163.367
R380 B.n323 B.n31 163.367
R381 B.n318 B.n31 163.367
R382 B.n318 B.n317 163.367
R383 B.n317 B.n316 163.367
R384 B.n316 B.n35 163.367
R385 B.n312 B.n35 163.367
R386 B.n312 B.n311 163.367
R387 B.n311 B.n310 163.367
R388 B.n310 B.n37 163.367
R389 B.n306 B.n37 163.367
R390 B.n306 B.n305 163.367
R391 B.n305 B.n304 163.367
R392 B.n304 B.n39 163.367
R393 B.n300 B.n39 163.367
R394 B.n300 B.n299 163.367
R395 B.n299 B.n298 163.367
R396 B.n298 B.n41 163.367
R397 B.n294 B.n41 163.367
R398 B.n294 B.n293 163.367
R399 B.n293 B.n292 163.367
R400 B.n292 B.n43 163.367
R401 B.n288 B.n43 163.367
R402 B.n288 B.n287 163.367
R403 B.n287 B.n286 163.367
R404 B.n187 B.n79 59.5399
R405 B.n86 B.n85 59.5399
R406 B.n26 B.n25 59.5399
R407 B.n321 B.n33 59.5399
R408 B.n373 B.n12 28.8785
R409 B.n285 B.n284 28.8785
R410 B.n224 B.n223 28.8785
R411 B.n135 B.n98 28.8785
R412 B.n79 B.n78 25.7944
R413 B.n85 B.n84 25.7944
R414 B.n25 B.n24 25.7944
R415 B.n33 B.n32 25.7944
R416 B B.n403 18.0485
R417 B.n369 B.n12 10.6151
R418 B.n369 B.n368 10.6151
R419 B.n368 B.n367 10.6151
R420 B.n367 B.n14 10.6151
R421 B.n363 B.n14 10.6151
R422 B.n363 B.n362 10.6151
R423 B.n362 B.n361 10.6151
R424 B.n361 B.n16 10.6151
R425 B.n357 B.n16 10.6151
R426 B.n357 B.n356 10.6151
R427 B.n356 B.n355 10.6151
R428 B.n355 B.n18 10.6151
R429 B.n351 B.n18 10.6151
R430 B.n351 B.n350 10.6151
R431 B.n350 B.n349 10.6151
R432 B.n349 B.n20 10.6151
R433 B.n345 B.n20 10.6151
R434 B.n345 B.n344 10.6151
R435 B.n344 B.n343 10.6151
R436 B.n343 B.n22 10.6151
R437 B.n339 B.n22 10.6151
R438 B.n339 B.n338 10.6151
R439 B.n338 B.n337 10.6151
R440 B.n334 B.n333 10.6151
R441 B.n333 B.n332 10.6151
R442 B.n332 B.n28 10.6151
R443 B.n328 B.n28 10.6151
R444 B.n328 B.n327 10.6151
R445 B.n327 B.n326 10.6151
R446 B.n326 B.n30 10.6151
R447 B.n322 B.n30 10.6151
R448 B.n320 B.n319 10.6151
R449 B.n319 B.n34 10.6151
R450 B.n315 B.n34 10.6151
R451 B.n315 B.n314 10.6151
R452 B.n314 B.n313 10.6151
R453 B.n313 B.n36 10.6151
R454 B.n309 B.n36 10.6151
R455 B.n309 B.n308 10.6151
R456 B.n308 B.n307 10.6151
R457 B.n307 B.n38 10.6151
R458 B.n303 B.n38 10.6151
R459 B.n303 B.n302 10.6151
R460 B.n302 B.n301 10.6151
R461 B.n301 B.n40 10.6151
R462 B.n297 B.n40 10.6151
R463 B.n297 B.n296 10.6151
R464 B.n296 B.n295 10.6151
R465 B.n295 B.n42 10.6151
R466 B.n291 B.n42 10.6151
R467 B.n291 B.n290 10.6151
R468 B.n290 B.n289 10.6151
R469 B.n289 B.n44 10.6151
R470 B.n285 B.n44 10.6151
R471 B.n225 B.n224 10.6151
R472 B.n225 B.n64 10.6151
R473 B.n229 B.n64 10.6151
R474 B.n230 B.n229 10.6151
R475 B.n231 B.n230 10.6151
R476 B.n231 B.n62 10.6151
R477 B.n235 B.n62 10.6151
R478 B.n236 B.n235 10.6151
R479 B.n237 B.n236 10.6151
R480 B.n237 B.n60 10.6151
R481 B.n241 B.n60 10.6151
R482 B.n242 B.n241 10.6151
R483 B.n243 B.n242 10.6151
R484 B.n243 B.n58 10.6151
R485 B.n247 B.n58 10.6151
R486 B.n248 B.n247 10.6151
R487 B.n249 B.n248 10.6151
R488 B.n249 B.n56 10.6151
R489 B.n253 B.n56 10.6151
R490 B.n254 B.n253 10.6151
R491 B.n255 B.n254 10.6151
R492 B.n255 B.n54 10.6151
R493 B.n259 B.n54 10.6151
R494 B.n260 B.n259 10.6151
R495 B.n261 B.n260 10.6151
R496 B.n261 B.n52 10.6151
R497 B.n265 B.n52 10.6151
R498 B.n266 B.n265 10.6151
R499 B.n267 B.n266 10.6151
R500 B.n267 B.n50 10.6151
R501 B.n271 B.n50 10.6151
R502 B.n272 B.n271 10.6151
R503 B.n273 B.n272 10.6151
R504 B.n273 B.n48 10.6151
R505 B.n277 B.n48 10.6151
R506 B.n278 B.n277 10.6151
R507 B.n279 B.n278 10.6151
R508 B.n279 B.n46 10.6151
R509 B.n283 B.n46 10.6151
R510 B.n284 B.n283 10.6151
R511 B.n139 B.n98 10.6151
R512 B.n140 B.n139 10.6151
R513 B.n141 B.n140 10.6151
R514 B.n141 B.n96 10.6151
R515 B.n145 B.n96 10.6151
R516 B.n146 B.n145 10.6151
R517 B.n147 B.n146 10.6151
R518 B.n147 B.n94 10.6151
R519 B.n151 B.n94 10.6151
R520 B.n152 B.n151 10.6151
R521 B.n153 B.n152 10.6151
R522 B.n153 B.n92 10.6151
R523 B.n157 B.n92 10.6151
R524 B.n158 B.n157 10.6151
R525 B.n159 B.n158 10.6151
R526 B.n159 B.n90 10.6151
R527 B.n163 B.n90 10.6151
R528 B.n164 B.n163 10.6151
R529 B.n165 B.n164 10.6151
R530 B.n165 B.n88 10.6151
R531 B.n169 B.n88 10.6151
R532 B.n170 B.n169 10.6151
R533 B.n171 B.n170 10.6151
R534 B.n175 B.n174 10.6151
R535 B.n176 B.n175 10.6151
R536 B.n176 B.n82 10.6151
R537 B.n180 B.n82 10.6151
R538 B.n181 B.n180 10.6151
R539 B.n182 B.n181 10.6151
R540 B.n182 B.n80 10.6151
R541 B.n186 B.n80 10.6151
R542 B.n189 B.n188 10.6151
R543 B.n189 B.n76 10.6151
R544 B.n193 B.n76 10.6151
R545 B.n194 B.n193 10.6151
R546 B.n195 B.n194 10.6151
R547 B.n195 B.n74 10.6151
R548 B.n199 B.n74 10.6151
R549 B.n200 B.n199 10.6151
R550 B.n201 B.n200 10.6151
R551 B.n201 B.n72 10.6151
R552 B.n205 B.n72 10.6151
R553 B.n206 B.n205 10.6151
R554 B.n207 B.n206 10.6151
R555 B.n207 B.n70 10.6151
R556 B.n211 B.n70 10.6151
R557 B.n212 B.n211 10.6151
R558 B.n213 B.n212 10.6151
R559 B.n213 B.n68 10.6151
R560 B.n217 B.n68 10.6151
R561 B.n218 B.n217 10.6151
R562 B.n219 B.n218 10.6151
R563 B.n219 B.n66 10.6151
R564 B.n223 B.n66 10.6151
R565 B.n135 B.n134 10.6151
R566 B.n134 B.n133 10.6151
R567 B.n133 B.n100 10.6151
R568 B.n129 B.n100 10.6151
R569 B.n129 B.n128 10.6151
R570 B.n128 B.n127 10.6151
R571 B.n127 B.n102 10.6151
R572 B.n123 B.n102 10.6151
R573 B.n123 B.n122 10.6151
R574 B.n122 B.n121 10.6151
R575 B.n121 B.n104 10.6151
R576 B.n117 B.n104 10.6151
R577 B.n117 B.n116 10.6151
R578 B.n116 B.n115 10.6151
R579 B.n115 B.n106 10.6151
R580 B.n111 B.n106 10.6151
R581 B.n111 B.n110 10.6151
R582 B.n110 B.n109 10.6151
R583 B.n109 B.n0 10.6151
R584 B.n399 B.n1 10.6151
R585 B.n399 B.n398 10.6151
R586 B.n398 B.n397 10.6151
R587 B.n397 B.n4 10.6151
R588 B.n393 B.n4 10.6151
R589 B.n393 B.n392 10.6151
R590 B.n392 B.n391 10.6151
R591 B.n391 B.n6 10.6151
R592 B.n387 B.n6 10.6151
R593 B.n387 B.n386 10.6151
R594 B.n386 B.n385 10.6151
R595 B.n385 B.n8 10.6151
R596 B.n381 B.n8 10.6151
R597 B.n381 B.n380 10.6151
R598 B.n380 B.n379 10.6151
R599 B.n379 B.n10 10.6151
R600 B.n375 B.n10 10.6151
R601 B.n375 B.n374 10.6151
R602 B.n374 B.n373 10.6151
R603 B.n334 B.n26 6.5566
R604 B.n322 B.n321 6.5566
R605 B.n174 B.n86 6.5566
R606 B.n187 B.n186 6.5566
R607 B.n337 B.n26 4.05904
R608 B.n321 B.n320 4.05904
R609 B.n171 B.n86 4.05904
R610 B.n188 B.n187 4.05904
R611 B.n403 B.n0 2.81026
R612 B.n403 B.n1 2.81026
R613 VP.n0 VP.t2 199.117
R614 VP.n0 VP.t3 199.03
R615 VP.n2 VP.t0 180.51
R616 VP.n3 VP.t1 180.51
R617 VP.n4 VP.n3 80.6037
R618 VP.n2 VP.n1 80.6037
R619 VP.n1 VP.n0 68.0032
R620 VP.n3 VP.n2 48.2005
R621 VP.n4 VP.n1 0.380177
R622 VP VP.n4 0.146778
R623 VDD1 VDD1.n1 128.417
R624 VDD1 VDD1.n0 95.7518
R625 VDD1.n0 VDD1.t0 5.55691
R626 VDD1.n0 VDD1.t3 5.55691
R627 VDD1.n1 VDD1.t1 5.55691
R628 VDD1.n1 VDD1.t2 5.55691
R629 VTAIL.n238 VTAIL.n237 756.745
R630 VTAIL.n28 VTAIL.n27 756.745
R631 VTAIL.n58 VTAIL.n57 756.745
R632 VTAIL.n88 VTAIL.n87 756.745
R633 VTAIL.n208 VTAIL.n207 756.745
R634 VTAIL.n178 VTAIL.n177 756.745
R635 VTAIL.n148 VTAIL.n147 756.745
R636 VTAIL.n118 VTAIL.n117 756.745
R637 VTAIL.n221 VTAIL.n220 585
R638 VTAIL.n223 VTAIL.n222 585
R639 VTAIL.n216 VTAIL.n215 585
R640 VTAIL.n229 VTAIL.n228 585
R641 VTAIL.n231 VTAIL.n230 585
R642 VTAIL.n212 VTAIL.n211 585
R643 VTAIL.n237 VTAIL.n236 585
R644 VTAIL.n11 VTAIL.n10 585
R645 VTAIL.n13 VTAIL.n12 585
R646 VTAIL.n6 VTAIL.n5 585
R647 VTAIL.n19 VTAIL.n18 585
R648 VTAIL.n21 VTAIL.n20 585
R649 VTAIL.n2 VTAIL.n1 585
R650 VTAIL.n27 VTAIL.n26 585
R651 VTAIL.n41 VTAIL.n40 585
R652 VTAIL.n43 VTAIL.n42 585
R653 VTAIL.n36 VTAIL.n35 585
R654 VTAIL.n49 VTAIL.n48 585
R655 VTAIL.n51 VTAIL.n50 585
R656 VTAIL.n32 VTAIL.n31 585
R657 VTAIL.n57 VTAIL.n56 585
R658 VTAIL.n71 VTAIL.n70 585
R659 VTAIL.n73 VTAIL.n72 585
R660 VTAIL.n66 VTAIL.n65 585
R661 VTAIL.n79 VTAIL.n78 585
R662 VTAIL.n81 VTAIL.n80 585
R663 VTAIL.n62 VTAIL.n61 585
R664 VTAIL.n87 VTAIL.n86 585
R665 VTAIL.n207 VTAIL.n206 585
R666 VTAIL.n182 VTAIL.n181 585
R667 VTAIL.n201 VTAIL.n200 585
R668 VTAIL.n199 VTAIL.n198 585
R669 VTAIL.n186 VTAIL.n185 585
R670 VTAIL.n193 VTAIL.n192 585
R671 VTAIL.n191 VTAIL.n190 585
R672 VTAIL.n177 VTAIL.n176 585
R673 VTAIL.n152 VTAIL.n151 585
R674 VTAIL.n171 VTAIL.n170 585
R675 VTAIL.n169 VTAIL.n168 585
R676 VTAIL.n156 VTAIL.n155 585
R677 VTAIL.n163 VTAIL.n162 585
R678 VTAIL.n161 VTAIL.n160 585
R679 VTAIL.n147 VTAIL.n146 585
R680 VTAIL.n122 VTAIL.n121 585
R681 VTAIL.n141 VTAIL.n140 585
R682 VTAIL.n139 VTAIL.n138 585
R683 VTAIL.n126 VTAIL.n125 585
R684 VTAIL.n133 VTAIL.n132 585
R685 VTAIL.n131 VTAIL.n130 585
R686 VTAIL.n117 VTAIL.n116 585
R687 VTAIL.n92 VTAIL.n91 585
R688 VTAIL.n111 VTAIL.n110 585
R689 VTAIL.n109 VTAIL.n108 585
R690 VTAIL.n96 VTAIL.n95 585
R691 VTAIL.n103 VTAIL.n102 585
R692 VTAIL.n101 VTAIL.n100 585
R693 VTAIL.n219 VTAIL.t1 329.175
R694 VTAIL.n9 VTAIL.t3 329.175
R695 VTAIL.n39 VTAIL.t6 329.175
R696 VTAIL.n69 VTAIL.t7 329.175
R697 VTAIL.n189 VTAIL.t4 329.175
R698 VTAIL.n159 VTAIL.t5 329.175
R699 VTAIL.n129 VTAIL.t0 329.175
R700 VTAIL.n99 VTAIL.t2 329.175
R701 VTAIL.n222 VTAIL.n221 171.744
R702 VTAIL.n222 VTAIL.n215 171.744
R703 VTAIL.n229 VTAIL.n215 171.744
R704 VTAIL.n230 VTAIL.n229 171.744
R705 VTAIL.n230 VTAIL.n211 171.744
R706 VTAIL.n237 VTAIL.n211 171.744
R707 VTAIL.n12 VTAIL.n11 171.744
R708 VTAIL.n12 VTAIL.n5 171.744
R709 VTAIL.n19 VTAIL.n5 171.744
R710 VTAIL.n20 VTAIL.n19 171.744
R711 VTAIL.n20 VTAIL.n1 171.744
R712 VTAIL.n27 VTAIL.n1 171.744
R713 VTAIL.n42 VTAIL.n41 171.744
R714 VTAIL.n42 VTAIL.n35 171.744
R715 VTAIL.n49 VTAIL.n35 171.744
R716 VTAIL.n50 VTAIL.n49 171.744
R717 VTAIL.n50 VTAIL.n31 171.744
R718 VTAIL.n57 VTAIL.n31 171.744
R719 VTAIL.n72 VTAIL.n71 171.744
R720 VTAIL.n72 VTAIL.n65 171.744
R721 VTAIL.n79 VTAIL.n65 171.744
R722 VTAIL.n80 VTAIL.n79 171.744
R723 VTAIL.n80 VTAIL.n61 171.744
R724 VTAIL.n87 VTAIL.n61 171.744
R725 VTAIL.n207 VTAIL.n181 171.744
R726 VTAIL.n200 VTAIL.n181 171.744
R727 VTAIL.n200 VTAIL.n199 171.744
R728 VTAIL.n199 VTAIL.n185 171.744
R729 VTAIL.n192 VTAIL.n185 171.744
R730 VTAIL.n192 VTAIL.n191 171.744
R731 VTAIL.n177 VTAIL.n151 171.744
R732 VTAIL.n170 VTAIL.n151 171.744
R733 VTAIL.n170 VTAIL.n169 171.744
R734 VTAIL.n169 VTAIL.n155 171.744
R735 VTAIL.n162 VTAIL.n155 171.744
R736 VTAIL.n162 VTAIL.n161 171.744
R737 VTAIL.n147 VTAIL.n121 171.744
R738 VTAIL.n140 VTAIL.n121 171.744
R739 VTAIL.n140 VTAIL.n139 171.744
R740 VTAIL.n139 VTAIL.n125 171.744
R741 VTAIL.n132 VTAIL.n125 171.744
R742 VTAIL.n132 VTAIL.n131 171.744
R743 VTAIL.n117 VTAIL.n91 171.744
R744 VTAIL.n110 VTAIL.n91 171.744
R745 VTAIL.n110 VTAIL.n109 171.744
R746 VTAIL.n109 VTAIL.n95 171.744
R747 VTAIL.n102 VTAIL.n95 171.744
R748 VTAIL.n102 VTAIL.n101 171.744
R749 VTAIL.n221 VTAIL.t1 85.8723
R750 VTAIL.n11 VTAIL.t3 85.8723
R751 VTAIL.n41 VTAIL.t6 85.8723
R752 VTAIL.n71 VTAIL.t7 85.8723
R753 VTAIL.n191 VTAIL.t4 85.8723
R754 VTAIL.n161 VTAIL.t5 85.8723
R755 VTAIL.n131 VTAIL.t0 85.8723
R756 VTAIL.n101 VTAIL.t2 85.8723
R757 VTAIL.n239 VTAIL.n238 35.0944
R758 VTAIL.n29 VTAIL.n28 35.0944
R759 VTAIL.n59 VTAIL.n58 35.0944
R760 VTAIL.n89 VTAIL.n88 35.0944
R761 VTAIL.n209 VTAIL.n208 35.0944
R762 VTAIL.n179 VTAIL.n178 35.0944
R763 VTAIL.n149 VTAIL.n148 35.0944
R764 VTAIL.n119 VTAIL.n118 35.0944
R765 VTAIL.n239 VTAIL.n209 18.5565
R766 VTAIL.n119 VTAIL.n89 18.5565
R767 VTAIL.n236 VTAIL.n210 12.0247
R768 VTAIL.n26 VTAIL.n0 12.0247
R769 VTAIL.n56 VTAIL.n30 12.0247
R770 VTAIL.n86 VTAIL.n60 12.0247
R771 VTAIL.n206 VTAIL.n180 12.0247
R772 VTAIL.n176 VTAIL.n150 12.0247
R773 VTAIL.n146 VTAIL.n120 12.0247
R774 VTAIL.n116 VTAIL.n90 12.0247
R775 VTAIL.n235 VTAIL.n212 11.249
R776 VTAIL.n25 VTAIL.n2 11.249
R777 VTAIL.n55 VTAIL.n32 11.249
R778 VTAIL.n85 VTAIL.n62 11.249
R779 VTAIL.n205 VTAIL.n182 11.249
R780 VTAIL.n175 VTAIL.n152 11.249
R781 VTAIL.n145 VTAIL.n122 11.249
R782 VTAIL.n115 VTAIL.n92 11.249
R783 VTAIL.n220 VTAIL.n219 10.722
R784 VTAIL.n10 VTAIL.n9 10.722
R785 VTAIL.n40 VTAIL.n39 10.722
R786 VTAIL.n70 VTAIL.n69 10.722
R787 VTAIL.n190 VTAIL.n189 10.722
R788 VTAIL.n160 VTAIL.n159 10.722
R789 VTAIL.n130 VTAIL.n129 10.722
R790 VTAIL.n100 VTAIL.n99 10.722
R791 VTAIL.n232 VTAIL.n231 10.4732
R792 VTAIL.n22 VTAIL.n21 10.4732
R793 VTAIL.n52 VTAIL.n51 10.4732
R794 VTAIL.n82 VTAIL.n81 10.4732
R795 VTAIL.n202 VTAIL.n201 10.4732
R796 VTAIL.n172 VTAIL.n171 10.4732
R797 VTAIL.n142 VTAIL.n141 10.4732
R798 VTAIL.n112 VTAIL.n111 10.4732
R799 VTAIL.n228 VTAIL.n214 9.69747
R800 VTAIL.n18 VTAIL.n4 9.69747
R801 VTAIL.n48 VTAIL.n34 9.69747
R802 VTAIL.n78 VTAIL.n64 9.69747
R803 VTAIL.n198 VTAIL.n184 9.69747
R804 VTAIL.n168 VTAIL.n154 9.69747
R805 VTAIL.n138 VTAIL.n124 9.69747
R806 VTAIL.n108 VTAIL.n94 9.69747
R807 VTAIL.n234 VTAIL.n210 9.45567
R808 VTAIL.n24 VTAIL.n0 9.45567
R809 VTAIL.n54 VTAIL.n30 9.45567
R810 VTAIL.n84 VTAIL.n60 9.45567
R811 VTAIL.n204 VTAIL.n180 9.45567
R812 VTAIL.n174 VTAIL.n150 9.45567
R813 VTAIL.n144 VTAIL.n120 9.45567
R814 VTAIL.n114 VTAIL.n90 9.45567
R815 VTAIL.n218 VTAIL.n217 9.3005
R816 VTAIL.n225 VTAIL.n224 9.3005
R817 VTAIL.n227 VTAIL.n226 9.3005
R818 VTAIL.n214 VTAIL.n213 9.3005
R819 VTAIL.n233 VTAIL.n232 9.3005
R820 VTAIL.n235 VTAIL.n234 9.3005
R821 VTAIL.n8 VTAIL.n7 9.3005
R822 VTAIL.n15 VTAIL.n14 9.3005
R823 VTAIL.n17 VTAIL.n16 9.3005
R824 VTAIL.n4 VTAIL.n3 9.3005
R825 VTAIL.n23 VTAIL.n22 9.3005
R826 VTAIL.n25 VTAIL.n24 9.3005
R827 VTAIL.n38 VTAIL.n37 9.3005
R828 VTAIL.n45 VTAIL.n44 9.3005
R829 VTAIL.n47 VTAIL.n46 9.3005
R830 VTAIL.n34 VTAIL.n33 9.3005
R831 VTAIL.n53 VTAIL.n52 9.3005
R832 VTAIL.n55 VTAIL.n54 9.3005
R833 VTAIL.n68 VTAIL.n67 9.3005
R834 VTAIL.n75 VTAIL.n74 9.3005
R835 VTAIL.n77 VTAIL.n76 9.3005
R836 VTAIL.n64 VTAIL.n63 9.3005
R837 VTAIL.n83 VTAIL.n82 9.3005
R838 VTAIL.n85 VTAIL.n84 9.3005
R839 VTAIL.n205 VTAIL.n204 9.3005
R840 VTAIL.n203 VTAIL.n202 9.3005
R841 VTAIL.n184 VTAIL.n183 9.3005
R842 VTAIL.n197 VTAIL.n196 9.3005
R843 VTAIL.n195 VTAIL.n194 9.3005
R844 VTAIL.n188 VTAIL.n187 9.3005
R845 VTAIL.n165 VTAIL.n164 9.3005
R846 VTAIL.n167 VTAIL.n166 9.3005
R847 VTAIL.n154 VTAIL.n153 9.3005
R848 VTAIL.n173 VTAIL.n172 9.3005
R849 VTAIL.n175 VTAIL.n174 9.3005
R850 VTAIL.n158 VTAIL.n157 9.3005
R851 VTAIL.n135 VTAIL.n134 9.3005
R852 VTAIL.n137 VTAIL.n136 9.3005
R853 VTAIL.n124 VTAIL.n123 9.3005
R854 VTAIL.n143 VTAIL.n142 9.3005
R855 VTAIL.n145 VTAIL.n144 9.3005
R856 VTAIL.n128 VTAIL.n127 9.3005
R857 VTAIL.n105 VTAIL.n104 9.3005
R858 VTAIL.n107 VTAIL.n106 9.3005
R859 VTAIL.n94 VTAIL.n93 9.3005
R860 VTAIL.n113 VTAIL.n112 9.3005
R861 VTAIL.n115 VTAIL.n114 9.3005
R862 VTAIL.n98 VTAIL.n97 9.3005
R863 VTAIL.n227 VTAIL.n216 8.92171
R864 VTAIL.n17 VTAIL.n6 8.92171
R865 VTAIL.n47 VTAIL.n36 8.92171
R866 VTAIL.n77 VTAIL.n66 8.92171
R867 VTAIL.n197 VTAIL.n186 8.92171
R868 VTAIL.n167 VTAIL.n156 8.92171
R869 VTAIL.n137 VTAIL.n126 8.92171
R870 VTAIL.n107 VTAIL.n96 8.92171
R871 VTAIL.n224 VTAIL.n223 8.14595
R872 VTAIL.n14 VTAIL.n13 8.14595
R873 VTAIL.n44 VTAIL.n43 8.14595
R874 VTAIL.n74 VTAIL.n73 8.14595
R875 VTAIL.n194 VTAIL.n193 8.14595
R876 VTAIL.n164 VTAIL.n163 8.14595
R877 VTAIL.n134 VTAIL.n133 8.14595
R878 VTAIL.n104 VTAIL.n103 8.14595
R879 VTAIL.n220 VTAIL.n218 7.3702
R880 VTAIL.n10 VTAIL.n8 7.3702
R881 VTAIL.n40 VTAIL.n38 7.3702
R882 VTAIL.n70 VTAIL.n68 7.3702
R883 VTAIL.n190 VTAIL.n188 7.3702
R884 VTAIL.n160 VTAIL.n158 7.3702
R885 VTAIL.n130 VTAIL.n128 7.3702
R886 VTAIL.n100 VTAIL.n98 7.3702
R887 VTAIL.n223 VTAIL.n218 5.81868
R888 VTAIL.n13 VTAIL.n8 5.81868
R889 VTAIL.n43 VTAIL.n38 5.81868
R890 VTAIL.n73 VTAIL.n68 5.81868
R891 VTAIL.n193 VTAIL.n188 5.81868
R892 VTAIL.n163 VTAIL.n158 5.81868
R893 VTAIL.n133 VTAIL.n128 5.81868
R894 VTAIL.n103 VTAIL.n98 5.81868
R895 VTAIL.n224 VTAIL.n216 5.04292
R896 VTAIL.n14 VTAIL.n6 5.04292
R897 VTAIL.n44 VTAIL.n36 5.04292
R898 VTAIL.n74 VTAIL.n66 5.04292
R899 VTAIL.n194 VTAIL.n186 5.04292
R900 VTAIL.n164 VTAIL.n156 5.04292
R901 VTAIL.n134 VTAIL.n126 5.04292
R902 VTAIL.n104 VTAIL.n96 5.04292
R903 VTAIL.n228 VTAIL.n227 4.26717
R904 VTAIL.n18 VTAIL.n17 4.26717
R905 VTAIL.n48 VTAIL.n47 4.26717
R906 VTAIL.n78 VTAIL.n77 4.26717
R907 VTAIL.n198 VTAIL.n197 4.26717
R908 VTAIL.n168 VTAIL.n167 4.26717
R909 VTAIL.n138 VTAIL.n137 4.26717
R910 VTAIL.n108 VTAIL.n107 4.26717
R911 VTAIL.n231 VTAIL.n214 3.49141
R912 VTAIL.n21 VTAIL.n4 3.49141
R913 VTAIL.n51 VTAIL.n34 3.49141
R914 VTAIL.n81 VTAIL.n64 3.49141
R915 VTAIL.n201 VTAIL.n184 3.49141
R916 VTAIL.n171 VTAIL.n154 3.49141
R917 VTAIL.n141 VTAIL.n124 3.49141
R918 VTAIL.n111 VTAIL.n94 3.49141
R919 VTAIL.n232 VTAIL.n212 2.71565
R920 VTAIL.n22 VTAIL.n2 2.71565
R921 VTAIL.n52 VTAIL.n32 2.71565
R922 VTAIL.n82 VTAIL.n62 2.71565
R923 VTAIL.n202 VTAIL.n182 2.71565
R924 VTAIL.n172 VTAIL.n152 2.71565
R925 VTAIL.n142 VTAIL.n122 2.71565
R926 VTAIL.n112 VTAIL.n92 2.71565
R927 VTAIL.n219 VTAIL.n217 2.4147
R928 VTAIL.n9 VTAIL.n7 2.4147
R929 VTAIL.n39 VTAIL.n37 2.4147
R930 VTAIL.n69 VTAIL.n67 2.4147
R931 VTAIL.n189 VTAIL.n187 2.4147
R932 VTAIL.n159 VTAIL.n157 2.4147
R933 VTAIL.n129 VTAIL.n127 2.4147
R934 VTAIL.n99 VTAIL.n97 2.4147
R935 VTAIL.n236 VTAIL.n235 1.93989
R936 VTAIL.n26 VTAIL.n25 1.93989
R937 VTAIL.n56 VTAIL.n55 1.93989
R938 VTAIL.n86 VTAIL.n85 1.93989
R939 VTAIL.n206 VTAIL.n205 1.93989
R940 VTAIL.n176 VTAIL.n175 1.93989
R941 VTAIL.n146 VTAIL.n145 1.93989
R942 VTAIL.n116 VTAIL.n115 1.93989
R943 VTAIL.n238 VTAIL.n210 1.16414
R944 VTAIL.n28 VTAIL.n0 1.16414
R945 VTAIL.n58 VTAIL.n30 1.16414
R946 VTAIL.n88 VTAIL.n60 1.16414
R947 VTAIL.n208 VTAIL.n180 1.16414
R948 VTAIL.n178 VTAIL.n150 1.16414
R949 VTAIL.n148 VTAIL.n120 1.16414
R950 VTAIL.n118 VTAIL.n90 1.16414
R951 VTAIL.n149 VTAIL.n119 1.14705
R952 VTAIL.n209 VTAIL.n179 1.14705
R953 VTAIL.n89 VTAIL.n59 1.14705
R954 VTAIL VTAIL.n29 0.631965
R955 VTAIL VTAIL.n239 0.515586
R956 VTAIL.n179 VTAIL.n149 0.470328
R957 VTAIL.n59 VTAIL.n29 0.470328
R958 VTAIL.n225 VTAIL.n217 0.155672
R959 VTAIL.n226 VTAIL.n225 0.155672
R960 VTAIL.n226 VTAIL.n213 0.155672
R961 VTAIL.n233 VTAIL.n213 0.155672
R962 VTAIL.n234 VTAIL.n233 0.155672
R963 VTAIL.n15 VTAIL.n7 0.155672
R964 VTAIL.n16 VTAIL.n15 0.155672
R965 VTAIL.n16 VTAIL.n3 0.155672
R966 VTAIL.n23 VTAIL.n3 0.155672
R967 VTAIL.n24 VTAIL.n23 0.155672
R968 VTAIL.n45 VTAIL.n37 0.155672
R969 VTAIL.n46 VTAIL.n45 0.155672
R970 VTAIL.n46 VTAIL.n33 0.155672
R971 VTAIL.n53 VTAIL.n33 0.155672
R972 VTAIL.n54 VTAIL.n53 0.155672
R973 VTAIL.n75 VTAIL.n67 0.155672
R974 VTAIL.n76 VTAIL.n75 0.155672
R975 VTAIL.n76 VTAIL.n63 0.155672
R976 VTAIL.n83 VTAIL.n63 0.155672
R977 VTAIL.n84 VTAIL.n83 0.155672
R978 VTAIL.n204 VTAIL.n203 0.155672
R979 VTAIL.n203 VTAIL.n183 0.155672
R980 VTAIL.n196 VTAIL.n183 0.155672
R981 VTAIL.n196 VTAIL.n195 0.155672
R982 VTAIL.n195 VTAIL.n187 0.155672
R983 VTAIL.n174 VTAIL.n173 0.155672
R984 VTAIL.n173 VTAIL.n153 0.155672
R985 VTAIL.n166 VTAIL.n153 0.155672
R986 VTAIL.n166 VTAIL.n165 0.155672
R987 VTAIL.n165 VTAIL.n157 0.155672
R988 VTAIL.n144 VTAIL.n143 0.155672
R989 VTAIL.n143 VTAIL.n123 0.155672
R990 VTAIL.n136 VTAIL.n123 0.155672
R991 VTAIL.n136 VTAIL.n135 0.155672
R992 VTAIL.n135 VTAIL.n127 0.155672
R993 VTAIL.n114 VTAIL.n113 0.155672
R994 VTAIL.n113 VTAIL.n93 0.155672
R995 VTAIL.n106 VTAIL.n93 0.155672
R996 VTAIL.n106 VTAIL.n105 0.155672
R997 VTAIL.n105 VTAIL.n97 0.155672
R998 VN.n0 VN.t1 199.117
R999 VN.n1 VN.t2 199.117
R1000 VN.n1 VN.t3 199.03
R1001 VN.n0 VN.t0 199.03
R1002 VN VN.n1 68.2887
R1003 VN VN.n0 31.2622
R1004 VDD2.n2 VDD2.n0 127.891
R1005 VDD2.n2 VDD2.n1 95.6936
R1006 VDD2.n1 VDD2.t0 5.55691
R1007 VDD2.n1 VDD2.t1 5.55691
R1008 VDD2.n0 VDD2.t2 5.55691
R1009 VDD2.n0 VDD2.t3 5.55691
R1010 VDD2 VDD2.n2 0.0586897
C0 VTAIL VP 1.92274f
C1 VDD1 VP 2.07771f
C2 VDD2 VP 0.292605f
C3 B VP 1.09258f
C4 VP VN 3.89981f
C5 w_n1768_n2138# VP 2.80535f
C6 VDD1 VTAIL 3.78709f
C7 VTAIL VDD2 3.83057f
C8 B VTAIL 2.29838f
C9 VTAIL VN 1.90863f
C10 VDD1 VDD2 0.638587f
C11 w_n1768_n2138# VTAIL 2.54871f
C12 B VDD1 0.813752f
C13 B VDD2 0.839886f
C14 VDD1 VN 0.147665f
C15 VDD2 VN 1.9331f
C16 B VN 0.729577f
C17 VDD1 w_n1768_n2138# 0.967312f
C18 w_n1768_n2138# VDD2 0.988032f
C19 B w_n1768_n2138# 5.55732f
C20 w_n1768_n2138# VN 2.58212f
C21 VDD2 VSUBS 0.524304f
C22 VDD1 VSUBS 4.014891f
C23 VTAIL VSUBS 0.51557f
C24 VN VSUBS 3.84679f
C25 VP VSUBS 1.169687f
C26 B VSUBS 2.368645f
C27 w_n1768_n2138# VSUBS 47.2056f
C28 VDD2.t2 VSUBS 0.08279f
C29 VDD2.t3 VSUBS 0.08279f
C30 VDD2.n0 VSUBS 0.78679f
C31 VDD2.t0 VSUBS 0.08279f
C32 VDD2.t1 VSUBS 0.08279f
C33 VDD2.n1 VSUBS 0.557661f
C34 VDD2.n2 VSUBS 2.05437f
C35 VN.t1 VSUBS 0.664606f
C36 VN.t0 VSUBS 0.664453f
C37 VN.n0 VSUBS 0.535584f
C38 VN.t2 VSUBS 0.664606f
C39 VN.t3 VSUBS 0.664453f
C40 VN.n1 VSUBS 1.27687f
C41 VTAIL.n0 VSUBS 0.011067f
C42 VTAIL.n1 VSUBS 0.024921f
C43 VTAIL.n2 VSUBS 0.011164f
C44 VTAIL.n3 VSUBS 0.019621f
C45 VTAIL.n4 VSUBS 0.010544f
C46 VTAIL.n5 VSUBS 0.024921f
C47 VTAIL.n6 VSUBS 0.011164f
C48 VTAIL.n7 VSUBS 0.434584f
C49 VTAIL.n8 VSUBS 0.010544f
C50 VTAIL.t3 VSUBS 0.053709f
C51 VTAIL.n9 VSUBS 0.100298f
C52 VTAIL.n10 VSUBS 0.018739f
C53 VTAIL.n11 VSUBS 0.018691f
C54 VTAIL.n12 VSUBS 0.024921f
C55 VTAIL.n13 VSUBS 0.011164f
C56 VTAIL.n14 VSUBS 0.010544f
C57 VTAIL.n15 VSUBS 0.019621f
C58 VTAIL.n16 VSUBS 0.019621f
C59 VTAIL.n17 VSUBS 0.010544f
C60 VTAIL.n18 VSUBS 0.011164f
C61 VTAIL.n19 VSUBS 0.024921f
C62 VTAIL.n20 VSUBS 0.024921f
C63 VTAIL.n21 VSUBS 0.011164f
C64 VTAIL.n22 VSUBS 0.010544f
C65 VTAIL.n23 VSUBS 0.019621f
C66 VTAIL.n24 VSUBS 0.050983f
C67 VTAIL.n25 VSUBS 0.010544f
C68 VTAIL.n26 VSUBS 0.011164f
C69 VTAIL.n27 VSUBS 0.055803f
C70 VTAIL.n28 VSUBS 0.03748f
C71 VTAIL.n29 VSUBS 0.08866f
C72 VTAIL.n30 VSUBS 0.011067f
C73 VTAIL.n31 VSUBS 0.024921f
C74 VTAIL.n32 VSUBS 0.011164f
C75 VTAIL.n33 VSUBS 0.019621f
C76 VTAIL.n34 VSUBS 0.010544f
C77 VTAIL.n35 VSUBS 0.024921f
C78 VTAIL.n36 VSUBS 0.011164f
C79 VTAIL.n37 VSUBS 0.434584f
C80 VTAIL.n38 VSUBS 0.010544f
C81 VTAIL.t6 VSUBS 0.053709f
C82 VTAIL.n39 VSUBS 0.100298f
C83 VTAIL.n40 VSUBS 0.018739f
C84 VTAIL.n41 VSUBS 0.018691f
C85 VTAIL.n42 VSUBS 0.024921f
C86 VTAIL.n43 VSUBS 0.011164f
C87 VTAIL.n44 VSUBS 0.010544f
C88 VTAIL.n45 VSUBS 0.019621f
C89 VTAIL.n46 VSUBS 0.019621f
C90 VTAIL.n47 VSUBS 0.010544f
C91 VTAIL.n48 VSUBS 0.011164f
C92 VTAIL.n49 VSUBS 0.024921f
C93 VTAIL.n50 VSUBS 0.024921f
C94 VTAIL.n51 VSUBS 0.011164f
C95 VTAIL.n52 VSUBS 0.010544f
C96 VTAIL.n53 VSUBS 0.019621f
C97 VTAIL.n54 VSUBS 0.050983f
C98 VTAIL.n55 VSUBS 0.010544f
C99 VTAIL.n56 VSUBS 0.011164f
C100 VTAIL.n57 VSUBS 0.055803f
C101 VTAIL.n58 VSUBS 0.03748f
C102 VTAIL.n59 VSUBS 0.121226f
C103 VTAIL.n60 VSUBS 0.011067f
C104 VTAIL.n61 VSUBS 0.024921f
C105 VTAIL.n62 VSUBS 0.011164f
C106 VTAIL.n63 VSUBS 0.019621f
C107 VTAIL.n64 VSUBS 0.010544f
C108 VTAIL.n65 VSUBS 0.024921f
C109 VTAIL.n66 VSUBS 0.011164f
C110 VTAIL.n67 VSUBS 0.434584f
C111 VTAIL.n68 VSUBS 0.010544f
C112 VTAIL.t7 VSUBS 0.053709f
C113 VTAIL.n69 VSUBS 0.100298f
C114 VTAIL.n70 VSUBS 0.018739f
C115 VTAIL.n71 VSUBS 0.018691f
C116 VTAIL.n72 VSUBS 0.024921f
C117 VTAIL.n73 VSUBS 0.011164f
C118 VTAIL.n74 VSUBS 0.010544f
C119 VTAIL.n75 VSUBS 0.019621f
C120 VTAIL.n76 VSUBS 0.019621f
C121 VTAIL.n77 VSUBS 0.010544f
C122 VTAIL.n78 VSUBS 0.011164f
C123 VTAIL.n79 VSUBS 0.024921f
C124 VTAIL.n80 VSUBS 0.024921f
C125 VTAIL.n81 VSUBS 0.011164f
C126 VTAIL.n82 VSUBS 0.010544f
C127 VTAIL.n83 VSUBS 0.019621f
C128 VTAIL.n84 VSUBS 0.050983f
C129 VTAIL.n85 VSUBS 0.010544f
C130 VTAIL.n86 VSUBS 0.011164f
C131 VTAIL.n87 VSUBS 0.055803f
C132 VTAIL.n88 VSUBS 0.03748f
C133 VTAIL.n89 VSUBS 0.749391f
C134 VTAIL.n90 VSUBS 0.011067f
C135 VTAIL.n91 VSUBS 0.024921f
C136 VTAIL.n92 VSUBS 0.011164f
C137 VTAIL.n93 VSUBS 0.019621f
C138 VTAIL.n94 VSUBS 0.010544f
C139 VTAIL.n95 VSUBS 0.024921f
C140 VTAIL.n96 VSUBS 0.011164f
C141 VTAIL.n97 VSUBS 0.434584f
C142 VTAIL.n98 VSUBS 0.010544f
C143 VTAIL.t2 VSUBS 0.053709f
C144 VTAIL.n99 VSUBS 0.100298f
C145 VTAIL.n100 VSUBS 0.018739f
C146 VTAIL.n101 VSUBS 0.018691f
C147 VTAIL.n102 VSUBS 0.024921f
C148 VTAIL.n103 VSUBS 0.011164f
C149 VTAIL.n104 VSUBS 0.010544f
C150 VTAIL.n105 VSUBS 0.019621f
C151 VTAIL.n106 VSUBS 0.019621f
C152 VTAIL.n107 VSUBS 0.010544f
C153 VTAIL.n108 VSUBS 0.011164f
C154 VTAIL.n109 VSUBS 0.024921f
C155 VTAIL.n110 VSUBS 0.024921f
C156 VTAIL.n111 VSUBS 0.011164f
C157 VTAIL.n112 VSUBS 0.010544f
C158 VTAIL.n113 VSUBS 0.019621f
C159 VTAIL.n114 VSUBS 0.050983f
C160 VTAIL.n115 VSUBS 0.010544f
C161 VTAIL.n116 VSUBS 0.011164f
C162 VTAIL.n117 VSUBS 0.055803f
C163 VTAIL.n118 VSUBS 0.03748f
C164 VTAIL.n119 VSUBS 0.749391f
C165 VTAIL.n120 VSUBS 0.011067f
C166 VTAIL.n121 VSUBS 0.024921f
C167 VTAIL.n122 VSUBS 0.011164f
C168 VTAIL.n123 VSUBS 0.019621f
C169 VTAIL.n124 VSUBS 0.010544f
C170 VTAIL.n125 VSUBS 0.024921f
C171 VTAIL.n126 VSUBS 0.011164f
C172 VTAIL.n127 VSUBS 0.434584f
C173 VTAIL.n128 VSUBS 0.010544f
C174 VTAIL.t0 VSUBS 0.053709f
C175 VTAIL.n129 VSUBS 0.100298f
C176 VTAIL.n130 VSUBS 0.018739f
C177 VTAIL.n131 VSUBS 0.018691f
C178 VTAIL.n132 VSUBS 0.024921f
C179 VTAIL.n133 VSUBS 0.011164f
C180 VTAIL.n134 VSUBS 0.010544f
C181 VTAIL.n135 VSUBS 0.019621f
C182 VTAIL.n136 VSUBS 0.019621f
C183 VTAIL.n137 VSUBS 0.010544f
C184 VTAIL.n138 VSUBS 0.011164f
C185 VTAIL.n139 VSUBS 0.024921f
C186 VTAIL.n140 VSUBS 0.024921f
C187 VTAIL.n141 VSUBS 0.011164f
C188 VTAIL.n142 VSUBS 0.010544f
C189 VTAIL.n143 VSUBS 0.019621f
C190 VTAIL.n144 VSUBS 0.050983f
C191 VTAIL.n145 VSUBS 0.010544f
C192 VTAIL.n146 VSUBS 0.011164f
C193 VTAIL.n147 VSUBS 0.055803f
C194 VTAIL.n148 VSUBS 0.03748f
C195 VTAIL.n149 VSUBS 0.121226f
C196 VTAIL.n150 VSUBS 0.011067f
C197 VTAIL.n151 VSUBS 0.024921f
C198 VTAIL.n152 VSUBS 0.011164f
C199 VTAIL.n153 VSUBS 0.019621f
C200 VTAIL.n154 VSUBS 0.010544f
C201 VTAIL.n155 VSUBS 0.024921f
C202 VTAIL.n156 VSUBS 0.011164f
C203 VTAIL.n157 VSUBS 0.434584f
C204 VTAIL.n158 VSUBS 0.010544f
C205 VTAIL.t5 VSUBS 0.053709f
C206 VTAIL.n159 VSUBS 0.100298f
C207 VTAIL.n160 VSUBS 0.018739f
C208 VTAIL.n161 VSUBS 0.018691f
C209 VTAIL.n162 VSUBS 0.024921f
C210 VTAIL.n163 VSUBS 0.011164f
C211 VTAIL.n164 VSUBS 0.010544f
C212 VTAIL.n165 VSUBS 0.019621f
C213 VTAIL.n166 VSUBS 0.019621f
C214 VTAIL.n167 VSUBS 0.010544f
C215 VTAIL.n168 VSUBS 0.011164f
C216 VTAIL.n169 VSUBS 0.024921f
C217 VTAIL.n170 VSUBS 0.024921f
C218 VTAIL.n171 VSUBS 0.011164f
C219 VTAIL.n172 VSUBS 0.010544f
C220 VTAIL.n173 VSUBS 0.019621f
C221 VTAIL.n174 VSUBS 0.050983f
C222 VTAIL.n175 VSUBS 0.010544f
C223 VTAIL.n176 VSUBS 0.011164f
C224 VTAIL.n177 VSUBS 0.055803f
C225 VTAIL.n178 VSUBS 0.03748f
C226 VTAIL.n179 VSUBS 0.121226f
C227 VTAIL.n180 VSUBS 0.011067f
C228 VTAIL.n181 VSUBS 0.024921f
C229 VTAIL.n182 VSUBS 0.011164f
C230 VTAIL.n183 VSUBS 0.019621f
C231 VTAIL.n184 VSUBS 0.010544f
C232 VTAIL.n185 VSUBS 0.024921f
C233 VTAIL.n186 VSUBS 0.011164f
C234 VTAIL.n187 VSUBS 0.434584f
C235 VTAIL.n188 VSUBS 0.010544f
C236 VTAIL.t4 VSUBS 0.053709f
C237 VTAIL.n189 VSUBS 0.100298f
C238 VTAIL.n190 VSUBS 0.018739f
C239 VTAIL.n191 VSUBS 0.018691f
C240 VTAIL.n192 VSUBS 0.024921f
C241 VTAIL.n193 VSUBS 0.011164f
C242 VTAIL.n194 VSUBS 0.010544f
C243 VTAIL.n195 VSUBS 0.019621f
C244 VTAIL.n196 VSUBS 0.019621f
C245 VTAIL.n197 VSUBS 0.010544f
C246 VTAIL.n198 VSUBS 0.011164f
C247 VTAIL.n199 VSUBS 0.024921f
C248 VTAIL.n200 VSUBS 0.024921f
C249 VTAIL.n201 VSUBS 0.011164f
C250 VTAIL.n202 VSUBS 0.010544f
C251 VTAIL.n203 VSUBS 0.019621f
C252 VTAIL.n204 VSUBS 0.050983f
C253 VTAIL.n205 VSUBS 0.010544f
C254 VTAIL.n206 VSUBS 0.011164f
C255 VTAIL.n207 VSUBS 0.055803f
C256 VTAIL.n208 VSUBS 0.03748f
C257 VTAIL.n209 VSUBS 0.74939f
C258 VTAIL.n210 VSUBS 0.011067f
C259 VTAIL.n211 VSUBS 0.024921f
C260 VTAIL.n212 VSUBS 0.011164f
C261 VTAIL.n213 VSUBS 0.019621f
C262 VTAIL.n214 VSUBS 0.010544f
C263 VTAIL.n215 VSUBS 0.024921f
C264 VTAIL.n216 VSUBS 0.011164f
C265 VTAIL.n217 VSUBS 0.434584f
C266 VTAIL.n218 VSUBS 0.010544f
C267 VTAIL.t1 VSUBS 0.053709f
C268 VTAIL.n219 VSUBS 0.100298f
C269 VTAIL.n220 VSUBS 0.018739f
C270 VTAIL.n221 VSUBS 0.018691f
C271 VTAIL.n222 VSUBS 0.024921f
C272 VTAIL.n223 VSUBS 0.011164f
C273 VTAIL.n224 VSUBS 0.010544f
C274 VTAIL.n225 VSUBS 0.019621f
C275 VTAIL.n226 VSUBS 0.019621f
C276 VTAIL.n227 VSUBS 0.010544f
C277 VTAIL.n228 VSUBS 0.011164f
C278 VTAIL.n229 VSUBS 0.024921f
C279 VTAIL.n230 VSUBS 0.024921f
C280 VTAIL.n231 VSUBS 0.011164f
C281 VTAIL.n232 VSUBS 0.010544f
C282 VTAIL.n233 VSUBS 0.019621f
C283 VTAIL.n234 VSUBS 0.050983f
C284 VTAIL.n235 VSUBS 0.010544f
C285 VTAIL.n236 VSUBS 0.011164f
C286 VTAIL.n237 VSUBS 0.055803f
C287 VTAIL.n238 VSUBS 0.03748f
C288 VTAIL.n239 VSUBS 0.709467f
C289 VDD1.t0 VSUBS 0.126344f
C290 VDD1.t3 VSUBS 0.126344f
C291 VDD1.n0 VSUBS 0.851356f
C292 VDD1.t1 VSUBS 0.126344f
C293 VDD1.t2 VSUBS 0.126344f
C294 VDD1.n1 VSUBS 1.21921f
C295 VP.t3 VSUBS 0.90692f
C296 VP.t2 VSUBS 0.907129f
C297 VP.n0 VSUBS 1.7233f
C298 VP.n1 VSUBS 2.60618f
C299 VP.t0 VSUBS 0.869478f
C300 VP.n2 VSUBS 0.40238f
C301 VP.t1 VSUBS 0.869478f
C302 VP.n3 VSUBS 0.40238f
C303 VP.n4 VSUBS 0.065031f
C304 B.n0 VSUBS 0.005819f
C305 B.n1 VSUBS 0.005819f
C306 B.n2 VSUBS 0.009202f
C307 B.n3 VSUBS 0.009202f
C308 B.n4 VSUBS 0.009202f
C309 B.n5 VSUBS 0.009202f
C310 B.n6 VSUBS 0.009202f
C311 B.n7 VSUBS 0.009202f
C312 B.n8 VSUBS 0.009202f
C313 B.n9 VSUBS 0.009202f
C314 B.n10 VSUBS 0.009202f
C315 B.n11 VSUBS 0.009202f
C316 B.n12 VSUBS 0.020507f
C317 B.n13 VSUBS 0.009202f
C318 B.n14 VSUBS 0.009202f
C319 B.n15 VSUBS 0.009202f
C320 B.n16 VSUBS 0.009202f
C321 B.n17 VSUBS 0.009202f
C322 B.n18 VSUBS 0.009202f
C323 B.n19 VSUBS 0.009202f
C324 B.n20 VSUBS 0.009202f
C325 B.n21 VSUBS 0.009202f
C326 B.n22 VSUBS 0.009202f
C327 B.n23 VSUBS 0.009202f
C328 B.t8 VSUBS 0.113825f
C329 B.t7 VSUBS 0.12982f
C330 B.t6 VSUBS 0.342882f
C331 B.n24 VSUBS 0.229458f
C332 B.n25 VSUBS 0.193621f
C333 B.n26 VSUBS 0.02132f
C334 B.n27 VSUBS 0.009202f
C335 B.n28 VSUBS 0.009202f
C336 B.n29 VSUBS 0.009202f
C337 B.n30 VSUBS 0.009202f
C338 B.n31 VSUBS 0.009202f
C339 B.t2 VSUBS 0.113828f
C340 B.t1 VSUBS 0.129822f
C341 B.t0 VSUBS 0.342882f
C342 B.n32 VSUBS 0.229455f
C343 B.n33 VSUBS 0.193618f
C344 B.n34 VSUBS 0.009202f
C345 B.n35 VSUBS 0.009202f
C346 B.n36 VSUBS 0.009202f
C347 B.n37 VSUBS 0.009202f
C348 B.n38 VSUBS 0.009202f
C349 B.n39 VSUBS 0.009202f
C350 B.n40 VSUBS 0.009202f
C351 B.n41 VSUBS 0.009202f
C352 B.n42 VSUBS 0.009202f
C353 B.n43 VSUBS 0.009202f
C354 B.n44 VSUBS 0.009202f
C355 B.n45 VSUBS 0.019278f
C356 B.n46 VSUBS 0.009202f
C357 B.n47 VSUBS 0.009202f
C358 B.n48 VSUBS 0.009202f
C359 B.n49 VSUBS 0.009202f
C360 B.n50 VSUBS 0.009202f
C361 B.n51 VSUBS 0.009202f
C362 B.n52 VSUBS 0.009202f
C363 B.n53 VSUBS 0.009202f
C364 B.n54 VSUBS 0.009202f
C365 B.n55 VSUBS 0.009202f
C366 B.n56 VSUBS 0.009202f
C367 B.n57 VSUBS 0.009202f
C368 B.n58 VSUBS 0.009202f
C369 B.n59 VSUBS 0.009202f
C370 B.n60 VSUBS 0.009202f
C371 B.n61 VSUBS 0.009202f
C372 B.n62 VSUBS 0.009202f
C373 B.n63 VSUBS 0.009202f
C374 B.n64 VSUBS 0.009202f
C375 B.n65 VSUBS 0.019278f
C376 B.n66 VSUBS 0.009202f
C377 B.n67 VSUBS 0.009202f
C378 B.n68 VSUBS 0.009202f
C379 B.n69 VSUBS 0.009202f
C380 B.n70 VSUBS 0.009202f
C381 B.n71 VSUBS 0.009202f
C382 B.n72 VSUBS 0.009202f
C383 B.n73 VSUBS 0.009202f
C384 B.n74 VSUBS 0.009202f
C385 B.n75 VSUBS 0.009202f
C386 B.n76 VSUBS 0.009202f
C387 B.n77 VSUBS 0.009202f
C388 B.t4 VSUBS 0.113828f
C389 B.t5 VSUBS 0.129822f
C390 B.t3 VSUBS 0.342882f
C391 B.n78 VSUBS 0.229455f
C392 B.n79 VSUBS 0.193618f
C393 B.n80 VSUBS 0.009202f
C394 B.n81 VSUBS 0.009202f
C395 B.n82 VSUBS 0.009202f
C396 B.n83 VSUBS 0.009202f
C397 B.t10 VSUBS 0.113825f
C398 B.t11 VSUBS 0.12982f
C399 B.t9 VSUBS 0.342882f
C400 B.n84 VSUBS 0.229458f
C401 B.n85 VSUBS 0.193621f
C402 B.n86 VSUBS 0.02132f
C403 B.n87 VSUBS 0.009202f
C404 B.n88 VSUBS 0.009202f
C405 B.n89 VSUBS 0.009202f
C406 B.n90 VSUBS 0.009202f
C407 B.n91 VSUBS 0.009202f
C408 B.n92 VSUBS 0.009202f
C409 B.n93 VSUBS 0.009202f
C410 B.n94 VSUBS 0.009202f
C411 B.n95 VSUBS 0.009202f
C412 B.n96 VSUBS 0.009202f
C413 B.n97 VSUBS 0.009202f
C414 B.n98 VSUBS 0.020507f
C415 B.n99 VSUBS 0.009202f
C416 B.n100 VSUBS 0.009202f
C417 B.n101 VSUBS 0.009202f
C418 B.n102 VSUBS 0.009202f
C419 B.n103 VSUBS 0.009202f
C420 B.n104 VSUBS 0.009202f
C421 B.n105 VSUBS 0.009202f
C422 B.n106 VSUBS 0.009202f
C423 B.n107 VSUBS 0.009202f
C424 B.n108 VSUBS 0.009202f
C425 B.n109 VSUBS 0.009202f
C426 B.n110 VSUBS 0.009202f
C427 B.n111 VSUBS 0.009202f
C428 B.n112 VSUBS 0.009202f
C429 B.n113 VSUBS 0.009202f
C430 B.n114 VSUBS 0.009202f
C431 B.n115 VSUBS 0.009202f
C432 B.n116 VSUBS 0.009202f
C433 B.n117 VSUBS 0.009202f
C434 B.n118 VSUBS 0.009202f
C435 B.n119 VSUBS 0.009202f
C436 B.n120 VSUBS 0.009202f
C437 B.n121 VSUBS 0.009202f
C438 B.n122 VSUBS 0.009202f
C439 B.n123 VSUBS 0.009202f
C440 B.n124 VSUBS 0.009202f
C441 B.n125 VSUBS 0.009202f
C442 B.n126 VSUBS 0.009202f
C443 B.n127 VSUBS 0.009202f
C444 B.n128 VSUBS 0.009202f
C445 B.n129 VSUBS 0.009202f
C446 B.n130 VSUBS 0.009202f
C447 B.n131 VSUBS 0.009202f
C448 B.n132 VSUBS 0.009202f
C449 B.n133 VSUBS 0.009202f
C450 B.n134 VSUBS 0.009202f
C451 B.n135 VSUBS 0.019278f
C452 B.n136 VSUBS 0.019278f
C453 B.n137 VSUBS 0.020507f
C454 B.n138 VSUBS 0.009202f
C455 B.n139 VSUBS 0.009202f
C456 B.n140 VSUBS 0.009202f
C457 B.n141 VSUBS 0.009202f
C458 B.n142 VSUBS 0.009202f
C459 B.n143 VSUBS 0.009202f
C460 B.n144 VSUBS 0.009202f
C461 B.n145 VSUBS 0.009202f
C462 B.n146 VSUBS 0.009202f
C463 B.n147 VSUBS 0.009202f
C464 B.n148 VSUBS 0.009202f
C465 B.n149 VSUBS 0.009202f
C466 B.n150 VSUBS 0.009202f
C467 B.n151 VSUBS 0.009202f
C468 B.n152 VSUBS 0.009202f
C469 B.n153 VSUBS 0.009202f
C470 B.n154 VSUBS 0.009202f
C471 B.n155 VSUBS 0.009202f
C472 B.n156 VSUBS 0.009202f
C473 B.n157 VSUBS 0.009202f
C474 B.n158 VSUBS 0.009202f
C475 B.n159 VSUBS 0.009202f
C476 B.n160 VSUBS 0.009202f
C477 B.n161 VSUBS 0.009202f
C478 B.n162 VSUBS 0.009202f
C479 B.n163 VSUBS 0.009202f
C480 B.n164 VSUBS 0.009202f
C481 B.n165 VSUBS 0.009202f
C482 B.n166 VSUBS 0.009202f
C483 B.n167 VSUBS 0.009202f
C484 B.n168 VSUBS 0.009202f
C485 B.n169 VSUBS 0.009202f
C486 B.n170 VSUBS 0.009202f
C487 B.n171 VSUBS 0.00636f
C488 B.n172 VSUBS 0.009202f
C489 B.n173 VSUBS 0.009202f
C490 B.n174 VSUBS 0.007443f
C491 B.n175 VSUBS 0.009202f
C492 B.n176 VSUBS 0.009202f
C493 B.n177 VSUBS 0.009202f
C494 B.n178 VSUBS 0.009202f
C495 B.n179 VSUBS 0.009202f
C496 B.n180 VSUBS 0.009202f
C497 B.n181 VSUBS 0.009202f
C498 B.n182 VSUBS 0.009202f
C499 B.n183 VSUBS 0.009202f
C500 B.n184 VSUBS 0.009202f
C501 B.n185 VSUBS 0.009202f
C502 B.n186 VSUBS 0.007443f
C503 B.n187 VSUBS 0.02132f
C504 B.n188 VSUBS 0.00636f
C505 B.n189 VSUBS 0.009202f
C506 B.n190 VSUBS 0.009202f
C507 B.n191 VSUBS 0.009202f
C508 B.n192 VSUBS 0.009202f
C509 B.n193 VSUBS 0.009202f
C510 B.n194 VSUBS 0.009202f
C511 B.n195 VSUBS 0.009202f
C512 B.n196 VSUBS 0.009202f
C513 B.n197 VSUBS 0.009202f
C514 B.n198 VSUBS 0.009202f
C515 B.n199 VSUBS 0.009202f
C516 B.n200 VSUBS 0.009202f
C517 B.n201 VSUBS 0.009202f
C518 B.n202 VSUBS 0.009202f
C519 B.n203 VSUBS 0.009202f
C520 B.n204 VSUBS 0.009202f
C521 B.n205 VSUBS 0.009202f
C522 B.n206 VSUBS 0.009202f
C523 B.n207 VSUBS 0.009202f
C524 B.n208 VSUBS 0.009202f
C525 B.n209 VSUBS 0.009202f
C526 B.n210 VSUBS 0.009202f
C527 B.n211 VSUBS 0.009202f
C528 B.n212 VSUBS 0.009202f
C529 B.n213 VSUBS 0.009202f
C530 B.n214 VSUBS 0.009202f
C531 B.n215 VSUBS 0.009202f
C532 B.n216 VSUBS 0.009202f
C533 B.n217 VSUBS 0.009202f
C534 B.n218 VSUBS 0.009202f
C535 B.n219 VSUBS 0.009202f
C536 B.n220 VSUBS 0.009202f
C537 B.n221 VSUBS 0.009202f
C538 B.n222 VSUBS 0.020507f
C539 B.n223 VSUBS 0.020507f
C540 B.n224 VSUBS 0.019278f
C541 B.n225 VSUBS 0.009202f
C542 B.n226 VSUBS 0.009202f
C543 B.n227 VSUBS 0.009202f
C544 B.n228 VSUBS 0.009202f
C545 B.n229 VSUBS 0.009202f
C546 B.n230 VSUBS 0.009202f
C547 B.n231 VSUBS 0.009202f
C548 B.n232 VSUBS 0.009202f
C549 B.n233 VSUBS 0.009202f
C550 B.n234 VSUBS 0.009202f
C551 B.n235 VSUBS 0.009202f
C552 B.n236 VSUBS 0.009202f
C553 B.n237 VSUBS 0.009202f
C554 B.n238 VSUBS 0.009202f
C555 B.n239 VSUBS 0.009202f
C556 B.n240 VSUBS 0.009202f
C557 B.n241 VSUBS 0.009202f
C558 B.n242 VSUBS 0.009202f
C559 B.n243 VSUBS 0.009202f
C560 B.n244 VSUBS 0.009202f
C561 B.n245 VSUBS 0.009202f
C562 B.n246 VSUBS 0.009202f
C563 B.n247 VSUBS 0.009202f
C564 B.n248 VSUBS 0.009202f
C565 B.n249 VSUBS 0.009202f
C566 B.n250 VSUBS 0.009202f
C567 B.n251 VSUBS 0.009202f
C568 B.n252 VSUBS 0.009202f
C569 B.n253 VSUBS 0.009202f
C570 B.n254 VSUBS 0.009202f
C571 B.n255 VSUBS 0.009202f
C572 B.n256 VSUBS 0.009202f
C573 B.n257 VSUBS 0.009202f
C574 B.n258 VSUBS 0.009202f
C575 B.n259 VSUBS 0.009202f
C576 B.n260 VSUBS 0.009202f
C577 B.n261 VSUBS 0.009202f
C578 B.n262 VSUBS 0.009202f
C579 B.n263 VSUBS 0.009202f
C580 B.n264 VSUBS 0.009202f
C581 B.n265 VSUBS 0.009202f
C582 B.n266 VSUBS 0.009202f
C583 B.n267 VSUBS 0.009202f
C584 B.n268 VSUBS 0.009202f
C585 B.n269 VSUBS 0.009202f
C586 B.n270 VSUBS 0.009202f
C587 B.n271 VSUBS 0.009202f
C588 B.n272 VSUBS 0.009202f
C589 B.n273 VSUBS 0.009202f
C590 B.n274 VSUBS 0.009202f
C591 B.n275 VSUBS 0.009202f
C592 B.n276 VSUBS 0.009202f
C593 B.n277 VSUBS 0.009202f
C594 B.n278 VSUBS 0.009202f
C595 B.n279 VSUBS 0.009202f
C596 B.n280 VSUBS 0.009202f
C597 B.n281 VSUBS 0.009202f
C598 B.n282 VSUBS 0.009202f
C599 B.n283 VSUBS 0.009202f
C600 B.n284 VSUBS 0.020507f
C601 B.n285 VSUBS 0.019278f
C602 B.n286 VSUBS 0.020507f
C603 B.n287 VSUBS 0.009202f
C604 B.n288 VSUBS 0.009202f
C605 B.n289 VSUBS 0.009202f
C606 B.n290 VSUBS 0.009202f
C607 B.n291 VSUBS 0.009202f
C608 B.n292 VSUBS 0.009202f
C609 B.n293 VSUBS 0.009202f
C610 B.n294 VSUBS 0.009202f
C611 B.n295 VSUBS 0.009202f
C612 B.n296 VSUBS 0.009202f
C613 B.n297 VSUBS 0.009202f
C614 B.n298 VSUBS 0.009202f
C615 B.n299 VSUBS 0.009202f
C616 B.n300 VSUBS 0.009202f
C617 B.n301 VSUBS 0.009202f
C618 B.n302 VSUBS 0.009202f
C619 B.n303 VSUBS 0.009202f
C620 B.n304 VSUBS 0.009202f
C621 B.n305 VSUBS 0.009202f
C622 B.n306 VSUBS 0.009202f
C623 B.n307 VSUBS 0.009202f
C624 B.n308 VSUBS 0.009202f
C625 B.n309 VSUBS 0.009202f
C626 B.n310 VSUBS 0.009202f
C627 B.n311 VSUBS 0.009202f
C628 B.n312 VSUBS 0.009202f
C629 B.n313 VSUBS 0.009202f
C630 B.n314 VSUBS 0.009202f
C631 B.n315 VSUBS 0.009202f
C632 B.n316 VSUBS 0.009202f
C633 B.n317 VSUBS 0.009202f
C634 B.n318 VSUBS 0.009202f
C635 B.n319 VSUBS 0.009202f
C636 B.n320 VSUBS 0.00636f
C637 B.n321 VSUBS 0.02132f
C638 B.n322 VSUBS 0.007443f
C639 B.n323 VSUBS 0.009202f
C640 B.n324 VSUBS 0.009202f
C641 B.n325 VSUBS 0.009202f
C642 B.n326 VSUBS 0.009202f
C643 B.n327 VSUBS 0.009202f
C644 B.n328 VSUBS 0.009202f
C645 B.n329 VSUBS 0.009202f
C646 B.n330 VSUBS 0.009202f
C647 B.n331 VSUBS 0.009202f
C648 B.n332 VSUBS 0.009202f
C649 B.n333 VSUBS 0.009202f
C650 B.n334 VSUBS 0.007443f
C651 B.n335 VSUBS 0.009202f
C652 B.n336 VSUBS 0.009202f
C653 B.n337 VSUBS 0.00636f
C654 B.n338 VSUBS 0.009202f
C655 B.n339 VSUBS 0.009202f
C656 B.n340 VSUBS 0.009202f
C657 B.n341 VSUBS 0.009202f
C658 B.n342 VSUBS 0.009202f
C659 B.n343 VSUBS 0.009202f
C660 B.n344 VSUBS 0.009202f
C661 B.n345 VSUBS 0.009202f
C662 B.n346 VSUBS 0.009202f
C663 B.n347 VSUBS 0.009202f
C664 B.n348 VSUBS 0.009202f
C665 B.n349 VSUBS 0.009202f
C666 B.n350 VSUBS 0.009202f
C667 B.n351 VSUBS 0.009202f
C668 B.n352 VSUBS 0.009202f
C669 B.n353 VSUBS 0.009202f
C670 B.n354 VSUBS 0.009202f
C671 B.n355 VSUBS 0.009202f
C672 B.n356 VSUBS 0.009202f
C673 B.n357 VSUBS 0.009202f
C674 B.n358 VSUBS 0.009202f
C675 B.n359 VSUBS 0.009202f
C676 B.n360 VSUBS 0.009202f
C677 B.n361 VSUBS 0.009202f
C678 B.n362 VSUBS 0.009202f
C679 B.n363 VSUBS 0.009202f
C680 B.n364 VSUBS 0.009202f
C681 B.n365 VSUBS 0.009202f
C682 B.n366 VSUBS 0.009202f
C683 B.n367 VSUBS 0.009202f
C684 B.n368 VSUBS 0.009202f
C685 B.n369 VSUBS 0.009202f
C686 B.n370 VSUBS 0.009202f
C687 B.n371 VSUBS 0.020507f
C688 B.n372 VSUBS 0.019278f
C689 B.n373 VSUBS 0.019278f
C690 B.n374 VSUBS 0.009202f
C691 B.n375 VSUBS 0.009202f
C692 B.n376 VSUBS 0.009202f
C693 B.n377 VSUBS 0.009202f
C694 B.n378 VSUBS 0.009202f
C695 B.n379 VSUBS 0.009202f
C696 B.n380 VSUBS 0.009202f
C697 B.n381 VSUBS 0.009202f
C698 B.n382 VSUBS 0.009202f
C699 B.n383 VSUBS 0.009202f
C700 B.n384 VSUBS 0.009202f
C701 B.n385 VSUBS 0.009202f
C702 B.n386 VSUBS 0.009202f
C703 B.n387 VSUBS 0.009202f
C704 B.n388 VSUBS 0.009202f
C705 B.n389 VSUBS 0.009202f
C706 B.n390 VSUBS 0.009202f
C707 B.n391 VSUBS 0.009202f
C708 B.n392 VSUBS 0.009202f
C709 B.n393 VSUBS 0.009202f
C710 B.n394 VSUBS 0.009202f
C711 B.n395 VSUBS 0.009202f
C712 B.n396 VSUBS 0.009202f
C713 B.n397 VSUBS 0.009202f
C714 B.n398 VSUBS 0.009202f
C715 B.n399 VSUBS 0.009202f
C716 B.n400 VSUBS 0.009202f
C717 B.n401 VSUBS 0.009202f
C718 B.n402 VSUBS 0.009202f
C719 B.n403 VSUBS 0.020836f
.ends

