* NGSPICE file created from diff_pair_sample_1171.ext - technology: sky130A

.subckt diff_pair_sample_1171 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t9 VN.t0 VTAIL.t16 w_n4666_n2018# sky130_fd_pr__pfet_01v8 ad=0.86625 pd=5.58 as=2.0475 ps=11.28 w=5.25 l=2.75
X1 VDD1.t9 VP.t0 VTAIL.t0 w_n4666_n2018# sky130_fd_pr__pfet_01v8 ad=0.86625 pd=5.58 as=2.0475 ps=11.28 w=5.25 l=2.75
X2 VDD1.t8 VP.t1 VTAIL.t2 w_n4666_n2018# sky130_fd_pr__pfet_01v8 ad=0.86625 pd=5.58 as=2.0475 ps=11.28 w=5.25 l=2.75
X3 VDD1.t7 VP.t2 VTAIL.t6 w_n4666_n2018# sky130_fd_pr__pfet_01v8 ad=2.0475 pd=11.28 as=0.86625 ps=5.58 w=5.25 l=2.75
X4 B.t11 B.t9 B.t10 w_n4666_n2018# sky130_fd_pr__pfet_01v8 ad=2.0475 pd=11.28 as=0 ps=0 w=5.25 l=2.75
X5 B.t8 B.t6 B.t7 w_n4666_n2018# sky130_fd_pr__pfet_01v8 ad=2.0475 pd=11.28 as=0 ps=0 w=5.25 l=2.75
X6 VDD2.t8 VN.t1 VTAIL.t14 w_n4666_n2018# sky130_fd_pr__pfet_01v8 ad=0.86625 pd=5.58 as=2.0475 ps=11.28 w=5.25 l=2.75
X7 VTAIL.t13 VN.t2 VDD2.t7 w_n4666_n2018# sky130_fd_pr__pfet_01v8 ad=0.86625 pd=5.58 as=0.86625 ps=5.58 w=5.25 l=2.75
X8 VTAIL.t18 VN.t3 VDD2.t6 w_n4666_n2018# sky130_fd_pr__pfet_01v8 ad=0.86625 pd=5.58 as=0.86625 ps=5.58 w=5.25 l=2.75
X9 VTAIL.t5 VP.t3 VDD1.t6 w_n4666_n2018# sky130_fd_pr__pfet_01v8 ad=0.86625 pd=5.58 as=0.86625 ps=5.58 w=5.25 l=2.75
X10 VDD2.t5 VN.t4 VTAIL.t10 w_n4666_n2018# sky130_fd_pr__pfet_01v8 ad=0.86625 pd=5.58 as=0.86625 ps=5.58 w=5.25 l=2.75
X11 VDD2.t4 VN.t5 VTAIL.t11 w_n4666_n2018# sky130_fd_pr__pfet_01v8 ad=2.0475 pd=11.28 as=0.86625 ps=5.58 w=5.25 l=2.75
X12 VTAIL.t19 VN.t6 VDD2.t3 w_n4666_n2018# sky130_fd_pr__pfet_01v8 ad=0.86625 pd=5.58 as=0.86625 ps=5.58 w=5.25 l=2.75
X13 VDD1.t5 VP.t4 VTAIL.t3 w_n4666_n2018# sky130_fd_pr__pfet_01v8 ad=2.0475 pd=11.28 as=0.86625 ps=5.58 w=5.25 l=2.75
X14 VDD1.t4 VP.t5 VTAIL.t7 w_n4666_n2018# sky130_fd_pr__pfet_01v8 ad=0.86625 pd=5.58 as=0.86625 ps=5.58 w=5.25 l=2.75
X15 VTAIL.t4 VP.t6 VDD1.t3 w_n4666_n2018# sky130_fd_pr__pfet_01v8 ad=0.86625 pd=5.58 as=0.86625 ps=5.58 w=5.25 l=2.75
X16 VDD2.t2 VN.t7 VTAIL.t12 w_n4666_n2018# sky130_fd_pr__pfet_01v8 ad=0.86625 pd=5.58 as=0.86625 ps=5.58 w=5.25 l=2.75
X17 VDD1.t2 VP.t7 VTAIL.t9 w_n4666_n2018# sky130_fd_pr__pfet_01v8 ad=0.86625 pd=5.58 as=0.86625 ps=5.58 w=5.25 l=2.75
X18 VTAIL.t1 VP.t8 VDD1.t1 w_n4666_n2018# sky130_fd_pr__pfet_01v8 ad=0.86625 pd=5.58 as=0.86625 ps=5.58 w=5.25 l=2.75
X19 VTAIL.t8 VP.t9 VDD1.t0 w_n4666_n2018# sky130_fd_pr__pfet_01v8 ad=0.86625 pd=5.58 as=0.86625 ps=5.58 w=5.25 l=2.75
X20 B.t5 B.t3 B.t4 w_n4666_n2018# sky130_fd_pr__pfet_01v8 ad=2.0475 pd=11.28 as=0 ps=0 w=5.25 l=2.75
X21 B.t2 B.t0 B.t1 w_n4666_n2018# sky130_fd_pr__pfet_01v8 ad=2.0475 pd=11.28 as=0 ps=0 w=5.25 l=2.75
X22 VDD2.t1 VN.t8 VTAIL.t15 w_n4666_n2018# sky130_fd_pr__pfet_01v8 ad=2.0475 pd=11.28 as=0.86625 ps=5.58 w=5.25 l=2.75
X23 VTAIL.t17 VN.t9 VDD2.t0 w_n4666_n2018# sky130_fd_pr__pfet_01v8 ad=0.86625 pd=5.58 as=0.86625 ps=5.58 w=5.25 l=2.75
R0 VN.n83 VN.n43 161.3
R1 VN.n82 VN.n81 161.3
R2 VN.n80 VN.n44 161.3
R3 VN.n79 VN.n78 161.3
R4 VN.n77 VN.n45 161.3
R5 VN.n76 VN.n75 161.3
R6 VN.n74 VN.n73 161.3
R7 VN.n72 VN.n47 161.3
R8 VN.n71 VN.n70 161.3
R9 VN.n69 VN.n48 161.3
R10 VN.n68 VN.n67 161.3
R11 VN.n66 VN.n49 161.3
R12 VN.n65 VN.n64 161.3
R13 VN.n63 VN.n50 161.3
R14 VN.n62 VN.n61 161.3
R15 VN.n60 VN.n51 161.3
R16 VN.n59 VN.n58 161.3
R17 VN.n57 VN.n52 161.3
R18 VN.n56 VN.n55 161.3
R19 VN.n40 VN.n0 161.3
R20 VN.n39 VN.n38 161.3
R21 VN.n37 VN.n1 161.3
R22 VN.n36 VN.n35 161.3
R23 VN.n34 VN.n2 161.3
R24 VN.n33 VN.n32 161.3
R25 VN.n31 VN.n30 161.3
R26 VN.n29 VN.n4 161.3
R27 VN.n28 VN.n27 161.3
R28 VN.n26 VN.n5 161.3
R29 VN.n25 VN.n24 161.3
R30 VN.n23 VN.n6 161.3
R31 VN.n22 VN.n21 161.3
R32 VN.n20 VN.n7 161.3
R33 VN.n19 VN.n18 161.3
R34 VN.n17 VN.n8 161.3
R35 VN.n16 VN.n15 161.3
R36 VN.n14 VN.n9 161.3
R37 VN.n13 VN.n12 161.3
R38 VN.n42 VN.n41 102.927
R39 VN.n85 VN.n84 102.927
R40 VN.n10 VN.t8 78.9128
R41 VN.n53 VN.t1 78.9128
R42 VN.n11 VN.n10 68.8984
R43 VN.n54 VN.n53 68.8984
R44 VN.n35 VN.n1 52.1486
R45 VN.n78 VN.n44 52.1486
R46 VN VN.n85 49.1194
R47 VN.n22 VN.t7 46.0096
R48 VN.n11 VN.t6 46.0096
R49 VN.n3 VN.t9 46.0096
R50 VN.n41 VN.t0 46.0096
R51 VN.n65 VN.t4 46.0096
R52 VN.n54 VN.t2 46.0096
R53 VN.n46 VN.t3 46.0096
R54 VN.n84 VN.t5 46.0096
R55 VN.n17 VN.n16 44.3785
R56 VN.n28 VN.n5 44.3785
R57 VN.n60 VN.n59 44.3785
R58 VN.n71 VN.n48 44.3785
R59 VN.n18 VN.n17 36.6083
R60 VN.n24 VN.n5 36.6083
R61 VN.n61 VN.n60 36.6083
R62 VN.n67 VN.n48 36.6083
R63 VN.n35 VN.n34 28.8382
R64 VN.n78 VN.n77 28.8382
R65 VN.n12 VN.n9 24.4675
R66 VN.n16 VN.n9 24.4675
R67 VN.n18 VN.n7 24.4675
R68 VN.n22 VN.n7 24.4675
R69 VN.n23 VN.n22 24.4675
R70 VN.n24 VN.n23 24.4675
R71 VN.n29 VN.n28 24.4675
R72 VN.n30 VN.n29 24.4675
R73 VN.n34 VN.n33 24.4675
R74 VN.n39 VN.n1 24.4675
R75 VN.n40 VN.n39 24.4675
R76 VN.n59 VN.n52 24.4675
R77 VN.n55 VN.n52 24.4675
R78 VN.n67 VN.n66 24.4675
R79 VN.n66 VN.n65 24.4675
R80 VN.n65 VN.n50 24.4675
R81 VN.n61 VN.n50 24.4675
R82 VN.n77 VN.n76 24.4675
R83 VN.n73 VN.n72 24.4675
R84 VN.n72 VN.n71 24.4675
R85 VN.n83 VN.n82 24.4675
R86 VN.n82 VN.n44 24.4675
R87 VN.n33 VN.n3 20.5528
R88 VN.n76 VN.n46 20.5528
R89 VN.n41 VN.n40 7.82994
R90 VN.n84 VN.n83 7.82994
R91 VN.n56 VN.n53 6.98708
R92 VN.n13 VN.n10 6.98708
R93 VN.n12 VN.n11 3.91522
R94 VN.n30 VN.n3 3.91522
R95 VN.n55 VN.n54 3.91522
R96 VN.n73 VN.n46 3.91522
R97 VN.n85 VN.n43 0.278367
R98 VN.n42 VN.n0 0.278367
R99 VN.n81 VN.n43 0.189894
R100 VN.n81 VN.n80 0.189894
R101 VN.n80 VN.n79 0.189894
R102 VN.n79 VN.n45 0.189894
R103 VN.n75 VN.n45 0.189894
R104 VN.n75 VN.n74 0.189894
R105 VN.n74 VN.n47 0.189894
R106 VN.n70 VN.n47 0.189894
R107 VN.n70 VN.n69 0.189894
R108 VN.n69 VN.n68 0.189894
R109 VN.n68 VN.n49 0.189894
R110 VN.n64 VN.n49 0.189894
R111 VN.n64 VN.n63 0.189894
R112 VN.n63 VN.n62 0.189894
R113 VN.n62 VN.n51 0.189894
R114 VN.n58 VN.n51 0.189894
R115 VN.n58 VN.n57 0.189894
R116 VN.n57 VN.n56 0.189894
R117 VN.n14 VN.n13 0.189894
R118 VN.n15 VN.n14 0.189894
R119 VN.n15 VN.n8 0.189894
R120 VN.n19 VN.n8 0.189894
R121 VN.n20 VN.n19 0.189894
R122 VN.n21 VN.n20 0.189894
R123 VN.n21 VN.n6 0.189894
R124 VN.n25 VN.n6 0.189894
R125 VN.n26 VN.n25 0.189894
R126 VN.n27 VN.n26 0.189894
R127 VN.n27 VN.n4 0.189894
R128 VN.n31 VN.n4 0.189894
R129 VN.n32 VN.n31 0.189894
R130 VN.n32 VN.n2 0.189894
R131 VN.n36 VN.n2 0.189894
R132 VN.n37 VN.n36 0.189894
R133 VN.n38 VN.n37 0.189894
R134 VN.n38 VN.n0 0.189894
R135 VN VN.n42 0.153454
R136 VTAIL.n120 VTAIL.n98 756.745
R137 VTAIL.n24 VTAIL.n2 756.745
R138 VTAIL.n92 VTAIL.n70 756.745
R139 VTAIL.n60 VTAIL.n38 756.745
R140 VTAIL.n106 VTAIL.n105 585
R141 VTAIL.n111 VTAIL.n110 585
R142 VTAIL.n113 VTAIL.n112 585
R143 VTAIL.n102 VTAIL.n101 585
R144 VTAIL.n119 VTAIL.n118 585
R145 VTAIL.n121 VTAIL.n120 585
R146 VTAIL.n10 VTAIL.n9 585
R147 VTAIL.n15 VTAIL.n14 585
R148 VTAIL.n17 VTAIL.n16 585
R149 VTAIL.n6 VTAIL.n5 585
R150 VTAIL.n23 VTAIL.n22 585
R151 VTAIL.n25 VTAIL.n24 585
R152 VTAIL.n93 VTAIL.n92 585
R153 VTAIL.n91 VTAIL.n90 585
R154 VTAIL.n74 VTAIL.n73 585
R155 VTAIL.n85 VTAIL.n84 585
R156 VTAIL.n83 VTAIL.n82 585
R157 VTAIL.n78 VTAIL.n77 585
R158 VTAIL.n61 VTAIL.n60 585
R159 VTAIL.n59 VTAIL.n58 585
R160 VTAIL.n42 VTAIL.n41 585
R161 VTAIL.n53 VTAIL.n52 585
R162 VTAIL.n51 VTAIL.n50 585
R163 VTAIL.n46 VTAIL.n45 585
R164 VTAIL.n107 VTAIL.t16 327.856
R165 VTAIL.n11 VTAIL.t0 327.856
R166 VTAIL.n79 VTAIL.t2 327.856
R167 VTAIL.n47 VTAIL.t14 327.856
R168 VTAIL.n111 VTAIL.n105 171.744
R169 VTAIL.n112 VTAIL.n111 171.744
R170 VTAIL.n112 VTAIL.n101 171.744
R171 VTAIL.n119 VTAIL.n101 171.744
R172 VTAIL.n120 VTAIL.n119 171.744
R173 VTAIL.n15 VTAIL.n9 171.744
R174 VTAIL.n16 VTAIL.n15 171.744
R175 VTAIL.n16 VTAIL.n5 171.744
R176 VTAIL.n23 VTAIL.n5 171.744
R177 VTAIL.n24 VTAIL.n23 171.744
R178 VTAIL.n92 VTAIL.n91 171.744
R179 VTAIL.n91 VTAIL.n73 171.744
R180 VTAIL.n84 VTAIL.n73 171.744
R181 VTAIL.n84 VTAIL.n83 171.744
R182 VTAIL.n83 VTAIL.n77 171.744
R183 VTAIL.n60 VTAIL.n59 171.744
R184 VTAIL.n59 VTAIL.n41 171.744
R185 VTAIL.n52 VTAIL.n41 171.744
R186 VTAIL.n52 VTAIL.n51 171.744
R187 VTAIL.n51 VTAIL.n45 171.744
R188 VTAIL.t16 VTAIL.n105 85.8723
R189 VTAIL.t0 VTAIL.n9 85.8723
R190 VTAIL.t2 VTAIL.n77 85.8723
R191 VTAIL.t14 VTAIL.n45 85.8723
R192 VTAIL.n69 VTAIL.n68 80.0703
R193 VTAIL.n67 VTAIL.n66 80.0703
R194 VTAIL.n37 VTAIL.n36 80.0703
R195 VTAIL.n35 VTAIL.n34 80.0703
R196 VTAIL.n127 VTAIL.n126 80.0702
R197 VTAIL.n1 VTAIL.n0 80.0702
R198 VTAIL.n31 VTAIL.n30 80.0702
R199 VTAIL.n33 VTAIL.n32 80.0702
R200 VTAIL.n125 VTAIL.n124 31.6035
R201 VTAIL.n29 VTAIL.n28 31.6035
R202 VTAIL.n97 VTAIL.n96 31.6035
R203 VTAIL.n65 VTAIL.n64 31.6035
R204 VTAIL.n35 VTAIL.n33 22.2031
R205 VTAIL.n125 VTAIL.n97 19.5479
R206 VTAIL.n107 VTAIL.n106 16.381
R207 VTAIL.n11 VTAIL.n10 16.381
R208 VTAIL.n79 VTAIL.n78 16.381
R209 VTAIL.n47 VTAIL.n46 16.381
R210 VTAIL.n110 VTAIL.n109 12.8005
R211 VTAIL.n14 VTAIL.n13 12.8005
R212 VTAIL.n82 VTAIL.n81 12.8005
R213 VTAIL.n50 VTAIL.n49 12.8005
R214 VTAIL.n113 VTAIL.n104 12.0247
R215 VTAIL.n17 VTAIL.n8 12.0247
R216 VTAIL.n85 VTAIL.n76 12.0247
R217 VTAIL.n53 VTAIL.n44 12.0247
R218 VTAIL.n114 VTAIL.n102 11.249
R219 VTAIL.n18 VTAIL.n6 11.249
R220 VTAIL.n86 VTAIL.n74 11.249
R221 VTAIL.n54 VTAIL.n42 11.249
R222 VTAIL.n118 VTAIL.n117 10.4732
R223 VTAIL.n22 VTAIL.n21 10.4732
R224 VTAIL.n90 VTAIL.n89 10.4732
R225 VTAIL.n58 VTAIL.n57 10.4732
R226 VTAIL.n121 VTAIL.n100 9.69747
R227 VTAIL.n25 VTAIL.n4 9.69747
R228 VTAIL.n93 VTAIL.n72 9.69747
R229 VTAIL.n61 VTAIL.n40 9.69747
R230 VTAIL.n124 VTAIL.n123 9.45567
R231 VTAIL.n28 VTAIL.n27 9.45567
R232 VTAIL.n96 VTAIL.n95 9.45567
R233 VTAIL.n64 VTAIL.n63 9.45567
R234 VTAIL.n123 VTAIL.n122 9.3005
R235 VTAIL.n100 VTAIL.n99 9.3005
R236 VTAIL.n117 VTAIL.n116 9.3005
R237 VTAIL.n115 VTAIL.n114 9.3005
R238 VTAIL.n104 VTAIL.n103 9.3005
R239 VTAIL.n109 VTAIL.n108 9.3005
R240 VTAIL.n27 VTAIL.n26 9.3005
R241 VTAIL.n4 VTAIL.n3 9.3005
R242 VTAIL.n21 VTAIL.n20 9.3005
R243 VTAIL.n19 VTAIL.n18 9.3005
R244 VTAIL.n8 VTAIL.n7 9.3005
R245 VTAIL.n13 VTAIL.n12 9.3005
R246 VTAIL.n95 VTAIL.n94 9.3005
R247 VTAIL.n72 VTAIL.n71 9.3005
R248 VTAIL.n89 VTAIL.n88 9.3005
R249 VTAIL.n87 VTAIL.n86 9.3005
R250 VTAIL.n76 VTAIL.n75 9.3005
R251 VTAIL.n81 VTAIL.n80 9.3005
R252 VTAIL.n63 VTAIL.n62 9.3005
R253 VTAIL.n40 VTAIL.n39 9.3005
R254 VTAIL.n57 VTAIL.n56 9.3005
R255 VTAIL.n55 VTAIL.n54 9.3005
R256 VTAIL.n44 VTAIL.n43 9.3005
R257 VTAIL.n49 VTAIL.n48 9.3005
R258 VTAIL.n122 VTAIL.n98 8.92171
R259 VTAIL.n26 VTAIL.n2 8.92171
R260 VTAIL.n94 VTAIL.n70 8.92171
R261 VTAIL.n62 VTAIL.n38 8.92171
R262 VTAIL.n126 VTAIL.t12 6.19193
R263 VTAIL.n126 VTAIL.t17 6.19193
R264 VTAIL.n0 VTAIL.t15 6.19193
R265 VTAIL.n0 VTAIL.t19 6.19193
R266 VTAIL.n30 VTAIL.t7 6.19193
R267 VTAIL.n30 VTAIL.t4 6.19193
R268 VTAIL.n32 VTAIL.t6 6.19193
R269 VTAIL.n32 VTAIL.t1 6.19193
R270 VTAIL.n68 VTAIL.t9 6.19193
R271 VTAIL.n68 VTAIL.t5 6.19193
R272 VTAIL.n66 VTAIL.t3 6.19193
R273 VTAIL.n66 VTAIL.t8 6.19193
R274 VTAIL.n36 VTAIL.t10 6.19193
R275 VTAIL.n36 VTAIL.t13 6.19193
R276 VTAIL.n34 VTAIL.t11 6.19193
R277 VTAIL.n34 VTAIL.t18 6.19193
R278 VTAIL.n124 VTAIL.n98 5.04292
R279 VTAIL.n28 VTAIL.n2 5.04292
R280 VTAIL.n96 VTAIL.n70 5.04292
R281 VTAIL.n64 VTAIL.n38 5.04292
R282 VTAIL.n122 VTAIL.n121 4.26717
R283 VTAIL.n26 VTAIL.n25 4.26717
R284 VTAIL.n94 VTAIL.n93 4.26717
R285 VTAIL.n62 VTAIL.n61 4.26717
R286 VTAIL.n80 VTAIL.n79 3.71853
R287 VTAIL.n48 VTAIL.n47 3.71853
R288 VTAIL.n108 VTAIL.n107 3.71853
R289 VTAIL.n12 VTAIL.n11 3.71853
R290 VTAIL.n118 VTAIL.n100 3.49141
R291 VTAIL.n22 VTAIL.n4 3.49141
R292 VTAIL.n90 VTAIL.n72 3.49141
R293 VTAIL.n58 VTAIL.n40 3.49141
R294 VTAIL.n117 VTAIL.n102 2.71565
R295 VTAIL.n21 VTAIL.n6 2.71565
R296 VTAIL.n89 VTAIL.n74 2.71565
R297 VTAIL.n57 VTAIL.n42 2.71565
R298 VTAIL.n37 VTAIL.n35 2.65567
R299 VTAIL.n65 VTAIL.n37 2.65567
R300 VTAIL.n69 VTAIL.n67 2.65567
R301 VTAIL.n97 VTAIL.n69 2.65567
R302 VTAIL.n33 VTAIL.n31 2.65567
R303 VTAIL.n31 VTAIL.n29 2.65567
R304 VTAIL.n127 VTAIL.n125 2.65567
R305 VTAIL VTAIL.n1 2.05007
R306 VTAIL.n114 VTAIL.n113 1.93989
R307 VTAIL.n18 VTAIL.n17 1.93989
R308 VTAIL.n86 VTAIL.n85 1.93989
R309 VTAIL.n54 VTAIL.n53 1.93989
R310 VTAIL.n67 VTAIL.n65 1.79791
R311 VTAIL.n29 VTAIL.n1 1.79791
R312 VTAIL.n110 VTAIL.n104 1.16414
R313 VTAIL.n14 VTAIL.n8 1.16414
R314 VTAIL.n82 VTAIL.n76 1.16414
R315 VTAIL.n50 VTAIL.n44 1.16414
R316 VTAIL VTAIL.n127 0.606103
R317 VTAIL.n109 VTAIL.n106 0.388379
R318 VTAIL.n13 VTAIL.n10 0.388379
R319 VTAIL.n81 VTAIL.n78 0.388379
R320 VTAIL.n49 VTAIL.n46 0.388379
R321 VTAIL.n108 VTAIL.n103 0.155672
R322 VTAIL.n115 VTAIL.n103 0.155672
R323 VTAIL.n116 VTAIL.n115 0.155672
R324 VTAIL.n116 VTAIL.n99 0.155672
R325 VTAIL.n123 VTAIL.n99 0.155672
R326 VTAIL.n12 VTAIL.n7 0.155672
R327 VTAIL.n19 VTAIL.n7 0.155672
R328 VTAIL.n20 VTAIL.n19 0.155672
R329 VTAIL.n20 VTAIL.n3 0.155672
R330 VTAIL.n27 VTAIL.n3 0.155672
R331 VTAIL.n95 VTAIL.n71 0.155672
R332 VTAIL.n88 VTAIL.n71 0.155672
R333 VTAIL.n88 VTAIL.n87 0.155672
R334 VTAIL.n87 VTAIL.n75 0.155672
R335 VTAIL.n80 VTAIL.n75 0.155672
R336 VTAIL.n63 VTAIL.n39 0.155672
R337 VTAIL.n56 VTAIL.n39 0.155672
R338 VTAIL.n56 VTAIL.n55 0.155672
R339 VTAIL.n55 VTAIL.n43 0.155672
R340 VTAIL.n48 VTAIL.n43 0.155672
R341 VDD2.n53 VDD2.n31 756.745
R342 VDD2.n22 VDD2.n0 756.745
R343 VDD2.n54 VDD2.n53 585
R344 VDD2.n52 VDD2.n51 585
R345 VDD2.n35 VDD2.n34 585
R346 VDD2.n46 VDD2.n45 585
R347 VDD2.n44 VDD2.n43 585
R348 VDD2.n39 VDD2.n38 585
R349 VDD2.n8 VDD2.n7 585
R350 VDD2.n13 VDD2.n12 585
R351 VDD2.n15 VDD2.n14 585
R352 VDD2.n4 VDD2.n3 585
R353 VDD2.n21 VDD2.n20 585
R354 VDD2.n23 VDD2.n22 585
R355 VDD2.n40 VDD2.t4 327.856
R356 VDD2.n9 VDD2.t1 327.856
R357 VDD2.n53 VDD2.n52 171.744
R358 VDD2.n52 VDD2.n34 171.744
R359 VDD2.n45 VDD2.n34 171.744
R360 VDD2.n45 VDD2.n44 171.744
R361 VDD2.n44 VDD2.n38 171.744
R362 VDD2.n13 VDD2.n7 171.744
R363 VDD2.n14 VDD2.n13 171.744
R364 VDD2.n14 VDD2.n3 171.744
R365 VDD2.n21 VDD2.n3 171.744
R366 VDD2.n22 VDD2.n21 171.744
R367 VDD2.n30 VDD2.n29 98.685
R368 VDD2 VDD2.n61 98.6821
R369 VDD2.n60 VDD2.n59 96.7491
R370 VDD2.n28 VDD2.n27 96.749
R371 VDD2.t4 VDD2.n38 85.8723
R372 VDD2.t1 VDD2.n7 85.8723
R373 VDD2.n28 VDD2.n26 50.9375
R374 VDD2.n58 VDD2.n57 48.2823
R375 VDD2.n58 VDD2.n30 40.8532
R376 VDD2.n40 VDD2.n39 16.381
R377 VDD2.n9 VDD2.n8 16.381
R378 VDD2.n43 VDD2.n42 12.8005
R379 VDD2.n12 VDD2.n11 12.8005
R380 VDD2.n46 VDD2.n37 12.0247
R381 VDD2.n15 VDD2.n6 12.0247
R382 VDD2.n47 VDD2.n35 11.249
R383 VDD2.n16 VDD2.n4 11.249
R384 VDD2.n51 VDD2.n50 10.4732
R385 VDD2.n20 VDD2.n19 10.4732
R386 VDD2.n54 VDD2.n33 9.69747
R387 VDD2.n23 VDD2.n2 9.69747
R388 VDD2.n57 VDD2.n56 9.45567
R389 VDD2.n26 VDD2.n25 9.45567
R390 VDD2.n56 VDD2.n55 9.3005
R391 VDD2.n33 VDD2.n32 9.3005
R392 VDD2.n50 VDD2.n49 9.3005
R393 VDD2.n48 VDD2.n47 9.3005
R394 VDD2.n37 VDD2.n36 9.3005
R395 VDD2.n42 VDD2.n41 9.3005
R396 VDD2.n25 VDD2.n24 9.3005
R397 VDD2.n2 VDD2.n1 9.3005
R398 VDD2.n19 VDD2.n18 9.3005
R399 VDD2.n17 VDD2.n16 9.3005
R400 VDD2.n6 VDD2.n5 9.3005
R401 VDD2.n11 VDD2.n10 9.3005
R402 VDD2.n55 VDD2.n31 8.92171
R403 VDD2.n24 VDD2.n0 8.92171
R404 VDD2.n61 VDD2.t7 6.19193
R405 VDD2.n61 VDD2.t8 6.19193
R406 VDD2.n59 VDD2.t6 6.19193
R407 VDD2.n59 VDD2.t5 6.19193
R408 VDD2.n29 VDD2.t0 6.19193
R409 VDD2.n29 VDD2.t9 6.19193
R410 VDD2.n27 VDD2.t3 6.19193
R411 VDD2.n27 VDD2.t2 6.19193
R412 VDD2.n57 VDD2.n31 5.04292
R413 VDD2.n26 VDD2.n0 5.04292
R414 VDD2.n55 VDD2.n54 4.26717
R415 VDD2.n24 VDD2.n23 4.26717
R416 VDD2.n41 VDD2.n40 3.71853
R417 VDD2.n10 VDD2.n9 3.71853
R418 VDD2.n51 VDD2.n33 3.49141
R419 VDD2.n20 VDD2.n2 3.49141
R420 VDD2.n50 VDD2.n35 2.71565
R421 VDD2.n19 VDD2.n4 2.71565
R422 VDD2.n60 VDD2.n58 2.65567
R423 VDD2.n47 VDD2.n46 1.93989
R424 VDD2.n16 VDD2.n15 1.93989
R425 VDD2.n43 VDD2.n37 1.16414
R426 VDD2.n12 VDD2.n6 1.16414
R427 VDD2 VDD2.n60 0.722483
R428 VDD2.n30 VDD2.n28 0.608947
R429 VDD2.n42 VDD2.n39 0.388379
R430 VDD2.n11 VDD2.n8 0.388379
R431 VDD2.n56 VDD2.n32 0.155672
R432 VDD2.n49 VDD2.n32 0.155672
R433 VDD2.n49 VDD2.n48 0.155672
R434 VDD2.n48 VDD2.n36 0.155672
R435 VDD2.n41 VDD2.n36 0.155672
R436 VDD2.n10 VDD2.n5 0.155672
R437 VDD2.n17 VDD2.n5 0.155672
R438 VDD2.n18 VDD2.n17 0.155672
R439 VDD2.n18 VDD2.n1 0.155672
R440 VDD2.n25 VDD2.n1 0.155672
R441 VP.n27 VP.n26 161.3
R442 VP.n28 VP.n23 161.3
R443 VP.n30 VP.n29 161.3
R444 VP.n31 VP.n22 161.3
R445 VP.n33 VP.n32 161.3
R446 VP.n34 VP.n21 161.3
R447 VP.n36 VP.n35 161.3
R448 VP.n37 VP.n20 161.3
R449 VP.n39 VP.n38 161.3
R450 VP.n40 VP.n19 161.3
R451 VP.n42 VP.n41 161.3
R452 VP.n43 VP.n18 161.3
R453 VP.n45 VP.n44 161.3
R454 VP.n47 VP.n46 161.3
R455 VP.n48 VP.n16 161.3
R456 VP.n50 VP.n49 161.3
R457 VP.n51 VP.n15 161.3
R458 VP.n53 VP.n52 161.3
R459 VP.n54 VP.n14 161.3
R460 VP.n96 VP.n0 161.3
R461 VP.n95 VP.n94 161.3
R462 VP.n93 VP.n1 161.3
R463 VP.n92 VP.n91 161.3
R464 VP.n90 VP.n2 161.3
R465 VP.n89 VP.n88 161.3
R466 VP.n87 VP.n86 161.3
R467 VP.n85 VP.n4 161.3
R468 VP.n84 VP.n83 161.3
R469 VP.n82 VP.n5 161.3
R470 VP.n81 VP.n80 161.3
R471 VP.n79 VP.n6 161.3
R472 VP.n78 VP.n77 161.3
R473 VP.n76 VP.n7 161.3
R474 VP.n75 VP.n74 161.3
R475 VP.n73 VP.n8 161.3
R476 VP.n72 VP.n71 161.3
R477 VP.n70 VP.n9 161.3
R478 VP.n69 VP.n68 161.3
R479 VP.n66 VP.n10 161.3
R480 VP.n65 VP.n64 161.3
R481 VP.n63 VP.n11 161.3
R482 VP.n62 VP.n61 161.3
R483 VP.n60 VP.n12 161.3
R484 VP.n59 VP.n58 161.3
R485 VP.n57 VP.n13 102.927
R486 VP.n98 VP.n97 102.927
R487 VP.n56 VP.n55 102.927
R488 VP.n24 VP.t4 78.9128
R489 VP.n25 VP.n24 68.8984
R490 VP.n61 VP.n11 52.1486
R491 VP.n91 VP.n1 52.1486
R492 VP.n49 VP.n15 52.1486
R493 VP.n57 VP.n56 48.8405
R494 VP.n78 VP.t5 46.0096
R495 VP.n13 VP.t2 46.0096
R496 VP.n67 VP.t8 46.0096
R497 VP.n3 VP.t6 46.0096
R498 VP.n97 VP.t0 46.0096
R499 VP.n36 VP.t7 46.0096
R500 VP.n55 VP.t1 46.0096
R501 VP.n17 VP.t3 46.0096
R502 VP.n25 VP.t9 46.0096
R503 VP.n73 VP.n72 44.3785
R504 VP.n84 VP.n5 44.3785
R505 VP.n42 VP.n19 44.3785
R506 VP.n31 VP.n30 44.3785
R507 VP.n74 VP.n73 36.6083
R508 VP.n80 VP.n5 36.6083
R509 VP.n38 VP.n19 36.6083
R510 VP.n32 VP.n31 36.6083
R511 VP.n65 VP.n11 28.8382
R512 VP.n91 VP.n90 28.8382
R513 VP.n49 VP.n48 28.8382
R514 VP.n60 VP.n59 24.4675
R515 VP.n61 VP.n60 24.4675
R516 VP.n66 VP.n65 24.4675
R517 VP.n68 VP.n9 24.4675
R518 VP.n72 VP.n9 24.4675
R519 VP.n74 VP.n7 24.4675
R520 VP.n78 VP.n7 24.4675
R521 VP.n79 VP.n78 24.4675
R522 VP.n80 VP.n79 24.4675
R523 VP.n85 VP.n84 24.4675
R524 VP.n86 VP.n85 24.4675
R525 VP.n90 VP.n89 24.4675
R526 VP.n95 VP.n1 24.4675
R527 VP.n96 VP.n95 24.4675
R528 VP.n53 VP.n15 24.4675
R529 VP.n54 VP.n53 24.4675
R530 VP.n43 VP.n42 24.4675
R531 VP.n44 VP.n43 24.4675
R532 VP.n48 VP.n47 24.4675
R533 VP.n32 VP.n21 24.4675
R534 VP.n36 VP.n21 24.4675
R535 VP.n37 VP.n36 24.4675
R536 VP.n38 VP.n37 24.4675
R537 VP.n26 VP.n23 24.4675
R538 VP.n30 VP.n23 24.4675
R539 VP.n67 VP.n66 20.5528
R540 VP.n89 VP.n3 20.5528
R541 VP.n47 VP.n17 20.5528
R542 VP.n59 VP.n13 7.82994
R543 VP.n97 VP.n96 7.82994
R544 VP.n55 VP.n54 7.82994
R545 VP.n27 VP.n24 6.98708
R546 VP.n68 VP.n67 3.91522
R547 VP.n86 VP.n3 3.91522
R548 VP.n44 VP.n17 3.91522
R549 VP.n26 VP.n25 3.91522
R550 VP.n56 VP.n14 0.278367
R551 VP.n58 VP.n57 0.278367
R552 VP.n98 VP.n0 0.278367
R553 VP.n28 VP.n27 0.189894
R554 VP.n29 VP.n28 0.189894
R555 VP.n29 VP.n22 0.189894
R556 VP.n33 VP.n22 0.189894
R557 VP.n34 VP.n33 0.189894
R558 VP.n35 VP.n34 0.189894
R559 VP.n35 VP.n20 0.189894
R560 VP.n39 VP.n20 0.189894
R561 VP.n40 VP.n39 0.189894
R562 VP.n41 VP.n40 0.189894
R563 VP.n41 VP.n18 0.189894
R564 VP.n45 VP.n18 0.189894
R565 VP.n46 VP.n45 0.189894
R566 VP.n46 VP.n16 0.189894
R567 VP.n50 VP.n16 0.189894
R568 VP.n51 VP.n50 0.189894
R569 VP.n52 VP.n51 0.189894
R570 VP.n52 VP.n14 0.189894
R571 VP.n58 VP.n12 0.189894
R572 VP.n62 VP.n12 0.189894
R573 VP.n63 VP.n62 0.189894
R574 VP.n64 VP.n63 0.189894
R575 VP.n64 VP.n10 0.189894
R576 VP.n69 VP.n10 0.189894
R577 VP.n70 VP.n69 0.189894
R578 VP.n71 VP.n70 0.189894
R579 VP.n71 VP.n8 0.189894
R580 VP.n75 VP.n8 0.189894
R581 VP.n76 VP.n75 0.189894
R582 VP.n77 VP.n76 0.189894
R583 VP.n77 VP.n6 0.189894
R584 VP.n81 VP.n6 0.189894
R585 VP.n82 VP.n81 0.189894
R586 VP.n83 VP.n82 0.189894
R587 VP.n83 VP.n4 0.189894
R588 VP.n87 VP.n4 0.189894
R589 VP.n88 VP.n87 0.189894
R590 VP.n88 VP.n2 0.189894
R591 VP.n92 VP.n2 0.189894
R592 VP.n93 VP.n92 0.189894
R593 VP.n94 VP.n93 0.189894
R594 VP.n94 VP.n0 0.189894
R595 VP VP.n98 0.153454
R596 VDD1.n22 VDD1.n0 756.745
R597 VDD1.n51 VDD1.n29 756.745
R598 VDD1.n23 VDD1.n22 585
R599 VDD1.n21 VDD1.n20 585
R600 VDD1.n4 VDD1.n3 585
R601 VDD1.n15 VDD1.n14 585
R602 VDD1.n13 VDD1.n12 585
R603 VDD1.n8 VDD1.n7 585
R604 VDD1.n37 VDD1.n36 585
R605 VDD1.n42 VDD1.n41 585
R606 VDD1.n44 VDD1.n43 585
R607 VDD1.n33 VDD1.n32 585
R608 VDD1.n50 VDD1.n49 585
R609 VDD1.n52 VDD1.n51 585
R610 VDD1.n9 VDD1.t5 327.856
R611 VDD1.n38 VDD1.t7 327.856
R612 VDD1.n22 VDD1.n21 171.744
R613 VDD1.n21 VDD1.n3 171.744
R614 VDD1.n14 VDD1.n3 171.744
R615 VDD1.n14 VDD1.n13 171.744
R616 VDD1.n13 VDD1.n7 171.744
R617 VDD1.n42 VDD1.n36 171.744
R618 VDD1.n43 VDD1.n42 171.744
R619 VDD1.n43 VDD1.n32 171.744
R620 VDD1.n50 VDD1.n32 171.744
R621 VDD1.n51 VDD1.n50 171.744
R622 VDD1.n59 VDD1.n58 98.685
R623 VDD1.n28 VDD1.n27 96.7491
R624 VDD1.n57 VDD1.n56 96.749
R625 VDD1.n61 VDD1.n60 96.7489
R626 VDD1.t5 VDD1.n7 85.8723
R627 VDD1.t7 VDD1.n36 85.8723
R628 VDD1.n28 VDD1.n26 50.9375
R629 VDD1.n57 VDD1.n55 50.9375
R630 VDD1.n61 VDD1.n59 42.7638
R631 VDD1.n9 VDD1.n8 16.381
R632 VDD1.n38 VDD1.n37 16.381
R633 VDD1.n12 VDD1.n11 12.8005
R634 VDD1.n41 VDD1.n40 12.8005
R635 VDD1.n15 VDD1.n6 12.0247
R636 VDD1.n44 VDD1.n35 12.0247
R637 VDD1.n16 VDD1.n4 11.249
R638 VDD1.n45 VDD1.n33 11.249
R639 VDD1.n20 VDD1.n19 10.4732
R640 VDD1.n49 VDD1.n48 10.4732
R641 VDD1.n23 VDD1.n2 9.69747
R642 VDD1.n52 VDD1.n31 9.69747
R643 VDD1.n26 VDD1.n25 9.45567
R644 VDD1.n55 VDD1.n54 9.45567
R645 VDD1.n25 VDD1.n24 9.3005
R646 VDD1.n2 VDD1.n1 9.3005
R647 VDD1.n19 VDD1.n18 9.3005
R648 VDD1.n17 VDD1.n16 9.3005
R649 VDD1.n6 VDD1.n5 9.3005
R650 VDD1.n11 VDD1.n10 9.3005
R651 VDD1.n54 VDD1.n53 9.3005
R652 VDD1.n31 VDD1.n30 9.3005
R653 VDD1.n48 VDD1.n47 9.3005
R654 VDD1.n46 VDD1.n45 9.3005
R655 VDD1.n35 VDD1.n34 9.3005
R656 VDD1.n40 VDD1.n39 9.3005
R657 VDD1.n24 VDD1.n0 8.92171
R658 VDD1.n53 VDD1.n29 8.92171
R659 VDD1.n60 VDD1.t6 6.19193
R660 VDD1.n60 VDD1.t8 6.19193
R661 VDD1.n27 VDD1.t0 6.19193
R662 VDD1.n27 VDD1.t2 6.19193
R663 VDD1.n58 VDD1.t3 6.19193
R664 VDD1.n58 VDD1.t9 6.19193
R665 VDD1.n56 VDD1.t1 6.19193
R666 VDD1.n56 VDD1.t4 6.19193
R667 VDD1.n26 VDD1.n0 5.04292
R668 VDD1.n55 VDD1.n29 5.04292
R669 VDD1.n24 VDD1.n23 4.26717
R670 VDD1.n53 VDD1.n52 4.26717
R671 VDD1.n10 VDD1.n9 3.71853
R672 VDD1.n39 VDD1.n38 3.71853
R673 VDD1.n20 VDD1.n2 3.49141
R674 VDD1.n49 VDD1.n31 3.49141
R675 VDD1.n19 VDD1.n4 2.71565
R676 VDD1.n48 VDD1.n33 2.71565
R677 VDD1.n16 VDD1.n15 1.93989
R678 VDD1.n45 VDD1.n44 1.93989
R679 VDD1 VDD1.n61 1.93369
R680 VDD1.n12 VDD1.n6 1.16414
R681 VDD1.n41 VDD1.n35 1.16414
R682 VDD1 VDD1.n28 0.722483
R683 VDD1.n59 VDD1.n57 0.608947
R684 VDD1.n11 VDD1.n8 0.388379
R685 VDD1.n40 VDD1.n37 0.388379
R686 VDD1.n25 VDD1.n1 0.155672
R687 VDD1.n18 VDD1.n1 0.155672
R688 VDD1.n18 VDD1.n17 0.155672
R689 VDD1.n17 VDD1.n5 0.155672
R690 VDD1.n10 VDD1.n5 0.155672
R691 VDD1.n39 VDD1.n34 0.155672
R692 VDD1.n46 VDD1.n34 0.155672
R693 VDD1.n47 VDD1.n46 0.155672
R694 VDD1.n47 VDD1.n30 0.155672
R695 VDD1.n54 VDD1.n30 0.155672
R696 B.n360 B.n127 585
R697 B.n359 B.n358 585
R698 B.n357 B.n128 585
R699 B.n356 B.n355 585
R700 B.n354 B.n129 585
R701 B.n353 B.n352 585
R702 B.n351 B.n130 585
R703 B.n350 B.n349 585
R704 B.n348 B.n131 585
R705 B.n347 B.n346 585
R706 B.n345 B.n132 585
R707 B.n344 B.n343 585
R708 B.n342 B.n133 585
R709 B.n341 B.n340 585
R710 B.n339 B.n134 585
R711 B.n338 B.n337 585
R712 B.n336 B.n135 585
R713 B.n335 B.n334 585
R714 B.n333 B.n136 585
R715 B.n332 B.n331 585
R716 B.n330 B.n137 585
R717 B.n329 B.n328 585
R718 B.n327 B.n326 585
R719 B.n325 B.n141 585
R720 B.n324 B.n323 585
R721 B.n322 B.n142 585
R722 B.n321 B.n320 585
R723 B.n319 B.n143 585
R724 B.n318 B.n317 585
R725 B.n316 B.n144 585
R726 B.n315 B.n314 585
R727 B.n312 B.n145 585
R728 B.n311 B.n310 585
R729 B.n309 B.n148 585
R730 B.n308 B.n307 585
R731 B.n306 B.n149 585
R732 B.n305 B.n304 585
R733 B.n303 B.n150 585
R734 B.n302 B.n301 585
R735 B.n300 B.n151 585
R736 B.n299 B.n298 585
R737 B.n297 B.n152 585
R738 B.n296 B.n295 585
R739 B.n294 B.n153 585
R740 B.n293 B.n292 585
R741 B.n291 B.n154 585
R742 B.n290 B.n289 585
R743 B.n288 B.n155 585
R744 B.n287 B.n286 585
R745 B.n285 B.n156 585
R746 B.n284 B.n283 585
R747 B.n282 B.n157 585
R748 B.n281 B.n280 585
R749 B.n362 B.n361 585
R750 B.n363 B.n126 585
R751 B.n365 B.n364 585
R752 B.n366 B.n125 585
R753 B.n368 B.n367 585
R754 B.n369 B.n124 585
R755 B.n371 B.n370 585
R756 B.n372 B.n123 585
R757 B.n374 B.n373 585
R758 B.n375 B.n122 585
R759 B.n377 B.n376 585
R760 B.n378 B.n121 585
R761 B.n380 B.n379 585
R762 B.n381 B.n120 585
R763 B.n383 B.n382 585
R764 B.n384 B.n119 585
R765 B.n386 B.n385 585
R766 B.n387 B.n118 585
R767 B.n389 B.n388 585
R768 B.n390 B.n117 585
R769 B.n392 B.n391 585
R770 B.n393 B.n116 585
R771 B.n395 B.n394 585
R772 B.n396 B.n115 585
R773 B.n398 B.n397 585
R774 B.n399 B.n114 585
R775 B.n401 B.n400 585
R776 B.n402 B.n113 585
R777 B.n404 B.n403 585
R778 B.n405 B.n112 585
R779 B.n407 B.n406 585
R780 B.n408 B.n111 585
R781 B.n410 B.n409 585
R782 B.n411 B.n110 585
R783 B.n413 B.n412 585
R784 B.n414 B.n109 585
R785 B.n416 B.n415 585
R786 B.n417 B.n108 585
R787 B.n419 B.n418 585
R788 B.n420 B.n107 585
R789 B.n422 B.n421 585
R790 B.n423 B.n106 585
R791 B.n425 B.n424 585
R792 B.n426 B.n105 585
R793 B.n428 B.n427 585
R794 B.n429 B.n104 585
R795 B.n431 B.n430 585
R796 B.n432 B.n103 585
R797 B.n434 B.n433 585
R798 B.n435 B.n102 585
R799 B.n437 B.n436 585
R800 B.n438 B.n101 585
R801 B.n440 B.n439 585
R802 B.n441 B.n100 585
R803 B.n443 B.n442 585
R804 B.n444 B.n99 585
R805 B.n446 B.n445 585
R806 B.n447 B.n98 585
R807 B.n449 B.n448 585
R808 B.n450 B.n97 585
R809 B.n452 B.n451 585
R810 B.n453 B.n96 585
R811 B.n455 B.n454 585
R812 B.n456 B.n95 585
R813 B.n458 B.n457 585
R814 B.n459 B.n94 585
R815 B.n461 B.n460 585
R816 B.n462 B.n93 585
R817 B.n464 B.n463 585
R818 B.n465 B.n92 585
R819 B.n467 B.n466 585
R820 B.n468 B.n91 585
R821 B.n470 B.n469 585
R822 B.n471 B.n90 585
R823 B.n473 B.n472 585
R824 B.n474 B.n89 585
R825 B.n476 B.n475 585
R826 B.n477 B.n88 585
R827 B.n479 B.n478 585
R828 B.n480 B.n87 585
R829 B.n482 B.n481 585
R830 B.n483 B.n86 585
R831 B.n485 B.n484 585
R832 B.n486 B.n85 585
R833 B.n488 B.n487 585
R834 B.n489 B.n84 585
R835 B.n491 B.n490 585
R836 B.n492 B.n83 585
R837 B.n494 B.n493 585
R838 B.n495 B.n82 585
R839 B.n497 B.n496 585
R840 B.n498 B.n81 585
R841 B.n500 B.n499 585
R842 B.n501 B.n80 585
R843 B.n503 B.n502 585
R844 B.n504 B.n79 585
R845 B.n506 B.n505 585
R846 B.n507 B.n78 585
R847 B.n509 B.n508 585
R848 B.n510 B.n77 585
R849 B.n512 B.n511 585
R850 B.n513 B.n76 585
R851 B.n515 B.n514 585
R852 B.n516 B.n75 585
R853 B.n518 B.n517 585
R854 B.n519 B.n74 585
R855 B.n521 B.n520 585
R856 B.n522 B.n73 585
R857 B.n524 B.n523 585
R858 B.n525 B.n72 585
R859 B.n527 B.n526 585
R860 B.n528 B.n71 585
R861 B.n530 B.n529 585
R862 B.n531 B.n70 585
R863 B.n533 B.n532 585
R864 B.n534 B.n69 585
R865 B.n536 B.n535 585
R866 B.n537 B.n68 585
R867 B.n539 B.n538 585
R868 B.n540 B.n67 585
R869 B.n542 B.n541 585
R870 B.n543 B.n66 585
R871 B.n545 B.n544 585
R872 B.n546 B.n65 585
R873 B.n548 B.n547 585
R874 B.n549 B.n64 585
R875 B.n630 B.n33 585
R876 B.n629 B.n628 585
R877 B.n627 B.n34 585
R878 B.n626 B.n625 585
R879 B.n624 B.n35 585
R880 B.n623 B.n622 585
R881 B.n621 B.n36 585
R882 B.n620 B.n619 585
R883 B.n618 B.n37 585
R884 B.n617 B.n616 585
R885 B.n615 B.n38 585
R886 B.n614 B.n613 585
R887 B.n612 B.n39 585
R888 B.n611 B.n610 585
R889 B.n609 B.n40 585
R890 B.n608 B.n607 585
R891 B.n606 B.n41 585
R892 B.n605 B.n604 585
R893 B.n603 B.n42 585
R894 B.n602 B.n601 585
R895 B.n600 B.n43 585
R896 B.n599 B.n598 585
R897 B.n597 B.n596 585
R898 B.n595 B.n47 585
R899 B.n594 B.n593 585
R900 B.n592 B.n48 585
R901 B.n591 B.n590 585
R902 B.n589 B.n49 585
R903 B.n588 B.n587 585
R904 B.n586 B.n50 585
R905 B.n585 B.n584 585
R906 B.n582 B.n51 585
R907 B.n581 B.n580 585
R908 B.n579 B.n54 585
R909 B.n578 B.n577 585
R910 B.n576 B.n55 585
R911 B.n575 B.n574 585
R912 B.n573 B.n56 585
R913 B.n572 B.n571 585
R914 B.n570 B.n57 585
R915 B.n569 B.n568 585
R916 B.n567 B.n58 585
R917 B.n566 B.n565 585
R918 B.n564 B.n59 585
R919 B.n563 B.n562 585
R920 B.n561 B.n60 585
R921 B.n560 B.n559 585
R922 B.n558 B.n61 585
R923 B.n557 B.n556 585
R924 B.n555 B.n62 585
R925 B.n554 B.n553 585
R926 B.n552 B.n63 585
R927 B.n551 B.n550 585
R928 B.n632 B.n631 585
R929 B.n633 B.n32 585
R930 B.n635 B.n634 585
R931 B.n636 B.n31 585
R932 B.n638 B.n637 585
R933 B.n639 B.n30 585
R934 B.n641 B.n640 585
R935 B.n642 B.n29 585
R936 B.n644 B.n643 585
R937 B.n645 B.n28 585
R938 B.n647 B.n646 585
R939 B.n648 B.n27 585
R940 B.n650 B.n649 585
R941 B.n651 B.n26 585
R942 B.n653 B.n652 585
R943 B.n654 B.n25 585
R944 B.n656 B.n655 585
R945 B.n657 B.n24 585
R946 B.n659 B.n658 585
R947 B.n660 B.n23 585
R948 B.n662 B.n661 585
R949 B.n663 B.n22 585
R950 B.n665 B.n664 585
R951 B.n666 B.n21 585
R952 B.n668 B.n667 585
R953 B.n669 B.n20 585
R954 B.n671 B.n670 585
R955 B.n672 B.n19 585
R956 B.n674 B.n673 585
R957 B.n675 B.n18 585
R958 B.n677 B.n676 585
R959 B.n678 B.n17 585
R960 B.n680 B.n679 585
R961 B.n681 B.n16 585
R962 B.n683 B.n682 585
R963 B.n684 B.n15 585
R964 B.n686 B.n685 585
R965 B.n687 B.n14 585
R966 B.n689 B.n688 585
R967 B.n690 B.n13 585
R968 B.n692 B.n691 585
R969 B.n693 B.n12 585
R970 B.n695 B.n694 585
R971 B.n696 B.n11 585
R972 B.n698 B.n697 585
R973 B.n699 B.n10 585
R974 B.n701 B.n700 585
R975 B.n702 B.n9 585
R976 B.n704 B.n703 585
R977 B.n705 B.n8 585
R978 B.n707 B.n706 585
R979 B.n708 B.n7 585
R980 B.n710 B.n709 585
R981 B.n711 B.n6 585
R982 B.n713 B.n712 585
R983 B.n714 B.n5 585
R984 B.n716 B.n715 585
R985 B.n717 B.n4 585
R986 B.n719 B.n718 585
R987 B.n720 B.n3 585
R988 B.n722 B.n721 585
R989 B.n723 B.n0 585
R990 B.n2 B.n1 585
R991 B.n189 B.n188 585
R992 B.n191 B.n190 585
R993 B.n192 B.n187 585
R994 B.n194 B.n193 585
R995 B.n195 B.n186 585
R996 B.n197 B.n196 585
R997 B.n198 B.n185 585
R998 B.n200 B.n199 585
R999 B.n201 B.n184 585
R1000 B.n203 B.n202 585
R1001 B.n204 B.n183 585
R1002 B.n206 B.n205 585
R1003 B.n207 B.n182 585
R1004 B.n209 B.n208 585
R1005 B.n210 B.n181 585
R1006 B.n212 B.n211 585
R1007 B.n213 B.n180 585
R1008 B.n215 B.n214 585
R1009 B.n216 B.n179 585
R1010 B.n218 B.n217 585
R1011 B.n219 B.n178 585
R1012 B.n221 B.n220 585
R1013 B.n222 B.n177 585
R1014 B.n224 B.n223 585
R1015 B.n225 B.n176 585
R1016 B.n227 B.n226 585
R1017 B.n228 B.n175 585
R1018 B.n230 B.n229 585
R1019 B.n231 B.n174 585
R1020 B.n233 B.n232 585
R1021 B.n234 B.n173 585
R1022 B.n236 B.n235 585
R1023 B.n237 B.n172 585
R1024 B.n239 B.n238 585
R1025 B.n240 B.n171 585
R1026 B.n242 B.n241 585
R1027 B.n243 B.n170 585
R1028 B.n245 B.n244 585
R1029 B.n246 B.n169 585
R1030 B.n248 B.n247 585
R1031 B.n249 B.n168 585
R1032 B.n251 B.n250 585
R1033 B.n252 B.n167 585
R1034 B.n254 B.n253 585
R1035 B.n255 B.n166 585
R1036 B.n257 B.n256 585
R1037 B.n258 B.n165 585
R1038 B.n260 B.n259 585
R1039 B.n261 B.n164 585
R1040 B.n263 B.n262 585
R1041 B.n264 B.n163 585
R1042 B.n266 B.n265 585
R1043 B.n267 B.n162 585
R1044 B.n269 B.n268 585
R1045 B.n270 B.n161 585
R1046 B.n272 B.n271 585
R1047 B.n273 B.n160 585
R1048 B.n275 B.n274 585
R1049 B.n276 B.n159 585
R1050 B.n278 B.n277 585
R1051 B.n279 B.n158 585
R1052 B.n280 B.n279 502.111
R1053 B.n362 B.n127 502.111
R1054 B.n550 B.n549 502.111
R1055 B.n632 B.n33 502.111
R1056 B.n138 B.t7 314.8
R1057 B.n52 B.t11 314.8
R1058 B.n146 B.t4 314.8
R1059 B.n44 B.t2 314.8
R1060 B.n725 B.n724 256.663
R1061 B.n139 B.t8 255.066
R1062 B.n53 B.t10 255.066
R1063 B.n147 B.t5 255.066
R1064 B.n45 B.t1 255.066
R1065 B.n146 B.t3 254.272
R1066 B.n138 B.t6 254.272
R1067 B.n52 B.t9 254.272
R1068 B.n44 B.t0 254.272
R1069 B.n724 B.n723 235.042
R1070 B.n724 B.n2 235.042
R1071 B.n280 B.n157 163.367
R1072 B.n284 B.n157 163.367
R1073 B.n285 B.n284 163.367
R1074 B.n286 B.n285 163.367
R1075 B.n286 B.n155 163.367
R1076 B.n290 B.n155 163.367
R1077 B.n291 B.n290 163.367
R1078 B.n292 B.n291 163.367
R1079 B.n292 B.n153 163.367
R1080 B.n296 B.n153 163.367
R1081 B.n297 B.n296 163.367
R1082 B.n298 B.n297 163.367
R1083 B.n298 B.n151 163.367
R1084 B.n302 B.n151 163.367
R1085 B.n303 B.n302 163.367
R1086 B.n304 B.n303 163.367
R1087 B.n304 B.n149 163.367
R1088 B.n308 B.n149 163.367
R1089 B.n309 B.n308 163.367
R1090 B.n310 B.n309 163.367
R1091 B.n310 B.n145 163.367
R1092 B.n315 B.n145 163.367
R1093 B.n316 B.n315 163.367
R1094 B.n317 B.n316 163.367
R1095 B.n317 B.n143 163.367
R1096 B.n321 B.n143 163.367
R1097 B.n322 B.n321 163.367
R1098 B.n323 B.n322 163.367
R1099 B.n323 B.n141 163.367
R1100 B.n327 B.n141 163.367
R1101 B.n328 B.n327 163.367
R1102 B.n328 B.n137 163.367
R1103 B.n332 B.n137 163.367
R1104 B.n333 B.n332 163.367
R1105 B.n334 B.n333 163.367
R1106 B.n334 B.n135 163.367
R1107 B.n338 B.n135 163.367
R1108 B.n339 B.n338 163.367
R1109 B.n340 B.n339 163.367
R1110 B.n340 B.n133 163.367
R1111 B.n344 B.n133 163.367
R1112 B.n345 B.n344 163.367
R1113 B.n346 B.n345 163.367
R1114 B.n346 B.n131 163.367
R1115 B.n350 B.n131 163.367
R1116 B.n351 B.n350 163.367
R1117 B.n352 B.n351 163.367
R1118 B.n352 B.n129 163.367
R1119 B.n356 B.n129 163.367
R1120 B.n357 B.n356 163.367
R1121 B.n358 B.n357 163.367
R1122 B.n358 B.n127 163.367
R1123 B.n549 B.n548 163.367
R1124 B.n548 B.n65 163.367
R1125 B.n544 B.n65 163.367
R1126 B.n544 B.n543 163.367
R1127 B.n543 B.n542 163.367
R1128 B.n542 B.n67 163.367
R1129 B.n538 B.n67 163.367
R1130 B.n538 B.n537 163.367
R1131 B.n537 B.n536 163.367
R1132 B.n536 B.n69 163.367
R1133 B.n532 B.n69 163.367
R1134 B.n532 B.n531 163.367
R1135 B.n531 B.n530 163.367
R1136 B.n530 B.n71 163.367
R1137 B.n526 B.n71 163.367
R1138 B.n526 B.n525 163.367
R1139 B.n525 B.n524 163.367
R1140 B.n524 B.n73 163.367
R1141 B.n520 B.n73 163.367
R1142 B.n520 B.n519 163.367
R1143 B.n519 B.n518 163.367
R1144 B.n518 B.n75 163.367
R1145 B.n514 B.n75 163.367
R1146 B.n514 B.n513 163.367
R1147 B.n513 B.n512 163.367
R1148 B.n512 B.n77 163.367
R1149 B.n508 B.n77 163.367
R1150 B.n508 B.n507 163.367
R1151 B.n507 B.n506 163.367
R1152 B.n506 B.n79 163.367
R1153 B.n502 B.n79 163.367
R1154 B.n502 B.n501 163.367
R1155 B.n501 B.n500 163.367
R1156 B.n500 B.n81 163.367
R1157 B.n496 B.n81 163.367
R1158 B.n496 B.n495 163.367
R1159 B.n495 B.n494 163.367
R1160 B.n494 B.n83 163.367
R1161 B.n490 B.n83 163.367
R1162 B.n490 B.n489 163.367
R1163 B.n489 B.n488 163.367
R1164 B.n488 B.n85 163.367
R1165 B.n484 B.n85 163.367
R1166 B.n484 B.n483 163.367
R1167 B.n483 B.n482 163.367
R1168 B.n482 B.n87 163.367
R1169 B.n478 B.n87 163.367
R1170 B.n478 B.n477 163.367
R1171 B.n477 B.n476 163.367
R1172 B.n476 B.n89 163.367
R1173 B.n472 B.n89 163.367
R1174 B.n472 B.n471 163.367
R1175 B.n471 B.n470 163.367
R1176 B.n470 B.n91 163.367
R1177 B.n466 B.n91 163.367
R1178 B.n466 B.n465 163.367
R1179 B.n465 B.n464 163.367
R1180 B.n464 B.n93 163.367
R1181 B.n460 B.n93 163.367
R1182 B.n460 B.n459 163.367
R1183 B.n459 B.n458 163.367
R1184 B.n458 B.n95 163.367
R1185 B.n454 B.n95 163.367
R1186 B.n454 B.n453 163.367
R1187 B.n453 B.n452 163.367
R1188 B.n452 B.n97 163.367
R1189 B.n448 B.n97 163.367
R1190 B.n448 B.n447 163.367
R1191 B.n447 B.n446 163.367
R1192 B.n446 B.n99 163.367
R1193 B.n442 B.n99 163.367
R1194 B.n442 B.n441 163.367
R1195 B.n441 B.n440 163.367
R1196 B.n440 B.n101 163.367
R1197 B.n436 B.n101 163.367
R1198 B.n436 B.n435 163.367
R1199 B.n435 B.n434 163.367
R1200 B.n434 B.n103 163.367
R1201 B.n430 B.n103 163.367
R1202 B.n430 B.n429 163.367
R1203 B.n429 B.n428 163.367
R1204 B.n428 B.n105 163.367
R1205 B.n424 B.n105 163.367
R1206 B.n424 B.n423 163.367
R1207 B.n423 B.n422 163.367
R1208 B.n422 B.n107 163.367
R1209 B.n418 B.n107 163.367
R1210 B.n418 B.n417 163.367
R1211 B.n417 B.n416 163.367
R1212 B.n416 B.n109 163.367
R1213 B.n412 B.n109 163.367
R1214 B.n412 B.n411 163.367
R1215 B.n411 B.n410 163.367
R1216 B.n410 B.n111 163.367
R1217 B.n406 B.n111 163.367
R1218 B.n406 B.n405 163.367
R1219 B.n405 B.n404 163.367
R1220 B.n404 B.n113 163.367
R1221 B.n400 B.n113 163.367
R1222 B.n400 B.n399 163.367
R1223 B.n399 B.n398 163.367
R1224 B.n398 B.n115 163.367
R1225 B.n394 B.n115 163.367
R1226 B.n394 B.n393 163.367
R1227 B.n393 B.n392 163.367
R1228 B.n392 B.n117 163.367
R1229 B.n388 B.n117 163.367
R1230 B.n388 B.n387 163.367
R1231 B.n387 B.n386 163.367
R1232 B.n386 B.n119 163.367
R1233 B.n382 B.n119 163.367
R1234 B.n382 B.n381 163.367
R1235 B.n381 B.n380 163.367
R1236 B.n380 B.n121 163.367
R1237 B.n376 B.n121 163.367
R1238 B.n376 B.n375 163.367
R1239 B.n375 B.n374 163.367
R1240 B.n374 B.n123 163.367
R1241 B.n370 B.n123 163.367
R1242 B.n370 B.n369 163.367
R1243 B.n369 B.n368 163.367
R1244 B.n368 B.n125 163.367
R1245 B.n364 B.n125 163.367
R1246 B.n364 B.n363 163.367
R1247 B.n363 B.n362 163.367
R1248 B.n628 B.n33 163.367
R1249 B.n628 B.n627 163.367
R1250 B.n627 B.n626 163.367
R1251 B.n626 B.n35 163.367
R1252 B.n622 B.n35 163.367
R1253 B.n622 B.n621 163.367
R1254 B.n621 B.n620 163.367
R1255 B.n620 B.n37 163.367
R1256 B.n616 B.n37 163.367
R1257 B.n616 B.n615 163.367
R1258 B.n615 B.n614 163.367
R1259 B.n614 B.n39 163.367
R1260 B.n610 B.n39 163.367
R1261 B.n610 B.n609 163.367
R1262 B.n609 B.n608 163.367
R1263 B.n608 B.n41 163.367
R1264 B.n604 B.n41 163.367
R1265 B.n604 B.n603 163.367
R1266 B.n603 B.n602 163.367
R1267 B.n602 B.n43 163.367
R1268 B.n598 B.n43 163.367
R1269 B.n598 B.n597 163.367
R1270 B.n597 B.n47 163.367
R1271 B.n593 B.n47 163.367
R1272 B.n593 B.n592 163.367
R1273 B.n592 B.n591 163.367
R1274 B.n591 B.n49 163.367
R1275 B.n587 B.n49 163.367
R1276 B.n587 B.n586 163.367
R1277 B.n586 B.n585 163.367
R1278 B.n585 B.n51 163.367
R1279 B.n580 B.n51 163.367
R1280 B.n580 B.n579 163.367
R1281 B.n579 B.n578 163.367
R1282 B.n578 B.n55 163.367
R1283 B.n574 B.n55 163.367
R1284 B.n574 B.n573 163.367
R1285 B.n573 B.n572 163.367
R1286 B.n572 B.n57 163.367
R1287 B.n568 B.n57 163.367
R1288 B.n568 B.n567 163.367
R1289 B.n567 B.n566 163.367
R1290 B.n566 B.n59 163.367
R1291 B.n562 B.n59 163.367
R1292 B.n562 B.n561 163.367
R1293 B.n561 B.n560 163.367
R1294 B.n560 B.n61 163.367
R1295 B.n556 B.n61 163.367
R1296 B.n556 B.n555 163.367
R1297 B.n555 B.n554 163.367
R1298 B.n554 B.n63 163.367
R1299 B.n550 B.n63 163.367
R1300 B.n633 B.n632 163.367
R1301 B.n634 B.n633 163.367
R1302 B.n634 B.n31 163.367
R1303 B.n638 B.n31 163.367
R1304 B.n639 B.n638 163.367
R1305 B.n640 B.n639 163.367
R1306 B.n640 B.n29 163.367
R1307 B.n644 B.n29 163.367
R1308 B.n645 B.n644 163.367
R1309 B.n646 B.n645 163.367
R1310 B.n646 B.n27 163.367
R1311 B.n650 B.n27 163.367
R1312 B.n651 B.n650 163.367
R1313 B.n652 B.n651 163.367
R1314 B.n652 B.n25 163.367
R1315 B.n656 B.n25 163.367
R1316 B.n657 B.n656 163.367
R1317 B.n658 B.n657 163.367
R1318 B.n658 B.n23 163.367
R1319 B.n662 B.n23 163.367
R1320 B.n663 B.n662 163.367
R1321 B.n664 B.n663 163.367
R1322 B.n664 B.n21 163.367
R1323 B.n668 B.n21 163.367
R1324 B.n669 B.n668 163.367
R1325 B.n670 B.n669 163.367
R1326 B.n670 B.n19 163.367
R1327 B.n674 B.n19 163.367
R1328 B.n675 B.n674 163.367
R1329 B.n676 B.n675 163.367
R1330 B.n676 B.n17 163.367
R1331 B.n680 B.n17 163.367
R1332 B.n681 B.n680 163.367
R1333 B.n682 B.n681 163.367
R1334 B.n682 B.n15 163.367
R1335 B.n686 B.n15 163.367
R1336 B.n687 B.n686 163.367
R1337 B.n688 B.n687 163.367
R1338 B.n688 B.n13 163.367
R1339 B.n692 B.n13 163.367
R1340 B.n693 B.n692 163.367
R1341 B.n694 B.n693 163.367
R1342 B.n694 B.n11 163.367
R1343 B.n698 B.n11 163.367
R1344 B.n699 B.n698 163.367
R1345 B.n700 B.n699 163.367
R1346 B.n700 B.n9 163.367
R1347 B.n704 B.n9 163.367
R1348 B.n705 B.n704 163.367
R1349 B.n706 B.n705 163.367
R1350 B.n706 B.n7 163.367
R1351 B.n710 B.n7 163.367
R1352 B.n711 B.n710 163.367
R1353 B.n712 B.n711 163.367
R1354 B.n712 B.n5 163.367
R1355 B.n716 B.n5 163.367
R1356 B.n717 B.n716 163.367
R1357 B.n718 B.n717 163.367
R1358 B.n718 B.n3 163.367
R1359 B.n722 B.n3 163.367
R1360 B.n723 B.n722 163.367
R1361 B.n189 B.n2 163.367
R1362 B.n190 B.n189 163.367
R1363 B.n190 B.n187 163.367
R1364 B.n194 B.n187 163.367
R1365 B.n195 B.n194 163.367
R1366 B.n196 B.n195 163.367
R1367 B.n196 B.n185 163.367
R1368 B.n200 B.n185 163.367
R1369 B.n201 B.n200 163.367
R1370 B.n202 B.n201 163.367
R1371 B.n202 B.n183 163.367
R1372 B.n206 B.n183 163.367
R1373 B.n207 B.n206 163.367
R1374 B.n208 B.n207 163.367
R1375 B.n208 B.n181 163.367
R1376 B.n212 B.n181 163.367
R1377 B.n213 B.n212 163.367
R1378 B.n214 B.n213 163.367
R1379 B.n214 B.n179 163.367
R1380 B.n218 B.n179 163.367
R1381 B.n219 B.n218 163.367
R1382 B.n220 B.n219 163.367
R1383 B.n220 B.n177 163.367
R1384 B.n224 B.n177 163.367
R1385 B.n225 B.n224 163.367
R1386 B.n226 B.n225 163.367
R1387 B.n226 B.n175 163.367
R1388 B.n230 B.n175 163.367
R1389 B.n231 B.n230 163.367
R1390 B.n232 B.n231 163.367
R1391 B.n232 B.n173 163.367
R1392 B.n236 B.n173 163.367
R1393 B.n237 B.n236 163.367
R1394 B.n238 B.n237 163.367
R1395 B.n238 B.n171 163.367
R1396 B.n242 B.n171 163.367
R1397 B.n243 B.n242 163.367
R1398 B.n244 B.n243 163.367
R1399 B.n244 B.n169 163.367
R1400 B.n248 B.n169 163.367
R1401 B.n249 B.n248 163.367
R1402 B.n250 B.n249 163.367
R1403 B.n250 B.n167 163.367
R1404 B.n254 B.n167 163.367
R1405 B.n255 B.n254 163.367
R1406 B.n256 B.n255 163.367
R1407 B.n256 B.n165 163.367
R1408 B.n260 B.n165 163.367
R1409 B.n261 B.n260 163.367
R1410 B.n262 B.n261 163.367
R1411 B.n262 B.n163 163.367
R1412 B.n266 B.n163 163.367
R1413 B.n267 B.n266 163.367
R1414 B.n268 B.n267 163.367
R1415 B.n268 B.n161 163.367
R1416 B.n272 B.n161 163.367
R1417 B.n273 B.n272 163.367
R1418 B.n274 B.n273 163.367
R1419 B.n274 B.n159 163.367
R1420 B.n278 B.n159 163.367
R1421 B.n279 B.n278 163.367
R1422 B.n147 B.n146 59.7338
R1423 B.n139 B.n138 59.7338
R1424 B.n53 B.n52 59.7338
R1425 B.n45 B.n44 59.7338
R1426 B.n313 B.n147 59.5399
R1427 B.n140 B.n139 59.5399
R1428 B.n583 B.n53 59.5399
R1429 B.n46 B.n45 59.5399
R1430 B.n631 B.n630 32.6249
R1431 B.n551 B.n64 32.6249
R1432 B.n361 B.n360 32.6249
R1433 B.n281 B.n158 32.6249
R1434 B B.n725 18.0485
R1435 B.n631 B.n32 10.6151
R1436 B.n635 B.n32 10.6151
R1437 B.n636 B.n635 10.6151
R1438 B.n637 B.n636 10.6151
R1439 B.n637 B.n30 10.6151
R1440 B.n641 B.n30 10.6151
R1441 B.n642 B.n641 10.6151
R1442 B.n643 B.n642 10.6151
R1443 B.n643 B.n28 10.6151
R1444 B.n647 B.n28 10.6151
R1445 B.n648 B.n647 10.6151
R1446 B.n649 B.n648 10.6151
R1447 B.n649 B.n26 10.6151
R1448 B.n653 B.n26 10.6151
R1449 B.n654 B.n653 10.6151
R1450 B.n655 B.n654 10.6151
R1451 B.n655 B.n24 10.6151
R1452 B.n659 B.n24 10.6151
R1453 B.n660 B.n659 10.6151
R1454 B.n661 B.n660 10.6151
R1455 B.n661 B.n22 10.6151
R1456 B.n665 B.n22 10.6151
R1457 B.n666 B.n665 10.6151
R1458 B.n667 B.n666 10.6151
R1459 B.n667 B.n20 10.6151
R1460 B.n671 B.n20 10.6151
R1461 B.n672 B.n671 10.6151
R1462 B.n673 B.n672 10.6151
R1463 B.n673 B.n18 10.6151
R1464 B.n677 B.n18 10.6151
R1465 B.n678 B.n677 10.6151
R1466 B.n679 B.n678 10.6151
R1467 B.n679 B.n16 10.6151
R1468 B.n683 B.n16 10.6151
R1469 B.n684 B.n683 10.6151
R1470 B.n685 B.n684 10.6151
R1471 B.n685 B.n14 10.6151
R1472 B.n689 B.n14 10.6151
R1473 B.n690 B.n689 10.6151
R1474 B.n691 B.n690 10.6151
R1475 B.n691 B.n12 10.6151
R1476 B.n695 B.n12 10.6151
R1477 B.n696 B.n695 10.6151
R1478 B.n697 B.n696 10.6151
R1479 B.n697 B.n10 10.6151
R1480 B.n701 B.n10 10.6151
R1481 B.n702 B.n701 10.6151
R1482 B.n703 B.n702 10.6151
R1483 B.n703 B.n8 10.6151
R1484 B.n707 B.n8 10.6151
R1485 B.n708 B.n707 10.6151
R1486 B.n709 B.n708 10.6151
R1487 B.n709 B.n6 10.6151
R1488 B.n713 B.n6 10.6151
R1489 B.n714 B.n713 10.6151
R1490 B.n715 B.n714 10.6151
R1491 B.n715 B.n4 10.6151
R1492 B.n719 B.n4 10.6151
R1493 B.n720 B.n719 10.6151
R1494 B.n721 B.n720 10.6151
R1495 B.n721 B.n0 10.6151
R1496 B.n630 B.n629 10.6151
R1497 B.n629 B.n34 10.6151
R1498 B.n625 B.n34 10.6151
R1499 B.n625 B.n624 10.6151
R1500 B.n624 B.n623 10.6151
R1501 B.n623 B.n36 10.6151
R1502 B.n619 B.n36 10.6151
R1503 B.n619 B.n618 10.6151
R1504 B.n618 B.n617 10.6151
R1505 B.n617 B.n38 10.6151
R1506 B.n613 B.n38 10.6151
R1507 B.n613 B.n612 10.6151
R1508 B.n612 B.n611 10.6151
R1509 B.n611 B.n40 10.6151
R1510 B.n607 B.n40 10.6151
R1511 B.n607 B.n606 10.6151
R1512 B.n606 B.n605 10.6151
R1513 B.n605 B.n42 10.6151
R1514 B.n601 B.n42 10.6151
R1515 B.n601 B.n600 10.6151
R1516 B.n600 B.n599 10.6151
R1517 B.n596 B.n595 10.6151
R1518 B.n595 B.n594 10.6151
R1519 B.n594 B.n48 10.6151
R1520 B.n590 B.n48 10.6151
R1521 B.n590 B.n589 10.6151
R1522 B.n589 B.n588 10.6151
R1523 B.n588 B.n50 10.6151
R1524 B.n584 B.n50 10.6151
R1525 B.n582 B.n581 10.6151
R1526 B.n581 B.n54 10.6151
R1527 B.n577 B.n54 10.6151
R1528 B.n577 B.n576 10.6151
R1529 B.n576 B.n575 10.6151
R1530 B.n575 B.n56 10.6151
R1531 B.n571 B.n56 10.6151
R1532 B.n571 B.n570 10.6151
R1533 B.n570 B.n569 10.6151
R1534 B.n569 B.n58 10.6151
R1535 B.n565 B.n58 10.6151
R1536 B.n565 B.n564 10.6151
R1537 B.n564 B.n563 10.6151
R1538 B.n563 B.n60 10.6151
R1539 B.n559 B.n60 10.6151
R1540 B.n559 B.n558 10.6151
R1541 B.n558 B.n557 10.6151
R1542 B.n557 B.n62 10.6151
R1543 B.n553 B.n62 10.6151
R1544 B.n553 B.n552 10.6151
R1545 B.n552 B.n551 10.6151
R1546 B.n547 B.n64 10.6151
R1547 B.n547 B.n546 10.6151
R1548 B.n546 B.n545 10.6151
R1549 B.n545 B.n66 10.6151
R1550 B.n541 B.n66 10.6151
R1551 B.n541 B.n540 10.6151
R1552 B.n540 B.n539 10.6151
R1553 B.n539 B.n68 10.6151
R1554 B.n535 B.n68 10.6151
R1555 B.n535 B.n534 10.6151
R1556 B.n534 B.n533 10.6151
R1557 B.n533 B.n70 10.6151
R1558 B.n529 B.n70 10.6151
R1559 B.n529 B.n528 10.6151
R1560 B.n528 B.n527 10.6151
R1561 B.n527 B.n72 10.6151
R1562 B.n523 B.n72 10.6151
R1563 B.n523 B.n522 10.6151
R1564 B.n522 B.n521 10.6151
R1565 B.n521 B.n74 10.6151
R1566 B.n517 B.n74 10.6151
R1567 B.n517 B.n516 10.6151
R1568 B.n516 B.n515 10.6151
R1569 B.n515 B.n76 10.6151
R1570 B.n511 B.n76 10.6151
R1571 B.n511 B.n510 10.6151
R1572 B.n510 B.n509 10.6151
R1573 B.n509 B.n78 10.6151
R1574 B.n505 B.n78 10.6151
R1575 B.n505 B.n504 10.6151
R1576 B.n504 B.n503 10.6151
R1577 B.n503 B.n80 10.6151
R1578 B.n499 B.n80 10.6151
R1579 B.n499 B.n498 10.6151
R1580 B.n498 B.n497 10.6151
R1581 B.n497 B.n82 10.6151
R1582 B.n493 B.n82 10.6151
R1583 B.n493 B.n492 10.6151
R1584 B.n492 B.n491 10.6151
R1585 B.n491 B.n84 10.6151
R1586 B.n487 B.n84 10.6151
R1587 B.n487 B.n486 10.6151
R1588 B.n486 B.n485 10.6151
R1589 B.n485 B.n86 10.6151
R1590 B.n481 B.n86 10.6151
R1591 B.n481 B.n480 10.6151
R1592 B.n480 B.n479 10.6151
R1593 B.n479 B.n88 10.6151
R1594 B.n475 B.n88 10.6151
R1595 B.n475 B.n474 10.6151
R1596 B.n474 B.n473 10.6151
R1597 B.n473 B.n90 10.6151
R1598 B.n469 B.n90 10.6151
R1599 B.n469 B.n468 10.6151
R1600 B.n468 B.n467 10.6151
R1601 B.n467 B.n92 10.6151
R1602 B.n463 B.n92 10.6151
R1603 B.n463 B.n462 10.6151
R1604 B.n462 B.n461 10.6151
R1605 B.n461 B.n94 10.6151
R1606 B.n457 B.n94 10.6151
R1607 B.n457 B.n456 10.6151
R1608 B.n456 B.n455 10.6151
R1609 B.n455 B.n96 10.6151
R1610 B.n451 B.n96 10.6151
R1611 B.n451 B.n450 10.6151
R1612 B.n450 B.n449 10.6151
R1613 B.n449 B.n98 10.6151
R1614 B.n445 B.n98 10.6151
R1615 B.n445 B.n444 10.6151
R1616 B.n444 B.n443 10.6151
R1617 B.n443 B.n100 10.6151
R1618 B.n439 B.n100 10.6151
R1619 B.n439 B.n438 10.6151
R1620 B.n438 B.n437 10.6151
R1621 B.n437 B.n102 10.6151
R1622 B.n433 B.n102 10.6151
R1623 B.n433 B.n432 10.6151
R1624 B.n432 B.n431 10.6151
R1625 B.n431 B.n104 10.6151
R1626 B.n427 B.n104 10.6151
R1627 B.n427 B.n426 10.6151
R1628 B.n426 B.n425 10.6151
R1629 B.n425 B.n106 10.6151
R1630 B.n421 B.n106 10.6151
R1631 B.n421 B.n420 10.6151
R1632 B.n420 B.n419 10.6151
R1633 B.n419 B.n108 10.6151
R1634 B.n415 B.n108 10.6151
R1635 B.n415 B.n414 10.6151
R1636 B.n414 B.n413 10.6151
R1637 B.n413 B.n110 10.6151
R1638 B.n409 B.n110 10.6151
R1639 B.n409 B.n408 10.6151
R1640 B.n408 B.n407 10.6151
R1641 B.n407 B.n112 10.6151
R1642 B.n403 B.n112 10.6151
R1643 B.n403 B.n402 10.6151
R1644 B.n402 B.n401 10.6151
R1645 B.n401 B.n114 10.6151
R1646 B.n397 B.n114 10.6151
R1647 B.n397 B.n396 10.6151
R1648 B.n396 B.n395 10.6151
R1649 B.n395 B.n116 10.6151
R1650 B.n391 B.n116 10.6151
R1651 B.n391 B.n390 10.6151
R1652 B.n390 B.n389 10.6151
R1653 B.n389 B.n118 10.6151
R1654 B.n385 B.n118 10.6151
R1655 B.n385 B.n384 10.6151
R1656 B.n384 B.n383 10.6151
R1657 B.n383 B.n120 10.6151
R1658 B.n379 B.n120 10.6151
R1659 B.n379 B.n378 10.6151
R1660 B.n378 B.n377 10.6151
R1661 B.n377 B.n122 10.6151
R1662 B.n373 B.n122 10.6151
R1663 B.n373 B.n372 10.6151
R1664 B.n372 B.n371 10.6151
R1665 B.n371 B.n124 10.6151
R1666 B.n367 B.n124 10.6151
R1667 B.n367 B.n366 10.6151
R1668 B.n366 B.n365 10.6151
R1669 B.n365 B.n126 10.6151
R1670 B.n361 B.n126 10.6151
R1671 B.n188 B.n1 10.6151
R1672 B.n191 B.n188 10.6151
R1673 B.n192 B.n191 10.6151
R1674 B.n193 B.n192 10.6151
R1675 B.n193 B.n186 10.6151
R1676 B.n197 B.n186 10.6151
R1677 B.n198 B.n197 10.6151
R1678 B.n199 B.n198 10.6151
R1679 B.n199 B.n184 10.6151
R1680 B.n203 B.n184 10.6151
R1681 B.n204 B.n203 10.6151
R1682 B.n205 B.n204 10.6151
R1683 B.n205 B.n182 10.6151
R1684 B.n209 B.n182 10.6151
R1685 B.n210 B.n209 10.6151
R1686 B.n211 B.n210 10.6151
R1687 B.n211 B.n180 10.6151
R1688 B.n215 B.n180 10.6151
R1689 B.n216 B.n215 10.6151
R1690 B.n217 B.n216 10.6151
R1691 B.n217 B.n178 10.6151
R1692 B.n221 B.n178 10.6151
R1693 B.n222 B.n221 10.6151
R1694 B.n223 B.n222 10.6151
R1695 B.n223 B.n176 10.6151
R1696 B.n227 B.n176 10.6151
R1697 B.n228 B.n227 10.6151
R1698 B.n229 B.n228 10.6151
R1699 B.n229 B.n174 10.6151
R1700 B.n233 B.n174 10.6151
R1701 B.n234 B.n233 10.6151
R1702 B.n235 B.n234 10.6151
R1703 B.n235 B.n172 10.6151
R1704 B.n239 B.n172 10.6151
R1705 B.n240 B.n239 10.6151
R1706 B.n241 B.n240 10.6151
R1707 B.n241 B.n170 10.6151
R1708 B.n245 B.n170 10.6151
R1709 B.n246 B.n245 10.6151
R1710 B.n247 B.n246 10.6151
R1711 B.n247 B.n168 10.6151
R1712 B.n251 B.n168 10.6151
R1713 B.n252 B.n251 10.6151
R1714 B.n253 B.n252 10.6151
R1715 B.n253 B.n166 10.6151
R1716 B.n257 B.n166 10.6151
R1717 B.n258 B.n257 10.6151
R1718 B.n259 B.n258 10.6151
R1719 B.n259 B.n164 10.6151
R1720 B.n263 B.n164 10.6151
R1721 B.n264 B.n263 10.6151
R1722 B.n265 B.n264 10.6151
R1723 B.n265 B.n162 10.6151
R1724 B.n269 B.n162 10.6151
R1725 B.n270 B.n269 10.6151
R1726 B.n271 B.n270 10.6151
R1727 B.n271 B.n160 10.6151
R1728 B.n275 B.n160 10.6151
R1729 B.n276 B.n275 10.6151
R1730 B.n277 B.n276 10.6151
R1731 B.n277 B.n158 10.6151
R1732 B.n282 B.n281 10.6151
R1733 B.n283 B.n282 10.6151
R1734 B.n283 B.n156 10.6151
R1735 B.n287 B.n156 10.6151
R1736 B.n288 B.n287 10.6151
R1737 B.n289 B.n288 10.6151
R1738 B.n289 B.n154 10.6151
R1739 B.n293 B.n154 10.6151
R1740 B.n294 B.n293 10.6151
R1741 B.n295 B.n294 10.6151
R1742 B.n295 B.n152 10.6151
R1743 B.n299 B.n152 10.6151
R1744 B.n300 B.n299 10.6151
R1745 B.n301 B.n300 10.6151
R1746 B.n301 B.n150 10.6151
R1747 B.n305 B.n150 10.6151
R1748 B.n306 B.n305 10.6151
R1749 B.n307 B.n306 10.6151
R1750 B.n307 B.n148 10.6151
R1751 B.n311 B.n148 10.6151
R1752 B.n312 B.n311 10.6151
R1753 B.n314 B.n144 10.6151
R1754 B.n318 B.n144 10.6151
R1755 B.n319 B.n318 10.6151
R1756 B.n320 B.n319 10.6151
R1757 B.n320 B.n142 10.6151
R1758 B.n324 B.n142 10.6151
R1759 B.n325 B.n324 10.6151
R1760 B.n326 B.n325 10.6151
R1761 B.n330 B.n329 10.6151
R1762 B.n331 B.n330 10.6151
R1763 B.n331 B.n136 10.6151
R1764 B.n335 B.n136 10.6151
R1765 B.n336 B.n335 10.6151
R1766 B.n337 B.n336 10.6151
R1767 B.n337 B.n134 10.6151
R1768 B.n341 B.n134 10.6151
R1769 B.n342 B.n341 10.6151
R1770 B.n343 B.n342 10.6151
R1771 B.n343 B.n132 10.6151
R1772 B.n347 B.n132 10.6151
R1773 B.n348 B.n347 10.6151
R1774 B.n349 B.n348 10.6151
R1775 B.n349 B.n130 10.6151
R1776 B.n353 B.n130 10.6151
R1777 B.n354 B.n353 10.6151
R1778 B.n355 B.n354 10.6151
R1779 B.n355 B.n128 10.6151
R1780 B.n359 B.n128 10.6151
R1781 B.n360 B.n359 10.6151
R1782 B.n725 B.n0 8.11757
R1783 B.n725 B.n1 8.11757
R1784 B.n596 B.n46 6.5566
R1785 B.n584 B.n583 6.5566
R1786 B.n314 B.n313 6.5566
R1787 B.n326 B.n140 6.5566
R1788 B.n599 B.n46 4.05904
R1789 B.n583 B.n582 4.05904
R1790 B.n313 B.n312 4.05904
R1791 B.n329 B.n140 4.05904
C0 VN B 1.28752f
C1 VP VN 7.36749f
C2 VDD2 VN 5.01754f
C3 VTAIL w_n4666_n2018# 2.28188f
C4 VTAIL VDD1 7.40201f
C5 VTAIL B 2.24587f
C6 VTAIL VP 6.26435f
C7 VDD1 w_n4666_n2018# 2.37531f
C8 VTAIL VDD2 7.4556f
C9 w_n4666_n2018# B 8.920191f
C10 VDD1 B 2.00392f
C11 VP w_n4666_n2018# 10.5198f
C12 VP VDD1 5.46317f
C13 VP B 2.31064f
C14 VDD2 w_n4666_n2018# 2.52639f
C15 VDD2 VDD1 2.27022f
C16 VTAIL VN 6.25017f
C17 VDD2 B 2.12784f
C18 VDD2 VP 0.606238f
C19 w_n4666_n2018# VN 9.91189f
C20 VDD1 VN 0.153546f
C21 VDD2 VSUBS 2.130569f
C22 VDD1 VSUBS 1.864551f
C23 VTAIL VSUBS 0.671884f
C24 VN VSUBS 7.616529f
C25 VP VSUBS 3.871306f
C26 B VSUBS 4.695043f
C27 w_n4666_n2018# VSUBS 0.117863p
C28 B.n0 VSUBS 0.010847f
C29 B.n1 VSUBS 0.010847f
C30 B.n2 VSUBS 0.016042f
C31 B.n3 VSUBS 0.012293f
C32 B.n4 VSUBS 0.012293f
C33 B.n5 VSUBS 0.012293f
C34 B.n6 VSUBS 0.012293f
C35 B.n7 VSUBS 0.012293f
C36 B.n8 VSUBS 0.012293f
C37 B.n9 VSUBS 0.012293f
C38 B.n10 VSUBS 0.012293f
C39 B.n11 VSUBS 0.012293f
C40 B.n12 VSUBS 0.012293f
C41 B.n13 VSUBS 0.012293f
C42 B.n14 VSUBS 0.012293f
C43 B.n15 VSUBS 0.012293f
C44 B.n16 VSUBS 0.012293f
C45 B.n17 VSUBS 0.012293f
C46 B.n18 VSUBS 0.012293f
C47 B.n19 VSUBS 0.012293f
C48 B.n20 VSUBS 0.012293f
C49 B.n21 VSUBS 0.012293f
C50 B.n22 VSUBS 0.012293f
C51 B.n23 VSUBS 0.012293f
C52 B.n24 VSUBS 0.012293f
C53 B.n25 VSUBS 0.012293f
C54 B.n26 VSUBS 0.012293f
C55 B.n27 VSUBS 0.012293f
C56 B.n28 VSUBS 0.012293f
C57 B.n29 VSUBS 0.012293f
C58 B.n30 VSUBS 0.012293f
C59 B.n31 VSUBS 0.012293f
C60 B.n32 VSUBS 0.012293f
C61 B.n33 VSUBS 0.02933f
C62 B.n34 VSUBS 0.012293f
C63 B.n35 VSUBS 0.012293f
C64 B.n36 VSUBS 0.012293f
C65 B.n37 VSUBS 0.012293f
C66 B.n38 VSUBS 0.012293f
C67 B.n39 VSUBS 0.012293f
C68 B.n40 VSUBS 0.012293f
C69 B.n41 VSUBS 0.012293f
C70 B.n42 VSUBS 0.012293f
C71 B.n43 VSUBS 0.012293f
C72 B.t1 VSUBS 0.134681f
C73 B.t2 VSUBS 0.178922f
C74 B.t0 VSUBS 1.20945f
C75 B.n44 VSUBS 0.307089f
C76 B.n45 VSUBS 0.250688f
C77 B.n46 VSUBS 0.028482f
C78 B.n47 VSUBS 0.012293f
C79 B.n48 VSUBS 0.012293f
C80 B.n49 VSUBS 0.012293f
C81 B.n50 VSUBS 0.012293f
C82 B.n51 VSUBS 0.012293f
C83 B.t10 VSUBS 0.134684f
C84 B.t11 VSUBS 0.178925f
C85 B.t9 VSUBS 1.20945f
C86 B.n52 VSUBS 0.307087f
C87 B.n53 VSUBS 0.250685f
C88 B.n54 VSUBS 0.012293f
C89 B.n55 VSUBS 0.012293f
C90 B.n56 VSUBS 0.012293f
C91 B.n57 VSUBS 0.012293f
C92 B.n58 VSUBS 0.012293f
C93 B.n59 VSUBS 0.012293f
C94 B.n60 VSUBS 0.012293f
C95 B.n61 VSUBS 0.012293f
C96 B.n62 VSUBS 0.012293f
C97 B.n63 VSUBS 0.012293f
C98 B.n64 VSUBS 0.02816f
C99 B.n65 VSUBS 0.012293f
C100 B.n66 VSUBS 0.012293f
C101 B.n67 VSUBS 0.012293f
C102 B.n68 VSUBS 0.012293f
C103 B.n69 VSUBS 0.012293f
C104 B.n70 VSUBS 0.012293f
C105 B.n71 VSUBS 0.012293f
C106 B.n72 VSUBS 0.012293f
C107 B.n73 VSUBS 0.012293f
C108 B.n74 VSUBS 0.012293f
C109 B.n75 VSUBS 0.012293f
C110 B.n76 VSUBS 0.012293f
C111 B.n77 VSUBS 0.012293f
C112 B.n78 VSUBS 0.012293f
C113 B.n79 VSUBS 0.012293f
C114 B.n80 VSUBS 0.012293f
C115 B.n81 VSUBS 0.012293f
C116 B.n82 VSUBS 0.012293f
C117 B.n83 VSUBS 0.012293f
C118 B.n84 VSUBS 0.012293f
C119 B.n85 VSUBS 0.012293f
C120 B.n86 VSUBS 0.012293f
C121 B.n87 VSUBS 0.012293f
C122 B.n88 VSUBS 0.012293f
C123 B.n89 VSUBS 0.012293f
C124 B.n90 VSUBS 0.012293f
C125 B.n91 VSUBS 0.012293f
C126 B.n92 VSUBS 0.012293f
C127 B.n93 VSUBS 0.012293f
C128 B.n94 VSUBS 0.012293f
C129 B.n95 VSUBS 0.012293f
C130 B.n96 VSUBS 0.012293f
C131 B.n97 VSUBS 0.012293f
C132 B.n98 VSUBS 0.012293f
C133 B.n99 VSUBS 0.012293f
C134 B.n100 VSUBS 0.012293f
C135 B.n101 VSUBS 0.012293f
C136 B.n102 VSUBS 0.012293f
C137 B.n103 VSUBS 0.012293f
C138 B.n104 VSUBS 0.012293f
C139 B.n105 VSUBS 0.012293f
C140 B.n106 VSUBS 0.012293f
C141 B.n107 VSUBS 0.012293f
C142 B.n108 VSUBS 0.012293f
C143 B.n109 VSUBS 0.012293f
C144 B.n110 VSUBS 0.012293f
C145 B.n111 VSUBS 0.012293f
C146 B.n112 VSUBS 0.012293f
C147 B.n113 VSUBS 0.012293f
C148 B.n114 VSUBS 0.012293f
C149 B.n115 VSUBS 0.012293f
C150 B.n116 VSUBS 0.012293f
C151 B.n117 VSUBS 0.012293f
C152 B.n118 VSUBS 0.012293f
C153 B.n119 VSUBS 0.012293f
C154 B.n120 VSUBS 0.012293f
C155 B.n121 VSUBS 0.012293f
C156 B.n122 VSUBS 0.012293f
C157 B.n123 VSUBS 0.012293f
C158 B.n124 VSUBS 0.012293f
C159 B.n125 VSUBS 0.012293f
C160 B.n126 VSUBS 0.012293f
C161 B.n127 VSUBS 0.02933f
C162 B.n128 VSUBS 0.012293f
C163 B.n129 VSUBS 0.012293f
C164 B.n130 VSUBS 0.012293f
C165 B.n131 VSUBS 0.012293f
C166 B.n132 VSUBS 0.012293f
C167 B.n133 VSUBS 0.012293f
C168 B.n134 VSUBS 0.012293f
C169 B.n135 VSUBS 0.012293f
C170 B.n136 VSUBS 0.012293f
C171 B.n137 VSUBS 0.012293f
C172 B.t8 VSUBS 0.134684f
C173 B.t7 VSUBS 0.178925f
C174 B.t6 VSUBS 1.20945f
C175 B.n138 VSUBS 0.307087f
C176 B.n139 VSUBS 0.250685f
C177 B.n140 VSUBS 0.028482f
C178 B.n141 VSUBS 0.012293f
C179 B.n142 VSUBS 0.012293f
C180 B.n143 VSUBS 0.012293f
C181 B.n144 VSUBS 0.012293f
C182 B.n145 VSUBS 0.012293f
C183 B.t5 VSUBS 0.134681f
C184 B.t4 VSUBS 0.178922f
C185 B.t3 VSUBS 1.20945f
C186 B.n146 VSUBS 0.307089f
C187 B.n147 VSUBS 0.250688f
C188 B.n148 VSUBS 0.012293f
C189 B.n149 VSUBS 0.012293f
C190 B.n150 VSUBS 0.012293f
C191 B.n151 VSUBS 0.012293f
C192 B.n152 VSUBS 0.012293f
C193 B.n153 VSUBS 0.012293f
C194 B.n154 VSUBS 0.012293f
C195 B.n155 VSUBS 0.012293f
C196 B.n156 VSUBS 0.012293f
C197 B.n157 VSUBS 0.012293f
C198 B.n158 VSUBS 0.02816f
C199 B.n159 VSUBS 0.012293f
C200 B.n160 VSUBS 0.012293f
C201 B.n161 VSUBS 0.012293f
C202 B.n162 VSUBS 0.012293f
C203 B.n163 VSUBS 0.012293f
C204 B.n164 VSUBS 0.012293f
C205 B.n165 VSUBS 0.012293f
C206 B.n166 VSUBS 0.012293f
C207 B.n167 VSUBS 0.012293f
C208 B.n168 VSUBS 0.012293f
C209 B.n169 VSUBS 0.012293f
C210 B.n170 VSUBS 0.012293f
C211 B.n171 VSUBS 0.012293f
C212 B.n172 VSUBS 0.012293f
C213 B.n173 VSUBS 0.012293f
C214 B.n174 VSUBS 0.012293f
C215 B.n175 VSUBS 0.012293f
C216 B.n176 VSUBS 0.012293f
C217 B.n177 VSUBS 0.012293f
C218 B.n178 VSUBS 0.012293f
C219 B.n179 VSUBS 0.012293f
C220 B.n180 VSUBS 0.012293f
C221 B.n181 VSUBS 0.012293f
C222 B.n182 VSUBS 0.012293f
C223 B.n183 VSUBS 0.012293f
C224 B.n184 VSUBS 0.012293f
C225 B.n185 VSUBS 0.012293f
C226 B.n186 VSUBS 0.012293f
C227 B.n187 VSUBS 0.012293f
C228 B.n188 VSUBS 0.012293f
C229 B.n189 VSUBS 0.012293f
C230 B.n190 VSUBS 0.012293f
C231 B.n191 VSUBS 0.012293f
C232 B.n192 VSUBS 0.012293f
C233 B.n193 VSUBS 0.012293f
C234 B.n194 VSUBS 0.012293f
C235 B.n195 VSUBS 0.012293f
C236 B.n196 VSUBS 0.012293f
C237 B.n197 VSUBS 0.012293f
C238 B.n198 VSUBS 0.012293f
C239 B.n199 VSUBS 0.012293f
C240 B.n200 VSUBS 0.012293f
C241 B.n201 VSUBS 0.012293f
C242 B.n202 VSUBS 0.012293f
C243 B.n203 VSUBS 0.012293f
C244 B.n204 VSUBS 0.012293f
C245 B.n205 VSUBS 0.012293f
C246 B.n206 VSUBS 0.012293f
C247 B.n207 VSUBS 0.012293f
C248 B.n208 VSUBS 0.012293f
C249 B.n209 VSUBS 0.012293f
C250 B.n210 VSUBS 0.012293f
C251 B.n211 VSUBS 0.012293f
C252 B.n212 VSUBS 0.012293f
C253 B.n213 VSUBS 0.012293f
C254 B.n214 VSUBS 0.012293f
C255 B.n215 VSUBS 0.012293f
C256 B.n216 VSUBS 0.012293f
C257 B.n217 VSUBS 0.012293f
C258 B.n218 VSUBS 0.012293f
C259 B.n219 VSUBS 0.012293f
C260 B.n220 VSUBS 0.012293f
C261 B.n221 VSUBS 0.012293f
C262 B.n222 VSUBS 0.012293f
C263 B.n223 VSUBS 0.012293f
C264 B.n224 VSUBS 0.012293f
C265 B.n225 VSUBS 0.012293f
C266 B.n226 VSUBS 0.012293f
C267 B.n227 VSUBS 0.012293f
C268 B.n228 VSUBS 0.012293f
C269 B.n229 VSUBS 0.012293f
C270 B.n230 VSUBS 0.012293f
C271 B.n231 VSUBS 0.012293f
C272 B.n232 VSUBS 0.012293f
C273 B.n233 VSUBS 0.012293f
C274 B.n234 VSUBS 0.012293f
C275 B.n235 VSUBS 0.012293f
C276 B.n236 VSUBS 0.012293f
C277 B.n237 VSUBS 0.012293f
C278 B.n238 VSUBS 0.012293f
C279 B.n239 VSUBS 0.012293f
C280 B.n240 VSUBS 0.012293f
C281 B.n241 VSUBS 0.012293f
C282 B.n242 VSUBS 0.012293f
C283 B.n243 VSUBS 0.012293f
C284 B.n244 VSUBS 0.012293f
C285 B.n245 VSUBS 0.012293f
C286 B.n246 VSUBS 0.012293f
C287 B.n247 VSUBS 0.012293f
C288 B.n248 VSUBS 0.012293f
C289 B.n249 VSUBS 0.012293f
C290 B.n250 VSUBS 0.012293f
C291 B.n251 VSUBS 0.012293f
C292 B.n252 VSUBS 0.012293f
C293 B.n253 VSUBS 0.012293f
C294 B.n254 VSUBS 0.012293f
C295 B.n255 VSUBS 0.012293f
C296 B.n256 VSUBS 0.012293f
C297 B.n257 VSUBS 0.012293f
C298 B.n258 VSUBS 0.012293f
C299 B.n259 VSUBS 0.012293f
C300 B.n260 VSUBS 0.012293f
C301 B.n261 VSUBS 0.012293f
C302 B.n262 VSUBS 0.012293f
C303 B.n263 VSUBS 0.012293f
C304 B.n264 VSUBS 0.012293f
C305 B.n265 VSUBS 0.012293f
C306 B.n266 VSUBS 0.012293f
C307 B.n267 VSUBS 0.012293f
C308 B.n268 VSUBS 0.012293f
C309 B.n269 VSUBS 0.012293f
C310 B.n270 VSUBS 0.012293f
C311 B.n271 VSUBS 0.012293f
C312 B.n272 VSUBS 0.012293f
C313 B.n273 VSUBS 0.012293f
C314 B.n274 VSUBS 0.012293f
C315 B.n275 VSUBS 0.012293f
C316 B.n276 VSUBS 0.012293f
C317 B.n277 VSUBS 0.012293f
C318 B.n278 VSUBS 0.012293f
C319 B.n279 VSUBS 0.02816f
C320 B.n280 VSUBS 0.02933f
C321 B.n281 VSUBS 0.02933f
C322 B.n282 VSUBS 0.012293f
C323 B.n283 VSUBS 0.012293f
C324 B.n284 VSUBS 0.012293f
C325 B.n285 VSUBS 0.012293f
C326 B.n286 VSUBS 0.012293f
C327 B.n287 VSUBS 0.012293f
C328 B.n288 VSUBS 0.012293f
C329 B.n289 VSUBS 0.012293f
C330 B.n290 VSUBS 0.012293f
C331 B.n291 VSUBS 0.012293f
C332 B.n292 VSUBS 0.012293f
C333 B.n293 VSUBS 0.012293f
C334 B.n294 VSUBS 0.012293f
C335 B.n295 VSUBS 0.012293f
C336 B.n296 VSUBS 0.012293f
C337 B.n297 VSUBS 0.012293f
C338 B.n298 VSUBS 0.012293f
C339 B.n299 VSUBS 0.012293f
C340 B.n300 VSUBS 0.012293f
C341 B.n301 VSUBS 0.012293f
C342 B.n302 VSUBS 0.012293f
C343 B.n303 VSUBS 0.012293f
C344 B.n304 VSUBS 0.012293f
C345 B.n305 VSUBS 0.012293f
C346 B.n306 VSUBS 0.012293f
C347 B.n307 VSUBS 0.012293f
C348 B.n308 VSUBS 0.012293f
C349 B.n309 VSUBS 0.012293f
C350 B.n310 VSUBS 0.012293f
C351 B.n311 VSUBS 0.012293f
C352 B.n312 VSUBS 0.008497f
C353 B.n313 VSUBS 0.028482f
C354 B.n314 VSUBS 0.009943f
C355 B.n315 VSUBS 0.012293f
C356 B.n316 VSUBS 0.012293f
C357 B.n317 VSUBS 0.012293f
C358 B.n318 VSUBS 0.012293f
C359 B.n319 VSUBS 0.012293f
C360 B.n320 VSUBS 0.012293f
C361 B.n321 VSUBS 0.012293f
C362 B.n322 VSUBS 0.012293f
C363 B.n323 VSUBS 0.012293f
C364 B.n324 VSUBS 0.012293f
C365 B.n325 VSUBS 0.012293f
C366 B.n326 VSUBS 0.009943f
C367 B.n327 VSUBS 0.012293f
C368 B.n328 VSUBS 0.012293f
C369 B.n329 VSUBS 0.008497f
C370 B.n330 VSUBS 0.012293f
C371 B.n331 VSUBS 0.012293f
C372 B.n332 VSUBS 0.012293f
C373 B.n333 VSUBS 0.012293f
C374 B.n334 VSUBS 0.012293f
C375 B.n335 VSUBS 0.012293f
C376 B.n336 VSUBS 0.012293f
C377 B.n337 VSUBS 0.012293f
C378 B.n338 VSUBS 0.012293f
C379 B.n339 VSUBS 0.012293f
C380 B.n340 VSUBS 0.012293f
C381 B.n341 VSUBS 0.012293f
C382 B.n342 VSUBS 0.012293f
C383 B.n343 VSUBS 0.012293f
C384 B.n344 VSUBS 0.012293f
C385 B.n345 VSUBS 0.012293f
C386 B.n346 VSUBS 0.012293f
C387 B.n347 VSUBS 0.012293f
C388 B.n348 VSUBS 0.012293f
C389 B.n349 VSUBS 0.012293f
C390 B.n350 VSUBS 0.012293f
C391 B.n351 VSUBS 0.012293f
C392 B.n352 VSUBS 0.012293f
C393 B.n353 VSUBS 0.012293f
C394 B.n354 VSUBS 0.012293f
C395 B.n355 VSUBS 0.012293f
C396 B.n356 VSUBS 0.012293f
C397 B.n357 VSUBS 0.012293f
C398 B.n358 VSUBS 0.012293f
C399 B.n359 VSUBS 0.012293f
C400 B.n360 VSUBS 0.027876f
C401 B.n361 VSUBS 0.029614f
C402 B.n362 VSUBS 0.02816f
C403 B.n363 VSUBS 0.012293f
C404 B.n364 VSUBS 0.012293f
C405 B.n365 VSUBS 0.012293f
C406 B.n366 VSUBS 0.012293f
C407 B.n367 VSUBS 0.012293f
C408 B.n368 VSUBS 0.012293f
C409 B.n369 VSUBS 0.012293f
C410 B.n370 VSUBS 0.012293f
C411 B.n371 VSUBS 0.012293f
C412 B.n372 VSUBS 0.012293f
C413 B.n373 VSUBS 0.012293f
C414 B.n374 VSUBS 0.012293f
C415 B.n375 VSUBS 0.012293f
C416 B.n376 VSUBS 0.012293f
C417 B.n377 VSUBS 0.012293f
C418 B.n378 VSUBS 0.012293f
C419 B.n379 VSUBS 0.012293f
C420 B.n380 VSUBS 0.012293f
C421 B.n381 VSUBS 0.012293f
C422 B.n382 VSUBS 0.012293f
C423 B.n383 VSUBS 0.012293f
C424 B.n384 VSUBS 0.012293f
C425 B.n385 VSUBS 0.012293f
C426 B.n386 VSUBS 0.012293f
C427 B.n387 VSUBS 0.012293f
C428 B.n388 VSUBS 0.012293f
C429 B.n389 VSUBS 0.012293f
C430 B.n390 VSUBS 0.012293f
C431 B.n391 VSUBS 0.012293f
C432 B.n392 VSUBS 0.012293f
C433 B.n393 VSUBS 0.012293f
C434 B.n394 VSUBS 0.012293f
C435 B.n395 VSUBS 0.012293f
C436 B.n396 VSUBS 0.012293f
C437 B.n397 VSUBS 0.012293f
C438 B.n398 VSUBS 0.012293f
C439 B.n399 VSUBS 0.012293f
C440 B.n400 VSUBS 0.012293f
C441 B.n401 VSUBS 0.012293f
C442 B.n402 VSUBS 0.012293f
C443 B.n403 VSUBS 0.012293f
C444 B.n404 VSUBS 0.012293f
C445 B.n405 VSUBS 0.012293f
C446 B.n406 VSUBS 0.012293f
C447 B.n407 VSUBS 0.012293f
C448 B.n408 VSUBS 0.012293f
C449 B.n409 VSUBS 0.012293f
C450 B.n410 VSUBS 0.012293f
C451 B.n411 VSUBS 0.012293f
C452 B.n412 VSUBS 0.012293f
C453 B.n413 VSUBS 0.012293f
C454 B.n414 VSUBS 0.012293f
C455 B.n415 VSUBS 0.012293f
C456 B.n416 VSUBS 0.012293f
C457 B.n417 VSUBS 0.012293f
C458 B.n418 VSUBS 0.012293f
C459 B.n419 VSUBS 0.012293f
C460 B.n420 VSUBS 0.012293f
C461 B.n421 VSUBS 0.012293f
C462 B.n422 VSUBS 0.012293f
C463 B.n423 VSUBS 0.012293f
C464 B.n424 VSUBS 0.012293f
C465 B.n425 VSUBS 0.012293f
C466 B.n426 VSUBS 0.012293f
C467 B.n427 VSUBS 0.012293f
C468 B.n428 VSUBS 0.012293f
C469 B.n429 VSUBS 0.012293f
C470 B.n430 VSUBS 0.012293f
C471 B.n431 VSUBS 0.012293f
C472 B.n432 VSUBS 0.012293f
C473 B.n433 VSUBS 0.012293f
C474 B.n434 VSUBS 0.012293f
C475 B.n435 VSUBS 0.012293f
C476 B.n436 VSUBS 0.012293f
C477 B.n437 VSUBS 0.012293f
C478 B.n438 VSUBS 0.012293f
C479 B.n439 VSUBS 0.012293f
C480 B.n440 VSUBS 0.012293f
C481 B.n441 VSUBS 0.012293f
C482 B.n442 VSUBS 0.012293f
C483 B.n443 VSUBS 0.012293f
C484 B.n444 VSUBS 0.012293f
C485 B.n445 VSUBS 0.012293f
C486 B.n446 VSUBS 0.012293f
C487 B.n447 VSUBS 0.012293f
C488 B.n448 VSUBS 0.012293f
C489 B.n449 VSUBS 0.012293f
C490 B.n450 VSUBS 0.012293f
C491 B.n451 VSUBS 0.012293f
C492 B.n452 VSUBS 0.012293f
C493 B.n453 VSUBS 0.012293f
C494 B.n454 VSUBS 0.012293f
C495 B.n455 VSUBS 0.012293f
C496 B.n456 VSUBS 0.012293f
C497 B.n457 VSUBS 0.012293f
C498 B.n458 VSUBS 0.012293f
C499 B.n459 VSUBS 0.012293f
C500 B.n460 VSUBS 0.012293f
C501 B.n461 VSUBS 0.012293f
C502 B.n462 VSUBS 0.012293f
C503 B.n463 VSUBS 0.012293f
C504 B.n464 VSUBS 0.012293f
C505 B.n465 VSUBS 0.012293f
C506 B.n466 VSUBS 0.012293f
C507 B.n467 VSUBS 0.012293f
C508 B.n468 VSUBS 0.012293f
C509 B.n469 VSUBS 0.012293f
C510 B.n470 VSUBS 0.012293f
C511 B.n471 VSUBS 0.012293f
C512 B.n472 VSUBS 0.012293f
C513 B.n473 VSUBS 0.012293f
C514 B.n474 VSUBS 0.012293f
C515 B.n475 VSUBS 0.012293f
C516 B.n476 VSUBS 0.012293f
C517 B.n477 VSUBS 0.012293f
C518 B.n478 VSUBS 0.012293f
C519 B.n479 VSUBS 0.012293f
C520 B.n480 VSUBS 0.012293f
C521 B.n481 VSUBS 0.012293f
C522 B.n482 VSUBS 0.012293f
C523 B.n483 VSUBS 0.012293f
C524 B.n484 VSUBS 0.012293f
C525 B.n485 VSUBS 0.012293f
C526 B.n486 VSUBS 0.012293f
C527 B.n487 VSUBS 0.012293f
C528 B.n488 VSUBS 0.012293f
C529 B.n489 VSUBS 0.012293f
C530 B.n490 VSUBS 0.012293f
C531 B.n491 VSUBS 0.012293f
C532 B.n492 VSUBS 0.012293f
C533 B.n493 VSUBS 0.012293f
C534 B.n494 VSUBS 0.012293f
C535 B.n495 VSUBS 0.012293f
C536 B.n496 VSUBS 0.012293f
C537 B.n497 VSUBS 0.012293f
C538 B.n498 VSUBS 0.012293f
C539 B.n499 VSUBS 0.012293f
C540 B.n500 VSUBS 0.012293f
C541 B.n501 VSUBS 0.012293f
C542 B.n502 VSUBS 0.012293f
C543 B.n503 VSUBS 0.012293f
C544 B.n504 VSUBS 0.012293f
C545 B.n505 VSUBS 0.012293f
C546 B.n506 VSUBS 0.012293f
C547 B.n507 VSUBS 0.012293f
C548 B.n508 VSUBS 0.012293f
C549 B.n509 VSUBS 0.012293f
C550 B.n510 VSUBS 0.012293f
C551 B.n511 VSUBS 0.012293f
C552 B.n512 VSUBS 0.012293f
C553 B.n513 VSUBS 0.012293f
C554 B.n514 VSUBS 0.012293f
C555 B.n515 VSUBS 0.012293f
C556 B.n516 VSUBS 0.012293f
C557 B.n517 VSUBS 0.012293f
C558 B.n518 VSUBS 0.012293f
C559 B.n519 VSUBS 0.012293f
C560 B.n520 VSUBS 0.012293f
C561 B.n521 VSUBS 0.012293f
C562 B.n522 VSUBS 0.012293f
C563 B.n523 VSUBS 0.012293f
C564 B.n524 VSUBS 0.012293f
C565 B.n525 VSUBS 0.012293f
C566 B.n526 VSUBS 0.012293f
C567 B.n527 VSUBS 0.012293f
C568 B.n528 VSUBS 0.012293f
C569 B.n529 VSUBS 0.012293f
C570 B.n530 VSUBS 0.012293f
C571 B.n531 VSUBS 0.012293f
C572 B.n532 VSUBS 0.012293f
C573 B.n533 VSUBS 0.012293f
C574 B.n534 VSUBS 0.012293f
C575 B.n535 VSUBS 0.012293f
C576 B.n536 VSUBS 0.012293f
C577 B.n537 VSUBS 0.012293f
C578 B.n538 VSUBS 0.012293f
C579 B.n539 VSUBS 0.012293f
C580 B.n540 VSUBS 0.012293f
C581 B.n541 VSUBS 0.012293f
C582 B.n542 VSUBS 0.012293f
C583 B.n543 VSUBS 0.012293f
C584 B.n544 VSUBS 0.012293f
C585 B.n545 VSUBS 0.012293f
C586 B.n546 VSUBS 0.012293f
C587 B.n547 VSUBS 0.012293f
C588 B.n548 VSUBS 0.012293f
C589 B.n549 VSUBS 0.02816f
C590 B.n550 VSUBS 0.02933f
C591 B.n551 VSUBS 0.02933f
C592 B.n552 VSUBS 0.012293f
C593 B.n553 VSUBS 0.012293f
C594 B.n554 VSUBS 0.012293f
C595 B.n555 VSUBS 0.012293f
C596 B.n556 VSUBS 0.012293f
C597 B.n557 VSUBS 0.012293f
C598 B.n558 VSUBS 0.012293f
C599 B.n559 VSUBS 0.012293f
C600 B.n560 VSUBS 0.012293f
C601 B.n561 VSUBS 0.012293f
C602 B.n562 VSUBS 0.012293f
C603 B.n563 VSUBS 0.012293f
C604 B.n564 VSUBS 0.012293f
C605 B.n565 VSUBS 0.012293f
C606 B.n566 VSUBS 0.012293f
C607 B.n567 VSUBS 0.012293f
C608 B.n568 VSUBS 0.012293f
C609 B.n569 VSUBS 0.012293f
C610 B.n570 VSUBS 0.012293f
C611 B.n571 VSUBS 0.012293f
C612 B.n572 VSUBS 0.012293f
C613 B.n573 VSUBS 0.012293f
C614 B.n574 VSUBS 0.012293f
C615 B.n575 VSUBS 0.012293f
C616 B.n576 VSUBS 0.012293f
C617 B.n577 VSUBS 0.012293f
C618 B.n578 VSUBS 0.012293f
C619 B.n579 VSUBS 0.012293f
C620 B.n580 VSUBS 0.012293f
C621 B.n581 VSUBS 0.012293f
C622 B.n582 VSUBS 0.008497f
C623 B.n583 VSUBS 0.028482f
C624 B.n584 VSUBS 0.009943f
C625 B.n585 VSUBS 0.012293f
C626 B.n586 VSUBS 0.012293f
C627 B.n587 VSUBS 0.012293f
C628 B.n588 VSUBS 0.012293f
C629 B.n589 VSUBS 0.012293f
C630 B.n590 VSUBS 0.012293f
C631 B.n591 VSUBS 0.012293f
C632 B.n592 VSUBS 0.012293f
C633 B.n593 VSUBS 0.012293f
C634 B.n594 VSUBS 0.012293f
C635 B.n595 VSUBS 0.012293f
C636 B.n596 VSUBS 0.009943f
C637 B.n597 VSUBS 0.012293f
C638 B.n598 VSUBS 0.012293f
C639 B.n599 VSUBS 0.008497f
C640 B.n600 VSUBS 0.012293f
C641 B.n601 VSUBS 0.012293f
C642 B.n602 VSUBS 0.012293f
C643 B.n603 VSUBS 0.012293f
C644 B.n604 VSUBS 0.012293f
C645 B.n605 VSUBS 0.012293f
C646 B.n606 VSUBS 0.012293f
C647 B.n607 VSUBS 0.012293f
C648 B.n608 VSUBS 0.012293f
C649 B.n609 VSUBS 0.012293f
C650 B.n610 VSUBS 0.012293f
C651 B.n611 VSUBS 0.012293f
C652 B.n612 VSUBS 0.012293f
C653 B.n613 VSUBS 0.012293f
C654 B.n614 VSUBS 0.012293f
C655 B.n615 VSUBS 0.012293f
C656 B.n616 VSUBS 0.012293f
C657 B.n617 VSUBS 0.012293f
C658 B.n618 VSUBS 0.012293f
C659 B.n619 VSUBS 0.012293f
C660 B.n620 VSUBS 0.012293f
C661 B.n621 VSUBS 0.012293f
C662 B.n622 VSUBS 0.012293f
C663 B.n623 VSUBS 0.012293f
C664 B.n624 VSUBS 0.012293f
C665 B.n625 VSUBS 0.012293f
C666 B.n626 VSUBS 0.012293f
C667 B.n627 VSUBS 0.012293f
C668 B.n628 VSUBS 0.012293f
C669 B.n629 VSUBS 0.012293f
C670 B.n630 VSUBS 0.02933f
C671 B.n631 VSUBS 0.02816f
C672 B.n632 VSUBS 0.02816f
C673 B.n633 VSUBS 0.012293f
C674 B.n634 VSUBS 0.012293f
C675 B.n635 VSUBS 0.012293f
C676 B.n636 VSUBS 0.012293f
C677 B.n637 VSUBS 0.012293f
C678 B.n638 VSUBS 0.012293f
C679 B.n639 VSUBS 0.012293f
C680 B.n640 VSUBS 0.012293f
C681 B.n641 VSUBS 0.012293f
C682 B.n642 VSUBS 0.012293f
C683 B.n643 VSUBS 0.012293f
C684 B.n644 VSUBS 0.012293f
C685 B.n645 VSUBS 0.012293f
C686 B.n646 VSUBS 0.012293f
C687 B.n647 VSUBS 0.012293f
C688 B.n648 VSUBS 0.012293f
C689 B.n649 VSUBS 0.012293f
C690 B.n650 VSUBS 0.012293f
C691 B.n651 VSUBS 0.012293f
C692 B.n652 VSUBS 0.012293f
C693 B.n653 VSUBS 0.012293f
C694 B.n654 VSUBS 0.012293f
C695 B.n655 VSUBS 0.012293f
C696 B.n656 VSUBS 0.012293f
C697 B.n657 VSUBS 0.012293f
C698 B.n658 VSUBS 0.012293f
C699 B.n659 VSUBS 0.012293f
C700 B.n660 VSUBS 0.012293f
C701 B.n661 VSUBS 0.012293f
C702 B.n662 VSUBS 0.012293f
C703 B.n663 VSUBS 0.012293f
C704 B.n664 VSUBS 0.012293f
C705 B.n665 VSUBS 0.012293f
C706 B.n666 VSUBS 0.012293f
C707 B.n667 VSUBS 0.012293f
C708 B.n668 VSUBS 0.012293f
C709 B.n669 VSUBS 0.012293f
C710 B.n670 VSUBS 0.012293f
C711 B.n671 VSUBS 0.012293f
C712 B.n672 VSUBS 0.012293f
C713 B.n673 VSUBS 0.012293f
C714 B.n674 VSUBS 0.012293f
C715 B.n675 VSUBS 0.012293f
C716 B.n676 VSUBS 0.012293f
C717 B.n677 VSUBS 0.012293f
C718 B.n678 VSUBS 0.012293f
C719 B.n679 VSUBS 0.012293f
C720 B.n680 VSUBS 0.012293f
C721 B.n681 VSUBS 0.012293f
C722 B.n682 VSUBS 0.012293f
C723 B.n683 VSUBS 0.012293f
C724 B.n684 VSUBS 0.012293f
C725 B.n685 VSUBS 0.012293f
C726 B.n686 VSUBS 0.012293f
C727 B.n687 VSUBS 0.012293f
C728 B.n688 VSUBS 0.012293f
C729 B.n689 VSUBS 0.012293f
C730 B.n690 VSUBS 0.012293f
C731 B.n691 VSUBS 0.012293f
C732 B.n692 VSUBS 0.012293f
C733 B.n693 VSUBS 0.012293f
C734 B.n694 VSUBS 0.012293f
C735 B.n695 VSUBS 0.012293f
C736 B.n696 VSUBS 0.012293f
C737 B.n697 VSUBS 0.012293f
C738 B.n698 VSUBS 0.012293f
C739 B.n699 VSUBS 0.012293f
C740 B.n700 VSUBS 0.012293f
C741 B.n701 VSUBS 0.012293f
C742 B.n702 VSUBS 0.012293f
C743 B.n703 VSUBS 0.012293f
C744 B.n704 VSUBS 0.012293f
C745 B.n705 VSUBS 0.012293f
C746 B.n706 VSUBS 0.012293f
C747 B.n707 VSUBS 0.012293f
C748 B.n708 VSUBS 0.012293f
C749 B.n709 VSUBS 0.012293f
C750 B.n710 VSUBS 0.012293f
C751 B.n711 VSUBS 0.012293f
C752 B.n712 VSUBS 0.012293f
C753 B.n713 VSUBS 0.012293f
C754 B.n714 VSUBS 0.012293f
C755 B.n715 VSUBS 0.012293f
C756 B.n716 VSUBS 0.012293f
C757 B.n717 VSUBS 0.012293f
C758 B.n718 VSUBS 0.012293f
C759 B.n719 VSUBS 0.012293f
C760 B.n720 VSUBS 0.012293f
C761 B.n721 VSUBS 0.012293f
C762 B.n722 VSUBS 0.012293f
C763 B.n723 VSUBS 0.016042f
C764 B.n724 VSUBS 0.017089f
C765 B.n725 VSUBS 0.033983f
C766 VDD1.n0 VSUBS 0.037506f
C767 VDD1.n1 VSUBS 0.035219f
C768 VDD1.n2 VSUBS 0.018925f
C769 VDD1.n3 VSUBS 0.044733f
C770 VDD1.n4 VSUBS 0.020039f
C771 VDD1.n5 VSUBS 0.035219f
C772 VDD1.n6 VSUBS 0.018925f
C773 VDD1.n7 VSUBS 0.033549f
C774 VDD1.n8 VSUBS 0.028414f
C775 VDD1.t5 VSUBS 0.096358f
C776 VDD1.n9 VSUBS 0.14827f
C777 VDD1.n10 VSUBS 0.687241f
C778 VDD1.n11 VSUBS 0.018925f
C779 VDD1.n12 VSUBS 0.020039f
C780 VDD1.n13 VSUBS 0.044733f
C781 VDD1.n14 VSUBS 0.044733f
C782 VDD1.n15 VSUBS 0.020039f
C783 VDD1.n16 VSUBS 0.018925f
C784 VDD1.n17 VSUBS 0.035219f
C785 VDD1.n18 VSUBS 0.035219f
C786 VDD1.n19 VSUBS 0.018925f
C787 VDD1.n20 VSUBS 0.020039f
C788 VDD1.n21 VSUBS 0.044733f
C789 VDD1.n22 VSUBS 0.104231f
C790 VDD1.n23 VSUBS 0.020039f
C791 VDD1.n24 VSUBS 0.018925f
C792 VDD1.n25 VSUBS 0.079964f
C793 VDD1.n26 VSUBS 0.095721f
C794 VDD1.t0 VSUBS 0.146115f
C795 VDD1.t2 VSUBS 0.146115f
C796 VDD1.n27 VSUBS 0.930512f
C797 VDD1.n28 VSUBS 1.28178f
C798 VDD1.n29 VSUBS 0.037506f
C799 VDD1.n30 VSUBS 0.035219f
C800 VDD1.n31 VSUBS 0.018925f
C801 VDD1.n32 VSUBS 0.044733f
C802 VDD1.n33 VSUBS 0.020039f
C803 VDD1.n34 VSUBS 0.035219f
C804 VDD1.n35 VSUBS 0.018925f
C805 VDD1.n36 VSUBS 0.033549f
C806 VDD1.n37 VSUBS 0.028414f
C807 VDD1.t7 VSUBS 0.096358f
C808 VDD1.n38 VSUBS 0.14827f
C809 VDD1.n39 VSUBS 0.687241f
C810 VDD1.n40 VSUBS 0.018925f
C811 VDD1.n41 VSUBS 0.020039f
C812 VDD1.n42 VSUBS 0.044733f
C813 VDD1.n43 VSUBS 0.044733f
C814 VDD1.n44 VSUBS 0.020039f
C815 VDD1.n45 VSUBS 0.018925f
C816 VDD1.n46 VSUBS 0.035219f
C817 VDD1.n47 VSUBS 0.035219f
C818 VDD1.n48 VSUBS 0.018925f
C819 VDD1.n49 VSUBS 0.020039f
C820 VDD1.n50 VSUBS 0.044733f
C821 VDD1.n51 VSUBS 0.104231f
C822 VDD1.n52 VSUBS 0.020039f
C823 VDD1.n53 VSUBS 0.018925f
C824 VDD1.n54 VSUBS 0.079964f
C825 VDD1.n55 VSUBS 0.095721f
C826 VDD1.t1 VSUBS 0.146115f
C827 VDD1.t4 VSUBS 0.146115f
C828 VDD1.n56 VSUBS 0.930507f
C829 VDD1.n57 VSUBS 1.27024f
C830 VDD1.t3 VSUBS 0.146115f
C831 VDD1.t9 VSUBS 0.146115f
C832 VDD1.n58 VSUBS 0.951794f
C833 VDD1.n59 VSUBS 4.06132f
C834 VDD1.t6 VSUBS 0.146115f
C835 VDD1.t8 VSUBS 0.146115f
C836 VDD1.n60 VSUBS 0.930507f
C837 VDD1.n61 VSUBS 4.08348f
C838 VP.n0 VSUBS 0.053996f
C839 VP.t0 VSUBS 1.55188f
C840 VP.n1 VSUBS 0.073527f
C841 VP.n2 VSUBS 0.040956f
C842 VP.t6 VSUBS 1.55188f
C843 VP.n3 VSUBS 0.590048f
C844 VP.n4 VSUBS 0.040956f
C845 VP.n5 VSUBS 0.033958f
C846 VP.n6 VSUBS 0.040956f
C847 VP.t5 VSUBS 1.55188f
C848 VP.n7 VSUBS 0.076331f
C849 VP.n8 VSUBS 0.040956f
C850 VP.n9 VSUBS 0.076331f
C851 VP.n10 VSUBS 0.040956f
C852 VP.t8 VSUBS 1.55188f
C853 VP.n11 VSUBS 0.041367f
C854 VP.n12 VSUBS 0.040956f
C855 VP.t2 VSUBS 1.55188f
C856 VP.n13 VSUBS 0.730767f
C857 VP.n14 VSUBS 0.053996f
C858 VP.t1 VSUBS 1.55188f
C859 VP.n15 VSUBS 0.073527f
C860 VP.n16 VSUBS 0.040956f
C861 VP.t3 VSUBS 1.55188f
C862 VP.n17 VSUBS 0.590048f
C863 VP.n18 VSUBS 0.040956f
C864 VP.n19 VSUBS 0.033958f
C865 VP.n20 VSUBS 0.040956f
C866 VP.t7 VSUBS 1.55188f
C867 VP.n21 VSUBS 0.076331f
C868 VP.n22 VSUBS 0.040956f
C869 VP.n23 VSUBS 0.076331f
C870 VP.t4 VSUBS 1.90728f
C871 VP.n24 VSUBS 0.681407f
C872 VP.t9 VSUBS 1.55188f
C873 VP.n25 VSUBS 0.700847f
C874 VP.n26 VSUBS 0.044675f
C875 VP.n27 VSUBS 0.402235f
C876 VP.n28 VSUBS 0.040956f
C877 VP.n29 VSUBS 0.040956f
C878 VP.n30 VSUBS 0.079371f
C879 VP.n31 VSUBS 0.033958f
C880 VP.n32 VSUBS 0.082577f
C881 VP.n33 VSUBS 0.040956f
C882 VP.n34 VSUBS 0.040956f
C883 VP.n35 VSUBS 0.040956f
C884 VP.n36 VSUBS 0.628694f
C885 VP.n37 VSUBS 0.076331f
C886 VP.n38 VSUBS 0.082577f
C887 VP.n39 VSUBS 0.040956f
C888 VP.n40 VSUBS 0.040956f
C889 VP.n41 VSUBS 0.040956f
C890 VP.n42 VSUBS 0.079371f
C891 VP.n43 VSUBS 0.076331f
C892 VP.n44 VSUBS 0.044675f
C893 VP.n45 VSUBS 0.040956f
C894 VP.n46 VSUBS 0.040956f
C895 VP.n47 VSUBS 0.070301f
C896 VP.n48 VSUBS 0.081012f
C897 VP.n49 VSUBS 0.041367f
C898 VP.n50 VSUBS 0.040956f
C899 VP.n51 VSUBS 0.040956f
C900 VP.n52 VSUBS 0.040956f
C901 VP.n53 VSUBS 0.076331f
C902 VP.n54 VSUBS 0.050705f
C903 VP.n55 VSUBS 0.730767f
C904 VP.n56 VSUBS 2.20616f
C905 VP.n57 VSUBS 2.23631f
C906 VP.n58 VSUBS 0.053996f
C907 VP.n59 VSUBS 0.050705f
C908 VP.n60 VSUBS 0.076331f
C909 VP.n61 VSUBS 0.073527f
C910 VP.n62 VSUBS 0.040956f
C911 VP.n63 VSUBS 0.040956f
C912 VP.n64 VSUBS 0.040956f
C913 VP.n65 VSUBS 0.081012f
C914 VP.n66 VSUBS 0.070301f
C915 VP.n67 VSUBS 0.590048f
C916 VP.n68 VSUBS 0.044675f
C917 VP.n69 VSUBS 0.040956f
C918 VP.n70 VSUBS 0.040956f
C919 VP.n71 VSUBS 0.040956f
C920 VP.n72 VSUBS 0.079371f
C921 VP.n73 VSUBS 0.033958f
C922 VP.n74 VSUBS 0.082577f
C923 VP.n75 VSUBS 0.040956f
C924 VP.n76 VSUBS 0.040956f
C925 VP.n77 VSUBS 0.040956f
C926 VP.n78 VSUBS 0.628694f
C927 VP.n79 VSUBS 0.076331f
C928 VP.n80 VSUBS 0.082577f
C929 VP.n81 VSUBS 0.040956f
C930 VP.n82 VSUBS 0.040956f
C931 VP.n83 VSUBS 0.040956f
C932 VP.n84 VSUBS 0.079371f
C933 VP.n85 VSUBS 0.076331f
C934 VP.n86 VSUBS 0.044675f
C935 VP.n87 VSUBS 0.040956f
C936 VP.n88 VSUBS 0.040956f
C937 VP.n89 VSUBS 0.070301f
C938 VP.n90 VSUBS 0.081012f
C939 VP.n91 VSUBS 0.041367f
C940 VP.n92 VSUBS 0.040956f
C941 VP.n93 VSUBS 0.040956f
C942 VP.n94 VSUBS 0.040956f
C943 VP.n95 VSUBS 0.076331f
C944 VP.n96 VSUBS 0.050705f
C945 VP.n97 VSUBS 0.730767f
C946 VP.n98 VSUBS 0.070912f
C947 VDD2.n0 VSUBS 0.037371f
C948 VDD2.n1 VSUBS 0.035093f
C949 VDD2.n2 VSUBS 0.018857f
C950 VDD2.n3 VSUBS 0.044572f
C951 VDD2.n4 VSUBS 0.019967f
C952 VDD2.n5 VSUBS 0.035093f
C953 VDD2.n6 VSUBS 0.018857f
C954 VDD2.n7 VSUBS 0.033429f
C955 VDD2.n8 VSUBS 0.028312f
C956 VDD2.t1 VSUBS 0.096012f
C957 VDD2.n9 VSUBS 0.147738f
C958 VDD2.n10 VSUBS 0.684773f
C959 VDD2.n11 VSUBS 0.018857f
C960 VDD2.n12 VSUBS 0.019967f
C961 VDD2.n13 VSUBS 0.044572f
C962 VDD2.n14 VSUBS 0.044572f
C963 VDD2.n15 VSUBS 0.019967f
C964 VDD2.n16 VSUBS 0.018857f
C965 VDD2.n17 VSUBS 0.035093f
C966 VDD2.n18 VSUBS 0.035093f
C967 VDD2.n19 VSUBS 0.018857f
C968 VDD2.n20 VSUBS 0.019967f
C969 VDD2.n21 VSUBS 0.044572f
C970 VDD2.n22 VSUBS 0.103857f
C971 VDD2.n23 VSUBS 0.019967f
C972 VDD2.n24 VSUBS 0.018857f
C973 VDD2.n25 VSUBS 0.079677f
C974 VDD2.n26 VSUBS 0.095377f
C975 VDD2.t3 VSUBS 0.14559f
C976 VDD2.t2 VSUBS 0.14559f
C977 VDD2.n27 VSUBS 0.927166f
C978 VDD2.n28 VSUBS 1.26568f
C979 VDD2.t0 VSUBS 0.14559f
C980 VDD2.t9 VSUBS 0.14559f
C981 VDD2.n29 VSUBS 0.948376f
C982 VDD2.n30 VSUBS 3.87356f
C983 VDD2.n31 VSUBS 0.037371f
C984 VDD2.n32 VSUBS 0.035093f
C985 VDD2.n33 VSUBS 0.018857f
C986 VDD2.n34 VSUBS 0.044572f
C987 VDD2.n35 VSUBS 0.019967f
C988 VDD2.n36 VSUBS 0.035093f
C989 VDD2.n37 VSUBS 0.018857f
C990 VDD2.n38 VSUBS 0.033429f
C991 VDD2.n39 VSUBS 0.028312f
C992 VDD2.t4 VSUBS 0.096012f
C993 VDD2.n40 VSUBS 0.147738f
C994 VDD2.n41 VSUBS 0.684773f
C995 VDD2.n42 VSUBS 0.018857f
C996 VDD2.n43 VSUBS 0.019967f
C997 VDD2.n44 VSUBS 0.044572f
C998 VDD2.n45 VSUBS 0.044572f
C999 VDD2.n46 VSUBS 0.019967f
C1000 VDD2.n47 VSUBS 0.018857f
C1001 VDD2.n48 VSUBS 0.035093f
C1002 VDD2.n49 VSUBS 0.035093f
C1003 VDD2.n50 VSUBS 0.018857f
C1004 VDD2.n51 VSUBS 0.019967f
C1005 VDD2.n52 VSUBS 0.044572f
C1006 VDD2.n53 VSUBS 0.103857f
C1007 VDD2.n54 VSUBS 0.019967f
C1008 VDD2.n55 VSUBS 0.018857f
C1009 VDD2.n56 VSUBS 0.079677f
C1010 VDD2.n57 VSUBS 0.076247f
C1011 VDD2.n58 VSUBS 3.39896f
C1012 VDD2.t6 VSUBS 0.14559f
C1013 VDD2.t5 VSUBS 0.14559f
C1014 VDD2.n59 VSUBS 0.927171f
C1015 VDD2.n60 VSUBS 0.929314f
C1016 VDD2.t7 VSUBS 0.14559f
C1017 VDD2.t8 VSUBS 0.14559f
C1018 VDD2.n61 VSUBS 0.948331f
C1019 VTAIL.t15 VSUBS 0.143736f
C1020 VTAIL.t19 VSUBS 0.143736f
C1021 VTAIL.n0 VSUBS 0.804153f
C1022 VTAIL.n1 VSUBS 1.03405f
C1023 VTAIL.n2 VSUBS 0.036896f
C1024 VTAIL.n3 VSUBS 0.034646f
C1025 VTAIL.n4 VSUBS 0.018617f
C1026 VTAIL.n5 VSUBS 0.044004f
C1027 VTAIL.n6 VSUBS 0.019712f
C1028 VTAIL.n7 VSUBS 0.034646f
C1029 VTAIL.n8 VSUBS 0.018617f
C1030 VTAIL.n9 VSUBS 0.033003f
C1031 VTAIL.n10 VSUBS 0.027952f
C1032 VTAIL.t0 VSUBS 0.094789f
C1033 VTAIL.n11 VSUBS 0.145857f
C1034 VTAIL.n12 VSUBS 0.676054f
C1035 VTAIL.n13 VSUBS 0.018617f
C1036 VTAIL.n14 VSUBS 0.019712f
C1037 VTAIL.n15 VSUBS 0.044004f
C1038 VTAIL.n16 VSUBS 0.044004f
C1039 VTAIL.n17 VSUBS 0.019712f
C1040 VTAIL.n18 VSUBS 0.018617f
C1041 VTAIL.n19 VSUBS 0.034646f
C1042 VTAIL.n20 VSUBS 0.034646f
C1043 VTAIL.n21 VSUBS 0.018617f
C1044 VTAIL.n22 VSUBS 0.019712f
C1045 VTAIL.n23 VSUBS 0.044004f
C1046 VTAIL.n24 VSUBS 0.102535f
C1047 VTAIL.n25 VSUBS 0.019712f
C1048 VTAIL.n26 VSUBS 0.018617f
C1049 VTAIL.n27 VSUBS 0.078663f
C1050 VTAIL.n28 VSUBS 0.051342f
C1051 VTAIL.n29 VSUBS 0.525864f
C1052 VTAIL.t7 VSUBS 0.143736f
C1053 VTAIL.t4 VSUBS 0.143736f
C1054 VTAIL.n30 VSUBS 0.804153f
C1055 VTAIL.n31 VSUBS 1.19742f
C1056 VTAIL.t6 VSUBS 0.143736f
C1057 VTAIL.t1 VSUBS 0.143736f
C1058 VTAIL.n32 VSUBS 0.804153f
C1059 VTAIL.n33 VSUBS 2.46972f
C1060 VTAIL.t11 VSUBS 0.143736f
C1061 VTAIL.t18 VSUBS 0.143736f
C1062 VTAIL.n34 VSUBS 0.804159f
C1063 VTAIL.n35 VSUBS 2.46971f
C1064 VTAIL.t10 VSUBS 0.143736f
C1065 VTAIL.t13 VSUBS 0.143736f
C1066 VTAIL.n36 VSUBS 0.804159f
C1067 VTAIL.n37 VSUBS 1.19741f
C1068 VTAIL.n38 VSUBS 0.036896f
C1069 VTAIL.n39 VSUBS 0.034646f
C1070 VTAIL.n40 VSUBS 0.018617f
C1071 VTAIL.n41 VSUBS 0.044004f
C1072 VTAIL.n42 VSUBS 0.019712f
C1073 VTAIL.n43 VSUBS 0.034646f
C1074 VTAIL.n44 VSUBS 0.018617f
C1075 VTAIL.n45 VSUBS 0.033003f
C1076 VTAIL.n46 VSUBS 0.027952f
C1077 VTAIL.t14 VSUBS 0.094789f
C1078 VTAIL.n47 VSUBS 0.145857f
C1079 VTAIL.n48 VSUBS 0.676054f
C1080 VTAIL.n49 VSUBS 0.018617f
C1081 VTAIL.n50 VSUBS 0.019712f
C1082 VTAIL.n51 VSUBS 0.044004f
C1083 VTAIL.n52 VSUBS 0.044004f
C1084 VTAIL.n53 VSUBS 0.019712f
C1085 VTAIL.n54 VSUBS 0.018617f
C1086 VTAIL.n55 VSUBS 0.034646f
C1087 VTAIL.n56 VSUBS 0.034646f
C1088 VTAIL.n57 VSUBS 0.018617f
C1089 VTAIL.n58 VSUBS 0.019712f
C1090 VTAIL.n59 VSUBS 0.044004f
C1091 VTAIL.n60 VSUBS 0.102535f
C1092 VTAIL.n61 VSUBS 0.019712f
C1093 VTAIL.n62 VSUBS 0.018617f
C1094 VTAIL.n63 VSUBS 0.078663f
C1095 VTAIL.n64 VSUBS 0.051342f
C1096 VTAIL.n65 VSUBS 0.525864f
C1097 VTAIL.t3 VSUBS 0.143736f
C1098 VTAIL.t8 VSUBS 0.143736f
C1099 VTAIL.n66 VSUBS 0.804159f
C1100 VTAIL.n67 VSUBS 1.10166f
C1101 VTAIL.t9 VSUBS 0.143736f
C1102 VTAIL.t5 VSUBS 0.143736f
C1103 VTAIL.n68 VSUBS 0.804159f
C1104 VTAIL.n69 VSUBS 1.19741f
C1105 VTAIL.n70 VSUBS 0.036896f
C1106 VTAIL.n71 VSUBS 0.034646f
C1107 VTAIL.n72 VSUBS 0.018617f
C1108 VTAIL.n73 VSUBS 0.044004f
C1109 VTAIL.n74 VSUBS 0.019712f
C1110 VTAIL.n75 VSUBS 0.034646f
C1111 VTAIL.n76 VSUBS 0.018617f
C1112 VTAIL.n77 VSUBS 0.033003f
C1113 VTAIL.n78 VSUBS 0.027952f
C1114 VTAIL.t2 VSUBS 0.094789f
C1115 VTAIL.n79 VSUBS 0.145857f
C1116 VTAIL.n80 VSUBS 0.676054f
C1117 VTAIL.n81 VSUBS 0.018617f
C1118 VTAIL.n82 VSUBS 0.019712f
C1119 VTAIL.n83 VSUBS 0.044004f
C1120 VTAIL.n84 VSUBS 0.044004f
C1121 VTAIL.n85 VSUBS 0.019712f
C1122 VTAIL.n86 VSUBS 0.018617f
C1123 VTAIL.n87 VSUBS 0.034646f
C1124 VTAIL.n88 VSUBS 0.034646f
C1125 VTAIL.n89 VSUBS 0.018617f
C1126 VTAIL.n90 VSUBS 0.019712f
C1127 VTAIL.n91 VSUBS 0.044004f
C1128 VTAIL.n92 VSUBS 0.102535f
C1129 VTAIL.n93 VSUBS 0.019712f
C1130 VTAIL.n94 VSUBS 0.018617f
C1131 VTAIL.n95 VSUBS 0.078663f
C1132 VTAIL.n96 VSUBS 0.051342f
C1133 VTAIL.n97 VSUBS 1.5975f
C1134 VTAIL.n98 VSUBS 0.036896f
C1135 VTAIL.n99 VSUBS 0.034646f
C1136 VTAIL.n100 VSUBS 0.018617f
C1137 VTAIL.n101 VSUBS 0.044004f
C1138 VTAIL.n102 VSUBS 0.019712f
C1139 VTAIL.n103 VSUBS 0.034646f
C1140 VTAIL.n104 VSUBS 0.018617f
C1141 VTAIL.n105 VSUBS 0.033003f
C1142 VTAIL.n106 VSUBS 0.027952f
C1143 VTAIL.t16 VSUBS 0.094789f
C1144 VTAIL.n107 VSUBS 0.145857f
C1145 VTAIL.n108 VSUBS 0.676054f
C1146 VTAIL.n109 VSUBS 0.018617f
C1147 VTAIL.n110 VSUBS 0.019712f
C1148 VTAIL.n111 VSUBS 0.044004f
C1149 VTAIL.n112 VSUBS 0.044004f
C1150 VTAIL.n113 VSUBS 0.019712f
C1151 VTAIL.n114 VSUBS 0.018617f
C1152 VTAIL.n115 VSUBS 0.034646f
C1153 VTAIL.n116 VSUBS 0.034646f
C1154 VTAIL.n117 VSUBS 0.018617f
C1155 VTAIL.n118 VSUBS 0.019712f
C1156 VTAIL.n119 VSUBS 0.044004f
C1157 VTAIL.n120 VSUBS 0.102535f
C1158 VTAIL.n121 VSUBS 0.019712f
C1159 VTAIL.n122 VSUBS 0.018617f
C1160 VTAIL.n123 VSUBS 0.078663f
C1161 VTAIL.n124 VSUBS 0.051342f
C1162 VTAIL.n125 VSUBS 1.5975f
C1163 VTAIL.t12 VSUBS 0.143736f
C1164 VTAIL.t17 VSUBS 0.143736f
C1165 VTAIL.n126 VSUBS 0.804153f
C1166 VTAIL.n127 VSUBS 0.968611f
C1167 VN.n0 VSUBS 0.048172f
C1168 VN.t0 VSUBS 1.3845f
C1169 VN.n1 VSUBS 0.065597f
C1170 VN.n2 VSUBS 0.036538f
C1171 VN.t9 VSUBS 1.3845f
C1172 VN.n3 VSUBS 0.526408f
C1173 VN.n4 VSUBS 0.036538f
C1174 VN.n5 VSUBS 0.030296f
C1175 VN.n6 VSUBS 0.036538f
C1176 VN.t7 VSUBS 1.3845f
C1177 VN.n7 VSUBS 0.068098f
C1178 VN.n8 VSUBS 0.036538f
C1179 VN.n9 VSUBS 0.068098f
C1180 VN.t8 VSUBS 1.70157f
C1181 VN.n10 VSUBS 0.607914f
C1182 VN.t6 VSUBS 1.3845f
C1183 VN.n11 VSUBS 0.625257f
C1184 VN.n12 VSUBS 0.039857f
C1185 VN.n13 VSUBS 0.358851f
C1186 VN.n14 VSUBS 0.036538f
C1187 VN.n15 VSUBS 0.036538f
C1188 VN.n16 VSUBS 0.070811f
C1189 VN.n17 VSUBS 0.030296f
C1190 VN.n18 VSUBS 0.073671f
C1191 VN.n19 VSUBS 0.036538f
C1192 VN.n20 VSUBS 0.036538f
C1193 VN.n21 VSUBS 0.036538f
C1194 VN.n22 VSUBS 0.560886f
C1195 VN.n23 VSUBS 0.068098f
C1196 VN.n24 VSUBS 0.073671f
C1197 VN.n25 VSUBS 0.036538f
C1198 VN.n26 VSUBS 0.036538f
C1199 VN.n27 VSUBS 0.036538f
C1200 VN.n28 VSUBS 0.070811f
C1201 VN.n29 VSUBS 0.068098f
C1202 VN.n30 VSUBS 0.039857f
C1203 VN.n31 VSUBS 0.036538f
C1204 VN.n32 VSUBS 0.036538f
C1205 VN.n33 VSUBS 0.062719f
C1206 VN.n34 VSUBS 0.072274f
C1207 VN.n35 VSUBS 0.036906f
C1208 VN.n36 VSUBS 0.036538f
C1209 VN.n37 VSUBS 0.036538f
C1210 VN.n38 VSUBS 0.036538f
C1211 VN.n39 VSUBS 0.068098f
C1212 VN.n40 VSUBS 0.045236f
C1213 VN.n41 VSUBS 0.65195f
C1214 VN.n42 VSUBS 0.063263f
C1215 VN.n43 VSUBS 0.048172f
C1216 VN.t5 VSUBS 1.3845f
C1217 VN.n44 VSUBS 0.065597f
C1218 VN.n45 VSUBS 0.036538f
C1219 VN.t3 VSUBS 1.3845f
C1220 VN.n46 VSUBS 0.526408f
C1221 VN.n47 VSUBS 0.036538f
C1222 VN.n48 VSUBS 0.030296f
C1223 VN.n49 VSUBS 0.036538f
C1224 VN.t4 VSUBS 1.3845f
C1225 VN.n50 VSUBS 0.068098f
C1226 VN.n51 VSUBS 0.036538f
C1227 VN.n52 VSUBS 0.068098f
C1228 VN.t1 VSUBS 1.70157f
C1229 VN.n53 VSUBS 0.607914f
C1230 VN.t2 VSUBS 1.3845f
C1231 VN.n54 VSUBS 0.625257f
C1232 VN.n55 VSUBS 0.039857f
C1233 VN.n56 VSUBS 0.358851f
C1234 VN.n57 VSUBS 0.036538f
C1235 VN.n58 VSUBS 0.036538f
C1236 VN.n59 VSUBS 0.070811f
C1237 VN.n60 VSUBS 0.030296f
C1238 VN.n61 VSUBS 0.073671f
C1239 VN.n62 VSUBS 0.036538f
C1240 VN.n63 VSUBS 0.036538f
C1241 VN.n64 VSUBS 0.036538f
C1242 VN.n65 VSUBS 0.560886f
C1243 VN.n66 VSUBS 0.068098f
C1244 VN.n67 VSUBS 0.073671f
C1245 VN.n68 VSUBS 0.036538f
C1246 VN.n69 VSUBS 0.036538f
C1247 VN.n70 VSUBS 0.036538f
C1248 VN.n71 VSUBS 0.070811f
C1249 VN.n72 VSUBS 0.068098f
C1250 VN.n73 VSUBS 0.039857f
C1251 VN.n74 VSUBS 0.036538f
C1252 VN.n75 VSUBS 0.036538f
C1253 VN.n76 VSUBS 0.062719f
C1254 VN.n77 VSUBS 0.072274f
C1255 VN.n78 VSUBS 0.036906f
C1256 VN.n79 VSUBS 0.036538f
C1257 VN.n80 VSUBS 0.036538f
C1258 VN.n81 VSUBS 0.036538f
C1259 VN.n82 VSUBS 0.068098f
C1260 VN.n83 VSUBS 0.045236f
C1261 VN.n84 VSUBS 0.65195f
C1262 VN.n85 VSUBS 1.98792f
.ends

