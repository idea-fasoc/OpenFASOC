* NGSPICE file created from diff_pair_sample_0045.ext - technology: sky130A

.subckt diff_pair_sample_0045 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t3 sky130_fd_pr__nfet_01v8 ad=4.7073 pd=24.92 as=0 ps=0 w=12.07 l=2.58
X1 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=4.7073 pd=24.92 as=0 ps=0 w=12.07 l=2.58
X2 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=4.7073 pd=24.92 as=0 ps=0 w=12.07 l=2.58
X3 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=4.7073 pd=24.92 as=0 ps=0 w=12.07 l=2.58
X4 VDD2.t1 VN.t0 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=4.7073 pd=24.92 as=4.7073 ps=24.92 w=12.07 l=2.58
X5 VDD2.t0 VN.t1 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=4.7073 pd=24.92 as=4.7073 ps=24.92 w=12.07 l=2.58
X6 VDD1.t1 VP.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=4.7073 pd=24.92 as=4.7073 ps=24.92 w=12.07 l=2.58
X7 VDD1.t0 VP.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=4.7073 pd=24.92 as=4.7073 ps=24.92 w=12.07 l=2.58
R0 B.n679 B.n678 585
R1 B.n680 B.n679 585
R2 B.n284 B.n95 585
R3 B.n283 B.n282 585
R4 B.n281 B.n280 585
R5 B.n279 B.n278 585
R6 B.n277 B.n276 585
R7 B.n275 B.n274 585
R8 B.n273 B.n272 585
R9 B.n271 B.n270 585
R10 B.n269 B.n268 585
R11 B.n267 B.n266 585
R12 B.n265 B.n264 585
R13 B.n263 B.n262 585
R14 B.n261 B.n260 585
R15 B.n259 B.n258 585
R16 B.n257 B.n256 585
R17 B.n255 B.n254 585
R18 B.n253 B.n252 585
R19 B.n251 B.n250 585
R20 B.n249 B.n248 585
R21 B.n247 B.n246 585
R22 B.n245 B.n244 585
R23 B.n243 B.n242 585
R24 B.n241 B.n240 585
R25 B.n239 B.n238 585
R26 B.n237 B.n236 585
R27 B.n235 B.n234 585
R28 B.n233 B.n232 585
R29 B.n231 B.n230 585
R30 B.n229 B.n228 585
R31 B.n227 B.n226 585
R32 B.n225 B.n224 585
R33 B.n223 B.n222 585
R34 B.n221 B.n220 585
R35 B.n219 B.n218 585
R36 B.n217 B.n216 585
R37 B.n215 B.n214 585
R38 B.n213 B.n212 585
R39 B.n211 B.n210 585
R40 B.n209 B.n208 585
R41 B.n207 B.n206 585
R42 B.n205 B.n204 585
R43 B.n202 B.n201 585
R44 B.n200 B.n199 585
R45 B.n198 B.n197 585
R46 B.n196 B.n195 585
R47 B.n194 B.n193 585
R48 B.n192 B.n191 585
R49 B.n190 B.n189 585
R50 B.n188 B.n187 585
R51 B.n186 B.n185 585
R52 B.n184 B.n183 585
R53 B.n182 B.n181 585
R54 B.n180 B.n179 585
R55 B.n178 B.n177 585
R56 B.n176 B.n175 585
R57 B.n174 B.n173 585
R58 B.n172 B.n171 585
R59 B.n170 B.n169 585
R60 B.n168 B.n167 585
R61 B.n166 B.n165 585
R62 B.n164 B.n163 585
R63 B.n162 B.n161 585
R64 B.n160 B.n159 585
R65 B.n158 B.n157 585
R66 B.n156 B.n155 585
R67 B.n154 B.n153 585
R68 B.n152 B.n151 585
R69 B.n150 B.n149 585
R70 B.n148 B.n147 585
R71 B.n146 B.n145 585
R72 B.n144 B.n143 585
R73 B.n142 B.n141 585
R74 B.n140 B.n139 585
R75 B.n138 B.n137 585
R76 B.n136 B.n135 585
R77 B.n134 B.n133 585
R78 B.n132 B.n131 585
R79 B.n130 B.n129 585
R80 B.n128 B.n127 585
R81 B.n126 B.n125 585
R82 B.n124 B.n123 585
R83 B.n122 B.n121 585
R84 B.n120 B.n119 585
R85 B.n118 B.n117 585
R86 B.n116 B.n115 585
R87 B.n114 B.n113 585
R88 B.n112 B.n111 585
R89 B.n110 B.n109 585
R90 B.n108 B.n107 585
R91 B.n106 B.n105 585
R92 B.n104 B.n103 585
R93 B.n102 B.n101 585
R94 B.n677 B.n48 585
R95 B.n681 B.n48 585
R96 B.n676 B.n47 585
R97 B.n682 B.n47 585
R98 B.n675 B.n674 585
R99 B.n674 B.n43 585
R100 B.n673 B.n42 585
R101 B.n688 B.n42 585
R102 B.n672 B.n41 585
R103 B.n689 B.n41 585
R104 B.n671 B.n40 585
R105 B.n690 B.n40 585
R106 B.n670 B.n669 585
R107 B.n669 B.n36 585
R108 B.n668 B.n35 585
R109 B.n696 B.n35 585
R110 B.n667 B.n34 585
R111 B.n697 B.n34 585
R112 B.n666 B.n33 585
R113 B.n698 B.n33 585
R114 B.n665 B.n664 585
R115 B.n664 B.n29 585
R116 B.n663 B.n28 585
R117 B.n704 B.n28 585
R118 B.n662 B.n27 585
R119 B.n705 B.n27 585
R120 B.n661 B.n26 585
R121 B.n706 B.n26 585
R122 B.n660 B.n659 585
R123 B.n659 B.n22 585
R124 B.n658 B.n21 585
R125 B.n712 B.n21 585
R126 B.n657 B.n20 585
R127 B.n713 B.n20 585
R128 B.n656 B.n19 585
R129 B.n714 B.n19 585
R130 B.n655 B.n654 585
R131 B.n654 B.n15 585
R132 B.n653 B.n14 585
R133 B.n720 B.n14 585
R134 B.n652 B.n13 585
R135 B.n721 B.n13 585
R136 B.n651 B.n12 585
R137 B.n722 B.n12 585
R138 B.n650 B.n649 585
R139 B.n649 B.n8 585
R140 B.n648 B.n7 585
R141 B.n728 B.n7 585
R142 B.n647 B.n6 585
R143 B.n729 B.n6 585
R144 B.n646 B.n5 585
R145 B.n730 B.n5 585
R146 B.n645 B.n644 585
R147 B.n644 B.n4 585
R148 B.n643 B.n285 585
R149 B.n643 B.n642 585
R150 B.n633 B.n286 585
R151 B.n287 B.n286 585
R152 B.n635 B.n634 585
R153 B.n636 B.n635 585
R154 B.n632 B.n292 585
R155 B.n292 B.n291 585
R156 B.n631 B.n630 585
R157 B.n630 B.n629 585
R158 B.n294 B.n293 585
R159 B.n295 B.n294 585
R160 B.n622 B.n621 585
R161 B.n623 B.n622 585
R162 B.n620 B.n300 585
R163 B.n300 B.n299 585
R164 B.n619 B.n618 585
R165 B.n618 B.n617 585
R166 B.n302 B.n301 585
R167 B.n303 B.n302 585
R168 B.n610 B.n609 585
R169 B.n611 B.n610 585
R170 B.n608 B.n308 585
R171 B.n308 B.n307 585
R172 B.n607 B.n606 585
R173 B.n606 B.n605 585
R174 B.n310 B.n309 585
R175 B.n311 B.n310 585
R176 B.n598 B.n597 585
R177 B.n599 B.n598 585
R178 B.n596 B.n316 585
R179 B.n316 B.n315 585
R180 B.n595 B.n594 585
R181 B.n594 B.n593 585
R182 B.n318 B.n317 585
R183 B.n319 B.n318 585
R184 B.n586 B.n585 585
R185 B.n587 B.n586 585
R186 B.n584 B.n324 585
R187 B.n324 B.n323 585
R188 B.n583 B.n582 585
R189 B.n582 B.n581 585
R190 B.n326 B.n325 585
R191 B.n327 B.n326 585
R192 B.n574 B.n573 585
R193 B.n575 B.n574 585
R194 B.n572 B.n332 585
R195 B.n332 B.n331 585
R196 B.n566 B.n565 585
R197 B.n564 B.n380 585
R198 B.n563 B.n379 585
R199 B.n568 B.n379 585
R200 B.n562 B.n561 585
R201 B.n560 B.n559 585
R202 B.n558 B.n557 585
R203 B.n556 B.n555 585
R204 B.n554 B.n553 585
R205 B.n552 B.n551 585
R206 B.n550 B.n549 585
R207 B.n548 B.n547 585
R208 B.n546 B.n545 585
R209 B.n544 B.n543 585
R210 B.n542 B.n541 585
R211 B.n540 B.n539 585
R212 B.n538 B.n537 585
R213 B.n536 B.n535 585
R214 B.n534 B.n533 585
R215 B.n532 B.n531 585
R216 B.n530 B.n529 585
R217 B.n528 B.n527 585
R218 B.n526 B.n525 585
R219 B.n524 B.n523 585
R220 B.n522 B.n521 585
R221 B.n520 B.n519 585
R222 B.n518 B.n517 585
R223 B.n516 B.n515 585
R224 B.n514 B.n513 585
R225 B.n512 B.n511 585
R226 B.n510 B.n509 585
R227 B.n508 B.n507 585
R228 B.n506 B.n505 585
R229 B.n504 B.n503 585
R230 B.n502 B.n501 585
R231 B.n500 B.n499 585
R232 B.n498 B.n497 585
R233 B.n496 B.n495 585
R234 B.n494 B.n493 585
R235 B.n492 B.n491 585
R236 B.n490 B.n489 585
R237 B.n488 B.n487 585
R238 B.n486 B.n485 585
R239 B.n483 B.n482 585
R240 B.n481 B.n480 585
R241 B.n479 B.n478 585
R242 B.n477 B.n476 585
R243 B.n475 B.n474 585
R244 B.n473 B.n472 585
R245 B.n471 B.n470 585
R246 B.n469 B.n468 585
R247 B.n467 B.n466 585
R248 B.n465 B.n464 585
R249 B.n463 B.n462 585
R250 B.n461 B.n460 585
R251 B.n459 B.n458 585
R252 B.n457 B.n456 585
R253 B.n455 B.n454 585
R254 B.n453 B.n452 585
R255 B.n451 B.n450 585
R256 B.n449 B.n448 585
R257 B.n447 B.n446 585
R258 B.n445 B.n444 585
R259 B.n443 B.n442 585
R260 B.n441 B.n440 585
R261 B.n439 B.n438 585
R262 B.n437 B.n436 585
R263 B.n435 B.n434 585
R264 B.n433 B.n432 585
R265 B.n431 B.n430 585
R266 B.n429 B.n428 585
R267 B.n427 B.n426 585
R268 B.n425 B.n424 585
R269 B.n423 B.n422 585
R270 B.n421 B.n420 585
R271 B.n419 B.n418 585
R272 B.n417 B.n416 585
R273 B.n415 B.n414 585
R274 B.n413 B.n412 585
R275 B.n411 B.n410 585
R276 B.n409 B.n408 585
R277 B.n407 B.n406 585
R278 B.n405 B.n404 585
R279 B.n403 B.n402 585
R280 B.n401 B.n400 585
R281 B.n399 B.n398 585
R282 B.n397 B.n396 585
R283 B.n395 B.n394 585
R284 B.n393 B.n392 585
R285 B.n391 B.n390 585
R286 B.n389 B.n388 585
R287 B.n387 B.n386 585
R288 B.n334 B.n333 585
R289 B.n571 B.n570 585
R290 B.n330 B.n329 585
R291 B.n331 B.n330 585
R292 B.n577 B.n576 585
R293 B.n576 B.n575 585
R294 B.n578 B.n328 585
R295 B.n328 B.n327 585
R296 B.n580 B.n579 585
R297 B.n581 B.n580 585
R298 B.n322 B.n321 585
R299 B.n323 B.n322 585
R300 B.n589 B.n588 585
R301 B.n588 B.n587 585
R302 B.n590 B.n320 585
R303 B.n320 B.n319 585
R304 B.n592 B.n591 585
R305 B.n593 B.n592 585
R306 B.n314 B.n313 585
R307 B.n315 B.n314 585
R308 B.n601 B.n600 585
R309 B.n600 B.n599 585
R310 B.n602 B.n312 585
R311 B.n312 B.n311 585
R312 B.n604 B.n603 585
R313 B.n605 B.n604 585
R314 B.n306 B.n305 585
R315 B.n307 B.n306 585
R316 B.n613 B.n612 585
R317 B.n612 B.n611 585
R318 B.n614 B.n304 585
R319 B.n304 B.n303 585
R320 B.n616 B.n615 585
R321 B.n617 B.n616 585
R322 B.n298 B.n297 585
R323 B.n299 B.n298 585
R324 B.n625 B.n624 585
R325 B.n624 B.n623 585
R326 B.n626 B.n296 585
R327 B.n296 B.n295 585
R328 B.n628 B.n627 585
R329 B.n629 B.n628 585
R330 B.n290 B.n289 585
R331 B.n291 B.n290 585
R332 B.n638 B.n637 585
R333 B.n637 B.n636 585
R334 B.n639 B.n288 585
R335 B.n288 B.n287 585
R336 B.n641 B.n640 585
R337 B.n642 B.n641 585
R338 B.n2 B.n0 585
R339 B.n4 B.n2 585
R340 B.n3 B.n1 585
R341 B.n729 B.n3 585
R342 B.n727 B.n726 585
R343 B.n728 B.n727 585
R344 B.n725 B.n9 585
R345 B.n9 B.n8 585
R346 B.n724 B.n723 585
R347 B.n723 B.n722 585
R348 B.n11 B.n10 585
R349 B.n721 B.n11 585
R350 B.n719 B.n718 585
R351 B.n720 B.n719 585
R352 B.n717 B.n16 585
R353 B.n16 B.n15 585
R354 B.n716 B.n715 585
R355 B.n715 B.n714 585
R356 B.n18 B.n17 585
R357 B.n713 B.n18 585
R358 B.n711 B.n710 585
R359 B.n712 B.n711 585
R360 B.n709 B.n23 585
R361 B.n23 B.n22 585
R362 B.n708 B.n707 585
R363 B.n707 B.n706 585
R364 B.n25 B.n24 585
R365 B.n705 B.n25 585
R366 B.n703 B.n702 585
R367 B.n704 B.n703 585
R368 B.n701 B.n30 585
R369 B.n30 B.n29 585
R370 B.n700 B.n699 585
R371 B.n699 B.n698 585
R372 B.n32 B.n31 585
R373 B.n697 B.n32 585
R374 B.n695 B.n694 585
R375 B.n696 B.n695 585
R376 B.n693 B.n37 585
R377 B.n37 B.n36 585
R378 B.n692 B.n691 585
R379 B.n691 B.n690 585
R380 B.n39 B.n38 585
R381 B.n689 B.n39 585
R382 B.n687 B.n686 585
R383 B.n688 B.n687 585
R384 B.n685 B.n44 585
R385 B.n44 B.n43 585
R386 B.n684 B.n683 585
R387 B.n683 B.n682 585
R388 B.n46 B.n45 585
R389 B.n681 B.n46 585
R390 B.n732 B.n731 585
R391 B.n731 B.n730 585
R392 B.n566 B.n330 554.963
R393 B.n101 B.n46 554.963
R394 B.n570 B.n332 554.963
R395 B.n679 B.n48 554.963
R396 B.n383 B.t9 339.803
R397 B.n96 B.t14 339.803
R398 B.n381 B.t12 339.803
R399 B.n98 B.t4 339.803
R400 B.n383 B.t6 320.764
R401 B.n381 B.t10 320.764
R402 B.n98 B.t2 320.764
R403 B.n96 B.t13 320.764
R404 B.n384 B.t8 283.365
R405 B.n97 B.t15 283.365
R406 B.n382 B.t11 283.365
R407 B.n99 B.t5 283.365
R408 B.n680 B.n94 256.663
R409 B.n680 B.n93 256.663
R410 B.n680 B.n92 256.663
R411 B.n680 B.n91 256.663
R412 B.n680 B.n90 256.663
R413 B.n680 B.n89 256.663
R414 B.n680 B.n88 256.663
R415 B.n680 B.n87 256.663
R416 B.n680 B.n86 256.663
R417 B.n680 B.n85 256.663
R418 B.n680 B.n84 256.663
R419 B.n680 B.n83 256.663
R420 B.n680 B.n82 256.663
R421 B.n680 B.n81 256.663
R422 B.n680 B.n80 256.663
R423 B.n680 B.n79 256.663
R424 B.n680 B.n78 256.663
R425 B.n680 B.n77 256.663
R426 B.n680 B.n76 256.663
R427 B.n680 B.n75 256.663
R428 B.n680 B.n74 256.663
R429 B.n680 B.n73 256.663
R430 B.n680 B.n72 256.663
R431 B.n680 B.n71 256.663
R432 B.n680 B.n70 256.663
R433 B.n680 B.n69 256.663
R434 B.n680 B.n68 256.663
R435 B.n680 B.n67 256.663
R436 B.n680 B.n66 256.663
R437 B.n680 B.n65 256.663
R438 B.n680 B.n64 256.663
R439 B.n680 B.n63 256.663
R440 B.n680 B.n62 256.663
R441 B.n680 B.n61 256.663
R442 B.n680 B.n60 256.663
R443 B.n680 B.n59 256.663
R444 B.n680 B.n58 256.663
R445 B.n680 B.n57 256.663
R446 B.n680 B.n56 256.663
R447 B.n680 B.n55 256.663
R448 B.n680 B.n54 256.663
R449 B.n680 B.n53 256.663
R450 B.n680 B.n52 256.663
R451 B.n680 B.n51 256.663
R452 B.n680 B.n50 256.663
R453 B.n680 B.n49 256.663
R454 B.n568 B.n567 256.663
R455 B.n568 B.n335 256.663
R456 B.n568 B.n336 256.663
R457 B.n568 B.n337 256.663
R458 B.n568 B.n338 256.663
R459 B.n568 B.n339 256.663
R460 B.n568 B.n340 256.663
R461 B.n568 B.n341 256.663
R462 B.n568 B.n342 256.663
R463 B.n568 B.n343 256.663
R464 B.n568 B.n344 256.663
R465 B.n568 B.n345 256.663
R466 B.n568 B.n346 256.663
R467 B.n568 B.n347 256.663
R468 B.n568 B.n348 256.663
R469 B.n568 B.n349 256.663
R470 B.n568 B.n350 256.663
R471 B.n568 B.n351 256.663
R472 B.n568 B.n352 256.663
R473 B.n568 B.n353 256.663
R474 B.n568 B.n354 256.663
R475 B.n568 B.n355 256.663
R476 B.n568 B.n356 256.663
R477 B.n568 B.n357 256.663
R478 B.n568 B.n358 256.663
R479 B.n568 B.n359 256.663
R480 B.n568 B.n360 256.663
R481 B.n568 B.n361 256.663
R482 B.n568 B.n362 256.663
R483 B.n568 B.n363 256.663
R484 B.n568 B.n364 256.663
R485 B.n568 B.n365 256.663
R486 B.n568 B.n366 256.663
R487 B.n568 B.n367 256.663
R488 B.n568 B.n368 256.663
R489 B.n568 B.n369 256.663
R490 B.n568 B.n370 256.663
R491 B.n568 B.n371 256.663
R492 B.n568 B.n372 256.663
R493 B.n568 B.n373 256.663
R494 B.n568 B.n374 256.663
R495 B.n568 B.n375 256.663
R496 B.n568 B.n376 256.663
R497 B.n568 B.n377 256.663
R498 B.n568 B.n378 256.663
R499 B.n569 B.n568 256.663
R500 B.n576 B.n330 163.367
R501 B.n576 B.n328 163.367
R502 B.n580 B.n328 163.367
R503 B.n580 B.n322 163.367
R504 B.n588 B.n322 163.367
R505 B.n588 B.n320 163.367
R506 B.n592 B.n320 163.367
R507 B.n592 B.n314 163.367
R508 B.n600 B.n314 163.367
R509 B.n600 B.n312 163.367
R510 B.n604 B.n312 163.367
R511 B.n604 B.n306 163.367
R512 B.n612 B.n306 163.367
R513 B.n612 B.n304 163.367
R514 B.n616 B.n304 163.367
R515 B.n616 B.n298 163.367
R516 B.n624 B.n298 163.367
R517 B.n624 B.n296 163.367
R518 B.n628 B.n296 163.367
R519 B.n628 B.n290 163.367
R520 B.n637 B.n290 163.367
R521 B.n637 B.n288 163.367
R522 B.n641 B.n288 163.367
R523 B.n641 B.n2 163.367
R524 B.n731 B.n2 163.367
R525 B.n731 B.n3 163.367
R526 B.n727 B.n3 163.367
R527 B.n727 B.n9 163.367
R528 B.n723 B.n9 163.367
R529 B.n723 B.n11 163.367
R530 B.n719 B.n11 163.367
R531 B.n719 B.n16 163.367
R532 B.n715 B.n16 163.367
R533 B.n715 B.n18 163.367
R534 B.n711 B.n18 163.367
R535 B.n711 B.n23 163.367
R536 B.n707 B.n23 163.367
R537 B.n707 B.n25 163.367
R538 B.n703 B.n25 163.367
R539 B.n703 B.n30 163.367
R540 B.n699 B.n30 163.367
R541 B.n699 B.n32 163.367
R542 B.n695 B.n32 163.367
R543 B.n695 B.n37 163.367
R544 B.n691 B.n37 163.367
R545 B.n691 B.n39 163.367
R546 B.n687 B.n39 163.367
R547 B.n687 B.n44 163.367
R548 B.n683 B.n44 163.367
R549 B.n683 B.n46 163.367
R550 B.n380 B.n379 163.367
R551 B.n561 B.n379 163.367
R552 B.n559 B.n558 163.367
R553 B.n555 B.n554 163.367
R554 B.n551 B.n550 163.367
R555 B.n547 B.n546 163.367
R556 B.n543 B.n542 163.367
R557 B.n539 B.n538 163.367
R558 B.n535 B.n534 163.367
R559 B.n531 B.n530 163.367
R560 B.n527 B.n526 163.367
R561 B.n523 B.n522 163.367
R562 B.n519 B.n518 163.367
R563 B.n515 B.n514 163.367
R564 B.n511 B.n510 163.367
R565 B.n507 B.n506 163.367
R566 B.n503 B.n502 163.367
R567 B.n499 B.n498 163.367
R568 B.n495 B.n494 163.367
R569 B.n491 B.n490 163.367
R570 B.n487 B.n486 163.367
R571 B.n482 B.n481 163.367
R572 B.n478 B.n477 163.367
R573 B.n474 B.n473 163.367
R574 B.n470 B.n469 163.367
R575 B.n466 B.n465 163.367
R576 B.n462 B.n461 163.367
R577 B.n458 B.n457 163.367
R578 B.n454 B.n453 163.367
R579 B.n450 B.n449 163.367
R580 B.n446 B.n445 163.367
R581 B.n442 B.n441 163.367
R582 B.n438 B.n437 163.367
R583 B.n434 B.n433 163.367
R584 B.n430 B.n429 163.367
R585 B.n426 B.n425 163.367
R586 B.n422 B.n421 163.367
R587 B.n418 B.n417 163.367
R588 B.n414 B.n413 163.367
R589 B.n410 B.n409 163.367
R590 B.n406 B.n405 163.367
R591 B.n402 B.n401 163.367
R592 B.n398 B.n397 163.367
R593 B.n394 B.n393 163.367
R594 B.n390 B.n389 163.367
R595 B.n386 B.n334 163.367
R596 B.n574 B.n332 163.367
R597 B.n574 B.n326 163.367
R598 B.n582 B.n326 163.367
R599 B.n582 B.n324 163.367
R600 B.n586 B.n324 163.367
R601 B.n586 B.n318 163.367
R602 B.n594 B.n318 163.367
R603 B.n594 B.n316 163.367
R604 B.n598 B.n316 163.367
R605 B.n598 B.n310 163.367
R606 B.n606 B.n310 163.367
R607 B.n606 B.n308 163.367
R608 B.n610 B.n308 163.367
R609 B.n610 B.n302 163.367
R610 B.n618 B.n302 163.367
R611 B.n618 B.n300 163.367
R612 B.n622 B.n300 163.367
R613 B.n622 B.n294 163.367
R614 B.n630 B.n294 163.367
R615 B.n630 B.n292 163.367
R616 B.n635 B.n292 163.367
R617 B.n635 B.n286 163.367
R618 B.n643 B.n286 163.367
R619 B.n644 B.n643 163.367
R620 B.n644 B.n5 163.367
R621 B.n6 B.n5 163.367
R622 B.n7 B.n6 163.367
R623 B.n649 B.n7 163.367
R624 B.n649 B.n12 163.367
R625 B.n13 B.n12 163.367
R626 B.n14 B.n13 163.367
R627 B.n654 B.n14 163.367
R628 B.n654 B.n19 163.367
R629 B.n20 B.n19 163.367
R630 B.n21 B.n20 163.367
R631 B.n659 B.n21 163.367
R632 B.n659 B.n26 163.367
R633 B.n27 B.n26 163.367
R634 B.n28 B.n27 163.367
R635 B.n664 B.n28 163.367
R636 B.n664 B.n33 163.367
R637 B.n34 B.n33 163.367
R638 B.n35 B.n34 163.367
R639 B.n669 B.n35 163.367
R640 B.n669 B.n40 163.367
R641 B.n41 B.n40 163.367
R642 B.n42 B.n41 163.367
R643 B.n674 B.n42 163.367
R644 B.n674 B.n47 163.367
R645 B.n48 B.n47 163.367
R646 B.n105 B.n104 163.367
R647 B.n109 B.n108 163.367
R648 B.n113 B.n112 163.367
R649 B.n117 B.n116 163.367
R650 B.n121 B.n120 163.367
R651 B.n125 B.n124 163.367
R652 B.n129 B.n128 163.367
R653 B.n133 B.n132 163.367
R654 B.n137 B.n136 163.367
R655 B.n141 B.n140 163.367
R656 B.n145 B.n144 163.367
R657 B.n149 B.n148 163.367
R658 B.n153 B.n152 163.367
R659 B.n157 B.n156 163.367
R660 B.n161 B.n160 163.367
R661 B.n165 B.n164 163.367
R662 B.n169 B.n168 163.367
R663 B.n173 B.n172 163.367
R664 B.n177 B.n176 163.367
R665 B.n181 B.n180 163.367
R666 B.n185 B.n184 163.367
R667 B.n189 B.n188 163.367
R668 B.n193 B.n192 163.367
R669 B.n197 B.n196 163.367
R670 B.n201 B.n200 163.367
R671 B.n206 B.n205 163.367
R672 B.n210 B.n209 163.367
R673 B.n214 B.n213 163.367
R674 B.n218 B.n217 163.367
R675 B.n222 B.n221 163.367
R676 B.n226 B.n225 163.367
R677 B.n230 B.n229 163.367
R678 B.n234 B.n233 163.367
R679 B.n238 B.n237 163.367
R680 B.n242 B.n241 163.367
R681 B.n246 B.n245 163.367
R682 B.n250 B.n249 163.367
R683 B.n254 B.n253 163.367
R684 B.n258 B.n257 163.367
R685 B.n262 B.n261 163.367
R686 B.n266 B.n265 163.367
R687 B.n270 B.n269 163.367
R688 B.n274 B.n273 163.367
R689 B.n278 B.n277 163.367
R690 B.n282 B.n281 163.367
R691 B.n679 B.n95 163.367
R692 B.n568 B.n331 88.1527
R693 B.n681 B.n680 88.1527
R694 B.n567 B.n566 71.676
R695 B.n561 B.n335 71.676
R696 B.n558 B.n336 71.676
R697 B.n554 B.n337 71.676
R698 B.n550 B.n338 71.676
R699 B.n546 B.n339 71.676
R700 B.n542 B.n340 71.676
R701 B.n538 B.n341 71.676
R702 B.n534 B.n342 71.676
R703 B.n530 B.n343 71.676
R704 B.n526 B.n344 71.676
R705 B.n522 B.n345 71.676
R706 B.n518 B.n346 71.676
R707 B.n514 B.n347 71.676
R708 B.n510 B.n348 71.676
R709 B.n506 B.n349 71.676
R710 B.n502 B.n350 71.676
R711 B.n498 B.n351 71.676
R712 B.n494 B.n352 71.676
R713 B.n490 B.n353 71.676
R714 B.n486 B.n354 71.676
R715 B.n481 B.n355 71.676
R716 B.n477 B.n356 71.676
R717 B.n473 B.n357 71.676
R718 B.n469 B.n358 71.676
R719 B.n465 B.n359 71.676
R720 B.n461 B.n360 71.676
R721 B.n457 B.n361 71.676
R722 B.n453 B.n362 71.676
R723 B.n449 B.n363 71.676
R724 B.n445 B.n364 71.676
R725 B.n441 B.n365 71.676
R726 B.n437 B.n366 71.676
R727 B.n433 B.n367 71.676
R728 B.n429 B.n368 71.676
R729 B.n425 B.n369 71.676
R730 B.n421 B.n370 71.676
R731 B.n417 B.n371 71.676
R732 B.n413 B.n372 71.676
R733 B.n409 B.n373 71.676
R734 B.n405 B.n374 71.676
R735 B.n401 B.n375 71.676
R736 B.n397 B.n376 71.676
R737 B.n393 B.n377 71.676
R738 B.n389 B.n378 71.676
R739 B.n569 B.n334 71.676
R740 B.n101 B.n49 71.676
R741 B.n105 B.n50 71.676
R742 B.n109 B.n51 71.676
R743 B.n113 B.n52 71.676
R744 B.n117 B.n53 71.676
R745 B.n121 B.n54 71.676
R746 B.n125 B.n55 71.676
R747 B.n129 B.n56 71.676
R748 B.n133 B.n57 71.676
R749 B.n137 B.n58 71.676
R750 B.n141 B.n59 71.676
R751 B.n145 B.n60 71.676
R752 B.n149 B.n61 71.676
R753 B.n153 B.n62 71.676
R754 B.n157 B.n63 71.676
R755 B.n161 B.n64 71.676
R756 B.n165 B.n65 71.676
R757 B.n169 B.n66 71.676
R758 B.n173 B.n67 71.676
R759 B.n177 B.n68 71.676
R760 B.n181 B.n69 71.676
R761 B.n185 B.n70 71.676
R762 B.n189 B.n71 71.676
R763 B.n193 B.n72 71.676
R764 B.n197 B.n73 71.676
R765 B.n201 B.n74 71.676
R766 B.n206 B.n75 71.676
R767 B.n210 B.n76 71.676
R768 B.n214 B.n77 71.676
R769 B.n218 B.n78 71.676
R770 B.n222 B.n79 71.676
R771 B.n226 B.n80 71.676
R772 B.n230 B.n81 71.676
R773 B.n234 B.n82 71.676
R774 B.n238 B.n83 71.676
R775 B.n242 B.n84 71.676
R776 B.n246 B.n85 71.676
R777 B.n250 B.n86 71.676
R778 B.n254 B.n87 71.676
R779 B.n258 B.n88 71.676
R780 B.n262 B.n89 71.676
R781 B.n266 B.n90 71.676
R782 B.n270 B.n91 71.676
R783 B.n274 B.n92 71.676
R784 B.n278 B.n93 71.676
R785 B.n282 B.n94 71.676
R786 B.n95 B.n94 71.676
R787 B.n281 B.n93 71.676
R788 B.n277 B.n92 71.676
R789 B.n273 B.n91 71.676
R790 B.n269 B.n90 71.676
R791 B.n265 B.n89 71.676
R792 B.n261 B.n88 71.676
R793 B.n257 B.n87 71.676
R794 B.n253 B.n86 71.676
R795 B.n249 B.n85 71.676
R796 B.n245 B.n84 71.676
R797 B.n241 B.n83 71.676
R798 B.n237 B.n82 71.676
R799 B.n233 B.n81 71.676
R800 B.n229 B.n80 71.676
R801 B.n225 B.n79 71.676
R802 B.n221 B.n78 71.676
R803 B.n217 B.n77 71.676
R804 B.n213 B.n76 71.676
R805 B.n209 B.n75 71.676
R806 B.n205 B.n74 71.676
R807 B.n200 B.n73 71.676
R808 B.n196 B.n72 71.676
R809 B.n192 B.n71 71.676
R810 B.n188 B.n70 71.676
R811 B.n184 B.n69 71.676
R812 B.n180 B.n68 71.676
R813 B.n176 B.n67 71.676
R814 B.n172 B.n66 71.676
R815 B.n168 B.n65 71.676
R816 B.n164 B.n64 71.676
R817 B.n160 B.n63 71.676
R818 B.n156 B.n62 71.676
R819 B.n152 B.n61 71.676
R820 B.n148 B.n60 71.676
R821 B.n144 B.n59 71.676
R822 B.n140 B.n58 71.676
R823 B.n136 B.n57 71.676
R824 B.n132 B.n56 71.676
R825 B.n128 B.n55 71.676
R826 B.n124 B.n54 71.676
R827 B.n120 B.n53 71.676
R828 B.n116 B.n52 71.676
R829 B.n112 B.n51 71.676
R830 B.n108 B.n50 71.676
R831 B.n104 B.n49 71.676
R832 B.n567 B.n380 71.676
R833 B.n559 B.n335 71.676
R834 B.n555 B.n336 71.676
R835 B.n551 B.n337 71.676
R836 B.n547 B.n338 71.676
R837 B.n543 B.n339 71.676
R838 B.n539 B.n340 71.676
R839 B.n535 B.n341 71.676
R840 B.n531 B.n342 71.676
R841 B.n527 B.n343 71.676
R842 B.n523 B.n344 71.676
R843 B.n519 B.n345 71.676
R844 B.n515 B.n346 71.676
R845 B.n511 B.n347 71.676
R846 B.n507 B.n348 71.676
R847 B.n503 B.n349 71.676
R848 B.n499 B.n350 71.676
R849 B.n495 B.n351 71.676
R850 B.n491 B.n352 71.676
R851 B.n487 B.n353 71.676
R852 B.n482 B.n354 71.676
R853 B.n478 B.n355 71.676
R854 B.n474 B.n356 71.676
R855 B.n470 B.n357 71.676
R856 B.n466 B.n358 71.676
R857 B.n462 B.n359 71.676
R858 B.n458 B.n360 71.676
R859 B.n454 B.n361 71.676
R860 B.n450 B.n362 71.676
R861 B.n446 B.n363 71.676
R862 B.n442 B.n364 71.676
R863 B.n438 B.n365 71.676
R864 B.n434 B.n366 71.676
R865 B.n430 B.n367 71.676
R866 B.n426 B.n368 71.676
R867 B.n422 B.n369 71.676
R868 B.n418 B.n370 71.676
R869 B.n414 B.n371 71.676
R870 B.n410 B.n372 71.676
R871 B.n406 B.n373 71.676
R872 B.n402 B.n374 71.676
R873 B.n398 B.n375 71.676
R874 B.n394 B.n376 71.676
R875 B.n390 B.n377 71.676
R876 B.n386 B.n378 71.676
R877 B.n570 B.n569 71.676
R878 B.n385 B.n384 59.5399
R879 B.n484 B.n382 59.5399
R880 B.n100 B.n99 59.5399
R881 B.n203 B.n97 59.5399
R882 B.n384 B.n383 56.4369
R883 B.n382 B.n381 56.4369
R884 B.n99 B.n98 56.4369
R885 B.n97 B.n96 56.4369
R886 B.n575 B.n331 43.1253
R887 B.n575 B.n327 43.1253
R888 B.n581 B.n327 43.1253
R889 B.n581 B.n323 43.1253
R890 B.n587 B.n323 43.1253
R891 B.n587 B.n319 43.1253
R892 B.n593 B.n319 43.1253
R893 B.n599 B.n315 43.1253
R894 B.n599 B.n311 43.1253
R895 B.n605 B.n311 43.1253
R896 B.n605 B.n307 43.1253
R897 B.n611 B.n307 43.1253
R898 B.n611 B.n303 43.1253
R899 B.n617 B.n303 43.1253
R900 B.n617 B.n299 43.1253
R901 B.n623 B.n299 43.1253
R902 B.n623 B.n295 43.1253
R903 B.n629 B.n295 43.1253
R904 B.n636 B.n291 43.1253
R905 B.n636 B.n287 43.1253
R906 B.n642 B.n287 43.1253
R907 B.n642 B.n4 43.1253
R908 B.n730 B.n4 43.1253
R909 B.n730 B.n729 43.1253
R910 B.n729 B.n728 43.1253
R911 B.n728 B.n8 43.1253
R912 B.n722 B.n8 43.1253
R913 B.n722 B.n721 43.1253
R914 B.n720 B.n15 43.1253
R915 B.n714 B.n15 43.1253
R916 B.n714 B.n713 43.1253
R917 B.n713 B.n712 43.1253
R918 B.n712 B.n22 43.1253
R919 B.n706 B.n22 43.1253
R920 B.n706 B.n705 43.1253
R921 B.n705 B.n704 43.1253
R922 B.n704 B.n29 43.1253
R923 B.n698 B.n29 43.1253
R924 B.n698 B.n697 43.1253
R925 B.n696 B.n36 43.1253
R926 B.n690 B.n36 43.1253
R927 B.n690 B.n689 43.1253
R928 B.n689 B.n688 43.1253
R929 B.n688 B.n43 43.1253
R930 B.n682 B.n43 43.1253
R931 B.n682 B.n681 43.1253
R932 B.t1 B.n291 38.0518
R933 B.n721 B.t0 38.0518
R934 B.n678 B.n677 36.059
R935 B.n102 B.n45 36.059
R936 B.n572 B.n571 36.059
R937 B.n565 B.n329 36.059
R938 B.t7 B.n315 27.9048
R939 B.n697 B.t3 27.9048
R940 B B.n732 18.0485
R941 B.n593 B.t7 15.221
R942 B.t3 B.n696 15.221
R943 B.n103 B.n102 10.6151
R944 B.n106 B.n103 10.6151
R945 B.n107 B.n106 10.6151
R946 B.n110 B.n107 10.6151
R947 B.n111 B.n110 10.6151
R948 B.n114 B.n111 10.6151
R949 B.n115 B.n114 10.6151
R950 B.n118 B.n115 10.6151
R951 B.n119 B.n118 10.6151
R952 B.n122 B.n119 10.6151
R953 B.n123 B.n122 10.6151
R954 B.n126 B.n123 10.6151
R955 B.n127 B.n126 10.6151
R956 B.n130 B.n127 10.6151
R957 B.n131 B.n130 10.6151
R958 B.n134 B.n131 10.6151
R959 B.n135 B.n134 10.6151
R960 B.n138 B.n135 10.6151
R961 B.n139 B.n138 10.6151
R962 B.n142 B.n139 10.6151
R963 B.n143 B.n142 10.6151
R964 B.n146 B.n143 10.6151
R965 B.n147 B.n146 10.6151
R966 B.n150 B.n147 10.6151
R967 B.n151 B.n150 10.6151
R968 B.n154 B.n151 10.6151
R969 B.n155 B.n154 10.6151
R970 B.n158 B.n155 10.6151
R971 B.n159 B.n158 10.6151
R972 B.n162 B.n159 10.6151
R973 B.n163 B.n162 10.6151
R974 B.n166 B.n163 10.6151
R975 B.n167 B.n166 10.6151
R976 B.n170 B.n167 10.6151
R977 B.n171 B.n170 10.6151
R978 B.n174 B.n171 10.6151
R979 B.n175 B.n174 10.6151
R980 B.n178 B.n175 10.6151
R981 B.n179 B.n178 10.6151
R982 B.n182 B.n179 10.6151
R983 B.n183 B.n182 10.6151
R984 B.n187 B.n186 10.6151
R985 B.n190 B.n187 10.6151
R986 B.n191 B.n190 10.6151
R987 B.n194 B.n191 10.6151
R988 B.n195 B.n194 10.6151
R989 B.n198 B.n195 10.6151
R990 B.n199 B.n198 10.6151
R991 B.n202 B.n199 10.6151
R992 B.n207 B.n204 10.6151
R993 B.n208 B.n207 10.6151
R994 B.n211 B.n208 10.6151
R995 B.n212 B.n211 10.6151
R996 B.n215 B.n212 10.6151
R997 B.n216 B.n215 10.6151
R998 B.n219 B.n216 10.6151
R999 B.n220 B.n219 10.6151
R1000 B.n223 B.n220 10.6151
R1001 B.n224 B.n223 10.6151
R1002 B.n227 B.n224 10.6151
R1003 B.n228 B.n227 10.6151
R1004 B.n231 B.n228 10.6151
R1005 B.n232 B.n231 10.6151
R1006 B.n235 B.n232 10.6151
R1007 B.n236 B.n235 10.6151
R1008 B.n239 B.n236 10.6151
R1009 B.n240 B.n239 10.6151
R1010 B.n243 B.n240 10.6151
R1011 B.n244 B.n243 10.6151
R1012 B.n247 B.n244 10.6151
R1013 B.n248 B.n247 10.6151
R1014 B.n251 B.n248 10.6151
R1015 B.n252 B.n251 10.6151
R1016 B.n255 B.n252 10.6151
R1017 B.n256 B.n255 10.6151
R1018 B.n259 B.n256 10.6151
R1019 B.n260 B.n259 10.6151
R1020 B.n263 B.n260 10.6151
R1021 B.n264 B.n263 10.6151
R1022 B.n267 B.n264 10.6151
R1023 B.n268 B.n267 10.6151
R1024 B.n271 B.n268 10.6151
R1025 B.n272 B.n271 10.6151
R1026 B.n275 B.n272 10.6151
R1027 B.n276 B.n275 10.6151
R1028 B.n279 B.n276 10.6151
R1029 B.n280 B.n279 10.6151
R1030 B.n283 B.n280 10.6151
R1031 B.n284 B.n283 10.6151
R1032 B.n678 B.n284 10.6151
R1033 B.n573 B.n572 10.6151
R1034 B.n573 B.n325 10.6151
R1035 B.n583 B.n325 10.6151
R1036 B.n584 B.n583 10.6151
R1037 B.n585 B.n584 10.6151
R1038 B.n585 B.n317 10.6151
R1039 B.n595 B.n317 10.6151
R1040 B.n596 B.n595 10.6151
R1041 B.n597 B.n596 10.6151
R1042 B.n597 B.n309 10.6151
R1043 B.n607 B.n309 10.6151
R1044 B.n608 B.n607 10.6151
R1045 B.n609 B.n608 10.6151
R1046 B.n609 B.n301 10.6151
R1047 B.n619 B.n301 10.6151
R1048 B.n620 B.n619 10.6151
R1049 B.n621 B.n620 10.6151
R1050 B.n621 B.n293 10.6151
R1051 B.n631 B.n293 10.6151
R1052 B.n632 B.n631 10.6151
R1053 B.n634 B.n632 10.6151
R1054 B.n634 B.n633 10.6151
R1055 B.n633 B.n285 10.6151
R1056 B.n645 B.n285 10.6151
R1057 B.n646 B.n645 10.6151
R1058 B.n647 B.n646 10.6151
R1059 B.n648 B.n647 10.6151
R1060 B.n650 B.n648 10.6151
R1061 B.n651 B.n650 10.6151
R1062 B.n652 B.n651 10.6151
R1063 B.n653 B.n652 10.6151
R1064 B.n655 B.n653 10.6151
R1065 B.n656 B.n655 10.6151
R1066 B.n657 B.n656 10.6151
R1067 B.n658 B.n657 10.6151
R1068 B.n660 B.n658 10.6151
R1069 B.n661 B.n660 10.6151
R1070 B.n662 B.n661 10.6151
R1071 B.n663 B.n662 10.6151
R1072 B.n665 B.n663 10.6151
R1073 B.n666 B.n665 10.6151
R1074 B.n667 B.n666 10.6151
R1075 B.n668 B.n667 10.6151
R1076 B.n670 B.n668 10.6151
R1077 B.n671 B.n670 10.6151
R1078 B.n672 B.n671 10.6151
R1079 B.n673 B.n672 10.6151
R1080 B.n675 B.n673 10.6151
R1081 B.n676 B.n675 10.6151
R1082 B.n677 B.n676 10.6151
R1083 B.n565 B.n564 10.6151
R1084 B.n564 B.n563 10.6151
R1085 B.n563 B.n562 10.6151
R1086 B.n562 B.n560 10.6151
R1087 B.n560 B.n557 10.6151
R1088 B.n557 B.n556 10.6151
R1089 B.n556 B.n553 10.6151
R1090 B.n553 B.n552 10.6151
R1091 B.n552 B.n549 10.6151
R1092 B.n549 B.n548 10.6151
R1093 B.n548 B.n545 10.6151
R1094 B.n545 B.n544 10.6151
R1095 B.n544 B.n541 10.6151
R1096 B.n541 B.n540 10.6151
R1097 B.n540 B.n537 10.6151
R1098 B.n537 B.n536 10.6151
R1099 B.n536 B.n533 10.6151
R1100 B.n533 B.n532 10.6151
R1101 B.n532 B.n529 10.6151
R1102 B.n529 B.n528 10.6151
R1103 B.n528 B.n525 10.6151
R1104 B.n525 B.n524 10.6151
R1105 B.n524 B.n521 10.6151
R1106 B.n521 B.n520 10.6151
R1107 B.n520 B.n517 10.6151
R1108 B.n517 B.n516 10.6151
R1109 B.n516 B.n513 10.6151
R1110 B.n513 B.n512 10.6151
R1111 B.n512 B.n509 10.6151
R1112 B.n509 B.n508 10.6151
R1113 B.n508 B.n505 10.6151
R1114 B.n505 B.n504 10.6151
R1115 B.n504 B.n501 10.6151
R1116 B.n501 B.n500 10.6151
R1117 B.n500 B.n497 10.6151
R1118 B.n497 B.n496 10.6151
R1119 B.n496 B.n493 10.6151
R1120 B.n493 B.n492 10.6151
R1121 B.n492 B.n489 10.6151
R1122 B.n489 B.n488 10.6151
R1123 B.n488 B.n485 10.6151
R1124 B.n483 B.n480 10.6151
R1125 B.n480 B.n479 10.6151
R1126 B.n479 B.n476 10.6151
R1127 B.n476 B.n475 10.6151
R1128 B.n475 B.n472 10.6151
R1129 B.n472 B.n471 10.6151
R1130 B.n471 B.n468 10.6151
R1131 B.n468 B.n467 10.6151
R1132 B.n464 B.n463 10.6151
R1133 B.n463 B.n460 10.6151
R1134 B.n460 B.n459 10.6151
R1135 B.n459 B.n456 10.6151
R1136 B.n456 B.n455 10.6151
R1137 B.n455 B.n452 10.6151
R1138 B.n452 B.n451 10.6151
R1139 B.n451 B.n448 10.6151
R1140 B.n448 B.n447 10.6151
R1141 B.n447 B.n444 10.6151
R1142 B.n444 B.n443 10.6151
R1143 B.n443 B.n440 10.6151
R1144 B.n440 B.n439 10.6151
R1145 B.n439 B.n436 10.6151
R1146 B.n436 B.n435 10.6151
R1147 B.n435 B.n432 10.6151
R1148 B.n432 B.n431 10.6151
R1149 B.n431 B.n428 10.6151
R1150 B.n428 B.n427 10.6151
R1151 B.n427 B.n424 10.6151
R1152 B.n424 B.n423 10.6151
R1153 B.n423 B.n420 10.6151
R1154 B.n420 B.n419 10.6151
R1155 B.n419 B.n416 10.6151
R1156 B.n416 B.n415 10.6151
R1157 B.n415 B.n412 10.6151
R1158 B.n412 B.n411 10.6151
R1159 B.n411 B.n408 10.6151
R1160 B.n408 B.n407 10.6151
R1161 B.n407 B.n404 10.6151
R1162 B.n404 B.n403 10.6151
R1163 B.n403 B.n400 10.6151
R1164 B.n400 B.n399 10.6151
R1165 B.n399 B.n396 10.6151
R1166 B.n396 B.n395 10.6151
R1167 B.n395 B.n392 10.6151
R1168 B.n392 B.n391 10.6151
R1169 B.n391 B.n388 10.6151
R1170 B.n388 B.n387 10.6151
R1171 B.n387 B.n333 10.6151
R1172 B.n571 B.n333 10.6151
R1173 B.n577 B.n329 10.6151
R1174 B.n578 B.n577 10.6151
R1175 B.n579 B.n578 10.6151
R1176 B.n579 B.n321 10.6151
R1177 B.n589 B.n321 10.6151
R1178 B.n590 B.n589 10.6151
R1179 B.n591 B.n590 10.6151
R1180 B.n591 B.n313 10.6151
R1181 B.n601 B.n313 10.6151
R1182 B.n602 B.n601 10.6151
R1183 B.n603 B.n602 10.6151
R1184 B.n603 B.n305 10.6151
R1185 B.n613 B.n305 10.6151
R1186 B.n614 B.n613 10.6151
R1187 B.n615 B.n614 10.6151
R1188 B.n615 B.n297 10.6151
R1189 B.n625 B.n297 10.6151
R1190 B.n626 B.n625 10.6151
R1191 B.n627 B.n626 10.6151
R1192 B.n627 B.n289 10.6151
R1193 B.n638 B.n289 10.6151
R1194 B.n639 B.n638 10.6151
R1195 B.n640 B.n639 10.6151
R1196 B.n640 B.n0 10.6151
R1197 B.n726 B.n1 10.6151
R1198 B.n726 B.n725 10.6151
R1199 B.n725 B.n724 10.6151
R1200 B.n724 B.n10 10.6151
R1201 B.n718 B.n10 10.6151
R1202 B.n718 B.n717 10.6151
R1203 B.n717 B.n716 10.6151
R1204 B.n716 B.n17 10.6151
R1205 B.n710 B.n17 10.6151
R1206 B.n710 B.n709 10.6151
R1207 B.n709 B.n708 10.6151
R1208 B.n708 B.n24 10.6151
R1209 B.n702 B.n24 10.6151
R1210 B.n702 B.n701 10.6151
R1211 B.n701 B.n700 10.6151
R1212 B.n700 B.n31 10.6151
R1213 B.n694 B.n31 10.6151
R1214 B.n694 B.n693 10.6151
R1215 B.n693 B.n692 10.6151
R1216 B.n692 B.n38 10.6151
R1217 B.n686 B.n38 10.6151
R1218 B.n686 B.n685 10.6151
R1219 B.n685 B.n684 10.6151
R1220 B.n684 B.n45 10.6151
R1221 B.n186 B.n100 6.5566
R1222 B.n203 B.n202 6.5566
R1223 B.n484 B.n483 6.5566
R1224 B.n467 B.n385 6.5566
R1225 B.n629 B.t1 5.07401
R1226 B.t0 B.n720 5.07401
R1227 B.n183 B.n100 4.05904
R1228 B.n204 B.n203 4.05904
R1229 B.n485 B.n484 4.05904
R1230 B.n464 B.n385 4.05904
R1231 B.n732 B.n0 2.81026
R1232 B.n732 B.n1 2.81026
R1233 VN VN.t0 206.671
R1234 VN VN.t1 162.254
R1235 VTAIL.n258 VTAIL.n198 289.615
R1236 VTAIL.n60 VTAIL.n0 289.615
R1237 VTAIL.n192 VTAIL.n132 289.615
R1238 VTAIL.n126 VTAIL.n66 289.615
R1239 VTAIL.n218 VTAIL.n217 185
R1240 VTAIL.n223 VTAIL.n222 185
R1241 VTAIL.n225 VTAIL.n224 185
R1242 VTAIL.n214 VTAIL.n213 185
R1243 VTAIL.n231 VTAIL.n230 185
R1244 VTAIL.n233 VTAIL.n232 185
R1245 VTAIL.n210 VTAIL.n209 185
R1246 VTAIL.n240 VTAIL.n239 185
R1247 VTAIL.n241 VTAIL.n208 185
R1248 VTAIL.n243 VTAIL.n242 185
R1249 VTAIL.n206 VTAIL.n205 185
R1250 VTAIL.n249 VTAIL.n248 185
R1251 VTAIL.n251 VTAIL.n250 185
R1252 VTAIL.n202 VTAIL.n201 185
R1253 VTAIL.n257 VTAIL.n256 185
R1254 VTAIL.n259 VTAIL.n258 185
R1255 VTAIL.n20 VTAIL.n19 185
R1256 VTAIL.n25 VTAIL.n24 185
R1257 VTAIL.n27 VTAIL.n26 185
R1258 VTAIL.n16 VTAIL.n15 185
R1259 VTAIL.n33 VTAIL.n32 185
R1260 VTAIL.n35 VTAIL.n34 185
R1261 VTAIL.n12 VTAIL.n11 185
R1262 VTAIL.n42 VTAIL.n41 185
R1263 VTAIL.n43 VTAIL.n10 185
R1264 VTAIL.n45 VTAIL.n44 185
R1265 VTAIL.n8 VTAIL.n7 185
R1266 VTAIL.n51 VTAIL.n50 185
R1267 VTAIL.n53 VTAIL.n52 185
R1268 VTAIL.n4 VTAIL.n3 185
R1269 VTAIL.n59 VTAIL.n58 185
R1270 VTAIL.n61 VTAIL.n60 185
R1271 VTAIL.n193 VTAIL.n192 185
R1272 VTAIL.n191 VTAIL.n190 185
R1273 VTAIL.n136 VTAIL.n135 185
R1274 VTAIL.n185 VTAIL.n184 185
R1275 VTAIL.n183 VTAIL.n182 185
R1276 VTAIL.n140 VTAIL.n139 185
R1277 VTAIL.n177 VTAIL.n176 185
R1278 VTAIL.n175 VTAIL.n142 185
R1279 VTAIL.n174 VTAIL.n173 185
R1280 VTAIL.n145 VTAIL.n143 185
R1281 VTAIL.n168 VTAIL.n167 185
R1282 VTAIL.n166 VTAIL.n165 185
R1283 VTAIL.n149 VTAIL.n148 185
R1284 VTAIL.n160 VTAIL.n159 185
R1285 VTAIL.n158 VTAIL.n157 185
R1286 VTAIL.n153 VTAIL.n152 185
R1287 VTAIL.n127 VTAIL.n126 185
R1288 VTAIL.n125 VTAIL.n124 185
R1289 VTAIL.n70 VTAIL.n69 185
R1290 VTAIL.n119 VTAIL.n118 185
R1291 VTAIL.n117 VTAIL.n116 185
R1292 VTAIL.n74 VTAIL.n73 185
R1293 VTAIL.n111 VTAIL.n110 185
R1294 VTAIL.n109 VTAIL.n76 185
R1295 VTAIL.n108 VTAIL.n107 185
R1296 VTAIL.n79 VTAIL.n77 185
R1297 VTAIL.n102 VTAIL.n101 185
R1298 VTAIL.n100 VTAIL.n99 185
R1299 VTAIL.n83 VTAIL.n82 185
R1300 VTAIL.n94 VTAIL.n93 185
R1301 VTAIL.n92 VTAIL.n91 185
R1302 VTAIL.n87 VTAIL.n86 185
R1303 VTAIL.n219 VTAIL.t3 149.524
R1304 VTAIL.n21 VTAIL.t1 149.524
R1305 VTAIL.n154 VTAIL.t0 149.524
R1306 VTAIL.n88 VTAIL.t2 149.524
R1307 VTAIL.n223 VTAIL.n217 104.615
R1308 VTAIL.n224 VTAIL.n223 104.615
R1309 VTAIL.n224 VTAIL.n213 104.615
R1310 VTAIL.n231 VTAIL.n213 104.615
R1311 VTAIL.n232 VTAIL.n231 104.615
R1312 VTAIL.n232 VTAIL.n209 104.615
R1313 VTAIL.n240 VTAIL.n209 104.615
R1314 VTAIL.n241 VTAIL.n240 104.615
R1315 VTAIL.n242 VTAIL.n241 104.615
R1316 VTAIL.n242 VTAIL.n205 104.615
R1317 VTAIL.n249 VTAIL.n205 104.615
R1318 VTAIL.n250 VTAIL.n249 104.615
R1319 VTAIL.n250 VTAIL.n201 104.615
R1320 VTAIL.n257 VTAIL.n201 104.615
R1321 VTAIL.n258 VTAIL.n257 104.615
R1322 VTAIL.n25 VTAIL.n19 104.615
R1323 VTAIL.n26 VTAIL.n25 104.615
R1324 VTAIL.n26 VTAIL.n15 104.615
R1325 VTAIL.n33 VTAIL.n15 104.615
R1326 VTAIL.n34 VTAIL.n33 104.615
R1327 VTAIL.n34 VTAIL.n11 104.615
R1328 VTAIL.n42 VTAIL.n11 104.615
R1329 VTAIL.n43 VTAIL.n42 104.615
R1330 VTAIL.n44 VTAIL.n43 104.615
R1331 VTAIL.n44 VTAIL.n7 104.615
R1332 VTAIL.n51 VTAIL.n7 104.615
R1333 VTAIL.n52 VTAIL.n51 104.615
R1334 VTAIL.n52 VTAIL.n3 104.615
R1335 VTAIL.n59 VTAIL.n3 104.615
R1336 VTAIL.n60 VTAIL.n59 104.615
R1337 VTAIL.n192 VTAIL.n191 104.615
R1338 VTAIL.n191 VTAIL.n135 104.615
R1339 VTAIL.n184 VTAIL.n135 104.615
R1340 VTAIL.n184 VTAIL.n183 104.615
R1341 VTAIL.n183 VTAIL.n139 104.615
R1342 VTAIL.n176 VTAIL.n139 104.615
R1343 VTAIL.n176 VTAIL.n175 104.615
R1344 VTAIL.n175 VTAIL.n174 104.615
R1345 VTAIL.n174 VTAIL.n143 104.615
R1346 VTAIL.n167 VTAIL.n143 104.615
R1347 VTAIL.n167 VTAIL.n166 104.615
R1348 VTAIL.n166 VTAIL.n148 104.615
R1349 VTAIL.n159 VTAIL.n148 104.615
R1350 VTAIL.n159 VTAIL.n158 104.615
R1351 VTAIL.n158 VTAIL.n152 104.615
R1352 VTAIL.n126 VTAIL.n125 104.615
R1353 VTAIL.n125 VTAIL.n69 104.615
R1354 VTAIL.n118 VTAIL.n69 104.615
R1355 VTAIL.n118 VTAIL.n117 104.615
R1356 VTAIL.n117 VTAIL.n73 104.615
R1357 VTAIL.n110 VTAIL.n73 104.615
R1358 VTAIL.n110 VTAIL.n109 104.615
R1359 VTAIL.n109 VTAIL.n108 104.615
R1360 VTAIL.n108 VTAIL.n77 104.615
R1361 VTAIL.n101 VTAIL.n77 104.615
R1362 VTAIL.n101 VTAIL.n100 104.615
R1363 VTAIL.n100 VTAIL.n82 104.615
R1364 VTAIL.n93 VTAIL.n82 104.615
R1365 VTAIL.n93 VTAIL.n92 104.615
R1366 VTAIL.n92 VTAIL.n86 104.615
R1367 VTAIL.t3 VTAIL.n217 52.3082
R1368 VTAIL.t1 VTAIL.n19 52.3082
R1369 VTAIL.t0 VTAIL.n152 52.3082
R1370 VTAIL.t2 VTAIL.n86 52.3082
R1371 VTAIL.n263 VTAIL.n262 31.2157
R1372 VTAIL.n65 VTAIL.n64 31.2157
R1373 VTAIL.n197 VTAIL.n196 31.2157
R1374 VTAIL.n131 VTAIL.n130 31.2157
R1375 VTAIL.n131 VTAIL.n65 27.7893
R1376 VTAIL.n263 VTAIL.n197 25.2807
R1377 VTAIL.n243 VTAIL.n208 13.1884
R1378 VTAIL.n45 VTAIL.n10 13.1884
R1379 VTAIL.n177 VTAIL.n142 13.1884
R1380 VTAIL.n111 VTAIL.n76 13.1884
R1381 VTAIL.n239 VTAIL.n238 12.8005
R1382 VTAIL.n244 VTAIL.n206 12.8005
R1383 VTAIL.n41 VTAIL.n40 12.8005
R1384 VTAIL.n46 VTAIL.n8 12.8005
R1385 VTAIL.n178 VTAIL.n140 12.8005
R1386 VTAIL.n173 VTAIL.n144 12.8005
R1387 VTAIL.n112 VTAIL.n74 12.8005
R1388 VTAIL.n107 VTAIL.n78 12.8005
R1389 VTAIL.n237 VTAIL.n210 12.0247
R1390 VTAIL.n248 VTAIL.n247 12.0247
R1391 VTAIL.n39 VTAIL.n12 12.0247
R1392 VTAIL.n50 VTAIL.n49 12.0247
R1393 VTAIL.n182 VTAIL.n181 12.0247
R1394 VTAIL.n172 VTAIL.n145 12.0247
R1395 VTAIL.n116 VTAIL.n115 12.0247
R1396 VTAIL.n106 VTAIL.n79 12.0247
R1397 VTAIL.n234 VTAIL.n233 11.249
R1398 VTAIL.n251 VTAIL.n204 11.249
R1399 VTAIL.n36 VTAIL.n35 11.249
R1400 VTAIL.n53 VTAIL.n6 11.249
R1401 VTAIL.n185 VTAIL.n138 11.249
R1402 VTAIL.n169 VTAIL.n168 11.249
R1403 VTAIL.n119 VTAIL.n72 11.249
R1404 VTAIL.n103 VTAIL.n102 11.249
R1405 VTAIL.n230 VTAIL.n212 10.4732
R1406 VTAIL.n252 VTAIL.n202 10.4732
R1407 VTAIL.n32 VTAIL.n14 10.4732
R1408 VTAIL.n54 VTAIL.n4 10.4732
R1409 VTAIL.n186 VTAIL.n136 10.4732
R1410 VTAIL.n165 VTAIL.n147 10.4732
R1411 VTAIL.n120 VTAIL.n70 10.4732
R1412 VTAIL.n99 VTAIL.n81 10.4732
R1413 VTAIL.n219 VTAIL.n218 10.2747
R1414 VTAIL.n21 VTAIL.n20 10.2747
R1415 VTAIL.n154 VTAIL.n153 10.2747
R1416 VTAIL.n88 VTAIL.n87 10.2747
R1417 VTAIL.n229 VTAIL.n214 9.69747
R1418 VTAIL.n256 VTAIL.n255 9.69747
R1419 VTAIL.n31 VTAIL.n16 9.69747
R1420 VTAIL.n58 VTAIL.n57 9.69747
R1421 VTAIL.n190 VTAIL.n189 9.69747
R1422 VTAIL.n164 VTAIL.n149 9.69747
R1423 VTAIL.n124 VTAIL.n123 9.69747
R1424 VTAIL.n98 VTAIL.n83 9.69747
R1425 VTAIL.n262 VTAIL.n261 9.45567
R1426 VTAIL.n64 VTAIL.n63 9.45567
R1427 VTAIL.n196 VTAIL.n195 9.45567
R1428 VTAIL.n130 VTAIL.n129 9.45567
R1429 VTAIL.n261 VTAIL.n260 9.3005
R1430 VTAIL.n200 VTAIL.n199 9.3005
R1431 VTAIL.n255 VTAIL.n254 9.3005
R1432 VTAIL.n253 VTAIL.n252 9.3005
R1433 VTAIL.n204 VTAIL.n203 9.3005
R1434 VTAIL.n247 VTAIL.n246 9.3005
R1435 VTAIL.n245 VTAIL.n244 9.3005
R1436 VTAIL.n221 VTAIL.n220 9.3005
R1437 VTAIL.n216 VTAIL.n215 9.3005
R1438 VTAIL.n227 VTAIL.n226 9.3005
R1439 VTAIL.n229 VTAIL.n228 9.3005
R1440 VTAIL.n212 VTAIL.n211 9.3005
R1441 VTAIL.n235 VTAIL.n234 9.3005
R1442 VTAIL.n237 VTAIL.n236 9.3005
R1443 VTAIL.n238 VTAIL.n207 9.3005
R1444 VTAIL.n63 VTAIL.n62 9.3005
R1445 VTAIL.n2 VTAIL.n1 9.3005
R1446 VTAIL.n57 VTAIL.n56 9.3005
R1447 VTAIL.n55 VTAIL.n54 9.3005
R1448 VTAIL.n6 VTAIL.n5 9.3005
R1449 VTAIL.n49 VTAIL.n48 9.3005
R1450 VTAIL.n47 VTAIL.n46 9.3005
R1451 VTAIL.n23 VTAIL.n22 9.3005
R1452 VTAIL.n18 VTAIL.n17 9.3005
R1453 VTAIL.n29 VTAIL.n28 9.3005
R1454 VTAIL.n31 VTAIL.n30 9.3005
R1455 VTAIL.n14 VTAIL.n13 9.3005
R1456 VTAIL.n37 VTAIL.n36 9.3005
R1457 VTAIL.n39 VTAIL.n38 9.3005
R1458 VTAIL.n40 VTAIL.n9 9.3005
R1459 VTAIL.n156 VTAIL.n155 9.3005
R1460 VTAIL.n151 VTAIL.n150 9.3005
R1461 VTAIL.n162 VTAIL.n161 9.3005
R1462 VTAIL.n164 VTAIL.n163 9.3005
R1463 VTAIL.n147 VTAIL.n146 9.3005
R1464 VTAIL.n170 VTAIL.n169 9.3005
R1465 VTAIL.n172 VTAIL.n171 9.3005
R1466 VTAIL.n144 VTAIL.n141 9.3005
R1467 VTAIL.n195 VTAIL.n194 9.3005
R1468 VTAIL.n134 VTAIL.n133 9.3005
R1469 VTAIL.n189 VTAIL.n188 9.3005
R1470 VTAIL.n187 VTAIL.n186 9.3005
R1471 VTAIL.n138 VTAIL.n137 9.3005
R1472 VTAIL.n181 VTAIL.n180 9.3005
R1473 VTAIL.n179 VTAIL.n178 9.3005
R1474 VTAIL.n90 VTAIL.n89 9.3005
R1475 VTAIL.n85 VTAIL.n84 9.3005
R1476 VTAIL.n96 VTAIL.n95 9.3005
R1477 VTAIL.n98 VTAIL.n97 9.3005
R1478 VTAIL.n81 VTAIL.n80 9.3005
R1479 VTAIL.n104 VTAIL.n103 9.3005
R1480 VTAIL.n106 VTAIL.n105 9.3005
R1481 VTAIL.n78 VTAIL.n75 9.3005
R1482 VTAIL.n129 VTAIL.n128 9.3005
R1483 VTAIL.n68 VTAIL.n67 9.3005
R1484 VTAIL.n123 VTAIL.n122 9.3005
R1485 VTAIL.n121 VTAIL.n120 9.3005
R1486 VTAIL.n72 VTAIL.n71 9.3005
R1487 VTAIL.n115 VTAIL.n114 9.3005
R1488 VTAIL.n113 VTAIL.n112 9.3005
R1489 VTAIL.n226 VTAIL.n225 8.92171
R1490 VTAIL.n259 VTAIL.n200 8.92171
R1491 VTAIL.n28 VTAIL.n27 8.92171
R1492 VTAIL.n61 VTAIL.n2 8.92171
R1493 VTAIL.n193 VTAIL.n134 8.92171
R1494 VTAIL.n161 VTAIL.n160 8.92171
R1495 VTAIL.n127 VTAIL.n68 8.92171
R1496 VTAIL.n95 VTAIL.n94 8.92171
R1497 VTAIL.n222 VTAIL.n216 8.14595
R1498 VTAIL.n260 VTAIL.n198 8.14595
R1499 VTAIL.n24 VTAIL.n18 8.14595
R1500 VTAIL.n62 VTAIL.n0 8.14595
R1501 VTAIL.n194 VTAIL.n132 8.14595
R1502 VTAIL.n157 VTAIL.n151 8.14595
R1503 VTAIL.n128 VTAIL.n66 8.14595
R1504 VTAIL.n91 VTAIL.n85 8.14595
R1505 VTAIL.n221 VTAIL.n218 7.3702
R1506 VTAIL.n23 VTAIL.n20 7.3702
R1507 VTAIL.n156 VTAIL.n153 7.3702
R1508 VTAIL.n90 VTAIL.n87 7.3702
R1509 VTAIL.n222 VTAIL.n221 5.81868
R1510 VTAIL.n262 VTAIL.n198 5.81868
R1511 VTAIL.n24 VTAIL.n23 5.81868
R1512 VTAIL.n64 VTAIL.n0 5.81868
R1513 VTAIL.n196 VTAIL.n132 5.81868
R1514 VTAIL.n157 VTAIL.n156 5.81868
R1515 VTAIL.n130 VTAIL.n66 5.81868
R1516 VTAIL.n91 VTAIL.n90 5.81868
R1517 VTAIL.n225 VTAIL.n216 5.04292
R1518 VTAIL.n260 VTAIL.n259 5.04292
R1519 VTAIL.n27 VTAIL.n18 5.04292
R1520 VTAIL.n62 VTAIL.n61 5.04292
R1521 VTAIL.n194 VTAIL.n193 5.04292
R1522 VTAIL.n160 VTAIL.n151 5.04292
R1523 VTAIL.n128 VTAIL.n127 5.04292
R1524 VTAIL.n94 VTAIL.n85 5.04292
R1525 VTAIL.n226 VTAIL.n214 4.26717
R1526 VTAIL.n256 VTAIL.n200 4.26717
R1527 VTAIL.n28 VTAIL.n16 4.26717
R1528 VTAIL.n58 VTAIL.n2 4.26717
R1529 VTAIL.n190 VTAIL.n134 4.26717
R1530 VTAIL.n161 VTAIL.n149 4.26717
R1531 VTAIL.n124 VTAIL.n68 4.26717
R1532 VTAIL.n95 VTAIL.n83 4.26717
R1533 VTAIL.n230 VTAIL.n229 3.49141
R1534 VTAIL.n255 VTAIL.n202 3.49141
R1535 VTAIL.n32 VTAIL.n31 3.49141
R1536 VTAIL.n57 VTAIL.n4 3.49141
R1537 VTAIL.n189 VTAIL.n136 3.49141
R1538 VTAIL.n165 VTAIL.n164 3.49141
R1539 VTAIL.n123 VTAIL.n70 3.49141
R1540 VTAIL.n99 VTAIL.n98 3.49141
R1541 VTAIL.n220 VTAIL.n219 2.84303
R1542 VTAIL.n22 VTAIL.n21 2.84303
R1543 VTAIL.n155 VTAIL.n154 2.84303
R1544 VTAIL.n89 VTAIL.n88 2.84303
R1545 VTAIL.n233 VTAIL.n212 2.71565
R1546 VTAIL.n252 VTAIL.n251 2.71565
R1547 VTAIL.n35 VTAIL.n14 2.71565
R1548 VTAIL.n54 VTAIL.n53 2.71565
R1549 VTAIL.n186 VTAIL.n185 2.71565
R1550 VTAIL.n168 VTAIL.n147 2.71565
R1551 VTAIL.n120 VTAIL.n119 2.71565
R1552 VTAIL.n102 VTAIL.n81 2.71565
R1553 VTAIL.n234 VTAIL.n210 1.93989
R1554 VTAIL.n248 VTAIL.n204 1.93989
R1555 VTAIL.n36 VTAIL.n12 1.93989
R1556 VTAIL.n50 VTAIL.n6 1.93989
R1557 VTAIL.n182 VTAIL.n138 1.93989
R1558 VTAIL.n169 VTAIL.n145 1.93989
R1559 VTAIL.n116 VTAIL.n72 1.93989
R1560 VTAIL.n103 VTAIL.n79 1.93989
R1561 VTAIL.n197 VTAIL.n131 1.72464
R1562 VTAIL.n239 VTAIL.n237 1.16414
R1563 VTAIL.n247 VTAIL.n206 1.16414
R1564 VTAIL.n41 VTAIL.n39 1.16414
R1565 VTAIL.n49 VTAIL.n8 1.16414
R1566 VTAIL.n181 VTAIL.n140 1.16414
R1567 VTAIL.n173 VTAIL.n172 1.16414
R1568 VTAIL.n115 VTAIL.n74 1.16414
R1569 VTAIL.n107 VTAIL.n106 1.16414
R1570 VTAIL VTAIL.n65 1.15567
R1571 VTAIL VTAIL.n263 0.569465
R1572 VTAIL.n238 VTAIL.n208 0.388379
R1573 VTAIL.n244 VTAIL.n243 0.388379
R1574 VTAIL.n40 VTAIL.n10 0.388379
R1575 VTAIL.n46 VTAIL.n45 0.388379
R1576 VTAIL.n178 VTAIL.n177 0.388379
R1577 VTAIL.n144 VTAIL.n142 0.388379
R1578 VTAIL.n112 VTAIL.n111 0.388379
R1579 VTAIL.n78 VTAIL.n76 0.388379
R1580 VTAIL.n220 VTAIL.n215 0.155672
R1581 VTAIL.n227 VTAIL.n215 0.155672
R1582 VTAIL.n228 VTAIL.n227 0.155672
R1583 VTAIL.n228 VTAIL.n211 0.155672
R1584 VTAIL.n235 VTAIL.n211 0.155672
R1585 VTAIL.n236 VTAIL.n235 0.155672
R1586 VTAIL.n236 VTAIL.n207 0.155672
R1587 VTAIL.n245 VTAIL.n207 0.155672
R1588 VTAIL.n246 VTAIL.n245 0.155672
R1589 VTAIL.n246 VTAIL.n203 0.155672
R1590 VTAIL.n253 VTAIL.n203 0.155672
R1591 VTAIL.n254 VTAIL.n253 0.155672
R1592 VTAIL.n254 VTAIL.n199 0.155672
R1593 VTAIL.n261 VTAIL.n199 0.155672
R1594 VTAIL.n22 VTAIL.n17 0.155672
R1595 VTAIL.n29 VTAIL.n17 0.155672
R1596 VTAIL.n30 VTAIL.n29 0.155672
R1597 VTAIL.n30 VTAIL.n13 0.155672
R1598 VTAIL.n37 VTAIL.n13 0.155672
R1599 VTAIL.n38 VTAIL.n37 0.155672
R1600 VTAIL.n38 VTAIL.n9 0.155672
R1601 VTAIL.n47 VTAIL.n9 0.155672
R1602 VTAIL.n48 VTAIL.n47 0.155672
R1603 VTAIL.n48 VTAIL.n5 0.155672
R1604 VTAIL.n55 VTAIL.n5 0.155672
R1605 VTAIL.n56 VTAIL.n55 0.155672
R1606 VTAIL.n56 VTAIL.n1 0.155672
R1607 VTAIL.n63 VTAIL.n1 0.155672
R1608 VTAIL.n195 VTAIL.n133 0.155672
R1609 VTAIL.n188 VTAIL.n133 0.155672
R1610 VTAIL.n188 VTAIL.n187 0.155672
R1611 VTAIL.n187 VTAIL.n137 0.155672
R1612 VTAIL.n180 VTAIL.n137 0.155672
R1613 VTAIL.n180 VTAIL.n179 0.155672
R1614 VTAIL.n179 VTAIL.n141 0.155672
R1615 VTAIL.n171 VTAIL.n141 0.155672
R1616 VTAIL.n171 VTAIL.n170 0.155672
R1617 VTAIL.n170 VTAIL.n146 0.155672
R1618 VTAIL.n163 VTAIL.n146 0.155672
R1619 VTAIL.n163 VTAIL.n162 0.155672
R1620 VTAIL.n162 VTAIL.n150 0.155672
R1621 VTAIL.n155 VTAIL.n150 0.155672
R1622 VTAIL.n129 VTAIL.n67 0.155672
R1623 VTAIL.n122 VTAIL.n67 0.155672
R1624 VTAIL.n122 VTAIL.n121 0.155672
R1625 VTAIL.n121 VTAIL.n71 0.155672
R1626 VTAIL.n114 VTAIL.n71 0.155672
R1627 VTAIL.n114 VTAIL.n113 0.155672
R1628 VTAIL.n113 VTAIL.n75 0.155672
R1629 VTAIL.n105 VTAIL.n75 0.155672
R1630 VTAIL.n105 VTAIL.n104 0.155672
R1631 VTAIL.n104 VTAIL.n80 0.155672
R1632 VTAIL.n97 VTAIL.n80 0.155672
R1633 VTAIL.n97 VTAIL.n96 0.155672
R1634 VTAIL.n96 VTAIL.n84 0.155672
R1635 VTAIL.n89 VTAIL.n84 0.155672
R1636 VDD2.n125 VDD2.n65 289.615
R1637 VDD2.n60 VDD2.n0 289.615
R1638 VDD2.n126 VDD2.n125 185
R1639 VDD2.n124 VDD2.n123 185
R1640 VDD2.n69 VDD2.n68 185
R1641 VDD2.n118 VDD2.n117 185
R1642 VDD2.n116 VDD2.n115 185
R1643 VDD2.n73 VDD2.n72 185
R1644 VDD2.n110 VDD2.n109 185
R1645 VDD2.n108 VDD2.n75 185
R1646 VDD2.n107 VDD2.n106 185
R1647 VDD2.n78 VDD2.n76 185
R1648 VDD2.n101 VDD2.n100 185
R1649 VDD2.n99 VDD2.n98 185
R1650 VDD2.n82 VDD2.n81 185
R1651 VDD2.n93 VDD2.n92 185
R1652 VDD2.n91 VDD2.n90 185
R1653 VDD2.n86 VDD2.n85 185
R1654 VDD2.n20 VDD2.n19 185
R1655 VDD2.n25 VDD2.n24 185
R1656 VDD2.n27 VDD2.n26 185
R1657 VDD2.n16 VDD2.n15 185
R1658 VDD2.n33 VDD2.n32 185
R1659 VDD2.n35 VDD2.n34 185
R1660 VDD2.n12 VDD2.n11 185
R1661 VDD2.n42 VDD2.n41 185
R1662 VDD2.n43 VDD2.n10 185
R1663 VDD2.n45 VDD2.n44 185
R1664 VDD2.n8 VDD2.n7 185
R1665 VDD2.n51 VDD2.n50 185
R1666 VDD2.n53 VDD2.n52 185
R1667 VDD2.n4 VDD2.n3 185
R1668 VDD2.n59 VDD2.n58 185
R1669 VDD2.n61 VDD2.n60 185
R1670 VDD2.n87 VDD2.t1 149.524
R1671 VDD2.n21 VDD2.t0 149.524
R1672 VDD2.n125 VDD2.n124 104.615
R1673 VDD2.n124 VDD2.n68 104.615
R1674 VDD2.n117 VDD2.n68 104.615
R1675 VDD2.n117 VDD2.n116 104.615
R1676 VDD2.n116 VDD2.n72 104.615
R1677 VDD2.n109 VDD2.n72 104.615
R1678 VDD2.n109 VDD2.n108 104.615
R1679 VDD2.n108 VDD2.n107 104.615
R1680 VDD2.n107 VDD2.n76 104.615
R1681 VDD2.n100 VDD2.n76 104.615
R1682 VDD2.n100 VDD2.n99 104.615
R1683 VDD2.n99 VDD2.n81 104.615
R1684 VDD2.n92 VDD2.n81 104.615
R1685 VDD2.n92 VDD2.n91 104.615
R1686 VDD2.n91 VDD2.n85 104.615
R1687 VDD2.n25 VDD2.n19 104.615
R1688 VDD2.n26 VDD2.n25 104.615
R1689 VDD2.n26 VDD2.n15 104.615
R1690 VDD2.n33 VDD2.n15 104.615
R1691 VDD2.n34 VDD2.n33 104.615
R1692 VDD2.n34 VDD2.n11 104.615
R1693 VDD2.n42 VDD2.n11 104.615
R1694 VDD2.n43 VDD2.n42 104.615
R1695 VDD2.n44 VDD2.n43 104.615
R1696 VDD2.n44 VDD2.n7 104.615
R1697 VDD2.n51 VDD2.n7 104.615
R1698 VDD2.n52 VDD2.n51 104.615
R1699 VDD2.n52 VDD2.n3 104.615
R1700 VDD2.n59 VDD2.n3 104.615
R1701 VDD2.n60 VDD2.n59 104.615
R1702 VDD2.n130 VDD2.n64 86.9763
R1703 VDD2.t1 VDD2.n85 52.3082
R1704 VDD2.t0 VDD2.n19 52.3082
R1705 VDD2.n130 VDD2.n129 47.8944
R1706 VDD2.n110 VDD2.n75 13.1884
R1707 VDD2.n45 VDD2.n10 13.1884
R1708 VDD2.n111 VDD2.n73 12.8005
R1709 VDD2.n106 VDD2.n77 12.8005
R1710 VDD2.n41 VDD2.n40 12.8005
R1711 VDD2.n46 VDD2.n8 12.8005
R1712 VDD2.n115 VDD2.n114 12.0247
R1713 VDD2.n105 VDD2.n78 12.0247
R1714 VDD2.n39 VDD2.n12 12.0247
R1715 VDD2.n50 VDD2.n49 12.0247
R1716 VDD2.n118 VDD2.n71 11.249
R1717 VDD2.n102 VDD2.n101 11.249
R1718 VDD2.n36 VDD2.n35 11.249
R1719 VDD2.n53 VDD2.n6 11.249
R1720 VDD2.n119 VDD2.n69 10.4732
R1721 VDD2.n98 VDD2.n80 10.4732
R1722 VDD2.n32 VDD2.n14 10.4732
R1723 VDD2.n54 VDD2.n4 10.4732
R1724 VDD2.n87 VDD2.n86 10.2747
R1725 VDD2.n21 VDD2.n20 10.2747
R1726 VDD2.n123 VDD2.n122 9.69747
R1727 VDD2.n97 VDD2.n82 9.69747
R1728 VDD2.n31 VDD2.n16 9.69747
R1729 VDD2.n58 VDD2.n57 9.69747
R1730 VDD2.n129 VDD2.n128 9.45567
R1731 VDD2.n64 VDD2.n63 9.45567
R1732 VDD2.n89 VDD2.n88 9.3005
R1733 VDD2.n84 VDD2.n83 9.3005
R1734 VDD2.n95 VDD2.n94 9.3005
R1735 VDD2.n97 VDD2.n96 9.3005
R1736 VDD2.n80 VDD2.n79 9.3005
R1737 VDD2.n103 VDD2.n102 9.3005
R1738 VDD2.n105 VDD2.n104 9.3005
R1739 VDD2.n77 VDD2.n74 9.3005
R1740 VDD2.n128 VDD2.n127 9.3005
R1741 VDD2.n67 VDD2.n66 9.3005
R1742 VDD2.n122 VDD2.n121 9.3005
R1743 VDD2.n120 VDD2.n119 9.3005
R1744 VDD2.n71 VDD2.n70 9.3005
R1745 VDD2.n114 VDD2.n113 9.3005
R1746 VDD2.n112 VDD2.n111 9.3005
R1747 VDD2.n63 VDD2.n62 9.3005
R1748 VDD2.n2 VDD2.n1 9.3005
R1749 VDD2.n57 VDD2.n56 9.3005
R1750 VDD2.n55 VDD2.n54 9.3005
R1751 VDD2.n6 VDD2.n5 9.3005
R1752 VDD2.n49 VDD2.n48 9.3005
R1753 VDD2.n47 VDD2.n46 9.3005
R1754 VDD2.n23 VDD2.n22 9.3005
R1755 VDD2.n18 VDD2.n17 9.3005
R1756 VDD2.n29 VDD2.n28 9.3005
R1757 VDD2.n31 VDD2.n30 9.3005
R1758 VDD2.n14 VDD2.n13 9.3005
R1759 VDD2.n37 VDD2.n36 9.3005
R1760 VDD2.n39 VDD2.n38 9.3005
R1761 VDD2.n40 VDD2.n9 9.3005
R1762 VDD2.n126 VDD2.n67 8.92171
R1763 VDD2.n94 VDD2.n93 8.92171
R1764 VDD2.n28 VDD2.n27 8.92171
R1765 VDD2.n61 VDD2.n2 8.92171
R1766 VDD2.n127 VDD2.n65 8.14595
R1767 VDD2.n90 VDD2.n84 8.14595
R1768 VDD2.n24 VDD2.n18 8.14595
R1769 VDD2.n62 VDD2.n0 8.14595
R1770 VDD2.n89 VDD2.n86 7.3702
R1771 VDD2.n23 VDD2.n20 7.3702
R1772 VDD2.n129 VDD2.n65 5.81868
R1773 VDD2.n90 VDD2.n89 5.81868
R1774 VDD2.n24 VDD2.n23 5.81868
R1775 VDD2.n64 VDD2.n0 5.81868
R1776 VDD2.n127 VDD2.n126 5.04292
R1777 VDD2.n93 VDD2.n84 5.04292
R1778 VDD2.n27 VDD2.n18 5.04292
R1779 VDD2.n62 VDD2.n61 5.04292
R1780 VDD2.n123 VDD2.n67 4.26717
R1781 VDD2.n94 VDD2.n82 4.26717
R1782 VDD2.n28 VDD2.n16 4.26717
R1783 VDD2.n58 VDD2.n2 4.26717
R1784 VDD2.n122 VDD2.n69 3.49141
R1785 VDD2.n98 VDD2.n97 3.49141
R1786 VDD2.n32 VDD2.n31 3.49141
R1787 VDD2.n57 VDD2.n4 3.49141
R1788 VDD2.n88 VDD2.n87 2.84303
R1789 VDD2.n22 VDD2.n21 2.84303
R1790 VDD2.n119 VDD2.n118 2.71565
R1791 VDD2.n101 VDD2.n80 2.71565
R1792 VDD2.n35 VDD2.n14 2.71565
R1793 VDD2.n54 VDD2.n53 2.71565
R1794 VDD2.n115 VDD2.n71 1.93989
R1795 VDD2.n102 VDD2.n78 1.93989
R1796 VDD2.n36 VDD2.n12 1.93989
R1797 VDD2.n50 VDD2.n6 1.93989
R1798 VDD2.n114 VDD2.n73 1.16414
R1799 VDD2.n106 VDD2.n105 1.16414
R1800 VDD2.n41 VDD2.n39 1.16414
R1801 VDD2.n49 VDD2.n8 1.16414
R1802 VDD2 VDD2.n130 0.685845
R1803 VDD2.n111 VDD2.n110 0.388379
R1804 VDD2.n77 VDD2.n75 0.388379
R1805 VDD2.n40 VDD2.n10 0.388379
R1806 VDD2.n46 VDD2.n45 0.388379
R1807 VDD2.n128 VDD2.n66 0.155672
R1808 VDD2.n121 VDD2.n66 0.155672
R1809 VDD2.n121 VDD2.n120 0.155672
R1810 VDD2.n120 VDD2.n70 0.155672
R1811 VDD2.n113 VDD2.n70 0.155672
R1812 VDD2.n113 VDD2.n112 0.155672
R1813 VDD2.n112 VDD2.n74 0.155672
R1814 VDD2.n104 VDD2.n74 0.155672
R1815 VDD2.n104 VDD2.n103 0.155672
R1816 VDD2.n103 VDD2.n79 0.155672
R1817 VDD2.n96 VDD2.n79 0.155672
R1818 VDD2.n96 VDD2.n95 0.155672
R1819 VDD2.n95 VDD2.n83 0.155672
R1820 VDD2.n88 VDD2.n83 0.155672
R1821 VDD2.n22 VDD2.n17 0.155672
R1822 VDD2.n29 VDD2.n17 0.155672
R1823 VDD2.n30 VDD2.n29 0.155672
R1824 VDD2.n30 VDD2.n13 0.155672
R1825 VDD2.n37 VDD2.n13 0.155672
R1826 VDD2.n38 VDD2.n37 0.155672
R1827 VDD2.n38 VDD2.n9 0.155672
R1828 VDD2.n47 VDD2.n9 0.155672
R1829 VDD2.n48 VDD2.n47 0.155672
R1830 VDD2.n48 VDD2.n5 0.155672
R1831 VDD2.n55 VDD2.n5 0.155672
R1832 VDD2.n56 VDD2.n55 0.155672
R1833 VDD2.n56 VDD2.n1 0.155672
R1834 VDD2.n63 VDD2.n1 0.155672
R1835 VP.n0 VP.t0 206.575
R1836 VP.n0 VP.t1 161.917
R1837 VP VP.n0 0.336784
R1838 VDD1.n60 VDD1.n0 289.615
R1839 VDD1.n125 VDD1.n65 289.615
R1840 VDD1.n61 VDD1.n60 185
R1841 VDD1.n59 VDD1.n58 185
R1842 VDD1.n4 VDD1.n3 185
R1843 VDD1.n53 VDD1.n52 185
R1844 VDD1.n51 VDD1.n50 185
R1845 VDD1.n8 VDD1.n7 185
R1846 VDD1.n45 VDD1.n44 185
R1847 VDD1.n43 VDD1.n10 185
R1848 VDD1.n42 VDD1.n41 185
R1849 VDD1.n13 VDD1.n11 185
R1850 VDD1.n36 VDD1.n35 185
R1851 VDD1.n34 VDD1.n33 185
R1852 VDD1.n17 VDD1.n16 185
R1853 VDD1.n28 VDD1.n27 185
R1854 VDD1.n26 VDD1.n25 185
R1855 VDD1.n21 VDD1.n20 185
R1856 VDD1.n85 VDD1.n84 185
R1857 VDD1.n90 VDD1.n89 185
R1858 VDD1.n92 VDD1.n91 185
R1859 VDD1.n81 VDD1.n80 185
R1860 VDD1.n98 VDD1.n97 185
R1861 VDD1.n100 VDD1.n99 185
R1862 VDD1.n77 VDD1.n76 185
R1863 VDD1.n107 VDD1.n106 185
R1864 VDD1.n108 VDD1.n75 185
R1865 VDD1.n110 VDD1.n109 185
R1866 VDD1.n73 VDD1.n72 185
R1867 VDD1.n116 VDD1.n115 185
R1868 VDD1.n118 VDD1.n117 185
R1869 VDD1.n69 VDD1.n68 185
R1870 VDD1.n124 VDD1.n123 185
R1871 VDD1.n126 VDD1.n125 185
R1872 VDD1.n22 VDD1.t1 149.524
R1873 VDD1.n86 VDD1.t0 149.524
R1874 VDD1.n60 VDD1.n59 104.615
R1875 VDD1.n59 VDD1.n3 104.615
R1876 VDD1.n52 VDD1.n3 104.615
R1877 VDD1.n52 VDD1.n51 104.615
R1878 VDD1.n51 VDD1.n7 104.615
R1879 VDD1.n44 VDD1.n7 104.615
R1880 VDD1.n44 VDD1.n43 104.615
R1881 VDD1.n43 VDD1.n42 104.615
R1882 VDD1.n42 VDD1.n11 104.615
R1883 VDD1.n35 VDD1.n11 104.615
R1884 VDD1.n35 VDD1.n34 104.615
R1885 VDD1.n34 VDD1.n16 104.615
R1886 VDD1.n27 VDD1.n16 104.615
R1887 VDD1.n27 VDD1.n26 104.615
R1888 VDD1.n26 VDD1.n20 104.615
R1889 VDD1.n90 VDD1.n84 104.615
R1890 VDD1.n91 VDD1.n90 104.615
R1891 VDD1.n91 VDD1.n80 104.615
R1892 VDD1.n98 VDD1.n80 104.615
R1893 VDD1.n99 VDD1.n98 104.615
R1894 VDD1.n99 VDD1.n76 104.615
R1895 VDD1.n107 VDD1.n76 104.615
R1896 VDD1.n108 VDD1.n107 104.615
R1897 VDD1.n109 VDD1.n108 104.615
R1898 VDD1.n109 VDD1.n72 104.615
R1899 VDD1.n116 VDD1.n72 104.615
R1900 VDD1.n117 VDD1.n116 104.615
R1901 VDD1.n117 VDD1.n68 104.615
R1902 VDD1.n124 VDD1.n68 104.615
R1903 VDD1.n125 VDD1.n124 104.615
R1904 VDD1 VDD1.n129 88.1283
R1905 VDD1.t1 VDD1.n20 52.3082
R1906 VDD1.t0 VDD1.n84 52.3082
R1907 VDD1 VDD1.n64 48.5798
R1908 VDD1.n45 VDD1.n10 13.1884
R1909 VDD1.n110 VDD1.n75 13.1884
R1910 VDD1.n46 VDD1.n8 12.8005
R1911 VDD1.n41 VDD1.n12 12.8005
R1912 VDD1.n106 VDD1.n105 12.8005
R1913 VDD1.n111 VDD1.n73 12.8005
R1914 VDD1.n50 VDD1.n49 12.0247
R1915 VDD1.n40 VDD1.n13 12.0247
R1916 VDD1.n104 VDD1.n77 12.0247
R1917 VDD1.n115 VDD1.n114 12.0247
R1918 VDD1.n53 VDD1.n6 11.249
R1919 VDD1.n37 VDD1.n36 11.249
R1920 VDD1.n101 VDD1.n100 11.249
R1921 VDD1.n118 VDD1.n71 11.249
R1922 VDD1.n54 VDD1.n4 10.4732
R1923 VDD1.n33 VDD1.n15 10.4732
R1924 VDD1.n97 VDD1.n79 10.4732
R1925 VDD1.n119 VDD1.n69 10.4732
R1926 VDD1.n22 VDD1.n21 10.2747
R1927 VDD1.n86 VDD1.n85 10.2747
R1928 VDD1.n58 VDD1.n57 9.69747
R1929 VDD1.n32 VDD1.n17 9.69747
R1930 VDD1.n96 VDD1.n81 9.69747
R1931 VDD1.n123 VDD1.n122 9.69747
R1932 VDD1.n64 VDD1.n63 9.45567
R1933 VDD1.n129 VDD1.n128 9.45567
R1934 VDD1.n24 VDD1.n23 9.3005
R1935 VDD1.n19 VDD1.n18 9.3005
R1936 VDD1.n30 VDD1.n29 9.3005
R1937 VDD1.n32 VDD1.n31 9.3005
R1938 VDD1.n15 VDD1.n14 9.3005
R1939 VDD1.n38 VDD1.n37 9.3005
R1940 VDD1.n40 VDD1.n39 9.3005
R1941 VDD1.n12 VDD1.n9 9.3005
R1942 VDD1.n63 VDD1.n62 9.3005
R1943 VDD1.n2 VDD1.n1 9.3005
R1944 VDD1.n57 VDD1.n56 9.3005
R1945 VDD1.n55 VDD1.n54 9.3005
R1946 VDD1.n6 VDD1.n5 9.3005
R1947 VDD1.n49 VDD1.n48 9.3005
R1948 VDD1.n47 VDD1.n46 9.3005
R1949 VDD1.n128 VDD1.n127 9.3005
R1950 VDD1.n67 VDD1.n66 9.3005
R1951 VDD1.n122 VDD1.n121 9.3005
R1952 VDD1.n120 VDD1.n119 9.3005
R1953 VDD1.n71 VDD1.n70 9.3005
R1954 VDD1.n114 VDD1.n113 9.3005
R1955 VDD1.n112 VDD1.n111 9.3005
R1956 VDD1.n88 VDD1.n87 9.3005
R1957 VDD1.n83 VDD1.n82 9.3005
R1958 VDD1.n94 VDD1.n93 9.3005
R1959 VDD1.n96 VDD1.n95 9.3005
R1960 VDD1.n79 VDD1.n78 9.3005
R1961 VDD1.n102 VDD1.n101 9.3005
R1962 VDD1.n104 VDD1.n103 9.3005
R1963 VDD1.n105 VDD1.n74 9.3005
R1964 VDD1.n61 VDD1.n2 8.92171
R1965 VDD1.n29 VDD1.n28 8.92171
R1966 VDD1.n93 VDD1.n92 8.92171
R1967 VDD1.n126 VDD1.n67 8.92171
R1968 VDD1.n62 VDD1.n0 8.14595
R1969 VDD1.n25 VDD1.n19 8.14595
R1970 VDD1.n89 VDD1.n83 8.14595
R1971 VDD1.n127 VDD1.n65 8.14595
R1972 VDD1.n24 VDD1.n21 7.3702
R1973 VDD1.n88 VDD1.n85 7.3702
R1974 VDD1.n64 VDD1.n0 5.81868
R1975 VDD1.n25 VDD1.n24 5.81868
R1976 VDD1.n89 VDD1.n88 5.81868
R1977 VDD1.n129 VDD1.n65 5.81868
R1978 VDD1.n62 VDD1.n61 5.04292
R1979 VDD1.n28 VDD1.n19 5.04292
R1980 VDD1.n92 VDD1.n83 5.04292
R1981 VDD1.n127 VDD1.n126 5.04292
R1982 VDD1.n58 VDD1.n2 4.26717
R1983 VDD1.n29 VDD1.n17 4.26717
R1984 VDD1.n93 VDD1.n81 4.26717
R1985 VDD1.n123 VDD1.n67 4.26717
R1986 VDD1.n57 VDD1.n4 3.49141
R1987 VDD1.n33 VDD1.n32 3.49141
R1988 VDD1.n97 VDD1.n96 3.49141
R1989 VDD1.n122 VDD1.n69 3.49141
R1990 VDD1.n23 VDD1.n22 2.84303
R1991 VDD1.n87 VDD1.n86 2.84303
R1992 VDD1.n54 VDD1.n53 2.71565
R1993 VDD1.n36 VDD1.n15 2.71565
R1994 VDD1.n100 VDD1.n79 2.71565
R1995 VDD1.n119 VDD1.n118 2.71565
R1996 VDD1.n50 VDD1.n6 1.93989
R1997 VDD1.n37 VDD1.n13 1.93989
R1998 VDD1.n101 VDD1.n77 1.93989
R1999 VDD1.n115 VDD1.n71 1.93989
R2000 VDD1.n49 VDD1.n8 1.16414
R2001 VDD1.n41 VDD1.n40 1.16414
R2002 VDD1.n106 VDD1.n104 1.16414
R2003 VDD1.n114 VDD1.n73 1.16414
R2004 VDD1.n46 VDD1.n45 0.388379
R2005 VDD1.n12 VDD1.n10 0.388379
R2006 VDD1.n105 VDD1.n75 0.388379
R2007 VDD1.n111 VDD1.n110 0.388379
R2008 VDD1.n63 VDD1.n1 0.155672
R2009 VDD1.n56 VDD1.n1 0.155672
R2010 VDD1.n56 VDD1.n55 0.155672
R2011 VDD1.n55 VDD1.n5 0.155672
R2012 VDD1.n48 VDD1.n5 0.155672
R2013 VDD1.n48 VDD1.n47 0.155672
R2014 VDD1.n47 VDD1.n9 0.155672
R2015 VDD1.n39 VDD1.n9 0.155672
R2016 VDD1.n39 VDD1.n38 0.155672
R2017 VDD1.n38 VDD1.n14 0.155672
R2018 VDD1.n31 VDD1.n14 0.155672
R2019 VDD1.n31 VDD1.n30 0.155672
R2020 VDD1.n30 VDD1.n18 0.155672
R2021 VDD1.n23 VDD1.n18 0.155672
R2022 VDD1.n87 VDD1.n82 0.155672
R2023 VDD1.n94 VDD1.n82 0.155672
R2024 VDD1.n95 VDD1.n94 0.155672
R2025 VDD1.n95 VDD1.n78 0.155672
R2026 VDD1.n102 VDD1.n78 0.155672
R2027 VDD1.n103 VDD1.n102 0.155672
R2028 VDD1.n103 VDD1.n74 0.155672
R2029 VDD1.n112 VDD1.n74 0.155672
R2030 VDD1.n113 VDD1.n112 0.155672
R2031 VDD1.n113 VDD1.n70 0.155672
R2032 VDD1.n120 VDD1.n70 0.155672
R2033 VDD1.n121 VDD1.n120 0.155672
R2034 VDD1.n121 VDD1.n66 0.155672
R2035 VDD1.n128 VDD1.n66 0.155672
C0 VN VTAIL 2.45218f
C1 VDD2 VN 2.79137f
C2 VDD1 VP 2.97293f
C3 VN VP 5.45609f
C4 VDD2 VTAIL 5.13309f
C5 VDD1 VN 0.148113f
C6 VP VTAIL 2.46647f
C7 VDD2 VP 0.332232f
C8 VDD1 VTAIL 5.08265f
C9 VDD2 VDD1 0.672209f
C10 VDD2 B 4.436134f
C11 VDD1 B 7.174f
C12 VTAIL B 7.383361f
C13 VN B 10.6896f
C14 VP B 6.368881f
C15 VDD1.n0 B 0.02813f
C16 VDD1.n1 B 0.020505f
C17 VDD1.n2 B 0.011019f
C18 VDD1.n3 B 0.026044f
C19 VDD1.n4 B 0.011667f
C20 VDD1.n5 B 0.020505f
C21 VDD1.n6 B 0.011019f
C22 VDD1.n7 B 0.026044f
C23 VDD1.n8 B 0.011667f
C24 VDD1.n9 B 0.020505f
C25 VDD1.n10 B 0.011343f
C26 VDD1.n11 B 0.026044f
C27 VDD1.n12 B 0.011019f
C28 VDD1.n13 B 0.011667f
C29 VDD1.n14 B 0.020505f
C30 VDD1.n15 B 0.011019f
C31 VDD1.n16 B 0.026044f
C32 VDD1.n17 B 0.011667f
C33 VDD1.n18 B 0.020505f
C34 VDD1.n19 B 0.011019f
C35 VDD1.n20 B 0.019533f
C36 VDD1.n21 B 0.018411f
C37 VDD1.t1 B 0.043995f
C38 VDD1.n22 B 0.148392f
C39 VDD1.n23 B 1.04084f
C40 VDD1.n24 B 0.011019f
C41 VDD1.n25 B 0.011667f
C42 VDD1.n26 B 0.026044f
C43 VDD1.n27 B 0.026044f
C44 VDD1.n28 B 0.011667f
C45 VDD1.n29 B 0.011019f
C46 VDD1.n30 B 0.020505f
C47 VDD1.n31 B 0.020505f
C48 VDD1.n32 B 0.011019f
C49 VDD1.n33 B 0.011667f
C50 VDD1.n34 B 0.026044f
C51 VDD1.n35 B 0.026044f
C52 VDD1.n36 B 0.011667f
C53 VDD1.n37 B 0.011019f
C54 VDD1.n38 B 0.020505f
C55 VDD1.n39 B 0.020505f
C56 VDD1.n40 B 0.011019f
C57 VDD1.n41 B 0.011667f
C58 VDD1.n42 B 0.026044f
C59 VDD1.n43 B 0.026044f
C60 VDD1.n44 B 0.026044f
C61 VDD1.n45 B 0.011343f
C62 VDD1.n46 B 0.011019f
C63 VDD1.n47 B 0.020505f
C64 VDD1.n48 B 0.020505f
C65 VDD1.n49 B 0.011019f
C66 VDD1.n50 B 0.011667f
C67 VDD1.n51 B 0.026044f
C68 VDD1.n52 B 0.026044f
C69 VDD1.n53 B 0.011667f
C70 VDD1.n54 B 0.011019f
C71 VDD1.n55 B 0.020505f
C72 VDD1.n56 B 0.020505f
C73 VDD1.n57 B 0.011019f
C74 VDD1.n58 B 0.011667f
C75 VDD1.n59 B 0.026044f
C76 VDD1.n60 B 0.055158f
C77 VDD1.n61 B 0.011667f
C78 VDD1.n62 B 0.011019f
C79 VDD1.n63 B 0.045996f
C80 VDD1.n64 B 0.046048f
C81 VDD1.n65 B 0.02813f
C82 VDD1.n66 B 0.020505f
C83 VDD1.n67 B 0.011019f
C84 VDD1.n68 B 0.026044f
C85 VDD1.n69 B 0.011667f
C86 VDD1.n70 B 0.020505f
C87 VDD1.n71 B 0.011019f
C88 VDD1.n72 B 0.026044f
C89 VDD1.n73 B 0.011667f
C90 VDD1.n74 B 0.020505f
C91 VDD1.n75 B 0.011343f
C92 VDD1.n76 B 0.026044f
C93 VDD1.n77 B 0.011667f
C94 VDD1.n78 B 0.020505f
C95 VDD1.n79 B 0.011019f
C96 VDD1.n80 B 0.026044f
C97 VDD1.n81 B 0.011667f
C98 VDD1.n82 B 0.020505f
C99 VDD1.n83 B 0.011019f
C100 VDD1.n84 B 0.019533f
C101 VDD1.n85 B 0.018411f
C102 VDD1.t0 B 0.043995f
C103 VDD1.n86 B 0.148392f
C104 VDD1.n87 B 1.04084f
C105 VDD1.n88 B 0.011019f
C106 VDD1.n89 B 0.011667f
C107 VDD1.n90 B 0.026044f
C108 VDD1.n91 B 0.026044f
C109 VDD1.n92 B 0.011667f
C110 VDD1.n93 B 0.011019f
C111 VDD1.n94 B 0.020505f
C112 VDD1.n95 B 0.020505f
C113 VDD1.n96 B 0.011019f
C114 VDD1.n97 B 0.011667f
C115 VDD1.n98 B 0.026044f
C116 VDD1.n99 B 0.026044f
C117 VDD1.n100 B 0.011667f
C118 VDD1.n101 B 0.011019f
C119 VDD1.n102 B 0.020505f
C120 VDD1.n103 B 0.020505f
C121 VDD1.n104 B 0.011019f
C122 VDD1.n105 B 0.011019f
C123 VDD1.n106 B 0.011667f
C124 VDD1.n107 B 0.026044f
C125 VDD1.n108 B 0.026044f
C126 VDD1.n109 B 0.026044f
C127 VDD1.n110 B 0.011343f
C128 VDD1.n111 B 0.011019f
C129 VDD1.n112 B 0.020505f
C130 VDD1.n113 B 0.020505f
C131 VDD1.n114 B 0.011019f
C132 VDD1.n115 B 0.011667f
C133 VDD1.n116 B 0.026044f
C134 VDD1.n117 B 0.026044f
C135 VDD1.n118 B 0.011667f
C136 VDD1.n119 B 0.011019f
C137 VDD1.n120 B 0.020505f
C138 VDD1.n121 B 0.020505f
C139 VDD1.n122 B 0.011019f
C140 VDD1.n123 B 0.011667f
C141 VDD1.n124 B 0.026044f
C142 VDD1.n125 B 0.055158f
C143 VDD1.n126 B 0.011667f
C144 VDD1.n127 B 0.011019f
C145 VDD1.n128 B 0.045996f
C146 VDD1.n129 B 0.649373f
C147 VP.t0 B 3.5942f
C148 VP.t1 B 3.07213f
C149 VP.n0 B 4.25758f
C150 VDD2.n0 B 0.027695f
C151 VDD2.n1 B 0.020188f
C152 VDD2.n2 B 0.010848f
C153 VDD2.n3 B 0.025641f
C154 VDD2.n4 B 0.011486f
C155 VDD2.n5 B 0.020188f
C156 VDD2.n6 B 0.010848f
C157 VDD2.n7 B 0.025641f
C158 VDD2.n8 B 0.011486f
C159 VDD2.n9 B 0.020188f
C160 VDD2.n10 B 0.011167f
C161 VDD2.n11 B 0.025641f
C162 VDD2.n12 B 0.011486f
C163 VDD2.n13 B 0.020188f
C164 VDD2.n14 B 0.010848f
C165 VDD2.n15 B 0.025641f
C166 VDD2.n16 B 0.011486f
C167 VDD2.n17 B 0.020188f
C168 VDD2.n18 B 0.010848f
C169 VDD2.n19 B 0.019231f
C170 VDD2.n20 B 0.018126f
C171 VDD2.t0 B 0.043313f
C172 VDD2.n21 B 0.146094f
C173 VDD2.n22 B 1.02472f
C174 VDD2.n23 B 0.010848f
C175 VDD2.n24 B 0.011486f
C176 VDD2.n25 B 0.025641f
C177 VDD2.n26 B 0.025641f
C178 VDD2.n27 B 0.011486f
C179 VDD2.n28 B 0.010848f
C180 VDD2.n29 B 0.020188f
C181 VDD2.n30 B 0.020188f
C182 VDD2.n31 B 0.010848f
C183 VDD2.n32 B 0.011486f
C184 VDD2.n33 B 0.025641f
C185 VDD2.n34 B 0.025641f
C186 VDD2.n35 B 0.011486f
C187 VDD2.n36 B 0.010848f
C188 VDD2.n37 B 0.020188f
C189 VDD2.n38 B 0.020188f
C190 VDD2.n39 B 0.010848f
C191 VDD2.n40 B 0.010848f
C192 VDD2.n41 B 0.011486f
C193 VDD2.n42 B 0.025641f
C194 VDD2.n43 B 0.025641f
C195 VDD2.n44 B 0.025641f
C196 VDD2.n45 B 0.011167f
C197 VDD2.n46 B 0.010848f
C198 VDD2.n47 B 0.020188f
C199 VDD2.n48 B 0.020188f
C200 VDD2.n49 B 0.010848f
C201 VDD2.n50 B 0.011486f
C202 VDD2.n51 B 0.025641f
C203 VDD2.n52 B 0.025641f
C204 VDD2.n53 B 0.011486f
C205 VDD2.n54 B 0.010848f
C206 VDD2.n55 B 0.020188f
C207 VDD2.n56 B 0.020188f
C208 VDD2.n57 B 0.010848f
C209 VDD2.n58 B 0.011486f
C210 VDD2.n59 B 0.025641f
C211 VDD2.n60 B 0.054304f
C212 VDD2.n61 B 0.011486f
C213 VDD2.n62 B 0.010848f
C214 VDD2.n63 B 0.045284f
C215 VDD2.n64 B 0.599446f
C216 VDD2.n65 B 0.027695f
C217 VDD2.n66 B 0.020188f
C218 VDD2.n67 B 0.010848f
C219 VDD2.n68 B 0.025641f
C220 VDD2.n69 B 0.011486f
C221 VDD2.n70 B 0.020188f
C222 VDD2.n71 B 0.010848f
C223 VDD2.n72 B 0.025641f
C224 VDD2.n73 B 0.011486f
C225 VDD2.n74 B 0.020188f
C226 VDD2.n75 B 0.011167f
C227 VDD2.n76 B 0.025641f
C228 VDD2.n77 B 0.010848f
C229 VDD2.n78 B 0.011486f
C230 VDD2.n79 B 0.020188f
C231 VDD2.n80 B 0.010848f
C232 VDD2.n81 B 0.025641f
C233 VDD2.n82 B 0.011486f
C234 VDD2.n83 B 0.020188f
C235 VDD2.n84 B 0.010848f
C236 VDD2.n85 B 0.019231f
C237 VDD2.n86 B 0.018126f
C238 VDD2.t1 B 0.043313f
C239 VDD2.n87 B 0.146094f
C240 VDD2.n88 B 1.02472f
C241 VDD2.n89 B 0.010848f
C242 VDD2.n90 B 0.011486f
C243 VDD2.n91 B 0.025641f
C244 VDD2.n92 B 0.025641f
C245 VDD2.n93 B 0.011486f
C246 VDD2.n94 B 0.010848f
C247 VDD2.n95 B 0.020188f
C248 VDD2.n96 B 0.020188f
C249 VDD2.n97 B 0.010848f
C250 VDD2.n98 B 0.011486f
C251 VDD2.n99 B 0.025641f
C252 VDD2.n100 B 0.025641f
C253 VDD2.n101 B 0.011486f
C254 VDD2.n102 B 0.010848f
C255 VDD2.n103 B 0.020188f
C256 VDD2.n104 B 0.020188f
C257 VDD2.n105 B 0.010848f
C258 VDD2.n106 B 0.011486f
C259 VDD2.n107 B 0.025641f
C260 VDD2.n108 B 0.025641f
C261 VDD2.n109 B 0.025641f
C262 VDD2.n110 B 0.011167f
C263 VDD2.n111 B 0.010848f
C264 VDD2.n112 B 0.020188f
C265 VDD2.n113 B 0.020188f
C266 VDD2.n114 B 0.010848f
C267 VDD2.n115 B 0.011486f
C268 VDD2.n116 B 0.025641f
C269 VDD2.n117 B 0.025641f
C270 VDD2.n118 B 0.011486f
C271 VDD2.n119 B 0.010848f
C272 VDD2.n120 B 0.020188f
C273 VDD2.n121 B 0.020188f
C274 VDD2.n122 B 0.010848f
C275 VDD2.n123 B 0.011486f
C276 VDD2.n124 B 0.025641f
C277 VDD2.n125 B 0.054304f
C278 VDD2.n126 B 0.011486f
C279 VDD2.n127 B 0.010848f
C280 VDD2.n128 B 0.045284f
C281 VDD2.n129 B 0.044169f
C282 VDD2.n130 B 2.46054f
C283 VTAIL.n0 B 0.028526f
C284 VTAIL.n1 B 0.020794f
C285 VTAIL.n2 B 0.011174f
C286 VTAIL.n3 B 0.02641f
C287 VTAIL.n4 B 0.011831f
C288 VTAIL.n5 B 0.020794f
C289 VTAIL.n6 B 0.011174f
C290 VTAIL.n7 B 0.02641f
C291 VTAIL.n8 B 0.011831f
C292 VTAIL.n9 B 0.020794f
C293 VTAIL.n10 B 0.011502f
C294 VTAIL.n11 B 0.02641f
C295 VTAIL.n12 B 0.011831f
C296 VTAIL.n13 B 0.020794f
C297 VTAIL.n14 B 0.011174f
C298 VTAIL.n15 B 0.02641f
C299 VTAIL.n16 B 0.011831f
C300 VTAIL.n17 B 0.020794f
C301 VTAIL.n18 B 0.011174f
C302 VTAIL.n19 B 0.019808f
C303 VTAIL.n20 B 0.01867f
C304 VTAIL.t1 B 0.044613f
C305 VTAIL.n21 B 0.15048f
C306 VTAIL.n22 B 1.05549f
C307 VTAIL.n23 B 0.011174f
C308 VTAIL.n24 B 0.011831f
C309 VTAIL.n25 B 0.02641f
C310 VTAIL.n26 B 0.02641f
C311 VTAIL.n27 B 0.011831f
C312 VTAIL.n28 B 0.011174f
C313 VTAIL.n29 B 0.020794f
C314 VTAIL.n30 B 0.020794f
C315 VTAIL.n31 B 0.011174f
C316 VTAIL.n32 B 0.011831f
C317 VTAIL.n33 B 0.02641f
C318 VTAIL.n34 B 0.02641f
C319 VTAIL.n35 B 0.011831f
C320 VTAIL.n36 B 0.011174f
C321 VTAIL.n37 B 0.020794f
C322 VTAIL.n38 B 0.020794f
C323 VTAIL.n39 B 0.011174f
C324 VTAIL.n40 B 0.011174f
C325 VTAIL.n41 B 0.011831f
C326 VTAIL.n42 B 0.02641f
C327 VTAIL.n43 B 0.02641f
C328 VTAIL.n44 B 0.02641f
C329 VTAIL.n45 B 0.011502f
C330 VTAIL.n46 B 0.011174f
C331 VTAIL.n47 B 0.020794f
C332 VTAIL.n48 B 0.020794f
C333 VTAIL.n49 B 0.011174f
C334 VTAIL.n50 B 0.011831f
C335 VTAIL.n51 B 0.02641f
C336 VTAIL.n52 B 0.02641f
C337 VTAIL.n53 B 0.011831f
C338 VTAIL.n54 B 0.011174f
C339 VTAIL.n55 B 0.020794f
C340 VTAIL.n56 B 0.020794f
C341 VTAIL.n57 B 0.011174f
C342 VTAIL.n58 B 0.011831f
C343 VTAIL.n59 B 0.02641f
C344 VTAIL.n60 B 0.055934f
C345 VTAIL.n61 B 0.011831f
C346 VTAIL.n62 B 0.011174f
C347 VTAIL.n63 B 0.046644f
C348 VTAIL.n64 B 0.031125f
C349 VTAIL.n65 B 1.41015f
C350 VTAIL.n66 B 0.028526f
C351 VTAIL.n67 B 0.020794f
C352 VTAIL.n68 B 0.011174f
C353 VTAIL.n69 B 0.02641f
C354 VTAIL.n70 B 0.011831f
C355 VTAIL.n71 B 0.020794f
C356 VTAIL.n72 B 0.011174f
C357 VTAIL.n73 B 0.02641f
C358 VTAIL.n74 B 0.011831f
C359 VTAIL.n75 B 0.020794f
C360 VTAIL.n76 B 0.011502f
C361 VTAIL.n77 B 0.02641f
C362 VTAIL.n78 B 0.011174f
C363 VTAIL.n79 B 0.011831f
C364 VTAIL.n80 B 0.020794f
C365 VTAIL.n81 B 0.011174f
C366 VTAIL.n82 B 0.02641f
C367 VTAIL.n83 B 0.011831f
C368 VTAIL.n84 B 0.020794f
C369 VTAIL.n85 B 0.011174f
C370 VTAIL.n86 B 0.019808f
C371 VTAIL.n87 B 0.01867f
C372 VTAIL.t2 B 0.044613f
C373 VTAIL.n88 B 0.15048f
C374 VTAIL.n89 B 1.05549f
C375 VTAIL.n90 B 0.011174f
C376 VTAIL.n91 B 0.011831f
C377 VTAIL.n92 B 0.02641f
C378 VTAIL.n93 B 0.02641f
C379 VTAIL.n94 B 0.011831f
C380 VTAIL.n95 B 0.011174f
C381 VTAIL.n96 B 0.020794f
C382 VTAIL.n97 B 0.020794f
C383 VTAIL.n98 B 0.011174f
C384 VTAIL.n99 B 0.011831f
C385 VTAIL.n100 B 0.02641f
C386 VTAIL.n101 B 0.02641f
C387 VTAIL.n102 B 0.011831f
C388 VTAIL.n103 B 0.011174f
C389 VTAIL.n104 B 0.020794f
C390 VTAIL.n105 B 0.020794f
C391 VTAIL.n106 B 0.011174f
C392 VTAIL.n107 B 0.011831f
C393 VTAIL.n108 B 0.02641f
C394 VTAIL.n109 B 0.02641f
C395 VTAIL.n110 B 0.02641f
C396 VTAIL.n111 B 0.011502f
C397 VTAIL.n112 B 0.011174f
C398 VTAIL.n113 B 0.020794f
C399 VTAIL.n114 B 0.020794f
C400 VTAIL.n115 B 0.011174f
C401 VTAIL.n116 B 0.011831f
C402 VTAIL.n117 B 0.02641f
C403 VTAIL.n118 B 0.02641f
C404 VTAIL.n119 B 0.011831f
C405 VTAIL.n120 B 0.011174f
C406 VTAIL.n121 B 0.020794f
C407 VTAIL.n122 B 0.020794f
C408 VTAIL.n123 B 0.011174f
C409 VTAIL.n124 B 0.011831f
C410 VTAIL.n125 B 0.02641f
C411 VTAIL.n126 B 0.055934f
C412 VTAIL.n127 B 0.011831f
C413 VTAIL.n128 B 0.011174f
C414 VTAIL.n129 B 0.046644f
C415 VTAIL.n130 B 0.031125f
C416 VTAIL.n131 B 1.44828f
C417 VTAIL.n132 B 0.028526f
C418 VTAIL.n133 B 0.020794f
C419 VTAIL.n134 B 0.011174f
C420 VTAIL.n135 B 0.02641f
C421 VTAIL.n136 B 0.011831f
C422 VTAIL.n137 B 0.020794f
C423 VTAIL.n138 B 0.011174f
C424 VTAIL.n139 B 0.02641f
C425 VTAIL.n140 B 0.011831f
C426 VTAIL.n141 B 0.020794f
C427 VTAIL.n142 B 0.011502f
C428 VTAIL.n143 B 0.02641f
C429 VTAIL.n144 B 0.011174f
C430 VTAIL.n145 B 0.011831f
C431 VTAIL.n146 B 0.020794f
C432 VTAIL.n147 B 0.011174f
C433 VTAIL.n148 B 0.02641f
C434 VTAIL.n149 B 0.011831f
C435 VTAIL.n150 B 0.020794f
C436 VTAIL.n151 B 0.011174f
C437 VTAIL.n152 B 0.019808f
C438 VTAIL.n153 B 0.01867f
C439 VTAIL.t0 B 0.044613f
C440 VTAIL.n154 B 0.15048f
C441 VTAIL.n155 B 1.05549f
C442 VTAIL.n156 B 0.011174f
C443 VTAIL.n157 B 0.011831f
C444 VTAIL.n158 B 0.02641f
C445 VTAIL.n159 B 0.02641f
C446 VTAIL.n160 B 0.011831f
C447 VTAIL.n161 B 0.011174f
C448 VTAIL.n162 B 0.020794f
C449 VTAIL.n163 B 0.020794f
C450 VTAIL.n164 B 0.011174f
C451 VTAIL.n165 B 0.011831f
C452 VTAIL.n166 B 0.02641f
C453 VTAIL.n167 B 0.02641f
C454 VTAIL.n168 B 0.011831f
C455 VTAIL.n169 B 0.011174f
C456 VTAIL.n170 B 0.020794f
C457 VTAIL.n171 B 0.020794f
C458 VTAIL.n172 B 0.011174f
C459 VTAIL.n173 B 0.011831f
C460 VTAIL.n174 B 0.02641f
C461 VTAIL.n175 B 0.02641f
C462 VTAIL.n176 B 0.02641f
C463 VTAIL.n177 B 0.011502f
C464 VTAIL.n178 B 0.011174f
C465 VTAIL.n179 B 0.020794f
C466 VTAIL.n180 B 0.020794f
C467 VTAIL.n181 B 0.011174f
C468 VTAIL.n182 B 0.011831f
C469 VTAIL.n183 B 0.02641f
C470 VTAIL.n184 B 0.02641f
C471 VTAIL.n185 B 0.011831f
C472 VTAIL.n186 B 0.011174f
C473 VTAIL.n187 B 0.020794f
C474 VTAIL.n188 B 0.020794f
C475 VTAIL.n189 B 0.011174f
C476 VTAIL.n190 B 0.011831f
C477 VTAIL.n191 B 0.02641f
C478 VTAIL.n192 B 0.055934f
C479 VTAIL.n193 B 0.011831f
C480 VTAIL.n194 B 0.011174f
C481 VTAIL.n195 B 0.046644f
C482 VTAIL.n196 B 0.031125f
C483 VTAIL.n197 B 1.28019f
C484 VTAIL.n198 B 0.028526f
C485 VTAIL.n199 B 0.020794f
C486 VTAIL.n200 B 0.011174f
C487 VTAIL.n201 B 0.02641f
C488 VTAIL.n202 B 0.011831f
C489 VTAIL.n203 B 0.020794f
C490 VTAIL.n204 B 0.011174f
C491 VTAIL.n205 B 0.02641f
C492 VTAIL.n206 B 0.011831f
C493 VTAIL.n207 B 0.020794f
C494 VTAIL.n208 B 0.011502f
C495 VTAIL.n209 B 0.02641f
C496 VTAIL.n210 B 0.011831f
C497 VTAIL.n211 B 0.020794f
C498 VTAIL.n212 B 0.011174f
C499 VTAIL.n213 B 0.02641f
C500 VTAIL.n214 B 0.011831f
C501 VTAIL.n215 B 0.020794f
C502 VTAIL.n216 B 0.011174f
C503 VTAIL.n217 B 0.019808f
C504 VTAIL.n218 B 0.01867f
C505 VTAIL.t3 B 0.044613f
C506 VTAIL.n219 B 0.15048f
C507 VTAIL.n220 B 1.05549f
C508 VTAIL.n221 B 0.011174f
C509 VTAIL.n222 B 0.011831f
C510 VTAIL.n223 B 0.02641f
C511 VTAIL.n224 B 0.02641f
C512 VTAIL.n225 B 0.011831f
C513 VTAIL.n226 B 0.011174f
C514 VTAIL.n227 B 0.020794f
C515 VTAIL.n228 B 0.020794f
C516 VTAIL.n229 B 0.011174f
C517 VTAIL.n230 B 0.011831f
C518 VTAIL.n231 B 0.02641f
C519 VTAIL.n232 B 0.02641f
C520 VTAIL.n233 B 0.011831f
C521 VTAIL.n234 B 0.011174f
C522 VTAIL.n235 B 0.020794f
C523 VTAIL.n236 B 0.020794f
C524 VTAIL.n237 B 0.011174f
C525 VTAIL.n238 B 0.011174f
C526 VTAIL.n239 B 0.011831f
C527 VTAIL.n240 B 0.02641f
C528 VTAIL.n241 B 0.02641f
C529 VTAIL.n242 B 0.02641f
C530 VTAIL.n243 B 0.011502f
C531 VTAIL.n244 B 0.011174f
C532 VTAIL.n245 B 0.020794f
C533 VTAIL.n246 B 0.020794f
C534 VTAIL.n247 B 0.011174f
C535 VTAIL.n248 B 0.011831f
C536 VTAIL.n249 B 0.02641f
C537 VTAIL.n250 B 0.02641f
C538 VTAIL.n251 B 0.011831f
C539 VTAIL.n252 B 0.011174f
C540 VTAIL.n253 B 0.020794f
C541 VTAIL.n254 B 0.020794f
C542 VTAIL.n255 B 0.011174f
C543 VTAIL.n256 B 0.011831f
C544 VTAIL.n257 B 0.02641f
C545 VTAIL.n258 B 0.055934f
C546 VTAIL.n259 B 0.011831f
C547 VTAIL.n260 B 0.011174f
C548 VTAIL.n261 B 0.046644f
C549 VTAIL.n262 B 0.031125f
C550 VTAIL.n263 B 1.20279f
C551 VN.t1 B 3.00593f
C552 VN.t0 B 3.51773f
.ends

