* NGSPICE file created from diff_pair_sample_0105.ext - technology: sky130A

.subckt diff_pair_sample_0105 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=2.33145 pd=14.46 as=5.5107 ps=29.04 w=14.13 l=0.61
X1 VTAIL.t3 VP.t1 VDD1.t6 B.t7 sky130_fd_pr__nfet_01v8 ad=5.5107 pd=29.04 as=2.33145 ps=14.46 w=14.13 l=0.61
X2 B.t21 B.t19 B.t20 B.t13 sky130_fd_pr__nfet_01v8 ad=5.5107 pd=29.04 as=0 ps=0 w=14.13 l=0.61
X3 VDD1.t5 VP.t2 VTAIL.t9 B.t6 sky130_fd_pr__nfet_01v8 ad=2.33145 pd=14.46 as=5.5107 ps=29.04 w=14.13 l=0.61
X4 VDD2.t7 VN.t0 VTAIL.t15 B.t3 sky130_fd_pr__nfet_01v8 ad=2.33145 pd=14.46 as=2.33145 ps=14.46 w=14.13 l=0.61
X5 VTAIL.t10 VN.t1 VDD2.t6 B.t7 sky130_fd_pr__nfet_01v8 ad=5.5107 pd=29.04 as=2.33145 ps=14.46 w=14.13 l=0.61
X6 VDD1.t4 VP.t3 VTAIL.t7 B.t5 sky130_fd_pr__nfet_01v8 ad=2.33145 pd=14.46 as=2.33145 ps=14.46 w=14.13 l=0.61
X7 VTAIL.t2 VP.t4 VDD1.t3 B.t4 sky130_fd_pr__nfet_01v8 ad=5.5107 pd=29.04 as=2.33145 ps=14.46 w=14.13 l=0.61
X8 B.t18 B.t16 B.t17 B.t9 sky130_fd_pr__nfet_01v8 ad=5.5107 pd=29.04 as=0 ps=0 w=14.13 l=0.61
X9 VDD2.t5 VN.t2 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.33145 pd=14.46 as=5.5107 ps=29.04 w=14.13 l=0.61
X10 VTAIL.t14 VN.t3 VDD2.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=5.5107 pd=29.04 as=2.33145 ps=14.46 w=14.13 l=0.61
X11 VDD2.t3 VN.t4 VTAIL.t13 B.t6 sky130_fd_pr__nfet_01v8 ad=2.33145 pd=14.46 as=5.5107 ps=29.04 w=14.13 l=0.61
X12 VTAIL.t8 VP.t5 VDD1.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=2.33145 pd=14.46 as=2.33145 ps=14.46 w=14.13 l=0.61
X13 VDD1.t1 VP.t6 VTAIL.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=2.33145 pd=14.46 as=2.33145 ps=14.46 w=14.13 l=0.61
X14 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=5.5107 pd=29.04 as=0 ps=0 w=14.13 l=0.61
X15 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=5.5107 pd=29.04 as=0 ps=0 w=14.13 l=0.61
X16 VTAIL.t6 VP.t7 VDD1.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=2.33145 pd=14.46 as=2.33145 ps=14.46 w=14.13 l=0.61
X17 VTAIL.t0 VN.t5 VDD2.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=2.33145 pd=14.46 as=2.33145 ps=14.46 w=14.13 l=0.61
X18 VTAIL.t12 VN.t6 VDD2.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=2.33145 pd=14.46 as=2.33145 ps=14.46 w=14.13 l=0.61
X19 VDD2.t0 VN.t7 VTAIL.t11 B.t5 sky130_fd_pr__nfet_01v8 ad=2.33145 pd=14.46 as=2.33145 ps=14.46 w=14.13 l=0.61
R0 VP.n3 VP.t1 649.865
R1 VP.n1 VP.t4 623.044
R2 VP.n10 VP.t6 623.044
R3 VP.n11 VP.t7 623.044
R4 VP.n12 VP.t2 623.044
R5 VP.n6 VP.t0 623.044
R6 VP.n5 VP.t5 623.044
R7 VP.n4 VP.t3 623.044
R8 VP.n13 VP.n12 161.3
R9 VP.n7 VP.n6 161.3
R10 VP.n8 VP.n1 161.3
R11 VP.n5 VP.n2 80.6037
R12 VP.n11 VP.n0 80.6037
R13 VP.n10 VP.n9 80.6037
R14 VP.n10 VP.n1 48.2005
R15 VP.n11 VP.n10 48.2005
R16 VP.n12 VP.n11 48.2005
R17 VP.n6 VP.n5 48.2005
R18 VP.n5 VP.n4 48.2005
R19 VP.n3 VP.n2 45.2318
R20 VP.n8 VP.n7 43.2505
R21 VP.n4 VP.n3 13.3799
R22 VP.n9 VP.n0 0.380177
R23 VP.n7 VP.n2 0.285035
R24 VP.n9 VP.n8 0.285035
R25 VP.n13 VP.n0 0.285035
R26 VP VP.n13 0.0516364
R27 VTAIL.n626 VTAIL.n554 289.615
R28 VTAIL.n74 VTAIL.n2 289.615
R29 VTAIL.n152 VTAIL.n80 289.615
R30 VTAIL.n232 VTAIL.n160 289.615
R31 VTAIL.n548 VTAIL.n476 289.615
R32 VTAIL.n468 VTAIL.n396 289.615
R33 VTAIL.n390 VTAIL.n318 289.615
R34 VTAIL.n310 VTAIL.n238 289.615
R35 VTAIL.n578 VTAIL.n577 185
R36 VTAIL.n583 VTAIL.n582 185
R37 VTAIL.n585 VTAIL.n584 185
R38 VTAIL.n574 VTAIL.n573 185
R39 VTAIL.n591 VTAIL.n590 185
R40 VTAIL.n593 VTAIL.n592 185
R41 VTAIL.n570 VTAIL.n569 185
R42 VTAIL.n599 VTAIL.n598 185
R43 VTAIL.n601 VTAIL.n600 185
R44 VTAIL.n566 VTAIL.n565 185
R45 VTAIL.n607 VTAIL.n606 185
R46 VTAIL.n609 VTAIL.n608 185
R47 VTAIL.n562 VTAIL.n561 185
R48 VTAIL.n615 VTAIL.n614 185
R49 VTAIL.n617 VTAIL.n616 185
R50 VTAIL.n558 VTAIL.n557 185
R51 VTAIL.n624 VTAIL.n623 185
R52 VTAIL.n625 VTAIL.n556 185
R53 VTAIL.n627 VTAIL.n626 185
R54 VTAIL.n26 VTAIL.n25 185
R55 VTAIL.n31 VTAIL.n30 185
R56 VTAIL.n33 VTAIL.n32 185
R57 VTAIL.n22 VTAIL.n21 185
R58 VTAIL.n39 VTAIL.n38 185
R59 VTAIL.n41 VTAIL.n40 185
R60 VTAIL.n18 VTAIL.n17 185
R61 VTAIL.n47 VTAIL.n46 185
R62 VTAIL.n49 VTAIL.n48 185
R63 VTAIL.n14 VTAIL.n13 185
R64 VTAIL.n55 VTAIL.n54 185
R65 VTAIL.n57 VTAIL.n56 185
R66 VTAIL.n10 VTAIL.n9 185
R67 VTAIL.n63 VTAIL.n62 185
R68 VTAIL.n65 VTAIL.n64 185
R69 VTAIL.n6 VTAIL.n5 185
R70 VTAIL.n72 VTAIL.n71 185
R71 VTAIL.n73 VTAIL.n4 185
R72 VTAIL.n75 VTAIL.n74 185
R73 VTAIL.n104 VTAIL.n103 185
R74 VTAIL.n109 VTAIL.n108 185
R75 VTAIL.n111 VTAIL.n110 185
R76 VTAIL.n100 VTAIL.n99 185
R77 VTAIL.n117 VTAIL.n116 185
R78 VTAIL.n119 VTAIL.n118 185
R79 VTAIL.n96 VTAIL.n95 185
R80 VTAIL.n125 VTAIL.n124 185
R81 VTAIL.n127 VTAIL.n126 185
R82 VTAIL.n92 VTAIL.n91 185
R83 VTAIL.n133 VTAIL.n132 185
R84 VTAIL.n135 VTAIL.n134 185
R85 VTAIL.n88 VTAIL.n87 185
R86 VTAIL.n141 VTAIL.n140 185
R87 VTAIL.n143 VTAIL.n142 185
R88 VTAIL.n84 VTAIL.n83 185
R89 VTAIL.n150 VTAIL.n149 185
R90 VTAIL.n151 VTAIL.n82 185
R91 VTAIL.n153 VTAIL.n152 185
R92 VTAIL.n184 VTAIL.n183 185
R93 VTAIL.n189 VTAIL.n188 185
R94 VTAIL.n191 VTAIL.n190 185
R95 VTAIL.n180 VTAIL.n179 185
R96 VTAIL.n197 VTAIL.n196 185
R97 VTAIL.n199 VTAIL.n198 185
R98 VTAIL.n176 VTAIL.n175 185
R99 VTAIL.n205 VTAIL.n204 185
R100 VTAIL.n207 VTAIL.n206 185
R101 VTAIL.n172 VTAIL.n171 185
R102 VTAIL.n213 VTAIL.n212 185
R103 VTAIL.n215 VTAIL.n214 185
R104 VTAIL.n168 VTAIL.n167 185
R105 VTAIL.n221 VTAIL.n220 185
R106 VTAIL.n223 VTAIL.n222 185
R107 VTAIL.n164 VTAIL.n163 185
R108 VTAIL.n230 VTAIL.n229 185
R109 VTAIL.n231 VTAIL.n162 185
R110 VTAIL.n233 VTAIL.n232 185
R111 VTAIL.n549 VTAIL.n548 185
R112 VTAIL.n547 VTAIL.n478 185
R113 VTAIL.n546 VTAIL.n545 185
R114 VTAIL.n481 VTAIL.n479 185
R115 VTAIL.n540 VTAIL.n539 185
R116 VTAIL.n538 VTAIL.n537 185
R117 VTAIL.n485 VTAIL.n484 185
R118 VTAIL.n532 VTAIL.n531 185
R119 VTAIL.n530 VTAIL.n529 185
R120 VTAIL.n489 VTAIL.n488 185
R121 VTAIL.n524 VTAIL.n523 185
R122 VTAIL.n522 VTAIL.n521 185
R123 VTAIL.n493 VTAIL.n492 185
R124 VTAIL.n516 VTAIL.n515 185
R125 VTAIL.n514 VTAIL.n513 185
R126 VTAIL.n497 VTAIL.n496 185
R127 VTAIL.n508 VTAIL.n507 185
R128 VTAIL.n506 VTAIL.n505 185
R129 VTAIL.n501 VTAIL.n500 185
R130 VTAIL.n469 VTAIL.n468 185
R131 VTAIL.n467 VTAIL.n398 185
R132 VTAIL.n466 VTAIL.n465 185
R133 VTAIL.n401 VTAIL.n399 185
R134 VTAIL.n460 VTAIL.n459 185
R135 VTAIL.n458 VTAIL.n457 185
R136 VTAIL.n405 VTAIL.n404 185
R137 VTAIL.n452 VTAIL.n451 185
R138 VTAIL.n450 VTAIL.n449 185
R139 VTAIL.n409 VTAIL.n408 185
R140 VTAIL.n444 VTAIL.n443 185
R141 VTAIL.n442 VTAIL.n441 185
R142 VTAIL.n413 VTAIL.n412 185
R143 VTAIL.n436 VTAIL.n435 185
R144 VTAIL.n434 VTAIL.n433 185
R145 VTAIL.n417 VTAIL.n416 185
R146 VTAIL.n428 VTAIL.n427 185
R147 VTAIL.n426 VTAIL.n425 185
R148 VTAIL.n421 VTAIL.n420 185
R149 VTAIL.n391 VTAIL.n390 185
R150 VTAIL.n389 VTAIL.n320 185
R151 VTAIL.n388 VTAIL.n387 185
R152 VTAIL.n323 VTAIL.n321 185
R153 VTAIL.n382 VTAIL.n381 185
R154 VTAIL.n380 VTAIL.n379 185
R155 VTAIL.n327 VTAIL.n326 185
R156 VTAIL.n374 VTAIL.n373 185
R157 VTAIL.n372 VTAIL.n371 185
R158 VTAIL.n331 VTAIL.n330 185
R159 VTAIL.n366 VTAIL.n365 185
R160 VTAIL.n364 VTAIL.n363 185
R161 VTAIL.n335 VTAIL.n334 185
R162 VTAIL.n358 VTAIL.n357 185
R163 VTAIL.n356 VTAIL.n355 185
R164 VTAIL.n339 VTAIL.n338 185
R165 VTAIL.n350 VTAIL.n349 185
R166 VTAIL.n348 VTAIL.n347 185
R167 VTAIL.n343 VTAIL.n342 185
R168 VTAIL.n311 VTAIL.n310 185
R169 VTAIL.n309 VTAIL.n240 185
R170 VTAIL.n308 VTAIL.n307 185
R171 VTAIL.n243 VTAIL.n241 185
R172 VTAIL.n302 VTAIL.n301 185
R173 VTAIL.n300 VTAIL.n299 185
R174 VTAIL.n247 VTAIL.n246 185
R175 VTAIL.n294 VTAIL.n293 185
R176 VTAIL.n292 VTAIL.n291 185
R177 VTAIL.n251 VTAIL.n250 185
R178 VTAIL.n286 VTAIL.n285 185
R179 VTAIL.n284 VTAIL.n283 185
R180 VTAIL.n255 VTAIL.n254 185
R181 VTAIL.n278 VTAIL.n277 185
R182 VTAIL.n276 VTAIL.n275 185
R183 VTAIL.n259 VTAIL.n258 185
R184 VTAIL.n270 VTAIL.n269 185
R185 VTAIL.n268 VTAIL.n267 185
R186 VTAIL.n263 VTAIL.n262 185
R187 VTAIL.n579 VTAIL.t1 147.659
R188 VTAIL.n27 VTAIL.t10 147.659
R189 VTAIL.n105 VTAIL.t9 147.659
R190 VTAIL.n185 VTAIL.t2 147.659
R191 VTAIL.n502 VTAIL.t5 147.659
R192 VTAIL.n422 VTAIL.t3 147.659
R193 VTAIL.n344 VTAIL.t13 147.659
R194 VTAIL.n264 VTAIL.t14 147.659
R195 VTAIL.n583 VTAIL.n577 104.615
R196 VTAIL.n584 VTAIL.n583 104.615
R197 VTAIL.n584 VTAIL.n573 104.615
R198 VTAIL.n591 VTAIL.n573 104.615
R199 VTAIL.n592 VTAIL.n591 104.615
R200 VTAIL.n592 VTAIL.n569 104.615
R201 VTAIL.n599 VTAIL.n569 104.615
R202 VTAIL.n600 VTAIL.n599 104.615
R203 VTAIL.n600 VTAIL.n565 104.615
R204 VTAIL.n607 VTAIL.n565 104.615
R205 VTAIL.n608 VTAIL.n607 104.615
R206 VTAIL.n608 VTAIL.n561 104.615
R207 VTAIL.n615 VTAIL.n561 104.615
R208 VTAIL.n616 VTAIL.n615 104.615
R209 VTAIL.n616 VTAIL.n557 104.615
R210 VTAIL.n624 VTAIL.n557 104.615
R211 VTAIL.n625 VTAIL.n624 104.615
R212 VTAIL.n626 VTAIL.n625 104.615
R213 VTAIL.n31 VTAIL.n25 104.615
R214 VTAIL.n32 VTAIL.n31 104.615
R215 VTAIL.n32 VTAIL.n21 104.615
R216 VTAIL.n39 VTAIL.n21 104.615
R217 VTAIL.n40 VTAIL.n39 104.615
R218 VTAIL.n40 VTAIL.n17 104.615
R219 VTAIL.n47 VTAIL.n17 104.615
R220 VTAIL.n48 VTAIL.n47 104.615
R221 VTAIL.n48 VTAIL.n13 104.615
R222 VTAIL.n55 VTAIL.n13 104.615
R223 VTAIL.n56 VTAIL.n55 104.615
R224 VTAIL.n56 VTAIL.n9 104.615
R225 VTAIL.n63 VTAIL.n9 104.615
R226 VTAIL.n64 VTAIL.n63 104.615
R227 VTAIL.n64 VTAIL.n5 104.615
R228 VTAIL.n72 VTAIL.n5 104.615
R229 VTAIL.n73 VTAIL.n72 104.615
R230 VTAIL.n74 VTAIL.n73 104.615
R231 VTAIL.n109 VTAIL.n103 104.615
R232 VTAIL.n110 VTAIL.n109 104.615
R233 VTAIL.n110 VTAIL.n99 104.615
R234 VTAIL.n117 VTAIL.n99 104.615
R235 VTAIL.n118 VTAIL.n117 104.615
R236 VTAIL.n118 VTAIL.n95 104.615
R237 VTAIL.n125 VTAIL.n95 104.615
R238 VTAIL.n126 VTAIL.n125 104.615
R239 VTAIL.n126 VTAIL.n91 104.615
R240 VTAIL.n133 VTAIL.n91 104.615
R241 VTAIL.n134 VTAIL.n133 104.615
R242 VTAIL.n134 VTAIL.n87 104.615
R243 VTAIL.n141 VTAIL.n87 104.615
R244 VTAIL.n142 VTAIL.n141 104.615
R245 VTAIL.n142 VTAIL.n83 104.615
R246 VTAIL.n150 VTAIL.n83 104.615
R247 VTAIL.n151 VTAIL.n150 104.615
R248 VTAIL.n152 VTAIL.n151 104.615
R249 VTAIL.n189 VTAIL.n183 104.615
R250 VTAIL.n190 VTAIL.n189 104.615
R251 VTAIL.n190 VTAIL.n179 104.615
R252 VTAIL.n197 VTAIL.n179 104.615
R253 VTAIL.n198 VTAIL.n197 104.615
R254 VTAIL.n198 VTAIL.n175 104.615
R255 VTAIL.n205 VTAIL.n175 104.615
R256 VTAIL.n206 VTAIL.n205 104.615
R257 VTAIL.n206 VTAIL.n171 104.615
R258 VTAIL.n213 VTAIL.n171 104.615
R259 VTAIL.n214 VTAIL.n213 104.615
R260 VTAIL.n214 VTAIL.n167 104.615
R261 VTAIL.n221 VTAIL.n167 104.615
R262 VTAIL.n222 VTAIL.n221 104.615
R263 VTAIL.n222 VTAIL.n163 104.615
R264 VTAIL.n230 VTAIL.n163 104.615
R265 VTAIL.n231 VTAIL.n230 104.615
R266 VTAIL.n232 VTAIL.n231 104.615
R267 VTAIL.n548 VTAIL.n547 104.615
R268 VTAIL.n547 VTAIL.n546 104.615
R269 VTAIL.n546 VTAIL.n479 104.615
R270 VTAIL.n539 VTAIL.n479 104.615
R271 VTAIL.n539 VTAIL.n538 104.615
R272 VTAIL.n538 VTAIL.n484 104.615
R273 VTAIL.n531 VTAIL.n484 104.615
R274 VTAIL.n531 VTAIL.n530 104.615
R275 VTAIL.n530 VTAIL.n488 104.615
R276 VTAIL.n523 VTAIL.n488 104.615
R277 VTAIL.n523 VTAIL.n522 104.615
R278 VTAIL.n522 VTAIL.n492 104.615
R279 VTAIL.n515 VTAIL.n492 104.615
R280 VTAIL.n515 VTAIL.n514 104.615
R281 VTAIL.n514 VTAIL.n496 104.615
R282 VTAIL.n507 VTAIL.n496 104.615
R283 VTAIL.n507 VTAIL.n506 104.615
R284 VTAIL.n506 VTAIL.n500 104.615
R285 VTAIL.n468 VTAIL.n467 104.615
R286 VTAIL.n467 VTAIL.n466 104.615
R287 VTAIL.n466 VTAIL.n399 104.615
R288 VTAIL.n459 VTAIL.n399 104.615
R289 VTAIL.n459 VTAIL.n458 104.615
R290 VTAIL.n458 VTAIL.n404 104.615
R291 VTAIL.n451 VTAIL.n404 104.615
R292 VTAIL.n451 VTAIL.n450 104.615
R293 VTAIL.n450 VTAIL.n408 104.615
R294 VTAIL.n443 VTAIL.n408 104.615
R295 VTAIL.n443 VTAIL.n442 104.615
R296 VTAIL.n442 VTAIL.n412 104.615
R297 VTAIL.n435 VTAIL.n412 104.615
R298 VTAIL.n435 VTAIL.n434 104.615
R299 VTAIL.n434 VTAIL.n416 104.615
R300 VTAIL.n427 VTAIL.n416 104.615
R301 VTAIL.n427 VTAIL.n426 104.615
R302 VTAIL.n426 VTAIL.n420 104.615
R303 VTAIL.n390 VTAIL.n389 104.615
R304 VTAIL.n389 VTAIL.n388 104.615
R305 VTAIL.n388 VTAIL.n321 104.615
R306 VTAIL.n381 VTAIL.n321 104.615
R307 VTAIL.n381 VTAIL.n380 104.615
R308 VTAIL.n380 VTAIL.n326 104.615
R309 VTAIL.n373 VTAIL.n326 104.615
R310 VTAIL.n373 VTAIL.n372 104.615
R311 VTAIL.n372 VTAIL.n330 104.615
R312 VTAIL.n365 VTAIL.n330 104.615
R313 VTAIL.n365 VTAIL.n364 104.615
R314 VTAIL.n364 VTAIL.n334 104.615
R315 VTAIL.n357 VTAIL.n334 104.615
R316 VTAIL.n357 VTAIL.n356 104.615
R317 VTAIL.n356 VTAIL.n338 104.615
R318 VTAIL.n349 VTAIL.n338 104.615
R319 VTAIL.n349 VTAIL.n348 104.615
R320 VTAIL.n348 VTAIL.n342 104.615
R321 VTAIL.n310 VTAIL.n309 104.615
R322 VTAIL.n309 VTAIL.n308 104.615
R323 VTAIL.n308 VTAIL.n241 104.615
R324 VTAIL.n301 VTAIL.n241 104.615
R325 VTAIL.n301 VTAIL.n300 104.615
R326 VTAIL.n300 VTAIL.n246 104.615
R327 VTAIL.n293 VTAIL.n246 104.615
R328 VTAIL.n293 VTAIL.n292 104.615
R329 VTAIL.n292 VTAIL.n250 104.615
R330 VTAIL.n285 VTAIL.n250 104.615
R331 VTAIL.n285 VTAIL.n284 104.615
R332 VTAIL.n284 VTAIL.n254 104.615
R333 VTAIL.n277 VTAIL.n254 104.615
R334 VTAIL.n277 VTAIL.n276 104.615
R335 VTAIL.n276 VTAIL.n258 104.615
R336 VTAIL.n269 VTAIL.n258 104.615
R337 VTAIL.n269 VTAIL.n268 104.615
R338 VTAIL.n268 VTAIL.n262 104.615
R339 VTAIL.t1 VTAIL.n577 52.3082
R340 VTAIL.t10 VTAIL.n25 52.3082
R341 VTAIL.t9 VTAIL.n103 52.3082
R342 VTAIL.t2 VTAIL.n183 52.3082
R343 VTAIL.t5 VTAIL.n500 52.3082
R344 VTAIL.t3 VTAIL.n420 52.3082
R345 VTAIL.t13 VTAIL.n342 52.3082
R346 VTAIL.t14 VTAIL.n262 52.3082
R347 VTAIL.n475 VTAIL.n474 48.4084
R348 VTAIL.n317 VTAIL.n316 48.4084
R349 VTAIL.n1 VTAIL.n0 48.4082
R350 VTAIL.n159 VTAIL.n158 48.4082
R351 VTAIL.n631 VTAIL.n630 36.2581
R352 VTAIL.n79 VTAIL.n78 36.2581
R353 VTAIL.n157 VTAIL.n156 36.2581
R354 VTAIL.n237 VTAIL.n236 36.2581
R355 VTAIL.n553 VTAIL.n552 36.2581
R356 VTAIL.n473 VTAIL.n472 36.2581
R357 VTAIL.n395 VTAIL.n394 36.2581
R358 VTAIL.n315 VTAIL.n314 36.2581
R359 VTAIL.n631 VTAIL.n553 25.3583
R360 VTAIL.n315 VTAIL.n237 25.3583
R361 VTAIL.n579 VTAIL.n578 15.6677
R362 VTAIL.n27 VTAIL.n26 15.6677
R363 VTAIL.n105 VTAIL.n104 15.6677
R364 VTAIL.n185 VTAIL.n184 15.6677
R365 VTAIL.n502 VTAIL.n501 15.6677
R366 VTAIL.n422 VTAIL.n421 15.6677
R367 VTAIL.n344 VTAIL.n343 15.6677
R368 VTAIL.n264 VTAIL.n263 15.6677
R369 VTAIL.n627 VTAIL.n556 13.1884
R370 VTAIL.n75 VTAIL.n4 13.1884
R371 VTAIL.n153 VTAIL.n82 13.1884
R372 VTAIL.n233 VTAIL.n162 13.1884
R373 VTAIL.n549 VTAIL.n478 13.1884
R374 VTAIL.n469 VTAIL.n398 13.1884
R375 VTAIL.n391 VTAIL.n320 13.1884
R376 VTAIL.n311 VTAIL.n240 13.1884
R377 VTAIL.n582 VTAIL.n581 12.8005
R378 VTAIL.n623 VTAIL.n622 12.8005
R379 VTAIL.n628 VTAIL.n554 12.8005
R380 VTAIL.n30 VTAIL.n29 12.8005
R381 VTAIL.n71 VTAIL.n70 12.8005
R382 VTAIL.n76 VTAIL.n2 12.8005
R383 VTAIL.n108 VTAIL.n107 12.8005
R384 VTAIL.n149 VTAIL.n148 12.8005
R385 VTAIL.n154 VTAIL.n80 12.8005
R386 VTAIL.n188 VTAIL.n187 12.8005
R387 VTAIL.n229 VTAIL.n228 12.8005
R388 VTAIL.n234 VTAIL.n160 12.8005
R389 VTAIL.n550 VTAIL.n476 12.8005
R390 VTAIL.n545 VTAIL.n480 12.8005
R391 VTAIL.n505 VTAIL.n504 12.8005
R392 VTAIL.n470 VTAIL.n396 12.8005
R393 VTAIL.n465 VTAIL.n400 12.8005
R394 VTAIL.n425 VTAIL.n424 12.8005
R395 VTAIL.n392 VTAIL.n318 12.8005
R396 VTAIL.n387 VTAIL.n322 12.8005
R397 VTAIL.n347 VTAIL.n346 12.8005
R398 VTAIL.n312 VTAIL.n238 12.8005
R399 VTAIL.n307 VTAIL.n242 12.8005
R400 VTAIL.n267 VTAIL.n266 12.8005
R401 VTAIL.n585 VTAIL.n576 12.0247
R402 VTAIL.n621 VTAIL.n558 12.0247
R403 VTAIL.n33 VTAIL.n24 12.0247
R404 VTAIL.n69 VTAIL.n6 12.0247
R405 VTAIL.n111 VTAIL.n102 12.0247
R406 VTAIL.n147 VTAIL.n84 12.0247
R407 VTAIL.n191 VTAIL.n182 12.0247
R408 VTAIL.n227 VTAIL.n164 12.0247
R409 VTAIL.n544 VTAIL.n481 12.0247
R410 VTAIL.n508 VTAIL.n499 12.0247
R411 VTAIL.n464 VTAIL.n401 12.0247
R412 VTAIL.n428 VTAIL.n419 12.0247
R413 VTAIL.n386 VTAIL.n323 12.0247
R414 VTAIL.n350 VTAIL.n341 12.0247
R415 VTAIL.n306 VTAIL.n243 12.0247
R416 VTAIL.n270 VTAIL.n261 12.0247
R417 VTAIL.n586 VTAIL.n574 11.249
R418 VTAIL.n618 VTAIL.n617 11.249
R419 VTAIL.n34 VTAIL.n22 11.249
R420 VTAIL.n66 VTAIL.n65 11.249
R421 VTAIL.n112 VTAIL.n100 11.249
R422 VTAIL.n144 VTAIL.n143 11.249
R423 VTAIL.n192 VTAIL.n180 11.249
R424 VTAIL.n224 VTAIL.n223 11.249
R425 VTAIL.n541 VTAIL.n540 11.249
R426 VTAIL.n509 VTAIL.n497 11.249
R427 VTAIL.n461 VTAIL.n460 11.249
R428 VTAIL.n429 VTAIL.n417 11.249
R429 VTAIL.n383 VTAIL.n382 11.249
R430 VTAIL.n351 VTAIL.n339 11.249
R431 VTAIL.n303 VTAIL.n302 11.249
R432 VTAIL.n271 VTAIL.n259 11.249
R433 VTAIL.n590 VTAIL.n589 10.4732
R434 VTAIL.n614 VTAIL.n560 10.4732
R435 VTAIL.n38 VTAIL.n37 10.4732
R436 VTAIL.n62 VTAIL.n8 10.4732
R437 VTAIL.n116 VTAIL.n115 10.4732
R438 VTAIL.n140 VTAIL.n86 10.4732
R439 VTAIL.n196 VTAIL.n195 10.4732
R440 VTAIL.n220 VTAIL.n166 10.4732
R441 VTAIL.n537 VTAIL.n483 10.4732
R442 VTAIL.n513 VTAIL.n512 10.4732
R443 VTAIL.n457 VTAIL.n403 10.4732
R444 VTAIL.n433 VTAIL.n432 10.4732
R445 VTAIL.n379 VTAIL.n325 10.4732
R446 VTAIL.n355 VTAIL.n354 10.4732
R447 VTAIL.n299 VTAIL.n245 10.4732
R448 VTAIL.n275 VTAIL.n274 10.4732
R449 VTAIL.n593 VTAIL.n572 9.69747
R450 VTAIL.n613 VTAIL.n562 9.69747
R451 VTAIL.n41 VTAIL.n20 9.69747
R452 VTAIL.n61 VTAIL.n10 9.69747
R453 VTAIL.n119 VTAIL.n98 9.69747
R454 VTAIL.n139 VTAIL.n88 9.69747
R455 VTAIL.n199 VTAIL.n178 9.69747
R456 VTAIL.n219 VTAIL.n168 9.69747
R457 VTAIL.n536 VTAIL.n485 9.69747
R458 VTAIL.n516 VTAIL.n495 9.69747
R459 VTAIL.n456 VTAIL.n405 9.69747
R460 VTAIL.n436 VTAIL.n415 9.69747
R461 VTAIL.n378 VTAIL.n327 9.69747
R462 VTAIL.n358 VTAIL.n337 9.69747
R463 VTAIL.n298 VTAIL.n247 9.69747
R464 VTAIL.n278 VTAIL.n257 9.69747
R465 VTAIL.n630 VTAIL.n629 9.45567
R466 VTAIL.n78 VTAIL.n77 9.45567
R467 VTAIL.n156 VTAIL.n155 9.45567
R468 VTAIL.n236 VTAIL.n235 9.45567
R469 VTAIL.n552 VTAIL.n551 9.45567
R470 VTAIL.n472 VTAIL.n471 9.45567
R471 VTAIL.n394 VTAIL.n393 9.45567
R472 VTAIL.n314 VTAIL.n313 9.45567
R473 VTAIL.n629 VTAIL.n628 9.3005
R474 VTAIL.n568 VTAIL.n567 9.3005
R475 VTAIL.n597 VTAIL.n596 9.3005
R476 VTAIL.n595 VTAIL.n594 9.3005
R477 VTAIL.n572 VTAIL.n571 9.3005
R478 VTAIL.n589 VTAIL.n588 9.3005
R479 VTAIL.n587 VTAIL.n586 9.3005
R480 VTAIL.n576 VTAIL.n575 9.3005
R481 VTAIL.n581 VTAIL.n580 9.3005
R482 VTAIL.n603 VTAIL.n602 9.3005
R483 VTAIL.n605 VTAIL.n604 9.3005
R484 VTAIL.n564 VTAIL.n563 9.3005
R485 VTAIL.n611 VTAIL.n610 9.3005
R486 VTAIL.n613 VTAIL.n612 9.3005
R487 VTAIL.n560 VTAIL.n559 9.3005
R488 VTAIL.n619 VTAIL.n618 9.3005
R489 VTAIL.n621 VTAIL.n620 9.3005
R490 VTAIL.n622 VTAIL.n555 9.3005
R491 VTAIL.n77 VTAIL.n76 9.3005
R492 VTAIL.n16 VTAIL.n15 9.3005
R493 VTAIL.n45 VTAIL.n44 9.3005
R494 VTAIL.n43 VTAIL.n42 9.3005
R495 VTAIL.n20 VTAIL.n19 9.3005
R496 VTAIL.n37 VTAIL.n36 9.3005
R497 VTAIL.n35 VTAIL.n34 9.3005
R498 VTAIL.n24 VTAIL.n23 9.3005
R499 VTAIL.n29 VTAIL.n28 9.3005
R500 VTAIL.n51 VTAIL.n50 9.3005
R501 VTAIL.n53 VTAIL.n52 9.3005
R502 VTAIL.n12 VTAIL.n11 9.3005
R503 VTAIL.n59 VTAIL.n58 9.3005
R504 VTAIL.n61 VTAIL.n60 9.3005
R505 VTAIL.n8 VTAIL.n7 9.3005
R506 VTAIL.n67 VTAIL.n66 9.3005
R507 VTAIL.n69 VTAIL.n68 9.3005
R508 VTAIL.n70 VTAIL.n3 9.3005
R509 VTAIL.n155 VTAIL.n154 9.3005
R510 VTAIL.n94 VTAIL.n93 9.3005
R511 VTAIL.n123 VTAIL.n122 9.3005
R512 VTAIL.n121 VTAIL.n120 9.3005
R513 VTAIL.n98 VTAIL.n97 9.3005
R514 VTAIL.n115 VTAIL.n114 9.3005
R515 VTAIL.n113 VTAIL.n112 9.3005
R516 VTAIL.n102 VTAIL.n101 9.3005
R517 VTAIL.n107 VTAIL.n106 9.3005
R518 VTAIL.n129 VTAIL.n128 9.3005
R519 VTAIL.n131 VTAIL.n130 9.3005
R520 VTAIL.n90 VTAIL.n89 9.3005
R521 VTAIL.n137 VTAIL.n136 9.3005
R522 VTAIL.n139 VTAIL.n138 9.3005
R523 VTAIL.n86 VTAIL.n85 9.3005
R524 VTAIL.n145 VTAIL.n144 9.3005
R525 VTAIL.n147 VTAIL.n146 9.3005
R526 VTAIL.n148 VTAIL.n81 9.3005
R527 VTAIL.n235 VTAIL.n234 9.3005
R528 VTAIL.n174 VTAIL.n173 9.3005
R529 VTAIL.n203 VTAIL.n202 9.3005
R530 VTAIL.n201 VTAIL.n200 9.3005
R531 VTAIL.n178 VTAIL.n177 9.3005
R532 VTAIL.n195 VTAIL.n194 9.3005
R533 VTAIL.n193 VTAIL.n192 9.3005
R534 VTAIL.n182 VTAIL.n181 9.3005
R535 VTAIL.n187 VTAIL.n186 9.3005
R536 VTAIL.n209 VTAIL.n208 9.3005
R537 VTAIL.n211 VTAIL.n210 9.3005
R538 VTAIL.n170 VTAIL.n169 9.3005
R539 VTAIL.n217 VTAIL.n216 9.3005
R540 VTAIL.n219 VTAIL.n218 9.3005
R541 VTAIL.n166 VTAIL.n165 9.3005
R542 VTAIL.n225 VTAIL.n224 9.3005
R543 VTAIL.n227 VTAIL.n226 9.3005
R544 VTAIL.n228 VTAIL.n161 9.3005
R545 VTAIL.n528 VTAIL.n527 9.3005
R546 VTAIL.n487 VTAIL.n486 9.3005
R547 VTAIL.n534 VTAIL.n533 9.3005
R548 VTAIL.n536 VTAIL.n535 9.3005
R549 VTAIL.n483 VTAIL.n482 9.3005
R550 VTAIL.n542 VTAIL.n541 9.3005
R551 VTAIL.n544 VTAIL.n543 9.3005
R552 VTAIL.n480 VTAIL.n477 9.3005
R553 VTAIL.n551 VTAIL.n550 9.3005
R554 VTAIL.n526 VTAIL.n525 9.3005
R555 VTAIL.n491 VTAIL.n490 9.3005
R556 VTAIL.n520 VTAIL.n519 9.3005
R557 VTAIL.n518 VTAIL.n517 9.3005
R558 VTAIL.n495 VTAIL.n494 9.3005
R559 VTAIL.n512 VTAIL.n511 9.3005
R560 VTAIL.n510 VTAIL.n509 9.3005
R561 VTAIL.n499 VTAIL.n498 9.3005
R562 VTAIL.n504 VTAIL.n503 9.3005
R563 VTAIL.n448 VTAIL.n447 9.3005
R564 VTAIL.n407 VTAIL.n406 9.3005
R565 VTAIL.n454 VTAIL.n453 9.3005
R566 VTAIL.n456 VTAIL.n455 9.3005
R567 VTAIL.n403 VTAIL.n402 9.3005
R568 VTAIL.n462 VTAIL.n461 9.3005
R569 VTAIL.n464 VTAIL.n463 9.3005
R570 VTAIL.n400 VTAIL.n397 9.3005
R571 VTAIL.n471 VTAIL.n470 9.3005
R572 VTAIL.n446 VTAIL.n445 9.3005
R573 VTAIL.n411 VTAIL.n410 9.3005
R574 VTAIL.n440 VTAIL.n439 9.3005
R575 VTAIL.n438 VTAIL.n437 9.3005
R576 VTAIL.n415 VTAIL.n414 9.3005
R577 VTAIL.n432 VTAIL.n431 9.3005
R578 VTAIL.n430 VTAIL.n429 9.3005
R579 VTAIL.n419 VTAIL.n418 9.3005
R580 VTAIL.n424 VTAIL.n423 9.3005
R581 VTAIL.n370 VTAIL.n369 9.3005
R582 VTAIL.n329 VTAIL.n328 9.3005
R583 VTAIL.n376 VTAIL.n375 9.3005
R584 VTAIL.n378 VTAIL.n377 9.3005
R585 VTAIL.n325 VTAIL.n324 9.3005
R586 VTAIL.n384 VTAIL.n383 9.3005
R587 VTAIL.n386 VTAIL.n385 9.3005
R588 VTAIL.n322 VTAIL.n319 9.3005
R589 VTAIL.n393 VTAIL.n392 9.3005
R590 VTAIL.n368 VTAIL.n367 9.3005
R591 VTAIL.n333 VTAIL.n332 9.3005
R592 VTAIL.n362 VTAIL.n361 9.3005
R593 VTAIL.n360 VTAIL.n359 9.3005
R594 VTAIL.n337 VTAIL.n336 9.3005
R595 VTAIL.n354 VTAIL.n353 9.3005
R596 VTAIL.n352 VTAIL.n351 9.3005
R597 VTAIL.n341 VTAIL.n340 9.3005
R598 VTAIL.n346 VTAIL.n345 9.3005
R599 VTAIL.n290 VTAIL.n289 9.3005
R600 VTAIL.n249 VTAIL.n248 9.3005
R601 VTAIL.n296 VTAIL.n295 9.3005
R602 VTAIL.n298 VTAIL.n297 9.3005
R603 VTAIL.n245 VTAIL.n244 9.3005
R604 VTAIL.n304 VTAIL.n303 9.3005
R605 VTAIL.n306 VTAIL.n305 9.3005
R606 VTAIL.n242 VTAIL.n239 9.3005
R607 VTAIL.n313 VTAIL.n312 9.3005
R608 VTAIL.n288 VTAIL.n287 9.3005
R609 VTAIL.n253 VTAIL.n252 9.3005
R610 VTAIL.n282 VTAIL.n281 9.3005
R611 VTAIL.n280 VTAIL.n279 9.3005
R612 VTAIL.n257 VTAIL.n256 9.3005
R613 VTAIL.n274 VTAIL.n273 9.3005
R614 VTAIL.n272 VTAIL.n271 9.3005
R615 VTAIL.n261 VTAIL.n260 9.3005
R616 VTAIL.n266 VTAIL.n265 9.3005
R617 VTAIL.n594 VTAIL.n570 8.92171
R618 VTAIL.n610 VTAIL.n609 8.92171
R619 VTAIL.n42 VTAIL.n18 8.92171
R620 VTAIL.n58 VTAIL.n57 8.92171
R621 VTAIL.n120 VTAIL.n96 8.92171
R622 VTAIL.n136 VTAIL.n135 8.92171
R623 VTAIL.n200 VTAIL.n176 8.92171
R624 VTAIL.n216 VTAIL.n215 8.92171
R625 VTAIL.n533 VTAIL.n532 8.92171
R626 VTAIL.n517 VTAIL.n493 8.92171
R627 VTAIL.n453 VTAIL.n452 8.92171
R628 VTAIL.n437 VTAIL.n413 8.92171
R629 VTAIL.n375 VTAIL.n374 8.92171
R630 VTAIL.n359 VTAIL.n335 8.92171
R631 VTAIL.n295 VTAIL.n294 8.92171
R632 VTAIL.n279 VTAIL.n255 8.92171
R633 VTAIL.n598 VTAIL.n597 8.14595
R634 VTAIL.n606 VTAIL.n564 8.14595
R635 VTAIL.n46 VTAIL.n45 8.14595
R636 VTAIL.n54 VTAIL.n12 8.14595
R637 VTAIL.n124 VTAIL.n123 8.14595
R638 VTAIL.n132 VTAIL.n90 8.14595
R639 VTAIL.n204 VTAIL.n203 8.14595
R640 VTAIL.n212 VTAIL.n170 8.14595
R641 VTAIL.n529 VTAIL.n487 8.14595
R642 VTAIL.n521 VTAIL.n520 8.14595
R643 VTAIL.n449 VTAIL.n407 8.14595
R644 VTAIL.n441 VTAIL.n440 8.14595
R645 VTAIL.n371 VTAIL.n329 8.14595
R646 VTAIL.n363 VTAIL.n362 8.14595
R647 VTAIL.n291 VTAIL.n249 8.14595
R648 VTAIL.n283 VTAIL.n282 8.14595
R649 VTAIL.n601 VTAIL.n568 7.3702
R650 VTAIL.n605 VTAIL.n566 7.3702
R651 VTAIL.n49 VTAIL.n16 7.3702
R652 VTAIL.n53 VTAIL.n14 7.3702
R653 VTAIL.n127 VTAIL.n94 7.3702
R654 VTAIL.n131 VTAIL.n92 7.3702
R655 VTAIL.n207 VTAIL.n174 7.3702
R656 VTAIL.n211 VTAIL.n172 7.3702
R657 VTAIL.n528 VTAIL.n489 7.3702
R658 VTAIL.n524 VTAIL.n491 7.3702
R659 VTAIL.n448 VTAIL.n409 7.3702
R660 VTAIL.n444 VTAIL.n411 7.3702
R661 VTAIL.n370 VTAIL.n331 7.3702
R662 VTAIL.n366 VTAIL.n333 7.3702
R663 VTAIL.n290 VTAIL.n251 7.3702
R664 VTAIL.n286 VTAIL.n253 7.3702
R665 VTAIL.n602 VTAIL.n601 6.59444
R666 VTAIL.n602 VTAIL.n566 6.59444
R667 VTAIL.n50 VTAIL.n49 6.59444
R668 VTAIL.n50 VTAIL.n14 6.59444
R669 VTAIL.n128 VTAIL.n127 6.59444
R670 VTAIL.n128 VTAIL.n92 6.59444
R671 VTAIL.n208 VTAIL.n207 6.59444
R672 VTAIL.n208 VTAIL.n172 6.59444
R673 VTAIL.n525 VTAIL.n489 6.59444
R674 VTAIL.n525 VTAIL.n524 6.59444
R675 VTAIL.n445 VTAIL.n409 6.59444
R676 VTAIL.n445 VTAIL.n444 6.59444
R677 VTAIL.n367 VTAIL.n331 6.59444
R678 VTAIL.n367 VTAIL.n366 6.59444
R679 VTAIL.n287 VTAIL.n251 6.59444
R680 VTAIL.n287 VTAIL.n286 6.59444
R681 VTAIL.n598 VTAIL.n568 5.81868
R682 VTAIL.n606 VTAIL.n605 5.81868
R683 VTAIL.n46 VTAIL.n16 5.81868
R684 VTAIL.n54 VTAIL.n53 5.81868
R685 VTAIL.n124 VTAIL.n94 5.81868
R686 VTAIL.n132 VTAIL.n131 5.81868
R687 VTAIL.n204 VTAIL.n174 5.81868
R688 VTAIL.n212 VTAIL.n211 5.81868
R689 VTAIL.n529 VTAIL.n528 5.81868
R690 VTAIL.n521 VTAIL.n491 5.81868
R691 VTAIL.n449 VTAIL.n448 5.81868
R692 VTAIL.n441 VTAIL.n411 5.81868
R693 VTAIL.n371 VTAIL.n370 5.81868
R694 VTAIL.n363 VTAIL.n333 5.81868
R695 VTAIL.n291 VTAIL.n290 5.81868
R696 VTAIL.n283 VTAIL.n253 5.81868
R697 VTAIL.n597 VTAIL.n570 5.04292
R698 VTAIL.n609 VTAIL.n564 5.04292
R699 VTAIL.n45 VTAIL.n18 5.04292
R700 VTAIL.n57 VTAIL.n12 5.04292
R701 VTAIL.n123 VTAIL.n96 5.04292
R702 VTAIL.n135 VTAIL.n90 5.04292
R703 VTAIL.n203 VTAIL.n176 5.04292
R704 VTAIL.n215 VTAIL.n170 5.04292
R705 VTAIL.n532 VTAIL.n487 5.04292
R706 VTAIL.n520 VTAIL.n493 5.04292
R707 VTAIL.n452 VTAIL.n407 5.04292
R708 VTAIL.n440 VTAIL.n413 5.04292
R709 VTAIL.n374 VTAIL.n329 5.04292
R710 VTAIL.n362 VTAIL.n335 5.04292
R711 VTAIL.n294 VTAIL.n249 5.04292
R712 VTAIL.n282 VTAIL.n255 5.04292
R713 VTAIL.n580 VTAIL.n579 4.38563
R714 VTAIL.n28 VTAIL.n27 4.38563
R715 VTAIL.n106 VTAIL.n105 4.38563
R716 VTAIL.n186 VTAIL.n185 4.38563
R717 VTAIL.n503 VTAIL.n502 4.38563
R718 VTAIL.n423 VTAIL.n422 4.38563
R719 VTAIL.n345 VTAIL.n344 4.38563
R720 VTAIL.n265 VTAIL.n264 4.38563
R721 VTAIL.n594 VTAIL.n593 4.26717
R722 VTAIL.n610 VTAIL.n562 4.26717
R723 VTAIL.n42 VTAIL.n41 4.26717
R724 VTAIL.n58 VTAIL.n10 4.26717
R725 VTAIL.n120 VTAIL.n119 4.26717
R726 VTAIL.n136 VTAIL.n88 4.26717
R727 VTAIL.n200 VTAIL.n199 4.26717
R728 VTAIL.n216 VTAIL.n168 4.26717
R729 VTAIL.n533 VTAIL.n485 4.26717
R730 VTAIL.n517 VTAIL.n516 4.26717
R731 VTAIL.n453 VTAIL.n405 4.26717
R732 VTAIL.n437 VTAIL.n436 4.26717
R733 VTAIL.n375 VTAIL.n327 4.26717
R734 VTAIL.n359 VTAIL.n358 4.26717
R735 VTAIL.n295 VTAIL.n247 4.26717
R736 VTAIL.n279 VTAIL.n278 4.26717
R737 VTAIL.n590 VTAIL.n572 3.49141
R738 VTAIL.n614 VTAIL.n613 3.49141
R739 VTAIL.n38 VTAIL.n20 3.49141
R740 VTAIL.n62 VTAIL.n61 3.49141
R741 VTAIL.n116 VTAIL.n98 3.49141
R742 VTAIL.n140 VTAIL.n139 3.49141
R743 VTAIL.n196 VTAIL.n178 3.49141
R744 VTAIL.n220 VTAIL.n219 3.49141
R745 VTAIL.n537 VTAIL.n536 3.49141
R746 VTAIL.n513 VTAIL.n495 3.49141
R747 VTAIL.n457 VTAIL.n456 3.49141
R748 VTAIL.n433 VTAIL.n415 3.49141
R749 VTAIL.n379 VTAIL.n378 3.49141
R750 VTAIL.n355 VTAIL.n337 3.49141
R751 VTAIL.n299 VTAIL.n298 3.49141
R752 VTAIL.n275 VTAIL.n257 3.49141
R753 VTAIL.n589 VTAIL.n574 2.71565
R754 VTAIL.n617 VTAIL.n560 2.71565
R755 VTAIL.n37 VTAIL.n22 2.71565
R756 VTAIL.n65 VTAIL.n8 2.71565
R757 VTAIL.n115 VTAIL.n100 2.71565
R758 VTAIL.n143 VTAIL.n86 2.71565
R759 VTAIL.n195 VTAIL.n180 2.71565
R760 VTAIL.n223 VTAIL.n166 2.71565
R761 VTAIL.n540 VTAIL.n483 2.71565
R762 VTAIL.n512 VTAIL.n497 2.71565
R763 VTAIL.n460 VTAIL.n403 2.71565
R764 VTAIL.n432 VTAIL.n417 2.71565
R765 VTAIL.n382 VTAIL.n325 2.71565
R766 VTAIL.n354 VTAIL.n339 2.71565
R767 VTAIL.n302 VTAIL.n245 2.71565
R768 VTAIL.n274 VTAIL.n259 2.71565
R769 VTAIL.n586 VTAIL.n585 1.93989
R770 VTAIL.n618 VTAIL.n558 1.93989
R771 VTAIL.n34 VTAIL.n33 1.93989
R772 VTAIL.n66 VTAIL.n6 1.93989
R773 VTAIL.n112 VTAIL.n111 1.93989
R774 VTAIL.n144 VTAIL.n84 1.93989
R775 VTAIL.n192 VTAIL.n191 1.93989
R776 VTAIL.n224 VTAIL.n164 1.93989
R777 VTAIL.n541 VTAIL.n481 1.93989
R778 VTAIL.n509 VTAIL.n508 1.93989
R779 VTAIL.n461 VTAIL.n401 1.93989
R780 VTAIL.n429 VTAIL.n428 1.93989
R781 VTAIL.n383 VTAIL.n323 1.93989
R782 VTAIL.n351 VTAIL.n350 1.93989
R783 VTAIL.n303 VTAIL.n243 1.93989
R784 VTAIL.n271 VTAIL.n270 1.93989
R785 VTAIL.n0 VTAIL.t11 1.40177
R786 VTAIL.n0 VTAIL.t0 1.40177
R787 VTAIL.n158 VTAIL.t4 1.40177
R788 VTAIL.n158 VTAIL.t6 1.40177
R789 VTAIL.n474 VTAIL.t7 1.40177
R790 VTAIL.n474 VTAIL.t8 1.40177
R791 VTAIL.n316 VTAIL.t15 1.40177
R792 VTAIL.n316 VTAIL.t12 1.40177
R793 VTAIL.n582 VTAIL.n576 1.16414
R794 VTAIL.n623 VTAIL.n621 1.16414
R795 VTAIL.n630 VTAIL.n554 1.16414
R796 VTAIL.n30 VTAIL.n24 1.16414
R797 VTAIL.n71 VTAIL.n69 1.16414
R798 VTAIL.n78 VTAIL.n2 1.16414
R799 VTAIL.n108 VTAIL.n102 1.16414
R800 VTAIL.n149 VTAIL.n147 1.16414
R801 VTAIL.n156 VTAIL.n80 1.16414
R802 VTAIL.n188 VTAIL.n182 1.16414
R803 VTAIL.n229 VTAIL.n227 1.16414
R804 VTAIL.n236 VTAIL.n160 1.16414
R805 VTAIL.n552 VTAIL.n476 1.16414
R806 VTAIL.n545 VTAIL.n544 1.16414
R807 VTAIL.n505 VTAIL.n499 1.16414
R808 VTAIL.n472 VTAIL.n396 1.16414
R809 VTAIL.n465 VTAIL.n464 1.16414
R810 VTAIL.n425 VTAIL.n419 1.16414
R811 VTAIL.n394 VTAIL.n318 1.16414
R812 VTAIL.n387 VTAIL.n386 1.16414
R813 VTAIL.n347 VTAIL.n341 1.16414
R814 VTAIL.n314 VTAIL.n238 1.16414
R815 VTAIL.n307 VTAIL.n306 1.16414
R816 VTAIL.n267 VTAIL.n261 1.16414
R817 VTAIL.n317 VTAIL.n315 0.810845
R818 VTAIL.n395 VTAIL.n317 0.810845
R819 VTAIL.n475 VTAIL.n473 0.810845
R820 VTAIL.n553 VTAIL.n475 0.810845
R821 VTAIL.n237 VTAIL.n159 0.810845
R822 VTAIL.n159 VTAIL.n157 0.810845
R823 VTAIL.n79 VTAIL.n1 0.810845
R824 VTAIL VTAIL.n631 0.752655
R825 VTAIL.n473 VTAIL.n395 0.470328
R826 VTAIL.n157 VTAIL.n79 0.470328
R827 VTAIL.n581 VTAIL.n578 0.388379
R828 VTAIL.n622 VTAIL.n556 0.388379
R829 VTAIL.n628 VTAIL.n627 0.388379
R830 VTAIL.n29 VTAIL.n26 0.388379
R831 VTAIL.n70 VTAIL.n4 0.388379
R832 VTAIL.n76 VTAIL.n75 0.388379
R833 VTAIL.n107 VTAIL.n104 0.388379
R834 VTAIL.n148 VTAIL.n82 0.388379
R835 VTAIL.n154 VTAIL.n153 0.388379
R836 VTAIL.n187 VTAIL.n184 0.388379
R837 VTAIL.n228 VTAIL.n162 0.388379
R838 VTAIL.n234 VTAIL.n233 0.388379
R839 VTAIL.n550 VTAIL.n549 0.388379
R840 VTAIL.n480 VTAIL.n478 0.388379
R841 VTAIL.n504 VTAIL.n501 0.388379
R842 VTAIL.n470 VTAIL.n469 0.388379
R843 VTAIL.n400 VTAIL.n398 0.388379
R844 VTAIL.n424 VTAIL.n421 0.388379
R845 VTAIL.n392 VTAIL.n391 0.388379
R846 VTAIL.n322 VTAIL.n320 0.388379
R847 VTAIL.n346 VTAIL.n343 0.388379
R848 VTAIL.n312 VTAIL.n311 0.388379
R849 VTAIL.n242 VTAIL.n240 0.388379
R850 VTAIL.n266 VTAIL.n263 0.388379
R851 VTAIL.n580 VTAIL.n575 0.155672
R852 VTAIL.n587 VTAIL.n575 0.155672
R853 VTAIL.n588 VTAIL.n587 0.155672
R854 VTAIL.n588 VTAIL.n571 0.155672
R855 VTAIL.n595 VTAIL.n571 0.155672
R856 VTAIL.n596 VTAIL.n595 0.155672
R857 VTAIL.n596 VTAIL.n567 0.155672
R858 VTAIL.n603 VTAIL.n567 0.155672
R859 VTAIL.n604 VTAIL.n603 0.155672
R860 VTAIL.n604 VTAIL.n563 0.155672
R861 VTAIL.n611 VTAIL.n563 0.155672
R862 VTAIL.n612 VTAIL.n611 0.155672
R863 VTAIL.n612 VTAIL.n559 0.155672
R864 VTAIL.n619 VTAIL.n559 0.155672
R865 VTAIL.n620 VTAIL.n619 0.155672
R866 VTAIL.n620 VTAIL.n555 0.155672
R867 VTAIL.n629 VTAIL.n555 0.155672
R868 VTAIL.n28 VTAIL.n23 0.155672
R869 VTAIL.n35 VTAIL.n23 0.155672
R870 VTAIL.n36 VTAIL.n35 0.155672
R871 VTAIL.n36 VTAIL.n19 0.155672
R872 VTAIL.n43 VTAIL.n19 0.155672
R873 VTAIL.n44 VTAIL.n43 0.155672
R874 VTAIL.n44 VTAIL.n15 0.155672
R875 VTAIL.n51 VTAIL.n15 0.155672
R876 VTAIL.n52 VTAIL.n51 0.155672
R877 VTAIL.n52 VTAIL.n11 0.155672
R878 VTAIL.n59 VTAIL.n11 0.155672
R879 VTAIL.n60 VTAIL.n59 0.155672
R880 VTAIL.n60 VTAIL.n7 0.155672
R881 VTAIL.n67 VTAIL.n7 0.155672
R882 VTAIL.n68 VTAIL.n67 0.155672
R883 VTAIL.n68 VTAIL.n3 0.155672
R884 VTAIL.n77 VTAIL.n3 0.155672
R885 VTAIL.n106 VTAIL.n101 0.155672
R886 VTAIL.n113 VTAIL.n101 0.155672
R887 VTAIL.n114 VTAIL.n113 0.155672
R888 VTAIL.n114 VTAIL.n97 0.155672
R889 VTAIL.n121 VTAIL.n97 0.155672
R890 VTAIL.n122 VTAIL.n121 0.155672
R891 VTAIL.n122 VTAIL.n93 0.155672
R892 VTAIL.n129 VTAIL.n93 0.155672
R893 VTAIL.n130 VTAIL.n129 0.155672
R894 VTAIL.n130 VTAIL.n89 0.155672
R895 VTAIL.n137 VTAIL.n89 0.155672
R896 VTAIL.n138 VTAIL.n137 0.155672
R897 VTAIL.n138 VTAIL.n85 0.155672
R898 VTAIL.n145 VTAIL.n85 0.155672
R899 VTAIL.n146 VTAIL.n145 0.155672
R900 VTAIL.n146 VTAIL.n81 0.155672
R901 VTAIL.n155 VTAIL.n81 0.155672
R902 VTAIL.n186 VTAIL.n181 0.155672
R903 VTAIL.n193 VTAIL.n181 0.155672
R904 VTAIL.n194 VTAIL.n193 0.155672
R905 VTAIL.n194 VTAIL.n177 0.155672
R906 VTAIL.n201 VTAIL.n177 0.155672
R907 VTAIL.n202 VTAIL.n201 0.155672
R908 VTAIL.n202 VTAIL.n173 0.155672
R909 VTAIL.n209 VTAIL.n173 0.155672
R910 VTAIL.n210 VTAIL.n209 0.155672
R911 VTAIL.n210 VTAIL.n169 0.155672
R912 VTAIL.n217 VTAIL.n169 0.155672
R913 VTAIL.n218 VTAIL.n217 0.155672
R914 VTAIL.n218 VTAIL.n165 0.155672
R915 VTAIL.n225 VTAIL.n165 0.155672
R916 VTAIL.n226 VTAIL.n225 0.155672
R917 VTAIL.n226 VTAIL.n161 0.155672
R918 VTAIL.n235 VTAIL.n161 0.155672
R919 VTAIL.n551 VTAIL.n477 0.155672
R920 VTAIL.n543 VTAIL.n477 0.155672
R921 VTAIL.n543 VTAIL.n542 0.155672
R922 VTAIL.n542 VTAIL.n482 0.155672
R923 VTAIL.n535 VTAIL.n482 0.155672
R924 VTAIL.n535 VTAIL.n534 0.155672
R925 VTAIL.n534 VTAIL.n486 0.155672
R926 VTAIL.n527 VTAIL.n486 0.155672
R927 VTAIL.n527 VTAIL.n526 0.155672
R928 VTAIL.n526 VTAIL.n490 0.155672
R929 VTAIL.n519 VTAIL.n490 0.155672
R930 VTAIL.n519 VTAIL.n518 0.155672
R931 VTAIL.n518 VTAIL.n494 0.155672
R932 VTAIL.n511 VTAIL.n494 0.155672
R933 VTAIL.n511 VTAIL.n510 0.155672
R934 VTAIL.n510 VTAIL.n498 0.155672
R935 VTAIL.n503 VTAIL.n498 0.155672
R936 VTAIL.n471 VTAIL.n397 0.155672
R937 VTAIL.n463 VTAIL.n397 0.155672
R938 VTAIL.n463 VTAIL.n462 0.155672
R939 VTAIL.n462 VTAIL.n402 0.155672
R940 VTAIL.n455 VTAIL.n402 0.155672
R941 VTAIL.n455 VTAIL.n454 0.155672
R942 VTAIL.n454 VTAIL.n406 0.155672
R943 VTAIL.n447 VTAIL.n406 0.155672
R944 VTAIL.n447 VTAIL.n446 0.155672
R945 VTAIL.n446 VTAIL.n410 0.155672
R946 VTAIL.n439 VTAIL.n410 0.155672
R947 VTAIL.n439 VTAIL.n438 0.155672
R948 VTAIL.n438 VTAIL.n414 0.155672
R949 VTAIL.n431 VTAIL.n414 0.155672
R950 VTAIL.n431 VTAIL.n430 0.155672
R951 VTAIL.n430 VTAIL.n418 0.155672
R952 VTAIL.n423 VTAIL.n418 0.155672
R953 VTAIL.n393 VTAIL.n319 0.155672
R954 VTAIL.n385 VTAIL.n319 0.155672
R955 VTAIL.n385 VTAIL.n384 0.155672
R956 VTAIL.n384 VTAIL.n324 0.155672
R957 VTAIL.n377 VTAIL.n324 0.155672
R958 VTAIL.n377 VTAIL.n376 0.155672
R959 VTAIL.n376 VTAIL.n328 0.155672
R960 VTAIL.n369 VTAIL.n328 0.155672
R961 VTAIL.n369 VTAIL.n368 0.155672
R962 VTAIL.n368 VTAIL.n332 0.155672
R963 VTAIL.n361 VTAIL.n332 0.155672
R964 VTAIL.n361 VTAIL.n360 0.155672
R965 VTAIL.n360 VTAIL.n336 0.155672
R966 VTAIL.n353 VTAIL.n336 0.155672
R967 VTAIL.n353 VTAIL.n352 0.155672
R968 VTAIL.n352 VTAIL.n340 0.155672
R969 VTAIL.n345 VTAIL.n340 0.155672
R970 VTAIL.n313 VTAIL.n239 0.155672
R971 VTAIL.n305 VTAIL.n239 0.155672
R972 VTAIL.n305 VTAIL.n304 0.155672
R973 VTAIL.n304 VTAIL.n244 0.155672
R974 VTAIL.n297 VTAIL.n244 0.155672
R975 VTAIL.n297 VTAIL.n296 0.155672
R976 VTAIL.n296 VTAIL.n248 0.155672
R977 VTAIL.n289 VTAIL.n248 0.155672
R978 VTAIL.n289 VTAIL.n288 0.155672
R979 VTAIL.n288 VTAIL.n252 0.155672
R980 VTAIL.n281 VTAIL.n252 0.155672
R981 VTAIL.n281 VTAIL.n280 0.155672
R982 VTAIL.n280 VTAIL.n256 0.155672
R983 VTAIL.n273 VTAIL.n256 0.155672
R984 VTAIL.n273 VTAIL.n272 0.155672
R985 VTAIL.n272 VTAIL.n260 0.155672
R986 VTAIL.n265 VTAIL.n260 0.155672
R987 VTAIL VTAIL.n1 0.0586897
R988 VDD1 VDD1.n0 65.5505
R989 VDD1.n3 VDD1.n2 65.4368
R990 VDD1.n3 VDD1.n1 65.4368
R991 VDD1.n5 VDD1.n4 65.087
R992 VDD1.n5 VDD1.n3 40.1259
R993 VDD1.n4 VDD1.t2 1.40177
R994 VDD1.n4 VDD1.t7 1.40177
R995 VDD1.n0 VDD1.t6 1.40177
R996 VDD1.n0 VDD1.t4 1.40177
R997 VDD1.n2 VDD1.t0 1.40177
R998 VDD1.n2 VDD1.t5 1.40177
R999 VDD1.n1 VDD1.t3 1.40177
R1000 VDD1.n1 VDD1.t1 1.40177
R1001 VDD1 VDD1.n5 0.347483
R1002 B.n174 B.t8 762.486
R1003 B.n168 B.t16 762.486
R1004 B.n69 B.t12 762.486
R1005 B.n75 B.t19 762.486
R1006 B.n505 B.n100 585
R1007 B.n100 B.n43 585
R1008 B.n507 B.n506 585
R1009 B.n509 B.n99 585
R1010 B.n512 B.n511 585
R1011 B.n513 B.n98 585
R1012 B.n515 B.n514 585
R1013 B.n517 B.n97 585
R1014 B.n520 B.n519 585
R1015 B.n521 B.n96 585
R1016 B.n523 B.n522 585
R1017 B.n525 B.n95 585
R1018 B.n528 B.n527 585
R1019 B.n529 B.n94 585
R1020 B.n531 B.n530 585
R1021 B.n533 B.n93 585
R1022 B.n536 B.n535 585
R1023 B.n537 B.n92 585
R1024 B.n539 B.n538 585
R1025 B.n541 B.n91 585
R1026 B.n544 B.n543 585
R1027 B.n545 B.n90 585
R1028 B.n547 B.n546 585
R1029 B.n549 B.n89 585
R1030 B.n552 B.n551 585
R1031 B.n553 B.n88 585
R1032 B.n555 B.n554 585
R1033 B.n557 B.n87 585
R1034 B.n560 B.n559 585
R1035 B.n561 B.n86 585
R1036 B.n563 B.n562 585
R1037 B.n565 B.n85 585
R1038 B.n568 B.n567 585
R1039 B.n569 B.n84 585
R1040 B.n571 B.n570 585
R1041 B.n573 B.n83 585
R1042 B.n576 B.n575 585
R1043 B.n577 B.n82 585
R1044 B.n579 B.n578 585
R1045 B.n581 B.n81 585
R1046 B.n584 B.n583 585
R1047 B.n585 B.n80 585
R1048 B.n587 B.n586 585
R1049 B.n589 B.n79 585
R1050 B.n592 B.n591 585
R1051 B.n593 B.n78 585
R1052 B.n595 B.n594 585
R1053 B.n597 B.n77 585
R1054 B.n600 B.n599 585
R1055 B.n602 B.n74 585
R1056 B.n604 B.n603 585
R1057 B.n606 B.n73 585
R1058 B.n609 B.n608 585
R1059 B.n610 B.n72 585
R1060 B.n612 B.n611 585
R1061 B.n614 B.n71 585
R1062 B.n617 B.n616 585
R1063 B.n618 B.n68 585
R1064 B.n621 B.n620 585
R1065 B.n623 B.n67 585
R1066 B.n626 B.n625 585
R1067 B.n627 B.n66 585
R1068 B.n629 B.n628 585
R1069 B.n631 B.n65 585
R1070 B.n634 B.n633 585
R1071 B.n635 B.n64 585
R1072 B.n637 B.n636 585
R1073 B.n639 B.n63 585
R1074 B.n642 B.n641 585
R1075 B.n643 B.n62 585
R1076 B.n645 B.n644 585
R1077 B.n647 B.n61 585
R1078 B.n650 B.n649 585
R1079 B.n651 B.n60 585
R1080 B.n653 B.n652 585
R1081 B.n655 B.n59 585
R1082 B.n658 B.n657 585
R1083 B.n659 B.n58 585
R1084 B.n661 B.n660 585
R1085 B.n663 B.n57 585
R1086 B.n666 B.n665 585
R1087 B.n667 B.n56 585
R1088 B.n669 B.n668 585
R1089 B.n671 B.n55 585
R1090 B.n674 B.n673 585
R1091 B.n675 B.n54 585
R1092 B.n677 B.n676 585
R1093 B.n679 B.n53 585
R1094 B.n682 B.n681 585
R1095 B.n683 B.n52 585
R1096 B.n685 B.n684 585
R1097 B.n687 B.n51 585
R1098 B.n690 B.n689 585
R1099 B.n691 B.n50 585
R1100 B.n693 B.n692 585
R1101 B.n695 B.n49 585
R1102 B.n698 B.n697 585
R1103 B.n699 B.n48 585
R1104 B.n701 B.n700 585
R1105 B.n703 B.n47 585
R1106 B.n706 B.n705 585
R1107 B.n707 B.n46 585
R1108 B.n709 B.n708 585
R1109 B.n711 B.n45 585
R1110 B.n714 B.n713 585
R1111 B.n715 B.n44 585
R1112 B.n504 B.n42 585
R1113 B.n718 B.n42 585
R1114 B.n503 B.n41 585
R1115 B.n719 B.n41 585
R1116 B.n502 B.n40 585
R1117 B.n720 B.n40 585
R1118 B.n501 B.n500 585
R1119 B.n500 B.n36 585
R1120 B.n499 B.n35 585
R1121 B.n726 B.n35 585
R1122 B.n498 B.n34 585
R1123 B.n727 B.n34 585
R1124 B.n497 B.n33 585
R1125 B.n728 B.n33 585
R1126 B.n496 B.n495 585
R1127 B.n495 B.n29 585
R1128 B.n494 B.n28 585
R1129 B.n734 B.n28 585
R1130 B.n493 B.n27 585
R1131 B.n735 B.n27 585
R1132 B.n492 B.n26 585
R1133 B.n736 B.n26 585
R1134 B.n491 B.n490 585
R1135 B.n490 B.n22 585
R1136 B.n489 B.n21 585
R1137 B.n742 B.n21 585
R1138 B.n488 B.n20 585
R1139 B.n743 B.n20 585
R1140 B.n487 B.n19 585
R1141 B.n744 B.n19 585
R1142 B.n486 B.n485 585
R1143 B.n485 B.n15 585
R1144 B.n484 B.n14 585
R1145 B.n750 B.n14 585
R1146 B.n483 B.n13 585
R1147 B.n751 B.n13 585
R1148 B.n482 B.n12 585
R1149 B.n752 B.n12 585
R1150 B.n481 B.n480 585
R1151 B.n480 B.n11 585
R1152 B.n479 B.n7 585
R1153 B.n758 B.n7 585
R1154 B.n478 B.n6 585
R1155 B.n759 B.n6 585
R1156 B.n477 B.n5 585
R1157 B.n760 B.n5 585
R1158 B.n476 B.n475 585
R1159 B.n475 B.n4 585
R1160 B.n474 B.n101 585
R1161 B.n474 B.n473 585
R1162 B.n463 B.n102 585
R1163 B.n466 B.n102 585
R1164 B.n465 B.n464 585
R1165 B.n467 B.n465 585
R1166 B.n462 B.n107 585
R1167 B.n107 B.n106 585
R1168 B.n461 B.n460 585
R1169 B.n460 B.n459 585
R1170 B.n109 B.n108 585
R1171 B.n110 B.n109 585
R1172 B.n452 B.n451 585
R1173 B.n453 B.n452 585
R1174 B.n450 B.n114 585
R1175 B.n118 B.n114 585
R1176 B.n449 B.n448 585
R1177 B.n448 B.n447 585
R1178 B.n116 B.n115 585
R1179 B.n117 B.n116 585
R1180 B.n440 B.n439 585
R1181 B.n441 B.n440 585
R1182 B.n438 B.n123 585
R1183 B.n123 B.n122 585
R1184 B.n437 B.n436 585
R1185 B.n436 B.n435 585
R1186 B.n125 B.n124 585
R1187 B.n126 B.n125 585
R1188 B.n428 B.n427 585
R1189 B.n429 B.n428 585
R1190 B.n426 B.n131 585
R1191 B.n131 B.n130 585
R1192 B.n425 B.n424 585
R1193 B.n424 B.n423 585
R1194 B.n133 B.n132 585
R1195 B.n134 B.n133 585
R1196 B.n416 B.n415 585
R1197 B.n417 B.n416 585
R1198 B.n414 B.n139 585
R1199 B.n139 B.n138 585
R1200 B.n413 B.n412 585
R1201 B.n412 B.n411 585
R1202 B.n408 B.n143 585
R1203 B.n407 B.n406 585
R1204 B.n404 B.n144 585
R1205 B.n404 B.n142 585
R1206 B.n403 B.n402 585
R1207 B.n401 B.n400 585
R1208 B.n399 B.n146 585
R1209 B.n397 B.n396 585
R1210 B.n395 B.n147 585
R1211 B.n394 B.n393 585
R1212 B.n391 B.n148 585
R1213 B.n389 B.n388 585
R1214 B.n387 B.n149 585
R1215 B.n386 B.n385 585
R1216 B.n383 B.n150 585
R1217 B.n381 B.n380 585
R1218 B.n379 B.n151 585
R1219 B.n378 B.n377 585
R1220 B.n375 B.n152 585
R1221 B.n373 B.n372 585
R1222 B.n371 B.n153 585
R1223 B.n370 B.n369 585
R1224 B.n367 B.n154 585
R1225 B.n365 B.n364 585
R1226 B.n363 B.n155 585
R1227 B.n362 B.n361 585
R1228 B.n359 B.n156 585
R1229 B.n357 B.n356 585
R1230 B.n355 B.n157 585
R1231 B.n354 B.n353 585
R1232 B.n351 B.n158 585
R1233 B.n349 B.n348 585
R1234 B.n347 B.n159 585
R1235 B.n346 B.n345 585
R1236 B.n343 B.n160 585
R1237 B.n341 B.n340 585
R1238 B.n339 B.n161 585
R1239 B.n338 B.n337 585
R1240 B.n335 B.n162 585
R1241 B.n333 B.n332 585
R1242 B.n331 B.n163 585
R1243 B.n330 B.n329 585
R1244 B.n327 B.n164 585
R1245 B.n325 B.n324 585
R1246 B.n323 B.n165 585
R1247 B.n322 B.n321 585
R1248 B.n319 B.n166 585
R1249 B.n317 B.n316 585
R1250 B.n315 B.n167 585
R1251 B.n313 B.n312 585
R1252 B.n310 B.n170 585
R1253 B.n308 B.n307 585
R1254 B.n306 B.n171 585
R1255 B.n305 B.n304 585
R1256 B.n302 B.n172 585
R1257 B.n300 B.n299 585
R1258 B.n298 B.n173 585
R1259 B.n297 B.n296 585
R1260 B.n294 B.n293 585
R1261 B.n292 B.n291 585
R1262 B.n290 B.n178 585
R1263 B.n288 B.n287 585
R1264 B.n286 B.n179 585
R1265 B.n285 B.n284 585
R1266 B.n282 B.n180 585
R1267 B.n280 B.n279 585
R1268 B.n278 B.n181 585
R1269 B.n277 B.n276 585
R1270 B.n274 B.n182 585
R1271 B.n272 B.n271 585
R1272 B.n270 B.n183 585
R1273 B.n269 B.n268 585
R1274 B.n266 B.n184 585
R1275 B.n264 B.n263 585
R1276 B.n262 B.n185 585
R1277 B.n261 B.n260 585
R1278 B.n258 B.n186 585
R1279 B.n256 B.n255 585
R1280 B.n254 B.n187 585
R1281 B.n253 B.n252 585
R1282 B.n250 B.n188 585
R1283 B.n248 B.n247 585
R1284 B.n246 B.n189 585
R1285 B.n245 B.n244 585
R1286 B.n242 B.n190 585
R1287 B.n240 B.n239 585
R1288 B.n238 B.n191 585
R1289 B.n237 B.n236 585
R1290 B.n234 B.n192 585
R1291 B.n232 B.n231 585
R1292 B.n230 B.n193 585
R1293 B.n229 B.n228 585
R1294 B.n226 B.n194 585
R1295 B.n224 B.n223 585
R1296 B.n222 B.n195 585
R1297 B.n221 B.n220 585
R1298 B.n218 B.n196 585
R1299 B.n216 B.n215 585
R1300 B.n214 B.n197 585
R1301 B.n213 B.n212 585
R1302 B.n210 B.n198 585
R1303 B.n208 B.n207 585
R1304 B.n206 B.n199 585
R1305 B.n205 B.n204 585
R1306 B.n202 B.n200 585
R1307 B.n141 B.n140 585
R1308 B.n410 B.n409 585
R1309 B.n411 B.n410 585
R1310 B.n137 B.n136 585
R1311 B.n138 B.n137 585
R1312 B.n419 B.n418 585
R1313 B.n418 B.n417 585
R1314 B.n420 B.n135 585
R1315 B.n135 B.n134 585
R1316 B.n422 B.n421 585
R1317 B.n423 B.n422 585
R1318 B.n129 B.n128 585
R1319 B.n130 B.n129 585
R1320 B.n431 B.n430 585
R1321 B.n430 B.n429 585
R1322 B.n432 B.n127 585
R1323 B.n127 B.n126 585
R1324 B.n434 B.n433 585
R1325 B.n435 B.n434 585
R1326 B.n121 B.n120 585
R1327 B.n122 B.n121 585
R1328 B.n443 B.n442 585
R1329 B.n442 B.n441 585
R1330 B.n444 B.n119 585
R1331 B.n119 B.n117 585
R1332 B.n446 B.n445 585
R1333 B.n447 B.n446 585
R1334 B.n113 B.n112 585
R1335 B.n118 B.n113 585
R1336 B.n455 B.n454 585
R1337 B.n454 B.n453 585
R1338 B.n456 B.n111 585
R1339 B.n111 B.n110 585
R1340 B.n458 B.n457 585
R1341 B.n459 B.n458 585
R1342 B.n105 B.n104 585
R1343 B.n106 B.n105 585
R1344 B.n469 B.n468 585
R1345 B.n468 B.n467 585
R1346 B.n470 B.n103 585
R1347 B.n466 B.n103 585
R1348 B.n472 B.n471 585
R1349 B.n473 B.n472 585
R1350 B.n2 B.n0 585
R1351 B.n4 B.n2 585
R1352 B.n3 B.n1 585
R1353 B.n759 B.n3 585
R1354 B.n757 B.n756 585
R1355 B.n758 B.n757 585
R1356 B.n755 B.n8 585
R1357 B.n11 B.n8 585
R1358 B.n754 B.n753 585
R1359 B.n753 B.n752 585
R1360 B.n10 B.n9 585
R1361 B.n751 B.n10 585
R1362 B.n749 B.n748 585
R1363 B.n750 B.n749 585
R1364 B.n747 B.n16 585
R1365 B.n16 B.n15 585
R1366 B.n746 B.n745 585
R1367 B.n745 B.n744 585
R1368 B.n18 B.n17 585
R1369 B.n743 B.n18 585
R1370 B.n741 B.n740 585
R1371 B.n742 B.n741 585
R1372 B.n739 B.n23 585
R1373 B.n23 B.n22 585
R1374 B.n738 B.n737 585
R1375 B.n737 B.n736 585
R1376 B.n25 B.n24 585
R1377 B.n735 B.n25 585
R1378 B.n733 B.n732 585
R1379 B.n734 B.n733 585
R1380 B.n731 B.n30 585
R1381 B.n30 B.n29 585
R1382 B.n730 B.n729 585
R1383 B.n729 B.n728 585
R1384 B.n32 B.n31 585
R1385 B.n727 B.n32 585
R1386 B.n725 B.n724 585
R1387 B.n726 B.n725 585
R1388 B.n723 B.n37 585
R1389 B.n37 B.n36 585
R1390 B.n722 B.n721 585
R1391 B.n721 B.n720 585
R1392 B.n39 B.n38 585
R1393 B.n719 B.n39 585
R1394 B.n717 B.n716 585
R1395 B.n718 B.n717 585
R1396 B.n762 B.n761 585
R1397 B.n761 B.n760 585
R1398 B.n410 B.n143 516.524
R1399 B.n717 B.n44 516.524
R1400 B.n412 B.n141 516.524
R1401 B.n100 B.n42 516.524
R1402 B.n174 B.t11 337.122
R1403 B.n75 B.t20 337.122
R1404 B.n168 B.t18 337.122
R1405 B.n69 B.t14 337.122
R1406 B.n175 B.t10 318.89
R1407 B.n76 B.t21 318.89
R1408 B.n169 B.t17 318.89
R1409 B.n70 B.t15 318.89
R1410 B.n508 B.n43 256.663
R1411 B.n510 B.n43 256.663
R1412 B.n516 B.n43 256.663
R1413 B.n518 B.n43 256.663
R1414 B.n524 B.n43 256.663
R1415 B.n526 B.n43 256.663
R1416 B.n532 B.n43 256.663
R1417 B.n534 B.n43 256.663
R1418 B.n540 B.n43 256.663
R1419 B.n542 B.n43 256.663
R1420 B.n548 B.n43 256.663
R1421 B.n550 B.n43 256.663
R1422 B.n556 B.n43 256.663
R1423 B.n558 B.n43 256.663
R1424 B.n564 B.n43 256.663
R1425 B.n566 B.n43 256.663
R1426 B.n572 B.n43 256.663
R1427 B.n574 B.n43 256.663
R1428 B.n580 B.n43 256.663
R1429 B.n582 B.n43 256.663
R1430 B.n588 B.n43 256.663
R1431 B.n590 B.n43 256.663
R1432 B.n596 B.n43 256.663
R1433 B.n598 B.n43 256.663
R1434 B.n605 B.n43 256.663
R1435 B.n607 B.n43 256.663
R1436 B.n613 B.n43 256.663
R1437 B.n615 B.n43 256.663
R1438 B.n622 B.n43 256.663
R1439 B.n624 B.n43 256.663
R1440 B.n630 B.n43 256.663
R1441 B.n632 B.n43 256.663
R1442 B.n638 B.n43 256.663
R1443 B.n640 B.n43 256.663
R1444 B.n646 B.n43 256.663
R1445 B.n648 B.n43 256.663
R1446 B.n654 B.n43 256.663
R1447 B.n656 B.n43 256.663
R1448 B.n662 B.n43 256.663
R1449 B.n664 B.n43 256.663
R1450 B.n670 B.n43 256.663
R1451 B.n672 B.n43 256.663
R1452 B.n678 B.n43 256.663
R1453 B.n680 B.n43 256.663
R1454 B.n686 B.n43 256.663
R1455 B.n688 B.n43 256.663
R1456 B.n694 B.n43 256.663
R1457 B.n696 B.n43 256.663
R1458 B.n702 B.n43 256.663
R1459 B.n704 B.n43 256.663
R1460 B.n710 B.n43 256.663
R1461 B.n712 B.n43 256.663
R1462 B.n405 B.n142 256.663
R1463 B.n145 B.n142 256.663
R1464 B.n398 B.n142 256.663
R1465 B.n392 B.n142 256.663
R1466 B.n390 B.n142 256.663
R1467 B.n384 B.n142 256.663
R1468 B.n382 B.n142 256.663
R1469 B.n376 B.n142 256.663
R1470 B.n374 B.n142 256.663
R1471 B.n368 B.n142 256.663
R1472 B.n366 B.n142 256.663
R1473 B.n360 B.n142 256.663
R1474 B.n358 B.n142 256.663
R1475 B.n352 B.n142 256.663
R1476 B.n350 B.n142 256.663
R1477 B.n344 B.n142 256.663
R1478 B.n342 B.n142 256.663
R1479 B.n336 B.n142 256.663
R1480 B.n334 B.n142 256.663
R1481 B.n328 B.n142 256.663
R1482 B.n326 B.n142 256.663
R1483 B.n320 B.n142 256.663
R1484 B.n318 B.n142 256.663
R1485 B.n311 B.n142 256.663
R1486 B.n309 B.n142 256.663
R1487 B.n303 B.n142 256.663
R1488 B.n301 B.n142 256.663
R1489 B.n295 B.n142 256.663
R1490 B.n177 B.n142 256.663
R1491 B.n289 B.n142 256.663
R1492 B.n283 B.n142 256.663
R1493 B.n281 B.n142 256.663
R1494 B.n275 B.n142 256.663
R1495 B.n273 B.n142 256.663
R1496 B.n267 B.n142 256.663
R1497 B.n265 B.n142 256.663
R1498 B.n259 B.n142 256.663
R1499 B.n257 B.n142 256.663
R1500 B.n251 B.n142 256.663
R1501 B.n249 B.n142 256.663
R1502 B.n243 B.n142 256.663
R1503 B.n241 B.n142 256.663
R1504 B.n235 B.n142 256.663
R1505 B.n233 B.n142 256.663
R1506 B.n227 B.n142 256.663
R1507 B.n225 B.n142 256.663
R1508 B.n219 B.n142 256.663
R1509 B.n217 B.n142 256.663
R1510 B.n211 B.n142 256.663
R1511 B.n209 B.n142 256.663
R1512 B.n203 B.n142 256.663
R1513 B.n201 B.n142 256.663
R1514 B.n410 B.n137 163.367
R1515 B.n418 B.n137 163.367
R1516 B.n418 B.n135 163.367
R1517 B.n422 B.n135 163.367
R1518 B.n422 B.n129 163.367
R1519 B.n430 B.n129 163.367
R1520 B.n430 B.n127 163.367
R1521 B.n434 B.n127 163.367
R1522 B.n434 B.n121 163.367
R1523 B.n442 B.n121 163.367
R1524 B.n442 B.n119 163.367
R1525 B.n446 B.n119 163.367
R1526 B.n446 B.n113 163.367
R1527 B.n454 B.n113 163.367
R1528 B.n454 B.n111 163.367
R1529 B.n458 B.n111 163.367
R1530 B.n458 B.n105 163.367
R1531 B.n468 B.n105 163.367
R1532 B.n468 B.n103 163.367
R1533 B.n472 B.n103 163.367
R1534 B.n472 B.n2 163.367
R1535 B.n761 B.n2 163.367
R1536 B.n761 B.n3 163.367
R1537 B.n757 B.n3 163.367
R1538 B.n757 B.n8 163.367
R1539 B.n753 B.n8 163.367
R1540 B.n753 B.n10 163.367
R1541 B.n749 B.n10 163.367
R1542 B.n749 B.n16 163.367
R1543 B.n745 B.n16 163.367
R1544 B.n745 B.n18 163.367
R1545 B.n741 B.n18 163.367
R1546 B.n741 B.n23 163.367
R1547 B.n737 B.n23 163.367
R1548 B.n737 B.n25 163.367
R1549 B.n733 B.n25 163.367
R1550 B.n733 B.n30 163.367
R1551 B.n729 B.n30 163.367
R1552 B.n729 B.n32 163.367
R1553 B.n725 B.n32 163.367
R1554 B.n725 B.n37 163.367
R1555 B.n721 B.n37 163.367
R1556 B.n721 B.n39 163.367
R1557 B.n717 B.n39 163.367
R1558 B.n406 B.n404 163.367
R1559 B.n404 B.n403 163.367
R1560 B.n400 B.n399 163.367
R1561 B.n397 B.n147 163.367
R1562 B.n393 B.n391 163.367
R1563 B.n389 B.n149 163.367
R1564 B.n385 B.n383 163.367
R1565 B.n381 B.n151 163.367
R1566 B.n377 B.n375 163.367
R1567 B.n373 B.n153 163.367
R1568 B.n369 B.n367 163.367
R1569 B.n365 B.n155 163.367
R1570 B.n361 B.n359 163.367
R1571 B.n357 B.n157 163.367
R1572 B.n353 B.n351 163.367
R1573 B.n349 B.n159 163.367
R1574 B.n345 B.n343 163.367
R1575 B.n341 B.n161 163.367
R1576 B.n337 B.n335 163.367
R1577 B.n333 B.n163 163.367
R1578 B.n329 B.n327 163.367
R1579 B.n325 B.n165 163.367
R1580 B.n321 B.n319 163.367
R1581 B.n317 B.n167 163.367
R1582 B.n312 B.n310 163.367
R1583 B.n308 B.n171 163.367
R1584 B.n304 B.n302 163.367
R1585 B.n300 B.n173 163.367
R1586 B.n296 B.n294 163.367
R1587 B.n291 B.n290 163.367
R1588 B.n288 B.n179 163.367
R1589 B.n284 B.n282 163.367
R1590 B.n280 B.n181 163.367
R1591 B.n276 B.n274 163.367
R1592 B.n272 B.n183 163.367
R1593 B.n268 B.n266 163.367
R1594 B.n264 B.n185 163.367
R1595 B.n260 B.n258 163.367
R1596 B.n256 B.n187 163.367
R1597 B.n252 B.n250 163.367
R1598 B.n248 B.n189 163.367
R1599 B.n244 B.n242 163.367
R1600 B.n240 B.n191 163.367
R1601 B.n236 B.n234 163.367
R1602 B.n232 B.n193 163.367
R1603 B.n228 B.n226 163.367
R1604 B.n224 B.n195 163.367
R1605 B.n220 B.n218 163.367
R1606 B.n216 B.n197 163.367
R1607 B.n212 B.n210 163.367
R1608 B.n208 B.n199 163.367
R1609 B.n204 B.n202 163.367
R1610 B.n412 B.n139 163.367
R1611 B.n416 B.n139 163.367
R1612 B.n416 B.n133 163.367
R1613 B.n424 B.n133 163.367
R1614 B.n424 B.n131 163.367
R1615 B.n428 B.n131 163.367
R1616 B.n428 B.n125 163.367
R1617 B.n436 B.n125 163.367
R1618 B.n436 B.n123 163.367
R1619 B.n440 B.n123 163.367
R1620 B.n440 B.n116 163.367
R1621 B.n448 B.n116 163.367
R1622 B.n448 B.n114 163.367
R1623 B.n452 B.n114 163.367
R1624 B.n452 B.n109 163.367
R1625 B.n460 B.n109 163.367
R1626 B.n460 B.n107 163.367
R1627 B.n465 B.n107 163.367
R1628 B.n465 B.n102 163.367
R1629 B.n474 B.n102 163.367
R1630 B.n475 B.n474 163.367
R1631 B.n475 B.n5 163.367
R1632 B.n6 B.n5 163.367
R1633 B.n7 B.n6 163.367
R1634 B.n480 B.n7 163.367
R1635 B.n480 B.n12 163.367
R1636 B.n13 B.n12 163.367
R1637 B.n14 B.n13 163.367
R1638 B.n485 B.n14 163.367
R1639 B.n485 B.n19 163.367
R1640 B.n20 B.n19 163.367
R1641 B.n21 B.n20 163.367
R1642 B.n490 B.n21 163.367
R1643 B.n490 B.n26 163.367
R1644 B.n27 B.n26 163.367
R1645 B.n28 B.n27 163.367
R1646 B.n495 B.n28 163.367
R1647 B.n495 B.n33 163.367
R1648 B.n34 B.n33 163.367
R1649 B.n35 B.n34 163.367
R1650 B.n500 B.n35 163.367
R1651 B.n500 B.n40 163.367
R1652 B.n41 B.n40 163.367
R1653 B.n42 B.n41 163.367
R1654 B.n713 B.n711 163.367
R1655 B.n709 B.n46 163.367
R1656 B.n705 B.n703 163.367
R1657 B.n701 B.n48 163.367
R1658 B.n697 B.n695 163.367
R1659 B.n693 B.n50 163.367
R1660 B.n689 B.n687 163.367
R1661 B.n685 B.n52 163.367
R1662 B.n681 B.n679 163.367
R1663 B.n677 B.n54 163.367
R1664 B.n673 B.n671 163.367
R1665 B.n669 B.n56 163.367
R1666 B.n665 B.n663 163.367
R1667 B.n661 B.n58 163.367
R1668 B.n657 B.n655 163.367
R1669 B.n653 B.n60 163.367
R1670 B.n649 B.n647 163.367
R1671 B.n645 B.n62 163.367
R1672 B.n641 B.n639 163.367
R1673 B.n637 B.n64 163.367
R1674 B.n633 B.n631 163.367
R1675 B.n629 B.n66 163.367
R1676 B.n625 B.n623 163.367
R1677 B.n621 B.n68 163.367
R1678 B.n616 B.n614 163.367
R1679 B.n612 B.n72 163.367
R1680 B.n608 B.n606 163.367
R1681 B.n604 B.n74 163.367
R1682 B.n599 B.n597 163.367
R1683 B.n595 B.n78 163.367
R1684 B.n591 B.n589 163.367
R1685 B.n587 B.n80 163.367
R1686 B.n583 B.n581 163.367
R1687 B.n579 B.n82 163.367
R1688 B.n575 B.n573 163.367
R1689 B.n571 B.n84 163.367
R1690 B.n567 B.n565 163.367
R1691 B.n563 B.n86 163.367
R1692 B.n559 B.n557 163.367
R1693 B.n555 B.n88 163.367
R1694 B.n551 B.n549 163.367
R1695 B.n547 B.n90 163.367
R1696 B.n543 B.n541 163.367
R1697 B.n539 B.n92 163.367
R1698 B.n535 B.n533 163.367
R1699 B.n531 B.n94 163.367
R1700 B.n527 B.n525 163.367
R1701 B.n523 B.n96 163.367
R1702 B.n519 B.n517 163.367
R1703 B.n515 B.n98 163.367
R1704 B.n511 B.n509 163.367
R1705 B.n507 B.n100 163.367
R1706 B.n405 B.n143 71.676
R1707 B.n403 B.n145 71.676
R1708 B.n399 B.n398 71.676
R1709 B.n392 B.n147 71.676
R1710 B.n391 B.n390 71.676
R1711 B.n384 B.n149 71.676
R1712 B.n383 B.n382 71.676
R1713 B.n376 B.n151 71.676
R1714 B.n375 B.n374 71.676
R1715 B.n368 B.n153 71.676
R1716 B.n367 B.n366 71.676
R1717 B.n360 B.n155 71.676
R1718 B.n359 B.n358 71.676
R1719 B.n352 B.n157 71.676
R1720 B.n351 B.n350 71.676
R1721 B.n344 B.n159 71.676
R1722 B.n343 B.n342 71.676
R1723 B.n336 B.n161 71.676
R1724 B.n335 B.n334 71.676
R1725 B.n328 B.n163 71.676
R1726 B.n327 B.n326 71.676
R1727 B.n320 B.n165 71.676
R1728 B.n319 B.n318 71.676
R1729 B.n311 B.n167 71.676
R1730 B.n310 B.n309 71.676
R1731 B.n303 B.n171 71.676
R1732 B.n302 B.n301 71.676
R1733 B.n295 B.n173 71.676
R1734 B.n294 B.n177 71.676
R1735 B.n290 B.n289 71.676
R1736 B.n283 B.n179 71.676
R1737 B.n282 B.n281 71.676
R1738 B.n275 B.n181 71.676
R1739 B.n274 B.n273 71.676
R1740 B.n267 B.n183 71.676
R1741 B.n266 B.n265 71.676
R1742 B.n259 B.n185 71.676
R1743 B.n258 B.n257 71.676
R1744 B.n251 B.n187 71.676
R1745 B.n250 B.n249 71.676
R1746 B.n243 B.n189 71.676
R1747 B.n242 B.n241 71.676
R1748 B.n235 B.n191 71.676
R1749 B.n234 B.n233 71.676
R1750 B.n227 B.n193 71.676
R1751 B.n226 B.n225 71.676
R1752 B.n219 B.n195 71.676
R1753 B.n218 B.n217 71.676
R1754 B.n211 B.n197 71.676
R1755 B.n210 B.n209 71.676
R1756 B.n203 B.n199 71.676
R1757 B.n202 B.n201 71.676
R1758 B.n712 B.n44 71.676
R1759 B.n711 B.n710 71.676
R1760 B.n704 B.n46 71.676
R1761 B.n703 B.n702 71.676
R1762 B.n696 B.n48 71.676
R1763 B.n695 B.n694 71.676
R1764 B.n688 B.n50 71.676
R1765 B.n687 B.n686 71.676
R1766 B.n680 B.n52 71.676
R1767 B.n679 B.n678 71.676
R1768 B.n672 B.n54 71.676
R1769 B.n671 B.n670 71.676
R1770 B.n664 B.n56 71.676
R1771 B.n663 B.n662 71.676
R1772 B.n656 B.n58 71.676
R1773 B.n655 B.n654 71.676
R1774 B.n648 B.n60 71.676
R1775 B.n647 B.n646 71.676
R1776 B.n640 B.n62 71.676
R1777 B.n639 B.n638 71.676
R1778 B.n632 B.n64 71.676
R1779 B.n631 B.n630 71.676
R1780 B.n624 B.n66 71.676
R1781 B.n623 B.n622 71.676
R1782 B.n615 B.n68 71.676
R1783 B.n614 B.n613 71.676
R1784 B.n607 B.n72 71.676
R1785 B.n606 B.n605 71.676
R1786 B.n598 B.n74 71.676
R1787 B.n597 B.n596 71.676
R1788 B.n590 B.n78 71.676
R1789 B.n589 B.n588 71.676
R1790 B.n582 B.n80 71.676
R1791 B.n581 B.n580 71.676
R1792 B.n574 B.n82 71.676
R1793 B.n573 B.n572 71.676
R1794 B.n566 B.n84 71.676
R1795 B.n565 B.n564 71.676
R1796 B.n558 B.n86 71.676
R1797 B.n557 B.n556 71.676
R1798 B.n550 B.n88 71.676
R1799 B.n549 B.n548 71.676
R1800 B.n542 B.n90 71.676
R1801 B.n541 B.n540 71.676
R1802 B.n534 B.n92 71.676
R1803 B.n533 B.n532 71.676
R1804 B.n526 B.n94 71.676
R1805 B.n525 B.n524 71.676
R1806 B.n518 B.n96 71.676
R1807 B.n517 B.n516 71.676
R1808 B.n510 B.n98 71.676
R1809 B.n509 B.n508 71.676
R1810 B.n508 B.n507 71.676
R1811 B.n511 B.n510 71.676
R1812 B.n516 B.n515 71.676
R1813 B.n519 B.n518 71.676
R1814 B.n524 B.n523 71.676
R1815 B.n527 B.n526 71.676
R1816 B.n532 B.n531 71.676
R1817 B.n535 B.n534 71.676
R1818 B.n540 B.n539 71.676
R1819 B.n543 B.n542 71.676
R1820 B.n548 B.n547 71.676
R1821 B.n551 B.n550 71.676
R1822 B.n556 B.n555 71.676
R1823 B.n559 B.n558 71.676
R1824 B.n564 B.n563 71.676
R1825 B.n567 B.n566 71.676
R1826 B.n572 B.n571 71.676
R1827 B.n575 B.n574 71.676
R1828 B.n580 B.n579 71.676
R1829 B.n583 B.n582 71.676
R1830 B.n588 B.n587 71.676
R1831 B.n591 B.n590 71.676
R1832 B.n596 B.n595 71.676
R1833 B.n599 B.n598 71.676
R1834 B.n605 B.n604 71.676
R1835 B.n608 B.n607 71.676
R1836 B.n613 B.n612 71.676
R1837 B.n616 B.n615 71.676
R1838 B.n622 B.n621 71.676
R1839 B.n625 B.n624 71.676
R1840 B.n630 B.n629 71.676
R1841 B.n633 B.n632 71.676
R1842 B.n638 B.n637 71.676
R1843 B.n641 B.n640 71.676
R1844 B.n646 B.n645 71.676
R1845 B.n649 B.n648 71.676
R1846 B.n654 B.n653 71.676
R1847 B.n657 B.n656 71.676
R1848 B.n662 B.n661 71.676
R1849 B.n665 B.n664 71.676
R1850 B.n670 B.n669 71.676
R1851 B.n673 B.n672 71.676
R1852 B.n678 B.n677 71.676
R1853 B.n681 B.n680 71.676
R1854 B.n686 B.n685 71.676
R1855 B.n689 B.n688 71.676
R1856 B.n694 B.n693 71.676
R1857 B.n697 B.n696 71.676
R1858 B.n702 B.n701 71.676
R1859 B.n705 B.n704 71.676
R1860 B.n710 B.n709 71.676
R1861 B.n713 B.n712 71.676
R1862 B.n406 B.n405 71.676
R1863 B.n400 B.n145 71.676
R1864 B.n398 B.n397 71.676
R1865 B.n393 B.n392 71.676
R1866 B.n390 B.n389 71.676
R1867 B.n385 B.n384 71.676
R1868 B.n382 B.n381 71.676
R1869 B.n377 B.n376 71.676
R1870 B.n374 B.n373 71.676
R1871 B.n369 B.n368 71.676
R1872 B.n366 B.n365 71.676
R1873 B.n361 B.n360 71.676
R1874 B.n358 B.n357 71.676
R1875 B.n353 B.n352 71.676
R1876 B.n350 B.n349 71.676
R1877 B.n345 B.n344 71.676
R1878 B.n342 B.n341 71.676
R1879 B.n337 B.n336 71.676
R1880 B.n334 B.n333 71.676
R1881 B.n329 B.n328 71.676
R1882 B.n326 B.n325 71.676
R1883 B.n321 B.n320 71.676
R1884 B.n318 B.n317 71.676
R1885 B.n312 B.n311 71.676
R1886 B.n309 B.n308 71.676
R1887 B.n304 B.n303 71.676
R1888 B.n301 B.n300 71.676
R1889 B.n296 B.n295 71.676
R1890 B.n291 B.n177 71.676
R1891 B.n289 B.n288 71.676
R1892 B.n284 B.n283 71.676
R1893 B.n281 B.n280 71.676
R1894 B.n276 B.n275 71.676
R1895 B.n273 B.n272 71.676
R1896 B.n268 B.n267 71.676
R1897 B.n265 B.n264 71.676
R1898 B.n260 B.n259 71.676
R1899 B.n257 B.n256 71.676
R1900 B.n252 B.n251 71.676
R1901 B.n249 B.n248 71.676
R1902 B.n244 B.n243 71.676
R1903 B.n241 B.n240 71.676
R1904 B.n236 B.n235 71.676
R1905 B.n233 B.n232 71.676
R1906 B.n228 B.n227 71.676
R1907 B.n225 B.n224 71.676
R1908 B.n220 B.n219 71.676
R1909 B.n217 B.n216 71.676
R1910 B.n212 B.n211 71.676
R1911 B.n209 B.n208 71.676
R1912 B.n204 B.n203 71.676
R1913 B.n201 B.n141 71.676
R1914 B.n411 B.n142 67.4573
R1915 B.n718 B.n43 67.4573
R1916 B.n176 B.n175 59.5399
R1917 B.n314 B.n169 59.5399
R1918 B.n619 B.n70 59.5399
R1919 B.n601 B.n76 59.5399
R1920 B.n411 B.n138 38.5473
R1921 B.n417 B.n138 38.5473
R1922 B.n417 B.n134 38.5473
R1923 B.n423 B.n134 38.5473
R1924 B.n429 B.n130 38.5473
R1925 B.n429 B.n126 38.5473
R1926 B.n435 B.n126 38.5473
R1927 B.n435 B.n122 38.5473
R1928 B.n441 B.n122 38.5473
R1929 B.n447 B.n117 38.5473
R1930 B.n447 B.n118 38.5473
R1931 B.n453 B.n110 38.5473
R1932 B.n459 B.n110 38.5473
R1933 B.n467 B.n106 38.5473
R1934 B.n467 B.n466 38.5473
R1935 B.n473 B.n4 38.5473
R1936 B.n760 B.n4 38.5473
R1937 B.n760 B.n759 38.5473
R1938 B.n759 B.n758 38.5473
R1939 B.n752 B.n11 38.5473
R1940 B.n752 B.n751 38.5473
R1941 B.n750 B.n15 38.5473
R1942 B.n744 B.n15 38.5473
R1943 B.n743 B.n742 38.5473
R1944 B.n742 B.n22 38.5473
R1945 B.n736 B.n735 38.5473
R1946 B.n735 B.n734 38.5473
R1947 B.n734 B.n29 38.5473
R1948 B.n728 B.n29 38.5473
R1949 B.n728 B.n727 38.5473
R1950 B.n726 B.n36 38.5473
R1951 B.n720 B.n36 38.5473
R1952 B.n720 B.n719 38.5473
R1953 B.n719 B.n718 38.5473
R1954 B.n473 B.t6 37.9804
R1955 B.n758 B.t7 37.9804
R1956 B.n716 B.n715 33.5615
R1957 B.n505 B.n504 33.5615
R1958 B.n413 B.n140 33.5615
R1959 B.n409 B.n408 33.5615
R1960 B.n423 B.t9 28.9106
R1961 B.t2 B.n106 28.9106
R1962 B.n751 B.t5 28.9106
R1963 B.t13 B.n726 28.9106
R1964 B.n441 B.t4 27.7768
R1965 B.n736 B.t1 27.7768
R1966 B.n453 B.t3 19.8407
R1967 B.n744 B.t0 19.8407
R1968 B.n118 B.t3 18.707
R1969 B.t0 B.n743 18.707
R1970 B.n175 B.n174 18.2308
R1971 B.n169 B.n168 18.2308
R1972 B.n70 B.n69 18.2308
R1973 B.n76 B.n75 18.2308
R1974 B B.n762 18.0485
R1975 B.t4 B.n117 10.7709
R1976 B.t1 B.n22 10.7709
R1977 B.n715 B.n714 10.6151
R1978 B.n714 B.n45 10.6151
R1979 B.n708 B.n45 10.6151
R1980 B.n708 B.n707 10.6151
R1981 B.n707 B.n706 10.6151
R1982 B.n706 B.n47 10.6151
R1983 B.n700 B.n47 10.6151
R1984 B.n700 B.n699 10.6151
R1985 B.n699 B.n698 10.6151
R1986 B.n698 B.n49 10.6151
R1987 B.n692 B.n49 10.6151
R1988 B.n692 B.n691 10.6151
R1989 B.n691 B.n690 10.6151
R1990 B.n690 B.n51 10.6151
R1991 B.n684 B.n51 10.6151
R1992 B.n684 B.n683 10.6151
R1993 B.n683 B.n682 10.6151
R1994 B.n682 B.n53 10.6151
R1995 B.n676 B.n53 10.6151
R1996 B.n676 B.n675 10.6151
R1997 B.n675 B.n674 10.6151
R1998 B.n674 B.n55 10.6151
R1999 B.n668 B.n55 10.6151
R2000 B.n668 B.n667 10.6151
R2001 B.n667 B.n666 10.6151
R2002 B.n666 B.n57 10.6151
R2003 B.n660 B.n57 10.6151
R2004 B.n660 B.n659 10.6151
R2005 B.n659 B.n658 10.6151
R2006 B.n658 B.n59 10.6151
R2007 B.n652 B.n59 10.6151
R2008 B.n652 B.n651 10.6151
R2009 B.n651 B.n650 10.6151
R2010 B.n650 B.n61 10.6151
R2011 B.n644 B.n61 10.6151
R2012 B.n644 B.n643 10.6151
R2013 B.n643 B.n642 10.6151
R2014 B.n642 B.n63 10.6151
R2015 B.n636 B.n63 10.6151
R2016 B.n636 B.n635 10.6151
R2017 B.n635 B.n634 10.6151
R2018 B.n634 B.n65 10.6151
R2019 B.n628 B.n65 10.6151
R2020 B.n628 B.n627 10.6151
R2021 B.n627 B.n626 10.6151
R2022 B.n626 B.n67 10.6151
R2023 B.n620 B.n67 10.6151
R2024 B.n618 B.n617 10.6151
R2025 B.n617 B.n71 10.6151
R2026 B.n611 B.n71 10.6151
R2027 B.n611 B.n610 10.6151
R2028 B.n610 B.n609 10.6151
R2029 B.n609 B.n73 10.6151
R2030 B.n603 B.n73 10.6151
R2031 B.n603 B.n602 10.6151
R2032 B.n600 B.n77 10.6151
R2033 B.n594 B.n77 10.6151
R2034 B.n594 B.n593 10.6151
R2035 B.n593 B.n592 10.6151
R2036 B.n592 B.n79 10.6151
R2037 B.n586 B.n79 10.6151
R2038 B.n586 B.n585 10.6151
R2039 B.n585 B.n584 10.6151
R2040 B.n584 B.n81 10.6151
R2041 B.n578 B.n81 10.6151
R2042 B.n578 B.n577 10.6151
R2043 B.n577 B.n576 10.6151
R2044 B.n576 B.n83 10.6151
R2045 B.n570 B.n83 10.6151
R2046 B.n570 B.n569 10.6151
R2047 B.n569 B.n568 10.6151
R2048 B.n568 B.n85 10.6151
R2049 B.n562 B.n85 10.6151
R2050 B.n562 B.n561 10.6151
R2051 B.n561 B.n560 10.6151
R2052 B.n560 B.n87 10.6151
R2053 B.n554 B.n87 10.6151
R2054 B.n554 B.n553 10.6151
R2055 B.n553 B.n552 10.6151
R2056 B.n552 B.n89 10.6151
R2057 B.n546 B.n89 10.6151
R2058 B.n546 B.n545 10.6151
R2059 B.n545 B.n544 10.6151
R2060 B.n544 B.n91 10.6151
R2061 B.n538 B.n91 10.6151
R2062 B.n538 B.n537 10.6151
R2063 B.n537 B.n536 10.6151
R2064 B.n536 B.n93 10.6151
R2065 B.n530 B.n93 10.6151
R2066 B.n530 B.n529 10.6151
R2067 B.n529 B.n528 10.6151
R2068 B.n528 B.n95 10.6151
R2069 B.n522 B.n95 10.6151
R2070 B.n522 B.n521 10.6151
R2071 B.n521 B.n520 10.6151
R2072 B.n520 B.n97 10.6151
R2073 B.n514 B.n97 10.6151
R2074 B.n514 B.n513 10.6151
R2075 B.n513 B.n512 10.6151
R2076 B.n512 B.n99 10.6151
R2077 B.n506 B.n99 10.6151
R2078 B.n506 B.n505 10.6151
R2079 B.n414 B.n413 10.6151
R2080 B.n415 B.n414 10.6151
R2081 B.n415 B.n132 10.6151
R2082 B.n425 B.n132 10.6151
R2083 B.n426 B.n425 10.6151
R2084 B.n427 B.n426 10.6151
R2085 B.n427 B.n124 10.6151
R2086 B.n437 B.n124 10.6151
R2087 B.n438 B.n437 10.6151
R2088 B.n439 B.n438 10.6151
R2089 B.n439 B.n115 10.6151
R2090 B.n449 B.n115 10.6151
R2091 B.n450 B.n449 10.6151
R2092 B.n451 B.n450 10.6151
R2093 B.n451 B.n108 10.6151
R2094 B.n461 B.n108 10.6151
R2095 B.n462 B.n461 10.6151
R2096 B.n464 B.n462 10.6151
R2097 B.n464 B.n463 10.6151
R2098 B.n463 B.n101 10.6151
R2099 B.n476 B.n101 10.6151
R2100 B.n477 B.n476 10.6151
R2101 B.n478 B.n477 10.6151
R2102 B.n479 B.n478 10.6151
R2103 B.n481 B.n479 10.6151
R2104 B.n482 B.n481 10.6151
R2105 B.n483 B.n482 10.6151
R2106 B.n484 B.n483 10.6151
R2107 B.n486 B.n484 10.6151
R2108 B.n487 B.n486 10.6151
R2109 B.n488 B.n487 10.6151
R2110 B.n489 B.n488 10.6151
R2111 B.n491 B.n489 10.6151
R2112 B.n492 B.n491 10.6151
R2113 B.n493 B.n492 10.6151
R2114 B.n494 B.n493 10.6151
R2115 B.n496 B.n494 10.6151
R2116 B.n497 B.n496 10.6151
R2117 B.n498 B.n497 10.6151
R2118 B.n499 B.n498 10.6151
R2119 B.n501 B.n499 10.6151
R2120 B.n502 B.n501 10.6151
R2121 B.n503 B.n502 10.6151
R2122 B.n504 B.n503 10.6151
R2123 B.n408 B.n407 10.6151
R2124 B.n407 B.n144 10.6151
R2125 B.n402 B.n144 10.6151
R2126 B.n402 B.n401 10.6151
R2127 B.n401 B.n146 10.6151
R2128 B.n396 B.n146 10.6151
R2129 B.n396 B.n395 10.6151
R2130 B.n395 B.n394 10.6151
R2131 B.n394 B.n148 10.6151
R2132 B.n388 B.n148 10.6151
R2133 B.n388 B.n387 10.6151
R2134 B.n387 B.n386 10.6151
R2135 B.n386 B.n150 10.6151
R2136 B.n380 B.n150 10.6151
R2137 B.n380 B.n379 10.6151
R2138 B.n379 B.n378 10.6151
R2139 B.n378 B.n152 10.6151
R2140 B.n372 B.n152 10.6151
R2141 B.n372 B.n371 10.6151
R2142 B.n371 B.n370 10.6151
R2143 B.n370 B.n154 10.6151
R2144 B.n364 B.n154 10.6151
R2145 B.n364 B.n363 10.6151
R2146 B.n363 B.n362 10.6151
R2147 B.n362 B.n156 10.6151
R2148 B.n356 B.n156 10.6151
R2149 B.n356 B.n355 10.6151
R2150 B.n355 B.n354 10.6151
R2151 B.n354 B.n158 10.6151
R2152 B.n348 B.n158 10.6151
R2153 B.n348 B.n347 10.6151
R2154 B.n347 B.n346 10.6151
R2155 B.n346 B.n160 10.6151
R2156 B.n340 B.n160 10.6151
R2157 B.n340 B.n339 10.6151
R2158 B.n339 B.n338 10.6151
R2159 B.n338 B.n162 10.6151
R2160 B.n332 B.n162 10.6151
R2161 B.n332 B.n331 10.6151
R2162 B.n331 B.n330 10.6151
R2163 B.n330 B.n164 10.6151
R2164 B.n324 B.n164 10.6151
R2165 B.n324 B.n323 10.6151
R2166 B.n323 B.n322 10.6151
R2167 B.n322 B.n166 10.6151
R2168 B.n316 B.n166 10.6151
R2169 B.n316 B.n315 10.6151
R2170 B.n313 B.n170 10.6151
R2171 B.n307 B.n170 10.6151
R2172 B.n307 B.n306 10.6151
R2173 B.n306 B.n305 10.6151
R2174 B.n305 B.n172 10.6151
R2175 B.n299 B.n172 10.6151
R2176 B.n299 B.n298 10.6151
R2177 B.n298 B.n297 10.6151
R2178 B.n293 B.n292 10.6151
R2179 B.n292 B.n178 10.6151
R2180 B.n287 B.n178 10.6151
R2181 B.n287 B.n286 10.6151
R2182 B.n286 B.n285 10.6151
R2183 B.n285 B.n180 10.6151
R2184 B.n279 B.n180 10.6151
R2185 B.n279 B.n278 10.6151
R2186 B.n278 B.n277 10.6151
R2187 B.n277 B.n182 10.6151
R2188 B.n271 B.n182 10.6151
R2189 B.n271 B.n270 10.6151
R2190 B.n270 B.n269 10.6151
R2191 B.n269 B.n184 10.6151
R2192 B.n263 B.n184 10.6151
R2193 B.n263 B.n262 10.6151
R2194 B.n262 B.n261 10.6151
R2195 B.n261 B.n186 10.6151
R2196 B.n255 B.n186 10.6151
R2197 B.n255 B.n254 10.6151
R2198 B.n254 B.n253 10.6151
R2199 B.n253 B.n188 10.6151
R2200 B.n247 B.n188 10.6151
R2201 B.n247 B.n246 10.6151
R2202 B.n246 B.n245 10.6151
R2203 B.n245 B.n190 10.6151
R2204 B.n239 B.n190 10.6151
R2205 B.n239 B.n238 10.6151
R2206 B.n238 B.n237 10.6151
R2207 B.n237 B.n192 10.6151
R2208 B.n231 B.n192 10.6151
R2209 B.n231 B.n230 10.6151
R2210 B.n230 B.n229 10.6151
R2211 B.n229 B.n194 10.6151
R2212 B.n223 B.n194 10.6151
R2213 B.n223 B.n222 10.6151
R2214 B.n222 B.n221 10.6151
R2215 B.n221 B.n196 10.6151
R2216 B.n215 B.n196 10.6151
R2217 B.n215 B.n214 10.6151
R2218 B.n214 B.n213 10.6151
R2219 B.n213 B.n198 10.6151
R2220 B.n207 B.n198 10.6151
R2221 B.n207 B.n206 10.6151
R2222 B.n206 B.n205 10.6151
R2223 B.n205 B.n200 10.6151
R2224 B.n200 B.n140 10.6151
R2225 B.n409 B.n136 10.6151
R2226 B.n419 B.n136 10.6151
R2227 B.n420 B.n419 10.6151
R2228 B.n421 B.n420 10.6151
R2229 B.n421 B.n128 10.6151
R2230 B.n431 B.n128 10.6151
R2231 B.n432 B.n431 10.6151
R2232 B.n433 B.n432 10.6151
R2233 B.n433 B.n120 10.6151
R2234 B.n443 B.n120 10.6151
R2235 B.n444 B.n443 10.6151
R2236 B.n445 B.n444 10.6151
R2237 B.n445 B.n112 10.6151
R2238 B.n455 B.n112 10.6151
R2239 B.n456 B.n455 10.6151
R2240 B.n457 B.n456 10.6151
R2241 B.n457 B.n104 10.6151
R2242 B.n469 B.n104 10.6151
R2243 B.n470 B.n469 10.6151
R2244 B.n471 B.n470 10.6151
R2245 B.n471 B.n0 10.6151
R2246 B.n756 B.n1 10.6151
R2247 B.n756 B.n755 10.6151
R2248 B.n755 B.n754 10.6151
R2249 B.n754 B.n9 10.6151
R2250 B.n748 B.n9 10.6151
R2251 B.n748 B.n747 10.6151
R2252 B.n747 B.n746 10.6151
R2253 B.n746 B.n17 10.6151
R2254 B.n740 B.n17 10.6151
R2255 B.n740 B.n739 10.6151
R2256 B.n739 B.n738 10.6151
R2257 B.n738 B.n24 10.6151
R2258 B.n732 B.n24 10.6151
R2259 B.n732 B.n731 10.6151
R2260 B.n731 B.n730 10.6151
R2261 B.n730 B.n31 10.6151
R2262 B.n724 B.n31 10.6151
R2263 B.n724 B.n723 10.6151
R2264 B.n723 B.n722 10.6151
R2265 B.n722 B.n38 10.6151
R2266 B.n716 B.n38 10.6151
R2267 B.t9 B.n130 9.63719
R2268 B.n459 B.t2 9.63719
R2269 B.t5 B.n750 9.63719
R2270 B.n727 B.t13 9.63719
R2271 B.n619 B.n618 6.5566
R2272 B.n602 B.n601 6.5566
R2273 B.n314 B.n313 6.5566
R2274 B.n297 B.n176 6.5566
R2275 B.n620 B.n619 4.05904
R2276 B.n601 B.n600 4.05904
R2277 B.n315 B.n314 4.05904
R2278 B.n293 B.n176 4.05904
R2279 B.n762 B.n0 2.81026
R2280 B.n762 B.n1 2.81026
R2281 B.n466 B.t6 0.567364
R2282 B.n11 B.t7 0.567364
R2283 VN.n1 VN.t1 649.865
R2284 VN.n7 VN.t4 649.865
R2285 VN.n2 VN.t7 623.044
R2286 VN.n3 VN.t5 623.044
R2287 VN.n4 VN.t2 623.044
R2288 VN.n8 VN.t6 623.044
R2289 VN.n9 VN.t0 623.044
R2290 VN.n10 VN.t3 623.044
R2291 VN.n5 VN.n4 161.3
R2292 VN.n11 VN.n10 161.3
R2293 VN.n9 VN.n6 80.6037
R2294 VN.n3 VN.n0 80.6037
R2295 VN.n3 VN.n2 48.2005
R2296 VN.n4 VN.n3 48.2005
R2297 VN.n9 VN.n8 48.2005
R2298 VN.n10 VN.n9 48.2005
R2299 VN.n7 VN.n6 45.2318
R2300 VN.n1 VN.n0 45.2318
R2301 VN VN.n11 43.6312
R2302 VN.n8 VN.n7 13.3799
R2303 VN.n2 VN.n1 13.3799
R2304 VN.n11 VN.n6 0.285035
R2305 VN.n5 VN.n0 0.285035
R2306 VN VN.n5 0.0516364
R2307 VDD2.n2 VDD2.n1 65.4368
R2308 VDD2.n2 VDD2.n0 65.4368
R2309 VDD2 VDD2.n5 65.4339
R2310 VDD2.n4 VDD2.n3 65.0871
R2311 VDD2.n4 VDD2.n2 39.5429
R2312 VDD2.n5 VDD2.t1 1.40177
R2313 VDD2.n5 VDD2.t3 1.40177
R2314 VDD2.n3 VDD2.t4 1.40177
R2315 VDD2.n3 VDD2.t7 1.40177
R2316 VDD2.n1 VDD2.t2 1.40177
R2317 VDD2.n1 VDD2.t5 1.40177
R2318 VDD2.n0 VDD2.t6 1.40177
R2319 VDD2.n0 VDD2.t0 1.40177
R2320 VDD2 VDD2.n4 0.463862
C0 VDD1 VDD2 0.78214f
C1 VP VDD2 0.307954f
C2 VN VDD2 5.95873f
C3 VP VDD1 6.11812f
C4 VTAIL VDD2 13.5625f
C5 VN VDD1 0.14817f
C6 VTAIL VDD1 13.5214f
C7 VP VN 5.62204f
C8 VP VTAIL 5.61093f
C9 VN VTAIL 5.59683f
C10 VDD2 B 3.572076f
C11 VDD1 B 3.794936f
C12 VTAIL B 10.028173f
C13 VN B 8.54405f
C14 VP B 6.419137f
C15 VDD2.t6 B 0.315511f
C16 VDD2.t0 B 0.315511f
C17 VDD2.n0 B 2.85028f
C18 VDD2.t2 B 0.315511f
C19 VDD2.t5 B 0.315511f
C20 VDD2.n1 B 2.85028f
C21 VDD2.n2 B 2.52972f
C22 VDD2.t4 B 0.315511f
C23 VDD2.t7 B 0.315511f
C24 VDD2.n3 B 2.84845f
C25 VDD2.n4 B 2.73263f
C26 VDD2.t1 B 0.315511f
C27 VDD2.t3 B 0.315511f
C28 VDD2.n5 B 2.85025f
C29 VN.n0 B 0.225856f
C30 VN.t1 B 1.14832f
C31 VN.n1 B 0.425099f
C32 VN.t7 B 1.13008f
C33 VN.n2 B 0.452411f
C34 VN.t5 B 1.13008f
C35 VN.n3 B 0.452411f
C36 VN.t2 B 1.13008f
C37 VN.n4 B 0.441953f
C38 VN.n5 B 0.051127f
C39 VN.n6 B 0.225856f
C40 VN.t6 B 1.13008f
C41 VN.t4 B 1.14832f
C42 VN.n7 B 0.425099f
C43 VN.n8 B 0.452411f
C44 VN.t0 B 1.13008f
C45 VN.n9 B 0.452411f
C46 VN.t3 B 1.13008f
C47 VN.n10 B 0.441953f
C48 VN.n11 B 2.04236f
C49 VDD1.t6 B 0.31384f
C50 VDD1.t4 B 0.31384f
C51 VDD1.n0 B 2.83584f
C52 VDD1.t3 B 0.31384f
C53 VDD1.t1 B 0.31384f
C54 VDD1.n1 B 2.83518f
C55 VDD1.t0 B 0.31384f
C56 VDD1.t5 B 0.31384f
C57 VDD1.n2 B 2.83518f
C58 VDD1.n3 B 2.57625f
C59 VDD1.t2 B 0.31384f
C60 VDD1.t7 B 0.31384f
C61 VDD1.n4 B 2.83335f
C62 VDD1.n5 B 2.75151f
C63 VTAIL.t11 B 0.226066f
C64 VTAIL.t0 B 0.226066f
C65 VTAIL.n0 B 1.98656f
C66 VTAIL.n1 B 0.245148f
C67 VTAIL.n2 B 0.028048f
C68 VTAIL.n3 B 0.020246f
C69 VTAIL.n4 B 0.011199f
C70 VTAIL.n5 B 0.025715f
C71 VTAIL.n6 B 0.011519f
C72 VTAIL.n7 B 0.020246f
C73 VTAIL.n8 B 0.010879f
C74 VTAIL.n9 B 0.025715f
C75 VTAIL.n10 B 0.011519f
C76 VTAIL.n11 B 0.020246f
C77 VTAIL.n12 B 0.010879f
C78 VTAIL.n13 B 0.025715f
C79 VTAIL.n14 B 0.011519f
C80 VTAIL.n15 B 0.020246f
C81 VTAIL.n16 B 0.010879f
C82 VTAIL.n17 B 0.025715f
C83 VTAIL.n18 B 0.011519f
C84 VTAIL.n19 B 0.020246f
C85 VTAIL.n20 B 0.010879f
C86 VTAIL.n21 B 0.025715f
C87 VTAIL.n22 B 0.011519f
C88 VTAIL.n23 B 0.020246f
C89 VTAIL.n24 B 0.010879f
C90 VTAIL.n25 B 0.019286f
C91 VTAIL.n26 B 0.01519f
C92 VTAIL.t10 B 0.04234f
C93 VTAIL.n27 B 0.127632f
C94 VTAIL.n28 B 1.23651f
C95 VTAIL.n29 B 0.010879f
C96 VTAIL.n30 B 0.011519f
C97 VTAIL.n31 B 0.025715f
C98 VTAIL.n32 B 0.025715f
C99 VTAIL.n33 B 0.011519f
C100 VTAIL.n34 B 0.010879f
C101 VTAIL.n35 B 0.020246f
C102 VTAIL.n36 B 0.020246f
C103 VTAIL.n37 B 0.010879f
C104 VTAIL.n38 B 0.011519f
C105 VTAIL.n39 B 0.025715f
C106 VTAIL.n40 B 0.025715f
C107 VTAIL.n41 B 0.011519f
C108 VTAIL.n42 B 0.010879f
C109 VTAIL.n43 B 0.020246f
C110 VTAIL.n44 B 0.020246f
C111 VTAIL.n45 B 0.010879f
C112 VTAIL.n46 B 0.011519f
C113 VTAIL.n47 B 0.025715f
C114 VTAIL.n48 B 0.025715f
C115 VTAIL.n49 B 0.011519f
C116 VTAIL.n50 B 0.010879f
C117 VTAIL.n51 B 0.020246f
C118 VTAIL.n52 B 0.020246f
C119 VTAIL.n53 B 0.010879f
C120 VTAIL.n54 B 0.011519f
C121 VTAIL.n55 B 0.025715f
C122 VTAIL.n56 B 0.025715f
C123 VTAIL.n57 B 0.011519f
C124 VTAIL.n58 B 0.010879f
C125 VTAIL.n59 B 0.020246f
C126 VTAIL.n60 B 0.020246f
C127 VTAIL.n61 B 0.010879f
C128 VTAIL.n62 B 0.011519f
C129 VTAIL.n63 B 0.025715f
C130 VTAIL.n64 B 0.025715f
C131 VTAIL.n65 B 0.011519f
C132 VTAIL.n66 B 0.010879f
C133 VTAIL.n67 B 0.020246f
C134 VTAIL.n68 B 0.020246f
C135 VTAIL.n69 B 0.010879f
C136 VTAIL.n70 B 0.010879f
C137 VTAIL.n71 B 0.011519f
C138 VTAIL.n72 B 0.025715f
C139 VTAIL.n73 B 0.025715f
C140 VTAIL.n74 B 0.054943f
C141 VTAIL.n75 B 0.011199f
C142 VTAIL.n76 B 0.010879f
C143 VTAIL.n77 B 0.052606f
C144 VTAIL.n78 B 0.030838f
C145 VTAIL.n79 B 0.104094f
C146 VTAIL.n80 B 0.028048f
C147 VTAIL.n81 B 0.020246f
C148 VTAIL.n82 B 0.011199f
C149 VTAIL.n83 B 0.025715f
C150 VTAIL.n84 B 0.011519f
C151 VTAIL.n85 B 0.020246f
C152 VTAIL.n86 B 0.010879f
C153 VTAIL.n87 B 0.025715f
C154 VTAIL.n88 B 0.011519f
C155 VTAIL.n89 B 0.020246f
C156 VTAIL.n90 B 0.010879f
C157 VTAIL.n91 B 0.025715f
C158 VTAIL.n92 B 0.011519f
C159 VTAIL.n93 B 0.020246f
C160 VTAIL.n94 B 0.010879f
C161 VTAIL.n95 B 0.025715f
C162 VTAIL.n96 B 0.011519f
C163 VTAIL.n97 B 0.020246f
C164 VTAIL.n98 B 0.010879f
C165 VTAIL.n99 B 0.025715f
C166 VTAIL.n100 B 0.011519f
C167 VTAIL.n101 B 0.020246f
C168 VTAIL.n102 B 0.010879f
C169 VTAIL.n103 B 0.019286f
C170 VTAIL.n104 B 0.01519f
C171 VTAIL.t9 B 0.04234f
C172 VTAIL.n105 B 0.127632f
C173 VTAIL.n106 B 1.23651f
C174 VTAIL.n107 B 0.010879f
C175 VTAIL.n108 B 0.011519f
C176 VTAIL.n109 B 0.025715f
C177 VTAIL.n110 B 0.025715f
C178 VTAIL.n111 B 0.011519f
C179 VTAIL.n112 B 0.010879f
C180 VTAIL.n113 B 0.020246f
C181 VTAIL.n114 B 0.020246f
C182 VTAIL.n115 B 0.010879f
C183 VTAIL.n116 B 0.011519f
C184 VTAIL.n117 B 0.025715f
C185 VTAIL.n118 B 0.025715f
C186 VTAIL.n119 B 0.011519f
C187 VTAIL.n120 B 0.010879f
C188 VTAIL.n121 B 0.020246f
C189 VTAIL.n122 B 0.020246f
C190 VTAIL.n123 B 0.010879f
C191 VTAIL.n124 B 0.011519f
C192 VTAIL.n125 B 0.025715f
C193 VTAIL.n126 B 0.025715f
C194 VTAIL.n127 B 0.011519f
C195 VTAIL.n128 B 0.010879f
C196 VTAIL.n129 B 0.020246f
C197 VTAIL.n130 B 0.020246f
C198 VTAIL.n131 B 0.010879f
C199 VTAIL.n132 B 0.011519f
C200 VTAIL.n133 B 0.025715f
C201 VTAIL.n134 B 0.025715f
C202 VTAIL.n135 B 0.011519f
C203 VTAIL.n136 B 0.010879f
C204 VTAIL.n137 B 0.020246f
C205 VTAIL.n138 B 0.020246f
C206 VTAIL.n139 B 0.010879f
C207 VTAIL.n140 B 0.011519f
C208 VTAIL.n141 B 0.025715f
C209 VTAIL.n142 B 0.025715f
C210 VTAIL.n143 B 0.011519f
C211 VTAIL.n144 B 0.010879f
C212 VTAIL.n145 B 0.020246f
C213 VTAIL.n146 B 0.020246f
C214 VTAIL.n147 B 0.010879f
C215 VTAIL.n148 B 0.010879f
C216 VTAIL.n149 B 0.011519f
C217 VTAIL.n150 B 0.025715f
C218 VTAIL.n151 B 0.025715f
C219 VTAIL.n152 B 0.054943f
C220 VTAIL.n153 B 0.011199f
C221 VTAIL.n154 B 0.010879f
C222 VTAIL.n155 B 0.052606f
C223 VTAIL.n156 B 0.030838f
C224 VTAIL.n157 B 0.104094f
C225 VTAIL.t4 B 0.226066f
C226 VTAIL.t6 B 0.226066f
C227 VTAIL.n158 B 1.98656f
C228 VTAIL.n159 B 0.294217f
C229 VTAIL.n160 B 0.028048f
C230 VTAIL.n161 B 0.020246f
C231 VTAIL.n162 B 0.011199f
C232 VTAIL.n163 B 0.025715f
C233 VTAIL.n164 B 0.011519f
C234 VTAIL.n165 B 0.020246f
C235 VTAIL.n166 B 0.010879f
C236 VTAIL.n167 B 0.025715f
C237 VTAIL.n168 B 0.011519f
C238 VTAIL.n169 B 0.020246f
C239 VTAIL.n170 B 0.010879f
C240 VTAIL.n171 B 0.025715f
C241 VTAIL.n172 B 0.011519f
C242 VTAIL.n173 B 0.020246f
C243 VTAIL.n174 B 0.010879f
C244 VTAIL.n175 B 0.025715f
C245 VTAIL.n176 B 0.011519f
C246 VTAIL.n177 B 0.020246f
C247 VTAIL.n178 B 0.010879f
C248 VTAIL.n179 B 0.025715f
C249 VTAIL.n180 B 0.011519f
C250 VTAIL.n181 B 0.020246f
C251 VTAIL.n182 B 0.010879f
C252 VTAIL.n183 B 0.019286f
C253 VTAIL.n184 B 0.01519f
C254 VTAIL.t2 B 0.04234f
C255 VTAIL.n185 B 0.127632f
C256 VTAIL.n186 B 1.23651f
C257 VTAIL.n187 B 0.010879f
C258 VTAIL.n188 B 0.011519f
C259 VTAIL.n189 B 0.025715f
C260 VTAIL.n190 B 0.025715f
C261 VTAIL.n191 B 0.011519f
C262 VTAIL.n192 B 0.010879f
C263 VTAIL.n193 B 0.020246f
C264 VTAIL.n194 B 0.020246f
C265 VTAIL.n195 B 0.010879f
C266 VTAIL.n196 B 0.011519f
C267 VTAIL.n197 B 0.025715f
C268 VTAIL.n198 B 0.025715f
C269 VTAIL.n199 B 0.011519f
C270 VTAIL.n200 B 0.010879f
C271 VTAIL.n201 B 0.020246f
C272 VTAIL.n202 B 0.020246f
C273 VTAIL.n203 B 0.010879f
C274 VTAIL.n204 B 0.011519f
C275 VTAIL.n205 B 0.025715f
C276 VTAIL.n206 B 0.025715f
C277 VTAIL.n207 B 0.011519f
C278 VTAIL.n208 B 0.010879f
C279 VTAIL.n209 B 0.020246f
C280 VTAIL.n210 B 0.020246f
C281 VTAIL.n211 B 0.010879f
C282 VTAIL.n212 B 0.011519f
C283 VTAIL.n213 B 0.025715f
C284 VTAIL.n214 B 0.025715f
C285 VTAIL.n215 B 0.011519f
C286 VTAIL.n216 B 0.010879f
C287 VTAIL.n217 B 0.020246f
C288 VTAIL.n218 B 0.020246f
C289 VTAIL.n219 B 0.010879f
C290 VTAIL.n220 B 0.011519f
C291 VTAIL.n221 B 0.025715f
C292 VTAIL.n222 B 0.025715f
C293 VTAIL.n223 B 0.011519f
C294 VTAIL.n224 B 0.010879f
C295 VTAIL.n225 B 0.020246f
C296 VTAIL.n226 B 0.020246f
C297 VTAIL.n227 B 0.010879f
C298 VTAIL.n228 B 0.010879f
C299 VTAIL.n229 B 0.011519f
C300 VTAIL.n230 B 0.025715f
C301 VTAIL.n231 B 0.025715f
C302 VTAIL.n232 B 0.054943f
C303 VTAIL.n233 B 0.011199f
C304 VTAIL.n234 B 0.010879f
C305 VTAIL.n235 B 0.052606f
C306 VTAIL.n236 B 0.030838f
C307 VTAIL.n237 B 1.19598f
C308 VTAIL.n238 B 0.028048f
C309 VTAIL.n239 B 0.020246f
C310 VTAIL.n240 B 0.011199f
C311 VTAIL.n241 B 0.025715f
C312 VTAIL.n242 B 0.010879f
C313 VTAIL.n243 B 0.011519f
C314 VTAIL.n244 B 0.020246f
C315 VTAIL.n245 B 0.010879f
C316 VTAIL.n246 B 0.025715f
C317 VTAIL.n247 B 0.011519f
C318 VTAIL.n248 B 0.020246f
C319 VTAIL.n249 B 0.010879f
C320 VTAIL.n250 B 0.025715f
C321 VTAIL.n251 B 0.011519f
C322 VTAIL.n252 B 0.020246f
C323 VTAIL.n253 B 0.010879f
C324 VTAIL.n254 B 0.025715f
C325 VTAIL.n255 B 0.011519f
C326 VTAIL.n256 B 0.020246f
C327 VTAIL.n257 B 0.010879f
C328 VTAIL.n258 B 0.025715f
C329 VTAIL.n259 B 0.011519f
C330 VTAIL.n260 B 0.020246f
C331 VTAIL.n261 B 0.010879f
C332 VTAIL.n262 B 0.019286f
C333 VTAIL.n263 B 0.01519f
C334 VTAIL.t14 B 0.04234f
C335 VTAIL.n264 B 0.127632f
C336 VTAIL.n265 B 1.23651f
C337 VTAIL.n266 B 0.010879f
C338 VTAIL.n267 B 0.011519f
C339 VTAIL.n268 B 0.025715f
C340 VTAIL.n269 B 0.025715f
C341 VTAIL.n270 B 0.011519f
C342 VTAIL.n271 B 0.010879f
C343 VTAIL.n272 B 0.020246f
C344 VTAIL.n273 B 0.020246f
C345 VTAIL.n274 B 0.010879f
C346 VTAIL.n275 B 0.011519f
C347 VTAIL.n276 B 0.025715f
C348 VTAIL.n277 B 0.025715f
C349 VTAIL.n278 B 0.011519f
C350 VTAIL.n279 B 0.010879f
C351 VTAIL.n280 B 0.020246f
C352 VTAIL.n281 B 0.020246f
C353 VTAIL.n282 B 0.010879f
C354 VTAIL.n283 B 0.011519f
C355 VTAIL.n284 B 0.025715f
C356 VTAIL.n285 B 0.025715f
C357 VTAIL.n286 B 0.011519f
C358 VTAIL.n287 B 0.010879f
C359 VTAIL.n288 B 0.020246f
C360 VTAIL.n289 B 0.020246f
C361 VTAIL.n290 B 0.010879f
C362 VTAIL.n291 B 0.011519f
C363 VTAIL.n292 B 0.025715f
C364 VTAIL.n293 B 0.025715f
C365 VTAIL.n294 B 0.011519f
C366 VTAIL.n295 B 0.010879f
C367 VTAIL.n296 B 0.020246f
C368 VTAIL.n297 B 0.020246f
C369 VTAIL.n298 B 0.010879f
C370 VTAIL.n299 B 0.011519f
C371 VTAIL.n300 B 0.025715f
C372 VTAIL.n301 B 0.025715f
C373 VTAIL.n302 B 0.011519f
C374 VTAIL.n303 B 0.010879f
C375 VTAIL.n304 B 0.020246f
C376 VTAIL.n305 B 0.020246f
C377 VTAIL.n306 B 0.010879f
C378 VTAIL.n307 B 0.011519f
C379 VTAIL.n308 B 0.025715f
C380 VTAIL.n309 B 0.025715f
C381 VTAIL.n310 B 0.054943f
C382 VTAIL.n311 B 0.011199f
C383 VTAIL.n312 B 0.010879f
C384 VTAIL.n313 B 0.052606f
C385 VTAIL.n314 B 0.030838f
C386 VTAIL.n315 B 1.19598f
C387 VTAIL.t15 B 0.226066f
C388 VTAIL.t12 B 0.226066f
C389 VTAIL.n316 B 1.98657f
C390 VTAIL.n317 B 0.294207f
C391 VTAIL.n318 B 0.028048f
C392 VTAIL.n319 B 0.020246f
C393 VTAIL.n320 B 0.011199f
C394 VTAIL.n321 B 0.025715f
C395 VTAIL.n322 B 0.010879f
C396 VTAIL.n323 B 0.011519f
C397 VTAIL.n324 B 0.020246f
C398 VTAIL.n325 B 0.010879f
C399 VTAIL.n326 B 0.025715f
C400 VTAIL.n327 B 0.011519f
C401 VTAIL.n328 B 0.020246f
C402 VTAIL.n329 B 0.010879f
C403 VTAIL.n330 B 0.025715f
C404 VTAIL.n331 B 0.011519f
C405 VTAIL.n332 B 0.020246f
C406 VTAIL.n333 B 0.010879f
C407 VTAIL.n334 B 0.025715f
C408 VTAIL.n335 B 0.011519f
C409 VTAIL.n336 B 0.020246f
C410 VTAIL.n337 B 0.010879f
C411 VTAIL.n338 B 0.025715f
C412 VTAIL.n339 B 0.011519f
C413 VTAIL.n340 B 0.020246f
C414 VTAIL.n341 B 0.010879f
C415 VTAIL.n342 B 0.019286f
C416 VTAIL.n343 B 0.01519f
C417 VTAIL.t13 B 0.04234f
C418 VTAIL.n344 B 0.127632f
C419 VTAIL.n345 B 1.23651f
C420 VTAIL.n346 B 0.010879f
C421 VTAIL.n347 B 0.011519f
C422 VTAIL.n348 B 0.025715f
C423 VTAIL.n349 B 0.025715f
C424 VTAIL.n350 B 0.011519f
C425 VTAIL.n351 B 0.010879f
C426 VTAIL.n352 B 0.020246f
C427 VTAIL.n353 B 0.020246f
C428 VTAIL.n354 B 0.010879f
C429 VTAIL.n355 B 0.011519f
C430 VTAIL.n356 B 0.025715f
C431 VTAIL.n357 B 0.025715f
C432 VTAIL.n358 B 0.011519f
C433 VTAIL.n359 B 0.010879f
C434 VTAIL.n360 B 0.020246f
C435 VTAIL.n361 B 0.020246f
C436 VTAIL.n362 B 0.010879f
C437 VTAIL.n363 B 0.011519f
C438 VTAIL.n364 B 0.025715f
C439 VTAIL.n365 B 0.025715f
C440 VTAIL.n366 B 0.011519f
C441 VTAIL.n367 B 0.010879f
C442 VTAIL.n368 B 0.020246f
C443 VTAIL.n369 B 0.020246f
C444 VTAIL.n370 B 0.010879f
C445 VTAIL.n371 B 0.011519f
C446 VTAIL.n372 B 0.025715f
C447 VTAIL.n373 B 0.025715f
C448 VTAIL.n374 B 0.011519f
C449 VTAIL.n375 B 0.010879f
C450 VTAIL.n376 B 0.020246f
C451 VTAIL.n377 B 0.020246f
C452 VTAIL.n378 B 0.010879f
C453 VTAIL.n379 B 0.011519f
C454 VTAIL.n380 B 0.025715f
C455 VTAIL.n381 B 0.025715f
C456 VTAIL.n382 B 0.011519f
C457 VTAIL.n383 B 0.010879f
C458 VTAIL.n384 B 0.020246f
C459 VTAIL.n385 B 0.020246f
C460 VTAIL.n386 B 0.010879f
C461 VTAIL.n387 B 0.011519f
C462 VTAIL.n388 B 0.025715f
C463 VTAIL.n389 B 0.025715f
C464 VTAIL.n390 B 0.054943f
C465 VTAIL.n391 B 0.011199f
C466 VTAIL.n392 B 0.010879f
C467 VTAIL.n393 B 0.052606f
C468 VTAIL.n394 B 0.030838f
C469 VTAIL.n395 B 0.104094f
C470 VTAIL.n396 B 0.028048f
C471 VTAIL.n397 B 0.020246f
C472 VTAIL.n398 B 0.011199f
C473 VTAIL.n399 B 0.025715f
C474 VTAIL.n400 B 0.010879f
C475 VTAIL.n401 B 0.011519f
C476 VTAIL.n402 B 0.020246f
C477 VTAIL.n403 B 0.010879f
C478 VTAIL.n404 B 0.025715f
C479 VTAIL.n405 B 0.011519f
C480 VTAIL.n406 B 0.020246f
C481 VTAIL.n407 B 0.010879f
C482 VTAIL.n408 B 0.025715f
C483 VTAIL.n409 B 0.011519f
C484 VTAIL.n410 B 0.020246f
C485 VTAIL.n411 B 0.010879f
C486 VTAIL.n412 B 0.025715f
C487 VTAIL.n413 B 0.011519f
C488 VTAIL.n414 B 0.020246f
C489 VTAIL.n415 B 0.010879f
C490 VTAIL.n416 B 0.025715f
C491 VTAIL.n417 B 0.011519f
C492 VTAIL.n418 B 0.020246f
C493 VTAIL.n419 B 0.010879f
C494 VTAIL.n420 B 0.019286f
C495 VTAIL.n421 B 0.01519f
C496 VTAIL.t3 B 0.04234f
C497 VTAIL.n422 B 0.127632f
C498 VTAIL.n423 B 1.23651f
C499 VTAIL.n424 B 0.010879f
C500 VTAIL.n425 B 0.011519f
C501 VTAIL.n426 B 0.025715f
C502 VTAIL.n427 B 0.025715f
C503 VTAIL.n428 B 0.011519f
C504 VTAIL.n429 B 0.010879f
C505 VTAIL.n430 B 0.020246f
C506 VTAIL.n431 B 0.020246f
C507 VTAIL.n432 B 0.010879f
C508 VTAIL.n433 B 0.011519f
C509 VTAIL.n434 B 0.025715f
C510 VTAIL.n435 B 0.025715f
C511 VTAIL.n436 B 0.011519f
C512 VTAIL.n437 B 0.010879f
C513 VTAIL.n438 B 0.020246f
C514 VTAIL.n439 B 0.020246f
C515 VTAIL.n440 B 0.010879f
C516 VTAIL.n441 B 0.011519f
C517 VTAIL.n442 B 0.025715f
C518 VTAIL.n443 B 0.025715f
C519 VTAIL.n444 B 0.011519f
C520 VTAIL.n445 B 0.010879f
C521 VTAIL.n446 B 0.020246f
C522 VTAIL.n447 B 0.020246f
C523 VTAIL.n448 B 0.010879f
C524 VTAIL.n449 B 0.011519f
C525 VTAIL.n450 B 0.025715f
C526 VTAIL.n451 B 0.025715f
C527 VTAIL.n452 B 0.011519f
C528 VTAIL.n453 B 0.010879f
C529 VTAIL.n454 B 0.020246f
C530 VTAIL.n455 B 0.020246f
C531 VTAIL.n456 B 0.010879f
C532 VTAIL.n457 B 0.011519f
C533 VTAIL.n458 B 0.025715f
C534 VTAIL.n459 B 0.025715f
C535 VTAIL.n460 B 0.011519f
C536 VTAIL.n461 B 0.010879f
C537 VTAIL.n462 B 0.020246f
C538 VTAIL.n463 B 0.020246f
C539 VTAIL.n464 B 0.010879f
C540 VTAIL.n465 B 0.011519f
C541 VTAIL.n466 B 0.025715f
C542 VTAIL.n467 B 0.025715f
C543 VTAIL.n468 B 0.054943f
C544 VTAIL.n469 B 0.011199f
C545 VTAIL.n470 B 0.010879f
C546 VTAIL.n471 B 0.052606f
C547 VTAIL.n472 B 0.030838f
C548 VTAIL.n473 B 0.104094f
C549 VTAIL.t7 B 0.226066f
C550 VTAIL.t8 B 0.226066f
C551 VTAIL.n474 B 1.98657f
C552 VTAIL.n475 B 0.294207f
C553 VTAIL.n476 B 0.028048f
C554 VTAIL.n477 B 0.020246f
C555 VTAIL.n478 B 0.011199f
C556 VTAIL.n479 B 0.025715f
C557 VTAIL.n480 B 0.010879f
C558 VTAIL.n481 B 0.011519f
C559 VTAIL.n482 B 0.020246f
C560 VTAIL.n483 B 0.010879f
C561 VTAIL.n484 B 0.025715f
C562 VTAIL.n485 B 0.011519f
C563 VTAIL.n486 B 0.020246f
C564 VTAIL.n487 B 0.010879f
C565 VTAIL.n488 B 0.025715f
C566 VTAIL.n489 B 0.011519f
C567 VTAIL.n490 B 0.020246f
C568 VTAIL.n491 B 0.010879f
C569 VTAIL.n492 B 0.025715f
C570 VTAIL.n493 B 0.011519f
C571 VTAIL.n494 B 0.020246f
C572 VTAIL.n495 B 0.010879f
C573 VTAIL.n496 B 0.025715f
C574 VTAIL.n497 B 0.011519f
C575 VTAIL.n498 B 0.020246f
C576 VTAIL.n499 B 0.010879f
C577 VTAIL.n500 B 0.019286f
C578 VTAIL.n501 B 0.01519f
C579 VTAIL.t5 B 0.04234f
C580 VTAIL.n502 B 0.127632f
C581 VTAIL.n503 B 1.23651f
C582 VTAIL.n504 B 0.010879f
C583 VTAIL.n505 B 0.011519f
C584 VTAIL.n506 B 0.025715f
C585 VTAIL.n507 B 0.025715f
C586 VTAIL.n508 B 0.011519f
C587 VTAIL.n509 B 0.010879f
C588 VTAIL.n510 B 0.020246f
C589 VTAIL.n511 B 0.020246f
C590 VTAIL.n512 B 0.010879f
C591 VTAIL.n513 B 0.011519f
C592 VTAIL.n514 B 0.025715f
C593 VTAIL.n515 B 0.025715f
C594 VTAIL.n516 B 0.011519f
C595 VTAIL.n517 B 0.010879f
C596 VTAIL.n518 B 0.020246f
C597 VTAIL.n519 B 0.020246f
C598 VTAIL.n520 B 0.010879f
C599 VTAIL.n521 B 0.011519f
C600 VTAIL.n522 B 0.025715f
C601 VTAIL.n523 B 0.025715f
C602 VTAIL.n524 B 0.011519f
C603 VTAIL.n525 B 0.010879f
C604 VTAIL.n526 B 0.020246f
C605 VTAIL.n527 B 0.020246f
C606 VTAIL.n528 B 0.010879f
C607 VTAIL.n529 B 0.011519f
C608 VTAIL.n530 B 0.025715f
C609 VTAIL.n531 B 0.025715f
C610 VTAIL.n532 B 0.011519f
C611 VTAIL.n533 B 0.010879f
C612 VTAIL.n534 B 0.020246f
C613 VTAIL.n535 B 0.020246f
C614 VTAIL.n536 B 0.010879f
C615 VTAIL.n537 B 0.011519f
C616 VTAIL.n538 B 0.025715f
C617 VTAIL.n539 B 0.025715f
C618 VTAIL.n540 B 0.011519f
C619 VTAIL.n541 B 0.010879f
C620 VTAIL.n542 B 0.020246f
C621 VTAIL.n543 B 0.020246f
C622 VTAIL.n544 B 0.010879f
C623 VTAIL.n545 B 0.011519f
C624 VTAIL.n546 B 0.025715f
C625 VTAIL.n547 B 0.025715f
C626 VTAIL.n548 B 0.054943f
C627 VTAIL.n549 B 0.011199f
C628 VTAIL.n550 B 0.010879f
C629 VTAIL.n551 B 0.052606f
C630 VTAIL.n552 B 0.030838f
C631 VTAIL.n553 B 1.19598f
C632 VTAIL.n554 B 0.028048f
C633 VTAIL.n555 B 0.020246f
C634 VTAIL.n556 B 0.011199f
C635 VTAIL.n557 B 0.025715f
C636 VTAIL.n558 B 0.011519f
C637 VTAIL.n559 B 0.020246f
C638 VTAIL.n560 B 0.010879f
C639 VTAIL.n561 B 0.025715f
C640 VTAIL.n562 B 0.011519f
C641 VTAIL.n563 B 0.020246f
C642 VTAIL.n564 B 0.010879f
C643 VTAIL.n565 B 0.025715f
C644 VTAIL.n566 B 0.011519f
C645 VTAIL.n567 B 0.020246f
C646 VTAIL.n568 B 0.010879f
C647 VTAIL.n569 B 0.025715f
C648 VTAIL.n570 B 0.011519f
C649 VTAIL.n571 B 0.020246f
C650 VTAIL.n572 B 0.010879f
C651 VTAIL.n573 B 0.025715f
C652 VTAIL.n574 B 0.011519f
C653 VTAIL.n575 B 0.020246f
C654 VTAIL.n576 B 0.010879f
C655 VTAIL.n577 B 0.019286f
C656 VTAIL.n578 B 0.01519f
C657 VTAIL.t1 B 0.04234f
C658 VTAIL.n579 B 0.127632f
C659 VTAIL.n580 B 1.23651f
C660 VTAIL.n581 B 0.010879f
C661 VTAIL.n582 B 0.011519f
C662 VTAIL.n583 B 0.025715f
C663 VTAIL.n584 B 0.025715f
C664 VTAIL.n585 B 0.011519f
C665 VTAIL.n586 B 0.010879f
C666 VTAIL.n587 B 0.020246f
C667 VTAIL.n588 B 0.020246f
C668 VTAIL.n589 B 0.010879f
C669 VTAIL.n590 B 0.011519f
C670 VTAIL.n591 B 0.025715f
C671 VTAIL.n592 B 0.025715f
C672 VTAIL.n593 B 0.011519f
C673 VTAIL.n594 B 0.010879f
C674 VTAIL.n595 B 0.020246f
C675 VTAIL.n596 B 0.020246f
C676 VTAIL.n597 B 0.010879f
C677 VTAIL.n598 B 0.011519f
C678 VTAIL.n599 B 0.025715f
C679 VTAIL.n600 B 0.025715f
C680 VTAIL.n601 B 0.011519f
C681 VTAIL.n602 B 0.010879f
C682 VTAIL.n603 B 0.020246f
C683 VTAIL.n604 B 0.020246f
C684 VTAIL.n605 B 0.010879f
C685 VTAIL.n606 B 0.011519f
C686 VTAIL.n607 B 0.025715f
C687 VTAIL.n608 B 0.025715f
C688 VTAIL.n609 B 0.011519f
C689 VTAIL.n610 B 0.010879f
C690 VTAIL.n611 B 0.020246f
C691 VTAIL.n612 B 0.020246f
C692 VTAIL.n613 B 0.010879f
C693 VTAIL.n614 B 0.011519f
C694 VTAIL.n615 B 0.025715f
C695 VTAIL.n616 B 0.025715f
C696 VTAIL.n617 B 0.011519f
C697 VTAIL.n618 B 0.010879f
C698 VTAIL.n619 B 0.020246f
C699 VTAIL.n620 B 0.020246f
C700 VTAIL.n621 B 0.010879f
C701 VTAIL.n622 B 0.010879f
C702 VTAIL.n623 B 0.011519f
C703 VTAIL.n624 B 0.025715f
C704 VTAIL.n625 B 0.025715f
C705 VTAIL.n626 B 0.054943f
C706 VTAIL.n627 B 0.011199f
C707 VTAIL.n628 B 0.010879f
C708 VTAIL.n629 B 0.052606f
C709 VTAIL.n630 B 0.030838f
C710 VTAIL.n631 B 1.19218f
C711 VP.n0 B 0.077504f
C712 VP.t4 B 1.14095f
C713 VP.n1 B 0.446203f
C714 VP.n2 B 0.228028f
C715 VP.t0 B 1.14095f
C716 VP.t5 B 1.14095f
C717 VP.t3 B 1.14095f
C718 VP.t1 B 1.15937f
C719 VP.n3 B 0.429187f
C720 VP.n4 B 0.456762f
C721 VP.n5 B 0.456762f
C722 VP.n6 B 0.446203f
C723 VP.n7 B 2.03151f
C724 VP.n8 B 2.07019f
C725 VP.n9 B 0.077504f
C726 VP.t6 B 1.14095f
C727 VP.n10 B 0.456762f
C728 VP.t7 B 1.14095f
C729 VP.n11 B 0.456762f
C730 VP.t2 B 1.14095f
C731 VP.n12 B 0.446203f
C732 VP.n13 B 0.051619f
.ends

