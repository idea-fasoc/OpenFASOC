* NGSPICE file created from diff_pair_sample_1597.ext - technology: sky130A

.subckt diff_pair_sample_1597 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=5.4717 pd=28.84 as=5.4717 ps=28.84 w=14.03 l=0.83
X1 VDD1.t1 VP.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=5.4717 pd=28.84 as=5.4717 ps=28.84 w=14.03 l=0.83
X2 VDD1.t0 VP.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=5.4717 pd=28.84 as=5.4717 ps=28.84 w=14.03 l=0.83
X3 VDD2.t0 VN.t1 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=5.4717 pd=28.84 as=5.4717 ps=28.84 w=14.03 l=0.83
X4 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=5.4717 pd=28.84 as=0 ps=0 w=14.03 l=0.83
X5 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=5.4717 pd=28.84 as=0 ps=0 w=14.03 l=0.83
X6 B.t8 B.t6 B.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=5.4717 pd=28.84 as=0 ps=0 w=14.03 l=0.83
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=5.4717 pd=28.84 as=0 ps=0 w=14.03 l=0.83
R0 VN VN.t0 658.192
R1 VN VN.t1 616.347
R2 VTAIL.n306 VTAIL.n234 289.615
R3 VTAIL.n72 VTAIL.n0 289.615
R4 VTAIL.n228 VTAIL.n156 289.615
R5 VTAIL.n150 VTAIL.n78 289.615
R6 VTAIL.n258 VTAIL.n257 185
R7 VTAIL.n263 VTAIL.n262 185
R8 VTAIL.n265 VTAIL.n264 185
R9 VTAIL.n254 VTAIL.n253 185
R10 VTAIL.n271 VTAIL.n270 185
R11 VTAIL.n273 VTAIL.n272 185
R12 VTAIL.n250 VTAIL.n249 185
R13 VTAIL.n279 VTAIL.n278 185
R14 VTAIL.n281 VTAIL.n280 185
R15 VTAIL.n246 VTAIL.n245 185
R16 VTAIL.n287 VTAIL.n286 185
R17 VTAIL.n289 VTAIL.n288 185
R18 VTAIL.n242 VTAIL.n241 185
R19 VTAIL.n295 VTAIL.n294 185
R20 VTAIL.n297 VTAIL.n296 185
R21 VTAIL.n238 VTAIL.n237 185
R22 VTAIL.n304 VTAIL.n303 185
R23 VTAIL.n305 VTAIL.n236 185
R24 VTAIL.n307 VTAIL.n306 185
R25 VTAIL.n24 VTAIL.n23 185
R26 VTAIL.n29 VTAIL.n28 185
R27 VTAIL.n31 VTAIL.n30 185
R28 VTAIL.n20 VTAIL.n19 185
R29 VTAIL.n37 VTAIL.n36 185
R30 VTAIL.n39 VTAIL.n38 185
R31 VTAIL.n16 VTAIL.n15 185
R32 VTAIL.n45 VTAIL.n44 185
R33 VTAIL.n47 VTAIL.n46 185
R34 VTAIL.n12 VTAIL.n11 185
R35 VTAIL.n53 VTAIL.n52 185
R36 VTAIL.n55 VTAIL.n54 185
R37 VTAIL.n8 VTAIL.n7 185
R38 VTAIL.n61 VTAIL.n60 185
R39 VTAIL.n63 VTAIL.n62 185
R40 VTAIL.n4 VTAIL.n3 185
R41 VTAIL.n70 VTAIL.n69 185
R42 VTAIL.n71 VTAIL.n2 185
R43 VTAIL.n73 VTAIL.n72 185
R44 VTAIL.n229 VTAIL.n228 185
R45 VTAIL.n227 VTAIL.n158 185
R46 VTAIL.n226 VTAIL.n225 185
R47 VTAIL.n161 VTAIL.n159 185
R48 VTAIL.n220 VTAIL.n219 185
R49 VTAIL.n218 VTAIL.n217 185
R50 VTAIL.n165 VTAIL.n164 185
R51 VTAIL.n212 VTAIL.n211 185
R52 VTAIL.n210 VTAIL.n209 185
R53 VTAIL.n169 VTAIL.n168 185
R54 VTAIL.n204 VTAIL.n203 185
R55 VTAIL.n202 VTAIL.n201 185
R56 VTAIL.n173 VTAIL.n172 185
R57 VTAIL.n196 VTAIL.n195 185
R58 VTAIL.n194 VTAIL.n193 185
R59 VTAIL.n177 VTAIL.n176 185
R60 VTAIL.n188 VTAIL.n187 185
R61 VTAIL.n186 VTAIL.n185 185
R62 VTAIL.n181 VTAIL.n180 185
R63 VTAIL.n151 VTAIL.n150 185
R64 VTAIL.n149 VTAIL.n80 185
R65 VTAIL.n148 VTAIL.n147 185
R66 VTAIL.n83 VTAIL.n81 185
R67 VTAIL.n142 VTAIL.n141 185
R68 VTAIL.n140 VTAIL.n139 185
R69 VTAIL.n87 VTAIL.n86 185
R70 VTAIL.n134 VTAIL.n133 185
R71 VTAIL.n132 VTAIL.n131 185
R72 VTAIL.n91 VTAIL.n90 185
R73 VTAIL.n126 VTAIL.n125 185
R74 VTAIL.n124 VTAIL.n123 185
R75 VTAIL.n95 VTAIL.n94 185
R76 VTAIL.n118 VTAIL.n117 185
R77 VTAIL.n116 VTAIL.n115 185
R78 VTAIL.n99 VTAIL.n98 185
R79 VTAIL.n110 VTAIL.n109 185
R80 VTAIL.n108 VTAIL.n107 185
R81 VTAIL.n103 VTAIL.n102 185
R82 VTAIL.n259 VTAIL.t3 147.659
R83 VTAIL.n25 VTAIL.t1 147.659
R84 VTAIL.n182 VTAIL.t0 147.659
R85 VTAIL.n104 VTAIL.t2 147.659
R86 VTAIL.n263 VTAIL.n257 104.615
R87 VTAIL.n264 VTAIL.n263 104.615
R88 VTAIL.n264 VTAIL.n253 104.615
R89 VTAIL.n271 VTAIL.n253 104.615
R90 VTAIL.n272 VTAIL.n271 104.615
R91 VTAIL.n272 VTAIL.n249 104.615
R92 VTAIL.n279 VTAIL.n249 104.615
R93 VTAIL.n280 VTAIL.n279 104.615
R94 VTAIL.n280 VTAIL.n245 104.615
R95 VTAIL.n287 VTAIL.n245 104.615
R96 VTAIL.n288 VTAIL.n287 104.615
R97 VTAIL.n288 VTAIL.n241 104.615
R98 VTAIL.n295 VTAIL.n241 104.615
R99 VTAIL.n296 VTAIL.n295 104.615
R100 VTAIL.n296 VTAIL.n237 104.615
R101 VTAIL.n304 VTAIL.n237 104.615
R102 VTAIL.n305 VTAIL.n304 104.615
R103 VTAIL.n306 VTAIL.n305 104.615
R104 VTAIL.n29 VTAIL.n23 104.615
R105 VTAIL.n30 VTAIL.n29 104.615
R106 VTAIL.n30 VTAIL.n19 104.615
R107 VTAIL.n37 VTAIL.n19 104.615
R108 VTAIL.n38 VTAIL.n37 104.615
R109 VTAIL.n38 VTAIL.n15 104.615
R110 VTAIL.n45 VTAIL.n15 104.615
R111 VTAIL.n46 VTAIL.n45 104.615
R112 VTAIL.n46 VTAIL.n11 104.615
R113 VTAIL.n53 VTAIL.n11 104.615
R114 VTAIL.n54 VTAIL.n53 104.615
R115 VTAIL.n54 VTAIL.n7 104.615
R116 VTAIL.n61 VTAIL.n7 104.615
R117 VTAIL.n62 VTAIL.n61 104.615
R118 VTAIL.n62 VTAIL.n3 104.615
R119 VTAIL.n70 VTAIL.n3 104.615
R120 VTAIL.n71 VTAIL.n70 104.615
R121 VTAIL.n72 VTAIL.n71 104.615
R122 VTAIL.n228 VTAIL.n227 104.615
R123 VTAIL.n227 VTAIL.n226 104.615
R124 VTAIL.n226 VTAIL.n159 104.615
R125 VTAIL.n219 VTAIL.n159 104.615
R126 VTAIL.n219 VTAIL.n218 104.615
R127 VTAIL.n218 VTAIL.n164 104.615
R128 VTAIL.n211 VTAIL.n164 104.615
R129 VTAIL.n211 VTAIL.n210 104.615
R130 VTAIL.n210 VTAIL.n168 104.615
R131 VTAIL.n203 VTAIL.n168 104.615
R132 VTAIL.n203 VTAIL.n202 104.615
R133 VTAIL.n202 VTAIL.n172 104.615
R134 VTAIL.n195 VTAIL.n172 104.615
R135 VTAIL.n195 VTAIL.n194 104.615
R136 VTAIL.n194 VTAIL.n176 104.615
R137 VTAIL.n187 VTAIL.n176 104.615
R138 VTAIL.n187 VTAIL.n186 104.615
R139 VTAIL.n186 VTAIL.n180 104.615
R140 VTAIL.n150 VTAIL.n149 104.615
R141 VTAIL.n149 VTAIL.n148 104.615
R142 VTAIL.n148 VTAIL.n81 104.615
R143 VTAIL.n141 VTAIL.n81 104.615
R144 VTAIL.n141 VTAIL.n140 104.615
R145 VTAIL.n140 VTAIL.n86 104.615
R146 VTAIL.n133 VTAIL.n86 104.615
R147 VTAIL.n133 VTAIL.n132 104.615
R148 VTAIL.n132 VTAIL.n90 104.615
R149 VTAIL.n125 VTAIL.n90 104.615
R150 VTAIL.n125 VTAIL.n124 104.615
R151 VTAIL.n124 VTAIL.n94 104.615
R152 VTAIL.n117 VTAIL.n94 104.615
R153 VTAIL.n117 VTAIL.n116 104.615
R154 VTAIL.n116 VTAIL.n98 104.615
R155 VTAIL.n109 VTAIL.n98 104.615
R156 VTAIL.n109 VTAIL.n108 104.615
R157 VTAIL.n108 VTAIL.n102 104.615
R158 VTAIL.t3 VTAIL.n257 52.3082
R159 VTAIL.t1 VTAIL.n23 52.3082
R160 VTAIL.t0 VTAIL.n180 52.3082
R161 VTAIL.t2 VTAIL.n102 52.3082
R162 VTAIL.n311 VTAIL.n310 34.3187
R163 VTAIL.n77 VTAIL.n76 34.3187
R164 VTAIL.n233 VTAIL.n232 34.3187
R165 VTAIL.n155 VTAIL.n154 34.3187
R166 VTAIL.n155 VTAIL.n77 26.4789
R167 VTAIL.n311 VTAIL.n233 25.4789
R168 VTAIL.n259 VTAIL.n258 15.6677
R169 VTAIL.n25 VTAIL.n24 15.6677
R170 VTAIL.n182 VTAIL.n181 15.6677
R171 VTAIL.n104 VTAIL.n103 15.6677
R172 VTAIL.n307 VTAIL.n236 13.1884
R173 VTAIL.n73 VTAIL.n2 13.1884
R174 VTAIL.n229 VTAIL.n158 13.1884
R175 VTAIL.n151 VTAIL.n80 13.1884
R176 VTAIL.n262 VTAIL.n261 12.8005
R177 VTAIL.n303 VTAIL.n302 12.8005
R178 VTAIL.n308 VTAIL.n234 12.8005
R179 VTAIL.n28 VTAIL.n27 12.8005
R180 VTAIL.n69 VTAIL.n68 12.8005
R181 VTAIL.n74 VTAIL.n0 12.8005
R182 VTAIL.n230 VTAIL.n156 12.8005
R183 VTAIL.n225 VTAIL.n160 12.8005
R184 VTAIL.n185 VTAIL.n184 12.8005
R185 VTAIL.n152 VTAIL.n78 12.8005
R186 VTAIL.n147 VTAIL.n82 12.8005
R187 VTAIL.n107 VTAIL.n106 12.8005
R188 VTAIL.n265 VTAIL.n256 12.0247
R189 VTAIL.n301 VTAIL.n238 12.0247
R190 VTAIL.n31 VTAIL.n22 12.0247
R191 VTAIL.n67 VTAIL.n4 12.0247
R192 VTAIL.n224 VTAIL.n161 12.0247
R193 VTAIL.n188 VTAIL.n179 12.0247
R194 VTAIL.n146 VTAIL.n83 12.0247
R195 VTAIL.n110 VTAIL.n101 12.0247
R196 VTAIL.n266 VTAIL.n254 11.249
R197 VTAIL.n298 VTAIL.n297 11.249
R198 VTAIL.n32 VTAIL.n20 11.249
R199 VTAIL.n64 VTAIL.n63 11.249
R200 VTAIL.n221 VTAIL.n220 11.249
R201 VTAIL.n189 VTAIL.n177 11.249
R202 VTAIL.n143 VTAIL.n142 11.249
R203 VTAIL.n111 VTAIL.n99 11.249
R204 VTAIL.n270 VTAIL.n269 10.4732
R205 VTAIL.n294 VTAIL.n240 10.4732
R206 VTAIL.n36 VTAIL.n35 10.4732
R207 VTAIL.n60 VTAIL.n6 10.4732
R208 VTAIL.n217 VTAIL.n163 10.4732
R209 VTAIL.n193 VTAIL.n192 10.4732
R210 VTAIL.n139 VTAIL.n85 10.4732
R211 VTAIL.n115 VTAIL.n114 10.4732
R212 VTAIL.n273 VTAIL.n252 9.69747
R213 VTAIL.n293 VTAIL.n242 9.69747
R214 VTAIL.n39 VTAIL.n18 9.69747
R215 VTAIL.n59 VTAIL.n8 9.69747
R216 VTAIL.n216 VTAIL.n165 9.69747
R217 VTAIL.n196 VTAIL.n175 9.69747
R218 VTAIL.n138 VTAIL.n87 9.69747
R219 VTAIL.n118 VTAIL.n97 9.69747
R220 VTAIL.n310 VTAIL.n309 9.45567
R221 VTAIL.n76 VTAIL.n75 9.45567
R222 VTAIL.n232 VTAIL.n231 9.45567
R223 VTAIL.n154 VTAIL.n153 9.45567
R224 VTAIL.n309 VTAIL.n308 9.3005
R225 VTAIL.n248 VTAIL.n247 9.3005
R226 VTAIL.n277 VTAIL.n276 9.3005
R227 VTAIL.n275 VTAIL.n274 9.3005
R228 VTAIL.n252 VTAIL.n251 9.3005
R229 VTAIL.n269 VTAIL.n268 9.3005
R230 VTAIL.n267 VTAIL.n266 9.3005
R231 VTAIL.n256 VTAIL.n255 9.3005
R232 VTAIL.n261 VTAIL.n260 9.3005
R233 VTAIL.n283 VTAIL.n282 9.3005
R234 VTAIL.n285 VTAIL.n284 9.3005
R235 VTAIL.n244 VTAIL.n243 9.3005
R236 VTAIL.n291 VTAIL.n290 9.3005
R237 VTAIL.n293 VTAIL.n292 9.3005
R238 VTAIL.n240 VTAIL.n239 9.3005
R239 VTAIL.n299 VTAIL.n298 9.3005
R240 VTAIL.n301 VTAIL.n300 9.3005
R241 VTAIL.n302 VTAIL.n235 9.3005
R242 VTAIL.n75 VTAIL.n74 9.3005
R243 VTAIL.n14 VTAIL.n13 9.3005
R244 VTAIL.n43 VTAIL.n42 9.3005
R245 VTAIL.n41 VTAIL.n40 9.3005
R246 VTAIL.n18 VTAIL.n17 9.3005
R247 VTAIL.n35 VTAIL.n34 9.3005
R248 VTAIL.n33 VTAIL.n32 9.3005
R249 VTAIL.n22 VTAIL.n21 9.3005
R250 VTAIL.n27 VTAIL.n26 9.3005
R251 VTAIL.n49 VTAIL.n48 9.3005
R252 VTAIL.n51 VTAIL.n50 9.3005
R253 VTAIL.n10 VTAIL.n9 9.3005
R254 VTAIL.n57 VTAIL.n56 9.3005
R255 VTAIL.n59 VTAIL.n58 9.3005
R256 VTAIL.n6 VTAIL.n5 9.3005
R257 VTAIL.n65 VTAIL.n64 9.3005
R258 VTAIL.n67 VTAIL.n66 9.3005
R259 VTAIL.n68 VTAIL.n1 9.3005
R260 VTAIL.n208 VTAIL.n207 9.3005
R261 VTAIL.n167 VTAIL.n166 9.3005
R262 VTAIL.n214 VTAIL.n213 9.3005
R263 VTAIL.n216 VTAIL.n215 9.3005
R264 VTAIL.n163 VTAIL.n162 9.3005
R265 VTAIL.n222 VTAIL.n221 9.3005
R266 VTAIL.n224 VTAIL.n223 9.3005
R267 VTAIL.n160 VTAIL.n157 9.3005
R268 VTAIL.n231 VTAIL.n230 9.3005
R269 VTAIL.n206 VTAIL.n205 9.3005
R270 VTAIL.n171 VTAIL.n170 9.3005
R271 VTAIL.n200 VTAIL.n199 9.3005
R272 VTAIL.n198 VTAIL.n197 9.3005
R273 VTAIL.n175 VTAIL.n174 9.3005
R274 VTAIL.n192 VTAIL.n191 9.3005
R275 VTAIL.n190 VTAIL.n189 9.3005
R276 VTAIL.n179 VTAIL.n178 9.3005
R277 VTAIL.n184 VTAIL.n183 9.3005
R278 VTAIL.n130 VTAIL.n129 9.3005
R279 VTAIL.n89 VTAIL.n88 9.3005
R280 VTAIL.n136 VTAIL.n135 9.3005
R281 VTAIL.n138 VTAIL.n137 9.3005
R282 VTAIL.n85 VTAIL.n84 9.3005
R283 VTAIL.n144 VTAIL.n143 9.3005
R284 VTAIL.n146 VTAIL.n145 9.3005
R285 VTAIL.n82 VTAIL.n79 9.3005
R286 VTAIL.n153 VTAIL.n152 9.3005
R287 VTAIL.n128 VTAIL.n127 9.3005
R288 VTAIL.n93 VTAIL.n92 9.3005
R289 VTAIL.n122 VTAIL.n121 9.3005
R290 VTAIL.n120 VTAIL.n119 9.3005
R291 VTAIL.n97 VTAIL.n96 9.3005
R292 VTAIL.n114 VTAIL.n113 9.3005
R293 VTAIL.n112 VTAIL.n111 9.3005
R294 VTAIL.n101 VTAIL.n100 9.3005
R295 VTAIL.n106 VTAIL.n105 9.3005
R296 VTAIL.n274 VTAIL.n250 8.92171
R297 VTAIL.n290 VTAIL.n289 8.92171
R298 VTAIL.n40 VTAIL.n16 8.92171
R299 VTAIL.n56 VTAIL.n55 8.92171
R300 VTAIL.n213 VTAIL.n212 8.92171
R301 VTAIL.n197 VTAIL.n173 8.92171
R302 VTAIL.n135 VTAIL.n134 8.92171
R303 VTAIL.n119 VTAIL.n95 8.92171
R304 VTAIL.n278 VTAIL.n277 8.14595
R305 VTAIL.n286 VTAIL.n244 8.14595
R306 VTAIL.n44 VTAIL.n43 8.14595
R307 VTAIL.n52 VTAIL.n10 8.14595
R308 VTAIL.n209 VTAIL.n167 8.14595
R309 VTAIL.n201 VTAIL.n200 8.14595
R310 VTAIL.n131 VTAIL.n89 8.14595
R311 VTAIL.n123 VTAIL.n122 8.14595
R312 VTAIL.n281 VTAIL.n248 7.3702
R313 VTAIL.n285 VTAIL.n246 7.3702
R314 VTAIL.n47 VTAIL.n14 7.3702
R315 VTAIL.n51 VTAIL.n12 7.3702
R316 VTAIL.n208 VTAIL.n169 7.3702
R317 VTAIL.n204 VTAIL.n171 7.3702
R318 VTAIL.n130 VTAIL.n91 7.3702
R319 VTAIL.n126 VTAIL.n93 7.3702
R320 VTAIL.n282 VTAIL.n281 6.59444
R321 VTAIL.n282 VTAIL.n246 6.59444
R322 VTAIL.n48 VTAIL.n47 6.59444
R323 VTAIL.n48 VTAIL.n12 6.59444
R324 VTAIL.n205 VTAIL.n169 6.59444
R325 VTAIL.n205 VTAIL.n204 6.59444
R326 VTAIL.n127 VTAIL.n91 6.59444
R327 VTAIL.n127 VTAIL.n126 6.59444
R328 VTAIL.n278 VTAIL.n248 5.81868
R329 VTAIL.n286 VTAIL.n285 5.81868
R330 VTAIL.n44 VTAIL.n14 5.81868
R331 VTAIL.n52 VTAIL.n51 5.81868
R332 VTAIL.n209 VTAIL.n208 5.81868
R333 VTAIL.n201 VTAIL.n171 5.81868
R334 VTAIL.n131 VTAIL.n130 5.81868
R335 VTAIL.n123 VTAIL.n93 5.81868
R336 VTAIL.n277 VTAIL.n250 5.04292
R337 VTAIL.n289 VTAIL.n244 5.04292
R338 VTAIL.n43 VTAIL.n16 5.04292
R339 VTAIL.n55 VTAIL.n10 5.04292
R340 VTAIL.n212 VTAIL.n167 5.04292
R341 VTAIL.n200 VTAIL.n173 5.04292
R342 VTAIL.n134 VTAIL.n89 5.04292
R343 VTAIL.n122 VTAIL.n95 5.04292
R344 VTAIL.n260 VTAIL.n259 4.38563
R345 VTAIL.n26 VTAIL.n25 4.38563
R346 VTAIL.n183 VTAIL.n182 4.38563
R347 VTAIL.n105 VTAIL.n104 4.38563
R348 VTAIL.n274 VTAIL.n273 4.26717
R349 VTAIL.n290 VTAIL.n242 4.26717
R350 VTAIL.n40 VTAIL.n39 4.26717
R351 VTAIL.n56 VTAIL.n8 4.26717
R352 VTAIL.n213 VTAIL.n165 4.26717
R353 VTAIL.n197 VTAIL.n196 4.26717
R354 VTAIL.n135 VTAIL.n87 4.26717
R355 VTAIL.n119 VTAIL.n118 4.26717
R356 VTAIL.n270 VTAIL.n252 3.49141
R357 VTAIL.n294 VTAIL.n293 3.49141
R358 VTAIL.n36 VTAIL.n18 3.49141
R359 VTAIL.n60 VTAIL.n59 3.49141
R360 VTAIL.n217 VTAIL.n216 3.49141
R361 VTAIL.n193 VTAIL.n175 3.49141
R362 VTAIL.n139 VTAIL.n138 3.49141
R363 VTAIL.n115 VTAIL.n97 3.49141
R364 VTAIL.n269 VTAIL.n254 2.71565
R365 VTAIL.n297 VTAIL.n240 2.71565
R366 VTAIL.n35 VTAIL.n20 2.71565
R367 VTAIL.n63 VTAIL.n6 2.71565
R368 VTAIL.n220 VTAIL.n163 2.71565
R369 VTAIL.n192 VTAIL.n177 2.71565
R370 VTAIL.n142 VTAIL.n85 2.71565
R371 VTAIL.n114 VTAIL.n99 2.71565
R372 VTAIL.n266 VTAIL.n265 1.93989
R373 VTAIL.n298 VTAIL.n238 1.93989
R374 VTAIL.n32 VTAIL.n31 1.93989
R375 VTAIL.n64 VTAIL.n4 1.93989
R376 VTAIL.n221 VTAIL.n161 1.93989
R377 VTAIL.n189 VTAIL.n188 1.93989
R378 VTAIL.n143 VTAIL.n83 1.93989
R379 VTAIL.n111 VTAIL.n110 1.93989
R380 VTAIL.n262 VTAIL.n256 1.16414
R381 VTAIL.n303 VTAIL.n301 1.16414
R382 VTAIL.n310 VTAIL.n234 1.16414
R383 VTAIL.n28 VTAIL.n22 1.16414
R384 VTAIL.n69 VTAIL.n67 1.16414
R385 VTAIL.n76 VTAIL.n0 1.16414
R386 VTAIL.n232 VTAIL.n156 1.16414
R387 VTAIL.n225 VTAIL.n224 1.16414
R388 VTAIL.n185 VTAIL.n179 1.16414
R389 VTAIL.n154 VTAIL.n78 1.16414
R390 VTAIL.n147 VTAIL.n146 1.16414
R391 VTAIL.n107 VTAIL.n101 1.16414
R392 VTAIL.n233 VTAIL.n155 0.970328
R393 VTAIL VTAIL.n77 0.778517
R394 VTAIL.n261 VTAIL.n258 0.388379
R395 VTAIL.n302 VTAIL.n236 0.388379
R396 VTAIL.n308 VTAIL.n307 0.388379
R397 VTAIL.n27 VTAIL.n24 0.388379
R398 VTAIL.n68 VTAIL.n2 0.388379
R399 VTAIL.n74 VTAIL.n73 0.388379
R400 VTAIL.n230 VTAIL.n229 0.388379
R401 VTAIL.n160 VTAIL.n158 0.388379
R402 VTAIL.n184 VTAIL.n181 0.388379
R403 VTAIL.n152 VTAIL.n151 0.388379
R404 VTAIL.n82 VTAIL.n80 0.388379
R405 VTAIL.n106 VTAIL.n103 0.388379
R406 VTAIL VTAIL.n311 0.19231
R407 VTAIL.n260 VTAIL.n255 0.155672
R408 VTAIL.n267 VTAIL.n255 0.155672
R409 VTAIL.n268 VTAIL.n267 0.155672
R410 VTAIL.n268 VTAIL.n251 0.155672
R411 VTAIL.n275 VTAIL.n251 0.155672
R412 VTAIL.n276 VTAIL.n275 0.155672
R413 VTAIL.n276 VTAIL.n247 0.155672
R414 VTAIL.n283 VTAIL.n247 0.155672
R415 VTAIL.n284 VTAIL.n283 0.155672
R416 VTAIL.n284 VTAIL.n243 0.155672
R417 VTAIL.n291 VTAIL.n243 0.155672
R418 VTAIL.n292 VTAIL.n291 0.155672
R419 VTAIL.n292 VTAIL.n239 0.155672
R420 VTAIL.n299 VTAIL.n239 0.155672
R421 VTAIL.n300 VTAIL.n299 0.155672
R422 VTAIL.n300 VTAIL.n235 0.155672
R423 VTAIL.n309 VTAIL.n235 0.155672
R424 VTAIL.n26 VTAIL.n21 0.155672
R425 VTAIL.n33 VTAIL.n21 0.155672
R426 VTAIL.n34 VTAIL.n33 0.155672
R427 VTAIL.n34 VTAIL.n17 0.155672
R428 VTAIL.n41 VTAIL.n17 0.155672
R429 VTAIL.n42 VTAIL.n41 0.155672
R430 VTAIL.n42 VTAIL.n13 0.155672
R431 VTAIL.n49 VTAIL.n13 0.155672
R432 VTAIL.n50 VTAIL.n49 0.155672
R433 VTAIL.n50 VTAIL.n9 0.155672
R434 VTAIL.n57 VTAIL.n9 0.155672
R435 VTAIL.n58 VTAIL.n57 0.155672
R436 VTAIL.n58 VTAIL.n5 0.155672
R437 VTAIL.n65 VTAIL.n5 0.155672
R438 VTAIL.n66 VTAIL.n65 0.155672
R439 VTAIL.n66 VTAIL.n1 0.155672
R440 VTAIL.n75 VTAIL.n1 0.155672
R441 VTAIL.n231 VTAIL.n157 0.155672
R442 VTAIL.n223 VTAIL.n157 0.155672
R443 VTAIL.n223 VTAIL.n222 0.155672
R444 VTAIL.n222 VTAIL.n162 0.155672
R445 VTAIL.n215 VTAIL.n162 0.155672
R446 VTAIL.n215 VTAIL.n214 0.155672
R447 VTAIL.n214 VTAIL.n166 0.155672
R448 VTAIL.n207 VTAIL.n166 0.155672
R449 VTAIL.n207 VTAIL.n206 0.155672
R450 VTAIL.n206 VTAIL.n170 0.155672
R451 VTAIL.n199 VTAIL.n170 0.155672
R452 VTAIL.n199 VTAIL.n198 0.155672
R453 VTAIL.n198 VTAIL.n174 0.155672
R454 VTAIL.n191 VTAIL.n174 0.155672
R455 VTAIL.n191 VTAIL.n190 0.155672
R456 VTAIL.n190 VTAIL.n178 0.155672
R457 VTAIL.n183 VTAIL.n178 0.155672
R458 VTAIL.n153 VTAIL.n79 0.155672
R459 VTAIL.n145 VTAIL.n79 0.155672
R460 VTAIL.n145 VTAIL.n144 0.155672
R461 VTAIL.n144 VTAIL.n84 0.155672
R462 VTAIL.n137 VTAIL.n84 0.155672
R463 VTAIL.n137 VTAIL.n136 0.155672
R464 VTAIL.n136 VTAIL.n88 0.155672
R465 VTAIL.n129 VTAIL.n88 0.155672
R466 VTAIL.n129 VTAIL.n128 0.155672
R467 VTAIL.n128 VTAIL.n92 0.155672
R468 VTAIL.n121 VTAIL.n92 0.155672
R469 VTAIL.n121 VTAIL.n120 0.155672
R470 VTAIL.n120 VTAIL.n96 0.155672
R471 VTAIL.n113 VTAIL.n96 0.155672
R472 VTAIL.n113 VTAIL.n112 0.155672
R473 VTAIL.n112 VTAIL.n100 0.155672
R474 VTAIL.n105 VTAIL.n100 0.155672
R475 VDD2.n149 VDD2.n77 289.615
R476 VDD2.n72 VDD2.n0 289.615
R477 VDD2.n150 VDD2.n149 185
R478 VDD2.n148 VDD2.n79 185
R479 VDD2.n147 VDD2.n146 185
R480 VDD2.n82 VDD2.n80 185
R481 VDD2.n141 VDD2.n140 185
R482 VDD2.n139 VDD2.n138 185
R483 VDD2.n86 VDD2.n85 185
R484 VDD2.n133 VDD2.n132 185
R485 VDD2.n131 VDD2.n130 185
R486 VDD2.n90 VDD2.n89 185
R487 VDD2.n125 VDD2.n124 185
R488 VDD2.n123 VDD2.n122 185
R489 VDD2.n94 VDD2.n93 185
R490 VDD2.n117 VDD2.n116 185
R491 VDD2.n115 VDD2.n114 185
R492 VDD2.n98 VDD2.n97 185
R493 VDD2.n109 VDD2.n108 185
R494 VDD2.n107 VDD2.n106 185
R495 VDD2.n102 VDD2.n101 185
R496 VDD2.n24 VDD2.n23 185
R497 VDD2.n29 VDD2.n28 185
R498 VDD2.n31 VDD2.n30 185
R499 VDD2.n20 VDD2.n19 185
R500 VDD2.n37 VDD2.n36 185
R501 VDD2.n39 VDD2.n38 185
R502 VDD2.n16 VDD2.n15 185
R503 VDD2.n45 VDD2.n44 185
R504 VDD2.n47 VDD2.n46 185
R505 VDD2.n12 VDD2.n11 185
R506 VDD2.n53 VDD2.n52 185
R507 VDD2.n55 VDD2.n54 185
R508 VDD2.n8 VDD2.n7 185
R509 VDD2.n61 VDD2.n60 185
R510 VDD2.n63 VDD2.n62 185
R511 VDD2.n4 VDD2.n3 185
R512 VDD2.n70 VDD2.n69 185
R513 VDD2.n71 VDD2.n2 185
R514 VDD2.n73 VDD2.n72 185
R515 VDD2.n103 VDD2.t1 147.659
R516 VDD2.n25 VDD2.t0 147.659
R517 VDD2.n149 VDD2.n148 104.615
R518 VDD2.n148 VDD2.n147 104.615
R519 VDD2.n147 VDD2.n80 104.615
R520 VDD2.n140 VDD2.n80 104.615
R521 VDD2.n140 VDD2.n139 104.615
R522 VDD2.n139 VDD2.n85 104.615
R523 VDD2.n132 VDD2.n85 104.615
R524 VDD2.n132 VDD2.n131 104.615
R525 VDD2.n131 VDD2.n89 104.615
R526 VDD2.n124 VDD2.n89 104.615
R527 VDD2.n124 VDD2.n123 104.615
R528 VDD2.n123 VDD2.n93 104.615
R529 VDD2.n116 VDD2.n93 104.615
R530 VDD2.n116 VDD2.n115 104.615
R531 VDD2.n115 VDD2.n97 104.615
R532 VDD2.n108 VDD2.n97 104.615
R533 VDD2.n108 VDD2.n107 104.615
R534 VDD2.n107 VDD2.n101 104.615
R535 VDD2.n29 VDD2.n23 104.615
R536 VDD2.n30 VDD2.n29 104.615
R537 VDD2.n30 VDD2.n19 104.615
R538 VDD2.n37 VDD2.n19 104.615
R539 VDD2.n38 VDD2.n37 104.615
R540 VDD2.n38 VDD2.n15 104.615
R541 VDD2.n45 VDD2.n15 104.615
R542 VDD2.n46 VDD2.n45 104.615
R543 VDD2.n46 VDD2.n11 104.615
R544 VDD2.n53 VDD2.n11 104.615
R545 VDD2.n54 VDD2.n53 104.615
R546 VDD2.n54 VDD2.n7 104.615
R547 VDD2.n61 VDD2.n7 104.615
R548 VDD2.n62 VDD2.n61 104.615
R549 VDD2.n62 VDD2.n3 104.615
R550 VDD2.n70 VDD2.n3 104.615
R551 VDD2.n71 VDD2.n70 104.615
R552 VDD2.n72 VDD2.n71 104.615
R553 VDD2.n154 VDD2.n76 88.769
R554 VDD2.t1 VDD2.n101 52.3082
R555 VDD2.t0 VDD2.n23 52.3082
R556 VDD2.n154 VDD2.n153 50.9975
R557 VDD2.n103 VDD2.n102 15.6677
R558 VDD2.n25 VDD2.n24 15.6677
R559 VDD2.n150 VDD2.n79 13.1884
R560 VDD2.n73 VDD2.n2 13.1884
R561 VDD2.n151 VDD2.n77 12.8005
R562 VDD2.n146 VDD2.n81 12.8005
R563 VDD2.n106 VDD2.n105 12.8005
R564 VDD2.n28 VDD2.n27 12.8005
R565 VDD2.n69 VDD2.n68 12.8005
R566 VDD2.n74 VDD2.n0 12.8005
R567 VDD2.n145 VDD2.n82 12.0247
R568 VDD2.n109 VDD2.n100 12.0247
R569 VDD2.n31 VDD2.n22 12.0247
R570 VDD2.n67 VDD2.n4 12.0247
R571 VDD2.n142 VDD2.n141 11.249
R572 VDD2.n110 VDD2.n98 11.249
R573 VDD2.n32 VDD2.n20 11.249
R574 VDD2.n64 VDD2.n63 11.249
R575 VDD2.n138 VDD2.n84 10.4732
R576 VDD2.n114 VDD2.n113 10.4732
R577 VDD2.n36 VDD2.n35 10.4732
R578 VDD2.n60 VDD2.n6 10.4732
R579 VDD2.n137 VDD2.n86 9.69747
R580 VDD2.n117 VDD2.n96 9.69747
R581 VDD2.n39 VDD2.n18 9.69747
R582 VDD2.n59 VDD2.n8 9.69747
R583 VDD2.n153 VDD2.n152 9.45567
R584 VDD2.n76 VDD2.n75 9.45567
R585 VDD2.n129 VDD2.n128 9.3005
R586 VDD2.n88 VDD2.n87 9.3005
R587 VDD2.n135 VDD2.n134 9.3005
R588 VDD2.n137 VDD2.n136 9.3005
R589 VDD2.n84 VDD2.n83 9.3005
R590 VDD2.n143 VDD2.n142 9.3005
R591 VDD2.n145 VDD2.n144 9.3005
R592 VDD2.n81 VDD2.n78 9.3005
R593 VDD2.n152 VDD2.n151 9.3005
R594 VDD2.n127 VDD2.n126 9.3005
R595 VDD2.n92 VDD2.n91 9.3005
R596 VDD2.n121 VDD2.n120 9.3005
R597 VDD2.n119 VDD2.n118 9.3005
R598 VDD2.n96 VDD2.n95 9.3005
R599 VDD2.n113 VDD2.n112 9.3005
R600 VDD2.n111 VDD2.n110 9.3005
R601 VDD2.n100 VDD2.n99 9.3005
R602 VDD2.n105 VDD2.n104 9.3005
R603 VDD2.n75 VDD2.n74 9.3005
R604 VDD2.n14 VDD2.n13 9.3005
R605 VDD2.n43 VDD2.n42 9.3005
R606 VDD2.n41 VDD2.n40 9.3005
R607 VDD2.n18 VDD2.n17 9.3005
R608 VDD2.n35 VDD2.n34 9.3005
R609 VDD2.n33 VDD2.n32 9.3005
R610 VDD2.n22 VDD2.n21 9.3005
R611 VDD2.n27 VDD2.n26 9.3005
R612 VDD2.n49 VDD2.n48 9.3005
R613 VDD2.n51 VDD2.n50 9.3005
R614 VDD2.n10 VDD2.n9 9.3005
R615 VDD2.n57 VDD2.n56 9.3005
R616 VDD2.n59 VDD2.n58 9.3005
R617 VDD2.n6 VDD2.n5 9.3005
R618 VDD2.n65 VDD2.n64 9.3005
R619 VDD2.n67 VDD2.n66 9.3005
R620 VDD2.n68 VDD2.n1 9.3005
R621 VDD2.n134 VDD2.n133 8.92171
R622 VDD2.n118 VDD2.n94 8.92171
R623 VDD2.n40 VDD2.n16 8.92171
R624 VDD2.n56 VDD2.n55 8.92171
R625 VDD2.n130 VDD2.n88 8.14595
R626 VDD2.n122 VDD2.n121 8.14595
R627 VDD2.n44 VDD2.n43 8.14595
R628 VDD2.n52 VDD2.n10 8.14595
R629 VDD2.n129 VDD2.n90 7.3702
R630 VDD2.n125 VDD2.n92 7.3702
R631 VDD2.n47 VDD2.n14 7.3702
R632 VDD2.n51 VDD2.n12 7.3702
R633 VDD2.n126 VDD2.n90 6.59444
R634 VDD2.n126 VDD2.n125 6.59444
R635 VDD2.n48 VDD2.n47 6.59444
R636 VDD2.n48 VDD2.n12 6.59444
R637 VDD2.n130 VDD2.n129 5.81868
R638 VDD2.n122 VDD2.n92 5.81868
R639 VDD2.n44 VDD2.n14 5.81868
R640 VDD2.n52 VDD2.n51 5.81868
R641 VDD2.n133 VDD2.n88 5.04292
R642 VDD2.n121 VDD2.n94 5.04292
R643 VDD2.n43 VDD2.n16 5.04292
R644 VDD2.n55 VDD2.n10 5.04292
R645 VDD2.n104 VDD2.n103 4.38563
R646 VDD2.n26 VDD2.n25 4.38563
R647 VDD2.n134 VDD2.n86 4.26717
R648 VDD2.n118 VDD2.n117 4.26717
R649 VDD2.n40 VDD2.n39 4.26717
R650 VDD2.n56 VDD2.n8 4.26717
R651 VDD2.n138 VDD2.n137 3.49141
R652 VDD2.n114 VDD2.n96 3.49141
R653 VDD2.n36 VDD2.n18 3.49141
R654 VDD2.n60 VDD2.n59 3.49141
R655 VDD2.n141 VDD2.n84 2.71565
R656 VDD2.n113 VDD2.n98 2.71565
R657 VDD2.n35 VDD2.n20 2.71565
R658 VDD2.n63 VDD2.n6 2.71565
R659 VDD2.n142 VDD2.n82 1.93989
R660 VDD2.n110 VDD2.n109 1.93989
R661 VDD2.n32 VDD2.n31 1.93989
R662 VDD2.n64 VDD2.n4 1.93989
R663 VDD2.n153 VDD2.n77 1.16414
R664 VDD2.n146 VDD2.n145 1.16414
R665 VDD2.n106 VDD2.n100 1.16414
R666 VDD2.n28 VDD2.n22 1.16414
R667 VDD2.n69 VDD2.n67 1.16414
R668 VDD2.n76 VDD2.n0 1.16414
R669 VDD2.n151 VDD2.n150 0.388379
R670 VDD2.n81 VDD2.n79 0.388379
R671 VDD2.n105 VDD2.n102 0.388379
R672 VDD2.n27 VDD2.n24 0.388379
R673 VDD2.n68 VDD2.n2 0.388379
R674 VDD2.n74 VDD2.n73 0.388379
R675 VDD2 VDD2.n154 0.30869
R676 VDD2.n152 VDD2.n78 0.155672
R677 VDD2.n144 VDD2.n78 0.155672
R678 VDD2.n144 VDD2.n143 0.155672
R679 VDD2.n143 VDD2.n83 0.155672
R680 VDD2.n136 VDD2.n83 0.155672
R681 VDD2.n136 VDD2.n135 0.155672
R682 VDD2.n135 VDD2.n87 0.155672
R683 VDD2.n128 VDD2.n87 0.155672
R684 VDD2.n128 VDD2.n127 0.155672
R685 VDD2.n127 VDD2.n91 0.155672
R686 VDD2.n120 VDD2.n91 0.155672
R687 VDD2.n120 VDD2.n119 0.155672
R688 VDD2.n119 VDD2.n95 0.155672
R689 VDD2.n112 VDD2.n95 0.155672
R690 VDD2.n112 VDD2.n111 0.155672
R691 VDD2.n111 VDD2.n99 0.155672
R692 VDD2.n104 VDD2.n99 0.155672
R693 VDD2.n26 VDD2.n21 0.155672
R694 VDD2.n33 VDD2.n21 0.155672
R695 VDD2.n34 VDD2.n33 0.155672
R696 VDD2.n34 VDD2.n17 0.155672
R697 VDD2.n41 VDD2.n17 0.155672
R698 VDD2.n42 VDD2.n41 0.155672
R699 VDD2.n42 VDD2.n13 0.155672
R700 VDD2.n49 VDD2.n13 0.155672
R701 VDD2.n50 VDD2.n49 0.155672
R702 VDD2.n50 VDD2.n9 0.155672
R703 VDD2.n57 VDD2.n9 0.155672
R704 VDD2.n58 VDD2.n57 0.155672
R705 VDD2.n58 VDD2.n5 0.155672
R706 VDD2.n65 VDD2.n5 0.155672
R707 VDD2.n66 VDD2.n65 0.155672
R708 VDD2.n66 VDD2.n1 0.155672
R709 VDD2.n75 VDD2.n1 0.155672
R710 B.n379 B.t13 608.995
R711 B.n377 B.t9 608.995
R712 B.n88 B.t2 608.995
R713 B.n86 B.t6 608.995
R714 B.n656 B.n655 585
R715 B.n657 B.n656 585
R716 B.n294 B.n84 585
R717 B.n293 B.n292 585
R718 B.n291 B.n290 585
R719 B.n289 B.n288 585
R720 B.n287 B.n286 585
R721 B.n285 B.n284 585
R722 B.n283 B.n282 585
R723 B.n281 B.n280 585
R724 B.n279 B.n278 585
R725 B.n277 B.n276 585
R726 B.n275 B.n274 585
R727 B.n273 B.n272 585
R728 B.n271 B.n270 585
R729 B.n269 B.n268 585
R730 B.n267 B.n266 585
R731 B.n265 B.n264 585
R732 B.n263 B.n262 585
R733 B.n261 B.n260 585
R734 B.n259 B.n258 585
R735 B.n257 B.n256 585
R736 B.n255 B.n254 585
R737 B.n253 B.n252 585
R738 B.n251 B.n250 585
R739 B.n249 B.n248 585
R740 B.n247 B.n246 585
R741 B.n245 B.n244 585
R742 B.n243 B.n242 585
R743 B.n241 B.n240 585
R744 B.n239 B.n238 585
R745 B.n237 B.n236 585
R746 B.n235 B.n234 585
R747 B.n233 B.n232 585
R748 B.n231 B.n230 585
R749 B.n229 B.n228 585
R750 B.n227 B.n226 585
R751 B.n225 B.n224 585
R752 B.n223 B.n222 585
R753 B.n221 B.n220 585
R754 B.n219 B.n218 585
R755 B.n217 B.n216 585
R756 B.n215 B.n214 585
R757 B.n213 B.n212 585
R758 B.n211 B.n210 585
R759 B.n209 B.n208 585
R760 B.n207 B.n206 585
R761 B.n205 B.n204 585
R762 B.n203 B.n202 585
R763 B.n200 B.n199 585
R764 B.n198 B.n197 585
R765 B.n196 B.n195 585
R766 B.n194 B.n193 585
R767 B.n192 B.n191 585
R768 B.n190 B.n189 585
R769 B.n188 B.n187 585
R770 B.n186 B.n185 585
R771 B.n184 B.n183 585
R772 B.n182 B.n181 585
R773 B.n180 B.n179 585
R774 B.n178 B.n177 585
R775 B.n176 B.n175 585
R776 B.n174 B.n173 585
R777 B.n172 B.n171 585
R778 B.n170 B.n169 585
R779 B.n168 B.n167 585
R780 B.n166 B.n165 585
R781 B.n164 B.n163 585
R782 B.n162 B.n161 585
R783 B.n160 B.n159 585
R784 B.n158 B.n157 585
R785 B.n156 B.n155 585
R786 B.n154 B.n153 585
R787 B.n152 B.n151 585
R788 B.n150 B.n149 585
R789 B.n148 B.n147 585
R790 B.n146 B.n145 585
R791 B.n144 B.n143 585
R792 B.n142 B.n141 585
R793 B.n140 B.n139 585
R794 B.n138 B.n137 585
R795 B.n136 B.n135 585
R796 B.n134 B.n133 585
R797 B.n132 B.n131 585
R798 B.n130 B.n129 585
R799 B.n128 B.n127 585
R800 B.n126 B.n125 585
R801 B.n124 B.n123 585
R802 B.n122 B.n121 585
R803 B.n120 B.n119 585
R804 B.n118 B.n117 585
R805 B.n116 B.n115 585
R806 B.n114 B.n113 585
R807 B.n112 B.n111 585
R808 B.n110 B.n109 585
R809 B.n108 B.n107 585
R810 B.n106 B.n105 585
R811 B.n104 B.n103 585
R812 B.n102 B.n101 585
R813 B.n100 B.n99 585
R814 B.n98 B.n97 585
R815 B.n96 B.n95 585
R816 B.n94 B.n93 585
R817 B.n92 B.n91 585
R818 B.n32 B.n31 585
R819 B.n660 B.n659 585
R820 B.n654 B.n85 585
R821 B.n85 B.n29 585
R822 B.n653 B.n28 585
R823 B.n664 B.n28 585
R824 B.n652 B.n27 585
R825 B.n665 B.n27 585
R826 B.n651 B.n26 585
R827 B.n666 B.n26 585
R828 B.n650 B.n649 585
R829 B.n649 B.n22 585
R830 B.n648 B.n21 585
R831 B.n672 B.n21 585
R832 B.n647 B.n20 585
R833 B.n673 B.n20 585
R834 B.n646 B.n19 585
R835 B.n674 B.n19 585
R836 B.n645 B.n644 585
R837 B.n644 B.n15 585
R838 B.n643 B.n14 585
R839 B.n680 B.n14 585
R840 B.n642 B.n13 585
R841 B.n681 B.n13 585
R842 B.n641 B.n12 585
R843 B.n682 B.n12 585
R844 B.n640 B.n639 585
R845 B.n639 B.n8 585
R846 B.n638 B.n7 585
R847 B.n688 B.n7 585
R848 B.n637 B.n6 585
R849 B.n689 B.n6 585
R850 B.n636 B.n5 585
R851 B.n690 B.n5 585
R852 B.n635 B.n634 585
R853 B.n634 B.n4 585
R854 B.n633 B.n295 585
R855 B.n633 B.n632 585
R856 B.n623 B.n296 585
R857 B.n297 B.n296 585
R858 B.n625 B.n624 585
R859 B.n626 B.n625 585
R860 B.n622 B.n302 585
R861 B.n302 B.n301 585
R862 B.n621 B.n620 585
R863 B.n620 B.n619 585
R864 B.n304 B.n303 585
R865 B.n305 B.n304 585
R866 B.n612 B.n611 585
R867 B.n613 B.n612 585
R868 B.n610 B.n310 585
R869 B.n310 B.n309 585
R870 B.n609 B.n608 585
R871 B.n608 B.n607 585
R872 B.n312 B.n311 585
R873 B.n313 B.n312 585
R874 B.n600 B.n599 585
R875 B.n601 B.n600 585
R876 B.n598 B.n318 585
R877 B.n318 B.n317 585
R878 B.n597 B.n596 585
R879 B.n596 B.n595 585
R880 B.n320 B.n319 585
R881 B.n321 B.n320 585
R882 B.n591 B.n590 585
R883 B.n324 B.n323 585
R884 B.n587 B.n586 585
R885 B.n588 B.n587 585
R886 B.n585 B.n376 585
R887 B.n584 B.n583 585
R888 B.n582 B.n581 585
R889 B.n580 B.n579 585
R890 B.n578 B.n577 585
R891 B.n576 B.n575 585
R892 B.n574 B.n573 585
R893 B.n572 B.n571 585
R894 B.n570 B.n569 585
R895 B.n568 B.n567 585
R896 B.n566 B.n565 585
R897 B.n564 B.n563 585
R898 B.n562 B.n561 585
R899 B.n560 B.n559 585
R900 B.n558 B.n557 585
R901 B.n556 B.n555 585
R902 B.n554 B.n553 585
R903 B.n552 B.n551 585
R904 B.n550 B.n549 585
R905 B.n548 B.n547 585
R906 B.n546 B.n545 585
R907 B.n544 B.n543 585
R908 B.n542 B.n541 585
R909 B.n540 B.n539 585
R910 B.n538 B.n537 585
R911 B.n536 B.n535 585
R912 B.n534 B.n533 585
R913 B.n532 B.n531 585
R914 B.n530 B.n529 585
R915 B.n528 B.n527 585
R916 B.n526 B.n525 585
R917 B.n524 B.n523 585
R918 B.n522 B.n521 585
R919 B.n520 B.n519 585
R920 B.n518 B.n517 585
R921 B.n516 B.n515 585
R922 B.n514 B.n513 585
R923 B.n512 B.n511 585
R924 B.n510 B.n509 585
R925 B.n508 B.n507 585
R926 B.n506 B.n505 585
R927 B.n504 B.n503 585
R928 B.n502 B.n501 585
R929 B.n500 B.n499 585
R930 B.n498 B.n497 585
R931 B.n495 B.n494 585
R932 B.n493 B.n492 585
R933 B.n491 B.n490 585
R934 B.n489 B.n488 585
R935 B.n487 B.n486 585
R936 B.n485 B.n484 585
R937 B.n483 B.n482 585
R938 B.n481 B.n480 585
R939 B.n479 B.n478 585
R940 B.n477 B.n476 585
R941 B.n475 B.n474 585
R942 B.n473 B.n472 585
R943 B.n471 B.n470 585
R944 B.n469 B.n468 585
R945 B.n467 B.n466 585
R946 B.n465 B.n464 585
R947 B.n463 B.n462 585
R948 B.n461 B.n460 585
R949 B.n459 B.n458 585
R950 B.n457 B.n456 585
R951 B.n455 B.n454 585
R952 B.n453 B.n452 585
R953 B.n451 B.n450 585
R954 B.n449 B.n448 585
R955 B.n447 B.n446 585
R956 B.n445 B.n444 585
R957 B.n443 B.n442 585
R958 B.n441 B.n440 585
R959 B.n439 B.n438 585
R960 B.n437 B.n436 585
R961 B.n435 B.n434 585
R962 B.n433 B.n432 585
R963 B.n431 B.n430 585
R964 B.n429 B.n428 585
R965 B.n427 B.n426 585
R966 B.n425 B.n424 585
R967 B.n423 B.n422 585
R968 B.n421 B.n420 585
R969 B.n419 B.n418 585
R970 B.n417 B.n416 585
R971 B.n415 B.n414 585
R972 B.n413 B.n412 585
R973 B.n411 B.n410 585
R974 B.n409 B.n408 585
R975 B.n407 B.n406 585
R976 B.n405 B.n404 585
R977 B.n403 B.n402 585
R978 B.n401 B.n400 585
R979 B.n399 B.n398 585
R980 B.n397 B.n396 585
R981 B.n395 B.n394 585
R982 B.n393 B.n392 585
R983 B.n391 B.n390 585
R984 B.n389 B.n388 585
R985 B.n387 B.n386 585
R986 B.n385 B.n384 585
R987 B.n383 B.n382 585
R988 B.n592 B.n322 585
R989 B.n322 B.n321 585
R990 B.n594 B.n593 585
R991 B.n595 B.n594 585
R992 B.n316 B.n315 585
R993 B.n317 B.n316 585
R994 B.n603 B.n602 585
R995 B.n602 B.n601 585
R996 B.n604 B.n314 585
R997 B.n314 B.n313 585
R998 B.n606 B.n605 585
R999 B.n607 B.n606 585
R1000 B.n308 B.n307 585
R1001 B.n309 B.n308 585
R1002 B.n615 B.n614 585
R1003 B.n614 B.n613 585
R1004 B.n616 B.n306 585
R1005 B.n306 B.n305 585
R1006 B.n618 B.n617 585
R1007 B.n619 B.n618 585
R1008 B.n300 B.n299 585
R1009 B.n301 B.n300 585
R1010 B.n628 B.n627 585
R1011 B.n627 B.n626 585
R1012 B.n629 B.n298 585
R1013 B.n298 B.n297 585
R1014 B.n631 B.n630 585
R1015 B.n632 B.n631 585
R1016 B.n2 B.n0 585
R1017 B.n4 B.n2 585
R1018 B.n3 B.n1 585
R1019 B.n689 B.n3 585
R1020 B.n687 B.n686 585
R1021 B.n688 B.n687 585
R1022 B.n685 B.n9 585
R1023 B.n9 B.n8 585
R1024 B.n684 B.n683 585
R1025 B.n683 B.n682 585
R1026 B.n11 B.n10 585
R1027 B.n681 B.n11 585
R1028 B.n679 B.n678 585
R1029 B.n680 B.n679 585
R1030 B.n677 B.n16 585
R1031 B.n16 B.n15 585
R1032 B.n676 B.n675 585
R1033 B.n675 B.n674 585
R1034 B.n18 B.n17 585
R1035 B.n673 B.n18 585
R1036 B.n671 B.n670 585
R1037 B.n672 B.n671 585
R1038 B.n669 B.n23 585
R1039 B.n23 B.n22 585
R1040 B.n668 B.n667 585
R1041 B.n667 B.n666 585
R1042 B.n25 B.n24 585
R1043 B.n665 B.n25 585
R1044 B.n663 B.n662 585
R1045 B.n664 B.n663 585
R1046 B.n661 B.n30 585
R1047 B.n30 B.n29 585
R1048 B.n692 B.n691 585
R1049 B.n691 B.n690 585
R1050 B.n590 B.n322 478.086
R1051 B.n659 B.n30 478.086
R1052 B.n382 B.n320 478.086
R1053 B.n656 B.n85 478.086
R1054 B.n379 B.t15 339.449
R1055 B.n86 B.t7 339.449
R1056 B.n377 B.t12 339.449
R1057 B.n88 B.t4 339.449
R1058 B.n380 B.t14 316.952
R1059 B.n87 B.t8 316.952
R1060 B.n378 B.t11 316.952
R1061 B.n89 B.t5 316.952
R1062 B.n657 B.n83 256.663
R1063 B.n657 B.n82 256.663
R1064 B.n657 B.n81 256.663
R1065 B.n657 B.n80 256.663
R1066 B.n657 B.n79 256.663
R1067 B.n657 B.n78 256.663
R1068 B.n657 B.n77 256.663
R1069 B.n657 B.n76 256.663
R1070 B.n657 B.n75 256.663
R1071 B.n657 B.n74 256.663
R1072 B.n657 B.n73 256.663
R1073 B.n657 B.n72 256.663
R1074 B.n657 B.n71 256.663
R1075 B.n657 B.n70 256.663
R1076 B.n657 B.n69 256.663
R1077 B.n657 B.n68 256.663
R1078 B.n657 B.n67 256.663
R1079 B.n657 B.n66 256.663
R1080 B.n657 B.n65 256.663
R1081 B.n657 B.n64 256.663
R1082 B.n657 B.n63 256.663
R1083 B.n657 B.n62 256.663
R1084 B.n657 B.n61 256.663
R1085 B.n657 B.n60 256.663
R1086 B.n657 B.n59 256.663
R1087 B.n657 B.n58 256.663
R1088 B.n657 B.n57 256.663
R1089 B.n657 B.n56 256.663
R1090 B.n657 B.n55 256.663
R1091 B.n657 B.n54 256.663
R1092 B.n657 B.n53 256.663
R1093 B.n657 B.n52 256.663
R1094 B.n657 B.n51 256.663
R1095 B.n657 B.n50 256.663
R1096 B.n657 B.n49 256.663
R1097 B.n657 B.n48 256.663
R1098 B.n657 B.n47 256.663
R1099 B.n657 B.n46 256.663
R1100 B.n657 B.n45 256.663
R1101 B.n657 B.n44 256.663
R1102 B.n657 B.n43 256.663
R1103 B.n657 B.n42 256.663
R1104 B.n657 B.n41 256.663
R1105 B.n657 B.n40 256.663
R1106 B.n657 B.n39 256.663
R1107 B.n657 B.n38 256.663
R1108 B.n657 B.n37 256.663
R1109 B.n657 B.n36 256.663
R1110 B.n657 B.n35 256.663
R1111 B.n657 B.n34 256.663
R1112 B.n657 B.n33 256.663
R1113 B.n658 B.n657 256.663
R1114 B.n589 B.n588 256.663
R1115 B.n588 B.n325 256.663
R1116 B.n588 B.n326 256.663
R1117 B.n588 B.n327 256.663
R1118 B.n588 B.n328 256.663
R1119 B.n588 B.n329 256.663
R1120 B.n588 B.n330 256.663
R1121 B.n588 B.n331 256.663
R1122 B.n588 B.n332 256.663
R1123 B.n588 B.n333 256.663
R1124 B.n588 B.n334 256.663
R1125 B.n588 B.n335 256.663
R1126 B.n588 B.n336 256.663
R1127 B.n588 B.n337 256.663
R1128 B.n588 B.n338 256.663
R1129 B.n588 B.n339 256.663
R1130 B.n588 B.n340 256.663
R1131 B.n588 B.n341 256.663
R1132 B.n588 B.n342 256.663
R1133 B.n588 B.n343 256.663
R1134 B.n588 B.n344 256.663
R1135 B.n588 B.n345 256.663
R1136 B.n588 B.n346 256.663
R1137 B.n588 B.n347 256.663
R1138 B.n588 B.n348 256.663
R1139 B.n588 B.n349 256.663
R1140 B.n588 B.n350 256.663
R1141 B.n588 B.n351 256.663
R1142 B.n588 B.n352 256.663
R1143 B.n588 B.n353 256.663
R1144 B.n588 B.n354 256.663
R1145 B.n588 B.n355 256.663
R1146 B.n588 B.n356 256.663
R1147 B.n588 B.n357 256.663
R1148 B.n588 B.n358 256.663
R1149 B.n588 B.n359 256.663
R1150 B.n588 B.n360 256.663
R1151 B.n588 B.n361 256.663
R1152 B.n588 B.n362 256.663
R1153 B.n588 B.n363 256.663
R1154 B.n588 B.n364 256.663
R1155 B.n588 B.n365 256.663
R1156 B.n588 B.n366 256.663
R1157 B.n588 B.n367 256.663
R1158 B.n588 B.n368 256.663
R1159 B.n588 B.n369 256.663
R1160 B.n588 B.n370 256.663
R1161 B.n588 B.n371 256.663
R1162 B.n588 B.n372 256.663
R1163 B.n588 B.n373 256.663
R1164 B.n588 B.n374 256.663
R1165 B.n588 B.n375 256.663
R1166 B.n594 B.n322 163.367
R1167 B.n594 B.n316 163.367
R1168 B.n602 B.n316 163.367
R1169 B.n602 B.n314 163.367
R1170 B.n606 B.n314 163.367
R1171 B.n606 B.n308 163.367
R1172 B.n614 B.n308 163.367
R1173 B.n614 B.n306 163.367
R1174 B.n618 B.n306 163.367
R1175 B.n618 B.n300 163.367
R1176 B.n627 B.n300 163.367
R1177 B.n627 B.n298 163.367
R1178 B.n631 B.n298 163.367
R1179 B.n631 B.n2 163.367
R1180 B.n691 B.n2 163.367
R1181 B.n691 B.n3 163.367
R1182 B.n687 B.n3 163.367
R1183 B.n687 B.n9 163.367
R1184 B.n683 B.n9 163.367
R1185 B.n683 B.n11 163.367
R1186 B.n679 B.n11 163.367
R1187 B.n679 B.n16 163.367
R1188 B.n675 B.n16 163.367
R1189 B.n675 B.n18 163.367
R1190 B.n671 B.n18 163.367
R1191 B.n671 B.n23 163.367
R1192 B.n667 B.n23 163.367
R1193 B.n667 B.n25 163.367
R1194 B.n663 B.n25 163.367
R1195 B.n663 B.n30 163.367
R1196 B.n587 B.n324 163.367
R1197 B.n587 B.n376 163.367
R1198 B.n583 B.n582 163.367
R1199 B.n579 B.n578 163.367
R1200 B.n575 B.n574 163.367
R1201 B.n571 B.n570 163.367
R1202 B.n567 B.n566 163.367
R1203 B.n563 B.n562 163.367
R1204 B.n559 B.n558 163.367
R1205 B.n555 B.n554 163.367
R1206 B.n551 B.n550 163.367
R1207 B.n547 B.n546 163.367
R1208 B.n543 B.n542 163.367
R1209 B.n539 B.n538 163.367
R1210 B.n535 B.n534 163.367
R1211 B.n531 B.n530 163.367
R1212 B.n527 B.n526 163.367
R1213 B.n523 B.n522 163.367
R1214 B.n519 B.n518 163.367
R1215 B.n515 B.n514 163.367
R1216 B.n511 B.n510 163.367
R1217 B.n507 B.n506 163.367
R1218 B.n503 B.n502 163.367
R1219 B.n499 B.n498 163.367
R1220 B.n494 B.n493 163.367
R1221 B.n490 B.n489 163.367
R1222 B.n486 B.n485 163.367
R1223 B.n482 B.n481 163.367
R1224 B.n478 B.n477 163.367
R1225 B.n474 B.n473 163.367
R1226 B.n470 B.n469 163.367
R1227 B.n466 B.n465 163.367
R1228 B.n462 B.n461 163.367
R1229 B.n458 B.n457 163.367
R1230 B.n454 B.n453 163.367
R1231 B.n450 B.n449 163.367
R1232 B.n446 B.n445 163.367
R1233 B.n442 B.n441 163.367
R1234 B.n438 B.n437 163.367
R1235 B.n434 B.n433 163.367
R1236 B.n430 B.n429 163.367
R1237 B.n426 B.n425 163.367
R1238 B.n422 B.n421 163.367
R1239 B.n418 B.n417 163.367
R1240 B.n414 B.n413 163.367
R1241 B.n410 B.n409 163.367
R1242 B.n406 B.n405 163.367
R1243 B.n402 B.n401 163.367
R1244 B.n398 B.n397 163.367
R1245 B.n394 B.n393 163.367
R1246 B.n390 B.n389 163.367
R1247 B.n386 B.n385 163.367
R1248 B.n596 B.n320 163.367
R1249 B.n596 B.n318 163.367
R1250 B.n600 B.n318 163.367
R1251 B.n600 B.n312 163.367
R1252 B.n608 B.n312 163.367
R1253 B.n608 B.n310 163.367
R1254 B.n612 B.n310 163.367
R1255 B.n612 B.n304 163.367
R1256 B.n620 B.n304 163.367
R1257 B.n620 B.n302 163.367
R1258 B.n625 B.n302 163.367
R1259 B.n625 B.n296 163.367
R1260 B.n633 B.n296 163.367
R1261 B.n634 B.n633 163.367
R1262 B.n634 B.n5 163.367
R1263 B.n6 B.n5 163.367
R1264 B.n7 B.n6 163.367
R1265 B.n639 B.n7 163.367
R1266 B.n639 B.n12 163.367
R1267 B.n13 B.n12 163.367
R1268 B.n14 B.n13 163.367
R1269 B.n644 B.n14 163.367
R1270 B.n644 B.n19 163.367
R1271 B.n20 B.n19 163.367
R1272 B.n21 B.n20 163.367
R1273 B.n649 B.n21 163.367
R1274 B.n649 B.n26 163.367
R1275 B.n27 B.n26 163.367
R1276 B.n28 B.n27 163.367
R1277 B.n85 B.n28 163.367
R1278 B.n91 B.n32 163.367
R1279 B.n95 B.n94 163.367
R1280 B.n99 B.n98 163.367
R1281 B.n103 B.n102 163.367
R1282 B.n107 B.n106 163.367
R1283 B.n111 B.n110 163.367
R1284 B.n115 B.n114 163.367
R1285 B.n119 B.n118 163.367
R1286 B.n123 B.n122 163.367
R1287 B.n127 B.n126 163.367
R1288 B.n131 B.n130 163.367
R1289 B.n135 B.n134 163.367
R1290 B.n139 B.n138 163.367
R1291 B.n143 B.n142 163.367
R1292 B.n147 B.n146 163.367
R1293 B.n151 B.n150 163.367
R1294 B.n155 B.n154 163.367
R1295 B.n159 B.n158 163.367
R1296 B.n163 B.n162 163.367
R1297 B.n167 B.n166 163.367
R1298 B.n171 B.n170 163.367
R1299 B.n175 B.n174 163.367
R1300 B.n179 B.n178 163.367
R1301 B.n183 B.n182 163.367
R1302 B.n187 B.n186 163.367
R1303 B.n191 B.n190 163.367
R1304 B.n195 B.n194 163.367
R1305 B.n199 B.n198 163.367
R1306 B.n204 B.n203 163.367
R1307 B.n208 B.n207 163.367
R1308 B.n212 B.n211 163.367
R1309 B.n216 B.n215 163.367
R1310 B.n220 B.n219 163.367
R1311 B.n224 B.n223 163.367
R1312 B.n228 B.n227 163.367
R1313 B.n232 B.n231 163.367
R1314 B.n236 B.n235 163.367
R1315 B.n240 B.n239 163.367
R1316 B.n244 B.n243 163.367
R1317 B.n248 B.n247 163.367
R1318 B.n252 B.n251 163.367
R1319 B.n256 B.n255 163.367
R1320 B.n260 B.n259 163.367
R1321 B.n264 B.n263 163.367
R1322 B.n268 B.n267 163.367
R1323 B.n272 B.n271 163.367
R1324 B.n276 B.n275 163.367
R1325 B.n280 B.n279 163.367
R1326 B.n284 B.n283 163.367
R1327 B.n288 B.n287 163.367
R1328 B.n292 B.n291 163.367
R1329 B.n656 B.n84 163.367
R1330 B.n590 B.n589 71.676
R1331 B.n376 B.n325 71.676
R1332 B.n582 B.n326 71.676
R1333 B.n578 B.n327 71.676
R1334 B.n574 B.n328 71.676
R1335 B.n570 B.n329 71.676
R1336 B.n566 B.n330 71.676
R1337 B.n562 B.n331 71.676
R1338 B.n558 B.n332 71.676
R1339 B.n554 B.n333 71.676
R1340 B.n550 B.n334 71.676
R1341 B.n546 B.n335 71.676
R1342 B.n542 B.n336 71.676
R1343 B.n538 B.n337 71.676
R1344 B.n534 B.n338 71.676
R1345 B.n530 B.n339 71.676
R1346 B.n526 B.n340 71.676
R1347 B.n522 B.n341 71.676
R1348 B.n518 B.n342 71.676
R1349 B.n514 B.n343 71.676
R1350 B.n510 B.n344 71.676
R1351 B.n506 B.n345 71.676
R1352 B.n502 B.n346 71.676
R1353 B.n498 B.n347 71.676
R1354 B.n493 B.n348 71.676
R1355 B.n489 B.n349 71.676
R1356 B.n485 B.n350 71.676
R1357 B.n481 B.n351 71.676
R1358 B.n477 B.n352 71.676
R1359 B.n473 B.n353 71.676
R1360 B.n469 B.n354 71.676
R1361 B.n465 B.n355 71.676
R1362 B.n461 B.n356 71.676
R1363 B.n457 B.n357 71.676
R1364 B.n453 B.n358 71.676
R1365 B.n449 B.n359 71.676
R1366 B.n445 B.n360 71.676
R1367 B.n441 B.n361 71.676
R1368 B.n437 B.n362 71.676
R1369 B.n433 B.n363 71.676
R1370 B.n429 B.n364 71.676
R1371 B.n425 B.n365 71.676
R1372 B.n421 B.n366 71.676
R1373 B.n417 B.n367 71.676
R1374 B.n413 B.n368 71.676
R1375 B.n409 B.n369 71.676
R1376 B.n405 B.n370 71.676
R1377 B.n401 B.n371 71.676
R1378 B.n397 B.n372 71.676
R1379 B.n393 B.n373 71.676
R1380 B.n389 B.n374 71.676
R1381 B.n385 B.n375 71.676
R1382 B.n659 B.n658 71.676
R1383 B.n91 B.n33 71.676
R1384 B.n95 B.n34 71.676
R1385 B.n99 B.n35 71.676
R1386 B.n103 B.n36 71.676
R1387 B.n107 B.n37 71.676
R1388 B.n111 B.n38 71.676
R1389 B.n115 B.n39 71.676
R1390 B.n119 B.n40 71.676
R1391 B.n123 B.n41 71.676
R1392 B.n127 B.n42 71.676
R1393 B.n131 B.n43 71.676
R1394 B.n135 B.n44 71.676
R1395 B.n139 B.n45 71.676
R1396 B.n143 B.n46 71.676
R1397 B.n147 B.n47 71.676
R1398 B.n151 B.n48 71.676
R1399 B.n155 B.n49 71.676
R1400 B.n159 B.n50 71.676
R1401 B.n163 B.n51 71.676
R1402 B.n167 B.n52 71.676
R1403 B.n171 B.n53 71.676
R1404 B.n175 B.n54 71.676
R1405 B.n179 B.n55 71.676
R1406 B.n183 B.n56 71.676
R1407 B.n187 B.n57 71.676
R1408 B.n191 B.n58 71.676
R1409 B.n195 B.n59 71.676
R1410 B.n199 B.n60 71.676
R1411 B.n204 B.n61 71.676
R1412 B.n208 B.n62 71.676
R1413 B.n212 B.n63 71.676
R1414 B.n216 B.n64 71.676
R1415 B.n220 B.n65 71.676
R1416 B.n224 B.n66 71.676
R1417 B.n228 B.n67 71.676
R1418 B.n232 B.n68 71.676
R1419 B.n236 B.n69 71.676
R1420 B.n240 B.n70 71.676
R1421 B.n244 B.n71 71.676
R1422 B.n248 B.n72 71.676
R1423 B.n252 B.n73 71.676
R1424 B.n256 B.n74 71.676
R1425 B.n260 B.n75 71.676
R1426 B.n264 B.n76 71.676
R1427 B.n268 B.n77 71.676
R1428 B.n272 B.n78 71.676
R1429 B.n276 B.n79 71.676
R1430 B.n280 B.n80 71.676
R1431 B.n284 B.n81 71.676
R1432 B.n288 B.n82 71.676
R1433 B.n292 B.n83 71.676
R1434 B.n84 B.n83 71.676
R1435 B.n291 B.n82 71.676
R1436 B.n287 B.n81 71.676
R1437 B.n283 B.n80 71.676
R1438 B.n279 B.n79 71.676
R1439 B.n275 B.n78 71.676
R1440 B.n271 B.n77 71.676
R1441 B.n267 B.n76 71.676
R1442 B.n263 B.n75 71.676
R1443 B.n259 B.n74 71.676
R1444 B.n255 B.n73 71.676
R1445 B.n251 B.n72 71.676
R1446 B.n247 B.n71 71.676
R1447 B.n243 B.n70 71.676
R1448 B.n239 B.n69 71.676
R1449 B.n235 B.n68 71.676
R1450 B.n231 B.n67 71.676
R1451 B.n227 B.n66 71.676
R1452 B.n223 B.n65 71.676
R1453 B.n219 B.n64 71.676
R1454 B.n215 B.n63 71.676
R1455 B.n211 B.n62 71.676
R1456 B.n207 B.n61 71.676
R1457 B.n203 B.n60 71.676
R1458 B.n198 B.n59 71.676
R1459 B.n194 B.n58 71.676
R1460 B.n190 B.n57 71.676
R1461 B.n186 B.n56 71.676
R1462 B.n182 B.n55 71.676
R1463 B.n178 B.n54 71.676
R1464 B.n174 B.n53 71.676
R1465 B.n170 B.n52 71.676
R1466 B.n166 B.n51 71.676
R1467 B.n162 B.n50 71.676
R1468 B.n158 B.n49 71.676
R1469 B.n154 B.n48 71.676
R1470 B.n150 B.n47 71.676
R1471 B.n146 B.n46 71.676
R1472 B.n142 B.n45 71.676
R1473 B.n138 B.n44 71.676
R1474 B.n134 B.n43 71.676
R1475 B.n130 B.n42 71.676
R1476 B.n126 B.n41 71.676
R1477 B.n122 B.n40 71.676
R1478 B.n118 B.n39 71.676
R1479 B.n114 B.n38 71.676
R1480 B.n110 B.n37 71.676
R1481 B.n106 B.n36 71.676
R1482 B.n102 B.n35 71.676
R1483 B.n98 B.n34 71.676
R1484 B.n94 B.n33 71.676
R1485 B.n658 B.n32 71.676
R1486 B.n589 B.n324 71.676
R1487 B.n583 B.n325 71.676
R1488 B.n579 B.n326 71.676
R1489 B.n575 B.n327 71.676
R1490 B.n571 B.n328 71.676
R1491 B.n567 B.n329 71.676
R1492 B.n563 B.n330 71.676
R1493 B.n559 B.n331 71.676
R1494 B.n555 B.n332 71.676
R1495 B.n551 B.n333 71.676
R1496 B.n547 B.n334 71.676
R1497 B.n543 B.n335 71.676
R1498 B.n539 B.n336 71.676
R1499 B.n535 B.n337 71.676
R1500 B.n531 B.n338 71.676
R1501 B.n527 B.n339 71.676
R1502 B.n523 B.n340 71.676
R1503 B.n519 B.n341 71.676
R1504 B.n515 B.n342 71.676
R1505 B.n511 B.n343 71.676
R1506 B.n507 B.n344 71.676
R1507 B.n503 B.n345 71.676
R1508 B.n499 B.n346 71.676
R1509 B.n494 B.n347 71.676
R1510 B.n490 B.n348 71.676
R1511 B.n486 B.n349 71.676
R1512 B.n482 B.n350 71.676
R1513 B.n478 B.n351 71.676
R1514 B.n474 B.n352 71.676
R1515 B.n470 B.n353 71.676
R1516 B.n466 B.n354 71.676
R1517 B.n462 B.n355 71.676
R1518 B.n458 B.n356 71.676
R1519 B.n454 B.n357 71.676
R1520 B.n450 B.n358 71.676
R1521 B.n446 B.n359 71.676
R1522 B.n442 B.n360 71.676
R1523 B.n438 B.n361 71.676
R1524 B.n434 B.n362 71.676
R1525 B.n430 B.n363 71.676
R1526 B.n426 B.n364 71.676
R1527 B.n422 B.n365 71.676
R1528 B.n418 B.n366 71.676
R1529 B.n414 B.n367 71.676
R1530 B.n410 B.n368 71.676
R1531 B.n406 B.n369 71.676
R1532 B.n402 B.n370 71.676
R1533 B.n398 B.n371 71.676
R1534 B.n394 B.n372 71.676
R1535 B.n390 B.n373 71.676
R1536 B.n386 B.n374 71.676
R1537 B.n382 B.n375 71.676
R1538 B.n588 B.n321 67.7366
R1539 B.n657 B.n29 67.7366
R1540 B.n381 B.n380 59.5399
R1541 B.n496 B.n378 59.5399
R1542 B.n90 B.n89 59.5399
R1543 B.n201 B.n87 59.5399
R1544 B.n595 B.n321 38.7068
R1545 B.n595 B.n317 38.7068
R1546 B.n601 B.n317 38.7068
R1547 B.n601 B.n313 38.7068
R1548 B.n607 B.n313 38.7068
R1549 B.n613 B.n309 38.7068
R1550 B.n613 B.n305 38.7068
R1551 B.n619 B.n305 38.7068
R1552 B.n619 B.n301 38.7068
R1553 B.n626 B.n301 38.7068
R1554 B.n632 B.n297 38.7068
R1555 B.n632 B.n4 38.7068
R1556 B.n690 B.n4 38.7068
R1557 B.n690 B.n689 38.7068
R1558 B.n689 B.n688 38.7068
R1559 B.n688 B.n8 38.7068
R1560 B.n682 B.n681 38.7068
R1561 B.n681 B.n680 38.7068
R1562 B.n680 B.n15 38.7068
R1563 B.n674 B.n15 38.7068
R1564 B.n674 B.n673 38.7068
R1565 B.n672 B.n22 38.7068
R1566 B.n666 B.n22 38.7068
R1567 B.n666 B.n665 38.7068
R1568 B.n665 B.n664 38.7068
R1569 B.n664 B.n29 38.7068
R1570 B.t10 B.n309 35.8608
R1571 B.n673 B.t3 35.8608
R1572 B.n661 B.n660 31.0639
R1573 B.n655 B.n654 31.0639
R1574 B.n383 B.n319 31.0639
R1575 B.n592 B.n591 31.0639
R1576 B.n626 B.t1 26.7534
R1577 B.n682 B.t0 26.7534
R1578 B.n380 B.n379 22.4975
R1579 B.n378 B.n377 22.4975
R1580 B.n89 B.n88 22.4975
R1581 B.n87 B.n86 22.4975
R1582 B B.n692 18.0485
R1583 B.t1 B.n297 11.9539
R1584 B.t0 B.n8 11.9539
R1585 B.n660 B.n31 10.6151
R1586 B.n92 B.n31 10.6151
R1587 B.n93 B.n92 10.6151
R1588 B.n96 B.n93 10.6151
R1589 B.n97 B.n96 10.6151
R1590 B.n100 B.n97 10.6151
R1591 B.n101 B.n100 10.6151
R1592 B.n104 B.n101 10.6151
R1593 B.n105 B.n104 10.6151
R1594 B.n108 B.n105 10.6151
R1595 B.n109 B.n108 10.6151
R1596 B.n112 B.n109 10.6151
R1597 B.n113 B.n112 10.6151
R1598 B.n116 B.n113 10.6151
R1599 B.n117 B.n116 10.6151
R1600 B.n120 B.n117 10.6151
R1601 B.n121 B.n120 10.6151
R1602 B.n124 B.n121 10.6151
R1603 B.n125 B.n124 10.6151
R1604 B.n128 B.n125 10.6151
R1605 B.n129 B.n128 10.6151
R1606 B.n132 B.n129 10.6151
R1607 B.n133 B.n132 10.6151
R1608 B.n136 B.n133 10.6151
R1609 B.n137 B.n136 10.6151
R1610 B.n140 B.n137 10.6151
R1611 B.n141 B.n140 10.6151
R1612 B.n144 B.n141 10.6151
R1613 B.n145 B.n144 10.6151
R1614 B.n148 B.n145 10.6151
R1615 B.n149 B.n148 10.6151
R1616 B.n152 B.n149 10.6151
R1617 B.n153 B.n152 10.6151
R1618 B.n156 B.n153 10.6151
R1619 B.n157 B.n156 10.6151
R1620 B.n160 B.n157 10.6151
R1621 B.n161 B.n160 10.6151
R1622 B.n164 B.n161 10.6151
R1623 B.n165 B.n164 10.6151
R1624 B.n168 B.n165 10.6151
R1625 B.n169 B.n168 10.6151
R1626 B.n172 B.n169 10.6151
R1627 B.n173 B.n172 10.6151
R1628 B.n176 B.n173 10.6151
R1629 B.n177 B.n176 10.6151
R1630 B.n180 B.n177 10.6151
R1631 B.n181 B.n180 10.6151
R1632 B.n185 B.n184 10.6151
R1633 B.n188 B.n185 10.6151
R1634 B.n189 B.n188 10.6151
R1635 B.n192 B.n189 10.6151
R1636 B.n193 B.n192 10.6151
R1637 B.n196 B.n193 10.6151
R1638 B.n197 B.n196 10.6151
R1639 B.n200 B.n197 10.6151
R1640 B.n205 B.n202 10.6151
R1641 B.n206 B.n205 10.6151
R1642 B.n209 B.n206 10.6151
R1643 B.n210 B.n209 10.6151
R1644 B.n213 B.n210 10.6151
R1645 B.n214 B.n213 10.6151
R1646 B.n217 B.n214 10.6151
R1647 B.n218 B.n217 10.6151
R1648 B.n221 B.n218 10.6151
R1649 B.n222 B.n221 10.6151
R1650 B.n225 B.n222 10.6151
R1651 B.n226 B.n225 10.6151
R1652 B.n229 B.n226 10.6151
R1653 B.n230 B.n229 10.6151
R1654 B.n233 B.n230 10.6151
R1655 B.n234 B.n233 10.6151
R1656 B.n237 B.n234 10.6151
R1657 B.n238 B.n237 10.6151
R1658 B.n241 B.n238 10.6151
R1659 B.n242 B.n241 10.6151
R1660 B.n245 B.n242 10.6151
R1661 B.n246 B.n245 10.6151
R1662 B.n249 B.n246 10.6151
R1663 B.n250 B.n249 10.6151
R1664 B.n253 B.n250 10.6151
R1665 B.n254 B.n253 10.6151
R1666 B.n257 B.n254 10.6151
R1667 B.n258 B.n257 10.6151
R1668 B.n261 B.n258 10.6151
R1669 B.n262 B.n261 10.6151
R1670 B.n265 B.n262 10.6151
R1671 B.n266 B.n265 10.6151
R1672 B.n269 B.n266 10.6151
R1673 B.n270 B.n269 10.6151
R1674 B.n273 B.n270 10.6151
R1675 B.n274 B.n273 10.6151
R1676 B.n277 B.n274 10.6151
R1677 B.n278 B.n277 10.6151
R1678 B.n281 B.n278 10.6151
R1679 B.n282 B.n281 10.6151
R1680 B.n285 B.n282 10.6151
R1681 B.n286 B.n285 10.6151
R1682 B.n289 B.n286 10.6151
R1683 B.n290 B.n289 10.6151
R1684 B.n293 B.n290 10.6151
R1685 B.n294 B.n293 10.6151
R1686 B.n655 B.n294 10.6151
R1687 B.n597 B.n319 10.6151
R1688 B.n598 B.n597 10.6151
R1689 B.n599 B.n598 10.6151
R1690 B.n599 B.n311 10.6151
R1691 B.n609 B.n311 10.6151
R1692 B.n610 B.n609 10.6151
R1693 B.n611 B.n610 10.6151
R1694 B.n611 B.n303 10.6151
R1695 B.n621 B.n303 10.6151
R1696 B.n622 B.n621 10.6151
R1697 B.n624 B.n622 10.6151
R1698 B.n624 B.n623 10.6151
R1699 B.n623 B.n295 10.6151
R1700 B.n635 B.n295 10.6151
R1701 B.n636 B.n635 10.6151
R1702 B.n637 B.n636 10.6151
R1703 B.n638 B.n637 10.6151
R1704 B.n640 B.n638 10.6151
R1705 B.n641 B.n640 10.6151
R1706 B.n642 B.n641 10.6151
R1707 B.n643 B.n642 10.6151
R1708 B.n645 B.n643 10.6151
R1709 B.n646 B.n645 10.6151
R1710 B.n647 B.n646 10.6151
R1711 B.n648 B.n647 10.6151
R1712 B.n650 B.n648 10.6151
R1713 B.n651 B.n650 10.6151
R1714 B.n652 B.n651 10.6151
R1715 B.n653 B.n652 10.6151
R1716 B.n654 B.n653 10.6151
R1717 B.n591 B.n323 10.6151
R1718 B.n586 B.n323 10.6151
R1719 B.n586 B.n585 10.6151
R1720 B.n585 B.n584 10.6151
R1721 B.n584 B.n581 10.6151
R1722 B.n581 B.n580 10.6151
R1723 B.n580 B.n577 10.6151
R1724 B.n577 B.n576 10.6151
R1725 B.n576 B.n573 10.6151
R1726 B.n573 B.n572 10.6151
R1727 B.n572 B.n569 10.6151
R1728 B.n569 B.n568 10.6151
R1729 B.n568 B.n565 10.6151
R1730 B.n565 B.n564 10.6151
R1731 B.n564 B.n561 10.6151
R1732 B.n561 B.n560 10.6151
R1733 B.n560 B.n557 10.6151
R1734 B.n557 B.n556 10.6151
R1735 B.n556 B.n553 10.6151
R1736 B.n553 B.n552 10.6151
R1737 B.n552 B.n549 10.6151
R1738 B.n549 B.n548 10.6151
R1739 B.n548 B.n545 10.6151
R1740 B.n545 B.n544 10.6151
R1741 B.n544 B.n541 10.6151
R1742 B.n541 B.n540 10.6151
R1743 B.n540 B.n537 10.6151
R1744 B.n537 B.n536 10.6151
R1745 B.n536 B.n533 10.6151
R1746 B.n533 B.n532 10.6151
R1747 B.n532 B.n529 10.6151
R1748 B.n529 B.n528 10.6151
R1749 B.n528 B.n525 10.6151
R1750 B.n525 B.n524 10.6151
R1751 B.n524 B.n521 10.6151
R1752 B.n521 B.n520 10.6151
R1753 B.n520 B.n517 10.6151
R1754 B.n517 B.n516 10.6151
R1755 B.n516 B.n513 10.6151
R1756 B.n513 B.n512 10.6151
R1757 B.n512 B.n509 10.6151
R1758 B.n509 B.n508 10.6151
R1759 B.n508 B.n505 10.6151
R1760 B.n505 B.n504 10.6151
R1761 B.n504 B.n501 10.6151
R1762 B.n501 B.n500 10.6151
R1763 B.n500 B.n497 10.6151
R1764 B.n495 B.n492 10.6151
R1765 B.n492 B.n491 10.6151
R1766 B.n491 B.n488 10.6151
R1767 B.n488 B.n487 10.6151
R1768 B.n487 B.n484 10.6151
R1769 B.n484 B.n483 10.6151
R1770 B.n483 B.n480 10.6151
R1771 B.n480 B.n479 10.6151
R1772 B.n476 B.n475 10.6151
R1773 B.n475 B.n472 10.6151
R1774 B.n472 B.n471 10.6151
R1775 B.n471 B.n468 10.6151
R1776 B.n468 B.n467 10.6151
R1777 B.n467 B.n464 10.6151
R1778 B.n464 B.n463 10.6151
R1779 B.n463 B.n460 10.6151
R1780 B.n460 B.n459 10.6151
R1781 B.n459 B.n456 10.6151
R1782 B.n456 B.n455 10.6151
R1783 B.n455 B.n452 10.6151
R1784 B.n452 B.n451 10.6151
R1785 B.n451 B.n448 10.6151
R1786 B.n448 B.n447 10.6151
R1787 B.n447 B.n444 10.6151
R1788 B.n444 B.n443 10.6151
R1789 B.n443 B.n440 10.6151
R1790 B.n440 B.n439 10.6151
R1791 B.n439 B.n436 10.6151
R1792 B.n436 B.n435 10.6151
R1793 B.n435 B.n432 10.6151
R1794 B.n432 B.n431 10.6151
R1795 B.n431 B.n428 10.6151
R1796 B.n428 B.n427 10.6151
R1797 B.n427 B.n424 10.6151
R1798 B.n424 B.n423 10.6151
R1799 B.n423 B.n420 10.6151
R1800 B.n420 B.n419 10.6151
R1801 B.n419 B.n416 10.6151
R1802 B.n416 B.n415 10.6151
R1803 B.n415 B.n412 10.6151
R1804 B.n412 B.n411 10.6151
R1805 B.n411 B.n408 10.6151
R1806 B.n408 B.n407 10.6151
R1807 B.n407 B.n404 10.6151
R1808 B.n404 B.n403 10.6151
R1809 B.n403 B.n400 10.6151
R1810 B.n400 B.n399 10.6151
R1811 B.n399 B.n396 10.6151
R1812 B.n396 B.n395 10.6151
R1813 B.n395 B.n392 10.6151
R1814 B.n392 B.n391 10.6151
R1815 B.n391 B.n388 10.6151
R1816 B.n388 B.n387 10.6151
R1817 B.n387 B.n384 10.6151
R1818 B.n384 B.n383 10.6151
R1819 B.n593 B.n592 10.6151
R1820 B.n593 B.n315 10.6151
R1821 B.n603 B.n315 10.6151
R1822 B.n604 B.n603 10.6151
R1823 B.n605 B.n604 10.6151
R1824 B.n605 B.n307 10.6151
R1825 B.n615 B.n307 10.6151
R1826 B.n616 B.n615 10.6151
R1827 B.n617 B.n616 10.6151
R1828 B.n617 B.n299 10.6151
R1829 B.n628 B.n299 10.6151
R1830 B.n629 B.n628 10.6151
R1831 B.n630 B.n629 10.6151
R1832 B.n630 B.n0 10.6151
R1833 B.n686 B.n1 10.6151
R1834 B.n686 B.n685 10.6151
R1835 B.n685 B.n684 10.6151
R1836 B.n684 B.n10 10.6151
R1837 B.n678 B.n10 10.6151
R1838 B.n678 B.n677 10.6151
R1839 B.n677 B.n676 10.6151
R1840 B.n676 B.n17 10.6151
R1841 B.n670 B.n17 10.6151
R1842 B.n670 B.n669 10.6151
R1843 B.n669 B.n668 10.6151
R1844 B.n668 B.n24 10.6151
R1845 B.n662 B.n24 10.6151
R1846 B.n662 B.n661 10.6151
R1847 B.n184 B.n90 7.18099
R1848 B.n201 B.n200 7.18099
R1849 B.n496 B.n495 7.18099
R1850 B.n479 B.n381 7.18099
R1851 B.n181 B.n90 3.43465
R1852 B.n202 B.n201 3.43465
R1853 B.n497 B.n496 3.43465
R1854 B.n476 B.n381 3.43465
R1855 B.n607 B.t10 2.84655
R1856 B.t3 B.n672 2.84655
R1857 B.n692 B.n0 2.81026
R1858 B.n692 B.n1 2.81026
R1859 VP.n0 VP.t1 657.812
R1860 VP.n0 VP.t0 616.297
R1861 VP VP.n0 0.0516364
R1862 VDD1.n72 VDD1.n0 289.615
R1863 VDD1.n149 VDD1.n77 289.615
R1864 VDD1.n73 VDD1.n72 185
R1865 VDD1.n71 VDD1.n2 185
R1866 VDD1.n70 VDD1.n69 185
R1867 VDD1.n5 VDD1.n3 185
R1868 VDD1.n64 VDD1.n63 185
R1869 VDD1.n62 VDD1.n61 185
R1870 VDD1.n9 VDD1.n8 185
R1871 VDD1.n56 VDD1.n55 185
R1872 VDD1.n54 VDD1.n53 185
R1873 VDD1.n13 VDD1.n12 185
R1874 VDD1.n48 VDD1.n47 185
R1875 VDD1.n46 VDD1.n45 185
R1876 VDD1.n17 VDD1.n16 185
R1877 VDD1.n40 VDD1.n39 185
R1878 VDD1.n38 VDD1.n37 185
R1879 VDD1.n21 VDD1.n20 185
R1880 VDD1.n32 VDD1.n31 185
R1881 VDD1.n30 VDD1.n29 185
R1882 VDD1.n25 VDD1.n24 185
R1883 VDD1.n101 VDD1.n100 185
R1884 VDD1.n106 VDD1.n105 185
R1885 VDD1.n108 VDD1.n107 185
R1886 VDD1.n97 VDD1.n96 185
R1887 VDD1.n114 VDD1.n113 185
R1888 VDD1.n116 VDD1.n115 185
R1889 VDD1.n93 VDD1.n92 185
R1890 VDD1.n122 VDD1.n121 185
R1891 VDD1.n124 VDD1.n123 185
R1892 VDD1.n89 VDD1.n88 185
R1893 VDD1.n130 VDD1.n129 185
R1894 VDD1.n132 VDD1.n131 185
R1895 VDD1.n85 VDD1.n84 185
R1896 VDD1.n138 VDD1.n137 185
R1897 VDD1.n140 VDD1.n139 185
R1898 VDD1.n81 VDD1.n80 185
R1899 VDD1.n147 VDD1.n146 185
R1900 VDD1.n148 VDD1.n79 185
R1901 VDD1.n150 VDD1.n149 185
R1902 VDD1.n26 VDD1.t0 147.659
R1903 VDD1.n102 VDD1.t1 147.659
R1904 VDD1.n72 VDD1.n71 104.615
R1905 VDD1.n71 VDD1.n70 104.615
R1906 VDD1.n70 VDD1.n3 104.615
R1907 VDD1.n63 VDD1.n3 104.615
R1908 VDD1.n63 VDD1.n62 104.615
R1909 VDD1.n62 VDD1.n8 104.615
R1910 VDD1.n55 VDD1.n8 104.615
R1911 VDD1.n55 VDD1.n54 104.615
R1912 VDD1.n54 VDD1.n12 104.615
R1913 VDD1.n47 VDD1.n12 104.615
R1914 VDD1.n47 VDD1.n46 104.615
R1915 VDD1.n46 VDD1.n16 104.615
R1916 VDD1.n39 VDD1.n16 104.615
R1917 VDD1.n39 VDD1.n38 104.615
R1918 VDD1.n38 VDD1.n20 104.615
R1919 VDD1.n31 VDD1.n20 104.615
R1920 VDD1.n31 VDD1.n30 104.615
R1921 VDD1.n30 VDD1.n24 104.615
R1922 VDD1.n106 VDD1.n100 104.615
R1923 VDD1.n107 VDD1.n106 104.615
R1924 VDD1.n107 VDD1.n96 104.615
R1925 VDD1.n114 VDD1.n96 104.615
R1926 VDD1.n115 VDD1.n114 104.615
R1927 VDD1.n115 VDD1.n92 104.615
R1928 VDD1.n122 VDD1.n92 104.615
R1929 VDD1.n123 VDD1.n122 104.615
R1930 VDD1.n123 VDD1.n88 104.615
R1931 VDD1.n130 VDD1.n88 104.615
R1932 VDD1.n131 VDD1.n130 104.615
R1933 VDD1.n131 VDD1.n84 104.615
R1934 VDD1.n138 VDD1.n84 104.615
R1935 VDD1.n139 VDD1.n138 104.615
R1936 VDD1.n139 VDD1.n80 104.615
R1937 VDD1.n147 VDD1.n80 104.615
R1938 VDD1.n148 VDD1.n147 104.615
R1939 VDD1.n149 VDD1.n148 104.615
R1940 VDD1 VDD1.n153 89.5438
R1941 VDD1.t0 VDD1.n24 52.3082
R1942 VDD1.t1 VDD1.n100 52.3082
R1943 VDD1 VDD1.n76 51.3057
R1944 VDD1.n26 VDD1.n25 15.6677
R1945 VDD1.n102 VDD1.n101 15.6677
R1946 VDD1.n73 VDD1.n2 13.1884
R1947 VDD1.n150 VDD1.n79 13.1884
R1948 VDD1.n74 VDD1.n0 12.8005
R1949 VDD1.n69 VDD1.n4 12.8005
R1950 VDD1.n29 VDD1.n28 12.8005
R1951 VDD1.n105 VDD1.n104 12.8005
R1952 VDD1.n146 VDD1.n145 12.8005
R1953 VDD1.n151 VDD1.n77 12.8005
R1954 VDD1.n68 VDD1.n5 12.0247
R1955 VDD1.n32 VDD1.n23 12.0247
R1956 VDD1.n108 VDD1.n99 12.0247
R1957 VDD1.n144 VDD1.n81 12.0247
R1958 VDD1.n65 VDD1.n64 11.249
R1959 VDD1.n33 VDD1.n21 11.249
R1960 VDD1.n109 VDD1.n97 11.249
R1961 VDD1.n141 VDD1.n140 11.249
R1962 VDD1.n61 VDD1.n7 10.4732
R1963 VDD1.n37 VDD1.n36 10.4732
R1964 VDD1.n113 VDD1.n112 10.4732
R1965 VDD1.n137 VDD1.n83 10.4732
R1966 VDD1.n60 VDD1.n9 9.69747
R1967 VDD1.n40 VDD1.n19 9.69747
R1968 VDD1.n116 VDD1.n95 9.69747
R1969 VDD1.n136 VDD1.n85 9.69747
R1970 VDD1.n76 VDD1.n75 9.45567
R1971 VDD1.n153 VDD1.n152 9.45567
R1972 VDD1.n52 VDD1.n51 9.3005
R1973 VDD1.n11 VDD1.n10 9.3005
R1974 VDD1.n58 VDD1.n57 9.3005
R1975 VDD1.n60 VDD1.n59 9.3005
R1976 VDD1.n7 VDD1.n6 9.3005
R1977 VDD1.n66 VDD1.n65 9.3005
R1978 VDD1.n68 VDD1.n67 9.3005
R1979 VDD1.n4 VDD1.n1 9.3005
R1980 VDD1.n75 VDD1.n74 9.3005
R1981 VDD1.n50 VDD1.n49 9.3005
R1982 VDD1.n15 VDD1.n14 9.3005
R1983 VDD1.n44 VDD1.n43 9.3005
R1984 VDD1.n42 VDD1.n41 9.3005
R1985 VDD1.n19 VDD1.n18 9.3005
R1986 VDD1.n36 VDD1.n35 9.3005
R1987 VDD1.n34 VDD1.n33 9.3005
R1988 VDD1.n23 VDD1.n22 9.3005
R1989 VDD1.n28 VDD1.n27 9.3005
R1990 VDD1.n152 VDD1.n151 9.3005
R1991 VDD1.n91 VDD1.n90 9.3005
R1992 VDD1.n120 VDD1.n119 9.3005
R1993 VDD1.n118 VDD1.n117 9.3005
R1994 VDD1.n95 VDD1.n94 9.3005
R1995 VDD1.n112 VDD1.n111 9.3005
R1996 VDD1.n110 VDD1.n109 9.3005
R1997 VDD1.n99 VDD1.n98 9.3005
R1998 VDD1.n104 VDD1.n103 9.3005
R1999 VDD1.n126 VDD1.n125 9.3005
R2000 VDD1.n128 VDD1.n127 9.3005
R2001 VDD1.n87 VDD1.n86 9.3005
R2002 VDD1.n134 VDD1.n133 9.3005
R2003 VDD1.n136 VDD1.n135 9.3005
R2004 VDD1.n83 VDD1.n82 9.3005
R2005 VDD1.n142 VDD1.n141 9.3005
R2006 VDD1.n144 VDD1.n143 9.3005
R2007 VDD1.n145 VDD1.n78 9.3005
R2008 VDD1.n57 VDD1.n56 8.92171
R2009 VDD1.n41 VDD1.n17 8.92171
R2010 VDD1.n117 VDD1.n93 8.92171
R2011 VDD1.n133 VDD1.n132 8.92171
R2012 VDD1.n53 VDD1.n11 8.14595
R2013 VDD1.n45 VDD1.n44 8.14595
R2014 VDD1.n121 VDD1.n120 8.14595
R2015 VDD1.n129 VDD1.n87 8.14595
R2016 VDD1.n52 VDD1.n13 7.3702
R2017 VDD1.n48 VDD1.n15 7.3702
R2018 VDD1.n124 VDD1.n91 7.3702
R2019 VDD1.n128 VDD1.n89 7.3702
R2020 VDD1.n49 VDD1.n13 6.59444
R2021 VDD1.n49 VDD1.n48 6.59444
R2022 VDD1.n125 VDD1.n124 6.59444
R2023 VDD1.n125 VDD1.n89 6.59444
R2024 VDD1.n53 VDD1.n52 5.81868
R2025 VDD1.n45 VDD1.n15 5.81868
R2026 VDD1.n121 VDD1.n91 5.81868
R2027 VDD1.n129 VDD1.n128 5.81868
R2028 VDD1.n56 VDD1.n11 5.04292
R2029 VDD1.n44 VDD1.n17 5.04292
R2030 VDD1.n120 VDD1.n93 5.04292
R2031 VDD1.n132 VDD1.n87 5.04292
R2032 VDD1.n27 VDD1.n26 4.38563
R2033 VDD1.n103 VDD1.n102 4.38563
R2034 VDD1.n57 VDD1.n9 4.26717
R2035 VDD1.n41 VDD1.n40 4.26717
R2036 VDD1.n117 VDD1.n116 4.26717
R2037 VDD1.n133 VDD1.n85 4.26717
R2038 VDD1.n61 VDD1.n60 3.49141
R2039 VDD1.n37 VDD1.n19 3.49141
R2040 VDD1.n113 VDD1.n95 3.49141
R2041 VDD1.n137 VDD1.n136 3.49141
R2042 VDD1.n64 VDD1.n7 2.71565
R2043 VDD1.n36 VDD1.n21 2.71565
R2044 VDD1.n112 VDD1.n97 2.71565
R2045 VDD1.n140 VDD1.n83 2.71565
R2046 VDD1.n65 VDD1.n5 1.93989
R2047 VDD1.n33 VDD1.n32 1.93989
R2048 VDD1.n109 VDD1.n108 1.93989
R2049 VDD1.n141 VDD1.n81 1.93989
R2050 VDD1.n76 VDD1.n0 1.16414
R2051 VDD1.n69 VDD1.n68 1.16414
R2052 VDD1.n29 VDD1.n23 1.16414
R2053 VDD1.n105 VDD1.n99 1.16414
R2054 VDD1.n146 VDD1.n144 1.16414
R2055 VDD1.n153 VDD1.n77 1.16414
R2056 VDD1.n74 VDD1.n73 0.388379
R2057 VDD1.n4 VDD1.n2 0.388379
R2058 VDD1.n28 VDD1.n25 0.388379
R2059 VDD1.n104 VDD1.n101 0.388379
R2060 VDD1.n145 VDD1.n79 0.388379
R2061 VDD1.n151 VDD1.n150 0.388379
R2062 VDD1.n75 VDD1.n1 0.155672
R2063 VDD1.n67 VDD1.n1 0.155672
R2064 VDD1.n67 VDD1.n66 0.155672
R2065 VDD1.n66 VDD1.n6 0.155672
R2066 VDD1.n59 VDD1.n6 0.155672
R2067 VDD1.n59 VDD1.n58 0.155672
R2068 VDD1.n58 VDD1.n10 0.155672
R2069 VDD1.n51 VDD1.n10 0.155672
R2070 VDD1.n51 VDD1.n50 0.155672
R2071 VDD1.n50 VDD1.n14 0.155672
R2072 VDD1.n43 VDD1.n14 0.155672
R2073 VDD1.n43 VDD1.n42 0.155672
R2074 VDD1.n42 VDD1.n18 0.155672
R2075 VDD1.n35 VDD1.n18 0.155672
R2076 VDD1.n35 VDD1.n34 0.155672
R2077 VDD1.n34 VDD1.n22 0.155672
R2078 VDD1.n27 VDD1.n22 0.155672
R2079 VDD1.n103 VDD1.n98 0.155672
R2080 VDD1.n110 VDD1.n98 0.155672
R2081 VDD1.n111 VDD1.n110 0.155672
R2082 VDD1.n111 VDD1.n94 0.155672
R2083 VDD1.n118 VDD1.n94 0.155672
R2084 VDD1.n119 VDD1.n118 0.155672
R2085 VDD1.n119 VDD1.n90 0.155672
R2086 VDD1.n126 VDD1.n90 0.155672
R2087 VDD1.n127 VDD1.n126 0.155672
R2088 VDD1.n127 VDD1.n86 0.155672
R2089 VDD1.n134 VDD1.n86 0.155672
R2090 VDD1.n135 VDD1.n134 0.155672
R2091 VDD1.n135 VDD1.n82 0.155672
R2092 VDD1.n142 VDD1.n82 0.155672
R2093 VDD1.n143 VDD1.n142 0.155672
R2094 VDD1.n143 VDD1.n78 0.155672
R2095 VDD1.n152 VDD1.n78 0.155672
C0 VTAIL VP 1.86147f
C1 VDD1 VP 2.52974f
C2 VDD2 VP 0.260692f
C3 VN VP 4.99642f
C4 VTAIL VDD1 6.17953f
C5 VTAIL VDD2 6.21369f
C6 VDD1 VDD2 0.475358f
C7 VTAIL VN 1.84682f
C8 VDD1 VN 0.148648f
C9 VN VDD2 2.4225f
C10 VDD2 B 4.168831f
C11 VDD1 B 6.77415f
C12 VTAIL B 7.220294f
C13 VN B 8.589311f
C14 VP B 4.323363f
C15 VDD1.n0 B 0.027165f
C16 VDD1.n1 B 0.020613f
C17 VDD1.n2 B 0.011402f
C18 VDD1.n3 B 0.026181f
C19 VDD1.n4 B 0.011076f
C20 VDD1.n5 B 0.011728f
C21 VDD1.n6 B 0.020613f
C22 VDD1.n7 B 0.011076f
C23 VDD1.n8 B 0.026181f
C24 VDD1.n9 B 0.011728f
C25 VDD1.n10 B 0.020613f
C26 VDD1.n11 B 0.011076f
C27 VDD1.n12 B 0.026181f
C28 VDD1.n13 B 0.011728f
C29 VDD1.n14 B 0.020613f
C30 VDD1.n15 B 0.011076f
C31 VDD1.n16 B 0.026181f
C32 VDD1.n17 B 0.011728f
C33 VDD1.n18 B 0.020613f
C34 VDD1.n19 B 0.011076f
C35 VDD1.n20 B 0.026181f
C36 VDD1.n21 B 0.011728f
C37 VDD1.n22 B 0.020613f
C38 VDD1.n23 B 0.011076f
C39 VDD1.n24 B 0.019635f
C40 VDD1.n25 B 0.015466f
C41 VDD1.t0 B 0.0431f
C42 VDD1.n26 B 0.129428f
C43 VDD1.n27 B 1.24946f
C44 VDD1.n28 B 0.011076f
C45 VDD1.n29 B 0.011728f
C46 VDD1.n30 B 0.026181f
C47 VDD1.n31 B 0.026181f
C48 VDD1.n32 B 0.011728f
C49 VDD1.n33 B 0.011076f
C50 VDD1.n34 B 0.020613f
C51 VDD1.n35 B 0.020613f
C52 VDD1.n36 B 0.011076f
C53 VDD1.n37 B 0.011728f
C54 VDD1.n38 B 0.026181f
C55 VDD1.n39 B 0.026181f
C56 VDD1.n40 B 0.011728f
C57 VDD1.n41 B 0.011076f
C58 VDD1.n42 B 0.020613f
C59 VDD1.n43 B 0.020613f
C60 VDD1.n44 B 0.011076f
C61 VDD1.n45 B 0.011728f
C62 VDD1.n46 B 0.026181f
C63 VDD1.n47 B 0.026181f
C64 VDD1.n48 B 0.011728f
C65 VDD1.n49 B 0.011076f
C66 VDD1.n50 B 0.020613f
C67 VDD1.n51 B 0.020613f
C68 VDD1.n52 B 0.011076f
C69 VDD1.n53 B 0.011728f
C70 VDD1.n54 B 0.026181f
C71 VDD1.n55 B 0.026181f
C72 VDD1.n56 B 0.011728f
C73 VDD1.n57 B 0.011076f
C74 VDD1.n58 B 0.020613f
C75 VDD1.n59 B 0.020613f
C76 VDD1.n60 B 0.011076f
C77 VDD1.n61 B 0.011728f
C78 VDD1.n62 B 0.026181f
C79 VDD1.n63 B 0.026181f
C80 VDD1.n64 B 0.011728f
C81 VDD1.n65 B 0.011076f
C82 VDD1.n66 B 0.020613f
C83 VDD1.n67 B 0.020613f
C84 VDD1.n68 B 0.011076f
C85 VDD1.n69 B 0.011728f
C86 VDD1.n70 B 0.026181f
C87 VDD1.n71 B 0.026181f
C88 VDD1.n72 B 0.05348f
C89 VDD1.n73 B 0.011402f
C90 VDD1.n74 B 0.011076f
C91 VDD1.n75 B 0.050743f
C92 VDD1.n76 B 0.04427f
C93 VDD1.n77 B 0.027165f
C94 VDD1.n78 B 0.020613f
C95 VDD1.n79 B 0.011402f
C96 VDD1.n80 B 0.026181f
C97 VDD1.n81 B 0.011728f
C98 VDD1.n82 B 0.020613f
C99 VDD1.n83 B 0.011076f
C100 VDD1.n84 B 0.026181f
C101 VDD1.n85 B 0.011728f
C102 VDD1.n86 B 0.020613f
C103 VDD1.n87 B 0.011076f
C104 VDD1.n88 B 0.026181f
C105 VDD1.n89 B 0.011728f
C106 VDD1.n90 B 0.020613f
C107 VDD1.n91 B 0.011076f
C108 VDD1.n92 B 0.026181f
C109 VDD1.n93 B 0.011728f
C110 VDD1.n94 B 0.020613f
C111 VDD1.n95 B 0.011076f
C112 VDD1.n96 B 0.026181f
C113 VDD1.n97 B 0.011728f
C114 VDD1.n98 B 0.020613f
C115 VDD1.n99 B 0.011076f
C116 VDD1.n100 B 0.019635f
C117 VDD1.n101 B 0.015466f
C118 VDD1.t1 B 0.0431f
C119 VDD1.n102 B 0.129428f
C120 VDD1.n103 B 1.24946f
C121 VDD1.n104 B 0.011076f
C122 VDD1.n105 B 0.011728f
C123 VDD1.n106 B 0.026181f
C124 VDD1.n107 B 0.026181f
C125 VDD1.n108 B 0.011728f
C126 VDD1.n109 B 0.011076f
C127 VDD1.n110 B 0.020613f
C128 VDD1.n111 B 0.020613f
C129 VDD1.n112 B 0.011076f
C130 VDD1.n113 B 0.011728f
C131 VDD1.n114 B 0.026181f
C132 VDD1.n115 B 0.026181f
C133 VDD1.n116 B 0.011728f
C134 VDD1.n117 B 0.011076f
C135 VDD1.n118 B 0.020613f
C136 VDD1.n119 B 0.020613f
C137 VDD1.n120 B 0.011076f
C138 VDD1.n121 B 0.011728f
C139 VDD1.n122 B 0.026181f
C140 VDD1.n123 B 0.026181f
C141 VDD1.n124 B 0.011728f
C142 VDD1.n125 B 0.011076f
C143 VDD1.n126 B 0.020613f
C144 VDD1.n127 B 0.020613f
C145 VDD1.n128 B 0.011076f
C146 VDD1.n129 B 0.011728f
C147 VDD1.n130 B 0.026181f
C148 VDD1.n131 B 0.026181f
C149 VDD1.n132 B 0.011728f
C150 VDD1.n133 B 0.011076f
C151 VDD1.n134 B 0.020613f
C152 VDD1.n135 B 0.020613f
C153 VDD1.n136 B 0.011076f
C154 VDD1.n137 B 0.011728f
C155 VDD1.n138 B 0.026181f
C156 VDD1.n139 B 0.026181f
C157 VDD1.n140 B 0.011728f
C158 VDD1.n141 B 0.011076f
C159 VDD1.n142 B 0.020613f
C160 VDD1.n143 B 0.020613f
C161 VDD1.n144 B 0.011076f
C162 VDD1.n145 B 0.011076f
C163 VDD1.n146 B 0.011728f
C164 VDD1.n147 B 0.026181f
C165 VDD1.n148 B 0.026181f
C166 VDD1.n149 B 0.05348f
C167 VDD1.n150 B 0.011402f
C168 VDD1.n151 B 0.011076f
C169 VDD1.n152 B 0.050743f
C170 VDD1.n153 B 0.585325f
C171 VP.t1 B 1.70856f
C172 VP.t0 B 1.57231f
C173 VP.n0 B 4.20065f
C174 VDD2.n0 B 0.02709f
C175 VDD2.n1 B 0.020556f
C176 VDD2.n2 B 0.011371f
C177 VDD2.n3 B 0.026108f
C178 VDD2.n4 B 0.011696f
C179 VDD2.n5 B 0.020556f
C180 VDD2.n6 B 0.011046f
C181 VDD2.n7 B 0.026108f
C182 VDD2.n8 B 0.011696f
C183 VDD2.n9 B 0.020556f
C184 VDD2.n10 B 0.011046f
C185 VDD2.n11 B 0.026108f
C186 VDD2.n12 B 0.011696f
C187 VDD2.n13 B 0.020556f
C188 VDD2.n14 B 0.011046f
C189 VDD2.n15 B 0.026108f
C190 VDD2.n16 B 0.011696f
C191 VDD2.n17 B 0.020556f
C192 VDD2.n18 B 0.011046f
C193 VDD2.n19 B 0.026108f
C194 VDD2.n20 B 0.011696f
C195 VDD2.n21 B 0.020556f
C196 VDD2.n22 B 0.011046f
C197 VDD2.n23 B 0.019581f
C198 VDD2.n24 B 0.015423f
C199 VDD2.t0 B 0.042981f
C200 VDD2.n25 B 0.12907f
C201 VDD2.n26 B 1.246f
C202 VDD2.n27 B 0.011046f
C203 VDD2.n28 B 0.011696f
C204 VDD2.n29 B 0.026108f
C205 VDD2.n30 B 0.026108f
C206 VDD2.n31 B 0.011696f
C207 VDD2.n32 B 0.011046f
C208 VDD2.n33 B 0.020556f
C209 VDD2.n34 B 0.020556f
C210 VDD2.n35 B 0.011046f
C211 VDD2.n36 B 0.011696f
C212 VDD2.n37 B 0.026108f
C213 VDD2.n38 B 0.026108f
C214 VDD2.n39 B 0.011696f
C215 VDD2.n40 B 0.011046f
C216 VDD2.n41 B 0.020556f
C217 VDD2.n42 B 0.020556f
C218 VDD2.n43 B 0.011046f
C219 VDD2.n44 B 0.011696f
C220 VDD2.n45 B 0.026108f
C221 VDD2.n46 B 0.026108f
C222 VDD2.n47 B 0.011696f
C223 VDD2.n48 B 0.011046f
C224 VDD2.n49 B 0.020556f
C225 VDD2.n50 B 0.020556f
C226 VDD2.n51 B 0.011046f
C227 VDD2.n52 B 0.011696f
C228 VDD2.n53 B 0.026108f
C229 VDD2.n54 B 0.026108f
C230 VDD2.n55 B 0.011696f
C231 VDD2.n56 B 0.011046f
C232 VDD2.n57 B 0.020556f
C233 VDD2.n58 B 0.020556f
C234 VDD2.n59 B 0.011046f
C235 VDD2.n60 B 0.011696f
C236 VDD2.n61 B 0.026108f
C237 VDD2.n62 B 0.026108f
C238 VDD2.n63 B 0.011696f
C239 VDD2.n64 B 0.011046f
C240 VDD2.n65 B 0.020556f
C241 VDD2.n66 B 0.020556f
C242 VDD2.n67 B 0.011046f
C243 VDD2.n68 B 0.011046f
C244 VDD2.n69 B 0.011696f
C245 VDD2.n70 B 0.026108f
C246 VDD2.n71 B 0.026108f
C247 VDD2.n72 B 0.053331f
C248 VDD2.n73 B 0.011371f
C249 VDD2.n74 B 0.011046f
C250 VDD2.n75 B 0.050602f
C251 VDD2.n76 B 0.55508f
C252 VDD2.n77 B 0.02709f
C253 VDD2.n78 B 0.020556f
C254 VDD2.n79 B 0.011371f
C255 VDD2.n80 B 0.026108f
C256 VDD2.n81 B 0.011046f
C257 VDD2.n82 B 0.011696f
C258 VDD2.n83 B 0.020556f
C259 VDD2.n84 B 0.011046f
C260 VDD2.n85 B 0.026108f
C261 VDD2.n86 B 0.011696f
C262 VDD2.n87 B 0.020556f
C263 VDD2.n88 B 0.011046f
C264 VDD2.n89 B 0.026108f
C265 VDD2.n90 B 0.011696f
C266 VDD2.n91 B 0.020556f
C267 VDD2.n92 B 0.011046f
C268 VDD2.n93 B 0.026108f
C269 VDD2.n94 B 0.011696f
C270 VDD2.n95 B 0.020556f
C271 VDD2.n96 B 0.011046f
C272 VDD2.n97 B 0.026108f
C273 VDD2.n98 B 0.011696f
C274 VDD2.n99 B 0.020556f
C275 VDD2.n100 B 0.011046f
C276 VDD2.n101 B 0.019581f
C277 VDD2.n102 B 0.015423f
C278 VDD2.t1 B 0.042981f
C279 VDD2.n103 B 0.12907f
C280 VDD2.n104 B 1.246f
C281 VDD2.n105 B 0.011046f
C282 VDD2.n106 B 0.011696f
C283 VDD2.n107 B 0.026108f
C284 VDD2.n108 B 0.026108f
C285 VDD2.n109 B 0.011696f
C286 VDD2.n110 B 0.011046f
C287 VDD2.n111 B 0.020556f
C288 VDD2.n112 B 0.020556f
C289 VDD2.n113 B 0.011046f
C290 VDD2.n114 B 0.011696f
C291 VDD2.n115 B 0.026108f
C292 VDD2.n116 B 0.026108f
C293 VDD2.n117 B 0.011696f
C294 VDD2.n118 B 0.011046f
C295 VDD2.n119 B 0.020556f
C296 VDD2.n120 B 0.020556f
C297 VDD2.n121 B 0.011046f
C298 VDD2.n122 B 0.011696f
C299 VDD2.n123 B 0.026108f
C300 VDD2.n124 B 0.026108f
C301 VDD2.n125 B 0.011696f
C302 VDD2.n126 B 0.011046f
C303 VDD2.n127 B 0.020556f
C304 VDD2.n128 B 0.020556f
C305 VDD2.n129 B 0.011046f
C306 VDD2.n130 B 0.011696f
C307 VDD2.n131 B 0.026108f
C308 VDD2.n132 B 0.026108f
C309 VDD2.n133 B 0.011696f
C310 VDD2.n134 B 0.011046f
C311 VDD2.n135 B 0.020556f
C312 VDD2.n136 B 0.020556f
C313 VDD2.n137 B 0.011046f
C314 VDD2.n138 B 0.011696f
C315 VDD2.n139 B 0.026108f
C316 VDD2.n140 B 0.026108f
C317 VDD2.n141 B 0.011696f
C318 VDD2.n142 B 0.011046f
C319 VDD2.n143 B 0.020556f
C320 VDD2.n144 B 0.020556f
C321 VDD2.n145 B 0.011046f
C322 VDD2.n146 B 0.011696f
C323 VDD2.n147 B 0.026108f
C324 VDD2.n148 B 0.026108f
C325 VDD2.n149 B 0.053331f
C326 VDD2.n150 B 0.011371f
C327 VDD2.n151 B 0.011046f
C328 VDD2.n152 B 0.050602f
C329 VDD2.n153 B 0.043776f
C330 VDD2.n154 B 2.41603f
C331 VTAIL.n0 B 0.020687f
C332 VTAIL.n1 B 0.015697f
C333 VTAIL.n2 B 0.008683f
C334 VTAIL.n3 B 0.019937f
C335 VTAIL.n4 B 0.008931f
C336 VTAIL.n5 B 0.015697f
C337 VTAIL.n6 B 0.008435f
C338 VTAIL.n7 B 0.019937f
C339 VTAIL.n8 B 0.008931f
C340 VTAIL.n9 B 0.015697f
C341 VTAIL.n10 B 0.008435f
C342 VTAIL.n11 B 0.019937f
C343 VTAIL.n12 B 0.008931f
C344 VTAIL.n13 B 0.015697f
C345 VTAIL.n14 B 0.008435f
C346 VTAIL.n15 B 0.019937f
C347 VTAIL.n16 B 0.008931f
C348 VTAIL.n17 B 0.015697f
C349 VTAIL.n18 B 0.008435f
C350 VTAIL.n19 B 0.019937f
C351 VTAIL.n20 B 0.008931f
C352 VTAIL.n21 B 0.015697f
C353 VTAIL.n22 B 0.008435f
C354 VTAIL.n23 B 0.014953f
C355 VTAIL.n24 B 0.011778f
C356 VTAIL.t1 B 0.032822f
C357 VTAIL.n25 B 0.098563f
C358 VTAIL.n26 B 0.951506f
C359 VTAIL.n27 B 0.008435f
C360 VTAIL.n28 B 0.008931f
C361 VTAIL.n29 B 0.019937f
C362 VTAIL.n30 B 0.019937f
C363 VTAIL.n31 B 0.008931f
C364 VTAIL.n32 B 0.008435f
C365 VTAIL.n33 B 0.015697f
C366 VTAIL.n34 B 0.015697f
C367 VTAIL.n35 B 0.008435f
C368 VTAIL.n36 B 0.008931f
C369 VTAIL.n37 B 0.019937f
C370 VTAIL.n38 B 0.019937f
C371 VTAIL.n39 B 0.008931f
C372 VTAIL.n40 B 0.008435f
C373 VTAIL.n41 B 0.015697f
C374 VTAIL.n42 B 0.015697f
C375 VTAIL.n43 B 0.008435f
C376 VTAIL.n44 B 0.008931f
C377 VTAIL.n45 B 0.019937f
C378 VTAIL.n46 B 0.019937f
C379 VTAIL.n47 B 0.008931f
C380 VTAIL.n48 B 0.008435f
C381 VTAIL.n49 B 0.015697f
C382 VTAIL.n50 B 0.015697f
C383 VTAIL.n51 B 0.008435f
C384 VTAIL.n52 B 0.008931f
C385 VTAIL.n53 B 0.019937f
C386 VTAIL.n54 B 0.019937f
C387 VTAIL.n55 B 0.008931f
C388 VTAIL.n56 B 0.008435f
C389 VTAIL.n57 B 0.015697f
C390 VTAIL.n58 B 0.015697f
C391 VTAIL.n59 B 0.008435f
C392 VTAIL.n60 B 0.008931f
C393 VTAIL.n61 B 0.019937f
C394 VTAIL.n62 B 0.019937f
C395 VTAIL.n63 B 0.008931f
C396 VTAIL.n64 B 0.008435f
C397 VTAIL.n65 B 0.015697f
C398 VTAIL.n66 B 0.015697f
C399 VTAIL.n67 B 0.008435f
C400 VTAIL.n68 B 0.008435f
C401 VTAIL.n69 B 0.008931f
C402 VTAIL.n70 B 0.019937f
C403 VTAIL.n71 B 0.019937f
C404 VTAIL.n72 B 0.040726f
C405 VTAIL.n73 B 0.008683f
C406 VTAIL.n74 B 0.008435f
C407 VTAIL.n75 B 0.038642f
C408 VTAIL.n76 B 0.022608f
C409 VTAIL.n77 B 0.981113f
C410 VTAIL.n78 B 0.020687f
C411 VTAIL.n79 B 0.015697f
C412 VTAIL.n80 B 0.008683f
C413 VTAIL.n81 B 0.019937f
C414 VTAIL.n82 B 0.008435f
C415 VTAIL.n83 B 0.008931f
C416 VTAIL.n84 B 0.015697f
C417 VTAIL.n85 B 0.008435f
C418 VTAIL.n86 B 0.019937f
C419 VTAIL.n87 B 0.008931f
C420 VTAIL.n88 B 0.015697f
C421 VTAIL.n89 B 0.008435f
C422 VTAIL.n90 B 0.019937f
C423 VTAIL.n91 B 0.008931f
C424 VTAIL.n92 B 0.015697f
C425 VTAIL.n93 B 0.008435f
C426 VTAIL.n94 B 0.019937f
C427 VTAIL.n95 B 0.008931f
C428 VTAIL.n96 B 0.015697f
C429 VTAIL.n97 B 0.008435f
C430 VTAIL.n98 B 0.019937f
C431 VTAIL.n99 B 0.008931f
C432 VTAIL.n100 B 0.015697f
C433 VTAIL.n101 B 0.008435f
C434 VTAIL.n102 B 0.014953f
C435 VTAIL.n103 B 0.011778f
C436 VTAIL.t2 B 0.032822f
C437 VTAIL.n104 B 0.098563f
C438 VTAIL.n105 B 0.951506f
C439 VTAIL.n106 B 0.008435f
C440 VTAIL.n107 B 0.008931f
C441 VTAIL.n108 B 0.019937f
C442 VTAIL.n109 B 0.019937f
C443 VTAIL.n110 B 0.008931f
C444 VTAIL.n111 B 0.008435f
C445 VTAIL.n112 B 0.015697f
C446 VTAIL.n113 B 0.015697f
C447 VTAIL.n114 B 0.008435f
C448 VTAIL.n115 B 0.008931f
C449 VTAIL.n116 B 0.019937f
C450 VTAIL.n117 B 0.019937f
C451 VTAIL.n118 B 0.008931f
C452 VTAIL.n119 B 0.008435f
C453 VTAIL.n120 B 0.015697f
C454 VTAIL.n121 B 0.015697f
C455 VTAIL.n122 B 0.008435f
C456 VTAIL.n123 B 0.008931f
C457 VTAIL.n124 B 0.019937f
C458 VTAIL.n125 B 0.019937f
C459 VTAIL.n126 B 0.008931f
C460 VTAIL.n127 B 0.008435f
C461 VTAIL.n128 B 0.015697f
C462 VTAIL.n129 B 0.015697f
C463 VTAIL.n130 B 0.008435f
C464 VTAIL.n131 B 0.008931f
C465 VTAIL.n132 B 0.019937f
C466 VTAIL.n133 B 0.019937f
C467 VTAIL.n134 B 0.008931f
C468 VTAIL.n135 B 0.008435f
C469 VTAIL.n136 B 0.015697f
C470 VTAIL.n137 B 0.015697f
C471 VTAIL.n138 B 0.008435f
C472 VTAIL.n139 B 0.008931f
C473 VTAIL.n140 B 0.019937f
C474 VTAIL.n141 B 0.019937f
C475 VTAIL.n142 B 0.008931f
C476 VTAIL.n143 B 0.008435f
C477 VTAIL.n144 B 0.015697f
C478 VTAIL.n145 B 0.015697f
C479 VTAIL.n146 B 0.008435f
C480 VTAIL.n147 B 0.008931f
C481 VTAIL.n148 B 0.019937f
C482 VTAIL.n149 B 0.019937f
C483 VTAIL.n150 B 0.040726f
C484 VTAIL.n151 B 0.008683f
C485 VTAIL.n152 B 0.008435f
C486 VTAIL.n153 B 0.038642f
C487 VTAIL.n154 B 0.022608f
C488 VTAIL.n155 B 0.990815f
C489 VTAIL.n156 B 0.020687f
C490 VTAIL.n157 B 0.015697f
C491 VTAIL.n158 B 0.008683f
C492 VTAIL.n159 B 0.019937f
C493 VTAIL.n160 B 0.008435f
C494 VTAIL.n161 B 0.008931f
C495 VTAIL.n162 B 0.015697f
C496 VTAIL.n163 B 0.008435f
C497 VTAIL.n164 B 0.019937f
C498 VTAIL.n165 B 0.008931f
C499 VTAIL.n166 B 0.015697f
C500 VTAIL.n167 B 0.008435f
C501 VTAIL.n168 B 0.019937f
C502 VTAIL.n169 B 0.008931f
C503 VTAIL.n170 B 0.015697f
C504 VTAIL.n171 B 0.008435f
C505 VTAIL.n172 B 0.019937f
C506 VTAIL.n173 B 0.008931f
C507 VTAIL.n174 B 0.015697f
C508 VTAIL.n175 B 0.008435f
C509 VTAIL.n176 B 0.019937f
C510 VTAIL.n177 B 0.008931f
C511 VTAIL.n178 B 0.015697f
C512 VTAIL.n179 B 0.008435f
C513 VTAIL.n180 B 0.014953f
C514 VTAIL.n181 B 0.011778f
C515 VTAIL.t0 B 0.032822f
C516 VTAIL.n182 B 0.098563f
C517 VTAIL.n183 B 0.951506f
C518 VTAIL.n184 B 0.008435f
C519 VTAIL.n185 B 0.008931f
C520 VTAIL.n186 B 0.019937f
C521 VTAIL.n187 B 0.019937f
C522 VTAIL.n188 B 0.008931f
C523 VTAIL.n189 B 0.008435f
C524 VTAIL.n190 B 0.015697f
C525 VTAIL.n191 B 0.015697f
C526 VTAIL.n192 B 0.008435f
C527 VTAIL.n193 B 0.008931f
C528 VTAIL.n194 B 0.019937f
C529 VTAIL.n195 B 0.019937f
C530 VTAIL.n196 B 0.008931f
C531 VTAIL.n197 B 0.008435f
C532 VTAIL.n198 B 0.015697f
C533 VTAIL.n199 B 0.015697f
C534 VTAIL.n200 B 0.008435f
C535 VTAIL.n201 B 0.008931f
C536 VTAIL.n202 B 0.019937f
C537 VTAIL.n203 B 0.019937f
C538 VTAIL.n204 B 0.008931f
C539 VTAIL.n205 B 0.008435f
C540 VTAIL.n206 B 0.015697f
C541 VTAIL.n207 B 0.015697f
C542 VTAIL.n208 B 0.008435f
C543 VTAIL.n209 B 0.008931f
C544 VTAIL.n210 B 0.019937f
C545 VTAIL.n211 B 0.019937f
C546 VTAIL.n212 B 0.008931f
C547 VTAIL.n213 B 0.008435f
C548 VTAIL.n214 B 0.015697f
C549 VTAIL.n215 B 0.015697f
C550 VTAIL.n216 B 0.008435f
C551 VTAIL.n217 B 0.008931f
C552 VTAIL.n218 B 0.019937f
C553 VTAIL.n219 B 0.019937f
C554 VTAIL.n220 B 0.008931f
C555 VTAIL.n221 B 0.008435f
C556 VTAIL.n222 B 0.015697f
C557 VTAIL.n223 B 0.015697f
C558 VTAIL.n224 B 0.008435f
C559 VTAIL.n225 B 0.008931f
C560 VTAIL.n226 B 0.019937f
C561 VTAIL.n227 B 0.019937f
C562 VTAIL.n228 B 0.040726f
C563 VTAIL.n229 B 0.008683f
C564 VTAIL.n230 B 0.008435f
C565 VTAIL.n231 B 0.038642f
C566 VTAIL.n232 B 0.022608f
C567 VTAIL.n233 B 0.940234f
C568 VTAIL.n234 B 0.020687f
C569 VTAIL.n235 B 0.015697f
C570 VTAIL.n236 B 0.008683f
C571 VTAIL.n237 B 0.019937f
C572 VTAIL.n238 B 0.008931f
C573 VTAIL.n239 B 0.015697f
C574 VTAIL.n240 B 0.008435f
C575 VTAIL.n241 B 0.019937f
C576 VTAIL.n242 B 0.008931f
C577 VTAIL.n243 B 0.015697f
C578 VTAIL.n244 B 0.008435f
C579 VTAIL.n245 B 0.019937f
C580 VTAIL.n246 B 0.008931f
C581 VTAIL.n247 B 0.015697f
C582 VTAIL.n248 B 0.008435f
C583 VTAIL.n249 B 0.019937f
C584 VTAIL.n250 B 0.008931f
C585 VTAIL.n251 B 0.015697f
C586 VTAIL.n252 B 0.008435f
C587 VTAIL.n253 B 0.019937f
C588 VTAIL.n254 B 0.008931f
C589 VTAIL.n255 B 0.015697f
C590 VTAIL.n256 B 0.008435f
C591 VTAIL.n257 B 0.014953f
C592 VTAIL.n258 B 0.011778f
C593 VTAIL.t3 B 0.032822f
C594 VTAIL.n259 B 0.098563f
C595 VTAIL.n260 B 0.951506f
C596 VTAIL.n261 B 0.008435f
C597 VTAIL.n262 B 0.008931f
C598 VTAIL.n263 B 0.019937f
C599 VTAIL.n264 B 0.019937f
C600 VTAIL.n265 B 0.008931f
C601 VTAIL.n266 B 0.008435f
C602 VTAIL.n267 B 0.015697f
C603 VTAIL.n268 B 0.015697f
C604 VTAIL.n269 B 0.008435f
C605 VTAIL.n270 B 0.008931f
C606 VTAIL.n271 B 0.019937f
C607 VTAIL.n272 B 0.019937f
C608 VTAIL.n273 B 0.008931f
C609 VTAIL.n274 B 0.008435f
C610 VTAIL.n275 B 0.015697f
C611 VTAIL.n276 B 0.015697f
C612 VTAIL.n277 B 0.008435f
C613 VTAIL.n278 B 0.008931f
C614 VTAIL.n279 B 0.019937f
C615 VTAIL.n280 B 0.019937f
C616 VTAIL.n281 B 0.008931f
C617 VTAIL.n282 B 0.008435f
C618 VTAIL.n283 B 0.015697f
C619 VTAIL.n284 B 0.015697f
C620 VTAIL.n285 B 0.008435f
C621 VTAIL.n286 B 0.008931f
C622 VTAIL.n287 B 0.019937f
C623 VTAIL.n288 B 0.019937f
C624 VTAIL.n289 B 0.008931f
C625 VTAIL.n290 B 0.008435f
C626 VTAIL.n291 B 0.015697f
C627 VTAIL.n292 B 0.015697f
C628 VTAIL.n293 B 0.008435f
C629 VTAIL.n294 B 0.008931f
C630 VTAIL.n295 B 0.019937f
C631 VTAIL.n296 B 0.019937f
C632 VTAIL.n297 B 0.008931f
C633 VTAIL.n298 B 0.008435f
C634 VTAIL.n299 B 0.015697f
C635 VTAIL.n300 B 0.015697f
C636 VTAIL.n301 B 0.008435f
C637 VTAIL.n302 B 0.008435f
C638 VTAIL.n303 B 0.008931f
C639 VTAIL.n304 B 0.019937f
C640 VTAIL.n305 B 0.019937f
C641 VTAIL.n306 B 0.040726f
C642 VTAIL.n307 B 0.008683f
C643 VTAIL.n308 B 0.008435f
C644 VTAIL.n309 B 0.038642f
C645 VTAIL.n310 B 0.022608f
C646 VTAIL.n311 B 0.900882f
C647 VN.t1 B 1.53894f
C648 VN.t0 B 1.67517f
.ends

