* NGSPICE file created from diff_pair_sample_1588.ext - technology: sky130A

.subckt diff_pair_sample_1588 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VP.t0 VDD1.t0 w_n1876_n1932# sky130_fd_pr__pfet_01v8 ad=1.8798 pd=10.42 as=0.7953 ps=5.15 w=4.82 l=1.18
X1 B.t11 B.t9 B.t10 w_n1876_n1932# sky130_fd_pr__pfet_01v8 ad=1.8798 pd=10.42 as=0 ps=0 w=4.82 l=1.18
X2 B.t8 B.t6 B.t7 w_n1876_n1932# sky130_fd_pr__pfet_01v8 ad=1.8798 pd=10.42 as=0 ps=0 w=4.82 l=1.18
X3 VDD2.t3 VN.t0 VTAIL.t3 w_n1876_n1932# sky130_fd_pr__pfet_01v8 ad=0.7953 pd=5.15 as=1.8798 ps=10.42 w=4.82 l=1.18
X4 VTAIL.t0 VN.t1 VDD2.t2 w_n1876_n1932# sky130_fd_pr__pfet_01v8 ad=1.8798 pd=10.42 as=0.7953 ps=5.15 w=4.82 l=1.18
X5 VDD1.t3 VP.t1 VTAIL.t6 w_n1876_n1932# sky130_fd_pr__pfet_01v8 ad=0.7953 pd=5.15 as=1.8798 ps=10.42 w=4.82 l=1.18
X6 VDD2.t1 VN.t2 VTAIL.t1 w_n1876_n1932# sky130_fd_pr__pfet_01v8 ad=0.7953 pd=5.15 as=1.8798 ps=10.42 w=4.82 l=1.18
X7 B.t5 B.t3 B.t4 w_n1876_n1932# sky130_fd_pr__pfet_01v8 ad=1.8798 pd=10.42 as=0 ps=0 w=4.82 l=1.18
X8 VDD1.t1 VP.t2 VTAIL.t5 w_n1876_n1932# sky130_fd_pr__pfet_01v8 ad=0.7953 pd=5.15 as=1.8798 ps=10.42 w=4.82 l=1.18
X9 VTAIL.t2 VN.t3 VDD2.t0 w_n1876_n1932# sky130_fd_pr__pfet_01v8 ad=1.8798 pd=10.42 as=0.7953 ps=5.15 w=4.82 l=1.18
X10 B.t2 B.t0 B.t1 w_n1876_n1932# sky130_fd_pr__pfet_01v8 ad=1.8798 pd=10.42 as=0 ps=0 w=4.82 l=1.18
X11 VTAIL.t4 VP.t3 VDD1.t2 w_n1876_n1932# sky130_fd_pr__pfet_01v8 ad=1.8798 pd=10.42 as=0.7953 ps=5.15 w=4.82 l=1.18
R0 VP.n4 VP.n3 173.351
R1 VP.n10 VP.n9 173.351
R2 VP.n8 VP.n0 161.3
R3 VP.n7 VP.n6 161.3
R4 VP.n5 VP.n1 161.3
R5 VP.n2 VP.t0 134.29
R6 VP.n2 VP.t1 134.071
R7 VP.n3 VP.t3 98.4429
R8 VP.n9 VP.t2 98.4429
R9 VP.n4 VP.n2 54.9517
R10 VP.n7 VP.n1 40.577
R11 VP.n8 VP.n7 40.577
R12 VP.n3 VP.n1 12.5423
R13 VP.n9 VP.n8 12.5423
R14 VP.n5 VP.n4 0.189894
R15 VP.n6 VP.n5 0.189894
R16 VP.n6 VP.n0 0.189894
R17 VP.n10 VP.n0 0.189894
R18 VP VP.n10 0.0516364
R19 VDD1 VDD1.n1 130.802
R20 VDD1 VDD1.n0 98.5594
R21 VDD1.n0 VDD1.t0 6.74428
R22 VDD1.n0 VDD1.t3 6.74428
R23 VDD1.n1 VDD1.t2 6.74428
R24 VDD1.n1 VDD1.t1 6.74428
R25 VTAIL.n5 VTAIL.t7 88.5663
R26 VTAIL.n4 VTAIL.t3 88.5663
R27 VTAIL.n3 VTAIL.t2 88.5663
R28 VTAIL.n7 VTAIL.t1 88.5662
R29 VTAIL.n0 VTAIL.t0 88.5662
R30 VTAIL.n1 VTAIL.t5 88.5662
R31 VTAIL.n2 VTAIL.t4 88.5662
R32 VTAIL.n6 VTAIL.t6 88.5662
R33 VTAIL.n7 VTAIL.n6 17.8238
R34 VTAIL.n3 VTAIL.n2 17.8238
R35 VTAIL.n4 VTAIL.n3 1.30222
R36 VTAIL.n6 VTAIL.n5 1.30222
R37 VTAIL.n2 VTAIL.n1 1.30222
R38 VTAIL VTAIL.n0 0.709552
R39 VTAIL VTAIL.n7 0.593172
R40 VTAIL.n5 VTAIL.n4 0.470328
R41 VTAIL.n1 VTAIL.n0 0.470328
R42 B.n211 B.n64 585
R43 B.n210 B.n209 585
R44 B.n208 B.n65 585
R45 B.n207 B.n206 585
R46 B.n205 B.n66 585
R47 B.n204 B.n203 585
R48 B.n202 B.n67 585
R49 B.n201 B.n200 585
R50 B.n199 B.n68 585
R51 B.n198 B.n197 585
R52 B.n196 B.n69 585
R53 B.n195 B.n194 585
R54 B.n193 B.n70 585
R55 B.n192 B.n191 585
R56 B.n190 B.n71 585
R57 B.n189 B.n188 585
R58 B.n187 B.n72 585
R59 B.n186 B.n185 585
R60 B.n184 B.n73 585
R61 B.n183 B.n182 585
R62 B.n181 B.n74 585
R63 B.n180 B.n179 585
R64 B.n175 B.n75 585
R65 B.n174 B.n173 585
R66 B.n172 B.n76 585
R67 B.n171 B.n170 585
R68 B.n169 B.n77 585
R69 B.n168 B.n167 585
R70 B.n166 B.n78 585
R71 B.n165 B.n164 585
R72 B.n162 B.n79 585
R73 B.n161 B.n160 585
R74 B.n159 B.n82 585
R75 B.n158 B.n157 585
R76 B.n156 B.n83 585
R77 B.n155 B.n154 585
R78 B.n153 B.n84 585
R79 B.n152 B.n151 585
R80 B.n150 B.n85 585
R81 B.n149 B.n148 585
R82 B.n147 B.n86 585
R83 B.n146 B.n145 585
R84 B.n144 B.n87 585
R85 B.n143 B.n142 585
R86 B.n141 B.n88 585
R87 B.n140 B.n139 585
R88 B.n138 B.n89 585
R89 B.n137 B.n136 585
R90 B.n135 B.n90 585
R91 B.n134 B.n133 585
R92 B.n132 B.n91 585
R93 B.n213 B.n212 585
R94 B.n214 B.n63 585
R95 B.n216 B.n215 585
R96 B.n217 B.n62 585
R97 B.n219 B.n218 585
R98 B.n220 B.n61 585
R99 B.n222 B.n221 585
R100 B.n223 B.n60 585
R101 B.n225 B.n224 585
R102 B.n226 B.n59 585
R103 B.n228 B.n227 585
R104 B.n229 B.n58 585
R105 B.n231 B.n230 585
R106 B.n232 B.n57 585
R107 B.n234 B.n233 585
R108 B.n235 B.n56 585
R109 B.n237 B.n236 585
R110 B.n238 B.n55 585
R111 B.n240 B.n239 585
R112 B.n241 B.n54 585
R113 B.n243 B.n242 585
R114 B.n244 B.n53 585
R115 B.n246 B.n245 585
R116 B.n247 B.n52 585
R117 B.n249 B.n248 585
R118 B.n250 B.n51 585
R119 B.n252 B.n251 585
R120 B.n253 B.n50 585
R121 B.n255 B.n254 585
R122 B.n256 B.n49 585
R123 B.n258 B.n257 585
R124 B.n259 B.n48 585
R125 B.n261 B.n260 585
R126 B.n262 B.n47 585
R127 B.n264 B.n263 585
R128 B.n265 B.n46 585
R129 B.n267 B.n266 585
R130 B.n268 B.n45 585
R131 B.n270 B.n269 585
R132 B.n271 B.n44 585
R133 B.n273 B.n272 585
R134 B.n274 B.n43 585
R135 B.n276 B.n275 585
R136 B.n277 B.n42 585
R137 B.n356 B.n355 585
R138 B.n354 B.n13 585
R139 B.n353 B.n352 585
R140 B.n351 B.n14 585
R141 B.n350 B.n349 585
R142 B.n348 B.n15 585
R143 B.n347 B.n346 585
R144 B.n345 B.n16 585
R145 B.n344 B.n343 585
R146 B.n342 B.n17 585
R147 B.n341 B.n340 585
R148 B.n339 B.n18 585
R149 B.n338 B.n337 585
R150 B.n336 B.n19 585
R151 B.n335 B.n334 585
R152 B.n333 B.n20 585
R153 B.n332 B.n331 585
R154 B.n330 B.n21 585
R155 B.n329 B.n328 585
R156 B.n327 B.n22 585
R157 B.n326 B.n325 585
R158 B.n323 B.n23 585
R159 B.n322 B.n321 585
R160 B.n320 B.n26 585
R161 B.n319 B.n318 585
R162 B.n317 B.n27 585
R163 B.n316 B.n315 585
R164 B.n314 B.n28 585
R165 B.n313 B.n312 585
R166 B.n311 B.n29 585
R167 B.n309 B.n308 585
R168 B.n307 B.n32 585
R169 B.n306 B.n305 585
R170 B.n304 B.n33 585
R171 B.n303 B.n302 585
R172 B.n301 B.n34 585
R173 B.n300 B.n299 585
R174 B.n298 B.n35 585
R175 B.n297 B.n296 585
R176 B.n295 B.n36 585
R177 B.n294 B.n293 585
R178 B.n292 B.n37 585
R179 B.n291 B.n290 585
R180 B.n289 B.n38 585
R181 B.n288 B.n287 585
R182 B.n286 B.n39 585
R183 B.n285 B.n284 585
R184 B.n283 B.n40 585
R185 B.n282 B.n281 585
R186 B.n280 B.n41 585
R187 B.n279 B.n278 585
R188 B.n357 B.n12 585
R189 B.n359 B.n358 585
R190 B.n360 B.n11 585
R191 B.n362 B.n361 585
R192 B.n363 B.n10 585
R193 B.n365 B.n364 585
R194 B.n366 B.n9 585
R195 B.n368 B.n367 585
R196 B.n369 B.n8 585
R197 B.n371 B.n370 585
R198 B.n372 B.n7 585
R199 B.n374 B.n373 585
R200 B.n375 B.n6 585
R201 B.n377 B.n376 585
R202 B.n378 B.n5 585
R203 B.n380 B.n379 585
R204 B.n381 B.n4 585
R205 B.n383 B.n382 585
R206 B.n384 B.n3 585
R207 B.n386 B.n385 585
R208 B.n387 B.n0 585
R209 B.n2 B.n1 585
R210 B.n102 B.n101 585
R211 B.n104 B.n103 585
R212 B.n105 B.n100 585
R213 B.n107 B.n106 585
R214 B.n108 B.n99 585
R215 B.n110 B.n109 585
R216 B.n111 B.n98 585
R217 B.n113 B.n112 585
R218 B.n114 B.n97 585
R219 B.n116 B.n115 585
R220 B.n117 B.n96 585
R221 B.n119 B.n118 585
R222 B.n120 B.n95 585
R223 B.n122 B.n121 585
R224 B.n123 B.n94 585
R225 B.n125 B.n124 585
R226 B.n126 B.n93 585
R227 B.n128 B.n127 585
R228 B.n129 B.n92 585
R229 B.n131 B.n130 585
R230 B.n130 B.n91 454.062
R231 B.n212 B.n211 454.062
R232 B.n278 B.n277 454.062
R233 B.n357 B.n356 454.062
R234 B.n80 B.t6 302.454
R235 B.n176 B.t3 302.454
R236 B.n30 B.t9 302.454
R237 B.n24 B.t0 302.454
R238 B.n389 B.n388 256.663
R239 B.n388 B.n387 235.042
R240 B.n388 B.n2 235.042
R241 B.n134 B.n91 163.367
R242 B.n135 B.n134 163.367
R243 B.n136 B.n135 163.367
R244 B.n136 B.n89 163.367
R245 B.n140 B.n89 163.367
R246 B.n141 B.n140 163.367
R247 B.n142 B.n141 163.367
R248 B.n142 B.n87 163.367
R249 B.n146 B.n87 163.367
R250 B.n147 B.n146 163.367
R251 B.n148 B.n147 163.367
R252 B.n148 B.n85 163.367
R253 B.n152 B.n85 163.367
R254 B.n153 B.n152 163.367
R255 B.n154 B.n153 163.367
R256 B.n154 B.n83 163.367
R257 B.n158 B.n83 163.367
R258 B.n159 B.n158 163.367
R259 B.n160 B.n159 163.367
R260 B.n160 B.n79 163.367
R261 B.n165 B.n79 163.367
R262 B.n166 B.n165 163.367
R263 B.n167 B.n166 163.367
R264 B.n167 B.n77 163.367
R265 B.n171 B.n77 163.367
R266 B.n172 B.n171 163.367
R267 B.n173 B.n172 163.367
R268 B.n173 B.n75 163.367
R269 B.n180 B.n75 163.367
R270 B.n181 B.n180 163.367
R271 B.n182 B.n181 163.367
R272 B.n182 B.n73 163.367
R273 B.n186 B.n73 163.367
R274 B.n187 B.n186 163.367
R275 B.n188 B.n187 163.367
R276 B.n188 B.n71 163.367
R277 B.n192 B.n71 163.367
R278 B.n193 B.n192 163.367
R279 B.n194 B.n193 163.367
R280 B.n194 B.n69 163.367
R281 B.n198 B.n69 163.367
R282 B.n199 B.n198 163.367
R283 B.n200 B.n199 163.367
R284 B.n200 B.n67 163.367
R285 B.n204 B.n67 163.367
R286 B.n205 B.n204 163.367
R287 B.n206 B.n205 163.367
R288 B.n206 B.n65 163.367
R289 B.n210 B.n65 163.367
R290 B.n211 B.n210 163.367
R291 B.n277 B.n276 163.367
R292 B.n276 B.n43 163.367
R293 B.n272 B.n43 163.367
R294 B.n272 B.n271 163.367
R295 B.n271 B.n270 163.367
R296 B.n270 B.n45 163.367
R297 B.n266 B.n45 163.367
R298 B.n266 B.n265 163.367
R299 B.n265 B.n264 163.367
R300 B.n264 B.n47 163.367
R301 B.n260 B.n47 163.367
R302 B.n260 B.n259 163.367
R303 B.n259 B.n258 163.367
R304 B.n258 B.n49 163.367
R305 B.n254 B.n49 163.367
R306 B.n254 B.n253 163.367
R307 B.n253 B.n252 163.367
R308 B.n252 B.n51 163.367
R309 B.n248 B.n51 163.367
R310 B.n248 B.n247 163.367
R311 B.n247 B.n246 163.367
R312 B.n246 B.n53 163.367
R313 B.n242 B.n53 163.367
R314 B.n242 B.n241 163.367
R315 B.n241 B.n240 163.367
R316 B.n240 B.n55 163.367
R317 B.n236 B.n55 163.367
R318 B.n236 B.n235 163.367
R319 B.n235 B.n234 163.367
R320 B.n234 B.n57 163.367
R321 B.n230 B.n57 163.367
R322 B.n230 B.n229 163.367
R323 B.n229 B.n228 163.367
R324 B.n228 B.n59 163.367
R325 B.n224 B.n59 163.367
R326 B.n224 B.n223 163.367
R327 B.n223 B.n222 163.367
R328 B.n222 B.n61 163.367
R329 B.n218 B.n61 163.367
R330 B.n218 B.n217 163.367
R331 B.n217 B.n216 163.367
R332 B.n216 B.n63 163.367
R333 B.n212 B.n63 163.367
R334 B.n356 B.n13 163.367
R335 B.n352 B.n13 163.367
R336 B.n352 B.n351 163.367
R337 B.n351 B.n350 163.367
R338 B.n350 B.n15 163.367
R339 B.n346 B.n15 163.367
R340 B.n346 B.n345 163.367
R341 B.n345 B.n344 163.367
R342 B.n344 B.n17 163.367
R343 B.n340 B.n17 163.367
R344 B.n340 B.n339 163.367
R345 B.n339 B.n338 163.367
R346 B.n338 B.n19 163.367
R347 B.n334 B.n19 163.367
R348 B.n334 B.n333 163.367
R349 B.n333 B.n332 163.367
R350 B.n332 B.n21 163.367
R351 B.n328 B.n21 163.367
R352 B.n328 B.n327 163.367
R353 B.n327 B.n326 163.367
R354 B.n326 B.n23 163.367
R355 B.n321 B.n23 163.367
R356 B.n321 B.n320 163.367
R357 B.n320 B.n319 163.367
R358 B.n319 B.n27 163.367
R359 B.n315 B.n27 163.367
R360 B.n315 B.n314 163.367
R361 B.n314 B.n313 163.367
R362 B.n313 B.n29 163.367
R363 B.n308 B.n29 163.367
R364 B.n308 B.n307 163.367
R365 B.n307 B.n306 163.367
R366 B.n306 B.n33 163.367
R367 B.n302 B.n33 163.367
R368 B.n302 B.n301 163.367
R369 B.n301 B.n300 163.367
R370 B.n300 B.n35 163.367
R371 B.n296 B.n35 163.367
R372 B.n296 B.n295 163.367
R373 B.n295 B.n294 163.367
R374 B.n294 B.n37 163.367
R375 B.n290 B.n37 163.367
R376 B.n290 B.n289 163.367
R377 B.n289 B.n288 163.367
R378 B.n288 B.n39 163.367
R379 B.n284 B.n39 163.367
R380 B.n284 B.n283 163.367
R381 B.n283 B.n282 163.367
R382 B.n282 B.n41 163.367
R383 B.n278 B.n41 163.367
R384 B.n358 B.n357 163.367
R385 B.n358 B.n11 163.367
R386 B.n362 B.n11 163.367
R387 B.n363 B.n362 163.367
R388 B.n364 B.n363 163.367
R389 B.n364 B.n9 163.367
R390 B.n368 B.n9 163.367
R391 B.n369 B.n368 163.367
R392 B.n370 B.n369 163.367
R393 B.n370 B.n7 163.367
R394 B.n374 B.n7 163.367
R395 B.n375 B.n374 163.367
R396 B.n376 B.n375 163.367
R397 B.n376 B.n5 163.367
R398 B.n380 B.n5 163.367
R399 B.n381 B.n380 163.367
R400 B.n382 B.n381 163.367
R401 B.n382 B.n3 163.367
R402 B.n386 B.n3 163.367
R403 B.n387 B.n386 163.367
R404 B.n101 B.n2 163.367
R405 B.n104 B.n101 163.367
R406 B.n105 B.n104 163.367
R407 B.n106 B.n105 163.367
R408 B.n106 B.n99 163.367
R409 B.n110 B.n99 163.367
R410 B.n111 B.n110 163.367
R411 B.n112 B.n111 163.367
R412 B.n112 B.n97 163.367
R413 B.n116 B.n97 163.367
R414 B.n117 B.n116 163.367
R415 B.n118 B.n117 163.367
R416 B.n118 B.n95 163.367
R417 B.n122 B.n95 163.367
R418 B.n123 B.n122 163.367
R419 B.n124 B.n123 163.367
R420 B.n124 B.n93 163.367
R421 B.n128 B.n93 163.367
R422 B.n129 B.n128 163.367
R423 B.n130 B.n129 163.367
R424 B.n176 B.t4 145.21
R425 B.n30 B.t11 145.21
R426 B.n80 B.t7 145.207
R427 B.n24 B.t2 145.207
R428 B.n177 B.t5 115.925
R429 B.n31 B.t10 115.925
R430 B.n81 B.t8 115.921
R431 B.n25 B.t1 115.921
R432 B.n163 B.n81 59.5399
R433 B.n178 B.n177 59.5399
R434 B.n310 B.n31 59.5399
R435 B.n324 B.n25 59.5399
R436 B.n213 B.n64 29.5029
R437 B.n355 B.n12 29.5029
R438 B.n279 B.n42 29.5029
R439 B.n132 B.n131 29.5029
R440 B.n81 B.n80 29.2853
R441 B.n177 B.n176 29.2853
R442 B.n31 B.n30 29.2853
R443 B.n25 B.n24 29.2853
R444 B B.n389 18.0485
R445 B.n359 B.n12 10.6151
R446 B.n360 B.n359 10.6151
R447 B.n361 B.n360 10.6151
R448 B.n361 B.n10 10.6151
R449 B.n365 B.n10 10.6151
R450 B.n366 B.n365 10.6151
R451 B.n367 B.n366 10.6151
R452 B.n367 B.n8 10.6151
R453 B.n371 B.n8 10.6151
R454 B.n372 B.n371 10.6151
R455 B.n373 B.n372 10.6151
R456 B.n373 B.n6 10.6151
R457 B.n377 B.n6 10.6151
R458 B.n378 B.n377 10.6151
R459 B.n379 B.n378 10.6151
R460 B.n379 B.n4 10.6151
R461 B.n383 B.n4 10.6151
R462 B.n384 B.n383 10.6151
R463 B.n385 B.n384 10.6151
R464 B.n385 B.n0 10.6151
R465 B.n355 B.n354 10.6151
R466 B.n354 B.n353 10.6151
R467 B.n353 B.n14 10.6151
R468 B.n349 B.n14 10.6151
R469 B.n349 B.n348 10.6151
R470 B.n348 B.n347 10.6151
R471 B.n347 B.n16 10.6151
R472 B.n343 B.n16 10.6151
R473 B.n343 B.n342 10.6151
R474 B.n342 B.n341 10.6151
R475 B.n341 B.n18 10.6151
R476 B.n337 B.n18 10.6151
R477 B.n337 B.n336 10.6151
R478 B.n336 B.n335 10.6151
R479 B.n335 B.n20 10.6151
R480 B.n331 B.n20 10.6151
R481 B.n331 B.n330 10.6151
R482 B.n330 B.n329 10.6151
R483 B.n329 B.n22 10.6151
R484 B.n325 B.n22 10.6151
R485 B.n323 B.n322 10.6151
R486 B.n322 B.n26 10.6151
R487 B.n318 B.n26 10.6151
R488 B.n318 B.n317 10.6151
R489 B.n317 B.n316 10.6151
R490 B.n316 B.n28 10.6151
R491 B.n312 B.n28 10.6151
R492 B.n312 B.n311 10.6151
R493 B.n309 B.n32 10.6151
R494 B.n305 B.n32 10.6151
R495 B.n305 B.n304 10.6151
R496 B.n304 B.n303 10.6151
R497 B.n303 B.n34 10.6151
R498 B.n299 B.n34 10.6151
R499 B.n299 B.n298 10.6151
R500 B.n298 B.n297 10.6151
R501 B.n297 B.n36 10.6151
R502 B.n293 B.n36 10.6151
R503 B.n293 B.n292 10.6151
R504 B.n292 B.n291 10.6151
R505 B.n291 B.n38 10.6151
R506 B.n287 B.n38 10.6151
R507 B.n287 B.n286 10.6151
R508 B.n286 B.n285 10.6151
R509 B.n285 B.n40 10.6151
R510 B.n281 B.n40 10.6151
R511 B.n281 B.n280 10.6151
R512 B.n280 B.n279 10.6151
R513 B.n275 B.n42 10.6151
R514 B.n275 B.n274 10.6151
R515 B.n274 B.n273 10.6151
R516 B.n273 B.n44 10.6151
R517 B.n269 B.n44 10.6151
R518 B.n269 B.n268 10.6151
R519 B.n268 B.n267 10.6151
R520 B.n267 B.n46 10.6151
R521 B.n263 B.n46 10.6151
R522 B.n263 B.n262 10.6151
R523 B.n262 B.n261 10.6151
R524 B.n261 B.n48 10.6151
R525 B.n257 B.n48 10.6151
R526 B.n257 B.n256 10.6151
R527 B.n256 B.n255 10.6151
R528 B.n255 B.n50 10.6151
R529 B.n251 B.n50 10.6151
R530 B.n251 B.n250 10.6151
R531 B.n250 B.n249 10.6151
R532 B.n249 B.n52 10.6151
R533 B.n245 B.n52 10.6151
R534 B.n245 B.n244 10.6151
R535 B.n244 B.n243 10.6151
R536 B.n243 B.n54 10.6151
R537 B.n239 B.n54 10.6151
R538 B.n239 B.n238 10.6151
R539 B.n238 B.n237 10.6151
R540 B.n237 B.n56 10.6151
R541 B.n233 B.n56 10.6151
R542 B.n233 B.n232 10.6151
R543 B.n232 B.n231 10.6151
R544 B.n231 B.n58 10.6151
R545 B.n227 B.n58 10.6151
R546 B.n227 B.n226 10.6151
R547 B.n226 B.n225 10.6151
R548 B.n225 B.n60 10.6151
R549 B.n221 B.n60 10.6151
R550 B.n221 B.n220 10.6151
R551 B.n220 B.n219 10.6151
R552 B.n219 B.n62 10.6151
R553 B.n215 B.n62 10.6151
R554 B.n215 B.n214 10.6151
R555 B.n214 B.n213 10.6151
R556 B.n102 B.n1 10.6151
R557 B.n103 B.n102 10.6151
R558 B.n103 B.n100 10.6151
R559 B.n107 B.n100 10.6151
R560 B.n108 B.n107 10.6151
R561 B.n109 B.n108 10.6151
R562 B.n109 B.n98 10.6151
R563 B.n113 B.n98 10.6151
R564 B.n114 B.n113 10.6151
R565 B.n115 B.n114 10.6151
R566 B.n115 B.n96 10.6151
R567 B.n119 B.n96 10.6151
R568 B.n120 B.n119 10.6151
R569 B.n121 B.n120 10.6151
R570 B.n121 B.n94 10.6151
R571 B.n125 B.n94 10.6151
R572 B.n126 B.n125 10.6151
R573 B.n127 B.n126 10.6151
R574 B.n127 B.n92 10.6151
R575 B.n131 B.n92 10.6151
R576 B.n133 B.n132 10.6151
R577 B.n133 B.n90 10.6151
R578 B.n137 B.n90 10.6151
R579 B.n138 B.n137 10.6151
R580 B.n139 B.n138 10.6151
R581 B.n139 B.n88 10.6151
R582 B.n143 B.n88 10.6151
R583 B.n144 B.n143 10.6151
R584 B.n145 B.n144 10.6151
R585 B.n145 B.n86 10.6151
R586 B.n149 B.n86 10.6151
R587 B.n150 B.n149 10.6151
R588 B.n151 B.n150 10.6151
R589 B.n151 B.n84 10.6151
R590 B.n155 B.n84 10.6151
R591 B.n156 B.n155 10.6151
R592 B.n157 B.n156 10.6151
R593 B.n157 B.n82 10.6151
R594 B.n161 B.n82 10.6151
R595 B.n162 B.n161 10.6151
R596 B.n164 B.n78 10.6151
R597 B.n168 B.n78 10.6151
R598 B.n169 B.n168 10.6151
R599 B.n170 B.n169 10.6151
R600 B.n170 B.n76 10.6151
R601 B.n174 B.n76 10.6151
R602 B.n175 B.n174 10.6151
R603 B.n179 B.n175 10.6151
R604 B.n183 B.n74 10.6151
R605 B.n184 B.n183 10.6151
R606 B.n185 B.n184 10.6151
R607 B.n185 B.n72 10.6151
R608 B.n189 B.n72 10.6151
R609 B.n190 B.n189 10.6151
R610 B.n191 B.n190 10.6151
R611 B.n191 B.n70 10.6151
R612 B.n195 B.n70 10.6151
R613 B.n196 B.n195 10.6151
R614 B.n197 B.n196 10.6151
R615 B.n197 B.n68 10.6151
R616 B.n201 B.n68 10.6151
R617 B.n202 B.n201 10.6151
R618 B.n203 B.n202 10.6151
R619 B.n203 B.n66 10.6151
R620 B.n207 B.n66 10.6151
R621 B.n208 B.n207 10.6151
R622 B.n209 B.n208 10.6151
R623 B.n209 B.n64 10.6151
R624 B.n389 B.n0 8.11757
R625 B.n389 B.n1 8.11757
R626 B.n324 B.n323 6.5566
R627 B.n311 B.n310 6.5566
R628 B.n164 B.n163 6.5566
R629 B.n179 B.n178 6.5566
R630 B.n325 B.n324 4.05904
R631 B.n310 B.n309 4.05904
R632 B.n163 B.n162 4.05904
R633 B.n178 B.n74 4.05904
R634 VN.n0 VN.t1 134.29
R635 VN.n1 VN.t0 134.29
R636 VN.n0 VN.t2 134.071
R637 VN.n1 VN.t3 134.071
R638 VN VN.n1 55.3324
R639 VN VN.n0 18.5938
R640 VDD2.n2 VDD2.n0 130.276
R641 VDD2.n2 VDD2.n1 98.5012
R642 VDD2.n1 VDD2.t0 6.74428
R643 VDD2.n1 VDD2.t3 6.74428
R644 VDD2.n0 VDD2.t2 6.74428
R645 VDD2.n0 VDD2.t1 6.74428
R646 VDD2 VDD2.n2 0.0586897
C0 VDD2 VP 0.308251f
C1 VDD1 VP 1.89975f
C2 VTAIL VN 1.79847f
C3 VP B 1.14738f
C4 VTAIL w_n1876_n1932# 2.29058f
C5 VDD2 VDD1 0.679573f
C6 VP VN 3.83831f
C7 VDD2 B 0.846807f
C8 VDD1 B 0.817732f
C9 VP w_n1876_n1932# 3.02169f
C10 VDD2 VN 1.74393f
C11 VDD1 VN 0.151701f
C12 VDD2 w_n1876_n1932# 0.996949f
C13 VTAIL VP 1.81258f
C14 B VN 0.759829f
C15 VDD1 w_n1876_n1932# 0.972619f
C16 B w_n1876_n1932# 5.48822f
C17 VDD2 VTAIL 3.41157f
C18 VDD1 VTAIL 3.36688f
C19 VN w_n1876_n1932# 2.7842f
C20 VTAIL B 2.07456f
C21 VDD2 VSUBS 0.515394f
C22 VDD1 VSUBS 2.77539f
C23 VTAIL VSUBS 0.485174f
C24 VN VSUBS 3.81085f
C25 VP VSUBS 1.166238f
C26 B VSUBS 2.325109f
C27 w_n1876_n1932# VSUBS 45.4517f
C28 VDD2.t2 VSUBS 0.068082f
C29 VDD2.t1 VSUBS 0.068082f
C30 VDD2.n0 VSUBS 0.633635f
C31 VDD2.t0 VSUBS 0.068082f
C32 VDD2.t3 VSUBS 0.068082f
C33 VDD2.n1 VSUBS 0.421744f
C34 VDD2.n2 VSUBS 1.99347f
C35 VN.t1 VSUBS 0.657933f
C36 VN.t2 VSUBS 0.657316f
C37 VN.n0 VSUBS 0.556656f
C38 VN.t0 VSUBS 0.657933f
C39 VN.t3 VSUBS 0.657316f
C40 VN.n1 VSUBS 1.49249f
C41 B.n0 VSUBS 0.008367f
C42 B.n1 VSUBS 0.008367f
C43 B.n2 VSUBS 0.012374f
C44 B.n3 VSUBS 0.009483f
C45 B.n4 VSUBS 0.009483f
C46 B.n5 VSUBS 0.009483f
C47 B.n6 VSUBS 0.009483f
C48 B.n7 VSUBS 0.009483f
C49 B.n8 VSUBS 0.009483f
C50 B.n9 VSUBS 0.009483f
C51 B.n10 VSUBS 0.009483f
C52 B.n11 VSUBS 0.009483f
C53 B.n12 VSUBS 0.020037f
C54 B.n13 VSUBS 0.009483f
C55 B.n14 VSUBS 0.009483f
C56 B.n15 VSUBS 0.009483f
C57 B.n16 VSUBS 0.009483f
C58 B.n17 VSUBS 0.009483f
C59 B.n18 VSUBS 0.009483f
C60 B.n19 VSUBS 0.009483f
C61 B.n20 VSUBS 0.009483f
C62 B.n21 VSUBS 0.009483f
C63 B.n22 VSUBS 0.009483f
C64 B.n23 VSUBS 0.009483f
C65 B.t1 VSUBS 0.180827f
C66 B.t2 VSUBS 0.195556f
C67 B.t0 VSUBS 0.352417f
C68 B.n24 VSUBS 0.117137f
C69 B.n25 VSUBS 0.086559f
C70 B.n26 VSUBS 0.009483f
C71 B.n27 VSUBS 0.009483f
C72 B.n28 VSUBS 0.009483f
C73 B.n29 VSUBS 0.009483f
C74 B.t10 VSUBS 0.180827f
C75 B.t11 VSUBS 0.195556f
C76 B.t9 VSUBS 0.352417f
C77 B.n30 VSUBS 0.117138f
C78 B.n31 VSUBS 0.086559f
C79 B.n32 VSUBS 0.009483f
C80 B.n33 VSUBS 0.009483f
C81 B.n34 VSUBS 0.009483f
C82 B.n35 VSUBS 0.009483f
C83 B.n36 VSUBS 0.009483f
C84 B.n37 VSUBS 0.009483f
C85 B.n38 VSUBS 0.009483f
C86 B.n39 VSUBS 0.009483f
C87 B.n40 VSUBS 0.009483f
C88 B.n41 VSUBS 0.009483f
C89 B.n42 VSUBS 0.020037f
C90 B.n43 VSUBS 0.009483f
C91 B.n44 VSUBS 0.009483f
C92 B.n45 VSUBS 0.009483f
C93 B.n46 VSUBS 0.009483f
C94 B.n47 VSUBS 0.009483f
C95 B.n48 VSUBS 0.009483f
C96 B.n49 VSUBS 0.009483f
C97 B.n50 VSUBS 0.009483f
C98 B.n51 VSUBS 0.009483f
C99 B.n52 VSUBS 0.009483f
C100 B.n53 VSUBS 0.009483f
C101 B.n54 VSUBS 0.009483f
C102 B.n55 VSUBS 0.009483f
C103 B.n56 VSUBS 0.009483f
C104 B.n57 VSUBS 0.009483f
C105 B.n58 VSUBS 0.009483f
C106 B.n59 VSUBS 0.009483f
C107 B.n60 VSUBS 0.009483f
C108 B.n61 VSUBS 0.009483f
C109 B.n62 VSUBS 0.009483f
C110 B.n63 VSUBS 0.009483f
C111 B.n64 VSUBS 0.020279f
C112 B.n65 VSUBS 0.009483f
C113 B.n66 VSUBS 0.009483f
C114 B.n67 VSUBS 0.009483f
C115 B.n68 VSUBS 0.009483f
C116 B.n69 VSUBS 0.009483f
C117 B.n70 VSUBS 0.009483f
C118 B.n71 VSUBS 0.009483f
C119 B.n72 VSUBS 0.009483f
C120 B.n73 VSUBS 0.009483f
C121 B.n74 VSUBS 0.006554f
C122 B.n75 VSUBS 0.009483f
C123 B.n76 VSUBS 0.009483f
C124 B.n77 VSUBS 0.009483f
C125 B.n78 VSUBS 0.009483f
C126 B.n79 VSUBS 0.009483f
C127 B.t8 VSUBS 0.180827f
C128 B.t7 VSUBS 0.195556f
C129 B.t6 VSUBS 0.352417f
C130 B.n80 VSUBS 0.117137f
C131 B.n81 VSUBS 0.086559f
C132 B.n82 VSUBS 0.009483f
C133 B.n83 VSUBS 0.009483f
C134 B.n84 VSUBS 0.009483f
C135 B.n85 VSUBS 0.009483f
C136 B.n86 VSUBS 0.009483f
C137 B.n87 VSUBS 0.009483f
C138 B.n88 VSUBS 0.009483f
C139 B.n89 VSUBS 0.009483f
C140 B.n90 VSUBS 0.009483f
C141 B.n91 VSUBS 0.021519f
C142 B.n92 VSUBS 0.009483f
C143 B.n93 VSUBS 0.009483f
C144 B.n94 VSUBS 0.009483f
C145 B.n95 VSUBS 0.009483f
C146 B.n96 VSUBS 0.009483f
C147 B.n97 VSUBS 0.009483f
C148 B.n98 VSUBS 0.009483f
C149 B.n99 VSUBS 0.009483f
C150 B.n100 VSUBS 0.009483f
C151 B.n101 VSUBS 0.009483f
C152 B.n102 VSUBS 0.009483f
C153 B.n103 VSUBS 0.009483f
C154 B.n104 VSUBS 0.009483f
C155 B.n105 VSUBS 0.009483f
C156 B.n106 VSUBS 0.009483f
C157 B.n107 VSUBS 0.009483f
C158 B.n108 VSUBS 0.009483f
C159 B.n109 VSUBS 0.009483f
C160 B.n110 VSUBS 0.009483f
C161 B.n111 VSUBS 0.009483f
C162 B.n112 VSUBS 0.009483f
C163 B.n113 VSUBS 0.009483f
C164 B.n114 VSUBS 0.009483f
C165 B.n115 VSUBS 0.009483f
C166 B.n116 VSUBS 0.009483f
C167 B.n117 VSUBS 0.009483f
C168 B.n118 VSUBS 0.009483f
C169 B.n119 VSUBS 0.009483f
C170 B.n120 VSUBS 0.009483f
C171 B.n121 VSUBS 0.009483f
C172 B.n122 VSUBS 0.009483f
C173 B.n123 VSUBS 0.009483f
C174 B.n124 VSUBS 0.009483f
C175 B.n125 VSUBS 0.009483f
C176 B.n126 VSUBS 0.009483f
C177 B.n127 VSUBS 0.009483f
C178 B.n128 VSUBS 0.009483f
C179 B.n129 VSUBS 0.009483f
C180 B.n130 VSUBS 0.020037f
C181 B.n131 VSUBS 0.020037f
C182 B.n132 VSUBS 0.021519f
C183 B.n133 VSUBS 0.009483f
C184 B.n134 VSUBS 0.009483f
C185 B.n135 VSUBS 0.009483f
C186 B.n136 VSUBS 0.009483f
C187 B.n137 VSUBS 0.009483f
C188 B.n138 VSUBS 0.009483f
C189 B.n139 VSUBS 0.009483f
C190 B.n140 VSUBS 0.009483f
C191 B.n141 VSUBS 0.009483f
C192 B.n142 VSUBS 0.009483f
C193 B.n143 VSUBS 0.009483f
C194 B.n144 VSUBS 0.009483f
C195 B.n145 VSUBS 0.009483f
C196 B.n146 VSUBS 0.009483f
C197 B.n147 VSUBS 0.009483f
C198 B.n148 VSUBS 0.009483f
C199 B.n149 VSUBS 0.009483f
C200 B.n150 VSUBS 0.009483f
C201 B.n151 VSUBS 0.009483f
C202 B.n152 VSUBS 0.009483f
C203 B.n153 VSUBS 0.009483f
C204 B.n154 VSUBS 0.009483f
C205 B.n155 VSUBS 0.009483f
C206 B.n156 VSUBS 0.009483f
C207 B.n157 VSUBS 0.009483f
C208 B.n158 VSUBS 0.009483f
C209 B.n159 VSUBS 0.009483f
C210 B.n160 VSUBS 0.009483f
C211 B.n161 VSUBS 0.009483f
C212 B.n162 VSUBS 0.006554f
C213 B.n163 VSUBS 0.02197f
C214 B.n164 VSUBS 0.00767f
C215 B.n165 VSUBS 0.009483f
C216 B.n166 VSUBS 0.009483f
C217 B.n167 VSUBS 0.009483f
C218 B.n168 VSUBS 0.009483f
C219 B.n169 VSUBS 0.009483f
C220 B.n170 VSUBS 0.009483f
C221 B.n171 VSUBS 0.009483f
C222 B.n172 VSUBS 0.009483f
C223 B.n173 VSUBS 0.009483f
C224 B.n174 VSUBS 0.009483f
C225 B.n175 VSUBS 0.009483f
C226 B.t5 VSUBS 0.180827f
C227 B.t4 VSUBS 0.195556f
C228 B.t3 VSUBS 0.352417f
C229 B.n176 VSUBS 0.117138f
C230 B.n177 VSUBS 0.086559f
C231 B.n178 VSUBS 0.02197f
C232 B.n179 VSUBS 0.00767f
C233 B.n180 VSUBS 0.009483f
C234 B.n181 VSUBS 0.009483f
C235 B.n182 VSUBS 0.009483f
C236 B.n183 VSUBS 0.009483f
C237 B.n184 VSUBS 0.009483f
C238 B.n185 VSUBS 0.009483f
C239 B.n186 VSUBS 0.009483f
C240 B.n187 VSUBS 0.009483f
C241 B.n188 VSUBS 0.009483f
C242 B.n189 VSUBS 0.009483f
C243 B.n190 VSUBS 0.009483f
C244 B.n191 VSUBS 0.009483f
C245 B.n192 VSUBS 0.009483f
C246 B.n193 VSUBS 0.009483f
C247 B.n194 VSUBS 0.009483f
C248 B.n195 VSUBS 0.009483f
C249 B.n196 VSUBS 0.009483f
C250 B.n197 VSUBS 0.009483f
C251 B.n198 VSUBS 0.009483f
C252 B.n199 VSUBS 0.009483f
C253 B.n200 VSUBS 0.009483f
C254 B.n201 VSUBS 0.009483f
C255 B.n202 VSUBS 0.009483f
C256 B.n203 VSUBS 0.009483f
C257 B.n204 VSUBS 0.009483f
C258 B.n205 VSUBS 0.009483f
C259 B.n206 VSUBS 0.009483f
C260 B.n207 VSUBS 0.009483f
C261 B.n208 VSUBS 0.009483f
C262 B.n209 VSUBS 0.009483f
C263 B.n210 VSUBS 0.009483f
C264 B.n211 VSUBS 0.021519f
C265 B.n212 VSUBS 0.020037f
C266 B.n213 VSUBS 0.021277f
C267 B.n214 VSUBS 0.009483f
C268 B.n215 VSUBS 0.009483f
C269 B.n216 VSUBS 0.009483f
C270 B.n217 VSUBS 0.009483f
C271 B.n218 VSUBS 0.009483f
C272 B.n219 VSUBS 0.009483f
C273 B.n220 VSUBS 0.009483f
C274 B.n221 VSUBS 0.009483f
C275 B.n222 VSUBS 0.009483f
C276 B.n223 VSUBS 0.009483f
C277 B.n224 VSUBS 0.009483f
C278 B.n225 VSUBS 0.009483f
C279 B.n226 VSUBS 0.009483f
C280 B.n227 VSUBS 0.009483f
C281 B.n228 VSUBS 0.009483f
C282 B.n229 VSUBS 0.009483f
C283 B.n230 VSUBS 0.009483f
C284 B.n231 VSUBS 0.009483f
C285 B.n232 VSUBS 0.009483f
C286 B.n233 VSUBS 0.009483f
C287 B.n234 VSUBS 0.009483f
C288 B.n235 VSUBS 0.009483f
C289 B.n236 VSUBS 0.009483f
C290 B.n237 VSUBS 0.009483f
C291 B.n238 VSUBS 0.009483f
C292 B.n239 VSUBS 0.009483f
C293 B.n240 VSUBS 0.009483f
C294 B.n241 VSUBS 0.009483f
C295 B.n242 VSUBS 0.009483f
C296 B.n243 VSUBS 0.009483f
C297 B.n244 VSUBS 0.009483f
C298 B.n245 VSUBS 0.009483f
C299 B.n246 VSUBS 0.009483f
C300 B.n247 VSUBS 0.009483f
C301 B.n248 VSUBS 0.009483f
C302 B.n249 VSUBS 0.009483f
C303 B.n250 VSUBS 0.009483f
C304 B.n251 VSUBS 0.009483f
C305 B.n252 VSUBS 0.009483f
C306 B.n253 VSUBS 0.009483f
C307 B.n254 VSUBS 0.009483f
C308 B.n255 VSUBS 0.009483f
C309 B.n256 VSUBS 0.009483f
C310 B.n257 VSUBS 0.009483f
C311 B.n258 VSUBS 0.009483f
C312 B.n259 VSUBS 0.009483f
C313 B.n260 VSUBS 0.009483f
C314 B.n261 VSUBS 0.009483f
C315 B.n262 VSUBS 0.009483f
C316 B.n263 VSUBS 0.009483f
C317 B.n264 VSUBS 0.009483f
C318 B.n265 VSUBS 0.009483f
C319 B.n266 VSUBS 0.009483f
C320 B.n267 VSUBS 0.009483f
C321 B.n268 VSUBS 0.009483f
C322 B.n269 VSUBS 0.009483f
C323 B.n270 VSUBS 0.009483f
C324 B.n271 VSUBS 0.009483f
C325 B.n272 VSUBS 0.009483f
C326 B.n273 VSUBS 0.009483f
C327 B.n274 VSUBS 0.009483f
C328 B.n275 VSUBS 0.009483f
C329 B.n276 VSUBS 0.009483f
C330 B.n277 VSUBS 0.020037f
C331 B.n278 VSUBS 0.021519f
C332 B.n279 VSUBS 0.021519f
C333 B.n280 VSUBS 0.009483f
C334 B.n281 VSUBS 0.009483f
C335 B.n282 VSUBS 0.009483f
C336 B.n283 VSUBS 0.009483f
C337 B.n284 VSUBS 0.009483f
C338 B.n285 VSUBS 0.009483f
C339 B.n286 VSUBS 0.009483f
C340 B.n287 VSUBS 0.009483f
C341 B.n288 VSUBS 0.009483f
C342 B.n289 VSUBS 0.009483f
C343 B.n290 VSUBS 0.009483f
C344 B.n291 VSUBS 0.009483f
C345 B.n292 VSUBS 0.009483f
C346 B.n293 VSUBS 0.009483f
C347 B.n294 VSUBS 0.009483f
C348 B.n295 VSUBS 0.009483f
C349 B.n296 VSUBS 0.009483f
C350 B.n297 VSUBS 0.009483f
C351 B.n298 VSUBS 0.009483f
C352 B.n299 VSUBS 0.009483f
C353 B.n300 VSUBS 0.009483f
C354 B.n301 VSUBS 0.009483f
C355 B.n302 VSUBS 0.009483f
C356 B.n303 VSUBS 0.009483f
C357 B.n304 VSUBS 0.009483f
C358 B.n305 VSUBS 0.009483f
C359 B.n306 VSUBS 0.009483f
C360 B.n307 VSUBS 0.009483f
C361 B.n308 VSUBS 0.009483f
C362 B.n309 VSUBS 0.006554f
C363 B.n310 VSUBS 0.02197f
C364 B.n311 VSUBS 0.00767f
C365 B.n312 VSUBS 0.009483f
C366 B.n313 VSUBS 0.009483f
C367 B.n314 VSUBS 0.009483f
C368 B.n315 VSUBS 0.009483f
C369 B.n316 VSUBS 0.009483f
C370 B.n317 VSUBS 0.009483f
C371 B.n318 VSUBS 0.009483f
C372 B.n319 VSUBS 0.009483f
C373 B.n320 VSUBS 0.009483f
C374 B.n321 VSUBS 0.009483f
C375 B.n322 VSUBS 0.009483f
C376 B.n323 VSUBS 0.00767f
C377 B.n324 VSUBS 0.02197f
C378 B.n325 VSUBS 0.006554f
C379 B.n326 VSUBS 0.009483f
C380 B.n327 VSUBS 0.009483f
C381 B.n328 VSUBS 0.009483f
C382 B.n329 VSUBS 0.009483f
C383 B.n330 VSUBS 0.009483f
C384 B.n331 VSUBS 0.009483f
C385 B.n332 VSUBS 0.009483f
C386 B.n333 VSUBS 0.009483f
C387 B.n334 VSUBS 0.009483f
C388 B.n335 VSUBS 0.009483f
C389 B.n336 VSUBS 0.009483f
C390 B.n337 VSUBS 0.009483f
C391 B.n338 VSUBS 0.009483f
C392 B.n339 VSUBS 0.009483f
C393 B.n340 VSUBS 0.009483f
C394 B.n341 VSUBS 0.009483f
C395 B.n342 VSUBS 0.009483f
C396 B.n343 VSUBS 0.009483f
C397 B.n344 VSUBS 0.009483f
C398 B.n345 VSUBS 0.009483f
C399 B.n346 VSUBS 0.009483f
C400 B.n347 VSUBS 0.009483f
C401 B.n348 VSUBS 0.009483f
C402 B.n349 VSUBS 0.009483f
C403 B.n350 VSUBS 0.009483f
C404 B.n351 VSUBS 0.009483f
C405 B.n352 VSUBS 0.009483f
C406 B.n353 VSUBS 0.009483f
C407 B.n354 VSUBS 0.009483f
C408 B.n355 VSUBS 0.021519f
C409 B.n356 VSUBS 0.021519f
C410 B.n357 VSUBS 0.020037f
C411 B.n358 VSUBS 0.009483f
C412 B.n359 VSUBS 0.009483f
C413 B.n360 VSUBS 0.009483f
C414 B.n361 VSUBS 0.009483f
C415 B.n362 VSUBS 0.009483f
C416 B.n363 VSUBS 0.009483f
C417 B.n364 VSUBS 0.009483f
C418 B.n365 VSUBS 0.009483f
C419 B.n366 VSUBS 0.009483f
C420 B.n367 VSUBS 0.009483f
C421 B.n368 VSUBS 0.009483f
C422 B.n369 VSUBS 0.009483f
C423 B.n370 VSUBS 0.009483f
C424 B.n371 VSUBS 0.009483f
C425 B.n372 VSUBS 0.009483f
C426 B.n373 VSUBS 0.009483f
C427 B.n374 VSUBS 0.009483f
C428 B.n375 VSUBS 0.009483f
C429 B.n376 VSUBS 0.009483f
C430 B.n377 VSUBS 0.009483f
C431 B.n378 VSUBS 0.009483f
C432 B.n379 VSUBS 0.009483f
C433 B.n380 VSUBS 0.009483f
C434 B.n381 VSUBS 0.009483f
C435 B.n382 VSUBS 0.009483f
C436 B.n383 VSUBS 0.009483f
C437 B.n384 VSUBS 0.009483f
C438 B.n385 VSUBS 0.009483f
C439 B.n386 VSUBS 0.009483f
C440 B.n387 VSUBS 0.012374f
C441 B.n388 VSUBS 0.013182f
C442 B.n389 VSUBS 0.026213f
C443 VTAIL.t0 VSUBS 0.591132f
C444 VTAIL.n0 VSUBS 0.466064f
C445 VTAIL.t5 VSUBS 0.591132f
C446 VTAIL.n1 VSUBS 0.50518f
C447 VTAIL.t4 VSUBS 0.591132f
C448 VTAIL.n2 VSUBS 1.11256f
C449 VTAIL.t2 VSUBS 0.591135f
C450 VTAIL.n3 VSUBS 1.11255f
C451 VTAIL.t3 VSUBS 0.591135f
C452 VTAIL.n4 VSUBS 0.505177f
C453 VTAIL.t7 VSUBS 0.591135f
C454 VTAIL.n5 VSUBS 0.505177f
C455 VTAIL.t6 VSUBS 0.591132f
C456 VTAIL.n6 VSUBS 1.11256f
C457 VTAIL.t1 VSUBS 0.591132f
C458 VTAIL.n7 VSUBS 1.06576f
C459 VDD1.t0 VSUBS 0.066785f
C460 VDD1.t3 VSUBS 0.066785f
C461 VDD1.n0 VSUBS 0.413917f
C462 VDD1.t2 VSUBS 0.066785f
C463 VDD1.t1 VSUBS 0.066785f
C464 VDD1.n1 VSUBS 0.633019f
C465 VP.n0 VSUBS 0.039448f
C466 VP.t2 VSUBS 0.585292f
C467 VP.n1 VSUBS 0.060294f
C468 VP.t0 VSUBS 0.683398f
C469 VP.t1 VSUBS 0.682757f
C470 VP.n2 VSUBS 1.52954f
C471 VP.t3 VSUBS 0.585292f
C472 VP.n3 VSUBS 0.309405f
C473 VP.n4 VSUBS 1.79529f
C474 VP.n5 VSUBS 0.039448f
C475 VP.n6 VSUBS 0.039448f
C476 VP.n7 VSUBS 0.031861f
C477 VP.n8 VSUBS 0.060294f
C478 VP.n9 VSUBS 0.309405f
C479 VP.n10 VSUBS 0.035329f
.ends

