* NGSPICE file created from diff_pair_sample_0682.ext - technology: sky130A

.subckt diff_pair_sample_0682 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VP.t0 VDD1.t0 B.t5 sky130_fd_pr__nfet_01v8 ad=0.57585 pd=3.82 as=0.57585 ps=3.82 w=3.49 l=0.3
X1 VDD2.t7 VN.t0 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=0.57585 pd=3.82 as=0.57585 ps=3.82 w=3.49 l=0.3
X2 VTAIL.t14 VP.t1 VDD1.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=1.3611 pd=7.76 as=0.57585 ps=3.82 w=3.49 l=0.3
X3 VDD2.t6 VN.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.57585 pd=3.82 as=1.3611 ps=7.76 w=3.49 l=0.3
X4 VDD2.t5 VN.t2 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=0.57585 pd=3.82 as=0.57585 ps=3.82 w=3.49 l=0.3
X5 VTAIL.t13 VP.t2 VDD1.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=1.3611 pd=7.76 as=0.57585 ps=3.82 w=3.49 l=0.3
X6 B.t21 B.t19 B.t20 B.t16 sky130_fd_pr__nfet_01v8 ad=1.3611 pd=7.76 as=0 ps=0 w=3.49 l=0.3
X7 VDD1.t3 VP.t3 VTAIL.t12 B.t1 sky130_fd_pr__nfet_01v8 ad=0.57585 pd=3.82 as=1.3611 ps=7.76 w=3.49 l=0.3
X8 VDD1.t4 VP.t4 VTAIL.t11 B.t6 sky130_fd_pr__nfet_01v8 ad=0.57585 pd=3.82 as=0.57585 ps=3.82 w=3.49 l=0.3
X9 VDD1.t5 VP.t5 VTAIL.t10 B.t7 sky130_fd_pr__nfet_01v8 ad=0.57585 pd=3.82 as=0.57585 ps=3.82 w=3.49 l=0.3
X10 VTAIL.t2 VN.t3 VDD2.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=0.57585 pd=3.82 as=0.57585 ps=3.82 w=3.49 l=0.3
X11 VTAIL.t3 VN.t4 VDD2.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.3611 pd=7.76 as=0.57585 ps=3.82 w=3.49 l=0.3
X12 VTAIL.t4 VN.t5 VDD2.t2 B.t4 sky130_fd_pr__nfet_01v8 ad=1.3611 pd=7.76 as=0.57585 ps=3.82 w=3.49 l=0.3
X13 VDD2.t1 VN.t6 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.57585 pd=3.82 as=1.3611 ps=7.76 w=3.49 l=0.3
X14 B.t18 B.t15 B.t17 B.t16 sky130_fd_pr__nfet_01v8 ad=1.3611 pd=7.76 as=0 ps=0 w=3.49 l=0.3
X15 VTAIL.t9 VP.t6 VDD1.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=0.57585 pd=3.82 as=0.57585 ps=3.82 w=3.49 l=0.3
X16 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=1.3611 pd=7.76 as=0 ps=0 w=3.49 l=0.3
X17 VTAIL.t5 VN.t7 VDD2.t0 B.t5 sky130_fd_pr__nfet_01v8 ad=0.57585 pd=3.82 as=0.57585 ps=3.82 w=3.49 l=0.3
X18 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=1.3611 pd=7.76 as=0 ps=0 w=3.49 l=0.3
X19 VDD1.t7 VP.t7 VTAIL.t8 B.t0 sky130_fd_pr__nfet_01v8 ad=0.57585 pd=3.82 as=1.3611 ps=7.76 w=3.49 l=0.3
R0 VP.n17 VP.t3 414.082
R1 VP.n11 VP.t1 414.082
R2 VP.n4 VP.t2 414.082
R3 VP.n9 VP.t7 414.082
R4 VP.n16 VP.t0 385.601
R5 VP.n1 VP.t4 385.601
R6 VP.n3 VP.t5 385.601
R7 VP.n8 VP.t6 385.601
R8 VP.n5 VP.n4 161.489
R9 VP.n18 VP.n17 161.3
R10 VP.n6 VP.n5 161.3
R11 VP.n7 VP.n2 161.3
R12 VP.n10 VP.n9 161.3
R13 VP.n15 VP.n0 161.3
R14 VP.n14 VP.n13 161.3
R15 VP.n12 VP.n11 161.3
R16 VP.n15 VP.n14 73.0308
R17 VP.n7 VP.n6 73.0308
R18 VP.n11 VP.n1 63.5369
R19 VP.n17 VP.n16 63.5369
R20 VP.n4 VP.n3 63.5369
R21 VP.n9 VP.n8 63.5369
R22 VP.n12 VP.n10 33.6899
R23 VP.n14 VP.n1 9.49444
R24 VP.n16 VP.n15 9.49444
R25 VP.n6 VP.n3 9.49444
R26 VP.n8 VP.n7 9.49444
R27 VP.n5 VP.n2 0.189894
R28 VP.n10 VP.n2 0.189894
R29 VP.n13 VP.n12 0.189894
R30 VP.n13 VP.n0 0.189894
R31 VP.n18 VP.n0 0.189894
R32 VP VP.n18 0.0516364
R33 VDD1 VDD1.n0 75.8843
R34 VDD1.n3 VDD1.n2 75.7706
R35 VDD1.n3 VDD1.n1 75.7706
R36 VDD1.n5 VDD1.n4 75.5545
R37 VDD1.n5 VDD1.n3 29.7509
R38 VDD1.n4 VDD1.t6 5.67385
R39 VDD1.n4 VDD1.t7 5.67385
R40 VDD1.n0 VDD1.t2 5.67385
R41 VDD1.n0 VDD1.t5 5.67385
R42 VDD1.n2 VDD1.t0 5.67385
R43 VDD1.n2 VDD1.t3 5.67385
R44 VDD1.n1 VDD1.t1 5.67385
R45 VDD1.n1 VDD1.t4 5.67385
R46 VDD1 VDD1.n5 0.213862
R47 VTAIL.n11 VTAIL.t13 64.549
R48 VTAIL.n10 VTAIL.t1 64.549
R49 VTAIL.n7 VTAIL.t4 64.549
R50 VTAIL.n15 VTAIL.t0 64.549
R51 VTAIL.n2 VTAIL.t3 64.549
R52 VTAIL.n3 VTAIL.t12 64.549
R53 VTAIL.n6 VTAIL.t14 64.549
R54 VTAIL.n14 VTAIL.t8 64.549
R55 VTAIL.n13 VTAIL.n12 58.8758
R56 VTAIL.n9 VTAIL.n8 58.8758
R57 VTAIL.n1 VTAIL.n0 58.8756
R58 VTAIL.n5 VTAIL.n4 58.8756
R59 VTAIL.n15 VTAIL.n14 15.9186
R60 VTAIL.n7 VTAIL.n6 15.9186
R61 VTAIL.n0 VTAIL.t7 5.67385
R62 VTAIL.n0 VTAIL.t2 5.67385
R63 VTAIL.n4 VTAIL.t11 5.67385
R64 VTAIL.n4 VTAIL.t15 5.67385
R65 VTAIL.n12 VTAIL.t10 5.67385
R66 VTAIL.n12 VTAIL.t9 5.67385
R67 VTAIL.n8 VTAIL.t6 5.67385
R68 VTAIL.n8 VTAIL.t5 5.67385
R69 VTAIL.n9 VTAIL.n7 0.543603
R70 VTAIL.n10 VTAIL.n9 0.543603
R71 VTAIL.n13 VTAIL.n11 0.543603
R72 VTAIL.n14 VTAIL.n13 0.543603
R73 VTAIL.n6 VTAIL.n5 0.543603
R74 VTAIL.n5 VTAIL.n3 0.543603
R75 VTAIL.n2 VTAIL.n1 0.543603
R76 VTAIL VTAIL.n15 0.485414
R77 VTAIL.n11 VTAIL.n10 0.470328
R78 VTAIL.n3 VTAIL.n2 0.470328
R79 VTAIL VTAIL.n1 0.0586897
R80 B.n368 B.n367 585
R81 B.n369 B.n368 585
R82 B.n145 B.n56 585
R83 B.n144 B.n143 585
R84 B.n142 B.n141 585
R85 B.n140 B.n139 585
R86 B.n138 B.n137 585
R87 B.n136 B.n135 585
R88 B.n134 B.n133 585
R89 B.n132 B.n131 585
R90 B.n130 B.n129 585
R91 B.n128 B.n127 585
R92 B.n126 B.n125 585
R93 B.n124 B.n123 585
R94 B.n122 B.n121 585
R95 B.n120 B.n119 585
R96 B.n118 B.n117 585
R97 B.n116 B.n115 585
R98 B.n114 B.n113 585
R99 B.n112 B.n111 585
R100 B.n110 B.n109 585
R101 B.n108 B.n107 585
R102 B.n106 B.n105 585
R103 B.n104 B.n103 585
R104 B.n102 B.n101 585
R105 B.n100 B.n99 585
R106 B.n98 B.n97 585
R107 B.n95 B.n94 585
R108 B.n93 B.n92 585
R109 B.n91 B.n90 585
R110 B.n89 B.n88 585
R111 B.n87 B.n86 585
R112 B.n85 B.n84 585
R113 B.n83 B.n82 585
R114 B.n81 B.n80 585
R115 B.n79 B.n78 585
R116 B.n77 B.n76 585
R117 B.n75 B.n74 585
R118 B.n73 B.n72 585
R119 B.n71 B.n70 585
R120 B.n69 B.n68 585
R121 B.n67 B.n66 585
R122 B.n65 B.n64 585
R123 B.n63 B.n62 585
R124 B.n366 B.n34 585
R125 B.n370 B.n34 585
R126 B.n365 B.n33 585
R127 B.n371 B.n33 585
R128 B.n364 B.n363 585
R129 B.n363 B.n29 585
R130 B.n362 B.n28 585
R131 B.n377 B.n28 585
R132 B.n361 B.n27 585
R133 B.n378 B.n27 585
R134 B.n360 B.n26 585
R135 B.n379 B.n26 585
R136 B.n359 B.n358 585
R137 B.n358 B.n22 585
R138 B.n357 B.n21 585
R139 B.n385 B.n21 585
R140 B.n356 B.n20 585
R141 B.n386 B.n20 585
R142 B.n355 B.n19 585
R143 B.n387 B.n19 585
R144 B.n354 B.n353 585
R145 B.n353 B.n15 585
R146 B.n352 B.n14 585
R147 B.n393 B.n14 585
R148 B.n351 B.n13 585
R149 B.n394 B.n13 585
R150 B.n350 B.n12 585
R151 B.n395 B.n12 585
R152 B.n349 B.n348 585
R153 B.n348 B.n347 585
R154 B.n346 B.n345 585
R155 B.n346 B.n8 585
R156 B.n344 B.n7 585
R157 B.n402 B.n7 585
R158 B.n343 B.n6 585
R159 B.n403 B.n6 585
R160 B.n342 B.n5 585
R161 B.n404 B.n5 585
R162 B.n341 B.n340 585
R163 B.n340 B.n4 585
R164 B.n339 B.n146 585
R165 B.n339 B.n338 585
R166 B.n328 B.n147 585
R167 B.n331 B.n147 585
R168 B.n330 B.n329 585
R169 B.n332 B.n330 585
R170 B.n327 B.n152 585
R171 B.n152 B.n151 585
R172 B.n326 B.n325 585
R173 B.n325 B.n324 585
R174 B.n154 B.n153 585
R175 B.n155 B.n154 585
R176 B.n317 B.n316 585
R177 B.n318 B.n317 585
R178 B.n315 B.n160 585
R179 B.n160 B.n159 585
R180 B.n314 B.n313 585
R181 B.n313 B.n312 585
R182 B.n162 B.n161 585
R183 B.n163 B.n162 585
R184 B.n305 B.n304 585
R185 B.n306 B.n305 585
R186 B.n303 B.n167 585
R187 B.n171 B.n167 585
R188 B.n302 B.n301 585
R189 B.n301 B.n300 585
R190 B.n169 B.n168 585
R191 B.n170 B.n169 585
R192 B.n293 B.n292 585
R193 B.n294 B.n293 585
R194 B.n291 B.n176 585
R195 B.n176 B.n175 585
R196 B.n285 B.n284 585
R197 B.n283 B.n199 585
R198 B.n282 B.n198 585
R199 B.n287 B.n198 585
R200 B.n281 B.n280 585
R201 B.n279 B.n278 585
R202 B.n277 B.n276 585
R203 B.n275 B.n274 585
R204 B.n273 B.n272 585
R205 B.n271 B.n270 585
R206 B.n269 B.n268 585
R207 B.n267 B.n266 585
R208 B.n265 B.n264 585
R209 B.n263 B.n262 585
R210 B.n261 B.n260 585
R211 B.n259 B.n258 585
R212 B.n257 B.n256 585
R213 B.n255 B.n254 585
R214 B.n253 B.n252 585
R215 B.n251 B.n250 585
R216 B.n249 B.n248 585
R217 B.n247 B.n246 585
R218 B.n245 B.n244 585
R219 B.n243 B.n242 585
R220 B.n241 B.n240 585
R221 B.n239 B.n238 585
R222 B.n237 B.n236 585
R223 B.n234 B.n233 585
R224 B.n232 B.n231 585
R225 B.n230 B.n229 585
R226 B.n228 B.n227 585
R227 B.n226 B.n225 585
R228 B.n224 B.n223 585
R229 B.n222 B.n221 585
R230 B.n220 B.n219 585
R231 B.n218 B.n217 585
R232 B.n216 B.n215 585
R233 B.n214 B.n213 585
R234 B.n212 B.n211 585
R235 B.n210 B.n209 585
R236 B.n208 B.n207 585
R237 B.n206 B.n205 585
R238 B.n178 B.n177 585
R239 B.n290 B.n289 585
R240 B.n174 B.n173 585
R241 B.n175 B.n174 585
R242 B.n296 B.n295 585
R243 B.n295 B.n294 585
R244 B.n297 B.n172 585
R245 B.n172 B.n170 585
R246 B.n299 B.n298 585
R247 B.n300 B.n299 585
R248 B.n166 B.n165 585
R249 B.n171 B.n166 585
R250 B.n308 B.n307 585
R251 B.n307 B.n306 585
R252 B.n309 B.n164 585
R253 B.n164 B.n163 585
R254 B.n311 B.n310 585
R255 B.n312 B.n311 585
R256 B.n158 B.n157 585
R257 B.n159 B.n158 585
R258 B.n320 B.n319 585
R259 B.n319 B.n318 585
R260 B.n321 B.n156 585
R261 B.n156 B.n155 585
R262 B.n323 B.n322 585
R263 B.n324 B.n323 585
R264 B.n150 B.n149 585
R265 B.n151 B.n150 585
R266 B.n334 B.n333 585
R267 B.n333 B.n332 585
R268 B.n335 B.n148 585
R269 B.n331 B.n148 585
R270 B.n337 B.n336 585
R271 B.n338 B.n337 585
R272 B.n3 B.n0 585
R273 B.n4 B.n3 585
R274 B.n401 B.n1 585
R275 B.n402 B.n401 585
R276 B.n400 B.n399 585
R277 B.n400 B.n8 585
R278 B.n398 B.n9 585
R279 B.n347 B.n9 585
R280 B.n397 B.n396 585
R281 B.n396 B.n395 585
R282 B.n11 B.n10 585
R283 B.n394 B.n11 585
R284 B.n392 B.n391 585
R285 B.n393 B.n392 585
R286 B.n390 B.n16 585
R287 B.n16 B.n15 585
R288 B.n389 B.n388 585
R289 B.n388 B.n387 585
R290 B.n18 B.n17 585
R291 B.n386 B.n18 585
R292 B.n384 B.n383 585
R293 B.n385 B.n384 585
R294 B.n382 B.n23 585
R295 B.n23 B.n22 585
R296 B.n381 B.n380 585
R297 B.n380 B.n379 585
R298 B.n25 B.n24 585
R299 B.n378 B.n25 585
R300 B.n376 B.n375 585
R301 B.n377 B.n376 585
R302 B.n374 B.n30 585
R303 B.n30 B.n29 585
R304 B.n373 B.n372 585
R305 B.n372 B.n371 585
R306 B.n32 B.n31 585
R307 B.n370 B.n32 585
R308 B.n405 B.n404 585
R309 B.n403 B.n2 585
R310 B.n60 B.t8 496.63
R311 B.n57 B.t12 496.63
R312 B.n203 B.t15 496.63
R313 B.n200 B.t19 496.63
R314 B.n62 B.n32 458.866
R315 B.n368 B.n34 458.866
R316 B.n289 B.n176 458.866
R317 B.n285 B.n174 458.866
R318 B.n369 B.n55 256.663
R319 B.n369 B.n54 256.663
R320 B.n369 B.n53 256.663
R321 B.n369 B.n52 256.663
R322 B.n369 B.n51 256.663
R323 B.n369 B.n50 256.663
R324 B.n369 B.n49 256.663
R325 B.n369 B.n48 256.663
R326 B.n369 B.n47 256.663
R327 B.n369 B.n46 256.663
R328 B.n369 B.n45 256.663
R329 B.n369 B.n44 256.663
R330 B.n369 B.n43 256.663
R331 B.n369 B.n42 256.663
R332 B.n369 B.n41 256.663
R333 B.n369 B.n40 256.663
R334 B.n369 B.n39 256.663
R335 B.n369 B.n38 256.663
R336 B.n369 B.n37 256.663
R337 B.n369 B.n36 256.663
R338 B.n369 B.n35 256.663
R339 B.n287 B.n286 256.663
R340 B.n287 B.n179 256.663
R341 B.n287 B.n180 256.663
R342 B.n287 B.n181 256.663
R343 B.n287 B.n182 256.663
R344 B.n287 B.n183 256.663
R345 B.n287 B.n184 256.663
R346 B.n287 B.n185 256.663
R347 B.n287 B.n186 256.663
R348 B.n287 B.n187 256.663
R349 B.n287 B.n188 256.663
R350 B.n287 B.n189 256.663
R351 B.n287 B.n190 256.663
R352 B.n287 B.n191 256.663
R353 B.n287 B.n192 256.663
R354 B.n287 B.n193 256.663
R355 B.n287 B.n194 256.663
R356 B.n287 B.n195 256.663
R357 B.n287 B.n196 256.663
R358 B.n287 B.n197 256.663
R359 B.n288 B.n287 256.663
R360 B.n407 B.n406 256.663
R361 B.n66 B.n65 163.367
R362 B.n70 B.n69 163.367
R363 B.n74 B.n73 163.367
R364 B.n78 B.n77 163.367
R365 B.n82 B.n81 163.367
R366 B.n86 B.n85 163.367
R367 B.n90 B.n89 163.367
R368 B.n94 B.n93 163.367
R369 B.n99 B.n98 163.367
R370 B.n103 B.n102 163.367
R371 B.n107 B.n106 163.367
R372 B.n111 B.n110 163.367
R373 B.n115 B.n114 163.367
R374 B.n119 B.n118 163.367
R375 B.n123 B.n122 163.367
R376 B.n127 B.n126 163.367
R377 B.n131 B.n130 163.367
R378 B.n135 B.n134 163.367
R379 B.n139 B.n138 163.367
R380 B.n143 B.n142 163.367
R381 B.n368 B.n56 163.367
R382 B.n293 B.n176 163.367
R383 B.n293 B.n169 163.367
R384 B.n301 B.n169 163.367
R385 B.n301 B.n167 163.367
R386 B.n305 B.n167 163.367
R387 B.n305 B.n162 163.367
R388 B.n313 B.n162 163.367
R389 B.n313 B.n160 163.367
R390 B.n317 B.n160 163.367
R391 B.n317 B.n154 163.367
R392 B.n325 B.n154 163.367
R393 B.n325 B.n152 163.367
R394 B.n330 B.n152 163.367
R395 B.n330 B.n147 163.367
R396 B.n339 B.n147 163.367
R397 B.n340 B.n339 163.367
R398 B.n340 B.n5 163.367
R399 B.n6 B.n5 163.367
R400 B.n7 B.n6 163.367
R401 B.n346 B.n7 163.367
R402 B.n348 B.n346 163.367
R403 B.n348 B.n12 163.367
R404 B.n13 B.n12 163.367
R405 B.n14 B.n13 163.367
R406 B.n353 B.n14 163.367
R407 B.n353 B.n19 163.367
R408 B.n20 B.n19 163.367
R409 B.n21 B.n20 163.367
R410 B.n358 B.n21 163.367
R411 B.n358 B.n26 163.367
R412 B.n27 B.n26 163.367
R413 B.n28 B.n27 163.367
R414 B.n363 B.n28 163.367
R415 B.n363 B.n33 163.367
R416 B.n34 B.n33 163.367
R417 B.n199 B.n198 163.367
R418 B.n280 B.n198 163.367
R419 B.n278 B.n277 163.367
R420 B.n274 B.n273 163.367
R421 B.n270 B.n269 163.367
R422 B.n266 B.n265 163.367
R423 B.n262 B.n261 163.367
R424 B.n258 B.n257 163.367
R425 B.n254 B.n253 163.367
R426 B.n250 B.n249 163.367
R427 B.n246 B.n245 163.367
R428 B.n242 B.n241 163.367
R429 B.n238 B.n237 163.367
R430 B.n233 B.n232 163.367
R431 B.n229 B.n228 163.367
R432 B.n225 B.n224 163.367
R433 B.n221 B.n220 163.367
R434 B.n217 B.n216 163.367
R435 B.n213 B.n212 163.367
R436 B.n209 B.n208 163.367
R437 B.n205 B.n178 163.367
R438 B.n295 B.n174 163.367
R439 B.n295 B.n172 163.367
R440 B.n299 B.n172 163.367
R441 B.n299 B.n166 163.367
R442 B.n307 B.n166 163.367
R443 B.n307 B.n164 163.367
R444 B.n311 B.n164 163.367
R445 B.n311 B.n158 163.367
R446 B.n319 B.n158 163.367
R447 B.n319 B.n156 163.367
R448 B.n323 B.n156 163.367
R449 B.n323 B.n150 163.367
R450 B.n333 B.n150 163.367
R451 B.n333 B.n148 163.367
R452 B.n337 B.n148 163.367
R453 B.n337 B.n3 163.367
R454 B.n405 B.n3 163.367
R455 B.n401 B.n2 163.367
R456 B.n401 B.n400 163.367
R457 B.n400 B.n9 163.367
R458 B.n396 B.n9 163.367
R459 B.n396 B.n11 163.367
R460 B.n392 B.n11 163.367
R461 B.n392 B.n16 163.367
R462 B.n388 B.n16 163.367
R463 B.n388 B.n18 163.367
R464 B.n384 B.n18 163.367
R465 B.n384 B.n23 163.367
R466 B.n380 B.n23 163.367
R467 B.n380 B.n25 163.367
R468 B.n376 B.n25 163.367
R469 B.n376 B.n30 163.367
R470 B.n372 B.n30 163.367
R471 B.n372 B.n32 163.367
R472 B.n287 B.n175 144.325
R473 B.n370 B.n369 144.325
R474 B.n57 B.t13 86.5986
R475 B.n203 B.t18 86.5986
R476 B.n60 B.t10 86.5956
R477 B.n200 B.t21 86.5956
R478 B.n294 B.n175 85.3399
R479 B.n294 B.n170 85.3399
R480 B.n300 B.n170 85.3399
R481 B.n300 B.n171 85.3399
R482 B.n306 B.n163 85.3399
R483 B.n312 B.n163 85.3399
R484 B.n312 B.n159 85.3399
R485 B.n318 B.n159 85.3399
R486 B.n324 B.n155 85.3399
R487 B.n332 B.n151 85.3399
R488 B.n338 B.n4 85.3399
R489 B.n404 B.n4 85.3399
R490 B.n404 B.n403 85.3399
R491 B.n403 B.n402 85.3399
R492 B.n402 B.n8 85.3399
R493 B.n395 B.n394 85.3399
R494 B.n393 B.n15 85.3399
R495 B.n387 B.n386 85.3399
R496 B.n386 B.n385 85.3399
R497 B.n385 B.n22 85.3399
R498 B.n379 B.n22 85.3399
R499 B.n378 B.n377 85.3399
R500 B.n377 B.n29 85.3399
R501 B.n371 B.n29 85.3399
R502 B.n371 B.n370 85.3399
R503 B.n331 B.t1 82.8299
R504 B.n347 B.t3 82.8299
R505 B.t5 B.n331 75.3
R506 B.n347 B.t7 75.3
R507 B.n58 B.t14 74.3804
R508 B.n204 B.t17 74.3804
R509 B.n61 B.t11 74.3775
R510 B.n201 B.t20 74.3775
R511 B.n62 B.n35 71.676
R512 B.n66 B.n36 71.676
R513 B.n70 B.n37 71.676
R514 B.n74 B.n38 71.676
R515 B.n78 B.n39 71.676
R516 B.n82 B.n40 71.676
R517 B.n86 B.n41 71.676
R518 B.n90 B.n42 71.676
R519 B.n94 B.n43 71.676
R520 B.n99 B.n44 71.676
R521 B.n103 B.n45 71.676
R522 B.n107 B.n46 71.676
R523 B.n111 B.n47 71.676
R524 B.n115 B.n48 71.676
R525 B.n119 B.n49 71.676
R526 B.n123 B.n50 71.676
R527 B.n127 B.n51 71.676
R528 B.n131 B.n52 71.676
R529 B.n135 B.n53 71.676
R530 B.n139 B.n54 71.676
R531 B.n143 B.n55 71.676
R532 B.n56 B.n55 71.676
R533 B.n142 B.n54 71.676
R534 B.n138 B.n53 71.676
R535 B.n134 B.n52 71.676
R536 B.n130 B.n51 71.676
R537 B.n126 B.n50 71.676
R538 B.n122 B.n49 71.676
R539 B.n118 B.n48 71.676
R540 B.n114 B.n47 71.676
R541 B.n110 B.n46 71.676
R542 B.n106 B.n45 71.676
R543 B.n102 B.n44 71.676
R544 B.n98 B.n43 71.676
R545 B.n93 B.n42 71.676
R546 B.n89 B.n41 71.676
R547 B.n85 B.n40 71.676
R548 B.n81 B.n39 71.676
R549 B.n77 B.n38 71.676
R550 B.n73 B.n37 71.676
R551 B.n69 B.n36 71.676
R552 B.n65 B.n35 71.676
R553 B.n286 B.n285 71.676
R554 B.n280 B.n179 71.676
R555 B.n277 B.n180 71.676
R556 B.n273 B.n181 71.676
R557 B.n269 B.n182 71.676
R558 B.n265 B.n183 71.676
R559 B.n261 B.n184 71.676
R560 B.n257 B.n185 71.676
R561 B.n253 B.n186 71.676
R562 B.n249 B.n187 71.676
R563 B.n245 B.n188 71.676
R564 B.n241 B.n189 71.676
R565 B.n237 B.n190 71.676
R566 B.n232 B.n191 71.676
R567 B.n228 B.n192 71.676
R568 B.n224 B.n193 71.676
R569 B.n220 B.n194 71.676
R570 B.n216 B.n195 71.676
R571 B.n212 B.n196 71.676
R572 B.n208 B.n197 71.676
R573 B.n288 B.n178 71.676
R574 B.n286 B.n199 71.676
R575 B.n278 B.n179 71.676
R576 B.n274 B.n180 71.676
R577 B.n270 B.n181 71.676
R578 B.n266 B.n182 71.676
R579 B.n262 B.n183 71.676
R580 B.n258 B.n184 71.676
R581 B.n254 B.n185 71.676
R582 B.n250 B.n186 71.676
R583 B.n246 B.n187 71.676
R584 B.n242 B.n188 71.676
R585 B.n238 B.n189 71.676
R586 B.n233 B.n190 71.676
R587 B.n229 B.n191 71.676
R588 B.n225 B.n192 71.676
R589 B.n221 B.n193 71.676
R590 B.n217 B.n194 71.676
R591 B.n213 B.n195 71.676
R592 B.n209 B.n196 71.676
R593 B.n205 B.n197 71.676
R594 B.n289 B.n288 71.676
R595 B.n406 B.n405 71.676
R596 B.n406 B.n2 71.676
R597 B.t6 B.n151 62.7501
R598 B.n394 B.t2 62.7501
R599 B.n96 B.n61 59.5399
R600 B.n59 B.n58 59.5399
R601 B.n235 B.n204 59.5399
R602 B.n202 B.n201 59.5399
R603 B.n306 B.t16 55.2201
R604 B.n379 B.t9 55.2201
R605 B.t4 B.n155 50.2002
R606 B.t0 B.n15 50.2002
R607 B.n318 B.t4 35.1403
R608 B.n387 B.t0 35.1403
R609 B.n171 B.t16 30.1203
R610 B.t9 B.n378 30.1203
R611 B.n284 B.n173 29.8151
R612 B.n291 B.n290 29.8151
R613 B.n367 B.n366 29.8151
R614 B.n63 B.n31 29.8151
R615 B.n324 B.t6 22.5903
R616 B.t2 B.n393 22.5903
R617 B B.n407 18.0485
R618 B.n61 B.n60 12.2187
R619 B.n58 B.n57 12.2187
R620 B.n204 B.n203 12.2187
R621 B.n201 B.n200 12.2187
R622 B.n296 B.n173 10.6151
R623 B.n297 B.n296 10.6151
R624 B.n298 B.n297 10.6151
R625 B.n298 B.n165 10.6151
R626 B.n308 B.n165 10.6151
R627 B.n309 B.n308 10.6151
R628 B.n310 B.n309 10.6151
R629 B.n310 B.n157 10.6151
R630 B.n320 B.n157 10.6151
R631 B.n321 B.n320 10.6151
R632 B.n322 B.n321 10.6151
R633 B.n322 B.n149 10.6151
R634 B.n334 B.n149 10.6151
R635 B.n335 B.n334 10.6151
R636 B.n336 B.n335 10.6151
R637 B.n336 B.n0 10.6151
R638 B.n284 B.n283 10.6151
R639 B.n283 B.n282 10.6151
R640 B.n282 B.n281 10.6151
R641 B.n281 B.n279 10.6151
R642 B.n279 B.n276 10.6151
R643 B.n276 B.n275 10.6151
R644 B.n275 B.n272 10.6151
R645 B.n272 B.n271 10.6151
R646 B.n271 B.n268 10.6151
R647 B.n268 B.n267 10.6151
R648 B.n267 B.n264 10.6151
R649 B.n264 B.n263 10.6151
R650 B.n263 B.n260 10.6151
R651 B.n260 B.n259 10.6151
R652 B.n259 B.n256 10.6151
R653 B.n256 B.n255 10.6151
R654 B.n252 B.n251 10.6151
R655 B.n251 B.n248 10.6151
R656 B.n248 B.n247 10.6151
R657 B.n247 B.n244 10.6151
R658 B.n244 B.n243 10.6151
R659 B.n243 B.n240 10.6151
R660 B.n240 B.n239 10.6151
R661 B.n239 B.n236 10.6151
R662 B.n234 B.n231 10.6151
R663 B.n231 B.n230 10.6151
R664 B.n230 B.n227 10.6151
R665 B.n227 B.n226 10.6151
R666 B.n226 B.n223 10.6151
R667 B.n223 B.n222 10.6151
R668 B.n222 B.n219 10.6151
R669 B.n219 B.n218 10.6151
R670 B.n218 B.n215 10.6151
R671 B.n215 B.n214 10.6151
R672 B.n214 B.n211 10.6151
R673 B.n211 B.n210 10.6151
R674 B.n210 B.n207 10.6151
R675 B.n207 B.n206 10.6151
R676 B.n206 B.n177 10.6151
R677 B.n290 B.n177 10.6151
R678 B.n292 B.n291 10.6151
R679 B.n292 B.n168 10.6151
R680 B.n302 B.n168 10.6151
R681 B.n303 B.n302 10.6151
R682 B.n304 B.n303 10.6151
R683 B.n304 B.n161 10.6151
R684 B.n314 B.n161 10.6151
R685 B.n315 B.n314 10.6151
R686 B.n316 B.n315 10.6151
R687 B.n316 B.n153 10.6151
R688 B.n326 B.n153 10.6151
R689 B.n327 B.n326 10.6151
R690 B.n329 B.n327 10.6151
R691 B.n329 B.n328 10.6151
R692 B.n328 B.n146 10.6151
R693 B.n341 B.n146 10.6151
R694 B.n342 B.n341 10.6151
R695 B.n343 B.n342 10.6151
R696 B.n344 B.n343 10.6151
R697 B.n345 B.n344 10.6151
R698 B.n349 B.n345 10.6151
R699 B.n350 B.n349 10.6151
R700 B.n351 B.n350 10.6151
R701 B.n352 B.n351 10.6151
R702 B.n354 B.n352 10.6151
R703 B.n355 B.n354 10.6151
R704 B.n356 B.n355 10.6151
R705 B.n357 B.n356 10.6151
R706 B.n359 B.n357 10.6151
R707 B.n360 B.n359 10.6151
R708 B.n361 B.n360 10.6151
R709 B.n362 B.n361 10.6151
R710 B.n364 B.n362 10.6151
R711 B.n365 B.n364 10.6151
R712 B.n366 B.n365 10.6151
R713 B.n399 B.n1 10.6151
R714 B.n399 B.n398 10.6151
R715 B.n398 B.n397 10.6151
R716 B.n397 B.n10 10.6151
R717 B.n391 B.n10 10.6151
R718 B.n391 B.n390 10.6151
R719 B.n390 B.n389 10.6151
R720 B.n389 B.n17 10.6151
R721 B.n383 B.n17 10.6151
R722 B.n383 B.n382 10.6151
R723 B.n382 B.n381 10.6151
R724 B.n381 B.n24 10.6151
R725 B.n375 B.n24 10.6151
R726 B.n375 B.n374 10.6151
R727 B.n374 B.n373 10.6151
R728 B.n373 B.n31 10.6151
R729 B.n64 B.n63 10.6151
R730 B.n67 B.n64 10.6151
R731 B.n68 B.n67 10.6151
R732 B.n71 B.n68 10.6151
R733 B.n72 B.n71 10.6151
R734 B.n75 B.n72 10.6151
R735 B.n76 B.n75 10.6151
R736 B.n79 B.n76 10.6151
R737 B.n80 B.n79 10.6151
R738 B.n83 B.n80 10.6151
R739 B.n84 B.n83 10.6151
R740 B.n87 B.n84 10.6151
R741 B.n88 B.n87 10.6151
R742 B.n91 B.n88 10.6151
R743 B.n92 B.n91 10.6151
R744 B.n95 B.n92 10.6151
R745 B.n100 B.n97 10.6151
R746 B.n101 B.n100 10.6151
R747 B.n104 B.n101 10.6151
R748 B.n105 B.n104 10.6151
R749 B.n108 B.n105 10.6151
R750 B.n109 B.n108 10.6151
R751 B.n112 B.n109 10.6151
R752 B.n113 B.n112 10.6151
R753 B.n117 B.n116 10.6151
R754 B.n120 B.n117 10.6151
R755 B.n121 B.n120 10.6151
R756 B.n124 B.n121 10.6151
R757 B.n125 B.n124 10.6151
R758 B.n128 B.n125 10.6151
R759 B.n129 B.n128 10.6151
R760 B.n132 B.n129 10.6151
R761 B.n133 B.n132 10.6151
R762 B.n136 B.n133 10.6151
R763 B.n137 B.n136 10.6151
R764 B.n140 B.n137 10.6151
R765 B.n141 B.n140 10.6151
R766 B.n144 B.n141 10.6151
R767 B.n145 B.n144 10.6151
R768 B.n367 B.n145 10.6151
R769 B.n332 B.t5 10.0404
R770 B.n395 B.t7 10.0404
R771 B.n407 B.n0 8.11757
R772 B.n407 B.n1 8.11757
R773 B.n252 B.n202 6.5566
R774 B.n236 B.n235 6.5566
R775 B.n97 B.n96 6.5566
R776 B.n113 B.n59 6.5566
R777 B.n255 B.n202 4.05904
R778 B.n235 B.n234 4.05904
R779 B.n96 B.n95 4.05904
R780 B.n116 B.n59 4.05904
R781 B.n338 B.t1 2.51048
R782 B.t3 B.n8 2.51048
R783 VN.n7 VN.t1 414.082
R784 VN.n2 VN.t4 414.082
R785 VN.n16 VN.t5 414.082
R786 VN.n11 VN.t6 414.082
R787 VN.n6 VN.t3 385.601
R788 VN.n1 VN.t2 385.601
R789 VN.n15 VN.t0 385.601
R790 VN.n10 VN.t7 385.601
R791 VN.n12 VN.n11 161.489
R792 VN.n3 VN.n2 161.489
R793 VN.n8 VN.n7 161.3
R794 VN.n17 VN.n16 161.3
R795 VN.n14 VN.n9 161.3
R796 VN.n13 VN.n12 161.3
R797 VN.n5 VN.n0 161.3
R798 VN.n4 VN.n3 161.3
R799 VN.n5 VN.n4 73.0308
R800 VN.n14 VN.n13 73.0308
R801 VN.n2 VN.n1 63.5369
R802 VN.n7 VN.n6 63.5369
R803 VN.n16 VN.n15 63.5369
R804 VN.n11 VN.n10 63.5369
R805 VN VN.n17 34.0706
R806 VN.n4 VN.n1 9.49444
R807 VN.n6 VN.n5 9.49444
R808 VN.n15 VN.n14 9.49444
R809 VN.n13 VN.n10 9.49444
R810 VN.n17 VN.n9 0.189894
R811 VN.n12 VN.n9 0.189894
R812 VN.n3 VN.n0 0.189894
R813 VN.n8 VN.n0 0.189894
R814 VN VN.n8 0.0516364
R815 VDD2.n2 VDD2.n1 75.7706
R816 VDD2.n2 VDD2.n0 75.7706
R817 VDD2 VDD2.n5 75.7678
R818 VDD2.n4 VDD2.n3 75.5546
R819 VDD2.n4 VDD2.n2 29.1679
R820 VDD2.n5 VDD2.t0 5.67385
R821 VDD2.n5 VDD2.t1 5.67385
R822 VDD2.n3 VDD2.t2 5.67385
R823 VDD2.n3 VDD2.t7 5.67385
R824 VDD2.n1 VDD2.t4 5.67385
R825 VDD2.n1 VDD2.t6 5.67385
R826 VDD2.n0 VDD2.t3 5.67385
R827 VDD2.n0 VDD2.t5 5.67385
R828 VDD2 VDD2.n4 0.330241
C0 VTAIL VDD1 6.03032f
C1 VDD2 VN 1.22066f
C2 VDD2 VP 0.279799f
C3 VP VN 3.28236f
C4 VDD2 VDD1 0.631433f
C5 VDD2 VTAIL 6.06932f
C6 VDD1 VN 0.15204f
C7 VDD1 VP 1.34778f
C8 VTAIL VN 1.20572f
C9 VTAIL VP 1.21983f
C10 VDD2 B 2.367347f
C11 VDD1 B 2.534059f
C12 VTAIL B 3.717475f
C13 VN B 5.39412f
C14 VP B 4.381881f
C15 VDD2.t3 B 0.072055f
C16 VDD2.t5 B 0.072055f
C17 VDD2.n0 B 0.553667f
C18 VDD2.t4 B 0.072055f
C19 VDD2.t6 B 0.072055f
C20 VDD2.n1 B 0.553667f
C21 VDD2.n2 B 1.47235f
C22 VDD2.t2 B 0.072055f
C23 VDD2.t7 B 0.072055f
C24 VDD2.n3 B 0.55288f
C25 VDD2.n4 B 1.51897f
C26 VDD2.t0 B 0.072055f
C27 VDD2.t1 B 0.072055f
C28 VDD2.n5 B 0.553648f
C29 VN.n0 B 0.031574f
C30 VN.t3 B 0.095387f
C31 VN.t2 B 0.095387f
C32 VN.n1 B 0.052206f
C33 VN.t4 B 0.098972f
C34 VN.n2 B 0.061571f
C35 VN.n3 B 0.066805f
C36 VN.n4 B 0.011739f
C37 VN.n5 B 0.011739f
C38 VN.n6 B 0.052206f
C39 VN.t1 B 0.098972f
C40 VN.n7 B 0.06153f
C41 VN.n8 B 0.024469f
C42 VN.n9 B 0.031574f
C43 VN.t5 B 0.098972f
C44 VN.t0 B 0.095387f
C45 VN.t7 B 0.095387f
C46 VN.n10 B 0.052206f
C47 VN.t6 B 0.098972f
C48 VN.n11 B 0.061571f
C49 VN.n12 B 0.066805f
C50 VN.n13 B 0.011739f
C51 VN.n14 B 0.011739f
C52 VN.n15 B 0.052206f
C53 VN.n16 B 0.06153f
C54 VN.n17 B 0.893921f
C55 VTAIL.t7 B 0.061171f
C56 VTAIL.t2 B 0.061171f
C57 VTAIL.n0 B 0.422649f
C58 VTAIL.n1 B 0.228667f
C59 VTAIL.t3 B 0.543044f
C60 VTAIL.n2 B 0.304522f
C61 VTAIL.t12 B 0.543044f
C62 VTAIL.n3 B 0.304522f
C63 VTAIL.t11 B 0.061171f
C64 VTAIL.t15 B 0.061171f
C65 VTAIL.n4 B 0.422649f
C66 VTAIL.n5 B 0.263323f
C67 VTAIL.t14 B 0.543044f
C68 VTAIL.n6 B 0.826076f
C69 VTAIL.t4 B 0.543047f
C70 VTAIL.n7 B 0.826072f
C71 VTAIL.t6 B 0.061171f
C72 VTAIL.t5 B 0.061171f
C73 VTAIL.n8 B 0.422651f
C74 VTAIL.n9 B 0.263321f
C75 VTAIL.t1 B 0.543047f
C76 VTAIL.n10 B 0.304518f
C77 VTAIL.t13 B 0.543047f
C78 VTAIL.n11 B 0.304518f
C79 VTAIL.t10 B 0.061171f
C80 VTAIL.t9 B 0.061171f
C81 VTAIL.n12 B 0.422651f
C82 VTAIL.n13 B 0.263321f
C83 VTAIL.t8 B 0.543044f
C84 VTAIL.n14 B 0.826076f
C85 VTAIL.t0 B 0.543044f
C86 VTAIL.n15 B 0.821917f
C87 VDD1.t2 B 0.06977f
C88 VDD1.t5 B 0.06977f
C89 VDD1.n0 B 0.53654f
C90 VDD1.t1 B 0.06977f
C91 VDD1.t4 B 0.06977f
C92 VDD1.n1 B 0.53611f
C93 VDD1.t0 B 0.06977f
C94 VDD1.t3 B 0.06977f
C95 VDD1.n2 B 0.53611f
C96 VDD1.n3 B 1.48023f
C97 VDD1.t6 B 0.06977f
C98 VDD1.t7 B 0.06977f
C99 VDD1.n4 B 0.535345f
C100 VDD1.n5 B 1.50018f
C101 VP.n0 B 0.032005f
C102 VP.t0 B 0.096688f
C103 VP.t4 B 0.096688f
C104 VP.n1 B 0.052918f
C105 VP.n2 B 0.032005f
C106 VP.t6 B 0.096688f
C107 VP.t5 B 0.096688f
C108 VP.n3 B 0.052918f
C109 VP.t2 B 0.100321f
C110 VP.n4 B 0.06241f
C111 VP.n5 B 0.067716f
C112 VP.n6 B 0.0119f
C113 VP.n7 B 0.0119f
C114 VP.n8 B 0.052918f
C115 VP.t7 B 0.100321f
C116 VP.n9 B 0.062369f
C117 VP.n10 B 0.884773f
C118 VP.t1 B 0.100321f
C119 VP.n11 B 0.062369f
C120 VP.n12 B 0.918922f
C121 VP.n13 B 0.032005f
C122 VP.n14 B 0.0119f
C123 VP.n15 B 0.0119f
C124 VP.n16 B 0.052918f
C125 VP.t3 B 0.100321f
C126 VP.n17 B 0.062369f
C127 VP.n18 B 0.024802f
.ends

