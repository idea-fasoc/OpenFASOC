* NGSPICE file created from diff_pair_sample_1168.ext - technology: sky130A

.subckt diff_pair_sample_1168 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=6.2946 pd=33.06 as=6.2946 ps=33.06 w=16.14 l=3.24
X1 B.t15 B.t13 B.t14 B.t3 sky130_fd_pr__nfet_01v8 ad=6.2946 pd=33.06 as=0 ps=0 w=16.14 l=3.24
X2 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=6.2946 pd=33.06 as=0 ps=0 w=16.14 l=3.24
X3 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=6.2946 pd=33.06 as=0 ps=0 w=16.14 l=3.24
X4 VDD1.t0 VP.t1 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=6.2946 pd=33.06 as=6.2946 ps=33.06 w=16.14 l=3.24
X5 VDD2.t1 VN.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=6.2946 pd=33.06 as=6.2946 ps=33.06 w=16.14 l=3.24
X6 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=6.2946 pd=33.06 as=0 ps=0 w=16.14 l=3.24
X7 VDD2.t0 VN.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=6.2946 pd=33.06 as=6.2946 ps=33.06 w=16.14 l=3.24
R0 VP.n0 VP.t0 208.389
R1 VP.n0 VP.t1 158.899
R2 VP VP.n0 0.526373
R3 VTAIL.n354 VTAIL.n270 289.615
R4 VTAIL.n84 VTAIL.n0 289.615
R5 VTAIL.n264 VTAIL.n180 289.615
R6 VTAIL.n174 VTAIL.n90 289.615
R7 VTAIL.n298 VTAIL.n297 185
R8 VTAIL.n303 VTAIL.n302 185
R9 VTAIL.n305 VTAIL.n304 185
R10 VTAIL.n294 VTAIL.n293 185
R11 VTAIL.n311 VTAIL.n310 185
R12 VTAIL.n313 VTAIL.n312 185
R13 VTAIL.n290 VTAIL.n289 185
R14 VTAIL.n319 VTAIL.n318 185
R15 VTAIL.n321 VTAIL.n320 185
R16 VTAIL.n286 VTAIL.n285 185
R17 VTAIL.n327 VTAIL.n326 185
R18 VTAIL.n329 VTAIL.n328 185
R19 VTAIL.n282 VTAIL.n281 185
R20 VTAIL.n335 VTAIL.n334 185
R21 VTAIL.n337 VTAIL.n336 185
R22 VTAIL.n278 VTAIL.n277 185
R23 VTAIL.n344 VTAIL.n343 185
R24 VTAIL.n345 VTAIL.n276 185
R25 VTAIL.n347 VTAIL.n346 185
R26 VTAIL.n274 VTAIL.n273 185
R27 VTAIL.n353 VTAIL.n352 185
R28 VTAIL.n355 VTAIL.n354 185
R29 VTAIL.n28 VTAIL.n27 185
R30 VTAIL.n33 VTAIL.n32 185
R31 VTAIL.n35 VTAIL.n34 185
R32 VTAIL.n24 VTAIL.n23 185
R33 VTAIL.n41 VTAIL.n40 185
R34 VTAIL.n43 VTAIL.n42 185
R35 VTAIL.n20 VTAIL.n19 185
R36 VTAIL.n49 VTAIL.n48 185
R37 VTAIL.n51 VTAIL.n50 185
R38 VTAIL.n16 VTAIL.n15 185
R39 VTAIL.n57 VTAIL.n56 185
R40 VTAIL.n59 VTAIL.n58 185
R41 VTAIL.n12 VTAIL.n11 185
R42 VTAIL.n65 VTAIL.n64 185
R43 VTAIL.n67 VTAIL.n66 185
R44 VTAIL.n8 VTAIL.n7 185
R45 VTAIL.n74 VTAIL.n73 185
R46 VTAIL.n75 VTAIL.n6 185
R47 VTAIL.n77 VTAIL.n76 185
R48 VTAIL.n4 VTAIL.n3 185
R49 VTAIL.n83 VTAIL.n82 185
R50 VTAIL.n85 VTAIL.n84 185
R51 VTAIL.n265 VTAIL.n264 185
R52 VTAIL.n263 VTAIL.n262 185
R53 VTAIL.n184 VTAIL.n183 185
R54 VTAIL.n257 VTAIL.n256 185
R55 VTAIL.n255 VTAIL.n186 185
R56 VTAIL.n254 VTAIL.n253 185
R57 VTAIL.n189 VTAIL.n187 185
R58 VTAIL.n248 VTAIL.n247 185
R59 VTAIL.n246 VTAIL.n245 185
R60 VTAIL.n193 VTAIL.n192 185
R61 VTAIL.n240 VTAIL.n239 185
R62 VTAIL.n238 VTAIL.n237 185
R63 VTAIL.n197 VTAIL.n196 185
R64 VTAIL.n232 VTAIL.n231 185
R65 VTAIL.n230 VTAIL.n229 185
R66 VTAIL.n201 VTAIL.n200 185
R67 VTAIL.n224 VTAIL.n223 185
R68 VTAIL.n222 VTAIL.n221 185
R69 VTAIL.n205 VTAIL.n204 185
R70 VTAIL.n216 VTAIL.n215 185
R71 VTAIL.n214 VTAIL.n213 185
R72 VTAIL.n209 VTAIL.n208 185
R73 VTAIL.n175 VTAIL.n174 185
R74 VTAIL.n173 VTAIL.n172 185
R75 VTAIL.n94 VTAIL.n93 185
R76 VTAIL.n167 VTAIL.n166 185
R77 VTAIL.n165 VTAIL.n96 185
R78 VTAIL.n164 VTAIL.n163 185
R79 VTAIL.n99 VTAIL.n97 185
R80 VTAIL.n158 VTAIL.n157 185
R81 VTAIL.n156 VTAIL.n155 185
R82 VTAIL.n103 VTAIL.n102 185
R83 VTAIL.n150 VTAIL.n149 185
R84 VTAIL.n148 VTAIL.n147 185
R85 VTAIL.n107 VTAIL.n106 185
R86 VTAIL.n142 VTAIL.n141 185
R87 VTAIL.n140 VTAIL.n139 185
R88 VTAIL.n111 VTAIL.n110 185
R89 VTAIL.n134 VTAIL.n133 185
R90 VTAIL.n132 VTAIL.n131 185
R91 VTAIL.n115 VTAIL.n114 185
R92 VTAIL.n126 VTAIL.n125 185
R93 VTAIL.n124 VTAIL.n123 185
R94 VTAIL.n119 VTAIL.n118 185
R95 VTAIL.n299 VTAIL.t0 147.659
R96 VTAIL.n29 VTAIL.t2 147.659
R97 VTAIL.n210 VTAIL.t3 147.659
R98 VTAIL.n120 VTAIL.t1 147.659
R99 VTAIL.n303 VTAIL.n297 104.615
R100 VTAIL.n304 VTAIL.n303 104.615
R101 VTAIL.n304 VTAIL.n293 104.615
R102 VTAIL.n311 VTAIL.n293 104.615
R103 VTAIL.n312 VTAIL.n311 104.615
R104 VTAIL.n312 VTAIL.n289 104.615
R105 VTAIL.n319 VTAIL.n289 104.615
R106 VTAIL.n320 VTAIL.n319 104.615
R107 VTAIL.n320 VTAIL.n285 104.615
R108 VTAIL.n327 VTAIL.n285 104.615
R109 VTAIL.n328 VTAIL.n327 104.615
R110 VTAIL.n328 VTAIL.n281 104.615
R111 VTAIL.n335 VTAIL.n281 104.615
R112 VTAIL.n336 VTAIL.n335 104.615
R113 VTAIL.n336 VTAIL.n277 104.615
R114 VTAIL.n344 VTAIL.n277 104.615
R115 VTAIL.n345 VTAIL.n344 104.615
R116 VTAIL.n346 VTAIL.n345 104.615
R117 VTAIL.n346 VTAIL.n273 104.615
R118 VTAIL.n353 VTAIL.n273 104.615
R119 VTAIL.n354 VTAIL.n353 104.615
R120 VTAIL.n33 VTAIL.n27 104.615
R121 VTAIL.n34 VTAIL.n33 104.615
R122 VTAIL.n34 VTAIL.n23 104.615
R123 VTAIL.n41 VTAIL.n23 104.615
R124 VTAIL.n42 VTAIL.n41 104.615
R125 VTAIL.n42 VTAIL.n19 104.615
R126 VTAIL.n49 VTAIL.n19 104.615
R127 VTAIL.n50 VTAIL.n49 104.615
R128 VTAIL.n50 VTAIL.n15 104.615
R129 VTAIL.n57 VTAIL.n15 104.615
R130 VTAIL.n58 VTAIL.n57 104.615
R131 VTAIL.n58 VTAIL.n11 104.615
R132 VTAIL.n65 VTAIL.n11 104.615
R133 VTAIL.n66 VTAIL.n65 104.615
R134 VTAIL.n66 VTAIL.n7 104.615
R135 VTAIL.n74 VTAIL.n7 104.615
R136 VTAIL.n75 VTAIL.n74 104.615
R137 VTAIL.n76 VTAIL.n75 104.615
R138 VTAIL.n76 VTAIL.n3 104.615
R139 VTAIL.n83 VTAIL.n3 104.615
R140 VTAIL.n84 VTAIL.n83 104.615
R141 VTAIL.n264 VTAIL.n263 104.615
R142 VTAIL.n263 VTAIL.n183 104.615
R143 VTAIL.n256 VTAIL.n183 104.615
R144 VTAIL.n256 VTAIL.n255 104.615
R145 VTAIL.n255 VTAIL.n254 104.615
R146 VTAIL.n254 VTAIL.n187 104.615
R147 VTAIL.n247 VTAIL.n187 104.615
R148 VTAIL.n247 VTAIL.n246 104.615
R149 VTAIL.n246 VTAIL.n192 104.615
R150 VTAIL.n239 VTAIL.n192 104.615
R151 VTAIL.n239 VTAIL.n238 104.615
R152 VTAIL.n238 VTAIL.n196 104.615
R153 VTAIL.n231 VTAIL.n196 104.615
R154 VTAIL.n231 VTAIL.n230 104.615
R155 VTAIL.n230 VTAIL.n200 104.615
R156 VTAIL.n223 VTAIL.n200 104.615
R157 VTAIL.n223 VTAIL.n222 104.615
R158 VTAIL.n222 VTAIL.n204 104.615
R159 VTAIL.n215 VTAIL.n204 104.615
R160 VTAIL.n215 VTAIL.n214 104.615
R161 VTAIL.n214 VTAIL.n208 104.615
R162 VTAIL.n174 VTAIL.n173 104.615
R163 VTAIL.n173 VTAIL.n93 104.615
R164 VTAIL.n166 VTAIL.n93 104.615
R165 VTAIL.n166 VTAIL.n165 104.615
R166 VTAIL.n165 VTAIL.n164 104.615
R167 VTAIL.n164 VTAIL.n97 104.615
R168 VTAIL.n157 VTAIL.n97 104.615
R169 VTAIL.n157 VTAIL.n156 104.615
R170 VTAIL.n156 VTAIL.n102 104.615
R171 VTAIL.n149 VTAIL.n102 104.615
R172 VTAIL.n149 VTAIL.n148 104.615
R173 VTAIL.n148 VTAIL.n106 104.615
R174 VTAIL.n141 VTAIL.n106 104.615
R175 VTAIL.n141 VTAIL.n140 104.615
R176 VTAIL.n140 VTAIL.n110 104.615
R177 VTAIL.n133 VTAIL.n110 104.615
R178 VTAIL.n133 VTAIL.n132 104.615
R179 VTAIL.n132 VTAIL.n114 104.615
R180 VTAIL.n125 VTAIL.n114 104.615
R181 VTAIL.n125 VTAIL.n124 104.615
R182 VTAIL.n124 VTAIL.n118 104.615
R183 VTAIL.t0 VTAIL.n297 52.3082
R184 VTAIL.t2 VTAIL.n27 52.3082
R185 VTAIL.t3 VTAIL.n208 52.3082
R186 VTAIL.t1 VTAIL.n118 52.3082
R187 VTAIL.n359 VTAIL.n358 33.349
R188 VTAIL.n89 VTAIL.n88 33.349
R189 VTAIL.n269 VTAIL.n268 33.349
R190 VTAIL.n179 VTAIL.n178 33.349
R191 VTAIL.n179 VTAIL.n89 32.4358
R192 VTAIL.n359 VTAIL.n269 29.3583
R193 VTAIL.n299 VTAIL.n298 15.6677
R194 VTAIL.n29 VTAIL.n28 15.6677
R195 VTAIL.n210 VTAIL.n209 15.6677
R196 VTAIL.n120 VTAIL.n119 15.6677
R197 VTAIL.n347 VTAIL.n276 13.1884
R198 VTAIL.n77 VTAIL.n6 13.1884
R199 VTAIL.n257 VTAIL.n186 13.1884
R200 VTAIL.n167 VTAIL.n96 13.1884
R201 VTAIL.n302 VTAIL.n301 12.8005
R202 VTAIL.n343 VTAIL.n342 12.8005
R203 VTAIL.n348 VTAIL.n274 12.8005
R204 VTAIL.n32 VTAIL.n31 12.8005
R205 VTAIL.n73 VTAIL.n72 12.8005
R206 VTAIL.n78 VTAIL.n4 12.8005
R207 VTAIL.n258 VTAIL.n184 12.8005
R208 VTAIL.n253 VTAIL.n188 12.8005
R209 VTAIL.n213 VTAIL.n212 12.8005
R210 VTAIL.n168 VTAIL.n94 12.8005
R211 VTAIL.n163 VTAIL.n98 12.8005
R212 VTAIL.n123 VTAIL.n122 12.8005
R213 VTAIL.n305 VTAIL.n296 12.0247
R214 VTAIL.n341 VTAIL.n278 12.0247
R215 VTAIL.n352 VTAIL.n351 12.0247
R216 VTAIL.n35 VTAIL.n26 12.0247
R217 VTAIL.n71 VTAIL.n8 12.0247
R218 VTAIL.n82 VTAIL.n81 12.0247
R219 VTAIL.n262 VTAIL.n261 12.0247
R220 VTAIL.n252 VTAIL.n189 12.0247
R221 VTAIL.n216 VTAIL.n207 12.0247
R222 VTAIL.n172 VTAIL.n171 12.0247
R223 VTAIL.n162 VTAIL.n99 12.0247
R224 VTAIL.n126 VTAIL.n117 12.0247
R225 VTAIL.n306 VTAIL.n294 11.249
R226 VTAIL.n338 VTAIL.n337 11.249
R227 VTAIL.n355 VTAIL.n272 11.249
R228 VTAIL.n36 VTAIL.n24 11.249
R229 VTAIL.n68 VTAIL.n67 11.249
R230 VTAIL.n85 VTAIL.n2 11.249
R231 VTAIL.n265 VTAIL.n182 11.249
R232 VTAIL.n249 VTAIL.n248 11.249
R233 VTAIL.n217 VTAIL.n205 11.249
R234 VTAIL.n175 VTAIL.n92 11.249
R235 VTAIL.n159 VTAIL.n158 11.249
R236 VTAIL.n127 VTAIL.n115 11.249
R237 VTAIL.n310 VTAIL.n309 10.4732
R238 VTAIL.n334 VTAIL.n280 10.4732
R239 VTAIL.n356 VTAIL.n270 10.4732
R240 VTAIL.n40 VTAIL.n39 10.4732
R241 VTAIL.n64 VTAIL.n10 10.4732
R242 VTAIL.n86 VTAIL.n0 10.4732
R243 VTAIL.n266 VTAIL.n180 10.4732
R244 VTAIL.n245 VTAIL.n191 10.4732
R245 VTAIL.n221 VTAIL.n220 10.4732
R246 VTAIL.n176 VTAIL.n90 10.4732
R247 VTAIL.n155 VTAIL.n101 10.4732
R248 VTAIL.n131 VTAIL.n130 10.4732
R249 VTAIL.n313 VTAIL.n292 9.69747
R250 VTAIL.n333 VTAIL.n282 9.69747
R251 VTAIL.n43 VTAIL.n22 9.69747
R252 VTAIL.n63 VTAIL.n12 9.69747
R253 VTAIL.n244 VTAIL.n193 9.69747
R254 VTAIL.n224 VTAIL.n203 9.69747
R255 VTAIL.n154 VTAIL.n103 9.69747
R256 VTAIL.n134 VTAIL.n113 9.69747
R257 VTAIL.n358 VTAIL.n357 9.45567
R258 VTAIL.n88 VTAIL.n87 9.45567
R259 VTAIL.n268 VTAIL.n267 9.45567
R260 VTAIL.n178 VTAIL.n177 9.45567
R261 VTAIL.n357 VTAIL.n356 9.3005
R262 VTAIL.n272 VTAIL.n271 9.3005
R263 VTAIL.n351 VTAIL.n350 9.3005
R264 VTAIL.n349 VTAIL.n348 9.3005
R265 VTAIL.n288 VTAIL.n287 9.3005
R266 VTAIL.n317 VTAIL.n316 9.3005
R267 VTAIL.n315 VTAIL.n314 9.3005
R268 VTAIL.n292 VTAIL.n291 9.3005
R269 VTAIL.n309 VTAIL.n308 9.3005
R270 VTAIL.n307 VTAIL.n306 9.3005
R271 VTAIL.n296 VTAIL.n295 9.3005
R272 VTAIL.n301 VTAIL.n300 9.3005
R273 VTAIL.n323 VTAIL.n322 9.3005
R274 VTAIL.n325 VTAIL.n324 9.3005
R275 VTAIL.n284 VTAIL.n283 9.3005
R276 VTAIL.n331 VTAIL.n330 9.3005
R277 VTAIL.n333 VTAIL.n332 9.3005
R278 VTAIL.n280 VTAIL.n279 9.3005
R279 VTAIL.n339 VTAIL.n338 9.3005
R280 VTAIL.n341 VTAIL.n340 9.3005
R281 VTAIL.n342 VTAIL.n275 9.3005
R282 VTAIL.n87 VTAIL.n86 9.3005
R283 VTAIL.n2 VTAIL.n1 9.3005
R284 VTAIL.n81 VTAIL.n80 9.3005
R285 VTAIL.n79 VTAIL.n78 9.3005
R286 VTAIL.n18 VTAIL.n17 9.3005
R287 VTAIL.n47 VTAIL.n46 9.3005
R288 VTAIL.n45 VTAIL.n44 9.3005
R289 VTAIL.n22 VTAIL.n21 9.3005
R290 VTAIL.n39 VTAIL.n38 9.3005
R291 VTAIL.n37 VTAIL.n36 9.3005
R292 VTAIL.n26 VTAIL.n25 9.3005
R293 VTAIL.n31 VTAIL.n30 9.3005
R294 VTAIL.n53 VTAIL.n52 9.3005
R295 VTAIL.n55 VTAIL.n54 9.3005
R296 VTAIL.n14 VTAIL.n13 9.3005
R297 VTAIL.n61 VTAIL.n60 9.3005
R298 VTAIL.n63 VTAIL.n62 9.3005
R299 VTAIL.n10 VTAIL.n9 9.3005
R300 VTAIL.n69 VTAIL.n68 9.3005
R301 VTAIL.n71 VTAIL.n70 9.3005
R302 VTAIL.n72 VTAIL.n5 9.3005
R303 VTAIL.n236 VTAIL.n235 9.3005
R304 VTAIL.n195 VTAIL.n194 9.3005
R305 VTAIL.n242 VTAIL.n241 9.3005
R306 VTAIL.n244 VTAIL.n243 9.3005
R307 VTAIL.n191 VTAIL.n190 9.3005
R308 VTAIL.n250 VTAIL.n249 9.3005
R309 VTAIL.n252 VTAIL.n251 9.3005
R310 VTAIL.n188 VTAIL.n185 9.3005
R311 VTAIL.n267 VTAIL.n266 9.3005
R312 VTAIL.n182 VTAIL.n181 9.3005
R313 VTAIL.n261 VTAIL.n260 9.3005
R314 VTAIL.n259 VTAIL.n258 9.3005
R315 VTAIL.n234 VTAIL.n233 9.3005
R316 VTAIL.n199 VTAIL.n198 9.3005
R317 VTAIL.n228 VTAIL.n227 9.3005
R318 VTAIL.n226 VTAIL.n225 9.3005
R319 VTAIL.n203 VTAIL.n202 9.3005
R320 VTAIL.n220 VTAIL.n219 9.3005
R321 VTAIL.n218 VTAIL.n217 9.3005
R322 VTAIL.n207 VTAIL.n206 9.3005
R323 VTAIL.n212 VTAIL.n211 9.3005
R324 VTAIL.n146 VTAIL.n145 9.3005
R325 VTAIL.n105 VTAIL.n104 9.3005
R326 VTAIL.n152 VTAIL.n151 9.3005
R327 VTAIL.n154 VTAIL.n153 9.3005
R328 VTAIL.n101 VTAIL.n100 9.3005
R329 VTAIL.n160 VTAIL.n159 9.3005
R330 VTAIL.n162 VTAIL.n161 9.3005
R331 VTAIL.n98 VTAIL.n95 9.3005
R332 VTAIL.n177 VTAIL.n176 9.3005
R333 VTAIL.n92 VTAIL.n91 9.3005
R334 VTAIL.n171 VTAIL.n170 9.3005
R335 VTAIL.n169 VTAIL.n168 9.3005
R336 VTAIL.n144 VTAIL.n143 9.3005
R337 VTAIL.n109 VTAIL.n108 9.3005
R338 VTAIL.n138 VTAIL.n137 9.3005
R339 VTAIL.n136 VTAIL.n135 9.3005
R340 VTAIL.n113 VTAIL.n112 9.3005
R341 VTAIL.n130 VTAIL.n129 9.3005
R342 VTAIL.n128 VTAIL.n127 9.3005
R343 VTAIL.n117 VTAIL.n116 9.3005
R344 VTAIL.n122 VTAIL.n121 9.3005
R345 VTAIL.n314 VTAIL.n290 8.92171
R346 VTAIL.n330 VTAIL.n329 8.92171
R347 VTAIL.n44 VTAIL.n20 8.92171
R348 VTAIL.n60 VTAIL.n59 8.92171
R349 VTAIL.n241 VTAIL.n240 8.92171
R350 VTAIL.n225 VTAIL.n201 8.92171
R351 VTAIL.n151 VTAIL.n150 8.92171
R352 VTAIL.n135 VTAIL.n111 8.92171
R353 VTAIL.n318 VTAIL.n317 8.14595
R354 VTAIL.n326 VTAIL.n284 8.14595
R355 VTAIL.n48 VTAIL.n47 8.14595
R356 VTAIL.n56 VTAIL.n14 8.14595
R357 VTAIL.n237 VTAIL.n195 8.14595
R358 VTAIL.n229 VTAIL.n228 8.14595
R359 VTAIL.n147 VTAIL.n105 8.14595
R360 VTAIL.n139 VTAIL.n138 8.14595
R361 VTAIL.n321 VTAIL.n288 7.3702
R362 VTAIL.n325 VTAIL.n286 7.3702
R363 VTAIL.n51 VTAIL.n18 7.3702
R364 VTAIL.n55 VTAIL.n16 7.3702
R365 VTAIL.n236 VTAIL.n197 7.3702
R366 VTAIL.n232 VTAIL.n199 7.3702
R367 VTAIL.n146 VTAIL.n107 7.3702
R368 VTAIL.n142 VTAIL.n109 7.3702
R369 VTAIL.n322 VTAIL.n321 6.59444
R370 VTAIL.n322 VTAIL.n286 6.59444
R371 VTAIL.n52 VTAIL.n51 6.59444
R372 VTAIL.n52 VTAIL.n16 6.59444
R373 VTAIL.n233 VTAIL.n197 6.59444
R374 VTAIL.n233 VTAIL.n232 6.59444
R375 VTAIL.n143 VTAIL.n107 6.59444
R376 VTAIL.n143 VTAIL.n142 6.59444
R377 VTAIL.n318 VTAIL.n288 5.81868
R378 VTAIL.n326 VTAIL.n325 5.81868
R379 VTAIL.n48 VTAIL.n18 5.81868
R380 VTAIL.n56 VTAIL.n55 5.81868
R381 VTAIL.n237 VTAIL.n236 5.81868
R382 VTAIL.n229 VTAIL.n199 5.81868
R383 VTAIL.n147 VTAIL.n146 5.81868
R384 VTAIL.n139 VTAIL.n109 5.81868
R385 VTAIL.n317 VTAIL.n290 5.04292
R386 VTAIL.n329 VTAIL.n284 5.04292
R387 VTAIL.n47 VTAIL.n20 5.04292
R388 VTAIL.n59 VTAIL.n14 5.04292
R389 VTAIL.n240 VTAIL.n195 5.04292
R390 VTAIL.n228 VTAIL.n201 5.04292
R391 VTAIL.n150 VTAIL.n105 5.04292
R392 VTAIL.n138 VTAIL.n111 5.04292
R393 VTAIL.n300 VTAIL.n299 4.38563
R394 VTAIL.n30 VTAIL.n29 4.38563
R395 VTAIL.n211 VTAIL.n210 4.38563
R396 VTAIL.n121 VTAIL.n120 4.38563
R397 VTAIL.n314 VTAIL.n313 4.26717
R398 VTAIL.n330 VTAIL.n282 4.26717
R399 VTAIL.n44 VTAIL.n43 4.26717
R400 VTAIL.n60 VTAIL.n12 4.26717
R401 VTAIL.n241 VTAIL.n193 4.26717
R402 VTAIL.n225 VTAIL.n224 4.26717
R403 VTAIL.n151 VTAIL.n103 4.26717
R404 VTAIL.n135 VTAIL.n134 4.26717
R405 VTAIL.n310 VTAIL.n292 3.49141
R406 VTAIL.n334 VTAIL.n333 3.49141
R407 VTAIL.n358 VTAIL.n270 3.49141
R408 VTAIL.n40 VTAIL.n22 3.49141
R409 VTAIL.n64 VTAIL.n63 3.49141
R410 VTAIL.n88 VTAIL.n0 3.49141
R411 VTAIL.n268 VTAIL.n180 3.49141
R412 VTAIL.n245 VTAIL.n244 3.49141
R413 VTAIL.n221 VTAIL.n203 3.49141
R414 VTAIL.n178 VTAIL.n90 3.49141
R415 VTAIL.n155 VTAIL.n154 3.49141
R416 VTAIL.n131 VTAIL.n113 3.49141
R417 VTAIL.n309 VTAIL.n294 2.71565
R418 VTAIL.n337 VTAIL.n280 2.71565
R419 VTAIL.n356 VTAIL.n355 2.71565
R420 VTAIL.n39 VTAIL.n24 2.71565
R421 VTAIL.n67 VTAIL.n10 2.71565
R422 VTAIL.n86 VTAIL.n85 2.71565
R423 VTAIL.n266 VTAIL.n265 2.71565
R424 VTAIL.n248 VTAIL.n191 2.71565
R425 VTAIL.n220 VTAIL.n205 2.71565
R426 VTAIL.n176 VTAIL.n175 2.71565
R427 VTAIL.n158 VTAIL.n101 2.71565
R428 VTAIL.n130 VTAIL.n115 2.71565
R429 VTAIL.n269 VTAIL.n179 2.00912
R430 VTAIL.n306 VTAIL.n305 1.93989
R431 VTAIL.n338 VTAIL.n278 1.93989
R432 VTAIL.n352 VTAIL.n272 1.93989
R433 VTAIL.n36 VTAIL.n35 1.93989
R434 VTAIL.n68 VTAIL.n8 1.93989
R435 VTAIL.n82 VTAIL.n2 1.93989
R436 VTAIL.n262 VTAIL.n182 1.93989
R437 VTAIL.n249 VTAIL.n189 1.93989
R438 VTAIL.n217 VTAIL.n216 1.93989
R439 VTAIL.n172 VTAIL.n92 1.93989
R440 VTAIL.n159 VTAIL.n99 1.93989
R441 VTAIL.n127 VTAIL.n126 1.93989
R442 VTAIL VTAIL.n89 1.29791
R443 VTAIL.n302 VTAIL.n296 1.16414
R444 VTAIL.n343 VTAIL.n341 1.16414
R445 VTAIL.n351 VTAIL.n274 1.16414
R446 VTAIL.n32 VTAIL.n26 1.16414
R447 VTAIL.n73 VTAIL.n71 1.16414
R448 VTAIL.n81 VTAIL.n4 1.16414
R449 VTAIL.n261 VTAIL.n184 1.16414
R450 VTAIL.n253 VTAIL.n252 1.16414
R451 VTAIL.n213 VTAIL.n207 1.16414
R452 VTAIL.n171 VTAIL.n94 1.16414
R453 VTAIL.n163 VTAIL.n162 1.16414
R454 VTAIL.n123 VTAIL.n117 1.16414
R455 VTAIL VTAIL.n359 0.711707
R456 VTAIL.n301 VTAIL.n298 0.388379
R457 VTAIL.n342 VTAIL.n276 0.388379
R458 VTAIL.n348 VTAIL.n347 0.388379
R459 VTAIL.n31 VTAIL.n28 0.388379
R460 VTAIL.n72 VTAIL.n6 0.388379
R461 VTAIL.n78 VTAIL.n77 0.388379
R462 VTAIL.n258 VTAIL.n257 0.388379
R463 VTAIL.n188 VTAIL.n186 0.388379
R464 VTAIL.n212 VTAIL.n209 0.388379
R465 VTAIL.n168 VTAIL.n167 0.388379
R466 VTAIL.n98 VTAIL.n96 0.388379
R467 VTAIL.n122 VTAIL.n119 0.388379
R468 VTAIL.n300 VTAIL.n295 0.155672
R469 VTAIL.n307 VTAIL.n295 0.155672
R470 VTAIL.n308 VTAIL.n307 0.155672
R471 VTAIL.n308 VTAIL.n291 0.155672
R472 VTAIL.n315 VTAIL.n291 0.155672
R473 VTAIL.n316 VTAIL.n315 0.155672
R474 VTAIL.n316 VTAIL.n287 0.155672
R475 VTAIL.n323 VTAIL.n287 0.155672
R476 VTAIL.n324 VTAIL.n323 0.155672
R477 VTAIL.n324 VTAIL.n283 0.155672
R478 VTAIL.n331 VTAIL.n283 0.155672
R479 VTAIL.n332 VTAIL.n331 0.155672
R480 VTAIL.n332 VTAIL.n279 0.155672
R481 VTAIL.n339 VTAIL.n279 0.155672
R482 VTAIL.n340 VTAIL.n339 0.155672
R483 VTAIL.n340 VTAIL.n275 0.155672
R484 VTAIL.n349 VTAIL.n275 0.155672
R485 VTAIL.n350 VTAIL.n349 0.155672
R486 VTAIL.n350 VTAIL.n271 0.155672
R487 VTAIL.n357 VTAIL.n271 0.155672
R488 VTAIL.n30 VTAIL.n25 0.155672
R489 VTAIL.n37 VTAIL.n25 0.155672
R490 VTAIL.n38 VTAIL.n37 0.155672
R491 VTAIL.n38 VTAIL.n21 0.155672
R492 VTAIL.n45 VTAIL.n21 0.155672
R493 VTAIL.n46 VTAIL.n45 0.155672
R494 VTAIL.n46 VTAIL.n17 0.155672
R495 VTAIL.n53 VTAIL.n17 0.155672
R496 VTAIL.n54 VTAIL.n53 0.155672
R497 VTAIL.n54 VTAIL.n13 0.155672
R498 VTAIL.n61 VTAIL.n13 0.155672
R499 VTAIL.n62 VTAIL.n61 0.155672
R500 VTAIL.n62 VTAIL.n9 0.155672
R501 VTAIL.n69 VTAIL.n9 0.155672
R502 VTAIL.n70 VTAIL.n69 0.155672
R503 VTAIL.n70 VTAIL.n5 0.155672
R504 VTAIL.n79 VTAIL.n5 0.155672
R505 VTAIL.n80 VTAIL.n79 0.155672
R506 VTAIL.n80 VTAIL.n1 0.155672
R507 VTAIL.n87 VTAIL.n1 0.155672
R508 VTAIL.n267 VTAIL.n181 0.155672
R509 VTAIL.n260 VTAIL.n181 0.155672
R510 VTAIL.n260 VTAIL.n259 0.155672
R511 VTAIL.n259 VTAIL.n185 0.155672
R512 VTAIL.n251 VTAIL.n185 0.155672
R513 VTAIL.n251 VTAIL.n250 0.155672
R514 VTAIL.n250 VTAIL.n190 0.155672
R515 VTAIL.n243 VTAIL.n190 0.155672
R516 VTAIL.n243 VTAIL.n242 0.155672
R517 VTAIL.n242 VTAIL.n194 0.155672
R518 VTAIL.n235 VTAIL.n194 0.155672
R519 VTAIL.n235 VTAIL.n234 0.155672
R520 VTAIL.n234 VTAIL.n198 0.155672
R521 VTAIL.n227 VTAIL.n198 0.155672
R522 VTAIL.n227 VTAIL.n226 0.155672
R523 VTAIL.n226 VTAIL.n202 0.155672
R524 VTAIL.n219 VTAIL.n202 0.155672
R525 VTAIL.n219 VTAIL.n218 0.155672
R526 VTAIL.n218 VTAIL.n206 0.155672
R527 VTAIL.n211 VTAIL.n206 0.155672
R528 VTAIL.n177 VTAIL.n91 0.155672
R529 VTAIL.n170 VTAIL.n91 0.155672
R530 VTAIL.n170 VTAIL.n169 0.155672
R531 VTAIL.n169 VTAIL.n95 0.155672
R532 VTAIL.n161 VTAIL.n95 0.155672
R533 VTAIL.n161 VTAIL.n160 0.155672
R534 VTAIL.n160 VTAIL.n100 0.155672
R535 VTAIL.n153 VTAIL.n100 0.155672
R536 VTAIL.n153 VTAIL.n152 0.155672
R537 VTAIL.n152 VTAIL.n104 0.155672
R538 VTAIL.n145 VTAIL.n104 0.155672
R539 VTAIL.n145 VTAIL.n144 0.155672
R540 VTAIL.n144 VTAIL.n108 0.155672
R541 VTAIL.n137 VTAIL.n108 0.155672
R542 VTAIL.n137 VTAIL.n136 0.155672
R543 VTAIL.n136 VTAIL.n112 0.155672
R544 VTAIL.n129 VTAIL.n112 0.155672
R545 VTAIL.n129 VTAIL.n128 0.155672
R546 VTAIL.n128 VTAIL.n116 0.155672
R547 VTAIL.n121 VTAIL.n116 0.155672
R548 VDD1.n84 VDD1.n0 289.615
R549 VDD1.n173 VDD1.n89 289.615
R550 VDD1.n85 VDD1.n84 185
R551 VDD1.n83 VDD1.n82 185
R552 VDD1.n4 VDD1.n3 185
R553 VDD1.n77 VDD1.n76 185
R554 VDD1.n75 VDD1.n6 185
R555 VDD1.n74 VDD1.n73 185
R556 VDD1.n9 VDD1.n7 185
R557 VDD1.n68 VDD1.n67 185
R558 VDD1.n66 VDD1.n65 185
R559 VDD1.n13 VDD1.n12 185
R560 VDD1.n60 VDD1.n59 185
R561 VDD1.n58 VDD1.n57 185
R562 VDD1.n17 VDD1.n16 185
R563 VDD1.n52 VDD1.n51 185
R564 VDD1.n50 VDD1.n49 185
R565 VDD1.n21 VDD1.n20 185
R566 VDD1.n44 VDD1.n43 185
R567 VDD1.n42 VDD1.n41 185
R568 VDD1.n25 VDD1.n24 185
R569 VDD1.n36 VDD1.n35 185
R570 VDD1.n34 VDD1.n33 185
R571 VDD1.n29 VDD1.n28 185
R572 VDD1.n117 VDD1.n116 185
R573 VDD1.n122 VDD1.n121 185
R574 VDD1.n124 VDD1.n123 185
R575 VDD1.n113 VDD1.n112 185
R576 VDD1.n130 VDD1.n129 185
R577 VDD1.n132 VDD1.n131 185
R578 VDD1.n109 VDD1.n108 185
R579 VDD1.n138 VDD1.n137 185
R580 VDD1.n140 VDD1.n139 185
R581 VDD1.n105 VDD1.n104 185
R582 VDD1.n146 VDD1.n145 185
R583 VDD1.n148 VDD1.n147 185
R584 VDD1.n101 VDD1.n100 185
R585 VDD1.n154 VDD1.n153 185
R586 VDD1.n156 VDD1.n155 185
R587 VDD1.n97 VDD1.n96 185
R588 VDD1.n163 VDD1.n162 185
R589 VDD1.n164 VDD1.n95 185
R590 VDD1.n166 VDD1.n165 185
R591 VDD1.n93 VDD1.n92 185
R592 VDD1.n172 VDD1.n171 185
R593 VDD1.n174 VDD1.n173 185
R594 VDD1.n30 VDD1.t1 147.659
R595 VDD1.n118 VDD1.t0 147.659
R596 VDD1.n84 VDD1.n83 104.615
R597 VDD1.n83 VDD1.n3 104.615
R598 VDD1.n76 VDD1.n3 104.615
R599 VDD1.n76 VDD1.n75 104.615
R600 VDD1.n75 VDD1.n74 104.615
R601 VDD1.n74 VDD1.n7 104.615
R602 VDD1.n67 VDD1.n7 104.615
R603 VDD1.n67 VDD1.n66 104.615
R604 VDD1.n66 VDD1.n12 104.615
R605 VDD1.n59 VDD1.n12 104.615
R606 VDD1.n59 VDD1.n58 104.615
R607 VDD1.n58 VDD1.n16 104.615
R608 VDD1.n51 VDD1.n16 104.615
R609 VDD1.n51 VDD1.n50 104.615
R610 VDD1.n50 VDD1.n20 104.615
R611 VDD1.n43 VDD1.n20 104.615
R612 VDD1.n43 VDD1.n42 104.615
R613 VDD1.n42 VDD1.n24 104.615
R614 VDD1.n35 VDD1.n24 104.615
R615 VDD1.n35 VDD1.n34 104.615
R616 VDD1.n34 VDD1.n28 104.615
R617 VDD1.n122 VDD1.n116 104.615
R618 VDD1.n123 VDD1.n122 104.615
R619 VDD1.n123 VDD1.n112 104.615
R620 VDD1.n130 VDD1.n112 104.615
R621 VDD1.n131 VDD1.n130 104.615
R622 VDD1.n131 VDD1.n108 104.615
R623 VDD1.n138 VDD1.n108 104.615
R624 VDD1.n139 VDD1.n138 104.615
R625 VDD1.n139 VDD1.n104 104.615
R626 VDD1.n146 VDD1.n104 104.615
R627 VDD1.n147 VDD1.n146 104.615
R628 VDD1.n147 VDD1.n100 104.615
R629 VDD1.n154 VDD1.n100 104.615
R630 VDD1.n155 VDD1.n154 104.615
R631 VDD1.n155 VDD1.n96 104.615
R632 VDD1.n163 VDD1.n96 104.615
R633 VDD1.n164 VDD1.n163 104.615
R634 VDD1.n165 VDD1.n164 104.615
R635 VDD1.n165 VDD1.n92 104.615
R636 VDD1.n172 VDD1.n92 104.615
R637 VDD1.n173 VDD1.n172 104.615
R638 VDD1 VDD1.n177 95.0504
R639 VDD1.t1 VDD1.n28 52.3082
R640 VDD1.t0 VDD1.n116 52.3082
R641 VDD1 VDD1.n88 50.8554
R642 VDD1.n30 VDD1.n29 15.6677
R643 VDD1.n118 VDD1.n117 15.6677
R644 VDD1.n77 VDD1.n6 13.1884
R645 VDD1.n166 VDD1.n95 13.1884
R646 VDD1.n78 VDD1.n4 12.8005
R647 VDD1.n73 VDD1.n8 12.8005
R648 VDD1.n33 VDD1.n32 12.8005
R649 VDD1.n121 VDD1.n120 12.8005
R650 VDD1.n162 VDD1.n161 12.8005
R651 VDD1.n167 VDD1.n93 12.8005
R652 VDD1.n82 VDD1.n81 12.0247
R653 VDD1.n72 VDD1.n9 12.0247
R654 VDD1.n36 VDD1.n27 12.0247
R655 VDD1.n124 VDD1.n115 12.0247
R656 VDD1.n160 VDD1.n97 12.0247
R657 VDD1.n171 VDD1.n170 12.0247
R658 VDD1.n85 VDD1.n2 11.249
R659 VDD1.n69 VDD1.n68 11.249
R660 VDD1.n37 VDD1.n25 11.249
R661 VDD1.n125 VDD1.n113 11.249
R662 VDD1.n157 VDD1.n156 11.249
R663 VDD1.n174 VDD1.n91 11.249
R664 VDD1.n86 VDD1.n0 10.4732
R665 VDD1.n65 VDD1.n11 10.4732
R666 VDD1.n41 VDD1.n40 10.4732
R667 VDD1.n129 VDD1.n128 10.4732
R668 VDD1.n153 VDD1.n99 10.4732
R669 VDD1.n175 VDD1.n89 10.4732
R670 VDD1.n64 VDD1.n13 9.69747
R671 VDD1.n44 VDD1.n23 9.69747
R672 VDD1.n132 VDD1.n111 9.69747
R673 VDD1.n152 VDD1.n101 9.69747
R674 VDD1.n88 VDD1.n87 9.45567
R675 VDD1.n177 VDD1.n176 9.45567
R676 VDD1.n56 VDD1.n55 9.3005
R677 VDD1.n15 VDD1.n14 9.3005
R678 VDD1.n62 VDD1.n61 9.3005
R679 VDD1.n64 VDD1.n63 9.3005
R680 VDD1.n11 VDD1.n10 9.3005
R681 VDD1.n70 VDD1.n69 9.3005
R682 VDD1.n72 VDD1.n71 9.3005
R683 VDD1.n8 VDD1.n5 9.3005
R684 VDD1.n87 VDD1.n86 9.3005
R685 VDD1.n2 VDD1.n1 9.3005
R686 VDD1.n81 VDD1.n80 9.3005
R687 VDD1.n79 VDD1.n78 9.3005
R688 VDD1.n54 VDD1.n53 9.3005
R689 VDD1.n19 VDD1.n18 9.3005
R690 VDD1.n48 VDD1.n47 9.3005
R691 VDD1.n46 VDD1.n45 9.3005
R692 VDD1.n23 VDD1.n22 9.3005
R693 VDD1.n40 VDD1.n39 9.3005
R694 VDD1.n38 VDD1.n37 9.3005
R695 VDD1.n27 VDD1.n26 9.3005
R696 VDD1.n32 VDD1.n31 9.3005
R697 VDD1.n176 VDD1.n175 9.3005
R698 VDD1.n91 VDD1.n90 9.3005
R699 VDD1.n170 VDD1.n169 9.3005
R700 VDD1.n168 VDD1.n167 9.3005
R701 VDD1.n107 VDD1.n106 9.3005
R702 VDD1.n136 VDD1.n135 9.3005
R703 VDD1.n134 VDD1.n133 9.3005
R704 VDD1.n111 VDD1.n110 9.3005
R705 VDD1.n128 VDD1.n127 9.3005
R706 VDD1.n126 VDD1.n125 9.3005
R707 VDD1.n115 VDD1.n114 9.3005
R708 VDD1.n120 VDD1.n119 9.3005
R709 VDD1.n142 VDD1.n141 9.3005
R710 VDD1.n144 VDD1.n143 9.3005
R711 VDD1.n103 VDD1.n102 9.3005
R712 VDD1.n150 VDD1.n149 9.3005
R713 VDD1.n152 VDD1.n151 9.3005
R714 VDD1.n99 VDD1.n98 9.3005
R715 VDD1.n158 VDD1.n157 9.3005
R716 VDD1.n160 VDD1.n159 9.3005
R717 VDD1.n161 VDD1.n94 9.3005
R718 VDD1.n61 VDD1.n60 8.92171
R719 VDD1.n45 VDD1.n21 8.92171
R720 VDD1.n133 VDD1.n109 8.92171
R721 VDD1.n149 VDD1.n148 8.92171
R722 VDD1.n57 VDD1.n15 8.14595
R723 VDD1.n49 VDD1.n48 8.14595
R724 VDD1.n137 VDD1.n136 8.14595
R725 VDD1.n145 VDD1.n103 8.14595
R726 VDD1.n56 VDD1.n17 7.3702
R727 VDD1.n52 VDD1.n19 7.3702
R728 VDD1.n140 VDD1.n107 7.3702
R729 VDD1.n144 VDD1.n105 7.3702
R730 VDD1.n53 VDD1.n17 6.59444
R731 VDD1.n53 VDD1.n52 6.59444
R732 VDD1.n141 VDD1.n140 6.59444
R733 VDD1.n141 VDD1.n105 6.59444
R734 VDD1.n57 VDD1.n56 5.81868
R735 VDD1.n49 VDD1.n19 5.81868
R736 VDD1.n137 VDD1.n107 5.81868
R737 VDD1.n145 VDD1.n144 5.81868
R738 VDD1.n60 VDD1.n15 5.04292
R739 VDD1.n48 VDD1.n21 5.04292
R740 VDD1.n136 VDD1.n109 5.04292
R741 VDD1.n148 VDD1.n103 5.04292
R742 VDD1.n31 VDD1.n30 4.38563
R743 VDD1.n119 VDD1.n118 4.38563
R744 VDD1.n61 VDD1.n13 4.26717
R745 VDD1.n45 VDD1.n44 4.26717
R746 VDD1.n133 VDD1.n132 4.26717
R747 VDD1.n149 VDD1.n101 4.26717
R748 VDD1.n88 VDD1.n0 3.49141
R749 VDD1.n65 VDD1.n64 3.49141
R750 VDD1.n41 VDD1.n23 3.49141
R751 VDD1.n129 VDD1.n111 3.49141
R752 VDD1.n153 VDD1.n152 3.49141
R753 VDD1.n177 VDD1.n89 3.49141
R754 VDD1.n86 VDD1.n85 2.71565
R755 VDD1.n68 VDD1.n11 2.71565
R756 VDD1.n40 VDD1.n25 2.71565
R757 VDD1.n128 VDD1.n113 2.71565
R758 VDD1.n156 VDD1.n99 2.71565
R759 VDD1.n175 VDD1.n174 2.71565
R760 VDD1.n82 VDD1.n2 1.93989
R761 VDD1.n69 VDD1.n9 1.93989
R762 VDD1.n37 VDD1.n36 1.93989
R763 VDD1.n125 VDD1.n124 1.93989
R764 VDD1.n157 VDD1.n97 1.93989
R765 VDD1.n171 VDD1.n91 1.93989
R766 VDD1.n81 VDD1.n4 1.16414
R767 VDD1.n73 VDD1.n72 1.16414
R768 VDD1.n33 VDD1.n27 1.16414
R769 VDD1.n121 VDD1.n115 1.16414
R770 VDD1.n162 VDD1.n160 1.16414
R771 VDD1.n170 VDD1.n93 1.16414
R772 VDD1.n78 VDD1.n77 0.388379
R773 VDD1.n8 VDD1.n6 0.388379
R774 VDD1.n32 VDD1.n29 0.388379
R775 VDD1.n120 VDD1.n117 0.388379
R776 VDD1.n161 VDD1.n95 0.388379
R777 VDD1.n167 VDD1.n166 0.388379
R778 VDD1.n87 VDD1.n1 0.155672
R779 VDD1.n80 VDD1.n1 0.155672
R780 VDD1.n80 VDD1.n79 0.155672
R781 VDD1.n79 VDD1.n5 0.155672
R782 VDD1.n71 VDD1.n5 0.155672
R783 VDD1.n71 VDD1.n70 0.155672
R784 VDD1.n70 VDD1.n10 0.155672
R785 VDD1.n63 VDD1.n10 0.155672
R786 VDD1.n63 VDD1.n62 0.155672
R787 VDD1.n62 VDD1.n14 0.155672
R788 VDD1.n55 VDD1.n14 0.155672
R789 VDD1.n55 VDD1.n54 0.155672
R790 VDD1.n54 VDD1.n18 0.155672
R791 VDD1.n47 VDD1.n18 0.155672
R792 VDD1.n47 VDD1.n46 0.155672
R793 VDD1.n46 VDD1.n22 0.155672
R794 VDD1.n39 VDD1.n22 0.155672
R795 VDD1.n39 VDD1.n38 0.155672
R796 VDD1.n38 VDD1.n26 0.155672
R797 VDD1.n31 VDD1.n26 0.155672
R798 VDD1.n119 VDD1.n114 0.155672
R799 VDD1.n126 VDD1.n114 0.155672
R800 VDD1.n127 VDD1.n126 0.155672
R801 VDD1.n127 VDD1.n110 0.155672
R802 VDD1.n134 VDD1.n110 0.155672
R803 VDD1.n135 VDD1.n134 0.155672
R804 VDD1.n135 VDD1.n106 0.155672
R805 VDD1.n142 VDD1.n106 0.155672
R806 VDD1.n143 VDD1.n142 0.155672
R807 VDD1.n143 VDD1.n102 0.155672
R808 VDD1.n150 VDD1.n102 0.155672
R809 VDD1.n151 VDD1.n150 0.155672
R810 VDD1.n151 VDD1.n98 0.155672
R811 VDD1.n158 VDD1.n98 0.155672
R812 VDD1.n159 VDD1.n158 0.155672
R813 VDD1.n159 VDD1.n94 0.155672
R814 VDD1.n168 VDD1.n94 0.155672
R815 VDD1.n169 VDD1.n168 0.155672
R816 VDD1.n169 VDD1.n90 0.155672
R817 VDD1.n176 VDD1.n90 0.155672
R818 B.n831 B.n830 585
R819 B.n832 B.n831 585
R820 B.n351 B.n114 585
R821 B.n350 B.n349 585
R822 B.n348 B.n347 585
R823 B.n346 B.n345 585
R824 B.n344 B.n343 585
R825 B.n342 B.n341 585
R826 B.n340 B.n339 585
R827 B.n338 B.n337 585
R828 B.n336 B.n335 585
R829 B.n334 B.n333 585
R830 B.n332 B.n331 585
R831 B.n330 B.n329 585
R832 B.n328 B.n327 585
R833 B.n326 B.n325 585
R834 B.n324 B.n323 585
R835 B.n322 B.n321 585
R836 B.n320 B.n319 585
R837 B.n318 B.n317 585
R838 B.n316 B.n315 585
R839 B.n314 B.n313 585
R840 B.n312 B.n311 585
R841 B.n310 B.n309 585
R842 B.n308 B.n307 585
R843 B.n306 B.n305 585
R844 B.n304 B.n303 585
R845 B.n302 B.n301 585
R846 B.n300 B.n299 585
R847 B.n298 B.n297 585
R848 B.n296 B.n295 585
R849 B.n294 B.n293 585
R850 B.n292 B.n291 585
R851 B.n290 B.n289 585
R852 B.n288 B.n287 585
R853 B.n286 B.n285 585
R854 B.n284 B.n283 585
R855 B.n282 B.n281 585
R856 B.n280 B.n279 585
R857 B.n278 B.n277 585
R858 B.n276 B.n275 585
R859 B.n274 B.n273 585
R860 B.n272 B.n271 585
R861 B.n270 B.n269 585
R862 B.n268 B.n267 585
R863 B.n266 B.n265 585
R864 B.n264 B.n263 585
R865 B.n262 B.n261 585
R866 B.n260 B.n259 585
R867 B.n258 B.n257 585
R868 B.n256 B.n255 585
R869 B.n254 B.n253 585
R870 B.n252 B.n251 585
R871 B.n250 B.n249 585
R872 B.n248 B.n247 585
R873 B.n245 B.n244 585
R874 B.n243 B.n242 585
R875 B.n241 B.n240 585
R876 B.n239 B.n238 585
R877 B.n237 B.n236 585
R878 B.n235 B.n234 585
R879 B.n233 B.n232 585
R880 B.n231 B.n230 585
R881 B.n229 B.n228 585
R882 B.n227 B.n226 585
R883 B.n225 B.n224 585
R884 B.n223 B.n222 585
R885 B.n221 B.n220 585
R886 B.n219 B.n218 585
R887 B.n217 B.n216 585
R888 B.n215 B.n214 585
R889 B.n213 B.n212 585
R890 B.n211 B.n210 585
R891 B.n209 B.n208 585
R892 B.n207 B.n206 585
R893 B.n205 B.n204 585
R894 B.n203 B.n202 585
R895 B.n201 B.n200 585
R896 B.n199 B.n198 585
R897 B.n197 B.n196 585
R898 B.n195 B.n194 585
R899 B.n193 B.n192 585
R900 B.n191 B.n190 585
R901 B.n189 B.n188 585
R902 B.n187 B.n186 585
R903 B.n185 B.n184 585
R904 B.n183 B.n182 585
R905 B.n181 B.n180 585
R906 B.n179 B.n178 585
R907 B.n177 B.n176 585
R908 B.n175 B.n174 585
R909 B.n173 B.n172 585
R910 B.n171 B.n170 585
R911 B.n169 B.n168 585
R912 B.n167 B.n166 585
R913 B.n165 B.n164 585
R914 B.n163 B.n162 585
R915 B.n161 B.n160 585
R916 B.n159 B.n158 585
R917 B.n157 B.n156 585
R918 B.n155 B.n154 585
R919 B.n153 B.n152 585
R920 B.n151 B.n150 585
R921 B.n149 B.n148 585
R922 B.n147 B.n146 585
R923 B.n145 B.n144 585
R924 B.n143 B.n142 585
R925 B.n141 B.n140 585
R926 B.n139 B.n138 585
R927 B.n137 B.n136 585
R928 B.n135 B.n134 585
R929 B.n133 B.n132 585
R930 B.n131 B.n130 585
R931 B.n129 B.n128 585
R932 B.n127 B.n126 585
R933 B.n125 B.n124 585
R934 B.n123 B.n122 585
R935 B.n121 B.n120 585
R936 B.n829 B.n55 585
R937 B.n833 B.n55 585
R938 B.n828 B.n54 585
R939 B.n834 B.n54 585
R940 B.n827 B.n826 585
R941 B.n826 B.n50 585
R942 B.n825 B.n49 585
R943 B.n840 B.n49 585
R944 B.n824 B.n48 585
R945 B.n841 B.n48 585
R946 B.n823 B.n47 585
R947 B.n842 B.n47 585
R948 B.n822 B.n821 585
R949 B.n821 B.n43 585
R950 B.n820 B.n42 585
R951 B.n848 B.n42 585
R952 B.n819 B.n41 585
R953 B.n849 B.n41 585
R954 B.n818 B.n40 585
R955 B.n850 B.n40 585
R956 B.n817 B.n816 585
R957 B.n816 B.n36 585
R958 B.n815 B.n35 585
R959 B.n856 B.n35 585
R960 B.n814 B.n34 585
R961 B.n857 B.n34 585
R962 B.n813 B.n33 585
R963 B.n858 B.n33 585
R964 B.n812 B.n811 585
R965 B.n811 B.n29 585
R966 B.n810 B.n28 585
R967 B.n864 B.n28 585
R968 B.n809 B.n27 585
R969 B.n865 B.n27 585
R970 B.n808 B.n26 585
R971 B.n866 B.n26 585
R972 B.n807 B.n806 585
R973 B.n806 B.n22 585
R974 B.n805 B.n21 585
R975 B.n872 B.n21 585
R976 B.n804 B.n20 585
R977 B.n873 B.n20 585
R978 B.n803 B.n19 585
R979 B.n874 B.n19 585
R980 B.n802 B.n801 585
R981 B.n801 B.n18 585
R982 B.n800 B.n14 585
R983 B.n880 B.n14 585
R984 B.n799 B.n13 585
R985 B.n881 B.n13 585
R986 B.n798 B.n12 585
R987 B.n882 B.n12 585
R988 B.n797 B.n796 585
R989 B.n796 B.n8 585
R990 B.n795 B.n7 585
R991 B.n888 B.n7 585
R992 B.n794 B.n6 585
R993 B.n889 B.n6 585
R994 B.n793 B.n5 585
R995 B.n890 B.n5 585
R996 B.n792 B.n791 585
R997 B.n791 B.n4 585
R998 B.n790 B.n352 585
R999 B.n790 B.n789 585
R1000 B.n780 B.n353 585
R1001 B.n354 B.n353 585
R1002 B.n782 B.n781 585
R1003 B.n783 B.n782 585
R1004 B.n779 B.n359 585
R1005 B.n359 B.n358 585
R1006 B.n778 B.n777 585
R1007 B.n777 B.n776 585
R1008 B.n361 B.n360 585
R1009 B.n769 B.n361 585
R1010 B.n768 B.n767 585
R1011 B.n770 B.n768 585
R1012 B.n766 B.n366 585
R1013 B.n366 B.n365 585
R1014 B.n765 B.n764 585
R1015 B.n764 B.n763 585
R1016 B.n368 B.n367 585
R1017 B.n369 B.n368 585
R1018 B.n756 B.n755 585
R1019 B.n757 B.n756 585
R1020 B.n754 B.n374 585
R1021 B.n374 B.n373 585
R1022 B.n753 B.n752 585
R1023 B.n752 B.n751 585
R1024 B.n376 B.n375 585
R1025 B.n377 B.n376 585
R1026 B.n744 B.n743 585
R1027 B.n745 B.n744 585
R1028 B.n742 B.n382 585
R1029 B.n382 B.n381 585
R1030 B.n741 B.n740 585
R1031 B.n740 B.n739 585
R1032 B.n384 B.n383 585
R1033 B.n385 B.n384 585
R1034 B.n732 B.n731 585
R1035 B.n733 B.n732 585
R1036 B.n730 B.n389 585
R1037 B.n393 B.n389 585
R1038 B.n729 B.n728 585
R1039 B.n728 B.n727 585
R1040 B.n391 B.n390 585
R1041 B.n392 B.n391 585
R1042 B.n720 B.n719 585
R1043 B.n721 B.n720 585
R1044 B.n718 B.n398 585
R1045 B.n398 B.n397 585
R1046 B.n717 B.n716 585
R1047 B.n716 B.n715 585
R1048 B.n400 B.n399 585
R1049 B.n401 B.n400 585
R1050 B.n708 B.n707 585
R1051 B.n709 B.n708 585
R1052 B.n706 B.n406 585
R1053 B.n406 B.n405 585
R1054 B.n700 B.n699 585
R1055 B.n698 B.n466 585
R1056 B.n697 B.n465 585
R1057 B.n702 B.n465 585
R1058 B.n696 B.n695 585
R1059 B.n694 B.n693 585
R1060 B.n692 B.n691 585
R1061 B.n690 B.n689 585
R1062 B.n688 B.n687 585
R1063 B.n686 B.n685 585
R1064 B.n684 B.n683 585
R1065 B.n682 B.n681 585
R1066 B.n680 B.n679 585
R1067 B.n678 B.n677 585
R1068 B.n676 B.n675 585
R1069 B.n674 B.n673 585
R1070 B.n672 B.n671 585
R1071 B.n670 B.n669 585
R1072 B.n668 B.n667 585
R1073 B.n666 B.n665 585
R1074 B.n664 B.n663 585
R1075 B.n662 B.n661 585
R1076 B.n660 B.n659 585
R1077 B.n658 B.n657 585
R1078 B.n656 B.n655 585
R1079 B.n654 B.n653 585
R1080 B.n652 B.n651 585
R1081 B.n650 B.n649 585
R1082 B.n648 B.n647 585
R1083 B.n646 B.n645 585
R1084 B.n644 B.n643 585
R1085 B.n642 B.n641 585
R1086 B.n640 B.n639 585
R1087 B.n638 B.n637 585
R1088 B.n636 B.n635 585
R1089 B.n634 B.n633 585
R1090 B.n632 B.n631 585
R1091 B.n630 B.n629 585
R1092 B.n628 B.n627 585
R1093 B.n626 B.n625 585
R1094 B.n624 B.n623 585
R1095 B.n622 B.n621 585
R1096 B.n620 B.n619 585
R1097 B.n618 B.n617 585
R1098 B.n616 B.n615 585
R1099 B.n614 B.n613 585
R1100 B.n612 B.n611 585
R1101 B.n610 B.n609 585
R1102 B.n608 B.n607 585
R1103 B.n606 B.n605 585
R1104 B.n604 B.n603 585
R1105 B.n602 B.n601 585
R1106 B.n600 B.n599 585
R1107 B.n598 B.n597 585
R1108 B.n596 B.n595 585
R1109 B.n593 B.n592 585
R1110 B.n591 B.n590 585
R1111 B.n589 B.n588 585
R1112 B.n587 B.n586 585
R1113 B.n585 B.n584 585
R1114 B.n583 B.n582 585
R1115 B.n581 B.n580 585
R1116 B.n579 B.n578 585
R1117 B.n577 B.n576 585
R1118 B.n575 B.n574 585
R1119 B.n573 B.n572 585
R1120 B.n571 B.n570 585
R1121 B.n569 B.n568 585
R1122 B.n567 B.n566 585
R1123 B.n565 B.n564 585
R1124 B.n563 B.n562 585
R1125 B.n561 B.n560 585
R1126 B.n559 B.n558 585
R1127 B.n557 B.n556 585
R1128 B.n555 B.n554 585
R1129 B.n553 B.n552 585
R1130 B.n551 B.n550 585
R1131 B.n549 B.n548 585
R1132 B.n547 B.n546 585
R1133 B.n545 B.n544 585
R1134 B.n543 B.n542 585
R1135 B.n541 B.n540 585
R1136 B.n539 B.n538 585
R1137 B.n537 B.n536 585
R1138 B.n535 B.n534 585
R1139 B.n533 B.n532 585
R1140 B.n531 B.n530 585
R1141 B.n529 B.n528 585
R1142 B.n527 B.n526 585
R1143 B.n525 B.n524 585
R1144 B.n523 B.n522 585
R1145 B.n521 B.n520 585
R1146 B.n519 B.n518 585
R1147 B.n517 B.n516 585
R1148 B.n515 B.n514 585
R1149 B.n513 B.n512 585
R1150 B.n511 B.n510 585
R1151 B.n509 B.n508 585
R1152 B.n507 B.n506 585
R1153 B.n505 B.n504 585
R1154 B.n503 B.n502 585
R1155 B.n501 B.n500 585
R1156 B.n499 B.n498 585
R1157 B.n497 B.n496 585
R1158 B.n495 B.n494 585
R1159 B.n493 B.n492 585
R1160 B.n491 B.n490 585
R1161 B.n489 B.n488 585
R1162 B.n487 B.n486 585
R1163 B.n485 B.n484 585
R1164 B.n483 B.n482 585
R1165 B.n481 B.n480 585
R1166 B.n479 B.n478 585
R1167 B.n477 B.n476 585
R1168 B.n475 B.n474 585
R1169 B.n473 B.n472 585
R1170 B.n408 B.n407 585
R1171 B.n705 B.n704 585
R1172 B.n404 B.n403 585
R1173 B.n405 B.n404 585
R1174 B.n711 B.n710 585
R1175 B.n710 B.n709 585
R1176 B.n712 B.n402 585
R1177 B.n402 B.n401 585
R1178 B.n714 B.n713 585
R1179 B.n715 B.n714 585
R1180 B.n396 B.n395 585
R1181 B.n397 B.n396 585
R1182 B.n723 B.n722 585
R1183 B.n722 B.n721 585
R1184 B.n724 B.n394 585
R1185 B.n394 B.n392 585
R1186 B.n726 B.n725 585
R1187 B.n727 B.n726 585
R1188 B.n388 B.n387 585
R1189 B.n393 B.n388 585
R1190 B.n735 B.n734 585
R1191 B.n734 B.n733 585
R1192 B.n736 B.n386 585
R1193 B.n386 B.n385 585
R1194 B.n738 B.n737 585
R1195 B.n739 B.n738 585
R1196 B.n380 B.n379 585
R1197 B.n381 B.n380 585
R1198 B.n747 B.n746 585
R1199 B.n746 B.n745 585
R1200 B.n748 B.n378 585
R1201 B.n378 B.n377 585
R1202 B.n750 B.n749 585
R1203 B.n751 B.n750 585
R1204 B.n372 B.n371 585
R1205 B.n373 B.n372 585
R1206 B.n759 B.n758 585
R1207 B.n758 B.n757 585
R1208 B.n760 B.n370 585
R1209 B.n370 B.n369 585
R1210 B.n762 B.n761 585
R1211 B.n763 B.n762 585
R1212 B.n364 B.n363 585
R1213 B.n365 B.n364 585
R1214 B.n772 B.n771 585
R1215 B.n771 B.n770 585
R1216 B.n773 B.n362 585
R1217 B.n769 B.n362 585
R1218 B.n775 B.n774 585
R1219 B.n776 B.n775 585
R1220 B.n357 B.n356 585
R1221 B.n358 B.n357 585
R1222 B.n785 B.n784 585
R1223 B.n784 B.n783 585
R1224 B.n786 B.n355 585
R1225 B.n355 B.n354 585
R1226 B.n788 B.n787 585
R1227 B.n789 B.n788 585
R1228 B.n2 B.n0 585
R1229 B.n4 B.n2 585
R1230 B.n3 B.n1 585
R1231 B.n889 B.n3 585
R1232 B.n887 B.n886 585
R1233 B.n888 B.n887 585
R1234 B.n885 B.n9 585
R1235 B.n9 B.n8 585
R1236 B.n884 B.n883 585
R1237 B.n883 B.n882 585
R1238 B.n11 B.n10 585
R1239 B.n881 B.n11 585
R1240 B.n879 B.n878 585
R1241 B.n880 B.n879 585
R1242 B.n877 B.n15 585
R1243 B.n18 B.n15 585
R1244 B.n876 B.n875 585
R1245 B.n875 B.n874 585
R1246 B.n17 B.n16 585
R1247 B.n873 B.n17 585
R1248 B.n871 B.n870 585
R1249 B.n872 B.n871 585
R1250 B.n869 B.n23 585
R1251 B.n23 B.n22 585
R1252 B.n868 B.n867 585
R1253 B.n867 B.n866 585
R1254 B.n25 B.n24 585
R1255 B.n865 B.n25 585
R1256 B.n863 B.n862 585
R1257 B.n864 B.n863 585
R1258 B.n861 B.n30 585
R1259 B.n30 B.n29 585
R1260 B.n860 B.n859 585
R1261 B.n859 B.n858 585
R1262 B.n32 B.n31 585
R1263 B.n857 B.n32 585
R1264 B.n855 B.n854 585
R1265 B.n856 B.n855 585
R1266 B.n853 B.n37 585
R1267 B.n37 B.n36 585
R1268 B.n852 B.n851 585
R1269 B.n851 B.n850 585
R1270 B.n39 B.n38 585
R1271 B.n849 B.n39 585
R1272 B.n847 B.n846 585
R1273 B.n848 B.n847 585
R1274 B.n845 B.n44 585
R1275 B.n44 B.n43 585
R1276 B.n844 B.n843 585
R1277 B.n843 B.n842 585
R1278 B.n46 B.n45 585
R1279 B.n841 B.n46 585
R1280 B.n839 B.n838 585
R1281 B.n840 B.n839 585
R1282 B.n837 B.n51 585
R1283 B.n51 B.n50 585
R1284 B.n836 B.n835 585
R1285 B.n835 B.n834 585
R1286 B.n53 B.n52 585
R1287 B.n833 B.n53 585
R1288 B.n892 B.n891 585
R1289 B.n891 B.n890 585
R1290 B.n700 B.n404 530.939
R1291 B.n120 B.n53 530.939
R1292 B.n704 B.n406 530.939
R1293 B.n831 B.n55 530.939
R1294 B.n469 B.t12 422.683
R1295 B.n115 B.t4 422.683
R1296 B.n467 B.t9 422.683
R1297 B.n117 B.t14 422.683
R1298 B.n470 B.t11 353.447
R1299 B.n116 B.t5 353.447
R1300 B.n468 B.t8 353.447
R1301 B.n118 B.t15 353.447
R1302 B.n469 B.t10 328.899
R1303 B.n467 B.t6 328.899
R1304 B.n117 B.t13 328.899
R1305 B.n115 B.t2 328.899
R1306 B.n832 B.n113 256.663
R1307 B.n832 B.n112 256.663
R1308 B.n832 B.n111 256.663
R1309 B.n832 B.n110 256.663
R1310 B.n832 B.n109 256.663
R1311 B.n832 B.n108 256.663
R1312 B.n832 B.n107 256.663
R1313 B.n832 B.n106 256.663
R1314 B.n832 B.n105 256.663
R1315 B.n832 B.n104 256.663
R1316 B.n832 B.n103 256.663
R1317 B.n832 B.n102 256.663
R1318 B.n832 B.n101 256.663
R1319 B.n832 B.n100 256.663
R1320 B.n832 B.n99 256.663
R1321 B.n832 B.n98 256.663
R1322 B.n832 B.n97 256.663
R1323 B.n832 B.n96 256.663
R1324 B.n832 B.n95 256.663
R1325 B.n832 B.n94 256.663
R1326 B.n832 B.n93 256.663
R1327 B.n832 B.n92 256.663
R1328 B.n832 B.n91 256.663
R1329 B.n832 B.n90 256.663
R1330 B.n832 B.n89 256.663
R1331 B.n832 B.n88 256.663
R1332 B.n832 B.n87 256.663
R1333 B.n832 B.n86 256.663
R1334 B.n832 B.n85 256.663
R1335 B.n832 B.n84 256.663
R1336 B.n832 B.n83 256.663
R1337 B.n832 B.n82 256.663
R1338 B.n832 B.n81 256.663
R1339 B.n832 B.n80 256.663
R1340 B.n832 B.n79 256.663
R1341 B.n832 B.n78 256.663
R1342 B.n832 B.n77 256.663
R1343 B.n832 B.n76 256.663
R1344 B.n832 B.n75 256.663
R1345 B.n832 B.n74 256.663
R1346 B.n832 B.n73 256.663
R1347 B.n832 B.n72 256.663
R1348 B.n832 B.n71 256.663
R1349 B.n832 B.n70 256.663
R1350 B.n832 B.n69 256.663
R1351 B.n832 B.n68 256.663
R1352 B.n832 B.n67 256.663
R1353 B.n832 B.n66 256.663
R1354 B.n832 B.n65 256.663
R1355 B.n832 B.n64 256.663
R1356 B.n832 B.n63 256.663
R1357 B.n832 B.n62 256.663
R1358 B.n832 B.n61 256.663
R1359 B.n832 B.n60 256.663
R1360 B.n832 B.n59 256.663
R1361 B.n832 B.n58 256.663
R1362 B.n832 B.n57 256.663
R1363 B.n832 B.n56 256.663
R1364 B.n702 B.n701 256.663
R1365 B.n702 B.n409 256.663
R1366 B.n702 B.n410 256.663
R1367 B.n702 B.n411 256.663
R1368 B.n702 B.n412 256.663
R1369 B.n702 B.n413 256.663
R1370 B.n702 B.n414 256.663
R1371 B.n702 B.n415 256.663
R1372 B.n702 B.n416 256.663
R1373 B.n702 B.n417 256.663
R1374 B.n702 B.n418 256.663
R1375 B.n702 B.n419 256.663
R1376 B.n702 B.n420 256.663
R1377 B.n702 B.n421 256.663
R1378 B.n702 B.n422 256.663
R1379 B.n702 B.n423 256.663
R1380 B.n702 B.n424 256.663
R1381 B.n702 B.n425 256.663
R1382 B.n702 B.n426 256.663
R1383 B.n702 B.n427 256.663
R1384 B.n702 B.n428 256.663
R1385 B.n702 B.n429 256.663
R1386 B.n702 B.n430 256.663
R1387 B.n702 B.n431 256.663
R1388 B.n702 B.n432 256.663
R1389 B.n702 B.n433 256.663
R1390 B.n702 B.n434 256.663
R1391 B.n702 B.n435 256.663
R1392 B.n702 B.n436 256.663
R1393 B.n702 B.n437 256.663
R1394 B.n702 B.n438 256.663
R1395 B.n702 B.n439 256.663
R1396 B.n702 B.n440 256.663
R1397 B.n702 B.n441 256.663
R1398 B.n702 B.n442 256.663
R1399 B.n702 B.n443 256.663
R1400 B.n702 B.n444 256.663
R1401 B.n702 B.n445 256.663
R1402 B.n702 B.n446 256.663
R1403 B.n702 B.n447 256.663
R1404 B.n702 B.n448 256.663
R1405 B.n702 B.n449 256.663
R1406 B.n702 B.n450 256.663
R1407 B.n702 B.n451 256.663
R1408 B.n702 B.n452 256.663
R1409 B.n702 B.n453 256.663
R1410 B.n702 B.n454 256.663
R1411 B.n702 B.n455 256.663
R1412 B.n702 B.n456 256.663
R1413 B.n702 B.n457 256.663
R1414 B.n702 B.n458 256.663
R1415 B.n702 B.n459 256.663
R1416 B.n702 B.n460 256.663
R1417 B.n702 B.n461 256.663
R1418 B.n702 B.n462 256.663
R1419 B.n702 B.n463 256.663
R1420 B.n702 B.n464 256.663
R1421 B.n703 B.n702 256.663
R1422 B.n710 B.n404 163.367
R1423 B.n710 B.n402 163.367
R1424 B.n714 B.n402 163.367
R1425 B.n714 B.n396 163.367
R1426 B.n722 B.n396 163.367
R1427 B.n722 B.n394 163.367
R1428 B.n726 B.n394 163.367
R1429 B.n726 B.n388 163.367
R1430 B.n734 B.n388 163.367
R1431 B.n734 B.n386 163.367
R1432 B.n738 B.n386 163.367
R1433 B.n738 B.n380 163.367
R1434 B.n746 B.n380 163.367
R1435 B.n746 B.n378 163.367
R1436 B.n750 B.n378 163.367
R1437 B.n750 B.n372 163.367
R1438 B.n758 B.n372 163.367
R1439 B.n758 B.n370 163.367
R1440 B.n762 B.n370 163.367
R1441 B.n762 B.n364 163.367
R1442 B.n771 B.n364 163.367
R1443 B.n771 B.n362 163.367
R1444 B.n775 B.n362 163.367
R1445 B.n775 B.n357 163.367
R1446 B.n784 B.n357 163.367
R1447 B.n784 B.n355 163.367
R1448 B.n788 B.n355 163.367
R1449 B.n788 B.n2 163.367
R1450 B.n891 B.n2 163.367
R1451 B.n891 B.n3 163.367
R1452 B.n887 B.n3 163.367
R1453 B.n887 B.n9 163.367
R1454 B.n883 B.n9 163.367
R1455 B.n883 B.n11 163.367
R1456 B.n879 B.n11 163.367
R1457 B.n879 B.n15 163.367
R1458 B.n875 B.n15 163.367
R1459 B.n875 B.n17 163.367
R1460 B.n871 B.n17 163.367
R1461 B.n871 B.n23 163.367
R1462 B.n867 B.n23 163.367
R1463 B.n867 B.n25 163.367
R1464 B.n863 B.n25 163.367
R1465 B.n863 B.n30 163.367
R1466 B.n859 B.n30 163.367
R1467 B.n859 B.n32 163.367
R1468 B.n855 B.n32 163.367
R1469 B.n855 B.n37 163.367
R1470 B.n851 B.n37 163.367
R1471 B.n851 B.n39 163.367
R1472 B.n847 B.n39 163.367
R1473 B.n847 B.n44 163.367
R1474 B.n843 B.n44 163.367
R1475 B.n843 B.n46 163.367
R1476 B.n839 B.n46 163.367
R1477 B.n839 B.n51 163.367
R1478 B.n835 B.n51 163.367
R1479 B.n835 B.n53 163.367
R1480 B.n466 B.n465 163.367
R1481 B.n695 B.n465 163.367
R1482 B.n693 B.n692 163.367
R1483 B.n689 B.n688 163.367
R1484 B.n685 B.n684 163.367
R1485 B.n681 B.n680 163.367
R1486 B.n677 B.n676 163.367
R1487 B.n673 B.n672 163.367
R1488 B.n669 B.n668 163.367
R1489 B.n665 B.n664 163.367
R1490 B.n661 B.n660 163.367
R1491 B.n657 B.n656 163.367
R1492 B.n653 B.n652 163.367
R1493 B.n649 B.n648 163.367
R1494 B.n645 B.n644 163.367
R1495 B.n641 B.n640 163.367
R1496 B.n637 B.n636 163.367
R1497 B.n633 B.n632 163.367
R1498 B.n629 B.n628 163.367
R1499 B.n625 B.n624 163.367
R1500 B.n621 B.n620 163.367
R1501 B.n617 B.n616 163.367
R1502 B.n613 B.n612 163.367
R1503 B.n609 B.n608 163.367
R1504 B.n605 B.n604 163.367
R1505 B.n601 B.n600 163.367
R1506 B.n597 B.n596 163.367
R1507 B.n592 B.n591 163.367
R1508 B.n588 B.n587 163.367
R1509 B.n584 B.n583 163.367
R1510 B.n580 B.n579 163.367
R1511 B.n576 B.n575 163.367
R1512 B.n572 B.n571 163.367
R1513 B.n568 B.n567 163.367
R1514 B.n564 B.n563 163.367
R1515 B.n560 B.n559 163.367
R1516 B.n556 B.n555 163.367
R1517 B.n552 B.n551 163.367
R1518 B.n548 B.n547 163.367
R1519 B.n544 B.n543 163.367
R1520 B.n540 B.n539 163.367
R1521 B.n536 B.n535 163.367
R1522 B.n532 B.n531 163.367
R1523 B.n528 B.n527 163.367
R1524 B.n524 B.n523 163.367
R1525 B.n520 B.n519 163.367
R1526 B.n516 B.n515 163.367
R1527 B.n512 B.n511 163.367
R1528 B.n508 B.n507 163.367
R1529 B.n504 B.n503 163.367
R1530 B.n500 B.n499 163.367
R1531 B.n496 B.n495 163.367
R1532 B.n492 B.n491 163.367
R1533 B.n488 B.n487 163.367
R1534 B.n484 B.n483 163.367
R1535 B.n480 B.n479 163.367
R1536 B.n476 B.n475 163.367
R1537 B.n472 B.n408 163.367
R1538 B.n708 B.n406 163.367
R1539 B.n708 B.n400 163.367
R1540 B.n716 B.n400 163.367
R1541 B.n716 B.n398 163.367
R1542 B.n720 B.n398 163.367
R1543 B.n720 B.n391 163.367
R1544 B.n728 B.n391 163.367
R1545 B.n728 B.n389 163.367
R1546 B.n732 B.n389 163.367
R1547 B.n732 B.n384 163.367
R1548 B.n740 B.n384 163.367
R1549 B.n740 B.n382 163.367
R1550 B.n744 B.n382 163.367
R1551 B.n744 B.n376 163.367
R1552 B.n752 B.n376 163.367
R1553 B.n752 B.n374 163.367
R1554 B.n756 B.n374 163.367
R1555 B.n756 B.n368 163.367
R1556 B.n764 B.n368 163.367
R1557 B.n764 B.n366 163.367
R1558 B.n768 B.n366 163.367
R1559 B.n768 B.n361 163.367
R1560 B.n777 B.n361 163.367
R1561 B.n777 B.n359 163.367
R1562 B.n782 B.n359 163.367
R1563 B.n782 B.n353 163.367
R1564 B.n790 B.n353 163.367
R1565 B.n791 B.n790 163.367
R1566 B.n791 B.n5 163.367
R1567 B.n6 B.n5 163.367
R1568 B.n7 B.n6 163.367
R1569 B.n796 B.n7 163.367
R1570 B.n796 B.n12 163.367
R1571 B.n13 B.n12 163.367
R1572 B.n14 B.n13 163.367
R1573 B.n801 B.n14 163.367
R1574 B.n801 B.n19 163.367
R1575 B.n20 B.n19 163.367
R1576 B.n21 B.n20 163.367
R1577 B.n806 B.n21 163.367
R1578 B.n806 B.n26 163.367
R1579 B.n27 B.n26 163.367
R1580 B.n28 B.n27 163.367
R1581 B.n811 B.n28 163.367
R1582 B.n811 B.n33 163.367
R1583 B.n34 B.n33 163.367
R1584 B.n35 B.n34 163.367
R1585 B.n816 B.n35 163.367
R1586 B.n816 B.n40 163.367
R1587 B.n41 B.n40 163.367
R1588 B.n42 B.n41 163.367
R1589 B.n821 B.n42 163.367
R1590 B.n821 B.n47 163.367
R1591 B.n48 B.n47 163.367
R1592 B.n49 B.n48 163.367
R1593 B.n826 B.n49 163.367
R1594 B.n826 B.n54 163.367
R1595 B.n55 B.n54 163.367
R1596 B.n124 B.n123 163.367
R1597 B.n128 B.n127 163.367
R1598 B.n132 B.n131 163.367
R1599 B.n136 B.n135 163.367
R1600 B.n140 B.n139 163.367
R1601 B.n144 B.n143 163.367
R1602 B.n148 B.n147 163.367
R1603 B.n152 B.n151 163.367
R1604 B.n156 B.n155 163.367
R1605 B.n160 B.n159 163.367
R1606 B.n164 B.n163 163.367
R1607 B.n168 B.n167 163.367
R1608 B.n172 B.n171 163.367
R1609 B.n176 B.n175 163.367
R1610 B.n180 B.n179 163.367
R1611 B.n184 B.n183 163.367
R1612 B.n188 B.n187 163.367
R1613 B.n192 B.n191 163.367
R1614 B.n196 B.n195 163.367
R1615 B.n200 B.n199 163.367
R1616 B.n204 B.n203 163.367
R1617 B.n208 B.n207 163.367
R1618 B.n212 B.n211 163.367
R1619 B.n216 B.n215 163.367
R1620 B.n220 B.n219 163.367
R1621 B.n224 B.n223 163.367
R1622 B.n228 B.n227 163.367
R1623 B.n232 B.n231 163.367
R1624 B.n236 B.n235 163.367
R1625 B.n240 B.n239 163.367
R1626 B.n244 B.n243 163.367
R1627 B.n249 B.n248 163.367
R1628 B.n253 B.n252 163.367
R1629 B.n257 B.n256 163.367
R1630 B.n261 B.n260 163.367
R1631 B.n265 B.n264 163.367
R1632 B.n269 B.n268 163.367
R1633 B.n273 B.n272 163.367
R1634 B.n277 B.n276 163.367
R1635 B.n281 B.n280 163.367
R1636 B.n285 B.n284 163.367
R1637 B.n289 B.n288 163.367
R1638 B.n293 B.n292 163.367
R1639 B.n297 B.n296 163.367
R1640 B.n301 B.n300 163.367
R1641 B.n305 B.n304 163.367
R1642 B.n309 B.n308 163.367
R1643 B.n313 B.n312 163.367
R1644 B.n317 B.n316 163.367
R1645 B.n321 B.n320 163.367
R1646 B.n325 B.n324 163.367
R1647 B.n329 B.n328 163.367
R1648 B.n333 B.n332 163.367
R1649 B.n337 B.n336 163.367
R1650 B.n341 B.n340 163.367
R1651 B.n345 B.n344 163.367
R1652 B.n349 B.n348 163.367
R1653 B.n831 B.n114 163.367
R1654 B.n701 B.n700 71.676
R1655 B.n695 B.n409 71.676
R1656 B.n692 B.n410 71.676
R1657 B.n688 B.n411 71.676
R1658 B.n684 B.n412 71.676
R1659 B.n680 B.n413 71.676
R1660 B.n676 B.n414 71.676
R1661 B.n672 B.n415 71.676
R1662 B.n668 B.n416 71.676
R1663 B.n664 B.n417 71.676
R1664 B.n660 B.n418 71.676
R1665 B.n656 B.n419 71.676
R1666 B.n652 B.n420 71.676
R1667 B.n648 B.n421 71.676
R1668 B.n644 B.n422 71.676
R1669 B.n640 B.n423 71.676
R1670 B.n636 B.n424 71.676
R1671 B.n632 B.n425 71.676
R1672 B.n628 B.n426 71.676
R1673 B.n624 B.n427 71.676
R1674 B.n620 B.n428 71.676
R1675 B.n616 B.n429 71.676
R1676 B.n612 B.n430 71.676
R1677 B.n608 B.n431 71.676
R1678 B.n604 B.n432 71.676
R1679 B.n600 B.n433 71.676
R1680 B.n596 B.n434 71.676
R1681 B.n591 B.n435 71.676
R1682 B.n587 B.n436 71.676
R1683 B.n583 B.n437 71.676
R1684 B.n579 B.n438 71.676
R1685 B.n575 B.n439 71.676
R1686 B.n571 B.n440 71.676
R1687 B.n567 B.n441 71.676
R1688 B.n563 B.n442 71.676
R1689 B.n559 B.n443 71.676
R1690 B.n555 B.n444 71.676
R1691 B.n551 B.n445 71.676
R1692 B.n547 B.n446 71.676
R1693 B.n543 B.n447 71.676
R1694 B.n539 B.n448 71.676
R1695 B.n535 B.n449 71.676
R1696 B.n531 B.n450 71.676
R1697 B.n527 B.n451 71.676
R1698 B.n523 B.n452 71.676
R1699 B.n519 B.n453 71.676
R1700 B.n515 B.n454 71.676
R1701 B.n511 B.n455 71.676
R1702 B.n507 B.n456 71.676
R1703 B.n503 B.n457 71.676
R1704 B.n499 B.n458 71.676
R1705 B.n495 B.n459 71.676
R1706 B.n491 B.n460 71.676
R1707 B.n487 B.n461 71.676
R1708 B.n483 B.n462 71.676
R1709 B.n479 B.n463 71.676
R1710 B.n475 B.n464 71.676
R1711 B.n703 B.n408 71.676
R1712 B.n120 B.n56 71.676
R1713 B.n124 B.n57 71.676
R1714 B.n128 B.n58 71.676
R1715 B.n132 B.n59 71.676
R1716 B.n136 B.n60 71.676
R1717 B.n140 B.n61 71.676
R1718 B.n144 B.n62 71.676
R1719 B.n148 B.n63 71.676
R1720 B.n152 B.n64 71.676
R1721 B.n156 B.n65 71.676
R1722 B.n160 B.n66 71.676
R1723 B.n164 B.n67 71.676
R1724 B.n168 B.n68 71.676
R1725 B.n172 B.n69 71.676
R1726 B.n176 B.n70 71.676
R1727 B.n180 B.n71 71.676
R1728 B.n184 B.n72 71.676
R1729 B.n188 B.n73 71.676
R1730 B.n192 B.n74 71.676
R1731 B.n196 B.n75 71.676
R1732 B.n200 B.n76 71.676
R1733 B.n204 B.n77 71.676
R1734 B.n208 B.n78 71.676
R1735 B.n212 B.n79 71.676
R1736 B.n216 B.n80 71.676
R1737 B.n220 B.n81 71.676
R1738 B.n224 B.n82 71.676
R1739 B.n228 B.n83 71.676
R1740 B.n232 B.n84 71.676
R1741 B.n236 B.n85 71.676
R1742 B.n240 B.n86 71.676
R1743 B.n244 B.n87 71.676
R1744 B.n249 B.n88 71.676
R1745 B.n253 B.n89 71.676
R1746 B.n257 B.n90 71.676
R1747 B.n261 B.n91 71.676
R1748 B.n265 B.n92 71.676
R1749 B.n269 B.n93 71.676
R1750 B.n273 B.n94 71.676
R1751 B.n277 B.n95 71.676
R1752 B.n281 B.n96 71.676
R1753 B.n285 B.n97 71.676
R1754 B.n289 B.n98 71.676
R1755 B.n293 B.n99 71.676
R1756 B.n297 B.n100 71.676
R1757 B.n301 B.n101 71.676
R1758 B.n305 B.n102 71.676
R1759 B.n309 B.n103 71.676
R1760 B.n313 B.n104 71.676
R1761 B.n317 B.n105 71.676
R1762 B.n321 B.n106 71.676
R1763 B.n325 B.n107 71.676
R1764 B.n329 B.n108 71.676
R1765 B.n333 B.n109 71.676
R1766 B.n337 B.n110 71.676
R1767 B.n341 B.n111 71.676
R1768 B.n345 B.n112 71.676
R1769 B.n349 B.n113 71.676
R1770 B.n114 B.n113 71.676
R1771 B.n348 B.n112 71.676
R1772 B.n344 B.n111 71.676
R1773 B.n340 B.n110 71.676
R1774 B.n336 B.n109 71.676
R1775 B.n332 B.n108 71.676
R1776 B.n328 B.n107 71.676
R1777 B.n324 B.n106 71.676
R1778 B.n320 B.n105 71.676
R1779 B.n316 B.n104 71.676
R1780 B.n312 B.n103 71.676
R1781 B.n308 B.n102 71.676
R1782 B.n304 B.n101 71.676
R1783 B.n300 B.n100 71.676
R1784 B.n296 B.n99 71.676
R1785 B.n292 B.n98 71.676
R1786 B.n288 B.n97 71.676
R1787 B.n284 B.n96 71.676
R1788 B.n280 B.n95 71.676
R1789 B.n276 B.n94 71.676
R1790 B.n272 B.n93 71.676
R1791 B.n268 B.n92 71.676
R1792 B.n264 B.n91 71.676
R1793 B.n260 B.n90 71.676
R1794 B.n256 B.n89 71.676
R1795 B.n252 B.n88 71.676
R1796 B.n248 B.n87 71.676
R1797 B.n243 B.n86 71.676
R1798 B.n239 B.n85 71.676
R1799 B.n235 B.n84 71.676
R1800 B.n231 B.n83 71.676
R1801 B.n227 B.n82 71.676
R1802 B.n223 B.n81 71.676
R1803 B.n219 B.n80 71.676
R1804 B.n215 B.n79 71.676
R1805 B.n211 B.n78 71.676
R1806 B.n207 B.n77 71.676
R1807 B.n203 B.n76 71.676
R1808 B.n199 B.n75 71.676
R1809 B.n195 B.n74 71.676
R1810 B.n191 B.n73 71.676
R1811 B.n187 B.n72 71.676
R1812 B.n183 B.n71 71.676
R1813 B.n179 B.n70 71.676
R1814 B.n175 B.n69 71.676
R1815 B.n171 B.n68 71.676
R1816 B.n167 B.n67 71.676
R1817 B.n163 B.n66 71.676
R1818 B.n159 B.n65 71.676
R1819 B.n155 B.n64 71.676
R1820 B.n151 B.n63 71.676
R1821 B.n147 B.n62 71.676
R1822 B.n143 B.n61 71.676
R1823 B.n139 B.n60 71.676
R1824 B.n135 B.n59 71.676
R1825 B.n131 B.n58 71.676
R1826 B.n127 B.n57 71.676
R1827 B.n123 B.n56 71.676
R1828 B.n701 B.n466 71.676
R1829 B.n693 B.n409 71.676
R1830 B.n689 B.n410 71.676
R1831 B.n685 B.n411 71.676
R1832 B.n681 B.n412 71.676
R1833 B.n677 B.n413 71.676
R1834 B.n673 B.n414 71.676
R1835 B.n669 B.n415 71.676
R1836 B.n665 B.n416 71.676
R1837 B.n661 B.n417 71.676
R1838 B.n657 B.n418 71.676
R1839 B.n653 B.n419 71.676
R1840 B.n649 B.n420 71.676
R1841 B.n645 B.n421 71.676
R1842 B.n641 B.n422 71.676
R1843 B.n637 B.n423 71.676
R1844 B.n633 B.n424 71.676
R1845 B.n629 B.n425 71.676
R1846 B.n625 B.n426 71.676
R1847 B.n621 B.n427 71.676
R1848 B.n617 B.n428 71.676
R1849 B.n613 B.n429 71.676
R1850 B.n609 B.n430 71.676
R1851 B.n605 B.n431 71.676
R1852 B.n601 B.n432 71.676
R1853 B.n597 B.n433 71.676
R1854 B.n592 B.n434 71.676
R1855 B.n588 B.n435 71.676
R1856 B.n584 B.n436 71.676
R1857 B.n580 B.n437 71.676
R1858 B.n576 B.n438 71.676
R1859 B.n572 B.n439 71.676
R1860 B.n568 B.n440 71.676
R1861 B.n564 B.n441 71.676
R1862 B.n560 B.n442 71.676
R1863 B.n556 B.n443 71.676
R1864 B.n552 B.n444 71.676
R1865 B.n548 B.n445 71.676
R1866 B.n544 B.n446 71.676
R1867 B.n540 B.n447 71.676
R1868 B.n536 B.n448 71.676
R1869 B.n532 B.n449 71.676
R1870 B.n528 B.n450 71.676
R1871 B.n524 B.n451 71.676
R1872 B.n520 B.n452 71.676
R1873 B.n516 B.n453 71.676
R1874 B.n512 B.n454 71.676
R1875 B.n508 B.n455 71.676
R1876 B.n504 B.n456 71.676
R1877 B.n500 B.n457 71.676
R1878 B.n496 B.n458 71.676
R1879 B.n492 B.n459 71.676
R1880 B.n488 B.n460 71.676
R1881 B.n484 B.n461 71.676
R1882 B.n480 B.n462 71.676
R1883 B.n476 B.n463 71.676
R1884 B.n472 B.n464 71.676
R1885 B.n704 B.n703 71.676
R1886 B.n470 B.n469 69.2369
R1887 B.n468 B.n467 69.2369
R1888 B.n118 B.n117 69.2369
R1889 B.n116 B.n115 69.2369
R1890 B.n702 B.n405 67.2898
R1891 B.n833 B.n832 67.2898
R1892 B.n471 B.n470 59.5399
R1893 B.n594 B.n468 59.5399
R1894 B.n119 B.n118 59.5399
R1895 B.n246 B.n116 59.5399
R1896 B.n709 B.n405 34.9293
R1897 B.n709 B.n401 34.9293
R1898 B.n715 B.n401 34.9293
R1899 B.n715 B.n397 34.9293
R1900 B.n721 B.n397 34.9293
R1901 B.n721 B.n392 34.9293
R1902 B.n727 B.n392 34.9293
R1903 B.n727 B.n393 34.9293
R1904 B.n733 B.n385 34.9293
R1905 B.n739 B.n385 34.9293
R1906 B.n739 B.n381 34.9293
R1907 B.n745 B.n381 34.9293
R1908 B.n745 B.n377 34.9293
R1909 B.n751 B.n377 34.9293
R1910 B.n751 B.n373 34.9293
R1911 B.n757 B.n373 34.9293
R1912 B.n757 B.n369 34.9293
R1913 B.n763 B.n369 34.9293
R1914 B.n763 B.n365 34.9293
R1915 B.n770 B.n365 34.9293
R1916 B.n770 B.n769 34.9293
R1917 B.n776 B.n358 34.9293
R1918 B.n783 B.n358 34.9293
R1919 B.n783 B.n354 34.9293
R1920 B.n789 B.n354 34.9293
R1921 B.n789 B.n4 34.9293
R1922 B.n890 B.n4 34.9293
R1923 B.n890 B.n889 34.9293
R1924 B.n889 B.n888 34.9293
R1925 B.n888 B.n8 34.9293
R1926 B.n882 B.n8 34.9293
R1927 B.n882 B.n881 34.9293
R1928 B.n881 B.n880 34.9293
R1929 B.n874 B.n18 34.9293
R1930 B.n874 B.n873 34.9293
R1931 B.n873 B.n872 34.9293
R1932 B.n872 B.n22 34.9293
R1933 B.n866 B.n22 34.9293
R1934 B.n866 B.n865 34.9293
R1935 B.n865 B.n864 34.9293
R1936 B.n864 B.n29 34.9293
R1937 B.n858 B.n29 34.9293
R1938 B.n858 B.n857 34.9293
R1939 B.n857 B.n856 34.9293
R1940 B.n856 B.n36 34.9293
R1941 B.n850 B.n36 34.9293
R1942 B.n849 B.n848 34.9293
R1943 B.n848 B.n43 34.9293
R1944 B.n842 B.n43 34.9293
R1945 B.n842 B.n841 34.9293
R1946 B.n841 B.n840 34.9293
R1947 B.n840 B.n50 34.9293
R1948 B.n834 B.n50 34.9293
R1949 B.n834 B.n833 34.9293
R1950 B.n121 B.n52 34.4981
R1951 B.n830 B.n829 34.4981
R1952 B.n706 B.n705 34.4981
R1953 B.n699 B.n403 34.4981
R1954 B.n776 B.t1 29.7927
R1955 B.n880 B.t0 29.7927
R1956 B.n733 B.t7 19.5195
R1957 B.n850 B.t3 19.5195
R1958 B B.n892 18.0485
R1959 B.n393 B.t7 15.4103
R1960 B.t3 B.n849 15.4103
R1961 B.n122 B.n121 10.6151
R1962 B.n125 B.n122 10.6151
R1963 B.n126 B.n125 10.6151
R1964 B.n129 B.n126 10.6151
R1965 B.n130 B.n129 10.6151
R1966 B.n133 B.n130 10.6151
R1967 B.n134 B.n133 10.6151
R1968 B.n137 B.n134 10.6151
R1969 B.n138 B.n137 10.6151
R1970 B.n141 B.n138 10.6151
R1971 B.n142 B.n141 10.6151
R1972 B.n145 B.n142 10.6151
R1973 B.n146 B.n145 10.6151
R1974 B.n149 B.n146 10.6151
R1975 B.n150 B.n149 10.6151
R1976 B.n153 B.n150 10.6151
R1977 B.n154 B.n153 10.6151
R1978 B.n157 B.n154 10.6151
R1979 B.n158 B.n157 10.6151
R1980 B.n161 B.n158 10.6151
R1981 B.n162 B.n161 10.6151
R1982 B.n165 B.n162 10.6151
R1983 B.n166 B.n165 10.6151
R1984 B.n169 B.n166 10.6151
R1985 B.n170 B.n169 10.6151
R1986 B.n173 B.n170 10.6151
R1987 B.n174 B.n173 10.6151
R1988 B.n177 B.n174 10.6151
R1989 B.n178 B.n177 10.6151
R1990 B.n181 B.n178 10.6151
R1991 B.n182 B.n181 10.6151
R1992 B.n185 B.n182 10.6151
R1993 B.n186 B.n185 10.6151
R1994 B.n189 B.n186 10.6151
R1995 B.n190 B.n189 10.6151
R1996 B.n193 B.n190 10.6151
R1997 B.n194 B.n193 10.6151
R1998 B.n197 B.n194 10.6151
R1999 B.n198 B.n197 10.6151
R2000 B.n201 B.n198 10.6151
R2001 B.n202 B.n201 10.6151
R2002 B.n205 B.n202 10.6151
R2003 B.n206 B.n205 10.6151
R2004 B.n209 B.n206 10.6151
R2005 B.n210 B.n209 10.6151
R2006 B.n213 B.n210 10.6151
R2007 B.n214 B.n213 10.6151
R2008 B.n217 B.n214 10.6151
R2009 B.n218 B.n217 10.6151
R2010 B.n221 B.n218 10.6151
R2011 B.n222 B.n221 10.6151
R2012 B.n225 B.n222 10.6151
R2013 B.n226 B.n225 10.6151
R2014 B.n230 B.n229 10.6151
R2015 B.n233 B.n230 10.6151
R2016 B.n234 B.n233 10.6151
R2017 B.n237 B.n234 10.6151
R2018 B.n238 B.n237 10.6151
R2019 B.n241 B.n238 10.6151
R2020 B.n242 B.n241 10.6151
R2021 B.n245 B.n242 10.6151
R2022 B.n250 B.n247 10.6151
R2023 B.n251 B.n250 10.6151
R2024 B.n254 B.n251 10.6151
R2025 B.n255 B.n254 10.6151
R2026 B.n258 B.n255 10.6151
R2027 B.n259 B.n258 10.6151
R2028 B.n262 B.n259 10.6151
R2029 B.n263 B.n262 10.6151
R2030 B.n266 B.n263 10.6151
R2031 B.n267 B.n266 10.6151
R2032 B.n270 B.n267 10.6151
R2033 B.n271 B.n270 10.6151
R2034 B.n274 B.n271 10.6151
R2035 B.n275 B.n274 10.6151
R2036 B.n278 B.n275 10.6151
R2037 B.n279 B.n278 10.6151
R2038 B.n282 B.n279 10.6151
R2039 B.n283 B.n282 10.6151
R2040 B.n286 B.n283 10.6151
R2041 B.n287 B.n286 10.6151
R2042 B.n290 B.n287 10.6151
R2043 B.n291 B.n290 10.6151
R2044 B.n294 B.n291 10.6151
R2045 B.n295 B.n294 10.6151
R2046 B.n298 B.n295 10.6151
R2047 B.n299 B.n298 10.6151
R2048 B.n302 B.n299 10.6151
R2049 B.n303 B.n302 10.6151
R2050 B.n306 B.n303 10.6151
R2051 B.n307 B.n306 10.6151
R2052 B.n310 B.n307 10.6151
R2053 B.n311 B.n310 10.6151
R2054 B.n314 B.n311 10.6151
R2055 B.n315 B.n314 10.6151
R2056 B.n318 B.n315 10.6151
R2057 B.n319 B.n318 10.6151
R2058 B.n322 B.n319 10.6151
R2059 B.n323 B.n322 10.6151
R2060 B.n326 B.n323 10.6151
R2061 B.n327 B.n326 10.6151
R2062 B.n330 B.n327 10.6151
R2063 B.n331 B.n330 10.6151
R2064 B.n334 B.n331 10.6151
R2065 B.n335 B.n334 10.6151
R2066 B.n338 B.n335 10.6151
R2067 B.n339 B.n338 10.6151
R2068 B.n342 B.n339 10.6151
R2069 B.n343 B.n342 10.6151
R2070 B.n346 B.n343 10.6151
R2071 B.n347 B.n346 10.6151
R2072 B.n350 B.n347 10.6151
R2073 B.n351 B.n350 10.6151
R2074 B.n830 B.n351 10.6151
R2075 B.n707 B.n706 10.6151
R2076 B.n707 B.n399 10.6151
R2077 B.n717 B.n399 10.6151
R2078 B.n718 B.n717 10.6151
R2079 B.n719 B.n718 10.6151
R2080 B.n719 B.n390 10.6151
R2081 B.n729 B.n390 10.6151
R2082 B.n730 B.n729 10.6151
R2083 B.n731 B.n730 10.6151
R2084 B.n731 B.n383 10.6151
R2085 B.n741 B.n383 10.6151
R2086 B.n742 B.n741 10.6151
R2087 B.n743 B.n742 10.6151
R2088 B.n743 B.n375 10.6151
R2089 B.n753 B.n375 10.6151
R2090 B.n754 B.n753 10.6151
R2091 B.n755 B.n754 10.6151
R2092 B.n755 B.n367 10.6151
R2093 B.n765 B.n367 10.6151
R2094 B.n766 B.n765 10.6151
R2095 B.n767 B.n766 10.6151
R2096 B.n767 B.n360 10.6151
R2097 B.n778 B.n360 10.6151
R2098 B.n779 B.n778 10.6151
R2099 B.n781 B.n779 10.6151
R2100 B.n781 B.n780 10.6151
R2101 B.n780 B.n352 10.6151
R2102 B.n792 B.n352 10.6151
R2103 B.n793 B.n792 10.6151
R2104 B.n794 B.n793 10.6151
R2105 B.n795 B.n794 10.6151
R2106 B.n797 B.n795 10.6151
R2107 B.n798 B.n797 10.6151
R2108 B.n799 B.n798 10.6151
R2109 B.n800 B.n799 10.6151
R2110 B.n802 B.n800 10.6151
R2111 B.n803 B.n802 10.6151
R2112 B.n804 B.n803 10.6151
R2113 B.n805 B.n804 10.6151
R2114 B.n807 B.n805 10.6151
R2115 B.n808 B.n807 10.6151
R2116 B.n809 B.n808 10.6151
R2117 B.n810 B.n809 10.6151
R2118 B.n812 B.n810 10.6151
R2119 B.n813 B.n812 10.6151
R2120 B.n814 B.n813 10.6151
R2121 B.n815 B.n814 10.6151
R2122 B.n817 B.n815 10.6151
R2123 B.n818 B.n817 10.6151
R2124 B.n819 B.n818 10.6151
R2125 B.n820 B.n819 10.6151
R2126 B.n822 B.n820 10.6151
R2127 B.n823 B.n822 10.6151
R2128 B.n824 B.n823 10.6151
R2129 B.n825 B.n824 10.6151
R2130 B.n827 B.n825 10.6151
R2131 B.n828 B.n827 10.6151
R2132 B.n829 B.n828 10.6151
R2133 B.n699 B.n698 10.6151
R2134 B.n698 B.n697 10.6151
R2135 B.n697 B.n696 10.6151
R2136 B.n696 B.n694 10.6151
R2137 B.n694 B.n691 10.6151
R2138 B.n691 B.n690 10.6151
R2139 B.n690 B.n687 10.6151
R2140 B.n687 B.n686 10.6151
R2141 B.n686 B.n683 10.6151
R2142 B.n683 B.n682 10.6151
R2143 B.n682 B.n679 10.6151
R2144 B.n679 B.n678 10.6151
R2145 B.n678 B.n675 10.6151
R2146 B.n675 B.n674 10.6151
R2147 B.n674 B.n671 10.6151
R2148 B.n671 B.n670 10.6151
R2149 B.n670 B.n667 10.6151
R2150 B.n667 B.n666 10.6151
R2151 B.n666 B.n663 10.6151
R2152 B.n663 B.n662 10.6151
R2153 B.n662 B.n659 10.6151
R2154 B.n659 B.n658 10.6151
R2155 B.n658 B.n655 10.6151
R2156 B.n655 B.n654 10.6151
R2157 B.n654 B.n651 10.6151
R2158 B.n651 B.n650 10.6151
R2159 B.n650 B.n647 10.6151
R2160 B.n647 B.n646 10.6151
R2161 B.n646 B.n643 10.6151
R2162 B.n643 B.n642 10.6151
R2163 B.n642 B.n639 10.6151
R2164 B.n639 B.n638 10.6151
R2165 B.n638 B.n635 10.6151
R2166 B.n635 B.n634 10.6151
R2167 B.n634 B.n631 10.6151
R2168 B.n631 B.n630 10.6151
R2169 B.n630 B.n627 10.6151
R2170 B.n627 B.n626 10.6151
R2171 B.n626 B.n623 10.6151
R2172 B.n623 B.n622 10.6151
R2173 B.n622 B.n619 10.6151
R2174 B.n619 B.n618 10.6151
R2175 B.n618 B.n615 10.6151
R2176 B.n615 B.n614 10.6151
R2177 B.n614 B.n611 10.6151
R2178 B.n611 B.n610 10.6151
R2179 B.n610 B.n607 10.6151
R2180 B.n607 B.n606 10.6151
R2181 B.n606 B.n603 10.6151
R2182 B.n603 B.n602 10.6151
R2183 B.n602 B.n599 10.6151
R2184 B.n599 B.n598 10.6151
R2185 B.n598 B.n595 10.6151
R2186 B.n593 B.n590 10.6151
R2187 B.n590 B.n589 10.6151
R2188 B.n589 B.n586 10.6151
R2189 B.n586 B.n585 10.6151
R2190 B.n585 B.n582 10.6151
R2191 B.n582 B.n581 10.6151
R2192 B.n581 B.n578 10.6151
R2193 B.n578 B.n577 10.6151
R2194 B.n574 B.n573 10.6151
R2195 B.n573 B.n570 10.6151
R2196 B.n570 B.n569 10.6151
R2197 B.n569 B.n566 10.6151
R2198 B.n566 B.n565 10.6151
R2199 B.n565 B.n562 10.6151
R2200 B.n562 B.n561 10.6151
R2201 B.n561 B.n558 10.6151
R2202 B.n558 B.n557 10.6151
R2203 B.n557 B.n554 10.6151
R2204 B.n554 B.n553 10.6151
R2205 B.n553 B.n550 10.6151
R2206 B.n550 B.n549 10.6151
R2207 B.n549 B.n546 10.6151
R2208 B.n546 B.n545 10.6151
R2209 B.n545 B.n542 10.6151
R2210 B.n542 B.n541 10.6151
R2211 B.n541 B.n538 10.6151
R2212 B.n538 B.n537 10.6151
R2213 B.n537 B.n534 10.6151
R2214 B.n534 B.n533 10.6151
R2215 B.n533 B.n530 10.6151
R2216 B.n530 B.n529 10.6151
R2217 B.n529 B.n526 10.6151
R2218 B.n526 B.n525 10.6151
R2219 B.n525 B.n522 10.6151
R2220 B.n522 B.n521 10.6151
R2221 B.n521 B.n518 10.6151
R2222 B.n518 B.n517 10.6151
R2223 B.n517 B.n514 10.6151
R2224 B.n514 B.n513 10.6151
R2225 B.n513 B.n510 10.6151
R2226 B.n510 B.n509 10.6151
R2227 B.n509 B.n506 10.6151
R2228 B.n506 B.n505 10.6151
R2229 B.n505 B.n502 10.6151
R2230 B.n502 B.n501 10.6151
R2231 B.n501 B.n498 10.6151
R2232 B.n498 B.n497 10.6151
R2233 B.n497 B.n494 10.6151
R2234 B.n494 B.n493 10.6151
R2235 B.n493 B.n490 10.6151
R2236 B.n490 B.n489 10.6151
R2237 B.n489 B.n486 10.6151
R2238 B.n486 B.n485 10.6151
R2239 B.n485 B.n482 10.6151
R2240 B.n482 B.n481 10.6151
R2241 B.n481 B.n478 10.6151
R2242 B.n478 B.n477 10.6151
R2243 B.n477 B.n474 10.6151
R2244 B.n474 B.n473 10.6151
R2245 B.n473 B.n407 10.6151
R2246 B.n705 B.n407 10.6151
R2247 B.n711 B.n403 10.6151
R2248 B.n712 B.n711 10.6151
R2249 B.n713 B.n712 10.6151
R2250 B.n713 B.n395 10.6151
R2251 B.n723 B.n395 10.6151
R2252 B.n724 B.n723 10.6151
R2253 B.n725 B.n724 10.6151
R2254 B.n725 B.n387 10.6151
R2255 B.n735 B.n387 10.6151
R2256 B.n736 B.n735 10.6151
R2257 B.n737 B.n736 10.6151
R2258 B.n737 B.n379 10.6151
R2259 B.n747 B.n379 10.6151
R2260 B.n748 B.n747 10.6151
R2261 B.n749 B.n748 10.6151
R2262 B.n749 B.n371 10.6151
R2263 B.n759 B.n371 10.6151
R2264 B.n760 B.n759 10.6151
R2265 B.n761 B.n760 10.6151
R2266 B.n761 B.n363 10.6151
R2267 B.n772 B.n363 10.6151
R2268 B.n773 B.n772 10.6151
R2269 B.n774 B.n773 10.6151
R2270 B.n774 B.n356 10.6151
R2271 B.n785 B.n356 10.6151
R2272 B.n786 B.n785 10.6151
R2273 B.n787 B.n786 10.6151
R2274 B.n787 B.n0 10.6151
R2275 B.n886 B.n1 10.6151
R2276 B.n886 B.n885 10.6151
R2277 B.n885 B.n884 10.6151
R2278 B.n884 B.n10 10.6151
R2279 B.n878 B.n10 10.6151
R2280 B.n878 B.n877 10.6151
R2281 B.n877 B.n876 10.6151
R2282 B.n876 B.n16 10.6151
R2283 B.n870 B.n16 10.6151
R2284 B.n870 B.n869 10.6151
R2285 B.n869 B.n868 10.6151
R2286 B.n868 B.n24 10.6151
R2287 B.n862 B.n24 10.6151
R2288 B.n862 B.n861 10.6151
R2289 B.n861 B.n860 10.6151
R2290 B.n860 B.n31 10.6151
R2291 B.n854 B.n31 10.6151
R2292 B.n854 B.n853 10.6151
R2293 B.n853 B.n852 10.6151
R2294 B.n852 B.n38 10.6151
R2295 B.n846 B.n38 10.6151
R2296 B.n846 B.n845 10.6151
R2297 B.n845 B.n844 10.6151
R2298 B.n844 B.n45 10.6151
R2299 B.n838 B.n45 10.6151
R2300 B.n838 B.n837 10.6151
R2301 B.n837 B.n836 10.6151
R2302 B.n836 B.n52 10.6151
R2303 B.n229 B.n119 6.5566
R2304 B.n246 B.n245 6.5566
R2305 B.n594 B.n593 6.5566
R2306 B.n577 B.n471 6.5566
R2307 B.n769 B.t1 5.13709
R2308 B.n18 B.t0 5.13709
R2309 B.n226 B.n119 4.05904
R2310 B.n247 B.n246 4.05904
R2311 B.n595 B.n594 4.05904
R2312 B.n574 B.n471 4.05904
R2313 B.n892 B.n0 2.81026
R2314 B.n892 B.n1 2.81026
R2315 VN VN.t0 208.297
R2316 VN VN.t1 159.425
R2317 VDD2.n173 VDD2.n89 289.615
R2318 VDD2.n84 VDD2.n0 289.615
R2319 VDD2.n174 VDD2.n173 185
R2320 VDD2.n172 VDD2.n171 185
R2321 VDD2.n93 VDD2.n92 185
R2322 VDD2.n166 VDD2.n165 185
R2323 VDD2.n164 VDD2.n95 185
R2324 VDD2.n163 VDD2.n162 185
R2325 VDD2.n98 VDD2.n96 185
R2326 VDD2.n157 VDD2.n156 185
R2327 VDD2.n155 VDD2.n154 185
R2328 VDD2.n102 VDD2.n101 185
R2329 VDD2.n149 VDD2.n148 185
R2330 VDD2.n147 VDD2.n146 185
R2331 VDD2.n106 VDD2.n105 185
R2332 VDD2.n141 VDD2.n140 185
R2333 VDD2.n139 VDD2.n138 185
R2334 VDD2.n110 VDD2.n109 185
R2335 VDD2.n133 VDD2.n132 185
R2336 VDD2.n131 VDD2.n130 185
R2337 VDD2.n114 VDD2.n113 185
R2338 VDD2.n125 VDD2.n124 185
R2339 VDD2.n123 VDD2.n122 185
R2340 VDD2.n118 VDD2.n117 185
R2341 VDD2.n28 VDD2.n27 185
R2342 VDD2.n33 VDD2.n32 185
R2343 VDD2.n35 VDD2.n34 185
R2344 VDD2.n24 VDD2.n23 185
R2345 VDD2.n41 VDD2.n40 185
R2346 VDD2.n43 VDD2.n42 185
R2347 VDD2.n20 VDD2.n19 185
R2348 VDD2.n49 VDD2.n48 185
R2349 VDD2.n51 VDD2.n50 185
R2350 VDD2.n16 VDD2.n15 185
R2351 VDD2.n57 VDD2.n56 185
R2352 VDD2.n59 VDD2.n58 185
R2353 VDD2.n12 VDD2.n11 185
R2354 VDD2.n65 VDD2.n64 185
R2355 VDD2.n67 VDD2.n66 185
R2356 VDD2.n8 VDD2.n7 185
R2357 VDD2.n74 VDD2.n73 185
R2358 VDD2.n75 VDD2.n6 185
R2359 VDD2.n77 VDD2.n76 185
R2360 VDD2.n4 VDD2.n3 185
R2361 VDD2.n83 VDD2.n82 185
R2362 VDD2.n85 VDD2.n84 185
R2363 VDD2.n119 VDD2.t1 147.659
R2364 VDD2.n29 VDD2.t0 147.659
R2365 VDD2.n173 VDD2.n172 104.615
R2366 VDD2.n172 VDD2.n92 104.615
R2367 VDD2.n165 VDD2.n92 104.615
R2368 VDD2.n165 VDD2.n164 104.615
R2369 VDD2.n164 VDD2.n163 104.615
R2370 VDD2.n163 VDD2.n96 104.615
R2371 VDD2.n156 VDD2.n96 104.615
R2372 VDD2.n156 VDD2.n155 104.615
R2373 VDD2.n155 VDD2.n101 104.615
R2374 VDD2.n148 VDD2.n101 104.615
R2375 VDD2.n148 VDD2.n147 104.615
R2376 VDD2.n147 VDD2.n105 104.615
R2377 VDD2.n140 VDD2.n105 104.615
R2378 VDD2.n140 VDD2.n139 104.615
R2379 VDD2.n139 VDD2.n109 104.615
R2380 VDD2.n132 VDD2.n109 104.615
R2381 VDD2.n132 VDD2.n131 104.615
R2382 VDD2.n131 VDD2.n113 104.615
R2383 VDD2.n124 VDD2.n113 104.615
R2384 VDD2.n124 VDD2.n123 104.615
R2385 VDD2.n123 VDD2.n117 104.615
R2386 VDD2.n33 VDD2.n27 104.615
R2387 VDD2.n34 VDD2.n33 104.615
R2388 VDD2.n34 VDD2.n23 104.615
R2389 VDD2.n41 VDD2.n23 104.615
R2390 VDD2.n42 VDD2.n41 104.615
R2391 VDD2.n42 VDD2.n19 104.615
R2392 VDD2.n49 VDD2.n19 104.615
R2393 VDD2.n50 VDD2.n49 104.615
R2394 VDD2.n50 VDD2.n15 104.615
R2395 VDD2.n57 VDD2.n15 104.615
R2396 VDD2.n58 VDD2.n57 104.615
R2397 VDD2.n58 VDD2.n11 104.615
R2398 VDD2.n65 VDD2.n11 104.615
R2399 VDD2.n66 VDD2.n65 104.615
R2400 VDD2.n66 VDD2.n7 104.615
R2401 VDD2.n74 VDD2.n7 104.615
R2402 VDD2.n75 VDD2.n74 104.615
R2403 VDD2.n76 VDD2.n75 104.615
R2404 VDD2.n76 VDD2.n3 104.615
R2405 VDD2.n83 VDD2.n3 104.615
R2406 VDD2.n84 VDD2.n83 104.615
R2407 VDD2.n178 VDD2.n88 93.7562
R2408 VDD2.t1 VDD2.n117 52.3082
R2409 VDD2.t0 VDD2.n27 52.3082
R2410 VDD2.n178 VDD2.n177 50.0278
R2411 VDD2.n119 VDD2.n118 15.6677
R2412 VDD2.n29 VDD2.n28 15.6677
R2413 VDD2.n166 VDD2.n95 13.1884
R2414 VDD2.n77 VDD2.n6 13.1884
R2415 VDD2.n167 VDD2.n93 12.8005
R2416 VDD2.n162 VDD2.n97 12.8005
R2417 VDD2.n122 VDD2.n121 12.8005
R2418 VDD2.n32 VDD2.n31 12.8005
R2419 VDD2.n73 VDD2.n72 12.8005
R2420 VDD2.n78 VDD2.n4 12.8005
R2421 VDD2.n171 VDD2.n170 12.0247
R2422 VDD2.n161 VDD2.n98 12.0247
R2423 VDD2.n125 VDD2.n116 12.0247
R2424 VDD2.n35 VDD2.n26 12.0247
R2425 VDD2.n71 VDD2.n8 12.0247
R2426 VDD2.n82 VDD2.n81 12.0247
R2427 VDD2.n174 VDD2.n91 11.249
R2428 VDD2.n158 VDD2.n157 11.249
R2429 VDD2.n126 VDD2.n114 11.249
R2430 VDD2.n36 VDD2.n24 11.249
R2431 VDD2.n68 VDD2.n67 11.249
R2432 VDD2.n85 VDD2.n2 11.249
R2433 VDD2.n175 VDD2.n89 10.4732
R2434 VDD2.n154 VDD2.n100 10.4732
R2435 VDD2.n130 VDD2.n129 10.4732
R2436 VDD2.n40 VDD2.n39 10.4732
R2437 VDD2.n64 VDD2.n10 10.4732
R2438 VDD2.n86 VDD2.n0 10.4732
R2439 VDD2.n153 VDD2.n102 9.69747
R2440 VDD2.n133 VDD2.n112 9.69747
R2441 VDD2.n43 VDD2.n22 9.69747
R2442 VDD2.n63 VDD2.n12 9.69747
R2443 VDD2.n177 VDD2.n176 9.45567
R2444 VDD2.n88 VDD2.n87 9.45567
R2445 VDD2.n145 VDD2.n144 9.3005
R2446 VDD2.n104 VDD2.n103 9.3005
R2447 VDD2.n151 VDD2.n150 9.3005
R2448 VDD2.n153 VDD2.n152 9.3005
R2449 VDD2.n100 VDD2.n99 9.3005
R2450 VDD2.n159 VDD2.n158 9.3005
R2451 VDD2.n161 VDD2.n160 9.3005
R2452 VDD2.n97 VDD2.n94 9.3005
R2453 VDD2.n176 VDD2.n175 9.3005
R2454 VDD2.n91 VDD2.n90 9.3005
R2455 VDD2.n170 VDD2.n169 9.3005
R2456 VDD2.n168 VDD2.n167 9.3005
R2457 VDD2.n143 VDD2.n142 9.3005
R2458 VDD2.n108 VDD2.n107 9.3005
R2459 VDD2.n137 VDD2.n136 9.3005
R2460 VDD2.n135 VDD2.n134 9.3005
R2461 VDD2.n112 VDD2.n111 9.3005
R2462 VDD2.n129 VDD2.n128 9.3005
R2463 VDD2.n127 VDD2.n126 9.3005
R2464 VDD2.n116 VDD2.n115 9.3005
R2465 VDD2.n121 VDD2.n120 9.3005
R2466 VDD2.n87 VDD2.n86 9.3005
R2467 VDD2.n2 VDD2.n1 9.3005
R2468 VDD2.n81 VDD2.n80 9.3005
R2469 VDD2.n79 VDD2.n78 9.3005
R2470 VDD2.n18 VDD2.n17 9.3005
R2471 VDD2.n47 VDD2.n46 9.3005
R2472 VDD2.n45 VDD2.n44 9.3005
R2473 VDD2.n22 VDD2.n21 9.3005
R2474 VDD2.n39 VDD2.n38 9.3005
R2475 VDD2.n37 VDD2.n36 9.3005
R2476 VDD2.n26 VDD2.n25 9.3005
R2477 VDD2.n31 VDD2.n30 9.3005
R2478 VDD2.n53 VDD2.n52 9.3005
R2479 VDD2.n55 VDD2.n54 9.3005
R2480 VDD2.n14 VDD2.n13 9.3005
R2481 VDD2.n61 VDD2.n60 9.3005
R2482 VDD2.n63 VDD2.n62 9.3005
R2483 VDD2.n10 VDD2.n9 9.3005
R2484 VDD2.n69 VDD2.n68 9.3005
R2485 VDD2.n71 VDD2.n70 9.3005
R2486 VDD2.n72 VDD2.n5 9.3005
R2487 VDD2.n150 VDD2.n149 8.92171
R2488 VDD2.n134 VDD2.n110 8.92171
R2489 VDD2.n44 VDD2.n20 8.92171
R2490 VDD2.n60 VDD2.n59 8.92171
R2491 VDD2.n146 VDD2.n104 8.14595
R2492 VDD2.n138 VDD2.n137 8.14595
R2493 VDD2.n48 VDD2.n47 8.14595
R2494 VDD2.n56 VDD2.n14 8.14595
R2495 VDD2.n145 VDD2.n106 7.3702
R2496 VDD2.n141 VDD2.n108 7.3702
R2497 VDD2.n51 VDD2.n18 7.3702
R2498 VDD2.n55 VDD2.n16 7.3702
R2499 VDD2.n142 VDD2.n106 6.59444
R2500 VDD2.n142 VDD2.n141 6.59444
R2501 VDD2.n52 VDD2.n51 6.59444
R2502 VDD2.n52 VDD2.n16 6.59444
R2503 VDD2.n146 VDD2.n145 5.81868
R2504 VDD2.n138 VDD2.n108 5.81868
R2505 VDD2.n48 VDD2.n18 5.81868
R2506 VDD2.n56 VDD2.n55 5.81868
R2507 VDD2.n149 VDD2.n104 5.04292
R2508 VDD2.n137 VDD2.n110 5.04292
R2509 VDD2.n47 VDD2.n20 5.04292
R2510 VDD2.n59 VDD2.n14 5.04292
R2511 VDD2.n120 VDD2.n119 4.38563
R2512 VDD2.n30 VDD2.n29 4.38563
R2513 VDD2.n150 VDD2.n102 4.26717
R2514 VDD2.n134 VDD2.n133 4.26717
R2515 VDD2.n44 VDD2.n43 4.26717
R2516 VDD2.n60 VDD2.n12 4.26717
R2517 VDD2.n177 VDD2.n89 3.49141
R2518 VDD2.n154 VDD2.n153 3.49141
R2519 VDD2.n130 VDD2.n112 3.49141
R2520 VDD2.n40 VDD2.n22 3.49141
R2521 VDD2.n64 VDD2.n63 3.49141
R2522 VDD2.n88 VDD2.n0 3.49141
R2523 VDD2.n175 VDD2.n174 2.71565
R2524 VDD2.n157 VDD2.n100 2.71565
R2525 VDD2.n129 VDD2.n114 2.71565
R2526 VDD2.n39 VDD2.n24 2.71565
R2527 VDD2.n67 VDD2.n10 2.71565
R2528 VDD2.n86 VDD2.n85 2.71565
R2529 VDD2.n171 VDD2.n91 1.93989
R2530 VDD2.n158 VDD2.n98 1.93989
R2531 VDD2.n126 VDD2.n125 1.93989
R2532 VDD2.n36 VDD2.n35 1.93989
R2533 VDD2.n68 VDD2.n8 1.93989
R2534 VDD2.n82 VDD2.n2 1.93989
R2535 VDD2.n170 VDD2.n93 1.16414
R2536 VDD2.n162 VDD2.n161 1.16414
R2537 VDD2.n122 VDD2.n116 1.16414
R2538 VDD2.n32 VDD2.n26 1.16414
R2539 VDD2.n73 VDD2.n71 1.16414
R2540 VDD2.n81 VDD2.n4 1.16414
R2541 VDD2 VDD2.n178 0.828086
R2542 VDD2.n167 VDD2.n166 0.388379
R2543 VDD2.n97 VDD2.n95 0.388379
R2544 VDD2.n121 VDD2.n118 0.388379
R2545 VDD2.n31 VDD2.n28 0.388379
R2546 VDD2.n72 VDD2.n6 0.388379
R2547 VDD2.n78 VDD2.n77 0.388379
R2548 VDD2.n176 VDD2.n90 0.155672
R2549 VDD2.n169 VDD2.n90 0.155672
R2550 VDD2.n169 VDD2.n168 0.155672
R2551 VDD2.n168 VDD2.n94 0.155672
R2552 VDD2.n160 VDD2.n94 0.155672
R2553 VDD2.n160 VDD2.n159 0.155672
R2554 VDD2.n159 VDD2.n99 0.155672
R2555 VDD2.n152 VDD2.n99 0.155672
R2556 VDD2.n152 VDD2.n151 0.155672
R2557 VDD2.n151 VDD2.n103 0.155672
R2558 VDD2.n144 VDD2.n103 0.155672
R2559 VDD2.n144 VDD2.n143 0.155672
R2560 VDD2.n143 VDD2.n107 0.155672
R2561 VDD2.n136 VDD2.n107 0.155672
R2562 VDD2.n136 VDD2.n135 0.155672
R2563 VDD2.n135 VDD2.n111 0.155672
R2564 VDD2.n128 VDD2.n111 0.155672
R2565 VDD2.n128 VDD2.n127 0.155672
R2566 VDD2.n127 VDD2.n115 0.155672
R2567 VDD2.n120 VDD2.n115 0.155672
R2568 VDD2.n30 VDD2.n25 0.155672
R2569 VDD2.n37 VDD2.n25 0.155672
R2570 VDD2.n38 VDD2.n37 0.155672
R2571 VDD2.n38 VDD2.n21 0.155672
R2572 VDD2.n45 VDD2.n21 0.155672
R2573 VDD2.n46 VDD2.n45 0.155672
R2574 VDD2.n46 VDD2.n17 0.155672
R2575 VDD2.n53 VDD2.n17 0.155672
R2576 VDD2.n54 VDD2.n53 0.155672
R2577 VDD2.n54 VDD2.n13 0.155672
R2578 VDD2.n61 VDD2.n13 0.155672
R2579 VDD2.n62 VDD2.n61 0.155672
R2580 VDD2.n62 VDD2.n9 0.155672
R2581 VDD2.n69 VDD2.n9 0.155672
R2582 VDD2.n70 VDD2.n69 0.155672
R2583 VDD2.n70 VDD2.n5 0.155672
R2584 VDD2.n79 VDD2.n5 0.155672
R2585 VDD2.n80 VDD2.n79 0.155672
R2586 VDD2.n80 VDD2.n1 0.155672
R2587 VDD2.n87 VDD2.n1 0.155672
C0 VP VTAIL 3.30061f
C1 VDD2 VN 3.76834f
C2 VP VDD2 0.360561f
C3 VDD2 VTAIL 6.29118f
C4 VDD1 VN 0.14875f
C5 VP VDD1 3.97729f
C6 VDD1 VTAIL 6.23646f
C7 VDD1 VDD2 0.752943f
C8 VP VN 6.52221f
C9 VN VTAIL 3.28632f
C10 VDD2 B 5.395097f
C11 VDD1 B 8.56177f
C12 VTAIL B 9.365909f
C13 VN B 12.31886f
C14 VP B 7.481413f
C15 VDD2.n0 B 0.027524f
C16 VDD2.n1 B 0.020162f
C17 VDD2.n2 B 0.010834f
C18 VDD2.n3 B 0.025608f
C19 VDD2.n4 B 0.011472f
C20 VDD2.n5 B 0.020162f
C21 VDD2.n6 B 0.011153f
C22 VDD2.n7 B 0.025608f
C23 VDD2.n8 B 0.011472f
C24 VDD2.n9 B 0.020162f
C25 VDD2.n10 B 0.010834f
C26 VDD2.n11 B 0.025608f
C27 VDD2.n12 B 0.011472f
C28 VDD2.n13 B 0.020162f
C29 VDD2.n14 B 0.010834f
C30 VDD2.n15 B 0.025608f
C31 VDD2.n16 B 0.011472f
C32 VDD2.n17 B 0.020162f
C33 VDD2.n18 B 0.010834f
C34 VDD2.n19 B 0.025608f
C35 VDD2.n20 B 0.011472f
C36 VDD2.n21 B 0.020162f
C37 VDD2.n22 B 0.010834f
C38 VDD2.n23 B 0.025608f
C39 VDD2.n24 B 0.011472f
C40 VDD2.n25 B 0.020162f
C41 VDD2.n26 B 0.010834f
C42 VDD2.n27 B 0.019206f
C43 VDD2.n28 B 0.015128f
C44 VDD2.t0 B 0.042304f
C45 VDD2.n29 B 0.137265f
C46 VDD2.n30 B 1.41712f
C47 VDD2.n31 B 0.010834f
C48 VDD2.n32 B 0.011472f
C49 VDD2.n33 B 0.025608f
C50 VDD2.n34 B 0.025608f
C51 VDD2.n35 B 0.011472f
C52 VDD2.n36 B 0.010834f
C53 VDD2.n37 B 0.020162f
C54 VDD2.n38 B 0.020162f
C55 VDD2.n39 B 0.010834f
C56 VDD2.n40 B 0.011472f
C57 VDD2.n41 B 0.025608f
C58 VDD2.n42 B 0.025608f
C59 VDD2.n43 B 0.011472f
C60 VDD2.n44 B 0.010834f
C61 VDD2.n45 B 0.020162f
C62 VDD2.n46 B 0.020162f
C63 VDD2.n47 B 0.010834f
C64 VDD2.n48 B 0.011472f
C65 VDD2.n49 B 0.025608f
C66 VDD2.n50 B 0.025608f
C67 VDD2.n51 B 0.011472f
C68 VDD2.n52 B 0.010834f
C69 VDD2.n53 B 0.020162f
C70 VDD2.n54 B 0.020162f
C71 VDD2.n55 B 0.010834f
C72 VDD2.n56 B 0.011472f
C73 VDD2.n57 B 0.025608f
C74 VDD2.n58 B 0.025608f
C75 VDD2.n59 B 0.011472f
C76 VDD2.n60 B 0.010834f
C77 VDD2.n61 B 0.020162f
C78 VDD2.n62 B 0.020162f
C79 VDD2.n63 B 0.010834f
C80 VDD2.n64 B 0.011472f
C81 VDD2.n65 B 0.025608f
C82 VDD2.n66 B 0.025608f
C83 VDD2.n67 B 0.011472f
C84 VDD2.n68 B 0.010834f
C85 VDD2.n69 B 0.020162f
C86 VDD2.n70 B 0.020162f
C87 VDD2.n71 B 0.010834f
C88 VDD2.n72 B 0.010834f
C89 VDD2.n73 B 0.011472f
C90 VDD2.n74 B 0.025608f
C91 VDD2.n75 B 0.025608f
C92 VDD2.n76 B 0.025608f
C93 VDD2.n77 B 0.011153f
C94 VDD2.n78 B 0.010834f
C95 VDD2.n79 B 0.020162f
C96 VDD2.n80 B 0.020162f
C97 VDD2.n81 B 0.010834f
C98 VDD2.n82 B 0.011472f
C99 VDD2.n83 B 0.025608f
C100 VDD2.n84 B 0.053994f
C101 VDD2.n85 B 0.011472f
C102 VDD2.n86 B 0.010834f
C103 VDD2.n87 B 0.048257f
C104 VDD2.n88 B 0.742526f
C105 VDD2.n89 B 0.027524f
C106 VDD2.n90 B 0.020162f
C107 VDD2.n91 B 0.010834f
C108 VDD2.n92 B 0.025608f
C109 VDD2.n93 B 0.011472f
C110 VDD2.n94 B 0.020162f
C111 VDD2.n95 B 0.011153f
C112 VDD2.n96 B 0.025608f
C113 VDD2.n97 B 0.010834f
C114 VDD2.n98 B 0.011472f
C115 VDD2.n99 B 0.020162f
C116 VDD2.n100 B 0.010834f
C117 VDD2.n101 B 0.025608f
C118 VDD2.n102 B 0.011472f
C119 VDD2.n103 B 0.020162f
C120 VDD2.n104 B 0.010834f
C121 VDD2.n105 B 0.025608f
C122 VDD2.n106 B 0.011472f
C123 VDD2.n107 B 0.020162f
C124 VDD2.n108 B 0.010834f
C125 VDD2.n109 B 0.025608f
C126 VDD2.n110 B 0.011472f
C127 VDD2.n111 B 0.020162f
C128 VDD2.n112 B 0.010834f
C129 VDD2.n113 B 0.025608f
C130 VDD2.n114 B 0.011472f
C131 VDD2.n115 B 0.020162f
C132 VDD2.n116 B 0.010834f
C133 VDD2.n117 B 0.019206f
C134 VDD2.n118 B 0.015128f
C135 VDD2.t1 B 0.042304f
C136 VDD2.n119 B 0.137265f
C137 VDD2.n120 B 1.41712f
C138 VDD2.n121 B 0.010834f
C139 VDD2.n122 B 0.011472f
C140 VDD2.n123 B 0.025608f
C141 VDD2.n124 B 0.025608f
C142 VDD2.n125 B 0.011472f
C143 VDD2.n126 B 0.010834f
C144 VDD2.n127 B 0.020162f
C145 VDD2.n128 B 0.020162f
C146 VDD2.n129 B 0.010834f
C147 VDD2.n130 B 0.011472f
C148 VDD2.n131 B 0.025608f
C149 VDD2.n132 B 0.025608f
C150 VDD2.n133 B 0.011472f
C151 VDD2.n134 B 0.010834f
C152 VDD2.n135 B 0.020162f
C153 VDD2.n136 B 0.020162f
C154 VDD2.n137 B 0.010834f
C155 VDD2.n138 B 0.011472f
C156 VDD2.n139 B 0.025608f
C157 VDD2.n140 B 0.025608f
C158 VDD2.n141 B 0.011472f
C159 VDD2.n142 B 0.010834f
C160 VDD2.n143 B 0.020162f
C161 VDD2.n144 B 0.020162f
C162 VDD2.n145 B 0.010834f
C163 VDD2.n146 B 0.011472f
C164 VDD2.n147 B 0.025608f
C165 VDD2.n148 B 0.025608f
C166 VDD2.n149 B 0.011472f
C167 VDD2.n150 B 0.010834f
C168 VDD2.n151 B 0.020162f
C169 VDD2.n152 B 0.020162f
C170 VDD2.n153 B 0.010834f
C171 VDD2.n154 B 0.011472f
C172 VDD2.n155 B 0.025608f
C173 VDD2.n156 B 0.025608f
C174 VDD2.n157 B 0.011472f
C175 VDD2.n158 B 0.010834f
C176 VDD2.n159 B 0.020162f
C177 VDD2.n160 B 0.020162f
C178 VDD2.n161 B 0.010834f
C179 VDD2.n162 B 0.011472f
C180 VDD2.n163 B 0.025608f
C181 VDD2.n164 B 0.025608f
C182 VDD2.n165 B 0.025608f
C183 VDD2.n166 B 0.011153f
C184 VDD2.n167 B 0.010834f
C185 VDD2.n168 B 0.020162f
C186 VDD2.n169 B 0.020162f
C187 VDD2.n170 B 0.010834f
C188 VDD2.n171 B 0.011472f
C189 VDD2.n172 B 0.025608f
C190 VDD2.n173 B 0.053994f
C191 VDD2.n174 B 0.011472f
C192 VDD2.n175 B 0.010834f
C193 VDD2.n176 B 0.048257f
C194 VDD2.n177 B 0.044023f
C195 VDD2.n178 B 2.91148f
C196 VN.t1 B 4.08289f
C197 VN.t0 B 4.71814f
C198 VDD1.n0 B 0.027593f
C199 VDD1.n1 B 0.020213f
C200 VDD1.n2 B 0.010862f
C201 VDD1.n3 B 0.025673f
C202 VDD1.n4 B 0.0115f
C203 VDD1.n5 B 0.020213f
C204 VDD1.n6 B 0.011181f
C205 VDD1.n7 B 0.025673f
C206 VDD1.n8 B 0.010862f
C207 VDD1.n9 B 0.0115f
C208 VDD1.n10 B 0.020213f
C209 VDD1.n11 B 0.010862f
C210 VDD1.n12 B 0.025673f
C211 VDD1.n13 B 0.0115f
C212 VDD1.n14 B 0.020213f
C213 VDD1.n15 B 0.010862f
C214 VDD1.n16 B 0.025673f
C215 VDD1.n17 B 0.0115f
C216 VDD1.n18 B 0.020213f
C217 VDD1.n19 B 0.010862f
C218 VDD1.n20 B 0.025673f
C219 VDD1.n21 B 0.0115f
C220 VDD1.n22 B 0.020213f
C221 VDD1.n23 B 0.010862f
C222 VDD1.n24 B 0.025673f
C223 VDD1.n25 B 0.0115f
C224 VDD1.n26 B 0.020213f
C225 VDD1.n27 B 0.010862f
C226 VDD1.n28 B 0.019255f
C227 VDD1.n29 B 0.015166f
C228 VDD1.t1 B 0.04241f
C229 VDD1.n30 B 0.13761f
C230 VDD1.n31 B 1.42068f
C231 VDD1.n32 B 0.010862f
C232 VDD1.n33 B 0.0115f
C233 VDD1.n34 B 0.025673f
C234 VDD1.n35 B 0.025673f
C235 VDD1.n36 B 0.0115f
C236 VDD1.n37 B 0.010862f
C237 VDD1.n38 B 0.020213f
C238 VDD1.n39 B 0.020213f
C239 VDD1.n40 B 0.010862f
C240 VDD1.n41 B 0.0115f
C241 VDD1.n42 B 0.025673f
C242 VDD1.n43 B 0.025673f
C243 VDD1.n44 B 0.0115f
C244 VDD1.n45 B 0.010862f
C245 VDD1.n46 B 0.020213f
C246 VDD1.n47 B 0.020213f
C247 VDD1.n48 B 0.010862f
C248 VDD1.n49 B 0.0115f
C249 VDD1.n50 B 0.025673f
C250 VDD1.n51 B 0.025673f
C251 VDD1.n52 B 0.0115f
C252 VDD1.n53 B 0.010862f
C253 VDD1.n54 B 0.020213f
C254 VDD1.n55 B 0.020213f
C255 VDD1.n56 B 0.010862f
C256 VDD1.n57 B 0.0115f
C257 VDD1.n58 B 0.025673f
C258 VDD1.n59 B 0.025673f
C259 VDD1.n60 B 0.0115f
C260 VDD1.n61 B 0.010862f
C261 VDD1.n62 B 0.020213f
C262 VDD1.n63 B 0.020213f
C263 VDD1.n64 B 0.010862f
C264 VDD1.n65 B 0.0115f
C265 VDD1.n66 B 0.025673f
C266 VDD1.n67 B 0.025673f
C267 VDD1.n68 B 0.0115f
C268 VDD1.n69 B 0.010862f
C269 VDD1.n70 B 0.020213f
C270 VDD1.n71 B 0.020213f
C271 VDD1.n72 B 0.010862f
C272 VDD1.n73 B 0.0115f
C273 VDD1.n74 B 0.025673f
C274 VDD1.n75 B 0.025673f
C275 VDD1.n76 B 0.025673f
C276 VDD1.n77 B 0.011181f
C277 VDD1.n78 B 0.010862f
C278 VDD1.n79 B 0.020213f
C279 VDD1.n80 B 0.020213f
C280 VDD1.n81 B 0.010862f
C281 VDD1.n82 B 0.0115f
C282 VDD1.n83 B 0.025673f
C283 VDD1.n84 B 0.05413f
C284 VDD1.n85 B 0.0115f
C285 VDD1.n86 B 0.010862f
C286 VDD1.n87 B 0.048378f
C287 VDD1.n88 B 0.045659f
C288 VDD1.n89 B 0.027593f
C289 VDD1.n90 B 0.020213f
C290 VDD1.n91 B 0.010862f
C291 VDD1.n92 B 0.025673f
C292 VDD1.n93 B 0.0115f
C293 VDD1.n94 B 0.020213f
C294 VDD1.n95 B 0.011181f
C295 VDD1.n96 B 0.025673f
C296 VDD1.n97 B 0.0115f
C297 VDD1.n98 B 0.020213f
C298 VDD1.n99 B 0.010862f
C299 VDD1.n100 B 0.025673f
C300 VDD1.n101 B 0.0115f
C301 VDD1.n102 B 0.020213f
C302 VDD1.n103 B 0.010862f
C303 VDD1.n104 B 0.025673f
C304 VDD1.n105 B 0.0115f
C305 VDD1.n106 B 0.020213f
C306 VDD1.n107 B 0.010862f
C307 VDD1.n108 B 0.025673f
C308 VDD1.n109 B 0.0115f
C309 VDD1.n110 B 0.020213f
C310 VDD1.n111 B 0.010862f
C311 VDD1.n112 B 0.025673f
C312 VDD1.n113 B 0.0115f
C313 VDD1.n114 B 0.020213f
C314 VDD1.n115 B 0.010862f
C315 VDD1.n116 B 0.019255f
C316 VDD1.n117 B 0.015166f
C317 VDD1.t0 B 0.04241f
C318 VDD1.n118 B 0.13761f
C319 VDD1.n119 B 1.42068f
C320 VDD1.n120 B 0.010862f
C321 VDD1.n121 B 0.0115f
C322 VDD1.n122 B 0.025673f
C323 VDD1.n123 B 0.025673f
C324 VDD1.n124 B 0.0115f
C325 VDD1.n125 B 0.010862f
C326 VDD1.n126 B 0.020213f
C327 VDD1.n127 B 0.020213f
C328 VDD1.n128 B 0.010862f
C329 VDD1.n129 B 0.0115f
C330 VDD1.n130 B 0.025673f
C331 VDD1.n131 B 0.025673f
C332 VDD1.n132 B 0.0115f
C333 VDD1.n133 B 0.010862f
C334 VDD1.n134 B 0.020213f
C335 VDD1.n135 B 0.020213f
C336 VDD1.n136 B 0.010862f
C337 VDD1.n137 B 0.0115f
C338 VDD1.n138 B 0.025673f
C339 VDD1.n139 B 0.025673f
C340 VDD1.n140 B 0.0115f
C341 VDD1.n141 B 0.010862f
C342 VDD1.n142 B 0.020213f
C343 VDD1.n143 B 0.020213f
C344 VDD1.n144 B 0.010862f
C345 VDD1.n145 B 0.0115f
C346 VDD1.n146 B 0.025673f
C347 VDD1.n147 B 0.025673f
C348 VDD1.n148 B 0.0115f
C349 VDD1.n149 B 0.010862f
C350 VDD1.n150 B 0.020213f
C351 VDD1.n151 B 0.020213f
C352 VDD1.n152 B 0.010862f
C353 VDD1.n153 B 0.0115f
C354 VDD1.n154 B 0.025673f
C355 VDD1.n155 B 0.025673f
C356 VDD1.n156 B 0.0115f
C357 VDD1.n157 B 0.010862f
C358 VDD1.n158 B 0.020213f
C359 VDD1.n159 B 0.020213f
C360 VDD1.n160 B 0.010862f
C361 VDD1.n161 B 0.010862f
C362 VDD1.n162 B 0.0115f
C363 VDD1.n163 B 0.025673f
C364 VDD1.n164 B 0.025673f
C365 VDD1.n165 B 0.025673f
C366 VDD1.n166 B 0.011181f
C367 VDD1.n167 B 0.010862f
C368 VDD1.n168 B 0.020213f
C369 VDD1.n169 B 0.020213f
C370 VDD1.n170 B 0.010862f
C371 VDD1.n171 B 0.0115f
C372 VDD1.n172 B 0.025673f
C373 VDD1.n173 B 0.05413f
C374 VDD1.n174 B 0.0115f
C375 VDD1.n175 B 0.010862f
C376 VDD1.n176 B 0.048378f
C377 VDD1.n177 B 0.791201f
C378 VTAIL.n0 B 0.027493f
C379 VTAIL.n1 B 0.02014f
C380 VTAIL.n2 B 0.010822f
C381 VTAIL.n3 B 0.02558f
C382 VTAIL.n4 B 0.011459f
C383 VTAIL.n5 B 0.02014f
C384 VTAIL.n6 B 0.011141f
C385 VTAIL.n7 B 0.02558f
C386 VTAIL.n8 B 0.011459f
C387 VTAIL.n9 B 0.02014f
C388 VTAIL.n10 B 0.010822f
C389 VTAIL.n11 B 0.02558f
C390 VTAIL.n12 B 0.011459f
C391 VTAIL.n13 B 0.02014f
C392 VTAIL.n14 B 0.010822f
C393 VTAIL.n15 B 0.02558f
C394 VTAIL.n16 B 0.011459f
C395 VTAIL.n17 B 0.02014f
C396 VTAIL.n18 B 0.010822f
C397 VTAIL.n19 B 0.02558f
C398 VTAIL.n20 B 0.011459f
C399 VTAIL.n21 B 0.02014f
C400 VTAIL.n22 B 0.010822f
C401 VTAIL.n23 B 0.02558f
C402 VTAIL.n24 B 0.011459f
C403 VTAIL.n25 B 0.02014f
C404 VTAIL.n26 B 0.010822f
C405 VTAIL.n27 B 0.019185f
C406 VTAIL.n28 B 0.015111f
C407 VTAIL.t2 B 0.042257f
C408 VTAIL.n29 B 0.137112f
C409 VTAIL.n30 B 1.41554f
C410 VTAIL.n31 B 0.010822f
C411 VTAIL.n32 B 0.011459f
C412 VTAIL.n33 B 0.02558f
C413 VTAIL.n34 B 0.02558f
C414 VTAIL.n35 B 0.011459f
C415 VTAIL.n36 B 0.010822f
C416 VTAIL.n37 B 0.02014f
C417 VTAIL.n38 B 0.02014f
C418 VTAIL.n39 B 0.010822f
C419 VTAIL.n40 B 0.011459f
C420 VTAIL.n41 B 0.02558f
C421 VTAIL.n42 B 0.02558f
C422 VTAIL.n43 B 0.011459f
C423 VTAIL.n44 B 0.010822f
C424 VTAIL.n45 B 0.02014f
C425 VTAIL.n46 B 0.02014f
C426 VTAIL.n47 B 0.010822f
C427 VTAIL.n48 B 0.011459f
C428 VTAIL.n49 B 0.02558f
C429 VTAIL.n50 B 0.02558f
C430 VTAIL.n51 B 0.011459f
C431 VTAIL.n52 B 0.010822f
C432 VTAIL.n53 B 0.02014f
C433 VTAIL.n54 B 0.02014f
C434 VTAIL.n55 B 0.010822f
C435 VTAIL.n56 B 0.011459f
C436 VTAIL.n57 B 0.02558f
C437 VTAIL.n58 B 0.02558f
C438 VTAIL.n59 B 0.011459f
C439 VTAIL.n60 B 0.010822f
C440 VTAIL.n61 B 0.02014f
C441 VTAIL.n62 B 0.02014f
C442 VTAIL.n63 B 0.010822f
C443 VTAIL.n64 B 0.011459f
C444 VTAIL.n65 B 0.02558f
C445 VTAIL.n66 B 0.02558f
C446 VTAIL.n67 B 0.011459f
C447 VTAIL.n68 B 0.010822f
C448 VTAIL.n69 B 0.02014f
C449 VTAIL.n70 B 0.02014f
C450 VTAIL.n71 B 0.010822f
C451 VTAIL.n72 B 0.010822f
C452 VTAIL.n73 B 0.011459f
C453 VTAIL.n74 B 0.02558f
C454 VTAIL.n75 B 0.02558f
C455 VTAIL.n76 B 0.02558f
C456 VTAIL.n77 B 0.011141f
C457 VTAIL.n78 B 0.010822f
C458 VTAIL.n79 B 0.02014f
C459 VTAIL.n80 B 0.02014f
C460 VTAIL.n81 B 0.010822f
C461 VTAIL.n82 B 0.011459f
C462 VTAIL.n83 B 0.02558f
C463 VTAIL.n84 B 0.053934f
C464 VTAIL.n85 B 0.011459f
C465 VTAIL.n86 B 0.010822f
C466 VTAIL.n87 B 0.048203f
C467 VTAIL.n88 B 0.03008f
C468 VTAIL.n89 B 1.67827f
C469 VTAIL.n90 B 0.027493f
C470 VTAIL.n91 B 0.02014f
C471 VTAIL.n92 B 0.010822f
C472 VTAIL.n93 B 0.02558f
C473 VTAIL.n94 B 0.011459f
C474 VTAIL.n95 B 0.02014f
C475 VTAIL.n96 B 0.011141f
C476 VTAIL.n97 B 0.02558f
C477 VTAIL.n98 B 0.010822f
C478 VTAIL.n99 B 0.011459f
C479 VTAIL.n100 B 0.02014f
C480 VTAIL.n101 B 0.010822f
C481 VTAIL.n102 B 0.02558f
C482 VTAIL.n103 B 0.011459f
C483 VTAIL.n104 B 0.02014f
C484 VTAIL.n105 B 0.010822f
C485 VTAIL.n106 B 0.02558f
C486 VTAIL.n107 B 0.011459f
C487 VTAIL.n108 B 0.02014f
C488 VTAIL.n109 B 0.010822f
C489 VTAIL.n110 B 0.02558f
C490 VTAIL.n111 B 0.011459f
C491 VTAIL.n112 B 0.02014f
C492 VTAIL.n113 B 0.010822f
C493 VTAIL.n114 B 0.02558f
C494 VTAIL.n115 B 0.011459f
C495 VTAIL.n116 B 0.02014f
C496 VTAIL.n117 B 0.010822f
C497 VTAIL.n118 B 0.019185f
C498 VTAIL.n119 B 0.015111f
C499 VTAIL.t1 B 0.042257f
C500 VTAIL.n120 B 0.137112f
C501 VTAIL.n121 B 1.41554f
C502 VTAIL.n122 B 0.010822f
C503 VTAIL.n123 B 0.011459f
C504 VTAIL.n124 B 0.02558f
C505 VTAIL.n125 B 0.02558f
C506 VTAIL.n126 B 0.011459f
C507 VTAIL.n127 B 0.010822f
C508 VTAIL.n128 B 0.02014f
C509 VTAIL.n129 B 0.02014f
C510 VTAIL.n130 B 0.010822f
C511 VTAIL.n131 B 0.011459f
C512 VTAIL.n132 B 0.02558f
C513 VTAIL.n133 B 0.02558f
C514 VTAIL.n134 B 0.011459f
C515 VTAIL.n135 B 0.010822f
C516 VTAIL.n136 B 0.02014f
C517 VTAIL.n137 B 0.02014f
C518 VTAIL.n138 B 0.010822f
C519 VTAIL.n139 B 0.011459f
C520 VTAIL.n140 B 0.02558f
C521 VTAIL.n141 B 0.02558f
C522 VTAIL.n142 B 0.011459f
C523 VTAIL.n143 B 0.010822f
C524 VTAIL.n144 B 0.02014f
C525 VTAIL.n145 B 0.02014f
C526 VTAIL.n146 B 0.010822f
C527 VTAIL.n147 B 0.011459f
C528 VTAIL.n148 B 0.02558f
C529 VTAIL.n149 B 0.02558f
C530 VTAIL.n150 B 0.011459f
C531 VTAIL.n151 B 0.010822f
C532 VTAIL.n152 B 0.02014f
C533 VTAIL.n153 B 0.02014f
C534 VTAIL.n154 B 0.010822f
C535 VTAIL.n155 B 0.011459f
C536 VTAIL.n156 B 0.02558f
C537 VTAIL.n157 B 0.02558f
C538 VTAIL.n158 B 0.011459f
C539 VTAIL.n159 B 0.010822f
C540 VTAIL.n160 B 0.02014f
C541 VTAIL.n161 B 0.02014f
C542 VTAIL.n162 B 0.010822f
C543 VTAIL.n163 B 0.011459f
C544 VTAIL.n164 B 0.02558f
C545 VTAIL.n165 B 0.02558f
C546 VTAIL.n166 B 0.02558f
C547 VTAIL.n167 B 0.011141f
C548 VTAIL.n168 B 0.010822f
C549 VTAIL.n169 B 0.02014f
C550 VTAIL.n170 B 0.02014f
C551 VTAIL.n171 B 0.010822f
C552 VTAIL.n172 B 0.011459f
C553 VTAIL.n173 B 0.02558f
C554 VTAIL.n174 B 0.053934f
C555 VTAIL.n175 B 0.011459f
C556 VTAIL.n176 B 0.010822f
C557 VTAIL.n177 B 0.048203f
C558 VTAIL.n178 B 0.03008f
C559 VTAIL.n179 B 1.72443f
C560 VTAIL.n180 B 0.027493f
C561 VTAIL.n181 B 0.02014f
C562 VTAIL.n182 B 0.010822f
C563 VTAIL.n183 B 0.02558f
C564 VTAIL.n184 B 0.011459f
C565 VTAIL.n185 B 0.02014f
C566 VTAIL.n186 B 0.011141f
C567 VTAIL.n187 B 0.02558f
C568 VTAIL.n188 B 0.010822f
C569 VTAIL.n189 B 0.011459f
C570 VTAIL.n190 B 0.02014f
C571 VTAIL.n191 B 0.010822f
C572 VTAIL.n192 B 0.02558f
C573 VTAIL.n193 B 0.011459f
C574 VTAIL.n194 B 0.02014f
C575 VTAIL.n195 B 0.010822f
C576 VTAIL.n196 B 0.02558f
C577 VTAIL.n197 B 0.011459f
C578 VTAIL.n198 B 0.02014f
C579 VTAIL.n199 B 0.010822f
C580 VTAIL.n200 B 0.02558f
C581 VTAIL.n201 B 0.011459f
C582 VTAIL.n202 B 0.02014f
C583 VTAIL.n203 B 0.010822f
C584 VTAIL.n204 B 0.02558f
C585 VTAIL.n205 B 0.011459f
C586 VTAIL.n206 B 0.02014f
C587 VTAIL.n207 B 0.010822f
C588 VTAIL.n208 B 0.019185f
C589 VTAIL.n209 B 0.015111f
C590 VTAIL.t3 B 0.042257f
C591 VTAIL.n210 B 0.137112f
C592 VTAIL.n211 B 1.41554f
C593 VTAIL.n212 B 0.010822f
C594 VTAIL.n213 B 0.011459f
C595 VTAIL.n214 B 0.02558f
C596 VTAIL.n215 B 0.02558f
C597 VTAIL.n216 B 0.011459f
C598 VTAIL.n217 B 0.010822f
C599 VTAIL.n218 B 0.02014f
C600 VTAIL.n219 B 0.02014f
C601 VTAIL.n220 B 0.010822f
C602 VTAIL.n221 B 0.011459f
C603 VTAIL.n222 B 0.02558f
C604 VTAIL.n223 B 0.02558f
C605 VTAIL.n224 B 0.011459f
C606 VTAIL.n225 B 0.010822f
C607 VTAIL.n226 B 0.02014f
C608 VTAIL.n227 B 0.02014f
C609 VTAIL.n228 B 0.010822f
C610 VTAIL.n229 B 0.011459f
C611 VTAIL.n230 B 0.02558f
C612 VTAIL.n231 B 0.02558f
C613 VTAIL.n232 B 0.011459f
C614 VTAIL.n233 B 0.010822f
C615 VTAIL.n234 B 0.02014f
C616 VTAIL.n235 B 0.02014f
C617 VTAIL.n236 B 0.010822f
C618 VTAIL.n237 B 0.011459f
C619 VTAIL.n238 B 0.02558f
C620 VTAIL.n239 B 0.02558f
C621 VTAIL.n240 B 0.011459f
C622 VTAIL.n241 B 0.010822f
C623 VTAIL.n242 B 0.02014f
C624 VTAIL.n243 B 0.02014f
C625 VTAIL.n244 B 0.010822f
C626 VTAIL.n245 B 0.011459f
C627 VTAIL.n246 B 0.02558f
C628 VTAIL.n247 B 0.02558f
C629 VTAIL.n248 B 0.011459f
C630 VTAIL.n249 B 0.010822f
C631 VTAIL.n250 B 0.02014f
C632 VTAIL.n251 B 0.02014f
C633 VTAIL.n252 B 0.010822f
C634 VTAIL.n253 B 0.011459f
C635 VTAIL.n254 B 0.02558f
C636 VTAIL.n255 B 0.02558f
C637 VTAIL.n256 B 0.02558f
C638 VTAIL.n257 B 0.011141f
C639 VTAIL.n258 B 0.010822f
C640 VTAIL.n259 B 0.02014f
C641 VTAIL.n260 B 0.02014f
C642 VTAIL.n261 B 0.010822f
C643 VTAIL.n262 B 0.011459f
C644 VTAIL.n263 B 0.02558f
C645 VTAIL.n264 B 0.053934f
C646 VTAIL.n265 B 0.011459f
C647 VTAIL.n266 B 0.010822f
C648 VTAIL.n267 B 0.048203f
C649 VTAIL.n268 B 0.03008f
C650 VTAIL.n269 B 1.52471f
C651 VTAIL.n270 B 0.027493f
C652 VTAIL.n271 B 0.02014f
C653 VTAIL.n272 B 0.010822f
C654 VTAIL.n273 B 0.02558f
C655 VTAIL.n274 B 0.011459f
C656 VTAIL.n275 B 0.02014f
C657 VTAIL.n276 B 0.011141f
C658 VTAIL.n277 B 0.02558f
C659 VTAIL.n278 B 0.011459f
C660 VTAIL.n279 B 0.02014f
C661 VTAIL.n280 B 0.010822f
C662 VTAIL.n281 B 0.02558f
C663 VTAIL.n282 B 0.011459f
C664 VTAIL.n283 B 0.02014f
C665 VTAIL.n284 B 0.010822f
C666 VTAIL.n285 B 0.02558f
C667 VTAIL.n286 B 0.011459f
C668 VTAIL.n287 B 0.02014f
C669 VTAIL.n288 B 0.010822f
C670 VTAIL.n289 B 0.02558f
C671 VTAIL.n290 B 0.011459f
C672 VTAIL.n291 B 0.02014f
C673 VTAIL.n292 B 0.010822f
C674 VTAIL.n293 B 0.02558f
C675 VTAIL.n294 B 0.011459f
C676 VTAIL.n295 B 0.02014f
C677 VTAIL.n296 B 0.010822f
C678 VTAIL.n297 B 0.019185f
C679 VTAIL.n298 B 0.015111f
C680 VTAIL.t0 B 0.042257f
C681 VTAIL.n299 B 0.137112f
C682 VTAIL.n300 B 1.41554f
C683 VTAIL.n301 B 0.010822f
C684 VTAIL.n302 B 0.011459f
C685 VTAIL.n303 B 0.02558f
C686 VTAIL.n304 B 0.02558f
C687 VTAIL.n305 B 0.011459f
C688 VTAIL.n306 B 0.010822f
C689 VTAIL.n307 B 0.02014f
C690 VTAIL.n308 B 0.02014f
C691 VTAIL.n309 B 0.010822f
C692 VTAIL.n310 B 0.011459f
C693 VTAIL.n311 B 0.02558f
C694 VTAIL.n312 B 0.02558f
C695 VTAIL.n313 B 0.011459f
C696 VTAIL.n314 B 0.010822f
C697 VTAIL.n315 B 0.02014f
C698 VTAIL.n316 B 0.02014f
C699 VTAIL.n317 B 0.010822f
C700 VTAIL.n318 B 0.011459f
C701 VTAIL.n319 B 0.02558f
C702 VTAIL.n320 B 0.02558f
C703 VTAIL.n321 B 0.011459f
C704 VTAIL.n322 B 0.010822f
C705 VTAIL.n323 B 0.02014f
C706 VTAIL.n324 B 0.02014f
C707 VTAIL.n325 B 0.010822f
C708 VTAIL.n326 B 0.011459f
C709 VTAIL.n327 B 0.02558f
C710 VTAIL.n328 B 0.02558f
C711 VTAIL.n329 B 0.011459f
C712 VTAIL.n330 B 0.010822f
C713 VTAIL.n331 B 0.02014f
C714 VTAIL.n332 B 0.02014f
C715 VTAIL.n333 B 0.010822f
C716 VTAIL.n334 B 0.011459f
C717 VTAIL.n335 B 0.02558f
C718 VTAIL.n336 B 0.02558f
C719 VTAIL.n337 B 0.011459f
C720 VTAIL.n338 B 0.010822f
C721 VTAIL.n339 B 0.02014f
C722 VTAIL.n340 B 0.02014f
C723 VTAIL.n341 B 0.010822f
C724 VTAIL.n342 B 0.010822f
C725 VTAIL.n343 B 0.011459f
C726 VTAIL.n344 B 0.02558f
C727 VTAIL.n345 B 0.02558f
C728 VTAIL.n346 B 0.02558f
C729 VTAIL.n347 B 0.011141f
C730 VTAIL.n348 B 0.010822f
C731 VTAIL.n349 B 0.02014f
C732 VTAIL.n350 B 0.02014f
C733 VTAIL.n351 B 0.010822f
C734 VTAIL.n352 B 0.011459f
C735 VTAIL.n353 B 0.02558f
C736 VTAIL.n354 B 0.053934f
C737 VTAIL.n355 B 0.011459f
C738 VTAIL.n356 B 0.010822f
C739 VTAIL.n357 B 0.048203f
C740 VTAIL.n358 B 0.03008f
C741 VTAIL.n359 B 1.44051f
C742 VP.t0 B 4.80061f
C743 VP.t1 B 4.14973f
C744 VP.n0 B 4.7594f
.ends

