* NGSPICE file created from diff_pair_sample_1673.ext - technology: sky130A

.subckt diff_pair_sample_1673 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t3 VP.t0 VTAIL.t6 w_n3166_n4838# sky130_fd_pr__pfet_01v8 ad=3.19275 pd=19.68 as=7.5465 ps=39.48 w=19.35 l=3.33
X1 VTAIL.t7 VP.t1 VDD1.t2 w_n3166_n4838# sky130_fd_pr__pfet_01v8 ad=7.5465 pd=39.48 as=3.19275 ps=19.68 w=19.35 l=3.33
X2 B.t11 B.t9 B.t10 w_n3166_n4838# sky130_fd_pr__pfet_01v8 ad=7.5465 pd=39.48 as=0 ps=0 w=19.35 l=3.33
X3 B.t8 B.t6 B.t7 w_n3166_n4838# sky130_fd_pr__pfet_01v8 ad=7.5465 pd=39.48 as=0 ps=0 w=19.35 l=3.33
X4 VTAIL.t5 VP.t2 VDD1.t1 w_n3166_n4838# sky130_fd_pr__pfet_01v8 ad=7.5465 pd=39.48 as=3.19275 ps=19.68 w=19.35 l=3.33
X5 VDD2.t3 VN.t0 VTAIL.t2 w_n3166_n4838# sky130_fd_pr__pfet_01v8 ad=3.19275 pd=19.68 as=7.5465 ps=39.48 w=19.35 l=3.33
X6 B.t5 B.t3 B.t4 w_n3166_n4838# sky130_fd_pr__pfet_01v8 ad=7.5465 pd=39.48 as=0 ps=0 w=19.35 l=3.33
X7 VDD1.t0 VP.t3 VTAIL.t4 w_n3166_n4838# sky130_fd_pr__pfet_01v8 ad=3.19275 pd=19.68 as=7.5465 ps=39.48 w=19.35 l=3.33
X8 B.t2 B.t0 B.t1 w_n3166_n4838# sky130_fd_pr__pfet_01v8 ad=7.5465 pd=39.48 as=0 ps=0 w=19.35 l=3.33
X9 VTAIL.t3 VN.t1 VDD2.t2 w_n3166_n4838# sky130_fd_pr__pfet_01v8 ad=7.5465 pd=39.48 as=3.19275 ps=19.68 w=19.35 l=3.33
X10 VTAIL.t1 VN.t2 VDD2.t1 w_n3166_n4838# sky130_fd_pr__pfet_01v8 ad=7.5465 pd=39.48 as=3.19275 ps=19.68 w=19.35 l=3.33
X11 VDD2.t0 VN.t3 VTAIL.t0 w_n3166_n4838# sky130_fd_pr__pfet_01v8 ad=3.19275 pd=19.68 as=7.5465 ps=39.48 w=19.35 l=3.33
R0 VP.n5 VP.t2 175.043
R1 VP.n5 VP.t3 173.917
R2 VP.n17 VP.n16 161.3
R3 VP.n15 VP.n1 161.3
R4 VP.n14 VP.n13 161.3
R5 VP.n12 VP.n2 161.3
R6 VP.n11 VP.n10 161.3
R7 VP.n9 VP.n3 161.3
R8 VP.n8 VP.n7 161.3
R9 VP.n4 VP.t1 140.042
R10 VP.n0 VP.t0 140.042
R11 VP.n6 VP.n4 73.9192
R12 VP.n18 VP.n0 73.9192
R13 VP.n6 VP.n5 56.6561
R14 VP.n10 VP.n2 40.4934
R15 VP.n14 VP.n2 40.4934
R16 VP.n9 VP.n8 24.4675
R17 VP.n10 VP.n9 24.4675
R18 VP.n15 VP.n14 24.4675
R19 VP.n16 VP.n15 24.4675
R20 VP.n8 VP.n4 16.1487
R21 VP.n16 VP.n0 16.1487
R22 VP.n7 VP.n6 0.354971
R23 VP.n18 VP.n17 0.354971
R24 VP VP.n18 0.26696
R25 VP.n7 VP.n3 0.189894
R26 VP.n11 VP.n3 0.189894
R27 VP.n12 VP.n11 0.189894
R28 VP.n13 VP.n12 0.189894
R29 VP.n13 VP.n1 0.189894
R30 VP.n17 VP.n1 0.189894
R31 VTAIL.n5 VTAIL.t5 53.8268
R32 VTAIL.n4 VTAIL.t2 53.8268
R33 VTAIL.n3 VTAIL.t1 53.8268
R34 VTAIL.n7 VTAIL.t0 53.8265
R35 VTAIL.n0 VTAIL.t3 53.8265
R36 VTAIL.n1 VTAIL.t6 53.8265
R37 VTAIL.n2 VTAIL.t7 53.8265
R38 VTAIL.n6 VTAIL.t4 53.8265
R39 VTAIL.n7 VTAIL.n6 32.2031
R40 VTAIL.n3 VTAIL.n2 32.2031
R41 VTAIL.n4 VTAIL.n3 3.15567
R42 VTAIL.n6 VTAIL.n5 3.15567
R43 VTAIL.n2 VTAIL.n1 3.15567
R44 VTAIL VTAIL.n0 1.63628
R45 VTAIL VTAIL.n7 1.5199
R46 VTAIL.n5 VTAIL.n4 0.470328
R47 VTAIL.n1 VTAIL.n0 0.470328
R48 VDD1 VDD1.n1 119.212
R49 VDD1 VDD1.n0 68.8837
R50 VDD1.n0 VDD1.t1 1.68034
R51 VDD1.n0 VDD1.t0 1.68034
R52 VDD1.n1 VDD1.t2 1.68034
R53 VDD1.n1 VDD1.t3 1.68034
R54 B.n491 B.n136 585
R55 B.n490 B.n489 585
R56 B.n488 B.n137 585
R57 B.n487 B.n486 585
R58 B.n485 B.n138 585
R59 B.n484 B.n483 585
R60 B.n482 B.n139 585
R61 B.n481 B.n480 585
R62 B.n479 B.n140 585
R63 B.n478 B.n477 585
R64 B.n476 B.n141 585
R65 B.n475 B.n474 585
R66 B.n473 B.n142 585
R67 B.n472 B.n471 585
R68 B.n470 B.n143 585
R69 B.n469 B.n468 585
R70 B.n467 B.n144 585
R71 B.n466 B.n465 585
R72 B.n464 B.n145 585
R73 B.n463 B.n462 585
R74 B.n461 B.n146 585
R75 B.n460 B.n459 585
R76 B.n458 B.n147 585
R77 B.n457 B.n456 585
R78 B.n455 B.n148 585
R79 B.n454 B.n453 585
R80 B.n452 B.n149 585
R81 B.n451 B.n450 585
R82 B.n449 B.n150 585
R83 B.n448 B.n447 585
R84 B.n446 B.n151 585
R85 B.n445 B.n444 585
R86 B.n443 B.n152 585
R87 B.n442 B.n441 585
R88 B.n440 B.n153 585
R89 B.n439 B.n438 585
R90 B.n437 B.n154 585
R91 B.n436 B.n435 585
R92 B.n434 B.n155 585
R93 B.n433 B.n432 585
R94 B.n431 B.n156 585
R95 B.n430 B.n429 585
R96 B.n428 B.n157 585
R97 B.n427 B.n426 585
R98 B.n425 B.n158 585
R99 B.n424 B.n423 585
R100 B.n422 B.n159 585
R101 B.n421 B.n420 585
R102 B.n419 B.n160 585
R103 B.n418 B.n417 585
R104 B.n416 B.n161 585
R105 B.n415 B.n414 585
R106 B.n413 B.n162 585
R107 B.n412 B.n411 585
R108 B.n410 B.n163 585
R109 B.n409 B.n408 585
R110 B.n407 B.n164 585
R111 B.n406 B.n405 585
R112 B.n404 B.n165 585
R113 B.n403 B.n402 585
R114 B.n401 B.n166 585
R115 B.n400 B.n399 585
R116 B.n398 B.n167 585
R117 B.n397 B.n396 585
R118 B.n392 B.n168 585
R119 B.n391 B.n390 585
R120 B.n389 B.n169 585
R121 B.n388 B.n387 585
R122 B.n386 B.n170 585
R123 B.n385 B.n384 585
R124 B.n383 B.n171 585
R125 B.n382 B.n381 585
R126 B.n380 B.n172 585
R127 B.n378 B.n377 585
R128 B.n376 B.n175 585
R129 B.n375 B.n374 585
R130 B.n373 B.n176 585
R131 B.n372 B.n371 585
R132 B.n370 B.n177 585
R133 B.n369 B.n368 585
R134 B.n367 B.n178 585
R135 B.n366 B.n365 585
R136 B.n364 B.n179 585
R137 B.n363 B.n362 585
R138 B.n361 B.n180 585
R139 B.n360 B.n359 585
R140 B.n358 B.n181 585
R141 B.n357 B.n356 585
R142 B.n355 B.n182 585
R143 B.n354 B.n353 585
R144 B.n352 B.n183 585
R145 B.n351 B.n350 585
R146 B.n349 B.n184 585
R147 B.n348 B.n347 585
R148 B.n346 B.n185 585
R149 B.n345 B.n344 585
R150 B.n343 B.n186 585
R151 B.n342 B.n341 585
R152 B.n340 B.n187 585
R153 B.n339 B.n338 585
R154 B.n337 B.n188 585
R155 B.n336 B.n335 585
R156 B.n334 B.n189 585
R157 B.n333 B.n332 585
R158 B.n331 B.n190 585
R159 B.n330 B.n329 585
R160 B.n328 B.n191 585
R161 B.n327 B.n326 585
R162 B.n325 B.n192 585
R163 B.n324 B.n323 585
R164 B.n322 B.n193 585
R165 B.n321 B.n320 585
R166 B.n319 B.n194 585
R167 B.n318 B.n317 585
R168 B.n316 B.n195 585
R169 B.n315 B.n314 585
R170 B.n313 B.n196 585
R171 B.n312 B.n311 585
R172 B.n310 B.n197 585
R173 B.n309 B.n308 585
R174 B.n307 B.n198 585
R175 B.n306 B.n305 585
R176 B.n304 B.n199 585
R177 B.n303 B.n302 585
R178 B.n301 B.n200 585
R179 B.n300 B.n299 585
R180 B.n298 B.n201 585
R181 B.n297 B.n296 585
R182 B.n295 B.n202 585
R183 B.n294 B.n293 585
R184 B.n292 B.n203 585
R185 B.n291 B.n290 585
R186 B.n289 B.n204 585
R187 B.n288 B.n287 585
R188 B.n286 B.n205 585
R189 B.n285 B.n284 585
R190 B.n493 B.n492 585
R191 B.n494 B.n135 585
R192 B.n496 B.n495 585
R193 B.n497 B.n134 585
R194 B.n499 B.n498 585
R195 B.n500 B.n133 585
R196 B.n502 B.n501 585
R197 B.n503 B.n132 585
R198 B.n505 B.n504 585
R199 B.n506 B.n131 585
R200 B.n508 B.n507 585
R201 B.n509 B.n130 585
R202 B.n511 B.n510 585
R203 B.n512 B.n129 585
R204 B.n514 B.n513 585
R205 B.n515 B.n128 585
R206 B.n517 B.n516 585
R207 B.n518 B.n127 585
R208 B.n520 B.n519 585
R209 B.n521 B.n126 585
R210 B.n523 B.n522 585
R211 B.n524 B.n125 585
R212 B.n526 B.n525 585
R213 B.n527 B.n124 585
R214 B.n529 B.n528 585
R215 B.n530 B.n123 585
R216 B.n532 B.n531 585
R217 B.n533 B.n122 585
R218 B.n535 B.n534 585
R219 B.n536 B.n121 585
R220 B.n538 B.n537 585
R221 B.n539 B.n120 585
R222 B.n541 B.n540 585
R223 B.n542 B.n119 585
R224 B.n544 B.n543 585
R225 B.n545 B.n118 585
R226 B.n547 B.n546 585
R227 B.n548 B.n117 585
R228 B.n550 B.n549 585
R229 B.n551 B.n116 585
R230 B.n553 B.n552 585
R231 B.n554 B.n115 585
R232 B.n556 B.n555 585
R233 B.n557 B.n114 585
R234 B.n559 B.n558 585
R235 B.n560 B.n113 585
R236 B.n562 B.n561 585
R237 B.n563 B.n112 585
R238 B.n565 B.n564 585
R239 B.n566 B.n111 585
R240 B.n568 B.n567 585
R241 B.n569 B.n110 585
R242 B.n571 B.n570 585
R243 B.n572 B.n109 585
R244 B.n574 B.n573 585
R245 B.n575 B.n108 585
R246 B.n577 B.n576 585
R247 B.n578 B.n107 585
R248 B.n580 B.n579 585
R249 B.n581 B.n106 585
R250 B.n583 B.n582 585
R251 B.n584 B.n105 585
R252 B.n586 B.n585 585
R253 B.n587 B.n104 585
R254 B.n589 B.n588 585
R255 B.n590 B.n103 585
R256 B.n592 B.n591 585
R257 B.n593 B.n102 585
R258 B.n595 B.n594 585
R259 B.n596 B.n101 585
R260 B.n598 B.n597 585
R261 B.n599 B.n100 585
R262 B.n601 B.n600 585
R263 B.n602 B.n99 585
R264 B.n604 B.n603 585
R265 B.n605 B.n98 585
R266 B.n607 B.n606 585
R267 B.n608 B.n97 585
R268 B.n610 B.n609 585
R269 B.n611 B.n96 585
R270 B.n613 B.n612 585
R271 B.n614 B.n95 585
R272 B.n819 B.n22 585
R273 B.n818 B.n817 585
R274 B.n816 B.n23 585
R275 B.n815 B.n814 585
R276 B.n813 B.n24 585
R277 B.n812 B.n811 585
R278 B.n810 B.n25 585
R279 B.n809 B.n808 585
R280 B.n807 B.n26 585
R281 B.n806 B.n805 585
R282 B.n804 B.n27 585
R283 B.n803 B.n802 585
R284 B.n801 B.n28 585
R285 B.n800 B.n799 585
R286 B.n798 B.n29 585
R287 B.n797 B.n796 585
R288 B.n795 B.n30 585
R289 B.n794 B.n793 585
R290 B.n792 B.n31 585
R291 B.n791 B.n790 585
R292 B.n789 B.n32 585
R293 B.n788 B.n787 585
R294 B.n786 B.n33 585
R295 B.n785 B.n784 585
R296 B.n783 B.n34 585
R297 B.n782 B.n781 585
R298 B.n780 B.n35 585
R299 B.n779 B.n778 585
R300 B.n777 B.n36 585
R301 B.n776 B.n775 585
R302 B.n774 B.n37 585
R303 B.n773 B.n772 585
R304 B.n771 B.n38 585
R305 B.n770 B.n769 585
R306 B.n768 B.n39 585
R307 B.n767 B.n766 585
R308 B.n765 B.n40 585
R309 B.n764 B.n763 585
R310 B.n762 B.n41 585
R311 B.n761 B.n760 585
R312 B.n759 B.n42 585
R313 B.n758 B.n757 585
R314 B.n756 B.n43 585
R315 B.n755 B.n754 585
R316 B.n753 B.n44 585
R317 B.n752 B.n751 585
R318 B.n750 B.n45 585
R319 B.n749 B.n748 585
R320 B.n747 B.n46 585
R321 B.n746 B.n745 585
R322 B.n744 B.n47 585
R323 B.n743 B.n742 585
R324 B.n741 B.n48 585
R325 B.n740 B.n739 585
R326 B.n738 B.n49 585
R327 B.n737 B.n736 585
R328 B.n735 B.n50 585
R329 B.n734 B.n733 585
R330 B.n732 B.n51 585
R331 B.n731 B.n730 585
R332 B.n729 B.n52 585
R333 B.n728 B.n727 585
R334 B.n726 B.n53 585
R335 B.n724 B.n723 585
R336 B.n722 B.n56 585
R337 B.n721 B.n720 585
R338 B.n719 B.n57 585
R339 B.n718 B.n717 585
R340 B.n716 B.n58 585
R341 B.n715 B.n714 585
R342 B.n713 B.n59 585
R343 B.n712 B.n711 585
R344 B.n710 B.n60 585
R345 B.n709 B.n708 585
R346 B.n707 B.n61 585
R347 B.n706 B.n705 585
R348 B.n704 B.n65 585
R349 B.n703 B.n702 585
R350 B.n701 B.n66 585
R351 B.n700 B.n699 585
R352 B.n698 B.n67 585
R353 B.n697 B.n696 585
R354 B.n695 B.n68 585
R355 B.n694 B.n693 585
R356 B.n692 B.n69 585
R357 B.n691 B.n690 585
R358 B.n689 B.n70 585
R359 B.n688 B.n687 585
R360 B.n686 B.n71 585
R361 B.n685 B.n684 585
R362 B.n683 B.n72 585
R363 B.n682 B.n681 585
R364 B.n680 B.n73 585
R365 B.n679 B.n678 585
R366 B.n677 B.n74 585
R367 B.n676 B.n675 585
R368 B.n674 B.n75 585
R369 B.n673 B.n672 585
R370 B.n671 B.n76 585
R371 B.n670 B.n669 585
R372 B.n668 B.n77 585
R373 B.n667 B.n666 585
R374 B.n665 B.n78 585
R375 B.n664 B.n663 585
R376 B.n662 B.n79 585
R377 B.n661 B.n660 585
R378 B.n659 B.n80 585
R379 B.n658 B.n657 585
R380 B.n656 B.n81 585
R381 B.n655 B.n654 585
R382 B.n653 B.n82 585
R383 B.n652 B.n651 585
R384 B.n650 B.n83 585
R385 B.n649 B.n648 585
R386 B.n647 B.n84 585
R387 B.n646 B.n645 585
R388 B.n644 B.n85 585
R389 B.n643 B.n642 585
R390 B.n641 B.n86 585
R391 B.n640 B.n639 585
R392 B.n638 B.n87 585
R393 B.n637 B.n636 585
R394 B.n635 B.n88 585
R395 B.n634 B.n633 585
R396 B.n632 B.n89 585
R397 B.n631 B.n630 585
R398 B.n629 B.n90 585
R399 B.n628 B.n627 585
R400 B.n626 B.n91 585
R401 B.n625 B.n624 585
R402 B.n623 B.n92 585
R403 B.n622 B.n621 585
R404 B.n620 B.n93 585
R405 B.n619 B.n618 585
R406 B.n617 B.n94 585
R407 B.n616 B.n615 585
R408 B.n821 B.n820 585
R409 B.n822 B.n21 585
R410 B.n824 B.n823 585
R411 B.n825 B.n20 585
R412 B.n827 B.n826 585
R413 B.n828 B.n19 585
R414 B.n830 B.n829 585
R415 B.n831 B.n18 585
R416 B.n833 B.n832 585
R417 B.n834 B.n17 585
R418 B.n836 B.n835 585
R419 B.n837 B.n16 585
R420 B.n839 B.n838 585
R421 B.n840 B.n15 585
R422 B.n842 B.n841 585
R423 B.n843 B.n14 585
R424 B.n845 B.n844 585
R425 B.n846 B.n13 585
R426 B.n848 B.n847 585
R427 B.n849 B.n12 585
R428 B.n851 B.n850 585
R429 B.n852 B.n11 585
R430 B.n854 B.n853 585
R431 B.n855 B.n10 585
R432 B.n857 B.n856 585
R433 B.n858 B.n9 585
R434 B.n860 B.n859 585
R435 B.n861 B.n8 585
R436 B.n863 B.n862 585
R437 B.n864 B.n7 585
R438 B.n866 B.n865 585
R439 B.n867 B.n6 585
R440 B.n869 B.n868 585
R441 B.n870 B.n5 585
R442 B.n872 B.n871 585
R443 B.n873 B.n4 585
R444 B.n875 B.n874 585
R445 B.n876 B.n3 585
R446 B.n878 B.n877 585
R447 B.n879 B.n0 585
R448 B.n2 B.n1 585
R449 B.n226 B.n225 585
R450 B.n228 B.n227 585
R451 B.n229 B.n224 585
R452 B.n231 B.n230 585
R453 B.n232 B.n223 585
R454 B.n234 B.n233 585
R455 B.n235 B.n222 585
R456 B.n237 B.n236 585
R457 B.n238 B.n221 585
R458 B.n240 B.n239 585
R459 B.n241 B.n220 585
R460 B.n243 B.n242 585
R461 B.n244 B.n219 585
R462 B.n246 B.n245 585
R463 B.n247 B.n218 585
R464 B.n249 B.n248 585
R465 B.n250 B.n217 585
R466 B.n252 B.n251 585
R467 B.n253 B.n216 585
R468 B.n255 B.n254 585
R469 B.n256 B.n215 585
R470 B.n258 B.n257 585
R471 B.n259 B.n214 585
R472 B.n261 B.n260 585
R473 B.n262 B.n213 585
R474 B.n264 B.n263 585
R475 B.n265 B.n212 585
R476 B.n267 B.n266 585
R477 B.n268 B.n211 585
R478 B.n270 B.n269 585
R479 B.n271 B.n210 585
R480 B.n273 B.n272 585
R481 B.n274 B.n209 585
R482 B.n276 B.n275 585
R483 B.n277 B.n208 585
R484 B.n279 B.n278 585
R485 B.n280 B.n207 585
R486 B.n282 B.n281 585
R487 B.n283 B.n206 585
R488 B.n285 B.n206 487.695
R489 B.n493 B.n136 487.695
R490 B.n615 B.n614 487.695
R491 B.n820 B.n819 487.695
R492 B.n173 B.t3 348.976
R493 B.n393 B.t0 348.976
R494 B.n62 B.t9 348.976
R495 B.n54 B.t6 348.976
R496 B.n881 B.n880 256.663
R497 B.n880 B.n879 235.042
R498 B.n880 B.n2 235.042
R499 B.n393 B.t1 183.073
R500 B.n62 B.t11 183.073
R501 B.n173 B.t4 183.048
R502 B.n54 B.t8 183.048
R503 B.n286 B.n285 163.367
R504 B.n287 B.n286 163.367
R505 B.n287 B.n204 163.367
R506 B.n291 B.n204 163.367
R507 B.n292 B.n291 163.367
R508 B.n293 B.n292 163.367
R509 B.n293 B.n202 163.367
R510 B.n297 B.n202 163.367
R511 B.n298 B.n297 163.367
R512 B.n299 B.n298 163.367
R513 B.n299 B.n200 163.367
R514 B.n303 B.n200 163.367
R515 B.n304 B.n303 163.367
R516 B.n305 B.n304 163.367
R517 B.n305 B.n198 163.367
R518 B.n309 B.n198 163.367
R519 B.n310 B.n309 163.367
R520 B.n311 B.n310 163.367
R521 B.n311 B.n196 163.367
R522 B.n315 B.n196 163.367
R523 B.n316 B.n315 163.367
R524 B.n317 B.n316 163.367
R525 B.n317 B.n194 163.367
R526 B.n321 B.n194 163.367
R527 B.n322 B.n321 163.367
R528 B.n323 B.n322 163.367
R529 B.n323 B.n192 163.367
R530 B.n327 B.n192 163.367
R531 B.n328 B.n327 163.367
R532 B.n329 B.n328 163.367
R533 B.n329 B.n190 163.367
R534 B.n333 B.n190 163.367
R535 B.n334 B.n333 163.367
R536 B.n335 B.n334 163.367
R537 B.n335 B.n188 163.367
R538 B.n339 B.n188 163.367
R539 B.n340 B.n339 163.367
R540 B.n341 B.n340 163.367
R541 B.n341 B.n186 163.367
R542 B.n345 B.n186 163.367
R543 B.n346 B.n345 163.367
R544 B.n347 B.n346 163.367
R545 B.n347 B.n184 163.367
R546 B.n351 B.n184 163.367
R547 B.n352 B.n351 163.367
R548 B.n353 B.n352 163.367
R549 B.n353 B.n182 163.367
R550 B.n357 B.n182 163.367
R551 B.n358 B.n357 163.367
R552 B.n359 B.n358 163.367
R553 B.n359 B.n180 163.367
R554 B.n363 B.n180 163.367
R555 B.n364 B.n363 163.367
R556 B.n365 B.n364 163.367
R557 B.n365 B.n178 163.367
R558 B.n369 B.n178 163.367
R559 B.n370 B.n369 163.367
R560 B.n371 B.n370 163.367
R561 B.n371 B.n176 163.367
R562 B.n375 B.n176 163.367
R563 B.n376 B.n375 163.367
R564 B.n377 B.n376 163.367
R565 B.n377 B.n172 163.367
R566 B.n382 B.n172 163.367
R567 B.n383 B.n382 163.367
R568 B.n384 B.n383 163.367
R569 B.n384 B.n170 163.367
R570 B.n388 B.n170 163.367
R571 B.n389 B.n388 163.367
R572 B.n390 B.n389 163.367
R573 B.n390 B.n168 163.367
R574 B.n397 B.n168 163.367
R575 B.n398 B.n397 163.367
R576 B.n399 B.n398 163.367
R577 B.n399 B.n166 163.367
R578 B.n403 B.n166 163.367
R579 B.n404 B.n403 163.367
R580 B.n405 B.n404 163.367
R581 B.n405 B.n164 163.367
R582 B.n409 B.n164 163.367
R583 B.n410 B.n409 163.367
R584 B.n411 B.n410 163.367
R585 B.n411 B.n162 163.367
R586 B.n415 B.n162 163.367
R587 B.n416 B.n415 163.367
R588 B.n417 B.n416 163.367
R589 B.n417 B.n160 163.367
R590 B.n421 B.n160 163.367
R591 B.n422 B.n421 163.367
R592 B.n423 B.n422 163.367
R593 B.n423 B.n158 163.367
R594 B.n427 B.n158 163.367
R595 B.n428 B.n427 163.367
R596 B.n429 B.n428 163.367
R597 B.n429 B.n156 163.367
R598 B.n433 B.n156 163.367
R599 B.n434 B.n433 163.367
R600 B.n435 B.n434 163.367
R601 B.n435 B.n154 163.367
R602 B.n439 B.n154 163.367
R603 B.n440 B.n439 163.367
R604 B.n441 B.n440 163.367
R605 B.n441 B.n152 163.367
R606 B.n445 B.n152 163.367
R607 B.n446 B.n445 163.367
R608 B.n447 B.n446 163.367
R609 B.n447 B.n150 163.367
R610 B.n451 B.n150 163.367
R611 B.n452 B.n451 163.367
R612 B.n453 B.n452 163.367
R613 B.n453 B.n148 163.367
R614 B.n457 B.n148 163.367
R615 B.n458 B.n457 163.367
R616 B.n459 B.n458 163.367
R617 B.n459 B.n146 163.367
R618 B.n463 B.n146 163.367
R619 B.n464 B.n463 163.367
R620 B.n465 B.n464 163.367
R621 B.n465 B.n144 163.367
R622 B.n469 B.n144 163.367
R623 B.n470 B.n469 163.367
R624 B.n471 B.n470 163.367
R625 B.n471 B.n142 163.367
R626 B.n475 B.n142 163.367
R627 B.n476 B.n475 163.367
R628 B.n477 B.n476 163.367
R629 B.n477 B.n140 163.367
R630 B.n481 B.n140 163.367
R631 B.n482 B.n481 163.367
R632 B.n483 B.n482 163.367
R633 B.n483 B.n138 163.367
R634 B.n487 B.n138 163.367
R635 B.n488 B.n487 163.367
R636 B.n489 B.n488 163.367
R637 B.n489 B.n136 163.367
R638 B.n614 B.n613 163.367
R639 B.n613 B.n96 163.367
R640 B.n609 B.n96 163.367
R641 B.n609 B.n608 163.367
R642 B.n608 B.n607 163.367
R643 B.n607 B.n98 163.367
R644 B.n603 B.n98 163.367
R645 B.n603 B.n602 163.367
R646 B.n602 B.n601 163.367
R647 B.n601 B.n100 163.367
R648 B.n597 B.n100 163.367
R649 B.n597 B.n596 163.367
R650 B.n596 B.n595 163.367
R651 B.n595 B.n102 163.367
R652 B.n591 B.n102 163.367
R653 B.n591 B.n590 163.367
R654 B.n590 B.n589 163.367
R655 B.n589 B.n104 163.367
R656 B.n585 B.n104 163.367
R657 B.n585 B.n584 163.367
R658 B.n584 B.n583 163.367
R659 B.n583 B.n106 163.367
R660 B.n579 B.n106 163.367
R661 B.n579 B.n578 163.367
R662 B.n578 B.n577 163.367
R663 B.n577 B.n108 163.367
R664 B.n573 B.n108 163.367
R665 B.n573 B.n572 163.367
R666 B.n572 B.n571 163.367
R667 B.n571 B.n110 163.367
R668 B.n567 B.n110 163.367
R669 B.n567 B.n566 163.367
R670 B.n566 B.n565 163.367
R671 B.n565 B.n112 163.367
R672 B.n561 B.n112 163.367
R673 B.n561 B.n560 163.367
R674 B.n560 B.n559 163.367
R675 B.n559 B.n114 163.367
R676 B.n555 B.n114 163.367
R677 B.n555 B.n554 163.367
R678 B.n554 B.n553 163.367
R679 B.n553 B.n116 163.367
R680 B.n549 B.n116 163.367
R681 B.n549 B.n548 163.367
R682 B.n548 B.n547 163.367
R683 B.n547 B.n118 163.367
R684 B.n543 B.n118 163.367
R685 B.n543 B.n542 163.367
R686 B.n542 B.n541 163.367
R687 B.n541 B.n120 163.367
R688 B.n537 B.n120 163.367
R689 B.n537 B.n536 163.367
R690 B.n536 B.n535 163.367
R691 B.n535 B.n122 163.367
R692 B.n531 B.n122 163.367
R693 B.n531 B.n530 163.367
R694 B.n530 B.n529 163.367
R695 B.n529 B.n124 163.367
R696 B.n525 B.n124 163.367
R697 B.n525 B.n524 163.367
R698 B.n524 B.n523 163.367
R699 B.n523 B.n126 163.367
R700 B.n519 B.n126 163.367
R701 B.n519 B.n518 163.367
R702 B.n518 B.n517 163.367
R703 B.n517 B.n128 163.367
R704 B.n513 B.n128 163.367
R705 B.n513 B.n512 163.367
R706 B.n512 B.n511 163.367
R707 B.n511 B.n130 163.367
R708 B.n507 B.n130 163.367
R709 B.n507 B.n506 163.367
R710 B.n506 B.n505 163.367
R711 B.n505 B.n132 163.367
R712 B.n501 B.n132 163.367
R713 B.n501 B.n500 163.367
R714 B.n500 B.n499 163.367
R715 B.n499 B.n134 163.367
R716 B.n495 B.n134 163.367
R717 B.n495 B.n494 163.367
R718 B.n494 B.n493 163.367
R719 B.n819 B.n818 163.367
R720 B.n818 B.n23 163.367
R721 B.n814 B.n23 163.367
R722 B.n814 B.n813 163.367
R723 B.n813 B.n812 163.367
R724 B.n812 B.n25 163.367
R725 B.n808 B.n25 163.367
R726 B.n808 B.n807 163.367
R727 B.n807 B.n806 163.367
R728 B.n806 B.n27 163.367
R729 B.n802 B.n27 163.367
R730 B.n802 B.n801 163.367
R731 B.n801 B.n800 163.367
R732 B.n800 B.n29 163.367
R733 B.n796 B.n29 163.367
R734 B.n796 B.n795 163.367
R735 B.n795 B.n794 163.367
R736 B.n794 B.n31 163.367
R737 B.n790 B.n31 163.367
R738 B.n790 B.n789 163.367
R739 B.n789 B.n788 163.367
R740 B.n788 B.n33 163.367
R741 B.n784 B.n33 163.367
R742 B.n784 B.n783 163.367
R743 B.n783 B.n782 163.367
R744 B.n782 B.n35 163.367
R745 B.n778 B.n35 163.367
R746 B.n778 B.n777 163.367
R747 B.n777 B.n776 163.367
R748 B.n776 B.n37 163.367
R749 B.n772 B.n37 163.367
R750 B.n772 B.n771 163.367
R751 B.n771 B.n770 163.367
R752 B.n770 B.n39 163.367
R753 B.n766 B.n39 163.367
R754 B.n766 B.n765 163.367
R755 B.n765 B.n764 163.367
R756 B.n764 B.n41 163.367
R757 B.n760 B.n41 163.367
R758 B.n760 B.n759 163.367
R759 B.n759 B.n758 163.367
R760 B.n758 B.n43 163.367
R761 B.n754 B.n43 163.367
R762 B.n754 B.n753 163.367
R763 B.n753 B.n752 163.367
R764 B.n752 B.n45 163.367
R765 B.n748 B.n45 163.367
R766 B.n748 B.n747 163.367
R767 B.n747 B.n746 163.367
R768 B.n746 B.n47 163.367
R769 B.n742 B.n47 163.367
R770 B.n742 B.n741 163.367
R771 B.n741 B.n740 163.367
R772 B.n740 B.n49 163.367
R773 B.n736 B.n49 163.367
R774 B.n736 B.n735 163.367
R775 B.n735 B.n734 163.367
R776 B.n734 B.n51 163.367
R777 B.n730 B.n51 163.367
R778 B.n730 B.n729 163.367
R779 B.n729 B.n728 163.367
R780 B.n728 B.n53 163.367
R781 B.n723 B.n53 163.367
R782 B.n723 B.n722 163.367
R783 B.n722 B.n721 163.367
R784 B.n721 B.n57 163.367
R785 B.n717 B.n57 163.367
R786 B.n717 B.n716 163.367
R787 B.n716 B.n715 163.367
R788 B.n715 B.n59 163.367
R789 B.n711 B.n59 163.367
R790 B.n711 B.n710 163.367
R791 B.n710 B.n709 163.367
R792 B.n709 B.n61 163.367
R793 B.n705 B.n61 163.367
R794 B.n705 B.n704 163.367
R795 B.n704 B.n703 163.367
R796 B.n703 B.n66 163.367
R797 B.n699 B.n66 163.367
R798 B.n699 B.n698 163.367
R799 B.n698 B.n697 163.367
R800 B.n697 B.n68 163.367
R801 B.n693 B.n68 163.367
R802 B.n693 B.n692 163.367
R803 B.n692 B.n691 163.367
R804 B.n691 B.n70 163.367
R805 B.n687 B.n70 163.367
R806 B.n687 B.n686 163.367
R807 B.n686 B.n685 163.367
R808 B.n685 B.n72 163.367
R809 B.n681 B.n72 163.367
R810 B.n681 B.n680 163.367
R811 B.n680 B.n679 163.367
R812 B.n679 B.n74 163.367
R813 B.n675 B.n74 163.367
R814 B.n675 B.n674 163.367
R815 B.n674 B.n673 163.367
R816 B.n673 B.n76 163.367
R817 B.n669 B.n76 163.367
R818 B.n669 B.n668 163.367
R819 B.n668 B.n667 163.367
R820 B.n667 B.n78 163.367
R821 B.n663 B.n78 163.367
R822 B.n663 B.n662 163.367
R823 B.n662 B.n661 163.367
R824 B.n661 B.n80 163.367
R825 B.n657 B.n80 163.367
R826 B.n657 B.n656 163.367
R827 B.n656 B.n655 163.367
R828 B.n655 B.n82 163.367
R829 B.n651 B.n82 163.367
R830 B.n651 B.n650 163.367
R831 B.n650 B.n649 163.367
R832 B.n649 B.n84 163.367
R833 B.n645 B.n84 163.367
R834 B.n645 B.n644 163.367
R835 B.n644 B.n643 163.367
R836 B.n643 B.n86 163.367
R837 B.n639 B.n86 163.367
R838 B.n639 B.n638 163.367
R839 B.n638 B.n637 163.367
R840 B.n637 B.n88 163.367
R841 B.n633 B.n88 163.367
R842 B.n633 B.n632 163.367
R843 B.n632 B.n631 163.367
R844 B.n631 B.n90 163.367
R845 B.n627 B.n90 163.367
R846 B.n627 B.n626 163.367
R847 B.n626 B.n625 163.367
R848 B.n625 B.n92 163.367
R849 B.n621 B.n92 163.367
R850 B.n621 B.n620 163.367
R851 B.n620 B.n619 163.367
R852 B.n619 B.n94 163.367
R853 B.n615 B.n94 163.367
R854 B.n820 B.n21 163.367
R855 B.n824 B.n21 163.367
R856 B.n825 B.n824 163.367
R857 B.n826 B.n825 163.367
R858 B.n826 B.n19 163.367
R859 B.n830 B.n19 163.367
R860 B.n831 B.n830 163.367
R861 B.n832 B.n831 163.367
R862 B.n832 B.n17 163.367
R863 B.n836 B.n17 163.367
R864 B.n837 B.n836 163.367
R865 B.n838 B.n837 163.367
R866 B.n838 B.n15 163.367
R867 B.n842 B.n15 163.367
R868 B.n843 B.n842 163.367
R869 B.n844 B.n843 163.367
R870 B.n844 B.n13 163.367
R871 B.n848 B.n13 163.367
R872 B.n849 B.n848 163.367
R873 B.n850 B.n849 163.367
R874 B.n850 B.n11 163.367
R875 B.n854 B.n11 163.367
R876 B.n855 B.n854 163.367
R877 B.n856 B.n855 163.367
R878 B.n856 B.n9 163.367
R879 B.n860 B.n9 163.367
R880 B.n861 B.n860 163.367
R881 B.n862 B.n861 163.367
R882 B.n862 B.n7 163.367
R883 B.n866 B.n7 163.367
R884 B.n867 B.n866 163.367
R885 B.n868 B.n867 163.367
R886 B.n868 B.n5 163.367
R887 B.n872 B.n5 163.367
R888 B.n873 B.n872 163.367
R889 B.n874 B.n873 163.367
R890 B.n874 B.n3 163.367
R891 B.n878 B.n3 163.367
R892 B.n879 B.n878 163.367
R893 B.n226 B.n2 163.367
R894 B.n227 B.n226 163.367
R895 B.n227 B.n224 163.367
R896 B.n231 B.n224 163.367
R897 B.n232 B.n231 163.367
R898 B.n233 B.n232 163.367
R899 B.n233 B.n222 163.367
R900 B.n237 B.n222 163.367
R901 B.n238 B.n237 163.367
R902 B.n239 B.n238 163.367
R903 B.n239 B.n220 163.367
R904 B.n243 B.n220 163.367
R905 B.n244 B.n243 163.367
R906 B.n245 B.n244 163.367
R907 B.n245 B.n218 163.367
R908 B.n249 B.n218 163.367
R909 B.n250 B.n249 163.367
R910 B.n251 B.n250 163.367
R911 B.n251 B.n216 163.367
R912 B.n255 B.n216 163.367
R913 B.n256 B.n255 163.367
R914 B.n257 B.n256 163.367
R915 B.n257 B.n214 163.367
R916 B.n261 B.n214 163.367
R917 B.n262 B.n261 163.367
R918 B.n263 B.n262 163.367
R919 B.n263 B.n212 163.367
R920 B.n267 B.n212 163.367
R921 B.n268 B.n267 163.367
R922 B.n269 B.n268 163.367
R923 B.n269 B.n210 163.367
R924 B.n273 B.n210 163.367
R925 B.n274 B.n273 163.367
R926 B.n275 B.n274 163.367
R927 B.n275 B.n208 163.367
R928 B.n279 B.n208 163.367
R929 B.n280 B.n279 163.367
R930 B.n281 B.n280 163.367
R931 B.n281 B.n206 163.367
R932 B.n394 B.t2 112.091
R933 B.n63 B.t10 112.091
R934 B.n174 B.t5 112.067
R935 B.n55 B.t7 112.067
R936 B.n174 B.n173 70.9823
R937 B.n394 B.n393 70.9823
R938 B.n63 B.n62 70.9823
R939 B.n55 B.n54 70.9823
R940 B.n379 B.n174 59.5399
R941 B.n395 B.n394 59.5399
R942 B.n64 B.n63 59.5399
R943 B.n725 B.n55 59.5399
R944 B.n821 B.n22 31.6883
R945 B.n616 B.n95 31.6883
R946 B.n492 B.n491 31.6883
R947 B.n284 B.n283 31.6883
R948 B B.n881 18.0485
R949 B.n822 B.n821 10.6151
R950 B.n823 B.n822 10.6151
R951 B.n823 B.n20 10.6151
R952 B.n827 B.n20 10.6151
R953 B.n828 B.n827 10.6151
R954 B.n829 B.n828 10.6151
R955 B.n829 B.n18 10.6151
R956 B.n833 B.n18 10.6151
R957 B.n834 B.n833 10.6151
R958 B.n835 B.n834 10.6151
R959 B.n835 B.n16 10.6151
R960 B.n839 B.n16 10.6151
R961 B.n840 B.n839 10.6151
R962 B.n841 B.n840 10.6151
R963 B.n841 B.n14 10.6151
R964 B.n845 B.n14 10.6151
R965 B.n846 B.n845 10.6151
R966 B.n847 B.n846 10.6151
R967 B.n847 B.n12 10.6151
R968 B.n851 B.n12 10.6151
R969 B.n852 B.n851 10.6151
R970 B.n853 B.n852 10.6151
R971 B.n853 B.n10 10.6151
R972 B.n857 B.n10 10.6151
R973 B.n858 B.n857 10.6151
R974 B.n859 B.n858 10.6151
R975 B.n859 B.n8 10.6151
R976 B.n863 B.n8 10.6151
R977 B.n864 B.n863 10.6151
R978 B.n865 B.n864 10.6151
R979 B.n865 B.n6 10.6151
R980 B.n869 B.n6 10.6151
R981 B.n870 B.n869 10.6151
R982 B.n871 B.n870 10.6151
R983 B.n871 B.n4 10.6151
R984 B.n875 B.n4 10.6151
R985 B.n876 B.n875 10.6151
R986 B.n877 B.n876 10.6151
R987 B.n877 B.n0 10.6151
R988 B.n817 B.n22 10.6151
R989 B.n817 B.n816 10.6151
R990 B.n816 B.n815 10.6151
R991 B.n815 B.n24 10.6151
R992 B.n811 B.n24 10.6151
R993 B.n811 B.n810 10.6151
R994 B.n810 B.n809 10.6151
R995 B.n809 B.n26 10.6151
R996 B.n805 B.n26 10.6151
R997 B.n805 B.n804 10.6151
R998 B.n804 B.n803 10.6151
R999 B.n803 B.n28 10.6151
R1000 B.n799 B.n28 10.6151
R1001 B.n799 B.n798 10.6151
R1002 B.n798 B.n797 10.6151
R1003 B.n797 B.n30 10.6151
R1004 B.n793 B.n30 10.6151
R1005 B.n793 B.n792 10.6151
R1006 B.n792 B.n791 10.6151
R1007 B.n791 B.n32 10.6151
R1008 B.n787 B.n32 10.6151
R1009 B.n787 B.n786 10.6151
R1010 B.n786 B.n785 10.6151
R1011 B.n785 B.n34 10.6151
R1012 B.n781 B.n34 10.6151
R1013 B.n781 B.n780 10.6151
R1014 B.n780 B.n779 10.6151
R1015 B.n779 B.n36 10.6151
R1016 B.n775 B.n36 10.6151
R1017 B.n775 B.n774 10.6151
R1018 B.n774 B.n773 10.6151
R1019 B.n773 B.n38 10.6151
R1020 B.n769 B.n38 10.6151
R1021 B.n769 B.n768 10.6151
R1022 B.n768 B.n767 10.6151
R1023 B.n767 B.n40 10.6151
R1024 B.n763 B.n40 10.6151
R1025 B.n763 B.n762 10.6151
R1026 B.n762 B.n761 10.6151
R1027 B.n761 B.n42 10.6151
R1028 B.n757 B.n42 10.6151
R1029 B.n757 B.n756 10.6151
R1030 B.n756 B.n755 10.6151
R1031 B.n755 B.n44 10.6151
R1032 B.n751 B.n44 10.6151
R1033 B.n751 B.n750 10.6151
R1034 B.n750 B.n749 10.6151
R1035 B.n749 B.n46 10.6151
R1036 B.n745 B.n46 10.6151
R1037 B.n745 B.n744 10.6151
R1038 B.n744 B.n743 10.6151
R1039 B.n743 B.n48 10.6151
R1040 B.n739 B.n48 10.6151
R1041 B.n739 B.n738 10.6151
R1042 B.n738 B.n737 10.6151
R1043 B.n737 B.n50 10.6151
R1044 B.n733 B.n50 10.6151
R1045 B.n733 B.n732 10.6151
R1046 B.n732 B.n731 10.6151
R1047 B.n731 B.n52 10.6151
R1048 B.n727 B.n52 10.6151
R1049 B.n727 B.n726 10.6151
R1050 B.n724 B.n56 10.6151
R1051 B.n720 B.n56 10.6151
R1052 B.n720 B.n719 10.6151
R1053 B.n719 B.n718 10.6151
R1054 B.n718 B.n58 10.6151
R1055 B.n714 B.n58 10.6151
R1056 B.n714 B.n713 10.6151
R1057 B.n713 B.n712 10.6151
R1058 B.n712 B.n60 10.6151
R1059 B.n708 B.n707 10.6151
R1060 B.n707 B.n706 10.6151
R1061 B.n706 B.n65 10.6151
R1062 B.n702 B.n65 10.6151
R1063 B.n702 B.n701 10.6151
R1064 B.n701 B.n700 10.6151
R1065 B.n700 B.n67 10.6151
R1066 B.n696 B.n67 10.6151
R1067 B.n696 B.n695 10.6151
R1068 B.n695 B.n694 10.6151
R1069 B.n694 B.n69 10.6151
R1070 B.n690 B.n69 10.6151
R1071 B.n690 B.n689 10.6151
R1072 B.n689 B.n688 10.6151
R1073 B.n688 B.n71 10.6151
R1074 B.n684 B.n71 10.6151
R1075 B.n684 B.n683 10.6151
R1076 B.n683 B.n682 10.6151
R1077 B.n682 B.n73 10.6151
R1078 B.n678 B.n73 10.6151
R1079 B.n678 B.n677 10.6151
R1080 B.n677 B.n676 10.6151
R1081 B.n676 B.n75 10.6151
R1082 B.n672 B.n75 10.6151
R1083 B.n672 B.n671 10.6151
R1084 B.n671 B.n670 10.6151
R1085 B.n670 B.n77 10.6151
R1086 B.n666 B.n77 10.6151
R1087 B.n666 B.n665 10.6151
R1088 B.n665 B.n664 10.6151
R1089 B.n664 B.n79 10.6151
R1090 B.n660 B.n79 10.6151
R1091 B.n660 B.n659 10.6151
R1092 B.n659 B.n658 10.6151
R1093 B.n658 B.n81 10.6151
R1094 B.n654 B.n81 10.6151
R1095 B.n654 B.n653 10.6151
R1096 B.n653 B.n652 10.6151
R1097 B.n652 B.n83 10.6151
R1098 B.n648 B.n83 10.6151
R1099 B.n648 B.n647 10.6151
R1100 B.n647 B.n646 10.6151
R1101 B.n646 B.n85 10.6151
R1102 B.n642 B.n85 10.6151
R1103 B.n642 B.n641 10.6151
R1104 B.n641 B.n640 10.6151
R1105 B.n640 B.n87 10.6151
R1106 B.n636 B.n87 10.6151
R1107 B.n636 B.n635 10.6151
R1108 B.n635 B.n634 10.6151
R1109 B.n634 B.n89 10.6151
R1110 B.n630 B.n89 10.6151
R1111 B.n630 B.n629 10.6151
R1112 B.n629 B.n628 10.6151
R1113 B.n628 B.n91 10.6151
R1114 B.n624 B.n91 10.6151
R1115 B.n624 B.n623 10.6151
R1116 B.n623 B.n622 10.6151
R1117 B.n622 B.n93 10.6151
R1118 B.n618 B.n93 10.6151
R1119 B.n618 B.n617 10.6151
R1120 B.n617 B.n616 10.6151
R1121 B.n612 B.n95 10.6151
R1122 B.n612 B.n611 10.6151
R1123 B.n611 B.n610 10.6151
R1124 B.n610 B.n97 10.6151
R1125 B.n606 B.n97 10.6151
R1126 B.n606 B.n605 10.6151
R1127 B.n605 B.n604 10.6151
R1128 B.n604 B.n99 10.6151
R1129 B.n600 B.n99 10.6151
R1130 B.n600 B.n599 10.6151
R1131 B.n599 B.n598 10.6151
R1132 B.n598 B.n101 10.6151
R1133 B.n594 B.n101 10.6151
R1134 B.n594 B.n593 10.6151
R1135 B.n593 B.n592 10.6151
R1136 B.n592 B.n103 10.6151
R1137 B.n588 B.n103 10.6151
R1138 B.n588 B.n587 10.6151
R1139 B.n587 B.n586 10.6151
R1140 B.n586 B.n105 10.6151
R1141 B.n582 B.n105 10.6151
R1142 B.n582 B.n581 10.6151
R1143 B.n581 B.n580 10.6151
R1144 B.n580 B.n107 10.6151
R1145 B.n576 B.n107 10.6151
R1146 B.n576 B.n575 10.6151
R1147 B.n575 B.n574 10.6151
R1148 B.n574 B.n109 10.6151
R1149 B.n570 B.n109 10.6151
R1150 B.n570 B.n569 10.6151
R1151 B.n569 B.n568 10.6151
R1152 B.n568 B.n111 10.6151
R1153 B.n564 B.n111 10.6151
R1154 B.n564 B.n563 10.6151
R1155 B.n563 B.n562 10.6151
R1156 B.n562 B.n113 10.6151
R1157 B.n558 B.n113 10.6151
R1158 B.n558 B.n557 10.6151
R1159 B.n557 B.n556 10.6151
R1160 B.n556 B.n115 10.6151
R1161 B.n552 B.n115 10.6151
R1162 B.n552 B.n551 10.6151
R1163 B.n551 B.n550 10.6151
R1164 B.n550 B.n117 10.6151
R1165 B.n546 B.n117 10.6151
R1166 B.n546 B.n545 10.6151
R1167 B.n545 B.n544 10.6151
R1168 B.n544 B.n119 10.6151
R1169 B.n540 B.n119 10.6151
R1170 B.n540 B.n539 10.6151
R1171 B.n539 B.n538 10.6151
R1172 B.n538 B.n121 10.6151
R1173 B.n534 B.n121 10.6151
R1174 B.n534 B.n533 10.6151
R1175 B.n533 B.n532 10.6151
R1176 B.n532 B.n123 10.6151
R1177 B.n528 B.n123 10.6151
R1178 B.n528 B.n527 10.6151
R1179 B.n527 B.n526 10.6151
R1180 B.n526 B.n125 10.6151
R1181 B.n522 B.n125 10.6151
R1182 B.n522 B.n521 10.6151
R1183 B.n521 B.n520 10.6151
R1184 B.n520 B.n127 10.6151
R1185 B.n516 B.n127 10.6151
R1186 B.n516 B.n515 10.6151
R1187 B.n515 B.n514 10.6151
R1188 B.n514 B.n129 10.6151
R1189 B.n510 B.n129 10.6151
R1190 B.n510 B.n509 10.6151
R1191 B.n509 B.n508 10.6151
R1192 B.n508 B.n131 10.6151
R1193 B.n504 B.n131 10.6151
R1194 B.n504 B.n503 10.6151
R1195 B.n503 B.n502 10.6151
R1196 B.n502 B.n133 10.6151
R1197 B.n498 B.n133 10.6151
R1198 B.n498 B.n497 10.6151
R1199 B.n497 B.n496 10.6151
R1200 B.n496 B.n135 10.6151
R1201 B.n492 B.n135 10.6151
R1202 B.n225 B.n1 10.6151
R1203 B.n228 B.n225 10.6151
R1204 B.n229 B.n228 10.6151
R1205 B.n230 B.n229 10.6151
R1206 B.n230 B.n223 10.6151
R1207 B.n234 B.n223 10.6151
R1208 B.n235 B.n234 10.6151
R1209 B.n236 B.n235 10.6151
R1210 B.n236 B.n221 10.6151
R1211 B.n240 B.n221 10.6151
R1212 B.n241 B.n240 10.6151
R1213 B.n242 B.n241 10.6151
R1214 B.n242 B.n219 10.6151
R1215 B.n246 B.n219 10.6151
R1216 B.n247 B.n246 10.6151
R1217 B.n248 B.n247 10.6151
R1218 B.n248 B.n217 10.6151
R1219 B.n252 B.n217 10.6151
R1220 B.n253 B.n252 10.6151
R1221 B.n254 B.n253 10.6151
R1222 B.n254 B.n215 10.6151
R1223 B.n258 B.n215 10.6151
R1224 B.n259 B.n258 10.6151
R1225 B.n260 B.n259 10.6151
R1226 B.n260 B.n213 10.6151
R1227 B.n264 B.n213 10.6151
R1228 B.n265 B.n264 10.6151
R1229 B.n266 B.n265 10.6151
R1230 B.n266 B.n211 10.6151
R1231 B.n270 B.n211 10.6151
R1232 B.n271 B.n270 10.6151
R1233 B.n272 B.n271 10.6151
R1234 B.n272 B.n209 10.6151
R1235 B.n276 B.n209 10.6151
R1236 B.n277 B.n276 10.6151
R1237 B.n278 B.n277 10.6151
R1238 B.n278 B.n207 10.6151
R1239 B.n282 B.n207 10.6151
R1240 B.n283 B.n282 10.6151
R1241 B.n284 B.n205 10.6151
R1242 B.n288 B.n205 10.6151
R1243 B.n289 B.n288 10.6151
R1244 B.n290 B.n289 10.6151
R1245 B.n290 B.n203 10.6151
R1246 B.n294 B.n203 10.6151
R1247 B.n295 B.n294 10.6151
R1248 B.n296 B.n295 10.6151
R1249 B.n296 B.n201 10.6151
R1250 B.n300 B.n201 10.6151
R1251 B.n301 B.n300 10.6151
R1252 B.n302 B.n301 10.6151
R1253 B.n302 B.n199 10.6151
R1254 B.n306 B.n199 10.6151
R1255 B.n307 B.n306 10.6151
R1256 B.n308 B.n307 10.6151
R1257 B.n308 B.n197 10.6151
R1258 B.n312 B.n197 10.6151
R1259 B.n313 B.n312 10.6151
R1260 B.n314 B.n313 10.6151
R1261 B.n314 B.n195 10.6151
R1262 B.n318 B.n195 10.6151
R1263 B.n319 B.n318 10.6151
R1264 B.n320 B.n319 10.6151
R1265 B.n320 B.n193 10.6151
R1266 B.n324 B.n193 10.6151
R1267 B.n325 B.n324 10.6151
R1268 B.n326 B.n325 10.6151
R1269 B.n326 B.n191 10.6151
R1270 B.n330 B.n191 10.6151
R1271 B.n331 B.n330 10.6151
R1272 B.n332 B.n331 10.6151
R1273 B.n332 B.n189 10.6151
R1274 B.n336 B.n189 10.6151
R1275 B.n337 B.n336 10.6151
R1276 B.n338 B.n337 10.6151
R1277 B.n338 B.n187 10.6151
R1278 B.n342 B.n187 10.6151
R1279 B.n343 B.n342 10.6151
R1280 B.n344 B.n343 10.6151
R1281 B.n344 B.n185 10.6151
R1282 B.n348 B.n185 10.6151
R1283 B.n349 B.n348 10.6151
R1284 B.n350 B.n349 10.6151
R1285 B.n350 B.n183 10.6151
R1286 B.n354 B.n183 10.6151
R1287 B.n355 B.n354 10.6151
R1288 B.n356 B.n355 10.6151
R1289 B.n356 B.n181 10.6151
R1290 B.n360 B.n181 10.6151
R1291 B.n361 B.n360 10.6151
R1292 B.n362 B.n361 10.6151
R1293 B.n362 B.n179 10.6151
R1294 B.n366 B.n179 10.6151
R1295 B.n367 B.n366 10.6151
R1296 B.n368 B.n367 10.6151
R1297 B.n368 B.n177 10.6151
R1298 B.n372 B.n177 10.6151
R1299 B.n373 B.n372 10.6151
R1300 B.n374 B.n373 10.6151
R1301 B.n374 B.n175 10.6151
R1302 B.n378 B.n175 10.6151
R1303 B.n381 B.n380 10.6151
R1304 B.n381 B.n171 10.6151
R1305 B.n385 B.n171 10.6151
R1306 B.n386 B.n385 10.6151
R1307 B.n387 B.n386 10.6151
R1308 B.n387 B.n169 10.6151
R1309 B.n391 B.n169 10.6151
R1310 B.n392 B.n391 10.6151
R1311 B.n396 B.n392 10.6151
R1312 B.n400 B.n167 10.6151
R1313 B.n401 B.n400 10.6151
R1314 B.n402 B.n401 10.6151
R1315 B.n402 B.n165 10.6151
R1316 B.n406 B.n165 10.6151
R1317 B.n407 B.n406 10.6151
R1318 B.n408 B.n407 10.6151
R1319 B.n408 B.n163 10.6151
R1320 B.n412 B.n163 10.6151
R1321 B.n413 B.n412 10.6151
R1322 B.n414 B.n413 10.6151
R1323 B.n414 B.n161 10.6151
R1324 B.n418 B.n161 10.6151
R1325 B.n419 B.n418 10.6151
R1326 B.n420 B.n419 10.6151
R1327 B.n420 B.n159 10.6151
R1328 B.n424 B.n159 10.6151
R1329 B.n425 B.n424 10.6151
R1330 B.n426 B.n425 10.6151
R1331 B.n426 B.n157 10.6151
R1332 B.n430 B.n157 10.6151
R1333 B.n431 B.n430 10.6151
R1334 B.n432 B.n431 10.6151
R1335 B.n432 B.n155 10.6151
R1336 B.n436 B.n155 10.6151
R1337 B.n437 B.n436 10.6151
R1338 B.n438 B.n437 10.6151
R1339 B.n438 B.n153 10.6151
R1340 B.n442 B.n153 10.6151
R1341 B.n443 B.n442 10.6151
R1342 B.n444 B.n443 10.6151
R1343 B.n444 B.n151 10.6151
R1344 B.n448 B.n151 10.6151
R1345 B.n449 B.n448 10.6151
R1346 B.n450 B.n449 10.6151
R1347 B.n450 B.n149 10.6151
R1348 B.n454 B.n149 10.6151
R1349 B.n455 B.n454 10.6151
R1350 B.n456 B.n455 10.6151
R1351 B.n456 B.n147 10.6151
R1352 B.n460 B.n147 10.6151
R1353 B.n461 B.n460 10.6151
R1354 B.n462 B.n461 10.6151
R1355 B.n462 B.n145 10.6151
R1356 B.n466 B.n145 10.6151
R1357 B.n467 B.n466 10.6151
R1358 B.n468 B.n467 10.6151
R1359 B.n468 B.n143 10.6151
R1360 B.n472 B.n143 10.6151
R1361 B.n473 B.n472 10.6151
R1362 B.n474 B.n473 10.6151
R1363 B.n474 B.n141 10.6151
R1364 B.n478 B.n141 10.6151
R1365 B.n479 B.n478 10.6151
R1366 B.n480 B.n479 10.6151
R1367 B.n480 B.n139 10.6151
R1368 B.n484 B.n139 10.6151
R1369 B.n485 B.n484 10.6151
R1370 B.n486 B.n485 10.6151
R1371 B.n486 B.n137 10.6151
R1372 B.n490 B.n137 10.6151
R1373 B.n491 B.n490 10.6151
R1374 B.n726 B.n725 9.36635
R1375 B.n708 B.n64 9.36635
R1376 B.n379 B.n378 9.36635
R1377 B.n395 B.n167 9.36635
R1378 B.n881 B.n0 8.11757
R1379 B.n881 B.n1 8.11757
R1380 B.n725 B.n724 1.24928
R1381 B.n64 B.n60 1.24928
R1382 B.n380 B.n379 1.24928
R1383 B.n396 B.n395 1.24928
R1384 VN.n1 VN.t0 175.044
R1385 VN.n0 VN.t1 175.044
R1386 VN.n0 VN.t3 173.917
R1387 VN.n1 VN.t2 173.917
R1388 VN VN.n1 56.8214
R1389 VN VN.n0 2.44645
R1390 VDD2.n2 VDD2.n0 118.688
R1391 VDD2.n2 VDD2.n1 68.8255
R1392 VDD2.n1 VDD2.t1 1.68034
R1393 VDD2.n1 VDD2.t3 1.68034
R1394 VDD2.n0 VDD2.t2 1.68034
R1395 VDD2.n0 VDD2.t0 1.68034
R1396 VDD2 VDD2.n2 0.0586897
C0 VDD1 w_n3166_n4838# 1.78531f
C1 VDD2 VP 0.440603f
C2 VP w_n3166_n4838# 6.04258f
C3 VDD2 w_n3166_n4838# 1.85755f
C4 B VTAIL 7.75339f
C5 VTAIL VN 7.45106f
C6 B VN 1.33364f
C7 VDD1 VTAIL 7.18217f
C8 B VDD1 1.58877f
C9 VDD1 VN 0.149506f
C10 VTAIL VP 7.46516f
C11 B VP 2.0155f
C12 VP VN 8.07749f
C13 VDD2 VTAIL 7.24128f
C14 B VDD2 1.65302f
C15 VDD2 VN 7.77792f
C16 VTAIL w_n3166_n4838# 5.61475f
C17 B w_n3166_n4838# 12.2037f
C18 VDD1 VP 8.068089f
C19 VN w_n3166_n4838# 5.63373f
C20 VDD2 VDD1 1.19746f
C21 VDD2 VSUBS 1.243257f
C22 VDD1 VSUBS 7.081229f
C23 VTAIL VSUBS 1.641981f
C24 VN VSUBS 6.10355f
C25 VP VSUBS 2.94583f
C26 B VSUBS 5.525983f
C27 w_n3166_n4838# VSUBS 0.187111p
C28 VDD2.t2 VSUBS 0.405786f
C29 VDD2.t0 VSUBS 0.405786f
C30 VDD2.n0 VSUBS 4.4554f
C31 VDD2.t1 VSUBS 0.405786f
C32 VDD2.t3 VSUBS 0.405786f
C33 VDD2.n1 VSUBS 3.40175f
C34 VDD2.n2 VSUBS 5.2442f
C35 VN.t3 VSUBS 4.81239f
C36 VN.t1 VSUBS 4.82314f
C37 VN.n0 VSUBS 2.98073f
C38 VN.t2 VSUBS 4.81239f
C39 VN.t0 VSUBS 4.82314f
C40 VN.n1 VSUBS 4.77541f
C41 B.n0 VSUBS 0.00539f
C42 B.n1 VSUBS 0.00539f
C43 B.n2 VSUBS 0.007971f
C44 B.n3 VSUBS 0.006108f
C45 B.n4 VSUBS 0.006108f
C46 B.n5 VSUBS 0.006108f
C47 B.n6 VSUBS 0.006108f
C48 B.n7 VSUBS 0.006108f
C49 B.n8 VSUBS 0.006108f
C50 B.n9 VSUBS 0.006108f
C51 B.n10 VSUBS 0.006108f
C52 B.n11 VSUBS 0.006108f
C53 B.n12 VSUBS 0.006108f
C54 B.n13 VSUBS 0.006108f
C55 B.n14 VSUBS 0.006108f
C56 B.n15 VSUBS 0.006108f
C57 B.n16 VSUBS 0.006108f
C58 B.n17 VSUBS 0.006108f
C59 B.n18 VSUBS 0.006108f
C60 B.n19 VSUBS 0.006108f
C61 B.n20 VSUBS 0.006108f
C62 B.n21 VSUBS 0.006108f
C63 B.n22 VSUBS 0.014295f
C64 B.n23 VSUBS 0.006108f
C65 B.n24 VSUBS 0.006108f
C66 B.n25 VSUBS 0.006108f
C67 B.n26 VSUBS 0.006108f
C68 B.n27 VSUBS 0.006108f
C69 B.n28 VSUBS 0.006108f
C70 B.n29 VSUBS 0.006108f
C71 B.n30 VSUBS 0.006108f
C72 B.n31 VSUBS 0.006108f
C73 B.n32 VSUBS 0.006108f
C74 B.n33 VSUBS 0.006108f
C75 B.n34 VSUBS 0.006108f
C76 B.n35 VSUBS 0.006108f
C77 B.n36 VSUBS 0.006108f
C78 B.n37 VSUBS 0.006108f
C79 B.n38 VSUBS 0.006108f
C80 B.n39 VSUBS 0.006108f
C81 B.n40 VSUBS 0.006108f
C82 B.n41 VSUBS 0.006108f
C83 B.n42 VSUBS 0.006108f
C84 B.n43 VSUBS 0.006108f
C85 B.n44 VSUBS 0.006108f
C86 B.n45 VSUBS 0.006108f
C87 B.n46 VSUBS 0.006108f
C88 B.n47 VSUBS 0.006108f
C89 B.n48 VSUBS 0.006108f
C90 B.n49 VSUBS 0.006108f
C91 B.n50 VSUBS 0.006108f
C92 B.n51 VSUBS 0.006108f
C93 B.n52 VSUBS 0.006108f
C94 B.n53 VSUBS 0.006108f
C95 B.t7 VSUBS 0.572847f
C96 B.t8 VSUBS 0.594902f
C97 B.t6 VSUBS 2.52727f
C98 B.n54 VSUBS 0.3623f
C99 B.n55 VSUBS 0.065588f
C100 B.n56 VSUBS 0.006108f
C101 B.n57 VSUBS 0.006108f
C102 B.n58 VSUBS 0.006108f
C103 B.n59 VSUBS 0.006108f
C104 B.n60 VSUBS 0.003414f
C105 B.n61 VSUBS 0.006108f
C106 B.t10 VSUBS 0.572824f
C107 B.t11 VSUBS 0.594885f
C108 B.t9 VSUBS 2.52727f
C109 B.n62 VSUBS 0.362317f
C110 B.n63 VSUBS 0.065611f
C111 B.n64 VSUBS 0.014152f
C112 B.n65 VSUBS 0.006108f
C113 B.n66 VSUBS 0.006108f
C114 B.n67 VSUBS 0.006108f
C115 B.n68 VSUBS 0.006108f
C116 B.n69 VSUBS 0.006108f
C117 B.n70 VSUBS 0.006108f
C118 B.n71 VSUBS 0.006108f
C119 B.n72 VSUBS 0.006108f
C120 B.n73 VSUBS 0.006108f
C121 B.n74 VSUBS 0.006108f
C122 B.n75 VSUBS 0.006108f
C123 B.n76 VSUBS 0.006108f
C124 B.n77 VSUBS 0.006108f
C125 B.n78 VSUBS 0.006108f
C126 B.n79 VSUBS 0.006108f
C127 B.n80 VSUBS 0.006108f
C128 B.n81 VSUBS 0.006108f
C129 B.n82 VSUBS 0.006108f
C130 B.n83 VSUBS 0.006108f
C131 B.n84 VSUBS 0.006108f
C132 B.n85 VSUBS 0.006108f
C133 B.n86 VSUBS 0.006108f
C134 B.n87 VSUBS 0.006108f
C135 B.n88 VSUBS 0.006108f
C136 B.n89 VSUBS 0.006108f
C137 B.n90 VSUBS 0.006108f
C138 B.n91 VSUBS 0.006108f
C139 B.n92 VSUBS 0.006108f
C140 B.n93 VSUBS 0.006108f
C141 B.n94 VSUBS 0.006108f
C142 B.n95 VSUBS 0.013732f
C143 B.n96 VSUBS 0.006108f
C144 B.n97 VSUBS 0.006108f
C145 B.n98 VSUBS 0.006108f
C146 B.n99 VSUBS 0.006108f
C147 B.n100 VSUBS 0.006108f
C148 B.n101 VSUBS 0.006108f
C149 B.n102 VSUBS 0.006108f
C150 B.n103 VSUBS 0.006108f
C151 B.n104 VSUBS 0.006108f
C152 B.n105 VSUBS 0.006108f
C153 B.n106 VSUBS 0.006108f
C154 B.n107 VSUBS 0.006108f
C155 B.n108 VSUBS 0.006108f
C156 B.n109 VSUBS 0.006108f
C157 B.n110 VSUBS 0.006108f
C158 B.n111 VSUBS 0.006108f
C159 B.n112 VSUBS 0.006108f
C160 B.n113 VSUBS 0.006108f
C161 B.n114 VSUBS 0.006108f
C162 B.n115 VSUBS 0.006108f
C163 B.n116 VSUBS 0.006108f
C164 B.n117 VSUBS 0.006108f
C165 B.n118 VSUBS 0.006108f
C166 B.n119 VSUBS 0.006108f
C167 B.n120 VSUBS 0.006108f
C168 B.n121 VSUBS 0.006108f
C169 B.n122 VSUBS 0.006108f
C170 B.n123 VSUBS 0.006108f
C171 B.n124 VSUBS 0.006108f
C172 B.n125 VSUBS 0.006108f
C173 B.n126 VSUBS 0.006108f
C174 B.n127 VSUBS 0.006108f
C175 B.n128 VSUBS 0.006108f
C176 B.n129 VSUBS 0.006108f
C177 B.n130 VSUBS 0.006108f
C178 B.n131 VSUBS 0.006108f
C179 B.n132 VSUBS 0.006108f
C180 B.n133 VSUBS 0.006108f
C181 B.n134 VSUBS 0.006108f
C182 B.n135 VSUBS 0.006108f
C183 B.n136 VSUBS 0.014295f
C184 B.n137 VSUBS 0.006108f
C185 B.n138 VSUBS 0.006108f
C186 B.n139 VSUBS 0.006108f
C187 B.n140 VSUBS 0.006108f
C188 B.n141 VSUBS 0.006108f
C189 B.n142 VSUBS 0.006108f
C190 B.n143 VSUBS 0.006108f
C191 B.n144 VSUBS 0.006108f
C192 B.n145 VSUBS 0.006108f
C193 B.n146 VSUBS 0.006108f
C194 B.n147 VSUBS 0.006108f
C195 B.n148 VSUBS 0.006108f
C196 B.n149 VSUBS 0.006108f
C197 B.n150 VSUBS 0.006108f
C198 B.n151 VSUBS 0.006108f
C199 B.n152 VSUBS 0.006108f
C200 B.n153 VSUBS 0.006108f
C201 B.n154 VSUBS 0.006108f
C202 B.n155 VSUBS 0.006108f
C203 B.n156 VSUBS 0.006108f
C204 B.n157 VSUBS 0.006108f
C205 B.n158 VSUBS 0.006108f
C206 B.n159 VSUBS 0.006108f
C207 B.n160 VSUBS 0.006108f
C208 B.n161 VSUBS 0.006108f
C209 B.n162 VSUBS 0.006108f
C210 B.n163 VSUBS 0.006108f
C211 B.n164 VSUBS 0.006108f
C212 B.n165 VSUBS 0.006108f
C213 B.n166 VSUBS 0.006108f
C214 B.n167 VSUBS 0.005749f
C215 B.n168 VSUBS 0.006108f
C216 B.n169 VSUBS 0.006108f
C217 B.n170 VSUBS 0.006108f
C218 B.n171 VSUBS 0.006108f
C219 B.n172 VSUBS 0.006108f
C220 B.t5 VSUBS 0.572847f
C221 B.t4 VSUBS 0.594902f
C222 B.t3 VSUBS 2.52727f
C223 B.n173 VSUBS 0.3623f
C224 B.n174 VSUBS 0.065588f
C225 B.n175 VSUBS 0.006108f
C226 B.n176 VSUBS 0.006108f
C227 B.n177 VSUBS 0.006108f
C228 B.n178 VSUBS 0.006108f
C229 B.n179 VSUBS 0.006108f
C230 B.n180 VSUBS 0.006108f
C231 B.n181 VSUBS 0.006108f
C232 B.n182 VSUBS 0.006108f
C233 B.n183 VSUBS 0.006108f
C234 B.n184 VSUBS 0.006108f
C235 B.n185 VSUBS 0.006108f
C236 B.n186 VSUBS 0.006108f
C237 B.n187 VSUBS 0.006108f
C238 B.n188 VSUBS 0.006108f
C239 B.n189 VSUBS 0.006108f
C240 B.n190 VSUBS 0.006108f
C241 B.n191 VSUBS 0.006108f
C242 B.n192 VSUBS 0.006108f
C243 B.n193 VSUBS 0.006108f
C244 B.n194 VSUBS 0.006108f
C245 B.n195 VSUBS 0.006108f
C246 B.n196 VSUBS 0.006108f
C247 B.n197 VSUBS 0.006108f
C248 B.n198 VSUBS 0.006108f
C249 B.n199 VSUBS 0.006108f
C250 B.n200 VSUBS 0.006108f
C251 B.n201 VSUBS 0.006108f
C252 B.n202 VSUBS 0.006108f
C253 B.n203 VSUBS 0.006108f
C254 B.n204 VSUBS 0.006108f
C255 B.n205 VSUBS 0.006108f
C256 B.n206 VSUBS 0.013732f
C257 B.n207 VSUBS 0.006108f
C258 B.n208 VSUBS 0.006108f
C259 B.n209 VSUBS 0.006108f
C260 B.n210 VSUBS 0.006108f
C261 B.n211 VSUBS 0.006108f
C262 B.n212 VSUBS 0.006108f
C263 B.n213 VSUBS 0.006108f
C264 B.n214 VSUBS 0.006108f
C265 B.n215 VSUBS 0.006108f
C266 B.n216 VSUBS 0.006108f
C267 B.n217 VSUBS 0.006108f
C268 B.n218 VSUBS 0.006108f
C269 B.n219 VSUBS 0.006108f
C270 B.n220 VSUBS 0.006108f
C271 B.n221 VSUBS 0.006108f
C272 B.n222 VSUBS 0.006108f
C273 B.n223 VSUBS 0.006108f
C274 B.n224 VSUBS 0.006108f
C275 B.n225 VSUBS 0.006108f
C276 B.n226 VSUBS 0.006108f
C277 B.n227 VSUBS 0.006108f
C278 B.n228 VSUBS 0.006108f
C279 B.n229 VSUBS 0.006108f
C280 B.n230 VSUBS 0.006108f
C281 B.n231 VSUBS 0.006108f
C282 B.n232 VSUBS 0.006108f
C283 B.n233 VSUBS 0.006108f
C284 B.n234 VSUBS 0.006108f
C285 B.n235 VSUBS 0.006108f
C286 B.n236 VSUBS 0.006108f
C287 B.n237 VSUBS 0.006108f
C288 B.n238 VSUBS 0.006108f
C289 B.n239 VSUBS 0.006108f
C290 B.n240 VSUBS 0.006108f
C291 B.n241 VSUBS 0.006108f
C292 B.n242 VSUBS 0.006108f
C293 B.n243 VSUBS 0.006108f
C294 B.n244 VSUBS 0.006108f
C295 B.n245 VSUBS 0.006108f
C296 B.n246 VSUBS 0.006108f
C297 B.n247 VSUBS 0.006108f
C298 B.n248 VSUBS 0.006108f
C299 B.n249 VSUBS 0.006108f
C300 B.n250 VSUBS 0.006108f
C301 B.n251 VSUBS 0.006108f
C302 B.n252 VSUBS 0.006108f
C303 B.n253 VSUBS 0.006108f
C304 B.n254 VSUBS 0.006108f
C305 B.n255 VSUBS 0.006108f
C306 B.n256 VSUBS 0.006108f
C307 B.n257 VSUBS 0.006108f
C308 B.n258 VSUBS 0.006108f
C309 B.n259 VSUBS 0.006108f
C310 B.n260 VSUBS 0.006108f
C311 B.n261 VSUBS 0.006108f
C312 B.n262 VSUBS 0.006108f
C313 B.n263 VSUBS 0.006108f
C314 B.n264 VSUBS 0.006108f
C315 B.n265 VSUBS 0.006108f
C316 B.n266 VSUBS 0.006108f
C317 B.n267 VSUBS 0.006108f
C318 B.n268 VSUBS 0.006108f
C319 B.n269 VSUBS 0.006108f
C320 B.n270 VSUBS 0.006108f
C321 B.n271 VSUBS 0.006108f
C322 B.n272 VSUBS 0.006108f
C323 B.n273 VSUBS 0.006108f
C324 B.n274 VSUBS 0.006108f
C325 B.n275 VSUBS 0.006108f
C326 B.n276 VSUBS 0.006108f
C327 B.n277 VSUBS 0.006108f
C328 B.n278 VSUBS 0.006108f
C329 B.n279 VSUBS 0.006108f
C330 B.n280 VSUBS 0.006108f
C331 B.n281 VSUBS 0.006108f
C332 B.n282 VSUBS 0.006108f
C333 B.n283 VSUBS 0.013732f
C334 B.n284 VSUBS 0.014295f
C335 B.n285 VSUBS 0.014295f
C336 B.n286 VSUBS 0.006108f
C337 B.n287 VSUBS 0.006108f
C338 B.n288 VSUBS 0.006108f
C339 B.n289 VSUBS 0.006108f
C340 B.n290 VSUBS 0.006108f
C341 B.n291 VSUBS 0.006108f
C342 B.n292 VSUBS 0.006108f
C343 B.n293 VSUBS 0.006108f
C344 B.n294 VSUBS 0.006108f
C345 B.n295 VSUBS 0.006108f
C346 B.n296 VSUBS 0.006108f
C347 B.n297 VSUBS 0.006108f
C348 B.n298 VSUBS 0.006108f
C349 B.n299 VSUBS 0.006108f
C350 B.n300 VSUBS 0.006108f
C351 B.n301 VSUBS 0.006108f
C352 B.n302 VSUBS 0.006108f
C353 B.n303 VSUBS 0.006108f
C354 B.n304 VSUBS 0.006108f
C355 B.n305 VSUBS 0.006108f
C356 B.n306 VSUBS 0.006108f
C357 B.n307 VSUBS 0.006108f
C358 B.n308 VSUBS 0.006108f
C359 B.n309 VSUBS 0.006108f
C360 B.n310 VSUBS 0.006108f
C361 B.n311 VSUBS 0.006108f
C362 B.n312 VSUBS 0.006108f
C363 B.n313 VSUBS 0.006108f
C364 B.n314 VSUBS 0.006108f
C365 B.n315 VSUBS 0.006108f
C366 B.n316 VSUBS 0.006108f
C367 B.n317 VSUBS 0.006108f
C368 B.n318 VSUBS 0.006108f
C369 B.n319 VSUBS 0.006108f
C370 B.n320 VSUBS 0.006108f
C371 B.n321 VSUBS 0.006108f
C372 B.n322 VSUBS 0.006108f
C373 B.n323 VSUBS 0.006108f
C374 B.n324 VSUBS 0.006108f
C375 B.n325 VSUBS 0.006108f
C376 B.n326 VSUBS 0.006108f
C377 B.n327 VSUBS 0.006108f
C378 B.n328 VSUBS 0.006108f
C379 B.n329 VSUBS 0.006108f
C380 B.n330 VSUBS 0.006108f
C381 B.n331 VSUBS 0.006108f
C382 B.n332 VSUBS 0.006108f
C383 B.n333 VSUBS 0.006108f
C384 B.n334 VSUBS 0.006108f
C385 B.n335 VSUBS 0.006108f
C386 B.n336 VSUBS 0.006108f
C387 B.n337 VSUBS 0.006108f
C388 B.n338 VSUBS 0.006108f
C389 B.n339 VSUBS 0.006108f
C390 B.n340 VSUBS 0.006108f
C391 B.n341 VSUBS 0.006108f
C392 B.n342 VSUBS 0.006108f
C393 B.n343 VSUBS 0.006108f
C394 B.n344 VSUBS 0.006108f
C395 B.n345 VSUBS 0.006108f
C396 B.n346 VSUBS 0.006108f
C397 B.n347 VSUBS 0.006108f
C398 B.n348 VSUBS 0.006108f
C399 B.n349 VSUBS 0.006108f
C400 B.n350 VSUBS 0.006108f
C401 B.n351 VSUBS 0.006108f
C402 B.n352 VSUBS 0.006108f
C403 B.n353 VSUBS 0.006108f
C404 B.n354 VSUBS 0.006108f
C405 B.n355 VSUBS 0.006108f
C406 B.n356 VSUBS 0.006108f
C407 B.n357 VSUBS 0.006108f
C408 B.n358 VSUBS 0.006108f
C409 B.n359 VSUBS 0.006108f
C410 B.n360 VSUBS 0.006108f
C411 B.n361 VSUBS 0.006108f
C412 B.n362 VSUBS 0.006108f
C413 B.n363 VSUBS 0.006108f
C414 B.n364 VSUBS 0.006108f
C415 B.n365 VSUBS 0.006108f
C416 B.n366 VSUBS 0.006108f
C417 B.n367 VSUBS 0.006108f
C418 B.n368 VSUBS 0.006108f
C419 B.n369 VSUBS 0.006108f
C420 B.n370 VSUBS 0.006108f
C421 B.n371 VSUBS 0.006108f
C422 B.n372 VSUBS 0.006108f
C423 B.n373 VSUBS 0.006108f
C424 B.n374 VSUBS 0.006108f
C425 B.n375 VSUBS 0.006108f
C426 B.n376 VSUBS 0.006108f
C427 B.n377 VSUBS 0.006108f
C428 B.n378 VSUBS 0.005749f
C429 B.n379 VSUBS 0.014152f
C430 B.n380 VSUBS 0.003414f
C431 B.n381 VSUBS 0.006108f
C432 B.n382 VSUBS 0.006108f
C433 B.n383 VSUBS 0.006108f
C434 B.n384 VSUBS 0.006108f
C435 B.n385 VSUBS 0.006108f
C436 B.n386 VSUBS 0.006108f
C437 B.n387 VSUBS 0.006108f
C438 B.n388 VSUBS 0.006108f
C439 B.n389 VSUBS 0.006108f
C440 B.n390 VSUBS 0.006108f
C441 B.n391 VSUBS 0.006108f
C442 B.n392 VSUBS 0.006108f
C443 B.t2 VSUBS 0.572824f
C444 B.t1 VSUBS 0.594885f
C445 B.t0 VSUBS 2.52727f
C446 B.n393 VSUBS 0.362317f
C447 B.n394 VSUBS 0.065611f
C448 B.n395 VSUBS 0.014152f
C449 B.n396 VSUBS 0.003414f
C450 B.n397 VSUBS 0.006108f
C451 B.n398 VSUBS 0.006108f
C452 B.n399 VSUBS 0.006108f
C453 B.n400 VSUBS 0.006108f
C454 B.n401 VSUBS 0.006108f
C455 B.n402 VSUBS 0.006108f
C456 B.n403 VSUBS 0.006108f
C457 B.n404 VSUBS 0.006108f
C458 B.n405 VSUBS 0.006108f
C459 B.n406 VSUBS 0.006108f
C460 B.n407 VSUBS 0.006108f
C461 B.n408 VSUBS 0.006108f
C462 B.n409 VSUBS 0.006108f
C463 B.n410 VSUBS 0.006108f
C464 B.n411 VSUBS 0.006108f
C465 B.n412 VSUBS 0.006108f
C466 B.n413 VSUBS 0.006108f
C467 B.n414 VSUBS 0.006108f
C468 B.n415 VSUBS 0.006108f
C469 B.n416 VSUBS 0.006108f
C470 B.n417 VSUBS 0.006108f
C471 B.n418 VSUBS 0.006108f
C472 B.n419 VSUBS 0.006108f
C473 B.n420 VSUBS 0.006108f
C474 B.n421 VSUBS 0.006108f
C475 B.n422 VSUBS 0.006108f
C476 B.n423 VSUBS 0.006108f
C477 B.n424 VSUBS 0.006108f
C478 B.n425 VSUBS 0.006108f
C479 B.n426 VSUBS 0.006108f
C480 B.n427 VSUBS 0.006108f
C481 B.n428 VSUBS 0.006108f
C482 B.n429 VSUBS 0.006108f
C483 B.n430 VSUBS 0.006108f
C484 B.n431 VSUBS 0.006108f
C485 B.n432 VSUBS 0.006108f
C486 B.n433 VSUBS 0.006108f
C487 B.n434 VSUBS 0.006108f
C488 B.n435 VSUBS 0.006108f
C489 B.n436 VSUBS 0.006108f
C490 B.n437 VSUBS 0.006108f
C491 B.n438 VSUBS 0.006108f
C492 B.n439 VSUBS 0.006108f
C493 B.n440 VSUBS 0.006108f
C494 B.n441 VSUBS 0.006108f
C495 B.n442 VSUBS 0.006108f
C496 B.n443 VSUBS 0.006108f
C497 B.n444 VSUBS 0.006108f
C498 B.n445 VSUBS 0.006108f
C499 B.n446 VSUBS 0.006108f
C500 B.n447 VSUBS 0.006108f
C501 B.n448 VSUBS 0.006108f
C502 B.n449 VSUBS 0.006108f
C503 B.n450 VSUBS 0.006108f
C504 B.n451 VSUBS 0.006108f
C505 B.n452 VSUBS 0.006108f
C506 B.n453 VSUBS 0.006108f
C507 B.n454 VSUBS 0.006108f
C508 B.n455 VSUBS 0.006108f
C509 B.n456 VSUBS 0.006108f
C510 B.n457 VSUBS 0.006108f
C511 B.n458 VSUBS 0.006108f
C512 B.n459 VSUBS 0.006108f
C513 B.n460 VSUBS 0.006108f
C514 B.n461 VSUBS 0.006108f
C515 B.n462 VSUBS 0.006108f
C516 B.n463 VSUBS 0.006108f
C517 B.n464 VSUBS 0.006108f
C518 B.n465 VSUBS 0.006108f
C519 B.n466 VSUBS 0.006108f
C520 B.n467 VSUBS 0.006108f
C521 B.n468 VSUBS 0.006108f
C522 B.n469 VSUBS 0.006108f
C523 B.n470 VSUBS 0.006108f
C524 B.n471 VSUBS 0.006108f
C525 B.n472 VSUBS 0.006108f
C526 B.n473 VSUBS 0.006108f
C527 B.n474 VSUBS 0.006108f
C528 B.n475 VSUBS 0.006108f
C529 B.n476 VSUBS 0.006108f
C530 B.n477 VSUBS 0.006108f
C531 B.n478 VSUBS 0.006108f
C532 B.n479 VSUBS 0.006108f
C533 B.n480 VSUBS 0.006108f
C534 B.n481 VSUBS 0.006108f
C535 B.n482 VSUBS 0.006108f
C536 B.n483 VSUBS 0.006108f
C537 B.n484 VSUBS 0.006108f
C538 B.n485 VSUBS 0.006108f
C539 B.n486 VSUBS 0.006108f
C540 B.n487 VSUBS 0.006108f
C541 B.n488 VSUBS 0.006108f
C542 B.n489 VSUBS 0.006108f
C543 B.n490 VSUBS 0.006108f
C544 B.n491 VSUBS 0.013551f
C545 B.n492 VSUBS 0.014476f
C546 B.n493 VSUBS 0.013732f
C547 B.n494 VSUBS 0.006108f
C548 B.n495 VSUBS 0.006108f
C549 B.n496 VSUBS 0.006108f
C550 B.n497 VSUBS 0.006108f
C551 B.n498 VSUBS 0.006108f
C552 B.n499 VSUBS 0.006108f
C553 B.n500 VSUBS 0.006108f
C554 B.n501 VSUBS 0.006108f
C555 B.n502 VSUBS 0.006108f
C556 B.n503 VSUBS 0.006108f
C557 B.n504 VSUBS 0.006108f
C558 B.n505 VSUBS 0.006108f
C559 B.n506 VSUBS 0.006108f
C560 B.n507 VSUBS 0.006108f
C561 B.n508 VSUBS 0.006108f
C562 B.n509 VSUBS 0.006108f
C563 B.n510 VSUBS 0.006108f
C564 B.n511 VSUBS 0.006108f
C565 B.n512 VSUBS 0.006108f
C566 B.n513 VSUBS 0.006108f
C567 B.n514 VSUBS 0.006108f
C568 B.n515 VSUBS 0.006108f
C569 B.n516 VSUBS 0.006108f
C570 B.n517 VSUBS 0.006108f
C571 B.n518 VSUBS 0.006108f
C572 B.n519 VSUBS 0.006108f
C573 B.n520 VSUBS 0.006108f
C574 B.n521 VSUBS 0.006108f
C575 B.n522 VSUBS 0.006108f
C576 B.n523 VSUBS 0.006108f
C577 B.n524 VSUBS 0.006108f
C578 B.n525 VSUBS 0.006108f
C579 B.n526 VSUBS 0.006108f
C580 B.n527 VSUBS 0.006108f
C581 B.n528 VSUBS 0.006108f
C582 B.n529 VSUBS 0.006108f
C583 B.n530 VSUBS 0.006108f
C584 B.n531 VSUBS 0.006108f
C585 B.n532 VSUBS 0.006108f
C586 B.n533 VSUBS 0.006108f
C587 B.n534 VSUBS 0.006108f
C588 B.n535 VSUBS 0.006108f
C589 B.n536 VSUBS 0.006108f
C590 B.n537 VSUBS 0.006108f
C591 B.n538 VSUBS 0.006108f
C592 B.n539 VSUBS 0.006108f
C593 B.n540 VSUBS 0.006108f
C594 B.n541 VSUBS 0.006108f
C595 B.n542 VSUBS 0.006108f
C596 B.n543 VSUBS 0.006108f
C597 B.n544 VSUBS 0.006108f
C598 B.n545 VSUBS 0.006108f
C599 B.n546 VSUBS 0.006108f
C600 B.n547 VSUBS 0.006108f
C601 B.n548 VSUBS 0.006108f
C602 B.n549 VSUBS 0.006108f
C603 B.n550 VSUBS 0.006108f
C604 B.n551 VSUBS 0.006108f
C605 B.n552 VSUBS 0.006108f
C606 B.n553 VSUBS 0.006108f
C607 B.n554 VSUBS 0.006108f
C608 B.n555 VSUBS 0.006108f
C609 B.n556 VSUBS 0.006108f
C610 B.n557 VSUBS 0.006108f
C611 B.n558 VSUBS 0.006108f
C612 B.n559 VSUBS 0.006108f
C613 B.n560 VSUBS 0.006108f
C614 B.n561 VSUBS 0.006108f
C615 B.n562 VSUBS 0.006108f
C616 B.n563 VSUBS 0.006108f
C617 B.n564 VSUBS 0.006108f
C618 B.n565 VSUBS 0.006108f
C619 B.n566 VSUBS 0.006108f
C620 B.n567 VSUBS 0.006108f
C621 B.n568 VSUBS 0.006108f
C622 B.n569 VSUBS 0.006108f
C623 B.n570 VSUBS 0.006108f
C624 B.n571 VSUBS 0.006108f
C625 B.n572 VSUBS 0.006108f
C626 B.n573 VSUBS 0.006108f
C627 B.n574 VSUBS 0.006108f
C628 B.n575 VSUBS 0.006108f
C629 B.n576 VSUBS 0.006108f
C630 B.n577 VSUBS 0.006108f
C631 B.n578 VSUBS 0.006108f
C632 B.n579 VSUBS 0.006108f
C633 B.n580 VSUBS 0.006108f
C634 B.n581 VSUBS 0.006108f
C635 B.n582 VSUBS 0.006108f
C636 B.n583 VSUBS 0.006108f
C637 B.n584 VSUBS 0.006108f
C638 B.n585 VSUBS 0.006108f
C639 B.n586 VSUBS 0.006108f
C640 B.n587 VSUBS 0.006108f
C641 B.n588 VSUBS 0.006108f
C642 B.n589 VSUBS 0.006108f
C643 B.n590 VSUBS 0.006108f
C644 B.n591 VSUBS 0.006108f
C645 B.n592 VSUBS 0.006108f
C646 B.n593 VSUBS 0.006108f
C647 B.n594 VSUBS 0.006108f
C648 B.n595 VSUBS 0.006108f
C649 B.n596 VSUBS 0.006108f
C650 B.n597 VSUBS 0.006108f
C651 B.n598 VSUBS 0.006108f
C652 B.n599 VSUBS 0.006108f
C653 B.n600 VSUBS 0.006108f
C654 B.n601 VSUBS 0.006108f
C655 B.n602 VSUBS 0.006108f
C656 B.n603 VSUBS 0.006108f
C657 B.n604 VSUBS 0.006108f
C658 B.n605 VSUBS 0.006108f
C659 B.n606 VSUBS 0.006108f
C660 B.n607 VSUBS 0.006108f
C661 B.n608 VSUBS 0.006108f
C662 B.n609 VSUBS 0.006108f
C663 B.n610 VSUBS 0.006108f
C664 B.n611 VSUBS 0.006108f
C665 B.n612 VSUBS 0.006108f
C666 B.n613 VSUBS 0.006108f
C667 B.n614 VSUBS 0.013732f
C668 B.n615 VSUBS 0.014295f
C669 B.n616 VSUBS 0.014295f
C670 B.n617 VSUBS 0.006108f
C671 B.n618 VSUBS 0.006108f
C672 B.n619 VSUBS 0.006108f
C673 B.n620 VSUBS 0.006108f
C674 B.n621 VSUBS 0.006108f
C675 B.n622 VSUBS 0.006108f
C676 B.n623 VSUBS 0.006108f
C677 B.n624 VSUBS 0.006108f
C678 B.n625 VSUBS 0.006108f
C679 B.n626 VSUBS 0.006108f
C680 B.n627 VSUBS 0.006108f
C681 B.n628 VSUBS 0.006108f
C682 B.n629 VSUBS 0.006108f
C683 B.n630 VSUBS 0.006108f
C684 B.n631 VSUBS 0.006108f
C685 B.n632 VSUBS 0.006108f
C686 B.n633 VSUBS 0.006108f
C687 B.n634 VSUBS 0.006108f
C688 B.n635 VSUBS 0.006108f
C689 B.n636 VSUBS 0.006108f
C690 B.n637 VSUBS 0.006108f
C691 B.n638 VSUBS 0.006108f
C692 B.n639 VSUBS 0.006108f
C693 B.n640 VSUBS 0.006108f
C694 B.n641 VSUBS 0.006108f
C695 B.n642 VSUBS 0.006108f
C696 B.n643 VSUBS 0.006108f
C697 B.n644 VSUBS 0.006108f
C698 B.n645 VSUBS 0.006108f
C699 B.n646 VSUBS 0.006108f
C700 B.n647 VSUBS 0.006108f
C701 B.n648 VSUBS 0.006108f
C702 B.n649 VSUBS 0.006108f
C703 B.n650 VSUBS 0.006108f
C704 B.n651 VSUBS 0.006108f
C705 B.n652 VSUBS 0.006108f
C706 B.n653 VSUBS 0.006108f
C707 B.n654 VSUBS 0.006108f
C708 B.n655 VSUBS 0.006108f
C709 B.n656 VSUBS 0.006108f
C710 B.n657 VSUBS 0.006108f
C711 B.n658 VSUBS 0.006108f
C712 B.n659 VSUBS 0.006108f
C713 B.n660 VSUBS 0.006108f
C714 B.n661 VSUBS 0.006108f
C715 B.n662 VSUBS 0.006108f
C716 B.n663 VSUBS 0.006108f
C717 B.n664 VSUBS 0.006108f
C718 B.n665 VSUBS 0.006108f
C719 B.n666 VSUBS 0.006108f
C720 B.n667 VSUBS 0.006108f
C721 B.n668 VSUBS 0.006108f
C722 B.n669 VSUBS 0.006108f
C723 B.n670 VSUBS 0.006108f
C724 B.n671 VSUBS 0.006108f
C725 B.n672 VSUBS 0.006108f
C726 B.n673 VSUBS 0.006108f
C727 B.n674 VSUBS 0.006108f
C728 B.n675 VSUBS 0.006108f
C729 B.n676 VSUBS 0.006108f
C730 B.n677 VSUBS 0.006108f
C731 B.n678 VSUBS 0.006108f
C732 B.n679 VSUBS 0.006108f
C733 B.n680 VSUBS 0.006108f
C734 B.n681 VSUBS 0.006108f
C735 B.n682 VSUBS 0.006108f
C736 B.n683 VSUBS 0.006108f
C737 B.n684 VSUBS 0.006108f
C738 B.n685 VSUBS 0.006108f
C739 B.n686 VSUBS 0.006108f
C740 B.n687 VSUBS 0.006108f
C741 B.n688 VSUBS 0.006108f
C742 B.n689 VSUBS 0.006108f
C743 B.n690 VSUBS 0.006108f
C744 B.n691 VSUBS 0.006108f
C745 B.n692 VSUBS 0.006108f
C746 B.n693 VSUBS 0.006108f
C747 B.n694 VSUBS 0.006108f
C748 B.n695 VSUBS 0.006108f
C749 B.n696 VSUBS 0.006108f
C750 B.n697 VSUBS 0.006108f
C751 B.n698 VSUBS 0.006108f
C752 B.n699 VSUBS 0.006108f
C753 B.n700 VSUBS 0.006108f
C754 B.n701 VSUBS 0.006108f
C755 B.n702 VSUBS 0.006108f
C756 B.n703 VSUBS 0.006108f
C757 B.n704 VSUBS 0.006108f
C758 B.n705 VSUBS 0.006108f
C759 B.n706 VSUBS 0.006108f
C760 B.n707 VSUBS 0.006108f
C761 B.n708 VSUBS 0.005749f
C762 B.n709 VSUBS 0.006108f
C763 B.n710 VSUBS 0.006108f
C764 B.n711 VSUBS 0.006108f
C765 B.n712 VSUBS 0.006108f
C766 B.n713 VSUBS 0.006108f
C767 B.n714 VSUBS 0.006108f
C768 B.n715 VSUBS 0.006108f
C769 B.n716 VSUBS 0.006108f
C770 B.n717 VSUBS 0.006108f
C771 B.n718 VSUBS 0.006108f
C772 B.n719 VSUBS 0.006108f
C773 B.n720 VSUBS 0.006108f
C774 B.n721 VSUBS 0.006108f
C775 B.n722 VSUBS 0.006108f
C776 B.n723 VSUBS 0.006108f
C777 B.n724 VSUBS 0.003414f
C778 B.n725 VSUBS 0.014152f
C779 B.n726 VSUBS 0.005749f
C780 B.n727 VSUBS 0.006108f
C781 B.n728 VSUBS 0.006108f
C782 B.n729 VSUBS 0.006108f
C783 B.n730 VSUBS 0.006108f
C784 B.n731 VSUBS 0.006108f
C785 B.n732 VSUBS 0.006108f
C786 B.n733 VSUBS 0.006108f
C787 B.n734 VSUBS 0.006108f
C788 B.n735 VSUBS 0.006108f
C789 B.n736 VSUBS 0.006108f
C790 B.n737 VSUBS 0.006108f
C791 B.n738 VSUBS 0.006108f
C792 B.n739 VSUBS 0.006108f
C793 B.n740 VSUBS 0.006108f
C794 B.n741 VSUBS 0.006108f
C795 B.n742 VSUBS 0.006108f
C796 B.n743 VSUBS 0.006108f
C797 B.n744 VSUBS 0.006108f
C798 B.n745 VSUBS 0.006108f
C799 B.n746 VSUBS 0.006108f
C800 B.n747 VSUBS 0.006108f
C801 B.n748 VSUBS 0.006108f
C802 B.n749 VSUBS 0.006108f
C803 B.n750 VSUBS 0.006108f
C804 B.n751 VSUBS 0.006108f
C805 B.n752 VSUBS 0.006108f
C806 B.n753 VSUBS 0.006108f
C807 B.n754 VSUBS 0.006108f
C808 B.n755 VSUBS 0.006108f
C809 B.n756 VSUBS 0.006108f
C810 B.n757 VSUBS 0.006108f
C811 B.n758 VSUBS 0.006108f
C812 B.n759 VSUBS 0.006108f
C813 B.n760 VSUBS 0.006108f
C814 B.n761 VSUBS 0.006108f
C815 B.n762 VSUBS 0.006108f
C816 B.n763 VSUBS 0.006108f
C817 B.n764 VSUBS 0.006108f
C818 B.n765 VSUBS 0.006108f
C819 B.n766 VSUBS 0.006108f
C820 B.n767 VSUBS 0.006108f
C821 B.n768 VSUBS 0.006108f
C822 B.n769 VSUBS 0.006108f
C823 B.n770 VSUBS 0.006108f
C824 B.n771 VSUBS 0.006108f
C825 B.n772 VSUBS 0.006108f
C826 B.n773 VSUBS 0.006108f
C827 B.n774 VSUBS 0.006108f
C828 B.n775 VSUBS 0.006108f
C829 B.n776 VSUBS 0.006108f
C830 B.n777 VSUBS 0.006108f
C831 B.n778 VSUBS 0.006108f
C832 B.n779 VSUBS 0.006108f
C833 B.n780 VSUBS 0.006108f
C834 B.n781 VSUBS 0.006108f
C835 B.n782 VSUBS 0.006108f
C836 B.n783 VSUBS 0.006108f
C837 B.n784 VSUBS 0.006108f
C838 B.n785 VSUBS 0.006108f
C839 B.n786 VSUBS 0.006108f
C840 B.n787 VSUBS 0.006108f
C841 B.n788 VSUBS 0.006108f
C842 B.n789 VSUBS 0.006108f
C843 B.n790 VSUBS 0.006108f
C844 B.n791 VSUBS 0.006108f
C845 B.n792 VSUBS 0.006108f
C846 B.n793 VSUBS 0.006108f
C847 B.n794 VSUBS 0.006108f
C848 B.n795 VSUBS 0.006108f
C849 B.n796 VSUBS 0.006108f
C850 B.n797 VSUBS 0.006108f
C851 B.n798 VSUBS 0.006108f
C852 B.n799 VSUBS 0.006108f
C853 B.n800 VSUBS 0.006108f
C854 B.n801 VSUBS 0.006108f
C855 B.n802 VSUBS 0.006108f
C856 B.n803 VSUBS 0.006108f
C857 B.n804 VSUBS 0.006108f
C858 B.n805 VSUBS 0.006108f
C859 B.n806 VSUBS 0.006108f
C860 B.n807 VSUBS 0.006108f
C861 B.n808 VSUBS 0.006108f
C862 B.n809 VSUBS 0.006108f
C863 B.n810 VSUBS 0.006108f
C864 B.n811 VSUBS 0.006108f
C865 B.n812 VSUBS 0.006108f
C866 B.n813 VSUBS 0.006108f
C867 B.n814 VSUBS 0.006108f
C868 B.n815 VSUBS 0.006108f
C869 B.n816 VSUBS 0.006108f
C870 B.n817 VSUBS 0.006108f
C871 B.n818 VSUBS 0.006108f
C872 B.n819 VSUBS 0.014295f
C873 B.n820 VSUBS 0.013732f
C874 B.n821 VSUBS 0.013732f
C875 B.n822 VSUBS 0.006108f
C876 B.n823 VSUBS 0.006108f
C877 B.n824 VSUBS 0.006108f
C878 B.n825 VSUBS 0.006108f
C879 B.n826 VSUBS 0.006108f
C880 B.n827 VSUBS 0.006108f
C881 B.n828 VSUBS 0.006108f
C882 B.n829 VSUBS 0.006108f
C883 B.n830 VSUBS 0.006108f
C884 B.n831 VSUBS 0.006108f
C885 B.n832 VSUBS 0.006108f
C886 B.n833 VSUBS 0.006108f
C887 B.n834 VSUBS 0.006108f
C888 B.n835 VSUBS 0.006108f
C889 B.n836 VSUBS 0.006108f
C890 B.n837 VSUBS 0.006108f
C891 B.n838 VSUBS 0.006108f
C892 B.n839 VSUBS 0.006108f
C893 B.n840 VSUBS 0.006108f
C894 B.n841 VSUBS 0.006108f
C895 B.n842 VSUBS 0.006108f
C896 B.n843 VSUBS 0.006108f
C897 B.n844 VSUBS 0.006108f
C898 B.n845 VSUBS 0.006108f
C899 B.n846 VSUBS 0.006108f
C900 B.n847 VSUBS 0.006108f
C901 B.n848 VSUBS 0.006108f
C902 B.n849 VSUBS 0.006108f
C903 B.n850 VSUBS 0.006108f
C904 B.n851 VSUBS 0.006108f
C905 B.n852 VSUBS 0.006108f
C906 B.n853 VSUBS 0.006108f
C907 B.n854 VSUBS 0.006108f
C908 B.n855 VSUBS 0.006108f
C909 B.n856 VSUBS 0.006108f
C910 B.n857 VSUBS 0.006108f
C911 B.n858 VSUBS 0.006108f
C912 B.n859 VSUBS 0.006108f
C913 B.n860 VSUBS 0.006108f
C914 B.n861 VSUBS 0.006108f
C915 B.n862 VSUBS 0.006108f
C916 B.n863 VSUBS 0.006108f
C917 B.n864 VSUBS 0.006108f
C918 B.n865 VSUBS 0.006108f
C919 B.n866 VSUBS 0.006108f
C920 B.n867 VSUBS 0.006108f
C921 B.n868 VSUBS 0.006108f
C922 B.n869 VSUBS 0.006108f
C923 B.n870 VSUBS 0.006108f
C924 B.n871 VSUBS 0.006108f
C925 B.n872 VSUBS 0.006108f
C926 B.n873 VSUBS 0.006108f
C927 B.n874 VSUBS 0.006108f
C928 B.n875 VSUBS 0.006108f
C929 B.n876 VSUBS 0.006108f
C930 B.n877 VSUBS 0.006108f
C931 B.n878 VSUBS 0.006108f
C932 B.n879 VSUBS 0.007971f
C933 B.n880 VSUBS 0.008491f
C934 B.n881 VSUBS 0.016886f
C935 VDD1.t1 VSUBS 0.411215f
C936 VDD1.t0 VSUBS 0.411215f
C937 VDD1.n0 VSUBS 3.44795f
C938 VDD1.t2 VSUBS 0.411215f
C939 VDD1.t3 VSUBS 0.411215f
C940 VDD1.n1 VSUBS 4.54366f
C941 VTAIL.t3 VSUBS 3.57264f
C942 VTAIL.n0 VSUBS 0.813492f
C943 VTAIL.t6 VSUBS 3.57264f
C944 VTAIL.n1 VSUBS 0.923519f
C945 VTAIL.t7 VSUBS 3.57264f
C946 VTAIL.n2 VSUBS 2.63121f
C947 VTAIL.t1 VSUBS 3.57264f
C948 VTAIL.n3 VSUBS 2.6312f
C949 VTAIL.t2 VSUBS 3.57264f
C950 VTAIL.n4 VSUBS 0.923513f
C951 VTAIL.t5 VSUBS 3.57264f
C952 VTAIL.n5 VSUBS 0.923513f
C953 VTAIL.t4 VSUBS 3.57264f
C954 VTAIL.n6 VSUBS 2.63121f
C955 VTAIL.t0 VSUBS 3.57264f
C956 VTAIL.n7 VSUBS 2.51275f
C957 VP.t0 VSUBS 4.8991f
C958 VP.n0 VSUBS 1.79925f
C959 VP.n1 VSUBS 0.027606f
C960 VP.n2 VSUBS 0.022316f
C961 VP.n3 VSUBS 0.027606f
C962 VP.t1 VSUBS 4.8991f
C963 VP.n4 VSUBS 1.79925f
C964 VP.t2 VSUBS 5.27864f
C965 VP.t3 VSUBS 5.26688f
C966 VP.n5 VSUBS 5.21563f
C967 VP.n6 VSUBS 1.86996f
C968 VP.n7 VSUBS 0.044555f
C969 VP.n8 VSUBS 0.042813f
C970 VP.n9 VSUBS 0.05145f
C971 VP.n10 VSUBS 0.054866f
C972 VP.n11 VSUBS 0.027606f
C973 VP.n12 VSUBS 0.027606f
C974 VP.n13 VSUBS 0.027606f
C975 VP.n14 VSUBS 0.054866f
C976 VP.n15 VSUBS 0.05145f
C977 VP.n16 VSUBS 0.042813f
C978 VP.n17 VSUBS 0.044555f
C979 VP.n18 VSUBS 0.065438f
.ends

