* NGSPICE file created from diff_pair_sample_0221.ext - technology: sky130A

.subckt diff_pair_sample_0221 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2626_n1462# sky130_fd_pr__pfet_01v8 ad=0.9633 pd=5.72 as=0 ps=0 w=2.47 l=3.81
X1 B.t8 B.t6 B.t7 w_n2626_n1462# sky130_fd_pr__pfet_01v8 ad=0.9633 pd=5.72 as=0 ps=0 w=2.47 l=3.81
X2 B.t5 B.t3 B.t4 w_n2626_n1462# sky130_fd_pr__pfet_01v8 ad=0.9633 pd=5.72 as=0 ps=0 w=2.47 l=3.81
X3 VDD1.t1 VP.t0 VTAIL.t3 w_n2626_n1462# sky130_fd_pr__pfet_01v8 ad=0.9633 pd=5.72 as=0.9633 ps=5.72 w=2.47 l=3.81
X4 VDD2.t1 VN.t0 VTAIL.t1 w_n2626_n1462# sky130_fd_pr__pfet_01v8 ad=0.9633 pd=5.72 as=0.9633 ps=5.72 w=2.47 l=3.81
X5 VDD1.t0 VP.t1 VTAIL.t2 w_n2626_n1462# sky130_fd_pr__pfet_01v8 ad=0.9633 pd=5.72 as=0.9633 ps=5.72 w=2.47 l=3.81
X6 VDD2.t0 VN.t1 VTAIL.t0 w_n2626_n1462# sky130_fd_pr__pfet_01v8 ad=0.9633 pd=5.72 as=0.9633 ps=5.72 w=2.47 l=3.81
X7 B.t2 B.t0 B.t1 w_n2626_n1462# sky130_fd_pr__pfet_01v8 ad=0.9633 pd=5.72 as=0 ps=0 w=2.47 l=3.81
R0 B.n215 B.n214 585
R1 B.n213 B.n74 585
R2 B.n212 B.n211 585
R3 B.n210 B.n75 585
R4 B.n209 B.n208 585
R5 B.n207 B.n76 585
R6 B.n206 B.n205 585
R7 B.n204 B.n77 585
R8 B.n203 B.n202 585
R9 B.n201 B.n78 585
R10 B.n200 B.n199 585
R11 B.n198 B.n79 585
R12 B.n197 B.n196 585
R13 B.n195 B.n80 585
R14 B.n194 B.n193 585
R15 B.n189 B.n81 585
R16 B.n188 B.n187 585
R17 B.n186 B.n82 585
R18 B.n185 B.n184 585
R19 B.n183 B.n83 585
R20 B.n182 B.n181 585
R21 B.n180 B.n84 585
R22 B.n179 B.n178 585
R23 B.n176 B.n85 585
R24 B.n175 B.n174 585
R25 B.n173 B.n88 585
R26 B.n172 B.n171 585
R27 B.n170 B.n89 585
R28 B.n169 B.n168 585
R29 B.n167 B.n90 585
R30 B.n166 B.n165 585
R31 B.n164 B.n91 585
R32 B.n163 B.n162 585
R33 B.n161 B.n92 585
R34 B.n160 B.n159 585
R35 B.n158 B.n93 585
R36 B.n157 B.n156 585
R37 B.n216 B.n73 585
R38 B.n218 B.n217 585
R39 B.n219 B.n72 585
R40 B.n221 B.n220 585
R41 B.n222 B.n71 585
R42 B.n224 B.n223 585
R43 B.n225 B.n70 585
R44 B.n227 B.n226 585
R45 B.n228 B.n69 585
R46 B.n230 B.n229 585
R47 B.n231 B.n68 585
R48 B.n233 B.n232 585
R49 B.n234 B.n67 585
R50 B.n236 B.n235 585
R51 B.n237 B.n66 585
R52 B.n239 B.n238 585
R53 B.n240 B.n65 585
R54 B.n242 B.n241 585
R55 B.n243 B.n64 585
R56 B.n245 B.n244 585
R57 B.n246 B.n63 585
R58 B.n248 B.n247 585
R59 B.n249 B.n62 585
R60 B.n251 B.n250 585
R61 B.n252 B.n61 585
R62 B.n254 B.n253 585
R63 B.n255 B.n60 585
R64 B.n257 B.n256 585
R65 B.n258 B.n59 585
R66 B.n260 B.n259 585
R67 B.n261 B.n58 585
R68 B.n263 B.n262 585
R69 B.n264 B.n57 585
R70 B.n266 B.n265 585
R71 B.n267 B.n56 585
R72 B.n269 B.n268 585
R73 B.n270 B.n55 585
R74 B.n272 B.n271 585
R75 B.n273 B.n54 585
R76 B.n275 B.n274 585
R77 B.n276 B.n53 585
R78 B.n278 B.n277 585
R79 B.n279 B.n52 585
R80 B.n281 B.n280 585
R81 B.n282 B.n51 585
R82 B.n284 B.n283 585
R83 B.n285 B.n50 585
R84 B.n287 B.n286 585
R85 B.n288 B.n49 585
R86 B.n290 B.n289 585
R87 B.n291 B.n48 585
R88 B.n293 B.n292 585
R89 B.n294 B.n47 585
R90 B.n296 B.n295 585
R91 B.n297 B.n46 585
R92 B.n299 B.n298 585
R93 B.n300 B.n45 585
R94 B.n302 B.n301 585
R95 B.n303 B.n44 585
R96 B.n305 B.n304 585
R97 B.n306 B.n43 585
R98 B.n308 B.n307 585
R99 B.n309 B.n42 585
R100 B.n311 B.n310 585
R101 B.n312 B.n41 585
R102 B.n314 B.n313 585
R103 B.n371 B.n18 585
R104 B.n370 B.n369 585
R105 B.n368 B.n19 585
R106 B.n367 B.n366 585
R107 B.n365 B.n20 585
R108 B.n364 B.n363 585
R109 B.n362 B.n21 585
R110 B.n361 B.n360 585
R111 B.n359 B.n22 585
R112 B.n358 B.n357 585
R113 B.n356 B.n23 585
R114 B.n355 B.n354 585
R115 B.n353 B.n24 585
R116 B.n352 B.n351 585
R117 B.n349 B.n25 585
R118 B.n348 B.n347 585
R119 B.n346 B.n28 585
R120 B.n345 B.n344 585
R121 B.n343 B.n29 585
R122 B.n342 B.n341 585
R123 B.n340 B.n30 585
R124 B.n339 B.n338 585
R125 B.n337 B.n31 585
R126 B.n335 B.n334 585
R127 B.n333 B.n34 585
R128 B.n332 B.n331 585
R129 B.n330 B.n35 585
R130 B.n329 B.n328 585
R131 B.n327 B.n36 585
R132 B.n326 B.n325 585
R133 B.n324 B.n37 585
R134 B.n323 B.n322 585
R135 B.n321 B.n38 585
R136 B.n320 B.n319 585
R137 B.n318 B.n39 585
R138 B.n317 B.n316 585
R139 B.n315 B.n40 585
R140 B.n373 B.n372 585
R141 B.n374 B.n17 585
R142 B.n376 B.n375 585
R143 B.n377 B.n16 585
R144 B.n379 B.n378 585
R145 B.n380 B.n15 585
R146 B.n382 B.n381 585
R147 B.n383 B.n14 585
R148 B.n385 B.n384 585
R149 B.n386 B.n13 585
R150 B.n388 B.n387 585
R151 B.n389 B.n12 585
R152 B.n391 B.n390 585
R153 B.n392 B.n11 585
R154 B.n394 B.n393 585
R155 B.n395 B.n10 585
R156 B.n397 B.n396 585
R157 B.n398 B.n9 585
R158 B.n400 B.n399 585
R159 B.n401 B.n8 585
R160 B.n403 B.n402 585
R161 B.n404 B.n7 585
R162 B.n406 B.n405 585
R163 B.n407 B.n6 585
R164 B.n409 B.n408 585
R165 B.n410 B.n5 585
R166 B.n412 B.n411 585
R167 B.n413 B.n4 585
R168 B.n415 B.n414 585
R169 B.n416 B.n3 585
R170 B.n418 B.n417 585
R171 B.n419 B.n0 585
R172 B.n2 B.n1 585
R173 B.n110 B.n109 585
R174 B.n112 B.n111 585
R175 B.n113 B.n108 585
R176 B.n115 B.n114 585
R177 B.n116 B.n107 585
R178 B.n118 B.n117 585
R179 B.n119 B.n106 585
R180 B.n121 B.n120 585
R181 B.n122 B.n105 585
R182 B.n124 B.n123 585
R183 B.n125 B.n104 585
R184 B.n127 B.n126 585
R185 B.n128 B.n103 585
R186 B.n130 B.n129 585
R187 B.n131 B.n102 585
R188 B.n133 B.n132 585
R189 B.n134 B.n101 585
R190 B.n136 B.n135 585
R191 B.n137 B.n100 585
R192 B.n139 B.n138 585
R193 B.n140 B.n99 585
R194 B.n142 B.n141 585
R195 B.n143 B.n98 585
R196 B.n145 B.n144 585
R197 B.n146 B.n97 585
R198 B.n148 B.n147 585
R199 B.n149 B.n96 585
R200 B.n151 B.n150 585
R201 B.n152 B.n95 585
R202 B.n154 B.n153 585
R203 B.n155 B.n94 585
R204 B.n156 B.n155 473.281
R205 B.n214 B.n73 473.281
R206 B.n315 B.n314 473.281
R207 B.n372 B.n371 473.281
R208 B.n190 B.t10 303.961
R209 B.n32 B.t8 303.961
R210 B.n86 B.t4 303.961
R211 B.n26 B.t2 303.961
R212 B.n421 B.n420 256.663
R213 B.n420 B.n419 235.042
R214 B.n420 B.n2 235.042
R215 B.n86 B.t3 224.976
R216 B.n190 B.t9 224.976
R217 B.n32 B.t6 224.976
R218 B.n26 B.t0 224.976
R219 B.n191 B.t11 223.669
R220 B.n33 B.t7 223.669
R221 B.n87 B.t5 223.669
R222 B.n27 B.t1 223.669
R223 B.n156 B.n93 163.367
R224 B.n160 B.n93 163.367
R225 B.n161 B.n160 163.367
R226 B.n162 B.n161 163.367
R227 B.n162 B.n91 163.367
R228 B.n166 B.n91 163.367
R229 B.n167 B.n166 163.367
R230 B.n168 B.n167 163.367
R231 B.n168 B.n89 163.367
R232 B.n172 B.n89 163.367
R233 B.n173 B.n172 163.367
R234 B.n174 B.n173 163.367
R235 B.n174 B.n85 163.367
R236 B.n179 B.n85 163.367
R237 B.n180 B.n179 163.367
R238 B.n181 B.n180 163.367
R239 B.n181 B.n83 163.367
R240 B.n185 B.n83 163.367
R241 B.n186 B.n185 163.367
R242 B.n187 B.n186 163.367
R243 B.n187 B.n81 163.367
R244 B.n194 B.n81 163.367
R245 B.n195 B.n194 163.367
R246 B.n196 B.n195 163.367
R247 B.n196 B.n79 163.367
R248 B.n200 B.n79 163.367
R249 B.n201 B.n200 163.367
R250 B.n202 B.n201 163.367
R251 B.n202 B.n77 163.367
R252 B.n206 B.n77 163.367
R253 B.n207 B.n206 163.367
R254 B.n208 B.n207 163.367
R255 B.n208 B.n75 163.367
R256 B.n212 B.n75 163.367
R257 B.n213 B.n212 163.367
R258 B.n214 B.n213 163.367
R259 B.n314 B.n41 163.367
R260 B.n310 B.n41 163.367
R261 B.n310 B.n309 163.367
R262 B.n309 B.n308 163.367
R263 B.n308 B.n43 163.367
R264 B.n304 B.n43 163.367
R265 B.n304 B.n303 163.367
R266 B.n303 B.n302 163.367
R267 B.n302 B.n45 163.367
R268 B.n298 B.n45 163.367
R269 B.n298 B.n297 163.367
R270 B.n297 B.n296 163.367
R271 B.n296 B.n47 163.367
R272 B.n292 B.n47 163.367
R273 B.n292 B.n291 163.367
R274 B.n291 B.n290 163.367
R275 B.n290 B.n49 163.367
R276 B.n286 B.n49 163.367
R277 B.n286 B.n285 163.367
R278 B.n285 B.n284 163.367
R279 B.n284 B.n51 163.367
R280 B.n280 B.n51 163.367
R281 B.n280 B.n279 163.367
R282 B.n279 B.n278 163.367
R283 B.n278 B.n53 163.367
R284 B.n274 B.n53 163.367
R285 B.n274 B.n273 163.367
R286 B.n273 B.n272 163.367
R287 B.n272 B.n55 163.367
R288 B.n268 B.n55 163.367
R289 B.n268 B.n267 163.367
R290 B.n267 B.n266 163.367
R291 B.n266 B.n57 163.367
R292 B.n262 B.n57 163.367
R293 B.n262 B.n261 163.367
R294 B.n261 B.n260 163.367
R295 B.n260 B.n59 163.367
R296 B.n256 B.n59 163.367
R297 B.n256 B.n255 163.367
R298 B.n255 B.n254 163.367
R299 B.n254 B.n61 163.367
R300 B.n250 B.n61 163.367
R301 B.n250 B.n249 163.367
R302 B.n249 B.n248 163.367
R303 B.n248 B.n63 163.367
R304 B.n244 B.n63 163.367
R305 B.n244 B.n243 163.367
R306 B.n243 B.n242 163.367
R307 B.n242 B.n65 163.367
R308 B.n238 B.n65 163.367
R309 B.n238 B.n237 163.367
R310 B.n237 B.n236 163.367
R311 B.n236 B.n67 163.367
R312 B.n232 B.n67 163.367
R313 B.n232 B.n231 163.367
R314 B.n231 B.n230 163.367
R315 B.n230 B.n69 163.367
R316 B.n226 B.n69 163.367
R317 B.n226 B.n225 163.367
R318 B.n225 B.n224 163.367
R319 B.n224 B.n71 163.367
R320 B.n220 B.n71 163.367
R321 B.n220 B.n219 163.367
R322 B.n219 B.n218 163.367
R323 B.n218 B.n73 163.367
R324 B.n371 B.n370 163.367
R325 B.n370 B.n19 163.367
R326 B.n366 B.n19 163.367
R327 B.n366 B.n365 163.367
R328 B.n365 B.n364 163.367
R329 B.n364 B.n21 163.367
R330 B.n360 B.n21 163.367
R331 B.n360 B.n359 163.367
R332 B.n359 B.n358 163.367
R333 B.n358 B.n23 163.367
R334 B.n354 B.n23 163.367
R335 B.n354 B.n353 163.367
R336 B.n353 B.n352 163.367
R337 B.n352 B.n25 163.367
R338 B.n347 B.n25 163.367
R339 B.n347 B.n346 163.367
R340 B.n346 B.n345 163.367
R341 B.n345 B.n29 163.367
R342 B.n341 B.n29 163.367
R343 B.n341 B.n340 163.367
R344 B.n340 B.n339 163.367
R345 B.n339 B.n31 163.367
R346 B.n334 B.n31 163.367
R347 B.n334 B.n333 163.367
R348 B.n333 B.n332 163.367
R349 B.n332 B.n35 163.367
R350 B.n328 B.n35 163.367
R351 B.n328 B.n327 163.367
R352 B.n327 B.n326 163.367
R353 B.n326 B.n37 163.367
R354 B.n322 B.n37 163.367
R355 B.n322 B.n321 163.367
R356 B.n321 B.n320 163.367
R357 B.n320 B.n39 163.367
R358 B.n316 B.n39 163.367
R359 B.n316 B.n315 163.367
R360 B.n372 B.n17 163.367
R361 B.n376 B.n17 163.367
R362 B.n377 B.n376 163.367
R363 B.n378 B.n377 163.367
R364 B.n378 B.n15 163.367
R365 B.n382 B.n15 163.367
R366 B.n383 B.n382 163.367
R367 B.n384 B.n383 163.367
R368 B.n384 B.n13 163.367
R369 B.n388 B.n13 163.367
R370 B.n389 B.n388 163.367
R371 B.n390 B.n389 163.367
R372 B.n390 B.n11 163.367
R373 B.n394 B.n11 163.367
R374 B.n395 B.n394 163.367
R375 B.n396 B.n395 163.367
R376 B.n396 B.n9 163.367
R377 B.n400 B.n9 163.367
R378 B.n401 B.n400 163.367
R379 B.n402 B.n401 163.367
R380 B.n402 B.n7 163.367
R381 B.n406 B.n7 163.367
R382 B.n407 B.n406 163.367
R383 B.n408 B.n407 163.367
R384 B.n408 B.n5 163.367
R385 B.n412 B.n5 163.367
R386 B.n413 B.n412 163.367
R387 B.n414 B.n413 163.367
R388 B.n414 B.n3 163.367
R389 B.n418 B.n3 163.367
R390 B.n419 B.n418 163.367
R391 B.n109 B.n2 163.367
R392 B.n112 B.n109 163.367
R393 B.n113 B.n112 163.367
R394 B.n114 B.n113 163.367
R395 B.n114 B.n107 163.367
R396 B.n118 B.n107 163.367
R397 B.n119 B.n118 163.367
R398 B.n120 B.n119 163.367
R399 B.n120 B.n105 163.367
R400 B.n124 B.n105 163.367
R401 B.n125 B.n124 163.367
R402 B.n126 B.n125 163.367
R403 B.n126 B.n103 163.367
R404 B.n130 B.n103 163.367
R405 B.n131 B.n130 163.367
R406 B.n132 B.n131 163.367
R407 B.n132 B.n101 163.367
R408 B.n136 B.n101 163.367
R409 B.n137 B.n136 163.367
R410 B.n138 B.n137 163.367
R411 B.n138 B.n99 163.367
R412 B.n142 B.n99 163.367
R413 B.n143 B.n142 163.367
R414 B.n144 B.n143 163.367
R415 B.n144 B.n97 163.367
R416 B.n148 B.n97 163.367
R417 B.n149 B.n148 163.367
R418 B.n150 B.n149 163.367
R419 B.n150 B.n95 163.367
R420 B.n154 B.n95 163.367
R421 B.n155 B.n154 163.367
R422 B.n87 B.n86 80.2914
R423 B.n191 B.n190 80.2914
R424 B.n33 B.n32 80.2914
R425 B.n27 B.n26 80.2914
R426 B.n177 B.n87 59.5399
R427 B.n192 B.n191 59.5399
R428 B.n336 B.n33 59.5399
R429 B.n350 B.n27 59.5399
R430 B.n373 B.n18 30.7517
R431 B.n313 B.n40 30.7517
R432 B.n216 B.n215 30.7517
R433 B.n157 B.n94 30.7517
R434 B B.n421 18.0485
R435 B.n374 B.n373 10.6151
R436 B.n375 B.n374 10.6151
R437 B.n375 B.n16 10.6151
R438 B.n379 B.n16 10.6151
R439 B.n380 B.n379 10.6151
R440 B.n381 B.n380 10.6151
R441 B.n381 B.n14 10.6151
R442 B.n385 B.n14 10.6151
R443 B.n386 B.n385 10.6151
R444 B.n387 B.n386 10.6151
R445 B.n387 B.n12 10.6151
R446 B.n391 B.n12 10.6151
R447 B.n392 B.n391 10.6151
R448 B.n393 B.n392 10.6151
R449 B.n393 B.n10 10.6151
R450 B.n397 B.n10 10.6151
R451 B.n398 B.n397 10.6151
R452 B.n399 B.n398 10.6151
R453 B.n399 B.n8 10.6151
R454 B.n403 B.n8 10.6151
R455 B.n404 B.n403 10.6151
R456 B.n405 B.n404 10.6151
R457 B.n405 B.n6 10.6151
R458 B.n409 B.n6 10.6151
R459 B.n410 B.n409 10.6151
R460 B.n411 B.n410 10.6151
R461 B.n411 B.n4 10.6151
R462 B.n415 B.n4 10.6151
R463 B.n416 B.n415 10.6151
R464 B.n417 B.n416 10.6151
R465 B.n417 B.n0 10.6151
R466 B.n369 B.n18 10.6151
R467 B.n369 B.n368 10.6151
R468 B.n368 B.n367 10.6151
R469 B.n367 B.n20 10.6151
R470 B.n363 B.n20 10.6151
R471 B.n363 B.n362 10.6151
R472 B.n362 B.n361 10.6151
R473 B.n361 B.n22 10.6151
R474 B.n357 B.n22 10.6151
R475 B.n357 B.n356 10.6151
R476 B.n356 B.n355 10.6151
R477 B.n355 B.n24 10.6151
R478 B.n351 B.n24 10.6151
R479 B.n349 B.n348 10.6151
R480 B.n348 B.n28 10.6151
R481 B.n344 B.n28 10.6151
R482 B.n344 B.n343 10.6151
R483 B.n343 B.n342 10.6151
R484 B.n342 B.n30 10.6151
R485 B.n338 B.n30 10.6151
R486 B.n338 B.n337 10.6151
R487 B.n335 B.n34 10.6151
R488 B.n331 B.n34 10.6151
R489 B.n331 B.n330 10.6151
R490 B.n330 B.n329 10.6151
R491 B.n329 B.n36 10.6151
R492 B.n325 B.n36 10.6151
R493 B.n325 B.n324 10.6151
R494 B.n324 B.n323 10.6151
R495 B.n323 B.n38 10.6151
R496 B.n319 B.n38 10.6151
R497 B.n319 B.n318 10.6151
R498 B.n318 B.n317 10.6151
R499 B.n317 B.n40 10.6151
R500 B.n313 B.n312 10.6151
R501 B.n312 B.n311 10.6151
R502 B.n311 B.n42 10.6151
R503 B.n307 B.n42 10.6151
R504 B.n307 B.n306 10.6151
R505 B.n306 B.n305 10.6151
R506 B.n305 B.n44 10.6151
R507 B.n301 B.n44 10.6151
R508 B.n301 B.n300 10.6151
R509 B.n300 B.n299 10.6151
R510 B.n299 B.n46 10.6151
R511 B.n295 B.n46 10.6151
R512 B.n295 B.n294 10.6151
R513 B.n294 B.n293 10.6151
R514 B.n293 B.n48 10.6151
R515 B.n289 B.n48 10.6151
R516 B.n289 B.n288 10.6151
R517 B.n288 B.n287 10.6151
R518 B.n287 B.n50 10.6151
R519 B.n283 B.n50 10.6151
R520 B.n283 B.n282 10.6151
R521 B.n282 B.n281 10.6151
R522 B.n281 B.n52 10.6151
R523 B.n277 B.n52 10.6151
R524 B.n277 B.n276 10.6151
R525 B.n276 B.n275 10.6151
R526 B.n275 B.n54 10.6151
R527 B.n271 B.n54 10.6151
R528 B.n271 B.n270 10.6151
R529 B.n270 B.n269 10.6151
R530 B.n269 B.n56 10.6151
R531 B.n265 B.n56 10.6151
R532 B.n265 B.n264 10.6151
R533 B.n264 B.n263 10.6151
R534 B.n263 B.n58 10.6151
R535 B.n259 B.n58 10.6151
R536 B.n259 B.n258 10.6151
R537 B.n258 B.n257 10.6151
R538 B.n257 B.n60 10.6151
R539 B.n253 B.n60 10.6151
R540 B.n253 B.n252 10.6151
R541 B.n252 B.n251 10.6151
R542 B.n251 B.n62 10.6151
R543 B.n247 B.n62 10.6151
R544 B.n247 B.n246 10.6151
R545 B.n246 B.n245 10.6151
R546 B.n245 B.n64 10.6151
R547 B.n241 B.n64 10.6151
R548 B.n241 B.n240 10.6151
R549 B.n240 B.n239 10.6151
R550 B.n239 B.n66 10.6151
R551 B.n235 B.n66 10.6151
R552 B.n235 B.n234 10.6151
R553 B.n234 B.n233 10.6151
R554 B.n233 B.n68 10.6151
R555 B.n229 B.n68 10.6151
R556 B.n229 B.n228 10.6151
R557 B.n228 B.n227 10.6151
R558 B.n227 B.n70 10.6151
R559 B.n223 B.n70 10.6151
R560 B.n223 B.n222 10.6151
R561 B.n222 B.n221 10.6151
R562 B.n221 B.n72 10.6151
R563 B.n217 B.n72 10.6151
R564 B.n217 B.n216 10.6151
R565 B.n110 B.n1 10.6151
R566 B.n111 B.n110 10.6151
R567 B.n111 B.n108 10.6151
R568 B.n115 B.n108 10.6151
R569 B.n116 B.n115 10.6151
R570 B.n117 B.n116 10.6151
R571 B.n117 B.n106 10.6151
R572 B.n121 B.n106 10.6151
R573 B.n122 B.n121 10.6151
R574 B.n123 B.n122 10.6151
R575 B.n123 B.n104 10.6151
R576 B.n127 B.n104 10.6151
R577 B.n128 B.n127 10.6151
R578 B.n129 B.n128 10.6151
R579 B.n129 B.n102 10.6151
R580 B.n133 B.n102 10.6151
R581 B.n134 B.n133 10.6151
R582 B.n135 B.n134 10.6151
R583 B.n135 B.n100 10.6151
R584 B.n139 B.n100 10.6151
R585 B.n140 B.n139 10.6151
R586 B.n141 B.n140 10.6151
R587 B.n141 B.n98 10.6151
R588 B.n145 B.n98 10.6151
R589 B.n146 B.n145 10.6151
R590 B.n147 B.n146 10.6151
R591 B.n147 B.n96 10.6151
R592 B.n151 B.n96 10.6151
R593 B.n152 B.n151 10.6151
R594 B.n153 B.n152 10.6151
R595 B.n153 B.n94 10.6151
R596 B.n158 B.n157 10.6151
R597 B.n159 B.n158 10.6151
R598 B.n159 B.n92 10.6151
R599 B.n163 B.n92 10.6151
R600 B.n164 B.n163 10.6151
R601 B.n165 B.n164 10.6151
R602 B.n165 B.n90 10.6151
R603 B.n169 B.n90 10.6151
R604 B.n170 B.n169 10.6151
R605 B.n171 B.n170 10.6151
R606 B.n171 B.n88 10.6151
R607 B.n175 B.n88 10.6151
R608 B.n176 B.n175 10.6151
R609 B.n178 B.n84 10.6151
R610 B.n182 B.n84 10.6151
R611 B.n183 B.n182 10.6151
R612 B.n184 B.n183 10.6151
R613 B.n184 B.n82 10.6151
R614 B.n188 B.n82 10.6151
R615 B.n189 B.n188 10.6151
R616 B.n193 B.n189 10.6151
R617 B.n197 B.n80 10.6151
R618 B.n198 B.n197 10.6151
R619 B.n199 B.n198 10.6151
R620 B.n199 B.n78 10.6151
R621 B.n203 B.n78 10.6151
R622 B.n204 B.n203 10.6151
R623 B.n205 B.n204 10.6151
R624 B.n205 B.n76 10.6151
R625 B.n209 B.n76 10.6151
R626 B.n210 B.n209 10.6151
R627 B.n211 B.n210 10.6151
R628 B.n211 B.n74 10.6151
R629 B.n215 B.n74 10.6151
R630 B.n421 B.n0 8.11757
R631 B.n421 B.n1 8.11757
R632 B.n350 B.n349 6.5566
R633 B.n337 B.n336 6.5566
R634 B.n178 B.n177 6.5566
R635 B.n193 B.n192 6.5566
R636 B.n351 B.n350 4.05904
R637 B.n336 B.n335 4.05904
R638 B.n177 B.n176 4.05904
R639 B.n192 B.n80 4.05904
R640 VP.n0 VP.t0 91.307
R641 VP.n0 VP.t1 50.6615
R642 VP VP.n0 0.621237
R643 VTAIL.n42 VTAIL.n36 756.745
R644 VTAIL.n6 VTAIL.n0 756.745
R645 VTAIL.n30 VTAIL.n24 756.745
R646 VTAIL.n18 VTAIL.n12 756.745
R647 VTAIL.n41 VTAIL.n40 585
R648 VTAIL.n43 VTAIL.n42 585
R649 VTAIL.n5 VTAIL.n4 585
R650 VTAIL.n7 VTAIL.n6 585
R651 VTAIL.n31 VTAIL.n30 585
R652 VTAIL.n29 VTAIL.n28 585
R653 VTAIL.n19 VTAIL.n18 585
R654 VTAIL.n17 VTAIL.n16 585
R655 VTAIL.n39 VTAIL.t1 355.474
R656 VTAIL.n3 VTAIL.t2 355.474
R657 VTAIL.n27 VTAIL.t3 355.474
R658 VTAIL.n15 VTAIL.t0 355.474
R659 VTAIL.n42 VTAIL.n41 171.744
R660 VTAIL.n6 VTAIL.n5 171.744
R661 VTAIL.n30 VTAIL.n29 171.744
R662 VTAIL.n18 VTAIL.n17 171.744
R663 VTAIL.n41 VTAIL.t1 85.8723
R664 VTAIL.n5 VTAIL.t2 85.8723
R665 VTAIL.n29 VTAIL.t3 85.8723
R666 VTAIL.n17 VTAIL.t0 85.8723
R667 VTAIL.n47 VTAIL.n46 33.5429
R668 VTAIL.n11 VTAIL.n10 33.5429
R669 VTAIL.n35 VTAIL.n34 33.5429
R670 VTAIL.n23 VTAIL.n22 33.5429
R671 VTAIL.n23 VTAIL.n11 21.6341
R672 VTAIL.n47 VTAIL.n35 18.0652
R673 VTAIL.n40 VTAIL.n39 15.8418
R674 VTAIL.n4 VTAIL.n3 15.8418
R675 VTAIL.n28 VTAIL.n27 15.8418
R676 VTAIL.n16 VTAIL.n15 15.8418
R677 VTAIL.n43 VTAIL.n38 12.8005
R678 VTAIL.n7 VTAIL.n2 12.8005
R679 VTAIL.n31 VTAIL.n26 12.8005
R680 VTAIL.n19 VTAIL.n14 12.8005
R681 VTAIL.n44 VTAIL.n36 12.0247
R682 VTAIL.n8 VTAIL.n0 12.0247
R683 VTAIL.n32 VTAIL.n24 12.0247
R684 VTAIL.n20 VTAIL.n12 12.0247
R685 VTAIL.n46 VTAIL.n45 9.45567
R686 VTAIL.n10 VTAIL.n9 9.45567
R687 VTAIL.n34 VTAIL.n33 9.45567
R688 VTAIL.n22 VTAIL.n21 9.45567
R689 VTAIL.n45 VTAIL.n44 9.3005
R690 VTAIL.n38 VTAIL.n37 9.3005
R691 VTAIL.n9 VTAIL.n8 9.3005
R692 VTAIL.n2 VTAIL.n1 9.3005
R693 VTAIL.n33 VTAIL.n32 9.3005
R694 VTAIL.n26 VTAIL.n25 9.3005
R695 VTAIL.n21 VTAIL.n20 9.3005
R696 VTAIL.n14 VTAIL.n13 9.3005
R697 VTAIL.n27 VTAIL.n25 4.29255
R698 VTAIL.n15 VTAIL.n13 4.29255
R699 VTAIL.n39 VTAIL.n37 4.29255
R700 VTAIL.n3 VTAIL.n1 4.29255
R701 VTAIL.n35 VTAIL.n23 2.25481
R702 VTAIL.n46 VTAIL.n36 1.93989
R703 VTAIL.n10 VTAIL.n0 1.93989
R704 VTAIL.n34 VTAIL.n24 1.93989
R705 VTAIL.n22 VTAIL.n12 1.93989
R706 VTAIL VTAIL.n11 1.42076
R707 VTAIL.n44 VTAIL.n43 1.16414
R708 VTAIL.n8 VTAIL.n7 1.16414
R709 VTAIL.n32 VTAIL.n31 1.16414
R710 VTAIL.n20 VTAIL.n19 1.16414
R711 VTAIL VTAIL.n47 0.834552
R712 VTAIL.n40 VTAIL.n38 0.388379
R713 VTAIL.n4 VTAIL.n2 0.388379
R714 VTAIL.n28 VTAIL.n26 0.388379
R715 VTAIL.n16 VTAIL.n14 0.388379
R716 VTAIL.n45 VTAIL.n37 0.155672
R717 VTAIL.n9 VTAIL.n1 0.155672
R718 VTAIL.n33 VTAIL.n25 0.155672
R719 VTAIL.n21 VTAIL.n13 0.155672
R720 VDD1.n6 VDD1.n0 756.745
R721 VDD1.n17 VDD1.n11 756.745
R722 VDD1.n7 VDD1.n6 585
R723 VDD1.n5 VDD1.n4 585
R724 VDD1.n16 VDD1.n15 585
R725 VDD1.n18 VDD1.n17 585
R726 VDD1.n3 VDD1.t1 355.474
R727 VDD1.n14 VDD1.t0 355.474
R728 VDD1.n6 VDD1.n5 171.744
R729 VDD1.n17 VDD1.n16 171.744
R730 VDD1.n5 VDD1.t1 85.8723
R731 VDD1.n16 VDD1.t0 85.8723
R732 VDD1 VDD1.n21 84.5655
R733 VDD1 VDD1.n10 51.1721
R734 VDD1.n4 VDD1.n3 15.8418
R735 VDD1.n15 VDD1.n14 15.8418
R736 VDD1.n7 VDD1.n2 12.8005
R737 VDD1.n18 VDD1.n13 12.8005
R738 VDD1.n8 VDD1.n0 12.0247
R739 VDD1.n19 VDD1.n11 12.0247
R740 VDD1.n10 VDD1.n9 9.45567
R741 VDD1.n21 VDD1.n20 9.45567
R742 VDD1.n9 VDD1.n8 9.3005
R743 VDD1.n2 VDD1.n1 9.3005
R744 VDD1.n20 VDD1.n19 9.3005
R745 VDD1.n13 VDD1.n12 9.3005
R746 VDD1.n3 VDD1.n1 4.29255
R747 VDD1.n14 VDD1.n12 4.29255
R748 VDD1.n10 VDD1.n0 1.93989
R749 VDD1.n21 VDD1.n11 1.93989
R750 VDD1.n8 VDD1.n7 1.16414
R751 VDD1.n19 VDD1.n18 1.16414
R752 VDD1.n4 VDD1.n2 0.388379
R753 VDD1.n15 VDD1.n13 0.388379
R754 VDD1.n9 VDD1.n1 0.155672
R755 VDD1.n20 VDD1.n12 0.155672
R756 VN VN.t1 91.1193
R757 VN VN.t0 51.2822
R758 VDD2.n17 VDD2.n11 756.745
R759 VDD2.n6 VDD2.n0 756.745
R760 VDD2.n18 VDD2.n17 585
R761 VDD2.n16 VDD2.n15 585
R762 VDD2.n5 VDD2.n4 585
R763 VDD2.n7 VDD2.n6 585
R764 VDD2.n14 VDD2.t0 355.474
R765 VDD2.n3 VDD2.t1 355.474
R766 VDD2.n17 VDD2.n16 171.744
R767 VDD2.n6 VDD2.n5 171.744
R768 VDD2.n16 VDD2.t0 85.8723
R769 VDD2.n5 VDD2.t1 85.8723
R770 VDD2.n22 VDD2.n10 83.1484
R771 VDD2.n22 VDD2.n21 50.2217
R772 VDD2.n15 VDD2.n14 15.8418
R773 VDD2.n4 VDD2.n3 15.8418
R774 VDD2.n18 VDD2.n13 12.8005
R775 VDD2.n7 VDD2.n2 12.8005
R776 VDD2.n19 VDD2.n11 12.0247
R777 VDD2.n8 VDD2.n0 12.0247
R778 VDD2.n21 VDD2.n20 9.45567
R779 VDD2.n10 VDD2.n9 9.45567
R780 VDD2.n20 VDD2.n19 9.3005
R781 VDD2.n13 VDD2.n12 9.3005
R782 VDD2.n9 VDD2.n8 9.3005
R783 VDD2.n2 VDD2.n1 9.3005
R784 VDD2.n14 VDD2.n12 4.29255
R785 VDD2.n3 VDD2.n1 4.29255
R786 VDD2.n21 VDD2.n11 1.93989
R787 VDD2.n10 VDD2.n0 1.93989
R788 VDD2.n19 VDD2.n18 1.16414
R789 VDD2.n8 VDD2.n7 1.16414
R790 VDD2 VDD2.n22 0.950931
R791 VDD2.n15 VDD2.n13 0.388379
R792 VDD2.n4 VDD2.n2 0.388379
R793 VDD2.n20 VDD2.n12 0.155672
R794 VDD2.n9 VDD2.n1 0.155672
C0 VTAIL B 1.70971f
C1 VTAIL VDD2 3.00311f
C2 VP VN 4.26762f
C3 VP VDD1 1.04388f
C4 VN VDD1 0.154361f
C5 w_n2626_n1462# VTAIL 1.4579f
C6 B VP 1.66484f
C7 B VN 1.10634f
C8 B VDD1 1.09362f
C9 VP VDD2 0.389637f
C10 VDD2 VN 0.810153f
C11 VDD2 VDD1 0.808495f
C12 B VDD2 1.13495f
C13 w_n2626_n1462# VP 3.88518f
C14 w_n2626_n1462# VN 3.55135f
C15 w_n2626_n1462# VDD1 1.262f
C16 w_n2626_n1462# B 7.48746f
C17 w_n2626_n1462# VDD2 1.30214f
C18 VTAIL VP 1.2204f
C19 VTAIL VN 1.20616f
C20 VTAIL VDD1 2.94195f
C21 VDD2 VSUBS 0.687017f
C22 VDD1 VSUBS 2.577103f
C23 VTAIL VSUBS 0.425776f
C24 VN VSUBS 6.194269f
C25 VP VSUBS 1.579219f
C26 B VSUBS 3.773052f
C27 w_n2626_n1462# VSUBS 48.812103f
C28 VDD2.n0 VSUBS 0.018605f
C29 VDD2.n1 VSUBS 0.124714f
C30 VDD2.n2 VSUBS 0.009617f
C31 VDD2.t1 VSUBS 0.050278f
C32 VDD2.n3 VSUBS 0.058922f
C33 VDD2.n4 VSUBS 0.013403f
C34 VDD2.n5 VSUBS 0.017049f
C35 VDD2.n6 VSUBS 0.051417f
C36 VDD2.n7 VSUBS 0.010183f
C37 VDD2.n8 VSUBS 0.009617f
C38 VDD2.n9 VSUBS 0.043081f
C39 VDD2.n10 VSUBS 0.349516f
C40 VDD2.n11 VSUBS 0.018605f
C41 VDD2.n12 VSUBS 0.124714f
C42 VDD2.n13 VSUBS 0.009617f
C43 VDD2.t0 VSUBS 0.050278f
C44 VDD2.n14 VSUBS 0.058922f
C45 VDD2.n15 VSUBS 0.013403f
C46 VDD2.n16 VSUBS 0.017049f
C47 VDD2.n17 VSUBS 0.051417f
C48 VDD2.n18 VSUBS 0.010183f
C49 VDD2.n19 VSUBS 0.009617f
C50 VDD2.n20 VSUBS 0.043081f
C51 VDD2.n21 VSUBS 0.038093f
C52 VDD2.n22 VSUBS 1.6404f
C53 VN.t0 VSUBS 1.54565f
C54 VN.t1 VSUBS 2.58821f
C55 VDD1.n0 VSUBS 0.017597f
C56 VDD1.n1 VSUBS 0.117957f
C57 VDD1.n2 VSUBS 0.009096f
C58 VDD1.t1 VSUBS 0.047554f
C59 VDD1.n3 VSUBS 0.05573f
C60 VDD1.n4 VSUBS 0.012677f
C61 VDD1.n5 VSUBS 0.016125f
C62 VDD1.n6 VSUBS 0.048632f
C63 VDD1.n7 VSUBS 0.009631f
C64 VDD1.n8 VSUBS 0.009096f
C65 VDD1.n9 VSUBS 0.040747f
C66 VDD1.n10 VSUBS 0.037615f
C67 VDD1.n11 VSUBS 0.017597f
C68 VDD1.n12 VSUBS 0.117957f
C69 VDD1.n13 VSUBS 0.009096f
C70 VDD1.t0 VSUBS 0.047554f
C71 VDD1.n14 VSUBS 0.05573f
C72 VDD1.n15 VSUBS 0.012677f
C73 VDD1.n16 VSUBS 0.016125f
C74 VDD1.n17 VSUBS 0.048632f
C75 VDD1.n18 VSUBS 0.009631f
C76 VDD1.n19 VSUBS 0.009096f
C77 VDD1.n20 VSUBS 0.040747f
C78 VDD1.n21 VSUBS 0.363368f
C79 VTAIL.n0 VSUBS 0.021891f
C80 VTAIL.n1 VSUBS 0.146746f
C81 VTAIL.n2 VSUBS 0.011316f
C82 VTAIL.t2 VSUBS 0.059161f
C83 VTAIL.n3 VSUBS 0.069331f
C84 VTAIL.n4 VSUBS 0.015771f
C85 VTAIL.n5 VSUBS 0.020061f
C86 VTAIL.n6 VSUBS 0.060501f
C87 VTAIL.n7 VSUBS 0.011982f
C88 VTAIL.n8 VSUBS 0.011316f
C89 VTAIL.n9 VSUBS 0.050692f
C90 VTAIL.n10 VSUBS 0.030297f
C91 VTAIL.n11 VSUBS 1.03043f
C92 VTAIL.n12 VSUBS 0.021891f
C93 VTAIL.n13 VSUBS 0.146746f
C94 VTAIL.n14 VSUBS 0.011316f
C95 VTAIL.t0 VSUBS 0.059161f
C96 VTAIL.n15 VSUBS 0.069331f
C97 VTAIL.n16 VSUBS 0.015771f
C98 VTAIL.n17 VSUBS 0.020061f
C99 VTAIL.n18 VSUBS 0.060501f
C100 VTAIL.n19 VSUBS 0.011982f
C101 VTAIL.n20 VSUBS 0.011316f
C102 VTAIL.n21 VSUBS 0.050692f
C103 VTAIL.n22 VSUBS 0.030297f
C104 VTAIL.n23 VSUBS 1.08702f
C105 VTAIL.n24 VSUBS 0.021891f
C106 VTAIL.n25 VSUBS 0.146746f
C107 VTAIL.n26 VSUBS 0.011316f
C108 VTAIL.t3 VSUBS 0.059161f
C109 VTAIL.n27 VSUBS 0.069331f
C110 VTAIL.n28 VSUBS 0.015771f
C111 VTAIL.n29 VSUBS 0.020061f
C112 VTAIL.n30 VSUBS 0.060501f
C113 VTAIL.n31 VSUBS 0.011982f
C114 VTAIL.n32 VSUBS 0.011316f
C115 VTAIL.n33 VSUBS 0.050692f
C116 VTAIL.n34 VSUBS 0.030297f
C117 VTAIL.n35 VSUBS 0.844841f
C118 VTAIL.n36 VSUBS 0.021891f
C119 VTAIL.n37 VSUBS 0.146746f
C120 VTAIL.n38 VSUBS 0.011316f
C121 VTAIL.t1 VSUBS 0.059161f
C122 VTAIL.n39 VSUBS 0.069331f
C123 VTAIL.n40 VSUBS 0.015771f
C124 VTAIL.n41 VSUBS 0.020061f
C125 VTAIL.n42 VSUBS 0.060501f
C126 VTAIL.n43 VSUBS 0.011982f
C127 VTAIL.n44 VSUBS 0.011316f
C128 VTAIL.n45 VSUBS 0.050692f
C129 VTAIL.n46 VSUBS 0.030297f
C130 VTAIL.n47 VSUBS 0.748464f
C131 VP.t0 VSUBS 2.70906f
C132 VP.t1 VSUBS 1.60933f
C133 VP.n0 VSUBS 3.68653f
C134 B.n0 VSUBS 0.007615f
C135 B.n1 VSUBS 0.007615f
C136 B.n2 VSUBS 0.011262f
C137 B.n3 VSUBS 0.00863f
C138 B.n4 VSUBS 0.00863f
C139 B.n5 VSUBS 0.00863f
C140 B.n6 VSUBS 0.00863f
C141 B.n7 VSUBS 0.00863f
C142 B.n8 VSUBS 0.00863f
C143 B.n9 VSUBS 0.00863f
C144 B.n10 VSUBS 0.00863f
C145 B.n11 VSUBS 0.00863f
C146 B.n12 VSUBS 0.00863f
C147 B.n13 VSUBS 0.00863f
C148 B.n14 VSUBS 0.00863f
C149 B.n15 VSUBS 0.00863f
C150 B.n16 VSUBS 0.00863f
C151 B.n17 VSUBS 0.00863f
C152 B.n18 VSUBS 0.020012f
C153 B.n19 VSUBS 0.00863f
C154 B.n20 VSUBS 0.00863f
C155 B.n21 VSUBS 0.00863f
C156 B.n22 VSUBS 0.00863f
C157 B.n23 VSUBS 0.00863f
C158 B.n24 VSUBS 0.00863f
C159 B.n25 VSUBS 0.00863f
C160 B.t1 VSUBS 0.047144f
C161 B.t2 VSUBS 0.071599f
C162 B.t0 VSUBS 0.571878f
C163 B.n26 VSUBS 0.127887f
C164 B.n27 VSUBS 0.104888f
C165 B.n28 VSUBS 0.00863f
C166 B.n29 VSUBS 0.00863f
C167 B.n30 VSUBS 0.00863f
C168 B.n31 VSUBS 0.00863f
C169 B.t7 VSUBS 0.047145f
C170 B.t8 VSUBS 0.071599f
C171 B.t6 VSUBS 0.571878f
C172 B.n32 VSUBS 0.127887f
C173 B.n33 VSUBS 0.104887f
C174 B.n34 VSUBS 0.00863f
C175 B.n35 VSUBS 0.00863f
C176 B.n36 VSUBS 0.00863f
C177 B.n37 VSUBS 0.00863f
C178 B.n38 VSUBS 0.00863f
C179 B.n39 VSUBS 0.00863f
C180 B.n40 VSUBS 0.020012f
C181 B.n41 VSUBS 0.00863f
C182 B.n42 VSUBS 0.00863f
C183 B.n43 VSUBS 0.00863f
C184 B.n44 VSUBS 0.00863f
C185 B.n45 VSUBS 0.00863f
C186 B.n46 VSUBS 0.00863f
C187 B.n47 VSUBS 0.00863f
C188 B.n48 VSUBS 0.00863f
C189 B.n49 VSUBS 0.00863f
C190 B.n50 VSUBS 0.00863f
C191 B.n51 VSUBS 0.00863f
C192 B.n52 VSUBS 0.00863f
C193 B.n53 VSUBS 0.00863f
C194 B.n54 VSUBS 0.00863f
C195 B.n55 VSUBS 0.00863f
C196 B.n56 VSUBS 0.00863f
C197 B.n57 VSUBS 0.00863f
C198 B.n58 VSUBS 0.00863f
C199 B.n59 VSUBS 0.00863f
C200 B.n60 VSUBS 0.00863f
C201 B.n61 VSUBS 0.00863f
C202 B.n62 VSUBS 0.00863f
C203 B.n63 VSUBS 0.00863f
C204 B.n64 VSUBS 0.00863f
C205 B.n65 VSUBS 0.00863f
C206 B.n66 VSUBS 0.00863f
C207 B.n67 VSUBS 0.00863f
C208 B.n68 VSUBS 0.00863f
C209 B.n69 VSUBS 0.00863f
C210 B.n70 VSUBS 0.00863f
C211 B.n71 VSUBS 0.00863f
C212 B.n72 VSUBS 0.00863f
C213 B.n73 VSUBS 0.018823f
C214 B.n74 VSUBS 0.00863f
C215 B.n75 VSUBS 0.00863f
C216 B.n76 VSUBS 0.00863f
C217 B.n77 VSUBS 0.00863f
C218 B.n78 VSUBS 0.00863f
C219 B.n79 VSUBS 0.00863f
C220 B.n80 VSUBS 0.005965f
C221 B.n81 VSUBS 0.00863f
C222 B.n82 VSUBS 0.00863f
C223 B.n83 VSUBS 0.00863f
C224 B.n84 VSUBS 0.00863f
C225 B.n85 VSUBS 0.00863f
C226 B.t5 VSUBS 0.047144f
C227 B.t4 VSUBS 0.071599f
C228 B.t3 VSUBS 0.571878f
C229 B.n86 VSUBS 0.127887f
C230 B.n87 VSUBS 0.104888f
C231 B.n88 VSUBS 0.00863f
C232 B.n89 VSUBS 0.00863f
C233 B.n90 VSUBS 0.00863f
C234 B.n91 VSUBS 0.00863f
C235 B.n92 VSUBS 0.00863f
C236 B.n93 VSUBS 0.00863f
C237 B.n94 VSUBS 0.018823f
C238 B.n95 VSUBS 0.00863f
C239 B.n96 VSUBS 0.00863f
C240 B.n97 VSUBS 0.00863f
C241 B.n98 VSUBS 0.00863f
C242 B.n99 VSUBS 0.00863f
C243 B.n100 VSUBS 0.00863f
C244 B.n101 VSUBS 0.00863f
C245 B.n102 VSUBS 0.00863f
C246 B.n103 VSUBS 0.00863f
C247 B.n104 VSUBS 0.00863f
C248 B.n105 VSUBS 0.00863f
C249 B.n106 VSUBS 0.00863f
C250 B.n107 VSUBS 0.00863f
C251 B.n108 VSUBS 0.00863f
C252 B.n109 VSUBS 0.00863f
C253 B.n110 VSUBS 0.00863f
C254 B.n111 VSUBS 0.00863f
C255 B.n112 VSUBS 0.00863f
C256 B.n113 VSUBS 0.00863f
C257 B.n114 VSUBS 0.00863f
C258 B.n115 VSUBS 0.00863f
C259 B.n116 VSUBS 0.00863f
C260 B.n117 VSUBS 0.00863f
C261 B.n118 VSUBS 0.00863f
C262 B.n119 VSUBS 0.00863f
C263 B.n120 VSUBS 0.00863f
C264 B.n121 VSUBS 0.00863f
C265 B.n122 VSUBS 0.00863f
C266 B.n123 VSUBS 0.00863f
C267 B.n124 VSUBS 0.00863f
C268 B.n125 VSUBS 0.00863f
C269 B.n126 VSUBS 0.00863f
C270 B.n127 VSUBS 0.00863f
C271 B.n128 VSUBS 0.00863f
C272 B.n129 VSUBS 0.00863f
C273 B.n130 VSUBS 0.00863f
C274 B.n131 VSUBS 0.00863f
C275 B.n132 VSUBS 0.00863f
C276 B.n133 VSUBS 0.00863f
C277 B.n134 VSUBS 0.00863f
C278 B.n135 VSUBS 0.00863f
C279 B.n136 VSUBS 0.00863f
C280 B.n137 VSUBS 0.00863f
C281 B.n138 VSUBS 0.00863f
C282 B.n139 VSUBS 0.00863f
C283 B.n140 VSUBS 0.00863f
C284 B.n141 VSUBS 0.00863f
C285 B.n142 VSUBS 0.00863f
C286 B.n143 VSUBS 0.00863f
C287 B.n144 VSUBS 0.00863f
C288 B.n145 VSUBS 0.00863f
C289 B.n146 VSUBS 0.00863f
C290 B.n147 VSUBS 0.00863f
C291 B.n148 VSUBS 0.00863f
C292 B.n149 VSUBS 0.00863f
C293 B.n150 VSUBS 0.00863f
C294 B.n151 VSUBS 0.00863f
C295 B.n152 VSUBS 0.00863f
C296 B.n153 VSUBS 0.00863f
C297 B.n154 VSUBS 0.00863f
C298 B.n155 VSUBS 0.018823f
C299 B.n156 VSUBS 0.020012f
C300 B.n157 VSUBS 0.020012f
C301 B.n158 VSUBS 0.00863f
C302 B.n159 VSUBS 0.00863f
C303 B.n160 VSUBS 0.00863f
C304 B.n161 VSUBS 0.00863f
C305 B.n162 VSUBS 0.00863f
C306 B.n163 VSUBS 0.00863f
C307 B.n164 VSUBS 0.00863f
C308 B.n165 VSUBS 0.00863f
C309 B.n166 VSUBS 0.00863f
C310 B.n167 VSUBS 0.00863f
C311 B.n168 VSUBS 0.00863f
C312 B.n169 VSUBS 0.00863f
C313 B.n170 VSUBS 0.00863f
C314 B.n171 VSUBS 0.00863f
C315 B.n172 VSUBS 0.00863f
C316 B.n173 VSUBS 0.00863f
C317 B.n174 VSUBS 0.00863f
C318 B.n175 VSUBS 0.00863f
C319 B.n176 VSUBS 0.005965f
C320 B.n177 VSUBS 0.019995f
C321 B.n178 VSUBS 0.00698f
C322 B.n179 VSUBS 0.00863f
C323 B.n180 VSUBS 0.00863f
C324 B.n181 VSUBS 0.00863f
C325 B.n182 VSUBS 0.00863f
C326 B.n183 VSUBS 0.00863f
C327 B.n184 VSUBS 0.00863f
C328 B.n185 VSUBS 0.00863f
C329 B.n186 VSUBS 0.00863f
C330 B.n187 VSUBS 0.00863f
C331 B.n188 VSUBS 0.00863f
C332 B.n189 VSUBS 0.00863f
C333 B.t11 VSUBS 0.047145f
C334 B.t10 VSUBS 0.071599f
C335 B.t9 VSUBS 0.571878f
C336 B.n190 VSUBS 0.127887f
C337 B.n191 VSUBS 0.104887f
C338 B.n192 VSUBS 0.019995f
C339 B.n193 VSUBS 0.00698f
C340 B.n194 VSUBS 0.00863f
C341 B.n195 VSUBS 0.00863f
C342 B.n196 VSUBS 0.00863f
C343 B.n197 VSUBS 0.00863f
C344 B.n198 VSUBS 0.00863f
C345 B.n199 VSUBS 0.00863f
C346 B.n200 VSUBS 0.00863f
C347 B.n201 VSUBS 0.00863f
C348 B.n202 VSUBS 0.00863f
C349 B.n203 VSUBS 0.00863f
C350 B.n204 VSUBS 0.00863f
C351 B.n205 VSUBS 0.00863f
C352 B.n206 VSUBS 0.00863f
C353 B.n207 VSUBS 0.00863f
C354 B.n208 VSUBS 0.00863f
C355 B.n209 VSUBS 0.00863f
C356 B.n210 VSUBS 0.00863f
C357 B.n211 VSUBS 0.00863f
C358 B.n212 VSUBS 0.00863f
C359 B.n213 VSUBS 0.00863f
C360 B.n214 VSUBS 0.020012f
C361 B.n215 VSUBS 0.018929f
C362 B.n216 VSUBS 0.019907f
C363 B.n217 VSUBS 0.00863f
C364 B.n218 VSUBS 0.00863f
C365 B.n219 VSUBS 0.00863f
C366 B.n220 VSUBS 0.00863f
C367 B.n221 VSUBS 0.00863f
C368 B.n222 VSUBS 0.00863f
C369 B.n223 VSUBS 0.00863f
C370 B.n224 VSUBS 0.00863f
C371 B.n225 VSUBS 0.00863f
C372 B.n226 VSUBS 0.00863f
C373 B.n227 VSUBS 0.00863f
C374 B.n228 VSUBS 0.00863f
C375 B.n229 VSUBS 0.00863f
C376 B.n230 VSUBS 0.00863f
C377 B.n231 VSUBS 0.00863f
C378 B.n232 VSUBS 0.00863f
C379 B.n233 VSUBS 0.00863f
C380 B.n234 VSUBS 0.00863f
C381 B.n235 VSUBS 0.00863f
C382 B.n236 VSUBS 0.00863f
C383 B.n237 VSUBS 0.00863f
C384 B.n238 VSUBS 0.00863f
C385 B.n239 VSUBS 0.00863f
C386 B.n240 VSUBS 0.00863f
C387 B.n241 VSUBS 0.00863f
C388 B.n242 VSUBS 0.00863f
C389 B.n243 VSUBS 0.00863f
C390 B.n244 VSUBS 0.00863f
C391 B.n245 VSUBS 0.00863f
C392 B.n246 VSUBS 0.00863f
C393 B.n247 VSUBS 0.00863f
C394 B.n248 VSUBS 0.00863f
C395 B.n249 VSUBS 0.00863f
C396 B.n250 VSUBS 0.00863f
C397 B.n251 VSUBS 0.00863f
C398 B.n252 VSUBS 0.00863f
C399 B.n253 VSUBS 0.00863f
C400 B.n254 VSUBS 0.00863f
C401 B.n255 VSUBS 0.00863f
C402 B.n256 VSUBS 0.00863f
C403 B.n257 VSUBS 0.00863f
C404 B.n258 VSUBS 0.00863f
C405 B.n259 VSUBS 0.00863f
C406 B.n260 VSUBS 0.00863f
C407 B.n261 VSUBS 0.00863f
C408 B.n262 VSUBS 0.00863f
C409 B.n263 VSUBS 0.00863f
C410 B.n264 VSUBS 0.00863f
C411 B.n265 VSUBS 0.00863f
C412 B.n266 VSUBS 0.00863f
C413 B.n267 VSUBS 0.00863f
C414 B.n268 VSUBS 0.00863f
C415 B.n269 VSUBS 0.00863f
C416 B.n270 VSUBS 0.00863f
C417 B.n271 VSUBS 0.00863f
C418 B.n272 VSUBS 0.00863f
C419 B.n273 VSUBS 0.00863f
C420 B.n274 VSUBS 0.00863f
C421 B.n275 VSUBS 0.00863f
C422 B.n276 VSUBS 0.00863f
C423 B.n277 VSUBS 0.00863f
C424 B.n278 VSUBS 0.00863f
C425 B.n279 VSUBS 0.00863f
C426 B.n280 VSUBS 0.00863f
C427 B.n281 VSUBS 0.00863f
C428 B.n282 VSUBS 0.00863f
C429 B.n283 VSUBS 0.00863f
C430 B.n284 VSUBS 0.00863f
C431 B.n285 VSUBS 0.00863f
C432 B.n286 VSUBS 0.00863f
C433 B.n287 VSUBS 0.00863f
C434 B.n288 VSUBS 0.00863f
C435 B.n289 VSUBS 0.00863f
C436 B.n290 VSUBS 0.00863f
C437 B.n291 VSUBS 0.00863f
C438 B.n292 VSUBS 0.00863f
C439 B.n293 VSUBS 0.00863f
C440 B.n294 VSUBS 0.00863f
C441 B.n295 VSUBS 0.00863f
C442 B.n296 VSUBS 0.00863f
C443 B.n297 VSUBS 0.00863f
C444 B.n298 VSUBS 0.00863f
C445 B.n299 VSUBS 0.00863f
C446 B.n300 VSUBS 0.00863f
C447 B.n301 VSUBS 0.00863f
C448 B.n302 VSUBS 0.00863f
C449 B.n303 VSUBS 0.00863f
C450 B.n304 VSUBS 0.00863f
C451 B.n305 VSUBS 0.00863f
C452 B.n306 VSUBS 0.00863f
C453 B.n307 VSUBS 0.00863f
C454 B.n308 VSUBS 0.00863f
C455 B.n309 VSUBS 0.00863f
C456 B.n310 VSUBS 0.00863f
C457 B.n311 VSUBS 0.00863f
C458 B.n312 VSUBS 0.00863f
C459 B.n313 VSUBS 0.018823f
C460 B.n314 VSUBS 0.018823f
C461 B.n315 VSUBS 0.020012f
C462 B.n316 VSUBS 0.00863f
C463 B.n317 VSUBS 0.00863f
C464 B.n318 VSUBS 0.00863f
C465 B.n319 VSUBS 0.00863f
C466 B.n320 VSUBS 0.00863f
C467 B.n321 VSUBS 0.00863f
C468 B.n322 VSUBS 0.00863f
C469 B.n323 VSUBS 0.00863f
C470 B.n324 VSUBS 0.00863f
C471 B.n325 VSUBS 0.00863f
C472 B.n326 VSUBS 0.00863f
C473 B.n327 VSUBS 0.00863f
C474 B.n328 VSUBS 0.00863f
C475 B.n329 VSUBS 0.00863f
C476 B.n330 VSUBS 0.00863f
C477 B.n331 VSUBS 0.00863f
C478 B.n332 VSUBS 0.00863f
C479 B.n333 VSUBS 0.00863f
C480 B.n334 VSUBS 0.00863f
C481 B.n335 VSUBS 0.005965f
C482 B.n336 VSUBS 0.019995f
C483 B.n337 VSUBS 0.00698f
C484 B.n338 VSUBS 0.00863f
C485 B.n339 VSUBS 0.00863f
C486 B.n340 VSUBS 0.00863f
C487 B.n341 VSUBS 0.00863f
C488 B.n342 VSUBS 0.00863f
C489 B.n343 VSUBS 0.00863f
C490 B.n344 VSUBS 0.00863f
C491 B.n345 VSUBS 0.00863f
C492 B.n346 VSUBS 0.00863f
C493 B.n347 VSUBS 0.00863f
C494 B.n348 VSUBS 0.00863f
C495 B.n349 VSUBS 0.00698f
C496 B.n350 VSUBS 0.019995f
C497 B.n351 VSUBS 0.005965f
C498 B.n352 VSUBS 0.00863f
C499 B.n353 VSUBS 0.00863f
C500 B.n354 VSUBS 0.00863f
C501 B.n355 VSUBS 0.00863f
C502 B.n356 VSUBS 0.00863f
C503 B.n357 VSUBS 0.00863f
C504 B.n358 VSUBS 0.00863f
C505 B.n359 VSUBS 0.00863f
C506 B.n360 VSUBS 0.00863f
C507 B.n361 VSUBS 0.00863f
C508 B.n362 VSUBS 0.00863f
C509 B.n363 VSUBS 0.00863f
C510 B.n364 VSUBS 0.00863f
C511 B.n365 VSUBS 0.00863f
C512 B.n366 VSUBS 0.00863f
C513 B.n367 VSUBS 0.00863f
C514 B.n368 VSUBS 0.00863f
C515 B.n369 VSUBS 0.00863f
C516 B.n370 VSUBS 0.00863f
C517 B.n371 VSUBS 0.020012f
C518 B.n372 VSUBS 0.018823f
C519 B.n373 VSUBS 0.018823f
C520 B.n374 VSUBS 0.00863f
C521 B.n375 VSUBS 0.00863f
C522 B.n376 VSUBS 0.00863f
C523 B.n377 VSUBS 0.00863f
C524 B.n378 VSUBS 0.00863f
C525 B.n379 VSUBS 0.00863f
C526 B.n380 VSUBS 0.00863f
C527 B.n381 VSUBS 0.00863f
C528 B.n382 VSUBS 0.00863f
C529 B.n383 VSUBS 0.00863f
C530 B.n384 VSUBS 0.00863f
C531 B.n385 VSUBS 0.00863f
C532 B.n386 VSUBS 0.00863f
C533 B.n387 VSUBS 0.00863f
C534 B.n388 VSUBS 0.00863f
C535 B.n389 VSUBS 0.00863f
C536 B.n390 VSUBS 0.00863f
C537 B.n391 VSUBS 0.00863f
C538 B.n392 VSUBS 0.00863f
C539 B.n393 VSUBS 0.00863f
C540 B.n394 VSUBS 0.00863f
C541 B.n395 VSUBS 0.00863f
C542 B.n396 VSUBS 0.00863f
C543 B.n397 VSUBS 0.00863f
C544 B.n398 VSUBS 0.00863f
C545 B.n399 VSUBS 0.00863f
C546 B.n400 VSUBS 0.00863f
C547 B.n401 VSUBS 0.00863f
C548 B.n402 VSUBS 0.00863f
C549 B.n403 VSUBS 0.00863f
C550 B.n404 VSUBS 0.00863f
C551 B.n405 VSUBS 0.00863f
C552 B.n406 VSUBS 0.00863f
C553 B.n407 VSUBS 0.00863f
C554 B.n408 VSUBS 0.00863f
C555 B.n409 VSUBS 0.00863f
C556 B.n410 VSUBS 0.00863f
C557 B.n411 VSUBS 0.00863f
C558 B.n412 VSUBS 0.00863f
C559 B.n413 VSUBS 0.00863f
C560 B.n414 VSUBS 0.00863f
C561 B.n415 VSUBS 0.00863f
C562 B.n416 VSUBS 0.00863f
C563 B.n417 VSUBS 0.00863f
C564 B.n418 VSUBS 0.00863f
C565 B.n419 VSUBS 0.011262f
C566 B.n420 VSUBS 0.011997f
C567 B.n421 VSUBS 0.023857f
.ends

