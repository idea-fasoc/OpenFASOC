* NGSPICE file created from diff_pair_sample_0317.ext - technology: sky130A

.subckt diff_pair_sample_0317 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t19 VN.t0 VDD2.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=0.8646 pd=5.57 as=0.8646 ps=5.57 w=5.24 l=3.19
X1 VDD1.t9 VP.t0 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.8646 pd=5.57 as=2.0436 ps=11.26 w=5.24 l=3.19
X2 VTAIL.t18 VN.t1 VDD2.t9 B.t9 sky130_fd_pr__nfet_01v8 ad=0.8646 pd=5.57 as=0.8646 ps=5.57 w=5.24 l=3.19
X3 VTAIL.t17 VN.t2 VDD2.t5 B.t6 sky130_fd_pr__nfet_01v8 ad=0.8646 pd=5.57 as=0.8646 ps=5.57 w=5.24 l=3.19
X4 VDD2.t8 VN.t3 VTAIL.t16 B.t3 sky130_fd_pr__nfet_01v8 ad=0.8646 pd=5.57 as=2.0436 ps=11.26 w=5.24 l=3.19
X5 VDD1.t8 VP.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.8646 pd=5.57 as=0.8646 ps=5.57 w=5.24 l=3.19
X6 VDD2.t4 VN.t4 VTAIL.t15 B.t1 sky130_fd_pr__nfet_01v8 ad=0.8646 pd=5.57 as=0.8646 ps=5.57 w=5.24 l=3.19
X7 VTAIL.t14 VN.t5 VDD2.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=0.8646 pd=5.57 as=0.8646 ps=5.57 w=5.24 l=3.19
X8 VDD2.t0 VN.t6 VTAIL.t13 B.t2 sky130_fd_pr__nfet_01v8 ad=2.0436 pd=11.26 as=0.8646 ps=5.57 w=5.24 l=3.19
X9 B.t23 B.t21 B.t22 B.t15 sky130_fd_pr__nfet_01v8 ad=2.0436 pd=11.26 as=0 ps=0 w=5.24 l=3.19
X10 VDD1.t7 VP.t2 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.0436 pd=11.26 as=0.8646 ps=5.57 w=5.24 l=3.19
X11 B.t20 B.t18 B.t19 B.t11 sky130_fd_pr__nfet_01v8 ad=2.0436 pd=11.26 as=0 ps=0 w=5.24 l=3.19
X12 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=2.0436 pd=11.26 as=0 ps=0 w=5.24 l=3.19
X13 VDD1.t6 VP.t3 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=0.8646 pd=5.57 as=0.8646 ps=5.57 w=5.24 l=3.19
X14 VDD2.t1 VN.t7 VTAIL.t12 B.t8 sky130_fd_pr__nfet_01v8 ad=0.8646 pd=5.57 as=2.0436 ps=11.26 w=5.24 l=3.19
X15 VTAIL.t0 VP.t4 VDD1.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=0.8646 pd=5.57 as=0.8646 ps=5.57 w=5.24 l=3.19
X16 VDD1.t4 VP.t5 VTAIL.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=0.8646 pd=5.57 as=2.0436 ps=11.26 w=5.24 l=3.19
X17 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=2.0436 pd=11.26 as=0 ps=0 w=5.24 l=3.19
X18 VDD1.t3 VP.t6 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=2.0436 pd=11.26 as=0.8646 ps=5.57 w=5.24 l=3.19
X19 VTAIL.t7 VP.t7 VDD1.t2 B.t7 sky130_fd_pr__nfet_01v8 ad=0.8646 pd=5.57 as=0.8646 ps=5.57 w=5.24 l=3.19
X20 VTAIL.t6 VP.t8 VDD1.t1 B.t6 sky130_fd_pr__nfet_01v8 ad=0.8646 pd=5.57 as=0.8646 ps=5.57 w=5.24 l=3.19
X21 VTAIL.t9 VP.t9 VDD1.t0 B.t9 sky130_fd_pr__nfet_01v8 ad=0.8646 pd=5.57 as=0.8646 ps=5.57 w=5.24 l=3.19
X22 VDD2.t2 VN.t8 VTAIL.t11 B.t4 sky130_fd_pr__nfet_01v8 ad=2.0436 pd=11.26 as=0.8646 ps=5.57 w=5.24 l=3.19
X23 VDD2.t6 VN.t9 VTAIL.t10 B.t5 sky130_fd_pr__nfet_01v8 ad=0.8646 pd=5.57 as=0.8646 ps=5.57 w=5.24 l=3.19
R0 VN.n94 VN.n93 161.3
R1 VN.n92 VN.n49 161.3
R2 VN.n91 VN.n90 161.3
R3 VN.n89 VN.n50 161.3
R4 VN.n88 VN.n87 161.3
R5 VN.n86 VN.n51 161.3
R6 VN.n85 VN.n84 161.3
R7 VN.n83 VN.n82 161.3
R8 VN.n81 VN.n53 161.3
R9 VN.n80 VN.n79 161.3
R10 VN.n78 VN.n54 161.3
R11 VN.n77 VN.n76 161.3
R12 VN.n75 VN.n55 161.3
R13 VN.n74 VN.n73 161.3
R14 VN.n72 VN.n71 161.3
R15 VN.n70 VN.n57 161.3
R16 VN.n69 VN.n68 161.3
R17 VN.n67 VN.n58 161.3
R18 VN.n66 VN.n65 161.3
R19 VN.n64 VN.n59 161.3
R20 VN.n63 VN.n62 161.3
R21 VN.n46 VN.n45 161.3
R22 VN.n44 VN.n1 161.3
R23 VN.n43 VN.n42 161.3
R24 VN.n41 VN.n2 161.3
R25 VN.n40 VN.n39 161.3
R26 VN.n38 VN.n3 161.3
R27 VN.n37 VN.n36 161.3
R28 VN.n35 VN.n34 161.3
R29 VN.n33 VN.n5 161.3
R30 VN.n32 VN.n31 161.3
R31 VN.n30 VN.n6 161.3
R32 VN.n29 VN.n28 161.3
R33 VN.n27 VN.n7 161.3
R34 VN.n26 VN.n25 161.3
R35 VN.n24 VN.n23 161.3
R36 VN.n22 VN.n9 161.3
R37 VN.n21 VN.n20 161.3
R38 VN.n19 VN.n10 161.3
R39 VN.n18 VN.n17 161.3
R40 VN.n16 VN.n11 161.3
R41 VN.n15 VN.n14 161.3
R42 VN.n47 VN.n0 75.9823
R43 VN.n95 VN.n48 75.9823
R44 VN.n61 VN.t7 72.5791
R45 VN.n13 VN.t6 72.5791
R46 VN.n13 VN.n12 61.1843
R47 VN.n61 VN.n60 61.1843
R48 VN VN.n95 51.4451
R49 VN.n43 VN.n2 43.4833
R50 VN.n91 VN.n50 43.4833
R51 VN.n17 VN.n10 41.5458
R52 VN.n32 VN.n6 41.5458
R53 VN.n65 VN.n58 41.5458
R54 VN.n80 VN.n54 41.5458
R55 VN.n21 VN.n10 39.6083
R56 VN.n28 VN.n6 39.6083
R57 VN.n69 VN.n58 39.6083
R58 VN.n76 VN.n54 39.6083
R59 VN.n12 VN.t1 39.588
R60 VN.n8 VN.t4 39.588
R61 VN.n4 VN.t0 39.588
R62 VN.n0 VN.t3 39.588
R63 VN.n60 VN.t2 39.588
R64 VN.n56 VN.t9 39.588
R65 VN.n52 VN.t5 39.588
R66 VN.n48 VN.t8 39.588
R67 VN.n39 VN.n2 37.6707
R68 VN.n87 VN.n50 37.6707
R69 VN.n16 VN.n15 24.5923
R70 VN.n17 VN.n16 24.5923
R71 VN.n22 VN.n21 24.5923
R72 VN.n23 VN.n22 24.5923
R73 VN.n27 VN.n26 24.5923
R74 VN.n28 VN.n27 24.5923
R75 VN.n33 VN.n32 24.5923
R76 VN.n34 VN.n33 24.5923
R77 VN.n38 VN.n37 24.5923
R78 VN.n39 VN.n38 24.5923
R79 VN.n44 VN.n43 24.5923
R80 VN.n45 VN.n44 24.5923
R81 VN.n65 VN.n64 24.5923
R82 VN.n64 VN.n63 24.5923
R83 VN.n76 VN.n75 24.5923
R84 VN.n75 VN.n74 24.5923
R85 VN.n71 VN.n70 24.5923
R86 VN.n70 VN.n69 24.5923
R87 VN.n87 VN.n86 24.5923
R88 VN.n86 VN.n85 24.5923
R89 VN.n82 VN.n81 24.5923
R90 VN.n81 VN.n80 24.5923
R91 VN.n93 VN.n92 24.5923
R92 VN.n92 VN.n91 24.5923
R93 VN.n45 VN.n0 14.2638
R94 VN.n93 VN.n48 14.2638
R95 VN.n15 VN.n12 13.2801
R96 VN.n34 VN.n4 13.2801
R97 VN.n63 VN.n60 13.2801
R98 VN.n82 VN.n52 13.2801
R99 VN.n23 VN.n8 12.2964
R100 VN.n26 VN.n8 12.2964
R101 VN.n74 VN.n56 12.2964
R102 VN.n71 VN.n56 12.2964
R103 VN.n37 VN.n4 11.3127
R104 VN.n85 VN.n52 11.3127
R105 VN.n62 VN.n61 4.16722
R106 VN.n14 VN.n13 4.16722
R107 VN.n95 VN.n94 0.354861
R108 VN.n47 VN.n46 0.354861
R109 VN VN.n47 0.267071
R110 VN.n94 VN.n49 0.189894
R111 VN.n90 VN.n49 0.189894
R112 VN.n90 VN.n89 0.189894
R113 VN.n89 VN.n88 0.189894
R114 VN.n88 VN.n51 0.189894
R115 VN.n84 VN.n51 0.189894
R116 VN.n84 VN.n83 0.189894
R117 VN.n83 VN.n53 0.189894
R118 VN.n79 VN.n53 0.189894
R119 VN.n79 VN.n78 0.189894
R120 VN.n78 VN.n77 0.189894
R121 VN.n77 VN.n55 0.189894
R122 VN.n73 VN.n55 0.189894
R123 VN.n73 VN.n72 0.189894
R124 VN.n72 VN.n57 0.189894
R125 VN.n68 VN.n57 0.189894
R126 VN.n68 VN.n67 0.189894
R127 VN.n67 VN.n66 0.189894
R128 VN.n66 VN.n59 0.189894
R129 VN.n62 VN.n59 0.189894
R130 VN.n14 VN.n11 0.189894
R131 VN.n18 VN.n11 0.189894
R132 VN.n19 VN.n18 0.189894
R133 VN.n20 VN.n19 0.189894
R134 VN.n20 VN.n9 0.189894
R135 VN.n24 VN.n9 0.189894
R136 VN.n25 VN.n24 0.189894
R137 VN.n25 VN.n7 0.189894
R138 VN.n29 VN.n7 0.189894
R139 VN.n30 VN.n29 0.189894
R140 VN.n31 VN.n30 0.189894
R141 VN.n31 VN.n5 0.189894
R142 VN.n35 VN.n5 0.189894
R143 VN.n36 VN.n35 0.189894
R144 VN.n36 VN.n3 0.189894
R145 VN.n40 VN.n3 0.189894
R146 VN.n41 VN.n40 0.189894
R147 VN.n42 VN.n41 0.189894
R148 VN.n42 VN.n1 0.189894
R149 VN.n46 VN.n1 0.189894
R150 VDD2.n53 VDD2.n31 289.615
R151 VDD2.n22 VDD2.n0 289.615
R152 VDD2.n54 VDD2.n53 185
R153 VDD2.n52 VDD2.n51 185
R154 VDD2.n35 VDD2.n34 185
R155 VDD2.n46 VDD2.n45 185
R156 VDD2.n44 VDD2.n43 185
R157 VDD2.n39 VDD2.n38 185
R158 VDD2.n8 VDD2.n7 185
R159 VDD2.n13 VDD2.n12 185
R160 VDD2.n15 VDD2.n14 185
R161 VDD2.n4 VDD2.n3 185
R162 VDD2.n21 VDD2.n20 185
R163 VDD2.n23 VDD2.n22 185
R164 VDD2.n40 VDD2.t2 147.672
R165 VDD2.n9 VDD2.t0 147.672
R166 VDD2.n53 VDD2.n52 104.615
R167 VDD2.n52 VDD2.n34 104.615
R168 VDD2.n45 VDD2.n34 104.615
R169 VDD2.n45 VDD2.n44 104.615
R170 VDD2.n44 VDD2.n38 104.615
R171 VDD2.n13 VDD2.n7 104.615
R172 VDD2.n14 VDD2.n13 104.615
R173 VDD2.n14 VDD2.n3 104.615
R174 VDD2.n21 VDD2.n3 104.615
R175 VDD2.n22 VDD2.n21 104.615
R176 VDD2.n30 VDD2.n29 70.0999
R177 VDD2 VDD2.n61 70.097
R178 VDD2.n60 VDD2.n59 67.8795
R179 VDD2.n28 VDD2.n27 67.8794
R180 VDD2.t2 VDD2.n38 52.3082
R181 VDD2.t0 VDD2.n7 52.3082
R182 VDD2.n28 VDD2.n26 51.1229
R183 VDD2.n58 VDD2.n57 48.0884
R184 VDD2.n58 VDD2.n30 42.6463
R185 VDD2.n40 VDD2.n39 15.6666
R186 VDD2.n9 VDD2.n8 15.6666
R187 VDD2.n43 VDD2.n42 12.8005
R188 VDD2.n12 VDD2.n11 12.8005
R189 VDD2.n46 VDD2.n37 12.0247
R190 VDD2.n15 VDD2.n6 12.0247
R191 VDD2.n47 VDD2.n35 11.249
R192 VDD2.n16 VDD2.n4 11.249
R193 VDD2.n51 VDD2.n50 10.4732
R194 VDD2.n20 VDD2.n19 10.4732
R195 VDD2.n54 VDD2.n33 9.69747
R196 VDD2.n23 VDD2.n2 9.69747
R197 VDD2.n57 VDD2.n56 9.45567
R198 VDD2.n26 VDD2.n25 9.45567
R199 VDD2.n56 VDD2.n55 9.3005
R200 VDD2.n33 VDD2.n32 9.3005
R201 VDD2.n50 VDD2.n49 9.3005
R202 VDD2.n48 VDD2.n47 9.3005
R203 VDD2.n37 VDD2.n36 9.3005
R204 VDD2.n42 VDD2.n41 9.3005
R205 VDD2.n25 VDD2.n24 9.3005
R206 VDD2.n2 VDD2.n1 9.3005
R207 VDD2.n19 VDD2.n18 9.3005
R208 VDD2.n17 VDD2.n16 9.3005
R209 VDD2.n6 VDD2.n5 9.3005
R210 VDD2.n11 VDD2.n10 9.3005
R211 VDD2.n55 VDD2.n31 8.92171
R212 VDD2.n24 VDD2.n0 8.92171
R213 VDD2.n57 VDD2.n31 5.04292
R214 VDD2.n26 VDD2.n0 5.04292
R215 VDD2.n41 VDD2.n40 4.38687
R216 VDD2.n10 VDD2.n9 4.38687
R217 VDD2.n55 VDD2.n54 4.26717
R218 VDD2.n24 VDD2.n23 4.26717
R219 VDD2.n61 VDD2.t5 3.77913
R220 VDD2.n61 VDD2.t1 3.77913
R221 VDD2.n59 VDD2.t3 3.77913
R222 VDD2.n59 VDD2.t6 3.77913
R223 VDD2.n29 VDD2.t7 3.77913
R224 VDD2.n29 VDD2.t8 3.77913
R225 VDD2.n27 VDD2.t9 3.77913
R226 VDD2.n27 VDD2.t4 3.77913
R227 VDD2.n51 VDD2.n33 3.49141
R228 VDD2.n20 VDD2.n2 3.49141
R229 VDD2.n60 VDD2.n58 3.03498
R230 VDD2.n50 VDD2.n35 2.71565
R231 VDD2.n19 VDD2.n4 2.71565
R232 VDD2.n47 VDD2.n46 1.93989
R233 VDD2.n16 VDD2.n15 1.93989
R234 VDD2.n43 VDD2.n37 1.16414
R235 VDD2.n12 VDD2.n6 1.16414
R236 VDD2 VDD2.n60 0.81731
R237 VDD2.n30 VDD2.n28 0.703775
R238 VDD2.n42 VDD2.n39 0.388379
R239 VDD2.n11 VDD2.n8 0.388379
R240 VDD2.n56 VDD2.n32 0.155672
R241 VDD2.n49 VDD2.n32 0.155672
R242 VDD2.n49 VDD2.n48 0.155672
R243 VDD2.n48 VDD2.n36 0.155672
R244 VDD2.n41 VDD2.n36 0.155672
R245 VDD2.n10 VDD2.n5 0.155672
R246 VDD2.n17 VDD2.n5 0.155672
R247 VDD2.n18 VDD2.n17 0.155672
R248 VDD2.n18 VDD2.n1 0.155672
R249 VDD2.n25 VDD2.n1 0.155672
R250 VTAIL.n120 VTAIL.n98 289.615
R251 VTAIL.n24 VTAIL.n2 289.615
R252 VTAIL.n92 VTAIL.n70 289.615
R253 VTAIL.n60 VTAIL.n38 289.615
R254 VTAIL.n106 VTAIL.n105 185
R255 VTAIL.n111 VTAIL.n110 185
R256 VTAIL.n113 VTAIL.n112 185
R257 VTAIL.n102 VTAIL.n101 185
R258 VTAIL.n119 VTAIL.n118 185
R259 VTAIL.n121 VTAIL.n120 185
R260 VTAIL.n10 VTAIL.n9 185
R261 VTAIL.n15 VTAIL.n14 185
R262 VTAIL.n17 VTAIL.n16 185
R263 VTAIL.n6 VTAIL.n5 185
R264 VTAIL.n23 VTAIL.n22 185
R265 VTAIL.n25 VTAIL.n24 185
R266 VTAIL.n93 VTAIL.n92 185
R267 VTAIL.n91 VTAIL.n90 185
R268 VTAIL.n74 VTAIL.n73 185
R269 VTAIL.n85 VTAIL.n84 185
R270 VTAIL.n83 VTAIL.n82 185
R271 VTAIL.n78 VTAIL.n77 185
R272 VTAIL.n61 VTAIL.n60 185
R273 VTAIL.n59 VTAIL.n58 185
R274 VTAIL.n42 VTAIL.n41 185
R275 VTAIL.n53 VTAIL.n52 185
R276 VTAIL.n51 VTAIL.n50 185
R277 VTAIL.n46 VTAIL.n45 185
R278 VTAIL.n107 VTAIL.t16 147.672
R279 VTAIL.n11 VTAIL.t8 147.672
R280 VTAIL.n79 VTAIL.t3 147.672
R281 VTAIL.n47 VTAIL.t12 147.672
R282 VTAIL.n111 VTAIL.n105 104.615
R283 VTAIL.n112 VTAIL.n111 104.615
R284 VTAIL.n112 VTAIL.n101 104.615
R285 VTAIL.n119 VTAIL.n101 104.615
R286 VTAIL.n120 VTAIL.n119 104.615
R287 VTAIL.n15 VTAIL.n9 104.615
R288 VTAIL.n16 VTAIL.n15 104.615
R289 VTAIL.n16 VTAIL.n5 104.615
R290 VTAIL.n23 VTAIL.n5 104.615
R291 VTAIL.n24 VTAIL.n23 104.615
R292 VTAIL.n92 VTAIL.n91 104.615
R293 VTAIL.n91 VTAIL.n73 104.615
R294 VTAIL.n84 VTAIL.n73 104.615
R295 VTAIL.n84 VTAIL.n83 104.615
R296 VTAIL.n83 VTAIL.n77 104.615
R297 VTAIL.n60 VTAIL.n59 104.615
R298 VTAIL.n59 VTAIL.n41 104.615
R299 VTAIL.n52 VTAIL.n41 104.615
R300 VTAIL.n52 VTAIL.n51 104.615
R301 VTAIL.n51 VTAIL.n45 104.615
R302 VTAIL.t16 VTAIL.n105 52.3082
R303 VTAIL.t8 VTAIL.n9 52.3082
R304 VTAIL.t3 VTAIL.n77 52.3082
R305 VTAIL.t12 VTAIL.n45 52.3082
R306 VTAIL.n69 VTAIL.n68 51.2007
R307 VTAIL.n67 VTAIL.n66 51.2007
R308 VTAIL.n37 VTAIL.n36 51.2007
R309 VTAIL.n35 VTAIL.n34 51.2007
R310 VTAIL.n127 VTAIL.n126 51.2006
R311 VTAIL.n1 VTAIL.n0 51.2006
R312 VTAIL.n31 VTAIL.n30 51.2006
R313 VTAIL.n33 VTAIL.n32 51.2006
R314 VTAIL.n125 VTAIL.n124 31.4096
R315 VTAIL.n29 VTAIL.n28 31.4096
R316 VTAIL.n97 VTAIL.n96 31.4096
R317 VTAIL.n65 VTAIL.n64 31.4096
R318 VTAIL.n35 VTAIL.n33 22.9531
R319 VTAIL.n125 VTAIL.n97 19.9186
R320 VTAIL.n107 VTAIL.n106 15.6666
R321 VTAIL.n11 VTAIL.n10 15.6666
R322 VTAIL.n79 VTAIL.n78 15.6666
R323 VTAIL.n47 VTAIL.n46 15.6666
R324 VTAIL.n110 VTAIL.n109 12.8005
R325 VTAIL.n14 VTAIL.n13 12.8005
R326 VTAIL.n82 VTAIL.n81 12.8005
R327 VTAIL.n50 VTAIL.n49 12.8005
R328 VTAIL.n113 VTAIL.n104 12.0247
R329 VTAIL.n17 VTAIL.n8 12.0247
R330 VTAIL.n85 VTAIL.n76 12.0247
R331 VTAIL.n53 VTAIL.n44 12.0247
R332 VTAIL.n114 VTAIL.n102 11.249
R333 VTAIL.n18 VTAIL.n6 11.249
R334 VTAIL.n86 VTAIL.n74 11.249
R335 VTAIL.n54 VTAIL.n42 11.249
R336 VTAIL.n118 VTAIL.n117 10.4732
R337 VTAIL.n22 VTAIL.n21 10.4732
R338 VTAIL.n90 VTAIL.n89 10.4732
R339 VTAIL.n58 VTAIL.n57 10.4732
R340 VTAIL.n121 VTAIL.n100 9.69747
R341 VTAIL.n25 VTAIL.n4 9.69747
R342 VTAIL.n93 VTAIL.n72 9.69747
R343 VTAIL.n61 VTAIL.n40 9.69747
R344 VTAIL.n124 VTAIL.n123 9.45567
R345 VTAIL.n28 VTAIL.n27 9.45567
R346 VTAIL.n96 VTAIL.n95 9.45567
R347 VTAIL.n64 VTAIL.n63 9.45567
R348 VTAIL.n123 VTAIL.n122 9.3005
R349 VTAIL.n100 VTAIL.n99 9.3005
R350 VTAIL.n117 VTAIL.n116 9.3005
R351 VTAIL.n115 VTAIL.n114 9.3005
R352 VTAIL.n104 VTAIL.n103 9.3005
R353 VTAIL.n109 VTAIL.n108 9.3005
R354 VTAIL.n27 VTAIL.n26 9.3005
R355 VTAIL.n4 VTAIL.n3 9.3005
R356 VTAIL.n21 VTAIL.n20 9.3005
R357 VTAIL.n19 VTAIL.n18 9.3005
R358 VTAIL.n8 VTAIL.n7 9.3005
R359 VTAIL.n13 VTAIL.n12 9.3005
R360 VTAIL.n95 VTAIL.n94 9.3005
R361 VTAIL.n72 VTAIL.n71 9.3005
R362 VTAIL.n89 VTAIL.n88 9.3005
R363 VTAIL.n87 VTAIL.n86 9.3005
R364 VTAIL.n76 VTAIL.n75 9.3005
R365 VTAIL.n81 VTAIL.n80 9.3005
R366 VTAIL.n63 VTAIL.n62 9.3005
R367 VTAIL.n40 VTAIL.n39 9.3005
R368 VTAIL.n57 VTAIL.n56 9.3005
R369 VTAIL.n55 VTAIL.n54 9.3005
R370 VTAIL.n44 VTAIL.n43 9.3005
R371 VTAIL.n49 VTAIL.n48 9.3005
R372 VTAIL.n122 VTAIL.n98 8.92171
R373 VTAIL.n26 VTAIL.n2 8.92171
R374 VTAIL.n94 VTAIL.n70 8.92171
R375 VTAIL.n62 VTAIL.n38 8.92171
R376 VTAIL.n124 VTAIL.n98 5.04292
R377 VTAIL.n28 VTAIL.n2 5.04292
R378 VTAIL.n96 VTAIL.n70 5.04292
R379 VTAIL.n64 VTAIL.n38 5.04292
R380 VTAIL.n108 VTAIL.n107 4.38687
R381 VTAIL.n12 VTAIL.n11 4.38687
R382 VTAIL.n80 VTAIL.n79 4.38687
R383 VTAIL.n48 VTAIL.n47 4.38687
R384 VTAIL.n122 VTAIL.n121 4.26717
R385 VTAIL.n26 VTAIL.n25 4.26717
R386 VTAIL.n94 VTAIL.n93 4.26717
R387 VTAIL.n62 VTAIL.n61 4.26717
R388 VTAIL.n126 VTAIL.t15 3.77913
R389 VTAIL.n126 VTAIL.t19 3.77913
R390 VTAIL.n0 VTAIL.t13 3.77913
R391 VTAIL.n0 VTAIL.t18 3.77913
R392 VTAIL.n30 VTAIL.t5 3.77913
R393 VTAIL.n30 VTAIL.t6 3.77913
R394 VTAIL.n32 VTAIL.t4 3.77913
R395 VTAIL.n32 VTAIL.t0 3.77913
R396 VTAIL.n68 VTAIL.t1 3.77913
R397 VTAIL.n68 VTAIL.t7 3.77913
R398 VTAIL.n66 VTAIL.t2 3.77913
R399 VTAIL.n66 VTAIL.t9 3.77913
R400 VTAIL.n36 VTAIL.t10 3.77913
R401 VTAIL.n36 VTAIL.t17 3.77913
R402 VTAIL.n34 VTAIL.t11 3.77913
R403 VTAIL.n34 VTAIL.t14 3.77913
R404 VTAIL.n118 VTAIL.n100 3.49141
R405 VTAIL.n22 VTAIL.n4 3.49141
R406 VTAIL.n90 VTAIL.n72 3.49141
R407 VTAIL.n58 VTAIL.n40 3.49141
R408 VTAIL.n37 VTAIL.n35 3.03498
R409 VTAIL.n65 VTAIL.n37 3.03498
R410 VTAIL.n69 VTAIL.n67 3.03498
R411 VTAIL.n97 VTAIL.n69 3.03498
R412 VTAIL.n33 VTAIL.n31 3.03498
R413 VTAIL.n31 VTAIL.n29 3.03498
R414 VTAIL.n127 VTAIL.n125 3.03498
R415 VTAIL.n117 VTAIL.n102 2.71565
R416 VTAIL.n21 VTAIL.n6 2.71565
R417 VTAIL.n89 VTAIL.n74 2.71565
R418 VTAIL.n57 VTAIL.n42 2.71565
R419 VTAIL VTAIL.n1 2.33455
R420 VTAIL.n67 VTAIL.n65 1.98757
R421 VTAIL.n29 VTAIL.n1 1.98757
R422 VTAIL.n114 VTAIL.n113 1.93989
R423 VTAIL.n18 VTAIL.n17 1.93989
R424 VTAIL.n86 VTAIL.n85 1.93989
R425 VTAIL.n54 VTAIL.n53 1.93989
R426 VTAIL.n110 VTAIL.n104 1.16414
R427 VTAIL.n14 VTAIL.n8 1.16414
R428 VTAIL.n82 VTAIL.n76 1.16414
R429 VTAIL.n50 VTAIL.n44 1.16414
R430 VTAIL VTAIL.n127 0.700931
R431 VTAIL.n109 VTAIL.n106 0.388379
R432 VTAIL.n13 VTAIL.n10 0.388379
R433 VTAIL.n81 VTAIL.n78 0.388379
R434 VTAIL.n49 VTAIL.n46 0.388379
R435 VTAIL.n108 VTAIL.n103 0.155672
R436 VTAIL.n115 VTAIL.n103 0.155672
R437 VTAIL.n116 VTAIL.n115 0.155672
R438 VTAIL.n116 VTAIL.n99 0.155672
R439 VTAIL.n123 VTAIL.n99 0.155672
R440 VTAIL.n12 VTAIL.n7 0.155672
R441 VTAIL.n19 VTAIL.n7 0.155672
R442 VTAIL.n20 VTAIL.n19 0.155672
R443 VTAIL.n20 VTAIL.n3 0.155672
R444 VTAIL.n27 VTAIL.n3 0.155672
R445 VTAIL.n95 VTAIL.n71 0.155672
R446 VTAIL.n88 VTAIL.n71 0.155672
R447 VTAIL.n88 VTAIL.n87 0.155672
R448 VTAIL.n87 VTAIL.n75 0.155672
R449 VTAIL.n80 VTAIL.n75 0.155672
R450 VTAIL.n63 VTAIL.n39 0.155672
R451 VTAIL.n56 VTAIL.n39 0.155672
R452 VTAIL.n56 VTAIL.n55 0.155672
R453 VTAIL.n55 VTAIL.n43 0.155672
R454 VTAIL.n48 VTAIL.n43 0.155672
R455 B.n734 B.n733 585
R456 B.n734 B.n127 585
R457 B.n737 B.n736 585
R458 B.n738 B.n158 585
R459 B.n740 B.n739 585
R460 B.n742 B.n157 585
R461 B.n745 B.n744 585
R462 B.n746 B.n156 585
R463 B.n748 B.n747 585
R464 B.n750 B.n155 585
R465 B.n753 B.n752 585
R466 B.n754 B.n154 585
R467 B.n756 B.n755 585
R468 B.n758 B.n153 585
R469 B.n761 B.n760 585
R470 B.n762 B.n152 585
R471 B.n764 B.n763 585
R472 B.n766 B.n151 585
R473 B.n769 B.n768 585
R474 B.n770 B.n150 585
R475 B.n772 B.n771 585
R476 B.n774 B.n149 585
R477 B.n777 B.n776 585
R478 B.n779 B.n146 585
R479 B.n781 B.n780 585
R480 B.n783 B.n145 585
R481 B.n786 B.n785 585
R482 B.n787 B.n144 585
R483 B.n789 B.n788 585
R484 B.n791 B.n143 585
R485 B.n793 B.n792 585
R486 B.n795 B.n794 585
R487 B.n798 B.n797 585
R488 B.n799 B.n138 585
R489 B.n801 B.n800 585
R490 B.n803 B.n137 585
R491 B.n806 B.n805 585
R492 B.n807 B.n136 585
R493 B.n809 B.n808 585
R494 B.n811 B.n135 585
R495 B.n814 B.n813 585
R496 B.n815 B.n134 585
R497 B.n817 B.n816 585
R498 B.n819 B.n133 585
R499 B.n822 B.n821 585
R500 B.n823 B.n132 585
R501 B.n825 B.n824 585
R502 B.n827 B.n131 585
R503 B.n830 B.n829 585
R504 B.n831 B.n130 585
R505 B.n833 B.n832 585
R506 B.n835 B.n129 585
R507 B.n838 B.n837 585
R508 B.n839 B.n128 585
R509 B.n732 B.n126 585
R510 B.n842 B.n126 585
R511 B.n731 B.n125 585
R512 B.n843 B.n125 585
R513 B.n730 B.n124 585
R514 B.n844 B.n124 585
R515 B.n729 B.n728 585
R516 B.n728 B.n120 585
R517 B.n727 B.n119 585
R518 B.n850 B.n119 585
R519 B.n726 B.n118 585
R520 B.n851 B.n118 585
R521 B.n725 B.n117 585
R522 B.n852 B.n117 585
R523 B.n724 B.n723 585
R524 B.n723 B.n113 585
R525 B.n722 B.n112 585
R526 B.n858 B.n112 585
R527 B.n721 B.n111 585
R528 B.n859 B.n111 585
R529 B.n720 B.n110 585
R530 B.n860 B.n110 585
R531 B.n719 B.n718 585
R532 B.n718 B.n106 585
R533 B.n717 B.n105 585
R534 B.n866 B.n105 585
R535 B.n716 B.n104 585
R536 B.n867 B.n104 585
R537 B.n715 B.n103 585
R538 B.n868 B.n103 585
R539 B.n714 B.n713 585
R540 B.n713 B.n99 585
R541 B.n712 B.n98 585
R542 B.n874 B.n98 585
R543 B.n711 B.n97 585
R544 B.n875 B.n97 585
R545 B.n710 B.n96 585
R546 B.n876 B.n96 585
R547 B.n709 B.n708 585
R548 B.n708 B.n92 585
R549 B.n707 B.n91 585
R550 B.n882 B.n91 585
R551 B.n706 B.n90 585
R552 B.n883 B.n90 585
R553 B.n705 B.n89 585
R554 B.n884 B.n89 585
R555 B.n704 B.n703 585
R556 B.n703 B.n85 585
R557 B.n702 B.n84 585
R558 B.n890 B.n84 585
R559 B.n701 B.n83 585
R560 B.n891 B.n83 585
R561 B.n700 B.n82 585
R562 B.n892 B.n82 585
R563 B.n699 B.n698 585
R564 B.n698 B.n78 585
R565 B.n697 B.n77 585
R566 B.n898 B.n77 585
R567 B.n696 B.n76 585
R568 B.n899 B.n76 585
R569 B.n695 B.n75 585
R570 B.n900 B.n75 585
R571 B.n694 B.n693 585
R572 B.n693 B.n71 585
R573 B.n692 B.n70 585
R574 B.n906 B.n70 585
R575 B.n691 B.n69 585
R576 B.n907 B.n69 585
R577 B.n690 B.n68 585
R578 B.n908 B.n68 585
R579 B.n689 B.n688 585
R580 B.n688 B.n64 585
R581 B.n687 B.n63 585
R582 B.n914 B.n63 585
R583 B.n686 B.n62 585
R584 B.n915 B.n62 585
R585 B.n685 B.n61 585
R586 B.n916 B.n61 585
R587 B.n684 B.n683 585
R588 B.n683 B.n57 585
R589 B.n682 B.n56 585
R590 B.n922 B.n56 585
R591 B.n681 B.n55 585
R592 B.n923 B.n55 585
R593 B.n680 B.n54 585
R594 B.n924 B.n54 585
R595 B.n679 B.n678 585
R596 B.n678 B.n50 585
R597 B.n677 B.n49 585
R598 B.n930 B.n49 585
R599 B.n676 B.n48 585
R600 B.n931 B.n48 585
R601 B.n675 B.n47 585
R602 B.n932 B.n47 585
R603 B.n674 B.n673 585
R604 B.n673 B.n43 585
R605 B.n672 B.n42 585
R606 B.n938 B.n42 585
R607 B.n671 B.n41 585
R608 B.n939 B.n41 585
R609 B.n670 B.n40 585
R610 B.n940 B.n40 585
R611 B.n669 B.n668 585
R612 B.n668 B.n36 585
R613 B.n667 B.n35 585
R614 B.n946 B.n35 585
R615 B.n666 B.n34 585
R616 B.n947 B.n34 585
R617 B.n665 B.n33 585
R618 B.n948 B.n33 585
R619 B.n664 B.n663 585
R620 B.n663 B.n29 585
R621 B.n662 B.n28 585
R622 B.n954 B.n28 585
R623 B.n661 B.n27 585
R624 B.n955 B.n27 585
R625 B.n660 B.n26 585
R626 B.n956 B.n26 585
R627 B.n659 B.n658 585
R628 B.n658 B.n22 585
R629 B.n657 B.n21 585
R630 B.n962 B.n21 585
R631 B.n656 B.n20 585
R632 B.n963 B.n20 585
R633 B.n655 B.n19 585
R634 B.n964 B.n19 585
R635 B.n654 B.n653 585
R636 B.n653 B.n18 585
R637 B.n652 B.n14 585
R638 B.n970 B.n14 585
R639 B.n651 B.n13 585
R640 B.n971 B.n13 585
R641 B.n650 B.n12 585
R642 B.n972 B.n12 585
R643 B.n649 B.n648 585
R644 B.n648 B.n8 585
R645 B.n647 B.n7 585
R646 B.n978 B.n7 585
R647 B.n646 B.n6 585
R648 B.n979 B.n6 585
R649 B.n645 B.n5 585
R650 B.n980 B.n5 585
R651 B.n644 B.n643 585
R652 B.n643 B.n4 585
R653 B.n642 B.n159 585
R654 B.n642 B.n641 585
R655 B.n632 B.n160 585
R656 B.n161 B.n160 585
R657 B.n634 B.n633 585
R658 B.n635 B.n634 585
R659 B.n631 B.n166 585
R660 B.n166 B.n165 585
R661 B.n630 B.n629 585
R662 B.n629 B.n628 585
R663 B.n168 B.n167 585
R664 B.n621 B.n168 585
R665 B.n620 B.n619 585
R666 B.n622 B.n620 585
R667 B.n618 B.n173 585
R668 B.n173 B.n172 585
R669 B.n617 B.n616 585
R670 B.n616 B.n615 585
R671 B.n175 B.n174 585
R672 B.n176 B.n175 585
R673 B.n608 B.n607 585
R674 B.n609 B.n608 585
R675 B.n606 B.n181 585
R676 B.n181 B.n180 585
R677 B.n605 B.n604 585
R678 B.n604 B.n603 585
R679 B.n183 B.n182 585
R680 B.n184 B.n183 585
R681 B.n596 B.n595 585
R682 B.n597 B.n596 585
R683 B.n594 B.n189 585
R684 B.n189 B.n188 585
R685 B.n593 B.n592 585
R686 B.n592 B.n591 585
R687 B.n191 B.n190 585
R688 B.n192 B.n191 585
R689 B.n584 B.n583 585
R690 B.n585 B.n584 585
R691 B.n582 B.n197 585
R692 B.n197 B.n196 585
R693 B.n581 B.n580 585
R694 B.n580 B.n579 585
R695 B.n199 B.n198 585
R696 B.n200 B.n199 585
R697 B.n572 B.n571 585
R698 B.n573 B.n572 585
R699 B.n570 B.n205 585
R700 B.n205 B.n204 585
R701 B.n569 B.n568 585
R702 B.n568 B.n567 585
R703 B.n207 B.n206 585
R704 B.n208 B.n207 585
R705 B.n560 B.n559 585
R706 B.n561 B.n560 585
R707 B.n558 B.n213 585
R708 B.n213 B.n212 585
R709 B.n557 B.n556 585
R710 B.n556 B.n555 585
R711 B.n215 B.n214 585
R712 B.n216 B.n215 585
R713 B.n548 B.n547 585
R714 B.n549 B.n548 585
R715 B.n546 B.n221 585
R716 B.n221 B.n220 585
R717 B.n545 B.n544 585
R718 B.n544 B.n543 585
R719 B.n223 B.n222 585
R720 B.n224 B.n223 585
R721 B.n536 B.n535 585
R722 B.n537 B.n536 585
R723 B.n534 B.n229 585
R724 B.n229 B.n228 585
R725 B.n533 B.n532 585
R726 B.n532 B.n531 585
R727 B.n231 B.n230 585
R728 B.n232 B.n231 585
R729 B.n524 B.n523 585
R730 B.n525 B.n524 585
R731 B.n522 B.n237 585
R732 B.n237 B.n236 585
R733 B.n521 B.n520 585
R734 B.n520 B.n519 585
R735 B.n239 B.n238 585
R736 B.n240 B.n239 585
R737 B.n512 B.n511 585
R738 B.n513 B.n512 585
R739 B.n510 B.n245 585
R740 B.n245 B.n244 585
R741 B.n509 B.n508 585
R742 B.n508 B.n507 585
R743 B.n247 B.n246 585
R744 B.n248 B.n247 585
R745 B.n500 B.n499 585
R746 B.n501 B.n500 585
R747 B.n498 B.n252 585
R748 B.n256 B.n252 585
R749 B.n497 B.n496 585
R750 B.n496 B.n495 585
R751 B.n254 B.n253 585
R752 B.n255 B.n254 585
R753 B.n488 B.n487 585
R754 B.n489 B.n488 585
R755 B.n486 B.n261 585
R756 B.n261 B.n260 585
R757 B.n485 B.n484 585
R758 B.n484 B.n483 585
R759 B.n263 B.n262 585
R760 B.n264 B.n263 585
R761 B.n476 B.n475 585
R762 B.n477 B.n476 585
R763 B.n474 B.n269 585
R764 B.n269 B.n268 585
R765 B.n473 B.n472 585
R766 B.n472 B.n471 585
R767 B.n271 B.n270 585
R768 B.n272 B.n271 585
R769 B.n464 B.n463 585
R770 B.n465 B.n464 585
R771 B.n462 B.n277 585
R772 B.n277 B.n276 585
R773 B.n461 B.n460 585
R774 B.n460 B.n459 585
R775 B.n279 B.n278 585
R776 B.n280 B.n279 585
R777 B.n452 B.n451 585
R778 B.n453 B.n452 585
R779 B.n450 B.n285 585
R780 B.n285 B.n284 585
R781 B.n449 B.n448 585
R782 B.n448 B.n447 585
R783 B.n287 B.n286 585
R784 B.n288 B.n287 585
R785 B.n440 B.n439 585
R786 B.n441 B.n440 585
R787 B.n438 B.n293 585
R788 B.n293 B.n292 585
R789 B.n437 B.n436 585
R790 B.n436 B.n435 585
R791 B.n432 B.n297 585
R792 B.n431 B.n430 585
R793 B.n428 B.n298 585
R794 B.n428 B.n296 585
R795 B.n427 B.n426 585
R796 B.n425 B.n424 585
R797 B.n423 B.n300 585
R798 B.n421 B.n420 585
R799 B.n419 B.n301 585
R800 B.n418 B.n417 585
R801 B.n415 B.n302 585
R802 B.n413 B.n412 585
R803 B.n411 B.n303 585
R804 B.n410 B.n409 585
R805 B.n407 B.n304 585
R806 B.n405 B.n404 585
R807 B.n403 B.n305 585
R808 B.n402 B.n401 585
R809 B.n399 B.n306 585
R810 B.n397 B.n396 585
R811 B.n395 B.n307 585
R812 B.n394 B.n393 585
R813 B.n391 B.n308 585
R814 B.n389 B.n388 585
R815 B.n387 B.n309 585
R816 B.n386 B.n385 585
R817 B.n383 B.n313 585
R818 B.n381 B.n380 585
R819 B.n379 B.n314 585
R820 B.n378 B.n377 585
R821 B.n375 B.n315 585
R822 B.n373 B.n372 585
R823 B.n370 B.n316 585
R824 B.n369 B.n368 585
R825 B.n366 B.n319 585
R826 B.n364 B.n363 585
R827 B.n362 B.n320 585
R828 B.n361 B.n360 585
R829 B.n358 B.n321 585
R830 B.n356 B.n355 585
R831 B.n354 B.n322 585
R832 B.n353 B.n352 585
R833 B.n350 B.n323 585
R834 B.n348 B.n347 585
R835 B.n346 B.n324 585
R836 B.n345 B.n344 585
R837 B.n342 B.n325 585
R838 B.n340 B.n339 585
R839 B.n338 B.n326 585
R840 B.n337 B.n336 585
R841 B.n334 B.n327 585
R842 B.n332 B.n331 585
R843 B.n330 B.n329 585
R844 B.n295 B.n294 585
R845 B.n434 B.n433 585
R846 B.n435 B.n434 585
R847 B.n291 B.n290 585
R848 B.n292 B.n291 585
R849 B.n443 B.n442 585
R850 B.n442 B.n441 585
R851 B.n444 B.n289 585
R852 B.n289 B.n288 585
R853 B.n446 B.n445 585
R854 B.n447 B.n446 585
R855 B.n283 B.n282 585
R856 B.n284 B.n283 585
R857 B.n455 B.n454 585
R858 B.n454 B.n453 585
R859 B.n456 B.n281 585
R860 B.n281 B.n280 585
R861 B.n458 B.n457 585
R862 B.n459 B.n458 585
R863 B.n275 B.n274 585
R864 B.n276 B.n275 585
R865 B.n467 B.n466 585
R866 B.n466 B.n465 585
R867 B.n468 B.n273 585
R868 B.n273 B.n272 585
R869 B.n470 B.n469 585
R870 B.n471 B.n470 585
R871 B.n267 B.n266 585
R872 B.n268 B.n267 585
R873 B.n479 B.n478 585
R874 B.n478 B.n477 585
R875 B.n480 B.n265 585
R876 B.n265 B.n264 585
R877 B.n482 B.n481 585
R878 B.n483 B.n482 585
R879 B.n259 B.n258 585
R880 B.n260 B.n259 585
R881 B.n491 B.n490 585
R882 B.n490 B.n489 585
R883 B.n492 B.n257 585
R884 B.n257 B.n255 585
R885 B.n494 B.n493 585
R886 B.n495 B.n494 585
R887 B.n251 B.n250 585
R888 B.n256 B.n251 585
R889 B.n503 B.n502 585
R890 B.n502 B.n501 585
R891 B.n504 B.n249 585
R892 B.n249 B.n248 585
R893 B.n506 B.n505 585
R894 B.n507 B.n506 585
R895 B.n243 B.n242 585
R896 B.n244 B.n243 585
R897 B.n515 B.n514 585
R898 B.n514 B.n513 585
R899 B.n516 B.n241 585
R900 B.n241 B.n240 585
R901 B.n518 B.n517 585
R902 B.n519 B.n518 585
R903 B.n235 B.n234 585
R904 B.n236 B.n235 585
R905 B.n527 B.n526 585
R906 B.n526 B.n525 585
R907 B.n528 B.n233 585
R908 B.n233 B.n232 585
R909 B.n530 B.n529 585
R910 B.n531 B.n530 585
R911 B.n227 B.n226 585
R912 B.n228 B.n227 585
R913 B.n539 B.n538 585
R914 B.n538 B.n537 585
R915 B.n540 B.n225 585
R916 B.n225 B.n224 585
R917 B.n542 B.n541 585
R918 B.n543 B.n542 585
R919 B.n219 B.n218 585
R920 B.n220 B.n219 585
R921 B.n551 B.n550 585
R922 B.n550 B.n549 585
R923 B.n552 B.n217 585
R924 B.n217 B.n216 585
R925 B.n554 B.n553 585
R926 B.n555 B.n554 585
R927 B.n211 B.n210 585
R928 B.n212 B.n211 585
R929 B.n563 B.n562 585
R930 B.n562 B.n561 585
R931 B.n564 B.n209 585
R932 B.n209 B.n208 585
R933 B.n566 B.n565 585
R934 B.n567 B.n566 585
R935 B.n203 B.n202 585
R936 B.n204 B.n203 585
R937 B.n575 B.n574 585
R938 B.n574 B.n573 585
R939 B.n576 B.n201 585
R940 B.n201 B.n200 585
R941 B.n578 B.n577 585
R942 B.n579 B.n578 585
R943 B.n195 B.n194 585
R944 B.n196 B.n195 585
R945 B.n587 B.n586 585
R946 B.n586 B.n585 585
R947 B.n588 B.n193 585
R948 B.n193 B.n192 585
R949 B.n590 B.n589 585
R950 B.n591 B.n590 585
R951 B.n187 B.n186 585
R952 B.n188 B.n187 585
R953 B.n599 B.n598 585
R954 B.n598 B.n597 585
R955 B.n600 B.n185 585
R956 B.n185 B.n184 585
R957 B.n602 B.n601 585
R958 B.n603 B.n602 585
R959 B.n179 B.n178 585
R960 B.n180 B.n179 585
R961 B.n611 B.n610 585
R962 B.n610 B.n609 585
R963 B.n612 B.n177 585
R964 B.n177 B.n176 585
R965 B.n614 B.n613 585
R966 B.n615 B.n614 585
R967 B.n171 B.n170 585
R968 B.n172 B.n171 585
R969 B.n624 B.n623 585
R970 B.n623 B.n622 585
R971 B.n625 B.n169 585
R972 B.n621 B.n169 585
R973 B.n627 B.n626 585
R974 B.n628 B.n627 585
R975 B.n164 B.n163 585
R976 B.n165 B.n164 585
R977 B.n637 B.n636 585
R978 B.n636 B.n635 585
R979 B.n638 B.n162 585
R980 B.n162 B.n161 585
R981 B.n640 B.n639 585
R982 B.n641 B.n640 585
R983 B.n2 B.n0 585
R984 B.n4 B.n2 585
R985 B.n3 B.n1 585
R986 B.n979 B.n3 585
R987 B.n977 B.n976 585
R988 B.n978 B.n977 585
R989 B.n975 B.n9 585
R990 B.n9 B.n8 585
R991 B.n974 B.n973 585
R992 B.n973 B.n972 585
R993 B.n11 B.n10 585
R994 B.n971 B.n11 585
R995 B.n969 B.n968 585
R996 B.n970 B.n969 585
R997 B.n967 B.n15 585
R998 B.n18 B.n15 585
R999 B.n966 B.n965 585
R1000 B.n965 B.n964 585
R1001 B.n17 B.n16 585
R1002 B.n963 B.n17 585
R1003 B.n961 B.n960 585
R1004 B.n962 B.n961 585
R1005 B.n959 B.n23 585
R1006 B.n23 B.n22 585
R1007 B.n958 B.n957 585
R1008 B.n957 B.n956 585
R1009 B.n25 B.n24 585
R1010 B.n955 B.n25 585
R1011 B.n953 B.n952 585
R1012 B.n954 B.n953 585
R1013 B.n951 B.n30 585
R1014 B.n30 B.n29 585
R1015 B.n950 B.n949 585
R1016 B.n949 B.n948 585
R1017 B.n32 B.n31 585
R1018 B.n947 B.n32 585
R1019 B.n945 B.n944 585
R1020 B.n946 B.n945 585
R1021 B.n943 B.n37 585
R1022 B.n37 B.n36 585
R1023 B.n942 B.n941 585
R1024 B.n941 B.n940 585
R1025 B.n39 B.n38 585
R1026 B.n939 B.n39 585
R1027 B.n937 B.n936 585
R1028 B.n938 B.n937 585
R1029 B.n935 B.n44 585
R1030 B.n44 B.n43 585
R1031 B.n934 B.n933 585
R1032 B.n933 B.n932 585
R1033 B.n46 B.n45 585
R1034 B.n931 B.n46 585
R1035 B.n929 B.n928 585
R1036 B.n930 B.n929 585
R1037 B.n927 B.n51 585
R1038 B.n51 B.n50 585
R1039 B.n926 B.n925 585
R1040 B.n925 B.n924 585
R1041 B.n53 B.n52 585
R1042 B.n923 B.n53 585
R1043 B.n921 B.n920 585
R1044 B.n922 B.n921 585
R1045 B.n919 B.n58 585
R1046 B.n58 B.n57 585
R1047 B.n918 B.n917 585
R1048 B.n917 B.n916 585
R1049 B.n60 B.n59 585
R1050 B.n915 B.n60 585
R1051 B.n913 B.n912 585
R1052 B.n914 B.n913 585
R1053 B.n911 B.n65 585
R1054 B.n65 B.n64 585
R1055 B.n910 B.n909 585
R1056 B.n909 B.n908 585
R1057 B.n67 B.n66 585
R1058 B.n907 B.n67 585
R1059 B.n905 B.n904 585
R1060 B.n906 B.n905 585
R1061 B.n903 B.n72 585
R1062 B.n72 B.n71 585
R1063 B.n902 B.n901 585
R1064 B.n901 B.n900 585
R1065 B.n74 B.n73 585
R1066 B.n899 B.n74 585
R1067 B.n897 B.n896 585
R1068 B.n898 B.n897 585
R1069 B.n895 B.n79 585
R1070 B.n79 B.n78 585
R1071 B.n894 B.n893 585
R1072 B.n893 B.n892 585
R1073 B.n81 B.n80 585
R1074 B.n891 B.n81 585
R1075 B.n889 B.n888 585
R1076 B.n890 B.n889 585
R1077 B.n887 B.n86 585
R1078 B.n86 B.n85 585
R1079 B.n886 B.n885 585
R1080 B.n885 B.n884 585
R1081 B.n88 B.n87 585
R1082 B.n883 B.n88 585
R1083 B.n881 B.n880 585
R1084 B.n882 B.n881 585
R1085 B.n879 B.n93 585
R1086 B.n93 B.n92 585
R1087 B.n878 B.n877 585
R1088 B.n877 B.n876 585
R1089 B.n95 B.n94 585
R1090 B.n875 B.n95 585
R1091 B.n873 B.n872 585
R1092 B.n874 B.n873 585
R1093 B.n871 B.n100 585
R1094 B.n100 B.n99 585
R1095 B.n870 B.n869 585
R1096 B.n869 B.n868 585
R1097 B.n102 B.n101 585
R1098 B.n867 B.n102 585
R1099 B.n865 B.n864 585
R1100 B.n866 B.n865 585
R1101 B.n863 B.n107 585
R1102 B.n107 B.n106 585
R1103 B.n862 B.n861 585
R1104 B.n861 B.n860 585
R1105 B.n109 B.n108 585
R1106 B.n859 B.n109 585
R1107 B.n857 B.n856 585
R1108 B.n858 B.n857 585
R1109 B.n855 B.n114 585
R1110 B.n114 B.n113 585
R1111 B.n854 B.n853 585
R1112 B.n853 B.n852 585
R1113 B.n116 B.n115 585
R1114 B.n851 B.n116 585
R1115 B.n849 B.n848 585
R1116 B.n850 B.n849 585
R1117 B.n847 B.n121 585
R1118 B.n121 B.n120 585
R1119 B.n846 B.n845 585
R1120 B.n845 B.n844 585
R1121 B.n123 B.n122 585
R1122 B.n843 B.n123 585
R1123 B.n841 B.n840 585
R1124 B.n842 B.n841 585
R1125 B.n982 B.n981 585
R1126 B.n981 B.n980 585
R1127 B.n434 B.n297 540.549
R1128 B.n841 B.n128 540.549
R1129 B.n436 B.n295 540.549
R1130 B.n734 B.n126 540.549
R1131 B.n735 B.n127 256.663
R1132 B.n741 B.n127 256.663
R1133 B.n743 B.n127 256.663
R1134 B.n749 B.n127 256.663
R1135 B.n751 B.n127 256.663
R1136 B.n757 B.n127 256.663
R1137 B.n759 B.n127 256.663
R1138 B.n765 B.n127 256.663
R1139 B.n767 B.n127 256.663
R1140 B.n773 B.n127 256.663
R1141 B.n775 B.n127 256.663
R1142 B.n782 B.n127 256.663
R1143 B.n784 B.n127 256.663
R1144 B.n790 B.n127 256.663
R1145 B.n142 B.n127 256.663
R1146 B.n796 B.n127 256.663
R1147 B.n802 B.n127 256.663
R1148 B.n804 B.n127 256.663
R1149 B.n810 B.n127 256.663
R1150 B.n812 B.n127 256.663
R1151 B.n818 B.n127 256.663
R1152 B.n820 B.n127 256.663
R1153 B.n826 B.n127 256.663
R1154 B.n828 B.n127 256.663
R1155 B.n834 B.n127 256.663
R1156 B.n836 B.n127 256.663
R1157 B.n429 B.n296 256.663
R1158 B.n299 B.n296 256.663
R1159 B.n422 B.n296 256.663
R1160 B.n416 B.n296 256.663
R1161 B.n414 B.n296 256.663
R1162 B.n408 B.n296 256.663
R1163 B.n406 B.n296 256.663
R1164 B.n400 B.n296 256.663
R1165 B.n398 B.n296 256.663
R1166 B.n392 B.n296 256.663
R1167 B.n390 B.n296 256.663
R1168 B.n384 B.n296 256.663
R1169 B.n382 B.n296 256.663
R1170 B.n376 B.n296 256.663
R1171 B.n374 B.n296 256.663
R1172 B.n367 B.n296 256.663
R1173 B.n365 B.n296 256.663
R1174 B.n359 B.n296 256.663
R1175 B.n357 B.n296 256.663
R1176 B.n351 B.n296 256.663
R1177 B.n349 B.n296 256.663
R1178 B.n343 B.n296 256.663
R1179 B.n341 B.n296 256.663
R1180 B.n335 B.n296 256.663
R1181 B.n333 B.n296 256.663
R1182 B.n328 B.n296 256.663
R1183 B.n317 B.t18 248.38
R1184 B.n310 B.t10 248.38
R1185 B.n139 B.t21 248.38
R1186 B.n147 B.t14 248.38
R1187 B.n317 B.t20 234.065
R1188 B.n147 B.t16 234.065
R1189 B.n310 B.t13 234.065
R1190 B.n139 B.t22 234.065
R1191 B.n318 B.t19 165.798
R1192 B.n148 B.t17 165.798
R1193 B.n311 B.t12 165.798
R1194 B.n140 B.t23 165.798
R1195 B.n434 B.n291 163.367
R1196 B.n442 B.n291 163.367
R1197 B.n442 B.n289 163.367
R1198 B.n446 B.n289 163.367
R1199 B.n446 B.n283 163.367
R1200 B.n454 B.n283 163.367
R1201 B.n454 B.n281 163.367
R1202 B.n458 B.n281 163.367
R1203 B.n458 B.n275 163.367
R1204 B.n466 B.n275 163.367
R1205 B.n466 B.n273 163.367
R1206 B.n470 B.n273 163.367
R1207 B.n470 B.n267 163.367
R1208 B.n478 B.n267 163.367
R1209 B.n478 B.n265 163.367
R1210 B.n482 B.n265 163.367
R1211 B.n482 B.n259 163.367
R1212 B.n490 B.n259 163.367
R1213 B.n490 B.n257 163.367
R1214 B.n494 B.n257 163.367
R1215 B.n494 B.n251 163.367
R1216 B.n502 B.n251 163.367
R1217 B.n502 B.n249 163.367
R1218 B.n506 B.n249 163.367
R1219 B.n506 B.n243 163.367
R1220 B.n514 B.n243 163.367
R1221 B.n514 B.n241 163.367
R1222 B.n518 B.n241 163.367
R1223 B.n518 B.n235 163.367
R1224 B.n526 B.n235 163.367
R1225 B.n526 B.n233 163.367
R1226 B.n530 B.n233 163.367
R1227 B.n530 B.n227 163.367
R1228 B.n538 B.n227 163.367
R1229 B.n538 B.n225 163.367
R1230 B.n542 B.n225 163.367
R1231 B.n542 B.n219 163.367
R1232 B.n550 B.n219 163.367
R1233 B.n550 B.n217 163.367
R1234 B.n554 B.n217 163.367
R1235 B.n554 B.n211 163.367
R1236 B.n562 B.n211 163.367
R1237 B.n562 B.n209 163.367
R1238 B.n566 B.n209 163.367
R1239 B.n566 B.n203 163.367
R1240 B.n574 B.n203 163.367
R1241 B.n574 B.n201 163.367
R1242 B.n578 B.n201 163.367
R1243 B.n578 B.n195 163.367
R1244 B.n586 B.n195 163.367
R1245 B.n586 B.n193 163.367
R1246 B.n590 B.n193 163.367
R1247 B.n590 B.n187 163.367
R1248 B.n598 B.n187 163.367
R1249 B.n598 B.n185 163.367
R1250 B.n602 B.n185 163.367
R1251 B.n602 B.n179 163.367
R1252 B.n610 B.n179 163.367
R1253 B.n610 B.n177 163.367
R1254 B.n614 B.n177 163.367
R1255 B.n614 B.n171 163.367
R1256 B.n623 B.n171 163.367
R1257 B.n623 B.n169 163.367
R1258 B.n627 B.n169 163.367
R1259 B.n627 B.n164 163.367
R1260 B.n636 B.n164 163.367
R1261 B.n636 B.n162 163.367
R1262 B.n640 B.n162 163.367
R1263 B.n640 B.n2 163.367
R1264 B.n981 B.n2 163.367
R1265 B.n981 B.n3 163.367
R1266 B.n977 B.n3 163.367
R1267 B.n977 B.n9 163.367
R1268 B.n973 B.n9 163.367
R1269 B.n973 B.n11 163.367
R1270 B.n969 B.n11 163.367
R1271 B.n969 B.n15 163.367
R1272 B.n965 B.n15 163.367
R1273 B.n965 B.n17 163.367
R1274 B.n961 B.n17 163.367
R1275 B.n961 B.n23 163.367
R1276 B.n957 B.n23 163.367
R1277 B.n957 B.n25 163.367
R1278 B.n953 B.n25 163.367
R1279 B.n953 B.n30 163.367
R1280 B.n949 B.n30 163.367
R1281 B.n949 B.n32 163.367
R1282 B.n945 B.n32 163.367
R1283 B.n945 B.n37 163.367
R1284 B.n941 B.n37 163.367
R1285 B.n941 B.n39 163.367
R1286 B.n937 B.n39 163.367
R1287 B.n937 B.n44 163.367
R1288 B.n933 B.n44 163.367
R1289 B.n933 B.n46 163.367
R1290 B.n929 B.n46 163.367
R1291 B.n929 B.n51 163.367
R1292 B.n925 B.n51 163.367
R1293 B.n925 B.n53 163.367
R1294 B.n921 B.n53 163.367
R1295 B.n921 B.n58 163.367
R1296 B.n917 B.n58 163.367
R1297 B.n917 B.n60 163.367
R1298 B.n913 B.n60 163.367
R1299 B.n913 B.n65 163.367
R1300 B.n909 B.n65 163.367
R1301 B.n909 B.n67 163.367
R1302 B.n905 B.n67 163.367
R1303 B.n905 B.n72 163.367
R1304 B.n901 B.n72 163.367
R1305 B.n901 B.n74 163.367
R1306 B.n897 B.n74 163.367
R1307 B.n897 B.n79 163.367
R1308 B.n893 B.n79 163.367
R1309 B.n893 B.n81 163.367
R1310 B.n889 B.n81 163.367
R1311 B.n889 B.n86 163.367
R1312 B.n885 B.n86 163.367
R1313 B.n885 B.n88 163.367
R1314 B.n881 B.n88 163.367
R1315 B.n881 B.n93 163.367
R1316 B.n877 B.n93 163.367
R1317 B.n877 B.n95 163.367
R1318 B.n873 B.n95 163.367
R1319 B.n873 B.n100 163.367
R1320 B.n869 B.n100 163.367
R1321 B.n869 B.n102 163.367
R1322 B.n865 B.n102 163.367
R1323 B.n865 B.n107 163.367
R1324 B.n861 B.n107 163.367
R1325 B.n861 B.n109 163.367
R1326 B.n857 B.n109 163.367
R1327 B.n857 B.n114 163.367
R1328 B.n853 B.n114 163.367
R1329 B.n853 B.n116 163.367
R1330 B.n849 B.n116 163.367
R1331 B.n849 B.n121 163.367
R1332 B.n845 B.n121 163.367
R1333 B.n845 B.n123 163.367
R1334 B.n841 B.n123 163.367
R1335 B.n430 B.n428 163.367
R1336 B.n428 B.n427 163.367
R1337 B.n424 B.n423 163.367
R1338 B.n421 B.n301 163.367
R1339 B.n417 B.n415 163.367
R1340 B.n413 B.n303 163.367
R1341 B.n409 B.n407 163.367
R1342 B.n405 B.n305 163.367
R1343 B.n401 B.n399 163.367
R1344 B.n397 B.n307 163.367
R1345 B.n393 B.n391 163.367
R1346 B.n389 B.n309 163.367
R1347 B.n385 B.n383 163.367
R1348 B.n381 B.n314 163.367
R1349 B.n377 B.n375 163.367
R1350 B.n373 B.n316 163.367
R1351 B.n368 B.n366 163.367
R1352 B.n364 B.n320 163.367
R1353 B.n360 B.n358 163.367
R1354 B.n356 B.n322 163.367
R1355 B.n352 B.n350 163.367
R1356 B.n348 B.n324 163.367
R1357 B.n344 B.n342 163.367
R1358 B.n340 B.n326 163.367
R1359 B.n336 B.n334 163.367
R1360 B.n332 B.n329 163.367
R1361 B.n436 B.n293 163.367
R1362 B.n440 B.n293 163.367
R1363 B.n440 B.n287 163.367
R1364 B.n448 B.n287 163.367
R1365 B.n448 B.n285 163.367
R1366 B.n452 B.n285 163.367
R1367 B.n452 B.n279 163.367
R1368 B.n460 B.n279 163.367
R1369 B.n460 B.n277 163.367
R1370 B.n464 B.n277 163.367
R1371 B.n464 B.n271 163.367
R1372 B.n472 B.n271 163.367
R1373 B.n472 B.n269 163.367
R1374 B.n476 B.n269 163.367
R1375 B.n476 B.n263 163.367
R1376 B.n484 B.n263 163.367
R1377 B.n484 B.n261 163.367
R1378 B.n488 B.n261 163.367
R1379 B.n488 B.n254 163.367
R1380 B.n496 B.n254 163.367
R1381 B.n496 B.n252 163.367
R1382 B.n500 B.n252 163.367
R1383 B.n500 B.n247 163.367
R1384 B.n508 B.n247 163.367
R1385 B.n508 B.n245 163.367
R1386 B.n512 B.n245 163.367
R1387 B.n512 B.n239 163.367
R1388 B.n520 B.n239 163.367
R1389 B.n520 B.n237 163.367
R1390 B.n524 B.n237 163.367
R1391 B.n524 B.n231 163.367
R1392 B.n532 B.n231 163.367
R1393 B.n532 B.n229 163.367
R1394 B.n536 B.n229 163.367
R1395 B.n536 B.n223 163.367
R1396 B.n544 B.n223 163.367
R1397 B.n544 B.n221 163.367
R1398 B.n548 B.n221 163.367
R1399 B.n548 B.n215 163.367
R1400 B.n556 B.n215 163.367
R1401 B.n556 B.n213 163.367
R1402 B.n560 B.n213 163.367
R1403 B.n560 B.n207 163.367
R1404 B.n568 B.n207 163.367
R1405 B.n568 B.n205 163.367
R1406 B.n572 B.n205 163.367
R1407 B.n572 B.n199 163.367
R1408 B.n580 B.n199 163.367
R1409 B.n580 B.n197 163.367
R1410 B.n584 B.n197 163.367
R1411 B.n584 B.n191 163.367
R1412 B.n592 B.n191 163.367
R1413 B.n592 B.n189 163.367
R1414 B.n596 B.n189 163.367
R1415 B.n596 B.n183 163.367
R1416 B.n604 B.n183 163.367
R1417 B.n604 B.n181 163.367
R1418 B.n608 B.n181 163.367
R1419 B.n608 B.n175 163.367
R1420 B.n616 B.n175 163.367
R1421 B.n616 B.n173 163.367
R1422 B.n620 B.n173 163.367
R1423 B.n620 B.n168 163.367
R1424 B.n629 B.n168 163.367
R1425 B.n629 B.n166 163.367
R1426 B.n634 B.n166 163.367
R1427 B.n634 B.n160 163.367
R1428 B.n642 B.n160 163.367
R1429 B.n643 B.n642 163.367
R1430 B.n643 B.n5 163.367
R1431 B.n6 B.n5 163.367
R1432 B.n7 B.n6 163.367
R1433 B.n648 B.n7 163.367
R1434 B.n648 B.n12 163.367
R1435 B.n13 B.n12 163.367
R1436 B.n14 B.n13 163.367
R1437 B.n653 B.n14 163.367
R1438 B.n653 B.n19 163.367
R1439 B.n20 B.n19 163.367
R1440 B.n21 B.n20 163.367
R1441 B.n658 B.n21 163.367
R1442 B.n658 B.n26 163.367
R1443 B.n27 B.n26 163.367
R1444 B.n28 B.n27 163.367
R1445 B.n663 B.n28 163.367
R1446 B.n663 B.n33 163.367
R1447 B.n34 B.n33 163.367
R1448 B.n35 B.n34 163.367
R1449 B.n668 B.n35 163.367
R1450 B.n668 B.n40 163.367
R1451 B.n41 B.n40 163.367
R1452 B.n42 B.n41 163.367
R1453 B.n673 B.n42 163.367
R1454 B.n673 B.n47 163.367
R1455 B.n48 B.n47 163.367
R1456 B.n49 B.n48 163.367
R1457 B.n678 B.n49 163.367
R1458 B.n678 B.n54 163.367
R1459 B.n55 B.n54 163.367
R1460 B.n56 B.n55 163.367
R1461 B.n683 B.n56 163.367
R1462 B.n683 B.n61 163.367
R1463 B.n62 B.n61 163.367
R1464 B.n63 B.n62 163.367
R1465 B.n688 B.n63 163.367
R1466 B.n688 B.n68 163.367
R1467 B.n69 B.n68 163.367
R1468 B.n70 B.n69 163.367
R1469 B.n693 B.n70 163.367
R1470 B.n693 B.n75 163.367
R1471 B.n76 B.n75 163.367
R1472 B.n77 B.n76 163.367
R1473 B.n698 B.n77 163.367
R1474 B.n698 B.n82 163.367
R1475 B.n83 B.n82 163.367
R1476 B.n84 B.n83 163.367
R1477 B.n703 B.n84 163.367
R1478 B.n703 B.n89 163.367
R1479 B.n90 B.n89 163.367
R1480 B.n91 B.n90 163.367
R1481 B.n708 B.n91 163.367
R1482 B.n708 B.n96 163.367
R1483 B.n97 B.n96 163.367
R1484 B.n98 B.n97 163.367
R1485 B.n713 B.n98 163.367
R1486 B.n713 B.n103 163.367
R1487 B.n104 B.n103 163.367
R1488 B.n105 B.n104 163.367
R1489 B.n718 B.n105 163.367
R1490 B.n718 B.n110 163.367
R1491 B.n111 B.n110 163.367
R1492 B.n112 B.n111 163.367
R1493 B.n723 B.n112 163.367
R1494 B.n723 B.n117 163.367
R1495 B.n118 B.n117 163.367
R1496 B.n119 B.n118 163.367
R1497 B.n728 B.n119 163.367
R1498 B.n728 B.n124 163.367
R1499 B.n125 B.n124 163.367
R1500 B.n126 B.n125 163.367
R1501 B.n837 B.n835 163.367
R1502 B.n833 B.n130 163.367
R1503 B.n829 B.n827 163.367
R1504 B.n825 B.n132 163.367
R1505 B.n821 B.n819 163.367
R1506 B.n817 B.n134 163.367
R1507 B.n813 B.n811 163.367
R1508 B.n809 B.n136 163.367
R1509 B.n805 B.n803 163.367
R1510 B.n801 B.n138 163.367
R1511 B.n797 B.n795 163.367
R1512 B.n792 B.n791 163.367
R1513 B.n789 B.n144 163.367
R1514 B.n785 B.n783 163.367
R1515 B.n781 B.n146 163.367
R1516 B.n776 B.n774 163.367
R1517 B.n772 B.n150 163.367
R1518 B.n768 B.n766 163.367
R1519 B.n764 B.n152 163.367
R1520 B.n760 B.n758 163.367
R1521 B.n756 B.n154 163.367
R1522 B.n752 B.n750 163.367
R1523 B.n748 B.n156 163.367
R1524 B.n744 B.n742 163.367
R1525 B.n740 B.n158 163.367
R1526 B.n736 B.n734 163.367
R1527 B.n435 B.n296 145.411
R1528 B.n842 B.n127 145.411
R1529 B.n429 B.n297 71.676
R1530 B.n427 B.n299 71.676
R1531 B.n423 B.n422 71.676
R1532 B.n416 B.n301 71.676
R1533 B.n415 B.n414 71.676
R1534 B.n408 B.n303 71.676
R1535 B.n407 B.n406 71.676
R1536 B.n400 B.n305 71.676
R1537 B.n399 B.n398 71.676
R1538 B.n392 B.n307 71.676
R1539 B.n391 B.n390 71.676
R1540 B.n384 B.n309 71.676
R1541 B.n383 B.n382 71.676
R1542 B.n376 B.n314 71.676
R1543 B.n375 B.n374 71.676
R1544 B.n367 B.n316 71.676
R1545 B.n366 B.n365 71.676
R1546 B.n359 B.n320 71.676
R1547 B.n358 B.n357 71.676
R1548 B.n351 B.n322 71.676
R1549 B.n350 B.n349 71.676
R1550 B.n343 B.n324 71.676
R1551 B.n342 B.n341 71.676
R1552 B.n335 B.n326 71.676
R1553 B.n334 B.n333 71.676
R1554 B.n329 B.n328 71.676
R1555 B.n836 B.n128 71.676
R1556 B.n835 B.n834 71.676
R1557 B.n828 B.n130 71.676
R1558 B.n827 B.n826 71.676
R1559 B.n820 B.n132 71.676
R1560 B.n819 B.n818 71.676
R1561 B.n812 B.n134 71.676
R1562 B.n811 B.n810 71.676
R1563 B.n804 B.n136 71.676
R1564 B.n803 B.n802 71.676
R1565 B.n796 B.n138 71.676
R1566 B.n795 B.n142 71.676
R1567 B.n791 B.n790 71.676
R1568 B.n784 B.n144 71.676
R1569 B.n783 B.n782 71.676
R1570 B.n775 B.n146 71.676
R1571 B.n774 B.n773 71.676
R1572 B.n767 B.n150 71.676
R1573 B.n766 B.n765 71.676
R1574 B.n759 B.n152 71.676
R1575 B.n758 B.n757 71.676
R1576 B.n751 B.n154 71.676
R1577 B.n750 B.n749 71.676
R1578 B.n743 B.n156 71.676
R1579 B.n742 B.n741 71.676
R1580 B.n735 B.n158 71.676
R1581 B.n736 B.n735 71.676
R1582 B.n741 B.n740 71.676
R1583 B.n744 B.n743 71.676
R1584 B.n749 B.n748 71.676
R1585 B.n752 B.n751 71.676
R1586 B.n757 B.n756 71.676
R1587 B.n760 B.n759 71.676
R1588 B.n765 B.n764 71.676
R1589 B.n768 B.n767 71.676
R1590 B.n773 B.n772 71.676
R1591 B.n776 B.n775 71.676
R1592 B.n782 B.n781 71.676
R1593 B.n785 B.n784 71.676
R1594 B.n790 B.n789 71.676
R1595 B.n792 B.n142 71.676
R1596 B.n797 B.n796 71.676
R1597 B.n802 B.n801 71.676
R1598 B.n805 B.n804 71.676
R1599 B.n810 B.n809 71.676
R1600 B.n813 B.n812 71.676
R1601 B.n818 B.n817 71.676
R1602 B.n821 B.n820 71.676
R1603 B.n826 B.n825 71.676
R1604 B.n829 B.n828 71.676
R1605 B.n834 B.n833 71.676
R1606 B.n837 B.n836 71.676
R1607 B.n430 B.n429 71.676
R1608 B.n424 B.n299 71.676
R1609 B.n422 B.n421 71.676
R1610 B.n417 B.n416 71.676
R1611 B.n414 B.n413 71.676
R1612 B.n409 B.n408 71.676
R1613 B.n406 B.n405 71.676
R1614 B.n401 B.n400 71.676
R1615 B.n398 B.n397 71.676
R1616 B.n393 B.n392 71.676
R1617 B.n390 B.n389 71.676
R1618 B.n385 B.n384 71.676
R1619 B.n382 B.n381 71.676
R1620 B.n377 B.n376 71.676
R1621 B.n374 B.n373 71.676
R1622 B.n368 B.n367 71.676
R1623 B.n365 B.n364 71.676
R1624 B.n360 B.n359 71.676
R1625 B.n357 B.n356 71.676
R1626 B.n352 B.n351 71.676
R1627 B.n349 B.n348 71.676
R1628 B.n344 B.n343 71.676
R1629 B.n341 B.n340 71.676
R1630 B.n336 B.n335 71.676
R1631 B.n333 B.n332 71.676
R1632 B.n328 B.n295 71.676
R1633 B.n435 B.n292 71.137
R1634 B.n441 B.n292 71.137
R1635 B.n441 B.n288 71.137
R1636 B.n447 B.n288 71.137
R1637 B.n447 B.n284 71.137
R1638 B.n453 B.n284 71.137
R1639 B.n453 B.n280 71.137
R1640 B.n459 B.n280 71.137
R1641 B.n465 B.n276 71.137
R1642 B.n465 B.n272 71.137
R1643 B.n471 B.n272 71.137
R1644 B.n471 B.n268 71.137
R1645 B.n477 B.n268 71.137
R1646 B.n477 B.n264 71.137
R1647 B.n483 B.n264 71.137
R1648 B.n483 B.n260 71.137
R1649 B.n489 B.n260 71.137
R1650 B.n489 B.n255 71.137
R1651 B.n495 B.n255 71.137
R1652 B.n495 B.n256 71.137
R1653 B.n501 B.n248 71.137
R1654 B.n507 B.n248 71.137
R1655 B.n507 B.n244 71.137
R1656 B.n513 B.n244 71.137
R1657 B.n513 B.n240 71.137
R1658 B.n519 B.n240 71.137
R1659 B.n519 B.n236 71.137
R1660 B.n525 B.n236 71.137
R1661 B.n525 B.n232 71.137
R1662 B.n531 B.n232 71.137
R1663 B.n537 B.n228 71.137
R1664 B.n537 B.n224 71.137
R1665 B.n543 B.n224 71.137
R1666 B.n543 B.n220 71.137
R1667 B.n549 B.n220 71.137
R1668 B.n549 B.n216 71.137
R1669 B.n555 B.n216 71.137
R1670 B.n555 B.n212 71.137
R1671 B.n561 B.n212 71.137
R1672 B.n567 B.n208 71.137
R1673 B.n567 B.n204 71.137
R1674 B.n573 B.n204 71.137
R1675 B.n573 B.n200 71.137
R1676 B.n579 B.n200 71.137
R1677 B.n579 B.n196 71.137
R1678 B.n585 B.n196 71.137
R1679 B.n585 B.n192 71.137
R1680 B.n591 B.n192 71.137
R1681 B.n597 B.n188 71.137
R1682 B.n597 B.n184 71.137
R1683 B.n603 B.n184 71.137
R1684 B.n603 B.n180 71.137
R1685 B.n609 B.n180 71.137
R1686 B.n609 B.n176 71.137
R1687 B.n615 B.n176 71.137
R1688 B.n615 B.n172 71.137
R1689 B.n622 B.n172 71.137
R1690 B.n622 B.n621 71.137
R1691 B.n628 B.n165 71.137
R1692 B.n635 B.n165 71.137
R1693 B.n635 B.n161 71.137
R1694 B.n641 B.n161 71.137
R1695 B.n641 B.n4 71.137
R1696 B.n980 B.n4 71.137
R1697 B.n980 B.n979 71.137
R1698 B.n979 B.n978 71.137
R1699 B.n978 B.n8 71.137
R1700 B.n972 B.n8 71.137
R1701 B.n972 B.n971 71.137
R1702 B.n971 B.n970 71.137
R1703 B.n964 B.n18 71.137
R1704 B.n964 B.n963 71.137
R1705 B.n963 B.n962 71.137
R1706 B.n962 B.n22 71.137
R1707 B.n956 B.n22 71.137
R1708 B.n956 B.n955 71.137
R1709 B.n955 B.n954 71.137
R1710 B.n954 B.n29 71.137
R1711 B.n948 B.n29 71.137
R1712 B.n948 B.n947 71.137
R1713 B.n946 B.n36 71.137
R1714 B.n940 B.n36 71.137
R1715 B.n940 B.n939 71.137
R1716 B.n939 B.n938 71.137
R1717 B.n938 B.n43 71.137
R1718 B.n932 B.n43 71.137
R1719 B.n932 B.n931 71.137
R1720 B.n931 B.n930 71.137
R1721 B.n930 B.n50 71.137
R1722 B.n924 B.n923 71.137
R1723 B.n923 B.n922 71.137
R1724 B.n922 B.n57 71.137
R1725 B.n916 B.n57 71.137
R1726 B.n916 B.n915 71.137
R1727 B.n915 B.n914 71.137
R1728 B.n914 B.n64 71.137
R1729 B.n908 B.n64 71.137
R1730 B.n908 B.n907 71.137
R1731 B.n906 B.n71 71.137
R1732 B.n900 B.n71 71.137
R1733 B.n900 B.n899 71.137
R1734 B.n899 B.n898 71.137
R1735 B.n898 B.n78 71.137
R1736 B.n892 B.n78 71.137
R1737 B.n892 B.n891 71.137
R1738 B.n891 B.n890 71.137
R1739 B.n890 B.n85 71.137
R1740 B.n884 B.n85 71.137
R1741 B.n883 B.n882 71.137
R1742 B.n882 B.n92 71.137
R1743 B.n876 B.n92 71.137
R1744 B.n876 B.n875 71.137
R1745 B.n875 B.n874 71.137
R1746 B.n874 B.n99 71.137
R1747 B.n868 B.n99 71.137
R1748 B.n868 B.n867 71.137
R1749 B.n867 B.n866 71.137
R1750 B.n866 B.n106 71.137
R1751 B.n860 B.n106 71.137
R1752 B.n860 B.n859 71.137
R1753 B.n858 B.n113 71.137
R1754 B.n852 B.n113 71.137
R1755 B.n852 B.n851 71.137
R1756 B.n851 B.n850 71.137
R1757 B.n850 B.n120 71.137
R1758 B.n844 B.n120 71.137
R1759 B.n844 B.n843 71.137
R1760 B.n843 B.n842 71.137
R1761 B.n318 B.n317 68.2672
R1762 B.n311 B.n310 68.2672
R1763 B.n140 B.n139 68.2672
R1764 B.n148 B.n147 68.2672
R1765 B.n591 B.t6 61.7219
R1766 B.t9 B.n946 61.7219
R1767 B.t0 B.n228 59.6296
R1768 B.n907 B.t7 59.6296
R1769 B.n371 B.n318 59.5399
R1770 B.n312 B.n311 59.5399
R1771 B.n141 B.n140 59.5399
R1772 B.n778 B.n148 59.5399
R1773 B.n256 B.t4 57.5373
R1774 B.t3 B.n883 57.5373
R1775 B.n628 B.t8 55.4451
R1776 B.n970 B.t2 55.4451
R1777 B.t11 B.n276 53.3529
R1778 B.n859 B.t15 53.3529
R1779 B.n561 B.t5 36.6149
R1780 B.n924 B.t1 36.6149
R1781 B.n840 B.n839 35.1225
R1782 B.n733 B.n732 35.1225
R1783 B.n437 B.n294 35.1225
R1784 B.n433 B.n432 35.1225
R1785 B.t5 B.n208 34.5226
R1786 B.t1 B.n50 34.5226
R1787 B B.n982 18.0485
R1788 B.n459 B.t11 17.7846
R1789 B.t15 B.n858 17.7846
R1790 B.n621 B.t8 15.6924
R1791 B.n18 B.t2 15.6924
R1792 B.n501 B.t4 13.6001
R1793 B.n884 B.t3 13.6001
R1794 B.n531 B.t0 11.5079
R1795 B.t7 B.n906 11.5079
R1796 B.n839 B.n838 10.6151
R1797 B.n838 B.n129 10.6151
R1798 B.n832 B.n129 10.6151
R1799 B.n832 B.n831 10.6151
R1800 B.n831 B.n830 10.6151
R1801 B.n830 B.n131 10.6151
R1802 B.n824 B.n131 10.6151
R1803 B.n824 B.n823 10.6151
R1804 B.n823 B.n822 10.6151
R1805 B.n822 B.n133 10.6151
R1806 B.n816 B.n133 10.6151
R1807 B.n816 B.n815 10.6151
R1808 B.n815 B.n814 10.6151
R1809 B.n814 B.n135 10.6151
R1810 B.n808 B.n135 10.6151
R1811 B.n808 B.n807 10.6151
R1812 B.n807 B.n806 10.6151
R1813 B.n806 B.n137 10.6151
R1814 B.n800 B.n137 10.6151
R1815 B.n800 B.n799 10.6151
R1816 B.n799 B.n798 10.6151
R1817 B.n794 B.n793 10.6151
R1818 B.n793 B.n143 10.6151
R1819 B.n788 B.n143 10.6151
R1820 B.n788 B.n787 10.6151
R1821 B.n787 B.n786 10.6151
R1822 B.n786 B.n145 10.6151
R1823 B.n780 B.n145 10.6151
R1824 B.n780 B.n779 10.6151
R1825 B.n777 B.n149 10.6151
R1826 B.n771 B.n149 10.6151
R1827 B.n771 B.n770 10.6151
R1828 B.n770 B.n769 10.6151
R1829 B.n769 B.n151 10.6151
R1830 B.n763 B.n151 10.6151
R1831 B.n763 B.n762 10.6151
R1832 B.n762 B.n761 10.6151
R1833 B.n761 B.n153 10.6151
R1834 B.n755 B.n153 10.6151
R1835 B.n755 B.n754 10.6151
R1836 B.n754 B.n753 10.6151
R1837 B.n753 B.n155 10.6151
R1838 B.n747 B.n155 10.6151
R1839 B.n747 B.n746 10.6151
R1840 B.n746 B.n745 10.6151
R1841 B.n745 B.n157 10.6151
R1842 B.n739 B.n157 10.6151
R1843 B.n739 B.n738 10.6151
R1844 B.n738 B.n737 10.6151
R1845 B.n737 B.n733 10.6151
R1846 B.n438 B.n437 10.6151
R1847 B.n439 B.n438 10.6151
R1848 B.n439 B.n286 10.6151
R1849 B.n449 B.n286 10.6151
R1850 B.n450 B.n449 10.6151
R1851 B.n451 B.n450 10.6151
R1852 B.n451 B.n278 10.6151
R1853 B.n461 B.n278 10.6151
R1854 B.n462 B.n461 10.6151
R1855 B.n463 B.n462 10.6151
R1856 B.n463 B.n270 10.6151
R1857 B.n473 B.n270 10.6151
R1858 B.n474 B.n473 10.6151
R1859 B.n475 B.n474 10.6151
R1860 B.n475 B.n262 10.6151
R1861 B.n485 B.n262 10.6151
R1862 B.n486 B.n485 10.6151
R1863 B.n487 B.n486 10.6151
R1864 B.n487 B.n253 10.6151
R1865 B.n497 B.n253 10.6151
R1866 B.n498 B.n497 10.6151
R1867 B.n499 B.n498 10.6151
R1868 B.n499 B.n246 10.6151
R1869 B.n509 B.n246 10.6151
R1870 B.n510 B.n509 10.6151
R1871 B.n511 B.n510 10.6151
R1872 B.n511 B.n238 10.6151
R1873 B.n521 B.n238 10.6151
R1874 B.n522 B.n521 10.6151
R1875 B.n523 B.n522 10.6151
R1876 B.n523 B.n230 10.6151
R1877 B.n533 B.n230 10.6151
R1878 B.n534 B.n533 10.6151
R1879 B.n535 B.n534 10.6151
R1880 B.n535 B.n222 10.6151
R1881 B.n545 B.n222 10.6151
R1882 B.n546 B.n545 10.6151
R1883 B.n547 B.n546 10.6151
R1884 B.n547 B.n214 10.6151
R1885 B.n557 B.n214 10.6151
R1886 B.n558 B.n557 10.6151
R1887 B.n559 B.n558 10.6151
R1888 B.n559 B.n206 10.6151
R1889 B.n569 B.n206 10.6151
R1890 B.n570 B.n569 10.6151
R1891 B.n571 B.n570 10.6151
R1892 B.n571 B.n198 10.6151
R1893 B.n581 B.n198 10.6151
R1894 B.n582 B.n581 10.6151
R1895 B.n583 B.n582 10.6151
R1896 B.n583 B.n190 10.6151
R1897 B.n593 B.n190 10.6151
R1898 B.n594 B.n593 10.6151
R1899 B.n595 B.n594 10.6151
R1900 B.n595 B.n182 10.6151
R1901 B.n605 B.n182 10.6151
R1902 B.n606 B.n605 10.6151
R1903 B.n607 B.n606 10.6151
R1904 B.n607 B.n174 10.6151
R1905 B.n617 B.n174 10.6151
R1906 B.n618 B.n617 10.6151
R1907 B.n619 B.n618 10.6151
R1908 B.n619 B.n167 10.6151
R1909 B.n630 B.n167 10.6151
R1910 B.n631 B.n630 10.6151
R1911 B.n633 B.n631 10.6151
R1912 B.n633 B.n632 10.6151
R1913 B.n632 B.n159 10.6151
R1914 B.n644 B.n159 10.6151
R1915 B.n645 B.n644 10.6151
R1916 B.n646 B.n645 10.6151
R1917 B.n647 B.n646 10.6151
R1918 B.n649 B.n647 10.6151
R1919 B.n650 B.n649 10.6151
R1920 B.n651 B.n650 10.6151
R1921 B.n652 B.n651 10.6151
R1922 B.n654 B.n652 10.6151
R1923 B.n655 B.n654 10.6151
R1924 B.n656 B.n655 10.6151
R1925 B.n657 B.n656 10.6151
R1926 B.n659 B.n657 10.6151
R1927 B.n660 B.n659 10.6151
R1928 B.n661 B.n660 10.6151
R1929 B.n662 B.n661 10.6151
R1930 B.n664 B.n662 10.6151
R1931 B.n665 B.n664 10.6151
R1932 B.n666 B.n665 10.6151
R1933 B.n667 B.n666 10.6151
R1934 B.n669 B.n667 10.6151
R1935 B.n670 B.n669 10.6151
R1936 B.n671 B.n670 10.6151
R1937 B.n672 B.n671 10.6151
R1938 B.n674 B.n672 10.6151
R1939 B.n675 B.n674 10.6151
R1940 B.n676 B.n675 10.6151
R1941 B.n677 B.n676 10.6151
R1942 B.n679 B.n677 10.6151
R1943 B.n680 B.n679 10.6151
R1944 B.n681 B.n680 10.6151
R1945 B.n682 B.n681 10.6151
R1946 B.n684 B.n682 10.6151
R1947 B.n685 B.n684 10.6151
R1948 B.n686 B.n685 10.6151
R1949 B.n687 B.n686 10.6151
R1950 B.n689 B.n687 10.6151
R1951 B.n690 B.n689 10.6151
R1952 B.n691 B.n690 10.6151
R1953 B.n692 B.n691 10.6151
R1954 B.n694 B.n692 10.6151
R1955 B.n695 B.n694 10.6151
R1956 B.n696 B.n695 10.6151
R1957 B.n697 B.n696 10.6151
R1958 B.n699 B.n697 10.6151
R1959 B.n700 B.n699 10.6151
R1960 B.n701 B.n700 10.6151
R1961 B.n702 B.n701 10.6151
R1962 B.n704 B.n702 10.6151
R1963 B.n705 B.n704 10.6151
R1964 B.n706 B.n705 10.6151
R1965 B.n707 B.n706 10.6151
R1966 B.n709 B.n707 10.6151
R1967 B.n710 B.n709 10.6151
R1968 B.n711 B.n710 10.6151
R1969 B.n712 B.n711 10.6151
R1970 B.n714 B.n712 10.6151
R1971 B.n715 B.n714 10.6151
R1972 B.n716 B.n715 10.6151
R1973 B.n717 B.n716 10.6151
R1974 B.n719 B.n717 10.6151
R1975 B.n720 B.n719 10.6151
R1976 B.n721 B.n720 10.6151
R1977 B.n722 B.n721 10.6151
R1978 B.n724 B.n722 10.6151
R1979 B.n725 B.n724 10.6151
R1980 B.n726 B.n725 10.6151
R1981 B.n727 B.n726 10.6151
R1982 B.n729 B.n727 10.6151
R1983 B.n730 B.n729 10.6151
R1984 B.n731 B.n730 10.6151
R1985 B.n732 B.n731 10.6151
R1986 B.n432 B.n431 10.6151
R1987 B.n431 B.n298 10.6151
R1988 B.n426 B.n298 10.6151
R1989 B.n426 B.n425 10.6151
R1990 B.n425 B.n300 10.6151
R1991 B.n420 B.n300 10.6151
R1992 B.n420 B.n419 10.6151
R1993 B.n419 B.n418 10.6151
R1994 B.n418 B.n302 10.6151
R1995 B.n412 B.n302 10.6151
R1996 B.n412 B.n411 10.6151
R1997 B.n411 B.n410 10.6151
R1998 B.n410 B.n304 10.6151
R1999 B.n404 B.n304 10.6151
R2000 B.n404 B.n403 10.6151
R2001 B.n403 B.n402 10.6151
R2002 B.n402 B.n306 10.6151
R2003 B.n396 B.n306 10.6151
R2004 B.n396 B.n395 10.6151
R2005 B.n395 B.n394 10.6151
R2006 B.n394 B.n308 10.6151
R2007 B.n388 B.n387 10.6151
R2008 B.n387 B.n386 10.6151
R2009 B.n386 B.n313 10.6151
R2010 B.n380 B.n313 10.6151
R2011 B.n380 B.n379 10.6151
R2012 B.n379 B.n378 10.6151
R2013 B.n378 B.n315 10.6151
R2014 B.n372 B.n315 10.6151
R2015 B.n370 B.n369 10.6151
R2016 B.n369 B.n319 10.6151
R2017 B.n363 B.n319 10.6151
R2018 B.n363 B.n362 10.6151
R2019 B.n362 B.n361 10.6151
R2020 B.n361 B.n321 10.6151
R2021 B.n355 B.n321 10.6151
R2022 B.n355 B.n354 10.6151
R2023 B.n354 B.n353 10.6151
R2024 B.n353 B.n323 10.6151
R2025 B.n347 B.n323 10.6151
R2026 B.n347 B.n346 10.6151
R2027 B.n346 B.n345 10.6151
R2028 B.n345 B.n325 10.6151
R2029 B.n339 B.n325 10.6151
R2030 B.n339 B.n338 10.6151
R2031 B.n338 B.n337 10.6151
R2032 B.n337 B.n327 10.6151
R2033 B.n331 B.n327 10.6151
R2034 B.n331 B.n330 10.6151
R2035 B.n330 B.n294 10.6151
R2036 B.n433 B.n290 10.6151
R2037 B.n443 B.n290 10.6151
R2038 B.n444 B.n443 10.6151
R2039 B.n445 B.n444 10.6151
R2040 B.n445 B.n282 10.6151
R2041 B.n455 B.n282 10.6151
R2042 B.n456 B.n455 10.6151
R2043 B.n457 B.n456 10.6151
R2044 B.n457 B.n274 10.6151
R2045 B.n467 B.n274 10.6151
R2046 B.n468 B.n467 10.6151
R2047 B.n469 B.n468 10.6151
R2048 B.n469 B.n266 10.6151
R2049 B.n479 B.n266 10.6151
R2050 B.n480 B.n479 10.6151
R2051 B.n481 B.n480 10.6151
R2052 B.n481 B.n258 10.6151
R2053 B.n491 B.n258 10.6151
R2054 B.n492 B.n491 10.6151
R2055 B.n493 B.n492 10.6151
R2056 B.n493 B.n250 10.6151
R2057 B.n503 B.n250 10.6151
R2058 B.n504 B.n503 10.6151
R2059 B.n505 B.n504 10.6151
R2060 B.n505 B.n242 10.6151
R2061 B.n515 B.n242 10.6151
R2062 B.n516 B.n515 10.6151
R2063 B.n517 B.n516 10.6151
R2064 B.n517 B.n234 10.6151
R2065 B.n527 B.n234 10.6151
R2066 B.n528 B.n527 10.6151
R2067 B.n529 B.n528 10.6151
R2068 B.n529 B.n226 10.6151
R2069 B.n539 B.n226 10.6151
R2070 B.n540 B.n539 10.6151
R2071 B.n541 B.n540 10.6151
R2072 B.n541 B.n218 10.6151
R2073 B.n551 B.n218 10.6151
R2074 B.n552 B.n551 10.6151
R2075 B.n553 B.n552 10.6151
R2076 B.n553 B.n210 10.6151
R2077 B.n563 B.n210 10.6151
R2078 B.n564 B.n563 10.6151
R2079 B.n565 B.n564 10.6151
R2080 B.n565 B.n202 10.6151
R2081 B.n575 B.n202 10.6151
R2082 B.n576 B.n575 10.6151
R2083 B.n577 B.n576 10.6151
R2084 B.n577 B.n194 10.6151
R2085 B.n587 B.n194 10.6151
R2086 B.n588 B.n587 10.6151
R2087 B.n589 B.n588 10.6151
R2088 B.n589 B.n186 10.6151
R2089 B.n599 B.n186 10.6151
R2090 B.n600 B.n599 10.6151
R2091 B.n601 B.n600 10.6151
R2092 B.n601 B.n178 10.6151
R2093 B.n611 B.n178 10.6151
R2094 B.n612 B.n611 10.6151
R2095 B.n613 B.n612 10.6151
R2096 B.n613 B.n170 10.6151
R2097 B.n624 B.n170 10.6151
R2098 B.n625 B.n624 10.6151
R2099 B.n626 B.n625 10.6151
R2100 B.n626 B.n163 10.6151
R2101 B.n637 B.n163 10.6151
R2102 B.n638 B.n637 10.6151
R2103 B.n639 B.n638 10.6151
R2104 B.n639 B.n0 10.6151
R2105 B.n976 B.n1 10.6151
R2106 B.n976 B.n975 10.6151
R2107 B.n975 B.n974 10.6151
R2108 B.n974 B.n10 10.6151
R2109 B.n968 B.n10 10.6151
R2110 B.n968 B.n967 10.6151
R2111 B.n967 B.n966 10.6151
R2112 B.n966 B.n16 10.6151
R2113 B.n960 B.n16 10.6151
R2114 B.n960 B.n959 10.6151
R2115 B.n959 B.n958 10.6151
R2116 B.n958 B.n24 10.6151
R2117 B.n952 B.n24 10.6151
R2118 B.n952 B.n951 10.6151
R2119 B.n951 B.n950 10.6151
R2120 B.n950 B.n31 10.6151
R2121 B.n944 B.n31 10.6151
R2122 B.n944 B.n943 10.6151
R2123 B.n943 B.n942 10.6151
R2124 B.n942 B.n38 10.6151
R2125 B.n936 B.n38 10.6151
R2126 B.n936 B.n935 10.6151
R2127 B.n935 B.n934 10.6151
R2128 B.n934 B.n45 10.6151
R2129 B.n928 B.n45 10.6151
R2130 B.n928 B.n927 10.6151
R2131 B.n927 B.n926 10.6151
R2132 B.n926 B.n52 10.6151
R2133 B.n920 B.n52 10.6151
R2134 B.n920 B.n919 10.6151
R2135 B.n919 B.n918 10.6151
R2136 B.n918 B.n59 10.6151
R2137 B.n912 B.n59 10.6151
R2138 B.n912 B.n911 10.6151
R2139 B.n911 B.n910 10.6151
R2140 B.n910 B.n66 10.6151
R2141 B.n904 B.n66 10.6151
R2142 B.n904 B.n903 10.6151
R2143 B.n903 B.n902 10.6151
R2144 B.n902 B.n73 10.6151
R2145 B.n896 B.n73 10.6151
R2146 B.n896 B.n895 10.6151
R2147 B.n895 B.n894 10.6151
R2148 B.n894 B.n80 10.6151
R2149 B.n888 B.n80 10.6151
R2150 B.n888 B.n887 10.6151
R2151 B.n887 B.n886 10.6151
R2152 B.n886 B.n87 10.6151
R2153 B.n880 B.n87 10.6151
R2154 B.n880 B.n879 10.6151
R2155 B.n879 B.n878 10.6151
R2156 B.n878 B.n94 10.6151
R2157 B.n872 B.n94 10.6151
R2158 B.n872 B.n871 10.6151
R2159 B.n871 B.n870 10.6151
R2160 B.n870 B.n101 10.6151
R2161 B.n864 B.n101 10.6151
R2162 B.n864 B.n863 10.6151
R2163 B.n863 B.n862 10.6151
R2164 B.n862 B.n108 10.6151
R2165 B.n856 B.n108 10.6151
R2166 B.n856 B.n855 10.6151
R2167 B.n855 B.n854 10.6151
R2168 B.n854 B.n115 10.6151
R2169 B.n848 B.n115 10.6151
R2170 B.n848 B.n847 10.6151
R2171 B.n847 B.n846 10.6151
R2172 B.n846 B.n122 10.6151
R2173 B.n840 B.n122 10.6151
R2174 B.t6 B.n188 9.41562
R2175 B.n947 B.t9 9.41562
R2176 B.n794 B.n141 6.5566
R2177 B.n779 B.n778 6.5566
R2178 B.n388 B.n312 6.5566
R2179 B.n372 B.n371 6.5566
R2180 B.n798 B.n141 4.05904
R2181 B.n778 B.n777 4.05904
R2182 B.n312 B.n308 4.05904
R2183 B.n371 B.n370 4.05904
R2184 B.n982 B.n0 2.81026
R2185 B.n982 B.n1 2.81026
R2186 VP.n32 VP.n31 161.3
R2187 VP.n33 VP.n28 161.3
R2188 VP.n35 VP.n34 161.3
R2189 VP.n36 VP.n27 161.3
R2190 VP.n38 VP.n37 161.3
R2191 VP.n39 VP.n26 161.3
R2192 VP.n41 VP.n40 161.3
R2193 VP.n43 VP.n42 161.3
R2194 VP.n44 VP.n24 161.3
R2195 VP.n46 VP.n45 161.3
R2196 VP.n47 VP.n23 161.3
R2197 VP.n49 VP.n48 161.3
R2198 VP.n50 VP.n22 161.3
R2199 VP.n52 VP.n51 161.3
R2200 VP.n54 VP.n53 161.3
R2201 VP.n55 VP.n20 161.3
R2202 VP.n57 VP.n56 161.3
R2203 VP.n58 VP.n19 161.3
R2204 VP.n60 VP.n59 161.3
R2205 VP.n61 VP.n18 161.3
R2206 VP.n63 VP.n62 161.3
R2207 VP.n109 VP.n108 161.3
R2208 VP.n107 VP.n1 161.3
R2209 VP.n106 VP.n105 161.3
R2210 VP.n104 VP.n2 161.3
R2211 VP.n103 VP.n102 161.3
R2212 VP.n101 VP.n3 161.3
R2213 VP.n100 VP.n99 161.3
R2214 VP.n98 VP.n97 161.3
R2215 VP.n96 VP.n5 161.3
R2216 VP.n95 VP.n94 161.3
R2217 VP.n93 VP.n6 161.3
R2218 VP.n92 VP.n91 161.3
R2219 VP.n90 VP.n7 161.3
R2220 VP.n89 VP.n88 161.3
R2221 VP.n87 VP.n86 161.3
R2222 VP.n85 VP.n9 161.3
R2223 VP.n84 VP.n83 161.3
R2224 VP.n82 VP.n10 161.3
R2225 VP.n81 VP.n80 161.3
R2226 VP.n79 VP.n11 161.3
R2227 VP.n78 VP.n77 161.3
R2228 VP.n76 VP.n75 161.3
R2229 VP.n74 VP.n13 161.3
R2230 VP.n73 VP.n72 161.3
R2231 VP.n71 VP.n14 161.3
R2232 VP.n70 VP.n69 161.3
R2233 VP.n68 VP.n15 161.3
R2234 VP.n67 VP.n66 161.3
R2235 VP.n65 VP.n16 75.9823
R2236 VP.n110 VP.n0 75.9823
R2237 VP.n64 VP.n17 75.9823
R2238 VP.n30 VP.t2 72.5789
R2239 VP.n30 VP.n29 61.1843
R2240 VP.n65 VP.n64 51.2799
R2241 VP.n69 VP.n14 43.4833
R2242 VP.n106 VP.n2 43.4833
R2243 VP.n60 VP.n19 43.4833
R2244 VP.n80 VP.n10 41.5458
R2245 VP.n95 VP.n6 41.5458
R2246 VP.n49 VP.n23 41.5458
R2247 VP.n34 VP.n27 41.5458
R2248 VP.n84 VP.n10 39.6083
R2249 VP.n91 VP.n6 39.6083
R2250 VP.n45 VP.n23 39.6083
R2251 VP.n38 VP.n27 39.6083
R2252 VP.n16 VP.t6 39.588
R2253 VP.n12 VP.t4 39.588
R2254 VP.n8 VP.t3 39.588
R2255 VP.n4 VP.t8 39.588
R2256 VP.n0 VP.t5 39.588
R2257 VP.n17 VP.t0 39.588
R2258 VP.n21 VP.t7 39.588
R2259 VP.n25 VP.t1 39.588
R2260 VP.n29 VP.t9 39.588
R2261 VP.n73 VP.n14 37.6707
R2262 VP.n102 VP.n2 37.6707
R2263 VP.n56 VP.n19 37.6707
R2264 VP.n68 VP.n67 24.5923
R2265 VP.n69 VP.n68 24.5923
R2266 VP.n74 VP.n73 24.5923
R2267 VP.n75 VP.n74 24.5923
R2268 VP.n79 VP.n78 24.5923
R2269 VP.n80 VP.n79 24.5923
R2270 VP.n85 VP.n84 24.5923
R2271 VP.n86 VP.n85 24.5923
R2272 VP.n90 VP.n89 24.5923
R2273 VP.n91 VP.n90 24.5923
R2274 VP.n96 VP.n95 24.5923
R2275 VP.n97 VP.n96 24.5923
R2276 VP.n101 VP.n100 24.5923
R2277 VP.n102 VP.n101 24.5923
R2278 VP.n107 VP.n106 24.5923
R2279 VP.n108 VP.n107 24.5923
R2280 VP.n61 VP.n60 24.5923
R2281 VP.n62 VP.n61 24.5923
R2282 VP.n50 VP.n49 24.5923
R2283 VP.n51 VP.n50 24.5923
R2284 VP.n55 VP.n54 24.5923
R2285 VP.n56 VP.n55 24.5923
R2286 VP.n39 VP.n38 24.5923
R2287 VP.n40 VP.n39 24.5923
R2288 VP.n44 VP.n43 24.5923
R2289 VP.n45 VP.n44 24.5923
R2290 VP.n33 VP.n32 24.5923
R2291 VP.n34 VP.n33 24.5923
R2292 VP.n67 VP.n16 14.2638
R2293 VP.n108 VP.n0 14.2638
R2294 VP.n62 VP.n17 14.2638
R2295 VP.n78 VP.n12 13.2801
R2296 VP.n97 VP.n4 13.2801
R2297 VP.n51 VP.n21 13.2801
R2298 VP.n32 VP.n29 13.2801
R2299 VP.n86 VP.n8 12.2964
R2300 VP.n89 VP.n8 12.2964
R2301 VP.n40 VP.n25 12.2964
R2302 VP.n43 VP.n25 12.2964
R2303 VP.n75 VP.n12 11.3127
R2304 VP.n100 VP.n4 11.3127
R2305 VP.n54 VP.n21 11.3127
R2306 VP.n31 VP.n30 4.1672
R2307 VP.n64 VP.n63 0.354861
R2308 VP.n66 VP.n65 0.354861
R2309 VP.n110 VP.n109 0.354861
R2310 VP VP.n110 0.267071
R2311 VP.n31 VP.n28 0.189894
R2312 VP.n35 VP.n28 0.189894
R2313 VP.n36 VP.n35 0.189894
R2314 VP.n37 VP.n36 0.189894
R2315 VP.n37 VP.n26 0.189894
R2316 VP.n41 VP.n26 0.189894
R2317 VP.n42 VP.n41 0.189894
R2318 VP.n42 VP.n24 0.189894
R2319 VP.n46 VP.n24 0.189894
R2320 VP.n47 VP.n46 0.189894
R2321 VP.n48 VP.n47 0.189894
R2322 VP.n48 VP.n22 0.189894
R2323 VP.n52 VP.n22 0.189894
R2324 VP.n53 VP.n52 0.189894
R2325 VP.n53 VP.n20 0.189894
R2326 VP.n57 VP.n20 0.189894
R2327 VP.n58 VP.n57 0.189894
R2328 VP.n59 VP.n58 0.189894
R2329 VP.n59 VP.n18 0.189894
R2330 VP.n63 VP.n18 0.189894
R2331 VP.n66 VP.n15 0.189894
R2332 VP.n70 VP.n15 0.189894
R2333 VP.n71 VP.n70 0.189894
R2334 VP.n72 VP.n71 0.189894
R2335 VP.n72 VP.n13 0.189894
R2336 VP.n76 VP.n13 0.189894
R2337 VP.n77 VP.n76 0.189894
R2338 VP.n77 VP.n11 0.189894
R2339 VP.n81 VP.n11 0.189894
R2340 VP.n82 VP.n81 0.189894
R2341 VP.n83 VP.n82 0.189894
R2342 VP.n83 VP.n9 0.189894
R2343 VP.n87 VP.n9 0.189894
R2344 VP.n88 VP.n87 0.189894
R2345 VP.n88 VP.n7 0.189894
R2346 VP.n92 VP.n7 0.189894
R2347 VP.n93 VP.n92 0.189894
R2348 VP.n94 VP.n93 0.189894
R2349 VP.n94 VP.n5 0.189894
R2350 VP.n98 VP.n5 0.189894
R2351 VP.n99 VP.n98 0.189894
R2352 VP.n99 VP.n3 0.189894
R2353 VP.n103 VP.n3 0.189894
R2354 VP.n104 VP.n103 0.189894
R2355 VP.n105 VP.n104 0.189894
R2356 VP.n105 VP.n1 0.189894
R2357 VP.n109 VP.n1 0.189894
R2358 VDD1.n22 VDD1.n0 289.615
R2359 VDD1.n51 VDD1.n29 289.615
R2360 VDD1.n23 VDD1.n22 185
R2361 VDD1.n21 VDD1.n20 185
R2362 VDD1.n4 VDD1.n3 185
R2363 VDD1.n15 VDD1.n14 185
R2364 VDD1.n13 VDD1.n12 185
R2365 VDD1.n8 VDD1.n7 185
R2366 VDD1.n37 VDD1.n36 185
R2367 VDD1.n42 VDD1.n41 185
R2368 VDD1.n44 VDD1.n43 185
R2369 VDD1.n33 VDD1.n32 185
R2370 VDD1.n50 VDD1.n49 185
R2371 VDD1.n52 VDD1.n51 185
R2372 VDD1.n9 VDD1.t7 147.672
R2373 VDD1.n38 VDD1.t3 147.672
R2374 VDD1.n22 VDD1.n21 104.615
R2375 VDD1.n21 VDD1.n3 104.615
R2376 VDD1.n14 VDD1.n3 104.615
R2377 VDD1.n14 VDD1.n13 104.615
R2378 VDD1.n13 VDD1.n7 104.615
R2379 VDD1.n42 VDD1.n36 104.615
R2380 VDD1.n43 VDD1.n42 104.615
R2381 VDD1.n43 VDD1.n32 104.615
R2382 VDD1.n50 VDD1.n32 104.615
R2383 VDD1.n51 VDD1.n50 104.615
R2384 VDD1.n59 VDD1.n58 70.0999
R2385 VDD1.n28 VDD1.n27 67.8795
R2386 VDD1.n61 VDD1.n60 67.8794
R2387 VDD1.n57 VDD1.n56 67.8794
R2388 VDD1.t7 VDD1.n7 52.3082
R2389 VDD1.t3 VDD1.n36 52.3082
R2390 VDD1.n28 VDD1.n26 51.1229
R2391 VDD1.n57 VDD1.n55 51.1229
R2392 VDD1.n61 VDD1.n59 44.7466
R2393 VDD1.n9 VDD1.n8 15.6666
R2394 VDD1.n38 VDD1.n37 15.6666
R2395 VDD1.n12 VDD1.n11 12.8005
R2396 VDD1.n41 VDD1.n40 12.8005
R2397 VDD1.n15 VDD1.n6 12.0247
R2398 VDD1.n44 VDD1.n35 12.0247
R2399 VDD1.n16 VDD1.n4 11.249
R2400 VDD1.n45 VDD1.n33 11.249
R2401 VDD1.n20 VDD1.n19 10.4732
R2402 VDD1.n49 VDD1.n48 10.4732
R2403 VDD1.n23 VDD1.n2 9.69747
R2404 VDD1.n52 VDD1.n31 9.69747
R2405 VDD1.n26 VDD1.n25 9.45567
R2406 VDD1.n55 VDD1.n54 9.45567
R2407 VDD1.n25 VDD1.n24 9.3005
R2408 VDD1.n2 VDD1.n1 9.3005
R2409 VDD1.n19 VDD1.n18 9.3005
R2410 VDD1.n17 VDD1.n16 9.3005
R2411 VDD1.n6 VDD1.n5 9.3005
R2412 VDD1.n11 VDD1.n10 9.3005
R2413 VDD1.n54 VDD1.n53 9.3005
R2414 VDD1.n31 VDD1.n30 9.3005
R2415 VDD1.n48 VDD1.n47 9.3005
R2416 VDD1.n46 VDD1.n45 9.3005
R2417 VDD1.n35 VDD1.n34 9.3005
R2418 VDD1.n40 VDD1.n39 9.3005
R2419 VDD1.n24 VDD1.n0 8.92171
R2420 VDD1.n53 VDD1.n29 8.92171
R2421 VDD1.n26 VDD1.n0 5.04292
R2422 VDD1.n55 VDD1.n29 5.04292
R2423 VDD1.n10 VDD1.n9 4.38687
R2424 VDD1.n39 VDD1.n38 4.38687
R2425 VDD1.n24 VDD1.n23 4.26717
R2426 VDD1.n53 VDD1.n52 4.26717
R2427 VDD1.n60 VDD1.t2 3.77913
R2428 VDD1.n60 VDD1.t9 3.77913
R2429 VDD1.n27 VDD1.t0 3.77913
R2430 VDD1.n27 VDD1.t8 3.77913
R2431 VDD1.n58 VDD1.t1 3.77913
R2432 VDD1.n58 VDD1.t4 3.77913
R2433 VDD1.n56 VDD1.t5 3.77913
R2434 VDD1.n56 VDD1.t6 3.77913
R2435 VDD1.n20 VDD1.n2 3.49141
R2436 VDD1.n49 VDD1.n31 3.49141
R2437 VDD1.n19 VDD1.n4 2.71565
R2438 VDD1.n48 VDD1.n33 2.71565
R2439 VDD1 VDD1.n61 2.21817
R2440 VDD1.n16 VDD1.n15 1.93989
R2441 VDD1.n45 VDD1.n44 1.93989
R2442 VDD1.n12 VDD1.n6 1.16414
R2443 VDD1.n41 VDD1.n35 1.16414
R2444 VDD1 VDD1.n28 0.81731
R2445 VDD1.n59 VDD1.n57 0.703775
R2446 VDD1.n11 VDD1.n8 0.388379
R2447 VDD1.n40 VDD1.n37 0.388379
R2448 VDD1.n25 VDD1.n1 0.155672
R2449 VDD1.n18 VDD1.n1 0.155672
R2450 VDD1.n18 VDD1.n17 0.155672
R2451 VDD1.n17 VDD1.n5 0.155672
R2452 VDD1.n10 VDD1.n5 0.155672
R2453 VDD1.n39 VDD1.n34 0.155672
R2454 VDD1.n46 VDD1.n34 0.155672
R2455 VDD1.n47 VDD1.n46 0.155672
R2456 VDD1.n47 VDD1.n30 0.155672
R2457 VDD1.n54 VDD1.n30 0.155672
C0 VP VN 8.01165f
C1 VP VDD1 5.64863f
C2 VP VDD2 0.662615f
C3 VN VDD1 0.154682f
C4 VP VTAIL 6.62537f
C5 VN VDD2 5.14801f
C6 VDD1 VDD2 2.5555f
C7 VN VTAIL 6.6112f
C8 VTAIL VDD1 7.78989f
C9 VTAIL VDD2 7.84661f
C10 VDD2 B 6.766477f
C11 VDD1 B 6.686366f
C12 VTAIL B 5.395571f
C13 VN B 20.243671f
C14 VP B 18.784994f
C15 VDD1.n0 B 0.037303f
C16 VDD1.n1 B 0.027599f
C17 VDD1.n2 B 0.01483f
C18 VDD1.n3 B 0.035054f
C19 VDD1.n4 B 0.015703f
C20 VDD1.n5 B 0.027599f
C21 VDD1.n6 B 0.01483f
C22 VDD1.n7 B 0.02629f
C23 VDD1.n8 B 0.020702f
C24 VDD1.t7 B 0.057193f
C25 VDD1.n9 B 0.113089f
C26 VDD1.n10 B 0.560188f
C27 VDD1.n11 B 0.01483f
C28 VDD1.n12 B 0.015703f
C29 VDD1.n13 B 0.035054f
C30 VDD1.n14 B 0.035054f
C31 VDD1.n15 B 0.015703f
C32 VDD1.n16 B 0.01483f
C33 VDD1.n17 B 0.027599f
C34 VDD1.n18 B 0.027599f
C35 VDD1.n19 B 0.01483f
C36 VDD1.n20 B 0.015703f
C37 VDD1.n21 B 0.035054f
C38 VDD1.n22 B 0.073251f
C39 VDD1.n23 B 0.015703f
C40 VDD1.n24 B 0.01483f
C41 VDD1.n25 B 0.062286f
C42 VDD1.n26 B 0.078859f
C43 VDD1.t0 B 0.114282f
C44 VDD1.t8 B 0.114282f
C45 VDD1.n27 B 0.936511f
C46 VDD1.n28 B 0.866635f
C47 VDD1.n29 B 0.037303f
C48 VDD1.n30 B 0.027599f
C49 VDD1.n31 B 0.01483f
C50 VDD1.n32 B 0.035054f
C51 VDD1.n33 B 0.015703f
C52 VDD1.n34 B 0.027599f
C53 VDD1.n35 B 0.01483f
C54 VDD1.n36 B 0.02629f
C55 VDD1.n37 B 0.020702f
C56 VDD1.t3 B 0.057193f
C57 VDD1.n38 B 0.113089f
C58 VDD1.n39 B 0.560188f
C59 VDD1.n40 B 0.01483f
C60 VDD1.n41 B 0.015703f
C61 VDD1.n42 B 0.035054f
C62 VDD1.n43 B 0.035054f
C63 VDD1.n44 B 0.015703f
C64 VDD1.n45 B 0.01483f
C65 VDD1.n46 B 0.027599f
C66 VDD1.n47 B 0.027599f
C67 VDD1.n48 B 0.01483f
C68 VDD1.n49 B 0.015703f
C69 VDD1.n50 B 0.035054f
C70 VDD1.n51 B 0.073251f
C71 VDD1.n52 B 0.015703f
C72 VDD1.n53 B 0.01483f
C73 VDD1.n54 B 0.062286f
C74 VDD1.n55 B 0.078859f
C75 VDD1.t5 B 0.114282f
C76 VDD1.t6 B 0.114282f
C77 VDD1.n56 B 0.936506f
C78 VDD1.n57 B 0.857452f
C79 VDD1.t1 B 0.114282f
C80 VDD1.t4 B 0.114282f
C81 VDD1.n58 B 0.958675f
C82 VDD1.n59 B 3.23558f
C83 VDD1.t2 B 0.114282f
C84 VDD1.t9 B 0.114282f
C85 VDD1.n60 B 0.936506f
C86 VDD1.n61 B 3.19348f
C87 VP.t5 B 0.99001f
C88 VP.n0 B 0.45797f
C89 VP.n1 B 0.022569f
C90 VP.n2 B 0.018489f
C91 VP.n3 B 0.022569f
C92 VP.t8 B 0.99001f
C93 VP.n4 B 0.373084f
C94 VP.n5 B 0.022569f
C95 VP.n6 B 0.018257f
C96 VP.n7 B 0.022569f
C97 VP.t3 B 0.99001f
C98 VP.n8 B 0.373084f
C99 VP.n9 B 0.022569f
C100 VP.n10 B 0.018257f
C101 VP.n11 B 0.022569f
C102 VP.t4 B 0.99001f
C103 VP.n12 B 0.373084f
C104 VP.n13 B 0.022569f
C105 VP.n14 B 0.018489f
C106 VP.n15 B 0.022569f
C107 VP.t6 B 0.99001f
C108 VP.n16 B 0.45797f
C109 VP.t0 B 0.99001f
C110 VP.n17 B 0.45797f
C111 VP.n18 B 0.022569f
C112 VP.n19 B 0.018489f
C113 VP.n20 B 0.022569f
C114 VP.t7 B 0.99001f
C115 VP.n21 B 0.373084f
C116 VP.n22 B 0.022569f
C117 VP.n23 B 0.018257f
C118 VP.n24 B 0.022569f
C119 VP.t1 B 0.99001f
C120 VP.n25 B 0.373084f
C121 VP.n26 B 0.022569f
C122 VP.n27 B 0.018257f
C123 VP.n28 B 0.022569f
C124 VP.t9 B 0.99001f
C125 VP.n29 B 0.44754f
C126 VP.t2 B 1.2309f
C127 VP.n30 B 0.427308f
C128 VP.n31 B 0.262224f
C129 VP.n32 B 0.032349f
C130 VP.n33 B 0.041853f
C131 VP.n34 B 0.044382f
C132 VP.n35 B 0.022569f
C133 VP.n36 B 0.022569f
C134 VP.n37 B 0.022569f
C135 VP.n38 B 0.04483f
C136 VP.n39 B 0.041853f
C137 VP.n40 B 0.031522f
C138 VP.n41 B 0.022569f
C139 VP.n42 B 0.022569f
C140 VP.n43 B 0.031522f
C141 VP.n44 B 0.041853f
C142 VP.n45 B 0.04483f
C143 VP.n46 B 0.022569f
C144 VP.n47 B 0.022569f
C145 VP.n48 B 0.022569f
C146 VP.n49 B 0.044382f
C147 VP.n50 B 0.041853f
C148 VP.n51 B 0.032349f
C149 VP.n52 B 0.022569f
C150 VP.n53 B 0.022569f
C151 VP.n54 B 0.030696f
C152 VP.n55 B 0.041853f
C153 VP.n56 B 0.045153f
C154 VP.n57 B 0.022569f
C155 VP.n58 B 0.022569f
C156 VP.n59 B 0.022569f
C157 VP.n60 B 0.043828f
C158 VP.n61 B 0.041853f
C159 VP.n62 B 0.033175f
C160 VP.n63 B 0.036421f
C161 VP.n64 B 1.32953f
C162 VP.n65 B 1.3454f
C163 VP.n66 B 0.036421f
C164 VP.n67 B 0.033175f
C165 VP.n68 B 0.041853f
C166 VP.n69 B 0.043828f
C167 VP.n70 B 0.022569f
C168 VP.n71 B 0.022569f
C169 VP.n72 B 0.022569f
C170 VP.n73 B 0.045153f
C171 VP.n74 B 0.041853f
C172 VP.n75 B 0.030696f
C173 VP.n76 B 0.022569f
C174 VP.n77 B 0.022569f
C175 VP.n78 B 0.032349f
C176 VP.n79 B 0.041853f
C177 VP.n80 B 0.044382f
C178 VP.n81 B 0.022569f
C179 VP.n82 B 0.022569f
C180 VP.n83 B 0.022569f
C181 VP.n84 B 0.04483f
C182 VP.n85 B 0.041853f
C183 VP.n86 B 0.031522f
C184 VP.n87 B 0.022569f
C185 VP.n88 B 0.022569f
C186 VP.n89 B 0.031522f
C187 VP.n90 B 0.041853f
C188 VP.n91 B 0.04483f
C189 VP.n92 B 0.022569f
C190 VP.n93 B 0.022569f
C191 VP.n94 B 0.022569f
C192 VP.n95 B 0.044382f
C193 VP.n96 B 0.041853f
C194 VP.n97 B 0.032349f
C195 VP.n98 B 0.022569f
C196 VP.n99 B 0.022569f
C197 VP.n100 B 0.030696f
C198 VP.n101 B 0.041853f
C199 VP.n102 B 0.045153f
C200 VP.n103 B 0.022569f
C201 VP.n104 B 0.022569f
C202 VP.n105 B 0.022569f
C203 VP.n106 B 0.043828f
C204 VP.n107 B 0.041853f
C205 VP.n108 B 0.033175f
C206 VP.n109 B 0.036421f
C207 VP.n110 B 0.053966f
C208 VTAIL.t13 B 0.125303f
C209 VTAIL.t18 B 0.125303f
C210 VTAIL.n0 B 0.949719f
C211 VTAIL.n1 B 0.699764f
C212 VTAIL.n2 B 0.040901f
C213 VTAIL.n3 B 0.030261f
C214 VTAIL.n4 B 0.016261f
C215 VTAIL.n5 B 0.038434f
C216 VTAIL.n6 B 0.017217f
C217 VTAIL.n7 B 0.030261f
C218 VTAIL.n8 B 0.016261f
C219 VTAIL.n9 B 0.028826f
C220 VTAIL.n10 B 0.022698f
C221 VTAIL.t8 B 0.062709f
C222 VTAIL.n11 B 0.123996f
C223 VTAIL.n12 B 0.614212f
C224 VTAIL.n13 B 0.016261f
C225 VTAIL.n14 B 0.017217f
C226 VTAIL.n15 B 0.038434f
C227 VTAIL.n16 B 0.038434f
C228 VTAIL.n17 B 0.017217f
C229 VTAIL.n18 B 0.016261f
C230 VTAIL.n19 B 0.030261f
C231 VTAIL.n20 B 0.030261f
C232 VTAIL.n21 B 0.016261f
C233 VTAIL.n22 B 0.017217f
C234 VTAIL.n23 B 0.038434f
C235 VTAIL.n24 B 0.080316f
C236 VTAIL.n25 B 0.017217f
C237 VTAIL.n26 B 0.016261f
C238 VTAIL.n27 B 0.068292f
C239 VTAIL.n28 B 0.044592f
C240 VTAIL.n29 B 0.514545f
C241 VTAIL.t5 B 0.125303f
C242 VTAIL.t6 B 0.125303f
C243 VTAIL.n30 B 0.949719f
C244 VTAIL.n31 B 0.87019f
C245 VTAIL.t4 B 0.125303f
C246 VTAIL.t0 B 0.125303f
C247 VTAIL.n32 B 0.949719f
C248 VTAIL.n33 B 2.01758f
C249 VTAIL.t11 B 0.125303f
C250 VTAIL.t14 B 0.125303f
C251 VTAIL.n34 B 0.949726f
C252 VTAIL.n35 B 2.01758f
C253 VTAIL.t10 B 0.125303f
C254 VTAIL.t17 B 0.125303f
C255 VTAIL.n36 B 0.949726f
C256 VTAIL.n37 B 0.870183f
C257 VTAIL.n38 B 0.040901f
C258 VTAIL.n39 B 0.030261f
C259 VTAIL.n40 B 0.016261f
C260 VTAIL.n41 B 0.038434f
C261 VTAIL.n42 B 0.017217f
C262 VTAIL.n43 B 0.030261f
C263 VTAIL.n44 B 0.016261f
C264 VTAIL.n45 B 0.028826f
C265 VTAIL.n46 B 0.022698f
C266 VTAIL.t12 B 0.062709f
C267 VTAIL.n47 B 0.123996f
C268 VTAIL.n48 B 0.614212f
C269 VTAIL.n49 B 0.016261f
C270 VTAIL.n50 B 0.017217f
C271 VTAIL.n51 B 0.038434f
C272 VTAIL.n52 B 0.038434f
C273 VTAIL.n53 B 0.017217f
C274 VTAIL.n54 B 0.016261f
C275 VTAIL.n55 B 0.030261f
C276 VTAIL.n56 B 0.030261f
C277 VTAIL.n57 B 0.016261f
C278 VTAIL.n58 B 0.017217f
C279 VTAIL.n59 B 0.038434f
C280 VTAIL.n60 B 0.080316f
C281 VTAIL.n61 B 0.017217f
C282 VTAIL.n62 B 0.016261f
C283 VTAIL.n63 B 0.068292f
C284 VTAIL.n64 B 0.044592f
C285 VTAIL.n65 B 0.514545f
C286 VTAIL.t2 B 0.125303f
C287 VTAIL.t9 B 0.125303f
C288 VTAIL.n66 B 0.949726f
C289 VTAIL.n67 B 0.768054f
C290 VTAIL.t1 B 0.125303f
C291 VTAIL.t7 B 0.125303f
C292 VTAIL.n68 B 0.949726f
C293 VTAIL.n69 B 0.870183f
C294 VTAIL.n70 B 0.040901f
C295 VTAIL.n71 B 0.030261f
C296 VTAIL.n72 B 0.016261f
C297 VTAIL.n73 B 0.038434f
C298 VTAIL.n74 B 0.017217f
C299 VTAIL.n75 B 0.030261f
C300 VTAIL.n76 B 0.016261f
C301 VTAIL.n77 B 0.028826f
C302 VTAIL.n78 B 0.022698f
C303 VTAIL.t3 B 0.062709f
C304 VTAIL.n79 B 0.123996f
C305 VTAIL.n80 B 0.614212f
C306 VTAIL.n81 B 0.016261f
C307 VTAIL.n82 B 0.017217f
C308 VTAIL.n83 B 0.038434f
C309 VTAIL.n84 B 0.038434f
C310 VTAIL.n85 B 0.017217f
C311 VTAIL.n86 B 0.016261f
C312 VTAIL.n87 B 0.030261f
C313 VTAIL.n88 B 0.030261f
C314 VTAIL.n89 B 0.016261f
C315 VTAIL.n90 B 0.017217f
C316 VTAIL.n91 B 0.038434f
C317 VTAIL.n92 B 0.080316f
C318 VTAIL.n93 B 0.017217f
C319 VTAIL.n94 B 0.016261f
C320 VTAIL.n95 B 0.068292f
C321 VTAIL.n96 B 0.044592f
C322 VTAIL.n97 B 1.46819f
C323 VTAIL.n98 B 0.040901f
C324 VTAIL.n99 B 0.030261f
C325 VTAIL.n100 B 0.016261f
C326 VTAIL.n101 B 0.038434f
C327 VTAIL.n102 B 0.017217f
C328 VTAIL.n103 B 0.030261f
C329 VTAIL.n104 B 0.016261f
C330 VTAIL.n105 B 0.028826f
C331 VTAIL.n106 B 0.022698f
C332 VTAIL.t16 B 0.062709f
C333 VTAIL.n107 B 0.123996f
C334 VTAIL.n108 B 0.614212f
C335 VTAIL.n109 B 0.016261f
C336 VTAIL.n110 B 0.017217f
C337 VTAIL.n111 B 0.038434f
C338 VTAIL.n112 B 0.038434f
C339 VTAIL.n113 B 0.017217f
C340 VTAIL.n114 B 0.016261f
C341 VTAIL.n115 B 0.030261f
C342 VTAIL.n116 B 0.030261f
C343 VTAIL.n117 B 0.016261f
C344 VTAIL.n118 B 0.017217f
C345 VTAIL.n119 B 0.038434f
C346 VTAIL.n120 B 0.080316f
C347 VTAIL.n121 B 0.017217f
C348 VTAIL.n122 B 0.016261f
C349 VTAIL.n123 B 0.068292f
C350 VTAIL.n124 B 0.044592f
C351 VTAIL.n125 B 1.46819f
C352 VTAIL.t15 B 0.125303f
C353 VTAIL.t19 B 0.125303f
C354 VTAIL.n126 B 0.949719f
C355 VTAIL.n127 B 0.642606f
C356 VDD2.n0 B 0.036369f
C357 VDD2.n1 B 0.026908f
C358 VDD2.n2 B 0.014459f
C359 VDD2.n3 B 0.034176f
C360 VDD2.n4 B 0.01531f
C361 VDD2.n5 B 0.026908f
C362 VDD2.n6 B 0.014459f
C363 VDD2.n7 B 0.025632f
C364 VDD2.n8 B 0.020184f
C365 VDD2.t0 B 0.055761f
C366 VDD2.n9 B 0.110258f
C367 VDD2.n10 B 0.546161f
C368 VDD2.n11 B 0.014459f
C369 VDD2.n12 B 0.01531f
C370 VDD2.n13 B 0.034176f
C371 VDD2.n14 B 0.034176f
C372 VDD2.n15 B 0.01531f
C373 VDD2.n16 B 0.014459f
C374 VDD2.n17 B 0.026908f
C375 VDD2.n18 B 0.026908f
C376 VDD2.n19 B 0.014459f
C377 VDD2.n20 B 0.01531f
C378 VDD2.n21 B 0.034176f
C379 VDD2.n22 B 0.071417f
C380 VDD2.n23 B 0.01531f
C381 VDD2.n24 B 0.014459f
C382 VDD2.n25 B 0.060726f
C383 VDD2.n26 B 0.076885f
C384 VDD2.t9 B 0.11142f
C385 VDD2.t4 B 0.11142f
C386 VDD2.n27 B 0.913058f
C387 VDD2.n28 B 0.835983f
C388 VDD2.t7 B 0.11142f
C389 VDD2.t8 B 0.11142f
C390 VDD2.n29 B 0.934672f
C391 VDD2.n30 B 3.00919f
C392 VDD2.n31 B 0.036369f
C393 VDD2.n32 B 0.026908f
C394 VDD2.n33 B 0.014459f
C395 VDD2.n34 B 0.034176f
C396 VDD2.n35 B 0.01531f
C397 VDD2.n36 B 0.026908f
C398 VDD2.n37 B 0.014459f
C399 VDD2.n38 B 0.025632f
C400 VDD2.n39 B 0.020184f
C401 VDD2.t2 B 0.055761f
C402 VDD2.n40 B 0.110258f
C403 VDD2.n41 B 0.546161f
C404 VDD2.n42 B 0.014459f
C405 VDD2.n43 B 0.01531f
C406 VDD2.n44 B 0.034176f
C407 VDD2.n45 B 0.034176f
C408 VDD2.n46 B 0.01531f
C409 VDD2.n47 B 0.014459f
C410 VDD2.n48 B 0.026908f
C411 VDD2.n49 B 0.026908f
C412 VDD2.n50 B 0.014459f
C413 VDD2.n51 B 0.01531f
C414 VDD2.n52 B 0.034176f
C415 VDD2.n53 B 0.071417f
C416 VDD2.n54 B 0.01531f
C417 VDD2.n55 B 0.014459f
C418 VDD2.n56 B 0.060726f
C419 VDD2.n57 B 0.058242f
C420 VDD2.n58 B 2.79178f
C421 VDD2.t3 B 0.11142f
C422 VDD2.t6 B 0.11142f
C423 VDD2.n59 B 0.913062f
C424 VDD2.n60 B 0.549507f
C425 VDD2.t5 B 0.11142f
C426 VDD2.t1 B 0.11142f
C427 VDD2.n61 B 0.934628f
C428 VN.t3 B 0.963991f
C429 VN.n0 B 0.445934f
C430 VN.n1 B 0.021976f
C431 VN.n2 B 0.018003f
C432 VN.n3 B 0.021976f
C433 VN.t0 B 0.963991f
C434 VN.n4 B 0.363278f
C435 VN.n5 B 0.021976f
C436 VN.n6 B 0.017777f
C437 VN.n7 B 0.021976f
C438 VN.t4 B 0.963991f
C439 VN.n8 B 0.363278f
C440 VN.n9 B 0.021976f
C441 VN.n10 B 0.017777f
C442 VN.n11 B 0.021976f
C443 VN.t1 B 0.963991f
C444 VN.n12 B 0.435778f
C445 VN.t6 B 1.19856f
C446 VN.n13 B 0.416077f
C447 VN.n14 B 0.255332f
C448 VN.n15 B 0.031498f
C449 VN.n16 B 0.040753f
C450 VN.n17 B 0.043216f
C451 VN.n18 B 0.021976f
C452 VN.n19 B 0.021976f
C453 VN.n20 B 0.021976f
C454 VN.n21 B 0.043651f
C455 VN.n22 B 0.040753f
C456 VN.n23 B 0.030694f
C457 VN.n24 B 0.021976f
C458 VN.n25 B 0.021976f
C459 VN.n26 B 0.030694f
C460 VN.n27 B 0.040753f
C461 VN.n28 B 0.043651f
C462 VN.n29 B 0.021976f
C463 VN.n30 B 0.021976f
C464 VN.n31 B 0.021976f
C465 VN.n32 B 0.043216f
C466 VN.n33 B 0.040753f
C467 VN.n34 B 0.031498f
C468 VN.n35 B 0.021976f
C469 VN.n36 B 0.021976f
C470 VN.n37 B 0.029889f
C471 VN.n38 B 0.040753f
C472 VN.n39 B 0.043966f
C473 VN.n40 B 0.021976f
C474 VN.n41 B 0.021976f
C475 VN.n42 B 0.021976f
C476 VN.n43 B 0.042676f
C477 VN.n44 B 0.040753f
C478 VN.n45 B 0.032303f
C479 VN.n46 B 0.035464f
C480 VN.n47 B 0.052548f
C481 VN.t8 B 0.963991f
C482 VN.n48 B 0.445934f
C483 VN.n49 B 0.021976f
C484 VN.n50 B 0.018003f
C485 VN.n51 B 0.021976f
C486 VN.t5 B 0.963991f
C487 VN.n52 B 0.363278f
C488 VN.n53 B 0.021976f
C489 VN.n54 B 0.017777f
C490 VN.n55 B 0.021976f
C491 VN.t9 B 0.963991f
C492 VN.n56 B 0.363278f
C493 VN.n57 B 0.021976f
C494 VN.n58 B 0.017777f
C495 VN.n59 B 0.021976f
C496 VN.t2 B 0.963991f
C497 VN.n60 B 0.435778f
C498 VN.t7 B 1.19856f
C499 VN.n61 B 0.416077f
C500 VN.n62 B 0.255332f
C501 VN.n63 B 0.031498f
C502 VN.n64 B 0.040753f
C503 VN.n65 B 0.043216f
C504 VN.n66 B 0.021976f
C505 VN.n67 B 0.021976f
C506 VN.n68 B 0.021976f
C507 VN.n69 B 0.043651f
C508 VN.n70 B 0.040753f
C509 VN.n71 B 0.030694f
C510 VN.n72 B 0.021976f
C511 VN.n73 B 0.021976f
C512 VN.n74 B 0.030694f
C513 VN.n75 B 0.040753f
C514 VN.n76 B 0.043651f
C515 VN.n77 B 0.021976f
C516 VN.n78 B 0.021976f
C517 VN.n79 B 0.021976f
C518 VN.n80 B 0.043216f
C519 VN.n81 B 0.040753f
C520 VN.n82 B 0.031498f
C521 VN.n83 B 0.021976f
C522 VN.n84 B 0.021976f
C523 VN.n85 B 0.029889f
C524 VN.n86 B 0.040753f
C525 VN.n87 B 0.043966f
C526 VN.n88 B 0.021976f
C527 VN.n89 B 0.021976f
C528 VN.n90 B 0.021976f
C529 VN.n91 B 0.042676f
C530 VN.n92 B 0.040753f
C531 VN.n93 B 0.032303f
C532 VN.n94 B 0.035464f
C533 VN.n95 B 1.3035f
.ends

