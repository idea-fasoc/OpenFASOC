* NGSPICE file created from diff_pair_sample_1565.ext - technology: sky130A

.subckt diff_pair_sample_1565 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t5 VP.t0 VDD1.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=5.5302 pd=29.14 as=2.3397 ps=14.51 w=14.18 l=2.49
X1 B.t17 B.t15 B.t16 B.t9 sky130_fd_pr__nfet_01v8 ad=5.5302 pd=29.14 as=0 ps=0 w=14.18 l=2.49
X2 VDD2.t3 VN.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.3397 pd=14.51 as=5.5302 ps=29.14 w=14.18 l=2.49
X3 VDD1.t1 VP.t1 VTAIL.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=2.3397 pd=14.51 as=5.5302 ps=29.14 w=14.18 l=2.49
X4 VTAIL.t0 VN.t1 VDD2.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=5.5302 pd=29.14 as=2.3397 ps=14.51 w=14.18 l=2.49
X5 VTAIL.t6 VN.t2 VDD2.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=5.5302 pd=29.14 as=2.3397 ps=14.51 w=14.18 l=2.49
X6 VDD2.t0 VN.t3 VTAIL.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=2.3397 pd=14.51 as=5.5302 ps=29.14 w=14.18 l=2.49
X7 VTAIL.t3 VP.t2 VDD1.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=5.5302 pd=29.14 as=2.3397 ps=14.51 w=14.18 l=2.49
X8 B.t14 B.t12 B.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=5.5302 pd=29.14 as=0 ps=0 w=14.18 l=2.49
X9 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=5.5302 pd=29.14 as=0 ps=0 w=14.18 l=2.49
X10 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=5.5302 pd=29.14 as=0 ps=0 w=14.18 l=2.49
X11 VDD1.t3 VP.t3 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.3397 pd=14.51 as=5.5302 ps=29.14 w=14.18 l=2.49
R0 VP.n4 VP.t2 172.669
R1 VP.n4 VP.t1 171.912
R2 VP.n14 VP.n0 161.3
R3 VP.n13 VP.n12 161.3
R4 VP.n11 VP.n1 161.3
R5 VP.n10 VP.n9 161.3
R6 VP.n8 VP.n2 161.3
R7 VP.n7 VP.n6 161.3
R8 VP.n3 VP.t0 137.244
R9 VP.n15 VP.t3 137.244
R10 VP.n5 VP.n3 103.038
R11 VP.n16 VP.n15 103.038
R12 VP.n9 VP.n1 56.5617
R13 VP.n5 VP.n4 52.1011
R14 VP.n8 VP.n7 24.5923
R15 VP.n9 VP.n8 24.5923
R16 VP.n13 VP.n1 24.5923
R17 VP.n14 VP.n13 24.5923
R18 VP.n7 VP.n3 7.86989
R19 VP.n15 VP.n14 7.86989
R20 VP.n6 VP.n5 0.278335
R21 VP.n16 VP.n0 0.278335
R22 VP.n6 VP.n2 0.189894
R23 VP.n10 VP.n2 0.189894
R24 VP.n11 VP.n10 0.189894
R25 VP.n12 VP.n11 0.189894
R26 VP.n12 VP.n0 0.189894
R27 VP VP.n16 0.153485
R28 VDD1 VDD1.n1 103.246
R29 VDD1 VDD1.n0 59.547
R30 VDD1.n0 VDD1.t0 1.39683
R31 VDD1.n0 VDD1.t1 1.39683
R32 VDD1.n1 VDD1.t2 1.39683
R33 VDD1.n1 VDD1.t3 1.39683
R34 VTAIL.n618 VTAIL.n546 289.615
R35 VTAIL.n72 VTAIL.n0 289.615
R36 VTAIL.n150 VTAIL.n78 289.615
R37 VTAIL.n228 VTAIL.n156 289.615
R38 VTAIL.n540 VTAIL.n468 289.615
R39 VTAIL.n462 VTAIL.n390 289.615
R40 VTAIL.n384 VTAIL.n312 289.615
R41 VTAIL.n306 VTAIL.n234 289.615
R42 VTAIL.n570 VTAIL.n569 185
R43 VTAIL.n575 VTAIL.n574 185
R44 VTAIL.n577 VTAIL.n576 185
R45 VTAIL.n566 VTAIL.n565 185
R46 VTAIL.n583 VTAIL.n582 185
R47 VTAIL.n585 VTAIL.n584 185
R48 VTAIL.n562 VTAIL.n561 185
R49 VTAIL.n592 VTAIL.n591 185
R50 VTAIL.n593 VTAIL.n560 185
R51 VTAIL.n595 VTAIL.n594 185
R52 VTAIL.n558 VTAIL.n557 185
R53 VTAIL.n601 VTAIL.n600 185
R54 VTAIL.n603 VTAIL.n602 185
R55 VTAIL.n554 VTAIL.n553 185
R56 VTAIL.n609 VTAIL.n608 185
R57 VTAIL.n611 VTAIL.n610 185
R58 VTAIL.n550 VTAIL.n549 185
R59 VTAIL.n617 VTAIL.n616 185
R60 VTAIL.n619 VTAIL.n618 185
R61 VTAIL.n24 VTAIL.n23 185
R62 VTAIL.n29 VTAIL.n28 185
R63 VTAIL.n31 VTAIL.n30 185
R64 VTAIL.n20 VTAIL.n19 185
R65 VTAIL.n37 VTAIL.n36 185
R66 VTAIL.n39 VTAIL.n38 185
R67 VTAIL.n16 VTAIL.n15 185
R68 VTAIL.n46 VTAIL.n45 185
R69 VTAIL.n47 VTAIL.n14 185
R70 VTAIL.n49 VTAIL.n48 185
R71 VTAIL.n12 VTAIL.n11 185
R72 VTAIL.n55 VTAIL.n54 185
R73 VTAIL.n57 VTAIL.n56 185
R74 VTAIL.n8 VTAIL.n7 185
R75 VTAIL.n63 VTAIL.n62 185
R76 VTAIL.n65 VTAIL.n64 185
R77 VTAIL.n4 VTAIL.n3 185
R78 VTAIL.n71 VTAIL.n70 185
R79 VTAIL.n73 VTAIL.n72 185
R80 VTAIL.n102 VTAIL.n101 185
R81 VTAIL.n107 VTAIL.n106 185
R82 VTAIL.n109 VTAIL.n108 185
R83 VTAIL.n98 VTAIL.n97 185
R84 VTAIL.n115 VTAIL.n114 185
R85 VTAIL.n117 VTAIL.n116 185
R86 VTAIL.n94 VTAIL.n93 185
R87 VTAIL.n124 VTAIL.n123 185
R88 VTAIL.n125 VTAIL.n92 185
R89 VTAIL.n127 VTAIL.n126 185
R90 VTAIL.n90 VTAIL.n89 185
R91 VTAIL.n133 VTAIL.n132 185
R92 VTAIL.n135 VTAIL.n134 185
R93 VTAIL.n86 VTAIL.n85 185
R94 VTAIL.n141 VTAIL.n140 185
R95 VTAIL.n143 VTAIL.n142 185
R96 VTAIL.n82 VTAIL.n81 185
R97 VTAIL.n149 VTAIL.n148 185
R98 VTAIL.n151 VTAIL.n150 185
R99 VTAIL.n180 VTAIL.n179 185
R100 VTAIL.n185 VTAIL.n184 185
R101 VTAIL.n187 VTAIL.n186 185
R102 VTAIL.n176 VTAIL.n175 185
R103 VTAIL.n193 VTAIL.n192 185
R104 VTAIL.n195 VTAIL.n194 185
R105 VTAIL.n172 VTAIL.n171 185
R106 VTAIL.n202 VTAIL.n201 185
R107 VTAIL.n203 VTAIL.n170 185
R108 VTAIL.n205 VTAIL.n204 185
R109 VTAIL.n168 VTAIL.n167 185
R110 VTAIL.n211 VTAIL.n210 185
R111 VTAIL.n213 VTAIL.n212 185
R112 VTAIL.n164 VTAIL.n163 185
R113 VTAIL.n219 VTAIL.n218 185
R114 VTAIL.n221 VTAIL.n220 185
R115 VTAIL.n160 VTAIL.n159 185
R116 VTAIL.n227 VTAIL.n226 185
R117 VTAIL.n229 VTAIL.n228 185
R118 VTAIL.n541 VTAIL.n540 185
R119 VTAIL.n539 VTAIL.n538 185
R120 VTAIL.n472 VTAIL.n471 185
R121 VTAIL.n533 VTAIL.n532 185
R122 VTAIL.n531 VTAIL.n530 185
R123 VTAIL.n476 VTAIL.n475 185
R124 VTAIL.n525 VTAIL.n524 185
R125 VTAIL.n523 VTAIL.n522 185
R126 VTAIL.n480 VTAIL.n479 185
R127 VTAIL.n517 VTAIL.n516 185
R128 VTAIL.n515 VTAIL.n482 185
R129 VTAIL.n514 VTAIL.n513 185
R130 VTAIL.n485 VTAIL.n483 185
R131 VTAIL.n508 VTAIL.n507 185
R132 VTAIL.n506 VTAIL.n505 185
R133 VTAIL.n489 VTAIL.n488 185
R134 VTAIL.n500 VTAIL.n499 185
R135 VTAIL.n498 VTAIL.n497 185
R136 VTAIL.n493 VTAIL.n492 185
R137 VTAIL.n463 VTAIL.n462 185
R138 VTAIL.n461 VTAIL.n460 185
R139 VTAIL.n394 VTAIL.n393 185
R140 VTAIL.n455 VTAIL.n454 185
R141 VTAIL.n453 VTAIL.n452 185
R142 VTAIL.n398 VTAIL.n397 185
R143 VTAIL.n447 VTAIL.n446 185
R144 VTAIL.n445 VTAIL.n444 185
R145 VTAIL.n402 VTAIL.n401 185
R146 VTAIL.n439 VTAIL.n438 185
R147 VTAIL.n437 VTAIL.n404 185
R148 VTAIL.n436 VTAIL.n435 185
R149 VTAIL.n407 VTAIL.n405 185
R150 VTAIL.n430 VTAIL.n429 185
R151 VTAIL.n428 VTAIL.n427 185
R152 VTAIL.n411 VTAIL.n410 185
R153 VTAIL.n422 VTAIL.n421 185
R154 VTAIL.n420 VTAIL.n419 185
R155 VTAIL.n415 VTAIL.n414 185
R156 VTAIL.n385 VTAIL.n384 185
R157 VTAIL.n383 VTAIL.n382 185
R158 VTAIL.n316 VTAIL.n315 185
R159 VTAIL.n377 VTAIL.n376 185
R160 VTAIL.n375 VTAIL.n374 185
R161 VTAIL.n320 VTAIL.n319 185
R162 VTAIL.n369 VTAIL.n368 185
R163 VTAIL.n367 VTAIL.n366 185
R164 VTAIL.n324 VTAIL.n323 185
R165 VTAIL.n361 VTAIL.n360 185
R166 VTAIL.n359 VTAIL.n326 185
R167 VTAIL.n358 VTAIL.n357 185
R168 VTAIL.n329 VTAIL.n327 185
R169 VTAIL.n352 VTAIL.n351 185
R170 VTAIL.n350 VTAIL.n349 185
R171 VTAIL.n333 VTAIL.n332 185
R172 VTAIL.n344 VTAIL.n343 185
R173 VTAIL.n342 VTAIL.n341 185
R174 VTAIL.n337 VTAIL.n336 185
R175 VTAIL.n307 VTAIL.n306 185
R176 VTAIL.n305 VTAIL.n304 185
R177 VTAIL.n238 VTAIL.n237 185
R178 VTAIL.n299 VTAIL.n298 185
R179 VTAIL.n297 VTAIL.n296 185
R180 VTAIL.n242 VTAIL.n241 185
R181 VTAIL.n291 VTAIL.n290 185
R182 VTAIL.n289 VTAIL.n288 185
R183 VTAIL.n246 VTAIL.n245 185
R184 VTAIL.n283 VTAIL.n282 185
R185 VTAIL.n281 VTAIL.n248 185
R186 VTAIL.n280 VTAIL.n279 185
R187 VTAIL.n251 VTAIL.n249 185
R188 VTAIL.n274 VTAIL.n273 185
R189 VTAIL.n272 VTAIL.n271 185
R190 VTAIL.n255 VTAIL.n254 185
R191 VTAIL.n266 VTAIL.n265 185
R192 VTAIL.n264 VTAIL.n263 185
R193 VTAIL.n259 VTAIL.n258 185
R194 VTAIL.n571 VTAIL.t1 149.524
R195 VTAIL.n25 VTAIL.t0 149.524
R196 VTAIL.n103 VTAIL.t2 149.524
R197 VTAIL.n181 VTAIL.t5 149.524
R198 VTAIL.n494 VTAIL.t4 149.524
R199 VTAIL.n416 VTAIL.t3 149.524
R200 VTAIL.n338 VTAIL.t7 149.524
R201 VTAIL.n260 VTAIL.t6 149.524
R202 VTAIL.n575 VTAIL.n569 104.615
R203 VTAIL.n576 VTAIL.n575 104.615
R204 VTAIL.n576 VTAIL.n565 104.615
R205 VTAIL.n583 VTAIL.n565 104.615
R206 VTAIL.n584 VTAIL.n583 104.615
R207 VTAIL.n584 VTAIL.n561 104.615
R208 VTAIL.n592 VTAIL.n561 104.615
R209 VTAIL.n593 VTAIL.n592 104.615
R210 VTAIL.n594 VTAIL.n593 104.615
R211 VTAIL.n594 VTAIL.n557 104.615
R212 VTAIL.n601 VTAIL.n557 104.615
R213 VTAIL.n602 VTAIL.n601 104.615
R214 VTAIL.n602 VTAIL.n553 104.615
R215 VTAIL.n609 VTAIL.n553 104.615
R216 VTAIL.n610 VTAIL.n609 104.615
R217 VTAIL.n610 VTAIL.n549 104.615
R218 VTAIL.n617 VTAIL.n549 104.615
R219 VTAIL.n618 VTAIL.n617 104.615
R220 VTAIL.n29 VTAIL.n23 104.615
R221 VTAIL.n30 VTAIL.n29 104.615
R222 VTAIL.n30 VTAIL.n19 104.615
R223 VTAIL.n37 VTAIL.n19 104.615
R224 VTAIL.n38 VTAIL.n37 104.615
R225 VTAIL.n38 VTAIL.n15 104.615
R226 VTAIL.n46 VTAIL.n15 104.615
R227 VTAIL.n47 VTAIL.n46 104.615
R228 VTAIL.n48 VTAIL.n47 104.615
R229 VTAIL.n48 VTAIL.n11 104.615
R230 VTAIL.n55 VTAIL.n11 104.615
R231 VTAIL.n56 VTAIL.n55 104.615
R232 VTAIL.n56 VTAIL.n7 104.615
R233 VTAIL.n63 VTAIL.n7 104.615
R234 VTAIL.n64 VTAIL.n63 104.615
R235 VTAIL.n64 VTAIL.n3 104.615
R236 VTAIL.n71 VTAIL.n3 104.615
R237 VTAIL.n72 VTAIL.n71 104.615
R238 VTAIL.n107 VTAIL.n101 104.615
R239 VTAIL.n108 VTAIL.n107 104.615
R240 VTAIL.n108 VTAIL.n97 104.615
R241 VTAIL.n115 VTAIL.n97 104.615
R242 VTAIL.n116 VTAIL.n115 104.615
R243 VTAIL.n116 VTAIL.n93 104.615
R244 VTAIL.n124 VTAIL.n93 104.615
R245 VTAIL.n125 VTAIL.n124 104.615
R246 VTAIL.n126 VTAIL.n125 104.615
R247 VTAIL.n126 VTAIL.n89 104.615
R248 VTAIL.n133 VTAIL.n89 104.615
R249 VTAIL.n134 VTAIL.n133 104.615
R250 VTAIL.n134 VTAIL.n85 104.615
R251 VTAIL.n141 VTAIL.n85 104.615
R252 VTAIL.n142 VTAIL.n141 104.615
R253 VTAIL.n142 VTAIL.n81 104.615
R254 VTAIL.n149 VTAIL.n81 104.615
R255 VTAIL.n150 VTAIL.n149 104.615
R256 VTAIL.n185 VTAIL.n179 104.615
R257 VTAIL.n186 VTAIL.n185 104.615
R258 VTAIL.n186 VTAIL.n175 104.615
R259 VTAIL.n193 VTAIL.n175 104.615
R260 VTAIL.n194 VTAIL.n193 104.615
R261 VTAIL.n194 VTAIL.n171 104.615
R262 VTAIL.n202 VTAIL.n171 104.615
R263 VTAIL.n203 VTAIL.n202 104.615
R264 VTAIL.n204 VTAIL.n203 104.615
R265 VTAIL.n204 VTAIL.n167 104.615
R266 VTAIL.n211 VTAIL.n167 104.615
R267 VTAIL.n212 VTAIL.n211 104.615
R268 VTAIL.n212 VTAIL.n163 104.615
R269 VTAIL.n219 VTAIL.n163 104.615
R270 VTAIL.n220 VTAIL.n219 104.615
R271 VTAIL.n220 VTAIL.n159 104.615
R272 VTAIL.n227 VTAIL.n159 104.615
R273 VTAIL.n228 VTAIL.n227 104.615
R274 VTAIL.n540 VTAIL.n539 104.615
R275 VTAIL.n539 VTAIL.n471 104.615
R276 VTAIL.n532 VTAIL.n471 104.615
R277 VTAIL.n532 VTAIL.n531 104.615
R278 VTAIL.n531 VTAIL.n475 104.615
R279 VTAIL.n524 VTAIL.n475 104.615
R280 VTAIL.n524 VTAIL.n523 104.615
R281 VTAIL.n523 VTAIL.n479 104.615
R282 VTAIL.n516 VTAIL.n479 104.615
R283 VTAIL.n516 VTAIL.n515 104.615
R284 VTAIL.n515 VTAIL.n514 104.615
R285 VTAIL.n514 VTAIL.n483 104.615
R286 VTAIL.n507 VTAIL.n483 104.615
R287 VTAIL.n507 VTAIL.n506 104.615
R288 VTAIL.n506 VTAIL.n488 104.615
R289 VTAIL.n499 VTAIL.n488 104.615
R290 VTAIL.n499 VTAIL.n498 104.615
R291 VTAIL.n498 VTAIL.n492 104.615
R292 VTAIL.n462 VTAIL.n461 104.615
R293 VTAIL.n461 VTAIL.n393 104.615
R294 VTAIL.n454 VTAIL.n393 104.615
R295 VTAIL.n454 VTAIL.n453 104.615
R296 VTAIL.n453 VTAIL.n397 104.615
R297 VTAIL.n446 VTAIL.n397 104.615
R298 VTAIL.n446 VTAIL.n445 104.615
R299 VTAIL.n445 VTAIL.n401 104.615
R300 VTAIL.n438 VTAIL.n401 104.615
R301 VTAIL.n438 VTAIL.n437 104.615
R302 VTAIL.n437 VTAIL.n436 104.615
R303 VTAIL.n436 VTAIL.n405 104.615
R304 VTAIL.n429 VTAIL.n405 104.615
R305 VTAIL.n429 VTAIL.n428 104.615
R306 VTAIL.n428 VTAIL.n410 104.615
R307 VTAIL.n421 VTAIL.n410 104.615
R308 VTAIL.n421 VTAIL.n420 104.615
R309 VTAIL.n420 VTAIL.n414 104.615
R310 VTAIL.n384 VTAIL.n383 104.615
R311 VTAIL.n383 VTAIL.n315 104.615
R312 VTAIL.n376 VTAIL.n315 104.615
R313 VTAIL.n376 VTAIL.n375 104.615
R314 VTAIL.n375 VTAIL.n319 104.615
R315 VTAIL.n368 VTAIL.n319 104.615
R316 VTAIL.n368 VTAIL.n367 104.615
R317 VTAIL.n367 VTAIL.n323 104.615
R318 VTAIL.n360 VTAIL.n323 104.615
R319 VTAIL.n360 VTAIL.n359 104.615
R320 VTAIL.n359 VTAIL.n358 104.615
R321 VTAIL.n358 VTAIL.n327 104.615
R322 VTAIL.n351 VTAIL.n327 104.615
R323 VTAIL.n351 VTAIL.n350 104.615
R324 VTAIL.n350 VTAIL.n332 104.615
R325 VTAIL.n343 VTAIL.n332 104.615
R326 VTAIL.n343 VTAIL.n342 104.615
R327 VTAIL.n342 VTAIL.n336 104.615
R328 VTAIL.n306 VTAIL.n305 104.615
R329 VTAIL.n305 VTAIL.n237 104.615
R330 VTAIL.n298 VTAIL.n237 104.615
R331 VTAIL.n298 VTAIL.n297 104.615
R332 VTAIL.n297 VTAIL.n241 104.615
R333 VTAIL.n290 VTAIL.n241 104.615
R334 VTAIL.n290 VTAIL.n289 104.615
R335 VTAIL.n289 VTAIL.n245 104.615
R336 VTAIL.n282 VTAIL.n245 104.615
R337 VTAIL.n282 VTAIL.n281 104.615
R338 VTAIL.n281 VTAIL.n280 104.615
R339 VTAIL.n280 VTAIL.n249 104.615
R340 VTAIL.n273 VTAIL.n249 104.615
R341 VTAIL.n273 VTAIL.n272 104.615
R342 VTAIL.n272 VTAIL.n254 104.615
R343 VTAIL.n265 VTAIL.n254 104.615
R344 VTAIL.n265 VTAIL.n264 104.615
R345 VTAIL.n264 VTAIL.n258 104.615
R346 VTAIL.t1 VTAIL.n569 52.3082
R347 VTAIL.t0 VTAIL.n23 52.3082
R348 VTAIL.t2 VTAIL.n101 52.3082
R349 VTAIL.t5 VTAIL.n179 52.3082
R350 VTAIL.t4 VTAIL.n492 52.3082
R351 VTAIL.t3 VTAIL.n414 52.3082
R352 VTAIL.t7 VTAIL.n336 52.3082
R353 VTAIL.t6 VTAIL.n258 52.3082
R354 VTAIL.n623 VTAIL.n622 30.246
R355 VTAIL.n77 VTAIL.n76 30.246
R356 VTAIL.n155 VTAIL.n154 30.246
R357 VTAIL.n233 VTAIL.n232 30.246
R358 VTAIL.n545 VTAIL.n544 30.246
R359 VTAIL.n467 VTAIL.n466 30.246
R360 VTAIL.n389 VTAIL.n388 30.246
R361 VTAIL.n311 VTAIL.n310 30.246
R362 VTAIL.n623 VTAIL.n545 27.0221
R363 VTAIL.n311 VTAIL.n233 27.0221
R364 VTAIL.n595 VTAIL.n560 13.1884
R365 VTAIL.n49 VTAIL.n14 13.1884
R366 VTAIL.n127 VTAIL.n92 13.1884
R367 VTAIL.n205 VTAIL.n170 13.1884
R368 VTAIL.n517 VTAIL.n482 13.1884
R369 VTAIL.n439 VTAIL.n404 13.1884
R370 VTAIL.n361 VTAIL.n326 13.1884
R371 VTAIL.n283 VTAIL.n248 13.1884
R372 VTAIL.n591 VTAIL.n590 12.8005
R373 VTAIL.n596 VTAIL.n558 12.8005
R374 VTAIL.n45 VTAIL.n44 12.8005
R375 VTAIL.n50 VTAIL.n12 12.8005
R376 VTAIL.n123 VTAIL.n122 12.8005
R377 VTAIL.n128 VTAIL.n90 12.8005
R378 VTAIL.n201 VTAIL.n200 12.8005
R379 VTAIL.n206 VTAIL.n168 12.8005
R380 VTAIL.n518 VTAIL.n480 12.8005
R381 VTAIL.n513 VTAIL.n484 12.8005
R382 VTAIL.n440 VTAIL.n402 12.8005
R383 VTAIL.n435 VTAIL.n406 12.8005
R384 VTAIL.n362 VTAIL.n324 12.8005
R385 VTAIL.n357 VTAIL.n328 12.8005
R386 VTAIL.n284 VTAIL.n246 12.8005
R387 VTAIL.n279 VTAIL.n250 12.8005
R388 VTAIL.n589 VTAIL.n562 12.0247
R389 VTAIL.n600 VTAIL.n599 12.0247
R390 VTAIL.n43 VTAIL.n16 12.0247
R391 VTAIL.n54 VTAIL.n53 12.0247
R392 VTAIL.n121 VTAIL.n94 12.0247
R393 VTAIL.n132 VTAIL.n131 12.0247
R394 VTAIL.n199 VTAIL.n172 12.0247
R395 VTAIL.n210 VTAIL.n209 12.0247
R396 VTAIL.n522 VTAIL.n521 12.0247
R397 VTAIL.n512 VTAIL.n485 12.0247
R398 VTAIL.n444 VTAIL.n443 12.0247
R399 VTAIL.n434 VTAIL.n407 12.0247
R400 VTAIL.n366 VTAIL.n365 12.0247
R401 VTAIL.n356 VTAIL.n329 12.0247
R402 VTAIL.n288 VTAIL.n287 12.0247
R403 VTAIL.n278 VTAIL.n251 12.0247
R404 VTAIL.n586 VTAIL.n585 11.249
R405 VTAIL.n603 VTAIL.n556 11.249
R406 VTAIL.n40 VTAIL.n39 11.249
R407 VTAIL.n57 VTAIL.n10 11.249
R408 VTAIL.n118 VTAIL.n117 11.249
R409 VTAIL.n135 VTAIL.n88 11.249
R410 VTAIL.n196 VTAIL.n195 11.249
R411 VTAIL.n213 VTAIL.n166 11.249
R412 VTAIL.n525 VTAIL.n478 11.249
R413 VTAIL.n509 VTAIL.n508 11.249
R414 VTAIL.n447 VTAIL.n400 11.249
R415 VTAIL.n431 VTAIL.n430 11.249
R416 VTAIL.n369 VTAIL.n322 11.249
R417 VTAIL.n353 VTAIL.n352 11.249
R418 VTAIL.n291 VTAIL.n244 11.249
R419 VTAIL.n275 VTAIL.n274 11.249
R420 VTAIL.n582 VTAIL.n564 10.4732
R421 VTAIL.n604 VTAIL.n554 10.4732
R422 VTAIL.n36 VTAIL.n18 10.4732
R423 VTAIL.n58 VTAIL.n8 10.4732
R424 VTAIL.n114 VTAIL.n96 10.4732
R425 VTAIL.n136 VTAIL.n86 10.4732
R426 VTAIL.n192 VTAIL.n174 10.4732
R427 VTAIL.n214 VTAIL.n164 10.4732
R428 VTAIL.n526 VTAIL.n476 10.4732
R429 VTAIL.n505 VTAIL.n487 10.4732
R430 VTAIL.n448 VTAIL.n398 10.4732
R431 VTAIL.n427 VTAIL.n409 10.4732
R432 VTAIL.n370 VTAIL.n320 10.4732
R433 VTAIL.n349 VTAIL.n331 10.4732
R434 VTAIL.n292 VTAIL.n242 10.4732
R435 VTAIL.n271 VTAIL.n253 10.4732
R436 VTAIL.n571 VTAIL.n570 10.2747
R437 VTAIL.n25 VTAIL.n24 10.2747
R438 VTAIL.n103 VTAIL.n102 10.2747
R439 VTAIL.n181 VTAIL.n180 10.2747
R440 VTAIL.n494 VTAIL.n493 10.2747
R441 VTAIL.n416 VTAIL.n415 10.2747
R442 VTAIL.n338 VTAIL.n337 10.2747
R443 VTAIL.n260 VTAIL.n259 10.2747
R444 VTAIL.n581 VTAIL.n566 9.69747
R445 VTAIL.n608 VTAIL.n607 9.69747
R446 VTAIL.n35 VTAIL.n20 9.69747
R447 VTAIL.n62 VTAIL.n61 9.69747
R448 VTAIL.n113 VTAIL.n98 9.69747
R449 VTAIL.n140 VTAIL.n139 9.69747
R450 VTAIL.n191 VTAIL.n176 9.69747
R451 VTAIL.n218 VTAIL.n217 9.69747
R452 VTAIL.n530 VTAIL.n529 9.69747
R453 VTAIL.n504 VTAIL.n489 9.69747
R454 VTAIL.n452 VTAIL.n451 9.69747
R455 VTAIL.n426 VTAIL.n411 9.69747
R456 VTAIL.n374 VTAIL.n373 9.69747
R457 VTAIL.n348 VTAIL.n333 9.69747
R458 VTAIL.n296 VTAIL.n295 9.69747
R459 VTAIL.n270 VTAIL.n255 9.69747
R460 VTAIL.n622 VTAIL.n621 9.45567
R461 VTAIL.n76 VTAIL.n75 9.45567
R462 VTAIL.n154 VTAIL.n153 9.45567
R463 VTAIL.n232 VTAIL.n231 9.45567
R464 VTAIL.n544 VTAIL.n543 9.45567
R465 VTAIL.n466 VTAIL.n465 9.45567
R466 VTAIL.n388 VTAIL.n387 9.45567
R467 VTAIL.n310 VTAIL.n309 9.45567
R468 VTAIL.n548 VTAIL.n547 9.3005
R469 VTAIL.n621 VTAIL.n620 9.3005
R470 VTAIL.n613 VTAIL.n612 9.3005
R471 VTAIL.n552 VTAIL.n551 9.3005
R472 VTAIL.n607 VTAIL.n606 9.3005
R473 VTAIL.n605 VTAIL.n604 9.3005
R474 VTAIL.n556 VTAIL.n555 9.3005
R475 VTAIL.n599 VTAIL.n598 9.3005
R476 VTAIL.n597 VTAIL.n596 9.3005
R477 VTAIL.n573 VTAIL.n572 9.3005
R478 VTAIL.n568 VTAIL.n567 9.3005
R479 VTAIL.n579 VTAIL.n578 9.3005
R480 VTAIL.n581 VTAIL.n580 9.3005
R481 VTAIL.n564 VTAIL.n563 9.3005
R482 VTAIL.n587 VTAIL.n586 9.3005
R483 VTAIL.n589 VTAIL.n588 9.3005
R484 VTAIL.n590 VTAIL.n559 9.3005
R485 VTAIL.n615 VTAIL.n614 9.3005
R486 VTAIL.n2 VTAIL.n1 9.3005
R487 VTAIL.n75 VTAIL.n74 9.3005
R488 VTAIL.n67 VTAIL.n66 9.3005
R489 VTAIL.n6 VTAIL.n5 9.3005
R490 VTAIL.n61 VTAIL.n60 9.3005
R491 VTAIL.n59 VTAIL.n58 9.3005
R492 VTAIL.n10 VTAIL.n9 9.3005
R493 VTAIL.n53 VTAIL.n52 9.3005
R494 VTAIL.n51 VTAIL.n50 9.3005
R495 VTAIL.n27 VTAIL.n26 9.3005
R496 VTAIL.n22 VTAIL.n21 9.3005
R497 VTAIL.n33 VTAIL.n32 9.3005
R498 VTAIL.n35 VTAIL.n34 9.3005
R499 VTAIL.n18 VTAIL.n17 9.3005
R500 VTAIL.n41 VTAIL.n40 9.3005
R501 VTAIL.n43 VTAIL.n42 9.3005
R502 VTAIL.n44 VTAIL.n13 9.3005
R503 VTAIL.n69 VTAIL.n68 9.3005
R504 VTAIL.n80 VTAIL.n79 9.3005
R505 VTAIL.n153 VTAIL.n152 9.3005
R506 VTAIL.n145 VTAIL.n144 9.3005
R507 VTAIL.n84 VTAIL.n83 9.3005
R508 VTAIL.n139 VTAIL.n138 9.3005
R509 VTAIL.n137 VTAIL.n136 9.3005
R510 VTAIL.n88 VTAIL.n87 9.3005
R511 VTAIL.n131 VTAIL.n130 9.3005
R512 VTAIL.n129 VTAIL.n128 9.3005
R513 VTAIL.n105 VTAIL.n104 9.3005
R514 VTAIL.n100 VTAIL.n99 9.3005
R515 VTAIL.n111 VTAIL.n110 9.3005
R516 VTAIL.n113 VTAIL.n112 9.3005
R517 VTAIL.n96 VTAIL.n95 9.3005
R518 VTAIL.n119 VTAIL.n118 9.3005
R519 VTAIL.n121 VTAIL.n120 9.3005
R520 VTAIL.n122 VTAIL.n91 9.3005
R521 VTAIL.n147 VTAIL.n146 9.3005
R522 VTAIL.n158 VTAIL.n157 9.3005
R523 VTAIL.n231 VTAIL.n230 9.3005
R524 VTAIL.n223 VTAIL.n222 9.3005
R525 VTAIL.n162 VTAIL.n161 9.3005
R526 VTAIL.n217 VTAIL.n216 9.3005
R527 VTAIL.n215 VTAIL.n214 9.3005
R528 VTAIL.n166 VTAIL.n165 9.3005
R529 VTAIL.n209 VTAIL.n208 9.3005
R530 VTAIL.n207 VTAIL.n206 9.3005
R531 VTAIL.n183 VTAIL.n182 9.3005
R532 VTAIL.n178 VTAIL.n177 9.3005
R533 VTAIL.n189 VTAIL.n188 9.3005
R534 VTAIL.n191 VTAIL.n190 9.3005
R535 VTAIL.n174 VTAIL.n173 9.3005
R536 VTAIL.n197 VTAIL.n196 9.3005
R537 VTAIL.n199 VTAIL.n198 9.3005
R538 VTAIL.n200 VTAIL.n169 9.3005
R539 VTAIL.n225 VTAIL.n224 9.3005
R540 VTAIL.n470 VTAIL.n469 9.3005
R541 VTAIL.n537 VTAIL.n536 9.3005
R542 VTAIL.n535 VTAIL.n534 9.3005
R543 VTAIL.n474 VTAIL.n473 9.3005
R544 VTAIL.n529 VTAIL.n528 9.3005
R545 VTAIL.n527 VTAIL.n526 9.3005
R546 VTAIL.n478 VTAIL.n477 9.3005
R547 VTAIL.n521 VTAIL.n520 9.3005
R548 VTAIL.n519 VTAIL.n518 9.3005
R549 VTAIL.n484 VTAIL.n481 9.3005
R550 VTAIL.n512 VTAIL.n511 9.3005
R551 VTAIL.n510 VTAIL.n509 9.3005
R552 VTAIL.n487 VTAIL.n486 9.3005
R553 VTAIL.n504 VTAIL.n503 9.3005
R554 VTAIL.n502 VTAIL.n501 9.3005
R555 VTAIL.n491 VTAIL.n490 9.3005
R556 VTAIL.n496 VTAIL.n495 9.3005
R557 VTAIL.n543 VTAIL.n542 9.3005
R558 VTAIL.n418 VTAIL.n417 9.3005
R559 VTAIL.n413 VTAIL.n412 9.3005
R560 VTAIL.n424 VTAIL.n423 9.3005
R561 VTAIL.n426 VTAIL.n425 9.3005
R562 VTAIL.n409 VTAIL.n408 9.3005
R563 VTAIL.n432 VTAIL.n431 9.3005
R564 VTAIL.n434 VTAIL.n433 9.3005
R565 VTAIL.n406 VTAIL.n403 9.3005
R566 VTAIL.n465 VTAIL.n464 9.3005
R567 VTAIL.n392 VTAIL.n391 9.3005
R568 VTAIL.n459 VTAIL.n458 9.3005
R569 VTAIL.n457 VTAIL.n456 9.3005
R570 VTAIL.n396 VTAIL.n395 9.3005
R571 VTAIL.n451 VTAIL.n450 9.3005
R572 VTAIL.n449 VTAIL.n448 9.3005
R573 VTAIL.n400 VTAIL.n399 9.3005
R574 VTAIL.n443 VTAIL.n442 9.3005
R575 VTAIL.n441 VTAIL.n440 9.3005
R576 VTAIL.n340 VTAIL.n339 9.3005
R577 VTAIL.n335 VTAIL.n334 9.3005
R578 VTAIL.n346 VTAIL.n345 9.3005
R579 VTAIL.n348 VTAIL.n347 9.3005
R580 VTAIL.n331 VTAIL.n330 9.3005
R581 VTAIL.n354 VTAIL.n353 9.3005
R582 VTAIL.n356 VTAIL.n355 9.3005
R583 VTAIL.n328 VTAIL.n325 9.3005
R584 VTAIL.n387 VTAIL.n386 9.3005
R585 VTAIL.n314 VTAIL.n313 9.3005
R586 VTAIL.n381 VTAIL.n380 9.3005
R587 VTAIL.n379 VTAIL.n378 9.3005
R588 VTAIL.n318 VTAIL.n317 9.3005
R589 VTAIL.n373 VTAIL.n372 9.3005
R590 VTAIL.n371 VTAIL.n370 9.3005
R591 VTAIL.n322 VTAIL.n321 9.3005
R592 VTAIL.n365 VTAIL.n364 9.3005
R593 VTAIL.n363 VTAIL.n362 9.3005
R594 VTAIL.n262 VTAIL.n261 9.3005
R595 VTAIL.n257 VTAIL.n256 9.3005
R596 VTAIL.n268 VTAIL.n267 9.3005
R597 VTAIL.n270 VTAIL.n269 9.3005
R598 VTAIL.n253 VTAIL.n252 9.3005
R599 VTAIL.n276 VTAIL.n275 9.3005
R600 VTAIL.n278 VTAIL.n277 9.3005
R601 VTAIL.n250 VTAIL.n247 9.3005
R602 VTAIL.n309 VTAIL.n308 9.3005
R603 VTAIL.n236 VTAIL.n235 9.3005
R604 VTAIL.n303 VTAIL.n302 9.3005
R605 VTAIL.n301 VTAIL.n300 9.3005
R606 VTAIL.n240 VTAIL.n239 9.3005
R607 VTAIL.n295 VTAIL.n294 9.3005
R608 VTAIL.n293 VTAIL.n292 9.3005
R609 VTAIL.n244 VTAIL.n243 9.3005
R610 VTAIL.n287 VTAIL.n286 9.3005
R611 VTAIL.n285 VTAIL.n284 9.3005
R612 VTAIL.n578 VTAIL.n577 8.92171
R613 VTAIL.n611 VTAIL.n552 8.92171
R614 VTAIL.n32 VTAIL.n31 8.92171
R615 VTAIL.n65 VTAIL.n6 8.92171
R616 VTAIL.n110 VTAIL.n109 8.92171
R617 VTAIL.n143 VTAIL.n84 8.92171
R618 VTAIL.n188 VTAIL.n187 8.92171
R619 VTAIL.n221 VTAIL.n162 8.92171
R620 VTAIL.n533 VTAIL.n474 8.92171
R621 VTAIL.n501 VTAIL.n500 8.92171
R622 VTAIL.n455 VTAIL.n396 8.92171
R623 VTAIL.n423 VTAIL.n422 8.92171
R624 VTAIL.n377 VTAIL.n318 8.92171
R625 VTAIL.n345 VTAIL.n344 8.92171
R626 VTAIL.n299 VTAIL.n240 8.92171
R627 VTAIL.n267 VTAIL.n266 8.92171
R628 VTAIL.n574 VTAIL.n568 8.14595
R629 VTAIL.n612 VTAIL.n550 8.14595
R630 VTAIL.n622 VTAIL.n546 8.14595
R631 VTAIL.n28 VTAIL.n22 8.14595
R632 VTAIL.n66 VTAIL.n4 8.14595
R633 VTAIL.n76 VTAIL.n0 8.14595
R634 VTAIL.n106 VTAIL.n100 8.14595
R635 VTAIL.n144 VTAIL.n82 8.14595
R636 VTAIL.n154 VTAIL.n78 8.14595
R637 VTAIL.n184 VTAIL.n178 8.14595
R638 VTAIL.n222 VTAIL.n160 8.14595
R639 VTAIL.n232 VTAIL.n156 8.14595
R640 VTAIL.n544 VTAIL.n468 8.14595
R641 VTAIL.n534 VTAIL.n472 8.14595
R642 VTAIL.n497 VTAIL.n491 8.14595
R643 VTAIL.n466 VTAIL.n390 8.14595
R644 VTAIL.n456 VTAIL.n394 8.14595
R645 VTAIL.n419 VTAIL.n413 8.14595
R646 VTAIL.n388 VTAIL.n312 8.14595
R647 VTAIL.n378 VTAIL.n316 8.14595
R648 VTAIL.n341 VTAIL.n335 8.14595
R649 VTAIL.n310 VTAIL.n234 8.14595
R650 VTAIL.n300 VTAIL.n238 8.14595
R651 VTAIL.n263 VTAIL.n257 8.14595
R652 VTAIL.n573 VTAIL.n570 7.3702
R653 VTAIL.n616 VTAIL.n615 7.3702
R654 VTAIL.n620 VTAIL.n619 7.3702
R655 VTAIL.n27 VTAIL.n24 7.3702
R656 VTAIL.n70 VTAIL.n69 7.3702
R657 VTAIL.n74 VTAIL.n73 7.3702
R658 VTAIL.n105 VTAIL.n102 7.3702
R659 VTAIL.n148 VTAIL.n147 7.3702
R660 VTAIL.n152 VTAIL.n151 7.3702
R661 VTAIL.n183 VTAIL.n180 7.3702
R662 VTAIL.n226 VTAIL.n225 7.3702
R663 VTAIL.n230 VTAIL.n229 7.3702
R664 VTAIL.n542 VTAIL.n541 7.3702
R665 VTAIL.n538 VTAIL.n537 7.3702
R666 VTAIL.n496 VTAIL.n493 7.3702
R667 VTAIL.n464 VTAIL.n463 7.3702
R668 VTAIL.n460 VTAIL.n459 7.3702
R669 VTAIL.n418 VTAIL.n415 7.3702
R670 VTAIL.n386 VTAIL.n385 7.3702
R671 VTAIL.n382 VTAIL.n381 7.3702
R672 VTAIL.n340 VTAIL.n337 7.3702
R673 VTAIL.n308 VTAIL.n307 7.3702
R674 VTAIL.n304 VTAIL.n303 7.3702
R675 VTAIL.n262 VTAIL.n259 7.3702
R676 VTAIL.n616 VTAIL.n548 6.59444
R677 VTAIL.n619 VTAIL.n548 6.59444
R678 VTAIL.n70 VTAIL.n2 6.59444
R679 VTAIL.n73 VTAIL.n2 6.59444
R680 VTAIL.n148 VTAIL.n80 6.59444
R681 VTAIL.n151 VTAIL.n80 6.59444
R682 VTAIL.n226 VTAIL.n158 6.59444
R683 VTAIL.n229 VTAIL.n158 6.59444
R684 VTAIL.n541 VTAIL.n470 6.59444
R685 VTAIL.n538 VTAIL.n470 6.59444
R686 VTAIL.n463 VTAIL.n392 6.59444
R687 VTAIL.n460 VTAIL.n392 6.59444
R688 VTAIL.n385 VTAIL.n314 6.59444
R689 VTAIL.n382 VTAIL.n314 6.59444
R690 VTAIL.n307 VTAIL.n236 6.59444
R691 VTAIL.n304 VTAIL.n236 6.59444
R692 VTAIL.n574 VTAIL.n573 5.81868
R693 VTAIL.n615 VTAIL.n550 5.81868
R694 VTAIL.n620 VTAIL.n546 5.81868
R695 VTAIL.n28 VTAIL.n27 5.81868
R696 VTAIL.n69 VTAIL.n4 5.81868
R697 VTAIL.n74 VTAIL.n0 5.81868
R698 VTAIL.n106 VTAIL.n105 5.81868
R699 VTAIL.n147 VTAIL.n82 5.81868
R700 VTAIL.n152 VTAIL.n78 5.81868
R701 VTAIL.n184 VTAIL.n183 5.81868
R702 VTAIL.n225 VTAIL.n160 5.81868
R703 VTAIL.n230 VTAIL.n156 5.81868
R704 VTAIL.n542 VTAIL.n468 5.81868
R705 VTAIL.n537 VTAIL.n472 5.81868
R706 VTAIL.n497 VTAIL.n496 5.81868
R707 VTAIL.n464 VTAIL.n390 5.81868
R708 VTAIL.n459 VTAIL.n394 5.81868
R709 VTAIL.n419 VTAIL.n418 5.81868
R710 VTAIL.n386 VTAIL.n312 5.81868
R711 VTAIL.n381 VTAIL.n316 5.81868
R712 VTAIL.n341 VTAIL.n340 5.81868
R713 VTAIL.n308 VTAIL.n234 5.81868
R714 VTAIL.n303 VTAIL.n238 5.81868
R715 VTAIL.n263 VTAIL.n262 5.81868
R716 VTAIL.n577 VTAIL.n568 5.04292
R717 VTAIL.n612 VTAIL.n611 5.04292
R718 VTAIL.n31 VTAIL.n22 5.04292
R719 VTAIL.n66 VTAIL.n65 5.04292
R720 VTAIL.n109 VTAIL.n100 5.04292
R721 VTAIL.n144 VTAIL.n143 5.04292
R722 VTAIL.n187 VTAIL.n178 5.04292
R723 VTAIL.n222 VTAIL.n221 5.04292
R724 VTAIL.n534 VTAIL.n533 5.04292
R725 VTAIL.n500 VTAIL.n491 5.04292
R726 VTAIL.n456 VTAIL.n455 5.04292
R727 VTAIL.n422 VTAIL.n413 5.04292
R728 VTAIL.n378 VTAIL.n377 5.04292
R729 VTAIL.n344 VTAIL.n335 5.04292
R730 VTAIL.n300 VTAIL.n299 5.04292
R731 VTAIL.n266 VTAIL.n257 5.04292
R732 VTAIL.n578 VTAIL.n566 4.26717
R733 VTAIL.n608 VTAIL.n552 4.26717
R734 VTAIL.n32 VTAIL.n20 4.26717
R735 VTAIL.n62 VTAIL.n6 4.26717
R736 VTAIL.n110 VTAIL.n98 4.26717
R737 VTAIL.n140 VTAIL.n84 4.26717
R738 VTAIL.n188 VTAIL.n176 4.26717
R739 VTAIL.n218 VTAIL.n162 4.26717
R740 VTAIL.n530 VTAIL.n474 4.26717
R741 VTAIL.n501 VTAIL.n489 4.26717
R742 VTAIL.n452 VTAIL.n396 4.26717
R743 VTAIL.n423 VTAIL.n411 4.26717
R744 VTAIL.n374 VTAIL.n318 4.26717
R745 VTAIL.n345 VTAIL.n333 4.26717
R746 VTAIL.n296 VTAIL.n240 4.26717
R747 VTAIL.n267 VTAIL.n255 4.26717
R748 VTAIL.n582 VTAIL.n581 3.49141
R749 VTAIL.n607 VTAIL.n554 3.49141
R750 VTAIL.n36 VTAIL.n35 3.49141
R751 VTAIL.n61 VTAIL.n8 3.49141
R752 VTAIL.n114 VTAIL.n113 3.49141
R753 VTAIL.n139 VTAIL.n86 3.49141
R754 VTAIL.n192 VTAIL.n191 3.49141
R755 VTAIL.n217 VTAIL.n164 3.49141
R756 VTAIL.n529 VTAIL.n476 3.49141
R757 VTAIL.n505 VTAIL.n504 3.49141
R758 VTAIL.n451 VTAIL.n398 3.49141
R759 VTAIL.n427 VTAIL.n426 3.49141
R760 VTAIL.n373 VTAIL.n320 3.49141
R761 VTAIL.n349 VTAIL.n348 3.49141
R762 VTAIL.n295 VTAIL.n242 3.49141
R763 VTAIL.n271 VTAIL.n270 3.49141
R764 VTAIL.n572 VTAIL.n571 2.84303
R765 VTAIL.n26 VTAIL.n25 2.84303
R766 VTAIL.n104 VTAIL.n103 2.84303
R767 VTAIL.n182 VTAIL.n181 2.84303
R768 VTAIL.n417 VTAIL.n416 2.84303
R769 VTAIL.n339 VTAIL.n338 2.84303
R770 VTAIL.n261 VTAIL.n260 2.84303
R771 VTAIL.n495 VTAIL.n494 2.84303
R772 VTAIL.n585 VTAIL.n564 2.71565
R773 VTAIL.n604 VTAIL.n603 2.71565
R774 VTAIL.n39 VTAIL.n18 2.71565
R775 VTAIL.n58 VTAIL.n57 2.71565
R776 VTAIL.n117 VTAIL.n96 2.71565
R777 VTAIL.n136 VTAIL.n135 2.71565
R778 VTAIL.n195 VTAIL.n174 2.71565
R779 VTAIL.n214 VTAIL.n213 2.71565
R780 VTAIL.n526 VTAIL.n525 2.71565
R781 VTAIL.n508 VTAIL.n487 2.71565
R782 VTAIL.n448 VTAIL.n447 2.71565
R783 VTAIL.n430 VTAIL.n409 2.71565
R784 VTAIL.n370 VTAIL.n369 2.71565
R785 VTAIL.n352 VTAIL.n331 2.71565
R786 VTAIL.n292 VTAIL.n291 2.71565
R787 VTAIL.n274 VTAIL.n253 2.71565
R788 VTAIL.n389 VTAIL.n311 2.43153
R789 VTAIL.n545 VTAIL.n467 2.43153
R790 VTAIL.n233 VTAIL.n155 2.43153
R791 VTAIL.n586 VTAIL.n562 1.93989
R792 VTAIL.n600 VTAIL.n556 1.93989
R793 VTAIL.n40 VTAIL.n16 1.93989
R794 VTAIL.n54 VTAIL.n10 1.93989
R795 VTAIL.n118 VTAIL.n94 1.93989
R796 VTAIL.n132 VTAIL.n88 1.93989
R797 VTAIL.n196 VTAIL.n172 1.93989
R798 VTAIL.n210 VTAIL.n166 1.93989
R799 VTAIL.n522 VTAIL.n478 1.93989
R800 VTAIL.n509 VTAIL.n485 1.93989
R801 VTAIL.n444 VTAIL.n400 1.93989
R802 VTAIL.n431 VTAIL.n407 1.93989
R803 VTAIL.n366 VTAIL.n322 1.93989
R804 VTAIL.n353 VTAIL.n329 1.93989
R805 VTAIL.n288 VTAIL.n244 1.93989
R806 VTAIL.n275 VTAIL.n251 1.93989
R807 VTAIL VTAIL.n77 1.27421
R808 VTAIL.n591 VTAIL.n589 1.16414
R809 VTAIL.n599 VTAIL.n558 1.16414
R810 VTAIL.n45 VTAIL.n43 1.16414
R811 VTAIL.n53 VTAIL.n12 1.16414
R812 VTAIL.n123 VTAIL.n121 1.16414
R813 VTAIL.n131 VTAIL.n90 1.16414
R814 VTAIL.n201 VTAIL.n199 1.16414
R815 VTAIL.n209 VTAIL.n168 1.16414
R816 VTAIL.n521 VTAIL.n480 1.16414
R817 VTAIL.n513 VTAIL.n512 1.16414
R818 VTAIL.n443 VTAIL.n402 1.16414
R819 VTAIL.n435 VTAIL.n434 1.16414
R820 VTAIL.n365 VTAIL.n324 1.16414
R821 VTAIL.n357 VTAIL.n356 1.16414
R822 VTAIL.n287 VTAIL.n246 1.16414
R823 VTAIL.n279 VTAIL.n278 1.16414
R824 VTAIL VTAIL.n623 1.15783
R825 VTAIL.n467 VTAIL.n389 0.470328
R826 VTAIL.n155 VTAIL.n77 0.470328
R827 VTAIL.n590 VTAIL.n560 0.388379
R828 VTAIL.n596 VTAIL.n595 0.388379
R829 VTAIL.n44 VTAIL.n14 0.388379
R830 VTAIL.n50 VTAIL.n49 0.388379
R831 VTAIL.n122 VTAIL.n92 0.388379
R832 VTAIL.n128 VTAIL.n127 0.388379
R833 VTAIL.n200 VTAIL.n170 0.388379
R834 VTAIL.n206 VTAIL.n205 0.388379
R835 VTAIL.n518 VTAIL.n517 0.388379
R836 VTAIL.n484 VTAIL.n482 0.388379
R837 VTAIL.n440 VTAIL.n439 0.388379
R838 VTAIL.n406 VTAIL.n404 0.388379
R839 VTAIL.n362 VTAIL.n361 0.388379
R840 VTAIL.n328 VTAIL.n326 0.388379
R841 VTAIL.n284 VTAIL.n283 0.388379
R842 VTAIL.n250 VTAIL.n248 0.388379
R843 VTAIL.n572 VTAIL.n567 0.155672
R844 VTAIL.n579 VTAIL.n567 0.155672
R845 VTAIL.n580 VTAIL.n579 0.155672
R846 VTAIL.n580 VTAIL.n563 0.155672
R847 VTAIL.n587 VTAIL.n563 0.155672
R848 VTAIL.n588 VTAIL.n587 0.155672
R849 VTAIL.n588 VTAIL.n559 0.155672
R850 VTAIL.n597 VTAIL.n559 0.155672
R851 VTAIL.n598 VTAIL.n597 0.155672
R852 VTAIL.n598 VTAIL.n555 0.155672
R853 VTAIL.n605 VTAIL.n555 0.155672
R854 VTAIL.n606 VTAIL.n605 0.155672
R855 VTAIL.n606 VTAIL.n551 0.155672
R856 VTAIL.n613 VTAIL.n551 0.155672
R857 VTAIL.n614 VTAIL.n613 0.155672
R858 VTAIL.n614 VTAIL.n547 0.155672
R859 VTAIL.n621 VTAIL.n547 0.155672
R860 VTAIL.n26 VTAIL.n21 0.155672
R861 VTAIL.n33 VTAIL.n21 0.155672
R862 VTAIL.n34 VTAIL.n33 0.155672
R863 VTAIL.n34 VTAIL.n17 0.155672
R864 VTAIL.n41 VTAIL.n17 0.155672
R865 VTAIL.n42 VTAIL.n41 0.155672
R866 VTAIL.n42 VTAIL.n13 0.155672
R867 VTAIL.n51 VTAIL.n13 0.155672
R868 VTAIL.n52 VTAIL.n51 0.155672
R869 VTAIL.n52 VTAIL.n9 0.155672
R870 VTAIL.n59 VTAIL.n9 0.155672
R871 VTAIL.n60 VTAIL.n59 0.155672
R872 VTAIL.n60 VTAIL.n5 0.155672
R873 VTAIL.n67 VTAIL.n5 0.155672
R874 VTAIL.n68 VTAIL.n67 0.155672
R875 VTAIL.n68 VTAIL.n1 0.155672
R876 VTAIL.n75 VTAIL.n1 0.155672
R877 VTAIL.n104 VTAIL.n99 0.155672
R878 VTAIL.n111 VTAIL.n99 0.155672
R879 VTAIL.n112 VTAIL.n111 0.155672
R880 VTAIL.n112 VTAIL.n95 0.155672
R881 VTAIL.n119 VTAIL.n95 0.155672
R882 VTAIL.n120 VTAIL.n119 0.155672
R883 VTAIL.n120 VTAIL.n91 0.155672
R884 VTAIL.n129 VTAIL.n91 0.155672
R885 VTAIL.n130 VTAIL.n129 0.155672
R886 VTAIL.n130 VTAIL.n87 0.155672
R887 VTAIL.n137 VTAIL.n87 0.155672
R888 VTAIL.n138 VTAIL.n137 0.155672
R889 VTAIL.n138 VTAIL.n83 0.155672
R890 VTAIL.n145 VTAIL.n83 0.155672
R891 VTAIL.n146 VTAIL.n145 0.155672
R892 VTAIL.n146 VTAIL.n79 0.155672
R893 VTAIL.n153 VTAIL.n79 0.155672
R894 VTAIL.n182 VTAIL.n177 0.155672
R895 VTAIL.n189 VTAIL.n177 0.155672
R896 VTAIL.n190 VTAIL.n189 0.155672
R897 VTAIL.n190 VTAIL.n173 0.155672
R898 VTAIL.n197 VTAIL.n173 0.155672
R899 VTAIL.n198 VTAIL.n197 0.155672
R900 VTAIL.n198 VTAIL.n169 0.155672
R901 VTAIL.n207 VTAIL.n169 0.155672
R902 VTAIL.n208 VTAIL.n207 0.155672
R903 VTAIL.n208 VTAIL.n165 0.155672
R904 VTAIL.n215 VTAIL.n165 0.155672
R905 VTAIL.n216 VTAIL.n215 0.155672
R906 VTAIL.n216 VTAIL.n161 0.155672
R907 VTAIL.n223 VTAIL.n161 0.155672
R908 VTAIL.n224 VTAIL.n223 0.155672
R909 VTAIL.n224 VTAIL.n157 0.155672
R910 VTAIL.n231 VTAIL.n157 0.155672
R911 VTAIL.n543 VTAIL.n469 0.155672
R912 VTAIL.n536 VTAIL.n469 0.155672
R913 VTAIL.n536 VTAIL.n535 0.155672
R914 VTAIL.n535 VTAIL.n473 0.155672
R915 VTAIL.n528 VTAIL.n473 0.155672
R916 VTAIL.n528 VTAIL.n527 0.155672
R917 VTAIL.n527 VTAIL.n477 0.155672
R918 VTAIL.n520 VTAIL.n477 0.155672
R919 VTAIL.n520 VTAIL.n519 0.155672
R920 VTAIL.n519 VTAIL.n481 0.155672
R921 VTAIL.n511 VTAIL.n481 0.155672
R922 VTAIL.n511 VTAIL.n510 0.155672
R923 VTAIL.n510 VTAIL.n486 0.155672
R924 VTAIL.n503 VTAIL.n486 0.155672
R925 VTAIL.n503 VTAIL.n502 0.155672
R926 VTAIL.n502 VTAIL.n490 0.155672
R927 VTAIL.n495 VTAIL.n490 0.155672
R928 VTAIL.n465 VTAIL.n391 0.155672
R929 VTAIL.n458 VTAIL.n391 0.155672
R930 VTAIL.n458 VTAIL.n457 0.155672
R931 VTAIL.n457 VTAIL.n395 0.155672
R932 VTAIL.n450 VTAIL.n395 0.155672
R933 VTAIL.n450 VTAIL.n449 0.155672
R934 VTAIL.n449 VTAIL.n399 0.155672
R935 VTAIL.n442 VTAIL.n399 0.155672
R936 VTAIL.n442 VTAIL.n441 0.155672
R937 VTAIL.n441 VTAIL.n403 0.155672
R938 VTAIL.n433 VTAIL.n403 0.155672
R939 VTAIL.n433 VTAIL.n432 0.155672
R940 VTAIL.n432 VTAIL.n408 0.155672
R941 VTAIL.n425 VTAIL.n408 0.155672
R942 VTAIL.n425 VTAIL.n424 0.155672
R943 VTAIL.n424 VTAIL.n412 0.155672
R944 VTAIL.n417 VTAIL.n412 0.155672
R945 VTAIL.n387 VTAIL.n313 0.155672
R946 VTAIL.n380 VTAIL.n313 0.155672
R947 VTAIL.n380 VTAIL.n379 0.155672
R948 VTAIL.n379 VTAIL.n317 0.155672
R949 VTAIL.n372 VTAIL.n317 0.155672
R950 VTAIL.n372 VTAIL.n371 0.155672
R951 VTAIL.n371 VTAIL.n321 0.155672
R952 VTAIL.n364 VTAIL.n321 0.155672
R953 VTAIL.n364 VTAIL.n363 0.155672
R954 VTAIL.n363 VTAIL.n325 0.155672
R955 VTAIL.n355 VTAIL.n325 0.155672
R956 VTAIL.n355 VTAIL.n354 0.155672
R957 VTAIL.n354 VTAIL.n330 0.155672
R958 VTAIL.n347 VTAIL.n330 0.155672
R959 VTAIL.n347 VTAIL.n346 0.155672
R960 VTAIL.n346 VTAIL.n334 0.155672
R961 VTAIL.n339 VTAIL.n334 0.155672
R962 VTAIL.n309 VTAIL.n235 0.155672
R963 VTAIL.n302 VTAIL.n235 0.155672
R964 VTAIL.n302 VTAIL.n301 0.155672
R965 VTAIL.n301 VTAIL.n239 0.155672
R966 VTAIL.n294 VTAIL.n239 0.155672
R967 VTAIL.n294 VTAIL.n293 0.155672
R968 VTAIL.n293 VTAIL.n243 0.155672
R969 VTAIL.n286 VTAIL.n243 0.155672
R970 VTAIL.n286 VTAIL.n285 0.155672
R971 VTAIL.n285 VTAIL.n247 0.155672
R972 VTAIL.n277 VTAIL.n247 0.155672
R973 VTAIL.n277 VTAIL.n276 0.155672
R974 VTAIL.n276 VTAIL.n252 0.155672
R975 VTAIL.n269 VTAIL.n252 0.155672
R976 VTAIL.n269 VTAIL.n268 0.155672
R977 VTAIL.n268 VTAIL.n256 0.155672
R978 VTAIL.n261 VTAIL.n256 0.155672
R979 B.n807 B.n806 585
R980 B.n330 B.n115 585
R981 B.n329 B.n328 585
R982 B.n327 B.n326 585
R983 B.n325 B.n324 585
R984 B.n323 B.n322 585
R985 B.n321 B.n320 585
R986 B.n319 B.n318 585
R987 B.n317 B.n316 585
R988 B.n315 B.n314 585
R989 B.n313 B.n312 585
R990 B.n311 B.n310 585
R991 B.n309 B.n308 585
R992 B.n307 B.n306 585
R993 B.n305 B.n304 585
R994 B.n303 B.n302 585
R995 B.n301 B.n300 585
R996 B.n299 B.n298 585
R997 B.n297 B.n296 585
R998 B.n295 B.n294 585
R999 B.n293 B.n292 585
R1000 B.n291 B.n290 585
R1001 B.n289 B.n288 585
R1002 B.n287 B.n286 585
R1003 B.n285 B.n284 585
R1004 B.n283 B.n282 585
R1005 B.n281 B.n280 585
R1006 B.n279 B.n278 585
R1007 B.n277 B.n276 585
R1008 B.n275 B.n274 585
R1009 B.n273 B.n272 585
R1010 B.n271 B.n270 585
R1011 B.n269 B.n268 585
R1012 B.n267 B.n266 585
R1013 B.n265 B.n264 585
R1014 B.n263 B.n262 585
R1015 B.n261 B.n260 585
R1016 B.n259 B.n258 585
R1017 B.n257 B.n256 585
R1018 B.n255 B.n254 585
R1019 B.n253 B.n252 585
R1020 B.n251 B.n250 585
R1021 B.n249 B.n248 585
R1022 B.n247 B.n246 585
R1023 B.n245 B.n244 585
R1024 B.n243 B.n242 585
R1025 B.n241 B.n240 585
R1026 B.n239 B.n238 585
R1027 B.n237 B.n236 585
R1028 B.n235 B.n234 585
R1029 B.n233 B.n232 585
R1030 B.n231 B.n230 585
R1031 B.n229 B.n228 585
R1032 B.n227 B.n226 585
R1033 B.n225 B.n224 585
R1034 B.n223 B.n222 585
R1035 B.n221 B.n220 585
R1036 B.n219 B.n218 585
R1037 B.n217 B.n216 585
R1038 B.n215 B.n214 585
R1039 B.n213 B.n212 585
R1040 B.n211 B.n210 585
R1041 B.n209 B.n208 585
R1042 B.n207 B.n206 585
R1043 B.n205 B.n204 585
R1044 B.n203 B.n202 585
R1045 B.n201 B.n200 585
R1046 B.n199 B.n198 585
R1047 B.n197 B.n196 585
R1048 B.n195 B.n194 585
R1049 B.n193 B.n192 585
R1050 B.n191 B.n190 585
R1051 B.n189 B.n188 585
R1052 B.n187 B.n186 585
R1053 B.n185 B.n184 585
R1054 B.n183 B.n182 585
R1055 B.n181 B.n180 585
R1056 B.n179 B.n178 585
R1057 B.n177 B.n176 585
R1058 B.n175 B.n174 585
R1059 B.n173 B.n172 585
R1060 B.n171 B.n170 585
R1061 B.n169 B.n168 585
R1062 B.n167 B.n166 585
R1063 B.n165 B.n164 585
R1064 B.n163 B.n162 585
R1065 B.n161 B.n160 585
R1066 B.n159 B.n158 585
R1067 B.n157 B.n156 585
R1068 B.n155 B.n154 585
R1069 B.n153 B.n152 585
R1070 B.n151 B.n150 585
R1071 B.n149 B.n148 585
R1072 B.n147 B.n146 585
R1073 B.n145 B.n144 585
R1074 B.n143 B.n142 585
R1075 B.n141 B.n140 585
R1076 B.n139 B.n138 585
R1077 B.n137 B.n136 585
R1078 B.n135 B.n134 585
R1079 B.n133 B.n132 585
R1080 B.n131 B.n130 585
R1081 B.n129 B.n128 585
R1082 B.n127 B.n126 585
R1083 B.n125 B.n124 585
R1084 B.n123 B.n122 585
R1085 B.n805 B.n62 585
R1086 B.n810 B.n62 585
R1087 B.n804 B.n61 585
R1088 B.n811 B.n61 585
R1089 B.n803 B.n802 585
R1090 B.n802 B.n57 585
R1091 B.n801 B.n56 585
R1092 B.n817 B.n56 585
R1093 B.n800 B.n55 585
R1094 B.n818 B.n55 585
R1095 B.n799 B.n54 585
R1096 B.n819 B.n54 585
R1097 B.n798 B.n797 585
R1098 B.n797 B.n50 585
R1099 B.n796 B.n49 585
R1100 B.n825 B.n49 585
R1101 B.n795 B.n48 585
R1102 B.n826 B.n48 585
R1103 B.n794 B.n47 585
R1104 B.n827 B.n47 585
R1105 B.n793 B.n792 585
R1106 B.n792 B.n43 585
R1107 B.n791 B.n42 585
R1108 B.n833 B.n42 585
R1109 B.n790 B.n41 585
R1110 B.n834 B.n41 585
R1111 B.n789 B.n40 585
R1112 B.n835 B.n40 585
R1113 B.n788 B.n787 585
R1114 B.n787 B.n36 585
R1115 B.n786 B.n35 585
R1116 B.n841 B.n35 585
R1117 B.n785 B.n34 585
R1118 B.n842 B.n34 585
R1119 B.n784 B.n33 585
R1120 B.n843 B.n33 585
R1121 B.n783 B.n782 585
R1122 B.n782 B.n32 585
R1123 B.n781 B.n28 585
R1124 B.n849 B.n28 585
R1125 B.n780 B.n27 585
R1126 B.n850 B.n27 585
R1127 B.n779 B.n26 585
R1128 B.n851 B.n26 585
R1129 B.n778 B.n777 585
R1130 B.n777 B.n22 585
R1131 B.n776 B.n21 585
R1132 B.n857 B.n21 585
R1133 B.n775 B.n20 585
R1134 B.n858 B.n20 585
R1135 B.n774 B.n19 585
R1136 B.n859 B.n19 585
R1137 B.n773 B.n772 585
R1138 B.n772 B.n15 585
R1139 B.n771 B.n14 585
R1140 B.n865 B.n14 585
R1141 B.n770 B.n13 585
R1142 B.n866 B.n13 585
R1143 B.n769 B.n12 585
R1144 B.n867 B.n12 585
R1145 B.n768 B.n767 585
R1146 B.n767 B.n8 585
R1147 B.n766 B.n7 585
R1148 B.n873 B.n7 585
R1149 B.n765 B.n6 585
R1150 B.n874 B.n6 585
R1151 B.n764 B.n5 585
R1152 B.n875 B.n5 585
R1153 B.n763 B.n762 585
R1154 B.n762 B.n4 585
R1155 B.n761 B.n331 585
R1156 B.n761 B.n760 585
R1157 B.n751 B.n332 585
R1158 B.n333 B.n332 585
R1159 B.n753 B.n752 585
R1160 B.n754 B.n753 585
R1161 B.n750 B.n338 585
R1162 B.n338 B.n337 585
R1163 B.n749 B.n748 585
R1164 B.n748 B.n747 585
R1165 B.n340 B.n339 585
R1166 B.n341 B.n340 585
R1167 B.n740 B.n739 585
R1168 B.n741 B.n740 585
R1169 B.n738 B.n346 585
R1170 B.n346 B.n345 585
R1171 B.n737 B.n736 585
R1172 B.n736 B.n735 585
R1173 B.n348 B.n347 585
R1174 B.n349 B.n348 585
R1175 B.n728 B.n727 585
R1176 B.n729 B.n728 585
R1177 B.n726 B.n354 585
R1178 B.n354 B.n353 585
R1179 B.n725 B.n724 585
R1180 B.n724 B.n723 585
R1181 B.n356 B.n355 585
R1182 B.n716 B.n356 585
R1183 B.n715 B.n714 585
R1184 B.n717 B.n715 585
R1185 B.n713 B.n361 585
R1186 B.n361 B.n360 585
R1187 B.n712 B.n711 585
R1188 B.n711 B.n710 585
R1189 B.n363 B.n362 585
R1190 B.n364 B.n363 585
R1191 B.n703 B.n702 585
R1192 B.n704 B.n703 585
R1193 B.n701 B.n369 585
R1194 B.n369 B.n368 585
R1195 B.n700 B.n699 585
R1196 B.n699 B.n698 585
R1197 B.n371 B.n370 585
R1198 B.n372 B.n371 585
R1199 B.n691 B.n690 585
R1200 B.n692 B.n691 585
R1201 B.n689 B.n377 585
R1202 B.n377 B.n376 585
R1203 B.n688 B.n687 585
R1204 B.n687 B.n686 585
R1205 B.n379 B.n378 585
R1206 B.n380 B.n379 585
R1207 B.n679 B.n678 585
R1208 B.n680 B.n679 585
R1209 B.n677 B.n385 585
R1210 B.n385 B.n384 585
R1211 B.n676 B.n675 585
R1212 B.n675 B.n674 585
R1213 B.n387 B.n386 585
R1214 B.n388 B.n387 585
R1215 B.n667 B.n666 585
R1216 B.n668 B.n667 585
R1217 B.n665 B.n393 585
R1218 B.n393 B.n392 585
R1219 B.n660 B.n659 585
R1220 B.n658 B.n448 585
R1221 B.n657 B.n447 585
R1222 B.n662 B.n447 585
R1223 B.n656 B.n655 585
R1224 B.n654 B.n653 585
R1225 B.n652 B.n651 585
R1226 B.n650 B.n649 585
R1227 B.n648 B.n647 585
R1228 B.n646 B.n645 585
R1229 B.n644 B.n643 585
R1230 B.n642 B.n641 585
R1231 B.n640 B.n639 585
R1232 B.n638 B.n637 585
R1233 B.n636 B.n635 585
R1234 B.n634 B.n633 585
R1235 B.n632 B.n631 585
R1236 B.n630 B.n629 585
R1237 B.n628 B.n627 585
R1238 B.n626 B.n625 585
R1239 B.n624 B.n623 585
R1240 B.n622 B.n621 585
R1241 B.n620 B.n619 585
R1242 B.n618 B.n617 585
R1243 B.n616 B.n615 585
R1244 B.n614 B.n613 585
R1245 B.n612 B.n611 585
R1246 B.n610 B.n609 585
R1247 B.n608 B.n607 585
R1248 B.n606 B.n605 585
R1249 B.n604 B.n603 585
R1250 B.n602 B.n601 585
R1251 B.n600 B.n599 585
R1252 B.n598 B.n597 585
R1253 B.n596 B.n595 585
R1254 B.n594 B.n593 585
R1255 B.n592 B.n591 585
R1256 B.n590 B.n589 585
R1257 B.n588 B.n587 585
R1258 B.n586 B.n585 585
R1259 B.n584 B.n583 585
R1260 B.n582 B.n581 585
R1261 B.n580 B.n579 585
R1262 B.n578 B.n577 585
R1263 B.n576 B.n575 585
R1264 B.n574 B.n573 585
R1265 B.n572 B.n571 585
R1266 B.n570 B.n569 585
R1267 B.n568 B.n567 585
R1268 B.n565 B.n564 585
R1269 B.n563 B.n562 585
R1270 B.n561 B.n560 585
R1271 B.n559 B.n558 585
R1272 B.n557 B.n556 585
R1273 B.n555 B.n554 585
R1274 B.n553 B.n552 585
R1275 B.n551 B.n550 585
R1276 B.n549 B.n548 585
R1277 B.n547 B.n546 585
R1278 B.n544 B.n543 585
R1279 B.n542 B.n541 585
R1280 B.n540 B.n539 585
R1281 B.n538 B.n537 585
R1282 B.n536 B.n535 585
R1283 B.n534 B.n533 585
R1284 B.n532 B.n531 585
R1285 B.n530 B.n529 585
R1286 B.n528 B.n527 585
R1287 B.n526 B.n525 585
R1288 B.n524 B.n523 585
R1289 B.n522 B.n521 585
R1290 B.n520 B.n519 585
R1291 B.n518 B.n517 585
R1292 B.n516 B.n515 585
R1293 B.n514 B.n513 585
R1294 B.n512 B.n511 585
R1295 B.n510 B.n509 585
R1296 B.n508 B.n507 585
R1297 B.n506 B.n505 585
R1298 B.n504 B.n503 585
R1299 B.n502 B.n501 585
R1300 B.n500 B.n499 585
R1301 B.n498 B.n497 585
R1302 B.n496 B.n495 585
R1303 B.n494 B.n493 585
R1304 B.n492 B.n491 585
R1305 B.n490 B.n489 585
R1306 B.n488 B.n487 585
R1307 B.n486 B.n485 585
R1308 B.n484 B.n483 585
R1309 B.n482 B.n481 585
R1310 B.n480 B.n479 585
R1311 B.n478 B.n477 585
R1312 B.n476 B.n475 585
R1313 B.n474 B.n473 585
R1314 B.n472 B.n471 585
R1315 B.n470 B.n469 585
R1316 B.n468 B.n467 585
R1317 B.n466 B.n465 585
R1318 B.n464 B.n463 585
R1319 B.n462 B.n461 585
R1320 B.n460 B.n459 585
R1321 B.n458 B.n457 585
R1322 B.n456 B.n455 585
R1323 B.n454 B.n453 585
R1324 B.n395 B.n394 585
R1325 B.n664 B.n663 585
R1326 B.n663 B.n662 585
R1327 B.n391 B.n390 585
R1328 B.n392 B.n391 585
R1329 B.n670 B.n669 585
R1330 B.n669 B.n668 585
R1331 B.n671 B.n389 585
R1332 B.n389 B.n388 585
R1333 B.n673 B.n672 585
R1334 B.n674 B.n673 585
R1335 B.n383 B.n382 585
R1336 B.n384 B.n383 585
R1337 B.n682 B.n681 585
R1338 B.n681 B.n680 585
R1339 B.n683 B.n381 585
R1340 B.n381 B.n380 585
R1341 B.n685 B.n684 585
R1342 B.n686 B.n685 585
R1343 B.n375 B.n374 585
R1344 B.n376 B.n375 585
R1345 B.n694 B.n693 585
R1346 B.n693 B.n692 585
R1347 B.n695 B.n373 585
R1348 B.n373 B.n372 585
R1349 B.n697 B.n696 585
R1350 B.n698 B.n697 585
R1351 B.n367 B.n366 585
R1352 B.n368 B.n367 585
R1353 B.n706 B.n705 585
R1354 B.n705 B.n704 585
R1355 B.n707 B.n365 585
R1356 B.n365 B.n364 585
R1357 B.n709 B.n708 585
R1358 B.n710 B.n709 585
R1359 B.n359 B.n358 585
R1360 B.n360 B.n359 585
R1361 B.n719 B.n718 585
R1362 B.n718 B.n717 585
R1363 B.n720 B.n357 585
R1364 B.n716 B.n357 585
R1365 B.n722 B.n721 585
R1366 B.n723 B.n722 585
R1367 B.n352 B.n351 585
R1368 B.n353 B.n352 585
R1369 B.n731 B.n730 585
R1370 B.n730 B.n729 585
R1371 B.n732 B.n350 585
R1372 B.n350 B.n349 585
R1373 B.n734 B.n733 585
R1374 B.n735 B.n734 585
R1375 B.n344 B.n343 585
R1376 B.n345 B.n344 585
R1377 B.n743 B.n742 585
R1378 B.n742 B.n741 585
R1379 B.n744 B.n342 585
R1380 B.n342 B.n341 585
R1381 B.n746 B.n745 585
R1382 B.n747 B.n746 585
R1383 B.n336 B.n335 585
R1384 B.n337 B.n336 585
R1385 B.n756 B.n755 585
R1386 B.n755 B.n754 585
R1387 B.n757 B.n334 585
R1388 B.n334 B.n333 585
R1389 B.n759 B.n758 585
R1390 B.n760 B.n759 585
R1391 B.n2 B.n0 585
R1392 B.n4 B.n2 585
R1393 B.n3 B.n1 585
R1394 B.n874 B.n3 585
R1395 B.n872 B.n871 585
R1396 B.n873 B.n872 585
R1397 B.n870 B.n9 585
R1398 B.n9 B.n8 585
R1399 B.n869 B.n868 585
R1400 B.n868 B.n867 585
R1401 B.n11 B.n10 585
R1402 B.n866 B.n11 585
R1403 B.n864 B.n863 585
R1404 B.n865 B.n864 585
R1405 B.n862 B.n16 585
R1406 B.n16 B.n15 585
R1407 B.n861 B.n860 585
R1408 B.n860 B.n859 585
R1409 B.n18 B.n17 585
R1410 B.n858 B.n18 585
R1411 B.n856 B.n855 585
R1412 B.n857 B.n856 585
R1413 B.n854 B.n23 585
R1414 B.n23 B.n22 585
R1415 B.n853 B.n852 585
R1416 B.n852 B.n851 585
R1417 B.n25 B.n24 585
R1418 B.n850 B.n25 585
R1419 B.n848 B.n847 585
R1420 B.n849 B.n848 585
R1421 B.n846 B.n29 585
R1422 B.n32 B.n29 585
R1423 B.n845 B.n844 585
R1424 B.n844 B.n843 585
R1425 B.n31 B.n30 585
R1426 B.n842 B.n31 585
R1427 B.n840 B.n839 585
R1428 B.n841 B.n840 585
R1429 B.n838 B.n37 585
R1430 B.n37 B.n36 585
R1431 B.n837 B.n836 585
R1432 B.n836 B.n835 585
R1433 B.n39 B.n38 585
R1434 B.n834 B.n39 585
R1435 B.n832 B.n831 585
R1436 B.n833 B.n832 585
R1437 B.n830 B.n44 585
R1438 B.n44 B.n43 585
R1439 B.n829 B.n828 585
R1440 B.n828 B.n827 585
R1441 B.n46 B.n45 585
R1442 B.n826 B.n46 585
R1443 B.n824 B.n823 585
R1444 B.n825 B.n824 585
R1445 B.n822 B.n51 585
R1446 B.n51 B.n50 585
R1447 B.n821 B.n820 585
R1448 B.n820 B.n819 585
R1449 B.n53 B.n52 585
R1450 B.n818 B.n53 585
R1451 B.n816 B.n815 585
R1452 B.n817 B.n816 585
R1453 B.n814 B.n58 585
R1454 B.n58 B.n57 585
R1455 B.n813 B.n812 585
R1456 B.n812 B.n811 585
R1457 B.n60 B.n59 585
R1458 B.n810 B.n60 585
R1459 B.n877 B.n876 585
R1460 B.n876 B.n875 585
R1461 B.n660 B.n391 468.476
R1462 B.n122 B.n60 468.476
R1463 B.n663 B.n393 468.476
R1464 B.n807 B.n62 468.476
R1465 B.n451 B.t14 374.551
R1466 B.n116 B.t16 374.551
R1467 B.n449 B.t7 374.551
R1468 B.n119 B.t10 374.551
R1469 B.n451 B.t12 345.12
R1470 B.n449 B.t4 345.12
R1471 B.n119 B.t8 345.12
R1472 B.n116 B.t15 345.12
R1473 B.n452 B.t13 319.861
R1474 B.n117 B.t17 319.861
R1475 B.n450 B.t6 319.861
R1476 B.n120 B.t11 319.861
R1477 B.n809 B.n808 256.663
R1478 B.n809 B.n114 256.663
R1479 B.n809 B.n113 256.663
R1480 B.n809 B.n112 256.663
R1481 B.n809 B.n111 256.663
R1482 B.n809 B.n110 256.663
R1483 B.n809 B.n109 256.663
R1484 B.n809 B.n108 256.663
R1485 B.n809 B.n107 256.663
R1486 B.n809 B.n106 256.663
R1487 B.n809 B.n105 256.663
R1488 B.n809 B.n104 256.663
R1489 B.n809 B.n103 256.663
R1490 B.n809 B.n102 256.663
R1491 B.n809 B.n101 256.663
R1492 B.n809 B.n100 256.663
R1493 B.n809 B.n99 256.663
R1494 B.n809 B.n98 256.663
R1495 B.n809 B.n97 256.663
R1496 B.n809 B.n96 256.663
R1497 B.n809 B.n95 256.663
R1498 B.n809 B.n94 256.663
R1499 B.n809 B.n93 256.663
R1500 B.n809 B.n92 256.663
R1501 B.n809 B.n91 256.663
R1502 B.n809 B.n90 256.663
R1503 B.n809 B.n89 256.663
R1504 B.n809 B.n88 256.663
R1505 B.n809 B.n87 256.663
R1506 B.n809 B.n86 256.663
R1507 B.n809 B.n85 256.663
R1508 B.n809 B.n84 256.663
R1509 B.n809 B.n83 256.663
R1510 B.n809 B.n82 256.663
R1511 B.n809 B.n81 256.663
R1512 B.n809 B.n80 256.663
R1513 B.n809 B.n79 256.663
R1514 B.n809 B.n78 256.663
R1515 B.n809 B.n77 256.663
R1516 B.n809 B.n76 256.663
R1517 B.n809 B.n75 256.663
R1518 B.n809 B.n74 256.663
R1519 B.n809 B.n73 256.663
R1520 B.n809 B.n72 256.663
R1521 B.n809 B.n71 256.663
R1522 B.n809 B.n70 256.663
R1523 B.n809 B.n69 256.663
R1524 B.n809 B.n68 256.663
R1525 B.n809 B.n67 256.663
R1526 B.n809 B.n66 256.663
R1527 B.n809 B.n65 256.663
R1528 B.n809 B.n64 256.663
R1529 B.n809 B.n63 256.663
R1530 B.n662 B.n661 256.663
R1531 B.n662 B.n396 256.663
R1532 B.n662 B.n397 256.663
R1533 B.n662 B.n398 256.663
R1534 B.n662 B.n399 256.663
R1535 B.n662 B.n400 256.663
R1536 B.n662 B.n401 256.663
R1537 B.n662 B.n402 256.663
R1538 B.n662 B.n403 256.663
R1539 B.n662 B.n404 256.663
R1540 B.n662 B.n405 256.663
R1541 B.n662 B.n406 256.663
R1542 B.n662 B.n407 256.663
R1543 B.n662 B.n408 256.663
R1544 B.n662 B.n409 256.663
R1545 B.n662 B.n410 256.663
R1546 B.n662 B.n411 256.663
R1547 B.n662 B.n412 256.663
R1548 B.n662 B.n413 256.663
R1549 B.n662 B.n414 256.663
R1550 B.n662 B.n415 256.663
R1551 B.n662 B.n416 256.663
R1552 B.n662 B.n417 256.663
R1553 B.n662 B.n418 256.663
R1554 B.n662 B.n419 256.663
R1555 B.n662 B.n420 256.663
R1556 B.n662 B.n421 256.663
R1557 B.n662 B.n422 256.663
R1558 B.n662 B.n423 256.663
R1559 B.n662 B.n424 256.663
R1560 B.n662 B.n425 256.663
R1561 B.n662 B.n426 256.663
R1562 B.n662 B.n427 256.663
R1563 B.n662 B.n428 256.663
R1564 B.n662 B.n429 256.663
R1565 B.n662 B.n430 256.663
R1566 B.n662 B.n431 256.663
R1567 B.n662 B.n432 256.663
R1568 B.n662 B.n433 256.663
R1569 B.n662 B.n434 256.663
R1570 B.n662 B.n435 256.663
R1571 B.n662 B.n436 256.663
R1572 B.n662 B.n437 256.663
R1573 B.n662 B.n438 256.663
R1574 B.n662 B.n439 256.663
R1575 B.n662 B.n440 256.663
R1576 B.n662 B.n441 256.663
R1577 B.n662 B.n442 256.663
R1578 B.n662 B.n443 256.663
R1579 B.n662 B.n444 256.663
R1580 B.n662 B.n445 256.663
R1581 B.n662 B.n446 256.663
R1582 B.n669 B.n391 163.367
R1583 B.n669 B.n389 163.367
R1584 B.n673 B.n389 163.367
R1585 B.n673 B.n383 163.367
R1586 B.n681 B.n383 163.367
R1587 B.n681 B.n381 163.367
R1588 B.n685 B.n381 163.367
R1589 B.n685 B.n375 163.367
R1590 B.n693 B.n375 163.367
R1591 B.n693 B.n373 163.367
R1592 B.n697 B.n373 163.367
R1593 B.n697 B.n367 163.367
R1594 B.n705 B.n367 163.367
R1595 B.n705 B.n365 163.367
R1596 B.n709 B.n365 163.367
R1597 B.n709 B.n359 163.367
R1598 B.n718 B.n359 163.367
R1599 B.n718 B.n357 163.367
R1600 B.n722 B.n357 163.367
R1601 B.n722 B.n352 163.367
R1602 B.n730 B.n352 163.367
R1603 B.n730 B.n350 163.367
R1604 B.n734 B.n350 163.367
R1605 B.n734 B.n344 163.367
R1606 B.n742 B.n344 163.367
R1607 B.n742 B.n342 163.367
R1608 B.n746 B.n342 163.367
R1609 B.n746 B.n336 163.367
R1610 B.n755 B.n336 163.367
R1611 B.n755 B.n334 163.367
R1612 B.n759 B.n334 163.367
R1613 B.n759 B.n2 163.367
R1614 B.n876 B.n2 163.367
R1615 B.n876 B.n3 163.367
R1616 B.n872 B.n3 163.367
R1617 B.n872 B.n9 163.367
R1618 B.n868 B.n9 163.367
R1619 B.n868 B.n11 163.367
R1620 B.n864 B.n11 163.367
R1621 B.n864 B.n16 163.367
R1622 B.n860 B.n16 163.367
R1623 B.n860 B.n18 163.367
R1624 B.n856 B.n18 163.367
R1625 B.n856 B.n23 163.367
R1626 B.n852 B.n23 163.367
R1627 B.n852 B.n25 163.367
R1628 B.n848 B.n25 163.367
R1629 B.n848 B.n29 163.367
R1630 B.n844 B.n29 163.367
R1631 B.n844 B.n31 163.367
R1632 B.n840 B.n31 163.367
R1633 B.n840 B.n37 163.367
R1634 B.n836 B.n37 163.367
R1635 B.n836 B.n39 163.367
R1636 B.n832 B.n39 163.367
R1637 B.n832 B.n44 163.367
R1638 B.n828 B.n44 163.367
R1639 B.n828 B.n46 163.367
R1640 B.n824 B.n46 163.367
R1641 B.n824 B.n51 163.367
R1642 B.n820 B.n51 163.367
R1643 B.n820 B.n53 163.367
R1644 B.n816 B.n53 163.367
R1645 B.n816 B.n58 163.367
R1646 B.n812 B.n58 163.367
R1647 B.n812 B.n60 163.367
R1648 B.n448 B.n447 163.367
R1649 B.n655 B.n447 163.367
R1650 B.n653 B.n652 163.367
R1651 B.n649 B.n648 163.367
R1652 B.n645 B.n644 163.367
R1653 B.n641 B.n640 163.367
R1654 B.n637 B.n636 163.367
R1655 B.n633 B.n632 163.367
R1656 B.n629 B.n628 163.367
R1657 B.n625 B.n624 163.367
R1658 B.n621 B.n620 163.367
R1659 B.n617 B.n616 163.367
R1660 B.n613 B.n612 163.367
R1661 B.n609 B.n608 163.367
R1662 B.n605 B.n604 163.367
R1663 B.n601 B.n600 163.367
R1664 B.n597 B.n596 163.367
R1665 B.n593 B.n592 163.367
R1666 B.n589 B.n588 163.367
R1667 B.n585 B.n584 163.367
R1668 B.n581 B.n580 163.367
R1669 B.n577 B.n576 163.367
R1670 B.n573 B.n572 163.367
R1671 B.n569 B.n568 163.367
R1672 B.n564 B.n563 163.367
R1673 B.n560 B.n559 163.367
R1674 B.n556 B.n555 163.367
R1675 B.n552 B.n551 163.367
R1676 B.n548 B.n547 163.367
R1677 B.n543 B.n542 163.367
R1678 B.n539 B.n538 163.367
R1679 B.n535 B.n534 163.367
R1680 B.n531 B.n530 163.367
R1681 B.n527 B.n526 163.367
R1682 B.n523 B.n522 163.367
R1683 B.n519 B.n518 163.367
R1684 B.n515 B.n514 163.367
R1685 B.n511 B.n510 163.367
R1686 B.n507 B.n506 163.367
R1687 B.n503 B.n502 163.367
R1688 B.n499 B.n498 163.367
R1689 B.n495 B.n494 163.367
R1690 B.n491 B.n490 163.367
R1691 B.n487 B.n486 163.367
R1692 B.n483 B.n482 163.367
R1693 B.n479 B.n478 163.367
R1694 B.n475 B.n474 163.367
R1695 B.n471 B.n470 163.367
R1696 B.n467 B.n466 163.367
R1697 B.n463 B.n462 163.367
R1698 B.n459 B.n458 163.367
R1699 B.n455 B.n454 163.367
R1700 B.n663 B.n395 163.367
R1701 B.n667 B.n393 163.367
R1702 B.n667 B.n387 163.367
R1703 B.n675 B.n387 163.367
R1704 B.n675 B.n385 163.367
R1705 B.n679 B.n385 163.367
R1706 B.n679 B.n379 163.367
R1707 B.n687 B.n379 163.367
R1708 B.n687 B.n377 163.367
R1709 B.n691 B.n377 163.367
R1710 B.n691 B.n371 163.367
R1711 B.n699 B.n371 163.367
R1712 B.n699 B.n369 163.367
R1713 B.n703 B.n369 163.367
R1714 B.n703 B.n363 163.367
R1715 B.n711 B.n363 163.367
R1716 B.n711 B.n361 163.367
R1717 B.n715 B.n361 163.367
R1718 B.n715 B.n356 163.367
R1719 B.n724 B.n356 163.367
R1720 B.n724 B.n354 163.367
R1721 B.n728 B.n354 163.367
R1722 B.n728 B.n348 163.367
R1723 B.n736 B.n348 163.367
R1724 B.n736 B.n346 163.367
R1725 B.n740 B.n346 163.367
R1726 B.n740 B.n340 163.367
R1727 B.n748 B.n340 163.367
R1728 B.n748 B.n338 163.367
R1729 B.n753 B.n338 163.367
R1730 B.n753 B.n332 163.367
R1731 B.n761 B.n332 163.367
R1732 B.n762 B.n761 163.367
R1733 B.n762 B.n5 163.367
R1734 B.n6 B.n5 163.367
R1735 B.n7 B.n6 163.367
R1736 B.n767 B.n7 163.367
R1737 B.n767 B.n12 163.367
R1738 B.n13 B.n12 163.367
R1739 B.n14 B.n13 163.367
R1740 B.n772 B.n14 163.367
R1741 B.n772 B.n19 163.367
R1742 B.n20 B.n19 163.367
R1743 B.n21 B.n20 163.367
R1744 B.n777 B.n21 163.367
R1745 B.n777 B.n26 163.367
R1746 B.n27 B.n26 163.367
R1747 B.n28 B.n27 163.367
R1748 B.n782 B.n28 163.367
R1749 B.n782 B.n33 163.367
R1750 B.n34 B.n33 163.367
R1751 B.n35 B.n34 163.367
R1752 B.n787 B.n35 163.367
R1753 B.n787 B.n40 163.367
R1754 B.n41 B.n40 163.367
R1755 B.n42 B.n41 163.367
R1756 B.n792 B.n42 163.367
R1757 B.n792 B.n47 163.367
R1758 B.n48 B.n47 163.367
R1759 B.n49 B.n48 163.367
R1760 B.n797 B.n49 163.367
R1761 B.n797 B.n54 163.367
R1762 B.n55 B.n54 163.367
R1763 B.n56 B.n55 163.367
R1764 B.n802 B.n56 163.367
R1765 B.n802 B.n61 163.367
R1766 B.n62 B.n61 163.367
R1767 B.n126 B.n125 163.367
R1768 B.n130 B.n129 163.367
R1769 B.n134 B.n133 163.367
R1770 B.n138 B.n137 163.367
R1771 B.n142 B.n141 163.367
R1772 B.n146 B.n145 163.367
R1773 B.n150 B.n149 163.367
R1774 B.n154 B.n153 163.367
R1775 B.n158 B.n157 163.367
R1776 B.n162 B.n161 163.367
R1777 B.n166 B.n165 163.367
R1778 B.n170 B.n169 163.367
R1779 B.n174 B.n173 163.367
R1780 B.n178 B.n177 163.367
R1781 B.n182 B.n181 163.367
R1782 B.n186 B.n185 163.367
R1783 B.n190 B.n189 163.367
R1784 B.n194 B.n193 163.367
R1785 B.n198 B.n197 163.367
R1786 B.n202 B.n201 163.367
R1787 B.n206 B.n205 163.367
R1788 B.n210 B.n209 163.367
R1789 B.n214 B.n213 163.367
R1790 B.n218 B.n217 163.367
R1791 B.n222 B.n221 163.367
R1792 B.n226 B.n225 163.367
R1793 B.n230 B.n229 163.367
R1794 B.n234 B.n233 163.367
R1795 B.n238 B.n237 163.367
R1796 B.n242 B.n241 163.367
R1797 B.n246 B.n245 163.367
R1798 B.n250 B.n249 163.367
R1799 B.n254 B.n253 163.367
R1800 B.n258 B.n257 163.367
R1801 B.n262 B.n261 163.367
R1802 B.n266 B.n265 163.367
R1803 B.n270 B.n269 163.367
R1804 B.n274 B.n273 163.367
R1805 B.n278 B.n277 163.367
R1806 B.n282 B.n281 163.367
R1807 B.n286 B.n285 163.367
R1808 B.n290 B.n289 163.367
R1809 B.n294 B.n293 163.367
R1810 B.n298 B.n297 163.367
R1811 B.n302 B.n301 163.367
R1812 B.n306 B.n305 163.367
R1813 B.n310 B.n309 163.367
R1814 B.n314 B.n313 163.367
R1815 B.n318 B.n317 163.367
R1816 B.n322 B.n321 163.367
R1817 B.n326 B.n325 163.367
R1818 B.n328 B.n115 163.367
R1819 B.n661 B.n660 71.676
R1820 B.n655 B.n396 71.676
R1821 B.n652 B.n397 71.676
R1822 B.n648 B.n398 71.676
R1823 B.n644 B.n399 71.676
R1824 B.n640 B.n400 71.676
R1825 B.n636 B.n401 71.676
R1826 B.n632 B.n402 71.676
R1827 B.n628 B.n403 71.676
R1828 B.n624 B.n404 71.676
R1829 B.n620 B.n405 71.676
R1830 B.n616 B.n406 71.676
R1831 B.n612 B.n407 71.676
R1832 B.n608 B.n408 71.676
R1833 B.n604 B.n409 71.676
R1834 B.n600 B.n410 71.676
R1835 B.n596 B.n411 71.676
R1836 B.n592 B.n412 71.676
R1837 B.n588 B.n413 71.676
R1838 B.n584 B.n414 71.676
R1839 B.n580 B.n415 71.676
R1840 B.n576 B.n416 71.676
R1841 B.n572 B.n417 71.676
R1842 B.n568 B.n418 71.676
R1843 B.n563 B.n419 71.676
R1844 B.n559 B.n420 71.676
R1845 B.n555 B.n421 71.676
R1846 B.n551 B.n422 71.676
R1847 B.n547 B.n423 71.676
R1848 B.n542 B.n424 71.676
R1849 B.n538 B.n425 71.676
R1850 B.n534 B.n426 71.676
R1851 B.n530 B.n427 71.676
R1852 B.n526 B.n428 71.676
R1853 B.n522 B.n429 71.676
R1854 B.n518 B.n430 71.676
R1855 B.n514 B.n431 71.676
R1856 B.n510 B.n432 71.676
R1857 B.n506 B.n433 71.676
R1858 B.n502 B.n434 71.676
R1859 B.n498 B.n435 71.676
R1860 B.n494 B.n436 71.676
R1861 B.n490 B.n437 71.676
R1862 B.n486 B.n438 71.676
R1863 B.n482 B.n439 71.676
R1864 B.n478 B.n440 71.676
R1865 B.n474 B.n441 71.676
R1866 B.n470 B.n442 71.676
R1867 B.n466 B.n443 71.676
R1868 B.n462 B.n444 71.676
R1869 B.n458 B.n445 71.676
R1870 B.n454 B.n446 71.676
R1871 B.n122 B.n63 71.676
R1872 B.n126 B.n64 71.676
R1873 B.n130 B.n65 71.676
R1874 B.n134 B.n66 71.676
R1875 B.n138 B.n67 71.676
R1876 B.n142 B.n68 71.676
R1877 B.n146 B.n69 71.676
R1878 B.n150 B.n70 71.676
R1879 B.n154 B.n71 71.676
R1880 B.n158 B.n72 71.676
R1881 B.n162 B.n73 71.676
R1882 B.n166 B.n74 71.676
R1883 B.n170 B.n75 71.676
R1884 B.n174 B.n76 71.676
R1885 B.n178 B.n77 71.676
R1886 B.n182 B.n78 71.676
R1887 B.n186 B.n79 71.676
R1888 B.n190 B.n80 71.676
R1889 B.n194 B.n81 71.676
R1890 B.n198 B.n82 71.676
R1891 B.n202 B.n83 71.676
R1892 B.n206 B.n84 71.676
R1893 B.n210 B.n85 71.676
R1894 B.n214 B.n86 71.676
R1895 B.n218 B.n87 71.676
R1896 B.n222 B.n88 71.676
R1897 B.n226 B.n89 71.676
R1898 B.n230 B.n90 71.676
R1899 B.n234 B.n91 71.676
R1900 B.n238 B.n92 71.676
R1901 B.n242 B.n93 71.676
R1902 B.n246 B.n94 71.676
R1903 B.n250 B.n95 71.676
R1904 B.n254 B.n96 71.676
R1905 B.n258 B.n97 71.676
R1906 B.n262 B.n98 71.676
R1907 B.n266 B.n99 71.676
R1908 B.n270 B.n100 71.676
R1909 B.n274 B.n101 71.676
R1910 B.n278 B.n102 71.676
R1911 B.n282 B.n103 71.676
R1912 B.n286 B.n104 71.676
R1913 B.n290 B.n105 71.676
R1914 B.n294 B.n106 71.676
R1915 B.n298 B.n107 71.676
R1916 B.n302 B.n108 71.676
R1917 B.n306 B.n109 71.676
R1918 B.n310 B.n110 71.676
R1919 B.n314 B.n111 71.676
R1920 B.n318 B.n112 71.676
R1921 B.n322 B.n113 71.676
R1922 B.n326 B.n114 71.676
R1923 B.n808 B.n115 71.676
R1924 B.n808 B.n807 71.676
R1925 B.n328 B.n114 71.676
R1926 B.n325 B.n113 71.676
R1927 B.n321 B.n112 71.676
R1928 B.n317 B.n111 71.676
R1929 B.n313 B.n110 71.676
R1930 B.n309 B.n109 71.676
R1931 B.n305 B.n108 71.676
R1932 B.n301 B.n107 71.676
R1933 B.n297 B.n106 71.676
R1934 B.n293 B.n105 71.676
R1935 B.n289 B.n104 71.676
R1936 B.n285 B.n103 71.676
R1937 B.n281 B.n102 71.676
R1938 B.n277 B.n101 71.676
R1939 B.n273 B.n100 71.676
R1940 B.n269 B.n99 71.676
R1941 B.n265 B.n98 71.676
R1942 B.n261 B.n97 71.676
R1943 B.n257 B.n96 71.676
R1944 B.n253 B.n95 71.676
R1945 B.n249 B.n94 71.676
R1946 B.n245 B.n93 71.676
R1947 B.n241 B.n92 71.676
R1948 B.n237 B.n91 71.676
R1949 B.n233 B.n90 71.676
R1950 B.n229 B.n89 71.676
R1951 B.n225 B.n88 71.676
R1952 B.n221 B.n87 71.676
R1953 B.n217 B.n86 71.676
R1954 B.n213 B.n85 71.676
R1955 B.n209 B.n84 71.676
R1956 B.n205 B.n83 71.676
R1957 B.n201 B.n82 71.676
R1958 B.n197 B.n81 71.676
R1959 B.n193 B.n80 71.676
R1960 B.n189 B.n79 71.676
R1961 B.n185 B.n78 71.676
R1962 B.n181 B.n77 71.676
R1963 B.n177 B.n76 71.676
R1964 B.n173 B.n75 71.676
R1965 B.n169 B.n74 71.676
R1966 B.n165 B.n73 71.676
R1967 B.n161 B.n72 71.676
R1968 B.n157 B.n71 71.676
R1969 B.n153 B.n70 71.676
R1970 B.n149 B.n69 71.676
R1971 B.n145 B.n68 71.676
R1972 B.n141 B.n67 71.676
R1973 B.n137 B.n66 71.676
R1974 B.n133 B.n65 71.676
R1975 B.n129 B.n64 71.676
R1976 B.n125 B.n63 71.676
R1977 B.n661 B.n448 71.676
R1978 B.n653 B.n396 71.676
R1979 B.n649 B.n397 71.676
R1980 B.n645 B.n398 71.676
R1981 B.n641 B.n399 71.676
R1982 B.n637 B.n400 71.676
R1983 B.n633 B.n401 71.676
R1984 B.n629 B.n402 71.676
R1985 B.n625 B.n403 71.676
R1986 B.n621 B.n404 71.676
R1987 B.n617 B.n405 71.676
R1988 B.n613 B.n406 71.676
R1989 B.n609 B.n407 71.676
R1990 B.n605 B.n408 71.676
R1991 B.n601 B.n409 71.676
R1992 B.n597 B.n410 71.676
R1993 B.n593 B.n411 71.676
R1994 B.n589 B.n412 71.676
R1995 B.n585 B.n413 71.676
R1996 B.n581 B.n414 71.676
R1997 B.n577 B.n415 71.676
R1998 B.n573 B.n416 71.676
R1999 B.n569 B.n417 71.676
R2000 B.n564 B.n418 71.676
R2001 B.n560 B.n419 71.676
R2002 B.n556 B.n420 71.676
R2003 B.n552 B.n421 71.676
R2004 B.n548 B.n422 71.676
R2005 B.n543 B.n423 71.676
R2006 B.n539 B.n424 71.676
R2007 B.n535 B.n425 71.676
R2008 B.n531 B.n426 71.676
R2009 B.n527 B.n427 71.676
R2010 B.n523 B.n428 71.676
R2011 B.n519 B.n429 71.676
R2012 B.n515 B.n430 71.676
R2013 B.n511 B.n431 71.676
R2014 B.n507 B.n432 71.676
R2015 B.n503 B.n433 71.676
R2016 B.n499 B.n434 71.676
R2017 B.n495 B.n435 71.676
R2018 B.n491 B.n436 71.676
R2019 B.n487 B.n437 71.676
R2020 B.n483 B.n438 71.676
R2021 B.n479 B.n439 71.676
R2022 B.n475 B.n440 71.676
R2023 B.n471 B.n441 71.676
R2024 B.n467 B.n442 71.676
R2025 B.n463 B.n443 71.676
R2026 B.n459 B.n444 71.676
R2027 B.n455 B.n445 71.676
R2028 B.n446 B.n395 71.676
R2029 B.n662 B.n392 69.5456
R2030 B.n810 B.n809 69.5456
R2031 B.n545 B.n452 59.5399
R2032 B.n566 B.n450 59.5399
R2033 B.n121 B.n120 59.5399
R2034 B.n118 B.n117 59.5399
R2035 B.n452 B.n451 54.6914
R2036 B.n450 B.n449 54.6914
R2037 B.n120 B.n119 54.6914
R2038 B.n117 B.n116 54.6914
R2039 B.n668 B.n392 38.4482
R2040 B.n668 B.n388 38.4482
R2041 B.n674 B.n388 38.4482
R2042 B.n674 B.n384 38.4482
R2043 B.n680 B.n384 38.4482
R2044 B.n680 B.n380 38.4482
R2045 B.n686 B.n380 38.4482
R2046 B.n692 B.n376 38.4482
R2047 B.n692 B.n372 38.4482
R2048 B.n698 B.n372 38.4482
R2049 B.n698 B.n368 38.4482
R2050 B.n704 B.n368 38.4482
R2051 B.n704 B.n364 38.4482
R2052 B.n710 B.n364 38.4482
R2053 B.n710 B.n360 38.4482
R2054 B.n717 B.n360 38.4482
R2055 B.n717 B.n716 38.4482
R2056 B.n723 B.n353 38.4482
R2057 B.n729 B.n353 38.4482
R2058 B.n729 B.n349 38.4482
R2059 B.n735 B.n349 38.4482
R2060 B.n735 B.n345 38.4482
R2061 B.n741 B.n345 38.4482
R2062 B.n741 B.n341 38.4482
R2063 B.n747 B.n341 38.4482
R2064 B.n754 B.n337 38.4482
R2065 B.n754 B.n333 38.4482
R2066 B.n760 B.n333 38.4482
R2067 B.n760 B.n4 38.4482
R2068 B.n875 B.n4 38.4482
R2069 B.n875 B.n874 38.4482
R2070 B.n874 B.n873 38.4482
R2071 B.n873 B.n8 38.4482
R2072 B.n867 B.n8 38.4482
R2073 B.n867 B.n866 38.4482
R2074 B.n865 B.n15 38.4482
R2075 B.n859 B.n15 38.4482
R2076 B.n859 B.n858 38.4482
R2077 B.n858 B.n857 38.4482
R2078 B.n857 B.n22 38.4482
R2079 B.n851 B.n22 38.4482
R2080 B.n851 B.n850 38.4482
R2081 B.n850 B.n849 38.4482
R2082 B.n843 B.n32 38.4482
R2083 B.n843 B.n842 38.4482
R2084 B.n842 B.n841 38.4482
R2085 B.n841 B.n36 38.4482
R2086 B.n835 B.n36 38.4482
R2087 B.n835 B.n834 38.4482
R2088 B.n834 B.n833 38.4482
R2089 B.n833 B.n43 38.4482
R2090 B.n827 B.n43 38.4482
R2091 B.n827 B.n826 38.4482
R2092 B.n825 B.n50 38.4482
R2093 B.n819 B.n50 38.4482
R2094 B.n819 B.n818 38.4482
R2095 B.n818 B.n817 38.4482
R2096 B.n817 B.n57 38.4482
R2097 B.n811 B.n57 38.4482
R2098 B.n811 B.n810 38.4482
R2099 B.n716 B.t3 36.752
R2100 B.n32 B.t1 36.752
R2101 B.n123 B.n59 30.4395
R2102 B.n806 B.n805 30.4395
R2103 B.n665 B.n664 30.4395
R2104 B.n659 B.n390 30.4395
R2105 B.t2 B.n337 28.8363
R2106 B.n866 B.t0 28.8363
R2107 B.t5 B.n376 20.9206
R2108 B.n826 B.t9 20.9206
R2109 B B.n877 18.0485
R2110 B.n686 B.t5 17.5281
R2111 B.t9 B.n825 17.5281
R2112 B.n124 B.n123 10.6151
R2113 B.n127 B.n124 10.6151
R2114 B.n128 B.n127 10.6151
R2115 B.n131 B.n128 10.6151
R2116 B.n132 B.n131 10.6151
R2117 B.n135 B.n132 10.6151
R2118 B.n136 B.n135 10.6151
R2119 B.n139 B.n136 10.6151
R2120 B.n140 B.n139 10.6151
R2121 B.n143 B.n140 10.6151
R2122 B.n144 B.n143 10.6151
R2123 B.n147 B.n144 10.6151
R2124 B.n148 B.n147 10.6151
R2125 B.n151 B.n148 10.6151
R2126 B.n152 B.n151 10.6151
R2127 B.n155 B.n152 10.6151
R2128 B.n156 B.n155 10.6151
R2129 B.n159 B.n156 10.6151
R2130 B.n160 B.n159 10.6151
R2131 B.n163 B.n160 10.6151
R2132 B.n164 B.n163 10.6151
R2133 B.n167 B.n164 10.6151
R2134 B.n168 B.n167 10.6151
R2135 B.n171 B.n168 10.6151
R2136 B.n172 B.n171 10.6151
R2137 B.n175 B.n172 10.6151
R2138 B.n176 B.n175 10.6151
R2139 B.n179 B.n176 10.6151
R2140 B.n180 B.n179 10.6151
R2141 B.n183 B.n180 10.6151
R2142 B.n184 B.n183 10.6151
R2143 B.n187 B.n184 10.6151
R2144 B.n188 B.n187 10.6151
R2145 B.n191 B.n188 10.6151
R2146 B.n192 B.n191 10.6151
R2147 B.n195 B.n192 10.6151
R2148 B.n196 B.n195 10.6151
R2149 B.n199 B.n196 10.6151
R2150 B.n200 B.n199 10.6151
R2151 B.n203 B.n200 10.6151
R2152 B.n204 B.n203 10.6151
R2153 B.n207 B.n204 10.6151
R2154 B.n208 B.n207 10.6151
R2155 B.n211 B.n208 10.6151
R2156 B.n212 B.n211 10.6151
R2157 B.n215 B.n212 10.6151
R2158 B.n216 B.n215 10.6151
R2159 B.n220 B.n219 10.6151
R2160 B.n223 B.n220 10.6151
R2161 B.n224 B.n223 10.6151
R2162 B.n227 B.n224 10.6151
R2163 B.n228 B.n227 10.6151
R2164 B.n231 B.n228 10.6151
R2165 B.n232 B.n231 10.6151
R2166 B.n235 B.n232 10.6151
R2167 B.n236 B.n235 10.6151
R2168 B.n240 B.n239 10.6151
R2169 B.n243 B.n240 10.6151
R2170 B.n244 B.n243 10.6151
R2171 B.n247 B.n244 10.6151
R2172 B.n248 B.n247 10.6151
R2173 B.n251 B.n248 10.6151
R2174 B.n252 B.n251 10.6151
R2175 B.n255 B.n252 10.6151
R2176 B.n256 B.n255 10.6151
R2177 B.n259 B.n256 10.6151
R2178 B.n260 B.n259 10.6151
R2179 B.n263 B.n260 10.6151
R2180 B.n264 B.n263 10.6151
R2181 B.n267 B.n264 10.6151
R2182 B.n268 B.n267 10.6151
R2183 B.n271 B.n268 10.6151
R2184 B.n272 B.n271 10.6151
R2185 B.n275 B.n272 10.6151
R2186 B.n276 B.n275 10.6151
R2187 B.n279 B.n276 10.6151
R2188 B.n280 B.n279 10.6151
R2189 B.n283 B.n280 10.6151
R2190 B.n284 B.n283 10.6151
R2191 B.n287 B.n284 10.6151
R2192 B.n288 B.n287 10.6151
R2193 B.n291 B.n288 10.6151
R2194 B.n292 B.n291 10.6151
R2195 B.n295 B.n292 10.6151
R2196 B.n296 B.n295 10.6151
R2197 B.n299 B.n296 10.6151
R2198 B.n300 B.n299 10.6151
R2199 B.n303 B.n300 10.6151
R2200 B.n304 B.n303 10.6151
R2201 B.n307 B.n304 10.6151
R2202 B.n308 B.n307 10.6151
R2203 B.n311 B.n308 10.6151
R2204 B.n312 B.n311 10.6151
R2205 B.n315 B.n312 10.6151
R2206 B.n316 B.n315 10.6151
R2207 B.n319 B.n316 10.6151
R2208 B.n320 B.n319 10.6151
R2209 B.n323 B.n320 10.6151
R2210 B.n324 B.n323 10.6151
R2211 B.n327 B.n324 10.6151
R2212 B.n329 B.n327 10.6151
R2213 B.n330 B.n329 10.6151
R2214 B.n806 B.n330 10.6151
R2215 B.n666 B.n665 10.6151
R2216 B.n666 B.n386 10.6151
R2217 B.n676 B.n386 10.6151
R2218 B.n677 B.n676 10.6151
R2219 B.n678 B.n677 10.6151
R2220 B.n678 B.n378 10.6151
R2221 B.n688 B.n378 10.6151
R2222 B.n689 B.n688 10.6151
R2223 B.n690 B.n689 10.6151
R2224 B.n690 B.n370 10.6151
R2225 B.n700 B.n370 10.6151
R2226 B.n701 B.n700 10.6151
R2227 B.n702 B.n701 10.6151
R2228 B.n702 B.n362 10.6151
R2229 B.n712 B.n362 10.6151
R2230 B.n713 B.n712 10.6151
R2231 B.n714 B.n713 10.6151
R2232 B.n714 B.n355 10.6151
R2233 B.n725 B.n355 10.6151
R2234 B.n726 B.n725 10.6151
R2235 B.n727 B.n726 10.6151
R2236 B.n727 B.n347 10.6151
R2237 B.n737 B.n347 10.6151
R2238 B.n738 B.n737 10.6151
R2239 B.n739 B.n738 10.6151
R2240 B.n739 B.n339 10.6151
R2241 B.n749 B.n339 10.6151
R2242 B.n750 B.n749 10.6151
R2243 B.n752 B.n750 10.6151
R2244 B.n752 B.n751 10.6151
R2245 B.n751 B.n331 10.6151
R2246 B.n763 B.n331 10.6151
R2247 B.n764 B.n763 10.6151
R2248 B.n765 B.n764 10.6151
R2249 B.n766 B.n765 10.6151
R2250 B.n768 B.n766 10.6151
R2251 B.n769 B.n768 10.6151
R2252 B.n770 B.n769 10.6151
R2253 B.n771 B.n770 10.6151
R2254 B.n773 B.n771 10.6151
R2255 B.n774 B.n773 10.6151
R2256 B.n775 B.n774 10.6151
R2257 B.n776 B.n775 10.6151
R2258 B.n778 B.n776 10.6151
R2259 B.n779 B.n778 10.6151
R2260 B.n780 B.n779 10.6151
R2261 B.n781 B.n780 10.6151
R2262 B.n783 B.n781 10.6151
R2263 B.n784 B.n783 10.6151
R2264 B.n785 B.n784 10.6151
R2265 B.n786 B.n785 10.6151
R2266 B.n788 B.n786 10.6151
R2267 B.n789 B.n788 10.6151
R2268 B.n790 B.n789 10.6151
R2269 B.n791 B.n790 10.6151
R2270 B.n793 B.n791 10.6151
R2271 B.n794 B.n793 10.6151
R2272 B.n795 B.n794 10.6151
R2273 B.n796 B.n795 10.6151
R2274 B.n798 B.n796 10.6151
R2275 B.n799 B.n798 10.6151
R2276 B.n800 B.n799 10.6151
R2277 B.n801 B.n800 10.6151
R2278 B.n803 B.n801 10.6151
R2279 B.n804 B.n803 10.6151
R2280 B.n805 B.n804 10.6151
R2281 B.n659 B.n658 10.6151
R2282 B.n658 B.n657 10.6151
R2283 B.n657 B.n656 10.6151
R2284 B.n656 B.n654 10.6151
R2285 B.n654 B.n651 10.6151
R2286 B.n651 B.n650 10.6151
R2287 B.n650 B.n647 10.6151
R2288 B.n647 B.n646 10.6151
R2289 B.n646 B.n643 10.6151
R2290 B.n643 B.n642 10.6151
R2291 B.n642 B.n639 10.6151
R2292 B.n639 B.n638 10.6151
R2293 B.n638 B.n635 10.6151
R2294 B.n635 B.n634 10.6151
R2295 B.n634 B.n631 10.6151
R2296 B.n631 B.n630 10.6151
R2297 B.n630 B.n627 10.6151
R2298 B.n627 B.n626 10.6151
R2299 B.n626 B.n623 10.6151
R2300 B.n623 B.n622 10.6151
R2301 B.n622 B.n619 10.6151
R2302 B.n619 B.n618 10.6151
R2303 B.n618 B.n615 10.6151
R2304 B.n615 B.n614 10.6151
R2305 B.n614 B.n611 10.6151
R2306 B.n611 B.n610 10.6151
R2307 B.n610 B.n607 10.6151
R2308 B.n607 B.n606 10.6151
R2309 B.n606 B.n603 10.6151
R2310 B.n603 B.n602 10.6151
R2311 B.n602 B.n599 10.6151
R2312 B.n599 B.n598 10.6151
R2313 B.n598 B.n595 10.6151
R2314 B.n595 B.n594 10.6151
R2315 B.n594 B.n591 10.6151
R2316 B.n591 B.n590 10.6151
R2317 B.n590 B.n587 10.6151
R2318 B.n587 B.n586 10.6151
R2319 B.n586 B.n583 10.6151
R2320 B.n583 B.n582 10.6151
R2321 B.n582 B.n579 10.6151
R2322 B.n579 B.n578 10.6151
R2323 B.n578 B.n575 10.6151
R2324 B.n575 B.n574 10.6151
R2325 B.n574 B.n571 10.6151
R2326 B.n571 B.n570 10.6151
R2327 B.n570 B.n567 10.6151
R2328 B.n565 B.n562 10.6151
R2329 B.n562 B.n561 10.6151
R2330 B.n561 B.n558 10.6151
R2331 B.n558 B.n557 10.6151
R2332 B.n557 B.n554 10.6151
R2333 B.n554 B.n553 10.6151
R2334 B.n553 B.n550 10.6151
R2335 B.n550 B.n549 10.6151
R2336 B.n549 B.n546 10.6151
R2337 B.n544 B.n541 10.6151
R2338 B.n541 B.n540 10.6151
R2339 B.n540 B.n537 10.6151
R2340 B.n537 B.n536 10.6151
R2341 B.n536 B.n533 10.6151
R2342 B.n533 B.n532 10.6151
R2343 B.n532 B.n529 10.6151
R2344 B.n529 B.n528 10.6151
R2345 B.n528 B.n525 10.6151
R2346 B.n525 B.n524 10.6151
R2347 B.n524 B.n521 10.6151
R2348 B.n521 B.n520 10.6151
R2349 B.n520 B.n517 10.6151
R2350 B.n517 B.n516 10.6151
R2351 B.n516 B.n513 10.6151
R2352 B.n513 B.n512 10.6151
R2353 B.n512 B.n509 10.6151
R2354 B.n509 B.n508 10.6151
R2355 B.n508 B.n505 10.6151
R2356 B.n505 B.n504 10.6151
R2357 B.n504 B.n501 10.6151
R2358 B.n501 B.n500 10.6151
R2359 B.n500 B.n497 10.6151
R2360 B.n497 B.n496 10.6151
R2361 B.n496 B.n493 10.6151
R2362 B.n493 B.n492 10.6151
R2363 B.n492 B.n489 10.6151
R2364 B.n489 B.n488 10.6151
R2365 B.n488 B.n485 10.6151
R2366 B.n485 B.n484 10.6151
R2367 B.n484 B.n481 10.6151
R2368 B.n481 B.n480 10.6151
R2369 B.n480 B.n477 10.6151
R2370 B.n477 B.n476 10.6151
R2371 B.n476 B.n473 10.6151
R2372 B.n473 B.n472 10.6151
R2373 B.n472 B.n469 10.6151
R2374 B.n469 B.n468 10.6151
R2375 B.n468 B.n465 10.6151
R2376 B.n465 B.n464 10.6151
R2377 B.n464 B.n461 10.6151
R2378 B.n461 B.n460 10.6151
R2379 B.n460 B.n457 10.6151
R2380 B.n457 B.n456 10.6151
R2381 B.n456 B.n453 10.6151
R2382 B.n453 B.n394 10.6151
R2383 B.n664 B.n394 10.6151
R2384 B.n670 B.n390 10.6151
R2385 B.n671 B.n670 10.6151
R2386 B.n672 B.n671 10.6151
R2387 B.n672 B.n382 10.6151
R2388 B.n682 B.n382 10.6151
R2389 B.n683 B.n682 10.6151
R2390 B.n684 B.n683 10.6151
R2391 B.n684 B.n374 10.6151
R2392 B.n694 B.n374 10.6151
R2393 B.n695 B.n694 10.6151
R2394 B.n696 B.n695 10.6151
R2395 B.n696 B.n366 10.6151
R2396 B.n706 B.n366 10.6151
R2397 B.n707 B.n706 10.6151
R2398 B.n708 B.n707 10.6151
R2399 B.n708 B.n358 10.6151
R2400 B.n719 B.n358 10.6151
R2401 B.n720 B.n719 10.6151
R2402 B.n721 B.n720 10.6151
R2403 B.n721 B.n351 10.6151
R2404 B.n731 B.n351 10.6151
R2405 B.n732 B.n731 10.6151
R2406 B.n733 B.n732 10.6151
R2407 B.n733 B.n343 10.6151
R2408 B.n743 B.n343 10.6151
R2409 B.n744 B.n743 10.6151
R2410 B.n745 B.n744 10.6151
R2411 B.n745 B.n335 10.6151
R2412 B.n756 B.n335 10.6151
R2413 B.n757 B.n756 10.6151
R2414 B.n758 B.n757 10.6151
R2415 B.n758 B.n0 10.6151
R2416 B.n871 B.n1 10.6151
R2417 B.n871 B.n870 10.6151
R2418 B.n870 B.n869 10.6151
R2419 B.n869 B.n10 10.6151
R2420 B.n863 B.n10 10.6151
R2421 B.n863 B.n862 10.6151
R2422 B.n862 B.n861 10.6151
R2423 B.n861 B.n17 10.6151
R2424 B.n855 B.n17 10.6151
R2425 B.n855 B.n854 10.6151
R2426 B.n854 B.n853 10.6151
R2427 B.n853 B.n24 10.6151
R2428 B.n847 B.n24 10.6151
R2429 B.n847 B.n846 10.6151
R2430 B.n846 B.n845 10.6151
R2431 B.n845 B.n30 10.6151
R2432 B.n839 B.n30 10.6151
R2433 B.n839 B.n838 10.6151
R2434 B.n838 B.n837 10.6151
R2435 B.n837 B.n38 10.6151
R2436 B.n831 B.n38 10.6151
R2437 B.n831 B.n830 10.6151
R2438 B.n830 B.n829 10.6151
R2439 B.n829 B.n45 10.6151
R2440 B.n823 B.n45 10.6151
R2441 B.n823 B.n822 10.6151
R2442 B.n822 B.n821 10.6151
R2443 B.n821 B.n52 10.6151
R2444 B.n815 B.n52 10.6151
R2445 B.n815 B.n814 10.6151
R2446 B.n814 B.n813 10.6151
R2447 B.n813 B.n59 10.6151
R2448 B.n747 B.t2 9.61243
R2449 B.t0 B.n865 9.61243
R2450 B.n216 B.n121 9.36635
R2451 B.n239 B.n118 9.36635
R2452 B.n567 B.n566 9.36635
R2453 B.n545 B.n544 9.36635
R2454 B.n877 B.n0 2.81026
R2455 B.n877 B.n1 2.81026
R2456 B.n723 B.t3 1.69672
R2457 B.n849 B.t1 1.69672
R2458 B.n219 B.n121 1.24928
R2459 B.n236 B.n118 1.24928
R2460 B.n566 B.n565 1.24928
R2461 B.n546 B.n545 1.24928
R2462 VN.n0 VN.t1 172.669
R2463 VN.n1 VN.t3 172.669
R2464 VN.n0 VN.t0 171.912
R2465 VN.n1 VN.t2 171.912
R2466 VN VN.n1 52.38
R2467 VN VN.n0 4.53529
R2468 VDD2.n2 VDD2.n0 102.721
R2469 VDD2.n2 VDD2.n1 59.4888
R2470 VDD2.n1 VDD2.t1 1.39683
R2471 VDD2.n1 VDD2.t0 1.39683
R2472 VDD2.n0 VDD2.t2 1.39683
R2473 VDD2.n0 VDD2.t3 1.39683
R2474 VDD2 VDD2.n2 0.0586897
C0 VDD1 VDD2 1.00702f
C1 VN VTAIL 5.30998f
C2 VP VTAIL 5.32409f
C3 VP VN 6.51336f
C4 VDD1 VTAIL 5.91907f
C5 VDD2 VTAIL 5.97254f
C6 VDD1 VN 0.149367f
C7 VDD1 VP 5.74659f
C8 VDD2 VN 5.50889f
C9 VDD2 VP 0.387773f
C10 VDD2 B 3.868826f
C11 VDD1 B 8.15992f
C12 VTAIL B 11.320217f
C13 VN B 10.66825f
C14 VP B 8.848373f
C15 VDD2.t2 B 0.299155f
C16 VDD2.t3 B 0.299155f
C17 VDD2.n0 B 3.44945f
C18 VDD2.t1 B 0.299155f
C19 VDD2.t0 B 0.299155f
C20 VDD2.n1 B 2.68768f
C21 VDD2.n2 B 3.95138f
C22 VN.t1 B 2.678f
C23 VN.t0 B 2.67358f
C24 VN.n0 B 1.73076f
C25 VN.t3 B 2.678f
C26 VN.t2 B 2.67358f
C27 VN.n1 B 3.15392f
C28 VTAIL.n0 B 0.022503f
C29 VTAIL.n1 B 0.015858f
C30 VTAIL.n2 B 0.008521f
C31 VTAIL.n3 B 0.020141f
C32 VTAIL.n4 B 0.009022f
C33 VTAIL.n5 B 0.015858f
C34 VTAIL.n6 B 0.008521f
C35 VTAIL.n7 B 0.020141f
C36 VTAIL.n8 B 0.009022f
C37 VTAIL.n9 B 0.015858f
C38 VTAIL.n10 B 0.008521f
C39 VTAIL.n11 B 0.020141f
C40 VTAIL.n12 B 0.009022f
C41 VTAIL.n13 B 0.015858f
C42 VTAIL.n14 B 0.008772f
C43 VTAIL.n15 B 0.020141f
C44 VTAIL.n16 B 0.009022f
C45 VTAIL.n17 B 0.015858f
C46 VTAIL.n18 B 0.008521f
C47 VTAIL.n19 B 0.020141f
C48 VTAIL.n20 B 0.009022f
C49 VTAIL.n21 B 0.015858f
C50 VTAIL.n22 B 0.008521f
C51 VTAIL.n23 B 0.015106f
C52 VTAIL.n24 B 0.014238f
C53 VTAIL.t0 B 0.034203f
C54 VTAIL.n25 B 0.127603f
C55 VTAIL.n26 B 0.953745f
C56 VTAIL.n27 B 0.008521f
C57 VTAIL.n28 B 0.009022f
C58 VTAIL.n29 B 0.020141f
C59 VTAIL.n30 B 0.020141f
C60 VTAIL.n31 B 0.009022f
C61 VTAIL.n32 B 0.008521f
C62 VTAIL.n33 B 0.015858f
C63 VTAIL.n34 B 0.015858f
C64 VTAIL.n35 B 0.008521f
C65 VTAIL.n36 B 0.009022f
C66 VTAIL.n37 B 0.020141f
C67 VTAIL.n38 B 0.020141f
C68 VTAIL.n39 B 0.009022f
C69 VTAIL.n40 B 0.008521f
C70 VTAIL.n41 B 0.015858f
C71 VTAIL.n42 B 0.015858f
C72 VTAIL.n43 B 0.008521f
C73 VTAIL.n44 B 0.008521f
C74 VTAIL.n45 B 0.009022f
C75 VTAIL.n46 B 0.020141f
C76 VTAIL.n47 B 0.020141f
C77 VTAIL.n48 B 0.020141f
C78 VTAIL.n49 B 0.008772f
C79 VTAIL.n50 B 0.008521f
C80 VTAIL.n51 B 0.015858f
C81 VTAIL.n52 B 0.015858f
C82 VTAIL.n53 B 0.008521f
C83 VTAIL.n54 B 0.009022f
C84 VTAIL.n55 B 0.020141f
C85 VTAIL.n56 B 0.020141f
C86 VTAIL.n57 B 0.009022f
C87 VTAIL.n58 B 0.008521f
C88 VTAIL.n59 B 0.015858f
C89 VTAIL.n60 B 0.015858f
C90 VTAIL.n61 B 0.008521f
C91 VTAIL.n62 B 0.009022f
C92 VTAIL.n63 B 0.020141f
C93 VTAIL.n64 B 0.020141f
C94 VTAIL.n65 B 0.009022f
C95 VTAIL.n66 B 0.008521f
C96 VTAIL.n67 B 0.015858f
C97 VTAIL.n68 B 0.015858f
C98 VTAIL.n69 B 0.008521f
C99 VTAIL.n70 B 0.009022f
C100 VTAIL.n71 B 0.020141f
C101 VTAIL.n72 B 0.04398f
C102 VTAIL.n73 B 0.009022f
C103 VTAIL.n74 B 0.008521f
C104 VTAIL.n75 B 0.034488f
C105 VTAIL.n76 B 0.024579f
C106 VTAIL.n77 B 0.101411f
C107 VTAIL.n78 B 0.022503f
C108 VTAIL.n79 B 0.015858f
C109 VTAIL.n80 B 0.008521f
C110 VTAIL.n81 B 0.020141f
C111 VTAIL.n82 B 0.009022f
C112 VTAIL.n83 B 0.015858f
C113 VTAIL.n84 B 0.008521f
C114 VTAIL.n85 B 0.020141f
C115 VTAIL.n86 B 0.009022f
C116 VTAIL.n87 B 0.015858f
C117 VTAIL.n88 B 0.008521f
C118 VTAIL.n89 B 0.020141f
C119 VTAIL.n90 B 0.009022f
C120 VTAIL.n91 B 0.015858f
C121 VTAIL.n92 B 0.008772f
C122 VTAIL.n93 B 0.020141f
C123 VTAIL.n94 B 0.009022f
C124 VTAIL.n95 B 0.015858f
C125 VTAIL.n96 B 0.008521f
C126 VTAIL.n97 B 0.020141f
C127 VTAIL.n98 B 0.009022f
C128 VTAIL.n99 B 0.015858f
C129 VTAIL.n100 B 0.008521f
C130 VTAIL.n101 B 0.015106f
C131 VTAIL.n102 B 0.014238f
C132 VTAIL.t2 B 0.034203f
C133 VTAIL.n103 B 0.127603f
C134 VTAIL.n104 B 0.953745f
C135 VTAIL.n105 B 0.008521f
C136 VTAIL.n106 B 0.009022f
C137 VTAIL.n107 B 0.020141f
C138 VTAIL.n108 B 0.020141f
C139 VTAIL.n109 B 0.009022f
C140 VTAIL.n110 B 0.008521f
C141 VTAIL.n111 B 0.015858f
C142 VTAIL.n112 B 0.015858f
C143 VTAIL.n113 B 0.008521f
C144 VTAIL.n114 B 0.009022f
C145 VTAIL.n115 B 0.020141f
C146 VTAIL.n116 B 0.020141f
C147 VTAIL.n117 B 0.009022f
C148 VTAIL.n118 B 0.008521f
C149 VTAIL.n119 B 0.015858f
C150 VTAIL.n120 B 0.015858f
C151 VTAIL.n121 B 0.008521f
C152 VTAIL.n122 B 0.008521f
C153 VTAIL.n123 B 0.009022f
C154 VTAIL.n124 B 0.020141f
C155 VTAIL.n125 B 0.020141f
C156 VTAIL.n126 B 0.020141f
C157 VTAIL.n127 B 0.008772f
C158 VTAIL.n128 B 0.008521f
C159 VTAIL.n129 B 0.015858f
C160 VTAIL.n130 B 0.015858f
C161 VTAIL.n131 B 0.008521f
C162 VTAIL.n132 B 0.009022f
C163 VTAIL.n133 B 0.020141f
C164 VTAIL.n134 B 0.020141f
C165 VTAIL.n135 B 0.009022f
C166 VTAIL.n136 B 0.008521f
C167 VTAIL.n137 B 0.015858f
C168 VTAIL.n138 B 0.015858f
C169 VTAIL.n139 B 0.008521f
C170 VTAIL.n140 B 0.009022f
C171 VTAIL.n141 B 0.020141f
C172 VTAIL.n142 B 0.020141f
C173 VTAIL.n143 B 0.009022f
C174 VTAIL.n144 B 0.008521f
C175 VTAIL.n145 B 0.015858f
C176 VTAIL.n146 B 0.015858f
C177 VTAIL.n147 B 0.008521f
C178 VTAIL.n148 B 0.009022f
C179 VTAIL.n149 B 0.020141f
C180 VTAIL.n150 B 0.04398f
C181 VTAIL.n151 B 0.009022f
C182 VTAIL.n152 B 0.008521f
C183 VTAIL.n153 B 0.034488f
C184 VTAIL.n154 B 0.024579f
C185 VTAIL.n155 B 0.160547f
C186 VTAIL.n156 B 0.022503f
C187 VTAIL.n157 B 0.015858f
C188 VTAIL.n158 B 0.008521f
C189 VTAIL.n159 B 0.020141f
C190 VTAIL.n160 B 0.009022f
C191 VTAIL.n161 B 0.015858f
C192 VTAIL.n162 B 0.008521f
C193 VTAIL.n163 B 0.020141f
C194 VTAIL.n164 B 0.009022f
C195 VTAIL.n165 B 0.015858f
C196 VTAIL.n166 B 0.008521f
C197 VTAIL.n167 B 0.020141f
C198 VTAIL.n168 B 0.009022f
C199 VTAIL.n169 B 0.015858f
C200 VTAIL.n170 B 0.008772f
C201 VTAIL.n171 B 0.020141f
C202 VTAIL.n172 B 0.009022f
C203 VTAIL.n173 B 0.015858f
C204 VTAIL.n174 B 0.008521f
C205 VTAIL.n175 B 0.020141f
C206 VTAIL.n176 B 0.009022f
C207 VTAIL.n177 B 0.015858f
C208 VTAIL.n178 B 0.008521f
C209 VTAIL.n179 B 0.015106f
C210 VTAIL.n180 B 0.014238f
C211 VTAIL.t5 B 0.034203f
C212 VTAIL.n181 B 0.127603f
C213 VTAIL.n182 B 0.953745f
C214 VTAIL.n183 B 0.008521f
C215 VTAIL.n184 B 0.009022f
C216 VTAIL.n185 B 0.020141f
C217 VTAIL.n186 B 0.020141f
C218 VTAIL.n187 B 0.009022f
C219 VTAIL.n188 B 0.008521f
C220 VTAIL.n189 B 0.015858f
C221 VTAIL.n190 B 0.015858f
C222 VTAIL.n191 B 0.008521f
C223 VTAIL.n192 B 0.009022f
C224 VTAIL.n193 B 0.020141f
C225 VTAIL.n194 B 0.020141f
C226 VTAIL.n195 B 0.009022f
C227 VTAIL.n196 B 0.008521f
C228 VTAIL.n197 B 0.015858f
C229 VTAIL.n198 B 0.015858f
C230 VTAIL.n199 B 0.008521f
C231 VTAIL.n200 B 0.008521f
C232 VTAIL.n201 B 0.009022f
C233 VTAIL.n202 B 0.020141f
C234 VTAIL.n203 B 0.020141f
C235 VTAIL.n204 B 0.020141f
C236 VTAIL.n205 B 0.008772f
C237 VTAIL.n206 B 0.008521f
C238 VTAIL.n207 B 0.015858f
C239 VTAIL.n208 B 0.015858f
C240 VTAIL.n209 B 0.008521f
C241 VTAIL.n210 B 0.009022f
C242 VTAIL.n211 B 0.020141f
C243 VTAIL.n212 B 0.020141f
C244 VTAIL.n213 B 0.009022f
C245 VTAIL.n214 B 0.008521f
C246 VTAIL.n215 B 0.015858f
C247 VTAIL.n216 B 0.015858f
C248 VTAIL.n217 B 0.008521f
C249 VTAIL.n218 B 0.009022f
C250 VTAIL.n219 B 0.020141f
C251 VTAIL.n220 B 0.020141f
C252 VTAIL.n221 B 0.009022f
C253 VTAIL.n222 B 0.008521f
C254 VTAIL.n223 B 0.015858f
C255 VTAIL.n224 B 0.015858f
C256 VTAIL.n225 B 0.008521f
C257 VTAIL.n226 B 0.009022f
C258 VTAIL.n227 B 0.020141f
C259 VTAIL.n228 B 0.04398f
C260 VTAIL.n229 B 0.009022f
C261 VTAIL.n230 B 0.008521f
C262 VTAIL.n231 B 0.034488f
C263 VTAIL.n232 B 0.024579f
C264 VTAIL.n233 B 1.10077f
C265 VTAIL.n234 B 0.022503f
C266 VTAIL.n235 B 0.015858f
C267 VTAIL.n236 B 0.008521f
C268 VTAIL.n237 B 0.020141f
C269 VTAIL.n238 B 0.009022f
C270 VTAIL.n239 B 0.015858f
C271 VTAIL.n240 B 0.008521f
C272 VTAIL.n241 B 0.020141f
C273 VTAIL.n242 B 0.009022f
C274 VTAIL.n243 B 0.015858f
C275 VTAIL.n244 B 0.008521f
C276 VTAIL.n245 B 0.020141f
C277 VTAIL.n246 B 0.009022f
C278 VTAIL.n247 B 0.015858f
C279 VTAIL.n248 B 0.008772f
C280 VTAIL.n249 B 0.020141f
C281 VTAIL.n250 B 0.008521f
C282 VTAIL.n251 B 0.009022f
C283 VTAIL.n252 B 0.015858f
C284 VTAIL.n253 B 0.008521f
C285 VTAIL.n254 B 0.020141f
C286 VTAIL.n255 B 0.009022f
C287 VTAIL.n256 B 0.015858f
C288 VTAIL.n257 B 0.008521f
C289 VTAIL.n258 B 0.015106f
C290 VTAIL.n259 B 0.014238f
C291 VTAIL.t6 B 0.034203f
C292 VTAIL.n260 B 0.127602f
C293 VTAIL.n261 B 0.953744f
C294 VTAIL.n262 B 0.008521f
C295 VTAIL.n263 B 0.009022f
C296 VTAIL.n264 B 0.020141f
C297 VTAIL.n265 B 0.020141f
C298 VTAIL.n266 B 0.009022f
C299 VTAIL.n267 B 0.008521f
C300 VTAIL.n268 B 0.015858f
C301 VTAIL.n269 B 0.015858f
C302 VTAIL.n270 B 0.008521f
C303 VTAIL.n271 B 0.009022f
C304 VTAIL.n272 B 0.020141f
C305 VTAIL.n273 B 0.020141f
C306 VTAIL.n274 B 0.009022f
C307 VTAIL.n275 B 0.008521f
C308 VTAIL.n276 B 0.015858f
C309 VTAIL.n277 B 0.015858f
C310 VTAIL.n278 B 0.008521f
C311 VTAIL.n279 B 0.009022f
C312 VTAIL.n280 B 0.020141f
C313 VTAIL.n281 B 0.020141f
C314 VTAIL.n282 B 0.020141f
C315 VTAIL.n283 B 0.008772f
C316 VTAIL.n284 B 0.008521f
C317 VTAIL.n285 B 0.015858f
C318 VTAIL.n286 B 0.015858f
C319 VTAIL.n287 B 0.008521f
C320 VTAIL.n288 B 0.009022f
C321 VTAIL.n289 B 0.020141f
C322 VTAIL.n290 B 0.020141f
C323 VTAIL.n291 B 0.009022f
C324 VTAIL.n292 B 0.008521f
C325 VTAIL.n293 B 0.015858f
C326 VTAIL.n294 B 0.015858f
C327 VTAIL.n295 B 0.008521f
C328 VTAIL.n296 B 0.009022f
C329 VTAIL.n297 B 0.020141f
C330 VTAIL.n298 B 0.020141f
C331 VTAIL.n299 B 0.009022f
C332 VTAIL.n300 B 0.008521f
C333 VTAIL.n301 B 0.015858f
C334 VTAIL.n302 B 0.015858f
C335 VTAIL.n303 B 0.008521f
C336 VTAIL.n304 B 0.009022f
C337 VTAIL.n305 B 0.020141f
C338 VTAIL.n306 B 0.04398f
C339 VTAIL.n307 B 0.009022f
C340 VTAIL.n308 B 0.008521f
C341 VTAIL.n309 B 0.034488f
C342 VTAIL.n310 B 0.024579f
C343 VTAIL.n311 B 1.10077f
C344 VTAIL.n312 B 0.022503f
C345 VTAIL.n313 B 0.015858f
C346 VTAIL.n314 B 0.008521f
C347 VTAIL.n315 B 0.020141f
C348 VTAIL.n316 B 0.009022f
C349 VTAIL.n317 B 0.015858f
C350 VTAIL.n318 B 0.008521f
C351 VTAIL.n319 B 0.020141f
C352 VTAIL.n320 B 0.009022f
C353 VTAIL.n321 B 0.015858f
C354 VTAIL.n322 B 0.008521f
C355 VTAIL.n323 B 0.020141f
C356 VTAIL.n324 B 0.009022f
C357 VTAIL.n325 B 0.015858f
C358 VTAIL.n326 B 0.008772f
C359 VTAIL.n327 B 0.020141f
C360 VTAIL.n328 B 0.008521f
C361 VTAIL.n329 B 0.009022f
C362 VTAIL.n330 B 0.015858f
C363 VTAIL.n331 B 0.008521f
C364 VTAIL.n332 B 0.020141f
C365 VTAIL.n333 B 0.009022f
C366 VTAIL.n334 B 0.015858f
C367 VTAIL.n335 B 0.008521f
C368 VTAIL.n336 B 0.015106f
C369 VTAIL.n337 B 0.014238f
C370 VTAIL.t7 B 0.034203f
C371 VTAIL.n338 B 0.127602f
C372 VTAIL.n339 B 0.953744f
C373 VTAIL.n340 B 0.008521f
C374 VTAIL.n341 B 0.009022f
C375 VTAIL.n342 B 0.020141f
C376 VTAIL.n343 B 0.020141f
C377 VTAIL.n344 B 0.009022f
C378 VTAIL.n345 B 0.008521f
C379 VTAIL.n346 B 0.015858f
C380 VTAIL.n347 B 0.015858f
C381 VTAIL.n348 B 0.008521f
C382 VTAIL.n349 B 0.009022f
C383 VTAIL.n350 B 0.020141f
C384 VTAIL.n351 B 0.020141f
C385 VTAIL.n352 B 0.009022f
C386 VTAIL.n353 B 0.008521f
C387 VTAIL.n354 B 0.015858f
C388 VTAIL.n355 B 0.015858f
C389 VTAIL.n356 B 0.008521f
C390 VTAIL.n357 B 0.009022f
C391 VTAIL.n358 B 0.020141f
C392 VTAIL.n359 B 0.020141f
C393 VTAIL.n360 B 0.020141f
C394 VTAIL.n361 B 0.008772f
C395 VTAIL.n362 B 0.008521f
C396 VTAIL.n363 B 0.015858f
C397 VTAIL.n364 B 0.015858f
C398 VTAIL.n365 B 0.008521f
C399 VTAIL.n366 B 0.009022f
C400 VTAIL.n367 B 0.020141f
C401 VTAIL.n368 B 0.020141f
C402 VTAIL.n369 B 0.009022f
C403 VTAIL.n370 B 0.008521f
C404 VTAIL.n371 B 0.015858f
C405 VTAIL.n372 B 0.015858f
C406 VTAIL.n373 B 0.008521f
C407 VTAIL.n374 B 0.009022f
C408 VTAIL.n375 B 0.020141f
C409 VTAIL.n376 B 0.020141f
C410 VTAIL.n377 B 0.009022f
C411 VTAIL.n378 B 0.008521f
C412 VTAIL.n379 B 0.015858f
C413 VTAIL.n380 B 0.015858f
C414 VTAIL.n381 B 0.008521f
C415 VTAIL.n382 B 0.009022f
C416 VTAIL.n383 B 0.020141f
C417 VTAIL.n384 B 0.04398f
C418 VTAIL.n385 B 0.009022f
C419 VTAIL.n386 B 0.008521f
C420 VTAIL.n387 B 0.034488f
C421 VTAIL.n388 B 0.024579f
C422 VTAIL.n389 B 0.160547f
C423 VTAIL.n390 B 0.022503f
C424 VTAIL.n391 B 0.015858f
C425 VTAIL.n392 B 0.008521f
C426 VTAIL.n393 B 0.020141f
C427 VTAIL.n394 B 0.009022f
C428 VTAIL.n395 B 0.015858f
C429 VTAIL.n396 B 0.008521f
C430 VTAIL.n397 B 0.020141f
C431 VTAIL.n398 B 0.009022f
C432 VTAIL.n399 B 0.015858f
C433 VTAIL.n400 B 0.008521f
C434 VTAIL.n401 B 0.020141f
C435 VTAIL.n402 B 0.009022f
C436 VTAIL.n403 B 0.015858f
C437 VTAIL.n404 B 0.008772f
C438 VTAIL.n405 B 0.020141f
C439 VTAIL.n406 B 0.008521f
C440 VTAIL.n407 B 0.009022f
C441 VTAIL.n408 B 0.015858f
C442 VTAIL.n409 B 0.008521f
C443 VTAIL.n410 B 0.020141f
C444 VTAIL.n411 B 0.009022f
C445 VTAIL.n412 B 0.015858f
C446 VTAIL.n413 B 0.008521f
C447 VTAIL.n414 B 0.015106f
C448 VTAIL.n415 B 0.014238f
C449 VTAIL.t3 B 0.034203f
C450 VTAIL.n416 B 0.127602f
C451 VTAIL.n417 B 0.953744f
C452 VTAIL.n418 B 0.008521f
C453 VTAIL.n419 B 0.009022f
C454 VTAIL.n420 B 0.020141f
C455 VTAIL.n421 B 0.020141f
C456 VTAIL.n422 B 0.009022f
C457 VTAIL.n423 B 0.008521f
C458 VTAIL.n424 B 0.015858f
C459 VTAIL.n425 B 0.015858f
C460 VTAIL.n426 B 0.008521f
C461 VTAIL.n427 B 0.009022f
C462 VTAIL.n428 B 0.020141f
C463 VTAIL.n429 B 0.020141f
C464 VTAIL.n430 B 0.009022f
C465 VTAIL.n431 B 0.008521f
C466 VTAIL.n432 B 0.015858f
C467 VTAIL.n433 B 0.015858f
C468 VTAIL.n434 B 0.008521f
C469 VTAIL.n435 B 0.009022f
C470 VTAIL.n436 B 0.020141f
C471 VTAIL.n437 B 0.020141f
C472 VTAIL.n438 B 0.020141f
C473 VTAIL.n439 B 0.008772f
C474 VTAIL.n440 B 0.008521f
C475 VTAIL.n441 B 0.015858f
C476 VTAIL.n442 B 0.015858f
C477 VTAIL.n443 B 0.008521f
C478 VTAIL.n444 B 0.009022f
C479 VTAIL.n445 B 0.020141f
C480 VTAIL.n446 B 0.020141f
C481 VTAIL.n447 B 0.009022f
C482 VTAIL.n448 B 0.008521f
C483 VTAIL.n449 B 0.015858f
C484 VTAIL.n450 B 0.015858f
C485 VTAIL.n451 B 0.008521f
C486 VTAIL.n452 B 0.009022f
C487 VTAIL.n453 B 0.020141f
C488 VTAIL.n454 B 0.020141f
C489 VTAIL.n455 B 0.009022f
C490 VTAIL.n456 B 0.008521f
C491 VTAIL.n457 B 0.015858f
C492 VTAIL.n458 B 0.015858f
C493 VTAIL.n459 B 0.008521f
C494 VTAIL.n460 B 0.009022f
C495 VTAIL.n461 B 0.020141f
C496 VTAIL.n462 B 0.04398f
C497 VTAIL.n463 B 0.009022f
C498 VTAIL.n464 B 0.008521f
C499 VTAIL.n465 B 0.034488f
C500 VTAIL.n466 B 0.024579f
C501 VTAIL.n467 B 0.160547f
C502 VTAIL.n468 B 0.022503f
C503 VTAIL.n469 B 0.015858f
C504 VTAIL.n470 B 0.008521f
C505 VTAIL.n471 B 0.020141f
C506 VTAIL.n472 B 0.009022f
C507 VTAIL.n473 B 0.015858f
C508 VTAIL.n474 B 0.008521f
C509 VTAIL.n475 B 0.020141f
C510 VTAIL.n476 B 0.009022f
C511 VTAIL.n477 B 0.015858f
C512 VTAIL.n478 B 0.008521f
C513 VTAIL.n479 B 0.020141f
C514 VTAIL.n480 B 0.009022f
C515 VTAIL.n481 B 0.015858f
C516 VTAIL.n482 B 0.008772f
C517 VTAIL.n483 B 0.020141f
C518 VTAIL.n484 B 0.008521f
C519 VTAIL.n485 B 0.009022f
C520 VTAIL.n486 B 0.015858f
C521 VTAIL.n487 B 0.008521f
C522 VTAIL.n488 B 0.020141f
C523 VTAIL.n489 B 0.009022f
C524 VTAIL.n490 B 0.015858f
C525 VTAIL.n491 B 0.008521f
C526 VTAIL.n492 B 0.015106f
C527 VTAIL.n493 B 0.014238f
C528 VTAIL.t4 B 0.034203f
C529 VTAIL.n494 B 0.127603f
C530 VTAIL.n495 B 0.953745f
C531 VTAIL.n496 B 0.008521f
C532 VTAIL.n497 B 0.009022f
C533 VTAIL.n498 B 0.020141f
C534 VTAIL.n499 B 0.020141f
C535 VTAIL.n500 B 0.009022f
C536 VTAIL.n501 B 0.008521f
C537 VTAIL.n502 B 0.015858f
C538 VTAIL.n503 B 0.015858f
C539 VTAIL.n504 B 0.008521f
C540 VTAIL.n505 B 0.009022f
C541 VTAIL.n506 B 0.020141f
C542 VTAIL.n507 B 0.020141f
C543 VTAIL.n508 B 0.009022f
C544 VTAIL.n509 B 0.008521f
C545 VTAIL.n510 B 0.015858f
C546 VTAIL.n511 B 0.015858f
C547 VTAIL.n512 B 0.008521f
C548 VTAIL.n513 B 0.009022f
C549 VTAIL.n514 B 0.020141f
C550 VTAIL.n515 B 0.020141f
C551 VTAIL.n516 B 0.020141f
C552 VTAIL.n517 B 0.008772f
C553 VTAIL.n518 B 0.008521f
C554 VTAIL.n519 B 0.015858f
C555 VTAIL.n520 B 0.015858f
C556 VTAIL.n521 B 0.008521f
C557 VTAIL.n522 B 0.009022f
C558 VTAIL.n523 B 0.020141f
C559 VTAIL.n524 B 0.020141f
C560 VTAIL.n525 B 0.009022f
C561 VTAIL.n526 B 0.008521f
C562 VTAIL.n527 B 0.015858f
C563 VTAIL.n528 B 0.015858f
C564 VTAIL.n529 B 0.008521f
C565 VTAIL.n530 B 0.009022f
C566 VTAIL.n531 B 0.020141f
C567 VTAIL.n532 B 0.020141f
C568 VTAIL.n533 B 0.009022f
C569 VTAIL.n534 B 0.008521f
C570 VTAIL.n535 B 0.015858f
C571 VTAIL.n536 B 0.015858f
C572 VTAIL.n537 B 0.008521f
C573 VTAIL.n538 B 0.009022f
C574 VTAIL.n539 B 0.020141f
C575 VTAIL.n540 B 0.04398f
C576 VTAIL.n541 B 0.009022f
C577 VTAIL.n542 B 0.008521f
C578 VTAIL.n543 B 0.034488f
C579 VTAIL.n544 B 0.024579f
C580 VTAIL.n545 B 1.10077f
C581 VTAIL.n546 B 0.022503f
C582 VTAIL.n547 B 0.015858f
C583 VTAIL.n548 B 0.008521f
C584 VTAIL.n549 B 0.020141f
C585 VTAIL.n550 B 0.009022f
C586 VTAIL.n551 B 0.015858f
C587 VTAIL.n552 B 0.008521f
C588 VTAIL.n553 B 0.020141f
C589 VTAIL.n554 B 0.009022f
C590 VTAIL.n555 B 0.015858f
C591 VTAIL.n556 B 0.008521f
C592 VTAIL.n557 B 0.020141f
C593 VTAIL.n558 B 0.009022f
C594 VTAIL.n559 B 0.015858f
C595 VTAIL.n560 B 0.008772f
C596 VTAIL.n561 B 0.020141f
C597 VTAIL.n562 B 0.009022f
C598 VTAIL.n563 B 0.015858f
C599 VTAIL.n564 B 0.008521f
C600 VTAIL.n565 B 0.020141f
C601 VTAIL.n566 B 0.009022f
C602 VTAIL.n567 B 0.015858f
C603 VTAIL.n568 B 0.008521f
C604 VTAIL.n569 B 0.015106f
C605 VTAIL.n570 B 0.014238f
C606 VTAIL.t1 B 0.034203f
C607 VTAIL.n571 B 0.127603f
C608 VTAIL.n572 B 0.953745f
C609 VTAIL.n573 B 0.008521f
C610 VTAIL.n574 B 0.009022f
C611 VTAIL.n575 B 0.020141f
C612 VTAIL.n576 B 0.020141f
C613 VTAIL.n577 B 0.009022f
C614 VTAIL.n578 B 0.008521f
C615 VTAIL.n579 B 0.015858f
C616 VTAIL.n580 B 0.015858f
C617 VTAIL.n581 B 0.008521f
C618 VTAIL.n582 B 0.009022f
C619 VTAIL.n583 B 0.020141f
C620 VTAIL.n584 B 0.020141f
C621 VTAIL.n585 B 0.009022f
C622 VTAIL.n586 B 0.008521f
C623 VTAIL.n587 B 0.015858f
C624 VTAIL.n588 B 0.015858f
C625 VTAIL.n589 B 0.008521f
C626 VTAIL.n590 B 0.008521f
C627 VTAIL.n591 B 0.009022f
C628 VTAIL.n592 B 0.020141f
C629 VTAIL.n593 B 0.020141f
C630 VTAIL.n594 B 0.020141f
C631 VTAIL.n595 B 0.008772f
C632 VTAIL.n596 B 0.008521f
C633 VTAIL.n597 B 0.015858f
C634 VTAIL.n598 B 0.015858f
C635 VTAIL.n599 B 0.008521f
C636 VTAIL.n600 B 0.009022f
C637 VTAIL.n601 B 0.020141f
C638 VTAIL.n602 B 0.020141f
C639 VTAIL.n603 B 0.009022f
C640 VTAIL.n604 B 0.008521f
C641 VTAIL.n605 B 0.015858f
C642 VTAIL.n606 B 0.015858f
C643 VTAIL.n607 B 0.008521f
C644 VTAIL.n608 B 0.009022f
C645 VTAIL.n609 B 0.020141f
C646 VTAIL.n610 B 0.020141f
C647 VTAIL.n611 B 0.009022f
C648 VTAIL.n612 B 0.008521f
C649 VTAIL.n613 B 0.015858f
C650 VTAIL.n614 B 0.015858f
C651 VTAIL.n615 B 0.008521f
C652 VTAIL.n616 B 0.009022f
C653 VTAIL.n617 B 0.020141f
C654 VTAIL.n618 B 0.04398f
C655 VTAIL.n619 B 0.009022f
C656 VTAIL.n620 B 0.008521f
C657 VTAIL.n621 B 0.034488f
C658 VTAIL.n622 B 0.024579f
C659 VTAIL.n623 B 1.03569f
C660 VDD1.t0 B 0.299191f
C661 VDD1.t1 B 0.299191f
C662 VDD1.n0 B 2.68844f
C663 VDD1.t2 B 0.299191f
C664 VDD1.t3 B 0.299191f
C665 VDD1.n1 B 3.47763f
C666 VP.n0 B 0.034132f
C667 VP.t3 B 2.50161f
C668 VP.n1 B 0.037635f
C669 VP.n2 B 0.02589f
C670 VP.t0 B 2.50161f
C671 VP.n3 B 0.957092f
C672 VP.t1 B 2.71011f
C673 VP.t2 B 2.71459f
C674 VP.n4 B 3.18346f
C675 VP.n5 B 1.49535f
C676 VP.n6 B 0.034132f
C677 VP.n7 B 0.031894f
C678 VP.n8 B 0.048011f
C679 VP.n9 B 0.037635f
C680 VP.n10 B 0.02589f
C681 VP.n11 B 0.02589f
C682 VP.n12 B 0.02589f
C683 VP.n13 B 0.048011f
C684 VP.n14 B 0.031894f
C685 VP.n15 B 0.957092f
C686 VP.n16 B 0.042519f
.ends

