* NGSPICE file created from diff_pair_sample_1020.ext - technology: sky130A

.subckt diff_pair_sample_1020 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t2 w_n2286_n1704# sky130_fd_pr__pfet_01v8 ad=1.4352 pd=8.14 as=1.4352 ps=8.14 w=3.68 l=2.96
X1 VDD1.t0 VP.t1 VTAIL.t1 w_n2286_n1704# sky130_fd_pr__pfet_01v8 ad=1.4352 pd=8.14 as=1.4352 ps=8.14 w=3.68 l=2.96
X2 B.t11 B.t9 B.t10 w_n2286_n1704# sky130_fd_pr__pfet_01v8 ad=1.4352 pd=8.14 as=0 ps=0 w=3.68 l=2.96
X3 VDD2.t1 VN.t0 VTAIL.t3 w_n2286_n1704# sky130_fd_pr__pfet_01v8 ad=1.4352 pd=8.14 as=1.4352 ps=8.14 w=3.68 l=2.96
X4 VDD2.t0 VN.t1 VTAIL.t0 w_n2286_n1704# sky130_fd_pr__pfet_01v8 ad=1.4352 pd=8.14 as=1.4352 ps=8.14 w=3.68 l=2.96
X5 B.t8 B.t6 B.t7 w_n2286_n1704# sky130_fd_pr__pfet_01v8 ad=1.4352 pd=8.14 as=0 ps=0 w=3.68 l=2.96
X6 B.t5 B.t3 B.t4 w_n2286_n1704# sky130_fd_pr__pfet_01v8 ad=1.4352 pd=8.14 as=0 ps=0 w=3.68 l=2.96
X7 B.t2 B.t0 B.t1 w_n2286_n1704# sky130_fd_pr__pfet_01v8 ad=1.4352 pd=8.14 as=0 ps=0 w=3.68 l=2.96
R0 VP.n0 VP.t1 110.409
R1 VP.n0 VP.t0 71.1004
R2 VP VP.n0 0.431812
R3 VTAIL.n1 VTAIL.t3 115.942
R4 VTAIL.n3 VTAIL.t0 115.942
R5 VTAIL.n0 VTAIL.t2 115.942
R6 VTAIL.n2 VTAIL.t1 115.942
R7 VTAIL.n1 VTAIL.n0 21.2117
R8 VTAIL.n3 VTAIL.n2 18.3755
R9 VTAIL.n2 VTAIL.n1 1.88843
R10 VTAIL VTAIL.n0 1.23757
R11 VTAIL VTAIL.n3 0.651362
R12 VDD1 VDD1.t1 166.357
R13 VDD1 VDD1.t0 133.387
R14 B.n215 B.n70 585
R15 B.n214 B.n213 585
R16 B.n212 B.n71 585
R17 B.n211 B.n210 585
R18 B.n209 B.n72 585
R19 B.n208 B.n207 585
R20 B.n206 B.n73 585
R21 B.n205 B.n204 585
R22 B.n203 B.n74 585
R23 B.n202 B.n201 585
R24 B.n200 B.n75 585
R25 B.n199 B.n198 585
R26 B.n197 B.n76 585
R27 B.n196 B.n195 585
R28 B.n194 B.n77 585
R29 B.n193 B.n192 585
R30 B.n191 B.n78 585
R31 B.n190 B.n189 585
R32 B.n185 B.n79 585
R33 B.n184 B.n183 585
R34 B.n182 B.n80 585
R35 B.n181 B.n180 585
R36 B.n179 B.n81 585
R37 B.n178 B.n177 585
R38 B.n176 B.n82 585
R39 B.n175 B.n174 585
R40 B.n173 B.n83 585
R41 B.n171 B.n170 585
R42 B.n169 B.n86 585
R43 B.n168 B.n167 585
R44 B.n166 B.n87 585
R45 B.n165 B.n164 585
R46 B.n163 B.n88 585
R47 B.n162 B.n161 585
R48 B.n160 B.n89 585
R49 B.n159 B.n158 585
R50 B.n157 B.n90 585
R51 B.n156 B.n155 585
R52 B.n154 B.n91 585
R53 B.n153 B.n152 585
R54 B.n151 B.n92 585
R55 B.n150 B.n149 585
R56 B.n148 B.n93 585
R57 B.n147 B.n146 585
R58 B.n217 B.n216 585
R59 B.n218 B.n69 585
R60 B.n220 B.n219 585
R61 B.n221 B.n68 585
R62 B.n223 B.n222 585
R63 B.n224 B.n67 585
R64 B.n226 B.n225 585
R65 B.n227 B.n66 585
R66 B.n229 B.n228 585
R67 B.n230 B.n65 585
R68 B.n232 B.n231 585
R69 B.n233 B.n64 585
R70 B.n235 B.n234 585
R71 B.n236 B.n63 585
R72 B.n238 B.n237 585
R73 B.n239 B.n62 585
R74 B.n241 B.n240 585
R75 B.n242 B.n61 585
R76 B.n244 B.n243 585
R77 B.n245 B.n60 585
R78 B.n247 B.n246 585
R79 B.n248 B.n59 585
R80 B.n250 B.n249 585
R81 B.n251 B.n58 585
R82 B.n253 B.n252 585
R83 B.n254 B.n57 585
R84 B.n256 B.n255 585
R85 B.n257 B.n56 585
R86 B.n259 B.n258 585
R87 B.n260 B.n55 585
R88 B.n262 B.n261 585
R89 B.n263 B.n54 585
R90 B.n265 B.n264 585
R91 B.n266 B.n53 585
R92 B.n268 B.n267 585
R93 B.n269 B.n52 585
R94 B.n271 B.n270 585
R95 B.n272 B.n51 585
R96 B.n274 B.n273 585
R97 B.n275 B.n50 585
R98 B.n277 B.n276 585
R99 B.n278 B.n49 585
R100 B.n280 B.n279 585
R101 B.n281 B.n48 585
R102 B.n283 B.n282 585
R103 B.n284 B.n47 585
R104 B.n286 B.n285 585
R105 B.n287 B.n46 585
R106 B.n289 B.n288 585
R107 B.n290 B.n45 585
R108 B.n292 B.n291 585
R109 B.n293 B.n44 585
R110 B.n295 B.n294 585
R111 B.n296 B.n43 585
R112 B.n298 B.n297 585
R113 B.n299 B.n42 585
R114 B.n367 B.n366 585
R115 B.n365 B.n16 585
R116 B.n364 B.n363 585
R117 B.n362 B.n17 585
R118 B.n361 B.n360 585
R119 B.n359 B.n18 585
R120 B.n358 B.n357 585
R121 B.n356 B.n19 585
R122 B.n355 B.n354 585
R123 B.n353 B.n20 585
R124 B.n352 B.n351 585
R125 B.n350 B.n21 585
R126 B.n349 B.n348 585
R127 B.n347 B.n22 585
R128 B.n346 B.n345 585
R129 B.n344 B.n23 585
R130 B.n343 B.n342 585
R131 B.n341 B.n340 585
R132 B.n339 B.n27 585
R133 B.n338 B.n337 585
R134 B.n336 B.n28 585
R135 B.n335 B.n334 585
R136 B.n333 B.n29 585
R137 B.n332 B.n331 585
R138 B.n330 B.n30 585
R139 B.n329 B.n328 585
R140 B.n327 B.n31 585
R141 B.n325 B.n324 585
R142 B.n323 B.n34 585
R143 B.n322 B.n321 585
R144 B.n320 B.n35 585
R145 B.n319 B.n318 585
R146 B.n317 B.n36 585
R147 B.n316 B.n315 585
R148 B.n314 B.n37 585
R149 B.n313 B.n312 585
R150 B.n311 B.n38 585
R151 B.n310 B.n309 585
R152 B.n308 B.n39 585
R153 B.n307 B.n306 585
R154 B.n305 B.n40 585
R155 B.n304 B.n303 585
R156 B.n302 B.n41 585
R157 B.n301 B.n300 585
R158 B.n368 B.n15 585
R159 B.n370 B.n369 585
R160 B.n371 B.n14 585
R161 B.n373 B.n372 585
R162 B.n374 B.n13 585
R163 B.n376 B.n375 585
R164 B.n377 B.n12 585
R165 B.n379 B.n378 585
R166 B.n380 B.n11 585
R167 B.n382 B.n381 585
R168 B.n383 B.n10 585
R169 B.n385 B.n384 585
R170 B.n386 B.n9 585
R171 B.n388 B.n387 585
R172 B.n389 B.n8 585
R173 B.n391 B.n390 585
R174 B.n392 B.n7 585
R175 B.n394 B.n393 585
R176 B.n395 B.n6 585
R177 B.n397 B.n396 585
R178 B.n398 B.n5 585
R179 B.n400 B.n399 585
R180 B.n401 B.n4 585
R181 B.n403 B.n402 585
R182 B.n404 B.n3 585
R183 B.n406 B.n405 585
R184 B.n407 B.n0 585
R185 B.n2 B.n1 585
R186 B.n108 B.n107 585
R187 B.n109 B.n106 585
R188 B.n111 B.n110 585
R189 B.n112 B.n105 585
R190 B.n114 B.n113 585
R191 B.n115 B.n104 585
R192 B.n117 B.n116 585
R193 B.n118 B.n103 585
R194 B.n120 B.n119 585
R195 B.n121 B.n102 585
R196 B.n123 B.n122 585
R197 B.n124 B.n101 585
R198 B.n126 B.n125 585
R199 B.n127 B.n100 585
R200 B.n129 B.n128 585
R201 B.n130 B.n99 585
R202 B.n132 B.n131 585
R203 B.n133 B.n98 585
R204 B.n135 B.n134 585
R205 B.n136 B.n97 585
R206 B.n138 B.n137 585
R207 B.n139 B.n96 585
R208 B.n141 B.n140 585
R209 B.n142 B.n95 585
R210 B.n144 B.n143 585
R211 B.n145 B.n94 585
R212 B.n146 B.n145 482.89
R213 B.n216 B.n215 482.89
R214 B.n300 B.n299 482.89
R215 B.n366 B.n15 482.89
R216 B.n409 B.n408 256.663
R217 B.n84 B.t9 238.494
R218 B.n186 B.t6 238.494
R219 B.n32 B.t0 238.494
R220 B.n24 B.t3 238.494
R221 B.n408 B.n407 235.042
R222 B.n408 B.n2 235.042
R223 B.n186 B.t7 195.137
R224 B.n32 B.t2 195.137
R225 B.n84 B.t10 195.136
R226 B.n24 B.t5 195.136
R227 B.n146 B.n93 163.367
R228 B.n150 B.n93 163.367
R229 B.n151 B.n150 163.367
R230 B.n152 B.n151 163.367
R231 B.n152 B.n91 163.367
R232 B.n156 B.n91 163.367
R233 B.n157 B.n156 163.367
R234 B.n158 B.n157 163.367
R235 B.n158 B.n89 163.367
R236 B.n162 B.n89 163.367
R237 B.n163 B.n162 163.367
R238 B.n164 B.n163 163.367
R239 B.n164 B.n87 163.367
R240 B.n168 B.n87 163.367
R241 B.n169 B.n168 163.367
R242 B.n170 B.n169 163.367
R243 B.n170 B.n83 163.367
R244 B.n175 B.n83 163.367
R245 B.n176 B.n175 163.367
R246 B.n177 B.n176 163.367
R247 B.n177 B.n81 163.367
R248 B.n181 B.n81 163.367
R249 B.n182 B.n181 163.367
R250 B.n183 B.n182 163.367
R251 B.n183 B.n79 163.367
R252 B.n190 B.n79 163.367
R253 B.n191 B.n190 163.367
R254 B.n192 B.n191 163.367
R255 B.n192 B.n77 163.367
R256 B.n196 B.n77 163.367
R257 B.n197 B.n196 163.367
R258 B.n198 B.n197 163.367
R259 B.n198 B.n75 163.367
R260 B.n202 B.n75 163.367
R261 B.n203 B.n202 163.367
R262 B.n204 B.n203 163.367
R263 B.n204 B.n73 163.367
R264 B.n208 B.n73 163.367
R265 B.n209 B.n208 163.367
R266 B.n210 B.n209 163.367
R267 B.n210 B.n71 163.367
R268 B.n214 B.n71 163.367
R269 B.n215 B.n214 163.367
R270 B.n299 B.n298 163.367
R271 B.n298 B.n43 163.367
R272 B.n294 B.n43 163.367
R273 B.n294 B.n293 163.367
R274 B.n293 B.n292 163.367
R275 B.n292 B.n45 163.367
R276 B.n288 B.n45 163.367
R277 B.n288 B.n287 163.367
R278 B.n287 B.n286 163.367
R279 B.n286 B.n47 163.367
R280 B.n282 B.n47 163.367
R281 B.n282 B.n281 163.367
R282 B.n281 B.n280 163.367
R283 B.n280 B.n49 163.367
R284 B.n276 B.n49 163.367
R285 B.n276 B.n275 163.367
R286 B.n275 B.n274 163.367
R287 B.n274 B.n51 163.367
R288 B.n270 B.n51 163.367
R289 B.n270 B.n269 163.367
R290 B.n269 B.n268 163.367
R291 B.n268 B.n53 163.367
R292 B.n264 B.n53 163.367
R293 B.n264 B.n263 163.367
R294 B.n263 B.n262 163.367
R295 B.n262 B.n55 163.367
R296 B.n258 B.n55 163.367
R297 B.n258 B.n257 163.367
R298 B.n257 B.n256 163.367
R299 B.n256 B.n57 163.367
R300 B.n252 B.n57 163.367
R301 B.n252 B.n251 163.367
R302 B.n251 B.n250 163.367
R303 B.n250 B.n59 163.367
R304 B.n246 B.n59 163.367
R305 B.n246 B.n245 163.367
R306 B.n245 B.n244 163.367
R307 B.n244 B.n61 163.367
R308 B.n240 B.n61 163.367
R309 B.n240 B.n239 163.367
R310 B.n239 B.n238 163.367
R311 B.n238 B.n63 163.367
R312 B.n234 B.n63 163.367
R313 B.n234 B.n233 163.367
R314 B.n233 B.n232 163.367
R315 B.n232 B.n65 163.367
R316 B.n228 B.n65 163.367
R317 B.n228 B.n227 163.367
R318 B.n227 B.n226 163.367
R319 B.n226 B.n67 163.367
R320 B.n222 B.n67 163.367
R321 B.n222 B.n221 163.367
R322 B.n221 B.n220 163.367
R323 B.n220 B.n69 163.367
R324 B.n216 B.n69 163.367
R325 B.n366 B.n365 163.367
R326 B.n365 B.n364 163.367
R327 B.n364 B.n17 163.367
R328 B.n360 B.n17 163.367
R329 B.n360 B.n359 163.367
R330 B.n359 B.n358 163.367
R331 B.n358 B.n19 163.367
R332 B.n354 B.n19 163.367
R333 B.n354 B.n353 163.367
R334 B.n353 B.n352 163.367
R335 B.n352 B.n21 163.367
R336 B.n348 B.n21 163.367
R337 B.n348 B.n347 163.367
R338 B.n347 B.n346 163.367
R339 B.n346 B.n23 163.367
R340 B.n342 B.n23 163.367
R341 B.n342 B.n341 163.367
R342 B.n341 B.n27 163.367
R343 B.n337 B.n27 163.367
R344 B.n337 B.n336 163.367
R345 B.n336 B.n335 163.367
R346 B.n335 B.n29 163.367
R347 B.n331 B.n29 163.367
R348 B.n331 B.n330 163.367
R349 B.n330 B.n329 163.367
R350 B.n329 B.n31 163.367
R351 B.n324 B.n31 163.367
R352 B.n324 B.n323 163.367
R353 B.n323 B.n322 163.367
R354 B.n322 B.n35 163.367
R355 B.n318 B.n35 163.367
R356 B.n318 B.n317 163.367
R357 B.n317 B.n316 163.367
R358 B.n316 B.n37 163.367
R359 B.n312 B.n37 163.367
R360 B.n312 B.n311 163.367
R361 B.n311 B.n310 163.367
R362 B.n310 B.n39 163.367
R363 B.n306 B.n39 163.367
R364 B.n306 B.n305 163.367
R365 B.n305 B.n304 163.367
R366 B.n304 B.n41 163.367
R367 B.n300 B.n41 163.367
R368 B.n370 B.n15 163.367
R369 B.n371 B.n370 163.367
R370 B.n372 B.n371 163.367
R371 B.n372 B.n13 163.367
R372 B.n376 B.n13 163.367
R373 B.n377 B.n376 163.367
R374 B.n378 B.n377 163.367
R375 B.n378 B.n11 163.367
R376 B.n382 B.n11 163.367
R377 B.n383 B.n382 163.367
R378 B.n384 B.n383 163.367
R379 B.n384 B.n9 163.367
R380 B.n388 B.n9 163.367
R381 B.n389 B.n388 163.367
R382 B.n390 B.n389 163.367
R383 B.n390 B.n7 163.367
R384 B.n394 B.n7 163.367
R385 B.n395 B.n394 163.367
R386 B.n396 B.n395 163.367
R387 B.n396 B.n5 163.367
R388 B.n400 B.n5 163.367
R389 B.n401 B.n400 163.367
R390 B.n402 B.n401 163.367
R391 B.n402 B.n3 163.367
R392 B.n406 B.n3 163.367
R393 B.n407 B.n406 163.367
R394 B.n108 B.n2 163.367
R395 B.n109 B.n108 163.367
R396 B.n110 B.n109 163.367
R397 B.n110 B.n105 163.367
R398 B.n114 B.n105 163.367
R399 B.n115 B.n114 163.367
R400 B.n116 B.n115 163.367
R401 B.n116 B.n103 163.367
R402 B.n120 B.n103 163.367
R403 B.n121 B.n120 163.367
R404 B.n122 B.n121 163.367
R405 B.n122 B.n101 163.367
R406 B.n126 B.n101 163.367
R407 B.n127 B.n126 163.367
R408 B.n128 B.n127 163.367
R409 B.n128 B.n99 163.367
R410 B.n132 B.n99 163.367
R411 B.n133 B.n132 163.367
R412 B.n134 B.n133 163.367
R413 B.n134 B.n97 163.367
R414 B.n138 B.n97 163.367
R415 B.n139 B.n138 163.367
R416 B.n140 B.n139 163.367
R417 B.n140 B.n95 163.367
R418 B.n144 B.n95 163.367
R419 B.n145 B.n144 163.367
R420 B.n187 B.t8 131.332
R421 B.n33 B.t1 131.332
R422 B.n85 B.t11 131.329
R423 B.n25 B.t4 131.329
R424 B.n85 B.n84 63.8066
R425 B.n187 B.n186 63.8066
R426 B.n33 B.n32 63.8066
R427 B.n25 B.n24 63.8066
R428 B.n172 B.n85 59.5399
R429 B.n188 B.n187 59.5399
R430 B.n326 B.n33 59.5399
R431 B.n26 B.n25 59.5399
R432 B.n368 B.n367 31.3761
R433 B.n301 B.n42 31.3761
R434 B.n217 B.n70 31.3761
R435 B.n147 B.n94 31.3761
R436 B B.n409 18.0485
R437 B.n369 B.n368 10.6151
R438 B.n369 B.n14 10.6151
R439 B.n373 B.n14 10.6151
R440 B.n374 B.n373 10.6151
R441 B.n375 B.n374 10.6151
R442 B.n375 B.n12 10.6151
R443 B.n379 B.n12 10.6151
R444 B.n380 B.n379 10.6151
R445 B.n381 B.n380 10.6151
R446 B.n381 B.n10 10.6151
R447 B.n385 B.n10 10.6151
R448 B.n386 B.n385 10.6151
R449 B.n387 B.n386 10.6151
R450 B.n387 B.n8 10.6151
R451 B.n391 B.n8 10.6151
R452 B.n392 B.n391 10.6151
R453 B.n393 B.n392 10.6151
R454 B.n393 B.n6 10.6151
R455 B.n397 B.n6 10.6151
R456 B.n398 B.n397 10.6151
R457 B.n399 B.n398 10.6151
R458 B.n399 B.n4 10.6151
R459 B.n403 B.n4 10.6151
R460 B.n404 B.n403 10.6151
R461 B.n405 B.n404 10.6151
R462 B.n405 B.n0 10.6151
R463 B.n367 B.n16 10.6151
R464 B.n363 B.n16 10.6151
R465 B.n363 B.n362 10.6151
R466 B.n362 B.n361 10.6151
R467 B.n361 B.n18 10.6151
R468 B.n357 B.n18 10.6151
R469 B.n357 B.n356 10.6151
R470 B.n356 B.n355 10.6151
R471 B.n355 B.n20 10.6151
R472 B.n351 B.n20 10.6151
R473 B.n351 B.n350 10.6151
R474 B.n350 B.n349 10.6151
R475 B.n349 B.n22 10.6151
R476 B.n345 B.n22 10.6151
R477 B.n345 B.n344 10.6151
R478 B.n344 B.n343 10.6151
R479 B.n340 B.n339 10.6151
R480 B.n339 B.n338 10.6151
R481 B.n338 B.n28 10.6151
R482 B.n334 B.n28 10.6151
R483 B.n334 B.n333 10.6151
R484 B.n333 B.n332 10.6151
R485 B.n332 B.n30 10.6151
R486 B.n328 B.n30 10.6151
R487 B.n328 B.n327 10.6151
R488 B.n325 B.n34 10.6151
R489 B.n321 B.n34 10.6151
R490 B.n321 B.n320 10.6151
R491 B.n320 B.n319 10.6151
R492 B.n319 B.n36 10.6151
R493 B.n315 B.n36 10.6151
R494 B.n315 B.n314 10.6151
R495 B.n314 B.n313 10.6151
R496 B.n313 B.n38 10.6151
R497 B.n309 B.n38 10.6151
R498 B.n309 B.n308 10.6151
R499 B.n308 B.n307 10.6151
R500 B.n307 B.n40 10.6151
R501 B.n303 B.n40 10.6151
R502 B.n303 B.n302 10.6151
R503 B.n302 B.n301 10.6151
R504 B.n297 B.n42 10.6151
R505 B.n297 B.n296 10.6151
R506 B.n296 B.n295 10.6151
R507 B.n295 B.n44 10.6151
R508 B.n291 B.n44 10.6151
R509 B.n291 B.n290 10.6151
R510 B.n290 B.n289 10.6151
R511 B.n289 B.n46 10.6151
R512 B.n285 B.n46 10.6151
R513 B.n285 B.n284 10.6151
R514 B.n284 B.n283 10.6151
R515 B.n283 B.n48 10.6151
R516 B.n279 B.n48 10.6151
R517 B.n279 B.n278 10.6151
R518 B.n278 B.n277 10.6151
R519 B.n277 B.n50 10.6151
R520 B.n273 B.n50 10.6151
R521 B.n273 B.n272 10.6151
R522 B.n272 B.n271 10.6151
R523 B.n271 B.n52 10.6151
R524 B.n267 B.n52 10.6151
R525 B.n267 B.n266 10.6151
R526 B.n266 B.n265 10.6151
R527 B.n265 B.n54 10.6151
R528 B.n261 B.n54 10.6151
R529 B.n261 B.n260 10.6151
R530 B.n260 B.n259 10.6151
R531 B.n259 B.n56 10.6151
R532 B.n255 B.n56 10.6151
R533 B.n255 B.n254 10.6151
R534 B.n254 B.n253 10.6151
R535 B.n253 B.n58 10.6151
R536 B.n249 B.n58 10.6151
R537 B.n249 B.n248 10.6151
R538 B.n248 B.n247 10.6151
R539 B.n247 B.n60 10.6151
R540 B.n243 B.n60 10.6151
R541 B.n243 B.n242 10.6151
R542 B.n242 B.n241 10.6151
R543 B.n241 B.n62 10.6151
R544 B.n237 B.n62 10.6151
R545 B.n237 B.n236 10.6151
R546 B.n236 B.n235 10.6151
R547 B.n235 B.n64 10.6151
R548 B.n231 B.n64 10.6151
R549 B.n231 B.n230 10.6151
R550 B.n230 B.n229 10.6151
R551 B.n229 B.n66 10.6151
R552 B.n225 B.n66 10.6151
R553 B.n225 B.n224 10.6151
R554 B.n224 B.n223 10.6151
R555 B.n223 B.n68 10.6151
R556 B.n219 B.n68 10.6151
R557 B.n219 B.n218 10.6151
R558 B.n218 B.n217 10.6151
R559 B.n107 B.n1 10.6151
R560 B.n107 B.n106 10.6151
R561 B.n111 B.n106 10.6151
R562 B.n112 B.n111 10.6151
R563 B.n113 B.n112 10.6151
R564 B.n113 B.n104 10.6151
R565 B.n117 B.n104 10.6151
R566 B.n118 B.n117 10.6151
R567 B.n119 B.n118 10.6151
R568 B.n119 B.n102 10.6151
R569 B.n123 B.n102 10.6151
R570 B.n124 B.n123 10.6151
R571 B.n125 B.n124 10.6151
R572 B.n125 B.n100 10.6151
R573 B.n129 B.n100 10.6151
R574 B.n130 B.n129 10.6151
R575 B.n131 B.n130 10.6151
R576 B.n131 B.n98 10.6151
R577 B.n135 B.n98 10.6151
R578 B.n136 B.n135 10.6151
R579 B.n137 B.n136 10.6151
R580 B.n137 B.n96 10.6151
R581 B.n141 B.n96 10.6151
R582 B.n142 B.n141 10.6151
R583 B.n143 B.n142 10.6151
R584 B.n143 B.n94 10.6151
R585 B.n148 B.n147 10.6151
R586 B.n149 B.n148 10.6151
R587 B.n149 B.n92 10.6151
R588 B.n153 B.n92 10.6151
R589 B.n154 B.n153 10.6151
R590 B.n155 B.n154 10.6151
R591 B.n155 B.n90 10.6151
R592 B.n159 B.n90 10.6151
R593 B.n160 B.n159 10.6151
R594 B.n161 B.n160 10.6151
R595 B.n161 B.n88 10.6151
R596 B.n165 B.n88 10.6151
R597 B.n166 B.n165 10.6151
R598 B.n167 B.n166 10.6151
R599 B.n167 B.n86 10.6151
R600 B.n171 B.n86 10.6151
R601 B.n174 B.n173 10.6151
R602 B.n174 B.n82 10.6151
R603 B.n178 B.n82 10.6151
R604 B.n179 B.n178 10.6151
R605 B.n180 B.n179 10.6151
R606 B.n180 B.n80 10.6151
R607 B.n184 B.n80 10.6151
R608 B.n185 B.n184 10.6151
R609 B.n189 B.n185 10.6151
R610 B.n193 B.n78 10.6151
R611 B.n194 B.n193 10.6151
R612 B.n195 B.n194 10.6151
R613 B.n195 B.n76 10.6151
R614 B.n199 B.n76 10.6151
R615 B.n200 B.n199 10.6151
R616 B.n201 B.n200 10.6151
R617 B.n201 B.n74 10.6151
R618 B.n205 B.n74 10.6151
R619 B.n206 B.n205 10.6151
R620 B.n207 B.n206 10.6151
R621 B.n207 B.n72 10.6151
R622 B.n211 B.n72 10.6151
R623 B.n212 B.n211 10.6151
R624 B.n213 B.n212 10.6151
R625 B.n213 B.n70 10.6151
R626 B.n343 B.n26 9.36635
R627 B.n326 B.n325 9.36635
R628 B.n172 B.n171 9.36635
R629 B.n188 B.n78 9.36635
R630 B.n409 B.n0 8.11757
R631 B.n409 B.n1 8.11757
R632 B.n340 B.n26 1.24928
R633 B.n327 B.n326 1.24928
R634 B.n173 B.n172 1.24928
R635 B.n189 B.n188 1.24928
R636 VN VN.t0 110.41
R637 VN VN.t1 71.5317
R638 VDD2.n0 VDD2.t0 165.125
R639 VDD2.n0 VDD2.t1 132.619
R640 VDD2 VDD2.n0 0.767741
C0 VDD1 w_n2286_n1704# 1.24492f
C1 VTAIL B 1.84139f
C2 VN VP 4.08553f
C3 VDD1 VN 0.153084f
C4 VDD2 VP 0.35281f
C5 VDD2 VDD1 0.717407f
C6 VP B 1.48609f
C7 VN w_n2286_n1704# 3.02341f
C8 VDD1 B 1.09091f
C9 VDD2 w_n2286_n1704# 1.27484f
C10 VTAIL VP 1.2631f
C11 VDD1 VTAIL 2.97485f
C12 VDD2 VN 1.04699f
C13 B w_n2286_n1704# 6.88403f
C14 VTAIL w_n2286_n1704# 1.57871f
C15 VN B 1.0049f
C16 VDD1 VP 1.2452f
C17 VDD2 B 1.12438f
C18 VTAIL VN 1.24894f
C19 VDD2 VTAIL 3.02993f
C20 VP w_n2286_n1704# 3.31406f
C21 VDD2 VSUBS 0.620568f
C22 VDD1 VSUBS 2.86849f
C23 VTAIL VSUBS 0.436531f
C24 VN VSUBS 5.48807f
C25 VP VSUBS 1.351315f
C26 B VSUBS 3.291311f
C27 w_n2286_n1704# VSUBS 49.1307f
C28 VDD2.t0 VSUBS 0.547296f
C29 VDD2.t1 VSUBS 0.368504f
C30 VDD2.n0 VSUBS 1.97087f
C31 VN.t1 VSUBS 1.52221f
C32 VN.t0 VSUBS 2.22982f
C33 B.n0 VSUBS 0.006463f
C34 B.n1 VSUBS 0.006463f
C35 B.n2 VSUBS 0.009559f
C36 B.n3 VSUBS 0.007325f
C37 B.n4 VSUBS 0.007325f
C38 B.n5 VSUBS 0.007325f
C39 B.n6 VSUBS 0.007325f
C40 B.n7 VSUBS 0.007325f
C41 B.n8 VSUBS 0.007325f
C42 B.n9 VSUBS 0.007325f
C43 B.n10 VSUBS 0.007325f
C44 B.n11 VSUBS 0.007325f
C45 B.n12 VSUBS 0.007325f
C46 B.n13 VSUBS 0.007325f
C47 B.n14 VSUBS 0.007325f
C48 B.n15 VSUBS 0.016246f
C49 B.n16 VSUBS 0.007325f
C50 B.n17 VSUBS 0.007325f
C51 B.n18 VSUBS 0.007325f
C52 B.n19 VSUBS 0.007325f
C53 B.n20 VSUBS 0.007325f
C54 B.n21 VSUBS 0.007325f
C55 B.n22 VSUBS 0.007325f
C56 B.n23 VSUBS 0.007325f
C57 B.t4 VSUBS 0.098384f
C58 B.t5 VSUBS 0.118755f
C59 B.t3 VSUBS 0.552511f
C60 B.n24 VSUBS 0.096036f
C61 B.n25 VSUBS 0.072748f
C62 B.n26 VSUBS 0.016971f
C63 B.n27 VSUBS 0.007325f
C64 B.n28 VSUBS 0.007325f
C65 B.n29 VSUBS 0.007325f
C66 B.n30 VSUBS 0.007325f
C67 B.n31 VSUBS 0.007325f
C68 B.t1 VSUBS 0.098384f
C69 B.t2 VSUBS 0.118755f
C70 B.t0 VSUBS 0.552511f
C71 B.n32 VSUBS 0.096036f
C72 B.n33 VSUBS 0.072748f
C73 B.n34 VSUBS 0.007325f
C74 B.n35 VSUBS 0.007325f
C75 B.n36 VSUBS 0.007325f
C76 B.n37 VSUBS 0.007325f
C77 B.n38 VSUBS 0.007325f
C78 B.n39 VSUBS 0.007325f
C79 B.n40 VSUBS 0.007325f
C80 B.n41 VSUBS 0.007325f
C81 B.n42 VSUBS 0.016246f
C82 B.n43 VSUBS 0.007325f
C83 B.n44 VSUBS 0.007325f
C84 B.n45 VSUBS 0.007325f
C85 B.n46 VSUBS 0.007325f
C86 B.n47 VSUBS 0.007325f
C87 B.n48 VSUBS 0.007325f
C88 B.n49 VSUBS 0.007325f
C89 B.n50 VSUBS 0.007325f
C90 B.n51 VSUBS 0.007325f
C91 B.n52 VSUBS 0.007325f
C92 B.n53 VSUBS 0.007325f
C93 B.n54 VSUBS 0.007325f
C94 B.n55 VSUBS 0.007325f
C95 B.n56 VSUBS 0.007325f
C96 B.n57 VSUBS 0.007325f
C97 B.n58 VSUBS 0.007325f
C98 B.n59 VSUBS 0.007325f
C99 B.n60 VSUBS 0.007325f
C100 B.n61 VSUBS 0.007325f
C101 B.n62 VSUBS 0.007325f
C102 B.n63 VSUBS 0.007325f
C103 B.n64 VSUBS 0.007325f
C104 B.n65 VSUBS 0.007325f
C105 B.n66 VSUBS 0.007325f
C106 B.n67 VSUBS 0.007325f
C107 B.n68 VSUBS 0.007325f
C108 B.n69 VSUBS 0.007325f
C109 B.n70 VSUBS 0.016246f
C110 B.n71 VSUBS 0.007325f
C111 B.n72 VSUBS 0.007325f
C112 B.n73 VSUBS 0.007325f
C113 B.n74 VSUBS 0.007325f
C114 B.n75 VSUBS 0.007325f
C115 B.n76 VSUBS 0.007325f
C116 B.n77 VSUBS 0.007325f
C117 B.n78 VSUBS 0.006894f
C118 B.n79 VSUBS 0.007325f
C119 B.n80 VSUBS 0.007325f
C120 B.n81 VSUBS 0.007325f
C121 B.n82 VSUBS 0.007325f
C122 B.n83 VSUBS 0.007325f
C123 B.t11 VSUBS 0.098384f
C124 B.t10 VSUBS 0.118755f
C125 B.t9 VSUBS 0.552511f
C126 B.n84 VSUBS 0.096036f
C127 B.n85 VSUBS 0.072748f
C128 B.n86 VSUBS 0.007325f
C129 B.n87 VSUBS 0.007325f
C130 B.n88 VSUBS 0.007325f
C131 B.n89 VSUBS 0.007325f
C132 B.n90 VSUBS 0.007325f
C133 B.n91 VSUBS 0.007325f
C134 B.n92 VSUBS 0.007325f
C135 B.n93 VSUBS 0.007325f
C136 B.n94 VSUBS 0.016246f
C137 B.n95 VSUBS 0.007325f
C138 B.n96 VSUBS 0.007325f
C139 B.n97 VSUBS 0.007325f
C140 B.n98 VSUBS 0.007325f
C141 B.n99 VSUBS 0.007325f
C142 B.n100 VSUBS 0.007325f
C143 B.n101 VSUBS 0.007325f
C144 B.n102 VSUBS 0.007325f
C145 B.n103 VSUBS 0.007325f
C146 B.n104 VSUBS 0.007325f
C147 B.n105 VSUBS 0.007325f
C148 B.n106 VSUBS 0.007325f
C149 B.n107 VSUBS 0.007325f
C150 B.n108 VSUBS 0.007325f
C151 B.n109 VSUBS 0.007325f
C152 B.n110 VSUBS 0.007325f
C153 B.n111 VSUBS 0.007325f
C154 B.n112 VSUBS 0.007325f
C155 B.n113 VSUBS 0.007325f
C156 B.n114 VSUBS 0.007325f
C157 B.n115 VSUBS 0.007325f
C158 B.n116 VSUBS 0.007325f
C159 B.n117 VSUBS 0.007325f
C160 B.n118 VSUBS 0.007325f
C161 B.n119 VSUBS 0.007325f
C162 B.n120 VSUBS 0.007325f
C163 B.n121 VSUBS 0.007325f
C164 B.n122 VSUBS 0.007325f
C165 B.n123 VSUBS 0.007325f
C166 B.n124 VSUBS 0.007325f
C167 B.n125 VSUBS 0.007325f
C168 B.n126 VSUBS 0.007325f
C169 B.n127 VSUBS 0.007325f
C170 B.n128 VSUBS 0.007325f
C171 B.n129 VSUBS 0.007325f
C172 B.n130 VSUBS 0.007325f
C173 B.n131 VSUBS 0.007325f
C174 B.n132 VSUBS 0.007325f
C175 B.n133 VSUBS 0.007325f
C176 B.n134 VSUBS 0.007325f
C177 B.n135 VSUBS 0.007325f
C178 B.n136 VSUBS 0.007325f
C179 B.n137 VSUBS 0.007325f
C180 B.n138 VSUBS 0.007325f
C181 B.n139 VSUBS 0.007325f
C182 B.n140 VSUBS 0.007325f
C183 B.n141 VSUBS 0.007325f
C184 B.n142 VSUBS 0.007325f
C185 B.n143 VSUBS 0.007325f
C186 B.n144 VSUBS 0.007325f
C187 B.n145 VSUBS 0.016246f
C188 B.n146 VSUBS 0.017147f
C189 B.n147 VSUBS 0.017147f
C190 B.n148 VSUBS 0.007325f
C191 B.n149 VSUBS 0.007325f
C192 B.n150 VSUBS 0.007325f
C193 B.n151 VSUBS 0.007325f
C194 B.n152 VSUBS 0.007325f
C195 B.n153 VSUBS 0.007325f
C196 B.n154 VSUBS 0.007325f
C197 B.n155 VSUBS 0.007325f
C198 B.n156 VSUBS 0.007325f
C199 B.n157 VSUBS 0.007325f
C200 B.n158 VSUBS 0.007325f
C201 B.n159 VSUBS 0.007325f
C202 B.n160 VSUBS 0.007325f
C203 B.n161 VSUBS 0.007325f
C204 B.n162 VSUBS 0.007325f
C205 B.n163 VSUBS 0.007325f
C206 B.n164 VSUBS 0.007325f
C207 B.n165 VSUBS 0.007325f
C208 B.n166 VSUBS 0.007325f
C209 B.n167 VSUBS 0.007325f
C210 B.n168 VSUBS 0.007325f
C211 B.n169 VSUBS 0.007325f
C212 B.n170 VSUBS 0.007325f
C213 B.n171 VSUBS 0.006894f
C214 B.n172 VSUBS 0.016971f
C215 B.n173 VSUBS 0.004093f
C216 B.n174 VSUBS 0.007325f
C217 B.n175 VSUBS 0.007325f
C218 B.n176 VSUBS 0.007325f
C219 B.n177 VSUBS 0.007325f
C220 B.n178 VSUBS 0.007325f
C221 B.n179 VSUBS 0.007325f
C222 B.n180 VSUBS 0.007325f
C223 B.n181 VSUBS 0.007325f
C224 B.n182 VSUBS 0.007325f
C225 B.n183 VSUBS 0.007325f
C226 B.n184 VSUBS 0.007325f
C227 B.n185 VSUBS 0.007325f
C228 B.t8 VSUBS 0.098384f
C229 B.t7 VSUBS 0.118755f
C230 B.t6 VSUBS 0.552511f
C231 B.n186 VSUBS 0.096036f
C232 B.n187 VSUBS 0.072748f
C233 B.n188 VSUBS 0.016971f
C234 B.n189 VSUBS 0.004093f
C235 B.n190 VSUBS 0.007325f
C236 B.n191 VSUBS 0.007325f
C237 B.n192 VSUBS 0.007325f
C238 B.n193 VSUBS 0.007325f
C239 B.n194 VSUBS 0.007325f
C240 B.n195 VSUBS 0.007325f
C241 B.n196 VSUBS 0.007325f
C242 B.n197 VSUBS 0.007325f
C243 B.n198 VSUBS 0.007325f
C244 B.n199 VSUBS 0.007325f
C245 B.n200 VSUBS 0.007325f
C246 B.n201 VSUBS 0.007325f
C247 B.n202 VSUBS 0.007325f
C248 B.n203 VSUBS 0.007325f
C249 B.n204 VSUBS 0.007325f
C250 B.n205 VSUBS 0.007325f
C251 B.n206 VSUBS 0.007325f
C252 B.n207 VSUBS 0.007325f
C253 B.n208 VSUBS 0.007325f
C254 B.n209 VSUBS 0.007325f
C255 B.n210 VSUBS 0.007325f
C256 B.n211 VSUBS 0.007325f
C257 B.n212 VSUBS 0.007325f
C258 B.n213 VSUBS 0.007325f
C259 B.n214 VSUBS 0.007325f
C260 B.n215 VSUBS 0.017147f
C261 B.n216 VSUBS 0.016246f
C262 B.n217 VSUBS 0.017147f
C263 B.n218 VSUBS 0.007325f
C264 B.n219 VSUBS 0.007325f
C265 B.n220 VSUBS 0.007325f
C266 B.n221 VSUBS 0.007325f
C267 B.n222 VSUBS 0.007325f
C268 B.n223 VSUBS 0.007325f
C269 B.n224 VSUBS 0.007325f
C270 B.n225 VSUBS 0.007325f
C271 B.n226 VSUBS 0.007325f
C272 B.n227 VSUBS 0.007325f
C273 B.n228 VSUBS 0.007325f
C274 B.n229 VSUBS 0.007325f
C275 B.n230 VSUBS 0.007325f
C276 B.n231 VSUBS 0.007325f
C277 B.n232 VSUBS 0.007325f
C278 B.n233 VSUBS 0.007325f
C279 B.n234 VSUBS 0.007325f
C280 B.n235 VSUBS 0.007325f
C281 B.n236 VSUBS 0.007325f
C282 B.n237 VSUBS 0.007325f
C283 B.n238 VSUBS 0.007325f
C284 B.n239 VSUBS 0.007325f
C285 B.n240 VSUBS 0.007325f
C286 B.n241 VSUBS 0.007325f
C287 B.n242 VSUBS 0.007325f
C288 B.n243 VSUBS 0.007325f
C289 B.n244 VSUBS 0.007325f
C290 B.n245 VSUBS 0.007325f
C291 B.n246 VSUBS 0.007325f
C292 B.n247 VSUBS 0.007325f
C293 B.n248 VSUBS 0.007325f
C294 B.n249 VSUBS 0.007325f
C295 B.n250 VSUBS 0.007325f
C296 B.n251 VSUBS 0.007325f
C297 B.n252 VSUBS 0.007325f
C298 B.n253 VSUBS 0.007325f
C299 B.n254 VSUBS 0.007325f
C300 B.n255 VSUBS 0.007325f
C301 B.n256 VSUBS 0.007325f
C302 B.n257 VSUBS 0.007325f
C303 B.n258 VSUBS 0.007325f
C304 B.n259 VSUBS 0.007325f
C305 B.n260 VSUBS 0.007325f
C306 B.n261 VSUBS 0.007325f
C307 B.n262 VSUBS 0.007325f
C308 B.n263 VSUBS 0.007325f
C309 B.n264 VSUBS 0.007325f
C310 B.n265 VSUBS 0.007325f
C311 B.n266 VSUBS 0.007325f
C312 B.n267 VSUBS 0.007325f
C313 B.n268 VSUBS 0.007325f
C314 B.n269 VSUBS 0.007325f
C315 B.n270 VSUBS 0.007325f
C316 B.n271 VSUBS 0.007325f
C317 B.n272 VSUBS 0.007325f
C318 B.n273 VSUBS 0.007325f
C319 B.n274 VSUBS 0.007325f
C320 B.n275 VSUBS 0.007325f
C321 B.n276 VSUBS 0.007325f
C322 B.n277 VSUBS 0.007325f
C323 B.n278 VSUBS 0.007325f
C324 B.n279 VSUBS 0.007325f
C325 B.n280 VSUBS 0.007325f
C326 B.n281 VSUBS 0.007325f
C327 B.n282 VSUBS 0.007325f
C328 B.n283 VSUBS 0.007325f
C329 B.n284 VSUBS 0.007325f
C330 B.n285 VSUBS 0.007325f
C331 B.n286 VSUBS 0.007325f
C332 B.n287 VSUBS 0.007325f
C333 B.n288 VSUBS 0.007325f
C334 B.n289 VSUBS 0.007325f
C335 B.n290 VSUBS 0.007325f
C336 B.n291 VSUBS 0.007325f
C337 B.n292 VSUBS 0.007325f
C338 B.n293 VSUBS 0.007325f
C339 B.n294 VSUBS 0.007325f
C340 B.n295 VSUBS 0.007325f
C341 B.n296 VSUBS 0.007325f
C342 B.n297 VSUBS 0.007325f
C343 B.n298 VSUBS 0.007325f
C344 B.n299 VSUBS 0.016246f
C345 B.n300 VSUBS 0.017147f
C346 B.n301 VSUBS 0.017147f
C347 B.n302 VSUBS 0.007325f
C348 B.n303 VSUBS 0.007325f
C349 B.n304 VSUBS 0.007325f
C350 B.n305 VSUBS 0.007325f
C351 B.n306 VSUBS 0.007325f
C352 B.n307 VSUBS 0.007325f
C353 B.n308 VSUBS 0.007325f
C354 B.n309 VSUBS 0.007325f
C355 B.n310 VSUBS 0.007325f
C356 B.n311 VSUBS 0.007325f
C357 B.n312 VSUBS 0.007325f
C358 B.n313 VSUBS 0.007325f
C359 B.n314 VSUBS 0.007325f
C360 B.n315 VSUBS 0.007325f
C361 B.n316 VSUBS 0.007325f
C362 B.n317 VSUBS 0.007325f
C363 B.n318 VSUBS 0.007325f
C364 B.n319 VSUBS 0.007325f
C365 B.n320 VSUBS 0.007325f
C366 B.n321 VSUBS 0.007325f
C367 B.n322 VSUBS 0.007325f
C368 B.n323 VSUBS 0.007325f
C369 B.n324 VSUBS 0.007325f
C370 B.n325 VSUBS 0.006894f
C371 B.n326 VSUBS 0.016971f
C372 B.n327 VSUBS 0.004093f
C373 B.n328 VSUBS 0.007325f
C374 B.n329 VSUBS 0.007325f
C375 B.n330 VSUBS 0.007325f
C376 B.n331 VSUBS 0.007325f
C377 B.n332 VSUBS 0.007325f
C378 B.n333 VSUBS 0.007325f
C379 B.n334 VSUBS 0.007325f
C380 B.n335 VSUBS 0.007325f
C381 B.n336 VSUBS 0.007325f
C382 B.n337 VSUBS 0.007325f
C383 B.n338 VSUBS 0.007325f
C384 B.n339 VSUBS 0.007325f
C385 B.n340 VSUBS 0.004093f
C386 B.n341 VSUBS 0.007325f
C387 B.n342 VSUBS 0.007325f
C388 B.n343 VSUBS 0.006894f
C389 B.n344 VSUBS 0.007325f
C390 B.n345 VSUBS 0.007325f
C391 B.n346 VSUBS 0.007325f
C392 B.n347 VSUBS 0.007325f
C393 B.n348 VSUBS 0.007325f
C394 B.n349 VSUBS 0.007325f
C395 B.n350 VSUBS 0.007325f
C396 B.n351 VSUBS 0.007325f
C397 B.n352 VSUBS 0.007325f
C398 B.n353 VSUBS 0.007325f
C399 B.n354 VSUBS 0.007325f
C400 B.n355 VSUBS 0.007325f
C401 B.n356 VSUBS 0.007325f
C402 B.n357 VSUBS 0.007325f
C403 B.n358 VSUBS 0.007325f
C404 B.n359 VSUBS 0.007325f
C405 B.n360 VSUBS 0.007325f
C406 B.n361 VSUBS 0.007325f
C407 B.n362 VSUBS 0.007325f
C408 B.n363 VSUBS 0.007325f
C409 B.n364 VSUBS 0.007325f
C410 B.n365 VSUBS 0.007325f
C411 B.n366 VSUBS 0.017147f
C412 B.n367 VSUBS 0.017147f
C413 B.n368 VSUBS 0.016246f
C414 B.n369 VSUBS 0.007325f
C415 B.n370 VSUBS 0.007325f
C416 B.n371 VSUBS 0.007325f
C417 B.n372 VSUBS 0.007325f
C418 B.n373 VSUBS 0.007325f
C419 B.n374 VSUBS 0.007325f
C420 B.n375 VSUBS 0.007325f
C421 B.n376 VSUBS 0.007325f
C422 B.n377 VSUBS 0.007325f
C423 B.n378 VSUBS 0.007325f
C424 B.n379 VSUBS 0.007325f
C425 B.n380 VSUBS 0.007325f
C426 B.n381 VSUBS 0.007325f
C427 B.n382 VSUBS 0.007325f
C428 B.n383 VSUBS 0.007325f
C429 B.n384 VSUBS 0.007325f
C430 B.n385 VSUBS 0.007325f
C431 B.n386 VSUBS 0.007325f
C432 B.n387 VSUBS 0.007325f
C433 B.n388 VSUBS 0.007325f
C434 B.n389 VSUBS 0.007325f
C435 B.n390 VSUBS 0.007325f
C436 B.n391 VSUBS 0.007325f
C437 B.n392 VSUBS 0.007325f
C438 B.n393 VSUBS 0.007325f
C439 B.n394 VSUBS 0.007325f
C440 B.n395 VSUBS 0.007325f
C441 B.n396 VSUBS 0.007325f
C442 B.n397 VSUBS 0.007325f
C443 B.n398 VSUBS 0.007325f
C444 B.n399 VSUBS 0.007325f
C445 B.n400 VSUBS 0.007325f
C446 B.n401 VSUBS 0.007325f
C447 B.n402 VSUBS 0.007325f
C448 B.n403 VSUBS 0.007325f
C449 B.n404 VSUBS 0.007325f
C450 B.n405 VSUBS 0.007325f
C451 B.n406 VSUBS 0.007325f
C452 B.n407 VSUBS 0.009559f
C453 B.n408 VSUBS 0.010182f
C454 B.n409 VSUBS 0.020249f
C455 VDD1.t0 VSUBS 0.363002f
C456 VDD1.t1 VSUBS 0.552662f
C457 VTAIL.t2 VSUBS 0.388741f
C458 VTAIL.n0 VSUBS 1.15739f
C459 VTAIL.t3 VSUBS 0.388743f
C460 VTAIL.n1 VSUBS 1.19652f
C461 VTAIL.t1 VSUBS 0.388741f
C462 VTAIL.n2 VSUBS 1.02599f
C463 VTAIL.t0 VSUBS 0.388741f
C464 VTAIL.n3 VSUBS 0.95161f
C465 VP.t0 VSUBS 1.59576f
C466 VP.t1 VSUBS 2.33817f
C467 VP.n0 VSUBS 3.34427f
.ends

