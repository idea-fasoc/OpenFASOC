* NGSPICE file created from diff_pair_sample_1575.ext - technology: sky130A

.subckt diff_pair_sample_1575 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VN.t0 VDD2.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.8892 pd=5.34 as=0.3762 ps=2.61 w=2.28 l=1.88
X1 B.t17 B.t15 B.t16 B.t5 sky130_fd_pr__nfet_01v8 ad=0.8892 pd=5.34 as=0 ps=0 w=2.28 l=1.88
X2 VTAIL.t0 VP.t0 VDD1.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=0.8892 pd=5.34 as=0.3762 ps=2.61 w=2.28 l=1.88
X3 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=0.8892 pd=5.34 as=0 ps=0 w=2.28 l=1.88
X4 VDD1.t2 VP.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.3762 pd=2.61 as=0.8892 ps=5.34 w=2.28 l=1.88
X5 VDD2.t1 VN.t1 VTAIL.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=0.3762 pd=2.61 as=0.8892 ps=5.34 w=2.28 l=1.88
X6 VDD1.t1 VP.t2 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.3762 pd=2.61 as=0.8892 ps=5.34 w=2.28 l=1.88
X7 VDD2.t3 VN.t2 VTAIL.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=0.3762 pd=2.61 as=0.8892 ps=5.34 w=2.28 l=1.88
X8 VTAIL.t4 VN.t3 VDD2.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.8892 pd=5.34 as=0.3762 ps=2.61 w=2.28 l=1.88
X9 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=0.8892 pd=5.34 as=0 ps=0 w=2.28 l=1.88
X10 VTAIL.t2 VP.t3 VDD1.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=0.8892 pd=5.34 as=0.3762 ps=2.61 w=2.28 l=1.88
X11 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=0.8892 pd=5.34 as=0 ps=0 w=2.28 l=1.88
R0 VN.n0 VN.t0 67.0251
R1 VN.n1 VN.t2 67.0251
R2 VN.n0 VN.t1 66.586
R3 VN.n1 VN.t3 66.586
R4 VN VN.n1 46.1902
R5 VN VN.n0 9.10304
R6 VDD2.n2 VDD2.n0 126.802
R7 VDD2.n2 VDD2.n1 95.407
R8 VDD2.n1 VDD2.t2 8.68471
R9 VDD2.n1 VDD2.t3 8.68471
R10 VDD2.n0 VDD2.t0 8.68471
R11 VDD2.n0 VDD2.t1 8.68471
R12 VDD2 VDD2.n2 0.0586897
R13 VTAIL.n7 VTAIL.t6 87.4124
R14 VTAIL.n0 VTAIL.t7 87.4124
R15 VTAIL.n1 VTAIL.t3 87.4124
R16 VTAIL.n2 VTAIL.t2 87.4124
R17 VTAIL.n6 VTAIL.t1 87.4124
R18 VTAIL.n5 VTAIL.t0 87.4123
R19 VTAIL.n4 VTAIL.t5 87.4123
R20 VTAIL.n3 VTAIL.t4 87.4123
R21 VTAIL.n7 VTAIL.n6 16.2376
R22 VTAIL.n3 VTAIL.n2 16.2376
R23 VTAIL.n4 VTAIL.n3 1.90567
R24 VTAIL.n6 VTAIL.n5 1.90567
R25 VTAIL.n2 VTAIL.n1 1.90567
R26 VTAIL VTAIL.n0 1.01128
R27 VTAIL VTAIL.n7 0.894897
R28 VTAIL.n5 VTAIL.n4 0.470328
R29 VTAIL.n1 VTAIL.n0 0.470328
R30 B.n409 B.n408 585
R31 B.n143 B.n71 585
R32 B.n142 B.n141 585
R33 B.n140 B.n139 585
R34 B.n138 B.n137 585
R35 B.n136 B.n135 585
R36 B.n134 B.n133 585
R37 B.n132 B.n131 585
R38 B.n130 B.n129 585
R39 B.n128 B.n127 585
R40 B.n126 B.n125 585
R41 B.n124 B.n123 585
R42 B.n122 B.n121 585
R43 B.n119 B.n118 585
R44 B.n117 B.n116 585
R45 B.n115 B.n114 585
R46 B.n113 B.n112 585
R47 B.n111 B.n110 585
R48 B.n109 B.n108 585
R49 B.n107 B.n106 585
R50 B.n105 B.n104 585
R51 B.n103 B.n102 585
R52 B.n101 B.n100 585
R53 B.n98 B.n97 585
R54 B.n96 B.n95 585
R55 B.n94 B.n93 585
R56 B.n92 B.n91 585
R57 B.n90 B.n89 585
R58 B.n88 B.n87 585
R59 B.n86 B.n85 585
R60 B.n84 B.n83 585
R61 B.n82 B.n81 585
R62 B.n80 B.n79 585
R63 B.n78 B.n77 585
R64 B.n54 B.n53 585
R65 B.n414 B.n413 585
R66 B.n407 B.n72 585
R67 B.n72 B.n51 585
R68 B.n406 B.n50 585
R69 B.n418 B.n50 585
R70 B.n405 B.n49 585
R71 B.n419 B.n49 585
R72 B.n404 B.n48 585
R73 B.n420 B.n48 585
R74 B.n403 B.n402 585
R75 B.n402 B.n44 585
R76 B.n401 B.n43 585
R77 B.n426 B.n43 585
R78 B.n400 B.n42 585
R79 B.n427 B.n42 585
R80 B.n399 B.n41 585
R81 B.n428 B.n41 585
R82 B.n398 B.n397 585
R83 B.n397 B.n37 585
R84 B.n396 B.n36 585
R85 B.n434 B.n36 585
R86 B.n395 B.n35 585
R87 B.n435 B.n35 585
R88 B.n394 B.n34 585
R89 B.n436 B.n34 585
R90 B.n393 B.n392 585
R91 B.n392 B.n30 585
R92 B.n391 B.n29 585
R93 B.n442 B.n29 585
R94 B.n390 B.n28 585
R95 B.n443 B.n28 585
R96 B.n389 B.n27 585
R97 B.n444 B.n27 585
R98 B.n388 B.n387 585
R99 B.n387 B.n26 585
R100 B.n386 B.n22 585
R101 B.n450 B.n22 585
R102 B.n385 B.n21 585
R103 B.n451 B.n21 585
R104 B.n384 B.n20 585
R105 B.n452 B.n20 585
R106 B.n383 B.n382 585
R107 B.n382 B.n16 585
R108 B.n381 B.n15 585
R109 B.n458 B.n15 585
R110 B.n380 B.n14 585
R111 B.n459 B.n14 585
R112 B.n379 B.n13 585
R113 B.n460 B.n13 585
R114 B.n378 B.n377 585
R115 B.n377 B.n12 585
R116 B.n376 B.n375 585
R117 B.n376 B.n8 585
R118 B.n374 B.n7 585
R119 B.n467 B.n7 585
R120 B.n373 B.n6 585
R121 B.n468 B.n6 585
R122 B.n372 B.n5 585
R123 B.n469 B.n5 585
R124 B.n371 B.n370 585
R125 B.n370 B.n4 585
R126 B.n369 B.n144 585
R127 B.n369 B.n368 585
R128 B.n359 B.n145 585
R129 B.n146 B.n145 585
R130 B.n361 B.n360 585
R131 B.n362 B.n361 585
R132 B.n358 B.n150 585
R133 B.n154 B.n150 585
R134 B.n357 B.n356 585
R135 B.n356 B.n355 585
R136 B.n152 B.n151 585
R137 B.n153 B.n152 585
R138 B.n348 B.n347 585
R139 B.n349 B.n348 585
R140 B.n346 B.n159 585
R141 B.n159 B.n158 585
R142 B.n345 B.n344 585
R143 B.n344 B.n343 585
R144 B.n161 B.n160 585
R145 B.n336 B.n161 585
R146 B.n335 B.n334 585
R147 B.n337 B.n335 585
R148 B.n333 B.n166 585
R149 B.n166 B.n165 585
R150 B.n332 B.n331 585
R151 B.n331 B.n330 585
R152 B.n168 B.n167 585
R153 B.n169 B.n168 585
R154 B.n323 B.n322 585
R155 B.n324 B.n323 585
R156 B.n321 B.n174 585
R157 B.n174 B.n173 585
R158 B.n320 B.n319 585
R159 B.n319 B.n318 585
R160 B.n176 B.n175 585
R161 B.n177 B.n176 585
R162 B.n311 B.n310 585
R163 B.n312 B.n311 585
R164 B.n309 B.n181 585
R165 B.n185 B.n181 585
R166 B.n308 B.n307 585
R167 B.n307 B.n306 585
R168 B.n183 B.n182 585
R169 B.n184 B.n183 585
R170 B.n299 B.n298 585
R171 B.n300 B.n299 585
R172 B.n297 B.n190 585
R173 B.n190 B.n189 585
R174 B.n296 B.n295 585
R175 B.n295 B.n294 585
R176 B.n192 B.n191 585
R177 B.n193 B.n192 585
R178 B.n290 B.n289 585
R179 B.n196 B.n195 585
R180 B.n286 B.n285 585
R181 B.n287 B.n286 585
R182 B.n284 B.n214 585
R183 B.n283 B.n282 585
R184 B.n281 B.n280 585
R185 B.n279 B.n278 585
R186 B.n277 B.n276 585
R187 B.n275 B.n274 585
R188 B.n273 B.n272 585
R189 B.n271 B.n270 585
R190 B.n269 B.n268 585
R191 B.n267 B.n266 585
R192 B.n265 B.n264 585
R193 B.n263 B.n262 585
R194 B.n261 B.n260 585
R195 B.n259 B.n258 585
R196 B.n257 B.n256 585
R197 B.n255 B.n254 585
R198 B.n253 B.n252 585
R199 B.n251 B.n250 585
R200 B.n249 B.n248 585
R201 B.n247 B.n246 585
R202 B.n245 B.n244 585
R203 B.n243 B.n242 585
R204 B.n241 B.n240 585
R205 B.n239 B.n238 585
R206 B.n237 B.n236 585
R207 B.n235 B.n234 585
R208 B.n233 B.n232 585
R209 B.n231 B.n230 585
R210 B.n229 B.n228 585
R211 B.n227 B.n226 585
R212 B.n225 B.n224 585
R213 B.n223 B.n222 585
R214 B.n221 B.n213 585
R215 B.n287 B.n213 585
R216 B.n291 B.n194 585
R217 B.n194 B.n193 585
R218 B.n293 B.n292 585
R219 B.n294 B.n293 585
R220 B.n188 B.n187 585
R221 B.n189 B.n188 585
R222 B.n302 B.n301 585
R223 B.n301 B.n300 585
R224 B.n303 B.n186 585
R225 B.n186 B.n184 585
R226 B.n305 B.n304 585
R227 B.n306 B.n305 585
R228 B.n180 B.n179 585
R229 B.n185 B.n180 585
R230 B.n314 B.n313 585
R231 B.n313 B.n312 585
R232 B.n315 B.n178 585
R233 B.n178 B.n177 585
R234 B.n317 B.n316 585
R235 B.n318 B.n317 585
R236 B.n172 B.n171 585
R237 B.n173 B.n172 585
R238 B.n326 B.n325 585
R239 B.n325 B.n324 585
R240 B.n327 B.n170 585
R241 B.n170 B.n169 585
R242 B.n329 B.n328 585
R243 B.n330 B.n329 585
R244 B.n164 B.n163 585
R245 B.n165 B.n164 585
R246 B.n339 B.n338 585
R247 B.n338 B.n337 585
R248 B.n340 B.n162 585
R249 B.n336 B.n162 585
R250 B.n342 B.n341 585
R251 B.n343 B.n342 585
R252 B.n157 B.n156 585
R253 B.n158 B.n157 585
R254 B.n351 B.n350 585
R255 B.n350 B.n349 585
R256 B.n352 B.n155 585
R257 B.n155 B.n153 585
R258 B.n354 B.n353 585
R259 B.n355 B.n354 585
R260 B.n149 B.n148 585
R261 B.n154 B.n149 585
R262 B.n364 B.n363 585
R263 B.n363 B.n362 585
R264 B.n365 B.n147 585
R265 B.n147 B.n146 585
R266 B.n367 B.n366 585
R267 B.n368 B.n367 585
R268 B.n3 B.n0 585
R269 B.n4 B.n3 585
R270 B.n466 B.n1 585
R271 B.n467 B.n466 585
R272 B.n465 B.n464 585
R273 B.n465 B.n8 585
R274 B.n463 B.n9 585
R275 B.n12 B.n9 585
R276 B.n462 B.n461 585
R277 B.n461 B.n460 585
R278 B.n11 B.n10 585
R279 B.n459 B.n11 585
R280 B.n457 B.n456 585
R281 B.n458 B.n457 585
R282 B.n455 B.n17 585
R283 B.n17 B.n16 585
R284 B.n454 B.n453 585
R285 B.n453 B.n452 585
R286 B.n19 B.n18 585
R287 B.n451 B.n19 585
R288 B.n449 B.n448 585
R289 B.n450 B.n449 585
R290 B.n447 B.n23 585
R291 B.n26 B.n23 585
R292 B.n446 B.n445 585
R293 B.n445 B.n444 585
R294 B.n25 B.n24 585
R295 B.n443 B.n25 585
R296 B.n441 B.n440 585
R297 B.n442 B.n441 585
R298 B.n439 B.n31 585
R299 B.n31 B.n30 585
R300 B.n438 B.n437 585
R301 B.n437 B.n436 585
R302 B.n33 B.n32 585
R303 B.n435 B.n33 585
R304 B.n433 B.n432 585
R305 B.n434 B.n433 585
R306 B.n431 B.n38 585
R307 B.n38 B.n37 585
R308 B.n430 B.n429 585
R309 B.n429 B.n428 585
R310 B.n40 B.n39 585
R311 B.n427 B.n40 585
R312 B.n425 B.n424 585
R313 B.n426 B.n425 585
R314 B.n423 B.n45 585
R315 B.n45 B.n44 585
R316 B.n422 B.n421 585
R317 B.n421 B.n420 585
R318 B.n47 B.n46 585
R319 B.n419 B.n47 585
R320 B.n417 B.n416 585
R321 B.n418 B.n417 585
R322 B.n415 B.n52 585
R323 B.n52 B.n51 585
R324 B.n470 B.n469 585
R325 B.n468 B.n2 585
R326 B.n413 B.n52 487.695
R327 B.n409 B.n72 487.695
R328 B.n213 B.n192 487.695
R329 B.n289 B.n194 487.695
R330 B.n411 B.n410 256.663
R331 B.n411 B.n70 256.663
R332 B.n411 B.n69 256.663
R333 B.n411 B.n68 256.663
R334 B.n411 B.n67 256.663
R335 B.n411 B.n66 256.663
R336 B.n411 B.n65 256.663
R337 B.n411 B.n64 256.663
R338 B.n411 B.n63 256.663
R339 B.n411 B.n62 256.663
R340 B.n411 B.n61 256.663
R341 B.n411 B.n60 256.663
R342 B.n411 B.n59 256.663
R343 B.n411 B.n58 256.663
R344 B.n411 B.n57 256.663
R345 B.n411 B.n56 256.663
R346 B.n411 B.n55 256.663
R347 B.n412 B.n411 256.663
R348 B.n288 B.n287 256.663
R349 B.n287 B.n197 256.663
R350 B.n287 B.n198 256.663
R351 B.n287 B.n199 256.663
R352 B.n287 B.n200 256.663
R353 B.n287 B.n201 256.663
R354 B.n287 B.n202 256.663
R355 B.n287 B.n203 256.663
R356 B.n287 B.n204 256.663
R357 B.n287 B.n205 256.663
R358 B.n287 B.n206 256.663
R359 B.n287 B.n207 256.663
R360 B.n287 B.n208 256.663
R361 B.n287 B.n209 256.663
R362 B.n287 B.n210 256.663
R363 B.n287 B.n211 256.663
R364 B.n287 B.n212 256.663
R365 B.n472 B.n471 256.663
R366 B.n75 B.t15 235.85
R367 B.n73 B.t4 235.85
R368 B.n218 B.t12 235.85
R369 B.n215 B.t8 235.85
R370 B.n287 B.n193 190.736
R371 B.n411 B.n51 190.736
R372 B.n77 B.n54 163.367
R373 B.n81 B.n80 163.367
R374 B.n85 B.n84 163.367
R375 B.n89 B.n88 163.367
R376 B.n93 B.n92 163.367
R377 B.n97 B.n96 163.367
R378 B.n102 B.n101 163.367
R379 B.n106 B.n105 163.367
R380 B.n110 B.n109 163.367
R381 B.n114 B.n113 163.367
R382 B.n118 B.n117 163.367
R383 B.n123 B.n122 163.367
R384 B.n127 B.n126 163.367
R385 B.n131 B.n130 163.367
R386 B.n135 B.n134 163.367
R387 B.n139 B.n138 163.367
R388 B.n141 B.n71 163.367
R389 B.n295 B.n192 163.367
R390 B.n295 B.n190 163.367
R391 B.n299 B.n190 163.367
R392 B.n299 B.n183 163.367
R393 B.n307 B.n183 163.367
R394 B.n307 B.n181 163.367
R395 B.n311 B.n181 163.367
R396 B.n311 B.n176 163.367
R397 B.n319 B.n176 163.367
R398 B.n319 B.n174 163.367
R399 B.n323 B.n174 163.367
R400 B.n323 B.n168 163.367
R401 B.n331 B.n168 163.367
R402 B.n331 B.n166 163.367
R403 B.n335 B.n166 163.367
R404 B.n335 B.n161 163.367
R405 B.n344 B.n161 163.367
R406 B.n344 B.n159 163.367
R407 B.n348 B.n159 163.367
R408 B.n348 B.n152 163.367
R409 B.n356 B.n152 163.367
R410 B.n356 B.n150 163.367
R411 B.n361 B.n150 163.367
R412 B.n361 B.n145 163.367
R413 B.n369 B.n145 163.367
R414 B.n370 B.n369 163.367
R415 B.n370 B.n5 163.367
R416 B.n6 B.n5 163.367
R417 B.n7 B.n6 163.367
R418 B.n376 B.n7 163.367
R419 B.n377 B.n376 163.367
R420 B.n377 B.n13 163.367
R421 B.n14 B.n13 163.367
R422 B.n15 B.n14 163.367
R423 B.n382 B.n15 163.367
R424 B.n382 B.n20 163.367
R425 B.n21 B.n20 163.367
R426 B.n22 B.n21 163.367
R427 B.n387 B.n22 163.367
R428 B.n387 B.n27 163.367
R429 B.n28 B.n27 163.367
R430 B.n29 B.n28 163.367
R431 B.n392 B.n29 163.367
R432 B.n392 B.n34 163.367
R433 B.n35 B.n34 163.367
R434 B.n36 B.n35 163.367
R435 B.n397 B.n36 163.367
R436 B.n397 B.n41 163.367
R437 B.n42 B.n41 163.367
R438 B.n43 B.n42 163.367
R439 B.n402 B.n43 163.367
R440 B.n402 B.n48 163.367
R441 B.n49 B.n48 163.367
R442 B.n50 B.n49 163.367
R443 B.n72 B.n50 163.367
R444 B.n286 B.n196 163.367
R445 B.n286 B.n214 163.367
R446 B.n282 B.n281 163.367
R447 B.n278 B.n277 163.367
R448 B.n274 B.n273 163.367
R449 B.n270 B.n269 163.367
R450 B.n266 B.n265 163.367
R451 B.n262 B.n261 163.367
R452 B.n258 B.n257 163.367
R453 B.n254 B.n253 163.367
R454 B.n250 B.n249 163.367
R455 B.n246 B.n245 163.367
R456 B.n242 B.n241 163.367
R457 B.n238 B.n237 163.367
R458 B.n234 B.n233 163.367
R459 B.n230 B.n229 163.367
R460 B.n226 B.n225 163.367
R461 B.n222 B.n213 163.367
R462 B.n293 B.n194 163.367
R463 B.n293 B.n188 163.367
R464 B.n301 B.n188 163.367
R465 B.n301 B.n186 163.367
R466 B.n305 B.n186 163.367
R467 B.n305 B.n180 163.367
R468 B.n313 B.n180 163.367
R469 B.n313 B.n178 163.367
R470 B.n317 B.n178 163.367
R471 B.n317 B.n172 163.367
R472 B.n325 B.n172 163.367
R473 B.n325 B.n170 163.367
R474 B.n329 B.n170 163.367
R475 B.n329 B.n164 163.367
R476 B.n338 B.n164 163.367
R477 B.n338 B.n162 163.367
R478 B.n342 B.n162 163.367
R479 B.n342 B.n157 163.367
R480 B.n350 B.n157 163.367
R481 B.n350 B.n155 163.367
R482 B.n354 B.n155 163.367
R483 B.n354 B.n149 163.367
R484 B.n363 B.n149 163.367
R485 B.n363 B.n147 163.367
R486 B.n367 B.n147 163.367
R487 B.n367 B.n3 163.367
R488 B.n470 B.n3 163.367
R489 B.n466 B.n2 163.367
R490 B.n466 B.n465 163.367
R491 B.n465 B.n9 163.367
R492 B.n461 B.n9 163.367
R493 B.n461 B.n11 163.367
R494 B.n457 B.n11 163.367
R495 B.n457 B.n17 163.367
R496 B.n453 B.n17 163.367
R497 B.n453 B.n19 163.367
R498 B.n449 B.n19 163.367
R499 B.n449 B.n23 163.367
R500 B.n445 B.n23 163.367
R501 B.n445 B.n25 163.367
R502 B.n441 B.n25 163.367
R503 B.n441 B.n31 163.367
R504 B.n437 B.n31 163.367
R505 B.n437 B.n33 163.367
R506 B.n433 B.n33 163.367
R507 B.n433 B.n38 163.367
R508 B.n429 B.n38 163.367
R509 B.n429 B.n40 163.367
R510 B.n425 B.n40 163.367
R511 B.n425 B.n45 163.367
R512 B.n421 B.n45 163.367
R513 B.n421 B.n47 163.367
R514 B.n417 B.n47 163.367
R515 B.n417 B.n52 163.367
R516 B.n73 B.t6 129.804
R517 B.n218 B.t14 129.804
R518 B.n75 B.t16 129.804
R519 B.n215 B.t11 129.804
R520 B.n294 B.n193 99.0078
R521 B.n294 B.n189 99.0078
R522 B.n300 B.n189 99.0078
R523 B.n300 B.n184 99.0078
R524 B.n306 B.n184 99.0078
R525 B.n306 B.n185 99.0078
R526 B.n312 B.n177 99.0078
R527 B.n318 B.n177 99.0078
R528 B.n318 B.n173 99.0078
R529 B.n324 B.n173 99.0078
R530 B.n324 B.n169 99.0078
R531 B.n330 B.n169 99.0078
R532 B.n330 B.n165 99.0078
R533 B.n337 B.n165 99.0078
R534 B.n337 B.n336 99.0078
R535 B.n343 B.n158 99.0078
R536 B.n349 B.n158 99.0078
R537 B.n349 B.n153 99.0078
R538 B.n355 B.n153 99.0078
R539 B.n355 B.n154 99.0078
R540 B.n362 B.n146 99.0078
R541 B.n368 B.n146 99.0078
R542 B.n368 B.n4 99.0078
R543 B.n469 B.n4 99.0078
R544 B.n469 B.n468 99.0078
R545 B.n468 B.n467 99.0078
R546 B.n467 B.n8 99.0078
R547 B.n12 B.n8 99.0078
R548 B.n460 B.n12 99.0078
R549 B.n459 B.n458 99.0078
R550 B.n458 B.n16 99.0078
R551 B.n452 B.n16 99.0078
R552 B.n452 B.n451 99.0078
R553 B.n451 B.n450 99.0078
R554 B.n444 B.n26 99.0078
R555 B.n444 B.n443 99.0078
R556 B.n443 B.n442 99.0078
R557 B.n442 B.n30 99.0078
R558 B.n436 B.n30 99.0078
R559 B.n436 B.n435 99.0078
R560 B.n435 B.n434 99.0078
R561 B.n434 B.n37 99.0078
R562 B.n428 B.n37 99.0078
R563 B.n427 B.n426 99.0078
R564 B.n426 B.n44 99.0078
R565 B.n420 B.n44 99.0078
R566 B.n420 B.n419 99.0078
R567 B.n419 B.n418 99.0078
R568 B.n418 B.n51 99.0078
R569 B.n74 B.t7 86.9435
R570 B.n219 B.t13 86.9435
R571 B.n76 B.t17 86.9432
R572 B.n216 B.t10 86.9432
R573 B.n343 B.t2 84.4479
R574 B.n450 B.t1 84.4479
R575 B.n413 B.n412 71.676
R576 B.n77 B.n55 71.676
R577 B.n81 B.n56 71.676
R578 B.n85 B.n57 71.676
R579 B.n89 B.n58 71.676
R580 B.n93 B.n59 71.676
R581 B.n97 B.n60 71.676
R582 B.n102 B.n61 71.676
R583 B.n106 B.n62 71.676
R584 B.n110 B.n63 71.676
R585 B.n114 B.n64 71.676
R586 B.n118 B.n65 71.676
R587 B.n123 B.n66 71.676
R588 B.n127 B.n67 71.676
R589 B.n131 B.n68 71.676
R590 B.n135 B.n69 71.676
R591 B.n139 B.n70 71.676
R592 B.n410 B.n71 71.676
R593 B.n410 B.n409 71.676
R594 B.n141 B.n70 71.676
R595 B.n138 B.n69 71.676
R596 B.n134 B.n68 71.676
R597 B.n130 B.n67 71.676
R598 B.n126 B.n66 71.676
R599 B.n122 B.n65 71.676
R600 B.n117 B.n64 71.676
R601 B.n113 B.n63 71.676
R602 B.n109 B.n62 71.676
R603 B.n105 B.n61 71.676
R604 B.n101 B.n60 71.676
R605 B.n96 B.n59 71.676
R606 B.n92 B.n58 71.676
R607 B.n88 B.n57 71.676
R608 B.n84 B.n56 71.676
R609 B.n80 B.n55 71.676
R610 B.n412 B.n54 71.676
R611 B.n289 B.n288 71.676
R612 B.n214 B.n197 71.676
R613 B.n281 B.n198 71.676
R614 B.n277 B.n199 71.676
R615 B.n273 B.n200 71.676
R616 B.n269 B.n201 71.676
R617 B.n265 B.n202 71.676
R618 B.n261 B.n203 71.676
R619 B.n257 B.n204 71.676
R620 B.n253 B.n205 71.676
R621 B.n249 B.n206 71.676
R622 B.n245 B.n207 71.676
R623 B.n241 B.n208 71.676
R624 B.n237 B.n209 71.676
R625 B.n233 B.n210 71.676
R626 B.n229 B.n211 71.676
R627 B.n225 B.n212 71.676
R628 B.n288 B.n196 71.676
R629 B.n282 B.n197 71.676
R630 B.n278 B.n198 71.676
R631 B.n274 B.n199 71.676
R632 B.n270 B.n200 71.676
R633 B.n266 B.n201 71.676
R634 B.n262 B.n202 71.676
R635 B.n258 B.n203 71.676
R636 B.n254 B.n204 71.676
R637 B.n250 B.n205 71.676
R638 B.n246 B.n206 71.676
R639 B.n242 B.n207 71.676
R640 B.n238 B.n208 71.676
R641 B.n234 B.n209 71.676
R642 B.n230 B.n210 71.676
R643 B.n226 B.n211 71.676
R644 B.n222 B.n212 71.676
R645 B.n471 B.n470 71.676
R646 B.n471 B.n2 71.676
R647 B.n154 B.t3 64.064
R648 B.t0 B.n459 64.064
R649 B.n99 B.n76 59.5399
R650 B.n120 B.n74 59.5399
R651 B.n220 B.n219 59.5399
R652 B.n217 B.n216 59.5399
R653 B.n312 B.t9 55.3281
R654 B.n428 B.t5 55.3281
R655 B.n185 B.t9 43.6802
R656 B.t5 B.n427 43.6802
R657 B.n76 B.n75 42.8611
R658 B.n74 B.n73 42.8611
R659 B.n219 B.n218 42.8611
R660 B.n216 B.n215 42.8611
R661 B.n362 B.t3 34.9442
R662 B.n460 B.t0 34.9442
R663 B.n291 B.n290 31.6883
R664 B.n221 B.n191 31.6883
R665 B.n408 B.n407 31.6883
R666 B.n415 B.n414 31.6883
R667 B B.n472 18.0485
R668 B.n336 B.t2 14.5604
R669 B.n26 B.t1 14.5604
R670 B.n292 B.n291 10.6151
R671 B.n292 B.n187 10.6151
R672 B.n302 B.n187 10.6151
R673 B.n303 B.n302 10.6151
R674 B.n304 B.n303 10.6151
R675 B.n304 B.n179 10.6151
R676 B.n314 B.n179 10.6151
R677 B.n315 B.n314 10.6151
R678 B.n316 B.n315 10.6151
R679 B.n316 B.n171 10.6151
R680 B.n326 B.n171 10.6151
R681 B.n327 B.n326 10.6151
R682 B.n328 B.n327 10.6151
R683 B.n328 B.n163 10.6151
R684 B.n339 B.n163 10.6151
R685 B.n340 B.n339 10.6151
R686 B.n341 B.n340 10.6151
R687 B.n341 B.n156 10.6151
R688 B.n351 B.n156 10.6151
R689 B.n352 B.n351 10.6151
R690 B.n353 B.n352 10.6151
R691 B.n353 B.n148 10.6151
R692 B.n364 B.n148 10.6151
R693 B.n365 B.n364 10.6151
R694 B.n366 B.n365 10.6151
R695 B.n366 B.n0 10.6151
R696 B.n290 B.n195 10.6151
R697 B.n285 B.n195 10.6151
R698 B.n285 B.n284 10.6151
R699 B.n284 B.n283 10.6151
R700 B.n283 B.n280 10.6151
R701 B.n280 B.n279 10.6151
R702 B.n279 B.n276 10.6151
R703 B.n276 B.n275 10.6151
R704 B.n275 B.n272 10.6151
R705 B.n272 B.n271 10.6151
R706 B.n271 B.n268 10.6151
R707 B.n268 B.n267 10.6151
R708 B.n264 B.n263 10.6151
R709 B.n263 B.n260 10.6151
R710 B.n260 B.n259 10.6151
R711 B.n259 B.n256 10.6151
R712 B.n256 B.n255 10.6151
R713 B.n255 B.n252 10.6151
R714 B.n252 B.n251 10.6151
R715 B.n251 B.n248 10.6151
R716 B.n248 B.n247 10.6151
R717 B.n244 B.n243 10.6151
R718 B.n243 B.n240 10.6151
R719 B.n240 B.n239 10.6151
R720 B.n239 B.n236 10.6151
R721 B.n236 B.n235 10.6151
R722 B.n235 B.n232 10.6151
R723 B.n232 B.n231 10.6151
R724 B.n231 B.n228 10.6151
R725 B.n228 B.n227 10.6151
R726 B.n227 B.n224 10.6151
R727 B.n224 B.n223 10.6151
R728 B.n223 B.n221 10.6151
R729 B.n296 B.n191 10.6151
R730 B.n297 B.n296 10.6151
R731 B.n298 B.n297 10.6151
R732 B.n298 B.n182 10.6151
R733 B.n308 B.n182 10.6151
R734 B.n309 B.n308 10.6151
R735 B.n310 B.n309 10.6151
R736 B.n310 B.n175 10.6151
R737 B.n320 B.n175 10.6151
R738 B.n321 B.n320 10.6151
R739 B.n322 B.n321 10.6151
R740 B.n322 B.n167 10.6151
R741 B.n332 B.n167 10.6151
R742 B.n333 B.n332 10.6151
R743 B.n334 B.n333 10.6151
R744 B.n334 B.n160 10.6151
R745 B.n345 B.n160 10.6151
R746 B.n346 B.n345 10.6151
R747 B.n347 B.n346 10.6151
R748 B.n347 B.n151 10.6151
R749 B.n357 B.n151 10.6151
R750 B.n358 B.n357 10.6151
R751 B.n360 B.n358 10.6151
R752 B.n360 B.n359 10.6151
R753 B.n359 B.n144 10.6151
R754 B.n371 B.n144 10.6151
R755 B.n372 B.n371 10.6151
R756 B.n373 B.n372 10.6151
R757 B.n374 B.n373 10.6151
R758 B.n375 B.n374 10.6151
R759 B.n378 B.n375 10.6151
R760 B.n379 B.n378 10.6151
R761 B.n380 B.n379 10.6151
R762 B.n381 B.n380 10.6151
R763 B.n383 B.n381 10.6151
R764 B.n384 B.n383 10.6151
R765 B.n385 B.n384 10.6151
R766 B.n386 B.n385 10.6151
R767 B.n388 B.n386 10.6151
R768 B.n389 B.n388 10.6151
R769 B.n390 B.n389 10.6151
R770 B.n391 B.n390 10.6151
R771 B.n393 B.n391 10.6151
R772 B.n394 B.n393 10.6151
R773 B.n395 B.n394 10.6151
R774 B.n396 B.n395 10.6151
R775 B.n398 B.n396 10.6151
R776 B.n399 B.n398 10.6151
R777 B.n400 B.n399 10.6151
R778 B.n401 B.n400 10.6151
R779 B.n403 B.n401 10.6151
R780 B.n404 B.n403 10.6151
R781 B.n405 B.n404 10.6151
R782 B.n406 B.n405 10.6151
R783 B.n407 B.n406 10.6151
R784 B.n464 B.n1 10.6151
R785 B.n464 B.n463 10.6151
R786 B.n463 B.n462 10.6151
R787 B.n462 B.n10 10.6151
R788 B.n456 B.n10 10.6151
R789 B.n456 B.n455 10.6151
R790 B.n455 B.n454 10.6151
R791 B.n454 B.n18 10.6151
R792 B.n448 B.n18 10.6151
R793 B.n448 B.n447 10.6151
R794 B.n447 B.n446 10.6151
R795 B.n446 B.n24 10.6151
R796 B.n440 B.n24 10.6151
R797 B.n440 B.n439 10.6151
R798 B.n439 B.n438 10.6151
R799 B.n438 B.n32 10.6151
R800 B.n432 B.n32 10.6151
R801 B.n432 B.n431 10.6151
R802 B.n431 B.n430 10.6151
R803 B.n430 B.n39 10.6151
R804 B.n424 B.n39 10.6151
R805 B.n424 B.n423 10.6151
R806 B.n423 B.n422 10.6151
R807 B.n422 B.n46 10.6151
R808 B.n416 B.n46 10.6151
R809 B.n416 B.n415 10.6151
R810 B.n414 B.n53 10.6151
R811 B.n78 B.n53 10.6151
R812 B.n79 B.n78 10.6151
R813 B.n82 B.n79 10.6151
R814 B.n83 B.n82 10.6151
R815 B.n86 B.n83 10.6151
R816 B.n87 B.n86 10.6151
R817 B.n90 B.n87 10.6151
R818 B.n91 B.n90 10.6151
R819 B.n94 B.n91 10.6151
R820 B.n95 B.n94 10.6151
R821 B.n98 B.n95 10.6151
R822 B.n103 B.n100 10.6151
R823 B.n104 B.n103 10.6151
R824 B.n107 B.n104 10.6151
R825 B.n108 B.n107 10.6151
R826 B.n111 B.n108 10.6151
R827 B.n112 B.n111 10.6151
R828 B.n115 B.n112 10.6151
R829 B.n116 B.n115 10.6151
R830 B.n119 B.n116 10.6151
R831 B.n124 B.n121 10.6151
R832 B.n125 B.n124 10.6151
R833 B.n128 B.n125 10.6151
R834 B.n129 B.n128 10.6151
R835 B.n132 B.n129 10.6151
R836 B.n133 B.n132 10.6151
R837 B.n136 B.n133 10.6151
R838 B.n137 B.n136 10.6151
R839 B.n140 B.n137 10.6151
R840 B.n142 B.n140 10.6151
R841 B.n143 B.n142 10.6151
R842 B.n408 B.n143 10.6151
R843 B.n267 B.n217 9.36635
R844 B.n244 B.n220 9.36635
R845 B.n99 B.n98 9.36635
R846 B.n121 B.n120 9.36635
R847 B.n472 B.n0 8.11757
R848 B.n472 B.n1 8.11757
R849 B.n264 B.n217 1.24928
R850 B.n247 B.n220 1.24928
R851 B.n100 B.n99 1.24928
R852 B.n120 B.n119 1.24928
R853 VP.n5 VP.n4 180.728
R854 VP.n14 VP.n13 180.728
R855 VP.n12 VP.n0 161.3
R856 VP.n11 VP.n10 161.3
R857 VP.n9 VP.n1 161.3
R858 VP.n8 VP.n7 161.3
R859 VP.n6 VP.n2 161.3
R860 VP.n3 VP.t0 67.0251
R861 VP.n3 VP.t1 66.586
R862 VP.n4 VP.n3 45.8095
R863 VP.n7 VP.n1 40.577
R864 VP.n11 VP.n1 40.577
R865 VP.n5 VP.t3 29.2282
R866 VP.n13 VP.t2 29.2282
R867 VP.n7 VP.n6 24.5923
R868 VP.n12 VP.n11 24.5923
R869 VP.n6 VP.n5 5.16479
R870 VP.n13 VP.n12 5.16479
R871 VP.n4 VP.n2 0.189894
R872 VP.n8 VP.n2 0.189894
R873 VP.n9 VP.n8 0.189894
R874 VP.n10 VP.n9 0.189894
R875 VP.n10 VP.n0 0.189894
R876 VP.n14 VP.n0 0.189894
R877 VP VP.n14 0.0516364
R878 VDD1 VDD1.n1 127.328
R879 VDD1 VDD1.n0 95.4652
R880 VDD1.n0 VDD1.t3 8.68471
R881 VDD1.n0 VDD1.t2 8.68471
R882 VDD1.n1 VDD1.t0 8.68471
R883 VDD1.n1 VDD1.t1 8.68471
C0 VP VTAIL 1.48297f
C1 VP VDD1 1.3018f
C2 VP VN 3.87271f
C3 VDD2 VTAIL 2.80547f
C4 VDD2 VDD1 0.851886f
C5 VDD2 VN 1.10228f
C6 VTAIL VDD1 2.75609f
C7 VP VDD2 0.354849f
C8 VN VTAIL 1.46886f
C9 VN VDD1 0.153995f
C10 VDD2 B 2.546196f
C11 VDD1 B 4.64559f
C12 VTAIL B 3.57173f
C13 VN B 7.817581f
C14 VP B 6.531845f
C15 VDD1.t3 B 0.035206f
C16 VDD1.t2 B 0.035206f
C17 VDD1.n0 B 0.24054f
C18 VDD1.t0 B 0.035206f
C19 VDD1.t1 B 0.035206f
C20 VDD1.n1 B 0.42865f
C21 VP.n0 B 0.023666f
C22 VP.t2 B 0.242724f
C23 VP.n1 B 0.019114f
C24 VP.n2 B 0.023666f
C25 VP.t3 B 0.242724f
C26 VP.t0 B 0.375651f
C27 VP.t1 B 0.374187f
C28 VP.n3 B 1.0042f
C29 VP.n4 B 0.988004f
C30 VP.n5 B 0.174352f
C31 VP.n6 B 0.02677f
C32 VP.n7 B 0.046788f
C33 VP.n8 B 0.023666f
C34 VP.n9 B 0.023666f
C35 VP.n10 B 0.023666f
C36 VP.n11 B 0.046788f
C37 VP.n12 B 0.02677f
C38 VP.n13 B 0.174352f
C39 VP.n14 B 0.025317f
C40 VTAIL.t7 B 0.232067f
C41 VTAIL.n0 B 0.222208f
C42 VTAIL.t3 B 0.232067f
C43 VTAIL.n1 B 0.268942f
C44 VTAIL.t2 B 0.232067f
C45 VTAIL.n2 B 0.666923f
C46 VTAIL.t4 B 0.232069f
C47 VTAIL.n3 B 0.666922f
C48 VTAIL.t5 B 0.232069f
C49 VTAIL.n4 B 0.268941f
C50 VTAIL.t0 B 0.232069f
C51 VTAIL.n5 B 0.268941f
C52 VTAIL.t1 B 0.232067f
C53 VTAIL.n6 B 0.666923f
C54 VTAIL.t6 B 0.232067f
C55 VTAIL.n7 B 0.614108f
C56 VDD2.t0 B 0.036137f
C57 VDD2.t1 B 0.036137f
C58 VDD2.n0 B 0.427461f
C59 VDD2.t2 B 0.036137f
C60 VDD2.t3 B 0.036137f
C61 VDD2.n1 B 0.246731f
C62 VDD2.n2 B 1.85381f
C63 VN.t0 B 0.372474f
C64 VN.t1 B 0.371022f
C65 VN.n0 B 0.254336f
C66 VN.t2 B 0.372474f
C67 VN.t3 B 0.371022f
C68 VN.n1 B 1.0097f
.ends

