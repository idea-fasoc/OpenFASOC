* NGSPICE file created from diff_pair_sample_1657.ext - technology: sky130A

.subckt diff_pair_sample_1657 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t5 w_n3146_n3140# sky130_fd_pr__pfet_01v8 ad=4.2354 pd=22.5 as=1.7919 ps=11.19 w=10.86 l=2.39
X1 B.t11 B.t9 B.t10 w_n3146_n3140# sky130_fd_pr__pfet_01v8 ad=4.2354 pd=22.5 as=0 ps=0 w=10.86 l=2.39
X2 VDD2.t5 VN.t0 VTAIL.t0 w_n3146_n3140# sky130_fd_pr__pfet_01v8 ad=4.2354 pd=22.5 as=1.7919 ps=11.19 w=10.86 l=2.39
X3 B.t8 B.t6 B.t7 w_n3146_n3140# sky130_fd_pr__pfet_01v8 ad=4.2354 pd=22.5 as=0 ps=0 w=10.86 l=2.39
X4 VTAIL.t10 VP.t1 VDD1.t4 w_n3146_n3140# sky130_fd_pr__pfet_01v8 ad=1.7919 pd=11.19 as=1.7919 ps=11.19 w=10.86 l=2.39
X5 VDD2.t4 VN.t1 VTAIL.t4 w_n3146_n3140# sky130_fd_pr__pfet_01v8 ad=4.2354 pd=22.5 as=1.7919 ps=11.19 w=10.86 l=2.39
X6 VTAIL.t11 VN.t2 VDD2.t3 w_n3146_n3140# sky130_fd_pr__pfet_01v8 ad=1.7919 pd=11.19 as=1.7919 ps=11.19 w=10.86 l=2.39
X7 VTAIL.t9 VP.t2 VDD1.t3 w_n3146_n3140# sky130_fd_pr__pfet_01v8 ad=1.7919 pd=11.19 as=1.7919 ps=11.19 w=10.86 l=2.39
X8 VDD2.t2 VN.t3 VTAIL.t2 w_n3146_n3140# sky130_fd_pr__pfet_01v8 ad=1.7919 pd=11.19 as=4.2354 ps=22.5 w=10.86 l=2.39
X9 VDD1.t2 VP.t3 VTAIL.t8 w_n3146_n3140# sky130_fd_pr__pfet_01v8 ad=1.7919 pd=11.19 as=4.2354 ps=22.5 w=10.86 l=2.39
X10 VDD1.t1 VP.t4 VTAIL.t7 w_n3146_n3140# sky130_fd_pr__pfet_01v8 ad=4.2354 pd=22.5 as=1.7919 ps=11.19 w=10.86 l=2.39
X11 VTAIL.t1 VN.t4 VDD2.t1 w_n3146_n3140# sky130_fd_pr__pfet_01v8 ad=1.7919 pd=11.19 as=1.7919 ps=11.19 w=10.86 l=2.39
X12 B.t5 B.t3 B.t4 w_n3146_n3140# sky130_fd_pr__pfet_01v8 ad=4.2354 pd=22.5 as=0 ps=0 w=10.86 l=2.39
X13 B.t2 B.t0 B.t1 w_n3146_n3140# sky130_fd_pr__pfet_01v8 ad=4.2354 pd=22.5 as=0 ps=0 w=10.86 l=2.39
X14 VDD2.t0 VN.t5 VTAIL.t3 w_n3146_n3140# sky130_fd_pr__pfet_01v8 ad=1.7919 pd=11.19 as=4.2354 ps=22.5 w=10.86 l=2.39
X15 VDD1.t0 VP.t5 VTAIL.t6 w_n3146_n3140# sky130_fd_pr__pfet_01v8 ad=1.7919 pd=11.19 as=4.2354 ps=22.5 w=10.86 l=2.39
R0 VP.n11 VP.n8 161.3
R1 VP.n13 VP.n12 161.3
R2 VP.n14 VP.n7 161.3
R3 VP.n16 VP.n15 161.3
R4 VP.n17 VP.n6 161.3
R5 VP.n37 VP.n0 161.3
R6 VP.n36 VP.n35 161.3
R7 VP.n34 VP.n1 161.3
R8 VP.n33 VP.n32 161.3
R9 VP.n31 VP.n2 161.3
R10 VP.n30 VP.n29 161.3
R11 VP.n28 VP.n3 161.3
R12 VP.n27 VP.n26 161.3
R13 VP.n25 VP.n4 161.3
R14 VP.n24 VP.n23 161.3
R15 VP.n22 VP.n5 161.3
R16 VP.n9 VP.t0 143.528
R17 VP.n30 VP.t2 109.51
R18 VP.n20 VP.t4 109.51
R19 VP.n38 VP.t5 109.51
R20 VP.n10 VP.t1 109.51
R21 VP.n18 VP.t3 109.51
R22 VP.n21 VP.n20 100.088
R23 VP.n39 VP.n38 100.088
R24 VP.n19 VP.n18 100.088
R25 VP.n26 VP.n25 54.1398
R26 VP.n32 VP.n1 54.1398
R27 VP.n12 VP.n7 54.1398
R28 VP.n10 VP.n9 48.0647
R29 VP.n21 VP.n19 46.9694
R30 VP.n25 VP.n24 27.0143
R31 VP.n36 VP.n1 27.0143
R32 VP.n16 VP.n7 27.0143
R33 VP.n24 VP.n5 24.5923
R34 VP.n26 VP.n3 24.5923
R35 VP.n30 VP.n3 24.5923
R36 VP.n31 VP.n30 24.5923
R37 VP.n32 VP.n31 24.5923
R38 VP.n37 VP.n36 24.5923
R39 VP.n17 VP.n16 24.5923
R40 VP.n11 VP.n10 24.5923
R41 VP.n12 VP.n11 24.5923
R42 VP.n20 VP.n5 10.8209
R43 VP.n38 VP.n37 10.8209
R44 VP.n18 VP.n17 10.8209
R45 VP.n9 VP.n8 6.7696
R46 VP.n19 VP.n6 0.278335
R47 VP.n22 VP.n21 0.278335
R48 VP.n39 VP.n0 0.278335
R49 VP.n13 VP.n8 0.189894
R50 VP.n14 VP.n13 0.189894
R51 VP.n15 VP.n14 0.189894
R52 VP.n15 VP.n6 0.189894
R53 VP.n23 VP.n22 0.189894
R54 VP.n23 VP.n4 0.189894
R55 VP.n27 VP.n4 0.189894
R56 VP.n28 VP.n27 0.189894
R57 VP.n29 VP.n28 0.189894
R58 VP.n29 VP.n2 0.189894
R59 VP.n33 VP.n2 0.189894
R60 VP.n34 VP.n33 0.189894
R61 VP.n35 VP.n34 0.189894
R62 VP.n35 VP.n0 0.189894
R63 VP VP.n39 0.153485
R64 VTAIL.n234 VTAIL.n182 756.745
R65 VTAIL.n54 VTAIL.n2 756.745
R66 VTAIL.n176 VTAIL.n124 756.745
R67 VTAIL.n116 VTAIL.n64 756.745
R68 VTAIL.n201 VTAIL.n200 585
R69 VTAIL.n198 VTAIL.n197 585
R70 VTAIL.n207 VTAIL.n206 585
R71 VTAIL.n209 VTAIL.n208 585
R72 VTAIL.n194 VTAIL.n193 585
R73 VTAIL.n215 VTAIL.n214 585
R74 VTAIL.n218 VTAIL.n217 585
R75 VTAIL.n216 VTAIL.n190 585
R76 VTAIL.n223 VTAIL.n189 585
R77 VTAIL.n225 VTAIL.n224 585
R78 VTAIL.n227 VTAIL.n226 585
R79 VTAIL.n186 VTAIL.n185 585
R80 VTAIL.n233 VTAIL.n232 585
R81 VTAIL.n235 VTAIL.n234 585
R82 VTAIL.n21 VTAIL.n20 585
R83 VTAIL.n18 VTAIL.n17 585
R84 VTAIL.n27 VTAIL.n26 585
R85 VTAIL.n29 VTAIL.n28 585
R86 VTAIL.n14 VTAIL.n13 585
R87 VTAIL.n35 VTAIL.n34 585
R88 VTAIL.n38 VTAIL.n37 585
R89 VTAIL.n36 VTAIL.n10 585
R90 VTAIL.n43 VTAIL.n9 585
R91 VTAIL.n45 VTAIL.n44 585
R92 VTAIL.n47 VTAIL.n46 585
R93 VTAIL.n6 VTAIL.n5 585
R94 VTAIL.n53 VTAIL.n52 585
R95 VTAIL.n55 VTAIL.n54 585
R96 VTAIL.n177 VTAIL.n176 585
R97 VTAIL.n175 VTAIL.n174 585
R98 VTAIL.n128 VTAIL.n127 585
R99 VTAIL.n169 VTAIL.n168 585
R100 VTAIL.n167 VTAIL.n166 585
R101 VTAIL.n165 VTAIL.n131 585
R102 VTAIL.n135 VTAIL.n132 585
R103 VTAIL.n160 VTAIL.n159 585
R104 VTAIL.n158 VTAIL.n157 585
R105 VTAIL.n137 VTAIL.n136 585
R106 VTAIL.n152 VTAIL.n151 585
R107 VTAIL.n150 VTAIL.n149 585
R108 VTAIL.n141 VTAIL.n140 585
R109 VTAIL.n144 VTAIL.n143 585
R110 VTAIL.n117 VTAIL.n116 585
R111 VTAIL.n115 VTAIL.n114 585
R112 VTAIL.n68 VTAIL.n67 585
R113 VTAIL.n109 VTAIL.n108 585
R114 VTAIL.n107 VTAIL.n106 585
R115 VTAIL.n105 VTAIL.n71 585
R116 VTAIL.n75 VTAIL.n72 585
R117 VTAIL.n100 VTAIL.n99 585
R118 VTAIL.n98 VTAIL.n97 585
R119 VTAIL.n77 VTAIL.n76 585
R120 VTAIL.n92 VTAIL.n91 585
R121 VTAIL.n90 VTAIL.n89 585
R122 VTAIL.n81 VTAIL.n80 585
R123 VTAIL.n84 VTAIL.n83 585
R124 VTAIL.t8 VTAIL.n142 329.038
R125 VTAIL.t2 VTAIL.n82 329.038
R126 VTAIL.t3 VTAIL.n199 329.038
R127 VTAIL.t6 VTAIL.n19 329.038
R128 VTAIL.n200 VTAIL.n197 171.744
R129 VTAIL.n207 VTAIL.n197 171.744
R130 VTAIL.n208 VTAIL.n207 171.744
R131 VTAIL.n208 VTAIL.n193 171.744
R132 VTAIL.n215 VTAIL.n193 171.744
R133 VTAIL.n217 VTAIL.n215 171.744
R134 VTAIL.n217 VTAIL.n216 171.744
R135 VTAIL.n216 VTAIL.n189 171.744
R136 VTAIL.n225 VTAIL.n189 171.744
R137 VTAIL.n226 VTAIL.n225 171.744
R138 VTAIL.n226 VTAIL.n185 171.744
R139 VTAIL.n233 VTAIL.n185 171.744
R140 VTAIL.n234 VTAIL.n233 171.744
R141 VTAIL.n20 VTAIL.n17 171.744
R142 VTAIL.n27 VTAIL.n17 171.744
R143 VTAIL.n28 VTAIL.n27 171.744
R144 VTAIL.n28 VTAIL.n13 171.744
R145 VTAIL.n35 VTAIL.n13 171.744
R146 VTAIL.n37 VTAIL.n35 171.744
R147 VTAIL.n37 VTAIL.n36 171.744
R148 VTAIL.n36 VTAIL.n9 171.744
R149 VTAIL.n45 VTAIL.n9 171.744
R150 VTAIL.n46 VTAIL.n45 171.744
R151 VTAIL.n46 VTAIL.n5 171.744
R152 VTAIL.n53 VTAIL.n5 171.744
R153 VTAIL.n54 VTAIL.n53 171.744
R154 VTAIL.n176 VTAIL.n175 171.744
R155 VTAIL.n175 VTAIL.n127 171.744
R156 VTAIL.n168 VTAIL.n127 171.744
R157 VTAIL.n168 VTAIL.n167 171.744
R158 VTAIL.n167 VTAIL.n131 171.744
R159 VTAIL.n135 VTAIL.n131 171.744
R160 VTAIL.n159 VTAIL.n135 171.744
R161 VTAIL.n159 VTAIL.n158 171.744
R162 VTAIL.n158 VTAIL.n136 171.744
R163 VTAIL.n151 VTAIL.n136 171.744
R164 VTAIL.n151 VTAIL.n150 171.744
R165 VTAIL.n150 VTAIL.n140 171.744
R166 VTAIL.n143 VTAIL.n140 171.744
R167 VTAIL.n116 VTAIL.n115 171.744
R168 VTAIL.n115 VTAIL.n67 171.744
R169 VTAIL.n108 VTAIL.n67 171.744
R170 VTAIL.n108 VTAIL.n107 171.744
R171 VTAIL.n107 VTAIL.n71 171.744
R172 VTAIL.n75 VTAIL.n71 171.744
R173 VTAIL.n99 VTAIL.n75 171.744
R174 VTAIL.n99 VTAIL.n98 171.744
R175 VTAIL.n98 VTAIL.n76 171.744
R176 VTAIL.n91 VTAIL.n76 171.744
R177 VTAIL.n91 VTAIL.n90 171.744
R178 VTAIL.n90 VTAIL.n80 171.744
R179 VTAIL.n83 VTAIL.n80 171.744
R180 VTAIL.n200 VTAIL.t3 85.8723
R181 VTAIL.n20 VTAIL.t6 85.8723
R182 VTAIL.n143 VTAIL.t8 85.8723
R183 VTAIL.n83 VTAIL.t2 85.8723
R184 VTAIL.n123 VTAIL.n122 62.6783
R185 VTAIL.n63 VTAIL.n62 62.6783
R186 VTAIL.n1 VTAIL.n0 62.6781
R187 VTAIL.n61 VTAIL.n60 62.6781
R188 VTAIL.n239 VTAIL.n238 35.6763
R189 VTAIL.n59 VTAIL.n58 35.6763
R190 VTAIL.n181 VTAIL.n180 35.6763
R191 VTAIL.n121 VTAIL.n120 35.6763
R192 VTAIL.n63 VTAIL.n61 26.4186
R193 VTAIL.n239 VTAIL.n181 24.0738
R194 VTAIL.n224 VTAIL.n223 13.1884
R195 VTAIL.n44 VTAIL.n43 13.1884
R196 VTAIL.n166 VTAIL.n165 13.1884
R197 VTAIL.n106 VTAIL.n105 13.1884
R198 VTAIL.n222 VTAIL.n190 12.8005
R199 VTAIL.n227 VTAIL.n188 12.8005
R200 VTAIL.n42 VTAIL.n10 12.8005
R201 VTAIL.n47 VTAIL.n8 12.8005
R202 VTAIL.n169 VTAIL.n130 12.8005
R203 VTAIL.n164 VTAIL.n132 12.8005
R204 VTAIL.n109 VTAIL.n70 12.8005
R205 VTAIL.n104 VTAIL.n72 12.8005
R206 VTAIL.n219 VTAIL.n218 12.0247
R207 VTAIL.n228 VTAIL.n186 12.0247
R208 VTAIL.n39 VTAIL.n38 12.0247
R209 VTAIL.n48 VTAIL.n6 12.0247
R210 VTAIL.n170 VTAIL.n128 12.0247
R211 VTAIL.n161 VTAIL.n160 12.0247
R212 VTAIL.n110 VTAIL.n68 12.0247
R213 VTAIL.n101 VTAIL.n100 12.0247
R214 VTAIL.n214 VTAIL.n192 11.249
R215 VTAIL.n232 VTAIL.n231 11.249
R216 VTAIL.n34 VTAIL.n12 11.249
R217 VTAIL.n52 VTAIL.n51 11.249
R218 VTAIL.n174 VTAIL.n173 11.249
R219 VTAIL.n157 VTAIL.n134 11.249
R220 VTAIL.n114 VTAIL.n113 11.249
R221 VTAIL.n97 VTAIL.n74 11.249
R222 VTAIL.n201 VTAIL.n199 10.7239
R223 VTAIL.n21 VTAIL.n19 10.7239
R224 VTAIL.n144 VTAIL.n142 10.7239
R225 VTAIL.n84 VTAIL.n82 10.7239
R226 VTAIL.n213 VTAIL.n194 10.4732
R227 VTAIL.n235 VTAIL.n184 10.4732
R228 VTAIL.n33 VTAIL.n14 10.4732
R229 VTAIL.n55 VTAIL.n4 10.4732
R230 VTAIL.n177 VTAIL.n126 10.4732
R231 VTAIL.n156 VTAIL.n137 10.4732
R232 VTAIL.n117 VTAIL.n66 10.4732
R233 VTAIL.n96 VTAIL.n77 10.4732
R234 VTAIL.n210 VTAIL.n209 9.69747
R235 VTAIL.n236 VTAIL.n182 9.69747
R236 VTAIL.n30 VTAIL.n29 9.69747
R237 VTAIL.n56 VTAIL.n2 9.69747
R238 VTAIL.n178 VTAIL.n124 9.69747
R239 VTAIL.n153 VTAIL.n152 9.69747
R240 VTAIL.n118 VTAIL.n64 9.69747
R241 VTAIL.n93 VTAIL.n92 9.69747
R242 VTAIL.n238 VTAIL.n237 9.45567
R243 VTAIL.n58 VTAIL.n57 9.45567
R244 VTAIL.n180 VTAIL.n179 9.45567
R245 VTAIL.n120 VTAIL.n119 9.45567
R246 VTAIL.n237 VTAIL.n236 9.3005
R247 VTAIL.n184 VTAIL.n183 9.3005
R248 VTAIL.n231 VTAIL.n230 9.3005
R249 VTAIL.n229 VTAIL.n228 9.3005
R250 VTAIL.n188 VTAIL.n187 9.3005
R251 VTAIL.n203 VTAIL.n202 9.3005
R252 VTAIL.n205 VTAIL.n204 9.3005
R253 VTAIL.n196 VTAIL.n195 9.3005
R254 VTAIL.n211 VTAIL.n210 9.3005
R255 VTAIL.n213 VTAIL.n212 9.3005
R256 VTAIL.n192 VTAIL.n191 9.3005
R257 VTAIL.n220 VTAIL.n219 9.3005
R258 VTAIL.n222 VTAIL.n221 9.3005
R259 VTAIL.n57 VTAIL.n56 9.3005
R260 VTAIL.n4 VTAIL.n3 9.3005
R261 VTAIL.n51 VTAIL.n50 9.3005
R262 VTAIL.n49 VTAIL.n48 9.3005
R263 VTAIL.n8 VTAIL.n7 9.3005
R264 VTAIL.n23 VTAIL.n22 9.3005
R265 VTAIL.n25 VTAIL.n24 9.3005
R266 VTAIL.n16 VTAIL.n15 9.3005
R267 VTAIL.n31 VTAIL.n30 9.3005
R268 VTAIL.n33 VTAIL.n32 9.3005
R269 VTAIL.n12 VTAIL.n11 9.3005
R270 VTAIL.n40 VTAIL.n39 9.3005
R271 VTAIL.n42 VTAIL.n41 9.3005
R272 VTAIL.n146 VTAIL.n145 9.3005
R273 VTAIL.n148 VTAIL.n147 9.3005
R274 VTAIL.n139 VTAIL.n138 9.3005
R275 VTAIL.n154 VTAIL.n153 9.3005
R276 VTAIL.n156 VTAIL.n155 9.3005
R277 VTAIL.n134 VTAIL.n133 9.3005
R278 VTAIL.n162 VTAIL.n161 9.3005
R279 VTAIL.n164 VTAIL.n163 9.3005
R280 VTAIL.n179 VTAIL.n178 9.3005
R281 VTAIL.n126 VTAIL.n125 9.3005
R282 VTAIL.n173 VTAIL.n172 9.3005
R283 VTAIL.n171 VTAIL.n170 9.3005
R284 VTAIL.n130 VTAIL.n129 9.3005
R285 VTAIL.n86 VTAIL.n85 9.3005
R286 VTAIL.n88 VTAIL.n87 9.3005
R287 VTAIL.n79 VTAIL.n78 9.3005
R288 VTAIL.n94 VTAIL.n93 9.3005
R289 VTAIL.n96 VTAIL.n95 9.3005
R290 VTAIL.n74 VTAIL.n73 9.3005
R291 VTAIL.n102 VTAIL.n101 9.3005
R292 VTAIL.n104 VTAIL.n103 9.3005
R293 VTAIL.n119 VTAIL.n118 9.3005
R294 VTAIL.n66 VTAIL.n65 9.3005
R295 VTAIL.n113 VTAIL.n112 9.3005
R296 VTAIL.n111 VTAIL.n110 9.3005
R297 VTAIL.n70 VTAIL.n69 9.3005
R298 VTAIL.n206 VTAIL.n196 8.92171
R299 VTAIL.n26 VTAIL.n16 8.92171
R300 VTAIL.n149 VTAIL.n139 8.92171
R301 VTAIL.n89 VTAIL.n79 8.92171
R302 VTAIL.n205 VTAIL.n198 8.14595
R303 VTAIL.n25 VTAIL.n18 8.14595
R304 VTAIL.n148 VTAIL.n141 8.14595
R305 VTAIL.n88 VTAIL.n81 8.14595
R306 VTAIL.n202 VTAIL.n201 7.3702
R307 VTAIL.n22 VTAIL.n21 7.3702
R308 VTAIL.n145 VTAIL.n144 7.3702
R309 VTAIL.n85 VTAIL.n84 7.3702
R310 VTAIL.n202 VTAIL.n198 5.81868
R311 VTAIL.n22 VTAIL.n18 5.81868
R312 VTAIL.n145 VTAIL.n141 5.81868
R313 VTAIL.n85 VTAIL.n81 5.81868
R314 VTAIL.n206 VTAIL.n205 5.04292
R315 VTAIL.n26 VTAIL.n25 5.04292
R316 VTAIL.n149 VTAIL.n148 5.04292
R317 VTAIL.n89 VTAIL.n88 5.04292
R318 VTAIL.n209 VTAIL.n196 4.26717
R319 VTAIL.n238 VTAIL.n182 4.26717
R320 VTAIL.n29 VTAIL.n16 4.26717
R321 VTAIL.n58 VTAIL.n2 4.26717
R322 VTAIL.n180 VTAIL.n124 4.26717
R323 VTAIL.n152 VTAIL.n139 4.26717
R324 VTAIL.n120 VTAIL.n64 4.26717
R325 VTAIL.n92 VTAIL.n79 4.26717
R326 VTAIL.n210 VTAIL.n194 3.49141
R327 VTAIL.n236 VTAIL.n235 3.49141
R328 VTAIL.n30 VTAIL.n14 3.49141
R329 VTAIL.n56 VTAIL.n55 3.49141
R330 VTAIL.n178 VTAIL.n177 3.49141
R331 VTAIL.n153 VTAIL.n137 3.49141
R332 VTAIL.n118 VTAIL.n117 3.49141
R333 VTAIL.n93 VTAIL.n77 3.49141
R334 VTAIL.n0 VTAIL.t0 2.99359
R335 VTAIL.n0 VTAIL.t11 2.99359
R336 VTAIL.n60 VTAIL.t7 2.99359
R337 VTAIL.n60 VTAIL.t9 2.99359
R338 VTAIL.n122 VTAIL.t5 2.99359
R339 VTAIL.n122 VTAIL.t10 2.99359
R340 VTAIL.n62 VTAIL.t4 2.99359
R341 VTAIL.n62 VTAIL.t1 2.99359
R342 VTAIL.n214 VTAIL.n213 2.71565
R343 VTAIL.n232 VTAIL.n184 2.71565
R344 VTAIL.n34 VTAIL.n33 2.71565
R345 VTAIL.n52 VTAIL.n4 2.71565
R346 VTAIL.n174 VTAIL.n126 2.71565
R347 VTAIL.n157 VTAIL.n156 2.71565
R348 VTAIL.n114 VTAIL.n66 2.71565
R349 VTAIL.n97 VTAIL.n96 2.71565
R350 VTAIL.n203 VTAIL.n199 2.41282
R351 VTAIL.n23 VTAIL.n19 2.41282
R352 VTAIL.n146 VTAIL.n142 2.41282
R353 VTAIL.n86 VTAIL.n82 2.41282
R354 VTAIL.n121 VTAIL.n63 2.34533
R355 VTAIL.n181 VTAIL.n123 2.34533
R356 VTAIL.n61 VTAIL.n59 2.34533
R357 VTAIL.n218 VTAIL.n192 1.93989
R358 VTAIL.n231 VTAIL.n186 1.93989
R359 VTAIL.n38 VTAIL.n12 1.93989
R360 VTAIL.n51 VTAIL.n6 1.93989
R361 VTAIL.n173 VTAIL.n128 1.93989
R362 VTAIL.n160 VTAIL.n134 1.93989
R363 VTAIL.n113 VTAIL.n68 1.93989
R364 VTAIL.n100 VTAIL.n74 1.93989
R365 VTAIL VTAIL.n239 1.70093
R366 VTAIL.n123 VTAIL.n121 1.64274
R367 VTAIL.n59 VTAIL.n1 1.64274
R368 VTAIL.n219 VTAIL.n190 1.16414
R369 VTAIL.n228 VTAIL.n227 1.16414
R370 VTAIL.n39 VTAIL.n10 1.16414
R371 VTAIL.n48 VTAIL.n47 1.16414
R372 VTAIL.n170 VTAIL.n169 1.16414
R373 VTAIL.n161 VTAIL.n132 1.16414
R374 VTAIL.n110 VTAIL.n109 1.16414
R375 VTAIL.n101 VTAIL.n72 1.16414
R376 VTAIL VTAIL.n1 0.644897
R377 VTAIL.n223 VTAIL.n222 0.388379
R378 VTAIL.n224 VTAIL.n188 0.388379
R379 VTAIL.n43 VTAIL.n42 0.388379
R380 VTAIL.n44 VTAIL.n8 0.388379
R381 VTAIL.n166 VTAIL.n130 0.388379
R382 VTAIL.n165 VTAIL.n164 0.388379
R383 VTAIL.n106 VTAIL.n70 0.388379
R384 VTAIL.n105 VTAIL.n104 0.388379
R385 VTAIL.n204 VTAIL.n203 0.155672
R386 VTAIL.n204 VTAIL.n195 0.155672
R387 VTAIL.n211 VTAIL.n195 0.155672
R388 VTAIL.n212 VTAIL.n211 0.155672
R389 VTAIL.n212 VTAIL.n191 0.155672
R390 VTAIL.n220 VTAIL.n191 0.155672
R391 VTAIL.n221 VTAIL.n220 0.155672
R392 VTAIL.n221 VTAIL.n187 0.155672
R393 VTAIL.n229 VTAIL.n187 0.155672
R394 VTAIL.n230 VTAIL.n229 0.155672
R395 VTAIL.n230 VTAIL.n183 0.155672
R396 VTAIL.n237 VTAIL.n183 0.155672
R397 VTAIL.n24 VTAIL.n23 0.155672
R398 VTAIL.n24 VTAIL.n15 0.155672
R399 VTAIL.n31 VTAIL.n15 0.155672
R400 VTAIL.n32 VTAIL.n31 0.155672
R401 VTAIL.n32 VTAIL.n11 0.155672
R402 VTAIL.n40 VTAIL.n11 0.155672
R403 VTAIL.n41 VTAIL.n40 0.155672
R404 VTAIL.n41 VTAIL.n7 0.155672
R405 VTAIL.n49 VTAIL.n7 0.155672
R406 VTAIL.n50 VTAIL.n49 0.155672
R407 VTAIL.n50 VTAIL.n3 0.155672
R408 VTAIL.n57 VTAIL.n3 0.155672
R409 VTAIL.n179 VTAIL.n125 0.155672
R410 VTAIL.n172 VTAIL.n125 0.155672
R411 VTAIL.n172 VTAIL.n171 0.155672
R412 VTAIL.n171 VTAIL.n129 0.155672
R413 VTAIL.n163 VTAIL.n129 0.155672
R414 VTAIL.n163 VTAIL.n162 0.155672
R415 VTAIL.n162 VTAIL.n133 0.155672
R416 VTAIL.n155 VTAIL.n133 0.155672
R417 VTAIL.n155 VTAIL.n154 0.155672
R418 VTAIL.n154 VTAIL.n138 0.155672
R419 VTAIL.n147 VTAIL.n138 0.155672
R420 VTAIL.n147 VTAIL.n146 0.155672
R421 VTAIL.n119 VTAIL.n65 0.155672
R422 VTAIL.n112 VTAIL.n65 0.155672
R423 VTAIL.n112 VTAIL.n111 0.155672
R424 VTAIL.n111 VTAIL.n69 0.155672
R425 VTAIL.n103 VTAIL.n69 0.155672
R426 VTAIL.n103 VTAIL.n102 0.155672
R427 VTAIL.n102 VTAIL.n73 0.155672
R428 VTAIL.n95 VTAIL.n73 0.155672
R429 VTAIL.n95 VTAIL.n94 0.155672
R430 VTAIL.n94 VTAIL.n78 0.155672
R431 VTAIL.n87 VTAIL.n78 0.155672
R432 VTAIL.n87 VTAIL.n86 0.155672
R433 VDD1.n52 VDD1.n0 756.745
R434 VDD1.n109 VDD1.n57 756.745
R435 VDD1.n53 VDD1.n52 585
R436 VDD1.n51 VDD1.n50 585
R437 VDD1.n4 VDD1.n3 585
R438 VDD1.n45 VDD1.n44 585
R439 VDD1.n43 VDD1.n42 585
R440 VDD1.n41 VDD1.n7 585
R441 VDD1.n11 VDD1.n8 585
R442 VDD1.n36 VDD1.n35 585
R443 VDD1.n34 VDD1.n33 585
R444 VDD1.n13 VDD1.n12 585
R445 VDD1.n28 VDD1.n27 585
R446 VDD1.n26 VDD1.n25 585
R447 VDD1.n17 VDD1.n16 585
R448 VDD1.n20 VDD1.n19 585
R449 VDD1.n76 VDD1.n75 585
R450 VDD1.n73 VDD1.n72 585
R451 VDD1.n82 VDD1.n81 585
R452 VDD1.n84 VDD1.n83 585
R453 VDD1.n69 VDD1.n68 585
R454 VDD1.n90 VDD1.n89 585
R455 VDD1.n93 VDD1.n92 585
R456 VDD1.n91 VDD1.n65 585
R457 VDD1.n98 VDD1.n64 585
R458 VDD1.n100 VDD1.n99 585
R459 VDD1.n102 VDD1.n101 585
R460 VDD1.n61 VDD1.n60 585
R461 VDD1.n108 VDD1.n107 585
R462 VDD1.n110 VDD1.n109 585
R463 VDD1.t5 VDD1.n18 329.038
R464 VDD1.t1 VDD1.n74 329.038
R465 VDD1.n52 VDD1.n51 171.744
R466 VDD1.n51 VDD1.n3 171.744
R467 VDD1.n44 VDD1.n3 171.744
R468 VDD1.n44 VDD1.n43 171.744
R469 VDD1.n43 VDD1.n7 171.744
R470 VDD1.n11 VDD1.n7 171.744
R471 VDD1.n35 VDD1.n11 171.744
R472 VDD1.n35 VDD1.n34 171.744
R473 VDD1.n34 VDD1.n12 171.744
R474 VDD1.n27 VDD1.n12 171.744
R475 VDD1.n27 VDD1.n26 171.744
R476 VDD1.n26 VDD1.n16 171.744
R477 VDD1.n19 VDD1.n16 171.744
R478 VDD1.n75 VDD1.n72 171.744
R479 VDD1.n82 VDD1.n72 171.744
R480 VDD1.n83 VDD1.n82 171.744
R481 VDD1.n83 VDD1.n68 171.744
R482 VDD1.n90 VDD1.n68 171.744
R483 VDD1.n92 VDD1.n90 171.744
R484 VDD1.n92 VDD1.n91 171.744
R485 VDD1.n91 VDD1.n64 171.744
R486 VDD1.n100 VDD1.n64 171.744
R487 VDD1.n101 VDD1.n100 171.744
R488 VDD1.n101 VDD1.n60 171.744
R489 VDD1.n108 VDD1.n60 171.744
R490 VDD1.n109 VDD1.n108 171.744
R491 VDD1.n19 VDD1.t5 85.8723
R492 VDD1.n75 VDD1.t1 85.8723
R493 VDD1.n115 VDD1.n114 79.8878
R494 VDD1.n117 VDD1.n116 79.3569
R495 VDD1 VDD1.n56 54.1719
R496 VDD1.n115 VDD1.n113 54.0583
R497 VDD1.n117 VDD1.n115 42.4535
R498 VDD1.n42 VDD1.n41 13.1884
R499 VDD1.n99 VDD1.n98 13.1884
R500 VDD1.n45 VDD1.n6 12.8005
R501 VDD1.n40 VDD1.n8 12.8005
R502 VDD1.n97 VDD1.n65 12.8005
R503 VDD1.n102 VDD1.n63 12.8005
R504 VDD1.n46 VDD1.n4 12.0247
R505 VDD1.n37 VDD1.n36 12.0247
R506 VDD1.n94 VDD1.n93 12.0247
R507 VDD1.n103 VDD1.n61 12.0247
R508 VDD1.n50 VDD1.n49 11.249
R509 VDD1.n33 VDD1.n10 11.249
R510 VDD1.n89 VDD1.n67 11.249
R511 VDD1.n107 VDD1.n106 11.249
R512 VDD1.n20 VDD1.n18 10.7239
R513 VDD1.n76 VDD1.n74 10.7239
R514 VDD1.n53 VDD1.n2 10.4732
R515 VDD1.n32 VDD1.n13 10.4732
R516 VDD1.n88 VDD1.n69 10.4732
R517 VDD1.n110 VDD1.n59 10.4732
R518 VDD1.n54 VDD1.n0 9.69747
R519 VDD1.n29 VDD1.n28 9.69747
R520 VDD1.n85 VDD1.n84 9.69747
R521 VDD1.n111 VDD1.n57 9.69747
R522 VDD1.n56 VDD1.n55 9.45567
R523 VDD1.n113 VDD1.n112 9.45567
R524 VDD1.n22 VDD1.n21 9.3005
R525 VDD1.n24 VDD1.n23 9.3005
R526 VDD1.n15 VDD1.n14 9.3005
R527 VDD1.n30 VDD1.n29 9.3005
R528 VDD1.n32 VDD1.n31 9.3005
R529 VDD1.n10 VDD1.n9 9.3005
R530 VDD1.n38 VDD1.n37 9.3005
R531 VDD1.n40 VDD1.n39 9.3005
R532 VDD1.n55 VDD1.n54 9.3005
R533 VDD1.n2 VDD1.n1 9.3005
R534 VDD1.n49 VDD1.n48 9.3005
R535 VDD1.n47 VDD1.n46 9.3005
R536 VDD1.n6 VDD1.n5 9.3005
R537 VDD1.n112 VDD1.n111 9.3005
R538 VDD1.n59 VDD1.n58 9.3005
R539 VDD1.n106 VDD1.n105 9.3005
R540 VDD1.n104 VDD1.n103 9.3005
R541 VDD1.n63 VDD1.n62 9.3005
R542 VDD1.n78 VDD1.n77 9.3005
R543 VDD1.n80 VDD1.n79 9.3005
R544 VDD1.n71 VDD1.n70 9.3005
R545 VDD1.n86 VDD1.n85 9.3005
R546 VDD1.n88 VDD1.n87 9.3005
R547 VDD1.n67 VDD1.n66 9.3005
R548 VDD1.n95 VDD1.n94 9.3005
R549 VDD1.n97 VDD1.n96 9.3005
R550 VDD1.n25 VDD1.n15 8.92171
R551 VDD1.n81 VDD1.n71 8.92171
R552 VDD1.n24 VDD1.n17 8.14595
R553 VDD1.n80 VDD1.n73 8.14595
R554 VDD1.n21 VDD1.n20 7.3702
R555 VDD1.n77 VDD1.n76 7.3702
R556 VDD1.n21 VDD1.n17 5.81868
R557 VDD1.n77 VDD1.n73 5.81868
R558 VDD1.n25 VDD1.n24 5.04292
R559 VDD1.n81 VDD1.n80 5.04292
R560 VDD1.n56 VDD1.n0 4.26717
R561 VDD1.n28 VDD1.n15 4.26717
R562 VDD1.n84 VDD1.n71 4.26717
R563 VDD1.n113 VDD1.n57 4.26717
R564 VDD1.n54 VDD1.n53 3.49141
R565 VDD1.n29 VDD1.n13 3.49141
R566 VDD1.n85 VDD1.n69 3.49141
R567 VDD1.n111 VDD1.n110 3.49141
R568 VDD1.n116 VDD1.t4 2.99359
R569 VDD1.n116 VDD1.t2 2.99359
R570 VDD1.n114 VDD1.t3 2.99359
R571 VDD1.n114 VDD1.t0 2.99359
R572 VDD1.n50 VDD1.n2 2.71565
R573 VDD1.n33 VDD1.n32 2.71565
R574 VDD1.n89 VDD1.n88 2.71565
R575 VDD1.n107 VDD1.n59 2.71565
R576 VDD1.n22 VDD1.n18 2.41282
R577 VDD1.n78 VDD1.n74 2.41282
R578 VDD1.n49 VDD1.n4 1.93989
R579 VDD1.n36 VDD1.n10 1.93989
R580 VDD1.n93 VDD1.n67 1.93989
R581 VDD1.n106 VDD1.n61 1.93989
R582 VDD1.n46 VDD1.n45 1.16414
R583 VDD1.n37 VDD1.n8 1.16414
R584 VDD1.n94 VDD1.n65 1.16414
R585 VDD1.n103 VDD1.n102 1.16414
R586 VDD1 VDD1.n117 0.528517
R587 VDD1.n42 VDD1.n6 0.388379
R588 VDD1.n41 VDD1.n40 0.388379
R589 VDD1.n98 VDD1.n97 0.388379
R590 VDD1.n99 VDD1.n63 0.388379
R591 VDD1.n55 VDD1.n1 0.155672
R592 VDD1.n48 VDD1.n1 0.155672
R593 VDD1.n48 VDD1.n47 0.155672
R594 VDD1.n47 VDD1.n5 0.155672
R595 VDD1.n39 VDD1.n5 0.155672
R596 VDD1.n39 VDD1.n38 0.155672
R597 VDD1.n38 VDD1.n9 0.155672
R598 VDD1.n31 VDD1.n9 0.155672
R599 VDD1.n31 VDD1.n30 0.155672
R600 VDD1.n30 VDD1.n14 0.155672
R601 VDD1.n23 VDD1.n14 0.155672
R602 VDD1.n23 VDD1.n22 0.155672
R603 VDD1.n79 VDD1.n78 0.155672
R604 VDD1.n79 VDD1.n70 0.155672
R605 VDD1.n86 VDD1.n70 0.155672
R606 VDD1.n87 VDD1.n86 0.155672
R607 VDD1.n87 VDD1.n66 0.155672
R608 VDD1.n95 VDD1.n66 0.155672
R609 VDD1.n96 VDD1.n95 0.155672
R610 VDD1.n96 VDD1.n62 0.155672
R611 VDD1.n104 VDD1.n62 0.155672
R612 VDD1.n105 VDD1.n104 0.155672
R613 VDD1.n105 VDD1.n58 0.155672
R614 VDD1.n112 VDD1.n58 0.155672
R615 B.n488 B.n69 585
R616 B.n490 B.n489 585
R617 B.n491 B.n68 585
R618 B.n493 B.n492 585
R619 B.n494 B.n67 585
R620 B.n496 B.n495 585
R621 B.n497 B.n66 585
R622 B.n499 B.n498 585
R623 B.n500 B.n65 585
R624 B.n502 B.n501 585
R625 B.n503 B.n64 585
R626 B.n505 B.n504 585
R627 B.n506 B.n63 585
R628 B.n508 B.n507 585
R629 B.n509 B.n62 585
R630 B.n511 B.n510 585
R631 B.n512 B.n61 585
R632 B.n514 B.n513 585
R633 B.n515 B.n60 585
R634 B.n517 B.n516 585
R635 B.n518 B.n59 585
R636 B.n520 B.n519 585
R637 B.n521 B.n58 585
R638 B.n523 B.n522 585
R639 B.n524 B.n57 585
R640 B.n526 B.n525 585
R641 B.n527 B.n56 585
R642 B.n529 B.n528 585
R643 B.n530 B.n55 585
R644 B.n532 B.n531 585
R645 B.n533 B.n54 585
R646 B.n535 B.n534 585
R647 B.n536 B.n53 585
R648 B.n538 B.n537 585
R649 B.n539 B.n52 585
R650 B.n541 B.n540 585
R651 B.n542 B.n51 585
R652 B.n544 B.n543 585
R653 B.n546 B.n545 585
R654 B.n547 B.n47 585
R655 B.n549 B.n548 585
R656 B.n550 B.n46 585
R657 B.n552 B.n551 585
R658 B.n553 B.n45 585
R659 B.n555 B.n554 585
R660 B.n556 B.n44 585
R661 B.n558 B.n557 585
R662 B.n559 B.n41 585
R663 B.n562 B.n561 585
R664 B.n563 B.n40 585
R665 B.n565 B.n564 585
R666 B.n566 B.n39 585
R667 B.n568 B.n567 585
R668 B.n569 B.n38 585
R669 B.n571 B.n570 585
R670 B.n572 B.n37 585
R671 B.n574 B.n573 585
R672 B.n575 B.n36 585
R673 B.n577 B.n576 585
R674 B.n578 B.n35 585
R675 B.n580 B.n579 585
R676 B.n581 B.n34 585
R677 B.n583 B.n582 585
R678 B.n584 B.n33 585
R679 B.n586 B.n585 585
R680 B.n587 B.n32 585
R681 B.n589 B.n588 585
R682 B.n590 B.n31 585
R683 B.n592 B.n591 585
R684 B.n593 B.n30 585
R685 B.n595 B.n594 585
R686 B.n596 B.n29 585
R687 B.n598 B.n597 585
R688 B.n599 B.n28 585
R689 B.n601 B.n600 585
R690 B.n602 B.n27 585
R691 B.n604 B.n603 585
R692 B.n605 B.n26 585
R693 B.n607 B.n606 585
R694 B.n608 B.n25 585
R695 B.n610 B.n609 585
R696 B.n611 B.n24 585
R697 B.n613 B.n612 585
R698 B.n614 B.n23 585
R699 B.n616 B.n615 585
R700 B.n617 B.n22 585
R701 B.n487 B.n486 585
R702 B.n485 B.n70 585
R703 B.n484 B.n483 585
R704 B.n482 B.n71 585
R705 B.n481 B.n480 585
R706 B.n479 B.n72 585
R707 B.n478 B.n477 585
R708 B.n476 B.n73 585
R709 B.n475 B.n474 585
R710 B.n473 B.n74 585
R711 B.n472 B.n471 585
R712 B.n470 B.n75 585
R713 B.n469 B.n468 585
R714 B.n467 B.n76 585
R715 B.n466 B.n465 585
R716 B.n464 B.n77 585
R717 B.n463 B.n462 585
R718 B.n461 B.n78 585
R719 B.n460 B.n459 585
R720 B.n458 B.n79 585
R721 B.n457 B.n456 585
R722 B.n455 B.n80 585
R723 B.n454 B.n453 585
R724 B.n452 B.n81 585
R725 B.n451 B.n450 585
R726 B.n449 B.n82 585
R727 B.n448 B.n447 585
R728 B.n446 B.n83 585
R729 B.n445 B.n444 585
R730 B.n443 B.n84 585
R731 B.n442 B.n441 585
R732 B.n440 B.n85 585
R733 B.n439 B.n438 585
R734 B.n437 B.n86 585
R735 B.n436 B.n435 585
R736 B.n434 B.n87 585
R737 B.n433 B.n432 585
R738 B.n431 B.n88 585
R739 B.n430 B.n429 585
R740 B.n428 B.n89 585
R741 B.n427 B.n426 585
R742 B.n425 B.n90 585
R743 B.n424 B.n423 585
R744 B.n422 B.n91 585
R745 B.n421 B.n420 585
R746 B.n419 B.n92 585
R747 B.n418 B.n417 585
R748 B.n416 B.n93 585
R749 B.n415 B.n414 585
R750 B.n413 B.n94 585
R751 B.n412 B.n411 585
R752 B.n410 B.n95 585
R753 B.n409 B.n408 585
R754 B.n407 B.n96 585
R755 B.n406 B.n405 585
R756 B.n404 B.n97 585
R757 B.n403 B.n402 585
R758 B.n401 B.n98 585
R759 B.n400 B.n399 585
R760 B.n398 B.n99 585
R761 B.n397 B.n396 585
R762 B.n395 B.n100 585
R763 B.n394 B.n393 585
R764 B.n392 B.n101 585
R765 B.n391 B.n390 585
R766 B.n389 B.n102 585
R767 B.n388 B.n387 585
R768 B.n386 B.n103 585
R769 B.n385 B.n384 585
R770 B.n383 B.n104 585
R771 B.n382 B.n381 585
R772 B.n380 B.n105 585
R773 B.n379 B.n378 585
R774 B.n377 B.n106 585
R775 B.n376 B.n375 585
R776 B.n374 B.n107 585
R777 B.n373 B.n372 585
R778 B.n371 B.n108 585
R779 B.n370 B.n369 585
R780 B.n368 B.n109 585
R781 B.n367 B.n366 585
R782 B.n236 B.n157 585
R783 B.n238 B.n237 585
R784 B.n239 B.n156 585
R785 B.n241 B.n240 585
R786 B.n242 B.n155 585
R787 B.n244 B.n243 585
R788 B.n245 B.n154 585
R789 B.n247 B.n246 585
R790 B.n248 B.n153 585
R791 B.n250 B.n249 585
R792 B.n251 B.n152 585
R793 B.n253 B.n252 585
R794 B.n254 B.n151 585
R795 B.n256 B.n255 585
R796 B.n257 B.n150 585
R797 B.n259 B.n258 585
R798 B.n260 B.n149 585
R799 B.n262 B.n261 585
R800 B.n263 B.n148 585
R801 B.n265 B.n264 585
R802 B.n266 B.n147 585
R803 B.n268 B.n267 585
R804 B.n269 B.n146 585
R805 B.n271 B.n270 585
R806 B.n272 B.n145 585
R807 B.n274 B.n273 585
R808 B.n275 B.n144 585
R809 B.n277 B.n276 585
R810 B.n278 B.n143 585
R811 B.n280 B.n279 585
R812 B.n281 B.n142 585
R813 B.n283 B.n282 585
R814 B.n284 B.n141 585
R815 B.n286 B.n285 585
R816 B.n287 B.n140 585
R817 B.n289 B.n288 585
R818 B.n290 B.n139 585
R819 B.n292 B.n291 585
R820 B.n294 B.n293 585
R821 B.n295 B.n135 585
R822 B.n297 B.n296 585
R823 B.n298 B.n134 585
R824 B.n300 B.n299 585
R825 B.n301 B.n133 585
R826 B.n303 B.n302 585
R827 B.n304 B.n132 585
R828 B.n306 B.n305 585
R829 B.n307 B.n129 585
R830 B.n310 B.n309 585
R831 B.n311 B.n128 585
R832 B.n313 B.n312 585
R833 B.n314 B.n127 585
R834 B.n316 B.n315 585
R835 B.n317 B.n126 585
R836 B.n319 B.n318 585
R837 B.n320 B.n125 585
R838 B.n322 B.n321 585
R839 B.n323 B.n124 585
R840 B.n325 B.n324 585
R841 B.n326 B.n123 585
R842 B.n328 B.n327 585
R843 B.n329 B.n122 585
R844 B.n331 B.n330 585
R845 B.n332 B.n121 585
R846 B.n334 B.n333 585
R847 B.n335 B.n120 585
R848 B.n337 B.n336 585
R849 B.n338 B.n119 585
R850 B.n340 B.n339 585
R851 B.n341 B.n118 585
R852 B.n343 B.n342 585
R853 B.n344 B.n117 585
R854 B.n346 B.n345 585
R855 B.n347 B.n116 585
R856 B.n349 B.n348 585
R857 B.n350 B.n115 585
R858 B.n352 B.n351 585
R859 B.n353 B.n114 585
R860 B.n355 B.n354 585
R861 B.n356 B.n113 585
R862 B.n358 B.n357 585
R863 B.n359 B.n112 585
R864 B.n361 B.n360 585
R865 B.n362 B.n111 585
R866 B.n364 B.n363 585
R867 B.n365 B.n110 585
R868 B.n235 B.n234 585
R869 B.n233 B.n158 585
R870 B.n232 B.n231 585
R871 B.n230 B.n159 585
R872 B.n229 B.n228 585
R873 B.n227 B.n160 585
R874 B.n226 B.n225 585
R875 B.n224 B.n161 585
R876 B.n223 B.n222 585
R877 B.n221 B.n162 585
R878 B.n220 B.n219 585
R879 B.n218 B.n163 585
R880 B.n217 B.n216 585
R881 B.n215 B.n164 585
R882 B.n214 B.n213 585
R883 B.n212 B.n165 585
R884 B.n211 B.n210 585
R885 B.n209 B.n166 585
R886 B.n208 B.n207 585
R887 B.n206 B.n167 585
R888 B.n205 B.n204 585
R889 B.n203 B.n168 585
R890 B.n202 B.n201 585
R891 B.n200 B.n169 585
R892 B.n199 B.n198 585
R893 B.n197 B.n170 585
R894 B.n196 B.n195 585
R895 B.n194 B.n171 585
R896 B.n193 B.n192 585
R897 B.n191 B.n172 585
R898 B.n190 B.n189 585
R899 B.n188 B.n173 585
R900 B.n187 B.n186 585
R901 B.n185 B.n174 585
R902 B.n184 B.n183 585
R903 B.n182 B.n175 585
R904 B.n181 B.n180 585
R905 B.n179 B.n176 585
R906 B.n178 B.n177 585
R907 B.n2 B.n0 585
R908 B.n677 B.n1 585
R909 B.n676 B.n675 585
R910 B.n674 B.n3 585
R911 B.n673 B.n672 585
R912 B.n671 B.n4 585
R913 B.n670 B.n669 585
R914 B.n668 B.n5 585
R915 B.n667 B.n666 585
R916 B.n665 B.n6 585
R917 B.n664 B.n663 585
R918 B.n662 B.n7 585
R919 B.n661 B.n660 585
R920 B.n659 B.n8 585
R921 B.n658 B.n657 585
R922 B.n656 B.n9 585
R923 B.n655 B.n654 585
R924 B.n653 B.n10 585
R925 B.n652 B.n651 585
R926 B.n650 B.n11 585
R927 B.n649 B.n648 585
R928 B.n647 B.n12 585
R929 B.n646 B.n645 585
R930 B.n644 B.n13 585
R931 B.n643 B.n642 585
R932 B.n641 B.n14 585
R933 B.n640 B.n639 585
R934 B.n638 B.n15 585
R935 B.n637 B.n636 585
R936 B.n635 B.n16 585
R937 B.n634 B.n633 585
R938 B.n632 B.n17 585
R939 B.n631 B.n630 585
R940 B.n629 B.n18 585
R941 B.n628 B.n627 585
R942 B.n626 B.n19 585
R943 B.n625 B.n624 585
R944 B.n623 B.n20 585
R945 B.n622 B.n621 585
R946 B.n620 B.n21 585
R947 B.n619 B.n618 585
R948 B.n679 B.n678 585
R949 B.n234 B.n157 526.135
R950 B.n618 B.n617 526.135
R951 B.n366 B.n365 526.135
R952 B.n486 B.n69 526.135
R953 B.n130 B.t2 408.058
R954 B.n48 B.t7 408.058
R955 B.n136 B.t5 408.058
R956 B.n42 B.t10 408.058
R957 B.n131 B.t1 355.308
R958 B.n49 B.t8 355.308
R959 B.n137 B.t4 355.308
R960 B.n43 B.t11 355.308
R961 B.n130 B.t0 317.216
R962 B.n136 B.t3 317.216
R963 B.n42 B.t9 317.216
R964 B.n48 B.t6 317.216
R965 B.n234 B.n233 163.367
R966 B.n233 B.n232 163.367
R967 B.n232 B.n159 163.367
R968 B.n228 B.n159 163.367
R969 B.n228 B.n227 163.367
R970 B.n227 B.n226 163.367
R971 B.n226 B.n161 163.367
R972 B.n222 B.n161 163.367
R973 B.n222 B.n221 163.367
R974 B.n221 B.n220 163.367
R975 B.n220 B.n163 163.367
R976 B.n216 B.n163 163.367
R977 B.n216 B.n215 163.367
R978 B.n215 B.n214 163.367
R979 B.n214 B.n165 163.367
R980 B.n210 B.n165 163.367
R981 B.n210 B.n209 163.367
R982 B.n209 B.n208 163.367
R983 B.n208 B.n167 163.367
R984 B.n204 B.n167 163.367
R985 B.n204 B.n203 163.367
R986 B.n203 B.n202 163.367
R987 B.n202 B.n169 163.367
R988 B.n198 B.n169 163.367
R989 B.n198 B.n197 163.367
R990 B.n197 B.n196 163.367
R991 B.n196 B.n171 163.367
R992 B.n192 B.n171 163.367
R993 B.n192 B.n191 163.367
R994 B.n191 B.n190 163.367
R995 B.n190 B.n173 163.367
R996 B.n186 B.n173 163.367
R997 B.n186 B.n185 163.367
R998 B.n185 B.n184 163.367
R999 B.n184 B.n175 163.367
R1000 B.n180 B.n175 163.367
R1001 B.n180 B.n179 163.367
R1002 B.n179 B.n178 163.367
R1003 B.n178 B.n2 163.367
R1004 B.n678 B.n2 163.367
R1005 B.n678 B.n677 163.367
R1006 B.n677 B.n676 163.367
R1007 B.n676 B.n3 163.367
R1008 B.n672 B.n3 163.367
R1009 B.n672 B.n671 163.367
R1010 B.n671 B.n670 163.367
R1011 B.n670 B.n5 163.367
R1012 B.n666 B.n5 163.367
R1013 B.n666 B.n665 163.367
R1014 B.n665 B.n664 163.367
R1015 B.n664 B.n7 163.367
R1016 B.n660 B.n7 163.367
R1017 B.n660 B.n659 163.367
R1018 B.n659 B.n658 163.367
R1019 B.n658 B.n9 163.367
R1020 B.n654 B.n9 163.367
R1021 B.n654 B.n653 163.367
R1022 B.n653 B.n652 163.367
R1023 B.n652 B.n11 163.367
R1024 B.n648 B.n11 163.367
R1025 B.n648 B.n647 163.367
R1026 B.n647 B.n646 163.367
R1027 B.n646 B.n13 163.367
R1028 B.n642 B.n13 163.367
R1029 B.n642 B.n641 163.367
R1030 B.n641 B.n640 163.367
R1031 B.n640 B.n15 163.367
R1032 B.n636 B.n15 163.367
R1033 B.n636 B.n635 163.367
R1034 B.n635 B.n634 163.367
R1035 B.n634 B.n17 163.367
R1036 B.n630 B.n17 163.367
R1037 B.n630 B.n629 163.367
R1038 B.n629 B.n628 163.367
R1039 B.n628 B.n19 163.367
R1040 B.n624 B.n19 163.367
R1041 B.n624 B.n623 163.367
R1042 B.n623 B.n622 163.367
R1043 B.n622 B.n21 163.367
R1044 B.n618 B.n21 163.367
R1045 B.n238 B.n157 163.367
R1046 B.n239 B.n238 163.367
R1047 B.n240 B.n239 163.367
R1048 B.n240 B.n155 163.367
R1049 B.n244 B.n155 163.367
R1050 B.n245 B.n244 163.367
R1051 B.n246 B.n245 163.367
R1052 B.n246 B.n153 163.367
R1053 B.n250 B.n153 163.367
R1054 B.n251 B.n250 163.367
R1055 B.n252 B.n251 163.367
R1056 B.n252 B.n151 163.367
R1057 B.n256 B.n151 163.367
R1058 B.n257 B.n256 163.367
R1059 B.n258 B.n257 163.367
R1060 B.n258 B.n149 163.367
R1061 B.n262 B.n149 163.367
R1062 B.n263 B.n262 163.367
R1063 B.n264 B.n263 163.367
R1064 B.n264 B.n147 163.367
R1065 B.n268 B.n147 163.367
R1066 B.n269 B.n268 163.367
R1067 B.n270 B.n269 163.367
R1068 B.n270 B.n145 163.367
R1069 B.n274 B.n145 163.367
R1070 B.n275 B.n274 163.367
R1071 B.n276 B.n275 163.367
R1072 B.n276 B.n143 163.367
R1073 B.n280 B.n143 163.367
R1074 B.n281 B.n280 163.367
R1075 B.n282 B.n281 163.367
R1076 B.n282 B.n141 163.367
R1077 B.n286 B.n141 163.367
R1078 B.n287 B.n286 163.367
R1079 B.n288 B.n287 163.367
R1080 B.n288 B.n139 163.367
R1081 B.n292 B.n139 163.367
R1082 B.n293 B.n292 163.367
R1083 B.n293 B.n135 163.367
R1084 B.n297 B.n135 163.367
R1085 B.n298 B.n297 163.367
R1086 B.n299 B.n298 163.367
R1087 B.n299 B.n133 163.367
R1088 B.n303 B.n133 163.367
R1089 B.n304 B.n303 163.367
R1090 B.n305 B.n304 163.367
R1091 B.n305 B.n129 163.367
R1092 B.n310 B.n129 163.367
R1093 B.n311 B.n310 163.367
R1094 B.n312 B.n311 163.367
R1095 B.n312 B.n127 163.367
R1096 B.n316 B.n127 163.367
R1097 B.n317 B.n316 163.367
R1098 B.n318 B.n317 163.367
R1099 B.n318 B.n125 163.367
R1100 B.n322 B.n125 163.367
R1101 B.n323 B.n322 163.367
R1102 B.n324 B.n323 163.367
R1103 B.n324 B.n123 163.367
R1104 B.n328 B.n123 163.367
R1105 B.n329 B.n328 163.367
R1106 B.n330 B.n329 163.367
R1107 B.n330 B.n121 163.367
R1108 B.n334 B.n121 163.367
R1109 B.n335 B.n334 163.367
R1110 B.n336 B.n335 163.367
R1111 B.n336 B.n119 163.367
R1112 B.n340 B.n119 163.367
R1113 B.n341 B.n340 163.367
R1114 B.n342 B.n341 163.367
R1115 B.n342 B.n117 163.367
R1116 B.n346 B.n117 163.367
R1117 B.n347 B.n346 163.367
R1118 B.n348 B.n347 163.367
R1119 B.n348 B.n115 163.367
R1120 B.n352 B.n115 163.367
R1121 B.n353 B.n352 163.367
R1122 B.n354 B.n353 163.367
R1123 B.n354 B.n113 163.367
R1124 B.n358 B.n113 163.367
R1125 B.n359 B.n358 163.367
R1126 B.n360 B.n359 163.367
R1127 B.n360 B.n111 163.367
R1128 B.n364 B.n111 163.367
R1129 B.n365 B.n364 163.367
R1130 B.n366 B.n109 163.367
R1131 B.n370 B.n109 163.367
R1132 B.n371 B.n370 163.367
R1133 B.n372 B.n371 163.367
R1134 B.n372 B.n107 163.367
R1135 B.n376 B.n107 163.367
R1136 B.n377 B.n376 163.367
R1137 B.n378 B.n377 163.367
R1138 B.n378 B.n105 163.367
R1139 B.n382 B.n105 163.367
R1140 B.n383 B.n382 163.367
R1141 B.n384 B.n383 163.367
R1142 B.n384 B.n103 163.367
R1143 B.n388 B.n103 163.367
R1144 B.n389 B.n388 163.367
R1145 B.n390 B.n389 163.367
R1146 B.n390 B.n101 163.367
R1147 B.n394 B.n101 163.367
R1148 B.n395 B.n394 163.367
R1149 B.n396 B.n395 163.367
R1150 B.n396 B.n99 163.367
R1151 B.n400 B.n99 163.367
R1152 B.n401 B.n400 163.367
R1153 B.n402 B.n401 163.367
R1154 B.n402 B.n97 163.367
R1155 B.n406 B.n97 163.367
R1156 B.n407 B.n406 163.367
R1157 B.n408 B.n407 163.367
R1158 B.n408 B.n95 163.367
R1159 B.n412 B.n95 163.367
R1160 B.n413 B.n412 163.367
R1161 B.n414 B.n413 163.367
R1162 B.n414 B.n93 163.367
R1163 B.n418 B.n93 163.367
R1164 B.n419 B.n418 163.367
R1165 B.n420 B.n419 163.367
R1166 B.n420 B.n91 163.367
R1167 B.n424 B.n91 163.367
R1168 B.n425 B.n424 163.367
R1169 B.n426 B.n425 163.367
R1170 B.n426 B.n89 163.367
R1171 B.n430 B.n89 163.367
R1172 B.n431 B.n430 163.367
R1173 B.n432 B.n431 163.367
R1174 B.n432 B.n87 163.367
R1175 B.n436 B.n87 163.367
R1176 B.n437 B.n436 163.367
R1177 B.n438 B.n437 163.367
R1178 B.n438 B.n85 163.367
R1179 B.n442 B.n85 163.367
R1180 B.n443 B.n442 163.367
R1181 B.n444 B.n443 163.367
R1182 B.n444 B.n83 163.367
R1183 B.n448 B.n83 163.367
R1184 B.n449 B.n448 163.367
R1185 B.n450 B.n449 163.367
R1186 B.n450 B.n81 163.367
R1187 B.n454 B.n81 163.367
R1188 B.n455 B.n454 163.367
R1189 B.n456 B.n455 163.367
R1190 B.n456 B.n79 163.367
R1191 B.n460 B.n79 163.367
R1192 B.n461 B.n460 163.367
R1193 B.n462 B.n461 163.367
R1194 B.n462 B.n77 163.367
R1195 B.n466 B.n77 163.367
R1196 B.n467 B.n466 163.367
R1197 B.n468 B.n467 163.367
R1198 B.n468 B.n75 163.367
R1199 B.n472 B.n75 163.367
R1200 B.n473 B.n472 163.367
R1201 B.n474 B.n473 163.367
R1202 B.n474 B.n73 163.367
R1203 B.n478 B.n73 163.367
R1204 B.n479 B.n478 163.367
R1205 B.n480 B.n479 163.367
R1206 B.n480 B.n71 163.367
R1207 B.n484 B.n71 163.367
R1208 B.n485 B.n484 163.367
R1209 B.n486 B.n485 163.367
R1210 B.n617 B.n616 163.367
R1211 B.n616 B.n23 163.367
R1212 B.n612 B.n23 163.367
R1213 B.n612 B.n611 163.367
R1214 B.n611 B.n610 163.367
R1215 B.n610 B.n25 163.367
R1216 B.n606 B.n25 163.367
R1217 B.n606 B.n605 163.367
R1218 B.n605 B.n604 163.367
R1219 B.n604 B.n27 163.367
R1220 B.n600 B.n27 163.367
R1221 B.n600 B.n599 163.367
R1222 B.n599 B.n598 163.367
R1223 B.n598 B.n29 163.367
R1224 B.n594 B.n29 163.367
R1225 B.n594 B.n593 163.367
R1226 B.n593 B.n592 163.367
R1227 B.n592 B.n31 163.367
R1228 B.n588 B.n31 163.367
R1229 B.n588 B.n587 163.367
R1230 B.n587 B.n586 163.367
R1231 B.n586 B.n33 163.367
R1232 B.n582 B.n33 163.367
R1233 B.n582 B.n581 163.367
R1234 B.n581 B.n580 163.367
R1235 B.n580 B.n35 163.367
R1236 B.n576 B.n35 163.367
R1237 B.n576 B.n575 163.367
R1238 B.n575 B.n574 163.367
R1239 B.n574 B.n37 163.367
R1240 B.n570 B.n37 163.367
R1241 B.n570 B.n569 163.367
R1242 B.n569 B.n568 163.367
R1243 B.n568 B.n39 163.367
R1244 B.n564 B.n39 163.367
R1245 B.n564 B.n563 163.367
R1246 B.n563 B.n562 163.367
R1247 B.n562 B.n41 163.367
R1248 B.n557 B.n41 163.367
R1249 B.n557 B.n556 163.367
R1250 B.n556 B.n555 163.367
R1251 B.n555 B.n45 163.367
R1252 B.n551 B.n45 163.367
R1253 B.n551 B.n550 163.367
R1254 B.n550 B.n549 163.367
R1255 B.n549 B.n47 163.367
R1256 B.n545 B.n47 163.367
R1257 B.n545 B.n544 163.367
R1258 B.n544 B.n51 163.367
R1259 B.n540 B.n51 163.367
R1260 B.n540 B.n539 163.367
R1261 B.n539 B.n538 163.367
R1262 B.n538 B.n53 163.367
R1263 B.n534 B.n53 163.367
R1264 B.n534 B.n533 163.367
R1265 B.n533 B.n532 163.367
R1266 B.n532 B.n55 163.367
R1267 B.n528 B.n55 163.367
R1268 B.n528 B.n527 163.367
R1269 B.n527 B.n526 163.367
R1270 B.n526 B.n57 163.367
R1271 B.n522 B.n57 163.367
R1272 B.n522 B.n521 163.367
R1273 B.n521 B.n520 163.367
R1274 B.n520 B.n59 163.367
R1275 B.n516 B.n59 163.367
R1276 B.n516 B.n515 163.367
R1277 B.n515 B.n514 163.367
R1278 B.n514 B.n61 163.367
R1279 B.n510 B.n61 163.367
R1280 B.n510 B.n509 163.367
R1281 B.n509 B.n508 163.367
R1282 B.n508 B.n63 163.367
R1283 B.n504 B.n63 163.367
R1284 B.n504 B.n503 163.367
R1285 B.n503 B.n502 163.367
R1286 B.n502 B.n65 163.367
R1287 B.n498 B.n65 163.367
R1288 B.n498 B.n497 163.367
R1289 B.n497 B.n496 163.367
R1290 B.n496 B.n67 163.367
R1291 B.n492 B.n67 163.367
R1292 B.n492 B.n491 163.367
R1293 B.n491 B.n490 163.367
R1294 B.n490 B.n69 163.367
R1295 B.n308 B.n131 59.5399
R1296 B.n138 B.n137 59.5399
R1297 B.n560 B.n43 59.5399
R1298 B.n50 B.n49 59.5399
R1299 B.n131 B.n130 52.752
R1300 B.n137 B.n136 52.752
R1301 B.n43 B.n42 52.752
R1302 B.n49 B.n48 52.752
R1303 B.n619 B.n22 34.1859
R1304 B.n488 B.n487 34.1859
R1305 B.n367 B.n110 34.1859
R1306 B.n236 B.n235 34.1859
R1307 B B.n679 18.0485
R1308 B.n615 B.n22 10.6151
R1309 B.n615 B.n614 10.6151
R1310 B.n614 B.n613 10.6151
R1311 B.n613 B.n24 10.6151
R1312 B.n609 B.n24 10.6151
R1313 B.n609 B.n608 10.6151
R1314 B.n608 B.n607 10.6151
R1315 B.n607 B.n26 10.6151
R1316 B.n603 B.n26 10.6151
R1317 B.n603 B.n602 10.6151
R1318 B.n602 B.n601 10.6151
R1319 B.n601 B.n28 10.6151
R1320 B.n597 B.n28 10.6151
R1321 B.n597 B.n596 10.6151
R1322 B.n596 B.n595 10.6151
R1323 B.n595 B.n30 10.6151
R1324 B.n591 B.n30 10.6151
R1325 B.n591 B.n590 10.6151
R1326 B.n590 B.n589 10.6151
R1327 B.n589 B.n32 10.6151
R1328 B.n585 B.n32 10.6151
R1329 B.n585 B.n584 10.6151
R1330 B.n584 B.n583 10.6151
R1331 B.n583 B.n34 10.6151
R1332 B.n579 B.n34 10.6151
R1333 B.n579 B.n578 10.6151
R1334 B.n578 B.n577 10.6151
R1335 B.n577 B.n36 10.6151
R1336 B.n573 B.n36 10.6151
R1337 B.n573 B.n572 10.6151
R1338 B.n572 B.n571 10.6151
R1339 B.n571 B.n38 10.6151
R1340 B.n567 B.n38 10.6151
R1341 B.n567 B.n566 10.6151
R1342 B.n566 B.n565 10.6151
R1343 B.n565 B.n40 10.6151
R1344 B.n561 B.n40 10.6151
R1345 B.n559 B.n558 10.6151
R1346 B.n558 B.n44 10.6151
R1347 B.n554 B.n44 10.6151
R1348 B.n554 B.n553 10.6151
R1349 B.n553 B.n552 10.6151
R1350 B.n552 B.n46 10.6151
R1351 B.n548 B.n46 10.6151
R1352 B.n548 B.n547 10.6151
R1353 B.n547 B.n546 10.6151
R1354 B.n543 B.n542 10.6151
R1355 B.n542 B.n541 10.6151
R1356 B.n541 B.n52 10.6151
R1357 B.n537 B.n52 10.6151
R1358 B.n537 B.n536 10.6151
R1359 B.n536 B.n535 10.6151
R1360 B.n535 B.n54 10.6151
R1361 B.n531 B.n54 10.6151
R1362 B.n531 B.n530 10.6151
R1363 B.n530 B.n529 10.6151
R1364 B.n529 B.n56 10.6151
R1365 B.n525 B.n56 10.6151
R1366 B.n525 B.n524 10.6151
R1367 B.n524 B.n523 10.6151
R1368 B.n523 B.n58 10.6151
R1369 B.n519 B.n58 10.6151
R1370 B.n519 B.n518 10.6151
R1371 B.n518 B.n517 10.6151
R1372 B.n517 B.n60 10.6151
R1373 B.n513 B.n60 10.6151
R1374 B.n513 B.n512 10.6151
R1375 B.n512 B.n511 10.6151
R1376 B.n511 B.n62 10.6151
R1377 B.n507 B.n62 10.6151
R1378 B.n507 B.n506 10.6151
R1379 B.n506 B.n505 10.6151
R1380 B.n505 B.n64 10.6151
R1381 B.n501 B.n64 10.6151
R1382 B.n501 B.n500 10.6151
R1383 B.n500 B.n499 10.6151
R1384 B.n499 B.n66 10.6151
R1385 B.n495 B.n66 10.6151
R1386 B.n495 B.n494 10.6151
R1387 B.n494 B.n493 10.6151
R1388 B.n493 B.n68 10.6151
R1389 B.n489 B.n68 10.6151
R1390 B.n489 B.n488 10.6151
R1391 B.n368 B.n367 10.6151
R1392 B.n369 B.n368 10.6151
R1393 B.n369 B.n108 10.6151
R1394 B.n373 B.n108 10.6151
R1395 B.n374 B.n373 10.6151
R1396 B.n375 B.n374 10.6151
R1397 B.n375 B.n106 10.6151
R1398 B.n379 B.n106 10.6151
R1399 B.n380 B.n379 10.6151
R1400 B.n381 B.n380 10.6151
R1401 B.n381 B.n104 10.6151
R1402 B.n385 B.n104 10.6151
R1403 B.n386 B.n385 10.6151
R1404 B.n387 B.n386 10.6151
R1405 B.n387 B.n102 10.6151
R1406 B.n391 B.n102 10.6151
R1407 B.n392 B.n391 10.6151
R1408 B.n393 B.n392 10.6151
R1409 B.n393 B.n100 10.6151
R1410 B.n397 B.n100 10.6151
R1411 B.n398 B.n397 10.6151
R1412 B.n399 B.n398 10.6151
R1413 B.n399 B.n98 10.6151
R1414 B.n403 B.n98 10.6151
R1415 B.n404 B.n403 10.6151
R1416 B.n405 B.n404 10.6151
R1417 B.n405 B.n96 10.6151
R1418 B.n409 B.n96 10.6151
R1419 B.n410 B.n409 10.6151
R1420 B.n411 B.n410 10.6151
R1421 B.n411 B.n94 10.6151
R1422 B.n415 B.n94 10.6151
R1423 B.n416 B.n415 10.6151
R1424 B.n417 B.n416 10.6151
R1425 B.n417 B.n92 10.6151
R1426 B.n421 B.n92 10.6151
R1427 B.n422 B.n421 10.6151
R1428 B.n423 B.n422 10.6151
R1429 B.n423 B.n90 10.6151
R1430 B.n427 B.n90 10.6151
R1431 B.n428 B.n427 10.6151
R1432 B.n429 B.n428 10.6151
R1433 B.n429 B.n88 10.6151
R1434 B.n433 B.n88 10.6151
R1435 B.n434 B.n433 10.6151
R1436 B.n435 B.n434 10.6151
R1437 B.n435 B.n86 10.6151
R1438 B.n439 B.n86 10.6151
R1439 B.n440 B.n439 10.6151
R1440 B.n441 B.n440 10.6151
R1441 B.n441 B.n84 10.6151
R1442 B.n445 B.n84 10.6151
R1443 B.n446 B.n445 10.6151
R1444 B.n447 B.n446 10.6151
R1445 B.n447 B.n82 10.6151
R1446 B.n451 B.n82 10.6151
R1447 B.n452 B.n451 10.6151
R1448 B.n453 B.n452 10.6151
R1449 B.n453 B.n80 10.6151
R1450 B.n457 B.n80 10.6151
R1451 B.n458 B.n457 10.6151
R1452 B.n459 B.n458 10.6151
R1453 B.n459 B.n78 10.6151
R1454 B.n463 B.n78 10.6151
R1455 B.n464 B.n463 10.6151
R1456 B.n465 B.n464 10.6151
R1457 B.n465 B.n76 10.6151
R1458 B.n469 B.n76 10.6151
R1459 B.n470 B.n469 10.6151
R1460 B.n471 B.n470 10.6151
R1461 B.n471 B.n74 10.6151
R1462 B.n475 B.n74 10.6151
R1463 B.n476 B.n475 10.6151
R1464 B.n477 B.n476 10.6151
R1465 B.n477 B.n72 10.6151
R1466 B.n481 B.n72 10.6151
R1467 B.n482 B.n481 10.6151
R1468 B.n483 B.n482 10.6151
R1469 B.n483 B.n70 10.6151
R1470 B.n487 B.n70 10.6151
R1471 B.n237 B.n236 10.6151
R1472 B.n237 B.n156 10.6151
R1473 B.n241 B.n156 10.6151
R1474 B.n242 B.n241 10.6151
R1475 B.n243 B.n242 10.6151
R1476 B.n243 B.n154 10.6151
R1477 B.n247 B.n154 10.6151
R1478 B.n248 B.n247 10.6151
R1479 B.n249 B.n248 10.6151
R1480 B.n249 B.n152 10.6151
R1481 B.n253 B.n152 10.6151
R1482 B.n254 B.n253 10.6151
R1483 B.n255 B.n254 10.6151
R1484 B.n255 B.n150 10.6151
R1485 B.n259 B.n150 10.6151
R1486 B.n260 B.n259 10.6151
R1487 B.n261 B.n260 10.6151
R1488 B.n261 B.n148 10.6151
R1489 B.n265 B.n148 10.6151
R1490 B.n266 B.n265 10.6151
R1491 B.n267 B.n266 10.6151
R1492 B.n267 B.n146 10.6151
R1493 B.n271 B.n146 10.6151
R1494 B.n272 B.n271 10.6151
R1495 B.n273 B.n272 10.6151
R1496 B.n273 B.n144 10.6151
R1497 B.n277 B.n144 10.6151
R1498 B.n278 B.n277 10.6151
R1499 B.n279 B.n278 10.6151
R1500 B.n279 B.n142 10.6151
R1501 B.n283 B.n142 10.6151
R1502 B.n284 B.n283 10.6151
R1503 B.n285 B.n284 10.6151
R1504 B.n285 B.n140 10.6151
R1505 B.n289 B.n140 10.6151
R1506 B.n290 B.n289 10.6151
R1507 B.n291 B.n290 10.6151
R1508 B.n295 B.n294 10.6151
R1509 B.n296 B.n295 10.6151
R1510 B.n296 B.n134 10.6151
R1511 B.n300 B.n134 10.6151
R1512 B.n301 B.n300 10.6151
R1513 B.n302 B.n301 10.6151
R1514 B.n302 B.n132 10.6151
R1515 B.n306 B.n132 10.6151
R1516 B.n307 B.n306 10.6151
R1517 B.n309 B.n128 10.6151
R1518 B.n313 B.n128 10.6151
R1519 B.n314 B.n313 10.6151
R1520 B.n315 B.n314 10.6151
R1521 B.n315 B.n126 10.6151
R1522 B.n319 B.n126 10.6151
R1523 B.n320 B.n319 10.6151
R1524 B.n321 B.n320 10.6151
R1525 B.n321 B.n124 10.6151
R1526 B.n325 B.n124 10.6151
R1527 B.n326 B.n325 10.6151
R1528 B.n327 B.n326 10.6151
R1529 B.n327 B.n122 10.6151
R1530 B.n331 B.n122 10.6151
R1531 B.n332 B.n331 10.6151
R1532 B.n333 B.n332 10.6151
R1533 B.n333 B.n120 10.6151
R1534 B.n337 B.n120 10.6151
R1535 B.n338 B.n337 10.6151
R1536 B.n339 B.n338 10.6151
R1537 B.n339 B.n118 10.6151
R1538 B.n343 B.n118 10.6151
R1539 B.n344 B.n343 10.6151
R1540 B.n345 B.n344 10.6151
R1541 B.n345 B.n116 10.6151
R1542 B.n349 B.n116 10.6151
R1543 B.n350 B.n349 10.6151
R1544 B.n351 B.n350 10.6151
R1545 B.n351 B.n114 10.6151
R1546 B.n355 B.n114 10.6151
R1547 B.n356 B.n355 10.6151
R1548 B.n357 B.n356 10.6151
R1549 B.n357 B.n112 10.6151
R1550 B.n361 B.n112 10.6151
R1551 B.n362 B.n361 10.6151
R1552 B.n363 B.n362 10.6151
R1553 B.n363 B.n110 10.6151
R1554 B.n235 B.n158 10.6151
R1555 B.n231 B.n158 10.6151
R1556 B.n231 B.n230 10.6151
R1557 B.n230 B.n229 10.6151
R1558 B.n229 B.n160 10.6151
R1559 B.n225 B.n160 10.6151
R1560 B.n225 B.n224 10.6151
R1561 B.n224 B.n223 10.6151
R1562 B.n223 B.n162 10.6151
R1563 B.n219 B.n162 10.6151
R1564 B.n219 B.n218 10.6151
R1565 B.n218 B.n217 10.6151
R1566 B.n217 B.n164 10.6151
R1567 B.n213 B.n164 10.6151
R1568 B.n213 B.n212 10.6151
R1569 B.n212 B.n211 10.6151
R1570 B.n211 B.n166 10.6151
R1571 B.n207 B.n166 10.6151
R1572 B.n207 B.n206 10.6151
R1573 B.n206 B.n205 10.6151
R1574 B.n205 B.n168 10.6151
R1575 B.n201 B.n168 10.6151
R1576 B.n201 B.n200 10.6151
R1577 B.n200 B.n199 10.6151
R1578 B.n199 B.n170 10.6151
R1579 B.n195 B.n170 10.6151
R1580 B.n195 B.n194 10.6151
R1581 B.n194 B.n193 10.6151
R1582 B.n193 B.n172 10.6151
R1583 B.n189 B.n172 10.6151
R1584 B.n189 B.n188 10.6151
R1585 B.n188 B.n187 10.6151
R1586 B.n187 B.n174 10.6151
R1587 B.n183 B.n174 10.6151
R1588 B.n183 B.n182 10.6151
R1589 B.n182 B.n181 10.6151
R1590 B.n181 B.n176 10.6151
R1591 B.n177 B.n176 10.6151
R1592 B.n177 B.n0 10.6151
R1593 B.n675 B.n1 10.6151
R1594 B.n675 B.n674 10.6151
R1595 B.n674 B.n673 10.6151
R1596 B.n673 B.n4 10.6151
R1597 B.n669 B.n4 10.6151
R1598 B.n669 B.n668 10.6151
R1599 B.n668 B.n667 10.6151
R1600 B.n667 B.n6 10.6151
R1601 B.n663 B.n6 10.6151
R1602 B.n663 B.n662 10.6151
R1603 B.n662 B.n661 10.6151
R1604 B.n661 B.n8 10.6151
R1605 B.n657 B.n8 10.6151
R1606 B.n657 B.n656 10.6151
R1607 B.n656 B.n655 10.6151
R1608 B.n655 B.n10 10.6151
R1609 B.n651 B.n10 10.6151
R1610 B.n651 B.n650 10.6151
R1611 B.n650 B.n649 10.6151
R1612 B.n649 B.n12 10.6151
R1613 B.n645 B.n12 10.6151
R1614 B.n645 B.n644 10.6151
R1615 B.n644 B.n643 10.6151
R1616 B.n643 B.n14 10.6151
R1617 B.n639 B.n14 10.6151
R1618 B.n639 B.n638 10.6151
R1619 B.n638 B.n637 10.6151
R1620 B.n637 B.n16 10.6151
R1621 B.n633 B.n16 10.6151
R1622 B.n633 B.n632 10.6151
R1623 B.n632 B.n631 10.6151
R1624 B.n631 B.n18 10.6151
R1625 B.n627 B.n18 10.6151
R1626 B.n627 B.n626 10.6151
R1627 B.n626 B.n625 10.6151
R1628 B.n625 B.n20 10.6151
R1629 B.n621 B.n20 10.6151
R1630 B.n621 B.n620 10.6151
R1631 B.n620 B.n619 10.6151
R1632 B.n561 B.n560 9.36635
R1633 B.n543 B.n50 9.36635
R1634 B.n291 B.n138 9.36635
R1635 B.n309 B.n308 9.36635
R1636 B.n679 B.n0 2.81026
R1637 B.n679 B.n1 2.81026
R1638 B.n560 B.n559 1.24928
R1639 B.n546 B.n50 1.24928
R1640 B.n294 B.n138 1.24928
R1641 B.n308 B.n307 1.24928
R1642 VN.n25 VN.n14 161.3
R1643 VN.n24 VN.n23 161.3
R1644 VN.n22 VN.n15 161.3
R1645 VN.n21 VN.n20 161.3
R1646 VN.n19 VN.n16 161.3
R1647 VN.n11 VN.n0 161.3
R1648 VN.n10 VN.n9 161.3
R1649 VN.n8 VN.n1 161.3
R1650 VN.n7 VN.n6 161.3
R1651 VN.n5 VN.n2 161.3
R1652 VN.n3 VN.t0 143.528
R1653 VN.n17 VN.t3 143.528
R1654 VN.n4 VN.t2 109.51
R1655 VN.n12 VN.t5 109.51
R1656 VN.n18 VN.t4 109.51
R1657 VN.n26 VN.t1 109.51
R1658 VN.n13 VN.n12 100.088
R1659 VN.n27 VN.n26 100.088
R1660 VN.n6 VN.n1 54.1398
R1661 VN.n20 VN.n15 54.1398
R1662 VN.n4 VN.n3 48.0647
R1663 VN.n18 VN.n17 48.0647
R1664 VN VN.n27 47.2482
R1665 VN.n10 VN.n1 27.0143
R1666 VN.n24 VN.n15 27.0143
R1667 VN.n5 VN.n4 24.5923
R1668 VN.n6 VN.n5 24.5923
R1669 VN.n11 VN.n10 24.5923
R1670 VN.n20 VN.n19 24.5923
R1671 VN.n19 VN.n18 24.5923
R1672 VN.n25 VN.n24 24.5923
R1673 VN.n12 VN.n11 10.8209
R1674 VN.n26 VN.n25 10.8209
R1675 VN.n17 VN.n16 6.7696
R1676 VN.n3 VN.n2 6.7696
R1677 VN.n27 VN.n14 0.278335
R1678 VN.n13 VN.n0 0.278335
R1679 VN.n23 VN.n14 0.189894
R1680 VN.n23 VN.n22 0.189894
R1681 VN.n22 VN.n21 0.189894
R1682 VN.n21 VN.n16 0.189894
R1683 VN.n7 VN.n2 0.189894
R1684 VN.n8 VN.n7 0.189894
R1685 VN.n9 VN.n8 0.189894
R1686 VN.n9 VN.n0 0.189894
R1687 VN VN.n13 0.153485
R1688 VDD2.n111 VDD2.n59 756.745
R1689 VDD2.n52 VDD2.n0 756.745
R1690 VDD2.n112 VDD2.n111 585
R1691 VDD2.n110 VDD2.n109 585
R1692 VDD2.n63 VDD2.n62 585
R1693 VDD2.n104 VDD2.n103 585
R1694 VDD2.n102 VDD2.n101 585
R1695 VDD2.n100 VDD2.n66 585
R1696 VDD2.n70 VDD2.n67 585
R1697 VDD2.n95 VDD2.n94 585
R1698 VDD2.n93 VDD2.n92 585
R1699 VDD2.n72 VDD2.n71 585
R1700 VDD2.n87 VDD2.n86 585
R1701 VDD2.n85 VDD2.n84 585
R1702 VDD2.n76 VDD2.n75 585
R1703 VDD2.n79 VDD2.n78 585
R1704 VDD2.n19 VDD2.n18 585
R1705 VDD2.n16 VDD2.n15 585
R1706 VDD2.n25 VDD2.n24 585
R1707 VDD2.n27 VDD2.n26 585
R1708 VDD2.n12 VDD2.n11 585
R1709 VDD2.n33 VDD2.n32 585
R1710 VDD2.n36 VDD2.n35 585
R1711 VDD2.n34 VDD2.n8 585
R1712 VDD2.n41 VDD2.n7 585
R1713 VDD2.n43 VDD2.n42 585
R1714 VDD2.n45 VDD2.n44 585
R1715 VDD2.n4 VDD2.n3 585
R1716 VDD2.n51 VDD2.n50 585
R1717 VDD2.n53 VDD2.n52 585
R1718 VDD2.t4 VDD2.n77 329.038
R1719 VDD2.t5 VDD2.n17 329.038
R1720 VDD2.n111 VDD2.n110 171.744
R1721 VDD2.n110 VDD2.n62 171.744
R1722 VDD2.n103 VDD2.n62 171.744
R1723 VDD2.n103 VDD2.n102 171.744
R1724 VDD2.n102 VDD2.n66 171.744
R1725 VDD2.n70 VDD2.n66 171.744
R1726 VDD2.n94 VDD2.n70 171.744
R1727 VDD2.n94 VDD2.n93 171.744
R1728 VDD2.n93 VDD2.n71 171.744
R1729 VDD2.n86 VDD2.n71 171.744
R1730 VDD2.n86 VDD2.n85 171.744
R1731 VDD2.n85 VDD2.n75 171.744
R1732 VDD2.n78 VDD2.n75 171.744
R1733 VDD2.n18 VDD2.n15 171.744
R1734 VDD2.n25 VDD2.n15 171.744
R1735 VDD2.n26 VDD2.n25 171.744
R1736 VDD2.n26 VDD2.n11 171.744
R1737 VDD2.n33 VDD2.n11 171.744
R1738 VDD2.n35 VDD2.n33 171.744
R1739 VDD2.n35 VDD2.n34 171.744
R1740 VDD2.n34 VDD2.n7 171.744
R1741 VDD2.n43 VDD2.n7 171.744
R1742 VDD2.n44 VDD2.n43 171.744
R1743 VDD2.n44 VDD2.n3 171.744
R1744 VDD2.n51 VDD2.n3 171.744
R1745 VDD2.n52 VDD2.n51 171.744
R1746 VDD2.n78 VDD2.t4 85.8723
R1747 VDD2.n18 VDD2.t5 85.8723
R1748 VDD2.n58 VDD2.n57 79.8878
R1749 VDD2 VDD2.n117 79.8849
R1750 VDD2.n58 VDD2.n56 54.0583
R1751 VDD2.n116 VDD2.n115 52.355
R1752 VDD2.n116 VDD2.n58 40.6981
R1753 VDD2.n101 VDD2.n100 13.1884
R1754 VDD2.n42 VDD2.n41 13.1884
R1755 VDD2.n104 VDD2.n65 12.8005
R1756 VDD2.n99 VDD2.n67 12.8005
R1757 VDD2.n40 VDD2.n8 12.8005
R1758 VDD2.n45 VDD2.n6 12.8005
R1759 VDD2.n105 VDD2.n63 12.0247
R1760 VDD2.n96 VDD2.n95 12.0247
R1761 VDD2.n37 VDD2.n36 12.0247
R1762 VDD2.n46 VDD2.n4 12.0247
R1763 VDD2.n109 VDD2.n108 11.249
R1764 VDD2.n92 VDD2.n69 11.249
R1765 VDD2.n32 VDD2.n10 11.249
R1766 VDD2.n50 VDD2.n49 11.249
R1767 VDD2.n79 VDD2.n77 10.7239
R1768 VDD2.n19 VDD2.n17 10.7239
R1769 VDD2.n112 VDD2.n61 10.4732
R1770 VDD2.n91 VDD2.n72 10.4732
R1771 VDD2.n31 VDD2.n12 10.4732
R1772 VDD2.n53 VDD2.n2 10.4732
R1773 VDD2.n113 VDD2.n59 9.69747
R1774 VDD2.n88 VDD2.n87 9.69747
R1775 VDD2.n28 VDD2.n27 9.69747
R1776 VDD2.n54 VDD2.n0 9.69747
R1777 VDD2.n115 VDD2.n114 9.45567
R1778 VDD2.n56 VDD2.n55 9.45567
R1779 VDD2.n81 VDD2.n80 9.3005
R1780 VDD2.n83 VDD2.n82 9.3005
R1781 VDD2.n74 VDD2.n73 9.3005
R1782 VDD2.n89 VDD2.n88 9.3005
R1783 VDD2.n91 VDD2.n90 9.3005
R1784 VDD2.n69 VDD2.n68 9.3005
R1785 VDD2.n97 VDD2.n96 9.3005
R1786 VDD2.n99 VDD2.n98 9.3005
R1787 VDD2.n114 VDD2.n113 9.3005
R1788 VDD2.n61 VDD2.n60 9.3005
R1789 VDD2.n108 VDD2.n107 9.3005
R1790 VDD2.n106 VDD2.n105 9.3005
R1791 VDD2.n65 VDD2.n64 9.3005
R1792 VDD2.n55 VDD2.n54 9.3005
R1793 VDD2.n2 VDD2.n1 9.3005
R1794 VDD2.n49 VDD2.n48 9.3005
R1795 VDD2.n47 VDD2.n46 9.3005
R1796 VDD2.n6 VDD2.n5 9.3005
R1797 VDD2.n21 VDD2.n20 9.3005
R1798 VDD2.n23 VDD2.n22 9.3005
R1799 VDD2.n14 VDD2.n13 9.3005
R1800 VDD2.n29 VDD2.n28 9.3005
R1801 VDD2.n31 VDD2.n30 9.3005
R1802 VDD2.n10 VDD2.n9 9.3005
R1803 VDD2.n38 VDD2.n37 9.3005
R1804 VDD2.n40 VDD2.n39 9.3005
R1805 VDD2.n84 VDD2.n74 8.92171
R1806 VDD2.n24 VDD2.n14 8.92171
R1807 VDD2.n83 VDD2.n76 8.14595
R1808 VDD2.n23 VDD2.n16 8.14595
R1809 VDD2.n80 VDD2.n79 7.3702
R1810 VDD2.n20 VDD2.n19 7.3702
R1811 VDD2.n80 VDD2.n76 5.81868
R1812 VDD2.n20 VDD2.n16 5.81868
R1813 VDD2.n84 VDD2.n83 5.04292
R1814 VDD2.n24 VDD2.n23 5.04292
R1815 VDD2.n115 VDD2.n59 4.26717
R1816 VDD2.n87 VDD2.n74 4.26717
R1817 VDD2.n27 VDD2.n14 4.26717
R1818 VDD2.n56 VDD2.n0 4.26717
R1819 VDD2.n113 VDD2.n112 3.49141
R1820 VDD2.n88 VDD2.n72 3.49141
R1821 VDD2.n28 VDD2.n12 3.49141
R1822 VDD2.n54 VDD2.n53 3.49141
R1823 VDD2.n117 VDD2.t1 2.99359
R1824 VDD2.n117 VDD2.t2 2.99359
R1825 VDD2.n57 VDD2.t3 2.99359
R1826 VDD2.n57 VDD2.t0 2.99359
R1827 VDD2.n109 VDD2.n61 2.71565
R1828 VDD2.n92 VDD2.n91 2.71565
R1829 VDD2.n32 VDD2.n31 2.71565
R1830 VDD2.n50 VDD2.n2 2.71565
R1831 VDD2.n81 VDD2.n77 2.41282
R1832 VDD2.n21 VDD2.n17 2.41282
R1833 VDD2.n108 VDD2.n63 1.93989
R1834 VDD2.n95 VDD2.n69 1.93989
R1835 VDD2.n36 VDD2.n10 1.93989
R1836 VDD2.n49 VDD2.n4 1.93989
R1837 VDD2 VDD2.n116 1.81731
R1838 VDD2.n105 VDD2.n104 1.16414
R1839 VDD2.n96 VDD2.n67 1.16414
R1840 VDD2.n37 VDD2.n8 1.16414
R1841 VDD2.n46 VDD2.n45 1.16414
R1842 VDD2.n101 VDD2.n65 0.388379
R1843 VDD2.n100 VDD2.n99 0.388379
R1844 VDD2.n41 VDD2.n40 0.388379
R1845 VDD2.n42 VDD2.n6 0.388379
R1846 VDD2.n114 VDD2.n60 0.155672
R1847 VDD2.n107 VDD2.n60 0.155672
R1848 VDD2.n107 VDD2.n106 0.155672
R1849 VDD2.n106 VDD2.n64 0.155672
R1850 VDD2.n98 VDD2.n64 0.155672
R1851 VDD2.n98 VDD2.n97 0.155672
R1852 VDD2.n97 VDD2.n68 0.155672
R1853 VDD2.n90 VDD2.n68 0.155672
R1854 VDD2.n90 VDD2.n89 0.155672
R1855 VDD2.n89 VDD2.n73 0.155672
R1856 VDD2.n82 VDD2.n73 0.155672
R1857 VDD2.n82 VDD2.n81 0.155672
R1858 VDD2.n22 VDD2.n21 0.155672
R1859 VDD2.n22 VDD2.n13 0.155672
R1860 VDD2.n29 VDD2.n13 0.155672
R1861 VDD2.n30 VDD2.n29 0.155672
R1862 VDD2.n30 VDD2.n9 0.155672
R1863 VDD2.n38 VDD2.n9 0.155672
R1864 VDD2.n39 VDD2.n38 0.155672
R1865 VDD2.n39 VDD2.n5 0.155672
R1866 VDD2.n47 VDD2.n5 0.155672
R1867 VDD2.n48 VDD2.n47 0.155672
R1868 VDD2.n48 VDD2.n1 0.155672
R1869 VDD2.n55 VDD2.n1 0.155672
C0 w_n3146_n3140# VDD1 2.16157f
C1 B VP 1.79009f
C2 VP VN 6.50842f
C3 VTAIL VDD1 7.27759f
C4 VP VDD2 0.440787f
C5 B w_n3146_n3140# 9.06637f
C6 w_n3146_n3140# VN 5.88325f
C7 B VTAIL 3.3552f
C8 VTAIL VN 6.1775f
C9 B VDD1 1.94865f
C10 w_n3146_n3140# VDD2 2.23997f
C11 VDD1 VN 0.150811f
C12 VTAIL VDD2 7.32706f
C13 VDD1 VDD2 1.32525f
C14 B VN 1.11304f
C15 B VDD2 2.01771f
C16 VDD2 VN 6.01935f
C17 w_n3146_n3140# VP 6.2894f
C18 VTAIL VP 6.19178f
C19 VDD1 VP 6.30629f
C20 VTAIL w_n3146_n3140# 2.79972f
C21 VDD2 VSUBS 1.811235f
C22 VDD1 VSUBS 1.688467f
C23 VTAIL VSUBS 1.108774f
C24 VN VSUBS 5.58368f
C25 VP VSUBS 2.729487f
C26 B VSUBS 4.331182f
C27 w_n3146_n3140# VSUBS 0.121826p
C28 VDD2.n0 VSUBS 0.03201f
C29 VDD2.n1 VSUBS 0.028153f
C30 VDD2.n2 VSUBS 0.015128f
C31 VDD2.n3 VSUBS 0.035757f
C32 VDD2.n4 VSUBS 0.016018f
C33 VDD2.n5 VSUBS 0.028153f
C34 VDD2.n6 VSUBS 0.015128f
C35 VDD2.n7 VSUBS 0.035757f
C36 VDD2.n8 VSUBS 0.016018f
C37 VDD2.n9 VSUBS 0.028153f
C38 VDD2.n10 VSUBS 0.015128f
C39 VDD2.n11 VSUBS 0.035757f
C40 VDD2.n12 VSUBS 0.016018f
C41 VDD2.n13 VSUBS 0.028153f
C42 VDD2.n14 VSUBS 0.015128f
C43 VDD2.n15 VSUBS 0.035757f
C44 VDD2.n16 VSUBS 0.016018f
C45 VDD2.n17 VSUBS 0.207223f
C46 VDD2.t5 VSUBS 0.076961f
C47 VDD2.n18 VSUBS 0.026818f
C48 VDD2.n19 VSUBS 0.026899f
C49 VDD2.n20 VSUBS 0.015128f
C50 VDD2.n21 VSUBS 1.24259f
C51 VDD2.n22 VSUBS 0.028153f
C52 VDD2.n23 VSUBS 0.015128f
C53 VDD2.n24 VSUBS 0.016018f
C54 VDD2.n25 VSUBS 0.035757f
C55 VDD2.n26 VSUBS 0.035757f
C56 VDD2.n27 VSUBS 0.016018f
C57 VDD2.n28 VSUBS 0.015128f
C58 VDD2.n29 VSUBS 0.028153f
C59 VDD2.n30 VSUBS 0.028153f
C60 VDD2.n31 VSUBS 0.015128f
C61 VDD2.n32 VSUBS 0.016018f
C62 VDD2.n33 VSUBS 0.035757f
C63 VDD2.n34 VSUBS 0.035757f
C64 VDD2.n35 VSUBS 0.035757f
C65 VDD2.n36 VSUBS 0.016018f
C66 VDD2.n37 VSUBS 0.015128f
C67 VDD2.n38 VSUBS 0.028153f
C68 VDD2.n39 VSUBS 0.028153f
C69 VDD2.n40 VSUBS 0.015128f
C70 VDD2.n41 VSUBS 0.015573f
C71 VDD2.n42 VSUBS 0.015573f
C72 VDD2.n43 VSUBS 0.035757f
C73 VDD2.n44 VSUBS 0.035757f
C74 VDD2.n45 VSUBS 0.016018f
C75 VDD2.n46 VSUBS 0.015128f
C76 VDD2.n47 VSUBS 0.028153f
C77 VDD2.n48 VSUBS 0.028153f
C78 VDD2.n49 VSUBS 0.015128f
C79 VDD2.n50 VSUBS 0.016018f
C80 VDD2.n51 VSUBS 0.035757f
C81 VDD2.n52 VSUBS 0.090229f
C82 VDD2.n53 VSUBS 0.016018f
C83 VDD2.n54 VSUBS 0.015128f
C84 VDD2.n55 VSUBS 0.071997f
C85 VDD2.n56 VSUBS 0.071845f
C86 VDD2.t3 VSUBS 0.241605f
C87 VDD2.t0 VSUBS 0.241605f
C88 VDD2.n57 VSUBS 1.86933f
C89 VDD2.n58 VSUBS 3.11273f
C90 VDD2.n59 VSUBS 0.03201f
C91 VDD2.n60 VSUBS 0.028153f
C92 VDD2.n61 VSUBS 0.015128f
C93 VDD2.n62 VSUBS 0.035757f
C94 VDD2.n63 VSUBS 0.016018f
C95 VDD2.n64 VSUBS 0.028153f
C96 VDD2.n65 VSUBS 0.015128f
C97 VDD2.n66 VSUBS 0.035757f
C98 VDD2.n67 VSUBS 0.016018f
C99 VDD2.n68 VSUBS 0.028153f
C100 VDD2.n69 VSUBS 0.015128f
C101 VDD2.n70 VSUBS 0.035757f
C102 VDD2.n71 VSUBS 0.035757f
C103 VDD2.n72 VSUBS 0.016018f
C104 VDD2.n73 VSUBS 0.028153f
C105 VDD2.n74 VSUBS 0.015128f
C106 VDD2.n75 VSUBS 0.035757f
C107 VDD2.n76 VSUBS 0.016018f
C108 VDD2.n77 VSUBS 0.207223f
C109 VDD2.t4 VSUBS 0.076961f
C110 VDD2.n78 VSUBS 0.026818f
C111 VDD2.n79 VSUBS 0.026899f
C112 VDD2.n80 VSUBS 0.015128f
C113 VDD2.n81 VSUBS 1.24259f
C114 VDD2.n82 VSUBS 0.028153f
C115 VDD2.n83 VSUBS 0.015128f
C116 VDD2.n84 VSUBS 0.016018f
C117 VDD2.n85 VSUBS 0.035757f
C118 VDD2.n86 VSUBS 0.035757f
C119 VDD2.n87 VSUBS 0.016018f
C120 VDD2.n88 VSUBS 0.015128f
C121 VDD2.n89 VSUBS 0.028153f
C122 VDD2.n90 VSUBS 0.028153f
C123 VDD2.n91 VSUBS 0.015128f
C124 VDD2.n92 VSUBS 0.016018f
C125 VDD2.n93 VSUBS 0.035757f
C126 VDD2.n94 VSUBS 0.035757f
C127 VDD2.n95 VSUBS 0.016018f
C128 VDD2.n96 VSUBS 0.015128f
C129 VDD2.n97 VSUBS 0.028153f
C130 VDD2.n98 VSUBS 0.028153f
C131 VDD2.n99 VSUBS 0.015128f
C132 VDD2.n100 VSUBS 0.015573f
C133 VDD2.n101 VSUBS 0.015573f
C134 VDD2.n102 VSUBS 0.035757f
C135 VDD2.n103 VSUBS 0.035757f
C136 VDD2.n104 VSUBS 0.016018f
C137 VDD2.n105 VSUBS 0.015128f
C138 VDD2.n106 VSUBS 0.028153f
C139 VDD2.n107 VSUBS 0.028153f
C140 VDD2.n108 VSUBS 0.015128f
C141 VDD2.n109 VSUBS 0.016018f
C142 VDD2.n110 VSUBS 0.035757f
C143 VDD2.n111 VSUBS 0.090229f
C144 VDD2.n112 VSUBS 0.016018f
C145 VDD2.n113 VSUBS 0.015128f
C146 VDD2.n114 VSUBS 0.071997f
C147 VDD2.n115 VSUBS 0.065132f
C148 VDD2.n116 VSUBS 2.72433f
C149 VDD2.t1 VSUBS 0.241605f
C150 VDD2.t2 VSUBS 0.241605f
C151 VDD2.n117 VSUBS 1.86929f
C152 VN.n0 VSUBS 0.04312f
C153 VN.t5 VSUBS 2.30617f
C154 VN.n1 VSUBS 0.035618f
C155 VN.n2 VSUBS 0.309205f
C156 VN.t2 VSUBS 2.30617f
C157 VN.t0 VSUBS 2.54647f
C158 VN.n3 VSUBS 0.886572f
C159 VN.n4 VSUBS 0.929869f
C160 VN.n5 VSUBS 0.060655f
C161 VN.n6 VSUBS 0.05706f
C162 VN.n7 VSUBS 0.032709f
C163 VN.n8 VSUBS 0.032709f
C164 VN.n9 VSUBS 0.032709f
C165 VN.n10 VSUBS 0.063071f
C166 VN.n11 VSUBS 0.043887f
C167 VN.n12 VSUBS 0.924133f
C168 VN.n13 VSUBS 0.05046f
C169 VN.n14 VSUBS 0.04312f
C170 VN.t1 VSUBS 2.30617f
C171 VN.n15 VSUBS 0.035618f
C172 VN.n16 VSUBS 0.309205f
C173 VN.t4 VSUBS 2.30617f
C174 VN.t3 VSUBS 2.54647f
C175 VN.n17 VSUBS 0.886572f
C176 VN.n18 VSUBS 0.929869f
C177 VN.n19 VSUBS 0.060655f
C178 VN.n20 VSUBS 0.05706f
C179 VN.n21 VSUBS 0.032709f
C180 VN.n22 VSUBS 0.032709f
C181 VN.n23 VSUBS 0.032709f
C182 VN.n24 VSUBS 0.063071f
C183 VN.n25 VSUBS 0.043887f
C184 VN.n26 VSUBS 0.924133f
C185 VN.n27 VSUBS 1.6721f
C186 B.n0 VSUBS 0.004737f
C187 B.n1 VSUBS 0.004737f
C188 B.n2 VSUBS 0.007491f
C189 B.n3 VSUBS 0.007491f
C190 B.n4 VSUBS 0.007491f
C191 B.n5 VSUBS 0.007491f
C192 B.n6 VSUBS 0.007491f
C193 B.n7 VSUBS 0.007491f
C194 B.n8 VSUBS 0.007491f
C195 B.n9 VSUBS 0.007491f
C196 B.n10 VSUBS 0.007491f
C197 B.n11 VSUBS 0.007491f
C198 B.n12 VSUBS 0.007491f
C199 B.n13 VSUBS 0.007491f
C200 B.n14 VSUBS 0.007491f
C201 B.n15 VSUBS 0.007491f
C202 B.n16 VSUBS 0.007491f
C203 B.n17 VSUBS 0.007491f
C204 B.n18 VSUBS 0.007491f
C205 B.n19 VSUBS 0.007491f
C206 B.n20 VSUBS 0.007491f
C207 B.n21 VSUBS 0.007491f
C208 B.n22 VSUBS 0.01851f
C209 B.n23 VSUBS 0.007491f
C210 B.n24 VSUBS 0.007491f
C211 B.n25 VSUBS 0.007491f
C212 B.n26 VSUBS 0.007491f
C213 B.n27 VSUBS 0.007491f
C214 B.n28 VSUBS 0.007491f
C215 B.n29 VSUBS 0.007491f
C216 B.n30 VSUBS 0.007491f
C217 B.n31 VSUBS 0.007491f
C218 B.n32 VSUBS 0.007491f
C219 B.n33 VSUBS 0.007491f
C220 B.n34 VSUBS 0.007491f
C221 B.n35 VSUBS 0.007491f
C222 B.n36 VSUBS 0.007491f
C223 B.n37 VSUBS 0.007491f
C224 B.n38 VSUBS 0.007491f
C225 B.n39 VSUBS 0.007491f
C226 B.n40 VSUBS 0.007491f
C227 B.n41 VSUBS 0.007491f
C228 B.t11 VSUBS 0.199281f
C229 B.t10 VSUBS 0.23035f
C230 B.t9 VSUBS 1.26577f
C231 B.n42 VSUBS 0.368277f
C232 B.n43 VSUBS 0.251017f
C233 B.n44 VSUBS 0.007491f
C234 B.n45 VSUBS 0.007491f
C235 B.n46 VSUBS 0.007491f
C236 B.n47 VSUBS 0.007491f
C237 B.t8 VSUBS 0.199284f
C238 B.t7 VSUBS 0.230353f
C239 B.t6 VSUBS 1.26577f
C240 B.n48 VSUBS 0.368275f
C241 B.n49 VSUBS 0.251014f
C242 B.n50 VSUBS 0.017356f
C243 B.n51 VSUBS 0.007491f
C244 B.n52 VSUBS 0.007491f
C245 B.n53 VSUBS 0.007491f
C246 B.n54 VSUBS 0.007491f
C247 B.n55 VSUBS 0.007491f
C248 B.n56 VSUBS 0.007491f
C249 B.n57 VSUBS 0.007491f
C250 B.n58 VSUBS 0.007491f
C251 B.n59 VSUBS 0.007491f
C252 B.n60 VSUBS 0.007491f
C253 B.n61 VSUBS 0.007491f
C254 B.n62 VSUBS 0.007491f
C255 B.n63 VSUBS 0.007491f
C256 B.n64 VSUBS 0.007491f
C257 B.n65 VSUBS 0.007491f
C258 B.n66 VSUBS 0.007491f
C259 B.n67 VSUBS 0.007491f
C260 B.n68 VSUBS 0.007491f
C261 B.n69 VSUBS 0.01851f
C262 B.n70 VSUBS 0.007491f
C263 B.n71 VSUBS 0.007491f
C264 B.n72 VSUBS 0.007491f
C265 B.n73 VSUBS 0.007491f
C266 B.n74 VSUBS 0.007491f
C267 B.n75 VSUBS 0.007491f
C268 B.n76 VSUBS 0.007491f
C269 B.n77 VSUBS 0.007491f
C270 B.n78 VSUBS 0.007491f
C271 B.n79 VSUBS 0.007491f
C272 B.n80 VSUBS 0.007491f
C273 B.n81 VSUBS 0.007491f
C274 B.n82 VSUBS 0.007491f
C275 B.n83 VSUBS 0.007491f
C276 B.n84 VSUBS 0.007491f
C277 B.n85 VSUBS 0.007491f
C278 B.n86 VSUBS 0.007491f
C279 B.n87 VSUBS 0.007491f
C280 B.n88 VSUBS 0.007491f
C281 B.n89 VSUBS 0.007491f
C282 B.n90 VSUBS 0.007491f
C283 B.n91 VSUBS 0.007491f
C284 B.n92 VSUBS 0.007491f
C285 B.n93 VSUBS 0.007491f
C286 B.n94 VSUBS 0.007491f
C287 B.n95 VSUBS 0.007491f
C288 B.n96 VSUBS 0.007491f
C289 B.n97 VSUBS 0.007491f
C290 B.n98 VSUBS 0.007491f
C291 B.n99 VSUBS 0.007491f
C292 B.n100 VSUBS 0.007491f
C293 B.n101 VSUBS 0.007491f
C294 B.n102 VSUBS 0.007491f
C295 B.n103 VSUBS 0.007491f
C296 B.n104 VSUBS 0.007491f
C297 B.n105 VSUBS 0.007491f
C298 B.n106 VSUBS 0.007491f
C299 B.n107 VSUBS 0.007491f
C300 B.n108 VSUBS 0.007491f
C301 B.n109 VSUBS 0.007491f
C302 B.n110 VSUBS 0.01851f
C303 B.n111 VSUBS 0.007491f
C304 B.n112 VSUBS 0.007491f
C305 B.n113 VSUBS 0.007491f
C306 B.n114 VSUBS 0.007491f
C307 B.n115 VSUBS 0.007491f
C308 B.n116 VSUBS 0.007491f
C309 B.n117 VSUBS 0.007491f
C310 B.n118 VSUBS 0.007491f
C311 B.n119 VSUBS 0.007491f
C312 B.n120 VSUBS 0.007491f
C313 B.n121 VSUBS 0.007491f
C314 B.n122 VSUBS 0.007491f
C315 B.n123 VSUBS 0.007491f
C316 B.n124 VSUBS 0.007491f
C317 B.n125 VSUBS 0.007491f
C318 B.n126 VSUBS 0.007491f
C319 B.n127 VSUBS 0.007491f
C320 B.n128 VSUBS 0.007491f
C321 B.n129 VSUBS 0.007491f
C322 B.t1 VSUBS 0.199284f
C323 B.t2 VSUBS 0.230353f
C324 B.t0 VSUBS 1.26577f
C325 B.n130 VSUBS 0.368275f
C326 B.n131 VSUBS 0.251014f
C327 B.n132 VSUBS 0.007491f
C328 B.n133 VSUBS 0.007491f
C329 B.n134 VSUBS 0.007491f
C330 B.n135 VSUBS 0.007491f
C331 B.t4 VSUBS 0.199281f
C332 B.t5 VSUBS 0.23035f
C333 B.t3 VSUBS 1.26577f
C334 B.n136 VSUBS 0.368277f
C335 B.n137 VSUBS 0.251017f
C336 B.n138 VSUBS 0.017356f
C337 B.n139 VSUBS 0.007491f
C338 B.n140 VSUBS 0.007491f
C339 B.n141 VSUBS 0.007491f
C340 B.n142 VSUBS 0.007491f
C341 B.n143 VSUBS 0.007491f
C342 B.n144 VSUBS 0.007491f
C343 B.n145 VSUBS 0.007491f
C344 B.n146 VSUBS 0.007491f
C345 B.n147 VSUBS 0.007491f
C346 B.n148 VSUBS 0.007491f
C347 B.n149 VSUBS 0.007491f
C348 B.n150 VSUBS 0.007491f
C349 B.n151 VSUBS 0.007491f
C350 B.n152 VSUBS 0.007491f
C351 B.n153 VSUBS 0.007491f
C352 B.n154 VSUBS 0.007491f
C353 B.n155 VSUBS 0.007491f
C354 B.n156 VSUBS 0.007491f
C355 B.n157 VSUBS 0.01851f
C356 B.n158 VSUBS 0.007491f
C357 B.n159 VSUBS 0.007491f
C358 B.n160 VSUBS 0.007491f
C359 B.n161 VSUBS 0.007491f
C360 B.n162 VSUBS 0.007491f
C361 B.n163 VSUBS 0.007491f
C362 B.n164 VSUBS 0.007491f
C363 B.n165 VSUBS 0.007491f
C364 B.n166 VSUBS 0.007491f
C365 B.n167 VSUBS 0.007491f
C366 B.n168 VSUBS 0.007491f
C367 B.n169 VSUBS 0.007491f
C368 B.n170 VSUBS 0.007491f
C369 B.n171 VSUBS 0.007491f
C370 B.n172 VSUBS 0.007491f
C371 B.n173 VSUBS 0.007491f
C372 B.n174 VSUBS 0.007491f
C373 B.n175 VSUBS 0.007491f
C374 B.n176 VSUBS 0.007491f
C375 B.n177 VSUBS 0.007491f
C376 B.n178 VSUBS 0.007491f
C377 B.n179 VSUBS 0.007491f
C378 B.n180 VSUBS 0.007491f
C379 B.n181 VSUBS 0.007491f
C380 B.n182 VSUBS 0.007491f
C381 B.n183 VSUBS 0.007491f
C382 B.n184 VSUBS 0.007491f
C383 B.n185 VSUBS 0.007491f
C384 B.n186 VSUBS 0.007491f
C385 B.n187 VSUBS 0.007491f
C386 B.n188 VSUBS 0.007491f
C387 B.n189 VSUBS 0.007491f
C388 B.n190 VSUBS 0.007491f
C389 B.n191 VSUBS 0.007491f
C390 B.n192 VSUBS 0.007491f
C391 B.n193 VSUBS 0.007491f
C392 B.n194 VSUBS 0.007491f
C393 B.n195 VSUBS 0.007491f
C394 B.n196 VSUBS 0.007491f
C395 B.n197 VSUBS 0.007491f
C396 B.n198 VSUBS 0.007491f
C397 B.n199 VSUBS 0.007491f
C398 B.n200 VSUBS 0.007491f
C399 B.n201 VSUBS 0.007491f
C400 B.n202 VSUBS 0.007491f
C401 B.n203 VSUBS 0.007491f
C402 B.n204 VSUBS 0.007491f
C403 B.n205 VSUBS 0.007491f
C404 B.n206 VSUBS 0.007491f
C405 B.n207 VSUBS 0.007491f
C406 B.n208 VSUBS 0.007491f
C407 B.n209 VSUBS 0.007491f
C408 B.n210 VSUBS 0.007491f
C409 B.n211 VSUBS 0.007491f
C410 B.n212 VSUBS 0.007491f
C411 B.n213 VSUBS 0.007491f
C412 B.n214 VSUBS 0.007491f
C413 B.n215 VSUBS 0.007491f
C414 B.n216 VSUBS 0.007491f
C415 B.n217 VSUBS 0.007491f
C416 B.n218 VSUBS 0.007491f
C417 B.n219 VSUBS 0.007491f
C418 B.n220 VSUBS 0.007491f
C419 B.n221 VSUBS 0.007491f
C420 B.n222 VSUBS 0.007491f
C421 B.n223 VSUBS 0.007491f
C422 B.n224 VSUBS 0.007491f
C423 B.n225 VSUBS 0.007491f
C424 B.n226 VSUBS 0.007491f
C425 B.n227 VSUBS 0.007491f
C426 B.n228 VSUBS 0.007491f
C427 B.n229 VSUBS 0.007491f
C428 B.n230 VSUBS 0.007491f
C429 B.n231 VSUBS 0.007491f
C430 B.n232 VSUBS 0.007491f
C431 B.n233 VSUBS 0.007491f
C432 B.n234 VSUBS 0.017624f
C433 B.n235 VSUBS 0.017624f
C434 B.n236 VSUBS 0.01851f
C435 B.n237 VSUBS 0.007491f
C436 B.n238 VSUBS 0.007491f
C437 B.n239 VSUBS 0.007491f
C438 B.n240 VSUBS 0.007491f
C439 B.n241 VSUBS 0.007491f
C440 B.n242 VSUBS 0.007491f
C441 B.n243 VSUBS 0.007491f
C442 B.n244 VSUBS 0.007491f
C443 B.n245 VSUBS 0.007491f
C444 B.n246 VSUBS 0.007491f
C445 B.n247 VSUBS 0.007491f
C446 B.n248 VSUBS 0.007491f
C447 B.n249 VSUBS 0.007491f
C448 B.n250 VSUBS 0.007491f
C449 B.n251 VSUBS 0.007491f
C450 B.n252 VSUBS 0.007491f
C451 B.n253 VSUBS 0.007491f
C452 B.n254 VSUBS 0.007491f
C453 B.n255 VSUBS 0.007491f
C454 B.n256 VSUBS 0.007491f
C455 B.n257 VSUBS 0.007491f
C456 B.n258 VSUBS 0.007491f
C457 B.n259 VSUBS 0.007491f
C458 B.n260 VSUBS 0.007491f
C459 B.n261 VSUBS 0.007491f
C460 B.n262 VSUBS 0.007491f
C461 B.n263 VSUBS 0.007491f
C462 B.n264 VSUBS 0.007491f
C463 B.n265 VSUBS 0.007491f
C464 B.n266 VSUBS 0.007491f
C465 B.n267 VSUBS 0.007491f
C466 B.n268 VSUBS 0.007491f
C467 B.n269 VSUBS 0.007491f
C468 B.n270 VSUBS 0.007491f
C469 B.n271 VSUBS 0.007491f
C470 B.n272 VSUBS 0.007491f
C471 B.n273 VSUBS 0.007491f
C472 B.n274 VSUBS 0.007491f
C473 B.n275 VSUBS 0.007491f
C474 B.n276 VSUBS 0.007491f
C475 B.n277 VSUBS 0.007491f
C476 B.n278 VSUBS 0.007491f
C477 B.n279 VSUBS 0.007491f
C478 B.n280 VSUBS 0.007491f
C479 B.n281 VSUBS 0.007491f
C480 B.n282 VSUBS 0.007491f
C481 B.n283 VSUBS 0.007491f
C482 B.n284 VSUBS 0.007491f
C483 B.n285 VSUBS 0.007491f
C484 B.n286 VSUBS 0.007491f
C485 B.n287 VSUBS 0.007491f
C486 B.n288 VSUBS 0.007491f
C487 B.n289 VSUBS 0.007491f
C488 B.n290 VSUBS 0.007491f
C489 B.n291 VSUBS 0.007051f
C490 B.n292 VSUBS 0.007491f
C491 B.n293 VSUBS 0.007491f
C492 B.n294 VSUBS 0.004186f
C493 B.n295 VSUBS 0.007491f
C494 B.n296 VSUBS 0.007491f
C495 B.n297 VSUBS 0.007491f
C496 B.n298 VSUBS 0.007491f
C497 B.n299 VSUBS 0.007491f
C498 B.n300 VSUBS 0.007491f
C499 B.n301 VSUBS 0.007491f
C500 B.n302 VSUBS 0.007491f
C501 B.n303 VSUBS 0.007491f
C502 B.n304 VSUBS 0.007491f
C503 B.n305 VSUBS 0.007491f
C504 B.n306 VSUBS 0.007491f
C505 B.n307 VSUBS 0.004186f
C506 B.n308 VSUBS 0.017356f
C507 B.n309 VSUBS 0.007051f
C508 B.n310 VSUBS 0.007491f
C509 B.n311 VSUBS 0.007491f
C510 B.n312 VSUBS 0.007491f
C511 B.n313 VSUBS 0.007491f
C512 B.n314 VSUBS 0.007491f
C513 B.n315 VSUBS 0.007491f
C514 B.n316 VSUBS 0.007491f
C515 B.n317 VSUBS 0.007491f
C516 B.n318 VSUBS 0.007491f
C517 B.n319 VSUBS 0.007491f
C518 B.n320 VSUBS 0.007491f
C519 B.n321 VSUBS 0.007491f
C520 B.n322 VSUBS 0.007491f
C521 B.n323 VSUBS 0.007491f
C522 B.n324 VSUBS 0.007491f
C523 B.n325 VSUBS 0.007491f
C524 B.n326 VSUBS 0.007491f
C525 B.n327 VSUBS 0.007491f
C526 B.n328 VSUBS 0.007491f
C527 B.n329 VSUBS 0.007491f
C528 B.n330 VSUBS 0.007491f
C529 B.n331 VSUBS 0.007491f
C530 B.n332 VSUBS 0.007491f
C531 B.n333 VSUBS 0.007491f
C532 B.n334 VSUBS 0.007491f
C533 B.n335 VSUBS 0.007491f
C534 B.n336 VSUBS 0.007491f
C535 B.n337 VSUBS 0.007491f
C536 B.n338 VSUBS 0.007491f
C537 B.n339 VSUBS 0.007491f
C538 B.n340 VSUBS 0.007491f
C539 B.n341 VSUBS 0.007491f
C540 B.n342 VSUBS 0.007491f
C541 B.n343 VSUBS 0.007491f
C542 B.n344 VSUBS 0.007491f
C543 B.n345 VSUBS 0.007491f
C544 B.n346 VSUBS 0.007491f
C545 B.n347 VSUBS 0.007491f
C546 B.n348 VSUBS 0.007491f
C547 B.n349 VSUBS 0.007491f
C548 B.n350 VSUBS 0.007491f
C549 B.n351 VSUBS 0.007491f
C550 B.n352 VSUBS 0.007491f
C551 B.n353 VSUBS 0.007491f
C552 B.n354 VSUBS 0.007491f
C553 B.n355 VSUBS 0.007491f
C554 B.n356 VSUBS 0.007491f
C555 B.n357 VSUBS 0.007491f
C556 B.n358 VSUBS 0.007491f
C557 B.n359 VSUBS 0.007491f
C558 B.n360 VSUBS 0.007491f
C559 B.n361 VSUBS 0.007491f
C560 B.n362 VSUBS 0.007491f
C561 B.n363 VSUBS 0.007491f
C562 B.n364 VSUBS 0.007491f
C563 B.n365 VSUBS 0.01851f
C564 B.n366 VSUBS 0.017624f
C565 B.n367 VSUBS 0.017624f
C566 B.n368 VSUBS 0.007491f
C567 B.n369 VSUBS 0.007491f
C568 B.n370 VSUBS 0.007491f
C569 B.n371 VSUBS 0.007491f
C570 B.n372 VSUBS 0.007491f
C571 B.n373 VSUBS 0.007491f
C572 B.n374 VSUBS 0.007491f
C573 B.n375 VSUBS 0.007491f
C574 B.n376 VSUBS 0.007491f
C575 B.n377 VSUBS 0.007491f
C576 B.n378 VSUBS 0.007491f
C577 B.n379 VSUBS 0.007491f
C578 B.n380 VSUBS 0.007491f
C579 B.n381 VSUBS 0.007491f
C580 B.n382 VSUBS 0.007491f
C581 B.n383 VSUBS 0.007491f
C582 B.n384 VSUBS 0.007491f
C583 B.n385 VSUBS 0.007491f
C584 B.n386 VSUBS 0.007491f
C585 B.n387 VSUBS 0.007491f
C586 B.n388 VSUBS 0.007491f
C587 B.n389 VSUBS 0.007491f
C588 B.n390 VSUBS 0.007491f
C589 B.n391 VSUBS 0.007491f
C590 B.n392 VSUBS 0.007491f
C591 B.n393 VSUBS 0.007491f
C592 B.n394 VSUBS 0.007491f
C593 B.n395 VSUBS 0.007491f
C594 B.n396 VSUBS 0.007491f
C595 B.n397 VSUBS 0.007491f
C596 B.n398 VSUBS 0.007491f
C597 B.n399 VSUBS 0.007491f
C598 B.n400 VSUBS 0.007491f
C599 B.n401 VSUBS 0.007491f
C600 B.n402 VSUBS 0.007491f
C601 B.n403 VSUBS 0.007491f
C602 B.n404 VSUBS 0.007491f
C603 B.n405 VSUBS 0.007491f
C604 B.n406 VSUBS 0.007491f
C605 B.n407 VSUBS 0.007491f
C606 B.n408 VSUBS 0.007491f
C607 B.n409 VSUBS 0.007491f
C608 B.n410 VSUBS 0.007491f
C609 B.n411 VSUBS 0.007491f
C610 B.n412 VSUBS 0.007491f
C611 B.n413 VSUBS 0.007491f
C612 B.n414 VSUBS 0.007491f
C613 B.n415 VSUBS 0.007491f
C614 B.n416 VSUBS 0.007491f
C615 B.n417 VSUBS 0.007491f
C616 B.n418 VSUBS 0.007491f
C617 B.n419 VSUBS 0.007491f
C618 B.n420 VSUBS 0.007491f
C619 B.n421 VSUBS 0.007491f
C620 B.n422 VSUBS 0.007491f
C621 B.n423 VSUBS 0.007491f
C622 B.n424 VSUBS 0.007491f
C623 B.n425 VSUBS 0.007491f
C624 B.n426 VSUBS 0.007491f
C625 B.n427 VSUBS 0.007491f
C626 B.n428 VSUBS 0.007491f
C627 B.n429 VSUBS 0.007491f
C628 B.n430 VSUBS 0.007491f
C629 B.n431 VSUBS 0.007491f
C630 B.n432 VSUBS 0.007491f
C631 B.n433 VSUBS 0.007491f
C632 B.n434 VSUBS 0.007491f
C633 B.n435 VSUBS 0.007491f
C634 B.n436 VSUBS 0.007491f
C635 B.n437 VSUBS 0.007491f
C636 B.n438 VSUBS 0.007491f
C637 B.n439 VSUBS 0.007491f
C638 B.n440 VSUBS 0.007491f
C639 B.n441 VSUBS 0.007491f
C640 B.n442 VSUBS 0.007491f
C641 B.n443 VSUBS 0.007491f
C642 B.n444 VSUBS 0.007491f
C643 B.n445 VSUBS 0.007491f
C644 B.n446 VSUBS 0.007491f
C645 B.n447 VSUBS 0.007491f
C646 B.n448 VSUBS 0.007491f
C647 B.n449 VSUBS 0.007491f
C648 B.n450 VSUBS 0.007491f
C649 B.n451 VSUBS 0.007491f
C650 B.n452 VSUBS 0.007491f
C651 B.n453 VSUBS 0.007491f
C652 B.n454 VSUBS 0.007491f
C653 B.n455 VSUBS 0.007491f
C654 B.n456 VSUBS 0.007491f
C655 B.n457 VSUBS 0.007491f
C656 B.n458 VSUBS 0.007491f
C657 B.n459 VSUBS 0.007491f
C658 B.n460 VSUBS 0.007491f
C659 B.n461 VSUBS 0.007491f
C660 B.n462 VSUBS 0.007491f
C661 B.n463 VSUBS 0.007491f
C662 B.n464 VSUBS 0.007491f
C663 B.n465 VSUBS 0.007491f
C664 B.n466 VSUBS 0.007491f
C665 B.n467 VSUBS 0.007491f
C666 B.n468 VSUBS 0.007491f
C667 B.n469 VSUBS 0.007491f
C668 B.n470 VSUBS 0.007491f
C669 B.n471 VSUBS 0.007491f
C670 B.n472 VSUBS 0.007491f
C671 B.n473 VSUBS 0.007491f
C672 B.n474 VSUBS 0.007491f
C673 B.n475 VSUBS 0.007491f
C674 B.n476 VSUBS 0.007491f
C675 B.n477 VSUBS 0.007491f
C676 B.n478 VSUBS 0.007491f
C677 B.n479 VSUBS 0.007491f
C678 B.n480 VSUBS 0.007491f
C679 B.n481 VSUBS 0.007491f
C680 B.n482 VSUBS 0.007491f
C681 B.n483 VSUBS 0.007491f
C682 B.n484 VSUBS 0.007491f
C683 B.n485 VSUBS 0.007491f
C684 B.n486 VSUBS 0.017624f
C685 B.n487 VSUBS 0.018469f
C686 B.n488 VSUBS 0.017665f
C687 B.n489 VSUBS 0.007491f
C688 B.n490 VSUBS 0.007491f
C689 B.n491 VSUBS 0.007491f
C690 B.n492 VSUBS 0.007491f
C691 B.n493 VSUBS 0.007491f
C692 B.n494 VSUBS 0.007491f
C693 B.n495 VSUBS 0.007491f
C694 B.n496 VSUBS 0.007491f
C695 B.n497 VSUBS 0.007491f
C696 B.n498 VSUBS 0.007491f
C697 B.n499 VSUBS 0.007491f
C698 B.n500 VSUBS 0.007491f
C699 B.n501 VSUBS 0.007491f
C700 B.n502 VSUBS 0.007491f
C701 B.n503 VSUBS 0.007491f
C702 B.n504 VSUBS 0.007491f
C703 B.n505 VSUBS 0.007491f
C704 B.n506 VSUBS 0.007491f
C705 B.n507 VSUBS 0.007491f
C706 B.n508 VSUBS 0.007491f
C707 B.n509 VSUBS 0.007491f
C708 B.n510 VSUBS 0.007491f
C709 B.n511 VSUBS 0.007491f
C710 B.n512 VSUBS 0.007491f
C711 B.n513 VSUBS 0.007491f
C712 B.n514 VSUBS 0.007491f
C713 B.n515 VSUBS 0.007491f
C714 B.n516 VSUBS 0.007491f
C715 B.n517 VSUBS 0.007491f
C716 B.n518 VSUBS 0.007491f
C717 B.n519 VSUBS 0.007491f
C718 B.n520 VSUBS 0.007491f
C719 B.n521 VSUBS 0.007491f
C720 B.n522 VSUBS 0.007491f
C721 B.n523 VSUBS 0.007491f
C722 B.n524 VSUBS 0.007491f
C723 B.n525 VSUBS 0.007491f
C724 B.n526 VSUBS 0.007491f
C725 B.n527 VSUBS 0.007491f
C726 B.n528 VSUBS 0.007491f
C727 B.n529 VSUBS 0.007491f
C728 B.n530 VSUBS 0.007491f
C729 B.n531 VSUBS 0.007491f
C730 B.n532 VSUBS 0.007491f
C731 B.n533 VSUBS 0.007491f
C732 B.n534 VSUBS 0.007491f
C733 B.n535 VSUBS 0.007491f
C734 B.n536 VSUBS 0.007491f
C735 B.n537 VSUBS 0.007491f
C736 B.n538 VSUBS 0.007491f
C737 B.n539 VSUBS 0.007491f
C738 B.n540 VSUBS 0.007491f
C739 B.n541 VSUBS 0.007491f
C740 B.n542 VSUBS 0.007491f
C741 B.n543 VSUBS 0.007051f
C742 B.n544 VSUBS 0.007491f
C743 B.n545 VSUBS 0.007491f
C744 B.n546 VSUBS 0.004186f
C745 B.n547 VSUBS 0.007491f
C746 B.n548 VSUBS 0.007491f
C747 B.n549 VSUBS 0.007491f
C748 B.n550 VSUBS 0.007491f
C749 B.n551 VSUBS 0.007491f
C750 B.n552 VSUBS 0.007491f
C751 B.n553 VSUBS 0.007491f
C752 B.n554 VSUBS 0.007491f
C753 B.n555 VSUBS 0.007491f
C754 B.n556 VSUBS 0.007491f
C755 B.n557 VSUBS 0.007491f
C756 B.n558 VSUBS 0.007491f
C757 B.n559 VSUBS 0.004186f
C758 B.n560 VSUBS 0.017356f
C759 B.n561 VSUBS 0.007051f
C760 B.n562 VSUBS 0.007491f
C761 B.n563 VSUBS 0.007491f
C762 B.n564 VSUBS 0.007491f
C763 B.n565 VSUBS 0.007491f
C764 B.n566 VSUBS 0.007491f
C765 B.n567 VSUBS 0.007491f
C766 B.n568 VSUBS 0.007491f
C767 B.n569 VSUBS 0.007491f
C768 B.n570 VSUBS 0.007491f
C769 B.n571 VSUBS 0.007491f
C770 B.n572 VSUBS 0.007491f
C771 B.n573 VSUBS 0.007491f
C772 B.n574 VSUBS 0.007491f
C773 B.n575 VSUBS 0.007491f
C774 B.n576 VSUBS 0.007491f
C775 B.n577 VSUBS 0.007491f
C776 B.n578 VSUBS 0.007491f
C777 B.n579 VSUBS 0.007491f
C778 B.n580 VSUBS 0.007491f
C779 B.n581 VSUBS 0.007491f
C780 B.n582 VSUBS 0.007491f
C781 B.n583 VSUBS 0.007491f
C782 B.n584 VSUBS 0.007491f
C783 B.n585 VSUBS 0.007491f
C784 B.n586 VSUBS 0.007491f
C785 B.n587 VSUBS 0.007491f
C786 B.n588 VSUBS 0.007491f
C787 B.n589 VSUBS 0.007491f
C788 B.n590 VSUBS 0.007491f
C789 B.n591 VSUBS 0.007491f
C790 B.n592 VSUBS 0.007491f
C791 B.n593 VSUBS 0.007491f
C792 B.n594 VSUBS 0.007491f
C793 B.n595 VSUBS 0.007491f
C794 B.n596 VSUBS 0.007491f
C795 B.n597 VSUBS 0.007491f
C796 B.n598 VSUBS 0.007491f
C797 B.n599 VSUBS 0.007491f
C798 B.n600 VSUBS 0.007491f
C799 B.n601 VSUBS 0.007491f
C800 B.n602 VSUBS 0.007491f
C801 B.n603 VSUBS 0.007491f
C802 B.n604 VSUBS 0.007491f
C803 B.n605 VSUBS 0.007491f
C804 B.n606 VSUBS 0.007491f
C805 B.n607 VSUBS 0.007491f
C806 B.n608 VSUBS 0.007491f
C807 B.n609 VSUBS 0.007491f
C808 B.n610 VSUBS 0.007491f
C809 B.n611 VSUBS 0.007491f
C810 B.n612 VSUBS 0.007491f
C811 B.n613 VSUBS 0.007491f
C812 B.n614 VSUBS 0.007491f
C813 B.n615 VSUBS 0.007491f
C814 B.n616 VSUBS 0.007491f
C815 B.n617 VSUBS 0.01851f
C816 B.n618 VSUBS 0.017624f
C817 B.n619 VSUBS 0.017624f
C818 B.n620 VSUBS 0.007491f
C819 B.n621 VSUBS 0.007491f
C820 B.n622 VSUBS 0.007491f
C821 B.n623 VSUBS 0.007491f
C822 B.n624 VSUBS 0.007491f
C823 B.n625 VSUBS 0.007491f
C824 B.n626 VSUBS 0.007491f
C825 B.n627 VSUBS 0.007491f
C826 B.n628 VSUBS 0.007491f
C827 B.n629 VSUBS 0.007491f
C828 B.n630 VSUBS 0.007491f
C829 B.n631 VSUBS 0.007491f
C830 B.n632 VSUBS 0.007491f
C831 B.n633 VSUBS 0.007491f
C832 B.n634 VSUBS 0.007491f
C833 B.n635 VSUBS 0.007491f
C834 B.n636 VSUBS 0.007491f
C835 B.n637 VSUBS 0.007491f
C836 B.n638 VSUBS 0.007491f
C837 B.n639 VSUBS 0.007491f
C838 B.n640 VSUBS 0.007491f
C839 B.n641 VSUBS 0.007491f
C840 B.n642 VSUBS 0.007491f
C841 B.n643 VSUBS 0.007491f
C842 B.n644 VSUBS 0.007491f
C843 B.n645 VSUBS 0.007491f
C844 B.n646 VSUBS 0.007491f
C845 B.n647 VSUBS 0.007491f
C846 B.n648 VSUBS 0.007491f
C847 B.n649 VSUBS 0.007491f
C848 B.n650 VSUBS 0.007491f
C849 B.n651 VSUBS 0.007491f
C850 B.n652 VSUBS 0.007491f
C851 B.n653 VSUBS 0.007491f
C852 B.n654 VSUBS 0.007491f
C853 B.n655 VSUBS 0.007491f
C854 B.n656 VSUBS 0.007491f
C855 B.n657 VSUBS 0.007491f
C856 B.n658 VSUBS 0.007491f
C857 B.n659 VSUBS 0.007491f
C858 B.n660 VSUBS 0.007491f
C859 B.n661 VSUBS 0.007491f
C860 B.n662 VSUBS 0.007491f
C861 B.n663 VSUBS 0.007491f
C862 B.n664 VSUBS 0.007491f
C863 B.n665 VSUBS 0.007491f
C864 B.n666 VSUBS 0.007491f
C865 B.n667 VSUBS 0.007491f
C866 B.n668 VSUBS 0.007491f
C867 B.n669 VSUBS 0.007491f
C868 B.n670 VSUBS 0.007491f
C869 B.n671 VSUBS 0.007491f
C870 B.n672 VSUBS 0.007491f
C871 B.n673 VSUBS 0.007491f
C872 B.n674 VSUBS 0.007491f
C873 B.n675 VSUBS 0.007491f
C874 B.n676 VSUBS 0.007491f
C875 B.n677 VSUBS 0.007491f
C876 B.n678 VSUBS 0.007491f
C877 B.n679 VSUBS 0.016963f
C878 VDD1.n0 VSUBS 0.02873f
C879 VDD1.n1 VSUBS 0.025268f
C880 VDD1.n2 VSUBS 0.013578f
C881 VDD1.n3 VSUBS 0.032093f
C882 VDD1.n4 VSUBS 0.014377f
C883 VDD1.n5 VSUBS 0.025268f
C884 VDD1.n6 VSUBS 0.013578f
C885 VDD1.n7 VSUBS 0.032093f
C886 VDD1.n8 VSUBS 0.014377f
C887 VDD1.n9 VSUBS 0.025268f
C888 VDD1.n10 VSUBS 0.013578f
C889 VDD1.n11 VSUBS 0.032093f
C890 VDD1.n12 VSUBS 0.032093f
C891 VDD1.n13 VSUBS 0.014377f
C892 VDD1.n14 VSUBS 0.025268f
C893 VDD1.n15 VSUBS 0.013578f
C894 VDD1.n16 VSUBS 0.032093f
C895 VDD1.n17 VSUBS 0.014377f
C896 VDD1.n18 VSUBS 0.185988f
C897 VDD1.t5 VSUBS 0.069074f
C898 VDD1.n19 VSUBS 0.02407f
C899 VDD1.n20 VSUBS 0.024142f
C900 VDD1.n21 VSUBS 0.013578f
C901 VDD1.n22 VSUBS 1.11525f
C902 VDD1.n23 VSUBS 0.025268f
C903 VDD1.n24 VSUBS 0.013578f
C904 VDD1.n25 VSUBS 0.014377f
C905 VDD1.n26 VSUBS 0.032093f
C906 VDD1.n27 VSUBS 0.032093f
C907 VDD1.n28 VSUBS 0.014377f
C908 VDD1.n29 VSUBS 0.013578f
C909 VDD1.n30 VSUBS 0.025268f
C910 VDD1.n31 VSUBS 0.025268f
C911 VDD1.n32 VSUBS 0.013578f
C912 VDD1.n33 VSUBS 0.014377f
C913 VDD1.n34 VSUBS 0.032093f
C914 VDD1.n35 VSUBS 0.032093f
C915 VDD1.n36 VSUBS 0.014377f
C916 VDD1.n37 VSUBS 0.013578f
C917 VDD1.n38 VSUBS 0.025268f
C918 VDD1.n39 VSUBS 0.025268f
C919 VDD1.n40 VSUBS 0.013578f
C920 VDD1.n41 VSUBS 0.013977f
C921 VDD1.n42 VSUBS 0.013977f
C922 VDD1.n43 VSUBS 0.032093f
C923 VDD1.n44 VSUBS 0.032093f
C924 VDD1.n45 VSUBS 0.014377f
C925 VDD1.n46 VSUBS 0.013578f
C926 VDD1.n47 VSUBS 0.025268f
C927 VDD1.n48 VSUBS 0.025268f
C928 VDD1.n49 VSUBS 0.013578f
C929 VDD1.n50 VSUBS 0.014377f
C930 VDD1.n51 VSUBS 0.032093f
C931 VDD1.n52 VSUBS 0.080983f
C932 VDD1.n53 VSUBS 0.014377f
C933 VDD1.n54 VSUBS 0.013578f
C934 VDD1.n55 VSUBS 0.064619f
C935 VDD1.n56 VSUBS 0.06517f
C936 VDD1.n57 VSUBS 0.02873f
C937 VDD1.n58 VSUBS 0.025268f
C938 VDD1.n59 VSUBS 0.013578f
C939 VDD1.n60 VSUBS 0.032093f
C940 VDD1.n61 VSUBS 0.014377f
C941 VDD1.n62 VSUBS 0.025268f
C942 VDD1.n63 VSUBS 0.013578f
C943 VDD1.n64 VSUBS 0.032093f
C944 VDD1.n65 VSUBS 0.014377f
C945 VDD1.n66 VSUBS 0.025268f
C946 VDD1.n67 VSUBS 0.013578f
C947 VDD1.n68 VSUBS 0.032093f
C948 VDD1.n69 VSUBS 0.014377f
C949 VDD1.n70 VSUBS 0.025268f
C950 VDD1.n71 VSUBS 0.013578f
C951 VDD1.n72 VSUBS 0.032093f
C952 VDD1.n73 VSUBS 0.014377f
C953 VDD1.n74 VSUBS 0.185988f
C954 VDD1.t1 VSUBS 0.069074f
C955 VDD1.n75 VSUBS 0.02407f
C956 VDD1.n76 VSUBS 0.024142f
C957 VDD1.n77 VSUBS 0.013578f
C958 VDD1.n78 VSUBS 1.11525f
C959 VDD1.n79 VSUBS 0.025268f
C960 VDD1.n80 VSUBS 0.013578f
C961 VDD1.n81 VSUBS 0.014377f
C962 VDD1.n82 VSUBS 0.032093f
C963 VDD1.n83 VSUBS 0.032093f
C964 VDD1.n84 VSUBS 0.014377f
C965 VDD1.n85 VSUBS 0.013578f
C966 VDD1.n86 VSUBS 0.025268f
C967 VDD1.n87 VSUBS 0.025268f
C968 VDD1.n88 VSUBS 0.013578f
C969 VDD1.n89 VSUBS 0.014377f
C970 VDD1.n90 VSUBS 0.032093f
C971 VDD1.n91 VSUBS 0.032093f
C972 VDD1.n92 VSUBS 0.032093f
C973 VDD1.n93 VSUBS 0.014377f
C974 VDD1.n94 VSUBS 0.013578f
C975 VDD1.n95 VSUBS 0.025268f
C976 VDD1.n96 VSUBS 0.025268f
C977 VDD1.n97 VSUBS 0.013578f
C978 VDD1.n98 VSUBS 0.013977f
C979 VDD1.n99 VSUBS 0.013977f
C980 VDD1.n100 VSUBS 0.032093f
C981 VDD1.n101 VSUBS 0.032093f
C982 VDD1.n102 VSUBS 0.014377f
C983 VDD1.n103 VSUBS 0.013578f
C984 VDD1.n104 VSUBS 0.025268f
C985 VDD1.n105 VSUBS 0.025268f
C986 VDD1.n106 VSUBS 0.013578f
C987 VDD1.n107 VSUBS 0.014377f
C988 VDD1.n108 VSUBS 0.032093f
C989 VDD1.n109 VSUBS 0.080983f
C990 VDD1.n110 VSUBS 0.014377f
C991 VDD1.n111 VSUBS 0.013578f
C992 VDD1.n112 VSUBS 0.064619f
C993 VDD1.n113 VSUBS 0.064483f
C994 VDD1.t3 VSUBS 0.216847f
C995 VDD1.t0 VSUBS 0.216847f
C996 VDD1.n114 VSUBS 1.67777f
C997 VDD1.n115 VSUBS 2.91282f
C998 VDD1.t4 VSUBS 0.216847f
C999 VDD1.t2 VSUBS 0.216847f
C1000 VDD1.n116 VSUBS 1.67312f
C1001 VDD1.n117 VSUBS 2.91786f
C1002 VTAIL.t0 VSUBS 0.252819f
C1003 VTAIL.t11 VSUBS 0.252819f
C1004 VTAIL.n0 VSUBS 1.81115f
C1005 VTAIL.n1 VSUBS 0.846441f
C1006 VTAIL.n2 VSUBS 0.033495f
C1007 VTAIL.n3 VSUBS 0.029459f
C1008 VTAIL.n4 VSUBS 0.01583f
C1009 VTAIL.n5 VSUBS 0.037417f
C1010 VTAIL.n6 VSUBS 0.016762f
C1011 VTAIL.n7 VSUBS 0.029459f
C1012 VTAIL.n8 VSUBS 0.01583f
C1013 VTAIL.n9 VSUBS 0.037417f
C1014 VTAIL.n10 VSUBS 0.016762f
C1015 VTAIL.n11 VSUBS 0.029459f
C1016 VTAIL.n12 VSUBS 0.01583f
C1017 VTAIL.n13 VSUBS 0.037417f
C1018 VTAIL.n14 VSUBS 0.016762f
C1019 VTAIL.n15 VSUBS 0.029459f
C1020 VTAIL.n16 VSUBS 0.01583f
C1021 VTAIL.n17 VSUBS 0.037417f
C1022 VTAIL.n18 VSUBS 0.016762f
C1023 VTAIL.n19 VSUBS 0.21684f
C1024 VTAIL.t6 VSUBS 0.080533f
C1025 VTAIL.n20 VSUBS 0.028063f
C1026 VTAIL.n21 VSUBS 0.028147f
C1027 VTAIL.n22 VSUBS 0.01583f
C1028 VTAIL.n23 VSUBS 1.30026f
C1029 VTAIL.n24 VSUBS 0.029459f
C1030 VTAIL.n25 VSUBS 0.01583f
C1031 VTAIL.n26 VSUBS 0.016762f
C1032 VTAIL.n27 VSUBS 0.037417f
C1033 VTAIL.n28 VSUBS 0.037417f
C1034 VTAIL.n29 VSUBS 0.016762f
C1035 VTAIL.n30 VSUBS 0.01583f
C1036 VTAIL.n31 VSUBS 0.029459f
C1037 VTAIL.n32 VSUBS 0.029459f
C1038 VTAIL.n33 VSUBS 0.01583f
C1039 VTAIL.n34 VSUBS 0.016762f
C1040 VTAIL.n35 VSUBS 0.037417f
C1041 VTAIL.n36 VSUBS 0.037417f
C1042 VTAIL.n37 VSUBS 0.037417f
C1043 VTAIL.n38 VSUBS 0.016762f
C1044 VTAIL.n39 VSUBS 0.01583f
C1045 VTAIL.n40 VSUBS 0.029459f
C1046 VTAIL.n41 VSUBS 0.029459f
C1047 VTAIL.n42 VSUBS 0.01583f
C1048 VTAIL.n43 VSUBS 0.016296f
C1049 VTAIL.n44 VSUBS 0.016296f
C1050 VTAIL.n45 VSUBS 0.037417f
C1051 VTAIL.n46 VSUBS 0.037417f
C1052 VTAIL.n47 VSUBS 0.016762f
C1053 VTAIL.n48 VSUBS 0.01583f
C1054 VTAIL.n49 VSUBS 0.029459f
C1055 VTAIL.n50 VSUBS 0.029459f
C1056 VTAIL.n51 VSUBS 0.01583f
C1057 VTAIL.n52 VSUBS 0.016762f
C1058 VTAIL.n53 VSUBS 0.037417f
C1059 VTAIL.n54 VSUBS 0.094417f
C1060 VTAIL.n55 VSUBS 0.016762f
C1061 VTAIL.n56 VSUBS 0.01583f
C1062 VTAIL.n57 VSUBS 0.075338f
C1063 VTAIL.n58 VSUBS 0.047864f
C1064 VTAIL.n59 VSUBS 0.407732f
C1065 VTAIL.t7 VSUBS 0.252819f
C1066 VTAIL.t9 VSUBS 0.252819f
C1067 VTAIL.n60 VSUBS 1.81115f
C1068 VTAIL.n61 VSUBS 2.586f
C1069 VTAIL.t4 VSUBS 0.252819f
C1070 VTAIL.t1 VSUBS 0.252819f
C1071 VTAIL.n62 VSUBS 1.81116f
C1072 VTAIL.n63 VSUBS 2.58599f
C1073 VTAIL.n64 VSUBS 0.033495f
C1074 VTAIL.n65 VSUBS 0.029459f
C1075 VTAIL.n66 VSUBS 0.01583f
C1076 VTAIL.n67 VSUBS 0.037417f
C1077 VTAIL.n68 VSUBS 0.016762f
C1078 VTAIL.n69 VSUBS 0.029459f
C1079 VTAIL.n70 VSUBS 0.01583f
C1080 VTAIL.n71 VSUBS 0.037417f
C1081 VTAIL.n72 VSUBS 0.016762f
C1082 VTAIL.n73 VSUBS 0.029459f
C1083 VTAIL.n74 VSUBS 0.01583f
C1084 VTAIL.n75 VSUBS 0.037417f
C1085 VTAIL.n76 VSUBS 0.037417f
C1086 VTAIL.n77 VSUBS 0.016762f
C1087 VTAIL.n78 VSUBS 0.029459f
C1088 VTAIL.n79 VSUBS 0.01583f
C1089 VTAIL.n80 VSUBS 0.037417f
C1090 VTAIL.n81 VSUBS 0.016762f
C1091 VTAIL.n82 VSUBS 0.21684f
C1092 VTAIL.t2 VSUBS 0.080533f
C1093 VTAIL.n83 VSUBS 0.028063f
C1094 VTAIL.n84 VSUBS 0.028147f
C1095 VTAIL.n85 VSUBS 0.01583f
C1096 VTAIL.n86 VSUBS 1.30026f
C1097 VTAIL.n87 VSUBS 0.029459f
C1098 VTAIL.n88 VSUBS 0.01583f
C1099 VTAIL.n89 VSUBS 0.016762f
C1100 VTAIL.n90 VSUBS 0.037417f
C1101 VTAIL.n91 VSUBS 0.037417f
C1102 VTAIL.n92 VSUBS 0.016762f
C1103 VTAIL.n93 VSUBS 0.01583f
C1104 VTAIL.n94 VSUBS 0.029459f
C1105 VTAIL.n95 VSUBS 0.029459f
C1106 VTAIL.n96 VSUBS 0.01583f
C1107 VTAIL.n97 VSUBS 0.016762f
C1108 VTAIL.n98 VSUBS 0.037417f
C1109 VTAIL.n99 VSUBS 0.037417f
C1110 VTAIL.n100 VSUBS 0.016762f
C1111 VTAIL.n101 VSUBS 0.01583f
C1112 VTAIL.n102 VSUBS 0.029459f
C1113 VTAIL.n103 VSUBS 0.029459f
C1114 VTAIL.n104 VSUBS 0.01583f
C1115 VTAIL.n105 VSUBS 0.016296f
C1116 VTAIL.n106 VSUBS 0.016296f
C1117 VTAIL.n107 VSUBS 0.037417f
C1118 VTAIL.n108 VSUBS 0.037417f
C1119 VTAIL.n109 VSUBS 0.016762f
C1120 VTAIL.n110 VSUBS 0.01583f
C1121 VTAIL.n111 VSUBS 0.029459f
C1122 VTAIL.n112 VSUBS 0.029459f
C1123 VTAIL.n113 VSUBS 0.01583f
C1124 VTAIL.n114 VSUBS 0.016762f
C1125 VTAIL.n115 VSUBS 0.037417f
C1126 VTAIL.n116 VSUBS 0.094417f
C1127 VTAIL.n117 VSUBS 0.016762f
C1128 VTAIL.n118 VSUBS 0.01583f
C1129 VTAIL.n119 VSUBS 0.075338f
C1130 VTAIL.n120 VSUBS 0.047864f
C1131 VTAIL.n121 VSUBS 0.407732f
C1132 VTAIL.t5 VSUBS 0.252819f
C1133 VTAIL.t10 VSUBS 0.252819f
C1134 VTAIL.n122 VSUBS 1.81116f
C1135 VTAIL.n123 VSUBS 1.00784f
C1136 VTAIL.n124 VSUBS 0.033495f
C1137 VTAIL.n125 VSUBS 0.029459f
C1138 VTAIL.n126 VSUBS 0.01583f
C1139 VTAIL.n127 VSUBS 0.037417f
C1140 VTAIL.n128 VSUBS 0.016762f
C1141 VTAIL.n129 VSUBS 0.029459f
C1142 VTAIL.n130 VSUBS 0.01583f
C1143 VTAIL.n131 VSUBS 0.037417f
C1144 VTAIL.n132 VSUBS 0.016762f
C1145 VTAIL.n133 VSUBS 0.029459f
C1146 VTAIL.n134 VSUBS 0.01583f
C1147 VTAIL.n135 VSUBS 0.037417f
C1148 VTAIL.n136 VSUBS 0.037417f
C1149 VTAIL.n137 VSUBS 0.016762f
C1150 VTAIL.n138 VSUBS 0.029459f
C1151 VTAIL.n139 VSUBS 0.01583f
C1152 VTAIL.n140 VSUBS 0.037417f
C1153 VTAIL.n141 VSUBS 0.016762f
C1154 VTAIL.n142 VSUBS 0.21684f
C1155 VTAIL.t8 VSUBS 0.080533f
C1156 VTAIL.n143 VSUBS 0.028063f
C1157 VTAIL.n144 VSUBS 0.028147f
C1158 VTAIL.n145 VSUBS 0.01583f
C1159 VTAIL.n146 VSUBS 1.30026f
C1160 VTAIL.n147 VSUBS 0.029459f
C1161 VTAIL.n148 VSUBS 0.01583f
C1162 VTAIL.n149 VSUBS 0.016762f
C1163 VTAIL.n150 VSUBS 0.037417f
C1164 VTAIL.n151 VSUBS 0.037417f
C1165 VTAIL.n152 VSUBS 0.016762f
C1166 VTAIL.n153 VSUBS 0.01583f
C1167 VTAIL.n154 VSUBS 0.029459f
C1168 VTAIL.n155 VSUBS 0.029459f
C1169 VTAIL.n156 VSUBS 0.01583f
C1170 VTAIL.n157 VSUBS 0.016762f
C1171 VTAIL.n158 VSUBS 0.037417f
C1172 VTAIL.n159 VSUBS 0.037417f
C1173 VTAIL.n160 VSUBS 0.016762f
C1174 VTAIL.n161 VSUBS 0.01583f
C1175 VTAIL.n162 VSUBS 0.029459f
C1176 VTAIL.n163 VSUBS 0.029459f
C1177 VTAIL.n164 VSUBS 0.01583f
C1178 VTAIL.n165 VSUBS 0.016296f
C1179 VTAIL.n166 VSUBS 0.016296f
C1180 VTAIL.n167 VSUBS 0.037417f
C1181 VTAIL.n168 VSUBS 0.037417f
C1182 VTAIL.n169 VSUBS 0.016762f
C1183 VTAIL.n170 VSUBS 0.01583f
C1184 VTAIL.n171 VSUBS 0.029459f
C1185 VTAIL.n172 VSUBS 0.029459f
C1186 VTAIL.n173 VSUBS 0.01583f
C1187 VTAIL.n174 VSUBS 0.016762f
C1188 VTAIL.n175 VSUBS 0.037417f
C1189 VTAIL.n176 VSUBS 0.094417f
C1190 VTAIL.n177 VSUBS 0.016762f
C1191 VTAIL.n178 VSUBS 0.01583f
C1192 VTAIL.n179 VSUBS 0.075338f
C1193 VTAIL.n180 VSUBS 0.047864f
C1194 VTAIL.n181 VSUBS 1.76329f
C1195 VTAIL.n182 VSUBS 0.033495f
C1196 VTAIL.n183 VSUBS 0.029459f
C1197 VTAIL.n184 VSUBS 0.01583f
C1198 VTAIL.n185 VSUBS 0.037417f
C1199 VTAIL.n186 VSUBS 0.016762f
C1200 VTAIL.n187 VSUBS 0.029459f
C1201 VTAIL.n188 VSUBS 0.01583f
C1202 VTAIL.n189 VSUBS 0.037417f
C1203 VTAIL.n190 VSUBS 0.016762f
C1204 VTAIL.n191 VSUBS 0.029459f
C1205 VTAIL.n192 VSUBS 0.01583f
C1206 VTAIL.n193 VSUBS 0.037417f
C1207 VTAIL.n194 VSUBS 0.016762f
C1208 VTAIL.n195 VSUBS 0.029459f
C1209 VTAIL.n196 VSUBS 0.01583f
C1210 VTAIL.n197 VSUBS 0.037417f
C1211 VTAIL.n198 VSUBS 0.016762f
C1212 VTAIL.n199 VSUBS 0.21684f
C1213 VTAIL.t3 VSUBS 0.080533f
C1214 VTAIL.n200 VSUBS 0.028063f
C1215 VTAIL.n201 VSUBS 0.028147f
C1216 VTAIL.n202 VSUBS 0.01583f
C1217 VTAIL.n203 VSUBS 1.30026f
C1218 VTAIL.n204 VSUBS 0.029459f
C1219 VTAIL.n205 VSUBS 0.01583f
C1220 VTAIL.n206 VSUBS 0.016762f
C1221 VTAIL.n207 VSUBS 0.037417f
C1222 VTAIL.n208 VSUBS 0.037417f
C1223 VTAIL.n209 VSUBS 0.016762f
C1224 VTAIL.n210 VSUBS 0.01583f
C1225 VTAIL.n211 VSUBS 0.029459f
C1226 VTAIL.n212 VSUBS 0.029459f
C1227 VTAIL.n213 VSUBS 0.01583f
C1228 VTAIL.n214 VSUBS 0.016762f
C1229 VTAIL.n215 VSUBS 0.037417f
C1230 VTAIL.n216 VSUBS 0.037417f
C1231 VTAIL.n217 VSUBS 0.037417f
C1232 VTAIL.n218 VSUBS 0.016762f
C1233 VTAIL.n219 VSUBS 0.01583f
C1234 VTAIL.n220 VSUBS 0.029459f
C1235 VTAIL.n221 VSUBS 0.029459f
C1236 VTAIL.n222 VSUBS 0.01583f
C1237 VTAIL.n223 VSUBS 0.016296f
C1238 VTAIL.n224 VSUBS 0.016296f
C1239 VTAIL.n225 VSUBS 0.037417f
C1240 VTAIL.n226 VSUBS 0.037417f
C1241 VTAIL.n227 VSUBS 0.016762f
C1242 VTAIL.n228 VSUBS 0.01583f
C1243 VTAIL.n229 VSUBS 0.029459f
C1244 VTAIL.n230 VSUBS 0.029459f
C1245 VTAIL.n231 VSUBS 0.01583f
C1246 VTAIL.n232 VSUBS 0.016762f
C1247 VTAIL.n233 VSUBS 0.037417f
C1248 VTAIL.n234 VSUBS 0.094417f
C1249 VTAIL.n235 VSUBS 0.016762f
C1250 VTAIL.n236 VSUBS 0.01583f
C1251 VTAIL.n237 VSUBS 0.075338f
C1252 VTAIL.n238 VSUBS 0.047864f
C1253 VTAIL.n239 VSUBS 1.70212f
C1254 VP.n0 VSUBS 0.044431f
C1255 VP.t5 VSUBS 2.37623f
C1256 VP.n1 VSUBS 0.0367f
C1257 VP.n2 VSUBS 0.033702f
C1258 VP.t2 VSUBS 2.37623f
C1259 VP.n3 VSUBS 0.062498f
C1260 VP.n4 VSUBS 0.033702f
C1261 VP.n5 VSUBS 0.04522f
C1262 VP.n6 VSUBS 0.044431f
C1263 VP.t3 VSUBS 2.37623f
C1264 VP.n7 VSUBS 0.0367f
C1265 VP.n8 VSUBS 0.318599f
C1266 VP.t1 VSUBS 2.37623f
C1267 VP.t0 VSUBS 2.62383f
C1268 VP.n9 VSUBS 0.913507f
C1269 VP.n10 VSUBS 0.95812f
C1270 VP.n11 VSUBS 0.062498f
C1271 VP.n12 VSUBS 0.058793f
C1272 VP.n13 VSUBS 0.033702f
C1273 VP.n14 VSUBS 0.033702f
C1274 VP.n15 VSUBS 0.033702f
C1275 VP.n16 VSUBS 0.064987f
C1276 VP.n17 VSUBS 0.04522f
C1277 VP.n18 VSUBS 0.952209f
C1278 VP.n19 VSUBS 1.7046f
C1279 VP.t4 VSUBS 2.37623f
C1280 VP.n20 VSUBS 0.952209f
C1281 VP.n21 VSUBS 1.73047f
C1282 VP.n22 VSUBS 0.044431f
C1283 VP.n23 VSUBS 0.033702f
C1284 VP.n24 VSUBS 0.064987f
C1285 VP.n25 VSUBS 0.0367f
C1286 VP.n26 VSUBS 0.058793f
C1287 VP.n27 VSUBS 0.033702f
C1288 VP.n28 VSUBS 0.033702f
C1289 VP.n29 VSUBS 0.033702f
C1290 VP.n30 VSUBS 0.879656f
C1291 VP.n31 VSUBS 0.062498f
C1292 VP.n32 VSUBS 0.058793f
C1293 VP.n33 VSUBS 0.033702f
C1294 VP.n34 VSUBS 0.033702f
C1295 VP.n35 VSUBS 0.033702f
C1296 VP.n36 VSUBS 0.064987f
C1297 VP.n37 VSUBS 0.04522f
C1298 VP.n38 VSUBS 0.952209f
C1299 VP.n39 VSUBS 0.051993f
.ends

