* NGSPICE file created from diff_pair_sample_0274.ext - technology: sky130A

.subckt diff_pair_sample_0274 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VN.t0 VDD2.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=4.524 pd=23.98 as=1.914 ps=11.93 w=11.6 l=1.19
X1 B.t17 B.t15 B.t16 B.t9 sky130_fd_pr__nfet_01v8 ad=4.524 pd=23.98 as=0 ps=0 w=11.6 l=1.19
X2 VDD1.t3 VP.t0 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.914 pd=11.93 as=4.524 ps=23.98 w=11.6 l=1.19
X3 VDD1.t2 VP.t1 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.914 pd=11.93 as=4.524 ps=23.98 w=11.6 l=1.19
X4 B.t14 B.t12 B.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=4.524 pd=23.98 as=0 ps=0 w=11.6 l=1.19
X5 VTAIL.t6 VN.t1 VDD2.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=4.524 pd=23.98 as=1.914 ps=11.93 w=11.6 l=1.19
X6 VTAIL.t0 VP.t2 VDD1.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=4.524 pd=23.98 as=1.914 ps=11.93 w=11.6 l=1.19
X7 VDD2.t2 VN.t2 VTAIL.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=1.914 pd=11.93 as=4.524 ps=23.98 w=11.6 l=1.19
X8 VDD2.t0 VN.t3 VTAIL.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=1.914 pd=11.93 as=4.524 ps=23.98 w=11.6 l=1.19
X9 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=4.524 pd=23.98 as=0 ps=0 w=11.6 l=1.19
X10 VTAIL.t1 VP.t3 VDD1.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=4.524 pd=23.98 as=1.914 ps=11.93 w=11.6 l=1.19
X11 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=4.524 pd=23.98 as=0 ps=0 w=11.6 l=1.19
R0 VN.n0 VN.t0 270.916
R1 VN.n1 VN.t3 270.916
R2 VN.n0 VN.t2 270.697
R3 VN.n1 VN.t1 270.697
R4 VN VN.n1 60.4544
R5 VN VN.n0 18.5416
R6 VDD2.n2 VDD2.n0 102.855
R7 VDD2.n2 VDD2.n1 65.2087
R8 VDD2.n1 VDD2.t3 1.7074
R9 VDD2.n1 VDD2.t0 1.7074
R10 VDD2.n0 VDD2.t1 1.7074
R11 VDD2.n0 VDD2.t2 1.7074
R12 VDD2 VDD2.n2 0.0586897
R13 VTAIL.n5 VTAIL.t0 50.2379
R14 VTAIL.n4 VTAIL.t4 50.2379
R15 VTAIL.n3 VTAIL.t6 50.2379
R16 VTAIL.n7 VTAIL.t5 50.237
R17 VTAIL.n0 VTAIL.t7 50.237
R18 VTAIL.n1 VTAIL.t2 50.237
R19 VTAIL.n2 VTAIL.t1 50.237
R20 VTAIL.n6 VTAIL.t3 50.2368
R21 VTAIL.n7 VTAIL.n6 23.6772
R22 VTAIL.n3 VTAIL.n2 23.6772
R23 VTAIL.n4 VTAIL.n3 1.31084
R24 VTAIL.n6 VTAIL.n5 1.31084
R25 VTAIL.n2 VTAIL.n1 1.31084
R26 VTAIL VTAIL.n0 0.713862
R27 VTAIL VTAIL.n7 0.597483
R28 VTAIL.n5 VTAIL.n4 0.470328
R29 VTAIL.n1 VTAIL.n0 0.470328
R30 B.n634 B.n633 585
R31 B.n269 B.n86 585
R32 B.n268 B.n267 585
R33 B.n266 B.n265 585
R34 B.n264 B.n263 585
R35 B.n262 B.n261 585
R36 B.n260 B.n259 585
R37 B.n258 B.n257 585
R38 B.n256 B.n255 585
R39 B.n254 B.n253 585
R40 B.n252 B.n251 585
R41 B.n250 B.n249 585
R42 B.n248 B.n247 585
R43 B.n246 B.n245 585
R44 B.n244 B.n243 585
R45 B.n242 B.n241 585
R46 B.n240 B.n239 585
R47 B.n238 B.n237 585
R48 B.n236 B.n235 585
R49 B.n234 B.n233 585
R50 B.n232 B.n231 585
R51 B.n230 B.n229 585
R52 B.n228 B.n227 585
R53 B.n226 B.n225 585
R54 B.n224 B.n223 585
R55 B.n222 B.n221 585
R56 B.n220 B.n219 585
R57 B.n218 B.n217 585
R58 B.n216 B.n215 585
R59 B.n214 B.n213 585
R60 B.n212 B.n211 585
R61 B.n210 B.n209 585
R62 B.n208 B.n207 585
R63 B.n206 B.n205 585
R64 B.n204 B.n203 585
R65 B.n202 B.n201 585
R66 B.n200 B.n199 585
R67 B.n198 B.n197 585
R68 B.n196 B.n195 585
R69 B.n194 B.n193 585
R70 B.n192 B.n191 585
R71 B.n190 B.n189 585
R72 B.n188 B.n187 585
R73 B.n186 B.n185 585
R74 B.n184 B.n183 585
R75 B.n182 B.n181 585
R76 B.n180 B.n179 585
R77 B.n178 B.n177 585
R78 B.n176 B.n175 585
R79 B.n174 B.n173 585
R80 B.n172 B.n171 585
R81 B.n170 B.n169 585
R82 B.n168 B.n167 585
R83 B.n166 B.n165 585
R84 B.n164 B.n163 585
R85 B.n162 B.n161 585
R86 B.n160 B.n159 585
R87 B.n158 B.n157 585
R88 B.n156 B.n155 585
R89 B.n154 B.n153 585
R90 B.n152 B.n151 585
R91 B.n150 B.n149 585
R92 B.n148 B.n147 585
R93 B.n146 B.n145 585
R94 B.n144 B.n143 585
R95 B.n142 B.n141 585
R96 B.n140 B.n139 585
R97 B.n138 B.n137 585
R98 B.n136 B.n135 585
R99 B.n134 B.n133 585
R100 B.n132 B.n131 585
R101 B.n130 B.n129 585
R102 B.n128 B.n127 585
R103 B.n126 B.n125 585
R104 B.n124 B.n123 585
R105 B.n122 B.n121 585
R106 B.n120 B.n119 585
R107 B.n118 B.n117 585
R108 B.n116 B.n115 585
R109 B.n114 B.n113 585
R110 B.n112 B.n111 585
R111 B.n110 B.n109 585
R112 B.n108 B.n107 585
R113 B.n106 B.n105 585
R114 B.n104 B.n103 585
R115 B.n102 B.n101 585
R116 B.n100 B.n99 585
R117 B.n98 B.n97 585
R118 B.n96 B.n95 585
R119 B.n94 B.n93 585
R120 B.n632 B.n41 585
R121 B.n637 B.n41 585
R122 B.n631 B.n40 585
R123 B.n638 B.n40 585
R124 B.n630 B.n629 585
R125 B.n629 B.n36 585
R126 B.n628 B.n35 585
R127 B.n644 B.n35 585
R128 B.n627 B.n34 585
R129 B.n645 B.n34 585
R130 B.n626 B.n33 585
R131 B.n646 B.n33 585
R132 B.n625 B.n624 585
R133 B.n624 B.n29 585
R134 B.n623 B.n28 585
R135 B.n652 B.n28 585
R136 B.n622 B.n27 585
R137 B.n653 B.n27 585
R138 B.n621 B.n26 585
R139 B.n654 B.n26 585
R140 B.n620 B.n619 585
R141 B.n619 B.n22 585
R142 B.n618 B.n21 585
R143 B.n660 B.n21 585
R144 B.n617 B.n20 585
R145 B.n661 B.n20 585
R146 B.n616 B.n19 585
R147 B.n662 B.n19 585
R148 B.n615 B.n614 585
R149 B.n614 B.n15 585
R150 B.n613 B.n14 585
R151 B.n668 B.n14 585
R152 B.n612 B.n13 585
R153 B.n669 B.n13 585
R154 B.n611 B.n12 585
R155 B.n670 B.n12 585
R156 B.n610 B.n609 585
R157 B.n609 B.n608 585
R158 B.n607 B.n606 585
R159 B.n607 B.n8 585
R160 B.n605 B.n7 585
R161 B.n677 B.n7 585
R162 B.n604 B.n6 585
R163 B.n678 B.n6 585
R164 B.n603 B.n5 585
R165 B.n679 B.n5 585
R166 B.n602 B.n601 585
R167 B.n601 B.n4 585
R168 B.n600 B.n270 585
R169 B.n600 B.n599 585
R170 B.n590 B.n271 585
R171 B.n272 B.n271 585
R172 B.n592 B.n591 585
R173 B.n593 B.n592 585
R174 B.n589 B.n277 585
R175 B.n277 B.n276 585
R176 B.n588 B.n587 585
R177 B.n587 B.n586 585
R178 B.n279 B.n278 585
R179 B.n280 B.n279 585
R180 B.n579 B.n578 585
R181 B.n580 B.n579 585
R182 B.n577 B.n285 585
R183 B.n285 B.n284 585
R184 B.n576 B.n575 585
R185 B.n575 B.n574 585
R186 B.n287 B.n286 585
R187 B.n288 B.n287 585
R188 B.n567 B.n566 585
R189 B.n568 B.n567 585
R190 B.n565 B.n293 585
R191 B.n293 B.n292 585
R192 B.n564 B.n563 585
R193 B.n563 B.n562 585
R194 B.n295 B.n294 585
R195 B.n296 B.n295 585
R196 B.n555 B.n554 585
R197 B.n556 B.n555 585
R198 B.n553 B.n301 585
R199 B.n301 B.n300 585
R200 B.n552 B.n551 585
R201 B.n551 B.n550 585
R202 B.n303 B.n302 585
R203 B.n304 B.n303 585
R204 B.n543 B.n542 585
R205 B.n544 B.n543 585
R206 B.n541 B.n309 585
R207 B.n309 B.n308 585
R208 B.n536 B.n535 585
R209 B.n534 B.n356 585
R210 B.n533 B.n355 585
R211 B.n538 B.n355 585
R212 B.n532 B.n531 585
R213 B.n530 B.n529 585
R214 B.n528 B.n527 585
R215 B.n526 B.n525 585
R216 B.n524 B.n523 585
R217 B.n522 B.n521 585
R218 B.n520 B.n519 585
R219 B.n518 B.n517 585
R220 B.n516 B.n515 585
R221 B.n514 B.n513 585
R222 B.n512 B.n511 585
R223 B.n510 B.n509 585
R224 B.n508 B.n507 585
R225 B.n506 B.n505 585
R226 B.n504 B.n503 585
R227 B.n502 B.n501 585
R228 B.n500 B.n499 585
R229 B.n498 B.n497 585
R230 B.n496 B.n495 585
R231 B.n494 B.n493 585
R232 B.n492 B.n491 585
R233 B.n490 B.n489 585
R234 B.n488 B.n487 585
R235 B.n486 B.n485 585
R236 B.n484 B.n483 585
R237 B.n482 B.n481 585
R238 B.n480 B.n479 585
R239 B.n478 B.n477 585
R240 B.n476 B.n475 585
R241 B.n474 B.n473 585
R242 B.n472 B.n471 585
R243 B.n470 B.n469 585
R244 B.n468 B.n467 585
R245 B.n466 B.n465 585
R246 B.n464 B.n463 585
R247 B.n462 B.n461 585
R248 B.n460 B.n459 585
R249 B.n457 B.n456 585
R250 B.n455 B.n454 585
R251 B.n453 B.n452 585
R252 B.n451 B.n450 585
R253 B.n449 B.n448 585
R254 B.n447 B.n446 585
R255 B.n445 B.n444 585
R256 B.n443 B.n442 585
R257 B.n441 B.n440 585
R258 B.n439 B.n438 585
R259 B.n436 B.n435 585
R260 B.n434 B.n433 585
R261 B.n432 B.n431 585
R262 B.n430 B.n429 585
R263 B.n428 B.n427 585
R264 B.n426 B.n425 585
R265 B.n424 B.n423 585
R266 B.n422 B.n421 585
R267 B.n420 B.n419 585
R268 B.n418 B.n417 585
R269 B.n416 B.n415 585
R270 B.n414 B.n413 585
R271 B.n412 B.n411 585
R272 B.n410 B.n409 585
R273 B.n408 B.n407 585
R274 B.n406 B.n405 585
R275 B.n404 B.n403 585
R276 B.n402 B.n401 585
R277 B.n400 B.n399 585
R278 B.n398 B.n397 585
R279 B.n396 B.n395 585
R280 B.n394 B.n393 585
R281 B.n392 B.n391 585
R282 B.n390 B.n389 585
R283 B.n388 B.n387 585
R284 B.n386 B.n385 585
R285 B.n384 B.n383 585
R286 B.n382 B.n381 585
R287 B.n380 B.n379 585
R288 B.n378 B.n377 585
R289 B.n376 B.n375 585
R290 B.n374 B.n373 585
R291 B.n372 B.n371 585
R292 B.n370 B.n369 585
R293 B.n368 B.n367 585
R294 B.n366 B.n365 585
R295 B.n364 B.n363 585
R296 B.n362 B.n361 585
R297 B.n311 B.n310 585
R298 B.n540 B.n539 585
R299 B.n539 B.n538 585
R300 B.n307 B.n306 585
R301 B.n308 B.n307 585
R302 B.n546 B.n545 585
R303 B.n545 B.n544 585
R304 B.n547 B.n305 585
R305 B.n305 B.n304 585
R306 B.n549 B.n548 585
R307 B.n550 B.n549 585
R308 B.n299 B.n298 585
R309 B.n300 B.n299 585
R310 B.n558 B.n557 585
R311 B.n557 B.n556 585
R312 B.n559 B.n297 585
R313 B.n297 B.n296 585
R314 B.n561 B.n560 585
R315 B.n562 B.n561 585
R316 B.n291 B.n290 585
R317 B.n292 B.n291 585
R318 B.n570 B.n569 585
R319 B.n569 B.n568 585
R320 B.n571 B.n289 585
R321 B.n289 B.n288 585
R322 B.n573 B.n572 585
R323 B.n574 B.n573 585
R324 B.n283 B.n282 585
R325 B.n284 B.n283 585
R326 B.n582 B.n581 585
R327 B.n581 B.n580 585
R328 B.n583 B.n281 585
R329 B.n281 B.n280 585
R330 B.n585 B.n584 585
R331 B.n586 B.n585 585
R332 B.n275 B.n274 585
R333 B.n276 B.n275 585
R334 B.n595 B.n594 585
R335 B.n594 B.n593 585
R336 B.n596 B.n273 585
R337 B.n273 B.n272 585
R338 B.n598 B.n597 585
R339 B.n599 B.n598 585
R340 B.n3 B.n0 585
R341 B.n4 B.n3 585
R342 B.n676 B.n1 585
R343 B.n677 B.n676 585
R344 B.n675 B.n674 585
R345 B.n675 B.n8 585
R346 B.n673 B.n9 585
R347 B.n608 B.n9 585
R348 B.n672 B.n671 585
R349 B.n671 B.n670 585
R350 B.n11 B.n10 585
R351 B.n669 B.n11 585
R352 B.n667 B.n666 585
R353 B.n668 B.n667 585
R354 B.n665 B.n16 585
R355 B.n16 B.n15 585
R356 B.n664 B.n663 585
R357 B.n663 B.n662 585
R358 B.n18 B.n17 585
R359 B.n661 B.n18 585
R360 B.n659 B.n658 585
R361 B.n660 B.n659 585
R362 B.n657 B.n23 585
R363 B.n23 B.n22 585
R364 B.n656 B.n655 585
R365 B.n655 B.n654 585
R366 B.n25 B.n24 585
R367 B.n653 B.n25 585
R368 B.n651 B.n650 585
R369 B.n652 B.n651 585
R370 B.n649 B.n30 585
R371 B.n30 B.n29 585
R372 B.n648 B.n647 585
R373 B.n647 B.n646 585
R374 B.n32 B.n31 585
R375 B.n645 B.n32 585
R376 B.n643 B.n642 585
R377 B.n644 B.n643 585
R378 B.n641 B.n37 585
R379 B.n37 B.n36 585
R380 B.n640 B.n639 585
R381 B.n639 B.n638 585
R382 B.n39 B.n38 585
R383 B.n637 B.n39 585
R384 B.n680 B.n679 585
R385 B.n678 B.n2 585
R386 B.n93 B.n39 540.549
R387 B.n634 B.n41 540.549
R388 B.n539 B.n309 540.549
R389 B.n536 B.n307 540.549
R390 B.n90 B.t4 438.99
R391 B.n87 B.t12 438.99
R392 B.n359 B.t15 438.99
R393 B.n357 B.t8 438.99
R394 B.n636 B.n635 256.663
R395 B.n636 B.n85 256.663
R396 B.n636 B.n84 256.663
R397 B.n636 B.n83 256.663
R398 B.n636 B.n82 256.663
R399 B.n636 B.n81 256.663
R400 B.n636 B.n80 256.663
R401 B.n636 B.n79 256.663
R402 B.n636 B.n78 256.663
R403 B.n636 B.n77 256.663
R404 B.n636 B.n76 256.663
R405 B.n636 B.n75 256.663
R406 B.n636 B.n74 256.663
R407 B.n636 B.n73 256.663
R408 B.n636 B.n72 256.663
R409 B.n636 B.n71 256.663
R410 B.n636 B.n70 256.663
R411 B.n636 B.n69 256.663
R412 B.n636 B.n68 256.663
R413 B.n636 B.n67 256.663
R414 B.n636 B.n66 256.663
R415 B.n636 B.n65 256.663
R416 B.n636 B.n64 256.663
R417 B.n636 B.n63 256.663
R418 B.n636 B.n62 256.663
R419 B.n636 B.n61 256.663
R420 B.n636 B.n60 256.663
R421 B.n636 B.n59 256.663
R422 B.n636 B.n58 256.663
R423 B.n636 B.n57 256.663
R424 B.n636 B.n56 256.663
R425 B.n636 B.n55 256.663
R426 B.n636 B.n54 256.663
R427 B.n636 B.n53 256.663
R428 B.n636 B.n52 256.663
R429 B.n636 B.n51 256.663
R430 B.n636 B.n50 256.663
R431 B.n636 B.n49 256.663
R432 B.n636 B.n48 256.663
R433 B.n636 B.n47 256.663
R434 B.n636 B.n46 256.663
R435 B.n636 B.n45 256.663
R436 B.n636 B.n44 256.663
R437 B.n636 B.n43 256.663
R438 B.n636 B.n42 256.663
R439 B.n538 B.n537 256.663
R440 B.n538 B.n312 256.663
R441 B.n538 B.n313 256.663
R442 B.n538 B.n314 256.663
R443 B.n538 B.n315 256.663
R444 B.n538 B.n316 256.663
R445 B.n538 B.n317 256.663
R446 B.n538 B.n318 256.663
R447 B.n538 B.n319 256.663
R448 B.n538 B.n320 256.663
R449 B.n538 B.n321 256.663
R450 B.n538 B.n322 256.663
R451 B.n538 B.n323 256.663
R452 B.n538 B.n324 256.663
R453 B.n538 B.n325 256.663
R454 B.n538 B.n326 256.663
R455 B.n538 B.n327 256.663
R456 B.n538 B.n328 256.663
R457 B.n538 B.n329 256.663
R458 B.n538 B.n330 256.663
R459 B.n538 B.n331 256.663
R460 B.n538 B.n332 256.663
R461 B.n538 B.n333 256.663
R462 B.n538 B.n334 256.663
R463 B.n538 B.n335 256.663
R464 B.n538 B.n336 256.663
R465 B.n538 B.n337 256.663
R466 B.n538 B.n338 256.663
R467 B.n538 B.n339 256.663
R468 B.n538 B.n340 256.663
R469 B.n538 B.n341 256.663
R470 B.n538 B.n342 256.663
R471 B.n538 B.n343 256.663
R472 B.n538 B.n344 256.663
R473 B.n538 B.n345 256.663
R474 B.n538 B.n346 256.663
R475 B.n538 B.n347 256.663
R476 B.n538 B.n348 256.663
R477 B.n538 B.n349 256.663
R478 B.n538 B.n350 256.663
R479 B.n538 B.n351 256.663
R480 B.n538 B.n352 256.663
R481 B.n538 B.n353 256.663
R482 B.n538 B.n354 256.663
R483 B.n682 B.n681 256.663
R484 B.n97 B.n96 163.367
R485 B.n101 B.n100 163.367
R486 B.n105 B.n104 163.367
R487 B.n109 B.n108 163.367
R488 B.n113 B.n112 163.367
R489 B.n117 B.n116 163.367
R490 B.n121 B.n120 163.367
R491 B.n125 B.n124 163.367
R492 B.n129 B.n128 163.367
R493 B.n133 B.n132 163.367
R494 B.n137 B.n136 163.367
R495 B.n141 B.n140 163.367
R496 B.n145 B.n144 163.367
R497 B.n149 B.n148 163.367
R498 B.n153 B.n152 163.367
R499 B.n157 B.n156 163.367
R500 B.n161 B.n160 163.367
R501 B.n165 B.n164 163.367
R502 B.n169 B.n168 163.367
R503 B.n173 B.n172 163.367
R504 B.n177 B.n176 163.367
R505 B.n181 B.n180 163.367
R506 B.n185 B.n184 163.367
R507 B.n189 B.n188 163.367
R508 B.n193 B.n192 163.367
R509 B.n197 B.n196 163.367
R510 B.n201 B.n200 163.367
R511 B.n205 B.n204 163.367
R512 B.n209 B.n208 163.367
R513 B.n213 B.n212 163.367
R514 B.n217 B.n216 163.367
R515 B.n221 B.n220 163.367
R516 B.n225 B.n224 163.367
R517 B.n229 B.n228 163.367
R518 B.n233 B.n232 163.367
R519 B.n237 B.n236 163.367
R520 B.n241 B.n240 163.367
R521 B.n245 B.n244 163.367
R522 B.n249 B.n248 163.367
R523 B.n253 B.n252 163.367
R524 B.n257 B.n256 163.367
R525 B.n261 B.n260 163.367
R526 B.n265 B.n264 163.367
R527 B.n267 B.n86 163.367
R528 B.n543 B.n309 163.367
R529 B.n543 B.n303 163.367
R530 B.n551 B.n303 163.367
R531 B.n551 B.n301 163.367
R532 B.n555 B.n301 163.367
R533 B.n555 B.n295 163.367
R534 B.n563 B.n295 163.367
R535 B.n563 B.n293 163.367
R536 B.n567 B.n293 163.367
R537 B.n567 B.n287 163.367
R538 B.n575 B.n287 163.367
R539 B.n575 B.n285 163.367
R540 B.n579 B.n285 163.367
R541 B.n579 B.n279 163.367
R542 B.n587 B.n279 163.367
R543 B.n587 B.n277 163.367
R544 B.n592 B.n277 163.367
R545 B.n592 B.n271 163.367
R546 B.n600 B.n271 163.367
R547 B.n601 B.n600 163.367
R548 B.n601 B.n5 163.367
R549 B.n6 B.n5 163.367
R550 B.n7 B.n6 163.367
R551 B.n607 B.n7 163.367
R552 B.n609 B.n607 163.367
R553 B.n609 B.n12 163.367
R554 B.n13 B.n12 163.367
R555 B.n14 B.n13 163.367
R556 B.n614 B.n14 163.367
R557 B.n614 B.n19 163.367
R558 B.n20 B.n19 163.367
R559 B.n21 B.n20 163.367
R560 B.n619 B.n21 163.367
R561 B.n619 B.n26 163.367
R562 B.n27 B.n26 163.367
R563 B.n28 B.n27 163.367
R564 B.n624 B.n28 163.367
R565 B.n624 B.n33 163.367
R566 B.n34 B.n33 163.367
R567 B.n35 B.n34 163.367
R568 B.n629 B.n35 163.367
R569 B.n629 B.n40 163.367
R570 B.n41 B.n40 163.367
R571 B.n356 B.n355 163.367
R572 B.n531 B.n355 163.367
R573 B.n529 B.n528 163.367
R574 B.n525 B.n524 163.367
R575 B.n521 B.n520 163.367
R576 B.n517 B.n516 163.367
R577 B.n513 B.n512 163.367
R578 B.n509 B.n508 163.367
R579 B.n505 B.n504 163.367
R580 B.n501 B.n500 163.367
R581 B.n497 B.n496 163.367
R582 B.n493 B.n492 163.367
R583 B.n489 B.n488 163.367
R584 B.n485 B.n484 163.367
R585 B.n481 B.n480 163.367
R586 B.n477 B.n476 163.367
R587 B.n473 B.n472 163.367
R588 B.n469 B.n468 163.367
R589 B.n465 B.n464 163.367
R590 B.n461 B.n460 163.367
R591 B.n456 B.n455 163.367
R592 B.n452 B.n451 163.367
R593 B.n448 B.n447 163.367
R594 B.n444 B.n443 163.367
R595 B.n440 B.n439 163.367
R596 B.n435 B.n434 163.367
R597 B.n431 B.n430 163.367
R598 B.n427 B.n426 163.367
R599 B.n423 B.n422 163.367
R600 B.n419 B.n418 163.367
R601 B.n415 B.n414 163.367
R602 B.n411 B.n410 163.367
R603 B.n407 B.n406 163.367
R604 B.n403 B.n402 163.367
R605 B.n399 B.n398 163.367
R606 B.n395 B.n394 163.367
R607 B.n391 B.n390 163.367
R608 B.n387 B.n386 163.367
R609 B.n383 B.n382 163.367
R610 B.n379 B.n378 163.367
R611 B.n375 B.n374 163.367
R612 B.n371 B.n370 163.367
R613 B.n367 B.n366 163.367
R614 B.n363 B.n362 163.367
R615 B.n539 B.n311 163.367
R616 B.n545 B.n307 163.367
R617 B.n545 B.n305 163.367
R618 B.n549 B.n305 163.367
R619 B.n549 B.n299 163.367
R620 B.n557 B.n299 163.367
R621 B.n557 B.n297 163.367
R622 B.n561 B.n297 163.367
R623 B.n561 B.n291 163.367
R624 B.n569 B.n291 163.367
R625 B.n569 B.n289 163.367
R626 B.n573 B.n289 163.367
R627 B.n573 B.n283 163.367
R628 B.n581 B.n283 163.367
R629 B.n581 B.n281 163.367
R630 B.n585 B.n281 163.367
R631 B.n585 B.n275 163.367
R632 B.n594 B.n275 163.367
R633 B.n594 B.n273 163.367
R634 B.n598 B.n273 163.367
R635 B.n598 B.n3 163.367
R636 B.n680 B.n3 163.367
R637 B.n676 B.n2 163.367
R638 B.n676 B.n675 163.367
R639 B.n675 B.n9 163.367
R640 B.n671 B.n9 163.367
R641 B.n671 B.n11 163.367
R642 B.n667 B.n11 163.367
R643 B.n667 B.n16 163.367
R644 B.n663 B.n16 163.367
R645 B.n663 B.n18 163.367
R646 B.n659 B.n18 163.367
R647 B.n659 B.n23 163.367
R648 B.n655 B.n23 163.367
R649 B.n655 B.n25 163.367
R650 B.n651 B.n25 163.367
R651 B.n651 B.n30 163.367
R652 B.n647 B.n30 163.367
R653 B.n647 B.n32 163.367
R654 B.n643 B.n32 163.367
R655 B.n643 B.n37 163.367
R656 B.n639 B.n37 163.367
R657 B.n639 B.n39 163.367
R658 B.n87 B.t13 98.1008
R659 B.n359 B.t17 98.1008
R660 B.n90 B.t6 98.0861
R661 B.n357 B.t11 98.0861
R662 B.n538 B.n308 81.482
R663 B.n637 B.n636 81.482
R664 B.n93 B.n42 71.676
R665 B.n97 B.n43 71.676
R666 B.n101 B.n44 71.676
R667 B.n105 B.n45 71.676
R668 B.n109 B.n46 71.676
R669 B.n113 B.n47 71.676
R670 B.n117 B.n48 71.676
R671 B.n121 B.n49 71.676
R672 B.n125 B.n50 71.676
R673 B.n129 B.n51 71.676
R674 B.n133 B.n52 71.676
R675 B.n137 B.n53 71.676
R676 B.n141 B.n54 71.676
R677 B.n145 B.n55 71.676
R678 B.n149 B.n56 71.676
R679 B.n153 B.n57 71.676
R680 B.n157 B.n58 71.676
R681 B.n161 B.n59 71.676
R682 B.n165 B.n60 71.676
R683 B.n169 B.n61 71.676
R684 B.n173 B.n62 71.676
R685 B.n177 B.n63 71.676
R686 B.n181 B.n64 71.676
R687 B.n185 B.n65 71.676
R688 B.n189 B.n66 71.676
R689 B.n193 B.n67 71.676
R690 B.n197 B.n68 71.676
R691 B.n201 B.n69 71.676
R692 B.n205 B.n70 71.676
R693 B.n209 B.n71 71.676
R694 B.n213 B.n72 71.676
R695 B.n217 B.n73 71.676
R696 B.n221 B.n74 71.676
R697 B.n225 B.n75 71.676
R698 B.n229 B.n76 71.676
R699 B.n233 B.n77 71.676
R700 B.n237 B.n78 71.676
R701 B.n241 B.n79 71.676
R702 B.n245 B.n80 71.676
R703 B.n249 B.n81 71.676
R704 B.n253 B.n82 71.676
R705 B.n257 B.n83 71.676
R706 B.n261 B.n84 71.676
R707 B.n265 B.n85 71.676
R708 B.n635 B.n86 71.676
R709 B.n635 B.n634 71.676
R710 B.n267 B.n85 71.676
R711 B.n264 B.n84 71.676
R712 B.n260 B.n83 71.676
R713 B.n256 B.n82 71.676
R714 B.n252 B.n81 71.676
R715 B.n248 B.n80 71.676
R716 B.n244 B.n79 71.676
R717 B.n240 B.n78 71.676
R718 B.n236 B.n77 71.676
R719 B.n232 B.n76 71.676
R720 B.n228 B.n75 71.676
R721 B.n224 B.n74 71.676
R722 B.n220 B.n73 71.676
R723 B.n216 B.n72 71.676
R724 B.n212 B.n71 71.676
R725 B.n208 B.n70 71.676
R726 B.n204 B.n69 71.676
R727 B.n200 B.n68 71.676
R728 B.n196 B.n67 71.676
R729 B.n192 B.n66 71.676
R730 B.n188 B.n65 71.676
R731 B.n184 B.n64 71.676
R732 B.n180 B.n63 71.676
R733 B.n176 B.n62 71.676
R734 B.n172 B.n61 71.676
R735 B.n168 B.n60 71.676
R736 B.n164 B.n59 71.676
R737 B.n160 B.n58 71.676
R738 B.n156 B.n57 71.676
R739 B.n152 B.n56 71.676
R740 B.n148 B.n55 71.676
R741 B.n144 B.n54 71.676
R742 B.n140 B.n53 71.676
R743 B.n136 B.n52 71.676
R744 B.n132 B.n51 71.676
R745 B.n128 B.n50 71.676
R746 B.n124 B.n49 71.676
R747 B.n120 B.n48 71.676
R748 B.n116 B.n47 71.676
R749 B.n112 B.n46 71.676
R750 B.n108 B.n45 71.676
R751 B.n104 B.n44 71.676
R752 B.n100 B.n43 71.676
R753 B.n96 B.n42 71.676
R754 B.n537 B.n536 71.676
R755 B.n531 B.n312 71.676
R756 B.n528 B.n313 71.676
R757 B.n524 B.n314 71.676
R758 B.n520 B.n315 71.676
R759 B.n516 B.n316 71.676
R760 B.n512 B.n317 71.676
R761 B.n508 B.n318 71.676
R762 B.n504 B.n319 71.676
R763 B.n500 B.n320 71.676
R764 B.n496 B.n321 71.676
R765 B.n492 B.n322 71.676
R766 B.n488 B.n323 71.676
R767 B.n484 B.n324 71.676
R768 B.n480 B.n325 71.676
R769 B.n476 B.n326 71.676
R770 B.n472 B.n327 71.676
R771 B.n468 B.n328 71.676
R772 B.n464 B.n329 71.676
R773 B.n460 B.n330 71.676
R774 B.n455 B.n331 71.676
R775 B.n451 B.n332 71.676
R776 B.n447 B.n333 71.676
R777 B.n443 B.n334 71.676
R778 B.n439 B.n335 71.676
R779 B.n434 B.n336 71.676
R780 B.n430 B.n337 71.676
R781 B.n426 B.n338 71.676
R782 B.n422 B.n339 71.676
R783 B.n418 B.n340 71.676
R784 B.n414 B.n341 71.676
R785 B.n410 B.n342 71.676
R786 B.n406 B.n343 71.676
R787 B.n402 B.n344 71.676
R788 B.n398 B.n345 71.676
R789 B.n394 B.n346 71.676
R790 B.n390 B.n347 71.676
R791 B.n386 B.n348 71.676
R792 B.n382 B.n349 71.676
R793 B.n378 B.n350 71.676
R794 B.n374 B.n351 71.676
R795 B.n370 B.n352 71.676
R796 B.n366 B.n353 71.676
R797 B.n362 B.n354 71.676
R798 B.n537 B.n356 71.676
R799 B.n529 B.n312 71.676
R800 B.n525 B.n313 71.676
R801 B.n521 B.n314 71.676
R802 B.n517 B.n315 71.676
R803 B.n513 B.n316 71.676
R804 B.n509 B.n317 71.676
R805 B.n505 B.n318 71.676
R806 B.n501 B.n319 71.676
R807 B.n497 B.n320 71.676
R808 B.n493 B.n321 71.676
R809 B.n489 B.n322 71.676
R810 B.n485 B.n323 71.676
R811 B.n481 B.n324 71.676
R812 B.n477 B.n325 71.676
R813 B.n473 B.n326 71.676
R814 B.n469 B.n327 71.676
R815 B.n465 B.n328 71.676
R816 B.n461 B.n329 71.676
R817 B.n456 B.n330 71.676
R818 B.n452 B.n331 71.676
R819 B.n448 B.n332 71.676
R820 B.n444 B.n333 71.676
R821 B.n440 B.n334 71.676
R822 B.n435 B.n335 71.676
R823 B.n431 B.n336 71.676
R824 B.n427 B.n337 71.676
R825 B.n423 B.n338 71.676
R826 B.n419 B.n339 71.676
R827 B.n415 B.n340 71.676
R828 B.n411 B.n341 71.676
R829 B.n407 B.n342 71.676
R830 B.n403 B.n343 71.676
R831 B.n399 B.n344 71.676
R832 B.n395 B.n345 71.676
R833 B.n391 B.n346 71.676
R834 B.n387 B.n347 71.676
R835 B.n383 B.n348 71.676
R836 B.n379 B.n349 71.676
R837 B.n375 B.n350 71.676
R838 B.n371 B.n351 71.676
R839 B.n367 B.n352 71.676
R840 B.n363 B.n353 71.676
R841 B.n354 B.n311 71.676
R842 B.n681 B.n680 71.676
R843 B.n681 B.n2 71.676
R844 B.n88 B.t14 68.6221
R845 B.n360 B.t16 68.6221
R846 B.n91 B.t7 68.6073
R847 B.n358 B.t10 68.6073
R848 B.n92 B.n91 59.5399
R849 B.n89 B.n88 59.5399
R850 B.n437 B.n360 59.5399
R851 B.n458 B.n358 59.5399
R852 B.n544 B.n308 44.3264
R853 B.n544 B.n304 44.3264
R854 B.n550 B.n304 44.3264
R855 B.n550 B.n300 44.3264
R856 B.n556 B.n300 44.3264
R857 B.n562 B.n296 44.3264
R858 B.n562 B.n292 44.3264
R859 B.n568 B.n292 44.3264
R860 B.n568 B.n288 44.3264
R861 B.n574 B.n288 44.3264
R862 B.n574 B.n284 44.3264
R863 B.n580 B.n284 44.3264
R864 B.n586 B.n280 44.3264
R865 B.n586 B.n276 44.3264
R866 B.n593 B.n276 44.3264
R867 B.n599 B.n272 44.3264
R868 B.n599 B.n4 44.3264
R869 B.n679 B.n4 44.3264
R870 B.n679 B.n678 44.3264
R871 B.n678 B.n677 44.3264
R872 B.n677 B.n8 44.3264
R873 B.n608 B.n8 44.3264
R874 B.n670 B.n669 44.3264
R875 B.n669 B.n668 44.3264
R876 B.n668 B.n15 44.3264
R877 B.n662 B.n661 44.3264
R878 B.n661 B.n660 44.3264
R879 B.n660 B.n22 44.3264
R880 B.n654 B.n22 44.3264
R881 B.n654 B.n653 44.3264
R882 B.n653 B.n652 44.3264
R883 B.n652 B.n29 44.3264
R884 B.n646 B.n645 44.3264
R885 B.n645 B.n644 44.3264
R886 B.n644 B.n36 44.3264
R887 B.n638 B.n36 44.3264
R888 B.n638 B.n637 44.3264
R889 B.t1 B.n280 35.8524
R890 B.t3 B.n15 35.8524
R891 B.n535 B.n306 35.1225
R892 B.n541 B.n540 35.1225
R893 B.n633 B.n632 35.1225
R894 B.n94 B.n38 35.1225
R895 B.n91 B.n90 29.4793
R896 B.n88 B.n87 29.4793
R897 B.n360 B.n359 29.4793
R898 B.n358 B.n357 29.4793
R899 B.n593 B.t2 29.3338
R900 B.n670 B.t0 29.3338
R901 B.n556 B.t9 22.8153
R902 B.n646 B.t5 22.8153
R903 B.t9 B.n296 21.5116
R904 B.t5 B.n29 21.5116
R905 B B.n682 18.0485
R906 B.t2 B.n272 14.9931
R907 B.n608 B.t0 14.9931
R908 B.n546 B.n306 10.6151
R909 B.n547 B.n546 10.6151
R910 B.n548 B.n547 10.6151
R911 B.n548 B.n298 10.6151
R912 B.n558 B.n298 10.6151
R913 B.n559 B.n558 10.6151
R914 B.n560 B.n559 10.6151
R915 B.n560 B.n290 10.6151
R916 B.n570 B.n290 10.6151
R917 B.n571 B.n570 10.6151
R918 B.n572 B.n571 10.6151
R919 B.n572 B.n282 10.6151
R920 B.n582 B.n282 10.6151
R921 B.n583 B.n582 10.6151
R922 B.n584 B.n583 10.6151
R923 B.n584 B.n274 10.6151
R924 B.n595 B.n274 10.6151
R925 B.n596 B.n595 10.6151
R926 B.n597 B.n596 10.6151
R927 B.n597 B.n0 10.6151
R928 B.n535 B.n534 10.6151
R929 B.n534 B.n533 10.6151
R930 B.n533 B.n532 10.6151
R931 B.n532 B.n530 10.6151
R932 B.n530 B.n527 10.6151
R933 B.n527 B.n526 10.6151
R934 B.n526 B.n523 10.6151
R935 B.n523 B.n522 10.6151
R936 B.n522 B.n519 10.6151
R937 B.n519 B.n518 10.6151
R938 B.n518 B.n515 10.6151
R939 B.n515 B.n514 10.6151
R940 B.n514 B.n511 10.6151
R941 B.n511 B.n510 10.6151
R942 B.n510 B.n507 10.6151
R943 B.n507 B.n506 10.6151
R944 B.n506 B.n503 10.6151
R945 B.n503 B.n502 10.6151
R946 B.n502 B.n499 10.6151
R947 B.n499 B.n498 10.6151
R948 B.n498 B.n495 10.6151
R949 B.n495 B.n494 10.6151
R950 B.n494 B.n491 10.6151
R951 B.n491 B.n490 10.6151
R952 B.n490 B.n487 10.6151
R953 B.n487 B.n486 10.6151
R954 B.n486 B.n483 10.6151
R955 B.n483 B.n482 10.6151
R956 B.n482 B.n479 10.6151
R957 B.n479 B.n478 10.6151
R958 B.n478 B.n475 10.6151
R959 B.n475 B.n474 10.6151
R960 B.n474 B.n471 10.6151
R961 B.n471 B.n470 10.6151
R962 B.n470 B.n467 10.6151
R963 B.n467 B.n466 10.6151
R964 B.n466 B.n463 10.6151
R965 B.n463 B.n462 10.6151
R966 B.n462 B.n459 10.6151
R967 B.n457 B.n454 10.6151
R968 B.n454 B.n453 10.6151
R969 B.n453 B.n450 10.6151
R970 B.n450 B.n449 10.6151
R971 B.n449 B.n446 10.6151
R972 B.n446 B.n445 10.6151
R973 B.n445 B.n442 10.6151
R974 B.n442 B.n441 10.6151
R975 B.n441 B.n438 10.6151
R976 B.n436 B.n433 10.6151
R977 B.n433 B.n432 10.6151
R978 B.n432 B.n429 10.6151
R979 B.n429 B.n428 10.6151
R980 B.n428 B.n425 10.6151
R981 B.n425 B.n424 10.6151
R982 B.n424 B.n421 10.6151
R983 B.n421 B.n420 10.6151
R984 B.n420 B.n417 10.6151
R985 B.n417 B.n416 10.6151
R986 B.n416 B.n413 10.6151
R987 B.n413 B.n412 10.6151
R988 B.n412 B.n409 10.6151
R989 B.n409 B.n408 10.6151
R990 B.n408 B.n405 10.6151
R991 B.n405 B.n404 10.6151
R992 B.n404 B.n401 10.6151
R993 B.n401 B.n400 10.6151
R994 B.n400 B.n397 10.6151
R995 B.n397 B.n396 10.6151
R996 B.n396 B.n393 10.6151
R997 B.n393 B.n392 10.6151
R998 B.n392 B.n389 10.6151
R999 B.n389 B.n388 10.6151
R1000 B.n388 B.n385 10.6151
R1001 B.n385 B.n384 10.6151
R1002 B.n384 B.n381 10.6151
R1003 B.n381 B.n380 10.6151
R1004 B.n380 B.n377 10.6151
R1005 B.n377 B.n376 10.6151
R1006 B.n376 B.n373 10.6151
R1007 B.n373 B.n372 10.6151
R1008 B.n372 B.n369 10.6151
R1009 B.n369 B.n368 10.6151
R1010 B.n368 B.n365 10.6151
R1011 B.n365 B.n364 10.6151
R1012 B.n364 B.n361 10.6151
R1013 B.n361 B.n310 10.6151
R1014 B.n540 B.n310 10.6151
R1015 B.n542 B.n541 10.6151
R1016 B.n542 B.n302 10.6151
R1017 B.n552 B.n302 10.6151
R1018 B.n553 B.n552 10.6151
R1019 B.n554 B.n553 10.6151
R1020 B.n554 B.n294 10.6151
R1021 B.n564 B.n294 10.6151
R1022 B.n565 B.n564 10.6151
R1023 B.n566 B.n565 10.6151
R1024 B.n566 B.n286 10.6151
R1025 B.n576 B.n286 10.6151
R1026 B.n577 B.n576 10.6151
R1027 B.n578 B.n577 10.6151
R1028 B.n578 B.n278 10.6151
R1029 B.n588 B.n278 10.6151
R1030 B.n589 B.n588 10.6151
R1031 B.n591 B.n589 10.6151
R1032 B.n591 B.n590 10.6151
R1033 B.n590 B.n270 10.6151
R1034 B.n602 B.n270 10.6151
R1035 B.n603 B.n602 10.6151
R1036 B.n604 B.n603 10.6151
R1037 B.n605 B.n604 10.6151
R1038 B.n606 B.n605 10.6151
R1039 B.n610 B.n606 10.6151
R1040 B.n611 B.n610 10.6151
R1041 B.n612 B.n611 10.6151
R1042 B.n613 B.n612 10.6151
R1043 B.n615 B.n613 10.6151
R1044 B.n616 B.n615 10.6151
R1045 B.n617 B.n616 10.6151
R1046 B.n618 B.n617 10.6151
R1047 B.n620 B.n618 10.6151
R1048 B.n621 B.n620 10.6151
R1049 B.n622 B.n621 10.6151
R1050 B.n623 B.n622 10.6151
R1051 B.n625 B.n623 10.6151
R1052 B.n626 B.n625 10.6151
R1053 B.n627 B.n626 10.6151
R1054 B.n628 B.n627 10.6151
R1055 B.n630 B.n628 10.6151
R1056 B.n631 B.n630 10.6151
R1057 B.n632 B.n631 10.6151
R1058 B.n674 B.n1 10.6151
R1059 B.n674 B.n673 10.6151
R1060 B.n673 B.n672 10.6151
R1061 B.n672 B.n10 10.6151
R1062 B.n666 B.n10 10.6151
R1063 B.n666 B.n665 10.6151
R1064 B.n665 B.n664 10.6151
R1065 B.n664 B.n17 10.6151
R1066 B.n658 B.n17 10.6151
R1067 B.n658 B.n657 10.6151
R1068 B.n657 B.n656 10.6151
R1069 B.n656 B.n24 10.6151
R1070 B.n650 B.n24 10.6151
R1071 B.n650 B.n649 10.6151
R1072 B.n649 B.n648 10.6151
R1073 B.n648 B.n31 10.6151
R1074 B.n642 B.n31 10.6151
R1075 B.n642 B.n641 10.6151
R1076 B.n641 B.n640 10.6151
R1077 B.n640 B.n38 10.6151
R1078 B.n95 B.n94 10.6151
R1079 B.n98 B.n95 10.6151
R1080 B.n99 B.n98 10.6151
R1081 B.n102 B.n99 10.6151
R1082 B.n103 B.n102 10.6151
R1083 B.n106 B.n103 10.6151
R1084 B.n107 B.n106 10.6151
R1085 B.n110 B.n107 10.6151
R1086 B.n111 B.n110 10.6151
R1087 B.n114 B.n111 10.6151
R1088 B.n115 B.n114 10.6151
R1089 B.n118 B.n115 10.6151
R1090 B.n119 B.n118 10.6151
R1091 B.n122 B.n119 10.6151
R1092 B.n123 B.n122 10.6151
R1093 B.n126 B.n123 10.6151
R1094 B.n127 B.n126 10.6151
R1095 B.n130 B.n127 10.6151
R1096 B.n131 B.n130 10.6151
R1097 B.n134 B.n131 10.6151
R1098 B.n135 B.n134 10.6151
R1099 B.n138 B.n135 10.6151
R1100 B.n139 B.n138 10.6151
R1101 B.n142 B.n139 10.6151
R1102 B.n143 B.n142 10.6151
R1103 B.n146 B.n143 10.6151
R1104 B.n147 B.n146 10.6151
R1105 B.n150 B.n147 10.6151
R1106 B.n151 B.n150 10.6151
R1107 B.n154 B.n151 10.6151
R1108 B.n155 B.n154 10.6151
R1109 B.n158 B.n155 10.6151
R1110 B.n159 B.n158 10.6151
R1111 B.n162 B.n159 10.6151
R1112 B.n163 B.n162 10.6151
R1113 B.n166 B.n163 10.6151
R1114 B.n167 B.n166 10.6151
R1115 B.n170 B.n167 10.6151
R1116 B.n171 B.n170 10.6151
R1117 B.n175 B.n174 10.6151
R1118 B.n178 B.n175 10.6151
R1119 B.n179 B.n178 10.6151
R1120 B.n182 B.n179 10.6151
R1121 B.n183 B.n182 10.6151
R1122 B.n186 B.n183 10.6151
R1123 B.n187 B.n186 10.6151
R1124 B.n190 B.n187 10.6151
R1125 B.n191 B.n190 10.6151
R1126 B.n195 B.n194 10.6151
R1127 B.n198 B.n195 10.6151
R1128 B.n199 B.n198 10.6151
R1129 B.n202 B.n199 10.6151
R1130 B.n203 B.n202 10.6151
R1131 B.n206 B.n203 10.6151
R1132 B.n207 B.n206 10.6151
R1133 B.n210 B.n207 10.6151
R1134 B.n211 B.n210 10.6151
R1135 B.n214 B.n211 10.6151
R1136 B.n215 B.n214 10.6151
R1137 B.n218 B.n215 10.6151
R1138 B.n219 B.n218 10.6151
R1139 B.n222 B.n219 10.6151
R1140 B.n223 B.n222 10.6151
R1141 B.n226 B.n223 10.6151
R1142 B.n227 B.n226 10.6151
R1143 B.n230 B.n227 10.6151
R1144 B.n231 B.n230 10.6151
R1145 B.n234 B.n231 10.6151
R1146 B.n235 B.n234 10.6151
R1147 B.n238 B.n235 10.6151
R1148 B.n239 B.n238 10.6151
R1149 B.n242 B.n239 10.6151
R1150 B.n243 B.n242 10.6151
R1151 B.n246 B.n243 10.6151
R1152 B.n247 B.n246 10.6151
R1153 B.n250 B.n247 10.6151
R1154 B.n251 B.n250 10.6151
R1155 B.n254 B.n251 10.6151
R1156 B.n255 B.n254 10.6151
R1157 B.n258 B.n255 10.6151
R1158 B.n259 B.n258 10.6151
R1159 B.n262 B.n259 10.6151
R1160 B.n263 B.n262 10.6151
R1161 B.n266 B.n263 10.6151
R1162 B.n268 B.n266 10.6151
R1163 B.n269 B.n268 10.6151
R1164 B.n633 B.n269 10.6151
R1165 B.n459 B.n458 9.36635
R1166 B.n437 B.n436 9.36635
R1167 B.n171 B.n92 9.36635
R1168 B.n194 B.n89 9.36635
R1169 B.n580 B.t1 8.47457
R1170 B.n662 B.t3 8.47457
R1171 B.n682 B.n0 8.11757
R1172 B.n682 B.n1 8.11757
R1173 B.n458 B.n457 1.24928
R1174 B.n438 B.n437 1.24928
R1175 B.n174 B.n92 1.24928
R1176 B.n191 B.n89 1.24928
R1177 VP.n2 VP.t2 270.916
R1178 VP.n2 VP.t1 270.697
R1179 VP.n3 VP.t3 234.924
R1180 VP.n9 VP.t0 234.924
R1181 VP.n4 VP.n3 173.105
R1182 VP.n10 VP.n9 173.105
R1183 VP.n8 VP.n0 161.3
R1184 VP.n7 VP.n6 161.3
R1185 VP.n5 VP.n1 161.3
R1186 VP.n4 VP.n2 60.0738
R1187 VP.n7 VP.n1 40.577
R1188 VP.n8 VP.n7 40.577
R1189 VP.n3 VP.n1 12.7883
R1190 VP.n9 VP.n8 12.7883
R1191 VP.n5 VP.n4 0.189894
R1192 VP.n6 VP.n5 0.189894
R1193 VP.n6 VP.n0 0.189894
R1194 VP.n10 VP.n0 0.189894
R1195 VP VP.n10 0.0516364
R1196 VDD1 VDD1.n1 103.379
R1197 VDD1 VDD1.n0 65.2669
R1198 VDD1.n0 VDD1.t1 1.7074
R1199 VDD1.n0 VDD1.t2 1.7074
R1200 VDD1.n1 VDD1.t0 1.7074
R1201 VDD1.n1 VDD1.t3 1.7074
C0 VTAIL VP 3.49833f
C1 VN VTAIL 3.48422f
C2 VDD1 VP 3.93527f
C3 VN VDD1 0.147872f
C4 VN VP 5.10075f
C5 VDD2 VTAIL 5.69575f
C6 VDD2 VDD1 0.681986f
C7 VDD2 VP 0.304731f
C8 VDD2 VN 3.77879f
C9 VTAIL VDD1 5.651f
C10 VDD2 B 2.942922f
C11 VDD1 B 6.60716f
C12 VTAIL B 8.937229f
C13 VN B 8.40988f
C14 VP B 5.909324f
C15 VDD1.t1 B 0.247813f
C16 VDD1.t2 B 0.247813f
C17 VDD1.n0 B 2.21522f
C18 VDD1.t0 B 0.247813f
C19 VDD1.t3 B 0.247813f
C20 VDD1.n1 B 2.8091f
C21 VP.n0 B 0.040236f
C22 VP.t0 B 1.51181f
C23 VP.n1 B 0.061867f
C24 VP.t2 B 1.6023f
C25 VP.t1 B 1.60172f
C26 VP.n2 B 2.47232f
C27 VP.t3 B 1.51181f
C28 VP.n3 B 0.621774f
C29 VP.n4 B 2.22928f
C30 VP.n5 B 0.040236f
C31 VP.n6 B 0.040236f
C32 VP.n7 B 0.032497f
C33 VP.n8 B 0.061867f
C34 VP.n9 B 0.621774f
C35 VP.n10 B 0.036018f
C36 VTAIL.t7 B 1.62107f
C37 VTAIL.n0 B 0.259021f
C38 VTAIL.t2 B 1.62107f
C39 VTAIL.n1 B 0.289874f
C40 VTAIL.t1 B 1.62107f
C41 VTAIL.n2 B 1.06799f
C42 VTAIL.t6 B 1.62107f
C43 VTAIL.n3 B 1.06799f
C44 VTAIL.t4 B 1.62107f
C45 VTAIL.n4 B 0.289875f
C46 VTAIL.t0 B 1.62107f
C47 VTAIL.n5 B 0.289875f
C48 VTAIL.t3 B 1.62106f
C49 VTAIL.n6 B 1.068f
C50 VTAIL.t5 B 1.62107f
C51 VTAIL.n7 B 1.03113f
C52 VDD2.t1 B 0.247809f
C53 VDD2.t2 B 0.247809f
C54 VDD2.n0 B 2.78389f
C55 VDD2.t3 B 0.247809f
C56 VDD2.t0 B 0.247809f
C57 VDD2.n1 B 2.21488f
C58 VDD2.n2 B 3.39002f
C59 VN.t0 B 1.58232f
C60 VN.t2 B 1.58175f
C61 VN.n0 B 1.20672f
C62 VN.t3 B 1.58232f
C63 VN.t1 B 1.58175f
C64 VN.n1 B 2.46307f
.ends

