* NGSPICE file created from diff_pair_sample_1398.ext - technology: sky130A

.subckt diff_pair_sample_1398 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2302_n2160# sky130_fd_pr__pfet_01v8 ad=2.3244 pd=12.7 as=0 ps=0 w=5.96 l=3
X1 VDD2.t1 VN.t0 VTAIL.t3 w_n2302_n2160# sky130_fd_pr__pfet_01v8 ad=2.3244 pd=12.7 as=2.3244 ps=12.7 w=5.96 l=3
X2 VDD1.t1 VP.t0 VTAIL.t1 w_n2302_n2160# sky130_fd_pr__pfet_01v8 ad=2.3244 pd=12.7 as=2.3244 ps=12.7 w=5.96 l=3
X3 VDD2.t0 VN.t1 VTAIL.t2 w_n2302_n2160# sky130_fd_pr__pfet_01v8 ad=2.3244 pd=12.7 as=2.3244 ps=12.7 w=5.96 l=3
X4 VDD1.t0 VP.t1 VTAIL.t0 w_n2302_n2160# sky130_fd_pr__pfet_01v8 ad=2.3244 pd=12.7 as=2.3244 ps=12.7 w=5.96 l=3
X5 B.t8 B.t6 B.t7 w_n2302_n2160# sky130_fd_pr__pfet_01v8 ad=2.3244 pd=12.7 as=0 ps=0 w=5.96 l=3
X6 B.t5 B.t3 B.t4 w_n2302_n2160# sky130_fd_pr__pfet_01v8 ad=2.3244 pd=12.7 as=0 ps=0 w=5.96 l=3
X7 B.t2 B.t0 B.t1 w_n2302_n2160# sky130_fd_pr__pfet_01v8 ad=2.3244 pd=12.7 as=0 ps=0 w=5.96 l=3
R0 B.n248 B.n247 585
R1 B.n246 B.n77 585
R2 B.n245 B.n244 585
R3 B.n243 B.n78 585
R4 B.n242 B.n241 585
R5 B.n240 B.n79 585
R6 B.n239 B.n238 585
R7 B.n237 B.n80 585
R8 B.n236 B.n235 585
R9 B.n234 B.n81 585
R10 B.n233 B.n232 585
R11 B.n231 B.n82 585
R12 B.n230 B.n229 585
R13 B.n228 B.n83 585
R14 B.n227 B.n226 585
R15 B.n225 B.n84 585
R16 B.n224 B.n223 585
R17 B.n222 B.n85 585
R18 B.n221 B.n220 585
R19 B.n219 B.n86 585
R20 B.n218 B.n217 585
R21 B.n216 B.n87 585
R22 B.n215 B.n214 585
R23 B.n213 B.n88 585
R24 B.n212 B.n211 585
R25 B.n207 B.n89 585
R26 B.n206 B.n205 585
R27 B.n204 B.n90 585
R28 B.n203 B.n202 585
R29 B.n201 B.n91 585
R30 B.n200 B.n199 585
R31 B.n198 B.n92 585
R32 B.n197 B.n196 585
R33 B.n194 B.n93 585
R34 B.n193 B.n192 585
R35 B.n191 B.n96 585
R36 B.n190 B.n189 585
R37 B.n188 B.n97 585
R38 B.n187 B.n186 585
R39 B.n185 B.n98 585
R40 B.n184 B.n183 585
R41 B.n182 B.n99 585
R42 B.n181 B.n180 585
R43 B.n179 B.n100 585
R44 B.n178 B.n177 585
R45 B.n176 B.n101 585
R46 B.n175 B.n174 585
R47 B.n173 B.n102 585
R48 B.n172 B.n171 585
R49 B.n170 B.n103 585
R50 B.n169 B.n168 585
R51 B.n167 B.n104 585
R52 B.n166 B.n165 585
R53 B.n164 B.n105 585
R54 B.n163 B.n162 585
R55 B.n161 B.n106 585
R56 B.n160 B.n159 585
R57 B.n249 B.n76 585
R58 B.n251 B.n250 585
R59 B.n252 B.n75 585
R60 B.n254 B.n253 585
R61 B.n255 B.n74 585
R62 B.n257 B.n256 585
R63 B.n258 B.n73 585
R64 B.n260 B.n259 585
R65 B.n261 B.n72 585
R66 B.n263 B.n262 585
R67 B.n264 B.n71 585
R68 B.n266 B.n265 585
R69 B.n267 B.n70 585
R70 B.n269 B.n268 585
R71 B.n270 B.n69 585
R72 B.n272 B.n271 585
R73 B.n273 B.n68 585
R74 B.n275 B.n274 585
R75 B.n276 B.n67 585
R76 B.n278 B.n277 585
R77 B.n279 B.n66 585
R78 B.n281 B.n280 585
R79 B.n282 B.n65 585
R80 B.n284 B.n283 585
R81 B.n285 B.n64 585
R82 B.n287 B.n286 585
R83 B.n288 B.n63 585
R84 B.n290 B.n289 585
R85 B.n291 B.n62 585
R86 B.n293 B.n292 585
R87 B.n294 B.n61 585
R88 B.n296 B.n295 585
R89 B.n297 B.n60 585
R90 B.n299 B.n298 585
R91 B.n300 B.n59 585
R92 B.n302 B.n301 585
R93 B.n303 B.n58 585
R94 B.n305 B.n304 585
R95 B.n306 B.n57 585
R96 B.n308 B.n307 585
R97 B.n309 B.n56 585
R98 B.n311 B.n310 585
R99 B.n312 B.n55 585
R100 B.n314 B.n313 585
R101 B.n315 B.n54 585
R102 B.n317 B.n316 585
R103 B.n318 B.n53 585
R104 B.n320 B.n319 585
R105 B.n321 B.n52 585
R106 B.n323 B.n322 585
R107 B.n324 B.n51 585
R108 B.n326 B.n325 585
R109 B.n327 B.n50 585
R110 B.n329 B.n328 585
R111 B.n330 B.n49 585
R112 B.n332 B.n331 585
R113 B.n419 B.n418 585
R114 B.n417 B.n16 585
R115 B.n416 B.n415 585
R116 B.n414 B.n17 585
R117 B.n413 B.n412 585
R118 B.n411 B.n18 585
R119 B.n410 B.n409 585
R120 B.n408 B.n19 585
R121 B.n407 B.n406 585
R122 B.n405 B.n20 585
R123 B.n404 B.n403 585
R124 B.n402 B.n21 585
R125 B.n401 B.n400 585
R126 B.n399 B.n22 585
R127 B.n398 B.n397 585
R128 B.n396 B.n23 585
R129 B.n395 B.n394 585
R130 B.n393 B.n24 585
R131 B.n392 B.n391 585
R132 B.n390 B.n25 585
R133 B.n389 B.n388 585
R134 B.n387 B.n26 585
R135 B.n386 B.n385 585
R136 B.n384 B.n27 585
R137 B.n382 B.n381 585
R138 B.n380 B.n30 585
R139 B.n379 B.n378 585
R140 B.n377 B.n31 585
R141 B.n376 B.n375 585
R142 B.n374 B.n32 585
R143 B.n373 B.n372 585
R144 B.n371 B.n33 585
R145 B.n370 B.n369 585
R146 B.n368 B.n367 585
R147 B.n366 B.n37 585
R148 B.n365 B.n364 585
R149 B.n363 B.n38 585
R150 B.n362 B.n361 585
R151 B.n360 B.n39 585
R152 B.n359 B.n358 585
R153 B.n357 B.n40 585
R154 B.n356 B.n355 585
R155 B.n354 B.n41 585
R156 B.n353 B.n352 585
R157 B.n351 B.n42 585
R158 B.n350 B.n349 585
R159 B.n348 B.n43 585
R160 B.n347 B.n346 585
R161 B.n345 B.n44 585
R162 B.n344 B.n343 585
R163 B.n342 B.n45 585
R164 B.n341 B.n340 585
R165 B.n339 B.n46 585
R166 B.n338 B.n337 585
R167 B.n336 B.n47 585
R168 B.n335 B.n334 585
R169 B.n333 B.n48 585
R170 B.n420 B.n15 585
R171 B.n422 B.n421 585
R172 B.n423 B.n14 585
R173 B.n425 B.n424 585
R174 B.n426 B.n13 585
R175 B.n428 B.n427 585
R176 B.n429 B.n12 585
R177 B.n431 B.n430 585
R178 B.n432 B.n11 585
R179 B.n434 B.n433 585
R180 B.n435 B.n10 585
R181 B.n437 B.n436 585
R182 B.n438 B.n9 585
R183 B.n440 B.n439 585
R184 B.n441 B.n8 585
R185 B.n443 B.n442 585
R186 B.n444 B.n7 585
R187 B.n446 B.n445 585
R188 B.n447 B.n6 585
R189 B.n449 B.n448 585
R190 B.n450 B.n5 585
R191 B.n452 B.n451 585
R192 B.n453 B.n4 585
R193 B.n455 B.n454 585
R194 B.n456 B.n3 585
R195 B.n458 B.n457 585
R196 B.n459 B.n0 585
R197 B.n2 B.n1 585
R198 B.n121 B.n120 585
R199 B.n122 B.n119 585
R200 B.n124 B.n123 585
R201 B.n125 B.n118 585
R202 B.n127 B.n126 585
R203 B.n128 B.n117 585
R204 B.n130 B.n129 585
R205 B.n131 B.n116 585
R206 B.n133 B.n132 585
R207 B.n134 B.n115 585
R208 B.n136 B.n135 585
R209 B.n137 B.n114 585
R210 B.n139 B.n138 585
R211 B.n140 B.n113 585
R212 B.n142 B.n141 585
R213 B.n143 B.n112 585
R214 B.n145 B.n144 585
R215 B.n146 B.n111 585
R216 B.n148 B.n147 585
R217 B.n149 B.n110 585
R218 B.n151 B.n150 585
R219 B.n152 B.n109 585
R220 B.n154 B.n153 585
R221 B.n155 B.n108 585
R222 B.n157 B.n156 585
R223 B.n158 B.n107 585
R224 B.n160 B.n107 554.963
R225 B.n249 B.n248 554.963
R226 B.n333 B.n332 554.963
R227 B.n418 B.n15 554.963
R228 B.n208 B.t7 332
R229 B.n34 B.t5 332
R230 B.n94 B.t1 331.998
R231 B.n28 B.t11 331.998
R232 B.n209 B.t8 267.418
R233 B.n35 B.t4 267.418
R234 B.n95 B.t2 267.418
R235 B.n29 B.t10 267.418
R236 B.n461 B.n460 256.663
R237 B.n94 B.t0 256.459
R238 B.n208 B.t6 256.459
R239 B.n34 B.t3 256.459
R240 B.n28 B.t9 256.459
R241 B.n460 B.n459 235.042
R242 B.n460 B.n2 235.042
R243 B.n161 B.n160 163.367
R244 B.n162 B.n161 163.367
R245 B.n162 B.n105 163.367
R246 B.n166 B.n105 163.367
R247 B.n167 B.n166 163.367
R248 B.n168 B.n167 163.367
R249 B.n168 B.n103 163.367
R250 B.n172 B.n103 163.367
R251 B.n173 B.n172 163.367
R252 B.n174 B.n173 163.367
R253 B.n174 B.n101 163.367
R254 B.n178 B.n101 163.367
R255 B.n179 B.n178 163.367
R256 B.n180 B.n179 163.367
R257 B.n180 B.n99 163.367
R258 B.n184 B.n99 163.367
R259 B.n185 B.n184 163.367
R260 B.n186 B.n185 163.367
R261 B.n186 B.n97 163.367
R262 B.n190 B.n97 163.367
R263 B.n191 B.n190 163.367
R264 B.n192 B.n191 163.367
R265 B.n192 B.n93 163.367
R266 B.n197 B.n93 163.367
R267 B.n198 B.n197 163.367
R268 B.n199 B.n198 163.367
R269 B.n199 B.n91 163.367
R270 B.n203 B.n91 163.367
R271 B.n204 B.n203 163.367
R272 B.n205 B.n204 163.367
R273 B.n205 B.n89 163.367
R274 B.n212 B.n89 163.367
R275 B.n213 B.n212 163.367
R276 B.n214 B.n213 163.367
R277 B.n214 B.n87 163.367
R278 B.n218 B.n87 163.367
R279 B.n219 B.n218 163.367
R280 B.n220 B.n219 163.367
R281 B.n220 B.n85 163.367
R282 B.n224 B.n85 163.367
R283 B.n225 B.n224 163.367
R284 B.n226 B.n225 163.367
R285 B.n226 B.n83 163.367
R286 B.n230 B.n83 163.367
R287 B.n231 B.n230 163.367
R288 B.n232 B.n231 163.367
R289 B.n232 B.n81 163.367
R290 B.n236 B.n81 163.367
R291 B.n237 B.n236 163.367
R292 B.n238 B.n237 163.367
R293 B.n238 B.n79 163.367
R294 B.n242 B.n79 163.367
R295 B.n243 B.n242 163.367
R296 B.n244 B.n243 163.367
R297 B.n244 B.n77 163.367
R298 B.n248 B.n77 163.367
R299 B.n332 B.n49 163.367
R300 B.n328 B.n49 163.367
R301 B.n328 B.n327 163.367
R302 B.n327 B.n326 163.367
R303 B.n326 B.n51 163.367
R304 B.n322 B.n51 163.367
R305 B.n322 B.n321 163.367
R306 B.n321 B.n320 163.367
R307 B.n320 B.n53 163.367
R308 B.n316 B.n53 163.367
R309 B.n316 B.n315 163.367
R310 B.n315 B.n314 163.367
R311 B.n314 B.n55 163.367
R312 B.n310 B.n55 163.367
R313 B.n310 B.n309 163.367
R314 B.n309 B.n308 163.367
R315 B.n308 B.n57 163.367
R316 B.n304 B.n57 163.367
R317 B.n304 B.n303 163.367
R318 B.n303 B.n302 163.367
R319 B.n302 B.n59 163.367
R320 B.n298 B.n59 163.367
R321 B.n298 B.n297 163.367
R322 B.n297 B.n296 163.367
R323 B.n296 B.n61 163.367
R324 B.n292 B.n61 163.367
R325 B.n292 B.n291 163.367
R326 B.n291 B.n290 163.367
R327 B.n290 B.n63 163.367
R328 B.n286 B.n63 163.367
R329 B.n286 B.n285 163.367
R330 B.n285 B.n284 163.367
R331 B.n284 B.n65 163.367
R332 B.n280 B.n65 163.367
R333 B.n280 B.n279 163.367
R334 B.n279 B.n278 163.367
R335 B.n278 B.n67 163.367
R336 B.n274 B.n67 163.367
R337 B.n274 B.n273 163.367
R338 B.n273 B.n272 163.367
R339 B.n272 B.n69 163.367
R340 B.n268 B.n69 163.367
R341 B.n268 B.n267 163.367
R342 B.n267 B.n266 163.367
R343 B.n266 B.n71 163.367
R344 B.n262 B.n71 163.367
R345 B.n262 B.n261 163.367
R346 B.n261 B.n260 163.367
R347 B.n260 B.n73 163.367
R348 B.n256 B.n73 163.367
R349 B.n256 B.n255 163.367
R350 B.n255 B.n254 163.367
R351 B.n254 B.n75 163.367
R352 B.n250 B.n75 163.367
R353 B.n250 B.n249 163.367
R354 B.n418 B.n417 163.367
R355 B.n417 B.n416 163.367
R356 B.n416 B.n17 163.367
R357 B.n412 B.n17 163.367
R358 B.n412 B.n411 163.367
R359 B.n411 B.n410 163.367
R360 B.n410 B.n19 163.367
R361 B.n406 B.n19 163.367
R362 B.n406 B.n405 163.367
R363 B.n405 B.n404 163.367
R364 B.n404 B.n21 163.367
R365 B.n400 B.n21 163.367
R366 B.n400 B.n399 163.367
R367 B.n399 B.n398 163.367
R368 B.n398 B.n23 163.367
R369 B.n394 B.n23 163.367
R370 B.n394 B.n393 163.367
R371 B.n393 B.n392 163.367
R372 B.n392 B.n25 163.367
R373 B.n388 B.n25 163.367
R374 B.n388 B.n387 163.367
R375 B.n387 B.n386 163.367
R376 B.n386 B.n27 163.367
R377 B.n381 B.n27 163.367
R378 B.n381 B.n380 163.367
R379 B.n380 B.n379 163.367
R380 B.n379 B.n31 163.367
R381 B.n375 B.n31 163.367
R382 B.n375 B.n374 163.367
R383 B.n374 B.n373 163.367
R384 B.n373 B.n33 163.367
R385 B.n369 B.n33 163.367
R386 B.n369 B.n368 163.367
R387 B.n368 B.n37 163.367
R388 B.n364 B.n37 163.367
R389 B.n364 B.n363 163.367
R390 B.n363 B.n362 163.367
R391 B.n362 B.n39 163.367
R392 B.n358 B.n39 163.367
R393 B.n358 B.n357 163.367
R394 B.n357 B.n356 163.367
R395 B.n356 B.n41 163.367
R396 B.n352 B.n41 163.367
R397 B.n352 B.n351 163.367
R398 B.n351 B.n350 163.367
R399 B.n350 B.n43 163.367
R400 B.n346 B.n43 163.367
R401 B.n346 B.n345 163.367
R402 B.n345 B.n344 163.367
R403 B.n344 B.n45 163.367
R404 B.n340 B.n45 163.367
R405 B.n340 B.n339 163.367
R406 B.n339 B.n338 163.367
R407 B.n338 B.n47 163.367
R408 B.n334 B.n47 163.367
R409 B.n334 B.n333 163.367
R410 B.n422 B.n15 163.367
R411 B.n423 B.n422 163.367
R412 B.n424 B.n423 163.367
R413 B.n424 B.n13 163.367
R414 B.n428 B.n13 163.367
R415 B.n429 B.n428 163.367
R416 B.n430 B.n429 163.367
R417 B.n430 B.n11 163.367
R418 B.n434 B.n11 163.367
R419 B.n435 B.n434 163.367
R420 B.n436 B.n435 163.367
R421 B.n436 B.n9 163.367
R422 B.n440 B.n9 163.367
R423 B.n441 B.n440 163.367
R424 B.n442 B.n441 163.367
R425 B.n442 B.n7 163.367
R426 B.n446 B.n7 163.367
R427 B.n447 B.n446 163.367
R428 B.n448 B.n447 163.367
R429 B.n448 B.n5 163.367
R430 B.n452 B.n5 163.367
R431 B.n453 B.n452 163.367
R432 B.n454 B.n453 163.367
R433 B.n454 B.n3 163.367
R434 B.n458 B.n3 163.367
R435 B.n459 B.n458 163.367
R436 B.n120 B.n2 163.367
R437 B.n120 B.n119 163.367
R438 B.n124 B.n119 163.367
R439 B.n125 B.n124 163.367
R440 B.n126 B.n125 163.367
R441 B.n126 B.n117 163.367
R442 B.n130 B.n117 163.367
R443 B.n131 B.n130 163.367
R444 B.n132 B.n131 163.367
R445 B.n132 B.n115 163.367
R446 B.n136 B.n115 163.367
R447 B.n137 B.n136 163.367
R448 B.n138 B.n137 163.367
R449 B.n138 B.n113 163.367
R450 B.n142 B.n113 163.367
R451 B.n143 B.n142 163.367
R452 B.n144 B.n143 163.367
R453 B.n144 B.n111 163.367
R454 B.n148 B.n111 163.367
R455 B.n149 B.n148 163.367
R456 B.n150 B.n149 163.367
R457 B.n150 B.n109 163.367
R458 B.n154 B.n109 163.367
R459 B.n155 B.n154 163.367
R460 B.n156 B.n155 163.367
R461 B.n156 B.n107 163.367
R462 B.n95 B.n94 64.5823
R463 B.n209 B.n208 64.5823
R464 B.n35 B.n34 64.5823
R465 B.n29 B.n28 64.5823
R466 B.n195 B.n95 59.5399
R467 B.n210 B.n209 59.5399
R468 B.n36 B.n35 59.5399
R469 B.n383 B.n29 59.5399
R470 B.n420 B.n419 36.059
R471 B.n331 B.n48 36.059
R472 B.n247 B.n76 36.059
R473 B.n159 B.n158 36.059
R474 B B.n461 18.0485
R475 B.n421 B.n420 10.6151
R476 B.n421 B.n14 10.6151
R477 B.n425 B.n14 10.6151
R478 B.n426 B.n425 10.6151
R479 B.n427 B.n426 10.6151
R480 B.n427 B.n12 10.6151
R481 B.n431 B.n12 10.6151
R482 B.n432 B.n431 10.6151
R483 B.n433 B.n432 10.6151
R484 B.n433 B.n10 10.6151
R485 B.n437 B.n10 10.6151
R486 B.n438 B.n437 10.6151
R487 B.n439 B.n438 10.6151
R488 B.n439 B.n8 10.6151
R489 B.n443 B.n8 10.6151
R490 B.n444 B.n443 10.6151
R491 B.n445 B.n444 10.6151
R492 B.n445 B.n6 10.6151
R493 B.n449 B.n6 10.6151
R494 B.n450 B.n449 10.6151
R495 B.n451 B.n450 10.6151
R496 B.n451 B.n4 10.6151
R497 B.n455 B.n4 10.6151
R498 B.n456 B.n455 10.6151
R499 B.n457 B.n456 10.6151
R500 B.n457 B.n0 10.6151
R501 B.n419 B.n16 10.6151
R502 B.n415 B.n16 10.6151
R503 B.n415 B.n414 10.6151
R504 B.n414 B.n413 10.6151
R505 B.n413 B.n18 10.6151
R506 B.n409 B.n18 10.6151
R507 B.n409 B.n408 10.6151
R508 B.n408 B.n407 10.6151
R509 B.n407 B.n20 10.6151
R510 B.n403 B.n20 10.6151
R511 B.n403 B.n402 10.6151
R512 B.n402 B.n401 10.6151
R513 B.n401 B.n22 10.6151
R514 B.n397 B.n22 10.6151
R515 B.n397 B.n396 10.6151
R516 B.n396 B.n395 10.6151
R517 B.n395 B.n24 10.6151
R518 B.n391 B.n24 10.6151
R519 B.n391 B.n390 10.6151
R520 B.n390 B.n389 10.6151
R521 B.n389 B.n26 10.6151
R522 B.n385 B.n26 10.6151
R523 B.n385 B.n384 10.6151
R524 B.n382 B.n30 10.6151
R525 B.n378 B.n30 10.6151
R526 B.n378 B.n377 10.6151
R527 B.n377 B.n376 10.6151
R528 B.n376 B.n32 10.6151
R529 B.n372 B.n32 10.6151
R530 B.n372 B.n371 10.6151
R531 B.n371 B.n370 10.6151
R532 B.n367 B.n366 10.6151
R533 B.n366 B.n365 10.6151
R534 B.n365 B.n38 10.6151
R535 B.n361 B.n38 10.6151
R536 B.n361 B.n360 10.6151
R537 B.n360 B.n359 10.6151
R538 B.n359 B.n40 10.6151
R539 B.n355 B.n40 10.6151
R540 B.n355 B.n354 10.6151
R541 B.n354 B.n353 10.6151
R542 B.n353 B.n42 10.6151
R543 B.n349 B.n42 10.6151
R544 B.n349 B.n348 10.6151
R545 B.n348 B.n347 10.6151
R546 B.n347 B.n44 10.6151
R547 B.n343 B.n44 10.6151
R548 B.n343 B.n342 10.6151
R549 B.n342 B.n341 10.6151
R550 B.n341 B.n46 10.6151
R551 B.n337 B.n46 10.6151
R552 B.n337 B.n336 10.6151
R553 B.n336 B.n335 10.6151
R554 B.n335 B.n48 10.6151
R555 B.n331 B.n330 10.6151
R556 B.n330 B.n329 10.6151
R557 B.n329 B.n50 10.6151
R558 B.n325 B.n50 10.6151
R559 B.n325 B.n324 10.6151
R560 B.n324 B.n323 10.6151
R561 B.n323 B.n52 10.6151
R562 B.n319 B.n52 10.6151
R563 B.n319 B.n318 10.6151
R564 B.n318 B.n317 10.6151
R565 B.n317 B.n54 10.6151
R566 B.n313 B.n54 10.6151
R567 B.n313 B.n312 10.6151
R568 B.n312 B.n311 10.6151
R569 B.n311 B.n56 10.6151
R570 B.n307 B.n56 10.6151
R571 B.n307 B.n306 10.6151
R572 B.n306 B.n305 10.6151
R573 B.n305 B.n58 10.6151
R574 B.n301 B.n58 10.6151
R575 B.n301 B.n300 10.6151
R576 B.n300 B.n299 10.6151
R577 B.n299 B.n60 10.6151
R578 B.n295 B.n60 10.6151
R579 B.n295 B.n294 10.6151
R580 B.n294 B.n293 10.6151
R581 B.n293 B.n62 10.6151
R582 B.n289 B.n62 10.6151
R583 B.n289 B.n288 10.6151
R584 B.n288 B.n287 10.6151
R585 B.n287 B.n64 10.6151
R586 B.n283 B.n64 10.6151
R587 B.n283 B.n282 10.6151
R588 B.n282 B.n281 10.6151
R589 B.n281 B.n66 10.6151
R590 B.n277 B.n66 10.6151
R591 B.n277 B.n276 10.6151
R592 B.n276 B.n275 10.6151
R593 B.n275 B.n68 10.6151
R594 B.n271 B.n68 10.6151
R595 B.n271 B.n270 10.6151
R596 B.n270 B.n269 10.6151
R597 B.n269 B.n70 10.6151
R598 B.n265 B.n70 10.6151
R599 B.n265 B.n264 10.6151
R600 B.n264 B.n263 10.6151
R601 B.n263 B.n72 10.6151
R602 B.n259 B.n72 10.6151
R603 B.n259 B.n258 10.6151
R604 B.n258 B.n257 10.6151
R605 B.n257 B.n74 10.6151
R606 B.n253 B.n74 10.6151
R607 B.n253 B.n252 10.6151
R608 B.n252 B.n251 10.6151
R609 B.n251 B.n76 10.6151
R610 B.n121 B.n1 10.6151
R611 B.n122 B.n121 10.6151
R612 B.n123 B.n122 10.6151
R613 B.n123 B.n118 10.6151
R614 B.n127 B.n118 10.6151
R615 B.n128 B.n127 10.6151
R616 B.n129 B.n128 10.6151
R617 B.n129 B.n116 10.6151
R618 B.n133 B.n116 10.6151
R619 B.n134 B.n133 10.6151
R620 B.n135 B.n134 10.6151
R621 B.n135 B.n114 10.6151
R622 B.n139 B.n114 10.6151
R623 B.n140 B.n139 10.6151
R624 B.n141 B.n140 10.6151
R625 B.n141 B.n112 10.6151
R626 B.n145 B.n112 10.6151
R627 B.n146 B.n145 10.6151
R628 B.n147 B.n146 10.6151
R629 B.n147 B.n110 10.6151
R630 B.n151 B.n110 10.6151
R631 B.n152 B.n151 10.6151
R632 B.n153 B.n152 10.6151
R633 B.n153 B.n108 10.6151
R634 B.n157 B.n108 10.6151
R635 B.n158 B.n157 10.6151
R636 B.n159 B.n106 10.6151
R637 B.n163 B.n106 10.6151
R638 B.n164 B.n163 10.6151
R639 B.n165 B.n164 10.6151
R640 B.n165 B.n104 10.6151
R641 B.n169 B.n104 10.6151
R642 B.n170 B.n169 10.6151
R643 B.n171 B.n170 10.6151
R644 B.n171 B.n102 10.6151
R645 B.n175 B.n102 10.6151
R646 B.n176 B.n175 10.6151
R647 B.n177 B.n176 10.6151
R648 B.n177 B.n100 10.6151
R649 B.n181 B.n100 10.6151
R650 B.n182 B.n181 10.6151
R651 B.n183 B.n182 10.6151
R652 B.n183 B.n98 10.6151
R653 B.n187 B.n98 10.6151
R654 B.n188 B.n187 10.6151
R655 B.n189 B.n188 10.6151
R656 B.n189 B.n96 10.6151
R657 B.n193 B.n96 10.6151
R658 B.n194 B.n193 10.6151
R659 B.n196 B.n92 10.6151
R660 B.n200 B.n92 10.6151
R661 B.n201 B.n200 10.6151
R662 B.n202 B.n201 10.6151
R663 B.n202 B.n90 10.6151
R664 B.n206 B.n90 10.6151
R665 B.n207 B.n206 10.6151
R666 B.n211 B.n207 10.6151
R667 B.n215 B.n88 10.6151
R668 B.n216 B.n215 10.6151
R669 B.n217 B.n216 10.6151
R670 B.n217 B.n86 10.6151
R671 B.n221 B.n86 10.6151
R672 B.n222 B.n221 10.6151
R673 B.n223 B.n222 10.6151
R674 B.n223 B.n84 10.6151
R675 B.n227 B.n84 10.6151
R676 B.n228 B.n227 10.6151
R677 B.n229 B.n228 10.6151
R678 B.n229 B.n82 10.6151
R679 B.n233 B.n82 10.6151
R680 B.n234 B.n233 10.6151
R681 B.n235 B.n234 10.6151
R682 B.n235 B.n80 10.6151
R683 B.n239 B.n80 10.6151
R684 B.n240 B.n239 10.6151
R685 B.n241 B.n240 10.6151
R686 B.n241 B.n78 10.6151
R687 B.n245 B.n78 10.6151
R688 B.n246 B.n245 10.6151
R689 B.n247 B.n246 10.6151
R690 B.n461 B.n0 8.11757
R691 B.n461 B.n1 8.11757
R692 B.n383 B.n382 6.5566
R693 B.n370 B.n36 6.5566
R694 B.n196 B.n195 6.5566
R695 B.n211 B.n210 6.5566
R696 B.n384 B.n383 4.05904
R697 B.n367 B.n36 4.05904
R698 B.n195 B.n194 4.05904
R699 B.n210 B.n88 4.05904
R700 VN VN.t1 130.161
R701 VN VN.t0 89.4482
R702 VTAIL.n122 VTAIL.n96 756.745
R703 VTAIL.n26 VTAIL.n0 756.745
R704 VTAIL.n90 VTAIL.n64 756.745
R705 VTAIL.n58 VTAIL.n32 756.745
R706 VTAIL.n107 VTAIL.n106 585
R707 VTAIL.n104 VTAIL.n103 585
R708 VTAIL.n113 VTAIL.n112 585
R709 VTAIL.n115 VTAIL.n114 585
R710 VTAIL.n100 VTAIL.n99 585
R711 VTAIL.n121 VTAIL.n120 585
R712 VTAIL.n123 VTAIL.n122 585
R713 VTAIL.n11 VTAIL.n10 585
R714 VTAIL.n8 VTAIL.n7 585
R715 VTAIL.n17 VTAIL.n16 585
R716 VTAIL.n19 VTAIL.n18 585
R717 VTAIL.n4 VTAIL.n3 585
R718 VTAIL.n25 VTAIL.n24 585
R719 VTAIL.n27 VTAIL.n26 585
R720 VTAIL.n91 VTAIL.n90 585
R721 VTAIL.n89 VTAIL.n88 585
R722 VTAIL.n68 VTAIL.n67 585
R723 VTAIL.n83 VTAIL.n82 585
R724 VTAIL.n81 VTAIL.n80 585
R725 VTAIL.n72 VTAIL.n71 585
R726 VTAIL.n75 VTAIL.n74 585
R727 VTAIL.n59 VTAIL.n58 585
R728 VTAIL.n57 VTAIL.n56 585
R729 VTAIL.n36 VTAIL.n35 585
R730 VTAIL.n51 VTAIL.n50 585
R731 VTAIL.n49 VTAIL.n48 585
R732 VTAIL.n40 VTAIL.n39 585
R733 VTAIL.n43 VTAIL.n42 585
R734 VTAIL.t3 VTAIL.n105 327.601
R735 VTAIL.t1 VTAIL.n9 327.601
R736 VTAIL.t0 VTAIL.n73 327.601
R737 VTAIL.t2 VTAIL.n41 327.601
R738 VTAIL.n106 VTAIL.n103 171.744
R739 VTAIL.n113 VTAIL.n103 171.744
R740 VTAIL.n114 VTAIL.n113 171.744
R741 VTAIL.n114 VTAIL.n99 171.744
R742 VTAIL.n121 VTAIL.n99 171.744
R743 VTAIL.n122 VTAIL.n121 171.744
R744 VTAIL.n10 VTAIL.n7 171.744
R745 VTAIL.n17 VTAIL.n7 171.744
R746 VTAIL.n18 VTAIL.n17 171.744
R747 VTAIL.n18 VTAIL.n3 171.744
R748 VTAIL.n25 VTAIL.n3 171.744
R749 VTAIL.n26 VTAIL.n25 171.744
R750 VTAIL.n90 VTAIL.n89 171.744
R751 VTAIL.n89 VTAIL.n67 171.744
R752 VTAIL.n82 VTAIL.n67 171.744
R753 VTAIL.n82 VTAIL.n81 171.744
R754 VTAIL.n81 VTAIL.n71 171.744
R755 VTAIL.n74 VTAIL.n71 171.744
R756 VTAIL.n58 VTAIL.n57 171.744
R757 VTAIL.n57 VTAIL.n35 171.744
R758 VTAIL.n50 VTAIL.n35 171.744
R759 VTAIL.n50 VTAIL.n49 171.744
R760 VTAIL.n49 VTAIL.n39 171.744
R761 VTAIL.n42 VTAIL.n39 171.744
R762 VTAIL.n106 VTAIL.t3 85.8723
R763 VTAIL.n10 VTAIL.t1 85.8723
R764 VTAIL.n74 VTAIL.t0 85.8723
R765 VTAIL.n42 VTAIL.t2 85.8723
R766 VTAIL.n127 VTAIL.n126 31.4096
R767 VTAIL.n31 VTAIL.n30 31.4096
R768 VTAIL.n95 VTAIL.n94 31.4096
R769 VTAIL.n63 VTAIL.n62 31.4096
R770 VTAIL.n63 VTAIL.n31 23.2462
R771 VTAIL.n127 VTAIL.n95 20.3755
R772 VTAIL.n107 VTAIL.n105 16.3865
R773 VTAIL.n11 VTAIL.n9 16.3865
R774 VTAIL.n75 VTAIL.n73 16.3865
R775 VTAIL.n43 VTAIL.n41 16.3865
R776 VTAIL.n108 VTAIL.n104 12.8005
R777 VTAIL.n12 VTAIL.n8 12.8005
R778 VTAIL.n76 VTAIL.n72 12.8005
R779 VTAIL.n44 VTAIL.n40 12.8005
R780 VTAIL.n112 VTAIL.n111 12.0247
R781 VTAIL.n16 VTAIL.n15 12.0247
R782 VTAIL.n80 VTAIL.n79 12.0247
R783 VTAIL.n48 VTAIL.n47 12.0247
R784 VTAIL.n115 VTAIL.n102 11.249
R785 VTAIL.n19 VTAIL.n6 11.249
R786 VTAIL.n83 VTAIL.n70 11.249
R787 VTAIL.n51 VTAIL.n38 11.249
R788 VTAIL.n116 VTAIL.n100 10.4732
R789 VTAIL.n20 VTAIL.n4 10.4732
R790 VTAIL.n84 VTAIL.n68 10.4732
R791 VTAIL.n52 VTAIL.n36 10.4732
R792 VTAIL.n120 VTAIL.n119 9.69747
R793 VTAIL.n24 VTAIL.n23 9.69747
R794 VTAIL.n88 VTAIL.n87 9.69747
R795 VTAIL.n56 VTAIL.n55 9.69747
R796 VTAIL.n126 VTAIL.n125 9.45567
R797 VTAIL.n30 VTAIL.n29 9.45567
R798 VTAIL.n94 VTAIL.n93 9.45567
R799 VTAIL.n62 VTAIL.n61 9.45567
R800 VTAIL.n125 VTAIL.n124 9.3005
R801 VTAIL.n98 VTAIL.n97 9.3005
R802 VTAIL.n119 VTAIL.n118 9.3005
R803 VTAIL.n117 VTAIL.n116 9.3005
R804 VTAIL.n102 VTAIL.n101 9.3005
R805 VTAIL.n111 VTAIL.n110 9.3005
R806 VTAIL.n109 VTAIL.n108 9.3005
R807 VTAIL.n29 VTAIL.n28 9.3005
R808 VTAIL.n2 VTAIL.n1 9.3005
R809 VTAIL.n23 VTAIL.n22 9.3005
R810 VTAIL.n21 VTAIL.n20 9.3005
R811 VTAIL.n6 VTAIL.n5 9.3005
R812 VTAIL.n15 VTAIL.n14 9.3005
R813 VTAIL.n13 VTAIL.n12 9.3005
R814 VTAIL.n93 VTAIL.n92 9.3005
R815 VTAIL.n66 VTAIL.n65 9.3005
R816 VTAIL.n87 VTAIL.n86 9.3005
R817 VTAIL.n85 VTAIL.n84 9.3005
R818 VTAIL.n70 VTAIL.n69 9.3005
R819 VTAIL.n79 VTAIL.n78 9.3005
R820 VTAIL.n77 VTAIL.n76 9.3005
R821 VTAIL.n61 VTAIL.n60 9.3005
R822 VTAIL.n34 VTAIL.n33 9.3005
R823 VTAIL.n55 VTAIL.n54 9.3005
R824 VTAIL.n53 VTAIL.n52 9.3005
R825 VTAIL.n38 VTAIL.n37 9.3005
R826 VTAIL.n47 VTAIL.n46 9.3005
R827 VTAIL.n45 VTAIL.n44 9.3005
R828 VTAIL.n123 VTAIL.n98 8.92171
R829 VTAIL.n27 VTAIL.n2 8.92171
R830 VTAIL.n91 VTAIL.n66 8.92171
R831 VTAIL.n59 VTAIL.n34 8.92171
R832 VTAIL.n124 VTAIL.n96 8.14595
R833 VTAIL.n28 VTAIL.n0 8.14595
R834 VTAIL.n92 VTAIL.n64 8.14595
R835 VTAIL.n60 VTAIL.n32 8.14595
R836 VTAIL.n126 VTAIL.n96 5.81868
R837 VTAIL.n30 VTAIL.n0 5.81868
R838 VTAIL.n94 VTAIL.n64 5.81868
R839 VTAIL.n62 VTAIL.n32 5.81868
R840 VTAIL.n124 VTAIL.n123 5.04292
R841 VTAIL.n28 VTAIL.n27 5.04292
R842 VTAIL.n92 VTAIL.n91 5.04292
R843 VTAIL.n60 VTAIL.n59 5.04292
R844 VTAIL.n120 VTAIL.n98 4.26717
R845 VTAIL.n24 VTAIL.n2 4.26717
R846 VTAIL.n88 VTAIL.n66 4.26717
R847 VTAIL.n56 VTAIL.n34 4.26717
R848 VTAIL.n77 VTAIL.n73 3.71286
R849 VTAIL.n45 VTAIL.n41 3.71286
R850 VTAIL.n109 VTAIL.n105 3.71286
R851 VTAIL.n13 VTAIL.n9 3.71286
R852 VTAIL.n119 VTAIL.n100 3.49141
R853 VTAIL.n23 VTAIL.n4 3.49141
R854 VTAIL.n87 VTAIL.n68 3.49141
R855 VTAIL.n55 VTAIL.n36 3.49141
R856 VTAIL.n116 VTAIL.n115 2.71565
R857 VTAIL.n20 VTAIL.n19 2.71565
R858 VTAIL.n84 VTAIL.n83 2.71565
R859 VTAIL.n52 VTAIL.n51 2.71565
R860 VTAIL.n112 VTAIL.n102 1.93989
R861 VTAIL.n16 VTAIL.n6 1.93989
R862 VTAIL.n80 VTAIL.n70 1.93989
R863 VTAIL.n48 VTAIL.n38 1.93989
R864 VTAIL.n95 VTAIL.n63 1.90567
R865 VTAIL VTAIL.n31 1.24619
R866 VTAIL.n111 VTAIL.n104 1.16414
R867 VTAIL.n15 VTAIL.n8 1.16414
R868 VTAIL.n79 VTAIL.n72 1.16414
R869 VTAIL.n47 VTAIL.n40 1.16414
R870 VTAIL VTAIL.n127 0.659983
R871 VTAIL.n108 VTAIL.n107 0.388379
R872 VTAIL.n12 VTAIL.n11 0.388379
R873 VTAIL.n76 VTAIL.n75 0.388379
R874 VTAIL.n44 VTAIL.n43 0.388379
R875 VTAIL.n110 VTAIL.n109 0.155672
R876 VTAIL.n110 VTAIL.n101 0.155672
R877 VTAIL.n117 VTAIL.n101 0.155672
R878 VTAIL.n118 VTAIL.n117 0.155672
R879 VTAIL.n118 VTAIL.n97 0.155672
R880 VTAIL.n125 VTAIL.n97 0.155672
R881 VTAIL.n14 VTAIL.n13 0.155672
R882 VTAIL.n14 VTAIL.n5 0.155672
R883 VTAIL.n21 VTAIL.n5 0.155672
R884 VTAIL.n22 VTAIL.n21 0.155672
R885 VTAIL.n22 VTAIL.n1 0.155672
R886 VTAIL.n29 VTAIL.n1 0.155672
R887 VTAIL.n93 VTAIL.n65 0.155672
R888 VTAIL.n86 VTAIL.n65 0.155672
R889 VTAIL.n86 VTAIL.n85 0.155672
R890 VTAIL.n85 VTAIL.n69 0.155672
R891 VTAIL.n78 VTAIL.n69 0.155672
R892 VTAIL.n78 VTAIL.n77 0.155672
R893 VTAIL.n61 VTAIL.n33 0.155672
R894 VTAIL.n54 VTAIL.n33 0.155672
R895 VTAIL.n54 VTAIL.n53 0.155672
R896 VTAIL.n53 VTAIL.n37 0.155672
R897 VTAIL.n46 VTAIL.n37 0.155672
R898 VTAIL.n46 VTAIL.n45 0.155672
R899 VDD2.n57 VDD2.n31 756.745
R900 VDD2.n26 VDD2.n0 756.745
R901 VDD2.n58 VDD2.n57 585
R902 VDD2.n56 VDD2.n55 585
R903 VDD2.n35 VDD2.n34 585
R904 VDD2.n50 VDD2.n49 585
R905 VDD2.n48 VDD2.n47 585
R906 VDD2.n39 VDD2.n38 585
R907 VDD2.n42 VDD2.n41 585
R908 VDD2.n11 VDD2.n10 585
R909 VDD2.n8 VDD2.n7 585
R910 VDD2.n17 VDD2.n16 585
R911 VDD2.n19 VDD2.n18 585
R912 VDD2.n4 VDD2.n3 585
R913 VDD2.n25 VDD2.n24 585
R914 VDD2.n27 VDD2.n26 585
R915 VDD2.t0 VDD2.n40 327.601
R916 VDD2.t1 VDD2.n9 327.601
R917 VDD2.n57 VDD2.n56 171.744
R918 VDD2.n56 VDD2.n34 171.744
R919 VDD2.n49 VDD2.n34 171.744
R920 VDD2.n49 VDD2.n48 171.744
R921 VDD2.n48 VDD2.n38 171.744
R922 VDD2.n41 VDD2.n38 171.744
R923 VDD2.n10 VDD2.n7 171.744
R924 VDD2.n17 VDD2.n7 171.744
R925 VDD2.n18 VDD2.n17 171.744
R926 VDD2.n18 VDD2.n3 171.744
R927 VDD2.n25 VDD2.n3 171.744
R928 VDD2.n26 VDD2.n25 171.744
R929 VDD2.n41 VDD2.t0 85.8723
R930 VDD2.n10 VDD2.t1 85.8723
R931 VDD2.n62 VDD2.n30 82.6271
R932 VDD2.n62 VDD2.n61 48.0884
R933 VDD2.n42 VDD2.n40 16.3865
R934 VDD2.n11 VDD2.n9 16.3865
R935 VDD2.n43 VDD2.n39 12.8005
R936 VDD2.n12 VDD2.n8 12.8005
R937 VDD2.n47 VDD2.n46 12.0247
R938 VDD2.n16 VDD2.n15 12.0247
R939 VDD2.n50 VDD2.n37 11.249
R940 VDD2.n19 VDD2.n6 11.249
R941 VDD2.n51 VDD2.n35 10.4732
R942 VDD2.n20 VDD2.n4 10.4732
R943 VDD2.n55 VDD2.n54 9.69747
R944 VDD2.n24 VDD2.n23 9.69747
R945 VDD2.n61 VDD2.n60 9.45567
R946 VDD2.n30 VDD2.n29 9.45567
R947 VDD2.n60 VDD2.n59 9.3005
R948 VDD2.n33 VDD2.n32 9.3005
R949 VDD2.n54 VDD2.n53 9.3005
R950 VDD2.n52 VDD2.n51 9.3005
R951 VDD2.n37 VDD2.n36 9.3005
R952 VDD2.n46 VDD2.n45 9.3005
R953 VDD2.n44 VDD2.n43 9.3005
R954 VDD2.n29 VDD2.n28 9.3005
R955 VDD2.n2 VDD2.n1 9.3005
R956 VDD2.n23 VDD2.n22 9.3005
R957 VDD2.n21 VDD2.n20 9.3005
R958 VDD2.n6 VDD2.n5 9.3005
R959 VDD2.n15 VDD2.n14 9.3005
R960 VDD2.n13 VDD2.n12 9.3005
R961 VDD2.n58 VDD2.n33 8.92171
R962 VDD2.n27 VDD2.n2 8.92171
R963 VDD2.n59 VDD2.n31 8.14595
R964 VDD2.n28 VDD2.n0 8.14595
R965 VDD2.n61 VDD2.n31 5.81868
R966 VDD2.n30 VDD2.n0 5.81868
R967 VDD2.n59 VDD2.n58 5.04292
R968 VDD2.n28 VDD2.n27 5.04292
R969 VDD2.n55 VDD2.n33 4.26717
R970 VDD2.n24 VDD2.n2 4.26717
R971 VDD2.n44 VDD2.n40 3.71286
R972 VDD2.n13 VDD2.n9 3.71286
R973 VDD2.n54 VDD2.n35 3.49141
R974 VDD2.n23 VDD2.n4 3.49141
R975 VDD2.n51 VDD2.n50 2.71565
R976 VDD2.n20 VDD2.n19 2.71565
R977 VDD2.n47 VDD2.n37 1.93989
R978 VDD2.n16 VDD2.n6 1.93989
R979 VDD2.n46 VDD2.n39 1.16414
R980 VDD2.n15 VDD2.n8 1.16414
R981 VDD2 VDD2.n62 0.776362
R982 VDD2.n43 VDD2.n42 0.388379
R983 VDD2.n12 VDD2.n11 0.388379
R984 VDD2.n60 VDD2.n32 0.155672
R985 VDD2.n53 VDD2.n32 0.155672
R986 VDD2.n53 VDD2.n52 0.155672
R987 VDD2.n52 VDD2.n36 0.155672
R988 VDD2.n45 VDD2.n36 0.155672
R989 VDD2.n45 VDD2.n44 0.155672
R990 VDD2.n14 VDD2.n13 0.155672
R991 VDD2.n14 VDD2.n5 0.155672
R992 VDD2.n21 VDD2.n5 0.155672
R993 VDD2.n22 VDD2.n21 0.155672
R994 VDD2.n22 VDD2.n1 0.155672
R995 VDD2.n29 VDD2.n1 0.155672
R996 VP.n0 VP.t1 130.159
R997 VP.n0 VP.t0 89.0169
R998 VP VP.n0 0.431812
R999 VDD1.n26 VDD1.n0 756.745
R1000 VDD1.n57 VDD1.n31 756.745
R1001 VDD1.n27 VDD1.n26 585
R1002 VDD1.n25 VDD1.n24 585
R1003 VDD1.n4 VDD1.n3 585
R1004 VDD1.n19 VDD1.n18 585
R1005 VDD1.n17 VDD1.n16 585
R1006 VDD1.n8 VDD1.n7 585
R1007 VDD1.n11 VDD1.n10 585
R1008 VDD1.n42 VDD1.n41 585
R1009 VDD1.n39 VDD1.n38 585
R1010 VDD1.n48 VDD1.n47 585
R1011 VDD1.n50 VDD1.n49 585
R1012 VDD1.n35 VDD1.n34 585
R1013 VDD1.n56 VDD1.n55 585
R1014 VDD1.n58 VDD1.n57 585
R1015 VDD1.t0 VDD1.n9 327.601
R1016 VDD1.t1 VDD1.n40 327.601
R1017 VDD1.n26 VDD1.n25 171.744
R1018 VDD1.n25 VDD1.n3 171.744
R1019 VDD1.n18 VDD1.n3 171.744
R1020 VDD1.n18 VDD1.n17 171.744
R1021 VDD1.n17 VDD1.n7 171.744
R1022 VDD1.n10 VDD1.n7 171.744
R1023 VDD1.n41 VDD1.n38 171.744
R1024 VDD1.n48 VDD1.n38 171.744
R1025 VDD1.n49 VDD1.n48 171.744
R1026 VDD1.n49 VDD1.n34 171.744
R1027 VDD1.n56 VDD1.n34 171.744
R1028 VDD1.n57 VDD1.n56 171.744
R1029 VDD1.n10 VDD1.t0 85.8723
R1030 VDD1.n41 VDD1.t1 85.8723
R1031 VDD1 VDD1.n61 83.8696
R1032 VDD1 VDD1.n30 48.8642
R1033 VDD1.n11 VDD1.n9 16.3865
R1034 VDD1.n42 VDD1.n40 16.3865
R1035 VDD1.n12 VDD1.n8 12.8005
R1036 VDD1.n43 VDD1.n39 12.8005
R1037 VDD1.n16 VDD1.n15 12.0247
R1038 VDD1.n47 VDD1.n46 12.0247
R1039 VDD1.n19 VDD1.n6 11.249
R1040 VDD1.n50 VDD1.n37 11.249
R1041 VDD1.n20 VDD1.n4 10.4732
R1042 VDD1.n51 VDD1.n35 10.4732
R1043 VDD1.n24 VDD1.n23 9.69747
R1044 VDD1.n55 VDD1.n54 9.69747
R1045 VDD1.n30 VDD1.n29 9.45567
R1046 VDD1.n61 VDD1.n60 9.45567
R1047 VDD1.n29 VDD1.n28 9.3005
R1048 VDD1.n2 VDD1.n1 9.3005
R1049 VDD1.n23 VDD1.n22 9.3005
R1050 VDD1.n21 VDD1.n20 9.3005
R1051 VDD1.n6 VDD1.n5 9.3005
R1052 VDD1.n15 VDD1.n14 9.3005
R1053 VDD1.n13 VDD1.n12 9.3005
R1054 VDD1.n60 VDD1.n59 9.3005
R1055 VDD1.n33 VDD1.n32 9.3005
R1056 VDD1.n54 VDD1.n53 9.3005
R1057 VDD1.n52 VDD1.n51 9.3005
R1058 VDD1.n37 VDD1.n36 9.3005
R1059 VDD1.n46 VDD1.n45 9.3005
R1060 VDD1.n44 VDD1.n43 9.3005
R1061 VDD1.n27 VDD1.n2 8.92171
R1062 VDD1.n58 VDD1.n33 8.92171
R1063 VDD1.n28 VDD1.n0 8.14595
R1064 VDD1.n59 VDD1.n31 8.14595
R1065 VDD1.n30 VDD1.n0 5.81868
R1066 VDD1.n61 VDD1.n31 5.81868
R1067 VDD1.n28 VDD1.n27 5.04292
R1068 VDD1.n59 VDD1.n58 5.04292
R1069 VDD1.n24 VDD1.n2 4.26717
R1070 VDD1.n55 VDD1.n33 4.26717
R1071 VDD1.n13 VDD1.n9 3.71286
R1072 VDD1.n44 VDD1.n40 3.71286
R1073 VDD1.n23 VDD1.n4 3.49141
R1074 VDD1.n54 VDD1.n35 3.49141
R1075 VDD1.n20 VDD1.n19 2.71565
R1076 VDD1.n51 VDD1.n50 2.71565
R1077 VDD1.n16 VDD1.n6 1.93989
R1078 VDD1.n47 VDD1.n37 1.93989
R1079 VDD1.n15 VDD1.n8 1.16414
R1080 VDD1.n46 VDD1.n39 1.16414
R1081 VDD1.n12 VDD1.n11 0.388379
R1082 VDD1.n43 VDD1.n42 0.388379
R1083 VDD1.n29 VDD1.n1 0.155672
R1084 VDD1.n22 VDD1.n1 0.155672
R1085 VDD1.n22 VDD1.n21 0.155672
R1086 VDD1.n21 VDD1.n5 0.155672
R1087 VDD1.n14 VDD1.n5 0.155672
R1088 VDD1.n14 VDD1.n13 0.155672
R1089 VDD1.n45 VDD1.n44 0.155672
R1090 VDD1.n45 VDD1.n36 0.155672
R1091 VDD1.n52 VDD1.n36 0.155672
R1092 VDD1.n53 VDD1.n52 0.155672
R1093 VDD1.n53 VDD1.n32 0.155672
R1094 VDD1.n60 VDD1.n32 0.155672
C0 VDD2 VN 1.53949f
C1 VDD1 B 1.27811f
C2 w_n2302_n2160# VDD2 1.43982f
C3 w_n2302_n2160# VN 3.09907f
C4 VTAIL VDD2 3.63032f
C5 VTAIL VN 1.60743f
C6 w_n2302_n2160# VTAIL 1.91258f
C7 VDD2 VP 0.349767f
C8 VP VN 4.52008f
C9 w_n2302_n2160# VP 3.39316f
C10 VDD1 VDD2 0.722532f
C11 VDD1 VN 0.14864f
C12 w_n2302_n2160# VDD1 1.409f
C13 VTAIL VP 1.62161f
C14 VDD2 B 1.31175f
C15 VDD1 VTAIL 3.57542f
C16 VN B 1.04505f
C17 w_n2302_n2160# B 7.55991f
C18 VTAIL B 2.41226f
C19 VDD1 VP 1.7392f
C20 VP B 1.53016f
C21 VDD2 VSUBS 0.689172f
C22 VDD1 VSUBS 2.436873f
C23 VTAIL VSUBS 0.551785f
C24 VN VSUBS 5.50597f
C25 VP VSUBS 1.460014f
C26 B VSUBS 3.693032f
C27 w_n2302_n2160# VSUBS 62.071102f
C28 VDD1.n0 VSUBS 0.015637f
C29 VDD1.n1 VSUBS 0.01451f
C30 VDD1.n2 VSUBS 0.007797f
C31 VDD1.n3 VSUBS 0.018429f
C32 VDD1.n4 VSUBS 0.008256f
C33 VDD1.n5 VSUBS 0.01451f
C34 VDD1.n6 VSUBS 0.007797f
C35 VDD1.n7 VSUBS 0.018429f
C36 VDD1.n8 VSUBS 0.008256f
C37 VDD1.n9 VSUBS 0.063953f
C38 VDD1.t0 VSUBS 0.039512f
C39 VDD1.n10 VSUBS 0.013822f
C40 VDD1.n11 VSUBS 0.011718f
C41 VDD1.n12 VSUBS 0.007797f
C42 VDD1.n13 VSUBS 0.330277f
C43 VDD1.n14 VSUBS 0.01451f
C44 VDD1.n15 VSUBS 0.007797f
C45 VDD1.n16 VSUBS 0.008256f
C46 VDD1.n17 VSUBS 0.018429f
C47 VDD1.n18 VSUBS 0.018429f
C48 VDD1.n19 VSUBS 0.008256f
C49 VDD1.n20 VSUBS 0.007797f
C50 VDD1.n21 VSUBS 0.01451f
C51 VDD1.n22 VSUBS 0.01451f
C52 VDD1.n23 VSUBS 0.007797f
C53 VDD1.n24 VSUBS 0.008256f
C54 VDD1.n25 VSUBS 0.018429f
C55 VDD1.n26 VSUBS 0.043571f
C56 VDD1.n27 VSUBS 0.008256f
C57 VDD1.n28 VSUBS 0.007797f
C58 VDD1.n29 VSUBS 0.032746f
C59 VDD1.n30 VSUBS 0.032878f
C60 VDD1.n31 VSUBS 0.015637f
C61 VDD1.n32 VSUBS 0.01451f
C62 VDD1.n33 VSUBS 0.007797f
C63 VDD1.n34 VSUBS 0.018429f
C64 VDD1.n35 VSUBS 0.008256f
C65 VDD1.n36 VSUBS 0.01451f
C66 VDD1.n37 VSUBS 0.007797f
C67 VDD1.n38 VSUBS 0.018429f
C68 VDD1.n39 VSUBS 0.008256f
C69 VDD1.n40 VSUBS 0.063953f
C70 VDD1.t1 VSUBS 0.039512f
C71 VDD1.n41 VSUBS 0.013822f
C72 VDD1.n42 VSUBS 0.011718f
C73 VDD1.n43 VSUBS 0.007797f
C74 VDD1.n44 VSUBS 0.330277f
C75 VDD1.n45 VSUBS 0.01451f
C76 VDD1.n46 VSUBS 0.007797f
C77 VDD1.n47 VSUBS 0.008256f
C78 VDD1.n48 VSUBS 0.018429f
C79 VDD1.n49 VSUBS 0.018429f
C80 VDD1.n50 VSUBS 0.008256f
C81 VDD1.n51 VSUBS 0.007797f
C82 VDD1.n52 VSUBS 0.01451f
C83 VDD1.n53 VSUBS 0.01451f
C84 VDD1.n54 VSUBS 0.007797f
C85 VDD1.n55 VSUBS 0.008256f
C86 VDD1.n56 VSUBS 0.018429f
C87 VDD1.n57 VSUBS 0.043571f
C88 VDD1.n58 VSUBS 0.008256f
C89 VDD1.n59 VSUBS 0.007797f
C90 VDD1.n60 VSUBS 0.032746f
C91 VDD1.n61 VSUBS 0.352875f
C92 VP.t0 VSUBS 1.96494f
C93 VP.t1 VSUBS 2.58778f
C94 VP.n0 VSUBS 3.24792f
C95 VDD2.n0 VSUBS 0.015873f
C96 VDD2.n1 VSUBS 0.014729f
C97 VDD2.n2 VSUBS 0.007915f
C98 VDD2.n3 VSUBS 0.018708f
C99 VDD2.n4 VSUBS 0.00838f
C100 VDD2.n5 VSUBS 0.014729f
C101 VDD2.n6 VSUBS 0.007915f
C102 VDD2.n7 VSUBS 0.018708f
C103 VDD2.n8 VSUBS 0.00838f
C104 VDD2.n9 VSUBS 0.06492f
C105 VDD2.t1 VSUBS 0.040109f
C106 VDD2.n10 VSUBS 0.014031f
C107 VDD2.n11 VSUBS 0.011895f
C108 VDD2.n12 VSUBS 0.007915f
C109 VDD2.n13 VSUBS 0.335268f
C110 VDD2.n14 VSUBS 0.014729f
C111 VDD2.n15 VSUBS 0.007915f
C112 VDD2.n16 VSUBS 0.00838f
C113 VDD2.n17 VSUBS 0.018708f
C114 VDD2.n18 VSUBS 0.018708f
C115 VDD2.n19 VSUBS 0.00838f
C116 VDD2.n20 VSUBS 0.007915f
C117 VDD2.n21 VSUBS 0.014729f
C118 VDD2.n22 VSUBS 0.014729f
C119 VDD2.n23 VSUBS 0.007915f
C120 VDD2.n24 VSUBS 0.00838f
C121 VDD2.n25 VSUBS 0.018708f
C122 VDD2.n26 VSUBS 0.044229f
C123 VDD2.n27 VSUBS 0.00838f
C124 VDD2.n28 VSUBS 0.007915f
C125 VDD2.n29 VSUBS 0.033241f
C126 VDD2.n30 VSUBS 0.330517f
C127 VDD2.n31 VSUBS 0.015873f
C128 VDD2.n32 VSUBS 0.014729f
C129 VDD2.n33 VSUBS 0.007915f
C130 VDD2.n34 VSUBS 0.018708f
C131 VDD2.n35 VSUBS 0.00838f
C132 VDD2.n36 VSUBS 0.014729f
C133 VDD2.n37 VSUBS 0.007915f
C134 VDD2.n38 VSUBS 0.018708f
C135 VDD2.n39 VSUBS 0.00838f
C136 VDD2.n40 VSUBS 0.06492f
C137 VDD2.t0 VSUBS 0.040109f
C138 VDD2.n41 VSUBS 0.014031f
C139 VDD2.n42 VSUBS 0.011895f
C140 VDD2.n43 VSUBS 0.007915f
C141 VDD2.n44 VSUBS 0.335268f
C142 VDD2.n45 VSUBS 0.014729f
C143 VDD2.n46 VSUBS 0.007915f
C144 VDD2.n47 VSUBS 0.00838f
C145 VDD2.n48 VSUBS 0.018708f
C146 VDD2.n49 VSUBS 0.018708f
C147 VDD2.n50 VSUBS 0.00838f
C148 VDD2.n51 VSUBS 0.007915f
C149 VDD2.n52 VSUBS 0.014729f
C150 VDD2.n53 VSUBS 0.014729f
C151 VDD2.n54 VSUBS 0.007915f
C152 VDD2.n55 VSUBS 0.00838f
C153 VDD2.n56 VSUBS 0.018708f
C154 VDD2.n57 VSUBS 0.044229f
C155 VDD2.n58 VSUBS 0.00838f
C156 VDD2.n59 VSUBS 0.007915f
C157 VDD2.n60 VSUBS 0.033241f
C158 VDD2.n61 VSUBS 0.032347f
C159 VDD2.n62 VSUBS 1.4669f
C160 VTAIL.n0 VSUBS 0.023729f
C161 VTAIL.n1 VSUBS 0.022019f
C162 VTAIL.n2 VSUBS 0.011832f
C163 VTAIL.n3 VSUBS 0.027966f
C164 VTAIL.n4 VSUBS 0.012528f
C165 VTAIL.n5 VSUBS 0.022019f
C166 VTAIL.n6 VSUBS 0.011832f
C167 VTAIL.n7 VSUBS 0.027966f
C168 VTAIL.n8 VSUBS 0.012528f
C169 VTAIL.n9 VSUBS 0.097049f
C170 VTAIL.t1 VSUBS 0.059959f
C171 VTAIL.n10 VSUBS 0.020975f
C172 VTAIL.n11 VSUBS 0.017781f
C173 VTAIL.n12 VSUBS 0.011832f
C174 VTAIL.n13 VSUBS 0.501193f
C175 VTAIL.n14 VSUBS 0.022019f
C176 VTAIL.n15 VSUBS 0.011832f
C177 VTAIL.n16 VSUBS 0.012528f
C178 VTAIL.n17 VSUBS 0.027966f
C179 VTAIL.n18 VSUBS 0.027966f
C180 VTAIL.n19 VSUBS 0.012528f
C181 VTAIL.n20 VSUBS 0.011832f
C182 VTAIL.n21 VSUBS 0.022019f
C183 VTAIL.n22 VSUBS 0.022019f
C184 VTAIL.n23 VSUBS 0.011832f
C185 VTAIL.n24 VSUBS 0.012528f
C186 VTAIL.n25 VSUBS 0.027966f
C187 VTAIL.n26 VSUBS 0.066118f
C188 VTAIL.n27 VSUBS 0.012528f
C189 VTAIL.n28 VSUBS 0.011832f
C190 VTAIL.n29 VSUBS 0.049692f
C191 VTAIL.n30 VSUBS 0.033143f
C192 VTAIL.n31 VSUBS 1.17749f
C193 VTAIL.n32 VSUBS 0.023729f
C194 VTAIL.n33 VSUBS 0.022019f
C195 VTAIL.n34 VSUBS 0.011832f
C196 VTAIL.n35 VSUBS 0.027966f
C197 VTAIL.n36 VSUBS 0.012528f
C198 VTAIL.n37 VSUBS 0.022019f
C199 VTAIL.n38 VSUBS 0.011832f
C200 VTAIL.n39 VSUBS 0.027966f
C201 VTAIL.n40 VSUBS 0.012528f
C202 VTAIL.n41 VSUBS 0.097049f
C203 VTAIL.t2 VSUBS 0.059959f
C204 VTAIL.n42 VSUBS 0.020975f
C205 VTAIL.n43 VSUBS 0.017781f
C206 VTAIL.n44 VSUBS 0.011832f
C207 VTAIL.n45 VSUBS 0.501193f
C208 VTAIL.n46 VSUBS 0.022019f
C209 VTAIL.n47 VSUBS 0.011832f
C210 VTAIL.n48 VSUBS 0.012528f
C211 VTAIL.n49 VSUBS 0.027966f
C212 VTAIL.n50 VSUBS 0.027966f
C213 VTAIL.n51 VSUBS 0.012528f
C214 VTAIL.n52 VSUBS 0.011832f
C215 VTAIL.n53 VSUBS 0.022019f
C216 VTAIL.n54 VSUBS 0.022019f
C217 VTAIL.n55 VSUBS 0.011832f
C218 VTAIL.n56 VSUBS 0.012528f
C219 VTAIL.n57 VSUBS 0.027966f
C220 VTAIL.n58 VSUBS 0.066118f
C221 VTAIL.n59 VSUBS 0.012528f
C222 VTAIL.n60 VSUBS 0.011832f
C223 VTAIL.n61 VSUBS 0.049692f
C224 VTAIL.n62 VSUBS 0.033143f
C225 VTAIL.n63 VSUBS 1.22428f
C226 VTAIL.n64 VSUBS 0.023729f
C227 VTAIL.n65 VSUBS 0.022019f
C228 VTAIL.n66 VSUBS 0.011832f
C229 VTAIL.n67 VSUBS 0.027966f
C230 VTAIL.n68 VSUBS 0.012528f
C231 VTAIL.n69 VSUBS 0.022019f
C232 VTAIL.n70 VSUBS 0.011832f
C233 VTAIL.n71 VSUBS 0.027966f
C234 VTAIL.n72 VSUBS 0.012528f
C235 VTAIL.n73 VSUBS 0.097049f
C236 VTAIL.t0 VSUBS 0.059959f
C237 VTAIL.n74 VSUBS 0.020975f
C238 VTAIL.n75 VSUBS 0.017781f
C239 VTAIL.n76 VSUBS 0.011832f
C240 VTAIL.n77 VSUBS 0.501193f
C241 VTAIL.n78 VSUBS 0.022019f
C242 VTAIL.n79 VSUBS 0.011832f
C243 VTAIL.n80 VSUBS 0.012528f
C244 VTAIL.n81 VSUBS 0.027966f
C245 VTAIL.n82 VSUBS 0.027966f
C246 VTAIL.n83 VSUBS 0.012528f
C247 VTAIL.n84 VSUBS 0.011832f
C248 VTAIL.n85 VSUBS 0.022019f
C249 VTAIL.n86 VSUBS 0.022019f
C250 VTAIL.n87 VSUBS 0.011832f
C251 VTAIL.n88 VSUBS 0.012528f
C252 VTAIL.n89 VSUBS 0.027966f
C253 VTAIL.n90 VSUBS 0.066118f
C254 VTAIL.n91 VSUBS 0.012528f
C255 VTAIL.n92 VSUBS 0.011832f
C256 VTAIL.n93 VSUBS 0.049692f
C257 VTAIL.n94 VSUBS 0.033143f
C258 VTAIL.n95 VSUBS 1.02061f
C259 VTAIL.n96 VSUBS 0.023729f
C260 VTAIL.n97 VSUBS 0.022019f
C261 VTAIL.n98 VSUBS 0.011832f
C262 VTAIL.n99 VSUBS 0.027966f
C263 VTAIL.n100 VSUBS 0.012528f
C264 VTAIL.n101 VSUBS 0.022019f
C265 VTAIL.n102 VSUBS 0.011832f
C266 VTAIL.n103 VSUBS 0.027966f
C267 VTAIL.n104 VSUBS 0.012528f
C268 VTAIL.n105 VSUBS 0.097049f
C269 VTAIL.t3 VSUBS 0.059959f
C270 VTAIL.n106 VSUBS 0.020975f
C271 VTAIL.n107 VSUBS 0.017781f
C272 VTAIL.n108 VSUBS 0.011832f
C273 VTAIL.n109 VSUBS 0.501193f
C274 VTAIL.n110 VSUBS 0.022019f
C275 VTAIL.n111 VSUBS 0.011832f
C276 VTAIL.n112 VSUBS 0.012528f
C277 VTAIL.n113 VSUBS 0.027966f
C278 VTAIL.n114 VSUBS 0.027966f
C279 VTAIL.n115 VSUBS 0.012528f
C280 VTAIL.n116 VSUBS 0.011832f
C281 VTAIL.n117 VSUBS 0.022019f
C282 VTAIL.n118 VSUBS 0.022019f
C283 VTAIL.n119 VSUBS 0.011832f
C284 VTAIL.n120 VSUBS 0.012528f
C285 VTAIL.n121 VSUBS 0.027966f
C286 VTAIL.n122 VSUBS 0.066118f
C287 VTAIL.n123 VSUBS 0.012528f
C288 VTAIL.n124 VSUBS 0.011832f
C289 VTAIL.n125 VSUBS 0.049692f
C290 VTAIL.n126 VSUBS 0.033143f
C291 VTAIL.n127 VSUBS 0.932225f
C292 VN.t0 VSUBS 1.88206f
C293 VN.t1 VSUBS 2.47755f
C294 B.n0 VSUBS 0.006826f
C295 B.n1 VSUBS 0.006826f
C296 B.n2 VSUBS 0.010096f
C297 B.n3 VSUBS 0.007736f
C298 B.n4 VSUBS 0.007736f
C299 B.n5 VSUBS 0.007736f
C300 B.n6 VSUBS 0.007736f
C301 B.n7 VSUBS 0.007736f
C302 B.n8 VSUBS 0.007736f
C303 B.n9 VSUBS 0.007736f
C304 B.n10 VSUBS 0.007736f
C305 B.n11 VSUBS 0.007736f
C306 B.n12 VSUBS 0.007736f
C307 B.n13 VSUBS 0.007736f
C308 B.n14 VSUBS 0.007736f
C309 B.n15 VSUBS 0.018907f
C310 B.n16 VSUBS 0.007736f
C311 B.n17 VSUBS 0.007736f
C312 B.n18 VSUBS 0.007736f
C313 B.n19 VSUBS 0.007736f
C314 B.n20 VSUBS 0.007736f
C315 B.n21 VSUBS 0.007736f
C316 B.n22 VSUBS 0.007736f
C317 B.n23 VSUBS 0.007736f
C318 B.n24 VSUBS 0.007736f
C319 B.n25 VSUBS 0.007736f
C320 B.n26 VSUBS 0.007736f
C321 B.n27 VSUBS 0.007736f
C322 B.t10 VSUBS 0.09805f
C323 B.t11 VSUBS 0.129747f
C324 B.t9 VSUBS 0.941145f
C325 B.n28 VSUBS 0.218931f
C326 B.n29 VSUBS 0.173981f
C327 B.n30 VSUBS 0.007736f
C328 B.n31 VSUBS 0.007736f
C329 B.n32 VSUBS 0.007736f
C330 B.n33 VSUBS 0.007736f
C331 B.t4 VSUBS 0.098052f
C332 B.t5 VSUBS 0.129749f
C333 B.t3 VSUBS 0.941145f
C334 B.n34 VSUBS 0.21893f
C335 B.n35 VSUBS 0.173979f
C336 B.n36 VSUBS 0.017924f
C337 B.n37 VSUBS 0.007736f
C338 B.n38 VSUBS 0.007736f
C339 B.n39 VSUBS 0.007736f
C340 B.n40 VSUBS 0.007736f
C341 B.n41 VSUBS 0.007736f
C342 B.n42 VSUBS 0.007736f
C343 B.n43 VSUBS 0.007736f
C344 B.n44 VSUBS 0.007736f
C345 B.n45 VSUBS 0.007736f
C346 B.n46 VSUBS 0.007736f
C347 B.n47 VSUBS 0.007736f
C348 B.n48 VSUBS 0.019775f
C349 B.n49 VSUBS 0.007736f
C350 B.n50 VSUBS 0.007736f
C351 B.n51 VSUBS 0.007736f
C352 B.n52 VSUBS 0.007736f
C353 B.n53 VSUBS 0.007736f
C354 B.n54 VSUBS 0.007736f
C355 B.n55 VSUBS 0.007736f
C356 B.n56 VSUBS 0.007736f
C357 B.n57 VSUBS 0.007736f
C358 B.n58 VSUBS 0.007736f
C359 B.n59 VSUBS 0.007736f
C360 B.n60 VSUBS 0.007736f
C361 B.n61 VSUBS 0.007736f
C362 B.n62 VSUBS 0.007736f
C363 B.n63 VSUBS 0.007736f
C364 B.n64 VSUBS 0.007736f
C365 B.n65 VSUBS 0.007736f
C366 B.n66 VSUBS 0.007736f
C367 B.n67 VSUBS 0.007736f
C368 B.n68 VSUBS 0.007736f
C369 B.n69 VSUBS 0.007736f
C370 B.n70 VSUBS 0.007736f
C371 B.n71 VSUBS 0.007736f
C372 B.n72 VSUBS 0.007736f
C373 B.n73 VSUBS 0.007736f
C374 B.n74 VSUBS 0.007736f
C375 B.n75 VSUBS 0.007736f
C376 B.n76 VSUBS 0.019735f
C377 B.n77 VSUBS 0.007736f
C378 B.n78 VSUBS 0.007736f
C379 B.n79 VSUBS 0.007736f
C380 B.n80 VSUBS 0.007736f
C381 B.n81 VSUBS 0.007736f
C382 B.n82 VSUBS 0.007736f
C383 B.n83 VSUBS 0.007736f
C384 B.n84 VSUBS 0.007736f
C385 B.n85 VSUBS 0.007736f
C386 B.n86 VSUBS 0.007736f
C387 B.n87 VSUBS 0.007736f
C388 B.n88 VSUBS 0.005347f
C389 B.n89 VSUBS 0.007736f
C390 B.n90 VSUBS 0.007736f
C391 B.n91 VSUBS 0.007736f
C392 B.n92 VSUBS 0.007736f
C393 B.n93 VSUBS 0.007736f
C394 B.t2 VSUBS 0.09805f
C395 B.t1 VSUBS 0.129747f
C396 B.t0 VSUBS 0.941145f
C397 B.n94 VSUBS 0.218931f
C398 B.n95 VSUBS 0.173981f
C399 B.n96 VSUBS 0.007736f
C400 B.n97 VSUBS 0.007736f
C401 B.n98 VSUBS 0.007736f
C402 B.n99 VSUBS 0.007736f
C403 B.n100 VSUBS 0.007736f
C404 B.n101 VSUBS 0.007736f
C405 B.n102 VSUBS 0.007736f
C406 B.n103 VSUBS 0.007736f
C407 B.n104 VSUBS 0.007736f
C408 B.n105 VSUBS 0.007736f
C409 B.n106 VSUBS 0.007736f
C410 B.n107 VSUBS 0.018907f
C411 B.n108 VSUBS 0.007736f
C412 B.n109 VSUBS 0.007736f
C413 B.n110 VSUBS 0.007736f
C414 B.n111 VSUBS 0.007736f
C415 B.n112 VSUBS 0.007736f
C416 B.n113 VSUBS 0.007736f
C417 B.n114 VSUBS 0.007736f
C418 B.n115 VSUBS 0.007736f
C419 B.n116 VSUBS 0.007736f
C420 B.n117 VSUBS 0.007736f
C421 B.n118 VSUBS 0.007736f
C422 B.n119 VSUBS 0.007736f
C423 B.n120 VSUBS 0.007736f
C424 B.n121 VSUBS 0.007736f
C425 B.n122 VSUBS 0.007736f
C426 B.n123 VSUBS 0.007736f
C427 B.n124 VSUBS 0.007736f
C428 B.n125 VSUBS 0.007736f
C429 B.n126 VSUBS 0.007736f
C430 B.n127 VSUBS 0.007736f
C431 B.n128 VSUBS 0.007736f
C432 B.n129 VSUBS 0.007736f
C433 B.n130 VSUBS 0.007736f
C434 B.n131 VSUBS 0.007736f
C435 B.n132 VSUBS 0.007736f
C436 B.n133 VSUBS 0.007736f
C437 B.n134 VSUBS 0.007736f
C438 B.n135 VSUBS 0.007736f
C439 B.n136 VSUBS 0.007736f
C440 B.n137 VSUBS 0.007736f
C441 B.n138 VSUBS 0.007736f
C442 B.n139 VSUBS 0.007736f
C443 B.n140 VSUBS 0.007736f
C444 B.n141 VSUBS 0.007736f
C445 B.n142 VSUBS 0.007736f
C446 B.n143 VSUBS 0.007736f
C447 B.n144 VSUBS 0.007736f
C448 B.n145 VSUBS 0.007736f
C449 B.n146 VSUBS 0.007736f
C450 B.n147 VSUBS 0.007736f
C451 B.n148 VSUBS 0.007736f
C452 B.n149 VSUBS 0.007736f
C453 B.n150 VSUBS 0.007736f
C454 B.n151 VSUBS 0.007736f
C455 B.n152 VSUBS 0.007736f
C456 B.n153 VSUBS 0.007736f
C457 B.n154 VSUBS 0.007736f
C458 B.n155 VSUBS 0.007736f
C459 B.n156 VSUBS 0.007736f
C460 B.n157 VSUBS 0.007736f
C461 B.n158 VSUBS 0.018907f
C462 B.n159 VSUBS 0.019775f
C463 B.n160 VSUBS 0.019775f
C464 B.n161 VSUBS 0.007736f
C465 B.n162 VSUBS 0.007736f
C466 B.n163 VSUBS 0.007736f
C467 B.n164 VSUBS 0.007736f
C468 B.n165 VSUBS 0.007736f
C469 B.n166 VSUBS 0.007736f
C470 B.n167 VSUBS 0.007736f
C471 B.n168 VSUBS 0.007736f
C472 B.n169 VSUBS 0.007736f
C473 B.n170 VSUBS 0.007736f
C474 B.n171 VSUBS 0.007736f
C475 B.n172 VSUBS 0.007736f
C476 B.n173 VSUBS 0.007736f
C477 B.n174 VSUBS 0.007736f
C478 B.n175 VSUBS 0.007736f
C479 B.n176 VSUBS 0.007736f
C480 B.n177 VSUBS 0.007736f
C481 B.n178 VSUBS 0.007736f
C482 B.n179 VSUBS 0.007736f
C483 B.n180 VSUBS 0.007736f
C484 B.n181 VSUBS 0.007736f
C485 B.n182 VSUBS 0.007736f
C486 B.n183 VSUBS 0.007736f
C487 B.n184 VSUBS 0.007736f
C488 B.n185 VSUBS 0.007736f
C489 B.n186 VSUBS 0.007736f
C490 B.n187 VSUBS 0.007736f
C491 B.n188 VSUBS 0.007736f
C492 B.n189 VSUBS 0.007736f
C493 B.n190 VSUBS 0.007736f
C494 B.n191 VSUBS 0.007736f
C495 B.n192 VSUBS 0.007736f
C496 B.n193 VSUBS 0.007736f
C497 B.n194 VSUBS 0.005347f
C498 B.n195 VSUBS 0.017924f
C499 B.n196 VSUBS 0.006257f
C500 B.n197 VSUBS 0.007736f
C501 B.n198 VSUBS 0.007736f
C502 B.n199 VSUBS 0.007736f
C503 B.n200 VSUBS 0.007736f
C504 B.n201 VSUBS 0.007736f
C505 B.n202 VSUBS 0.007736f
C506 B.n203 VSUBS 0.007736f
C507 B.n204 VSUBS 0.007736f
C508 B.n205 VSUBS 0.007736f
C509 B.n206 VSUBS 0.007736f
C510 B.n207 VSUBS 0.007736f
C511 B.t8 VSUBS 0.098052f
C512 B.t7 VSUBS 0.129749f
C513 B.t6 VSUBS 0.941145f
C514 B.n208 VSUBS 0.21893f
C515 B.n209 VSUBS 0.173979f
C516 B.n210 VSUBS 0.017924f
C517 B.n211 VSUBS 0.006257f
C518 B.n212 VSUBS 0.007736f
C519 B.n213 VSUBS 0.007736f
C520 B.n214 VSUBS 0.007736f
C521 B.n215 VSUBS 0.007736f
C522 B.n216 VSUBS 0.007736f
C523 B.n217 VSUBS 0.007736f
C524 B.n218 VSUBS 0.007736f
C525 B.n219 VSUBS 0.007736f
C526 B.n220 VSUBS 0.007736f
C527 B.n221 VSUBS 0.007736f
C528 B.n222 VSUBS 0.007736f
C529 B.n223 VSUBS 0.007736f
C530 B.n224 VSUBS 0.007736f
C531 B.n225 VSUBS 0.007736f
C532 B.n226 VSUBS 0.007736f
C533 B.n227 VSUBS 0.007736f
C534 B.n228 VSUBS 0.007736f
C535 B.n229 VSUBS 0.007736f
C536 B.n230 VSUBS 0.007736f
C537 B.n231 VSUBS 0.007736f
C538 B.n232 VSUBS 0.007736f
C539 B.n233 VSUBS 0.007736f
C540 B.n234 VSUBS 0.007736f
C541 B.n235 VSUBS 0.007736f
C542 B.n236 VSUBS 0.007736f
C543 B.n237 VSUBS 0.007736f
C544 B.n238 VSUBS 0.007736f
C545 B.n239 VSUBS 0.007736f
C546 B.n240 VSUBS 0.007736f
C547 B.n241 VSUBS 0.007736f
C548 B.n242 VSUBS 0.007736f
C549 B.n243 VSUBS 0.007736f
C550 B.n244 VSUBS 0.007736f
C551 B.n245 VSUBS 0.007736f
C552 B.n246 VSUBS 0.007736f
C553 B.n247 VSUBS 0.018947f
C554 B.n248 VSUBS 0.019775f
C555 B.n249 VSUBS 0.018907f
C556 B.n250 VSUBS 0.007736f
C557 B.n251 VSUBS 0.007736f
C558 B.n252 VSUBS 0.007736f
C559 B.n253 VSUBS 0.007736f
C560 B.n254 VSUBS 0.007736f
C561 B.n255 VSUBS 0.007736f
C562 B.n256 VSUBS 0.007736f
C563 B.n257 VSUBS 0.007736f
C564 B.n258 VSUBS 0.007736f
C565 B.n259 VSUBS 0.007736f
C566 B.n260 VSUBS 0.007736f
C567 B.n261 VSUBS 0.007736f
C568 B.n262 VSUBS 0.007736f
C569 B.n263 VSUBS 0.007736f
C570 B.n264 VSUBS 0.007736f
C571 B.n265 VSUBS 0.007736f
C572 B.n266 VSUBS 0.007736f
C573 B.n267 VSUBS 0.007736f
C574 B.n268 VSUBS 0.007736f
C575 B.n269 VSUBS 0.007736f
C576 B.n270 VSUBS 0.007736f
C577 B.n271 VSUBS 0.007736f
C578 B.n272 VSUBS 0.007736f
C579 B.n273 VSUBS 0.007736f
C580 B.n274 VSUBS 0.007736f
C581 B.n275 VSUBS 0.007736f
C582 B.n276 VSUBS 0.007736f
C583 B.n277 VSUBS 0.007736f
C584 B.n278 VSUBS 0.007736f
C585 B.n279 VSUBS 0.007736f
C586 B.n280 VSUBS 0.007736f
C587 B.n281 VSUBS 0.007736f
C588 B.n282 VSUBS 0.007736f
C589 B.n283 VSUBS 0.007736f
C590 B.n284 VSUBS 0.007736f
C591 B.n285 VSUBS 0.007736f
C592 B.n286 VSUBS 0.007736f
C593 B.n287 VSUBS 0.007736f
C594 B.n288 VSUBS 0.007736f
C595 B.n289 VSUBS 0.007736f
C596 B.n290 VSUBS 0.007736f
C597 B.n291 VSUBS 0.007736f
C598 B.n292 VSUBS 0.007736f
C599 B.n293 VSUBS 0.007736f
C600 B.n294 VSUBS 0.007736f
C601 B.n295 VSUBS 0.007736f
C602 B.n296 VSUBS 0.007736f
C603 B.n297 VSUBS 0.007736f
C604 B.n298 VSUBS 0.007736f
C605 B.n299 VSUBS 0.007736f
C606 B.n300 VSUBS 0.007736f
C607 B.n301 VSUBS 0.007736f
C608 B.n302 VSUBS 0.007736f
C609 B.n303 VSUBS 0.007736f
C610 B.n304 VSUBS 0.007736f
C611 B.n305 VSUBS 0.007736f
C612 B.n306 VSUBS 0.007736f
C613 B.n307 VSUBS 0.007736f
C614 B.n308 VSUBS 0.007736f
C615 B.n309 VSUBS 0.007736f
C616 B.n310 VSUBS 0.007736f
C617 B.n311 VSUBS 0.007736f
C618 B.n312 VSUBS 0.007736f
C619 B.n313 VSUBS 0.007736f
C620 B.n314 VSUBS 0.007736f
C621 B.n315 VSUBS 0.007736f
C622 B.n316 VSUBS 0.007736f
C623 B.n317 VSUBS 0.007736f
C624 B.n318 VSUBS 0.007736f
C625 B.n319 VSUBS 0.007736f
C626 B.n320 VSUBS 0.007736f
C627 B.n321 VSUBS 0.007736f
C628 B.n322 VSUBS 0.007736f
C629 B.n323 VSUBS 0.007736f
C630 B.n324 VSUBS 0.007736f
C631 B.n325 VSUBS 0.007736f
C632 B.n326 VSUBS 0.007736f
C633 B.n327 VSUBS 0.007736f
C634 B.n328 VSUBS 0.007736f
C635 B.n329 VSUBS 0.007736f
C636 B.n330 VSUBS 0.007736f
C637 B.n331 VSUBS 0.018907f
C638 B.n332 VSUBS 0.018907f
C639 B.n333 VSUBS 0.019775f
C640 B.n334 VSUBS 0.007736f
C641 B.n335 VSUBS 0.007736f
C642 B.n336 VSUBS 0.007736f
C643 B.n337 VSUBS 0.007736f
C644 B.n338 VSUBS 0.007736f
C645 B.n339 VSUBS 0.007736f
C646 B.n340 VSUBS 0.007736f
C647 B.n341 VSUBS 0.007736f
C648 B.n342 VSUBS 0.007736f
C649 B.n343 VSUBS 0.007736f
C650 B.n344 VSUBS 0.007736f
C651 B.n345 VSUBS 0.007736f
C652 B.n346 VSUBS 0.007736f
C653 B.n347 VSUBS 0.007736f
C654 B.n348 VSUBS 0.007736f
C655 B.n349 VSUBS 0.007736f
C656 B.n350 VSUBS 0.007736f
C657 B.n351 VSUBS 0.007736f
C658 B.n352 VSUBS 0.007736f
C659 B.n353 VSUBS 0.007736f
C660 B.n354 VSUBS 0.007736f
C661 B.n355 VSUBS 0.007736f
C662 B.n356 VSUBS 0.007736f
C663 B.n357 VSUBS 0.007736f
C664 B.n358 VSUBS 0.007736f
C665 B.n359 VSUBS 0.007736f
C666 B.n360 VSUBS 0.007736f
C667 B.n361 VSUBS 0.007736f
C668 B.n362 VSUBS 0.007736f
C669 B.n363 VSUBS 0.007736f
C670 B.n364 VSUBS 0.007736f
C671 B.n365 VSUBS 0.007736f
C672 B.n366 VSUBS 0.007736f
C673 B.n367 VSUBS 0.005347f
C674 B.n368 VSUBS 0.007736f
C675 B.n369 VSUBS 0.007736f
C676 B.n370 VSUBS 0.006257f
C677 B.n371 VSUBS 0.007736f
C678 B.n372 VSUBS 0.007736f
C679 B.n373 VSUBS 0.007736f
C680 B.n374 VSUBS 0.007736f
C681 B.n375 VSUBS 0.007736f
C682 B.n376 VSUBS 0.007736f
C683 B.n377 VSUBS 0.007736f
C684 B.n378 VSUBS 0.007736f
C685 B.n379 VSUBS 0.007736f
C686 B.n380 VSUBS 0.007736f
C687 B.n381 VSUBS 0.007736f
C688 B.n382 VSUBS 0.006257f
C689 B.n383 VSUBS 0.017924f
C690 B.n384 VSUBS 0.005347f
C691 B.n385 VSUBS 0.007736f
C692 B.n386 VSUBS 0.007736f
C693 B.n387 VSUBS 0.007736f
C694 B.n388 VSUBS 0.007736f
C695 B.n389 VSUBS 0.007736f
C696 B.n390 VSUBS 0.007736f
C697 B.n391 VSUBS 0.007736f
C698 B.n392 VSUBS 0.007736f
C699 B.n393 VSUBS 0.007736f
C700 B.n394 VSUBS 0.007736f
C701 B.n395 VSUBS 0.007736f
C702 B.n396 VSUBS 0.007736f
C703 B.n397 VSUBS 0.007736f
C704 B.n398 VSUBS 0.007736f
C705 B.n399 VSUBS 0.007736f
C706 B.n400 VSUBS 0.007736f
C707 B.n401 VSUBS 0.007736f
C708 B.n402 VSUBS 0.007736f
C709 B.n403 VSUBS 0.007736f
C710 B.n404 VSUBS 0.007736f
C711 B.n405 VSUBS 0.007736f
C712 B.n406 VSUBS 0.007736f
C713 B.n407 VSUBS 0.007736f
C714 B.n408 VSUBS 0.007736f
C715 B.n409 VSUBS 0.007736f
C716 B.n410 VSUBS 0.007736f
C717 B.n411 VSUBS 0.007736f
C718 B.n412 VSUBS 0.007736f
C719 B.n413 VSUBS 0.007736f
C720 B.n414 VSUBS 0.007736f
C721 B.n415 VSUBS 0.007736f
C722 B.n416 VSUBS 0.007736f
C723 B.n417 VSUBS 0.007736f
C724 B.n418 VSUBS 0.019775f
C725 B.n419 VSUBS 0.019775f
C726 B.n420 VSUBS 0.018907f
C727 B.n421 VSUBS 0.007736f
C728 B.n422 VSUBS 0.007736f
C729 B.n423 VSUBS 0.007736f
C730 B.n424 VSUBS 0.007736f
C731 B.n425 VSUBS 0.007736f
C732 B.n426 VSUBS 0.007736f
C733 B.n427 VSUBS 0.007736f
C734 B.n428 VSUBS 0.007736f
C735 B.n429 VSUBS 0.007736f
C736 B.n430 VSUBS 0.007736f
C737 B.n431 VSUBS 0.007736f
C738 B.n432 VSUBS 0.007736f
C739 B.n433 VSUBS 0.007736f
C740 B.n434 VSUBS 0.007736f
C741 B.n435 VSUBS 0.007736f
C742 B.n436 VSUBS 0.007736f
C743 B.n437 VSUBS 0.007736f
C744 B.n438 VSUBS 0.007736f
C745 B.n439 VSUBS 0.007736f
C746 B.n440 VSUBS 0.007736f
C747 B.n441 VSUBS 0.007736f
C748 B.n442 VSUBS 0.007736f
C749 B.n443 VSUBS 0.007736f
C750 B.n444 VSUBS 0.007736f
C751 B.n445 VSUBS 0.007736f
C752 B.n446 VSUBS 0.007736f
C753 B.n447 VSUBS 0.007736f
C754 B.n448 VSUBS 0.007736f
C755 B.n449 VSUBS 0.007736f
C756 B.n450 VSUBS 0.007736f
C757 B.n451 VSUBS 0.007736f
C758 B.n452 VSUBS 0.007736f
C759 B.n453 VSUBS 0.007736f
C760 B.n454 VSUBS 0.007736f
C761 B.n455 VSUBS 0.007736f
C762 B.n456 VSUBS 0.007736f
C763 B.n457 VSUBS 0.007736f
C764 B.n458 VSUBS 0.007736f
C765 B.n459 VSUBS 0.010096f
C766 B.n460 VSUBS 0.010754f
C767 B.n461 VSUBS 0.021386f
.ends

