* NGSPICE file created from diff_pair_sample_1285.ext - technology: sky130A

.subckt diff_pair_sample_1285 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t3 VP.t0 VTAIL.t5 w_n2230_n1808# sky130_fd_pr__pfet_01v8 ad=0.693 pd=4.53 as=1.638 ps=9.18 w=4.2 l=1.77
X1 B.t11 B.t9 B.t10 w_n2230_n1808# sky130_fd_pr__pfet_01v8 ad=1.638 pd=9.18 as=0 ps=0 w=4.2 l=1.77
X2 VDD2.t3 VN.t0 VTAIL.t1 w_n2230_n1808# sky130_fd_pr__pfet_01v8 ad=0.693 pd=4.53 as=1.638 ps=9.18 w=4.2 l=1.77
X3 B.t8 B.t6 B.t7 w_n2230_n1808# sky130_fd_pr__pfet_01v8 ad=1.638 pd=9.18 as=0 ps=0 w=4.2 l=1.77
X4 VTAIL.t6 VP.t1 VDD1.t2 w_n2230_n1808# sky130_fd_pr__pfet_01v8 ad=1.638 pd=9.18 as=0.693 ps=4.53 w=4.2 l=1.77
X5 VDD1.t1 VP.t2 VTAIL.t7 w_n2230_n1808# sky130_fd_pr__pfet_01v8 ad=0.693 pd=4.53 as=1.638 ps=9.18 w=4.2 l=1.77
X6 VDD2.t2 VN.t1 VTAIL.t2 w_n2230_n1808# sky130_fd_pr__pfet_01v8 ad=0.693 pd=4.53 as=1.638 ps=9.18 w=4.2 l=1.77
X7 B.t5 B.t3 B.t4 w_n2230_n1808# sky130_fd_pr__pfet_01v8 ad=1.638 pd=9.18 as=0 ps=0 w=4.2 l=1.77
X8 VTAIL.t3 VN.t2 VDD2.t1 w_n2230_n1808# sky130_fd_pr__pfet_01v8 ad=1.638 pd=9.18 as=0.693 ps=4.53 w=4.2 l=1.77
X9 VTAIL.t0 VN.t3 VDD2.t0 w_n2230_n1808# sky130_fd_pr__pfet_01v8 ad=1.638 pd=9.18 as=0.693 ps=4.53 w=4.2 l=1.77
X10 VTAIL.t4 VP.t3 VDD1.t0 w_n2230_n1808# sky130_fd_pr__pfet_01v8 ad=1.638 pd=9.18 as=0.693 ps=4.53 w=4.2 l=1.77
X11 B.t2 B.t0 B.t1 w_n2230_n1808# sky130_fd_pr__pfet_01v8 ad=1.638 pd=9.18 as=0 ps=0 w=4.2 l=1.77
R0 VP.n5 VP.n4 183.434
R1 VP.n14 VP.n13 183.434
R2 VP.n12 VP.n0 161.3
R3 VP.n11 VP.n10 161.3
R4 VP.n9 VP.n1 161.3
R5 VP.n8 VP.n7 161.3
R6 VP.n6 VP.n2 161.3
R7 VP.n3 VP.t3 93.3598
R8 VP.n3 VP.t2 92.9312
R9 VP.n5 VP.t1 57.1869
R10 VP.n13 VP.t0 57.1869
R11 VP.n4 VP.n3 47.115
R12 VP.n7 VP.n1 40.577
R13 VP.n11 VP.n1 40.577
R14 VP.n7 VP.n6 24.5923
R15 VP.n12 VP.n11 24.5923
R16 VP.n6 VP.n5 2.45968
R17 VP.n13 VP.n12 2.45968
R18 VP.n4 VP.n2 0.189894
R19 VP.n8 VP.n2 0.189894
R20 VP.n9 VP.n8 0.189894
R21 VP.n10 VP.n9 0.189894
R22 VP.n10 VP.n0 0.189894
R23 VP.n14 VP.n0 0.189894
R24 VP VP.n14 0.0516364
R25 VTAIL.n5 VTAIL.t4 99.4471
R26 VTAIL.n4 VTAIL.t2 99.4471
R27 VTAIL.n3 VTAIL.t0 99.4471
R28 VTAIL.n7 VTAIL.t1 99.4469
R29 VTAIL.n0 VTAIL.t3 99.4469
R30 VTAIL.n1 VTAIL.t5 99.4469
R31 VTAIL.n2 VTAIL.t6 99.4469
R32 VTAIL.n6 VTAIL.t7 99.4469
R33 VTAIL.n7 VTAIL.n6 17.7979
R34 VTAIL.n3 VTAIL.n2 17.7979
R35 VTAIL.n4 VTAIL.n3 1.81084
R36 VTAIL.n6 VTAIL.n5 1.81084
R37 VTAIL.n2 VTAIL.n1 1.81084
R38 VTAIL VTAIL.n0 0.963862
R39 VTAIL VTAIL.n7 0.847483
R40 VTAIL.n5 VTAIL.n4 0.470328
R41 VTAIL.n1 VTAIL.n0 0.470328
R42 VDD1 VDD1.n1 141.678
R43 VDD1 VDD1.n0 108.445
R44 VDD1.n0 VDD1.t0 7.73979
R45 VDD1.n0 VDD1.t1 7.73979
R46 VDD1.n1 VDD1.t2 7.73979
R47 VDD1.n1 VDD1.t3 7.73979
R48 B.n220 B.n219 585
R49 B.n218 B.n71 585
R50 B.n217 B.n216 585
R51 B.n215 B.n72 585
R52 B.n214 B.n213 585
R53 B.n212 B.n73 585
R54 B.n211 B.n210 585
R55 B.n209 B.n74 585
R56 B.n208 B.n207 585
R57 B.n206 B.n75 585
R58 B.n205 B.n204 585
R59 B.n203 B.n76 585
R60 B.n202 B.n201 585
R61 B.n200 B.n77 585
R62 B.n199 B.n198 585
R63 B.n197 B.n78 585
R64 B.n196 B.n195 585
R65 B.n194 B.n79 585
R66 B.n193 B.n192 585
R67 B.n190 B.n80 585
R68 B.n189 B.n188 585
R69 B.n187 B.n83 585
R70 B.n186 B.n185 585
R71 B.n184 B.n84 585
R72 B.n183 B.n182 585
R73 B.n181 B.n85 585
R74 B.n180 B.n179 585
R75 B.n178 B.n86 585
R76 B.n176 B.n175 585
R77 B.n174 B.n89 585
R78 B.n173 B.n172 585
R79 B.n171 B.n90 585
R80 B.n170 B.n169 585
R81 B.n168 B.n91 585
R82 B.n167 B.n166 585
R83 B.n165 B.n92 585
R84 B.n164 B.n163 585
R85 B.n162 B.n93 585
R86 B.n161 B.n160 585
R87 B.n159 B.n94 585
R88 B.n158 B.n157 585
R89 B.n156 B.n95 585
R90 B.n155 B.n154 585
R91 B.n153 B.n96 585
R92 B.n152 B.n151 585
R93 B.n150 B.n97 585
R94 B.n149 B.n148 585
R95 B.n221 B.n70 585
R96 B.n223 B.n222 585
R97 B.n224 B.n69 585
R98 B.n226 B.n225 585
R99 B.n227 B.n68 585
R100 B.n229 B.n228 585
R101 B.n230 B.n67 585
R102 B.n232 B.n231 585
R103 B.n233 B.n66 585
R104 B.n235 B.n234 585
R105 B.n236 B.n65 585
R106 B.n238 B.n237 585
R107 B.n239 B.n64 585
R108 B.n241 B.n240 585
R109 B.n242 B.n63 585
R110 B.n244 B.n243 585
R111 B.n245 B.n62 585
R112 B.n247 B.n246 585
R113 B.n248 B.n61 585
R114 B.n250 B.n249 585
R115 B.n251 B.n60 585
R116 B.n253 B.n252 585
R117 B.n254 B.n59 585
R118 B.n256 B.n255 585
R119 B.n257 B.n58 585
R120 B.n259 B.n258 585
R121 B.n260 B.n57 585
R122 B.n262 B.n261 585
R123 B.n263 B.n56 585
R124 B.n265 B.n264 585
R125 B.n266 B.n55 585
R126 B.n268 B.n267 585
R127 B.n269 B.n54 585
R128 B.n271 B.n270 585
R129 B.n272 B.n53 585
R130 B.n274 B.n273 585
R131 B.n275 B.n52 585
R132 B.n277 B.n276 585
R133 B.n278 B.n51 585
R134 B.n280 B.n279 585
R135 B.n281 B.n50 585
R136 B.n283 B.n282 585
R137 B.n284 B.n49 585
R138 B.n286 B.n285 585
R139 B.n287 B.n48 585
R140 B.n289 B.n288 585
R141 B.n290 B.n47 585
R142 B.n292 B.n291 585
R143 B.n293 B.n46 585
R144 B.n295 B.n294 585
R145 B.n296 B.n45 585
R146 B.n298 B.n297 585
R147 B.n299 B.n44 585
R148 B.n301 B.n300 585
R149 B.n372 B.n15 585
R150 B.n371 B.n370 585
R151 B.n369 B.n16 585
R152 B.n368 B.n367 585
R153 B.n366 B.n17 585
R154 B.n365 B.n364 585
R155 B.n363 B.n18 585
R156 B.n362 B.n361 585
R157 B.n360 B.n19 585
R158 B.n359 B.n358 585
R159 B.n357 B.n20 585
R160 B.n356 B.n355 585
R161 B.n354 B.n21 585
R162 B.n353 B.n352 585
R163 B.n351 B.n22 585
R164 B.n350 B.n349 585
R165 B.n348 B.n23 585
R166 B.n347 B.n346 585
R167 B.n345 B.n24 585
R168 B.n344 B.n343 585
R169 B.n342 B.n25 585
R170 B.n341 B.n340 585
R171 B.n339 B.n29 585
R172 B.n338 B.n337 585
R173 B.n336 B.n30 585
R174 B.n335 B.n334 585
R175 B.n333 B.n31 585
R176 B.n332 B.n331 585
R177 B.n329 B.n32 585
R178 B.n328 B.n327 585
R179 B.n326 B.n35 585
R180 B.n325 B.n324 585
R181 B.n323 B.n36 585
R182 B.n322 B.n321 585
R183 B.n320 B.n37 585
R184 B.n319 B.n318 585
R185 B.n317 B.n38 585
R186 B.n316 B.n315 585
R187 B.n314 B.n39 585
R188 B.n313 B.n312 585
R189 B.n311 B.n40 585
R190 B.n310 B.n309 585
R191 B.n308 B.n41 585
R192 B.n307 B.n306 585
R193 B.n305 B.n42 585
R194 B.n304 B.n303 585
R195 B.n302 B.n43 585
R196 B.n374 B.n373 585
R197 B.n375 B.n14 585
R198 B.n377 B.n376 585
R199 B.n378 B.n13 585
R200 B.n380 B.n379 585
R201 B.n381 B.n12 585
R202 B.n383 B.n382 585
R203 B.n384 B.n11 585
R204 B.n386 B.n385 585
R205 B.n387 B.n10 585
R206 B.n389 B.n388 585
R207 B.n390 B.n9 585
R208 B.n392 B.n391 585
R209 B.n393 B.n8 585
R210 B.n395 B.n394 585
R211 B.n396 B.n7 585
R212 B.n398 B.n397 585
R213 B.n399 B.n6 585
R214 B.n401 B.n400 585
R215 B.n402 B.n5 585
R216 B.n404 B.n403 585
R217 B.n405 B.n4 585
R218 B.n407 B.n406 585
R219 B.n408 B.n3 585
R220 B.n410 B.n409 585
R221 B.n411 B.n0 585
R222 B.n2 B.n1 585
R223 B.n111 B.n110 585
R224 B.n113 B.n112 585
R225 B.n114 B.n109 585
R226 B.n116 B.n115 585
R227 B.n117 B.n108 585
R228 B.n119 B.n118 585
R229 B.n120 B.n107 585
R230 B.n122 B.n121 585
R231 B.n123 B.n106 585
R232 B.n125 B.n124 585
R233 B.n126 B.n105 585
R234 B.n128 B.n127 585
R235 B.n129 B.n104 585
R236 B.n131 B.n130 585
R237 B.n132 B.n103 585
R238 B.n134 B.n133 585
R239 B.n135 B.n102 585
R240 B.n137 B.n136 585
R241 B.n138 B.n101 585
R242 B.n140 B.n139 585
R243 B.n141 B.n100 585
R244 B.n143 B.n142 585
R245 B.n144 B.n99 585
R246 B.n146 B.n145 585
R247 B.n147 B.n98 585
R248 B.n149 B.n98 516.524
R249 B.n219 B.n70 516.524
R250 B.n302 B.n301 516.524
R251 B.n374 B.n15 516.524
R252 B.n87 B.t9 263.509
R253 B.n81 B.t6 263.509
R254 B.n33 B.t3 263.509
R255 B.n26 B.t0 263.509
R256 B.n413 B.n412 256.663
R257 B.n412 B.n411 235.042
R258 B.n412 B.n2 235.042
R259 B.n150 B.n149 163.367
R260 B.n151 B.n150 163.367
R261 B.n151 B.n96 163.367
R262 B.n155 B.n96 163.367
R263 B.n156 B.n155 163.367
R264 B.n157 B.n156 163.367
R265 B.n157 B.n94 163.367
R266 B.n161 B.n94 163.367
R267 B.n162 B.n161 163.367
R268 B.n163 B.n162 163.367
R269 B.n163 B.n92 163.367
R270 B.n167 B.n92 163.367
R271 B.n168 B.n167 163.367
R272 B.n169 B.n168 163.367
R273 B.n169 B.n90 163.367
R274 B.n173 B.n90 163.367
R275 B.n174 B.n173 163.367
R276 B.n175 B.n174 163.367
R277 B.n175 B.n86 163.367
R278 B.n180 B.n86 163.367
R279 B.n181 B.n180 163.367
R280 B.n182 B.n181 163.367
R281 B.n182 B.n84 163.367
R282 B.n186 B.n84 163.367
R283 B.n187 B.n186 163.367
R284 B.n188 B.n187 163.367
R285 B.n188 B.n80 163.367
R286 B.n193 B.n80 163.367
R287 B.n194 B.n193 163.367
R288 B.n195 B.n194 163.367
R289 B.n195 B.n78 163.367
R290 B.n199 B.n78 163.367
R291 B.n200 B.n199 163.367
R292 B.n201 B.n200 163.367
R293 B.n201 B.n76 163.367
R294 B.n205 B.n76 163.367
R295 B.n206 B.n205 163.367
R296 B.n207 B.n206 163.367
R297 B.n207 B.n74 163.367
R298 B.n211 B.n74 163.367
R299 B.n212 B.n211 163.367
R300 B.n213 B.n212 163.367
R301 B.n213 B.n72 163.367
R302 B.n217 B.n72 163.367
R303 B.n218 B.n217 163.367
R304 B.n219 B.n218 163.367
R305 B.n301 B.n44 163.367
R306 B.n297 B.n44 163.367
R307 B.n297 B.n296 163.367
R308 B.n296 B.n295 163.367
R309 B.n295 B.n46 163.367
R310 B.n291 B.n46 163.367
R311 B.n291 B.n290 163.367
R312 B.n290 B.n289 163.367
R313 B.n289 B.n48 163.367
R314 B.n285 B.n48 163.367
R315 B.n285 B.n284 163.367
R316 B.n284 B.n283 163.367
R317 B.n283 B.n50 163.367
R318 B.n279 B.n50 163.367
R319 B.n279 B.n278 163.367
R320 B.n278 B.n277 163.367
R321 B.n277 B.n52 163.367
R322 B.n273 B.n52 163.367
R323 B.n273 B.n272 163.367
R324 B.n272 B.n271 163.367
R325 B.n271 B.n54 163.367
R326 B.n267 B.n54 163.367
R327 B.n267 B.n266 163.367
R328 B.n266 B.n265 163.367
R329 B.n265 B.n56 163.367
R330 B.n261 B.n56 163.367
R331 B.n261 B.n260 163.367
R332 B.n260 B.n259 163.367
R333 B.n259 B.n58 163.367
R334 B.n255 B.n58 163.367
R335 B.n255 B.n254 163.367
R336 B.n254 B.n253 163.367
R337 B.n253 B.n60 163.367
R338 B.n249 B.n60 163.367
R339 B.n249 B.n248 163.367
R340 B.n248 B.n247 163.367
R341 B.n247 B.n62 163.367
R342 B.n243 B.n62 163.367
R343 B.n243 B.n242 163.367
R344 B.n242 B.n241 163.367
R345 B.n241 B.n64 163.367
R346 B.n237 B.n64 163.367
R347 B.n237 B.n236 163.367
R348 B.n236 B.n235 163.367
R349 B.n235 B.n66 163.367
R350 B.n231 B.n66 163.367
R351 B.n231 B.n230 163.367
R352 B.n230 B.n229 163.367
R353 B.n229 B.n68 163.367
R354 B.n225 B.n68 163.367
R355 B.n225 B.n224 163.367
R356 B.n224 B.n223 163.367
R357 B.n223 B.n70 163.367
R358 B.n370 B.n15 163.367
R359 B.n370 B.n369 163.367
R360 B.n369 B.n368 163.367
R361 B.n368 B.n17 163.367
R362 B.n364 B.n17 163.367
R363 B.n364 B.n363 163.367
R364 B.n363 B.n362 163.367
R365 B.n362 B.n19 163.367
R366 B.n358 B.n19 163.367
R367 B.n358 B.n357 163.367
R368 B.n357 B.n356 163.367
R369 B.n356 B.n21 163.367
R370 B.n352 B.n21 163.367
R371 B.n352 B.n351 163.367
R372 B.n351 B.n350 163.367
R373 B.n350 B.n23 163.367
R374 B.n346 B.n23 163.367
R375 B.n346 B.n345 163.367
R376 B.n345 B.n344 163.367
R377 B.n344 B.n25 163.367
R378 B.n340 B.n25 163.367
R379 B.n340 B.n339 163.367
R380 B.n339 B.n338 163.367
R381 B.n338 B.n30 163.367
R382 B.n334 B.n30 163.367
R383 B.n334 B.n333 163.367
R384 B.n333 B.n332 163.367
R385 B.n332 B.n32 163.367
R386 B.n327 B.n32 163.367
R387 B.n327 B.n326 163.367
R388 B.n326 B.n325 163.367
R389 B.n325 B.n36 163.367
R390 B.n321 B.n36 163.367
R391 B.n321 B.n320 163.367
R392 B.n320 B.n319 163.367
R393 B.n319 B.n38 163.367
R394 B.n315 B.n38 163.367
R395 B.n315 B.n314 163.367
R396 B.n314 B.n313 163.367
R397 B.n313 B.n40 163.367
R398 B.n309 B.n40 163.367
R399 B.n309 B.n308 163.367
R400 B.n308 B.n307 163.367
R401 B.n307 B.n42 163.367
R402 B.n303 B.n42 163.367
R403 B.n303 B.n302 163.367
R404 B.n375 B.n374 163.367
R405 B.n376 B.n375 163.367
R406 B.n376 B.n13 163.367
R407 B.n380 B.n13 163.367
R408 B.n381 B.n380 163.367
R409 B.n382 B.n381 163.367
R410 B.n382 B.n11 163.367
R411 B.n386 B.n11 163.367
R412 B.n387 B.n386 163.367
R413 B.n388 B.n387 163.367
R414 B.n388 B.n9 163.367
R415 B.n392 B.n9 163.367
R416 B.n393 B.n392 163.367
R417 B.n394 B.n393 163.367
R418 B.n394 B.n7 163.367
R419 B.n398 B.n7 163.367
R420 B.n399 B.n398 163.367
R421 B.n400 B.n399 163.367
R422 B.n400 B.n5 163.367
R423 B.n404 B.n5 163.367
R424 B.n405 B.n404 163.367
R425 B.n406 B.n405 163.367
R426 B.n406 B.n3 163.367
R427 B.n410 B.n3 163.367
R428 B.n411 B.n410 163.367
R429 B.n110 B.n2 163.367
R430 B.n113 B.n110 163.367
R431 B.n114 B.n113 163.367
R432 B.n115 B.n114 163.367
R433 B.n115 B.n108 163.367
R434 B.n119 B.n108 163.367
R435 B.n120 B.n119 163.367
R436 B.n121 B.n120 163.367
R437 B.n121 B.n106 163.367
R438 B.n125 B.n106 163.367
R439 B.n126 B.n125 163.367
R440 B.n127 B.n126 163.367
R441 B.n127 B.n104 163.367
R442 B.n131 B.n104 163.367
R443 B.n132 B.n131 163.367
R444 B.n133 B.n132 163.367
R445 B.n133 B.n102 163.367
R446 B.n137 B.n102 163.367
R447 B.n138 B.n137 163.367
R448 B.n139 B.n138 163.367
R449 B.n139 B.n100 163.367
R450 B.n143 B.n100 163.367
R451 B.n144 B.n143 163.367
R452 B.n145 B.n144 163.367
R453 B.n145 B.n98 163.367
R454 B.n81 B.t7 161.917
R455 B.n33 B.t5 161.917
R456 B.n87 B.t10 161.915
R457 B.n26 B.t2 161.915
R458 B.n82 B.t8 121.191
R459 B.n34 B.t4 121.191
R460 B.n88 B.t11 121.188
R461 B.n27 B.t1 121.188
R462 B.n177 B.n88 59.5399
R463 B.n191 B.n82 59.5399
R464 B.n330 B.n34 59.5399
R465 B.n28 B.n27 59.5399
R466 B.n88 B.n87 40.7278
R467 B.n82 B.n81 40.7278
R468 B.n34 B.n33 40.7278
R469 B.n27 B.n26 40.7278
R470 B.n373 B.n372 33.5615
R471 B.n300 B.n43 33.5615
R472 B.n221 B.n220 33.5615
R473 B.n148 B.n147 33.5615
R474 B B.n413 18.0485
R475 B.n373 B.n14 10.6151
R476 B.n377 B.n14 10.6151
R477 B.n378 B.n377 10.6151
R478 B.n379 B.n378 10.6151
R479 B.n379 B.n12 10.6151
R480 B.n383 B.n12 10.6151
R481 B.n384 B.n383 10.6151
R482 B.n385 B.n384 10.6151
R483 B.n385 B.n10 10.6151
R484 B.n389 B.n10 10.6151
R485 B.n390 B.n389 10.6151
R486 B.n391 B.n390 10.6151
R487 B.n391 B.n8 10.6151
R488 B.n395 B.n8 10.6151
R489 B.n396 B.n395 10.6151
R490 B.n397 B.n396 10.6151
R491 B.n397 B.n6 10.6151
R492 B.n401 B.n6 10.6151
R493 B.n402 B.n401 10.6151
R494 B.n403 B.n402 10.6151
R495 B.n403 B.n4 10.6151
R496 B.n407 B.n4 10.6151
R497 B.n408 B.n407 10.6151
R498 B.n409 B.n408 10.6151
R499 B.n409 B.n0 10.6151
R500 B.n372 B.n371 10.6151
R501 B.n371 B.n16 10.6151
R502 B.n367 B.n16 10.6151
R503 B.n367 B.n366 10.6151
R504 B.n366 B.n365 10.6151
R505 B.n365 B.n18 10.6151
R506 B.n361 B.n18 10.6151
R507 B.n361 B.n360 10.6151
R508 B.n360 B.n359 10.6151
R509 B.n359 B.n20 10.6151
R510 B.n355 B.n20 10.6151
R511 B.n355 B.n354 10.6151
R512 B.n354 B.n353 10.6151
R513 B.n353 B.n22 10.6151
R514 B.n349 B.n22 10.6151
R515 B.n349 B.n348 10.6151
R516 B.n348 B.n347 10.6151
R517 B.n347 B.n24 10.6151
R518 B.n343 B.n342 10.6151
R519 B.n342 B.n341 10.6151
R520 B.n341 B.n29 10.6151
R521 B.n337 B.n29 10.6151
R522 B.n337 B.n336 10.6151
R523 B.n336 B.n335 10.6151
R524 B.n335 B.n31 10.6151
R525 B.n331 B.n31 10.6151
R526 B.n329 B.n328 10.6151
R527 B.n328 B.n35 10.6151
R528 B.n324 B.n35 10.6151
R529 B.n324 B.n323 10.6151
R530 B.n323 B.n322 10.6151
R531 B.n322 B.n37 10.6151
R532 B.n318 B.n37 10.6151
R533 B.n318 B.n317 10.6151
R534 B.n317 B.n316 10.6151
R535 B.n316 B.n39 10.6151
R536 B.n312 B.n39 10.6151
R537 B.n312 B.n311 10.6151
R538 B.n311 B.n310 10.6151
R539 B.n310 B.n41 10.6151
R540 B.n306 B.n41 10.6151
R541 B.n306 B.n305 10.6151
R542 B.n305 B.n304 10.6151
R543 B.n304 B.n43 10.6151
R544 B.n300 B.n299 10.6151
R545 B.n299 B.n298 10.6151
R546 B.n298 B.n45 10.6151
R547 B.n294 B.n45 10.6151
R548 B.n294 B.n293 10.6151
R549 B.n293 B.n292 10.6151
R550 B.n292 B.n47 10.6151
R551 B.n288 B.n47 10.6151
R552 B.n288 B.n287 10.6151
R553 B.n287 B.n286 10.6151
R554 B.n286 B.n49 10.6151
R555 B.n282 B.n49 10.6151
R556 B.n282 B.n281 10.6151
R557 B.n281 B.n280 10.6151
R558 B.n280 B.n51 10.6151
R559 B.n276 B.n51 10.6151
R560 B.n276 B.n275 10.6151
R561 B.n275 B.n274 10.6151
R562 B.n274 B.n53 10.6151
R563 B.n270 B.n53 10.6151
R564 B.n270 B.n269 10.6151
R565 B.n269 B.n268 10.6151
R566 B.n268 B.n55 10.6151
R567 B.n264 B.n55 10.6151
R568 B.n264 B.n263 10.6151
R569 B.n263 B.n262 10.6151
R570 B.n262 B.n57 10.6151
R571 B.n258 B.n57 10.6151
R572 B.n258 B.n257 10.6151
R573 B.n257 B.n256 10.6151
R574 B.n256 B.n59 10.6151
R575 B.n252 B.n59 10.6151
R576 B.n252 B.n251 10.6151
R577 B.n251 B.n250 10.6151
R578 B.n250 B.n61 10.6151
R579 B.n246 B.n61 10.6151
R580 B.n246 B.n245 10.6151
R581 B.n245 B.n244 10.6151
R582 B.n244 B.n63 10.6151
R583 B.n240 B.n63 10.6151
R584 B.n240 B.n239 10.6151
R585 B.n239 B.n238 10.6151
R586 B.n238 B.n65 10.6151
R587 B.n234 B.n65 10.6151
R588 B.n234 B.n233 10.6151
R589 B.n233 B.n232 10.6151
R590 B.n232 B.n67 10.6151
R591 B.n228 B.n67 10.6151
R592 B.n228 B.n227 10.6151
R593 B.n227 B.n226 10.6151
R594 B.n226 B.n69 10.6151
R595 B.n222 B.n69 10.6151
R596 B.n222 B.n221 10.6151
R597 B.n111 B.n1 10.6151
R598 B.n112 B.n111 10.6151
R599 B.n112 B.n109 10.6151
R600 B.n116 B.n109 10.6151
R601 B.n117 B.n116 10.6151
R602 B.n118 B.n117 10.6151
R603 B.n118 B.n107 10.6151
R604 B.n122 B.n107 10.6151
R605 B.n123 B.n122 10.6151
R606 B.n124 B.n123 10.6151
R607 B.n124 B.n105 10.6151
R608 B.n128 B.n105 10.6151
R609 B.n129 B.n128 10.6151
R610 B.n130 B.n129 10.6151
R611 B.n130 B.n103 10.6151
R612 B.n134 B.n103 10.6151
R613 B.n135 B.n134 10.6151
R614 B.n136 B.n135 10.6151
R615 B.n136 B.n101 10.6151
R616 B.n140 B.n101 10.6151
R617 B.n141 B.n140 10.6151
R618 B.n142 B.n141 10.6151
R619 B.n142 B.n99 10.6151
R620 B.n146 B.n99 10.6151
R621 B.n147 B.n146 10.6151
R622 B.n148 B.n97 10.6151
R623 B.n152 B.n97 10.6151
R624 B.n153 B.n152 10.6151
R625 B.n154 B.n153 10.6151
R626 B.n154 B.n95 10.6151
R627 B.n158 B.n95 10.6151
R628 B.n159 B.n158 10.6151
R629 B.n160 B.n159 10.6151
R630 B.n160 B.n93 10.6151
R631 B.n164 B.n93 10.6151
R632 B.n165 B.n164 10.6151
R633 B.n166 B.n165 10.6151
R634 B.n166 B.n91 10.6151
R635 B.n170 B.n91 10.6151
R636 B.n171 B.n170 10.6151
R637 B.n172 B.n171 10.6151
R638 B.n172 B.n89 10.6151
R639 B.n176 B.n89 10.6151
R640 B.n179 B.n178 10.6151
R641 B.n179 B.n85 10.6151
R642 B.n183 B.n85 10.6151
R643 B.n184 B.n183 10.6151
R644 B.n185 B.n184 10.6151
R645 B.n185 B.n83 10.6151
R646 B.n189 B.n83 10.6151
R647 B.n190 B.n189 10.6151
R648 B.n192 B.n79 10.6151
R649 B.n196 B.n79 10.6151
R650 B.n197 B.n196 10.6151
R651 B.n198 B.n197 10.6151
R652 B.n198 B.n77 10.6151
R653 B.n202 B.n77 10.6151
R654 B.n203 B.n202 10.6151
R655 B.n204 B.n203 10.6151
R656 B.n204 B.n75 10.6151
R657 B.n208 B.n75 10.6151
R658 B.n209 B.n208 10.6151
R659 B.n210 B.n209 10.6151
R660 B.n210 B.n73 10.6151
R661 B.n214 B.n73 10.6151
R662 B.n215 B.n214 10.6151
R663 B.n216 B.n215 10.6151
R664 B.n216 B.n71 10.6151
R665 B.n220 B.n71 10.6151
R666 B.n413 B.n0 8.11757
R667 B.n413 B.n1 8.11757
R668 B.n343 B.n28 6.5566
R669 B.n331 B.n330 6.5566
R670 B.n178 B.n177 6.5566
R671 B.n191 B.n190 6.5566
R672 B.n28 B.n24 4.05904
R673 B.n330 B.n329 4.05904
R674 B.n177 B.n176 4.05904
R675 B.n192 B.n191 4.05904
R676 VN.n0 VN.t2 93.3598
R677 VN.n1 VN.t1 93.3598
R678 VN.n0 VN.t0 92.9312
R679 VN.n1 VN.t3 92.9312
R680 VN VN.n1 47.4957
R681 VN VN.n0 9.3707
R682 VDD2.n2 VDD2.n0 141.153
R683 VDD2.n2 VDD2.n1 108.386
R684 VDD2.n1 VDD2.t0 7.73979
R685 VDD2.n1 VDD2.t2 7.73979
R686 VDD2.n0 VDD2.t1 7.73979
R687 VDD2.n0 VDD2.t3 7.73979
R688 VDD2 VDD2.n2 0.0586897
C0 VDD1 w_n2230_n1808# 1.0769f
C1 B w_n2230_n1808# 6.04532f
C2 VDD1 VN 0.152555f
C3 VN B 0.86405f
C4 VDD2 VP 0.346176f
C5 VP VTAIL 1.97009f
C6 VDD2 VTAIL 3.29438f
C7 VDD1 B 0.905609f
C8 VP w_n2230_n1808# 3.75628f
C9 VDD2 w_n2230_n1808# 1.1141f
C10 w_n2230_n1808# VTAIL 2.14646f
C11 VN VP 4.15103f
C12 VDD2 VN 1.73775f
C13 VN VTAIL 1.95598f
C14 VDD1 VP 1.93044f
C15 VDD1 VDD2 0.824331f
C16 VDD1 VTAIL 3.24573f
C17 VN w_n2230_n1808# 3.47232f
C18 VP B 1.33227f
C19 VDD2 B 0.944297f
C20 B VTAIL 2.09705f
C21 VDD2 VSUBS 0.567105f
C22 VDD1 VSUBS 2.865364f
C23 VTAIL VSUBS 0.509899f
C24 VN VSUBS 4.09383f
C25 VP VSUBS 1.401301f
C26 B VSUBS 2.756358f
C27 w_n2230_n1808# VSUBS 50.710197f
C28 VDD2.t1 VSUBS 0.059628f
C29 VDD2.t3 VSUBS 0.059628f
C30 VDD2.n0 VSUBS 0.552937f
C31 VDD2.t0 VSUBS 0.059628f
C32 VDD2.t2 VSUBS 0.059628f
C33 VDD2.n1 VSUBS 0.35428f
C34 VDD2.n2 VSUBS 2.0456f
C35 VN.t2 VSUBS 0.861548f
C36 VN.t0 VSUBS 0.859484f
C37 VN.n0 VSUBS 0.620838f
C38 VN.t1 VSUBS 0.861548f
C39 VN.t3 VSUBS 0.859484f
C40 VN.n1 VSUBS 1.81785f
C41 B.n0 VSUBS 0.008324f
C42 B.n1 VSUBS 0.008324f
C43 B.n2 VSUBS 0.012311f
C44 B.n3 VSUBS 0.009434f
C45 B.n4 VSUBS 0.009434f
C46 B.n5 VSUBS 0.009434f
C47 B.n6 VSUBS 0.009434f
C48 B.n7 VSUBS 0.009434f
C49 B.n8 VSUBS 0.009434f
C50 B.n9 VSUBS 0.009434f
C51 B.n10 VSUBS 0.009434f
C52 B.n11 VSUBS 0.009434f
C53 B.n12 VSUBS 0.009434f
C54 B.n13 VSUBS 0.009434f
C55 B.n14 VSUBS 0.009434f
C56 B.n15 VSUBS 0.023149f
C57 B.n16 VSUBS 0.009434f
C58 B.n17 VSUBS 0.009434f
C59 B.n18 VSUBS 0.009434f
C60 B.n19 VSUBS 0.009434f
C61 B.n20 VSUBS 0.009434f
C62 B.n21 VSUBS 0.009434f
C63 B.n22 VSUBS 0.009434f
C64 B.n23 VSUBS 0.009434f
C65 B.n24 VSUBS 0.00652f
C66 B.n25 VSUBS 0.009434f
C67 B.t1 VSUBS 0.150845f
C68 B.t2 VSUBS 0.169659f
C69 B.t0 VSUBS 0.473155f
C70 B.n26 VSUBS 0.116739f
C71 B.n27 VSUBS 0.088251f
C72 B.n28 VSUBS 0.021857f
C73 B.n29 VSUBS 0.009434f
C74 B.n30 VSUBS 0.009434f
C75 B.n31 VSUBS 0.009434f
C76 B.n32 VSUBS 0.009434f
C77 B.t4 VSUBS 0.150845f
C78 B.t5 VSUBS 0.169659f
C79 B.t3 VSUBS 0.473155f
C80 B.n33 VSUBS 0.116739f
C81 B.n34 VSUBS 0.088251f
C82 B.n35 VSUBS 0.009434f
C83 B.n36 VSUBS 0.009434f
C84 B.n37 VSUBS 0.009434f
C85 B.n38 VSUBS 0.009434f
C86 B.n39 VSUBS 0.009434f
C87 B.n40 VSUBS 0.009434f
C88 B.n41 VSUBS 0.009434f
C89 B.n42 VSUBS 0.009434f
C90 B.n43 VSUBS 0.023149f
C91 B.n44 VSUBS 0.009434f
C92 B.n45 VSUBS 0.009434f
C93 B.n46 VSUBS 0.009434f
C94 B.n47 VSUBS 0.009434f
C95 B.n48 VSUBS 0.009434f
C96 B.n49 VSUBS 0.009434f
C97 B.n50 VSUBS 0.009434f
C98 B.n51 VSUBS 0.009434f
C99 B.n52 VSUBS 0.009434f
C100 B.n53 VSUBS 0.009434f
C101 B.n54 VSUBS 0.009434f
C102 B.n55 VSUBS 0.009434f
C103 B.n56 VSUBS 0.009434f
C104 B.n57 VSUBS 0.009434f
C105 B.n58 VSUBS 0.009434f
C106 B.n59 VSUBS 0.009434f
C107 B.n60 VSUBS 0.009434f
C108 B.n61 VSUBS 0.009434f
C109 B.n62 VSUBS 0.009434f
C110 B.n63 VSUBS 0.009434f
C111 B.n64 VSUBS 0.009434f
C112 B.n65 VSUBS 0.009434f
C113 B.n66 VSUBS 0.009434f
C114 B.n67 VSUBS 0.009434f
C115 B.n68 VSUBS 0.009434f
C116 B.n69 VSUBS 0.009434f
C117 B.n70 VSUBS 0.0218f
C118 B.n71 VSUBS 0.009434f
C119 B.n72 VSUBS 0.009434f
C120 B.n73 VSUBS 0.009434f
C121 B.n74 VSUBS 0.009434f
C122 B.n75 VSUBS 0.009434f
C123 B.n76 VSUBS 0.009434f
C124 B.n77 VSUBS 0.009434f
C125 B.n78 VSUBS 0.009434f
C126 B.n79 VSUBS 0.009434f
C127 B.n80 VSUBS 0.009434f
C128 B.t8 VSUBS 0.150845f
C129 B.t7 VSUBS 0.169659f
C130 B.t6 VSUBS 0.473155f
C131 B.n81 VSUBS 0.116739f
C132 B.n82 VSUBS 0.088251f
C133 B.n83 VSUBS 0.009434f
C134 B.n84 VSUBS 0.009434f
C135 B.n85 VSUBS 0.009434f
C136 B.n86 VSUBS 0.009434f
C137 B.t11 VSUBS 0.150845f
C138 B.t10 VSUBS 0.169659f
C139 B.t9 VSUBS 0.473155f
C140 B.n87 VSUBS 0.116739f
C141 B.n88 VSUBS 0.088251f
C142 B.n89 VSUBS 0.009434f
C143 B.n90 VSUBS 0.009434f
C144 B.n91 VSUBS 0.009434f
C145 B.n92 VSUBS 0.009434f
C146 B.n93 VSUBS 0.009434f
C147 B.n94 VSUBS 0.009434f
C148 B.n95 VSUBS 0.009434f
C149 B.n96 VSUBS 0.009434f
C150 B.n97 VSUBS 0.009434f
C151 B.n98 VSUBS 0.0218f
C152 B.n99 VSUBS 0.009434f
C153 B.n100 VSUBS 0.009434f
C154 B.n101 VSUBS 0.009434f
C155 B.n102 VSUBS 0.009434f
C156 B.n103 VSUBS 0.009434f
C157 B.n104 VSUBS 0.009434f
C158 B.n105 VSUBS 0.009434f
C159 B.n106 VSUBS 0.009434f
C160 B.n107 VSUBS 0.009434f
C161 B.n108 VSUBS 0.009434f
C162 B.n109 VSUBS 0.009434f
C163 B.n110 VSUBS 0.009434f
C164 B.n111 VSUBS 0.009434f
C165 B.n112 VSUBS 0.009434f
C166 B.n113 VSUBS 0.009434f
C167 B.n114 VSUBS 0.009434f
C168 B.n115 VSUBS 0.009434f
C169 B.n116 VSUBS 0.009434f
C170 B.n117 VSUBS 0.009434f
C171 B.n118 VSUBS 0.009434f
C172 B.n119 VSUBS 0.009434f
C173 B.n120 VSUBS 0.009434f
C174 B.n121 VSUBS 0.009434f
C175 B.n122 VSUBS 0.009434f
C176 B.n123 VSUBS 0.009434f
C177 B.n124 VSUBS 0.009434f
C178 B.n125 VSUBS 0.009434f
C179 B.n126 VSUBS 0.009434f
C180 B.n127 VSUBS 0.009434f
C181 B.n128 VSUBS 0.009434f
C182 B.n129 VSUBS 0.009434f
C183 B.n130 VSUBS 0.009434f
C184 B.n131 VSUBS 0.009434f
C185 B.n132 VSUBS 0.009434f
C186 B.n133 VSUBS 0.009434f
C187 B.n134 VSUBS 0.009434f
C188 B.n135 VSUBS 0.009434f
C189 B.n136 VSUBS 0.009434f
C190 B.n137 VSUBS 0.009434f
C191 B.n138 VSUBS 0.009434f
C192 B.n139 VSUBS 0.009434f
C193 B.n140 VSUBS 0.009434f
C194 B.n141 VSUBS 0.009434f
C195 B.n142 VSUBS 0.009434f
C196 B.n143 VSUBS 0.009434f
C197 B.n144 VSUBS 0.009434f
C198 B.n145 VSUBS 0.009434f
C199 B.n146 VSUBS 0.009434f
C200 B.n147 VSUBS 0.0218f
C201 B.n148 VSUBS 0.023149f
C202 B.n149 VSUBS 0.023149f
C203 B.n150 VSUBS 0.009434f
C204 B.n151 VSUBS 0.009434f
C205 B.n152 VSUBS 0.009434f
C206 B.n153 VSUBS 0.009434f
C207 B.n154 VSUBS 0.009434f
C208 B.n155 VSUBS 0.009434f
C209 B.n156 VSUBS 0.009434f
C210 B.n157 VSUBS 0.009434f
C211 B.n158 VSUBS 0.009434f
C212 B.n159 VSUBS 0.009434f
C213 B.n160 VSUBS 0.009434f
C214 B.n161 VSUBS 0.009434f
C215 B.n162 VSUBS 0.009434f
C216 B.n163 VSUBS 0.009434f
C217 B.n164 VSUBS 0.009434f
C218 B.n165 VSUBS 0.009434f
C219 B.n166 VSUBS 0.009434f
C220 B.n167 VSUBS 0.009434f
C221 B.n168 VSUBS 0.009434f
C222 B.n169 VSUBS 0.009434f
C223 B.n170 VSUBS 0.009434f
C224 B.n171 VSUBS 0.009434f
C225 B.n172 VSUBS 0.009434f
C226 B.n173 VSUBS 0.009434f
C227 B.n174 VSUBS 0.009434f
C228 B.n175 VSUBS 0.009434f
C229 B.n176 VSUBS 0.00652f
C230 B.n177 VSUBS 0.021857f
C231 B.n178 VSUBS 0.00763f
C232 B.n179 VSUBS 0.009434f
C233 B.n180 VSUBS 0.009434f
C234 B.n181 VSUBS 0.009434f
C235 B.n182 VSUBS 0.009434f
C236 B.n183 VSUBS 0.009434f
C237 B.n184 VSUBS 0.009434f
C238 B.n185 VSUBS 0.009434f
C239 B.n186 VSUBS 0.009434f
C240 B.n187 VSUBS 0.009434f
C241 B.n188 VSUBS 0.009434f
C242 B.n189 VSUBS 0.009434f
C243 B.n190 VSUBS 0.00763f
C244 B.n191 VSUBS 0.021857f
C245 B.n192 VSUBS 0.00652f
C246 B.n193 VSUBS 0.009434f
C247 B.n194 VSUBS 0.009434f
C248 B.n195 VSUBS 0.009434f
C249 B.n196 VSUBS 0.009434f
C250 B.n197 VSUBS 0.009434f
C251 B.n198 VSUBS 0.009434f
C252 B.n199 VSUBS 0.009434f
C253 B.n200 VSUBS 0.009434f
C254 B.n201 VSUBS 0.009434f
C255 B.n202 VSUBS 0.009434f
C256 B.n203 VSUBS 0.009434f
C257 B.n204 VSUBS 0.009434f
C258 B.n205 VSUBS 0.009434f
C259 B.n206 VSUBS 0.009434f
C260 B.n207 VSUBS 0.009434f
C261 B.n208 VSUBS 0.009434f
C262 B.n209 VSUBS 0.009434f
C263 B.n210 VSUBS 0.009434f
C264 B.n211 VSUBS 0.009434f
C265 B.n212 VSUBS 0.009434f
C266 B.n213 VSUBS 0.009434f
C267 B.n214 VSUBS 0.009434f
C268 B.n215 VSUBS 0.009434f
C269 B.n216 VSUBS 0.009434f
C270 B.n217 VSUBS 0.009434f
C271 B.n218 VSUBS 0.009434f
C272 B.n219 VSUBS 0.023149f
C273 B.n220 VSUBS 0.022065f
C274 B.n221 VSUBS 0.022885f
C275 B.n222 VSUBS 0.009434f
C276 B.n223 VSUBS 0.009434f
C277 B.n224 VSUBS 0.009434f
C278 B.n225 VSUBS 0.009434f
C279 B.n226 VSUBS 0.009434f
C280 B.n227 VSUBS 0.009434f
C281 B.n228 VSUBS 0.009434f
C282 B.n229 VSUBS 0.009434f
C283 B.n230 VSUBS 0.009434f
C284 B.n231 VSUBS 0.009434f
C285 B.n232 VSUBS 0.009434f
C286 B.n233 VSUBS 0.009434f
C287 B.n234 VSUBS 0.009434f
C288 B.n235 VSUBS 0.009434f
C289 B.n236 VSUBS 0.009434f
C290 B.n237 VSUBS 0.009434f
C291 B.n238 VSUBS 0.009434f
C292 B.n239 VSUBS 0.009434f
C293 B.n240 VSUBS 0.009434f
C294 B.n241 VSUBS 0.009434f
C295 B.n242 VSUBS 0.009434f
C296 B.n243 VSUBS 0.009434f
C297 B.n244 VSUBS 0.009434f
C298 B.n245 VSUBS 0.009434f
C299 B.n246 VSUBS 0.009434f
C300 B.n247 VSUBS 0.009434f
C301 B.n248 VSUBS 0.009434f
C302 B.n249 VSUBS 0.009434f
C303 B.n250 VSUBS 0.009434f
C304 B.n251 VSUBS 0.009434f
C305 B.n252 VSUBS 0.009434f
C306 B.n253 VSUBS 0.009434f
C307 B.n254 VSUBS 0.009434f
C308 B.n255 VSUBS 0.009434f
C309 B.n256 VSUBS 0.009434f
C310 B.n257 VSUBS 0.009434f
C311 B.n258 VSUBS 0.009434f
C312 B.n259 VSUBS 0.009434f
C313 B.n260 VSUBS 0.009434f
C314 B.n261 VSUBS 0.009434f
C315 B.n262 VSUBS 0.009434f
C316 B.n263 VSUBS 0.009434f
C317 B.n264 VSUBS 0.009434f
C318 B.n265 VSUBS 0.009434f
C319 B.n266 VSUBS 0.009434f
C320 B.n267 VSUBS 0.009434f
C321 B.n268 VSUBS 0.009434f
C322 B.n269 VSUBS 0.009434f
C323 B.n270 VSUBS 0.009434f
C324 B.n271 VSUBS 0.009434f
C325 B.n272 VSUBS 0.009434f
C326 B.n273 VSUBS 0.009434f
C327 B.n274 VSUBS 0.009434f
C328 B.n275 VSUBS 0.009434f
C329 B.n276 VSUBS 0.009434f
C330 B.n277 VSUBS 0.009434f
C331 B.n278 VSUBS 0.009434f
C332 B.n279 VSUBS 0.009434f
C333 B.n280 VSUBS 0.009434f
C334 B.n281 VSUBS 0.009434f
C335 B.n282 VSUBS 0.009434f
C336 B.n283 VSUBS 0.009434f
C337 B.n284 VSUBS 0.009434f
C338 B.n285 VSUBS 0.009434f
C339 B.n286 VSUBS 0.009434f
C340 B.n287 VSUBS 0.009434f
C341 B.n288 VSUBS 0.009434f
C342 B.n289 VSUBS 0.009434f
C343 B.n290 VSUBS 0.009434f
C344 B.n291 VSUBS 0.009434f
C345 B.n292 VSUBS 0.009434f
C346 B.n293 VSUBS 0.009434f
C347 B.n294 VSUBS 0.009434f
C348 B.n295 VSUBS 0.009434f
C349 B.n296 VSUBS 0.009434f
C350 B.n297 VSUBS 0.009434f
C351 B.n298 VSUBS 0.009434f
C352 B.n299 VSUBS 0.009434f
C353 B.n300 VSUBS 0.0218f
C354 B.n301 VSUBS 0.0218f
C355 B.n302 VSUBS 0.023149f
C356 B.n303 VSUBS 0.009434f
C357 B.n304 VSUBS 0.009434f
C358 B.n305 VSUBS 0.009434f
C359 B.n306 VSUBS 0.009434f
C360 B.n307 VSUBS 0.009434f
C361 B.n308 VSUBS 0.009434f
C362 B.n309 VSUBS 0.009434f
C363 B.n310 VSUBS 0.009434f
C364 B.n311 VSUBS 0.009434f
C365 B.n312 VSUBS 0.009434f
C366 B.n313 VSUBS 0.009434f
C367 B.n314 VSUBS 0.009434f
C368 B.n315 VSUBS 0.009434f
C369 B.n316 VSUBS 0.009434f
C370 B.n317 VSUBS 0.009434f
C371 B.n318 VSUBS 0.009434f
C372 B.n319 VSUBS 0.009434f
C373 B.n320 VSUBS 0.009434f
C374 B.n321 VSUBS 0.009434f
C375 B.n322 VSUBS 0.009434f
C376 B.n323 VSUBS 0.009434f
C377 B.n324 VSUBS 0.009434f
C378 B.n325 VSUBS 0.009434f
C379 B.n326 VSUBS 0.009434f
C380 B.n327 VSUBS 0.009434f
C381 B.n328 VSUBS 0.009434f
C382 B.n329 VSUBS 0.00652f
C383 B.n330 VSUBS 0.021857f
C384 B.n331 VSUBS 0.00763f
C385 B.n332 VSUBS 0.009434f
C386 B.n333 VSUBS 0.009434f
C387 B.n334 VSUBS 0.009434f
C388 B.n335 VSUBS 0.009434f
C389 B.n336 VSUBS 0.009434f
C390 B.n337 VSUBS 0.009434f
C391 B.n338 VSUBS 0.009434f
C392 B.n339 VSUBS 0.009434f
C393 B.n340 VSUBS 0.009434f
C394 B.n341 VSUBS 0.009434f
C395 B.n342 VSUBS 0.009434f
C396 B.n343 VSUBS 0.00763f
C397 B.n344 VSUBS 0.009434f
C398 B.n345 VSUBS 0.009434f
C399 B.n346 VSUBS 0.009434f
C400 B.n347 VSUBS 0.009434f
C401 B.n348 VSUBS 0.009434f
C402 B.n349 VSUBS 0.009434f
C403 B.n350 VSUBS 0.009434f
C404 B.n351 VSUBS 0.009434f
C405 B.n352 VSUBS 0.009434f
C406 B.n353 VSUBS 0.009434f
C407 B.n354 VSUBS 0.009434f
C408 B.n355 VSUBS 0.009434f
C409 B.n356 VSUBS 0.009434f
C410 B.n357 VSUBS 0.009434f
C411 B.n358 VSUBS 0.009434f
C412 B.n359 VSUBS 0.009434f
C413 B.n360 VSUBS 0.009434f
C414 B.n361 VSUBS 0.009434f
C415 B.n362 VSUBS 0.009434f
C416 B.n363 VSUBS 0.009434f
C417 B.n364 VSUBS 0.009434f
C418 B.n365 VSUBS 0.009434f
C419 B.n366 VSUBS 0.009434f
C420 B.n367 VSUBS 0.009434f
C421 B.n368 VSUBS 0.009434f
C422 B.n369 VSUBS 0.009434f
C423 B.n370 VSUBS 0.009434f
C424 B.n371 VSUBS 0.009434f
C425 B.n372 VSUBS 0.023149f
C426 B.n373 VSUBS 0.0218f
C427 B.n374 VSUBS 0.0218f
C428 B.n375 VSUBS 0.009434f
C429 B.n376 VSUBS 0.009434f
C430 B.n377 VSUBS 0.009434f
C431 B.n378 VSUBS 0.009434f
C432 B.n379 VSUBS 0.009434f
C433 B.n380 VSUBS 0.009434f
C434 B.n381 VSUBS 0.009434f
C435 B.n382 VSUBS 0.009434f
C436 B.n383 VSUBS 0.009434f
C437 B.n384 VSUBS 0.009434f
C438 B.n385 VSUBS 0.009434f
C439 B.n386 VSUBS 0.009434f
C440 B.n387 VSUBS 0.009434f
C441 B.n388 VSUBS 0.009434f
C442 B.n389 VSUBS 0.009434f
C443 B.n390 VSUBS 0.009434f
C444 B.n391 VSUBS 0.009434f
C445 B.n392 VSUBS 0.009434f
C446 B.n393 VSUBS 0.009434f
C447 B.n394 VSUBS 0.009434f
C448 B.n395 VSUBS 0.009434f
C449 B.n396 VSUBS 0.009434f
C450 B.n397 VSUBS 0.009434f
C451 B.n398 VSUBS 0.009434f
C452 B.n399 VSUBS 0.009434f
C453 B.n400 VSUBS 0.009434f
C454 B.n401 VSUBS 0.009434f
C455 B.n402 VSUBS 0.009434f
C456 B.n403 VSUBS 0.009434f
C457 B.n404 VSUBS 0.009434f
C458 B.n405 VSUBS 0.009434f
C459 B.n406 VSUBS 0.009434f
C460 B.n407 VSUBS 0.009434f
C461 B.n408 VSUBS 0.009434f
C462 B.n409 VSUBS 0.009434f
C463 B.n410 VSUBS 0.009434f
C464 B.n411 VSUBS 0.012311f
C465 B.n412 VSUBS 0.013114f
C466 B.n413 VSUBS 0.026078f
C467 VDD1.t0 VSUBS 0.056681f
C468 VDD1.t1 VSUBS 0.056681f
C469 VDD1.n0 VSUBS 0.336963f
C470 VDD1.t2 VSUBS 0.056681f
C471 VDD1.t3 VSUBS 0.056681f
C472 VDD1.n1 VSUBS 0.536101f
C473 VTAIL.t3 VSUBS 0.510461f
C474 VTAIL.n0 VSUBS 0.460733f
C475 VTAIL.t5 VSUBS 0.510461f
C476 VTAIL.n1 VSUBS 0.517813f
C477 VTAIL.t6 VSUBS 0.510461f
C478 VTAIL.n2 VSUBS 1.13626f
C479 VTAIL.t0 VSUBS 0.510463f
C480 VTAIL.n3 VSUBS 1.13626f
C481 VTAIL.t2 VSUBS 0.510463f
C482 VTAIL.n4 VSUBS 0.517811f
C483 VTAIL.t4 VSUBS 0.510463f
C484 VTAIL.n5 VSUBS 0.517811f
C485 VTAIL.t7 VSUBS 0.510461f
C486 VTAIL.n6 VSUBS 1.13626f
C487 VTAIL.t1 VSUBS 0.510461f
C488 VTAIL.n7 VSUBS 1.07134f
C489 VP.n0 VSUBS 0.037427f
C490 VP.t0 VSUBS 0.717861f
C491 VP.n1 VSUBS 0.030229f
C492 VP.n2 VSUBS 0.037427f
C493 VP.t1 VSUBS 0.717861f
C494 VP.t3 VSUBS 0.901002f
C495 VP.t2 VSUBS 0.898843f
C496 VP.n3 VSUBS 1.87878f
C497 VP.n4 VSUBS 1.63719f
C498 VP.n5 VSUBS 0.374493f
C499 VP.n6 VSUBS 0.038568f
C500 VP.n7 VSUBS 0.073995f
C501 VP.n8 VSUBS 0.037427f
C502 VP.n9 VSUBS 0.037427f
C503 VP.n10 VSUBS 0.037427f
C504 VP.n11 VSUBS 0.073995f
C505 VP.n12 VSUBS 0.038568f
C506 VP.n13 VSUBS 0.374493f
C507 VP.n14 VSUBS 0.040025f
.ends

