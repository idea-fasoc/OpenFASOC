* NGSPICE file created from diff_pair_sample_1011.ext - technology: sky130A

.subckt diff_pair_sample_1011 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=5.8305 pd=30.68 as=0 ps=0 w=14.95 l=3.03
X1 B.t12 B.t10 B.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=5.8305 pd=30.68 as=0 ps=0 w=14.95 l=3.03
X2 VDD2.t1 VN.t0 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=5.8305 pd=30.68 as=5.8305 ps=30.68 w=14.95 l=3.03
X3 VDD1.t1 VP.t0 VTAIL.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=5.8305 pd=30.68 as=5.8305 ps=30.68 w=14.95 l=3.03
X4 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=5.8305 pd=30.68 as=0 ps=0 w=14.95 l=3.03
X5 VDD2.t0 VN.t1 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=5.8305 pd=30.68 as=5.8305 ps=30.68 w=14.95 l=3.03
X6 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=5.8305 pd=30.68 as=0 ps=0 w=14.95 l=3.03
X7 VDD1.t0 VP.t1 VTAIL.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=5.8305 pd=30.68 as=5.8305 ps=30.68 w=14.95 l=3.03
R0 B.n786 B.n785 585
R1 B.n330 B.n109 585
R2 B.n329 B.n328 585
R3 B.n327 B.n326 585
R4 B.n325 B.n324 585
R5 B.n323 B.n322 585
R6 B.n321 B.n320 585
R7 B.n319 B.n318 585
R8 B.n317 B.n316 585
R9 B.n315 B.n314 585
R10 B.n313 B.n312 585
R11 B.n311 B.n310 585
R12 B.n309 B.n308 585
R13 B.n307 B.n306 585
R14 B.n305 B.n304 585
R15 B.n303 B.n302 585
R16 B.n301 B.n300 585
R17 B.n299 B.n298 585
R18 B.n297 B.n296 585
R19 B.n295 B.n294 585
R20 B.n293 B.n292 585
R21 B.n291 B.n290 585
R22 B.n289 B.n288 585
R23 B.n287 B.n286 585
R24 B.n285 B.n284 585
R25 B.n283 B.n282 585
R26 B.n281 B.n280 585
R27 B.n279 B.n278 585
R28 B.n277 B.n276 585
R29 B.n275 B.n274 585
R30 B.n273 B.n272 585
R31 B.n271 B.n270 585
R32 B.n269 B.n268 585
R33 B.n267 B.n266 585
R34 B.n265 B.n264 585
R35 B.n263 B.n262 585
R36 B.n261 B.n260 585
R37 B.n259 B.n258 585
R38 B.n257 B.n256 585
R39 B.n255 B.n254 585
R40 B.n253 B.n252 585
R41 B.n251 B.n250 585
R42 B.n249 B.n248 585
R43 B.n247 B.n246 585
R44 B.n245 B.n244 585
R45 B.n243 B.n242 585
R46 B.n241 B.n240 585
R47 B.n239 B.n238 585
R48 B.n237 B.n236 585
R49 B.n235 B.n234 585
R50 B.n233 B.n232 585
R51 B.n231 B.n230 585
R52 B.n229 B.n228 585
R53 B.n227 B.n226 585
R54 B.n225 B.n224 585
R55 B.n223 B.n222 585
R56 B.n221 B.n220 585
R57 B.n219 B.n218 585
R58 B.n217 B.n216 585
R59 B.n215 B.n214 585
R60 B.n213 B.n212 585
R61 B.n211 B.n210 585
R62 B.n209 B.n208 585
R63 B.n207 B.n206 585
R64 B.n205 B.n204 585
R65 B.n203 B.n202 585
R66 B.n201 B.n200 585
R67 B.n199 B.n198 585
R68 B.n197 B.n196 585
R69 B.n195 B.n194 585
R70 B.n193 B.n192 585
R71 B.n191 B.n190 585
R72 B.n189 B.n188 585
R73 B.n187 B.n186 585
R74 B.n185 B.n184 585
R75 B.n183 B.n182 585
R76 B.n181 B.n180 585
R77 B.n179 B.n178 585
R78 B.n177 B.n176 585
R79 B.n175 B.n174 585
R80 B.n173 B.n172 585
R81 B.n171 B.n170 585
R82 B.n169 B.n168 585
R83 B.n167 B.n166 585
R84 B.n165 B.n164 585
R85 B.n163 B.n162 585
R86 B.n161 B.n160 585
R87 B.n159 B.n158 585
R88 B.n157 B.n156 585
R89 B.n155 B.n154 585
R90 B.n153 B.n152 585
R91 B.n151 B.n150 585
R92 B.n149 B.n148 585
R93 B.n147 B.n146 585
R94 B.n145 B.n144 585
R95 B.n143 B.n142 585
R96 B.n141 B.n140 585
R97 B.n139 B.n138 585
R98 B.n137 B.n136 585
R99 B.n135 B.n134 585
R100 B.n133 B.n132 585
R101 B.n131 B.n130 585
R102 B.n129 B.n128 585
R103 B.n127 B.n126 585
R104 B.n125 B.n124 585
R105 B.n123 B.n122 585
R106 B.n121 B.n120 585
R107 B.n119 B.n118 585
R108 B.n117 B.n116 585
R109 B.n53 B.n52 585
R110 B.n784 B.n54 585
R111 B.n789 B.n54 585
R112 B.n783 B.n782 585
R113 B.n782 B.n50 585
R114 B.n781 B.n49 585
R115 B.n795 B.n49 585
R116 B.n780 B.n48 585
R117 B.n796 B.n48 585
R118 B.n779 B.n47 585
R119 B.n797 B.n47 585
R120 B.n778 B.n777 585
R121 B.n777 B.n43 585
R122 B.n776 B.n42 585
R123 B.n803 B.n42 585
R124 B.n775 B.n41 585
R125 B.n804 B.n41 585
R126 B.n774 B.n40 585
R127 B.n805 B.n40 585
R128 B.n773 B.n772 585
R129 B.n772 B.n36 585
R130 B.n771 B.n35 585
R131 B.n811 B.n35 585
R132 B.n770 B.n34 585
R133 B.n812 B.n34 585
R134 B.n769 B.n33 585
R135 B.n813 B.n33 585
R136 B.n768 B.n767 585
R137 B.n767 B.n29 585
R138 B.n766 B.n28 585
R139 B.n819 B.n28 585
R140 B.n765 B.n27 585
R141 B.n820 B.n27 585
R142 B.n764 B.n26 585
R143 B.n821 B.n26 585
R144 B.n763 B.n762 585
R145 B.n762 B.n22 585
R146 B.n761 B.n21 585
R147 B.n827 B.n21 585
R148 B.n760 B.n20 585
R149 B.n828 B.n20 585
R150 B.n759 B.n19 585
R151 B.n829 B.n19 585
R152 B.n758 B.n757 585
R153 B.n757 B.n18 585
R154 B.n756 B.n14 585
R155 B.n835 B.n14 585
R156 B.n755 B.n13 585
R157 B.n836 B.n13 585
R158 B.n754 B.n12 585
R159 B.n837 B.n12 585
R160 B.n753 B.n752 585
R161 B.n752 B.n8 585
R162 B.n751 B.n7 585
R163 B.n843 B.n7 585
R164 B.n750 B.n6 585
R165 B.n844 B.n6 585
R166 B.n749 B.n5 585
R167 B.n845 B.n5 585
R168 B.n748 B.n747 585
R169 B.n747 B.n4 585
R170 B.n746 B.n331 585
R171 B.n746 B.n745 585
R172 B.n736 B.n332 585
R173 B.n333 B.n332 585
R174 B.n738 B.n737 585
R175 B.n739 B.n738 585
R176 B.n735 B.n338 585
R177 B.n338 B.n337 585
R178 B.n734 B.n733 585
R179 B.n733 B.n732 585
R180 B.n340 B.n339 585
R181 B.n725 B.n340 585
R182 B.n724 B.n723 585
R183 B.n726 B.n724 585
R184 B.n722 B.n345 585
R185 B.n345 B.n344 585
R186 B.n721 B.n720 585
R187 B.n720 B.n719 585
R188 B.n347 B.n346 585
R189 B.n348 B.n347 585
R190 B.n712 B.n711 585
R191 B.n713 B.n712 585
R192 B.n710 B.n353 585
R193 B.n353 B.n352 585
R194 B.n709 B.n708 585
R195 B.n708 B.n707 585
R196 B.n355 B.n354 585
R197 B.n356 B.n355 585
R198 B.n700 B.n699 585
R199 B.n701 B.n700 585
R200 B.n698 B.n361 585
R201 B.n361 B.n360 585
R202 B.n697 B.n696 585
R203 B.n696 B.n695 585
R204 B.n363 B.n362 585
R205 B.n364 B.n363 585
R206 B.n688 B.n687 585
R207 B.n689 B.n688 585
R208 B.n686 B.n369 585
R209 B.n369 B.n368 585
R210 B.n685 B.n684 585
R211 B.n684 B.n683 585
R212 B.n371 B.n370 585
R213 B.n372 B.n371 585
R214 B.n676 B.n675 585
R215 B.n677 B.n676 585
R216 B.n674 B.n377 585
R217 B.n377 B.n376 585
R218 B.n673 B.n672 585
R219 B.n672 B.n671 585
R220 B.n379 B.n378 585
R221 B.n380 B.n379 585
R222 B.n664 B.n663 585
R223 B.n665 B.n664 585
R224 B.n383 B.n382 585
R225 B.n444 B.n442 585
R226 B.n445 B.n441 585
R227 B.n445 B.n384 585
R228 B.n448 B.n447 585
R229 B.n449 B.n440 585
R230 B.n451 B.n450 585
R231 B.n453 B.n439 585
R232 B.n456 B.n455 585
R233 B.n457 B.n438 585
R234 B.n459 B.n458 585
R235 B.n461 B.n437 585
R236 B.n464 B.n463 585
R237 B.n465 B.n436 585
R238 B.n467 B.n466 585
R239 B.n469 B.n435 585
R240 B.n472 B.n471 585
R241 B.n473 B.n434 585
R242 B.n475 B.n474 585
R243 B.n477 B.n433 585
R244 B.n480 B.n479 585
R245 B.n481 B.n432 585
R246 B.n483 B.n482 585
R247 B.n485 B.n431 585
R248 B.n488 B.n487 585
R249 B.n489 B.n430 585
R250 B.n491 B.n490 585
R251 B.n493 B.n429 585
R252 B.n496 B.n495 585
R253 B.n497 B.n428 585
R254 B.n499 B.n498 585
R255 B.n501 B.n427 585
R256 B.n504 B.n503 585
R257 B.n505 B.n426 585
R258 B.n507 B.n506 585
R259 B.n509 B.n425 585
R260 B.n512 B.n511 585
R261 B.n513 B.n424 585
R262 B.n515 B.n514 585
R263 B.n517 B.n423 585
R264 B.n520 B.n519 585
R265 B.n521 B.n422 585
R266 B.n523 B.n522 585
R267 B.n525 B.n421 585
R268 B.n528 B.n527 585
R269 B.n529 B.n420 585
R270 B.n531 B.n530 585
R271 B.n533 B.n419 585
R272 B.n536 B.n535 585
R273 B.n537 B.n418 585
R274 B.n542 B.n541 585
R275 B.n544 B.n417 585
R276 B.n547 B.n546 585
R277 B.n548 B.n416 585
R278 B.n550 B.n549 585
R279 B.n552 B.n415 585
R280 B.n555 B.n554 585
R281 B.n556 B.n414 585
R282 B.n558 B.n557 585
R283 B.n560 B.n413 585
R284 B.n563 B.n562 585
R285 B.n565 B.n410 585
R286 B.n567 B.n566 585
R287 B.n569 B.n409 585
R288 B.n572 B.n571 585
R289 B.n573 B.n408 585
R290 B.n575 B.n574 585
R291 B.n577 B.n407 585
R292 B.n580 B.n579 585
R293 B.n581 B.n406 585
R294 B.n583 B.n582 585
R295 B.n585 B.n405 585
R296 B.n588 B.n587 585
R297 B.n589 B.n404 585
R298 B.n591 B.n590 585
R299 B.n593 B.n403 585
R300 B.n596 B.n595 585
R301 B.n597 B.n402 585
R302 B.n599 B.n598 585
R303 B.n601 B.n401 585
R304 B.n604 B.n603 585
R305 B.n605 B.n400 585
R306 B.n607 B.n606 585
R307 B.n609 B.n399 585
R308 B.n612 B.n611 585
R309 B.n613 B.n398 585
R310 B.n615 B.n614 585
R311 B.n617 B.n397 585
R312 B.n620 B.n619 585
R313 B.n621 B.n396 585
R314 B.n623 B.n622 585
R315 B.n625 B.n395 585
R316 B.n628 B.n627 585
R317 B.n629 B.n394 585
R318 B.n631 B.n630 585
R319 B.n633 B.n393 585
R320 B.n636 B.n635 585
R321 B.n637 B.n392 585
R322 B.n639 B.n638 585
R323 B.n641 B.n391 585
R324 B.n644 B.n643 585
R325 B.n645 B.n390 585
R326 B.n647 B.n646 585
R327 B.n649 B.n389 585
R328 B.n652 B.n651 585
R329 B.n653 B.n388 585
R330 B.n655 B.n654 585
R331 B.n657 B.n387 585
R332 B.n658 B.n386 585
R333 B.n661 B.n660 585
R334 B.n662 B.n385 585
R335 B.n385 B.n384 585
R336 B.n667 B.n666 585
R337 B.n666 B.n665 585
R338 B.n668 B.n381 585
R339 B.n381 B.n380 585
R340 B.n670 B.n669 585
R341 B.n671 B.n670 585
R342 B.n375 B.n374 585
R343 B.n376 B.n375 585
R344 B.n679 B.n678 585
R345 B.n678 B.n677 585
R346 B.n680 B.n373 585
R347 B.n373 B.n372 585
R348 B.n682 B.n681 585
R349 B.n683 B.n682 585
R350 B.n367 B.n366 585
R351 B.n368 B.n367 585
R352 B.n691 B.n690 585
R353 B.n690 B.n689 585
R354 B.n692 B.n365 585
R355 B.n365 B.n364 585
R356 B.n694 B.n693 585
R357 B.n695 B.n694 585
R358 B.n359 B.n358 585
R359 B.n360 B.n359 585
R360 B.n703 B.n702 585
R361 B.n702 B.n701 585
R362 B.n704 B.n357 585
R363 B.n357 B.n356 585
R364 B.n706 B.n705 585
R365 B.n707 B.n706 585
R366 B.n351 B.n350 585
R367 B.n352 B.n351 585
R368 B.n715 B.n714 585
R369 B.n714 B.n713 585
R370 B.n716 B.n349 585
R371 B.n349 B.n348 585
R372 B.n718 B.n717 585
R373 B.n719 B.n718 585
R374 B.n343 B.n342 585
R375 B.n344 B.n343 585
R376 B.n728 B.n727 585
R377 B.n727 B.n726 585
R378 B.n729 B.n341 585
R379 B.n725 B.n341 585
R380 B.n731 B.n730 585
R381 B.n732 B.n731 585
R382 B.n336 B.n335 585
R383 B.n337 B.n336 585
R384 B.n741 B.n740 585
R385 B.n740 B.n739 585
R386 B.n742 B.n334 585
R387 B.n334 B.n333 585
R388 B.n744 B.n743 585
R389 B.n745 B.n744 585
R390 B.n2 B.n0 585
R391 B.n4 B.n2 585
R392 B.n3 B.n1 585
R393 B.n844 B.n3 585
R394 B.n842 B.n841 585
R395 B.n843 B.n842 585
R396 B.n840 B.n9 585
R397 B.n9 B.n8 585
R398 B.n839 B.n838 585
R399 B.n838 B.n837 585
R400 B.n11 B.n10 585
R401 B.n836 B.n11 585
R402 B.n834 B.n833 585
R403 B.n835 B.n834 585
R404 B.n832 B.n15 585
R405 B.n18 B.n15 585
R406 B.n831 B.n830 585
R407 B.n830 B.n829 585
R408 B.n17 B.n16 585
R409 B.n828 B.n17 585
R410 B.n826 B.n825 585
R411 B.n827 B.n826 585
R412 B.n824 B.n23 585
R413 B.n23 B.n22 585
R414 B.n823 B.n822 585
R415 B.n822 B.n821 585
R416 B.n25 B.n24 585
R417 B.n820 B.n25 585
R418 B.n818 B.n817 585
R419 B.n819 B.n818 585
R420 B.n816 B.n30 585
R421 B.n30 B.n29 585
R422 B.n815 B.n814 585
R423 B.n814 B.n813 585
R424 B.n32 B.n31 585
R425 B.n812 B.n32 585
R426 B.n810 B.n809 585
R427 B.n811 B.n810 585
R428 B.n808 B.n37 585
R429 B.n37 B.n36 585
R430 B.n807 B.n806 585
R431 B.n806 B.n805 585
R432 B.n39 B.n38 585
R433 B.n804 B.n39 585
R434 B.n802 B.n801 585
R435 B.n803 B.n802 585
R436 B.n800 B.n44 585
R437 B.n44 B.n43 585
R438 B.n799 B.n798 585
R439 B.n798 B.n797 585
R440 B.n46 B.n45 585
R441 B.n796 B.n46 585
R442 B.n794 B.n793 585
R443 B.n795 B.n794 585
R444 B.n792 B.n51 585
R445 B.n51 B.n50 585
R446 B.n791 B.n790 585
R447 B.n790 B.n789 585
R448 B.n847 B.n846 585
R449 B.n846 B.n845 585
R450 B.n666 B.n383 492.5
R451 B.n790 B.n53 492.5
R452 B.n664 B.n385 492.5
R453 B.n786 B.n54 492.5
R454 B.n411 B.t9 398.483
R455 B.n110 B.t4 398.483
R456 B.n538 B.t15 398.481
R457 B.n113 B.t11 398.481
R458 B.n412 B.t8 333.318
R459 B.n111 B.t5 333.318
R460 B.n539 B.t14 333.318
R461 B.n114 B.t12 333.318
R462 B.n411 B.t6 327.524
R463 B.n538 B.t13 327.524
R464 B.n113 B.t10 327.524
R465 B.n110 B.t2 327.524
R466 B.n788 B.n787 256.663
R467 B.n788 B.n108 256.663
R468 B.n788 B.n107 256.663
R469 B.n788 B.n106 256.663
R470 B.n788 B.n105 256.663
R471 B.n788 B.n104 256.663
R472 B.n788 B.n103 256.663
R473 B.n788 B.n102 256.663
R474 B.n788 B.n101 256.663
R475 B.n788 B.n100 256.663
R476 B.n788 B.n99 256.663
R477 B.n788 B.n98 256.663
R478 B.n788 B.n97 256.663
R479 B.n788 B.n96 256.663
R480 B.n788 B.n95 256.663
R481 B.n788 B.n94 256.663
R482 B.n788 B.n93 256.663
R483 B.n788 B.n92 256.663
R484 B.n788 B.n91 256.663
R485 B.n788 B.n90 256.663
R486 B.n788 B.n89 256.663
R487 B.n788 B.n88 256.663
R488 B.n788 B.n87 256.663
R489 B.n788 B.n86 256.663
R490 B.n788 B.n85 256.663
R491 B.n788 B.n84 256.663
R492 B.n788 B.n83 256.663
R493 B.n788 B.n82 256.663
R494 B.n788 B.n81 256.663
R495 B.n788 B.n80 256.663
R496 B.n788 B.n79 256.663
R497 B.n788 B.n78 256.663
R498 B.n788 B.n77 256.663
R499 B.n788 B.n76 256.663
R500 B.n788 B.n75 256.663
R501 B.n788 B.n74 256.663
R502 B.n788 B.n73 256.663
R503 B.n788 B.n72 256.663
R504 B.n788 B.n71 256.663
R505 B.n788 B.n70 256.663
R506 B.n788 B.n69 256.663
R507 B.n788 B.n68 256.663
R508 B.n788 B.n67 256.663
R509 B.n788 B.n66 256.663
R510 B.n788 B.n65 256.663
R511 B.n788 B.n64 256.663
R512 B.n788 B.n63 256.663
R513 B.n788 B.n62 256.663
R514 B.n788 B.n61 256.663
R515 B.n788 B.n60 256.663
R516 B.n788 B.n59 256.663
R517 B.n788 B.n58 256.663
R518 B.n788 B.n57 256.663
R519 B.n788 B.n56 256.663
R520 B.n788 B.n55 256.663
R521 B.n443 B.n384 256.663
R522 B.n446 B.n384 256.663
R523 B.n452 B.n384 256.663
R524 B.n454 B.n384 256.663
R525 B.n460 B.n384 256.663
R526 B.n462 B.n384 256.663
R527 B.n468 B.n384 256.663
R528 B.n470 B.n384 256.663
R529 B.n476 B.n384 256.663
R530 B.n478 B.n384 256.663
R531 B.n484 B.n384 256.663
R532 B.n486 B.n384 256.663
R533 B.n492 B.n384 256.663
R534 B.n494 B.n384 256.663
R535 B.n500 B.n384 256.663
R536 B.n502 B.n384 256.663
R537 B.n508 B.n384 256.663
R538 B.n510 B.n384 256.663
R539 B.n516 B.n384 256.663
R540 B.n518 B.n384 256.663
R541 B.n524 B.n384 256.663
R542 B.n526 B.n384 256.663
R543 B.n532 B.n384 256.663
R544 B.n534 B.n384 256.663
R545 B.n543 B.n384 256.663
R546 B.n545 B.n384 256.663
R547 B.n551 B.n384 256.663
R548 B.n553 B.n384 256.663
R549 B.n559 B.n384 256.663
R550 B.n561 B.n384 256.663
R551 B.n568 B.n384 256.663
R552 B.n570 B.n384 256.663
R553 B.n576 B.n384 256.663
R554 B.n578 B.n384 256.663
R555 B.n584 B.n384 256.663
R556 B.n586 B.n384 256.663
R557 B.n592 B.n384 256.663
R558 B.n594 B.n384 256.663
R559 B.n600 B.n384 256.663
R560 B.n602 B.n384 256.663
R561 B.n608 B.n384 256.663
R562 B.n610 B.n384 256.663
R563 B.n616 B.n384 256.663
R564 B.n618 B.n384 256.663
R565 B.n624 B.n384 256.663
R566 B.n626 B.n384 256.663
R567 B.n632 B.n384 256.663
R568 B.n634 B.n384 256.663
R569 B.n640 B.n384 256.663
R570 B.n642 B.n384 256.663
R571 B.n648 B.n384 256.663
R572 B.n650 B.n384 256.663
R573 B.n656 B.n384 256.663
R574 B.n659 B.n384 256.663
R575 B.n666 B.n381 163.367
R576 B.n670 B.n381 163.367
R577 B.n670 B.n375 163.367
R578 B.n678 B.n375 163.367
R579 B.n678 B.n373 163.367
R580 B.n682 B.n373 163.367
R581 B.n682 B.n367 163.367
R582 B.n690 B.n367 163.367
R583 B.n690 B.n365 163.367
R584 B.n694 B.n365 163.367
R585 B.n694 B.n359 163.367
R586 B.n702 B.n359 163.367
R587 B.n702 B.n357 163.367
R588 B.n706 B.n357 163.367
R589 B.n706 B.n351 163.367
R590 B.n714 B.n351 163.367
R591 B.n714 B.n349 163.367
R592 B.n718 B.n349 163.367
R593 B.n718 B.n343 163.367
R594 B.n727 B.n343 163.367
R595 B.n727 B.n341 163.367
R596 B.n731 B.n341 163.367
R597 B.n731 B.n336 163.367
R598 B.n740 B.n336 163.367
R599 B.n740 B.n334 163.367
R600 B.n744 B.n334 163.367
R601 B.n744 B.n2 163.367
R602 B.n846 B.n2 163.367
R603 B.n846 B.n3 163.367
R604 B.n842 B.n3 163.367
R605 B.n842 B.n9 163.367
R606 B.n838 B.n9 163.367
R607 B.n838 B.n11 163.367
R608 B.n834 B.n11 163.367
R609 B.n834 B.n15 163.367
R610 B.n830 B.n15 163.367
R611 B.n830 B.n17 163.367
R612 B.n826 B.n17 163.367
R613 B.n826 B.n23 163.367
R614 B.n822 B.n23 163.367
R615 B.n822 B.n25 163.367
R616 B.n818 B.n25 163.367
R617 B.n818 B.n30 163.367
R618 B.n814 B.n30 163.367
R619 B.n814 B.n32 163.367
R620 B.n810 B.n32 163.367
R621 B.n810 B.n37 163.367
R622 B.n806 B.n37 163.367
R623 B.n806 B.n39 163.367
R624 B.n802 B.n39 163.367
R625 B.n802 B.n44 163.367
R626 B.n798 B.n44 163.367
R627 B.n798 B.n46 163.367
R628 B.n794 B.n46 163.367
R629 B.n794 B.n51 163.367
R630 B.n790 B.n51 163.367
R631 B.n445 B.n444 163.367
R632 B.n447 B.n445 163.367
R633 B.n451 B.n440 163.367
R634 B.n455 B.n453 163.367
R635 B.n459 B.n438 163.367
R636 B.n463 B.n461 163.367
R637 B.n467 B.n436 163.367
R638 B.n471 B.n469 163.367
R639 B.n475 B.n434 163.367
R640 B.n479 B.n477 163.367
R641 B.n483 B.n432 163.367
R642 B.n487 B.n485 163.367
R643 B.n491 B.n430 163.367
R644 B.n495 B.n493 163.367
R645 B.n499 B.n428 163.367
R646 B.n503 B.n501 163.367
R647 B.n507 B.n426 163.367
R648 B.n511 B.n509 163.367
R649 B.n515 B.n424 163.367
R650 B.n519 B.n517 163.367
R651 B.n523 B.n422 163.367
R652 B.n527 B.n525 163.367
R653 B.n531 B.n420 163.367
R654 B.n535 B.n533 163.367
R655 B.n542 B.n418 163.367
R656 B.n546 B.n544 163.367
R657 B.n550 B.n416 163.367
R658 B.n554 B.n552 163.367
R659 B.n558 B.n414 163.367
R660 B.n562 B.n560 163.367
R661 B.n567 B.n410 163.367
R662 B.n571 B.n569 163.367
R663 B.n575 B.n408 163.367
R664 B.n579 B.n577 163.367
R665 B.n583 B.n406 163.367
R666 B.n587 B.n585 163.367
R667 B.n591 B.n404 163.367
R668 B.n595 B.n593 163.367
R669 B.n599 B.n402 163.367
R670 B.n603 B.n601 163.367
R671 B.n607 B.n400 163.367
R672 B.n611 B.n609 163.367
R673 B.n615 B.n398 163.367
R674 B.n619 B.n617 163.367
R675 B.n623 B.n396 163.367
R676 B.n627 B.n625 163.367
R677 B.n631 B.n394 163.367
R678 B.n635 B.n633 163.367
R679 B.n639 B.n392 163.367
R680 B.n643 B.n641 163.367
R681 B.n647 B.n390 163.367
R682 B.n651 B.n649 163.367
R683 B.n655 B.n388 163.367
R684 B.n658 B.n657 163.367
R685 B.n660 B.n385 163.367
R686 B.n664 B.n379 163.367
R687 B.n672 B.n379 163.367
R688 B.n672 B.n377 163.367
R689 B.n676 B.n377 163.367
R690 B.n676 B.n371 163.367
R691 B.n684 B.n371 163.367
R692 B.n684 B.n369 163.367
R693 B.n688 B.n369 163.367
R694 B.n688 B.n363 163.367
R695 B.n696 B.n363 163.367
R696 B.n696 B.n361 163.367
R697 B.n700 B.n361 163.367
R698 B.n700 B.n355 163.367
R699 B.n708 B.n355 163.367
R700 B.n708 B.n353 163.367
R701 B.n712 B.n353 163.367
R702 B.n712 B.n347 163.367
R703 B.n720 B.n347 163.367
R704 B.n720 B.n345 163.367
R705 B.n724 B.n345 163.367
R706 B.n724 B.n340 163.367
R707 B.n733 B.n340 163.367
R708 B.n733 B.n338 163.367
R709 B.n738 B.n338 163.367
R710 B.n738 B.n332 163.367
R711 B.n746 B.n332 163.367
R712 B.n747 B.n746 163.367
R713 B.n747 B.n5 163.367
R714 B.n6 B.n5 163.367
R715 B.n7 B.n6 163.367
R716 B.n752 B.n7 163.367
R717 B.n752 B.n12 163.367
R718 B.n13 B.n12 163.367
R719 B.n14 B.n13 163.367
R720 B.n757 B.n14 163.367
R721 B.n757 B.n19 163.367
R722 B.n20 B.n19 163.367
R723 B.n21 B.n20 163.367
R724 B.n762 B.n21 163.367
R725 B.n762 B.n26 163.367
R726 B.n27 B.n26 163.367
R727 B.n28 B.n27 163.367
R728 B.n767 B.n28 163.367
R729 B.n767 B.n33 163.367
R730 B.n34 B.n33 163.367
R731 B.n35 B.n34 163.367
R732 B.n772 B.n35 163.367
R733 B.n772 B.n40 163.367
R734 B.n41 B.n40 163.367
R735 B.n42 B.n41 163.367
R736 B.n777 B.n42 163.367
R737 B.n777 B.n47 163.367
R738 B.n48 B.n47 163.367
R739 B.n49 B.n48 163.367
R740 B.n782 B.n49 163.367
R741 B.n782 B.n54 163.367
R742 B.n118 B.n117 163.367
R743 B.n122 B.n121 163.367
R744 B.n126 B.n125 163.367
R745 B.n130 B.n129 163.367
R746 B.n134 B.n133 163.367
R747 B.n138 B.n137 163.367
R748 B.n142 B.n141 163.367
R749 B.n146 B.n145 163.367
R750 B.n150 B.n149 163.367
R751 B.n154 B.n153 163.367
R752 B.n158 B.n157 163.367
R753 B.n162 B.n161 163.367
R754 B.n166 B.n165 163.367
R755 B.n170 B.n169 163.367
R756 B.n174 B.n173 163.367
R757 B.n178 B.n177 163.367
R758 B.n182 B.n181 163.367
R759 B.n186 B.n185 163.367
R760 B.n190 B.n189 163.367
R761 B.n194 B.n193 163.367
R762 B.n198 B.n197 163.367
R763 B.n202 B.n201 163.367
R764 B.n206 B.n205 163.367
R765 B.n210 B.n209 163.367
R766 B.n214 B.n213 163.367
R767 B.n218 B.n217 163.367
R768 B.n222 B.n221 163.367
R769 B.n226 B.n225 163.367
R770 B.n230 B.n229 163.367
R771 B.n234 B.n233 163.367
R772 B.n238 B.n237 163.367
R773 B.n242 B.n241 163.367
R774 B.n246 B.n245 163.367
R775 B.n250 B.n249 163.367
R776 B.n254 B.n253 163.367
R777 B.n258 B.n257 163.367
R778 B.n262 B.n261 163.367
R779 B.n266 B.n265 163.367
R780 B.n270 B.n269 163.367
R781 B.n274 B.n273 163.367
R782 B.n278 B.n277 163.367
R783 B.n282 B.n281 163.367
R784 B.n286 B.n285 163.367
R785 B.n290 B.n289 163.367
R786 B.n294 B.n293 163.367
R787 B.n298 B.n297 163.367
R788 B.n302 B.n301 163.367
R789 B.n306 B.n305 163.367
R790 B.n310 B.n309 163.367
R791 B.n314 B.n313 163.367
R792 B.n318 B.n317 163.367
R793 B.n322 B.n321 163.367
R794 B.n326 B.n325 163.367
R795 B.n328 B.n109 163.367
R796 B.n443 B.n383 71.676
R797 B.n447 B.n446 71.676
R798 B.n452 B.n451 71.676
R799 B.n455 B.n454 71.676
R800 B.n460 B.n459 71.676
R801 B.n463 B.n462 71.676
R802 B.n468 B.n467 71.676
R803 B.n471 B.n470 71.676
R804 B.n476 B.n475 71.676
R805 B.n479 B.n478 71.676
R806 B.n484 B.n483 71.676
R807 B.n487 B.n486 71.676
R808 B.n492 B.n491 71.676
R809 B.n495 B.n494 71.676
R810 B.n500 B.n499 71.676
R811 B.n503 B.n502 71.676
R812 B.n508 B.n507 71.676
R813 B.n511 B.n510 71.676
R814 B.n516 B.n515 71.676
R815 B.n519 B.n518 71.676
R816 B.n524 B.n523 71.676
R817 B.n527 B.n526 71.676
R818 B.n532 B.n531 71.676
R819 B.n535 B.n534 71.676
R820 B.n543 B.n542 71.676
R821 B.n546 B.n545 71.676
R822 B.n551 B.n550 71.676
R823 B.n554 B.n553 71.676
R824 B.n559 B.n558 71.676
R825 B.n562 B.n561 71.676
R826 B.n568 B.n567 71.676
R827 B.n571 B.n570 71.676
R828 B.n576 B.n575 71.676
R829 B.n579 B.n578 71.676
R830 B.n584 B.n583 71.676
R831 B.n587 B.n586 71.676
R832 B.n592 B.n591 71.676
R833 B.n595 B.n594 71.676
R834 B.n600 B.n599 71.676
R835 B.n603 B.n602 71.676
R836 B.n608 B.n607 71.676
R837 B.n611 B.n610 71.676
R838 B.n616 B.n615 71.676
R839 B.n619 B.n618 71.676
R840 B.n624 B.n623 71.676
R841 B.n627 B.n626 71.676
R842 B.n632 B.n631 71.676
R843 B.n635 B.n634 71.676
R844 B.n640 B.n639 71.676
R845 B.n643 B.n642 71.676
R846 B.n648 B.n647 71.676
R847 B.n651 B.n650 71.676
R848 B.n656 B.n655 71.676
R849 B.n659 B.n658 71.676
R850 B.n55 B.n53 71.676
R851 B.n118 B.n56 71.676
R852 B.n122 B.n57 71.676
R853 B.n126 B.n58 71.676
R854 B.n130 B.n59 71.676
R855 B.n134 B.n60 71.676
R856 B.n138 B.n61 71.676
R857 B.n142 B.n62 71.676
R858 B.n146 B.n63 71.676
R859 B.n150 B.n64 71.676
R860 B.n154 B.n65 71.676
R861 B.n158 B.n66 71.676
R862 B.n162 B.n67 71.676
R863 B.n166 B.n68 71.676
R864 B.n170 B.n69 71.676
R865 B.n174 B.n70 71.676
R866 B.n178 B.n71 71.676
R867 B.n182 B.n72 71.676
R868 B.n186 B.n73 71.676
R869 B.n190 B.n74 71.676
R870 B.n194 B.n75 71.676
R871 B.n198 B.n76 71.676
R872 B.n202 B.n77 71.676
R873 B.n206 B.n78 71.676
R874 B.n210 B.n79 71.676
R875 B.n214 B.n80 71.676
R876 B.n218 B.n81 71.676
R877 B.n222 B.n82 71.676
R878 B.n226 B.n83 71.676
R879 B.n230 B.n84 71.676
R880 B.n234 B.n85 71.676
R881 B.n238 B.n86 71.676
R882 B.n242 B.n87 71.676
R883 B.n246 B.n88 71.676
R884 B.n250 B.n89 71.676
R885 B.n254 B.n90 71.676
R886 B.n258 B.n91 71.676
R887 B.n262 B.n92 71.676
R888 B.n266 B.n93 71.676
R889 B.n270 B.n94 71.676
R890 B.n274 B.n95 71.676
R891 B.n278 B.n96 71.676
R892 B.n282 B.n97 71.676
R893 B.n286 B.n98 71.676
R894 B.n290 B.n99 71.676
R895 B.n294 B.n100 71.676
R896 B.n298 B.n101 71.676
R897 B.n302 B.n102 71.676
R898 B.n306 B.n103 71.676
R899 B.n310 B.n104 71.676
R900 B.n314 B.n105 71.676
R901 B.n318 B.n106 71.676
R902 B.n322 B.n107 71.676
R903 B.n326 B.n108 71.676
R904 B.n787 B.n109 71.676
R905 B.n787 B.n786 71.676
R906 B.n328 B.n108 71.676
R907 B.n325 B.n107 71.676
R908 B.n321 B.n106 71.676
R909 B.n317 B.n105 71.676
R910 B.n313 B.n104 71.676
R911 B.n309 B.n103 71.676
R912 B.n305 B.n102 71.676
R913 B.n301 B.n101 71.676
R914 B.n297 B.n100 71.676
R915 B.n293 B.n99 71.676
R916 B.n289 B.n98 71.676
R917 B.n285 B.n97 71.676
R918 B.n281 B.n96 71.676
R919 B.n277 B.n95 71.676
R920 B.n273 B.n94 71.676
R921 B.n269 B.n93 71.676
R922 B.n265 B.n92 71.676
R923 B.n261 B.n91 71.676
R924 B.n257 B.n90 71.676
R925 B.n253 B.n89 71.676
R926 B.n249 B.n88 71.676
R927 B.n245 B.n87 71.676
R928 B.n241 B.n86 71.676
R929 B.n237 B.n85 71.676
R930 B.n233 B.n84 71.676
R931 B.n229 B.n83 71.676
R932 B.n225 B.n82 71.676
R933 B.n221 B.n81 71.676
R934 B.n217 B.n80 71.676
R935 B.n213 B.n79 71.676
R936 B.n209 B.n78 71.676
R937 B.n205 B.n77 71.676
R938 B.n201 B.n76 71.676
R939 B.n197 B.n75 71.676
R940 B.n193 B.n74 71.676
R941 B.n189 B.n73 71.676
R942 B.n185 B.n72 71.676
R943 B.n181 B.n71 71.676
R944 B.n177 B.n70 71.676
R945 B.n173 B.n69 71.676
R946 B.n169 B.n68 71.676
R947 B.n165 B.n67 71.676
R948 B.n161 B.n66 71.676
R949 B.n157 B.n65 71.676
R950 B.n153 B.n64 71.676
R951 B.n149 B.n63 71.676
R952 B.n145 B.n62 71.676
R953 B.n141 B.n61 71.676
R954 B.n137 B.n60 71.676
R955 B.n133 B.n59 71.676
R956 B.n129 B.n58 71.676
R957 B.n125 B.n57 71.676
R958 B.n121 B.n56 71.676
R959 B.n117 B.n55 71.676
R960 B.n444 B.n443 71.676
R961 B.n446 B.n440 71.676
R962 B.n453 B.n452 71.676
R963 B.n454 B.n438 71.676
R964 B.n461 B.n460 71.676
R965 B.n462 B.n436 71.676
R966 B.n469 B.n468 71.676
R967 B.n470 B.n434 71.676
R968 B.n477 B.n476 71.676
R969 B.n478 B.n432 71.676
R970 B.n485 B.n484 71.676
R971 B.n486 B.n430 71.676
R972 B.n493 B.n492 71.676
R973 B.n494 B.n428 71.676
R974 B.n501 B.n500 71.676
R975 B.n502 B.n426 71.676
R976 B.n509 B.n508 71.676
R977 B.n510 B.n424 71.676
R978 B.n517 B.n516 71.676
R979 B.n518 B.n422 71.676
R980 B.n525 B.n524 71.676
R981 B.n526 B.n420 71.676
R982 B.n533 B.n532 71.676
R983 B.n534 B.n418 71.676
R984 B.n544 B.n543 71.676
R985 B.n545 B.n416 71.676
R986 B.n552 B.n551 71.676
R987 B.n553 B.n414 71.676
R988 B.n560 B.n559 71.676
R989 B.n561 B.n410 71.676
R990 B.n569 B.n568 71.676
R991 B.n570 B.n408 71.676
R992 B.n577 B.n576 71.676
R993 B.n578 B.n406 71.676
R994 B.n585 B.n584 71.676
R995 B.n586 B.n404 71.676
R996 B.n593 B.n592 71.676
R997 B.n594 B.n402 71.676
R998 B.n601 B.n600 71.676
R999 B.n602 B.n400 71.676
R1000 B.n609 B.n608 71.676
R1001 B.n610 B.n398 71.676
R1002 B.n617 B.n616 71.676
R1003 B.n618 B.n396 71.676
R1004 B.n625 B.n624 71.676
R1005 B.n626 B.n394 71.676
R1006 B.n633 B.n632 71.676
R1007 B.n634 B.n392 71.676
R1008 B.n641 B.n640 71.676
R1009 B.n642 B.n390 71.676
R1010 B.n649 B.n648 71.676
R1011 B.n650 B.n388 71.676
R1012 B.n657 B.n656 71.676
R1013 B.n660 B.n659 71.676
R1014 B.n412 B.n411 65.1641
R1015 B.n539 B.n538 65.1641
R1016 B.n114 B.n113 65.1641
R1017 B.n111 B.n110 65.1641
R1018 B.n665 B.n384 62.5469
R1019 B.n789 B.n788 62.5469
R1020 B.n564 B.n412 59.5399
R1021 B.n540 B.n539 59.5399
R1022 B.n115 B.n114 59.5399
R1023 B.n112 B.n111 59.5399
R1024 B.n665 B.n380 36.9844
R1025 B.n671 B.n380 36.9844
R1026 B.n671 B.n376 36.9844
R1027 B.n677 B.n376 36.9844
R1028 B.n677 B.n372 36.9844
R1029 B.n683 B.n372 36.9844
R1030 B.n683 B.n368 36.9844
R1031 B.n689 B.n368 36.9844
R1032 B.n695 B.n364 36.9844
R1033 B.n695 B.n360 36.9844
R1034 B.n701 B.n360 36.9844
R1035 B.n701 B.n356 36.9844
R1036 B.n707 B.n356 36.9844
R1037 B.n707 B.n352 36.9844
R1038 B.n713 B.n352 36.9844
R1039 B.n713 B.n348 36.9844
R1040 B.n719 B.n348 36.9844
R1041 B.n719 B.n344 36.9844
R1042 B.n726 B.n344 36.9844
R1043 B.n726 B.n725 36.9844
R1044 B.n732 B.n337 36.9844
R1045 B.n739 B.n337 36.9844
R1046 B.n739 B.n333 36.9844
R1047 B.n745 B.n333 36.9844
R1048 B.n745 B.n4 36.9844
R1049 B.n845 B.n4 36.9844
R1050 B.n845 B.n844 36.9844
R1051 B.n844 B.n843 36.9844
R1052 B.n843 B.n8 36.9844
R1053 B.n837 B.n8 36.9844
R1054 B.n837 B.n836 36.9844
R1055 B.n836 B.n835 36.9844
R1056 B.n829 B.n18 36.9844
R1057 B.n829 B.n828 36.9844
R1058 B.n828 B.n827 36.9844
R1059 B.n827 B.n22 36.9844
R1060 B.n821 B.n22 36.9844
R1061 B.n821 B.n820 36.9844
R1062 B.n820 B.n819 36.9844
R1063 B.n819 B.n29 36.9844
R1064 B.n813 B.n29 36.9844
R1065 B.n813 B.n812 36.9844
R1066 B.n812 B.n811 36.9844
R1067 B.n811 B.n36 36.9844
R1068 B.n805 B.n804 36.9844
R1069 B.n804 B.n803 36.9844
R1070 B.n803 B.n43 36.9844
R1071 B.n797 B.n43 36.9844
R1072 B.n797 B.n796 36.9844
R1073 B.n796 B.n795 36.9844
R1074 B.n795 B.n50 36.9844
R1075 B.n789 B.n50 36.9844
R1076 B.n791 B.n52 32.0005
R1077 B.n785 B.n784 32.0005
R1078 B.n663 B.n662 32.0005
R1079 B.n667 B.n382 32.0005
R1080 B.t7 B.n364 23.3874
R1081 B.t3 B.n36 23.3874
R1082 B.n732 B.t0 20.1241
R1083 B.n835 B.t1 20.1241
R1084 B B.n847 18.0485
R1085 B.n725 B.t0 16.8608
R1086 B.n18 B.t1 16.8608
R1087 B.n689 B.t7 13.5975
R1088 B.n805 B.t3 13.5975
R1089 B.n116 B.n52 10.6151
R1090 B.n119 B.n116 10.6151
R1091 B.n120 B.n119 10.6151
R1092 B.n123 B.n120 10.6151
R1093 B.n124 B.n123 10.6151
R1094 B.n127 B.n124 10.6151
R1095 B.n128 B.n127 10.6151
R1096 B.n131 B.n128 10.6151
R1097 B.n132 B.n131 10.6151
R1098 B.n135 B.n132 10.6151
R1099 B.n136 B.n135 10.6151
R1100 B.n139 B.n136 10.6151
R1101 B.n140 B.n139 10.6151
R1102 B.n143 B.n140 10.6151
R1103 B.n144 B.n143 10.6151
R1104 B.n147 B.n144 10.6151
R1105 B.n148 B.n147 10.6151
R1106 B.n151 B.n148 10.6151
R1107 B.n152 B.n151 10.6151
R1108 B.n155 B.n152 10.6151
R1109 B.n156 B.n155 10.6151
R1110 B.n159 B.n156 10.6151
R1111 B.n160 B.n159 10.6151
R1112 B.n163 B.n160 10.6151
R1113 B.n164 B.n163 10.6151
R1114 B.n167 B.n164 10.6151
R1115 B.n168 B.n167 10.6151
R1116 B.n171 B.n168 10.6151
R1117 B.n172 B.n171 10.6151
R1118 B.n175 B.n172 10.6151
R1119 B.n176 B.n175 10.6151
R1120 B.n179 B.n176 10.6151
R1121 B.n180 B.n179 10.6151
R1122 B.n183 B.n180 10.6151
R1123 B.n184 B.n183 10.6151
R1124 B.n187 B.n184 10.6151
R1125 B.n188 B.n187 10.6151
R1126 B.n191 B.n188 10.6151
R1127 B.n192 B.n191 10.6151
R1128 B.n195 B.n192 10.6151
R1129 B.n196 B.n195 10.6151
R1130 B.n199 B.n196 10.6151
R1131 B.n200 B.n199 10.6151
R1132 B.n203 B.n200 10.6151
R1133 B.n204 B.n203 10.6151
R1134 B.n207 B.n204 10.6151
R1135 B.n208 B.n207 10.6151
R1136 B.n211 B.n208 10.6151
R1137 B.n212 B.n211 10.6151
R1138 B.n216 B.n215 10.6151
R1139 B.n219 B.n216 10.6151
R1140 B.n220 B.n219 10.6151
R1141 B.n223 B.n220 10.6151
R1142 B.n224 B.n223 10.6151
R1143 B.n227 B.n224 10.6151
R1144 B.n228 B.n227 10.6151
R1145 B.n231 B.n228 10.6151
R1146 B.n232 B.n231 10.6151
R1147 B.n236 B.n235 10.6151
R1148 B.n239 B.n236 10.6151
R1149 B.n240 B.n239 10.6151
R1150 B.n243 B.n240 10.6151
R1151 B.n244 B.n243 10.6151
R1152 B.n247 B.n244 10.6151
R1153 B.n248 B.n247 10.6151
R1154 B.n251 B.n248 10.6151
R1155 B.n252 B.n251 10.6151
R1156 B.n255 B.n252 10.6151
R1157 B.n256 B.n255 10.6151
R1158 B.n259 B.n256 10.6151
R1159 B.n260 B.n259 10.6151
R1160 B.n263 B.n260 10.6151
R1161 B.n264 B.n263 10.6151
R1162 B.n267 B.n264 10.6151
R1163 B.n268 B.n267 10.6151
R1164 B.n271 B.n268 10.6151
R1165 B.n272 B.n271 10.6151
R1166 B.n275 B.n272 10.6151
R1167 B.n276 B.n275 10.6151
R1168 B.n279 B.n276 10.6151
R1169 B.n280 B.n279 10.6151
R1170 B.n283 B.n280 10.6151
R1171 B.n284 B.n283 10.6151
R1172 B.n287 B.n284 10.6151
R1173 B.n288 B.n287 10.6151
R1174 B.n291 B.n288 10.6151
R1175 B.n292 B.n291 10.6151
R1176 B.n295 B.n292 10.6151
R1177 B.n296 B.n295 10.6151
R1178 B.n299 B.n296 10.6151
R1179 B.n300 B.n299 10.6151
R1180 B.n303 B.n300 10.6151
R1181 B.n304 B.n303 10.6151
R1182 B.n307 B.n304 10.6151
R1183 B.n308 B.n307 10.6151
R1184 B.n311 B.n308 10.6151
R1185 B.n312 B.n311 10.6151
R1186 B.n315 B.n312 10.6151
R1187 B.n316 B.n315 10.6151
R1188 B.n319 B.n316 10.6151
R1189 B.n320 B.n319 10.6151
R1190 B.n323 B.n320 10.6151
R1191 B.n324 B.n323 10.6151
R1192 B.n327 B.n324 10.6151
R1193 B.n329 B.n327 10.6151
R1194 B.n330 B.n329 10.6151
R1195 B.n785 B.n330 10.6151
R1196 B.n663 B.n378 10.6151
R1197 B.n673 B.n378 10.6151
R1198 B.n674 B.n673 10.6151
R1199 B.n675 B.n674 10.6151
R1200 B.n675 B.n370 10.6151
R1201 B.n685 B.n370 10.6151
R1202 B.n686 B.n685 10.6151
R1203 B.n687 B.n686 10.6151
R1204 B.n687 B.n362 10.6151
R1205 B.n697 B.n362 10.6151
R1206 B.n698 B.n697 10.6151
R1207 B.n699 B.n698 10.6151
R1208 B.n699 B.n354 10.6151
R1209 B.n709 B.n354 10.6151
R1210 B.n710 B.n709 10.6151
R1211 B.n711 B.n710 10.6151
R1212 B.n711 B.n346 10.6151
R1213 B.n721 B.n346 10.6151
R1214 B.n722 B.n721 10.6151
R1215 B.n723 B.n722 10.6151
R1216 B.n723 B.n339 10.6151
R1217 B.n734 B.n339 10.6151
R1218 B.n735 B.n734 10.6151
R1219 B.n737 B.n735 10.6151
R1220 B.n737 B.n736 10.6151
R1221 B.n736 B.n331 10.6151
R1222 B.n748 B.n331 10.6151
R1223 B.n749 B.n748 10.6151
R1224 B.n750 B.n749 10.6151
R1225 B.n751 B.n750 10.6151
R1226 B.n753 B.n751 10.6151
R1227 B.n754 B.n753 10.6151
R1228 B.n755 B.n754 10.6151
R1229 B.n756 B.n755 10.6151
R1230 B.n758 B.n756 10.6151
R1231 B.n759 B.n758 10.6151
R1232 B.n760 B.n759 10.6151
R1233 B.n761 B.n760 10.6151
R1234 B.n763 B.n761 10.6151
R1235 B.n764 B.n763 10.6151
R1236 B.n765 B.n764 10.6151
R1237 B.n766 B.n765 10.6151
R1238 B.n768 B.n766 10.6151
R1239 B.n769 B.n768 10.6151
R1240 B.n770 B.n769 10.6151
R1241 B.n771 B.n770 10.6151
R1242 B.n773 B.n771 10.6151
R1243 B.n774 B.n773 10.6151
R1244 B.n775 B.n774 10.6151
R1245 B.n776 B.n775 10.6151
R1246 B.n778 B.n776 10.6151
R1247 B.n779 B.n778 10.6151
R1248 B.n780 B.n779 10.6151
R1249 B.n781 B.n780 10.6151
R1250 B.n783 B.n781 10.6151
R1251 B.n784 B.n783 10.6151
R1252 B.n442 B.n382 10.6151
R1253 B.n442 B.n441 10.6151
R1254 B.n448 B.n441 10.6151
R1255 B.n449 B.n448 10.6151
R1256 B.n450 B.n449 10.6151
R1257 B.n450 B.n439 10.6151
R1258 B.n456 B.n439 10.6151
R1259 B.n457 B.n456 10.6151
R1260 B.n458 B.n457 10.6151
R1261 B.n458 B.n437 10.6151
R1262 B.n464 B.n437 10.6151
R1263 B.n465 B.n464 10.6151
R1264 B.n466 B.n465 10.6151
R1265 B.n466 B.n435 10.6151
R1266 B.n472 B.n435 10.6151
R1267 B.n473 B.n472 10.6151
R1268 B.n474 B.n473 10.6151
R1269 B.n474 B.n433 10.6151
R1270 B.n480 B.n433 10.6151
R1271 B.n481 B.n480 10.6151
R1272 B.n482 B.n481 10.6151
R1273 B.n482 B.n431 10.6151
R1274 B.n488 B.n431 10.6151
R1275 B.n489 B.n488 10.6151
R1276 B.n490 B.n489 10.6151
R1277 B.n490 B.n429 10.6151
R1278 B.n496 B.n429 10.6151
R1279 B.n497 B.n496 10.6151
R1280 B.n498 B.n497 10.6151
R1281 B.n498 B.n427 10.6151
R1282 B.n504 B.n427 10.6151
R1283 B.n505 B.n504 10.6151
R1284 B.n506 B.n505 10.6151
R1285 B.n506 B.n425 10.6151
R1286 B.n512 B.n425 10.6151
R1287 B.n513 B.n512 10.6151
R1288 B.n514 B.n513 10.6151
R1289 B.n514 B.n423 10.6151
R1290 B.n520 B.n423 10.6151
R1291 B.n521 B.n520 10.6151
R1292 B.n522 B.n521 10.6151
R1293 B.n522 B.n421 10.6151
R1294 B.n528 B.n421 10.6151
R1295 B.n529 B.n528 10.6151
R1296 B.n530 B.n529 10.6151
R1297 B.n530 B.n419 10.6151
R1298 B.n536 B.n419 10.6151
R1299 B.n537 B.n536 10.6151
R1300 B.n541 B.n537 10.6151
R1301 B.n547 B.n417 10.6151
R1302 B.n548 B.n547 10.6151
R1303 B.n549 B.n548 10.6151
R1304 B.n549 B.n415 10.6151
R1305 B.n555 B.n415 10.6151
R1306 B.n556 B.n555 10.6151
R1307 B.n557 B.n556 10.6151
R1308 B.n557 B.n413 10.6151
R1309 B.n563 B.n413 10.6151
R1310 B.n566 B.n565 10.6151
R1311 B.n566 B.n409 10.6151
R1312 B.n572 B.n409 10.6151
R1313 B.n573 B.n572 10.6151
R1314 B.n574 B.n573 10.6151
R1315 B.n574 B.n407 10.6151
R1316 B.n580 B.n407 10.6151
R1317 B.n581 B.n580 10.6151
R1318 B.n582 B.n581 10.6151
R1319 B.n582 B.n405 10.6151
R1320 B.n588 B.n405 10.6151
R1321 B.n589 B.n588 10.6151
R1322 B.n590 B.n589 10.6151
R1323 B.n590 B.n403 10.6151
R1324 B.n596 B.n403 10.6151
R1325 B.n597 B.n596 10.6151
R1326 B.n598 B.n597 10.6151
R1327 B.n598 B.n401 10.6151
R1328 B.n604 B.n401 10.6151
R1329 B.n605 B.n604 10.6151
R1330 B.n606 B.n605 10.6151
R1331 B.n606 B.n399 10.6151
R1332 B.n612 B.n399 10.6151
R1333 B.n613 B.n612 10.6151
R1334 B.n614 B.n613 10.6151
R1335 B.n614 B.n397 10.6151
R1336 B.n620 B.n397 10.6151
R1337 B.n621 B.n620 10.6151
R1338 B.n622 B.n621 10.6151
R1339 B.n622 B.n395 10.6151
R1340 B.n628 B.n395 10.6151
R1341 B.n629 B.n628 10.6151
R1342 B.n630 B.n629 10.6151
R1343 B.n630 B.n393 10.6151
R1344 B.n636 B.n393 10.6151
R1345 B.n637 B.n636 10.6151
R1346 B.n638 B.n637 10.6151
R1347 B.n638 B.n391 10.6151
R1348 B.n644 B.n391 10.6151
R1349 B.n645 B.n644 10.6151
R1350 B.n646 B.n645 10.6151
R1351 B.n646 B.n389 10.6151
R1352 B.n652 B.n389 10.6151
R1353 B.n653 B.n652 10.6151
R1354 B.n654 B.n653 10.6151
R1355 B.n654 B.n387 10.6151
R1356 B.n387 B.n386 10.6151
R1357 B.n661 B.n386 10.6151
R1358 B.n662 B.n661 10.6151
R1359 B.n668 B.n667 10.6151
R1360 B.n669 B.n668 10.6151
R1361 B.n669 B.n374 10.6151
R1362 B.n679 B.n374 10.6151
R1363 B.n680 B.n679 10.6151
R1364 B.n681 B.n680 10.6151
R1365 B.n681 B.n366 10.6151
R1366 B.n691 B.n366 10.6151
R1367 B.n692 B.n691 10.6151
R1368 B.n693 B.n692 10.6151
R1369 B.n693 B.n358 10.6151
R1370 B.n703 B.n358 10.6151
R1371 B.n704 B.n703 10.6151
R1372 B.n705 B.n704 10.6151
R1373 B.n705 B.n350 10.6151
R1374 B.n715 B.n350 10.6151
R1375 B.n716 B.n715 10.6151
R1376 B.n717 B.n716 10.6151
R1377 B.n717 B.n342 10.6151
R1378 B.n728 B.n342 10.6151
R1379 B.n729 B.n728 10.6151
R1380 B.n730 B.n729 10.6151
R1381 B.n730 B.n335 10.6151
R1382 B.n741 B.n335 10.6151
R1383 B.n742 B.n741 10.6151
R1384 B.n743 B.n742 10.6151
R1385 B.n743 B.n0 10.6151
R1386 B.n841 B.n1 10.6151
R1387 B.n841 B.n840 10.6151
R1388 B.n840 B.n839 10.6151
R1389 B.n839 B.n10 10.6151
R1390 B.n833 B.n10 10.6151
R1391 B.n833 B.n832 10.6151
R1392 B.n832 B.n831 10.6151
R1393 B.n831 B.n16 10.6151
R1394 B.n825 B.n16 10.6151
R1395 B.n825 B.n824 10.6151
R1396 B.n824 B.n823 10.6151
R1397 B.n823 B.n24 10.6151
R1398 B.n817 B.n24 10.6151
R1399 B.n817 B.n816 10.6151
R1400 B.n816 B.n815 10.6151
R1401 B.n815 B.n31 10.6151
R1402 B.n809 B.n31 10.6151
R1403 B.n809 B.n808 10.6151
R1404 B.n808 B.n807 10.6151
R1405 B.n807 B.n38 10.6151
R1406 B.n801 B.n38 10.6151
R1407 B.n801 B.n800 10.6151
R1408 B.n800 B.n799 10.6151
R1409 B.n799 B.n45 10.6151
R1410 B.n793 B.n45 10.6151
R1411 B.n793 B.n792 10.6151
R1412 B.n792 B.n791 10.6151
R1413 B.n212 B.n115 9.36635
R1414 B.n235 B.n112 9.36635
R1415 B.n541 B.n540 9.36635
R1416 B.n565 B.n564 9.36635
R1417 B.n847 B.n0 2.81026
R1418 B.n847 B.n1 2.81026
R1419 B.n215 B.n115 1.24928
R1420 B.n232 B.n112 1.24928
R1421 B.n540 B.n417 1.24928
R1422 B.n564 B.n563 1.24928
R1423 VN VN.t1 208.04
R1424 VN VN.t0 160.436
R1425 VTAIL.n322 VTAIL.n246 289.615
R1426 VTAIL.n76 VTAIL.n0 289.615
R1427 VTAIL.n240 VTAIL.n164 289.615
R1428 VTAIL.n158 VTAIL.n82 289.615
R1429 VTAIL.n273 VTAIL.n272 185
R1430 VTAIL.n270 VTAIL.n269 185
R1431 VTAIL.n279 VTAIL.n278 185
R1432 VTAIL.n281 VTAIL.n280 185
R1433 VTAIL.n266 VTAIL.n265 185
R1434 VTAIL.n287 VTAIL.n286 185
R1435 VTAIL.n290 VTAIL.n289 185
R1436 VTAIL.n288 VTAIL.n262 185
R1437 VTAIL.n295 VTAIL.n261 185
R1438 VTAIL.n297 VTAIL.n296 185
R1439 VTAIL.n299 VTAIL.n298 185
R1440 VTAIL.n258 VTAIL.n257 185
R1441 VTAIL.n305 VTAIL.n304 185
R1442 VTAIL.n307 VTAIL.n306 185
R1443 VTAIL.n254 VTAIL.n253 185
R1444 VTAIL.n313 VTAIL.n312 185
R1445 VTAIL.n315 VTAIL.n314 185
R1446 VTAIL.n250 VTAIL.n249 185
R1447 VTAIL.n321 VTAIL.n320 185
R1448 VTAIL.n323 VTAIL.n322 185
R1449 VTAIL.n27 VTAIL.n26 185
R1450 VTAIL.n24 VTAIL.n23 185
R1451 VTAIL.n33 VTAIL.n32 185
R1452 VTAIL.n35 VTAIL.n34 185
R1453 VTAIL.n20 VTAIL.n19 185
R1454 VTAIL.n41 VTAIL.n40 185
R1455 VTAIL.n44 VTAIL.n43 185
R1456 VTAIL.n42 VTAIL.n16 185
R1457 VTAIL.n49 VTAIL.n15 185
R1458 VTAIL.n51 VTAIL.n50 185
R1459 VTAIL.n53 VTAIL.n52 185
R1460 VTAIL.n12 VTAIL.n11 185
R1461 VTAIL.n59 VTAIL.n58 185
R1462 VTAIL.n61 VTAIL.n60 185
R1463 VTAIL.n8 VTAIL.n7 185
R1464 VTAIL.n67 VTAIL.n66 185
R1465 VTAIL.n69 VTAIL.n68 185
R1466 VTAIL.n4 VTAIL.n3 185
R1467 VTAIL.n75 VTAIL.n74 185
R1468 VTAIL.n77 VTAIL.n76 185
R1469 VTAIL.n241 VTAIL.n240 185
R1470 VTAIL.n239 VTAIL.n238 185
R1471 VTAIL.n168 VTAIL.n167 185
R1472 VTAIL.n233 VTAIL.n232 185
R1473 VTAIL.n231 VTAIL.n230 185
R1474 VTAIL.n172 VTAIL.n171 185
R1475 VTAIL.n225 VTAIL.n224 185
R1476 VTAIL.n223 VTAIL.n222 185
R1477 VTAIL.n176 VTAIL.n175 185
R1478 VTAIL.n217 VTAIL.n216 185
R1479 VTAIL.n215 VTAIL.n214 185
R1480 VTAIL.n213 VTAIL.n179 185
R1481 VTAIL.n183 VTAIL.n180 185
R1482 VTAIL.n208 VTAIL.n207 185
R1483 VTAIL.n206 VTAIL.n205 185
R1484 VTAIL.n185 VTAIL.n184 185
R1485 VTAIL.n200 VTAIL.n199 185
R1486 VTAIL.n198 VTAIL.n197 185
R1487 VTAIL.n189 VTAIL.n188 185
R1488 VTAIL.n192 VTAIL.n191 185
R1489 VTAIL.n159 VTAIL.n158 185
R1490 VTAIL.n157 VTAIL.n156 185
R1491 VTAIL.n86 VTAIL.n85 185
R1492 VTAIL.n151 VTAIL.n150 185
R1493 VTAIL.n149 VTAIL.n148 185
R1494 VTAIL.n90 VTAIL.n89 185
R1495 VTAIL.n143 VTAIL.n142 185
R1496 VTAIL.n141 VTAIL.n140 185
R1497 VTAIL.n94 VTAIL.n93 185
R1498 VTAIL.n135 VTAIL.n134 185
R1499 VTAIL.n133 VTAIL.n132 185
R1500 VTAIL.n131 VTAIL.n97 185
R1501 VTAIL.n101 VTAIL.n98 185
R1502 VTAIL.n126 VTAIL.n125 185
R1503 VTAIL.n124 VTAIL.n123 185
R1504 VTAIL.n103 VTAIL.n102 185
R1505 VTAIL.n118 VTAIL.n117 185
R1506 VTAIL.n116 VTAIL.n115 185
R1507 VTAIL.n107 VTAIL.n106 185
R1508 VTAIL.n110 VTAIL.n109 185
R1509 VTAIL.t3 VTAIL.n271 149.524
R1510 VTAIL.t1 VTAIL.n25 149.524
R1511 VTAIL.t0 VTAIL.n190 149.524
R1512 VTAIL.t2 VTAIL.n108 149.524
R1513 VTAIL.n272 VTAIL.n269 104.615
R1514 VTAIL.n279 VTAIL.n269 104.615
R1515 VTAIL.n280 VTAIL.n279 104.615
R1516 VTAIL.n280 VTAIL.n265 104.615
R1517 VTAIL.n287 VTAIL.n265 104.615
R1518 VTAIL.n289 VTAIL.n287 104.615
R1519 VTAIL.n289 VTAIL.n288 104.615
R1520 VTAIL.n288 VTAIL.n261 104.615
R1521 VTAIL.n297 VTAIL.n261 104.615
R1522 VTAIL.n298 VTAIL.n297 104.615
R1523 VTAIL.n298 VTAIL.n257 104.615
R1524 VTAIL.n305 VTAIL.n257 104.615
R1525 VTAIL.n306 VTAIL.n305 104.615
R1526 VTAIL.n306 VTAIL.n253 104.615
R1527 VTAIL.n313 VTAIL.n253 104.615
R1528 VTAIL.n314 VTAIL.n313 104.615
R1529 VTAIL.n314 VTAIL.n249 104.615
R1530 VTAIL.n321 VTAIL.n249 104.615
R1531 VTAIL.n322 VTAIL.n321 104.615
R1532 VTAIL.n26 VTAIL.n23 104.615
R1533 VTAIL.n33 VTAIL.n23 104.615
R1534 VTAIL.n34 VTAIL.n33 104.615
R1535 VTAIL.n34 VTAIL.n19 104.615
R1536 VTAIL.n41 VTAIL.n19 104.615
R1537 VTAIL.n43 VTAIL.n41 104.615
R1538 VTAIL.n43 VTAIL.n42 104.615
R1539 VTAIL.n42 VTAIL.n15 104.615
R1540 VTAIL.n51 VTAIL.n15 104.615
R1541 VTAIL.n52 VTAIL.n51 104.615
R1542 VTAIL.n52 VTAIL.n11 104.615
R1543 VTAIL.n59 VTAIL.n11 104.615
R1544 VTAIL.n60 VTAIL.n59 104.615
R1545 VTAIL.n60 VTAIL.n7 104.615
R1546 VTAIL.n67 VTAIL.n7 104.615
R1547 VTAIL.n68 VTAIL.n67 104.615
R1548 VTAIL.n68 VTAIL.n3 104.615
R1549 VTAIL.n75 VTAIL.n3 104.615
R1550 VTAIL.n76 VTAIL.n75 104.615
R1551 VTAIL.n240 VTAIL.n239 104.615
R1552 VTAIL.n239 VTAIL.n167 104.615
R1553 VTAIL.n232 VTAIL.n167 104.615
R1554 VTAIL.n232 VTAIL.n231 104.615
R1555 VTAIL.n231 VTAIL.n171 104.615
R1556 VTAIL.n224 VTAIL.n171 104.615
R1557 VTAIL.n224 VTAIL.n223 104.615
R1558 VTAIL.n223 VTAIL.n175 104.615
R1559 VTAIL.n216 VTAIL.n175 104.615
R1560 VTAIL.n216 VTAIL.n215 104.615
R1561 VTAIL.n215 VTAIL.n179 104.615
R1562 VTAIL.n183 VTAIL.n179 104.615
R1563 VTAIL.n207 VTAIL.n183 104.615
R1564 VTAIL.n207 VTAIL.n206 104.615
R1565 VTAIL.n206 VTAIL.n184 104.615
R1566 VTAIL.n199 VTAIL.n184 104.615
R1567 VTAIL.n199 VTAIL.n198 104.615
R1568 VTAIL.n198 VTAIL.n188 104.615
R1569 VTAIL.n191 VTAIL.n188 104.615
R1570 VTAIL.n158 VTAIL.n157 104.615
R1571 VTAIL.n157 VTAIL.n85 104.615
R1572 VTAIL.n150 VTAIL.n85 104.615
R1573 VTAIL.n150 VTAIL.n149 104.615
R1574 VTAIL.n149 VTAIL.n89 104.615
R1575 VTAIL.n142 VTAIL.n89 104.615
R1576 VTAIL.n142 VTAIL.n141 104.615
R1577 VTAIL.n141 VTAIL.n93 104.615
R1578 VTAIL.n134 VTAIL.n93 104.615
R1579 VTAIL.n134 VTAIL.n133 104.615
R1580 VTAIL.n133 VTAIL.n97 104.615
R1581 VTAIL.n101 VTAIL.n97 104.615
R1582 VTAIL.n125 VTAIL.n101 104.615
R1583 VTAIL.n125 VTAIL.n124 104.615
R1584 VTAIL.n124 VTAIL.n102 104.615
R1585 VTAIL.n117 VTAIL.n102 104.615
R1586 VTAIL.n117 VTAIL.n116 104.615
R1587 VTAIL.n116 VTAIL.n106 104.615
R1588 VTAIL.n109 VTAIL.n106 104.615
R1589 VTAIL.n272 VTAIL.t3 52.3082
R1590 VTAIL.n26 VTAIL.t1 52.3082
R1591 VTAIL.n191 VTAIL.t0 52.3082
R1592 VTAIL.n109 VTAIL.t2 52.3082
R1593 VTAIL.n327 VTAIL.n326 31.2157
R1594 VTAIL.n81 VTAIL.n80 31.2157
R1595 VTAIL.n245 VTAIL.n244 31.2157
R1596 VTAIL.n163 VTAIL.n162 31.2157
R1597 VTAIL.n163 VTAIL.n81 31.0479
R1598 VTAIL.n327 VTAIL.n245 28.1514
R1599 VTAIL.n296 VTAIL.n295 13.1884
R1600 VTAIL.n50 VTAIL.n49 13.1884
R1601 VTAIL.n214 VTAIL.n213 13.1884
R1602 VTAIL.n132 VTAIL.n131 13.1884
R1603 VTAIL.n294 VTAIL.n262 12.8005
R1604 VTAIL.n299 VTAIL.n260 12.8005
R1605 VTAIL.n48 VTAIL.n16 12.8005
R1606 VTAIL.n53 VTAIL.n14 12.8005
R1607 VTAIL.n217 VTAIL.n178 12.8005
R1608 VTAIL.n212 VTAIL.n180 12.8005
R1609 VTAIL.n135 VTAIL.n96 12.8005
R1610 VTAIL.n130 VTAIL.n98 12.8005
R1611 VTAIL.n291 VTAIL.n290 12.0247
R1612 VTAIL.n300 VTAIL.n258 12.0247
R1613 VTAIL.n45 VTAIL.n44 12.0247
R1614 VTAIL.n54 VTAIL.n12 12.0247
R1615 VTAIL.n218 VTAIL.n176 12.0247
R1616 VTAIL.n209 VTAIL.n208 12.0247
R1617 VTAIL.n136 VTAIL.n94 12.0247
R1618 VTAIL.n127 VTAIL.n126 12.0247
R1619 VTAIL.n286 VTAIL.n264 11.249
R1620 VTAIL.n304 VTAIL.n303 11.249
R1621 VTAIL.n40 VTAIL.n18 11.249
R1622 VTAIL.n58 VTAIL.n57 11.249
R1623 VTAIL.n222 VTAIL.n221 11.249
R1624 VTAIL.n205 VTAIL.n182 11.249
R1625 VTAIL.n140 VTAIL.n139 11.249
R1626 VTAIL.n123 VTAIL.n100 11.249
R1627 VTAIL.n285 VTAIL.n266 10.4732
R1628 VTAIL.n307 VTAIL.n256 10.4732
R1629 VTAIL.n39 VTAIL.n20 10.4732
R1630 VTAIL.n61 VTAIL.n10 10.4732
R1631 VTAIL.n225 VTAIL.n174 10.4732
R1632 VTAIL.n204 VTAIL.n185 10.4732
R1633 VTAIL.n143 VTAIL.n92 10.4732
R1634 VTAIL.n122 VTAIL.n103 10.4732
R1635 VTAIL.n273 VTAIL.n271 10.2747
R1636 VTAIL.n27 VTAIL.n25 10.2747
R1637 VTAIL.n192 VTAIL.n190 10.2747
R1638 VTAIL.n110 VTAIL.n108 10.2747
R1639 VTAIL.n282 VTAIL.n281 9.69747
R1640 VTAIL.n308 VTAIL.n254 9.69747
R1641 VTAIL.n36 VTAIL.n35 9.69747
R1642 VTAIL.n62 VTAIL.n8 9.69747
R1643 VTAIL.n226 VTAIL.n172 9.69747
R1644 VTAIL.n201 VTAIL.n200 9.69747
R1645 VTAIL.n144 VTAIL.n90 9.69747
R1646 VTAIL.n119 VTAIL.n118 9.69747
R1647 VTAIL.n326 VTAIL.n325 9.45567
R1648 VTAIL.n80 VTAIL.n79 9.45567
R1649 VTAIL.n244 VTAIL.n243 9.45567
R1650 VTAIL.n162 VTAIL.n161 9.45567
R1651 VTAIL.n319 VTAIL.n318 9.3005
R1652 VTAIL.n248 VTAIL.n247 9.3005
R1653 VTAIL.n325 VTAIL.n324 9.3005
R1654 VTAIL.n252 VTAIL.n251 9.3005
R1655 VTAIL.n311 VTAIL.n310 9.3005
R1656 VTAIL.n309 VTAIL.n308 9.3005
R1657 VTAIL.n256 VTAIL.n255 9.3005
R1658 VTAIL.n303 VTAIL.n302 9.3005
R1659 VTAIL.n301 VTAIL.n300 9.3005
R1660 VTAIL.n260 VTAIL.n259 9.3005
R1661 VTAIL.n275 VTAIL.n274 9.3005
R1662 VTAIL.n277 VTAIL.n276 9.3005
R1663 VTAIL.n268 VTAIL.n267 9.3005
R1664 VTAIL.n283 VTAIL.n282 9.3005
R1665 VTAIL.n285 VTAIL.n284 9.3005
R1666 VTAIL.n264 VTAIL.n263 9.3005
R1667 VTAIL.n292 VTAIL.n291 9.3005
R1668 VTAIL.n294 VTAIL.n293 9.3005
R1669 VTAIL.n317 VTAIL.n316 9.3005
R1670 VTAIL.n73 VTAIL.n72 9.3005
R1671 VTAIL.n2 VTAIL.n1 9.3005
R1672 VTAIL.n79 VTAIL.n78 9.3005
R1673 VTAIL.n6 VTAIL.n5 9.3005
R1674 VTAIL.n65 VTAIL.n64 9.3005
R1675 VTAIL.n63 VTAIL.n62 9.3005
R1676 VTAIL.n10 VTAIL.n9 9.3005
R1677 VTAIL.n57 VTAIL.n56 9.3005
R1678 VTAIL.n55 VTAIL.n54 9.3005
R1679 VTAIL.n14 VTAIL.n13 9.3005
R1680 VTAIL.n29 VTAIL.n28 9.3005
R1681 VTAIL.n31 VTAIL.n30 9.3005
R1682 VTAIL.n22 VTAIL.n21 9.3005
R1683 VTAIL.n37 VTAIL.n36 9.3005
R1684 VTAIL.n39 VTAIL.n38 9.3005
R1685 VTAIL.n18 VTAIL.n17 9.3005
R1686 VTAIL.n46 VTAIL.n45 9.3005
R1687 VTAIL.n48 VTAIL.n47 9.3005
R1688 VTAIL.n71 VTAIL.n70 9.3005
R1689 VTAIL.n166 VTAIL.n165 9.3005
R1690 VTAIL.n237 VTAIL.n236 9.3005
R1691 VTAIL.n235 VTAIL.n234 9.3005
R1692 VTAIL.n170 VTAIL.n169 9.3005
R1693 VTAIL.n229 VTAIL.n228 9.3005
R1694 VTAIL.n227 VTAIL.n226 9.3005
R1695 VTAIL.n174 VTAIL.n173 9.3005
R1696 VTAIL.n221 VTAIL.n220 9.3005
R1697 VTAIL.n219 VTAIL.n218 9.3005
R1698 VTAIL.n178 VTAIL.n177 9.3005
R1699 VTAIL.n212 VTAIL.n211 9.3005
R1700 VTAIL.n210 VTAIL.n209 9.3005
R1701 VTAIL.n182 VTAIL.n181 9.3005
R1702 VTAIL.n204 VTAIL.n203 9.3005
R1703 VTAIL.n202 VTAIL.n201 9.3005
R1704 VTAIL.n187 VTAIL.n186 9.3005
R1705 VTAIL.n196 VTAIL.n195 9.3005
R1706 VTAIL.n194 VTAIL.n193 9.3005
R1707 VTAIL.n243 VTAIL.n242 9.3005
R1708 VTAIL.n112 VTAIL.n111 9.3005
R1709 VTAIL.n114 VTAIL.n113 9.3005
R1710 VTAIL.n105 VTAIL.n104 9.3005
R1711 VTAIL.n120 VTAIL.n119 9.3005
R1712 VTAIL.n122 VTAIL.n121 9.3005
R1713 VTAIL.n100 VTAIL.n99 9.3005
R1714 VTAIL.n128 VTAIL.n127 9.3005
R1715 VTAIL.n130 VTAIL.n129 9.3005
R1716 VTAIL.n84 VTAIL.n83 9.3005
R1717 VTAIL.n161 VTAIL.n160 9.3005
R1718 VTAIL.n155 VTAIL.n154 9.3005
R1719 VTAIL.n153 VTAIL.n152 9.3005
R1720 VTAIL.n88 VTAIL.n87 9.3005
R1721 VTAIL.n147 VTAIL.n146 9.3005
R1722 VTAIL.n145 VTAIL.n144 9.3005
R1723 VTAIL.n92 VTAIL.n91 9.3005
R1724 VTAIL.n139 VTAIL.n138 9.3005
R1725 VTAIL.n137 VTAIL.n136 9.3005
R1726 VTAIL.n96 VTAIL.n95 9.3005
R1727 VTAIL.n278 VTAIL.n268 8.92171
R1728 VTAIL.n312 VTAIL.n311 8.92171
R1729 VTAIL.n326 VTAIL.n246 8.92171
R1730 VTAIL.n32 VTAIL.n22 8.92171
R1731 VTAIL.n66 VTAIL.n65 8.92171
R1732 VTAIL.n80 VTAIL.n0 8.92171
R1733 VTAIL.n244 VTAIL.n164 8.92171
R1734 VTAIL.n230 VTAIL.n229 8.92171
R1735 VTAIL.n197 VTAIL.n187 8.92171
R1736 VTAIL.n162 VTAIL.n82 8.92171
R1737 VTAIL.n148 VTAIL.n147 8.92171
R1738 VTAIL.n115 VTAIL.n105 8.92171
R1739 VTAIL.n277 VTAIL.n270 8.14595
R1740 VTAIL.n315 VTAIL.n252 8.14595
R1741 VTAIL.n324 VTAIL.n323 8.14595
R1742 VTAIL.n31 VTAIL.n24 8.14595
R1743 VTAIL.n69 VTAIL.n6 8.14595
R1744 VTAIL.n78 VTAIL.n77 8.14595
R1745 VTAIL.n242 VTAIL.n241 8.14595
R1746 VTAIL.n233 VTAIL.n170 8.14595
R1747 VTAIL.n196 VTAIL.n189 8.14595
R1748 VTAIL.n160 VTAIL.n159 8.14595
R1749 VTAIL.n151 VTAIL.n88 8.14595
R1750 VTAIL.n114 VTAIL.n107 8.14595
R1751 VTAIL.n274 VTAIL.n273 7.3702
R1752 VTAIL.n316 VTAIL.n250 7.3702
R1753 VTAIL.n320 VTAIL.n248 7.3702
R1754 VTAIL.n28 VTAIL.n27 7.3702
R1755 VTAIL.n70 VTAIL.n4 7.3702
R1756 VTAIL.n74 VTAIL.n2 7.3702
R1757 VTAIL.n238 VTAIL.n166 7.3702
R1758 VTAIL.n234 VTAIL.n168 7.3702
R1759 VTAIL.n193 VTAIL.n192 7.3702
R1760 VTAIL.n156 VTAIL.n84 7.3702
R1761 VTAIL.n152 VTAIL.n86 7.3702
R1762 VTAIL.n111 VTAIL.n110 7.3702
R1763 VTAIL.n319 VTAIL.n250 6.59444
R1764 VTAIL.n320 VTAIL.n319 6.59444
R1765 VTAIL.n73 VTAIL.n4 6.59444
R1766 VTAIL.n74 VTAIL.n73 6.59444
R1767 VTAIL.n238 VTAIL.n237 6.59444
R1768 VTAIL.n237 VTAIL.n168 6.59444
R1769 VTAIL.n156 VTAIL.n155 6.59444
R1770 VTAIL.n155 VTAIL.n86 6.59444
R1771 VTAIL.n274 VTAIL.n270 5.81868
R1772 VTAIL.n316 VTAIL.n315 5.81868
R1773 VTAIL.n323 VTAIL.n248 5.81868
R1774 VTAIL.n28 VTAIL.n24 5.81868
R1775 VTAIL.n70 VTAIL.n69 5.81868
R1776 VTAIL.n77 VTAIL.n2 5.81868
R1777 VTAIL.n241 VTAIL.n166 5.81868
R1778 VTAIL.n234 VTAIL.n233 5.81868
R1779 VTAIL.n193 VTAIL.n189 5.81868
R1780 VTAIL.n159 VTAIL.n84 5.81868
R1781 VTAIL.n152 VTAIL.n151 5.81868
R1782 VTAIL.n111 VTAIL.n107 5.81868
R1783 VTAIL.n278 VTAIL.n277 5.04292
R1784 VTAIL.n312 VTAIL.n252 5.04292
R1785 VTAIL.n324 VTAIL.n246 5.04292
R1786 VTAIL.n32 VTAIL.n31 5.04292
R1787 VTAIL.n66 VTAIL.n6 5.04292
R1788 VTAIL.n78 VTAIL.n0 5.04292
R1789 VTAIL.n242 VTAIL.n164 5.04292
R1790 VTAIL.n230 VTAIL.n170 5.04292
R1791 VTAIL.n197 VTAIL.n196 5.04292
R1792 VTAIL.n160 VTAIL.n82 5.04292
R1793 VTAIL.n148 VTAIL.n88 5.04292
R1794 VTAIL.n115 VTAIL.n114 5.04292
R1795 VTAIL.n281 VTAIL.n268 4.26717
R1796 VTAIL.n311 VTAIL.n254 4.26717
R1797 VTAIL.n35 VTAIL.n22 4.26717
R1798 VTAIL.n65 VTAIL.n8 4.26717
R1799 VTAIL.n229 VTAIL.n172 4.26717
R1800 VTAIL.n200 VTAIL.n187 4.26717
R1801 VTAIL.n147 VTAIL.n90 4.26717
R1802 VTAIL.n118 VTAIL.n105 4.26717
R1803 VTAIL.n282 VTAIL.n266 3.49141
R1804 VTAIL.n308 VTAIL.n307 3.49141
R1805 VTAIL.n36 VTAIL.n20 3.49141
R1806 VTAIL.n62 VTAIL.n61 3.49141
R1807 VTAIL.n226 VTAIL.n225 3.49141
R1808 VTAIL.n201 VTAIL.n185 3.49141
R1809 VTAIL.n144 VTAIL.n143 3.49141
R1810 VTAIL.n119 VTAIL.n103 3.49141
R1811 VTAIL.n275 VTAIL.n271 2.84303
R1812 VTAIL.n29 VTAIL.n25 2.84303
R1813 VTAIL.n194 VTAIL.n190 2.84303
R1814 VTAIL.n112 VTAIL.n108 2.84303
R1815 VTAIL.n286 VTAIL.n285 2.71565
R1816 VTAIL.n304 VTAIL.n256 2.71565
R1817 VTAIL.n40 VTAIL.n39 2.71565
R1818 VTAIL.n58 VTAIL.n10 2.71565
R1819 VTAIL.n222 VTAIL.n174 2.71565
R1820 VTAIL.n205 VTAIL.n204 2.71565
R1821 VTAIL.n140 VTAIL.n92 2.71565
R1822 VTAIL.n123 VTAIL.n122 2.71565
R1823 VTAIL.n290 VTAIL.n264 1.93989
R1824 VTAIL.n303 VTAIL.n258 1.93989
R1825 VTAIL.n44 VTAIL.n18 1.93989
R1826 VTAIL.n57 VTAIL.n12 1.93989
R1827 VTAIL.n221 VTAIL.n176 1.93989
R1828 VTAIL.n208 VTAIL.n182 1.93989
R1829 VTAIL.n139 VTAIL.n94 1.93989
R1830 VTAIL.n126 VTAIL.n100 1.93989
R1831 VTAIL.n245 VTAIL.n163 1.9186
R1832 VTAIL VTAIL.n81 1.25266
R1833 VTAIL.n291 VTAIL.n262 1.16414
R1834 VTAIL.n300 VTAIL.n299 1.16414
R1835 VTAIL.n45 VTAIL.n16 1.16414
R1836 VTAIL.n54 VTAIL.n53 1.16414
R1837 VTAIL.n218 VTAIL.n217 1.16414
R1838 VTAIL.n209 VTAIL.n180 1.16414
R1839 VTAIL.n136 VTAIL.n135 1.16414
R1840 VTAIL.n127 VTAIL.n98 1.16414
R1841 VTAIL VTAIL.n327 0.666448
R1842 VTAIL.n295 VTAIL.n294 0.388379
R1843 VTAIL.n296 VTAIL.n260 0.388379
R1844 VTAIL.n49 VTAIL.n48 0.388379
R1845 VTAIL.n50 VTAIL.n14 0.388379
R1846 VTAIL.n214 VTAIL.n178 0.388379
R1847 VTAIL.n213 VTAIL.n212 0.388379
R1848 VTAIL.n132 VTAIL.n96 0.388379
R1849 VTAIL.n131 VTAIL.n130 0.388379
R1850 VTAIL.n276 VTAIL.n275 0.155672
R1851 VTAIL.n276 VTAIL.n267 0.155672
R1852 VTAIL.n283 VTAIL.n267 0.155672
R1853 VTAIL.n284 VTAIL.n283 0.155672
R1854 VTAIL.n284 VTAIL.n263 0.155672
R1855 VTAIL.n292 VTAIL.n263 0.155672
R1856 VTAIL.n293 VTAIL.n292 0.155672
R1857 VTAIL.n293 VTAIL.n259 0.155672
R1858 VTAIL.n301 VTAIL.n259 0.155672
R1859 VTAIL.n302 VTAIL.n301 0.155672
R1860 VTAIL.n302 VTAIL.n255 0.155672
R1861 VTAIL.n309 VTAIL.n255 0.155672
R1862 VTAIL.n310 VTAIL.n309 0.155672
R1863 VTAIL.n310 VTAIL.n251 0.155672
R1864 VTAIL.n317 VTAIL.n251 0.155672
R1865 VTAIL.n318 VTAIL.n317 0.155672
R1866 VTAIL.n318 VTAIL.n247 0.155672
R1867 VTAIL.n325 VTAIL.n247 0.155672
R1868 VTAIL.n30 VTAIL.n29 0.155672
R1869 VTAIL.n30 VTAIL.n21 0.155672
R1870 VTAIL.n37 VTAIL.n21 0.155672
R1871 VTAIL.n38 VTAIL.n37 0.155672
R1872 VTAIL.n38 VTAIL.n17 0.155672
R1873 VTAIL.n46 VTAIL.n17 0.155672
R1874 VTAIL.n47 VTAIL.n46 0.155672
R1875 VTAIL.n47 VTAIL.n13 0.155672
R1876 VTAIL.n55 VTAIL.n13 0.155672
R1877 VTAIL.n56 VTAIL.n55 0.155672
R1878 VTAIL.n56 VTAIL.n9 0.155672
R1879 VTAIL.n63 VTAIL.n9 0.155672
R1880 VTAIL.n64 VTAIL.n63 0.155672
R1881 VTAIL.n64 VTAIL.n5 0.155672
R1882 VTAIL.n71 VTAIL.n5 0.155672
R1883 VTAIL.n72 VTAIL.n71 0.155672
R1884 VTAIL.n72 VTAIL.n1 0.155672
R1885 VTAIL.n79 VTAIL.n1 0.155672
R1886 VTAIL.n243 VTAIL.n165 0.155672
R1887 VTAIL.n236 VTAIL.n165 0.155672
R1888 VTAIL.n236 VTAIL.n235 0.155672
R1889 VTAIL.n235 VTAIL.n169 0.155672
R1890 VTAIL.n228 VTAIL.n169 0.155672
R1891 VTAIL.n228 VTAIL.n227 0.155672
R1892 VTAIL.n227 VTAIL.n173 0.155672
R1893 VTAIL.n220 VTAIL.n173 0.155672
R1894 VTAIL.n220 VTAIL.n219 0.155672
R1895 VTAIL.n219 VTAIL.n177 0.155672
R1896 VTAIL.n211 VTAIL.n177 0.155672
R1897 VTAIL.n211 VTAIL.n210 0.155672
R1898 VTAIL.n210 VTAIL.n181 0.155672
R1899 VTAIL.n203 VTAIL.n181 0.155672
R1900 VTAIL.n203 VTAIL.n202 0.155672
R1901 VTAIL.n202 VTAIL.n186 0.155672
R1902 VTAIL.n195 VTAIL.n186 0.155672
R1903 VTAIL.n195 VTAIL.n194 0.155672
R1904 VTAIL.n161 VTAIL.n83 0.155672
R1905 VTAIL.n154 VTAIL.n83 0.155672
R1906 VTAIL.n154 VTAIL.n153 0.155672
R1907 VTAIL.n153 VTAIL.n87 0.155672
R1908 VTAIL.n146 VTAIL.n87 0.155672
R1909 VTAIL.n146 VTAIL.n145 0.155672
R1910 VTAIL.n145 VTAIL.n91 0.155672
R1911 VTAIL.n138 VTAIL.n91 0.155672
R1912 VTAIL.n138 VTAIL.n137 0.155672
R1913 VTAIL.n137 VTAIL.n95 0.155672
R1914 VTAIL.n129 VTAIL.n95 0.155672
R1915 VTAIL.n129 VTAIL.n128 0.155672
R1916 VTAIL.n128 VTAIL.n99 0.155672
R1917 VTAIL.n121 VTAIL.n99 0.155672
R1918 VTAIL.n121 VTAIL.n120 0.155672
R1919 VTAIL.n120 VTAIL.n104 0.155672
R1920 VTAIL.n113 VTAIL.n104 0.155672
R1921 VTAIL.n113 VTAIL.n112 0.155672
R1922 VDD2.n157 VDD2.n81 289.615
R1923 VDD2.n76 VDD2.n0 289.615
R1924 VDD2.n158 VDD2.n157 185
R1925 VDD2.n156 VDD2.n155 185
R1926 VDD2.n85 VDD2.n84 185
R1927 VDD2.n150 VDD2.n149 185
R1928 VDD2.n148 VDD2.n147 185
R1929 VDD2.n89 VDD2.n88 185
R1930 VDD2.n142 VDD2.n141 185
R1931 VDD2.n140 VDD2.n139 185
R1932 VDD2.n93 VDD2.n92 185
R1933 VDD2.n134 VDD2.n133 185
R1934 VDD2.n132 VDD2.n131 185
R1935 VDD2.n130 VDD2.n96 185
R1936 VDD2.n100 VDD2.n97 185
R1937 VDD2.n125 VDD2.n124 185
R1938 VDD2.n123 VDD2.n122 185
R1939 VDD2.n102 VDD2.n101 185
R1940 VDD2.n117 VDD2.n116 185
R1941 VDD2.n115 VDD2.n114 185
R1942 VDD2.n106 VDD2.n105 185
R1943 VDD2.n109 VDD2.n108 185
R1944 VDD2.n27 VDD2.n26 185
R1945 VDD2.n24 VDD2.n23 185
R1946 VDD2.n33 VDD2.n32 185
R1947 VDD2.n35 VDD2.n34 185
R1948 VDD2.n20 VDD2.n19 185
R1949 VDD2.n41 VDD2.n40 185
R1950 VDD2.n44 VDD2.n43 185
R1951 VDD2.n42 VDD2.n16 185
R1952 VDD2.n49 VDD2.n15 185
R1953 VDD2.n51 VDD2.n50 185
R1954 VDD2.n53 VDD2.n52 185
R1955 VDD2.n12 VDD2.n11 185
R1956 VDD2.n59 VDD2.n58 185
R1957 VDD2.n61 VDD2.n60 185
R1958 VDD2.n8 VDD2.n7 185
R1959 VDD2.n67 VDD2.n66 185
R1960 VDD2.n69 VDD2.n68 185
R1961 VDD2.n4 VDD2.n3 185
R1962 VDD2.n75 VDD2.n74 185
R1963 VDD2.n77 VDD2.n76 185
R1964 VDD2.t0 VDD2.n107 149.524
R1965 VDD2.t1 VDD2.n25 149.524
R1966 VDD2.n157 VDD2.n156 104.615
R1967 VDD2.n156 VDD2.n84 104.615
R1968 VDD2.n149 VDD2.n84 104.615
R1969 VDD2.n149 VDD2.n148 104.615
R1970 VDD2.n148 VDD2.n88 104.615
R1971 VDD2.n141 VDD2.n88 104.615
R1972 VDD2.n141 VDD2.n140 104.615
R1973 VDD2.n140 VDD2.n92 104.615
R1974 VDD2.n133 VDD2.n92 104.615
R1975 VDD2.n133 VDD2.n132 104.615
R1976 VDD2.n132 VDD2.n96 104.615
R1977 VDD2.n100 VDD2.n96 104.615
R1978 VDD2.n124 VDD2.n100 104.615
R1979 VDD2.n124 VDD2.n123 104.615
R1980 VDD2.n123 VDD2.n101 104.615
R1981 VDD2.n116 VDD2.n101 104.615
R1982 VDD2.n116 VDD2.n115 104.615
R1983 VDD2.n115 VDD2.n105 104.615
R1984 VDD2.n108 VDD2.n105 104.615
R1985 VDD2.n26 VDD2.n23 104.615
R1986 VDD2.n33 VDD2.n23 104.615
R1987 VDD2.n34 VDD2.n33 104.615
R1988 VDD2.n34 VDD2.n19 104.615
R1989 VDD2.n41 VDD2.n19 104.615
R1990 VDD2.n43 VDD2.n41 104.615
R1991 VDD2.n43 VDD2.n42 104.615
R1992 VDD2.n42 VDD2.n15 104.615
R1993 VDD2.n51 VDD2.n15 104.615
R1994 VDD2.n52 VDD2.n51 104.615
R1995 VDD2.n52 VDD2.n11 104.615
R1996 VDD2.n59 VDD2.n11 104.615
R1997 VDD2.n60 VDD2.n59 104.615
R1998 VDD2.n60 VDD2.n7 104.615
R1999 VDD2.n67 VDD2.n7 104.615
R2000 VDD2.n68 VDD2.n67 104.615
R2001 VDD2.n68 VDD2.n3 104.615
R2002 VDD2.n75 VDD2.n3 104.615
R2003 VDD2.n76 VDD2.n75 104.615
R2004 VDD2.n162 VDD2.n80 90.2349
R2005 VDD2.n108 VDD2.t0 52.3082
R2006 VDD2.n26 VDD2.t1 52.3082
R2007 VDD2.n162 VDD2.n161 47.8944
R2008 VDD2.n131 VDD2.n130 13.1884
R2009 VDD2.n50 VDD2.n49 13.1884
R2010 VDD2.n134 VDD2.n95 12.8005
R2011 VDD2.n129 VDD2.n97 12.8005
R2012 VDD2.n48 VDD2.n16 12.8005
R2013 VDD2.n53 VDD2.n14 12.8005
R2014 VDD2.n135 VDD2.n93 12.0247
R2015 VDD2.n126 VDD2.n125 12.0247
R2016 VDD2.n45 VDD2.n44 12.0247
R2017 VDD2.n54 VDD2.n12 12.0247
R2018 VDD2.n139 VDD2.n138 11.249
R2019 VDD2.n122 VDD2.n99 11.249
R2020 VDD2.n40 VDD2.n18 11.249
R2021 VDD2.n58 VDD2.n57 11.249
R2022 VDD2.n142 VDD2.n91 10.4732
R2023 VDD2.n121 VDD2.n102 10.4732
R2024 VDD2.n39 VDD2.n20 10.4732
R2025 VDD2.n61 VDD2.n10 10.4732
R2026 VDD2.n109 VDD2.n107 10.2747
R2027 VDD2.n27 VDD2.n25 10.2747
R2028 VDD2.n143 VDD2.n89 9.69747
R2029 VDD2.n118 VDD2.n117 9.69747
R2030 VDD2.n36 VDD2.n35 9.69747
R2031 VDD2.n62 VDD2.n8 9.69747
R2032 VDD2.n161 VDD2.n160 9.45567
R2033 VDD2.n80 VDD2.n79 9.45567
R2034 VDD2.n83 VDD2.n82 9.3005
R2035 VDD2.n154 VDD2.n153 9.3005
R2036 VDD2.n152 VDD2.n151 9.3005
R2037 VDD2.n87 VDD2.n86 9.3005
R2038 VDD2.n146 VDD2.n145 9.3005
R2039 VDD2.n144 VDD2.n143 9.3005
R2040 VDD2.n91 VDD2.n90 9.3005
R2041 VDD2.n138 VDD2.n137 9.3005
R2042 VDD2.n136 VDD2.n135 9.3005
R2043 VDD2.n95 VDD2.n94 9.3005
R2044 VDD2.n129 VDD2.n128 9.3005
R2045 VDD2.n127 VDD2.n126 9.3005
R2046 VDD2.n99 VDD2.n98 9.3005
R2047 VDD2.n121 VDD2.n120 9.3005
R2048 VDD2.n119 VDD2.n118 9.3005
R2049 VDD2.n104 VDD2.n103 9.3005
R2050 VDD2.n113 VDD2.n112 9.3005
R2051 VDD2.n111 VDD2.n110 9.3005
R2052 VDD2.n160 VDD2.n159 9.3005
R2053 VDD2.n73 VDD2.n72 9.3005
R2054 VDD2.n2 VDD2.n1 9.3005
R2055 VDD2.n79 VDD2.n78 9.3005
R2056 VDD2.n6 VDD2.n5 9.3005
R2057 VDD2.n65 VDD2.n64 9.3005
R2058 VDD2.n63 VDD2.n62 9.3005
R2059 VDD2.n10 VDD2.n9 9.3005
R2060 VDD2.n57 VDD2.n56 9.3005
R2061 VDD2.n55 VDD2.n54 9.3005
R2062 VDD2.n14 VDD2.n13 9.3005
R2063 VDD2.n29 VDD2.n28 9.3005
R2064 VDD2.n31 VDD2.n30 9.3005
R2065 VDD2.n22 VDD2.n21 9.3005
R2066 VDD2.n37 VDD2.n36 9.3005
R2067 VDD2.n39 VDD2.n38 9.3005
R2068 VDD2.n18 VDD2.n17 9.3005
R2069 VDD2.n46 VDD2.n45 9.3005
R2070 VDD2.n48 VDD2.n47 9.3005
R2071 VDD2.n71 VDD2.n70 9.3005
R2072 VDD2.n161 VDD2.n81 8.92171
R2073 VDD2.n147 VDD2.n146 8.92171
R2074 VDD2.n114 VDD2.n104 8.92171
R2075 VDD2.n32 VDD2.n22 8.92171
R2076 VDD2.n66 VDD2.n65 8.92171
R2077 VDD2.n80 VDD2.n0 8.92171
R2078 VDD2.n159 VDD2.n158 8.14595
R2079 VDD2.n150 VDD2.n87 8.14595
R2080 VDD2.n113 VDD2.n106 8.14595
R2081 VDD2.n31 VDD2.n24 8.14595
R2082 VDD2.n69 VDD2.n6 8.14595
R2083 VDD2.n78 VDD2.n77 8.14595
R2084 VDD2.n155 VDD2.n83 7.3702
R2085 VDD2.n151 VDD2.n85 7.3702
R2086 VDD2.n110 VDD2.n109 7.3702
R2087 VDD2.n28 VDD2.n27 7.3702
R2088 VDD2.n70 VDD2.n4 7.3702
R2089 VDD2.n74 VDD2.n2 7.3702
R2090 VDD2.n155 VDD2.n154 6.59444
R2091 VDD2.n154 VDD2.n85 6.59444
R2092 VDD2.n73 VDD2.n4 6.59444
R2093 VDD2.n74 VDD2.n73 6.59444
R2094 VDD2.n158 VDD2.n83 5.81868
R2095 VDD2.n151 VDD2.n150 5.81868
R2096 VDD2.n110 VDD2.n106 5.81868
R2097 VDD2.n28 VDD2.n24 5.81868
R2098 VDD2.n70 VDD2.n69 5.81868
R2099 VDD2.n77 VDD2.n2 5.81868
R2100 VDD2.n159 VDD2.n81 5.04292
R2101 VDD2.n147 VDD2.n87 5.04292
R2102 VDD2.n114 VDD2.n113 5.04292
R2103 VDD2.n32 VDD2.n31 5.04292
R2104 VDD2.n66 VDD2.n6 5.04292
R2105 VDD2.n78 VDD2.n0 5.04292
R2106 VDD2.n146 VDD2.n89 4.26717
R2107 VDD2.n117 VDD2.n104 4.26717
R2108 VDD2.n35 VDD2.n22 4.26717
R2109 VDD2.n65 VDD2.n8 4.26717
R2110 VDD2.n143 VDD2.n142 3.49141
R2111 VDD2.n118 VDD2.n102 3.49141
R2112 VDD2.n36 VDD2.n20 3.49141
R2113 VDD2.n62 VDD2.n61 3.49141
R2114 VDD2.n29 VDD2.n25 2.84303
R2115 VDD2.n111 VDD2.n107 2.84303
R2116 VDD2.n139 VDD2.n91 2.71565
R2117 VDD2.n122 VDD2.n121 2.71565
R2118 VDD2.n40 VDD2.n39 2.71565
R2119 VDD2.n58 VDD2.n10 2.71565
R2120 VDD2.n138 VDD2.n93 1.93989
R2121 VDD2.n125 VDD2.n99 1.93989
R2122 VDD2.n44 VDD2.n18 1.93989
R2123 VDD2.n57 VDD2.n12 1.93989
R2124 VDD2.n135 VDD2.n134 1.16414
R2125 VDD2.n126 VDD2.n97 1.16414
R2126 VDD2.n45 VDD2.n16 1.16414
R2127 VDD2.n54 VDD2.n53 1.16414
R2128 VDD2 VDD2.n162 0.782828
R2129 VDD2.n131 VDD2.n95 0.388379
R2130 VDD2.n130 VDD2.n129 0.388379
R2131 VDD2.n49 VDD2.n48 0.388379
R2132 VDD2.n50 VDD2.n14 0.388379
R2133 VDD2.n160 VDD2.n82 0.155672
R2134 VDD2.n153 VDD2.n82 0.155672
R2135 VDD2.n153 VDD2.n152 0.155672
R2136 VDD2.n152 VDD2.n86 0.155672
R2137 VDD2.n145 VDD2.n86 0.155672
R2138 VDD2.n145 VDD2.n144 0.155672
R2139 VDD2.n144 VDD2.n90 0.155672
R2140 VDD2.n137 VDD2.n90 0.155672
R2141 VDD2.n137 VDD2.n136 0.155672
R2142 VDD2.n136 VDD2.n94 0.155672
R2143 VDD2.n128 VDD2.n94 0.155672
R2144 VDD2.n128 VDD2.n127 0.155672
R2145 VDD2.n127 VDD2.n98 0.155672
R2146 VDD2.n120 VDD2.n98 0.155672
R2147 VDD2.n120 VDD2.n119 0.155672
R2148 VDD2.n119 VDD2.n103 0.155672
R2149 VDD2.n112 VDD2.n103 0.155672
R2150 VDD2.n112 VDD2.n111 0.155672
R2151 VDD2.n30 VDD2.n29 0.155672
R2152 VDD2.n30 VDD2.n21 0.155672
R2153 VDD2.n37 VDD2.n21 0.155672
R2154 VDD2.n38 VDD2.n37 0.155672
R2155 VDD2.n38 VDD2.n17 0.155672
R2156 VDD2.n46 VDD2.n17 0.155672
R2157 VDD2.n47 VDD2.n46 0.155672
R2158 VDD2.n47 VDD2.n13 0.155672
R2159 VDD2.n55 VDD2.n13 0.155672
R2160 VDD2.n56 VDD2.n55 0.155672
R2161 VDD2.n56 VDD2.n9 0.155672
R2162 VDD2.n63 VDD2.n9 0.155672
R2163 VDD2.n64 VDD2.n63 0.155672
R2164 VDD2.n64 VDD2.n5 0.155672
R2165 VDD2.n71 VDD2.n5 0.155672
R2166 VDD2.n72 VDD2.n71 0.155672
R2167 VDD2.n72 VDD2.n1 0.155672
R2168 VDD2.n79 VDD2.n1 0.155672
R2169 VP.n0 VP.t1 208.037
R2170 VP.n0 VP.t0 160.006
R2171 VP VP.n0 0.431811
R2172 VDD1.n76 VDD1.n0 289.615
R2173 VDD1.n157 VDD1.n81 289.615
R2174 VDD1.n77 VDD1.n76 185
R2175 VDD1.n75 VDD1.n74 185
R2176 VDD1.n4 VDD1.n3 185
R2177 VDD1.n69 VDD1.n68 185
R2178 VDD1.n67 VDD1.n66 185
R2179 VDD1.n8 VDD1.n7 185
R2180 VDD1.n61 VDD1.n60 185
R2181 VDD1.n59 VDD1.n58 185
R2182 VDD1.n12 VDD1.n11 185
R2183 VDD1.n53 VDD1.n52 185
R2184 VDD1.n51 VDD1.n50 185
R2185 VDD1.n49 VDD1.n15 185
R2186 VDD1.n19 VDD1.n16 185
R2187 VDD1.n44 VDD1.n43 185
R2188 VDD1.n42 VDD1.n41 185
R2189 VDD1.n21 VDD1.n20 185
R2190 VDD1.n36 VDD1.n35 185
R2191 VDD1.n34 VDD1.n33 185
R2192 VDD1.n25 VDD1.n24 185
R2193 VDD1.n28 VDD1.n27 185
R2194 VDD1.n108 VDD1.n107 185
R2195 VDD1.n105 VDD1.n104 185
R2196 VDD1.n114 VDD1.n113 185
R2197 VDD1.n116 VDD1.n115 185
R2198 VDD1.n101 VDD1.n100 185
R2199 VDD1.n122 VDD1.n121 185
R2200 VDD1.n125 VDD1.n124 185
R2201 VDD1.n123 VDD1.n97 185
R2202 VDD1.n130 VDD1.n96 185
R2203 VDD1.n132 VDD1.n131 185
R2204 VDD1.n134 VDD1.n133 185
R2205 VDD1.n93 VDD1.n92 185
R2206 VDD1.n140 VDD1.n139 185
R2207 VDD1.n142 VDD1.n141 185
R2208 VDD1.n89 VDD1.n88 185
R2209 VDD1.n148 VDD1.n147 185
R2210 VDD1.n150 VDD1.n149 185
R2211 VDD1.n85 VDD1.n84 185
R2212 VDD1.n156 VDD1.n155 185
R2213 VDD1.n158 VDD1.n157 185
R2214 VDD1.t0 VDD1.n26 149.524
R2215 VDD1.t1 VDD1.n106 149.524
R2216 VDD1.n76 VDD1.n75 104.615
R2217 VDD1.n75 VDD1.n3 104.615
R2218 VDD1.n68 VDD1.n3 104.615
R2219 VDD1.n68 VDD1.n67 104.615
R2220 VDD1.n67 VDD1.n7 104.615
R2221 VDD1.n60 VDD1.n7 104.615
R2222 VDD1.n60 VDD1.n59 104.615
R2223 VDD1.n59 VDD1.n11 104.615
R2224 VDD1.n52 VDD1.n11 104.615
R2225 VDD1.n52 VDD1.n51 104.615
R2226 VDD1.n51 VDD1.n15 104.615
R2227 VDD1.n19 VDD1.n15 104.615
R2228 VDD1.n43 VDD1.n19 104.615
R2229 VDD1.n43 VDD1.n42 104.615
R2230 VDD1.n42 VDD1.n20 104.615
R2231 VDD1.n35 VDD1.n20 104.615
R2232 VDD1.n35 VDD1.n34 104.615
R2233 VDD1.n34 VDD1.n24 104.615
R2234 VDD1.n27 VDD1.n24 104.615
R2235 VDD1.n107 VDD1.n104 104.615
R2236 VDD1.n114 VDD1.n104 104.615
R2237 VDD1.n115 VDD1.n114 104.615
R2238 VDD1.n115 VDD1.n100 104.615
R2239 VDD1.n122 VDD1.n100 104.615
R2240 VDD1.n124 VDD1.n122 104.615
R2241 VDD1.n124 VDD1.n123 104.615
R2242 VDD1.n123 VDD1.n96 104.615
R2243 VDD1.n132 VDD1.n96 104.615
R2244 VDD1.n133 VDD1.n132 104.615
R2245 VDD1.n133 VDD1.n92 104.615
R2246 VDD1.n140 VDD1.n92 104.615
R2247 VDD1.n141 VDD1.n140 104.615
R2248 VDD1.n141 VDD1.n88 104.615
R2249 VDD1.n148 VDD1.n88 104.615
R2250 VDD1.n149 VDD1.n148 104.615
R2251 VDD1.n149 VDD1.n84 104.615
R2252 VDD1.n156 VDD1.n84 104.615
R2253 VDD1.n157 VDD1.n156 104.615
R2254 VDD1 VDD1.n161 91.4839
R2255 VDD1.n27 VDD1.t0 52.3082
R2256 VDD1.n107 VDD1.t1 52.3082
R2257 VDD1 VDD1.n80 48.6768
R2258 VDD1.n50 VDD1.n49 13.1884
R2259 VDD1.n131 VDD1.n130 13.1884
R2260 VDD1.n53 VDD1.n14 12.8005
R2261 VDD1.n48 VDD1.n16 12.8005
R2262 VDD1.n129 VDD1.n97 12.8005
R2263 VDD1.n134 VDD1.n95 12.8005
R2264 VDD1.n54 VDD1.n12 12.0247
R2265 VDD1.n45 VDD1.n44 12.0247
R2266 VDD1.n126 VDD1.n125 12.0247
R2267 VDD1.n135 VDD1.n93 12.0247
R2268 VDD1.n58 VDD1.n57 11.249
R2269 VDD1.n41 VDD1.n18 11.249
R2270 VDD1.n121 VDD1.n99 11.249
R2271 VDD1.n139 VDD1.n138 11.249
R2272 VDD1.n61 VDD1.n10 10.4732
R2273 VDD1.n40 VDD1.n21 10.4732
R2274 VDD1.n120 VDD1.n101 10.4732
R2275 VDD1.n142 VDD1.n91 10.4732
R2276 VDD1.n28 VDD1.n26 10.2747
R2277 VDD1.n108 VDD1.n106 10.2747
R2278 VDD1.n62 VDD1.n8 9.69747
R2279 VDD1.n37 VDD1.n36 9.69747
R2280 VDD1.n117 VDD1.n116 9.69747
R2281 VDD1.n143 VDD1.n89 9.69747
R2282 VDD1.n80 VDD1.n79 9.45567
R2283 VDD1.n161 VDD1.n160 9.45567
R2284 VDD1.n2 VDD1.n1 9.3005
R2285 VDD1.n73 VDD1.n72 9.3005
R2286 VDD1.n71 VDD1.n70 9.3005
R2287 VDD1.n6 VDD1.n5 9.3005
R2288 VDD1.n65 VDD1.n64 9.3005
R2289 VDD1.n63 VDD1.n62 9.3005
R2290 VDD1.n10 VDD1.n9 9.3005
R2291 VDD1.n57 VDD1.n56 9.3005
R2292 VDD1.n55 VDD1.n54 9.3005
R2293 VDD1.n14 VDD1.n13 9.3005
R2294 VDD1.n48 VDD1.n47 9.3005
R2295 VDD1.n46 VDD1.n45 9.3005
R2296 VDD1.n18 VDD1.n17 9.3005
R2297 VDD1.n40 VDD1.n39 9.3005
R2298 VDD1.n38 VDD1.n37 9.3005
R2299 VDD1.n23 VDD1.n22 9.3005
R2300 VDD1.n32 VDD1.n31 9.3005
R2301 VDD1.n30 VDD1.n29 9.3005
R2302 VDD1.n79 VDD1.n78 9.3005
R2303 VDD1.n154 VDD1.n153 9.3005
R2304 VDD1.n83 VDD1.n82 9.3005
R2305 VDD1.n160 VDD1.n159 9.3005
R2306 VDD1.n87 VDD1.n86 9.3005
R2307 VDD1.n146 VDD1.n145 9.3005
R2308 VDD1.n144 VDD1.n143 9.3005
R2309 VDD1.n91 VDD1.n90 9.3005
R2310 VDD1.n138 VDD1.n137 9.3005
R2311 VDD1.n136 VDD1.n135 9.3005
R2312 VDD1.n95 VDD1.n94 9.3005
R2313 VDD1.n110 VDD1.n109 9.3005
R2314 VDD1.n112 VDD1.n111 9.3005
R2315 VDD1.n103 VDD1.n102 9.3005
R2316 VDD1.n118 VDD1.n117 9.3005
R2317 VDD1.n120 VDD1.n119 9.3005
R2318 VDD1.n99 VDD1.n98 9.3005
R2319 VDD1.n127 VDD1.n126 9.3005
R2320 VDD1.n129 VDD1.n128 9.3005
R2321 VDD1.n152 VDD1.n151 9.3005
R2322 VDD1.n80 VDD1.n0 8.92171
R2323 VDD1.n66 VDD1.n65 8.92171
R2324 VDD1.n33 VDD1.n23 8.92171
R2325 VDD1.n113 VDD1.n103 8.92171
R2326 VDD1.n147 VDD1.n146 8.92171
R2327 VDD1.n161 VDD1.n81 8.92171
R2328 VDD1.n78 VDD1.n77 8.14595
R2329 VDD1.n69 VDD1.n6 8.14595
R2330 VDD1.n32 VDD1.n25 8.14595
R2331 VDD1.n112 VDD1.n105 8.14595
R2332 VDD1.n150 VDD1.n87 8.14595
R2333 VDD1.n159 VDD1.n158 8.14595
R2334 VDD1.n74 VDD1.n2 7.3702
R2335 VDD1.n70 VDD1.n4 7.3702
R2336 VDD1.n29 VDD1.n28 7.3702
R2337 VDD1.n109 VDD1.n108 7.3702
R2338 VDD1.n151 VDD1.n85 7.3702
R2339 VDD1.n155 VDD1.n83 7.3702
R2340 VDD1.n74 VDD1.n73 6.59444
R2341 VDD1.n73 VDD1.n4 6.59444
R2342 VDD1.n154 VDD1.n85 6.59444
R2343 VDD1.n155 VDD1.n154 6.59444
R2344 VDD1.n77 VDD1.n2 5.81868
R2345 VDD1.n70 VDD1.n69 5.81868
R2346 VDD1.n29 VDD1.n25 5.81868
R2347 VDD1.n109 VDD1.n105 5.81868
R2348 VDD1.n151 VDD1.n150 5.81868
R2349 VDD1.n158 VDD1.n83 5.81868
R2350 VDD1.n78 VDD1.n0 5.04292
R2351 VDD1.n66 VDD1.n6 5.04292
R2352 VDD1.n33 VDD1.n32 5.04292
R2353 VDD1.n113 VDD1.n112 5.04292
R2354 VDD1.n147 VDD1.n87 5.04292
R2355 VDD1.n159 VDD1.n81 5.04292
R2356 VDD1.n65 VDD1.n8 4.26717
R2357 VDD1.n36 VDD1.n23 4.26717
R2358 VDD1.n116 VDD1.n103 4.26717
R2359 VDD1.n146 VDD1.n89 4.26717
R2360 VDD1.n62 VDD1.n61 3.49141
R2361 VDD1.n37 VDD1.n21 3.49141
R2362 VDD1.n117 VDD1.n101 3.49141
R2363 VDD1.n143 VDD1.n142 3.49141
R2364 VDD1.n110 VDD1.n106 2.84303
R2365 VDD1.n30 VDD1.n26 2.84303
R2366 VDD1.n58 VDD1.n10 2.71565
R2367 VDD1.n41 VDD1.n40 2.71565
R2368 VDD1.n121 VDD1.n120 2.71565
R2369 VDD1.n139 VDD1.n91 2.71565
R2370 VDD1.n57 VDD1.n12 1.93989
R2371 VDD1.n44 VDD1.n18 1.93989
R2372 VDD1.n125 VDD1.n99 1.93989
R2373 VDD1.n138 VDD1.n93 1.93989
R2374 VDD1.n54 VDD1.n53 1.16414
R2375 VDD1.n45 VDD1.n16 1.16414
R2376 VDD1.n126 VDD1.n97 1.16414
R2377 VDD1.n135 VDD1.n134 1.16414
R2378 VDD1.n50 VDD1.n14 0.388379
R2379 VDD1.n49 VDD1.n48 0.388379
R2380 VDD1.n130 VDD1.n129 0.388379
R2381 VDD1.n131 VDD1.n95 0.388379
R2382 VDD1.n79 VDD1.n1 0.155672
R2383 VDD1.n72 VDD1.n1 0.155672
R2384 VDD1.n72 VDD1.n71 0.155672
R2385 VDD1.n71 VDD1.n5 0.155672
R2386 VDD1.n64 VDD1.n5 0.155672
R2387 VDD1.n64 VDD1.n63 0.155672
R2388 VDD1.n63 VDD1.n9 0.155672
R2389 VDD1.n56 VDD1.n9 0.155672
R2390 VDD1.n56 VDD1.n55 0.155672
R2391 VDD1.n55 VDD1.n13 0.155672
R2392 VDD1.n47 VDD1.n13 0.155672
R2393 VDD1.n47 VDD1.n46 0.155672
R2394 VDD1.n46 VDD1.n17 0.155672
R2395 VDD1.n39 VDD1.n17 0.155672
R2396 VDD1.n39 VDD1.n38 0.155672
R2397 VDD1.n38 VDD1.n22 0.155672
R2398 VDD1.n31 VDD1.n22 0.155672
R2399 VDD1.n31 VDD1.n30 0.155672
R2400 VDD1.n111 VDD1.n110 0.155672
R2401 VDD1.n111 VDD1.n102 0.155672
R2402 VDD1.n118 VDD1.n102 0.155672
R2403 VDD1.n119 VDD1.n118 0.155672
R2404 VDD1.n119 VDD1.n98 0.155672
R2405 VDD1.n127 VDD1.n98 0.155672
R2406 VDD1.n128 VDD1.n127 0.155672
R2407 VDD1.n128 VDD1.n94 0.155672
R2408 VDD1.n136 VDD1.n94 0.155672
R2409 VDD1.n137 VDD1.n136 0.155672
R2410 VDD1.n137 VDD1.n90 0.155672
R2411 VDD1.n144 VDD1.n90 0.155672
R2412 VDD1.n145 VDD1.n144 0.155672
R2413 VDD1.n145 VDD1.n86 0.155672
R2414 VDD1.n152 VDD1.n86 0.155672
R2415 VDD1.n153 VDD1.n152 0.155672
R2416 VDD1.n153 VDD1.n82 0.155672
R2417 VDD1.n160 VDD1.n82 0.155672
C0 VTAIL VDD1 5.89789f
C1 VN VTAIL 3.04281f
C2 VTAIL VDD2 5.95121f
C3 VP VDD1 3.67876f
C4 VN VP 6.20173f
C5 VP VDD2 0.351333f
C6 VTAIL VP 3.0571f
C7 VN VDD1 0.148319f
C8 VDD1 VDD2 0.7271f
C9 VN VDD2 3.47853f
C10 VDD2 B 5.109983f
C11 VDD1 B 8.139919f
C12 VTAIL B 8.775948f
C13 VN B 11.78707f
C14 VP B 7.123488f
C15 VDD1.n0 B 0.030074f
C16 VDD1.n1 B 0.020323f
C17 VDD1.n2 B 0.010921f
C18 VDD1.n3 B 0.025813f
C19 VDD1.n4 B 0.011563f
C20 VDD1.n5 B 0.020323f
C21 VDD1.n6 B 0.010921f
C22 VDD1.n7 B 0.025813f
C23 VDD1.n8 B 0.011563f
C24 VDD1.n9 B 0.020323f
C25 VDD1.n10 B 0.010921f
C26 VDD1.n11 B 0.025813f
C27 VDD1.n12 B 0.011563f
C28 VDD1.n13 B 0.020323f
C29 VDD1.n14 B 0.010921f
C30 VDD1.n15 B 0.025813f
C31 VDD1.n16 B 0.011563f
C32 VDD1.n17 B 0.020323f
C33 VDD1.n18 B 0.010921f
C34 VDD1.n19 B 0.025813f
C35 VDD1.n20 B 0.025813f
C36 VDD1.n21 B 0.011563f
C37 VDD1.n22 B 0.020323f
C38 VDD1.n23 B 0.010921f
C39 VDD1.n24 B 0.025813f
C40 VDD1.n25 B 0.011563f
C41 VDD1.n26 B 0.169544f
C42 VDD1.t0 B 0.043919f
C43 VDD1.n27 B 0.01936f
C44 VDD1.n28 B 0.018248f
C45 VDD1.n29 B 0.010921f
C46 VDD1.n30 B 1.29193f
C47 VDD1.n31 B 0.020323f
C48 VDD1.n32 B 0.010921f
C49 VDD1.n33 B 0.011563f
C50 VDD1.n34 B 0.025813f
C51 VDD1.n35 B 0.025813f
C52 VDD1.n36 B 0.011563f
C53 VDD1.n37 B 0.010921f
C54 VDD1.n38 B 0.020323f
C55 VDD1.n39 B 0.020323f
C56 VDD1.n40 B 0.010921f
C57 VDD1.n41 B 0.011563f
C58 VDD1.n42 B 0.025813f
C59 VDD1.n43 B 0.025813f
C60 VDD1.n44 B 0.011563f
C61 VDD1.n45 B 0.010921f
C62 VDD1.n46 B 0.020323f
C63 VDD1.n47 B 0.020323f
C64 VDD1.n48 B 0.010921f
C65 VDD1.n49 B 0.011242f
C66 VDD1.n50 B 0.011242f
C67 VDD1.n51 B 0.025813f
C68 VDD1.n52 B 0.025813f
C69 VDD1.n53 B 0.011563f
C70 VDD1.n54 B 0.010921f
C71 VDD1.n55 B 0.020323f
C72 VDD1.n56 B 0.020323f
C73 VDD1.n57 B 0.010921f
C74 VDD1.n58 B 0.011563f
C75 VDD1.n59 B 0.025813f
C76 VDD1.n60 B 0.025813f
C77 VDD1.n61 B 0.011563f
C78 VDD1.n62 B 0.010921f
C79 VDD1.n63 B 0.020323f
C80 VDD1.n64 B 0.020323f
C81 VDD1.n65 B 0.010921f
C82 VDD1.n66 B 0.011563f
C83 VDD1.n67 B 0.025813f
C84 VDD1.n68 B 0.025813f
C85 VDD1.n69 B 0.011563f
C86 VDD1.n70 B 0.010921f
C87 VDD1.n71 B 0.020323f
C88 VDD1.n72 B 0.020323f
C89 VDD1.n73 B 0.010921f
C90 VDD1.n74 B 0.011563f
C91 VDD1.n75 B 0.025813f
C92 VDD1.n76 B 0.058547f
C93 VDD1.n77 B 0.011563f
C94 VDD1.n78 B 0.010921f
C95 VDD1.n79 B 0.045588f
C96 VDD1.n80 B 0.048474f
C97 VDD1.n81 B 0.030074f
C98 VDD1.n82 B 0.020323f
C99 VDD1.n83 B 0.010921f
C100 VDD1.n84 B 0.025813f
C101 VDD1.n85 B 0.011563f
C102 VDD1.n86 B 0.020323f
C103 VDD1.n87 B 0.010921f
C104 VDD1.n88 B 0.025813f
C105 VDD1.n89 B 0.011563f
C106 VDD1.n90 B 0.020323f
C107 VDD1.n91 B 0.010921f
C108 VDD1.n92 B 0.025813f
C109 VDD1.n93 B 0.011563f
C110 VDD1.n94 B 0.020323f
C111 VDD1.n95 B 0.010921f
C112 VDD1.n96 B 0.025813f
C113 VDD1.n97 B 0.011563f
C114 VDD1.n98 B 0.020323f
C115 VDD1.n99 B 0.010921f
C116 VDD1.n100 B 0.025813f
C117 VDD1.n101 B 0.011563f
C118 VDD1.n102 B 0.020323f
C119 VDD1.n103 B 0.010921f
C120 VDD1.n104 B 0.025813f
C121 VDD1.n105 B 0.011563f
C122 VDD1.n106 B 0.169544f
C123 VDD1.t1 B 0.043919f
C124 VDD1.n107 B 0.01936f
C125 VDD1.n108 B 0.018248f
C126 VDD1.n109 B 0.010921f
C127 VDD1.n110 B 1.29193f
C128 VDD1.n111 B 0.020323f
C129 VDD1.n112 B 0.010921f
C130 VDD1.n113 B 0.011563f
C131 VDD1.n114 B 0.025813f
C132 VDD1.n115 B 0.025813f
C133 VDD1.n116 B 0.011563f
C134 VDD1.n117 B 0.010921f
C135 VDD1.n118 B 0.020323f
C136 VDD1.n119 B 0.020323f
C137 VDD1.n120 B 0.010921f
C138 VDD1.n121 B 0.011563f
C139 VDD1.n122 B 0.025813f
C140 VDD1.n123 B 0.025813f
C141 VDD1.n124 B 0.025813f
C142 VDD1.n125 B 0.011563f
C143 VDD1.n126 B 0.010921f
C144 VDD1.n127 B 0.020323f
C145 VDD1.n128 B 0.020323f
C146 VDD1.n129 B 0.010921f
C147 VDD1.n130 B 0.011242f
C148 VDD1.n131 B 0.011242f
C149 VDD1.n132 B 0.025813f
C150 VDD1.n133 B 0.025813f
C151 VDD1.n134 B 0.011563f
C152 VDD1.n135 B 0.010921f
C153 VDD1.n136 B 0.020323f
C154 VDD1.n137 B 0.020323f
C155 VDD1.n138 B 0.010921f
C156 VDD1.n139 B 0.011563f
C157 VDD1.n140 B 0.025813f
C158 VDD1.n141 B 0.025813f
C159 VDD1.n142 B 0.011563f
C160 VDD1.n143 B 0.010921f
C161 VDD1.n144 B 0.020323f
C162 VDD1.n145 B 0.020323f
C163 VDD1.n146 B 0.010921f
C164 VDD1.n147 B 0.011563f
C165 VDD1.n148 B 0.025813f
C166 VDD1.n149 B 0.025813f
C167 VDD1.n150 B 0.011563f
C168 VDD1.n151 B 0.010921f
C169 VDD1.n152 B 0.020323f
C170 VDD1.n153 B 0.020323f
C171 VDD1.n154 B 0.010921f
C172 VDD1.n155 B 0.011563f
C173 VDD1.n156 B 0.025813f
C174 VDD1.n157 B 0.058547f
C175 VDD1.n158 B 0.011563f
C176 VDD1.n159 B 0.010921f
C177 VDD1.n160 B 0.045588f
C178 VDD1.n161 B 0.762866f
C179 VP.t0 B 3.83862f
C180 VP.t1 B 4.45067f
C181 VP.n0 B 4.62637f
C182 VDD2.n0 B 0.029996f
C183 VDD2.n1 B 0.02027f
C184 VDD2.n2 B 0.010892f
C185 VDD2.n3 B 0.025745f
C186 VDD2.n4 B 0.011533f
C187 VDD2.n5 B 0.02027f
C188 VDD2.n6 B 0.010892f
C189 VDD2.n7 B 0.025745f
C190 VDD2.n8 B 0.011533f
C191 VDD2.n9 B 0.02027f
C192 VDD2.n10 B 0.010892f
C193 VDD2.n11 B 0.025745f
C194 VDD2.n12 B 0.011533f
C195 VDD2.n13 B 0.02027f
C196 VDD2.n14 B 0.010892f
C197 VDD2.n15 B 0.025745f
C198 VDD2.n16 B 0.011533f
C199 VDD2.n17 B 0.02027f
C200 VDD2.n18 B 0.010892f
C201 VDD2.n19 B 0.025745f
C202 VDD2.n20 B 0.011533f
C203 VDD2.n21 B 0.02027f
C204 VDD2.n22 B 0.010892f
C205 VDD2.n23 B 0.025745f
C206 VDD2.n24 B 0.011533f
C207 VDD2.n25 B 0.1691f
C208 VDD2.t1 B 0.043804f
C209 VDD2.n26 B 0.019309f
C210 VDD2.n27 B 0.0182f
C211 VDD2.n28 B 0.010892f
C212 VDD2.n29 B 1.28855f
C213 VDD2.n30 B 0.02027f
C214 VDD2.n31 B 0.010892f
C215 VDD2.n32 B 0.011533f
C216 VDD2.n33 B 0.025745f
C217 VDD2.n34 B 0.025745f
C218 VDD2.n35 B 0.011533f
C219 VDD2.n36 B 0.010892f
C220 VDD2.n37 B 0.02027f
C221 VDD2.n38 B 0.02027f
C222 VDD2.n39 B 0.010892f
C223 VDD2.n40 B 0.011533f
C224 VDD2.n41 B 0.025745f
C225 VDD2.n42 B 0.025745f
C226 VDD2.n43 B 0.025745f
C227 VDD2.n44 B 0.011533f
C228 VDD2.n45 B 0.010892f
C229 VDD2.n46 B 0.02027f
C230 VDD2.n47 B 0.02027f
C231 VDD2.n48 B 0.010892f
C232 VDD2.n49 B 0.011212f
C233 VDD2.n50 B 0.011212f
C234 VDD2.n51 B 0.025745f
C235 VDD2.n52 B 0.025745f
C236 VDD2.n53 B 0.011533f
C237 VDD2.n54 B 0.010892f
C238 VDD2.n55 B 0.02027f
C239 VDD2.n56 B 0.02027f
C240 VDD2.n57 B 0.010892f
C241 VDD2.n58 B 0.011533f
C242 VDD2.n59 B 0.025745f
C243 VDD2.n60 B 0.025745f
C244 VDD2.n61 B 0.011533f
C245 VDD2.n62 B 0.010892f
C246 VDD2.n63 B 0.02027f
C247 VDD2.n64 B 0.02027f
C248 VDD2.n65 B 0.010892f
C249 VDD2.n66 B 0.011533f
C250 VDD2.n67 B 0.025745f
C251 VDD2.n68 B 0.025745f
C252 VDD2.n69 B 0.011533f
C253 VDD2.n70 B 0.010892f
C254 VDD2.n71 B 0.02027f
C255 VDD2.n72 B 0.02027f
C256 VDD2.n73 B 0.010892f
C257 VDD2.n74 B 0.011533f
C258 VDD2.n75 B 0.025745f
C259 VDD2.n76 B 0.058394f
C260 VDD2.n77 B 0.011533f
C261 VDD2.n78 B 0.010892f
C262 VDD2.n79 B 0.045468f
C263 VDD2.n80 B 0.715522f
C264 VDD2.n81 B 0.029996f
C265 VDD2.n82 B 0.02027f
C266 VDD2.n83 B 0.010892f
C267 VDD2.n84 B 0.025745f
C268 VDD2.n85 B 0.011533f
C269 VDD2.n86 B 0.02027f
C270 VDD2.n87 B 0.010892f
C271 VDD2.n88 B 0.025745f
C272 VDD2.n89 B 0.011533f
C273 VDD2.n90 B 0.02027f
C274 VDD2.n91 B 0.010892f
C275 VDD2.n92 B 0.025745f
C276 VDD2.n93 B 0.011533f
C277 VDD2.n94 B 0.02027f
C278 VDD2.n95 B 0.010892f
C279 VDD2.n96 B 0.025745f
C280 VDD2.n97 B 0.011533f
C281 VDD2.n98 B 0.02027f
C282 VDD2.n99 B 0.010892f
C283 VDD2.n100 B 0.025745f
C284 VDD2.n101 B 0.025745f
C285 VDD2.n102 B 0.011533f
C286 VDD2.n103 B 0.02027f
C287 VDD2.n104 B 0.010892f
C288 VDD2.n105 B 0.025745f
C289 VDD2.n106 B 0.011533f
C290 VDD2.n107 B 0.1691f
C291 VDD2.t0 B 0.043804f
C292 VDD2.n108 B 0.019309f
C293 VDD2.n109 B 0.0182f
C294 VDD2.n110 B 0.010892f
C295 VDD2.n111 B 1.28855f
C296 VDD2.n112 B 0.02027f
C297 VDD2.n113 B 0.010892f
C298 VDD2.n114 B 0.011533f
C299 VDD2.n115 B 0.025745f
C300 VDD2.n116 B 0.025745f
C301 VDD2.n117 B 0.011533f
C302 VDD2.n118 B 0.010892f
C303 VDD2.n119 B 0.02027f
C304 VDD2.n120 B 0.02027f
C305 VDD2.n121 B 0.010892f
C306 VDD2.n122 B 0.011533f
C307 VDD2.n123 B 0.025745f
C308 VDD2.n124 B 0.025745f
C309 VDD2.n125 B 0.011533f
C310 VDD2.n126 B 0.010892f
C311 VDD2.n127 B 0.02027f
C312 VDD2.n128 B 0.02027f
C313 VDD2.n129 B 0.010892f
C314 VDD2.n130 B 0.011212f
C315 VDD2.n131 B 0.011212f
C316 VDD2.n132 B 0.025745f
C317 VDD2.n133 B 0.025745f
C318 VDD2.n134 B 0.011533f
C319 VDD2.n135 B 0.010892f
C320 VDD2.n136 B 0.02027f
C321 VDD2.n137 B 0.02027f
C322 VDD2.n138 B 0.010892f
C323 VDD2.n139 B 0.011533f
C324 VDD2.n140 B 0.025745f
C325 VDD2.n141 B 0.025745f
C326 VDD2.n142 B 0.011533f
C327 VDD2.n143 B 0.010892f
C328 VDD2.n144 B 0.02027f
C329 VDD2.n145 B 0.02027f
C330 VDD2.n146 B 0.010892f
C331 VDD2.n147 B 0.011533f
C332 VDD2.n148 B 0.025745f
C333 VDD2.n149 B 0.025745f
C334 VDD2.n150 B 0.011533f
C335 VDD2.n151 B 0.010892f
C336 VDD2.n152 B 0.02027f
C337 VDD2.n153 B 0.02027f
C338 VDD2.n154 B 0.010892f
C339 VDD2.n155 B 0.011533f
C340 VDD2.n156 B 0.025745f
C341 VDD2.n157 B 0.058394f
C342 VDD2.n158 B 0.011533f
C343 VDD2.n159 B 0.010892f
C344 VDD2.n160 B 0.045468f
C345 VDD2.n161 B 0.046911f
C346 VDD2.n162 B 2.77881f
C347 VTAIL.n0 B 0.030117f
C348 VTAIL.n1 B 0.020352f
C349 VTAIL.n2 B 0.010936f
C350 VTAIL.n3 B 0.025849f
C351 VTAIL.n4 B 0.01158f
C352 VTAIL.n5 B 0.020352f
C353 VTAIL.n6 B 0.010936f
C354 VTAIL.n7 B 0.025849f
C355 VTAIL.n8 B 0.01158f
C356 VTAIL.n9 B 0.020352f
C357 VTAIL.n10 B 0.010936f
C358 VTAIL.n11 B 0.025849f
C359 VTAIL.n12 B 0.01158f
C360 VTAIL.n13 B 0.020352f
C361 VTAIL.n14 B 0.010936f
C362 VTAIL.n15 B 0.025849f
C363 VTAIL.n16 B 0.01158f
C364 VTAIL.n17 B 0.020352f
C365 VTAIL.n18 B 0.010936f
C366 VTAIL.n19 B 0.025849f
C367 VTAIL.n20 B 0.01158f
C368 VTAIL.n21 B 0.020352f
C369 VTAIL.n22 B 0.010936f
C370 VTAIL.n23 B 0.025849f
C371 VTAIL.n24 B 0.01158f
C372 VTAIL.n25 B 0.169785f
C373 VTAIL.t1 B 0.043981f
C374 VTAIL.n26 B 0.019387f
C375 VTAIL.n27 B 0.018274f
C376 VTAIL.n28 B 0.010936f
C377 VTAIL.n29 B 1.29376f
C378 VTAIL.n30 B 0.020352f
C379 VTAIL.n31 B 0.010936f
C380 VTAIL.n32 B 0.01158f
C381 VTAIL.n33 B 0.025849f
C382 VTAIL.n34 B 0.025849f
C383 VTAIL.n35 B 0.01158f
C384 VTAIL.n36 B 0.010936f
C385 VTAIL.n37 B 0.020352f
C386 VTAIL.n38 B 0.020352f
C387 VTAIL.n39 B 0.010936f
C388 VTAIL.n40 B 0.01158f
C389 VTAIL.n41 B 0.025849f
C390 VTAIL.n42 B 0.025849f
C391 VTAIL.n43 B 0.025849f
C392 VTAIL.n44 B 0.01158f
C393 VTAIL.n45 B 0.010936f
C394 VTAIL.n46 B 0.020352f
C395 VTAIL.n47 B 0.020352f
C396 VTAIL.n48 B 0.010936f
C397 VTAIL.n49 B 0.011258f
C398 VTAIL.n50 B 0.011258f
C399 VTAIL.n51 B 0.025849f
C400 VTAIL.n52 B 0.025849f
C401 VTAIL.n53 B 0.01158f
C402 VTAIL.n54 B 0.010936f
C403 VTAIL.n55 B 0.020352f
C404 VTAIL.n56 B 0.020352f
C405 VTAIL.n57 B 0.010936f
C406 VTAIL.n58 B 0.01158f
C407 VTAIL.n59 B 0.025849f
C408 VTAIL.n60 B 0.025849f
C409 VTAIL.n61 B 0.01158f
C410 VTAIL.n62 B 0.010936f
C411 VTAIL.n63 B 0.020352f
C412 VTAIL.n64 B 0.020352f
C413 VTAIL.n65 B 0.010936f
C414 VTAIL.n66 B 0.01158f
C415 VTAIL.n67 B 0.025849f
C416 VTAIL.n68 B 0.025849f
C417 VTAIL.n69 B 0.01158f
C418 VTAIL.n70 B 0.010936f
C419 VTAIL.n71 B 0.020352f
C420 VTAIL.n72 B 0.020352f
C421 VTAIL.n73 B 0.010936f
C422 VTAIL.n74 B 0.01158f
C423 VTAIL.n75 B 0.025849f
C424 VTAIL.n76 B 0.058631f
C425 VTAIL.n77 B 0.01158f
C426 VTAIL.n78 B 0.010936f
C427 VTAIL.n79 B 0.045653f
C428 VTAIL.n80 B 0.033037f
C429 VTAIL.n81 B 1.60025f
C430 VTAIL.n82 B 0.030117f
C431 VTAIL.n83 B 0.020352f
C432 VTAIL.n84 B 0.010936f
C433 VTAIL.n85 B 0.025849f
C434 VTAIL.n86 B 0.01158f
C435 VTAIL.n87 B 0.020352f
C436 VTAIL.n88 B 0.010936f
C437 VTAIL.n89 B 0.025849f
C438 VTAIL.n90 B 0.01158f
C439 VTAIL.n91 B 0.020352f
C440 VTAIL.n92 B 0.010936f
C441 VTAIL.n93 B 0.025849f
C442 VTAIL.n94 B 0.01158f
C443 VTAIL.n95 B 0.020352f
C444 VTAIL.n96 B 0.010936f
C445 VTAIL.n97 B 0.025849f
C446 VTAIL.n98 B 0.01158f
C447 VTAIL.n99 B 0.020352f
C448 VTAIL.n100 B 0.010936f
C449 VTAIL.n101 B 0.025849f
C450 VTAIL.n102 B 0.025849f
C451 VTAIL.n103 B 0.01158f
C452 VTAIL.n104 B 0.020352f
C453 VTAIL.n105 B 0.010936f
C454 VTAIL.n106 B 0.025849f
C455 VTAIL.n107 B 0.01158f
C456 VTAIL.n108 B 0.169785f
C457 VTAIL.t2 B 0.043981f
C458 VTAIL.n109 B 0.019387f
C459 VTAIL.n110 B 0.018274f
C460 VTAIL.n111 B 0.010936f
C461 VTAIL.n112 B 1.29376f
C462 VTAIL.n113 B 0.020352f
C463 VTAIL.n114 B 0.010936f
C464 VTAIL.n115 B 0.01158f
C465 VTAIL.n116 B 0.025849f
C466 VTAIL.n117 B 0.025849f
C467 VTAIL.n118 B 0.01158f
C468 VTAIL.n119 B 0.010936f
C469 VTAIL.n120 B 0.020352f
C470 VTAIL.n121 B 0.020352f
C471 VTAIL.n122 B 0.010936f
C472 VTAIL.n123 B 0.01158f
C473 VTAIL.n124 B 0.025849f
C474 VTAIL.n125 B 0.025849f
C475 VTAIL.n126 B 0.01158f
C476 VTAIL.n127 B 0.010936f
C477 VTAIL.n128 B 0.020352f
C478 VTAIL.n129 B 0.020352f
C479 VTAIL.n130 B 0.010936f
C480 VTAIL.n131 B 0.011258f
C481 VTAIL.n132 B 0.011258f
C482 VTAIL.n133 B 0.025849f
C483 VTAIL.n134 B 0.025849f
C484 VTAIL.n135 B 0.01158f
C485 VTAIL.n136 B 0.010936f
C486 VTAIL.n137 B 0.020352f
C487 VTAIL.n138 B 0.020352f
C488 VTAIL.n139 B 0.010936f
C489 VTAIL.n140 B 0.01158f
C490 VTAIL.n141 B 0.025849f
C491 VTAIL.n142 B 0.025849f
C492 VTAIL.n143 B 0.01158f
C493 VTAIL.n144 B 0.010936f
C494 VTAIL.n145 B 0.020352f
C495 VTAIL.n146 B 0.020352f
C496 VTAIL.n147 B 0.010936f
C497 VTAIL.n148 B 0.01158f
C498 VTAIL.n149 B 0.025849f
C499 VTAIL.n150 B 0.025849f
C500 VTAIL.n151 B 0.01158f
C501 VTAIL.n152 B 0.010936f
C502 VTAIL.n153 B 0.020352f
C503 VTAIL.n154 B 0.020352f
C504 VTAIL.n155 B 0.010936f
C505 VTAIL.n156 B 0.01158f
C506 VTAIL.n157 B 0.025849f
C507 VTAIL.n158 B 0.058631f
C508 VTAIL.n159 B 0.01158f
C509 VTAIL.n160 B 0.010936f
C510 VTAIL.n161 B 0.045653f
C511 VTAIL.n162 B 0.033037f
C512 VTAIL.n163 B 1.64392f
C513 VTAIL.n164 B 0.030117f
C514 VTAIL.n165 B 0.020352f
C515 VTAIL.n166 B 0.010936f
C516 VTAIL.n167 B 0.025849f
C517 VTAIL.n168 B 0.01158f
C518 VTAIL.n169 B 0.020352f
C519 VTAIL.n170 B 0.010936f
C520 VTAIL.n171 B 0.025849f
C521 VTAIL.n172 B 0.01158f
C522 VTAIL.n173 B 0.020352f
C523 VTAIL.n174 B 0.010936f
C524 VTAIL.n175 B 0.025849f
C525 VTAIL.n176 B 0.01158f
C526 VTAIL.n177 B 0.020352f
C527 VTAIL.n178 B 0.010936f
C528 VTAIL.n179 B 0.025849f
C529 VTAIL.n180 B 0.01158f
C530 VTAIL.n181 B 0.020352f
C531 VTAIL.n182 B 0.010936f
C532 VTAIL.n183 B 0.025849f
C533 VTAIL.n184 B 0.025849f
C534 VTAIL.n185 B 0.01158f
C535 VTAIL.n186 B 0.020352f
C536 VTAIL.n187 B 0.010936f
C537 VTAIL.n188 B 0.025849f
C538 VTAIL.n189 B 0.01158f
C539 VTAIL.n190 B 0.169785f
C540 VTAIL.t0 B 0.043981f
C541 VTAIL.n191 B 0.019387f
C542 VTAIL.n192 B 0.018274f
C543 VTAIL.n193 B 0.010936f
C544 VTAIL.n194 B 1.29376f
C545 VTAIL.n195 B 0.020352f
C546 VTAIL.n196 B 0.010936f
C547 VTAIL.n197 B 0.01158f
C548 VTAIL.n198 B 0.025849f
C549 VTAIL.n199 B 0.025849f
C550 VTAIL.n200 B 0.01158f
C551 VTAIL.n201 B 0.010936f
C552 VTAIL.n202 B 0.020352f
C553 VTAIL.n203 B 0.020352f
C554 VTAIL.n204 B 0.010936f
C555 VTAIL.n205 B 0.01158f
C556 VTAIL.n206 B 0.025849f
C557 VTAIL.n207 B 0.025849f
C558 VTAIL.n208 B 0.01158f
C559 VTAIL.n209 B 0.010936f
C560 VTAIL.n210 B 0.020352f
C561 VTAIL.n211 B 0.020352f
C562 VTAIL.n212 B 0.010936f
C563 VTAIL.n213 B 0.011258f
C564 VTAIL.n214 B 0.011258f
C565 VTAIL.n215 B 0.025849f
C566 VTAIL.n216 B 0.025849f
C567 VTAIL.n217 B 0.01158f
C568 VTAIL.n218 B 0.010936f
C569 VTAIL.n219 B 0.020352f
C570 VTAIL.n220 B 0.020352f
C571 VTAIL.n221 B 0.010936f
C572 VTAIL.n222 B 0.01158f
C573 VTAIL.n223 B 0.025849f
C574 VTAIL.n224 B 0.025849f
C575 VTAIL.n225 B 0.01158f
C576 VTAIL.n226 B 0.010936f
C577 VTAIL.n227 B 0.020352f
C578 VTAIL.n228 B 0.020352f
C579 VTAIL.n229 B 0.010936f
C580 VTAIL.n230 B 0.01158f
C581 VTAIL.n231 B 0.025849f
C582 VTAIL.n232 B 0.025849f
C583 VTAIL.n233 B 0.01158f
C584 VTAIL.n234 B 0.010936f
C585 VTAIL.n235 B 0.020352f
C586 VTAIL.n236 B 0.020352f
C587 VTAIL.n237 B 0.010936f
C588 VTAIL.n238 B 0.01158f
C589 VTAIL.n239 B 0.025849f
C590 VTAIL.n240 B 0.058631f
C591 VTAIL.n241 B 0.01158f
C592 VTAIL.n242 B 0.010936f
C593 VTAIL.n243 B 0.045653f
C594 VTAIL.n244 B 0.033037f
C595 VTAIL.n245 B 1.45397f
C596 VTAIL.n246 B 0.030117f
C597 VTAIL.n247 B 0.020352f
C598 VTAIL.n248 B 0.010936f
C599 VTAIL.n249 B 0.025849f
C600 VTAIL.n250 B 0.01158f
C601 VTAIL.n251 B 0.020352f
C602 VTAIL.n252 B 0.010936f
C603 VTAIL.n253 B 0.025849f
C604 VTAIL.n254 B 0.01158f
C605 VTAIL.n255 B 0.020352f
C606 VTAIL.n256 B 0.010936f
C607 VTAIL.n257 B 0.025849f
C608 VTAIL.n258 B 0.01158f
C609 VTAIL.n259 B 0.020352f
C610 VTAIL.n260 B 0.010936f
C611 VTAIL.n261 B 0.025849f
C612 VTAIL.n262 B 0.01158f
C613 VTAIL.n263 B 0.020352f
C614 VTAIL.n264 B 0.010936f
C615 VTAIL.n265 B 0.025849f
C616 VTAIL.n266 B 0.01158f
C617 VTAIL.n267 B 0.020352f
C618 VTAIL.n268 B 0.010936f
C619 VTAIL.n269 B 0.025849f
C620 VTAIL.n270 B 0.01158f
C621 VTAIL.n271 B 0.169785f
C622 VTAIL.t3 B 0.043981f
C623 VTAIL.n272 B 0.019387f
C624 VTAIL.n273 B 0.018274f
C625 VTAIL.n274 B 0.010936f
C626 VTAIL.n275 B 1.29376f
C627 VTAIL.n276 B 0.020352f
C628 VTAIL.n277 B 0.010936f
C629 VTAIL.n278 B 0.01158f
C630 VTAIL.n279 B 0.025849f
C631 VTAIL.n280 B 0.025849f
C632 VTAIL.n281 B 0.01158f
C633 VTAIL.n282 B 0.010936f
C634 VTAIL.n283 B 0.020352f
C635 VTAIL.n284 B 0.020352f
C636 VTAIL.n285 B 0.010936f
C637 VTAIL.n286 B 0.01158f
C638 VTAIL.n287 B 0.025849f
C639 VTAIL.n288 B 0.025849f
C640 VTAIL.n289 B 0.025849f
C641 VTAIL.n290 B 0.01158f
C642 VTAIL.n291 B 0.010936f
C643 VTAIL.n292 B 0.020352f
C644 VTAIL.n293 B 0.020352f
C645 VTAIL.n294 B 0.010936f
C646 VTAIL.n295 B 0.011258f
C647 VTAIL.n296 B 0.011258f
C648 VTAIL.n297 B 0.025849f
C649 VTAIL.n298 B 0.025849f
C650 VTAIL.n299 B 0.01158f
C651 VTAIL.n300 B 0.010936f
C652 VTAIL.n301 B 0.020352f
C653 VTAIL.n302 B 0.020352f
C654 VTAIL.n303 B 0.010936f
C655 VTAIL.n304 B 0.01158f
C656 VTAIL.n305 B 0.025849f
C657 VTAIL.n306 B 0.025849f
C658 VTAIL.n307 B 0.01158f
C659 VTAIL.n308 B 0.010936f
C660 VTAIL.n309 B 0.020352f
C661 VTAIL.n310 B 0.020352f
C662 VTAIL.n311 B 0.010936f
C663 VTAIL.n312 B 0.01158f
C664 VTAIL.n313 B 0.025849f
C665 VTAIL.n314 B 0.025849f
C666 VTAIL.n315 B 0.01158f
C667 VTAIL.n316 B 0.010936f
C668 VTAIL.n317 B 0.020352f
C669 VTAIL.n318 B 0.020352f
C670 VTAIL.n319 B 0.010936f
C671 VTAIL.n320 B 0.01158f
C672 VTAIL.n321 B 0.025849f
C673 VTAIL.n322 B 0.058631f
C674 VTAIL.n323 B 0.01158f
C675 VTAIL.n324 B 0.010936f
C676 VTAIL.n325 B 0.045653f
C677 VTAIL.n326 B 0.033037f
C678 VTAIL.n327 B 1.37185f
C679 VN.t0 B 3.74189f
C680 VN.t1 B 4.33631f
.ends

