* NGSPICE file created from diff_pair_sample_0801.ext - technology: sky130A

.subckt diff_pair_sample_0801 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t18 VP.t0 VDD1.t5 w_n2926_n3438# sky130_fd_pr__pfet_01v8 ad=2.03775 pd=12.68 as=2.03775 ps=12.68 w=12.35 l=1.3
X1 VTAIL.t2 VN.t0 VDD2.t9 w_n2926_n3438# sky130_fd_pr__pfet_01v8 ad=2.03775 pd=12.68 as=2.03775 ps=12.68 w=12.35 l=1.3
X2 B.t11 B.t9 B.t10 w_n2926_n3438# sky130_fd_pr__pfet_01v8 ad=4.8165 pd=25.48 as=0 ps=0 w=12.35 l=1.3
X3 B.t8 B.t6 B.t7 w_n2926_n3438# sky130_fd_pr__pfet_01v8 ad=4.8165 pd=25.48 as=0 ps=0 w=12.35 l=1.3
X4 VDD1.t8 VP.t1 VTAIL.t17 w_n2926_n3438# sky130_fd_pr__pfet_01v8 ad=2.03775 pd=12.68 as=4.8165 ps=25.48 w=12.35 l=1.3
X5 VDD2.t8 VN.t1 VTAIL.t4 w_n2926_n3438# sky130_fd_pr__pfet_01v8 ad=4.8165 pd=25.48 as=2.03775 ps=12.68 w=12.35 l=1.3
X6 VTAIL.t16 VP.t2 VDD1.t2 w_n2926_n3438# sky130_fd_pr__pfet_01v8 ad=2.03775 pd=12.68 as=2.03775 ps=12.68 w=12.35 l=1.3
X7 VDD1.t7 VP.t3 VTAIL.t15 w_n2926_n3438# sky130_fd_pr__pfet_01v8 ad=2.03775 pd=12.68 as=4.8165 ps=25.48 w=12.35 l=1.3
X8 VTAIL.t14 VP.t4 VDD1.t9 w_n2926_n3438# sky130_fd_pr__pfet_01v8 ad=2.03775 pd=12.68 as=2.03775 ps=12.68 w=12.35 l=1.3
X9 VTAIL.t1 VN.t2 VDD2.t7 w_n2926_n3438# sky130_fd_pr__pfet_01v8 ad=2.03775 pd=12.68 as=2.03775 ps=12.68 w=12.35 l=1.3
X10 VDD2.t6 VN.t3 VTAIL.t3 w_n2926_n3438# sky130_fd_pr__pfet_01v8 ad=4.8165 pd=25.48 as=2.03775 ps=12.68 w=12.35 l=1.3
X11 VDD2.t5 VN.t4 VTAIL.t8 w_n2926_n3438# sky130_fd_pr__pfet_01v8 ad=2.03775 pd=12.68 as=4.8165 ps=25.48 w=12.35 l=1.3
X12 VDD1.t0 VP.t5 VTAIL.t13 w_n2926_n3438# sky130_fd_pr__pfet_01v8 ad=4.8165 pd=25.48 as=2.03775 ps=12.68 w=12.35 l=1.3
X13 B.t5 B.t3 B.t4 w_n2926_n3438# sky130_fd_pr__pfet_01v8 ad=4.8165 pd=25.48 as=0 ps=0 w=12.35 l=1.3
X14 VDD1.t6 VP.t6 VTAIL.t12 w_n2926_n3438# sky130_fd_pr__pfet_01v8 ad=2.03775 pd=12.68 as=2.03775 ps=12.68 w=12.35 l=1.3
X15 VTAIL.t0 VN.t5 VDD2.t4 w_n2926_n3438# sky130_fd_pr__pfet_01v8 ad=2.03775 pd=12.68 as=2.03775 ps=12.68 w=12.35 l=1.3
X16 VDD2.t3 VN.t6 VTAIL.t19 w_n2926_n3438# sky130_fd_pr__pfet_01v8 ad=2.03775 pd=12.68 as=2.03775 ps=12.68 w=12.35 l=1.3
X17 VDD1.t4 VP.t7 VTAIL.t11 w_n2926_n3438# sky130_fd_pr__pfet_01v8 ad=4.8165 pd=25.48 as=2.03775 ps=12.68 w=12.35 l=1.3
X18 VTAIL.t5 VN.t7 VDD2.t2 w_n2926_n3438# sky130_fd_pr__pfet_01v8 ad=2.03775 pd=12.68 as=2.03775 ps=12.68 w=12.35 l=1.3
X19 VTAIL.t10 VP.t8 VDD1.t3 w_n2926_n3438# sky130_fd_pr__pfet_01v8 ad=2.03775 pd=12.68 as=2.03775 ps=12.68 w=12.35 l=1.3
X20 B.t2 B.t0 B.t1 w_n2926_n3438# sky130_fd_pr__pfet_01v8 ad=4.8165 pd=25.48 as=0 ps=0 w=12.35 l=1.3
X21 VDD2.t1 VN.t8 VTAIL.t7 w_n2926_n3438# sky130_fd_pr__pfet_01v8 ad=2.03775 pd=12.68 as=4.8165 ps=25.48 w=12.35 l=1.3
X22 VDD2.t0 VN.t9 VTAIL.t6 w_n2926_n3438# sky130_fd_pr__pfet_01v8 ad=2.03775 pd=12.68 as=2.03775 ps=12.68 w=12.35 l=1.3
X23 VDD1.t1 VP.t9 VTAIL.t9 w_n2926_n3438# sky130_fd_pr__pfet_01v8 ad=2.03775 pd=12.68 as=2.03775 ps=12.68 w=12.35 l=1.3
R0 VP.n14 VP.t5 258.551
R1 VP.n3 VP.t9 228.951
R2 VP.n7 VP.t7 228.951
R3 VP.n5 VP.t2 228.951
R4 VP.n48 VP.t8 228.951
R5 VP.n55 VP.t3 228.951
R6 VP.n11 VP.t6 228.951
R7 VP.n31 VP.t1 228.951
R8 VP.n24 VP.t4 228.951
R9 VP.n13 VP.t0 228.951
R10 VP.n33 VP.n7 173.044
R11 VP.n56 VP.n55 173.044
R12 VP.n32 VP.n31 173.044
R13 VP.n16 VP.n15 161.3
R14 VP.n17 VP.n12 161.3
R15 VP.n19 VP.n18 161.3
R16 VP.n20 VP.n11 161.3
R17 VP.n22 VP.n21 161.3
R18 VP.n23 VP.n10 161.3
R19 VP.n26 VP.n25 161.3
R20 VP.n27 VP.n9 161.3
R21 VP.n29 VP.n28 161.3
R22 VP.n30 VP.n8 161.3
R23 VP.n54 VP.n0 161.3
R24 VP.n53 VP.n52 161.3
R25 VP.n51 VP.n1 161.3
R26 VP.n50 VP.n49 161.3
R27 VP.n47 VP.n2 161.3
R28 VP.n46 VP.n45 161.3
R29 VP.n44 VP.n3 161.3
R30 VP.n43 VP.n42 161.3
R31 VP.n41 VP.n4 161.3
R32 VP.n40 VP.n39 161.3
R33 VP.n38 VP.n37 161.3
R34 VP.n36 VP.n6 161.3
R35 VP.n35 VP.n34 161.3
R36 VP.n14 VP.n13 58.4685
R37 VP.n42 VP.n41 56.5193
R38 VP.n47 VP.n46 56.5193
R39 VP.n23 VP.n22 56.5193
R40 VP.n18 VP.n17 56.5193
R41 VP.n33 VP.n32 46.2316
R42 VP.n37 VP.n36 45.8354
R43 VP.n53 VP.n1 45.8354
R44 VP.n29 VP.n9 45.8354
R45 VP.n36 VP.n35 35.1514
R46 VP.n54 VP.n53 35.1514
R47 VP.n30 VP.n29 35.1514
R48 VP.n15 VP.n14 27.0985
R49 VP.n41 VP.n40 24.4675
R50 VP.n42 VP.n3 24.4675
R51 VP.n46 VP.n3 24.4675
R52 VP.n49 VP.n47 24.4675
R53 VP.n25 VP.n23 24.4675
R54 VP.n18 VP.n11 24.4675
R55 VP.n22 VP.n11 24.4675
R56 VP.n17 VP.n16 24.4675
R57 VP.n37 VP.n5 18.1061
R58 VP.n48 VP.n1 18.1061
R59 VP.n24 VP.n9 18.1061
R60 VP.n35 VP.n7 12.7233
R61 VP.n55 VP.n54 12.7233
R62 VP.n31 VP.n30 12.7233
R63 VP.n40 VP.n5 6.36192
R64 VP.n49 VP.n48 6.36192
R65 VP.n25 VP.n24 6.36192
R66 VP.n16 VP.n13 6.36192
R67 VP.n15 VP.n12 0.189894
R68 VP.n19 VP.n12 0.189894
R69 VP.n20 VP.n19 0.189894
R70 VP.n21 VP.n20 0.189894
R71 VP.n21 VP.n10 0.189894
R72 VP.n26 VP.n10 0.189894
R73 VP.n27 VP.n26 0.189894
R74 VP.n28 VP.n27 0.189894
R75 VP.n28 VP.n8 0.189894
R76 VP.n32 VP.n8 0.189894
R77 VP.n34 VP.n33 0.189894
R78 VP.n34 VP.n6 0.189894
R79 VP.n38 VP.n6 0.189894
R80 VP.n39 VP.n38 0.189894
R81 VP.n39 VP.n4 0.189894
R82 VP.n43 VP.n4 0.189894
R83 VP.n44 VP.n43 0.189894
R84 VP.n45 VP.n44 0.189894
R85 VP.n45 VP.n2 0.189894
R86 VP.n50 VP.n2 0.189894
R87 VP.n51 VP.n50 0.189894
R88 VP.n52 VP.n51 0.189894
R89 VP.n52 VP.n0 0.189894
R90 VP.n56 VP.n0 0.189894
R91 VP VP.n56 0.0516364
R92 VDD1.n1 VDD1.t0 81.5211
R93 VDD1.n3 VDD1.t4 81.5201
R94 VDD1.n5 VDD1.n4 78.4823
R95 VDD1.n1 VDD1.n0 77.484
R96 VDD1.n3 VDD1.n2 77.4838
R97 VDD1.n7 VDD1.n6 77.4828
R98 VDD1.n7 VDD1.n5 42.322
R99 VDD1.n6 VDD1.t9 2.63248
R100 VDD1.n6 VDD1.t8 2.63248
R101 VDD1.n0 VDD1.t5 2.63248
R102 VDD1.n0 VDD1.t6 2.63248
R103 VDD1.n4 VDD1.t3 2.63248
R104 VDD1.n4 VDD1.t7 2.63248
R105 VDD1.n2 VDD1.t2 2.63248
R106 VDD1.n2 VDD1.t1 2.63248
R107 VDD1 VDD1.n7 0.99619
R108 VDD1 VDD1.n1 0.409983
R109 VDD1.n5 VDD1.n3 0.296447
R110 VTAIL.n11 VTAIL.t8 63.4372
R111 VTAIL.n17 VTAIL.t7 63.4361
R112 VTAIL.n2 VTAIL.t15 63.4361
R113 VTAIL.n16 VTAIL.t17 63.436
R114 VTAIL.n15 VTAIL.n14 60.8052
R115 VTAIL.n13 VTAIL.n12 60.8052
R116 VTAIL.n10 VTAIL.n9 60.8052
R117 VTAIL.n8 VTAIL.n7 60.8052
R118 VTAIL.n19 VTAIL.n18 60.805
R119 VTAIL.n1 VTAIL.n0 60.805
R120 VTAIL.n4 VTAIL.n3 60.805
R121 VTAIL.n6 VTAIL.n5 60.805
R122 VTAIL.n8 VTAIL.n6 25.8238
R123 VTAIL.n17 VTAIL.n16 24.4186
R124 VTAIL.n18 VTAIL.t6 2.63248
R125 VTAIL.n18 VTAIL.t1 2.63248
R126 VTAIL.n0 VTAIL.t4 2.63248
R127 VTAIL.n0 VTAIL.t5 2.63248
R128 VTAIL.n3 VTAIL.t9 2.63248
R129 VTAIL.n3 VTAIL.t10 2.63248
R130 VTAIL.n5 VTAIL.t11 2.63248
R131 VTAIL.n5 VTAIL.t16 2.63248
R132 VTAIL.n14 VTAIL.t12 2.63248
R133 VTAIL.n14 VTAIL.t14 2.63248
R134 VTAIL.n12 VTAIL.t13 2.63248
R135 VTAIL.n12 VTAIL.t18 2.63248
R136 VTAIL.n9 VTAIL.t19 2.63248
R137 VTAIL.n9 VTAIL.t2 2.63248
R138 VTAIL.n7 VTAIL.t3 2.63248
R139 VTAIL.n7 VTAIL.t0 2.63248
R140 VTAIL.n10 VTAIL.n8 1.40567
R141 VTAIL.n11 VTAIL.n10 1.40567
R142 VTAIL.n15 VTAIL.n13 1.40567
R143 VTAIL.n16 VTAIL.n15 1.40567
R144 VTAIL.n6 VTAIL.n4 1.40567
R145 VTAIL.n4 VTAIL.n2 1.40567
R146 VTAIL.n19 VTAIL.n17 1.40567
R147 VTAIL.n13 VTAIL.n11 1.17291
R148 VTAIL.n2 VTAIL.n1 1.17291
R149 VTAIL VTAIL.n1 1.11257
R150 VTAIL VTAIL.n19 0.293603
R151 VN.n6 VN.t1 258.551
R152 VN.n32 VN.t4 258.551
R153 VN.n3 VN.t9 228.951
R154 VN.n5 VN.t7 228.951
R155 VN.n16 VN.t2 228.951
R156 VN.n23 VN.t8 228.951
R157 VN.n29 VN.t6 228.951
R158 VN.n31 VN.t0 228.951
R159 VN.n28 VN.t5 228.951
R160 VN.n48 VN.t3 228.951
R161 VN.n24 VN.n23 173.044
R162 VN.n49 VN.n48 173.044
R163 VN.n47 VN.n25 161.3
R164 VN.n46 VN.n45 161.3
R165 VN.n44 VN.n26 161.3
R166 VN.n43 VN.n42 161.3
R167 VN.n41 VN.n27 161.3
R168 VN.n40 VN.n39 161.3
R169 VN.n38 VN.n29 161.3
R170 VN.n37 VN.n36 161.3
R171 VN.n35 VN.n30 161.3
R172 VN.n34 VN.n33 161.3
R173 VN.n22 VN.n0 161.3
R174 VN.n21 VN.n20 161.3
R175 VN.n19 VN.n1 161.3
R176 VN.n18 VN.n17 161.3
R177 VN.n15 VN.n2 161.3
R178 VN.n14 VN.n13 161.3
R179 VN.n12 VN.n3 161.3
R180 VN.n11 VN.n10 161.3
R181 VN.n9 VN.n4 161.3
R182 VN.n8 VN.n7 161.3
R183 VN.n6 VN.n5 58.4685
R184 VN.n32 VN.n31 58.4685
R185 VN.n10 VN.n9 56.5193
R186 VN.n15 VN.n14 56.5193
R187 VN.n36 VN.n35 56.5193
R188 VN.n41 VN.n40 56.5193
R189 VN VN.n49 46.6122
R190 VN.n21 VN.n1 45.8354
R191 VN.n46 VN.n26 45.8354
R192 VN.n22 VN.n21 35.1514
R193 VN.n47 VN.n46 35.1514
R194 VN.n33 VN.n32 27.0985
R195 VN.n7 VN.n6 27.0985
R196 VN.n9 VN.n8 24.4675
R197 VN.n10 VN.n3 24.4675
R198 VN.n14 VN.n3 24.4675
R199 VN.n17 VN.n15 24.4675
R200 VN.n35 VN.n34 24.4675
R201 VN.n40 VN.n29 24.4675
R202 VN.n36 VN.n29 24.4675
R203 VN.n42 VN.n41 24.4675
R204 VN.n16 VN.n1 18.1061
R205 VN.n28 VN.n26 18.1061
R206 VN.n23 VN.n22 12.7233
R207 VN.n48 VN.n47 12.7233
R208 VN.n8 VN.n5 6.36192
R209 VN.n17 VN.n16 6.36192
R210 VN.n34 VN.n31 6.36192
R211 VN.n42 VN.n28 6.36192
R212 VN.n49 VN.n25 0.189894
R213 VN.n45 VN.n25 0.189894
R214 VN.n45 VN.n44 0.189894
R215 VN.n44 VN.n43 0.189894
R216 VN.n43 VN.n27 0.189894
R217 VN.n39 VN.n27 0.189894
R218 VN.n39 VN.n38 0.189894
R219 VN.n38 VN.n37 0.189894
R220 VN.n37 VN.n30 0.189894
R221 VN.n33 VN.n30 0.189894
R222 VN.n7 VN.n4 0.189894
R223 VN.n11 VN.n4 0.189894
R224 VN.n12 VN.n11 0.189894
R225 VN.n13 VN.n12 0.189894
R226 VN.n13 VN.n2 0.189894
R227 VN.n18 VN.n2 0.189894
R228 VN.n19 VN.n18 0.189894
R229 VN.n20 VN.n19 0.189894
R230 VN.n20 VN.n0 0.189894
R231 VN.n24 VN.n0 0.189894
R232 VN VN.n24 0.0516364
R233 VDD2.n1 VDD2.t8 81.5201
R234 VDD2.n4 VDD2.t6 80.116
R235 VDD2.n3 VDD2.n2 78.4823
R236 VDD2 VDD2.n7 78.4785
R237 VDD2.n6 VDD2.n5 77.484
R238 VDD2.n1 VDD2.n0 77.4838
R239 VDD2.n4 VDD2.n3 41.0364
R240 VDD2.n7 VDD2.t9 2.63248
R241 VDD2.n7 VDD2.t5 2.63248
R242 VDD2.n5 VDD2.t4 2.63248
R243 VDD2.n5 VDD2.t3 2.63248
R244 VDD2.n2 VDD2.t7 2.63248
R245 VDD2.n2 VDD2.t1 2.63248
R246 VDD2.n0 VDD2.t2 2.63248
R247 VDD2.n0 VDD2.t0 2.63248
R248 VDD2.n6 VDD2.n4 1.40567
R249 VDD2 VDD2.n6 0.409983
R250 VDD2.n3 VDD2.n1 0.296447
R251 B.n491 B.n72 585
R252 B.n493 B.n492 585
R253 B.n494 B.n71 585
R254 B.n496 B.n495 585
R255 B.n497 B.n70 585
R256 B.n499 B.n498 585
R257 B.n500 B.n69 585
R258 B.n502 B.n501 585
R259 B.n503 B.n68 585
R260 B.n505 B.n504 585
R261 B.n506 B.n67 585
R262 B.n508 B.n507 585
R263 B.n509 B.n66 585
R264 B.n511 B.n510 585
R265 B.n512 B.n65 585
R266 B.n514 B.n513 585
R267 B.n515 B.n64 585
R268 B.n517 B.n516 585
R269 B.n518 B.n63 585
R270 B.n520 B.n519 585
R271 B.n521 B.n62 585
R272 B.n523 B.n522 585
R273 B.n524 B.n61 585
R274 B.n526 B.n525 585
R275 B.n527 B.n60 585
R276 B.n529 B.n528 585
R277 B.n530 B.n59 585
R278 B.n532 B.n531 585
R279 B.n533 B.n58 585
R280 B.n535 B.n534 585
R281 B.n536 B.n57 585
R282 B.n538 B.n537 585
R283 B.n539 B.n56 585
R284 B.n541 B.n540 585
R285 B.n542 B.n55 585
R286 B.n544 B.n543 585
R287 B.n545 B.n54 585
R288 B.n547 B.n546 585
R289 B.n548 B.n53 585
R290 B.n550 B.n549 585
R291 B.n551 B.n52 585
R292 B.n553 B.n552 585
R293 B.n554 B.n49 585
R294 B.n557 B.n556 585
R295 B.n558 B.n48 585
R296 B.n560 B.n559 585
R297 B.n561 B.n47 585
R298 B.n563 B.n562 585
R299 B.n564 B.n46 585
R300 B.n566 B.n565 585
R301 B.n567 B.n45 585
R302 B.n569 B.n568 585
R303 B.n571 B.n570 585
R304 B.n572 B.n41 585
R305 B.n574 B.n573 585
R306 B.n575 B.n40 585
R307 B.n577 B.n576 585
R308 B.n578 B.n39 585
R309 B.n580 B.n579 585
R310 B.n581 B.n38 585
R311 B.n583 B.n582 585
R312 B.n584 B.n37 585
R313 B.n586 B.n585 585
R314 B.n587 B.n36 585
R315 B.n589 B.n588 585
R316 B.n590 B.n35 585
R317 B.n592 B.n591 585
R318 B.n593 B.n34 585
R319 B.n595 B.n594 585
R320 B.n596 B.n33 585
R321 B.n598 B.n597 585
R322 B.n599 B.n32 585
R323 B.n601 B.n600 585
R324 B.n602 B.n31 585
R325 B.n604 B.n603 585
R326 B.n605 B.n30 585
R327 B.n607 B.n606 585
R328 B.n608 B.n29 585
R329 B.n610 B.n609 585
R330 B.n611 B.n28 585
R331 B.n613 B.n612 585
R332 B.n614 B.n27 585
R333 B.n616 B.n615 585
R334 B.n617 B.n26 585
R335 B.n619 B.n618 585
R336 B.n620 B.n25 585
R337 B.n622 B.n621 585
R338 B.n623 B.n24 585
R339 B.n625 B.n624 585
R340 B.n626 B.n23 585
R341 B.n628 B.n627 585
R342 B.n629 B.n22 585
R343 B.n631 B.n630 585
R344 B.n632 B.n21 585
R345 B.n634 B.n633 585
R346 B.n490 B.n489 585
R347 B.n488 B.n73 585
R348 B.n487 B.n486 585
R349 B.n485 B.n74 585
R350 B.n484 B.n483 585
R351 B.n482 B.n75 585
R352 B.n481 B.n480 585
R353 B.n479 B.n76 585
R354 B.n478 B.n477 585
R355 B.n476 B.n77 585
R356 B.n475 B.n474 585
R357 B.n473 B.n78 585
R358 B.n472 B.n471 585
R359 B.n470 B.n79 585
R360 B.n469 B.n468 585
R361 B.n467 B.n80 585
R362 B.n466 B.n465 585
R363 B.n464 B.n81 585
R364 B.n463 B.n462 585
R365 B.n461 B.n82 585
R366 B.n460 B.n459 585
R367 B.n458 B.n83 585
R368 B.n457 B.n456 585
R369 B.n455 B.n84 585
R370 B.n454 B.n453 585
R371 B.n452 B.n85 585
R372 B.n451 B.n450 585
R373 B.n449 B.n86 585
R374 B.n448 B.n447 585
R375 B.n446 B.n87 585
R376 B.n445 B.n444 585
R377 B.n443 B.n88 585
R378 B.n442 B.n441 585
R379 B.n440 B.n89 585
R380 B.n439 B.n438 585
R381 B.n437 B.n90 585
R382 B.n436 B.n435 585
R383 B.n434 B.n91 585
R384 B.n433 B.n432 585
R385 B.n431 B.n92 585
R386 B.n430 B.n429 585
R387 B.n428 B.n93 585
R388 B.n427 B.n426 585
R389 B.n425 B.n94 585
R390 B.n424 B.n423 585
R391 B.n422 B.n95 585
R392 B.n421 B.n420 585
R393 B.n419 B.n96 585
R394 B.n418 B.n417 585
R395 B.n416 B.n97 585
R396 B.n415 B.n414 585
R397 B.n413 B.n98 585
R398 B.n412 B.n411 585
R399 B.n410 B.n99 585
R400 B.n409 B.n408 585
R401 B.n407 B.n100 585
R402 B.n406 B.n405 585
R403 B.n404 B.n101 585
R404 B.n403 B.n402 585
R405 B.n401 B.n102 585
R406 B.n400 B.n399 585
R407 B.n398 B.n103 585
R408 B.n397 B.n396 585
R409 B.n395 B.n104 585
R410 B.n394 B.n393 585
R411 B.n392 B.n105 585
R412 B.n391 B.n390 585
R413 B.n389 B.n106 585
R414 B.n388 B.n387 585
R415 B.n386 B.n107 585
R416 B.n385 B.n384 585
R417 B.n383 B.n108 585
R418 B.n382 B.n381 585
R419 B.n380 B.n109 585
R420 B.n379 B.n378 585
R421 B.n235 B.n234 585
R422 B.n236 B.n161 585
R423 B.n238 B.n237 585
R424 B.n239 B.n160 585
R425 B.n241 B.n240 585
R426 B.n242 B.n159 585
R427 B.n244 B.n243 585
R428 B.n245 B.n158 585
R429 B.n247 B.n246 585
R430 B.n248 B.n157 585
R431 B.n250 B.n249 585
R432 B.n251 B.n156 585
R433 B.n253 B.n252 585
R434 B.n254 B.n155 585
R435 B.n256 B.n255 585
R436 B.n257 B.n154 585
R437 B.n259 B.n258 585
R438 B.n260 B.n153 585
R439 B.n262 B.n261 585
R440 B.n263 B.n152 585
R441 B.n265 B.n264 585
R442 B.n266 B.n151 585
R443 B.n268 B.n267 585
R444 B.n269 B.n150 585
R445 B.n271 B.n270 585
R446 B.n272 B.n149 585
R447 B.n274 B.n273 585
R448 B.n275 B.n148 585
R449 B.n277 B.n276 585
R450 B.n278 B.n147 585
R451 B.n280 B.n279 585
R452 B.n281 B.n146 585
R453 B.n283 B.n282 585
R454 B.n284 B.n145 585
R455 B.n286 B.n285 585
R456 B.n287 B.n144 585
R457 B.n289 B.n288 585
R458 B.n290 B.n143 585
R459 B.n292 B.n291 585
R460 B.n293 B.n142 585
R461 B.n295 B.n294 585
R462 B.n296 B.n141 585
R463 B.n298 B.n297 585
R464 B.n300 B.n299 585
R465 B.n301 B.n137 585
R466 B.n303 B.n302 585
R467 B.n304 B.n136 585
R468 B.n306 B.n305 585
R469 B.n307 B.n135 585
R470 B.n309 B.n308 585
R471 B.n310 B.n134 585
R472 B.n312 B.n311 585
R473 B.n314 B.n131 585
R474 B.n316 B.n315 585
R475 B.n317 B.n130 585
R476 B.n319 B.n318 585
R477 B.n320 B.n129 585
R478 B.n322 B.n321 585
R479 B.n323 B.n128 585
R480 B.n325 B.n324 585
R481 B.n326 B.n127 585
R482 B.n328 B.n327 585
R483 B.n329 B.n126 585
R484 B.n331 B.n330 585
R485 B.n332 B.n125 585
R486 B.n334 B.n333 585
R487 B.n335 B.n124 585
R488 B.n337 B.n336 585
R489 B.n338 B.n123 585
R490 B.n340 B.n339 585
R491 B.n341 B.n122 585
R492 B.n343 B.n342 585
R493 B.n344 B.n121 585
R494 B.n346 B.n345 585
R495 B.n347 B.n120 585
R496 B.n349 B.n348 585
R497 B.n350 B.n119 585
R498 B.n352 B.n351 585
R499 B.n353 B.n118 585
R500 B.n355 B.n354 585
R501 B.n356 B.n117 585
R502 B.n358 B.n357 585
R503 B.n359 B.n116 585
R504 B.n361 B.n360 585
R505 B.n362 B.n115 585
R506 B.n364 B.n363 585
R507 B.n365 B.n114 585
R508 B.n367 B.n366 585
R509 B.n368 B.n113 585
R510 B.n370 B.n369 585
R511 B.n371 B.n112 585
R512 B.n373 B.n372 585
R513 B.n374 B.n111 585
R514 B.n376 B.n375 585
R515 B.n377 B.n110 585
R516 B.n233 B.n162 585
R517 B.n232 B.n231 585
R518 B.n230 B.n163 585
R519 B.n229 B.n228 585
R520 B.n227 B.n164 585
R521 B.n226 B.n225 585
R522 B.n224 B.n165 585
R523 B.n223 B.n222 585
R524 B.n221 B.n166 585
R525 B.n220 B.n219 585
R526 B.n218 B.n167 585
R527 B.n217 B.n216 585
R528 B.n215 B.n168 585
R529 B.n214 B.n213 585
R530 B.n212 B.n169 585
R531 B.n211 B.n210 585
R532 B.n209 B.n170 585
R533 B.n208 B.n207 585
R534 B.n206 B.n171 585
R535 B.n205 B.n204 585
R536 B.n203 B.n172 585
R537 B.n202 B.n201 585
R538 B.n200 B.n173 585
R539 B.n199 B.n198 585
R540 B.n197 B.n174 585
R541 B.n196 B.n195 585
R542 B.n194 B.n175 585
R543 B.n193 B.n192 585
R544 B.n191 B.n176 585
R545 B.n190 B.n189 585
R546 B.n188 B.n177 585
R547 B.n187 B.n186 585
R548 B.n185 B.n178 585
R549 B.n184 B.n183 585
R550 B.n182 B.n179 585
R551 B.n181 B.n180 585
R552 B.n2 B.n0 585
R553 B.n689 B.n1 585
R554 B.n688 B.n687 585
R555 B.n686 B.n3 585
R556 B.n685 B.n684 585
R557 B.n683 B.n4 585
R558 B.n682 B.n681 585
R559 B.n680 B.n5 585
R560 B.n679 B.n678 585
R561 B.n677 B.n6 585
R562 B.n676 B.n675 585
R563 B.n674 B.n7 585
R564 B.n673 B.n672 585
R565 B.n671 B.n8 585
R566 B.n670 B.n669 585
R567 B.n668 B.n9 585
R568 B.n667 B.n666 585
R569 B.n665 B.n10 585
R570 B.n664 B.n663 585
R571 B.n662 B.n11 585
R572 B.n661 B.n660 585
R573 B.n659 B.n12 585
R574 B.n658 B.n657 585
R575 B.n656 B.n13 585
R576 B.n655 B.n654 585
R577 B.n653 B.n14 585
R578 B.n652 B.n651 585
R579 B.n650 B.n15 585
R580 B.n649 B.n648 585
R581 B.n647 B.n16 585
R582 B.n646 B.n645 585
R583 B.n644 B.n17 585
R584 B.n643 B.n642 585
R585 B.n641 B.n18 585
R586 B.n640 B.n639 585
R587 B.n638 B.n19 585
R588 B.n637 B.n636 585
R589 B.n635 B.n20 585
R590 B.n691 B.n690 585
R591 B.n234 B.n233 468.476
R592 B.n635 B.n634 468.476
R593 B.n378 B.n377 468.476
R594 B.n491 B.n490 468.476
R595 B.n132 B.t0 433.558
R596 B.n138 B.t3 433.558
R597 B.n42 B.t9 433.558
R598 B.n50 B.t6 433.558
R599 B.n233 B.n232 163.367
R600 B.n232 B.n163 163.367
R601 B.n228 B.n163 163.367
R602 B.n228 B.n227 163.367
R603 B.n227 B.n226 163.367
R604 B.n226 B.n165 163.367
R605 B.n222 B.n165 163.367
R606 B.n222 B.n221 163.367
R607 B.n221 B.n220 163.367
R608 B.n220 B.n167 163.367
R609 B.n216 B.n167 163.367
R610 B.n216 B.n215 163.367
R611 B.n215 B.n214 163.367
R612 B.n214 B.n169 163.367
R613 B.n210 B.n169 163.367
R614 B.n210 B.n209 163.367
R615 B.n209 B.n208 163.367
R616 B.n208 B.n171 163.367
R617 B.n204 B.n171 163.367
R618 B.n204 B.n203 163.367
R619 B.n203 B.n202 163.367
R620 B.n202 B.n173 163.367
R621 B.n198 B.n173 163.367
R622 B.n198 B.n197 163.367
R623 B.n197 B.n196 163.367
R624 B.n196 B.n175 163.367
R625 B.n192 B.n175 163.367
R626 B.n192 B.n191 163.367
R627 B.n191 B.n190 163.367
R628 B.n190 B.n177 163.367
R629 B.n186 B.n177 163.367
R630 B.n186 B.n185 163.367
R631 B.n185 B.n184 163.367
R632 B.n184 B.n179 163.367
R633 B.n180 B.n179 163.367
R634 B.n180 B.n2 163.367
R635 B.n690 B.n2 163.367
R636 B.n690 B.n689 163.367
R637 B.n689 B.n688 163.367
R638 B.n688 B.n3 163.367
R639 B.n684 B.n3 163.367
R640 B.n684 B.n683 163.367
R641 B.n683 B.n682 163.367
R642 B.n682 B.n5 163.367
R643 B.n678 B.n5 163.367
R644 B.n678 B.n677 163.367
R645 B.n677 B.n676 163.367
R646 B.n676 B.n7 163.367
R647 B.n672 B.n7 163.367
R648 B.n672 B.n671 163.367
R649 B.n671 B.n670 163.367
R650 B.n670 B.n9 163.367
R651 B.n666 B.n9 163.367
R652 B.n666 B.n665 163.367
R653 B.n665 B.n664 163.367
R654 B.n664 B.n11 163.367
R655 B.n660 B.n11 163.367
R656 B.n660 B.n659 163.367
R657 B.n659 B.n658 163.367
R658 B.n658 B.n13 163.367
R659 B.n654 B.n13 163.367
R660 B.n654 B.n653 163.367
R661 B.n653 B.n652 163.367
R662 B.n652 B.n15 163.367
R663 B.n648 B.n15 163.367
R664 B.n648 B.n647 163.367
R665 B.n647 B.n646 163.367
R666 B.n646 B.n17 163.367
R667 B.n642 B.n17 163.367
R668 B.n642 B.n641 163.367
R669 B.n641 B.n640 163.367
R670 B.n640 B.n19 163.367
R671 B.n636 B.n19 163.367
R672 B.n636 B.n635 163.367
R673 B.n234 B.n161 163.367
R674 B.n238 B.n161 163.367
R675 B.n239 B.n238 163.367
R676 B.n240 B.n239 163.367
R677 B.n240 B.n159 163.367
R678 B.n244 B.n159 163.367
R679 B.n245 B.n244 163.367
R680 B.n246 B.n245 163.367
R681 B.n246 B.n157 163.367
R682 B.n250 B.n157 163.367
R683 B.n251 B.n250 163.367
R684 B.n252 B.n251 163.367
R685 B.n252 B.n155 163.367
R686 B.n256 B.n155 163.367
R687 B.n257 B.n256 163.367
R688 B.n258 B.n257 163.367
R689 B.n258 B.n153 163.367
R690 B.n262 B.n153 163.367
R691 B.n263 B.n262 163.367
R692 B.n264 B.n263 163.367
R693 B.n264 B.n151 163.367
R694 B.n268 B.n151 163.367
R695 B.n269 B.n268 163.367
R696 B.n270 B.n269 163.367
R697 B.n270 B.n149 163.367
R698 B.n274 B.n149 163.367
R699 B.n275 B.n274 163.367
R700 B.n276 B.n275 163.367
R701 B.n276 B.n147 163.367
R702 B.n280 B.n147 163.367
R703 B.n281 B.n280 163.367
R704 B.n282 B.n281 163.367
R705 B.n282 B.n145 163.367
R706 B.n286 B.n145 163.367
R707 B.n287 B.n286 163.367
R708 B.n288 B.n287 163.367
R709 B.n288 B.n143 163.367
R710 B.n292 B.n143 163.367
R711 B.n293 B.n292 163.367
R712 B.n294 B.n293 163.367
R713 B.n294 B.n141 163.367
R714 B.n298 B.n141 163.367
R715 B.n299 B.n298 163.367
R716 B.n299 B.n137 163.367
R717 B.n303 B.n137 163.367
R718 B.n304 B.n303 163.367
R719 B.n305 B.n304 163.367
R720 B.n305 B.n135 163.367
R721 B.n309 B.n135 163.367
R722 B.n310 B.n309 163.367
R723 B.n311 B.n310 163.367
R724 B.n311 B.n131 163.367
R725 B.n316 B.n131 163.367
R726 B.n317 B.n316 163.367
R727 B.n318 B.n317 163.367
R728 B.n318 B.n129 163.367
R729 B.n322 B.n129 163.367
R730 B.n323 B.n322 163.367
R731 B.n324 B.n323 163.367
R732 B.n324 B.n127 163.367
R733 B.n328 B.n127 163.367
R734 B.n329 B.n328 163.367
R735 B.n330 B.n329 163.367
R736 B.n330 B.n125 163.367
R737 B.n334 B.n125 163.367
R738 B.n335 B.n334 163.367
R739 B.n336 B.n335 163.367
R740 B.n336 B.n123 163.367
R741 B.n340 B.n123 163.367
R742 B.n341 B.n340 163.367
R743 B.n342 B.n341 163.367
R744 B.n342 B.n121 163.367
R745 B.n346 B.n121 163.367
R746 B.n347 B.n346 163.367
R747 B.n348 B.n347 163.367
R748 B.n348 B.n119 163.367
R749 B.n352 B.n119 163.367
R750 B.n353 B.n352 163.367
R751 B.n354 B.n353 163.367
R752 B.n354 B.n117 163.367
R753 B.n358 B.n117 163.367
R754 B.n359 B.n358 163.367
R755 B.n360 B.n359 163.367
R756 B.n360 B.n115 163.367
R757 B.n364 B.n115 163.367
R758 B.n365 B.n364 163.367
R759 B.n366 B.n365 163.367
R760 B.n366 B.n113 163.367
R761 B.n370 B.n113 163.367
R762 B.n371 B.n370 163.367
R763 B.n372 B.n371 163.367
R764 B.n372 B.n111 163.367
R765 B.n376 B.n111 163.367
R766 B.n377 B.n376 163.367
R767 B.n378 B.n109 163.367
R768 B.n382 B.n109 163.367
R769 B.n383 B.n382 163.367
R770 B.n384 B.n383 163.367
R771 B.n384 B.n107 163.367
R772 B.n388 B.n107 163.367
R773 B.n389 B.n388 163.367
R774 B.n390 B.n389 163.367
R775 B.n390 B.n105 163.367
R776 B.n394 B.n105 163.367
R777 B.n395 B.n394 163.367
R778 B.n396 B.n395 163.367
R779 B.n396 B.n103 163.367
R780 B.n400 B.n103 163.367
R781 B.n401 B.n400 163.367
R782 B.n402 B.n401 163.367
R783 B.n402 B.n101 163.367
R784 B.n406 B.n101 163.367
R785 B.n407 B.n406 163.367
R786 B.n408 B.n407 163.367
R787 B.n408 B.n99 163.367
R788 B.n412 B.n99 163.367
R789 B.n413 B.n412 163.367
R790 B.n414 B.n413 163.367
R791 B.n414 B.n97 163.367
R792 B.n418 B.n97 163.367
R793 B.n419 B.n418 163.367
R794 B.n420 B.n419 163.367
R795 B.n420 B.n95 163.367
R796 B.n424 B.n95 163.367
R797 B.n425 B.n424 163.367
R798 B.n426 B.n425 163.367
R799 B.n426 B.n93 163.367
R800 B.n430 B.n93 163.367
R801 B.n431 B.n430 163.367
R802 B.n432 B.n431 163.367
R803 B.n432 B.n91 163.367
R804 B.n436 B.n91 163.367
R805 B.n437 B.n436 163.367
R806 B.n438 B.n437 163.367
R807 B.n438 B.n89 163.367
R808 B.n442 B.n89 163.367
R809 B.n443 B.n442 163.367
R810 B.n444 B.n443 163.367
R811 B.n444 B.n87 163.367
R812 B.n448 B.n87 163.367
R813 B.n449 B.n448 163.367
R814 B.n450 B.n449 163.367
R815 B.n450 B.n85 163.367
R816 B.n454 B.n85 163.367
R817 B.n455 B.n454 163.367
R818 B.n456 B.n455 163.367
R819 B.n456 B.n83 163.367
R820 B.n460 B.n83 163.367
R821 B.n461 B.n460 163.367
R822 B.n462 B.n461 163.367
R823 B.n462 B.n81 163.367
R824 B.n466 B.n81 163.367
R825 B.n467 B.n466 163.367
R826 B.n468 B.n467 163.367
R827 B.n468 B.n79 163.367
R828 B.n472 B.n79 163.367
R829 B.n473 B.n472 163.367
R830 B.n474 B.n473 163.367
R831 B.n474 B.n77 163.367
R832 B.n478 B.n77 163.367
R833 B.n479 B.n478 163.367
R834 B.n480 B.n479 163.367
R835 B.n480 B.n75 163.367
R836 B.n484 B.n75 163.367
R837 B.n485 B.n484 163.367
R838 B.n486 B.n485 163.367
R839 B.n486 B.n73 163.367
R840 B.n490 B.n73 163.367
R841 B.n634 B.n21 163.367
R842 B.n630 B.n21 163.367
R843 B.n630 B.n629 163.367
R844 B.n629 B.n628 163.367
R845 B.n628 B.n23 163.367
R846 B.n624 B.n23 163.367
R847 B.n624 B.n623 163.367
R848 B.n623 B.n622 163.367
R849 B.n622 B.n25 163.367
R850 B.n618 B.n25 163.367
R851 B.n618 B.n617 163.367
R852 B.n617 B.n616 163.367
R853 B.n616 B.n27 163.367
R854 B.n612 B.n27 163.367
R855 B.n612 B.n611 163.367
R856 B.n611 B.n610 163.367
R857 B.n610 B.n29 163.367
R858 B.n606 B.n29 163.367
R859 B.n606 B.n605 163.367
R860 B.n605 B.n604 163.367
R861 B.n604 B.n31 163.367
R862 B.n600 B.n31 163.367
R863 B.n600 B.n599 163.367
R864 B.n599 B.n598 163.367
R865 B.n598 B.n33 163.367
R866 B.n594 B.n33 163.367
R867 B.n594 B.n593 163.367
R868 B.n593 B.n592 163.367
R869 B.n592 B.n35 163.367
R870 B.n588 B.n35 163.367
R871 B.n588 B.n587 163.367
R872 B.n587 B.n586 163.367
R873 B.n586 B.n37 163.367
R874 B.n582 B.n37 163.367
R875 B.n582 B.n581 163.367
R876 B.n581 B.n580 163.367
R877 B.n580 B.n39 163.367
R878 B.n576 B.n39 163.367
R879 B.n576 B.n575 163.367
R880 B.n575 B.n574 163.367
R881 B.n574 B.n41 163.367
R882 B.n570 B.n41 163.367
R883 B.n570 B.n569 163.367
R884 B.n569 B.n45 163.367
R885 B.n565 B.n45 163.367
R886 B.n565 B.n564 163.367
R887 B.n564 B.n563 163.367
R888 B.n563 B.n47 163.367
R889 B.n559 B.n47 163.367
R890 B.n559 B.n558 163.367
R891 B.n558 B.n557 163.367
R892 B.n557 B.n49 163.367
R893 B.n552 B.n49 163.367
R894 B.n552 B.n551 163.367
R895 B.n551 B.n550 163.367
R896 B.n550 B.n53 163.367
R897 B.n546 B.n53 163.367
R898 B.n546 B.n545 163.367
R899 B.n545 B.n544 163.367
R900 B.n544 B.n55 163.367
R901 B.n540 B.n55 163.367
R902 B.n540 B.n539 163.367
R903 B.n539 B.n538 163.367
R904 B.n538 B.n57 163.367
R905 B.n534 B.n57 163.367
R906 B.n534 B.n533 163.367
R907 B.n533 B.n532 163.367
R908 B.n532 B.n59 163.367
R909 B.n528 B.n59 163.367
R910 B.n528 B.n527 163.367
R911 B.n527 B.n526 163.367
R912 B.n526 B.n61 163.367
R913 B.n522 B.n61 163.367
R914 B.n522 B.n521 163.367
R915 B.n521 B.n520 163.367
R916 B.n520 B.n63 163.367
R917 B.n516 B.n63 163.367
R918 B.n516 B.n515 163.367
R919 B.n515 B.n514 163.367
R920 B.n514 B.n65 163.367
R921 B.n510 B.n65 163.367
R922 B.n510 B.n509 163.367
R923 B.n509 B.n508 163.367
R924 B.n508 B.n67 163.367
R925 B.n504 B.n67 163.367
R926 B.n504 B.n503 163.367
R927 B.n503 B.n502 163.367
R928 B.n502 B.n69 163.367
R929 B.n498 B.n69 163.367
R930 B.n498 B.n497 163.367
R931 B.n497 B.n496 163.367
R932 B.n496 B.n71 163.367
R933 B.n492 B.n71 163.367
R934 B.n492 B.n491 163.367
R935 B.n132 B.t2 140.773
R936 B.n50 B.t7 140.773
R937 B.n138 B.t5 140.757
R938 B.n42 B.t10 140.757
R939 B.n133 B.t1 109.16
R940 B.n51 B.t8 109.16
R941 B.n139 B.t4 109.145
R942 B.n43 B.t11 109.145
R943 B.n313 B.n133 59.5399
R944 B.n140 B.n139 59.5399
R945 B.n44 B.n43 59.5399
R946 B.n555 B.n51 59.5399
R947 B.n133 B.n132 31.6126
R948 B.n139 B.n138 31.6126
R949 B.n43 B.n42 31.6126
R950 B.n51 B.n50 31.6126
R951 B.n633 B.n20 30.4395
R952 B.n489 B.n72 30.4395
R953 B.n379 B.n110 30.4395
R954 B.n235 B.n162 30.4395
R955 B B.n691 18.0485
R956 B.n633 B.n632 10.6151
R957 B.n632 B.n631 10.6151
R958 B.n631 B.n22 10.6151
R959 B.n627 B.n22 10.6151
R960 B.n627 B.n626 10.6151
R961 B.n626 B.n625 10.6151
R962 B.n625 B.n24 10.6151
R963 B.n621 B.n24 10.6151
R964 B.n621 B.n620 10.6151
R965 B.n620 B.n619 10.6151
R966 B.n619 B.n26 10.6151
R967 B.n615 B.n26 10.6151
R968 B.n615 B.n614 10.6151
R969 B.n614 B.n613 10.6151
R970 B.n613 B.n28 10.6151
R971 B.n609 B.n28 10.6151
R972 B.n609 B.n608 10.6151
R973 B.n608 B.n607 10.6151
R974 B.n607 B.n30 10.6151
R975 B.n603 B.n30 10.6151
R976 B.n603 B.n602 10.6151
R977 B.n602 B.n601 10.6151
R978 B.n601 B.n32 10.6151
R979 B.n597 B.n32 10.6151
R980 B.n597 B.n596 10.6151
R981 B.n596 B.n595 10.6151
R982 B.n595 B.n34 10.6151
R983 B.n591 B.n34 10.6151
R984 B.n591 B.n590 10.6151
R985 B.n590 B.n589 10.6151
R986 B.n589 B.n36 10.6151
R987 B.n585 B.n36 10.6151
R988 B.n585 B.n584 10.6151
R989 B.n584 B.n583 10.6151
R990 B.n583 B.n38 10.6151
R991 B.n579 B.n38 10.6151
R992 B.n579 B.n578 10.6151
R993 B.n578 B.n577 10.6151
R994 B.n577 B.n40 10.6151
R995 B.n573 B.n40 10.6151
R996 B.n573 B.n572 10.6151
R997 B.n572 B.n571 10.6151
R998 B.n568 B.n567 10.6151
R999 B.n567 B.n566 10.6151
R1000 B.n566 B.n46 10.6151
R1001 B.n562 B.n46 10.6151
R1002 B.n562 B.n561 10.6151
R1003 B.n561 B.n560 10.6151
R1004 B.n560 B.n48 10.6151
R1005 B.n556 B.n48 10.6151
R1006 B.n554 B.n553 10.6151
R1007 B.n553 B.n52 10.6151
R1008 B.n549 B.n52 10.6151
R1009 B.n549 B.n548 10.6151
R1010 B.n548 B.n547 10.6151
R1011 B.n547 B.n54 10.6151
R1012 B.n543 B.n54 10.6151
R1013 B.n543 B.n542 10.6151
R1014 B.n542 B.n541 10.6151
R1015 B.n541 B.n56 10.6151
R1016 B.n537 B.n56 10.6151
R1017 B.n537 B.n536 10.6151
R1018 B.n536 B.n535 10.6151
R1019 B.n535 B.n58 10.6151
R1020 B.n531 B.n58 10.6151
R1021 B.n531 B.n530 10.6151
R1022 B.n530 B.n529 10.6151
R1023 B.n529 B.n60 10.6151
R1024 B.n525 B.n60 10.6151
R1025 B.n525 B.n524 10.6151
R1026 B.n524 B.n523 10.6151
R1027 B.n523 B.n62 10.6151
R1028 B.n519 B.n62 10.6151
R1029 B.n519 B.n518 10.6151
R1030 B.n518 B.n517 10.6151
R1031 B.n517 B.n64 10.6151
R1032 B.n513 B.n64 10.6151
R1033 B.n513 B.n512 10.6151
R1034 B.n512 B.n511 10.6151
R1035 B.n511 B.n66 10.6151
R1036 B.n507 B.n66 10.6151
R1037 B.n507 B.n506 10.6151
R1038 B.n506 B.n505 10.6151
R1039 B.n505 B.n68 10.6151
R1040 B.n501 B.n68 10.6151
R1041 B.n501 B.n500 10.6151
R1042 B.n500 B.n499 10.6151
R1043 B.n499 B.n70 10.6151
R1044 B.n495 B.n70 10.6151
R1045 B.n495 B.n494 10.6151
R1046 B.n494 B.n493 10.6151
R1047 B.n493 B.n72 10.6151
R1048 B.n380 B.n379 10.6151
R1049 B.n381 B.n380 10.6151
R1050 B.n381 B.n108 10.6151
R1051 B.n385 B.n108 10.6151
R1052 B.n386 B.n385 10.6151
R1053 B.n387 B.n386 10.6151
R1054 B.n387 B.n106 10.6151
R1055 B.n391 B.n106 10.6151
R1056 B.n392 B.n391 10.6151
R1057 B.n393 B.n392 10.6151
R1058 B.n393 B.n104 10.6151
R1059 B.n397 B.n104 10.6151
R1060 B.n398 B.n397 10.6151
R1061 B.n399 B.n398 10.6151
R1062 B.n399 B.n102 10.6151
R1063 B.n403 B.n102 10.6151
R1064 B.n404 B.n403 10.6151
R1065 B.n405 B.n404 10.6151
R1066 B.n405 B.n100 10.6151
R1067 B.n409 B.n100 10.6151
R1068 B.n410 B.n409 10.6151
R1069 B.n411 B.n410 10.6151
R1070 B.n411 B.n98 10.6151
R1071 B.n415 B.n98 10.6151
R1072 B.n416 B.n415 10.6151
R1073 B.n417 B.n416 10.6151
R1074 B.n417 B.n96 10.6151
R1075 B.n421 B.n96 10.6151
R1076 B.n422 B.n421 10.6151
R1077 B.n423 B.n422 10.6151
R1078 B.n423 B.n94 10.6151
R1079 B.n427 B.n94 10.6151
R1080 B.n428 B.n427 10.6151
R1081 B.n429 B.n428 10.6151
R1082 B.n429 B.n92 10.6151
R1083 B.n433 B.n92 10.6151
R1084 B.n434 B.n433 10.6151
R1085 B.n435 B.n434 10.6151
R1086 B.n435 B.n90 10.6151
R1087 B.n439 B.n90 10.6151
R1088 B.n440 B.n439 10.6151
R1089 B.n441 B.n440 10.6151
R1090 B.n441 B.n88 10.6151
R1091 B.n445 B.n88 10.6151
R1092 B.n446 B.n445 10.6151
R1093 B.n447 B.n446 10.6151
R1094 B.n447 B.n86 10.6151
R1095 B.n451 B.n86 10.6151
R1096 B.n452 B.n451 10.6151
R1097 B.n453 B.n452 10.6151
R1098 B.n453 B.n84 10.6151
R1099 B.n457 B.n84 10.6151
R1100 B.n458 B.n457 10.6151
R1101 B.n459 B.n458 10.6151
R1102 B.n459 B.n82 10.6151
R1103 B.n463 B.n82 10.6151
R1104 B.n464 B.n463 10.6151
R1105 B.n465 B.n464 10.6151
R1106 B.n465 B.n80 10.6151
R1107 B.n469 B.n80 10.6151
R1108 B.n470 B.n469 10.6151
R1109 B.n471 B.n470 10.6151
R1110 B.n471 B.n78 10.6151
R1111 B.n475 B.n78 10.6151
R1112 B.n476 B.n475 10.6151
R1113 B.n477 B.n476 10.6151
R1114 B.n477 B.n76 10.6151
R1115 B.n481 B.n76 10.6151
R1116 B.n482 B.n481 10.6151
R1117 B.n483 B.n482 10.6151
R1118 B.n483 B.n74 10.6151
R1119 B.n487 B.n74 10.6151
R1120 B.n488 B.n487 10.6151
R1121 B.n489 B.n488 10.6151
R1122 B.n236 B.n235 10.6151
R1123 B.n237 B.n236 10.6151
R1124 B.n237 B.n160 10.6151
R1125 B.n241 B.n160 10.6151
R1126 B.n242 B.n241 10.6151
R1127 B.n243 B.n242 10.6151
R1128 B.n243 B.n158 10.6151
R1129 B.n247 B.n158 10.6151
R1130 B.n248 B.n247 10.6151
R1131 B.n249 B.n248 10.6151
R1132 B.n249 B.n156 10.6151
R1133 B.n253 B.n156 10.6151
R1134 B.n254 B.n253 10.6151
R1135 B.n255 B.n254 10.6151
R1136 B.n255 B.n154 10.6151
R1137 B.n259 B.n154 10.6151
R1138 B.n260 B.n259 10.6151
R1139 B.n261 B.n260 10.6151
R1140 B.n261 B.n152 10.6151
R1141 B.n265 B.n152 10.6151
R1142 B.n266 B.n265 10.6151
R1143 B.n267 B.n266 10.6151
R1144 B.n267 B.n150 10.6151
R1145 B.n271 B.n150 10.6151
R1146 B.n272 B.n271 10.6151
R1147 B.n273 B.n272 10.6151
R1148 B.n273 B.n148 10.6151
R1149 B.n277 B.n148 10.6151
R1150 B.n278 B.n277 10.6151
R1151 B.n279 B.n278 10.6151
R1152 B.n279 B.n146 10.6151
R1153 B.n283 B.n146 10.6151
R1154 B.n284 B.n283 10.6151
R1155 B.n285 B.n284 10.6151
R1156 B.n285 B.n144 10.6151
R1157 B.n289 B.n144 10.6151
R1158 B.n290 B.n289 10.6151
R1159 B.n291 B.n290 10.6151
R1160 B.n291 B.n142 10.6151
R1161 B.n295 B.n142 10.6151
R1162 B.n296 B.n295 10.6151
R1163 B.n297 B.n296 10.6151
R1164 B.n301 B.n300 10.6151
R1165 B.n302 B.n301 10.6151
R1166 B.n302 B.n136 10.6151
R1167 B.n306 B.n136 10.6151
R1168 B.n307 B.n306 10.6151
R1169 B.n308 B.n307 10.6151
R1170 B.n308 B.n134 10.6151
R1171 B.n312 B.n134 10.6151
R1172 B.n315 B.n314 10.6151
R1173 B.n315 B.n130 10.6151
R1174 B.n319 B.n130 10.6151
R1175 B.n320 B.n319 10.6151
R1176 B.n321 B.n320 10.6151
R1177 B.n321 B.n128 10.6151
R1178 B.n325 B.n128 10.6151
R1179 B.n326 B.n325 10.6151
R1180 B.n327 B.n326 10.6151
R1181 B.n327 B.n126 10.6151
R1182 B.n331 B.n126 10.6151
R1183 B.n332 B.n331 10.6151
R1184 B.n333 B.n332 10.6151
R1185 B.n333 B.n124 10.6151
R1186 B.n337 B.n124 10.6151
R1187 B.n338 B.n337 10.6151
R1188 B.n339 B.n338 10.6151
R1189 B.n339 B.n122 10.6151
R1190 B.n343 B.n122 10.6151
R1191 B.n344 B.n343 10.6151
R1192 B.n345 B.n344 10.6151
R1193 B.n345 B.n120 10.6151
R1194 B.n349 B.n120 10.6151
R1195 B.n350 B.n349 10.6151
R1196 B.n351 B.n350 10.6151
R1197 B.n351 B.n118 10.6151
R1198 B.n355 B.n118 10.6151
R1199 B.n356 B.n355 10.6151
R1200 B.n357 B.n356 10.6151
R1201 B.n357 B.n116 10.6151
R1202 B.n361 B.n116 10.6151
R1203 B.n362 B.n361 10.6151
R1204 B.n363 B.n362 10.6151
R1205 B.n363 B.n114 10.6151
R1206 B.n367 B.n114 10.6151
R1207 B.n368 B.n367 10.6151
R1208 B.n369 B.n368 10.6151
R1209 B.n369 B.n112 10.6151
R1210 B.n373 B.n112 10.6151
R1211 B.n374 B.n373 10.6151
R1212 B.n375 B.n374 10.6151
R1213 B.n375 B.n110 10.6151
R1214 B.n231 B.n162 10.6151
R1215 B.n231 B.n230 10.6151
R1216 B.n230 B.n229 10.6151
R1217 B.n229 B.n164 10.6151
R1218 B.n225 B.n164 10.6151
R1219 B.n225 B.n224 10.6151
R1220 B.n224 B.n223 10.6151
R1221 B.n223 B.n166 10.6151
R1222 B.n219 B.n166 10.6151
R1223 B.n219 B.n218 10.6151
R1224 B.n218 B.n217 10.6151
R1225 B.n217 B.n168 10.6151
R1226 B.n213 B.n168 10.6151
R1227 B.n213 B.n212 10.6151
R1228 B.n212 B.n211 10.6151
R1229 B.n211 B.n170 10.6151
R1230 B.n207 B.n170 10.6151
R1231 B.n207 B.n206 10.6151
R1232 B.n206 B.n205 10.6151
R1233 B.n205 B.n172 10.6151
R1234 B.n201 B.n172 10.6151
R1235 B.n201 B.n200 10.6151
R1236 B.n200 B.n199 10.6151
R1237 B.n199 B.n174 10.6151
R1238 B.n195 B.n174 10.6151
R1239 B.n195 B.n194 10.6151
R1240 B.n194 B.n193 10.6151
R1241 B.n193 B.n176 10.6151
R1242 B.n189 B.n176 10.6151
R1243 B.n189 B.n188 10.6151
R1244 B.n188 B.n187 10.6151
R1245 B.n187 B.n178 10.6151
R1246 B.n183 B.n178 10.6151
R1247 B.n183 B.n182 10.6151
R1248 B.n182 B.n181 10.6151
R1249 B.n181 B.n0 10.6151
R1250 B.n687 B.n1 10.6151
R1251 B.n687 B.n686 10.6151
R1252 B.n686 B.n685 10.6151
R1253 B.n685 B.n4 10.6151
R1254 B.n681 B.n4 10.6151
R1255 B.n681 B.n680 10.6151
R1256 B.n680 B.n679 10.6151
R1257 B.n679 B.n6 10.6151
R1258 B.n675 B.n6 10.6151
R1259 B.n675 B.n674 10.6151
R1260 B.n674 B.n673 10.6151
R1261 B.n673 B.n8 10.6151
R1262 B.n669 B.n8 10.6151
R1263 B.n669 B.n668 10.6151
R1264 B.n668 B.n667 10.6151
R1265 B.n667 B.n10 10.6151
R1266 B.n663 B.n10 10.6151
R1267 B.n663 B.n662 10.6151
R1268 B.n662 B.n661 10.6151
R1269 B.n661 B.n12 10.6151
R1270 B.n657 B.n12 10.6151
R1271 B.n657 B.n656 10.6151
R1272 B.n656 B.n655 10.6151
R1273 B.n655 B.n14 10.6151
R1274 B.n651 B.n14 10.6151
R1275 B.n651 B.n650 10.6151
R1276 B.n650 B.n649 10.6151
R1277 B.n649 B.n16 10.6151
R1278 B.n645 B.n16 10.6151
R1279 B.n645 B.n644 10.6151
R1280 B.n644 B.n643 10.6151
R1281 B.n643 B.n18 10.6151
R1282 B.n639 B.n18 10.6151
R1283 B.n639 B.n638 10.6151
R1284 B.n638 B.n637 10.6151
R1285 B.n637 B.n20 10.6151
R1286 B.n568 B.n44 6.5566
R1287 B.n556 B.n555 6.5566
R1288 B.n300 B.n140 6.5566
R1289 B.n313 B.n312 6.5566
R1290 B.n571 B.n44 4.05904
R1291 B.n555 B.n554 4.05904
R1292 B.n297 B.n140 4.05904
R1293 B.n314 B.n313 4.05904
R1294 B.n691 B.n0 2.81026
R1295 B.n691 B.n1 2.81026
C0 VTAIL VDD1 11.555099f
C1 VDD1 w_n2926_n3438# 2.31468f
C2 VP VTAIL 9.16237f
C3 VP w_n2926_n3438# 6.24928f
C4 VDD1 VDD2 1.3438f
C5 VTAIL B 3.17287f
C6 w_n2926_n3438# B 8.458631f
C7 VDD1 VN 0.150322f
C8 VP VDD2 0.417879f
C9 VDD2 B 2.05239f
C10 VTAIL w_n2926_n3438# 3.10871f
C11 VP VN 6.54783f
C12 VN B 0.956505f
C13 VTAIL VDD2 11.595f
C14 VDD2 w_n2926_n3438# 2.3907f
C15 VTAIL VN 9.147901f
C16 VN w_n2926_n3438# 5.87234f
C17 VN VDD2 9.058889f
C18 VP VDD1 9.32216f
C19 VDD1 B 1.98509f
C20 VP B 1.58318f
C21 VDD2 VSUBS 1.661248f
C22 VDD1 VSUBS 1.409556f
C23 VTAIL VSUBS 0.989577f
C24 VN VSUBS 5.67264f
C25 VP VSUBS 2.585701f
C26 B VSUBS 3.783522f
C27 w_n2926_n3438# VSUBS 0.12377p
C28 B.n0 VSUBS 0.005097f
C29 B.n1 VSUBS 0.005097f
C30 B.n2 VSUBS 0.008061f
C31 B.n3 VSUBS 0.008061f
C32 B.n4 VSUBS 0.008061f
C33 B.n5 VSUBS 0.008061f
C34 B.n6 VSUBS 0.008061f
C35 B.n7 VSUBS 0.008061f
C36 B.n8 VSUBS 0.008061f
C37 B.n9 VSUBS 0.008061f
C38 B.n10 VSUBS 0.008061f
C39 B.n11 VSUBS 0.008061f
C40 B.n12 VSUBS 0.008061f
C41 B.n13 VSUBS 0.008061f
C42 B.n14 VSUBS 0.008061f
C43 B.n15 VSUBS 0.008061f
C44 B.n16 VSUBS 0.008061f
C45 B.n17 VSUBS 0.008061f
C46 B.n18 VSUBS 0.008061f
C47 B.n19 VSUBS 0.008061f
C48 B.n20 VSUBS 0.017583f
C49 B.n21 VSUBS 0.008061f
C50 B.n22 VSUBS 0.008061f
C51 B.n23 VSUBS 0.008061f
C52 B.n24 VSUBS 0.008061f
C53 B.n25 VSUBS 0.008061f
C54 B.n26 VSUBS 0.008061f
C55 B.n27 VSUBS 0.008061f
C56 B.n28 VSUBS 0.008061f
C57 B.n29 VSUBS 0.008061f
C58 B.n30 VSUBS 0.008061f
C59 B.n31 VSUBS 0.008061f
C60 B.n32 VSUBS 0.008061f
C61 B.n33 VSUBS 0.008061f
C62 B.n34 VSUBS 0.008061f
C63 B.n35 VSUBS 0.008061f
C64 B.n36 VSUBS 0.008061f
C65 B.n37 VSUBS 0.008061f
C66 B.n38 VSUBS 0.008061f
C67 B.n39 VSUBS 0.008061f
C68 B.n40 VSUBS 0.008061f
C69 B.n41 VSUBS 0.008061f
C70 B.t11 VSUBS 0.46488f
C71 B.t10 VSUBS 0.479481f
C72 B.t9 VSUBS 0.797993f
C73 B.n42 VSUBS 0.202672f
C74 B.n43 VSUBS 0.076507f
C75 B.n44 VSUBS 0.018677f
C76 B.n45 VSUBS 0.008061f
C77 B.n46 VSUBS 0.008061f
C78 B.n47 VSUBS 0.008061f
C79 B.n48 VSUBS 0.008061f
C80 B.n49 VSUBS 0.008061f
C81 B.t8 VSUBS 0.464871f
C82 B.t7 VSUBS 0.479472f
C83 B.t6 VSUBS 0.797993f
C84 B.n50 VSUBS 0.202681f
C85 B.n51 VSUBS 0.076516f
C86 B.n52 VSUBS 0.008061f
C87 B.n53 VSUBS 0.008061f
C88 B.n54 VSUBS 0.008061f
C89 B.n55 VSUBS 0.008061f
C90 B.n56 VSUBS 0.008061f
C91 B.n57 VSUBS 0.008061f
C92 B.n58 VSUBS 0.008061f
C93 B.n59 VSUBS 0.008061f
C94 B.n60 VSUBS 0.008061f
C95 B.n61 VSUBS 0.008061f
C96 B.n62 VSUBS 0.008061f
C97 B.n63 VSUBS 0.008061f
C98 B.n64 VSUBS 0.008061f
C99 B.n65 VSUBS 0.008061f
C100 B.n66 VSUBS 0.008061f
C101 B.n67 VSUBS 0.008061f
C102 B.n68 VSUBS 0.008061f
C103 B.n69 VSUBS 0.008061f
C104 B.n70 VSUBS 0.008061f
C105 B.n71 VSUBS 0.008061f
C106 B.n72 VSUBS 0.017433f
C107 B.n73 VSUBS 0.008061f
C108 B.n74 VSUBS 0.008061f
C109 B.n75 VSUBS 0.008061f
C110 B.n76 VSUBS 0.008061f
C111 B.n77 VSUBS 0.008061f
C112 B.n78 VSUBS 0.008061f
C113 B.n79 VSUBS 0.008061f
C114 B.n80 VSUBS 0.008061f
C115 B.n81 VSUBS 0.008061f
C116 B.n82 VSUBS 0.008061f
C117 B.n83 VSUBS 0.008061f
C118 B.n84 VSUBS 0.008061f
C119 B.n85 VSUBS 0.008061f
C120 B.n86 VSUBS 0.008061f
C121 B.n87 VSUBS 0.008061f
C122 B.n88 VSUBS 0.008061f
C123 B.n89 VSUBS 0.008061f
C124 B.n90 VSUBS 0.008061f
C125 B.n91 VSUBS 0.008061f
C126 B.n92 VSUBS 0.008061f
C127 B.n93 VSUBS 0.008061f
C128 B.n94 VSUBS 0.008061f
C129 B.n95 VSUBS 0.008061f
C130 B.n96 VSUBS 0.008061f
C131 B.n97 VSUBS 0.008061f
C132 B.n98 VSUBS 0.008061f
C133 B.n99 VSUBS 0.008061f
C134 B.n100 VSUBS 0.008061f
C135 B.n101 VSUBS 0.008061f
C136 B.n102 VSUBS 0.008061f
C137 B.n103 VSUBS 0.008061f
C138 B.n104 VSUBS 0.008061f
C139 B.n105 VSUBS 0.008061f
C140 B.n106 VSUBS 0.008061f
C141 B.n107 VSUBS 0.008061f
C142 B.n108 VSUBS 0.008061f
C143 B.n109 VSUBS 0.008061f
C144 B.n110 VSUBS 0.018455f
C145 B.n111 VSUBS 0.008061f
C146 B.n112 VSUBS 0.008061f
C147 B.n113 VSUBS 0.008061f
C148 B.n114 VSUBS 0.008061f
C149 B.n115 VSUBS 0.008061f
C150 B.n116 VSUBS 0.008061f
C151 B.n117 VSUBS 0.008061f
C152 B.n118 VSUBS 0.008061f
C153 B.n119 VSUBS 0.008061f
C154 B.n120 VSUBS 0.008061f
C155 B.n121 VSUBS 0.008061f
C156 B.n122 VSUBS 0.008061f
C157 B.n123 VSUBS 0.008061f
C158 B.n124 VSUBS 0.008061f
C159 B.n125 VSUBS 0.008061f
C160 B.n126 VSUBS 0.008061f
C161 B.n127 VSUBS 0.008061f
C162 B.n128 VSUBS 0.008061f
C163 B.n129 VSUBS 0.008061f
C164 B.n130 VSUBS 0.008061f
C165 B.n131 VSUBS 0.008061f
C166 B.t1 VSUBS 0.464871f
C167 B.t2 VSUBS 0.479472f
C168 B.t0 VSUBS 0.797993f
C169 B.n132 VSUBS 0.202681f
C170 B.n133 VSUBS 0.076516f
C171 B.n134 VSUBS 0.008061f
C172 B.n135 VSUBS 0.008061f
C173 B.n136 VSUBS 0.008061f
C174 B.n137 VSUBS 0.008061f
C175 B.t4 VSUBS 0.46488f
C176 B.t5 VSUBS 0.479481f
C177 B.t3 VSUBS 0.797993f
C178 B.n138 VSUBS 0.202672f
C179 B.n139 VSUBS 0.076507f
C180 B.n140 VSUBS 0.018677f
C181 B.n141 VSUBS 0.008061f
C182 B.n142 VSUBS 0.008061f
C183 B.n143 VSUBS 0.008061f
C184 B.n144 VSUBS 0.008061f
C185 B.n145 VSUBS 0.008061f
C186 B.n146 VSUBS 0.008061f
C187 B.n147 VSUBS 0.008061f
C188 B.n148 VSUBS 0.008061f
C189 B.n149 VSUBS 0.008061f
C190 B.n150 VSUBS 0.008061f
C191 B.n151 VSUBS 0.008061f
C192 B.n152 VSUBS 0.008061f
C193 B.n153 VSUBS 0.008061f
C194 B.n154 VSUBS 0.008061f
C195 B.n155 VSUBS 0.008061f
C196 B.n156 VSUBS 0.008061f
C197 B.n157 VSUBS 0.008061f
C198 B.n158 VSUBS 0.008061f
C199 B.n159 VSUBS 0.008061f
C200 B.n160 VSUBS 0.008061f
C201 B.n161 VSUBS 0.008061f
C202 B.n162 VSUBS 0.017583f
C203 B.n163 VSUBS 0.008061f
C204 B.n164 VSUBS 0.008061f
C205 B.n165 VSUBS 0.008061f
C206 B.n166 VSUBS 0.008061f
C207 B.n167 VSUBS 0.008061f
C208 B.n168 VSUBS 0.008061f
C209 B.n169 VSUBS 0.008061f
C210 B.n170 VSUBS 0.008061f
C211 B.n171 VSUBS 0.008061f
C212 B.n172 VSUBS 0.008061f
C213 B.n173 VSUBS 0.008061f
C214 B.n174 VSUBS 0.008061f
C215 B.n175 VSUBS 0.008061f
C216 B.n176 VSUBS 0.008061f
C217 B.n177 VSUBS 0.008061f
C218 B.n178 VSUBS 0.008061f
C219 B.n179 VSUBS 0.008061f
C220 B.n180 VSUBS 0.008061f
C221 B.n181 VSUBS 0.008061f
C222 B.n182 VSUBS 0.008061f
C223 B.n183 VSUBS 0.008061f
C224 B.n184 VSUBS 0.008061f
C225 B.n185 VSUBS 0.008061f
C226 B.n186 VSUBS 0.008061f
C227 B.n187 VSUBS 0.008061f
C228 B.n188 VSUBS 0.008061f
C229 B.n189 VSUBS 0.008061f
C230 B.n190 VSUBS 0.008061f
C231 B.n191 VSUBS 0.008061f
C232 B.n192 VSUBS 0.008061f
C233 B.n193 VSUBS 0.008061f
C234 B.n194 VSUBS 0.008061f
C235 B.n195 VSUBS 0.008061f
C236 B.n196 VSUBS 0.008061f
C237 B.n197 VSUBS 0.008061f
C238 B.n198 VSUBS 0.008061f
C239 B.n199 VSUBS 0.008061f
C240 B.n200 VSUBS 0.008061f
C241 B.n201 VSUBS 0.008061f
C242 B.n202 VSUBS 0.008061f
C243 B.n203 VSUBS 0.008061f
C244 B.n204 VSUBS 0.008061f
C245 B.n205 VSUBS 0.008061f
C246 B.n206 VSUBS 0.008061f
C247 B.n207 VSUBS 0.008061f
C248 B.n208 VSUBS 0.008061f
C249 B.n209 VSUBS 0.008061f
C250 B.n210 VSUBS 0.008061f
C251 B.n211 VSUBS 0.008061f
C252 B.n212 VSUBS 0.008061f
C253 B.n213 VSUBS 0.008061f
C254 B.n214 VSUBS 0.008061f
C255 B.n215 VSUBS 0.008061f
C256 B.n216 VSUBS 0.008061f
C257 B.n217 VSUBS 0.008061f
C258 B.n218 VSUBS 0.008061f
C259 B.n219 VSUBS 0.008061f
C260 B.n220 VSUBS 0.008061f
C261 B.n221 VSUBS 0.008061f
C262 B.n222 VSUBS 0.008061f
C263 B.n223 VSUBS 0.008061f
C264 B.n224 VSUBS 0.008061f
C265 B.n225 VSUBS 0.008061f
C266 B.n226 VSUBS 0.008061f
C267 B.n227 VSUBS 0.008061f
C268 B.n228 VSUBS 0.008061f
C269 B.n229 VSUBS 0.008061f
C270 B.n230 VSUBS 0.008061f
C271 B.n231 VSUBS 0.008061f
C272 B.n232 VSUBS 0.008061f
C273 B.n233 VSUBS 0.017583f
C274 B.n234 VSUBS 0.018455f
C275 B.n235 VSUBS 0.018455f
C276 B.n236 VSUBS 0.008061f
C277 B.n237 VSUBS 0.008061f
C278 B.n238 VSUBS 0.008061f
C279 B.n239 VSUBS 0.008061f
C280 B.n240 VSUBS 0.008061f
C281 B.n241 VSUBS 0.008061f
C282 B.n242 VSUBS 0.008061f
C283 B.n243 VSUBS 0.008061f
C284 B.n244 VSUBS 0.008061f
C285 B.n245 VSUBS 0.008061f
C286 B.n246 VSUBS 0.008061f
C287 B.n247 VSUBS 0.008061f
C288 B.n248 VSUBS 0.008061f
C289 B.n249 VSUBS 0.008061f
C290 B.n250 VSUBS 0.008061f
C291 B.n251 VSUBS 0.008061f
C292 B.n252 VSUBS 0.008061f
C293 B.n253 VSUBS 0.008061f
C294 B.n254 VSUBS 0.008061f
C295 B.n255 VSUBS 0.008061f
C296 B.n256 VSUBS 0.008061f
C297 B.n257 VSUBS 0.008061f
C298 B.n258 VSUBS 0.008061f
C299 B.n259 VSUBS 0.008061f
C300 B.n260 VSUBS 0.008061f
C301 B.n261 VSUBS 0.008061f
C302 B.n262 VSUBS 0.008061f
C303 B.n263 VSUBS 0.008061f
C304 B.n264 VSUBS 0.008061f
C305 B.n265 VSUBS 0.008061f
C306 B.n266 VSUBS 0.008061f
C307 B.n267 VSUBS 0.008061f
C308 B.n268 VSUBS 0.008061f
C309 B.n269 VSUBS 0.008061f
C310 B.n270 VSUBS 0.008061f
C311 B.n271 VSUBS 0.008061f
C312 B.n272 VSUBS 0.008061f
C313 B.n273 VSUBS 0.008061f
C314 B.n274 VSUBS 0.008061f
C315 B.n275 VSUBS 0.008061f
C316 B.n276 VSUBS 0.008061f
C317 B.n277 VSUBS 0.008061f
C318 B.n278 VSUBS 0.008061f
C319 B.n279 VSUBS 0.008061f
C320 B.n280 VSUBS 0.008061f
C321 B.n281 VSUBS 0.008061f
C322 B.n282 VSUBS 0.008061f
C323 B.n283 VSUBS 0.008061f
C324 B.n284 VSUBS 0.008061f
C325 B.n285 VSUBS 0.008061f
C326 B.n286 VSUBS 0.008061f
C327 B.n287 VSUBS 0.008061f
C328 B.n288 VSUBS 0.008061f
C329 B.n289 VSUBS 0.008061f
C330 B.n290 VSUBS 0.008061f
C331 B.n291 VSUBS 0.008061f
C332 B.n292 VSUBS 0.008061f
C333 B.n293 VSUBS 0.008061f
C334 B.n294 VSUBS 0.008061f
C335 B.n295 VSUBS 0.008061f
C336 B.n296 VSUBS 0.008061f
C337 B.n297 VSUBS 0.005572f
C338 B.n298 VSUBS 0.008061f
C339 B.n299 VSUBS 0.008061f
C340 B.n300 VSUBS 0.00652f
C341 B.n301 VSUBS 0.008061f
C342 B.n302 VSUBS 0.008061f
C343 B.n303 VSUBS 0.008061f
C344 B.n304 VSUBS 0.008061f
C345 B.n305 VSUBS 0.008061f
C346 B.n306 VSUBS 0.008061f
C347 B.n307 VSUBS 0.008061f
C348 B.n308 VSUBS 0.008061f
C349 B.n309 VSUBS 0.008061f
C350 B.n310 VSUBS 0.008061f
C351 B.n311 VSUBS 0.008061f
C352 B.n312 VSUBS 0.00652f
C353 B.n313 VSUBS 0.018677f
C354 B.n314 VSUBS 0.005572f
C355 B.n315 VSUBS 0.008061f
C356 B.n316 VSUBS 0.008061f
C357 B.n317 VSUBS 0.008061f
C358 B.n318 VSUBS 0.008061f
C359 B.n319 VSUBS 0.008061f
C360 B.n320 VSUBS 0.008061f
C361 B.n321 VSUBS 0.008061f
C362 B.n322 VSUBS 0.008061f
C363 B.n323 VSUBS 0.008061f
C364 B.n324 VSUBS 0.008061f
C365 B.n325 VSUBS 0.008061f
C366 B.n326 VSUBS 0.008061f
C367 B.n327 VSUBS 0.008061f
C368 B.n328 VSUBS 0.008061f
C369 B.n329 VSUBS 0.008061f
C370 B.n330 VSUBS 0.008061f
C371 B.n331 VSUBS 0.008061f
C372 B.n332 VSUBS 0.008061f
C373 B.n333 VSUBS 0.008061f
C374 B.n334 VSUBS 0.008061f
C375 B.n335 VSUBS 0.008061f
C376 B.n336 VSUBS 0.008061f
C377 B.n337 VSUBS 0.008061f
C378 B.n338 VSUBS 0.008061f
C379 B.n339 VSUBS 0.008061f
C380 B.n340 VSUBS 0.008061f
C381 B.n341 VSUBS 0.008061f
C382 B.n342 VSUBS 0.008061f
C383 B.n343 VSUBS 0.008061f
C384 B.n344 VSUBS 0.008061f
C385 B.n345 VSUBS 0.008061f
C386 B.n346 VSUBS 0.008061f
C387 B.n347 VSUBS 0.008061f
C388 B.n348 VSUBS 0.008061f
C389 B.n349 VSUBS 0.008061f
C390 B.n350 VSUBS 0.008061f
C391 B.n351 VSUBS 0.008061f
C392 B.n352 VSUBS 0.008061f
C393 B.n353 VSUBS 0.008061f
C394 B.n354 VSUBS 0.008061f
C395 B.n355 VSUBS 0.008061f
C396 B.n356 VSUBS 0.008061f
C397 B.n357 VSUBS 0.008061f
C398 B.n358 VSUBS 0.008061f
C399 B.n359 VSUBS 0.008061f
C400 B.n360 VSUBS 0.008061f
C401 B.n361 VSUBS 0.008061f
C402 B.n362 VSUBS 0.008061f
C403 B.n363 VSUBS 0.008061f
C404 B.n364 VSUBS 0.008061f
C405 B.n365 VSUBS 0.008061f
C406 B.n366 VSUBS 0.008061f
C407 B.n367 VSUBS 0.008061f
C408 B.n368 VSUBS 0.008061f
C409 B.n369 VSUBS 0.008061f
C410 B.n370 VSUBS 0.008061f
C411 B.n371 VSUBS 0.008061f
C412 B.n372 VSUBS 0.008061f
C413 B.n373 VSUBS 0.008061f
C414 B.n374 VSUBS 0.008061f
C415 B.n375 VSUBS 0.008061f
C416 B.n376 VSUBS 0.008061f
C417 B.n377 VSUBS 0.018455f
C418 B.n378 VSUBS 0.017583f
C419 B.n379 VSUBS 0.017583f
C420 B.n380 VSUBS 0.008061f
C421 B.n381 VSUBS 0.008061f
C422 B.n382 VSUBS 0.008061f
C423 B.n383 VSUBS 0.008061f
C424 B.n384 VSUBS 0.008061f
C425 B.n385 VSUBS 0.008061f
C426 B.n386 VSUBS 0.008061f
C427 B.n387 VSUBS 0.008061f
C428 B.n388 VSUBS 0.008061f
C429 B.n389 VSUBS 0.008061f
C430 B.n390 VSUBS 0.008061f
C431 B.n391 VSUBS 0.008061f
C432 B.n392 VSUBS 0.008061f
C433 B.n393 VSUBS 0.008061f
C434 B.n394 VSUBS 0.008061f
C435 B.n395 VSUBS 0.008061f
C436 B.n396 VSUBS 0.008061f
C437 B.n397 VSUBS 0.008061f
C438 B.n398 VSUBS 0.008061f
C439 B.n399 VSUBS 0.008061f
C440 B.n400 VSUBS 0.008061f
C441 B.n401 VSUBS 0.008061f
C442 B.n402 VSUBS 0.008061f
C443 B.n403 VSUBS 0.008061f
C444 B.n404 VSUBS 0.008061f
C445 B.n405 VSUBS 0.008061f
C446 B.n406 VSUBS 0.008061f
C447 B.n407 VSUBS 0.008061f
C448 B.n408 VSUBS 0.008061f
C449 B.n409 VSUBS 0.008061f
C450 B.n410 VSUBS 0.008061f
C451 B.n411 VSUBS 0.008061f
C452 B.n412 VSUBS 0.008061f
C453 B.n413 VSUBS 0.008061f
C454 B.n414 VSUBS 0.008061f
C455 B.n415 VSUBS 0.008061f
C456 B.n416 VSUBS 0.008061f
C457 B.n417 VSUBS 0.008061f
C458 B.n418 VSUBS 0.008061f
C459 B.n419 VSUBS 0.008061f
C460 B.n420 VSUBS 0.008061f
C461 B.n421 VSUBS 0.008061f
C462 B.n422 VSUBS 0.008061f
C463 B.n423 VSUBS 0.008061f
C464 B.n424 VSUBS 0.008061f
C465 B.n425 VSUBS 0.008061f
C466 B.n426 VSUBS 0.008061f
C467 B.n427 VSUBS 0.008061f
C468 B.n428 VSUBS 0.008061f
C469 B.n429 VSUBS 0.008061f
C470 B.n430 VSUBS 0.008061f
C471 B.n431 VSUBS 0.008061f
C472 B.n432 VSUBS 0.008061f
C473 B.n433 VSUBS 0.008061f
C474 B.n434 VSUBS 0.008061f
C475 B.n435 VSUBS 0.008061f
C476 B.n436 VSUBS 0.008061f
C477 B.n437 VSUBS 0.008061f
C478 B.n438 VSUBS 0.008061f
C479 B.n439 VSUBS 0.008061f
C480 B.n440 VSUBS 0.008061f
C481 B.n441 VSUBS 0.008061f
C482 B.n442 VSUBS 0.008061f
C483 B.n443 VSUBS 0.008061f
C484 B.n444 VSUBS 0.008061f
C485 B.n445 VSUBS 0.008061f
C486 B.n446 VSUBS 0.008061f
C487 B.n447 VSUBS 0.008061f
C488 B.n448 VSUBS 0.008061f
C489 B.n449 VSUBS 0.008061f
C490 B.n450 VSUBS 0.008061f
C491 B.n451 VSUBS 0.008061f
C492 B.n452 VSUBS 0.008061f
C493 B.n453 VSUBS 0.008061f
C494 B.n454 VSUBS 0.008061f
C495 B.n455 VSUBS 0.008061f
C496 B.n456 VSUBS 0.008061f
C497 B.n457 VSUBS 0.008061f
C498 B.n458 VSUBS 0.008061f
C499 B.n459 VSUBS 0.008061f
C500 B.n460 VSUBS 0.008061f
C501 B.n461 VSUBS 0.008061f
C502 B.n462 VSUBS 0.008061f
C503 B.n463 VSUBS 0.008061f
C504 B.n464 VSUBS 0.008061f
C505 B.n465 VSUBS 0.008061f
C506 B.n466 VSUBS 0.008061f
C507 B.n467 VSUBS 0.008061f
C508 B.n468 VSUBS 0.008061f
C509 B.n469 VSUBS 0.008061f
C510 B.n470 VSUBS 0.008061f
C511 B.n471 VSUBS 0.008061f
C512 B.n472 VSUBS 0.008061f
C513 B.n473 VSUBS 0.008061f
C514 B.n474 VSUBS 0.008061f
C515 B.n475 VSUBS 0.008061f
C516 B.n476 VSUBS 0.008061f
C517 B.n477 VSUBS 0.008061f
C518 B.n478 VSUBS 0.008061f
C519 B.n479 VSUBS 0.008061f
C520 B.n480 VSUBS 0.008061f
C521 B.n481 VSUBS 0.008061f
C522 B.n482 VSUBS 0.008061f
C523 B.n483 VSUBS 0.008061f
C524 B.n484 VSUBS 0.008061f
C525 B.n485 VSUBS 0.008061f
C526 B.n486 VSUBS 0.008061f
C527 B.n487 VSUBS 0.008061f
C528 B.n488 VSUBS 0.008061f
C529 B.n489 VSUBS 0.018605f
C530 B.n490 VSUBS 0.017583f
C531 B.n491 VSUBS 0.018455f
C532 B.n492 VSUBS 0.008061f
C533 B.n493 VSUBS 0.008061f
C534 B.n494 VSUBS 0.008061f
C535 B.n495 VSUBS 0.008061f
C536 B.n496 VSUBS 0.008061f
C537 B.n497 VSUBS 0.008061f
C538 B.n498 VSUBS 0.008061f
C539 B.n499 VSUBS 0.008061f
C540 B.n500 VSUBS 0.008061f
C541 B.n501 VSUBS 0.008061f
C542 B.n502 VSUBS 0.008061f
C543 B.n503 VSUBS 0.008061f
C544 B.n504 VSUBS 0.008061f
C545 B.n505 VSUBS 0.008061f
C546 B.n506 VSUBS 0.008061f
C547 B.n507 VSUBS 0.008061f
C548 B.n508 VSUBS 0.008061f
C549 B.n509 VSUBS 0.008061f
C550 B.n510 VSUBS 0.008061f
C551 B.n511 VSUBS 0.008061f
C552 B.n512 VSUBS 0.008061f
C553 B.n513 VSUBS 0.008061f
C554 B.n514 VSUBS 0.008061f
C555 B.n515 VSUBS 0.008061f
C556 B.n516 VSUBS 0.008061f
C557 B.n517 VSUBS 0.008061f
C558 B.n518 VSUBS 0.008061f
C559 B.n519 VSUBS 0.008061f
C560 B.n520 VSUBS 0.008061f
C561 B.n521 VSUBS 0.008061f
C562 B.n522 VSUBS 0.008061f
C563 B.n523 VSUBS 0.008061f
C564 B.n524 VSUBS 0.008061f
C565 B.n525 VSUBS 0.008061f
C566 B.n526 VSUBS 0.008061f
C567 B.n527 VSUBS 0.008061f
C568 B.n528 VSUBS 0.008061f
C569 B.n529 VSUBS 0.008061f
C570 B.n530 VSUBS 0.008061f
C571 B.n531 VSUBS 0.008061f
C572 B.n532 VSUBS 0.008061f
C573 B.n533 VSUBS 0.008061f
C574 B.n534 VSUBS 0.008061f
C575 B.n535 VSUBS 0.008061f
C576 B.n536 VSUBS 0.008061f
C577 B.n537 VSUBS 0.008061f
C578 B.n538 VSUBS 0.008061f
C579 B.n539 VSUBS 0.008061f
C580 B.n540 VSUBS 0.008061f
C581 B.n541 VSUBS 0.008061f
C582 B.n542 VSUBS 0.008061f
C583 B.n543 VSUBS 0.008061f
C584 B.n544 VSUBS 0.008061f
C585 B.n545 VSUBS 0.008061f
C586 B.n546 VSUBS 0.008061f
C587 B.n547 VSUBS 0.008061f
C588 B.n548 VSUBS 0.008061f
C589 B.n549 VSUBS 0.008061f
C590 B.n550 VSUBS 0.008061f
C591 B.n551 VSUBS 0.008061f
C592 B.n552 VSUBS 0.008061f
C593 B.n553 VSUBS 0.008061f
C594 B.n554 VSUBS 0.005572f
C595 B.n555 VSUBS 0.018677f
C596 B.n556 VSUBS 0.00652f
C597 B.n557 VSUBS 0.008061f
C598 B.n558 VSUBS 0.008061f
C599 B.n559 VSUBS 0.008061f
C600 B.n560 VSUBS 0.008061f
C601 B.n561 VSUBS 0.008061f
C602 B.n562 VSUBS 0.008061f
C603 B.n563 VSUBS 0.008061f
C604 B.n564 VSUBS 0.008061f
C605 B.n565 VSUBS 0.008061f
C606 B.n566 VSUBS 0.008061f
C607 B.n567 VSUBS 0.008061f
C608 B.n568 VSUBS 0.00652f
C609 B.n569 VSUBS 0.008061f
C610 B.n570 VSUBS 0.008061f
C611 B.n571 VSUBS 0.005572f
C612 B.n572 VSUBS 0.008061f
C613 B.n573 VSUBS 0.008061f
C614 B.n574 VSUBS 0.008061f
C615 B.n575 VSUBS 0.008061f
C616 B.n576 VSUBS 0.008061f
C617 B.n577 VSUBS 0.008061f
C618 B.n578 VSUBS 0.008061f
C619 B.n579 VSUBS 0.008061f
C620 B.n580 VSUBS 0.008061f
C621 B.n581 VSUBS 0.008061f
C622 B.n582 VSUBS 0.008061f
C623 B.n583 VSUBS 0.008061f
C624 B.n584 VSUBS 0.008061f
C625 B.n585 VSUBS 0.008061f
C626 B.n586 VSUBS 0.008061f
C627 B.n587 VSUBS 0.008061f
C628 B.n588 VSUBS 0.008061f
C629 B.n589 VSUBS 0.008061f
C630 B.n590 VSUBS 0.008061f
C631 B.n591 VSUBS 0.008061f
C632 B.n592 VSUBS 0.008061f
C633 B.n593 VSUBS 0.008061f
C634 B.n594 VSUBS 0.008061f
C635 B.n595 VSUBS 0.008061f
C636 B.n596 VSUBS 0.008061f
C637 B.n597 VSUBS 0.008061f
C638 B.n598 VSUBS 0.008061f
C639 B.n599 VSUBS 0.008061f
C640 B.n600 VSUBS 0.008061f
C641 B.n601 VSUBS 0.008061f
C642 B.n602 VSUBS 0.008061f
C643 B.n603 VSUBS 0.008061f
C644 B.n604 VSUBS 0.008061f
C645 B.n605 VSUBS 0.008061f
C646 B.n606 VSUBS 0.008061f
C647 B.n607 VSUBS 0.008061f
C648 B.n608 VSUBS 0.008061f
C649 B.n609 VSUBS 0.008061f
C650 B.n610 VSUBS 0.008061f
C651 B.n611 VSUBS 0.008061f
C652 B.n612 VSUBS 0.008061f
C653 B.n613 VSUBS 0.008061f
C654 B.n614 VSUBS 0.008061f
C655 B.n615 VSUBS 0.008061f
C656 B.n616 VSUBS 0.008061f
C657 B.n617 VSUBS 0.008061f
C658 B.n618 VSUBS 0.008061f
C659 B.n619 VSUBS 0.008061f
C660 B.n620 VSUBS 0.008061f
C661 B.n621 VSUBS 0.008061f
C662 B.n622 VSUBS 0.008061f
C663 B.n623 VSUBS 0.008061f
C664 B.n624 VSUBS 0.008061f
C665 B.n625 VSUBS 0.008061f
C666 B.n626 VSUBS 0.008061f
C667 B.n627 VSUBS 0.008061f
C668 B.n628 VSUBS 0.008061f
C669 B.n629 VSUBS 0.008061f
C670 B.n630 VSUBS 0.008061f
C671 B.n631 VSUBS 0.008061f
C672 B.n632 VSUBS 0.008061f
C673 B.n633 VSUBS 0.018455f
C674 B.n634 VSUBS 0.018455f
C675 B.n635 VSUBS 0.017583f
C676 B.n636 VSUBS 0.008061f
C677 B.n637 VSUBS 0.008061f
C678 B.n638 VSUBS 0.008061f
C679 B.n639 VSUBS 0.008061f
C680 B.n640 VSUBS 0.008061f
C681 B.n641 VSUBS 0.008061f
C682 B.n642 VSUBS 0.008061f
C683 B.n643 VSUBS 0.008061f
C684 B.n644 VSUBS 0.008061f
C685 B.n645 VSUBS 0.008061f
C686 B.n646 VSUBS 0.008061f
C687 B.n647 VSUBS 0.008061f
C688 B.n648 VSUBS 0.008061f
C689 B.n649 VSUBS 0.008061f
C690 B.n650 VSUBS 0.008061f
C691 B.n651 VSUBS 0.008061f
C692 B.n652 VSUBS 0.008061f
C693 B.n653 VSUBS 0.008061f
C694 B.n654 VSUBS 0.008061f
C695 B.n655 VSUBS 0.008061f
C696 B.n656 VSUBS 0.008061f
C697 B.n657 VSUBS 0.008061f
C698 B.n658 VSUBS 0.008061f
C699 B.n659 VSUBS 0.008061f
C700 B.n660 VSUBS 0.008061f
C701 B.n661 VSUBS 0.008061f
C702 B.n662 VSUBS 0.008061f
C703 B.n663 VSUBS 0.008061f
C704 B.n664 VSUBS 0.008061f
C705 B.n665 VSUBS 0.008061f
C706 B.n666 VSUBS 0.008061f
C707 B.n667 VSUBS 0.008061f
C708 B.n668 VSUBS 0.008061f
C709 B.n669 VSUBS 0.008061f
C710 B.n670 VSUBS 0.008061f
C711 B.n671 VSUBS 0.008061f
C712 B.n672 VSUBS 0.008061f
C713 B.n673 VSUBS 0.008061f
C714 B.n674 VSUBS 0.008061f
C715 B.n675 VSUBS 0.008061f
C716 B.n676 VSUBS 0.008061f
C717 B.n677 VSUBS 0.008061f
C718 B.n678 VSUBS 0.008061f
C719 B.n679 VSUBS 0.008061f
C720 B.n680 VSUBS 0.008061f
C721 B.n681 VSUBS 0.008061f
C722 B.n682 VSUBS 0.008061f
C723 B.n683 VSUBS 0.008061f
C724 B.n684 VSUBS 0.008061f
C725 B.n685 VSUBS 0.008061f
C726 B.n686 VSUBS 0.008061f
C727 B.n687 VSUBS 0.008061f
C728 B.n688 VSUBS 0.008061f
C729 B.n689 VSUBS 0.008061f
C730 B.n690 VSUBS 0.008061f
C731 B.n691 VSUBS 0.018253f
C732 VDD2.t8 VSUBS 2.81178f
C733 VDD2.t2 VSUBS 0.270399f
C734 VDD2.t0 VSUBS 0.270399f
C735 VDD2.n0 VSUBS 2.14785f
C736 VDD2.n1 VSUBS 1.35525f
C737 VDD2.t7 VSUBS 0.270399f
C738 VDD2.t1 VSUBS 0.270399f
C739 VDD2.n2 VSUBS 2.15704f
C740 VDD2.n3 VSUBS 2.75209f
C741 VDD2.t6 VSUBS 2.79941f
C742 VDD2.n4 VSUBS 3.21364f
C743 VDD2.t4 VSUBS 0.270399f
C744 VDD2.t3 VSUBS 0.270399f
C745 VDD2.n5 VSUBS 2.14786f
C746 VDD2.n6 VSUBS 0.657539f
C747 VDD2.t9 VSUBS 0.270399f
C748 VDD2.t5 VSUBS 0.270399f
C749 VDD2.n7 VSUBS 2.157f
C750 VN.n0 VSUBS 0.039918f
C751 VN.t8 VSUBS 1.7476f
C752 VN.n1 VSUBS 0.066903f
C753 VN.n2 VSUBS 0.039918f
C754 VN.t9 VSUBS 1.7476f
C755 VN.n3 VSUBS 0.67309f
C756 VN.n4 VSUBS 0.039918f
C757 VN.t7 VSUBS 1.7476f
C758 VN.n5 VSUBS 0.691623f
C759 VN.t1 VSUBS 1.83493f
C760 VN.n6 VSUBS 0.731146f
C761 VN.n7 VSUBS 0.210793f
C762 VN.n8 VSUBS 0.047217f
C763 VN.n9 VSUBS 0.051047f
C764 VN.n10 VSUBS 0.065508f
C765 VN.n11 VSUBS 0.039918f
C766 VN.n12 VSUBS 0.039918f
C767 VN.n13 VSUBS 0.039918f
C768 VN.n14 VSUBS 0.065508f
C769 VN.n15 VSUBS 0.051047f
C770 VN.t2 VSUBS 1.7476f
C771 VN.n16 VSUBS 0.635423f
C772 VN.n17 VSUBS 0.047217f
C773 VN.n18 VSUBS 0.039918f
C774 VN.n19 VSUBS 0.039918f
C775 VN.n20 VSUBS 0.039918f
C776 VN.n21 VSUBS 0.03385f
C777 VN.n22 VSUBS 0.063019f
C778 VN.n23 VSUBS 0.70888f
C779 VN.n24 VSUBS 0.036284f
C780 VN.n25 VSUBS 0.039918f
C781 VN.t3 VSUBS 1.7476f
C782 VN.n26 VSUBS 0.066903f
C783 VN.n27 VSUBS 0.039918f
C784 VN.t5 VSUBS 1.7476f
C785 VN.n28 VSUBS 0.635423f
C786 VN.t6 VSUBS 1.7476f
C787 VN.n29 VSUBS 0.67309f
C788 VN.n30 VSUBS 0.039918f
C789 VN.t0 VSUBS 1.7476f
C790 VN.n31 VSUBS 0.691623f
C791 VN.t4 VSUBS 1.83493f
C792 VN.n32 VSUBS 0.731146f
C793 VN.n33 VSUBS 0.210793f
C794 VN.n34 VSUBS 0.047217f
C795 VN.n35 VSUBS 0.051047f
C796 VN.n36 VSUBS 0.065508f
C797 VN.n37 VSUBS 0.039918f
C798 VN.n38 VSUBS 0.039918f
C799 VN.n39 VSUBS 0.039918f
C800 VN.n40 VSUBS 0.065508f
C801 VN.n41 VSUBS 0.051047f
C802 VN.n42 VSUBS 0.047217f
C803 VN.n43 VSUBS 0.039918f
C804 VN.n44 VSUBS 0.039918f
C805 VN.n45 VSUBS 0.039918f
C806 VN.n46 VSUBS 0.03385f
C807 VN.n47 VSUBS 0.063019f
C808 VN.n48 VSUBS 0.70888f
C809 VN.n49 VSUBS 1.95562f
C810 VTAIL.t4 VSUBS 0.274821f
C811 VTAIL.t5 VSUBS 0.274821f
C812 VTAIL.n0 VSUBS 2.04629f
C813 VTAIL.n1 VSUBS 0.809332f
C814 VTAIL.t15 VSUBS 2.69121f
C815 VTAIL.n2 VSUBS 0.940518f
C816 VTAIL.t9 VSUBS 0.274821f
C817 VTAIL.t10 VSUBS 0.274821f
C818 VTAIL.n3 VSUBS 2.04629f
C819 VTAIL.n4 VSUBS 0.857047f
C820 VTAIL.t11 VSUBS 0.274821f
C821 VTAIL.t16 VSUBS 0.274821f
C822 VTAIL.n5 VSUBS 2.04629f
C823 VTAIL.n6 VSUBS 2.3331f
C824 VTAIL.t3 VSUBS 0.274821f
C825 VTAIL.t0 VSUBS 0.274821f
C826 VTAIL.n7 VSUBS 2.0463f
C827 VTAIL.n8 VSUBS 2.33309f
C828 VTAIL.t19 VSUBS 0.274821f
C829 VTAIL.t2 VSUBS 0.274821f
C830 VTAIL.n9 VSUBS 2.0463f
C831 VTAIL.n10 VSUBS 0.857039f
C832 VTAIL.t8 VSUBS 2.69122f
C833 VTAIL.n11 VSUBS 0.940515f
C834 VTAIL.t13 VSUBS 0.274821f
C835 VTAIL.t18 VSUBS 0.274821f
C836 VTAIL.n12 VSUBS 2.0463f
C837 VTAIL.n13 VSUBS 0.835919f
C838 VTAIL.t12 VSUBS 0.274821f
C839 VTAIL.t14 VSUBS 0.274821f
C840 VTAIL.n14 VSUBS 2.0463f
C841 VTAIL.n15 VSUBS 0.857039f
C842 VTAIL.t17 VSUBS 2.69121f
C843 VTAIL.n16 VSUBS 2.3102f
C844 VTAIL.t7 VSUBS 2.69121f
C845 VTAIL.n17 VSUBS 2.31019f
C846 VTAIL.t6 VSUBS 0.274821f
C847 VTAIL.t1 VSUBS 0.274821f
C848 VTAIL.n18 VSUBS 2.04629f
C849 VTAIL.n19 VSUBS 0.756141f
C850 VDD1.t0 VSUBS 2.57816f
C851 VDD1.t5 VSUBS 0.247932f
C852 VDD1.t6 VSUBS 0.247932f
C853 VDD1.n0 VSUBS 1.9694f
C854 VDD1.n1 VSUBS 1.24994f
C855 VDD1.t4 VSUBS 2.57816f
C856 VDD1.t2 VSUBS 0.247932f
C857 VDD1.t1 VSUBS 0.247932f
C858 VDD1.n2 VSUBS 1.96939f
C859 VDD1.n3 VSUBS 1.24265f
C860 VDD1.t3 VSUBS 0.247932f
C861 VDD1.t7 VSUBS 0.247932f
C862 VDD1.n4 VSUBS 1.97781f
C863 VDD1.n5 VSUBS 2.61652f
C864 VDD1.t9 VSUBS 0.247932f
C865 VDD1.t8 VSUBS 0.247932f
C866 VDD1.n6 VSUBS 1.96939f
C867 VDD1.n7 VSUBS 2.9501f
C868 VP.n0 VSUBS 0.040776f
C869 VP.t3 VSUBS 1.78514f
C870 VP.n1 VSUBS 0.06834f
C871 VP.n2 VSUBS 0.040776f
C872 VP.t9 VSUBS 1.78514f
C873 VP.n3 VSUBS 0.687549f
C874 VP.n4 VSUBS 0.040776f
C875 VP.t2 VSUBS 1.78514f
C876 VP.n5 VSUBS 0.649072f
C877 VP.n6 VSUBS 0.040776f
C878 VP.t7 VSUBS 1.78514f
C879 VP.n7 VSUBS 0.724107f
C880 VP.n8 VSUBS 0.040776f
C881 VP.t1 VSUBS 1.78514f
C882 VP.n9 VSUBS 0.06834f
C883 VP.n10 VSUBS 0.040776f
C884 VP.t6 VSUBS 1.78514f
C885 VP.n11 VSUBS 0.687549f
C886 VP.n12 VSUBS 0.040776f
C887 VP.t0 VSUBS 1.78514f
C888 VP.n13 VSUBS 0.70648f
C889 VP.t5 VSUBS 1.87434f
C890 VP.n14 VSUBS 0.746852f
C891 VP.n15 VSUBS 0.215321f
C892 VP.n16 VSUBS 0.048231f
C893 VP.n17 VSUBS 0.052144f
C894 VP.n18 VSUBS 0.066915f
C895 VP.n19 VSUBS 0.040776f
C896 VP.n20 VSUBS 0.040776f
C897 VP.n21 VSUBS 0.040776f
C898 VP.n22 VSUBS 0.066915f
C899 VP.n23 VSUBS 0.052144f
C900 VP.t4 VSUBS 1.78514f
C901 VP.n24 VSUBS 0.649072f
C902 VP.n25 VSUBS 0.048231f
C903 VP.n26 VSUBS 0.040776f
C904 VP.n27 VSUBS 0.040776f
C905 VP.n28 VSUBS 0.040776f
C906 VP.n29 VSUBS 0.034577f
C907 VP.n30 VSUBS 0.064373f
C908 VP.n31 VSUBS 0.724107f
C909 VP.n32 VSUBS 1.97101f
C910 VP.n33 VSUBS 2.00272f
C911 VP.n34 VSUBS 0.040776f
C912 VP.n35 VSUBS 0.064373f
C913 VP.n36 VSUBS 0.034577f
C914 VP.n37 VSUBS 0.06834f
C915 VP.n38 VSUBS 0.040776f
C916 VP.n39 VSUBS 0.040776f
C917 VP.n40 VSUBS 0.048231f
C918 VP.n41 VSUBS 0.052144f
C919 VP.n42 VSUBS 0.066915f
C920 VP.n43 VSUBS 0.040776f
C921 VP.n44 VSUBS 0.040776f
C922 VP.n45 VSUBS 0.040776f
C923 VP.n46 VSUBS 0.066915f
C924 VP.n47 VSUBS 0.052144f
C925 VP.t8 VSUBS 1.78514f
C926 VP.n48 VSUBS 0.649072f
C927 VP.n49 VSUBS 0.048231f
C928 VP.n50 VSUBS 0.040776f
C929 VP.n51 VSUBS 0.040776f
C930 VP.n52 VSUBS 0.040776f
C931 VP.n53 VSUBS 0.034577f
C932 VP.n54 VSUBS 0.064373f
C933 VP.n55 VSUBS 0.724107f
C934 VP.n56 VSUBS 0.037063f
.ends

