* NGSPICE file created from diff_pair_sample_1417.ext - technology: sky130A

.subckt diff_pair_sample_1417 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t7 VN.t0 VTAIL.t12 B.t6 sky130_fd_pr__nfet_01v8 ad=2.63505 pd=16.3 as=2.63505 ps=16.3 w=15.97 l=1.37
X1 B.t21 B.t19 B.t20 B.t9 sky130_fd_pr__nfet_01v8 ad=6.2283 pd=32.72 as=0 ps=0 w=15.97 l=1.37
X2 VTAIL.t4 VP.t0 VDD1.t7 B.t4 sky130_fd_pr__nfet_01v8 ad=6.2283 pd=32.72 as=2.63505 ps=16.3 w=15.97 l=1.37
X3 B.t18 B.t16 B.t17 B.t13 sky130_fd_pr__nfet_01v8 ad=6.2283 pd=32.72 as=0 ps=0 w=15.97 l=1.37
X4 VTAIL.t5 VP.t1 VDD1.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=2.63505 pd=16.3 as=2.63505 ps=16.3 w=15.97 l=1.37
X5 VDD1.t5 VP.t2 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.63505 pd=16.3 as=2.63505 ps=16.3 w=15.97 l=1.37
X6 VTAIL.t2 VP.t3 VDD1.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=2.63505 pd=16.3 as=2.63505 ps=16.3 w=15.97 l=1.37
X7 VTAIL.t10 VN.t1 VDD2.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=6.2283 pd=32.72 as=2.63505 ps=16.3 w=15.97 l=1.37
X8 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=6.2283 pd=32.72 as=0 ps=0 w=15.97 l=1.37
X9 VDD1.t3 VP.t4 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=2.63505 pd=16.3 as=2.63505 ps=16.3 w=15.97 l=1.37
X10 VDD1.t2 VP.t5 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=2.63505 pd=16.3 as=6.2283 ps=32.72 w=15.97 l=1.37
X11 VTAIL.t15 VN.t2 VDD2.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.63505 pd=16.3 as=2.63505 ps=16.3 w=15.97 l=1.37
X12 VDD1.t1 VP.t6 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.63505 pd=16.3 as=6.2283 ps=32.72 w=15.97 l=1.37
X13 VDD2.t4 VN.t3 VTAIL.t8 B.t1 sky130_fd_pr__nfet_01v8 ad=2.63505 pd=16.3 as=6.2283 ps=32.72 w=15.97 l=1.37
X14 VDD2.t3 VN.t4 VTAIL.t9 B.t7 sky130_fd_pr__nfet_01v8 ad=2.63505 pd=16.3 as=6.2283 ps=32.72 w=15.97 l=1.37
X15 VTAIL.t11 VN.t5 VDD2.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.63505 pd=16.3 as=2.63505 ps=16.3 w=15.97 l=1.37
X16 VDD2.t1 VN.t6 VTAIL.t14 B.t3 sky130_fd_pr__nfet_01v8 ad=2.63505 pd=16.3 as=2.63505 ps=16.3 w=15.97 l=1.37
X17 VTAIL.t0 VP.t7 VDD1.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=6.2283 pd=32.72 as=2.63505 ps=16.3 w=15.97 l=1.37
X18 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=6.2283 pd=32.72 as=0 ps=0 w=15.97 l=1.37
X19 VTAIL.t13 VN.t7 VDD2.t0 B.t4 sky130_fd_pr__nfet_01v8 ad=6.2283 pd=32.72 as=2.63505 ps=16.3 w=15.97 l=1.37
R0 VN.n5 VN.t7 311.577
R1 VN.n25 VN.t4 311.577
R2 VN.n4 VN.t6 280.933
R3 VN.n10 VN.t2 280.933
R4 VN.n17 VN.t3 280.933
R5 VN.n24 VN.t5 280.933
R6 VN.n22 VN.t0 280.933
R7 VN.n36 VN.t1 280.933
R8 VN.n18 VN.n17 171.088
R9 VN.n37 VN.n36 171.088
R10 VN.n35 VN.n19 161.3
R11 VN.n34 VN.n33 161.3
R12 VN.n32 VN.n20 161.3
R13 VN.n31 VN.n30 161.3
R14 VN.n29 VN.n21 161.3
R15 VN.n28 VN.n27 161.3
R16 VN.n26 VN.n23 161.3
R17 VN.n16 VN.n0 161.3
R18 VN.n15 VN.n14 161.3
R19 VN.n13 VN.n1 161.3
R20 VN.n12 VN.n11 161.3
R21 VN.n9 VN.n2 161.3
R22 VN.n8 VN.n7 161.3
R23 VN.n6 VN.n3 161.3
R24 VN.n5 VN.n4 60.1408
R25 VN.n25 VN.n24 60.1408
R26 VN.n9 VN.n8 56.5193
R27 VN.n29 VN.n28 56.5193
R28 VN VN.n37 48.4948
R29 VN.n15 VN.n1 45.3497
R30 VN.n34 VN.n20 45.3497
R31 VN.n16 VN.n15 35.6371
R32 VN.n35 VN.n34 35.6371
R33 VN.n26 VN.n25 26.7826
R34 VN.n6 VN.n5 26.7826
R35 VN.n8 VN.n3 24.4675
R36 VN.n11 VN.n9 24.4675
R37 VN.n28 VN.n23 24.4675
R38 VN.n30 VN.n29 24.4675
R39 VN.n10 VN.n1 19.5741
R40 VN.n22 VN.n20 19.5741
R41 VN.n17 VN.n16 14.6807
R42 VN.n36 VN.n35 14.6807
R43 VN.n4 VN.n3 4.8939
R44 VN.n11 VN.n10 4.8939
R45 VN.n24 VN.n23 4.8939
R46 VN.n30 VN.n22 4.8939
R47 VN.n37 VN.n19 0.189894
R48 VN.n33 VN.n19 0.189894
R49 VN.n33 VN.n32 0.189894
R50 VN.n32 VN.n31 0.189894
R51 VN.n31 VN.n21 0.189894
R52 VN.n27 VN.n21 0.189894
R53 VN.n27 VN.n26 0.189894
R54 VN.n7 VN.n6 0.189894
R55 VN.n7 VN.n2 0.189894
R56 VN.n12 VN.n2 0.189894
R57 VN.n13 VN.n12 0.189894
R58 VN.n14 VN.n13 0.189894
R59 VN.n14 VN.n0 0.189894
R60 VN.n18 VN.n0 0.189894
R61 VN VN.n18 0.0516364
R62 VTAIL.n11 VTAIL.t4 43.6195
R63 VTAIL.n10 VTAIL.t9 43.6195
R64 VTAIL.n7 VTAIL.t10 43.6195
R65 VTAIL.n14 VTAIL.t1 43.6195
R66 VTAIL.n15 VTAIL.t8 43.6193
R67 VTAIL.n2 VTAIL.t13 43.6193
R68 VTAIL.n3 VTAIL.t7 43.6193
R69 VTAIL.n6 VTAIL.t0 43.6193
R70 VTAIL.n13 VTAIL.n12 42.3797
R71 VTAIL.n9 VTAIL.n8 42.3797
R72 VTAIL.n1 VTAIL.n0 42.3795
R73 VTAIL.n5 VTAIL.n4 42.3795
R74 VTAIL.n15 VTAIL.n14 27.5996
R75 VTAIL.n7 VTAIL.n6 27.5996
R76 VTAIL.n9 VTAIL.n7 1.46602
R77 VTAIL.n10 VTAIL.n9 1.46602
R78 VTAIL.n13 VTAIL.n11 1.46602
R79 VTAIL.n14 VTAIL.n13 1.46602
R80 VTAIL.n6 VTAIL.n5 1.46602
R81 VTAIL.n5 VTAIL.n3 1.46602
R82 VTAIL.n2 VTAIL.n1 1.46602
R83 VTAIL VTAIL.n15 1.40783
R84 VTAIL.n0 VTAIL.t14 1.24032
R85 VTAIL.n0 VTAIL.t15 1.24032
R86 VTAIL.n4 VTAIL.t6 1.24032
R87 VTAIL.n4 VTAIL.t2 1.24032
R88 VTAIL.n12 VTAIL.t3 1.24032
R89 VTAIL.n12 VTAIL.t5 1.24032
R90 VTAIL.n8 VTAIL.t12 1.24032
R91 VTAIL.n8 VTAIL.t11 1.24032
R92 VTAIL.n11 VTAIL.n10 0.470328
R93 VTAIL.n3 VTAIL.n2 0.470328
R94 VTAIL VTAIL.n1 0.0586897
R95 VDD2.n2 VDD2.n1 59.7357
R96 VDD2.n2 VDD2.n0 59.7357
R97 VDD2 VDD2.n5 59.733
R98 VDD2.n4 VDD2.n3 59.0585
R99 VDD2.n4 VDD2.n2 44.0774
R100 VDD2.n5 VDD2.t2 1.24032
R101 VDD2.n5 VDD2.t3 1.24032
R102 VDD2.n3 VDD2.t6 1.24032
R103 VDD2.n3 VDD2.t7 1.24032
R104 VDD2.n1 VDD2.t5 1.24032
R105 VDD2.n1 VDD2.t4 1.24032
R106 VDD2.n0 VDD2.t0 1.24032
R107 VDD2.n0 VDD2.t1 1.24032
R108 VDD2 VDD2.n4 0.791448
R109 B.n857 B.n856 585
R110 B.n355 B.n120 585
R111 B.n354 B.n353 585
R112 B.n352 B.n351 585
R113 B.n350 B.n349 585
R114 B.n348 B.n347 585
R115 B.n346 B.n345 585
R116 B.n344 B.n343 585
R117 B.n342 B.n341 585
R118 B.n340 B.n339 585
R119 B.n338 B.n337 585
R120 B.n336 B.n335 585
R121 B.n334 B.n333 585
R122 B.n332 B.n331 585
R123 B.n330 B.n329 585
R124 B.n328 B.n327 585
R125 B.n326 B.n325 585
R126 B.n324 B.n323 585
R127 B.n322 B.n321 585
R128 B.n320 B.n319 585
R129 B.n318 B.n317 585
R130 B.n316 B.n315 585
R131 B.n314 B.n313 585
R132 B.n312 B.n311 585
R133 B.n310 B.n309 585
R134 B.n308 B.n307 585
R135 B.n306 B.n305 585
R136 B.n304 B.n303 585
R137 B.n302 B.n301 585
R138 B.n300 B.n299 585
R139 B.n298 B.n297 585
R140 B.n296 B.n295 585
R141 B.n294 B.n293 585
R142 B.n292 B.n291 585
R143 B.n290 B.n289 585
R144 B.n288 B.n287 585
R145 B.n286 B.n285 585
R146 B.n284 B.n283 585
R147 B.n282 B.n281 585
R148 B.n280 B.n279 585
R149 B.n278 B.n277 585
R150 B.n276 B.n275 585
R151 B.n274 B.n273 585
R152 B.n272 B.n271 585
R153 B.n270 B.n269 585
R154 B.n268 B.n267 585
R155 B.n266 B.n265 585
R156 B.n264 B.n263 585
R157 B.n262 B.n261 585
R158 B.n260 B.n259 585
R159 B.n258 B.n257 585
R160 B.n256 B.n255 585
R161 B.n254 B.n253 585
R162 B.n251 B.n250 585
R163 B.n249 B.n248 585
R164 B.n247 B.n246 585
R165 B.n245 B.n244 585
R166 B.n243 B.n242 585
R167 B.n241 B.n240 585
R168 B.n239 B.n238 585
R169 B.n237 B.n236 585
R170 B.n235 B.n234 585
R171 B.n233 B.n232 585
R172 B.n230 B.n229 585
R173 B.n228 B.n227 585
R174 B.n226 B.n225 585
R175 B.n224 B.n223 585
R176 B.n222 B.n221 585
R177 B.n220 B.n219 585
R178 B.n218 B.n217 585
R179 B.n216 B.n215 585
R180 B.n214 B.n213 585
R181 B.n212 B.n211 585
R182 B.n210 B.n209 585
R183 B.n208 B.n207 585
R184 B.n206 B.n205 585
R185 B.n204 B.n203 585
R186 B.n202 B.n201 585
R187 B.n200 B.n199 585
R188 B.n198 B.n197 585
R189 B.n196 B.n195 585
R190 B.n194 B.n193 585
R191 B.n192 B.n191 585
R192 B.n190 B.n189 585
R193 B.n188 B.n187 585
R194 B.n186 B.n185 585
R195 B.n184 B.n183 585
R196 B.n182 B.n181 585
R197 B.n180 B.n179 585
R198 B.n178 B.n177 585
R199 B.n176 B.n175 585
R200 B.n174 B.n173 585
R201 B.n172 B.n171 585
R202 B.n170 B.n169 585
R203 B.n168 B.n167 585
R204 B.n166 B.n165 585
R205 B.n164 B.n163 585
R206 B.n162 B.n161 585
R207 B.n160 B.n159 585
R208 B.n158 B.n157 585
R209 B.n156 B.n155 585
R210 B.n154 B.n153 585
R211 B.n152 B.n151 585
R212 B.n150 B.n149 585
R213 B.n148 B.n147 585
R214 B.n146 B.n145 585
R215 B.n144 B.n143 585
R216 B.n142 B.n141 585
R217 B.n140 B.n139 585
R218 B.n138 B.n137 585
R219 B.n136 B.n135 585
R220 B.n134 B.n133 585
R221 B.n132 B.n131 585
R222 B.n130 B.n129 585
R223 B.n128 B.n127 585
R224 B.n126 B.n125 585
R225 B.n855 B.n62 585
R226 B.n860 B.n62 585
R227 B.n854 B.n61 585
R228 B.n861 B.n61 585
R229 B.n853 B.n852 585
R230 B.n852 B.n57 585
R231 B.n851 B.n56 585
R232 B.n867 B.n56 585
R233 B.n850 B.n55 585
R234 B.n868 B.n55 585
R235 B.n849 B.n54 585
R236 B.n869 B.n54 585
R237 B.n848 B.n847 585
R238 B.n847 B.n50 585
R239 B.n846 B.n49 585
R240 B.n875 B.n49 585
R241 B.n845 B.n48 585
R242 B.n876 B.n48 585
R243 B.n844 B.n47 585
R244 B.n877 B.n47 585
R245 B.n843 B.n842 585
R246 B.n842 B.n43 585
R247 B.n841 B.n42 585
R248 B.n883 B.n42 585
R249 B.n840 B.n41 585
R250 B.n884 B.n41 585
R251 B.n839 B.n40 585
R252 B.n885 B.n40 585
R253 B.n838 B.n837 585
R254 B.n837 B.n36 585
R255 B.n836 B.n35 585
R256 B.n891 B.n35 585
R257 B.n835 B.n34 585
R258 B.n892 B.n34 585
R259 B.n834 B.n33 585
R260 B.n893 B.n33 585
R261 B.n833 B.n832 585
R262 B.n832 B.n32 585
R263 B.n831 B.n28 585
R264 B.n899 B.n28 585
R265 B.n830 B.n27 585
R266 B.n900 B.n27 585
R267 B.n829 B.n26 585
R268 B.n901 B.n26 585
R269 B.n828 B.n827 585
R270 B.n827 B.n22 585
R271 B.n826 B.n21 585
R272 B.n907 B.n21 585
R273 B.n825 B.n20 585
R274 B.n908 B.n20 585
R275 B.n824 B.n19 585
R276 B.n909 B.n19 585
R277 B.n823 B.n822 585
R278 B.n822 B.n15 585
R279 B.n821 B.n14 585
R280 B.n915 B.n14 585
R281 B.n820 B.n13 585
R282 B.n916 B.n13 585
R283 B.n819 B.n12 585
R284 B.n917 B.n12 585
R285 B.n818 B.n817 585
R286 B.n817 B.n8 585
R287 B.n816 B.n7 585
R288 B.n923 B.n7 585
R289 B.n815 B.n6 585
R290 B.n924 B.n6 585
R291 B.n814 B.n5 585
R292 B.n925 B.n5 585
R293 B.n813 B.n812 585
R294 B.n812 B.n4 585
R295 B.n811 B.n356 585
R296 B.n811 B.n810 585
R297 B.n801 B.n357 585
R298 B.n358 B.n357 585
R299 B.n803 B.n802 585
R300 B.n804 B.n803 585
R301 B.n800 B.n362 585
R302 B.n366 B.n362 585
R303 B.n799 B.n798 585
R304 B.n798 B.n797 585
R305 B.n364 B.n363 585
R306 B.n365 B.n364 585
R307 B.n790 B.n789 585
R308 B.n791 B.n790 585
R309 B.n788 B.n371 585
R310 B.n371 B.n370 585
R311 B.n787 B.n786 585
R312 B.n786 B.n785 585
R313 B.n373 B.n372 585
R314 B.n374 B.n373 585
R315 B.n778 B.n777 585
R316 B.n779 B.n778 585
R317 B.n776 B.n379 585
R318 B.n379 B.n378 585
R319 B.n775 B.n774 585
R320 B.n774 B.n773 585
R321 B.n381 B.n380 585
R322 B.n766 B.n381 585
R323 B.n765 B.n764 585
R324 B.n767 B.n765 585
R325 B.n763 B.n386 585
R326 B.n386 B.n385 585
R327 B.n762 B.n761 585
R328 B.n761 B.n760 585
R329 B.n388 B.n387 585
R330 B.n389 B.n388 585
R331 B.n753 B.n752 585
R332 B.n754 B.n753 585
R333 B.n751 B.n394 585
R334 B.n394 B.n393 585
R335 B.n750 B.n749 585
R336 B.n749 B.n748 585
R337 B.n396 B.n395 585
R338 B.n397 B.n396 585
R339 B.n741 B.n740 585
R340 B.n742 B.n741 585
R341 B.n739 B.n402 585
R342 B.n402 B.n401 585
R343 B.n738 B.n737 585
R344 B.n737 B.n736 585
R345 B.n404 B.n403 585
R346 B.n405 B.n404 585
R347 B.n729 B.n728 585
R348 B.n730 B.n729 585
R349 B.n727 B.n410 585
R350 B.n410 B.n409 585
R351 B.n726 B.n725 585
R352 B.n725 B.n724 585
R353 B.n412 B.n411 585
R354 B.n413 B.n412 585
R355 B.n717 B.n716 585
R356 B.n718 B.n717 585
R357 B.n715 B.n418 585
R358 B.n418 B.n417 585
R359 B.n710 B.n709 585
R360 B.n708 B.n478 585
R361 B.n707 B.n477 585
R362 B.n712 B.n477 585
R363 B.n706 B.n705 585
R364 B.n704 B.n703 585
R365 B.n702 B.n701 585
R366 B.n700 B.n699 585
R367 B.n698 B.n697 585
R368 B.n696 B.n695 585
R369 B.n694 B.n693 585
R370 B.n692 B.n691 585
R371 B.n690 B.n689 585
R372 B.n688 B.n687 585
R373 B.n686 B.n685 585
R374 B.n684 B.n683 585
R375 B.n682 B.n681 585
R376 B.n680 B.n679 585
R377 B.n678 B.n677 585
R378 B.n676 B.n675 585
R379 B.n674 B.n673 585
R380 B.n672 B.n671 585
R381 B.n670 B.n669 585
R382 B.n668 B.n667 585
R383 B.n666 B.n665 585
R384 B.n664 B.n663 585
R385 B.n662 B.n661 585
R386 B.n660 B.n659 585
R387 B.n658 B.n657 585
R388 B.n656 B.n655 585
R389 B.n654 B.n653 585
R390 B.n652 B.n651 585
R391 B.n650 B.n649 585
R392 B.n648 B.n647 585
R393 B.n646 B.n645 585
R394 B.n644 B.n643 585
R395 B.n642 B.n641 585
R396 B.n640 B.n639 585
R397 B.n638 B.n637 585
R398 B.n636 B.n635 585
R399 B.n634 B.n633 585
R400 B.n632 B.n631 585
R401 B.n630 B.n629 585
R402 B.n628 B.n627 585
R403 B.n626 B.n625 585
R404 B.n624 B.n623 585
R405 B.n622 B.n621 585
R406 B.n620 B.n619 585
R407 B.n618 B.n617 585
R408 B.n616 B.n615 585
R409 B.n614 B.n613 585
R410 B.n612 B.n611 585
R411 B.n610 B.n609 585
R412 B.n608 B.n607 585
R413 B.n606 B.n605 585
R414 B.n604 B.n603 585
R415 B.n602 B.n601 585
R416 B.n600 B.n599 585
R417 B.n598 B.n597 585
R418 B.n596 B.n595 585
R419 B.n594 B.n593 585
R420 B.n592 B.n591 585
R421 B.n590 B.n589 585
R422 B.n588 B.n587 585
R423 B.n586 B.n585 585
R424 B.n584 B.n583 585
R425 B.n582 B.n581 585
R426 B.n580 B.n579 585
R427 B.n578 B.n577 585
R428 B.n576 B.n575 585
R429 B.n574 B.n573 585
R430 B.n572 B.n571 585
R431 B.n570 B.n569 585
R432 B.n568 B.n567 585
R433 B.n566 B.n565 585
R434 B.n564 B.n563 585
R435 B.n562 B.n561 585
R436 B.n560 B.n559 585
R437 B.n558 B.n557 585
R438 B.n556 B.n555 585
R439 B.n554 B.n553 585
R440 B.n552 B.n551 585
R441 B.n550 B.n549 585
R442 B.n548 B.n547 585
R443 B.n546 B.n545 585
R444 B.n544 B.n543 585
R445 B.n542 B.n541 585
R446 B.n540 B.n539 585
R447 B.n538 B.n537 585
R448 B.n536 B.n535 585
R449 B.n534 B.n533 585
R450 B.n532 B.n531 585
R451 B.n530 B.n529 585
R452 B.n528 B.n527 585
R453 B.n526 B.n525 585
R454 B.n524 B.n523 585
R455 B.n522 B.n521 585
R456 B.n520 B.n519 585
R457 B.n518 B.n517 585
R458 B.n516 B.n515 585
R459 B.n514 B.n513 585
R460 B.n512 B.n511 585
R461 B.n510 B.n509 585
R462 B.n508 B.n507 585
R463 B.n506 B.n505 585
R464 B.n504 B.n503 585
R465 B.n502 B.n501 585
R466 B.n500 B.n499 585
R467 B.n498 B.n497 585
R468 B.n496 B.n495 585
R469 B.n494 B.n493 585
R470 B.n492 B.n491 585
R471 B.n490 B.n489 585
R472 B.n488 B.n487 585
R473 B.n486 B.n485 585
R474 B.n420 B.n419 585
R475 B.n714 B.n713 585
R476 B.n713 B.n712 585
R477 B.n416 B.n415 585
R478 B.n417 B.n416 585
R479 B.n720 B.n719 585
R480 B.n719 B.n718 585
R481 B.n721 B.n414 585
R482 B.n414 B.n413 585
R483 B.n723 B.n722 585
R484 B.n724 B.n723 585
R485 B.n408 B.n407 585
R486 B.n409 B.n408 585
R487 B.n732 B.n731 585
R488 B.n731 B.n730 585
R489 B.n733 B.n406 585
R490 B.n406 B.n405 585
R491 B.n735 B.n734 585
R492 B.n736 B.n735 585
R493 B.n400 B.n399 585
R494 B.n401 B.n400 585
R495 B.n744 B.n743 585
R496 B.n743 B.n742 585
R497 B.n745 B.n398 585
R498 B.n398 B.n397 585
R499 B.n747 B.n746 585
R500 B.n748 B.n747 585
R501 B.n392 B.n391 585
R502 B.n393 B.n392 585
R503 B.n756 B.n755 585
R504 B.n755 B.n754 585
R505 B.n757 B.n390 585
R506 B.n390 B.n389 585
R507 B.n759 B.n758 585
R508 B.n760 B.n759 585
R509 B.n384 B.n383 585
R510 B.n385 B.n384 585
R511 B.n769 B.n768 585
R512 B.n768 B.n767 585
R513 B.n770 B.n382 585
R514 B.n766 B.n382 585
R515 B.n772 B.n771 585
R516 B.n773 B.n772 585
R517 B.n377 B.n376 585
R518 B.n378 B.n377 585
R519 B.n781 B.n780 585
R520 B.n780 B.n779 585
R521 B.n782 B.n375 585
R522 B.n375 B.n374 585
R523 B.n784 B.n783 585
R524 B.n785 B.n784 585
R525 B.n369 B.n368 585
R526 B.n370 B.n369 585
R527 B.n793 B.n792 585
R528 B.n792 B.n791 585
R529 B.n794 B.n367 585
R530 B.n367 B.n365 585
R531 B.n796 B.n795 585
R532 B.n797 B.n796 585
R533 B.n361 B.n360 585
R534 B.n366 B.n361 585
R535 B.n806 B.n805 585
R536 B.n805 B.n804 585
R537 B.n807 B.n359 585
R538 B.n359 B.n358 585
R539 B.n809 B.n808 585
R540 B.n810 B.n809 585
R541 B.n2 B.n0 585
R542 B.n4 B.n2 585
R543 B.n3 B.n1 585
R544 B.n924 B.n3 585
R545 B.n922 B.n921 585
R546 B.n923 B.n922 585
R547 B.n920 B.n9 585
R548 B.n9 B.n8 585
R549 B.n919 B.n918 585
R550 B.n918 B.n917 585
R551 B.n11 B.n10 585
R552 B.n916 B.n11 585
R553 B.n914 B.n913 585
R554 B.n915 B.n914 585
R555 B.n912 B.n16 585
R556 B.n16 B.n15 585
R557 B.n911 B.n910 585
R558 B.n910 B.n909 585
R559 B.n18 B.n17 585
R560 B.n908 B.n18 585
R561 B.n906 B.n905 585
R562 B.n907 B.n906 585
R563 B.n904 B.n23 585
R564 B.n23 B.n22 585
R565 B.n903 B.n902 585
R566 B.n902 B.n901 585
R567 B.n25 B.n24 585
R568 B.n900 B.n25 585
R569 B.n898 B.n897 585
R570 B.n899 B.n898 585
R571 B.n896 B.n29 585
R572 B.n32 B.n29 585
R573 B.n895 B.n894 585
R574 B.n894 B.n893 585
R575 B.n31 B.n30 585
R576 B.n892 B.n31 585
R577 B.n890 B.n889 585
R578 B.n891 B.n890 585
R579 B.n888 B.n37 585
R580 B.n37 B.n36 585
R581 B.n887 B.n886 585
R582 B.n886 B.n885 585
R583 B.n39 B.n38 585
R584 B.n884 B.n39 585
R585 B.n882 B.n881 585
R586 B.n883 B.n882 585
R587 B.n880 B.n44 585
R588 B.n44 B.n43 585
R589 B.n879 B.n878 585
R590 B.n878 B.n877 585
R591 B.n46 B.n45 585
R592 B.n876 B.n46 585
R593 B.n874 B.n873 585
R594 B.n875 B.n874 585
R595 B.n872 B.n51 585
R596 B.n51 B.n50 585
R597 B.n871 B.n870 585
R598 B.n870 B.n869 585
R599 B.n53 B.n52 585
R600 B.n868 B.n53 585
R601 B.n866 B.n865 585
R602 B.n867 B.n866 585
R603 B.n864 B.n58 585
R604 B.n58 B.n57 585
R605 B.n863 B.n862 585
R606 B.n862 B.n861 585
R607 B.n60 B.n59 585
R608 B.n860 B.n60 585
R609 B.n927 B.n926 585
R610 B.n926 B.n925 585
R611 B.n710 B.n416 530.939
R612 B.n125 B.n60 530.939
R613 B.n713 B.n418 530.939
R614 B.n857 B.n62 530.939
R615 B.n482 B.t8 485.853
R616 B.n479 B.t19 485.853
R617 B.n123 B.t16 485.853
R618 B.n121 B.t12 485.853
R619 B.n859 B.n858 256.663
R620 B.n859 B.n119 256.663
R621 B.n859 B.n118 256.663
R622 B.n859 B.n117 256.663
R623 B.n859 B.n116 256.663
R624 B.n859 B.n115 256.663
R625 B.n859 B.n114 256.663
R626 B.n859 B.n113 256.663
R627 B.n859 B.n112 256.663
R628 B.n859 B.n111 256.663
R629 B.n859 B.n110 256.663
R630 B.n859 B.n109 256.663
R631 B.n859 B.n108 256.663
R632 B.n859 B.n107 256.663
R633 B.n859 B.n106 256.663
R634 B.n859 B.n105 256.663
R635 B.n859 B.n104 256.663
R636 B.n859 B.n103 256.663
R637 B.n859 B.n102 256.663
R638 B.n859 B.n101 256.663
R639 B.n859 B.n100 256.663
R640 B.n859 B.n99 256.663
R641 B.n859 B.n98 256.663
R642 B.n859 B.n97 256.663
R643 B.n859 B.n96 256.663
R644 B.n859 B.n95 256.663
R645 B.n859 B.n94 256.663
R646 B.n859 B.n93 256.663
R647 B.n859 B.n92 256.663
R648 B.n859 B.n91 256.663
R649 B.n859 B.n90 256.663
R650 B.n859 B.n89 256.663
R651 B.n859 B.n88 256.663
R652 B.n859 B.n87 256.663
R653 B.n859 B.n86 256.663
R654 B.n859 B.n85 256.663
R655 B.n859 B.n84 256.663
R656 B.n859 B.n83 256.663
R657 B.n859 B.n82 256.663
R658 B.n859 B.n81 256.663
R659 B.n859 B.n80 256.663
R660 B.n859 B.n79 256.663
R661 B.n859 B.n78 256.663
R662 B.n859 B.n77 256.663
R663 B.n859 B.n76 256.663
R664 B.n859 B.n75 256.663
R665 B.n859 B.n74 256.663
R666 B.n859 B.n73 256.663
R667 B.n859 B.n72 256.663
R668 B.n859 B.n71 256.663
R669 B.n859 B.n70 256.663
R670 B.n859 B.n69 256.663
R671 B.n859 B.n68 256.663
R672 B.n859 B.n67 256.663
R673 B.n859 B.n66 256.663
R674 B.n859 B.n65 256.663
R675 B.n859 B.n64 256.663
R676 B.n859 B.n63 256.663
R677 B.n712 B.n711 256.663
R678 B.n712 B.n421 256.663
R679 B.n712 B.n422 256.663
R680 B.n712 B.n423 256.663
R681 B.n712 B.n424 256.663
R682 B.n712 B.n425 256.663
R683 B.n712 B.n426 256.663
R684 B.n712 B.n427 256.663
R685 B.n712 B.n428 256.663
R686 B.n712 B.n429 256.663
R687 B.n712 B.n430 256.663
R688 B.n712 B.n431 256.663
R689 B.n712 B.n432 256.663
R690 B.n712 B.n433 256.663
R691 B.n712 B.n434 256.663
R692 B.n712 B.n435 256.663
R693 B.n712 B.n436 256.663
R694 B.n712 B.n437 256.663
R695 B.n712 B.n438 256.663
R696 B.n712 B.n439 256.663
R697 B.n712 B.n440 256.663
R698 B.n712 B.n441 256.663
R699 B.n712 B.n442 256.663
R700 B.n712 B.n443 256.663
R701 B.n712 B.n444 256.663
R702 B.n712 B.n445 256.663
R703 B.n712 B.n446 256.663
R704 B.n712 B.n447 256.663
R705 B.n712 B.n448 256.663
R706 B.n712 B.n449 256.663
R707 B.n712 B.n450 256.663
R708 B.n712 B.n451 256.663
R709 B.n712 B.n452 256.663
R710 B.n712 B.n453 256.663
R711 B.n712 B.n454 256.663
R712 B.n712 B.n455 256.663
R713 B.n712 B.n456 256.663
R714 B.n712 B.n457 256.663
R715 B.n712 B.n458 256.663
R716 B.n712 B.n459 256.663
R717 B.n712 B.n460 256.663
R718 B.n712 B.n461 256.663
R719 B.n712 B.n462 256.663
R720 B.n712 B.n463 256.663
R721 B.n712 B.n464 256.663
R722 B.n712 B.n465 256.663
R723 B.n712 B.n466 256.663
R724 B.n712 B.n467 256.663
R725 B.n712 B.n468 256.663
R726 B.n712 B.n469 256.663
R727 B.n712 B.n470 256.663
R728 B.n712 B.n471 256.663
R729 B.n712 B.n472 256.663
R730 B.n712 B.n473 256.663
R731 B.n712 B.n474 256.663
R732 B.n712 B.n475 256.663
R733 B.n712 B.n476 256.663
R734 B.n719 B.n416 163.367
R735 B.n719 B.n414 163.367
R736 B.n723 B.n414 163.367
R737 B.n723 B.n408 163.367
R738 B.n731 B.n408 163.367
R739 B.n731 B.n406 163.367
R740 B.n735 B.n406 163.367
R741 B.n735 B.n400 163.367
R742 B.n743 B.n400 163.367
R743 B.n743 B.n398 163.367
R744 B.n747 B.n398 163.367
R745 B.n747 B.n392 163.367
R746 B.n755 B.n392 163.367
R747 B.n755 B.n390 163.367
R748 B.n759 B.n390 163.367
R749 B.n759 B.n384 163.367
R750 B.n768 B.n384 163.367
R751 B.n768 B.n382 163.367
R752 B.n772 B.n382 163.367
R753 B.n772 B.n377 163.367
R754 B.n780 B.n377 163.367
R755 B.n780 B.n375 163.367
R756 B.n784 B.n375 163.367
R757 B.n784 B.n369 163.367
R758 B.n792 B.n369 163.367
R759 B.n792 B.n367 163.367
R760 B.n796 B.n367 163.367
R761 B.n796 B.n361 163.367
R762 B.n805 B.n361 163.367
R763 B.n805 B.n359 163.367
R764 B.n809 B.n359 163.367
R765 B.n809 B.n2 163.367
R766 B.n926 B.n2 163.367
R767 B.n926 B.n3 163.367
R768 B.n922 B.n3 163.367
R769 B.n922 B.n9 163.367
R770 B.n918 B.n9 163.367
R771 B.n918 B.n11 163.367
R772 B.n914 B.n11 163.367
R773 B.n914 B.n16 163.367
R774 B.n910 B.n16 163.367
R775 B.n910 B.n18 163.367
R776 B.n906 B.n18 163.367
R777 B.n906 B.n23 163.367
R778 B.n902 B.n23 163.367
R779 B.n902 B.n25 163.367
R780 B.n898 B.n25 163.367
R781 B.n898 B.n29 163.367
R782 B.n894 B.n29 163.367
R783 B.n894 B.n31 163.367
R784 B.n890 B.n31 163.367
R785 B.n890 B.n37 163.367
R786 B.n886 B.n37 163.367
R787 B.n886 B.n39 163.367
R788 B.n882 B.n39 163.367
R789 B.n882 B.n44 163.367
R790 B.n878 B.n44 163.367
R791 B.n878 B.n46 163.367
R792 B.n874 B.n46 163.367
R793 B.n874 B.n51 163.367
R794 B.n870 B.n51 163.367
R795 B.n870 B.n53 163.367
R796 B.n866 B.n53 163.367
R797 B.n866 B.n58 163.367
R798 B.n862 B.n58 163.367
R799 B.n862 B.n60 163.367
R800 B.n478 B.n477 163.367
R801 B.n705 B.n477 163.367
R802 B.n703 B.n702 163.367
R803 B.n699 B.n698 163.367
R804 B.n695 B.n694 163.367
R805 B.n691 B.n690 163.367
R806 B.n687 B.n686 163.367
R807 B.n683 B.n682 163.367
R808 B.n679 B.n678 163.367
R809 B.n675 B.n674 163.367
R810 B.n671 B.n670 163.367
R811 B.n667 B.n666 163.367
R812 B.n663 B.n662 163.367
R813 B.n659 B.n658 163.367
R814 B.n655 B.n654 163.367
R815 B.n651 B.n650 163.367
R816 B.n647 B.n646 163.367
R817 B.n643 B.n642 163.367
R818 B.n639 B.n638 163.367
R819 B.n635 B.n634 163.367
R820 B.n631 B.n630 163.367
R821 B.n627 B.n626 163.367
R822 B.n623 B.n622 163.367
R823 B.n619 B.n618 163.367
R824 B.n615 B.n614 163.367
R825 B.n611 B.n610 163.367
R826 B.n607 B.n606 163.367
R827 B.n603 B.n602 163.367
R828 B.n599 B.n598 163.367
R829 B.n595 B.n594 163.367
R830 B.n591 B.n590 163.367
R831 B.n587 B.n586 163.367
R832 B.n583 B.n582 163.367
R833 B.n579 B.n578 163.367
R834 B.n575 B.n574 163.367
R835 B.n571 B.n570 163.367
R836 B.n567 B.n566 163.367
R837 B.n563 B.n562 163.367
R838 B.n559 B.n558 163.367
R839 B.n555 B.n554 163.367
R840 B.n551 B.n550 163.367
R841 B.n547 B.n546 163.367
R842 B.n543 B.n542 163.367
R843 B.n539 B.n538 163.367
R844 B.n535 B.n534 163.367
R845 B.n531 B.n530 163.367
R846 B.n527 B.n526 163.367
R847 B.n523 B.n522 163.367
R848 B.n519 B.n518 163.367
R849 B.n515 B.n514 163.367
R850 B.n511 B.n510 163.367
R851 B.n507 B.n506 163.367
R852 B.n503 B.n502 163.367
R853 B.n499 B.n498 163.367
R854 B.n495 B.n494 163.367
R855 B.n491 B.n490 163.367
R856 B.n487 B.n486 163.367
R857 B.n713 B.n420 163.367
R858 B.n717 B.n418 163.367
R859 B.n717 B.n412 163.367
R860 B.n725 B.n412 163.367
R861 B.n725 B.n410 163.367
R862 B.n729 B.n410 163.367
R863 B.n729 B.n404 163.367
R864 B.n737 B.n404 163.367
R865 B.n737 B.n402 163.367
R866 B.n741 B.n402 163.367
R867 B.n741 B.n396 163.367
R868 B.n749 B.n396 163.367
R869 B.n749 B.n394 163.367
R870 B.n753 B.n394 163.367
R871 B.n753 B.n388 163.367
R872 B.n761 B.n388 163.367
R873 B.n761 B.n386 163.367
R874 B.n765 B.n386 163.367
R875 B.n765 B.n381 163.367
R876 B.n774 B.n381 163.367
R877 B.n774 B.n379 163.367
R878 B.n778 B.n379 163.367
R879 B.n778 B.n373 163.367
R880 B.n786 B.n373 163.367
R881 B.n786 B.n371 163.367
R882 B.n790 B.n371 163.367
R883 B.n790 B.n364 163.367
R884 B.n798 B.n364 163.367
R885 B.n798 B.n362 163.367
R886 B.n803 B.n362 163.367
R887 B.n803 B.n357 163.367
R888 B.n811 B.n357 163.367
R889 B.n812 B.n811 163.367
R890 B.n812 B.n5 163.367
R891 B.n6 B.n5 163.367
R892 B.n7 B.n6 163.367
R893 B.n817 B.n7 163.367
R894 B.n817 B.n12 163.367
R895 B.n13 B.n12 163.367
R896 B.n14 B.n13 163.367
R897 B.n822 B.n14 163.367
R898 B.n822 B.n19 163.367
R899 B.n20 B.n19 163.367
R900 B.n21 B.n20 163.367
R901 B.n827 B.n21 163.367
R902 B.n827 B.n26 163.367
R903 B.n27 B.n26 163.367
R904 B.n28 B.n27 163.367
R905 B.n832 B.n28 163.367
R906 B.n832 B.n33 163.367
R907 B.n34 B.n33 163.367
R908 B.n35 B.n34 163.367
R909 B.n837 B.n35 163.367
R910 B.n837 B.n40 163.367
R911 B.n41 B.n40 163.367
R912 B.n42 B.n41 163.367
R913 B.n842 B.n42 163.367
R914 B.n842 B.n47 163.367
R915 B.n48 B.n47 163.367
R916 B.n49 B.n48 163.367
R917 B.n847 B.n49 163.367
R918 B.n847 B.n54 163.367
R919 B.n55 B.n54 163.367
R920 B.n56 B.n55 163.367
R921 B.n852 B.n56 163.367
R922 B.n852 B.n61 163.367
R923 B.n62 B.n61 163.367
R924 B.n129 B.n128 163.367
R925 B.n133 B.n132 163.367
R926 B.n137 B.n136 163.367
R927 B.n141 B.n140 163.367
R928 B.n145 B.n144 163.367
R929 B.n149 B.n148 163.367
R930 B.n153 B.n152 163.367
R931 B.n157 B.n156 163.367
R932 B.n161 B.n160 163.367
R933 B.n165 B.n164 163.367
R934 B.n169 B.n168 163.367
R935 B.n173 B.n172 163.367
R936 B.n177 B.n176 163.367
R937 B.n181 B.n180 163.367
R938 B.n185 B.n184 163.367
R939 B.n189 B.n188 163.367
R940 B.n193 B.n192 163.367
R941 B.n197 B.n196 163.367
R942 B.n201 B.n200 163.367
R943 B.n205 B.n204 163.367
R944 B.n209 B.n208 163.367
R945 B.n213 B.n212 163.367
R946 B.n217 B.n216 163.367
R947 B.n221 B.n220 163.367
R948 B.n225 B.n224 163.367
R949 B.n229 B.n228 163.367
R950 B.n234 B.n233 163.367
R951 B.n238 B.n237 163.367
R952 B.n242 B.n241 163.367
R953 B.n246 B.n245 163.367
R954 B.n250 B.n249 163.367
R955 B.n255 B.n254 163.367
R956 B.n259 B.n258 163.367
R957 B.n263 B.n262 163.367
R958 B.n267 B.n266 163.367
R959 B.n271 B.n270 163.367
R960 B.n275 B.n274 163.367
R961 B.n279 B.n278 163.367
R962 B.n283 B.n282 163.367
R963 B.n287 B.n286 163.367
R964 B.n291 B.n290 163.367
R965 B.n295 B.n294 163.367
R966 B.n299 B.n298 163.367
R967 B.n303 B.n302 163.367
R968 B.n307 B.n306 163.367
R969 B.n311 B.n310 163.367
R970 B.n315 B.n314 163.367
R971 B.n319 B.n318 163.367
R972 B.n323 B.n322 163.367
R973 B.n327 B.n326 163.367
R974 B.n331 B.n330 163.367
R975 B.n335 B.n334 163.367
R976 B.n339 B.n338 163.367
R977 B.n343 B.n342 163.367
R978 B.n347 B.n346 163.367
R979 B.n351 B.n350 163.367
R980 B.n353 B.n120 163.367
R981 B.n482 B.t11 106.754
R982 B.n121 B.t14 106.754
R983 B.n479 B.t21 106.734
R984 B.n123 B.t17 106.734
R985 B.n483 B.t10 73.7852
R986 B.n122 B.t15 73.7852
R987 B.n480 B.t20 73.7645
R988 B.n124 B.t18 73.7645
R989 B.n711 B.n710 71.676
R990 B.n705 B.n421 71.676
R991 B.n702 B.n422 71.676
R992 B.n698 B.n423 71.676
R993 B.n694 B.n424 71.676
R994 B.n690 B.n425 71.676
R995 B.n686 B.n426 71.676
R996 B.n682 B.n427 71.676
R997 B.n678 B.n428 71.676
R998 B.n674 B.n429 71.676
R999 B.n670 B.n430 71.676
R1000 B.n666 B.n431 71.676
R1001 B.n662 B.n432 71.676
R1002 B.n658 B.n433 71.676
R1003 B.n654 B.n434 71.676
R1004 B.n650 B.n435 71.676
R1005 B.n646 B.n436 71.676
R1006 B.n642 B.n437 71.676
R1007 B.n638 B.n438 71.676
R1008 B.n634 B.n439 71.676
R1009 B.n630 B.n440 71.676
R1010 B.n626 B.n441 71.676
R1011 B.n622 B.n442 71.676
R1012 B.n618 B.n443 71.676
R1013 B.n614 B.n444 71.676
R1014 B.n610 B.n445 71.676
R1015 B.n606 B.n446 71.676
R1016 B.n602 B.n447 71.676
R1017 B.n598 B.n448 71.676
R1018 B.n594 B.n449 71.676
R1019 B.n590 B.n450 71.676
R1020 B.n586 B.n451 71.676
R1021 B.n582 B.n452 71.676
R1022 B.n578 B.n453 71.676
R1023 B.n574 B.n454 71.676
R1024 B.n570 B.n455 71.676
R1025 B.n566 B.n456 71.676
R1026 B.n562 B.n457 71.676
R1027 B.n558 B.n458 71.676
R1028 B.n554 B.n459 71.676
R1029 B.n550 B.n460 71.676
R1030 B.n546 B.n461 71.676
R1031 B.n542 B.n462 71.676
R1032 B.n538 B.n463 71.676
R1033 B.n534 B.n464 71.676
R1034 B.n530 B.n465 71.676
R1035 B.n526 B.n466 71.676
R1036 B.n522 B.n467 71.676
R1037 B.n518 B.n468 71.676
R1038 B.n514 B.n469 71.676
R1039 B.n510 B.n470 71.676
R1040 B.n506 B.n471 71.676
R1041 B.n502 B.n472 71.676
R1042 B.n498 B.n473 71.676
R1043 B.n494 B.n474 71.676
R1044 B.n490 B.n475 71.676
R1045 B.n486 B.n476 71.676
R1046 B.n125 B.n63 71.676
R1047 B.n129 B.n64 71.676
R1048 B.n133 B.n65 71.676
R1049 B.n137 B.n66 71.676
R1050 B.n141 B.n67 71.676
R1051 B.n145 B.n68 71.676
R1052 B.n149 B.n69 71.676
R1053 B.n153 B.n70 71.676
R1054 B.n157 B.n71 71.676
R1055 B.n161 B.n72 71.676
R1056 B.n165 B.n73 71.676
R1057 B.n169 B.n74 71.676
R1058 B.n173 B.n75 71.676
R1059 B.n177 B.n76 71.676
R1060 B.n181 B.n77 71.676
R1061 B.n185 B.n78 71.676
R1062 B.n189 B.n79 71.676
R1063 B.n193 B.n80 71.676
R1064 B.n197 B.n81 71.676
R1065 B.n201 B.n82 71.676
R1066 B.n205 B.n83 71.676
R1067 B.n209 B.n84 71.676
R1068 B.n213 B.n85 71.676
R1069 B.n217 B.n86 71.676
R1070 B.n221 B.n87 71.676
R1071 B.n225 B.n88 71.676
R1072 B.n229 B.n89 71.676
R1073 B.n234 B.n90 71.676
R1074 B.n238 B.n91 71.676
R1075 B.n242 B.n92 71.676
R1076 B.n246 B.n93 71.676
R1077 B.n250 B.n94 71.676
R1078 B.n255 B.n95 71.676
R1079 B.n259 B.n96 71.676
R1080 B.n263 B.n97 71.676
R1081 B.n267 B.n98 71.676
R1082 B.n271 B.n99 71.676
R1083 B.n275 B.n100 71.676
R1084 B.n279 B.n101 71.676
R1085 B.n283 B.n102 71.676
R1086 B.n287 B.n103 71.676
R1087 B.n291 B.n104 71.676
R1088 B.n295 B.n105 71.676
R1089 B.n299 B.n106 71.676
R1090 B.n303 B.n107 71.676
R1091 B.n307 B.n108 71.676
R1092 B.n311 B.n109 71.676
R1093 B.n315 B.n110 71.676
R1094 B.n319 B.n111 71.676
R1095 B.n323 B.n112 71.676
R1096 B.n327 B.n113 71.676
R1097 B.n331 B.n114 71.676
R1098 B.n335 B.n115 71.676
R1099 B.n339 B.n116 71.676
R1100 B.n343 B.n117 71.676
R1101 B.n347 B.n118 71.676
R1102 B.n351 B.n119 71.676
R1103 B.n858 B.n120 71.676
R1104 B.n858 B.n857 71.676
R1105 B.n353 B.n119 71.676
R1106 B.n350 B.n118 71.676
R1107 B.n346 B.n117 71.676
R1108 B.n342 B.n116 71.676
R1109 B.n338 B.n115 71.676
R1110 B.n334 B.n114 71.676
R1111 B.n330 B.n113 71.676
R1112 B.n326 B.n112 71.676
R1113 B.n322 B.n111 71.676
R1114 B.n318 B.n110 71.676
R1115 B.n314 B.n109 71.676
R1116 B.n310 B.n108 71.676
R1117 B.n306 B.n107 71.676
R1118 B.n302 B.n106 71.676
R1119 B.n298 B.n105 71.676
R1120 B.n294 B.n104 71.676
R1121 B.n290 B.n103 71.676
R1122 B.n286 B.n102 71.676
R1123 B.n282 B.n101 71.676
R1124 B.n278 B.n100 71.676
R1125 B.n274 B.n99 71.676
R1126 B.n270 B.n98 71.676
R1127 B.n266 B.n97 71.676
R1128 B.n262 B.n96 71.676
R1129 B.n258 B.n95 71.676
R1130 B.n254 B.n94 71.676
R1131 B.n249 B.n93 71.676
R1132 B.n245 B.n92 71.676
R1133 B.n241 B.n91 71.676
R1134 B.n237 B.n90 71.676
R1135 B.n233 B.n89 71.676
R1136 B.n228 B.n88 71.676
R1137 B.n224 B.n87 71.676
R1138 B.n220 B.n86 71.676
R1139 B.n216 B.n85 71.676
R1140 B.n212 B.n84 71.676
R1141 B.n208 B.n83 71.676
R1142 B.n204 B.n82 71.676
R1143 B.n200 B.n81 71.676
R1144 B.n196 B.n80 71.676
R1145 B.n192 B.n79 71.676
R1146 B.n188 B.n78 71.676
R1147 B.n184 B.n77 71.676
R1148 B.n180 B.n76 71.676
R1149 B.n176 B.n75 71.676
R1150 B.n172 B.n74 71.676
R1151 B.n168 B.n73 71.676
R1152 B.n164 B.n72 71.676
R1153 B.n160 B.n71 71.676
R1154 B.n156 B.n70 71.676
R1155 B.n152 B.n69 71.676
R1156 B.n148 B.n68 71.676
R1157 B.n144 B.n67 71.676
R1158 B.n140 B.n66 71.676
R1159 B.n136 B.n65 71.676
R1160 B.n132 B.n64 71.676
R1161 B.n128 B.n63 71.676
R1162 B.n711 B.n478 71.676
R1163 B.n703 B.n421 71.676
R1164 B.n699 B.n422 71.676
R1165 B.n695 B.n423 71.676
R1166 B.n691 B.n424 71.676
R1167 B.n687 B.n425 71.676
R1168 B.n683 B.n426 71.676
R1169 B.n679 B.n427 71.676
R1170 B.n675 B.n428 71.676
R1171 B.n671 B.n429 71.676
R1172 B.n667 B.n430 71.676
R1173 B.n663 B.n431 71.676
R1174 B.n659 B.n432 71.676
R1175 B.n655 B.n433 71.676
R1176 B.n651 B.n434 71.676
R1177 B.n647 B.n435 71.676
R1178 B.n643 B.n436 71.676
R1179 B.n639 B.n437 71.676
R1180 B.n635 B.n438 71.676
R1181 B.n631 B.n439 71.676
R1182 B.n627 B.n440 71.676
R1183 B.n623 B.n441 71.676
R1184 B.n619 B.n442 71.676
R1185 B.n615 B.n443 71.676
R1186 B.n611 B.n444 71.676
R1187 B.n607 B.n445 71.676
R1188 B.n603 B.n446 71.676
R1189 B.n599 B.n447 71.676
R1190 B.n595 B.n448 71.676
R1191 B.n591 B.n449 71.676
R1192 B.n587 B.n450 71.676
R1193 B.n583 B.n451 71.676
R1194 B.n579 B.n452 71.676
R1195 B.n575 B.n453 71.676
R1196 B.n571 B.n454 71.676
R1197 B.n567 B.n455 71.676
R1198 B.n563 B.n456 71.676
R1199 B.n559 B.n457 71.676
R1200 B.n555 B.n458 71.676
R1201 B.n551 B.n459 71.676
R1202 B.n547 B.n460 71.676
R1203 B.n543 B.n461 71.676
R1204 B.n539 B.n462 71.676
R1205 B.n535 B.n463 71.676
R1206 B.n531 B.n464 71.676
R1207 B.n527 B.n465 71.676
R1208 B.n523 B.n466 71.676
R1209 B.n519 B.n467 71.676
R1210 B.n515 B.n468 71.676
R1211 B.n511 B.n469 71.676
R1212 B.n507 B.n470 71.676
R1213 B.n503 B.n471 71.676
R1214 B.n499 B.n472 71.676
R1215 B.n495 B.n473 71.676
R1216 B.n491 B.n474 71.676
R1217 B.n487 B.n475 71.676
R1218 B.n476 B.n420 71.676
R1219 B.n712 B.n417 67.8282
R1220 B.n860 B.n859 67.8282
R1221 B.n484 B.n483 59.5399
R1222 B.n481 B.n480 59.5399
R1223 B.n231 B.n124 59.5399
R1224 B.n252 B.n122 59.5399
R1225 B.n718 B.n417 35.2088
R1226 B.n718 B.n413 35.2088
R1227 B.n724 B.n413 35.2088
R1228 B.n724 B.n409 35.2088
R1229 B.n730 B.n409 35.2088
R1230 B.n736 B.n405 35.2088
R1231 B.n736 B.n401 35.2088
R1232 B.n742 B.n401 35.2088
R1233 B.n742 B.n397 35.2088
R1234 B.n748 B.n397 35.2088
R1235 B.n748 B.n393 35.2088
R1236 B.n754 B.n393 35.2088
R1237 B.n760 B.n389 35.2088
R1238 B.n760 B.n385 35.2088
R1239 B.n767 B.n385 35.2088
R1240 B.n767 B.n766 35.2088
R1241 B.n773 B.n378 35.2088
R1242 B.n779 B.n378 35.2088
R1243 B.n779 B.n374 35.2088
R1244 B.n785 B.n374 35.2088
R1245 B.n791 B.n370 35.2088
R1246 B.n791 B.n365 35.2088
R1247 B.n797 B.n365 35.2088
R1248 B.n797 B.n366 35.2088
R1249 B.n804 B.n358 35.2088
R1250 B.n810 B.n358 35.2088
R1251 B.n810 B.n4 35.2088
R1252 B.n925 B.n4 35.2088
R1253 B.n925 B.n924 35.2088
R1254 B.n924 B.n923 35.2088
R1255 B.n923 B.n8 35.2088
R1256 B.n917 B.n8 35.2088
R1257 B.n916 B.n915 35.2088
R1258 B.n915 B.n15 35.2088
R1259 B.n909 B.n15 35.2088
R1260 B.n909 B.n908 35.2088
R1261 B.n907 B.n22 35.2088
R1262 B.n901 B.n22 35.2088
R1263 B.n901 B.n900 35.2088
R1264 B.n900 B.n899 35.2088
R1265 B.n893 B.n32 35.2088
R1266 B.n893 B.n892 35.2088
R1267 B.n892 B.n891 35.2088
R1268 B.n891 B.n36 35.2088
R1269 B.n885 B.n884 35.2088
R1270 B.n884 B.n883 35.2088
R1271 B.n883 B.n43 35.2088
R1272 B.n877 B.n43 35.2088
R1273 B.n877 B.n876 35.2088
R1274 B.n876 B.n875 35.2088
R1275 B.n875 B.n50 35.2088
R1276 B.n869 B.n868 35.2088
R1277 B.n868 B.n867 35.2088
R1278 B.n867 B.n57 35.2088
R1279 B.n861 B.n57 35.2088
R1280 B.n861 B.n860 35.2088
R1281 B.n126 B.n59 34.4981
R1282 B.n856 B.n855 34.4981
R1283 B.n715 B.n714 34.4981
R1284 B.n709 B.n415 34.4981
R1285 B.n483 B.n482 32.9702
R1286 B.n480 B.n479 32.9702
R1287 B.n124 B.n123 32.9702
R1288 B.n122 B.n121 32.9702
R1289 B.n754 B.t0 31.5844
R1290 B.n766 B.t6 31.5844
R1291 B.n785 B.t2 31.5844
R1292 B.n366 B.t7 31.5844
R1293 B.t4 B.n916 31.5844
R1294 B.t3 B.n907 31.5844
R1295 B.n32 B.t5 31.5844
R1296 B.n885 B.t1 31.5844
R1297 B.n730 B.t9 24.3356
R1298 B.n869 B.t13 24.3356
R1299 B B.n927 18.0485
R1300 B.t9 B.n405 10.8736
R1301 B.t13 B.n50 10.8736
R1302 B.n127 B.n126 10.6151
R1303 B.n130 B.n127 10.6151
R1304 B.n131 B.n130 10.6151
R1305 B.n134 B.n131 10.6151
R1306 B.n135 B.n134 10.6151
R1307 B.n138 B.n135 10.6151
R1308 B.n139 B.n138 10.6151
R1309 B.n142 B.n139 10.6151
R1310 B.n143 B.n142 10.6151
R1311 B.n146 B.n143 10.6151
R1312 B.n147 B.n146 10.6151
R1313 B.n150 B.n147 10.6151
R1314 B.n151 B.n150 10.6151
R1315 B.n154 B.n151 10.6151
R1316 B.n155 B.n154 10.6151
R1317 B.n158 B.n155 10.6151
R1318 B.n159 B.n158 10.6151
R1319 B.n162 B.n159 10.6151
R1320 B.n163 B.n162 10.6151
R1321 B.n166 B.n163 10.6151
R1322 B.n167 B.n166 10.6151
R1323 B.n170 B.n167 10.6151
R1324 B.n171 B.n170 10.6151
R1325 B.n174 B.n171 10.6151
R1326 B.n175 B.n174 10.6151
R1327 B.n178 B.n175 10.6151
R1328 B.n179 B.n178 10.6151
R1329 B.n182 B.n179 10.6151
R1330 B.n183 B.n182 10.6151
R1331 B.n186 B.n183 10.6151
R1332 B.n187 B.n186 10.6151
R1333 B.n190 B.n187 10.6151
R1334 B.n191 B.n190 10.6151
R1335 B.n194 B.n191 10.6151
R1336 B.n195 B.n194 10.6151
R1337 B.n198 B.n195 10.6151
R1338 B.n199 B.n198 10.6151
R1339 B.n202 B.n199 10.6151
R1340 B.n203 B.n202 10.6151
R1341 B.n206 B.n203 10.6151
R1342 B.n207 B.n206 10.6151
R1343 B.n210 B.n207 10.6151
R1344 B.n211 B.n210 10.6151
R1345 B.n214 B.n211 10.6151
R1346 B.n215 B.n214 10.6151
R1347 B.n218 B.n215 10.6151
R1348 B.n219 B.n218 10.6151
R1349 B.n222 B.n219 10.6151
R1350 B.n223 B.n222 10.6151
R1351 B.n226 B.n223 10.6151
R1352 B.n227 B.n226 10.6151
R1353 B.n230 B.n227 10.6151
R1354 B.n235 B.n232 10.6151
R1355 B.n236 B.n235 10.6151
R1356 B.n239 B.n236 10.6151
R1357 B.n240 B.n239 10.6151
R1358 B.n243 B.n240 10.6151
R1359 B.n244 B.n243 10.6151
R1360 B.n247 B.n244 10.6151
R1361 B.n248 B.n247 10.6151
R1362 B.n251 B.n248 10.6151
R1363 B.n256 B.n253 10.6151
R1364 B.n257 B.n256 10.6151
R1365 B.n260 B.n257 10.6151
R1366 B.n261 B.n260 10.6151
R1367 B.n264 B.n261 10.6151
R1368 B.n265 B.n264 10.6151
R1369 B.n268 B.n265 10.6151
R1370 B.n269 B.n268 10.6151
R1371 B.n272 B.n269 10.6151
R1372 B.n273 B.n272 10.6151
R1373 B.n276 B.n273 10.6151
R1374 B.n277 B.n276 10.6151
R1375 B.n280 B.n277 10.6151
R1376 B.n281 B.n280 10.6151
R1377 B.n284 B.n281 10.6151
R1378 B.n285 B.n284 10.6151
R1379 B.n288 B.n285 10.6151
R1380 B.n289 B.n288 10.6151
R1381 B.n292 B.n289 10.6151
R1382 B.n293 B.n292 10.6151
R1383 B.n296 B.n293 10.6151
R1384 B.n297 B.n296 10.6151
R1385 B.n300 B.n297 10.6151
R1386 B.n301 B.n300 10.6151
R1387 B.n304 B.n301 10.6151
R1388 B.n305 B.n304 10.6151
R1389 B.n308 B.n305 10.6151
R1390 B.n309 B.n308 10.6151
R1391 B.n312 B.n309 10.6151
R1392 B.n313 B.n312 10.6151
R1393 B.n316 B.n313 10.6151
R1394 B.n317 B.n316 10.6151
R1395 B.n320 B.n317 10.6151
R1396 B.n321 B.n320 10.6151
R1397 B.n324 B.n321 10.6151
R1398 B.n325 B.n324 10.6151
R1399 B.n328 B.n325 10.6151
R1400 B.n329 B.n328 10.6151
R1401 B.n332 B.n329 10.6151
R1402 B.n333 B.n332 10.6151
R1403 B.n336 B.n333 10.6151
R1404 B.n337 B.n336 10.6151
R1405 B.n340 B.n337 10.6151
R1406 B.n341 B.n340 10.6151
R1407 B.n344 B.n341 10.6151
R1408 B.n345 B.n344 10.6151
R1409 B.n348 B.n345 10.6151
R1410 B.n349 B.n348 10.6151
R1411 B.n352 B.n349 10.6151
R1412 B.n354 B.n352 10.6151
R1413 B.n355 B.n354 10.6151
R1414 B.n856 B.n355 10.6151
R1415 B.n716 B.n715 10.6151
R1416 B.n716 B.n411 10.6151
R1417 B.n726 B.n411 10.6151
R1418 B.n727 B.n726 10.6151
R1419 B.n728 B.n727 10.6151
R1420 B.n728 B.n403 10.6151
R1421 B.n738 B.n403 10.6151
R1422 B.n739 B.n738 10.6151
R1423 B.n740 B.n739 10.6151
R1424 B.n740 B.n395 10.6151
R1425 B.n750 B.n395 10.6151
R1426 B.n751 B.n750 10.6151
R1427 B.n752 B.n751 10.6151
R1428 B.n752 B.n387 10.6151
R1429 B.n762 B.n387 10.6151
R1430 B.n763 B.n762 10.6151
R1431 B.n764 B.n763 10.6151
R1432 B.n764 B.n380 10.6151
R1433 B.n775 B.n380 10.6151
R1434 B.n776 B.n775 10.6151
R1435 B.n777 B.n776 10.6151
R1436 B.n777 B.n372 10.6151
R1437 B.n787 B.n372 10.6151
R1438 B.n788 B.n787 10.6151
R1439 B.n789 B.n788 10.6151
R1440 B.n789 B.n363 10.6151
R1441 B.n799 B.n363 10.6151
R1442 B.n800 B.n799 10.6151
R1443 B.n802 B.n800 10.6151
R1444 B.n802 B.n801 10.6151
R1445 B.n801 B.n356 10.6151
R1446 B.n813 B.n356 10.6151
R1447 B.n814 B.n813 10.6151
R1448 B.n815 B.n814 10.6151
R1449 B.n816 B.n815 10.6151
R1450 B.n818 B.n816 10.6151
R1451 B.n819 B.n818 10.6151
R1452 B.n820 B.n819 10.6151
R1453 B.n821 B.n820 10.6151
R1454 B.n823 B.n821 10.6151
R1455 B.n824 B.n823 10.6151
R1456 B.n825 B.n824 10.6151
R1457 B.n826 B.n825 10.6151
R1458 B.n828 B.n826 10.6151
R1459 B.n829 B.n828 10.6151
R1460 B.n830 B.n829 10.6151
R1461 B.n831 B.n830 10.6151
R1462 B.n833 B.n831 10.6151
R1463 B.n834 B.n833 10.6151
R1464 B.n835 B.n834 10.6151
R1465 B.n836 B.n835 10.6151
R1466 B.n838 B.n836 10.6151
R1467 B.n839 B.n838 10.6151
R1468 B.n840 B.n839 10.6151
R1469 B.n841 B.n840 10.6151
R1470 B.n843 B.n841 10.6151
R1471 B.n844 B.n843 10.6151
R1472 B.n845 B.n844 10.6151
R1473 B.n846 B.n845 10.6151
R1474 B.n848 B.n846 10.6151
R1475 B.n849 B.n848 10.6151
R1476 B.n850 B.n849 10.6151
R1477 B.n851 B.n850 10.6151
R1478 B.n853 B.n851 10.6151
R1479 B.n854 B.n853 10.6151
R1480 B.n855 B.n854 10.6151
R1481 B.n709 B.n708 10.6151
R1482 B.n708 B.n707 10.6151
R1483 B.n707 B.n706 10.6151
R1484 B.n706 B.n704 10.6151
R1485 B.n704 B.n701 10.6151
R1486 B.n701 B.n700 10.6151
R1487 B.n700 B.n697 10.6151
R1488 B.n697 B.n696 10.6151
R1489 B.n696 B.n693 10.6151
R1490 B.n693 B.n692 10.6151
R1491 B.n692 B.n689 10.6151
R1492 B.n689 B.n688 10.6151
R1493 B.n688 B.n685 10.6151
R1494 B.n685 B.n684 10.6151
R1495 B.n684 B.n681 10.6151
R1496 B.n681 B.n680 10.6151
R1497 B.n680 B.n677 10.6151
R1498 B.n677 B.n676 10.6151
R1499 B.n676 B.n673 10.6151
R1500 B.n673 B.n672 10.6151
R1501 B.n672 B.n669 10.6151
R1502 B.n669 B.n668 10.6151
R1503 B.n668 B.n665 10.6151
R1504 B.n665 B.n664 10.6151
R1505 B.n664 B.n661 10.6151
R1506 B.n661 B.n660 10.6151
R1507 B.n660 B.n657 10.6151
R1508 B.n657 B.n656 10.6151
R1509 B.n656 B.n653 10.6151
R1510 B.n653 B.n652 10.6151
R1511 B.n652 B.n649 10.6151
R1512 B.n649 B.n648 10.6151
R1513 B.n648 B.n645 10.6151
R1514 B.n645 B.n644 10.6151
R1515 B.n644 B.n641 10.6151
R1516 B.n641 B.n640 10.6151
R1517 B.n640 B.n637 10.6151
R1518 B.n637 B.n636 10.6151
R1519 B.n636 B.n633 10.6151
R1520 B.n633 B.n632 10.6151
R1521 B.n632 B.n629 10.6151
R1522 B.n629 B.n628 10.6151
R1523 B.n628 B.n625 10.6151
R1524 B.n625 B.n624 10.6151
R1525 B.n624 B.n621 10.6151
R1526 B.n621 B.n620 10.6151
R1527 B.n620 B.n617 10.6151
R1528 B.n617 B.n616 10.6151
R1529 B.n616 B.n613 10.6151
R1530 B.n613 B.n612 10.6151
R1531 B.n612 B.n609 10.6151
R1532 B.n609 B.n608 10.6151
R1533 B.n605 B.n604 10.6151
R1534 B.n604 B.n601 10.6151
R1535 B.n601 B.n600 10.6151
R1536 B.n600 B.n597 10.6151
R1537 B.n597 B.n596 10.6151
R1538 B.n596 B.n593 10.6151
R1539 B.n593 B.n592 10.6151
R1540 B.n592 B.n589 10.6151
R1541 B.n589 B.n588 10.6151
R1542 B.n585 B.n584 10.6151
R1543 B.n584 B.n581 10.6151
R1544 B.n581 B.n580 10.6151
R1545 B.n580 B.n577 10.6151
R1546 B.n577 B.n576 10.6151
R1547 B.n576 B.n573 10.6151
R1548 B.n573 B.n572 10.6151
R1549 B.n572 B.n569 10.6151
R1550 B.n569 B.n568 10.6151
R1551 B.n568 B.n565 10.6151
R1552 B.n565 B.n564 10.6151
R1553 B.n564 B.n561 10.6151
R1554 B.n561 B.n560 10.6151
R1555 B.n560 B.n557 10.6151
R1556 B.n557 B.n556 10.6151
R1557 B.n556 B.n553 10.6151
R1558 B.n553 B.n552 10.6151
R1559 B.n552 B.n549 10.6151
R1560 B.n549 B.n548 10.6151
R1561 B.n548 B.n545 10.6151
R1562 B.n545 B.n544 10.6151
R1563 B.n544 B.n541 10.6151
R1564 B.n541 B.n540 10.6151
R1565 B.n540 B.n537 10.6151
R1566 B.n537 B.n536 10.6151
R1567 B.n536 B.n533 10.6151
R1568 B.n533 B.n532 10.6151
R1569 B.n532 B.n529 10.6151
R1570 B.n529 B.n528 10.6151
R1571 B.n528 B.n525 10.6151
R1572 B.n525 B.n524 10.6151
R1573 B.n524 B.n521 10.6151
R1574 B.n521 B.n520 10.6151
R1575 B.n520 B.n517 10.6151
R1576 B.n517 B.n516 10.6151
R1577 B.n516 B.n513 10.6151
R1578 B.n513 B.n512 10.6151
R1579 B.n512 B.n509 10.6151
R1580 B.n509 B.n508 10.6151
R1581 B.n508 B.n505 10.6151
R1582 B.n505 B.n504 10.6151
R1583 B.n504 B.n501 10.6151
R1584 B.n501 B.n500 10.6151
R1585 B.n500 B.n497 10.6151
R1586 B.n497 B.n496 10.6151
R1587 B.n496 B.n493 10.6151
R1588 B.n493 B.n492 10.6151
R1589 B.n492 B.n489 10.6151
R1590 B.n489 B.n488 10.6151
R1591 B.n488 B.n485 10.6151
R1592 B.n485 B.n419 10.6151
R1593 B.n714 B.n419 10.6151
R1594 B.n720 B.n415 10.6151
R1595 B.n721 B.n720 10.6151
R1596 B.n722 B.n721 10.6151
R1597 B.n722 B.n407 10.6151
R1598 B.n732 B.n407 10.6151
R1599 B.n733 B.n732 10.6151
R1600 B.n734 B.n733 10.6151
R1601 B.n734 B.n399 10.6151
R1602 B.n744 B.n399 10.6151
R1603 B.n745 B.n744 10.6151
R1604 B.n746 B.n745 10.6151
R1605 B.n746 B.n391 10.6151
R1606 B.n756 B.n391 10.6151
R1607 B.n757 B.n756 10.6151
R1608 B.n758 B.n757 10.6151
R1609 B.n758 B.n383 10.6151
R1610 B.n769 B.n383 10.6151
R1611 B.n770 B.n769 10.6151
R1612 B.n771 B.n770 10.6151
R1613 B.n771 B.n376 10.6151
R1614 B.n781 B.n376 10.6151
R1615 B.n782 B.n781 10.6151
R1616 B.n783 B.n782 10.6151
R1617 B.n783 B.n368 10.6151
R1618 B.n793 B.n368 10.6151
R1619 B.n794 B.n793 10.6151
R1620 B.n795 B.n794 10.6151
R1621 B.n795 B.n360 10.6151
R1622 B.n806 B.n360 10.6151
R1623 B.n807 B.n806 10.6151
R1624 B.n808 B.n807 10.6151
R1625 B.n808 B.n0 10.6151
R1626 B.n921 B.n1 10.6151
R1627 B.n921 B.n920 10.6151
R1628 B.n920 B.n919 10.6151
R1629 B.n919 B.n10 10.6151
R1630 B.n913 B.n10 10.6151
R1631 B.n913 B.n912 10.6151
R1632 B.n912 B.n911 10.6151
R1633 B.n911 B.n17 10.6151
R1634 B.n905 B.n17 10.6151
R1635 B.n905 B.n904 10.6151
R1636 B.n904 B.n903 10.6151
R1637 B.n903 B.n24 10.6151
R1638 B.n897 B.n24 10.6151
R1639 B.n897 B.n896 10.6151
R1640 B.n896 B.n895 10.6151
R1641 B.n895 B.n30 10.6151
R1642 B.n889 B.n30 10.6151
R1643 B.n889 B.n888 10.6151
R1644 B.n888 B.n887 10.6151
R1645 B.n887 B.n38 10.6151
R1646 B.n881 B.n38 10.6151
R1647 B.n881 B.n880 10.6151
R1648 B.n880 B.n879 10.6151
R1649 B.n879 B.n45 10.6151
R1650 B.n873 B.n45 10.6151
R1651 B.n873 B.n872 10.6151
R1652 B.n872 B.n871 10.6151
R1653 B.n871 B.n52 10.6151
R1654 B.n865 B.n52 10.6151
R1655 B.n865 B.n864 10.6151
R1656 B.n864 B.n863 10.6151
R1657 B.n863 B.n59 10.6151
R1658 B.n231 B.n230 9.36635
R1659 B.n253 B.n252 9.36635
R1660 B.n608 B.n481 9.36635
R1661 B.n585 B.n484 9.36635
R1662 B.t0 B.n389 3.62488
R1663 B.n773 B.t6 3.62488
R1664 B.t2 B.n370 3.62488
R1665 B.n804 B.t7 3.62488
R1666 B.n917 B.t4 3.62488
R1667 B.n908 B.t3 3.62488
R1668 B.n899 B.t5 3.62488
R1669 B.t1 B.n36 3.62488
R1670 B.n927 B.n0 2.81026
R1671 B.n927 B.n1 2.81026
R1672 B.n232 B.n231 1.24928
R1673 B.n252 B.n251 1.24928
R1674 B.n605 B.n481 1.24928
R1675 B.n588 B.n484 1.24928
R1676 VP.n11 VP.t0 311.577
R1677 VP.n5 VP.t7 280.933
R1678 VP.n29 VP.t4 280.933
R1679 VP.n36 VP.t3 280.933
R1680 VP.n43 VP.t5 280.933
R1681 VP.n23 VP.t6 280.933
R1682 VP.n16 VP.t1 280.933
R1683 VP.n10 VP.t2 280.933
R1684 VP.n25 VP.n5 171.088
R1685 VP.n44 VP.n43 171.088
R1686 VP.n24 VP.n23 171.088
R1687 VP.n12 VP.n9 161.3
R1688 VP.n14 VP.n13 161.3
R1689 VP.n15 VP.n8 161.3
R1690 VP.n18 VP.n17 161.3
R1691 VP.n19 VP.n7 161.3
R1692 VP.n21 VP.n20 161.3
R1693 VP.n22 VP.n6 161.3
R1694 VP.n42 VP.n0 161.3
R1695 VP.n41 VP.n40 161.3
R1696 VP.n39 VP.n1 161.3
R1697 VP.n38 VP.n37 161.3
R1698 VP.n35 VP.n2 161.3
R1699 VP.n34 VP.n33 161.3
R1700 VP.n32 VP.n3 161.3
R1701 VP.n31 VP.n30 161.3
R1702 VP.n28 VP.n4 161.3
R1703 VP.n27 VP.n26 161.3
R1704 VP.n11 VP.n10 60.1408
R1705 VP.n35 VP.n34 56.5193
R1706 VP.n15 VP.n14 56.5193
R1707 VP.n25 VP.n24 48.1141
R1708 VP.n30 VP.n28 45.3497
R1709 VP.n41 VP.n1 45.3497
R1710 VP.n21 VP.n7 45.3497
R1711 VP.n28 VP.n27 35.6371
R1712 VP.n42 VP.n41 35.6371
R1713 VP.n22 VP.n21 35.6371
R1714 VP.n12 VP.n11 26.7826
R1715 VP.n34 VP.n3 24.4675
R1716 VP.n37 VP.n35 24.4675
R1717 VP.n17 VP.n15 24.4675
R1718 VP.n14 VP.n9 24.4675
R1719 VP.n30 VP.n29 19.5741
R1720 VP.n36 VP.n1 19.5741
R1721 VP.n16 VP.n7 19.5741
R1722 VP.n27 VP.n5 14.6807
R1723 VP.n43 VP.n42 14.6807
R1724 VP.n23 VP.n22 14.6807
R1725 VP.n29 VP.n3 4.8939
R1726 VP.n37 VP.n36 4.8939
R1727 VP.n17 VP.n16 4.8939
R1728 VP.n10 VP.n9 4.8939
R1729 VP.n13 VP.n12 0.189894
R1730 VP.n13 VP.n8 0.189894
R1731 VP.n18 VP.n8 0.189894
R1732 VP.n19 VP.n18 0.189894
R1733 VP.n20 VP.n19 0.189894
R1734 VP.n20 VP.n6 0.189894
R1735 VP.n24 VP.n6 0.189894
R1736 VP.n26 VP.n25 0.189894
R1737 VP.n26 VP.n4 0.189894
R1738 VP.n31 VP.n4 0.189894
R1739 VP.n32 VP.n31 0.189894
R1740 VP.n33 VP.n32 0.189894
R1741 VP.n33 VP.n2 0.189894
R1742 VP.n38 VP.n2 0.189894
R1743 VP.n39 VP.n38 0.189894
R1744 VP.n40 VP.n39 0.189894
R1745 VP.n40 VP.n0 0.189894
R1746 VP.n44 VP.n0 0.189894
R1747 VP VP.n44 0.0516364
R1748 VDD1 VDD1.n0 59.8494
R1749 VDD1.n3 VDD1.n2 59.7357
R1750 VDD1.n3 VDD1.n1 59.7357
R1751 VDD1.n5 VDD1.n4 59.0585
R1752 VDD1.n5 VDD1.n3 44.6604
R1753 VDD1.n4 VDD1.t6 1.24032
R1754 VDD1.n4 VDD1.t1 1.24032
R1755 VDD1.n0 VDD1.t7 1.24032
R1756 VDD1.n0 VDD1.t5 1.24032
R1757 VDD1.n2 VDD1.t4 1.24032
R1758 VDD1.n2 VDD1.t2 1.24032
R1759 VDD1.n1 VDD1.t0 1.24032
R1760 VDD1.n1 VDD1.t3 1.24032
R1761 VDD1 VDD1.n5 0.675069
C0 VP VDD2 0.388426f
C1 VN VP 6.8921f
C2 VDD2 VDD1 1.16031f
C3 VN VDD1 0.149144f
C4 VTAIL VDD2 10.647f
C5 VN VTAIL 9.47736f
C6 VP VDD1 9.88068f
C7 VN VDD2 9.64217f
C8 VTAIL VP 9.49147f
C9 VTAIL VDD1 10.6008f
C10 VDD2 B 4.445672f
C11 VDD1 B 4.752871f
C12 VTAIL B 11.848832f
C13 VN B 11.30362f
C14 VP B 9.521993f
C15 VDD1.t7 B 0.320061f
C16 VDD1.t5 B 0.320061f
C17 VDD1.n0 B 2.89764f
C18 VDD1.t0 B 0.320061f
C19 VDD1.t3 B 0.320061f
C20 VDD1.n1 B 2.89677f
C21 VDD1.t4 B 0.320061f
C22 VDD1.t2 B 0.320061f
C23 VDD1.n2 B 2.89677f
C24 VDD1.n3 B 2.92184f
C25 VDD1.t6 B 0.320061f
C26 VDD1.t1 B 0.320061f
C27 VDD1.n4 B 2.89219f
C28 VDD1.n5 B 2.90761f
C29 VP.n0 B 0.032348f
C30 VP.t5 B 1.94204f
C31 VP.n1 B 0.056253f
C32 VP.n2 B 0.032348f
C33 VP.n3 B 0.036477f
C34 VP.n4 B 0.032348f
C35 VP.t7 B 1.94204f
C36 VP.n5 B 0.757294f
C37 VP.n6 B 0.032348f
C38 VP.t6 B 1.94204f
C39 VP.n7 B 0.056253f
C40 VP.n8 B 0.032348f
C41 VP.n9 B 0.036477f
C42 VP.t0 B 2.02078f
C43 VP.t2 B 1.94204f
C44 VP.n10 B 0.737245f
C45 VP.n11 B 0.770793f
C46 VP.n12 B 0.173445f
C47 VP.n13 B 0.032348f
C48 VP.n14 B 0.047223f
C49 VP.n15 B 0.047223f
C50 VP.t1 B 1.94204f
C51 VP.n16 B 0.690912f
C52 VP.n17 B 0.036477f
C53 VP.n18 B 0.032348f
C54 VP.n19 B 0.032348f
C55 VP.n20 B 0.032348f
C56 VP.n21 B 0.027205f
C57 VP.n22 B 0.053419f
C58 VP.n23 B 0.757294f
C59 VP.n24 B 1.66295f
C60 VP.n25 B 1.68712f
C61 VP.n26 B 0.032348f
C62 VP.n27 B 0.053419f
C63 VP.n28 B 0.027205f
C64 VP.t4 B 1.94204f
C65 VP.n29 B 0.690912f
C66 VP.n30 B 0.056253f
C67 VP.n31 B 0.032348f
C68 VP.n32 B 0.032348f
C69 VP.n33 B 0.032348f
C70 VP.n34 B 0.047223f
C71 VP.n35 B 0.047223f
C72 VP.t3 B 1.94204f
C73 VP.n36 B 0.690912f
C74 VP.n37 B 0.036477f
C75 VP.n38 B 0.032348f
C76 VP.n39 B 0.032348f
C77 VP.n40 B 0.032348f
C78 VP.n41 B 0.027205f
C79 VP.n42 B 0.053419f
C80 VP.n43 B 0.757294f
C81 VP.n44 B 0.029097f
C82 VDD2.t0 B 0.316825f
C83 VDD2.t1 B 0.316825f
C84 VDD2.n0 B 2.86748f
C85 VDD2.t5 B 0.316825f
C86 VDD2.t4 B 0.316825f
C87 VDD2.n1 B 2.86748f
C88 VDD2.n2 B 2.83943f
C89 VDD2.t6 B 0.316825f
C90 VDD2.t7 B 0.316825f
C91 VDD2.n3 B 2.86295f
C92 VDD2.n4 B 2.84776f
C93 VDD2.t2 B 0.316825f
C94 VDD2.t3 B 0.316825f
C95 VDD2.n5 B 2.86745f
C96 VTAIL.t14 B 0.234461f
C97 VTAIL.t15 B 0.234461f
C98 VTAIL.n0 B 2.05728f
C99 VTAIL.n1 B 0.286894f
C100 VTAIL.t13 B 2.62673f
C101 VTAIL.n2 B 0.381524f
C102 VTAIL.t7 B 2.62673f
C103 VTAIL.n3 B 0.381524f
C104 VTAIL.t6 B 0.234461f
C105 VTAIL.t2 B 0.234461f
C106 VTAIL.n4 B 2.05728f
C107 VTAIL.n5 B 0.371143f
C108 VTAIL.t0 B 2.62673f
C109 VTAIL.n6 B 1.51767f
C110 VTAIL.t10 B 2.62674f
C111 VTAIL.n7 B 1.51766f
C112 VTAIL.t12 B 0.234461f
C113 VTAIL.t11 B 0.234461f
C114 VTAIL.n8 B 2.05729f
C115 VTAIL.n9 B 0.371136f
C116 VTAIL.t9 B 2.62674f
C117 VTAIL.n10 B 0.381517f
C118 VTAIL.t4 B 2.62674f
C119 VTAIL.n11 B 0.381517f
C120 VTAIL.t3 B 0.234461f
C121 VTAIL.t5 B 0.234461f
C122 VTAIL.n12 B 2.05729f
C123 VTAIL.n13 B 0.371136f
C124 VTAIL.t1 B 2.62674f
C125 VTAIL.n14 B 1.51766f
C126 VTAIL.t8 B 2.62673f
C127 VTAIL.n15 B 1.51418f
C128 VN.n0 B 0.031924f
C129 VN.t3 B 1.91657f
C130 VN.n1 B 0.055515f
C131 VN.n2 B 0.031924f
C132 VN.n3 B 0.035999f
C133 VN.t7 B 1.99428f
C134 VN.t6 B 1.91657f
C135 VN.n4 B 0.727578f
C136 VN.n5 B 0.760686f
C137 VN.n6 B 0.17117f
C138 VN.n7 B 0.031924f
C139 VN.n8 B 0.046604f
C140 VN.n9 B 0.046604f
C141 VN.t2 B 1.91657f
C142 VN.n10 B 0.681852f
C143 VN.n11 B 0.035999f
C144 VN.n12 B 0.031924f
C145 VN.n13 B 0.031924f
C146 VN.n14 B 0.031924f
C147 VN.n15 B 0.026848f
C148 VN.n16 B 0.052718f
C149 VN.n17 B 0.747363f
C150 VN.n18 B 0.028715f
C151 VN.n19 B 0.031924f
C152 VN.t1 B 1.91657f
C153 VN.n20 B 0.055515f
C154 VN.n21 B 0.031924f
C155 VN.t0 B 1.91657f
C156 VN.n22 B 0.681852f
C157 VN.n23 B 0.035999f
C158 VN.t4 B 1.99428f
C159 VN.t5 B 1.91657f
C160 VN.n24 B 0.727578f
C161 VN.n25 B 0.760686f
C162 VN.n26 B 0.17117f
C163 VN.n27 B 0.031924f
C164 VN.n28 B 0.046604f
C165 VN.n29 B 0.046604f
C166 VN.n30 B 0.035999f
C167 VN.n31 B 0.031924f
C168 VN.n32 B 0.031924f
C169 VN.n33 B 0.031924f
C170 VN.n34 B 0.026848f
C171 VN.n35 B 0.052718f
C172 VN.n36 B 0.747363f
C173 VN.n37 B 1.66194f
.ends

