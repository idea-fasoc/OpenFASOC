* NGSPICE file created from diff_pair_sample_1051.ext - technology: sky130A

.subckt diff_pair_sample_1051 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t19 VP.t0 VDD1.t7 B.t9 sky130_fd_pr__nfet_01v8 ad=0.3597 pd=2.51 as=0.3597 ps=2.51 w=2.18 l=3.39
X1 VDD2.t9 VN.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.8502 pd=5.14 as=0.3597 ps=2.51 w=2.18 l=3.39
X2 VTAIL.t18 VP.t1 VDD1.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.3597 pd=2.51 as=0.3597 ps=2.51 w=2.18 l=3.39
X3 VDD1.t3 VP.t2 VTAIL.t17 B.t0 sky130_fd_pr__nfet_01v8 ad=0.3597 pd=2.51 as=0.8502 ps=5.14 w=2.18 l=3.39
X4 VDD2.t8 VN.t1 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.3597 pd=2.51 as=0.3597 ps=2.51 w=2.18 l=3.39
X5 VTAIL.t16 VP.t3 VDD1.t9 B.t4 sky130_fd_pr__nfet_01v8 ad=0.3597 pd=2.51 as=0.3597 ps=2.51 w=2.18 l=3.39
X6 VTAIL.t4 VN.t2 VDD2.t7 B.t4 sky130_fd_pr__nfet_01v8 ad=0.3597 pd=2.51 as=0.3597 ps=2.51 w=2.18 l=3.39
X7 VDD1.t0 VP.t4 VTAIL.t15 B.t3 sky130_fd_pr__nfet_01v8 ad=0.3597 pd=2.51 as=0.3597 ps=2.51 w=2.18 l=3.39
X8 B.t23 B.t21 B.t22 B.t18 sky130_fd_pr__nfet_01v8 ad=0.8502 pd=5.14 as=0 ps=0 w=2.18 l=3.39
X9 VDD2.t6 VN.t3 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=0.8502 pd=5.14 as=0.3597 ps=2.51 w=2.18 l=3.39
X10 VTAIL.t8 VN.t4 VDD2.t5 B.t8 sky130_fd_pr__nfet_01v8 ad=0.3597 pd=2.51 as=0.3597 ps=2.51 w=2.18 l=3.39
X11 VDD1.t6 VP.t5 VTAIL.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=0.3597 pd=2.51 as=0.8502 ps=5.14 w=2.18 l=3.39
X12 VDD1.t8 VP.t6 VTAIL.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=0.8502 pd=5.14 as=0.3597 ps=2.51 w=2.18 l=3.39
X13 VDD2.t4 VN.t5 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.3597 pd=2.51 as=0.8502 ps=5.14 w=2.18 l=3.39
X14 VTAIL.t9 VN.t6 VDD2.t3 B.t9 sky130_fd_pr__nfet_01v8 ad=0.3597 pd=2.51 as=0.3597 ps=2.51 w=2.18 l=3.39
X15 VTAIL.t12 VP.t7 VDD1.t5 B.t8 sky130_fd_pr__nfet_01v8 ad=0.3597 pd=2.51 as=0.3597 ps=2.51 w=2.18 l=3.39
X16 VDD1.t4 VP.t8 VTAIL.t11 B.t6 sky130_fd_pr__nfet_01v8 ad=0.3597 pd=2.51 as=0.3597 ps=2.51 w=2.18 l=3.39
X17 B.t20 B.t17 B.t19 B.t18 sky130_fd_pr__nfet_01v8 ad=0.8502 pd=5.14 as=0 ps=0 w=2.18 l=3.39
X18 VDD2.t2 VN.t7 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=0.3597 pd=2.51 as=0.8502 ps=5.14 w=2.18 l=3.39
X19 VTAIL.t2 VN.t8 VDD2.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=0.3597 pd=2.51 as=0.3597 ps=2.51 w=2.18 l=3.39
X20 VDD1.t1 VP.t9 VTAIL.t10 B.t1 sky130_fd_pr__nfet_01v8 ad=0.8502 pd=5.14 as=0.3597 ps=2.51 w=2.18 l=3.39
X21 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=0.8502 pd=5.14 as=0 ps=0 w=2.18 l=3.39
X22 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=0.8502 pd=5.14 as=0 ps=0 w=2.18 l=3.39
X23 VDD2.t0 VN.t9 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=0.3597 pd=2.51 as=0.3597 ps=2.51 w=2.18 l=3.39
R0 VP.n32 VP.n31 161.3
R1 VP.n33 VP.n28 161.3
R2 VP.n35 VP.n34 161.3
R3 VP.n36 VP.n27 161.3
R4 VP.n38 VP.n37 161.3
R5 VP.n39 VP.n26 161.3
R6 VP.n41 VP.n40 161.3
R7 VP.n43 VP.n42 161.3
R8 VP.n44 VP.n24 161.3
R9 VP.n46 VP.n45 161.3
R10 VP.n47 VP.n23 161.3
R11 VP.n49 VP.n48 161.3
R12 VP.n50 VP.n22 161.3
R13 VP.n53 VP.n52 161.3
R14 VP.n54 VP.n21 161.3
R15 VP.n56 VP.n55 161.3
R16 VP.n57 VP.n20 161.3
R17 VP.n59 VP.n58 161.3
R18 VP.n60 VP.n19 161.3
R19 VP.n62 VP.n61 161.3
R20 VP.n63 VP.n18 161.3
R21 VP.n65 VP.n64 161.3
R22 VP.n115 VP.n114 161.3
R23 VP.n113 VP.n1 161.3
R24 VP.n112 VP.n111 161.3
R25 VP.n110 VP.n2 161.3
R26 VP.n109 VP.n108 161.3
R27 VP.n107 VP.n3 161.3
R28 VP.n106 VP.n105 161.3
R29 VP.n104 VP.n4 161.3
R30 VP.n103 VP.n102 161.3
R31 VP.n100 VP.n5 161.3
R32 VP.n99 VP.n98 161.3
R33 VP.n97 VP.n6 161.3
R34 VP.n96 VP.n95 161.3
R35 VP.n94 VP.n7 161.3
R36 VP.n93 VP.n92 161.3
R37 VP.n91 VP.n90 161.3
R38 VP.n89 VP.n9 161.3
R39 VP.n88 VP.n87 161.3
R40 VP.n86 VP.n10 161.3
R41 VP.n85 VP.n84 161.3
R42 VP.n83 VP.n11 161.3
R43 VP.n82 VP.n81 161.3
R44 VP.n80 VP.n79 161.3
R45 VP.n78 VP.n13 161.3
R46 VP.n77 VP.n76 161.3
R47 VP.n75 VP.n14 161.3
R48 VP.n74 VP.n73 161.3
R49 VP.n72 VP.n15 161.3
R50 VP.n71 VP.n70 161.3
R51 VP.n69 VP.n16 161.3
R52 VP.n68 VP.n67 80.6405
R53 VP.n116 VP.n0 80.6405
R54 VP.n66 VP.n17 80.6405
R55 VP.n73 VP.n14 56.4773
R56 VP.n108 VP.n2 56.4773
R57 VP.n58 VP.n19 56.4773
R58 VP.n30 VP.n29 51.4682
R59 VP.n84 VP.n10 51.1217
R60 VP.n99 VP.n6 51.1217
R61 VP.n49 VP.n23 51.1217
R62 VP.n34 VP.n27 51.1217
R63 VP.n68 VP.n66 50.0218
R64 VP.n30 VP.t6 48.6972
R65 VP.n88 VP.n10 29.6995
R66 VP.n95 VP.n6 29.6995
R67 VP.n45 VP.n23 29.6995
R68 VP.n38 VP.n27 29.6995
R69 VP.n71 VP.n16 24.3439
R70 VP.n72 VP.n71 24.3439
R71 VP.n73 VP.n72 24.3439
R72 VP.n77 VP.n14 24.3439
R73 VP.n78 VP.n77 24.3439
R74 VP.n79 VP.n78 24.3439
R75 VP.n83 VP.n82 24.3439
R76 VP.n84 VP.n83 24.3439
R77 VP.n89 VP.n88 24.3439
R78 VP.n90 VP.n89 24.3439
R79 VP.n94 VP.n93 24.3439
R80 VP.n95 VP.n94 24.3439
R81 VP.n100 VP.n99 24.3439
R82 VP.n102 VP.n100 24.3439
R83 VP.n106 VP.n4 24.3439
R84 VP.n107 VP.n106 24.3439
R85 VP.n108 VP.n107 24.3439
R86 VP.n112 VP.n2 24.3439
R87 VP.n113 VP.n112 24.3439
R88 VP.n114 VP.n113 24.3439
R89 VP.n62 VP.n19 24.3439
R90 VP.n63 VP.n62 24.3439
R91 VP.n64 VP.n63 24.3439
R92 VP.n50 VP.n49 24.3439
R93 VP.n52 VP.n50 24.3439
R94 VP.n56 VP.n21 24.3439
R95 VP.n57 VP.n56 24.3439
R96 VP.n58 VP.n57 24.3439
R97 VP.n39 VP.n38 24.3439
R98 VP.n40 VP.n39 24.3439
R99 VP.n44 VP.n43 24.3439
R100 VP.n45 VP.n44 24.3439
R101 VP.n33 VP.n32 24.3439
R102 VP.n34 VP.n33 24.3439
R103 VP.n82 VP.n12 22.8833
R104 VP.n102 VP.n101 22.8833
R105 VP.n52 VP.n51 22.8833
R106 VP.n32 VP.n29 22.8833
R107 VP.n67 VP.t9 15.4984
R108 VP.n12 VP.t7 15.4984
R109 VP.n8 VP.t4 15.4984
R110 VP.n101 VP.t3 15.4984
R111 VP.n0 VP.t2 15.4984
R112 VP.n17 VP.t5 15.4984
R113 VP.n51 VP.t0 15.4984
R114 VP.n25 VP.t8 15.4984
R115 VP.n29 VP.t1 15.4984
R116 VP.n90 VP.n8 12.1722
R117 VP.n93 VP.n8 12.1722
R118 VP.n40 VP.n25 12.1722
R119 VP.n43 VP.n25 12.1722
R120 VP.n67 VP.n16 9.251
R121 VP.n114 VP.n0 9.251
R122 VP.n64 VP.n17 9.251
R123 VP.n31 VP.n30 3.19273
R124 VP.n79 VP.n12 1.46111
R125 VP.n101 VP.n4 1.46111
R126 VP.n51 VP.n21 1.46111
R127 VP.n66 VP.n65 0.355081
R128 VP.n69 VP.n68 0.355081
R129 VP.n116 VP.n115 0.355081
R130 VP VP.n116 0.26685
R131 VP.n31 VP.n28 0.189894
R132 VP.n35 VP.n28 0.189894
R133 VP.n36 VP.n35 0.189894
R134 VP.n37 VP.n36 0.189894
R135 VP.n37 VP.n26 0.189894
R136 VP.n41 VP.n26 0.189894
R137 VP.n42 VP.n41 0.189894
R138 VP.n42 VP.n24 0.189894
R139 VP.n46 VP.n24 0.189894
R140 VP.n47 VP.n46 0.189894
R141 VP.n48 VP.n47 0.189894
R142 VP.n48 VP.n22 0.189894
R143 VP.n53 VP.n22 0.189894
R144 VP.n54 VP.n53 0.189894
R145 VP.n55 VP.n54 0.189894
R146 VP.n55 VP.n20 0.189894
R147 VP.n59 VP.n20 0.189894
R148 VP.n60 VP.n59 0.189894
R149 VP.n61 VP.n60 0.189894
R150 VP.n61 VP.n18 0.189894
R151 VP.n65 VP.n18 0.189894
R152 VP.n70 VP.n69 0.189894
R153 VP.n70 VP.n15 0.189894
R154 VP.n74 VP.n15 0.189894
R155 VP.n75 VP.n74 0.189894
R156 VP.n76 VP.n75 0.189894
R157 VP.n76 VP.n13 0.189894
R158 VP.n80 VP.n13 0.189894
R159 VP.n81 VP.n80 0.189894
R160 VP.n81 VP.n11 0.189894
R161 VP.n85 VP.n11 0.189894
R162 VP.n86 VP.n85 0.189894
R163 VP.n87 VP.n86 0.189894
R164 VP.n87 VP.n9 0.189894
R165 VP.n91 VP.n9 0.189894
R166 VP.n92 VP.n91 0.189894
R167 VP.n92 VP.n7 0.189894
R168 VP.n96 VP.n7 0.189894
R169 VP.n97 VP.n96 0.189894
R170 VP.n98 VP.n97 0.189894
R171 VP.n98 VP.n5 0.189894
R172 VP.n103 VP.n5 0.189894
R173 VP.n104 VP.n103 0.189894
R174 VP.n105 VP.n104 0.189894
R175 VP.n105 VP.n3 0.189894
R176 VP.n109 VP.n3 0.189894
R177 VP.n110 VP.n109 0.189894
R178 VP.n111 VP.n110 0.189894
R179 VP.n111 VP.n1 0.189894
R180 VP.n115 VP.n1 0.189894
R181 VDD1.n3 VDD1.t1 105.757
R182 VDD1.n1 VDD1.t8 105.757
R183 VDD1.n5 VDD1.n4 95.8172
R184 VDD1.n1 VDD1.n0 93.4677
R185 VDD1.n7 VDD1.n6 93.4676
R186 VDD1.n3 VDD1.n2 93.4674
R187 VDD1.n7 VDD1.n5 43.0138
R188 VDD1.n6 VDD1.t7 9.08307
R189 VDD1.n6 VDD1.t6 9.08307
R190 VDD1.n0 VDD1.t2 9.08307
R191 VDD1.n0 VDD1.t4 9.08307
R192 VDD1.n4 VDD1.t9 9.08307
R193 VDD1.n4 VDD1.t3 9.08307
R194 VDD1.n2 VDD1.t5 9.08307
R195 VDD1.n2 VDD1.t0 9.08307
R196 VDD1 VDD1.n7 2.34748
R197 VDD1 VDD1.n1 0.860414
R198 VDD1.n5 VDD1.n3 0.746878
R199 VTAIL.n17 VTAIL.t7 85.8714
R200 VTAIL.n2 VTAIL.t17 85.8714
R201 VTAIL.n16 VTAIL.t14 85.8714
R202 VTAIL.n11 VTAIL.t0 85.8713
R203 VTAIL.n15 VTAIL.n14 76.7889
R204 VTAIL.n13 VTAIL.n12 76.7889
R205 VTAIL.n10 VTAIL.n9 76.7889
R206 VTAIL.n8 VTAIL.n7 76.7889
R207 VTAIL.n19 VTAIL.n18 76.7886
R208 VTAIL.n1 VTAIL.n0 76.7886
R209 VTAIL.n4 VTAIL.n3 76.7886
R210 VTAIL.n6 VTAIL.n5 76.7886
R211 VTAIL.n8 VTAIL.n6 20.66
R212 VTAIL.n17 VTAIL.n16 17.4531
R213 VTAIL.n18 VTAIL.t6 9.08307
R214 VTAIL.n18 VTAIL.t9 9.08307
R215 VTAIL.n0 VTAIL.t5 9.08307
R216 VTAIL.n0 VTAIL.t2 9.08307
R217 VTAIL.n3 VTAIL.t15 9.08307
R218 VTAIL.n3 VTAIL.t16 9.08307
R219 VTAIL.n5 VTAIL.t10 9.08307
R220 VTAIL.n5 VTAIL.t12 9.08307
R221 VTAIL.n14 VTAIL.t11 9.08307
R222 VTAIL.n14 VTAIL.t19 9.08307
R223 VTAIL.n12 VTAIL.t13 9.08307
R224 VTAIL.n12 VTAIL.t18 9.08307
R225 VTAIL.n9 VTAIL.t3 9.08307
R226 VTAIL.n9 VTAIL.t4 9.08307
R227 VTAIL.n7 VTAIL.t1 9.08307
R228 VTAIL.n7 VTAIL.t8 9.08307
R229 VTAIL.n10 VTAIL.n8 3.2074
R230 VTAIL.n11 VTAIL.n10 3.2074
R231 VTAIL.n15 VTAIL.n13 3.2074
R232 VTAIL.n16 VTAIL.n15 3.2074
R233 VTAIL.n6 VTAIL.n4 3.2074
R234 VTAIL.n4 VTAIL.n2 3.2074
R235 VTAIL.n19 VTAIL.n17 3.2074
R236 VTAIL VTAIL.n1 2.46386
R237 VTAIL.n13 VTAIL.n11 2.07378
R238 VTAIL.n2 VTAIL.n1 2.07378
R239 VTAIL VTAIL.n19 0.744035
R240 B.n776 B.n775 585
R241 B.n777 B.n776 585
R242 B.n224 B.n151 585
R243 B.n223 B.n222 585
R244 B.n221 B.n220 585
R245 B.n219 B.n218 585
R246 B.n217 B.n216 585
R247 B.n215 B.n214 585
R248 B.n213 B.n212 585
R249 B.n211 B.n210 585
R250 B.n209 B.n208 585
R251 B.n207 B.n206 585
R252 B.n205 B.n204 585
R253 B.n203 B.n202 585
R254 B.n201 B.n200 585
R255 B.n199 B.n198 585
R256 B.n197 B.n196 585
R257 B.n195 B.n194 585
R258 B.n193 B.n192 585
R259 B.n191 B.n190 585
R260 B.n189 B.n188 585
R261 B.n187 B.n186 585
R262 B.n185 B.n184 585
R263 B.n182 B.n181 585
R264 B.n180 B.n179 585
R265 B.n178 B.n177 585
R266 B.n176 B.n175 585
R267 B.n174 B.n173 585
R268 B.n172 B.n171 585
R269 B.n170 B.n169 585
R270 B.n168 B.n167 585
R271 B.n166 B.n165 585
R272 B.n164 B.n163 585
R273 B.n162 B.n161 585
R274 B.n160 B.n159 585
R275 B.n158 B.n157 585
R276 B.n774 B.n133 585
R277 B.n778 B.n133 585
R278 B.n773 B.n132 585
R279 B.n779 B.n132 585
R280 B.n772 B.n771 585
R281 B.n771 B.n128 585
R282 B.n770 B.n127 585
R283 B.n785 B.n127 585
R284 B.n769 B.n126 585
R285 B.n786 B.n126 585
R286 B.n768 B.n125 585
R287 B.n787 B.n125 585
R288 B.n767 B.n766 585
R289 B.n766 B.n121 585
R290 B.n765 B.n120 585
R291 B.n793 B.n120 585
R292 B.n764 B.n119 585
R293 B.n794 B.n119 585
R294 B.n763 B.n118 585
R295 B.n795 B.n118 585
R296 B.n762 B.n761 585
R297 B.n761 B.n114 585
R298 B.n760 B.n113 585
R299 B.n801 B.n113 585
R300 B.n759 B.n112 585
R301 B.n802 B.n112 585
R302 B.n758 B.n111 585
R303 B.n803 B.n111 585
R304 B.n757 B.n756 585
R305 B.n756 B.n107 585
R306 B.n755 B.n106 585
R307 B.n809 B.n106 585
R308 B.n754 B.n105 585
R309 B.n810 B.n105 585
R310 B.n753 B.n104 585
R311 B.n811 B.n104 585
R312 B.n752 B.n751 585
R313 B.n751 B.n100 585
R314 B.n750 B.n99 585
R315 B.n817 B.n99 585
R316 B.n749 B.n98 585
R317 B.n818 B.n98 585
R318 B.n748 B.n97 585
R319 B.n819 B.n97 585
R320 B.n747 B.n746 585
R321 B.n746 B.n96 585
R322 B.n745 B.n92 585
R323 B.n825 B.n92 585
R324 B.n744 B.n91 585
R325 B.n826 B.n91 585
R326 B.n743 B.n90 585
R327 B.n827 B.n90 585
R328 B.n742 B.n741 585
R329 B.n741 B.n86 585
R330 B.n740 B.n85 585
R331 B.n833 B.n85 585
R332 B.n739 B.n84 585
R333 B.n834 B.n84 585
R334 B.n738 B.n83 585
R335 B.n835 B.n83 585
R336 B.n737 B.n736 585
R337 B.n736 B.n79 585
R338 B.n735 B.n78 585
R339 B.n841 B.n78 585
R340 B.n734 B.n77 585
R341 B.n842 B.n77 585
R342 B.n733 B.n76 585
R343 B.n843 B.n76 585
R344 B.n732 B.n731 585
R345 B.n731 B.n72 585
R346 B.n730 B.n71 585
R347 B.n849 B.n71 585
R348 B.n729 B.n70 585
R349 B.n850 B.n70 585
R350 B.n728 B.n69 585
R351 B.n851 B.n69 585
R352 B.n727 B.n726 585
R353 B.n726 B.n65 585
R354 B.n725 B.n64 585
R355 B.n857 B.n64 585
R356 B.n724 B.n63 585
R357 B.n858 B.n63 585
R358 B.n723 B.n62 585
R359 B.n859 B.n62 585
R360 B.n722 B.n721 585
R361 B.n721 B.n58 585
R362 B.n720 B.n57 585
R363 B.n865 B.n57 585
R364 B.n719 B.n56 585
R365 B.n866 B.n56 585
R366 B.n718 B.n55 585
R367 B.n867 B.n55 585
R368 B.n717 B.n716 585
R369 B.n716 B.n51 585
R370 B.n715 B.n50 585
R371 B.n873 B.n50 585
R372 B.n714 B.n49 585
R373 B.n874 B.n49 585
R374 B.n713 B.n48 585
R375 B.n875 B.n48 585
R376 B.n712 B.n711 585
R377 B.n711 B.n44 585
R378 B.n710 B.n43 585
R379 B.n881 B.n43 585
R380 B.n709 B.n42 585
R381 B.n882 B.n42 585
R382 B.n708 B.n41 585
R383 B.n883 B.n41 585
R384 B.n707 B.n706 585
R385 B.n706 B.n37 585
R386 B.n705 B.n36 585
R387 B.n889 B.n36 585
R388 B.n704 B.n35 585
R389 B.n890 B.n35 585
R390 B.n703 B.n34 585
R391 B.n891 B.n34 585
R392 B.n702 B.n701 585
R393 B.n701 B.n30 585
R394 B.n700 B.n29 585
R395 B.n897 B.n29 585
R396 B.n699 B.n28 585
R397 B.n898 B.n28 585
R398 B.n698 B.n27 585
R399 B.n899 B.n27 585
R400 B.n697 B.n696 585
R401 B.n696 B.n23 585
R402 B.n695 B.n22 585
R403 B.n905 B.n22 585
R404 B.n694 B.n21 585
R405 B.n906 B.n21 585
R406 B.n693 B.n20 585
R407 B.n907 B.n20 585
R408 B.n692 B.n691 585
R409 B.n691 B.n19 585
R410 B.n690 B.n15 585
R411 B.n913 B.n15 585
R412 B.n689 B.n14 585
R413 B.n914 B.n14 585
R414 B.n688 B.n13 585
R415 B.n915 B.n13 585
R416 B.n687 B.n686 585
R417 B.n686 B.n12 585
R418 B.n685 B.n684 585
R419 B.n685 B.n8 585
R420 B.n683 B.n7 585
R421 B.n922 B.n7 585
R422 B.n682 B.n6 585
R423 B.n923 B.n6 585
R424 B.n681 B.n5 585
R425 B.n924 B.n5 585
R426 B.n680 B.n679 585
R427 B.n679 B.n4 585
R428 B.n678 B.n225 585
R429 B.n678 B.n677 585
R430 B.n668 B.n226 585
R431 B.n227 B.n226 585
R432 B.n670 B.n669 585
R433 B.n671 B.n670 585
R434 B.n667 B.n232 585
R435 B.n232 B.n231 585
R436 B.n666 B.n665 585
R437 B.n665 B.n664 585
R438 B.n234 B.n233 585
R439 B.n657 B.n234 585
R440 B.n656 B.n655 585
R441 B.n658 B.n656 585
R442 B.n654 B.n239 585
R443 B.n239 B.n238 585
R444 B.n653 B.n652 585
R445 B.n652 B.n651 585
R446 B.n241 B.n240 585
R447 B.n242 B.n241 585
R448 B.n644 B.n643 585
R449 B.n645 B.n644 585
R450 B.n642 B.n247 585
R451 B.n247 B.n246 585
R452 B.n641 B.n640 585
R453 B.n640 B.n639 585
R454 B.n249 B.n248 585
R455 B.n250 B.n249 585
R456 B.n632 B.n631 585
R457 B.n633 B.n632 585
R458 B.n630 B.n255 585
R459 B.n255 B.n254 585
R460 B.n629 B.n628 585
R461 B.n628 B.n627 585
R462 B.n257 B.n256 585
R463 B.n258 B.n257 585
R464 B.n620 B.n619 585
R465 B.n621 B.n620 585
R466 B.n618 B.n263 585
R467 B.n263 B.n262 585
R468 B.n617 B.n616 585
R469 B.n616 B.n615 585
R470 B.n265 B.n264 585
R471 B.n266 B.n265 585
R472 B.n608 B.n607 585
R473 B.n609 B.n608 585
R474 B.n606 B.n271 585
R475 B.n271 B.n270 585
R476 B.n605 B.n604 585
R477 B.n604 B.n603 585
R478 B.n273 B.n272 585
R479 B.n274 B.n273 585
R480 B.n596 B.n595 585
R481 B.n597 B.n596 585
R482 B.n594 B.n278 585
R483 B.n282 B.n278 585
R484 B.n593 B.n592 585
R485 B.n592 B.n591 585
R486 B.n280 B.n279 585
R487 B.n281 B.n280 585
R488 B.n584 B.n583 585
R489 B.n585 B.n584 585
R490 B.n582 B.n287 585
R491 B.n287 B.n286 585
R492 B.n581 B.n580 585
R493 B.n580 B.n579 585
R494 B.n289 B.n288 585
R495 B.n290 B.n289 585
R496 B.n572 B.n571 585
R497 B.n573 B.n572 585
R498 B.n570 B.n295 585
R499 B.n295 B.n294 585
R500 B.n569 B.n568 585
R501 B.n568 B.n567 585
R502 B.n297 B.n296 585
R503 B.n298 B.n297 585
R504 B.n560 B.n559 585
R505 B.n561 B.n560 585
R506 B.n558 B.n303 585
R507 B.n303 B.n302 585
R508 B.n557 B.n556 585
R509 B.n556 B.n555 585
R510 B.n305 B.n304 585
R511 B.n306 B.n305 585
R512 B.n548 B.n547 585
R513 B.n549 B.n548 585
R514 B.n546 B.n311 585
R515 B.n311 B.n310 585
R516 B.n545 B.n544 585
R517 B.n544 B.n543 585
R518 B.n313 B.n312 585
R519 B.n314 B.n313 585
R520 B.n536 B.n535 585
R521 B.n537 B.n536 585
R522 B.n534 B.n319 585
R523 B.n319 B.n318 585
R524 B.n533 B.n532 585
R525 B.n532 B.n531 585
R526 B.n321 B.n320 585
R527 B.n524 B.n321 585
R528 B.n523 B.n522 585
R529 B.n525 B.n523 585
R530 B.n521 B.n326 585
R531 B.n326 B.n325 585
R532 B.n520 B.n519 585
R533 B.n519 B.n518 585
R534 B.n328 B.n327 585
R535 B.n329 B.n328 585
R536 B.n511 B.n510 585
R537 B.n512 B.n511 585
R538 B.n509 B.n334 585
R539 B.n334 B.n333 585
R540 B.n508 B.n507 585
R541 B.n507 B.n506 585
R542 B.n336 B.n335 585
R543 B.n337 B.n336 585
R544 B.n499 B.n498 585
R545 B.n500 B.n499 585
R546 B.n497 B.n342 585
R547 B.n342 B.n341 585
R548 B.n496 B.n495 585
R549 B.n495 B.n494 585
R550 B.n344 B.n343 585
R551 B.n345 B.n344 585
R552 B.n487 B.n486 585
R553 B.n488 B.n487 585
R554 B.n485 B.n349 585
R555 B.n353 B.n349 585
R556 B.n484 B.n483 585
R557 B.n483 B.n482 585
R558 B.n351 B.n350 585
R559 B.n352 B.n351 585
R560 B.n475 B.n474 585
R561 B.n476 B.n475 585
R562 B.n473 B.n358 585
R563 B.n358 B.n357 585
R564 B.n472 B.n471 585
R565 B.n471 B.n470 585
R566 B.n360 B.n359 585
R567 B.n361 B.n360 585
R568 B.n463 B.n462 585
R569 B.n464 B.n463 585
R570 B.n461 B.n366 585
R571 B.n366 B.n365 585
R572 B.n455 B.n454 585
R573 B.n453 B.n385 585
R574 B.n452 B.n384 585
R575 B.n457 B.n384 585
R576 B.n451 B.n450 585
R577 B.n449 B.n448 585
R578 B.n447 B.n446 585
R579 B.n445 B.n444 585
R580 B.n443 B.n442 585
R581 B.n441 B.n440 585
R582 B.n439 B.n438 585
R583 B.n437 B.n436 585
R584 B.n435 B.n434 585
R585 B.n433 B.n432 585
R586 B.n431 B.n430 585
R587 B.n429 B.n428 585
R588 B.n427 B.n426 585
R589 B.n425 B.n424 585
R590 B.n423 B.n422 585
R591 B.n421 B.n420 585
R592 B.n419 B.n418 585
R593 B.n417 B.n416 585
R594 B.n415 B.n414 585
R595 B.n412 B.n411 585
R596 B.n410 B.n409 585
R597 B.n408 B.n407 585
R598 B.n406 B.n405 585
R599 B.n404 B.n403 585
R600 B.n402 B.n401 585
R601 B.n400 B.n399 585
R602 B.n398 B.n397 585
R603 B.n396 B.n395 585
R604 B.n394 B.n393 585
R605 B.n392 B.n391 585
R606 B.n368 B.n367 585
R607 B.n460 B.n459 585
R608 B.n364 B.n363 585
R609 B.n365 B.n364 585
R610 B.n466 B.n465 585
R611 B.n465 B.n464 585
R612 B.n467 B.n362 585
R613 B.n362 B.n361 585
R614 B.n469 B.n468 585
R615 B.n470 B.n469 585
R616 B.n356 B.n355 585
R617 B.n357 B.n356 585
R618 B.n478 B.n477 585
R619 B.n477 B.n476 585
R620 B.n479 B.n354 585
R621 B.n354 B.n352 585
R622 B.n481 B.n480 585
R623 B.n482 B.n481 585
R624 B.n348 B.n347 585
R625 B.n353 B.n348 585
R626 B.n490 B.n489 585
R627 B.n489 B.n488 585
R628 B.n491 B.n346 585
R629 B.n346 B.n345 585
R630 B.n493 B.n492 585
R631 B.n494 B.n493 585
R632 B.n340 B.n339 585
R633 B.n341 B.n340 585
R634 B.n502 B.n501 585
R635 B.n501 B.n500 585
R636 B.n503 B.n338 585
R637 B.n338 B.n337 585
R638 B.n505 B.n504 585
R639 B.n506 B.n505 585
R640 B.n332 B.n331 585
R641 B.n333 B.n332 585
R642 B.n514 B.n513 585
R643 B.n513 B.n512 585
R644 B.n515 B.n330 585
R645 B.n330 B.n329 585
R646 B.n517 B.n516 585
R647 B.n518 B.n517 585
R648 B.n324 B.n323 585
R649 B.n325 B.n324 585
R650 B.n527 B.n526 585
R651 B.n526 B.n525 585
R652 B.n528 B.n322 585
R653 B.n524 B.n322 585
R654 B.n530 B.n529 585
R655 B.n531 B.n530 585
R656 B.n317 B.n316 585
R657 B.n318 B.n317 585
R658 B.n539 B.n538 585
R659 B.n538 B.n537 585
R660 B.n540 B.n315 585
R661 B.n315 B.n314 585
R662 B.n542 B.n541 585
R663 B.n543 B.n542 585
R664 B.n309 B.n308 585
R665 B.n310 B.n309 585
R666 B.n551 B.n550 585
R667 B.n550 B.n549 585
R668 B.n552 B.n307 585
R669 B.n307 B.n306 585
R670 B.n554 B.n553 585
R671 B.n555 B.n554 585
R672 B.n301 B.n300 585
R673 B.n302 B.n301 585
R674 B.n563 B.n562 585
R675 B.n562 B.n561 585
R676 B.n564 B.n299 585
R677 B.n299 B.n298 585
R678 B.n566 B.n565 585
R679 B.n567 B.n566 585
R680 B.n293 B.n292 585
R681 B.n294 B.n293 585
R682 B.n575 B.n574 585
R683 B.n574 B.n573 585
R684 B.n576 B.n291 585
R685 B.n291 B.n290 585
R686 B.n578 B.n577 585
R687 B.n579 B.n578 585
R688 B.n285 B.n284 585
R689 B.n286 B.n285 585
R690 B.n587 B.n586 585
R691 B.n586 B.n585 585
R692 B.n588 B.n283 585
R693 B.n283 B.n281 585
R694 B.n590 B.n589 585
R695 B.n591 B.n590 585
R696 B.n277 B.n276 585
R697 B.n282 B.n277 585
R698 B.n599 B.n598 585
R699 B.n598 B.n597 585
R700 B.n600 B.n275 585
R701 B.n275 B.n274 585
R702 B.n602 B.n601 585
R703 B.n603 B.n602 585
R704 B.n269 B.n268 585
R705 B.n270 B.n269 585
R706 B.n611 B.n610 585
R707 B.n610 B.n609 585
R708 B.n612 B.n267 585
R709 B.n267 B.n266 585
R710 B.n614 B.n613 585
R711 B.n615 B.n614 585
R712 B.n261 B.n260 585
R713 B.n262 B.n261 585
R714 B.n623 B.n622 585
R715 B.n622 B.n621 585
R716 B.n624 B.n259 585
R717 B.n259 B.n258 585
R718 B.n626 B.n625 585
R719 B.n627 B.n626 585
R720 B.n253 B.n252 585
R721 B.n254 B.n253 585
R722 B.n635 B.n634 585
R723 B.n634 B.n633 585
R724 B.n636 B.n251 585
R725 B.n251 B.n250 585
R726 B.n638 B.n637 585
R727 B.n639 B.n638 585
R728 B.n245 B.n244 585
R729 B.n246 B.n245 585
R730 B.n647 B.n646 585
R731 B.n646 B.n645 585
R732 B.n648 B.n243 585
R733 B.n243 B.n242 585
R734 B.n650 B.n649 585
R735 B.n651 B.n650 585
R736 B.n237 B.n236 585
R737 B.n238 B.n237 585
R738 B.n660 B.n659 585
R739 B.n659 B.n658 585
R740 B.n661 B.n235 585
R741 B.n657 B.n235 585
R742 B.n663 B.n662 585
R743 B.n664 B.n663 585
R744 B.n230 B.n229 585
R745 B.n231 B.n230 585
R746 B.n673 B.n672 585
R747 B.n672 B.n671 585
R748 B.n674 B.n228 585
R749 B.n228 B.n227 585
R750 B.n676 B.n675 585
R751 B.n677 B.n676 585
R752 B.n3 B.n0 585
R753 B.n4 B.n3 585
R754 B.n921 B.n1 585
R755 B.n922 B.n921 585
R756 B.n920 B.n919 585
R757 B.n920 B.n8 585
R758 B.n918 B.n9 585
R759 B.n12 B.n9 585
R760 B.n917 B.n916 585
R761 B.n916 B.n915 585
R762 B.n11 B.n10 585
R763 B.n914 B.n11 585
R764 B.n912 B.n911 585
R765 B.n913 B.n912 585
R766 B.n910 B.n16 585
R767 B.n19 B.n16 585
R768 B.n909 B.n908 585
R769 B.n908 B.n907 585
R770 B.n18 B.n17 585
R771 B.n906 B.n18 585
R772 B.n904 B.n903 585
R773 B.n905 B.n904 585
R774 B.n902 B.n24 585
R775 B.n24 B.n23 585
R776 B.n901 B.n900 585
R777 B.n900 B.n899 585
R778 B.n26 B.n25 585
R779 B.n898 B.n26 585
R780 B.n896 B.n895 585
R781 B.n897 B.n896 585
R782 B.n894 B.n31 585
R783 B.n31 B.n30 585
R784 B.n893 B.n892 585
R785 B.n892 B.n891 585
R786 B.n33 B.n32 585
R787 B.n890 B.n33 585
R788 B.n888 B.n887 585
R789 B.n889 B.n888 585
R790 B.n886 B.n38 585
R791 B.n38 B.n37 585
R792 B.n885 B.n884 585
R793 B.n884 B.n883 585
R794 B.n40 B.n39 585
R795 B.n882 B.n40 585
R796 B.n880 B.n879 585
R797 B.n881 B.n880 585
R798 B.n878 B.n45 585
R799 B.n45 B.n44 585
R800 B.n877 B.n876 585
R801 B.n876 B.n875 585
R802 B.n47 B.n46 585
R803 B.n874 B.n47 585
R804 B.n872 B.n871 585
R805 B.n873 B.n872 585
R806 B.n870 B.n52 585
R807 B.n52 B.n51 585
R808 B.n869 B.n868 585
R809 B.n868 B.n867 585
R810 B.n54 B.n53 585
R811 B.n866 B.n54 585
R812 B.n864 B.n863 585
R813 B.n865 B.n864 585
R814 B.n862 B.n59 585
R815 B.n59 B.n58 585
R816 B.n861 B.n860 585
R817 B.n860 B.n859 585
R818 B.n61 B.n60 585
R819 B.n858 B.n61 585
R820 B.n856 B.n855 585
R821 B.n857 B.n856 585
R822 B.n854 B.n66 585
R823 B.n66 B.n65 585
R824 B.n853 B.n852 585
R825 B.n852 B.n851 585
R826 B.n68 B.n67 585
R827 B.n850 B.n68 585
R828 B.n848 B.n847 585
R829 B.n849 B.n848 585
R830 B.n846 B.n73 585
R831 B.n73 B.n72 585
R832 B.n845 B.n844 585
R833 B.n844 B.n843 585
R834 B.n75 B.n74 585
R835 B.n842 B.n75 585
R836 B.n840 B.n839 585
R837 B.n841 B.n840 585
R838 B.n838 B.n80 585
R839 B.n80 B.n79 585
R840 B.n837 B.n836 585
R841 B.n836 B.n835 585
R842 B.n82 B.n81 585
R843 B.n834 B.n82 585
R844 B.n832 B.n831 585
R845 B.n833 B.n832 585
R846 B.n830 B.n87 585
R847 B.n87 B.n86 585
R848 B.n829 B.n828 585
R849 B.n828 B.n827 585
R850 B.n89 B.n88 585
R851 B.n826 B.n89 585
R852 B.n824 B.n823 585
R853 B.n825 B.n824 585
R854 B.n822 B.n93 585
R855 B.n96 B.n93 585
R856 B.n821 B.n820 585
R857 B.n820 B.n819 585
R858 B.n95 B.n94 585
R859 B.n818 B.n95 585
R860 B.n816 B.n815 585
R861 B.n817 B.n816 585
R862 B.n814 B.n101 585
R863 B.n101 B.n100 585
R864 B.n813 B.n812 585
R865 B.n812 B.n811 585
R866 B.n103 B.n102 585
R867 B.n810 B.n103 585
R868 B.n808 B.n807 585
R869 B.n809 B.n808 585
R870 B.n806 B.n108 585
R871 B.n108 B.n107 585
R872 B.n805 B.n804 585
R873 B.n804 B.n803 585
R874 B.n110 B.n109 585
R875 B.n802 B.n110 585
R876 B.n800 B.n799 585
R877 B.n801 B.n800 585
R878 B.n798 B.n115 585
R879 B.n115 B.n114 585
R880 B.n797 B.n796 585
R881 B.n796 B.n795 585
R882 B.n117 B.n116 585
R883 B.n794 B.n117 585
R884 B.n792 B.n791 585
R885 B.n793 B.n792 585
R886 B.n790 B.n122 585
R887 B.n122 B.n121 585
R888 B.n789 B.n788 585
R889 B.n788 B.n787 585
R890 B.n124 B.n123 585
R891 B.n786 B.n124 585
R892 B.n784 B.n783 585
R893 B.n785 B.n784 585
R894 B.n782 B.n129 585
R895 B.n129 B.n128 585
R896 B.n781 B.n780 585
R897 B.n780 B.n779 585
R898 B.n131 B.n130 585
R899 B.n778 B.n131 585
R900 B.n925 B.n924 585
R901 B.n923 B.n2 585
R902 B.n157 B.n131 545.355
R903 B.n776 B.n133 545.355
R904 B.n459 B.n366 545.355
R905 B.n455 B.n364 545.355
R906 B.n777 B.n150 256.663
R907 B.n777 B.n149 256.663
R908 B.n777 B.n148 256.663
R909 B.n777 B.n147 256.663
R910 B.n777 B.n146 256.663
R911 B.n777 B.n145 256.663
R912 B.n777 B.n144 256.663
R913 B.n777 B.n143 256.663
R914 B.n777 B.n142 256.663
R915 B.n777 B.n141 256.663
R916 B.n777 B.n140 256.663
R917 B.n777 B.n139 256.663
R918 B.n777 B.n138 256.663
R919 B.n777 B.n137 256.663
R920 B.n777 B.n136 256.663
R921 B.n777 B.n135 256.663
R922 B.n777 B.n134 256.663
R923 B.n457 B.n456 256.663
R924 B.n457 B.n369 256.663
R925 B.n457 B.n370 256.663
R926 B.n457 B.n371 256.663
R927 B.n457 B.n372 256.663
R928 B.n457 B.n373 256.663
R929 B.n457 B.n374 256.663
R930 B.n457 B.n375 256.663
R931 B.n457 B.n376 256.663
R932 B.n457 B.n377 256.663
R933 B.n457 B.n378 256.663
R934 B.n457 B.n379 256.663
R935 B.n457 B.n380 256.663
R936 B.n457 B.n381 256.663
R937 B.n457 B.n382 256.663
R938 B.n457 B.n383 256.663
R939 B.n458 B.n457 256.663
R940 B.n927 B.n926 256.663
R941 B.n155 B.t17 224.49
R942 B.n152 B.t21 224.49
R943 B.n389 B.t10 224.49
R944 B.n386 B.t14 224.49
R945 B.n457 B.n365 208.048
R946 B.n778 B.n777 208.048
R947 B.n161 B.n160 163.367
R948 B.n165 B.n164 163.367
R949 B.n169 B.n168 163.367
R950 B.n173 B.n172 163.367
R951 B.n177 B.n176 163.367
R952 B.n181 B.n180 163.367
R953 B.n186 B.n185 163.367
R954 B.n190 B.n189 163.367
R955 B.n194 B.n193 163.367
R956 B.n198 B.n197 163.367
R957 B.n202 B.n201 163.367
R958 B.n206 B.n205 163.367
R959 B.n210 B.n209 163.367
R960 B.n214 B.n213 163.367
R961 B.n218 B.n217 163.367
R962 B.n222 B.n221 163.367
R963 B.n776 B.n151 163.367
R964 B.n463 B.n366 163.367
R965 B.n463 B.n360 163.367
R966 B.n471 B.n360 163.367
R967 B.n471 B.n358 163.367
R968 B.n475 B.n358 163.367
R969 B.n475 B.n351 163.367
R970 B.n483 B.n351 163.367
R971 B.n483 B.n349 163.367
R972 B.n487 B.n349 163.367
R973 B.n487 B.n344 163.367
R974 B.n495 B.n344 163.367
R975 B.n495 B.n342 163.367
R976 B.n499 B.n342 163.367
R977 B.n499 B.n336 163.367
R978 B.n507 B.n336 163.367
R979 B.n507 B.n334 163.367
R980 B.n511 B.n334 163.367
R981 B.n511 B.n328 163.367
R982 B.n519 B.n328 163.367
R983 B.n519 B.n326 163.367
R984 B.n523 B.n326 163.367
R985 B.n523 B.n321 163.367
R986 B.n532 B.n321 163.367
R987 B.n532 B.n319 163.367
R988 B.n536 B.n319 163.367
R989 B.n536 B.n313 163.367
R990 B.n544 B.n313 163.367
R991 B.n544 B.n311 163.367
R992 B.n548 B.n311 163.367
R993 B.n548 B.n305 163.367
R994 B.n556 B.n305 163.367
R995 B.n556 B.n303 163.367
R996 B.n560 B.n303 163.367
R997 B.n560 B.n297 163.367
R998 B.n568 B.n297 163.367
R999 B.n568 B.n295 163.367
R1000 B.n572 B.n295 163.367
R1001 B.n572 B.n289 163.367
R1002 B.n580 B.n289 163.367
R1003 B.n580 B.n287 163.367
R1004 B.n584 B.n287 163.367
R1005 B.n584 B.n280 163.367
R1006 B.n592 B.n280 163.367
R1007 B.n592 B.n278 163.367
R1008 B.n596 B.n278 163.367
R1009 B.n596 B.n273 163.367
R1010 B.n604 B.n273 163.367
R1011 B.n604 B.n271 163.367
R1012 B.n608 B.n271 163.367
R1013 B.n608 B.n265 163.367
R1014 B.n616 B.n265 163.367
R1015 B.n616 B.n263 163.367
R1016 B.n620 B.n263 163.367
R1017 B.n620 B.n257 163.367
R1018 B.n628 B.n257 163.367
R1019 B.n628 B.n255 163.367
R1020 B.n632 B.n255 163.367
R1021 B.n632 B.n249 163.367
R1022 B.n640 B.n249 163.367
R1023 B.n640 B.n247 163.367
R1024 B.n644 B.n247 163.367
R1025 B.n644 B.n241 163.367
R1026 B.n652 B.n241 163.367
R1027 B.n652 B.n239 163.367
R1028 B.n656 B.n239 163.367
R1029 B.n656 B.n234 163.367
R1030 B.n665 B.n234 163.367
R1031 B.n665 B.n232 163.367
R1032 B.n670 B.n232 163.367
R1033 B.n670 B.n226 163.367
R1034 B.n678 B.n226 163.367
R1035 B.n679 B.n678 163.367
R1036 B.n679 B.n5 163.367
R1037 B.n6 B.n5 163.367
R1038 B.n7 B.n6 163.367
R1039 B.n685 B.n7 163.367
R1040 B.n686 B.n685 163.367
R1041 B.n686 B.n13 163.367
R1042 B.n14 B.n13 163.367
R1043 B.n15 B.n14 163.367
R1044 B.n691 B.n15 163.367
R1045 B.n691 B.n20 163.367
R1046 B.n21 B.n20 163.367
R1047 B.n22 B.n21 163.367
R1048 B.n696 B.n22 163.367
R1049 B.n696 B.n27 163.367
R1050 B.n28 B.n27 163.367
R1051 B.n29 B.n28 163.367
R1052 B.n701 B.n29 163.367
R1053 B.n701 B.n34 163.367
R1054 B.n35 B.n34 163.367
R1055 B.n36 B.n35 163.367
R1056 B.n706 B.n36 163.367
R1057 B.n706 B.n41 163.367
R1058 B.n42 B.n41 163.367
R1059 B.n43 B.n42 163.367
R1060 B.n711 B.n43 163.367
R1061 B.n711 B.n48 163.367
R1062 B.n49 B.n48 163.367
R1063 B.n50 B.n49 163.367
R1064 B.n716 B.n50 163.367
R1065 B.n716 B.n55 163.367
R1066 B.n56 B.n55 163.367
R1067 B.n57 B.n56 163.367
R1068 B.n721 B.n57 163.367
R1069 B.n721 B.n62 163.367
R1070 B.n63 B.n62 163.367
R1071 B.n64 B.n63 163.367
R1072 B.n726 B.n64 163.367
R1073 B.n726 B.n69 163.367
R1074 B.n70 B.n69 163.367
R1075 B.n71 B.n70 163.367
R1076 B.n731 B.n71 163.367
R1077 B.n731 B.n76 163.367
R1078 B.n77 B.n76 163.367
R1079 B.n78 B.n77 163.367
R1080 B.n736 B.n78 163.367
R1081 B.n736 B.n83 163.367
R1082 B.n84 B.n83 163.367
R1083 B.n85 B.n84 163.367
R1084 B.n741 B.n85 163.367
R1085 B.n741 B.n90 163.367
R1086 B.n91 B.n90 163.367
R1087 B.n92 B.n91 163.367
R1088 B.n746 B.n92 163.367
R1089 B.n746 B.n97 163.367
R1090 B.n98 B.n97 163.367
R1091 B.n99 B.n98 163.367
R1092 B.n751 B.n99 163.367
R1093 B.n751 B.n104 163.367
R1094 B.n105 B.n104 163.367
R1095 B.n106 B.n105 163.367
R1096 B.n756 B.n106 163.367
R1097 B.n756 B.n111 163.367
R1098 B.n112 B.n111 163.367
R1099 B.n113 B.n112 163.367
R1100 B.n761 B.n113 163.367
R1101 B.n761 B.n118 163.367
R1102 B.n119 B.n118 163.367
R1103 B.n120 B.n119 163.367
R1104 B.n766 B.n120 163.367
R1105 B.n766 B.n125 163.367
R1106 B.n126 B.n125 163.367
R1107 B.n127 B.n126 163.367
R1108 B.n771 B.n127 163.367
R1109 B.n771 B.n132 163.367
R1110 B.n133 B.n132 163.367
R1111 B.n385 B.n384 163.367
R1112 B.n450 B.n384 163.367
R1113 B.n448 B.n447 163.367
R1114 B.n444 B.n443 163.367
R1115 B.n440 B.n439 163.367
R1116 B.n436 B.n435 163.367
R1117 B.n432 B.n431 163.367
R1118 B.n428 B.n427 163.367
R1119 B.n424 B.n423 163.367
R1120 B.n420 B.n419 163.367
R1121 B.n416 B.n415 163.367
R1122 B.n411 B.n410 163.367
R1123 B.n407 B.n406 163.367
R1124 B.n403 B.n402 163.367
R1125 B.n399 B.n398 163.367
R1126 B.n395 B.n394 163.367
R1127 B.n391 B.n368 163.367
R1128 B.n465 B.n364 163.367
R1129 B.n465 B.n362 163.367
R1130 B.n469 B.n362 163.367
R1131 B.n469 B.n356 163.367
R1132 B.n477 B.n356 163.367
R1133 B.n477 B.n354 163.367
R1134 B.n481 B.n354 163.367
R1135 B.n481 B.n348 163.367
R1136 B.n489 B.n348 163.367
R1137 B.n489 B.n346 163.367
R1138 B.n493 B.n346 163.367
R1139 B.n493 B.n340 163.367
R1140 B.n501 B.n340 163.367
R1141 B.n501 B.n338 163.367
R1142 B.n505 B.n338 163.367
R1143 B.n505 B.n332 163.367
R1144 B.n513 B.n332 163.367
R1145 B.n513 B.n330 163.367
R1146 B.n517 B.n330 163.367
R1147 B.n517 B.n324 163.367
R1148 B.n526 B.n324 163.367
R1149 B.n526 B.n322 163.367
R1150 B.n530 B.n322 163.367
R1151 B.n530 B.n317 163.367
R1152 B.n538 B.n317 163.367
R1153 B.n538 B.n315 163.367
R1154 B.n542 B.n315 163.367
R1155 B.n542 B.n309 163.367
R1156 B.n550 B.n309 163.367
R1157 B.n550 B.n307 163.367
R1158 B.n554 B.n307 163.367
R1159 B.n554 B.n301 163.367
R1160 B.n562 B.n301 163.367
R1161 B.n562 B.n299 163.367
R1162 B.n566 B.n299 163.367
R1163 B.n566 B.n293 163.367
R1164 B.n574 B.n293 163.367
R1165 B.n574 B.n291 163.367
R1166 B.n578 B.n291 163.367
R1167 B.n578 B.n285 163.367
R1168 B.n586 B.n285 163.367
R1169 B.n586 B.n283 163.367
R1170 B.n590 B.n283 163.367
R1171 B.n590 B.n277 163.367
R1172 B.n598 B.n277 163.367
R1173 B.n598 B.n275 163.367
R1174 B.n602 B.n275 163.367
R1175 B.n602 B.n269 163.367
R1176 B.n610 B.n269 163.367
R1177 B.n610 B.n267 163.367
R1178 B.n614 B.n267 163.367
R1179 B.n614 B.n261 163.367
R1180 B.n622 B.n261 163.367
R1181 B.n622 B.n259 163.367
R1182 B.n626 B.n259 163.367
R1183 B.n626 B.n253 163.367
R1184 B.n634 B.n253 163.367
R1185 B.n634 B.n251 163.367
R1186 B.n638 B.n251 163.367
R1187 B.n638 B.n245 163.367
R1188 B.n646 B.n245 163.367
R1189 B.n646 B.n243 163.367
R1190 B.n650 B.n243 163.367
R1191 B.n650 B.n237 163.367
R1192 B.n659 B.n237 163.367
R1193 B.n659 B.n235 163.367
R1194 B.n663 B.n235 163.367
R1195 B.n663 B.n230 163.367
R1196 B.n672 B.n230 163.367
R1197 B.n672 B.n228 163.367
R1198 B.n676 B.n228 163.367
R1199 B.n676 B.n3 163.367
R1200 B.n925 B.n3 163.367
R1201 B.n921 B.n2 163.367
R1202 B.n921 B.n920 163.367
R1203 B.n920 B.n9 163.367
R1204 B.n916 B.n9 163.367
R1205 B.n916 B.n11 163.367
R1206 B.n912 B.n11 163.367
R1207 B.n912 B.n16 163.367
R1208 B.n908 B.n16 163.367
R1209 B.n908 B.n18 163.367
R1210 B.n904 B.n18 163.367
R1211 B.n904 B.n24 163.367
R1212 B.n900 B.n24 163.367
R1213 B.n900 B.n26 163.367
R1214 B.n896 B.n26 163.367
R1215 B.n896 B.n31 163.367
R1216 B.n892 B.n31 163.367
R1217 B.n892 B.n33 163.367
R1218 B.n888 B.n33 163.367
R1219 B.n888 B.n38 163.367
R1220 B.n884 B.n38 163.367
R1221 B.n884 B.n40 163.367
R1222 B.n880 B.n40 163.367
R1223 B.n880 B.n45 163.367
R1224 B.n876 B.n45 163.367
R1225 B.n876 B.n47 163.367
R1226 B.n872 B.n47 163.367
R1227 B.n872 B.n52 163.367
R1228 B.n868 B.n52 163.367
R1229 B.n868 B.n54 163.367
R1230 B.n864 B.n54 163.367
R1231 B.n864 B.n59 163.367
R1232 B.n860 B.n59 163.367
R1233 B.n860 B.n61 163.367
R1234 B.n856 B.n61 163.367
R1235 B.n856 B.n66 163.367
R1236 B.n852 B.n66 163.367
R1237 B.n852 B.n68 163.367
R1238 B.n848 B.n68 163.367
R1239 B.n848 B.n73 163.367
R1240 B.n844 B.n73 163.367
R1241 B.n844 B.n75 163.367
R1242 B.n840 B.n75 163.367
R1243 B.n840 B.n80 163.367
R1244 B.n836 B.n80 163.367
R1245 B.n836 B.n82 163.367
R1246 B.n832 B.n82 163.367
R1247 B.n832 B.n87 163.367
R1248 B.n828 B.n87 163.367
R1249 B.n828 B.n89 163.367
R1250 B.n824 B.n89 163.367
R1251 B.n824 B.n93 163.367
R1252 B.n820 B.n93 163.367
R1253 B.n820 B.n95 163.367
R1254 B.n816 B.n95 163.367
R1255 B.n816 B.n101 163.367
R1256 B.n812 B.n101 163.367
R1257 B.n812 B.n103 163.367
R1258 B.n808 B.n103 163.367
R1259 B.n808 B.n108 163.367
R1260 B.n804 B.n108 163.367
R1261 B.n804 B.n110 163.367
R1262 B.n800 B.n110 163.367
R1263 B.n800 B.n115 163.367
R1264 B.n796 B.n115 163.367
R1265 B.n796 B.n117 163.367
R1266 B.n792 B.n117 163.367
R1267 B.n792 B.n122 163.367
R1268 B.n788 B.n122 163.367
R1269 B.n788 B.n124 163.367
R1270 B.n784 B.n124 163.367
R1271 B.n784 B.n129 163.367
R1272 B.n780 B.n129 163.367
R1273 B.n780 B.n131 163.367
R1274 B.n152 B.t22 157.548
R1275 B.n389 B.t13 157.548
R1276 B.n155 B.t19 157.548
R1277 B.n386 B.t16 157.548
R1278 B.n464 B.n365 100.335
R1279 B.n464 B.n361 100.335
R1280 B.n470 B.n361 100.335
R1281 B.n470 B.n357 100.335
R1282 B.n476 B.n357 100.335
R1283 B.n476 B.n352 100.335
R1284 B.n482 B.n352 100.335
R1285 B.n482 B.n353 100.335
R1286 B.n488 B.n345 100.335
R1287 B.n494 B.n345 100.335
R1288 B.n494 B.n341 100.335
R1289 B.n500 B.n341 100.335
R1290 B.n500 B.n337 100.335
R1291 B.n506 B.n337 100.335
R1292 B.n506 B.n333 100.335
R1293 B.n512 B.n333 100.335
R1294 B.n512 B.n329 100.335
R1295 B.n518 B.n329 100.335
R1296 B.n518 B.n325 100.335
R1297 B.n525 B.n325 100.335
R1298 B.n525 B.n524 100.335
R1299 B.n531 B.n318 100.335
R1300 B.n537 B.n318 100.335
R1301 B.n537 B.n314 100.335
R1302 B.n543 B.n314 100.335
R1303 B.n543 B.n310 100.335
R1304 B.n549 B.n310 100.335
R1305 B.n549 B.n306 100.335
R1306 B.n555 B.n306 100.335
R1307 B.n555 B.n302 100.335
R1308 B.n561 B.n302 100.335
R1309 B.n567 B.n298 100.335
R1310 B.n567 B.n294 100.335
R1311 B.n573 B.n294 100.335
R1312 B.n573 B.n290 100.335
R1313 B.n579 B.n290 100.335
R1314 B.n579 B.n286 100.335
R1315 B.n585 B.n286 100.335
R1316 B.n585 B.n281 100.335
R1317 B.n591 B.n281 100.335
R1318 B.n591 B.n282 100.335
R1319 B.n597 B.n274 100.335
R1320 B.n603 B.n274 100.335
R1321 B.n603 B.n270 100.335
R1322 B.n609 B.n270 100.335
R1323 B.n609 B.n266 100.335
R1324 B.n615 B.n266 100.335
R1325 B.n615 B.n262 100.335
R1326 B.n621 B.n262 100.335
R1327 B.n621 B.n258 100.335
R1328 B.n627 B.n258 100.335
R1329 B.n633 B.n254 100.335
R1330 B.n633 B.n250 100.335
R1331 B.n639 B.n250 100.335
R1332 B.n639 B.n246 100.335
R1333 B.n645 B.n246 100.335
R1334 B.n645 B.n242 100.335
R1335 B.n651 B.n242 100.335
R1336 B.n651 B.n238 100.335
R1337 B.n658 B.n238 100.335
R1338 B.n658 B.n657 100.335
R1339 B.n664 B.n231 100.335
R1340 B.n671 B.n231 100.335
R1341 B.n671 B.n227 100.335
R1342 B.n677 B.n227 100.335
R1343 B.n677 B.n4 100.335
R1344 B.n924 B.n4 100.335
R1345 B.n924 B.n923 100.335
R1346 B.n923 B.n922 100.335
R1347 B.n922 B.n8 100.335
R1348 B.n12 B.n8 100.335
R1349 B.n915 B.n12 100.335
R1350 B.n915 B.n914 100.335
R1351 B.n914 B.n913 100.335
R1352 B.n907 B.n19 100.335
R1353 B.n907 B.n906 100.335
R1354 B.n906 B.n905 100.335
R1355 B.n905 B.n23 100.335
R1356 B.n899 B.n23 100.335
R1357 B.n899 B.n898 100.335
R1358 B.n898 B.n897 100.335
R1359 B.n897 B.n30 100.335
R1360 B.n891 B.n30 100.335
R1361 B.n891 B.n890 100.335
R1362 B.n889 B.n37 100.335
R1363 B.n883 B.n37 100.335
R1364 B.n883 B.n882 100.335
R1365 B.n882 B.n881 100.335
R1366 B.n881 B.n44 100.335
R1367 B.n875 B.n44 100.335
R1368 B.n875 B.n874 100.335
R1369 B.n874 B.n873 100.335
R1370 B.n873 B.n51 100.335
R1371 B.n867 B.n51 100.335
R1372 B.n866 B.n865 100.335
R1373 B.n865 B.n58 100.335
R1374 B.n859 B.n58 100.335
R1375 B.n859 B.n858 100.335
R1376 B.n858 B.n857 100.335
R1377 B.n857 B.n65 100.335
R1378 B.n851 B.n65 100.335
R1379 B.n851 B.n850 100.335
R1380 B.n850 B.n849 100.335
R1381 B.n849 B.n72 100.335
R1382 B.n843 B.n842 100.335
R1383 B.n842 B.n841 100.335
R1384 B.n841 B.n79 100.335
R1385 B.n835 B.n79 100.335
R1386 B.n835 B.n834 100.335
R1387 B.n834 B.n833 100.335
R1388 B.n833 B.n86 100.335
R1389 B.n827 B.n86 100.335
R1390 B.n827 B.n826 100.335
R1391 B.n826 B.n825 100.335
R1392 B.n819 B.n96 100.335
R1393 B.n819 B.n818 100.335
R1394 B.n818 B.n817 100.335
R1395 B.n817 B.n100 100.335
R1396 B.n811 B.n100 100.335
R1397 B.n811 B.n810 100.335
R1398 B.n810 B.n809 100.335
R1399 B.n809 B.n107 100.335
R1400 B.n803 B.n107 100.335
R1401 B.n803 B.n802 100.335
R1402 B.n802 B.n801 100.335
R1403 B.n801 B.n114 100.335
R1404 B.n795 B.n114 100.335
R1405 B.n794 B.n793 100.335
R1406 B.n793 B.n121 100.335
R1407 B.n787 B.n121 100.335
R1408 B.n787 B.n786 100.335
R1409 B.n786 B.n785 100.335
R1410 B.n785 B.n128 100.335
R1411 B.n779 B.n128 100.335
R1412 B.n779 B.n778 100.335
R1413 B.n153 B.t23 85.4025
R1414 B.n390 B.t12 85.4025
R1415 B.n156 B.t20 85.4022
R1416 B.n387 B.t15 85.4022
R1417 B.n156 B.n155 72.146
R1418 B.n153 B.n152 72.146
R1419 B.n390 B.n389 72.146
R1420 B.n387 B.n386 72.146
R1421 B.n157 B.n134 71.676
R1422 B.n161 B.n135 71.676
R1423 B.n165 B.n136 71.676
R1424 B.n169 B.n137 71.676
R1425 B.n173 B.n138 71.676
R1426 B.n177 B.n139 71.676
R1427 B.n181 B.n140 71.676
R1428 B.n186 B.n141 71.676
R1429 B.n190 B.n142 71.676
R1430 B.n194 B.n143 71.676
R1431 B.n198 B.n144 71.676
R1432 B.n202 B.n145 71.676
R1433 B.n206 B.n146 71.676
R1434 B.n210 B.n147 71.676
R1435 B.n214 B.n148 71.676
R1436 B.n218 B.n149 71.676
R1437 B.n222 B.n150 71.676
R1438 B.n151 B.n150 71.676
R1439 B.n221 B.n149 71.676
R1440 B.n217 B.n148 71.676
R1441 B.n213 B.n147 71.676
R1442 B.n209 B.n146 71.676
R1443 B.n205 B.n145 71.676
R1444 B.n201 B.n144 71.676
R1445 B.n197 B.n143 71.676
R1446 B.n193 B.n142 71.676
R1447 B.n189 B.n141 71.676
R1448 B.n185 B.n140 71.676
R1449 B.n180 B.n139 71.676
R1450 B.n176 B.n138 71.676
R1451 B.n172 B.n137 71.676
R1452 B.n168 B.n136 71.676
R1453 B.n164 B.n135 71.676
R1454 B.n160 B.n134 71.676
R1455 B.n456 B.n455 71.676
R1456 B.n450 B.n369 71.676
R1457 B.n447 B.n370 71.676
R1458 B.n443 B.n371 71.676
R1459 B.n439 B.n372 71.676
R1460 B.n435 B.n373 71.676
R1461 B.n431 B.n374 71.676
R1462 B.n427 B.n375 71.676
R1463 B.n423 B.n376 71.676
R1464 B.n419 B.n377 71.676
R1465 B.n415 B.n378 71.676
R1466 B.n410 B.n379 71.676
R1467 B.n406 B.n380 71.676
R1468 B.n402 B.n381 71.676
R1469 B.n398 B.n382 71.676
R1470 B.n394 B.n383 71.676
R1471 B.n458 B.n368 71.676
R1472 B.n456 B.n385 71.676
R1473 B.n448 B.n369 71.676
R1474 B.n444 B.n370 71.676
R1475 B.n440 B.n371 71.676
R1476 B.n436 B.n372 71.676
R1477 B.n432 B.n373 71.676
R1478 B.n428 B.n374 71.676
R1479 B.n424 B.n375 71.676
R1480 B.n420 B.n376 71.676
R1481 B.n416 B.n377 71.676
R1482 B.n411 B.n378 71.676
R1483 B.n407 B.n379 71.676
R1484 B.n403 B.n380 71.676
R1485 B.n399 B.n381 71.676
R1486 B.n395 B.n382 71.676
R1487 B.n391 B.n383 71.676
R1488 B.n459 B.n458 71.676
R1489 B.n926 B.n925 71.676
R1490 B.n926 B.n2 71.676
R1491 B.n524 B.t1 66.3989
R1492 B.n96 B.t7 66.3989
R1493 B.n561 B.t8 60.4968
R1494 B.n843 B.t9 60.4968
R1495 B.n183 B.n156 59.5399
R1496 B.n154 B.n153 59.5399
R1497 B.n413 B.n390 59.5399
R1498 B.n388 B.n387 59.5399
R1499 B.n664 B.t0 57.5458
R1500 B.n913 B.t5 57.5458
R1501 B.n282 B.t3 54.5947
R1502 B.t6 B.n866 54.5947
R1503 B.n353 B.t11 51.6437
R1504 B.t4 B.n254 51.6437
R1505 B.n890 B.t2 51.6437
R1506 B.t18 B.n794 51.6437
R1507 B.n488 B.t11 48.6927
R1508 B.n627 B.t4 48.6927
R1509 B.t2 B.n889 48.6927
R1510 B.n795 B.t18 48.6927
R1511 B.n597 B.t3 45.7416
R1512 B.n867 B.t6 45.7416
R1513 B.n657 B.t0 42.7906
R1514 B.n19 B.t5 42.7906
R1515 B.t8 B.n298 39.8395
R1516 B.t9 B.n72 39.8395
R1517 B.n454 B.n363 35.4346
R1518 B.n461 B.n460 35.4346
R1519 B.n775 B.n774 35.4346
R1520 B.n158 B.n130 35.4346
R1521 B.n531 B.t1 33.9375
R1522 B.n825 B.t7 33.9375
R1523 B B.n927 18.0485
R1524 B.n466 B.n363 10.6151
R1525 B.n467 B.n466 10.6151
R1526 B.n468 B.n467 10.6151
R1527 B.n468 B.n355 10.6151
R1528 B.n478 B.n355 10.6151
R1529 B.n479 B.n478 10.6151
R1530 B.n480 B.n479 10.6151
R1531 B.n480 B.n347 10.6151
R1532 B.n490 B.n347 10.6151
R1533 B.n491 B.n490 10.6151
R1534 B.n492 B.n491 10.6151
R1535 B.n492 B.n339 10.6151
R1536 B.n502 B.n339 10.6151
R1537 B.n503 B.n502 10.6151
R1538 B.n504 B.n503 10.6151
R1539 B.n504 B.n331 10.6151
R1540 B.n514 B.n331 10.6151
R1541 B.n515 B.n514 10.6151
R1542 B.n516 B.n515 10.6151
R1543 B.n516 B.n323 10.6151
R1544 B.n527 B.n323 10.6151
R1545 B.n528 B.n527 10.6151
R1546 B.n529 B.n528 10.6151
R1547 B.n529 B.n316 10.6151
R1548 B.n539 B.n316 10.6151
R1549 B.n540 B.n539 10.6151
R1550 B.n541 B.n540 10.6151
R1551 B.n541 B.n308 10.6151
R1552 B.n551 B.n308 10.6151
R1553 B.n552 B.n551 10.6151
R1554 B.n553 B.n552 10.6151
R1555 B.n553 B.n300 10.6151
R1556 B.n563 B.n300 10.6151
R1557 B.n564 B.n563 10.6151
R1558 B.n565 B.n564 10.6151
R1559 B.n565 B.n292 10.6151
R1560 B.n575 B.n292 10.6151
R1561 B.n576 B.n575 10.6151
R1562 B.n577 B.n576 10.6151
R1563 B.n577 B.n284 10.6151
R1564 B.n587 B.n284 10.6151
R1565 B.n588 B.n587 10.6151
R1566 B.n589 B.n588 10.6151
R1567 B.n589 B.n276 10.6151
R1568 B.n599 B.n276 10.6151
R1569 B.n600 B.n599 10.6151
R1570 B.n601 B.n600 10.6151
R1571 B.n601 B.n268 10.6151
R1572 B.n611 B.n268 10.6151
R1573 B.n612 B.n611 10.6151
R1574 B.n613 B.n612 10.6151
R1575 B.n613 B.n260 10.6151
R1576 B.n623 B.n260 10.6151
R1577 B.n624 B.n623 10.6151
R1578 B.n625 B.n624 10.6151
R1579 B.n625 B.n252 10.6151
R1580 B.n635 B.n252 10.6151
R1581 B.n636 B.n635 10.6151
R1582 B.n637 B.n636 10.6151
R1583 B.n637 B.n244 10.6151
R1584 B.n647 B.n244 10.6151
R1585 B.n648 B.n647 10.6151
R1586 B.n649 B.n648 10.6151
R1587 B.n649 B.n236 10.6151
R1588 B.n660 B.n236 10.6151
R1589 B.n661 B.n660 10.6151
R1590 B.n662 B.n661 10.6151
R1591 B.n662 B.n229 10.6151
R1592 B.n673 B.n229 10.6151
R1593 B.n674 B.n673 10.6151
R1594 B.n675 B.n674 10.6151
R1595 B.n675 B.n0 10.6151
R1596 B.n454 B.n453 10.6151
R1597 B.n453 B.n452 10.6151
R1598 B.n452 B.n451 10.6151
R1599 B.n451 B.n449 10.6151
R1600 B.n449 B.n446 10.6151
R1601 B.n446 B.n445 10.6151
R1602 B.n445 B.n442 10.6151
R1603 B.n442 B.n441 10.6151
R1604 B.n441 B.n438 10.6151
R1605 B.n438 B.n437 10.6151
R1606 B.n437 B.n434 10.6151
R1607 B.n434 B.n433 10.6151
R1608 B.n430 B.n429 10.6151
R1609 B.n429 B.n426 10.6151
R1610 B.n426 B.n425 10.6151
R1611 B.n425 B.n422 10.6151
R1612 B.n422 B.n421 10.6151
R1613 B.n421 B.n418 10.6151
R1614 B.n418 B.n417 10.6151
R1615 B.n417 B.n414 10.6151
R1616 B.n412 B.n409 10.6151
R1617 B.n409 B.n408 10.6151
R1618 B.n408 B.n405 10.6151
R1619 B.n405 B.n404 10.6151
R1620 B.n404 B.n401 10.6151
R1621 B.n401 B.n400 10.6151
R1622 B.n400 B.n397 10.6151
R1623 B.n397 B.n396 10.6151
R1624 B.n396 B.n393 10.6151
R1625 B.n393 B.n392 10.6151
R1626 B.n392 B.n367 10.6151
R1627 B.n460 B.n367 10.6151
R1628 B.n462 B.n461 10.6151
R1629 B.n462 B.n359 10.6151
R1630 B.n472 B.n359 10.6151
R1631 B.n473 B.n472 10.6151
R1632 B.n474 B.n473 10.6151
R1633 B.n474 B.n350 10.6151
R1634 B.n484 B.n350 10.6151
R1635 B.n485 B.n484 10.6151
R1636 B.n486 B.n485 10.6151
R1637 B.n486 B.n343 10.6151
R1638 B.n496 B.n343 10.6151
R1639 B.n497 B.n496 10.6151
R1640 B.n498 B.n497 10.6151
R1641 B.n498 B.n335 10.6151
R1642 B.n508 B.n335 10.6151
R1643 B.n509 B.n508 10.6151
R1644 B.n510 B.n509 10.6151
R1645 B.n510 B.n327 10.6151
R1646 B.n520 B.n327 10.6151
R1647 B.n521 B.n520 10.6151
R1648 B.n522 B.n521 10.6151
R1649 B.n522 B.n320 10.6151
R1650 B.n533 B.n320 10.6151
R1651 B.n534 B.n533 10.6151
R1652 B.n535 B.n534 10.6151
R1653 B.n535 B.n312 10.6151
R1654 B.n545 B.n312 10.6151
R1655 B.n546 B.n545 10.6151
R1656 B.n547 B.n546 10.6151
R1657 B.n547 B.n304 10.6151
R1658 B.n557 B.n304 10.6151
R1659 B.n558 B.n557 10.6151
R1660 B.n559 B.n558 10.6151
R1661 B.n559 B.n296 10.6151
R1662 B.n569 B.n296 10.6151
R1663 B.n570 B.n569 10.6151
R1664 B.n571 B.n570 10.6151
R1665 B.n571 B.n288 10.6151
R1666 B.n581 B.n288 10.6151
R1667 B.n582 B.n581 10.6151
R1668 B.n583 B.n582 10.6151
R1669 B.n583 B.n279 10.6151
R1670 B.n593 B.n279 10.6151
R1671 B.n594 B.n593 10.6151
R1672 B.n595 B.n594 10.6151
R1673 B.n595 B.n272 10.6151
R1674 B.n605 B.n272 10.6151
R1675 B.n606 B.n605 10.6151
R1676 B.n607 B.n606 10.6151
R1677 B.n607 B.n264 10.6151
R1678 B.n617 B.n264 10.6151
R1679 B.n618 B.n617 10.6151
R1680 B.n619 B.n618 10.6151
R1681 B.n619 B.n256 10.6151
R1682 B.n629 B.n256 10.6151
R1683 B.n630 B.n629 10.6151
R1684 B.n631 B.n630 10.6151
R1685 B.n631 B.n248 10.6151
R1686 B.n641 B.n248 10.6151
R1687 B.n642 B.n641 10.6151
R1688 B.n643 B.n642 10.6151
R1689 B.n643 B.n240 10.6151
R1690 B.n653 B.n240 10.6151
R1691 B.n654 B.n653 10.6151
R1692 B.n655 B.n654 10.6151
R1693 B.n655 B.n233 10.6151
R1694 B.n666 B.n233 10.6151
R1695 B.n667 B.n666 10.6151
R1696 B.n669 B.n667 10.6151
R1697 B.n669 B.n668 10.6151
R1698 B.n668 B.n225 10.6151
R1699 B.n680 B.n225 10.6151
R1700 B.n681 B.n680 10.6151
R1701 B.n682 B.n681 10.6151
R1702 B.n683 B.n682 10.6151
R1703 B.n684 B.n683 10.6151
R1704 B.n687 B.n684 10.6151
R1705 B.n688 B.n687 10.6151
R1706 B.n689 B.n688 10.6151
R1707 B.n690 B.n689 10.6151
R1708 B.n692 B.n690 10.6151
R1709 B.n693 B.n692 10.6151
R1710 B.n694 B.n693 10.6151
R1711 B.n695 B.n694 10.6151
R1712 B.n697 B.n695 10.6151
R1713 B.n698 B.n697 10.6151
R1714 B.n699 B.n698 10.6151
R1715 B.n700 B.n699 10.6151
R1716 B.n702 B.n700 10.6151
R1717 B.n703 B.n702 10.6151
R1718 B.n704 B.n703 10.6151
R1719 B.n705 B.n704 10.6151
R1720 B.n707 B.n705 10.6151
R1721 B.n708 B.n707 10.6151
R1722 B.n709 B.n708 10.6151
R1723 B.n710 B.n709 10.6151
R1724 B.n712 B.n710 10.6151
R1725 B.n713 B.n712 10.6151
R1726 B.n714 B.n713 10.6151
R1727 B.n715 B.n714 10.6151
R1728 B.n717 B.n715 10.6151
R1729 B.n718 B.n717 10.6151
R1730 B.n719 B.n718 10.6151
R1731 B.n720 B.n719 10.6151
R1732 B.n722 B.n720 10.6151
R1733 B.n723 B.n722 10.6151
R1734 B.n724 B.n723 10.6151
R1735 B.n725 B.n724 10.6151
R1736 B.n727 B.n725 10.6151
R1737 B.n728 B.n727 10.6151
R1738 B.n729 B.n728 10.6151
R1739 B.n730 B.n729 10.6151
R1740 B.n732 B.n730 10.6151
R1741 B.n733 B.n732 10.6151
R1742 B.n734 B.n733 10.6151
R1743 B.n735 B.n734 10.6151
R1744 B.n737 B.n735 10.6151
R1745 B.n738 B.n737 10.6151
R1746 B.n739 B.n738 10.6151
R1747 B.n740 B.n739 10.6151
R1748 B.n742 B.n740 10.6151
R1749 B.n743 B.n742 10.6151
R1750 B.n744 B.n743 10.6151
R1751 B.n745 B.n744 10.6151
R1752 B.n747 B.n745 10.6151
R1753 B.n748 B.n747 10.6151
R1754 B.n749 B.n748 10.6151
R1755 B.n750 B.n749 10.6151
R1756 B.n752 B.n750 10.6151
R1757 B.n753 B.n752 10.6151
R1758 B.n754 B.n753 10.6151
R1759 B.n755 B.n754 10.6151
R1760 B.n757 B.n755 10.6151
R1761 B.n758 B.n757 10.6151
R1762 B.n759 B.n758 10.6151
R1763 B.n760 B.n759 10.6151
R1764 B.n762 B.n760 10.6151
R1765 B.n763 B.n762 10.6151
R1766 B.n764 B.n763 10.6151
R1767 B.n765 B.n764 10.6151
R1768 B.n767 B.n765 10.6151
R1769 B.n768 B.n767 10.6151
R1770 B.n769 B.n768 10.6151
R1771 B.n770 B.n769 10.6151
R1772 B.n772 B.n770 10.6151
R1773 B.n773 B.n772 10.6151
R1774 B.n774 B.n773 10.6151
R1775 B.n919 B.n1 10.6151
R1776 B.n919 B.n918 10.6151
R1777 B.n918 B.n917 10.6151
R1778 B.n917 B.n10 10.6151
R1779 B.n911 B.n10 10.6151
R1780 B.n911 B.n910 10.6151
R1781 B.n910 B.n909 10.6151
R1782 B.n909 B.n17 10.6151
R1783 B.n903 B.n17 10.6151
R1784 B.n903 B.n902 10.6151
R1785 B.n902 B.n901 10.6151
R1786 B.n901 B.n25 10.6151
R1787 B.n895 B.n25 10.6151
R1788 B.n895 B.n894 10.6151
R1789 B.n894 B.n893 10.6151
R1790 B.n893 B.n32 10.6151
R1791 B.n887 B.n32 10.6151
R1792 B.n887 B.n886 10.6151
R1793 B.n886 B.n885 10.6151
R1794 B.n885 B.n39 10.6151
R1795 B.n879 B.n39 10.6151
R1796 B.n879 B.n878 10.6151
R1797 B.n878 B.n877 10.6151
R1798 B.n877 B.n46 10.6151
R1799 B.n871 B.n46 10.6151
R1800 B.n871 B.n870 10.6151
R1801 B.n870 B.n869 10.6151
R1802 B.n869 B.n53 10.6151
R1803 B.n863 B.n53 10.6151
R1804 B.n863 B.n862 10.6151
R1805 B.n862 B.n861 10.6151
R1806 B.n861 B.n60 10.6151
R1807 B.n855 B.n60 10.6151
R1808 B.n855 B.n854 10.6151
R1809 B.n854 B.n853 10.6151
R1810 B.n853 B.n67 10.6151
R1811 B.n847 B.n67 10.6151
R1812 B.n847 B.n846 10.6151
R1813 B.n846 B.n845 10.6151
R1814 B.n845 B.n74 10.6151
R1815 B.n839 B.n74 10.6151
R1816 B.n839 B.n838 10.6151
R1817 B.n838 B.n837 10.6151
R1818 B.n837 B.n81 10.6151
R1819 B.n831 B.n81 10.6151
R1820 B.n831 B.n830 10.6151
R1821 B.n830 B.n829 10.6151
R1822 B.n829 B.n88 10.6151
R1823 B.n823 B.n88 10.6151
R1824 B.n823 B.n822 10.6151
R1825 B.n822 B.n821 10.6151
R1826 B.n821 B.n94 10.6151
R1827 B.n815 B.n94 10.6151
R1828 B.n815 B.n814 10.6151
R1829 B.n814 B.n813 10.6151
R1830 B.n813 B.n102 10.6151
R1831 B.n807 B.n102 10.6151
R1832 B.n807 B.n806 10.6151
R1833 B.n806 B.n805 10.6151
R1834 B.n805 B.n109 10.6151
R1835 B.n799 B.n109 10.6151
R1836 B.n799 B.n798 10.6151
R1837 B.n798 B.n797 10.6151
R1838 B.n797 B.n116 10.6151
R1839 B.n791 B.n116 10.6151
R1840 B.n791 B.n790 10.6151
R1841 B.n790 B.n789 10.6151
R1842 B.n789 B.n123 10.6151
R1843 B.n783 B.n123 10.6151
R1844 B.n783 B.n782 10.6151
R1845 B.n782 B.n781 10.6151
R1846 B.n781 B.n130 10.6151
R1847 B.n159 B.n158 10.6151
R1848 B.n162 B.n159 10.6151
R1849 B.n163 B.n162 10.6151
R1850 B.n166 B.n163 10.6151
R1851 B.n167 B.n166 10.6151
R1852 B.n170 B.n167 10.6151
R1853 B.n171 B.n170 10.6151
R1854 B.n174 B.n171 10.6151
R1855 B.n175 B.n174 10.6151
R1856 B.n178 B.n175 10.6151
R1857 B.n179 B.n178 10.6151
R1858 B.n182 B.n179 10.6151
R1859 B.n187 B.n184 10.6151
R1860 B.n188 B.n187 10.6151
R1861 B.n191 B.n188 10.6151
R1862 B.n192 B.n191 10.6151
R1863 B.n195 B.n192 10.6151
R1864 B.n196 B.n195 10.6151
R1865 B.n199 B.n196 10.6151
R1866 B.n200 B.n199 10.6151
R1867 B.n204 B.n203 10.6151
R1868 B.n207 B.n204 10.6151
R1869 B.n208 B.n207 10.6151
R1870 B.n211 B.n208 10.6151
R1871 B.n212 B.n211 10.6151
R1872 B.n215 B.n212 10.6151
R1873 B.n216 B.n215 10.6151
R1874 B.n219 B.n216 10.6151
R1875 B.n220 B.n219 10.6151
R1876 B.n223 B.n220 10.6151
R1877 B.n224 B.n223 10.6151
R1878 B.n775 B.n224 10.6151
R1879 B.n927 B.n0 8.11757
R1880 B.n927 B.n1 8.11757
R1881 B.n430 B.n388 6.5566
R1882 B.n414 B.n413 6.5566
R1883 B.n184 B.n183 6.5566
R1884 B.n200 B.n154 6.5566
R1885 B.n433 B.n388 4.05904
R1886 B.n413 B.n412 4.05904
R1887 B.n183 B.n182 4.05904
R1888 B.n203 B.n154 4.05904
R1889 VN.n98 VN.n97 161.3
R1890 VN.n96 VN.n51 161.3
R1891 VN.n95 VN.n94 161.3
R1892 VN.n93 VN.n52 161.3
R1893 VN.n92 VN.n91 161.3
R1894 VN.n90 VN.n53 161.3
R1895 VN.n89 VN.n88 161.3
R1896 VN.n87 VN.n54 161.3
R1897 VN.n86 VN.n85 161.3
R1898 VN.n84 VN.n55 161.3
R1899 VN.n83 VN.n82 161.3
R1900 VN.n81 VN.n57 161.3
R1901 VN.n80 VN.n79 161.3
R1902 VN.n78 VN.n58 161.3
R1903 VN.n77 VN.n76 161.3
R1904 VN.n75 VN.n74 161.3
R1905 VN.n73 VN.n60 161.3
R1906 VN.n72 VN.n71 161.3
R1907 VN.n70 VN.n61 161.3
R1908 VN.n69 VN.n68 161.3
R1909 VN.n67 VN.n62 161.3
R1910 VN.n66 VN.n65 161.3
R1911 VN.n48 VN.n47 161.3
R1912 VN.n46 VN.n1 161.3
R1913 VN.n45 VN.n44 161.3
R1914 VN.n43 VN.n2 161.3
R1915 VN.n42 VN.n41 161.3
R1916 VN.n40 VN.n3 161.3
R1917 VN.n39 VN.n38 161.3
R1918 VN.n37 VN.n4 161.3
R1919 VN.n36 VN.n35 161.3
R1920 VN.n33 VN.n5 161.3
R1921 VN.n32 VN.n31 161.3
R1922 VN.n30 VN.n6 161.3
R1923 VN.n29 VN.n28 161.3
R1924 VN.n27 VN.n7 161.3
R1925 VN.n26 VN.n25 161.3
R1926 VN.n24 VN.n23 161.3
R1927 VN.n22 VN.n9 161.3
R1928 VN.n21 VN.n20 161.3
R1929 VN.n19 VN.n10 161.3
R1930 VN.n18 VN.n17 161.3
R1931 VN.n16 VN.n11 161.3
R1932 VN.n15 VN.n14 161.3
R1933 VN.n49 VN.n0 80.6405
R1934 VN.n99 VN.n50 80.6405
R1935 VN.n41 VN.n2 56.4773
R1936 VN.n91 VN.n52 56.4773
R1937 VN.n13 VN.n12 51.4682
R1938 VN.n64 VN.n63 51.4682
R1939 VN.n17 VN.n10 51.1217
R1940 VN.n32 VN.n6 51.1217
R1941 VN.n68 VN.n61 51.1217
R1942 VN.n83 VN.n57 51.1217
R1943 VN VN.n99 50.1873
R1944 VN.n64 VN.t5 48.6974
R1945 VN.n13 VN.t3 48.6974
R1946 VN.n21 VN.n10 29.6995
R1947 VN.n28 VN.n6 29.6995
R1948 VN.n72 VN.n61 29.6995
R1949 VN.n79 VN.n57 29.6995
R1950 VN.n16 VN.n15 24.3439
R1951 VN.n17 VN.n16 24.3439
R1952 VN.n22 VN.n21 24.3439
R1953 VN.n23 VN.n22 24.3439
R1954 VN.n27 VN.n26 24.3439
R1955 VN.n28 VN.n27 24.3439
R1956 VN.n33 VN.n32 24.3439
R1957 VN.n35 VN.n33 24.3439
R1958 VN.n39 VN.n4 24.3439
R1959 VN.n40 VN.n39 24.3439
R1960 VN.n41 VN.n40 24.3439
R1961 VN.n45 VN.n2 24.3439
R1962 VN.n46 VN.n45 24.3439
R1963 VN.n47 VN.n46 24.3439
R1964 VN.n68 VN.n67 24.3439
R1965 VN.n67 VN.n66 24.3439
R1966 VN.n79 VN.n78 24.3439
R1967 VN.n78 VN.n77 24.3439
R1968 VN.n74 VN.n73 24.3439
R1969 VN.n73 VN.n72 24.3439
R1970 VN.n91 VN.n90 24.3439
R1971 VN.n90 VN.n89 24.3439
R1972 VN.n89 VN.n54 24.3439
R1973 VN.n85 VN.n84 24.3439
R1974 VN.n84 VN.n83 24.3439
R1975 VN.n97 VN.n96 24.3439
R1976 VN.n96 VN.n95 24.3439
R1977 VN.n95 VN.n52 24.3439
R1978 VN.n15 VN.n12 22.8833
R1979 VN.n35 VN.n34 22.8833
R1980 VN.n66 VN.n63 22.8833
R1981 VN.n85 VN.n56 22.8833
R1982 VN.n12 VN.t8 15.4984
R1983 VN.n8 VN.t9 15.4984
R1984 VN.n34 VN.t6 15.4984
R1985 VN.n0 VN.t7 15.4984
R1986 VN.n63 VN.t2 15.4984
R1987 VN.n59 VN.t1 15.4984
R1988 VN.n56 VN.t4 15.4984
R1989 VN.n50 VN.t0 15.4984
R1990 VN.n23 VN.n8 12.1722
R1991 VN.n26 VN.n8 12.1722
R1992 VN.n77 VN.n59 12.1722
R1993 VN.n74 VN.n59 12.1722
R1994 VN.n47 VN.n0 9.251
R1995 VN.n97 VN.n50 9.251
R1996 VN.n14 VN.n13 3.19274
R1997 VN.n65 VN.n64 3.19274
R1998 VN.n34 VN.n4 1.46111
R1999 VN.n56 VN.n54 1.46111
R2000 VN.n99 VN.n98 0.355081
R2001 VN.n49 VN.n48 0.355081
R2002 VN VN.n49 0.26685
R2003 VN.n98 VN.n51 0.189894
R2004 VN.n94 VN.n51 0.189894
R2005 VN.n94 VN.n93 0.189894
R2006 VN.n93 VN.n92 0.189894
R2007 VN.n92 VN.n53 0.189894
R2008 VN.n88 VN.n53 0.189894
R2009 VN.n88 VN.n87 0.189894
R2010 VN.n87 VN.n86 0.189894
R2011 VN.n86 VN.n55 0.189894
R2012 VN.n82 VN.n55 0.189894
R2013 VN.n82 VN.n81 0.189894
R2014 VN.n81 VN.n80 0.189894
R2015 VN.n80 VN.n58 0.189894
R2016 VN.n76 VN.n58 0.189894
R2017 VN.n76 VN.n75 0.189894
R2018 VN.n75 VN.n60 0.189894
R2019 VN.n71 VN.n60 0.189894
R2020 VN.n71 VN.n70 0.189894
R2021 VN.n70 VN.n69 0.189894
R2022 VN.n69 VN.n62 0.189894
R2023 VN.n65 VN.n62 0.189894
R2024 VN.n14 VN.n11 0.189894
R2025 VN.n18 VN.n11 0.189894
R2026 VN.n19 VN.n18 0.189894
R2027 VN.n20 VN.n19 0.189894
R2028 VN.n20 VN.n9 0.189894
R2029 VN.n24 VN.n9 0.189894
R2030 VN.n25 VN.n24 0.189894
R2031 VN.n25 VN.n7 0.189894
R2032 VN.n29 VN.n7 0.189894
R2033 VN.n30 VN.n29 0.189894
R2034 VN.n31 VN.n30 0.189894
R2035 VN.n31 VN.n5 0.189894
R2036 VN.n36 VN.n5 0.189894
R2037 VN.n37 VN.n36 0.189894
R2038 VN.n38 VN.n37 0.189894
R2039 VN.n38 VN.n3 0.189894
R2040 VN.n42 VN.n3 0.189894
R2041 VN.n43 VN.n42 0.189894
R2042 VN.n44 VN.n43 0.189894
R2043 VN.n44 VN.n1 0.189894
R2044 VN.n48 VN.n1 0.189894
R2045 VDD2.n1 VDD2.t6 105.757
R2046 VDD2.n4 VDD2.t9 102.55
R2047 VDD2.n3 VDD2.n2 95.8172
R2048 VDD2 VDD2.n7 95.8146
R2049 VDD2.n6 VDD2.n5 93.4677
R2050 VDD2.n1 VDD2.n0 93.4674
R2051 VDD2.n4 VDD2.n3 40.8274
R2052 VDD2.n7 VDD2.t7 9.08307
R2053 VDD2.n7 VDD2.t4 9.08307
R2054 VDD2.n5 VDD2.t5 9.08307
R2055 VDD2.n5 VDD2.t8 9.08307
R2056 VDD2.n2 VDD2.t3 9.08307
R2057 VDD2.n2 VDD2.t2 9.08307
R2058 VDD2.n0 VDD2.t1 9.08307
R2059 VDD2.n0 VDD2.t0 9.08307
R2060 VDD2.n6 VDD2.n4 3.2074
R2061 VDD2 VDD2.n6 0.860414
R2062 VDD2.n3 VDD2.n1 0.746878
C0 VP VTAIL 4.32218f
C1 VDD1 VTAIL 6.73445f
C2 VDD2 VTAIL 6.79312f
C3 VP VDD1 3.00181f
C4 VP VDD2 0.691116f
C5 VDD1 VDD2 2.6886f
C6 VN VTAIL 4.30805f
C7 VP VN 7.76369f
C8 VDD1 VN 0.161081f
C9 VDD2 VN 2.47623f
C10 VDD2 B 6.55283f
C11 VDD1 B 6.406865f
C12 VTAIL B 4.227341f
C13 VN B 21.18586f
C14 VP B 19.50872f
C15 VDD2.t6 B 0.471776f
C16 VDD2.t1 B 0.051773f
C17 VDD2.t0 B 0.051773f
C18 VDD2.n0 B 0.352135f
C19 VDD2.n1 B 1.16192f
C20 VDD2.t3 B 0.051773f
C21 VDD2.t2 B 0.051773f
C22 VDD2.n2 B 0.370957f
C23 VDD2.n3 B 3.2498f
C24 VDD2.t9 B 0.454228f
C25 VDD2.n4 B 3.13247f
C26 VDD2.t5 B 0.051773f
C27 VDD2.t8 B 0.051773f
C28 VDD2.n5 B 0.352136f
C29 VDD2.n6 B 0.610797f
C30 VDD2.t7 B 0.051773f
C31 VDD2.t4 B 0.051773f
C32 VDD2.n7 B 0.37092f
C33 VN.t7 B 0.461779f
C34 VN.n0 B 0.304259f
C35 VN.n1 B 0.026321f
C36 VN.n2 B 0.032682f
C37 VN.n3 B 0.026321f
C38 VN.n4 B 0.02642f
C39 VN.n5 B 0.026321f
C40 VN.n6 B 0.025732f
C41 VN.n7 B 0.026321f
C42 VN.t9 B 0.461779f
C43 VN.n8 B 0.206053f
C44 VN.n9 B 0.026321f
C45 VN.n10 B 0.025732f
C46 VN.n11 B 0.026321f
C47 VN.t8 B 0.461779f
C48 VN.n12 B 0.3085f
C49 VN.t3 B 0.73474f
C50 VN.n13 B 0.315363f
C51 VN.n14 B 0.322339f
C52 VN.n15 B 0.047841f
C53 VN.n16 B 0.049302f
C54 VN.n17 B 0.048027f
C55 VN.n18 B 0.026321f
C56 VN.n19 B 0.026321f
C57 VN.n20 B 0.026321f
C58 VN.n21 B 0.052726f
C59 VN.n22 B 0.049302f
C60 VN.n23 B 0.037131f
C61 VN.n24 B 0.026321f
C62 VN.n25 B 0.026321f
C63 VN.n26 B 0.037131f
C64 VN.n27 B 0.049302f
C65 VN.n28 B 0.052726f
C66 VN.n29 B 0.026321f
C67 VN.n30 B 0.026321f
C68 VN.n31 B 0.026321f
C69 VN.n32 B 0.048027f
C70 VN.n33 B 0.049302f
C71 VN.t6 B 0.461779f
C72 VN.n34 B 0.206053f
C73 VN.n35 B 0.047841f
C74 VN.n36 B 0.026321f
C75 VN.n37 B 0.026321f
C76 VN.n38 B 0.026321f
C77 VN.n39 B 0.049302f
C78 VN.n40 B 0.049302f
C79 VN.n41 B 0.044501f
C80 VN.n42 B 0.026321f
C81 VN.n43 B 0.026321f
C82 VN.n44 B 0.026321f
C83 VN.n45 B 0.049302f
C84 VN.n46 B 0.049302f
C85 VN.n47 B 0.03421f
C86 VN.n48 B 0.042489f
C87 VN.n49 B 0.070023f
C88 VN.t0 B 0.461779f
C89 VN.n50 B 0.304259f
C90 VN.n51 B 0.026321f
C91 VN.n52 B 0.032682f
C92 VN.n53 B 0.026321f
C93 VN.n54 B 0.02642f
C94 VN.n55 B 0.026321f
C95 VN.t4 B 0.461779f
C96 VN.n56 B 0.206053f
C97 VN.n57 B 0.025732f
C98 VN.n58 B 0.026321f
C99 VN.t1 B 0.461779f
C100 VN.n59 B 0.206053f
C101 VN.n60 B 0.026321f
C102 VN.n61 B 0.025732f
C103 VN.n62 B 0.026321f
C104 VN.t2 B 0.461779f
C105 VN.n63 B 0.3085f
C106 VN.t5 B 0.73474f
C107 VN.n64 B 0.315363f
C108 VN.n65 B 0.322339f
C109 VN.n66 B 0.047841f
C110 VN.n67 B 0.049302f
C111 VN.n68 B 0.048027f
C112 VN.n69 B 0.026321f
C113 VN.n70 B 0.026321f
C114 VN.n71 B 0.026321f
C115 VN.n72 B 0.052726f
C116 VN.n73 B 0.049302f
C117 VN.n74 B 0.037131f
C118 VN.n75 B 0.026321f
C119 VN.n76 B 0.026321f
C120 VN.n77 B 0.037131f
C121 VN.n78 B 0.049302f
C122 VN.n79 B 0.052726f
C123 VN.n80 B 0.026321f
C124 VN.n81 B 0.026321f
C125 VN.n82 B 0.026321f
C126 VN.n83 B 0.048027f
C127 VN.n84 B 0.049302f
C128 VN.n85 B 0.047841f
C129 VN.n86 B 0.026321f
C130 VN.n87 B 0.026321f
C131 VN.n88 B 0.026321f
C132 VN.n89 B 0.049302f
C133 VN.n90 B 0.049302f
C134 VN.n91 B 0.044501f
C135 VN.n92 B 0.026321f
C136 VN.n93 B 0.026321f
C137 VN.n94 B 0.026321f
C138 VN.n95 B 0.049302f
C139 VN.n96 B 0.049302f
C140 VN.n97 B 0.03421f
C141 VN.n98 B 0.042489f
C142 VN.n99 B 1.51437f
C143 VTAIL.t5 B 0.06454f
C144 VTAIL.t2 B 0.06454f
C145 VTAIL.n0 B 0.381767f
C146 VTAIL.n1 B 0.824403f
C147 VTAIL.t17 B 0.505613f
C148 VTAIL.n2 B 0.966333f
C149 VTAIL.t15 B 0.06454f
C150 VTAIL.t16 B 0.06454f
C151 VTAIL.n3 B 0.381767f
C152 VTAIL.n4 B 1.05101f
C153 VTAIL.t10 B 0.06454f
C154 VTAIL.t12 B 0.06454f
C155 VTAIL.n5 B 0.381767f
C156 VTAIL.n6 B 2.17392f
C157 VTAIL.t1 B 0.06454f
C158 VTAIL.t8 B 0.06454f
C159 VTAIL.n7 B 0.381768f
C160 VTAIL.n8 B 2.17392f
C161 VTAIL.t3 B 0.06454f
C162 VTAIL.t4 B 0.06454f
C163 VTAIL.n9 B 0.381768f
C164 VTAIL.n10 B 1.05101f
C165 VTAIL.t0 B 0.505616f
C166 VTAIL.n11 B 0.96633f
C167 VTAIL.t13 B 0.06454f
C168 VTAIL.t18 B 0.06454f
C169 VTAIL.n12 B 0.381768f
C170 VTAIL.n13 B 0.91416f
C171 VTAIL.t11 B 0.06454f
C172 VTAIL.t19 B 0.06454f
C173 VTAIL.n14 B 0.381768f
C174 VTAIL.n15 B 1.05101f
C175 VTAIL.t14 B 0.505613f
C176 VTAIL.n16 B 1.83896f
C177 VTAIL.t7 B 0.505613f
C178 VTAIL.n17 B 1.83896f
C179 VTAIL.t6 B 0.06454f
C180 VTAIL.t9 B 0.06454f
C181 VTAIL.n18 B 0.381767f
C182 VTAIL.n19 B 0.753637f
C183 VDD1.t8 B 0.483035f
C184 VDD1.t2 B 0.053009f
C185 VDD1.t4 B 0.053009f
C186 VDD1.n0 B 0.360538f
C187 VDD1.n1 B 1.19995f
C188 VDD1.t1 B 0.483033f
C189 VDD1.t5 B 0.053009f
C190 VDD1.t0 B 0.053009f
C191 VDD1.n2 B 0.360538f
C192 VDD1.n3 B 1.18965f
C193 VDD1.t9 B 0.053009f
C194 VDD1.t3 B 0.053009f
C195 VDD1.n4 B 0.379809f
C196 VDD1.n5 B 3.49581f
C197 VDD1.t7 B 0.053009f
C198 VDD1.t6 B 0.053009f
C199 VDD1.n6 B 0.360537f
C200 VDD1.n7 B 3.34507f
C201 VP.t2 B 0.478807f
C202 VP.n0 B 0.315479f
C203 VP.n1 B 0.027292f
C204 VP.n2 B 0.033887f
C205 VP.n3 B 0.027292f
C206 VP.n4 B 0.027395f
C207 VP.n5 B 0.027292f
C208 VP.n6 B 0.026681f
C209 VP.n7 B 0.027292f
C210 VP.t4 B 0.478807f
C211 VP.n8 B 0.213651f
C212 VP.n9 B 0.027292f
C213 VP.n10 B 0.026681f
C214 VP.n11 B 0.027292f
C215 VP.t7 B 0.478807f
C216 VP.n12 B 0.213651f
C217 VP.n13 B 0.027292f
C218 VP.n14 B 0.046142f
C219 VP.n15 B 0.027292f
C220 VP.n16 B 0.035471f
C221 VP.t5 B 0.478807f
C222 VP.n17 B 0.315479f
C223 VP.n18 B 0.027292f
C224 VP.n19 B 0.033887f
C225 VP.n20 B 0.027292f
C226 VP.n21 B 0.027395f
C227 VP.n22 B 0.027292f
C228 VP.n23 B 0.026681f
C229 VP.n24 B 0.027292f
C230 VP.t8 B 0.478807f
C231 VP.n25 B 0.213651f
C232 VP.n26 B 0.027292f
C233 VP.n27 B 0.026681f
C234 VP.n28 B 0.027292f
C235 VP.t1 B 0.478807f
C236 VP.n29 B 0.319876f
C237 VP.t6 B 0.761832f
C238 VP.n30 B 0.326992f
C239 VP.n31 B 0.334226f
C240 VP.n32 B 0.049605f
C241 VP.n33 B 0.05112f
C242 VP.n34 B 0.049798f
C243 VP.n35 B 0.027292f
C244 VP.n36 B 0.027292f
C245 VP.n37 B 0.027292f
C246 VP.n38 B 0.05467f
C247 VP.n39 B 0.05112f
C248 VP.n40 B 0.0385f
C249 VP.n41 B 0.027292f
C250 VP.n42 B 0.027292f
C251 VP.n43 B 0.0385f
C252 VP.n44 B 0.05112f
C253 VP.n45 B 0.05467f
C254 VP.n46 B 0.027292f
C255 VP.n47 B 0.027292f
C256 VP.n48 B 0.027292f
C257 VP.n49 B 0.049798f
C258 VP.n50 B 0.05112f
C259 VP.t0 B 0.478807f
C260 VP.n51 B 0.213651f
C261 VP.n52 B 0.049605f
C262 VP.n53 B 0.027292f
C263 VP.n54 B 0.027292f
C264 VP.n55 B 0.027292f
C265 VP.n56 B 0.05112f
C266 VP.n57 B 0.05112f
C267 VP.n58 B 0.046142f
C268 VP.n59 B 0.027292f
C269 VP.n60 B 0.027292f
C270 VP.n61 B 0.027292f
C271 VP.n62 B 0.05112f
C272 VP.n63 B 0.05112f
C273 VP.n64 B 0.035471f
C274 VP.n65 B 0.044055f
C275 VP.n66 B 1.55904f
C276 VP.t9 B 0.478807f
C277 VP.n67 B 0.315479f
C278 VP.n68 B 1.57859f
C279 VP.n69 B 0.044055f
C280 VP.n70 B 0.027292f
C281 VP.n71 B 0.05112f
C282 VP.n72 B 0.05112f
C283 VP.n73 B 0.033887f
C284 VP.n74 B 0.027292f
C285 VP.n75 B 0.027292f
C286 VP.n76 B 0.027292f
C287 VP.n77 B 0.05112f
C288 VP.n78 B 0.05112f
C289 VP.n79 B 0.027395f
C290 VP.n80 B 0.027292f
C291 VP.n81 B 0.027292f
C292 VP.n82 B 0.049605f
C293 VP.n83 B 0.05112f
C294 VP.n84 B 0.049798f
C295 VP.n85 B 0.027292f
C296 VP.n86 B 0.027292f
C297 VP.n87 B 0.027292f
C298 VP.n88 B 0.05467f
C299 VP.n89 B 0.05112f
C300 VP.n90 B 0.0385f
C301 VP.n91 B 0.027292f
C302 VP.n92 B 0.027292f
C303 VP.n93 B 0.0385f
C304 VP.n94 B 0.05112f
C305 VP.n95 B 0.05467f
C306 VP.n96 B 0.027292f
C307 VP.n97 B 0.027292f
C308 VP.n98 B 0.027292f
C309 VP.n99 B 0.049798f
C310 VP.n100 B 0.05112f
C311 VP.t3 B 0.478807f
C312 VP.n101 B 0.213651f
C313 VP.n102 B 0.049605f
C314 VP.n103 B 0.027292f
C315 VP.n104 B 0.027292f
C316 VP.n105 B 0.027292f
C317 VP.n106 B 0.05112f
C318 VP.n107 B 0.05112f
C319 VP.n108 B 0.046142f
C320 VP.n109 B 0.027292f
C321 VP.n110 B 0.027292f
C322 VP.n111 B 0.027292f
C323 VP.n112 B 0.05112f
C324 VP.n113 B 0.05112f
C325 VP.n114 B 0.035471f
C326 VP.n115 B 0.044055f
C327 VP.n116 B 0.072605f
.ends

