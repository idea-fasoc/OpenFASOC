* NGSPICE file created from diff_pair_sample_0997.ext - technology: sky130A

.subckt diff_pair_sample_0997 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t18 VP.t0 VDD1.t9 w_n4594_n3194# sky130_fd_pr__pfet_01v8 ad=1.83645 pd=11.46 as=1.83645 ps=11.46 w=11.13 l=2.69
X1 B.t11 B.t9 B.t10 w_n4594_n3194# sky130_fd_pr__pfet_01v8 ad=4.3407 pd=23.04 as=0 ps=0 w=11.13 l=2.69
X2 B.t8 B.t6 B.t7 w_n4594_n3194# sky130_fd_pr__pfet_01v8 ad=4.3407 pd=23.04 as=0 ps=0 w=11.13 l=2.69
X3 VTAIL.t17 VP.t1 VDD1.t0 w_n4594_n3194# sky130_fd_pr__pfet_01v8 ad=1.83645 pd=11.46 as=1.83645 ps=11.46 w=11.13 l=2.69
X4 B.t5 B.t3 B.t4 w_n4594_n3194# sky130_fd_pr__pfet_01v8 ad=4.3407 pd=23.04 as=0 ps=0 w=11.13 l=2.69
X5 VDD1.t6 VP.t2 VTAIL.t16 w_n4594_n3194# sky130_fd_pr__pfet_01v8 ad=1.83645 pd=11.46 as=1.83645 ps=11.46 w=11.13 l=2.69
X6 VTAIL.t19 VN.t0 VDD2.t9 w_n4594_n3194# sky130_fd_pr__pfet_01v8 ad=1.83645 pd=11.46 as=1.83645 ps=11.46 w=11.13 l=2.69
X7 VDD1.t2 VP.t3 VTAIL.t15 w_n4594_n3194# sky130_fd_pr__pfet_01v8 ad=4.3407 pd=23.04 as=1.83645 ps=11.46 w=11.13 l=2.69
X8 VTAIL.t14 VP.t4 VDD1.t1 w_n4594_n3194# sky130_fd_pr__pfet_01v8 ad=1.83645 pd=11.46 as=1.83645 ps=11.46 w=11.13 l=2.69
X9 B.t2 B.t0 B.t1 w_n4594_n3194# sky130_fd_pr__pfet_01v8 ad=4.3407 pd=23.04 as=0 ps=0 w=11.13 l=2.69
X10 VDD2.t8 VN.t1 VTAIL.t4 w_n4594_n3194# sky130_fd_pr__pfet_01v8 ad=1.83645 pd=11.46 as=1.83645 ps=11.46 w=11.13 l=2.69
X11 VTAIL.t8 VN.t2 VDD2.t7 w_n4594_n3194# sky130_fd_pr__pfet_01v8 ad=1.83645 pd=11.46 as=1.83645 ps=11.46 w=11.13 l=2.69
X12 VDD2.t6 VN.t3 VTAIL.t6 w_n4594_n3194# sky130_fd_pr__pfet_01v8 ad=1.83645 pd=11.46 as=4.3407 ps=23.04 w=11.13 l=2.69
X13 VTAIL.t3 VN.t4 VDD2.t5 w_n4594_n3194# sky130_fd_pr__pfet_01v8 ad=1.83645 pd=11.46 as=1.83645 ps=11.46 w=11.13 l=2.69
X14 VDD1.t7 VP.t5 VTAIL.t13 w_n4594_n3194# sky130_fd_pr__pfet_01v8 ad=4.3407 pd=23.04 as=1.83645 ps=11.46 w=11.13 l=2.69
X15 VDD2.t4 VN.t5 VTAIL.t1 w_n4594_n3194# sky130_fd_pr__pfet_01v8 ad=4.3407 pd=23.04 as=1.83645 ps=11.46 w=11.13 l=2.69
X16 VDD1.t5 VP.t6 VTAIL.t12 w_n4594_n3194# sky130_fd_pr__pfet_01v8 ad=1.83645 pd=11.46 as=4.3407 ps=23.04 w=11.13 l=2.69
X17 VTAIL.t7 VN.t6 VDD2.t3 w_n4594_n3194# sky130_fd_pr__pfet_01v8 ad=1.83645 pd=11.46 as=1.83645 ps=11.46 w=11.13 l=2.69
X18 VDD2.t2 VN.t7 VTAIL.t2 w_n4594_n3194# sky130_fd_pr__pfet_01v8 ad=1.83645 pd=11.46 as=1.83645 ps=11.46 w=11.13 l=2.69
X19 VDD2.t1 VN.t8 VTAIL.t5 w_n4594_n3194# sky130_fd_pr__pfet_01v8 ad=1.83645 pd=11.46 as=4.3407 ps=23.04 w=11.13 l=2.69
X20 VDD1.t8 VP.t7 VTAIL.t11 w_n4594_n3194# sky130_fd_pr__pfet_01v8 ad=1.83645 pd=11.46 as=4.3407 ps=23.04 w=11.13 l=2.69
X21 VTAIL.t10 VP.t8 VDD1.t3 w_n4594_n3194# sky130_fd_pr__pfet_01v8 ad=1.83645 pd=11.46 as=1.83645 ps=11.46 w=11.13 l=2.69
X22 VDD1.t4 VP.t9 VTAIL.t9 w_n4594_n3194# sky130_fd_pr__pfet_01v8 ad=1.83645 pd=11.46 as=1.83645 ps=11.46 w=11.13 l=2.69
X23 VDD2.t0 VN.t9 VTAIL.t0 w_n4594_n3194# sky130_fd_pr__pfet_01v8 ad=4.3407 pd=23.04 as=1.83645 ps=11.46 w=11.13 l=2.69
R0 VP.n27 VP.n26 161.3
R1 VP.n28 VP.n23 161.3
R2 VP.n30 VP.n29 161.3
R3 VP.n31 VP.n22 161.3
R4 VP.n33 VP.n32 161.3
R5 VP.n34 VP.n21 161.3
R6 VP.n36 VP.n35 161.3
R7 VP.n37 VP.n20 161.3
R8 VP.n39 VP.n38 161.3
R9 VP.n40 VP.n19 161.3
R10 VP.n42 VP.n41 161.3
R11 VP.n43 VP.n18 161.3
R12 VP.n45 VP.n44 161.3
R13 VP.n47 VP.n46 161.3
R14 VP.n48 VP.n16 161.3
R15 VP.n50 VP.n49 161.3
R16 VP.n51 VP.n15 161.3
R17 VP.n53 VP.n52 161.3
R18 VP.n54 VP.n14 161.3
R19 VP.n96 VP.n0 161.3
R20 VP.n95 VP.n94 161.3
R21 VP.n93 VP.n1 161.3
R22 VP.n92 VP.n91 161.3
R23 VP.n90 VP.n2 161.3
R24 VP.n89 VP.n88 161.3
R25 VP.n87 VP.n86 161.3
R26 VP.n85 VP.n4 161.3
R27 VP.n84 VP.n83 161.3
R28 VP.n82 VP.n5 161.3
R29 VP.n81 VP.n80 161.3
R30 VP.n79 VP.n6 161.3
R31 VP.n78 VP.n77 161.3
R32 VP.n76 VP.n7 161.3
R33 VP.n75 VP.n74 161.3
R34 VP.n73 VP.n8 161.3
R35 VP.n72 VP.n71 161.3
R36 VP.n70 VP.n9 161.3
R37 VP.n69 VP.n68 161.3
R38 VP.n66 VP.n10 161.3
R39 VP.n65 VP.n64 161.3
R40 VP.n63 VP.n11 161.3
R41 VP.n62 VP.n61 161.3
R42 VP.n60 VP.n12 161.3
R43 VP.n59 VP.n58 161.3
R44 VP.n24 VP.t5 130.427
R45 VP.n57 VP.n13 108.799
R46 VP.n98 VP.n97 108.799
R47 VP.n56 VP.n55 108.799
R48 VP.n78 VP.t9 99.7154
R49 VP.n13 VP.t3 99.7154
R50 VP.n67 VP.t1 99.7154
R51 VP.n3 VP.t0 99.7154
R52 VP.n97 VP.t7 99.7154
R53 VP.n36 VP.t2 99.7154
R54 VP.n55 VP.t6 99.7154
R55 VP.n17 VP.t8 99.7154
R56 VP.n25 VP.t4 99.7154
R57 VP.n25 VP.n24 72.37
R58 VP.n57 VP.n56 52.8632
R59 VP.n61 VP.n11 43.4072
R60 VP.n91 VP.n1 43.4072
R61 VP.n49 VP.n15 43.4072
R62 VP.n73 VP.n72 41.4647
R63 VP.n84 VP.n5 41.4647
R64 VP.n42 VP.n19 41.4647
R65 VP.n31 VP.n30 41.4647
R66 VP.n74 VP.n73 39.5221
R67 VP.n80 VP.n5 39.5221
R68 VP.n38 VP.n19 39.5221
R69 VP.n32 VP.n31 39.5221
R70 VP.n65 VP.n11 37.5796
R71 VP.n91 VP.n90 37.5796
R72 VP.n49 VP.n48 37.5796
R73 VP.n60 VP.n59 24.4675
R74 VP.n61 VP.n60 24.4675
R75 VP.n66 VP.n65 24.4675
R76 VP.n68 VP.n9 24.4675
R77 VP.n72 VP.n9 24.4675
R78 VP.n74 VP.n7 24.4675
R79 VP.n78 VP.n7 24.4675
R80 VP.n79 VP.n78 24.4675
R81 VP.n80 VP.n79 24.4675
R82 VP.n85 VP.n84 24.4675
R83 VP.n86 VP.n85 24.4675
R84 VP.n90 VP.n89 24.4675
R85 VP.n95 VP.n1 24.4675
R86 VP.n96 VP.n95 24.4675
R87 VP.n53 VP.n15 24.4675
R88 VP.n54 VP.n53 24.4675
R89 VP.n43 VP.n42 24.4675
R90 VP.n44 VP.n43 24.4675
R91 VP.n48 VP.n47 24.4675
R92 VP.n32 VP.n21 24.4675
R93 VP.n36 VP.n21 24.4675
R94 VP.n37 VP.n36 24.4675
R95 VP.n38 VP.n37 24.4675
R96 VP.n26 VP.n23 24.4675
R97 VP.n30 VP.n23 24.4675
R98 VP.n67 VP.n66 23.4888
R99 VP.n89 VP.n3 23.4888
R100 VP.n47 VP.n17 23.4888
R101 VP.n27 VP.n24 7.37486
R102 VP.n59 VP.n13 1.95786
R103 VP.n97 VP.n96 1.95786
R104 VP.n55 VP.n54 1.95786
R105 VP.n68 VP.n67 0.97918
R106 VP.n86 VP.n3 0.97918
R107 VP.n44 VP.n17 0.97918
R108 VP.n26 VP.n25 0.97918
R109 VP.n56 VP.n14 0.278367
R110 VP.n58 VP.n57 0.278367
R111 VP.n98 VP.n0 0.278367
R112 VP.n28 VP.n27 0.189894
R113 VP.n29 VP.n28 0.189894
R114 VP.n29 VP.n22 0.189894
R115 VP.n33 VP.n22 0.189894
R116 VP.n34 VP.n33 0.189894
R117 VP.n35 VP.n34 0.189894
R118 VP.n35 VP.n20 0.189894
R119 VP.n39 VP.n20 0.189894
R120 VP.n40 VP.n39 0.189894
R121 VP.n41 VP.n40 0.189894
R122 VP.n41 VP.n18 0.189894
R123 VP.n45 VP.n18 0.189894
R124 VP.n46 VP.n45 0.189894
R125 VP.n46 VP.n16 0.189894
R126 VP.n50 VP.n16 0.189894
R127 VP.n51 VP.n50 0.189894
R128 VP.n52 VP.n51 0.189894
R129 VP.n52 VP.n14 0.189894
R130 VP.n58 VP.n12 0.189894
R131 VP.n62 VP.n12 0.189894
R132 VP.n63 VP.n62 0.189894
R133 VP.n64 VP.n63 0.189894
R134 VP.n64 VP.n10 0.189894
R135 VP.n69 VP.n10 0.189894
R136 VP.n70 VP.n69 0.189894
R137 VP.n71 VP.n70 0.189894
R138 VP.n71 VP.n8 0.189894
R139 VP.n75 VP.n8 0.189894
R140 VP.n76 VP.n75 0.189894
R141 VP.n77 VP.n76 0.189894
R142 VP.n77 VP.n6 0.189894
R143 VP.n81 VP.n6 0.189894
R144 VP.n82 VP.n81 0.189894
R145 VP.n83 VP.n82 0.189894
R146 VP.n83 VP.n4 0.189894
R147 VP.n87 VP.n4 0.189894
R148 VP.n88 VP.n87 0.189894
R149 VP.n88 VP.n2 0.189894
R150 VP.n92 VP.n2 0.189894
R151 VP.n93 VP.n92 0.189894
R152 VP.n94 VP.n93 0.189894
R153 VP.n94 VP.n0 0.189894
R154 VP VP.n98 0.153454
R155 VDD1.n1 VDD1.t7 82.5744
R156 VDD1.n3 VDD1.t2 82.5743
R157 VDD1.n5 VDD1.n4 78.9475
R158 VDD1.n1 VDD1.n0 77.0505
R159 VDD1.n7 VDD1.n6 77.0503
R160 VDD1.n3 VDD1.n2 77.0503
R161 VDD1.n7 VDD1.n5 47.5612
R162 VDD1.n6 VDD1.t3 2.92099
R163 VDD1.n6 VDD1.t5 2.92099
R164 VDD1.n0 VDD1.t1 2.92099
R165 VDD1.n0 VDD1.t6 2.92099
R166 VDD1.n4 VDD1.t9 2.92099
R167 VDD1.n4 VDD1.t8 2.92099
R168 VDD1.n2 VDD1.t0 2.92099
R169 VDD1.n2 VDD1.t4 2.92099
R170 VDD1 VDD1.n7 1.8949
R171 VDD1 VDD1.n1 0.709552
R172 VDD1.n5 VDD1.n3 0.596016
R173 VTAIL.n11 VTAIL.t6 63.2921
R174 VTAIL.n17 VTAIL.t5 63.292
R175 VTAIL.n2 VTAIL.t11 63.292
R176 VTAIL.n16 VTAIL.t12 63.292
R177 VTAIL.n15 VTAIL.n14 60.3717
R178 VTAIL.n13 VTAIL.n12 60.3717
R179 VTAIL.n10 VTAIL.n9 60.3717
R180 VTAIL.n8 VTAIL.n7 60.3717
R181 VTAIL.n19 VTAIL.n18 60.3715
R182 VTAIL.n1 VTAIL.n0 60.3715
R183 VTAIL.n4 VTAIL.n3 60.3715
R184 VTAIL.n6 VTAIL.n5 60.3715
R185 VTAIL.n8 VTAIL.n6 27.1686
R186 VTAIL.n17 VTAIL.n16 24.5652
R187 VTAIL.n18 VTAIL.t2 2.92099
R188 VTAIL.n18 VTAIL.t7 2.92099
R189 VTAIL.n0 VTAIL.t1 2.92099
R190 VTAIL.n0 VTAIL.t3 2.92099
R191 VTAIL.n3 VTAIL.t9 2.92099
R192 VTAIL.n3 VTAIL.t18 2.92099
R193 VTAIL.n5 VTAIL.t15 2.92099
R194 VTAIL.n5 VTAIL.t17 2.92099
R195 VTAIL.n14 VTAIL.t16 2.92099
R196 VTAIL.n14 VTAIL.t10 2.92099
R197 VTAIL.n12 VTAIL.t13 2.92099
R198 VTAIL.n12 VTAIL.t14 2.92099
R199 VTAIL.n9 VTAIL.t4 2.92099
R200 VTAIL.n9 VTAIL.t8 2.92099
R201 VTAIL.n7 VTAIL.t0 2.92099
R202 VTAIL.n7 VTAIL.t19 2.92099
R203 VTAIL.n10 VTAIL.n8 2.60395
R204 VTAIL.n11 VTAIL.n10 2.60395
R205 VTAIL.n15 VTAIL.n13 2.60395
R206 VTAIL.n16 VTAIL.n15 2.60395
R207 VTAIL.n6 VTAIL.n4 2.60395
R208 VTAIL.n4 VTAIL.n2 2.60395
R209 VTAIL.n19 VTAIL.n17 2.60395
R210 VTAIL VTAIL.n1 2.01128
R211 VTAIL.n13 VTAIL.n11 1.77205
R212 VTAIL.n2 VTAIL.n1 1.77205
R213 VTAIL VTAIL.n19 0.593172
R214 B.n444 B.n143 585
R215 B.n443 B.n442 585
R216 B.n441 B.n144 585
R217 B.n440 B.n439 585
R218 B.n438 B.n145 585
R219 B.n437 B.n436 585
R220 B.n435 B.n146 585
R221 B.n434 B.n433 585
R222 B.n432 B.n147 585
R223 B.n431 B.n430 585
R224 B.n429 B.n148 585
R225 B.n428 B.n427 585
R226 B.n426 B.n149 585
R227 B.n425 B.n424 585
R228 B.n423 B.n150 585
R229 B.n422 B.n421 585
R230 B.n420 B.n151 585
R231 B.n419 B.n418 585
R232 B.n417 B.n152 585
R233 B.n416 B.n415 585
R234 B.n414 B.n153 585
R235 B.n413 B.n412 585
R236 B.n411 B.n154 585
R237 B.n410 B.n409 585
R238 B.n408 B.n155 585
R239 B.n407 B.n406 585
R240 B.n405 B.n156 585
R241 B.n404 B.n403 585
R242 B.n402 B.n157 585
R243 B.n401 B.n400 585
R244 B.n399 B.n158 585
R245 B.n398 B.n397 585
R246 B.n396 B.n159 585
R247 B.n395 B.n394 585
R248 B.n393 B.n160 585
R249 B.n392 B.n391 585
R250 B.n390 B.n161 585
R251 B.n389 B.n388 585
R252 B.n387 B.n162 585
R253 B.n386 B.n385 585
R254 B.n381 B.n163 585
R255 B.n380 B.n379 585
R256 B.n378 B.n164 585
R257 B.n377 B.n376 585
R258 B.n375 B.n165 585
R259 B.n374 B.n373 585
R260 B.n372 B.n166 585
R261 B.n371 B.n370 585
R262 B.n369 B.n167 585
R263 B.n367 B.n366 585
R264 B.n365 B.n170 585
R265 B.n364 B.n363 585
R266 B.n362 B.n171 585
R267 B.n361 B.n360 585
R268 B.n359 B.n172 585
R269 B.n358 B.n357 585
R270 B.n356 B.n173 585
R271 B.n355 B.n354 585
R272 B.n353 B.n174 585
R273 B.n352 B.n351 585
R274 B.n350 B.n175 585
R275 B.n349 B.n348 585
R276 B.n347 B.n176 585
R277 B.n346 B.n345 585
R278 B.n344 B.n177 585
R279 B.n343 B.n342 585
R280 B.n341 B.n178 585
R281 B.n340 B.n339 585
R282 B.n338 B.n179 585
R283 B.n337 B.n336 585
R284 B.n335 B.n180 585
R285 B.n334 B.n333 585
R286 B.n332 B.n181 585
R287 B.n331 B.n330 585
R288 B.n329 B.n182 585
R289 B.n328 B.n327 585
R290 B.n326 B.n183 585
R291 B.n325 B.n324 585
R292 B.n323 B.n184 585
R293 B.n322 B.n321 585
R294 B.n320 B.n185 585
R295 B.n319 B.n318 585
R296 B.n317 B.n186 585
R297 B.n316 B.n315 585
R298 B.n314 B.n187 585
R299 B.n313 B.n312 585
R300 B.n311 B.n188 585
R301 B.n310 B.n309 585
R302 B.n446 B.n445 585
R303 B.n447 B.n142 585
R304 B.n449 B.n448 585
R305 B.n450 B.n141 585
R306 B.n452 B.n451 585
R307 B.n453 B.n140 585
R308 B.n455 B.n454 585
R309 B.n456 B.n139 585
R310 B.n458 B.n457 585
R311 B.n459 B.n138 585
R312 B.n461 B.n460 585
R313 B.n462 B.n137 585
R314 B.n464 B.n463 585
R315 B.n465 B.n136 585
R316 B.n467 B.n466 585
R317 B.n468 B.n135 585
R318 B.n470 B.n469 585
R319 B.n471 B.n134 585
R320 B.n473 B.n472 585
R321 B.n474 B.n133 585
R322 B.n476 B.n475 585
R323 B.n477 B.n132 585
R324 B.n479 B.n478 585
R325 B.n480 B.n131 585
R326 B.n482 B.n481 585
R327 B.n483 B.n130 585
R328 B.n485 B.n484 585
R329 B.n486 B.n129 585
R330 B.n488 B.n487 585
R331 B.n489 B.n128 585
R332 B.n491 B.n490 585
R333 B.n492 B.n127 585
R334 B.n494 B.n493 585
R335 B.n495 B.n126 585
R336 B.n497 B.n496 585
R337 B.n498 B.n125 585
R338 B.n500 B.n499 585
R339 B.n501 B.n124 585
R340 B.n503 B.n502 585
R341 B.n504 B.n123 585
R342 B.n506 B.n505 585
R343 B.n507 B.n122 585
R344 B.n509 B.n508 585
R345 B.n510 B.n121 585
R346 B.n512 B.n511 585
R347 B.n513 B.n120 585
R348 B.n515 B.n514 585
R349 B.n516 B.n119 585
R350 B.n518 B.n517 585
R351 B.n519 B.n118 585
R352 B.n521 B.n520 585
R353 B.n522 B.n117 585
R354 B.n524 B.n523 585
R355 B.n525 B.n116 585
R356 B.n527 B.n526 585
R357 B.n528 B.n115 585
R358 B.n530 B.n529 585
R359 B.n531 B.n114 585
R360 B.n533 B.n532 585
R361 B.n534 B.n113 585
R362 B.n536 B.n535 585
R363 B.n537 B.n112 585
R364 B.n539 B.n538 585
R365 B.n540 B.n111 585
R366 B.n542 B.n541 585
R367 B.n543 B.n110 585
R368 B.n545 B.n544 585
R369 B.n546 B.n109 585
R370 B.n548 B.n547 585
R371 B.n549 B.n108 585
R372 B.n551 B.n550 585
R373 B.n552 B.n107 585
R374 B.n554 B.n553 585
R375 B.n555 B.n106 585
R376 B.n557 B.n556 585
R377 B.n558 B.n105 585
R378 B.n560 B.n559 585
R379 B.n561 B.n104 585
R380 B.n563 B.n562 585
R381 B.n564 B.n103 585
R382 B.n566 B.n565 585
R383 B.n567 B.n102 585
R384 B.n569 B.n568 585
R385 B.n570 B.n101 585
R386 B.n572 B.n571 585
R387 B.n573 B.n100 585
R388 B.n575 B.n574 585
R389 B.n576 B.n99 585
R390 B.n578 B.n577 585
R391 B.n579 B.n98 585
R392 B.n581 B.n580 585
R393 B.n582 B.n97 585
R394 B.n584 B.n583 585
R395 B.n585 B.n96 585
R396 B.n587 B.n586 585
R397 B.n588 B.n95 585
R398 B.n590 B.n589 585
R399 B.n591 B.n94 585
R400 B.n593 B.n592 585
R401 B.n594 B.n93 585
R402 B.n596 B.n595 585
R403 B.n597 B.n92 585
R404 B.n599 B.n598 585
R405 B.n600 B.n91 585
R406 B.n602 B.n601 585
R407 B.n603 B.n90 585
R408 B.n605 B.n604 585
R409 B.n606 B.n89 585
R410 B.n608 B.n607 585
R411 B.n609 B.n88 585
R412 B.n611 B.n610 585
R413 B.n612 B.n87 585
R414 B.n614 B.n613 585
R415 B.n615 B.n86 585
R416 B.n617 B.n616 585
R417 B.n618 B.n85 585
R418 B.n620 B.n619 585
R419 B.n621 B.n84 585
R420 B.n623 B.n622 585
R421 B.n624 B.n83 585
R422 B.n626 B.n625 585
R423 B.n627 B.n82 585
R424 B.n629 B.n628 585
R425 B.n630 B.n81 585
R426 B.n764 B.n763 585
R427 B.n762 B.n33 585
R428 B.n761 B.n760 585
R429 B.n759 B.n34 585
R430 B.n758 B.n757 585
R431 B.n756 B.n35 585
R432 B.n755 B.n754 585
R433 B.n753 B.n36 585
R434 B.n752 B.n751 585
R435 B.n750 B.n37 585
R436 B.n749 B.n748 585
R437 B.n747 B.n38 585
R438 B.n746 B.n745 585
R439 B.n744 B.n39 585
R440 B.n743 B.n742 585
R441 B.n741 B.n40 585
R442 B.n740 B.n739 585
R443 B.n738 B.n41 585
R444 B.n737 B.n736 585
R445 B.n735 B.n42 585
R446 B.n734 B.n733 585
R447 B.n732 B.n43 585
R448 B.n731 B.n730 585
R449 B.n729 B.n44 585
R450 B.n728 B.n727 585
R451 B.n726 B.n45 585
R452 B.n725 B.n724 585
R453 B.n723 B.n46 585
R454 B.n722 B.n721 585
R455 B.n720 B.n47 585
R456 B.n719 B.n718 585
R457 B.n717 B.n48 585
R458 B.n716 B.n715 585
R459 B.n714 B.n49 585
R460 B.n713 B.n712 585
R461 B.n711 B.n50 585
R462 B.n710 B.n709 585
R463 B.n708 B.n51 585
R464 B.n707 B.n706 585
R465 B.n705 B.n704 585
R466 B.n703 B.n55 585
R467 B.n702 B.n701 585
R468 B.n700 B.n56 585
R469 B.n699 B.n698 585
R470 B.n697 B.n57 585
R471 B.n696 B.n695 585
R472 B.n694 B.n58 585
R473 B.n693 B.n692 585
R474 B.n691 B.n59 585
R475 B.n689 B.n688 585
R476 B.n687 B.n62 585
R477 B.n686 B.n685 585
R478 B.n684 B.n63 585
R479 B.n683 B.n682 585
R480 B.n681 B.n64 585
R481 B.n680 B.n679 585
R482 B.n678 B.n65 585
R483 B.n677 B.n676 585
R484 B.n675 B.n66 585
R485 B.n674 B.n673 585
R486 B.n672 B.n67 585
R487 B.n671 B.n670 585
R488 B.n669 B.n68 585
R489 B.n668 B.n667 585
R490 B.n666 B.n69 585
R491 B.n665 B.n664 585
R492 B.n663 B.n70 585
R493 B.n662 B.n661 585
R494 B.n660 B.n71 585
R495 B.n659 B.n658 585
R496 B.n657 B.n72 585
R497 B.n656 B.n655 585
R498 B.n654 B.n73 585
R499 B.n653 B.n652 585
R500 B.n651 B.n74 585
R501 B.n650 B.n649 585
R502 B.n648 B.n75 585
R503 B.n647 B.n646 585
R504 B.n645 B.n76 585
R505 B.n644 B.n643 585
R506 B.n642 B.n77 585
R507 B.n641 B.n640 585
R508 B.n639 B.n78 585
R509 B.n638 B.n637 585
R510 B.n636 B.n79 585
R511 B.n635 B.n634 585
R512 B.n633 B.n80 585
R513 B.n632 B.n631 585
R514 B.n765 B.n32 585
R515 B.n767 B.n766 585
R516 B.n768 B.n31 585
R517 B.n770 B.n769 585
R518 B.n771 B.n30 585
R519 B.n773 B.n772 585
R520 B.n774 B.n29 585
R521 B.n776 B.n775 585
R522 B.n777 B.n28 585
R523 B.n779 B.n778 585
R524 B.n780 B.n27 585
R525 B.n782 B.n781 585
R526 B.n783 B.n26 585
R527 B.n785 B.n784 585
R528 B.n786 B.n25 585
R529 B.n788 B.n787 585
R530 B.n789 B.n24 585
R531 B.n791 B.n790 585
R532 B.n792 B.n23 585
R533 B.n794 B.n793 585
R534 B.n795 B.n22 585
R535 B.n797 B.n796 585
R536 B.n798 B.n21 585
R537 B.n800 B.n799 585
R538 B.n801 B.n20 585
R539 B.n803 B.n802 585
R540 B.n804 B.n19 585
R541 B.n806 B.n805 585
R542 B.n807 B.n18 585
R543 B.n809 B.n808 585
R544 B.n810 B.n17 585
R545 B.n812 B.n811 585
R546 B.n813 B.n16 585
R547 B.n815 B.n814 585
R548 B.n816 B.n15 585
R549 B.n818 B.n817 585
R550 B.n819 B.n14 585
R551 B.n821 B.n820 585
R552 B.n822 B.n13 585
R553 B.n824 B.n823 585
R554 B.n825 B.n12 585
R555 B.n827 B.n826 585
R556 B.n828 B.n11 585
R557 B.n830 B.n829 585
R558 B.n831 B.n10 585
R559 B.n833 B.n832 585
R560 B.n834 B.n9 585
R561 B.n836 B.n835 585
R562 B.n837 B.n8 585
R563 B.n839 B.n838 585
R564 B.n840 B.n7 585
R565 B.n842 B.n841 585
R566 B.n843 B.n6 585
R567 B.n845 B.n844 585
R568 B.n846 B.n5 585
R569 B.n848 B.n847 585
R570 B.n849 B.n4 585
R571 B.n851 B.n850 585
R572 B.n852 B.n3 585
R573 B.n854 B.n853 585
R574 B.n855 B.n0 585
R575 B.n2 B.n1 585
R576 B.n220 B.n219 585
R577 B.n221 B.n218 585
R578 B.n223 B.n222 585
R579 B.n224 B.n217 585
R580 B.n226 B.n225 585
R581 B.n227 B.n216 585
R582 B.n229 B.n228 585
R583 B.n230 B.n215 585
R584 B.n232 B.n231 585
R585 B.n233 B.n214 585
R586 B.n235 B.n234 585
R587 B.n236 B.n213 585
R588 B.n238 B.n237 585
R589 B.n239 B.n212 585
R590 B.n241 B.n240 585
R591 B.n242 B.n211 585
R592 B.n244 B.n243 585
R593 B.n245 B.n210 585
R594 B.n247 B.n246 585
R595 B.n248 B.n209 585
R596 B.n250 B.n249 585
R597 B.n251 B.n208 585
R598 B.n253 B.n252 585
R599 B.n254 B.n207 585
R600 B.n256 B.n255 585
R601 B.n257 B.n206 585
R602 B.n259 B.n258 585
R603 B.n260 B.n205 585
R604 B.n262 B.n261 585
R605 B.n263 B.n204 585
R606 B.n265 B.n264 585
R607 B.n266 B.n203 585
R608 B.n268 B.n267 585
R609 B.n269 B.n202 585
R610 B.n271 B.n270 585
R611 B.n272 B.n201 585
R612 B.n274 B.n273 585
R613 B.n275 B.n200 585
R614 B.n277 B.n276 585
R615 B.n278 B.n199 585
R616 B.n280 B.n279 585
R617 B.n281 B.n198 585
R618 B.n283 B.n282 585
R619 B.n284 B.n197 585
R620 B.n286 B.n285 585
R621 B.n287 B.n196 585
R622 B.n289 B.n288 585
R623 B.n290 B.n195 585
R624 B.n292 B.n291 585
R625 B.n293 B.n194 585
R626 B.n295 B.n294 585
R627 B.n296 B.n193 585
R628 B.n298 B.n297 585
R629 B.n299 B.n192 585
R630 B.n301 B.n300 585
R631 B.n302 B.n191 585
R632 B.n304 B.n303 585
R633 B.n305 B.n190 585
R634 B.n307 B.n306 585
R635 B.n308 B.n189 585
R636 B.n310 B.n189 458.866
R637 B.n446 B.n143 458.866
R638 B.n632 B.n81 458.866
R639 B.n765 B.n764 458.866
R640 B.n168 B.t3 307.894
R641 B.n382 B.t0 307.894
R642 B.n60 B.t6 307.894
R643 B.n52 B.t9 307.894
R644 B.n857 B.n856 256.663
R645 B.n856 B.n855 235.042
R646 B.n856 B.n2 235.042
R647 B.n382 B.t1 170.743
R648 B.n60 B.t8 170.743
R649 B.n168 B.t4 170.73
R650 B.n52 B.t11 170.73
R651 B.n311 B.n310 163.367
R652 B.n312 B.n311 163.367
R653 B.n312 B.n187 163.367
R654 B.n316 B.n187 163.367
R655 B.n317 B.n316 163.367
R656 B.n318 B.n317 163.367
R657 B.n318 B.n185 163.367
R658 B.n322 B.n185 163.367
R659 B.n323 B.n322 163.367
R660 B.n324 B.n323 163.367
R661 B.n324 B.n183 163.367
R662 B.n328 B.n183 163.367
R663 B.n329 B.n328 163.367
R664 B.n330 B.n329 163.367
R665 B.n330 B.n181 163.367
R666 B.n334 B.n181 163.367
R667 B.n335 B.n334 163.367
R668 B.n336 B.n335 163.367
R669 B.n336 B.n179 163.367
R670 B.n340 B.n179 163.367
R671 B.n341 B.n340 163.367
R672 B.n342 B.n341 163.367
R673 B.n342 B.n177 163.367
R674 B.n346 B.n177 163.367
R675 B.n347 B.n346 163.367
R676 B.n348 B.n347 163.367
R677 B.n348 B.n175 163.367
R678 B.n352 B.n175 163.367
R679 B.n353 B.n352 163.367
R680 B.n354 B.n353 163.367
R681 B.n354 B.n173 163.367
R682 B.n358 B.n173 163.367
R683 B.n359 B.n358 163.367
R684 B.n360 B.n359 163.367
R685 B.n360 B.n171 163.367
R686 B.n364 B.n171 163.367
R687 B.n365 B.n364 163.367
R688 B.n366 B.n365 163.367
R689 B.n366 B.n167 163.367
R690 B.n371 B.n167 163.367
R691 B.n372 B.n371 163.367
R692 B.n373 B.n372 163.367
R693 B.n373 B.n165 163.367
R694 B.n377 B.n165 163.367
R695 B.n378 B.n377 163.367
R696 B.n379 B.n378 163.367
R697 B.n379 B.n163 163.367
R698 B.n386 B.n163 163.367
R699 B.n387 B.n386 163.367
R700 B.n388 B.n387 163.367
R701 B.n388 B.n161 163.367
R702 B.n392 B.n161 163.367
R703 B.n393 B.n392 163.367
R704 B.n394 B.n393 163.367
R705 B.n394 B.n159 163.367
R706 B.n398 B.n159 163.367
R707 B.n399 B.n398 163.367
R708 B.n400 B.n399 163.367
R709 B.n400 B.n157 163.367
R710 B.n404 B.n157 163.367
R711 B.n405 B.n404 163.367
R712 B.n406 B.n405 163.367
R713 B.n406 B.n155 163.367
R714 B.n410 B.n155 163.367
R715 B.n411 B.n410 163.367
R716 B.n412 B.n411 163.367
R717 B.n412 B.n153 163.367
R718 B.n416 B.n153 163.367
R719 B.n417 B.n416 163.367
R720 B.n418 B.n417 163.367
R721 B.n418 B.n151 163.367
R722 B.n422 B.n151 163.367
R723 B.n423 B.n422 163.367
R724 B.n424 B.n423 163.367
R725 B.n424 B.n149 163.367
R726 B.n428 B.n149 163.367
R727 B.n429 B.n428 163.367
R728 B.n430 B.n429 163.367
R729 B.n430 B.n147 163.367
R730 B.n434 B.n147 163.367
R731 B.n435 B.n434 163.367
R732 B.n436 B.n435 163.367
R733 B.n436 B.n145 163.367
R734 B.n440 B.n145 163.367
R735 B.n441 B.n440 163.367
R736 B.n442 B.n441 163.367
R737 B.n442 B.n143 163.367
R738 B.n628 B.n81 163.367
R739 B.n628 B.n627 163.367
R740 B.n627 B.n626 163.367
R741 B.n626 B.n83 163.367
R742 B.n622 B.n83 163.367
R743 B.n622 B.n621 163.367
R744 B.n621 B.n620 163.367
R745 B.n620 B.n85 163.367
R746 B.n616 B.n85 163.367
R747 B.n616 B.n615 163.367
R748 B.n615 B.n614 163.367
R749 B.n614 B.n87 163.367
R750 B.n610 B.n87 163.367
R751 B.n610 B.n609 163.367
R752 B.n609 B.n608 163.367
R753 B.n608 B.n89 163.367
R754 B.n604 B.n89 163.367
R755 B.n604 B.n603 163.367
R756 B.n603 B.n602 163.367
R757 B.n602 B.n91 163.367
R758 B.n598 B.n91 163.367
R759 B.n598 B.n597 163.367
R760 B.n597 B.n596 163.367
R761 B.n596 B.n93 163.367
R762 B.n592 B.n93 163.367
R763 B.n592 B.n591 163.367
R764 B.n591 B.n590 163.367
R765 B.n590 B.n95 163.367
R766 B.n586 B.n95 163.367
R767 B.n586 B.n585 163.367
R768 B.n585 B.n584 163.367
R769 B.n584 B.n97 163.367
R770 B.n580 B.n97 163.367
R771 B.n580 B.n579 163.367
R772 B.n579 B.n578 163.367
R773 B.n578 B.n99 163.367
R774 B.n574 B.n99 163.367
R775 B.n574 B.n573 163.367
R776 B.n573 B.n572 163.367
R777 B.n572 B.n101 163.367
R778 B.n568 B.n101 163.367
R779 B.n568 B.n567 163.367
R780 B.n567 B.n566 163.367
R781 B.n566 B.n103 163.367
R782 B.n562 B.n103 163.367
R783 B.n562 B.n561 163.367
R784 B.n561 B.n560 163.367
R785 B.n560 B.n105 163.367
R786 B.n556 B.n105 163.367
R787 B.n556 B.n555 163.367
R788 B.n555 B.n554 163.367
R789 B.n554 B.n107 163.367
R790 B.n550 B.n107 163.367
R791 B.n550 B.n549 163.367
R792 B.n549 B.n548 163.367
R793 B.n548 B.n109 163.367
R794 B.n544 B.n109 163.367
R795 B.n544 B.n543 163.367
R796 B.n543 B.n542 163.367
R797 B.n542 B.n111 163.367
R798 B.n538 B.n111 163.367
R799 B.n538 B.n537 163.367
R800 B.n537 B.n536 163.367
R801 B.n536 B.n113 163.367
R802 B.n532 B.n113 163.367
R803 B.n532 B.n531 163.367
R804 B.n531 B.n530 163.367
R805 B.n530 B.n115 163.367
R806 B.n526 B.n115 163.367
R807 B.n526 B.n525 163.367
R808 B.n525 B.n524 163.367
R809 B.n524 B.n117 163.367
R810 B.n520 B.n117 163.367
R811 B.n520 B.n519 163.367
R812 B.n519 B.n518 163.367
R813 B.n518 B.n119 163.367
R814 B.n514 B.n119 163.367
R815 B.n514 B.n513 163.367
R816 B.n513 B.n512 163.367
R817 B.n512 B.n121 163.367
R818 B.n508 B.n121 163.367
R819 B.n508 B.n507 163.367
R820 B.n507 B.n506 163.367
R821 B.n506 B.n123 163.367
R822 B.n502 B.n123 163.367
R823 B.n502 B.n501 163.367
R824 B.n501 B.n500 163.367
R825 B.n500 B.n125 163.367
R826 B.n496 B.n125 163.367
R827 B.n496 B.n495 163.367
R828 B.n495 B.n494 163.367
R829 B.n494 B.n127 163.367
R830 B.n490 B.n127 163.367
R831 B.n490 B.n489 163.367
R832 B.n489 B.n488 163.367
R833 B.n488 B.n129 163.367
R834 B.n484 B.n129 163.367
R835 B.n484 B.n483 163.367
R836 B.n483 B.n482 163.367
R837 B.n482 B.n131 163.367
R838 B.n478 B.n131 163.367
R839 B.n478 B.n477 163.367
R840 B.n477 B.n476 163.367
R841 B.n476 B.n133 163.367
R842 B.n472 B.n133 163.367
R843 B.n472 B.n471 163.367
R844 B.n471 B.n470 163.367
R845 B.n470 B.n135 163.367
R846 B.n466 B.n135 163.367
R847 B.n466 B.n465 163.367
R848 B.n465 B.n464 163.367
R849 B.n464 B.n137 163.367
R850 B.n460 B.n137 163.367
R851 B.n460 B.n459 163.367
R852 B.n459 B.n458 163.367
R853 B.n458 B.n139 163.367
R854 B.n454 B.n139 163.367
R855 B.n454 B.n453 163.367
R856 B.n453 B.n452 163.367
R857 B.n452 B.n141 163.367
R858 B.n448 B.n141 163.367
R859 B.n448 B.n447 163.367
R860 B.n447 B.n446 163.367
R861 B.n764 B.n33 163.367
R862 B.n760 B.n33 163.367
R863 B.n760 B.n759 163.367
R864 B.n759 B.n758 163.367
R865 B.n758 B.n35 163.367
R866 B.n754 B.n35 163.367
R867 B.n754 B.n753 163.367
R868 B.n753 B.n752 163.367
R869 B.n752 B.n37 163.367
R870 B.n748 B.n37 163.367
R871 B.n748 B.n747 163.367
R872 B.n747 B.n746 163.367
R873 B.n746 B.n39 163.367
R874 B.n742 B.n39 163.367
R875 B.n742 B.n741 163.367
R876 B.n741 B.n740 163.367
R877 B.n740 B.n41 163.367
R878 B.n736 B.n41 163.367
R879 B.n736 B.n735 163.367
R880 B.n735 B.n734 163.367
R881 B.n734 B.n43 163.367
R882 B.n730 B.n43 163.367
R883 B.n730 B.n729 163.367
R884 B.n729 B.n728 163.367
R885 B.n728 B.n45 163.367
R886 B.n724 B.n45 163.367
R887 B.n724 B.n723 163.367
R888 B.n723 B.n722 163.367
R889 B.n722 B.n47 163.367
R890 B.n718 B.n47 163.367
R891 B.n718 B.n717 163.367
R892 B.n717 B.n716 163.367
R893 B.n716 B.n49 163.367
R894 B.n712 B.n49 163.367
R895 B.n712 B.n711 163.367
R896 B.n711 B.n710 163.367
R897 B.n710 B.n51 163.367
R898 B.n706 B.n51 163.367
R899 B.n706 B.n705 163.367
R900 B.n705 B.n55 163.367
R901 B.n701 B.n55 163.367
R902 B.n701 B.n700 163.367
R903 B.n700 B.n699 163.367
R904 B.n699 B.n57 163.367
R905 B.n695 B.n57 163.367
R906 B.n695 B.n694 163.367
R907 B.n694 B.n693 163.367
R908 B.n693 B.n59 163.367
R909 B.n688 B.n59 163.367
R910 B.n688 B.n687 163.367
R911 B.n687 B.n686 163.367
R912 B.n686 B.n63 163.367
R913 B.n682 B.n63 163.367
R914 B.n682 B.n681 163.367
R915 B.n681 B.n680 163.367
R916 B.n680 B.n65 163.367
R917 B.n676 B.n65 163.367
R918 B.n676 B.n675 163.367
R919 B.n675 B.n674 163.367
R920 B.n674 B.n67 163.367
R921 B.n670 B.n67 163.367
R922 B.n670 B.n669 163.367
R923 B.n669 B.n668 163.367
R924 B.n668 B.n69 163.367
R925 B.n664 B.n69 163.367
R926 B.n664 B.n663 163.367
R927 B.n663 B.n662 163.367
R928 B.n662 B.n71 163.367
R929 B.n658 B.n71 163.367
R930 B.n658 B.n657 163.367
R931 B.n657 B.n656 163.367
R932 B.n656 B.n73 163.367
R933 B.n652 B.n73 163.367
R934 B.n652 B.n651 163.367
R935 B.n651 B.n650 163.367
R936 B.n650 B.n75 163.367
R937 B.n646 B.n75 163.367
R938 B.n646 B.n645 163.367
R939 B.n645 B.n644 163.367
R940 B.n644 B.n77 163.367
R941 B.n640 B.n77 163.367
R942 B.n640 B.n639 163.367
R943 B.n639 B.n638 163.367
R944 B.n638 B.n79 163.367
R945 B.n634 B.n79 163.367
R946 B.n634 B.n633 163.367
R947 B.n633 B.n632 163.367
R948 B.n766 B.n765 163.367
R949 B.n766 B.n31 163.367
R950 B.n770 B.n31 163.367
R951 B.n771 B.n770 163.367
R952 B.n772 B.n771 163.367
R953 B.n772 B.n29 163.367
R954 B.n776 B.n29 163.367
R955 B.n777 B.n776 163.367
R956 B.n778 B.n777 163.367
R957 B.n778 B.n27 163.367
R958 B.n782 B.n27 163.367
R959 B.n783 B.n782 163.367
R960 B.n784 B.n783 163.367
R961 B.n784 B.n25 163.367
R962 B.n788 B.n25 163.367
R963 B.n789 B.n788 163.367
R964 B.n790 B.n789 163.367
R965 B.n790 B.n23 163.367
R966 B.n794 B.n23 163.367
R967 B.n795 B.n794 163.367
R968 B.n796 B.n795 163.367
R969 B.n796 B.n21 163.367
R970 B.n800 B.n21 163.367
R971 B.n801 B.n800 163.367
R972 B.n802 B.n801 163.367
R973 B.n802 B.n19 163.367
R974 B.n806 B.n19 163.367
R975 B.n807 B.n806 163.367
R976 B.n808 B.n807 163.367
R977 B.n808 B.n17 163.367
R978 B.n812 B.n17 163.367
R979 B.n813 B.n812 163.367
R980 B.n814 B.n813 163.367
R981 B.n814 B.n15 163.367
R982 B.n818 B.n15 163.367
R983 B.n819 B.n818 163.367
R984 B.n820 B.n819 163.367
R985 B.n820 B.n13 163.367
R986 B.n824 B.n13 163.367
R987 B.n825 B.n824 163.367
R988 B.n826 B.n825 163.367
R989 B.n826 B.n11 163.367
R990 B.n830 B.n11 163.367
R991 B.n831 B.n830 163.367
R992 B.n832 B.n831 163.367
R993 B.n832 B.n9 163.367
R994 B.n836 B.n9 163.367
R995 B.n837 B.n836 163.367
R996 B.n838 B.n837 163.367
R997 B.n838 B.n7 163.367
R998 B.n842 B.n7 163.367
R999 B.n843 B.n842 163.367
R1000 B.n844 B.n843 163.367
R1001 B.n844 B.n5 163.367
R1002 B.n848 B.n5 163.367
R1003 B.n849 B.n848 163.367
R1004 B.n850 B.n849 163.367
R1005 B.n850 B.n3 163.367
R1006 B.n854 B.n3 163.367
R1007 B.n855 B.n854 163.367
R1008 B.n220 B.n2 163.367
R1009 B.n221 B.n220 163.367
R1010 B.n222 B.n221 163.367
R1011 B.n222 B.n217 163.367
R1012 B.n226 B.n217 163.367
R1013 B.n227 B.n226 163.367
R1014 B.n228 B.n227 163.367
R1015 B.n228 B.n215 163.367
R1016 B.n232 B.n215 163.367
R1017 B.n233 B.n232 163.367
R1018 B.n234 B.n233 163.367
R1019 B.n234 B.n213 163.367
R1020 B.n238 B.n213 163.367
R1021 B.n239 B.n238 163.367
R1022 B.n240 B.n239 163.367
R1023 B.n240 B.n211 163.367
R1024 B.n244 B.n211 163.367
R1025 B.n245 B.n244 163.367
R1026 B.n246 B.n245 163.367
R1027 B.n246 B.n209 163.367
R1028 B.n250 B.n209 163.367
R1029 B.n251 B.n250 163.367
R1030 B.n252 B.n251 163.367
R1031 B.n252 B.n207 163.367
R1032 B.n256 B.n207 163.367
R1033 B.n257 B.n256 163.367
R1034 B.n258 B.n257 163.367
R1035 B.n258 B.n205 163.367
R1036 B.n262 B.n205 163.367
R1037 B.n263 B.n262 163.367
R1038 B.n264 B.n263 163.367
R1039 B.n264 B.n203 163.367
R1040 B.n268 B.n203 163.367
R1041 B.n269 B.n268 163.367
R1042 B.n270 B.n269 163.367
R1043 B.n270 B.n201 163.367
R1044 B.n274 B.n201 163.367
R1045 B.n275 B.n274 163.367
R1046 B.n276 B.n275 163.367
R1047 B.n276 B.n199 163.367
R1048 B.n280 B.n199 163.367
R1049 B.n281 B.n280 163.367
R1050 B.n282 B.n281 163.367
R1051 B.n282 B.n197 163.367
R1052 B.n286 B.n197 163.367
R1053 B.n287 B.n286 163.367
R1054 B.n288 B.n287 163.367
R1055 B.n288 B.n195 163.367
R1056 B.n292 B.n195 163.367
R1057 B.n293 B.n292 163.367
R1058 B.n294 B.n293 163.367
R1059 B.n294 B.n193 163.367
R1060 B.n298 B.n193 163.367
R1061 B.n299 B.n298 163.367
R1062 B.n300 B.n299 163.367
R1063 B.n300 B.n191 163.367
R1064 B.n304 B.n191 163.367
R1065 B.n305 B.n304 163.367
R1066 B.n306 B.n305 163.367
R1067 B.n306 B.n189 163.367
R1068 B.n383 B.t2 112.174
R1069 B.n61 B.t7 112.174
R1070 B.n169 B.t5 112.16
R1071 B.n53 B.t10 112.16
R1072 B.n368 B.n169 59.5399
R1073 B.n384 B.n383 59.5399
R1074 B.n690 B.n61 59.5399
R1075 B.n54 B.n53 59.5399
R1076 B.n169 B.n168 58.5702
R1077 B.n383 B.n382 58.5702
R1078 B.n61 B.n60 58.5702
R1079 B.n53 B.n52 58.5702
R1080 B.n763 B.n32 29.8151
R1081 B.n631 B.n630 29.8151
R1082 B.n445 B.n444 29.8151
R1083 B.n309 B.n308 29.8151
R1084 B B.n857 18.0485
R1085 B.n767 B.n32 10.6151
R1086 B.n768 B.n767 10.6151
R1087 B.n769 B.n768 10.6151
R1088 B.n769 B.n30 10.6151
R1089 B.n773 B.n30 10.6151
R1090 B.n774 B.n773 10.6151
R1091 B.n775 B.n774 10.6151
R1092 B.n775 B.n28 10.6151
R1093 B.n779 B.n28 10.6151
R1094 B.n780 B.n779 10.6151
R1095 B.n781 B.n780 10.6151
R1096 B.n781 B.n26 10.6151
R1097 B.n785 B.n26 10.6151
R1098 B.n786 B.n785 10.6151
R1099 B.n787 B.n786 10.6151
R1100 B.n787 B.n24 10.6151
R1101 B.n791 B.n24 10.6151
R1102 B.n792 B.n791 10.6151
R1103 B.n793 B.n792 10.6151
R1104 B.n793 B.n22 10.6151
R1105 B.n797 B.n22 10.6151
R1106 B.n798 B.n797 10.6151
R1107 B.n799 B.n798 10.6151
R1108 B.n799 B.n20 10.6151
R1109 B.n803 B.n20 10.6151
R1110 B.n804 B.n803 10.6151
R1111 B.n805 B.n804 10.6151
R1112 B.n805 B.n18 10.6151
R1113 B.n809 B.n18 10.6151
R1114 B.n810 B.n809 10.6151
R1115 B.n811 B.n810 10.6151
R1116 B.n811 B.n16 10.6151
R1117 B.n815 B.n16 10.6151
R1118 B.n816 B.n815 10.6151
R1119 B.n817 B.n816 10.6151
R1120 B.n817 B.n14 10.6151
R1121 B.n821 B.n14 10.6151
R1122 B.n822 B.n821 10.6151
R1123 B.n823 B.n822 10.6151
R1124 B.n823 B.n12 10.6151
R1125 B.n827 B.n12 10.6151
R1126 B.n828 B.n827 10.6151
R1127 B.n829 B.n828 10.6151
R1128 B.n829 B.n10 10.6151
R1129 B.n833 B.n10 10.6151
R1130 B.n834 B.n833 10.6151
R1131 B.n835 B.n834 10.6151
R1132 B.n835 B.n8 10.6151
R1133 B.n839 B.n8 10.6151
R1134 B.n840 B.n839 10.6151
R1135 B.n841 B.n840 10.6151
R1136 B.n841 B.n6 10.6151
R1137 B.n845 B.n6 10.6151
R1138 B.n846 B.n845 10.6151
R1139 B.n847 B.n846 10.6151
R1140 B.n847 B.n4 10.6151
R1141 B.n851 B.n4 10.6151
R1142 B.n852 B.n851 10.6151
R1143 B.n853 B.n852 10.6151
R1144 B.n853 B.n0 10.6151
R1145 B.n763 B.n762 10.6151
R1146 B.n762 B.n761 10.6151
R1147 B.n761 B.n34 10.6151
R1148 B.n757 B.n34 10.6151
R1149 B.n757 B.n756 10.6151
R1150 B.n756 B.n755 10.6151
R1151 B.n755 B.n36 10.6151
R1152 B.n751 B.n36 10.6151
R1153 B.n751 B.n750 10.6151
R1154 B.n750 B.n749 10.6151
R1155 B.n749 B.n38 10.6151
R1156 B.n745 B.n38 10.6151
R1157 B.n745 B.n744 10.6151
R1158 B.n744 B.n743 10.6151
R1159 B.n743 B.n40 10.6151
R1160 B.n739 B.n40 10.6151
R1161 B.n739 B.n738 10.6151
R1162 B.n738 B.n737 10.6151
R1163 B.n737 B.n42 10.6151
R1164 B.n733 B.n42 10.6151
R1165 B.n733 B.n732 10.6151
R1166 B.n732 B.n731 10.6151
R1167 B.n731 B.n44 10.6151
R1168 B.n727 B.n44 10.6151
R1169 B.n727 B.n726 10.6151
R1170 B.n726 B.n725 10.6151
R1171 B.n725 B.n46 10.6151
R1172 B.n721 B.n46 10.6151
R1173 B.n721 B.n720 10.6151
R1174 B.n720 B.n719 10.6151
R1175 B.n719 B.n48 10.6151
R1176 B.n715 B.n48 10.6151
R1177 B.n715 B.n714 10.6151
R1178 B.n714 B.n713 10.6151
R1179 B.n713 B.n50 10.6151
R1180 B.n709 B.n50 10.6151
R1181 B.n709 B.n708 10.6151
R1182 B.n708 B.n707 10.6151
R1183 B.n704 B.n703 10.6151
R1184 B.n703 B.n702 10.6151
R1185 B.n702 B.n56 10.6151
R1186 B.n698 B.n56 10.6151
R1187 B.n698 B.n697 10.6151
R1188 B.n697 B.n696 10.6151
R1189 B.n696 B.n58 10.6151
R1190 B.n692 B.n58 10.6151
R1191 B.n692 B.n691 10.6151
R1192 B.n689 B.n62 10.6151
R1193 B.n685 B.n62 10.6151
R1194 B.n685 B.n684 10.6151
R1195 B.n684 B.n683 10.6151
R1196 B.n683 B.n64 10.6151
R1197 B.n679 B.n64 10.6151
R1198 B.n679 B.n678 10.6151
R1199 B.n678 B.n677 10.6151
R1200 B.n677 B.n66 10.6151
R1201 B.n673 B.n66 10.6151
R1202 B.n673 B.n672 10.6151
R1203 B.n672 B.n671 10.6151
R1204 B.n671 B.n68 10.6151
R1205 B.n667 B.n68 10.6151
R1206 B.n667 B.n666 10.6151
R1207 B.n666 B.n665 10.6151
R1208 B.n665 B.n70 10.6151
R1209 B.n661 B.n70 10.6151
R1210 B.n661 B.n660 10.6151
R1211 B.n660 B.n659 10.6151
R1212 B.n659 B.n72 10.6151
R1213 B.n655 B.n72 10.6151
R1214 B.n655 B.n654 10.6151
R1215 B.n654 B.n653 10.6151
R1216 B.n653 B.n74 10.6151
R1217 B.n649 B.n74 10.6151
R1218 B.n649 B.n648 10.6151
R1219 B.n648 B.n647 10.6151
R1220 B.n647 B.n76 10.6151
R1221 B.n643 B.n76 10.6151
R1222 B.n643 B.n642 10.6151
R1223 B.n642 B.n641 10.6151
R1224 B.n641 B.n78 10.6151
R1225 B.n637 B.n78 10.6151
R1226 B.n637 B.n636 10.6151
R1227 B.n636 B.n635 10.6151
R1228 B.n635 B.n80 10.6151
R1229 B.n631 B.n80 10.6151
R1230 B.n630 B.n629 10.6151
R1231 B.n629 B.n82 10.6151
R1232 B.n625 B.n82 10.6151
R1233 B.n625 B.n624 10.6151
R1234 B.n624 B.n623 10.6151
R1235 B.n623 B.n84 10.6151
R1236 B.n619 B.n84 10.6151
R1237 B.n619 B.n618 10.6151
R1238 B.n618 B.n617 10.6151
R1239 B.n617 B.n86 10.6151
R1240 B.n613 B.n86 10.6151
R1241 B.n613 B.n612 10.6151
R1242 B.n612 B.n611 10.6151
R1243 B.n611 B.n88 10.6151
R1244 B.n607 B.n88 10.6151
R1245 B.n607 B.n606 10.6151
R1246 B.n606 B.n605 10.6151
R1247 B.n605 B.n90 10.6151
R1248 B.n601 B.n90 10.6151
R1249 B.n601 B.n600 10.6151
R1250 B.n600 B.n599 10.6151
R1251 B.n599 B.n92 10.6151
R1252 B.n595 B.n92 10.6151
R1253 B.n595 B.n594 10.6151
R1254 B.n594 B.n593 10.6151
R1255 B.n593 B.n94 10.6151
R1256 B.n589 B.n94 10.6151
R1257 B.n589 B.n588 10.6151
R1258 B.n588 B.n587 10.6151
R1259 B.n587 B.n96 10.6151
R1260 B.n583 B.n96 10.6151
R1261 B.n583 B.n582 10.6151
R1262 B.n582 B.n581 10.6151
R1263 B.n581 B.n98 10.6151
R1264 B.n577 B.n98 10.6151
R1265 B.n577 B.n576 10.6151
R1266 B.n576 B.n575 10.6151
R1267 B.n575 B.n100 10.6151
R1268 B.n571 B.n100 10.6151
R1269 B.n571 B.n570 10.6151
R1270 B.n570 B.n569 10.6151
R1271 B.n569 B.n102 10.6151
R1272 B.n565 B.n102 10.6151
R1273 B.n565 B.n564 10.6151
R1274 B.n564 B.n563 10.6151
R1275 B.n563 B.n104 10.6151
R1276 B.n559 B.n104 10.6151
R1277 B.n559 B.n558 10.6151
R1278 B.n558 B.n557 10.6151
R1279 B.n557 B.n106 10.6151
R1280 B.n553 B.n106 10.6151
R1281 B.n553 B.n552 10.6151
R1282 B.n552 B.n551 10.6151
R1283 B.n551 B.n108 10.6151
R1284 B.n547 B.n108 10.6151
R1285 B.n547 B.n546 10.6151
R1286 B.n546 B.n545 10.6151
R1287 B.n545 B.n110 10.6151
R1288 B.n541 B.n110 10.6151
R1289 B.n541 B.n540 10.6151
R1290 B.n540 B.n539 10.6151
R1291 B.n539 B.n112 10.6151
R1292 B.n535 B.n112 10.6151
R1293 B.n535 B.n534 10.6151
R1294 B.n534 B.n533 10.6151
R1295 B.n533 B.n114 10.6151
R1296 B.n529 B.n114 10.6151
R1297 B.n529 B.n528 10.6151
R1298 B.n528 B.n527 10.6151
R1299 B.n527 B.n116 10.6151
R1300 B.n523 B.n116 10.6151
R1301 B.n523 B.n522 10.6151
R1302 B.n522 B.n521 10.6151
R1303 B.n521 B.n118 10.6151
R1304 B.n517 B.n118 10.6151
R1305 B.n517 B.n516 10.6151
R1306 B.n516 B.n515 10.6151
R1307 B.n515 B.n120 10.6151
R1308 B.n511 B.n120 10.6151
R1309 B.n511 B.n510 10.6151
R1310 B.n510 B.n509 10.6151
R1311 B.n509 B.n122 10.6151
R1312 B.n505 B.n122 10.6151
R1313 B.n505 B.n504 10.6151
R1314 B.n504 B.n503 10.6151
R1315 B.n503 B.n124 10.6151
R1316 B.n499 B.n124 10.6151
R1317 B.n499 B.n498 10.6151
R1318 B.n498 B.n497 10.6151
R1319 B.n497 B.n126 10.6151
R1320 B.n493 B.n126 10.6151
R1321 B.n493 B.n492 10.6151
R1322 B.n492 B.n491 10.6151
R1323 B.n491 B.n128 10.6151
R1324 B.n487 B.n128 10.6151
R1325 B.n487 B.n486 10.6151
R1326 B.n486 B.n485 10.6151
R1327 B.n485 B.n130 10.6151
R1328 B.n481 B.n130 10.6151
R1329 B.n481 B.n480 10.6151
R1330 B.n480 B.n479 10.6151
R1331 B.n479 B.n132 10.6151
R1332 B.n475 B.n132 10.6151
R1333 B.n475 B.n474 10.6151
R1334 B.n474 B.n473 10.6151
R1335 B.n473 B.n134 10.6151
R1336 B.n469 B.n134 10.6151
R1337 B.n469 B.n468 10.6151
R1338 B.n468 B.n467 10.6151
R1339 B.n467 B.n136 10.6151
R1340 B.n463 B.n136 10.6151
R1341 B.n463 B.n462 10.6151
R1342 B.n462 B.n461 10.6151
R1343 B.n461 B.n138 10.6151
R1344 B.n457 B.n138 10.6151
R1345 B.n457 B.n456 10.6151
R1346 B.n456 B.n455 10.6151
R1347 B.n455 B.n140 10.6151
R1348 B.n451 B.n140 10.6151
R1349 B.n451 B.n450 10.6151
R1350 B.n450 B.n449 10.6151
R1351 B.n449 B.n142 10.6151
R1352 B.n445 B.n142 10.6151
R1353 B.n219 B.n1 10.6151
R1354 B.n219 B.n218 10.6151
R1355 B.n223 B.n218 10.6151
R1356 B.n224 B.n223 10.6151
R1357 B.n225 B.n224 10.6151
R1358 B.n225 B.n216 10.6151
R1359 B.n229 B.n216 10.6151
R1360 B.n230 B.n229 10.6151
R1361 B.n231 B.n230 10.6151
R1362 B.n231 B.n214 10.6151
R1363 B.n235 B.n214 10.6151
R1364 B.n236 B.n235 10.6151
R1365 B.n237 B.n236 10.6151
R1366 B.n237 B.n212 10.6151
R1367 B.n241 B.n212 10.6151
R1368 B.n242 B.n241 10.6151
R1369 B.n243 B.n242 10.6151
R1370 B.n243 B.n210 10.6151
R1371 B.n247 B.n210 10.6151
R1372 B.n248 B.n247 10.6151
R1373 B.n249 B.n248 10.6151
R1374 B.n249 B.n208 10.6151
R1375 B.n253 B.n208 10.6151
R1376 B.n254 B.n253 10.6151
R1377 B.n255 B.n254 10.6151
R1378 B.n255 B.n206 10.6151
R1379 B.n259 B.n206 10.6151
R1380 B.n260 B.n259 10.6151
R1381 B.n261 B.n260 10.6151
R1382 B.n261 B.n204 10.6151
R1383 B.n265 B.n204 10.6151
R1384 B.n266 B.n265 10.6151
R1385 B.n267 B.n266 10.6151
R1386 B.n267 B.n202 10.6151
R1387 B.n271 B.n202 10.6151
R1388 B.n272 B.n271 10.6151
R1389 B.n273 B.n272 10.6151
R1390 B.n273 B.n200 10.6151
R1391 B.n277 B.n200 10.6151
R1392 B.n278 B.n277 10.6151
R1393 B.n279 B.n278 10.6151
R1394 B.n279 B.n198 10.6151
R1395 B.n283 B.n198 10.6151
R1396 B.n284 B.n283 10.6151
R1397 B.n285 B.n284 10.6151
R1398 B.n285 B.n196 10.6151
R1399 B.n289 B.n196 10.6151
R1400 B.n290 B.n289 10.6151
R1401 B.n291 B.n290 10.6151
R1402 B.n291 B.n194 10.6151
R1403 B.n295 B.n194 10.6151
R1404 B.n296 B.n295 10.6151
R1405 B.n297 B.n296 10.6151
R1406 B.n297 B.n192 10.6151
R1407 B.n301 B.n192 10.6151
R1408 B.n302 B.n301 10.6151
R1409 B.n303 B.n302 10.6151
R1410 B.n303 B.n190 10.6151
R1411 B.n307 B.n190 10.6151
R1412 B.n308 B.n307 10.6151
R1413 B.n309 B.n188 10.6151
R1414 B.n313 B.n188 10.6151
R1415 B.n314 B.n313 10.6151
R1416 B.n315 B.n314 10.6151
R1417 B.n315 B.n186 10.6151
R1418 B.n319 B.n186 10.6151
R1419 B.n320 B.n319 10.6151
R1420 B.n321 B.n320 10.6151
R1421 B.n321 B.n184 10.6151
R1422 B.n325 B.n184 10.6151
R1423 B.n326 B.n325 10.6151
R1424 B.n327 B.n326 10.6151
R1425 B.n327 B.n182 10.6151
R1426 B.n331 B.n182 10.6151
R1427 B.n332 B.n331 10.6151
R1428 B.n333 B.n332 10.6151
R1429 B.n333 B.n180 10.6151
R1430 B.n337 B.n180 10.6151
R1431 B.n338 B.n337 10.6151
R1432 B.n339 B.n338 10.6151
R1433 B.n339 B.n178 10.6151
R1434 B.n343 B.n178 10.6151
R1435 B.n344 B.n343 10.6151
R1436 B.n345 B.n344 10.6151
R1437 B.n345 B.n176 10.6151
R1438 B.n349 B.n176 10.6151
R1439 B.n350 B.n349 10.6151
R1440 B.n351 B.n350 10.6151
R1441 B.n351 B.n174 10.6151
R1442 B.n355 B.n174 10.6151
R1443 B.n356 B.n355 10.6151
R1444 B.n357 B.n356 10.6151
R1445 B.n357 B.n172 10.6151
R1446 B.n361 B.n172 10.6151
R1447 B.n362 B.n361 10.6151
R1448 B.n363 B.n362 10.6151
R1449 B.n363 B.n170 10.6151
R1450 B.n367 B.n170 10.6151
R1451 B.n370 B.n369 10.6151
R1452 B.n370 B.n166 10.6151
R1453 B.n374 B.n166 10.6151
R1454 B.n375 B.n374 10.6151
R1455 B.n376 B.n375 10.6151
R1456 B.n376 B.n164 10.6151
R1457 B.n380 B.n164 10.6151
R1458 B.n381 B.n380 10.6151
R1459 B.n385 B.n381 10.6151
R1460 B.n389 B.n162 10.6151
R1461 B.n390 B.n389 10.6151
R1462 B.n391 B.n390 10.6151
R1463 B.n391 B.n160 10.6151
R1464 B.n395 B.n160 10.6151
R1465 B.n396 B.n395 10.6151
R1466 B.n397 B.n396 10.6151
R1467 B.n397 B.n158 10.6151
R1468 B.n401 B.n158 10.6151
R1469 B.n402 B.n401 10.6151
R1470 B.n403 B.n402 10.6151
R1471 B.n403 B.n156 10.6151
R1472 B.n407 B.n156 10.6151
R1473 B.n408 B.n407 10.6151
R1474 B.n409 B.n408 10.6151
R1475 B.n409 B.n154 10.6151
R1476 B.n413 B.n154 10.6151
R1477 B.n414 B.n413 10.6151
R1478 B.n415 B.n414 10.6151
R1479 B.n415 B.n152 10.6151
R1480 B.n419 B.n152 10.6151
R1481 B.n420 B.n419 10.6151
R1482 B.n421 B.n420 10.6151
R1483 B.n421 B.n150 10.6151
R1484 B.n425 B.n150 10.6151
R1485 B.n426 B.n425 10.6151
R1486 B.n427 B.n426 10.6151
R1487 B.n427 B.n148 10.6151
R1488 B.n431 B.n148 10.6151
R1489 B.n432 B.n431 10.6151
R1490 B.n433 B.n432 10.6151
R1491 B.n433 B.n146 10.6151
R1492 B.n437 B.n146 10.6151
R1493 B.n438 B.n437 10.6151
R1494 B.n439 B.n438 10.6151
R1495 B.n439 B.n144 10.6151
R1496 B.n443 B.n144 10.6151
R1497 B.n444 B.n443 10.6151
R1498 B.n707 B.n54 9.36635
R1499 B.n690 B.n689 9.36635
R1500 B.n368 B.n367 9.36635
R1501 B.n384 B.n162 9.36635
R1502 B.n857 B.n0 8.11757
R1503 B.n857 B.n1 8.11757
R1504 B.n704 B.n54 1.24928
R1505 B.n691 B.n690 1.24928
R1506 B.n369 B.n368 1.24928
R1507 B.n385 B.n384 1.24928
R1508 VN.n83 VN.n43 161.3
R1509 VN.n82 VN.n81 161.3
R1510 VN.n80 VN.n44 161.3
R1511 VN.n79 VN.n78 161.3
R1512 VN.n77 VN.n45 161.3
R1513 VN.n76 VN.n75 161.3
R1514 VN.n74 VN.n73 161.3
R1515 VN.n72 VN.n47 161.3
R1516 VN.n71 VN.n70 161.3
R1517 VN.n69 VN.n48 161.3
R1518 VN.n68 VN.n67 161.3
R1519 VN.n66 VN.n49 161.3
R1520 VN.n65 VN.n64 161.3
R1521 VN.n63 VN.n50 161.3
R1522 VN.n62 VN.n61 161.3
R1523 VN.n60 VN.n51 161.3
R1524 VN.n59 VN.n58 161.3
R1525 VN.n57 VN.n52 161.3
R1526 VN.n56 VN.n55 161.3
R1527 VN.n40 VN.n0 161.3
R1528 VN.n39 VN.n38 161.3
R1529 VN.n37 VN.n1 161.3
R1530 VN.n36 VN.n35 161.3
R1531 VN.n34 VN.n2 161.3
R1532 VN.n33 VN.n32 161.3
R1533 VN.n31 VN.n30 161.3
R1534 VN.n29 VN.n4 161.3
R1535 VN.n28 VN.n27 161.3
R1536 VN.n26 VN.n5 161.3
R1537 VN.n25 VN.n24 161.3
R1538 VN.n23 VN.n6 161.3
R1539 VN.n22 VN.n21 161.3
R1540 VN.n20 VN.n7 161.3
R1541 VN.n19 VN.n18 161.3
R1542 VN.n17 VN.n8 161.3
R1543 VN.n16 VN.n15 161.3
R1544 VN.n14 VN.n9 161.3
R1545 VN.n13 VN.n12 161.3
R1546 VN.n10 VN.t5 130.427
R1547 VN.n53 VN.t3 130.427
R1548 VN.n42 VN.n41 108.799
R1549 VN.n85 VN.n84 108.799
R1550 VN.n22 VN.t7 99.7154
R1551 VN.n11 VN.t4 99.7154
R1552 VN.n3 VN.t6 99.7154
R1553 VN.n41 VN.t8 99.7154
R1554 VN.n65 VN.t1 99.7154
R1555 VN.n54 VN.t2 99.7154
R1556 VN.n46 VN.t0 99.7154
R1557 VN.n84 VN.t9 99.7154
R1558 VN.n11 VN.n10 72.37
R1559 VN.n54 VN.n53 72.37
R1560 VN VN.n85 53.1421
R1561 VN.n35 VN.n1 43.4072
R1562 VN.n78 VN.n44 43.4072
R1563 VN.n17 VN.n16 41.4647
R1564 VN.n28 VN.n5 41.4647
R1565 VN.n60 VN.n59 41.4647
R1566 VN.n71 VN.n48 41.4647
R1567 VN.n18 VN.n17 39.5221
R1568 VN.n24 VN.n5 39.5221
R1569 VN.n61 VN.n60 39.5221
R1570 VN.n67 VN.n48 39.5221
R1571 VN.n35 VN.n34 37.5796
R1572 VN.n78 VN.n77 37.5796
R1573 VN.n12 VN.n9 24.4675
R1574 VN.n16 VN.n9 24.4675
R1575 VN.n18 VN.n7 24.4675
R1576 VN.n22 VN.n7 24.4675
R1577 VN.n23 VN.n22 24.4675
R1578 VN.n24 VN.n23 24.4675
R1579 VN.n29 VN.n28 24.4675
R1580 VN.n30 VN.n29 24.4675
R1581 VN.n34 VN.n33 24.4675
R1582 VN.n39 VN.n1 24.4675
R1583 VN.n40 VN.n39 24.4675
R1584 VN.n59 VN.n52 24.4675
R1585 VN.n55 VN.n52 24.4675
R1586 VN.n67 VN.n66 24.4675
R1587 VN.n66 VN.n65 24.4675
R1588 VN.n65 VN.n50 24.4675
R1589 VN.n61 VN.n50 24.4675
R1590 VN.n77 VN.n76 24.4675
R1591 VN.n73 VN.n72 24.4675
R1592 VN.n72 VN.n71 24.4675
R1593 VN.n83 VN.n82 24.4675
R1594 VN.n82 VN.n44 24.4675
R1595 VN.n33 VN.n3 23.4888
R1596 VN.n76 VN.n46 23.4888
R1597 VN.n56 VN.n53 7.37486
R1598 VN.n13 VN.n10 7.37486
R1599 VN.n41 VN.n40 1.95786
R1600 VN.n84 VN.n83 1.95786
R1601 VN.n12 VN.n11 0.97918
R1602 VN.n30 VN.n3 0.97918
R1603 VN.n55 VN.n54 0.97918
R1604 VN.n73 VN.n46 0.97918
R1605 VN.n85 VN.n43 0.278367
R1606 VN.n42 VN.n0 0.278367
R1607 VN.n81 VN.n43 0.189894
R1608 VN.n81 VN.n80 0.189894
R1609 VN.n80 VN.n79 0.189894
R1610 VN.n79 VN.n45 0.189894
R1611 VN.n75 VN.n45 0.189894
R1612 VN.n75 VN.n74 0.189894
R1613 VN.n74 VN.n47 0.189894
R1614 VN.n70 VN.n47 0.189894
R1615 VN.n70 VN.n69 0.189894
R1616 VN.n69 VN.n68 0.189894
R1617 VN.n68 VN.n49 0.189894
R1618 VN.n64 VN.n49 0.189894
R1619 VN.n64 VN.n63 0.189894
R1620 VN.n63 VN.n62 0.189894
R1621 VN.n62 VN.n51 0.189894
R1622 VN.n58 VN.n51 0.189894
R1623 VN.n58 VN.n57 0.189894
R1624 VN.n57 VN.n56 0.189894
R1625 VN.n14 VN.n13 0.189894
R1626 VN.n15 VN.n14 0.189894
R1627 VN.n15 VN.n8 0.189894
R1628 VN.n19 VN.n8 0.189894
R1629 VN.n20 VN.n19 0.189894
R1630 VN.n21 VN.n20 0.189894
R1631 VN.n21 VN.n6 0.189894
R1632 VN.n25 VN.n6 0.189894
R1633 VN.n26 VN.n25 0.189894
R1634 VN.n27 VN.n26 0.189894
R1635 VN.n27 VN.n4 0.189894
R1636 VN.n31 VN.n4 0.189894
R1637 VN.n32 VN.n31 0.189894
R1638 VN.n32 VN.n2 0.189894
R1639 VN.n36 VN.n2 0.189894
R1640 VN.n37 VN.n36 0.189894
R1641 VN.n38 VN.n37 0.189894
R1642 VN.n38 VN.n0 0.189894
R1643 VN VN.n42 0.153454
R1644 VDD2.n1 VDD2.t4 82.5743
R1645 VDD2.n4 VDD2.t0 79.9709
R1646 VDD2.n3 VDD2.n2 78.9475
R1647 VDD2 VDD2.n7 78.9447
R1648 VDD2.n6 VDD2.n5 77.0505
R1649 VDD2.n1 VDD2.n0 77.0503
R1650 VDD2.n4 VDD2.n3 45.6765
R1651 VDD2.n7 VDD2.t7 2.92099
R1652 VDD2.n7 VDD2.t6 2.92099
R1653 VDD2.n5 VDD2.t9 2.92099
R1654 VDD2.n5 VDD2.t8 2.92099
R1655 VDD2.n2 VDD2.t3 2.92099
R1656 VDD2.n2 VDD2.t1 2.92099
R1657 VDD2.n0 VDD2.t5 2.92099
R1658 VDD2.n0 VDD2.t2 2.92099
R1659 VDD2.n6 VDD2.n4 2.60395
R1660 VDD2 VDD2.n6 0.709552
R1661 VDD2.n3 VDD2.n1 0.596016
C0 w_n4594_n3194# B 10.4545f
C1 VP B 2.30274f
C2 VTAIL w_n4594_n3194# 3.09053f
C3 VDD1 B 2.44669f
C4 VTAIL VP 10.7382f
C5 VDD2 B 2.56811f
C6 VTAIL VDD1 10.019401f
C7 VTAIL VDD2 10.0712f
C8 w_n4594_n3194# VP 10.4509f
C9 VDD1 w_n4594_n3194# 2.75689f
C10 VN B 1.29601f
C11 VDD1 VP 10.4443f
C12 w_n4594_n3194# VDD2 2.90511f
C13 VP VDD2 0.594622f
C14 VTAIL VN 10.723901f
C15 VDD1 VDD2 2.2303f
C16 VTAIL B 3.57204f
C17 VN w_n4594_n3194# 9.852469f
C18 VN VP 8.372869f
C19 VDD1 VN 0.153196f
C20 VN VDD2 10.0066f
C21 VDD2 VSUBS 2.189784f
C22 VDD1 VSUBS 1.974162f
C23 VTAIL VSUBS 1.289329f
C24 VN VSUBS 7.789751f
C25 VP VSUBS 4.309474f
C26 B VSUBS 5.406625f
C27 w_n4594_n3194# VSUBS 0.180875p
C28 VDD2.t4 VSUBS 2.74477f
C29 VDD2.t5 VSUBS 0.268682f
C30 VDD2.t2 VSUBS 0.268682f
C31 VDD2.n0 VSUBS 2.07576f
C32 VDD2.n1 VSUBS 1.76545f
C33 VDD2.t3 VSUBS 0.268682f
C34 VDD2.t1 VSUBS 0.268682f
C35 VDD2.n2 VSUBS 2.10013f
C36 VDD2.n3 VSUBS 3.84544f
C37 VDD2.t0 VSUBS 2.71578f
C38 VDD2.n4 VSUBS 4.09727f
C39 VDD2.t9 VSUBS 0.268682f
C40 VDD2.t8 VSUBS 0.268682f
C41 VDD2.n5 VSUBS 2.07576f
C42 VDD2.n6 VSUBS 0.884578f
C43 VDD2.t7 VSUBS 0.268682f
C44 VDD2.t6 VSUBS 0.268682f
C45 VDD2.n7 VSUBS 2.10008f
C46 VN.n0 VSUBS 0.037447f
C47 VN.t8 VSUBS 2.31181f
C48 VN.n1 VSUBS 0.055443f
C49 VN.n2 VSUBS 0.028403f
C50 VN.t6 VSUBS 2.31181f
C51 VN.n3 VSUBS 0.820531f
C52 VN.n4 VSUBS 0.028403f
C53 VN.n5 VSUBS 0.022998f
C54 VN.n6 VSUBS 0.028403f
C55 VN.t7 VSUBS 2.31181f
C56 VN.n7 VSUBS 0.052937f
C57 VN.n8 VSUBS 0.028403f
C58 VN.n9 VSUBS 0.052937f
C59 VN.t5 VSUBS 2.54651f
C60 VN.n10 VSUBS 0.883097f
C61 VN.t4 VSUBS 2.31181f
C62 VN.n11 VSUBS 0.894524f
C63 VN.n12 VSUBS 0.027847f
C64 VN.n13 VSUBS 0.276585f
C65 VN.n14 VSUBS 0.028403f
C66 VN.n15 VSUBS 0.028403f
C67 VN.n16 VSUBS 0.056149f
C68 VN.n17 VSUBS 0.022998f
C69 VN.n18 VSUBS 0.056718f
C70 VN.n19 VSUBS 0.028403f
C71 VN.n20 VSUBS 0.028403f
C72 VN.n21 VSUBS 0.028403f
C73 VN.n22 VSUBS 0.847332f
C74 VN.n23 VSUBS 0.052937f
C75 VN.n24 VSUBS 0.056718f
C76 VN.n25 VSUBS 0.028403f
C77 VN.n26 VSUBS 0.028403f
C78 VN.n27 VSUBS 0.028403f
C79 VN.n28 VSUBS 0.056149f
C80 VN.n29 VSUBS 0.052937f
C81 VN.n30 VSUBS 0.027847f
C82 VN.n31 VSUBS 0.028403f
C83 VN.n32 VSUBS 0.028403f
C84 VN.n33 VSUBS 0.051891f
C85 VN.n34 VSUBS 0.057129f
C86 VN.n35 VSUBS 0.023292f
C87 VN.n36 VSUBS 0.028403f
C88 VN.n37 VSUBS 0.028403f
C89 VN.n38 VSUBS 0.028403f
C90 VN.n39 VSUBS 0.052937f
C91 VN.n40 VSUBS 0.028892f
C92 VN.n41 VSUBS 0.907031f
C93 VN.n42 VSUBS 0.052236f
C94 VN.n43 VSUBS 0.037447f
C95 VN.t9 VSUBS 2.31181f
C96 VN.n44 VSUBS 0.055443f
C97 VN.n45 VSUBS 0.028403f
C98 VN.t0 VSUBS 2.31181f
C99 VN.n46 VSUBS 0.820531f
C100 VN.n47 VSUBS 0.028403f
C101 VN.n48 VSUBS 0.022998f
C102 VN.n49 VSUBS 0.028403f
C103 VN.t1 VSUBS 2.31181f
C104 VN.n50 VSUBS 0.052937f
C105 VN.n51 VSUBS 0.028403f
C106 VN.n52 VSUBS 0.052937f
C107 VN.t3 VSUBS 2.54651f
C108 VN.n53 VSUBS 0.883097f
C109 VN.t2 VSUBS 2.31181f
C110 VN.n54 VSUBS 0.894524f
C111 VN.n55 VSUBS 0.027847f
C112 VN.n56 VSUBS 0.276585f
C113 VN.n57 VSUBS 0.028403f
C114 VN.n58 VSUBS 0.028403f
C115 VN.n59 VSUBS 0.056149f
C116 VN.n60 VSUBS 0.022998f
C117 VN.n61 VSUBS 0.056718f
C118 VN.n62 VSUBS 0.028403f
C119 VN.n63 VSUBS 0.028403f
C120 VN.n64 VSUBS 0.028403f
C121 VN.n65 VSUBS 0.847332f
C122 VN.n66 VSUBS 0.052937f
C123 VN.n67 VSUBS 0.056718f
C124 VN.n68 VSUBS 0.028403f
C125 VN.n69 VSUBS 0.028403f
C126 VN.n70 VSUBS 0.028403f
C127 VN.n71 VSUBS 0.056149f
C128 VN.n72 VSUBS 0.052937f
C129 VN.n73 VSUBS 0.027847f
C130 VN.n74 VSUBS 0.028403f
C131 VN.n75 VSUBS 0.028403f
C132 VN.n76 VSUBS 0.051891f
C133 VN.n77 VSUBS 0.057129f
C134 VN.n78 VSUBS 0.023292f
C135 VN.n79 VSUBS 0.028403f
C136 VN.n80 VSUBS 0.028403f
C137 VN.n81 VSUBS 0.028403f
C138 VN.n82 VSUBS 0.052937f
C139 VN.n83 VSUBS 0.028892f
C140 VN.n84 VSUBS 0.907031f
C141 VN.n85 VSUBS 1.7336f
C142 B.n0 VSUBS 0.008427f
C143 B.n1 VSUBS 0.008427f
C144 B.n2 VSUBS 0.012463f
C145 B.n3 VSUBS 0.009551f
C146 B.n4 VSUBS 0.009551f
C147 B.n5 VSUBS 0.009551f
C148 B.n6 VSUBS 0.009551f
C149 B.n7 VSUBS 0.009551f
C150 B.n8 VSUBS 0.009551f
C151 B.n9 VSUBS 0.009551f
C152 B.n10 VSUBS 0.009551f
C153 B.n11 VSUBS 0.009551f
C154 B.n12 VSUBS 0.009551f
C155 B.n13 VSUBS 0.009551f
C156 B.n14 VSUBS 0.009551f
C157 B.n15 VSUBS 0.009551f
C158 B.n16 VSUBS 0.009551f
C159 B.n17 VSUBS 0.009551f
C160 B.n18 VSUBS 0.009551f
C161 B.n19 VSUBS 0.009551f
C162 B.n20 VSUBS 0.009551f
C163 B.n21 VSUBS 0.009551f
C164 B.n22 VSUBS 0.009551f
C165 B.n23 VSUBS 0.009551f
C166 B.n24 VSUBS 0.009551f
C167 B.n25 VSUBS 0.009551f
C168 B.n26 VSUBS 0.009551f
C169 B.n27 VSUBS 0.009551f
C170 B.n28 VSUBS 0.009551f
C171 B.n29 VSUBS 0.009551f
C172 B.n30 VSUBS 0.009551f
C173 B.n31 VSUBS 0.009551f
C174 B.n32 VSUBS 0.02042f
C175 B.n33 VSUBS 0.009551f
C176 B.n34 VSUBS 0.009551f
C177 B.n35 VSUBS 0.009551f
C178 B.n36 VSUBS 0.009551f
C179 B.n37 VSUBS 0.009551f
C180 B.n38 VSUBS 0.009551f
C181 B.n39 VSUBS 0.009551f
C182 B.n40 VSUBS 0.009551f
C183 B.n41 VSUBS 0.009551f
C184 B.n42 VSUBS 0.009551f
C185 B.n43 VSUBS 0.009551f
C186 B.n44 VSUBS 0.009551f
C187 B.n45 VSUBS 0.009551f
C188 B.n46 VSUBS 0.009551f
C189 B.n47 VSUBS 0.009551f
C190 B.n48 VSUBS 0.009551f
C191 B.n49 VSUBS 0.009551f
C192 B.n50 VSUBS 0.009551f
C193 B.n51 VSUBS 0.009551f
C194 B.t10 VSUBS 0.490743f
C195 B.t11 VSUBS 0.519819f
C196 B.t9 VSUBS 1.87339f
C197 B.n52 VSUBS 0.275185f
C198 B.n53 VSUBS 0.098377f
C199 B.n54 VSUBS 0.022128f
C200 B.n55 VSUBS 0.009551f
C201 B.n56 VSUBS 0.009551f
C202 B.n57 VSUBS 0.009551f
C203 B.n58 VSUBS 0.009551f
C204 B.n59 VSUBS 0.009551f
C205 B.t7 VSUBS 0.490735f
C206 B.t8 VSUBS 0.519811f
C207 B.t6 VSUBS 1.87339f
C208 B.n60 VSUBS 0.275193f
C209 B.n61 VSUBS 0.098385f
C210 B.n62 VSUBS 0.009551f
C211 B.n63 VSUBS 0.009551f
C212 B.n64 VSUBS 0.009551f
C213 B.n65 VSUBS 0.009551f
C214 B.n66 VSUBS 0.009551f
C215 B.n67 VSUBS 0.009551f
C216 B.n68 VSUBS 0.009551f
C217 B.n69 VSUBS 0.009551f
C218 B.n70 VSUBS 0.009551f
C219 B.n71 VSUBS 0.009551f
C220 B.n72 VSUBS 0.009551f
C221 B.n73 VSUBS 0.009551f
C222 B.n74 VSUBS 0.009551f
C223 B.n75 VSUBS 0.009551f
C224 B.n76 VSUBS 0.009551f
C225 B.n77 VSUBS 0.009551f
C226 B.n78 VSUBS 0.009551f
C227 B.n79 VSUBS 0.009551f
C228 B.n80 VSUBS 0.009551f
C229 B.n81 VSUBS 0.02042f
C230 B.n82 VSUBS 0.009551f
C231 B.n83 VSUBS 0.009551f
C232 B.n84 VSUBS 0.009551f
C233 B.n85 VSUBS 0.009551f
C234 B.n86 VSUBS 0.009551f
C235 B.n87 VSUBS 0.009551f
C236 B.n88 VSUBS 0.009551f
C237 B.n89 VSUBS 0.009551f
C238 B.n90 VSUBS 0.009551f
C239 B.n91 VSUBS 0.009551f
C240 B.n92 VSUBS 0.009551f
C241 B.n93 VSUBS 0.009551f
C242 B.n94 VSUBS 0.009551f
C243 B.n95 VSUBS 0.009551f
C244 B.n96 VSUBS 0.009551f
C245 B.n97 VSUBS 0.009551f
C246 B.n98 VSUBS 0.009551f
C247 B.n99 VSUBS 0.009551f
C248 B.n100 VSUBS 0.009551f
C249 B.n101 VSUBS 0.009551f
C250 B.n102 VSUBS 0.009551f
C251 B.n103 VSUBS 0.009551f
C252 B.n104 VSUBS 0.009551f
C253 B.n105 VSUBS 0.009551f
C254 B.n106 VSUBS 0.009551f
C255 B.n107 VSUBS 0.009551f
C256 B.n108 VSUBS 0.009551f
C257 B.n109 VSUBS 0.009551f
C258 B.n110 VSUBS 0.009551f
C259 B.n111 VSUBS 0.009551f
C260 B.n112 VSUBS 0.009551f
C261 B.n113 VSUBS 0.009551f
C262 B.n114 VSUBS 0.009551f
C263 B.n115 VSUBS 0.009551f
C264 B.n116 VSUBS 0.009551f
C265 B.n117 VSUBS 0.009551f
C266 B.n118 VSUBS 0.009551f
C267 B.n119 VSUBS 0.009551f
C268 B.n120 VSUBS 0.009551f
C269 B.n121 VSUBS 0.009551f
C270 B.n122 VSUBS 0.009551f
C271 B.n123 VSUBS 0.009551f
C272 B.n124 VSUBS 0.009551f
C273 B.n125 VSUBS 0.009551f
C274 B.n126 VSUBS 0.009551f
C275 B.n127 VSUBS 0.009551f
C276 B.n128 VSUBS 0.009551f
C277 B.n129 VSUBS 0.009551f
C278 B.n130 VSUBS 0.009551f
C279 B.n131 VSUBS 0.009551f
C280 B.n132 VSUBS 0.009551f
C281 B.n133 VSUBS 0.009551f
C282 B.n134 VSUBS 0.009551f
C283 B.n135 VSUBS 0.009551f
C284 B.n136 VSUBS 0.009551f
C285 B.n137 VSUBS 0.009551f
C286 B.n138 VSUBS 0.009551f
C287 B.n139 VSUBS 0.009551f
C288 B.n140 VSUBS 0.009551f
C289 B.n141 VSUBS 0.009551f
C290 B.n142 VSUBS 0.009551f
C291 B.n143 VSUBS 0.021716f
C292 B.n144 VSUBS 0.009551f
C293 B.n145 VSUBS 0.009551f
C294 B.n146 VSUBS 0.009551f
C295 B.n147 VSUBS 0.009551f
C296 B.n148 VSUBS 0.009551f
C297 B.n149 VSUBS 0.009551f
C298 B.n150 VSUBS 0.009551f
C299 B.n151 VSUBS 0.009551f
C300 B.n152 VSUBS 0.009551f
C301 B.n153 VSUBS 0.009551f
C302 B.n154 VSUBS 0.009551f
C303 B.n155 VSUBS 0.009551f
C304 B.n156 VSUBS 0.009551f
C305 B.n157 VSUBS 0.009551f
C306 B.n158 VSUBS 0.009551f
C307 B.n159 VSUBS 0.009551f
C308 B.n160 VSUBS 0.009551f
C309 B.n161 VSUBS 0.009551f
C310 B.n162 VSUBS 0.008989f
C311 B.n163 VSUBS 0.009551f
C312 B.n164 VSUBS 0.009551f
C313 B.n165 VSUBS 0.009551f
C314 B.n166 VSUBS 0.009551f
C315 B.n167 VSUBS 0.009551f
C316 B.t5 VSUBS 0.490743f
C317 B.t4 VSUBS 0.519819f
C318 B.t3 VSUBS 1.87339f
C319 B.n168 VSUBS 0.275185f
C320 B.n169 VSUBS 0.098377f
C321 B.n170 VSUBS 0.009551f
C322 B.n171 VSUBS 0.009551f
C323 B.n172 VSUBS 0.009551f
C324 B.n173 VSUBS 0.009551f
C325 B.n174 VSUBS 0.009551f
C326 B.n175 VSUBS 0.009551f
C327 B.n176 VSUBS 0.009551f
C328 B.n177 VSUBS 0.009551f
C329 B.n178 VSUBS 0.009551f
C330 B.n179 VSUBS 0.009551f
C331 B.n180 VSUBS 0.009551f
C332 B.n181 VSUBS 0.009551f
C333 B.n182 VSUBS 0.009551f
C334 B.n183 VSUBS 0.009551f
C335 B.n184 VSUBS 0.009551f
C336 B.n185 VSUBS 0.009551f
C337 B.n186 VSUBS 0.009551f
C338 B.n187 VSUBS 0.009551f
C339 B.n188 VSUBS 0.009551f
C340 B.n189 VSUBS 0.02042f
C341 B.n190 VSUBS 0.009551f
C342 B.n191 VSUBS 0.009551f
C343 B.n192 VSUBS 0.009551f
C344 B.n193 VSUBS 0.009551f
C345 B.n194 VSUBS 0.009551f
C346 B.n195 VSUBS 0.009551f
C347 B.n196 VSUBS 0.009551f
C348 B.n197 VSUBS 0.009551f
C349 B.n198 VSUBS 0.009551f
C350 B.n199 VSUBS 0.009551f
C351 B.n200 VSUBS 0.009551f
C352 B.n201 VSUBS 0.009551f
C353 B.n202 VSUBS 0.009551f
C354 B.n203 VSUBS 0.009551f
C355 B.n204 VSUBS 0.009551f
C356 B.n205 VSUBS 0.009551f
C357 B.n206 VSUBS 0.009551f
C358 B.n207 VSUBS 0.009551f
C359 B.n208 VSUBS 0.009551f
C360 B.n209 VSUBS 0.009551f
C361 B.n210 VSUBS 0.009551f
C362 B.n211 VSUBS 0.009551f
C363 B.n212 VSUBS 0.009551f
C364 B.n213 VSUBS 0.009551f
C365 B.n214 VSUBS 0.009551f
C366 B.n215 VSUBS 0.009551f
C367 B.n216 VSUBS 0.009551f
C368 B.n217 VSUBS 0.009551f
C369 B.n218 VSUBS 0.009551f
C370 B.n219 VSUBS 0.009551f
C371 B.n220 VSUBS 0.009551f
C372 B.n221 VSUBS 0.009551f
C373 B.n222 VSUBS 0.009551f
C374 B.n223 VSUBS 0.009551f
C375 B.n224 VSUBS 0.009551f
C376 B.n225 VSUBS 0.009551f
C377 B.n226 VSUBS 0.009551f
C378 B.n227 VSUBS 0.009551f
C379 B.n228 VSUBS 0.009551f
C380 B.n229 VSUBS 0.009551f
C381 B.n230 VSUBS 0.009551f
C382 B.n231 VSUBS 0.009551f
C383 B.n232 VSUBS 0.009551f
C384 B.n233 VSUBS 0.009551f
C385 B.n234 VSUBS 0.009551f
C386 B.n235 VSUBS 0.009551f
C387 B.n236 VSUBS 0.009551f
C388 B.n237 VSUBS 0.009551f
C389 B.n238 VSUBS 0.009551f
C390 B.n239 VSUBS 0.009551f
C391 B.n240 VSUBS 0.009551f
C392 B.n241 VSUBS 0.009551f
C393 B.n242 VSUBS 0.009551f
C394 B.n243 VSUBS 0.009551f
C395 B.n244 VSUBS 0.009551f
C396 B.n245 VSUBS 0.009551f
C397 B.n246 VSUBS 0.009551f
C398 B.n247 VSUBS 0.009551f
C399 B.n248 VSUBS 0.009551f
C400 B.n249 VSUBS 0.009551f
C401 B.n250 VSUBS 0.009551f
C402 B.n251 VSUBS 0.009551f
C403 B.n252 VSUBS 0.009551f
C404 B.n253 VSUBS 0.009551f
C405 B.n254 VSUBS 0.009551f
C406 B.n255 VSUBS 0.009551f
C407 B.n256 VSUBS 0.009551f
C408 B.n257 VSUBS 0.009551f
C409 B.n258 VSUBS 0.009551f
C410 B.n259 VSUBS 0.009551f
C411 B.n260 VSUBS 0.009551f
C412 B.n261 VSUBS 0.009551f
C413 B.n262 VSUBS 0.009551f
C414 B.n263 VSUBS 0.009551f
C415 B.n264 VSUBS 0.009551f
C416 B.n265 VSUBS 0.009551f
C417 B.n266 VSUBS 0.009551f
C418 B.n267 VSUBS 0.009551f
C419 B.n268 VSUBS 0.009551f
C420 B.n269 VSUBS 0.009551f
C421 B.n270 VSUBS 0.009551f
C422 B.n271 VSUBS 0.009551f
C423 B.n272 VSUBS 0.009551f
C424 B.n273 VSUBS 0.009551f
C425 B.n274 VSUBS 0.009551f
C426 B.n275 VSUBS 0.009551f
C427 B.n276 VSUBS 0.009551f
C428 B.n277 VSUBS 0.009551f
C429 B.n278 VSUBS 0.009551f
C430 B.n279 VSUBS 0.009551f
C431 B.n280 VSUBS 0.009551f
C432 B.n281 VSUBS 0.009551f
C433 B.n282 VSUBS 0.009551f
C434 B.n283 VSUBS 0.009551f
C435 B.n284 VSUBS 0.009551f
C436 B.n285 VSUBS 0.009551f
C437 B.n286 VSUBS 0.009551f
C438 B.n287 VSUBS 0.009551f
C439 B.n288 VSUBS 0.009551f
C440 B.n289 VSUBS 0.009551f
C441 B.n290 VSUBS 0.009551f
C442 B.n291 VSUBS 0.009551f
C443 B.n292 VSUBS 0.009551f
C444 B.n293 VSUBS 0.009551f
C445 B.n294 VSUBS 0.009551f
C446 B.n295 VSUBS 0.009551f
C447 B.n296 VSUBS 0.009551f
C448 B.n297 VSUBS 0.009551f
C449 B.n298 VSUBS 0.009551f
C450 B.n299 VSUBS 0.009551f
C451 B.n300 VSUBS 0.009551f
C452 B.n301 VSUBS 0.009551f
C453 B.n302 VSUBS 0.009551f
C454 B.n303 VSUBS 0.009551f
C455 B.n304 VSUBS 0.009551f
C456 B.n305 VSUBS 0.009551f
C457 B.n306 VSUBS 0.009551f
C458 B.n307 VSUBS 0.009551f
C459 B.n308 VSUBS 0.02042f
C460 B.n309 VSUBS 0.021716f
C461 B.n310 VSUBS 0.021716f
C462 B.n311 VSUBS 0.009551f
C463 B.n312 VSUBS 0.009551f
C464 B.n313 VSUBS 0.009551f
C465 B.n314 VSUBS 0.009551f
C466 B.n315 VSUBS 0.009551f
C467 B.n316 VSUBS 0.009551f
C468 B.n317 VSUBS 0.009551f
C469 B.n318 VSUBS 0.009551f
C470 B.n319 VSUBS 0.009551f
C471 B.n320 VSUBS 0.009551f
C472 B.n321 VSUBS 0.009551f
C473 B.n322 VSUBS 0.009551f
C474 B.n323 VSUBS 0.009551f
C475 B.n324 VSUBS 0.009551f
C476 B.n325 VSUBS 0.009551f
C477 B.n326 VSUBS 0.009551f
C478 B.n327 VSUBS 0.009551f
C479 B.n328 VSUBS 0.009551f
C480 B.n329 VSUBS 0.009551f
C481 B.n330 VSUBS 0.009551f
C482 B.n331 VSUBS 0.009551f
C483 B.n332 VSUBS 0.009551f
C484 B.n333 VSUBS 0.009551f
C485 B.n334 VSUBS 0.009551f
C486 B.n335 VSUBS 0.009551f
C487 B.n336 VSUBS 0.009551f
C488 B.n337 VSUBS 0.009551f
C489 B.n338 VSUBS 0.009551f
C490 B.n339 VSUBS 0.009551f
C491 B.n340 VSUBS 0.009551f
C492 B.n341 VSUBS 0.009551f
C493 B.n342 VSUBS 0.009551f
C494 B.n343 VSUBS 0.009551f
C495 B.n344 VSUBS 0.009551f
C496 B.n345 VSUBS 0.009551f
C497 B.n346 VSUBS 0.009551f
C498 B.n347 VSUBS 0.009551f
C499 B.n348 VSUBS 0.009551f
C500 B.n349 VSUBS 0.009551f
C501 B.n350 VSUBS 0.009551f
C502 B.n351 VSUBS 0.009551f
C503 B.n352 VSUBS 0.009551f
C504 B.n353 VSUBS 0.009551f
C505 B.n354 VSUBS 0.009551f
C506 B.n355 VSUBS 0.009551f
C507 B.n356 VSUBS 0.009551f
C508 B.n357 VSUBS 0.009551f
C509 B.n358 VSUBS 0.009551f
C510 B.n359 VSUBS 0.009551f
C511 B.n360 VSUBS 0.009551f
C512 B.n361 VSUBS 0.009551f
C513 B.n362 VSUBS 0.009551f
C514 B.n363 VSUBS 0.009551f
C515 B.n364 VSUBS 0.009551f
C516 B.n365 VSUBS 0.009551f
C517 B.n366 VSUBS 0.009551f
C518 B.n367 VSUBS 0.008989f
C519 B.n368 VSUBS 0.022128f
C520 B.n369 VSUBS 0.005337f
C521 B.n370 VSUBS 0.009551f
C522 B.n371 VSUBS 0.009551f
C523 B.n372 VSUBS 0.009551f
C524 B.n373 VSUBS 0.009551f
C525 B.n374 VSUBS 0.009551f
C526 B.n375 VSUBS 0.009551f
C527 B.n376 VSUBS 0.009551f
C528 B.n377 VSUBS 0.009551f
C529 B.n378 VSUBS 0.009551f
C530 B.n379 VSUBS 0.009551f
C531 B.n380 VSUBS 0.009551f
C532 B.n381 VSUBS 0.009551f
C533 B.t2 VSUBS 0.490735f
C534 B.t1 VSUBS 0.519811f
C535 B.t0 VSUBS 1.87339f
C536 B.n382 VSUBS 0.275193f
C537 B.n383 VSUBS 0.098385f
C538 B.n384 VSUBS 0.022128f
C539 B.n385 VSUBS 0.005337f
C540 B.n386 VSUBS 0.009551f
C541 B.n387 VSUBS 0.009551f
C542 B.n388 VSUBS 0.009551f
C543 B.n389 VSUBS 0.009551f
C544 B.n390 VSUBS 0.009551f
C545 B.n391 VSUBS 0.009551f
C546 B.n392 VSUBS 0.009551f
C547 B.n393 VSUBS 0.009551f
C548 B.n394 VSUBS 0.009551f
C549 B.n395 VSUBS 0.009551f
C550 B.n396 VSUBS 0.009551f
C551 B.n397 VSUBS 0.009551f
C552 B.n398 VSUBS 0.009551f
C553 B.n399 VSUBS 0.009551f
C554 B.n400 VSUBS 0.009551f
C555 B.n401 VSUBS 0.009551f
C556 B.n402 VSUBS 0.009551f
C557 B.n403 VSUBS 0.009551f
C558 B.n404 VSUBS 0.009551f
C559 B.n405 VSUBS 0.009551f
C560 B.n406 VSUBS 0.009551f
C561 B.n407 VSUBS 0.009551f
C562 B.n408 VSUBS 0.009551f
C563 B.n409 VSUBS 0.009551f
C564 B.n410 VSUBS 0.009551f
C565 B.n411 VSUBS 0.009551f
C566 B.n412 VSUBS 0.009551f
C567 B.n413 VSUBS 0.009551f
C568 B.n414 VSUBS 0.009551f
C569 B.n415 VSUBS 0.009551f
C570 B.n416 VSUBS 0.009551f
C571 B.n417 VSUBS 0.009551f
C572 B.n418 VSUBS 0.009551f
C573 B.n419 VSUBS 0.009551f
C574 B.n420 VSUBS 0.009551f
C575 B.n421 VSUBS 0.009551f
C576 B.n422 VSUBS 0.009551f
C577 B.n423 VSUBS 0.009551f
C578 B.n424 VSUBS 0.009551f
C579 B.n425 VSUBS 0.009551f
C580 B.n426 VSUBS 0.009551f
C581 B.n427 VSUBS 0.009551f
C582 B.n428 VSUBS 0.009551f
C583 B.n429 VSUBS 0.009551f
C584 B.n430 VSUBS 0.009551f
C585 B.n431 VSUBS 0.009551f
C586 B.n432 VSUBS 0.009551f
C587 B.n433 VSUBS 0.009551f
C588 B.n434 VSUBS 0.009551f
C589 B.n435 VSUBS 0.009551f
C590 B.n436 VSUBS 0.009551f
C591 B.n437 VSUBS 0.009551f
C592 B.n438 VSUBS 0.009551f
C593 B.n439 VSUBS 0.009551f
C594 B.n440 VSUBS 0.009551f
C595 B.n441 VSUBS 0.009551f
C596 B.n442 VSUBS 0.009551f
C597 B.n443 VSUBS 0.009551f
C598 B.n444 VSUBS 0.02048f
C599 B.n445 VSUBS 0.021656f
C600 B.n446 VSUBS 0.02042f
C601 B.n447 VSUBS 0.009551f
C602 B.n448 VSUBS 0.009551f
C603 B.n449 VSUBS 0.009551f
C604 B.n450 VSUBS 0.009551f
C605 B.n451 VSUBS 0.009551f
C606 B.n452 VSUBS 0.009551f
C607 B.n453 VSUBS 0.009551f
C608 B.n454 VSUBS 0.009551f
C609 B.n455 VSUBS 0.009551f
C610 B.n456 VSUBS 0.009551f
C611 B.n457 VSUBS 0.009551f
C612 B.n458 VSUBS 0.009551f
C613 B.n459 VSUBS 0.009551f
C614 B.n460 VSUBS 0.009551f
C615 B.n461 VSUBS 0.009551f
C616 B.n462 VSUBS 0.009551f
C617 B.n463 VSUBS 0.009551f
C618 B.n464 VSUBS 0.009551f
C619 B.n465 VSUBS 0.009551f
C620 B.n466 VSUBS 0.009551f
C621 B.n467 VSUBS 0.009551f
C622 B.n468 VSUBS 0.009551f
C623 B.n469 VSUBS 0.009551f
C624 B.n470 VSUBS 0.009551f
C625 B.n471 VSUBS 0.009551f
C626 B.n472 VSUBS 0.009551f
C627 B.n473 VSUBS 0.009551f
C628 B.n474 VSUBS 0.009551f
C629 B.n475 VSUBS 0.009551f
C630 B.n476 VSUBS 0.009551f
C631 B.n477 VSUBS 0.009551f
C632 B.n478 VSUBS 0.009551f
C633 B.n479 VSUBS 0.009551f
C634 B.n480 VSUBS 0.009551f
C635 B.n481 VSUBS 0.009551f
C636 B.n482 VSUBS 0.009551f
C637 B.n483 VSUBS 0.009551f
C638 B.n484 VSUBS 0.009551f
C639 B.n485 VSUBS 0.009551f
C640 B.n486 VSUBS 0.009551f
C641 B.n487 VSUBS 0.009551f
C642 B.n488 VSUBS 0.009551f
C643 B.n489 VSUBS 0.009551f
C644 B.n490 VSUBS 0.009551f
C645 B.n491 VSUBS 0.009551f
C646 B.n492 VSUBS 0.009551f
C647 B.n493 VSUBS 0.009551f
C648 B.n494 VSUBS 0.009551f
C649 B.n495 VSUBS 0.009551f
C650 B.n496 VSUBS 0.009551f
C651 B.n497 VSUBS 0.009551f
C652 B.n498 VSUBS 0.009551f
C653 B.n499 VSUBS 0.009551f
C654 B.n500 VSUBS 0.009551f
C655 B.n501 VSUBS 0.009551f
C656 B.n502 VSUBS 0.009551f
C657 B.n503 VSUBS 0.009551f
C658 B.n504 VSUBS 0.009551f
C659 B.n505 VSUBS 0.009551f
C660 B.n506 VSUBS 0.009551f
C661 B.n507 VSUBS 0.009551f
C662 B.n508 VSUBS 0.009551f
C663 B.n509 VSUBS 0.009551f
C664 B.n510 VSUBS 0.009551f
C665 B.n511 VSUBS 0.009551f
C666 B.n512 VSUBS 0.009551f
C667 B.n513 VSUBS 0.009551f
C668 B.n514 VSUBS 0.009551f
C669 B.n515 VSUBS 0.009551f
C670 B.n516 VSUBS 0.009551f
C671 B.n517 VSUBS 0.009551f
C672 B.n518 VSUBS 0.009551f
C673 B.n519 VSUBS 0.009551f
C674 B.n520 VSUBS 0.009551f
C675 B.n521 VSUBS 0.009551f
C676 B.n522 VSUBS 0.009551f
C677 B.n523 VSUBS 0.009551f
C678 B.n524 VSUBS 0.009551f
C679 B.n525 VSUBS 0.009551f
C680 B.n526 VSUBS 0.009551f
C681 B.n527 VSUBS 0.009551f
C682 B.n528 VSUBS 0.009551f
C683 B.n529 VSUBS 0.009551f
C684 B.n530 VSUBS 0.009551f
C685 B.n531 VSUBS 0.009551f
C686 B.n532 VSUBS 0.009551f
C687 B.n533 VSUBS 0.009551f
C688 B.n534 VSUBS 0.009551f
C689 B.n535 VSUBS 0.009551f
C690 B.n536 VSUBS 0.009551f
C691 B.n537 VSUBS 0.009551f
C692 B.n538 VSUBS 0.009551f
C693 B.n539 VSUBS 0.009551f
C694 B.n540 VSUBS 0.009551f
C695 B.n541 VSUBS 0.009551f
C696 B.n542 VSUBS 0.009551f
C697 B.n543 VSUBS 0.009551f
C698 B.n544 VSUBS 0.009551f
C699 B.n545 VSUBS 0.009551f
C700 B.n546 VSUBS 0.009551f
C701 B.n547 VSUBS 0.009551f
C702 B.n548 VSUBS 0.009551f
C703 B.n549 VSUBS 0.009551f
C704 B.n550 VSUBS 0.009551f
C705 B.n551 VSUBS 0.009551f
C706 B.n552 VSUBS 0.009551f
C707 B.n553 VSUBS 0.009551f
C708 B.n554 VSUBS 0.009551f
C709 B.n555 VSUBS 0.009551f
C710 B.n556 VSUBS 0.009551f
C711 B.n557 VSUBS 0.009551f
C712 B.n558 VSUBS 0.009551f
C713 B.n559 VSUBS 0.009551f
C714 B.n560 VSUBS 0.009551f
C715 B.n561 VSUBS 0.009551f
C716 B.n562 VSUBS 0.009551f
C717 B.n563 VSUBS 0.009551f
C718 B.n564 VSUBS 0.009551f
C719 B.n565 VSUBS 0.009551f
C720 B.n566 VSUBS 0.009551f
C721 B.n567 VSUBS 0.009551f
C722 B.n568 VSUBS 0.009551f
C723 B.n569 VSUBS 0.009551f
C724 B.n570 VSUBS 0.009551f
C725 B.n571 VSUBS 0.009551f
C726 B.n572 VSUBS 0.009551f
C727 B.n573 VSUBS 0.009551f
C728 B.n574 VSUBS 0.009551f
C729 B.n575 VSUBS 0.009551f
C730 B.n576 VSUBS 0.009551f
C731 B.n577 VSUBS 0.009551f
C732 B.n578 VSUBS 0.009551f
C733 B.n579 VSUBS 0.009551f
C734 B.n580 VSUBS 0.009551f
C735 B.n581 VSUBS 0.009551f
C736 B.n582 VSUBS 0.009551f
C737 B.n583 VSUBS 0.009551f
C738 B.n584 VSUBS 0.009551f
C739 B.n585 VSUBS 0.009551f
C740 B.n586 VSUBS 0.009551f
C741 B.n587 VSUBS 0.009551f
C742 B.n588 VSUBS 0.009551f
C743 B.n589 VSUBS 0.009551f
C744 B.n590 VSUBS 0.009551f
C745 B.n591 VSUBS 0.009551f
C746 B.n592 VSUBS 0.009551f
C747 B.n593 VSUBS 0.009551f
C748 B.n594 VSUBS 0.009551f
C749 B.n595 VSUBS 0.009551f
C750 B.n596 VSUBS 0.009551f
C751 B.n597 VSUBS 0.009551f
C752 B.n598 VSUBS 0.009551f
C753 B.n599 VSUBS 0.009551f
C754 B.n600 VSUBS 0.009551f
C755 B.n601 VSUBS 0.009551f
C756 B.n602 VSUBS 0.009551f
C757 B.n603 VSUBS 0.009551f
C758 B.n604 VSUBS 0.009551f
C759 B.n605 VSUBS 0.009551f
C760 B.n606 VSUBS 0.009551f
C761 B.n607 VSUBS 0.009551f
C762 B.n608 VSUBS 0.009551f
C763 B.n609 VSUBS 0.009551f
C764 B.n610 VSUBS 0.009551f
C765 B.n611 VSUBS 0.009551f
C766 B.n612 VSUBS 0.009551f
C767 B.n613 VSUBS 0.009551f
C768 B.n614 VSUBS 0.009551f
C769 B.n615 VSUBS 0.009551f
C770 B.n616 VSUBS 0.009551f
C771 B.n617 VSUBS 0.009551f
C772 B.n618 VSUBS 0.009551f
C773 B.n619 VSUBS 0.009551f
C774 B.n620 VSUBS 0.009551f
C775 B.n621 VSUBS 0.009551f
C776 B.n622 VSUBS 0.009551f
C777 B.n623 VSUBS 0.009551f
C778 B.n624 VSUBS 0.009551f
C779 B.n625 VSUBS 0.009551f
C780 B.n626 VSUBS 0.009551f
C781 B.n627 VSUBS 0.009551f
C782 B.n628 VSUBS 0.009551f
C783 B.n629 VSUBS 0.009551f
C784 B.n630 VSUBS 0.02042f
C785 B.n631 VSUBS 0.021716f
C786 B.n632 VSUBS 0.021716f
C787 B.n633 VSUBS 0.009551f
C788 B.n634 VSUBS 0.009551f
C789 B.n635 VSUBS 0.009551f
C790 B.n636 VSUBS 0.009551f
C791 B.n637 VSUBS 0.009551f
C792 B.n638 VSUBS 0.009551f
C793 B.n639 VSUBS 0.009551f
C794 B.n640 VSUBS 0.009551f
C795 B.n641 VSUBS 0.009551f
C796 B.n642 VSUBS 0.009551f
C797 B.n643 VSUBS 0.009551f
C798 B.n644 VSUBS 0.009551f
C799 B.n645 VSUBS 0.009551f
C800 B.n646 VSUBS 0.009551f
C801 B.n647 VSUBS 0.009551f
C802 B.n648 VSUBS 0.009551f
C803 B.n649 VSUBS 0.009551f
C804 B.n650 VSUBS 0.009551f
C805 B.n651 VSUBS 0.009551f
C806 B.n652 VSUBS 0.009551f
C807 B.n653 VSUBS 0.009551f
C808 B.n654 VSUBS 0.009551f
C809 B.n655 VSUBS 0.009551f
C810 B.n656 VSUBS 0.009551f
C811 B.n657 VSUBS 0.009551f
C812 B.n658 VSUBS 0.009551f
C813 B.n659 VSUBS 0.009551f
C814 B.n660 VSUBS 0.009551f
C815 B.n661 VSUBS 0.009551f
C816 B.n662 VSUBS 0.009551f
C817 B.n663 VSUBS 0.009551f
C818 B.n664 VSUBS 0.009551f
C819 B.n665 VSUBS 0.009551f
C820 B.n666 VSUBS 0.009551f
C821 B.n667 VSUBS 0.009551f
C822 B.n668 VSUBS 0.009551f
C823 B.n669 VSUBS 0.009551f
C824 B.n670 VSUBS 0.009551f
C825 B.n671 VSUBS 0.009551f
C826 B.n672 VSUBS 0.009551f
C827 B.n673 VSUBS 0.009551f
C828 B.n674 VSUBS 0.009551f
C829 B.n675 VSUBS 0.009551f
C830 B.n676 VSUBS 0.009551f
C831 B.n677 VSUBS 0.009551f
C832 B.n678 VSUBS 0.009551f
C833 B.n679 VSUBS 0.009551f
C834 B.n680 VSUBS 0.009551f
C835 B.n681 VSUBS 0.009551f
C836 B.n682 VSUBS 0.009551f
C837 B.n683 VSUBS 0.009551f
C838 B.n684 VSUBS 0.009551f
C839 B.n685 VSUBS 0.009551f
C840 B.n686 VSUBS 0.009551f
C841 B.n687 VSUBS 0.009551f
C842 B.n688 VSUBS 0.009551f
C843 B.n689 VSUBS 0.008989f
C844 B.n690 VSUBS 0.022128f
C845 B.n691 VSUBS 0.005337f
C846 B.n692 VSUBS 0.009551f
C847 B.n693 VSUBS 0.009551f
C848 B.n694 VSUBS 0.009551f
C849 B.n695 VSUBS 0.009551f
C850 B.n696 VSUBS 0.009551f
C851 B.n697 VSUBS 0.009551f
C852 B.n698 VSUBS 0.009551f
C853 B.n699 VSUBS 0.009551f
C854 B.n700 VSUBS 0.009551f
C855 B.n701 VSUBS 0.009551f
C856 B.n702 VSUBS 0.009551f
C857 B.n703 VSUBS 0.009551f
C858 B.n704 VSUBS 0.005337f
C859 B.n705 VSUBS 0.009551f
C860 B.n706 VSUBS 0.009551f
C861 B.n707 VSUBS 0.008989f
C862 B.n708 VSUBS 0.009551f
C863 B.n709 VSUBS 0.009551f
C864 B.n710 VSUBS 0.009551f
C865 B.n711 VSUBS 0.009551f
C866 B.n712 VSUBS 0.009551f
C867 B.n713 VSUBS 0.009551f
C868 B.n714 VSUBS 0.009551f
C869 B.n715 VSUBS 0.009551f
C870 B.n716 VSUBS 0.009551f
C871 B.n717 VSUBS 0.009551f
C872 B.n718 VSUBS 0.009551f
C873 B.n719 VSUBS 0.009551f
C874 B.n720 VSUBS 0.009551f
C875 B.n721 VSUBS 0.009551f
C876 B.n722 VSUBS 0.009551f
C877 B.n723 VSUBS 0.009551f
C878 B.n724 VSUBS 0.009551f
C879 B.n725 VSUBS 0.009551f
C880 B.n726 VSUBS 0.009551f
C881 B.n727 VSUBS 0.009551f
C882 B.n728 VSUBS 0.009551f
C883 B.n729 VSUBS 0.009551f
C884 B.n730 VSUBS 0.009551f
C885 B.n731 VSUBS 0.009551f
C886 B.n732 VSUBS 0.009551f
C887 B.n733 VSUBS 0.009551f
C888 B.n734 VSUBS 0.009551f
C889 B.n735 VSUBS 0.009551f
C890 B.n736 VSUBS 0.009551f
C891 B.n737 VSUBS 0.009551f
C892 B.n738 VSUBS 0.009551f
C893 B.n739 VSUBS 0.009551f
C894 B.n740 VSUBS 0.009551f
C895 B.n741 VSUBS 0.009551f
C896 B.n742 VSUBS 0.009551f
C897 B.n743 VSUBS 0.009551f
C898 B.n744 VSUBS 0.009551f
C899 B.n745 VSUBS 0.009551f
C900 B.n746 VSUBS 0.009551f
C901 B.n747 VSUBS 0.009551f
C902 B.n748 VSUBS 0.009551f
C903 B.n749 VSUBS 0.009551f
C904 B.n750 VSUBS 0.009551f
C905 B.n751 VSUBS 0.009551f
C906 B.n752 VSUBS 0.009551f
C907 B.n753 VSUBS 0.009551f
C908 B.n754 VSUBS 0.009551f
C909 B.n755 VSUBS 0.009551f
C910 B.n756 VSUBS 0.009551f
C911 B.n757 VSUBS 0.009551f
C912 B.n758 VSUBS 0.009551f
C913 B.n759 VSUBS 0.009551f
C914 B.n760 VSUBS 0.009551f
C915 B.n761 VSUBS 0.009551f
C916 B.n762 VSUBS 0.009551f
C917 B.n763 VSUBS 0.021716f
C918 B.n764 VSUBS 0.021716f
C919 B.n765 VSUBS 0.02042f
C920 B.n766 VSUBS 0.009551f
C921 B.n767 VSUBS 0.009551f
C922 B.n768 VSUBS 0.009551f
C923 B.n769 VSUBS 0.009551f
C924 B.n770 VSUBS 0.009551f
C925 B.n771 VSUBS 0.009551f
C926 B.n772 VSUBS 0.009551f
C927 B.n773 VSUBS 0.009551f
C928 B.n774 VSUBS 0.009551f
C929 B.n775 VSUBS 0.009551f
C930 B.n776 VSUBS 0.009551f
C931 B.n777 VSUBS 0.009551f
C932 B.n778 VSUBS 0.009551f
C933 B.n779 VSUBS 0.009551f
C934 B.n780 VSUBS 0.009551f
C935 B.n781 VSUBS 0.009551f
C936 B.n782 VSUBS 0.009551f
C937 B.n783 VSUBS 0.009551f
C938 B.n784 VSUBS 0.009551f
C939 B.n785 VSUBS 0.009551f
C940 B.n786 VSUBS 0.009551f
C941 B.n787 VSUBS 0.009551f
C942 B.n788 VSUBS 0.009551f
C943 B.n789 VSUBS 0.009551f
C944 B.n790 VSUBS 0.009551f
C945 B.n791 VSUBS 0.009551f
C946 B.n792 VSUBS 0.009551f
C947 B.n793 VSUBS 0.009551f
C948 B.n794 VSUBS 0.009551f
C949 B.n795 VSUBS 0.009551f
C950 B.n796 VSUBS 0.009551f
C951 B.n797 VSUBS 0.009551f
C952 B.n798 VSUBS 0.009551f
C953 B.n799 VSUBS 0.009551f
C954 B.n800 VSUBS 0.009551f
C955 B.n801 VSUBS 0.009551f
C956 B.n802 VSUBS 0.009551f
C957 B.n803 VSUBS 0.009551f
C958 B.n804 VSUBS 0.009551f
C959 B.n805 VSUBS 0.009551f
C960 B.n806 VSUBS 0.009551f
C961 B.n807 VSUBS 0.009551f
C962 B.n808 VSUBS 0.009551f
C963 B.n809 VSUBS 0.009551f
C964 B.n810 VSUBS 0.009551f
C965 B.n811 VSUBS 0.009551f
C966 B.n812 VSUBS 0.009551f
C967 B.n813 VSUBS 0.009551f
C968 B.n814 VSUBS 0.009551f
C969 B.n815 VSUBS 0.009551f
C970 B.n816 VSUBS 0.009551f
C971 B.n817 VSUBS 0.009551f
C972 B.n818 VSUBS 0.009551f
C973 B.n819 VSUBS 0.009551f
C974 B.n820 VSUBS 0.009551f
C975 B.n821 VSUBS 0.009551f
C976 B.n822 VSUBS 0.009551f
C977 B.n823 VSUBS 0.009551f
C978 B.n824 VSUBS 0.009551f
C979 B.n825 VSUBS 0.009551f
C980 B.n826 VSUBS 0.009551f
C981 B.n827 VSUBS 0.009551f
C982 B.n828 VSUBS 0.009551f
C983 B.n829 VSUBS 0.009551f
C984 B.n830 VSUBS 0.009551f
C985 B.n831 VSUBS 0.009551f
C986 B.n832 VSUBS 0.009551f
C987 B.n833 VSUBS 0.009551f
C988 B.n834 VSUBS 0.009551f
C989 B.n835 VSUBS 0.009551f
C990 B.n836 VSUBS 0.009551f
C991 B.n837 VSUBS 0.009551f
C992 B.n838 VSUBS 0.009551f
C993 B.n839 VSUBS 0.009551f
C994 B.n840 VSUBS 0.009551f
C995 B.n841 VSUBS 0.009551f
C996 B.n842 VSUBS 0.009551f
C997 B.n843 VSUBS 0.009551f
C998 B.n844 VSUBS 0.009551f
C999 B.n845 VSUBS 0.009551f
C1000 B.n846 VSUBS 0.009551f
C1001 B.n847 VSUBS 0.009551f
C1002 B.n848 VSUBS 0.009551f
C1003 B.n849 VSUBS 0.009551f
C1004 B.n850 VSUBS 0.009551f
C1005 B.n851 VSUBS 0.009551f
C1006 B.n852 VSUBS 0.009551f
C1007 B.n853 VSUBS 0.009551f
C1008 B.n854 VSUBS 0.009551f
C1009 B.n855 VSUBS 0.012463f
C1010 B.n856 VSUBS 0.013277f
C1011 B.n857 VSUBS 0.026402f
C1012 VTAIL.t1 VSUBS 0.258409f
C1013 VTAIL.t3 VSUBS 0.258409f
C1014 VTAIL.n0 VSUBS 1.84953f
C1015 VTAIL.n1 VSUBS 1.00217f
C1016 VTAIL.t11 VSUBS 2.44834f
C1017 VTAIL.n2 VSUBS 1.16422f
C1018 VTAIL.t9 VSUBS 0.258409f
C1019 VTAIL.t18 VSUBS 0.258409f
C1020 VTAIL.n3 VSUBS 1.84953f
C1021 VTAIL.n4 VSUBS 1.13703f
C1022 VTAIL.t15 VSUBS 0.258409f
C1023 VTAIL.t17 VSUBS 0.258409f
C1024 VTAIL.n5 VSUBS 1.84953f
C1025 VTAIL.n6 VSUBS 2.69094f
C1026 VTAIL.t0 VSUBS 0.258409f
C1027 VTAIL.t19 VSUBS 0.258409f
C1028 VTAIL.n7 VSUBS 1.84954f
C1029 VTAIL.n8 VSUBS 2.69094f
C1030 VTAIL.t4 VSUBS 0.258409f
C1031 VTAIL.t8 VSUBS 0.258409f
C1032 VTAIL.n9 VSUBS 1.84954f
C1033 VTAIL.n10 VSUBS 1.13702f
C1034 VTAIL.t6 VSUBS 2.44836f
C1035 VTAIL.n11 VSUBS 1.1642f
C1036 VTAIL.t13 VSUBS 0.258409f
C1037 VTAIL.t14 VSUBS 0.258409f
C1038 VTAIL.n12 VSUBS 1.84954f
C1039 VTAIL.n13 VSUBS 1.05827f
C1040 VTAIL.t16 VSUBS 0.258409f
C1041 VTAIL.t10 VSUBS 0.258409f
C1042 VTAIL.n14 VSUBS 1.84954f
C1043 VTAIL.n15 VSUBS 1.13702f
C1044 VTAIL.t12 VSUBS 2.44834f
C1045 VTAIL.n16 VSUBS 2.55042f
C1046 VTAIL.t5 VSUBS 2.44834f
C1047 VTAIL.n17 VSUBS 2.55042f
C1048 VTAIL.t2 VSUBS 0.258409f
C1049 VTAIL.t7 VSUBS 0.258409f
C1050 VTAIL.n18 VSUBS 1.84953f
C1051 VTAIL.n19 VSUBS 0.946669f
C1052 VDD1.t7 VSUBS 2.73369f
C1053 VDD1.t1 VSUBS 0.267596f
C1054 VDD1.t6 VSUBS 0.267596f
C1055 VDD1.n0 VSUBS 2.06737f
C1056 VDD1.n1 VSUBS 1.76824f
C1057 VDD1.t2 VSUBS 2.73368f
C1058 VDD1.t0 VSUBS 0.267596f
C1059 VDD1.t4 VSUBS 0.267596f
C1060 VDD1.n2 VSUBS 2.06737f
C1061 VDD1.n3 VSUBS 1.75831f
C1062 VDD1.t9 VSUBS 0.267596f
C1063 VDD1.t8 VSUBS 0.267596f
C1064 VDD1.n4 VSUBS 2.09164f
C1065 VDD1.n5 VSUBS 3.9843f
C1066 VDD1.t3 VSUBS 0.267596f
C1067 VDD1.t5 VSUBS 0.267596f
C1068 VDD1.n6 VSUBS 2.06736f
C1069 VDD1.n7 VSUBS 4.13204f
C1070 VP.n0 VSUBS 0.040657f
C1071 VP.t7 VSUBS 2.51f
C1072 VP.n1 VSUBS 0.060196f
C1073 VP.n2 VSUBS 0.030838f
C1074 VP.t0 VSUBS 2.51f
C1075 VP.n3 VSUBS 0.890872f
C1076 VP.n4 VSUBS 0.030838f
C1077 VP.n5 VSUBS 0.024969f
C1078 VP.n6 VSUBS 0.030838f
C1079 VP.t9 VSUBS 2.51f
C1080 VP.n7 VSUBS 0.057475f
C1081 VP.n8 VSUBS 0.030838f
C1082 VP.n9 VSUBS 0.057475f
C1083 VP.n10 VSUBS 0.030838f
C1084 VP.t1 VSUBS 2.51f
C1085 VP.n11 VSUBS 0.025288f
C1086 VP.n12 VSUBS 0.030838f
C1087 VP.t3 VSUBS 2.51f
C1088 VP.n13 VSUBS 0.984788f
C1089 VP.n14 VSUBS 0.040657f
C1090 VP.t6 VSUBS 2.51f
C1091 VP.n15 VSUBS 0.060196f
C1092 VP.n16 VSUBS 0.030838f
C1093 VP.t8 VSUBS 2.51f
C1094 VP.n17 VSUBS 0.890872f
C1095 VP.n18 VSUBS 0.030838f
C1096 VP.n19 VSUBS 0.024969f
C1097 VP.n20 VSUBS 0.030838f
C1098 VP.t2 VSUBS 2.51f
C1099 VP.n21 VSUBS 0.057475f
C1100 VP.n22 VSUBS 0.030838f
C1101 VP.n23 VSUBS 0.057475f
C1102 VP.t5 VSUBS 2.76481f
C1103 VP.n24 VSUBS 0.958802f
C1104 VP.t4 VSUBS 2.51f
C1105 VP.n25 VSUBS 0.971209f
C1106 VP.n26 VSUBS 0.030234f
C1107 VP.n27 VSUBS 0.300296f
C1108 VP.n28 VSUBS 0.030838f
C1109 VP.n29 VSUBS 0.030838f
C1110 VP.n30 VSUBS 0.060962f
C1111 VP.n31 VSUBS 0.024969f
C1112 VP.n32 VSUBS 0.06158f
C1113 VP.n33 VSUBS 0.030838f
C1114 VP.n34 VSUBS 0.030838f
C1115 VP.n35 VSUBS 0.030838f
C1116 VP.n36 VSUBS 0.919971f
C1117 VP.n37 VSUBS 0.057475f
C1118 VP.n38 VSUBS 0.06158f
C1119 VP.n39 VSUBS 0.030838f
C1120 VP.n40 VSUBS 0.030838f
C1121 VP.n41 VSUBS 0.030838f
C1122 VP.n42 VSUBS 0.060962f
C1123 VP.n43 VSUBS 0.057475f
C1124 VP.n44 VSUBS 0.030234f
C1125 VP.n45 VSUBS 0.030838f
C1126 VP.n46 VSUBS 0.030838f
C1127 VP.n47 VSUBS 0.05634f
C1128 VP.n48 VSUBS 0.062027f
C1129 VP.n49 VSUBS 0.025288f
C1130 VP.n50 VSUBS 0.030838f
C1131 VP.n51 VSUBS 0.030838f
C1132 VP.n52 VSUBS 0.030838f
C1133 VP.n53 VSUBS 0.057475f
C1134 VP.n54 VSUBS 0.031369f
C1135 VP.n55 VSUBS 0.984788f
C1136 VP.n56 VSUBS 1.86578f
C1137 VP.n57 VSUBS 1.88675f
C1138 VP.n58 VSUBS 0.040657f
C1139 VP.n59 VSUBS 0.031369f
C1140 VP.n60 VSUBS 0.057475f
C1141 VP.n61 VSUBS 0.060196f
C1142 VP.n62 VSUBS 0.030838f
C1143 VP.n63 VSUBS 0.030838f
C1144 VP.n64 VSUBS 0.030838f
C1145 VP.n65 VSUBS 0.062027f
C1146 VP.n66 VSUBS 0.05634f
C1147 VP.n67 VSUBS 0.890872f
C1148 VP.n68 VSUBS 0.030234f
C1149 VP.n69 VSUBS 0.030838f
C1150 VP.n70 VSUBS 0.030838f
C1151 VP.n71 VSUBS 0.030838f
C1152 VP.n72 VSUBS 0.060962f
C1153 VP.n73 VSUBS 0.024969f
C1154 VP.n74 VSUBS 0.06158f
C1155 VP.n75 VSUBS 0.030838f
C1156 VP.n76 VSUBS 0.030838f
C1157 VP.n77 VSUBS 0.030838f
C1158 VP.n78 VSUBS 0.919971f
C1159 VP.n79 VSUBS 0.057475f
C1160 VP.n80 VSUBS 0.06158f
C1161 VP.n81 VSUBS 0.030838f
C1162 VP.n82 VSUBS 0.030838f
C1163 VP.n83 VSUBS 0.030838f
C1164 VP.n84 VSUBS 0.060962f
C1165 VP.n85 VSUBS 0.057475f
C1166 VP.n86 VSUBS 0.030234f
C1167 VP.n87 VSUBS 0.030838f
C1168 VP.n88 VSUBS 0.030838f
C1169 VP.n89 VSUBS 0.05634f
C1170 VP.n90 VSUBS 0.062027f
C1171 VP.n91 VSUBS 0.025288f
C1172 VP.n92 VSUBS 0.030838f
C1173 VP.n93 VSUBS 0.030838f
C1174 VP.n94 VSUBS 0.030838f
C1175 VP.n95 VSUBS 0.057475f
C1176 VP.n96 VSUBS 0.031369f
C1177 VP.n97 VSUBS 0.984788f
C1178 VP.n98 VSUBS 0.056714f
.ends

