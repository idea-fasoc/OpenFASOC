* NGSPICE file created from diff_pair_sample_1793.ext - technology: sky130A

.subckt diff_pair_sample_1793 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t19 VP.t0 VDD1.t3 w_n4486_n4508# sky130_fd_pr__pfet_01v8 ad=2.9205 pd=18.03 as=2.9205 ps=18.03 w=17.7 l=2.6
X1 VTAIL.t18 VP.t1 VDD1.t2 w_n4486_n4508# sky130_fd_pr__pfet_01v8 ad=2.9205 pd=18.03 as=2.9205 ps=18.03 w=17.7 l=2.6
X2 B.t11 B.t9 B.t10 w_n4486_n4508# sky130_fd_pr__pfet_01v8 ad=6.903 pd=36.18 as=0 ps=0 w=17.7 l=2.6
X3 VDD2.t9 VN.t0 VTAIL.t7 w_n4486_n4508# sky130_fd_pr__pfet_01v8 ad=2.9205 pd=18.03 as=2.9205 ps=18.03 w=17.7 l=2.6
X4 VDD2.t8 VN.t1 VTAIL.t6 w_n4486_n4508# sky130_fd_pr__pfet_01v8 ad=2.9205 pd=18.03 as=6.903 ps=36.18 w=17.7 l=2.6
X5 VDD2.t7 VN.t2 VTAIL.t4 w_n4486_n4508# sky130_fd_pr__pfet_01v8 ad=6.903 pd=36.18 as=2.9205 ps=18.03 w=17.7 l=2.6
X6 B.t8 B.t6 B.t7 w_n4486_n4508# sky130_fd_pr__pfet_01v8 ad=6.903 pd=36.18 as=0 ps=0 w=17.7 l=2.6
X7 B.t5 B.t3 B.t4 w_n4486_n4508# sky130_fd_pr__pfet_01v8 ad=6.903 pd=36.18 as=0 ps=0 w=17.7 l=2.6
X8 B.t2 B.t0 B.t1 w_n4486_n4508# sky130_fd_pr__pfet_01v8 ad=6.903 pd=36.18 as=0 ps=0 w=17.7 l=2.6
X9 VDD2.t6 VN.t3 VTAIL.t5 w_n4486_n4508# sky130_fd_pr__pfet_01v8 ad=6.903 pd=36.18 as=2.9205 ps=18.03 w=17.7 l=2.6
X10 VTAIL.t9 VN.t4 VDD2.t5 w_n4486_n4508# sky130_fd_pr__pfet_01v8 ad=2.9205 pd=18.03 as=2.9205 ps=18.03 w=17.7 l=2.6
X11 VDD2.t4 VN.t5 VTAIL.t3 w_n4486_n4508# sky130_fd_pr__pfet_01v8 ad=2.9205 pd=18.03 as=2.9205 ps=18.03 w=17.7 l=2.6
X12 VTAIL.t0 VN.t6 VDD2.t3 w_n4486_n4508# sky130_fd_pr__pfet_01v8 ad=2.9205 pd=18.03 as=2.9205 ps=18.03 w=17.7 l=2.6
X13 VTAIL.t17 VP.t2 VDD1.t1 w_n4486_n4508# sky130_fd_pr__pfet_01v8 ad=2.9205 pd=18.03 as=2.9205 ps=18.03 w=17.7 l=2.6
X14 VDD1.t0 VP.t3 VTAIL.t16 w_n4486_n4508# sky130_fd_pr__pfet_01v8 ad=6.903 pd=36.18 as=2.9205 ps=18.03 w=17.7 l=2.6
X15 VDD1.t7 VP.t4 VTAIL.t15 w_n4486_n4508# sky130_fd_pr__pfet_01v8 ad=6.903 pd=36.18 as=2.9205 ps=18.03 w=17.7 l=2.6
X16 VTAIL.t8 VN.t7 VDD2.t2 w_n4486_n4508# sky130_fd_pr__pfet_01v8 ad=2.9205 pd=18.03 as=2.9205 ps=18.03 w=17.7 l=2.6
X17 VDD2.t1 VN.t8 VTAIL.t2 w_n4486_n4508# sky130_fd_pr__pfet_01v8 ad=2.9205 pd=18.03 as=6.903 ps=36.18 w=17.7 l=2.6
X18 VTAIL.t14 VP.t5 VDD1.t6 w_n4486_n4508# sky130_fd_pr__pfet_01v8 ad=2.9205 pd=18.03 as=2.9205 ps=18.03 w=17.7 l=2.6
X19 VDD1.t9 VP.t6 VTAIL.t13 w_n4486_n4508# sky130_fd_pr__pfet_01v8 ad=2.9205 pd=18.03 as=2.9205 ps=18.03 w=17.7 l=2.6
X20 VDD1.t8 VP.t7 VTAIL.t12 w_n4486_n4508# sky130_fd_pr__pfet_01v8 ad=2.9205 pd=18.03 as=2.9205 ps=18.03 w=17.7 l=2.6
X21 VDD1.t5 VP.t8 VTAIL.t11 w_n4486_n4508# sky130_fd_pr__pfet_01v8 ad=2.9205 pd=18.03 as=6.903 ps=36.18 w=17.7 l=2.6
X22 VTAIL.t1 VN.t9 VDD2.t0 w_n4486_n4508# sky130_fd_pr__pfet_01v8 ad=2.9205 pd=18.03 as=2.9205 ps=18.03 w=17.7 l=2.6
X23 VDD1.t4 VP.t9 VTAIL.t10 w_n4486_n4508# sky130_fd_pr__pfet_01v8 ad=2.9205 pd=18.03 as=6.903 ps=36.18 w=17.7 l=2.6
R0 VP.n24 VP.t4 196.298
R1 VP.n56 VP.t3 164.065
R2 VP.n64 VP.t5 164.065
R3 VP.n76 VP.t6 164.065
R4 VP.n3 VP.t1 164.065
R5 VP.n95 VP.t9 164.065
R6 VP.n53 VP.t8 164.065
R7 VP.n16 VP.t2 164.065
R8 VP.n34 VP.t7 164.065
R9 VP.n23 VP.t0 164.065
R10 VP.n25 VP.n22 161.3
R11 VP.n27 VP.n26 161.3
R12 VP.n28 VP.n21 161.3
R13 VP.n30 VP.n29 161.3
R14 VP.n31 VP.n20 161.3
R15 VP.n33 VP.n32 161.3
R16 VP.n35 VP.n19 161.3
R17 VP.n37 VP.n36 161.3
R18 VP.n38 VP.n18 161.3
R19 VP.n40 VP.n39 161.3
R20 VP.n41 VP.n17 161.3
R21 VP.n43 VP.n42 161.3
R22 VP.n45 VP.n44 161.3
R23 VP.n46 VP.n15 161.3
R24 VP.n48 VP.n47 161.3
R25 VP.n49 VP.n14 161.3
R26 VP.n51 VP.n50 161.3
R27 VP.n52 VP.n13 161.3
R28 VP.n94 VP.n0 161.3
R29 VP.n93 VP.n92 161.3
R30 VP.n91 VP.n1 161.3
R31 VP.n90 VP.n89 161.3
R32 VP.n88 VP.n2 161.3
R33 VP.n87 VP.n86 161.3
R34 VP.n85 VP.n84 161.3
R35 VP.n83 VP.n4 161.3
R36 VP.n82 VP.n81 161.3
R37 VP.n80 VP.n5 161.3
R38 VP.n79 VP.n78 161.3
R39 VP.n77 VP.n6 161.3
R40 VP.n75 VP.n74 161.3
R41 VP.n73 VP.n7 161.3
R42 VP.n72 VP.n71 161.3
R43 VP.n70 VP.n8 161.3
R44 VP.n69 VP.n68 161.3
R45 VP.n67 VP.n9 161.3
R46 VP.n66 VP.n65 161.3
R47 VP.n63 VP.n10 161.3
R48 VP.n62 VP.n61 161.3
R49 VP.n60 VP.n11 161.3
R50 VP.n59 VP.n58 161.3
R51 VP.n57 VP.n12 161.3
R52 VP.n56 VP.n55 105.499
R53 VP.n96 VP.n95 105.499
R54 VP.n54 VP.n53 105.499
R55 VP.n24 VP.n23 63.762
R56 VP.n55 VP.n54 57.3822
R57 VP.n71 VP.n70 56.5617
R58 VP.n40 VP.n18 56.5617
R59 VP.n82 VP.n5 56.5617
R60 VP.n29 VP.n28 56.5617
R61 VP.n62 VP.n11 54.6242
R62 VP.n89 VP.n1 54.6242
R63 VP.n47 VP.n14 54.6242
R64 VP.n63 VP.n62 26.5299
R65 VP.n89 VP.n88 26.5299
R66 VP.n47 VP.n46 26.5299
R67 VP.n58 VP.n57 24.5923
R68 VP.n58 VP.n11 24.5923
R69 VP.n65 VP.n63 24.5923
R70 VP.n69 VP.n9 24.5923
R71 VP.n70 VP.n69 24.5923
R72 VP.n71 VP.n7 24.5923
R73 VP.n75 VP.n7 24.5923
R74 VP.n78 VP.n77 24.5923
R75 VP.n78 VP.n5 24.5923
R76 VP.n83 VP.n82 24.5923
R77 VP.n84 VP.n83 24.5923
R78 VP.n88 VP.n87 24.5923
R79 VP.n93 VP.n1 24.5923
R80 VP.n94 VP.n93 24.5923
R81 VP.n51 VP.n14 24.5923
R82 VP.n52 VP.n51 24.5923
R83 VP.n41 VP.n40 24.5923
R84 VP.n42 VP.n41 24.5923
R85 VP.n46 VP.n45 24.5923
R86 VP.n29 VP.n20 24.5923
R87 VP.n33 VP.n20 24.5923
R88 VP.n36 VP.n35 24.5923
R89 VP.n36 VP.n18 24.5923
R90 VP.n27 VP.n22 24.5923
R91 VP.n28 VP.n27 24.5923
R92 VP.n65 VP.n64 15.7393
R93 VP.n87 VP.n3 15.7393
R94 VP.n45 VP.n16 15.7393
R95 VP.n76 VP.n75 12.2964
R96 VP.n77 VP.n76 12.2964
R97 VP.n34 VP.n33 12.2964
R98 VP.n35 VP.n34 12.2964
R99 VP.n64 VP.n9 8.85356
R100 VP.n84 VP.n3 8.85356
R101 VP.n42 VP.n16 8.85356
R102 VP.n23 VP.n22 8.85356
R103 VP.n25 VP.n24 7.12066
R104 VP.n57 VP.n56 5.4107
R105 VP.n95 VP.n94 5.4107
R106 VP.n53 VP.n52 5.4107
R107 VP.n54 VP.n13 0.278335
R108 VP.n55 VP.n12 0.278335
R109 VP.n96 VP.n0 0.278335
R110 VP.n26 VP.n25 0.189894
R111 VP.n26 VP.n21 0.189894
R112 VP.n30 VP.n21 0.189894
R113 VP.n31 VP.n30 0.189894
R114 VP.n32 VP.n31 0.189894
R115 VP.n32 VP.n19 0.189894
R116 VP.n37 VP.n19 0.189894
R117 VP.n38 VP.n37 0.189894
R118 VP.n39 VP.n38 0.189894
R119 VP.n39 VP.n17 0.189894
R120 VP.n43 VP.n17 0.189894
R121 VP.n44 VP.n43 0.189894
R122 VP.n44 VP.n15 0.189894
R123 VP.n48 VP.n15 0.189894
R124 VP.n49 VP.n48 0.189894
R125 VP.n50 VP.n49 0.189894
R126 VP.n50 VP.n13 0.189894
R127 VP.n59 VP.n12 0.189894
R128 VP.n60 VP.n59 0.189894
R129 VP.n61 VP.n60 0.189894
R130 VP.n61 VP.n10 0.189894
R131 VP.n66 VP.n10 0.189894
R132 VP.n67 VP.n66 0.189894
R133 VP.n68 VP.n67 0.189894
R134 VP.n68 VP.n8 0.189894
R135 VP.n72 VP.n8 0.189894
R136 VP.n73 VP.n72 0.189894
R137 VP.n74 VP.n73 0.189894
R138 VP.n74 VP.n6 0.189894
R139 VP.n79 VP.n6 0.189894
R140 VP.n80 VP.n79 0.189894
R141 VP.n81 VP.n80 0.189894
R142 VP.n81 VP.n4 0.189894
R143 VP.n85 VP.n4 0.189894
R144 VP.n86 VP.n85 0.189894
R145 VP.n86 VP.n2 0.189894
R146 VP.n90 VP.n2 0.189894
R147 VP.n91 VP.n90 0.189894
R148 VP.n92 VP.n91 0.189894
R149 VP.n92 VP.n0 0.189894
R150 VP VP.n96 0.153485
R151 VDD1.n1 VDD1.t7 76.3276
R152 VDD1.n3 VDD1.t0 76.3266
R153 VDD1.n5 VDD1.n4 73.8033
R154 VDD1.n1 VDD1.n0 71.9653
R155 VDD1.n3 VDD1.n2 71.9643
R156 VDD1.n7 VDD1.n6 71.9642
R157 VDD1.n7 VDD1.n5 52.8177
R158 VDD1.n6 VDD1.t1 1.83694
R159 VDD1.n6 VDD1.t5 1.83694
R160 VDD1.n0 VDD1.t3 1.83694
R161 VDD1.n0 VDD1.t8 1.83694
R162 VDD1.n4 VDD1.t2 1.83694
R163 VDD1.n4 VDD1.t4 1.83694
R164 VDD1.n2 VDD1.t6 1.83694
R165 VDD1.n2 VDD1.t9 1.83694
R166 VDD1 VDD1.n7 1.83671
R167 VDD1 VDD1.n1 0.690155
R168 VDD1.n5 VDD1.n3 0.576619
R169 VTAIL.n11 VTAIL.t2 57.1229
R170 VTAIL.n17 VTAIL.t6 57.122
R171 VTAIL.n2 VTAIL.t10 57.122
R172 VTAIL.n16 VTAIL.t11 57.1218
R173 VTAIL.n15 VTAIL.n14 55.2865
R174 VTAIL.n13 VTAIL.n12 55.2865
R175 VTAIL.n10 VTAIL.n9 55.2865
R176 VTAIL.n8 VTAIL.n7 55.2865
R177 VTAIL.n19 VTAIL.n18 55.2855
R178 VTAIL.n1 VTAIL.n0 55.2855
R179 VTAIL.n4 VTAIL.n3 55.2855
R180 VTAIL.n6 VTAIL.n5 55.2855
R181 VTAIL.n8 VTAIL.n6 32.6772
R182 VTAIL.n17 VTAIL.n16 30.1514
R183 VTAIL.n10 VTAIL.n8 2.52636
R184 VTAIL.n11 VTAIL.n10 2.52636
R185 VTAIL.n15 VTAIL.n13 2.52636
R186 VTAIL.n16 VTAIL.n15 2.52636
R187 VTAIL.n6 VTAIL.n4 2.52636
R188 VTAIL.n4 VTAIL.n2 2.52636
R189 VTAIL.n19 VTAIL.n17 2.52636
R190 VTAIL VTAIL.n1 1.95309
R191 VTAIL.n18 VTAIL.t3 1.83694
R192 VTAIL.n18 VTAIL.t0 1.83694
R193 VTAIL.n0 VTAIL.t5 1.83694
R194 VTAIL.n0 VTAIL.t8 1.83694
R195 VTAIL.n3 VTAIL.t13 1.83694
R196 VTAIL.n3 VTAIL.t18 1.83694
R197 VTAIL.n5 VTAIL.t16 1.83694
R198 VTAIL.n5 VTAIL.t14 1.83694
R199 VTAIL.n14 VTAIL.t12 1.83694
R200 VTAIL.n14 VTAIL.t17 1.83694
R201 VTAIL.n12 VTAIL.t15 1.83694
R202 VTAIL.n12 VTAIL.t19 1.83694
R203 VTAIL.n9 VTAIL.t7 1.83694
R204 VTAIL.n9 VTAIL.t9 1.83694
R205 VTAIL.n7 VTAIL.t4 1.83694
R206 VTAIL.n7 VTAIL.t1 1.83694
R207 VTAIL.n13 VTAIL.n11 1.73326
R208 VTAIL.n2 VTAIL.n1 1.73326
R209 VTAIL VTAIL.n19 0.573776
R210 B.n718 B.n99 585
R211 B.n720 B.n719 585
R212 B.n721 B.n98 585
R213 B.n723 B.n722 585
R214 B.n724 B.n97 585
R215 B.n726 B.n725 585
R216 B.n727 B.n96 585
R217 B.n729 B.n728 585
R218 B.n730 B.n95 585
R219 B.n732 B.n731 585
R220 B.n733 B.n94 585
R221 B.n735 B.n734 585
R222 B.n736 B.n93 585
R223 B.n738 B.n737 585
R224 B.n739 B.n92 585
R225 B.n741 B.n740 585
R226 B.n742 B.n91 585
R227 B.n744 B.n743 585
R228 B.n745 B.n90 585
R229 B.n747 B.n746 585
R230 B.n748 B.n89 585
R231 B.n750 B.n749 585
R232 B.n751 B.n88 585
R233 B.n753 B.n752 585
R234 B.n754 B.n87 585
R235 B.n756 B.n755 585
R236 B.n757 B.n86 585
R237 B.n759 B.n758 585
R238 B.n760 B.n85 585
R239 B.n762 B.n761 585
R240 B.n763 B.n84 585
R241 B.n765 B.n764 585
R242 B.n766 B.n83 585
R243 B.n768 B.n767 585
R244 B.n769 B.n82 585
R245 B.n771 B.n770 585
R246 B.n772 B.n81 585
R247 B.n774 B.n773 585
R248 B.n775 B.n80 585
R249 B.n777 B.n776 585
R250 B.n778 B.n79 585
R251 B.n780 B.n779 585
R252 B.n781 B.n78 585
R253 B.n783 B.n782 585
R254 B.n784 B.n77 585
R255 B.n786 B.n785 585
R256 B.n787 B.n76 585
R257 B.n789 B.n788 585
R258 B.n790 B.n75 585
R259 B.n792 B.n791 585
R260 B.n793 B.n74 585
R261 B.n795 B.n794 585
R262 B.n796 B.n73 585
R263 B.n798 B.n797 585
R264 B.n799 B.n72 585
R265 B.n801 B.n800 585
R266 B.n802 B.n71 585
R267 B.n804 B.n803 585
R268 B.n806 B.n805 585
R269 B.n807 B.n67 585
R270 B.n809 B.n808 585
R271 B.n810 B.n66 585
R272 B.n812 B.n811 585
R273 B.n813 B.n65 585
R274 B.n815 B.n814 585
R275 B.n816 B.n64 585
R276 B.n818 B.n817 585
R277 B.n819 B.n61 585
R278 B.n822 B.n821 585
R279 B.n823 B.n60 585
R280 B.n825 B.n824 585
R281 B.n826 B.n59 585
R282 B.n828 B.n827 585
R283 B.n829 B.n58 585
R284 B.n831 B.n830 585
R285 B.n832 B.n57 585
R286 B.n834 B.n833 585
R287 B.n835 B.n56 585
R288 B.n837 B.n836 585
R289 B.n838 B.n55 585
R290 B.n840 B.n839 585
R291 B.n841 B.n54 585
R292 B.n843 B.n842 585
R293 B.n844 B.n53 585
R294 B.n846 B.n845 585
R295 B.n847 B.n52 585
R296 B.n849 B.n848 585
R297 B.n850 B.n51 585
R298 B.n852 B.n851 585
R299 B.n853 B.n50 585
R300 B.n855 B.n854 585
R301 B.n856 B.n49 585
R302 B.n858 B.n857 585
R303 B.n859 B.n48 585
R304 B.n861 B.n860 585
R305 B.n862 B.n47 585
R306 B.n864 B.n863 585
R307 B.n865 B.n46 585
R308 B.n867 B.n866 585
R309 B.n868 B.n45 585
R310 B.n870 B.n869 585
R311 B.n871 B.n44 585
R312 B.n873 B.n872 585
R313 B.n874 B.n43 585
R314 B.n876 B.n875 585
R315 B.n877 B.n42 585
R316 B.n879 B.n878 585
R317 B.n880 B.n41 585
R318 B.n882 B.n881 585
R319 B.n883 B.n40 585
R320 B.n885 B.n884 585
R321 B.n886 B.n39 585
R322 B.n888 B.n887 585
R323 B.n889 B.n38 585
R324 B.n891 B.n890 585
R325 B.n892 B.n37 585
R326 B.n894 B.n893 585
R327 B.n895 B.n36 585
R328 B.n897 B.n896 585
R329 B.n898 B.n35 585
R330 B.n900 B.n899 585
R331 B.n901 B.n34 585
R332 B.n903 B.n902 585
R333 B.n904 B.n33 585
R334 B.n906 B.n905 585
R335 B.n907 B.n32 585
R336 B.n717 B.n716 585
R337 B.n715 B.n100 585
R338 B.n714 B.n713 585
R339 B.n712 B.n101 585
R340 B.n711 B.n710 585
R341 B.n709 B.n102 585
R342 B.n708 B.n707 585
R343 B.n706 B.n103 585
R344 B.n705 B.n704 585
R345 B.n703 B.n104 585
R346 B.n702 B.n701 585
R347 B.n700 B.n105 585
R348 B.n699 B.n698 585
R349 B.n697 B.n106 585
R350 B.n696 B.n695 585
R351 B.n694 B.n107 585
R352 B.n693 B.n692 585
R353 B.n691 B.n108 585
R354 B.n690 B.n689 585
R355 B.n688 B.n109 585
R356 B.n687 B.n686 585
R357 B.n685 B.n110 585
R358 B.n684 B.n683 585
R359 B.n682 B.n111 585
R360 B.n681 B.n680 585
R361 B.n679 B.n112 585
R362 B.n678 B.n677 585
R363 B.n676 B.n113 585
R364 B.n675 B.n674 585
R365 B.n673 B.n114 585
R366 B.n672 B.n671 585
R367 B.n670 B.n115 585
R368 B.n669 B.n668 585
R369 B.n667 B.n116 585
R370 B.n666 B.n665 585
R371 B.n664 B.n117 585
R372 B.n663 B.n662 585
R373 B.n661 B.n118 585
R374 B.n660 B.n659 585
R375 B.n658 B.n119 585
R376 B.n657 B.n656 585
R377 B.n655 B.n120 585
R378 B.n654 B.n653 585
R379 B.n652 B.n121 585
R380 B.n651 B.n650 585
R381 B.n649 B.n122 585
R382 B.n648 B.n647 585
R383 B.n646 B.n123 585
R384 B.n645 B.n644 585
R385 B.n643 B.n124 585
R386 B.n642 B.n641 585
R387 B.n640 B.n125 585
R388 B.n639 B.n638 585
R389 B.n637 B.n126 585
R390 B.n636 B.n635 585
R391 B.n634 B.n127 585
R392 B.n633 B.n632 585
R393 B.n631 B.n128 585
R394 B.n630 B.n629 585
R395 B.n628 B.n129 585
R396 B.n627 B.n626 585
R397 B.n625 B.n130 585
R398 B.n624 B.n623 585
R399 B.n622 B.n131 585
R400 B.n621 B.n620 585
R401 B.n619 B.n132 585
R402 B.n618 B.n617 585
R403 B.n616 B.n133 585
R404 B.n615 B.n614 585
R405 B.n613 B.n134 585
R406 B.n612 B.n611 585
R407 B.n610 B.n135 585
R408 B.n609 B.n608 585
R409 B.n607 B.n136 585
R410 B.n606 B.n605 585
R411 B.n604 B.n137 585
R412 B.n603 B.n602 585
R413 B.n601 B.n138 585
R414 B.n600 B.n599 585
R415 B.n598 B.n139 585
R416 B.n597 B.n596 585
R417 B.n595 B.n140 585
R418 B.n594 B.n593 585
R419 B.n592 B.n141 585
R420 B.n591 B.n590 585
R421 B.n589 B.n142 585
R422 B.n588 B.n587 585
R423 B.n586 B.n143 585
R424 B.n585 B.n584 585
R425 B.n583 B.n144 585
R426 B.n582 B.n581 585
R427 B.n580 B.n145 585
R428 B.n579 B.n578 585
R429 B.n577 B.n146 585
R430 B.n576 B.n575 585
R431 B.n574 B.n147 585
R432 B.n573 B.n572 585
R433 B.n571 B.n148 585
R434 B.n570 B.n569 585
R435 B.n568 B.n149 585
R436 B.n567 B.n566 585
R437 B.n565 B.n150 585
R438 B.n564 B.n563 585
R439 B.n562 B.n151 585
R440 B.n561 B.n560 585
R441 B.n559 B.n152 585
R442 B.n558 B.n557 585
R443 B.n556 B.n153 585
R444 B.n555 B.n554 585
R445 B.n553 B.n154 585
R446 B.n552 B.n551 585
R447 B.n550 B.n155 585
R448 B.n549 B.n548 585
R449 B.n547 B.n156 585
R450 B.n546 B.n545 585
R451 B.n544 B.n157 585
R452 B.n543 B.n542 585
R453 B.n541 B.n158 585
R454 B.n540 B.n539 585
R455 B.n538 B.n159 585
R456 B.n537 B.n536 585
R457 B.n346 B.n227 585
R458 B.n348 B.n347 585
R459 B.n349 B.n226 585
R460 B.n351 B.n350 585
R461 B.n352 B.n225 585
R462 B.n354 B.n353 585
R463 B.n355 B.n224 585
R464 B.n357 B.n356 585
R465 B.n358 B.n223 585
R466 B.n360 B.n359 585
R467 B.n361 B.n222 585
R468 B.n363 B.n362 585
R469 B.n364 B.n221 585
R470 B.n366 B.n365 585
R471 B.n367 B.n220 585
R472 B.n369 B.n368 585
R473 B.n370 B.n219 585
R474 B.n372 B.n371 585
R475 B.n373 B.n218 585
R476 B.n375 B.n374 585
R477 B.n376 B.n217 585
R478 B.n378 B.n377 585
R479 B.n379 B.n216 585
R480 B.n381 B.n380 585
R481 B.n382 B.n215 585
R482 B.n384 B.n383 585
R483 B.n385 B.n214 585
R484 B.n387 B.n386 585
R485 B.n388 B.n213 585
R486 B.n390 B.n389 585
R487 B.n391 B.n212 585
R488 B.n393 B.n392 585
R489 B.n394 B.n211 585
R490 B.n396 B.n395 585
R491 B.n397 B.n210 585
R492 B.n399 B.n398 585
R493 B.n400 B.n209 585
R494 B.n402 B.n401 585
R495 B.n403 B.n208 585
R496 B.n405 B.n404 585
R497 B.n406 B.n207 585
R498 B.n408 B.n407 585
R499 B.n409 B.n206 585
R500 B.n411 B.n410 585
R501 B.n412 B.n205 585
R502 B.n414 B.n413 585
R503 B.n415 B.n204 585
R504 B.n417 B.n416 585
R505 B.n418 B.n203 585
R506 B.n420 B.n419 585
R507 B.n421 B.n202 585
R508 B.n423 B.n422 585
R509 B.n424 B.n201 585
R510 B.n426 B.n425 585
R511 B.n427 B.n200 585
R512 B.n429 B.n428 585
R513 B.n430 B.n199 585
R514 B.n432 B.n431 585
R515 B.n434 B.n433 585
R516 B.n435 B.n195 585
R517 B.n437 B.n436 585
R518 B.n438 B.n194 585
R519 B.n440 B.n439 585
R520 B.n441 B.n193 585
R521 B.n443 B.n442 585
R522 B.n444 B.n192 585
R523 B.n446 B.n445 585
R524 B.n447 B.n189 585
R525 B.n450 B.n449 585
R526 B.n451 B.n188 585
R527 B.n453 B.n452 585
R528 B.n454 B.n187 585
R529 B.n456 B.n455 585
R530 B.n457 B.n186 585
R531 B.n459 B.n458 585
R532 B.n460 B.n185 585
R533 B.n462 B.n461 585
R534 B.n463 B.n184 585
R535 B.n465 B.n464 585
R536 B.n466 B.n183 585
R537 B.n468 B.n467 585
R538 B.n469 B.n182 585
R539 B.n471 B.n470 585
R540 B.n472 B.n181 585
R541 B.n474 B.n473 585
R542 B.n475 B.n180 585
R543 B.n477 B.n476 585
R544 B.n478 B.n179 585
R545 B.n480 B.n479 585
R546 B.n481 B.n178 585
R547 B.n483 B.n482 585
R548 B.n484 B.n177 585
R549 B.n486 B.n485 585
R550 B.n487 B.n176 585
R551 B.n489 B.n488 585
R552 B.n490 B.n175 585
R553 B.n492 B.n491 585
R554 B.n493 B.n174 585
R555 B.n495 B.n494 585
R556 B.n496 B.n173 585
R557 B.n498 B.n497 585
R558 B.n499 B.n172 585
R559 B.n501 B.n500 585
R560 B.n502 B.n171 585
R561 B.n504 B.n503 585
R562 B.n505 B.n170 585
R563 B.n507 B.n506 585
R564 B.n508 B.n169 585
R565 B.n510 B.n509 585
R566 B.n511 B.n168 585
R567 B.n513 B.n512 585
R568 B.n514 B.n167 585
R569 B.n516 B.n515 585
R570 B.n517 B.n166 585
R571 B.n519 B.n518 585
R572 B.n520 B.n165 585
R573 B.n522 B.n521 585
R574 B.n523 B.n164 585
R575 B.n525 B.n524 585
R576 B.n526 B.n163 585
R577 B.n528 B.n527 585
R578 B.n529 B.n162 585
R579 B.n531 B.n530 585
R580 B.n532 B.n161 585
R581 B.n534 B.n533 585
R582 B.n535 B.n160 585
R583 B.n345 B.n344 585
R584 B.n343 B.n228 585
R585 B.n342 B.n341 585
R586 B.n340 B.n229 585
R587 B.n339 B.n338 585
R588 B.n337 B.n230 585
R589 B.n336 B.n335 585
R590 B.n334 B.n231 585
R591 B.n333 B.n332 585
R592 B.n331 B.n232 585
R593 B.n330 B.n329 585
R594 B.n328 B.n233 585
R595 B.n327 B.n326 585
R596 B.n325 B.n234 585
R597 B.n324 B.n323 585
R598 B.n322 B.n235 585
R599 B.n321 B.n320 585
R600 B.n319 B.n236 585
R601 B.n318 B.n317 585
R602 B.n316 B.n237 585
R603 B.n315 B.n314 585
R604 B.n313 B.n238 585
R605 B.n312 B.n311 585
R606 B.n310 B.n239 585
R607 B.n309 B.n308 585
R608 B.n307 B.n240 585
R609 B.n306 B.n305 585
R610 B.n304 B.n241 585
R611 B.n303 B.n302 585
R612 B.n301 B.n242 585
R613 B.n300 B.n299 585
R614 B.n298 B.n243 585
R615 B.n297 B.n296 585
R616 B.n295 B.n244 585
R617 B.n294 B.n293 585
R618 B.n292 B.n245 585
R619 B.n291 B.n290 585
R620 B.n289 B.n246 585
R621 B.n288 B.n287 585
R622 B.n286 B.n247 585
R623 B.n285 B.n284 585
R624 B.n283 B.n248 585
R625 B.n282 B.n281 585
R626 B.n280 B.n249 585
R627 B.n279 B.n278 585
R628 B.n277 B.n250 585
R629 B.n276 B.n275 585
R630 B.n274 B.n251 585
R631 B.n273 B.n272 585
R632 B.n271 B.n252 585
R633 B.n270 B.n269 585
R634 B.n268 B.n253 585
R635 B.n267 B.n266 585
R636 B.n265 B.n254 585
R637 B.n264 B.n263 585
R638 B.n262 B.n255 585
R639 B.n261 B.n260 585
R640 B.n259 B.n256 585
R641 B.n258 B.n257 585
R642 B.n2 B.n0 585
R643 B.n997 B.n1 585
R644 B.n996 B.n995 585
R645 B.n994 B.n3 585
R646 B.n993 B.n992 585
R647 B.n991 B.n4 585
R648 B.n990 B.n989 585
R649 B.n988 B.n5 585
R650 B.n987 B.n986 585
R651 B.n985 B.n6 585
R652 B.n984 B.n983 585
R653 B.n982 B.n7 585
R654 B.n981 B.n980 585
R655 B.n979 B.n8 585
R656 B.n978 B.n977 585
R657 B.n976 B.n9 585
R658 B.n975 B.n974 585
R659 B.n973 B.n10 585
R660 B.n972 B.n971 585
R661 B.n970 B.n11 585
R662 B.n969 B.n968 585
R663 B.n967 B.n12 585
R664 B.n966 B.n965 585
R665 B.n964 B.n13 585
R666 B.n963 B.n962 585
R667 B.n961 B.n14 585
R668 B.n960 B.n959 585
R669 B.n958 B.n15 585
R670 B.n957 B.n956 585
R671 B.n955 B.n16 585
R672 B.n954 B.n953 585
R673 B.n952 B.n17 585
R674 B.n951 B.n950 585
R675 B.n949 B.n18 585
R676 B.n948 B.n947 585
R677 B.n946 B.n19 585
R678 B.n945 B.n944 585
R679 B.n943 B.n20 585
R680 B.n942 B.n941 585
R681 B.n940 B.n21 585
R682 B.n939 B.n938 585
R683 B.n937 B.n22 585
R684 B.n936 B.n935 585
R685 B.n934 B.n23 585
R686 B.n933 B.n932 585
R687 B.n931 B.n24 585
R688 B.n930 B.n929 585
R689 B.n928 B.n25 585
R690 B.n927 B.n926 585
R691 B.n925 B.n26 585
R692 B.n924 B.n923 585
R693 B.n922 B.n27 585
R694 B.n921 B.n920 585
R695 B.n919 B.n28 585
R696 B.n918 B.n917 585
R697 B.n916 B.n29 585
R698 B.n915 B.n914 585
R699 B.n913 B.n30 585
R700 B.n912 B.n911 585
R701 B.n910 B.n31 585
R702 B.n909 B.n908 585
R703 B.n999 B.n998 585
R704 B.n344 B.n227 497.305
R705 B.n908 B.n907 497.305
R706 B.n536 B.n535 497.305
R707 B.n716 B.n99 497.305
R708 B.n190 B.t9 372.113
R709 B.n196 B.t6 372.113
R710 B.n62 B.t0 372.113
R711 B.n68 B.t3 372.113
R712 B.n190 B.t11 163.446
R713 B.n68 B.t4 163.446
R714 B.n196 B.t8 163.423
R715 B.n62 B.t1 163.423
R716 B.n344 B.n343 163.367
R717 B.n343 B.n342 163.367
R718 B.n342 B.n229 163.367
R719 B.n338 B.n229 163.367
R720 B.n338 B.n337 163.367
R721 B.n337 B.n336 163.367
R722 B.n336 B.n231 163.367
R723 B.n332 B.n231 163.367
R724 B.n332 B.n331 163.367
R725 B.n331 B.n330 163.367
R726 B.n330 B.n233 163.367
R727 B.n326 B.n233 163.367
R728 B.n326 B.n325 163.367
R729 B.n325 B.n324 163.367
R730 B.n324 B.n235 163.367
R731 B.n320 B.n235 163.367
R732 B.n320 B.n319 163.367
R733 B.n319 B.n318 163.367
R734 B.n318 B.n237 163.367
R735 B.n314 B.n237 163.367
R736 B.n314 B.n313 163.367
R737 B.n313 B.n312 163.367
R738 B.n312 B.n239 163.367
R739 B.n308 B.n239 163.367
R740 B.n308 B.n307 163.367
R741 B.n307 B.n306 163.367
R742 B.n306 B.n241 163.367
R743 B.n302 B.n241 163.367
R744 B.n302 B.n301 163.367
R745 B.n301 B.n300 163.367
R746 B.n300 B.n243 163.367
R747 B.n296 B.n243 163.367
R748 B.n296 B.n295 163.367
R749 B.n295 B.n294 163.367
R750 B.n294 B.n245 163.367
R751 B.n290 B.n245 163.367
R752 B.n290 B.n289 163.367
R753 B.n289 B.n288 163.367
R754 B.n288 B.n247 163.367
R755 B.n284 B.n247 163.367
R756 B.n284 B.n283 163.367
R757 B.n283 B.n282 163.367
R758 B.n282 B.n249 163.367
R759 B.n278 B.n249 163.367
R760 B.n278 B.n277 163.367
R761 B.n277 B.n276 163.367
R762 B.n276 B.n251 163.367
R763 B.n272 B.n251 163.367
R764 B.n272 B.n271 163.367
R765 B.n271 B.n270 163.367
R766 B.n270 B.n253 163.367
R767 B.n266 B.n253 163.367
R768 B.n266 B.n265 163.367
R769 B.n265 B.n264 163.367
R770 B.n264 B.n255 163.367
R771 B.n260 B.n255 163.367
R772 B.n260 B.n259 163.367
R773 B.n259 B.n258 163.367
R774 B.n258 B.n2 163.367
R775 B.n998 B.n2 163.367
R776 B.n998 B.n997 163.367
R777 B.n997 B.n996 163.367
R778 B.n996 B.n3 163.367
R779 B.n992 B.n3 163.367
R780 B.n992 B.n991 163.367
R781 B.n991 B.n990 163.367
R782 B.n990 B.n5 163.367
R783 B.n986 B.n5 163.367
R784 B.n986 B.n985 163.367
R785 B.n985 B.n984 163.367
R786 B.n984 B.n7 163.367
R787 B.n980 B.n7 163.367
R788 B.n980 B.n979 163.367
R789 B.n979 B.n978 163.367
R790 B.n978 B.n9 163.367
R791 B.n974 B.n9 163.367
R792 B.n974 B.n973 163.367
R793 B.n973 B.n972 163.367
R794 B.n972 B.n11 163.367
R795 B.n968 B.n11 163.367
R796 B.n968 B.n967 163.367
R797 B.n967 B.n966 163.367
R798 B.n966 B.n13 163.367
R799 B.n962 B.n13 163.367
R800 B.n962 B.n961 163.367
R801 B.n961 B.n960 163.367
R802 B.n960 B.n15 163.367
R803 B.n956 B.n15 163.367
R804 B.n956 B.n955 163.367
R805 B.n955 B.n954 163.367
R806 B.n954 B.n17 163.367
R807 B.n950 B.n17 163.367
R808 B.n950 B.n949 163.367
R809 B.n949 B.n948 163.367
R810 B.n948 B.n19 163.367
R811 B.n944 B.n19 163.367
R812 B.n944 B.n943 163.367
R813 B.n943 B.n942 163.367
R814 B.n942 B.n21 163.367
R815 B.n938 B.n21 163.367
R816 B.n938 B.n937 163.367
R817 B.n937 B.n936 163.367
R818 B.n936 B.n23 163.367
R819 B.n932 B.n23 163.367
R820 B.n932 B.n931 163.367
R821 B.n931 B.n930 163.367
R822 B.n930 B.n25 163.367
R823 B.n926 B.n25 163.367
R824 B.n926 B.n925 163.367
R825 B.n925 B.n924 163.367
R826 B.n924 B.n27 163.367
R827 B.n920 B.n27 163.367
R828 B.n920 B.n919 163.367
R829 B.n919 B.n918 163.367
R830 B.n918 B.n29 163.367
R831 B.n914 B.n29 163.367
R832 B.n914 B.n913 163.367
R833 B.n913 B.n912 163.367
R834 B.n912 B.n31 163.367
R835 B.n908 B.n31 163.367
R836 B.n348 B.n227 163.367
R837 B.n349 B.n348 163.367
R838 B.n350 B.n349 163.367
R839 B.n350 B.n225 163.367
R840 B.n354 B.n225 163.367
R841 B.n355 B.n354 163.367
R842 B.n356 B.n355 163.367
R843 B.n356 B.n223 163.367
R844 B.n360 B.n223 163.367
R845 B.n361 B.n360 163.367
R846 B.n362 B.n361 163.367
R847 B.n362 B.n221 163.367
R848 B.n366 B.n221 163.367
R849 B.n367 B.n366 163.367
R850 B.n368 B.n367 163.367
R851 B.n368 B.n219 163.367
R852 B.n372 B.n219 163.367
R853 B.n373 B.n372 163.367
R854 B.n374 B.n373 163.367
R855 B.n374 B.n217 163.367
R856 B.n378 B.n217 163.367
R857 B.n379 B.n378 163.367
R858 B.n380 B.n379 163.367
R859 B.n380 B.n215 163.367
R860 B.n384 B.n215 163.367
R861 B.n385 B.n384 163.367
R862 B.n386 B.n385 163.367
R863 B.n386 B.n213 163.367
R864 B.n390 B.n213 163.367
R865 B.n391 B.n390 163.367
R866 B.n392 B.n391 163.367
R867 B.n392 B.n211 163.367
R868 B.n396 B.n211 163.367
R869 B.n397 B.n396 163.367
R870 B.n398 B.n397 163.367
R871 B.n398 B.n209 163.367
R872 B.n402 B.n209 163.367
R873 B.n403 B.n402 163.367
R874 B.n404 B.n403 163.367
R875 B.n404 B.n207 163.367
R876 B.n408 B.n207 163.367
R877 B.n409 B.n408 163.367
R878 B.n410 B.n409 163.367
R879 B.n410 B.n205 163.367
R880 B.n414 B.n205 163.367
R881 B.n415 B.n414 163.367
R882 B.n416 B.n415 163.367
R883 B.n416 B.n203 163.367
R884 B.n420 B.n203 163.367
R885 B.n421 B.n420 163.367
R886 B.n422 B.n421 163.367
R887 B.n422 B.n201 163.367
R888 B.n426 B.n201 163.367
R889 B.n427 B.n426 163.367
R890 B.n428 B.n427 163.367
R891 B.n428 B.n199 163.367
R892 B.n432 B.n199 163.367
R893 B.n433 B.n432 163.367
R894 B.n433 B.n195 163.367
R895 B.n437 B.n195 163.367
R896 B.n438 B.n437 163.367
R897 B.n439 B.n438 163.367
R898 B.n439 B.n193 163.367
R899 B.n443 B.n193 163.367
R900 B.n444 B.n443 163.367
R901 B.n445 B.n444 163.367
R902 B.n445 B.n189 163.367
R903 B.n450 B.n189 163.367
R904 B.n451 B.n450 163.367
R905 B.n452 B.n451 163.367
R906 B.n452 B.n187 163.367
R907 B.n456 B.n187 163.367
R908 B.n457 B.n456 163.367
R909 B.n458 B.n457 163.367
R910 B.n458 B.n185 163.367
R911 B.n462 B.n185 163.367
R912 B.n463 B.n462 163.367
R913 B.n464 B.n463 163.367
R914 B.n464 B.n183 163.367
R915 B.n468 B.n183 163.367
R916 B.n469 B.n468 163.367
R917 B.n470 B.n469 163.367
R918 B.n470 B.n181 163.367
R919 B.n474 B.n181 163.367
R920 B.n475 B.n474 163.367
R921 B.n476 B.n475 163.367
R922 B.n476 B.n179 163.367
R923 B.n480 B.n179 163.367
R924 B.n481 B.n480 163.367
R925 B.n482 B.n481 163.367
R926 B.n482 B.n177 163.367
R927 B.n486 B.n177 163.367
R928 B.n487 B.n486 163.367
R929 B.n488 B.n487 163.367
R930 B.n488 B.n175 163.367
R931 B.n492 B.n175 163.367
R932 B.n493 B.n492 163.367
R933 B.n494 B.n493 163.367
R934 B.n494 B.n173 163.367
R935 B.n498 B.n173 163.367
R936 B.n499 B.n498 163.367
R937 B.n500 B.n499 163.367
R938 B.n500 B.n171 163.367
R939 B.n504 B.n171 163.367
R940 B.n505 B.n504 163.367
R941 B.n506 B.n505 163.367
R942 B.n506 B.n169 163.367
R943 B.n510 B.n169 163.367
R944 B.n511 B.n510 163.367
R945 B.n512 B.n511 163.367
R946 B.n512 B.n167 163.367
R947 B.n516 B.n167 163.367
R948 B.n517 B.n516 163.367
R949 B.n518 B.n517 163.367
R950 B.n518 B.n165 163.367
R951 B.n522 B.n165 163.367
R952 B.n523 B.n522 163.367
R953 B.n524 B.n523 163.367
R954 B.n524 B.n163 163.367
R955 B.n528 B.n163 163.367
R956 B.n529 B.n528 163.367
R957 B.n530 B.n529 163.367
R958 B.n530 B.n161 163.367
R959 B.n534 B.n161 163.367
R960 B.n535 B.n534 163.367
R961 B.n536 B.n159 163.367
R962 B.n540 B.n159 163.367
R963 B.n541 B.n540 163.367
R964 B.n542 B.n541 163.367
R965 B.n542 B.n157 163.367
R966 B.n546 B.n157 163.367
R967 B.n547 B.n546 163.367
R968 B.n548 B.n547 163.367
R969 B.n548 B.n155 163.367
R970 B.n552 B.n155 163.367
R971 B.n553 B.n552 163.367
R972 B.n554 B.n553 163.367
R973 B.n554 B.n153 163.367
R974 B.n558 B.n153 163.367
R975 B.n559 B.n558 163.367
R976 B.n560 B.n559 163.367
R977 B.n560 B.n151 163.367
R978 B.n564 B.n151 163.367
R979 B.n565 B.n564 163.367
R980 B.n566 B.n565 163.367
R981 B.n566 B.n149 163.367
R982 B.n570 B.n149 163.367
R983 B.n571 B.n570 163.367
R984 B.n572 B.n571 163.367
R985 B.n572 B.n147 163.367
R986 B.n576 B.n147 163.367
R987 B.n577 B.n576 163.367
R988 B.n578 B.n577 163.367
R989 B.n578 B.n145 163.367
R990 B.n582 B.n145 163.367
R991 B.n583 B.n582 163.367
R992 B.n584 B.n583 163.367
R993 B.n584 B.n143 163.367
R994 B.n588 B.n143 163.367
R995 B.n589 B.n588 163.367
R996 B.n590 B.n589 163.367
R997 B.n590 B.n141 163.367
R998 B.n594 B.n141 163.367
R999 B.n595 B.n594 163.367
R1000 B.n596 B.n595 163.367
R1001 B.n596 B.n139 163.367
R1002 B.n600 B.n139 163.367
R1003 B.n601 B.n600 163.367
R1004 B.n602 B.n601 163.367
R1005 B.n602 B.n137 163.367
R1006 B.n606 B.n137 163.367
R1007 B.n607 B.n606 163.367
R1008 B.n608 B.n607 163.367
R1009 B.n608 B.n135 163.367
R1010 B.n612 B.n135 163.367
R1011 B.n613 B.n612 163.367
R1012 B.n614 B.n613 163.367
R1013 B.n614 B.n133 163.367
R1014 B.n618 B.n133 163.367
R1015 B.n619 B.n618 163.367
R1016 B.n620 B.n619 163.367
R1017 B.n620 B.n131 163.367
R1018 B.n624 B.n131 163.367
R1019 B.n625 B.n624 163.367
R1020 B.n626 B.n625 163.367
R1021 B.n626 B.n129 163.367
R1022 B.n630 B.n129 163.367
R1023 B.n631 B.n630 163.367
R1024 B.n632 B.n631 163.367
R1025 B.n632 B.n127 163.367
R1026 B.n636 B.n127 163.367
R1027 B.n637 B.n636 163.367
R1028 B.n638 B.n637 163.367
R1029 B.n638 B.n125 163.367
R1030 B.n642 B.n125 163.367
R1031 B.n643 B.n642 163.367
R1032 B.n644 B.n643 163.367
R1033 B.n644 B.n123 163.367
R1034 B.n648 B.n123 163.367
R1035 B.n649 B.n648 163.367
R1036 B.n650 B.n649 163.367
R1037 B.n650 B.n121 163.367
R1038 B.n654 B.n121 163.367
R1039 B.n655 B.n654 163.367
R1040 B.n656 B.n655 163.367
R1041 B.n656 B.n119 163.367
R1042 B.n660 B.n119 163.367
R1043 B.n661 B.n660 163.367
R1044 B.n662 B.n661 163.367
R1045 B.n662 B.n117 163.367
R1046 B.n666 B.n117 163.367
R1047 B.n667 B.n666 163.367
R1048 B.n668 B.n667 163.367
R1049 B.n668 B.n115 163.367
R1050 B.n672 B.n115 163.367
R1051 B.n673 B.n672 163.367
R1052 B.n674 B.n673 163.367
R1053 B.n674 B.n113 163.367
R1054 B.n678 B.n113 163.367
R1055 B.n679 B.n678 163.367
R1056 B.n680 B.n679 163.367
R1057 B.n680 B.n111 163.367
R1058 B.n684 B.n111 163.367
R1059 B.n685 B.n684 163.367
R1060 B.n686 B.n685 163.367
R1061 B.n686 B.n109 163.367
R1062 B.n690 B.n109 163.367
R1063 B.n691 B.n690 163.367
R1064 B.n692 B.n691 163.367
R1065 B.n692 B.n107 163.367
R1066 B.n696 B.n107 163.367
R1067 B.n697 B.n696 163.367
R1068 B.n698 B.n697 163.367
R1069 B.n698 B.n105 163.367
R1070 B.n702 B.n105 163.367
R1071 B.n703 B.n702 163.367
R1072 B.n704 B.n703 163.367
R1073 B.n704 B.n103 163.367
R1074 B.n708 B.n103 163.367
R1075 B.n709 B.n708 163.367
R1076 B.n710 B.n709 163.367
R1077 B.n710 B.n101 163.367
R1078 B.n714 B.n101 163.367
R1079 B.n715 B.n714 163.367
R1080 B.n716 B.n715 163.367
R1081 B.n907 B.n906 163.367
R1082 B.n906 B.n33 163.367
R1083 B.n902 B.n33 163.367
R1084 B.n902 B.n901 163.367
R1085 B.n901 B.n900 163.367
R1086 B.n900 B.n35 163.367
R1087 B.n896 B.n35 163.367
R1088 B.n896 B.n895 163.367
R1089 B.n895 B.n894 163.367
R1090 B.n894 B.n37 163.367
R1091 B.n890 B.n37 163.367
R1092 B.n890 B.n889 163.367
R1093 B.n889 B.n888 163.367
R1094 B.n888 B.n39 163.367
R1095 B.n884 B.n39 163.367
R1096 B.n884 B.n883 163.367
R1097 B.n883 B.n882 163.367
R1098 B.n882 B.n41 163.367
R1099 B.n878 B.n41 163.367
R1100 B.n878 B.n877 163.367
R1101 B.n877 B.n876 163.367
R1102 B.n876 B.n43 163.367
R1103 B.n872 B.n43 163.367
R1104 B.n872 B.n871 163.367
R1105 B.n871 B.n870 163.367
R1106 B.n870 B.n45 163.367
R1107 B.n866 B.n45 163.367
R1108 B.n866 B.n865 163.367
R1109 B.n865 B.n864 163.367
R1110 B.n864 B.n47 163.367
R1111 B.n860 B.n47 163.367
R1112 B.n860 B.n859 163.367
R1113 B.n859 B.n858 163.367
R1114 B.n858 B.n49 163.367
R1115 B.n854 B.n49 163.367
R1116 B.n854 B.n853 163.367
R1117 B.n853 B.n852 163.367
R1118 B.n852 B.n51 163.367
R1119 B.n848 B.n51 163.367
R1120 B.n848 B.n847 163.367
R1121 B.n847 B.n846 163.367
R1122 B.n846 B.n53 163.367
R1123 B.n842 B.n53 163.367
R1124 B.n842 B.n841 163.367
R1125 B.n841 B.n840 163.367
R1126 B.n840 B.n55 163.367
R1127 B.n836 B.n55 163.367
R1128 B.n836 B.n835 163.367
R1129 B.n835 B.n834 163.367
R1130 B.n834 B.n57 163.367
R1131 B.n830 B.n57 163.367
R1132 B.n830 B.n829 163.367
R1133 B.n829 B.n828 163.367
R1134 B.n828 B.n59 163.367
R1135 B.n824 B.n59 163.367
R1136 B.n824 B.n823 163.367
R1137 B.n823 B.n822 163.367
R1138 B.n822 B.n61 163.367
R1139 B.n817 B.n61 163.367
R1140 B.n817 B.n816 163.367
R1141 B.n816 B.n815 163.367
R1142 B.n815 B.n65 163.367
R1143 B.n811 B.n65 163.367
R1144 B.n811 B.n810 163.367
R1145 B.n810 B.n809 163.367
R1146 B.n809 B.n67 163.367
R1147 B.n805 B.n67 163.367
R1148 B.n805 B.n804 163.367
R1149 B.n804 B.n71 163.367
R1150 B.n800 B.n71 163.367
R1151 B.n800 B.n799 163.367
R1152 B.n799 B.n798 163.367
R1153 B.n798 B.n73 163.367
R1154 B.n794 B.n73 163.367
R1155 B.n794 B.n793 163.367
R1156 B.n793 B.n792 163.367
R1157 B.n792 B.n75 163.367
R1158 B.n788 B.n75 163.367
R1159 B.n788 B.n787 163.367
R1160 B.n787 B.n786 163.367
R1161 B.n786 B.n77 163.367
R1162 B.n782 B.n77 163.367
R1163 B.n782 B.n781 163.367
R1164 B.n781 B.n780 163.367
R1165 B.n780 B.n79 163.367
R1166 B.n776 B.n79 163.367
R1167 B.n776 B.n775 163.367
R1168 B.n775 B.n774 163.367
R1169 B.n774 B.n81 163.367
R1170 B.n770 B.n81 163.367
R1171 B.n770 B.n769 163.367
R1172 B.n769 B.n768 163.367
R1173 B.n768 B.n83 163.367
R1174 B.n764 B.n83 163.367
R1175 B.n764 B.n763 163.367
R1176 B.n763 B.n762 163.367
R1177 B.n762 B.n85 163.367
R1178 B.n758 B.n85 163.367
R1179 B.n758 B.n757 163.367
R1180 B.n757 B.n756 163.367
R1181 B.n756 B.n87 163.367
R1182 B.n752 B.n87 163.367
R1183 B.n752 B.n751 163.367
R1184 B.n751 B.n750 163.367
R1185 B.n750 B.n89 163.367
R1186 B.n746 B.n89 163.367
R1187 B.n746 B.n745 163.367
R1188 B.n745 B.n744 163.367
R1189 B.n744 B.n91 163.367
R1190 B.n740 B.n91 163.367
R1191 B.n740 B.n739 163.367
R1192 B.n739 B.n738 163.367
R1193 B.n738 B.n93 163.367
R1194 B.n734 B.n93 163.367
R1195 B.n734 B.n733 163.367
R1196 B.n733 B.n732 163.367
R1197 B.n732 B.n95 163.367
R1198 B.n728 B.n95 163.367
R1199 B.n728 B.n727 163.367
R1200 B.n727 B.n726 163.367
R1201 B.n726 B.n97 163.367
R1202 B.n722 B.n97 163.367
R1203 B.n722 B.n721 163.367
R1204 B.n721 B.n720 163.367
R1205 B.n720 B.n99 163.367
R1206 B.n191 B.t10 106.623
R1207 B.n69 B.t5 106.623
R1208 B.n197 B.t7 106.6
R1209 B.n63 B.t2 106.6
R1210 B.n448 B.n191 59.5399
R1211 B.n198 B.n197 59.5399
R1212 B.n820 B.n63 59.5399
R1213 B.n70 B.n69 59.5399
R1214 B.n191 B.n190 56.8247
R1215 B.n197 B.n196 56.8247
R1216 B.n63 B.n62 56.8247
R1217 B.n69 B.n68 56.8247
R1218 B.n909 B.n32 32.3127
R1219 B.n718 B.n717 32.3127
R1220 B.n537 B.n160 32.3127
R1221 B.n346 B.n345 32.3127
R1222 B B.n999 18.0485
R1223 B.n905 B.n32 10.6151
R1224 B.n905 B.n904 10.6151
R1225 B.n904 B.n903 10.6151
R1226 B.n903 B.n34 10.6151
R1227 B.n899 B.n34 10.6151
R1228 B.n899 B.n898 10.6151
R1229 B.n898 B.n897 10.6151
R1230 B.n897 B.n36 10.6151
R1231 B.n893 B.n36 10.6151
R1232 B.n893 B.n892 10.6151
R1233 B.n892 B.n891 10.6151
R1234 B.n891 B.n38 10.6151
R1235 B.n887 B.n38 10.6151
R1236 B.n887 B.n886 10.6151
R1237 B.n886 B.n885 10.6151
R1238 B.n885 B.n40 10.6151
R1239 B.n881 B.n40 10.6151
R1240 B.n881 B.n880 10.6151
R1241 B.n880 B.n879 10.6151
R1242 B.n879 B.n42 10.6151
R1243 B.n875 B.n42 10.6151
R1244 B.n875 B.n874 10.6151
R1245 B.n874 B.n873 10.6151
R1246 B.n873 B.n44 10.6151
R1247 B.n869 B.n44 10.6151
R1248 B.n869 B.n868 10.6151
R1249 B.n868 B.n867 10.6151
R1250 B.n867 B.n46 10.6151
R1251 B.n863 B.n46 10.6151
R1252 B.n863 B.n862 10.6151
R1253 B.n862 B.n861 10.6151
R1254 B.n861 B.n48 10.6151
R1255 B.n857 B.n48 10.6151
R1256 B.n857 B.n856 10.6151
R1257 B.n856 B.n855 10.6151
R1258 B.n855 B.n50 10.6151
R1259 B.n851 B.n50 10.6151
R1260 B.n851 B.n850 10.6151
R1261 B.n850 B.n849 10.6151
R1262 B.n849 B.n52 10.6151
R1263 B.n845 B.n52 10.6151
R1264 B.n845 B.n844 10.6151
R1265 B.n844 B.n843 10.6151
R1266 B.n843 B.n54 10.6151
R1267 B.n839 B.n54 10.6151
R1268 B.n839 B.n838 10.6151
R1269 B.n838 B.n837 10.6151
R1270 B.n837 B.n56 10.6151
R1271 B.n833 B.n56 10.6151
R1272 B.n833 B.n832 10.6151
R1273 B.n832 B.n831 10.6151
R1274 B.n831 B.n58 10.6151
R1275 B.n827 B.n58 10.6151
R1276 B.n827 B.n826 10.6151
R1277 B.n826 B.n825 10.6151
R1278 B.n825 B.n60 10.6151
R1279 B.n821 B.n60 10.6151
R1280 B.n819 B.n818 10.6151
R1281 B.n818 B.n64 10.6151
R1282 B.n814 B.n64 10.6151
R1283 B.n814 B.n813 10.6151
R1284 B.n813 B.n812 10.6151
R1285 B.n812 B.n66 10.6151
R1286 B.n808 B.n66 10.6151
R1287 B.n808 B.n807 10.6151
R1288 B.n807 B.n806 10.6151
R1289 B.n803 B.n802 10.6151
R1290 B.n802 B.n801 10.6151
R1291 B.n801 B.n72 10.6151
R1292 B.n797 B.n72 10.6151
R1293 B.n797 B.n796 10.6151
R1294 B.n796 B.n795 10.6151
R1295 B.n795 B.n74 10.6151
R1296 B.n791 B.n74 10.6151
R1297 B.n791 B.n790 10.6151
R1298 B.n790 B.n789 10.6151
R1299 B.n789 B.n76 10.6151
R1300 B.n785 B.n76 10.6151
R1301 B.n785 B.n784 10.6151
R1302 B.n784 B.n783 10.6151
R1303 B.n783 B.n78 10.6151
R1304 B.n779 B.n78 10.6151
R1305 B.n779 B.n778 10.6151
R1306 B.n778 B.n777 10.6151
R1307 B.n777 B.n80 10.6151
R1308 B.n773 B.n80 10.6151
R1309 B.n773 B.n772 10.6151
R1310 B.n772 B.n771 10.6151
R1311 B.n771 B.n82 10.6151
R1312 B.n767 B.n82 10.6151
R1313 B.n767 B.n766 10.6151
R1314 B.n766 B.n765 10.6151
R1315 B.n765 B.n84 10.6151
R1316 B.n761 B.n84 10.6151
R1317 B.n761 B.n760 10.6151
R1318 B.n760 B.n759 10.6151
R1319 B.n759 B.n86 10.6151
R1320 B.n755 B.n86 10.6151
R1321 B.n755 B.n754 10.6151
R1322 B.n754 B.n753 10.6151
R1323 B.n753 B.n88 10.6151
R1324 B.n749 B.n88 10.6151
R1325 B.n749 B.n748 10.6151
R1326 B.n748 B.n747 10.6151
R1327 B.n747 B.n90 10.6151
R1328 B.n743 B.n90 10.6151
R1329 B.n743 B.n742 10.6151
R1330 B.n742 B.n741 10.6151
R1331 B.n741 B.n92 10.6151
R1332 B.n737 B.n92 10.6151
R1333 B.n737 B.n736 10.6151
R1334 B.n736 B.n735 10.6151
R1335 B.n735 B.n94 10.6151
R1336 B.n731 B.n94 10.6151
R1337 B.n731 B.n730 10.6151
R1338 B.n730 B.n729 10.6151
R1339 B.n729 B.n96 10.6151
R1340 B.n725 B.n96 10.6151
R1341 B.n725 B.n724 10.6151
R1342 B.n724 B.n723 10.6151
R1343 B.n723 B.n98 10.6151
R1344 B.n719 B.n98 10.6151
R1345 B.n719 B.n718 10.6151
R1346 B.n538 B.n537 10.6151
R1347 B.n539 B.n538 10.6151
R1348 B.n539 B.n158 10.6151
R1349 B.n543 B.n158 10.6151
R1350 B.n544 B.n543 10.6151
R1351 B.n545 B.n544 10.6151
R1352 B.n545 B.n156 10.6151
R1353 B.n549 B.n156 10.6151
R1354 B.n550 B.n549 10.6151
R1355 B.n551 B.n550 10.6151
R1356 B.n551 B.n154 10.6151
R1357 B.n555 B.n154 10.6151
R1358 B.n556 B.n555 10.6151
R1359 B.n557 B.n556 10.6151
R1360 B.n557 B.n152 10.6151
R1361 B.n561 B.n152 10.6151
R1362 B.n562 B.n561 10.6151
R1363 B.n563 B.n562 10.6151
R1364 B.n563 B.n150 10.6151
R1365 B.n567 B.n150 10.6151
R1366 B.n568 B.n567 10.6151
R1367 B.n569 B.n568 10.6151
R1368 B.n569 B.n148 10.6151
R1369 B.n573 B.n148 10.6151
R1370 B.n574 B.n573 10.6151
R1371 B.n575 B.n574 10.6151
R1372 B.n575 B.n146 10.6151
R1373 B.n579 B.n146 10.6151
R1374 B.n580 B.n579 10.6151
R1375 B.n581 B.n580 10.6151
R1376 B.n581 B.n144 10.6151
R1377 B.n585 B.n144 10.6151
R1378 B.n586 B.n585 10.6151
R1379 B.n587 B.n586 10.6151
R1380 B.n587 B.n142 10.6151
R1381 B.n591 B.n142 10.6151
R1382 B.n592 B.n591 10.6151
R1383 B.n593 B.n592 10.6151
R1384 B.n593 B.n140 10.6151
R1385 B.n597 B.n140 10.6151
R1386 B.n598 B.n597 10.6151
R1387 B.n599 B.n598 10.6151
R1388 B.n599 B.n138 10.6151
R1389 B.n603 B.n138 10.6151
R1390 B.n604 B.n603 10.6151
R1391 B.n605 B.n604 10.6151
R1392 B.n605 B.n136 10.6151
R1393 B.n609 B.n136 10.6151
R1394 B.n610 B.n609 10.6151
R1395 B.n611 B.n610 10.6151
R1396 B.n611 B.n134 10.6151
R1397 B.n615 B.n134 10.6151
R1398 B.n616 B.n615 10.6151
R1399 B.n617 B.n616 10.6151
R1400 B.n617 B.n132 10.6151
R1401 B.n621 B.n132 10.6151
R1402 B.n622 B.n621 10.6151
R1403 B.n623 B.n622 10.6151
R1404 B.n623 B.n130 10.6151
R1405 B.n627 B.n130 10.6151
R1406 B.n628 B.n627 10.6151
R1407 B.n629 B.n628 10.6151
R1408 B.n629 B.n128 10.6151
R1409 B.n633 B.n128 10.6151
R1410 B.n634 B.n633 10.6151
R1411 B.n635 B.n634 10.6151
R1412 B.n635 B.n126 10.6151
R1413 B.n639 B.n126 10.6151
R1414 B.n640 B.n639 10.6151
R1415 B.n641 B.n640 10.6151
R1416 B.n641 B.n124 10.6151
R1417 B.n645 B.n124 10.6151
R1418 B.n646 B.n645 10.6151
R1419 B.n647 B.n646 10.6151
R1420 B.n647 B.n122 10.6151
R1421 B.n651 B.n122 10.6151
R1422 B.n652 B.n651 10.6151
R1423 B.n653 B.n652 10.6151
R1424 B.n653 B.n120 10.6151
R1425 B.n657 B.n120 10.6151
R1426 B.n658 B.n657 10.6151
R1427 B.n659 B.n658 10.6151
R1428 B.n659 B.n118 10.6151
R1429 B.n663 B.n118 10.6151
R1430 B.n664 B.n663 10.6151
R1431 B.n665 B.n664 10.6151
R1432 B.n665 B.n116 10.6151
R1433 B.n669 B.n116 10.6151
R1434 B.n670 B.n669 10.6151
R1435 B.n671 B.n670 10.6151
R1436 B.n671 B.n114 10.6151
R1437 B.n675 B.n114 10.6151
R1438 B.n676 B.n675 10.6151
R1439 B.n677 B.n676 10.6151
R1440 B.n677 B.n112 10.6151
R1441 B.n681 B.n112 10.6151
R1442 B.n682 B.n681 10.6151
R1443 B.n683 B.n682 10.6151
R1444 B.n683 B.n110 10.6151
R1445 B.n687 B.n110 10.6151
R1446 B.n688 B.n687 10.6151
R1447 B.n689 B.n688 10.6151
R1448 B.n689 B.n108 10.6151
R1449 B.n693 B.n108 10.6151
R1450 B.n694 B.n693 10.6151
R1451 B.n695 B.n694 10.6151
R1452 B.n695 B.n106 10.6151
R1453 B.n699 B.n106 10.6151
R1454 B.n700 B.n699 10.6151
R1455 B.n701 B.n700 10.6151
R1456 B.n701 B.n104 10.6151
R1457 B.n705 B.n104 10.6151
R1458 B.n706 B.n705 10.6151
R1459 B.n707 B.n706 10.6151
R1460 B.n707 B.n102 10.6151
R1461 B.n711 B.n102 10.6151
R1462 B.n712 B.n711 10.6151
R1463 B.n713 B.n712 10.6151
R1464 B.n713 B.n100 10.6151
R1465 B.n717 B.n100 10.6151
R1466 B.n347 B.n346 10.6151
R1467 B.n347 B.n226 10.6151
R1468 B.n351 B.n226 10.6151
R1469 B.n352 B.n351 10.6151
R1470 B.n353 B.n352 10.6151
R1471 B.n353 B.n224 10.6151
R1472 B.n357 B.n224 10.6151
R1473 B.n358 B.n357 10.6151
R1474 B.n359 B.n358 10.6151
R1475 B.n359 B.n222 10.6151
R1476 B.n363 B.n222 10.6151
R1477 B.n364 B.n363 10.6151
R1478 B.n365 B.n364 10.6151
R1479 B.n365 B.n220 10.6151
R1480 B.n369 B.n220 10.6151
R1481 B.n370 B.n369 10.6151
R1482 B.n371 B.n370 10.6151
R1483 B.n371 B.n218 10.6151
R1484 B.n375 B.n218 10.6151
R1485 B.n376 B.n375 10.6151
R1486 B.n377 B.n376 10.6151
R1487 B.n377 B.n216 10.6151
R1488 B.n381 B.n216 10.6151
R1489 B.n382 B.n381 10.6151
R1490 B.n383 B.n382 10.6151
R1491 B.n383 B.n214 10.6151
R1492 B.n387 B.n214 10.6151
R1493 B.n388 B.n387 10.6151
R1494 B.n389 B.n388 10.6151
R1495 B.n389 B.n212 10.6151
R1496 B.n393 B.n212 10.6151
R1497 B.n394 B.n393 10.6151
R1498 B.n395 B.n394 10.6151
R1499 B.n395 B.n210 10.6151
R1500 B.n399 B.n210 10.6151
R1501 B.n400 B.n399 10.6151
R1502 B.n401 B.n400 10.6151
R1503 B.n401 B.n208 10.6151
R1504 B.n405 B.n208 10.6151
R1505 B.n406 B.n405 10.6151
R1506 B.n407 B.n406 10.6151
R1507 B.n407 B.n206 10.6151
R1508 B.n411 B.n206 10.6151
R1509 B.n412 B.n411 10.6151
R1510 B.n413 B.n412 10.6151
R1511 B.n413 B.n204 10.6151
R1512 B.n417 B.n204 10.6151
R1513 B.n418 B.n417 10.6151
R1514 B.n419 B.n418 10.6151
R1515 B.n419 B.n202 10.6151
R1516 B.n423 B.n202 10.6151
R1517 B.n424 B.n423 10.6151
R1518 B.n425 B.n424 10.6151
R1519 B.n425 B.n200 10.6151
R1520 B.n429 B.n200 10.6151
R1521 B.n430 B.n429 10.6151
R1522 B.n431 B.n430 10.6151
R1523 B.n435 B.n434 10.6151
R1524 B.n436 B.n435 10.6151
R1525 B.n436 B.n194 10.6151
R1526 B.n440 B.n194 10.6151
R1527 B.n441 B.n440 10.6151
R1528 B.n442 B.n441 10.6151
R1529 B.n442 B.n192 10.6151
R1530 B.n446 B.n192 10.6151
R1531 B.n447 B.n446 10.6151
R1532 B.n449 B.n188 10.6151
R1533 B.n453 B.n188 10.6151
R1534 B.n454 B.n453 10.6151
R1535 B.n455 B.n454 10.6151
R1536 B.n455 B.n186 10.6151
R1537 B.n459 B.n186 10.6151
R1538 B.n460 B.n459 10.6151
R1539 B.n461 B.n460 10.6151
R1540 B.n461 B.n184 10.6151
R1541 B.n465 B.n184 10.6151
R1542 B.n466 B.n465 10.6151
R1543 B.n467 B.n466 10.6151
R1544 B.n467 B.n182 10.6151
R1545 B.n471 B.n182 10.6151
R1546 B.n472 B.n471 10.6151
R1547 B.n473 B.n472 10.6151
R1548 B.n473 B.n180 10.6151
R1549 B.n477 B.n180 10.6151
R1550 B.n478 B.n477 10.6151
R1551 B.n479 B.n478 10.6151
R1552 B.n479 B.n178 10.6151
R1553 B.n483 B.n178 10.6151
R1554 B.n484 B.n483 10.6151
R1555 B.n485 B.n484 10.6151
R1556 B.n485 B.n176 10.6151
R1557 B.n489 B.n176 10.6151
R1558 B.n490 B.n489 10.6151
R1559 B.n491 B.n490 10.6151
R1560 B.n491 B.n174 10.6151
R1561 B.n495 B.n174 10.6151
R1562 B.n496 B.n495 10.6151
R1563 B.n497 B.n496 10.6151
R1564 B.n497 B.n172 10.6151
R1565 B.n501 B.n172 10.6151
R1566 B.n502 B.n501 10.6151
R1567 B.n503 B.n502 10.6151
R1568 B.n503 B.n170 10.6151
R1569 B.n507 B.n170 10.6151
R1570 B.n508 B.n507 10.6151
R1571 B.n509 B.n508 10.6151
R1572 B.n509 B.n168 10.6151
R1573 B.n513 B.n168 10.6151
R1574 B.n514 B.n513 10.6151
R1575 B.n515 B.n514 10.6151
R1576 B.n515 B.n166 10.6151
R1577 B.n519 B.n166 10.6151
R1578 B.n520 B.n519 10.6151
R1579 B.n521 B.n520 10.6151
R1580 B.n521 B.n164 10.6151
R1581 B.n525 B.n164 10.6151
R1582 B.n526 B.n525 10.6151
R1583 B.n527 B.n526 10.6151
R1584 B.n527 B.n162 10.6151
R1585 B.n531 B.n162 10.6151
R1586 B.n532 B.n531 10.6151
R1587 B.n533 B.n532 10.6151
R1588 B.n533 B.n160 10.6151
R1589 B.n345 B.n228 10.6151
R1590 B.n341 B.n228 10.6151
R1591 B.n341 B.n340 10.6151
R1592 B.n340 B.n339 10.6151
R1593 B.n339 B.n230 10.6151
R1594 B.n335 B.n230 10.6151
R1595 B.n335 B.n334 10.6151
R1596 B.n334 B.n333 10.6151
R1597 B.n333 B.n232 10.6151
R1598 B.n329 B.n232 10.6151
R1599 B.n329 B.n328 10.6151
R1600 B.n328 B.n327 10.6151
R1601 B.n327 B.n234 10.6151
R1602 B.n323 B.n234 10.6151
R1603 B.n323 B.n322 10.6151
R1604 B.n322 B.n321 10.6151
R1605 B.n321 B.n236 10.6151
R1606 B.n317 B.n236 10.6151
R1607 B.n317 B.n316 10.6151
R1608 B.n316 B.n315 10.6151
R1609 B.n315 B.n238 10.6151
R1610 B.n311 B.n238 10.6151
R1611 B.n311 B.n310 10.6151
R1612 B.n310 B.n309 10.6151
R1613 B.n309 B.n240 10.6151
R1614 B.n305 B.n240 10.6151
R1615 B.n305 B.n304 10.6151
R1616 B.n304 B.n303 10.6151
R1617 B.n303 B.n242 10.6151
R1618 B.n299 B.n242 10.6151
R1619 B.n299 B.n298 10.6151
R1620 B.n298 B.n297 10.6151
R1621 B.n297 B.n244 10.6151
R1622 B.n293 B.n244 10.6151
R1623 B.n293 B.n292 10.6151
R1624 B.n292 B.n291 10.6151
R1625 B.n291 B.n246 10.6151
R1626 B.n287 B.n246 10.6151
R1627 B.n287 B.n286 10.6151
R1628 B.n286 B.n285 10.6151
R1629 B.n285 B.n248 10.6151
R1630 B.n281 B.n248 10.6151
R1631 B.n281 B.n280 10.6151
R1632 B.n280 B.n279 10.6151
R1633 B.n279 B.n250 10.6151
R1634 B.n275 B.n250 10.6151
R1635 B.n275 B.n274 10.6151
R1636 B.n274 B.n273 10.6151
R1637 B.n273 B.n252 10.6151
R1638 B.n269 B.n252 10.6151
R1639 B.n269 B.n268 10.6151
R1640 B.n268 B.n267 10.6151
R1641 B.n267 B.n254 10.6151
R1642 B.n263 B.n254 10.6151
R1643 B.n263 B.n262 10.6151
R1644 B.n262 B.n261 10.6151
R1645 B.n261 B.n256 10.6151
R1646 B.n257 B.n256 10.6151
R1647 B.n257 B.n0 10.6151
R1648 B.n995 B.n1 10.6151
R1649 B.n995 B.n994 10.6151
R1650 B.n994 B.n993 10.6151
R1651 B.n993 B.n4 10.6151
R1652 B.n989 B.n4 10.6151
R1653 B.n989 B.n988 10.6151
R1654 B.n988 B.n987 10.6151
R1655 B.n987 B.n6 10.6151
R1656 B.n983 B.n6 10.6151
R1657 B.n983 B.n982 10.6151
R1658 B.n982 B.n981 10.6151
R1659 B.n981 B.n8 10.6151
R1660 B.n977 B.n8 10.6151
R1661 B.n977 B.n976 10.6151
R1662 B.n976 B.n975 10.6151
R1663 B.n975 B.n10 10.6151
R1664 B.n971 B.n10 10.6151
R1665 B.n971 B.n970 10.6151
R1666 B.n970 B.n969 10.6151
R1667 B.n969 B.n12 10.6151
R1668 B.n965 B.n12 10.6151
R1669 B.n965 B.n964 10.6151
R1670 B.n964 B.n963 10.6151
R1671 B.n963 B.n14 10.6151
R1672 B.n959 B.n14 10.6151
R1673 B.n959 B.n958 10.6151
R1674 B.n958 B.n957 10.6151
R1675 B.n957 B.n16 10.6151
R1676 B.n953 B.n16 10.6151
R1677 B.n953 B.n952 10.6151
R1678 B.n952 B.n951 10.6151
R1679 B.n951 B.n18 10.6151
R1680 B.n947 B.n18 10.6151
R1681 B.n947 B.n946 10.6151
R1682 B.n946 B.n945 10.6151
R1683 B.n945 B.n20 10.6151
R1684 B.n941 B.n20 10.6151
R1685 B.n941 B.n940 10.6151
R1686 B.n940 B.n939 10.6151
R1687 B.n939 B.n22 10.6151
R1688 B.n935 B.n22 10.6151
R1689 B.n935 B.n934 10.6151
R1690 B.n934 B.n933 10.6151
R1691 B.n933 B.n24 10.6151
R1692 B.n929 B.n24 10.6151
R1693 B.n929 B.n928 10.6151
R1694 B.n928 B.n927 10.6151
R1695 B.n927 B.n26 10.6151
R1696 B.n923 B.n26 10.6151
R1697 B.n923 B.n922 10.6151
R1698 B.n922 B.n921 10.6151
R1699 B.n921 B.n28 10.6151
R1700 B.n917 B.n28 10.6151
R1701 B.n917 B.n916 10.6151
R1702 B.n916 B.n915 10.6151
R1703 B.n915 B.n30 10.6151
R1704 B.n911 B.n30 10.6151
R1705 B.n911 B.n910 10.6151
R1706 B.n910 B.n909 10.6151
R1707 B.n821 B.n820 9.36635
R1708 B.n803 B.n70 9.36635
R1709 B.n431 B.n198 9.36635
R1710 B.n449 B.n448 9.36635
R1711 B.n999 B.n0 2.81026
R1712 B.n999 B.n1 2.81026
R1713 B.n820 B.n819 1.24928
R1714 B.n806 B.n70 1.24928
R1715 B.n434 B.n198 1.24928
R1716 B.n448 B.n447 1.24928
R1717 VN.n11 VN.t3 196.298
R1718 VN.n53 VN.t8 196.298
R1719 VN.n10 VN.t7 164.065
R1720 VN.n21 VN.t5 164.065
R1721 VN.n3 VN.t6 164.065
R1722 VN.n40 VN.t1 164.065
R1723 VN.n52 VN.t4 164.065
R1724 VN.n63 VN.t0 164.065
R1725 VN.n45 VN.t9 164.065
R1726 VN.n82 VN.t2 164.065
R1727 VN.n81 VN.n42 161.3
R1728 VN.n80 VN.n79 161.3
R1729 VN.n78 VN.n43 161.3
R1730 VN.n77 VN.n76 161.3
R1731 VN.n75 VN.n44 161.3
R1732 VN.n74 VN.n73 161.3
R1733 VN.n72 VN.n71 161.3
R1734 VN.n70 VN.n46 161.3
R1735 VN.n69 VN.n68 161.3
R1736 VN.n67 VN.n47 161.3
R1737 VN.n66 VN.n65 161.3
R1738 VN.n64 VN.n48 161.3
R1739 VN.n62 VN.n61 161.3
R1740 VN.n60 VN.n49 161.3
R1741 VN.n59 VN.n58 161.3
R1742 VN.n57 VN.n50 161.3
R1743 VN.n56 VN.n55 161.3
R1744 VN.n54 VN.n51 161.3
R1745 VN.n39 VN.n0 161.3
R1746 VN.n38 VN.n37 161.3
R1747 VN.n36 VN.n1 161.3
R1748 VN.n35 VN.n34 161.3
R1749 VN.n33 VN.n2 161.3
R1750 VN.n32 VN.n31 161.3
R1751 VN.n30 VN.n29 161.3
R1752 VN.n28 VN.n4 161.3
R1753 VN.n27 VN.n26 161.3
R1754 VN.n25 VN.n5 161.3
R1755 VN.n24 VN.n23 161.3
R1756 VN.n22 VN.n6 161.3
R1757 VN.n20 VN.n19 161.3
R1758 VN.n18 VN.n7 161.3
R1759 VN.n17 VN.n16 161.3
R1760 VN.n15 VN.n8 161.3
R1761 VN.n14 VN.n13 161.3
R1762 VN.n12 VN.n9 161.3
R1763 VN.n41 VN.n40 105.499
R1764 VN.n83 VN.n82 105.499
R1765 VN.n11 VN.n10 63.762
R1766 VN.n53 VN.n52 63.762
R1767 VN VN.n83 57.6611
R1768 VN.n16 VN.n15 56.5617
R1769 VN.n58 VN.n57 56.5617
R1770 VN.n27 VN.n5 56.5617
R1771 VN.n69 VN.n47 56.5617
R1772 VN.n34 VN.n1 54.6242
R1773 VN.n76 VN.n43 54.6242
R1774 VN.n34 VN.n33 26.5299
R1775 VN.n76 VN.n75 26.5299
R1776 VN.n14 VN.n9 24.5923
R1777 VN.n15 VN.n14 24.5923
R1778 VN.n16 VN.n7 24.5923
R1779 VN.n20 VN.n7 24.5923
R1780 VN.n23 VN.n22 24.5923
R1781 VN.n23 VN.n5 24.5923
R1782 VN.n28 VN.n27 24.5923
R1783 VN.n29 VN.n28 24.5923
R1784 VN.n33 VN.n32 24.5923
R1785 VN.n38 VN.n1 24.5923
R1786 VN.n39 VN.n38 24.5923
R1787 VN.n57 VN.n56 24.5923
R1788 VN.n56 VN.n51 24.5923
R1789 VN.n65 VN.n47 24.5923
R1790 VN.n65 VN.n64 24.5923
R1791 VN.n62 VN.n49 24.5923
R1792 VN.n58 VN.n49 24.5923
R1793 VN.n75 VN.n74 24.5923
R1794 VN.n71 VN.n70 24.5923
R1795 VN.n70 VN.n69 24.5923
R1796 VN.n81 VN.n80 24.5923
R1797 VN.n80 VN.n43 24.5923
R1798 VN.n32 VN.n3 15.7393
R1799 VN.n74 VN.n45 15.7393
R1800 VN.n21 VN.n20 12.2964
R1801 VN.n22 VN.n21 12.2964
R1802 VN.n64 VN.n63 12.2964
R1803 VN.n63 VN.n62 12.2964
R1804 VN.n10 VN.n9 8.85356
R1805 VN.n29 VN.n3 8.85356
R1806 VN.n52 VN.n51 8.85356
R1807 VN.n71 VN.n45 8.85356
R1808 VN.n54 VN.n53 7.12066
R1809 VN.n12 VN.n11 7.12066
R1810 VN.n40 VN.n39 5.4107
R1811 VN.n82 VN.n81 5.4107
R1812 VN.n83 VN.n42 0.278335
R1813 VN.n41 VN.n0 0.278335
R1814 VN.n79 VN.n42 0.189894
R1815 VN.n79 VN.n78 0.189894
R1816 VN.n78 VN.n77 0.189894
R1817 VN.n77 VN.n44 0.189894
R1818 VN.n73 VN.n44 0.189894
R1819 VN.n73 VN.n72 0.189894
R1820 VN.n72 VN.n46 0.189894
R1821 VN.n68 VN.n46 0.189894
R1822 VN.n68 VN.n67 0.189894
R1823 VN.n67 VN.n66 0.189894
R1824 VN.n66 VN.n48 0.189894
R1825 VN.n61 VN.n48 0.189894
R1826 VN.n61 VN.n60 0.189894
R1827 VN.n60 VN.n59 0.189894
R1828 VN.n59 VN.n50 0.189894
R1829 VN.n55 VN.n50 0.189894
R1830 VN.n55 VN.n54 0.189894
R1831 VN.n13 VN.n12 0.189894
R1832 VN.n13 VN.n8 0.189894
R1833 VN.n17 VN.n8 0.189894
R1834 VN.n18 VN.n17 0.189894
R1835 VN.n19 VN.n18 0.189894
R1836 VN.n19 VN.n6 0.189894
R1837 VN.n24 VN.n6 0.189894
R1838 VN.n25 VN.n24 0.189894
R1839 VN.n26 VN.n25 0.189894
R1840 VN.n26 VN.n4 0.189894
R1841 VN.n30 VN.n4 0.189894
R1842 VN.n31 VN.n30 0.189894
R1843 VN.n31 VN.n2 0.189894
R1844 VN.n35 VN.n2 0.189894
R1845 VN.n36 VN.n35 0.189894
R1846 VN.n37 VN.n36 0.189894
R1847 VN.n37 VN.n0 0.189894
R1848 VN VN.n41 0.153485
R1849 VDD2.n1 VDD2.t6 76.3266
R1850 VDD2.n3 VDD2.n2 73.8033
R1851 VDD2.n4 VDD2.t7 73.8017
R1852 VDD2 VDD2.n7 73.8004
R1853 VDD2.n6 VDD2.n5 71.9653
R1854 VDD2.n1 VDD2.n0 71.9643
R1855 VDD2.n4 VDD2.n3 50.9718
R1856 VDD2.n6 VDD2.n4 2.52636
R1857 VDD2.n7 VDD2.t5 1.83694
R1858 VDD2.n7 VDD2.t1 1.83694
R1859 VDD2.n5 VDD2.t0 1.83694
R1860 VDD2.n5 VDD2.t9 1.83694
R1861 VDD2.n2 VDD2.t3 1.83694
R1862 VDD2.n2 VDD2.t8 1.83694
R1863 VDD2.n0 VDD2.t2 1.83694
R1864 VDD2.n0 VDD2.t4 1.83694
R1865 VDD2 VDD2.n6 0.690155
R1866 VDD2.n3 VDD2.n1 0.576619
C0 VDD2 VP 0.584482f
C1 VDD2 VN 15.488201f
C2 VTAIL VP 15.889299f
C3 VDD2 VDD1 2.17587f
C4 w_n4486_n4508# B 12.145201f
C5 VTAIL VN 15.8749f
C6 VTAIL VDD1 13.021501f
C7 VDD2 VTAIL 13.071199f
C8 w_n4486_n4508# VP 10.2734f
C9 B VP 2.33617f
C10 VN w_n4486_n4508# 9.689361f
C11 VN B 1.35405f
C12 w_n4486_n4508# VDD1 3.18688f
C13 B VDD1 2.93065f
C14 VDD2 w_n4486_n4508# 3.33043f
C15 VDD2 B 3.04857f
C16 VTAIL w_n4486_n4508# 4.00983f
C17 VTAIL B 5.00816f
C18 VN VP 9.44909f
C19 VP VDD1 15.914001f
C20 VN VDD1 0.153807f
C21 VDD2 VSUBS 2.27584f
C22 VDD1 VSUBS 2.112327f
C23 VTAIL VSUBS 1.490927f
C24 VN VSUBS 7.89326f
C25 VP VSUBS 4.442738f
C26 B VSUBS 5.84942f
C27 w_n4486_n4508# VSUBS 0.247358p
C28 VDD2.t6 VSUBS 4.32701f
C29 VDD2.t2 VSUBS 0.396755f
C30 VDD2.t4 VSUBS 0.396755f
C31 VDD2.n0 VSUBS 3.3156f
C32 VDD2.n1 VSUBS 1.66112f
C33 VDD2.t3 VSUBS 0.396755f
C34 VDD2.t8 VSUBS 0.396755f
C35 VDD2.n2 VSUBS 3.33909f
C36 VDD2.n3 VSUBS 3.99456f
C37 VDD2.t7 VSUBS 4.2981f
C38 VDD2.n4 VSUBS 4.36088f
C39 VDD2.t0 VSUBS 0.396755f
C40 VDD2.t9 VSUBS 0.396755f
C41 VDD2.n5 VSUBS 3.3156f
C42 VDD2.n6 VSUBS 0.825664f
C43 VDD2.t5 VSUBS 0.396755f
C44 VDD2.t1 VSUBS 0.396755f
C45 VDD2.n7 VSUBS 3.33902f
C46 VN.n0 VSUBS 0.033561f
C47 VN.t1 VSUBS 3.2214f
C48 VN.n1 VSUBS 0.044133f
C49 VN.n2 VSUBS 0.025457f
C50 VN.t6 VSUBS 3.2214f
C51 VN.n3 VSUBS 1.11772f
C52 VN.n4 VSUBS 0.025457f
C53 VN.n5 VSUBS 0.034541f
C54 VN.n6 VSUBS 0.025457f
C55 VN.t5 VSUBS 3.2214f
C56 VN.n7 VSUBS 0.047208f
C57 VN.n8 VSUBS 0.025457f
C58 VN.n9 VSUBS 0.032293f
C59 VN.t3 VSUBS 3.43034f
C60 VN.t7 VSUBS 3.2214f
C61 VN.n10 VSUBS 1.18764f
C62 VN.n11 VSUBS 1.16772f
C63 VN.n12 VSUBS 0.245748f
C64 VN.n13 VSUBS 0.025457f
C65 VN.n14 VSUBS 0.047208f
C66 VN.n15 VSUBS 0.039471f
C67 VN.n16 VSUBS 0.034541f
C68 VN.n17 VSUBS 0.025457f
C69 VN.n18 VSUBS 0.025457f
C70 VN.n19 VSUBS 0.025457f
C71 VN.n20 VSUBS 0.035556f
C72 VN.n21 VSUBS 1.11772f
C73 VN.n22 VSUBS 0.035556f
C74 VN.n23 VSUBS 0.047208f
C75 VN.n24 VSUBS 0.025457f
C76 VN.n25 VSUBS 0.025457f
C77 VN.n26 VSUBS 0.025457f
C78 VN.n27 VSUBS 0.039471f
C79 VN.n28 VSUBS 0.047208f
C80 VN.n29 VSUBS 0.032293f
C81 VN.n30 VSUBS 0.025457f
C82 VN.n31 VSUBS 0.025457f
C83 VN.n32 VSUBS 0.038818f
C84 VN.n33 VSUBS 0.048774f
C85 VN.n34 VSUBS 0.028313f
C86 VN.n35 VSUBS 0.025457f
C87 VN.n36 VSUBS 0.025457f
C88 VN.n37 VSUBS 0.025457f
C89 VN.n38 VSUBS 0.047208f
C90 VN.n39 VSUBS 0.02903f
C91 VN.n40 VSUBS 1.19625f
C92 VN.n41 VSUBS 0.044147f
C93 VN.n42 VSUBS 0.033561f
C94 VN.t2 VSUBS 3.2214f
C95 VN.n43 VSUBS 0.044133f
C96 VN.n44 VSUBS 0.025457f
C97 VN.t9 VSUBS 3.2214f
C98 VN.n45 VSUBS 1.11772f
C99 VN.n46 VSUBS 0.025457f
C100 VN.n47 VSUBS 0.034541f
C101 VN.n48 VSUBS 0.025457f
C102 VN.t0 VSUBS 3.2214f
C103 VN.n49 VSUBS 0.047208f
C104 VN.n50 VSUBS 0.025457f
C105 VN.n51 VSUBS 0.032293f
C106 VN.t8 VSUBS 3.43034f
C107 VN.t4 VSUBS 3.2214f
C108 VN.n52 VSUBS 1.18764f
C109 VN.n53 VSUBS 1.16772f
C110 VN.n54 VSUBS 0.245748f
C111 VN.n55 VSUBS 0.025457f
C112 VN.n56 VSUBS 0.047208f
C113 VN.n57 VSUBS 0.039471f
C114 VN.n58 VSUBS 0.034541f
C115 VN.n59 VSUBS 0.025457f
C116 VN.n60 VSUBS 0.025457f
C117 VN.n61 VSUBS 0.025457f
C118 VN.n62 VSUBS 0.035556f
C119 VN.n63 VSUBS 1.11772f
C120 VN.n64 VSUBS 0.035556f
C121 VN.n65 VSUBS 0.047208f
C122 VN.n66 VSUBS 0.025457f
C123 VN.n67 VSUBS 0.025457f
C124 VN.n68 VSUBS 0.025457f
C125 VN.n69 VSUBS 0.039471f
C126 VN.n70 VSUBS 0.047208f
C127 VN.n71 VSUBS 0.032293f
C128 VN.n72 VSUBS 0.025457f
C129 VN.n73 VSUBS 0.025457f
C130 VN.n74 VSUBS 0.038818f
C131 VN.n75 VSUBS 0.048774f
C132 VN.n76 VSUBS 0.028313f
C133 VN.n77 VSUBS 0.025457f
C134 VN.n78 VSUBS 0.025457f
C135 VN.n79 VSUBS 0.025457f
C136 VN.n80 VSUBS 0.047208f
C137 VN.n81 VSUBS 0.02903f
C138 VN.n82 VSUBS 1.19625f
C139 VN.n83 VSUBS 1.73907f
C140 B.n0 VSUBS 0.005137f
C141 B.n1 VSUBS 0.005137f
C142 B.n2 VSUBS 0.008123f
C143 B.n3 VSUBS 0.008123f
C144 B.n4 VSUBS 0.008123f
C145 B.n5 VSUBS 0.008123f
C146 B.n6 VSUBS 0.008123f
C147 B.n7 VSUBS 0.008123f
C148 B.n8 VSUBS 0.008123f
C149 B.n9 VSUBS 0.008123f
C150 B.n10 VSUBS 0.008123f
C151 B.n11 VSUBS 0.008123f
C152 B.n12 VSUBS 0.008123f
C153 B.n13 VSUBS 0.008123f
C154 B.n14 VSUBS 0.008123f
C155 B.n15 VSUBS 0.008123f
C156 B.n16 VSUBS 0.008123f
C157 B.n17 VSUBS 0.008123f
C158 B.n18 VSUBS 0.008123f
C159 B.n19 VSUBS 0.008123f
C160 B.n20 VSUBS 0.008123f
C161 B.n21 VSUBS 0.008123f
C162 B.n22 VSUBS 0.008123f
C163 B.n23 VSUBS 0.008123f
C164 B.n24 VSUBS 0.008123f
C165 B.n25 VSUBS 0.008123f
C166 B.n26 VSUBS 0.008123f
C167 B.n27 VSUBS 0.008123f
C168 B.n28 VSUBS 0.008123f
C169 B.n29 VSUBS 0.008123f
C170 B.n30 VSUBS 0.008123f
C171 B.n31 VSUBS 0.008123f
C172 B.n32 VSUBS 0.019052f
C173 B.n33 VSUBS 0.008123f
C174 B.n34 VSUBS 0.008123f
C175 B.n35 VSUBS 0.008123f
C176 B.n36 VSUBS 0.008123f
C177 B.n37 VSUBS 0.008123f
C178 B.n38 VSUBS 0.008123f
C179 B.n39 VSUBS 0.008123f
C180 B.n40 VSUBS 0.008123f
C181 B.n41 VSUBS 0.008123f
C182 B.n42 VSUBS 0.008123f
C183 B.n43 VSUBS 0.008123f
C184 B.n44 VSUBS 0.008123f
C185 B.n45 VSUBS 0.008123f
C186 B.n46 VSUBS 0.008123f
C187 B.n47 VSUBS 0.008123f
C188 B.n48 VSUBS 0.008123f
C189 B.n49 VSUBS 0.008123f
C190 B.n50 VSUBS 0.008123f
C191 B.n51 VSUBS 0.008123f
C192 B.n52 VSUBS 0.008123f
C193 B.n53 VSUBS 0.008123f
C194 B.n54 VSUBS 0.008123f
C195 B.n55 VSUBS 0.008123f
C196 B.n56 VSUBS 0.008123f
C197 B.n57 VSUBS 0.008123f
C198 B.n58 VSUBS 0.008123f
C199 B.n59 VSUBS 0.008123f
C200 B.n60 VSUBS 0.008123f
C201 B.n61 VSUBS 0.008123f
C202 B.t2 VSUBS 0.692556f
C203 B.t1 VSUBS 0.717637f
C204 B.t0 VSUBS 2.3716f
C205 B.n62 VSUBS 0.391662f
C206 B.n63 VSUBS 0.083719f
C207 B.n64 VSUBS 0.008123f
C208 B.n65 VSUBS 0.008123f
C209 B.n66 VSUBS 0.008123f
C210 B.n67 VSUBS 0.008123f
C211 B.t5 VSUBS 0.69253f
C212 B.t4 VSUBS 0.717617f
C213 B.t3 VSUBS 2.3716f
C214 B.n68 VSUBS 0.391682f
C215 B.n69 VSUBS 0.083745f
C216 B.n70 VSUBS 0.018821f
C217 B.n71 VSUBS 0.008123f
C218 B.n72 VSUBS 0.008123f
C219 B.n73 VSUBS 0.008123f
C220 B.n74 VSUBS 0.008123f
C221 B.n75 VSUBS 0.008123f
C222 B.n76 VSUBS 0.008123f
C223 B.n77 VSUBS 0.008123f
C224 B.n78 VSUBS 0.008123f
C225 B.n79 VSUBS 0.008123f
C226 B.n80 VSUBS 0.008123f
C227 B.n81 VSUBS 0.008123f
C228 B.n82 VSUBS 0.008123f
C229 B.n83 VSUBS 0.008123f
C230 B.n84 VSUBS 0.008123f
C231 B.n85 VSUBS 0.008123f
C232 B.n86 VSUBS 0.008123f
C233 B.n87 VSUBS 0.008123f
C234 B.n88 VSUBS 0.008123f
C235 B.n89 VSUBS 0.008123f
C236 B.n90 VSUBS 0.008123f
C237 B.n91 VSUBS 0.008123f
C238 B.n92 VSUBS 0.008123f
C239 B.n93 VSUBS 0.008123f
C240 B.n94 VSUBS 0.008123f
C241 B.n95 VSUBS 0.008123f
C242 B.n96 VSUBS 0.008123f
C243 B.n97 VSUBS 0.008123f
C244 B.n98 VSUBS 0.008123f
C245 B.n99 VSUBS 0.019052f
C246 B.n100 VSUBS 0.008123f
C247 B.n101 VSUBS 0.008123f
C248 B.n102 VSUBS 0.008123f
C249 B.n103 VSUBS 0.008123f
C250 B.n104 VSUBS 0.008123f
C251 B.n105 VSUBS 0.008123f
C252 B.n106 VSUBS 0.008123f
C253 B.n107 VSUBS 0.008123f
C254 B.n108 VSUBS 0.008123f
C255 B.n109 VSUBS 0.008123f
C256 B.n110 VSUBS 0.008123f
C257 B.n111 VSUBS 0.008123f
C258 B.n112 VSUBS 0.008123f
C259 B.n113 VSUBS 0.008123f
C260 B.n114 VSUBS 0.008123f
C261 B.n115 VSUBS 0.008123f
C262 B.n116 VSUBS 0.008123f
C263 B.n117 VSUBS 0.008123f
C264 B.n118 VSUBS 0.008123f
C265 B.n119 VSUBS 0.008123f
C266 B.n120 VSUBS 0.008123f
C267 B.n121 VSUBS 0.008123f
C268 B.n122 VSUBS 0.008123f
C269 B.n123 VSUBS 0.008123f
C270 B.n124 VSUBS 0.008123f
C271 B.n125 VSUBS 0.008123f
C272 B.n126 VSUBS 0.008123f
C273 B.n127 VSUBS 0.008123f
C274 B.n128 VSUBS 0.008123f
C275 B.n129 VSUBS 0.008123f
C276 B.n130 VSUBS 0.008123f
C277 B.n131 VSUBS 0.008123f
C278 B.n132 VSUBS 0.008123f
C279 B.n133 VSUBS 0.008123f
C280 B.n134 VSUBS 0.008123f
C281 B.n135 VSUBS 0.008123f
C282 B.n136 VSUBS 0.008123f
C283 B.n137 VSUBS 0.008123f
C284 B.n138 VSUBS 0.008123f
C285 B.n139 VSUBS 0.008123f
C286 B.n140 VSUBS 0.008123f
C287 B.n141 VSUBS 0.008123f
C288 B.n142 VSUBS 0.008123f
C289 B.n143 VSUBS 0.008123f
C290 B.n144 VSUBS 0.008123f
C291 B.n145 VSUBS 0.008123f
C292 B.n146 VSUBS 0.008123f
C293 B.n147 VSUBS 0.008123f
C294 B.n148 VSUBS 0.008123f
C295 B.n149 VSUBS 0.008123f
C296 B.n150 VSUBS 0.008123f
C297 B.n151 VSUBS 0.008123f
C298 B.n152 VSUBS 0.008123f
C299 B.n153 VSUBS 0.008123f
C300 B.n154 VSUBS 0.008123f
C301 B.n155 VSUBS 0.008123f
C302 B.n156 VSUBS 0.008123f
C303 B.n157 VSUBS 0.008123f
C304 B.n158 VSUBS 0.008123f
C305 B.n159 VSUBS 0.008123f
C306 B.n160 VSUBS 0.019052f
C307 B.n161 VSUBS 0.008123f
C308 B.n162 VSUBS 0.008123f
C309 B.n163 VSUBS 0.008123f
C310 B.n164 VSUBS 0.008123f
C311 B.n165 VSUBS 0.008123f
C312 B.n166 VSUBS 0.008123f
C313 B.n167 VSUBS 0.008123f
C314 B.n168 VSUBS 0.008123f
C315 B.n169 VSUBS 0.008123f
C316 B.n170 VSUBS 0.008123f
C317 B.n171 VSUBS 0.008123f
C318 B.n172 VSUBS 0.008123f
C319 B.n173 VSUBS 0.008123f
C320 B.n174 VSUBS 0.008123f
C321 B.n175 VSUBS 0.008123f
C322 B.n176 VSUBS 0.008123f
C323 B.n177 VSUBS 0.008123f
C324 B.n178 VSUBS 0.008123f
C325 B.n179 VSUBS 0.008123f
C326 B.n180 VSUBS 0.008123f
C327 B.n181 VSUBS 0.008123f
C328 B.n182 VSUBS 0.008123f
C329 B.n183 VSUBS 0.008123f
C330 B.n184 VSUBS 0.008123f
C331 B.n185 VSUBS 0.008123f
C332 B.n186 VSUBS 0.008123f
C333 B.n187 VSUBS 0.008123f
C334 B.n188 VSUBS 0.008123f
C335 B.n189 VSUBS 0.008123f
C336 B.t10 VSUBS 0.69253f
C337 B.t11 VSUBS 0.717617f
C338 B.t9 VSUBS 2.3716f
C339 B.n190 VSUBS 0.391682f
C340 B.n191 VSUBS 0.083745f
C341 B.n192 VSUBS 0.008123f
C342 B.n193 VSUBS 0.008123f
C343 B.n194 VSUBS 0.008123f
C344 B.n195 VSUBS 0.008123f
C345 B.t7 VSUBS 0.692556f
C346 B.t8 VSUBS 0.717637f
C347 B.t6 VSUBS 2.3716f
C348 B.n196 VSUBS 0.391662f
C349 B.n197 VSUBS 0.083719f
C350 B.n198 VSUBS 0.018821f
C351 B.n199 VSUBS 0.008123f
C352 B.n200 VSUBS 0.008123f
C353 B.n201 VSUBS 0.008123f
C354 B.n202 VSUBS 0.008123f
C355 B.n203 VSUBS 0.008123f
C356 B.n204 VSUBS 0.008123f
C357 B.n205 VSUBS 0.008123f
C358 B.n206 VSUBS 0.008123f
C359 B.n207 VSUBS 0.008123f
C360 B.n208 VSUBS 0.008123f
C361 B.n209 VSUBS 0.008123f
C362 B.n210 VSUBS 0.008123f
C363 B.n211 VSUBS 0.008123f
C364 B.n212 VSUBS 0.008123f
C365 B.n213 VSUBS 0.008123f
C366 B.n214 VSUBS 0.008123f
C367 B.n215 VSUBS 0.008123f
C368 B.n216 VSUBS 0.008123f
C369 B.n217 VSUBS 0.008123f
C370 B.n218 VSUBS 0.008123f
C371 B.n219 VSUBS 0.008123f
C372 B.n220 VSUBS 0.008123f
C373 B.n221 VSUBS 0.008123f
C374 B.n222 VSUBS 0.008123f
C375 B.n223 VSUBS 0.008123f
C376 B.n224 VSUBS 0.008123f
C377 B.n225 VSUBS 0.008123f
C378 B.n226 VSUBS 0.008123f
C379 B.n227 VSUBS 0.019052f
C380 B.n228 VSUBS 0.008123f
C381 B.n229 VSUBS 0.008123f
C382 B.n230 VSUBS 0.008123f
C383 B.n231 VSUBS 0.008123f
C384 B.n232 VSUBS 0.008123f
C385 B.n233 VSUBS 0.008123f
C386 B.n234 VSUBS 0.008123f
C387 B.n235 VSUBS 0.008123f
C388 B.n236 VSUBS 0.008123f
C389 B.n237 VSUBS 0.008123f
C390 B.n238 VSUBS 0.008123f
C391 B.n239 VSUBS 0.008123f
C392 B.n240 VSUBS 0.008123f
C393 B.n241 VSUBS 0.008123f
C394 B.n242 VSUBS 0.008123f
C395 B.n243 VSUBS 0.008123f
C396 B.n244 VSUBS 0.008123f
C397 B.n245 VSUBS 0.008123f
C398 B.n246 VSUBS 0.008123f
C399 B.n247 VSUBS 0.008123f
C400 B.n248 VSUBS 0.008123f
C401 B.n249 VSUBS 0.008123f
C402 B.n250 VSUBS 0.008123f
C403 B.n251 VSUBS 0.008123f
C404 B.n252 VSUBS 0.008123f
C405 B.n253 VSUBS 0.008123f
C406 B.n254 VSUBS 0.008123f
C407 B.n255 VSUBS 0.008123f
C408 B.n256 VSUBS 0.008123f
C409 B.n257 VSUBS 0.008123f
C410 B.n258 VSUBS 0.008123f
C411 B.n259 VSUBS 0.008123f
C412 B.n260 VSUBS 0.008123f
C413 B.n261 VSUBS 0.008123f
C414 B.n262 VSUBS 0.008123f
C415 B.n263 VSUBS 0.008123f
C416 B.n264 VSUBS 0.008123f
C417 B.n265 VSUBS 0.008123f
C418 B.n266 VSUBS 0.008123f
C419 B.n267 VSUBS 0.008123f
C420 B.n268 VSUBS 0.008123f
C421 B.n269 VSUBS 0.008123f
C422 B.n270 VSUBS 0.008123f
C423 B.n271 VSUBS 0.008123f
C424 B.n272 VSUBS 0.008123f
C425 B.n273 VSUBS 0.008123f
C426 B.n274 VSUBS 0.008123f
C427 B.n275 VSUBS 0.008123f
C428 B.n276 VSUBS 0.008123f
C429 B.n277 VSUBS 0.008123f
C430 B.n278 VSUBS 0.008123f
C431 B.n279 VSUBS 0.008123f
C432 B.n280 VSUBS 0.008123f
C433 B.n281 VSUBS 0.008123f
C434 B.n282 VSUBS 0.008123f
C435 B.n283 VSUBS 0.008123f
C436 B.n284 VSUBS 0.008123f
C437 B.n285 VSUBS 0.008123f
C438 B.n286 VSUBS 0.008123f
C439 B.n287 VSUBS 0.008123f
C440 B.n288 VSUBS 0.008123f
C441 B.n289 VSUBS 0.008123f
C442 B.n290 VSUBS 0.008123f
C443 B.n291 VSUBS 0.008123f
C444 B.n292 VSUBS 0.008123f
C445 B.n293 VSUBS 0.008123f
C446 B.n294 VSUBS 0.008123f
C447 B.n295 VSUBS 0.008123f
C448 B.n296 VSUBS 0.008123f
C449 B.n297 VSUBS 0.008123f
C450 B.n298 VSUBS 0.008123f
C451 B.n299 VSUBS 0.008123f
C452 B.n300 VSUBS 0.008123f
C453 B.n301 VSUBS 0.008123f
C454 B.n302 VSUBS 0.008123f
C455 B.n303 VSUBS 0.008123f
C456 B.n304 VSUBS 0.008123f
C457 B.n305 VSUBS 0.008123f
C458 B.n306 VSUBS 0.008123f
C459 B.n307 VSUBS 0.008123f
C460 B.n308 VSUBS 0.008123f
C461 B.n309 VSUBS 0.008123f
C462 B.n310 VSUBS 0.008123f
C463 B.n311 VSUBS 0.008123f
C464 B.n312 VSUBS 0.008123f
C465 B.n313 VSUBS 0.008123f
C466 B.n314 VSUBS 0.008123f
C467 B.n315 VSUBS 0.008123f
C468 B.n316 VSUBS 0.008123f
C469 B.n317 VSUBS 0.008123f
C470 B.n318 VSUBS 0.008123f
C471 B.n319 VSUBS 0.008123f
C472 B.n320 VSUBS 0.008123f
C473 B.n321 VSUBS 0.008123f
C474 B.n322 VSUBS 0.008123f
C475 B.n323 VSUBS 0.008123f
C476 B.n324 VSUBS 0.008123f
C477 B.n325 VSUBS 0.008123f
C478 B.n326 VSUBS 0.008123f
C479 B.n327 VSUBS 0.008123f
C480 B.n328 VSUBS 0.008123f
C481 B.n329 VSUBS 0.008123f
C482 B.n330 VSUBS 0.008123f
C483 B.n331 VSUBS 0.008123f
C484 B.n332 VSUBS 0.008123f
C485 B.n333 VSUBS 0.008123f
C486 B.n334 VSUBS 0.008123f
C487 B.n335 VSUBS 0.008123f
C488 B.n336 VSUBS 0.008123f
C489 B.n337 VSUBS 0.008123f
C490 B.n338 VSUBS 0.008123f
C491 B.n339 VSUBS 0.008123f
C492 B.n340 VSUBS 0.008123f
C493 B.n341 VSUBS 0.008123f
C494 B.n342 VSUBS 0.008123f
C495 B.n343 VSUBS 0.008123f
C496 B.n344 VSUBS 0.018697f
C497 B.n345 VSUBS 0.018697f
C498 B.n346 VSUBS 0.019052f
C499 B.n347 VSUBS 0.008123f
C500 B.n348 VSUBS 0.008123f
C501 B.n349 VSUBS 0.008123f
C502 B.n350 VSUBS 0.008123f
C503 B.n351 VSUBS 0.008123f
C504 B.n352 VSUBS 0.008123f
C505 B.n353 VSUBS 0.008123f
C506 B.n354 VSUBS 0.008123f
C507 B.n355 VSUBS 0.008123f
C508 B.n356 VSUBS 0.008123f
C509 B.n357 VSUBS 0.008123f
C510 B.n358 VSUBS 0.008123f
C511 B.n359 VSUBS 0.008123f
C512 B.n360 VSUBS 0.008123f
C513 B.n361 VSUBS 0.008123f
C514 B.n362 VSUBS 0.008123f
C515 B.n363 VSUBS 0.008123f
C516 B.n364 VSUBS 0.008123f
C517 B.n365 VSUBS 0.008123f
C518 B.n366 VSUBS 0.008123f
C519 B.n367 VSUBS 0.008123f
C520 B.n368 VSUBS 0.008123f
C521 B.n369 VSUBS 0.008123f
C522 B.n370 VSUBS 0.008123f
C523 B.n371 VSUBS 0.008123f
C524 B.n372 VSUBS 0.008123f
C525 B.n373 VSUBS 0.008123f
C526 B.n374 VSUBS 0.008123f
C527 B.n375 VSUBS 0.008123f
C528 B.n376 VSUBS 0.008123f
C529 B.n377 VSUBS 0.008123f
C530 B.n378 VSUBS 0.008123f
C531 B.n379 VSUBS 0.008123f
C532 B.n380 VSUBS 0.008123f
C533 B.n381 VSUBS 0.008123f
C534 B.n382 VSUBS 0.008123f
C535 B.n383 VSUBS 0.008123f
C536 B.n384 VSUBS 0.008123f
C537 B.n385 VSUBS 0.008123f
C538 B.n386 VSUBS 0.008123f
C539 B.n387 VSUBS 0.008123f
C540 B.n388 VSUBS 0.008123f
C541 B.n389 VSUBS 0.008123f
C542 B.n390 VSUBS 0.008123f
C543 B.n391 VSUBS 0.008123f
C544 B.n392 VSUBS 0.008123f
C545 B.n393 VSUBS 0.008123f
C546 B.n394 VSUBS 0.008123f
C547 B.n395 VSUBS 0.008123f
C548 B.n396 VSUBS 0.008123f
C549 B.n397 VSUBS 0.008123f
C550 B.n398 VSUBS 0.008123f
C551 B.n399 VSUBS 0.008123f
C552 B.n400 VSUBS 0.008123f
C553 B.n401 VSUBS 0.008123f
C554 B.n402 VSUBS 0.008123f
C555 B.n403 VSUBS 0.008123f
C556 B.n404 VSUBS 0.008123f
C557 B.n405 VSUBS 0.008123f
C558 B.n406 VSUBS 0.008123f
C559 B.n407 VSUBS 0.008123f
C560 B.n408 VSUBS 0.008123f
C561 B.n409 VSUBS 0.008123f
C562 B.n410 VSUBS 0.008123f
C563 B.n411 VSUBS 0.008123f
C564 B.n412 VSUBS 0.008123f
C565 B.n413 VSUBS 0.008123f
C566 B.n414 VSUBS 0.008123f
C567 B.n415 VSUBS 0.008123f
C568 B.n416 VSUBS 0.008123f
C569 B.n417 VSUBS 0.008123f
C570 B.n418 VSUBS 0.008123f
C571 B.n419 VSUBS 0.008123f
C572 B.n420 VSUBS 0.008123f
C573 B.n421 VSUBS 0.008123f
C574 B.n422 VSUBS 0.008123f
C575 B.n423 VSUBS 0.008123f
C576 B.n424 VSUBS 0.008123f
C577 B.n425 VSUBS 0.008123f
C578 B.n426 VSUBS 0.008123f
C579 B.n427 VSUBS 0.008123f
C580 B.n428 VSUBS 0.008123f
C581 B.n429 VSUBS 0.008123f
C582 B.n430 VSUBS 0.008123f
C583 B.n431 VSUBS 0.007645f
C584 B.n432 VSUBS 0.008123f
C585 B.n433 VSUBS 0.008123f
C586 B.n434 VSUBS 0.004539f
C587 B.n435 VSUBS 0.008123f
C588 B.n436 VSUBS 0.008123f
C589 B.n437 VSUBS 0.008123f
C590 B.n438 VSUBS 0.008123f
C591 B.n439 VSUBS 0.008123f
C592 B.n440 VSUBS 0.008123f
C593 B.n441 VSUBS 0.008123f
C594 B.n442 VSUBS 0.008123f
C595 B.n443 VSUBS 0.008123f
C596 B.n444 VSUBS 0.008123f
C597 B.n445 VSUBS 0.008123f
C598 B.n446 VSUBS 0.008123f
C599 B.n447 VSUBS 0.004539f
C600 B.n448 VSUBS 0.018821f
C601 B.n449 VSUBS 0.007645f
C602 B.n450 VSUBS 0.008123f
C603 B.n451 VSUBS 0.008123f
C604 B.n452 VSUBS 0.008123f
C605 B.n453 VSUBS 0.008123f
C606 B.n454 VSUBS 0.008123f
C607 B.n455 VSUBS 0.008123f
C608 B.n456 VSUBS 0.008123f
C609 B.n457 VSUBS 0.008123f
C610 B.n458 VSUBS 0.008123f
C611 B.n459 VSUBS 0.008123f
C612 B.n460 VSUBS 0.008123f
C613 B.n461 VSUBS 0.008123f
C614 B.n462 VSUBS 0.008123f
C615 B.n463 VSUBS 0.008123f
C616 B.n464 VSUBS 0.008123f
C617 B.n465 VSUBS 0.008123f
C618 B.n466 VSUBS 0.008123f
C619 B.n467 VSUBS 0.008123f
C620 B.n468 VSUBS 0.008123f
C621 B.n469 VSUBS 0.008123f
C622 B.n470 VSUBS 0.008123f
C623 B.n471 VSUBS 0.008123f
C624 B.n472 VSUBS 0.008123f
C625 B.n473 VSUBS 0.008123f
C626 B.n474 VSUBS 0.008123f
C627 B.n475 VSUBS 0.008123f
C628 B.n476 VSUBS 0.008123f
C629 B.n477 VSUBS 0.008123f
C630 B.n478 VSUBS 0.008123f
C631 B.n479 VSUBS 0.008123f
C632 B.n480 VSUBS 0.008123f
C633 B.n481 VSUBS 0.008123f
C634 B.n482 VSUBS 0.008123f
C635 B.n483 VSUBS 0.008123f
C636 B.n484 VSUBS 0.008123f
C637 B.n485 VSUBS 0.008123f
C638 B.n486 VSUBS 0.008123f
C639 B.n487 VSUBS 0.008123f
C640 B.n488 VSUBS 0.008123f
C641 B.n489 VSUBS 0.008123f
C642 B.n490 VSUBS 0.008123f
C643 B.n491 VSUBS 0.008123f
C644 B.n492 VSUBS 0.008123f
C645 B.n493 VSUBS 0.008123f
C646 B.n494 VSUBS 0.008123f
C647 B.n495 VSUBS 0.008123f
C648 B.n496 VSUBS 0.008123f
C649 B.n497 VSUBS 0.008123f
C650 B.n498 VSUBS 0.008123f
C651 B.n499 VSUBS 0.008123f
C652 B.n500 VSUBS 0.008123f
C653 B.n501 VSUBS 0.008123f
C654 B.n502 VSUBS 0.008123f
C655 B.n503 VSUBS 0.008123f
C656 B.n504 VSUBS 0.008123f
C657 B.n505 VSUBS 0.008123f
C658 B.n506 VSUBS 0.008123f
C659 B.n507 VSUBS 0.008123f
C660 B.n508 VSUBS 0.008123f
C661 B.n509 VSUBS 0.008123f
C662 B.n510 VSUBS 0.008123f
C663 B.n511 VSUBS 0.008123f
C664 B.n512 VSUBS 0.008123f
C665 B.n513 VSUBS 0.008123f
C666 B.n514 VSUBS 0.008123f
C667 B.n515 VSUBS 0.008123f
C668 B.n516 VSUBS 0.008123f
C669 B.n517 VSUBS 0.008123f
C670 B.n518 VSUBS 0.008123f
C671 B.n519 VSUBS 0.008123f
C672 B.n520 VSUBS 0.008123f
C673 B.n521 VSUBS 0.008123f
C674 B.n522 VSUBS 0.008123f
C675 B.n523 VSUBS 0.008123f
C676 B.n524 VSUBS 0.008123f
C677 B.n525 VSUBS 0.008123f
C678 B.n526 VSUBS 0.008123f
C679 B.n527 VSUBS 0.008123f
C680 B.n528 VSUBS 0.008123f
C681 B.n529 VSUBS 0.008123f
C682 B.n530 VSUBS 0.008123f
C683 B.n531 VSUBS 0.008123f
C684 B.n532 VSUBS 0.008123f
C685 B.n533 VSUBS 0.008123f
C686 B.n534 VSUBS 0.008123f
C687 B.n535 VSUBS 0.019052f
C688 B.n536 VSUBS 0.018697f
C689 B.n537 VSUBS 0.018697f
C690 B.n538 VSUBS 0.008123f
C691 B.n539 VSUBS 0.008123f
C692 B.n540 VSUBS 0.008123f
C693 B.n541 VSUBS 0.008123f
C694 B.n542 VSUBS 0.008123f
C695 B.n543 VSUBS 0.008123f
C696 B.n544 VSUBS 0.008123f
C697 B.n545 VSUBS 0.008123f
C698 B.n546 VSUBS 0.008123f
C699 B.n547 VSUBS 0.008123f
C700 B.n548 VSUBS 0.008123f
C701 B.n549 VSUBS 0.008123f
C702 B.n550 VSUBS 0.008123f
C703 B.n551 VSUBS 0.008123f
C704 B.n552 VSUBS 0.008123f
C705 B.n553 VSUBS 0.008123f
C706 B.n554 VSUBS 0.008123f
C707 B.n555 VSUBS 0.008123f
C708 B.n556 VSUBS 0.008123f
C709 B.n557 VSUBS 0.008123f
C710 B.n558 VSUBS 0.008123f
C711 B.n559 VSUBS 0.008123f
C712 B.n560 VSUBS 0.008123f
C713 B.n561 VSUBS 0.008123f
C714 B.n562 VSUBS 0.008123f
C715 B.n563 VSUBS 0.008123f
C716 B.n564 VSUBS 0.008123f
C717 B.n565 VSUBS 0.008123f
C718 B.n566 VSUBS 0.008123f
C719 B.n567 VSUBS 0.008123f
C720 B.n568 VSUBS 0.008123f
C721 B.n569 VSUBS 0.008123f
C722 B.n570 VSUBS 0.008123f
C723 B.n571 VSUBS 0.008123f
C724 B.n572 VSUBS 0.008123f
C725 B.n573 VSUBS 0.008123f
C726 B.n574 VSUBS 0.008123f
C727 B.n575 VSUBS 0.008123f
C728 B.n576 VSUBS 0.008123f
C729 B.n577 VSUBS 0.008123f
C730 B.n578 VSUBS 0.008123f
C731 B.n579 VSUBS 0.008123f
C732 B.n580 VSUBS 0.008123f
C733 B.n581 VSUBS 0.008123f
C734 B.n582 VSUBS 0.008123f
C735 B.n583 VSUBS 0.008123f
C736 B.n584 VSUBS 0.008123f
C737 B.n585 VSUBS 0.008123f
C738 B.n586 VSUBS 0.008123f
C739 B.n587 VSUBS 0.008123f
C740 B.n588 VSUBS 0.008123f
C741 B.n589 VSUBS 0.008123f
C742 B.n590 VSUBS 0.008123f
C743 B.n591 VSUBS 0.008123f
C744 B.n592 VSUBS 0.008123f
C745 B.n593 VSUBS 0.008123f
C746 B.n594 VSUBS 0.008123f
C747 B.n595 VSUBS 0.008123f
C748 B.n596 VSUBS 0.008123f
C749 B.n597 VSUBS 0.008123f
C750 B.n598 VSUBS 0.008123f
C751 B.n599 VSUBS 0.008123f
C752 B.n600 VSUBS 0.008123f
C753 B.n601 VSUBS 0.008123f
C754 B.n602 VSUBS 0.008123f
C755 B.n603 VSUBS 0.008123f
C756 B.n604 VSUBS 0.008123f
C757 B.n605 VSUBS 0.008123f
C758 B.n606 VSUBS 0.008123f
C759 B.n607 VSUBS 0.008123f
C760 B.n608 VSUBS 0.008123f
C761 B.n609 VSUBS 0.008123f
C762 B.n610 VSUBS 0.008123f
C763 B.n611 VSUBS 0.008123f
C764 B.n612 VSUBS 0.008123f
C765 B.n613 VSUBS 0.008123f
C766 B.n614 VSUBS 0.008123f
C767 B.n615 VSUBS 0.008123f
C768 B.n616 VSUBS 0.008123f
C769 B.n617 VSUBS 0.008123f
C770 B.n618 VSUBS 0.008123f
C771 B.n619 VSUBS 0.008123f
C772 B.n620 VSUBS 0.008123f
C773 B.n621 VSUBS 0.008123f
C774 B.n622 VSUBS 0.008123f
C775 B.n623 VSUBS 0.008123f
C776 B.n624 VSUBS 0.008123f
C777 B.n625 VSUBS 0.008123f
C778 B.n626 VSUBS 0.008123f
C779 B.n627 VSUBS 0.008123f
C780 B.n628 VSUBS 0.008123f
C781 B.n629 VSUBS 0.008123f
C782 B.n630 VSUBS 0.008123f
C783 B.n631 VSUBS 0.008123f
C784 B.n632 VSUBS 0.008123f
C785 B.n633 VSUBS 0.008123f
C786 B.n634 VSUBS 0.008123f
C787 B.n635 VSUBS 0.008123f
C788 B.n636 VSUBS 0.008123f
C789 B.n637 VSUBS 0.008123f
C790 B.n638 VSUBS 0.008123f
C791 B.n639 VSUBS 0.008123f
C792 B.n640 VSUBS 0.008123f
C793 B.n641 VSUBS 0.008123f
C794 B.n642 VSUBS 0.008123f
C795 B.n643 VSUBS 0.008123f
C796 B.n644 VSUBS 0.008123f
C797 B.n645 VSUBS 0.008123f
C798 B.n646 VSUBS 0.008123f
C799 B.n647 VSUBS 0.008123f
C800 B.n648 VSUBS 0.008123f
C801 B.n649 VSUBS 0.008123f
C802 B.n650 VSUBS 0.008123f
C803 B.n651 VSUBS 0.008123f
C804 B.n652 VSUBS 0.008123f
C805 B.n653 VSUBS 0.008123f
C806 B.n654 VSUBS 0.008123f
C807 B.n655 VSUBS 0.008123f
C808 B.n656 VSUBS 0.008123f
C809 B.n657 VSUBS 0.008123f
C810 B.n658 VSUBS 0.008123f
C811 B.n659 VSUBS 0.008123f
C812 B.n660 VSUBS 0.008123f
C813 B.n661 VSUBS 0.008123f
C814 B.n662 VSUBS 0.008123f
C815 B.n663 VSUBS 0.008123f
C816 B.n664 VSUBS 0.008123f
C817 B.n665 VSUBS 0.008123f
C818 B.n666 VSUBS 0.008123f
C819 B.n667 VSUBS 0.008123f
C820 B.n668 VSUBS 0.008123f
C821 B.n669 VSUBS 0.008123f
C822 B.n670 VSUBS 0.008123f
C823 B.n671 VSUBS 0.008123f
C824 B.n672 VSUBS 0.008123f
C825 B.n673 VSUBS 0.008123f
C826 B.n674 VSUBS 0.008123f
C827 B.n675 VSUBS 0.008123f
C828 B.n676 VSUBS 0.008123f
C829 B.n677 VSUBS 0.008123f
C830 B.n678 VSUBS 0.008123f
C831 B.n679 VSUBS 0.008123f
C832 B.n680 VSUBS 0.008123f
C833 B.n681 VSUBS 0.008123f
C834 B.n682 VSUBS 0.008123f
C835 B.n683 VSUBS 0.008123f
C836 B.n684 VSUBS 0.008123f
C837 B.n685 VSUBS 0.008123f
C838 B.n686 VSUBS 0.008123f
C839 B.n687 VSUBS 0.008123f
C840 B.n688 VSUBS 0.008123f
C841 B.n689 VSUBS 0.008123f
C842 B.n690 VSUBS 0.008123f
C843 B.n691 VSUBS 0.008123f
C844 B.n692 VSUBS 0.008123f
C845 B.n693 VSUBS 0.008123f
C846 B.n694 VSUBS 0.008123f
C847 B.n695 VSUBS 0.008123f
C848 B.n696 VSUBS 0.008123f
C849 B.n697 VSUBS 0.008123f
C850 B.n698 VSUBS 0.008123f
C851 B.n699 VSUBS 0.008123f
C852 B.n700 VSUBS 0.008123f
C853 B.n701 VSUBS 0.008123f
C854 B.n702 VSUBS 0.008123f
C855 B.n703 VSUBS 0.008123f
C856 B.n704 VSUBS 0.008123f
C857 B.n705 VSUBS 0.008123f
C858 B.n706 VSUBS 0.008123f
C859 B.n707 VSUBS 0.008123f
C860 B.n708 VSUBS 0.008123f
C861 B.n709 VSUBS 0.008123f
C862 B.n710 VSUBS 0.008123f
C863 B.n711 VSUBS 0.008123f
C864 B.n712 VSUBS 0.008123f
C865 B.n713 VSUBS 0.008123f
C866 B.n714 VSUBS 0.008123f
C867 B.n715 VSUBS 0.008123f
C868 B.n716 VSUBS 0.018697f
C869 B.n717 VSUBS 0.019667f
C870 B.n718 VSUBS 0.018082f
C871 B.n719 VSUBS 0.008123f
C872 B.n720 VSUBS 0.008123f
C873 B.n721 VSUBS 0.008123f
C874 B.n722 VSUBS 0.008123f
C875 B.n723 VSUBS 0.008123f
C876 B.n724 VSUBS 0.008123f
C877 B.n725 VSUBS 0.008123f
C878 B.n726 VSUBS 0.008123f
C879 B.n727 VSUBS 0.008123f
C880 B.n728 VSUBS 0.008123f
C881 B.n729 VSUBS 0.008123f
C882 B.n730 VSUBS 0.008123f
C883 B.n731 VSUBS 0.008123f
C884 B.n732 VSUBS 0.008123f
C885 B.n733 VSUBS 0.008123f
C886 B.n734 VSUBS 0.008123f
C887 B.n735 VSUBS 0.008123f
C888 B.n736 VSUBS 0.008123f
C889 B.n737 VSUBS 0.008123f
C890 B.n738 VSUBS 0.008123f
C891 B.n739 VSUBS 0.008123f
C892 B.n740 VSUBS 0.008123f
C893 B.n741 VSUBS 0.008123f
C894 B.n742 VSUBS 0.008123f
C895 B.n743 VSUBS 0.008123f
C896 B.n744 VSUBS 0.008123f
C897 B.n745 VSUBS 0.008123f
C898 B.n746 VSUBS 0.008123f
C899 B.n747 VSUBS 0.008123f
C900 B.n748 VSUBS 0.008123f
C901 B.n749 VSUBS 0.008123f
C902 B.n750 VSUBS 0.008123f
C903 B.n751 VSUBS 0.008123f
C904 B.n752 VSUBS 0.008123f
C905 B.n753 VSUBS 0.008123f
C906 B.n754 VSUBS 0.008123f
C907 B.n755 VSUBS 0.008123f
C908 B.n756 VSUBS 0.008123f
C909 B.n757 VSUBS 0.008123f
C910 B.n758 VSUBS 0.008123f
C911 B.n759 VSUBS 0.008123f
C912 B.n760 VSUBS 0.008123f
C913 B.n761 VSUBS 0.008123f
C914 B.n762 VSUBS 0.008123f
C915 B.n763 VSUBS 0.008123f
C916 B.n764 VSUBS 0.008123f
C917 B.n765 VSUBS 0.008123f
C918 B.n766 VSUBS 0.008123f
C919 B.n767 VSUBS 0.008123f
C920 B.n768 VSUBS 0.008123f
C921 B.n769 VSUBS 0.008123f
C922 B.n770 VSUBS 0.008123f
C923 B.n771 VSUBS 0.008123f
C924 B.n772 VSUBS 0.008123f
C925 B.n773 VSUBS 0.008123f
C926 B.n774 VSUBS 0.008123f
C927 B.n775 VSUBS 0.008123f
C928 B.n776 VSUBS 0.008123f
C929 B.n777 VSUBS 0.008123f
C930 B.n778 VSUBS 0.008123f
C931 B.n779 VSUBS 0.008123f
C932 B.n780 VSUBS 0.008123f
C933 B.n781 VSUBS 0.008123f
C934 B.n782 VSUBS 0.008123f
C935 B.n783 VSUBS 0.008123f
C936 B.n784 VSUBS 0.008123f
C937 B.n785 VSUBS 0.008123f
C938 B.n786 VSUBS 0.008123f
C939 B.n787 VSUBS 0.008123f
C940 B.n788 VSUBS 0.008123f
C941 B.n789 VSUBS 0.008123f
C942 B.n790 VSUBS 0.008123f
C943 B.n791 VSUBS 0.008123f
C944 B.n792 VSUBS 0.008123f
C945 B.n793 VSUBS 0.008123f
C946 B.n794 VSUBS 0.008123f
C947 B.n795 VSUBS 0.008123f
C948 B.n796 VSUBS 0.008123f
C949 B.n797 VSUBS 0.008123f
C950 B.n798 VSUBS 0.008123f
C951 B.n799 VSUBS 0.008123f
C952 B.n800 VSUBS 0.008123f
C953 B.n801 VSUBS 0.008123f
C954 B.n802 VSUBS 0.008123f
C955 B.n803 VSUBS 0.007645f
C956 B.n804 VSUBS 0.008123f
C957 B.n805 VSUBS 0.008123f
C958 B.n806 VSUBS 0.004539f
C959 B.n807 VSUBS 0.008123f
C960 B.n808 VSUBS 0.008123f
C961 B.n809 VSUBS 0.008123f
C962 B.n810 VSUBS 0.008123f
C963 B.n811 VSUBS 0.008123f
C964 B.n812 VSUBS 0.008123f
C965 B.n813 VSUBS 0.008123f
C966 B.n814 VSUBS 0.008123f
C967 B.n815 VSUBS 0.008123f
C968 B.n816 VSUBS 0.008123f
C969 B.n817 VSUBS 0.008123f
C970 B.n818 VSUBS 0.008123f
C971 B.n819 VSUBS 0.004539f
C972 B.n820 VSUBS 0.018821f
C973 B.n821 VSUBS 0.007645f
C974 B.n822 VSUBS 0.008123f
C975 B.n823 VSUBS 0.008123f
C976 B.n824 VSUBS 0.008123f
C977 B.n825 VSUBS 0.008123f
C978 B.n826 VSUBS 0.008123f
C979 B.n827 VSUBS 0.008123f
C980 B.n828 VSUBS 0.008123f
C981 B.n829 VSUBS 0.008123f
C982 B.n830 VSUBS 0.008123f
C983 B.n831 VSUBS 0.008123f
C984 B.n832 VSUBS 0.008123f
C985 B.n833 VSUBS 0.008123f
C986 B.n834 VSUBS 0.008123f
C987 B.n835 VSUBS 0.008123f
C988 B.n836 VSUBS 0.008123f
C989 B.n837 VSUBS 0.008123f
C990 B.n838 VSUBS 0.008123f
C991 B.n839 VSUBS 0.008123f
C992 B.n840 VSUBS 0.008123f
C993 B.n841 VSUBS 0.008123f
C994 B.n842 VSUBS 0.008123f
C995 B.n843 VSUBS 0.008123f
C996 B.n844 VSUBS 0.008123f
C997 B.n845 VSUBS 0.008123f
C998 B.n846 VSUBS 0.008123f
C999 B.n847 VSUBS 0.008123f
C1000 B.n848 VSUBS 0.008123f
C1001 B.n849 VSUBS 0.008123f
C1002 B.n850 VSUBS 0.008123f
C1003 B.n851 VSUBS 0.008123f
C1004 B.n852 VSUBS 0.008123f
C1005 B.n853 VSUBS 0.008123f
C1006 B.n854 VSUBS 0.008123f
C1007 B.n855 VSUBS 0.008123f
C1008 B.n856 VSUBS 0.008123f
C1009 B.n857 VSUBS 0.008123f
C1010 B.n858 VSUBS 0.008123f
C1011 B.n859 VSUBS 0.008123f
C1012 B.n860 VSUBS 0.008123f
C1013 B.n861 VSUBS 0.008123f
C1014 B.n862 VSUBS 0.008123f
C1015 B.n863 VSUBS 0.008123f
C1016 B.n864 VSUBS 0.008123f
C1017 B.n865 VSUBS 0.008123f
C1018 B.n866 VSUBS 0.008123f
C1019 B.n867 VSUBS 0.008123f
C1020 B.n868 VSUBS 0.008123f
C1021 B.n869 VSUBS 0.008123f
C1022 B.n870 VSUBS 0.008123f
C1023 B.n871 VSUBS 0.008123f
C1024 B.n872 VSUBS 0.008123f
C1025 B.n873 VSUBS 0.008123f
C1026 B.n874 VSUBS 0.008123f
C1027 B.n875 VSUBS 0.008123f
C1028 B.n876 VSUBS 0.008123f
C1029 B.n877 VSUBS 0.008123f
C1030 B.n878 VSUBS 0.008123f
C1031 B.n879 VSUBS 0.008123f
C1032 B.n880 VSUBS 0.008123f
C1033 B.n881 VSUBS 0.008123f
C1034 B.n882 VSUBS 0.008123f
C1035 B.n883 VSUBS 0.008123f
C1036 B.n884 VSUBS 0.008123f
C1037 B.n885 VSUBS 0.008123f
C1038 B.n886 VSUBS 0.008123f
C1039 B.n887 VSUBS 0.008123f
C1040 B.n888 VSUBS 0.008123f
C1041 B.n889 VSUBS 0.008123f
C1042 B.n890 VSUBS 0.008123f
C1043 B.n891 VSUBS 0.008123f
C1044 B.n892 VSUBS 0.008123f
C1045 B.n893 VSUBS 0.008123f
C1046 B.n894 VSUBS 0.008123f
C1047 B.n895 VSUBS 0.008123f
C1048 B.n896 VSUBS 0.008123f
C1049 B.n897 VSUBS 0.008123f
C1050 B.n898 VSUBS 0.008123f
C1051 B.n899 VSUBS 0.008123f
C1052 B.n900 VSUBS 0.008123f
C1053 B.n901 VSUBS 0.008123f
C1054 B.n902 VSUBS 0.008123f
C1055 B.n903 VSUBS 0.008123f
C1056 B.n904 VSUBS 0.008123f
C1057 B.n905 VSUBS 0.008123f
C1058 B.n906 VSUBS 0.008123f
C1059 B.n907 VSUBS 0.019052f
C1060 B.n908 VSUBS 0.018697f
C1061 B.n909 VSUBS 0.018697f
C1062 B.n910 VSUBS 0.008123f
C1063 B.n911 VSUBS 0.008123f
C1064 B.n912 VSUBS 0.008123f
C1065 B.n913 VSUBS 0.008123f
C1066 B.n914 VSUBS 0.008123f
C1067 B.n915 VSUBS 0.008123f
C1068 B.n916 VSUBS 0.008123f
C1069 B.n917 VSUBS 0.008123f
C1070 B.n918 VSUBS 0.008123f
C1071 B.n919 VSUBS 0.008123f
C1072 B.n920 VSUBS 0.008123f
C1073 B.n921 VSUBS 0.008123f
C1074 B.n922 VSUBS 0.008123f
C1075 B.n923 VSUBS 0.008123f
C1076 B.n924 VSUBS 0.008123f
C1077 B.n925 VSUBS 0.008123f
C1078 B.n926 VSUBS 0.008123f
C1079 B.n927 VSUBS 0.008123f
C1080 B.n928 VSUBS 0.008123f
C1081 B.n929 VSUBS 0.008123f
C1082 B.n930 VSUBS 0.008123f
C1083 B.n931 VSUBS 0.008123f
C1084 B.n932 VSUBS 0.008123f
C1085 B.n933 VSUBS 0.008123f
C1086 B.n934 VSUBS 0.008123f
C1087 B.n935 VSUBS 0.008123f
C1088 B.n936 VSUBS 0.008123f
C1089 B.n937 VSUBS 0.008123f
C1090 B.n938 VSUBS 0.008123f
C1091 B.n939 VSUBS 0.008123f
C1092 B.n940 VSUBS 0.008123f
C1093 B.n941 VSUBS 0.008123f
C1094 B.n942 VSUBS 0.008123f
C1095 B.n943 VSUBS 0.008123f
C1096 B.n944 VSUBS 0.008123f
C1097 B.n945 VSUBS 0.008123f
C1098 B.n946 VSUBS 0.008123f
C1099 B.n947 VSUBS 0.008123f
C1100 B.n948 VSUBS 0.008123f
C1101 B.n949 VSUBS 0.008123f
C1102 B.n950 VSUBS 0.008123f
C1103 B.n951 VSUBS 0.008123f
C1104 B.n952 VSUBS 0.008123f
C1105 B.n953 VSUBS 0.008123f
C1106 B.n954 VSUBS 0.008123f
C1107 B.n955 VSUBS 0.008123f
C1108 B.n956 VSUBS 0.008123f
C1109 B.n957 VSUBS 0.008123f
C1110 B.n958 VSUBS 0.008123f
C1111 B.n959 VSUBS 0.008123f
C1112 B.n960 VSUBS 0.008123f
C1113 B.n961 VSUBS 0.008123f
C1114 B.n962 VSUBS 0.008123f
C1115 B.n963 VSUBS 0.008123f
C1116 B.n964 VSUBS 0.008123f
C1117 B.n965 VSUBS 0.008123f
C1118 B.n966 VSUBS 0.008123f
C1119 B.n967 VSUBS 0.008123f
C1120 B.n968 VSUBS 0.008123f
C1121 B.n969 VSUBS 0.008123f
C1122 B.n970 VSUBS 0.008123f
C1123 B.n971 VSUBS 0.008123f
C1124 B.n972 VSUBS 0.008123f
C1125 B.n973 VSUBS 0.008123f
C1126 B.n974 VSUBS 0.008123f
C1127 B.n975 VSUBS 0.008123f
C1128 B.n976 VSUBS 0.008123f
C1129 B.n977 VSUBS 0.008123f
C1130 B.n978 VSUBS 0.008123f
C1131 B.n979 VSUBS 0.008123f
C1132 B.n980 VSUBS 0.008123f
C1133 B.n981 VSUBS 0.008123f
C1134 B.n982 VSUBS 0.008123f
C1135 B.n983 VSUBS 0.008123f
C1136 B.n984 VSUBS 0.008123f
C1137 B.n985 VSUBS 0.008123f
C1138 B.n986 VSUBS 0.008123f
C1139 B.n987 VSUBS 0.008123f
C1140 B.n988 VSUBS 0.008123f
C1141 B.n989 VSUBS 0.008123f
C1142 B.n990 VSUBS 0.008123f
C1143 B.n991 VSUBS 0.008123f
C1144 B.n992 VSUBS 0.008123f
C1145 B.n993 VSUBS 0.008123f
C1146 B.n994 VSUBS 0.008123f
C1147 B.n995 VSUBS 0.008123f
C1148 B.n996 VSUBS 0.008123f
C1149 B.n997 VSUBS 0.008123f
C1150 B.n998 VSUBS 0.008123f
C1151 B.n999 VSUBS 0.018394f
C1152 VTAIL.t5 VSUBS 0.383488f
C1153 VTAIL.t8 VSUBS 0.383488f
C1154 VTAIL.n0 VSUBS 3.05125f
C1155 VTAIL.n1 VSUBS 0.955776f
C1156 VTAIL.t10 VSUBS 3.97773f
C1157 VTAIL.n2 VSUBS 1.12582f
C1158 VTAIL.t13 VSUBS 0.383488f
C1159 VTAIL.t18 VSUBS 0.383488f
C1160 VTAIL.n3 VSUBS 3.05125f
C1161 VTAIL.n4 VSUBS 1.07649f
C1162 VTAIL.t16 VSUBS 0.383488f
C1163 VTAIL.t14 VSUBS 0.383488f
C1164 VTAIL.n5 VSUBS 3.05125f
C1165 VTAIL.n6 VSUBS 3.02009f
C1166 VTAIL.t4 VSUBS 0.383488f
C1167 VTAIL.t1 VSUBS 0.383488f
C1168 VTAIL.n7 VSUBS 3.05124f
C1169 VTAIL.n8 VSUBS 3.02009f
C1170 VTAIL.t7 VSUBS 0.383488f
C1171 VTAIL.t9 VSUBS 0.383488f
C1172 VTAIL.n9 VSUBS 3.05124f
C1173 VTAIL.n10 VSUBS 1.07649f
C1174 VTAIL.t2 VSUBS 3.97774f
C1175 VTAIL.n11 VSUBS 1.12581f
C1176 VTAIL.t15 VSUBS 0.383488f
C1177 VTAIL.t19 VSUBS 0.383488f
C1178 VTAIL.n12 VSUBS 3.05124f
C1179 VTAIL.n13 VSUBS 1.00643f
C1180 VTAIL.t12 VSUBS 0.383488f
C1181 VTAIL.t17 VSUBS 0.383488f
C1182 VTAIL.n14 VSUBS 3.05124f
C1183 VTAIL.n15 VSUBS 1.07649f
C1184 VTAIL.t11 VSUBS 3.97771f
C1185 VTAIL.n16 VSUBS 2.91635f
C1186 VTAIL.t6 VSUBS 3.97773f
C1187 VTAIL.n17 VSUBS 2.91634f
C1188 VTAIL.t3 VSUBS 0.383488f
C1189 VTAIL.t0 VSUBS 0.383488f
C1190 VTAIL.n18 VSUBS 3.05125f
C1191 VTAIL.n19 VSUBS 0.903988f
C1192 VDD1.t7 VSUBS 4.32646f
C1193 VDD1.t3 VSUBS 0.396704f
C1194 VDD1.t8 VSUBS 0.396704f
C1195 VDD1.n0 VSUBS 3.31517f
C1196 VDD1.n1 VSUBS 1.67015f
C1197 VDD1.t0 VSUBS 4.32645f
C1198 VDD1.t6 VSUBS 0.396704f
C1199 VDD1.t9 VSUBS 0.396704f
C1200 VDD1.n2 VSUBS 3.31518f
C1201 VDD1.n3 VSUBS 1.66091f
C1202 VDD1.t2 VSUBS 0.396704f
C1203 VDD1.t4 VSUBS 0.396704f
C1204 VDD1.n4 VSUBS 3.33866f
C1205 VDD1.n5 VSUBS 4.13981f
C1206 VDD1.t1 VSUBS 0.396704f
C1207 VDD1.t5 VSUBS 0.396704f
C1208 VDD1.n6 VSUBS 3.31516f
C1209 VDD1.n7 VSUBS 4.38759f
C1210 VP.n0 VSUBS 0.035779f
C1211 VP.t9 VSUBS 3.43434f
C1212 VP.n1 VSUBS 0.04705f
C1213 VP.n2 VSUBS 0.02714f
C1214 VP.t1 VSUBS 3.43434f
C1215 VP.n3 VSUBS 1.1916f
C1216 VP.n4 VSUBS 0.02714f
C1217 VP.n5 VSUBS 0.036824f
C1218 VP.n6 VSUBS 0.02714f
C1219 VP.t6 VSUBS 3.43434f
C1220 VP.n7 VSUBS 0.050329f
C1221 VP.n8 VSUBS 0.02714f
C1222 VP.n9 VSUBS 0.034427f
C1223 VP.n10 VSUBS 0.02714f
C1224 VP.n11 VSUBS 0.04705f
C1225 VP.n12 VSUBS 0.035779f
C1226 VP.t3 VSUBS 3.43434f
C1227 VP.n13 VSUBS 0.035779f
C1228 VP.t8 VSUBS 3.43434f
C1229 VP.n14 VSUBS 0.04705f
C1230 VP.n15 VSUBS 0.02714f
C1231 VP.t2 VSUBS 3.43434f
C1232 VP.n16 VSUBS 1.1916f
C1233 VP.n17 VSUBS 0.02714f
C1234 VP.n18 VSUBS 0.036824f
C1235 VP.n19 VSUBS 0.02714f
C1236 VP.t7 VSUBS 3.43434f
C1237 VP.n20 VSUBS 0.050329f
C1238 VP.n21 VSUBS 0.02714f
C1239 VP.n22 VSUBS 0.034427f
C1240 VP.t4 VSUBS 3.65709f
C1241 VP.t0 VSUBS 3.43434f
C1242 VP.n23 VSUBS 1.26615f
C1243 VP.n24 VSUBS 1.24491f
C1244 VP.n25 VSUBS 0.261993f
C1245 VP.n26 VSUBS 0.02714f
C1246 VP.n27 VSUBS 0.050329f
C1247 VP.n28 VSUBS 0.042081f
C1248 VP.n29 VSUBS 0.036824f
C1249 VP.n30 VSUBS 0.02714f
C1250 VP.n31 VSUBS 0.02714f
C1251 VP.n32 VSUBS 0.02714f
C1252 VP.n33 VSUBS 0.037906f
C1253 VP.n34 VSUBS 1.1916f
C1254 VP.n35 VSUBS 0.037906f
C1255 VP.n36 VSUBS 0.050329f
C1256 VP.n37 VSUBS 0.02714f
C1257 VP.n38 VSUBS 0.02714f
C1258 VP.n39 VSUBS 0.02714f
C1259 VP.n40 VSUBS 0.042081f
C1260 VP.n41 VSUBS 0.050329f
C1261 VP.n42 VSUBS 0.034427f
C1262 VP.n43 VSUBS 0.02714f
C1263 VP.n44 VSUBS 0.02714f
C1264 VP.n45 VSUBS 0.041384f
C1265 VP.n46 VSUBS 0.051998f
C1266 VP.n47 VSUBS 0.030185f
C1267 VP.n48 VSUBS 0.02714f
C1268 VP.n49 VSUBS 0.02714f
C1269 VP.n50 VSUBS 0.02714f
C1270 VP.n51 VSUBS 0.050329f
C1271 VP.n52 VSUBS 0.030949f
C1272 VP.n53 VSUBS 1.27532f
C1273 VP.n54 VSUBS 1.83974f
C1274 VP.n55 VSUBS 1.85679f
C1275 VP.n56 VSUBS 1.27532f
C1276 VP.n57 VSUBS 0.030949f
C1277 VP.n58 VSUBS 0.050329f
C1278 VP.n59 VSUBS 0.02714f
C1279 VP.n60 VSUBS 0.02714f
C1280 VP.n61 VSUBS 0.02714f
C1281 VP.n62 VSUBS 0.030185f
C1282 VP.n63 VSUBS 0.051998f
C1283 VP.t5 VSUBS 3.43434f
C1284 VP.n64 VSUBS 1.1916f
C1285 VP.n65 VSUBS 0.041384f
C1286 VP.n66 VSUBS 0.02714f
C1287 VP.n67 VSUBS 0.02714f
C1288 VP.n68 VSUBS 0.02714f
C1289 VP.n69 VSUBS 0.050329f
C1290 VP.n70 VSUBS 0.042081f
C1291 VP.n71 VSUBS 0.036824f
C1292 VP.n72 VSUBS 0.02714f
C1293 VP.n73 VSUBS 0.02714f
C1294 VP.n74 VSUBS 0.02714f
C1295 VP.n75 VSUBS 0.037906f
C1296 VP.n76 VSUBS 1.1916f
C1297 VP.n77 VSUBS 0.037906f
C1298 VP.n78 VSUBS 0.050329f
C1299 VP.n79 VSUBS 0.02714f
C1300 VP.n80 VSUBS 0.02714f
C1301 VP.n81 VSUBS 0.02714f
C1302 VP.n82 VSUBS 0.042081f
C1303 VP.n83 VSUBS 0.050329f
C1304 VP.n84 VSUBS 0.034427f
C1305 VP.n85 VSUBS 0.02714f
C1306 VP.n86 VSUBS 0.02714f
C1307 VP.n87 VSUBS 0.041384f
C1308 VP.n88 VSUBS 0.051998f
C1309 VP.n89 VSUBS 0.030185f
C1310 VP.n90 VSUBS 0.02714f
C1311 VP.n91 VSUBS 0.02714f
C1312 VP.n92 VSUBS 0.02714f
C1313 VP.n93 VSUBS 0.050329f
C1314 VP.n94 VSUBS 0.030949f
C1315 VP.n95 VSUBS 1.27532f
C1316 VP.n96 VSUBS 0.047066f
.ends

