* NGSPICE file created from diff_pair_sample_1387.ext - technology: sky130A

.subckt diff_pair_sample_1387 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t13 w_n3970_n3374# sky130_fd_pr__pfet_01v8 ad=1.98495 pd=12.36 as=4.6917 ps=24.84 w=12.03 l=2.67
X1 VTAIL.t14 VP.t1 VDD1.t6 w_n3970_n3374# sky130_fd_pr__pfet_01v8 ad=1.98495 pd=12.36 as=1.98495 ps=12.36 w=12.03 l=2.67
X2 VDD2.t7 VN.t0 VTAIL.t1 w_n3970_n3374# sky130_fd_pr__pfet_01v8 ad=1.98495 pd=12.36 as=1.98495 ps=12.36 w=12.03 l=2.67
X3 VTAIL.t2 VN.t1 VDD2.t6 w_n3970_n3374# sky130_fd_pr__pfet_01v8 ad=4.6917 pd=24.84 as=1.98495 ps=12.36 w=12.03 l=2.67
X4 B.t11 B.t9 B.t10 w_n3970_n3374# sky130_fd_pr__pfet_01v8 ad=4.6917 pd=24.84 as=0 ps=0 w=12.03 l=2.67
X5 B.t8 B.t6 B.t7 w_n3970_n3374# sky130_fd_pr__pfet_01v8 ad=4.6917 pd=24.84 as=0 ps=0 w=12.03 l=2.67
X6 VTAIL.t9 VP.t2 VDD1.t5 w_n3970_n3374# sky130_fd_pr__pfet_01v8 ad=1.98495 pd=12.36 as=1.98495 ps=12.36 w=12.03 l=2.67
X7 VDD2.t5 VN.t2 VTAIL.t3 w_n3970_n3374# sky130_fd_pr__pfet_01v8 ad=1.98495 pd=12.36 as=4.6917 ps=24.84 w=12.03 l=2.67
X8 VDD1.t4 VP.t3 VTAIL.t15 w_n3970_n3374# sky130_fd_pr__pfet_01v8 ad=1.98495 pd=12.36 as=1.98495 ps=12.36 w=12.03 l=2.67
X9 B.t5 B.t3 B.t4 w_n3970_n3374# sky130_fd_pr__pfet_01v8 ad=4.6917 pd=24.84 as=0 ps=0 w=12.03 l=2.67
X10 VTAIL.t5 VN.t3 VDD2.t4 w_n3970_n3374# sky130_fd_pr__pfet_01v8 ad=1.98495 pd=12.36 as=1.98495 ps=12.36 w=12.03 l=2.67
X11 B.t2 B.t0 B.t1 w_n3970_n3374# sky130_fd_pr__pfet_01v8 ad=4.6917 pd=24.84 as=0 ps=0 w=12.03 l=2.67
X12 VTAIL.t7 VN.t4 VDD2.t3 w_n3970_n3374# sky130_fd_pr__pfet_01v8 ad=1.98495 pd=12.36 as=1.98495 ps=12.36 w=12.03 l=2.67
X13 VTAIL.t0 VN.t5 VDD2.t2 w_n3970_n3374# sky130_fd_pr__pfet_01v8 ad=4.6917 pd=24.84 as=1.98495 ps=12.36 w=12.03 l=2.67
X14 VTAIL.t11 VP.t4 VDD1.t3 w_n3970_n3374# sky130_fd_pr__pfet_01v8 ad=4.6917 pd=24.84 as=1.98495 ps=12.36 w=12.03 l=2.67
X15 VDD1.t2 VP.t5 VTAIL.t10 w_n3970_n3374# sky130_fd_pr__pfet_01v8 ad=1.98495 pd=12.36 as=4.6917 ps=24.84 w=12.03 l=2.67
X16 VDD1.t1 VP.t6 VTAIL.t8 w_n3970_n3374# sky130_fd_pr__pfet_01v8 ad=1.98495 pd=12.36 as=1.98495 ps=12.36 w=12.03 l=2.67
X17 VDD2.t1 VN.t6 VTAIL.t6 w_n3970_n3374# sky130_fd_pr__pfet_01v8 ad=1.98495 pd=12.36 as=4.6917 ps=24.84 w=12.03 l=2.67
X18 VDD2.t0 VN.t7 VTAIL.t4 w_n3970_n3374# sky130_fd_pr__pfet_01v8 ad=1.98495 pd=12.36 as=1.98495 ps=12.36 w=12.03 l=2.67
X19 VTAIL.t12 VP.t7 VDD1.t0 w_n3970_n3374# sky130_fd_pr__pfet_01v8 ad=4.6917 pd=24.84 as=1.98495 ps=12.36 w=12.03 l=2.67
R0 VP.n18 VP.n17 161.3
R1 VP.n19 VP.n14 161.3
R2 VP.n21 VP.n20 161.3
R3 VP.n22 VP.n13 161.3
R4 VP.n24 VP.n23 161.3
R5 VP.n25 VP.n12 161.3
R6 VP.n27 VP.n26 161.3
R7 VP.n28 VP.n11 161.3
R8 VP.n30 VP.n29 161.3
R9 VP.n31 VP.n10 161.3
R10 VP.n33 VP.n32 161.3
R11 VP.n62 VP.n61 161.3
R12 VP.n60 VP.n1 161.3
R13 VP.n59 VP.n58 161.3
R14 VP.n57 VP.n2 161.3
R15 VP.n56 VP.n55 161.3
R16 VP.n54 VP.n3 161.3
R17 VP.n53 VP.n52 161.3
R18 VP.n51 VP.n4 161.3
R19 VP.n50 VP.n49 161.3
R20 VP.n48 VP.n5 161.3
R21 VP.n47 VP.n46 161.3
R22 VP.n45 VP.n6 161.3
R23 VP.n44 VP.n43 161.3
R24 VP.n42 VP.n7 161.3
R25 VP.n41 VP.n40 161.3
R26 VP.n39 VP.n8 161.3
R27 VP.n38 VP.n37 161.3
R28 VP.n16 VP.t4 140.736
R29 VP.n0 VP.t5 108.585
R30 VP.n54 VP.t2 108.585
R31 VP.n6 VP.t3 108.585
R32 VP.n36 VP.t7 108.585
R33 VP.n15 VP.t6 108.585
R34 VP.n25 VP.t1 108.585
R35 VP.n9 VP.t0 108.585
R36 VP.n34 VP.n9 65.6004
R37 VP.n63 VP.n0 65.6004
R38 VP.n36 VP.n35 65.6004
R39 VP.n35 VP.n34 51.3554
R40 VP.n16 VP.n15 48.9289
R41 VP.n41 VP.n8 40.4934
R42 VP.n42 VP.n41 40.4934
R43 VP.n49 VP.n48 40.4934
R44 VP.n49 VP.n4 40.4934
R45 VP.n59 VP.n2 40.4934
R46 VP.n60 VP.n59 40.4934
R47 VP.n31 VP.n30 40.4934
R48 VP.n30 VP.n11 40.4934
R49 VP.n20 VP.n13 40.4934
R50 VP.n20 VP.n19 40.4934
R51 VP.n37 VP.n36 24.4675
R52 VP.n37 VP.n8 24.4675
R53 VP.n43 VP.n42 24.4675
R54 VP.n43 VP.n6 24.4675
R55 VP.n47 VP.n6 24.4675
R56 VP.n48 VP.n47 24.4675
R57 VP.n53 VP.n4 24.4675
R58 VP.n54 VP.n53 24.4675
R59 VP.n55 VP.n54 24.4675
R60 VP.n55 VP.n2 24.4675
R61 VP.n61 VP.n60 24.4675
R62 VP.n61 VP.n0 24.4675
R63 VP.n32 VP.n31 24.4675
R64 VP.n32 VP.n9 24.4675
R65 VP.n24 VP.n13 24.4675
R66 VP.n25 VP.n24 24.4675
R67 VP.n26 VP.n25 24.4675
R68 VP.n26 VP.n11 24.4675
R69 VP.n18 VP.n15 24.4675
R70 VP.n19 VP.n18 24.4675
R71 VP.n17 VP.n16 5.18913
R72 VP.n34 VP.n33 0.354971
R73 VP.n38 VP.n35 0.354971
R74 VP.n63 VP.n62 0.354971
R75 VP VP.n63 0.26696
R76 VP.n17 VP.n14 0.189894
R77 VP.n21 VP.n14 0.189894
R78 VP.n22 VP.n21 0.189894
R79 VP.n23 VP.n22 0.189894
R80 VP.n23 VP.n12 0.189894
R81 VP.n27 VP.n12 0.189894
R82 VP.n28 VP.n27 0.189894
R83 VP.n29 VP.n28 0.189894
R84 VP.n29 VP.n10 0.189894
R85 VP.n33 VP.n10 0.189894
R86 VP.n39 VP.n38 0.189894
R87 VP.n40 VP.n39 0.189894
R88 VP.n40 VP.n7 0.189894
R89 VP.n44 VP.n7 0.189894
R90 VP.n45 VP.n44 0.189894
R91 VP.n46 VP.n45 0.189894
R92 VP.n46 VP.n5 0.189894
R93 VP.n50 VP.n5 0.189894
R94 VP.n51 VP.n50 0.189894
R95 VP.n52 VP.n51 0.189894
R96 VP.n52 VP.n3 0.189894
R97 VP.n56 VP.n3 0.189894
R98 VP.n57 VP.n56 0.189894
R99 VP.n58 VP.n57 0.189894
R100 VP.n58 VP.n1 0.189894
R101 VP.n62 VP.n1 0.189894
R102 VTAIL.n530 VTAIL.n470 756.745
R103 VTAIL.n62 VTAIL.n2 756.745
R104 VTAIL.n128 VTAIL.n68 756.745
R105 VTAIL.n196 VTAIL.n136 756.745
R106 VTAIL.n464 VTAIL.n404 756.745
R107 VTAIL.n396 VTAIL.n336 756.745
R108 VTAIL.n330 VTAIL.n270 756.745
R109 VTAIL.n262 VTAIL.n202 756.745
R110 VTAIL.n490 VTAIL.n489 585
R111 VTAIL.n495 VTAIL.n494 585
R112 VTAIL.n497 VTAIL.n496 585
R113 VTAIL.n486 VTAIL.n485 585
R114 VTAIL.n503 VTAIL.n502 585
R115 VTAIL.n505 VTAIL.n504 585
R116 VTAIL.n482 VTAIL.n481 585
R117 VTAIL.n512 VTAIL.n511 585
R118 VTAIL.n513 VTAIL.n480 585
R119 VTAIL.n515 VTAIL.n514 585
R120 VTAIL.n478 VTAIL.n477 585
R121 VTAIL.n521 VTAIL.n520 585
R122 VTAIL.n523 VTAIL.n522 585
R123 VTAIL.n474 VTAIL.n473 585
R124 VTAIL.n529 VTAIL.n528 585
R125 VTAIL.n531 VTAIL.n530 585
R126 VTAIL.n22 VTAIL.n21 585
R127 VTAIL.n27 VTAIL.n26 585
R128 VTAIL.n29 VTAIL.n28 585
R129 VTAIL.n18 VTAIL.n17 585
R130 VTAIL.n35 VTAIL.n34 585
R131 VTAIL.n37 VTAIL.n36 585
R132 VTAIL.n14 VTAIL.n13 585
R133 VTAIL.n44 VTAIL.n43 585
R134 VTAIL.n45 VTAIL.n12 585
R135 VTAIL.n47 VTAIL.n46 585
R136 VTAIL.n10 VTAIL.n9 585
R137 VTAIL.n53 VTAIL.n52 585
R138 VTAIL.n55 VTAIL.n54 585
R139 VTAIL.n6 VTAIL.n5 585
R140 VTAIL.n61 VTAIL.n60 585
R141 VTAIL.n63 VTAIL.n62 585
R142 VTAIL.n88 VTAIL.n87 585
R143 VTAIL.n93 VTAIL.n92 585
R144 VTAIL.n95 VTAIL.n94 585
R145 VTAIL.n84 VTAIL.n83 585
R146 VTAIL.n101 VTAIL.n100 585
R147 VTAIL.n103 VTAIL.n102 585
R148 VTAIL.n80 VTAIL.n79 585
R149 VTAIL.n110 VTAIL.n109 585
R150 VTAIL.n111 VTAIL.n78 585
R151 VTAIL.n113 VTAIL.n112 585
R152 VTAIL.n76 VTAIL.n75 585
R153 VTAIL.n119 VTAIL.n118 585
R154 VTAIL.n121 VTAIL.n120 585
R155 VTAIL.n72 VTAIL.n71 585
R156 VTAIL.n127 VTAIL.n126 585
R157 VTAIL.n129 VTAIL.n128 585
R158 VTAIL.n156 VTAIL.n155 585
R159 VTAIL.n161 VTAIL.n160 585
R160 VTAIL.n163 VTAIL.n162 585
R161 VTAIL.n152 VTAIL.n151 585
R162 VTAIL.n169 VTAIL.n168 585
R163 VTAIL.n171 VTAIL.n170 585
R164 VTAIL.n148 VTAIL.n147 585
R165 VTAIL.n178 VTAIL.n177 585
R166 VTAIL.n179 VTAIL.n146 585
R167 VTAIL.n181 VTAIL.n180 585
R168 VTAIL.n144 VTAIL.n143 585
R169 VTAIL.n187 VTAIL.n186 585
R170 VTAIL.n189 VTAIL.n188 585
R171 VTAIL.n140 VTAIL.n139 585
R172 VTAIL.n195 VTAIL.n194 585
R173 VTAIL.n197 VTAIL.n196 585
R174 VTAIL.n465 VTAIL.n464 585
R175 VTAIL.n463 VTAIL.n462 585
R176 VTAIL.n408 VTAIL.n407 585
R177 VTAIL.n457 VTAIL.n456 585
R178 VTAIL.n455 VTAIL.n454 585
R179 VTAIL.n412 VTAIL.n411 585
R180 VTAIL.n449 VTAIL.n448 585
R181 VTAIL.n447 VTAIL.n414 585
R182 VTAIL.n446 VTAIL.n445 585
R183 VTAIL.n417 VTAIL.n415 585
R184 VTAIL.n440 VTAIL.n439 585
R185 VTAIL.n438 VTAIL.n437 585
R186 VTAIL.n421 VTAIL.n420 585
R187 VTAIL.n432 VTAIL.n431 585
R188 VTAIL.n430 VTAIL.n429 585
R189 VTAIL.n425 VTAIL.n424 585
R190 VTAIL.n397 VTAIL.n396 585
R191 VTAIL.n395 VTAIL.n394 585
R192 VTAIL.n340 VTAIL.n339 585
R193 VTAIL.n389 VTAIL.n388 585
R194 VTAIL.n387 VTAIL.n386 585
R195 VTAIL.n344 VTAIL.n343 585
R196 VTAIL.n381 VTAIL.n380 585
R197 VTAIL.n379 VTAIL.n346 585
R198 VTAIL.n378 VTAIL.n377 585
R199 VTAIL.n349 VTAIL.n347 585
R200 VTAIL.n372 VTAIL.n371 585
R201 VTAIL.n370 VTAIL.n369 585
R202 VTAIL.n353 VTAIL.n352 585
R203 VTAIL.n364 VTAIL.n363 585
R204 VTAIL.n362 VTAIL.n361 585
R205 VTAIL.n357 VTAIL.n356 585
R206 VTAIL.n331 VTAIL.n330 585
R207 VTAIL.n329 VTAIL.n328 585
R208 VTAIL.n274 VTAIL.n273 585
R209 VTAIL.n323 VTAIL.n322 585
R210 VTAIL.n321 VTAIL.n320 585
R211 VTAIL.n278 VTAIL.n277 585
R212 VTAIL.n315 VTAIL.n314 585
R213 VTAIL.n313 VTAIL.n280 585
R214 VTAIL.n312 VTAIL.n311 585
R215 VTAIL.n283 VTAIL.n281 585
R216 VTAIL.n306 VTAIL.n305 585
R217 VTAIL.n304 VTAIL.n303 585
R218 VTAIL.n287 VTAIL.n286 585
R219 VTAIL.n298 VTAIL.n297 585
R220 VTAIL.n296 VTAIL.n295 585
R221 VTAIL.n291 VTAIL.n290 585
R222 VTAIL.n263 VTAIL.n262 585
R223 VTAIL.n261 VTAIL.n260 585
R224 VTAIL.n206 VTAIL.n205 585
R225 VTAIL.n255 VTAIL.n254 585
R226 VTAIL.n253 VTAIL.n252 585
R227 VTAIL.n210 VTAIL.n209 585
R228 VTAIL.n247 VTAIL.n246 585
R229 VTAIL.n245 VTAIL.n212 585
R230 VTAIL.n244 VTAIL.n243 585
R231 VTAIL.n215 VTAIL.n213 585
R232 VTAIL.n238 VTAIL.n237 585
R233 VTAIL.n236 VTAIL.n235 585
R234 VTAIL.n219 VTAIL.n218 585
R235 VTAIL.n230 VTAIL.n229 585
R236 VTAIL.n228 VTAIL.n227 585
R237 VTAIL.n223 VTAIL.n222 585
R238 VTAIL.n491 VTAIL.t6 329.036
R239 VTAIL.n23 VTAIL.t0 329.036
R240 VTAIL.n89 VTAIL.t10 329.036
R241 VTAIL.n157 VTAIL.t12 329.036
R242 VTAIL.n426 VTAIL.t13 329.036
R243 VTAIL.n358 VTAIL.t11 329.036
R244 VTAIL.n292 VTAIL.t3 329.036
R245 VTAIL.n224 VTAIL.t2 329.036
R246 VTAIL.n495 VTAIL.n489 171.744
R247 VTAIL.n496 VTAIL.n495 171.744
R248 VTAIL.n496 VTAIL.n485 171.744
R249 VTAIL.n503 VTAIL.n485 171.744
R250 VTAIL.n504 VTAIL.n503 171.744
R251 VTAIL.n504 VTAIL.n481 171.744
R252 VTAIL.n512 VTAIL.n481 171.744
R253 VTAIL.n513 VTAIL.n512 171.744
R254 VTAIL.n514 VTAIL.n513 171.744
R255 VTAIL.n514 VTAIL.n477 171.744
R256 VTAIL.n521 VTAIL.n477 171.744
R257 VTAIL.n522 VTAIL.n521 171.744
R258 VTAIL.n522 VTAIL.n473 171.744
R259 VTAIL.n529 VTAIL.n473 171.744
R260 VTAIL.n530 VTAIL.n529 171.744
R261 VTAIL.n27 VTAIL.n21 171.744
R262 VTAIL.n28 VTAIL.n27 171.744
R263 VTAIL.n28 VTAIL.n17 171.744
R264 VTAIL.n35 VTAIL.n17 171.744
R265 VTAIL.n36 VTAIL.n35 171.744
R266 VTAIL.n36 VTAIL.n13 171.744
R267 VTAIL.n44 VTAIL.n13 171.744
R268 VTAIL.n45 VTAIL.n44 171.744
R269 VTAIL.n46 VTAIL.n45 171.744
R270 VTAIL.n46 VTAIL.n9 171.744
R271 VTAIL.n53 VTAIL.n9 171.744
R272 VTAIL.n54 VTAIL.n53 171.744
R273 VTAIL.n54 VTAIL.n5 171.744
R274 VTAIL.n61 VTAIL.n5 171.744
R275 VTAIL.n62 VTAIL.n61 171.744
R276 VTAIL.n93 VTAIL.n87 171.744
R277 VTAIL.n94 VTAIL.n93 171.744
R278 VTAIL.n94 VTAIL.n83 171.744
R279 VTAIL.n101 VTAIL.n83 171.744
R280 VTAIL.n102 VTAIL.n101 171.744
R281 VTAIL.n102 VTAIL.n79 171.744
R282 VTAIL.n110 VTAIL.n79 171.744
R283 VTAIL.n111 VTAIL.n110 171.744
R284 VTAIL.n112 VTAIL.n111 171.744
R285 VTAIL.n112 VTAIL.n75 171.744
R286 VTAIL.n119 VTAIL.n75 171.744
R287 VTAIL.n120 VTAIL.n119 171.744
R288 VTAIL.n120 VTAIL.n71 171.744
R289 VTAIL.n127 VTAIL.n71 171.744
R290 VTAIL.n128 VTAIL.n127 171.744
R291 VTAIL.n161 VTAIL.n155 171.744
R292 VTAIL.n162 VTAIL.n161 171.744
R293 VTAIL.n162 VTAIL.n151 171.744
R294 VTAIL.n169 VTAIL.n151 171.744
R295 VTAIL.n170 VTAIL.n169 171.744
R296 VTAIL.n170 VTAIL.n147 171.744
R297 VTAIL.n178 VTAIL.n147 171.744
R298 VTAIL.n179 VTAIL.n178 171.744
R299 VTAIL.n180 VTAIL.n179 171.744
R300 VTAIL.n180 VTAIL.n143 171.744
R301 VTAIL.n187 VTAIL.n143 171.744
R302 VTAIL.n188 VTAIL.n187 171.744
R303 VTAIL.n188 VTAIL.n139 171.744
R304 VTAIL.n195 VTAIL.n139 171.744
R305 VTAIL.n196 VTAIL.n195 171.744
R306 VTAIL.n464 VTAIL.n463 171.744
R307 VTAIL.n463 VTAIL.n407 171.744
R308 VTAIL.n456 VTAIL.n407 171.744
R309 VTAIL.n456 VTAIL.n455 171.744
R310 VTAIL.n455 VTAIL.n411 171.744
R311 VTAIL.n448 VTAIL.n411 171.744
R312 VTAIL.n448 VTAIL.n447 171.744
R313 VTAIL.n447 VTAIL.n446 171.744
R314 VTAIL.n446 VTAIL.n415 171.744
R315 VTAIL.n439 VTAIL.n415 171.744
R316 VTAIL.n439 VTAIL.n438 171.744
R317 VTAIL.n438 VTAIL.n420 171.744
R318 VTAIL.n431 VTAIL.n420 171.744
R319 VTAIL.n431 VTAIL.n430 171.744
R320 VTAIL.n430 VTAIL.n424 171.744
R321 VTAIL.n396 VTAIL.n395 171.744
R322 VTAIL.n395 VTAIL.n339 171.744
R323 VTAIL.n388 VTAIL.n339 171.744
R324 VTAIL.n388 VTAIL.n387 171.744
R325 VTAIL.n387 VTAIL.n343 171.744
R326 VTAIL.n380 VTAIL.n343 171.744
R327 VTAIL.n380 VTAIL.n379 171.744
R328 VTAIL.n379 VTAIL.n378 171.744
R329 VTAIL.n378 VTAIL.n347 171.744
R330 VTAIL.n371 VTAIL.n347 171.744
R331 VTAIL.n371 VTAIL.n370 171.744
R332 VTAIL.n370 VTAIL.n352 171.744
R333 VTAIL.n363 VTAIL.n352 171.744
R334 VTAIL.n363 VTAIL.n362 171.744
R335 VTAIL.n362 VTAIL.n356 171.744
R336 VTAIL.n330 VTAIL.n329 171.744
R337 VTAIL.n329 VTAIL.n273 171.744
R338 VTAIL.n322 VTAIL.n273 171.744
R339 VTAIL.n322 VTAIL.n321 171.744
R340 VTAIL.n321 VTAIL.n277 171.744
R341 VTAIL.n314 VTAIL.n277 171.744
R342 VTAIL.n314 VTAIL.n313 171.744
R343 VTAIL.n313 VTAIL.n312 171.744
R344 VTAIL.n312 VTAIL.n281 171.744
R345 VTAIL.n305 VTAIL.n281 171.744
R346 VTAIL.n305 VTAIL.n304 171.744
R347 VTAIL.n304 VTAIL.n286 171.744
R348 VTAIL.n297 VTAIL.n286 171.744
R349 VTAIL.n297 VTAIL.n296 171.744
R350 VTAIL.n296 VTAIL.n290 171.744
R351 VTAIL.n262 VTAIL.n261 171.744
R352 VTAIL.n261 VTAIL.n205 171.744
R353 VTAIL.n254 VTAIL.n205 171.744
R354 VTAIL.n254 VTAIL.n253 171.744
R355 VTAIL.n253 VTAIL.n209 171.744
R356 VTAIL.n246 VTAIL.n209 171.744
R357 VTAIL.n246 VTAIL.n245 171.744
R358 VTAIL.n245 VTAIL.n244 171.744
R359 VTAIL.n244 VTAIL.n213 171.744
R360 VTAIL.n237 VTAIL.n213 171.744
R361 VTAIL.n237 VTAIL.n236 171.744
R362 VTAIL.n236 VTAIL.n218 171.744
R363 VTAIL.n229 VTAIL.n218 171.744
R364 VTAIL.n229 VTAIL.n228 171.744
R365 VTAIL.n228 VTAIL.n222 171.744
R366 VTAIL.t6 VTAIL.n489 85.8723
R367 VTAIL.t0 VTAIL.n21 85.8723
R368 VTAIL.t10 VTAIL.n87 85.8723
R369 VTAIL.t12 VTAIL.n155 85.8723
R370 VTAIL.t13 VTAIL.n424 85.8723
R371 VTAIL.t11 VTAIL.n356 85.8723
R372 VTAIL.t3 VTAIL.n290 85.8723
R373 VTAIL.t2 VTAIL.n222 85.8723
R374 VTAIL.n403 VTAIL.n402 55.415
R375 VTAIL.n269 VTAIL.n268 55.415
R376 VTAIL.n1 VTAIL.n0 55.4148
R377 VTAIL.n135 VTAIL.n134 55.4148
R378 VTAIL.n535 VTAIL.n534 30.4399
R379 VTAIL.n67 VTAIL.n66 30.4399
R380 VTAIL.n133 VTAIL.n132 30.4399
R381 VTAIL.n201 VTAIL.n200 30.4399
R382 VTAIL.n469 VTAIL.n468 30.4399
R383 VTAIL.n401 VTAIL.n400 30.4399
R384 VTAIL.n335 VTAIL.n334 30.4399
R385 VTAIL.n267 VTAIL.n266 30.4399
R386 VTAIL.n535 VTAIL.n469 25.3238
R387 VTAIL.n267 VTAIL.n201 25.3238
R388 VTAIL.n515 VTAIL.n480 13.1884
R389 VTAIL.n47 VTAIL.n12 13.1884
R390 VTAIL.n113 VTAIL.n78 13.1884
R391 VTAIL.n181 VTAIL.n146 13.1884
R392 VTAIL.n449 VTAIL.n414 13.1884
R393 VTAIL.n381 VTAIL.n346 13.1884
R394 VTAIL.n315 VTAIL.n280 13.1884
R395 VTAIL.n247 VTAIL.n212 13.1884
R396 VTAIL.n511 VTAIL.n510 12.8005
R397 VTAIL.n516 VTAIL.n478 12.8005
R398 VTAIL.n43 VTAIL.n42 12.8005
R399 VTAIL.n48 VTAIL.n10 12.8005
R400 VTAIL.n109 VTAIL.n108 12.8005
R401 VTAIL.n114 VTAIL.n76 12.8005
R402 VTAIL.n177 VTAIL.n176 12.8005
R403 VTAIL.n182 VTAIL.n144 12.8005
R404 VTAIL.n450 VTAIL.n412 12.8005
R405 VTAIL.n445 VTAIL.n416 12.8005
R406 VTAIL.n382 VTAIL.n344 12.8005
R407 VTAIL.n377 VTAIL.n348 12.8005
R408 VTAIL.n316 VTAIL.n278 12.8005
R409 VTAIL.n311 VTAIL.n282 12.8005
R410 VTAIL.n248 VTAIL.n210 12.8005
R411 VTAIL.n243 VTAIL.n214 12.8005
R412 VTAIL.n509 VTAIL.n482 12.0247
R413 VTAIL.n520 VTAIL.n519 12.0247
R414 VTAIL.n41 VTAIL.n14 12.0247
R415 VTAIL.n52 VTAIL.n51 12.0247
R416 VTAIL.n107 VTAIL.n80 12.0247
R417 VTAIL.n118 VTAIL.n117 12.0247
R418 VTAIL.n175 VTAIL.n148 12.0247
R419 VTAIL.n186 VTAIL.n185 12.0247
R420 VTAIL.n454 VTAIL.n453 12.0247
R421 VTAIL.n444 VTAIL.n417 12.0247
R422 VTAIL.n386 VTAIL.n385 12.0247
R423 VTAIL.n376 VTAIL.n349 12.0247
R424 VTAIL.n320 VTAIL.n319 12.0247
R425 VTAIL.n310 VTAIL.n283 12.0247
R426 VTAIL.n252 VTAIL.n251 12.0247
R427 VTAIL.n242 VTAIL.n215 12.0247
R428 VTAIL.n506 VTAIL.n505 11.249
R429 VTAIL.n523 VTAIL.n476 11.249
R430 VTAIL.n38 VTAIL.n37 11.249
R431 VTAIL.n55 VTAIL.n8 11.249
R432 VTAIL.n104 VTAIL.n103 11.249
R433 VTAIL.n121 VTAIL.n74 11.249
R434 VTAIL.n172 VTAIL.n171 11.249
R435 VTAIL.n189 VTAIL.n142 11.249
R436 VTAIL.n457 VTAIL.n410 11.249
R437 VTAIL.n441 VTAIL.n440 11.249
R438 VTAIL.n389 VTAIL.n342 11.249
R439 VTAIL.n373 VTAIL.n372 11.249
R440 VTAIL.n323 VTAIL.n276 11.249
R441 VTAIL.n307 VTAIL.n306 11.249
R442 VTAIL.n255 VTAIL.n208 11.249
R443 VTAIL.n239 VTAIL.n238 11.249
R444 VTAIL.n491 VTAIL.n490 10.7239
R445 VTAIL.n23 VTAIL.n22 10.7239
R446 VTAIL.n89 VTAIL.n88 10.7239
R447 VTAIL.n157 VTAIL.n156 10.7239
R448 VTAIL.n426 VTAIL.n425 10.7239
R449 VTAIL.n358 VTAIL.n357 10.7239
R450 VTAIL.n292 VTAIL.n291 10.7239
R451 VTAIL.n224 VTAIL.n223 10.7239
R452 VTAIL.n502 VTAIL.n484 10.4732
R453 VTAIL.n524 VTAIL.n474 10.4732
R454 VTAIL.n34 VTAIL.n16 10.4732
R455 VTAIL.n56 VTAIL.n6 10.4732
R456 VTAIL.n100 VTAIL.n82 10.4732
R457 VTAIL.n122 VTAIL.n72 10.4732
R458 VTAIL.n168 VTAIL.n150 10.4732
R459 VTAIL.n190 VTAIL.n140 10.4732
R460 VTAIL.n458 VTAIL.n408 10.4732
R461 VTAIL.n437 VTAIL.n419 10.4732
R462 VTAIL.n390 VTAIL.n340 10.4732
R463 VTAIL.n369 VTAIL.n351 10.4732
R464 VTAIL.n324 VTAIL.n274 10.4732
R465 VTAIL.n303 VTAIL.n285 10.4732
R466 VTAIL.n256 VTAIL.n206 10.4732
R467 VTAIL.n235 VTAIL.n217 10.4732
R468 VTAIL.n501 VTAIL.n486 9.69747
R469 VTAIL.n528 VTAIL.n527 9.69747
R470 VTAIL.n33 VTAIL.n18 9.69747
R471 VTAIL.n60 VTAIL.n59 9.69747
R472 VTAIL.n99 VTAIL.n84 9.69747
R473 VTAIL.n126 VTAIL.n125 9.69747
R474 VTAIL.n167 VTAIL.n152 9.69747
R475 VTAIL.n194 VTAIL.n193 9.69747
R476 VTAIL.n462 VTAIL.n461 9.69747
R477 VTAIL.n436 VTAIL.n421 9.69747
R478 VTAIL.n394 VTAIL.n393 9.69747
R479 VTAIL.n368 VTAIL.n353 9.69747
R480 VTAIL.n328 VTAIL.n327 9.69747
R481 VTAIL.n302 VTAIL.n287 9.69747
R482 VTAIL.n260 VTAIL.n259 9.69747
R483 VTAIL.n234 VTAIL.n219 9.69747
R484 VTAIL.n534 VTAIL.n533 9.45567
R485 VTAIL.n66 VTAIL.n65 9.45567
R486 VTAIL.n132 VTAIL.n131 9.45567
R487 VTAIL.n200 VTAIL.n199 9.45567
R488 VTAIL.n468 VTAIL.n467 9.45567
R489 VTAIL.n400 VTAIL.n399 9.45567
R490 VTAIL.n334 VTAIL.n333 9.45567
R491 VTAIL.n266 VTAIL.n265 9.45567
R492 VTAIL.n533 VTAIL.n532 9.3005
R493 VTAIL.n472 VTAIL.n471 9.3005
R494 VTAIL.n527 VTAIL.n526 9.3005
R495 VTAIL.n525 VTAIL.n524 9.3005
R496 VTAIL.n476 VTAIL.n475 9.3005
R497 VTAIL.n519 VTAIL.n518 9.3005
R498 VTAIL.n517 VTAIL.n516 9.3005
R499 VTAIL.n493 VTAIL.n492 9.3005
R500 VTAIL.n488 VTAIL.n487 9.3005
R501 VTAIL.n499 VTAIL.n498 9.3005
R502 VTAIL.n501 VTAIL.n500 9.3005
R503 VTAIL.n484 VTAIL.n483 9.3005
R504 VTAIL.n507 VTAIL.n506 9.3005
R505 VTAIL.n509 VTAIL.n508 9.3005
R506 VTAIL.n510 VTAIL.n479 9.3005
R507 VTAIL.n65 VTAIL.n64 9.3005
R508 VTAIL.n4 VTAIL.n3 9.3005
R509 VTAIL.n59 VTAIL.n58 9.3005
R510 VTAIL.n57 VTAIL.n56 9.3005
R511 VTAIL.n8 VTAIL.n7 9.3005
R512 VTAIL.n51 VTAIL.n50 9.3005
R513 VTAIL.n49 VTAIL.n48 9.3005
R514 VTAIL.n25 VTAIL.n24 9.3005
R515 VTAIL.n20 VTAIL.n19 9.3005
R516 VTAIL.n31 VTAIL.n30 9.3005
R517 VTAIL.n33 VTAIL.n32 9.3005
R518 VTAIL.n16 VTAIL.n15 9.3005
R519 VTAIL.n39 VTAIL.n38 9.3005
R520 VTAIL.n41 VTAIL.n40 9.3005
R521 VTAIL.n42 VTAIL.n11 9.3005
R522 VTAIL.n131 VTAIL.n130 9.3005
R523 VTAIL.n70 VTAIL.n69 9.3005
R524 VTAIL.n125 VTAIL.n124 9.3005
R525 VTAIL.n123 VTAIL.n122 9.3005
R526 VTAIL.n74 VTAIL.n73 9.3005
R527 VTAIL.n117 VTAIL.n116 9.3005
R528 VTAIL.n115 VTAIL.n114 9.3005
R529 VTAIL.n91 VTAIL.n90 9.3005
R530 VTAIL.n86 VTAIL.n85 9.3005
R531 VTAIL.n97 VTAIL.n96 9.3005
R532 VTAIL.n99 VTAIL.n98 9.3005
R533 VTAIL.n82 VTAIL.n81 9.3005
R534 VTAIL.n105 VTAIL.n104 9.3005
R535 VTAIL.n107 VTAIL.n106 9.3005
R536 VTAIL.n108 VTAIL.n77 9.3005
R537 VTAIL.n199 VTAIL.n198 9.3005
R538 VTAIL.n138 VTAIL.n137 9.3005
R539 VTAIL.n193 VTAIL.n192 9.3005
R540 VTAIL.n191 VTAIL.n190 9.3005
R541 VTAIL.n142 VTAIL.n141 9.3005
R542 VTAIL.n185 VTAIL.n184 9.3005
R543 VTAIL.n183 VTAIL.n182 9.3005
R544 VTAIL.n159 VTAIL.n158 9.3005
R545 VTAIL.n154 VTAIL.n153 9.3005
R546 VTAIL.n165 VTAIL.n164 9.3005
R547 VTAIL.n167 VTAIL.n166 9.3005
R548 VTAIL.n150 VTAIL.n149 9.3005
R549 VTAIL.n173 VTAIL.n172 9.3005
R550 VTAIL.n175 VTAIL.n174 9.3005
R551 VTAIL.n176 VTAIL.n145 9.3005
R552 VTAIL.n428 VTAIL.n427 9.3005
R553 VTAIL.n423 VTAIL.n422 9.3005
R554 VTAIL.n434 VTAIL.n433 9.3005
R555 VTAIL.n436 VTAIL.n435 9.3005
R556 VTAIL.n419 VTAIL.n418 9.3005
R557 VTAIL.n442 VTAIL.n441 9.3005
R558 VTAIL.n444 VTAIL.n443 9.3005
R559 VTAIL.n416 VTAIL.n413 9.3005
R560 VTAIL.n467 VTAIL.n466 9.3005
R561 VTAIL.n406 VTAIL.n405 9.3005
R562 VTAIL.n461 VTAIL.n460 9.3005
R563 VTAIL.n459 VTAIL.n458 9.3005
R564 VTAIL.n410 VTAIL.n409 9.3005
R565 VTAIL.n453 VTAIL.n452 9.3005
R566 VTAIL.n451 VTAIL.n450 9.3005
R567 VTAIL.n360 VTAIL.n359 9.3005
R568 VTAIL.n355 VTAIL.n354 9.3005
R569 VTAIL.n366 VTAIL.n365 9.3005
R570 VTAIL.n368 VTAIL.n367 9.3005
R571 VTAIL.n351 VTAIL.n350 9.3005
R572 VTAIL.n374 VTAIL.n373 9.3005
R573 VTAIL.n376 VTAIL.n375 9.3005
R574 VTAIL.n348 VTAIL.n345 9.3005
R575 VTAIL.n399 VTAIL.n398 9.3005
R576 VTAIL.n338 VTAIL.n337 9.3005
R577 VTAIL.n393 VTAIL.n392 9.3005
R578 VTAIL.n391 VTAIL.n390 9.3005
R579 VTAIL.n342 VTAIL.n341 9.3005
R580 VTAIL.n385 VTAIL.n384 9.3005
R581 VTAIL.n383 VTAIL.n382 9.3005
R582 VTAIL.n294 VTAIL.n293 9.3005
R583 VTAIL.n289 VTAIL.n288 9.3005
R584 VTAIL.n300 VTAIL.n299 9.3005
R585 VTAIL.n302 VTAIL.n301 9.3005
R586 VTAIL.n285 VTAIL.n284 9.3005
R587 VTAIL.n308 VTAIL.n307 9.3005
R588 VTAIL.n310 VTAIL.n309 9.3005
R589 VTAIL.n282 VTAIL.n279 9.3005
R590 VTAIL.n333 VTAIL.n332 9.3005
R591 VTAIL.n272 VTAIL.n271 9.3005
R592 VTAIL.n327 VTAIL.n326 9.3005
R593 VTAIL.n325 VTAIL.n324 9.3005
R594 VTAIL.n276 VTAIL.n275 9.3005
R595 VTAIL.n319 VTAIL.n318 9.3005
R596 VTAIL.n317 VTAIL.n316 9.3005
R597 VTAIL.n226 VTAIL.n225 9.3005
R598 VTAIL.n221 VTAIL.n220 9.3005
R599 VTAIL.n232 VTAIL.n231 9.3005
R600 VTAIL.n234 VTAIL.n233 9.3005
R601 VTAIL.n217 VTAIL.n216 9.3005
R602 VTAIL.n240 VTAIL.n239 9.3005
R603 VTAIL.n242 VTAIL.n241 9.3005
R604 VTAIL.n214 VTAIL.n211 9.3005
R605 VTAIL.n265 VTAIL.n264 9.3005
R606 VTAIL.n204 VTAIL.n203 9.3005
R607 VTAIL.n259 VTAIL.n258 9.3005
R608 VTAIL.n257 VTAIL.n256 9.3005
R609 VTAIL.n208 VTAIL.n207 9.3005
R610 VTAIL.n251 VTAIL.n250 9.3005
R611 VTAIL.n249 VTAIL.n248 9.3005
R612 VTAIL.n498 VTAIL.n497 8.92171
R613 VTAIL.n531 VTAIL.n472 8.92171
R614 VTAIL.n30 VTAIL.n29 8.92171
R615 VTAIL.n63 VTAIL.n4 8.92171
R616 VTAIL.n96 VTAIL.n95 8.92171
R617 VTAIL.n129 VTAIL.n70 8.92171
R618 VTAIL.n164 VTAIL.n163 8.92171
R619 VTAIL.n197 VTAIL.n138 8.92171
R620 VTAIL.n465 VTAIL.n406 8.92171
R621 VTAIL.n433 VTAIL.n432 8.92171
R622 VTAIL.n397 VTAIL.n338 8.92171
R623 VTAIL.n365 VTAIL.n364 8.92171
R624 VTAIL.n331 VTAIL.n272 8.92171
R625 VTAIL.n299 VTAIL.n298 8.92171
R626 VTAIL.n263 VTAIL.n204 8.92171
R627 VTAIL.n231 VTAIL.n230 8.92171
R628 VTAIL.n494 VTAIL.n488 8.14595
R629 VTAIL.n532 VTAIL.n470 8.14595
R630 VTAIL.n26 VTAIL.n20 8.14595
R631 VTAIL.n64 VTAIL.n2 8.14595
R632 VTAIL.n92 VTAIL.n86 8.14595
R633 VTAIL.n130 VTAIL.n68 8.14595
R634 VTAIL.n160 VTAIL.n154 8.14595
R635 VTAIL.n198 VTAIL.n136 8.14595
R636 VTAIL.n466 VTAIL.n404 8.14595
R637 VTAIL.n429 VTAIL.n423 8.14595
R638 VTAIL.n398 VTAIL.n336 8.14595
R639 VTAIL.n361 VTAIL.n355 8.14595
R640 VTAIL.n332 VTAIL.n270 8.14595
R641 VTAIL.n295 VTAIL.n289 8.14595
R642 VTAIL.n264 VTAIL.n202 8.14595
R643 VTAIL.n227 VTAIL.n221 8.14595
R644 VTAIL.n493 VTAIL.n490 7.3702
R645 VTAIL.n25 VTAIL.n22 7.3702
R646 VTAIL.n91 VTAIL.n88 7.3702
R647 VTAIL.n159 VTAIL.n156 7.3702
R648 VTAIL.n428 VTAIL.n425 7.3702
R649 VTAIL.n360 VTAIL.n357 7.3702
R650 VTAIL.n294 VTAIL.n291 7.3702
R651 VTAIL.n226 VTAIL.n223 7.3702
R652 VTAIL.n494 VTAIL.n493 5.81868
R653 VTAIL.n534 VTAIL.n470 5.81868
R654 VTAIL.n26 VTAIL.n25 5.81868
R655 VTAIL.n66 VTAIL.n2 5.81868
R656 VTAIL.n92 VTAIL.n91 5.81868
R657 VTAIL.n132 VTAIL.n68 5.81868
R658 VTAIL.n160 VTAIL.n159 5.81868
R659 VTAIL.n200 VTAIL.n136 5.81868
R660 VTAIL.n468 VTAIL.n404 5.81868
R661 VTAIL.n429 VTAIL.n428 5.81868
R662 VTAIL.n400 VTAIL.n336 5.81868
R663 VTAIL.n361 VTAIL.n360 5.81868
R664 VTAIL.n334 VTAIL.n270 5.81868
R665 VTAIL.n295 VTAIL.n294 5.81868
R666 VTAIL.n266 VTAIL.n202 5.81868
R667 VTAIL.n227 VTAIL.n226 5.81868
R668 VTAIL.n497 VTAIL.n488 5.04292
R669 VTAIL.n532 VTAIL.n531 5.04292
R670 VTAIL.n29 VTAIL.n20 5.04292
R671 VTAIL.n64 VTAIL.n63 5.04292
R672 VTAIL.n95 VTAIL.n86 5.04292
R673 VTAIL.n130 VTAIL.n129 5.04292
R674 VTAIL.n163 VTAIL.n154 5.04292
R675 VTAIL.n198 VTAIL.n197 5.04292
R676 VTAIL.n466 VTAIL.n465 5.04292
R677 VTAIL.n432 VTAIL.n423 5.04292
R678 VTAIL.n398 VTAIL.n397 5.04292
R679 VTAIL.n364 VTAIL.n355 5.04292
R680 VTAIL.n332 VTAIL.n331 5.04292
R681 VTAIL.n298 VTAIL.n289 5.04292
R682 VTAIL.n264 VTAIL.n263 5.04292
R683 VTAIL.n230 VTAIL.n221 5.04292
R684 VTAIL.n498 VTAIL.n486 4.26717
R685 VTAIL.n528 VTAIL.n472 4.26717
R686 VTAIL.n30 VTAIL.n18 4.26717
R687 VTAIL.n60 VTAIL.n4 4.26717
R688 VTAIL.n96 VTAIL.n84 4.26717
R689 VTAIL.n126 VTAIL.n70 4.26717
R690 VTAIL.n164 VTAIL.n152 4.26717
R691 VTAIL.n194 VTAIL.n138 4.26717
R692 VTAIL.n462 VTAIL.n406 4.26717
R693 VTAIL.n433 VTAIL.n421 4.26717
R694 VTAIL.n394 VTAIL.n338 4.26717
R695 VTAIL.n365 VTAIL.n353 4.26717
R696 VTAIL.n328 VTAIL.n272 4.26717
R697 VTAIL.n299 VTAIL.n287 4.26717
R698 VTAIL.n260 VTAIL.n204 4.26717
R699 VTAIL.n231 VTAIL.n219 4.26717
R700 VTAIL.n502 VTAIL.n501 3.49141
R701 VTAIL.n527 VTAIL.n474 3.49141
R702 VTAIL.n34 VTAIL.n33 3.49141
R703 VTAIL.n59 VTAIL.n6 3.49141
R704 VTAIL.n100 VTAIL.n99 3.49141
R705 VTAIL.n125 VTAIL.n72 3.49141
R706 VTAIL.n168 VTAIL.n167 3.49141
R707 VTAIL.n193 VTAIL.n140 3.49141
R708 VTAIL.n461 VTAIL.n408 3.49141
R709 VTAIL.n437 VTAIL.n436 3.49141
R710 VTAIL.n393 VTAIL.n340 3.49141
R711 VTAIL.n369 VTAIL.n368 3.49141
R712 VTAIL.n327 VTAIL.n274 3.49141
R713 VTAIL.n303 VTAIL.n302 3.49141
R714 VTAIL.n259 VTAIL.n206 3.49141
R715 VTAIL.n235 VTAIL.n234 3.49141
R716 VTAIL.n505 VTAIL.n484 2.71565
R717 VTAIL.n524 VTAIL.n523 2.71565
R718 VTAIL.n37 VTAIL.n16 2.71565
R719 VTAIL.n56 VTAIL.n55 2.71565
R720 VTAIL.n103 VTAIL.n82 2.71565
R721 VTAIL.n122 VTAIL.n121 2.71565
R722 VTAIL.n171 VTAIL.n150 2.71565
R723 VTAIL.n190 VTAIL.n189 2.71565
R724 VTAIL.n458 VTAIL.n457 2.71565
R725 VTAIL.n440 VTAIL.n419 2.71565
R726 VTAIL.n390 VTAIL.n389 2.71565
R727 VTAIL.n372 VTAIL.n351 2.71565
R728 VTAIL.n324 VTAIL.n323 2.71565
R729 VTAIL.n306 VTAIL.n285 2.71565
R730 VTAIL.n256 VTAIL.n255 2.71565
R731 VTAIL.n238 VTAIL.n217 2.71565
R732 VTAIL.n0 VTAIL.t1 2.7025
R733 VTAIL.n0 VTAIL.t5 2.7025
R734 VTAIL.n134 VTAIL.t15 2.7025
R735 VTAIL.n134 VTAIL.t9 2.7025
R736 VTAIL.n402 VTAIL.t8 2.7025
R737 VTAIL.n402 VTAIL.t14 2.7025
R738 VTAIL.n268 VTAIL.t4 2.7025
R739 VTAIL.n268 VTAIL.t7 2.7025
R740 VTAIL.n269 VTAIL.n267 2.58671
R741 VTAIL.n335 VTAIL.n269 2.58671
R742 VTAIL.n403 VTAIL.n401 2.58671
R743 VTAIL.n469 VTAIL.n403 2.58671
R744 VTAIL.n201 VTAIL.n135 2.58671
R745 VTAIL.n135 VTAIL.n133 2.58671
R746 VTAIL.n67 VTAIL.n1 2.58671
R747 VTAIL VTAIL.n535 2.52852
R748 VTAIL.n427 VTAIL.n426 2.41282
R749 VTAIL.n359 VTAIL.n358 2.41282
R750 VTAIL.n293 VTAIL.n292 2.41282
R751 VTAIL.n225 VTAIL.n224 2.41282
R752 VTAIL.n492 VTAIL.n491 2.41282
R753 VTAIL.n24 VTAIL.n23 2.41282
R754 VTAIL.n90 VTAIL.n89 2.41282
R755 VTAIL.n158 VTAIL.n157 2.41282
R756 VTAIL.n506 VTAIL.n482 1.93989
R757 VTAIL.n520 VTAIL.n476 1.93989
R758 VTAIL.n38 VTAIL.n14 1.93989
R759 VTAIL.n52 VTAIL.n8 1.93989
R760 VTAIL.n104 VTAIL.n80 1.93989
R761 VTAIL.n118 VTAIL.n74 1.93989
R762 VTAIL.n172 VTAIL.n148 1.93989
R763 VTAIL.n186 VTAIL.n142 1.93989
R764 VTAIL.n454 VTAIL.n410 1.93989
R765 VTAIL.n441 VTAIL.n417 1.93989
R766 VTAIL.n386 VTAIL.n342 1.93989
R767 VTAIL.n373 VTAIL.n349 1.93989
R768 VTAIL.n320 VTAIL.n276 1.93989
R769 VTAIL.n307 VTAIL.n283 1.93989
R770 VTAIL.n252 VTAIL.n208 1.93989
R771 VTAIL.n239 VTAIL.n215 1.93989
R772 VTAIL.n511 VTAIL.n509 1.16414
R773 VTAIL.n519 VTAIL.n478 1.16414
R774 VTAIL.n43 VTAIL.n41 1.16414
R775 VTAIL.n51 VTAIL.n10 1.16414
R776 VTAIL.n109 VTAIL.n107 1.16414
R777 VTAIL.n117 VTAIL.n76 1.16414
R778 VTAIL.n177 VTAIL.n175 1.16414
R779 VTAIL.n185 VTAIL.n144 1.16414
R780 VTAIL.n453 VTAIL.n412 1.16414
R781 VTAIL.n445 VTAIL.n444 1.16414
R782 VTAIL.n385 VTAIL.n344 1.16414
R783 VTAIL.n377 VTAIL.n376 1.16414
R784 VTAIL.n319 VTAIL.n278 1.16414
R785 VTAIL.n311 VTAIL.n310 1.16414
R786 VTAIL.n251 VTAIL.n210 1.16414
R787 VTAIL.n243 VTAIL.n242 1.16414
R788 VTAIL.n401 VTAIL.n335 0.470328
R789 VTAIL.n133 VTAIL.n67 0.470328
R790 VTAIL.n510 VTAIL.n480 0.388379
R791 VTAIL.n516 VTAIL.n515 0.388379
R792 VTAIL.n42 VTAIL.n12 0.388379
R793 VTAIL.n48 VTAIL.n47 0.388379
R794 VTAIL.n108 VTAIL.n78 0.388379
R795 VTAIL.n114 VTAIL.n113 0.388379
R796 VTAIL.n176 VTAIL.n146 0.388379
R797 VTAIL.n182 VTAIL.n181 0.388379
R798 VTAIL.n450 VTAIL.n449 0.388379
R799 VTAIL.n416 VTAIL.n414 0.388379
R800 VTAIL.n382 VTAIL.n381 0.388379
R801 VTAIL.n348 VTAIL.n346 0.388379
R802 VTAIL.n316 VTAIL.n315 0.388379
R803 VTAIL.n282 VTAIL.n280 0.388379
R804 VTAIL.n248 VTAIL.n247 0.388379
R805 VTAIL.n214 VTAIL.n212 0.388379
R806 VTAIL.n492 VTAIL.n487 0.155672
R807 VTAIL.n499 VTAIL.n487 0.155672
R808 VTAIL.n500 VTAIL.n499 0.155672
R809 VTAIL.n500 VTAIL.n483 0.155672
R810 VTAIL.n507 VTAIL.n483 0.155672
R811 VTAIL.n508 VTAIL.n507 0.155672
R812 VTAIL.n508 VTAIL.n479 0.155672
R813 VTAIL.n517 VTAIL.n479 0.155672
R814 VTAIL.n518 VTAIL.n517 0.155672
R815 VTAIL.n518 VTAIL.n475 0.155672
R816 VTAIL.n525 VTAIL.n475 0.155672
R817 VTAIL.n526 VTAIL.n525 0.155672
R818 VTAIL.n526 VTAIL.n471 0.155672
R819 VTAIL.n533 VTAIL.n471 0.155672
R820 VTAIL.n24 VTAIL.n19 0.155672
R821 VTAIL.n31 VTAIL.n19 0.155672
R822 VTAIL.n32 VTAIL.n31 0.155672
R823 VTAIL.n32 VTAIL.n15 0.155672
R824 VTAIL.n39 VTAIL.n15 0.155672
R825 VTAIL.n40 VTAIL.n39 0.155672
R826 VTAIL.n40 VTAIL.n11 0.155672
R827 VTAIL.n49 VTAIL.n11 0.155672
R828 VTAIL.n50 VTAIL.n49 0.155672
R829 VTAIL.n50 VTAIL.n7 0.155672
R830 VTAIL.n57 VTAIL.n7 0.155672
R831 VTAIL.n58 VTAIL.n57 0.155672
R832 VTAIL.n58 VTAIL.n3 0.155672
R833 VTAIL.n65 VTAIL.n3 0.155672
R834 VTAIL.n90 VTAIL.n85 0.155672
R835 VTAIL.n97 VTAIL.n85 0.155672
R836 VTAIL.n98 VTAIL.n97 0.155672
R837 VTAIL.n98 VTAIL.n81 0.155672
R838 VTAIL.n105 VTAIL.n81 0.155672
R839 VTAIL.n106 VTAIL.n105 0.155672
R840 VTAIL.n106 VTAIL.n77 0.155672
R841 VTAIL.n115 VTAIL.n77 0.155672
R842 VTAIL.n116 VTAIL.n115 0.155672
R843 VTAIL.n116 VTAIL.n73 0.155672
R844 VTAIL.n123 VTAIL.n73 0.155672
R845 VTAIL.n124 VTAIL.n123 0.155672
R846 VTAIL.n124 VTAIL.n69 0.155672
R847 VTAIL.n131 VTAIL.n69 0.155672
R848 VTAIL.n158 VTAIL.n153 0.155672
R849 VTAIL.n165 VTAIL.n153 0.155672
R850 VTAIL.n166 VTAIL.n165 0.155672
R851 VTAIL.n166 VTAIL.n149 0.155672
R852 VTAIL.n173 VTAIL.n149 0.155672
R853 VTAIL.n174 VTAIL.n173 0.155672
R854 VTAIL.n174 VTAIL.n145 0.155672
R855 VTAIL.n183 VTAIL.n145 0.155672
R856 VTAIL.n184 VTAIL.n183 0.155672
R857 VTAIL.n184 VTAIL.n141 0.155672
R858 VTAIL.n191 VTAIL.n141 0.155672
R859 VTAIL.n192 VTAIL.n191 0.155672
R860 VTAIL.n192 VTAIL.n137 0.155672
R861 VTAIL.n199 VTAIL.n137 0.155672
R862 VTAIL.n467 VTAIL.n405 0.155672
R863 VTAIL.n460 VTAIL.n405 0.155672
R864 VTAIL.n460 VTAIL.n459 0.155672
R865 VTAIL.n459 VTAIL.n409 0.155672
R866 VTAIL.n452 VTAIL.n409 0.155672
R867 VTAIL.n452 VTAIL.n451 0.155672
R868 VTAIL.n451 VTAIL.n413 0.155672
R869 VTAIL.n443 VTAIL.n413 0.155672
R870 VTAIL.n443 VTAIL.n442 0.155672
R871 VTAIL.n442 VTAIL.n418 0.155672
R872 VTAIL.n435 VTAIL.n418 0.155672
R873 VTAIL.n435 VTAIL.n434 0.155672
R874 VTAIL.n434 VTAIL.n422 0.155672
R875 VTAIL.n427 VTAIL.n422 0.155672
R876 VTAIL.n399 VTAIL.n337 0.155672
R877 VTAIL.n392 VTAIL.n337 0.155672
R878 VTAIL.n392 VTAIL.n391 0.155672
R879 VTAIL.n391 VTAIL.n341 0.155672
R880 VTAIL.n384 VTAIL.n341 0.155672
R881 VTAIL.n384 VTAIL.n383 0.155672
R882 VTAIL.n383 VTAIL.n345 0.155672
R883 VTAIL.n375 VTAIL.n345 0.155672
R884 VTAIL.n375 VTAIL.n374 0.155672
R885 VTAIL.n374 VTAIL.n350 0.155672
R886 VTAIL.n367 VTAIL.n350 0.155672
R887 VTAIL.n367 VTAIL.n366 0.155672
R888 VTAIL.n366 VTAIL.n354 0.155672
R889 VTAIL.n359 VTAIL.n354 0.155672
R890 VTAIL.n333 VTAIL.n271 0.155672
R891 VTAIL.n326 VTAIL.n271 0.155672
R892 VTAIL.n326 VTAIL.n325 0.155672
R893 VTAIL.n325 VTAIL.n275 0.155672
R894 VTAIL.n318 VTAIL.n275 0.155672
R895 VTAIL.n318 VTAIL.n317 0.155672
R896 VTAIL.n317 VTAIL.n279 0.155672
R897 VTAIL.n309 VTAIL.n279 0.155672
R898 VTAIL.n309 VTAIL.n308 0.155672
R899 VTAIL.n308 VTAIL.n284 0.155672
R900 VTAIL.n301 VTAIL.n284 0.155672
R901 VTAIL.n301 VTAIL.n300 0.155672
R902 VTAIL.n300 VTAIL.n288 0.155672
R903 VTAIL.n293 VTAIL.n288 0.155672
R904 VTAIL.n265 VTAIL.n203 0.155672
R905 VTAIL.n258 VTAIL.n203 0.155672
R906 VTAIL.n258 VTAIL.n257 0.155672
R907 VTAIL.n257 VTAIL.n207 0.155672
R908 VTAIL.n250 VTAIL.n207 0.155672
R909 VTAIL.n250 VTAIL.n249 0.155672
R910 VTAIL.n249 VTAIL.n211 0.155672
R911 VTAIL.n241 VTAIL.n211 0.155672
R912 VTAIL.n241 VTAIL.n240 0.155672
R913 VTAIL.n240 VTAIL.n216 0.155672
R914 VTAIL.n233 VTAIL.n216 0.155672
R915 VTAIL.n233 VTAIL.n232 0.155672
R916 VTAIL.n232 VTAIL.n220 0.155672
R917 VTAIL.n225 VTAIL.n220 0.155672
R918 VTAIL VTAIL.n1 0.0586897
R919 VDD1 VDD1.n0 73.4451
R920 VDD1.n3 VDD1.n2 73.3313
R921 VDD1.n3 VDD1.n1 73.3313
R922 VDD1.n5 VDD1.n4 72.0936
R923 VDD1.n5 VDD1.n3 46.3069
R924 VDD1.n4 VDD1.t6 2.7025
R925 VDD1.n4 VDD1.t7 2.7025
R926 VDD1.n0 VDD1.t3 2.7025
R927 VDD1.n0 VDD1.t1 2.7025
R928 VDD1.n2 VDD1.t5 2.7025
R929 VDD1.n2 VDD1.t2 2.7025
R930 VDD1.n1 VDD1.t0 2.7025
R931 VDD1.n1 VDD1.t4 2.7025
R932 VDD1 VDD1.n5 1.23541
R933 VN.n50 VN.n49 161.3
R934 VN.n48 VN.n27 161.3
R935 VN.n47 VN.n46 161.3
R936 VN.n45 VN.n28 161.3
R937 VN.n44 VN.n43 161.3
R938 VN.n42 VN.n29 161.3
R939 VN.n41 VN.n40 161.3
R940 VN.n39 VN.n30 161.3
R941 VN.n38 VN.n37 161.3
R942 VN.n36 VN.n31 161.3
R943 VN.n35 VN.n34 161.3
R944 VN.n24 VN.n23 161.3
R945 VN.n22 VN.n1 161.3
R946 VN.n21 VN.n20 161.3
R947 VN.n19 VN.n2 161.3
R948 VN.n18 VN.n17 161.3
R949 VN.n16 VN.n3 161.3
R950 VN.n15 VN.n14 161.3
R951 VN.n13 VN.n4 161.3
R952 VN.n12 VN.n11 161.3
R953 VN.n10 VN.n5 161.3
R954 VN.n9 VN.n8 161.3
R955 VN.n7 VN.t5 140.736
R956 VN.n33 VN.t2 140.736
R957 VN.n0 VN.t6 108.585
R958 VN.n16 VN.t3 108.585
R959 VN.n6 VN.t0 108.585
R960 VN.n26 VN.t1 108.585
R961 VN.n42 VN.t7 108.585
R962 VN.n32 VN.t4 108.585
R963 VN.n51 VN.n26 65.6004
R964 VN.n25 VN.n0 65.6004
R965 VN VN.n51 51.5207
R966 VN.n33 VN.n32 48.9288
R967 VN.n7 VN.n6 48.9288
R968 VN.n11 VN.n10 40.4934
R969 VN.n11 VN.n4 40.4934
R970 VN.n21 VN.n2 40.4934
R971 VN.n22 VN.n21 40.4934
R972 VN.n37 VN.n36 40.4934
R973 VN.n37 VN.n30 40.4934
R974 VN.n47 VN.n28 40.4934
R975 VN.n48 VN.n47 40.4934
R976 VN.n9 VN.n6 24.4675
R977 VN.n10 VN.n9 24.4675
R978 VN.n15 VN.n4 24.4675
R979 VN.n16 VN.n15 24.4675
R980 VN.n17 VN.n16 24.4675
R981 VN.n17 VN.n2 24.4675
R982 VN.n23 VN.n22 24.4675
R983 VN.n23 VN.n0 24.4675
R984 VN.n36 VN.n35 24.4675
R985 VN.n35 VN.n32 24.4675
R986 VN.n43 VN.n28 24.4675
R987 VN.n43 VN.n42 24.4675
R988 VN.n42 VN.n41 24.4675
R989 VN.n41 VN.n30 24.4675
R990 VN.n49 VN.n26 24.4675
R991 VN.n49 VN.n48 24.4675
R992 VN.n34 VN.n33 5.18917
R993 VN.n8 VN.n7 5.18917
R994 VN.n51 VN.n50 0.354971
R995 VN.n25 VN.n24 0.354971
R996 VN VN.n25 0.26696
R997 VN.n50 VN.n27 0.189894
R998 VN.n46 VN.n27 0.189894
R999 VN.n46 VN.n45 0.189894
R1000 VN.n45 VN.n44 0.189894
R1001 VN.n44 VN.n29 0.189894
R1002 VN.n40 VN.n29 0.189894
R1003 VN.n40 VN.n39 0.189894
R1004 VN.n39 VN.n38 0.189894
R1005 VN.n38 VN.n31 0.189894
R1006 VN.n34 VN.n31 0.189894
R1007 VN.n8 VN.n5 0.189894
R1008 VN.n12 VN.n5 0.189894
R1009 VN.n13 VN.n12 0.189894
R1010 VN.n14 VN.n13 0.189894
R1011 VN.n14 VN.n3 0.189894
R1012 VN.n18 VN.n3 0.189894
R1013 VN.n19 VN.n18 0.189894
R1014 VN.n20 VN.n19 0.189894
R1015 VN.n20 VN.n1 0.189894
R1016 VN.n24 VN.n1 0.189894
R1017 VDD2.n2 VDD2.n1 73.3313
R1018 VDD2.n2 VDD2.n0 73.3313
R1019 VDD2 VDD2.n5 73.3285
R1020 VDD2.n4 VDD2.n3 72.0938
R1021 VDD2.n4 VDD2.n2 45.7239
R1022 VDD2.n5 VDD2.t3 2.7025
R1023 VDD2.n5 VDD2.t5 2.7025
R1024 VDD2.n3 VDD2.t6 2.7025
R1025 VDD2.n3 VDD2.t0 2.7025
R1026 VDD2.n1 VDD2.t4 2.7025
R1027 VDD2.n1 VDD2.t1 2.7025
R1028 VDD2.n0 VDD2.t2 2.7025
R1029 VDD2.n0 VDD2.t7 2.7025
R1030 VDD2 VDD2.n4 1.35179
R1031 B.n583 B.n78 585
R1032 B.n585 B.n584 585
R1033 B.n586 B.n77 585
R1034 B.n588 B.n587 585
R1035 B.n589 B.n76 585
R1036 B.n591 B.n590 585
R1037 B.n592 B.n75 585
R1038 B.n594 B.n593 585
R1039 B.n595 B.n74 585
R1040 B.n597 B.n596 585
R1041 B.n598 B.n73 585
R1042 B.n600 B.n599 585
R1043 B.n601 B.n72 585
R1044 B.n603 B.n602 585
R1045 B.n604 B.n71 585
R1046 B.n606 B.n605 585
R1047 B.n607 B.n70 585
R1048 B.n609 B.n608 585
R1049 B.n610 B.n69 585
R1050 B.n612 B.n611 585
R1051 B.n613 B.n68 585
R1052 B.n615 B.n614 585
R1053 B.n616 B.n67 585
R1054 B.n618 B.n617 585
R1055 B.n619 B.n66 585
R1056 B.n621 B.n620 585
R1057 B.n622 B.n65 585
R1058 B.n624 B.n623 585
R1059 B.n625 B.n64 585
R1060 B.n627 B.n626 585
R1061 B.n628 B.n63 585
R1062 B.n630 B.n629 585
R1063 B.n631 B.n62 585
R1064 B.n633 B.n632 585
R1065 B.n634 B.n61 585
R1066 B.n636 B.n635 585
R1067 B.n637 B.n60 585
R1068 B.n639 B.n638 585
R1069 B.n640 B.n59 585
R1070 B.n642 B.n641 585
R1071 B.n643 B.n58 585
R1072 B.n645 B.n644 585
R1073 B.n647 B.n55 585
R1074 B.n649 B.n648 585
R1075 B.n650 B.n54 585
R1076 B.n652 B.n651 585
R1077 B.n653 B.n53 585
R1078 B.n655 B.n654 585
R1079 B.n656 B.n52 585
R1080 B.n658 B.n657 585
R1081 B.n659 B.n49 585
R1082 B.n662 B.n661 585
R1083 B.n663 B.n48 585
R1084 B.n665 B.n664 585
R1085 B.n666 B.n47 585
R1086 B.n668 B.n667 585
R1087 B.n669 B.n46 585
R1088 B.n671 B.n670 585
R1089 B.n672 B.n45 585
R1090 B.n674 B.n673 585
R1091 B.n675 B.n44 585
R1092 B.n677 B.n676 585
R1093 B.n678 B.n43 585
R1094 B.n680 B.n679 585
R1095 B.n681 B.n42 585
R1096 B.n683 B.n682 585
R1097 B.n684 B.n41 585
R1098 B.n686 B.n685 585
R1099 B.n687 B.n40 585
R1100 B.n689 B.n688 585
R1101 B.n690 B.n39 585
R1102 B.n692 B.n691 585
R1103 B.n693 B.n38 585
R1104 B.n695 B.n694 585
R1105 B.n696 B.n37 585
R1106 B.n698 B.n697 585
R1107 B.n699 B.n36 585
R1108 B.n701 B.n700 585
R1109 B.n702 B.n35 585
R1110 B.n704 B.n703 585
R1111 B.n705 B.n34 585
R1112 B.n707 B.n706 585
R1113 B.n708 B.n33 585
R1114 B.n710 B.n709 585
R1115 B.n711 B.n32 585
R1116 B.n713 B.n712 585
R1117 B.n714 B.n31 585
R1118 B.n716 B.n715 585
R1119 B.n717 B.n30 585
R1120 B.n719 B.n718 585
R1121 B.n720 B.n29 585
R1122 B.n722 B.n721 585
R1123 B.n723 B.n28 585
R1124 B.n582 B.n581 585
R1125 B.n580 B.n79 585
R1126 B.n579 B.n578 585
R1127 B.n577 B.n80 585
R1128 B.n576 B.n575 585
R1129 B.n574 B.n81 585
R1130 B.n573 B.n572 585
R1131 B.n571 B.n82 585
R1132 B.n570 B.n569 585
R1133 B.n568 B.n83 585
R1134 B.n567 B.n566 585
R1135 B.n565 B.n84 585
R1136 B.n564 B.n563 585
R1137 B.n562 B.n85 585
R1138 B.n561 B.n560 585
R1139 B.n559 B.n86 585
R1140 B.n558 B.n557 585
R1141 B.n556 B.n87 585
R1142 B.n555 B.n554 585
R1143 B.n553 B.n88 585
R1144 B.n552 B.n551 585
R1145 B.n550 B.n89 585
R1146 B.n549 B.n548 585
R1147 B.n547 B.n90 585
R1148 B.n546 B.n545 585
R1149 B.n544 B.n91 585
R1150 B.n543 B.n542 585
R1151 B.n541 B.n92 585
R1152 B.n540 B.n539 585
R1153 B.n538 B.n93 585
R1154 B.n537 B.n536 585
R1155 B.n535 B.n94 585
R1156 B.n534 B.n533 585
R1157 B.n532 B.n95 585
R1158 B.n531 B.n530 585
R1159 B.n529 B.n96 585
R1160 B.n528 B.n527 585
R1161 B.n526 B.n97 585
R1162 B.n525 B.n524 585
R1163 B.n523 B.n98 585
R1164 B.n522 B.n521 585
R1165 B.n520 B.n99 585
R1166 B.n519 B.n518 585
R1167 B.n517 B.n100 585
R1168 B.n516 B.n515 585
R1169 B.n514 B.n101 585
R1170 B.n513 B.n512 585
R1171 B.n511 B.n102 585
R1172 B.n510 B.n509 585
R1173 B.n508 B.n103 585
R1174 B.n507 B.n506 585
R1175 B.n505 B.n104 585
R1176 B.n504 B.n503 585
R1177 B.n502 B.n105 585
R1178 B.n501 B.n500 585
R1179 B.n499 B.n106 585
R1180 B.n498 B.n497 585
R1181 B.n496 B.n107 585
R1182 B.n495 B.n494 585
R1183 B.n493 B.n108 585
R1184 B.n492 B.n491 585
R1185 B.n490 B.n109 585
R1186 B.n489 B.n488 585
R1187 B.n487 B.n110 585
R1188 B.n486 B.n485 585
R1189 B.n484 B.n111 585
R1190 B.n483 B.n482 585
R1191 B.n481 B.n112 585
R1192 B.n480 B.n479 585
R1193 B.n478 B.n113 585
R1194 B.n477 B.n476 585
R1195 B.n475 B.n114 585
R1196 B.n474 B.n473 585
R1197 B.n472 B.n115 585
R1198 B.n471 B.n470 585
R1199 B.n469 B.n116 585
R1200 B.n468 B.n467 585
R1201 B.n466 B.n117 585
R1202 B.n465 B.n464 585
R1203 B.n463 B.n118 585
R1204 B.n462 B.n461 585
R1205 B.n460 B.n119 585
R1206 B.n459 B.n458 585
R1207 B.n457 B.n120 585
R1208 B.n456 B.n455 585
R1209 B.n454 B.n121 585
R1210 B.n453 B.n452 585
R1211 B.n451 B.n122 585
R1212 B.n450 B.n449 585
R1213 B.n448 B.n123 585
R1214 B.n447 B.n446 585
R1215 B.n445 B.n124 585
R1216 B.n444 B.n443 585
R1217 B.n442 B.n125 585
R1218 B.n441 B.n440 585
R1219 B.n439 B.n126 585
R1220 B.n438 B.n437 585
R1221 B.n436 B.n127 585
R1222 B.n435 B.n434 585
R1223 B.n433 B.n128 585
R1224 B.n432 B.n431 585
R1225 B.n430 B.n129 585
R1226 B.n429 B.n428 585
R1227 B.n427 B.n130 585
R1228 B.n426 B.n425 585
R1229 B.n285 B.n284 585
R1230 B.n286 B.n181 585
R1231 B.n288 B.n287 585
R1232 B.n289 B.n180 585
R1233 B.n291 B.n290 585
R1234 B.n292 B.n179 585
R1235 B.n294 B.n293 585
R1236 B.n295 B.n178 585
R1237 B.n297 B.n296 585
R1238 B.n298 B.n177 585
R1239 B.n300 B.n299 585
R1240 B.n301 B.n176 585
R1241 B.n303 B.n302 585
R1242 B.n304 B.n175 585
R1243 B.n306 B.n305 585
R1244 B.n307 B.n174 585
R1245 B.n309 B.n308 585
R1246 B.n310 B.n173 585
R1247 B.n312 B.n311 585
R1248 B.n313 B.n172 585
R1249 B.n315 B.n314 585
R1250 B.n316 B.n171 585
R1251 B.n318 B.n317 585
R1252 B.n319 B.n170 585
R1253 B.n321 B.n320 585
R1254 B.n322 B.n169 585
R1255 B.n324 B.n323 585
R1256 B.n325 B.n168 585
R1257 B.n327 B.n326 585
R1258 B.n328 B.n167 585
R1259 B.n330 B.n329 585
R1260 B.n331 B.n166 585
R1261 B.n333 B.n332 585
R1262 B.n334 B.n165 585
R1263 B.n336 B.n335 585
R1264 B.n337 B.n164 585
R1265 B.n339 B.n338 585
R1266 B.n340 B.n163 585
R1267 B.n342 B.n341 585
R1268 B.n343 B.n162 585
R1269 B.n345 B.n344 585
R1270 B.n346 B.n159 585
R1271 B.n349 B.n348 585
R1272 B.n350 B.n158 585
R1273 B.n352 B.n351 585
R1274 B.n353 B.n157 585
R1275 B.n355 B.n354 585
R1276 B.n356 B.n156 585
R1277 B.n358 B.n357 585
R1278 B.n359 B.n155 585
R1279 B.n361 B.n360 585
R1280 B.n363 B.n362 585
R1281 B.n364 B.n151 585
R1282 B.n366 B.n365 585
R1283 B.n367 B.n150 585
R1284 B.n369 B.n368 585
R1285 B.n370 B.n149 585
R1286 B.n372 B.n371 585
R1287 B.n373 B.n148 585
R1288 B.n375 B.n374 585
R1289 B.n376 B.n147 585
R1290 B.n378 B.n377 585
R1291 B.n379 B.n146 585
R1292 B.n381 B.n380 585
R1293 B.n382 B.n145 585
R1294 B.n384 B.n383 585
R1295 B.n385 B.n144 585
R1296 B.n387 B.n386 585
R1297 B.n388 B.n143 585
R1298 B.n390 B.n389 585
R1299 B.n391 B.n142 585
R1300 B.n393 B.n392 585
R1301 B.n394 B.n141 585
R1302 B.n396 B.n395 585
R1303 B.n397 B.n140 585
R1304 B.n399 B.n398 585
R1305 B.n400 B.n139 585
R1306 B.n402 B.n401 585
R1307 B.n403 B.n138 585
R1308 B.n405 B.n404 585
R1309 B.n406 B.n137 585
R1310 B.n408 B.n407 585
R1311 B.n409 B.n136 585
R1312 B.n411 B.n410 585
R1313 B.n412 B.n135 585
R1314 B.n414 B.n413 585
R1315 B.n415 B.n134 585
R1316 B.n417 B.n416 585
R1317 B.n418 B.n133 585
R1318 B.n420 B.n419 585
R1319 B.n421 B.n132 585
R1320 B.n423 B.n422 585
R1321 B.n424 B.n131 585
R1322 B.n283 B.n182 585
R1323 B.n282 B.n281 585
R1324 B.n280 B.n183 585
R1325 B.n279 B.n278 585
R1326 B.n277 B.n184 585
R1327 B.n276 B.n275 585
R1328 B.n274 B.n185 585
R1329 B.n273 B.n272 585
R1330 B.n271 B.n186 585
R1331 B.n270 B.n269 585
R1332 B.n268 B.n187 585
R1333 B.n267 B.n266 585
R1334 B.n265 B.n188 585
R1335 B.n264 B.n263 585
R1336 B.n262 B.n189 585
R1337 B.n261 B.n260 585
R1338 B.n259 B.n190 585
R1339 B.n258 B.n257 585
R1340 B.n256 B.n191 585
R1341 B.n255 B.n254 585
R1342 B.n253 B.n192 585
R1343 B.n252 B.n251 585
R1344 B.n250 B.n193 585
R1345 B.n249 B.n248 585
R1346 B.n247 B.n194 585
R1347 B.n246 B.n245 585
R1348 B.n244 B.n195 585
R1349 B.n243 B.n242 585
R1350 B.n241 B.n196 585
R1351 B.n240 B.n239 585
R1352 B.n238 B.n197 585
R1353 B.n237 B.n236 585
R1354 B.n235 B.n198 585
R1355 B.n234 B.n233 585
R1356 B.n232 B.n199 585
R1357 B.n231 B.n230 585
R1358 B.n229 B.n200 585
R1359 B.n228 B.n227 585
R1360 B.n226 B.n201 585
R1361 B.n225 B.n224 585
R1362 B.n223 B.n202 585
R1363 B.n222 B.n221 585
R1364 B.n220 B.n203 585
R1365 B.n219 B.n218 585
R1366 B.n217 B.n204 585
R1367 B.n216 B.n215 585
R1368 B.n214 B.n205 585
R1369 B.n213 B.n212 585
R1370 B.n211 B.n206 585
R1371 B.n210 B.n209 585
R1372 B.n208 B.n207 585
R1373 B.n2 B.n0 585
R1374 B.n801 B.n1 585
R1375 B.n800 B.n799 585
R1376 B.n798 B.n3 585
R1377 B.n797 B.n796 585
R1378 B.n795 B.n4 585
R1379 B.n794 B.n793 585
R1380 B.n792 B.n5 585
R1381 B.n791 B.n790 585
R1382 B.n789 B.n6 585
R1383 B.n788 B.n787 585
R1384 B.n786 B.n7 585
R1385 B.n785 B.n784 585
R1386 B.n783 B.n8 585
R1387 B.n782 B.n781 585
R1388 B.n780 B.n9 585
R1389 B.n779 B.n778 585
R1390 B.n777 B.n10 585
R1391 B.n776 B.n775 585
R1392 B.n774 B.n11 585
R1393 B.n773 B.n772 585
R1394 B.n771 B.n12 585
R1395 B.n770 B.n769 585
R1396 B.n768 B.n13 585
R1397 B.n767 B.n766 585
R1398 B.n765 B.n14 585
R1399 B.n764 B.n763 585
R1400 B.n762 B.n15 585
R1401 B.n761 B.n760 585
R1402 B.n759 B.n16 585
R1403 B.n758 B.n757 585
R1404 B.n756 B.n17 585
R1405 B.n755 B.n754 585
R1406 B.n753 B.n18 585
R1407 B.n752 B.n751 585
R1408 B.n750 B.n19 585
R1409 B.n749 B.n748 585
R1410 B.n747 B.n20 585
R1411 B.n746 B.n745 585
R1412 B.n744 B.n21 585
R1413 B.n743 B.n742 585
R1414 B.n741 B.n22 585
R1415 B.n740 B.n739 585
R1416 B.n738 B.n23 585
R1417 B.n737 B.n736 585
R1418 B.n735 B.n24 585
R1419 B.n734 B.n733 585
R1420 B.n732 B.n25 585
R1421 B.n731 B.n730 585
R1422 B.n729 B.n26 585
R1423 B.n728 B.n727 585
R1424 B.n726 B.n27 585
R1425 B.n725 B.n724 585
R1426 B.n803 B.n802 585
R1427 B.n284 B.n283 535.745
R1428 B.n724 B.n723 535.745
R1429 B.n426 B.n131 535.745
R1430 B.n583 B.n582 535.745
R1431 B.n152 B.t8 434.293
R1432 B.n56 B.t10 434.293
R1433 B.n160 B.t2 434.293
R1434 B.n50 B.t4 434.293
R1435 B.n153 B.t7 376.111
R1436 B.n57 B.t11 376.111
R1437 B.n161 B.t1 376.111
R1438 B.n51 B.t5 376.111
R1439 B.n152 B.t6 316.736
R1440 B.n160 B.t0 316.736
R1441 B.n50 B.t3 316.736
R1442 B.n56 B.t9 316.736
R1443 B.n283 B.n282 163.367
R1444 B.n282 B.n183 163.367
R1445 B.n278 B.n183 163.367
R1446 B.n278 B.n277 163.367
R1447 B.n277 B.n276 163.367
R1448 B.n276 B.n185 163.367
R1449 B.n272 B.n185 163.367
R1450 B.n272 B.n271 163.367
R1451 B.n271 B.n270 163.367
R1452 B.n270 B.n187 163.367
R1453 B.n266 B.n187 163.367
R1454 B.n266 B.n265 163.367
R1455 B.n265 B.n264 163.367
R1456 B.n264 B.n189 163.367
R1457 B.n260 B.n189 163.367
R1458 B.n260 B.n259 163.367
R1459 B.n259 B.n258 163.367
R1460 B.n258 B.n191 163.367
R1461 B.n254 B.n191 163.367
R1462 B.n254 B.n253 163.367
R1463 B.n253 B.n252 163.367
R1464 B.n252 B.n193 163.367
R1465 B.n248 B.n193 163.367
R1466 B.n248 B.n247 163.367
R1467 B.n247 B.n246 163.367
R1468 B.n246 B.n195 163.367
R1469 B.n242 B.n195 163.367
R1470 B.n242 B.n241 163.367
R1471 B.n241 B.n240 163.367
R1472 B.n240 B.n197 163.367
R1473 B.n236 B.n197 163.367
R1474 B.n236 B.n235 163.367
R1475 B.n235 B.n234 163.367
R1476 B.n234 B.n199 163.367
R1477 B.n230 B.n199 163.367
R1478 B.n230 B.n229 163.367
R1479 B.n229 B.n228 163.367
R1480 B.n228 B.n201 163.367
R1481 B.n224 B.n201 163.367
R1482 B.n224 B.n223 163.367
R1483 B.n223 B.n222 163.367
R1484 B.n222 B.n203 163.367
R1485 B.n218 B.n203 163.367
R1486 B.n218 B.n217 163.367
R1487 B.n217 B.n216 163.367
R1488 B.n216 B.n205 163.367
R1489 B.n212 B.n205 163.367
R1490 B.n212 B.n211 163.367
R1491 B.n211 B.n210 163.367
R1492 B.n210 B.n207 163.367
R1493 B.n207 B.n2 163.367
R1494 B.n802 B.n2 163.367
R1495 B.n802 B.n801 163.367
R1496 B.n801 B.n800 163.367
R1497 B.n800 B.n3 163.367
R1498 B.n796 B.n3 163.367
R1499 B.n796 B.n795 163.367
R1500 B.n795 B.n794 163.367
R1501 B.n794 B.n5 163.367
R1502 B.n790 B.n5 163.367
R1503 B.n790 B.n789 163.367
R1504 B.n789 B.n788 163.367
R1505 B.n788 B.n7 163.367
R1506 B.n784 B.n7 163.367
R1507 B.n784 B.n783 163.367
R1508 B.n783 B.n782 163.367
R1509 B.n782 B.n9 163.367
R1510 B.n778 B.n9 163.367
R1511 B.n778 B.n777 163.367
R1512 B.n777 B.n776 163.367
R1513 B.n776 B.n11 163.367
R1514 B.n772 B.n11 163.367
R1515 B.n772 B.n771 163.367
R1516 B.n771 B.n770 163.367
R1517 B.n770 B.n13 163.367
R1518 B.n766 B.n13 163.367
R1519 B.n766 B.n765 163.367
R1520 B.n765 B.n764 163.367
R1521 B.n764 B.n15 163.367
R1522 B.n760 B.n15 163.367
R1523 B.n760 B.n759 163.367
R1524 B.n759 B.n758 163.367
R1525 B.n758 B.n17 163.367
R1526 B.n754 B.n17 163.367
R1527 B.n754 B.n753 163.367
R1528 B.n753 B.n752 163.367
R1529 B.n752 B.n19 163.367
R1530 B.n748 B.n19 163.367
R1531 B.n748 B.n747 163.367
R1532 B.n747 B.n746 163.367
R1533 B.n746 B.n21 163.367
R1534 B.n742 B.n21 163.367
R1535 B.n742 B.n741 163.367
R1536 B.n741 B.n740 163.367
R1537 B.n740 B.n23 163.367
R1538 B.n736 B.n23 163.367
R1539 B.n736 B.n735 163.367
R1540 B.n735 B.n734 163.367
R1541 B.n734 B.n25 163.367
R1542 B.n730 B.n25 163.367
R1543 B.n730 B.n729 163.367
R1544 B.n729 B.n728 163.367
R1545 B.n728 B.n27 163.367
R1546 B.n724 B.n27 163.367
R1547 B.n284 B.n181 163.367
R1548 B.n288 B.n181 163.367
R1549 B.n289 B.n288 163.367
R1550 B.n290 B.n289 163.367
R1551 B.n290 B.n179 163.367
R1552 B.n294 B.n179 163.367
R1553 B.n295 B.n294 163.367
R1554 B.n296 B.n295 163.367
R1555 B.n296 B.n177 163.367
R1556 B.n300 B.n177 163.367
R1557 B.n301 B.n300 163.367
R1558 B.n302 B.n301 163.367
R1559 B.n302 B.n175 163.367
R1560 B.n306 B.n175 163.367
R1561 B.n307 B.n306 163.367
R1562 B.n308 B.n307 163.367
R1563 B.n308 B.n173 163.367
R1564 B.n312 B.n173 163.367
R1565 B.n313 B.n312 163.367
R1566 B.n314 B.n313 163.367
R1567 B.n314 B.n171 163.367
R1568 B.n318 B.n171 163.367
R1569 B.n319 B.n318 163.367
R1570 B.n320 B.n319 163.367
R1571 B.n320 B.n169 163.367
R1572 B.n324 B.n169 163.367
R1573 B.n325 B.n324 163.367
R1574 B.n326 B.n325 163.367
R1575 B.n326 B.n167 163.367
R1576 B.n330 B.n167 163.367
R1577 B.n331 B.n330 163.367
R1578 B.n332 B.n331 163.367
R1579 B.n332 B.n165 163.367
R1580 B.n336 B.n165 163.367
R1581 B.n337 B.n336 163.367
R1582 B.n338 B.n337 163.367
R1583 B.n338 B.n163 163.367
R1584 B.n342 B.n163 163.367
R1585 B.n343 B.n342 163.367
R1586 B.n344 B.n343 163.367
R1587 B.n344 B.n159 163.367
R1588 B.n349 B.n159 163.367
R1589 B.n350 B.n349 163.367
R1590 B.n351 B.n350 163.367
R1591 B.n351 B.n157 163.367
R1592 B.n355 B.n157 163.367
R1593 B.n356 B.n355 163.367
R1594 B.n357 B.n356 163.367
R1595 B.n357 B.n155 163.367
R1596 B.n361 B.n155 163.367
R1597 B.n362 B.n361 163.367
R1598 B.n362 B.n151 163.367
R1599 B.n366 B.n151 163.367
R1600 B.n367 B.n366 163.367
R1601 B.n368 B.n367 163.367
R1602 B.n368 B.n149 163.367
R1603 B.n372 B.n149 163.367
R1604 B.n373 B.n372 163.367
R1605 B.n374 B.n373 163.367
R1606 B.n374 B.n147 163.367
R1607 B.n378 B.n147 163.367
R1608 B.n379 B.n378 163.367
R1609 B.n380 B.n379 163.367
R1610 B.n380 B.n145 163.367
R1611 B.n384 B.n145 163.367
R1612 B.n385 B.n384 163.367
R1613 B.n386 B.n385 163.367
R1614 B.n386 B.n143 163.367
R1615 B.n390 B.n143 163.367
R1616 B.n391 B.n390 163.367
R1617 B.n392 B.n391 163.367
R1618 B.n392 B.n141 163.367
R1619 B.n396 B.n141 163.367
R1620 B.n397 B.n396 163.367
R1621 B.n398 B.n397 163.367
R1622 B.n398 B.n139 163.367
R1623 B.n402 B.n139 163.367
R1624 B.n403 B.n402 163.367
R1625 B.n404 B.n403 163.367
R1626 B.n404 B.n137 163.367
R1627 B.n408 B.n137 163.367
R1628 B.n409 B.n408 163.367
R1629 B.n410 B.n409 163.367
R1630 B.n410 B.n135 163.367
R1631 B.n414 B.n135 163.367
R1632 B.n415 B.n414 163.367
R1633 B.n416 B.n415 163.367
R1634 B.n416 B.n133 163.367
R1635 B.n420 B.n133 163.367
R1636 B.n421 B.n420 163.367
R1637 B.n422 B.n421 163.367
R1638 B.n422 B.n131 163.367
R1639 B.n427 B.n426 163.367
R1640 B.n428 B.n427 163.367
R1641 B.n428 B.n129 163.367
R1642 B.n432 B.n129 163.367
R1643 B.n433 B.n432 163.367
R1644 B.n434 B.n433 163.367
R1645 B.n434 B.n127 163.367
R1646 B.n438 B.n127 163.367
R1647 B.n439 B.n438 163.367
R1648 B.n440 B.n439 163.367
R1649 B.n440 B.n125 163.367
R1650 B.n444 B.n125 163.367
R1651 B.n445 B.n444 163.367
R1652 B.n446 B.n445 163.367
R1653 B.n446 B.n123 163.367
R1654 B.n450 B.n123 163.367
R1655 B.n451 B.n450 163.367
R1656 B.n452 B.n451 163.367
R1657 B.n452 B.n121 163.367
R1658 B.n456 B.n121 163.367
R1659 B.n457 B.n456 163.367
R1660 B.n458 B.n457 163.367
R1661 B.n458 B.n119 163.367
R1662 B.n462 B.n119 163.367
R1663 B.n463 B.n462 163.367
R1664 B.n464 B.n463 163.367
R1665 B.n464 B.n117 163.367
R1666 B.n468 B.n117 163.367
R1667 B.n469 B.n468 163.367
R1668 B.n470 B.n469 163.367
R1669 B.n470 B.n115 163.367
R1670 B.n474 B.n115 163.367
R1671 B.n475 B.n474 163.367
R1672 B.n476 B.n475 163.367
R1673 B.n476 B.n113 163.367
R1674 B.n480 B.n113 163.367
R1675 B.n481 B.n480 163.367
R1676 B.n482 B.n481 163.367
R1677 B.n482 B.n111 163.367
R1678 B.n486 B.n111 163.367
R1679 B.n487 B.n486 163.367
R1680 B.n488 B.n487 163.367
R1681 B.n488 B.n109 163.367
R1682 B.n492 B.n109 163.367
R1683 B.n493 B.n492 163.367
R1684 B.n494 B.n493 163.367
R1685 B.n494 B.n107 163.367
R1686 B.n498 B.n107 163.367
R1687 B.n499 B.n498 163.367
R1688 B.n500 B.n499 163.367
R1689 B.n500 B.n105 163.367
R1690 B.n504 B.n105 163.367
R1691 B.n505 B.n504 163.367
R1692 B.n506 B.n505 163.367
R1693 B.n506 B.n103 163.367
R1694 B.n510 B.n103 163.367
R1695 B.n511 B.n510 163.367
R1696 B.n512 B.n511 163.367
R1697 B.n512 B.n101 163.367
R1698 B.n516 B.n101 163.367
R1699 B.n517 B.n516 163.367
R1700 B.n518 B.n517 163.367
R1701 B.n518 B.n99 163.367
R1702 B.n522 B.n99 163.367
R1703 B.n523 B.n522 163.367
R1704 B.n524 B.n523 163.367
R1705 B.n524 B.n97 163.367
R1706 B.n528 B.n97 163.367
R1707 B.n529 B.n528 163.367
R1708 B.n530 B.n529 163.367
R1709 B.n530 B.n95 163.367
R1710 B.n534 B.n95 163.367
R1711 B.n535 B.n534 163.367
R1712 B.n536 B.n535 163.367
R1713 B.n536 B.n93 163.367
R1714 B.n540 B.n93 163.367
R1715 B.n541 B.n540 163.367
R1716 B.n542 B.n541 163.367
R1717 B.n542 B.n91 163.367
R1718 B.n546 B.n91 163.367
R1719 B.n547 B.n546 163.367
R1720 B.n548 B.n547 163.367
R1721 B.n548 B.n89 163.367
R1722 B.n552 B.n89 163.367
R1723 B.n553 B.n552 163.367
R1724 B.n554 B.n553 163.367
R1725 B.n554 B.n87 163.367
R1726 B.n558 B.n87 163.367
R1727 B.n559 B.n558 163.367
R1728 B.n560 B.n559 163.367
R1729 B.n560 B.n85 163.367
R1730 B.n564 B.n85 163.367
R1731 B.n565 B.n564 163.367
R1732 B.n566 B.n565 163.367
R1733 B.n566 B.n83 163.367
R1734 B.n570 B.n83 163.367
R1735 B.n571 B.n570 163.367
R1736 B.n572 B.n571 163.367
R1737 B.n572 B.n81 163.367
R1738 B.n576 B.n81 163.367
R1739 B.n577 B.n576 163.367
R1740 B.n578 B.n577 163.367
R1741 B.n578 B.n79 163.367
R1742 B.n582 B.n79 163.367
R1743 B.n723 B.n722 163.367
R1744 B.n722 B.n29 163.367
R1745 B.n718 B.n29 163.367
R1746 B.n718 B.n717 163.367
R1747 B.n717 B.n716 163.367
R1748 B.n716 B.n31 163.367
R1749 B.n712 B.n31 163.367
R1750 B.n712 B.n711 163.367
R1751 B.n711 B.n710 163.367
R1752 B.n710 B.n33 163.367
R1753 B.n706 B.n33 163.367
R1754 B.n706 B.n705 163.367
R1755 B.n705 B.n704 163.367
R1756 B.n704 B.n35 163.367
R1757 B.n700 B.n35 163.367
R1758 B.n700 B.n699 163.367
R1759 B.n699 B.n698 163.367
R1760 B.n698 B.n37 163.367
R1761 B.n694 B.n37 163.367
R1762 B.n694 B.n693 163.367
R1763 B.n693 B.n692 163.367
R1764 B.n692 B.n39 163.367
R1765 B.n688 B.n39 163.367
R1766 B.n688 B.n687 163.367
R1767 B.n687 B.n686 163.367
R1768 B.n686 B.n41 163.367
R1769 B.n682 B.n41 163.367
R1770 B.n682 B.n681 163.367
R1771 B.n681 B.n680 163.367
R1772 B.n680 B.n43 163.367
R1773 B.n676 B.n43 163.367
R1774 B.n676 B.n675 163.367
R1775 B.n675 B.n674 163.367
R1776 B.n674 B.n45 163.367
R1777 B.n670 B.n45 163.367
R1778 B.n670 B.n669 163.367
R1779 B.n669 B.n668 163.367
R1780 B.n668 B.n47 163.367
R1781 B.n664 B.n47 163.367
R1782 B.n664 B.n663 163.367
R1783 B.n663 B.n662 163.367
R1784 B.n662 B.n49 163.367
R1785 B.n657 B.n49 163.367
R1786 B.n657 B.n656 163.367
R1787 B.n656 B.n655 163.367
R1788 B.n655 B.n53 163.367
R1789 B.n651 B.n53 163.367
R1790 B.n651 B.n650 163.367
R1791 B.n650 B.n649 163.367
R1792 B.n649 B.n55 163.367
R1793 B.n644 B.n55 163.367
R1794 B.n644 B.n643 163.367
R1795 B.n643 B.n642 163.367
R1796 B.n642 B.n59 163.367
R1797 B.n638 B.n59 163.367
R1798 B.n638 B.n637 163.367
R1799 B.n637 B.n636 163.367
R1800 B.n636 B.n61 163.367
R1801 B.n632 B.n61 163.367
R1802 B.n632 B.n631 163.367
R1803 B.n631 B.n630 163.367
R1804 B.n630 B.n63 163.367
R1805 B.n626 B.n63 163.367
R1806 B.n626 B.n625 163.367
R1807 B.n625 B.n624 163.367
R1808 B.n624 B.n65 163.367
R1809 B.n620 B.n65 163.367
R1810 B.n620 B.n619 163.367
R1811 B.n619 B.n618 163.367
R1812 B.n618 B.n67 163.367
R1813 B.n614 B.n67 163.367
R1814 B.n614 B.n613 163.367
R1815 B.n613 B.n612 163.367
R1816 B.n612 B.n69 163.367
R1817 B.n608 B.n69 163.367
R1818 B.n608 B.n607 163.367
R1819 B.n607 B.n606 163.367
R1820 B.n606 B.n71 163.367
R1821 B.n602 B.n71 163.367
R1822 B.n602 B.n601 163.367
R1823 B.n601 B.n600 163.367
R1824 B.n600 B.n73 163.367
R1825 B.n596 B.n73 163.367
R1826 B.n596 B.n595 163.367
R1827 B.n595 B.n594 163.367
R1828 B.n594 B.n75 163.367
R1829 B.n590 B.n75 163.367
R1830 B.n590 B.n589 163.367
R1831 B.n589 B.n588 163.367
R1832 B.n588 B.n77 163.367
R1833 B.n584 B.n77 163.367
R1834 B.n584 B.n583 163.367
R1835 B.n154 B.n153 59.5399
R1836 B.n347 B.n161 59.5399
R1837 B.n660 B.n51 59.5399
R1838 B.n646 B.n57 59.5399
R1839 B.n153 B.n152 58.1823
R1840 B.n161 B.n160 58.1823
R1841 B.n51 B.n50 58.1823
R1842 B.n57 B.n56 58.1823
R1843 B.n725 B.n28 34.8103
R1844 B.n581 B.n78 34.8103
R1845 B.n425 B.n424 34.8103
R1846 B.n285 B.n182 34.8103
R1847 B B.n803 18.0485
R1848 B.n721 B.n28 10.6151
R1849 B.n721 B.n720 10.6151
R1850 B.n720 B.n719 10.6151
R1851 B.n719 B.n30 10.6151
R1852 B.n715 B.n30 10.6151
R1853 B.n715 B.n714 10.6151
R1854 B.n714 B.n713 10.6151
R1855 B.n713 B.n32 10.6151
R1856 B.n709 B.n32 10.6151
R1857 B.n709 B.n708 10.6151
R1858 B.n708 B.n707 10.6151
R1859 B.n707 B.n34 10.6151
R1860 B.n703 B.n34 10.6151
R1861 B.n703 B.n702 10.6151
R1862 B.n702 B.n701 10.6151
R1863 B.n701 B.n36 10.6151
R1864 B.n697 B.n36 10.6151
R1865 B.n697 B.n696 10.6151
R1866 B.n696 B.n695 10.6151
R1867 B.n695 B.n38 10.6151
R1868 B.n691 B.n38 10.6151
R1869 B.n691 B.n690 10.6151
R1870 B.n690 B.n689 10.6151
R1871 B.n689 B.n40 10.6151
R1872 B.n685 B.n40 10.6151
R1873 B.n685 B.n684 10.6151
R1874 B.n684 B.n683 10.6151
R1875 B.n683 B.n42 10.6151
R1876 B.n679 B.n42 10.6151
R1877 B.n679 B.n678 10.6151
R1878 B.n678 B.n677 10.6151
R1879 B.n677 B.n44 10.6151
R1880 B.n673 B.n44 10.6151
R1881 B.n673 B.n672 10.6151
R1882 B.n672 B.n671 10.6151
R1883 B.n671 B.n46 10.6151
R1884 B.n667 B.n46 10.6151
R1885 B.n667 B.n666 10.6151
R1886 B.n666 B.n665 10.6151
R1887 B.n665 B.n48 10.6151
R1888 B.n661 B.n48 10.6151
R1889 B.n659 B.n658 10.6151
R1890 B.n658 B.n52 10.6151
R1891 B.n654 B.n52 10.6151
R1892 B.n654 B.n653 10.6151
R1893 B.n653 B.n652 10.6151
R1894 B.n652 B.n54 10.6151
R1895 B.n648 B.n54 10.6151
R1896 B.n648 B.n647 10.6151
R1897 B.n645 B.n58 10.6151
R1898 B.n641 B.n58 10.6151
R1899 B.n641 B.n640 10.6151
R1900 B.n640 B.n639 10.6151
R1901 B.n639 B.n60 10.6151
R1902 B.n635 B.n60 10.6151
R1903 B.n635 B.n634 10.6151
R1904 B.n634 B.n633 10.6151
R1905 B.n633 B.n62 10.6151
R1906 B.n629 B.n62 10.6151
R1907 B.n629 B.n628 10.6151
R1908 B.n628 B.n627 10.6151
R1909 B.n627 B.n64 10.6151
R1910 B.n623 B.n64 10.6151
R1911 B.n623 B.n622 10.6151
R1912 B.n622 B.n621 10.6151
R1913 B.n621 B.n66 10.6151
R1914 B.n617 B.n66 10.6151
R1915 B.n617 B.n616 10.6151
R1916 B.n616 B.n615 10.6151
R1917 B.n615 B.n68 10.6151
R1918 B.n611 B.n68 10.6151
R1919 B.n611 B.n610 10.6151
R1920 B.n610 B.n609 10.6151
R1921 B.n609 B.n70 10.6151
R1922 B.n605 B.n70 10.6151
R1923 B.n605 B.n604 10.6151
R1924 B.n604 B.n603 10.6151
R1925 B.n603 B.n72 10.6151
R1926 B.n599 B.n72 10.6151
R1927 B.n599 B.n598 10.6151
R1928 B.n598 B.n597 10.6151
R1929 B.n597 B.n74 10.6151
R1930 B.n593 B.n74 10.6151
R1931 B.n593 B.n592 10.6151
R1932 B.n592 B.n591 10.6151
R1933 B.n591 B.n76 10.6151
R1934 B.n587 B.n76 10.6151
R1935 B.n587 B.n586 10.6151
R1936 B.n586 B.n585 10.6151
R1937 B.n585 B.n78 10.6151
R1938 B.n425 B.n130 10.6151
R1939 B.n429 B.n130 10.6151
R1940 B.n430 B.n429 10.6151
R1941 B.n431 B.n430 10.6151
R1942 B.n431 B.n128 10.6151
R1943 B.n435 B.n128 10.6151
R1944 B.n436 B.n435 10.6151
R1945 B.n437 B.n436 10.6151
R1946 B.n437 B.n126 10.6151
R1947 B.n441 B.n126 10.6151
R1948 B.n442 B.n441 10.6151
R1949 B.n443 B.n442 10.6151
R1950 B.n443 B.n124 10.6151
R1951 B.n447 B.n124 10.6151
R1952 B.n448 B.n447 10.6151
R1953 B.n449 B.n448 10.6151
R1954 B.n449 B.n122 10.6151
R1955 B.n453 B.n122 10.6151
R1956 B.n454 B.n453 10.6151
R1957 B.n455 B.n454 10.6151
R1958 B.n455 B.n120 10.6151
R1959 B.n459 B.n120 10.6151
R1960 B.n460 B.n459 10.6151
R1961 B.n461 B.n460 10.6151
R1962 B.n461 B.n118 10.6151
R1963 B.n465 B.n118 10.6151
R1964 B.n466 B.n465 10.6151
R1965 B.n467 B.n466 10.6151
R1966 B.n467 B.n116 10.6151
R1967 B.n471 B.n116 10.6151
R1968 B.n472 B.n471 10.6151
R1969 B.n473 B.n472 10.6151
R1970 B.n473 B.n114 10.6151
R1971 B.n477 B.n114 10.6151
R1972 B.n478 B.n477 10.6151
R1973 B.n479 B.n478 10.6151
R1974 B.n479 B.n112 10.6151
R1975 B.n483 B.n112 10.6151
R1976 B.n484 B.n483 10.6151
R1977 B.n485 B.n484 10.6151
R1978 B.n485 B.n110 10.6151
R1979 B.n489 B.n110 10.6151
R1980 B.n490 B.n489 10.6151
R1981 B.n491 B.n490 10.6151
R1982 B.n491 B.n108 10.6151
R1983 B.n495 B.n108 10.6151
R1984 B.n496 B.n495 10.6151
R1985 B.n497 B.n496 10.6151
R1986 B.n497 B.n106 10.6151
R1987 B.n501 B.n106 10.6151
R1988 B.n502 B.n501 10.6151
R1989 B.n503 B.n502 10.6151
R1990 B.n503 B.n104 10.6151
R1991 B.n507 B.n104 10.6151
R1992 B.n508 B.n507 10.6151
R1993 B.n509 B.n508 10.6151
R1994 B.n509 B.n102 10.6151
R1995 B.n513 B.n102 10.6151
R1996 B.n514 B.n513 10.6151
R1997 B.n515 B.n514 10.6151
R1998 B.n515 B.n100 10.6151
R1999 B.n519 B.n100 10.6151
R2000 B.n520 B.n519 10.6151
R2001 B.n521 B.n520 10.6151
R2002 B.n521 B.n98 10.6151
R2003 B.n525 B.n98 10.6151
R2004 B.n526 B.n525 10.6151
R2005 B.n527 B.n526 10.6151
R2006 B.n527 B.n96 10.6151
R2007 B.n531 B.n96 10.6151
R2008 B.n532 B.n531 10.6151
R2009 B.n533 B.n532 10.6151
R2010 B.n533 B.n94 10.6151
R2011 B.n537 B.n94 10.6151
R2012 B.n538 B.n537 10.6151
R2013 B.n539 B.n538 10.6151
R2014 B.n539 B.n92 10.6151
R2015 B.n543 B.n92 10.6151
R2016 B.n544 B.n543 10.6151
R2017 B.n545 B.n544 10.6151
R2018 B.n545 B.n90 10.6151
R2019 B.n549 B.n90 10.6151
R2020 B.n550 B.n549 10.6151
R2021 B.n551 B.n550 10.6151
R2022 B.n551 B.n88 10.6151
R2023 B.n555 B.n88 10.6151
R2024 B.n556 B.n555 10.6151
R2025 B.n557 B.n556 10.6151
R2026 B.n557 B.n86 10.6151
R2027 B.n561 B.n86 10.6151
R2028 B.n562 B.n561 10.6151
R2029 B.n563 B.n562 10.6151
R2030 B.n563 B.n84 10.6151
R2031 B.n567 B.n84 10.6151
R2032 B.n568 B.n567 10.6151
R2033 B.n569 B.n568 10.6151
R2034 B.n569 B.n82 10.6151
R2035 B.n573 B.n82 10.6151
R2036 B.n574 B.n573 10.6151
R2037 B.n575 B.n574 10.6151
R2038 B.n575 B.n80 10.6151
R2039 B.n579 B.n80 10.6151
R2040 B.n580 B.n579 10.6151
R2041 B.n581 B.n580 10.6151
R2042 B.n286 B.n285 10.6151
R2043 B.n287 B.n286 10.6151
R2044 B.n287 B.n180 10.6151
R2045 B.n291 B.n180 10.6151
R2046 B.n292 B.n291 10.6151
R2047 B.n293 B.n292 10.6151
R2048 B.n293 B.n178 10.6151
R2049 B.n297 B.n178 10.6151
R2050 B.n298 B.n297 10.6151
R2051 B.n299 B.n298 10.6151
R2052 B.n299 B.n176 10.6151
R2053 B.n303 B.n176 10.6151
R2054 B.n304 B.n303 10.6151
R2055 B.n305 B.n304 10.6151
R2056 B.n305 B.n174 10.6151
R2057 B.n309 B.n174 10.6151
R2058 B.n310 B.n309 10.6151
R2059 B.n311 B.n310 10.6151
R2060 B.n311 B.n172 10.6151
R2061 B.n315 B.n172 10.6151
R2062 B.n316 B.n315 10.6151
R2063 B.n317 B.n316 10.6151
R2064 B.n317 B.n170 10.6151
R2065 B.n321 B.n170 10.6151
R2066 B.n322 B.n321 10.6151
R2067 B.n323 B.n322 10.6151
R2068 B.n323 B.n168 10.6151
R2069 B.n327 B.n168 10.6151
R2070 B.n328 B.n327 10.6151
R2071 B.n329 B.n328 10.6151
R2072 B.n329 B.n166 10.6151
R2073 B.n333 B.n166 10.6151
R2074 B.n334 B.n333 10.6151
R2075 B.n335 B.n334 10.6151
R2076 B.n335 B.n164 10.6151
R2077 B.n339 B.n164 10.6151
R2078 B.n340 B.n339 10.6151
R2079 B.n341 B.n340 10.6151
R2080 B.n341 B.n162 10.6151
R2081 B.n345 B.n162 10.6151
R2082 B.n346 B.n345 10.6151
R2083 B.n348 B.n158 10.6151
R2084 B.n352 B.n158 10.6151
R2085 B.n353 B.n352 10.6151
R2086 B.n354 B.n353 10.6151
R2087 B.n354 B.n156 10.6151
R2088 B.n358 B.n156 10.6151
R2089 B.n359 B.n358 10.6151
R2090 B.n360 B.n359 10.6151
R2091 B.n364 B.n363 10.6151
R2092 B.n365 B.n364 10.6151
R2093 B.n365 B.n150 10.6151
R2094 B.n369 B.n150 10.6151
R2095 B.n370 B.n369 10.6151
R2096 B.n371 B.n370 10.6151
R2097 B.n371 B.n148 10.6151
R2098 B.n375 B.n148 10.6151
R2099 B.n376 B.n375 10.6151
R2100 B.n377 B.n376 10.6151
R2101 B.n377 B.n146 10.6151
R2102 B.n381 B.n146 10.6151
R2103 B.n382 B.n381 10.6151
R2104 B.n383 B.n382 10.6151
R2105 B.n383 B.n144 10.6151
R2106 B.n387 B.n144 10.6151
R2107 B.n388 B.n387 10.6151
R2108 B.n389 B.n388 10.6151
R2109 B.n389 B.n142 10.6151
R2110 B.n393 B.n142 10.6151
R2111 B.n394 B.n393 10.6151
R2112 B.n395 B.n394 10.6151
R2113 B.n395 B.n140 10.6151
R2114 B.n399 B.n140 10.6151
R2115 B.n400 B.n399 10.6151
R2116 B.n401 B.n400 10.6151
R2117 B.n401 B.n138 10.6151
R2118 B.n405 B.n138 10.6151
R2119 B.n406 B.n405 10.6151
R2120 B.n407 B.n406 10.6151
R2121 B.n407 B.n136 10.6151
R2122 B.n411 B.n136 10.6151
R2123 B.n412 B.n411 10.6151
R2124 B.n413 B.n412 10.6151
R2125 B.n413 B.n134 10.6151
R2126 B.n417 B.n134 10.6151
R2127 B.n418 B.n417 10.6151
R2128 B.n419 B.n418 10.6151
R2129 B.n419 B.n132 10.6151
R2130 B.n423 B.n132 10.6151
R2131 B.n424 B.n423 10.6151
R2132 B.n281 B.n182 10.6151
R2133 B.n281 B.n280 10.6151
R2134 B.n280 B.n279 10.6151
R2135 B.n279 B.n184 10.6151
R2136 B.n275 B.n184 10.6151
R2137 B.n275 B.n274 10.6151
R2138 B.n274 B.n273 10.6151
R2139 B.n273 B.n186 10.6151
R2140 B.n269 B.n186 10.6151
R2141 B.n269 B.n268 10.6151
R2142 B.n268 B.n267 10.6151
R2143 B.n267 B.n188 10.6151
R2144 B.n263 B.n188 10.6151
R2145 B.n263 B.n262 10.6151
R2146 B.n262 B.n261 10.6151
R2147 B.n261 B.n190 10.6151
R2148 B.n257 B.n190 10.6151
R2149 B.n257 B.n256 10.6151
R2150 B.n256 B.n255 10.6151
R2151 B.n255 B.n192 10.6151
R2152 B.n251 B.n192 10.6151
R2153 B.n251 B.n250 10.6151
R2154 B.n250 B.n249 10.6151
R2155 B.n249 B.n194 10.6151
R2156 B.n245 B.n194 10.6151
R2157 B.n245 B.n244 10.6151
R2158 B.n244 B.n243 10.6151
R2159 B.n243 B.n196 10.6151
R2160 B.n239 B.n196 10.6151
R2161 B.n239 B.n238 10.6151
R2162 B.n238 B.n237 10.6151
R2163 B.n237 B.n198 10.6151
R2164 B.n233 B.n198 10.6151
R2165 B.n233 B.n232 10.6151
R2166 B.n232 B.n231 10.6151
R2167 B.n231 B.n200 10.6151
R2168 B.n227 B.n200 10.6151
R2169 B.n227 B.n226 10.6151
R2170 B.n226 B.n225 10.6151
R2171 B.n225 B.n202 10.6151
R2172 B.n221 B.n202 10.6151
R2173 B.n221 B.n220 10.6151
R2174 B.n220 B.n219 10.6151
R2175 B.n219 B.n204 10.6151
R2176 B.n215 B.n204 10.6151
R2177 B.n215 B.n214 10.6151
R2178 B.n214 B.n213 10.6151
R2179 B.n213 B.n206 10.6151
R2180 B.n209 B.n206 10.6151
R2181 B.n209 B.n208 10.6151
R2182 B.n208 B.n0 10.6151
R2183 B.n799 B.n1 10.6151
R2184 B.n799 B.n798 10.6151
R2185 B.n798 B.n797 10.6151
R2186 B.n797 B.n4 10.6151
R2187 B.n793 B.n4 10.6151
R2188 B.n793 B.n792 10.6151
R2189 B.n792 B.n791 10.6151
R2190 B.n791 B.n6 10.6151
R2191 B.n787 B.n6 10.6151
R2192 B.n787 B.n786 10.6151
R2193 B.n786 B.n785 10.6151
R2194 B.n785 B.n8 10.6151
R2195 B.n781 B.n8 10.6151
R2196 B.n781 B.n780 10.6151
R2197 B.n780 B.n779 10.6151
R2198 B.n779 B.n10 10.6151
R2199 B.n775 B.n10 10.6151
R2200 B.n775 B.n774 10.6151
R2201 B.n774 B.n773 10.6151
R2202 B.n773 B.n12 10.6151
R2203 B.n769 B.n12 10.6151
R2204 B.n769 B.n768 10.6151
R2205 B.n768 B.n767 10.6151
R2206 B.n767 B.n14 10.6151
R2207 B.n763 B.n14 10.6151
R2208 B.n763 B.n762 10.6151
R2209 B.n762 B.n761 10.6151
R2210 B.n761 B.n16 10.6151
R2211 B.n757 B.n16 10.6151
R2212 B.n757 B.n756 10.6151
R2213 B.n756 B.n755 10.6151
R2214 B.n755 B.n18 10.6151
R2215 B.n751 B.n18 10.6151
R2216 B.n751 B.n750 10.6151
R2217 B.n750 B.n749 10.6151
R2218 B.n749 B.n20 10.6151
R2219 B.n745 B.n20 10.6151
R2220 B.n745 B.n744 10.6151
R2221 B.n744 B.n743 10.6151
R2222 B.n743 B.n22 10.6151
R2223 B.n739 B.n22 10.6151
R2224 B.n739 B.n738 10.6151
R2225 B.n738 B.n737 10.6151
R2226 B.n737 B.n24 10.6151
R2227 B.n733 B.n24 10.6151
R2228 B.n733 B.n732 10.6151
R2229 B.n732 B.n731 10.6151
R2230 B.n731 B.n26 10.6151
R2231 B.n727 B.n26 10.6151
R2232 B.n727 B.n726 10.6151
R2233 B.n726 B.n725 10.6151
R2234 B.n660 B.n659 6.5566
R2235 B.n647 B.n646 6.5566
R2236 B.n348 B.n347 6.5566
R2237 B.n360 B.n154 6.5566
R2238 B.n661 B.n660 4.05904
R2239 B.n646 B.n645 4.05904
R2240 B.n347 B.n346 4.05904
R2241 B.n363 B.n154 4.05904
R2242 B.n803 B.n0 2.81026
R2243 B.n803 B.n1 2.81026
C0 VTAIL w_n3970_n3374# 4.21654f
C1 B VDD1 1.6705f
C2 w_n3970_n3374# VP 8.633551f
C3 VTAIL VP 9.19348f
C4 VN B 1.24187f
C5 B VDD2 1.76873f
C6 w_n3970_n3374# B 10.2315f
C7 VTAIL B 5.02509f
C8 B VP 2.10655f
C9 VN VDD1 0.151361f
C10 VDD1 VDD2 1.81036f
C11 VN VDD2 8.76905f
C12 w_n3970_n3374# VDD1 1.97077f
C13 VTAIL VDD1 8.10263f
C14 VN w_n3970_n3374# 8.11796f
C15 VN VTAIL 9.17937f
C16 w_n3970_n3374# VDD2 2.08841f
C17 VTAIL VDD2 8.15751f
C18 VP VDD1 9.14289f
C19 VN VP 7.75819f
C20 VP VDD2 0.526626f
C21 VDD2 VSUBS 1.93309f
C22 VDD1 VSUBS 2.471109f
C23 VTAIL VSUBS 1.350221f
C24 VN VSUBS 6.84855f
C25 VP VSUBS 3.67176f
C26 B VSUBS 5.08649f
C27 w_n3970_n3374# VSUBS 0.164882p
C28 B.n0 VSUBS 0.004781f
C29 B.n1 VSUBS 0.004781f
C30 B.n2 VSUBS 0.007561f
C31 B.n3 VSUBS 0.007561f
C32 B.n4 VSUBS 0.007561f
C33 B.n5 VSUBS 0.007561f
C34 B.n6 VSUBS 0.007561f
C35 B.n7 VSUBS 0.007561f
C36 B.n8 VSUBS 0.007561f
C37 B.n9 VSUBS 0.007561f
C38 B.n10 VSUBS 0.007561f
C39 B.n11 VSUBS 0.007561f
C40 B.n12 VSUBS 0.007561f
C41 B.n13 VSUBS 0.007561f
C42 B.n14 VSUBS 0.007561f
C43 B.n15 VSUBS 0.007561f
C44 B.n16 VSUBS 0.007561f
C45 B.n17 VSUBS 0.007561f
C46 B.n18 VSUBS 0.007561f
C47 B.n19 VSUBS 0.007561f
C48 B.n20 VSUBS 0.007561f
C49 B.n21 VSUBS 0.007561f
C50 B.n22 VSUBS 0.007561f
C51 B.n23 VSUBS 0.007561f
C52 B.n24 VSUBS 0.007561f
C53 B.n25 VSUBS 0.007561f
C54 B.n26 VSUBS 0.007561f
C55 B.n27 VSUBS 0.007561f
C56 B.n28 VSUBS 0.019021f
C57 B.n29 VSUBS 0.007561f
C58 B.n30 VSUBS 0.007561f
C59 B.n31 VSUBS 0.007561f
C60 B.n32 VSUBS 0.007561f
C61 B.n33 VSUBS 0.007561f
C62 B.n34 VSUBS 0.007561f
C63 B.n35 VSUBS 0.007561f
C64 B.n36 VSUBS 0.007561f
C65 B.n37 VSUBS 0.007561f
C66 B.n38 VSUBS 0.007561f
C67 B.n39 VSUBS 0.007561f
C68 B.n40 VSUBS 0.007561f
C69 B.n41 VSUBS 0.007561f
C70 B.n42 VSUBS 0.007561f
C71 B.n43 VSUBS 0.007561f
C72 B.n44 VSUBS 0.007561f
C73 B.n45 VSUBS 0.007561f
C74 B.n46 VSUBS 0.007561f
C75 B.n47 VSUBS 0.007561f
C76 B.n48 VSUBS 0.007561f
C77 B.n49 VSUBS 0.007561f
C78 B.t5 VSUBS 0.228589f
C79 B.t4 VSUBS 0.263701f
C80 B.t3 VSUBS 1.58291f
C81 B.n50 VSUBS 0.419075f
C82 B.n51 VSUBS 0.27287f
C83 B.n52 VSUBS 0.007561f
C84 B.n53 VSUBS 0.007561f
C85 B.n54 VSUBS 0.007561f
C86 B.n55 VSUBS 0.007561f
C87 B.t11 VSUBS 0.228592f
C88 B.t10 VSUBS 0.263703f
C89 B.t9 VSUBS 1.58291f
C90 B.n56 VSUBS 0.419072f
C91 B.n57 VSUBS 0.272867f
C92 B.n58 VSUBS 0.007561f
C93 B.n59 VSUBS 0.007561f
C94 B.n60 VSUBS 0.007561f
C95 B.n61 VSUBS 0.007561f
C96 B.n62 VSUBS 0.007561f
C97 B.n63 VSUBS 0.007561f
C98 B.n64 VSUBS 0.007561f
C99 B.n65 VSUBS 0.007561f
C100 B.n66 VSUBS 0.007561f
C101 B.n67 VSUBS 0.007561f
C102 B.n68 VSUBS 0.007561f
C103 B.n69 VSUBS 0.007561f
C104 B.n70 VSUBS 0.007561f
C105 B.n71 VSUBS 0.007561f
C106 B.n72 VSUBS 0.007561f
C107 B.n73 VSUBS 0.007561f
C108 B.n74 VSUBS 0.007561f
C109 B.n75 VSUBS 0.007561f
C110 B.n76 VSUBS 0.007561f
C111 B.n77 VSUBS 0.007561f
C112 B.n78 VSUBS 0.018182f
C113 B.n79 VSUBS 0.007561f
C114 B.n80 VSUBS 0.007561f
C115 B.n81 VSUBS 0.007561f
C116 B.n82 VSUBS 0.007561f
C117 B.n83 VSUBS 0.007561f
C118 B.n84 VSUBS 0.007561f
C119 B.n85 VSUBS 0.007561f
C120 B.n86 VSUBS 0.007561f
C121 B.n87 VSUBS 0.007561f
C122 B.n88 VSUBS 0.007561f
C123 B.n89 VSUBS 0.007561f
C124 B.n90 VSUBS 0.007561f
C125 B.n91 VSUBS 0.007561f
C126 B.n92 VSUBS 0.007561f
C127 B.n93 VSUBS 0.007561f
C128 B.n94 VSUBS 0.007561f
C129 B.n95 VSUBS 0.007561f
C130 B.n96 VSUBS 0.007561f
C131 B.n97 VSUBS 0.007561f
C132 B.n98 VSUBS 0.007561f
C133 B.n99 VSUBS 0.007561f
C134 B.n100 VSUBS 0.007561f
C135 B.n101 VSUBS 0.007561f
C136 B.n102 VSUBS 0.007561f
C137 B.n103 VSUBS 0.007561f
C138 B.n104 VSUBS 0.007561f
C139 B.n105 VSUBS 0.007561f
C140 B.n106 VSUBS 0.007561f
C141 B.n107 VSUBS 0.007561f
C142 B.n108 VSUBS 0.007561f
C143 B.n109 VSUBS 0.007561f
C144 B.n110 VSUBS 0.007561f
C145 B.n111 VSUBS 0.007561f
C146 B.n112 VSUBS 0.007561f
C147 B.n113 VSUBS 0.007561f
C148 B.n114 VSUBS 0.007561f
C149 B.n115 VSUBS 0.007561f
C150 B.n116 VSUBS 0.007561f
C151 B.n117 VSUBS 0.007561f
C152 B.n118 VSUBS 0.007561f
C153 B.n119 VSUBS 0.007561f
C154 B.n120 VSUBS 0.007561f
C155 B.n121 VSUBS 0.007561f
C156 B.n122 VSUBS 0.007561f
C157 B.n123 VSUBS 0.007561f
C158 B.n124 VSUBS 0.007561f
C159 B.n125 VSUBS 0.007561f
C160 B.n126 VSUBS 0.007561f
C161 B.n127 VSUBS 0.007561f
C162 B.n128 VSUBS 0.007561f
C163 B.n129 VSUBS 0.007561f
C164 B.n130 VSUBS 0.007561f
C165 B.n131 VSUBS 0.019021f
C166 B.n132 VSUBS 0.007561f
C167 B.n133 VSUBS 0.007561f
C168 B.n134 VSUBS 0.007561f
C169 B.n135 VSUBS 0.007561f
C170 B.n136 VSUBS 0.007561f
C171 B.n137 VSUBS 0.007561f
C172 B.n138 VSUBS 0.007561f
C173 B.n139 VSUBS 0.007561f
C174 B.n140 VSUBS 0.007561f
C175 B.n141 VSUBS 0.007561f
C176 B.n142 VSUBS 0.007561f
C177 B.n143 VSUBS 0.007561f
C178 B.n144 VSUBS 0.007561f
C179 B.n145 VSUBS 0.007561f
C180 B.n146 VSUBS 0.007561f
C181 B.n147 VSUBS 0.007561f
C182 B.n148 VSUBS 0.007561f
C183 B.n149 VSUBS 0.007561f
C184 B.n150 VSUBS 0.007561f
C185 B.n151 VSUBS 0.007561f
C186 B.t7 VSUBS 0.228592f
C187 B.t8 VSUBS 0.263703f
C188 B.t6 VSUBS 1.58291f
C189 B.n152 VSUBS 0.419072f
C190 B.n153 VSUBS 0.272867f
C191 B.n154 VSUBS 0.017519f
C192 B.n155 VSUBS 0.007561f
C193 B.n156 VSUBS 0.007561f
C194 B.n157 VSUBS 0.007561f
C195 B.n158 VSUBS 0.007561f
C196 B.n159 VSUBS 0.007561f
C197 B.t1 VSUBS 0.228589f
C198 B.t2 VSUBS 0.263701f
C199 B.t0 VSUBS 1.58291f
C200 B.n160 VSUBS 0.419075f
C201 B.n161 VSUBS 0.27287f
C202 B.n162 VSUBS 0.007561f
C203 B.n163 VSUBS 0.007561f
C204 B.n164 VSUBS 0.007561f
C205 B.n165 VSUBS 0.007561f
C206 B.n166 VSUBS 0.007561f
C207 B.n167 VSUBS 0.007561f
C208 B.n168 VSUBS 0.007561f
C209 B.n169 VSUBS 0.007561f
C210 B.n170 VSUBS 0.007561f
C211 B.n171 VSUBS 0.007561f
C212 B.n172 VSUBS 0.007561f
C213 B.n173 VSUBS 0.007561f
C214 B.n174 VSUBS 0.007561f
C215 B.n175 VSUBS 0.007561f
C216 B.n176 VSUBS 0.007561f
C217 B.n177 VSUBS 0.007561f
C218 B.n178 VSUBS 0.007561f
C219 B.n179 VSUBS 0.007561f
C220 B.n180 VSUBS 0.007561f
C221 B.n181 VSUBS 0.007561f
C222 B.n182 VSUBS 0.017896f
C223 B.n183 VSUBS 0.007561f
C224 B.n184 VSUBS 0.007561f
C225 B.n185 VSUBS 0.007561f
C226 B.n186 VSUBS 0.007561f
C227 B.n187 VSUBS 0.007561f
C228 B.n188 VSUBS 0.007561f
C229 B.n189 VSUBS 0.007561f
C230 B.n190 VSUBS 0.007561f
C231 B.n191 VSUBS 0.007561f
C232 B.n192 VSUBS 0.007561f
C233 B.n193 VSUBS 0.007561f
C234 B.n194 VSUBS 0.007561f
C235 B.n195 VSUBS 0.007561f
C236 B.n196 VSUBS 0.007561f
C237 B.n197 VSUBS 0.007561f
C238 B.n198 VSUBS 0.007561f
C239 B.n199 VSUBS 0.007561f
C240 B.n200 VSUBS 0.007561f
C241 B.n201 VSUBS 0.007561f
C242 B.n202 VSUBS 0.007561f
C243 B.n203 VSUBS 0.007561f
C244 B.n204 VSUBS 0.007561f
C245 B.n205 VSUBS 0.007561f
C246 B.n206 VSUBS 0.007561f
C247 B.n207 VSUBS 0.007561f
C248 B.n208 VSUBS 0.007561f
C249 B.n209 VSUBS 0.007561f
C250 B.n210 VSUBS 0.007561f
C251 B.n211 VSUBS 0.007561f
C252 B.n212 VSUBS 0.007561f
C253 B.n213 VSUBS 0.007561f
C254 B.n214 VSUBS 0.007561f
C255 B.n215 VSUBS 0.007561f
C256 B.n216 VSUBS 0.007561f
C257 B.n217 VSUBS 0.007561f
C258 B.n218 VSUBS 0.007561f
C259 B.n219 VSUBS 0.007561f
C260 B.n220 VSUBS 0.007561f
C261 B.n221 VSUBS 0.007561f
C262 B.n222 VSUBS 0.007561f
C263 B.n223 VSUBS 0.007561f
C264 B.n224 VSUBS 0.007561f
C265 B.n225 VSUBS 0.007561f
C266 B.n226 VSUBS 0.007561f
C267 B.n227 VSUBS 0.007561f
C268 B.n228 VSUBS 0.007561f
C269 B.n229 VSUBS 0.007561f
C270 B.n230 VSUBS 0.007561f
C271 B.n231 VSUBS 0.007561f
C272 B.n232 VSUBS 0.007561f
C273 B.n233 VSUBS 0.007561f
C274 B.n234 VSUBS 0.007561f
C275 B.n235 VSUBS 0.007561f
C276 B.n236 VSUBS 0.007561f
C277 B.n237 VSUBS 0.007561f
C278 B.n238 VSUBS 0.007561f
C279 B.n239 VSUBS 0.007561f
C280 B.n240 VSUBS 0.007561f
C281 B.n241 VSUBS 0.007561f
C282 B.n242 VSUBS 0.007561f
C283 B.n243 VSUBS 0.007561f
C284 B.n244 VSUBS 0.007561f
C285 B.n245 VSUBS 0.007561f
C286 B.n246 VSUBS 0.007561f
C287 B.n247 VSUBS 0.007561f
C288 B.n248 VSUBS 0.007561f
C289 B.n249 VSUBS 0.007561f
C290 B.n250 VSUBS 0.007561f
C291 B.n251 VSUBS 0.007561f
C292 B.n252 VSUBS 0.007561f
C293 B.n253 VSUBS 0.007561f
C294 B.n254 VSUBS 0.007561f
C295 B.n255 VSUBS 0.007561f
C296 B.n256 VSUBS 0.007561f
C297 B.n257 VSUBS 0.007561f
C298 B.n258 VSUBS 0.007561f
C299 B.n259 VSUBS 0.007561f
C300 B.n260 VSUBS 0.007561f
C301 B.n261 VSUBS 0.007561f
C302 B.n262 VSUBS 0.007561f
C303 B.n263 VSUBS 0.007561f
C304 B.n264 VSUBS 0.007561f
C305 B.n265 VSUBS 0.007561f
C306 B.n266 VSUBS 0.007561f
C307 B.n267 VSUBS 0.007561f
C308 B.n268 VSUBS 0.007561f
C309 B.n269 VSUBS 0.007561f
C310 B.n270 VSUBS 0.007561f
C311 B.n271 VSUBS 0.007561f
C312 B.n272 VSUBS 0.007561f
C313 B.n273 VSUBS 0.007561f
C314 B.n274 VSUBS 0.007561f
C315 B.n275 VSUBS 0.007561f
C316 B.n276 VSUBS 0.007561f
C317 B.n277 VSUBS 0.007561f
C318 B.n278 VSUBS 0.007561f
C319 B.n279 VSUBS 0.007561f
C320 B.n280 VSUBS 0.007561f
C321 B.n281 VSUBS 0.007561f
C322 B.n282 VSUBS 0.007561f
C323 B.n283 VSUBS 0.017896f
C324 B.n284 VSUBS 0.019021f
C325 B.n285 VSUBS 0.019021f
C326 B.n286 VSUBS 0.007561f
C327 B.n287 VSUBS 0.007561f
C328 B.n288 VSUBS 0.007561f
C329 B.n289 VSUBS 0.007561f
C330 B.n290 VSUBS 0.007561f
C331 B.n291 VSUBS 0.007561f
C332 B.n292 VSUBS 0.007561f
C333 B.n293 VSUBS 0.007561f
C334 B.n294 VSUBS 0.007561f
C335 B.n295 VSUBS 0.007561f
C336 B.n296 VSUBS 0.007561f
C337 B.n297 VSUBS 0.007561f
C338 B.n298 VSUBS 0.007561f
C339 B.n299 VSUBS 0.007561f
C340 B.n300 VSUBS 0.007561f
C341 B.n301 VSUBS 0.007561f
C342 B.n302 VSUBS 0.007561f
C343 B.n303 VSUBS 0.007561f
C344 B.n304 VSUBS 0.007561f
C345 B.n305 VSUBS 0.007561f
C346 B.n306 VSUBS 0.007561f
C347 B.n307 VSUBS 0.007561f
C348 B.n308 VSUBS 0.007561f
C349 B.n309 VSUBS 0.007561f
C350 B.n310 VSUBS 0.007561f
C351 B.n311 VSUBS 0.007561f
C352 B.n312 VSUBS 0.007561f
C353 B.n313 VSUBS 0.007561f
C354 B.n314 VSUBS 0.007561f
C355 B.n315 VSUBS 0.007561f
C356 B.n316 VSUBS 0.007561f
C357 B.n317 VSUBS 0.007561f
C358 B.n318 VSUBS 0.007561f
C359 B.n319 VSUBS 0.007561f
C360 B.n320 VSUBS 0.007561f
C361 B.n321 VSUBS 0.007561f
C362 B.n322 VSUBS 0.007561f
C363 B.n323 VSUBS 0.007561f
C364 B.n324 VSUBS 0.007561f
C365 B.n325 VSUBS 0.007561f
C366 B.n326 VSUBS 0.007561f
C367 B.n327 VSUBS 0.007561f
C368 B.n328 VSUBS 0.007561f
C369 B.n329 VSUBS 0.007561f
C370 B.n330 VSUBS 0.007561f
C371 B.n331 VSUBS 0.007561f
C372 B.n332 VSUBS 0.007561f
C373 B.n333 VSUBS 0.007561f
C374 B.n334 VSUBS 0.007561f
C375 B.n335 VSUBS 0.007561f
C376 B.n336 VSUBS 0.007561f
C377 B.n337 VSUBS 0.007561f
C378 B.n338 VSUBS 0.007561f
C379 B.n339 VSUBS 0.007561f
C380 B.n340 VSUBS 0.007561f
C381 B.n341 VSUBS 0.007561f
C382 B.n342 VSUBS 0.007561f
C383 B.n343 VSUBS 0.007561f
C384 B.n344 VSUBS 0.007561f
C385 B.n345 VSUBS 0.007561f
C386 B.n346 VSUBS 0.005226f
C387 B.n347 VSUBS 0.017519f
C388 B.n348 VSUBS 0.006116f
C389 B.n349 VSUBS 0.007561f
C390 B.n350 VSUBS 0.007561f
C391 B.n351 VSUBS 0.007561f
C392 B.n352 VSUBS 0.007561f
C393 B.n353 VSUBS 0.007561f
C394 B.n354 VSUBS 0.007561f
C395 B.n355 VSUBS 0.007561f
C396 B.n356 VSUBS 0.007561f
C397 B.n357 VSUBS 0.007561f
C398 B.n358 VSUBS 0.007561f
C399 B.n359 VSUBS 0.007561f
C400 B.n360 VSUBS 0.006116f
C401 B.n361 VSUBS 0.007561f
C402 B.n362 VSUBS 0.007561f
C403 B.n363 VSUBS 0.005226f
C404 B.n364 VSUBS 0.007561f
C405 B.n365 VSUBS 0.007561f
C406 B.n366 VSUBS 0.007561f
C407 B.n367 VSUBS 0.007561f
C408 B.n368 VSUBS 0.007561f
C409 B.n369 VSUBS 0.007561f
C410 B.n370 VSUBS 0.007561f
C411 B.n371 VSUBS 0.007561f
C412 B.n372 VSUBS 0.007561f
C413 B.n373 VSUBS 0.007561f
C414 B.n374 VSUBS 0.007561f
C415 B.n375 VSUBS 0.007561f
C416 B.n376 VSUBS 0.007561f
C417 B.n377 VSUBS 0.007561f
C418 B.n378 VSUBS 0.007561f
C419 B.n379 VSUBS 0.007561f
C420 B.n380 VSUBS 0.007561f
C421 B.n381 VSUBS 0.007561f
C422 B.n382 VSUBS 0.007561f
C423 B.n383 VSUBS 0.007561f
C424 B.n384 VSUBS 0.007561f
C425 B.n385 VSUBS 0.007561f
C426 B.n386 VSUBS 0.007561f
C427 B.n387 VSUBS 0.007561f
C428 B.n388 VSUBS 0.007561f
C429 B.n389 VSUBS 0.007561f
C430 B.n390 VSUBS 0.007561f
C431 B.n391 VSUBS 0.007561f
C432 B.n392 VSUBS 0.007561f
C433 B.n393 VSUBS 0.007561f
C434 B.n394 VSUBS 0.007561f
C435 B.n395 VSUBS 0.007561f
C436 B.n396 VSUBS 0.007561f
C437 B.n397 VSUBS 0.007561f
C438 B.n398 VSUBS 0.007561f
C439 B.n399 VSUBS 0.007561f
C440 B.n400 VSUBS 0.007561f
C441 B.n401 VSUBS 0.007561f
C442 B.n402 VSUBS 0.007561f
C443 B.n403 VSUBS 0.007561f
C444 B.n404 VSUBS 0.007561f
C445 B.n405 VSUBS 0.007561f
C446 B.n406 VSUBS 0.007561f
C447 B.n407 VSUBS 0.007561f
C448 B.n408 VSUBS 0.007561f
C449 B.n409 VSUBS 0.007561f
C450 B.n410 VSUBS 0.007561f
C451 B.n411 VSUBS 0.007561f
C452 B.n412 VSUBS 0.007561f
C453 B.n413 VSUBS 0.007561f
C454 B.n414 VSUBS 0.007561f
C455 B.n415 VSUBS 0.007561f
C456 B.n416 VSUBS 0.007561f
C457 B.n417 VSUBS 0.007561f
C458 B.n418 VSUBS 0.007561f
C459 B.n419 VSUBS 0.007561f
C460 B.n420 VSUBS 0.007561f
C461 B.n421 VSUBS 0.007561f
C462 B.n422 VSUBS 0.007561f
C463 B.n423 VSUBS 0.007561f
C464 B.n424 VSUBS 0.019021f
C465 B.n425 VSUBS 0.017896f
C466 B.n426 VSUBS 0.017896f
C467 B.n427 VSUBS 0.007561f
C468 B.n428 VSUBS 0.007561f
C469 B.n429 VSUBS 0.007561f
C470 B.n430 VSUBS 0.007561f
C471 B.n431 VSUBS 0.007561f
C472 B.n432 VSUBS 0.007561f
C473 B.n433 VSUBS 0.007561f
C474 B.n434 VSUBS 0.007561f
C475 B.n435 VSUBS 0.007561f
C476 B.n436 VSUBS 0.007561f
C477 B.n437 VSUBS 0.007561f
C478 B.n438 VSUBS 0.007561f
C479 B.n439 VSUBS 0.007561f
C480 B.n440 VSUBS 0.007561f
C481 B.n441 VSUBS 0.007561f
C482 B.n442 VSUBS 0.007561f
C483 B.n443 VSUBS 0.007561f
C484 B.n444 VSUBS 0.007561f
C485 B.n445 VSUBS 0.007561f
C486 B.n446 VSUBS 0.007561f
C487 B.n447 VSUBS 0.007561f
C488 B.n448 VSUBS 0.007561f
C489 B.n449 VSUBS 0.007561f
C490 B.n450 VSUBS 0.007561f
C491 B.n451 VSUBS 0.007561f
C492 B.n452 VSUBS 0.007561f
C493 B.n453 VSUBS 0.007561f
C494 B.n454 VSUBS 0.007561f
C495 B.n455 VSUBS 0.007561f
C496 B.n456 VSUBS 0.007561f
C497 B.n457 VSUBS 0.007561f
C498 B.n458 VSUBS 0.007561f
C499 B.n459 VSUBS 0.007561f
C500 B.n460 VSUBS 0.007561f
C501 B.n461 VSUBS 0.007561f
C502 B.n462 VSUBS 0.007561f
C503 B.n463 VSUBS 0.007561f
C504 B.n464 VSUBS 0.007561f
C505 B.n465 VSUBS 0.007561f
C506 B.n466 VSUBS 0.007561f
C507 B.n467 VSUBS 0.007561f
C508 B.n468 VSUBS 0.007561f
C509 B.n469 VSUBS 0.007561f
C510 B.n470 VSUBS 0.007561f
C511 B.n471 VSUBS 0.007561f
C512 B.n472 VSUBS 0.007561f
C513 B.n473 VSUBS 0.007561f
C514 B.n474 VSUBS 0.007561f
C515 B.n475 VSUBS 0.007561f
C516 B.n476 VSUBS 0.007561f
C517 B.n477 VSUBS 0.007561f
C518 B.n478 VSUBS 0.007561f
C519 B.n479 VSUBS 0.007561f
C520 B.n480 VSUBS 0.007561f
C521 B.n481 VSUBS 0.007561f
C522 B.n482 VSUBS 0.007561f
C523 B.n483 VSUBS 0.007561f
C524 B.n484 VSUBS 0.007561f
C525 B.n485 VSUBS 0.007561f
C526 B.n486 VSUBS 0.007561f
C527 B.n487 VSUBS 0.007561f
C528 B.n488 VSUBS 0.007561f
C529 B.n489 VSUBS 0.007561f
C530 B.n490 VSUBS 0.007561f
C531 B.n491 VSUBS 0.007561f
C532 B.n492 VSUBS 0.007561f
C533 B.n493 VSUBS 0.007561f
C534 B.n494 VSUBS 0.007561f
C535 B.n495 VSUBS 0.007561f
C536 B.n496 VSUBS 0.007561f
C537 B.n497 VSUBS 0.007561f
C538 B.n498 VSUBS 0.007561f
C539 B.n499 VSUBS 0.007561f
C540 B.n500 VSUBS 0.007561f
C541 B.n501 VSUBS 0.007561f
C542 B.n502 VSUBS 0.007561f
C543 B.n503 VSUBS 0.007561f
C544 B.n504 VSUBS 0.007561f
C545 B.n505 VSUBS 0.007561f
C546 B.n506 VSUBS 0.007561f
C547 B.n507 VSUBS 0.007561f
C548 B.n508 VSUBS 0.007561f
C549 B.n509 VSUBS 0.007561f
C550 B.n510 VSUBS 0.007561f
C551 B.n511 VSUBS 0.007561f
C552 B.n512 VSUBS 0.007561f
C553 B.n513 VSUBS 0.007561f
C554 B.n514 VSUBS 0.007561f
C555 B.n515 VSUBS 0.007561f
C556 B.n516 VSUBS 0.007561f
C557 B.n517 VSUBS 0.007561f
C558 B.n518 VSUBS 0.007561f
C559 B.n519 VSUBS 0.007561f
C560 B.n520 VSUBS 0.007561f
C561 B.n521 VSUBS 0.007561f
C562 B.n522 VSUBS 0.007561f
C563 B.n523 VSUBS 0.007561f
C564 B.n524 VSUBS 0.007561f
C565 B.n525 VSUBS 0.007561f
C566 B.n526 VSUBS 0.007561f
C567 B.n527 VSUBS 0.007561f
C568 B.n528 VSUBS 0.007561f
C569 B.n529 VSUBS 0.007561f
C570 B.n530 VSUBS 0.007561f
C571 B.n531 VSUBS 0.007561f
C572 B.n532 VSUBS 0.007561f
C573 B.n533 VSUBS 0.007561f
C574 B.n534 VSUBS 0.007561f
C575 B.n535 VSUBS 0.007561f
C576 B.n536 VSUBS 0.007561f
C577 B.n537 VSUBS 0.007561f
C578 B.n538 VSUBS 0.007561f
C579 B.n539 VSUBS 0.007561f
C580 B.n540 VSUBS 0.007561f
C581 B.n541 VSUBS 0.007561f
C582 B.n542 VSUBS 0.007561f
C583 B.n543 VSUBS 0.007561f
C584 B.n544 VSUBS 0.007561f
C585 B.n545 VSUBS 0.007561f
C586 B.n546 VSUBS 0.007561f
C587 B.n547 VSUBS 0.007561f
C588 B.n548 VSUBS 0.007561f
C589 B.n549 VSUBS 0.007561f
C590 B.n550 VSUBS 0.007561f
C591 B.n551 VSUBS 0.007561f
C592 B.n552 VSUBS 0.007561f
C593 B.n553 VSUBS 0.007561f
C594 B.n554 VSUBS 0.007561f
C595 B.n555 VSUBS 0.007561f
C596 B.n556 VSUBS 0.007561f
C597 B.n557 VSUBS 0.007561f
C598 B.n558 VSUBS 0.007561f
C599 B.n559 VSUBS 0.007561f
C600 B.n560 VSUBS 0.007561f
C601 B.n561 VSUBS 0.007561f
C602 B.n562 VSUBS 0.007561f
C603 B.n563 VSUBS 0.007561f
C604 B.n564 VSUBS 0.007561f
C605 B.n565 VSUBS 0.007561f
C606 B.n566 VSUBS 0.007561f
C607 B.n567 VSUBS 0.007561f
C608 B.n568 VSUBS 0.007561f
C609 B.n569 VSUBS 0.007561f
C610 B.n570 VSUBS 0.007561f
C611 B.n571 VSUBS 0.007561f
C612 B.n572 VSUBS 0.007561f
C613 B.n573 VSUBS 0.007561f
C614 B.n574 VSUBS 0.007561f
C615 B.n575 VSUBS 0.007561f
C616 B.n576 VSUBS 0.007561f
C617 B.n577 VSUBS 0.007561f
C618 B.n578 VSUBS 0.007561f
C619 B.n579 VSUBS 0.007561f
C620 B.n580 VSUBS 0.007561f
C621 B.n581 VSUBS 0.018735f
C622 B.n582 VSUBS 0.017896f
C623 B.n583 VSUBS 0.019021f
C624 B.n584 VSUBS 0.007561f
C625 B.n585 VSUBS 0.007561f
C626 B.n586 VSUBS 0.007561f
C627 B.n587 VSUBS 0.007561f
C628 B.n588 VSUBS 0.007561f
C629 B.n589 VSUBS 0.007561f
C630 B.n590 VSUBS 0.007561f
C631 B.n591 VSUBS 0.007561f
C632 B.n592 VSUBS 0.007561f
C633 B.n593 VSUBS 0.007561f
C634 B.n594 VSUBS 0.007561f
C635 B.n595 VSUBS 0.007561f
C636 B.n596 VSUBS 0.007561f
C637 B.n597 VSUBS 0.007561f
C638 B.n598 VSUBS 0.007561f
C639 B.n599 VSUBS 0.007561f
C640 B.n600 VSUBS 0.007561f
C641 B.n601 VSUBS 0.007561f
C642 B.n602 VSUBS 0.007561f
C643 B.n603 VSUBS 0.007561f
C644 B.n604 VSUBS 0.007561f
C645 B.n605 VSUBS 0.007561f
C646 B.n606 VSUBS 0.007561f
C647 B.n607 VSUBS 0.007561f
C648 B.n608 VSUBS 0.007561f
C649 B.n609 VSUBS 0.007561f
C650 B.n610 VSUBS 0.007561f
C651 B.n611 VSUBS 0.007561f
C652 B.n612 VSUBS 0.007561f
C653 B.n613 VSUBS 0.007561f
C654 B.n614 VSUBS 0.007561f
C655 B.n615 VSUBS 0.007561f
C656 B.n616 VSUBS 0.007561f
C657 B.n617 VSUBS 0.007561f
C658 B.n618 VSUBS 0.007561f
C659 B.n619 VSUBS 0.007561f
C660 B.n620 VSUBS 0.007561f
C661 B.n621 VSUBS 0.007561f
C662 B.n622 VSUBS 0.007561f
C663 B.n623 VSUBS 0.007561f
C664 B.n624 VSUBS 0.007561f
C665 B.n625 VSUBS 0.007561f
C666 B.n626 VSUBS 0.007561f
C667 B.n627 VSUBS 0.007561f
C668 B.n628 VSUBS 0.007561f
C669 B.n629 VSUBS 0.007561f
C670 B.n630 VSUBS 0.007561f
C671 B.n631 VSUBS 0.007561f
C672 B.n632 VSUBS 0.007561f
C673 B.n633 VSUBS 0.007561f
C674 B.n634 VSUBS 0.007561f
C675 B.n635 VSUBS 0.007561f
C676 B.n636 VSUBS 0.007561f
C677 B.n637 VSUBS 0.007561f
C678 B.n638 VSUBS 0.007561f
C679 B.n639 VSUBS 0.007561f
C680 B.n640 VSUBS 0.007561f
C681 B.n641 VSUBS 0.007561f
C682 B.n642 VSUBS 0.007561f
C683 B.n643 VSUBS 0.007561f
C684 B.n644 VSUBS 0.007561f
C685 B.n645 VSUBS 0.005226f
C686 B.n646 VSUBS 0.017519f
C687 B.n647 VSUBS 0.006116f
C688 B.n648 VSUBS 0.007561f
C689 B.n649 VSUBS 0.007561f
C690 B.n650 VSUBS 0.007561f
C691 B.n651 VSUBS 0.007561f
C692 B.n652 VSUBS 0.007561f
C693 B.n653 VSUBS 0.007561f
C694 B.n654 VSUBS 0.007561f
C695 B.n655 VSUBS 0.007561f
C696 B.n656 VSUBS 0.007561f
C697 B.n657 VSUBS 0.007561f
C698 B.n658 VSUBS 0.007561f
C699 B.n659 VSUBS 0.006116f
C700 B.n660 VSUBS 0.017519f
C701 B.n661 VSUBS 0.005226f
C702 B.n662 VSUBS 0.007561f
C703 B.n663 VSUBS 0.007561f
C704 B.n664 VSUBS 0.007561f
C705 B.n665 VSUBS 0.007561f
C706 B.n666 VSUBS 0.007561f
C707 B.n667 VSUBS 0.007561f
C708 B.n668 VSUBS 0.007561f
C709 B.n669 VSUBS 0.007561f
C710 B.n670 VSUBS 0.007561f
C711 B.n671 VSUBS 0.007561f
C712 B.n672 VSUBS 0.007561f
C713 B.n673 VSUBS 0.007561f
C714 B.n674 VSUBS 0.007561f
C715 B.n675 VSUBS 0.007561f
C716 B.n676 VSUBS 0.007561f
C717 B.n677 VSUBS 0.007561f
C718 B.n678 VSUBS 0.007561f
C719 B.n679 VSUBS 0.007561f
C720 B.n680 VSUBS 0.007561f
C721 B.n681 VSUBS 0.007561f
C722 B.n682 VSUBS 0.007561f
C723 B.n683 VSUBS 0.007561f
C724 B.n684 VSUBS 0.007561f
C725 B.n685 VSUBS 0.007561f
C726 B.n686 VSUBS 0.007561f
C727 B.n687 VSUBS 0.007561f
C728 B.n688 VSUBS 0.007561f
C729 B.n689 VSUBS 0.007561f
C730 B.n690 VSUBS 0.007561f
C731 B.n691 VSUBS 0.007561f
C732 B.n692 VSUBS 0.007561f
C733 B.n693 VSUBS 0.007561f
C734 B.n694 VSUBS 0.007561f
C735 B.n695 VSUBS 0.007561f
C736 B.n696 VSUBS 0.007561f
C737 B.n697 VSUBS 0.007561f
C738 B.n698 VSUBS 0.007561f
C739 B.n699 VSUBS 0.007561f
C740 B.n700 VSUBS 0.007561f
C741 B.n701 VSUBS 0.007561f
C742 B.n702 VSUBS 0.007561f
C743 B.n703 VSUBS 0.007561f
C744 B.n704 VSUBS 0.007561f
C745 B.n705 VSUBS 0.007561f
C746 B.n706 VSUBS 0.007561f
C747 B.n707 VSUBS 0.007561f
C748 B.n708 VSUBS 0.007561f
C749 B.n709 VSUBS 0.007561f
C750 B.n710 VSUBS 0.007561f
C751 B.n711 VSUBS 0.007561f
C752 B.n712 VSUBS 0.007561f
C753 B.n713 VSUBS 0.007561f
C754 B.n714 VSUBS 0.007561f
C755 B.n715 VSUBS 0.007561f
C756 B.n716 VSUBS 0.007561f
C757 B.n717 VSUBS 0.007561f
C758 B.n718 VSUBS 0.007561f
C759 B.n719 VSUBS 0.007561f
C760 B.n720 VSUBS 0.007561f
C761 B.n721 VSUBS 0.007561f
C762 B.n722 VSUBS 0.007561f
C763 B.n723 VSUBS 0.019021f
C764 B.n724 VSUBS 0.017896f
C765 B.n725 VSUBS 0.017896f
C766 B.n726 VSUBS 0.007561f
C767 B.n727 VSUBS 0.007561f
C768 B.n728 VSUBS 0.007561f
C769 B.n729 VSUBS 0.007561f
C770 B.n730 VSUBS 0.007561f
C771 B.n731 VSUBS 0.007561f
C772 B.n732 VSUBS 0.007561f
C773 B.n733 VSUBS 0.007561f
C774 B.n734 VSUBS 0.007561f
C775 B.n735 VSUBS 0.007561f
C776 B.n736 VSUBS 0.007561f
C777 B.n737 VSUBS 0.007561f
C778 B.n738 VSUBS 0.007561f
C779 B.n739 VSUBS 0.007561f
C780 B.n740 VSUBS 0.007561f
C781 B.n741 VSUBS 0.007561f
C782 B.n742 VSUBS 0.007561f
C783 B.n743 VSUBS 0.007561f
C784 B.n744 VSUBS 0.007561f
C785 B.n745 VSUBS 0.007561f
C786 B.n746 VSUBS 0.007561f
C787 B.n747 VSUBS 0.007561f
C788 B.n748 VSUBS 0.007561f
C789 B.n749 VSUBS 0.007561f
C790 B.n750 VSUBS 0.007561f
C791 B.n751 VSUBS 0.007561f
C792 B.n752 VSUBS 0.007561f
C793 B.n753 VSUBS 0.007561f
C794 B.n754 VSUBS 0.007561f
C795 B.n755 VSUBS 0.007561f
C796 B.n756 VSUBS 0.007561f
C797 B.n757 VSUBS 0.007561f
C798 B.n758 VSUBS 0.007561f
C799 B.n759 VSUBS 0.007561f
C800 B.n760 VSUBS 0.007561f
C801 B.n761 VSUBS 0.007561f
C802 B.n762 VSUBS 0.007561f
C803 B.n763 VSUBS 0.007561f
C804 B.n764 VSUBS 0.007561f
C805 B.n765 VSUBS 0.007561f
C806 B.n766 VSUBS 0.007561f
C807 B.n767 VSUBS 0.007561f
C808 B.n768 VSUBS 0.007561f
C809 B.n769 VSUBS 0.007561f
C810 B.n770 VSUBS 0.007561f
C811 B.n771 VSUBS 0.007561f
C812 B.n772 VSUBS 0.007561f
C813 B.n773 VSUBS 0.007561f
C814 B.n774 VSUBS 0.007561f
C815 B.n775 VSUBS 0.007561f
C816 B.n776 VSUBS 0.007561f
C817 B.n777 VSUBS 0.007561f
C818 B.n778 VSUBS 0.007561f
C819 B.n779 VSUBS 0.007561f
C820 B.n780 VSUBS 0.007561f
C821 B.n781 VSUBS 0.007561f
C822 B.n782 VSUBS 0.007561f
C823 B.n783 VSUBS 0.007561f
C824 B.n784 VSUBS 0.007561f
C825 B.n785 VSUBS 0.007561f
C826 B.n786 VSUBS 0.007561f
C827 B.n787 VSUBS 0.007561f
C828 B.n788 VSUBS 0.007561f
C829 B.n789 VSUBS 0.007561f
C830 B.n790 VSUBS 0.007561f
C831 B.n791 VSUBS 0.007561f
C832 B.n792 VSUBS 0.007561f
C833 B.n793 VSUBS 0.007561f
C834 B.n794 VSUBS 0.007561f
C835 B.n795 VSUBS 0.007561f
C836 B.n796 VSUBS 0.007561f
C837 B.n797 VSUBS 0.007561f
C838 B.n798 VSUBS 0.007561f
C839 B.n799 VSUBS 0.007561f
C840 B.n800 VSUBS 0.007561f
C841 B.n801 VSUBS 0.007561f
C842 B.n802 VSUBS 0.007561f
C843 B.n803 VSUBS 0.017121f
C844 VDD2.t2 VSUBS 0.260471f
C845 VDD2.t7 VSUBS 0.260471f
C846 VDD2.n0 VSUBS 2.04055f
C847 VDD2.t4 VSUBS 0.260471f
C848 VDD2.t1 VSUBS 0.260471f
C849 VDD2.n1 VSUBS 2.04055f
C850 VDD2.n2 VSUBS 4.22538f
C851 VDD2.t6 VSUBS 0.260471f
C852 VDD2.t0 VSUBS 0.260471f
C853 VDD2.n3 VSUBS 2.02585f
C854 VDD2.n4 VSUBS 3.55906f
C855 VDD2.t3 VSUBS 0.260471f
C856 VDD2.t5 VSUBS 0.260471f
C857 VDD2.n5 VSUBS 2.0405f
C858 VN.t6 VSUBS 2.51347f
C859 VN.n0 VSUBS 0.999211f
C860 VN.n1 VSUBS 0.028718f
C861 VN.n2 VSUBS 0.057078f
C862 VN.n3 VSUBS 0.028718f
C863 VN.t3 VSUBS 2.51347f
C864 VN.n4 VSUBS 0.057078f
C865 VN.n5 VSUBS 0.028718f
C866 VN.t0 VSUBS 2.51347f
C867 VN.n6 VSUBS 0.989077f
C868 VN.t5 VSUBS 2.75867f
C869 VN.n7 VSUBS 0.949684f
C870 VN.n8 VSUBS 0.297136f
C871 VN.n9 VSUBS 0.053524f
C872 VN.n10 VSUBS 0.057078f
C873 VN.n11 VSUBS 0.023216f
C874 VN.n12 VSUBS 0.028718f
C875 VN.n13 VSUBS 0.028718f
C876 VN.n14 VSUBS 0.028718f
C877 VN.n15 VSUBS 0.053524f
C878 VN.n16 VSUBS 0.915225f
C879 VN.n17 VSUBS 0.053524f
C880 VN.n18 VSUBS 0.028718f
C881 VN.n19 VSUBS 0.028718f
C882 VN.n20 VSUBS 0.028718f
C883 VN.n21 VSUBS 0.023216f
C884 VN.n22 VSUBS 0.057078f
C885 VN.n23 VSUBS 0.053524f
C886 VN.n24 VSUBS 0.046351f
C887 VN.n25 VSUBS 0.050987f
C888 VN.t1 VSUBS 2.51347f
C889 VN.n26 VSUBS 0.999211f
C890 VN.n27 VSUBS 0.028718f
C891 VN.n28 VSUBS 0.057078f
C892 VN.n29 VSUBS 0.028718f
C893 VN.t7 VSUBS 2.51347f
C894 VN.n30 VSUBS 0.057078f
C895 VN.n31 VSUBS 0.028718f
C896 VN.t4 VSUBS 2.51347f
C897 VN.n32 VSUBS 0.989077f
C898 VN.t2 VSUBS 2.75867f
C899 VN.n33 VSUBS 0.949684f
C900 VN.n34 VSUBS 0.297136f
C901 VN.n35 VSUBS 0.053524f
C902 VN.n36 VSUBS 0.057078f
C903 VN.n37 VSUBS 0.023216f
C904 VN.n38 VSUBS 0.028718f
C905 VN.n39 VSUBS 0.028718f
C906 VN.n40 VSUBS 0.028718f
C907 VN.n41 VSUBS 0.053524f
C908 VN.n42 VSUBS 0.915225f
C909 VN.n43 VSUBS 0.053524f
C910 VN.n44 VSUBS 0.028718f
C911 VN.n45 VSUBS 0.028718f
C912 VN.n46 VSUBS 0.028718f
C913 VN.n47 VSUBS 0.023216f
C914 VN.n48 VSUBS 0.057078f
C915 VN.n49 VSUBS 0.053524f
C916 VN.n50 VSUBS 0.046351f
C917 VN.n51 VSUBS 1.68833f
C918 VDD1.t3 VSUBS 0.233324f
C919 VDD1.t1 VSUBS 0.233324f
C920 VDD1.n0 VSUBS 1.82923f
C921 VDD1.t0 VSUBS 0.233324f
C922 VDD1.t4 VSUBS 0.233324f
C923 VDD1.n1 VSUBS 1.82788f
C924 VDD1.t5 VSUBS 0.233324f
C925 VDD1.t2 VSUBS 0.233324f
C926 VDD1.n2 VSUBS 1.82788f
C927 VDD1.n3 VSUBS 3.83608f
C928 VDD1.t6 VSUBS 0.233324f
C929 VDD1.t7 VSUBS 0.233324f
C930 VDD1.n4 VSUBS 1.8147f
C931 VDD1.n5 VSUBS 3.2185f
C932 VTAIL.t1 VSUBS 0.239313f
C933 VTAIL.t5 VSUBS 0.239313f
C934 VTAIL.n0 VSUBS 1.71829f
C935 VTAIL.n1 VSUBS 0.80315f
C936 VTAIL.n2 VSUBS 0.026595f
C937 VTAIL.n3 VSUBS 0.025174f
C938 VTAIL.n4 VSUBS 0.013527f
C939 VTAIL.n5 VSUBS 0.031974f
C940 VTAIL.n6 VSUBS 0.014323f
C941 VTAIL.n7 VSUBS 0.025174f
C942 VTAIL.n8 VSUBS 0.013527f
C943 VTAIL.n9 VSUBS 0.031974f
C944 VTAIL.n10 VSUBS 0.014323f
C945 VTAIL.n11 VSUBS 0.025174f
C946 VTAIL.n12 VSUBS 0.013925f
C947 VTAIL.n13 VSUBS 0.031974f
C948 VTAIL.n14 VSUBS 0.014323f
C949 VTAIL.n15 VSUBS 0.025174f
C950 VTAIL.n16 VSUBS 0.013527f
C951 VTAIL.n17 VSUBS 0.031974f
C952 VTAIL.n18 VSUBS 0.014323f
C953 VTAIL.n19 VSUBS 0.025174f
C954 VTAIL.n20 VSUBS 0.013527f
C955 VTAIL.n21 VSUBS 0.02398f
C956 VTAIL.n22 VSUBS 0.024052f
C957 VTAIL.t0 VSUBS 0.068901f
C958 VTAIL.n23 VSUBS 0.198599f
C959 VTAIL.n24 VSUBS 1.24018f
C960 VTAIL.n25 VSUBS 0.013527f
C961 VTAIL.n26 VSUBS 0.014323f
C962 VTAIL.n27 VSUBS 0.031974f
C963 VTAIL.n28 VSUBS 0.031974f
C964 VTAIL.n29 VSUBS 0.014323f
C965 VTAIL.n30 VSUBS 0.013527f
C966 VTAIL.n31 VSUBS 0.025174f
C967 VTAIL.n32 VSUBS 0.025174f
C968 VTAIL.n33 VSUBS 0.013527f
C969 VTAIL.n34 VSUBS 0.014323f
C970 VTAIL.n35 VSUBS 0.031974f
C971 VTAIL.n36 VSUBS 0.031974f
C972 VTAIL.n37 VSUBS 0.014323f
C973 VTAIL.n38 VSUBS 0.013527f
C974 VTAIL.n39 VSUBS 0.025174f
C975 VTAIL.n40 VSUBS 0.025174f
C976 VTAIL.n41 VSUBS 0.013527f
C977 VTAIL.n42 VSUBS 0.013527f
C978 VTAIL.n43 VSUBS 0.014323f
C979 VTAIL.n44 VSUBS 0.031974f
C980 VTAIL.n45 VSUBS 0.031974f
C981 VTAIL.n46 VSUBS 0.031974f
C982 VTAIL.n47 VSUBS 0.013925f
C983 VTAIL.n48 VSUBS 0.013527f
C984 VTAIL.n49 VSUBS 0.025174f
C985 VTAIL.n50 VSUBS 0.025174f
C986 VTAIL.n51 VSUBS 0.013527f
C987 VTAIL.n52 VSUBS 0.014323f
C988 VTAIL.n53 VSUBS 0.031974f
C989 VTAIL.n54 VSUBS 0.031974f
C990 VTAIL.n55 VSUBS 0.014323f
C991 VTAIL.n56 VSUBS 0.013527f
C992 VTAIL.n57 VSUBS 0.025174f
C993 VTAIL.n58 VSUBS 0.025174f
C994 VTAIL.n59 VSUBS 0.013527f
C995 VTAIL.n60 VSUBS 0.014323f
C996 VTAIL.n61 VSUBS 0.031974f
C997 VTAIL.n62 VSUBS 0.073775f
C998 VTAIL.n63 VSUBS 0.014323f
C999 VTAIL.n64 VSUBS 0.013527f
C1000 VTAIL.n65 VSUBS 0.055093f
C1001 VTAIL.n66 VSUBS 0.036842f
C1002 VTAIL.n67 VSUBS 0.267647f
C1003 VTAIL.n68 VSUBS 0.026595f
C1004 VTAIL.n69 VSUBS 0.025174f
C1005 VTAIL.n70 VSUBS 0.013527f
C1006 VTAIL.n71 VSUBS 0.031974f
C1007 VTAIL.n72 VSUBS 0.014323f
C1008 VTAIL.n73 VSUBS 0.025174f
C1009 VTAIL.n74 VSUBS 0.013527f
C1010 VTAIL.n75 VSUBS 0.031974f
C1011 VTAIL.n76 VSUBS 0.014323f
C1012 VTAIL.n77 VSUBS 0.025174f
C1013 VTAIL.n78 VSUBS 0.013925f
C1014 VTAIL.n79 VSUBS 0.031974f
C1015 VTAIL.n80 VSUBS 0.014323f
C1016 VTAIL.n81 VSUBS 0.025174f
C1017 VTAIL.n82 VSUBS 0.013527f
C1018 VTAIL.n83 VSUBS 0.031974f
C1019 VTAIL.n84 VSUBS 0.014323f
C1020 VTAIL.n85 VSUBS 0.025174f
C1021 VTAIL.n86 VSUBS 0.013527f
C1022 VTAIL.n87 VSUBS 0.02398f
C1023 VTAIL.n88 VSUBS 0.024052f
C1024 VTAIL.t10 VSUBS 0.068901f
C1025 VTAIL.n89 VSUBS 0.198599f
C1026 VTAIL.n90 VSUBS 1.24018f
C1027 VTAIL.n91 VSUBS 0.013527f
C1028 VTAIL.n92 VSUBS 0.014323f
C1029 VTAIL.n93 VSUBS 0.031974f
C1030 VTAIL.n94 VSUBS 0.031974f
C1031 VTAIL.n95 VSUBS 0.014323f
C1032 VTAIL.n96 VSUBS 0.013527f
C1033 VTAIL.n97 VSUBS 0.025174f
C1034 VTAIL.n98 VSUBS 0.025174f
C1035 VTAIL.n99 VSUBS 0.013527f
C1036 VTAIL.n100 VSUBS 0.014323f
C1037 VTAIL.n101 VSUBS 0.031974f
C1038 VTAIL.n102 VSUBS 0.031974f
C1039 VTAIL.n103 VSUBS 0.014323f
C1040 VTAIL.n104 VSUBS 0.013527f
C1041 VTAIL.n105 VSUBS 0.025174f
C1042 VTAIL.n106 VSUBS 0.025174f
C1043 VTAIL.n107 VSUBS 0.013527f
C1044 VTAIL.n108 VSUBS 0.013527f
C1045 VTAIL.n109 VSUBS 0.014323f
C1046 VTAIL.n110 VSUBS 0.031974f
C1047 VTAIL.n111 VSUBS 0.031974f
C1048 VTAIL.n112 VSUBS 0.031974f
C1049 VTAIL.n113 VSUBS 0.013925f
C1050 VTAIL.n114 VSUBS 0.013527f
C1051 VTAIL.n115 VSUBS 0.025174f
C1052 VTAIL.n116 VSUBS 0.025174f
C1053 VTAIL.n117 VSUBS 0.013527f
C1054 VTAIL.n118 VSUBS 0.014323f
C1055 VTAIL.n119 VSUBS 0.031974f
C1056 VTAIL.n120 VSUBS 0.031974f
C1057 VTAIL.n121 VSUBS 0.014323f
C1058 VTAIL.n122 VSUBS 0.013527f
C1059 VTAIL.n123 VSUBS 0.025174f
C1060 VTAIL.n124 VSUBS 0.025174f
C1061 VTAIL.n125 VSUBS 0.013527f
C1062 VTAIL.n126 VSUBS 0.014323f
C1063 VTAIL.n127 VSUBS 0.031974f
C1064 VTAIL.n128 VSUBS 0.073775f
C1065 VTAIL.n129 VSUBS 0.014323f
C1066 VTAIL.n130 VSUBS 0.013527f
C1067 VTAIL.n131 VSUBS 0.055093f
C1068 VTAIL.n132 VSUBS 0.036842f
C1069 VTAIL.n133 VSUBS 0.267647f
C1070 VTAIL.t15 VSUBS 0.239313f
C1071 VTAIL.t9 VSUBS 0.239313f
C1072 VTAIL.n134 VSUBS 1.71829f
C1073 VTAIL.n135 VSUBS 1.00821f
C1074 VTAIL.n136 VSUBS 0.026595f
C1075 VTAIL.n137 VSUBS 0.025174f
C1076 VTAIL.n138 VSUBS 0.013527f
C1077 VTAIL.n139 VSUBS 0.031974f
C1078 VTAIL.n140 VSUBS 0.014323f
C1079 VTAIL.n141 VSUBS 0.025174f
C1080 VTAIL.n142 VSUBS 0.013527f
C1081 VTAIL.n143 VSUBS 0.031974f
C1082 VTAIL.n144 VSUBS 0.014323f
C1083 VTAIL.n145 VSUBS 0.025174f
C1084 VTAIL.n146 VSUBS 0.013925f
C1085 VTAIL.n147 VSUBS 0.031974f
C1086 VTAIL.n148 VSUBS 0.014323f
C1087 VTAIL.n149 VSUBS 0.025174f
C1088 VTAIL.n150 VSUBS 0.013527f
C1089 VTAIL.n151 VSUBS 0.031974f
C1090 VTAIL.n152 VSUBS 0.014323f
C1091 VTAIL.n153 VSUBS 0.025174f
C1092 VTAIL.n154 VSUBS 0.013527f
C1093 VTAIL.n155 VSUBS 0.02398f
C1094 VTAIL.n156 VSUBS 0.024052f
C1095 VTAIL.t12 VSUBS 0.068901f
C1096 VTAIL.n157 VSUBS 0.198599f
C1097 VTAIL.n158 VSUBS 1.24018f
C1098 VTAIL.n159 VSUBS 0.013527f
C1099 VTAIL.n160 VSUBS 0.014323f
C1100 VTAIL.n161 VSUBS 0.031974f
C1101 VTAIL.n162 VSUBS 0.031974f
C1102 VTAIL.n163 VSUBS 0.014323f
C1103 VTAIL.n164 VSUBS 0.013527f
C1104 VTAIL.n165 VSUBS 0.025174f
C1105 VTAIL.n166 VSUBS 0.025174f
C1106 VTAIL.n167 VSUBS 0.013527f
C1107 VTAIL.n168 VSUBS 0.014323f
C1108 VTAIL.n169 VSUBS 0.031974f
C1109 VTAIL.n170 VSUBS 0.031974f
C1110 VTAIL.n171 VSUBS 0.014323f
C1111 VTAIL.n172 VSUBS 0.013527f
C1112 VTAIL.n173 VSUBS 0.025174f
C1113 VTAIL.n174 VSUBS 0.025174f
C1114 VTAIL.n175 VSUBS 0.013527f
C1115 VTAIL.n176 VSUBS 0.013527f
C1116 VTAIL.n177 VSUBS 0.014323f
C1117 VTAIL.n178 VSUBS 0.031974f
C1118 VTAIL.n179 VSUBS 0.031974f
C1119 VTAIL.n180 VSUBS 0.031974f
C1120 VTAIL.n181 VSUBS 0.013925f
C1121 VTAIL.n182 VSUBS 0.013527f
C1122 VTAIL.n183 VSUBS 0.025174f
C1123 VTAIL.n184 VSUBS 0.025174f
C1124 VTAIL.n185 VSUBS 0.013527f
C1125 VTAIL.n186 VSUBS 0.014323f
C1126 VTAIL.n187 VSUBS 0.031974f
C1127 VTAIL.n188 VSUBS 0.031974f
C1128 VTAIL.n189 VSUBS 0.014323f
C1129 VTAIL.n190 VSUBS 0.013527f
C1130 VTAIL.n191 VSUBS 0.025174f
C1131 VTAIL.n192 VSUBS 0.025174f
C1132 VTAIL.n193 VSUBS 0.013527f
C1133 VTAIL.n194 VSUBS 0.014323f
C1134 VTAIL.n195 VSUBS 0.031974f
C1135 VTAIL.n196 VSUBS 0.073775f
C1136 VTAIL.n197 VSUBS 0.014323f
C1137 VTAIL.n198 VSUBS 0.013527f
C1138 VTAIL.n199 VSUBS 0.055093f
C1139 VTAIL.n200 VSUBS 0.036842f
C1140 VTAIL.n201 VSUBS 1.6225f
C1141 VTAIL.n202 VSUBS 0.026595f
C1142 VTAIL.n203 VSUBS 0.025174f
C1143 VTAIL.n204 VSUBS 0.013527f
C1144 VTAIL.n205 VSUBS 0.031974f
C1145 VTAIL.n206 VSUBS 0.014323f
C1146 VTAIL.n207 VSUBS 0.025174f
C1147 VTAIL.n208 VSUBS 0.013527f
C1148 VTAIL.n209 VSUBS 0.031974f
C1149 VTAIL.n210 VSUBS 0.014323f
C1150 VTAIL.n211 VSUBS 0.025174f
C1151 VTAIL.n212 VSUBS 0.013925f
C1152 VTAIL.n213 VSUBS 0.031974f
C1153 VTAIL.n214 VSUBS 0.013527f
C1154 VTAIL.n215 VSUBS 0.014323f
C1155 VTAIL.n216 VSUBS 0.025174f
C1156 VTAIL.n217 VSUBS 0.013527f
C1157 VTAIL.n218 VSUBS 0.031974f
C1158 VTAIL.n219 VSUBS 0.014323f
C1159 VTAIL.n220 VSUBS 0.025174f
C1160 VTAIL.n221 VSUBS 0.013527f
C1161 VTAIL.n222 VSUBS 0.02398f
C1162 VTAIL.n223 VSUBS 0.024052f
C1163 VTAIL.t2 VSUBS 0.068901f
C1164 VTAIL.n224 VSUBS 0.198599f
C1165 VTAIL.n225 VSUBS 1.24018f
C1166 VTAIL.n226 VSUBS 0.013527f
C1167 VTAIL.n227 VSUBS 0.014323f
C1168 VTAIL.n228 VSUBS 0.031974f
C1169 VTAIL.n229 VSUBS 0.031974f
C1170 VTAIL.n230 VSUBS 0.014323f
C1171 VTAIL.n231 VSUBS 0.013527f
C1172 VTAIL.n232 VSUBS 0.025174f
C1173 VTAIL.n233 VSUBS 0.025174f
C1174 VTAIL.n234 VSUBS 0.013527f
C1175 VTAIL.n235 VSUBS 0.014323f
C1176 VTAIL.n236 VSUBS 0.031974f
C1177 VTAIL.n237 VSUBS 0.031974f
C1178 VTAIL.n238 VSUBS 0.014323f
C1179 VTAIL.n239 VSUBS 0.013527f
C1180 VTAIL.n240 VSUBS 0.025174f
C1181 VTAIL.n241 VSUBS 0.025174f
C1182 VTAIL.n242 VSUBS 0.013527f
C1183 VTAIL.n243 VSUBS 0.014323f
C1184 VTAIL.n244 VSUBS 0.031974f
C1185 VTAIL.n245 VSUBS 0.031974f
C1186 VTAIL.n246 VSUBS 0.031974f
C1187 VTAIL.n247 VSUBS 0.013925f
C1188 VTAIL.n248 VSUBS 0.013527f
C1189 VTAIL.n249 VSUBS 0.025174f
C1190 VTAIL.n250 VSUBS 0.025174f
C1191 VTAIL.n251 VSUBS 0.013527f
C1192 VTAIL.n252 VSUBS 0.014323f
C1193 VTAIL.n253 VSUBS 0.031974f
C1194 VTAIL.n254 VSUBS 0.031974f
C1195 VTAIL.n255 VSUBS 0.014323f
C1196 VTAIL.n256 VSUBS 0.013527f
C1197 VTAIL.n257 VSUBS 0.025174f
C1198 VTAIL.n258 VSUBS 0.025174f
C1199 VTAIL.n259 VSUBS 0.013527f
C1200 VTAIL.n260 VSUBS 0.014323f
C1201 VTAIL.n261 VSUBS 0.031974f
C1202 VTAIL.n262 VSUBS 0.073775f
C1203 VTAIL.n263 VSUBS 0.014323f
C1204 VTAIL.n264 VSUBS 0.013527f
C1205 VTAIL.n265 VSUBS 0.055093f
C1206 VTAIL.n266 VSUBS 0.036842f
C1207 VTAIL.n267 VSUBS 1.6225f
C1208 VTAIL.t4 VSUBS 0.239313f
C1209 VTAIL.t7 VSUBS 0.239313f
C1210 VTAIL.n268 VSUBS 1.71831f
C1211 VTAIL.n269 VSUBS 1.0082f
C1212 VTAIL.n270 VSUBS 0.026595f
C1213 VTAIL.n271 VSUBS 0.025174f
C1214 VTAIL.n272 VSUBS 0.013527f
C1215 VTAIL.n273 VSUBS 0.031974f
C1216 VTAIL.n274 VSUBS 0.014323f
C1217 VTAIL.n275 VSUBS 0.025174f
C1218 VTAIL.n276 VSUBS 0.013527f
C1219 VTAIL.n277 VSUBS 0.031974f
C1220 VTAIL.n278 VSUBS 0.014323f
C1221 VTAIL.n279 VSUBS 0.025174f
C1222 VTAIL.n280 VSUBS 0.013925f
C1223 VTAIL.n281 VSUBS 0.031974f
C1224 VTAIL.n282 VSUBS 0.013527f
C1225 VTAIL.n283 VSUBS 0.014323f
C1226 VTAIL.n284 VSUBS 0.025174f
C1227 VTAIL.n285 VSUBS 0.013527f
C1228 VTAIL.n286 VSUBS 0.031974f
C1229 VTAIL.n287 VSUBS 0.014323f
C1230 VTAIL.n288 VSUBS 0.025174f
C1231 VTAIL.n289 VSUBS 0.013527f
C1232 VTAIL.n290 VSUBS 0.02398f
C1233 VTAIL.n291 VSUBS 0.024052f
C1234 VTAIL.t3 VSUBS 0.068901f
C1235 VTAIL.n292 VSUBS 0.198599f
C1236 VTAIL.n293 VSUBS 1.24018f
C1237 VTAIL.n294 VSUBS 0.013527f
C1238 VTAIL.n295 VSUBS 0.014323f
C1239 VTAIL.n296 VSUBS 0.031974f
C1240 VTAIL.n297 VSUBS 0.031974f
C1241 VTAIL.n298 VSUBS 0.014323f
C1242 VTAIL.n299 VSUBS 0.013527f
C1243 VTAIL.n300 VSUBS 0.025174f
C1244 VTAIL.n301 VSUBS 0.025174f
C1245 VTAIL.n302 VSUBS 0.013527f
C1246 VTAIL.n303 VSUBS 0.014323f
C1247 VTAIL.n304 VSUBS 0.031974f
C1248 VTAIL.n305 VSUBS 0.031974f
C1249 VTAIL.n306 VSUBS 0.014323f
C1250 VTAIL.n307 VSUBS 0.013527f
C1251 VTAIL.n308 VSUBS 0.025174f
C1252 VTAIL.n309 VSUBS 0.025174f
C1253 VTAIL.n310 VSUBS 0.013527f
C1254 VTAIL.n311 VSUBS 0.014323f
C1255 VTAIL.n312 VSUBS 0.031974f
C1256 VTAIL.n313 VSUBS 0.031974f
C1257 VTAIL.n314 VSUBS 0.031974f
C1258 VTAIL.n315 VSUBS 0.013925f
C1259 VTAIL.n316 VSUBS 0.013527f
C1260 VTAIL.n317 VSUBS 0.025174f
C1261 VTAIL.n318 VSUBS 0.025174f
C1262 VTAIL.n319 VSUBS 0.013527f
C1263 VTAIL.n320 VSUBS 0.014323f
C1264 VTAIL.n321 VSUBS 0.031974f
C1265 VTAIL.n322 VSUBS 0.031974f
C1266 VTAIL.n323 VSUBS 0.014323f
C1267 VTAIL.n324 VSUBS 0.013527f
C1268 VTAIL.n325 VSUBS 0.025174f
C1269 VTAIL.n326 VSUBS 0.025174f
C1270 VTAIL.n327 VSUBS 0.013527f
C1271 VTAIL.n328 VSUBS 0.014323f
C1272 VTAIL.n329 VSUBS 0.031974f
C1273 VTAIL.n330 VSUBS 0.073775f
C1274 VTAIL.n331 VSUBS 0.014323f
C1275 VTAIL.n332 VSUBS 0.013527f
C1276 VTAIL.n333 VSUBS 0.055093f
C1277 VTAIL.n334 VSUBS 0.036842f
C1278 VTAIL.n335 VSUBS 0.267647f
C1279 VTAIL.n336 VSUBS 0.026595f
C1280 VTAIL.n337 VSUBS 0.025174f
C1281 VTAIL.n338 VSUBS 0.013527f
C1282 VTAIL.n339 VSUBS 0.031974f
C1283 VTAIL.n340 VSUBS 0.014323f
C1284 VTAIL.n341 VSUBS 0.025174f
C1285 VTAIL.n342 VSUBS 0.013527f
C1286 VTAIL.n343 VSUBS 0.031974f
C1287 VTAIL.n344 VSUBS 0.014323f
C1288 VTAIL.n345 VSUBS 0.025174f
C1289 VTAIL.n346 VSUBS 0.013925f
C1290 VTAIL.n347 VSUBS 0.031974f
C1291 VTAIL.n348 VSUBS 0.013527f
C1292 VTAIL.n349 VSUBS 0.014323f
C1293 VTAIL.n350 VSUBS 0.025174f
C1294 VTAIL.n351 VSUBS 0.013527f
C1295 VTAIL.n352 VSUBS 0.031974f
C1296 VTAIL.n353 VSUBS 0.014323f
C1297 VTAIL.n354 VSUBS 0.025174f
C1298 VTAIL.n355 VSUBS 0.013527f
C1299 VTAIL.n356 VSUBS 0.02398f
C1300 VTAIL.n357 VSUBS 0.024052f
C1301 VTAIL.t11 VSUBS 0.068901f
C1302 VTAIL.n358 VSUBS 0.198599f
C1303 VTAIL.n359 VSUBS 1.24018f
C1304 VTAIL.n360 VSUBS 0.013527f
C1305 VTAIL.n361 VSUBS 0.014323f
C1306 VTAIL.n362 VSUBS 0.031974f
C1307 VTAIL.n363 VSUBS 0.031974f
C1308 VTAIL.n364 VSUBS 0.014323f
C1309 VTAIL.n365 VSUBS 0.013527f
C1310 VTAIL.n366 VSUBS 0.025174f
C1311 VTAIL.n367 VSUBS 0.025174f
C1312 VTAIL.n368 VSUBS 0.013527f
C1313 VTAIL.n369 VSUBS 0.014323f
C1314 VTAIL.n370 VSUBS 0.031974f
C1315 VTAIL.n371 VSUBS 0.031974f
C1316 VTAIL.n372 VSUBS 0.014323f
C1317 VTAIL.n373 VSUBS 0.013527f
C1318 VTAIL.n374 VSUBS 0.025174f
C1319 VTAIL.n375 VSUBS 0.025174f
C1320 VTAIL.n376 VSUBS 0.013527f
C1321 VTAIL.n377 VSUBS 0.014323f
C1322 VTAIL.n378 VSUBS 0.031974f
C1323 VTAIL.n379 VSUBS 0.031974f
C1324 VTAIL.n380 VSUBS 0.031974f
C1325 VTAIL.n381 VSUBS 0.013925f
C1326 VTAIL.n382 VSUBS 0.013527f
C1327 VTAIL.n383 VSUBS 0.025174f
C1328 VTAIL.n384 VSUBS 0.025174f
C1329 VTAIL.n385 VSUBS 0.013527f
C1330 VTAIL.n386 VSUBS 0.014323f
C1331 VTAIL.n387 VSUBS 0.031974f
C1332 VTAIL.n388 VSUBS 0.031974f
C1333 VTAIL.n389 VSUBS 0.014323f
C1334 VTAIL.n390 VSUBS 0.013527f
C1335 VTAIL.n391 VSUBS 0.025174f
C1336 VTAIL.n392 VSUBS 0.025174f
C1337 VTAIL.n393 VSUBS 0.013527f
C1338 VTAIL.n394 VSUBS 0.014323f
C1339 VTAIL.n395 VSUBS 0.031974f
C1340 VTAIL.n396 VSUBS 0.073775f
C1341 VTAIL.n397 VSUBS 0.014323f
C1342 VTAIL.n398 VSUBS 0.013527f
C1343 VTAIL.n399 VSUBS 0.055093f
C1344 VTAIL.n400 VSUBS 0.036842f
C1345 VTAIL.n401 VSUBS 0.267647f
C1346 VTAIL.t8 VSUBS 0.239313f
C1347 VTAIL.t14 VSUBS 0.239313f
C1348 VTAIL.n402 VSUBS 1.71831f
C1349 VTAIL.n403 VSUBS 1.0082f
C1350 VTAIL.n404 VSUBS 0.026595f
C1351 VTAIL.n405 VSUBS 0.025174f
C1352 VTAIL.n406 VSUBS 0.013527f
C1353 VTAIL.n407 VSUBS 0.031974f
C1354 VTAIL.n408 VSUBS 0.014323f
C1355 VTAIL.n409 VSUBS 0.025174f
C1356 VTAIL.n410 VSUBS 0.013527f
C1357 VTAIL.n411 VSUBS 0.031974f
C1358 VTAIL.n412 VSUBS 0.014323f
C1359 VTAIL.n413 VSUBS 0.025174f
C1360 VTAIL.n414 VSUBS 0.013925f
C1361 VTAIL.n415 VSUBS 0.031974f
C1362 VTAIL.n416 VSUBS 0.013527f
C1363 VTAIL.n417 VSUBS 0.014323f
C1364 VTAIL.n418 VSUBS 0.025174f
C1365 VTAIL.n419 VSUBS 0.013527f
C1366 VTAIL.n420 VSUBS 0.031974f
C1367 VTAIL.n421 VSUBS 0.014323f
C1368 VTAIL.n422 VSUBS 0.025174f
C1369 VTAIL.n423 VSUBS 0.013527f
C1370 VTAIL.n424 VSUBS 0.02398f
C1371 VTAIL.n425 VSUBS 0.024052f
C1372 VTAIL.t13 VSUBS 0.068901f
C1373 VTAIL.n426 VSUBS 0.198599f
C1374 VTAIL.n427 VSUBS 1.24018f
C1375 VTAIL.n428 VSUBS 0.013527f
C1376 VTAIL.n429 VSUBS 0.014323f
C1377 VTAIL.n430 VSUBS 0.031974f
C1378 VTAIL.n431 VSUBS 0.031974f
C1379 VTAIL.n432 VSUBS 0.014323f
C1380 VTAIL.n433 VSUBS 0.013527f
C1381 VTAIL.n434 VSUBS 0.025174f
C1382 VTAIL.n435 VSUBS 0.025174f
C1383 VTAIL.n436 VSUBS 0.013527f
C1384 VTAIL.n437 VSUBS 0.014323f
C1385 VTAIL.n438 VSUBS 0.031974f
C1386 VTAIL.n439 VSUBS 0.031974f
C1387 VTAIL.n440 VSUBS 0.014323f
C1388 VTAIL.n441 VSUBS 0.013527f
C1389 VTAIL.n442 VSUBS 0.025174f
C1390 VTAIL.n443 VSUBS 0.025174f
C1391 VTAIL.n444 VSUBS 0.013527f
C1392 VTAIL.n445 VSUBS 0.014323f
C1393 VTAIL.n446 VSUBS 0.031974f
C1394 VTAIL.n447 VSUBS 0.031974f
C1395 VTAIL.n448 VSUBS 0.031974f
C1396 VTAIL.n449 VSUBS 0.013925f
C1397 VTAIL.n450 VSUBS 0.013527f
C1398 VTAIL.n451 VSUBS 0.025174f
C1399 VTAIL.n452 VSUBS 0.025174f
C1400 VTAIL.n453 VSUBS 0.013527f
C1401 VTAIL.n454 VSUBS 0.014323f
C1402 VTAIL.n455 VSUBS 0.031974f
C1403 VTAIL.n456 VSUBS 0.031974f
C1404 VTAIL.n457 VSUBS 0.014323f
C1405 VTAIL.n458 VSUBS 0.013527f
C1406 VTAIL.n459 VSUBS 0.025174f
C1407 VTAIL.n460 VSUBS 0.025174f
C1408 VTAIL.n461 VSUBS 0.013527f
C1409 VTAIL.n462 VSUBS 0.014323f
C1410 VTAIL.n463 VSUBS 0.031974f
C1411 VTAIL.n464 VSUBS 0.073775f
C1412 VTAIL.n465 VSUBS 0.014323f
C1413 VTAIL.n466 VSUBS 0.013527f
C1414 VTAIL.n467 VSUBS 0.055093f
C1415 VTAIL.n468 VSUBS 0.036842f
C1416 VTAIL.n469 VSUBS 1.6225f
C1417 VTAIL.n470 VSUBS 0.026595f
C1418 VTAIL.n471 VSUBS 0.025174f
C1419 VTAIL.n472 VSUBS 0.013527f
C1420 VTAIL.n473 VSUBS 0.031974f
C1421 VTAIL.n474 VSUBS 0.014323f
C1422 VTAIL.n475 VSUBS 0.025174f
C1423 VTAIL.n476 VSUBS 0.013527f
C1424 VTAIL.n477 VSUBS 0.031974f
C1425 VTAIL.n478 VSUBS 0.014323f
C1426 VTAIL.n479 VSUBS 0.025174f
C1427 VTAIL.n480 VSUBS 0.013925f
C1428 VTAIL.n481 VSUBS 0.031974f
C1429 VTAIL.n482 VSUBS 0.014323f
C1430 VTAIL.n483 VSUBS 0.025174f
C1431 VTAIL.n484 VSUBS 0.013527f
C1432 VTAIL.n485 VSUBS 0.031974f
C1433 VTAIL.n486 VSUBS 0.014323f
C1434 VTAIL.n487 VSUBS 0.025174f
C1435 VTAIL.n488 VSUBS 0.013527f
C1436 VTAIL.n489 VSUBS 0.02398f
C1437 VTAIL.n490 VSUBS 0.024052f
C1438 VTAIL.t6 VSUBS 0.068901f
C1439 VTAIL.n491 VSUBS 0.198599f
C1440 VTAIL.n492 VSUBS 1.24018f
C1441 VTAIL.n493 VSUBS 0.013527f
C1442 VTAIL.n494 VSUBS 0.014323f
C1443 VTAIL.n495 VSUBS 0.031974f
C1444 VTAIL.n496 VSUBS 0.031974f
C1445 VTAIL.n497 VSUBS 0.014323f
C1446 VTAIL.n498 VSUBS 0.013527f
C1447 VTAIL.n499 VSUBS 0.025174f
C1448 VTAIL.n500 VSUBS 0.025174f
C1449 VTAIL.n501 VSUBS 0.013527f
C1450 VTAIL.n502 VSUBS 0.014323f
C1451 VTAIL.n503 VSUBS 0.031974f
C1452 VTAIL.n504 VSUBS 0.031974f
C1453 VTAIL.n505 VSUBS 0.014323f
C1454 VTAIL.n506 VSUBS 0.013527f
C1455 VTAIL.n507 VSUBS 0.025174f
C1456 VTAIL.n508 VSUBS 0.025174f
C1457 VTAIL.n509 VSUBS 0.013527f
C1458 VTAIL.n510 VSUBS 0.013527f
C1459 VTAIL.n511 VSUBS 0.014323f
C1460 VTAIL.n512 VSUBS 0.031974f
C1461 VTAIL.n513 VSUBS 0.031974f
C1462 VTAIL.n514 VSUBS 0.031974f
C1463 VTAIL.n515 VSUBS 0.013925f
C1464 VTAIL.n516 VSUBS 0.013527f
C1465 VTAIL.n517 VSUBS 0.025174f
C1466 VTAIL.n518 VSUBS 0.025174f
C1467 VTAIL.n519 VSUBS 0.013527f
C1468 VTAIL.n520 VSUBS 0.014323f
C1469 VTAIL.n521 VSUBS 0.031974f
C1470 VTAIL.n522 VSUBS 0.031974f
C1471 VTAIL.n523 VSUBS 0.014323f
C1472 VTAIL.n524 VSUBS 0.013527f
C1473 VTAIL.n525 VSUBS 0.025174f
C1474 VTAIL.n526 VSUBS 0.025174f
C1475 VTAIL.n527 VSUBS 0.013527f
C1476 VTAIL.n528 VSUBS 0.014323f
C1477 VTAIL.n529 VSUBS 0.031974f
C1478 VTAIL.n530 VSUBS 0.073775f
C1479 VTAIL.n531 VSUBS 0.014323f
C1480 VTAIL.n532 VSUBS 0.013527f
C1481 VTAIL.n533 VSUBS 0.055093f
C1482 VTAIL.n534 VSUBS 0.036842f
C1483 VTAIL.n535 VSUBS 1.61778f
C1484 VP.t5 VSUBS 2.73174f
C1485 VP.n0 VSUBS 1.08598f
C1486 VP.n1 VSUBS 0.031212f
C1487 VP.n2 VSUBS 0.062034f
C1488 VP.n3 VSUBS 0.031212f
C1489 VP.t2 VSUBS 2.73174f
C1490 VP.n4 VSUBS 0.062034f
C1491 VP.n5 VSUBS 0.031212f
C1492 VP.t3 VSUBS 2.73174f
C1493 VP.n6 VSUBS 0.994703f
C1494 VP.n7 VSUBS 0.031212f
C1495 VP.n8 VSUBS 0.062034f
C1496 VP.t0 VSUBS 2.73174f
C1497 VP.n9 VSUBS 1.08598f
C1498 VP.n10 VSUBS 0.031212f
C1499 VP.n11 VSUBS 0.062034f
C1500 VP.n12 VSUBS 0.031212f
C1501 VP.t1 VSUBS 2.73174f
C1502 VP.n13 VSUBS 0.062034f
C1503 VP.n14 VSUBS 0.031212f
C1504 VP.t6 VSUBS 2.73174f
C1505 VP.n15 VSUBS 1.07497f
C1506 VP.t4 VSUBS 2.99823f
C1507 VP.n16 VSUBS 1.03216f
C1508 VP.n17 VSUBS 0.32294f
C1509 VP.n18 VSUBS 0.058172f
C1510 VP.n19 VSUBS 0.062034f
C1511 VP.n20 VSUBS 0.025232f
C1512 VP.n21 VSUBS 0.031212f
C1513 VP.n22 VSUBS 0.031212f
C1514 VP.n23 VSUBS 0.031212f
C1515 VP.n24 VSUBS 0.058172f
C1516 VP.n25 VSUBS 0.994703f
C1517 VP.n26 VSUBS 0.058172f
C1518 VP.n27 VSUBS 0.031212f
C1519 VP.n28 VSUBS 0.031212f
C1520 VP.n29 VSUBS 0.031212f
C1521 VP.n30 VSUBS 0.025232f
C1522 VP.n31 VSUBS 0.062034f
C1523 VP.n32 VSUBS 0.058172f
C1524 VP.n33 VSUBS 0.050376f
C1525 VP.n34 VSUBS 1.82228f
C1526 VP.n35 VSUBS 1.84413f
C1527 VP.t7 VSUBS 2.73174f
C1528 VP.n36 VSUBS 1.08598f
C1529 VP.n37 VSUBS 0.058172f
C1530 VP.n38 VSUBS 0.050376f
C1531 VP.n39 VSUBS 0.031212f
C1532 VP.n40 VSUBS 0.031212f
C1533 VP.n41 VSUBS 0.025232f
C1534 VP.n42 VSUBS 0.062034f
C1535 VP.n43 VSUBS 0.058172f
C1536 VP.n44 VSUBS 0.031212f
C1537 VP.n45 VSUBS 0.031212f
C1538 VP.n46 VSUBS 0.031212f
C1539 VP.n47 VSUBS 0.058172f
C1540 VP.n48 VSUBS 0.062034f
C1541 VP.n49 VSUBS 0.025232f
C1542 VP.n50 VSUBS 0.031212f
C1543 VP.n51 VSUBS 0.031212f
C1544 VP.n52 VSUBS 0.031212f
C1545 VP.n53 VSUBS 0.058172f
C1546 VP.n54 VSUBS 0.994703f
C1547 VP.n55 VSUBS 0.058172f
C1548 VP.n56 VSUBS 0.031212f
C1549 VP.n57 VSUBS 0.031212f
C1550 VP.n58 VSUBS 0.031212f
C1551 VP.n59 VSUBS 0.025232f
C1552 VP.n60 VSUBS 0.062034f
C1553 VP.n61 VSUBS 0.058172f
C1554 VP.n62 VSUBS 0.050376f
C1555 VP.n63 VSUBS 0.055414f
.ends

