* NGSPICE file created from diff_pair_sample_1536.ext - technology: sky130A

.subckt diff_pair_sample_1536 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VN.t0 VDD2.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=4.7814 pd=25.3 as=2.0229 ps=12.59 w=12.26 l=0.67
X1 VTAIL.t6 VN.t1 VDD2.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=4.7814 pd=25.3 as=2.0229 ps=12.59 w=12.26 l=0.67
X2 VTAIL.t0 VP.t0 VDD1.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=4.7814 pd=25.3 as=2.0229 ps=12.59 w=12.26 l=0.67
X3 B.t17 B.t15 B.t16 B.t5 sky130_fd_pr__nfet_01v8 ad=4.7814 pd=25.3 as=0 ps=0 w=12.26 l=0.67
X4 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=4.7814 pd=25.3 as=0 ps=0 w=12.26 l=0.67
X5 VDD1.t2 VP.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.0229 pd=12.59 as=4.7814 ps=25.3 w=12.26 l=0.67
X6 VTAIL.t3 VP.t2 VDD1.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=4.7814 pd=25.3 as=2.0229 ps=12.59 w=12.26 l=0.67
X7 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=4.7814 pd=25.3 as=0 ps=0 w=12.26 l=0.67
X8 VDD2.t3 VN.t2 VTAIL.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=2.0229 pd=12.59 as=4.7814 ps=25.3 w=12.26 l=0.67
X9 VDD1.t0 VP.t3 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.0229 pd=12.59 as=4.7814 ps=25.3 w=12.26 l=0.67
X10 VDD2.t2 VN.t3 VTAIL.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=2.0229 pd=12.59 as=4.7814 ps=25.3 w=12.26 l=0.67
X11 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=4.7814 pd=25.3 as=0 ps=0 w=12.26 l=0.67
R0 VN.n0 VN.t1 520.622
R1 VN.n1 VN.t2 520.622
R2 VN.n0 VN.t3 520.572
R3 VN.n1 VN.t0 520.572
R4 VN VN.n1 85.5352
R5 VN VN.n0 44.7132
R6 VDD2.n2 VDD2.n0 100.829
R7 VDD2.n2 VDD2.n1 63.9577
R8 VDD2.n1 VDD2.t1 1.61551
R9 VDD2.n1 VDD2.t3 1.61551
R10 VDD2.n0 VDD2.t0 1.61551
R11 VDD2.n0 VDD2.t2 1.61551
R12 VDD2 VDD2.n2 0.0586897
R13 VTAIL.n5 VTAIL.t0 48.8951
R14 VTAIL.n4 VTAIL.t5 48.8951
R15 VTAIL.n3 VTAIL.t7 48.8951
R16 VTAIL.n7 VTAIL.t4 48.8941
R17 VTAIL.n0 VTAIL.t6 48.8941
R18 VTAIL.n1 VTAIL.t2 48.8941
R19 VTAIL.n2 VTAIL.t3 48.8941
R20 VTAIL.n6 VTAIL.t1 48.8939
R21 VTAIL.n7 VTAIL.n6 23.7979
R22 VTAIL.n3 VTAIL.n2 23.7979
R23 VTAIL.n4 VTAIL.n3 0.862569
R24 VTAIL.n6 VTAIL.n5 0.862569
R25 VTAIL.n2 VTAIL.n1 0.862569
R26 VTAIL VTAIL.n0 0.489724
R27 VTAIL.n5 VTAIL.n4 0.470328
R28 VTAIL.n1 VTAIL.n0 0.470328
R29 VTAIL VTAIL.n7 0.373345
R30 B.n355 B.t15 644.345
R31 B.n353 B.t4 644.345
R32 B.n85 B.t12 644.345
R33 B.n82 B.t8 644.345
R34 B.n619 B.n618 585
R35 B.n272 B.n81 585
R36 B.n271 B.n270 585
R37 B.n269 B.n268 585
R38 B.n267 B.n266 585
R39 B.n265 B.n264 585
R40 B.n263 B.n262 585
R41 B.n261 B.n260 585
R42 B.n259 B.n258 585
R43 B.n257 B.n256 585
R44 B.n255 B.n254 585
R45 B.n253 B.n252 585
R46 B.n251 B.n250 585
R47 B.n249 B.n248 585
R48 B.n247 B.n246 585
R49 B.n245 B.n244 585
R50 B.n243 B.n242 585
R51 B.n241 B.n240 585
R52 B.n239 B.n238 585
R53 B.n237 B.n236 585
R54 B.n235 B.n234 585
R55 B.n233 B.n232 585
R56 B.n231 B.n230 585
R57 B.n229 B.n228 585
R58 B.n227 B.n226 585
R59 B.n225 B.n224 585
R60 B.n223 B.n222 585
R61 B.n221 B.n220 585
R62 B.n219 B.n218 585
R63 B.n217 B.n216 585
R64 B.n215 B.n214 585
R65 B.n213 B.n212 585
R66 B.n211 B.n210 585
R67 B.n209 B.n208 585
R68 B.n207 B.n206 585
R69 B.n205 B.n204 585
R70 B.n203 B.n202 585
R71 B.n201 B.n200 585
R72 B.n199 B.n198 585
R73 B.n197 B.n196 585
R74 B.n195 B.n194 585
R75 B.n193 B.n192 585
R76 B.n191 B.n190 585
R77 B.n189 B.n188 585
R78 B.n187 B.n186 585
R79 B.n185 B.n184 585
R80 B.n183 B.n182 585
R81 B.n181 B.n180 585
R82 B.n179 B.n178 585
R83 B.n177 B.n176 585
R84 B.n175 B.n174 585
R85 B.n173 B.n172 585
R86 B.n171 B.n170 585
R87 B.n169 B.n168 585
R88 B.n167 B.n166 585
R89 B.n165 B.n164 585
R90 B.n163 B.n162 585
R91 B.n161 B.n160 585
R92 B.n159 B.n158 585
R93 B.n157 B.n156 585
R94 B.n155 B.n154 585
R95 B.n153 B.n152 585
R96 B.n151 B.n150 585
R97 B.n149 B.n148 585
R98 B.n147 B.n146 585
R99 B.n145 B.n144 585
R100 B.n143 B.n142 585
R101 B.n141 B.n140 585
R102 B.n139 B.n138 585
R103 B.n137 B.n136 585
R104 B.n135 B.n134 585
R105 B.n133 B.n132 585
R106 B.n131 B.n130 585
R107 B.n129 B.n128 585
R108 B.n127 B.n126 585
R109 B.n125 B.n124 585
R110 B.n123 B.n122 585
R111 B.n121 B.n120 585
R112 B.n119 B.n118 585
R113 B.n117 B.n116 585
R114 B.n115 B.n114 585
R115 B.n113 B.n112 585
R116 B.n111 B.n110 585
R117 B.n109 B.n108 585
R118 B.n107 B.n106 585
R119 B.n105 B.n104 585
R120 B.n103 B.n102 585
R121 B.n101 B.n100 585
R122 B.n99 B.n98 585
R123 B.n97 B.n96 585
R124 B.n95 B.n94 585
R125 B.n93 B.n92 585
R126 B.n91 B.n90 585
R127 B.n89 B.n88 585
R128 B.n617 B.n34 585
R129 B.n622 B.n34 585
R130 B.n616 B.n33 585
R131 B.n623 B.n33 585
R132 B.n615 B.n614 585
R133 B.n614 B.n29 585
R134 B.n613 B.n28 585
R135 B.n629 B.n28 585
R136 B.n612 B.n27 585
R137 B.n630 B.n27 585
R138 B.n611 B.n26 585
R139 B.n631 B.n26 585
R140 B.n610 B.n609 585
R141 B.n609 B.n22 585
R142 B.n608 B.n21 585
R143 B.n637 B.n21 585
R144 B.n607 B.n20 585
R145 B.n638 B.n20 585
R146 B.n606 B.n19 585
R147 B.n639 B.n19 585
R148 B.n605 B.n604 585
R149 B.n604 B.n18 585
R150 B.n603 B.n14 585
R151 B.n645 B.n14 585
R152 B.n602 B.n13 585
R153 B.n646 B.n13 585
R154 B.n601 B.n12 585
R155 B.n647 B.n12 585
R156 B.n600 B.n599 585
R157 B.n599 B.n8 585
R158 B.n598 B.n7 585
R159 B.n653 B.n7 585
R160 B.n597 B.n6 585
R161 B.n654 B.n6 585
R162 B.n596 B.n5 585
R163 B.n655 B.n5 585
R164 B.n595 B.n594 585
R165 B.n594 B.n4 585
R166 B.n593 B.n273 585
R167 B.n593 B.n592 585
R168 B.n583 B.n274 585
R169 B.n275 B.n274 585
R170 B.n585 B.n584 585
R171 B.n586 B.n585 585
R172 B.n582 B.n280 585
R173 B.n280 B.n279 585
R174 B.n581 B.n580 585
R175 B.n580 B.n579 585
R176 B.n282 B.n281 585
R177 B.n572 B.n282 585
R178 B.n571 B.n570 585
R179 B.n573 B.n571 585
R180 B.n569 B.n287 585
R181 B.n287 B.n286 585
R182 B.n568 B.n567 585
R183 B.n567 B.n566 585
R184 B.n289 B.n288 585
R185 B.n290 B.n289 585
R186 B.n559 B.n558 585
R187 B.n560 B.n559 585
R188 B.n557 B.n294 585
R189 B.n298 B.n294 585
R190 B.n556 B.n555 585
R191 B.n555 B.n554 585
R192 B.n296 B.n295 585
R193 B.n297 B.n296 585
R194 B.n547 B.n546 585
R195 B.n548 B.n547 585
R196 B.n545 B.n303 585
R197 B.n303 B.n302 585
R198 B.n540 B.n539 585
R199 B.n538 B.n352 585
R200 B.n537 B.n351 585
R201 B.n542 B.n351 585
R202 B.n536 B.n535 585
R203 B.n534 B.n533 585
R204 B.n532 B.n531 585
R205 B.n530 B.n529 585
R206 B.n528 B.n527 585
R207 B.n526 B.n525 585
R208 B.n524 B.n523 585
R209 B.n522 B.n521 585
R210 B.n520 B.n519 585
R211 B.n518 B.n517 585
R212 B.n516 B.n515 585
R213 B.n514 B.n513 585
R214 B.n512 B.n511 585
R215 B.n510 B.n509 585
R216 B.n508 B.n507 585
R217 B.n506 B.n505 585
R218 B.n504 B.n503 585
R219 B.n502 B.n501 585
R220 B.n500 B.n499 585
R221 B.n498 B.n497 585
R222 B.n496 B.n495 585
R223 B.n494 B.n493 585
R224 B.n492 B.n491 585
R225 B.n490 B.n489 585
R226 B.n488 B.n487 585
R227 B.n486 B.n485 585
R228 B.n484 B.n483 585
R229 B.n482 B.n481 585
R230 B.n480 B.n479 585
R231 B.n478 B.n477 585
R232 B.n476 B.n475 585
R233 B.n474 B.n473 585
R234 B.n472 B.n471 585
R235 B.n470 B.n469 585
R236 B.n468 B.n467 585
R237 B.n466 B.n465 585
R238 B.n464 B.n463 585
R239 B.n462 B.n461 585
R240 B.n460 B.n459 585
R241 B.n457 B.n456 585
R242 B.n455 B.n454 585
R243 B.n453 B.n452 585
R244 B.n451 B.n450 585
R245 B.n449 B.n448 585
R246 B.n447 B.n446 585
R247 B.n445 B.n444 585
R248 B.n443 B.n442 585
R249 B.n441 B.n440 585
R250 B.n439 B.n438 585
R251 B.n436 B.n435 585
R252 B.n434 B.n433 585
R253 B.n432 B.n431 585
R254 B.n430 B.n429 585
R255 B.n428 B.n427 585
R256 B.n426 B.n425 585
R257 B.n424 B.n423 585
R258 B.n422 B.n421 585
R259 B.n420 B.n419 585
R260 B.n418 B.n417 585
R261 B.n416 B.n415 585
R262 B.n414 B.n413 585
R263 B.n412 B.n411 585
R264 B.n410 B.n409 585
R265 B.n408 B.n407 585
R266 B.n406 B.n405 585
R267 B.n404 B.n403 585
R268 B.n402 B.n401 585
R269 B.n400 B.n399 585
R270 B.n398 B.n397 585
R271 B.n396 B.n395 585
R272 B.n394 B.n393 585
R273 B.n392 B.n391 585
R274 B.n390 B.n389 585
R275 B.n388 B.n387 585
R276 B.n386 B.n385 585
R277 B.n384 B.n383 585
R278 B.n382 B.n381 585
R279 B.n380 B.n379 585
R280 B.n378 B.n377 585
R281 B.n376 B.n375 585
R282 B.n374 B.n373 585
R283 B.n372 B.n371 585
R284 B.n370 B.n369 585
R285 B.n368 B.n367 585
R286 B.n366 B.n365 585
R287 B.n364 B.n363 585
R288 B.n362 B.n361 585
R289 B.n360 B.n359 585
R290 B.n358 B.n357 585
R291 B.n305 B.n304 585
R292 B.n544 B.n543 585
R293 B.n543 B.n542 585
R294 B.n301 B.n300 585
R295 B.n302 B.n301 585
R296 B.n550 B.n549 585
R297 B.n549 B.n548 585
R298 B.n551 B.n299 585
R299 B.n299 B.n297 585
R300 B.n553 B.n552 585
R301 B.n554 B.n553 585
R302 B.n293 B.n292 585
R303 B.n298 B.n293 585
R304 B.n562 B.n561 585
R305 B.n561 B.n560 585
R306 B.n563 B.n291 585
R307 B.n291 B.n290 585
R308 B.n565 B.n564 585
R309 B.n566 B.n565 585
R310 B.n285 B.n284 585
R311 B.n286 B.n285 585
R312 B.n575 B.n574 585
R313 B.n574 B.n573 585
R314 B.n576 B.n283 585
R315 B.n572 B.n283 585
R316 B.n578 B.n577 585
R317 B.n579 B.n578 585
R318 B.n278 B.n277 585
R319 B.n279 B.n278 585
R320 B.n588 B.n587 585
R321 B.n587 B.n586 585
R322 B.n589 B.n276 585
R323 B.n276 B.n275 585
R324 B.n591 B.n590 585
R325 B.n592 B.n591 585
R326 B.n2 B.n0 585
R327 B.n4 B.n2 585
R328 B.n3 B.n1 585
R329 B.n654 B.n3 585
R330 B.n652 B.n651 585
R331 B.n653 B.n652 585
R332 B.n650 B.n9 585
R333 B.n9 B.n8 585
R334 B.n649 B.n648 585
R335 B.n648 B.n647 585
R336 B.n11 B.n10 585
R337 B.n646 B.n11 585
R338 B.n644 B.n643 585
R339 B.n645 B.n644 585
R340 B.n642 B.n15 585
R341 B.n18 B.n15 585
R342 B.n641 B.n640 585
R343 B.n640 B.n639 585
R344 B.n17 B.n16 585
R345 B.n638 B.n17 585
R346 B.n636 B.n635 585
R347 B.n637 B.n636 585
R348 B.n634 B.n23 585
R349 B.n23 B.n22 585
R350 B.n633 B.n632 585
R351 B.n632 B.n631 585
R352 B.n25 B.n24 585
R353 B.n630 B.n25 585
R354 B.n628 B.n627 585
R355 B.n629 B.n628 585
R356 B.n626 B.n30 585
R357 B.n30 B.n29 585
R358 B.n625 B.n624 585
R359 B.n624 B.n623 585
R360 B.n32 B.n31 585
R361 B.n622 B.n32 585
R362 B.n657 B.n656 585
R363 B.n656 B.n655 585
R364 B.n540 B.n301 516.524
R365 B.n88 B.n32 516.524
R366 B.n543 B.n303 516.524
R367 B.n619 B.n34 516.524
R368 B.n621 B.n620 256.663
R369 B.n621 B.n80 256.663
R370 B.n621 B.n79 256.663
R371 B.n621 B.n78 256.663
R372 B.n621 B.n77 256.663
R373 B.n621 B.n76 256.663
R374 B.n621 B.n75 256.663
R375 B.n621 B.n74 256.663
R376 B.n621 B.n73 256.663
R377 B.n621 B.n72 256.663
R378 B.n621 B.n71 256.663
R379 B.n621 B.n70 256.663
R380 B.n621 B.n69 256.663
R381 B.n621 B.n68 256.663
R382 B.n621 B.n67 256.663
R383 B.n621 B.n66 256.663
R384 B.n621 B.n65 256.663
R385 B.n621 B.n64 256.663
R386 B.n621 B.n63 256.663
R387 B.n621 B.n62 256.663
R388 B.n621 B.n61 256.663
R389 B.n621 B.n60 256.663
R390 B.n621 B.n59 256.663
R391 B.n621 B.n58 256.663
R392 B.n621 B.n57 256.663
R393 B.n621 B.n56 256.663
R394 B.n621 B.n55 256.663
R395 B.n621 B.n54 256.663
R396 B.n621 B.n53 256.663
R397 B.n621 B.n52 256.663
R398 B.n621 B.n51 256.663
R399 B.n621 B.n50 256.663
R400 B.n621 B.n49 256.663
R401 B.n621 B.n48 256.663
R402 B.n621 B.n47 256.663
R403 B.n621 B.n46 256.663
R404 B.n621 B.n45 256.663
R405 B.n621 B.n44 256.663
R406 B.n621 B.n43 256.663
R407 B.n621 B.n42 256.663
R408 B.n621 B.n41 256.663
R409 B.n621 B.n40 256.663
R410 B.n621 B.n39 256.663
R411 B.n621 B.n38 256.663
R412 B.n621 B.n37 256.663
R413 B.n621 B.n36 256.663
R414 B.n621 B.n35 256.663
R415 B.n542 B.n541 256.663
R416 B.n542 B.n306 256.663
R417 B.n542 B.n307 256.663
R418 B.n542 B.n308 256.663
R419 B.n542 B.n309 256.663
R420 B.n542 B.n310 256.663
R421 B.n542 B.n311 256.663
R422 B.n542 B.n312 256.663
R423 B.n542 B.n313 256.663
R424 B.n542 B.n314 256.663
R425 B.n542 B.n315 256.663
R426 B.n542 B.n316 256.663
R427 B.n542 B.n317 256.663
R428 B.n542 B.n318 256.663
R429 B.n542 B.n319 256.663
R430 B.n542 B.n320 256.663
R431 B.n542 B.n321 256.663
R432 B.n542 B.n322 256.663
R433 B.n542 B.n323 256.663
R434 B.n542 B.n324 256.663
R435 B.n542 B.n325 256.663
R436 B.n542 B.n326 256.663
R437 B.n542 B.n327 256.663
R438 B.n542 B.n328 256.663
R439 B.n542 B.n329 256.663
R440 B.n542 B.n330 256.663
R441 B.n542 B.n331 256.663
R442 B.n542 B.n332 256.663
R443 B.n542 B.n333 256.663
R444 B.n542 B.n334 256.663
R445 B.n542 B.n335 256.663
R446 B.n542 B.n336 256.663
R447 B.n542 B.n337 256.663
R448 B.n542 B.n338 256.663
R449 B.n542 B.n339 256.663
R450 B.n542 B.n340 256.663
R451 B.n542 B.n341 256.663
R452 B.n542 B.n342 256.663
R453 B.n542 B.n343 256.663
R454 B.n542 B.n344 256.663
R455 B.n542 B.n345 256.663
R456 B.n542 B.n346 256.663
R457 B.n542 B.n347 256.663
R458 B.n542 B.n348 256.663
R459 B.n542 B.n349 256.663
R460 B.n542 B.n350 256.663
R461 B.n549 B.n301 163.367
R462 B.n549 B.n299 163.367
R463 B.n553 B.n299 163.367
R464 B.n553 B.n293 163.367
R465 B.n561 B.n293 163.367
R466 B.n561 B.n291 163.367
R467 B.n565 B.n291 163.367
R468 B.n565 B.n285 163.367
R469 B.n574 B.n285 163.367
R470 B.n574 B.n283 163.367
R471 B.n578 B.n283 163.367
R472 B.n578 B.n278 163.367
R473 B.n587 B.n278 163.367
R474 B.n587 B.n276 163.367
R475 B.n591 B.n276 163.367
R476 B.n591 B.n2 163.367
R477 B.n656 B.n2 163.367
R478 B.n656 B.n3 163.367
R479 B.n652 B.n3 163.367
R480 B.n652 B.n9 163.367
R481 B.n648 B.n9 163.367
R482 B.n648 B.n11 163.367
R483 B.n644 B.n11 163.367
R484 B.n644 B.n15 163.367
R485 B.n640 B.n15 163.367
R486 B.n640 B.n17 163.367
R487 B.n636 B.n17 163.367
R488 B.n636 B.n23 163.367
R489 B.n632 B.n23 163.367
R490 B.n632 B.n25 163.367
R491 B.n628 B.n25 163.367
R492 B.n628 B.n30 163.367
R493 B.n624 B.n30 163.367
R494 B.n624 B.n32 163.367
R495 B.n352 B.n351 163.367
R496 B.n535 B.n351 163.367
R497 B.n533 B.n532 163.367
R498 B.n529 B.n528 163.367
R499 B.n525 B.n524 163.367
R500 B.n521 B.n520 163.367
R501 B.n517 B.n516 163.367
R502 B.n513 B.n512 163.367
R503 B.n509 B.n508 163.367
R504 B.n505 B.n504 163.367
R505 B.n501 B.n500 163.367
R506 B.n497 B.n496 163.367
R507 B.n493 B.n492 163.367
R508 B.n489 B.n488 163.367
R509 B.n485 B.n484 163.367
R510 B.n481 B.n480 163.367
R511 B.n477 B.n476 163.367
R512 B.n473 B.n472 163.367
R513 B.n469 B.n468 163.367
R514 B.n465 B.n464 163.367
R515 B.n461 B.n460 163.367
R516 B.n456 B.n455 163.367
R517 B.n452 B.n451 163.367
R518 B.n448 B.n447 163.367
R519 B.n444 B.n443 163.367
R520 B.n440 B.n439 163.367
R521 B.n435 B.n434 163.367
R522 B.n431 B.n430 163.367
R523 B.n427 B.n426 163.367
R524 B.n423 B.n422 163.367
R525 B.n419 B.n418 163.367
R526 B.n415 B.n414 163.367
R527 B.n411 B.n410 163.367
R528 B.n407 B.n406 163.367
R529 B.n403 B.n402 163.367
R530 B.n399 B.n398 163.367
R531 B.n395 B.n394 163.367
R532 B.n391 B.n390 163.367
R533 B.n387 B.n386 163.367
R534 B.n383 B.n382 163.367
R535 B.n379 B.n378 163.367
R536 B.n375 B.n374 163.367
R537 B.n371 B.n370 163.367
R538 B.n367 B.n366 163.367
R539 B.n363 B.n362 163.367
R540 B.n359 B.n358 163.367
R541 B.n543 B.n305 163.367
R542 B.n547 B.n303 163.367
R543 B.n547 B.n296 163.367
R544 B.n555 B.n296 163.367
R545 B.n555 B.n294 163.367
R546 B.n559 B.n294 163.367
R547 B.n559 B.n289 163.367
R548 B.n567 B.n289 163.367
R549 B.n567 B.n287 163.367
R550 B.n571 B.n287 163.367
R551 B.n571 B.n282 163.367
R552 B.n580 B.n282 163.367
R553 B.n580 B.n280 163.367
R554 B.n585 B.n280 163.367
R555 B.n585 B.n274 163.367
R556 B.n593 B.n274 163.367
R557 B.n594 B.n593 163.367
R558 B.n594 B.n5 163.367
R559 B.n6 B.n5 163.367
R560 B.n7 B.n6 163.367
R561 B.n599 B.n7 163.367
R562 B.n599 B.n12 163.367
R563 B.n13 B.n12 163.367
R564 B.n14 B.n13 163.367
R565 B.n604 B.n14 163.367
R566 B.n604 B.n19 163.367
R567 B.n20 B.n19 163.367
R568 B.n21 B.n20 163.367
R569 B.n609 B.n21 163.367
R570 B.n609 B.n26 163.367
R571 B.n27 B.n26 163.367
R572 B.n28 B.n27 163.367
R573 B.n614 B.n28 163.367
R574 B.n614 B.n33 163.367
R575 B.n34 B.n33 163.367
R576 B.n92 B.n91 163.367
R577 B.n96 B.n95 163.367
R578 B.n100 B.n99 163.367
R579 B.n104 B.n103 163.367
R580 B.n108 B.n107 163.367
R581 B.n112 B.n111 163.367
R582 B.n116 B.n115 163.367
R583 B.n120 B.n119 163.367
R584 B.n124 B.n123 163.367
R585 B.n128 B.n127 163.367
R586 B.n132 B.n131 163.367
R587 B.n136 B.n135 163.367
R588 B.n140 B.n139 163.367
R589 B.n144 B.n143 163.367
R590 B.n148 B.n147 163.367
R591 B.n152 B.n151 163.367
R592 B.n156 B.n155 163.367
R593 B.n160 B.n159 163.367
R594 B.n164 B.n163 163.367
R595 B.n168 B.n167 163.367
R596 B.n172 B.n171 163.367
R597 B.n176 B.n175 163.367
R598 B.n180 B.n179 163.367
R599 B.n184 B.n183 163.367
R600 B.n188 B.n187 163.367
R601 B.n192 B.n191 163.367
R602 B.n196 B.n195 163.367
R603 B.n200 B.n199 163.367
R604 B.n204 B.n203 163.367
R605 B.n208 B.n207 163.367
R606 B.n212 B.n211 163.367
R607 B.n216 B.n215 163.367
R608 B.n220 B.n219 163.367
R609 B.n224 B.n223 163.367
R610 B.n228 B.n227 163.367
R611 B.n232 B.n231 163.367
R612 B.n236 B.n235 163.367
R613 B.n240 B.n239 163.367
R614 B.n244 B.n243 163.367
R615 B.n248 B.n247 163.367
R616 B.n252 B.n251 163.367
R617 B.n256 B.n255 163.367
R618 B.n260 B.n259 163.367
R619 B.n264 B.n263 163.367
R620 B.n268 B.n267 163.367
R621 B.n270 B.n81 163.367
R622 B.n355 B.t17 87.5372
R623 B.n82 B.t10 87.5372
R624 B.n353 B.t7 87.5215
R625 B.n85 B.t13 87.5215
R626 B.n542 B.n302 74.6512
R627 B.n622 B.n621 74.6512
R628 B.n541 B.n540 71.676
R629 B.n535 B.n306 71.676
R630 B.n532 B.n307 71.676
R631 B.n528 B.n308 71.676
R632 B.n524 B.n309 71.676
R633 B.n520 B.n310 71.676
R634 B.n516 B.n311 71.676
R635 B.n512 B.n312 71.676
R636 B.n508 B.n313 71.676
R637 B.n504 B.n314 71.676
R638 B.n500 B.n315 71.676
R639 B.n496 B.n316 71.676
R640 B.n492 B.n317 71.676
R641 B.n488 B.n318 71.676
R642 B.n484 B.n319 71.676
R643 B.n480 B.n320 71.676
R644 B.n476 B.n321 71.676
R645 B.n472 B.n322 71.676
R646 B.n468 B.n323 71.676
R647 B.n464 B.n324 71.676
R648 B.n460 B.n325 71.676
R649 B.n455 B.n326 71.676
R650 B.n451 B.n327 71.676
R651 B.n447 B.n328 71.676
R652 B.n443 B.n329 71.676
R653 B.n439 B.n330 71.676
R654 B.n434 B.n331 71.676
R655 B.n430 B.n332 71.676
R656 B.n426 B.n333 71.676
R657 B.n422 B.n334 71.676
R658 B.n418 B.n335 71.676
R659 B.n414 B.n336 71.676
R660 B.n410 B.n337 71.676
R661 B.n406 B.n338 71.676
R662 B.n402 B.n339 71.676
R663 B.n398 B.n340 71.676
R664 B.n394 B.n341 71.676
R665 B.n390 B.n342 71.676
R666 B.n386 B.n343 71.676
R667 B.n382 B.n344 71.676
R668 B.n378 B.n345 71.676
R669 B.n374 B.n346 71.676
R670 B.n370 B.n347 71.676
R671 B.n366 B.n348 71.676
R672 B.n362 B.n349 71.676
R673 B.n358 B.n350 71.676
R674 B.n88 B.n35 71.676
R675 B.n92 B.n36 71.676
R676 B.n96 B.n37 71.676
R677 B.n100 B.n38 71.676
R678 B.n104 B.n39 71.676
R679 B.n108 B.n40 71.676
R680 B.n112 B.n41 71.676
R681 B.n116 B.n42 71.676
R682 B.n120 B.n43 71.676
R683 B.n124 B.n44 71.676
R684 B.n128 B.n45 71.676
R685 B.n132 B.n46 71.676
R686 B.n136 B.n47 71.676
R687 B.n140 B.n48 71.676
R688 B.n144 B.n49 71.676
R689 B.n148 B.n50 71.676
R690 B.n152 B.n51 71.676
R691 B.n156 B.n52 71.676
R692 B.n160 B.n53 71.676
R693 B.n164 B.n54 71.676
R694 B.n168 B.n55 71.676
R695 B.n172 B.n56 71.676
R696 B.n176 B.n57 71.676
R697 B.n180 B.n58 71.676
R698 B.n184 B.n59 71.676
R699 B.n188 B.n60 71.676
R700 B.n192 B.n61 71.676
R701 B.n196 B.n62 71.676
R702 B.n200 B.n63 71.676
R703 B.n204 B.n64 71.676
R704 B.n208 B.n65 71.676
R705 B.n212 B.n66 71.676
R706 B.n216 B.n67 71.676
R707 B.n220 B.n68 71.676
R708 B.n224 B.n69 71.676
R709 B.n228 B.n70 71.676
R710 B.n232 B.n71 71.676
R711 B.n236 B.n72 71.676
R712 B.n240 B.n73 71.676
R713 B.n244 B.n74 71.676
R714 B.n248 B.n75 71.676
R715 B.n252 B.n76 71.676
R716 B.n256 B.n77 71.676
R717 B.n260 B.n78 71.676
R718 B.n264 B.n79 71.676
R719 B.n268 B.n80 71.676
R720 B.n620 B.n81 71.676
R721 B.n620 B.n619 71.676
R722 B.n270 B.n80 71.676
R723 B.n267 B.n79 71.676
R724 B.n263 B.n78 71.676
R725 B.n259 B.n77 71.676
R726 B.n255 B.n76 71.676
R727 B.n251 B.n75 71.676
R728 B.n247 B.n74 71.676
R729 B.n243 B.n73 71.676
R730 B.n239 B.n72 71.676
R731 B.n235 B.n71 71.676
R732 B.n231 B.n70 71.676
R733 B.n227 B.n69 71.676
R734 B.n223 B.n68 71.676
R735 B.n219 B.n67 71.676
R736 B.n215 B.n66 71.676
R737 B.n211 B.n65 71.676
R738 B.n207 B.n64 71.676
R739 B.n203 B.n63 71.676
R740 B.n199 B.n62 71.676
R741 B.n195 B.n61 71.676
R742 B.n191 B.n60 71.676
R743 B.n187 B.n59 71.676
R744 B.n183 B.n58 71.676
R745 B.n179 B.n57 71.676
R746 B.n175 B.n56 71.676
R747 B.n171 B.n55 71.676
R748 B.n167 B.n54 71.676
R749 B.n163 B.n53 71.676
R750 B.n159 B.n52 71.676
R751 B.n155 B.n51 71.676
R752 B.n151 B.n50 71.676
R753 B.n147 B.n49 71.676
R754 B.n143 B.n48 71.676
R755 B.n139 B.n47 71.676
R756 B.n135 B.n46 71.676
R757 B.n131 B.n45 71.676
R758 B.n127 B.n44 71.676
R759 B.n123 B.n43 71.676
R760 B.n119 B.n42 71.676
R761 B.n115 B.n41 71.676
R762 B.n111 B.n40 71.676
R763 B.n107 B.n39 71.676
R764 B.n103 B.n38 71.676
R765 B.n99 B.n37 71.676
R766 B.n95 B.n36 71.676
R767 B.n91 B.n35 71.676
R768 B.n541 B.n352 71.676
R769 B.n533 B.n306 71.676
R770 B.n529 B.n307 71.676
R771 B.n525 B.n308 71.676
R772 B.n521 B.n309 71.676
R773 B.n517 B.n310 71.676
R774 B.n513 B.n311 71.676
R775 B.n509 B.n312 71.676
R776 B.n505 B.n313 71.676
R777 B.n501 B.n314 71.676
R778 B.n497 B.n315 71.676
R779 B.n493 B.n316 71.676
R780 B.n489 B.n317 71.676
R781 B.n485 B.n318 71.676
R782 B.n481 B.n319 71.676
R783 B.n477 B.n320 71.676
R784 B.n473 B.n321 71.676
R785 B.n469 B.n322 71.676
R786 B.n465 B.n323 71.676
R787 B.n461 B.n324 71.676
R788 B.n456 B.n325 71.676
R789 B.n452 B.n326 71.676
R790 B.n448 B.n327 71.676
R791 B.n444 B.n328 71.676
R792 B.n440 B.n329 71.676
R793 B.n435 B.n330 71.676
R794 B.n431 B.n331 71.676
R795 B.n427 B.n332 71.676
R796 B.n423 B.n333 71.676
R797 B.n419 B.n334 71.676
R798 B.n415 B.n335 71.676
R799 B.n411 B.n336 71.676
R800 B.n407 B.n337 71.676
R801 B.n403 B.n338 71.676
R802 B.n399 B.n339 71.676
R803 B.n395 B.n340 71.676
R804 B.n391 B.n341 71.676
R805 B.n387 B.n342 71.676
R806 B.n383 B.n343 71.676
R807 B.n379 B.n344 71.676
R808 B.n375 B.n345 71.676
R809 B.n371 B.n346 71.676
R810 B.n367 B.n347 71.676
R811 B.n363 B.n348 71.676
R812 B.n359 B.n349 71.676
R813 B.n350 B.n305 71.676
R814 B.n356 B.t16 68.1433
R815 B.n83 B.t11 68.1433
R816 B.n354 B.t6 68.1275
R817 B.n86 B.t14 68.1275
R818 B.n437 B.n356 59.5399
R819 B.n458 B.n354 59.5399
R820 B.n87 B.n86 59.5399
R821 B.n84 B.n83 59.5399
R822 B.n548 B.n302 42.658
R823 B.n548 B.n297 42.658
R824 B.n554 B.n297 42.658
R825 B.n554 B.n298 42.658
R826 B.n560 B.n290 42.658
R827 B.n566 B.n290 42.658
R828 B.n566 B.n286 42.658
R829 B.n573 B.n286 42.658
R830 B.n573 B.n572 42.658
R831 B.n579 B.n279 42.658
R832 B.n586 B.n279 42.658
R833 B.n592 B.n275 42.658
R834 B.n592 B.n4 42.658
R835 B.n655 B.n4 42.658
R836 B.n655 B.n654 42.658
R837 B.n654 B.n653 42.658
R838 B.n653 B.n8 42.658
R839 B.n647 B.n646 42.658
R840 B.n646 B.n645 42.658
R841 B.n639 B.n18 42.658
R842 B.n639 B.n638 42.658
R843 B.n638 B.n637 42.658
R844 B.n637 B.n22 42.658
R845 B.n631 B.n22 42.658
R846 B.n630 B.n629 42.658
R847 B.n629 B.n29 42.658
R848 B.n623 B.n29 42.658
R849 B.n623 B.n622 42.658
R850 B.n572 B.t3 42.0307
R851 B.n18 B.t1 42.0307
R852 B.n586 B.t2 39.5215
R853 B.n647 B.t0 39.5215
R854 B.n298 B.t5 35.7576
R855 B.t9 B.n630 35.7576
R856 B.n89 B.n31 33.5615
R857 B.n618 B.n617 33.5615
R858 B.n545 B.n544 33.5615
R859 B.n539 B.n300 33.5615
R860 B.n356 B.n355 19.3944
R861 B.n354 B.n353 19.3944
R862 B.n86 B.n85 19.3944
R863 B.n83 B.n82 19.3944
R864 B B.n657 18.0485
R865 B.n90 B.n89 10.6151
R866 B.n93 B.n90 10.6151
R867 B.n94 B.n93 10.6151
R868 B.n97 B.n94 10.6151
R869 B.n98 B.n97 10.6151
R870 B.n101 B.n98 10.6151
R871 B.n102 B.n101 10.6151
R872 B.n105 B.n102 10.6151
R873 B.n106 B.n105 10.6151
R874 B.n109 B.n106 10.6151
R875 B.n110 B.n109 10.6151
R876 B.n113 B.n110 10.6151
R877 B.n114 B.n113 10.6151
R878 B.n117 B.n114 10.6151
R879 B.n118 B.n117 10.6151
R880 B.n121 B.n118 10.6151
R881 B.n122 B.n121 10.6151
R882 B.n125 B.n122 10.6151
R883 B.n126 B.n125 10.6151
R884 B.n129 B.n126 10.6151
R885 B.n130 B.n129 10.6151
R886 B.n133 B.n130 10.6151
R887 B.n134 B.n133 10.6151
R888 B.n137 B.n134 10.6151
R889 B.n138 B.n137 10.6151
R890 B.n141 B.n138 10.6151
R891 B.n142 B.n141 10.6151
R892 B.n145 B.n142 10.6151
R893 B.n146 B.n145 10.6151
R894 B.n149 B.n146 10.6151
R895 B.n150 B.n149 10.6151
R896 B.n153 B.n150 10.6151
R897 B.n154 B.n153 10.6151
R898 B.n157 B.n154 10.6151
R899 B.n158 B.n157 10.6151
R900 B.n161 B.n158 10.6151
R901 B.n162 B.n161 10.6151
R902 B.n165 B.n162 10.6151
R903 B.n166 B.n165 10.6151
R904 B.n169 B.n166 10.6151
R905 B.n170 B.n169 10.6151
R906 B.n174 B.n173 10.6151
R907 B.n177 B.n174 10.6151
R908 B.n178 B.n177 10.6151
R909 B.n181 B.n178 10.6151
R910 B.n182 B.n181 10.6151
R911 B.n185 B.n182 10.6151
R912 B.n186 B.n185 10.6151
R913 B.n189 B.n186 10.6151
R914 B.n190 B.n189 10.6151
R915 B.n194 B.n193 10.6151
R916 B.n197 B.n194 10.6151
R917 B.n198 B.n197 10.6151
R918 B.n201 B.n198 10.6151
R919 B.n202 B.n201 10.6151
R920 B.n205 B.n202 10.6151
R921 B.n206 B.n205 10.6151
R922 B.n209 B.n206 10.6151
R923 B.n210 B.n209 10.6151
R924 B.n213 B.n210 10.6151
R925 B.n214 B.n213 10.6151
R926 B.n217 B.n214 10.6151
R927 B.n218 B.n217 10.6151
R928 B.n221 B.n218 10.6151
R929 B.n222 B.n221 10.6151
R930 B.n225 B.n222 10.6151
R931 B.n226 B.n225 10.6151
R932 B.n229 B.n226 10.6151
R933 B.n230 B.n229 10.6151
R934 B.n233 B.n230 10.6151
R935 B.n234 B.n233 10.6151
R936 B.n237 B.n234 10.6151
R937 B.n238 B.n237 10.6151
R938 B.n241 B.n238 10.6151
R939 B.n242 B.n241 10.6151
R940 B.n245 B.n242 10.6151
R941 B.n246 B.n245 10.6151
R942 B.n249 B.n246 10.6151
R943 B.n250 B.n249 10.6151
R944 B.n253 B.n250 10.6151
R945 B.n254 B.n253 10.6151
R946 B.n257 B.n254 10.6151
R947 B.n258 B.n257 10.6151
R948 B.n261 B.n258 10.6151
R949 B.n262 B.n261 10.6151
R950 B.n265 B.n262 10.6151
R951 B.n266 B.n265 10.6151
R952 B.n269 B.n266 10.6151
R953 B.n271 B.n269 10.6151
R954 B.n272 B.n271 10.6151
R955 B.n618 B.n272 10.6151
R956 B.n546 B.n545 10.6151
R957 B.n546 B.n295 10.6151
R958 B.n556 B.n295 10.6151
R959 B.n557 B.n556 10.6151
R960 B.n558 B.n557 10.6151
R961 B.n558 B.n288 10.6151
R962 B.n568 B.n288 10.6151
R963 B.n569 B.n568 10.6151
R964 B.n570 B.n569 10.6151
R965 B.n570 B.n281 10.6151
R966 B.n581 B.n281 10.6151
R967 B.n582 B.n581 10.6151
R968 B.n584 B.n582 10.6151
R969 B.n584 B.n583 10.6151
R970 B.n583 B.n273 10.6151
R971 B.n595 B.n273 10.6151
R972 B.n596 B.n595 10.6151
R973 B.n597 B.n596 10.6151
R974 B.n598 B.n597 10.6151
R975 B.n600 B.n598 10.6151
R976 B.n601 B.n600 10.6151
R977 B.n602 B.n601 10.6151
R978 B.n603 B.n602 10.6151
R979 B.n605 B.n603 10.6151
R980 B.n606 B.n605 10.6151
R981 B.n607 B.n606 10.6151
R982 B.n608 B.n607 10.6151
R983 B.n610 B.n608 10.6151
R984 B.n611 B.n610 10.6151
R985 B.n612 B.n611 10.6151
R986 B.n613 B.n612 10.6151
R987 B.n615 B.n613 10.6151
R988 B.n616 B.n615 10.6151
R989 B.n617 B.n616 10.6151
R990 B.n539 B.n538 10.6151
R991 B.n538 B.n537 10.6151
R992 B.n537 B.n536 10.6151
R993 B.n536 B.n534 10.6151
R994 B.n534 B.n531 10.6151
R995 B.n531 B.n530 10.6151
R996 B.n530 B.n527 10.6151
R997 B.n527 B.n526 10.6151
R998 B.n526 B.n523 10.6151
R999 B.n523 B.n522 10.6151
R1000 B.n522 B.n519 10.6151
R1001 B.n519 B.n518 10.6151
R1002 B.n518 B.n515 10.6151
R1003 B.n515 B.n514 10.6151
R1004 B.n514 B.n511 10.6151
R1005 B.n511 B.n510 10.6151
R1006 B.n510 B.n507 10.6151
R1007 B.n507 B.n506 10.6151
R1008 B.n506 B.n503 10.6151
R1009 B.n503 B.n502 10.6151
R1010 B.n502 B.n499 10.6151
R1011 B.n499 B.n498 10.6151
R1012 B.n498 B.n495 10.6151
R1013 B.n495 B.n494 10.6151
R1014 B.n494 B.n491 10.6151
R1015 B.n491 B.n490 10.6151
R1016 B.n490 B.n487 10.6151
R1017 B.n487 B.n486 10.6151
R1018 B.n486 B.n483 10.6151
R1019 B.n483 B.n482 10.6151
R1020 B.n482 B.n479 10.6151
R1021 B.n479 B.n478 10.6151
R1022 B.n478 B.n475 10.6151
R1023 B.n475 B.n474 10.6151
R1024 B.n474 B.n471 10.6151
R1025 B.n471 B.n470 10.6151
R1026 B.n470 B.n467 10.6151
R1027 B.n467 B.n466 10.6151
R1028 B.n466 B.n463 10.6151
R1029 B.n463 B.n462 10.6151
R1030 B.n462 B.n459 10.6151
R1031 B.n457 B.n454 10.6151
R1032 B.n454 B.n453 10.6151
R1033 B.n453 B.n450 10.6151
R1034 B.n450 B.n449 10.6151
R1035 B.n449 B.n446 10.6151
R1036 B.n446 B.n445 10.6151
R1037 B.n445 B.n442 10.6151
R1038 B.n442 B.n441 10.6151
R1039 B.n441 B.n438 10.6151
R1040 B.n436 B.n433 10.6151
R1041 B.n433 B.n432 10.6151
R1042 B.n432 B.n429 10.6151
R1043 B.n429 B.n428 10.6151
R1044 B.n428 B.n425 10.6151
R1045 B.n425 B.n424 10.6151
R1046 B.n424 B.n421 10.6151
R1047 B.n421 B.n420 10.6151
R1048 B.n420 B.n417 10.6151
R1049 B.n417 B.n416 10.6151
R1050 B.n416 B.n413 10.6151
R1051 B.n413 B.n412 10.6151
R1052 B.n412 B.n409 10.6151
R1053 B.n409 B.n408 10.6151
R1054 B.n408 B.n405 10.6151
R1055 B.n405 B.n404 10.6151
R1056 B.n404 B.n401 10.6151
R1057 B.n401 B.n400 10.6151
R1058 B.n400 B.n397 10.6151
R1059 B.n397 B.n396 10.6151
R1060 B.n396 B.n393 10.6151
R1061 B.n393 B.n392 10.6151
R1062 B.n392 B.n389 10.6151
R1063 B.n389 B.n388 10.6151
R1064 B.n388 B.n385 10.6151
R1065 B.n385 B.n384 10.6151
R1066 B.n384 B.n381 10.6151
R1067 B.n381 B.n380 10.6151
R1068 B.n380 B.n377 10.6151
R1069 B.n377 B.n376 10.6151
R1070 B.n376 B.n373 10.6151
R1071 B.n373 B.n372 10.6151
R1072 B.n372 B.n369 10.6151
R1073 B.n369 B.n368 10.6151
R1074 B.n368 B.n365 10.6151
R1075 B.n365 B.n364 10.6151
R1076 B.n364 B.n361 10.6151
R1077 B.n361 B.n360 10.6151
R1078 B.n360 B.n357 10.6151
R1079 B.n357 B.n304 10.6151
R1080 B.n544 B.n304 10.6151
R1081 B.n550 B.n300 10.6151
R1082 B.n551 B.n550 10.6151
R1083 B.n552 B.n551 10.6151
R1084 B.n552 B.n292 10.6151
R1085 B.n562 B.n292 10.6151
R1086 B.n563 B.n562 10.6151
R1087 B.n564 B.n563 10.6151
R1088 B.n564 B.n284 10.6151
R1089 B.n575 B.n284 10.6151
R1090 B.n576 B.n575 10.6151
R1091 B.n577 B.n576 10.6151
R1092 B.n577 B.n277 10.6151
R1093 B.n588 B.n277 10.6151
R1094 B.n589 B.n588 10.6151
R1095 B.n590 B.n589 10.6151
R1096 B.n590 B.n0 10.6151
R1097 B.n651 B.n1 10.6151
R1098 B.n651 B.n650 10.6151
R1099 B.n650 B.n649 10.6151
R1100 B.n649 B.n10 10.6151
R1101 B.n643 B.n10 10.6151
R1102 B.n643 B.n642 10.6151
R1103 B.n642 B.n641 10.6151
R1104 B.n641 B.n16 10.6151
R1105 B.n635 B.n16 10.6151
R1106 B.n635 B.n634 10.6151
R1107 B.n634 B.n633 10.6151
R1108 B.n633 B.n24 10.6151
R1109 B.n627 B.n24 10.6151
R1110 B.n627 B.n626 10.6151
R1111 B.n626 B.n625 10.6151
R1112 B.n625 B.n31 10.6151
R1113 B.n170 B.n87 9.36635
R1114 B.n193 B.n84 9.36635
R1115 B.n459 B.n458 9.36635
R1116 B.n437 B.n436 9.36635
R1117 B.n560 B.t5 6.90099
R1118 B.n631 B.t9 6.90099
R1119 B.t2 B.n275 3.13708
R1120 B.t0 B.n8 3.13708
R1121 B.n657 B.n0 2.81026
R1122 B.n657 B.n1 2.81026
R1123 B.n173 B.n87 1.24928
R1124 B.n190 B.n84 1.24928
R1125 B.n458 B.n457 1.24928
R1126 B.n438 B.n437 1.24928
R1127 B.n579 B.t3 0.627817
R1128 B.n645 B.t1 0.627817
R1129 VP.n1 VP.t0 520.622
R1130 VP.n1 VP.t1 520.572
R1131 VP.n3 VP.t2 499.625
R1132 VP.n5 VP.t3 499.625
R1133 VP.n6 VP.n5 161.3
R1134 VP.n4 VP.n0 161.3
R1135 VP.n3 VP.n2 161.3
R1136 VP.n2 VP.n1 85.1545
R1137 VP.n4 VP.n3 24.1005
R1138 VP.n5 VP.n4 24.1005
R1139 VP.n2 VP.n0 0.189894
R1140 VP.n6 VP.n0 0.189894
R1141 VP VP.n6 0.0516364
R1142 VDD1 VDD1.n1 101.353
R1143 VDD1 VDD1.n0 64.0159
R1144 VDD1.n0 VDD1.t3 1.61551
R1145 VDD1.n0 VDD1.t2 1.61551
R1146 VDD1.n1 VDD1.t1 1.61551
R1147 VDD1.n1 VDD1.t0 1.61551
C0 VDD2 VTAIL 7.05594f
C1 VDD1 VP 3.28525f
C2 VN VTAIL 2.74624f
C3 VDD2 VDD1 0.559564f
C4 VDD2 VP 0.271636f
C5 VDD1 VN 0.147395f
C6 VN VP 4.84904f
C7 VDD2 VN 3.16126f
C8 VDD1 VTAIL 7.01467f
C9 VP VTAIL 2.76035f
C10 VDD2 B 2.703276f
C11 VDD1 B 6.42966f
C12 VTAIL B 8.892317f
C13 VN B 8.13474f
C14 VP B 4.85386f
C15 VDD1.t3 B 0.274475f
C16 VDD1.t2 B 0.274475f
C17 VDD1.n0 B 2.45957f
C18 VDD1.t1 B 0.274475f
C19 VDD1.t0 B 0.274475f
C20 VDD1.n1 B 3.08632f
C21 VP.n0 B 0.050994f
C22 VP.t1 B 1.21308f
C23 VP.t0 B 1.21313f
C24 VP.n1 B 1.90709f
C25 VP.n2 B 3.11831f
C26 VP.t2 B 1.19398f
C27 VP.n3 B 0.470765f
C28 VP.n4 B 0.011571f
C29 VP.t3 B 1.19398f
C30 VP.n5 B 0.470765f
C31 VP.n6 B 0.039518f
C32 VTAIL.t6 B 1.76771f
C33 VTAIL.n0 B 0.259157f
C34 VTAIL.t2 B 1.76771f
C35 VTAIL.n1 B 0.278973f
C36 VTAIL.t3 B 1.76771f
C37 VTAIL.n2 B 1.0856f
C38 VTAIL.t7 B 1.76771f
C39 VTAIL.n3 B 1.0856f
C40 VTAIL.t5 B 1.76771f
C41 VTAIL.n4 B 0.278977f
C42 VTAIL.t0 B 1.76771f
C43 VTAIL.n5 B 0.278977f
C44 VTAIL.t1 B 1.76771f
C45 VTAIL.n6 B 1.08561f
C46 VTAIL.t4 B 1.76771f
C47 VTAIL.n7 B 1.0596f
C48 VDD2.t0 B 0.277292f
C49 VDD2.t2 B 0.277292f
C50 VDD2.n0 B 3.09113f
C51 VDD2.t1 B 0.277292f
C52 VDD2.t3 B 0.277292f
C53 VDD2.n1 B 2.48452f
C54 VDD2.n2 B 3.52951f
C55 VN.t1 B 1.18309f
C56 VN.t3 B 1.18304f
C57 VN.n0 B 0.892706f
C58 VN.t2 B 1.18309f
C59 VN.t0 B 1.18304f
C60 VN.n1 B 1.88025f
.ends

