* NGSPICE file created from opamp_sample_0012.ext - technology: sky130A

.subckt opamp_sample_0012 GND VOUT VDD VN VP CS_BIAS DIFFPAIR_BIAS
X0 GND.t87 CS_BIAS.t24 VOUT.t25 GND.t41 sky130_fd_pr__nfet_01v8 ad=1.4898 pd=8.42 as=0.6303 ps=4.15 w=3.82 l=2.21
X1 VOUT.t24 CS_BIAS.t25 GND.t86 GND.t24 sky130_fd_pr__nfet_01v8 ad=0.6303 pd=4.15 as=0.6303 ps=4.15 w=3.82 l=2.21
X2 GND.t233 GND.t231 GND.t232 GND.t145 sky130_fd_pr__nfet_01v8 ad=1.4898 pd=8.42 as=0 ps=0 w=3.82 l=2.21
X3 a_n16148_7944.t5 a_n10279_8682.t10 a_n4238_7449.t0 VDD.t35 sky130_fd_pr__pfet_01v8 ad=0.55275 pd=3.68 as=1.3065 ps=7.48 w=3.35 l=5.36
X4 CS_BIAS.t3 CS_BIAS.t2 GND.t85 GND.t24 sky130_fd_pr__nfet_01v8 ad=0.6303 pd=4.15 as=0.6303 ps=4.15 w=3.82 l=2.21
X5 GND.t230 GND.t228 GND.t229 GND.t89 sky130_fd_pr__nfet_01v8 ad=1.4898 pd=8.42 as=0 ps=0 w=3.82 l=2.21
X6 GND.t227 GND.t225 VP.t7 GND.t226 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X7 GND.t224 GND.t222 VN.t7 GND.t223 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X8 VDD.t105 VDD.t103 VDD.t104 VDD.t94 sky130_fd_pr__pfet_01v8 ad=1.3065 pd=7.48 as=0 ps=0 w=3.35 l=5.36
X9 a_n10279_8682.t0 VP.t8 a_n1140_n227.t2 GND.t0 sky130_fd_pr__nfet_01v8 ad=0.9282 pd=5.54 as=0.9282 ps=5.54 w=2.38 l=4.6
X10 VDD.t137 a_n16148_7944.t6 VOUT.t20 VDD.t108 sky130_fd_pr__pfet_01v8 ad=0.8151 pd=4.96 as=0.34485 ps=2.42 w=2.09 l=2.93
X11 VDD.t136 a_n16148_7944.t7 VOUT.t3 VDD.t106 sky130_fd_pr__pfet_01v8 ad=0.34485 pd=2.42 as=0.34485 ps=2.42 w=2.09 l=2.93
X12 VDD.t102 VDD.t100 VDD.t101 VDD.t90 sky130_fd_pr__pfet_01v8 ad=0.8151 pd=4.96 as=0 ps=0 w=2.09 l=2.93
X13 VOUT.t23 CS_BIAS.t26 GND.t84 GND.t14 sky130_fd_pr__nfet_01v8 ad=0.6303 pd=4.15 as=0.6303 ps=4.15 w=3.82 l=2.21
X14 CS_BIAS.t1 CS_BIAS.t0 GND.t83 GND.t14 sky130_fd_pr__nfet_01v8 ad=0.6303 pd=4.15 as=0.6303 ps=4.15 w=3.82 l=2.21
X15 GND.t82 CS_BIAS.t27 VOUT.t45 GND.t41 sky130_fd_pr__nfet_01v8 ad=1.4898 pd=8.42 as=0.6303 ps=4.15 w=3.82 l=2.21
X16 VOUT.t44 CS_BIAS.t28 GND.t81 GND.t39 sky130_fd_pr__nfet_01v8 ad=0.6303 pd=4.15 as=0.6303 ps=4.15 w=3.82 l=2.21
X17 VOUT.t43 CS_BIAS.t29 GND.t80 GND.t39 sky130_fd_pr__nfet_01v8 ad=0.6303 pd=4.15 as=0.6303 ps=4.15 w=3.82 l=2.21
X18 VOUT.t2 a_n16148_7944.t8 VDD.t135 VDD.t128 sky130_fd_pr__pfet_01v8 ad=0.34485 pd=2.42 as=0.8151 ps=4.96 w=2.09 l=2.93
X19 VDD.t134 a_n16148_7944.t9 VOUT.t10 VDD.t108 sky130_fd_pr__pfet_01v8 ad=0.8151 pd=4.96 as=0.34485 ps=2.42 w=2.09 l=2.93
X20 VOUT.t42 CS_BIAS.t30 GND.t79 GND.t14 sky130_fd_pr__nfet_01v8 ad=0.6303 pd=4.15 as=0.6303 ps=4.15 w=3.82 l=2.21
X21 GND.t78 CS_BIAS.t31 VOUT.t41 GND.t8 sky130_fd_pr__nfet_01v8 ad=0.6303 pd=4.15 as=0.6303 ps=4.15 w=3.82 l=2.21
X22 VDD.t133 a_n16148_7944.t10 VOUT.t18 VDD.t106 sky130_fd_pr__pfet_01v8 ad=0.34485 pd=2.42 as=0.34485 ps=2.42 w=2.09 l=2.93
X23 GND.t221 GND.t219 GND.t220 GND.t89 sky130_fd_pr__nfet_01v8 ad=1.4898 pd=8.42 as=0 ps=0 w=3.82 l=2.21
X24 VDD.t99 VDD.t97 VDD.t98 VDD.t90 sky130_fd_pr__pfet_01v8 ad=0.8151 pd=4.96 as=0 ps=0 w=2.09 l=2.93
X25 a_n16148_7944.t4 a_n10279_8682.t11 a_n4238_7449.t2 VDD.t17 sky130_fd_pr__pfet_01v8 ad=0.55275 pd=3.68 as=1.3065 ps=7.48 w=3.35 l=5.36
X26 VDD.t132 a_n16148_7944.t11 VOUT.t6 VDD.t125 sky130_fd_pr__pfet_01v8 ad=0.34485 pd=2.42 as=0.34485 ps=2.42 w=2.09 l=2.93
X27 a_n4238_7449.t5 a_n10279_8682.t12 VDD.t37 VDD.t36 sky130_fd_pr__pfet_01v8 ad=1.3065 pd=7.48 as=0.55275 ps=3.68 w=3.35 l=5.36
X28 GND.t218 GND.t216 GND.t217 GND.t145 sky130_fd_pr__nfet_01v8 ad=1.4898 pd=8.42 as=0 ps=0 w=3.82 l=2.21
X29 GND.t77 CS_BIAS.t32 VOUT.t40 GND.t11 sky130_fd_pr__nfet_01v8 ad=0.6303 pd=4.15 as=0.6303 ps=4.15 w=3.82 l=2.21
X30 GND.t215 GND.t213 GND.t214 GND.t109 sky130_fd_pr__nfet_01v8 ad=1.4898 pd=8.42 as=0 ps=0 w=3.82 l=2.21
X31 VOUT.t19 a_n16148_7944.t12 VDD.t131 VDD.t128 sky130_fd_pr__pfet_01v8 ad=0.34485 pd=2.42 as=0.8151 ps=4.96 w=2.09 l=2.93
X32 VDD.t96 VDD.t93 VDD.t95 VDD.t94 sky130_fd_pr__pfet_01v8 ad=1.3065 pd=7.48 as=0 ps=0 w=3.35 l=5.36
X33 GND.t212 GND.t210 GND.t211 GND.t122 sky130_fd_pr__nfet_01v8 ad=1.4898 pd=8.42 as=0 ps=0 w=3.82 l=2.21
X34 GND.t76 CS_BIAS.t33 VOUT.t31 GND.t11 sky130_fd_pr__nfet_01v8 ad=0.6303 pd=4.15 as=0.6303 ps=4.15 w=3.82 l=2.21
X35 VDD.t92 VDD.t89 VDD.t91 VDD.t90 sky130_fd_pr__pfet_01v8 ad=0.8151 pd=4.96 as=0 ps=0 w=2.09 l=2.93
X36 VOUT.t30 CS_BIAS.t34 GND.t75 GND.t24 sky130_fd_pr__nfet_01v8 ad=0.6303 pd=4.15 as=0.6303 ps=4.15 w=3.82 l=2.21
X37 VOUT.t29 CS_BIAS.t35 GND.t74 GND.t24 sky130_fd_pr__nfet_01v8 ad=0.6303 pd=4.15 as=0.6303 ps=4.15 w=3.82 l=2.21
X38 VDD.t130 a_n16148_7944.t13 VOUT.t5 VDD.t125 sky130_fd_pr__pfet_01v8 ad=0.34485 pd=2.42 as=0.34485 ps=2.42 w=2.09 l=2.93
X39 GND.t73 CS_BIAS.t36 VOUT.t28 GND.t31 sky130_fd_pr__nfet_01v8 ad=0.6303 pd=4.15 as=0.6303 ps=4.15 w=3.82 l=2.21
X40 GND.t72 CS_BIAS.t37 VOUT.t27 GND.t20 sky130_fd_pr__nfet_01v8 ad=0.6303 pd=4.15 as=0.6303 ps=4.15 w=3.82 l=2.21
X41 VOUT.t26 CS_BIAS.t38 GND.t71 GND.t16 sky130_fd_pr__nfet_01v8 ad=0.6303 pd=4.15 as=1.4898 ps=8.42 w=3.82 l=2.21
X42 a_n1140_n227.t0 DIFFPAIR_BIAS.t2 a_53_n2194# GND.t2 sky130_fd_pr__nfet_01v8 ad=0.8619 pd=5.2 as=0.8619 ps=5.2 w=2.21 l=3.05
X43 GND.t209 GND.t207 GND.t208 GND.t109 sky130_fd_pr__nfet_01v8 ad=1.4898 pd=8.42 as=0 ps=0 w=3.82 l=2.21
X44 VOUT.t4 a_n16148_7944.t14 VDD.t129 VDD.t128 sky130_fd_pr__pfet_01v8 ad=0.34485 pd=2.42 as=0.8151 ps=4.96 w=2.09 l=2.93
X45 VOUT.t67 CS_BIAS.t39 GND.t70 GND.t22 sky130_fd_pr__nfet_01v8 ad=0.6303 pd=4.15 as=0.6303 ps=4.15 w=3.82 l=2.21
X46 GND.t69 CS_BIAS.t40 VOUT.t66 GND.t4 sky130_fd_pr__nfet_01v8 ad=1.4898 pd=8.42 as=0.6303 ps=4.15 w=3.82 l=2.21
X47 a_n10357_8879.t3 a_n10279_8682.t8 a_n10279_8682.t9 VDD.t35 sky130_fd_pr__pfet_01v8 ad=0.55275 pd=3.68 as=1.3065 ps=7.48 w=3.35 l=5.36
X48 VN.t6 GND.t204 GND.t206 GND.t205 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X49 GND.t203 GND.t201 GND.t202 GND.t89 sky130_fd_pr__nfet_01v8 ad=1.4898 pd=8.42 as=0 ps=0 w=3.82 l=2.21
X50 VOUT.t17 a_n16148_7944.t15 VDD.t127 VDD.t122 sky130_fd_pr__pfet_01v8 ad=0.34485 pd=2.42 as=0.34485 ps=2.42 w=2.09 l=2.93
X51 VDD.t126 a_n16148_7944.t16 VOUT.t16 VDD.t125 sky130_fd_pr__pfet_01v8 ad=0.34485 pd=2.42 as=0.34485 ps=2.42 w=2.09 l=2.93
X52 GND.t200 GND.t198 GND.t199 GND.t89 sky130_fd_pr__nfet_01v8 ad=1.4898 pd=8.42 as=0 ps=0 w=3.82 l=2.21
X53 GND.t197 GND.t194 GND.t196 GND.t195 sky130_fd_pr__nfet_01v8 ad=0.8619 pd=5.2 as=0 ps=0 w=2.21 l=3.05
X54 GND.t193 GND.t191 GND.t192 GND.t145 sky130_fd_pr__nfet_01v8 ad=1.4898 pd=8.42 as=0 ps=0 w=3.82 l=2.21
X55 GND.t68 CS_BIAS.t41 VOUT.t65 GND.t20 sky130_fd_pr__nfet_01v8 ad=0.6303 pd=4.15 as=0.6303 ps=4.15 w=3.82 l=2.21
X56 VOUT.t64 CS_BIAS.t42 GND.t67 GND.t22 sky130_fd_pr__nfet_01v8 ad=0.6303 pd=4.15 as=0.6303 ps=4.15 w=3.82 l=2.21
X57 GND.t190 GND.t188 GND.t189 GND.t170 sky130_fd_pr__nfet_01v8 ad=0.9282 pd=5.54 as=0 ps=0 w=2.38 l=4.6
X58 GND.t66 CS_BIAS.t43 VOUT.t63 GND.t4 sky130_fd_pr__nfet_01v8 ad=1.4898 pd=8.42 as=0.6303 ps=4.15 w=3.82 l=2.21
X59 VDD.t34 a_n10279_8682.t13 a_n10357_8879.t11 VDD.t33 sky130_fd_pr__pfet_01v8 ad=0.55275 pd=3.68 as=1.3065 ps=7.48 w=3.35 l=5.36
X60 GND.t65 CS_BIAS.t16 CS_BIAS.t17 GND.t4 sky130_fd_pr__nfet_01v8 ad=1.4898 pd=8.42 as=0.6303 ps=4.15 w=3.82 l=2.21
X61 GND.t64 CS_BIAS.t44 VOUT.t62 GND.t41 sky130_fd_pr__nfet_01v8 ad=1.4898 pd=8.42 as=0.6303 ps=4.15 w=3.82 l=2.21
X62 a_n4238_7449.t9 a_n10279_8682.t14 a_n16148_7944.t3 VDD.t28 sky130_fd_pr__pfet_01v8 ad=1.3065 pd=7.48 as=0.55275 ps=3.68 w=3.35 l=5.36
X63 GND.t53 CS_BIAS.t18 CS_BIAS.t19 GND.t41 sky130_fd_pr__nfet_01v8 ad=1.4898 pd=8.42 as=0.6303 ps=4.15 w=3.82 l=2.21
X64 GND.t63 CS_BIAS.t45 VOUT.t61 GND.t4 sky130_fd_pr__nfet_01v8 ad=1.4898 pd=8.42 as=0.6303 ps=4.15 w=3.82 l=2.21
X65 GND.t62 CS_BIAS.t46 VOUT.t60 GND.t20 sky130_fd_pr__nfet_01v8 ad=0.6303 pd=4.15 as=0.6303 ps=4.15 w=3.82 l=2.21
X66 VN.t5 GND.t185 GND.t187 GND.t186 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X67 VOUT.t11 a_n16148_7944.t17 VDD.t124 VDD.t122 sky130_fd_pr__pfet_01v8 ad=0.34485 pd=2.42 as=0.34485 ps=2.42 w=2.09 l=2.93
X68 VP.t6 GND.t182 GND.t184 GND.t183 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X69 a_n4238_7449.t7 a_n10279_8682.t15 VDD.t32 VDD.t31 sky130_fd_pr__pfet_01v8 ad=0.55275 pd=3.68 as=0.55275 ps=3.68 w=3.35 l=5.36
X70 a_10485_8879# a_10485_8879# a_10485_8879# VDD.t0 sky130_fd_pr__pfet_01v8 ad=1.3065 pd=7.48 as=2.613 ps=14.96 w=3.35 l=5.36
X71 GND.t61 CS_BIAS.t47 VOUT.t59 GND.t31 sky130_fd_pr__nfet_01v8 ad=0.6303 pd=4.15 as=0.6303 ps=4.15 w=3.82 l=2.21
X72 VOUT.t58 CS_BIAS.t48 GND.t60 GND.t39 sky130_fd_pr__nfet_01v8 ad=0.6303 pd=4.15 as=0.6303 ps=4.15 w=3.82 l=2.21
X73 VOUT.t13 a_n16148_7944.t18 VDD.t123 VDD.t122 sky130_fd_pr__pfet_01v8 ad=0.34485 pd=2.42 as=0.34485 ps=2.42 w=2.09 l=2.93
X74 CS_BIAS.t15 CS_BIAS.t14 GND.t59 GND.t39 sky130_fd_pr__nfet_01v8 ad=0.6303 pd=4.15 as=0.6303 ps=4.15 w=3.82 l=2.21
X75 VOUT.t73 CS_BIAS.t49 GND.t58 GND.t6 sky130_fd_pr__nfet_01v8 ad=0.6303 pd=4.15 as=1.4898 ps=8.42 w=3.82 l=2.21
X76 VDD.t121 a_n16148_7944.t19 VOUT.t8 VDD.t117 sky130_fd_pr__pfet_01v8 ad=0.8151 pd=4.96 as=0.34485 ps=2.42 w=2.09 l=2.93
X77 VP.t5 GND.t179 GND.t181 GND.t180 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X78 VN.t4 GND.t176 GND.t178 GND.t177 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X79 VDD.t30 a_n10279_8682.t16 a_n4238_7449.t10 VDD.t29 sky130_fd_pr__pfet_01v8 ad=0.55275 pd=3.68 as=0.55275 ps=3.68 w=3.35 l=5.36
X80 VOUT.t72 CS_BIAS.t50 GND.t57 GND.t22 sky130_fd_pr__nfet_01v8 ad=0.6303 pd=4.15 as=0.6303 ps=4.15 w=3.82 l=2.21
X81 GND.t175 GND.t173 GND.t174 GND.t122 sky130_fd_pr__nfet_01v8 ad=1.4898 pd=8.42 as=0 ps=0 w=3.82 l=2.21
X82 VOUT.t71 CS_BIAS.t51 GND.t56 GND.t6 sky130_fd_pr__nfet_01v8 ad=0.6303 pd=4.15 as=1.4898 ps=8.42 w=3.82 l=2.21
X83 GND.t55 CS_BIAS.t52 VOUT.t70 GND.t41 sky130_fd_pr__nfet_01v8 ad=1.4898 pd=8.42 as=0.6303 ps=4.15 w=3.82 l=2.21
X84 VDD.t88 VDD.t86 VDD.t87 VDD.t50 sky130_fd_pr__pfet_01v8 ad=1.3065 pd=7.48 as=0 ps=0 w=3.35 l=5.36
X85 VOUT.t69 CS_BIAS.t53 GND.t54 GND.t39 sky130_fd_pr__nfet_01v8 ad=0.6303 pd=4.15 as=0.6303 ps=4.15 w=3.82 l=2.21
X86 VOUT.t84 a_n4238_7449.t12 sky130_fd_pr__cap_mim_m3_1 l=11.53 w=6.75
X87 GND.t172 GND.t169 GND.t171 GND.t170 sky130_fd_pr__nfet_01v8 ad=0.9282 pd=5.54 as=0 ps=0 w=2.38 l=4.6
X88 VDD.t85 VDD.t83 VDD.t84 VDD.t74 sky130_fd_pr__pfet_01v8 ad=0.8151 pd=4.96 as=0 ps=0 w=2.09 l=2.93
X89 a_n10279_8682.t1 VP.t9 a_n1140_n227.t1 GND.t1 sky130_fd_pr__nfet_01v8 ad=0.9282 pd=5.54 as=0.9282 ps=5.54 w=2.38 l=4.6
X90 VDD.t120 a_n16148_7944.t20 VOUT.t7 VDD.t117 sky130_fd_pr__pfet_01v8 ad=0.8151 pd=4.96 as=0.34485 ps=2.42 w=2.09 l=2.93
X91 VN.t3 GND.t166 GND.t168 GND.t167 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X92 VP.t4 GND.t163 GND.t165 GND.t164 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X93 VOUT.t79 CS_BIAS.t54 GND.t52 GND.t16 sky130_fd_pr__nfet_01v8 ad=0.6303 pd=4.15 as=1.4898 ps=8.42 w=3.82 l=2.21
X94 GND.t162 GND.t160 GND.t161 GND.t122 sky130_fd_pr__nfet_01v8 ad=1.4898 pd=8.42 as=0 ps=0 w=3.82 l=2.21
X95 GND.t159 GND.t157 GND.t158 GND.t145 sky130_fd_pr__nfet_01v8 ad=1.4898 pd=8.42 as=0 ps=0 w=3.82 l=2.21
X96 GND.t156 GND.t154 GND.t155 GND.t135 sky130_fd_pr__nfet_01v8 ad=0.9282 pd=5.54 as=0 ps=0 w=2.38 l=4.6
X97 a_n10279_8682.t7 a_n10279_8682.t6 a_n10357_8879.t2 VDD.t28 sky130_fd_pr__pfet_01v8 ad=1.3065 pd=7.48 as=0.55275 ps=3.68 w=3.35 l=5.36
X98 GND.t51 CS_BIAS.t55 VOUT.t78 GND.t8 sky130_fd_pr__nfet_01v8 ad=0.6303 pd=4.15 as=0.6303 ps=4.15 w=3.82 l=2.21
X99 VDD.t27 a_n10279_8682.t17 a_n10357_8879.t10 VDD.t26 sky130_fd_pr__pfet_01v8 ad=0.55275 pd=3.68 as=0.55275 ps=3.68 w=3.35 l=5.36
X100 VDD.t82 VDD.t80 VDD.t81 VDD.t74 sky130_fd_pr__pfet_01v8 ad=0.8151 pd=4.96 as=0 ps=0 w=2.09 l=2.93
X101 a_n10357_8879.t9 a_n10279_8682.t18 VDD.t25 VDD.t24 sky130_fd_pr__pfet_01v8 ad=1.3065 pd=7.48 as=0.55275 ps=3.68 w=3.35 l=5.36
X102 VOUT.t77 CS_BIAS.t56 GND.t50 GND.t6 sky130_fd_pr__nfet_01v8 ad=0.6303 pd=4.15 as=1.4898 ps=8.42 w=3.82 l=2.21
X103 VP.t3 GND.t151 GND.t153 GND.t152 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X104 VOUT.t76 CS_BIAS.t57 GND.t49 GND.t14 sky130_fd_pr__nfet_01v8 ad=0.6303 pd=4.15 as=0.6303 ps=4.15 w=3.82 l=2.21
X105 VOUT.t12 a_n16148_7944.t21 VDD.t119 VDD.t114 sky130_fd_pr__pfet_01v8 ad=0.34485 pd=2.42 as=0.34485 ps=2.42 w=2.09 l=2.93
X106 VDD.t118 a_n16148_7944.t22 VOUT.t0 VDD.t117 sky130_fd_pr__pfet_01v8 ad=0.8151 pd=4.96 as=0.34485 ps=2.42 w=2.09 l=2.93
X107 GND.t48 CS_BIAS.t58 VOUT.t75 GND.t31 sky130_fd_pr__nfet_01v8 ad=0.6303 pd=4.15 as=0.6303 ps=4.15 w=3.82 l=2.21
X108 VOUT.t85 a_n4238_7449.t12 sky130_fd_pr__cap_mim_m3_1 l=11.53 w=6.75
X109 GND.t150 GND.t148 GND.t149 GND.t145 sky130_fd_pr__nfet_01v8 ad=1.4898 pd=8.42 as=0 ps=0 w=3.82 l=2.21
X110 VDD.t79 VDD.t77 VDD.t78 VDD.t43 sky130_fd_pr__pfet_01v8 ad=1.3065 pd=7.48 as=0 ps=0 w=3.35 l=5.36
X111 a_n10357_8879.t8 a_n10279_8682.t19 VDD.t23 VDD.t22 sky130_fd_pr__pfet_01v8 ad=0.55275 pd=3.68 as=0.55275 ps=3.68 w=3.35 l=5.36
X112 GND.t147 GND.t144 GND.t146 GND.t145 sky130_fd_pr__nfet_01v8 ad=1.4898 pd=8.42 as=0 ps=0 w=3.82 l=2.21
X113 VDD.t76 VDD.t73 VDD.t75 VDD.t74 sky130_fd_pr__pfet_01v8 ad=0.8151 pd=4.96 as=0 ps=0 w=2.09 l=2.93
X114 GND.t143 GND.t141 GND.t142 GND.t109 sky130_fd_pr__nfet_01v8 ad=1.4898 pd=8.42 as=0 ps=0 w=3.82 l=2.21
X115 VOUT.t74 CS_BIAS.t59 GND.t47 GND.t16 sky130_fd_pr__nfet_01v8 ad=0.6303 pd=4.15 as=1.4898 ps=8.42 w=3.82 l=2.21
X116 VDD.t21 a_n10279_8682.t20 a_n4238_7449.t3 VDD.t20 sky130_fd_pr__pfet_01v8 ad=0.55275 pd=3.68 as=1.3065 ps=7.48 w=3.35 l=5.36
X117 GND.t46 CS_BIAS.t60 VOUT.t49 GND.t8 sky130_fd_pr__nfet_01v8 ad=0.6303 pd=4.15 as=0.6303 ps=4.15 w=3.82 l=2.21
X118 VOUT.t48 CS_BIAS.t61 GND.t45 GND.t14 sky130_fd_pr__nfet_01v8 ad=0.6303 pd=4.15 as=0.6303 ps=4.15 w=3.82 l=2.21
X119 VOUT.t14 a_n16148_7944.t23 VDD.t116 VDD.t114 sky130_fd_pr__pfet_01v8 ad=0.34485 pd=2.42 as=0.34485 ps=2.42 w=2.09 l=2.93
X120 GND.t44 CS_BIAS.t62 VOUT.t47 GND.t20 sky130_fd_pr__nfet_01v8 ad=0.6303 pd=4.15 as=0.6303 ps=4.15 w=3.82 l=2.21
X121 GND.t140 GND.t138 GND.t139 GND.t89 sky130_fd_pr__nfet_01v8 ad=1.4898 pd=8.42 as=0 ps=0 w=3.82 l=2.21
X122 GND.t43 CS_BIAS.t10 CS_BIAS.t11 GND.t20 sky130_fd_pr__nfet_01v8 ad=0.6303 pd=4.15 as=0.6303 ps=4.15 w=3.82 l=2.21
X123 a_n16148_7944.t1 VN.t8 a_n1140_n227.t4 GND.t1 sky130_fd_pr__nfet_01v8 ad=0.9282 pd=5.54 as=0.9282 ps=5.54 w=2.38 l=4.6
X124 GND.t42 CS_BIAS.t63 VOUT.t46 GND.t41 sky130_fd_pr__nfet_01v8 ad=1.4898 pd=8.42 as=0.6303 ps=4.15 w=3.82 l=2.21
X125 VOUT.t36 CS_BIAS.t64 GND.t40 GND.t39 sky130_fd_pr__nfet_01v8 ad=0.6303 pd=4.15 as=0.6303 ps=4.15 w=3.82 l=2.21
X126 VDD.t19 a_n10279_8682.t21 a_n4238_7449.t8 VDD.t18 sky130_fd_pr__pfet_01v8 ad=0.55275 pd=3.68 as=1.3065 ps=7.48 w=3.35 l=5.36
X127 GND.t38 CS_BIAS.t65 VOUT.t35 GND.t11 sky130_fd_pr__nfet_01v8 ad=0.6303 pd=4.15 as=0.6303 ps=4.15 w=3.82 l=2.21
X128 GND.t137 GND.t134 GND.t136 GND.t135 sky130_fd_pr__nfet_01v8 ad=0.9282 pd=5.54 as=0 ps=0 w=2.38 l=4.6
X129 a_n10357_8879.t1 a_n10279_8682.t4 a_n10279_8682.t5 VDD.t17 sky130_fd_pr__pfet_01v8 ad=0.55275 pd=3.68 as=1.3065 ps=7.48 w=3.35 l=5.36
X130 VOUT.t81 a_n16148_7944.t24 VDD.t115 VDD.t114 sky130_fd_pr__pfet_01v8 ad=0.34485 pd=2.42 as=0.34485 ps=2.42 w=2.09 l=2.93
X131 GND.t37 CS_BIAS.t66 VOUT.t34 GND.t11 sky130_fd_pr__nfet_01v8 ad=0.6303 pd=4.15 as=0.6303 ps=4.15 w=3.82 l=2.21
X132 VOUT.t33 CS_BIAS.t67 GND.t36 GND.t24 sky130_fd_pr__nfet_01v8 ad=0.6303 pd=4.15 as=0.6303 ps=4.15 w=3.82 l=2.21
X133 GND.t35 CS_BIAS.t68 VOUT.t32 GND.t31 sky130_fd_pr__nfet_01v8 ad=0.6303 pd=4.15 as=0.6303 ps=4.15 w=3.82 l=2.21
X134 GND.t34 CS_BIAS.t12 CS_BIAS.t13 GND.t31 sky130_fd_pr__nfet_01v8 ad=0.6303 pd=4.15 as=0.6303 ps=4.15 w=3.82 l=2.21
X135 VDD.t16 a_n10279_8682.t22 a_n10357_8879.t7 VDD.t15 sky130_fd_pr__pfet_01v8 ad=0.55275 pd=3.68 as=1.3065 ps=7.48 w=3.35 l=5.36
X136 VDD.t14 a_n10279_8682.t23 a_n4238_7449.t11 VDD.t13 sky130_fd_pr__pfet_01v8 ad=0.55275 pd=3.68 as=0.55275 ps=3.68 w=3.35 l=5.36
X137 VDD.t72 VDD.t70 VDD.t71 VDD.t61 sky130_fd_pr__pfet_01v8 ad=0.8151 pd=4.96 as=0 ps=0 w=2.09 l=2.93
X138 VOUT.t55 CS_BIAS.t69 GND.t33 GND.t16 sky130_fd_pr__nfet_01v8 ad=0.6303 pd=4.15 as=1.4898 ps=8.42 w=3.82 l=2.21
X139 GND.t32 CS_BIAS.t70 VOUT.t54 GND.t31 sky130_fd_pr__nfet_01v8 ad=0.6303 pd=4.15 as=0.6303 ps=4.15 w=3.82 l=2.21
X140 GND.t30 CS_BIAS.t71 VOUT.t53 GND.t8 sky130_fd_pr__nfet_01v8 ad=0.6303 pd=4.15 as=0.6303 ps=4.15 w=3.82 l=2.21
X141 VOUT.t52 CS_BIAS.t72 GND.t29 GND.t22 sky130_fd_pr__nfet_01v8 ad=0.6303 pd=4.15 as=0.6303 ps=4.15 w=3.82 l=2.21
X142 GND.t133 GND.t131 GND.t132 GND.t122 sky130_fd_pr__nfet_01v8 ad=1.4898 pd=8.42 as=0 ps=0 w=3.82 l=2.21
X143 VOUT.t39 CS_BIAS.t73 GND.t28 GND.t6 sky130_fd_pr__nfet_01v8 ad=0.6303 pd=4.15 as=1.4898 ps=8.42 w=3.82 l=2.21
X144 GND.t130 GND.t128 GND.t129 GND.t109 sky130_fd_pr__nfet_01v8 ad=1.4898 pd=8.42 as=0 ps=0 w=3.82 l=2.21
X145 CS_BIAS.t7 CS_BIAS.t6 GND.t27 GND.t22 sky130_fd_pr__nfet_01v8 ad=0.6303 pd=4.15 as=0.6303 ps=4.15 w=3.82 l=2.21
X146 CS_BIAS.t5 CS_BIAS.t4 GND.t26 GND.t6 sky130_fd_pr__nfet_01v8 ad=0.6303 pd=4.15 as=1.4898 ps=8.42 w=3.82 l=2.21
X147 GND.t127 GND.t125 GND.t126 GND.t122 sky130_fd_pr__nfet_01v8 ad=1.4898 pd=8.42 as=0 ps=0 w=3.82 l=2.21
X148 GND.t124 GND.t121 GND.t123 GND.t122 sky130_fd_pr__nfet_01v8 ad=1.4898 pd=8.42 as=0 ps=0 w=3.82 l=2.21
X149 a_n10279_8682.t3 a_n10279_8682.t2 a_n10357_8879.t0 VDD.t12 sky130_fd_pr__pfet_01v8 ad=1.3065 pd=7.48 as=0.55275 ps=3.68 w=3.35 l=5.36
X150 VOUT.t38 CS_BIAS.t74 GND.t25 GND.t24 sky130_fd_pr__nfet_01v8 ad=0.6303 pd=4.15 as=0.6303 ps=4.15 w=3.82 l=2.21
X151 VDD.t69 VDD.t67 VDD.t68 VDD.t61 sky130_fd_pr__pfet_01v8 ad=0.8151 pd=4.96 as=0 ps=0 w=2.09 l=2.93
X152 DIFFPAIR_BIAS.t1 DIFFPAIR_BIAS.t0 a_n819_n2194# GND.t3 sky130_fd_pr__nfet_01v8 ad=0.8619 pd=5.2 as=0.8619 ps=5.2 w=2.21 l=3.05
X153 VOUT.t82 a_n16148_7944.t25 VDD.t113 VDD.t110 sky130_fd_pr__pfet_01v8 ad=0.34485 pd=2.42 as=0.8151 ps=4.96 w=2.09 l=2.93
X154 VOUT.t37 CS_BIAS.t75 GND.t23 GND.t22 sky130_fd_pr__nfet_01v8 ad=0.6303 pd=4.15 as=0.6303 ps=4.15 w=3.82 l=2.21
X155 GND.t21 CS_BIAS.t76 VOUT.t50 GND.t20 sky130_fd_pr__nfet_01v8 ad=0.6303 pd=4.15 as=0.6303 ps=4.15 w=3.82 l=2.21
X156 VOUT.t56 CS_BIAS.t77 GND.t19 GND.t16 sky130_fd_pr__nfet_01v8 ad=0.6303 pd=4.15 as=1.4898 ps=8.42 w=3.82 l=2.21
X157 GND.t120 GND.t118 VP.t2 GND.t119 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X158 CS_BIAS.t9 CS_BIAS.t8 GND.t17 GND.t16 sky130_fd_pr__nfet_01v8 ad=0.6303 pd=4.15 as=1.4898 ps=8.42 w=3.82 l=2.21
X159 GND.t18 CS_BIAS.t78 VOUT.t57 GND.t4 sky130_fd_pr__nfet_01v8 ad=1.4898 pd=8.42 as=0.6303 ps=4.15 w=3.82 l=2.21
X160 VOUT.t51 CS_BIAS.t79 GND.t15 GND.t14 sky130_fd_pr__nfet_01v8 ad=0.6303 pd=4.15 as=0.6303 ps=4.15 w=3.82 l=2.21
X161 a_n4238_7449.t4 a_n10279_8682.t24 a_n16148_7944.t2 VDD.t12 sky130_fd_pr__pfet_01v8 ad=1.3065 pd=7.48 as=0.55275 ps=3.68 w=3.35 l=5.36
X162 VDD.t66 VDD.t64 VDD.t65 VDD.t54 sky130_fd_pr__pfet_01v8 ad=1.3065 pd=7.48 as=0 ps=0 w=3.35 l=5.36
X163 VDD.t63 VDD.t60 VDD.t62 VDD.t61 sky130_fd_pr__pfet_01v8 ad=0.8151 pd=4.96 as=0 ps=0 w=2.09 l=2.93
X164 VDD.t59 VDD.t57 VDD.t58 VDD.t39 sky130_fd_pr__pfet_01v8 ad=0.8151 pd=4.96 as=0 ps=0 w=2.09 l=2.93
X165 VOUT.t9 a_n16148_7944.t26 VDD.t112 VDD.t110 sky130_fd_pr__pfet_01v8 ad=0.34485 pd=2.42 as=0.8151 ps=4.96 w=2.09 l=2.93
X166 GND.t117 GND.t115 VN.t2 GND.t116 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X167 VDD.t56 VDD.t53 VDD.t55 VDD.t54 sky130_fd_pr__pfet_01v8 ad=1.3065 pd=7.48 as=0 ps=0 w=3.35 l=5.36
X168 a_n11713_8879# a_n11713_8879# a_n11713_8879# VDD.t1 sky130_fd_pr__pfet_01v8 ad=1.3065 pd=7.48 as=2.613 ps=14.96 w=3.35 l=5.36
X169 GND.t94 GND.t92 VP.t1 GND.t93 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X170 VDD.t52 VDD.t49 VDD.t51 VDD.t50 sky130_fd_pr__pfet_01v8 ad=1.3065 pd=7.48 as=0 ps=0 w=3.35 l=5.36
X171 GND.t114 GND.t112 GND.t113 GND.t109 sky130_fd_pr__nfet_01v8 ad=1.4898 pd=8.42 as=0 ps=0 w=3.82 l=2.21
X172 VDD.t48 VDD.t46 VDD.t47 VDD.t39 sky130_fd_pr__pfet_01v8 ad=0.8151 pd=4.96 as=0 ps=0 w=2.09 l=2.93
X173 VDD.t45 VDD.t42 VDD.t44 VDD.t43 sky130_fd_pr__pfet_01v8 ad=1.3065 pd=7.48 as=0 ps=0 w=3.35 l=5.36
X174 GND.t111 GND.t108 GND.t110 GND.t109 sky130_fd_pr__nfet_01v8 ad=1.4898 pd=8.42 as=0 ps=0 w=3.82 l=2.21
X175 a_n16148_7944.t0 VN.t9 a_n1140_n227.t3 GND.t0 sky130_fd_pr__nfet_01v8 ad=0.9282 pd=5.54 as=0.9282 ps=5.54 w=2.38 l=4.6
X176 VOUT.t1 a_n16148_7944.t27 VDD.t111 VDD.t110 sky130_fd_pr__pfet_01v8 ad=0.34485 pd=2.42 as=0.8151 ps=4.96 w=2.09 l=2.93
X177 GND.t107 GND.t105 VN.t1 GND.t106 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X178 GND.t104 GND.t102 VP.t0 GND.t103 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X179 GND.t13 CS_BIAS.t80 VOUT.t22 GND.t11 sky130_fd_pr__nfet_01v8 ad=0.6303 pd=4.15 as=0.6303 ps=4.15 w=3.82 l=2.21
X180 GND.t12 CS_BIAS.t22 CS_BIAS.t23 GND.t11 sky130_fd_pr__nfet_01v8 ad=0.6303 pd=4.15 as=0.6303 ps=4.15 w=3.82 l=2.21
X181 a_n10357_8879.t6 a_n10279_8682.t25 VDD.t11 VDD.t10 sky130_fd_pr__pfet_01v8 ad=1.3065 pd=7.48 as=0.55275 ps=3.68 w=3.35 l=5.36
X182 VDD.t41 VDD.t38 VDD.t40 VDD.t39 sky130_fd_pr__pfet_01v8 ad=0.8151 pd=4.96 as=0 ps=0 w=2.09 l=2.93
X183 GND.t101 GND.t98 GND.t100 GND.t99 sky130_fd_pr__nfet_01v8 ad=0.8619 pd=5.2 as=0 ps=0 w=2.21 l=3.05
X184 a_n4238_7449.t6 a_n10279_8682.t26 VDD.t9 VDD.t8 sky130_fd_pr__pfet_01v8 ad=0.55275 pd=3.68 as=0.55275 ps=3.68 w=3.35 l=5.36
X185 GND.t97 GND.t95 VN.t0 GND.t96 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X186 GND.t91 GND.t88 GND.t90 GND.t89 sky130_fd_pr__nfet_01v8 ad=1.4898 pd=8.42 as=0 ps=0 w=3.82 l=2.21
X187 GND.t10 CS_BIAS.t81 VOUT.t80 GND.t8 sky130_fd_pr__nfet_01v8 ad=0.6303 pd=4.15 as=0.6303 ps=4.15 w=3.82 l=2.21
X188 a_n10357_8879.t5 a_n10279_8682.t27 VDD.t7 VDD.t6 sky130_fd_pr__pfet_01v8 ad=0.55275 pd=3.68 as=0.55275 ps=3.68 w=3.35 l=5.36
X189 GND.t9 CS_BIAS.t20 CS_BIAS.t21 GND.t8 sky130_fd_pr__nfet_01v8 ad=0.6303 pd=4.15 as=0.6303 ps=4.15 w=3.82 l=2.21
X190 VDD.t109 a_n16148_7944.t28 VOUT.t15 VDD.t108 sky130_fd_pr__pfet_01v8 ad=0.8151 pd=4.96 as=0.34485 ps=2.42 w=2.09 l=2.93
X191 VDD.t107 a_n16148_7944.t29 VOUT.t83 VDD.t106 sky130_fd_pr__pfet_01v8 ad=0.34485 pd=2.42 as=0.34485 ps=2.42 w=2.09 l=2.93
X192 VDD.t5 a_n10279_8682.t28 a_n10357_8879.t4 VDD.t4 sky130_fd_pr__pfet_01v8 ad=0.55275 pd=3.68 as=0.55275 ps=3.68 w=3.35 l=5.36
X193 a_n4238_7449.t1 a_n10279_8682.t29 VDD.t3 VDD.t2 sky130_fd_pr__pfet_01v8 ad=1.3065 pd=7.48 as=0.55275 ps=3.68 w=3.35 l=5.36
X194 VOUT.t21 CS_BIAS.t82 GND.t7 GND.t6 sky130_fd_pr__nfet_01v8 ad=0.6303 pd=4.15 as=1.4898 ps=8.42 w=3.82 l=2.21
X195 GND.t5 CS_BIAS.t83 VOUT.t68 GND.t4 sky130_fd_pr__nfet_01v8 ad=1.4898 pd=8.42 as=0.6303 ps=4.15 w=3.82 l=2.21
R0 CS_BIAS.n287 CS_BIAS.n243 161.3
R1 CS_BIAS.n286 CS_BIAS.n285 161.3
R2 CS_BIAS.n284 CS_BIAS.n244 161.3
R3 CS_BIAS.n283 CS_BIAS.n282 161.3
R4 CS_BIAS.n281 CS_BIAS.n245 161.3
R5 CS_BIAS.n279 CS_BIAS.n278 161.3
R6 CS_BIAS.n277 CS_BIAS.n246 161.3
R7 CS_BIAS.n276 CS_BIAS.n275 161.3
R8 CS_BIAS.n274 CS_BIAS.n247 161.3
R9 CS_BIAS.n273 CS_BIAS.n272 161.3
R10 CS_BIAS.n271 CS_BIAS.n270 161.3
R11 CS_BIAS.n269 CS_BIAS.n249 161.3
R12 CS_BIAS.n268 CS_BIAS.n267 161.3
R13 CS_BIAS.n266 CS_BIAS.n250 161.3
R14 CS_BIAS.n265 CS_BIAS.n264 161.3
R15 CS_BIAS.n262 CS_BIAS.n251 161.3
R16 CS_BIAS.n261 CS_BIAS.n260 161.3
R17 CS_BIAS.n259 CS_BIAS.n252 161.3
R18 CS_BIAS.n258 CS_BIAS.n257 161.3
R19 CS_BIAS.n256 CS_BIAS.n253 161.3
R20 CS_BIAS.n208 CS_BIAS.n205 161.3
R21 CS_BIAS.n210 CS_BIAS.n209 161.3
R22 CS_BIAS.n211 CS_BIAS.n204 161.3
R23 CS_BIAS.n213 CS_BIAS.n212 161.3
R24 CS_BIAS.n214 CS_BIAS.n203 161.3
R25 CS_BIAS.n217 CS_BIAS.n216 161.3
R26 CS_BIAS.n218 CS_BIAS.n202 161.3
R27 CS_BIAS.n220 CS_BIAS.n219 161.3
R28 CS_BIAS.n221 CS_BIAS.n201 161.3
R29 CS_BIAS.n223 CS_BIAS.n222 161.3
R30 CS_BIAS.n225 CS_BIAS.n224 161.3
R31 CS_BIAS.n226 CS_BIAS.n199 161.3
R32 CS_BIAS.n228 CS_BIAS.n227 161.3
R33 CS_BIAS.n229 CS_BIAS.n198 161.3
R34 CS_BIAS.n231 CS_BIAS.n230 161.3
R35 CS_BIAS.n233 CS_BIAS.n197 161.3
R36 CS_BIAS.n235 CS_BIAS.n234 161.3
R37 CS_BIAS.n236 CS_BIAS.n196 161.3
R38 CS_BIAS.n238 CS_BIAS.n237 161.3
R39 CS_BIAS.n239 CS_BIAS.n195 161.3
R40 CS_BIAS.n160 CS_BIAS.n157 161.3
R41 CS_BIAS.n162 CS_BIAS.n161 161.3
R42 CS_BIAS.n163 CS_BIAS.n156 161.3
R43 CS_BIAS.n165 CS_BIAS.n164 161.3
R44 CS_BIAS.n166 CS_BIAS.n155 161.3
R45 CS_BIAS.n169 CS_BIAS.n168 161.3
R46 CS_BIAS.n170 CS_BIAS.n154 161.3
R47 CS_BIAS.n172 CS_BIAS.n171 161.3
R48 CS_BIAS.n173 CS_BIAS.n153 161.3
R49 CS_BIAS.n175 CS_BIAS.n174 161.3
R50 CS_BIAS.n177 CS_BIAS.n176 161.3
R51 CS_BIAS.n178 CS_BIAS.n151 161.3
R52 CS_BIAS.n180 CS_BIAS.n179 161.3
R53 CS_BIAS.n181 CS_BIAS.n150 161.3
R54 CS_BIAS.n183 CS_BIAS.n182 161.3
R55 CS_BIAS.n185 CS_BIAS.n149 161.3
R56 CS_BIAS.n187 CS_BIAS.n186 161.3
R57 CS_BIAS.n188 CS_BIAS.n148 161.3
R58 CS_BIAS.n190 CS_BIAS.n189 161.3
R59 CS_BIAS.n191 CS_BIAS.n147 161.3
R60 CS_BIAS.n112 CS_BIAS.n109 161.3
R61 CS_BIAS.n114 CS_BIAS.n113 161.3
R62 CS_BIAS.n115 CS_BIAS.n108 161.3
R63 CS_BIAS.n117 CS_BIAS.n116 161.3
R64 CS_BIAS.n118 CS_BIAS.n107 161.3
R65 CS_BIAS.n121 CS_BIAS.n120 161.3
R66 CS_BIAS.n122 CS_BIAS.n106 161.3
R67 CS_BIAS.n124 CS_BIAS.n123 161.3
R68 CS_BIAS.n125 CS_BIAS.n105 161.3
R69 CS_BIAS.n127 CS_BIAS.n126 161.3
R70 CS_BIAS.n129 CS_BIAS.n128 161.3
R71 CS_BIAS.n130 CS_BIAS.n103 161.3
R72 CS_BIAS.n132 CS_BIAS.n131 161.3
R73 CS_BIAS.n133 CS_BIAS.n102 161.3
R74 CS_BIAS.n135 CS_BIAS.n134 161.3
R75 CS_BIAS.n137 CS_BIAS.n101 161.3
R76 CS_BIAS.n139 CS_BIAS.n138 161.3
R77 CS_BIAS.n140 CS_BIAS.n100 161.3
R78 CS_BIAS.n142 CS_BIAS.n141 161.3
R79 CS_BIAS.n143 CS_BIAS.n99 161.3
R80 CS_BIAS.n21 CS_BIAS.n18 161.3
R81 CS_BIAS.n23 CS_BIAS.n22 161.3
R82 CS_BIAS.n24 CS_BIAS.n17 161.3
R83 CS_BIAS.n26 CS_BIAS.n25 161.3
R84 CS_BIAS.n27 CS_BIAS.n16 161.3
R85 CS_BIAS.n30 CS_BIAS.n29 161.3
R86 CS_BIAS.n31 CS_BIAS.n15 161.3
R87 CS_BIAS.n33 CS_BIAS.n32 161.3
R88 CS_BIAS.n34 CS_BIAS.n14 161.3
R89 CS_BIAS.n36 CS_BIAS.n35 161.3
R90 CS_BIAS.n38 CS_BIAS.n37 161.3
R91 CS_BIAS.n39 CS_BIAS.n12 161.3
R92 CS_BIAS.n41 CS_BIAS.n40 161.3
R93 CS_BIAS.n42 CS_BIAS.n11 161.3
R94 CS_BIAS.n44 CS_BIAS.n43 161.3
R95 CS_BIAS.n46 CS_BIAS.n10 161.3
R96 CS_BIAS.n48 CS_BIAS.n47 161.3
R97 CS_BIAS.n49 CS_BIAS.n9 161.3
R98 CS_BIAS.n51 CS_BIAS.n50 161.3
R99 CS_BIAS.n52 CS_BIAS.n8 161.3
R100 CS_BIAS.n65 CS_BIAS.n62 161.3
R101 CS_BIAS.n67 CS_BIAS.n66 161.3
R102 CS_BIAS.n68 CS_BIAS.n61 161.3
R103 CS_BIAS.n70 CS_BIAS.n69 161.3
R104 CS_BIAS.n71 CS_BIAS.n60 161.3
R105 CS_BIAS.n74 CS_BIAS.n73 161.3
R106 CS_BIAS.n75 CS_BIAS.n7 161.3
R107 CS_BIAS.n77 CS_BIAS.n76 161.3
R108 CS_BIAS.n78 CS_BIAS.n6 161.3
R109 CS_BIAS.n80 CS_BIAS.n79 161.3
R110 CS_BIAS.n82 CS_BIAS.n81 161.3
R111 CS_BIAS.n83 CS_BIAS.n4 161.3
R112 CS_BIAS.n85 CS_BIAS.n84 161.3
R113 CS_BIAS.n86 CS_BIAS.n3 161.3
R114 CS_BIAS.n88 CS_BIAS.n87 161.3
R115 CS_BIAS.n90 CS_BIAS.n2 161.3
R116 CS_BIAS.n92 CS_BIAS.n91 161.3
R117 CS_BIAS.n93 CS_BIAS.n1 161.3
R118 CS_BIAS.n95 CS_BIAS.n94 161.3
R119 CS_BIAS.n96 CS_BIAS.n0 161.3
R120 CS_BIAS.n578 CS_BIAS.n534 161.3
R121 CS_BIAS.n577 CS_BIAS.n576 161.3
R122 CS_BIAS.n575 CS_BIAS.n535 161.3
R123 CS_BIAS.n574 CS_BIAS.n573 161.3
R124 CS_BIAS.n572 CS_BIAS.n536 161.3
R125 CS_BIAS.n570 CS_BIAS.n569 161.3
R126 CS_BIAS.n568 CS_BIAS.n537 161.3
R127 CS_BIAS.n567 CS_BIAS.n566 161.3
R128 CS_BIAS.n565 CS_BIAS.n538 161.3
R129 CS_BIAS.n564 CS_BIAS.n563 161.3
R130 CS_BIAS.n562 CS_BIAS.n561 161.3
R131 CS_BIAS.n560 CS_BIAS.n540 161.3
R132 CS_BIAS.n559 CS_BIAS.n558 161.3
R133 CS_BIAS.n557 CS_BIAS.n541 161.3
R134 CS_BIAS.n556 CS_BIAS.n555 161.3
R135 CS_BIAS.n553 CS_BIAS.n542 161.3
R136 CS_BIAS.n552 CS_BIAS.n551 161.3
R137 CS_BIAS.n550 CS_BIAS.n543 161.3
R138 CS_BIAS.n549 CS_BIAS.n548 161.3
R139 CS_BIAS.n547 CS_BIAS.n544 161.3
R140 CS_BIAS.n530 CS_BIAS.n486 161.3
R141 CS_BIAS.n529 CS_BIAS.n528 161.3
R142 CS_BIAS.n527 CS_BIAS.n487 161.3
R143 CS_BIAS.n526 CS_BIAS.n525 161.3
R144 CS_BIAS.n524 CS_BIAS.n488 161.3
R145 CS_BIAS.n522 CS_BIAS.n521 161.3
R146 CS_BIAS.n520 CS_BIAS.n489 161.3
R147 CS_BIAS.n519 CS_BIAS.n518 161.3
R148 CS_BIAS.n517 CS_BIAS.n490 161.3
R149 CS_BIAS.n516 CS_BIAS.n515 161.3
R150 CS_BIAS.n514 CS_BIAS.n513 161.3
R151 CS_BIAS.n512 CS_BIAS.n492 161.3
R152 CS_BIAS.n511 CS_BIAS.n510 161.3
R153 CS_BIAS.n509 CS_BIAS.n493 161.3
R154 CS_BIAS.n508 CS_BIAS.n507 161.3
R155 CS_BIAS.n505 CS_BIAS.n494 161.3
R156 CS_BIAS.n504 CS_BIAS.n503 161.3
R157 CS_BIAS.n502 CS_BIAS.n495 161.3
R158 CS_BIAS.n501 CS_BIAS.n500 161.3
R159 CS_BIAS.n499 CS_BIAS.n496 161.3
R160 CS_BIAS.n482 CS_BIAS.n438 161.3
R161 CS_BIAS.n481 CS_BIAS.n480 161.3
R162 CS_BIAS.n479 CS_BIAS.n439 161.3
R163 CS_BIAS.n478 CS_BIAS.n477 161.3
R164 CS_BIAS.n476 CS_BIAS.n440 161.3
R165 CS_BIAS.n474 CS_BIAS.n473 161.3
R166 CS_BIAS.n472 CS_BIAS.n441 161.3
R167 CS_BIAS.n471 CS_BIAS.n470 161.3
R168 CS_BIAS.n469 CS_BIAS.n442 161.3
R169 CS_BIAS.n468 CS_BIAS.n467 161.3
R170 CS_BIAS.n466 CS_BIAS.n465 161.3
R171 CS_BIAS.n464 CS_BIAS.n444 161.3
R172 CS_BIAS.n463 CS_BIAS.n462 161.3
R173 CS_BIAS.n461 CS_BIAS.n445 161.3
R174 CS_BIAS.n460 CS_BIAS.n459 161.3
R175 CS_BIAS.n457 CS_BIAS.n446 161.3
R176 CS_BIAS.n456 CS_BIAS.n455 161.3
R177 CS_BIAS.n454 CS_BIAS.n447 161.3
R178 CS_BIAS.n453 CS_BIAS.n452 161.3
R179 CS_BIAS.n451 CS_BIAS.n448 161.3
R180 CS_BIAS.n434 CS_BIAS.n390 161.3
R181 CS_BIAS.n433 CS_BIAS.n432 161.3
R182 CS_BIAS.n431 CS_BIAS.n391 161.3
R183 CS_BIAS.n430 CS_BIAS.n429 161.3
R184 CS_BIAS.n428 CS_BIAS.n392 161.3
R185 CS_BIAS.n426 CS_BIAS.n425 161.3
R186 CS_BIAS.n424 CS_BIAS.n393 161.3
R187 CS_BIAS.n423 CS_BIAS.n422 161.3
R188 CS_BIAS.n421 CS_BIAS.n394 161.3
R189 CS_BIAS.n420 CS_BIAS.n419 161.3
R190 CS_BIAS.n418 CS_BIAS.n417 161.3
R191 CS_BIAS.n416 CS_BIAS.n396 161.3
R192 CS_BIAS.n415 CS_BIAS.n414 161.3
R193 CS_BIAS.n413 CS_BIAS.n397 161.3
R194 CS_BIAS.n412 CS_BIAS.n411 161.3
R195 CS_BIAS.n409 CS_BIAS.n398 161.3
R196 CS_BIAS.n408 CS_BIAS.n407 161.3
R197 CS_BIAS.n406 CS_BIAS.n399 161.3
R198 CS_BIAS.n405 CS_BIAS.n404 161.3
R199 CS_BIAS.n403 CS_BIAS.n400 161.3
R200 CS_BIAS.n361 CS_BIAS.n317 161.3
R201 CS_BIAS.n360 CS_BIAS.n359 161.3
R202 CS_BIAS.n358 CS_BIAS.n318 161.3
R203 CS_BIAS.n357 CS_BIAS.n356 161.3
R204 CS_BIAS.n355 CS_BIAS.n319 161.3
R205 CS_BIAS.n353 CS_BIAS.n352 161.3
R206 CS_BIAS.n351 CS_BIAS.n320 161.3
R207 CS_BIAS.n350 CS_BIAS.n349 161.3
R208 CS_BIAS.n348 CS_BIAS.n321 161.3
R209 CS_BIAS.n347 CS_BIAS.n346 161.3
R210 CS_BIAS.n345 CS_BIAS.n344 161.3
R211 CS_BIAS.n343 CS_BIAS.n323 161.3
R212 CS_BIAS.n342 CS_BIAS.n341 161.3
R213 CS_BIAS.n340 CS_BIAS.n324 161.3
R214 CS_BIAS.n339 CS_BIAS.n338 161.3
R215 CS_BIAS.n336 CS_BIAS.n325 161.3
R216 CS_BIAS.n335 CS_BIAS.n334 161.3
R217 CS_BIAS.n333 CS_BIAS.n326 161.3
R218 CS_BIAS.n332 CS_BIAS.n331 161.3
R219 CS_BIAS.n330 CS_BIAS.n327 161.3
R220 CS_BIAS.n314 CS_BIAS.n298 161.3
R221 CS_BIAS.n313 CS_BIAS.n312 161.3
R222 CS_BIAS.n310 CS_BIAS.n299 161.3
R223 CS_BIAS.n309 CS_BIAS.n308 161.3
R224 CS_BIAS.n307 CS_BIAS.n300 161.3
R225 CS_BIAS.n306 CS_BIAS.n305 161.3
R226 CS_BIAS.n304 CS_BIAS.n301 161.3
R227 CS_BIAS.n368 CS_BIAS.n367 161.3
R228 CS_BIAS.n387 CS_BIAS.n291 161.3
R229 CS_BIAS.n386 CS_BIAS.n385 161.3
R230 CS_BIAS.n384 CS_BIAS.n292 161.3
R231 CS_BIAS.n383 CS_BIAS.n382 161.3
R232 CS_BIAS.n381 CS_BIAS.n293 161.3
R233 CS_BIAS.n379 CS_BIAS.n378 161.3
R234 CS_BIAS.n377 CS_BIAS.n294 161.3
R235 CS_BIAS.n376 CS_BIAS.n375 161.3
R236 CS_BIAS.n374 CS_BIAS.n295 161.3
R237 CS_BIAS.n373 CS_BIAS.n372 161.3
R238 CS_BIAS.n371 CS_BIAS.n370 161.3
R239 CS_BIAS.n369 CS_BIAS.n297 161.3
R240 CS_BIAS.n289 CS_BIAS.n288 93.694
R241 CS_BIAS.n241 CS_BIAS.n240 93.694
R242 CS_BIAS.n193 CS_BIAS.n192 93.694
R243 CS_BIAS.n145 CS_BIAS.n144 93.694
R244 CS_BIAS.n54 CS_BIAS.n53 93.694
R245 CS_BIAS.n98 CS_BIAS.n97 93.694
R246 CS_BIAS.n580 CS_BIAS.n579 93.694
R247 CS_BIAS.n532 CS_BIAS.n531 93.694
R248 CS_BIAS.n484 CS_BIAS.n483 93.694
R249 CS_BIAS.n436 CS_BIAS.n435 93.694
R250 CS_BIAS.n363 CS_BIAS.n362 93.694
R251 CS_BIAS.n389 CS_BIAS.n388 93.694
R252 CS_BIAS.n59 CS_BIAS.n58 75.2357
R253 CS_BIAS.n366 CS_BIAS.n315 75.2357
R254 CS_BIAS.n254 CS_BIAS.t82 75.1476
R255 CS_BIAS.n545 CS_BIAS.t27 75.1476
R256 CS_BIAS.n497 CS_BIAS.t63 75.1476
R257 CS_BIAS.n449 CS_BIAS.t52 75.1476
R258 CS_BIAS.n401 CS_BIAS.t44 75.1476
R259 CS_BIAS.n328 CS_BIAS.t18 75.1476
R260 CS_BIAS.n302 CS_BIAS.t24 75.1476
R261 CS_BIAS.n206 CS_BIAS.t56 75.1476
R262 CS_BIAS.n158 CS_BIAS.t49 75.1476
R263 CS_BIAS.n110 CS_BIAS.t73 75.1476
R264 CS_BIAS.n19 CS_BIAS.t4 75.1476
R265 CS_BIAS.n63 CS_BIAS.t51 75.1476
R266 CS_BIAS.n59 CS_BIAS.n57 73.0762
R267 CS_BIAS.n56 CS_BIAS.n55 73.0762
R268 CS_BIAS.n366 CS_BIAS.n316 73.0762
R269 CS_BIAS.n365 CS_BIAS.n364 73.0762
R270 CS_BIAS.n207 CS_BIAS.n206 56.163
R271 CS_BIAS.n159 CS_BIAS.n158 56.163
R272 CS_BIAS.n111 CS_BIAS.n110 56.163
R273 CS_BIAS.n20 CS_BIAS.n19 56.163
R274 CS_BIAS.n64 CS_BIAS.n63 56.163
R275 CS_BIAS.n255 CS_BIAS.n254 56.163
R276 CS_BIAS.n546 CS_BIAS.n545 56.163
R277 CS_BIAS.n498 CS_BIAS.n497 56.163
R278 CS_BIAS.n450 CS_BIAS.n449 56.163
R279 CS_BIAS.n402 CS_BIAS.n401 56.163
R280 CS_BIAS.n329 CS_BIAS.n328 56.163
R281 CS_BIAS.n303 CS_BIAS.n302 56.163
R282 CS_BIAS.n286 CS_BIAS.n244 48.3272
R283 CS_BIAS.n238 CS_BIAS.n196 48.3272
R284 CS_BIAS.n190 CS_BIAS.n148 48.3272
R285 CS_BIAS.n142 CS_BIAS.n100 48.3272
R286 CS_BIAS.n51 CS_BIAS.n9 48.3272
R287 CS_BIAS.n95 CS_BIAS.n1 48.3272
R288 CS_BIAS.n577 CS_BIAS.n535 48.3272
R289 CS_BIAS.n529 CS_BIAS.n487 48.3272
R290 CS_BIAS.n481 CS_BIAS.n439 48.3272
R291 CS_BIAS.n433 CS_BIAS.n391 48.3272
R292 CS_BIAS.n360 CS_BIAS.n318 48.3272
R293 CS_BIAS.n386 CS_BIAS.n292 48.3272
R294 CS_BIAS.n257 CS_BIAS.n252 44.4521
R295 CS_BIAS.n275 CS_BIAS.n246 44.4521
R296 CS_BIAS.n227 CS_BIAS.n198 44.4521
R297 CS_BIAS.n209 CS_BIAS.n204 44.4521
R298 CS_BIAS.n179 CS_BIAS.n150 44.4521
R299 CS_BIAS.n161 CS_BIAS.n156 44.4521
R300 CS_BIAS.n131 CS_BIAS.n102 44.4521
R301 CS_BIAS.n113 CS_BIAS.n108 44.4521
R302 CS_BIAS.n40 CS_BIAS.n11 44.4521
R303 CS_BIAS.n22 CS_BIAS.n17 44.4521
R304 CS_BIAS.n84 CS_BIAS.n3 44.4521
R305 CS_BIAS.n66 CS_BIAS.n61 44.4521
R306 CS_BIAS.n548 CS_BIAS.n543 44.4521
R307 CS_BIAS.n566 CS_BIAS.n537 44.4521
R308 CS_BIAS.n500 CS_BIAS.n495 44.4521
R309 CS_BIAS.n518 CS_BIAS.n489 44.4521
R310 CS_BIAS.n452 CS_BIAS.n447 44.4521
R311 CS_BIAS.n470 CS_BIAS.n441 44.4521
R312 CS_BIAS.n404 CS_BIAS.n399 44.4521
R313 CS_BIAS.n422 CS_BIAS.n393 44.4521
R314 CS_BIAS.n331 CS_BIAS.n326 44.4521
R315 CS_BIAS.n349 CS_BIAS.n320 44.4521
R316 CS_BIAS.n375 CS_BIAS.n294 44.4521
R317 CS_BIAS.n305 CS_BIAS.n300 44.4521
R318 CS_BIAS.n255 CS_BIAS.t66 41.6575
R319 CS_BIAS.n263 CS_BIAS.t67 41.6575
R320 CS_BIAS.n248 CS_BIAS.t60 41.6575
R321 CS_BIAS.n280 CS_BIAS.t61 41.6575
R322 CS_BIAS.n288 CS_BIAS.t40 41.6575
R323 CS_BIAS.n240 CS_BIAS.t78 41.6575
R324 CS_BIAS.n232 CS_BIAS.t30 41.6575
R325 CS_BIAS.n200 CS_BIAS.t31 41.6575
R326 CS_BIAS.n215 CS_BIAS.t35 41.6575
R327 CS_BIAS.n207 CS_BIAS.t33 41.6575
R328 CS_BIAS.n192 CS_BIAS.t45 41.6575
R329 CS_BIAS.n184 CS_BIAS.t57 41.6575
R330 CS_BIAS.n152 CS_BIAS.t55 41.6575
R331 CS_BIAS.n167 CS_BIAS.t34 41.6575
R332 CS_BIAS.n159 CS_BIAS.t32 41.6575
R333 CS_BIAS.n144 CS_BIAS.t43 41.6575
R334 CS_BIAS.n136 CS_BIAS.t26 41.6575
R335 CS_BIAS.n104 CS_BIAS.t81 41.6575
R336 CS_BIAS.n119 CS_BIAS.t25 41.6575
R337 CS_BIAS.n111 CS_BIAS.t80 41.6575
R338 CS_BIAS.n53 CS_BIAS.t16 41.6575
R339 CS_BIAS.n45 CS_BIAS.t0 41.6575
R340 CS_BIAS.n13 CS_BIAS.t20 41.6575
R341 CS_BIAS.n28 CS_BIAS.t2 41.6575
R342 CS_BIAS.n20 CS_BIAS.t22 41.6575
R343 CS_BIAS.n97 CS_BIAS.t83 41.6575
R344 CS_BIAS.n89 CS_BIAS.t79 41.6575
R345 CS_BIAS.n5 CS_BIAS.t71 41.6575
R346 CS_BIAS.n72 CS_BIAS.t74 41.6575
R347 CS_BIAS.n64 CS_BIAS.t65 41.6575
R348 CS_BIAS.n546 CS_BIAS.t28 41.6575
R349 CS_BIAS.n554 CS_BIAS.t76 41.6575
R350 CS_BIAS.n539 CS_BIAS.t75 41.6575
R351 CS_BIAS.n571 CS_BIAS.t70 41.6575
R352 CS_BIAS.n579 CS_BIAS.t69 41.6575
R353 CS_BIAS.n498 CS_BIAS.t64 41.6575
R354 CS_BIAS.n506 CS_BIAS.t41 41.6575
R355 CS_BIAS.n491 CS_BIAS.t42 41.6575
R356 CS_BIAS.n523 CS_BIAS.t36 41.6575
R357 CS_BIAS.n531 CS_BIAS.t38 41.6575
R358 CS_BIAS.n450 CS_BIAS.t53 41.6575
R359 CS_BIAS.n458 CS_BIAS.t37 41.6575
R360 CS_BIAS.n443 CS_BIAS.t39 41.6575
R361 CS_BIAS.n475 CS_BIAS.t58 41.6575
R362 CS_BIAS.n483 CS_BIAS.t59 41.6575
R363 CS_BIAS.n402 CS_BIAS.t48 41.6575
R364 CS_BIAS.n410 CS_BIAS.t62 41.6575
R365 CS_BIAS.n395 CS_BIAS.t72 41.6575
R366 CS_BIAS.n427 CS_BIAS.t68 41.6575
R367 CS_BIAS.n435 CS_BIAS.t77 41.6575
R368 CS_BIAS.n329 CS_BIAS.t14 41.6575
R369 CS_BIAS.n337 CS_BIAS.t10 41.6575
R370 CS_BIAS.n322 CS_BIAS.t6 41.6575
R371 CS_BIAS.n354 CS_BIAS.t12 41.6575
R372 CS_BIAS.n362 CS_BIAS.t8 41.6575
R373 CS_BIAS.n388 CS_BIAS.t54 41.6575
R374 CS_BIAS.n380 CS_BIAS.t47 41.6575
R375 CS_BIAS.n296 CS_BIAS.t50 41.6575
R376 CS_BIAS.n303 CS_BIAS.t29 41.6575
R377 CS_BIAS.n311 CS_BIAS.t46 41.6575
R378 CS_BIAS.n268 CS_BIAS.n250 40.577
R379 CS_BIAS.n269 CS_BIAS.n268 40.577
R380 CS_BIAS.n221 CS_BIAS.n220 40.577
R381 CS_BIAS.n220 CS_BIAS.n202 40.577
R382 CS_BIAS.n173 CS_BIAS.n172 40.577
R383 CS_BIAS.n172 CS_BIAS.n154 40.577
R384 CS_BIAS.n125 CS_BIAS.n124 40.577
R385 CS_BIAS.n124 CS_BIAS.n106 40.577
R386 CS_BIAS.n34 CS_BIAS.n33 40.577
R387 CS_BIAS.n33 CS_BIAS.n15 40.577
R388 CS_BIAS.n78 CS_BIAS.n77 40.577
R389 CS_BIAS.n77 CS_BIAS.n7 40.577
R390 CS_BIAS.n559 CS_BIAS.n541 40.577
R391 CS_BIAS.n560 CS_BIAS.n559 40.577
R392 CS_BIAS.n511 CS_BIAS.n493 40.577
R393 CS_BIAS.n512 CS_BIAS.n511 40.577
R394 CS_BIAS.n463 CS_BIAS.n445 40.577
R395 CS_BIAS.n464 CS_BIAS.n463 40.577
R396 CS_BIAS.n415 CS_BIAS.n397 40.577
R397 CS_BIAS.n416 CS_BIAS.n415 40.577
R398 CS_BIAS.n342 CS_BIAS.n324 40.577
R399 CS_BIAS.n343 CS_BIAS.n342 40.577
R400 CS_BIAS.n369 CS_BIAS.n368 40.577
R401 CS_BIAS.n368 CS_BIAS.n298 40.577
R402 CS_BIAS.n261 CS_BIAS.n252 36.702
R403 CS_BIAS.n275 CS_BIAS.n274 36.702
R404 CS_BIAS.n227 CS_BIAS.n226 36.702
R405 CS_BIAS.n213 CS_BIAS.n204 36.702
R406 CS_BIAS.n179 CS_BIAS.n178 36.702
R407 CS_BIAS.n165 CS_BIAS.n156 36.702
R408 CS_BIAS.n131 CS_BIAS.n130 36.702
R409 CS_BIAS.n117 CS_BIAS.n108 36.702
R410 CS_BIAS.n40 CS_BIAS.n39 36.702
R411 CS_BIAS.n26 CS_BIAS.n17 36.702
R412 CS_BIAS.n84 CS_BIAS.n83 36.702
R413 CS_BIAS.n70 CS_BIAS.n61 36.702
R414 CS_BIAS.n552 CS_BIAS.n543 36.702
R415 CS_BIAS.n566 CS_BIAS.n565 36.702
R416 CS_BIAS.n504 CS_BIAS.n495 36.702
R417 CS_BIAS.n518 CS_BIAS.n517 36.702
R418 CS_BIAS.n456 CS_BIAS.n447 36.702
R419 CS_BIAS.n470 CS_BIAS.n469 36.702
R420 CS_BIAS.n408 CS_BIAS.n399 36.702
R421 CS_BIAS.n422 CS_BIAS.n421 36.702
R422 CS_BIAS.n335 CS_BIAS.n326 36.702
R423 CS_BIAS.n349 CS_BIAS.n348 36.702
R424 CS_BIAS.n375 CS_BIAS.n374 36.702
R425 CS_BIAS.n309 CS_BIAS.n300 36.702
R426 CS_BIAS.n282 CS_BIAS.n244 32.8269
R427 CS_BIAS.n234 CS_BIAS.n196 32.8269
R428 CS_BIAS.n186 CS_BIAS.n148 32.8269
R429 CS_BIAS.n138 CS_BIAS.n100 32.8269
R430 CS_BIAS.n47 CS_BIAS.n9 32.8269
R431 CS_BIAS.n91 CS_BIAS.n1 32.8269
R432 CS_BIAS.n573 CS_BIAS.n535 32.8269
R433 CS_BIAS.n525 CS_BIAS.n487 32.8269
R434 CS_BIAS.n477 CS_BIAS.n439 32.8269
R435 CS_BIAS.n429 CS_BIAS.n391 32.8269
R436 CS_BIAS.n356 CS_BIAS.n318 32.8269
R437 CS_BIAS.n382 CS_BIAS.n292 32.8269
R438 CS_BIAS.n257 CS_BIAS.n256 24.5923
R439 CS_BIAS.n264 CS_BIAS.n250 24.5923
R440 CS_BIAS.n262 CS_BIAS.n261 24.5923
R441 CS_BIAS.n274 CS_BIAS.n273 24.5923
R442 CS_BIAS.n270 CS_BIAS.n269 24.5923
R443 CS_BIAS.n282 CS_BIAS.n281 24.5923
R444 CS_BIAS.n279 CS_BIAS.n246 24.5923
R445 CS_BIAS.n287 CS_BIAS.n286 24.5923
R446 CS_BIAS.n239 CS_BIAS.n238 24.5923
R447 CS_BIAS.n234 CS_BIAS.n233 24.5923
R448 CS_BIAS.n231 CS_BIAS.n198 24.5923
R449 CS_BIAS.n226 CS_BIAS.n225 24.5923
R450 CS_BIAS.n222 CS_BIAS.n221 24.5923
R451 CS_BIAS.n216 CS_BIAS.n202 24.5923
R452 CS_BIAS.n214 CS_BIAS.n213 24.5923
R453 CS_BIAS.n209 CS_BIAS.n208 24.5923
R454 CS_BIAS.n191 CS_BIAS.n190 24.5923
R455 CS_BIAS.n186 CS_BIAS.n185 24.5923
R456 CS_BIAS.n183 CS_BIAS.n150 24.5923
R457 CS_BIAS.n178 CS_BIAS.n177 24.5923
R458 CS_BIAS.n174 CS_BIAS.n173 24.5923
R459 CS_BIAS.n168 CS_BIAS.n154 24.5923
R460 CS_BIAS.n166 CS_BIAS.n165 24.5923
R461 CS_BIAS.n161 CS_BIAS.n160 24.5923
R462 CS_BIAS.n143 CS_BIAS.n142 24.5923
R463 CS_BIAS.n138 CS_BIAS.n137 24.5923
R464 CS_BIAS.n135 CS_BIAS.n102 24.5923
R465 CS_BIAS.n130 CS_BIAS.n129 24.5923
R466 CS_BIAS.n126 CS_BIAS.n125 24.5923
R467 CS_BIAS.n120 CS_BIAS.n106 24.5923
R468 CS_BIAS.n118 CS_BIAS.n117 24.5923
R469 CS_BIAS.n113 CS_BIAS.n112 24.5923
R470 CS_BIAS.n52 CS_BIAS.n51 24.5923
R471 CS_BIAS.n47 CS_BIAS.n46 24.5923
R472 CS_BIAS.n44 CS_BIAS.n11 24.5923
R473 CS_BIAS.n39 CS_BIAS.n38 24.5923
R474 CS_BIAS.n35 CS_BIAS.n34 24.5923
R475 CS_BIAS.n29 CS_BIAS.n15 24.5923
R476 CS_BIAS.n27 CS_BIAS.n26 24.5923
R477 CS_BIAS.n22 CS_BIAS.n21 24.5923
R478 CS_BIAS.n96 CS_BIAS.n95 24.5923
R479 CS_BIAS.n91 CS_BIAS.n90 24.5923
R480 CS_BIAS.n88 CS_BIAS.n3 24.5923
R481 CS_BIAS.n83 CS_BIAS.n82 24.5923
R482 CS_BIAS.n79 CS_BIAS.n78 24.5923
R483 CS_BIAS.n73 CS_BIAS.n7 24.5923
R484 CS_BIAS.n71 CS_BIAS.n70 24.5923
R485 CS_BIAS.n66 CS_BIAS.n65 24.5923
R486 CS_BIAS.n548 CS_BIAS.n547 24.5923
R487 CS_BIAS.n553 CS_BIAS.n552 24.5923
R488 CS_BIAS.n555 CS_BIAS.n541 24.5923
R489 CS_BIAS.n561 CS_BIAS.n560 24.5923
R490 CS_BIAS.n565 CS_BIAS.n564 24.5923
R491 CS_BIAS.n570 CS_BIAS.n537 24.5923
R492 CS_BIAS.n573 CS_BIAS.n572 24.5923
R493 CS_BIAS.n578 CS_BIAS.n577 24.5923
R494 CS_BIAS.n500 CS_BIAS.n499 24.5923
R495 CS_BIAS.n505 CS_BIAS.n504 24.5923
R496 CS_BIAS.n507 CS_BIAS.n493 24.5923
R497 CS_BIAS.n513 CS_BIAS.n512 24.5923
R498 CS_BIAS.n517 CS_BIAS.n516 24.5923
R499 CS_BIAS.n522 CS_BIAS.n489 24.5923
R500 CS_BIAS.n525 CS_BIAS.n524 24.5923
R501 CS_BIAS.n530 CS_BIAS.n529 24.5923
R502 CS_BIAS.n452 CS_BIAS.n451 24.5923
R503 CS_BIAS.n457 CS_BIAS.n456 24.5923
R504 CS_BIAS.n459 CS_BIAS.n445 24.5923
R505 CS_BIAS.n465 CS_BIAS.n464 24.5923
R506 CS_BIAS.n469 CS_BIAS.n468 24.5923
R507 CS_BIAS.n474 CS_BIAS.n441 24.5923
R508 CS_BIAS.n477 CS_BIAS.n476 24.5923
R509 CS_BIAS.n482 CS_BIAS.n481 24.5923
R510 CS_BIAS.n404 CS_BIAS.n403 24.5923
R511 CS_BIAS.n409 CS_BIAS.n408 24.5923
R512 CS_BIAS.n411 CS_BIAS.n397 24.5923
R513 CS_BIAS.n417 CS_BIAS.n416 24.5923
R514 CS_BIAS.n421 CS_BIAS.n420 24.5923
R515 CS_BIAS.n426 CS_BIAS.n393 24.5923
R516 CS_BIAS.n429 CS_BIAS.n428 24.5923
R517 CS_BIAS.n434 CS_BIAS.n433 24.5923
R518 CS_BIAS.n331 CS_BIAS.n330 24.5923
R519 CS_BIAS.n336 CS_BIAS.n335 24.5923
R520 CS_BIAS.n338 CS_BIAS.n324 24.5923
R521 CS_BIAS.n344 CS_BIAS.n343 24.5923
R522 CS_BIAS.n348 CS_BIAS.n347 24.5923
R523 CS_BIAS.n353 CS_BIAS.n320 24.5923
R524 CS_BIAS.n356 CS_BIAS.n355 24.5923
R525 CS_BIAS.n361 CS_BIAS.n360 24.5923
R526 CS_BIAS.n387 CS_BIAS.n386 24.5923
R527 CS_BIAS.n379 CS_BIAS.n294 24.5923
R528 CS_BIAS.n382 CS_BIAS.n381 24.5923
R529 CS_BIAS.n370 CS_BIAS.n369 24.5923
R530 CS_BIAS.n374 CS_BIAS.n373 24.5923
R531 CS_BIAS.n305 CS_BIAS.n304 24.5923
R532 CS_BIAS.n310 CS_BIAS.n309 24.5923
R533 CS_BIAS.n312 CS_BIAS.n298 24.5923
R534 CS_BIAS.n288 CS_BIAS.n287 17.2148
R535 CS_BIAS.n240 CS_BIAS.n239 17.2148
R536 CS_BIAS.n192 CS_BIAS.n191 17.2148
R537 CS_BIAS.n144 CS_BIAS.n143 17.2148
R538 CS_BIAS.n53 CS_BIAS.n52 17.2148
R539 CS_BIAS.n97 CS_BIAS.n96 17.2148
R540 CS_BIAS.n579 CS_BIAS.n578 17.2148
R541 CS_BIAS.n531 CS_BIAS.n530 17.2148
R542 CS_BIAS.n483 CS_BIAS.n482 17.2148
R543 CS_BIAS.n435 CS_BIAS.n434 17.2148
R544 CS_BIAS.n362 CS_BIAS.n361 17.2148
R545 CS_BIAS.n388 CS_BIAS.n387 17.2148
R546 CS_BIAS.n256 CS_BIAS.n255 15.2474
R547 CS_BIAS.n280 CS_BIAS.n279 15.2474
R548 CS_BIAS.n232 CS_BIAS.n231 15.2474
R549 CS_BIAS.n208 CS_BIAS.n207 15.2474
R550 CS_BIAS.n184 CS_BIAS.n183 15.2474
R551 CS_BIAS.n160 CS_BIAS.n159 15.2474
R552 CS_BIAS.n136 CS_BIAS.n135 15.2474
R553 CS_BIAS.n112 CS_BIAS.n111 15.2474
R554 CS_BIAS.n45 CS_BIAS.n44 15.2474
R555 CS_BIAS.n21 CS_BIAS.n20 15.2474
R556 CS_BIAS.n89 CS_BIAS.n88 15.2474
R557 CS_BIAS.n65 CS_BIAS.n64 15.2474
R558 CS_BIAS.n547 CS_BIAS.n546 15.2474
R559 CS_BIAS.n571 CS_BIAS.n570 15.2474
R560 CS_BIAS.n499 CS_BIAS.n498 15.2474
R561 CS_BIAS.n523 CS_BIAS.n522 15.2474
R562 CS_BIAS.n451 CS_BIAS.n450 15.2474
R563 CS_BIAS.n475 CS_BIAS.n474 15.2474
R564 CS_BIAS.n403 CS_BIAS.n402 15.2474
R565 CS_BIAS.n427 CS_BIAS.n426 15.2474
R566 CS_BIAS.n330 CS_BIAS.n329 15.2474
R567 CS_BIAS.n354 CS_BIAS.n353 15.2474
R568 CS_BIAS.n380 CS_BIAS.n379 15.2474
R569 CS_BIAS.n304 CS_BIAS.n303 15.2474
R570 CS_BIAS.n264 CS_BIAS.n263 13.2801
R571 CS_BIAS.n270 CS_BIAS.n248 13.2801
R572 CS_BIAS.n222 CS_BIAS.n200 13.2801
R573 CS_BIAS.n216 CS_BIAS.n215 13.2801
R574 CS_BIAS.n174 CS_BIAS.n152 13.2801
R575 CS_BIAS.n168 CS_BIAS.n167 13.2801
R576 CS_BIAS.n126 CS_BIAS.n104 13.2801
R577 CS_BIAS.n120 CS_BIAS.n119 13.2801
R578 CS_BIAS.n35 CS_BIAS.n13 13.2801
R579 CS_BIAS.n29 CS_BIAS.n28 13.2801
R580 CS_BIAS.n79 CS_BIAS.n5 13.2801
R581 CS_BIAS.n73 CS_BIAS.n72 13.2801
R582 CS_BIAS.n555 CS_BIAS.n554 13.2801
R583 CS_BIAS.n561 CS_BIAS.n539 13.2801
R584 CS_BIAS.n507 CS_BIAS.n506 13.2801
R585 CS_BIAS.n513 CS_BIAS.n491 13.2801
R586 CS_BIAS.n459 CS_BIAS.n458 13.2801
R587 CS_BIAS.n465 CS_BIAS.n443 13.2801
R588 CS_BIAS.n411 CS_BIAS.n410 13.2801
R589 CS_BIAS.n417 CS_BIAS.n395 13.2801
R590 CS_BIAS.n338 CS_BIAS.n337 13.2801
R591 CS_BIAS.n344 CS_BIAS.n322 13.2801
R592 CS_BIAS.n370 CS_BIAS.n296 13.2801
R593 CS_BIAS.n312 CS_BIAS.n311 13.2801
R594 CS_BIAS.n56 CS_BIAS.n54 13.0109
R595 CS_BIAS.n365 CS_BIAS.n363 13.0109
R596 CS_BIAS.n263 CS_BIAS.n262 11.3127
R597 CS_BIAS.n273 CS_BIAS.n248 11.3127
R598 CS_BIAS.n225 CS_BIAS.n200 11.3127
R599 CS_BIAS.n215 CS_BIAS.n214 11.3127
R600 CS_BIAS.n177 CS_BIAS.n152 11.3127
R601 CS_BIAS.n167 CS_BIAS.n166 11.3127
R602 CS_BIAS.n129 CS_BIAS.n104 11.3127
R603 CS_BIAS.n119 CS_BIAS.n118 11.3127
R604 CS_BIAS.n38 CS_BIAS.n13 11.3127
R605 CS_BIAS.n28 CS_BIAS.n27 11.3127
R606 CS_BIAS.n82 CS_BIAS.n5 11.3127
R607 CS_BIAS.n72 CS_BIAS.n71 11.3127
R608 CS_BIAS.n554 CS_BIAS.n553 11.3127
R609 CS_BIAS.n564 CS_BIAS.n539 11.3127
R610 CS_BIAS.n506 CS_BIAS.n505 11.3127
R611 CS_BIAS.n516 CS_BIAS.n491 11.3127
R612 CS_BIAS.n458 CS_BIAS.n457 11.3127
R613 CS_BIAS.n468 CS_BIAS.n443 11.3127
R614 CS_BIAS.n410 CS_BIAS.n409 11.3127
R615 CS_BIAS.n420 CS_BIAS.n395 11.3127
R616 CS_BIAS.n337 CS_BIAS.n336 11.3127
R617 CS_BIAS.n347 CS_BIAS.n322 11.3127
R618 CS_BIAS.n373 CS_BIAS.n296 11.3127
R619 CS_BIAS.n311 CS_BIAS.n310 11.3127
R620 CS_BIAS.n76 CS_BIAS.n59 9.50363
R621 CS_BIAS.n367 CS_BIAS.n366 9.50363
R622 CS_BIAS.n281 CS_BIAS.n280 9.3454
R623 CS_BIAS.n233 CS_BIAS.n232 9.3454
R624 CS_BIAS.n185 CS_BIAS.n184 9.3454
R625 CS_BIAS.n137 CS_BIAS.n136 9.3454
R626 CS_BIAS.n46 CS_BIAS.n45 9.3454
R627 CS_BIAS.n90 CS_BIAS.n89 9.3454
R628 CS_BIAS.n572 CS_BIAS.n571 9.3454
R629 CS_BIAS.n524 CS_BIAS.n523 9.3454
R630 CS_BIAS.n476 CS_BIAS.n475 9.3454
R631 CS_BIAS.n428 CS_BIAS.n427 9.3454
R632 CS_BIAS.n355 CS_BIAS.n354 9.3454
R633 CS_BIAS.n381 CS_BIAS.n380 9.3454
R634 CS_BIAS.n254 CS_BIAS.n253 9.22054
R635 CS_BIAS.n206 CS_BIAS.n205 9.22054
R636 CS_BIAS.n158 CS_BIAS.n157 9.22054
R637 CS_BIAS.n110 CS_BIAS.n109 9.22054
R638 CS_BIAS.n19 CS_BIAS.n18 9.22054
R639 CS_BIAS.n63 CS_BIAS.n62 9.22054
R640 CS_BIAS.n545 CS_BIAS.n544 9.22054
R641 CS_BIAS.n497 CS_BIAS.n496 9.22054
R642 CS_BIAS.n449 CS_BIAS.n448 9.22054
R643 CS_BIAS.n401 CS_BIAS.n400 9.22054
R644 CS_BIAS.n328 CS_BIAS.n327 9.22054
R645 CS_BIAS.n302 CS_BIAS.n301 9.22054
R646 CS_BIAS.n582 CS_BIAS.n290 7.6798
R647 CS_BIAS.n146 CS_BIAS.n98 7.33152
R648 CS_BIAS.n437 CS_BIAS.n389 7.33152
R649 CS_BIAS.n582 CS_BIAS.n581 6.40861
R650 CS_BIAS CS_BIAS.n582 5.24691
R651 CS_BIAS.n57 CS_BIAS.t21 5.18375
R652 CS_BIAS.n57 CS_BIAS.t3 5.18375
R653 CS_BIAS.n58 CS_BIAS.t23 5.18375
R654 CS_BIAS.n58 CS_BIAS.t5 5.18375
R655 CS_BIAS.n55 CS_BIAS.t17 5.18375
R656 CS_BIAS.n55 CS_BIAS.t1 5.18375
R657 CS_BIAS.n316 CS_BIAS.t11 5.18375
R658 CS_BIAS.n316 CS_BIAS.t7 5.18375
R659 CS_BIAS.n364 CS_BIAS.t13 5.18375
R660 CS_BIAS.n364 CS_BIAS.t9 5.18375
R661 CS_BIAS.n315 CS_BIAS.t19 5.18375
R662 CS_BIAS.n315 CS_BIAS.t15 5.18375
R663 CS_BIAS.n290 CS_BIAS.n289 5.06447
R664 CS_BIAS.n242 CS_BIAS.n241 5.06447
R665 CS_BIAS.n194 CS_BIAS.n193 5.06447
R666 CS_BIAS.n146 CS_BIAS.n145 5.06447
R667 CS_BIAS.n581 CS_BIAS.n580 5.06447
R668 CS_BIAS.n533 CS_BIAS.n532 5.06447
R669 CS_BIAS.n485 CS_BIAS.n484 5.06447
R670 CS_BIAS.n437 CS_BIAS.n436 5.06447
R671 CS_BIAS.n194 CS_BIAS.n146 2.26755
R672 CS_BIAS.n242 CS_BIAS.n194 2.26755
R673 CS_BIAS.n290 CS_BIAS.n242 2.26755
R674 CS_BIAS.n485 CS_BIAS.n437 2.26755
R675 CS_BIAS.n533 CS_BIAS.n485 2.26755
R676 CS_BIAS.n581 CS_BIAS.n533 2.26755
R677 CS_BIAS.n59 CS_BIAS.n56 2.15998
R678 CS_BIAS.n366 CS_BIAS.n365 2.15998
R679 CS_BIAS.n289 CS_BIAS.n243 0.278335
R680 CS_BIAS.n241 CS_BIAS.n195 0.278335
R681 CS_BIAS.n193 CS_BIAS.n147 0.278335
R682 CS_BIAS.n145 CS_BIAS.n99 0.278335
R683 CS_BIAS.n54 CS_BIAS.n8 0.278335
R684 CS_BIAS.n98 CS_BIAS.n0 0.278335
R685 CS_BIAS.n580 CS_BIAS.n534 0.278335
R686 CS_BIAS.n532 CS_BIAS.n486 0.278335
R687 CS_BIAS.n484 CS_BIAS.n438 0.278335
R688 CS_BIAS.n436 CS_BIAS.n390 0.278335
R689 CS_BIAS.n363 CS_BIAS.n317 0.278335
R690 CS_BIAS.n389 CS_BIAS.n291 0.278335
R691 CS_BIAS.n285 CS_BIAS.n243 0.189894
R692 CS_BIAS.n285 CS_BIAS.n284 0.189894
R693 CS_BIAS.n284 CS_BIAS.n283 0.189894
R694 CS_BIAS.n283 CS_BIAS.n245 0.189894
R695 CS_BIAS.n278 CS_BIAS.n245 0.189894
R696 CS_BIAS.n278 CS_BIAS.n277 0.189894
R697 CS_BIAS.n277 CS_BIAS.n276 0.189894
R698 CS_BIAS.n276 CS_BIAS.n247 0.189894
R699 CS_BIAS.n272 CS_BIAS.n247 0.189894
R700 CS_BIAS.n272 CS_BIAS.n271 0.189894
R701 CS_BIAS.n271 CS_BIAS.n249 0.189894
R702 CS_BIAS.n267 CS_BIAS.n249 0.189894
R703 CS_BIAS.n267 CS_BIAS.n266 0.189894
R704 CS_BIAS.n266 CS_BIAS.n265 0.189894
R705 CS_BIAS.n265 CS_BIAS.n251 0.189894
R706 CS_BIAS.n260 CS_BIAS.n251 0.189894
R707 CS_BIAS.n260 CS_BIAS.n259 0.189894
R708 CS_BIAS.n259 CS_BIAS.n258 0.189894
R709 CS_BIAS.n258 CS_BIAS.n253 0.189894
R710 CS_BIAS.n237 CS_BIAS.n195 0.189894
R711 CS_BIAS.n237 CS_BIAS.n236 0.189894
R712 CS_BIAS.n236 CS_BIAS.n235 0.189894
R713 CS_BIAS.n235 CS_BIAS.n197 0.189894
R714 CS_BIAS.n230 CS_BIAS.n197 0.189894
R715 CS_BIAS.n230 CS_BIAS.n229 0.189894
R716 CS_BIAS.n229 CS_BIAS.n228 0.189894
R717 CS_BIAS.n228 CS_BIAS.n199 0.189894
R718 CS_BIAS.n224 CS_BIAS.n199 0.189894
R719 CS_BIAS.n224 CS_BIAS.n223 0.189894
R720 CS_BIAS.n223 CS_BIAS.n201 0.189894
R721 CS_BIAS.n219 CS_BIAS.n201 0.189894
R722 CS_BIAS.n219 CS_BIAS.n218 0.189894
R723 CS_BIAS.n218 CS_BIAS.n217 0.189894
R724 CS_BIAS.n217 CS_BIAS.n203 0.189894
R725 CS_BIAS.n212 CS_BIAS.n203 0.189894
R726 CS_BIAS.n212 CS_BIAS.n211 0.189894
R727 CS_BIAS.n211 CS_BIAS.n210 0.189894
R728 CS_BIAS.n210 CS_BIAS.n205 0.189894
R729 CS_BIAS.n189 CS_BIAS.n147 0.189894
R730 CS_BIAS.n189 CS_BIAS.n188 0.189894
R731 CS_BIAS.n188 CS_BIAS.n187 0.189894
R732 CS_BIAS.n187 CS_BIAS.n149 0.189894
R733 CS_BIAS.n182 CS_BIAS.n149 0.189894
R734 CS_BIAS.n182 CS_BIAS.n181 0.189894
R735 CS_BIAS.n181 CS_BIAS.n180 0.189894
R736 CS_BIAS.n180 CS_BIAS.n151 0.189894
R737 CS_BIAS.n176 CS_BIAS.n151 0.189894
R738 CS_BIAS.n176 CS_BIAS.n175 0.189894
R739 CS_BIAS.n175 CS_BIAS.n153 0.189894
R740 CS_BIAS.n171 CS_BIAS.n153 0.189894
R741 CS_BIAS.n171 CS_BIAS.n170 0.189894
R742 CS_BIAS.n170 CS_BIAS.n169 0.189894
R743 CS_BIAS.n169 CS_BIAS.n155 0.189894
R744 CS_BIAS.n164 CS_BIAS.n155 0.189894
R745 CS_BIAS.n164 CS_BIAS.n163 0.189894
R746 CS_BIAS.n163 CS_BIAS.n162 0.189894
R747 CS_BIAS.n162 CS_BIAS.n157 0.189894
R748 CS_BIAS.n141 CS_BIAS.n99 0.189894
R749 CS_BIAS.n141 CS_BIAS.n140 0.189894
R750 CS_BIAS.n140 CS_BIAS.n139 0.189894
R751 CS_BIAS.n139 CS_BIAS.n101 0.189894
R752 CS_BIAS.n134 CS_BIAS.n101 0.189894
R753 CS_BIAS.n134 CS_BIAS.n133 0.189894
R754 CS_BIAS.n133 CS_BIAS.n132 0.189894
R755 CS_BIAS.n132 CS_BIAS.n103 0.189894
R756 CS_BIAS.n128 CS_BIAS.n103 0.189894
R757 CS_BIAS.n128 CS_BIAS.n127 0.189894
R758 CS_BIAS.n127 CS_BIAS.n105 0.189894
R759 CS_BIAS.n123 CS_BIAS.n105 0.189894
R760 CS_BIAS.n123 CS_BIAS.n122 0.189894
R761 CS_BIAS.n122 CS_BIAS.n121 0.189894
R762 CS_BIAS.n121 CS_BIAS.n107 0.189894
R763 CS_BIAS.n116 CS_BIAS.n107 0.189894
R764 CS_BIAS.n116 CS_BIAS.n115 0.189894
R765 CS_BIAS.n115 CS_BIAS.n114 0.189894
R766 CS_BIAS.n114 CS_BIAS.n109 0.189894
R767 CS_BIAS.n50 CS_BIAS.n8 0.189894
R768 CS_BIAS.n50 CS_BIAS.n49 0.189894
R769 CS_BIAS.n49 CS_BIAS.n48 0.189894
R770 CS_BIAS.n48 CS_BIAS.n10 0.189894
R771 CS_BIAS.n43 CS_BIAS.n10 0.189894
R772 CS_BIAS.n43 CS_BIAS.n42 0.189894
R773 CS_BIAS.n42 CS_BIAS.n41 0.189894
R774 CS_BIAS.n41 CS_BIAS.n12 0.189894
R775 CS_BIAS.n37 CS_BIAS.n12 0.189894
R776 CS_BIAS.n37 CS_BIAS.n36 0.189894
R777 CS_BIAS.n36 CS_BIAS.n14 0.189894
R778 CS_BIAS.n32 CS_BIAS.n14 0.189894
R779 CS_BIAS.n32 CS_BIAS.n31 0.189894
R780 CS_BIAS.n31 CS_BIAS.n30 0.189894
R781 CS_BIAS.n30 CS_BIAS.n16 0.189894
R782 CS_BIAS.n25 CS_BIAS.n16 0.189894
R783 CS_BIAS.n25 CS_BIAS.n24 0.189894
R784 CS_BIAS.n24 CS_BIAS.n23 0.189894
R785 CS_BIAS.n23 CS_BIAS.n18 0.189894
R786 CS_BIAS.n75 CS_BIAS.n74 0.189894
R787 CS_BIAS.n74 CS_BIAS.n60 0.189894
R788 CS_BIAS.n69 CS_BIAS.n60 0.189894
R789 CS_BIAS.n69 CS_BIAS.n68 0.189894
R790 CS_BIAS.n68 CS_BIAS.n67 0.189894
R791 CS_BIAS.n67 CS_BIAS.n62 0.189894
R792 CS_BIAS.n94 CS_BIAS.n0 0.189894
R793 CS_BIAS.n94 CS_BIAS.n93 0.189894
R794 CS_BIAS.n93 CS_BIAS.n92 0.189894
R795 CS_BIAS.n92 CS_BIAS.n2 0.189894
R796 CS_BIAS.n87 CS_BIAS.n2 0.189894
R797 CS_BIAS.n87 CS_BIAS.n86 0.189894
R798 CS_BIAS.n86 CS_BIAS.n85 0.189894
R799 CS_BIAS.n85 CS_BIAS.n4 0.189894
R800 CS_BIAS.n81 CS_BIAS.n4 0.189894
R801 CS_BIAS.n81 CS_BIAS.n80 0.189894
R802 CS_BIAS.n80 CS_BIAS.n6 0.189894
R803 CS_BIAS.n549 CS_BIAS.n544 0.189894
R804 CS_BIAS.n550 CS_BIAS.n549 0.189894
R805 CS_BIAS.n551 CS_BIAS.n550 0.189894
R806 CS_BIAS.n551 CS_BIAS.n542 0.189894
R807 CS_BIAS.n556 CS_BIAS.n542 0.189894
R808 CS_BIAS.n557 CS_BIAS.n556 0.189894
R809 CS_BIAS.n558 CS_BIAS.n557 0.189894
R810 CS_BIAS.n558 CS_BIAS.n540 0.189894
R811 CS_BIAS.n562 CS_BIAS.n540 0.189894
R812 CS_BIAS.n563 CS_BIAS.n562 0.189894
R813 CS_BIAS.n563 CS_BIAS.n538 0.189894
R814 CS_BIAS.n567 CS_BIAS.n538 0.189894
R815 CS_BIAS.n568 CS_BIAS.n567 0.189894
R816 CS_BIAS.n569 CS_BIAS.n568 0.189894
R817 CS_BIAS.n569 CS_BIAS.n536 0.189894
R818 CS_BIAS.n574 CS_BIAS.n536 0.189894
R819 CS_BIAS.n575 CS_BIAS.n574 0.189894
R820 CS_BIAS.n576 CS_BIAS.n575 0.189894
R821 CS_BIAS.n576 CS_BIAS.n534 0.189894
R822 CS_BIAS.n501 CS_BIAS.n496 0.189894
R823 CS_BIAS.n502 CS_BIAS.n501 0.189894
R824 CS_BIAS.n503 CS_BIAS.n502 0.189894
R825 CS_BIAS.n503 CS_BIAS.n494 0.189894
R826 CS_BIAS.n508 CS_BIAS.n494 0.189894
R827 CS_BIAS.n509 CS_BIAS.n508 0.189894
R828 CS_BIAS.n510 CS_BIAS.n509 0.189894
R829 CS_BIAS.n510 CS_BIAS.n492 0.189894
R830 CS_BIAS.n514 CS_BIAS.n492 0.189894
R831 CS_BIAS.n515 CS_BIAS.n514 0.189894
R832 CS_BIAS.n515 CS_BIAS.n490 0.189894
R833 CS_BIAS.n519 CS_BIAS.n490 0.189894
R834 CS_BIAS.n520 CS_BIAS.n519 0.189894
R835 CS_BIAS.n521 CS_BIAS.n520 0.189894
R836 CS_BIAS.n521 CS_BIAS.n488 0.189894
R837 CS_BIAS.n526 CS_BIAS.n488 0.189894
R838 CS_BIAS.n527 CS_BIAS.n526 0.189894
R839 CS_BIAS.n528 CS_BIAS.n527 0.189894
R840 CS_BIAS.n528 CS_BIAS.n486 0.189894
R841 CS_BIAS.n453 CS_BIAS.n448 0.189894
R842 CS_BIAS.n454 CS_BIAS.n453 0.189894
R843 CS_BIAS.n455 CS_BIAS.n454 0.189894
R844 CS_BIAS.n455 CS_BIAS.n446 0.189894
R845 CS_BIAS.n460 CS_BIAS.n446 0.189894
R846 CS_BIAS.n461 CS_BIAS.n460 0.189894
R847 CS_BIAS.n462 CS_BIAS.n461 0.189894
R848 CS_BIAS.n462 CS_BIAS.n444 0.189894
R849 CS_BIAS.n466 CS_BIAS.n444 0.189894
R850 CS_BIAS.n467 CS_BIAS.n466 0.189894
R851 CS_BIAS.n467 CS_BIAS.n442 0.189894
R852 CS_BIAS.n471 CS_BIAS.n442 0.189894
R853 CS_BIAS.n472 CS_BIAS.n471 0.189894
R854 CS_BIAS.n473 CS_BIAS.n472 0.189894
R855 CS_BIAS.n473 CS_BIAS.n440 0.189894
R856 CS_BIAS.n478 CS_BIAS.n440 0.189894
R857 CS_BIAS.n479 CS_BIAS.n478 0.189894
R858 CS_BIAS.n480 CS_BIAS.n479 0.189894
R859 CS_BIAS.n480 CS_BIAS.n438 0.189894
R860 CS_BIAS.n405 CS_BIAS.n400 0.189894
R861 CS_BIAS.n406 CS_BIAS.n405 0.189894
R862 CS_BIAS.n407 CS_BIAS.n406 0.189894
R863 CS_BIAS.n407 CS_BIAS.n398 0.189894
R864 CS_BIAS.n412 CS_BIAS.n398 0.189894
R865 CS_BIAS.n413 CS_BIAS.n412 0.189894
R866 CS_BIAS.n414 CS_BIAS.n413 0.189894
R867 CS_BIAS.n414 CS_BIAS.n396 0.189894
R868 CS_BIAS.n418 CS_BIAS.n396 0.189894
R869 CS_BIAS.n419 CS_BIAS.n418 0.189894
R870 CS_BIAS.n419 CS_BIAS.n394 0.189894
R871 CS_BIAS.n423 CS_BIAS.n394 0.189894
R872 CS_BIAS.n424 CS_BIAS.n423 0.189894
R873 CS_BIAS.n425 CS_BIAS.n424 0.189894
R874 CS_BIAS.n425 CS_BIAS.n392 0.189894
R875 CS_BIAS.n430 CS_BIAS.n392 0.189894
R876 CS_BIAS.n431 CS_BIAS.n430 0.189894
R877 CS_BIAS.n432 CS_BIAS.n431 0.189894
R878 CS_BIAS.n432 CS_BIAS.n390 0.189894
R879 CS_BIAS.n332 CS_BIAS.n327 0.189894
R880 CS_BIAS.n333 CS_BIAS.n332 0.189894
R881 CS_BIAS.n334 CS_BIAS.n333 0.189894
R882 CS_BIAS.n334 CS_BIAS.n325 0.189894
R883 CS_BIAS.n339 CS_BIAS.n325 0.189894
R884 CS_BIAS.n340 CS_BIAS.n339 0.189894
R885 CS_BIAS.n341 CS_BIAS.n340 0.189894
R886 CS_BIAS.n341 CS_BIAS.n323 0.189894
R887 CS_BIAS.n345 CS_BIAS.n323 0.189894
R888 CS_BIAS.n346 CS_BIAS.n345 0.189894
R889 CS_BIAS.n346 CS_BIAS.n321 0.189894
R890 CS_BIAS.n350 CS_BIAS.n321 0.189894
R891 CS_BIAS.n351 CS_BIAS.n350 0.189894
R892 CS_BIAS.n352 CS_BIAS.n351 0.189894
R893 CS_BIAS.n352 CS_BIAS.n319 0.189894
R894 CS_BIAS.n357 CS_BIAS.n319 0.189894
R895 CS_BIAS.n358 CS_BIAS.n357 0.189894
R896 CS_BIAS.n359 CS_BIAS.n358 0.189894
R897 CS_BIAS.n359 CS_BIAS.n317 0.189894
R898 CS_BIAS.n306 CS_BIAS.n301 0.189894
R899 CS_BIAS.n307 CS_BIAS.n306 0.189894
R900 CS_BIAS.n308 CS_BIAS.n307 0.189894
R901 CS_BIAS.n308 CS_BIAS.n299 0.189894
R902 CS_BIAS.n313 CS_BIAS.n299 0.189894
R903 CS_BIAS.n314 CS_BIAS.n313 0.189894
R904 CS_BIAS.n371 CS_BIAS.n297 0.189894
R905 CS_BIAS.n372 CS_BIAS.n371 0.189894
R906 CS_BIAS.n372 CS_BIAS.n295 0.189894
R907 CS_BIAS.n376 CS_BIAS.n295 0.189894
R908 CS_BIAS.n377 CS_BIAS.n376 0.189894
R909 CS_BIAS.n378 CS_BIAS.n377 0.189894
R910 CS_BIAS.n378 CS_BIAS.n293 0.189894
R911 CS_BIAS.n383 CS_BIAS.n293 0.189894
R912 CS_BIAS.n384 CS_BIAS.n383 0.189894
R913 CS_BIAS.n385 CS_BIAS.n384 0.189894
R914 CS_BIAS.n385 CS_BIAS.n291 0.189894
R915 CS_BIAS.n76 CS_BIAS.n75 0.170955
R916 CS_BIAS.n76 CS_BIAS.n6 0.170955
R917 CS_BIAS.n367 CS_BIAS.n314 0.170955
R918 CS_BIAS.n367 CS_BIAS.n297 0.170955
R919 VOUT.n23 VOUT.n21 174.619
R920 VOUT.n19 VOUT.n17 174.619
R921 VOUT.n16 VOUT.n14 174.619
R922 VOUT.n9 VOUT.n7 174.619
R923 VOUT.n5 VOUT.n3 174.619
R924 VOUT.n2 VOUT.n0 174.619
R925 VOUT.n19 VOUT.n18 171.81
R926 VOUT.n16 VOUT.n15 171.81
R927 VOUT.n9 VOUT.n8 171.81
R928 VOUT.n5 VOUT.n4 171.81
R929 VOUT.n2 VOUT.n1 171.81
R930 VOUT.n23 VOUT.n22 171.81
R931 VOUT.n51 VOUT.n49 75.2659
R932 VOUT.n45 VOUT.n43 75.2659
R933 VOUT.n39 VOUT.n37 75.2659
R934 VOUT.n33 VOUT.n31 75.2659
R935 VOUT.n28 VOUT.n26 75.2659
R936 VOUT.n81 VOUT.n79 75.2659
R937 VOUT.n75 VOUT.n73 75.2659
R938 VOUT.n69 VOUT.n67 75.2659
R939 VOUT.n63 VOUT.n61 75.2659
R940 VOUT.n58 VOUT.n56 75.2659
R941 VOUT.n53 VOUT.n52 73.0762
R942 VOUT.n51 VOUT.n50 73.0762
R943 VOUT.n47 VOUT.n46 73.0762
R944 VOUT.n45 VOUT.n44 73.0762
R945 VOUT.n41 VOUT.n40 73.0762
R946 VOUT.n39 VOUT.n38 73.0762
R947 VOUT.n35 VOUT.n34 73.0762
R948 VOUT.n33 VOUT.n32 73.0762
R949 VOUT.n30 VOUT.n29 73.0762
R950 VOUT.n28 VOUT.n27 73.0762
R951 VOUT.n81 VOUT.n80 73.0762
R952 VOUT.n83 VOUT.n82 73.0762
R953 VOUT.n75 VOUT.n74 73.0762
R954 VOUT.n77 VOUT.n76 73.0762
R955 VOUT.n69 VOUT.n68 73.0762
R956 VOUT.n71 VOUT.n70 73.0762
R957 VOUT.n63 VOUT.n62 73.0762
R958 VOUT.n65 VOUT.n64 73.0762
R959 VOUT.n58 VOUT.n57 73.0762
R960 VOUT.n60 VOUT.n59 73.0762
R961 VOUT.n22 VOUT.t5 15.5531
R962 VOUT.n22 VOUT.t9 15.5531
R963 VOUT.n21 VOUT.t20 15.5531
R964 VOUT.n21 VOUT.t11 15.5531
R965 VOUT.n18 VOUT.t6 15.5531
R966 VOUT.n18 VOUT.t82 15.5531
R967 VOUT.n17 VOUT.t15 15.5531
R968 VOUT.n17 VOUT.t17 15.5531
R969 VOUT.n15 VOUT.t16 15.5531
R970 VOUT.n15 VOUT.t1 15.5531
R971 VOUT.n14 VOUT.t10 15.5531
R972 VOUT.n14 VOUT.t13 15.5531
R973 VOUT.n7 VOUT.t3 15.5531
R974 VOUT.n7 VOUT.t19 15.5531
R975 VOUT.n8 VOUT.t7 15.5531
R976 VOUT.n8 VOUT.t14 15.5531
R977 VOUT.n3 VOUT.t83 15.5531
R978 VOUT.n3 VOUT.t2 15.5531
R979 VOUT.n4 VOUT.t8 15.5531
R980 VOUT.n4 VOUT.t12 15.5531
R981 VOUT.n0 VOUT.t18 15.5531
R982 VOUT.n0 VOUT.t4 15.5531
R983 VOUT.n1 VOUT.t0 15.5531
R984 VOUT.n1 VOUT.t81 15.5531
R985 VOUT.n55 VOUT.n25 9.64653
R986 VOUT.n36 VOUT.n30 9.05869
R987 VOUT.n66 VOUT.n60 9.05869
R988 VOUT.n20 VOUT.n16 8.6255
R989 VOUT.n6 VOUT.n2 8.6255
R990 VOUT.n25 VOUT.n24 7.44929
R991 VOUT.n11 VOUT.n10 7.44929
R992 VOUT.n24 VOUT.n23 6.80653
R993 VOUT.n20 VOUT.n19 6.80653
R994 VOUT.n10 VOUT.n9 6.80653
R995 VOUT.n6 VOUT.n5 6.80653
R996 VOUT.n54 VOUT.n53 6.49619
R997 VOUT.n48 VOUT.n47 6.49619
R998 VOUT.n42 VOUT.n41 6.49619
R999 VOUT.n36 VOUT.n35 6.49619
R1000 VOUT.n84 VOUT.n83 6.49619
R1001 VOUT.n78 VOUT.n77 6.49619
R1002 VOUT.n72 VOUT.n71 6.49619
R1003 VOUT.n66 VOUT.n65 6.49619
R1004 VOUT.n55 VOUT.n54 5.58291
R1005 VOUT.n85 VOUT.n84 5.58291
R1006 VOUT.n25 VOUT.n11 5.24382
R1007 VOUT.n52 VOUT.t34 5.18375
R1008 VOUT.n52 VOUT.t21 5.18375
R1009 VOUT.n50 VOUT.t49 5.18375
R1010 VOUT.n50 VOUT.t33 5.18375
R1011 VOUT.n49 VOUT.t66 5.18375
R1012 VOUT.n49 VOUT.t48 5.18375
R1013 VOUT.n46 VOUT.t31 5.18375
R1014 VOUT.n46 VOUT.t77 5.18375
R1015 VOUT.n44 VOUT.t41 5.18375
R1016 VOUT.n44 VOUT.t29 5.18375
R1017 VOUT.n43 VOUT.t57 5.18375
R1018 VOUT.n43 VOUT.t42 5.18375
R1019 VOUT.n40 VOUT.t40 5.18375
R1020 VOUT.n40 VOUT.t73 5.18375
R1021 VOUT.n38 VOUT.t78 5.18375
R1022 VOUT.n38 VOUT.t30 5.18375
R1023 VOUT.n37 VOUT.t61 5.18375
R1024 VOUT.n37 VOUT.t76 5.18375
R1025 VOUT.n34 VOUT.t22 5.18375
R1026 VOUT.n34 VOUT.t39 5.18375
R1027 VOUT.n32 VOUT.t80 5.18375
R1028 VOUT.n32 VOUT.t24 5.18375
R1029 VOUT.n31 VOUT.t63 5.18375
R1030 VOUT.n31 VOUT.t23 5.18375
R1031 VOUT.n29 VOUT.t35 5.18375
R1032 VOUT.n29 VOUT.t71 5.18375
R1033 VOUT.n27 VOUT.t53 5.18375
R1034 VOUT.n27 VOUT.t38 5.18375
R1035 VOUT.n26 VOUT.t68 5.18375
R1036 VOUT.n26 VOUT.t51 5.18375
R1037 VOUT.n79 VOUT.t54 5.18375
R1038 VOUT.n79 VOUT.t55 5.18375
R1039 VOUT.n80 VOUT.t50 5.18375
R1040 VOUT.n80 VOUT.t37 5.18375
R1041 VOUT.n82 VOUT.t45 5.18375
R1042 VOUT.n82 VOUT.t44 5.18375
R1043 VOUT.n73 VOUT.t28 5.18375
R1044 VOUT.n73 VOUT.t26 5.18375
R1045 VOUT.n74 VOUT.t65 5.18375
R1046 VOUT.n74 VOUT.t64 5.18375
R1047 VOUT.n76 VOUT.t46 5.18375
R1048 VOUT.n76 VOUT.t36 5.18375
R1049 VOUT.n67 VOUT.t75 5.18375
R1050 VOUT.n67 VOUT.t74 5.18375
R1051 VOUT.n68 VOUT.t27 5.18375
R1052 VOUT.n68 VOUT.t67 5.18375
R1053 VOUT.n70 VOUT.t70 5.18375
R1054 VOUT.n70 VOUT.t69 5.18375
R1055 VOUT.n61 VOUT.t32 5.18375
R1056 VOUT.n61 VOUT.t56 5.18375
R1057 VOUT.n62 VOUT.t47 5.18375
R1058 VOUT.n62 VOUT.t52 5.18375
R1059 VOUT.n64 VOUT.t62 5.18375
R1060 VOUT.n64 VOUT.t58 5.18375
R1061 VOUT.n56 VOUT.t59 5.18375
R1062 VOUT.n56 VOUT.t79 5.18375
R1063 VOUT.n57 VOUT.t60 5.18375
R1064 VOUT.n57 VOUT.t72 5.18375
R1065 VOUT.n59 VOUT.t25 5.18375
R1066 VOUT.n59 VOUT.t43 5.18375
R1067 VOUT.n86 VOUT.n85 5.08887
R1068 VOUT.n86 VOUT.n11 4.53866
R1069 VOUT.n13 VOUT 3.0978
R1070 VOUT.n42 VOUT.n36 2.563
R1071 VOUT.n48 VOUT.n42 2.563
R1072 VOUT.n54 VOUT.n48 2.563
R1073 VOUT.n72 VOUT.n66 2.563
R1074 VOUT.n78 VOUT.n72 2.563
R1075 VOUT.n84 VOUT.n78 2.563
R1076 VOUT.n85 VOUT.n55 2.32825
R1077 VOUT.n53 VOUT.n51 2.19016
R1078 VOUT.n47 VOUT.n45 2.19016
R1079 VOUT.n41 VOUT.n39 2.19016
R1080 VOUT.n35 VOUT.n33 2.19016
R1081 VOUT.n30 VOUT.n28 2.19016
R1082 VOUT.n83 VOUT.n81 2.19016
R1083 VOUT.n77 VOUT.n75 2.19016
R1084 VOUT.n71 VOUT.n69 2.19016
R1085 VOUT.n65 VOUT.n63 2.19016
R1086 VOUT.n60 VOUT.n58 2.19016
R1087 VOUT.n24 VOUT.n20 1.81947
R1088 VOUT.n10 VOUT.n6 1.81947
R1089 VOUT.n13 VOUT.n12 0.361443
R1090 VOUT.n86 VOUT.n13 0.30083
R1091 VOUT.n12 VOUT.t84 0.115453
R1092 VOUT.n12 VOUT.t85 0.0486886
R1093 VOUT VOUT.n86 0.0099
R1094 GND.n6289 GND.n6288 2183.32
R1095 GND.n5331 GND.n5330 1044.86
R1096 GND.n3773 GND.n3202 725.538
R1097 GND.n3815 GND.n3313 725.538
R1098 GND.n4818 GND.n2963 725.538
R1099 GND.n4850 GND.n2966 725.538
R1100 GND.n6794 GND.n643 703.915
R1101 GND.n778 GND.n646 703.915
R1102 GND.n4275 GND.n4104 703.915
R1103 GND.n4266 GND.n3934 703.915
R1104 GND.n2278 GND.n1878 703.915
R1105 GND.n2534 GND.n1876 703.915
R1106 GND.n2846 GND.n1989 703.915
R1107 GND.n2876 GND.n1987 703.915
R1108 GND.n5417 GND.n1594 694.306
R1109 GND.n6287 GND.n1072 694.306
R1110 GND.n6401 GND.n1001 694.306
R1111 GND.n5322 GND.n1683 694.306
R1112 GND.n6792 GND.n648 684.696
R1113 GND.n756 GND.n645 684.696
R1114 GND.n4273 GND.n4272 684.696
R1115 GND.n4629 GND.n3926 684.696
R1116 GND.n5055 GND.n1991 684.696
R1117 GND.n5057 GND.n1985 684.696
R1118 GND.n2501 GND.n1875 684.696
R1119 GND.n5133 GND.n1879 684.696
R1120 GND.n5419 GND.n5418 680.317
R1121 GND.n5417 GND.n5416 585
R1122 GND.n5418 GND.n5417 585
R1123 GND.n5415 GND.n1596 585
R1124 GND.n1596 GND.n1595 585
R1125 GND.n5414 GND.n5413 585
R1126 GND.n5413 GND.n5412 585
R1127 GND.n1601 GND.n1600 585
R1128 GND.n5411 GND.n1601 585
R1129 GND.n5409 GND.n5408 585
R1130 GND.n5410 GND.n5409 585
R1131 GND.n5407 GND.n1603 585
R1132 GND.n1603 GND.n1602 585
R1133 GND.n5406 GND.n5405 585
R1134 GND.n5405 GND.n5404 585
R1135 GND.n1609 GND.n1608 585
R1136 GND.n5403 GND.n1609 585
R1137 GND.n5401 GND.n5400 585
R1138 GND.n5402 GND.n5401 585
R1139 GND.n5399 GND.n1611 585
R1140 GND.n1611 GND.n1610 585
R1141 GND.n5398 GND.n5397 585
R1142 GND.n5397 GND.n5396 585
R1143 GND.n1617 GND.n1616 585
R1144 GND.n5395 GND.n1617 585
R1145 GND.n5393 GND.n5392 585
R1146 GND.n5394 GND.n5393 585
R1147 GND.n5391 GND.n1619 585
R1148 GND.n1619 GND.n1618 585
R1149 GND.n5390 GND.n5389 585
R1150 GND.n5389 GND.n5388 585
R1151 GND.n1625 GND.n1624 585
R1152 GND.n5387 GND.n1625 585
R1153 GND.n5385 GND.n5384 585
R1154 GND.n5386 GND.n5385 585
R1155 GND.n5383 GND.n1627 585
R1156 GND.n1627 GND.n1626 585
R1157 GND.n5382 GND.n5381 585
R1158 GND.n5381 GND.n5380 585
R1159 GND.n1633 GND.n1632 585
R1160 GND.n5379 GND.n1633 585
R1161 GND.n5377 GND.n5376 585
R1162 GND.n5378 GND.n5377 585
R1163 GND.n5375 GND.n1635 585
R1164 GND.n1635 GND.n1634 585
R1165 GND.n5374 GND.n5373 585
R1166 GND.n5373 GND.n5372 585
R1167 GND.n1641 GND.n1640 585
R1168 GND.n5371 GND.n1641 585
R1169 GND.n5369 GND.n5368 585
R1170 GND.n5370 GND.n5369 585
R1171 GND.n5367 GND.n1643 585
R1172 GND.n1643 GND.n1642 585
R1173 GND.n5366 GND.n5365 585
R1174 GND.n5365 GND.n5364 585
R1175 GND.n1649 GND.n1648 585
R1176 GND.n5363 GND.n1649 585
R1177 GND.n5361 GND.n5360 585
R1178 GND.n5362 GND.n5361 585
R1179 GND.n5359 GND.n1651 585
R1180 GND.n1651 GND.n1650 585
R1181 GND.n5358 GND.n5357 585
R1182 GND.n5357 GND.n5356 585
R1183 GND.n1657 GND.n1656 585
R1184 GND.n5355 GND.n1657 585
R1185 GND.n5353 GND.n5352 585
R1186 GND.n5354 GND.n5353 585
R1187 GND.n5351 GND.n1659 585
R1188 GND.n1659 GND.n1658 585
R1189 GND.n5350 GND.n5349 585
R1190 GND.n5349 GND.n5348 585
R1191 GND.n1665 GND.n1664 585
R1192 GND.n5347 GND.n1665 585
R1193 GND.n5345 GND.n5344 585
R1194 GND.n5346 GND.n5345 585
R1195 GND.n5343 GND.n1667 585
R1196 GND.n1667 GND.n1666 585
R1197 GND.n5342 GND.n5341 585
R1198 GND.n5341 GND.n5340 585
R1199 GND.n1673 GND.n1672 585
R1200 GND.n5339 GND.n1673 585
R1201 GND.n5337 GND.n5336 585
R1202 GND.n5338 GND.n5337 585
R1203 GND.n5335 GND.n1675 585
R1204 GND.n1675 GND.n1674 585
R1205 GND.n5334 GND.n5333 585
R1206 GND.n5333 GND.n5332 585
R1207 GND.n1681 GND.n1680 585
R1208 GND.n5331 GND.n1681 585
R1209 GND.n1594 GND.n1593 585
R1210 GND.n5419 GND.n1594 585
R1211 GND.n5422 GND.n5421 585
R1212 GND.n5421 GND.n5420 585
R1213 GND.n1591 GND.n1590 585
R1214 GND.n1590 GND.n1589 585
R1215 GND.n5427 GND.n5426 585
R1216 GND.n5428 GND.n5427 585
R1217 GND.n1588 GND.n1587 585
R1218 GND.n5429 GND.n1588 585
R1219 GND.n5432 GND.n5431 585
R1220 GND.n5431 GND.n5430 585
R1221 GND.n1585 GND.n1584 585
R1222 GND.n1584 GND.n1583 585
R1223 GND.n5437 GND.n5436 585
R1224 GND.n5438 GND.n5437 585
R1225 GND.n1582 GND.n1581 585
R1226 GND.n5439 GND.n1582 585
R1227 GND.n5442 GND.n5441 585
R1228 GND.n5441 GND.n5440 585
R1229 GND.n1579 GND.n1578 585
R1230 GND.n1578 GND.n1577 585
R1231 GND.n5447 GND.n5446 585
R1232 GND.n5448 GND.n5447 585
R1233 GND.n1576 GND.n1575 585
R1234 GND.n5449 GND.n1576 585
R1235 GND.n5452 GND.n5451 585
R1236 GND.n5451 GND.n5450 585
R1237 GND.n1573 GND.n1572 585
R1238 GND.n1572 GND.n1571 585
R1239 GND.n5457 GND.n5456 585
R1240 GND.n5458 GND.n5457 585
R1241 GND.n1570 GND.n1569 585
R1242 GND.n5459 GND.n1570 585
R1243 GND.n5462 GND.n5461 585
R1244 GND.n5461 GND.n5460 585
R1245 GND.n1567 GND.n1566 585
R1246 GND.n1566 GND.n1565 585
R1247 GND.n5467 GND.n5466 585
R1248 GND.n5468 GND.n5467 585
R1249 GND.n1564 GND.n1563 585
R1250 GND.n5469 GND.n1564 585
R1251 GND.n5472 GND.n5471 585
R1252 GND.n5471 GND.n5470 585
R1253 GND.n1561 GND.n1560 585
R1254 GND.n1560 GND.n1559 585
R1255 GND.n5477 GND.n5476 585
R1256 GND.n5478 GND.n5477 585
R1257 GND.n1558 GND.n1557 585
R1258 GND.n5479 GND.n1558 585
R1259 GND.n5482 GND.n5481 585
R1260 GND.n5481 GND.n5480 585
R1261 GND.n1555 GND.n1554 585
R1262 GND.n1554 GND.n1553 585
R1263 GND.n5487 GND.n5486 585
R1264 GND.n5488 GND.n5487 585
R1265 GND.n1552 GND.n1551 585
R1266 GND.n5489 GND.n1552 585
R1267 GND.n5492 GND.n5491 585
R1268 GND.n5491 GND.n5490 585
R1269 GND.n1549 GND.n1548 585
R1270 GND.n1548 GND.n1547 585
R1271 GND.n5497 GND.n5496 585
R1272 GND.n5498 GND.n5497 585
R1273 GND.n1546 GND.n1545 585
R1274 GND.n5499 GND.n1546 585
R1275 GND.n5502 GND.n5501 585
R1276 GND.n5501 GND.n5500 585
R1277 GND.n1543 GND.n1542 585
R1278 GND.n1542 GND.n1541 585
R1279 GND.n5507 GND.n5506 585
R1280 GND.n5508 GND.n5507 585
R1281 GND.n1540 GND.n1539 585
R1282 GND.n5509 GND.n1540 585
R1283 GND.n5512 GND.n5511 585
R1284 GND.n5511 GND.n5510 585
R1285 GND.n1537 GND.n1536 585
R1286 GND.n1536 GND.n1535 585
R1287 GND.n5517 GND.n5516 585
R1288 GND.n5518 GND.n5517 585
R1289 GND.n1534 GND.n1533 585
R1290 GND.n5519 GND.n1534 585
R1291 GND.n5522 GND.n5521 585
R1292 GND.n5521 GND.n5520 585
R1293 GND.n1531 GND.n1530 585
R1294 GND.n1530 GND.n1529 585
R1295 GND.n5527 GND.n5526 585
R1296 GND.n5528 GND.n5527 585
R1297 GND.n1528 GND.n1527 585
R1298 GND.n5529 GND.n1528 585
R1299 GND.n5532 GND.n5531 585
R1300 GND.n5531 GND.n5530 585
R1301 GND.n1525 GND.n1524 585
R1302 GND.n1524 GND.n1523 585
R1303 GND.n5537 GND.n5536 585
R1304 GND.n5538 GND.n5537 585
R1305 GND.n1522 GND.n1521 585
R1306 GND.n5539 GND.n1522 585
R1307 GND.n5542 GND.n5541 585
R1308 GND.n5541 GND.n5540 585
R1309 GND.n1519 GND.n1518 585
R1310 GND.n1518 GND.n1517 585
R1311 GND.n5547 GND.n5546 585
R1312 GND.n5548 GND.n5547 585
R1313 GND.n1516 GND.n1515 585
R1314 GND.n5549 GND.n1516 585
R1315 GND.n5552 GND.n5551 585
R1316 GND.n5551 GND.n5550 585
R1317 GND.n1513 GND.n1512 585
R1318 GND.n1512 GND.n1511 585
R1319 GND.n5557 GND.n5556 585
R1320 GND.n5558 GND.n5557 585
R1321 GND.n1510 GND.n1509 585
R1322 GND.n5559 GND.n1510 585
R1323 GND.n5562 GND.n5561 585
R1324 GND.n5561 GND.n5560 585
R1325 GND.n1507 GND.n1506 585
R1326 GND.n1506 GND.n1505 585
R1327 GND.n5567 GND.n5566 585
R1328 GND.n5568 GND.n5567 585
R1329 GND.n1504 GND.n1503 585
R1330 GND.n5569 GND.n1504 585
R1331 GND.n5572 GND.n5571 585
R1332 GND.n5571 GND.n5570 585
R1333 GND.n1501 GND.n1500 585
R1334 GND.n1500 GND.n1499 585
R1335 GND.n5577 GND.n5576 585
R1336 GND.n5578 GND.n5577 585
R1337 GND.n1498 GND.n1497 585
R1338 GND.n5579 GND.n1498 585
R1339 GND.n5582 GND.n5581 585
R1340 GND.n5581 GND.n5580 585
R1341 GND.n1495 GND.n1494 585
R1342 GND.n1494 GND.n1493 585
R1343 GND.n5587 GND.n5586 585
R1344 GND.n5588 GND.n5587 585
R1345 GND.n1492 GND.n1491 585
R1346 GND.n5589 GND.n1492 585
R1347 GND.n5592 GND.n5591 585
R1348 GND.n5591 GND.n5590 585
R1349 GND.n1489 GND.n1488 585
R1350 GND.n1488 GND.n1487 585
R1351 GND.n5597 GND.n5596 585
R1352 GND.n5598 GND.n5597 585
R1353 GND.n1486 GND.n1485 585
R1354 GND.n5599 GND.n1486 585
R1355 GND.n5602 GND.n5601 585
R1356 GND.n5601 GND.n5600 585
R1357 GND.n1483 GND.n1482 585
R1358 GND.n1482 GND.n1481 585
R1359 GND.n5607 GND.n5606 585
R1360 GND.n5608 GND.n5607 585
R1361 GND.n1480 GND.n1479 585
R1362 GND.n5609 GND.n1480 585
R1363 GND.n5612 GND.n5611 585
R1364 GND.n5611 GND.n5610 585
R1365 GND.n1477 GND.n1476 585
R1366 GND.n1476 GND.n1475 585
R1367 GND.n5617 GND.n5616 585
R1368 GND.n5618 GND.n5617 585
R1369 GND.n1474 GND.n1473 585
R1370 GND.n5619 GND.n1474 585
R1371 GND.n5622 GND.n5621 585
R1372 GND.n5621 GND.n5620 585
R1373 GND.n1471 GND.n1470 585
R1374 GND.n1470 GND.n1469 585
R1375 GND.n5627 GND.n5626 585
R1376 GND.n5628 GND.n5627 585
R1377 GND.n1468 GND.n1467 585
R1378 GND.n5629 GND.n1468 585
R1379 GND.n5632 GND.n5631 585
R1380 GND.n5631 GND.n5630 585
R1381 GND.n1465 GND.n1464 585
R1382 GND.n1464 GND.n1463 585
R1383 GND.n5637 GND.n5636 585
R1384 GND.n5638 GND.n5637 585
R1385 GND.n1462 GND.n1461 585
R1386 GND.n5639 GND.n1462 585
R1387 GND.n5642 GND.n5641 585
R1388 GND.n5641 GND.n5640 585
R1389 GND.n1459 GND.n1458 585
R1390 GND.n1458 GND.n1457 585
R1391 GND.n5647 GND.n5646 585
R1392 GND.n5648 GND.n5647 585
R1393 GND.n1456 GND.n1455 585
R1394 GND.n5649 GND.n1456 585
R1395 GND.n5652 GND.n5651 585
R1396 GND.n5651 GND.n5650 585
R1397 GND.n1453 GND.n1452 585
R1398 GND.n1452 GND.n1451 585
R1399 GND.n5657 GND.n5656 585
R1400 GND.n5658 GND.n5657 585
R1401 GND.n1450 GND.n1449 585
R1402 GND.n5659 GND.n1450 585
R1403 GND.n5662 GND.n5661 585
R1404 GND.n5661 GND.n5660 585
R1405 GND.n1447 GND.n1446 585
R1406 GND.n1446 GND.n1445 585
R1407 GND.n5667 GND.n5666 585
R1408 GND.n5668 GND.n5667 585
R1409 GND.n1444 GND.n1443 585
R1410 GND.n5669 GND.n1444 585
R1411 GND.n5672 GND.n5671 585
R1412 GND.n5671 GND.n5670 585
R1413 GND.n1441 GND.n1440 585
R1414 GND.n1440 GND.n1439 585
R1415 GND.n5677 GND.n5676 585
R1416 GND.n5678 GND.n5677 585
R1417 GND.n1438 GND.n1437 585
R1418 GND.n5679 GND.n1438 585
R1419 GND.n5682 GND.n5681 585
R1420 GND.n5681 GND.n5680 585
R1421 GND.n1435 GND.n1434 585
R1422 GND.n1434 GND.n1433 585
R1423 GND.n5687 GND.n5686 585
R1424 GND.n5688 GND.n5687 585
R1425 GND.n1432 GND.n1431 585
R1426 GND.n5689 GND.n1432 585
R1427 GND.n5692 GND.n5691 585
R1428 GND.n5691 GND.n5690 585
R1429 GND.n1429 GND.n1428 585
R1430 GND.n1428 GND.n1427 585
R1431 GND.n5697 GND.n5696 585
R1432 GND.n5698 GND.n5697 585
R1433 GND.n1426 GND.n1425 585
R1434 GND.n5699 GND.n1426 585
R1435 GND.n5702 GND.n5701 585
R1436 GND.n5701 GND.n5700 585
R1437 GND.n1423 GND.n1422 585
R1438 GND.n1422 GND.n1421 585
R1439 GND.n5707 GND.n5706 585
R1440 GND.n5708 GND.n5707 585
R1441 GND.n1420 GND.n1419 585
R1442 GND.n5709 GND.n1420 585
R1443 GND.n5712 GND.n5711 585
R1444 GND.n5711 GND.n5710 585
R1445 GND.n1417 GND.n1416 585
R1446 GND.n1416 GND.n1415 585
R1447 GND.n5717 GND.n5716 585
R1448 GND.n5718 GND.n5717 585
R1449 GND.n1414 GND.n1413 585
R1450 GND.n5719 GND.n1414 585
R1451 GND.n5722 GND.n5721 585
R1452 GND.n5721 GND.n5720 585
R1453 GND.n1411 GND.n1410 585
R1454 GND.n1410 GND.n1409 585
R1455 GND.n5727 GND.n5726 585
R1456 GND.n5728 GND.n5727 585
R1457 GND.n1408 GND.n1407 585
R1458 GND.n5729 GND.n1408 585
R1459 GND.n5732 GND.n5731 585
R1460 GND.n5731 GND.n5730 585
R1461 GND.n1405 GND.n1404 585
R1462 GND.n1404 GND.n1403 585
R1463 GND.n5737 GND.n5736 585
R1464 GND.n5738 GND.n5737 585
R1465 GND.n1402 GND.n1401 585
R1466 GND.n5739 GND.n1402 585
R1467 GND.n5742 GND.n5741 585
R1468 GND.n5741 GND.n5740 585
R1469 GND.n1399 GND.n1398 585
R1470 GND.n1398 GND.n1397 585
R1471 GND.n5747 GND.n5746 585
R1472 GND.n5748 GND.n5747 585
R1473 GND.n1396 GND.n1395 585
R1474 GND.n5749 GND.n1396 585
R1475 GND.n5752 GND.n5751 585
R1476 GND.n5751 GND.n5750 585
R1477 GND.n1393 GND.n1392 585
R1478 GND.n1392 GND.n1391 585
R1479 GND.n5757 GND.n5756 585
R1480 GND.n5758 GND.n5757 585
R1481 GND.n1390 GND.n1389 585
R1482 GND.n5759 GND.n1390 585
R1483 GND.n5762 GND.n5761 585
R1484 GND.n5761 GND.n5760 585
R1485 GND.n1387 GND.n1386 585
R1486 GND.n1386 GND.n1385 585
R1487 GND.n5767 GND.n5766 585
R1488 GND.n5768 GND.n5767 585
R1489 GND.n1384 GND.n1383 585
R1490 GND.n5769 GND.n1384 585
R1491 GND.n5772 GND.n5771 585
R1492 GND.n5771 GND.n5770 585
R1493 GND.n1381 GND.n1380 585
R1494 GND.n1380 GND.n1379 585
R1495 GND.n5777 GND.n5776 585
R1496 GND.n5778 GND.n5777 585
R1497 GND.n1378 GND.n1377 585
R1498 GND.n5779 GND.n1378 585
R1499 GND.n5782 GND.n5781 585
R1500 GND.n5781 GND.n5780 585
R1501 GND.n1375 GND.n1374 585
R1502 GND.n1374 GND.n1373 585
R1503 GND.n5787 GND.n5786 585
R1504 GND.n5788 GND.n5787 585
R1505 GND.n1372 GND.n1371 585
R1506 GND.n5789 GND.n1372 585
R1507 GND.n5792 GND.n5791 585
R1508 GND.n5791 GND.n5790 585
R1509 GND.n1369 GND.n1368 585
R1510 GND.n1368 GND.n1367 585
R1511 GND.n5797 GND.n5796 585
R1512 GND.n5798 GND.n5797 585
R1513 GND.n1366 GND.n1365 585
R1514 GND.n5799 GND.n1366 585
R1515 GND.n5802 GND.n5801 585
R1516 GND.n5801 GND.n5800 585
R1517 GND.n1363 GND.n1362 585
R1518 GND.n1362 GND.n1361 585
R1519 GND.n5807 GND.n5806 585
R1520 GND.n5808 GND.n5807 585
R1521 GND.n1360 GND.n1359 585
R1522 GND.n5809 GND.n1360 585
R1523 GND.n5812 GND.n5811 585
R1524 GND.n5811 GND.n5810 585
R1525 GND.n1357 GND.n1356 585
R1526 GND.n1356 GND.n1355 585
R1527 GND.n5817 GND.n5816 585
R1528 GND.n5818 GND.n5817 585
R1529 GND.n1354 GND.n1353 585
R1530 GND.n5819 GND.n1354 585
R1531 GND.n5822 GND.n5821 585
R1532 GND.n5821 GND.n5820 585
R1533 GND.n1351 GND.n1350 585
R1534 GND.n1350 GND.n1349 585
R1535 GND.n5827 GND.n5826 585
R1536 GND.n5828 GND.n5827 585
R1537 GND.n1348 GND.n1347 585
R1538 GND.n5829 GND.n1348 585
R1539 GND.n5832 GND.n5831 585
R1540 GND.n5831 GND.n5830 585
R1541 GND.n1345 GND.n1344 585
R1542 GND.n1344 GND.n1343 585
R1543 GND.n5837 GND.n5836 585
R1544 GND.n5838 GND.n5837 585
R1545 GND.n1342 GND.n1341 585
R1546 GND.n5839 GND.n1342 585
R1547 GND.n5842 GND.n5841 585
R1548 GND.n5841 GND.n5840 585
R1549 GND.n1339 GND.n1338 585
R1550 GND.n1338 GND.n1337 585
R1551 GND.n5847 GND.n5846 585
R1552 GND.n5848 GND.n5847 585
R1553 GND.n1336 GND.n1335 585
R1554 GND.n5849 GND.n1336 585
R1555 GND.n5852 GND.n5851 585
R1556 GND.n5851 GND.n5850 585
R1557 GND.n1333 GND.n1332 585
R1558 GND.n1332 GND.n1331 585
R1559 GND.n5857 GND.n5856 585
R1560 GND.n5858 GND.n5857 585
R1561 GND.n1330 GND.n1329 585
R1562 GND.n5859 GND.n1330 585
R1563 GND.n5862 GND.n5861 585
R1564 GND.n5861 GND.n5860 585
R1565 GND.n1327 GND.n1326 585
R1566 GND.n1326 GND.n1325 585
R1567 GND.n5867 GND.n5866 585
R1568 GND.n5868 GND.n5867 585
R1569 GND.n1324 GND.n1323 585
R1570 GND.n5869 GND.n1324 585
R1571 GND.n5872 GND.n5871 585
R1572 GND.n5871 GND.n5870 585
R1573 GND.n1321 GND.n1320 585
R1574 GND.n1320 GND.n1319 585
R1575 GND.n5877 GND.n5876 585
R1576 GND.n5878 GND.n5877 585
R1577 GND.n1318 GND.n1317 585
R1578 GND.n5879 GND.n1318 585
R1579 GND.n5882 GND.n5881 585
R1580 GND.n5881 GND.n5880 585
R1581 GND.n1315 GND.n1314 585
R1582 GND.n1314 GND.n1313 585
R1583 GND.n5887 GND.n5886 585
R1584 GND.n5888 GND.n5887 585
R1585 GND.n1312 GND.n1311 585
R1586 GND.n5889 GND.n1312 585
R1587 GND.n5892 GND.n5891 585
R1588 GND.n5891 GND.n5890 585
R1589 GND.n1309 GND.n1308 585
R1590 GND.n1308 GND.n1307 585
R1591 GND.n5897 GND.n5896 585
R1592 GND.n5898 GND.n5897 585
R1593 GND.n1306 GND.n1305 585
R1594 GND.n5899 GND.n1306 585
R1595 GND.n5902 GND.n5901 585
R1596 GND.n5901 GND.n5900 585
R1597 GND.n1303 GND.n1302 585
R1598 GND.n1302 GND.n1301 585
R1599 GND.n5907 GND.n5906 585
R1600 GND.n5908 GND.n5907 585
R1601 GND.n1300 GND.n1299 585
R1602 GND.n5909 GND.n1300 585
R1603 GND.n5912 GND.n5911 585
R1604 GND.n5911 GND.n5910 585
R1605 GND.n1297 GND.n1296 585
R1606 GND.n1296 GND.n1295 585
R1607 GND.n5917 GND.n5916 585
R1608 GND.n5918 GND.n5917 585
R1609 GND.n1294 GND.n1293 585
R1610 GND.n5919 GND.n1294 585
R1611 GND.n5922 GND.n5921 585
R1612 GND.n5921 GND.n5920 585
R1613 GND.n1291 GND.n1290 585
R1614 GND.n1290 GND.n1289 585
R1615 GND.n5927 GND.n5926 585
R1616 GND.n5928 GND.n5927 585
R1617 GND.n1288 GND.n1287 585
R1618 GND.n5929 GND.n1288 585
R1619 GND.n5932 GND.n5931 585
R1620 GND.n5931 GND.n5930 585
R1621 GND.n1285 GND.n1284 585
R1622 GND.n1284 GND.n1283 585
R1623 GND.n5937 GND.n5936 585
R1624 GND.n5938 GND.n5937 585
R1625 GND.n1282 GND.n1281 585
R1626 GND.n5939 GND.n1282 585
R1627 GND.n5942 GND.n5941 585
R1628 GND.n5941 GND.n5940 585
R1629 GND.n1279 GND.n1278 585
R1630 GND.n1278 GND.n1277 585
R1631 GND.n5947 GND.n5946 585
R1632 GND.n5948 GND.n5947 585
R1633 GND.n1276 GND.n1275 585
R1634 GND.n5949 GND.n1276 585
R1635 GND.n5952 GND.n5951 585
R1636 GND.n5951 GND.n5950 585
R1637 GND.n1273 GND.n1272 585
R1638 GND.n1272 GND.n1271 585
R1639 GND.n5957 GND.n5956 585
R1640 GND.n5958 GND.n5957 585
R1641 GND.n1270 GND.n1269 585
R1642 GND.n5959 GND.n1270 585
R1643 GND.n5962 GND.n5961 585
R1644 GND.n5961 GND.n5960 585
R1645 GND.n1267 GND.n1266 585
R1646 GND.n1266 GND.n1265 585
R1647 GND.n5967 GND.n5966 585
R1648 GND.n5968 GND.n5967 585
R1649 GND.n1264 GND.n1263 585
R1650 GND.n5969 GND.n1264 585
R1651 GND.n5972 GND.n5971 585
R1652 GND.n5971 GND.n5970 585
R1653 GND.n1261 GND.n1260 585
R1654 GND.n1260 GND.n1259 585
R1655 GND.n5977 GND.n5976 585
R1656 GND.n5978 GND.n5977 585
R1657 GND.n1258 GND.n1257 585
R1658 GND.n5979 GND.n1258 585
R1659 GND.n5982 GND.n5981 585
R1660 GND.n5981 GND.n5980 585
R1661 GND.n1255 GND.n1254 585
R1662 GND.n1254 GND.n1253 585
R1663 GND.n5987 GND.n5986 585
R1664 GND.n5988 GND.n5987 585
R1665 GND.n1252 GND.n1251 585
R1666 GND.n5989 GND.n1252 585
R1667 GND.n5992 GND.n5991 585
R1668 GND.n5991 GND.n5990 585
R1669 GND.n1249 GND.n1248 585
R1670 GND.n1248 GND.n1247 585
R1671 GND.n5997 GND.n5996 585
R1672 GND.n5998 GND.n5997 585
R1673 GND.n1246 GND.n1245 585
R1674 GND.n5999 GND.n1246 585
R1675 GND.n6002 GND.n6001 585
R1676 GND.n6001 GND.n6000 585
R1677 GND.n1243 GND.n1242 585
R1678 GND.n1242 GND.n1241 585
R1679 GND.n6007 GND.n6006 585
R1680 GND.n6008 GND.n6007 585
R1681 GND.n1240 GND.n1239 585
R1682 GND.n6009 GND.n1240 585
R1683 GND.n6012 GND.n6011 585
R1684 GND.n6011 GND.n6010 585
R1685 GND.n1237 GND.n1236 585
R1686 GND.n1236 GND.n1235 585
R1687 GND.n6017 GND.n6016 585
R1688 GND.n6018 GND.n6017 585
R1689 GND.n1234 GND.n1233 585
R1690 GND.n6019 GND.n1234 585
R1691 GND.n6022 GND.n6021 585
R1692 GND.n6021 GND.n6020 585
R1693 GND.n1231 GND.n1230 585
R1694 GND.n1230 GND.n1229 585
R1695 GND.n6027 GND.n6026 585
R1696 GND.n6028 GND.n6027 585
R1697 GND.n1228 GND.n1227 585
R1698 GND.n6029 GND.n1228 585
R1699 GND.n6032 GND.n6031 585
R1700 GND.n6031 GND.n6030 585
R1701 GND.n1225 GND.n1224 585
R1702 GND.n1224 GND.n1223 585
R1703 GND.n6037 GND.n6036 585
R1704 GND.n6038 GND.n6037 585
R1705 GND.n1222 GND.n1221 585
R1706 GND.n6039 GND.n1222 585
R1707 GND.n6042 GND.n6041 585
R1708 GND.n6041 GND.n6040 585
R1709 GND.n1219 GND.n1218 585
R1710 GND.n1218 GND.n1217 585
R1711 GND.n6047 GND.n6046 585
R1712 GND.n6048 GND.n6047 585
R1713 GND.n1216 GND.n1215 585
R1714 GND.n6049 GND.n1216 585
R1715 GND.n6052 GND.n6051 585
R1716 GND.n6051 GND.n6050 585
R1717 GND.n1213 GND.n1212 585
R1718 GND.n1212 GND.n1211 585
R1719 GND.n6057 GND.n6056 585
R1720 GND.n6058 GND.n6057 585
R1721 GND.n1210 GND.n1209 585
R1722 GND.n6059 GND.n1210 585
R1723 GND.n6062 GND.n6061 585
R1724 GND.n6061 GND.n6060 585
R1725 GND.n1207 GND.n1206 585
R1726 GND.n1206 GND.n1205 585
R1727 GND.n6067 GND.n6066 585
R1728 GND.n6068 GND.n6067 585
R1729 GND.n1204 GND.n1203 585
R1730 GND.n6069 GND.n1204 585
R1731 GND.n6072 GND.n6071 585
R1732 GND.n6071 GND.n6070 585
R1733 GND.n1201 GND.n1200 585
R1734 GND.n1200 GND.n1199 585
R1735 GND.n6077 GND.n6076 585
R1736 GND.n6078 GND.n6077 585
R1737 GND.n1198 GND.n1197 585
R1738 GND.n6079 GND.n1198 585
R1739 GND.n6082 GND.n6081 585
R1740 GND.n6081 GND.n6080 585
R1741 GND.n1195 GND.n1194 585
R1742 GND.n1194 GND.n1193 585
R1743 GND.n6087 GND.n6086 585
R1744 GND.n6088 GND.n6087 585
R1745 GND.n1192 GND.n1191 585
R1746 GND.n6089 GND.n1192 585
R1747 GND.n6092 GND.n6091 585
R1748 GND.n6091 GND.n6090 585
R1749 GND.n1189 GND.n1188 585
R1750 GND.n1188 GND.n1187 585
R1751 GND.n6097 GND.n6096 585
R1752 GND.n6098 GND.n6097 585
R1753 GND.n1186 GND.n1185 585
R1754 GND.n6099 GND.n1186 585
R1755 GND.n6102 GND.n6101 585
R1756 GND.n6101 GND.n6100 585
R1757 GND.n1183 GND.n1182 585
R1758 GND.n1182 GND.n1181 585
R1759 GND.n6107 GND.n6106 585
R1760 GND.n6108 GND.n6107 585
R1761 GND.n1180 GND.n1179 585
R1762 GND.n6109 GND.n1180 585
R1763 GND.n6112 GND.n6111 585
R1764 GND.n6111 GND.n6110 585
R1765 GND.n1177 GND.n1176 585
R1766 GND.n1176 GND.n1175 585
R1767 GND.n6117 GND.n6116 585
R1768 GND.n6118 GND.n6117 585
R1769 GND.n1174 GND.n1173 585
R1770 GND.n6119 GND.n1174 585
R1771 GND.n6122 GND.n6121 585
R1772 GND.n6121 GND.n6120 585
R1773 GND.n1171 GND.n1170 585
R1774 GND.n1170 GND.n1169 585
R1775 GND.n6127 GND.n6126 585
R1776 GND.n6128 GND.n6127 585
R1777 GND.n1168 GND.n1167 585
R1778 GND.n6129 GND.n1168 585
R1779 GND.n6132 GND.n6131 585
R1780 GND.n6131 GND.n6130 585
R1781 GND.n1165 GND.n1164 585
R1782 GND.n1164 GND.n1163 585
R1783 GND.n6137 GND.n6136 585
R1784 GND.n6138 GND.n6137 585
R1785 GND.n1162 GND.n1161 585
R1786 GND.n6139 GND.n1162 585
R1787 GND.n6142 GND.n6141 585
R1788 GND.n6141 GND.n6140 585
R1789 GND.n1159 GND.n1158 585
R1790 GND.n1158 GND.n1157 585
R1791 GND.n6147 GND.n6146 585
R1792 GND.n6148 GND.n6147 585
R1793 GND.n1156 GND.n1155 585
R1794 GND.n6149 GND.n1156 585
R1795 GND.n6152 GND.n6151 585
R1796 GND.n6151 GND.n6150 585
R1797 GND.n1153 GND.n1152 585
R1798 GND.n1152 GND.n1151 585
R1799 GND.n6157 GND.n6156 585
R1800 GND.n6158 GND.n6157 585
R1801 GND.n1150 GND.n1149 585
R1802 GND.n6159 GND.n1150 585
R1803 GND.n6162 GND.n6161 585
R1804 GND.n6161 GND.n6160 585
R1805 GND.n1147 GND.n1146 585
R1806 GND.n1146 GND.n1145 585
R1807 GND.n6167 GND.n6166 585
R1808 GND.n6168 GND.n6167 585
R1809 GND.n1144 GND.n1143 585
R1810 GND.n6169 GND.n1144 585
R1811 GND.n6172 GND.n6171 585
R1812 GND.n6171 GND.n6170 585
R1813 GND.n1141 GND.n1140 585
R1814 GND.n1140 GND.n1139 585
R1815 GND.n6177 GND.n6176 585
R1816 GND.n6178 GND.n6177 585
R1817 GND.n1138 GND.n1137 585
R1818 GND.n6179 GND.n1138 585
R1819 GND.n6182 GND.n6181 585
R1820 GND.n6181 GND.n6180 585
R1821 GND.n1135 GND.n1134 585
R1822 GND.n1134 GND.n1133 585
R1823 GND.n6187 GND.n6186 585
R1824 GND.n6188 GND.n6187 585
R1825 GND.n1132 GND.n1131 585
R1826 GND.n6189 GND.n1132 585
R1827 GND.n6192 GND.n6191 585
R1828 GND.n6191 GND.n6190 585
R1829 GND.n1129 GND.n1128 585
R1830 GND.n1128 GND.n1127 585
R1831 GND.n6197 GND.n6196 585
R1832 GND.n6198 GND.n6197 585
R1833 GND.n1126 GND.n1125 585
R1834 GND.n6199 GND.n1126 585
R1835 GND.n6202 GND.n6201 585
R1836 GND.n6201 GND.n6200 585
R1837 GND.n1123 GND.n1122 585
R1838 GND.n1122 GND.n1121 585
R1839 GND.n6207 GND.n6206 585
R1840 GND.n6208 GND.n6207 585
R1841 GND.n1120 GND.n1119 585
R1842 GND.n6209 GND.n1120 585
R1843 GND.n6212 GND.n6211 585
R1844 GND.n6211 GND.n6210 585
R1845 GND.n1117 GND.n1116 585
R1846 GND.n1116 GND.n1115 585
R1847 GND.n6217 GND.n6216 585
R1848 GND.n6218 GND.n6217 585
R1849 GND.n1114 GND.n1113 585
R1850 GND.n6219 GND.n1114 585
R1851 GND.n6222 GND.n6221 585
R1852 GND.n6221 GND.n6220 585
R1853 GND.n1111 GND.n1110 585
R1854 GND.n1110 GND.n1109 585
R1855 GND.n6227 GND.n6226 585
R1856 GND.n6228 GND.n6227 585
R1857 GND.n1108 GND.n1107 585
R1858 GND.n6229 GND.n1108 585
R1859 GND.n6232 GND.n6231 585
R1860 GND.n6231 GND.n6230 585
R1861 GND.n1105 GND.n1104 585
R1862 GND.n1104 GND.n1103 585
R1863 GND.n6237 GND.n6236 585
R1864 GND.n6238 GND.n6237 585
R1865 GND.n1102 GND.n1101 585
R1866 GND.n6239 GND.n1102 585
R1867 GND.n6242 GND.n6241 585
R1868 GND.n6241 GND.n6240 585
R1869 GND.n1099 GND.n1098 585
R1870 GND.n1098 GND.n1097 585
R1871 GND.n6247 GND.n6246 585
R1872 GND.n6248 GND.n6247 585
R1873 GND.n1096 GND.n1095 585
R1874 GND.n6249 GND.n1096 585
R1875 GND.n6252 GND.n6251 585
R1876 GND.n6251 GND.n6250 585
R1877 GND.n1093 GND.n1092 585
R1878 GND.n1092 GND.n1091 585
R1879 GND.n6257 GND.n6256 585
R1880 GND.n6258 GND.n6257 585
R1881 GND.n1090 GND.n1089 585
R1882 GND.n6259 GND.n1090 585
R1883 GND.n6262 GND.n6261 585
R1884 GND.n6261 GND.n6260 585
R1885 GND.n1087 GND.n1086 585
R1886 GND.n1086 GND.n1085 585
R1887 GND.n6267 GND.n6266 585
R1888 GND.n6268 GND.n6267 585
R1889 GND.n1084 GND.n1083 585
R1890 GND.n6269 GND.n1084 585
R1891 GND.n6272 GND.n6271 585
R1892 GND.n6271 GND.n6270 585
R1893 GND.n1081 GND.n1080 585
R1894 GND.n1080 GND.n1079 585
R1895 GND.n6277 GND.n6276 585
R1896 GND.n6278 GND.n6277 585
R1897 GND.n1078 GND.n1077 585
R1898 GND.n6279 GND.n1078 585
R1899 GND.n6282 GND.n6281 585
R1900 GND.n6281 GND.n6280 585
R1901 GND.n1075 GND.n1074 585
R1902 GND.n1074 GND.n1073 585
R1903 GND.n6287 GND.n6286 585
R1904 GND.n6288 GND.n6287 585
R1905 GND.n6397 GND.n6396 585
R1906 GND.n6398 GND.n6397 585
R1907 GND.n1009 GND.n1008 585
R1908 GND.n1008 GND.n1007 585
R1909 GND.n6392 GND.n6391 585
R1910 GND.n6391 GND.n6390 585
R1911 GND.n1012 GND.n1011 585
R1912 GND.n6389 GND.n1012 585
R1913 GND.n6387 GND.n6386 585
R1914 GND.n6388 GND.n6387 585
R1915 GND.n1015 GND.n1014 585
R1916 GND.n1014 GND.n1013 585
R1917 GND.n6382 GND.n6381 585
R1918 GND.n6381 GND.n6380 585
R1919 GND.n1018 GND.n1017 585
R1920 GND.n6379 GND.n1018 585
R1921 GND.n6377 GND.n6376 585
R1922 GND.n6378 GND.n6377 585
R1923 GND.n1021 GND.n1020 585
R1924 GND.n1020 GND.n1019 585
R1925 GND.n6372 GND.n6371 585
R1926 GND.n6371 GND.n6370 585
R1927 GND.n1024 GND.n1023 585
R1928 GND.n6369 GND.n1024 585
R1929 GND.n6367 GND.n6366 585
R1930 GND.n6368 GND.n6367 585
R1931 GND.n1027 GND.n1026 585
R1932 GND.n1026 GND.n1025 585
R1933 GND.n6362 GND.n6361 585
R1934 GND.n6361 GND.n6360 585
R1935 GND.n1030 GND.n1029 585
R1936 GND.n6359 GND.n1030 585
R1937 GND.n6357 GND.n6356 585
R1938 GND.n6358 GND.n6357 585
R1939 GND.n1033 GND.n1032 585
R1940 GND.n1032 GND.n1031 585
R1941 GND.n6352 GND.n6351 585
R1942 GND.n6351 GND.n6350 585
R1943 GND.n1036 GND.n1035 585
R1944 GND.n6349 GND.n1036 585
R1945 GND.n6347 GND.n6346 585
R1946 GND.n6348 GND.n6347 585
R1947 GND.n1039 GND.n1038 585
R1948 GND.n1038 GND.n1037 585
R1949 GND.n6342 GND.n6341 585
R1950 GND.n6341 GND.n6340 585
R1951 GND.n1042 GND.n1041 585
R1952 GND.n6339 GND.n1042 585
R1953 GND.n6337 GND.n6336 585
R1954 GND.n6338 GND.n6337 585
R1955 GND.n1045 GND.n1044 585
R1956 GND.n1044 GND.n1043 585
R1957 GND.n6332 GND.n6331 585
R1958 GND.n6331 GND.n6330 585
R1959 GND.n1048 GND.n1047 585
R1960 GND.n6329 GND.n1048 585
R1961 GND.n6327 GND.n6326 585
R1962 GND.n6328 GND.n6327 585
R1963 GND.n1051 GND.n1050 585
R1964 GND.n1050 GND.n1049 585
R1965 GND.n6322 GND.n6321 585
R1966 GND.n6321 GND.n6320 585
R1967 GND.n1054 GND.n1053 585
R1968 GND.n6319 GND.n1054 585
R1969 GND.n6317 GND.n6316 585
R1970 GND.n6318 GND.n6317 585
R1971 GND.n1057 GND.n1056 585
R1972 GND.n1056 GND.n1055 585
R1973 GND.n6312 GND.n6311 585
R1974 GND.n6311 GND.n6310 585
R1975 GND.n1060 GND.n1059 585
R1976 GND.n6309 GND.n1060 585
R1977 GND.n6307 GND.n6306 585
R1978 GND.n6308 GND.n6307 585
R1979 GND.n1063 GND.n1062 585
R1980 GND.n1062 GND.n1061 585
R1981 GND.n6302 GND.n6301 585
R1982 GND.n6301 GND.n6300 585
R1983 GND.n1066 GND.n1065 585
R1984 GND.n6299 GND.n1066 585
R1985 GND.n6297 GND.n6296 585
R1986 GND.n6298 GND.n6297 585
R1987 GND.n1069 GND.n1068 585
R1988 GND.n1068 GND.n1067 585
R1989 GND.n6292 GND.n6291 585
R1990 GND.n6291 GND.n6290 585
R1991 GND.n1072 GND.n1071 585
R1992 GND.n6289 GND.n1072 585
R1993 GND.n6795 GND.n6794 585
R1994 GND.n6794 GND.n6793 585
R1995 GND.n6796 GND.n639 585
R1996 GND.n6648 GND.n639 585
R1997 GND.n6798 GND.n6797 585
R1998 GND.n6799 GND.n6798 585
R1999 GND.n623 GND.n622 585
R2000 GND.n6641 GND.n623 585
R2001 GND.n6807 GND.n6806 585
R2002 GND.n6806 GND.n6805 585
R2003 GND.n6808 GND.n618 585
R2004 GND.n6632 GND.n618 585
R2005 GND.n6810 GND.n6809 585
R2006 GND.n6811 GND.n6810 585
R2007 GND.n602 GND.n601 585
R2008 GND.n6626 GND.n602 585
R2009 GND.n6819 GND.n6818 585
R2010 GND.n6818 GND.n6817 585
R2011 GND.n6820 GND.n597 585
R2012 GND.n6618 GND.n597 585
R2013 GND.n6822 GND.n6821 585
R2014 GND.n6823 GND.n6822 585
R2015 GND.n582 GND.n581 585
R2016 GND.n6612 GND.n582 585
R2017 GND.n6831 GND.n6830 585
R2018 GND.n6830 GND.n6829 585
R2019 GND.n6832 GND.n577 585
R2020 GND.n4428 GND.n577 585
R2021 GND.n6834 GND.n6833 585
R2022 GND.n6835 GND.n6834 585
R2023 GND.n562 GND.n561 585
R2024 GND.n4434 GND.n562 585
R2025 GND.n6843 GND.n6842 585
R2026 GND.n6842 GND.n6841 585
R2027 GND.n6844 GND.n556 585
R2028 GND.n4440 GND.n556 585
R2029 GND.n6846 GND.n6845 585
R2030 GND.n6847 GND.n6846 585
R2031 GND.n557 GND.n555 585
R2032 GND.n4446 GND.n555 585
R2033 GND.n4458 GND.n4457 585
R2034 GND.n4457 GND.n4456 585
R2035 GND.n4459 GND.n4365 585
R2036 GND.n4452 GND.n4365 585
R2037 GND.n4461 GND.n4460 585
R2038 GND.n4462 GND.n4461 585
R2039 GND.n4053 GND.n536 585
R2040 GND.n6855 GND.n536 585
R2041 GND.n4470 GND.n4469 585
R2042 GND.n4469 GND.n4468 585
R2043 GND.n4471 GND.n4042 585
R2044 GND.n4479 GND.n4042 585
R2045 GND.n4473 GND.n4472 585
R2046 GND.n4474 GND.n4473 585
R2047 GND.n4049 GND.n4048 585
R2048 GND.n4048 GND.n4033 585
R2049 GND.n4025 GND.n4024 585
R2050 GND.n4488 GND.n4025 585
R2051 GND.n4495 GND.n4494 585
R2052 GND.n4494 GND.n4493 585
R2053 GND.n4496 GND.n4020 585
R2054 GND.n4349 GND.n4020 585
R2055 GND.n4498 GND.n4497 585
R2056 GND.n4499 GND.n4498 585
R2057 GND.n4004 GND.n4003 585
R2058 GND.n4330 GND.n4004 585
R2059 GND.n4507 GND.n4506 585
R2060 GND.n4506 GND.n4505 585
R2061 GND.n4508 GND.n3999 585
R2062 GND.n4323 GND.n3999 585
R2063 GND.n4510 GND.n4509 585
R2064 GND.n4511 GND.n4510 585
R2065 GND.n3983 GND.n3982 585
R2066 GND.n4315 GND.n3983 585
R2067 GND.n4519 GND.n4518 585
R2068 GND.n4518 GND.n4517 585
R2069 GND.n4520 GND.n3977 585
R2070 GND.n4308 GND.n3977 585
R2071 GND.n4522 GND.n4521 585
R2072 GND.n4523 GND.n4522 585
R2073 GND.n3978 GND.n3976 585
R2074 GND.n4300 GND.n3976 585
R2075 GND.n4295 GND.n3958 585
R2076 GND.n4529 GND.n3958 585
R2077 GND.n4294 GND.n4293 585
R2078 GND.n4293 GND.n3954 585
R2079 GND.n4292 GND.n4291 585
R2080 GND.n4292 GND.n3944 585
R2081 GND.n3937 GND.n3935 585
R2082 GND.n4537 GND.n3935 585
R2083 GND.n4543 GND.n4542 585
R2084 GND.n4544 GND.n4543 585
R2085 GND.n3936 GND.n3934 585
R2086 GND.n4274 GND.n3934 585
R2087 GND.n4267 GND.n4266 585
R2088 GND.n4265 GND.n4264 585
R2089 GND.n4263 GND.n4262 585
R2090 GND.n4261 GND.n4260 585
R2091 GND.n4259 GND.n4258 585
R2092 GND.n4257 GND.n4256 585
R2093 GND.n4255 GND.n4254 585
R2094 GND.n4253 GND.n4252 585
R2095 GND.n4251 GND.n4250 585
R2096 GND.n4249 GND.n4240 585
R2097 GND.n4244 GND.n4241 585
R2098 GND.n4245 GND.n4104 585
R2099 GND.n779 GND.n778 585
R2100 GND.n6655 GND.n774 585
R2101 GND.n6657 GND.n6656 585
R2102 GND.n6659 GND.n772 585
R2103 GND.n6661 GND.n6660 585
R2104 GND.n6662 GND.n766 585
R2105 GND.n6664 GND.n6663 585
R2106 GND.n6666 GND.n765 585
R2107 GND.n6667 GND.n764 585
R2108 GND.n6670 GND.n6669 585
R2109 GND.n6671 GND.n762 585
R2110 GND.n6672 GND.n643 585
R2111 GND.n6651 GND.n646 585
R2112 GND.n6793 GND.n646 585
R2113 GND.n6650 GND.n6649 585
R2114 GND.n6649 GND.n6648 585
R2115 GND.n783 GND.n637 585
R2116 GND.n6799 GND.n637 585
R2117 GND.n6640 GND.n6639 585
R2118 GND.n6641 GND.n6640 585
R2119 GND.n786 GND.n626 585
R2120 GND.n6805 GND.n626 585
R2121 GND.n6634 GND.n6633 585
R2122 GND.n6633 GND.n6632 585
R2123 GND.n788 GND.n616 585
R2124 GND.n6811 GND.n616 585
R2125 GND.n6625 GND.n6624 585
R2126 GND.n6626 GND.n6625 585
R2127 GND.n791 GND.n605 585
R2128 GND.n6817 GND.n605 585
R2129 GND.n6620 GND.n6619 585
R2130 GND.n6619 GND.n6618 585
R2131 GND.n793 GND.n595 585
R2132 GND.n6823 GND.n595 585
R2133 GND.n4424 GND.n796 585
R2134 GND.n6612 GND.n796 585
R2135 GND.n4425 GND.n585 585
R2136 GND.n6829 GND.n585 585
R2137 GND.n4427 GND.n4426 585
R2138 GND.n4428 GND.n4427 585
R2139 GND.n4418 GND.n575 585
R2140 GND.n6835 GND.n575 585
R2141 GND.n4436 GND.n4435 585
R2142 GND.n4435 GND.n4434 585
R2143 GND.n4437 GND.n565 585
R2144 GND.n6841 GND.n565 585
R2145 GND.n4439 GND.n4438 585
R2146 GND.n4440 GND.n4439 585
R2147 GND.n4410 GND.n553 585
R2148 GND.n6847 GND.n553 585
R2149 GND.n4448 GND.n4447 585
R2150 GND.n4447 GND.n4446 585
R2151 GND.n4449 GND.n4370 585
R2152 GND.n4456 GND.n4370 585
R2153 GND.n4451 GND.n4450 585
R2154 GND.n4452 GND.n4451 585
R2155 GND.n532 GND.n530 585
R2156 GND.n4462 GND.n532 585
R2157 GND.n6857 GND.n6856 585
R2158 GND.n6856 GND.n6855 585
R2159 GND.n531 GND.n529 585
R2160 GND.n4468 GND.n531 585
R2161 GND.n4341 GND.n4040 585
R2162 GND.n4479 GND.n4040 585
R2163 GND.n4342 GND.n4047 585
R2164 GND.n4474 GND.n4047 585
R2165 GND.n4344 GND.n4343 585
R2166 GND.n4343 GND.n4033 585
R2167 GND.n4345 GND.n4032 585
R2168 GND.n4488 GND.n4032 585
R2169 GND.n4346 GND.n4028 585
R2170 GND.n4493 GND.n4028 585
R2171 GND.n4348 GND.n4347 585
R2172 GND.n4349 GND.n4348 585
R2173 GND.n4091 GND.n4019 585
R2174 GND.n4499 GND.n4019 585
R2175 GND.n4332 GND.n4331 585
R2176 GND.n4331 GND.n4330 585
R2177 GND.n4093 GND.n4007 585
R2178 GND.n4505 GND.n4007 585
R2179 GND.n4322 GND.n4321 585
R2180 GND.n4323 GND.n4322 585
R2181 GND.n4095 GND.n3997 585
R2182 GND.n4511 GND.n3997 585
R2183 GND.n4317 GND.n4316 585
R2184 GND.n4316 GND.n4315 585
R2185 GND.n4097 GND.n3986 585
R2186 GND.n4517 GND.n3986 585
R2187 GND.n4307 GND.n4306 585
R2188 GND.n4308 GND.n4307 585
R2189 GND.n4099 GND.n3974 585
R2190 GND.n4523 GND.n3974 585
R2191 GND.n4302 GND.n4301 585
R2192 GND.n4301 GND.n4300 585
R2193 GND.n4285 GND.n3956 585
R2194 GND.n4529 GND.n3956 585
R2195 GND.n4284 GND.n4283 585
R2196 GND.n4283 GND.n3954 585
R2197 GND.n4282 GND.n4101 585
R2198 GND.n4282 GND.n3944 585
R2199 GND.n4278 GND.n3943 585
R2200 GND.n4537 GND.n3943 585
R2201 GND.n4277 GND.n3932 585
R2202 GND.n4544 GND.n3932 585
R2203 GND.n4276 GND.n4275 585
R2204 GND.n4275 GND.n4274 585
R2205 GND.n3202 GND.n3201 585
R2206 GND.n3816 GND.n3202 585
R2207 GND.n4702 GND.n4701 585
R2208 GND.n4701 GND.n4700 585
R2209 GND.n4703 GND.n3196 585
R2210 GND.t180 GND.n3196 585
R2211 GND.n4705 GND.n4704 585
R2212 GND.n4706 GND.n4705 585
R2213 GND.n3182 GND.n3181 585
R2214 GND.n3729 GND.n3182 585
R2215 GND.n4716 GND.n4715 585
R2216 GND.n4715 GND.n4714 585
R2217 GND.n4717 GND.n3176 585
R2218 GND.n3735 GND.n3176 585
R2219 GND.n4719 GND.n4718 585
R2220 GND.n4720 GND.n4719 585
R2221 GND.n3162 GND.n3161 585
R2222 GND.n3708 GND.n3162 585
R2223 GND.n4730 GND.n4729 585
R2224 GND.n4729 GND.n4728 585
R2225 GND.n4731 GND.n3151 585
R2226 GND.n3699 GND.n3151 585
R2227 GND.n4733 GND.n4732 585
R2228 GND.n4734 GND.n4733 585
R2229 GND.n3152 GND.n3150 585
R2230 GND.n3684 GND.n3150 585
R2231 GND.n3155 GND.n3154 585
R2232 GND.n3154 GND.n3131 585
R2233 GND.n3119 GND.n3118 585
R2234 GND.n3129 GND.n3119 585
R2235 GND.n4751 GND.n4750 585
R2236 GND.n4750 GND.n4749 585
R2237 GND.n4752 GND.n3108 585
R2238 GND.n3673 GND.n3108 585
R2239 GND.n4754 GND.n4753 585
R2240 GND.n4755 GND.n4754 585
R2241 GND.n3109 GND.n3107 585
R2242 GND.n3107 GND.n3097 585
R2243 GND.n3112 GND.n3111 585
R2244 GND.n3111 GND.n3095 585
R2245 GND.n3078 GND.n3077 585
R2246 GND.n3372 GND.n3078 585
R2247 GND.n4771 GND.n4770 585
R2248 GND.n4770 GND.n4769 585
R2249 GND.n4772 GND.n3064 585
R2250 GND.n3375 GND.n3064 585
R2251 GND.n4774 GND.n4773 585
R2252 GND.n4775 GND.n4774 585
R2253 GND.n3065 GND.n3063 585
R2254 GND.n3063 GND.n3053 585
R2255 GND.n3071 GND.n3070 585
R2256 GND.n3070 GND.n3051 585
R2257 GND.n3069 GND.n3068 585
R2258 GND.n3069 GND.n3037 585
R2259 GND.n3025 GND.n3024 585
R2260 GND.n3035 GND.n3025 585
R2261 GND.n4799 GND.n4798 585
R2262 GND.n4798 GND.n4797 585
R2263 GND.n4800 GND.n3010 585
R2264 GND.n3615 GND.n3010 585
R2265 GND.n4802 GND.n4801 585
R2266 GND.n4803 GND.n4802 585
R2267 GND.n3011 GND.n3009 585
R2268 GND.n3576 GND.n3009 585
R2269 GND.n3018 GND.n3017 585
R2270 GND.n3017 GND.n2997 585
R2271 GND.n3016 GND.n3015 585
R2272 GND.n3016 GND.n2995 585
R2273 GND.n3014 GND.n2966 585
R2274 GND.n4817 GND.n2966 585
R2275 GND.n4850 GND.n4849 585
R2276 GND.n4848 GND.n2965 585
R2277 GND.n4847 GND.n2964 585
R2278 GND.n4852 GND.n2964 585
R2279 GND.n4846 GND.n4845 585
R2280 GND.n4844 GND.n4843 585
R2281 GND.n4842 GND.n4841 585
R2282 GND.n4840 GND.n4839 585
R2283 GND.n4838 GND.n4837 585
R2284 GND.n4836 GND.n4835 585
R2285 GND.n4834 GND.n4833 585
R2286 GND.n4832 GND.n4831 585
R2287 GND.n4830 GND.n4829 585
R2288 GND.n4827 GND.n4826 585
R2289 GND.n4825 GND.n4824 585
R2290 GND.n4823 GND.n2983 585
R2291 GND.n2984 GND.n2963 585
R2292 GND.n4852 GND.n2963 585
R2293 GND.n3811 GND.n3313 585
R2294 GND.n3810 GND.n3809 585
R2295 GND.n3807 GND.n3755 585
R2296 GND.n3805 GND.n3804 585
R2297 GND.n3800 GND.n3756 585
R2298 GND.n3799 GND.n3798 585
R2299 GND.n3796 GND.n3761 585
R2300 GND.n3794 GND.n3793 585
R2301 GND.n3763 GND.n3762 585
R2302 GND.n3788 GND.n3787 585
R2303 GND.n3785 GND.n3765 585
R2304 GND.n3783 GND.n3782 585
R2305 GND.n3767 GND.n3766 585
R2306 GND.n3778 GND.n3777 585
R2307 GND.n3775 GND.n3769 585
R2308 GND.n3773 GND.n3772 585
R2309 GND.n3815 GND.n3814 585
R2310 GND.n3816 GND.n3815 585
R2311 GND.n3314 GND.n3204 585
R2312 GND.n4700 GND.n3204 585
R2313 GND.n3751 GND.n3750 585
R2314 GND.n3750 GND.t180 585
R2315 GND.n3316 GND.n3194 585
R2316 GND.n4706 GND.n3194 585
R2317 GND.n3731 GND.n3730 585
R2318 GND.n3730 GND.n3729 585
R2319 GND.n3732 GND.n3184 585
R2320 GND.n4714 GND.n3184 585
R2321 GND.n3734 GND.n3733 585
R2322 GND.n3735 GND.n3734 585
R2323 GND.n3345 GND.n3174 585
R2324 GND.n4720 GND.n3174 585
R2325 GND.n3707 GND.n3706 585
R2326 GND.n3708 GND.n3707 585
R2327 GND.n3351 GND.n3164 585
R2328 GND.n4728 GND.n3164 585
R2329 GND.n3701 GND.n3700 585
R2330 GND.n3700 GND.n3699 585
R2331 GND.n3353 GND.n3149 585
R2332 GND.n4734 GND.n3149 585
R2333 GND.n3683 GND.n3682 585
R2334 GND.n3684 GND.n3683 585
R2335 GND.n3364 GND.n3363 585
R2336 GND.n3363 GND.n3131 585
R2337 GND.n3678 GND.n3677 585
R2338 GND.n3677 GND.n3129 585
R2339 GND.n3676 GND.n3121 585
R2340 GND.n4749 GND.n3121 585
R2341 GND.n3675 GND.n3674 585
R2342 GND.n3674 GND.n3673 585
R2343 GND.n3366 GND.n3105 585
R2344 GND.n4755 GND.n3105 585
R2345 GND.n3598 GND.n3597 585
R2346 GND.n3598 GND.n3097 585
R2347 GND.n3599 GND.n3593 585
R2348 GND.n3599 GND.n3095 585
R2349 GND.n3601 GND.n3600 585
R2350 GND.n3600 GND.n3372 585
R2351 GND.n3602 GND.n3080 585
R2352 GND.n4769 GND.n3080 585
R2353 GND.n3604 GND.n3603 585
R2354 GND.n3603 GND.n3375 585
R2355 GND.n3605 GND.n3061 585
R2356 GND.n4775 GND.n3061 585
R2357 GND.n3606 GND.n3585 585
R2358 GND.n3585 GND.n3053 585
R2359 GND.n3608 GND.n3607 585
R2360 GND.n3608 GND.n3051 585
R2361 GND.n3609 GND.n3584 585
R2362 GND.n3609 GND.n3037 585
R2363 GND.n3611 GND.n3610 585
R2364 GND.n3610 GND.n3035 585
R2365 GND.n3612 GND.n3027 585
R2366 GND.n4797 GND.n3027 585
R2367 GND.n3614 GND.n3613 585
R2368 GND.n3615 GND.n3614 585
R2369 GND.n3383 GND.n3007 585
R2370 GND.n4803 GND.n3007 585
R2371 GND.n3578 GND.n3577 585
R2372 GND.n3577 GND.n3576 585
R2373 GND.n3386 GND.n3385 585
R2374 GND.n3386 GND.n2997 585
R2375 GND.n2987 GND.n2986 585
R2376 GND.n2995 GND.n2987 585
R2377 GND.n4819 GND.n4818 585
R2378 GND.n4818 GND.n4817 585
R2379 GND.n4669 GND.n4668 585
R2380 GND.n4670 GND.n4669 585
R2381 GND.n3247 GND.n3245 585
R2382 GND.n3245 GND.n3242 585
R2383 GND.n3841 GND.n3840 585
R2384 GND.n3842 GND.n3841 585
R2385 GND.n3231 GND.n3230 585
R2386 GND.n3234 GND.n3231 585
R2387 GND.n4680 GND.n4679 585
R2388 GND.n4679 GND.n4678 585
R2389 GND.n4681 GND.n3228 585
R2390 GND.n3232 GND.n3228 585
R2391 GND.n4683 GND.n4682 585
R2392 GND.n4684 GND.n4683 585
R2393 GND.n3229 GND.n3227 585
R2394 GND.n3227 GND.n3224 585
R2395 GND.n3828 GND.n3827 585
R2396 GND.n3829 GND.n3828 585
R2397 GND.n3826 GND.n3825 585
R2398 GND.n3825 GND.n3824 585
R2399 GND.n3211 GND.n3210 585
R2400 GND.n4692 GND.n3211 585
R2401 GND.n4695 GND.n4694 585
R2402 GND.n4694 GND.n4693 585
R2403 GND.n4696 GND.n3208 585
R2404 GND.n3816 GND.n3208 585
R2405 GND.n4698 GND.n4697 585
R2406 GND.n4699 GND.n4698 585
R2407 GND.n3209 GND.n3207 585
R2408 GND.n3207 GND.n3203 585
R2409 GND.n3318 GND.n3317 585
R2410 GND.n3319 GND.n3318 585
R2411 GND.n3191 GND.n3190 585
R2412 GND.n3195 GND.n3191 585
R2413 GND.n4709 GND.n4708 585
R2414 GND.n4708 GND.n4707 585
R2415 GND.n4710 GND.n3188 585
R2416 GND.n3728 GND.n3188 585
R2417 GND.n4712 GND.n4711 585
R2418 GND.n4713 GND.n4712 585
R2419 GND.n3189 GND.n3187 585
R2420 GND.n3187 GND.n3183 585
R2421 GND.n3343 GND.n3342 585
R2422 GND.n3344 GND.n3343 585
R2423 GND.n3171 GND.n3170 585
R2424 GND.n3175 GND.n3171 585
R2425 GND.n4723 GND.n4722 585
R2426 GND.n4722 GND.n4721 585
R2427 GND.n4724 GND.n3168 585
R2428 GND.n3709 GND.n3168 585
R2429 GND.n4726 GND.n4725 585
R2430 GND.n4727 GND.n4726 585
R2431 GND.n3169 GND.n3167 585
R2432 GND.n3698 GND.n3167 585
R2433 GND.n3689 GND.n3360 585
R2434 GND.n3360 GND.n3354 585
R2435 GND.n3691 GND.n3690 585
R2436 GND.n3692 GND.n3691 585
R2437 GND.n3688 GND.n3359 585
R2438 GND.n3359 GND.n3148 585
R2439 GND.n3687 GND.n3686 585
R2440 GND.n3686 GND.n3685 585
R2441 GND.n3128 GND.n3127 585
R2442 GND.n3662 GND.n3128 585
R2443 GND.n4744 GND.n4743 585
R2444 GND.n4743 GND.n4742 585
R2445 GND.n4745 GND.n3125 585
R2446 GND.n3666 GND.n3125 585
R2447 GND.n4747 GND.n4746 585
R2448 GND.n4748 GND.n4747 585
R2449 GND.n3126 GND.n3124 585
R2450 GND.n3672 GND.n3124 585
R2451 GND.n3102 GND.n3101 585
R2452 GND.n3368 GND.n3102 585
R2453 GND.n4757 GND.n4756 585
R2454 GND.n4756 GND.n4755 585
R2455 GND.n4758 GND.n3099 585
R2456 GND.n3656 GND.n3099 585
R2457 GND.n4760 GND.n4759 585
R2458 GND.n4761 GND.n4760 585
R2459 GND.n3100 GND.n3098 585
R2460 GND.n3652 GND.n3098 585
R2461 GND.n3649 GND.n3648 585
R2462 GND.n3650 GND.n3649 585
R2463 GND.n3647 GND.n3373 585
R2464 GND.n3373 GND.n3081 585
R2465 GND.n3646 GND.n3645 585
R2466 GND.n3645 GND.n3079 585
R2467 GND.n3644 GND.n3374 585
R2468 GND.n3644 GND.n3643 585
R2469 GND.n3058 GND.n3057 585
R2470 GND.n3376 GND.n3058 585
R2471 GND.n4778 GND.n4777 585
R2472 GND.n4777 GND.n4776 585
R2473 GND.n4779 GND.n3055 585
R2474 GND.n3632 GND.n3055 585
R2475 GND.n4781 GND.n4780 585
R2476 GND.n4782 GND.n4781 585
R2477 GND.n3056 GND.n3054 585
R2478 GND.n3628 GND.n3054 585
R2479 GND.n3034 GND.n3033 585
R2480 GND.n3626 GND.n3034 585
R2481 GND.n4792 GND.n4791 585
R2482 GND.n4791 GND.n4790 585
R2483 GND.n4793 GND.n3031 585
R2484 GND.n3620 GND.n3031 585
R2485 GND.n4795 GND.n4794 585
R2486 GND.n4796 GND.n4795 585
R2487 GND.n3032 GND.n3030 585
R2488 GND.n3616 GND.n3030 585
R2489 GND.n3569 GND.n3568 585
R2490 GND.n3569 GND.n3382 585
R2491 GND.n3571 GND.n3570 585
R2492 GND.n3570 GND.n3008 585
R2493 GND.n3572 GND.n3567 585
R2494 GND.n3567 GND.n3006 585
R2495 GND.n3574 GND.n3573 585
R2496 GND.n3575 GND.n3574 585
R2497 GND.n2994 GND.n2993 585
R2498 GND.n3388 GND.n2994 585
R2499 GND.n4813 GND.n4812 585
R2500 GND.n4812 GND.n4811 585
R2501 GND.n4814 GND.n2991 585
R2502 GND.n3557 GND.n2991 585
R2503 GND.n4816 GND.n4815 585
R2504 GND.n4817 GND.n4816 585
R2505 GND.n2992 GND.n2990 585
R2506 GND.n3553 GND.n2990 585
R2507 GND.n2954 GND.n2953 585
R2508 GND.n3542 GND.n2954 585
R2509 GND.n4855 GND.n4854 585
R2510 GND.n4854 GND.n4853 585
R2511 GND.n4856 GND.n2951 585
R2512 GND.n2951 GND.n2949 585
R2513 GND.n4858 GND.n4857 585
R2514 GND.n4859 GND.n4858 585
R2515 GND.n2952 GND.n2950 585
R2516 GND.n2950 GND.n2947 585
R2517 GND.n3531 GND.n3530 585
R2518 GND.n3532 GND.n3531 585
R2519 GND.n2936 GND.n2935 585
R2520 GND.n2939 GND.n2936 585
R2521 GND.n4868 GND.n4867 585
R2522 GND.n4867 GND.n4866 585
R2523 GND.n4869 GND.n2933 585
R2524 GND.n3523 GND.n2933 585
R2525 GND.n4871 GND.n4870 585
R2526 GND.n4872 GND.n4871 585
R2527 GND.n2934 GND.n2932 585
R2528 GND.n2932 GND.n2930 585
R2529 GND.n3451 GND.n3450 585
R2530 GND.n3454 GND.n3453 585
R2531 GND.n3455 GND.n3415 585
R2532 GND.n3415 GND.n2921 585
R2533 GND.n3457 GND.n3456 585
R2534 GND.n3459 GND.n3414 585
R2535 GND.n3462 GND.n3461 585
R2536 GND.n3463 GND.n3413 585
R2537 GND.n3465 GND.n3464 585
R2538 GND.n3467 GND.n3412 585
R2539 GND.n3470 GND.n3469 585
R2540 GND.n3471 GND.n3411 585
R2541 GND.n3473 GND.n3472 585
R2542 GND.n3475 GND.n3410 585
R2543 GND.n3478 GND.n3477 585
R2544 GND.n3479 GND.n3406 585
R2545 GND.n3481 GND.n3480 585
R2546 GND.n3483 GND.n3405 585
R2547 GND.n3484 GND.n3404 585
R2548 GND.n3486 GND.n3404 585
R2549 GND.n3489 GND.n3488 585
R2550 GND.n3490 GND.n3403 585
R2551 GND.n3492 GND.n3491 585
R2552 GND.n3494 GND.n3402 585
R2553 GND.n3497 GND.n3496 585
R2554 GND.n3498 GND.n3398 585
R2555 GND.n3500 GND.n3499 585
R2556 GND.n3502 GND.n3397 585
R2557 GND.n3505 GND.n3504 585
R2558 GND.n3506 GND.n3396 585
R2559 GND.n3508 GND.n3507 585
R2560 GND.n3510 GND.n3395 585
R2561 GND.n3513 GND.n3512 585
R2562 GND.n3514 GND.n3394 585
R2563 GND.n3516 GND.n3515 585
R2564 GND.n3518 GND.n3393 585
R2565 GND.n3519 GND.n3392 585
R2566 GND.n3519 GND.n2921 585
R2567 GND.n3849 GND.n3848 585
R2568 GND.n3850 GND.n3309 585
R2569 GND.n3852 GND.n3851 585
R2570 GND.n3854 GND.n3307 585
R2571 GND.n3856 GND.n3855 585
R2572 GND.n3857 GND.n3306 585
R2573 GND.n3859 GND.n3858 585
R2574 GND.n3861 GND.n3304 585
R2575 GND.n3863 GND.n3862 585
R2576 GND.n3864 GND.n3303 585
R2577 GND.n3866 GND.n3865 585
R2578 GND.n3868 GND.n3301 585
R2579 GND.n3870 GND.n3869 585
R2580 GND.n3872 GND.n3298 585
R2581 GND.n3874 GND.n3873 585
R2582 GND.n3876 GND.n3297 585
R2583 GND.n3877 GND.n3295 585
R2584 GND.n4637 GND.n3294 585
R2585 GND.n4639 GND.n4638 585
R2586 GND.n4641 GND.n3292 585
R2587 GND.n4643 GND.n4642 585
R2588 GND.n4645 GND.n3289 585
R2589 GND.n4647 GND.n4646 585
R2590 GND.n4649 GND.n3287 585
R2591 GND.n4651 GND.n4650 585
R2592 GND.n4652 GND.n3286 585
R2593 GND.n4654 GND.n4653 585
R2594 GND.n4656 GND.n3284 585
R2595 GND.n4658 GND.n4657 585
R2596 GND.n4659 GND.n3283 585
R2597 GND.n4661 GND.n4660 585
R2598 GND.n4663 GND.n3280 585
R2599 GND.n4665 GND.n4664 585
R2600 GND.n4666 GND.n3246 585
R2601 GND.n3846 GND.n3243 585
R2602 GND.n4670 GND.n3243 585
R2603 GND.n3845 GND.n3844 585
R2604 GND.n3844 GND.n3242 585
R2605 GND.n3843 GND.n3310 585
R2606 GND.n3843 GND.n3842 585
R2607 GND.n3838 GND.n3837 585
R2608 GND.n3838 GND.n3234 585
R2609 GND.n3836 GND.n3233 585
R2610 GND.n4678 GND.n3233 585
R2611 GND.n3835 GND.n3834 585
R2612 GND.n3834 GND.n3232 585
R2613 GND.n3833 GND.n3225 585
R2614 GND.n4684 GND.n3225 585
R2615 GND.n3832 GND.n3831 585
R2616 GND.n3831 GND.n3224 585
R2617 GND.n3830 GND.n3311 585
R2618 GND.n3830 GND.n3829 585
R2619 GND.n3822 GND.n3821 585
R2620 GND.n3824 GND.n3822 585
R2621 GND.n3820 GND.n3214 585
R2622 GND.n4692 GND.n3214 585
R2623 GND.n3819 GND.n3213 585
R2624 GND.n4693 GND.n3213 585
R2625 GND.n3818 GND.n3817 585
R2626 GND.n3817 GND.n3816 585
R2627 GND.n3312 GND.n3205 585
R2628 GND.n4699 GND.n3205 585
R2629 GND.n3721 GND.n3720 585
R2630 GND.n3721 GND.n3203 585
R2631 GND.n3722 GND.n3719 585
R2632 GND.n3722 GND.n3319 585
R2633 GND.n3724 GND.n3723 585
R2634 GND.n3723 GND.n3195 585
R2635 GND.n3725 GND.n3193 585
R2636 GND.n4707 GND.n3193 585
R2637 GND.n3727 GND.n3726 585
R2638 GND.n3728 GND.n3727 585
R2639 GND.n3718 GND.n3185 585
R2640 GND.n4713 GND.n3185 585
R2641 GND.n3717 GND.n3716 585
R2642 GND.n3716 GND.n3183 585
R2643 GND.n3715 GND.n3349 585
R2644 GND.n3715 GND.n3344 585
R2645 GND.n3714 GND.n3713 585
R2646 GND.n3714 GND.n3175 585
R2647 GND.n3712 GND.n3173 585
R2648 GND.n4721 GND.n3173 585
R2649 GND.n3711 GND.n3710 585
R2650 GND.n3710 GND.n3709 585
R2651 GND.n3350 GND.n3165 585
R2652 GND.n4727 GND.n3165 585
R2653 GND.n3697 GND.n3696 585
R2654 GND.n3698 GND.n3697 585
R2655 GND.n3695 GND.n3355 585
R2656 GND.n3355 GND.n3354 585
R2657 GND.n3694 GND.n3693 585
R2658 GND.n3693 GND.n3692 585
R2659 GND.n3357 GND.n3356 585
R2660 GND.n3357 GND.n3148 585
R2661 GND.n3661 GND.n3362 585
R2662 GND.n3685 GND.n3362 585
R2663 GND.n3664 GND.n3663 585
R2664 GND.n3663 GND.n3662 585
R2665 GND.n3665 GND.n3130 585
R2666 GND.n4742 GND.n3130 585
R2667 GND.n3668 GND.n3667 585
R2668 GND.n3667 GND.n3666 585
R2669 GND.n3669 GND.n3122 585
R2670 GND.n4748 GND.n3122 585
R2671 GND.n3671 GND.n3670 585
R2672 GND.n3672 GND.n3671 585
R2673 GND.n3660 GND.n3369 585
R2674 GND.n3369 GND.n3368 585
R2675 GND.n3659 GND.n3104 585
R2676 GND.n4755 GND.n3104 585
R2677 GND.n3658 GND.n3657 585
R2678 GND.n3657 GND.n3656 585
R2679 GND.n3655 GND.n3096 585
R2680 GND.n4761 GND.n3096 585
R2681 GND.n3654 GND.n3653 585
R2682 GND.n3653 GND.n3652 585
R2683 GND.n3371 GND.n3370 585
R2684 GND.n3650 GND.n3371 585
R2685 GND.n3638 GND.n3637 585
R2686 GND.n3637 GND.n3081 585
R2687 GND.n3639 GND.n3378 585
R2688 GND.n3378 GND.n3079 585
R2689 GND.n3641 GND.n3640 585
R2690 GND.n3643 GND.n3641 585
R2691 GND.n3636 GND.n3377 585
R2692 GND.n3377 GND.n3376 585
R2693 GND.n3635 GND.n3060 585
R2694 GND.n4776 GND.n3060 585
R2695 GND.n3634 GND.n3633 585
R2696 GND.n3633 GND.n3632 585
R2697 GND.n3631 GND.n3052 585
R2698 GND.n4782 GND.n3052 585
R2699 GND.n3630 GND.n3629 585
R2700 GND.n3629 GND.n3628 585
R2701 GND.n3625 GND.n3624 585
R2702 GND.n3626 GND.n3625 585
R2703 GND.n3623 GND.n3036 585
R2704 GND.n4790 GND.n3036 585
R2705 GND.n3622 GND.n3621 585
R2706 GND.n3621 GND.n3620 585
R2707 GND.n3619 GND.n3028 585
R2708 GND.n4796 GND.n3028 585
R2709 GND.n3618 GND.n3617 585
R2710 GND.n3617 GND.n3616 585
R2711 GND.n3380 GND.n3379 585
R2712 GND.n3382 GND.n3380 585
R2713 GND.n3563 GND.n3562 585
R2714 GND.n3562 GND.n3008 585
R2715 GND.n3564 GND.n3390 585
R2716 GND.n3390 GND.n3006 585
R2717 GND.n3566 GND.n3565 585
R2718 GND.n3575 GND.n3566 585
R2719 GND.n3561 GND.n3389 585
R2720 GND.n3389 GND.n3388 585
R2721 GND.n3560 GND.n2996 585
R2722 GND.n4811 GND.n2996 585
R2723 GND.n3559 GND.n3558 585
R2724 GND.n3558 GND.n3557 585
R2725 GND.n3556 GND.n2988 585
R2726 GND.n4817 GND.n2988 585
R2727 GND.n3555 GND.n3554 585
R2728 GND.n3554 GND.n3553 585
R2729 GND.n3541 GND.n3540 585
R2730 GND.n3542 GND.n3541 585
R2731 GND.n3539 GND.n2956 585
R2732 GND.n4853 GND.n2956 585
R2733 GND.n3538 GND.n3537 585
R2734 GND.n3537 GND.n2949 585
R2735 GND.n3536 GND.n2948 585
R2736 GND.n4859 GND.n2948 585
R2737 GND.n3535 GND.n3534 585
R2738 GND.n3534 GND.n2947 585
R2739 GND.n3533 GND.n3391 585
R2740 GND.n3533 GND.n3532 585
R2741 GND.n3528 GND.n3527 585
R2742 GND.n3528 GND.n2939 585
R2743 GND.n3526 GND.n2938 585
R2744 GND.n4866 GND.n2938 585
R2745 GND.n3525 GND.n3524 585
R2746 GND.n3524 GND.n3523 585
R2747 GND.n3522 GND.n2931 585
R2748 GND.n4872 GND.n2931 585
R2749 GND.n3521 GND.n3520 585
R2750 GND.n3520 GND.n2930 585
R2751 GND.n5055 GND.n5054 585
R2752 GND.n5056 GND.n5055 585
R2753 GND.n1992 GND.n1990 585
R2754 GND.n2908 GND.n1990 585
R2755 GND.n2901 GND.n2073 585
R2756 GND.n2073 GND.n2066 585
R2757 GND.n2903 GND.n2902 585
R2758 GND.n2904 GND.n2903 585
R2759 GND.n2074 GND.n2072 585
R2760 GND.n2837 GND.n2072 585
R2761 GND.n2896 GND.n2895 585
R2762 GND.n2895 GND.n2894 585
R2763 GND.n2077 GND.n2076 585
R2764 GND.n2891 GND.n2077 585
R2765 GND.n2821 GND.n2820 585
R2766 GND.n2822 GND.n2821 585
R2767 GND.n2098 GND.n2097 585
R2768 GND.n2097 GND.n2096 585
R2769 GND.n2816 GND.n2815 585
R2770 GND.n2815 GND.n2814 585
R2771 GND.n2101 GND.n2100 585
R2772 GND.n2810 GND.n2101 585
R2773 GND.n2795 GND.n2118 585
R2774 GND.n2711 GND.n2118 585
R2775 GND.n2797 GND.n2796 585
R2776 GND.n2798 GND.n2797 585
R2777 GND.n2119 GND.n2117 585
R2778 GND.n2785 GND.n2117 585
R2779 GND.n2790 GND.n2789 585
R2780 GND.n2789 GND.n2788 585
R2781 GND.n2122 GND.n2121 585
R2782 GND.n2782 GND.n2122 585
R2783 GND.n2770 GND.n2139 585
R2784 GND.n2731 GND.n2139 585
R2785 GND.n2772 GND.n2771 585
R2786 GND.n2773 GND.n2772 585
R2787 GND.n2140 GND.n2138 585
R2788 GND.n2698 GND.n2138 585
R2789 GND.n2694 GND.n2693 585
R2790 GND.n2695 GND.n2694 585
R2791 GND.n2176 GND.n2175 585
R2792 GND.n2742 GND.n2175 585
R2793 GND.n2746 GND.n2177 585
R2794 GND.n2746 GND.n2745 585
R2795 GND.n2749 GND.n2748 585
R2796 GND.n2750 GND.n2749 585
R2797 GND.n2747 GND.n2174 585
R2798 GND.n2174 GND.n2165 585
R2799 GND.n2173 GND.n2172 585
R2800 GND.n2173 GND.n2158 585
R2801 GND.n2171 GND.n2149 585
R2802 GND.n2759 GND.n2149 585
R2803 GND.n2764 GND.n2763 585
R2804 GND.n2763 GND.n2762 585
R2805 GND.n2765 GND.n2148 585
R2806 GND.n2652 GND.n2148 585
R2807 GND.n2201 GND.n2147 585
R2808 GND.n2651 GND.n2201 585
R2809 GND.n2672 GND.n2671 585
R2810 GND.n2673 GND.n2672 585
R2811 GND.n2670 GND.n2200 585
R2812 GND.n2214 GND.n2200 585
R2813 GND.n2206 GND.n2202 585
R2814 GND.n2661 GND.n2206 585
R2815 GND.n2666 GND.n2665 585
R2816 GND.n2665 GND.n2664 585
R2817 GND.n2205 GND.n2204 585
R2818 GND.n2635 GND.n2205 585
R2819 GND.n2621 GND.n2235 585
R2820 GND.n2235 GND.n2221 585
R2821 GND.n2623 GND.n2622 585
R2822 GND.n2624 GND.n2623 585
R2823 GND.n2236 GND.n2234 585
R2824 GND.n2611 GND.n2234 585
R2825 GND.n2616 GND.n2615 585
R2826 GND.n2615 GND.n2614 585
R2827 GND.n2239 GND.n2238 585
R2828 GND.n2609 GND.n2239 585
R2829 GND.n2597 GND.n2258 585
R2830 GND.n2258 GND.n2257 585
R2831 GND.n2599 GND.n2598 585
R2832 GND.n2600 GND.n2599 585
R2833 GND.n2259 GND.n2256 585
R2834 GND.n2587 GND.n2256 585
R2835 GND.n2592 GND.n2591 585
R2836 GND.n2591 GND.n2590 585
R2837 GND.n1885 GND.n1884 585
R2838 GND.n2262 GND.n1885 585
R2839 GND.n5130 GND.n5129 585
R2840 GND.n5129 GND.n5128 585
R2841 GND.n5131 GND.n1880 585
R2842 GND.n2540 GND.n1880 585
R2843 GND.n5133 GND.n5132 585
R2844 GND.n5134 GND.n5133 585
R2845 GND.n2343 GND.n1879 585
R2846 GND.n2342 GND.n2341 585
R2847 GND.n2348 GND.n2347 585
R2848 GND.n2350 GND.n2339 585
R2849 GND.n2353 GND.n2352 585
R2850 GND.n2337 GND.n2336 585
R2851 GND.n2358 GND.n2357 585
R2852 GND.n2360 GND.n2335 585
R2853 GND.n2363 GND.n2362 585
R2854 GND.n2333 GND.n2332 585
R2855 GND.n2370 GND.n2369 585
R2856 GND.n2372 GND.n2331 585
R2857 GND.n2375 GND.n2374 585
R2858 GND.n2329 GND.n2328 585
R2859 GND.n2380 GND.n2379 585
R2860 GND.n2382 GND.n2327 585
R2861 GND.n2385 GND.n2384 585
R2862 GND.n2325 GND.n2324 585
R2863 GND.n2390 GND.n2389 585
R2864 GND.n2392 GND.n2323 585
R2865 GND.n2395 GND.n2394 585
R2866 GND.n2321 GND.n2320 585
R2867 GND.n2402 GND.n2401 585
R2868 GND.n2404 GND.n2319 585
R2869 GND.n2407 GND.n2406 585
R2870 GND.n2317 GND.n2316 585
R2871 GND.n2412 GND.n2411 585
R2872 GND.n2414 GND.n2315 585
R2873 GND.n2417 GND.n2416 585
R2874 GND.n2313 GND.n2312 585
R2875 GND.n2422 GND.n2421 585
R2876 GND.n2424 GND.n2311 585
R2877 GND.n2427 GND.n2426 585
R2878 GND.n2309 GND.n2308 585
R2879 GND.n2435 GND.n2434 585
R2880 GND.n2437 GND.n2307 585
R2881 GND.n2440 GND.n2439 585
R2882 GND.n2305 GND.n2304 585
R2883 GND.n2445 GND.n2444 585
R2884 GND.n2447 GND.n2303 585
R2885 GND.n2450 GND.n2449 585
R2886 GND.n2301 GND.n2300 585
R2887 GND.n2455 GND.n2454 585
R2888 GND.n2457 GND.n2299 585
R2889 GND.n2460 GND.n2459 585
R2890 GND.n2297 GND.n2296 585
R2891 GND.n2468 GND.n2467 585
R2892 GND.n2470 GND.n2295 585
R2893 GND.n2473 GND.n2472 585
R2894 GND.n2293 GND.n2292 585
R2895 GND.n2478 GND.n2477 585
R2896 GND.n2480 GND.n2291 585
R2897 GND.n2483 GND.n2482 585
R2898 GND.n2289 GND.n2288 585
R2899 GND.n2488 GND.n2487 585
R2900 GND.n2490 GND.n2287 585
R2901 GND.n2493 GND.n2492 585
R2902 GND.n2285 GND.n2284 585
R2903 GND.n2498 GND.n2497 585
R2904 GND.n2500 GND.n2283 585
R2905 GND.n2502 GND.n2501 585
R2906 GND.n2501 GND.n1874 585
R2907 GND.n4959 GND.n1985 585
R2908 GND.n4960 GND.n4958 585
R2909 GND.n4956 GND.n4951 585
R2910 GND.n4964 GND.n4950 585
R2911 GND.n4965 GND.n4949 585
R2912 GND.n4966 GND.n4947 585
R2913 GND.n4946 GND.n4943 585
R2914 GND.n4970 GND.n4942 585
R2915 GND.n4971 GND.n4941 585
R2916 GND.n4972 GND.n4939 585
R2917 GND.n4938 GND.n4935 585
R2918 GND.n4976 GND.n4934 585
R2919 GND.n4977 GND.n4933 585
R2920 GND.n4978 GND.n4931 585
R2921 GND.n4930 GND.n4924 585
R2922 GND.n4982 GND.n4923 585
R2923 GND.n4983 GND.n4922 585
R2924 GND.n4984 GND.n4920 585
R2925 GND.n4919 GND.n4916 585
R2926 GND.n4988 GND.n4915 585
R2927 GND.n4989 GND.n4914 585
R2928 GND.n4990 GND.n4912 585
R2929 GND.n4911 GND.n4908 585
R2930 GND.n4994 GND.n4907 585
R2931 GND.n4995 GND.n4906 585
R2932 GND.n4996 GND.n4904 585
R2933 GND.n4999 GND.n4899 585
R2934 GND.n5000 GND.n4897 585
R2935 GND.n5001 GND.n4896 585
R2936 GND.n4891 GND.n4890 585
R2937 GND.n5006 GND.n5005 585
R2938 GND.n5008 GND.n4889 585
R2939 GND.n5009 GND.n4888 585
R2940 GND.n5013 GND.n5012 585
R2941 GND.n5014 GND.n2030 585
R2942 GND.n2050 GND.n2028 585
R2943 GND.n5018 GND.n2027 585
R2944 GND.n5019 GND.n2026 585
R2945 GND.n5020 GND.n2023 585
R2946 GND.n2047 GND.n2021 585
R2947 GND.n5024 GND.n2020 585
R2948 GND.n5025 GND.n2019 585
R2949 GND.n5026 GND.n2018 585
R2950 GND.n2044 GND.n2016 585
R2951 GND.n5030 GND.n2015 585
R2952 GND.n5031 GND.n2014 585
R2953 GND.n5032 GND.n2013 585
R2954 GND.n2041 GND.n2011 585
R2955 GND.n5036 GND.n2010 585
R2956 GND.n5037 GND.n2009 585
R2957 GND.n5038 GND.n2005 585
R2958 GND.n5039 GND.n2004 585
R2959 GND.n2037 GND.n2002 585
R2960 GND.n5043 GND.n2001 585
R2961 GND.n5044 GND.n2000 585
R2962 GND.n5045 GND.n1999 585
R2963 GND.n2034 GND.n1997 585
R2964 GND.n5049 GND.n1996 585
R2965 GND.n5050 GND.n1995 585
R2966 GND.n5051 GND.n1991 585
R2967 GND.n5058 GND.n5057 585
R2968 GND.n5057 GND.n5056 585
R2969 GND.n1984 GND.n1979 585
R2970 GND.n2908 GND.n1984 585
R2971 GND.n5062 GND.n1978 585
R2972 GND.n2066 GND.n1978 585
R2973 GND.n5063 GND.n1977 585
R2974 GND.n2904 GND.n1977 585
R2975 GND.n5064 GND.n1976 585
R2976 GND.n2837 GND.n1976 585
R2977 GND.n2079 GND.n1971 585
R2978 GND.n2894 GND.n2079 585
R2979 GND.n5068 GND.n1970 585
R2980 GND.n2891 GND.n1970 585
R2981 GND.n5069 GND.n1969 585
R2982 GND.n2822 GND.n1969 585
R2983 GND.n5070 GND.n1968 585
R2984 GND.n2096 GND.n1968 585
R2985 GND.n2103 GND.n1963 585
R2986 GND.n2814 GND.n2103 585
R2987 GND.n5074 GND.n1962 585
R2988 GND.n2810 GND.n1962 585
R2989 GND.n5075 GND.n1961 585
R2990 GND.n2711 GND.n1961 585
R2991 GND.n5076 GND.n1960 585
R2992 GND.n2798 GND.n1960 585
R2993 GND.n2784 GND.n1955 585
R2994 GND.n2785 GND.n2784 585
R2995 GND.n5080 GND.n1954 585
R2996 GND.n2788 GND.n1954 585
R2997 GND.n5081 GND.n1953 585
R2998 GND.n2782 GND.n1953 585
R2999 GND.n5082 GND.n1952 585
R3000 GND.n2731 GND.n1952 585
R3001 GND.n2135 GND.n1947 585
R3002 GND.n2773 GND.n2135 585
R3003 GND.n5086 GND.n1946 585
R3004 GND.n2698 GND.n1946 585
R3005 GND.n5087 GND.n1945 585
R3006 GND.n2695 GND.n1945 585
R3007 GND.n5088 GND.n1944 585
R3008 GND.n2742 GND.n1944 585
R3009 GND.n2178 GND.n1939 585
R3010 GND.n2745 GND.n2178 585
R3011 GND.n5092 GND.n1938 585
R3012 GND.n2750 GND.n1938 585
R3013 GND.n5093 GND.n1937 585
R3014 GND.n2165 GND.n1937 585
R3015 GND.n5094 GND.n1936 585
R3016 GND.n2158 GND.n1936 585
R3017 GND.n2156 GND.n1931 585
R3018 GND.n2759 GND.n2156 585
R3019 GND.n5098 GND.n1930 585
R3020 GND.n2762 GND.n1930 585
R3021 GND.n5099 GND.n1929 585
R3022 GND.n2652 GND.n1929 585
R3023 GND.n5100 GND.n1928 585
R3024 GND.n2651 GND.n1928 585
R3025 GND.n2197 GND.n1923 585
R3026 GND.n2673 GND.n2197 585
R3027 GND.n5104 GND.n1922 585
R3028 GND.n2214 GND.n1922 585
R3029 GND.n5105 GND.n1921 585
R3030 GND.n2661 GND.n1921 585
R3031 GND.n5106 GND.n1920 585
R3032 GND.n2664 GND.n1920 585
R3033 GND.n2222 GND.n1915 585
R3034 GND.n2635 GND.n2222 585
R3035 GND.n5110 GND.n1914 585
R3036 GND.n2221 GND.n1914 585
R3037 GND.n5111 GND.n1913 585
R3038 GND.n2624 GND.n1913 585
R3039 GND.n5112 GND.n1912 585
R3040 GND.n2611 GND.n1912 585
R3041 GND.n2241 GND.n1907 585
R3042 GND.n2614 GND.n2241 585
R3043 GND.n5116 GND.n1906 585
R3044 GND.n2609 GND.n1906 585
R3045 GND.n5117 GND.n1905 585
R3046 GND.n2257 GND.n1905 585
R3047 GND.n5118 GND.n1904 585
R3048 GND.n2600 GND.n1904 585
R3049 GND.n2586 GND.n1899 585
R3050 GND.n2587 GND.n2586 585
R3051 GND.n5122 GND.n1898 585
R3052 GND.n2590 GND.n1898 585
R3053 GND.n5123 GND.n1897 585
R3054 GND.n2262 GND.n1897 585
R3055 GND.n5124 GND.n1887 585
R3056 GND.n5128 GND.n1887 585
R3057 GND.n2539 GND.n1896 585
R3058 GND.n2540 GND.n2539 585
R3059 GND.n2505 GND.n1875 585
R3060 GND.n5134 GND.n1875 585
R3061 GND.n6792 GND.n6791 585
R3062 GND.n6793 GND.n6792 585
R3063 GND.n634 GND.n633 585
R3064 GND.n6648 GND.n634 585
R3065 GND.n6801 GND.n6800 585
R3066 GND.n6800 GND.n6799 585
R3067 GND.n6802 GND.n628 585
R3068 GND.n6641 GND.n628 585
R3069 GND.n6804 GND.n6803 585
R3070 GND.n6805 GND.n6804 585
R3071 GND.n613 GND.n612 585
R3072 GND.n6632 GND.n613 585
R3073 GND.n6813 GND.n6812 585
R3074 GND.n6812 GND.n6811 585
R3075 GND.n6814 GND.n607 585
R3076 GND.n6626 GND.n607 585
R3077 GND.n6816 GND.n6815 585
R3078 GND.n6817 GND.n6816 585
R3079 GND.n593 GND.n592 585
R3080 GND.n6618 GND.n593 585
R3081 GND.n6825 GND.n6824 585
R3082 GND.n6824 GND.n6823 585
R3083 GND.n6826 GND.n587 585
R3084 GND.n6612 GND.n587 585
R3085 GND.n6828 GND.n6827 585
R3086 GND.n6829 GND.n6828 585
R3087 GND.n572 GND.n571 585
R3088 GND.n4428 GND.n572 585
R3089 GND.n6837 GND.n6836 585
R3090 GND.n6836 GND.n6835 585
R3091 GND.n6838 GND.n567 585
R3092 GND.n4434 GND.n567 585
R3093 GND.n6840 GND.n6839 585
R3094 GND.n6841 GND.n6840 585
R3095 GND.n550 GND.n548 585
R3096 GND.n4440 GND.n550 585
R3097 GND.n6849 GND.n6848 585
R3098 GND.n6848 GND.n6847 585
R3099 GND.n549 GND.n547 585
R3100 GND.n4446 GND.n549 585
R3101 GND.n4455 GND.n4454 585
R3102 GND.n4456 GND.n4455 585
R3103 GND.n4453 GND.n540 585
R3104 GND.n4453 GND.n4452 585
R3105 GND.n6852 GND.n538 585
R3106 GND.n4462 GND.n538 585
R3107 GND.n6854 GND.n6853 585
R3108 GND.n6855 GND.n6854 585
R3109 GND.n4476 GND.n537 585
R3110 GND.n4468 GND.n537 585
R3111 GND.n4478 GND.n4477 585
R3112 GND.n4479 GND.n4478 585
R3113 GND.n4475 GND.n4044 585
R3114 GND.n4475 GND.n4474 585
R3115 GND.n4043 GND.n4030 585
R3116 GND.n4033 GND.n4030 585
R3117 GND.n4490 GND.n4489 585
R3118 GND.n4489 GND.n4488 585
R3119 GND.n4492 GND.n4491 585
R3120 GND.n4493 GND.n4492 585
R3121 GND.n4016 GND.n4015 585
R3122 GND.n4349 GND.n4016 585
R3123 GND.n4501 GND.n4500 585
R3124 GND.n4500 GND.n4499 585
R3125 GND.n4502 GND.n4009 585
R3126 GND.n4330 GND.n4009 585
R3127 GND.n4504 GND.n4503 585
R3128 GND.n4505 GND.n4504 585
R3129 GND.n3994 GND.n3993 585
R3130 GND.n4323 GND.n3994 585
R3131 GND.n4513 GND.n4512 585
R3132 GND.n4512 GND.n4511 585
R3133 GND.n4514 GND.n3988 585
R3134 GND.n4315 GND.n3988 585
R3135 GND.n4516 GND.n4515 585
R3136 GND.n4517 GND.n4516 585
R3137 GND.n3971 GND.n3970 585
R3138 GND.n4308 GND.n3971 585
R3139 GND.n4525 GND.n4524 585
R3140 GND.n4524 GND.n4523 585
R3141 GND.n4526 GND.n3960 585
R3142 GND.n4300 GND.n3960 585
R3143 GND.n4528 GND.n4527 585
R3144 GND.n4529 GND.n4528 585
R3145 GND.n3961 GND.n3959 585
R3146 GND.n3959 GND.n3954 585
R3147 GND.n3964 GND.n3963 585
R3148 GND.n3963 GND.n3944 585
R3149 GND.n3929 GND.n3928 585
R3150 GND.n4537 GND.n3929 585
R3151 GND.n4546 GND.n4545 585
R3152 GND.n4545 GND.n4544 585
R3153 GND.n4547 GND.n3926 585
R3154 GND.n4274 GND.n3926 585
R3155 GND.n4629 GND.n4628 585
R3156 GND.n4627 GND.n3925 585
R3157 GND.n4626 GND.n3924 585
R3158 GND.n4631 GND.n3924 585
R3159 GND.n4625 GND.n4624 585
R3160 GND.n4623 GND.n4622 585
R3161 GND.n4621 GND.n4620 585
R3162 GND.n4619 GND.n4618 585
R3163 GND.n4617 GND.n4616 585
R3164 GND.n4615 GND.n4614 585
R3165 GND.n4613 GND.n4612 585
R3166 GND.n4611 GND.n4559 585
R3167 GND.n4610 GND.n4609 585
R3168 GND.n4608 GND.n4607 585
R3169 GND.n4606 GND.n4605 585
R3170 GND.n4604 GND.n4603 585
R3171 GND.n4602 GND.n4601 585
R3172 GND.n4600 GND.n4599 585
R3173 GND.n4598 GND.n4597 585
R3174 GND.n4596 GND.n4595 585
R3175 GND.n4594 GND.n4593 585
R3176 GND.n4592 GND.n4591 585
R3177 GND.n4590 GND.n4589 585
R3178 GND.n4588 GND.n4574 585
R3179 GND.n4587 GND.n4586 585
R3180 GND.n4585 GND.n4584 585
R3181 GND.n4583 GND.n4582 585
R3182 GND.n3899 GND.n3880 585
R3183 GND.n4635 GND.n3882 585
R3184 GND.n4635 GND.n3881 585
R3185 GND.n4634 GND.n4633 585
R3186 GND.n3886 GND.n3885 585
R3187 GND.n4153 GND.n4152 585
R3188 GND.n4158 GND.n4157 585
R3189 GND.n4160 GND.n4159 585
R3190 GND.n4166 GND.n4165 585
R3191 GND.n4164 GND.n4150 585
R3192 GND.n4171 GND.n4170 585
R3193 GND.n4173 GND.n4172 585
R3194 GND.n4176 GND.n4175 585
R3195 GND.n4174 GND.n4148 585
R3196 GND.n4181 GND.n4180 585
R3197 GND.n4183 GND.n4182 585
R3198 GND.n4186 GND.n4185 585
R3199 GND.n4184 GND.n4146 585
R3200 GND.n4191 GND.n4190 585
R3201 GND.n4193 GND.n4192 585
R3202 GND.n4199 GND.n4198 585
R3203 GND.n4197 GND.n4144 585
R3204 GND.n4204 GND.n4203 585
R3205 GND.n4206 GND.n4205 585
R3206 GND.n4209 GND.n4208 585
R3207 GND.n4207 GND.n4142 585
R3208 GND.n4214 GND.n4213 585
R3209 GND.n4216 GND.n4215 585
R3210 GND.n4219 GND.n4218 585
R3211 GND.n4217 GND.n4140 585
R3212 GND.n4224 GND.n4223 585
R3213 GND.n4226 GND.n4225 585
R3214 GND.n4229 GND.n4228 585
R3215 GND.n4227 GND.n4138 585
R3216 GND.n4272 GND.n4271 585
R3217 GND.n757 GND.n756 585
R3218 GND.n6677 GND.n752 585
R3219 GND.n6679 GND.n6678 585
R3220 GND.n6681 GND.n750 585
R3221 GND.n6683 GND.n6682 585
R3222 GND.n6684 GND.n745 585
R3223 GND.n6686 GND.n6685 585
R3224 GND.n6688 GND.n743 585
R3225 GND.n6690 GND.n6689 585
R3226 GND.n6691 GND.n738 585
R3227 GND.n6693 GND.n6692 585
R3228 GND.n6695 GND.n736 585
R3229 GND.n6697 GND.n6696 585
R3230 GND.n6698 GND.n731 585
R3231 GND.n6703 GND.n6702 585
R3232 GND.n6705 GND.n729 585
R3233 GND.n6707 GND.n6706 585
R3234 GND.n6708 GND.n724 585
R3235 GND.n6710 GND.n6709 585
R3236 GND.n6712 GND.n722 585
R3237 GND.n6714 GND.n6713 585
R3238 GND.n6715 GND.n717 585
R3239 GND.n6717 GND.n6716 585
R3240 GND.n6719 GND.n715 585
R3241 GND.n6721 GND.n6720 585
R3242 GND.n6722 GND.n710 585
R3243 GND.n6727 GND.n6726 585
R3244 GND.n6729 GND.n708 585
R3245 GND.n6731 GND.n6730 585
R3246 GND.n6732 GND.n703 585
R3247 GND.n6734 GND.n6733 585
R3248 GND.n6736 GND.n701 585
R3249 GND.n6738 GND.n6737 585
R3250 GND.n6739 GND.n697 585
R3251 GND.n6741 GND.n6740 585
R3252 GND.n6743 GND.n695 585
R3253 GND.n6745 GND.n6744 585
R3254 GND.n690 GND.n689 585
R3255 GND.n6750 GND.n6749 585
R3256 GND.n6752 GND.n687 585
R3257 GND.n6754 GND.n6753 585
R3258 GND.n6755 GND.n682 585
R3259 GND.n6757 GND.n6756 585
R3260 GND.n6759 GND.n680 585
R3261 GND.n6761 GND.n6760 585
R3262 GND.n6762 GND.n676 585
R3263 GND.n6764 GND.n6763 585
R3264 GND.n6766 GND.n673 585
R3265 GND.n6768 GND.n6767 585
R3266 GND.n674 GND.n667 585
R3267 GND.n6772 GND.n671 585
R3268 GND.n6773 GND.n663 585
R3269 GND.n6775 GND.n6774 585
R3270 GND.n6777 GND.n661 585
R3271 GND.n6779 GND.n6778 585
R3272 GND.n6780 GND.n656 585
R3273 GND.n6782 GND.n6781 585
R3274 GND.n6784 GND.n653 585
R3275 GND.n6786 GND.n6785 585
R3276 GND.n6787 GND.n651 585
R3277 GND.n6788 GND.n648 585
R3278 GND.n655 GND.n648 585
R3279 GND.n6645 GND.n645 585
R3280 GND.n6793 GND.n645 585
R3281 GND.n6647 GND.n6646 585
R3282 GND.n6648 GND.n6647 585
R3283 GND.n6644 GND.n636 585
R3284 GND.n6799 GND.n636 585
R3285 GND.n6643 GND.n6642 585
R3286 GND.n6642 GND.n6641 585
R3287 GND.n784 GND.n625 585
R3288 GND.n6805 GND.n625 585
R3289 GND.n6631 GND.n6630 585
R3290 GND.n6632 GND.n6631 585
R3291 GND.n6629 GND.n615 585
R3292 GND.n6811 GND.n615 585
R3293 GND.n6628 GND.n6627 585
R3294 GND.n6627 GND.n6626 585
R3295 GND.n789 GND.n604 585
R3296 GND.n6817 GND.n604 585
R3297 GND.n6617 GND.n6616 585
R3298 GND.n6618 GND.n6617 585
R3299 GND.n6615 GND.n594 585
R3300 GND.n6823 GND.n594 585
R3301 GND.n6614 GND.n6613 585
R3302 GND.n6613 GND.n6612 585
R3303 GND.n794 GND.n584 585
R3304 GND.n6829 GND.n584 585
R3305 GND.n4430 GND.n4429 585
R3306 GND.n4429 GND.n4428 585
R3307 GND.n4431 GND.n574 585
R3308 GND.n6835 GND.n574 585
R3309 GND.n4433 GND.n4432 585
R3310 GND.n4434 GND.n4433 585
R3311 GND.n4413 GND.n564 585
R3312 GND.n6841 GND.n564 585
R3313 GND.n4442 GND.n4441 585
R3314 GND.n4441 GND.n4440 585
R3315 GND.n4443 GND.n552 585
R3316 GND.n6847 GND.n552 585
R3317 GND.n4445 GND.n4444 585
R3318 GND.n4446 GND.n4445 585
R3319 GND.n4411 GND.n4369 585
R3320 GND.n4456 GND.n4369 585
R3321 GND.n4363 GND.n4362 585
R3322 GND.n4452 GND.n4363 585
R3323 GND.n4464 GND.n4463 585
R3324 GND.n4463 GND.n4462 585
R3325 GND.n4465 GND.n534 585
R3326 GND.n6855 GND.n534 585
R3327 GND.n4467 GND.n4466 585
R3328 GND.n4468 GND.n4467 585
R3329 GND.n4359 GND.n4039 585
R3330 GND.n4479 GND.n4039 585
R3331 GND.n4358 GND.n4046 585
R3332 GND.n4474 GND.n4046 585
R3333 GND.n4357 GND.n4356 585
R3334 GND.n4356 GND.n4033 585
R3335 GND.n4353 GND.n4031 585
R3336 GND.n4488 GND.n4031 585
R3337 GND.n4352 GND.n4027 585
R3338 GND.n4493 GND.n4027 585
R3339 GND.n4351 GND.n4350 585
R3340 GND.n4350 GND.n4349 585
R3341 GND.n4054 GND.n4018 585
R3342 GND.n4499 GND.n4018 585
R3343 GND.n4329 GND.n4328 585
R3344 GND.n4330 GND.n4329 585
R3345 GND.n4326 GND.n4006 585
R3346 GND.n4505 GND.n4006 585
R3347 GND.n4325 GND.n4324 585
R3348 GND.n4324 GND.n4323 585
R3349 GND.n4094 GND.n3996 585
R3350 GND.n4511 GND.n3996 585
R3351 GND.n4314 GND.n4313 585
R3352 GND.n4315 GND.n4314 585
R3353 GND.n4311 GND.n3985 585
R3354 GND.n4517 GND.n3985 585
R3355 GND.n4310 GND.n4309 585
R3356 GND.n4309 GND.n4308 585
R3357 GND.n4098 GND.n3973 585
R3358 GND.n4523 GND.n3973 585
R3359 GND.n4299 GND.n4298 585
R3360 GND.n4300 GND.n4299 585
R3361 GND.n4286 GND.n3955 585
R3362 GND.n4529 GND.n3955 585
R3363 GND.n4288 GND.n4287 585
R3364 GND.n4287 GND.n3954 585
R3365 GND.n3942 GND.n3941 585
R3366 GND.n3944 GND.n3942 585
R3367 GND.n4539 GND.n4538 585
R3368 GND.n4538 GND.n4537 585
R3369 GND.n4540 GND.n3931 585
R3370 GND.n4544 GND.n3931 585
R3371 GND.n4273 GND.n3940 585
R3372 GND.n4274 GND.n4273 585
R3373 GND.n5328 GND.n5327 585
R3374 GND.n5326 GND.n1683 585
R3375 GND.n6402 GND.n6401 585
R3376 GND.n1006 GND.n1005 585
R3377 GND.n6405 GND.n1001 585
R3378 GND.n1001 GND.n1000 585
R3379 GND.n6407 GND.n6406 585
R3380 GND.n6408 GND.n6407 585
R3381 GND.n999 GND.n998 585
R3382 GND.n6409 GND.n999 585
R3383 GND.n6412 GND.n6411 585
R3384 GND.n6411 GND.n6410 585
R3385 GND.n6413 GND.n993 585
R3386 GND.n993 GND.n992 585
R3387 GND.n6415 GND.n6414 585
R3388 GND.n6416 GND.n6415 585
R3389 GND.n991 GND.n990 585
R3390 GND.n6417 GND.n991 585
R3391 GND.n6420 GND.n6419 585
R3392 GND.n6419 GND.n6418 585
R3393 GND.n6421 GND.n985 585
R3394 GND.n985 GND.n984 585
R3395 GND.n6423 GND.n6422 585
R3396 GND.n6424 GND.n6423 585
R3397 GND.n983 GND.n982 585
R3398 GND.n6425 GND.n983 585
R3399 GND.n6428 GND.n6427 585
R3400 GND.n6427 GND.n6426 585
R3401 GND.n6429 GND.n977 585
R3402 GND.n977 GND.n976 585
R3403 GND.n6431 GND.n6430 585
R3404 GND.n6432 GND.n6431 585
R3405 GND.n975 GND.n974 585
R3406 GND.n6433 GND.n975 585
R3407 GND.n6436 GND.n6435 585
R3408 GND.n6435 GND.n6434 585
R3409 GND.n6437 GND.n969 585
R3410 GND.n969 GND.n968 585
R3411 GND.n6439 GND.n6438 585
R3412 GND.n6440 GND.n6439 585
R3413 GND.n967 GND.n966 585
R3414 GND.n6441 GND.n967 585
R3415 GND.n6444 GND.n6443 585
R3416 GND.n6443 GND.n6442 585
R3417 GND.n6445 GND.n961 585
R3418 GND.n961 GND.n960 585
R3419 GND.n6447 GND.n6446 585
R3420 GND.n6448 GND.n6447 585
R3421 GND.n959 GND.n958 585
R3422 GND.n6449 GND.n959 585
R3423 GND.n6452 GND.n6451 585
R3424 GND.n6451 GND.n6450 585
R3425 GND.n6453 GND.n953 585
R3426 GND.n953 GND.n952 585
R3427 GND.n6455 GND.n6454 585
R3428 GND.n6456 GND.n6455 585
R3429 GND.n951 GND.n950 585
R3430 GND.n6457 GND.n951 585
R3431 GND.n6460 GND.n6459 585
R3432 GND.n6459 GND.n6458 585
R3433 GND.n6461 GND.n945 585
R3434 GND.n945 GND.n944 585
R3435 GND.n6463 GND.n6462 585
R3436 GND.n6464 GND.n6463 585
R3437 GND.n943 GND.n942 585
R3438 GND.n6465 GND.n943 585
R3439 GND.n6468 GND.n6467 585
R3440 GND.n6467 GND.n6466 585
R3441 GND.n6469 GND.n937 585
R3442 GND.n937 GND.n936 585
R3443 GND.n6471 GND.n6470 585
R3444 GND.n6472 GND.n6471 585
R3445 GND.n935 GND.n934 585
R3446 GND.n6473 GND.n935 585
R3447 GND.n6476 GND.n6475 585
R3448 GND.n6475 GND.n6474 585
R3449 GND.n6477 GND.n929 585
R3450 GND.n929 GND.n928 585
R3451 GND.n6479 GND.n6478 585
R3452 GND.n6480 GND.n6479 585
R3453 GND.n927 GND.n926 585
R3454 GND.n6481 GND.n927 585
R3455 GND.n6484 GND.n6483 585
R3456 GND.n6483 GND.n6482 585
R3457 GND.n6485 GND.n921 585
R3458 GND.n921 GND.n920 585
R3459 GND.n6487 GND.n6486 585
R3460 GND.n6488 GND.n6487 585
R3461 GND.n919 GND.n918 585
R3462 GND.n6489 GND.n919 585
R3463 GND.n6492 GND.n6491 585
R3464 GND.n6491 GND.n6490 585
R3465 GND.n6493 GND.n913 585
R3466 GND.n913 GND.n912 585
R3467 GND.n6495 GND.n6494 585
R3468 GND.n6496 GND.n6495 585
R3469 GND.n911 GND.n910 585
R3470 GND.n6497 GND.n911 585
R3471 GND.n6500 GND.n6499 585
R3472 GND.n6499 GND.n6498 585
R3473 GND.n6501 GND.n905 585
R3474 GND.n905 GND.n904 585
R3475 GND.n6503 GND.n6502 585
R3476 GND.n6504 GND.n6503 585
R3477 GND.n903 GND.n902 585
R3478 GND.n6505 GND.n903 585
R3479 GND.n6508 GND.n6507 585
R3480 GND.n6507 GND.n6506 585
R3481 GND.n6509 GND.n897 585
R3482 GND.n897 GND.n896 585
R3483 GND.n6511 GND.n6510 585
R3484 GND.n6512 GND.n6511 585
R3485 GND.n895 GND.n894 585
R3486 GND.n6513 GND.n895 585
R3487 GND.n6516 GND.n6515 585
R3488 GND.n6515 GND.n6514 585
R3489 GND.n6517 GND.n889 585
R3490 GND.n889 GND.n888 585
R3491 GND.n6519 GND.n6518 585
R3492 GND.n6520 GND.n6519 585
R3493 GND.n887 GND.n886 585
R3494 GND.n6521 GND.n887 585
R3495 GND.n6524 GND.n6523 585
R3496 GND.n6523 GND.n6522 585
R3497 GND.n6525 GND.n881 585
R3498 GND.n881 GND.n880 585
R3499 GND.n6527 GND.n6526 585
R3500 GND.n6528 GND.n6527 585
R3501 GND.n879 GND.n878 585
R3502 GND.n6529 GND.n879 585
R3503 GND.n6532 GND.n6531 585
R3504 GND.n6531 GND.n6530 585
R3505 GND.n6533 GND.n873 585
R3506 GND.n873 GND.n872 585
R3507 GND.n6535 GND.n6534 585
R3508 GND.n6536 GND.n6535 585
R3509 GND.n871 GND.n870 585
R3510 GND.n6537 GND.n871 585
R3511 GND.n6540 GND.n6539 585
R3512 GND.n6539 GND.n6538 585
R3513 GND.n6541 GND.n865 585
R3514 GND.n865 GND.n864 585
R3515 GND.n6543 GND.n6542 585
R3516 GND.n6544 GND.n6543 585
R3517 GND.n863 GND.n862 585
R3518 GND.n6545 GND.n863 585
R3519 GND.n6548 GND.n6547 585
R3520 GND.n6547 GND.n6546 585
R3521 GND.n6549 GND.n857 585
R3522 GND.n857 GND.n856 585
R3523 GND.n6551 GND.n6550 585
R3524 GND.n6552 GND.n6551 585
R3525 GND.n855 GND.n854 585
R3526 GND.n6553 GND.n855 585
R3527 GND.n6556 GND.n6555 585
R3528 GND.n6555 GND.n6554 585
R3529 GND.n6557 GND.n849 585
R3530 GND.n849 GND.n848 585
R3531 GND.n6559 GND.n6558 585
R3532 GND.n6560 GND.n6559 585
R3533 GND.n847 GND.n846 585
R3534 GND.n6561 GND.n847 585
R3535 GND.n6564 GND.n6563 585
R3536 GND.n6563 GND.n6562 585
R3537 GND.n6565 GND.n841 585
R3538 GND.n841 GND.n840 585
R3539 GND.n6567 GND.n6566 585
R3540 GND.n6568 GND.n6567 585
R3541 GND.n839 GND.n838 585
R3542 GND.n6569 GND.n839 585
R3543 GND.n6572 GND.n6571 585
R3544 GND.n6571 GND.n6570 585
R3545 GND.n6573 GND.n833 585
R3546 GND.n833 GND.n832 585
R3547 GND.n6575 GND.n6574 585
R3548 GND.n6576 GND.n6575 585
R3549 GND.n831 GND.n830 585
R3550 GND.n6577 GND.n831 585
R3551 GND.n6580 GND.n6579 585
R3552 GND.n6579 GND.n6578 585
R3553 GND.n6581 GND.n825 585
R3554 GND.n825 GND.n824 585
R3555 GND.n6583 GND.n6582 585
R3556 GND.n6584 GND.n6583 585
R3557 GND.n822 GND.n821 585
R3558 GND.n6585 GND.n822 585
R3559 GND.n6588 GND.n6587 585
R3560 GND.n6587 GND.n6586 585
R3561 GND.n6589 GND.n816 585
R3562 GND.n823 GND.n816 585
R3563 GND.n6592 GND.n6590 585
R3564 GND.n6592 GND.n6591 585
R3565 GND.n6593 GND.n815 585
R3566 GND.n6593 GND.n647 585
R3567 GND.n6595 GND.n6594 585
R3568 GND.n6594 GND.n644 585
R3569 GND.n6596 GND.n810 585
R3570 GND.n810 GND.n638 585
R3571 GND.n6598 GND.n6597 585
R3572 GND.n6598 GND.n635 585
R3573 GND.n6599 GND.n809 585
R3574 GND.n6599 GND.n627 585
R3575 GND.n6601 GND.n6600 585
R3576 GND.n6600 GND.n624 585
R3577 GND.n6602 GND.n804 585
R3578 GND.n804 GND.n617 585
R3579 GND.n6604 GND.n6603 585
R3580 GND.n6604 GND.n614 585
R3581 GND.n6605 GND.n803 585
R3582 GND.n6605 GND.n606 585
R3583 GND.n6607 GND.n6606 585
R3584 GND.n6606 GND.n603 585
R3585 GND.n6608 GND.n798 585
R3586 GND.n798 GND.n596 585
R3587 GND.n6610 GND.n6609 585
R3588 GND.n6611 GND.n6610 585
R3589 GND.n799 GND.n797 585
R3590 GND.n797 GND.n586 585
R3591 GND.n4393 GND.n4392 585
R3592 GND.n4393 GND.n583 585
R3593 GND.n4395 GND.n4394 585
R3594 GND.n4394 GND.n576 585
R3595 GND.n4396 GND.n4385 585
R3596 GND.n4385 GND.n573 585
R3597 GND.n4398 GND.n4397 585
R3598 GND.n4398 GND.n566 585
R3599 GND.n4399 GND.n4384 585
R3600 GND.n4399 GND.n563 585
R3601 GND.n4401 GND.n4400 585
R3602 GND.n4400 GND.n554 585
R3603 GND.n4402 GND.n4372 585
R3604 GND.n4372 GND.n551 585
R3605 GND.n4405 GND.n4404 585
R3606 GND.n4406 GND.n4405 585
R3607 GND.n4382 GND.n4371 585
R3608 GND.n4371 GND.n4368 585
R3609 GND.n4380 GND.n4379 585
R3610 GND.n4379 GND.n4364 585
R3611 GND.n4378 GND.n4373 585
R3612 GND.n4378 GND.n535 585
R3613 GND.n4377 GND.n4376 585
R3614 GND.n4377 GND.n533 585
R3615 GND.n4374 GND.n4038 585
R3616 GND.n4041 GND.n4038 585
R3617 GND.n4482 GND.n4481 585
R3618 GND.n4481 GND.n4480 585
R3619 GND.n4483 GND.n4035 585
R3620 GND.n4045 GND.n4035 585
R3621 GND.n4486 GND.n4485 585
R3622 GND.n4487 GND.n4486 585
R3623 GND.n4036 GND.n4034 585
R3624 GND.n4034 GND.n4029 585
R3625 GND.n4087 GND.n4056 585
R3626 GND.n4056 GND.n4026 585
R3627 GND.n4089 GND.n4088 585
R3628 GND.n4090 GND.n4089 585
R3629 GND.n4057 GND.n4055 585
R3630 GND.n4055 GND.n4017 585
R3631 GND.n4081 GND.n4080 585
R3632 GND.n4080 GND.n4008 585
R3633 GND.n4079 GND.n4059 585
R3634 GND.n4079 GND.n4005 585
R3635 GND.n4078 GND.n4077 585
R3636 GND.n4078 GND.n3998 585
R3637 GND.n4061 GND.n4060 585
R3638 GND.n4060 GND.n3995 585
R3639 GND.n4073 GND.n4072 585
R3640 GND.n4072 GND.n3987 585
R3641 GND.n4071 GND.n4063 585
R3642 GND.n4071 GND.n3984 585
R3643 GND.n4070 GND.n4069 585
R3644 GND.n4070 GND.n3975 585
R3645 GND.n4065 GND.n4064 585
R3646 GND.n4064 GND.n3972 585
R3647 GND.n3952 GND.n3951 585
R3648 GND.n3957 GND.n3952 585
R3649 GND.n4532 GND.n4531 585
R3650 GND.n4531 GND.n4530 585
R3651 GND.n4533 GND.n3946 585
R3652 GND.n3953 GND.n3946 585
R3653 GND.n4535 GND.n4534 585
R3654 GND.n4536 GND.n4535 585
R3655 GND.n3947 GND.n3945 585
R3656 GND.n3945 GND.n3933 585
R3657 GND.n4132 GND.n4106 585
R3658 GND.n4106 GND.n3930 585
R3659 GND.n4134 GND.n4133 585
R3660 GND.n4135 GND.n4134 585
R3661 GND.n4107 GND.n4105 585
R3662 GND.n4105 GND.n3923 585
R3663 GND.n4126 GND.n4125 585
R3664 GND.n4125 GND.n3887 585
R3665 GND.n4124 GND.n4109 585
R3666 GND.n4124 GND.n4123 585
R3667 GND.n4118 GND.n4110 585
R3668 GND.n4122 GND.n4110 585
R3669 GND.n4120 GND.n4119 585
R3670 GND.n4121 GND.n4120 585
R3671 GND.n4113 GND.n4112 585
R3672 GND.n4112 GND.n4111 585
R3673 GND.n3241 GND.n3240 585
R3674 GND.n3244 GND.n3241 585
R3675 GND.n4673 GND.n4672 585
R3676 GND.n4672 GND.n4671 585
R3677 GND.n4674 GND.n3235 585
R3678 GND.n3839 GND.n3235 585
R3679 GND.n4676 GND.n4675 585
R3680 GND.n4677 GND.n4676 585
R3681 GND.n3223 GND.n3222 585
R3682 GND.n3226 GND.n3223 585
R3683 GND.n4687 GND.n4686 585
R3684 GND.n4686 GND.n4685 585
R3685 GND.n4688 GND.n3217 585
R3686 GND.n3823 GND.n3217 585
R3687 GND.n4690 GND.n4689 585
R3688 GND.n4691 GND.n4690 585
R3689 GND.n3218 GND.n3216 585
R3690 GND.n3216 GND.n3212 585
R3691 GND.n3746 GND.n3322 585
R3692 GND.n3322 GND.n3206 585
R3693 GND.n3748 GND.n3747 585
R3694 GND.n3749 GND.n3748 585
R3695 GND.n3323 GND.n3321 585
R3696 GND.n3321 GND.n3320 585
R3697 GND.n3740 GND.n3739 585
R3698 GND.n3739 GND.n3192 585
R3699 GND.n3738 GND.n3325 585
R3700 GND.n3738 GND.n3186 585
R3701 GND.n3737 GND.n3340 585
R3702 GND.n3737 GND.n3736 585
R3703 GND.n3327 GND.n3326 585
R3704 GND.n3341 GND.n3326 585
R3705 GND.n3336 GND.n3335 585
R3706 GND.n3335 GND.n3172 585
R3707 GND.n3334 GND.n3329 585
R3708 GND.n3334 GND.n3166 585
R3709 GND.n3333 GND.n3332 585
R3710 GND.n3333 GND.n3163 585
R3711 GND.n3147 GND.n3146 585
R3712 GND.n3358 GND.n3147 585
R3713 GND.n4737 GND.n4736 585
R3714 GND.n4736 GND.n4735 585
R3715 GND.n4738 GND.n3133 585
R3716 GND.n3361 GND.n3133 585
R3717 GND.n4740 GND.n4739 585
R3718 GND.n4741 GND.n4740 585
R3719 GND.n3134 GND.n3132 585
R3720 GND.n3132 GND.n3123 585
R3721 GND.n3140 GND.n3139 585
R3722 GND.n3139 GND.n3120 585
R3723 GND.n3138 GND.n3137 585
R3724 GND.n3138 GND.n3106 585
R3725 GND.n3094 GND.n3093 585
R3726 GND.n3103 GND.n3094 585
R3727 GND.n4764 GND.n4763 585
R3728 GND.n4763 GND.n4762 585
R3729 GND.n4765 GND.n3083 585
R3730 GND.n3651 GND.n3083 585
R3731 GND.n4767 GND.n4766 585
R3732 GND.n4768 GND.n4767 585
R3733 GND.n3084 GND.n3082 585
R3734 GND.n3642 GND.n3082 585
R3735 GND.n3087 GND.n3086 585
R3736 GND.n3086 GND.n3062 585
R3737 GND.n3050 GND.n3049 585
R3738 GND.n3059 GND.n3050 585
R3739 GND.n4785 GND.n4784 585
R3740 GND.n4784 GND.n4783 585
R3741 GND.n4786 GND.n3039 585
R3742 GND.n3627 GND.n3039 585
R3743 GND.n4788 GND.n4787 585
R3744 GND.n4789 GND.n4788 585
R3745 GND.n3040 GND.n3038 585
R3746 GND.n3038 GND.n3029 585
R3747 GND.n3043 GND.n3042 585
R3748 GND.n3042 GND.n3026 585
R3749 GND.n3005 GND.n3004 585
R3750 GND.n3381 GND.n3005 585
R3751 GND.n4806 GND.n4805 585
R3752 GND.n4805 GND.n4804 585
R3753 GND.n4807 GND.n2999 585
R3754 GND.n3387 GND.n2999 585
R3755 GND.n4809 GND.n4808 585
R3756 GND.n4810 GND.n4809 585
R3757 GND.n3000 GND.n2998 585
R3758 GND.n2998 GND.n2989 585
R3759 GND.n3551 GND.n3550 585
R3760 GND.n3552 GND.n3551 585
R3761 GND.n3545 GND.n3544 585
R3762 GND.n3544 GND.n3543 585
R3763 GND.n2946 GND.n2945 585
R3764 GND.n2955 GND.n2946 585
R3765 GND.n4861 GND.n4860 585
R3766 GND.n4860 GND.t223 585
R3767 GND.n4862 GND.n2940 585
R3768 GND.n3529 GND.n2940 585
R3769 GND.n4864 GND.n4863 585
R3770 GND.n4865 GND.n4864 585
R3771 GND.n2928 GND.n2927 585
R3772 GND.n2937 GND.n2928 585
R3773 GND.n4875 GND.n4874 585
R3774 GND.n4874 GND.n4873 585
R3775 GND.n4876 GND.n2922 585
R3776 GND.n2929 GND.n2922 585
R3777 GND.n4878 GND.n4877 585
R3778 GND.n4879 GND.n4878 585
R3779 GND.n2920 GND.n2919 585
R3780 GND.n4880 GND.n2920 585
R3781 GND.n4883 GND.n4882 585
R3782 GND.n4882 GND.n4881 585
R3783 GND.n4884 GND.n2060 585
R3784 GND.n2060 GND.n2058 585
R3785 GND.n4886 GND.n4885 585
R3786 GND.n4887 GND.n4886 585
R3787 GND.n2061 GND.n2059 585
R3788 GND.n2059 GND.n2032 585
R3789 GND.n2913 GND.n2912 585
R3790 GND.n2912 GND.n1988 585
R3791 GND.n2911 GND.n2063 585
R3792 GND.n2911 GND.n1986 585
R3793 GND.n2910 GND.n2065 585
R3794 GND.n2910 GND.n2909 585
R3795 GND.n2833 GND.n2064 585
R3796 GND.n2071 GND.n2064 585
R3797 GND.n2835 GND.n2834 585
R3798 GND.n2836 GND.n2835 585
R3799 GND.n2091 GND.n2090 585
R3800 GND.n2090 GND.n2081 585
R3801 GND.n2827 GND.n2826 585
R3802 GND.n2826 GND.n2078 585
R3803 GND.n2825 GND.n2093 585
R3804 GND.n2825 GND.n2084 585
R3805 GND.n2824 GND.n2095 585
R3806 GND.n2824 GND.n2823 585
R3807 GND.n2720 GND.n2094 585
R3808 GND.n2105 GND.n2094 585
R3809 GND.n2722 GND.n2721 585
R3810 GND.n2721 GND.n2102 585
R3811 GND.n2723 GND.n2713 585
R3812 GND.n2713 GND.n2712 585
R3813 GND.n2725 GND.n2724 585
R3814 GND.n2725 GND.n2115 585
R3815 GND.n2726 GND.n2710 585
R3816 GND.n2726 GND.n2114 585
R3817 GND.n2728 GND.n2727 585
R3818 GND.n2727 GND.n2125 585
R3819 GND.n2729 GND.n2705 585
R3820 GND.n2705 GND.n2123 585
R3821 GND.n2733 GND.n2730 585
R3822 GND.n2733 GND.n2732 585
R3823 GND.n2734 GND.n2704 585
R3824 GND.n2734 GND.n2136 585
R3825 GND.n2736 GND.n2735 585
R3826 GND.n2735 GND.n2134 585
R3827 GND.n2737 GND.n2700 585
R3828 GND.n2700 GND.n2699 585
R3829 GND.n2740 GND.n2739 585
R3830 GND.n2741 GND.n2740 585
R3831 GND.n2702 GND.n2696 585
R3832 GND.n2696 GND.n2180 585
R3833 GND.n2163 GND.n2162 585
R3834 GND.n2167 GND.n2163 585
R3835 GND.n2753 GND.n2752 585
R3836 GND.n2752 GND.n2751 585
R3837 GND.n2755 GND.n2160 585
R3838 GND.n2164 GND.n2160 585
R3839 GND.n2757 GND.n2756 585
R3840 GND.n2758 GND.n2757 585
R3841 GND.n2647 GND.n2159 585
R3842 GND.n2159 GND.n2152 585
R3843 GND.n2649 GND.n2648 585
R3844 GND.n2649 GND.n2150 585
R3845 GND.n2654 GND.n2645 585
R3846 GND.n2654 GND.n2653 585
R3847 GND.n2656 GND.n2655 585
R3848 GND.n2655 GND.n2198 585
R3849 GND.n2657 GND.n2216 585
R3850 GND.n2216 GND.n2196 585
R3851 GND.n2659 GND.n2658 585
R3852 GND.n2660 GND.n2659 585
R3853 GND.n2217 GND.n2215 585
R3854 GND.n2215 GND.n2209 585
R3855 GND.n2639 GND.n2638 585
R3856 GND.n2638 GND.n2207 585
R3857 GND.n2637 GND.n2219 585
R3858 GND.n2637 GND.n2636 585
R3859 GND.n2573 GND.n2220 585
R3860 GND.n2230 GND.n2220 585
R3861 GND.n2575 GND.n2574 585
R3862 GND.n2574 GND.n2229 585
R3863 GND.n2576 GND.n2567 585
R3864 GND.n2567 GND.n2243 585
R3865 GND.n2578 GND.n2577 585
R3866 GND.n2578 GND.n2240 585
R3867 GND.n2579 GND.n2566 585
R3868 GND.n2579 GND.n2246 585
R3869 GND.n2581 GND.n2580 585
R3870 GND.n2580 GND.n2254 585
R3871 GND.n2582 GND.n2550 585
R3872 GND.n2550 GND.n2253 585
R3873 GND.n2584 GND.n2583 585
R3874 GND.n2585 GND.n2584 585
R3875 GND.n2551 GND.n2549 585
R3876 GND.n2549 GND.n2261 585
R3877 GND.n2560 GND.n2559 585
R3878 GND.n2559 GND.n1889 585
R3879 GND.n2558 GND.n2553 585
R3880 GND.n2558 GND.n1886 585
R3881 GND.n2557 GND.n2556 585
R3882 GND.n2557 GND.n1877 585
R3883 GND.n1873 GND.n1872 585
R3884 GND.n5135 GND.n1873 585
R3885 GND.n5138 GND.n5137 585
R3886 GND.n5137 GND.n5136 585
R3887 GND.n5139 GND.n1867 585
R3888 GND.n1867 GND.n1866 585
R3889 GND.n5141 GND.n5140 585
R3890 GND.n5142 GND.n5141 585
R3891 GND.n1865 GND.n1864 585
R3892 GND.n5143 GND.n1865 585
R3893 GND.n5146 GND.n5145 585
R3894 GND.n5145 GND.n5144 585
R3895 GND.n5147 GND.n1859 585
R3896 GND.n1859 GND.n1858 585
R3897 GND.n5149 GND.n5148 585
R3898 GND.n5150 GND.n5149 585
R3899 GND.n1857 GND.n1856 585
R3900 GND.n5151 GND.n1857 585
R3901 GND.n5154 GND.n5153 585
R3902 GND.n5153 GND.n5152 585
R3903 GND.n5155 GND.n1851 585
R3904 GND.n1851 GND.n1850 585
R3905 GND.n5157 GND.n5156 585
R3906 GND.n5158 GND.n5157 585
R3907 GND.n1849 GND.n1848 585
R3908 GND.n5159 GND.n1849 585
R3909 GND.n5162 GND.n5161 585
R3910 GND.n5161 GND.n5160 585
R3911 GND.n5163 GND.n1843 585
R3912 GND.n1843 GND.n1842 585
R3913 GND.n5165 GND.n5164 585
R3914 GND.n5166 GND.n5165 585
R3915 GND.n1841 GND.n1840 585
R3916 GND.n5167 GND.n1841 585
R3917 GND.n5170 GND.n5169 585
R3918 GND.n5169 GND.n5168 585
R3919 GND.n5171 GND.n1835 585
R3920 GND.n1835 GND.n1834 585
R3921 GND.n5173 GND.n5172 585
R3922 GND.n5174 GND.n5173 585
R3923 GND.n1833 GND.n1832 585
R3924 GND.n5175 GND.n1833 585
R3925 GND.n5178 GND.n5177 585
R3926 GND.n5177 GND.n5176 585
R3927 GND.n5179 GND.n1827 585
R3928 GND.n1827 GND.n1826 585
R3929 GND.n5181 GND.n5180 585
R3930 GND.n5182 GND.n5181 585
R3931 GND.n1825 GND.n1824 585
R3932 GND.n5183 GND.n1825 585
R3933 GND.n5186 GND.n5185 585
R3934 GND.n5185 GND.n5184 585
R3935 GND.n5187 GND.n1819 585
R3936 GND.n1819 GND.n1818 585
R3937 GND.n5189 GND.n5188 585
R3938 GND.n5190 GND.n5189 585
R3939 GND.n1817 GND.n1816 585
R3940 GND.n5191 GND.n1817 585
R3941 GND.n5194 GND.n5193 585
R3942 GND.n5193 GND.n5192 585
R3943 GND.n5195 GND.n1811 585
R3944 GND.n1811 GND.n1810 585
R3945 GND.n5197 GND.n5196 585
R3946 GND.n5198 GND.n5197 585
R3947 GND.n1809 GND.n1808 585
R3948 GND.n5199 GND.n1809 585
R3949 GND.n5202 GND.n5201 585
R3950 GND.n5201 GND.n5200 585
R3951 GND.n5203 GND.n1803 585
R3952 GND.n1803 GND.n1802 585
R3953 GND.n5205 GND.n5204 585
R3954 GND.n5206 GND.n5205 585
R3955 GND.n1801 GND.n1800 585
R3956 GND.n5207 GND.n1801 585
R3957 GND.n5210 GND.n5209 585
R3958 GND.n5209 GND.n5208 585
R3959 GND.n5211 GND.n1795 585
R3960 GND.n1795 GND.n1794 585
R3961 GND.n5213 GND.n5212 585
R3962 GND.n5214 GND.n5213 585
R3963 GND.n1793 GND.n1792 585
R3964 GND.n5215 GND.n1793 585
R3965 GND.n5218 GND.n5217 585
R3966 GND.n5217 GND.n5216 585
R3967 GND.n5219 GND.n1787 585
R3968 GND.n1787 GND.n1786 585
R3969 GND.n5221 GND.n5220 585
R3970 GND.n5222 GND.n5221 585
R3971 GND.n1785 GND.n1784 585
R3972 GND.n5223 GND.n1785 585
R3973 GND.n5226 GND.n5225 585
R3974 GND.n5225 GND.n5224 585
R3975 GND.n5227 GND.n1779 585
R3976 GND.n1779 GND.n1778 585
R3977 GND.n5229 GND.n5228 585
R3978 GND.n5230 GND.n5229 585
R3979 GND.n1777 GND.n1776 585
R3980 GND.n5231 GND.n1777 585
R3981 GND.n5234 GND.n5233 585
R3982 GND.n5233 GND.n5232 585
R3983 GND.n5235 GND.n1771 585
R3984 GND.n1771 GND.n1770 585
R3985 GND.n5237 GND.n5236 585
R3986 GND.n5238 GND.n5237 585
R3987 GND.n1769 GND.n1768 585
R3988 GND.n5239 GND.n1769 585
R3989 GND.n5242 GND.n5241 585
R3990 GND.n5241 GND.n5240 585
R3991 GND.n5243 GND.n1763 585
R3992 GND.n1763 GND.n1762 585
R3993 GND.n5245 GND.n5244 585
R3994 GND.n5246 GND.n5245 585
R3995 GND.n1761 GND.n1760 585
R3996 GND.n5247 GND.n1761 585
R3997 GND.n5250 GND.n5249 585
R3998 GND.n5249 GND.n5248 585
R3999 GND.n5251 GND.n1755 585
R4000 GND.n1755 GND.n1754 585
R4001 GND.n5253 GND.n5252 585
R4002 GND.n5254 GND.n5253 585
R4003 GND.n1753 GND.n1752 585
R4004 GND.n5255 GND.n1753 585
R4005 GND.n5258 GND.n5257 585
R4006 GND.n5257 GND.n5256 585
R4007 GND.n5259 GND.n1747 585
R4008 GND.n1747 GND.n1746 585
R4009 GND.n5261 GND.n5260 585
R4010 GND.n5262 GND.n5261 585
R4011 GND.n1745 GND.n1744 585
R4012 GND.n5263 GND.n1745 585
R4013 GND.n5266 GND.n5265 585
R4014 GND.n5265 GND.n5264 585
R4015 GND.n5267 GND.n1739 585
R4016 GND.n1739 GND.n1738 585
R4017 GND.n5269 GND.n5268 585
R4018 GND.n5270 GND.n5269 585
R4019 GND.n1737 GND.n1736 585
R4020 GND.n5271 GND.n1737 585
R4021 GND.n5274 GND.n5273 585
R4022 GND.n5273 GND.n5272 585
R4023 GND.n5275 GND.n1731 585
R4024 GND.n1731 GND.n1730 585
R4025 GND.n5277 GND.n5276 585
R4026 GND.n5278 GND.n5277 585
R4027 GND.n1729 GND.n1728 585
R4028 GND.n5279 GND.n1729 585
R4029 GND.n5282 GND.n5281 585
R4030 GND.n5281 GND.n5280 585
R4031 GND.n5283 GND.n1723 585
R4032 GND.n1723 GND.n1722 585
R4033 GND.n5285 GND.n5284 585
R4034 GND.n5286 GND.n5285 585
R4035 GND.n1721 GND.n1720 585
R4036 GND.n5287 GND.n1721 585
R4037 GND.n5290 GND.n5289 585
R4038 GND.n5289 GND.n5288 585
R4039 GND.n5291 GND.n1715 585
R4040 GND.n1715 GND.n1714 585
R4041 GND.n5293 GND.n5292 585
R4042 GND.n5294 GND.n5293 585
R4043 GND.n1713 GND.n1712 585
R4044 GND.n5295 GND.n1713 585
R4045 GND.n5298 GND.n5297 585
R4046 GND.n5297 GND.n5296 585
R4047 GND.n5299 GND.n1707 585
R4048 GND.n1707 GND.n1706 585
R4049 GND.n5301 GND.n5300 585
R4050 GND.n5302 GND.n5301 585
R4051 GND.n1705 GND.n1704 585
R4052 GND.n5303 GND.n1705 585
R4053 GND.n5306 GND.n5305 585
R4054 GND.n5305 GND.n5304 585
R4055 GND.n5307 GND.n1699 585
R4056 GND.n1699 GND.n1698 585
R4057 GND.n5309 GND.n5308 585
R4058 GND.n5310 GND.n5309 585
R4059 GND.n1697 GND.n1696 585
R4060 GND.n5311 GND.n1697 585
R4061 GND.n5314 GND.n5313 585
R4062 GND.n5313 GND.n5312 585
R4063 GND.n5315 GND.n1690 585
R4064 GND.n1690 GND.n1689 585
R4065 GND.n5317 GND.n5316 585
R4066 GND.n5318 GND.n5317 585
R4067 GND.n1691 GND.n1688 585
R4068 GND.n5319 GND.n1688 585
R4069 GND.n5321 GND.n1687 585
R4070 GND.n5321 GND.n5320 585
R4071 GND.n5323 GND.n5322 585
R4072 GND.n5322 GND.n1682 585
R4073 GND.n2279 GND.n2278 585
R4074 GND.n2278 GND.n1874 585
R4075 GND.n2511 GND.n2510 585
R4076 GND.n2513 GND.n2277 585
R4077 GND.n2516 GND.n2515 585
R4078 GND.n2275 GND.n2274 585
R4079 GND.n2521 GND.n2520 585
R4080 GND.n2523 GND.n2273 585
R4081 GND.n2526 GND.n2525 585
R4082 GND.n2271 GND.n2270 585
R4083 GND.n2531 GND.n2530 585
R4084 GND.n2533 GND.n2269 585
R4085 GND.n2535 GND.n2534 585
R4086 GND.n2534 GND.n1874 585
R4087 GND.n1989 GND.n1982 585
R4088 GND.n5056 GND.n1989 585
R4089 GND.n2907 GND.n1981 585
R4090 GND.n2908 GND.n2907 585
R4091 GND.n2906 GND.n1980 585
R4092 GND.n2906 GND.n2066 585
R4093 GND.n2905 GND.n2069 585
R4094 GND.n2905 GND.n2904 585
R4095 GND.n2068 GND.n1974 585
R4096 GND.n2837 GND.n2068 585
R4097 GND.n2893 GND.n1973 585
R4098 GND.n2894 GND.n2893 585
R4099 GND.n2892 GND.n1972 585
R4100 GND.n2892 GND.n2891 585
R4101 GND.n2083 GND.n2082 585
R4102 GND.n2822 GND.n2083 585
R4103 GND.n2812 GND.n1966 585
R4104 GND.n2812 GND.n2096 585
R4105 GND.n2813 GND.n1965 585
R4106 GND.n2814 GND.n2813 585
R4107 GND.n2811 GND.n1964 585
R4108 GND.n2811 GND.n2810 585
R4109 GND.n2107 GND.n2106 585
R4110 GND.n2711 GND.n2107 585
R4111 GND.n2116 GND.n1958 585
R4112 GND.n2798 GND.n2116 585
R4113 GND.n2786 GND.n1957 585
R4114 GND.n2786 GND.n2785 585
R4115 GND.n2787 GND.n1956 585
R4116 GND.n2788 GND.n2787 585
R4117 GND.n2783 GND.n2127 585
R4118 GND.n2783 GND.n2782 585
R4119 GND.n2126 GND.n1950 585
R4120 GND.n2731 GND.n2126 585
R4121 GND.n2137 GND.n1949 585
R4122 GND.n2773 GND.n2137 585
R4123 GND.n2697 GND.n1948 585
R4124 GND.n2698 GND.n2697 585
R4125 GND.n2182 GND.n2181 585
R4126 GND.n2695 GND.n2182 585
R4127 GND.n2743 GND.n1942 585
R4128 GND.n2743 GND.n2742 585
R4129 GND.n2744 GND.n1941 585
R4130 GND.n2745 GND.n2744 585
R4131 GND.n2170 GND.n1940 585
R4132 GND.n2750 GND.n2170 585
R4133 GND.n2169 GND.n2168 585
R4134 GND.n2169 GND.n2165 585
R4135 GND.n2155 GND.n1934 585
R4136 GND.n2158 GND.n2155 585
R4137 GND.n2760 GND.n1933 585
R4138 GND.n2760 GND.n2759 585
R4139 GND.n2761 GND.n1932 585
R4140 GND.n2762 GND.n2761 585
R4141 GND.n2154 GND.n2153 585
R4142 GND.n2652 GND.n2154 585
R4143 GND.n2650 GND.n1926 585
R4144 GND.n2651 GND.n2650 585
R4145 GND.n2199 GND.n1925 585
R4146 GND.n2673 GND.n2199 585
R4147 GND.n2211 GND.n1924 585
R4148 GND.n2214 GND.n2211 585
R4149 GND.n2662 GND.n2212 585
R4150 GND.n2662 GND.n2661 585
R4151 GND.n2663 GND.n1918 585
R4152 GND.n2664 GND.n2663 585
R4153 GND.n2210 GND.n1917 585
R4154 GND.n2635 GND.n2210 585
R4155 GND.n2231 GND.n1916 585
R4156 GND.n2231 GND.n2221 585
R4157 GND.n2233 GND.n2232 585
R4158 GND.n2624 GND.n2233 585
R4159 GND.n2612 GND.n1910 585
R4160 GND.n2612 GND.n2611 585
R4161 GND.n2613 GND.n1909 585
R4162 GND.n2614 GND.n2613 585
R4163 GND.n2610 GND.n1908 585
R4164 GND.n2610 GND.n2609 585
R4165 GND.n2245 GND.n2244 585
R4166 GND.n2257 GND.n2245 585
R4167 GND.n2255 GND.n1902 585
R4168 GND.n2600 GND.n2255 585
R4169 GND.n2588 GND.n1901 585
R4170 GND.n2588 GND.n2587 585
R4171 GND.n2589 GND.n1900 585
R4172 GND.n2590 GND.n2589 585
R4173 GND.n1893 GND.n1891 585
R4174 GND.n2262 GND.n1891 585
R4175 GND.n5127 GND.n5126 585
R4176 GND.n5128 GND.n5127 585
R4177 GND.n1892 GND.n1890 585
R4178 GND.n2540 GND.n1890 585
R4179 GND.n2504 GND.n1878 585
R4180 GND.n5134 GND.n1878 585
R4181 GND.n2877 GND.n2876 585
R4182 GND.n2875 GND.n2874 585
R4183 GND.n2873 GND.n2870 585
R4184 GND.n2864 GND.n2842 585
R4185 GND.n2866 GND.n2865 585
R4186 GND.n2863 GND.n2862 585
R4187 GND.n2861 GND.n2860 585
R4188 GND.n2854 GND.n2844 585
R4189 GND.n2856 GND.n2855 585
R4190 GND.n2853 GND.n2852 585
R4191 GND.n2851 GND.n2850 585
R4192 GND.n2847 GND.n2846 585
R4193 GND.n2879 GND.n1987 585
R4194 GND.n5056 GND.n1987 585
R4195 GND.n2840 GND.n2067 585
R4196 GND.n2908 GND.n2067 585
R4197 GND.n2883 GND.n2839 585
R4198 GND.n2839 GND.n2066 585
R4199 GND.n2884 GND.n2070 585
R4200 GND.n2904 GND.n2070 585
R4201 GND.n2885 GND.n2838 585
R4202 GND.n2838 GND.n2837 585
R4203 GND.n2087 GND.n2080 585
R4204 GND.n2894 GND.n2080 585
R4205 GND.n2890 GND.n2889 585
R4206 GND.n2891 GND.n2890 585
R4207 GND.n2086 GND.n2085 585
R4208 GND.n2822 GND.n2085 585
R4209 GND.n2804 GND.n2803 585
R4210 GND.n2803 GND.n2096 585
R4211 GND.n2110 GND.n2104 585
R4212 GND.n2814 GND.n2104 585
R4213 GND.n2809 GND.n2808 585
R4214 GND.n2810 GND.n2809 585
R4215 GND.n2109 GND.n2108 585
R4216 GND.n2711 GND.n2108 585
R4217 GND.n2800 GND.n2799 585
R4218 GND.n2799 GND.n2798 585
R4219 GND.n2113 GND.n2112 585
R4220 GND.n2785 GND.n2113 585
R4221 GND.n2130 GND.n2124 585
R4222 GND.n2788 GND.n2124 585
R4223 GND.n2781 GND.n2780 585
R4224 GND.n2782 GND.n2781 585
R4225 GND.n2129 GND.n2128 585
R4226 GND.n2731 GND.n2128 585
R4227 GND.n2775 GND.n2774 585
R4228 GND.n2774 GND.n2773 585
R4229 GND.n2133 GND.n2132 585
R4230 GND.n2698 GND.n2133 585
R4231 GND.n2692 GND.n2691 585
R4232 GND.n2695 GND.n2692 585
R4233 GND.n2184 GND.n2183 585
R4234 GND.n2742 GND.n2183 585
R4235 GND.n2687 GND.n2179 585
R4236 GND.n2745 GND.n2179 585
R4237 GND.n2686 GND.n2166 585
R4238 GND.n2750 GND.n2166 585
R4239 GND.n2685 GND.n2188 585
R4240 GND.n2188 GND.n2165 585
R4241 GND.n2187 GND.n2186 585
R4242 GND.n2187 GND.n2158 585
R4243 GND.n2681 GND.n2157 585
R4244 GND.n2759 GND.n2157 585
R4245 GND.n2680 GND.n2151 585
R4246 GND.n2762 GND.n2151 585
R4247 GND.n2679 GND.n2191 585
R4248 GND.n2652 GND.n2191 585
R4249 GND.n2195 GND.n2190 585
R4250 GND.n2651 GND.n2195 585
R4251 GND.n2675 GND.n2674 585
R4252 GND.n2674 GND.n2673 585
R4253 GND.n2194 GND.n2193 585
R4254 GND.n2214 GND.n2194 585
R4255 GND.n2629 GND.n2213 585
R4256 GND.n2661 GND.n2213 585
R4257 GND.n2225 GND.n2208 585
R4258 GND.n2664 GND.n2208 585
R4259 GND.n2634 GND.n2633 585
R4260 GND.n2635 GND.n2634 585
R4261 GND.n2224 GND.n2223 585
R4262 GND.n2223 GND.n2221 585
R4263 GND.n2626 GND.n2625 585
R4264 GND.n2625 GND.n2624 585
R4265 GND.n2228 GND.n2227 585
R4266 GND.n2611 GND.n2228 585
R4267 GND.n2249 GND.n2242 585
R4268 GND.n2614 GND.n2242 585
R4269 GND.n2608 GND.n2607 585
R4270 GND.n2609 GND.n2608 585
R4271 GND.n2248 GND.n2247 585
R4272 GND.n2257 GND.n2247 585
R4273 GND.n2602 GND.n2601 585
R4274 GND.n2601 GND.n2600 585
R4275 GND.n2252 GND.n2251 585
R4276 GND.n2587 GND.n2252 585
R4277 GND.n2548 GND.n2547 585
R4278 GND.n2590 GND.n2548 585
R4279 GND.n2264 GND.n2263 585
R4280 GND.n2263 GND.n2262 585
R4281 GND.n2543 GND.n1888 585
R4282 GND.n5128 GND.n1888 585
R4283 GND.n2542 GND.n2541 585
R4284 GND.n2541 GND.n2540 585
R4285 GND.n2538 GND.n1876 585
R4286 GND.n5134 GND.n1876 585
R4287 GND.n4669 GND.n3246 535.745
R4288 GND.n3848 GND.n3243 535.745
R4289 GND.n3520 GND.n3519 535.745
R4290 GND.n3451 GND.n2932 535.745
R4291 GND.n6399 GND.n6398 484.329
R4292 GND.n6290 GND.n6289 301.784
R4293 GND.n6290 GND.n1067 301.784
R4294 GND.n6298 GND.n1067 301.784
R4295 GND.n6299 GND.n6298 301.784
R4296 GND.n6300 GND.n6299 301.784
R4297 GND.n6300 GND.n1061 301.784
R4298 GND.n6308 GND.n1061 301.784
R4299 GND.n6309 GND.n6308 301.784
R4300 GND.n6310 GND.n6309 301.784
R4301 GND.n6310 GND.n1055 301.784
R4302 GND.n6318 GND.n1055 301.784
R4303 GND.n6319 GND.n6318 301.784
R4304 GND.n6320 GND.n6319 301.784
R4305 GND.n6320 GND.n1049 301.784
R4306 GND.n6328 GND.n1049 301.784
R4307 GND.n6329 GND.n6328 301.784
R4308 GND.n6330 GND.n6329 301.784
R4309 GND.n6330 GND.n1043 301.784
R4310 GND.n6338 GND.n1043 301.784
R4311 GND.n6339 GND.n6338 301.784
R4312 GND.n6340 GND.n6339 301.784
R4313 GND.n6340 GND.n1037 301.784
R4314 GND.n6348 GND.n1037 301.784
R4315 GND.n6349 GND.n6348 301.784
R4316 GND.n6350 GND.n6349 301.784
R4317 GND.n6350 GND.n1031 301.784
R4318 GND.n6358 GND.n1031 301.784
R4319 GND.n6359 GND.n6358 301.784
R4320 GND.n6360 GND.n6359 301.784
R4321 GND.n6360 GND.n1025 301.784
R4322 GND.n6368 GND.n1025 301.784
R4323 GND.n6369 GND.n6368 301.784
R4324 GND.n6370 GND.n6369 301.784
R4325 GND.n6370 GND.n1019 301.784
R4326 GND.n6378 GND.n1019 301.784
R4327 GND.n6379 GND.n6378 301.784
R4328 GND.n6380 GND.n6379 301.784
R4329 GND.n6380 GND.n1013 301.784
R4330 GND.n6388 GND.n1013 301.784
R4331 GND.n6389 GND.n6388 301.784
R4332 GND.n6390 GND.n6389 301.784
R4333 GND.n6390 GND.n1007 301.784
R4334 GND.n6398 GND.n1007 301.784
R4335 GND.n233 GND.n219 289.615
R4336 GND.n256 GND.n242 289.615
R4337 GND.n189 GND.n175 289.615
R4338 GND.n212 GND.n198 289.615
R4339 GND.n145 GND.n131 289.615
R4340 GND.n168 GND.n154 289.615
R4341 GND.n101 GND.n87 289.615
R4342 GND.n124 GND.n110 289.615
R4343 GND.n57 GND.n43 289.615
R4344 GND.n80 GND.n66 289.615
R4345 GND.n14 GND.n0 289.615
R4346 GND.n37 GND.n23 289.615
R4347 GND.n520 GND.n506 289.615
R4348 GND.n497 GND.n483 289.615
R4349 GND.n476 GND.n462 289.615
R4350 GND.n453 GND.n439 289.615
R4351 GND.n432 GND.n418 289.615
R4352 GND.n409 GND.n395 289.615
R4353 GND.n388 GND.n374 289.615
R4354 GND.n365 GND.n351 289.615
R4355 GND.n344 GND.n330 289.615
R4356 GND.n321 GND.n307 289.615
R4357 GND.n301 GND.n287 289.615
R4358 GND.n278 GND.n264 289.615
R4359 GND.n5420 GND.n5419 280.613
R4360 GND.n5420 GND.n1589 280.613
R4361 GND.n5428 GND.n1589 280.613
R4362 GND.n5429 GND.n5428 280.613
R4363 GND.n5430 GND.n5429 280.613
R4364 GND.n5430 GND.n1583 280.613
R4365 GND.n5438 GND.n1583 280.613
R4366 GND.n5439 GND.n5438 280.613
R4367 GND.n5440 GND.n5439 280.613
R4368 GND.n5440 GND.n1577 280.613
R4369 GND.n5448 GND.n1577 280.613
R4370 GND.n5449 GND.n5448 280.613
R4371 GND.n5450 GND.n5449 280.613
R4372 GND.n5450 GND.n1571 280.613
R4373 GND.n5458 GND.n1571 280.613
R4374 GND.n5459 GND.n5458 280.613
R4375 GND.n5460 GND.n5459 280.613
R4376 GND.n5460 GND.n1565 280.613
R4377 GND.n5468 GND.n1565 280.613
R4378 GND.n5469 GND.n5468 280.613
R4379 GND.n5470 GND.n5469 280.613
R4380 GND.n5470 GND.n1559 280.613
R4381 GND.n5478 GND.n1559 280.613
R4382 GND.n5479 GND.n5478 280.613
R4383 GND.n5480 GND.n5479 280.613
R4384 GND.n5480 GND.n1553 280.613
R4385 GND.n5488 GND.n1553 280.613
R4386 GND.n5489 GND.n5488 280.613
R4387 GND.n5490 GND.n5489 280.613
R4388 GND.n5490 GND.n1547 280.613
R4389 GND.n5498 GND.n1547 280.613
R4390 GND.n5499 GND.n5498 280.613
R4391 GND.n5500 GND.n5499 280.613
R4392 GND.n5500 GND.n1541 280.613
R4393 GND.n5508 GND.n1541 280.613
R4394 GND.n5509 GND.n5508 280.613
R4395 GND.n5510 GND.n5509 280.613
R4396 GND.n5510 GND.n1535 280.613
R4397 GND.n5518 GND.n1535 280.613
R4398 GND.n5519 GND.n5518 280.613
R4399 GND.n5520 GND.n5519 280.613
R4400 GND.n5520 GND.n1529 280.613
R4401 GND.n5528 GND.n1529 280.613
R4402 GND.n5529 GND.n5528 280.613
R4403 GND.n5530 GND.n5529 280.613
R4404 GND.n5530 GND.n1523 280.613
R4405 GND.n5538 GND.n1523 280.613
R4406 GND.n5539 GND.n5538 280.613
R4407 GND.n5540 GND.n5539 280.613
R4408 GND.n5540 GND.n1517 280.613
R4409 GND.n5548 GND.n1517 280.613
R4410 GND.n5549 GND.n5548 280.613
R4411 GND.n5550 GND.n5549 280.613
R4412 GND.n5550 GND.n1511 280.613
R4413 GND.n5558 GND.n1511 280.613
R4414 GND.n5559 GND.n5558 280.613
R4415 GND.n5560 GND.n5559 280.613
R4416 GND.n5560 GND.n1505 280.613
R4417 GND.n5568 GND.n1505 280.613
R4418 GND.n5569 GND.n5568 280.613
R4419 GND.n5570 GND.n5569 280.613
R4420 GND.n5570 GND.n1499 280.613
R4421 GND.n5578 GND.n1499 280.613
R4422 GND.n5579 GND.n5578 280.613
R4423 GND.n5580 GND.n5579 280.613
R4424 GND.n5580 GND.n1493 280.613
R4425 GND.n5588 GND.n1493 280.613
R4426 GND.n5589 GND.n5588 280.613
R4427 GND.n5590 GND.n5589 280.613
R4428 GND.n5590 GND.n1487 280.613
R4429 GND.n5598 GND.n1487 280.613
R4430 GND.n5599 GND.n5598 280.613
R4431 GND.n5600 GND.n5599 280.613
R4432 GND.n5600 GND.n1481 280.613
R4433 GND.n5608 GND.n1481 280.613
R4434 GND.n5609 GND.n5608 280.613
R4435 GND.n5610 GND.n5609 280.613
R4436 GND.n5610 GND.n1475 280.613
R4437 GND.n5618 GND.n1475 280.613
R4438 GND.n5619 GND.n5618 280.613
R4439 GND.n5620 GND.n5619 280.613
R4440 GND.n5620 GND.n1469 280.613
R4441 GND.n5628 GND.n1469 280.613
R4442 GND.n5629 GND.n5628 280.613
R4443 GND.n5630 GND.n5629 280.613
R4444 GND.n5630 GND.n1463 280.613
R4445 GND.n5638 GND.n1463 280.613
R4446 GND.n5639 GND.n5638 280.613
R4447 GND.n5640 GND.n5639 280.613
R4448 GND.n5640 GND.n1457 280.613
R4449 GND.n5648 GND.n1457 280.613
R4450 GND.n5649 GND.n5648 280.613
R4451 GND.n5650 GND.n5649 280.613
R4452 GND.n5650 GND.n1451 280.613
R4453 GND.n5658 GND.n1451 280.613
R4454 GND.n5659 GND.n5658 280.613
R4455 GND.n5660 GND.n5659 280.613
R4456 GND.n5660 GND.n1445 280.613
R4457 GND.n5668 GND.n1445 280.613
R4458 GND.n5669 GND.n5668 280.613
R4459 GND.n5670 GND.n5669 280.613
R4460 GND.n5670 GND.n1439 280.613
R4461 GND.n5678 GND.n1439 280.613
R4462 GND.n5679 GND.n5678 280.613
R4463 GND.n5680 GND.n5679 280.613
R4464 GND.n5680 GND.n1433 280.613
R4465 GND.n5688 GND.n1433 280.613
R4466 GND.n5689 GND.n5688 280.613
R4467 GND.n5690 GND.n5689 280.613
R4468 GND.n5690 GND.n1427 280.613
R4469 GND.n5698 GND.n1427 280.613
R4470 GND.n5699 GND.n5698 280.613
R4471 GND.n5700 GND.n5699 280.613
R4472 GND.n5700 GND.n1421 280.613
R4473 GND.n5708 GND.n1421 280.613
R4474 GND.n5709 GND.n5708 280.613
R4475 GND.n5710 GND.n5709 280.613
R4476 GND.n5710 GND.n1415 280.613
R4477 GND.n5718 GND.n1415 280.613
R4478 GND.n5719 GND.n5718 280.613
R4479 GND.n5720 GND.n5719 280.613
R4480 GND.n5720 GND.n1409 280.613
R4481 GND.n5728 GND.n1409 280.613
R4482 GND.n5729 GND.n5728 280.613
R4483 GND.n5730 GND.n5729 280.613
R4484 GND.n5730 GND.n1403 280.613
R4485 GND.n5738 GND.n1403 280.613
R4486 GND.n5739 GND.n5738 280.613
R4487 GND.n5740 GND.n5739 280.613
R4488 GND.n5740 GND.n1397 280.613
R4489 GND.n5748 GND.n1397 280.613
R4490 GND.n5749 GND.n5748 280.613
R4491 GND.n5750 GND.n5749 280.613
R4492 GND.n5750 GND.n1391 280.613
R4493 GND.n5758 GND.n1391 280.613
R4494 GND.n5759 GND.n5758 280.613
R4495 GND.n5760 GND.n5759 280.613
R4496 GND.n5760 GND.n1385 280.613
R4497 GND.n5768 GND.n1385 280.613
R4498 GND.n5769 GND.n5768 280.613
R4499 GND.n5770 GND.n5769 280.613
R4500 GND.n5770 GND.n1379 280.613
R4501 GND.n5778 GND.n1379 280.613
R4502 GND.n5779 GND.n5778 280.613
R4503 GND.n5780 GND.n5779 280.613
R4504 GND.n5780 GND.n1373 280.613
R4505 GND.n5788 GND.n1373 280.613
R4506 GND.n5789 GND.n5788 280.613
R4507 GND.n5790 GND.n5789 280.613
R4508 GND.n5790 GND.n1367 280.613
R4509 GND.n5798 GND.n1367 280.613
R4510 GND.n5799 GND.n5798 280.613
R4511 GND.n5800 GND.n5799 280.613
R4512 GND.n5800 GND.n1361 280.613
R4513 GND.n5808 GND.n1361 280.613
R4514 GND.n5809 GND.n5808 280.613
R4515 GND.n5810 GND.n5809 280.613
R4516 GND.n5810 GND.n1355 280.613
R4517 GND.n5818 GND.n1355 280.613
R4518 GND.n5819 GND.n5818 280.613
R4519 GND.n5820 GND.n5819 280.613
R4520 GND.n5820 GND.n1349 280.613
R4521 GND.n5828 GND.n1349 280.613
R4522 GND.n5829 GND.n5828 280.613
R4523 GND.n5830 GND.n5829 280.613
R4524 GND.n5830 GND.n1343 280.613
R4525 GND.n5838 GND.n1343 280.613
R4526 GND.n5839 GND.n5838 280.613
R4527 GND.n5840 GND.n5839 280.613
R4528 GND.n5840 GND.n1337 280.613
R4529 GND.n5848 GND.n1337 280.613
R4530 GND.n5849 GND.n5848 280.613
R4531 GND.n5850 GND.n5849 280.613
R4532 GND.n5850 GND.n1331 280.613
R4533 GND.n5858 GND.n1331 280.613
R4534 GND.n5859 GND.n5858 280.613
R4535 GND.n5860 GND.n5859 280.613
R4536 GND.n5860 GND.n1325 280.613
R4537 GND.n5868 GND.n1325 280.613
R4538 GND.n5869 GND.n5868 280.613
R4539 GND.n5870 GND.n5869 280.613
R4540 GND.n5870 GND.n1319 280.613
R4541 GND.n5878 GND.n1319 280.613
R4542 GND.n5879 GND.n5878 280.613
R4543 GND.n5880 GND.n5879 280.613
R4544 GND.n5880 GND.n1313 280.613
R4545 GND.n5888 GND.n1313 280.613
R4546 GND.n5889 GND.n5888 280.613
R4547 GND.n5890 GND.n5889 280.613
R4548 GND.n5890 GND.n1307 280.613
R4549 GND.n5898 GND.n1307 280.613
R4550 GND.n5899 GND.n5898 280.613
R4551 GND.n5900 GND.n5899 280.613
R4552 GND.n5900 GND.n1301 280.613
R4553 GND.n5908 GND.n1301 280.613
R4554 GND.n5909 GND.n5908 280.613
R4555 GND.n5910 GND.n5909 280.613
R4556 GND.n5910 GND.n1295 280.613
R4557 GND.n5918 GND.n1295 280.613
R4558 GND.n5919 GND.n5918 280.613
R4559 GND.n5920 GND.n5919 280.613
R4560 GND.n5920 GND.n1289 280.613
R4561 GND.n5928 GND.n1289 280.613
R4562 GND.n5929 GND.n5928 280.613
R4563 GND.n5930 GND.n5929 280.613
R4564 GND.n5930 GND.n1283 280.613
R4565 GND.n5938 GND.n1283 280.613
R4566 GND.n5939 GND.n5938 280.613
R4567 GND.n5940 GND.n5939 280.613
R4568 GND.n5940 GND.n1277 280.613
R4569 GND.n5948 GND.n1277 280.613
R4570 GND.n5949 GND.n5948 280.613
R4571 GND.n5950 GND.n5949 280.613
R4572 GND.n5950 GND.n1271 280.613
R4573 GND.n5958 GND.n1271 280.613
R4574 GND.n5959 GND.n5958 280.613
R4575 GND.n5960 GND.n5959 280.613
R4576 GND.n5960 GND.n1265 280.613
R4577 GND.n5968 GND.n1265 280.613
R4578 GND.n5969 GND.n5968 280.613
R4579 GND.n5970 GND.n5969 280.613
R4580 GND.n5970 GND.n1259 280.613
R4581 GND.n5978 GND.n1259 280.613
R4582 GND.n5979 GND.n5978 280.613
R4583 GND.n5980 GND.n5979 280.613
R4584 GND.n5980 GND.n1253 280.613
R4585 GND.n5988 GND.n1253 280.613
R4586 GND.n5989 GND.n5988 280.613
R4587 GND.n5990 GND.n5989 280.613
R4588 GND.n5990 GND.n1247 280.613
R4589 GND.n5998 GND.n1247 280.613
R4590 GND.n5999 GND.n5998 280.613
R4591 GND.n6000 GND.n5999 280.613
R4592 GND.n6000 GND.n1241 280.613
R4593 GND.n6008 GND.n1241 280.613
R4594 GND.n6009 GND.n6008 280.613
R4595 GND.n6010 GND.n6009 280.613
R4596 GND.n6010 GND.n1235 280.613
R4597 GND.n6018 GND.n1235 280.613
R4598 GND.n6019 GND.n6018 280.613
R4599 GND.n6020 GND.n6019 280.613
R4600 GND.n6020 GND.n1229 280.613
R4601 GND.n6028 GND.n1229 280.613
R4602 GND.n6029 GND.n6028 280.613
R4603 GND.n6030 GND.n6029 280.613
R4604 GND.n6030 GND.n1223 280.613
R4605 GND.n6038 GND.n1223 280.613
R4606 GND.n6039 GND.n6038 280.613
R4607 GND.n6040 GND.n6039 280.613
R4608 GND.n6040 GND.n1217 280.613
R4609 GND.n6048 GND.n1217 280.613
R4610 GND.n6049 GND.n6048 280.613
R4611 GND.n6050 GND.n6049 280.613
R4612 GND.n6050 GND.n1211 280.613
R4613 GND.n6058 GND.n1211 280.613
R4614 GND.n6059 GND.n6058 280.613
R4615 GND.n6060 GND.n6059 280.613
R4616 GND.n6060 GND.n1205 280.613
R4617 GND.n6068 GND.n1205 280.613
R4618 GND.n6069 GND.n6068 280.613
R4619 GND.n6070 GND.n6069 280.613
R4620 GND.n6070 GND.n1199 280.613
R4621 GND.n6078 GND.n1199 280.613
R4622 GND.n6079 GND.n6078 280.613
R4623 GND.n6080 GND.n6079 280.613
R4624 GND.n6080 GND.n1193 280.613
R4625 GND.n6088 GND.n1193 280.613
R4626 GND.n6089 GND.n6088 280.613
R4627 GND.n6090 GND.n6089 280.613
R4628 GND.n6090 GND.n1187 280.613
R4629 GND.n6098 GND.n1187 280.613
R4630 GND.n6099 GND.n6098 280.613
R4631 GND.n6100 GND.n6099 280.613
R4632 GND.n6100 GND.n1181 280.613
R4633 GND.n6108 GND.n1181 280.613
R4634 GND.n6109 GND.n6108 280.613
R4635 GND.n6110 GND.n6109 280.613
R4636 GND.n6110 GND.n1175 280.613
R4637 GND.n6118 GND.n1175 280.613
R4638 GND.n6119 GND.n6118 280.613
R4639 GND.n6120 GND.n6119 280.613
R4640 GND.n6120 GND.n1169 280.613
R4641 GND.n6128 GND.n1169 280.613
R4642 GND.n6129 GND.n6128 280.613
R4643 GND.n6130 GND.n6129 280.613
R4644 GND.n6130 GND.n1163 280.613
R4645 GND.n6138 GND.n1163 280.613
R4646 GND.n6139 GND.n6138 280.613
R4647 GND.n6140 GND.n6139 280.613
R4648 GND.n6140 GND.n1157 280.613
R4649 GND.n6148 GND.n1157 280.613
R4650 GND.n6149 GND.n6148 280.613
R4651 GND.n6150 GND.n6149 280.613
R4652 GND.n6150 GND.n1151 280.613
R4653 GND.n6158 GND.n1151 280.613
R4654 GND.n6159 GND.n6158 280.613
R4655 GND.n6160 GND.n6159 280.613
R4656 GND.n6160 GND.n1145 280.613
R4657 GND.n6168 GND.n1145 280.613
R4658 GND.n6169 GND.n6168 280.613
R4659 GND.n6170 GND.n6169 280.613
R4660 GND.n6170 GND.n1139 280.613
R4661 GND.n6178 GND.n1139 280.613
R4662 GND.n6179 GND.n6178 280.613
R4663 GND.n6180 GND.n6179 280.613
R4664 GND.n6180 GND.n1133 280.613
R4665 GND.n6188 GND.n1133 280.613
R4666 GND.n6189 GND.n6188 280.613
R4667 GND.n6190 GND.n6189 280.613
R4668 GND.n6190 GND.n1127 280.613
R4669 GND.n6198 GND.n1127 280.613
R4670 GND.n6199 GND.n6198 280.613
R4671 GND.n6200 GND.n6199 280.613
R4672 GND.n6200 GND.n1121 280.613
R4673 GND.n6208 GND.n1121 280.613
R4674 GND.n6209 GND.n6208 280.613
R4675 GND.n6210 GND.n6209 280.613
R4676 GND.n6210 GND.n1115 280.613
R4677 GND.n6218 GND.n1115 280.613
R4678 GND.n6219 GND.n6218 280.613
R4679 GND.n6220 GND.n6219 280.613
R4680 GND.n6220 GND.n1109 280.613
R4681 GND.n6228 GND.n1109 280.613
R4682 GND.n6229 GND.n6228 280.613
R4683 GND.n6230 GND.n6229 280.613
R4684 GND.n6230 GND.n1103 280.613
R4685 GND.n6238 GND.n1103 280.613
R4686 GND.n6239 GND.n6238 280.613
R4687 GND.n6240 GND.n6239 280.613
R4688 GND.n6240 GND.n1097 280.613
R4689 GND.n6248 GND.n1097 280.613
R4690 GND.n6249 GND.n6248 280.613
R4691 GND.n6250 GND.n6249 280.613
R4692 GND.n6250 GND.n1091 280.613
R4693 GND.n6258 GND.n1091 280.613
R4694 GND.n6259 GND.n6258 280.613
R4695 GND.n6260 GND.n6259 280.613
R4696 GND.n6260 GND.n1085 280.613
R4697 GND.n6268 GND.n1085 280.613
R4698 GND.n6269 GND.n6268 280.613
R4699 GND.n6270 GND.n6269 280.613
R4700 GND.n6270 GND.n1079 280.613
R4701 GND.n6278 GND.n1079 280.613
R4702 GND.n6279 GND.n6278 280.613
R4703 GND.n6280 GND.n6279 280.613
R4704 GND.n6280 GND.n1073 280.613
R4705 GND.n6288 GND.n1073 280.613
R4706 GND.n3452 GND.n2921 256.663
R4707 GND.n3458 GND.n2921 256.663
R4708 GND.n3460 GND.n2921 256.663
R4709 GND.n3466 GND.n2921 256.663
R4710 GND.n3468 GND.n2921 256.663
R4711 GND.n3474 GND.n2921 256.663
R4712 GND.n3476 GND.n2921 256.663
R4713 GND.n3482 GND.n2921 256.663
R4714 GND.n3485 GND.n2921 256.663
R4715 GND.n3487 GND.n2921 256.663
R4716 GND.n3493 GND.n2921 256.663
R4717 GND.n3495 GND.n2921 256.663
R4718 GND.n3501 GND.n2921 256.663
R4719 GND.n3503 GND.n2921 256.663
R4720 GND.n3509 GND.n2921 256.663
R4721 GND.n3511 GND.n2921 256.663
R4722 GND.n3517 GND.n2921 256.663
R4723 GND.n3847 GND.n3282 256.663
R4724 GND.n3853 GND.n3282 256.663
R4725 GND.n3308 GND.n3282 256.663
R4726 GND.n3860 GND.n3282 256.663
R4727 GND.n3305 GND.n3282 256.663
R4728 GND.n3867 GND.n3282 256.663
R4729 GND.n3302 GND.n3282 256.663
R4730 GND.n3875 GND.n3282 256.663
R4731 GND.n3878 GND.n3282 256.663
R4732 GND.n4636 GND.n3879 256.663
R4733 GND.n3296 GND.n3282 256.663
R4734 GND.n4640 GND.n3282 256.663
R4735 GND.n3293 GND.n3282 256.663
R4736 GND.n4648 GND.n3282 256.663
R4737 GND.n3288 GND.n3282 256.663
R4738 GND.n4655 GND.n3282 256.663
R4739 GND.n3285 GND.n3282 256.663
R4740 GND.n4662 GND.n3282 256.663
R4741 GND.n3282 GND.n3281 256.663
R4742 GND.n2871 GND.t121 249.029
R4743 GND.n2006 GND.t210 249.029
R4744 GND.n2024 GND.t131 249.029
R4745 GND.n4900 GND.t160 249.029
R4746 GND.n4926 GND.t125 249.029
R4747 GND.n4953 GND.t173 249.029
R4748 GND.n4561 GND.t157 249.029
R4749 GND.n4576 GND.t231 249.029
R4750 GND.n4161 GND.t216 249.029
R4751 GND.n4194 GND.t148 249.029
R4752 GND.n4136 GND.t191 249.029
R4753 GND.n758 GND.t141 249.029
R4754 GND.n6699 GND.t112 249.029
R4755 GND.n6723 GND.t207 249.029
R4756 GND.n691 GND.t128 249.029
R4757 GND.n668 GND.t213 249.029
R4758 GND.n780 GND.t108 249.029
R4759 GND.n4242 GND.t144 249.029
R4760 GND.n2367 GND.t138 249.029
R4761 GND.n2399 GND.t219 249.029
R4762 GND.n2431 GND.t228 249.029
R4763 GND.n2464 GND.t201 249.029
R4764 GND.n2281 GND.t88 249.029
R4765 GND.n2267 GND.t198 249.029
R4766 GND.n4631 GND.n3917 242.672
R4767 GND.n4631 GND.n3918 242.672
R4768 GND.n4631 GND.n3919 242.672
R4769 GND.n4631 GND.n3920 242.672
R4770 GND.n4631 GND.n3921 242.672
R4771 GND.n4631 GND.n3922 242.672
R4772 GND.n777 GND.n655 242.672
R4773 GND.n6658 GND.n655 242.672
R4774 GND.n773 GND.n655 242.672
R4775 GND.n6665 GND.n655 242.672
R4776 GND.n6668 GND.n655 242.672
R4777 GND.n761 GND.n655 242.672
R4778 GND.n4852 GND.n4851 242.672
R4779 GND.n4852 GND.n2957 242.672
R4780 GND.n4852 GND.n2958 242.672
R4781 GND.n4852 GND.n2959 242.672
R4782 GND.n4852 GND.n2960 242.672
R4783 GND.n4852 GND.n2961 242.672
R4784 GND.n4852 GND.n2962 242.672
R4785 GND.n3808 GND.n3215 242.672
R4786 GND.n3806 GND.n3215 242.672
R4787 GND.n3797 GND.n3215 242.672
R4788 GND.n3795 GND.n3215 242.672
R4789 GND.n3786 GND.n3215 242.672
R4790 GND.n3784 GND.n3215 242.672
R4791 GND.n3776 GND.n3215 242.672
R4792 GND.n3774 GND.n3215 242.672
R4793 GND.n2340 GND.n1874 242.672
R4794 GND.n2349 GND.n1874 242.672
R4795 GND.n2351 GND.n1874 242.672
R4796 GND.n2359 GND.n1874 242.672
R4797 GND.n2361 GND.n1874 242.672
R4798 GND.n2371 GND.n1874 242.672
R4799 GND.n2373 GND.n1874 242.672
R4800 GND.n2381 GND.n1874 242.672
R4801 GND.n2383 GND.n1874 242.672
R4802 GND.n2391 GND.n1874 242.672
R4803 GND.n2393 GND.n1874 242.672
R4804 GND.n2403 GND.n1874 242.672
R4805 GND.n2405 GND.n1874 242.672
R4806 GND.n2413 GND.n1874 242.672
R4807 GND.n2415 GND.n1874 242.672
R4808 GND.n2423 GND.n1874 242.672
R4809 GND.n2425 GND.n1874 242.672
R4810 GND.n2436 GND.n1874 242.672
R4811 GND.n2438 GND.n1874 242.672
R4812 GND.n2446 GND.n1874 242.672
R4813 GND.n2448 GND.n1874 242.672
R4814 GND.n2456 GND.n1874 242.672
R4815 GND.n2458 GND.n1874 242.672
R4816 GND.n2469 GND.n1874 242.672
R4817 GND.n2471 GND.n1874 242.672
R4818 GND.n2479 GND.n1874 242.672
R4819 GND.n2481 GND.n1874 242.672
R4820 GND.n2489 GND.n1874 242.672
R4821 GND.n2491 GND.n1874 242.672
R4822 GND.n2499 GND.n1874 242.672
R4823 GND.n4957 GND.n4888 242.672
R4824 GND.n4955 GND.n4888 242.672
R4825 GND.n4948 GND.n4888 242.672
R4826 GND.n4945 GND.n4888 242.672
R4827 GND.n4940 GND.n4888 242.672
R4828 GND.n4937 GND.n4888 242.672
R4829 GND.n4932 GND.n4888 242.672
R4830 GND.n4929 GND.n4888 242.672
R4831 GND.n4921 GND.n4888 242.672
R4832 GND.n4918 GND.n4888 242.672
R4833 GND.n4913 GND.n4888 242.672
R4834 GND.n4910 GND.n4888 242.672
R4835 GND.n4905 GND.n4888 242.672
R4836 GND.n4898 GND.n4888 242.672
R4837 GND.n4895 GND.n4888 242.672
R4838 GND.n5007 GND.n4888 242.672
R4839 GND.n5010 GND.n2031 242.672
R4840 GND.n5011 GND.n4888 242.672
R4841 GND.n4888 GND.n2051 242.672
R4842 GND.n4888 GND.n2049 242.672
R4843 GND.n4888 GND.n2048 242.672
R4844 GND.n4888 GND.n2046 242.672
R4845 GND.n4888 GND.n2045 242.672
R4846 GND.n4888 GND.n2043 242.672
R4847 GND.n4888 GND.n2042 242.672
R4848 GND.n4888 GND.n2040 242.672
R4849 GND.n4888 GND.n2039 242.672
R4850 GND.n4888 GND.n2038 242.672
R4851 GND.n4888 GND.n2036 242.672
R4852 GND.n4888 GND.n2035 242.672
R4853 GND.n4888 GND.n2033 242.672
R4854 GND.n4631 GND.n4630 242.672
R4855 GND.n4631 GND.n3888 242.672
R4856 GND.n4631 GND.n3889 242.672
R4857 GND.n4631 GND.n3890 242.672
R4858 GND.n4631 GND.n3891 242.672
R4859 GND.n4631 GND.n3892 242.672
R4860 GND.n4631 GND.n3893 242.672
R4861 GND.n4631 GND.n3894 242.672
R4862 GND.n4631 GND.n3895 242.672
R4863 GND.n4631 GND.n3896 242.672
R4864 GND.n4631 GND.n3897 242.672
R4865 GND.n4631 GND.n3898 242.672
R4866 GND.n4631 GND.n3900 242.672
R4867 GND.n4631 GND.n3901 242.672
R4868 GND.n4632 GND.n4631 242.672
R4869 GND.n4631 GND.n3902 242.672
R4870 GND.n4631 GND.n3903 242.672
R4871 GND.n4631 GND.n3904 242.672
R4872 GND.n4631 GND.n3905 242.672
R4873 GND.n4631 GND.n3906 242.672
R4874 GND.n4631 GND.n3907 242.672
R4875 GND.n4631 GND.n3908 242.672
R4876 GND.n4631 GND.n3909 242.672
R4877 GND.n4631 GND.n3910 242.672
R4878 GND.n4631 GND.n3911 242.672
R4879 GND.n4631 GND.n3912 242.672
R4880 GND.n4631 GND.n3913 242.672
R4881 GND.n4631 GND.n3914 242.672
R4882 GND.n4631 GND.n3915 242.672
R4883 GND.n4631 GND.n3916 242.672
R4884 GND.n755 GND.n655 242.672
R4885 GND.n6680 GND.n655 242.672
R4886 GND.n751 GND.n655 242.672
R4887 GND.n6687 GND.n655 242.672
R4888 GND.n744 GND.n655 242.672
R4889 GND.n6694 GND.n655 242.672
R4890 GND.n737 GND.n655 242.672
R4891 GND.n6704 GND.n655 242.672
R4892 GND.n730 GND.n655 242.672
R4893 GND.n6711 GND.n655 242.672
R4894 GND.n723 GND.n655 242.672
R4895 GND.n6718 GND.n655 242.672
R4896 GND.n716 GND.n655 242.672
R4897 GND.n6728 GND.n655 242.672
R4898 GND.n709 GND.n655 242.672
R4899 GND.n6735 GND.n655 242.672
R4900 GND.n702 GND.n655 242.672
R4901 GND.n6742 GND.n655 242.672
R4902 GND.n696 GND.n655 242.672
R4903 GND.n6751 GND.n655 242.672
R4904 GND.n688 GND.n655 242.672
R4905 GND.n6758 GND.n655 242.672
R4906 GND.n681 GND.n655 242.672
R4907 GND.n6765 GND.n655 242.672
R4908 GND.n675 GND.n655 242.672
R4909 GND.n670 GND.n655 242.672
R4910 GND.n6776 GND.n655 242.672
R4911 GND.n662 GND.n655 242.672
R4912 GND.n6783 GND.n655 242.672
R4913 GND.n655 GND.n654 242.672
R4914 GND.n5330 GND.n5329 242.672
R4915 GND.n6400 GND.n6399 242.672
R4916 GND.n2512 GND.n1874 242.672
R4917 GND.n2514 GND.n1874 242.672
R4918 GND.n2522 GND.n1874 242.672
R4919 GND.n2524 GND.n1874 242.672
R4920 GND.n2532 GND.n1874 242.672
R4921 GND.n4888 GND.n2057 242.672
R4922 GND.n4888 GND.n2056 242.672
R4923 GND.n4888 GND.n2055 242.672
R4924 GND.n4888 GND.n2054 242.672
R4925 GND.n4888 GND.n2053 242.672
R4926 GND.n4888 GND.n2052 242.672
R4927 GND.n3426 GND.n3424 240.849
R4928 GND.n3270 GND.n3268 240.849
R4929 GND.n651 GND.n648 240.244
R4930 GND.n6785 GND.n6784 240.244
R4931 GND.n6782 GND.n656 240.244
R4932 GND.n6778 GND.n6777 240.244
R4933 GND.n6775 GND.n663 240.244
R4934 GND.n674 GND.n671 240.244
R4935 GND.n6767 GND.n6766 240.244
R4936 GND.n6764 GND.n676 240.244
R4937 GND.n6760 GND.n6759 240.244
R4938 GND.n6757 GND.n682 240.244
R4939 GND.n6753 GND.n6752 240.244
R4940 GND.n6750 GND.n689 240.244
R4941 GND.n6744 GND.n6743 240.244
R4942 GND.n6741 GND.n697 240.244
R4943 GND.n6737 GND.n6736 240.244
R4944 GND.n6734 GND.n703 240.244
R4945 GND.n6730 GND.n6729 240.244
R4946 GND.n6727 GND.n710 240.244
R4947 GND.n6720 GND.n6719 240.244
R4948 GND.n6717 GND.n717 240.244
R4949 GND.n6713 GND.n6712 240.244
R4950 GND.n6710 GND.n724 240.244
R4951 GND.n6706 GND.n6705 240.244
R4952 GND.n6703 GND.n731 240.244
R4953 GND.n6696 GND.n6695 240.244
R4954 GND.n6693 GND.n738 240.244
R4955 GND.n6689 GND.n6688 240.244
R4956 GND.n6686 GND.n745 240.244
R4957 GND.n6682 GND.n6681 240.244
R4958 GND.n6679 GND.n752 240.244
R4959 GND.n4273 GND.n3931 240.244
R4960 GND.n4538 GND.n3931 240.244
R4961 GND.n4538 GND.n3942 240.244
R4962 GND.n4287 GND.n3942 240.244
R4963 GND.n4287 GND.n3955 240.244
R4964 GND.n4299 GND.n3955 240.244
R4965 GND.n4299 GND.n3973 240.244
R4966 GND.n4309 GND.n3973 240.244
R4967 GND.n4309 GND.n3985 240.244
R4968 GND.n4314 GND.n3985 240.244
R4969 GND.n4314 GND.n3996 240.244
R4970 GND.n4324 GND.n3996 240.244
R4971 GND.n4324 GND.n4006 240.244
R4972 GND.n4329 GND.n4006 240.244
R4973 GND.n4329 GND.n4018 240.244
R4974 GND.n4350 GND.n4018 240.244
R4975 GND.n4350 GND.n4027 240.244
R4976 GND.n4031 GND.n4027 240.244
R4977 GND.n4356 GND.n4031 240.244
R4978 GND.n4356 GND.n4046 240.244
R4979 GND.n4046 GND.n4039 240.244
R4980 GND.n4467 GND.n4039 240.244
R4981 GND.n4467 GND.n534 240.244
R4982 GND.n4463 GND.n534 240.244
R4983 GND.n4463 GND.n4363 240.244
R4984 GND.n4369 GND.n4363 240.244
R4985 GND.n4445 GND.n4369 240.244
R4986 GND.n4445 GND.n552 240.244
R4987 GND.n4441 GND.n552 240.244
R4988 GND.n4441 GND.n564 240.244
R4989 GND.n4433 GND.n564 240.244
R4990 GND.n4433 GND.n574 240.244
R4991 GND.n4429 GND.n574 240.244
R4992 GND.n4429 GND.n584 240.244
R4993 GND.n6613 GND.n584 240.244
R4994 GND.n6613 GND.n594 240.244
R4995 GND.n6617 GND.n594 240.244
R4996 GND.n6617 GND.n604 240.244
R4997 GND.n6627 GND.n604 240.244
R4998 GND.n6627 GND.n615 240.244
R4999 GND.n6631 GND.n615 240.244
R5000 GND.n6631 GND.n625 240.244
R5001 GND.n6642 GND.n625 240.244
R5002 GND.n6642 GND.n636 240.244
R5003 GND.n6647 GND.n636 240.244
R5004 GND.n6647 GND.n645 240.244
R5005 GND.n3925 GND.n3924 240.244
R5006 GND.n4624 GND.n3924 240.244
R5007 GND.n4622 GND.n4621 240.244
R5008 GND.n4618 GND.n4617 240.244
R5009 GND.n4614 GND.n4613 240.244
R5010 GND.n4609 GND.n4559 240.244
R5011 GND.n4607 GND.n4606 240.244
R5012 GND.n4603 GND.n4602 240.244
R5013 GND.n4599 GND.n4598 240.244
R5014 GND.n4595 GND.n4594 240.244
R5015 GND.n4591 GND.n4590 240.244
R5016 GND.n4586 GND.n4574 240.244
R5017 GND.n4584 GND.n4583 240.244
R5018 GND.n3899 GND.n3882 240.244
R5019 GND.n4633 GND.n3881 240.244
R5020 GND.n4152 GND.n3886 240.244
R5021 GND.n4159 GND.n4158 240.244
R5022 GND.n4165 GND.n4164 240.244
R5023 GND.n4172 GND.n4171 240.244
R5024 GND.n4175 GND.n4174 240.244
R5025 GND.n4182 GND.n4181 240.244
R5026 GND.n4185 GND.n4184 240.244
R5027 GND.n4192 GND.n4191 240.244
R5028 GND.n4198 GND.n4197 240.244
R5029 GND.n4205 GND.n4204 240.244
R5030 GND.n4208 GND.n4207 240.244
R5031 GND.n4215 GND.n4214 240.244
R5032 GND.n4218 GND.n4217 240.244
R5033 GND.n4225 GND.n4224 240.244
R5034 GND.n4228 GND.n4227 240.244
R5035 GND.n4545 GND.n3926 240.244
R5036 GND.n4545 GND.n3929 240.244
R5037 GND.n3963 GND.n3929 240.244
R5038 GND.n3963 GND.n3959 240.244
R5039 GND.n4528 GND.n3959 240.244
R5040 GND.n4528 GND.n3960 240.244
R5041 GND.n4524 GND.n3960 240.244
R5042 GND.n4524 GND.n3971 240.244
R5043 GND.n4516 GND.n3971 240.244
R5044 GND.n4516 GND.n3988 240.244
R5045 GND.n4512 GND.n3988 240.244
R5046 GND.n4512 GND.n3994 240.244
R5047 GND.n4504 GND.n3994 240.244
R5048 GND.n4504 GND.n4009 240.244
R5049 GND.n4500 GND.n4009 240.244
R5050 GND.n4500 GND.n4016 240.244
R5051 GND.n4492 GND.n4016 240.244
R5052 GND.n4492 GND.n4489 240.244
R5053 GND.n4489 GND.n4030 240.244
R5054 GND.n4475 GND.n4030 240.244
R5055 GND.n4478 GND.n4475 240.244
R5056 GND.n4478 GND.n537 240.244
R5057 GND.n6854 GND.n537 240.244
R5058 GND.n6854 GND.n538 240.244
R5059 GND.n4453 GND.n538 240.244
R5060 GND.n4455 GND.n4453 240.244
R5061 GND.n4455 GND.n549 240.244
R5062 GND.n6848 GND.n549 240.244
R5063 GND.n6848 GND.n550 240.244
R5064 GND.n6840 GND.n550 240.244
R5065 GND.n6840 GND.n567 240.244
R5066 GND.n6836 GND.n567 240.244
R5067 GND.n6836 GND.n572 240.244
R5068 GND.n6828 GND.n572 240.244
R5069 GND.n6828 GND.n587 240.244
R5070 GND.n6824 GND.n587 240.244
R5071 GND.n6824 GND.n593 240.244
R5072 GND.n6816 GND.n593 240.244
R5073 GND.n6816 GND.n607 240.244
R5074 GND.n6812 GND.n607 240.244
R5075 GND.n6812 GND.n613 240.244
R5076 GND.n6804 GND.n613 240.244
R5077 GND.n6804 GND.n628 240.244
R5078 GND.n6800 GND.n628 240.244
R5079 GND.n6800 GND.n634 240.244
R5080 GND.n6792 GND.n634 240.244
R5081 GND.n1996 GND.n1995 240.244
R5082 GND.n2034 GND.n1999 240.244
R5083 GND.n2001 GND.n2000 240.244
R5084 GND.n2037 GND.n2004 240.244
R5085 GND.n2009 GND.n2005 240.244
R5086 GND.n2041 GND.n2010 240.244
R5087 GND.n2014 GND.n2013 240.244
R5088 GND.n2044 GND.n2015 240.244
R5089 GND.n2019 GND.n2018 240.244
R5090 GND.n2047 GND.n2020 240.244
R5091 GND.n2026 GND.n2023 240.244
R5092 GND.n2050 GND.n2027 240.244
R5093 GND.n5012 GND.n2030 240.244
R5094 GND.n5009 GND.n5008 240.244
R5095 GND.n5006 GND.n4890 240.244
R5096 GND.n4897 GND.n4896 240.244
R5097 GND.n4904 GND.n4899 240.244
R5098 GND.n4907 GND.n4906 240.244
R5099 GND.n4912 GND.n4911 240.244
R5100 GND.n4915 GND.n4914 240.244
R5101 GND.n4920 GND.n4919 240.244
R5102 GND.n4923 GND.n4922 240.244
R5103 GND.n4931 GND.n4930 240.244
R5104 GND.n4934 GND.n4933 240.244
R5105 GND.n4939 GND.n4938 240.244
R5106 GND.n4942 GND.n4941 240.244
R5107 GND.n4947 GND.n4946 240.244
R5108 GND.n4950 GND.n4949 240.244
R5109 GND.n4958 GND.n4956 240.244
R5110 GND.n2539 GND.n1875 240.244
R5111 GND.n2539 GND.n1887 240.244
R5112 GND.n1897 GND.n1887 240.244
R5113 GND.n1898 GND.n1897 240.244
R5114 GND.n2586 GND.n1898 240.244
R5115 GND.n2586 GND.n1904 240.244
R5116 GND.n1905 GND.n1904 240.244
R5117 GND.n1906 GND.n1905 240.244
R5118 GND.n2241 GND.n1906 240.244
R5119 GND.n2241 GND.n1912 240.244
R5120 GND.n1913 GND.n1912 240.244
R5121 GND.n1914 GND.n1913 240.244
R5122 GND.n2222 GND.n1914 240.244
R5123 GND.n2222 GND.n1920 240.244
R5124 GND.n1921 GND.n1920 240.244
R5125 GND.n1922 GND.n1921 240.244
R5126 GND.n2197 GND.n1922 240.244
R5127 GND.n2197 GND.n1928 240.244
R5128 GND.n1929 GND.n1928 240.244
R5129 GND.n1930 GND.n1929 240.244
R5130 GND.n2156 GND.n1930 240.244
R5131 GND.n2156 GND.n1936 240.244
R5132 GND.n1937 GND.n1936 240.244
R5133 GND.n1938 GND.n1937 240.244
R5134 GND.n2178 GND.n1938 240.244
R5135 GND.n2178 GND.n1944 240.244
R5136 GND.n1945 GND.n1944 240.244
R5137 GND.n1946 GND.n1945 240.244
R5138 GND.n2135 GND.n1946 240.244
R5139 GND.n2135 GND.n1952 240.244
R5140 GND.n1953 GND.n1952 240.244
R5141 GND.n1954 GND.n1953 240.244
R5142 GND.n2784 GND.n1954 240.244
R5143 GND.n2784 GND.n1960 240.244
R5144 GND.n1961 GND.n1960 240.244
R5145 GND.n1962 GND.n1961 240.244
R5146 GND.n2103 GND.n1962 240.244
R5147 GND.n2103 GND.n1968 240.244
R5148 GND.n1969 GND.n1968 240.244
R5149 GND.n1970 GND.n1969 240.244
R5150 GND.n2079 GND.n1970 240.244
R5151 GND.n2079 GND.n1976 240.244
R5152 GND.n1977 GND.n1976 240.244
R5153 GND.n1978 GND.n1977 240.244
R5154 GND.n1984 GND.n1978 240.244
R5155 GND.n5057 GND.n1984 240.244
R5156 GND.n2348 GND.n2341 240.244
R5157 GND.n2352 GND.n2350 240.244
R5158 GND.n2358 GND.n2336 240.244
R5159 GND.n2362 GND.n2360 240.244
R5160 GND.n2370 GND.n2332 240.244
R5161 GND.n2374 GND.n2372 240.244
R5162 GND.n2380 GND.n2328 240.244
R5163 GND.n2384 GND.n2382 240.244
R5164 GND.n2390 GND.n2324 240.244
R5165 GND.n2394 GND.n2392 240.244
R5166 GND.n2402 GND.n2320 240.244
R5167 GND.n2406 GND.n2404 240.244
R5168 GND.n2412 GND.n2316 240.244
R5169 GND.n2416 GND.n2414 240.244
R5170 GND.n2422 GND.n2312 240.244
R5171 GND.n2426 GND.n2424 240.244
R5172 GND.n2435 GND.n2308 240.244
R5173 GND.n2439 GND.n2437 240.244
R5174 GND.n2445 GND.n2304 240.244
R5175 GND.n2449 GND.n2447 240.244
R5176 GND.n2455 GND.n2300 240.244
R5177 GND.n2459 GND.n2457 240.244
R5178 GND.n2468 GND.n2296 240.244
R5179 GND.n2472 GND.n2470 240.244
R5180 GND.n2478 GND.n2292 240.244
R5181 GND.n2482 GND.n2480 240.244
R5182 GND.n2488 GND.n2288 240.244
R5183 GND.n2492 GND.n2490 240.244
R5184 GND.n2498 GND.n2284 240.244
R5185 GND.n2501 GND.n2500 240.244
R5186 GND.n5133 GND.n1880 240.244
R5187 GND.n5129 GND.n1880 240.244
R5188 GND.n5129 GND.n1885 240.244
R5189 GND.n2591 GND.n1885 240.244
R5190 GND.n2591 GND.n2256 240.244
R5191 GND.n2599 GND.n2256 240.244
R5192 GND.n2599 GND.n2258 240.244
R5193 GND.n2258 GND.n2239 240.244
R5194 GND.n2615 GND.n2239 240.244
R5195 GND.n2615 GND.n2234 240.244
R5196 GND.n2623 GND.n2234 240.244
R5197 GND.n2623 GND.n2235 240.244
R5198 GND.n2235 GND.n2205 240.244
R5199 GND.n2665 GND.n2205 240.244
R5200 GND.n2665 GND.n2206 240.244
R5201 GND.n2206 GND.n2200 240.244
R5202 GND.n2672 GND.n2200 240.244
R5203 GND.n2672 GND.n2201 240.244
R5204 GND.n2201 GND.n2148 240.244
R5205 GND.n2763 GND.n2148 240.244
R5206 GND.n2763 GND.n2149 240.244
R5207 GND.n2173 GND.n2149 240.244
R5208 GND.n2174 GND.n2173 240.244
R5209 GND.n2749 GND.n2174 240.244
R5210 GND.n2749 GND.n2746 240.244
R5211 GND.n2746 GND.n2175 240.244
R5212 GND.n2694 GND.n2175 240.244
R5213 GND.n2694 GND.n2138 240.244
R5214 GND.n2772 GND.n2138 240.244
R5215 GND.n2772 GND.n2139 240.244
R5216 GND.n2139 GND.n2122 240.244
R5217 GND.n2789 GND.n2122 240.244
R5218 GND.n2789 GND.n2117 240.244
R5219 GND.n2797 GND.n2117 240.244
R5220 GND.n2797 GND.n2118 240.244
R5221 GND.n2118 GND.n2101 240.244
R5222 GND.n2815 GND.n2101 240.244
R5223 GND.n2815 GND.n2097 240.244
R5224 GND.n2821 GND.n2097 240.244
R5225 GND.n2821 GND.n2077 240.244
R5226 GND.n2895 GND.n2077 240.244
R5227 GND.n2895 GND.n2072 240.244
R5228 GND.n2903 GND.n2072 240.244
R5229 GND.n2903 GND.n2073 240.244
R5230 GND.n2073 GND.n1990 240.244
R5231 GND.n5055 GND.n1990 240.244
R5232 GND.n3777 GND.n3775 240.244
R5233 GND.n3783 GND.n3766 240.244
R5234 GND.n3787 GND.n3785 240.244
R5235 GND.n3794 GND.n3762 240.244
R5236 GND.n3798 GND.n3796 240.244
R5237 GND.n3805 GND.n3756 240.244
R5238 GND.n3809 GND.n3807 240.244
R5239 GND.n4818 GND.n2987 240.244
R5240 GND.n3386 GND.n2987 240.244
R5241 GND.n3577 GND.n3386 240.244
R5242 GND.n3577 GND.n3007 240.244
R5243 GND.n3614 GND.n3007 240.244
R5244 GND.n3614 GND.n3027 240.244
R5245 GND.n3610 GND.n3027 240.244
R5246 GND.n3610 GND.n3609 240.244
R5247 GND.n3609 GND.n3608 240.244
R5248 GND.n3608 GND.n3585 240.244
R5249 GND.n3585 GND.n3061 240.244
R5250 GND.n3603 GND.n3061 240.244
R5251 GND.n3603 GND.n3080 240.244
R5252 GND.n3600 GND.n3080 240.244
R5253 GND.n3600 GND.n3599 240.244
R5254 GND.n3599 GND.n3598 240.244
R5255 GND.n3598 GND.n3105 240.244
R5256 GND.n3674 GND.n3105 240.244
R5257 GND.n3674 GND.n3121 240.244
R5258 GND.n3677 GND.n3121 240.244
R5259 GND.n3677 GND.n3363 240.244
R5260 GND.n3683 GND.n3363 240.244
R5261 GND.n3683 GND.n3149 240.244
R5262 GND.n3700 GND.n3149 240.244
R5263 GND.n3700 GND.n3164 240.244
R5264 GND.n3707 GND.n3164 240.244
R5265 GND.n3707 GND.n3174 240.244
R5266 GND.n3734 GND.n3174 240.244
R5267 GND.n3734 GND.n3184 240.244
R5268 GND.n3730 GND.n3184 240.244
R5269 GND.n3730 GND.n3194 240.244
R5270 GND.n3750 GND.n3194 240.244
R5271 GND.n3750 GND.n3204 240.244
R5272 GND.n3815 GND.n3204 240.244
R5273 GND.n2965 GND.n2964 240.244
R5274 GND.n4845 GND.n2964 240.244
R5275 GND.n4843 GND.n4842 240.244
R5276 GND.n4839 GND.n4838 240.244
R5277 GND.n4835 GND.n4834 240.244
R5278 GND.n4831 GND.n4830 240.244
R5279 GND.n4826 GND.n4825 240.244
R5280 GND.n2983 GND.n2963 240.244
R5281 GND.n3016 GND.n2966 240.244
R5282 GND.n3017 GND.n3016 240.244
R5283 GND.n3017 GND.n3009 240.244
R5284 GND.n4802 GND.n3009 240.244
R5285 GND.n4802 GND.n3010 240.244
R5286 GND.n4798 GND.n3010 240.244
R5287 GND.n4798 GND.n3025 240.244
R5288 GND.n3069 GND.n3025 240.244
R5289 GND.n3070 GND.n3069 240.244
R5290 GND.n3070 GND.n3063 240.244
R5291 GND.n4774 GND.n3063 240.244
R5292 GND.n4774 GND.n3064 240.244
R5293 GND.n4770 GND.n3064 240.244
R5294 GND.n4770 GND.n3078 240.244
R5295 GND.n3111 GND.n3078 240.244
R5296 GND.n3111 GND.n3107 240.244
R5297 GND.n4754 GND.n3107 240.244
R5298 GND.n4754 GND.n3108 240.244
R5299 GND.n4750 GND.n3108 240.244
R5300 GND.n4750 GND.n3119 240.244
R5301 GND.n3154 GND.n3119 240.244
R5302 GND.n3154 GND.n3150 240.244
R5303 GND.n4733 GND.n3150 240.244
R5304 GND.n4733 GND.n3151 240.244
R5305 GND.n4729 GND.n3151 240.244
R5306 GND.n4729 GND.n3162 240.244
R5307 GND.n4719 GND.n3162 240.244
R5308 GND.n4719 GND.n3176 240.244
R5309 GND.n4715 GND.n3176 240.244
R5310 GND.n4715 GND.n3182 240.244
R5311 GND.n4705 GND.n3182 240.244
R5312 GND.n4705 GND.n3196 240.244
R5313 GND.n4701 GND.n3196 240.244
R5314 GND.n4701 GND.n3202 240.244
R5315 GND.n6669 GND.n762 240.244
R5316 GND.n6667 GND.n6666 240.244
R5317 GND.n6664 GND.n766 240.244
R5318 GND.n6660 GND.n6659 240.244
R5319 GND.n6657 GND.n774 240.244
R5320 GND.n4275 GND.n3932 240.244
R5321 GND.n3943 GND.n3932 240.244
R5322 GND.n4282 GND.n3943 240.244
R5323 GND.n4283 GND.n4282 240.244
R5324 GND.n4283 GND.n3956 240.244
R5325 GND.n4301 GND.n3956 240.244
R5326 GND.n4301 GND.n3974 240.244
R5327 GND.n4307 GND.n3974 240.244
R5328 GND.n4307 GND.n3986 240.244
R5329 GND.n4316 GND.n3986 240.244
R5330 GND.n4316 GND.n3997 240.244
R5331 GND.n4322 GND.n3997 240.244
R5332 GND.n4322 GND.n4007 240.244
R5333 GND.n4331 GND.n4007 240.244
R5334 GND.n4331 GND.n4019 240.244
R5335 GND.n4348 GND.n4019 240.244
R5336 GND.n4348 GND.n4028 240.244
R5337 GND.n4032 GND.n4028 240.244
R5338 GND.n4343 GND.n4032 240.244
R5339 GND.n4343 GND.n4047 240.244
R5340 GND.n4047 GND.n4040 240.244
R5341 GND.n4040 GND.n531 240.244
R5342 GND.n6856 GND.n531 240.244
R5343 GND.n6856 GND.n532 240.244
R5344 GND.n4451 GND.n532 240.244
R5345 GND.n4451 GND.n4370 240.244
R5346 GND.n4447 GND.n4370 240.244
R5347 GND.n4447 GND.n553 240.244
R5348 GND.n4439 GND.n553 240.244
R5349 GND.n4439 GND.n565 240.244
R5350 GND.n4435 GND.n565 240.244
R5351 GND.n4435 GND.n575 240.244
R5352 GND.n4427 GND.n575 240.244
R5353 GND.n4427 GND.n585 240.244
R5354 GND.n796 GND.n585 240.244
R5355 GND.n796 GND.n595 240.244
R5356 GND.n6619 GND.n595 240.244
R5357 GND.n6619 GND.n605 240.244
R5358 GND.n6625 GND.n605 240.244
R5359 GND.n6625 GND.n616 240.244
R5360 GND.n6633 GND.n616 240.244
R5361 GND.n6633 GND.n626 240.244
R5362 GND.n6640 GND.n626 240.244
R5363 GND.n6640 GND.n637 240.244
R5364 GND.n6649 GND.n637 240.244
R5365 GND.n6649 GND.n646 240.244
R5366 GND.n4264 GND.n4263 240.244
R5367 GND.n4260 GND.n4259 240.244
R5368 GND.n4256 GND.n4255 240.244
R5369 GND.n4252 GND.n4251 240.244
R5370 GND.n4241 GND.n4240 240.244
R5371 GND.n4543 GND.n3934 240.244
R5372 GND.n4543 GND.n3935 240.244
R5373 GND.n4292 GND.n3935 240.244
R5374 GND.n4293 GND.n4292 240.244
R5375 GND.n4293 GND.n3958 240.244
R5376 GND.n3976 GND.n3958 240.244
R5377 GND.n4522 GND.n3976 240.244
R5378 GND.n4522 GND.n3977 240.244
R5379 GND.n4518 GND.n3977 240.244
R5380 GND.n4518 GND.n3983 240.244
R5381 GND.n4510 GND.n3983 240.244
R5382 GND.n4510 GND.n3999 240.244
R5383 GND.n4506 GND.n3999 240.244
R5384 GND.n4506 GND.n4004 240.244
R5385 GND.n4498 GND.n4004 240.244
R5386 GND.n4498 GND.n4020 240.244
R5387 GND.n4494 GND.n4020 240.244
R5388 GND.n4494 GND.n4025 240.244
R5389 GND.n4048 GND.n4025 240.244
R5390 GND.n4473 GND.n4048 240.244
R5391 GND.n4473 GND.n4042 240.244
R5392 GND.n4469 GND.n4042 240.244
R5393 GND.n4469 GND.n536 240.244
R5394 GND.n4461 GND.n536 240.244
R5395 GND.n4461 GND.n4365 240.244
R5396 GND.n4457 GND.n4365 240.244
R5397 GND.n4457 GND.n555 240.244
R5398 GND.n6846 GND.n555 240.244
R5399 GND.n6846 GND.n556 240.244
R5400 GND.n6842 GND.n556 240.244
R5401 GND.n6842 GND.n562 240.244
R5402 GND.n6834 GND.n562 240.244
R5403 GND.n6834 GND.n577 240.244
R5404 GND.n6830 GND.n577 240.244
R5405 GND.n6830 GND.n582 240.244
R5406 GND.n6822 GND.n582 240.244
R5407 GND.n6822 GND.n597 240.244
R5408 GND.n6818 GND.n597 240.244
R5409 GND.n6818 GND.n602 240.244
R5410 GND.n6810 GND.n602 240.244
R5411 GND.n6810 GND.n618 240.244
R5412 GND.n6806 GND.n618 240.244
R5413 GND.n6806 GND.n623 240.244
R5414 GND.n6798 GND.n623 240.244
R5415 GND.n6798 GND.n639 240.244
R5416 GND.n6794 GND.n639 240.244
R5417 GND.n5421 GND.n1594 240.244
R5418 GND.n5421 GND.n1590 240.244
R5419 GND.n5427 GND.n1590 240.244
R5420 GND.n5427 GND.n1588 240.244
R5421 GND.n5431 GND.n1588 240.244
R5422 GND.n5431 GND.n1584 240.244
R5423 GND.n5437 GND.n1584 240.244
R5424 GND.n5437 GND.n1582 240.244
R5425 GND.n5441 GND.n1582 240.244
R5426 GND.n5441 GND.n1578 240.244
R5427 GND.n5447 GND.n1578 240.244
R5428 GND.n5447 GND.n1576 240.244
R5429 GND.n5451 GND.n1576 240.244
R5430 GND.n5451 GND.n1572 240.244
R5431 GND.n5457 GND.n1572 240.244
R5432 GND.n5457 GND.n1570 240.244
R5433 GND.n5461 GND.n1570 240.244
R5434 GND.n5461 GND.n1566 240.244
R5435 GND.n5467 GND.n1566 240.244
R5436 GND.n5467 GND.n1564 240.244
R5437 GND.n5471 GND.n1564 240.244
R5438 GND.n5471 GND.n1560 240.244
R5439 GND.n5477 GND.n1560 240.244
R5440 GND.n5477 GND.n1558 240.244
R5441 GND.n5481 GND.n1558 240.244
R5442 GND.n5481 GND.n1554 240.244
R5443 GND.n5487 GND.n1554 240.244
R5444 GND.n5487 GND.n1552 240.244
R5445 GND.n5491 GND.n1552 240.244
R5446 GND.n5491 GND.n1548 240.244
R5447 GND.n5497 GND.n1548 240.244
R5448 GND.n5497 GND.n1546 240.244
R5449 GND.n5501 GND.n1546 240.244
R5450 GND.n5501 GND.n1542 240.244
R5451 GND.n5507 GND.n1542 240.244
R5452 GND.n5507 GND.n1540 240.244
R5453 GND.n5511 GND.n1540 240.244
R5454 GND.n5511 GND.n1536 240.244
R5455 GND.n5517 GND.n1536 240.244
R5456 GND.n5517 GND.n1534 240.244
R5457 GND.n5521 GND.n1534 240.244
R5458 GND.n5521 GND.n1530 240.244
R5459 GND.n5527 GND.n1530 240.244
R5460 GND.n5527 GND.n1528 240.244
R5461 GND.n5531 GND.n1528 240.244
R5462 GND.n5531 GND.n1524 240.244
R5463 GND.n5537 GND.n1524 240.244
R5464 GND.n5537 GND.n1522 240.244
R5465 GND.n5541 GND.n1522 240.244
R5466 GND.n5541 GND.n1518 240.244
R5467 GND.n5547 GND.n1518 240.244
R5468 GND.n5547 GND.n1516 240.244
R5469 GND.n5551 GND.n1516 240.244
R5470 GND.n5551 GND.n1512 240.244
R5471 GND.n5557 GND.n1512 240.244
R5472 GND.n5557 GND.n1510 240.244
R5473 GND.n5561 GND.n1510 240.244
R5474 GND.n5561 GND.n1506 240.244
R5475 GND.n5567 GND.n1506 240.244
R5476 GND.n5567 GND.n1504 240.244
R5477 GND.n5571 GND.n1504 240.244
R5478 GND.n5571 GND.n1500 240.244
R5479 GND.n5577 GND.n1500 240.244
R5480 GND.n5577 GND.n1498 240.244
R5481 GND.n5581 GND.n1498 240.244
R5482 GND.n5581 GND.n1494 240.244
R5483 GND.n5587 GND.n1494 240.244
R5484 GND.n5587 GND.n1492 240.244
R5485 GND.n5591 GND.n1492 240.244
R5486 GND.n5591 GND.n1488 240.244
R5487 GND.n5597 GND.n1488 240.244
R5488 GND.n5597 GND.n1486 240.244
R5489 GND.n5601 GND.n1486 240.244
R5490 GND.n5601 GND.n1482 240.244
R5491 GND.n5607 GND.n1482 240.244
R5492 GND.n5607 GND.n1480 240.244
R5493 GND.n5611 GND.n1480 240.244
R5494 GND.n5611 GND.n1476 240.244
R5495 GND.n5617 GND.n1476 240.244
R5496 GND.n5617 GND.n1474 240.244
R5497 GND.n5621 GND.n1474 240.244
R5498 GND.n5621 GND.n1470 240.244
R5499 GND.n5627 GND.n1470 240.244
R5500 GND.n5627 GND.n1468 240.244
R5501 GND.n5631 GND.n1468 240.244
R5502 GND.n5631 GND.n1464 240.244
R5503 GND.n5637 GND.n1464 240.244
R5504 GND.n5637 GND.n1462 240.244
R5505 GND.n5641 GND.n1462 240.244
R5506 GND.n5641 GND.n1458 240.244
R5507 GND.n5647 GND.n1458 240.244
R5508 GND.n5647 GND.n1456 240.244
R5509 GND.n5651 GND.n1456 240.244
R5510 GND.n5651 GND.n1452 240.244
R5511 GND.n5657 GND.n1452 240.244
R5512 GND.n5657 GND.n1450 240.244
R5513 GND.n5661 GND.n1450 240.244
R5514 GND.n5661 GND.n1446 240.244
R5515 GND.n5667 GND.n1446 240.244
R5516 GND.n5667 GND.n1444 240.244
R5517 GND.n5671 GND.n1444 240.244
R5518 GND.n5671 GND.n1440 240.244
R5519 GND.n5677 GND.n1440 240.244
R5520 GND.n5677 GND.n1438 240.244
R5521 GND.n5681 GND.n1438 240.244
R5522 GND.n5681 GND.n1434 240.244
R5523 GND.n5687 GND.n1434 240.244
R5524 GND.n5687 GND.n1432 240.244
R5525 GND.n5691 GND.n1432 240.244
R5526 GND.n5691 GND.n1428 240.244
R5527 GND.n5697 GND.n1428 240.244
R5528 GND.n5697 GND.n1426 240.244
R5529 GND.n5701 GND.n1426 240.244
R5530 GND.n5701 GND.n1422 240.244
R5531 GND.n5707 GND.n1422 240.244
R5532 GND.n5707 GND.n1420 240.244
R5533 GND.n5711 GND.n1420 240.244
R5534 GND.n5711 GND.n1416 240.244
R5535 GND.n5717 GND.n1416 240.244
R5536 GND.n5717 GND.n1414 240.244
R5537 GND.n5721 GND.n1414 240.244
R5538 GND.n5721 GND.n1410 240.244
R5539 GND.n5727 GND.n1410 240.244
R5540 GND.n5727 GND.n1408 240.244
R5541 GND.n5731 GND.n1408 240.244
R5542 GND.n5731 GND.n1404 240.244
R5543 GND.n5737 GND.n1404 240.244
R5544 GND.n5737 GND.n1402 240.244
R5545 GND.n5741 GND.n1402 240.244
R5546 GND.n5741 GND.n1398 240.244
R5547 GND.n5747 GND.n1398 240.244
R5548 GND.n5747 GND.n1396 240.244
R5549 GND.n5751 GND.n1396 240.244
R5550 GND.n5751 GND.n1392 240.244
R5551 GND.n5757 GND.n1392 240.244
R5552 GND.n5757 GND.n1390 240.244
R5553 GND.n5761 GND.n1390 240.244
R5554 GND.n5761 GND.n1386 240.244
R5555 GND.n5767 GND.n1386 240.244
R5556 GND.n5767 GND.n1384 240.244
R5557 GND.n5771 GND.n1384 240.244
R5558 GND.n5771 GND.n1380 240.244
R5559 GND.n5777 GND.n1380 240.244
R5560 GND.n5777 GND.n1378 240.244
R5561 GND.n5781 GND.n1378 240.244
R5562 GND.n5781 GND.n1374 240.244
R5563 GND.n5787 GND.n1374 240.244
R5564 GND.n5787 GND.n1372 240.244
R5565 GND.n5791 GND.n1372 240.244
R5566 GND.n5791 GND.n1368 240.244
R5567 GND.n5797 GND.n1368 240.244
R5568 GND.n5797 GND.n1366 240.244
R5569 GND.n5801 GND.n1366 240.244
R5570 GND.n5801 GND.n1362 240.244
R5571 GND.n5807 GND.n1362 240.244
R5572 GND.n5807 GND.n1360 240.244
R5573 GND.n5811 GND.n1360 240.244
R5574 GND.n5811 GND.n1356 240.244
R5575 GND.n5817 GND.n1356 240.244
R5576 GND.n5817 GND.n1354 240.244
R5577 GND.n5821 GND.n1354 240.244
R5578 GND.n5821 GND.n1350 240.244
R5579 GND.n5827 GND.n1350 240.244
R5580 GND.n5827 GND.n1348 240.244
R5581 GND.n5831 GND.n1348 240.244
R5582 GND.n5831 GND.n1344 240.244
R5583 GND.n5837 GND.n1344 240.244
R5584 GND.n5837 GND.n1342 240.244
R5585 GND.n5841 GND.n1342 240.244
R5586 GND.n5841 GND.n1338 240.244
R5587 GND.n5847 GND.n1338 240.244
R5588 GND.n5847 GND.n1336 240.244
R5589 GND.n5851 GND.n1336 240.244
R5590 GND.n5851 GND.n1332 240.244
R5591 GND.n5857 GND.n1332 240.244
R5592 GND.n5857 GND.n1330 240.244
R5593 GND.n5861 GND.n1330 240.244
R5594 GND.n5861 GND.n1326 240.244
R5595 GND.n5867 GND.n1326 240.244
R5596 GND.n5867 GND.n1324 240.244
R5597 GND.n5871 GND.n1324 240.244
R5598 GND.n5871 GND.n1320 240.244
R5599 GND.n5877 GND.n1320 240.244
R5600 GND.n5877 GND.n1318 240.244
R5601 GND.n5881 GND.n1318 240.244
R5602 GND.n5881 GND.n1314 240.244
R5603 GND.n5887 GND.n1314 240.244
R5604 GND.n5887 GND.n1312 240.244
R5605 GND.n5891 GND.n1312 240.244
R5606 GND.n5891 GND.n1308 240.244
R5607 GND.n5897 GND.n1308 240.244
R5608 GND.n5897 GND.n1306 240.244
R5609 GND.n5901 GND.n1306 240.244
R5610 GND.n5901 GND.n1302 240.244
R5611 GND.n5907 GND.n1302 240.244
R5612 GND.n5907 GND.n1300 240.244
R5613 GND.n5911 GND.n1300 240.244
R5614 GND.n5911 GND.n1296 240.244
R5615 GND.n5917 GND.n1296 240.244
R5616 GND.n5917 GND.n1294 240.244
R5617 GND.n5921 GND.n1294 240.244
R5618 GND.n5921 GND.n1290 240.244
R5619 GND.n5927 GND.n1290 240.244
R5620 GND.n5927 GND.n1288 240.244
R5621 GND.n5931 GND.n1288 240.244
R5622 GND.n5931 GND.n1284 240.244
R5623 GND.n5937 GND.n1284 240.244
R5624 GND.n5937 GND.n1282 240.244
R5625 GND.n5941 GND.n1282 240.244
R5626 GND.n5941 GND.n1278 240.244
R5627 GND.n5947 GND.n1278 240.244
R5628 GND.n5947 GND.n1276 240.244
R5629 GND.n5951 GND.n1276 240.244
R5630 GND.n5951 GND.n1272 240.244
R5631 GND.n5957 GND.n1272 240.244
R5632 GND.n5957 GND.n1270 240.244
R5633 GND.n5961 GND.n1270 240.244
R5634 GND.n5961 GND.n1266 240.244
R5635 GND.n5967 GND.n1266 240.244
R5636 GND.n5967 GND.n1264 240.244
R5637 GND.n5971 GND.n1264 240.244
R5638 GND.n5971 GND.n1260 240.244
R5639 GND.n5977 GND.n1260 240.244
R5640 GND.n5977 GND.n1258 240.244
R5641 GND.n5981 GND.n1258 240.244
R5642 GND.n5981 GND.n1254 240.244
R5643 GND.n5987 GND.n1254 240.244
R5644 GND.n5987 GND.n1252 240.244
R5645 GND.n5991 GND.n1252 240.244
R5646 GND.n5991 GND.n1248 240.244
R5647 GND.n5997 GND.n1248 240.244
R5648 GND.n5997 GND.n1246 240.244
R5649 GND.n6001 GND.n1246 240.244
R5650 GND.n6001 GND.n1242 240.244
R5651 GND.n6007 GND.n1242 240.244
R5652 GND.n6007 GND.n1240 240.244
R5653 GND.n6011 GND.n1240 240.244
R5654 GND.n6011 GND.n1236 240.244
R5655 GND.n6017 GND.n1236 240.244
R5656 GND.n6017 GND.n1234 240.244
R5657 GND.n6021 GND.n1234 240.244
R5658 GND.n6021 GND.n1230 240.244
R5659 GND.n6027 GND.n1230 240.244
R5660 GND.n6027 GND.n1228 240.244
R5661 GND.n6031 GND.n1228 240.244
R5662 GND.n6031 GND.n1224 240.244
R5663 GND.n6037 GND.n1224 240.244
R5664 GND.n6037 GND.n1222 240.244
R5665 GND.n6041 GND.n1222 240.244
R5666 GND.n6041 GND.n1218 240.244
R5667 GND.n6047 GND.n1218 240.244
R5668 GND.n6047 GND.n1216 240.244
R5669 GND.n6051 GND.n1216 240.244
R5670 GND.n6051 GND.n1212 240.244
R5671 GND.n6057 GND.n1212 240.244
R5672 GND.n6057 GND.n1210 240.244
R5673 GND.n6061 GND.n1210 240.244
R5674 GND.n6061 GND.n1206 240.244
R5675 GND.n6067 GND.n1206 240.244
R5676 GND.n6067 GND.n1204 240.244
R5677 GND.n6071 GND.n1204 240.244
R5678 GND.n6071 GND.n1200 240.244
R5679 GND.n6077 GND.n1200 240.244
R5680 GND.n6077 GND.n1198 240.244
R5681 GND.n6081 GND.n1198 240.244
R5682 GND.n6081 GND.n1194 240.244
R5683 GND.n6087 GND.n1194 240.244
R5684 GND.n6087 GND.n1192 240.244
R5685 GND.n6091 GND.n1192 240.244
R5686 GND.n6091 GND.n1188 240.244
R5687 GND.n6097 GND.n1188 240.244
R5688 GND.n6097 GND.n1186 240.244
R5689 GND.n6101 GND.n1186 240.244
R5690 GND.n6101 GND.n1182 240.244
R5691 GND.n6107 GND.n1182 240.244
R5692 GND.n6107 GND.n1180 240.244
R5693 GND.n6111 GND.n1180 240.244
R5694 GND.n6111 GND.n1176 240.244
R5695 GND.n6117 GND.n1176 240.244
R5696 GND.n6117 GND.n1174 240.244
R5697 GND.n6121 GND.n1174 240.244
R5698 GND.n6121 GND.n1170 240.244
R5699 GND.n6127 GND.n1170 240.244
R5700 GND.n6127 GND.n1168 240.244
R5701 GND.n6131 GND.n1168 240.244
R5702 GND.n6131 GND.n1164 240.244
R5703 GND.n6137 GND.n1164 240.244
R5704 GND.n6137 GND.n1162 240.244
R5705 GND.n6141 GND.n1162 240.244
R5706 GND.n6141 GND.n1158 240.244
R5707 GND.n6147 GND.n1158 240.244
R5708 GND.n6147 GND.n1156 240.244
R5709 GND.n6151 GND.n1156 240.244
R5710 GND.n6151 GND.n1152 240.244
R5711 GND.n6157 GND.n1152 240.244
R5712 GND.n6157 GND.n1150 240.244
R5713 GND.n6161 GND.n1150 240.244
R5714 GND.n6161 GND.n1146 240.244
R5715 GND.n6167 GND.n1146 240.244
R5716 GND.n6167 GND.n1144 240.244
R5717 GND.n6171 GND.n1144 240.244
R5718 GND.n6171 GND.n1140 240.244
R5719 GND.n6177 GND.n1140 240.244
R5720 GND.n6177 GND.n1138 240.244
R5721 GND.n6181 GND.n1138 240.244
R5722 GND.n6181 GND.n1134 240.244
R5723 GND.n6187 GND.n1134 240.244
R5724 GND.n6187 GND.n1132 240.244
R5725 GND.n6191 GND.n1132 240.244
R5726 GND.n6191 GND.n1128 240.244
R5727 GND.n6197 GND.n1128 240.244
R5728 GND.n6197 GND.n1126 240.244
R5729 GND.n6201 GND.n1126 240.244
R5730 GND.n6201 GND.n1122 240.244
R5731 GND.n6207 GND.n1122 240.244
R5732 GND.n6207 GND.n1120 240.244
R5733 GND.n6211 GND.n1120 240.244
R5734 GND.n6211 GND.n1116 240.244
R5735 GND.n6217 GND.n1116 240.244
R5736 GND.n6217 GND.n1114 240.244
R5737 GND.n6221 GND.n1114 240.244
R5738 GND.n6221 GND.n1110 240.244
R5739 GND.n6227 GND.n1110 240.244
R5740 GND.n6227 GND.n1108 240.244
R5741 GND.n6231 GND.n1108 240.244
R5742 GND.n6231 GND.n1104 240.244
R5743 GND.n6237 GND.n1104 240.244
R5744 GND.n6237 GND.n1102 240.244
R5745 GND.n6241 GND.n1102 240.244
R5746 GND.n6241 GND.n1098 240.244
R5747 GND.n6247 GND.n1098 240.244
R5748 GND.n6247 GND.n1096 240.244
R5749 GND.n6251 GND.n1096 240.244
R5750 GND.n6251 GND.n1092 240.244
R5751 GND.n6257 GND.n1092 240.244
R5752 GND.n6257 GND.n1090 240.244
R5753 GND.n6261 GND.n1090 240.244
R5754 GND.n6261 GND.n1086 240.244
R5755 GND.n6267 GND.n1086 240.244
R5756 GND.n6267 GND.n1084 240.244
R5757 GND.n6271 GND.n1084 240.244
R5758 GND.n6271 GND.n1080 240.244
R5759 GND.n6277 GND.n1080 240.244
R5760 GND.n6277 GND.n1078 240.244
R5761 GND.n6281 GND.n1078 240.244
R5762 GND.n6281 GND.n1074 240.244
R5763 GND.n6287 GND.n1074 240.244
R5764 GND.n6291 GND.n1072 240.244
R5765 GND.n6291 GND.n1068 240.244
R5766 GND.n6297 GND.n1068 240.244
R5767 GND.n6297 GND.n1066 240.244
R5768 GND.n6301 GND.n1066 240.244
R5769 GND.n6301 GND.n1062 240.244
R5770 GND.n6307 GND.n1062 240.244
R5771 GND.n6307 GND.n1060 240.244
R5772 GND.n6311 GND.n1060 240.244
R5773 GND.n6311 GND.n1056 240.244
R5774 GND.n6317 GND.n1056 240.244
R5775 GND.n6317 GND.n1054 240.244
R5776 GND.n6321 GND.n1054 240.244
R5777 GND.n6321 GND.n1050 240.244
R5778 GND.n6327 GND.n1050 240.244
R5779 GND.n6327 GND.n1048 240.244
R5780 GND.n6331 GND.n1048 240.244
R5781 GND.n6331 GND.n1044 240.244
R5782 GND.n6337 GND.n1044 240.244
R5783 GND.n6337 GND.n1042 240.244
R5784 GND.n6341 GND.n1042 240.244
R5785 GND.n6341 GND.n1038 240.244
R5786 GND.n6347 GND.n1038 240.244
R5787 GND.n6347 GND.n1036 240.244
R5788 GND.n6351 GND.n1036 240.244
R5789 GND.n6351 GND.n1032 240.244
R5790 GND.n6357 GND.n1032 240.244
R5791 GND.n6357 GND.n1030 240.244
R5792 GND.n6361 GND.n1030 240.244
R5793 GND.n6361 GND.n1026 240.244
R5794 GND.n6367 GND.n1026 240.244
R5795 GND.n6367 GND.n1024 240.244
R5796 GND.n6371 GND.n1024 240.244
R5797 GND.n6371 GND.n1020 240.244
R5798 GND.n6377 GND.n1020 240.244
R5799 GND.n6377 GND.n1018 240.244
R5800 GND.n6381 GND.n1018 240.244
R5801 GND.n6381 GND.n1014 240.244
R5802 GND.n6387 GND.n1014 240.244
R5803 GND.n6387 GND.n1012 240.244
R5804 GND.n6391 GND.n1012 240.244
R5805 GND.n6391 GND.n1008 240.244
R5806 GND.n6397 GND.n1008 240.244
R5807 GND.n6397 GND.n1006 240.244
R5808 GND.n5322 GND.n5321 240.244
R5809 GND.n5321 GND.n1688 240.244
R5810 GND.n5317 GND.n1688 240.244
R5811 GND.n5317 GND.n1690 240.244
R5812 GND.n5313 GND.n1690 240.244
R5813 GND.n5313 GND.n1697 240.244
R5814 GND.n5309 GND.n1697 240.244
R5815 GND.n5309 GND.n1699 240.244
R5816 GND.n5305 GND.n1699 240.244
R5817 GND.n5305 GND.n1705 240.244
R5818 GND.n5301 GND.n1705 240.244
R5819 GND.n5301 GND.n1707 240.244
R5820 GND.n5297 GND.n1707 240.244
R5821 GND.n5297 GND.n1713 240.244
R5822 GND.n5293 GND.n1713 240.244
R5823 GND.n5293 GND.n1715 240.244
R5824 GND.n5289 GND.n1715 240.244
R5825 GND.n5289 GND.n1721 240.244
R5826 GND.n5285 GND.n1721 240.244
R5827 GND.n5285 GND.n1723 240.244
R5828 GND.n5281 GND.n1723 240.244
R5829 GND.n5281 GND.n1729 240.244
R5830 GND.n5277 GND.n1729 240.244
R5831 GND.n5277 GND.n1731 240.244
R5832 GND.n5273 GND.n1731 240.244
R5833 GND.n5273 GND.n1737 240.244
R5834 GND.n5269 GND.n1737 240.244
R5835 GND.n5269 GND.n1739 240.244
R5836 GND.n5265 GND.n1739 240.244
R5837 GND.n5265 GND.n1745 240.244
R5838 GND.n5261 GND.n1745 240.244
R5839 GND.n5261 GND.n1747 240.244
R5840 GND.n5257 GND.n1747 240.244
R5841 GND.n5257 GND.n1753 240.244
R5842 GND.n5253 GND.n1753 240.244
R5843 GND.n5253 GND.n1755 240.244
R5844 GND.n5249 GND.n1755 240.244
R5845 GND.n5249 GND.n1761 240.244
R5846 GND.n5245 GND.n1761 240.244
R5847 GND.n5245 GND.n1763 240.244
R5848 GND.n5241 GND.n1763 240.244
R5849 GND.n5241 GND.n1769 240.244
R5850 GND.n5237 GND.n1769 240.244
R5851 GND.n5237 GND.n1771 240.244
R5852 GND.n5233 GND.n1771 240.244
R5853 GND.n5233 GND.n1777 240.244
R5854 GND.n5229 GND.n1777 240.244
R5855 GND.n5229 GND.n1779 240.244
R5856 GND.n5225 GND.n1779 240.244
R5857 GND.n5225 GND.n1785 240.244
R5858 GND.n5221 GND.n1785 240.244
R5859 GND.n5221 GND.n1787 240.244
R5860 GND.n5217 GND.n1787 240.244
R5861 GND.n5217 GND.n1793 240.244
R5862 GND.n5213 GND.n1793 240.244
R5863 GND.n5213 GND.n1795 240.244
R5864 GND.n5209 GND.n1795 240.244
R5865 GND.n5209 GND.n1801 240.244
R5866 GND.n5205 GND.n1801 240.244
R5867 GND.n5205 GND.n1803 240.244
R5868 GND.n5201 GND.n1803 240.244
R5869 GND.n5201 GND.n1809 240.244
R5870 GND.n5197 GND.n1809 240.244
R5871 GND.n5197 GND.n1811 240.244
R5872 GND.n5193 GND.n1811 240.244
R5873 GND.n5193 GND.n1817 240.244
R5874 GND.n5189 GND.n1817 240.244
R5875 GND.n5189 GND.n1819 240.244
R5876 GND.n5185 GND.n1819 240.244
R5877 GND.n5185 GND.n1825 240.244
R5878 GND.n5181 GND.n1825 240.244
R5879 GND.n5181 GND.n1827 240.244
R5880 GND.n5177 GND.n1827 240.244
R5881 GND.n5177 GND.n1833 240.244
R5882 GND.n5173 GND.n1833 240.244
R5883 GND.n5173 GND.n1835 240.244
R5884 GND.n5169 GND.n1835 240.244
R5885 GND.n5169 GND.n1841 240.244
R5886 GND.n5165 GND.n1841 240.244
R5887 GND.n5165 GND.n1843 240.244
R5888 GND.n5161 GND.n1843 240.244
R5889 GND.n5161 GND.n1849 240.244
R5890 GND.n5157 GND.n1849 240.244
R5891 GND.n5157 GND.n1851 240.244
R5892 GND.n5153 GND.n1851 240.244
R5893 GND.n5153 GND.n1857 240.244
R5894 GND.n5149 GND.n1857 240.244
R5895 GND.n5149 GND.n1859 240.244
R5896 GND.n5145 GND.n1859 240.244
R5897 GND.n5145 GND.n1865 240.244
R5898 GND.n5141 GND.n1865 240.244
R5899 GND.n5141 GND.n1867 240.244
R5900 GND.n5137 GND.n1867 240.244
R5901 GND.n5137 GND.n1873 240.244
R5902 GND.n2557 GND.n1873 240.244
R5903 GND.n2558 GND.n2557 240.244
R5904 GND.n2559 GND.n2558 240.244
R5905 GND.n2559 GND.n2549 240.244
R5906 GND.n2584 GND.n2549 240.244
R5907 GND.n2584 GND.n2550 240.244
R5908 GND.n2580 GND.n2550 240.244
R5909 GND.n2580 GND.n2579 240.244
R5910 GND.n2579 GND.n2578 240.244
R5911 GND.n2578 GND.n2567 240.244
R5912 GND.n2574 GND.n2567 240.244
R5913 GND.n2574 GND.n2220 240.244
R5914 GND.n2637 GND.n2220 240.244
R5915 GND.n2638 GND.n2637 240.244
R5916 GND.n2638 GND.n2215 240.244
R5917 GND.n2659 GND.n2215 240.244
R5918 GND.n2659 GND.n2216 240.244
R5919 GND.n2655 GND.n2216 240.244
R5920 GND.n2655 GND.n2654 240.244
R5921 GND.n2654 GND.n2649 240.244
R5922 GND.n2649 GND.n2159 240.244
R5923 GND.n2757 GND.n2159 240.244
R5924 GND.n2757 GND.n2160 240.244
R5925 GND.n2752 GND.n2160 240.244
R5926 GND.n2752 GND.n2163 240.244
R5927 GND.n2696 GND.n2163 240.244
R5928 GND.n2740 GND.n2696 240.244
R5929 GND.n2740 GND.n2700 240.244
R5930 GND.n2735 GND.n2700 240.244
R5931 GND.n2735 GND.n2734 240.244
R5932 GND.n2734 GND.n2733 240.244
R5933 GND.n2733 GND.n2705 240.244
R5934 GND.n2727 GND.n2705 240.244
R5935 GND.n2727 GND.n2726 240.244
R5936 GND.n2726 GND.n2725 240.244
R5937 GND.n2725 GND.n2713 240.244
R5938 GND.n2721 GND.n2713 240.244
R5939 GND.n2721 GND.n2094 240.244
R5940 GND.n2824 GND.n2094 240.244
R5941 GND.n2825 GND.n2824 240.244
R5942 GND.n2826 GND.n2825 240.244
R5943 GND.n2826 GND.n2090 240.244
R5944 GND.n2835 GND.n2090 240.244
R5945 GND.n2835 GND.n2064 240.244
R5946 GND.n2910 GND.n2064 240.244
R5947 GND.n2911 GND.n2910 240.244
R5948 GND.n2912 GND.n2911 240.244
R5949 GND.n2912 GND.n2059 240.244
R5950 GND.n4886 GND.n2059 240.244
R5951 GND.n4886 GND.n2060 240.244
R5952 GND.n4882 GND.n2060 240.244
R5953 GND.n4882 GND.n2920 240.244
R5954 GND.n4878 GND.n2920 240.244
R5955 GND.n4878 GND.n2922 240.244
R5956 GND.n4874 GND.n2922 240.244
R5957 GND.n4874 GND.n2928 240.244
R5958 GND.n4864 GND.n2928 240.244
R5959 GND.n4864 GND.n2940 240.244
R5960 GND.n4860 GND.n2940 240.244
R5961 GND.n4860 GND.n2946 240.244
R5962 GND.n3544 GND.n2946 240.244
R5963 GND.n3551 GND.n3544 240.244
R5964 GND.n3551 GND.n2998 240.244
R5965 GND.n4809 GND.n2998 240.244
R5966 GND.n4809 GND.n2999 240.244
R5967 GND.n4805 GND.n2999 240.244
R5968 GND.n4805 GND.n3005 240.244
R5969 GND.n3042 GND.n3005 240.244
R5970 GND.n3042 GND.n3038 240.244
R5971 GND.n4788 GND.n3038 240.244
R5972 GND.n4788 GND.n3039 240.244
R5973 GND.n4784 GND.n3039 240.244
R5974 GND.n4784 GND.n3050 240.244
R5975 GND.n3086 GND.n3050 240.244
R5976 GND.n3086 GND.n3082 240.244
R5977 GND.n4767 GND.n3082 240.244
R5978 GND.n4767 GND.n3083 240.244
R5979 GND.n4763 GND.n3083 240.244
R5980 GND.n4763 GND.n3094 240.244
R5981 GND.n3138 GND.n3094 240.244
R5982 GND.n3139 GND.n3138 240.244
R5983 GND.n3139 GND.n3132 240.244
R5984 GND.n4740 GND.n3132 240.244
R5985 GND.n4740 GND.n3133 240.244
R5986 GND.n4736 GND.n3133 240.244
R5987 GND.n4736 GND.n3147 240.244
R5988 GND.n3333 GND.n3147 240.244
R5989 GND.n3334 GND.n3333 240.244
R5990 GND.n3335 GND.n3334 240.244
R5991 GND.n3335 GND.n3326 240.244
R5992 GND.n3737 GND.n3326 240.244
R5993 GND.n3738 GND.n3737 240.244
R5994 GND.n3739 GND.n3738 240.244
R5995 GND.n3739 GND.n3321 240.244
R5996 GND.n3748 GND.n3321 240.244
R5997 GND.n3748 GND.n3322 240.244
R5998 GND.n3322 GND.n3216 240.244
R5999 GND.n4690 GND.n3216 240.244
R6000 GND.n4690 GND.n3217 240.244
R6001 GND.n4686 GND.n3217 240.244
R6002 GND.n4686 GND.n3223 240.244
R6003 GND.n4676 GND.n3223 240.244
R6004 GND.n4676 GND.n3235 240.244
R6005 GND.n4672 GND.n3235 240.244
R6006 GND.n4672 GND.n3241 240.244
R6007 GND.n4112 GND.n3241 240.244
R6008 GND.n4120 GND.n4112 240.244
R6009 GND.n4120 GND.n4110 240.244
R6010 GND.n4124 GND.n4110 240.244
R6011 GND.n4125 GND.n4124 240.244
R6012 GND.n4125 GND.n4105 240.244
R6013 GND.n4134 GND.n4105 240.244
R6014 GND.n4134 GND.n4106 240.244
R6015 GND.n4106 GND.n3945 240.244
R6016 GND.n4535 GND.n3945 240.244
R6017 GND.n4535 GND.n3946 240.244
R6018 GND.n4531 GND.n3946 240.244
R6019 GND.n4531 GND.n3952 240.244
R6020 GND.n4064 GND.n3952 240.244
R6021 GND.n4070 GND.n4064 240.244
R6022 GND.n4071 GND.n4070 240.244
R6023 GND.n4072 GND.n4071 240.244
R6024 GND.n4072 GND.n4060 240.244
R6025 GND.n4078 GND.n4060 240.244
R6026 GND.n4079 GND.n4078 240.244
R6027 GND.n4080 GND.n4079 240.244
R6028 GND.n4080 GND.n4055 240.244
R6029 GND.n4089 GND.n4055 240.244
R6030 GND.n4089 GND.n4056 240.244
R6031 GND.n4056 GND.n4034 240.244
R6032 GND.n4486 GND.n4034 240.244
R6033 GND.n4486 GND.n4035 240.244
R6034 GND.n4481 GND.n4035 240.244
R6035 GND.n4481 GND.n4038 240.244
R6036 GND.n4377 GND.n4038 240.244
R6037 GND.n4378 GND.n4377 240.244
R6038 GND.n4379 GND.n4378 240.244
R6039 GND.n4379 GND.n4371 240.244
R6040 GND.n4405 GND.n4371 240.244
R6041 GND.n4405 GND.n4372 240.244
R6042 GND.n4400 GND.n4372 240.244
R6043 GND.n4400 GND.n4399 240.244
R6044 GND.n4399 GND.n4398 240.244
R6045 GND.n4398 GND.n4385 240.244
R6046 GND.n4394 GND.n4385 240.244
R6047 GND.n4394 GND.n4393 240.244
R6048 GND.n4393 GND.n797 240.244
R6049 GND.n6610 GND.n797 240.244
R6050 GND.n6610 GND.n798 240.244
R6051 GND.n6606 GND.n798 240.244
R6052 GND.n6606 GND.n6605 240.244
R6053 GND.n6605 GND.n6604 240.244
R6054 GND.n6604 GND.n804 240.244
R6055 GND.n6600 GND.n804 240.244
R6056 GND.n6600 GND.n6599 240.244
R6057 GND.n6599 GND.n6598 240.244
R6058 GND.n6598 GND.n810 240.244
R6059 GND.n6594 GND.n810 240.244
R6060 GND.n6594 GND.n6593 240.244
R6061 GND.n6593 GND.n6592 240.244
R6062 GND.n6592 GND.n816 240.244
R6063 GND.n6587 GND.n816 240.244
R6064 GND.n6587 GND.n822 240.244
R6065 GND.n6583 GND.n822 240.244
R6066 GND.n6583 GND.n825 240.244
R6067 GND.n6579 GND.n825 240.244
R6068 GND.n6579 GND.n831 240.244
R6069 GND.n6575 GND.n831 240.244
R6070 GND.n6575 GND.n833 240.244
R6071 GND.n6571 GND.n833 240.244
R6072 GND.n6571 GND.n839 240.244
R6073 GND.n6567 GND.n839 240.244
R6074 GND.n6567 GND.n841 240.244
R6075 GND.n6563 GND.n841 240.244
R6076 GND.n6563 GND.n847 240.244
R6077 GND.n6559 GND.n847 240.244
R6078 GND.n6559 GND.n849 240.244
R6079 GND.n6555 GND.n849 240.244
R6080 GND.n6555 GND.n855 240.244
R6081 GND.n6551 GND.n855 240.244
R6082 GND.n6551 GND.n857 240.244
R6083 GND.n6547 GND.n857 240.244
R6084 GND.n6547 GND.n863 240.244
R6085 GND.n6543 GND.n863 240.244
R6086 GND.n6543 GND.n865 240.244
R6087 GND.n6539 GND.n865 240.244
R6088 GND.n6539 GND.n871 240.244
R6089 GND.n6535 GND.n871 240.244
R6090 GND.n6535 GND.n873 240.244
R6091 GND.n6531 GND.n873 240.244
R6092 GND.n6531 GND.n879 240.244
R6093 GND.n6527 GND.n879 240.244
R6094 GND.n6527 GND.n881 240.244
R6095 GND.n6523 GND.n881 240.244
R6096 GND.n6523 GND.n887 240.244
R6097 GND.n6519 GND.n887 240.244
R6098 GND.n6519 GND.n889 240.244
R6099 GND.n6515 GND.n889 240.244
R6100 GND.n6515 GND.n895 240.244
R6101 GND.n6511 GND.n895 240.244
R6102 GND.n6511 GND.n897 240.244
R6103 GND.n6507 GND.n897 240.244
R6104 GND.n6507 GND.n903 240.244
R6105 GND.n6503 GND.n903 240.244
R6106 GND.n6503 GND.n905 240.244
R6107 GND.n6499 GND.n905 240.244
R6108 GND.n6499 GND.n911 240.244
R6109 GND.n6495 GND.n911 240.244
R6110 GND.n6495 GND.n913 240.244
R6111 GND.n6491 GND.n913 240.244
R6112 GND.n6491 GND.n919 240.244
R6113 GND.n6487 GND.n919 240.244
R6114 GND.n6487 GND.n921 240.244
R6115 GND.n6483 GND.n921 240.244
R6116 GND.n6483 GND.n927 240.244
R6117 GND.n6479 GND.n927 240.244
R6118 GND.n6479 GND.n929 240.244
R6119 GND.n6475 GND.n929 240.244
R6120 GND.n6475 GND.n935 240.244
R6121 GND.n6471 GND.n935 240.244
R6122 GND.n6471 GND.n937 240.244
R6123 GND.n6467 GND.n937 240.244
R6124 GND.n6467 GND.n943 240.244
R6125 GND.n6463 GND.n943 240.244
R6126 GND.n6463 GND.n945 240.244
R6127 GND.n6459 GND.n945 240.244
R6128 GND.n6459 GND.n951 240.244
R6129 GND.n6455 GND.n951 240.244
R6130 GND.n6455 GND.n953 240.244
R6131 GND.n6451 GND.n953 240.244
R6132 GND.n6451 GND.n959 240.244
R6133 GND.n6447 GND.n959 240.244
R6134 GND.n6447 GND.n961 240.244
R6135 GND.n6443 GND.n961 240.244
R6136 GND.n6443 GND.n967 240.244
R6137 GND.n6439 GND.n967 240.244
R6138 GND.n6439 GND.n969 240.244
R6139 GND.n6435 GND.n969 240.244
R6140 GND.n6435 GND.n975 240.244
R6141 GND.n6431 GND.n975 240.244
R6142 GND.n6431 GND.n977 240.244
R6143 GND.n6427 GND.n977 240.244
R6144 GND.n6427 GND.n983 240.244
R6145 GND.n6423 GND.n983 240.244
R6146 GND.n6423 GND.n985 240.244
R6147 GND.n6419 GND.n985 240.244
R6148 GND.n6419 GND.n991 240.244
R6149 GND.n6415 GND.n991 240.244
R6150 GND.n6415 GND.n993 240.244
R6151 GND.n6411 GND.n993 240.244
R6152 GND.n6411 GND.n999 240.244
R6153 GND.n6407 GND.n999 240.244
R6154 GND.n6407 GND.n1001 240.244
R6155 GND.n5417 GND.n1596 240.244
R6156 GND.n5413 GND.n1596 240.244
R6157 GND.n5413 GND.n1601 240.244
R6158 GND.n5409 GND.n1601 240.244
R6159 GND.n5409 GND.n1603 240.244
R6160 GND.n5405 GND.n1603 240.244
R6161 GND.n5405 GND.n1609 240.244
R6162 GND.n5401 GND.n1609 240.244
R6163 GND.n5401 GND.n1611 240.244
R6164 GND.n5397 GND.n1611 240.244
R6165 GND.n5397 GND.n1617 240.244
R6166 GND.n5393 GND.n1617 240.244
R6167 GND.n5393 GND.n1619 240.244
R6168 GND.n5389 GND.n1619 240.244
R6169 GND.n5389 GND.n1625 240.244
R6170 GND.n5385 GND.n1625 240.244
R6171 GND.n5385 GND.n1627 240.244
R6172 GND.n5381 GND.n1627 240.244
R6173 GND.n5381 GND.n1633 240.244
R6174 GND.n5377 GND.n1633 240.244
R6175 GND.n5377 GND.n1635 240.244
R6176 GND.n5373 GND.n1635 240.244
R6177 GND.n5373 GND.n1641 240.244
R6178 GND.n5369 GND.n1641 240.244
R6179 GND.n5369 GND.n1643 240.244
R6180 GND.n5365 GND.n1643 240.244
R6181 GND.n5365 GND.n1649 240.244
R6182 GND.n5361 GND.n1649 240.244
R6183 GND.n5361 GND.n1651 240.244
R6184 GND.n5357 GND.n1651 240.244
R6185 GND.n5357 GND.n1657 240.244
R6186 GND.n5353 GND.n1657 240.244
R6187 GND.n5353 GND.n1659 240.244
R6188 GND.n5349 GND.n1659 240.244
R6189 GND.n5349 GND.n1665 240.244
R6190 GND.n5345 GND.n1665 240.244
R6191 GND.n5345 GND.n1667 240.244
R6192 GND.n5341 GND.n1667 240.244
R6193 GND.n5341 GND.n1673 240.244
R6194 GND.n5337 GND.n1673 240.244
R6195 GND.n5337 GND.n1675 240.244
R6196 GND.n5333 GND.n1675 240.244
R6197 GND.n5333 GND.n1681 240.244
R6198 GND.n5328 GND.n1681 240.244
R6199 GND.n2511 GND.n2278 240.244
R6200 GND.n2515 GND.n2513 240.244
R6201 GND.n2521 GND.n2274 240.244
R6202 GND.n2525 GND.n2523 240.244
R6203 GND.n2531 GND.n2270 240.244
R6204 GND.n2534 GND.n2533 240.244
R6205 GND.n1890 GND.n1878 240.244
R6206 GND.n5127 GND.n1890 240.244
R6207 GND.n5127 GND.n1891 240.244
R6208 GND.n2589 GND.n1891 240.244
R6209 GND.n2589 GND.n2588 240.244
R6210 GND.n2588 GND.n2255 240.244
R6211 GND.n2255 GND.n2245 240.244
R6212 GND.n2610 GND.n2245 240.244
R6213 GND.n2613 GND.n2610 240.244
R6214 GND.n2613 GND.n2612 240.244
R6215 GND.n2612 GND.n2233 240.244
R6216 GND.n2233 GND.n2231 240.244
R6217 GND.n2231 GND.n2210 240.244
R6218 GND.n2663 GND.n2210 240.244
R6219 GND.n2663 GND.n2662 240.244
R6220 GND.n2662 GND.n2211 240.244
R6221 GND.n2211 GND.n2199 240.244
R6222 GND.n2650 GND.n2199 240.244
R6223 GND.n2650 GND.n2154 240.244
R6224 GND.n2761 GND.n2154 240.244
R6225 GND.n2761 GND.n2760 240.244
R6226 GND.n2760 GND.n2155 240.244
R6227 GND.n2169 GND.n2155 240.244
R6228 GND.n2170 GND.n2169 240.244
R6229 GND.n2744 GND.n2170 240.244
R6230 GND.n2744 GND.n2743 240.244
R6231 GND.n2743 GND.n2182 240.244
R6232 GND.n2697 GND.n2182 240.244
R6233 GND.n2697 GND.n2137 240.244
R6234 GND.n2137 GND.n2126 240.244
R6235 GND.n2783 GND.n2126 240.244
R6236 GND.n2787 GND.n2783 240.244
R6237 GND.n2787 GND.n2786 240.244
R6238 GND.n2786 GND.n2116 240.244
R6239 GND.n2116 GND.n2107 240.244
R6240 GND.n2811 GND.n2107 240.244
R6241 GND.n2813 GND.n2811 240.244
R6242 GND.n2813 GND.n2812 240.244
R6243 GND.n2812 GND.n2083 240.244
R6244 GND.n2892 GND.n2083 240.244
R6245 GND.n2893 GND.n2892 240.244
R6246 GND.n2893 GND.n2068 240.244
R6247 GND.n2905 GND.n2068 240.244
R6248 GND.n2906 GND.n2905 240.244
R6249 GND.n2907 GND.n2906 240.244
R6250 GND.n2907 GND.n1989 240.244
R6251 GND.n2852 GND.n2851 240.244
R6252 GND.n2855 GND.n2854 240.244
R6253 GND.n2862 GND.n2861 240.244
R6254 GND.n2865 GND.n2864 240.244
R6255 GND.n2874 GND.n2873 240.244
R6256 GND.n2541 GND.n1876 240.244
R6257 GND.n2541 GND.n1888 240.244
R6258 GND.n2263 GND.n1888 240.244
R6259 GND.n2548 GND.n2263 240.244
R6260 GND.n2548 GND.n2252 240.244
R6261 GND.n2601 GND.n2252 240.244
R6262 GND.n2601 GND.n2247 240.244
R6263 GND.n2608 GND.n2247 240.244
R6264 GND.n2608 GND.n2242 240.244
R6265 GND.n2242 GND.n2228 240.244
R6266 GND.n2625 GND.n2228 240.244
R6267 GND.n2625 GND.n2223 240.244
R6268 GND.n2634 GND.n2223 240.244
R6269 GND.n2634 GND.n2208 240.244
R6270 GND.n2213 GND.n2208 240.244
R6271 GND.n2213 GND.n2194 240.244
R6272 GND.n2674 GND.n2194 240.244
R6273 GND.n2674 GND.n2195 240.244
R6274 GND.n2195 GND.n2191 240.244
R6275 GND.n2191 GND.n2151 240.244
R6276 GND.n2157 GND.n2151 240.244
R6277 GND.n2187 GND.n2157 240.244
R6278 GND.n2188 GND.n2187 240.244
R6279 GND.n2188 GND.n2166 240.244
R6280 GND.n2179 GND.n2166 240.244
R6281 GND.n2183 GND.n2179 240.244
R6282 GND.n2692 GND.n2183 240.244
R6283 GND.n2692 GND.n2133 240.244
R6284 GND.n2774 GND.n2133 240.244
R6285 GND.n2774 GND.n2128 240.244
R6286 GND.n2781 GND.n2128 240.244
R6287 GND.n2781 GND.n2124 240.244
R6288 GND.n2124 GND.n2113 240.244
R6289 GND.n2799 GND.n2113 240.244
R6290 GND.n2799 GND.n2108 240.244
R6291 GND.n2809 GND.n2108 240.244
R6292 GND.n2809 GND.n2104 240.244
R6293 GND.n2803 GND.n2104 240.244
R6294 GND.n2803 GND.n2085 240.244
R6295 GND.n2890 GND.n2085 240.244
R6296 GND.n2890 GND.n2080 240.244
R6297 GND.n2838 GND.n2080 240.244
R6298 GND.n2838 GND.n2070 240.244
R6299 GND.n2839 GND.n2070 240.244
R6300 GND.n2839 GND.n2067 240.244
R6301 GND.n2067 GND.n1987 240.244
R6302 GND.n3428 GND.n3427 240.132
R6303 GND.n3426 GND.n3425 240.132
R6304 GND.n3272 GND.n3271 240.132
R6305 GND.n3270 GND.n3269 240.132
R6306 GND.n2979 GND.t194 226.101
R6307 GND.n3757 GND.t98 226.101
R6308 GND.n3407 GND.t154 210.121
R6309 GND.n3399 GND.t134 210.121
R6310 GND.n3299 GND.t169 210.121
R6311 GND.n3290 GND.t188 210.121
R6312 GND.n5011 GND.n5010 199.319
R6313 GND.n2871 GND.t123 191.03
R6314 GND.n2006 GND.t211 191.03
R6315 GND.n2024 GND.t132 191.03
R6316 GND.n4900 GND.t161 191.03
R6317 GND.n4926 GND.t126 191.03
R6318 GND.n4953 GND.t174 191.03
R6319 GND.n4561 GND.t159 191.03
R6320 GND.n4576 GND.t233 191.03
R6321 GND.n4161 GND.t218 191.03
R6322 GND.n4194 GND.t150 191.03
R6323 GND.n4136 GND.t193 191.03
R6324 GND.n758 GND.t142 191.03
R6325 GND.n6699 GND.t113 191.03
R6326 GND.n6723 GND.t208 191.03
R6327 GND.n691 GND.t129 191.03
R6328 GND.n668 GND.t214 191.03
R6329 GND.n780 GND.t110 191.03
R6330 GND.n4242 GND.t147 191.03
R6331 GND.n2367 GND.t140 191.03
R6332 GND.n2399 GND.t221 191.03
R6333 GND.n2431 GND.t230 191.03
R6334 GND.n2464 GND.t203 191.03
R6335 GND.n2281 GND.t91 191.03
R6336 GND.n2267 GND.t200 191.03
R6337 GND.n3429 GND.n3423 186.49
R6338 GND.n3273 GND.n3267 186.49
R6339 GND.n234 GND.n233 185
R6340 GND.n232 GND.n231 185
R6341 GND.n223 GND.n222 185
R6342 GND.n226 GND.n225 185
R6343 GND.n257 GND.n256 185
R6344 GND.n255 GND.n254 185
R6345 GND.n246 GND.n245 185
R6346 GND.n249 GND.n248 185
R6347 GND.n190 GND.n189 185
R6348 GND.n188 GND.n187 185
R6349 GND.n179 GND.n178 185
R6350 GND.n182 GND.n181 185
R6351 GND.n213 GND.n212 185
R6352 GND.n211 GND.n210 185
R6353 GND.n202 GND.n201 185
R6354 GND.n205 GND.n204 185
R6355 GND.n146 GND.n145 185
R6356 GND.n144 GND.n143 185
R6357 GND.n135 GND.n134 185
R6358 GND.n138 GND.n137 185
R6359 GND.n169 GND.n168 185
R6360 GND.n167 GND.n166 185
R6361 GND.n158 GND.n157 185
R6362 GND.n161 GND.n160 185
R6363 GND.n102 GND.n101 185
R6364 GND.n100 GND.n99 185
R6365 GND.n91 GND.n90 185
R6366 GND.n94 GND.n93 185
R6367 GND.n125 GND.n124 185
R6368 GND.n123 GND.n122 185
R6369 GND.n114 GND.n113 185
R6370 GND.n117 GND.n116 185
R6371 GND.n58 GND.n57 185
R6372 GND.n56 GND.n55 185
R6373 GND.n47 GND.n46 185
R6374 GND.n50 GND.n49 185
R6375 GND.n81 GND.n80 185
R6376 GND.n79 GND.n78 185
R6377 GND.n70 GND.n69 185
R6378 GND.n73 GND.n72 185
R6379 GND.n15 GND.n14 185
R6380 GND.n13 GND.n12 185
R6381 GND.n4 GND.n3 185
R6382 GND.n7 GND.n6 185
R6383 GND.n38 GND.n37 185
R6384 GND.n36 GND.n35 185
R6385 GND.n27 GND.n26 185
R6386 GND.n30 GND.n29 185
R6387 GND.n521 GND.n520 185
R6388 GND.n519 GND.n518 185
R6389 GND.n510 GND.n509 185
R6390 GND.n513 GND.n512 185
R6391 GND.n498 GND.n497 185
R6392 GND.n496 GND.n495 185
R6393 GND.n487 GND.n486 185
R6394 GND.n490 GND.n489 185
R6395 GND.n477 GND.n476 185
R6396 GND.n475 GND.n474 185
R6397 GND.n466 GND.n465 185
R6398 GND.n469 GND.n468 185
R6399 GND.n454 GND.n453 185
R6400 GND.n452 GND.n451 185
R6401 GND.n443 GND.n442 185
R6402 GND.n446 GND.n445 185
R6403 GND.n433 GND.n432 185
R6404 GND.n431 GND.n430 185
R6405 GND.n422 GND.n421 185
R6406 GND.n425 GND.n424 185
R6407 GND.n410 GND.n409 185
R6408 GND.n408 GND.n407 185
R6409 GND.n399 GND.n398 185
R6410 GND.n402 GND.n401 185
R6411 GND.n389 GND.n388 185
R6412 GND.n387 GND.n386 185
R6413 GND.n378 GND.n377 185
R6414 GND.n381 GND.n380 185
R6415 GND.n366 GND.n365 185
R6416 GND.n364 GND.n363 185
R6417 GND.n355 GND.n354 185
R6418 GND.n358 GND.n357 185
R6419 GND.n345 GND.n344 185
R6420 GND.n343 GND.n342 185
R6421 GND.n334 GND.n333 185
R6422 GND.n337 GND.n336 185
R6423 GND.n322 GND.n321 185
R6424 GND.n320 GND.n319 185
R6425 GND.n311 GND.n310 185
R6426 GND.n314 GND.n313 185
R6427 GND.n302 GND.n301 185
R6428 GND.n300 GND.n299 185
R6429 GND.n291 GND.n290 185
R6430 GND.n294 GND.n293 185
R6431 GND.n279 GND.n278 185
R6432 GND.n277 GND.n276 185
R6433 GND.n268 GND.n267 185
R6434 GND.n271 GND.n270 185
R6435 GND.n3399 GND.t137 184.131
R6436 GND.n3299 GND.t171 184.131
R6437 GND.n3407 GND.t156 184.13
R6438 GND.n3290 GND.t189 184.13
R6439 GND.n4664 GND.n4663 163.367
R6440 GND.n4661 GND.n3283 163.367
R6441 GND.n4657 GND.n4656 163.367
R6442 GND.n4654 GND.n3286 163.367
R6443 GND.n4650 GND.n4649 163.367
R6444 GND.n4647 GND.n3289 163.367
R6445 GND.n4642 GND.n4641 163.367
R6446 GND.n4639 GND.n3294 163.367
R6447 GND.n3877 GND.n3876 163.367
R6448 GND.n3874 GND.n3298 163.367
R6449 GND.n3869 GND.n3868 163.367
R6450 GND.n3866 GND.n3303 163.367
R6451 GND.n3862 GND.n3861 163.367
R6452 GND.n3859 GND.n3306 163.367
R6453 GND.n3855 GND.n3854 163.367
R6454 GND.n3852 GND.n3309 163.367
R6455 GND.n3520 GND.n2931 163.367
R6456 GND.n3524 GND.n2931 163.367
R6457 GND.n3524 GND.n2938 163.367
R6458 GND.n3528 GND.n2938 163.367
R6459 GND.n3533 GND.n3528 163.367
R6460 GND.n3534 GND.n3533 163.367
R6461 GND.n3534 GND.n2948 163.367
R6462 GND.n3537 GND.n2948 163.367
R6463 GND.n3537 GND.n2956 163.367
R6464 GND.n3541 GND.n2956 163.367
R6465 GND.n3554 GND.n3541 163.367
R6466 GND.n3554 GND.n2988 163.367
R6467 GND.n3558 GND.n2988 163.367
R6468 GND.n3558 GND.n2996 163.367
R6469 GND.n3389 GND.n2996 163.367
R6470 GND.n3566 GND.n3389 163.367
R6471 GND.n3566 GND.n3390 163.367
R6472 GND.n3562 GND.n3390 163.367
R6473 GND.n3562 GND.n3380 163.367
R6474 GND.n3617 GND.n3380 163.367
R6475 GND.n3617 GND.n3028 163.367
R6476 GND.n3621 GND.n3028 163.367
R6477 GND.n3621 GND.n3036 163.367
R6478 GND.n3625 GND.n3036 163.367
R6479 GND.n3629 GND.n3625 163.367
R6480 GND.n3629 GND.n3052 163.367
R6481 GND.n3633 GND.n3052 163.367
R6482 GND.n3633 GND.n3060 163.367
R6483 GND.n3377 GND.n3060 163.367
R6484 GND.n3641 GND.n3377 163.367
R6485 GND.n3641 GND.n3378 163.367
R6486 GND.n3637 GND.n3378 163.367
R6487 GND.n3637 GND.n3371 163.367
R6488 GND.n3653 GND.n3371 163.367
R6489 GND.n3653 GND.n3096 163.367
R6490 GND.n3657 GND.n3096 163.367
R6491 GND.n3657 GND.n3104 163.367
R6492 GND.n3369 GND.n3104 163.367
R6493 GND.n3671 GND.n3369 163.367
R6494 GND.n3671 GND.n3122 163.367
R6495 GND.n3667 GND.n3122 163.367
R6496 GND.n3667 GND.n3130 163.367
R6497 GND.n3663 GND.n3130 163.367
R6498 GND.n3663 GND.n3362 163.367
R6499 GND.n3362 GND.n3357 163.367
R6500 GND.n3693 GND.n3357 163.367
R6501 GND.n3693 GND.n3355 163.367
R6502 GND.n3697 GND.n3355 163.367
R6503 GND.n3697 GND.n3165 163.367
R6504 GND.n3710 GND.n3165 163.367
R6505 GND.n3710 GND.n3173 163.367
R6506 GND.n3714 GND.n3173 163.367
R6507 GND.n3715 GND.n3714 163.367
R6508 GND.n3716 GND.n3715 163.367
R6509 GND.n3716 GND.n3185 163.367
R6510 GND.n3727 GND.n3185 163.367
R6511 GND.n3727 GND.n3193 163.367
R6512 GND.n3723 GND.n3193 163.367
R6513 GND.n3723 GND.n3722 163.367
R6514 GND.n3722 GND.n3721 163.367
R6515 GND.n3721 GND.n3205 163.367
R6516 GND.n3817 GND.n3205 163.367
R6517 GND.n3817 GND.n3213 163.367
R6518 GND.n3214 GND.n3213 163.367
R6519 GND.n3822 GND.n3214 163.367
R6520 GND.n3830 GND.n3822 163.367
R6521 GND.n3831 GND.n3830 163.367
R6522 GND.n3831 GND.n3225 163.367
R6523 GND.n3834 GND.n3225 163.367
R6524 GND.n3834 GND.n3233 163.367
R6525 GND.n3838 GND.n3233 163.367
R6526 GND.n3843 GND.n3838 163.367
R6527 GND.n3844 GND.n3843 163.367
R6528 GND.n3844 GND.n3243 163.367
R6529 GND.n3453 GND.n3415 163.367
R6530 GND.n3457 GND.n3415 163.367
R6531 GND.n3461 GND.n3459 163.367
R6532 GND.n3465 GND.n3413 163.367
R6533 GND.n3469 GND.n3467 163.367
R6534 GND.n3473 GND.n3411 163.367
R6535 GND.n3477 GND.n3475 163.367
R6536 GND.n3481 GND.n3406 163.367
R6537 GND.n3484 GND.n3483 163.367
R6538 GND.n3488 GND.n3486 163.367
R6539 GND.n3492 GND.n3403 163.367
R6540 GND.n3496 GND.n3494 163.367
R6541 GND.n3500 GND.n3398 163.367
R6542 GND.n3504 GND.n3502 163.367
R6543 GND.n3508 GND.n3396 163.367
R6544 GND.n3512 GND.n3510 163.367
R6545 GND.n3516 GND.n3394 163.367
R6546 GND.n3519 GND.n3518 163.367
R6547 GND.n4871 GND.n2932 163.367
R6548 GND.n4871 GND.n2933 163.367
R6549 GND.n4867 GND.n2933 163.367
R6550 GND.n4867 GND.n2936 163.367
R6551 GND.n3531 GND.n2936 163.367
R6552 GND.n3531 GND.n2950 163.367
R6553 GND.n4858 GND.n2950 163.367
R6554 GND.n4858 GND.n2951 163.367
R6555 GND.n4854 GND.n2951 163.367
R6556 GND.n4854 GND.n2954 163.367
R6557 GND.n2990 GND.n2954 163.367
R6558 GND.n4816 GND.n2990 163.367
R6559 GND.n4816 GND.n2991 163.367
R6560 GND.n4812 GND.n2991 163.367
R6561 GND.n4812 GND.n2994 163.367
R6562 GND.n3574 GND.n2994 163.367
R6563 GND.n3574 GND.n3567 163.367
R6564 GND.n3570 GND.n3567 163.367
R6565 GND.n3570 GND.n3569 163.367
R6566 GND.n3569 GND.n3030 163.367
R6567 GND.n4795 GND.n3030 163.367
R6568 GND.n4795 GND.n3031 163.367
R6569 GND.n4791 GND.n3031 163.367
R6570 GND.n4791 GND.n3034 163.367
R6571 GND.n3054 GND.n3034 163.367
R6572 GND.n4781 GND.n3054 163.367
R6573 GND.n4781 GND.n3055 163.367
R6574 GND.n4777 GND.n3055 163.367
R6575 GND.n4777 GND.n3058 163.367
R6576 GND.n3644 GND.n3058 163.367
R6577 GND.n3645 GND.n3644 163.367
R6578 GND.n3645 GND.n3373 163.367
R6579 GND.n3649 GND.n3373 163.367
R6580 GND.n3649 GND.n3098 163.367
R6581 GND.n4760 GND.n3098 163.367
R6582 GND.n4760 GND.n3099 163.367
R6583 GND.n4756 GND.n3099 163.367
R6584 GND.n4756 GND.n3102 163.367
R6585 GND.n3124 GND.n3102 163.367
R6586 GND.n4747 GND.n3124 163.367
R6587 GND.n4747 GND.n3125 163.367
R6588 GND.n4743 GND.n3125 163.367
R6589 GND.n4743 GND.n3128 163.367
R6590 GND.n3686 GND.n3128 163.367
R6591 GND.n3686 GND.n3359 163.367
R6592 GND.n3691 GND.n3359 163.367
R6593 GND.n3691 GND.n3360 163.367
R6594 GND.n3360 GND.n3167 163.367
R6595 GND.n4726 GND.n3167 163.367
R6596 GND.n4726 GND.n3168 163.367
R6597 GND.n4722 GND.n3168 163.367
R6598 GND.n4722 GND.n3171 163.367
R6599 GND.n3343 GND.n3171 163.367
R6600 GND.n3343 GND.n3187 163.367
R6601 GND.n4712 GND.n3187 163.367
R6602 GND.n4712 GND.n3188 163.367
R6603 GND.n4708 GND.n3188 163.367
R6604 GND.n4708 GND.n3191 163.367
R6605 GND.n3318 GND.n3191 163.367
R6606 GND.n3318 GND.n3207 163.367
R6607 GND.n4698 GND.n3207 163.367
R6608 GND.n4698 GND.n3208 163.367
R6609 GND.n4694 GND.n3208 163.367
R6610 GND.n4694 GND.n3211 163.367
R6611 GND.n3825 GND.n3211 163.367
R6612 GND.n3828 GND.n3825 163.367
R6613 GND.n3828 GND.n3227 163.367
R6614 GND.n4683 GND.n3227 163.367
R6615 GND.n4683 GND.n3228 163.367
R6616 GND.n4679 GND.n3228 163.367
R6617 GND.n4679 GND.n3231 163.367
R6618 GND.n3841 GND.n3231 163.367
R6619 GND.n3841 GND.n3245 163.367
R6620 GND.n4669 GND.n3245 163.367
R6621 GND.n3279 GND.n3278 154.327
R6622 GND.n3254 GND.t179 152.625
R6623 GND.n3434 GND.n3433 152
R6624 GND.n3435 GND.n3421 152
R6625 GND.n3437 GND.n3436 152
R6626 GND.n3441 GND.n3440 152
R6627 GND.n3442 GND.n3418 152
R6628 GND.n3444 GND.n3443 152
R6629 GND.n3446 GND.n3416 152
R6630 GND.n3448 GND.n3447 152
R6631 GND.n3277 GND.n3248 152
R6632 GND.n3266 GND.n3249 152
R6633 GND.n3265 GND.n3264 152
R6634 GND.n3263 GND.n3250 152
R6635 GND.n3259 GND.n3258 152
R6636 GND.n3257 GND.n3252 152
R6637 GND.n3256 GND.n3255 152
R6638 GND.n2979 GND.t197 151.412
R6639 GND.n3757 GND.t100 151.412
R6640 GND.t17 GND.n224 147.888
R6641 GND.t53 GND.n247 147.888
R6642 GND.t52 GND.n180 147.888
R6643 GND.t87 GND.n203 147.888
R6644 GND.t19 GND.n136 147.888
R6645 GND.t64 GND.n159 147.888
R6646 GND.t47 GND.n92 147.888
R6647 GND.t55 GND.n115 147.888
R6648 GND.t71 GND.n48 147.888
R6649 GND.t42 GND.n71 147.888
R6650 GND.t33 GND.n5 147.888
R6651 GND.t82 GND.n28 147.888
R6652 GND.t26 GND.n511 147.888
R6653 GND.t65 GND.n488 147.888
R6654 GND.t56 GND.n467 147.888
R6655 GND.t5 GND.n444 147.888
R6656 GND.t28 GND.n423 147.888
R6657 GND.t66 GND.n400 147.888
R6658 GND.t58 GND.n379 147.888
R6659 GND.t63 GND.n356 147.888
R6660 GND.t50 GND.n335 147.888
R6661 GND.t18 GND.n312 147.888
R6662 GND.t7 GND.n292 147.888
R6663 GND.t69 GND.n269 147.888
R6664 GND.n3879 GND.n3296 143.351
R6665 GND.n3879 GND.n3878 143.351
R6666 GND.n2872 GND.t124 141.769
R6667 GND.n2007 GND.t212 141.769
R6668 GND.n2025 GND.t133 141.769
R6669 GND.n4901 GND.t162 141.769
R6670 GND.n4927 GND.t127 141.769
R6671 GND.n4954 GND.t175 141.769
R6672 GND.n4562 GND.t158 141.769
R6673 GND.n4577 GND.t232 141.769
R6674 GND.n4162 GND.t217 141.769
R6675 GND.n4195 GND.t149 141.769
R6676 GND.n4137 GND.t192 141.769
R6677 GND.n759 GND.t143 141.769
R6678 GND.n6700 GND.t114 141.769
R6679 GND.n6724 GND.t209 141.769
R6680 GND.n692 GND.t130 141.769
R6681 GND.n669 GND.t215 141.769
R6682 GND.n781 GND.t111 141.769
R6683 GND.n4243 GND.t146 141.769
R6684 GND.n2368 GND.t139 141.769
R6685 GND.n2400 GND.t220 141.769
R6686 GND.n2432 GND.t229 141.769
R6687 GND.n2465 GND.t202 141.769
R6688 GND.n2282 GND.t90 141.769
R6689 GND.n2268 GND.t199 141.769
R6690 GND.n3431 GND.t95 134.386
R6691 GND.n3447 GND.t185 126.766
R6692 GND.n3445 GND.t105 126.766
R6693 GND.n3418 GND.t166 126.766
R6694 GND.n3439 GND.t222 126.766
R6695 GND.n3438 GND.t204 126.766
R6696 GND.n3421 GND.t115 126.766
R6697 GND.n3432 GND.t176 126.766
R6698 GND.n3253 GND.t92 126.766
R6699 GND.n3257 GND.t151 126.766
R6700 GND.n3251 GND.t225 126.766
R6701 GND.n3262 GND.t163 126.766
R6702 GND.n3264 GND.t102 126.766
R6703 GND.n3276 GND.t182 126.766
R6704 GND.n3278 GND.t118 126.766
R6705 GND.n233 GND.n232 104.615
R6706 GND.n232 GND.n222 104.615
R6707 GND.n225 GND.n222 104.615
R6708 GND.n256 GND.n255 104.615
R6709 GND.n255 GND.n245 104.615
R6710 GND.n248 GND.n245 104.615
R6711 GND.n189 GND.n188 104.615
R6712 GND.n188 GND.n178 104.615
R6713 GND.n181 GND.n178 104.615
R6714 GND.n212 GND.n211 104.615
R6715 GND.n211 GND.n201 104.615
R6716 GND.n204 GND.n201 104.615
R6717 GND.n145 GND.n144 104.615
R6718 GND.n144 GND.n134 104.615
R6719 GND.n137 GND.n134 104.615
R6720 GND.n168 GND.n167 104.615
R6721 GND.n167 GND.n157 104.615
R6722 GND.n160 GND.n157 104.615
R6723 GND.n101 GND.n100 104.615
R6724 GND.n100 GND.n90 104.615
R6725 GND.n93 GND.n90 104.615
R6726 GND.n124 GND.n123 104.615
R6727 GND.n123 GND.n113 104.615
R6728 GND.n116 GND.n113 104.615
R6729 GND.n57 GND.n56 104.615
R6730 GND.n56 GND.n46 104.615
R6731 GND.n49 GND.n46 104.615
R6732 GND.n80 GND.n79 104.615
R6733 GND.n79 GND.n69 104.615
R6734 GND.n72 GND.n69 104.615
R6735 GND.n14 GND.n13 104.615
R6736 GND.n13 GND.n3 104.615
R6737 GND.n6 GND.n3 104.615
R6738 GND.n37 GND.n36 104.615
R6739 GND.n36 GND.n26 104.615
R6740 GND.n29 GND.n26 104.615
R6741 GND.n520 GND.n519 104.615
R6742 GND.n519 GND.n509 104.615
R6743 GND.n512 GND.n509 104.615
R6744 GND.n497 GND.n496 104.615
R6745 GND.n496 GND.n486 104.615
R6746 GND.n489 GND.n486 104.615
R6747 GND.n476 GND.n475 104.615
R6748 GND.n475 GND.n465 104.615
R6749 GND.n468 GND.n465 104.615
R6750 GND.n453 GND.n452 104.615
R6751 GND.n452 GND.n442 104.615
R6752 GND.n445 GND.n442 104.615
R6753 GND.n432 GND.n431 104.615
R6754 GND.n431 GND.n421 104.615
R6755 GND.n424 GND.n421 104.615
R6756 GND.n409 GND.n408 104.615
R6757 GND.n408 GND.n398 104.615
R6758 GND.n401 GND.n398 104.615
R6759 GND.n388 GND.n387 104.615
R6760 GND.n387 GND.n377 104.615
R6761 GND.n380 GND.n377 104.615
R6762 GND.n365 GND.n364 104.615
R6763 GND.n364 GND.n354 104.615
R6764 GND.n357 GND.n354 104.615
R6765 GND.n344 GND.n343 104.615
R6766 GND.n343 GND.n333 104.615
R6767 GND.n336 GND.n333 104.615
R6768 GND.n321 GND.n320 104.615
R6769 GND.n320 GND.n310 104.615
R6770 GND.n313 GND.n310 104.615
R6771 GND.n301 GND.n300 104.615
R6772 GND.n300 GND.n290 104.615
R6773 GND.n293 GND.n290 104.615
R6774 GND.n278 GND.n277 104.615
R6775 GND.n277 GND.n267 104.615
R6776 GND.n270 GND.n267 104.615
R6777 GND.n6785 GND.n654 99.6594
R6778 GND.n6783 GND.n6782 99.6594
R6779 GND.n6778 GND.n662 99.6594
R6780 GND.n6776 GND.n6775 99.6594
R6781 GND.n671 GND.n670 99.6594
R6782 GND.n6767 GND.n675 99.6594
R6783 GND.n6765 GND.n6764 99.6594
R6784 GND.n6760 GND.n681 99.6594
R6785 GND.n6758 GND.n6757 99.6594
R6786 GND.n6753 GND.n688 99.6594
R6787 GND.n6751 GND.n6750 99.6594
R6788 GND.n6744 GND.n696 99.6594
R6789 GND.n6742 GND.n6741 99.6594
R6790 GND.n6737 GND.n702 99.6594
R6791 GND.n6735 GND.n6734 99.6594
R6792 GND.n6730 GND.n709 99.6594
R6793 GND.n6728 GND.n6727 99.6594
R6794 GND.n6720 GND.n716 99.6594
R6795 GND.n6718 GND.n6717 99.6594
R6796 GND.n6713 GND.n723 99.6594
R6797 GND.n6711 GND.n6710 99.6594
R6798 GND.n6706 GND.n730 99.6594
R6799 GND.n6704 GND.n6703 99.6594
R6800 GND.n6696 GND.n737 99.6594
R6801 GND.n6694 GND.n6693 99.6594
R6802 GND.n6689 GND.n744 99.6594
R6803 GND.n6687 GND.n6686 99.6594
R6804 GND.n6682 GND.n751 99.6594
R6805 GND.n6680 GND.n6679 99.6594
R6806 GND.n756 GND.n755 99.6594
R6807 GND.n4630 GND.n4629 99.6594
R6808 GND.n4624 GND.n3888 99.6594
R6809 GND.n4621 GND.n3889 99.6594
R6810 GND.n4617 GND.n3890 99.6594
R6811 GND.n4613 GND.n3891 99.6594
R6812 GND.n4609 GND.n3892 99.6594
R6813 GND.n4606 GND.n3893 99.6594
R6814 GND.n4602 GND.n3894 99.6594
R6815 GND.n4598 GND.n3895 99.6594
R6816 GND.n4594 GND.n3896 99.6594
R6817 GND.n4590 GND.n3897 99.6594
R6818 GND.n4586 GND.n3898 99.6594
R6819 GND.n4583 GND.n3900 99.6594
R6820 GND.n3901 GND.n3882 99.6594
R6821 GND.n4633 GND.n4632 99.6594
R6822 GND.n4152 GND.n3902 99.6594
R6823 GND.n4159 GND.n3903 99.6594
R6824 GND.n4164 GND.n3904 99.6594
R6825 GND.n4172 GND.n3905 99.6594
R6826 GND.n4174 GND.n3906 99.6594
R6827 GND.n4182 GND.n3907 99.6594
R6828 GND.n4184 GND.n3908 99.6594
R6829 GND.n4192 GND.n3909 99.6594
R6830 GND.n4197 GND.n3910 99.6594
R6831 GND.n4205 GND.n3911 99.6594
R6832 GND.n4207 GND.n3912 99.6594
R6833 GND.n4215 GND.n3913 99.6594
R6834 GND.n4217 GND.n3914 99.6594
R6835 GND.n4225 GND.n3915 99.6594
R6836 GND.n4227 GND.n3916 99.6594
R6837 GND.n2033 GND.n1995 99.6594
R6838 GND.n2035 GND.n2034 99.6594
R6839 GND.n2036 GND.n2000 99.6594
R6840 GND.n2038 GND.n2037 99.6594
R6841 GND.n2039 GND.n2005 99.6594
R6842 GND.n2040 GND.n2010 99.6594
R6843 GND.n2042 GND.n2013 99.6594
R6844 GND.n2043 GND.n2015 99.6594
R6845 GND.n2045 GND.n2018 99.6594
R6846 GND.n2046 GND.n2020 99.6594
R6847 GND.n2048 GND.n2023 99.6594
R6848 GND.n2049 GND.n2027 99.6594
R6849 GND.n2051 GND.n2030 99.6594
R6850 GND.n5010 GND.n5009 99.6594
R6851 GND.n5007 GND.n5006 99.6594
R6852 GND.n4896 GND.n4895 99.6594
R6853 GND.n4899 GND.n4898 99.6594
R6854 GND.n4906 GND.n4905 99.6594
R6855 GND.n4911 GND.n4910 99.6594
R6856 GND.n4914 GND.n4913 99.6594
R6857 GND.n4919 GND.n4918 99.6594
R6858 GND.n4922 GND.n4921 99.6594
R6859 GND.n4930 GND.n4929 99.6594
R6860 GND.n4933 GND.n4932 99.6594
R6861 GND.n4938 GND.n4937 99.6594
R6862 GND.n4941 GND.n4940 99.6594
R6863 GND.n4946 GND.n4945 99.6594
R6864 GND.n4949 GND.n4948 99.6594
R6865 GND.n4956 GND.n4955 99.6594
R6866 GND.n4957 GND.n1985 99.6594
R6867 GND.n2340 GND.n1879 99.6594
R6868 GND.n2349 GND.n2348 99.6594
R6869 GND.n2352 GND.n2351 99.6594
R6870 GND.n2359 GND.n2358 99.6594
R6871 GND.n2362 GND.n2361 99.6594
R6872 GND.n2371 GND.n2370 99.6594
R6873 GND.n2374 GND.n2373 99.6594
R6874 GND.n2381 GND.n2380 99.6594
R6875 GND.n2384 GND.n2383 99.6594
R6876 GND.n2391 GND.n2390 99.6594
R6877 GND.n2394 GND.n2393 99.6594
R6878 GND.n2403 GND.n2402 99.6594
R6879 GND.n2406 GND.n2405 99.6594
R6880 GND.n2413 GND.n2412 99.6594
R6881 GND.n2416 GND.n2415 99.6594
R6882 GND.n2423 GND.n2422 99.6594
R6883 GND.n2426 GND.n2425 99.6594
R6884 GND.n2436 GND.n2435 99.6594
R6885 GND.n2439 GND.n2438 99.6594
R6886 GND.n2446 GND.n2445 99.6594
R6887 GND.n2449 GND.n2448 99.6594
R6888 GND.n2456 GND.n2455 99.6594
R6889 GND.n2459 GND.n2458 99.6594
R6890 GND.n2469 GND.n2468 99.6594
R6891 GND.n2472 GND.n2471 99.6594
R6892 GND.n2479 GND.n2478 99.6594
R6893 GND.n2482 GND.n2481 99.6594
R6894 GND.n2489 GND.n2488 99.6594
R6895 GND.n2492 GND.n2491 99.6594
R6896 GND.n2499 GND.n2498 99.6594
R6897 GND.n3775 GND.n3774 99.6594
R6898 GND.n3776 GND.n3766 99.6594
R6899 GND.n3785 GND.n3784 99.6594
R6900 GND.n3786 GND.n3762 99.6594
R6901 GND.n3796 GND.n3795 99.6594
R6902 GND.n3797 GND.n3756 99.6594
R6903 GND.n3807 GND.n3806 99.6594
R6904 GND.n3808 GND.n3313 99.6594
R6905 GND.n4851 GND.n4850 99.6594
R6906 GND.n4845 GND.n2957 99.6594
R6907 GND.n4842 GND.n2958 99.6594
R6908 GND.n4838 GND.n2959 99.6594
R6909 GND.n4834 GND.n2960 99.6594
R6910 GND.n4830 GND.n2961 99.6594
R6911 GND.n4825 GND.n2962 99.6594
R6912 GND.n762 GND.n761 99.6594
R6913 GND.n6668 GND.n6667 99.6594
R6914 GND.n6665 GND.n6664 99.6594
R6915 GND.n6660 GND.n773 99.6594
R6916 GND.n6658 GND.n6657 99.6594
R6917 GND.n778 GND.n777 99.6594
R6918 GND.n4266 GND.n3917 99.6594
R6919 GND.n4263 GND.n3918 99.6594
R6920 GND.n4259 GND.n3919 99.6594
R6921 GND.n4255 GND.n3920 99.6594
R6922 GND.n4251 GND.n3921 99.6594
R6923 GND.n4241 GND.n3922 99.6594
R6924 GND.n6401 GND.n6400 99.6594
R6925 GND.n5329 GND.n5328 99.6594
R6926 GND.n4264 GND.n3917 99.6594
R6927 GND.n4260 GND.n3918 99.6594
R6928 GND.n4256 GND.n3919 99.6594
R6929 GND.n4252 GND.n3920 99.6594
R6930 GND.n4240 GND.n3921 99.6594
R6931 GND.n4104 GND.n3922 99.6594
R6932 GND.n777 GND.n774 99.6594
R6933 GND.n6659 GND.n6658 99.6594
R6934 GND.n773 GND.n766 99.6594
R6935 GND.n6666 GND.n6665 99.6594
R6936 GND.n6669 GND.n6668 99.6594
R6937 GND.n761 GND.n643 99.6594
R6938 GND.n4851 GND.n2965 99.6594
R6939 GND.n4843 GND.n2957 99.6594
R6940 GND.n4839 GND.n2958 99.6594
R6941 GND.n4835 GND.n2959 99.6594
R6942 GND.n4831 GND.n2960 99.6594
R6943 GND.n4826 GND.n2961 99.6594
R6944 GND.n2983 GND.n2962 99.6594
R6945 GND.n3809 GND.n3808 99.6594
R6946 GND.n3806 GND.n3805 99.6594
R6947 GND.n3798 GND.n3797 99.6594
R6948 GND.n3795 GND.n3794 99.6594
R6949 GND.n3787 GND.n3786 99.6594
R6950 GND.n3784 GND.n3783 99.6594
R6951 GND.n3777 GND.n3776 99.6594
R6952 GND.n3774 GND.n3773 99.6594
R6953 GND.n2341 GND.n2340 99.6594
R6954 GND.n2350 GND.n2349 99.6594
R6955 GND.n2351 GND.n2336 99.6594
R6956 GND.n2360 GND.n2359 99.6594
R6957 GND.n2361 GND.n2332 99.6594
R6958 GND.n2372 GND.n2371 99.6594
R6959 GND.n2373 GND.n2328 99.6594
R6960 GND.n2382 GND.n2381 99.6594
R6961 GND.n2383 GND.n2324 99.6594
R6962 GND.n2392 GND.n2391 99.6594
R6963 GND.n2393 GND.n2320 99.6594
R6964 GND.n2404 GND.n2403 99.6594
R6965 GND.n2405 GND.n2316 99.6594
R6966 GND.n2414 GND.n2413 99.6594
R6967 GND.n2415 GND.n2312 99.6594
R6968 GND.n2424 GND.n2423 99.6594
R6969 GND.n2425 GND.n2308 99.6594
R6970 GND.n2437 GND.n2436 99.6594
R6971 GND.n2438 GND.n2304 99.6594
R6972 GND.n2447 GND.n2446 99.6594
R6973 GND.n2448 GND.n2300 99.6594
R6974 GND.n2457 GND.n2456 99.6594
R6975 GND.n2458 GND.n2296 99.6594
R6976 GND.n2470 GND.n2469 99.6594
R6977 GND.n2471 GND.n2292 99.6594
R6978 GND.n2480 GND.n2479 99.6594
R6979 GND.n2481 GND.n2288 99.6594
R6980 GND.n2490 GND.n2489 99.6594
R6981 GND.n2491 GND.n2284 99.6594
R6982 GND.n2500 GND.n2499 99.6594
R6983 GND.n4958 GND.n4957 99.6594
R6984 GND.n4955 GND.n4950 99.6594
R6985 GND.n4948 GND.n4947 99.6594
R6986 GND.n4945 GND.n4942 99.6594
R6987 GND.n4940 GND.n4939 99.6594
R6988 GND.n4937 GND.n4934 99.6594
R6989 GND.n4932 GND.n4931 99.6594
R6990 GND.n4929 GND.n4923 99.6594
R6991 GND.n4921 GND.n4920 99.6594
R6992 GND.n4918 GND.n4915 99.6594
R6993 GND.n4913 GND.n4912 99.6594
R6994 GND.n4910 GND.n4907 99.6594
R6995 GND.n4905 GND.n4904 99.6594
R6996 GND.n4898 GND.n4897 99.6594
R6997 GND.n4895 GND.n4890 99.6594
R6998 GND.n5008 GND.n5007 99.6594
R6999 GND.n5012 GND.n5011 99.6594
R7000 GND.n2051 GND.n2050 99.6594
R7001 GND.n2049 GND.n2026 99.6594
R7002 GND.n2048 GND.n2047 99.6594
R7003 GND.n2046 GND.n2019 99.6594
R7004 GND.n2045 GND.n2044 99.6594
R7005 GND.n2043 GND.n2014 99.6594
R7006 GND.n2042 GND.n2041 99.6594
R7007 GND.n2040 GND.n2009 99.6594
R7008 GND.n2039 GND.n2004 99.6594
R7009 GND.n2038 GND.n2001 99.6594
R7010 GND.n2036 GND.n1999 99.6594
R7011 GND.n2035 GND.n1996 99.6594
R7012 GND.n2033 GND.n1991 99.6594
R7013 GND.n4630 GND.n3925 99.6594
R7014 GND.n4622 GND.n3888 99.6594
R7015 GND.n4618 GND.n3889 99.6594
R7016 GND.n4614 GND.n3890 99.6594
R7017 GND.n4559 GND.n3891 99.6594
R7018 GND.n4607 GND.n3892 99.6594
R7019 GND.n4603 GND.n3893 99.6594
R7020 GND.n4599 GND.n3894 99.6594
R7021 GND.n4595 GND.n3895 99.6594
R7022 GND.n4591 GND.n3896 99.6594
R7023 GND.n4574 GND.n3897 99.6594
R7024 GND.n4584 GND.n3898 99.6594
R7025 GND.n3900 GND.n3899 99.6594
R7026 GND.n3901 GND.n3881 99.6594
R7027 GND.n4632 GND.n3886 99.6594
R7028 GND.n4158 GND.n3902 99.6594
R7029 GND.n4165 GND.n3903 99.6594
R7030 GND.n4171 GND.n3904 99.6594
R7031 GND.n4175 GND.n3905 99.6594
R7032 GND.n4181 GND.n3906 99.6594
R7033 GND.n4185 GND.n3907 99.6594
R7034 GND.n4191 GND.n3908 99.6594
R7035 GND.n4198 GND.n3909 99.6594
R7036 GND.n4204 GND.n3910 99.6594
R7037 GND.n4208 GND.n3911 99.6594
R7038 GND.n4214 GND.n3912 99.6594
R7039 GND.n4218 GND.n3913 99.6594
R7040 GND.n4224 GND.n3914 99.6594
R7041 GND.n4228 GND.n3915 99.6594
R7042 GND.n4272 GND.n3916 99.6594
R7043 GND.n755 GND.n752 99.6594
R7044 GND.n6681 GND.n6680 99.6594
R7045 GND.n751 GND.n745 99.6594
R7046 GND.n6688 GND.n6687 99.6594
R7047 GND.n744 GND.n738 99.6594
R7048 GND.n6695 GND.n6694 99.6594
R7049 GND.n737 GND.n731 99.6594
R7050 GND.n6705 GND.n6704 99.6594
R7051 GND.n730 GND.n724 99.6594
R7052 GND.n6712 GND.n6711 99.6594
R7053 GND.n723 GND.n717 99.6594
R7054 GND.n6719 GND.n6718 99.6594
R7055 GND.n716 GND.n710 99.6594
R7056 GND.n6729 GND.n6728 99.6594
R7057 GND.n709 GND.n703 99.6594
R7058 GND.n6736 GND.n6735 99.6594
R7059 GND.n702 GND.n697 99.6594
R7060 GND.n6743 GND.n6742 99.6594
R7061 GND.n696 GND.n689 99.6594
R7062 GND.n6752 GND.n6751 99.6594
R7063 GND.n688 GND.n682 99.6594
R7064 GND.n6759 GND.n6758 99.6594
R7065 GND.n681 GND.n676 99.6594
R7066 GND.n6766 GND.n6765 99.6594
R7067 GND.n675 GND.n674 99.6594
R7068 GND.n670 GND.n663 99.6594
R7069 GND.n6777 GND.n6776 99.6594
R7070 GND.n662 GND.n656 99.6594
R7071 GND.n6784 GND.n6783 99.6594
R7072 GND.n654 GND.n651 99.6594
R7073 GND.n5329 GND.n1683 99.6594
R7074 GND.n6400 GND.n1006 99.6594
R7075 GND.n2512 GND.n2511 99.6594
R7076 GND.n2515 GND.n2514 99.6594
R7077 GND.n2522 GND.n2521 99.6594
R7078 GND.n2525 GND.n2524 99.6594
R7079 GND.n2532 GND.n2531 99.6594
R7080 GND.n2513 GND.n2512 99.6594
R7081 GND.n2514 GND.n2274 99.6594
R7082 GND.n2523 GND.n2522 99.6594
R7083 GND.n2524 GND.n2270 99.6594
R7084 GND.n2533 GND.n2532 99.6594
R7085 GND.n2846 GND.n2052 99.6594
R7086 GND.n2852 GND.n2053 99.6594
R7087 GND.n2854 GND.n2054 99.6594
R7088 GND.n2862 GND.n2055 99.6594
R7089 GND.n2864 GND.n2056 99.6594
R7090 GND.n2874 GND.n2057 99.6594
R7091 GND.n2876 GND.n2057 99.6594
R7092 GND.n2873 GND.n2056 99.6594
R7093 GND.n2865 GND.n2055 99.6594
R7094 GND.n2861 GND.n2054 99.6594
R7095 GND.n2855 GND.n2053 99.6594
R7096 GND.n2851 GND.n2052 99.6594
R7097 GND.n3408 GND.n3407 95.6126
R7098 GND.n3400 GND.n3399 95.6126
R7099 GND.n3300 GND.n3299 95.6126
R7100 GND.n3291 GND.n3290 95.6126
R7101 GND.n3400 GND.t136 88.518
R7102 GND.n3300 GND.t172 88.518
R7103 GND.n3408 GND.t155 88.5177
R7104 GND.n3291 GND.t190 88.5177
R7105 GND.n2980 GND.t196 85.8607
R7106 GND.n3758 GND.t101 85.8607
R7107 GND.n3431 GND.n3430 77.8372
R7108 GND.n5418 GND.n1595 73.2972
R7109 GND.n5412 GND.n1595 73.2972
R7110 GND.n5412 GND.n5411 73.2972
R7111 GND.n5411 GND.n5410 73.2972
R7112 GND.n5410 GND.n1602 73.2972
R7113 GND.n5404 GND.n1602 73.2972
R7114 GND.n5404 GND.n5403 73.2972
R7115 GND.n5403 GND.n5402 73.2972
R7116 GND.n5402 GND.n1610 73.2972
R7117 GND.n5396 GND.n1610 73.2972
R7118 GND.n5396 GND.n5395 73.2972
R7119 GND.n5395 GND.n5394 73.2972
R7120 GND.n5394 GND.n1618 73.2972
R7121 GND.n5388 GND.n1618 73.2972
R7122 GND.n5388 GND.n5387 73.2972
R7123 GND.n5387 GND.n5386 73.2972
R7124 GND.n5386 GND.n1626 73.2972
R7125 GND.n5380 GND.n1626 73.2972
R7126 GND.n5380 GND.n5379 73.2972
R7127 GND.n5379 GND.n5378 73.2972
R7128 GND.n5378 GND.n1634 73.2972
R7129 GND.n5372 GND.n1634 73.2972
R7130 GND.n5372 GND.n5371 73.2972
R7131 GND.n5371 GND.n5370 73.2972
R7132 GND.n5370 GND.n1642 73.2972
R7133 GND.n5364 GND.n1642 73.2972
R7134 GND.n5364 GND.n5363 73.2972
R7135 GND.n5363 GND.n5362 73.2972
R7136 GND.n5362 GND.n1650 73.2972
R7137 GND.n5356 GND.n1650 73.2972
R7138 GND.n5356 GND.n5355 73.2972
R7139 GND.n5355 GND.n5354 73.2972
R7140 GND.n5354 GND.n1658 73.2972
R7141 GND.n5348 GND.n1658 73.2972
R7142 GND.n5348 GND.n5347 73.2972
R7143 GND.n5347 GND.n5346 73.2972
R7144 GND.n5346 GND.n1666 73.2972
R7145 GND.n5340 GND.n1666 73.2972
R7146 GND.n5340 GND.n5339 73.2972
R7147 GND.n5339 GND.n5338 73.2972
R7148 GND.n5338 GND.n1674 73.2972
R7149 GND.n5332 GND.n1674 73.2972
R7150 GND.n5332 GND.n5331 73.2972
R7151 GND.n3432 GND.n3422 72.8411
R7152 GND.n3438 GND.n3420 72.8411
R7153 GND.n3439 GND.n3419 72.8411
R7154 GND.n3445 GND.n3417 72.8411
R7155 GND.n3276 GND.n3275 72.8411
R7156 GND.n3262 GND.n3261 72.8411
R7157 GND.n3260 GND.n3251 72.8411
R7158 GND.n4664 GND.n3281 71.676
R7159 GND.n4662 GND.n4661 71.676
R7160 GND.n4657 GND.n3285 71.676
R7161 GND.n4655 GND.n4654 71.676
R7162 GND.n4650 GND.n3288 71.676
R7163 GND.n4648 GND.n4647 71.676
R7164 GND.n4642 GND.n3293 71.676
R7165 GND.n4640 GND.n4639 71.676
R7166 GND.n3878 GND.n3877 71.676
R7167 GND.n3875 GND.n3874 71.676
R7168 GND.n3869 GND.n3302 71.676
R7169 GND.n3867 GND.n3866 71.676
R7170 GND.n3862 GND.n3305 71.676
R7171 GND.n3860 GND.n3859 71.676
R7172 GND.n3855 GND.n3308 71.676
R7173 GND.n3853 GND.n3852 71.676
R7174 GND.n3848 GND.n3847 71.676
R7175 GND.n3452 GND.n3451 71.676
R7176 GND.n3458 GND.n3457 71.676
R7177 GND.n3461 GND.n3460 71.676
R7178 GND.n3466 GND.n3465 71.676
R7179 GND.n3469 GND.n3468 71.676
R7180 GND.n3474 GND.n3473 71.676
R7181 GND.n3477 GND.n3476 71.676
R7182 GND.n3482 GND.n3481 71.676
R7183 GND.n3485 GND.n3484 71.676
R7184 GND.n3488 GND.n3487 71.676
R7185 GND.n3493 GND.n3492 71.676
R7186 GND.n3496 GND.n3495 71.676
R7187 GND.n3501 GND.n3500 71.676
R7188 GND.n3504 GND.n3503 71.676
R7189 GND.n3509 GND.n3508 71.676
R7190 GND.n3512 GND.n3511 71.676
R7191 GND.n3517 GND.n3516 71.676
R7192 GND.n3453 GND.n3452 71.676
R7193 GND.n3459 GND.n3458 71.676
R7194 GND.n3460 GND.n3413 71.676
R7195 GND.n3467 GND.n3466 71.676
R7196 GND.n3468 GND.n3411 71.676
R7197 GND.n3475 GND.n3474 71.676
R7198 GND.n3476 GND.n3406 71.676
R7199 GND.n3483 GND.n3482 71.676
R7200 GND.n3486 GND.n3485 71.676
R7201 GND.n3487 GND.n3403 71.676
R7202 GND.n3494 GND.n3493 71.676
R7203 GND.n3495 GND.n3398 71.676
R7204 GND.n3502 GND.n3501 71.676
R7205 GND.n3503 GND.n3396 71.676
R7206 GND.n3510 GND.n3509 71.676
R7207 GND.n3511 GND.n3394 71.676
R7208 GND.n3518 GND.n3517 71.676
R7209 GND.n3847 GND.n3309 71.676
R7210 GND.n3854 GND.n3853 71.676
R7211 GND.n3308 GND.n3306 71.676
R7212 GND.n3861 GND.n3860 71.676
R7213 GND.n3305 GND.n3303 71.676
R7214 GND.n3868 GND.n3867 71.676
R7215 GND.n3302 GND.n3298 71.676
R7216 GND.n3876 GND.n3875 71.676
R7217 GND.n3296 GND.n3294 71.676
R7218 GND.n4641 GND.n4640 71.676
R7219 GND.n3293 GND.n3289 71.676
R7220 GND.n4649 GND.n4648 71.676
R7221 GND.n3288 GND.n3286 71.676
R7222 GND.n4656 GND.n4655 71.676
R7223 GND.n3285 GND.n3283 71.676
R7224 GND.n4663 GND.n4662 71.676
R7225 GND.n3281 GND.n3246 71.676
R7226 GND.n2980 GND.n2979 65.552
R7227 GND.n3758 GND.n3757 65.552
R7228 GND.n3449 GND.n3448 61.3137
R7229 GND.n5330 GND.n1682 59.7182
R7230 GND.n6399 GND.n1000 59.7182
R7231 GND.n3409 GND.n3408 59.5399
R7232 GND.n3401 GND.n3400 59.5399
R7233 GND.n3871 GND.n3300 59.5399
R7234 GND.n4644 GND.n3291 59.5399
R7235 GND.n239 GND.n238 56.3974
R7236 GND.n241 GND.n240 56.3974
R7237 GND.n195 GND.n194 56.3974
R7238 GND.n197 GND.n196 56.3974
R7239 GND.n151 GND.n150 56.3974
R7240 GND.n153 GND.n152 56.3974
R7241 GND.n107 GND.n106 56.3974
R7242 GND.n109 GND.n108 56.3974
R7243 GND.n63 GND.n62 56.3974
R7244 GND.n65 GND.n64 56.3974
R7245 GND.n20 GND.n19 56.3974
R7246 GND.n22 GND.n21 56.3974
R7247 GND.n505 GND.n504 56.3974
R7248 GND.n503 GND.n502 56.3974
R7249 GND.n461 GND.n460 56.3974
R7250 GND.n459 GND.n458 56.3974
R7251 GND.n417 GND.n416 56.3974
R7252 GND.n415 GND.n414 56.3974
R7253 GND.n373 GND.n372 56.3974
R7254 GND.n371 GND.n370 56.3974
R7255 GND.n329 GND.n328 56.3974
R7256 GND.n327 GND.n326 56.3974
R7257 GND.n286 GND.n285 56.3974
R7258 GND.n284 GND.n283 56.3974
R7259 GND.n3429 GND.n3428 54.358
R7260 GND.n3273 GND.n3272 54.358
R7261 GND.n3255 GND.n3254 52.8267
R7262 GND.n225 GND.t17 52.3082
R7263 GND.n248 GND.t53 52.3082
R7264 GND.n181 GND.t52 52.3082
R7265 GND.n204 GND.t87 52.3082
R7266 GND.n137 GND.t19 52.3082
R7267 GND.n160 GND.t64 52.3082
R7268 GND.n93 GND.t47 52.3082
R7269 GND.n116 GND.t55 52.3082
R7270 GND.n49 GND.t71 52.3082
R7271 GND.n72 GND.t42 52.3082
R7272 GND.n6 GND.t33 52.3082
R7273 GND.n29 GND.t82 52.3082
R7274 GND.n512 GND.t26 52.3082
R7275 GND.n489 GND.t65 52.3082
R7276 GND.n468 GND.t56 52.3082
R7277 GND.n445 GND.t5 52.3082
R7278 GND.n424 GND.t28 52.3082
R7279 GND.n401 GND.t66 52.3082
R7280 GND.n380 GND.t58 52.3082
R7281 GND.n357 GND.t63 52.3082
R7282 GND.n336 GND.t50 52.3082
R7283 GND.n313 GND.t18 52.3082
R7284 GND.n293 GND.t7 52.3082
R7285 GND.n270 GND.t69 52.3082
R7286 GND.n2872 GND.n2871 49.2611
R7287 GND.n2007 GND.n2006 49.2611
R7288 GND.n2025 GND.n2024 49.2611
R7289 GND.n4901 GND.n4900 49.2611
R7290 GND.n4927 GND.n4926 49.2611
R7291 GND.n4954 GND.n4953 49.2611
R7292 GND.n4562 GND.n4561 49.2611
R7293 GND.n4577 GND.n4576 49.2611
R7294 GND.n4162 GND.n4161 49.2611
R7295 GND.n4195 GND.n4194 49.2611
R7296 GND.n4137 GND.n4136 49.2611
R7297 GND.n759 GND.n758 49.2611
R7298 GND.n6700 GND.n6699 49.2611
R7299 GND.n6724 GND.n6723 49.2611
R7300 GND.n692 GND.n691 49.2611
R7301 GND.n669 GND.n668 49.2611
R7302 GND.n781 GND.n780 49.2611
R7303 GND.n4243 GND.n4242 49.2611
R7304 GND.n2368 GND.n2367 49.2611
R7305 GND.n2400 GND.n2399 49.2611
R7306 GND.n2432 GND.n2431 49.2611
R7307 GND.n2465 GND.n2464 49.2611
R7308 GND.n2282 GND.n2281 49.2611
R7309 GND.n2268 GND.n2267 49.2611
R7310 GND.n3439 GND.n3438 48.2005
R7311 GND.n3262 GND.n3251 48.2005
R7312 GND.n4667 GND.n3279 44.3322
R7313 GND.n3445 GND.n3444 43.0884
R7314 GND.n3433 GND.n3432 43.0884
R7315 GND.n3256 GND.n3253 43.0884
R7316 GND.n3276 GND.n3249 43.0884
R7317 GND.n2875 GND.n2872 42.2793
R7318 GND.n5037 GND.n2007 42.2793
R7319 GND.n5019 GND.n2025 42.2793
R7320 GND.n4902 GND.n4901 42.2793
R7321 GND.n4928 GND.n4927 42.2793
R7322 GND.n4960 GND.n4954 42.2793
R7323 GND.n4828 GND.n2980 42.2793
R7324 GND.n3759 GND.n3758 42.2793
R7325 GND.n4611 GND.n4562 42.2793
R7326 GND.n4588 GND.n4577 42.2793
R7327 GND.n4163 GND.n4162 42.2793
R7328 GND.n4196 GND.n4195 42.2793
R7329 GND.n4138 GND.n4137 42.2793
R7330 GND.n6677 GND.n759 42.2793
R7331 GND.n6701 GND.n6700 42.2793
R7332 GND.n6725 GND.n6724 42.2793
R7333 GND.n6749 GND.n692 42.2793
R7334 GND.n6772 GND.n669 42.2793
R7335 GND.n6655 GND.n781 42.2793
R7336 GND.n4244 GND.n4243 42.2793
R7337 GND.n2369 GND.n2368 42.2793
R7338 GND.n2401 GND.n2400 42.2793
R7339 GND.n2433 GND.n2432 42.2793
R7340 GND.n2466 GND.n2465 42.2793
R7341 GND.n2283 GND.n2282 42.2793
R7342 GND.n2269 GND.n2268 42.2793
R7343 GND.n3430 GND.n3429 41.6274
R7344 GND.n3274 GND.n3273 41.6274
R7345 GND.n3432 GND.n3431 39.875
R7346 GND.n3849 GND.n3846 34.8103
R7347 GND.n3521 GND.n3392 34.8103
R7348 GND.n5320 GND.n1682 34.1249
R7349 GND.n5320 GND.n5319 34.1249
R7350 GND.n5319 GND.n5318 34.1249
R7351 GND.n5318 GND.n1689 34.1249
R7352 GND.n5312 GND.n1689 34.1249
R7353 GND.n5312 GND.n5311 34.1249
R7354 GND.n5311 GND.n5310 34.1249
R7355 GND.n5310 GND.n1698 34.1249
R7356 GND.n5304 GND.n1698 34.1249
R7357 GND.n5304 GND.n5303 34.1249
R7358 GND.n5303 GND.n5302 34.1249
R7359 GND.n5302 GND.n1706 34.1249
R7360 GND.n5296 GND.n1706 34.1249
R7361 GND.n5296 GND.n5295 34.1249
R7362 GND.n5295 GND.n5294 34.1249
R7363 GND.n5294 GND.n1714 34.1249
R7364 GND.n5288 GND.n1714 34.1249
R7365 GND.n5288 GND.n5287 34.1249
R7366 GND.n5287 GND.n5286 34.1249
R7367 GND.n5286 GND.n1722 34.1249
R7368 GND.n5280 GND.n1722 34.1249
R7369 GND.n5280 GND.n5279 34.1249
R7370 GND.n5279 GND.n5278 34.1249
R7371 GND.n5278 GND.n1730 34.1249
R7372 GND.n5272 GND.n1730 34.1249
R7373 GND.n5272 GND.n5271 34.1249
R7374 GND.n5271 GND.n5270 34.1249
R7375 GND.n5270 GND.n1738 34.1249
R7376 GND.n5264 GND.n1738 34.1249
R7377 GND.n5264 GND.n5263 34.1249
R7378 GND.n5263 GND.n5262 34.1249
R7379 GND.n5262 GND.n1746 34.1249
R7380 GND.n5256 GND.n1746 34.1249
R7381 GND.n5256 GND.n5255 34.1249
R7382 GND.n5255 GND.n5254 34.1249
R7383 GND.n5254 GND.n1754 34.1249
R7384 GND.n5248 GND.n1754 34.1249
R7385 GND.n5248 GND.n5247 34.1249
R7386 GND.n5247 GND.n5246 34.1249
R7387 GND.n5246 GND.n1762 34.1249
R7388 GND.n5240 GND.n1762 34.1249
R7389 GND.n5240 GND.n5239 34.1249
R7390 GND.n5239 GND.n5238 34.1249
R7391 GND.n5238 GND.n1770 34.1249
R7392 GND.n5232 GND.n1770 34.1249
R7393 GND.n5232 GND.n5231 34.1249
R7394 GND.n5231 GND.n5230 34.1249
R7395 GND.n5230 GND.n1778 34.1249
R7396 GND.n5224 GND.n1778 34.1249
R7397 GND.n5224 GND.n5223 34.1249
R7398 GND.n5223 GND.n5222 34.1249
R7399 GND.n5222 GND.n1786 34.1249
R7400 GND.n5216 GND.n1786 34.1249
R7401 GND.n5216 GND.n5215 34.1249
R7402 GND.n5215 GND.n5214 34.1249
R7403 GND.n5214 GND.n1794 34.1249
R7404 GND.n5208 GND.n1794 34.1249
R7405 GND.n5208 GND.n5207 34.1249
R7406 GND.n5207 GND.n5206 34.1249
R7407 GND.n5206 GND.n1802 34.1249
R7408 GND.n5200 GND.n1802 34.1249
R7409 GND.n5200 GND.n5199 34.1249
R7410 GND.n5199 GND.n5198 34.1249
R7411 GND.n5198 GND.n1810 34.1249
R7412 GND.n5192 GND.n1810 34.1249
R7413 GND.n5192 GND.n5191 34.1249
R7414 GND.n5191 GND.n5190 34.1249
R7415 GND.n5190 GND.n1818 34.1249
R7416 GND.n5184 GND.n1818 34.1249
R7417 GND.n5184 GND.n5183 34.1249
R7418 GND.n5183 GND.n5182 34.1249
R7419 GND.n5182 GND.n1826 34.1249
R7420 GND.n5176 GND.n1826 34.1249
R7421 GND.n5176 GND.n5175 34.1249
R7422 GND.n5175 GND.n5174 34.1249
R7423 GND.n5174 GND.n1834 34.1249
R7424 GND.n5168 GND.n1834 34.1249
R7425 GND.n5168 GND.n5167 34.1249
R7426 GND.n5167 GND.n5166 34.1249
R7427 GND.n5166 GND.n1842 34.1249
R7428 GND.n5160 GND.n1842 34.1249
R7429 GND.n5160 GND.n5159 34.1249
R7430 GND.n5159 GND.n5158 34.1249
R7431 GND.n5158 GND.n1850 34.1249
R7432 GND.n5152 GND.n1850 34.1249
R7433 GND.n5152 GND.n5151 34.1249
R7434 GND.n5151 GND.n5150 34.1249
R7435 GND.n5150 GND.n1858 34.1249
R7436 GND.n5144 GND.n1858 34.1249
R7437 GND.n5144 GND.n5143 34.1249
R7438 GND.n5143 GND.n5142 34.1249
R7439 GND.n5142 GND.n1866 34.1249
R7440 GND.n5136 GND.n5135 34.1249
R7441 GND.n2032 GND.n1988 34.1249
R7442 GND.n4887 GND.n2058 34.1249
R7443 GND.n4881 GND.n2058 34.1249
R7444 GND.n4881 GND.n4880 34.1249
R7445 GND.n4880 GND.n4879 34.1249
R7446 GND.n4122 GND.n4121 34.1249
R7447 GND.n4123 GND.n4122 34.1249
R7448 GND.n4123 GND.n3887 34.1249
R7449 GND.n4135 GND.n3923 34.1249
R7450 GND.n6591 GND.n647 34.1249
R7451 GND.n6586 GND.n823 34.1249
R7452 GND.n6586 GND.n6585 34.1249
R7453 GND.n6585 GND.n6584 34.1249
R7454 GND.n6584 GND.n824 34.1249
R7455 GND.n6578 GND.n824 34.1249
R7456 GND.n6578 GND.n6577 34.1249
R7457 GND.n6577 GND.n6576 34.1249
R7458 GND.n6576 GND.n832 34.1249
R7459 GND.n6570 GND.n832 34.1249
R7460 GND.n6570 GND.n6569 34.1249
R7461 GND.n6569 GND.n6568 34.1249
R7462 GND.n6568 GND.n840 34.1249
R7463 GND.n6562 GND.n840 34.1249
R7464 GND.n6562 GND.n6561 34.1249
R7465 GND.n6561 GND.n6560 34.1249
R7466 GND.n6560 GND.n848 34.1249
R7467 GND.n6554 GND.n848 34.1249
R7468 GND.n6554 GND.n6553 34.1249
R7469 GND.n6553 GND.n6552 34.1249
R7470 GND.n6552 GND.n856 34.1249
R7471 GND.n6546 GND.n856 34.1249
R7472 GND.n6546 GND.n6545 34.1249
R7473 GND.n6545 GND.n6544 34.1249
R7474 GND.n6544 GND.n864 34.1249
R7475 GND.n6538 GND.n864 34.1249
R7476 GND.n6538 GND.n6537 34.1249
R7477 GND.n6537 GND.n6536 34.1249
R7478 GND.n6536 GND.n872 34.1249
R7479 GND.n6530 GND.n872 34.1249
R7480 GND.n6530 GND.n6529 34.1249
R7481 GND.n6529 GND.n6528 34.1249
R7482 GND.n6528 GND.n880 34.1249
R7483 GND.n6522 GND.n880 34.1249
R7484 GND.n6522 GND.n6521 34.1249
R7485 GND.n6521 GND.n6520 34.1249
R7486 GND.n6520 GND.n888 34.1249
R7487 GND.n6514 GND.n888 34.1249
R7488 GND.n6514 GND.n6513 34.1249
R7489 GND.n6513 GND.n6512 34.1249
R7490 GND.n6512 GND.n896 34.1249
R7491 GND.n6506 GND.n896 34.1249
R7492 GND.n6506 GND.n6505 34.1249
R7493 GND.n6505 GND.n6504 34.1249
R7494 GND.n6504 GND.n904 34.1249
R7495 GND.n6498 GND.n904 34.1249
R7496 GND.n6498 GND.n6497 34.1249
R7497 GND.n6497 GND.n6496 34.1249
R7498 GND.n6496 GND.n912 34.1249
R7499 GND.n6490 GND.n912 34.1249
R7500 GND.n6490 GND.n6489 34.1249
R7501 GND.n6489 GND.n6488 34.1249
R7502 GND.n6488 GND.n920 34.1249
R7503 GND.n6482 GND.n920 34.1249
R7504 GND.n6482 GND.n6481 34.1249
R7505 GND.n6481 GND.n6480 34.1249
R7506 GND.n6480 GND.n928 34.1249
R7507 GND.n6474 GND.n928 34.1249
R7508 GND.n6474 GND.n6473 34.1249
R7509 GND.n6473 GND.n6472 34.1249
R7510 GND.n6472 GND.n936 34.1249
R7511 GND.n6466 GND.n936 34.1249
R7512 GND.n6466 GND.n6465 34.1249
R7513 GND.n6465 GND.n6464 34.1249
R7514 GND.n6464 GND.n944 34.1249
R7515 GND.n6458 GND.n944 34.1249
R7516 GND.n6458 GND.n6457 34.1249
R7517 GND.n6457 GND.n6456 34.1249
R7518 GND.n6456 GND.n952 34.1249
R7519 GND.n6450 GND.n952 34.1249
R7520 GND.n6450 GND.n6449 34.1249
R7521 GND.n6449 GND.n6448 34.1249
R7522 GND.n6448 GND.n960 34.1249
R7523 GND.n6442 GND.n960 34.1249
R7524 GND.n6442 GND.n6441 34.1249
R7525 GND.n6441 GND.n6440 34.1249
R7526 GND.n6440 GND.n968 34.1249
R7527 GND.n6434 GND.n968 34.1249
R7528 GND.n6434 GND.n6433 34.1249
R7529 GND.n6433 GND.n6432 34.1249
R7530 GND.n6432 GND.n976 34.1249
R7531 GND.n6426 GND.n976 34.1249
R7532 GND.n6426 GND.n6425 34.1249
R7533 GND.n6425 GND.n6424 34.1249
R7534 GND.n6424 GND.n984 34.1249
R7535 GND.n6418 GND.n984 34.1249
R7536 GND.n6418 GND.n6417 34.1249
R7537 GND.n6417 GND.n6416 34.1249
R7538 GND.n6416 GND.n992 34.1249
R7539 GND.n6410 GND.n992 34.1249
R7540 GND.n6410 GND.n6409 34.1249
R7541 GND.n6409 GND.n6408 34.1249
R7542 GND.n6408 GND.n1000 34.1249
R7543 GND.n239 GND.n237 33.9871
R7544 GND.n195 GND.n193 33.9871
R7545 GND.n151 GND.n149 33.9871
R7546 GND.n107 GND.n105 33.9871
R7547 GND.n63 GND.n61 33.9871
R7548 GND.n20 GND.n18 33.9871
R7549 GND.n503 GND.n501 33.9871
R7550 GND.n459 GND.n457 33.9871
R7551 GND.n415 GND.n413 33.9871
R7552 GND.n371 GND.n369 33.9871
R7553 GND.n327 GND.n325 33.9871
R7554 GND.n284 GND.n282 33.9871
R7555 GND.n2929 GND.n2921 33.1012
R7556 GND.n3282 GND.n3244 33.1012
R7557 GND.n3446 GND.n3445 32.8641
R7558 GND.n3277 GND.n3276 32.8641
R7559 GND.n261 GND.n260 31.7975
R7560 GND.n217 GND.n216 31.7975
R7561 GND.n173 GND.n172 31.7975
R7562 GND.n129 GND.n128 31.7975
R7563 GND.n85 GND.n84 31.7975
R7564 GND.n42 GND.n41 31.7975
R7565 GND.n525 GND.n524 31.7975
R7566 GND.n481 GND.n480 31.7975
R7567 GND.n437 GND.n436 31.7975
R7568 GND.n393 GND.n392 31.7975
R7569 GND.n349 GND.n348 31.7975
R7570 GND.n306 GND.n305 31.7975
R7571 GND.n3404 GND.n2031 30.6565
R7572 GND.n4636 GND.n4635 30.6565
R7573 GND.n1874 GND.n1866 30.03
R7574 GND.n4121 GND.t119 30.03
R7575 GND.n823 GND.n655 30.03
R7576 GND.n3440 GND.n3439 27.0217
R7577 GND.n3438 GND.n3437 27.0217
R7578 GND.n3258 GND.n3251 27.0217
R7579 GND.n3263 GND.n3262 27.0217
R7580 GND.n4888 GND.n4887 25.935
R7581 GND.n4631 GND.n3887 25.935
R7582 GND.n3420 GND.n3419 25.8289
R7583 GND.n3261 GND.n3260 25.8289
R7584 GND.n4859 GND.n2949 23.2051
R7585 GND.n4678 GND.n3232 23.2051
R7586 GND.n3842 GND.n3242 23.2051
R7587 GND.n4873 GND.n2930 22.5226
R7588 GND.n4872 GND.t106 22.5226
R7589 GND.n3440 GND.n3418 21.1793
R7590 GND.n3437 GND.n3421 21.1793
R7591 GND.n3258 GND.n3257 21.1793
R7592 GND.n3264 GND.n3263 21.1793
R7593 GND.n4866 GND.n4865 21.1576
R7594 GND.n4677 GND.n3234 21.1576
R7595 GND.n3449 GND.n2934 20.4493
R7596 GND.n4668 GND.n4667 20.4493
R7597 GND.n3427 GND.t206 19.8005
R7598 GND.n3427 GND.t117 19.8005
R7599 GND.n3425 GND.t168 19.8005
R7600 GND.n3425 GND.t224 19.8005
R7601 GND.n3424 GND.t187 19.8005
R7602 GND.n3424 GND.t107 19.8005
R7603 GND.n3423 GND.t178 19.8005
R7604 GND.n3423 GND.t97 19.8005
R7605 GND.n3271 GND.t165 19.8005
R7606 GND.n3271 GND.t104 19.8005
R7607 GND.n3269 GND.t153 19.8005
R7608 GND.n3269 GND.t227 19.8005
R7609 GND.n3268 GND.t181 19.8005
R7610 GND.n3268 GND.t94 19.8005
R7611 GND.n3267 GND.t184 19.8005
R7612 GND.n3267 GND.t120 19.8005
R7613 GND.t223 GND.n2947 19.7927
R7614 GND.n4685 GND.n4684 19.7927
R7615 GND.n3417 GND.n3416 19.5087
R7616 GND.n3443 GND.n3417 19.5087
R7617 GND.n3441 GND.n3419 19.5087
R7618 GND.n3436 GND.n3420 19.5087
R7619 GND.n3434 GND.n3422 19.5087
R7620 GND.n3260 GND.n3259 19.5087
R7621 GND.n3261 GND.n3250 19.5087
R7622 GND.n3275 GND.n3266 19.5087
R7623 GND.n2850 GND.n2847 19.3944
R7624 GND.n2853 GND.n2850 19.3944
R7625 GND.n2856 GND.n2853 19.3944
R7626 GND.n2856 GND.n2844 19.3944
R7627 GND.n2860 GND.n2844 19.3944
R7628 GND.n2863 GND.n2860 19.3944
R7629 GND.n2866 GND.n2863 19.3944
R7630 GND.n2866 GND.n2842 19.3944
R7631 GND.n2870 GND.n2842 19.3944
R7632 GND.n2504 GND.n1892 19.3944
R7633 GND.n5126 GND.n1892 19.3944
R7634 GND.n5126 GND.n1893 19.3944
R7635 GND.n1900 GND.n1893 19.3944
R7636 GND.n1901 GND.n1900 19.3944
R7637 GND.n1902 GND.n1901 19.3944
R7638 GND.n2244 GND.n1902 19.3944
R7639 GND.n2244 GND.n1908 19.3944
R7640 GND.n1909 GND.n1908 19.3944
R7641 GND.n1910 GND.n1909 19.3944
R7642 GND.n2232 GND.n1910 19.3944
R7643 GND.n2232 GND.n1916 19.3944
R7644 GND.n1917 GND.n1916 19.3944
R7645 GND.n1918 GND.n1917 19.3944
R7646 GND.n2212 GND.n1918 19.3944
R7647 GND.n2212 GND.n1924 19.3944
R7648 GND.n1925 GND.n1924 19.3944
R7649 GND.n1926 GND.n1925 19.3944
R7650 GND.n2153 GND.n1926 19.3944
R7651 GND.n2153 GND.n1932 19.3944
R7652 GND.n1933 GND.n1932 19.3944
R7653 GND.n1934 GND.n1933 19.3944
R7654 GND.n2168 GND.n1934 19.3944
R7655 GND.n2168 GND.n1940 19.3944
R7656 GND.n1941 GND.n1940 19.3944
R7657 GND.n1942 GND.n1941 19.3944
R7658 GND.n2181 GND.n1942 19.3944
R7659 GND.n2181 GND.n1948 19.3944
R7660 GND.n1949 GND.n1948 19.3944
R7661 GND.n1950 GND.n1949 19.3944
R7662 GND.n2127 GND.n1950 19.3944
R7663 GND.n2127 GND.n1956 19.3944
R7664 GND.n1957 GND.n1956 19.3944
R7665 GND.n1958 GND.n1957 19.3944
R7666 GND.n2106 GND.n1958 19.3944
R7667 GND.n2106 GND.n1964 19.3944
R7668 GND.n1965 GND.n1964 19.3944
R7669 GND.n1966 GND.n1965 19.3944
R7670 GND.n2082 GND.n1966 19.3944
R7671 GND.n2082 GND.n1972 19.3944
R7672 GND.n1973 GND.n1972 19.3944
R7673 GND.n1974 GND.n1973 19.3944
R7674 GND.n2069 GND.n1974 19.3944
R7675 GND.n2069 GND.n1980 19.3944
R7676 GND.n1981 GND.n1980 19.3944
R7677 GND.n1982 GND.n1981 19.3944
R7678 GND.n2505 GND.n1896 19.3944
R7679 GND.n5124 GND.n1896 19.3944
R7680 GND.n5124 GND.n5123 19.3944
R7681 GND.n5123 GND.n5122 19.3944
R7682 GND.n5122 GND.n1899 19.3944
R7683 GND.n5118 GND.n1899 19.3944
R7684 GND.n5118 GND.n5117 19.3944
R7685 GND.n5117 GND.n5116 19.3944
R7686 GND.n5116 GND.n1907 19.3944
R7687 GND.n5112 GND.n1907 19.3944
R7688 GND.n5112 GND.n5111 19.3944
R7689 GND.n5111 GND.n5110 19.3944
R7690 GND.n5110 GND.n1915 19.3944
R7691 GND.n5106 GND.n1915 19.3944
R7692 GND.n5106 GND.n5105 19.3944
R7693 GND.n5105 GND.n5104 19.3944
R7694 GND.n5104 GND.n1923 19.3944
R7695 GND.n5100 GND.n1923 19.3944
R7696 GND.n5100 GND.n5099 19.3944
R7697 GND.n5099 GND.n5098 19.3944
R7698 GND.n5098 GND.n1931 19.3944
R7699 GND.n5094 GND.n1931 19.3944
R7700 GND.n5094 GND.n5093 19.3944
R7701 GND.n5093 GND.n5092 19.3944
R7702 GND.n5092 GND.n1939 19.3944
R7703 GND.n5088 GND.n1939 19.3944
R7704 GND.n5088 GND.n5087 19.3944
R7705 GND.n5087 GND.n5086 19.3944
R7706 GND.n5086 GND.n1947 19.3944
R7707 GND.n5082 GND.n1947 19.3944
R7708 GND.n5082 GND.n5081 19.3944
R7709 GND.n5081 GND.n5080 19.3944
R7710 GND.n5080 GND.n1955 19.3944
R7711 GND.n5076 GND.n1955 19.3944
R7712 GND.n5076 GND.n5075 19.3944
R7713 GND.n5075 GND.n5074 19.3944
R7714 GND.n5074 GND.n1963 19.3944
R7715 GND.n5070 GND.n1963 19.3944
R7716 GND.n5070 GND.n5069 19.3944
R7717 GND.n5069 GND.n5068 19.3944
R7718 GND.n5068 GND.n1971 19.3944
R7719 GND.n5064 GND.n1971 19.3944
R7720 GND.n5064 GND.n5063 19.3944
R7721 GND.n5063 GND.n5062 19.3944
R7722 GND.n5062 GND.n1979 19.3944
R7723 GND.n5058 GND.n1979 19.3944
R7724 GND.n5051 GND.n5050 19.3944
R7725 GND.n5050 GND.n5049 19.3944
R7726 GND.n5049 GND.n1997 19.3944
R7727 GND.n5045 GND.n1997 19.3944
R7728 GND.n5045 GND.n5044 19.3944
R7729 GND.n5044 GND.n5043 19.3944
R7730 GND.n5043 GND.n2002 19.3944
R7731 GND.n5039 GND.n2002 19.3944
R7732 GND.n5039 GND.n5038 19.3944
R7733 GND.n5036 GND.n2011 19.3944
R7734 GND.n5032 GND.n2011 19.3944
R7735 GND.n5032 GND.n5031 19.3944
R7736 GND.n5031 GND.n5030 19.3944
R7737 GND.n5030 GND.n2016 19.3944
R7738 GND.n5026 GND.n2016 19.3944
R7739 GND.n5026 GND.n5025 19.3944
R7740 GND.n5025 GND.n5024 19.3944
R7741 GND.n5024 GND.n2021 19.3944
R7742 GND.n5020 GND.n2021 19.3944
R7743 GND.n5018 GND.n2028 19.3944
R7744 GND.n5014 GND.n2028 19.3944
R7745 GND.n5014 GND.n5013 19.3944
R7746 GND.n5005 GND.n4889 19.3944
R7747 GND.n5005 GND.n4891 19.3944
R7748 GND.n5001 GND.n4891 19.3944
R7749 GND.n5001 GND.n5000 19.3944
R7750 GND.n5000 GND.n4999 19.3944
R7751 GND.n4996 GND.n4995 19.3944
R7752 GND.n4995 GND.n4994 19.3944
R7753 GND.n4994 GND.n4908 19.3944
R7754 GND.n4990 GND.n4908 19.3944
R7755 GND.n4990 GND.n4989 19.3944
R7756 GND.n4989 GND.n4988 19.3944
R7757 GND.n4988 GND.n4916 19.3944
R7758 GND.n4984 GND.n4916 19.3944
R7759 GND.n4984 GND.n4983 19.3944
R7760 GND.n4983 GND.n4982 19.3944
R7761 GND.n4982 GND.n4924 19.3944
R7762 GND.n4978 GND.n4977 19.3944
R7763 GND.n4977 GND.n4976 19.3944
R7764 GND.n4976 GND.n4935 19.3944
R7765 GND.n4972 GND.n4935 19.3944
R7766 GND.n4972 GND.n4971 19.3944
R7767 GND.n4971 GND.n4970 19.3944
R7768 GND.n4970 GND.n4943 19.3944
R7769 GND.n4966 GND.n4943 19.3944
R7770 GND.n4966 GND.n4965 19.3944
R7771 GND.n4965 GND.n4964 19.3944
R7772 GND.n4964 GND.n4951 19.3944
R7773 GND.n4849 GND.n4848 19.3944
R7774 GND.n4848 GND.n4847 19.3944
R7775 GND.n4847 GND.n4846 19.3944
R7776 GND.n4846 GND.n4844 19.3944
R7777 GND.n4844 GND.n4841 19.3944
R7778 GND.n4841 GND.n4840 19.3944
R7779 GND.n4840 GND.n4837 19.3944
R7780 GND.n4837 GND.n4836 19.3944
R7781 GND.n4836 GND.n4833 19.3944
R7782 GND.n4833 GND.n4832 19.3944
R7783 GND.n4832 GND.n4829 19.3944
R7784 GND.n4827 GND.n4824 19.3944
R7785 GND.n4824 GND.n4823 19.3944
R7786 GND.n4823 GND.n2984 19.3944
R7787 GND.n4819 GND.n2986 19.3944
R7788 GND.n3385 GND.n2986 19.3944
R7789 GND.n3578 GND.n3385 19.3944
R7790 GND.n3578 GND.n3383 19.3944
R7791 GND.n3613 GND.n3383 19.3944
R7792 GND.n3613 GND.n3612 19.3944
R7793 GND.n3612 GND.n3611 19.3944
R7794 GND.n3611 GND.n3584 19.3944
R7795 GND.n3607 GND.n3584 19.3944
R7796 GND.n3607 GND.n3606 19.3944
R7797 GND.n3606 GND.n3605 19.3944
R7798 GND.n3605 GND.n3604 19.3944
R7799 GND.n3604 GND.n3602 19.3944
R7800 GND.n3602 GND.n3601 19.3944
R7801 GND.n3601 GND.n3593 19.3944
R7802 GND.n3597 GND.n3593 19.3944
R7803 GND.n3597 GND.n3366 19.3944
R7804 GND.n3675 GND.n3366 19.3944
R7805 GND.n3676 GND.n3675 19.3944
R7806 GND.n3678 GND.n3676 19.3944
R7807 GND.n3678 GND.n3364 19.3944
R7808 GND.n3682 GND.n3364 19.3944
R7809 GND.n3682 GND.n3353 19.3944
R7810 GND.n3701 GND.n3353 19.3944
R7811 GND.n3701 GND.n3351 19.3944
R7812 GND.n3706 GND.n3351 19.3944
R7813 GND.n3706 GND.n3345 19.3944
R7814 GND.n3733 GND.n3345 19.3944
R7815 GND.n3733 GND.n3732 19.3944
R7816 GND.n3732 GND.n3731 19.3944
R7817 GND.n3731 GND.n3316 19.3944
R7818 GND.n3751 GND.n3316 19.3944
R7819 GND.n3751 GND.n3314 19.3944
R7820 GND.n3814 GND.n3314 19.3944
R7821 GND.n3804 GND.n3755 19.3944
R7822 GND.n3810 GND.n3755 19.3944
R7823 GND.n3811 GND.n3810 19.3944
R7824 GND.n3772 GND.n3769 19.3944
R7825 GND.n3778 GND.n3769 19.3944
R7826 GND.n3778 GND.n3767 19.3944
R7827 GND.n3782 GND.n3767 19.3944
R7828 GND.n3782 GND.n3765 19.3944
R7829 GND.n3788 GND.n3765 19.3944
R7830 GND.n3788 GND.n3763 19.3944
R7831 GND.n3793 GND.n3763 19.3944
R7832 GND.n3793 GND.n3761 19.3944
R7833 GND.n3799 GND.n3761 19.3944
R7834 GND.n3800 GND.n3799 19.3944
R7835 GND.n3015 GND.n3014 19.3944
R7836 GND.n3018 GND.n3015 19.3944
R7837 GND.n3018 GND.n3011 19.3944
R7838 GND.n4801 GND.n3011 19.3944
R7839 GND.n4801 GND.n4800 19.3944
R7840 GND.n4800 GND.n4799 19.3944
R7841 GND.n4799 GND.n3024 19.3944
R7842 GND.n3068 GND.n3024 19.3944
R7843 GND.n3071 GND.n3068 19.3944
R7844 GND.n3071 GND.n3065 19.3944
R7845 GND.n4773 GND.n3065 19.3944
R7846 GND.n4773 GND.n4772 19.3944
R7847 GND.n4772 GND.n4771 19.3944
R7848 GND.n4771 GND.n3077 19.3944
R7849 GND.n3112 GND.n3077 19.3944
R7850 GND.n3112 GND.n3109 19.3944
R7851 GND.n4753 GND.n3109 19.3944
R7852 GND.n4753 GND.n4752 19.3944
R7853 GND.n4752 GND.n4751 19.3944
R7854 GND.n4751 GND.n3118 19.3944
R7855 GND.n3155 GND.n3118 19.3944
R7856 GND.n3155 GND.n3152 19.3944
R7857 GND.n4732 GND.n3152 19.3944
R7858 GND.n4732 GND.n4731 19.3944
R7859 GND.n4731 GND.n4730 19.3944
R7860 GND.n4730 GND.n3161 19.3944
R7861 GND.n4718 GND.n3161 19.3944
R7862 GND.n4718 GND.n4717 19.3944
R7863 GND.n4717 GND.n4716 19.3944
R7864 GND.n4716 GND.n3181 19.3944
R7865 GND.n4704 GND.n3181 19.3944
R7866 GND.n4704 GND.n4703 19.3944
R7867 GND.n4703 GND.n4702 19.3944
R7868 GND.n4702 GND.n3201 19.3944
R7869 GND.n6292 GND.n1071 19.3944
R7870 GND.n6292 GND.n1069 19.3944
R7871 GND.n6296 GND.n1069 19.3944
R7872 GND.n6296 GND.n1065 19.3944
R7873 GND.n6302 GND.n1065 19.3944
R7874 GND.n6302 GND.n1063 19.3944
R7875 GND.n6306 GND.n1063 19.3944
R7876 GND.n6306 GND.n1059 19.3944
R7877 GND.n6312 GND.n1059 19.3944
R7878 GND.n6312 GND.n1057 19.3944
R7879 GND.n6316 GND.n1057 19.3944
R7880 GND.n6316 GND.n1053 19.3944
R7881 GND.n6322 GND.n1053 19.3944
R7882 GND.n6322 GND.n1051 19.3944
R7883 GND.n6326 GND.n1051 19.3944
R7884 GND.n6326 GND.n1047 19.3944
R7885 GND.n6332 GND.n1047 19.3944
R7886 GND.n6332 GND.n1045 19.3944
R7887 GND.n6336 GND.n1045 19.3944
R7888 GND.n6336 GND.n1041 19.3944
R7889 GND.n6342 GND.n1041 19.3944
R7890 GND.n6342 GND.n1039 19.3944
R7891 GND.n6346 GND.n1039 19.3944
R7892 GND.n6346 GND.n1035 19.3944
R7893 GND.n6352 GND.n1035 19.3944
R7894 GND.n6352 GND.n1033 19.3944
R7895 GND.n6356 GND.n1033 19.3944
R7896 GND.n6356 GND.n1029 19.3944
R7897 GND.n6362 GND.n1029 19.3944
R7898 GND.n6362 GND.n1027 19.3944
R7899 GND.n6366 GND.n1027 19.3944
R7900 GND.n6366 GND.n1023 19.3944
R7901 GND.n6372 GND.n1023 19.3944
R7902 GND.n6372 GND.n1021 19.3944
R7903 GND.n6376 GND.n1021 19.3944
R7904 GND.n6376 GND.n1017 19.3944
R7905 GND.n6382 GND.n1017 19.3944
R7906 GND.n6382 GND.n1015 19.3944
R7907 GND.n6386 GND.n1015 19.3944
R7908 GND.n6386 GND.n1011 19.3944
R7909 GND.n6392 GND.n1011 19.3944
R7910 GND.n6392 GND.n1009 19.3944
R7911 GND.n6396 GND.n1009 19.3944
R7912 GND.n6396 GND.n1005 19.3944
R7913 GND.n6402 GND.n1005 19.3944
R7914 GND.n5422 GND.n1593 19.3944
R7915 GND.n5422 GND.n1591 19.3944
R7916 GND.n5426 GND.n1591 19.3944
R7917 GND.n5426 GND.n1587 19.3944
R7918 GND.n5432 GND.n1587 19.3944
R7919 GND.n5432 GND.n1585 19.3944
R7920 GND.n5436 GND.n1585 19.3944
R7921 GND.n5436 GND.n1581 19.3944
R7922 GND.n5442 GND.n1581 19.3944
R7923 GND.n5442 GND.n1579 19.3944
R7924 GND.n5446 GND.n1579 19.3944
R7925 GND.n5446 GND.n1575 19.3944
R7926 GND.n5452 GND.n1575 19.3944
R7927 GND.n5452 GND.n1573 19.3944
R7928 GND.n5456 GND.n1573 19.3944
R7929 GND.n5456 GND.n1569 19.3944
R7930 GND.n5462 GND.n1569 19.3944
R7931 GND.n5462 GND.n1567 19.3944
R7932 GND.n5466 GND.n1567 19.3944
R7933 GND.n5466 GND.n1563 19.3944
R7934 GND.n5472 GND.n1563 19.3944
R7935 GND.n5472 GND.n1561 19.3944
R7936 GND.n5476 GND.n1561 19.3944
R7937 GND.n5476 GND.n1557 19.3944
R7938 GND.n5482 GND.n1557 19.3944
R7939 GND.n5482 GND.n1555 19.3944
R7940 GND.n5486 GND.n1555 19.3944
R7941 GND.n5486 GND.n1551 19.3944
R7942 GND.n5492 GND.n1551 19.3944
R7943 GND.n5492 GND.n1549 19.3944
R7944 GND.n5496 GND.n1549 19.3944
R7945 GND.n5496 GND.n1545 19.3944
R7946 GND.n5502 GND.n1545 19.3944
R7947 GND.n5502 GND.n1543 19.3944
R7948 GND.n5506 GND.n1543 19.3944
R7949 GND.n5506 GND.n1539 19.3944
R7950 GND.n5512 GND.n1539 19.3944
R7951 GND.n5512 GND.n1537 19.3944
R7952 GND.n5516 GND.n1537 19.3944
R7953 GND.n5516 GND.n1533 19.3944
R7954 GND.n5522 GND.n1533 19.3944
R7955 GND.n5522 GND.n1531 19.3944
R7956 GND.n5526 GND.n1531 19.3944
R7957 GND.n5526 GND.n1527 19.3944
R7958 GND.n5532 GND.n1527 19.3944
R7959 GND.n5532 GND.n1525 19.3944
R7960 GND.n5536 GND.n1525 19.3944
R7961 GND.n5536 GND.n1521 19.3944
R7962 GND.n5542 GND.n1521 19.3944
R7963 GND.n5542 GND.n1519 19.3944
R7964 GND.n5546 GND.n1519 19.3944
R7965 GND.n5546 GND.n1515 19.3944
R7966 GND.n5552 GND.n1515 19.3944
R7967 GND.n5552 GND.n1513 19.3944
R7968 GND.n5556 GND.n1513 19.3944
R7969 GND.n5556 GND.n1509 19.3944
R7970 GND.n5562 GND.n1509 19.3944
R7971 GND.n5562 GND.n1507 19.3944
R7972 GND.n5566 GND.n1507 19.3944
R7973 GND.n5566 GND.n1503 19.3944
R7974 GND.n5572 GND.n1503 19.3944
R7975 GND.n5572 GND.n1501 19.3944
R7976 GND.n5576 GND.n1501 19.3944
R7977 GND.n5576 GND.n1497 19.3944
R7978 GND.n5582 GND.n1497 19.3944
R7979 GND.n5582 GND.n1495 19.3944
R7980 GND.n5586 GND.n1495 19.3944
R7981 GND.n5586 GND.n1491 19.3944
R7982 GND.n5592 GND.n1491 19.3944
R7983 GND.n5592 GND.n1489 19.3944
R7984 GND.n5596 GND.n1489 19.3944
R7985 GND.n5596 GND.n1485 19.3944
R7986 GND.n5602 GND.n1485 19.3944
R7987 GND.n5602 GND.n1483 19.3944
R7988 GND.n5606 GND.n1483 19.3944
R7989 GND.n5606 GND.n1479 19.3944
R7990 GND.n5612 GND.n1479 19.3944
R7991 GND.n5612 GND.n1477 19.3944
R7992 GND.n5616 GND.n1477 19.3944
R7993 GND.n5616 GND.n1473 19.3944
R7994 GND.n5622 GND.n1473 19.3944
R7995 GND.n5622 GND.n1471 19.3944
R7996 GND.n5626 GND.n1471 19.3944
R7997 GND.n5626 GND.n1467 19.3944
R7998 GND.n5632 GND.n1467 19.3944
R7999 GND.n5632 GND.n1465 19.3944
R8000 GND.n5636 GND.n1465 19.3944
R8001 GND.n5636 GND.n1461 19.3944
R8002 GND.n5642 GND.n1461 19.3944
R8003 GND.n5642 GND.n1459 19.3944
R8004 GND.n5646 GND.n1459 19.3944
R8005 GND.n5646 GND.n1455 19.3944
R8006 GND.n5652 GND.n1455 19.3944
R8007 GND.n5652 GND.n1453 19.3944
R8008 GND.n5656 GND.n1453 19.3944
R8009 GND.n5656 GND.n1449 19.3944
R8010 GND.n5662 GND.n1449 19.3944
R8011 GND.n5662 GND.n1447 19.3944
R8012 GND.n5666 GND.n1447 19.3944
R8013 GND.n5666 GND.n1443 19.3944
R8014 GND.n5672 GND.n1443 19.3944
R8015 GND.n5672 GND.n1441 19.3944
R8016 GND.n5676 GND.n1441 19.3944
R8017 GND.n5676 GND.n1437 19.3944
R8018 GND.n5682 GND.n1437 19.3944
R8019 GND.n5682 GND.n1435 19.3944
R8020 GND.n5686 GND.n1435 19.3944
R8021 GND.n5686 GND.n1431 19.3944
R8022 GND.n5692 GND.n1431 19.3944
R8023 GND.n5692 GND.n1429 19.3944
R8024 GND.n5696 GND.n1429 19.3944
R8025 GND.n5696 GND.n1425 19.3944
R8026 GND.n5702 GND.n1425 19.3944
R8027 GND.n5702 GND.n1423 19.3944
R8028 GND.n5706 GND.n1423 19.3944
R8029 GND.n5706 GND.n1419 19.3944
R8030 GND.n5712 GND.n1419 19.3944
R8031 GND.n5712 GND.n1417 19.3944
R8032 GND.n5716 GND.n1417 19.3944
R8033 GND.n5716 GND.n1413 19.3944
R8034 GND.n5722 GND.n1413 19.3944
R8035 GND.n5722 GND.n1411 19.3944
R8036 GND.n5726 GND.n1411 19.3944
R8037 GND.n5726 GND.n1407 19.3944
R8038 GND.n5732 GND.n1407 19.3944
R8039 GND.n5732 GND.n1405 19.3944
R8040 GND.n5736 GND.n1405 19.3944
R8041 GND.n5736 GND.n1401 19.3944
R8042 GND.n5742 GND.n1401 19.3944
R8043 GND.n5742 GND.n1399 19.3944
R8044 GND.n5746 GND.n1399 19.3944
R8045 GND.n5746 GND.n1395 19.3944
R8046 GND.n5752 GND.n1395 19.3944
R8047 GND.n5752 GND.n1393 19.3944
R8048 GND.n5756 GND.n1393 19.3944
R8049 GND.n5756 GND.n1389 19.3944
R8050 GND.n5762 GND.n1389 19.3944
R8051 GND.n5762 GND.n1387 19.3944
R8052 GND.n5766 GND.n1387 19.3944
R8053 GND.n5766 GND.n1383 19.3944
R8054 GND.n5772 GND.n1383 19.3944
R8055 GND.n5772 GND.n1381 19.3944
R8056 GND.n5776 GND.n1381 19.3944
R8057 GND.n5776 GND.n1377 19.3944
R8058 GND.n5782 GND.n1377 19.3944
R8059 GND.n5782 GND.n1375 19.3944
R8060 GND.n5786 GND.n1375 19.3944
R8061 GND.n5786 GND.n1371 19.3944
R8062 GND.n5792 GND.n1371 19.3944
R8063 GND.n5792 GND.n1369 19.3944
R8064 GND.n5796 GND.n1369 19.3944
R8065 GND.n5796 GND.n1365 19.3944
R8066 GND.n5802 GND.n1365 19.3944
R8067 GND.n5802 GND.n1363 19.3944
R8068 GND.n5806 GND.n1363 19.3944
R8069 GND.n5806 GND.n1359 19.3944
R8070 GND.n5812 GND.n1359 19.3944
R8071 GND.n5812 GND.n1357 19.3944
R8072 GND.n5816 GND.n1357 19.3944
R8073 GND.n5816 GND.n1353 19.3944
R8074 GND.n5822 GND.n1353 19.3944
R8075 GND.n5822 GND.n1351 19.3944
R8076 GND.n5826 GND.n1351 19.3944
R8077 GND.n5826 GND.n1347 19.3944
R8078 GND.n5832 GND.n1347 19.3944
R8079 GND.n5832 GND.n1345 19.3944
R8080 GND.n5836 GND.n1345 19.3944
R8081 GND.n5836 GND.n1341 19.3944
R8082 GND.n5842 GND.n1341 19.3944
R8083 GND.n5842 GND.n1339 19.3944
R8084 GND.n5846 GND.n1339 19.3944
R8085 GND.n5846 GND.n1335 19.3944
R8086 GND.n5852 GND.n1335 19.3944
R8087 GND.n5852 GND.n1333 19.3944
R8088 GND.n5856 GND.n1333 19.3944
R8089 GND.n5856 GND.n1329 19.3944
R8090 GND.n5862 GND.n1329 19.3944
R8091 GND.n5862 GND.n1327 19.3944
R8092 GND.n5866 GND.n1327 19.3944
R8093 GND.n5866 GND.n1323 19.3944
R8094 GND.n5872 GND.n1323 19.3944
R8095 GND.n5872 GND.n1321 19.3944
R8096 GND.n5876 GND.n1321 19.3944
R8097 GND.n5876 GND.n1317 19.3944
R8098 GND.n5882 GND.n1317 19.3944
R8099 GND.n5882 GND.n1315 19.3944
R8100 GND.n5886 GND.n1315 19.3944
R8101 GND.n5886 GND.n1311 19.3944
R8102 GND.n5892 GND.n1311 19.3944
R8103 GND.n5892 GND.n1309 19.3944
R8104 GND.n5896 GND.n1309 19.3944
R8105 GND.n5896 GND.n1305 19.3944
R8106 GND.n5902 GND.n1305 19.3944
R8107 GND.n5902 GND.n1303 19.3944
R8108 GND.n5906 GND.n1303 19.3944
R8109 GND.n5906 GND.n1299 19.3944
R8110 GND.n5912 GND.n1299 19.3944
R8111 GND.n5912 GND.n1297 19.3944
R8112 GND.n5916 GND.n1297 19.3944
R8113 GND.n5916 GND.n1293 19.3944
R8114 GND.n5922 GND.n1293 19.3944
R8115 GND.n5922 GND.n1291 19.3944
R8116 GND.n5926 GND.n1291 19.3944
R8117 GND.n5926 GND.n1287 19.3944
R8118 GND.n5932 GND.n1287 19.3944
R8119 GND.n5932 GND.n1285 19.3944
R8120 GND.n5936 GND.n1285 19.3944
R8121 GND.n5936 GND.n1281 19.3944
R8122 GND.n5942 GND.n1281 19.3944
R8123 GND.n5942 GND.n1279 19.3944
R8124 GND.n5946 GND.n1279 19.3944
R8125 GND.n5946 GND.n1275 19.3944
R8126 GND.n5952 GND.n1275 19.3944
R8127 GND.n5952 GND.n1273 19.3944
R8128 GND.n5956 GND.n1273 19.3944
R8129 GND.n5956 GND.n1269 19.3944
R8130 GND.n5962 GND.n1269 19.3944
R8131 GND.n5962 GND.n1267 19.3944
R8132 GND.n5966 GND.n1267 19.3944
R8133 GND.n5966 GND.n1263 19.3944
R8134 GND.n5972 GND.n1263 19.3944
R8135 GND.n5972 GND.n1261 19.3944
R8136 GND.n5976 GND.n1261 19.3944
R8137 GND.n5976 GND.n1257 19.3944
R8138 GND.n5982 GND.n1257 19.3944
R8139 GND.n5982 GND.n1255 19.3944
R8140 GND.n5986 GND.n1255 19.3944
R8141 GND.n5986 GND.n1251 19.3944
R8142 GND.n5992 GND.n1251 19.3944
R8143 GND.n5992 GND.n1249 19.3944
R8144 GND.n5996 GND.n1249 19.3944
R8145 GND.n5996 GND.n1245 19.3944
R8146 GND.n6002 GND.n1245 19.3944
R8147 GND.n6002 GND.n1243 19.3944
R8148 GND.n6006 GND.n1243 19.3944
R8149 GND.n6006 GND.n1239 19.3944
R8150 GND.n6012 GND.n1239 19.3944
R8151 GND.n6012 GND.n1237 19.3944
R8152 GND.n6016 GND.n1237 19.3944
R8153 GND.n6016 GND.n1233 19.3944
R8154 GND.n6022 GND.n1233 19.3944
R8155 GND.n6022 GND.n1231 19.3944
R8156 GND.n6026 GND.n1231 19.3944
R8157 GND.n6026 GND.n1227 19.3944
R8158 GND.n6032 GND.n1227 19.3944
R8159 GND.n6032 GND.n1225 19.3944
R8160 GND.n6036 GND.n1225 19.3944
R8161 GND.n6036 GND.n1221 19.3944
R8162 GND.n6042 GND.n1221 19.3944
R8163 GND.n6042 GND.n1219 19.3944
R8164 GND.n6046 GND.n1219 19.3944
R8165 GND.n6046 GND.n1215 19.3944
R8166 GND.n6052 GND.n1215 19.3944
R8167 GND.n6052 GND.n1213 19.3944
R8168 GND.n6056 GND.n1213 19.3944
R8169 GND.n6056 GND.n1209 19.3944
R8170 GND.n6062 GND.n1209 19.3944
R8171 GND.n6062 GND.n1207 19.3944
R8172 GND.n6066 GND.n1207 19.3944
R8173 GND.n6066 GND.n1203 19.3944
R8174 GND.n6072 GND.n1203 19.3944
R8175 GND.n6072 GND.n1201 19.3944
R8176 GND.n6076 GND.n1201 19.3944
R8177 GND.n6076 GND.n1197 19.3944
R8178 GND.n6082 GND.n1197 19.3944
R8179 GND.n6082 GND.n1195 19.3944
R8180 GND.n6086 GND.n1195 19.3944
R8181 GND.n6086 GND.n1191 19.3944
R8182 GND.n6092 GND.n1191 19.3944
R8183 GND.n6092 GND.n1189 19.3944
R8184 GND.n6096 GND.n1189 19.3944
R8185 GND.n6096 GND.n1185 19.3944
R8186 GND.n6102 GND.n1185 19.3944
R8187 GND.n6102 GND.n1183 19.3944
R8188 GND.n6106 GND.n1183 19.3944
R8189 GND.n6106 GND.n1179 19.3944
R8190 GND.n6112 GND.n1179 19.3944
R8191 GND.n6112 GND.n1177 19.3944
R8192 GND.n6116 GND.n1177 19.3944
R8193 GND.n6116 GND.n1173 19.3944
R8194 GND.n6122 GND.n1173 19.3944
R8195 GND.n6122 GND.n1171 19.3944
R8196 GND.n6126 GND.n1171 19.3944
R8197 GND.n6126 GND.n1167 19.3944
R8198 GND.n6132 GND.n1167 19.3944
R8199 GND.n6132 GND.n1165 19.3944
R8200 GND.n6136 GND.n1165 19.3944
R8201 GND.n6136 GND.n1161 19.3944
R8202 GND.n6142 GND.n1161 19.3944
R8203 GND.n6142 GND.n1159 19.3944
R8204 GND.n6146 GND.n1159 19.3944
R8205 GND.n6146 GND.n1155 19.3944
R8206 GND.n6152 GND.n1155 19.3944
R8207 GND.n6152 GND.n1153 19.3944
R8208 GND.n6156 GND.n1153 19.3944
R8209 GND.n6156 GND.n1149 19.3944
R8210 GND.n6162 GND.n1149 19.3944
R8211 GND.n6162 GND.n1147 19.3944
R8212 GND.n6166 GND.n1147 19.3944
R8213 GND.n6166 GND.n1143 19.3944
R8214 GND.n6172 GND.n1143 19.3944
R8215 GND.n6172 GND.n1141 19.3944
R8216 GND.n6176 GND.n1141 19.3944
R8217 GND.n6176 GND.n1137 19.3944
R8218 GND.n6182 GND.n1137 19.3944
R8219 GND.n6182 GND.n1135 19.3944
R8220 GND.n6186 GND.n1135 19.3944
R8221 GND.n6186 GND.n1131 19.3944
R8222 GND.n6192 GND.n1131 19.3944
R8223 GND.n6192 GND.n1129 19.3944
R8224 GND.n6196 GND.n1129 19.3944
R8225 GND.n6196 GND.n1125 19.3944
R8226 GND.n6202 GND.n1125 19.3944
R8227 GND.n6202 GND.n1123 19.3944
R8228 GND.n6206 GND.n1123 19.3944
R8229 GND.n6206 GND.n1119 19.3944
R8230 GND.n6212 GND.n1119 19.3944
R8231 GND.n6212 GND.n1117 19.3944
R8232 GND.n6216 GND.n1117 19.3944
R8233 GND.n6216 GND.n1113 19.3944
R8234 GND.n6222 GND.n1113 19.3944
R8235 GND.n6222 GND.n1111 19.3944
R8236 GND.n6226 GND.n1111 19.3944
R8237 GND.n6226 GND.n1107 19.3944
R8238 GND.n6232 GND.n1107 19.3944
R8239 GND.n6232 GND.n1105 19.3944
R8240 GND.n6236 GND.n1105 19.3944
R8241 GND.n6236 GND.n1101 19.3944
R8242 GND.n6242 GND.n1101 19.3944
R8243 GND.n6242 GND.n1099 19.3944
R8244 GND.n6246 GND.n1099 19.3944
R8245 GND.n6246 GND.n1095 19.3944
R8246 GND.n6252 GND.n1095 19.3944
R8247 GND.n6252 GND.n1093 19.3944
R8248 GND.n6256 GND.n1093 19.3944
R8249 GND.n6256 GND.n1089 19.3944
R8250 GND.n6262 GND.n1089 19.3944
R8251 GND.n6262 GND.n1087 19.3944
R8252 GND.n6266 GND.n1087 19.3944
R8253 GND.n6266 GND.n1083 19.3944
R8254 GND.n6272 GND.n1083 19.3944
R8255 GND.n6272 GND.n1081 19.3944
R8256 GND.n6276 GND.n1081 19.3944
R8257 GND.n6276 GND.n1077 19.3944
R8258 GND.n6282 GND.n1077 19.3944
R8259 GND.n6282 GND.n1075 19.3944
R8260 GND.n6286 GND.n1075 19.3944
R8261 GND.n4628 GND.n4627 19.3944
R8262 GND.n4627 GND.n4626 19.3944
R8263 GND.n4626 GND.n4625 19.3944
R8264 GND.n4625 GND.n4623 19.3944
R8265 GND.n4623 GND.n4620 19.3944
R8266 GND.n4620 GND.n4619 19.3944
R8267 GND.n4619 GND.n4616 19.3944
R8268 GND.n4616 GND.n4615 19.3944
R8269 GND.n4615 GND.n4612 19.3944
R8270 GND.n4610 GND.n4608 19.3944
R8271 GND.n4608 GND.n4605 19.3944
R8272 GND.n4605 GND.n4604 19.3944
R8273 GND.n4604 GND.n4601 19.3944
R8274 GND.n4601 GND.n4600 19.3944
R8275 GND.n4600 GND.n4597 19.3944
R8276 GND.n4597 GND.n4596 19.3944
R8277 GND.n4596 GND.n4593 19.3944
R8278 GND.n4593 GND.n4592 19.3944
R8279 GND.n4592 GND.n4589 19.3944
R8280 GND.n4587 GND.n4585 19.3944
R8281 GND.n4585 GND.n4582 19.3944
R8282 GND.n4582 GND.n3880 19.3944
R8283 GND.n4634 GND.n3885 19.3944
R8284 GND.n4153 GND.n3885 19.3944
R8285 GND.n4157 GND.n4153 19.3944
R8286 GND.n4160 GND.n4157 19.3944
R8287 GND.n4166 GND.n4160 19.3944
R8288 GND.n4170 GND.n4150 19.3944
R8289 GND.n4173 GND.n4170 19.3944
R8290 GND.n4176 GND.n4173 19.3944
R8291 GND.n4176 GND.n4148 19.3944
R8292 GND.n4180 GND.n4148 19.3944
R8293 GND.n4183 GND.n4180 19.3944
R8294 GND.n4186 GND.n4183 19.3944
R8295 GND.n4186 GND.n4146 19.3944
R8296 GND.n4190 GND.n4146 19.3944
R8297 GND.n4193 GND.n4190 19.3944
R8298 GND.n4199 GND.n4193 19.3944
R8299 GND.n4203 GND.n4144 19.3944
R8300 GND.n4206 GND.n4203 19.3944
R8301 GND.n4209 GND.n4206 19.3944
R8302 GND.n4209 GND.n4142 19.3944
R8303 GND.n4213 GND.n4142 19.3944
R8304 GND.n4216 GND.n4213 19.3944
R8305 GND.n4219 GND.n4216 19.3944
R8306 GND.n4219 GND.n4140 19.3944
R8307 GND.n4223 GND.n4140 19.3944
R8308 GND.n4226 GND.n4223 19.3944
R8309 GND.n4229 GND.n4226 19.3944
R8310 GND.n4540 GND.n3940 19.3944
R8311 GND.n4540 GND.n4539 19.3944
R8312 GND.n4539 GND.n3941 19.3944
R8313 GND.n4288 GND.n3941 19.3944
R8314 GND.n4288 GND.n4286 19.3944
R8315 GND.n4298 GND.n4286 19.3944
R8316 GND.n4298 GND.n4098 19.3944
R8317 GND.n4310 GND.n4098 19.3944
R8318 GND.n4311 GND.n4310 19.3944
R8319 GND.n4313 GND.n4311 19.3944
R8320 GND.n4313 GND.n4094 19.3944
R8321 GND.n4325 GND.n4094 19.3944
R8322 GND.n4326 GND.n4325 19.3944
R8323 GND.n4328 GND.n4326 19.3944
R8324 GND.n4328 GND.n4054 19.3944
R8325 GND.n4351 GND.n4054 19.3944
R8326 GND.n4352 GND.n4351 19.3944
R8327 GND.n4353 GND.n4352 19.3944
R8328 GND.n4357 GND.n4353 19.3944
R8329 GND.n4358 GND.n4357 19.3944
R8330 GND.n4359 GND.n4358 19.3944
R8331 GND.n4466 GND.n4359 19.3944
R8332 GND.n4466 GND.n4465 19.3944
R8333 GND.n4465 GND.n4464 19.3944
R8334 GND.n4464 GND.n4362 19.3944
R8335 GND.n4411 GND.n4362 19.3944
R8336 GND.n4444 GND.n4411 19.3944
R8337 GND.n4444 GND.n4443 19.3944
R8338 GND.n4443 GND.n4442 19.3944
R8339 GND.n4442 GND.n4413 19.3944
R8340 GND.n4432 GND.n4413 19.3944
R8341 GND.n4432 GND.n4431 19.3944
R8342 GND.n4431 GND.n4430 19.3944
R8343 GND.n4430 GND.n794 19.3944
R8344 GND.n6614 GND.n794 19.3944
R8345 GND.n6615 GND.n6614 19.3944
R8346 GND.n6616 GND.n6615 19.3944
R8347 GND.n6616 GND.n789 19.3944
R8348 GND.n6628 GND.n789 19.3944
R8349 GND.n6629 GND.n6628 19.3944
R8350 GND.n6630 GND.n6629 19.3944
R8351 GND.n6630 GND.n784 19.3944
R8352 GND.n6643 GND.n784 19.3944
R8353 GND.n6644 GND.n6643 19.3944
R8354 GND.n6646 GND.n6644 19.3944
R8355 GND.n6646 GND.n6645 19.3944
R8356 GND.n4542 GND.n3936 19.3944
R8357 GND.n4542 GND.n3937 19.3944
R8358 GND.n4291 GND.n3937 19.3944
R8359 GND.n4294 GND.n4291 19.3944
R8360 GND.n4295 GND.n4294 19.3944
R8361 GND.n4295 GND.n3978 19.3944
R8362 GND.n4521 GND.n3978 19.3944
R8363 GND.n4521 GND.n4520 19.3944
R8364 GND.n4520 GND.n4519 19.3944
R8365 GND.n4519 GND.n3982 19.3944
R8366 GND.n4509 GND.n3982 19.3944
R8367 GND.n4509 GND.n4508 19.3944
R8368 GND.n4508 GND.n4507 19.3944
R8369 GND.n4507 GND.n4003 19.3944
R8370 GND.n4497 GND.n4003 19.3944
R8371 GND.n4497 GND.n4496 19.3944
R8372 GND.n4496 GND.n4495 19.3944
R8373 GND.n4495 GND.n4024 19.3944
R8374 GND.n4049 GND.n4024 19.3944
R8375 GND.n4472 GND.n4049 19.3944
R8376 GND.n4472 GND.n4471 19.3944
R8377 GND.n4471 GND.n4470 19.3944
R8378 GND.n4470 GND.n4053 19.3944
R8379 GND.n4460 GND.n4053 19.3944
R8380 GND.n4460 GND.n4459 19.3944
R8381 GND.n4459 GND.n4458 19.3944
R8382 GND.n4458 GND.n557 19.3944
R8383 GND.n6845 GND.n557 19.3944
R8384 GND.n6845 GND.n6844 19.3944
R8385 GND.n6844 GND.n6843 19.3944
R8386 GND.n6843 GND.n561 19.3944
R8387 GND.n6833 GND.n561 19.3944
R8388 GND.n6833 GND.n6832 19.3944
R8389 GND.n6832 GND.n6831 19.3944
R8390 GND.n6831 GND.n581 19.3944
R8391 GND.n6821 GND.n581 19.3944
R8392 GND.n6821 GND.n6820 19.3944
R8393 GND.n6820 GND.n6819 19.3944
R8394 GND.n6819 GND.n601 19.3944
R8395 GND.n6809 GND.n601 19.3944
R8396 GND.n6809 GND.n6808 19.3944
R8397 GND.n6808 GND.n6807 19.3944
R8398 GND.n6807 GND.n622 19.3944
R8399 GND.n6797 GND.n622 19.3944
R8400 GND.n6797 GND.n6796 19.3944
R8401 GND.n6796 GND.n6795 19.3944
R8402 GND.n6698 GND.n6697 19.3944
R8403 GND.n6697 GND.n736 19.3944
R8404 GND.n6692 GND.n736 19.3944
R8405 GND.n6692 GND.n6691 19.3944
R8406 GND.n6691 GND.n6690 19.3944
R8407 GND.n6690 GND.n743 19.3944
R8408 GND.n6685 GND.n743 19.3944
R8409 GND.n6685 GND.n6684 19.3944
R8410 GND.n6684 GND.n6683 19.3944
R8411 GND.n6683 GND.n750 19.3944
R8412 GND.n6678 GND.n750 19.3944
R8413 GND.n6722 GND.n6721 19.3944
R8414 GND.n6721 GND.n715 19.3944
R8415 GND.n6716 GND.n715 19.3944
R8416 GND.n6716 GND.n6715 19.3944
R8417 GND.n6715 GND.n6714 19.3944
R8418 GND.n6714 GND.n722 19.3944
R8419 GND.n6709 GND.n722 19.3944
R8420 GND.n6709 GND.n6708 19.3944
R8421 GND.n6708 GND.n6707 19.3944
R8422 GND.n6707 GND.n729 19.3944
R8423 GND.n6702 GND.n729 19.3944
R8424 GND.n6745 GND.n690 19.3944
R8425 GND.n6745 GND.n695 19.3944
R8426 GND.n6740 GND.n695 19.3944
R8427 GND.n6740 GND.n6739 19.3944
R8428 GND.n6739 GND.n6738 19.3944
R8429 GND.n6738 GND.n701 19.3944
R8430 GND.n6733 GND.n701 19.3944
R8431 GND.n6733 GND.n6732 19.3944
R8432 GND.n6732 GND.n6731 19.3944
R8433 GND.n6731 GND.n708 19.3944
R8434 GND.n6726 GND.n708 19.3944
R8435 GND.n6768 GND.n667 19.3944
R8436 GND.n6768 GND.n673 19.3944
R8437 GND.n6763 GND.n673 19.3944
R8438 GND.n6763 GND.n6762 19.3944
R8439 GND.n6762 GND.n6761 19.3944
R8440 GND.n6761 GND.n680 19.3944
R8441 GND.n6756 GND.n680 19.3944
R8442 GND.n6756 GND.n6755 19.3944
R8443 GND.n6755 GND.n6754 19.3944
R8444 GND.n6754 GND.n687 19.3944
R8445 GND.n6788 GND.n6787 19.3944
R8446 GND.n6787 GND.n6786 19.3944
R8447 GND.n6786 GND.n653 19.3944
R8448 GND.n6781 GND.n653 19.3944
R8449 GND.n6781 GND.n6780 19.3944
R8450 GND.n6780 GND.n6779 19.3944
R8451 GND.n6779 GND.n661 19.3944
R8452 GND.n6774 GND.n661 19.3944
R8453 GND.n6774 GND.n6773 19.3944
R8454 GND.n6672 GND.n6671 19.3944
R8455 GND.n6671 GND.n6670 19.3944
R8456 GND.n6670 GND.n764 19.3944
R8457 GND.n765 GND.n764 19.3944
R8458 GND.n6663 GND.n765 19.3944
R8459 GND.n6663 GND.n6662 19.3944
R8460 GND.n6662 GND.n6661 19.3944
R8461 GND.n6661 GND.n772 19.3944
R8462 GND.n6656 GND.n772 19.3944
R8463 GND.n4277 GND.n4276 19.3944
R8464 GND.n4278 GND.n4277 19.3944
R8465 GND.n4278 GND.n4101 19.3944
R8466 GND.n4284 GND.n4101 19.3944
R8467 GND.n4285 GND.n4284 19.3944
R8468 GND.n4302 GND.n4285 19.3944
R8469 GND.n4302 GND.n4099 19.3944
R8470 GND.n4306 GND.n4099 19.3944
R8471 GND.n4306 GND.n4097 19.3944
R8472 GND.n4317 GND.n4097 19.3944
R8473 GND.n4317 GND.n4095 19.3944
R8474 GND.n4321 GND.n4095 19.3944
R8475 GND.n4321 GND.n4093 19.3944
R8476 GND.n4332 GND.n4093 19.3944
R8477 GND.n4332 GND.n4091 19.3944
R8478 GND.n4347 GND.n4091 19.3944
R8479 GND.n4347 GND.n4346 19.3944
R8480 GND.n4346 GND.n4345 19.3944
R8481 GND.n4345 GND.n4344 19.3944
R8482 GND.n4344 GND.n4342 19.3944
R8483 GND.n4342 GND.n4341 19.3944
R8484 GND.n4341 GND.n529 19.3944
R8485 GND.n6857 GND.n529 19.3944
R8486 GND.n6857 GND.n530 19.3944
R8487 GND.n4450 GND.n530 19.3944
R8488 GND.n4450 GND.n4449 19.3944
R8489 GND.n4449 GND.n4448 19.3944
R8490 GND.n4448 GND.n4410 19.3944
R8491 GND.n4438 GND.n4410 19.3944
R8492 GND.n4438 GND.n4437 19.3944
R8493 GND.n4437 GND.n4436 19.3944
R8494 GND.n4436 GND.n4418 19.3944
R8495 GND.n4426 GND.n4418 19.3944
R8496 GND.n4426 GND.n4425 19.3944
R8497 GND.n4425 GND.n4424 19.3944
R8498 GND.n4424 GND.n793 19.3944
R8499 GND.n6620 GND.n793 19.3944
R8500 GND.n6620 GND.n791 19.3944
R8501 GND.n6624 GND.n791 19.3944
R8502 GND.n6624 GND.n788 19.3944
R8503 GND.n6634 GND.n788 19.3944
R8504 GND.n6634 GND.n786 19.3944
R8505 GND.n6639 GND.n786 19.3944
R8506 GND.n6639 GND.n783 19.3944
R8507 GND.n6650 GND.n783 19.3944
R8508 GND.n6651 GND.n6650 19.3944
R8509 GND.n4267 GND.n4265 19.3944
R8510 GND.n4265 GND.n4262 19.3944
R8511 GND.n4262 GND.n4261 19.3944
R8512 GND.n4261 GND.n4258 19.3944
R8513 GND.n4258 GND.n4257 19.3944
R8514 GND.n4257 GND.n4254 19.3944
R8515 GND.n4254 GND.n4253 19.3944
R8516 GND.n4253 GND.n4250 19.3944
R8517 GND.n4250 GND.n4249 19.3944
R8518 GND.n4547 GND.n4546 19.3944
R8519 GND.n4546 GND.n3928 19.3944
R8520 GND.n3964 GND.n3928 19.3944
R8521 GND.n3964 GND.n3961 19.3944
R8522 GND.n4527 GND.n3961 19.3944
R8523 GND.n4527 GND.n4526 19.3944
R8524 GND.n4526 GND.n4525 19.3944
R8525 GND.n4525 GND.n3970 19.3944
R8526 GND.n4515 GND.n3970 19.3944
R8527 GND.n4515 GND.n4514 19.3944
R8528 GND.n4514 GND.n4513 19.3944
R8529 GND.n4513 GND.n3993 19.3944
R8530 GND.n4503 GND.n3993 19.3944
R8531 GND.n4503 GND.n4502 19.3944
R8532 GND.n4502 GND.n4501 19.3944
R8533 GND.n4501 GND.n4015 19.3944
R8534 GND.n4491 GND.n4015 19.3944
R8535 GND.n4491 GND.n4490 19.3944
R8536 GND.n4044 GND.n4043 19.3944
R8537 GND.n4477 GND.n4476 19.3944
R8538 GND.n6853 GND.n6852 19.3944
R8539 GND.n4454 GND.n540 19.3944
R8540 GND.n6849 GND.n547 19.3944
R8541 GND.n6849 GND.n548 19.3944
R8542 GND.n6839 GND.n548 19.3944
R8543 GND.n6839 GND.n6838 19.3944
R8544 GND.n6838 GND.n6837 19.3944
R8545 GND.n6837 GND.n571 19.3944
R8546 GND.n6827 GND.n571 19.3944
R8547 GND.n6827 GND.n6826 19.3944
R8548 GND.n6826 GND.n6825 19.3944
R8549 GND.n6825 GND.n592 19.3944
R8550 GND.n6815 GND.n592 19.3944
R8551 GND.n6815 GND.n6814 19.3944
R8552 GND.n6814 GND.n6813 19.3944
R8553 GND.n6813 GND.n612 19.3944
R8554 GND.n6803 GND.n612 19.3944
R8555 GND.n6803 GND.n6802 19.3944
R8556 GND.n6802 GND.n6801 19.3944
R8557 GND.n6801 GND.n633 19.3944
R8558 GND.n6791 GND.n633 19.3944
R8559 GND.n5323 GND.n1687 19.3944
R8560 GND.n1691 GND.n1687 19.3944
R8561 GND.n5316 GND.n1691 19.3944
R8562 GND.n5316 GND.n5315 19.3944
R8563 GND.n5315 GND.n5314 19.3944
R8564 GND.n5314 GND.n1696 19.3944
R8565 GND.n5308 GND.n1696 19.3944
R8566 GND.n5308 GND.n5307 19.3944
R8567 GND.n5307 GND.n5306 19.3944
R8568 GND.n5306 GND.n1704 19.3944
R8569 GND.n5300 GND.n1704 19.3944
R8570 GND.n5300 GND.n5299 19.3944
R8571 GND.n5299 GND.n5298 19.3944
R8572 GND.n5298 GND.n1712 19.3944
R8573 GND.n5292 GND.n1712 19.3944
R8574 GND.n5292 GND.n5291 19.3944
R8575 GND.n5291 GND.n5290 19.3944
R8576 GND.n5290 GND.n1720 19.3944
R8577 GND.n5284 GND.n1720 19.3944
R8578 GND.n5284 GND.n5283 19.3944
R8579 GND.n5283 GND.n5282 19.3944
R8580 GND.n5282 GND.n1728 19.3944
R8581 GND.n5276 GND.n1728 19.3944
R8582 GND.n5276 GND.n5275 19.3944
R8583 GND.n5275 GND.n5274 19.3944
R8584 GND.n5274 GND.n1736 19.3944
R8585 GND.n5268 GND.n1736 19.3944
R8586 GND.n5268 GND.n5267 19.3944
R8587 GND.n5267 GND.n5266 19.3944
R8588 GND.n5266 GND.n1744 19.3944
R8589 GND.n5260 GND.n1744 19.3944
R8590 GND.n5260 GND.n5259 19.3944
R8591 GND.n5259 GND.n5258 19.3944
R8592 GND.n5258 GND.n1752 19.3944
R8593 GND.n5252 GND.n1752 19.3944
R8594 GND.n5252 GND.n5251 19.3944
R8595 GND.n5251 GND.n5250 19.3944
R8596 GND.n5250 GND.n1760 19.3944
R8597 GND.n5244 GND.n1760 19.3944
R8598 GND.n5244 GND.n5243 19.3944
R8599 GND.n5243 GND.n5242 19.3944
R8600 GND.n5242 GND.n1768 19.3944
R8601 GND.n5236 GND.n1768 19.3944
R8602 GND.n5236 GND.n5235 19.3944
R8603 GND.n5235 GND.n5234 19.3944
R8604 GND.n5234 GND.n1776 19.3944
R8605 GND.n5228 GND.n1776 19.3944
R8606 GND.n5228 GND.n5227 19.3944
R8607 GND.n5227 GND.n5226 19.3944
R8608 GND.n5226 GND.n1784 19.3944
R8609 GND.n5220 GND.n1784 19.3944
R8610 GND.n5220 GND.n5219 19.3944
R8611 GND.n5219 GND.n5218 19.3944
R8612 GND.n5218 GND.n1792 19.3944
R8613 GND.n5212 GND.n1792 19.3944
R8614 GND.n5212 GND.n5211 19.3944
R8615 GND.n5211 GND.n5210 19.3944
R8616 GND.n5210 GND.n1800 19.3944
R8617 GND.n5204 GND.n1800 19.3944
R8618 GND.n5204 GND.n5203 19.3944
R8619 GND.n5203 GND.n5202 19.3944
R8620 GND.n5202 GND.n1808 19.3944
R8621 GND.n5196 GND.n1808 19.3944
R8622 GND.n5196 GND.n5195 19.3944
R8623 GND.n5195 GND.n5194 19.3944
R8624 GND.n5194 GND.n1816 19.3944
R8625 GND.n5188 GND.n1816 19.3944
R8626 GND.n5188 GND.n5187 19.3944
R8627 GND.n5187 GND.n5186 19.3944
R8628 GND.n5186 GND.n1824 19.3944
R8629 GND.n5180 GND.n1824 19.3944
R8630 GND.n5180 GND.n5179 19.3944
R8631 GND.n5179 GND.n5178 19.3944
R8632 GND.n5178 GND.n1832 19.3944
R8633 GND.n5172 GND.n1832 19.3944
R8634 GND.n5172 GND.n5171 19.3944
R8635 GND.n5171 GND.n5170 19.3944
R8636 GND.n5170 GND.n1840 19.3944
R8637 GND.n5164 GND.n1840 19.3944
R8638 GND.n5164 GND.n5163 19.3944
R8639 GND.n5163 GND.n5162 19.3944
R8640 GND.n5162 GND.n1848 19.3944
R8641 GND.n5156 GND.n1848 19.3944
R8642 GND.n5156 GND.n5155 19.3944
R8643 GND.n5155 GND.n5154 19.3944
R8644 GND.n5154 GND.n1856 19.3944
R8645 GND.n5148 GND.n1856 19.3944
R8646 GND.n5148 GND.n5147 19.3944
R8647 GND.n5147 GND.n5146 19.3944
R8648 GND.n5146 GND.n1864 19.3944
R8649 GND.n5140 GND.n1864 19.3944
R8650 GND.n5140 GND.n5139 19.3944
R8651 GND.n5139 GND.n5138 19.3944
R8652 GND.n5138 GND.n1872 19.3944
R8653 GND.n2556 GND.n1872 19.3944
R8654 GND.n2556 GND.n2553 19.3944
R8655 GND.n2560 GND.n2553 19.3944
R8656 GND.n2560 GND.n2551 19.3944
R8657 GND.n2583 GND.n2551 19.3944
R8658 GND.n2583 GND.n2582 19.3944
R8659 GND.n2582 GND.n2581 19.3944
R8660 GND.n2581 GND.n2566 19.3944
R8661 GND.n2577 GND.n2566 19.3944
R8662 GND.n2577 GND.n2576 19.3944
R8663 GND.n2576 GND.n2575 19.3944
R8664 GND.n2575 GND.n2573 19.3944
R8665 GND.n2573 GND.n2219 19.3944
R8666 GND.n2639 GND.n2219 19.3944
R8667 GND.n2639 GND.n2217 19.3944
R8668 GND.n2658 GND.n2217 19.3944
R8669 GND.n2658 GND.n2657 19.3944
R8670 GND.n2657 GND.n2656 19.3944
R8671 GND.n2656 GND.n2645 19.3944
R8672 GND.n2648 GND.n2647 19.3944
R8673 GND.n2756 GND.n2755 19.3944
R8674 GND.n2753 GND.n2162 19.3944
R8675 GND.n2739 GND.n2702 19.3944
R8676 GND.n2737 GND.n2736 19.3944
R8677 GND.n2736 GND.n2704 19.3944
R8678 GND.n2730 GND.n2704 19.3944
R8679 GND.n2730 GND.n2729 19.3944
R8680 GND.n2729 GND.n2728 19.3944
R8681 GND.n2728 GND.n2710 19.3944
R8682 GND.n2724 GND.n2710 19.3944
R8683 GND.n2724 GND.n2723 19.3944
R8684 GND.n2723 GND.n2722 19.3944
R8685 GND.n2722 GND.n2720 19.3944
R8686 GND.n2720 GND.n2095 19.3944
R8687 GND.n2095 GND.n2093 19.3944
R8688 GND.n2827 GND.n2093 19.3944
R8689 GND.n2827 GND.n2091 19.3944
R8690 GND.n2834 GND.n2091 19.3944
R8691 GND.n2834 GND.n2833 19.3944
R8692 GND.n2833 GND.n2065 19.3944
R8693 GND.n2065 GND.n2063 19.3944
R8694 GND.n2913 GND.n2063 19.3944
R8695 GND.n2913 GND.n2061 19.3944
R8696 GND.n4885 GND.n2061 19.3944
R8697 GND.n4885 GND.n4884 19.3944
R8698 GND.n4884 GND.n4883 19.3944
R8699 GND.n4883 GND.n2919 19.3944
R8700 GND.n4877 GND.n2919 19.3944
R8701 GND.n4877 GND.n4876 19.3944
R8702 GND.n4876 GND.n4875 19.3944
R8703 GND.n4875 GND.n2927 19.3944
R8704 GND.n4863 GND.n2927 19.3944
R8705 GND.n4863 GND.n4862 19.3944
R8706 GND.n4862 GND.n4861 19.3944
R8707 GND.n4861 GND.n2945 19.3944
R8708 GND.n3545 GND.n2945 19.3944
R8709 GND.n3550 GND.n3545 19.3944
R8710 GND.n3550 GND.n3000 19.3944
R8711 GND.n4808 GND.n3000 19.3944
R8712 GND.n4808 GND.n4807 19.3944
R8713 GND.n4807 GND.n4806 19.3944
R8714 GND.n4806 GND.n3004 19.3944
R8715 GND.n3043 GND.n3004 19.3944
R8716 GND.n3043 GND.n3040 19.3944
R8717 GND.n4787 GND.n3040 19.3944
R8718 GND.n4787 GND.n4786 19.3944
R8719 GND.n4786 GND.n4785 19.3944
R8720 GND.n4785 GND.n3049 19.3944
R8721 GND.n3087 GND.n3049 19.3944
R8722 GND.n3087 GND.n3084 19.3944
R8723 GND.n4766 GND.n3084 19.3944
R8724 GND.n4766 GND.n4765 19.3944
R8725 GND.n4765 GND.n4764 19.3944
R8726 GND.n4764 GND.n3093 19.3944
R8727 GND.n3137 GND.n3093 19.3944
R8728 GND.n3140 GND.n3137 19.3944
R8729 GND.n3140 GND.n3134 19.3944
R8730 GND.n4739 GND.n3134 19.3944
R8731 GND.n4739 GND.n4738 19.3944
R8732 GND.n4738 GND.n4737 19.3944
R8733 GND.n4737 GND.n3146 19.3944
R8734 GND.n3332 GND.n3146 19.3944
R8735 GND.n3332 GND.n3329 19.3944
R8736 GND.n3336 GND.n3329 19.3944
R8737 GND.n3336 GND.n3327 19.3944
R8738 GND.n3340 GND.n3327 19.3944
R8739 GND.n3340 GND.n3325 19.3944
R8740 GND.n3740 GND.n3325 19.3944
R8741 GND.n3740 GND.n3323 19.3944
R8742 GND.n3747 GND.n3323 19.3944
R8743 GND.n3747 GND.n3746 19.3944
R8744 GND.n3746 GND.n3218 19.3944
R8745 GND.n4689 GND.n3218 19.3944
R8746 GND.n4689 GND.n4688 19.3944
R8747 GND.n4688 GND.n4687 19.3944
R8748 GND.n4687 GND.n3222 19.3944
R8749 GND.n4675 GND.n3222 19.3944
R8750 GND.n4675 GND.n4674 19.3944
R8751 GND.n4674 GND.n4673 19.3944
R8752 GND.n4673 GND.n3240 19.3944
R8753 GND.n4113 GND.n3240 19.3944
R8754 GND.n4119 GND.n4113 19.3944
R8755 GND.n4119 GND.n4118 19.3944
R8756 GND.n4118 GND.n4109 19.3944
R8757 GND.n4126 GND.n4109 19.3944
R8758 GND.n4126 GND.n4107 19.3944
R8759 GND.n4133 GND.n4107 19.3944
R8760 GND.n4133 GND.n4132 19.3944
R8761 GND.n4132 GND.n3947 19.3944
R8762 GND.n4534 GND.n3947 19.3944
R8763 GND.n4534 GND.n4533 19.3944
R8764 GND.n4533 GND.n4532 19.3944
R8765 GND.n4532 GND.n3951 19.3944
R8766 GND.n4065 GND.n3951 19.3944
R8767 GND.n4069 GND.n4065 19.3944
R8768 GND.n4069 GND.n4063 19.3944
R8769 GND.n4073 GND.n4063 19.3944
R8770 GND.n4073 GND.n4061 19.3944
R8771 GND.n4077 GND.n4061 19.3944
R8772 GND.n4077 GND.n4059 19.3944
R8773 GND.n4081 GND.n4059 19.3944
R8774 GND.n4081 GND.n4057 19.3944
R8775 GND.n4088 GND.n4057 19.3944
R8776 GND.n4088 GND.n4087 19.3944
R8777 GND.n4087 GND.n4036 19.3944
R8778 GND.n4485 GND.n4036 19.3944
R8779 GND.n4483 GND.n4482 19.3944
R8780 GND.n4376 GND.n4374 19.3944
R8781 GND.n4380 GND.n4373 19.3944
R8782 GND.n4404 GND.n4382 19.3944
R8783 GND.n4402 GND.n4401 19.3944
R8784 GND.n4401 GND.n4384 19.3944
R8785 GND.n4397 GND.n4384 19.3944
R8786 GND.n4397 GND.n4396 19.3944
R8787 GND.n4396 GND.n4395 19.3944
R8788 GND.n4395 GND.n4392 19.3944
R8789 GND.n4392 GND.n799 19.3944
R8790 GND.n6609 GND.n799 19.3944
R8791 GND.n6609 GND.n6608 19.3944
R8792 GND.n6608 GND.n6607 19.3944
R8793 GND.n6607 GND.n803 19.3944
R8794 GND.n6603 GND.n803 19.3944
R8795 GND.n6603 GND.n6602 19.3944
R8796 GND.n6602 GND.n6601 19.3944
R8797 GND.n6601 GND.n809 19.3944
R8798 GND.n6597 GND.n809 19.3944
R8799 GND.n6597 GND.n6596 19.3944
R8800 GND.n6596 GND.n6595 19.3944
R8801 GND.n6595 GND.n815 19.3944
R8802 GND.n6590 GND.n815 19.3944
R8803 GND.n6590 GND.n6589 19.3944
R8804 GND.n6589 GND.n6588 19.3944
R8805 GND.n6588 GND.n821 19.3944
R8806 GND.n6582 GND.n821 19.3944
R8807 GND.n6582 GND.n6581 19.3944
R8808 GND.n6581 GND.n6580 19.3944
R8809 GND.n6580 GND.n830 19.3944
R8810 GND.n6574 GND.n830 19.3944
R8811 GND.n6574 GND.n6573 19.3944
R8812 GND.n6573 GND.n6572 19.3944
R8813 GND.n6572 GND.n838 19.3944
R8814 GND.n6566 GND.n838 19.3944
R8815 GND.n6566 GND.n6565 19.3944
R8816 GND.n6565 GND.n6564 19.3944
R8817 GND.n6564 GND.n846 19.3944
R8818 GND.n6558 GND.n846 19.3944
R8819 GND.n6558 GND.n6557 19.3944
R8820 GND.n6557 GND.n6556 19.3944
R8821 GND.n6556 GND.n854 19.3944
R8822 GND.n6550 GND.n854 19.3944
R8823 GND.n6550 GND.n6549 19.3944
R8824 GND.n6549 GND.n6548 19.3944
R8825 GND.n6548 GND.n862 19.3944
R8826 GND.n6542 GND.n862 19.3944
R8827 GND.n6542 GND.n6541 19.3944
R8828 GND.n6541 GND.n6540 19.3944
R8829 GND.n6540 GND.n870 19.3944
R8830 GND.n6534 GND.n870 19.3944
R8831 GND.n6534 GND.n6533 19.3944
R8832 GND.n6533 GND.n6532 19.3944
R8833 GND.n6532 GND.n878 19.3944
R8834 GND.n6526 GND.n878 19.3944
R8835 GND.n6526 GND.n6525 19.3944
R8836 GND.n6525 GND.n6524 19.3944
R8837 GND.n6524 GND.n886 19.3944
R8838 GND.n6518 GND.n886 19.3944
R8839 GND.n6518 GND.n6517 19.3944
R8840 GND.n6517 GND.n6516 19.3944
R8841 GND.n6516 GND.n894 19.3944
R8842 GND.n6510 GND.n894 19.3944
R8843 GND.n6510 GND.n6509 19.3944
R8844 GND.n6509 GND.n6508 19.3944
R8845 GND.n6508 GND.n902 19.3944
R8846 GND.n6502 GND.n902 19.3944
R8847 GND.n6502 GND.n6501 19.3944
R8848 GND.n6501 GND.n6500 19.3944
R8849 GND.n6500 GND.n910 19.3944
R8850 GND.n6494 GND.n910 19.3944
R8851 GND.n6494 GND.n6493 19.3944
R8852 GND.n6493 GND.n6492 19.3944
R8853 GND.n6492 GND.n918 19.3944
R8854 GND.n6486 GND.n918 19.3944
R8855 GND.n6486 GND.n6485 19.3944
R8856 GND.n6485 GND.n6484 19.3944
R8857 GND.n6484 GND.n926 19.3944
R8858 GND.n6478 GND.n926 19.3944
R8859 GND.n6478 GND.n6477 19.3944
R8860 GND.n6477 GND.n6476 19.3944
R8861 GND.n6476 GND.n934 19.3944
R8862 GND.n6470 GND.n934 19.3944
R8863 GND.n6470 GND.n6469 19.3944
R8864 GND.n6469 GND.n6468 19.3944
R8865 GND.n6468 GND.n942 19.3944
R8866 GND.n6462 GND.n942 19.3944
R8867 GND.n6462 GND.n6461 19.3944
R8868 GND.n6461 GND.n6460 19.3944
R8869 GND.n6460 GND.n950 19.3944
R8870 GND.n6454 GND.n950 19.3944
R8871 GND.n6454 GND.n6453 19.3944
R8872 GND.n6453 GND.n6452 19.3944
R8873 GND.n6452 GND.n958 19.3944
R8874 GND.n6446 GND.n958 19.3944
R8875 GND.n6446 GND.n6445 19.3944
R8876 GND.n6445 GND.n6444 19.3944
R8877 GND.n6444 GND.n966 19.3944
R8878 GND.n6438 GND.n966 19.3944
R8879 GND.n6438 GND.n6437 19.3944
R8880 GND.n6437 GND.n6436 19.3944
R8881 GND.n6436 GND.n974 19.3944
R8882 GND.n6430 GND.n974 19.3944
R8883 GND.n6430 GND.n6429 19.3944
R8884 GND.n6429 GND.n6428 19.3944
R8885 GND.n6428 GND.n982 19.3944
R8886 GND.n6422 GND.n982 19.3944
R8887 GND.n6422 GND.n6421 19.3944
R8888 GND.n6421 GND.n6420 19.3944
R8889 GND.n6420 GND.n990 19.3944
R8890 GND.n6414 GND.n990 19.3944
R8891 GND.n6414 GND.n6413 19.3944
R8892 GND.n6413 GND.n6412 19.3944
R8893 GND.n6412 GND.n998 19.3944
R8894 GND.n6406 GND.n998 19.3944
R8895 GND.n6406 GND.n6405 19.3944
R8896 GND.n2343 GND.n2342 19.3944
R8897 GND.n2347 GND.n2342 19.3944
R8898 GND.n2347 GND.n2339 19.3944
R8899 GND.n2353 GND.n2339 19.3944
R8900 GND.n2353 GND.n2337 19.3944
R8901 GND.n2357 GND.n2337 19.3944
R8902 GND.n2357 GND.n2335 19.3944
R8903 GND.n2363 GND.n2335 19.3944
R8904 GND.n2363 GND.n2333 19.3944
R8905 GND.n2375 GND.n2331 19.3944
R8906 GND.n2375 GND.n2329 19.3944
R8907 GND.n2379 GND.n2329 19.3944
R8908 GND.n2379 GND.n2327 19.3944
R8909 GND.n2385 GND.n2327 19.3944
R8910 GND.n2385 GND.n2325 19.3944
R8911 GND.n2389 GND.n2325 19.3944
R8912 GND.n2389 GND.n2323 19.3944
R8913 GND.n2395 GND.n2323 19.3944
R8914 GND.n2395 GND.n2321 19.3944
R8915 GND.n2407 GND.n2319 19.3944
R8916 GND.n2407 GND.n2317 19.3944
R8917 GND.n2411 GND.n2317 19.3944
R8918 GND.n2411 GND.n2315 19.3944
R8919 GND.n2417 GND.n2315 19.3944
R8920 GND.n2417 GND.n2313 19.3944
R8921 GND.n2421 GND.n2313 19.3944
R8922 GND.n2421 GND.n2311 19.3944
R8923 GND.n2427 GND.n2311 19.3944
R8924 GND.n2427 GND.n2309 19.3944
R8925 GND.n2434 GND.n2309 19.3944
R8926 GND.n2440 GND.n2307 19.3944
R8927 GND.n2440 GND.n2305 19.3944
R8928 GND.n2444 GND.n2305 19.3944
R8929 GND.n2444 GND.n2303 19.3944
R8930 GND.n2450 GND.n2303 19.3944
R8931 GND.n2450 GND.n2301 19.3944
R8932 GND.n2454 GND.n2301 19.3944
R8933 GND.n2454 GND.n2299 19.3944
R8934 GND.n2460 GND.n2299 19.3944
R8935 GND.n2460 GND.n2297 19.3944
R8936 GND.n2467 GND.n2297 19.3944
R8937 GND.n2473 GND.n2295 19.3944
R8938 GND.n2473 GND.n2293 19.3944
R8939 GND.n2477 GND.n2293 19.3944
R8940 GND.n2477 GND.n2291 19.3944
R8941 GND.n2483 GND.n2291 19.3944
R8942 GND.n2483 GND.n2289 19.3944
R8943 GND.n2487 GND.n2289 19.3944
R8944 GND.n2487 GND.n2287 19.3944
R8945 GND.n2493 GND.n2287 19.3944
R8946 GND.n2493 GND.n2285 19.3944
R8947 GND.n2497 GND.n2285 19.3944
R8948 GND.n5132 GND.n5131 19.3944
R8949 GND.n5131 GND.n5130 19.3944
R8950 GND.n5130 GND.n1884 19.3944
R8951 GND.n2592 GND.n1884 19.3944
R8952 GND.n2592 GND.n2259 19.3944
R8953 GND.n2598 GND.n2259 19.3944
R8954 GND.n2598 GND.n2597 19.3944
R8955 GND.n2597 GND.n2238 19.3944
R8956 GND.n2616 GND.n2238 19.3944
R8957 GND.n2616 GND.n2236 19.3944
R8958 GND.n2622 GND.n2236 19.3944
R8959 GND.n2622 GND.n2621 19.3944
R8960 GND.n2621 GND.n2204 19.3944
R8961 GND.n2666 GND.n2204 19.3944
R8962 GND.n2666 GND.n2202 19.3944
R8963 GND.n2670 GND.n2202 19.3944
R8964 GND.n2671 GND.n2670 19.3944
R8965 GND.n2671 GND.n2147 19.3944
R8966 GND.n2765 GND.n2764 19.3944
R8967 GND.n2172 GND.n2171 19.3944
R8968 GND.n2748 GND.n2747 19.3944
R8969 GND.n2177 GND.n2176 19.3944
R8970 GND.n2693 GND.n2140 19.3944
R8971 GND.n2771 GND.n2140 19.3944
R8972 GND.n2771 GND.n2770 19.3944
R8973 GND.n2770 GND.n2121 19.3944
R8974 GND.n2790 GND.n2121 19.3944
R8975 GND.n2790 GND.n2119 19.3944
R8976 GND.n2796 GND.n2119 19.3944
R8977 GND.n2796 GND.n2795 19.3944
R8978 GND.n2795 GND.n2100 19.3944
R8979 GND.n2816 GND.n2100 19.3944
R8980 GND.n2816 GND.n2098 19.3944
R8981 GND.n2820 GND.n2098 19.3944
R8982 GND.n2820 GND.n2076 19.3944
R8983 GND.n2896 GND.n2076 19.3944
R8984 GND.n2896 GND.n2074 19.3944
R8985 GND.n2902 GND.n2074 19.3944
R8986 GND.n2902 GND.n2901 19.3944
R8987 GND.n2901 GND.n1992 19.3944
R8988 GND.n5054 GND.n1992 19.3944
R8989 GND.n5416 GND.n5415 19.3944
R8990 GND.n5415 GND.n5414 19.3944
R8991 GND.n5414 GND.n1600 19.3944
R8992 GND.n5408 GND.n1600 19.3944
R8993 GND.n5408 GND.n5407 19.3944
R8994 GND.n5407 GND.n5406 19.3944
R8995 GND.n5406 GND.n1608 19.3944
R8996 GND.n5400 GND.n1608 19.3944
R8997 GND.n5400 GND.n5399 19.3944
R8998 GND.n5399 GND.n5398 19.3944
R8999 GND.n5398 GND.n1616 19.3944
R9000 GND.n5392 GND.n1616 19.3944
R9001 GND.n5392 GND.n5391 19.3944
R9002 GND.n5391 GND.n5390 19.3944
R9003 GND.n5390 GND.n1624 19.3944
R9004 GND.n5384 GND.n1624 19.3944
R9005 GND.n5384 GND.n5383 19.3944
R9006 GND.n5383 GND.n5382 19.3944
R9007 GND.n5382 GND.n1632 19.3944
R9008 GND.n5376 GND.n1632 19.3944
R9009 GND.n5376 GND.n5375 19.3944
R9010 GND.n5375 GND.n5374 19.3944
R9011 GND.n5374 GND.n1640 19.3944
R9012 GND.n5368 GND.n1640 19.3944
R9013 GND.n5368 GND.n5367 19.3944
R9014 GND.n5367 GND.n5366 19.3944
R9015 GND.n5366 GND.n1648 19.3944
R9016 GND.n5360 GND.n1648 19.3944
R9017 GND.n5360 GND.n5359 19.3944
R9018 GND.n5359 GND.n5358 19.3944
R9019 GND.n5358 GND.n1656 19.3944
R9020 GND.n5352 GND.n1656 19.3944
R9021 GND.n5352 GND.n5351 19.3944
R9022 GND.n5351 GND.n5350 19.3944
R9023 GND.n5350 GND.n1664 19.3944
R9024 GND.n5344 GND.n1664 19.3944
R9025 GND.n5344 GND.n5343 19.3944
R9026 GND.n5343 GND.n5342 19.3944
R9027 GND.n5342 GND.n1672 19.3944
R9028 GND.n5336 GND.n1672 19.3944
R9029 GND.n5336 GND.n5335 19.3944
R9030 GND.n5335 GND.n5334 19.3944
R9031 GND.n5334 GND.n1680 19.3944
R9032 GND.n5327 GND.n1680 19.3944
R9033 GND.n5327 GND.n5326 19.3944
R9034 GND.n2510 GND.n2279 19.3944
R9035 GND.n2510 GND.n2277 19.3944
R9036 GND.n2516 GND.n2277 19.3944
R9037 GND.n2516 GND.n2275 19.3944
R9038 GND.n2520 GND.n2275 19.3944
R9039 GND.n2520 GND.n2273 19.3944
R9040 GND.n2526 GND.n2273 19.3944
R9041 GND.n2526 GND.n2271 19.3944
R9042 GND.n2530 GND.n2271 19.3944
R9043 GND.n2542 GND.n2538 19.3944
R9044 GND.n2543 GND.n2542 19.3944
R9045 GND.n2543 GND.n2264 19.3944
R9046 GND.n2547 GND.n2264 19.3944
R9047 GND.n2547 GND.n2251 19.3944
R9048 GND.n2602 GND.n2251 19.3944
R9049 GND.n2602 GND.n2248 19.3944
R9050 GND.n2607 GND.n2248 19.3944
R9051 GND.n2607 GND.n2249 19.3944
R9052 GND.n2249 GND.n2227 19.3944
R9053 GND.n2626 GND.n2227 19.3944
R9054 GND.n2626 GND.n2224 19.3944
R9055 GND.n2633 GND.n2224 19.3944
R9056 GND.n2633 GND.n2225 19.3944
R9057 GND.n2629 GND.n2225 19.3944
R9058 GND.n2629 GND.n2193 19.3944
R9059 GND.n2675 GND.n2193 19.3944
R9060 GND.n2675 GND.n2190 19.3944
R9061 GND.n2679 GND.n2190 19.3944
R9062 GND.n2680 GND.n2679 19.3944
R9063 GND.n2681 GND.n2680 19.3944
R9064 GND.n2681 GND.n2186 19.3944
R9065 GND.n2685 GND.n2186 19.3944
R9066 GND.n2686 GND.n2685 19.3944
R9067 GND.n2687 GND.n2686 19.3944
R9068 GND.n2687 GND.n2184 19.3944
R9069 GND.n2691 GND.n2184 19.3944
R9070 GND.n2691 GND.n2132 19.3944
R9071 GND.n2775 GND.n2132 19.3944
R9072 GND.n2775 GND.n2129 19.3944
R9073 GND.n2780 GND.n2129 19.3944
R9074 GND.n2780 GND.n2130 19.3944
R9075 GND.n2130 GND.n2112 19.3944
R9076 GND.n2800 GND.n2112 19.3944
R9077 GND.n2800 GND.n2109 19.3944
R9078 GND.n2808 GND.n2109 19.3944
R9079 GND.n2808 GND.n2110 19.3944
R9080 GND.n2804 GND.n2110 19.3944
R9081 GND.n2804 GND.n2086 19.3944
R9082 GND.n2889 GND.n2086 19.3944
R9083 GND.n2889 GND.n2087 19.3944
R9084 GND.n2885 GND.n2087 19.3944
R9085 GND.n2885 GND.n2884 19.3944
R9086 GND.n2884 GND.n2883 19.3944
R9087 GND.n2883 GND.n2840 19.3944
R9088 GND.n2879 GND.n2840 19.3944
R9089 GND.n5135 GND.n5134 19.1102
R9090 GND.n2540 GND.n1877 19.1102
R9091 GND.n5128 GND.n1886 19.1102
R9092 GND.n2262 GND.n1889 19.1102
R9093 GND.n2590 GND.n2261 19.1102
R9094 GND.n2587 GND.n2585 19.1102
R9095 GND.n2600 GND.n2253 19.1102
R9096 GND.n2257 GND.n2254 19.1102
R9097 GND.n2609 GND.n2246 19.1102
R9098 GND.n2614 GND.n2240 19.1102
R9099 GND.n2611 GND.n2243 19.1102
R9100 GND.n2624 GND.n2229 19.1102
R9101 GND.n2230 GND.n2221 19.1102
R9102 GND.n2636 GND.n2635 19.1102
R9103 GND.n2664 GND.n2207 19.1102
R9104 GND.n2661 GND.n2209 19.1102
R9105 GND.n2660 GND.n2214 19.1102
R9106 GND.n2673 GND.n2196 19.1102
R9107 GND.n2651 GND.n2198 19.1102
R9108 GND.n2653 GND.n2652 19.1102
R9109 GND.n2762 GND.n2150 19.1102
R9110 GND.n2758 GND.n2158 19.1102
R9111 GND.n2165 GND.n2164 19.1102
R9112 GND.n2751 GND.n2750 19.1102
R9113 GND.n2745 GND.n2167 19.1102
R9114 GND.n2741 GND.n2695 19.1102
R9115 GND.n2699 GND.n2698 19.1102
R9116 GND.n2773 GND.n2134 19.1102
R9117 GND.n2731 GND.n2136 19.1102
R9118 GND.n2788 GND.n2123 19.1102
R9119 GND.n2785 GND.n2125 19.1102
R9120 GND.n2798 GND.n2114 19.1102
R9121 GND.n2711 GND.n2115 19.1102
R9122 GND.n2814 GND.n2102 19.1102
R9123 GND.n2105 GND.n2096 19.1102
R9124 GND.n2823 GND.n2822 19.1102
R9125 GND.n2891 GND.n2084 19.1102
R9126 GND.n2894 GND.n2078 19.1102
R9127 GND.n2837 GND.n2081 19.1102
R9128 GND.n2071 GND.n2066 19.1102
R9129 GND.n2909 GND.n2908 19.1102
R9130 GND.n5056 GND.n1986 19.1102
R9131 GND.n4274 GND.n3930 19.1102
R9132 GND.n4544 GND.n3933 19.1102
R9133 GND.n4537 GND.n4536 19.1102
R9134 GND.n4530 GND.n3954 19.1102
R9135 GND.n4529 GND.n3957 19.1102
R9136 GND.n4300 GND.n3972 19.1102
R9137 GND.n4523 GND.n3975 19.1102
R9138 GND.n4308 GND.n3984 19.1102
R9139 GND.n4517 GND.n3987 19.1102
R9140 GND.n4511 GND.n3998 19.1102
R9141 GND.n4323 GND.n4005 19.1102
R9142 GND.n4505 GND.n4008 19.1102
R9143 GND.n4330 GND.n4017 19.1102
R9144 GND.n4349 GND.n4026 19.1102
R9145 GND.n4493 GND.n4029 19.1102
R9146 GND.n4488 GND.n4487 19.1102
R9147 GND.n4045 GND.n4033 19.1102
R9148 GND.n4479 GND.n4041 19.1102
R9149 GND.n4468 GND.n533 19.1102
R9150 GND.n6855 GND.n535 19.1102
R9151 GND.n4462 GND.n4364 19.1102
R9152 GND.n4456 GND.n4406 19.1102
R9153 GND.n4446 GND.n551 19.1102
R9154 GND.n6847 GND.n554 19.1102
R9155 GND.n4440 GND.n563 19.1102
R9156 GND.n6841 GND.n566 19.1102
R9157 GND.n4434 GND.n573 19.1102
R9158 GND.n6835 GND.n576 19.1102
R9159 GND.n4428 GND.n583 19.1102
R9160 GND.n6829 GND.n586 19.1102
R9161 GND.n6612 GND.n6611 19.1102
R9162 GND.n6823 GND.n596 19.1102
R9163 GND.n6618 GND.n603 19.1102
R9164 GND.n6817 GND.n606 19.1102
R9165 GND.n6626 GND.n614 19.1102
R9166 GND.n6811 GND.n617 19.1102
R9167 GND.n6632 GND.n624 19.1102
R9168 GND.n6805 GND.n627 19.1102
R9169 GND.n6641 GND.n635 19.1102
R9170 GND.n6799 GND.n638 19.1102
R9171 GND.n6648 GND.n644 19.1102
R9172 GND.n6793 GND.n647 19.1102
R9173 GND.n2759 GND.t20 18.4277
R9174 GND.n4452 GND.t24 18.4277
R9175 GND.n5013 GND.n2031 18.4247
R9176 GND.n4635 GND.n3880 18.4247
R9177 GND.n5020 GND.n5019 18.0369
R9178 GND.n4589 GND.n4588 18.0369
R9179 GND.n6749 GND.n687 18.0369
R9180 GND.n2401 GND.n2321 18.0369
R9181 GND.n2836 GND.t122 17.7452
R9182 GND.n3953 GND.t145 17.7452
R9183 GND.n4960 GND.n4959 17.455
R9184 GND.n4271 GND.n4138 17.455
R9185 GND.n6677 GND.n757 17.455
R9186 GND.n2502 GND.n2283 17.455
R9187 GND.n3430 GND.n3422 17.1814
R9188 GND.n3275 GND.n3274 17.1814
R9189 GND.n4817 GND.n2989 17.0627
R9190 GND.n4810 GND.n2997 17.0627
R9191 GND.n4797 GND.n3026 17.0627
R9192 GND.n4789 GND.n3037 17.0627
R9193 GND.n4783 GND.n3051 17.0627
R9194 GND.n4775 GND.n3062 17.0627
R9195 GND.n4769 GND.n4768 17.0627
R9196 GND.n4762 GND.n3095 17.0627
R9197 GND.n4755 GND.n3103 17.0627
R9198 GND.n4755 GND.n3106 17.0627
R9199 GND.n4749 GND.n3120 17.0627
R9200 GND.n4741 GND.n3131 17.0627
R9201 GND.n4735 GND.n4734 17.0627
R9202 GND.n4728 GND.n3163 17.0627
R9203 GND.n3708 GND.n3172 17.0627
R9204 GND.n3736 GND.n3735 17.0627
R9205 GND.t180 GND.n3749 17.0627
R9206 GND.n3816 GND.n3212 17.0627
R9207 GND.n4790 GND.n3035 16.3802
R9208 GND.n4782 GND.n3053 16.3802
R9209 GND.n3699 GND.n3698 16.3802
R9210 GND.n4721 GND.n4720 16.3802
R9211 GND.n2742 GND.t22 15.6977
R9212 GND.n4853 GND.n2955 15.6977
R9213 GND.n3388 GND.n3387 15.6977
R9214 GND.n3652 GND.n3651 15.6977
R9215 GND.n4748 GND.n3123 15.6977
R9216 GND.n3320 GND.n3319 15.6977
R9217 GND.n3824 GND.n3823 15.6977
R9218 GND.n4671 GND.t183 15.6977
R9219 GND.n4474 GND.t8 15.6977
R9220 GND.n226 GND.n224 15.6496
R9221 GND.n249 GND.n247 15.6496
R9222 GND.n182 GND.n180 15.6496
R9223 GND.n205 GND.n203 15.6496
R9224 GND.n138 GND.n136 15.6496
R9225 GND.n161 GND.n159 15.6496
R9226 GND.n94 GND.n92 15.6496
R9227 GND.n117 GND.n115 15.6496
R9228 GND.n50 GND.n48 15.6496
R9229 GND.n73 GND.n71 15.6496
R9230 GND.n7 GND.n5 15.6496
R9231 GND.n30 GND.n28 15.6496
R9232 GND.n513 GND.n511 15.6496
R9233 GND.n490 GND.n488 15.6496
R9234 GND.n469 GND.n467 15.6496
R9235 GND.n446 GND.n444 15.6496
R9236 GND.n425 GND.n423 15.6496
R9237 GND.n402 GND.n400 15.6496
R9238 GND.n381 GND.n379 15.6496
R9239 GND.n358 GND.n356 15.6496
R9240 GND.n337 GND.n335 15.6496
R9241 GND.n314 GND.n312 15.6496
R9242 GND.n294 GND.n292 15.6496
R9243 GND.n271 GND.n269 15.6496
R9244 GND.n3447 GND.n3446 15.3369
R9245 GND.n3278 GND.n3277 15.3369
R9246 GND.n5134 GND.n1877 15.0152
R9247 GND.n2540 GND.n1886 15.0152
R9248 GND.n5128 GND.n1889 15.0152
R9249 GND.n2590 GND.n2585 15.0152
R9250 GND.n2587 GND.n2253 15.0152
R9251 GND.n2600 GND.n2254 15.0152
R9252 GND.n2257 GND.n2246 15.0152
R9253 GND.n2609 GND.n2240 15.0152
R9254 GND.n2614 GND.n2243 15.0152
R9255 GND.n2624 GND.n2230 15.0152
R9256 GND.n2636 GND.n2221 15.0152
R9257 GND.n2635 GND.n2207 15.0152
R9258 GND.n2664 GND.n2209 15.0152
R9259 GND.n2214 GND.n2196 15.0152
R9260 GND.n2673 GND.n2198 15.0152
R9261 GND.n2653 GND.n2651 15.0152
R9262 GND.n2652 GND.n2150 15.0152
R9263 GND.n2762 GND.n2152 15.0152
R9264 GND.n2759 GND.n2758 15.0152
R9265 GND.n2164 GND.n2158 15.0152
R9266 GND.n2751 GND.n2165 15.0152
R9267 GND.n2750 GND.n2167 15.0152
R9268 GND.n2745 GND.n2180 15.0152
R9269 GND.n2742 GND.n2741 15.0152
R9270 GND.n2699 GND.n2695 15.0152
R9271 GND.n2698 GND.n2134 15.0152
R9272 GND.n2773 GND.n2136 15.0152
R9273 GND.n2732 GND.n2731 15.0152
R9274 GND.n2782 GND.n2123 15.0152
R9275 GND.n2788 GND.n2125 15.0152
R9276 GND.n2785 GND.n2114 15.0152
R9277 GND.n2798 GND.n2115 15.0152
R9278 GND.n2712 GND.n2711 15.0152
R9279 GND.n2810 GND.n2102 15.0152
R9280 GND.n2814 GND.n2105 15.0152
R9281 GND.n2823 GND.n2096 15.0152
R9282 GND.n2822 GND.n2084 15.0152
R9283 GND.n2891 GND.n2078 15.0152
R9284 GND.n2894 GND.n2081 15.0152
R9285 GND.n2837 GND.n2836 15.0152
R9286 GND.n2904 GND.n2071 15.0152
R9287 GND.n2909 GND.n2066 15.0152
R9288 GND.n2908 GND.n1986 15.0152
R9289 GND.n5056 GND.n1988 15.0152
R9290 GND.n3616 GND.n3615 15.0152
R9291 GND.n3376 GND.n3375 15.0152
R9292 GND.n3684 GND.n3148 15.0152
R9293 GND.n4714 GND.n3183 15.0152
R9294 GND.n4274 GND.n4135 15.0152
R9295 GND.n4544 GND.n3930 15.0152
R9296 GND.n4537 GND.n3933 15.0152
R9297 GND.n4536 GND.n3944 15.0152
R9298 GND.n3954 GND.n3953 15.0152
R9299 GND.n4530 GND.n4529 15.0152
R9300 GND.n4300 GND.n3957 15.0152
R9301 GND.n4523 GND.n3972 15.0152
R9302 GND.n4308 GND.n3975 15.0152
R9303 GND.n4517 GND.n3984 15.0152
R9304 GND.n4315 GND.n3987 15.0152
R9305 GND.n4511 GND.n3995 15.0152
R9306 GND.n4323 GND.n3998 15.0152
R9307 GND.n4505 GND.n4005 15.0152
R9308 GND.n4330 GND.n4008 15.0152
R9309 GND.n4499 GND.n4017 15.0152
R9310 GND.n4349 GND.n4090 15.0152
R9311 GND.n4493 GND.n4026 15.0152
R9312 GND.n4488 GND.n4029 15.0152
R9313 GND.n4487 GND.n4033 15.0152
R9314 GND.n4474 GND.n4045 15.0152
R9315 GND.n4480 GND.n4479 15.0152
R9316 GND.n4468 GND.n4041 15.0152
R9317 GND.n6855 GND.n533 15.0152
R9318 GND.n4462 GND.n535 15.0152
R9319 GND.n4452 GND.n4364 15.0152
R9320 GND.n4456 GND.n4368 15.0152
R9321 GND.n4446 GND.n4406 15.0152
R9322 GND.n6847 GND.n551 15.0152
R9323 GND.n4440 GND.n554 15.0152
R9324 GND.n6841 GND.n563 15.0152
R9325 GND.n6835 GND.n573 15.0152
R9326 GND.n4428 GND.n576 15.0152
R9327 GND.n6829 GND.n583 15.0152
R9328 GND.n6612 GND.n586 15.0152
R9329 GND.n6618 GND.n596 15.0152
R9330 GND.n6817 GND.n603 15.0152
R9331 GND.n6626 GND.n606 15.0152
R9332 GND.n6811 GND.n614 15.0152
R9333 GND.n6632 GND.n617 15.0152
R9334 GND.n6805 GND.n624 15.0152
R9335 GND.n6799 GND.n635 15.0152
R9336 GND.n6648 GND.n638 15.0152
R9337 GND.n6793 GND.n644 15.0152
R9338 GND.n5038 GND.n5037 14.7399
R9339 GND.n4612 GND.n4611 14.7399
R9340 GND.n6773 GND.n6772 14.7399
R9341 GND.n2369 GND.n2333 14.7399
R9342 GND.n3450 GND.n3449 14.3615
R9343 GND.n4667 GND.n4666 14.3615
R9344 GND.n3529 GND.n2947 14.3327
R9345 GND.n3381 GND.n3008 14.3327
R9346 GND.n3728 GND.n3186 14.3327
R9347 GND.t226 GND.n3224 14.3327
R9348 GND.n4684 GND.n3226 14.3327
R9349 GND.n3254 GND.n3253 13.9828
R9350 GND.t89 GND.n2261 13.6503
R9351 GND.n3532 GND.t167 13.6503
R9352 GND.n3372 GND.n3081 13.6503
R9353 GND.n4742 GND.n3129 13.6503
R9354 GND.n4707 GND.n4706 13.6503
R9355 GND.t109 GND.n627 13.6503
R9356 GND.n2875 GND.n2870 13.1884
R9357 GND.n3448 GND.n3416 13.1884
R9358 GND.n3443 GND.n3442 13.1884
R9359 GND.n3442 GND.n3441 13.1884
R9360 GND.n3436 GND.n3435 13.1884
R9361 GND.n3435 GND.n3434 13.1884
R9362 GND.n3255 GND.n3252 13.1884
R9363 GND.n3259 GND.n3252 13.1884
R9364 GND.n3265 GND.n3250 13.1884
R9365 GND.n3266 GND.n3265 13.1884
R9366 GND.n6656 GND.n6655 13.1884
R9367 GND.n4249 GND.n4244 13.1884
R9368 GND.n2530 GND.n2269 13.1884
R9369 GND.n2661 GND.t39 12.9678
R9370 GND.n2782 GND.t31 12.9678
R9371 GND.n4866 GND.n2937 12.9678
R9372 GND.n3553 GND.t135 12.9678
R9373 GND.n4796 GND.n3029 12.9678
R9374 GND.n4776 GND.n3059 12.9678
R9375 GND.n3692 GND.n3358 12.9678
R9376 GND.n3344 GND.n3341 12.9678
R9377 GND.n4693 GND.t170 12.9678
R9378 GND.n4499 GND.t14 12.9678
R9379 GND.n4434 GND.t11 12.9678
R9380 GND.n227 GND.n223 12.8005
R9381 GND.n250 GND.n246 12.8005
R9382 GND.n183 GND.n179 12.8005
R9383 GND.n206 GND.n202 12.8005
R9384 GND.n139 GND.n135 12.8005
R9385 GND.n162 GND.n158 12.8005
R9386 GND.n95 GND.n91 12.8005
R9387 GND.n118 GND.n114 12.8005
R9388 GND.n51 GND.n47 12.8005
R9389 GND.n74 GND.n70 12.8005
R9390 GND.n8 GND.n4 12.8005
R9391 GND.n31 GND.n27 12.8005
R9392 GND.n2877 GND.n2875 12.8005
R9393 GND.n6655 GND.n779 12.8005
R9394 GND.n514 GND.n510 12.8005
R9395 GND.n491 GND.n487 12.8005
R9396 GND.n470 GND.n466 12.8005
R9397 GND.n447 GND.n443 12.8005
R9398 GND.n426 GND.n422 12.8005
R9399 GND.n403 GND.n399 12.8005
R9400 GND.n382 GND.n378 12.8005
R9401 GND.n359 GND.n355 12.8005
R9402 GND.n338 GND.n334 12.8005
R9403 GND.n315 GND.n311 12.8005
R9404 GND.n295 GND.n291 12.8005
R9405 GND.n272 GND.n268 12.8005
R9406 GND.n4245 GND.n4244 12.8005
R9407 GND.n2535 GND.n2269 12.8005
R9408 GND.n4811 GND.n2995 12.2853
R9409 GND.n4761 GND.n3097 12.2853
R9410 GND.n3673 GND.n3672 12.2853
R9411 GND.n4700 GND.n3203 12.2853
R9412 GND.n4691 GND.n3215 12.2853
R9413 GND.n231 GND.n230 12.0247
R9414 GND.n254 GND.n253 12.0247
R9415 GND.n187 GND.n186 12.0247
R9416 GND.n210 GND.n209 12.0247
R9417 GND.n143 GND.n142 12.0247
R9418 GND.n166 GND.n165 12.0247
R9419 GND.n99 GND.n98 12.0247
R9420 GND.n122 GND.n121 12.0247
R9421 GND.n55 GND.n54 12.0247
R9422 GND.n78 GND.n77 12.0247
R9423 GND.n12 GND.n11 12.0247
R9424 GND.n35 GND.n34 12.0247
R9425 GND.n518 GND.n517 12.0247
R9426 GND.n495 GND.n494 12.0247
R9427 GND.n474 GND.n473 12.0247
R9428 GND.n451 GND.n450 12.0247
R9429 GND.n430 GND.n429 12.0247
R9430 GND.n407 GND.n406 12.0247
R9431 GND.n386 GND.n385 12.0247
R9432 GND.n363 GND.n362 12.0247
R9433 GND.n342 GND.n341 12.0247
R9434 GND.n319 GND.n318 12.0247
R9435 GND.n299 GND.n298 12.0247
R9436 GND.n276 GND.n275 12.0247
R9437 GND.n3543 GND.t205 11.6028
R9438 GND.n3627 GND.n3626 11.6028
R9439 GND.n3628 GND.n3627 11.6028
R9440 GND.n4727 GND.n3166 11.6028
R9441 GND.n3709 GND.n3166 11.6028
R9442 GND.n3816 GND.t93 11.6028
R9443 GND.n4670 GND.n3244 11.6028
R9444 GND.n234 GND.n221 11.249
R9445 GND.n257 GND.n244 11.249
R9446 GND.n190 GND.n177 11.249
R9447 GND.n213 GND.n200 11.249
R9448 GND.n146 GND.n133 11.249
R9449 GND.n169 GND.n156 11.249
R9450 GND.n102 GND.n89 11.249
R9451 GND.n125 GND.n112 11.249
R9452 GND.n58 GND.n45 11.249
R9453 GND.n81 GND.n68 11.249
R9454 GND.n15 GND.n2 11.249
R9455 GND.n38 GND.n25 11.249
R9456 GND.n5037 GND.n5036 11.249
R9457 GND.n4611 GND.n4610 11.249
R9458 GND.n6772 GND.n667 11.249
R9459 GND.n521 GND.n508 11.249
R9460 GND.n498 GND.n485 11.249
R9461 GND.n477 GND.n464 11.249
R9462 GND.n454 GND.n441 11.249
R9463 GND.n433 GND.n420 11.249
R9464 GND.n410 GND.n397 11.249
R9465 GND.n389 GND.n376 11.249
R9466 GND.n366 GND.n353 11.249
R9467 GND.n345 GND.n332 11.249
R9468 GND.n322 GND.n309 11.249
R9469 GND.n302 GND.n289 11.249
R9470 GND.n279 GND.n266 11.249
R9471 GND.n2369 GND.n2331 11.249
R9472 GND.n2930 GND.t186 10.9203
R9473 GND.n3552 GND.t116 10.9203
R9474 GND.n3557 GND.n2995 10.9203
R9475 GND.n3656 GND.n3097 10.9203
R9476 GND.n3673 GND.n3368 10.9203
R9477 GND.n4700 GND.n4699 10.9203
R9478 GND.n3279 GND.n3248 10.8611
R9479 GND.n3297 GND.n3295 10.6151
R9480 GND.n3873 GND.n3297 10.6151
R9481 GND.n3873 GND.n3872 10.6151
R9482 GND.n3870 GND.n3301 10.6151
R9483 GND.n3865 GND.n3301 10.6151
R9484 GND.n3865 GND.n3864 10.6151
R9485 GND.n3864 GND.n3863 10.6151
R9486 GND.n3863 GND.n3304 10.6151
R9487 GND.n3858 GND.n3304 10.6151
R9488 GND.n3858 GND.n3857 10.6151
R9489 GND.n3857 GND.n3856 10.6151
R9490 GND.n3856 GND.n3307 10.6151
R9491 GND.n3851 GND.n3307 10.6151
R9492 GND.n3851 GND.n3850 10.6151
R9493 GND.n3850 GND.n3849 10.6151
R9494 GND.n3522 GND.n3521 10.6151
R9495 GND.n3525 GND.n3522 10.6151
R9496 GND.n3526 GND.n3525 10.6151
R9497 GND.n3527 GND.n3526 10.6151
R9498 GND.n3527 GND.n3391 10.6151
R9499 GND.n3535 GND.n3391 10.6151
R9500 GND.n3536 GND.n3535 10.6151
R9501 GND.n3538 GND.n3536 10.6151
R9502 GND.n3539 GND.n3538 10.6151
R9503 GND.n3540 GND.n3539 10.6151
R9504 GND.n3555 GND.n3540 10.6151
R9505 GND.n3556 GND.n3555 10.6151
R9506 GND.n3559 GND.n3556 10.6151
R9507 GND.n3560 GND.n3559 10.6151
R9508 GND.n3561 GND.n3560 10.6151
R9509 GND.n3565 GND.n3561 10.6151
R9510 GND.n3565 GND.n3564 10.6151
R9511 GND.n3564 GND.n3563 10.6151
R9512 GND.n3563 GND.n3379 10.6151
R9513 GND.n3618 GND.n3379 10.6151
R9514 GND.n3619 GND.n3618 10.6151
R9515 GND.n3622 GND.n3619 10.6151
R9516 GND.n3623 GND.n3622 10.6151
R9517 GND.n3624 GND.n3623 10.6151
R9518 GND.n3630 GND.n3624 10.6151
R9519 GND.n3631 GND.n3630 10.6151
R9520 GND.n3634 GND.n3631 10.6151
R9521 GND.n3635 GND.n3634 10.6151
R9522 GND.n3636 GND.n3635 10.6151
R9523 GND.n3640 GND.n3636 10.6151
R9524 GND.n3640 GND.n3639 10.6151
R9525 GND.n3639 GND.n3638 10.6151
R9526 GND.n3638 GND.n3370 10.6151
R9527 GND.n3654 GND.n3370 10.6151
R9528 GND.n3655 GND.n3654 10.6151
R9529 GND.n3658 GND.n3655 10.6151
R9530 GND.n3659 GND.n3658 10.6151
R9531 GND.n3660 GND.n3659 10.6151
R9532 GND.n3670 GND.n3660 10.6151
R9533 GND.n3670 GND.n3669 10.6151
R9534 GND.n3669 GND.n3668 10.6151
R9535 GND.n3668 GND.n3665 10.6151
R9536 GND.n3665 GND.n3664 10.6151
R9537 GND.n3664 GND.n3661 10.6151
R9538 GND.n3661 GND.n3356 10.6151
R9539 GND.n3694 GND.n3356 10.6151
R9540 GND.n3695 GND.n3694 10.6151
R9541 GND.n3696 GND.n3695 10.6151
R9542 GND.n3696 GND.n3350 10.6151
R9543 GND.n3711 GND.n3350 10.6151
R9544 GND.n3712 GND.n3711 10.6151
R9545 GND.n3713 GND.n3712 10.6151
R9546 GND.n3713 GND.n3349 10.6151
R9547 GND.n3717 GND.n3349 10.6151
R9548 GND.n3718 GND.n3717 10.6151
R9549 GND.n3726 GND.n3718 10.6151
R9550 GND.n3726 GND.n3725 10.6151
R9551 GND.n3725 GND.n3724 10.6151
R9552 GND.n3724 GND.n3719 10.6151
R9553 GND.n3720 GND.n3719 10.6151
R9554 GND.n3720 GND.n3312 10.6151
R9555 GND.n3818 GND.n3312 10.6151
R9556 GND.n3819 GND.n3818 10.6151
R9557 GND.n3820 GND.n3819 10.6151
R9558 GND.n3821 GND.n3820 10.6151
R9559 GND.n3821 GND.n3311 10.6151
R9560 GND.n3832 GND.n3311 10.6151
R9561 GND.n3833 GND.n3832 10.6151
R9562 GND.n3835 GND.n3833 10.6151
R9563 GND.n3836 GND.n3835 10.6151
R9564 GND.n3837 GND.n3836 10.6151
R9565 GND.n3837 GND.n3310 10.6151
R9566 GND.n3845 GND.n3310 10.6151
R9567 GND.n3846 GND.n3845 10.6151
R9568 GND.n3490 GND.n3489 10.6151
R9569 GND.n3491 GND.n3490 10.6151
R9570 GND.n3491 GND.n3402 10.6151
R9571 GND.n3498 GND.n3497 10.6151
R9572 GND.n3499 GND.n3498 10.6151
R9573 GND.n3499 GND.n3397 10.6151
R9574 GND.n3505 GND.n3397 10.6151
R9575 GND.n3506 GND.n3505 10.6151
R9576 GND.n3507 GND.n3506 10.6151
R9577 GND.n3507 GND.n3395 10.6151
R9578 GND.n3513 GND.n3395 10.6151
R9579 GND.n3514 GND.n3513 10.6151
R9580 GND.n3515 GND.n3514 10.6151
R9581 GND.n3515 GND.n3393 10.6151
R9582 GND.n3393 GND.n3392 10.6151
R9583 GND.n3454 GND.n3450 10.6151
R9584 GND.n3455 GND.n3454 10.6151
R9585 GND.n3456 GND.n3455 10.6151
R9586 GND.n3456 GND.n3414 10.6151
R9587 GND.n3462 GND.n3414 10.6151
R9588 GND.n3463 GND.n3462 10.6151
R9589 GND.n3464 GND.n3463 10.6151
R9590 GND.n3464 GND.n3412 10.6151
R9591 GND.n3470 GND.n3412 10.6151
R9592 GND.n3471 GND.n3470 10.6151
R9593 GND.n3472 GND.n3471 10.6151
R9594 GND.n3472 GND.n3410 10.6151
R9595 GND.n3479 GND.n3478 10.6151
R9596 GND.n3480 GND.n3479 10.6151
R9597 GND.n3480 GND.n3405 10.6151
R9598 GND.n4666 GND.n4665 10.6151
R9599 GND.n4665 GND.n3280 10.6151
R9600 GND.n4660 GND.n3280 10.6151
R9601 GND.n4660 GND.n4659 10.6151
R9602 GND.n4659 GND.n4658 10.6151
R9603 GND.n4658 GND.n3284 10.6151
R9604 GND.n4653 GND.n3284 10.6151
R9605 GND.n4653 GND.n4652 10.6151
R9606 GND.n4652 GND.n4651 10.6151
R9607 GND.n4651 GND.n3287 10.6151
R9608 GND.n4646 GND.n3287 10.6151
R9609 GND.n4646 GND.n4645 10.6151
R9610 GND.n4643 GND.n3292 10.6151
R9611 GND.n4638 GND.n3292 10.6151
R9612 GND.n4638 GND.n4637 10.6151
R9613 GND.n4870 GND.n2934 10.6151
R9614 GND.n4870 GND.n4869 10.6151
R9615 GND.n4869 GND.n4868 10.6151
R9616 GND.n4868 GND.n2935 10.6151
R9617 GND.n3530 GND.n2935 10.6151
R9618 GND.n3530 GND.n2952 10.6151
R9619 GND.n4857 GND.n2952 10.6151
R9620 GND.n4857 GND.n4856 10.6151
R9621 GND.n4856 GND.n4855 10.6151
R9622 GND.n4855 GND.n2953 10.6151
R9623 GND.n2992 GND.n2953 10.6151
R9624 GND.n4815 GND.n2992 10.6151
R9625 GND.n4815 GND.n4814 10.6151
R9626 GND.n4814 GND.n4813 10.6151
R9627 GND.n4813 GND.n2993 10.6151
R9628 GND.n3573 GND.n2993 10.6151
R9629 GND.n3573 GND.n3572 10.6151
R9630 GND.n3572 GND.n3571 10.6151
R9631 GND.n3571 GND.n3568 10.6151
R9632 GND.n3568 GND.n3032 10.6151
R9633 GND.n4794 GND.n3032 10.6151
R9634 GND.n4794 GND.n4793 10.6151
R9635 GND.n4793 GND.n4792 10.6151
R9636 GND.n4792 GND.n3033 10.6151
R9637 GND.n3056 GND.n3033 10.6151
R9638 GND.n4780 GND.n3056 10.6151
R9639 GND.n4780 GND.n4779 10.6151
R9640 GND.n4779 GND.n4778 10.6151
R9641 GND.n4778 GND.n3057 10.6151
R9642 GND.n3374 GND.n3057 10.6151
R9643 GND.n3646 GND.n3374 10.6151
R9644 GND.n3647 GND.n3646 10.6151
R9645 GND.n3648 GND.n3647 10.6151
R9646 GND.n3648 GND.n3100 10.6151
R9647 GND.n4759 GND.n3100 10.6151
R9648 GND.n4759 GND.n4758 10.6151
R9649 GND.n4758 GND.n4757 10.6151
R9650 GND.n4757 GND.n3101 10.6151
R9651 GND.n3126 GND.n3101 10.6151
R9652 GND.n4746 GND.n3126 10.6151
R9653 GND.n4746 GND.n4745 10.6151
R9654 GND.n4745 GND.n4744 10.6151
R9655 GND.n4744 GND.n3127 10.6151
R9656 GND.n3687 GND.n3127 10.6151
R9657 GND.n3688 GND.n3687 10.6151
R9658 GND.n3690 GND.n3688 10.6151
R9659 GND.n3690 GND.n3689 10.6151
R9660 GND.n3689 GND.n3169 10.6151
R9661 GND.n4725 GND.n3169 10.6151
R9662 GND.n4725 GND.n4724 10.6151
R9663 GND.n4724 GND.n4723 10.6151
R9664 GND.n4723 GND.n3170 10.6151
R9665 GND.n3342 GND.n3170 10.6151
R9666 GND.n3342 GND.n3189 10.6151
R9667 GND.n4711 GND.n3189 10.6151
R9668 GND.n4711 GND.n4710 10.6151
R9669 GND.n4710 GND.n4709 10.6151
R9670 GND.n4709 GND.n3190 10.6151
R9671 GND.n3317 GND.n3190 10.6151
R9672 GND.n3317 GND.n3209 10.6151
R9673 GND.n4697 GND.n3209 10.6151
R9674 GND.n4697 GND.n4696 10.6151
R9675 GND.n4696 GND.n4695 10.6151
R9676 GND.n4695 GND.n3210 10.6151
R9677 GND.n3826 GND.n3210 10.6151
R9678 GND.n3827 GND.n3826 10.6151
R9679 GND.n3827 GND.n3229 10.6151
R9680 GND.n4682 GND.n3229 10.6151
R9681 GND.n4682 GND.n4681 10.6151
R9682 GND.n4681 GND.n4680 10.6151
R9683 GND.n4680 GND.n3230 10.6151
R9684 GND.n3840 GND.n3230 10.6151
R9685 GND.n3840 GND.n3247 10.6151
R9686 GND.n4668 GND.n3247 10.6151
R9687 GND.n235 GND.n219 10.4732
R9688 GND.n258 GND.n242 10.4732
R9689 GND.n191 GND.n175 10.4732
R9690 GND.n214 GND.n198 10.4732
R9691 GND.n147 GND.n131 10.4732
R9692 GND.n170 GND.n154 10.4732
R9693 GND.n103 GND.n87 10.4732
R9694 GND.n126 GND.n110 10.4732
R9695 GND.n59 GND.n43 10.4732
R9696 GND.n82 GND.n66 10.4732
R9697 GND.n16 GND.n0 10.4732
R9698 GND.n39 GND.n23 10.4732
R9699 GND.n522 GND.n506 10.4732
R9700 GND.n499 GND.n483 10.4732
R9701 GND.n478 GND.n462 10.4732
R9702 GND.n455 GND.n439 10.4732
R9703 GND.n434 GND.n418 10.4732
R9704 GND.n411 GND.n395 10.4732
R9705 GND.n390 GND.n374 10.4732
R9706 GND.n367 GND.n351 10.4732
R9707 GND.n346 GND.n330 10.4732
R9708 GND.n323 GND.n307 10.4732
R9709 GND.n303 GND.n287 10.4732
R9710 GND.n280 GND.n264 10.4732
R9711 GND.n2611 GND.t41 10.2378
R9712 GND.n2810 GND.t16 10.2378
R9713 GND.n3523 GND.n2937 10.2378
R9714 GND.n3542 GND.t135 10.2378
R9715 GND.t195 GND.n4803 10.2378
R9716 GND.n3620 GND.n3029 10.2378
R9717 GND.n3632 GND.n3059 10.2378
R9718 GND.n3358 GND.n3354 10.2378
R9719 GND.n3341 GND.n3175 10.2378
R9720 GND.n3729 GND.t99 10.2378
R9721 GND.n3842 GND.n3839 10.2378
R9722 GND.n4315 GND.t4 10.2378
R9723 GND.n6823 GND.t6 10.2378
R9724 GND.t167 GND.n2939 9.55533
R9725 GND.n3576 GND.n3575 9.55533
R9726 GND.t2 GND.n3079 9.55533
R9727 GND.n3650 GND.n3372 9.55533
R9728 GND.n3666 GND.n3129 9.55533
R9729 GND.n3662 GND.t3 9.55533
R9730 GND.n4706 GND.n3195 9.55533
R9731 GND.n237 GND.n236 9.45567
R9732 GND.n260 GND.n259 9.45567
R9733 GND.n193 GND.n192 9.45567
R9734 GND.n216 GND.n215 9.45567
R9735 GND.n149 GND.n148 9.45567
R9736 GND.n172 GND.n171 9.45567
R9737 GND.n105 GND.n104 9.45567
R9738 GND.n128 GND.n127 9.45567
R9739 GND.n61 GND.n60 9.45567
R9740 GND.n84 GND.n83 9.45567
R9741 GND.n18 GND.n17 9.45567
R9742 GND.n41 GND.n40 9.45567
R9743 GND.n524 GND.n523 9.45567
R9744 GND.n501 GND.n500 9.45567
R9745 GND.n480 GND.n479 9.45567
R9746 GND.n457 GND.n456 9.45567
R9747 GND.n436 GND.n435 9.45567
R9748 GND.n413 GND.n412 9.45567
R9749 GND.n392 GND.n391 9.45567
R9750 GND.n369 GND.n368 9.45567
R9751 GND.n348 GND.n347 9.45567
R9752 GND.n325 GND.n324 9.45567
R9753 GND.n305 GND.n304 9.45567
R9754 GND.n282 GND.n281 9.45567
R9755 GND.n3871 GND.n3870 9.36635
R9756 GND.n3497 GND.n3401 9.36635
R9757 GND.n3410 GND.n3409 9.36635
R9758 GND.n4645 GND.n4644 9.36635
R9759 GND.n236 GND.n235 9.3005
R9760 GND.n221 GND.n220 9.3005
R9761 GND.n230 GND.n229 9.3005
R9762 GND.n228 GND.n227 9.3005
R9763 GND.n259 GND.n258 9.3005
R9764 GND.n244 GND.n243 9.3005
R9765 GND.n253 GND.n252 9.3005
R9766 GND.n251 GND.n250 9.3005
R9767 GND.n192 GND.n191 9.3005
R9768 GND.n177 GND.n176 9.3005
R9769 GND.n186 GND.n185 9.3005
R9770 GND.n184 GND.n183 9.3005
R9771 GND.n215 GND.n214 9.3005
R9772 GND.n200 GND.n199 9.3005
R9773 GND.n209 GND.n208 9.3005
R9774 GND.n207 GND.n206 9.3005
R9775 GND.n148 GND.n147 9.3005
R9776 GND.n133 GND.n132 9.3005
R9777 GND.n142 GND.n141 9.3005
R9778 GND.n140 GND.n139 9.3005
R9779 GND.n171 GND.n170 9.3005
R9780 GND.n156 GND.n155 9.3005
R9781 GND.n165 GND.n164 9.3005
R9782 GND.n163 GND.n162 9.3005
R9783 GND.n104 GND.n103 9.3005
R9784 GND.n89 GND.n88 9.3005
R9785 GND.n98 GND.n97 9.3005
R9786 GND.n96 GND.n95 9.3005
R9787 GND.n127 GND.n126 9.3005
R9788 GND.n112 GND.n111 9.3005
R9789 GND.n121 GND.n120 9.3005
R9790 GND.n119 GND.n118 9.3005
R9791 GND.n60 GND.n59 9.3005
R9792 GND.n45 GND.n44 9.3005
R9793 GND.n54 GND.n53 9.3005
R9794 GND.n52 GND.n51 9.3005
R9795 GND.n83 GND.n82 9.3005
R9796 GND.n68 GND.n67 9.3005
R9797 GND.n77 GND.n76 9.3005
R9798 GND.n75 GND.n74 9.3005
R9799 GND.n17 GND.n16 9.3005
R9800 GND.n2 GND.n1 9.3005
R9801 GND.n11 GND.n10 9.3005
R9802 GND.n9 GND.n8 9.3005
R9803 GND.n40 GND.n39 9.3005
R9804 GND.n25 GND.n24 9.3005
R9805 GND.n34 GND.n33 9.3005
R9806 GND.n32 GND.n31 9.3005
R9807 GND.n3769 GND.n3768 9.3005
R9808 GND.n3779 GND.n3778 9.3005
R9809 GND.n3780 GND.n3767 9.3005
R9810 GND.n3782 GND.n3781 9.3005
R9811 GND.n3765 GND.n3764 9.3005
R9812 GND.n3789 GND.n3788 9.3005
R9813 GND.n3790 GND.n3763 9.3005
R9814 GND.n3793 GND.n3792 9.3005
R9815 GND.n3791 GND.n3761 9.3005
R9816 GND.n3799 GND.n3760 9.3005
R9817 GND.n3801 GND.n3800 9.3005
R9818 GND.n3804 GND.n3803 9.3005
R9819 GND.n3802 GND.n3755 9.3005
R9820 GND.n3810 GND.n3754 9.3005
R9821 GND.n3812 GND.n3811 9.3005
R9822 GND.n3772 GND.n3771 9.3005
R9823 GND.n2986 GND.n2985 9.3005
R9824 GND.n3385 GND.n3384 9.3005
R9825 GND.n3579 GND.n3578 9.3005
R9826 GND.n3580 GND.n3383 9.3005
R9827 GND.n3613 GND.n3581 9.3005
R9828 GND.n3612 GND.n3582 9.3005
R9829 GND.n3611 GND.n3583 9.3005
R9830 GND.n3586 GND.n3584 9.3005
R9831 GND.n3607 GND.n3587 9.3005
R9832 GND.n3606 GND.n3588 9.3005
R9833 GND.n3605 GND.n3589 9.3005
R9834 GND.n3604 GND.n3590 9.3005
R9835 GND.n3602 GND.n3591 9.3005
R9836 GND.n3601 GND.n3592 9.3005
R9837 GND.n3594 GND.n3593 9.3005
R9838 GND.n3597 GND.n3596 9.3005
R9839 GND.n3595 GND.n3366 9.3005
R9840 GND.n3675 GND.n3367 9.3005
R9841 GND.n3676 GND.n3365 9.3005
R9842 GND.n3679 GND.n3678 9.3005
R9843 GND.n3680 GND.n3364 9.3005
R9844 GND.n3682 GND.n3681 9.3005
R9845 GND.n3353 GND.n3352 9.3005
R9846 GND.n3702 GND.n3701 9.3005
R9847 GND.n3703 GND.n3351 9.3005
R9848 GND.n3706 GND.n3705 9.3005
R9849 GND.n3704 GND.n3345 9.3005
R9850 GND.n3733 GND.n3346 9.3005
R9851 GND.n3732 GND.n3347 9.3005
R9852 GND.n3731 GND.n3348 9.3005
R9853 GND.n3316 GND.n3315 9.3005
R9854 GND.n3752 GND.n3751 9.3005
R9855 GND.n3753 GND.n3314 9.3005
R9856 GND.n3814 GND.n3813 9.3005
R9857 GND.n4820 GND.n4819 9.3005
R9858 GND.n4823 GND.n4822 9.3005
R9859 GND.n4824 GND.n2982 9.3005
R9860 GND.n4827 GND.n2981 9.3005
R9861 GND.n4829 GND.n2978 9.3005
R9862 GND.n4832 GND.n2977 9.3005
R9863 GND.n4833 GND.n2976 9.3005
R9864 GND.n4836 GND.n2975 9.3005
R9865 GND.n4837 GND.n2974 9.3005
R9866 GND.n4840 GND.n2973 9.3005
R9867 GND.n4841 GND.n2972 9.3005
R9868 GND.n4844 GND.n2971 9.3005
R9869 GND.n4846 GND.n2970 9.3005
R9870 GND.n4847 GND.n2969 9.3005
R9871 GND.n4848 GND.n2968 9.3005
R9872 GND.n4849 GND.n2967 9.3005
R9873 GND.n4821 GND.n2984 9.3005
R9874 GND.n3015 GND.n3012 9.3005
R9875 GND.n3019 GND.n3018 9.3005
R9876 GND.n3020 GND.n3011 9.3005
R9877 GND.n4801 GND.n3021 9.3005
R9878 GND.n4800 GND.n3022 9.3005
R9879 GND.n4799 GND.n3023 9.3005
R9880 GND.n3066 GND.n3024 9.3005
R9881 GND.n3068 GND.n3067 9.3005
R9882 GND.n3072 GND.n3071 9.3005
R9883 GND.n3073 GND.n3065 9.3005
R9884 GND.n4773 GND.n3074 9.3005
R9885 GND.n4772 GND.n3075 9.3005
R9886 GND.n4771 GND.n3076 9.3005
R9887 GND.n3110 GND.n3077 9.3005
R9888 GND.n3113 GND.n3112 9.3005
R9889 GND.n3114 GND.n3109 9.3005
R9890 GND.n4753 GND.n3115 9.3005
R9891 GND.n4752 GND.n3116 9.3005
R9892 GND.n4751 GND.n3117 9.3005
R9893 GND.n3153 GND.n3118 9.3005
R9894 GND.n3156 GND.n3155 9.3005
R9895 GND.n3157 GND.n3152 9.3005
R9896 GND.n4732 GND.n3158 9.3005
R9897 GND.n4731 GND.n3159 9.3005
R9898 GND.n4730 GND.n3160 9.3005
R9899 GND.n3177 GND.n3161 9.3005
R9900 GND.n4718 GND.n3178 9.3005
R9901 GND.n4717 GND.n3179 9.3005
R9902 GND.n4716 GND.n3180 9.3005
R9903 GND.n3197 GND.n3181 9.3005
R9904 GND.n4704 GND.n3198 9.3005
R9905 GND.n4703 GND.n3199 9.3005
R9906 GND.n4702 GND.n3200 9.3005
R9907 GND.n3770 GND.n3201 9.3005
R9908 GND.n3014 GND.n3013 9.3005
R9909 GND.n1593 GND.n1592 9.3005
R9910 GND.n5423 GND.n5422 9.3005
R9911 GND.n5424 GND.n1591 9.3005
R9912 GND.n5426 GND.n5425 9.3005
R9913 GND.n1587 GND.n1586 9.3005
R9914 GND.n5433 GND.n5432 9.3005
R9915 GND.n5434 GND.n1585 9.3005
R9916 GND.n5436 GND.n5435 9.3005
R9917 GND.n1581 GND.n1580 9.3005
R9918 GND.n5443 GND.n5442 9.3005
R9919 GND.n5444 GND.n1579 9.3005
R9920 GND.n5446 GND.n5445 9.3005
R9921 GND.n1575 GND.n1574 9.3005
R9922 GND.n5453 GND.n5452 9.3005
R9923 GND.n5454 GND.n1573 9.3005
R9924 GND.n5456 GND.n5455 9.3005
R9925 GND.n1569 GND.n1568 9.3005
R9926 GND.n5463 GND.n5462 9.3005
R9927 GND.n5464 GND.n1567 9.3005
R9928 GND.n5466 GND.n5465 9.3005
R9929 GND.n1563 GND.n1562 9.3005
R9930 GND.n5473 GND.n5472 9.3005
R9931 GND.n5474 GND.n1561 9.3005
R9932 GND.n5476 GND.n5475 9.3005
R9933 GND.n1557 GND.n1556 9.3005
R9934 GND.n5483 GND.n5482 9.3005
R9935 GND.n5484 GND.n1555 9.3005
R9936 GND.n5486 GND.n5485 9.3005
R9937 GND.n1551 GND.n1550 9.3005
R9938 GND.n5493 GND.n5492 9.3005
R9939 GND.n5494 GND.n1549 9.3005
R9940 GND.n5496 GND.n5495 9.3005
R9941 GND.n1545 GND.n1544 9.3005
R9942 GND.n5503 GND.n5502 9.3005
R9943 GND.n5504 GND.n1543 9.3005
R9944 GND.n5506 GND.n5505 9.3005
R9945 GND.n1539 GND.n1538 9.3005
R9946 GND.n5513 GND.n5512 9.3005
R9947 GND.n5514 GND.n1537 9.3005
R9948 GND.n5516 GND.n5515 9.3005
R9949 GND.n1533 GND.n1532 9.3005
R9950 GND.n5523 GND.n5522 9.3005
R9951 GND.n5524 GND.n1531 9.3005
R9952 GND.n5526 GND.n5525 9.3005
R9953 GND.n1527 GND.n1526 9.3005
R9954 GND.n5533 GND.n5532 9.3005
R9955 GND.n5534 GND.n1525 9.3005
R9956 GND.n5536 GND.n5535 9.3005
R9957 GND.n1521 GND.n1520 9.3005
R9958 GND.n5543 GND.n5542 9.3005
R9959 GND.n5544 GND.n1519 9.3005
R9960 GND.n5546 GND.n5545 9.3005
R9961 GND.n1515 GND.n1514 9.3005
R9962 GND.n5553 GND.n5552 9.3005
R9963 GND.n5554 GND.n1513 9.3005
R9964 GND.n5556 GND.n5555 9.3005
R9965 GND.n1509 GND.n1508 9.3005
R9966 GND.n5563 GND.n5562 9.3005
R9967 GND.n5564 GND.n1507 9.3005
R9968 GND.n5566 GND.n5565 9.3005
R9969 GND.n1503 GND.n1502 9.3005
R9970 GND.n5573 GND.n5572 9.3005
R9971 GND.n5574 GND.n1501 9.3005
R9972 GND.n5576 GND.n5575 9.3005
R9973 GND.n1497 GND.n1496 9.3005
R9974 GND.n5583 GND.n5582 9.3005
R9975 GND.n5584 GND.n1495 9.3005
R9976 GND.n5586 GND.n5585 9.3005
R9977 GND.n1491 GND.n1490 9.3005
R9978 GND.n5593 GND.n5592 9.3005
R9979 GND.n5594 GND.n1489 9.3005
R9980 GND.n5596 GND.n5595 9.3005
R9981 GND.n1485 GND.n1484 9.3005
R9982 GND.n5603 GND.n5602 9.3005
R9983 GND.n5604 GND.n1483 9.3005
R9984 GND.n5606 GND.n5605 9.3005
R9985 GND.n1479 GND.n1478 9.3005
R9986 GND.n5613 GND.n5612 9.3005
R9987 GND.n5614 GND.n1477 9.3005
R9988 GND.n5616 GND.n5615 9.3005
R9989 GND.n1473 GND.n1472 9.3005
R9990 GND.n5623 GND.n5622 9.3005
R9991 GND.n5624 GND.n1471 9.3005
R9992 GND.n5626 GND.n5625 9.3005
R9993 GND.n1467 GND.n1466 9.3005
R9994 GND.n5633 GND.n5632 9.3005
R9995 GND.n5634 GND.n1465 9.3005
R9996 GND.n5636 GND.n5635 9.3005
R9997 GND.n1461 GND.n1460 9.3005
R9998 GND.n5643 GND.n5642 9.3005
R9999 GND.n5644 GND.n1459 9.3005
R10000 GND.n5646 GND.n5645 9.3005
R10001 GND.n1455 GND.n1454 9.3005
R10002 GND.n5653 GND.n5652 9.3005
R10003 GND.n5654 GND.n1453 9.3005
R10004 GND.n5656 GND.n5655 9.3005
R10005 GND.n1449 GND.n1448 9.3005
R10006 GND.n5663 GND.n5662 9.3005
R10007 GND.n5664 GND.n1447 9.3005
R10008 GND.n5666 GND.n5665 9.3005
R10009 GND.n1443 GND.n1442 9.3005
R10010 GND.n5673 GND.n5672 9.3005
R10011 GND.n5674 GND.n1441 9.3005
R10012 GND.n5676 GND.n5675 9.3005
R10013 GND.n1437 GND.n1436 9.3005
R10014 GND.n5683 GND.n5682 9.3005
R10015 GND.n5684 GND.n1435 9.3005
R10016 GND.n5686 GND.n5685 9.3005
R10017 GND.n1431 GND.n1430 9.3005
R10018 GND.n5693 GND.n5692 9.3005
R10019 GND.n5694 GND.n1429 9.3005
R10020 GND.n5696 GND.n5695 9.3005
R10021 GND.n1425 GND.n1424 9.3005
R10022 GND.n5703 GND.n5702 9.3005
R10023 GND.n5704 GND.n1423 9.3005
R10024 GND.n5706 GND.n5705 9.3005
R10025 GND.n1419 GND.n1418 9.3005
R10026 GND.n5713 GND.n5712 9.3005
R10027 GND.n5714 GND.n1417 9.3005
R10028 GND.n5716 GND.n5715 9.3005
R10029 GND.n1413 GND.n1412 9.3005
R10030 GND.n5723 GND.n5722 9.3005
R10031 GND.n5724 GND.n1411 9.3005
R10032 GND.n5726 GND.n5725 9.3005
R10033 GND.n1407 GND.n1406 9.3005
R10034 GND.n5733 GND.n5732 9.3005
R10035 GND.n5734 GND.n1405 9.3005
R10036 GND.n5736 GND.n5735 9.3005
R10037 GND.n1401 GND.n1400 9.3005
R10038 GND.n5743 GND.n5742 9.3005
R10039 GND.n5744 GND.n1399 9.3005
R10040 GND.n5746 GND.n5745 9.3005
R10041 GND.n1395 GND.n1394 9.3005
R10042 GND.n5753 GND.n5752 9.3005
R10043 GND.n5754 GND.n1393 9.3005
R10044 GND.n5756 GND.n5755 9.3005
R10045 GND.n1389 GND.n1388 9.3005
R10046 GND.n5763 GND.n5762 9.3005
R10047 GND.n5764 GND.n1387 9.3005
R10048 GND.n5766 GND.n5765 9.3005
R10049 GND.n1383 GND.n1382 9.3005
R10050 GND.n5773 GND.n5772 9.3005
R10051 GND.n5774 GND.n1381 9.3005
R10052 GND.n5776 GND.n5775 9.3005
R10053 GND.n1377 GND.n1376 9.3005
R10054 GND.n5783 GND.n5782 9.3005
R10055 GND.n5784 GND.n1375 9.3005
R10056 GND.n5786 GND.n5785 9.3005
R10057 GND.n1371 GND.n1370 9.3005
R10058 GND.n5793 GND.n5792 9.3005
R10059 GND.n5794 GND.n1369 9.3005
R10060 GND.n5796 GND.n5795 9.3005
R10061 GND.n1365 GND.n1364 9.3005
R10062 GND.n5803 GND.n5802 9.3005
R10063 GND.n5804 GND.n1363 9.3005
R10064 GND.n5806 GND.n5805 9.3005
R10065 GND.n1359 GND.n1358 9.3005
R10066 GND.n5813 GND.n5812 9.3005
R10067 GND.n5814 GND.n1357 9.3005
R10068 GND.n5816 GND.n5815 9.3005
R10069 GND.n1353 GND.n1352 9.3005
R10070 GND.n5823 GND.n5822 9.3005
R10071 GND.n5824 GND.n1351 9.3005
R10072 GND.n5826 GND.n5825 9.3005
R10073 GND.n1347 GND.n1346 9.3005
R10074 GND.n5833 GND.n5832 9.3005
R10075 GND.n5834 GND.n1345 9.3005
R10076 GND.n5836 GND.n5835 9.3005
R10077 GND.n1341 GND.n1340 9.3005
R10078 GND.n5843 GND.n5842 9.3005
R10079 GND.n5844 GND.n1339 9.3005
R10080 GND.n5846 GND.n5845 9.3005
R10081 GND.n1335 GND.n1334 9.3005
R10082 GND.n5853 GND.n5852 9.3005
R10083 GND.n5854 GND.n1333 9.3005
R10084 GND.n5856 GND.n5855 9.3005
R10085 GND.n1329 GND.n1328 9.3005
R10086 GND.n5863 GND.n5862 9.3005
R10087 GND.n5864 GND.n1327 9.3005
R10088 GND.n5866 GND.n5865 9.3005
R10089 GND.n1323 GND.n1322 9.3005
R10090 GND.n5873 GND.n5872 9.3005
R10091 GND.n5874 GND.n1321 9.3005
R10092 GND.n5876 GND.n5875 9.3005
R10093 GND.n1317 GND.n1316 9.3005
R10094 GND.n5883 GND.n5882 9.3005
R10095 GND.n5884 GND.n1315 9.3005
R10096 GND.n5886 GND.n5885 9.3005
R10097 GND.n1311 GND.n1310 9.3005
R10098 GND.n5893 GND.n5892 9.3005
R10099 GND.n5894 GND.n1309 9.3005
R10100 GND.n5896 GND.n5895 9.3005
R10101 GND.n1305 GND.n1304 9.3005
R10102 GND.n5903 GND.n5902 9.3005
R10103 GND.n5904 GND.n1303 9.3005
R10104 GND.n5906 GND.n5905 9.3005
R10105 GND.n1299 GND.n1298 9.3005
R10106 GND.n5913 GND.n5912 9.3005
R10107 GND.n5914 GND.n1297 9.3005
R10108 GND.n5916 GND.n5915 9.3005
R10109 GND.n1293 GND.n1292 9.3005
R10110 GND.n5923 GND.n5922 9.3005
R10111 GND.n5924 GND.n1291 9.3005
R10112 GND.n5926 GND.n5925 9.3005
R10113 GND.n1287 GND.n1286 9.3005
R10114 GND.n5933 GND.n5932 9.3005
R10115 GND.n5934 GND.n1285 9.3005
R10116 GND.n5936 GND.n5935 9.3005
R10117 GND.n1281 GND.n1280 9.3005
R10118 GND.n5943 GND.n5942 9.3005
R10119 GND.n5944 GND.n1279 9.3005
R10120 GND.n5946 GND.n5945 9.3005
R10121 GND.n1275 GND.n1274 9.3005
R10122 GND.n5953 GND.n5952 9.3005
R10123 GND.n5954 GND.n1273 9.3005
R10124 GND.n5956 GND.n5955 9.3005
R10125 GND.n1269 GND.n1268 9.3005
R10126 GND.n5963 GND.n5962 9.3005
R10127 GND.n5964 GND.n1267 9.3005
R10128 GND.n5966 GND.n5965 9.3005
R10129 GND.n1263 GND.n1262 9.3005
R10130 GND.n5973 GND.n5972 9.3005
R10131 GND.n5974 GND.n1261 9.3005
R10132 GND.n5976 GND.n5975 9.3005
R10133 GND.n1257 GND.n1256 9.3005
R10134 GND.n5983 GND.n5982 9.3005
R10135 GND.n5984 GND.n1255 9.3005
R10136 GND.n5986 GND.n5985 9.3005
R10137 GND.n1251 GND.n1250 9.3005
R10138 GND.n5993 GND.n5992 9.3005
R10139 GND.n5994 GND.n1249 9.3005
R10140 GND.n5996 GND.n5995 9.3005
R10141 GND.n1245 GND.n1244 9.3005
R10142 GND.n6003 GND.n6002 9.3005
R10143 GND.n6004 GND.n1243 9.3005
R10144 GND.n6006 GND.n6005 9.3005
R10145 GND.n1239 GND.n1238 9.3005
R10146 GND.n6013 GND.n6012 9.3005
R10147 GND.n6014 GND.n1237 9.3005
R10148 GND.n6016 GND.n6015 9.3005
R10149 GND.n1233 GND.n1232 9.3005
R10150 GND.n6023 GND.n6022 9.3005
R10151 GND.n6024 GND.n1231 9.3005
R10152 GND.n6026 GND.n6025 9.3005
R10153 GND.n1227 GND.n1226 9.3005
R10154 GND.n6033 GND.n6032 9.3005
R10155 GND.n6034 GND.n1225 9.3005
R10156 GND.n6036 GND.n6035 9.3005
R10157 GND.n1221 GND.n1220 9.3005
R10158 GND.n6043 GND.n6042 9.3005
R10159 GND.n6044 GND.n1219 9.3005
R10160 GND.n6046 GND.n6045 9.3005
R10161 GND.n1215 GND.n1214 9.3005
R10162 GND.n6053 GND.n6052 9.3005
R10163 GND.n6054 GND.n1213 9.3005
R10164 GND.n6056 GND.n6055 9.3005
R10165 GND.n1209 GND.n1208 9.3005
R10166 GND.n6063 GND.n6062 9.3005
R10167 GND.n6064 GND.n1207 9.3005
R10168 GND.n6066 GND.n6065 9.3005
R10169 GND.n1203 GND.n1202 9.3005
R10170 GND.n6073 GND.n6072 9.3005
R10171 GND.n6074 GND.n1201 9.3005
R10172 GND.n6076 GND.n6075 9.3005
R10173 GND.n1197 GND.n1196 9.3005
R10174 GND.n6083 GND.n6082 9.3005
R10175 GND.n6084 GND.n1195 9.3005
R10176 GND.n6086 GND.n6085 9.3005
R10177 GND.n1191 GND.n1190 9.3005
R10178 GND.n6093 GND.n6092 9.3005
R10179 GND.n6094 GND.n1189 9.3005
R10180 GND.n6096 GND.n6095 9.3005
R10181 GND.n1185 GND.n1184 9.3005
R10182 GND.n6103 GND.n6102 9.3005
R10183 GND.n6104 GND.n1183 9.3005
R10184 GND.n6106 GND.n6105 9.3005
R10185 GND.n1179 GND.n1178 9.3005
R10186 GND.n6113 GND.n6112 9.3005
R10187 GND.n6114 GND.n1177 9.3005
R10188 GND.n6116 GND.n6115 9.3005
R10189 GND.n1173 GND.n1172 9.3005
R10190 GND.n6123 GND.n6122 9.3005
R10191 GND.n6124 GND.n1171 9.3005
R10192 GND.n6126 GND.n6125 9.3005
R10193 GND.n1167 GND.n1166 9.3005
R10194 GND.n6133 GND.n6132 9.3005
R10195 GND.n6134 GND.n1165 9.3005
R10196 GND.n6136 GND.n6135 9.3005
R10197 GND.n1161 GND.n1160 9.3005
R10198 GND.n6143 GND.n6142 9.3005
R10199 GND.n6144 GND.n1159 9.3005
R10200 GND.n6146 GND.n6145 9.3005
R10201 GND.n1155 GND.n1154 9.3005
R10202 GND.n6153 GND.n6152 9.3005
R10203 GND.n6154 GND.n1153 9.3005
R10204 GND.n6156 GND.n6155 9.3005
R10205 GND.n1149 GND.n1148 9.3005
R10206 GND.n6163 GND.n6162 9.3005
R10207 GND.n6164 GND.n1147 9.3005
R10208 GND.n6166 GND.n6165 9.3005
R10209 GND.n1143 GND.n1142 9.3005
R10210 GND.n6173 GND.n6172 9.3005
R10211 GND.n6174 GND.n1141 9.3005
R10212 GND.n6176 GND.n6175 9.3005
R10213 GND.n1137 GND.n1136 9.3005
R10214 GND.n6183 GND.n6182 9.3005
R10215 GND.n6184 GND.n1135 9.3005
R10216 GND.n6186 GND.n6185 9.3005
R10217 GND.n1131 GND.n1130 9.3005
R10218 GND.n6193 GND.n6192 9.3005
R10219 GND.n6194 GND.n1129 9.3005
R10220 GND.n6196 GND.n6195 9.3005
R10221 GND.n1125 GND.n1124 9.3005
R10222 GND.n6203 GND.n6202 9.3005
R10223 GND.n6204 GND.n1123 9.3005
R10224 GND.n6206 GND.n6205 9.3005
R10225 GND.n1119 GND.n1118 9.3005
R10226 GND.n6213 GND.n6212 9.3005
R10227 GND.n6214 GND.n1117 9.3005
R10228 GND.n6216 GND.n6215 9.3005
R10229 GND.n1113 GND.n1112 9.3005
R10230 GND.n6223 GND.n6222 9.3005
R10231 GND.n6224 GND.n1111 9.3005
R10232 GND.n6226 GND.n6225 9.3005
R10233 GND.n1107 GND.n1106 9.3005
R10234 GND.n6233 GND.n6232 9.3005
R10235 GND.n6234 GND.n1105 9.3005
R10236 GND.n6236 GND.n6235 9.3005
R10237 GND.n1101 GND.n1100 9.3005
R10238 GND.n6243 GND.n6242 9.3005
R10239 GND.n6244 GND.n1099 9.3005
R10240 GND.n6246 GND.n6245 9.3005
R10241 GND.n1095 GND.n1094 9.3005
R10242 GND.n6253 GND.n6252 9.3005
R10243 GND.n6254 GND.n1093 9.3005
R10244 GND.n6256 GND.n6255 9.3005
R10245 GND.n1089 GND.n1088 9.3005
R10246 GND.n6263 GND.n6262 9.3005
R10247 GND.n6264 GND.n1087 9.3005
R10248 GND.n6266 GND.n6265 9.3005
R10249 GND.n1083 GND.n1082 9.3005
R10250 GND.n6273 GND.n6272 9.3005
R10251 GND.n6274 GND.n1081 9.3005
R10252 GND.n6276 GND.n6275 9.3005
R10253 GND.n1077 GND.n1076 9.3005
R10254 GND.n6283 GND.n6282 9.3005
R10255 GND.n6284 GND.n1075 9.3005
R10256 GND.n6286 GND.n6285 9.3005
R10257 GND.n6293 GND.n6292 9.3005
R10258 GND.n6294 GND.n1069 9.3005
R10259 GND.n6296 GND.n6295 9.3005
R10260 GND.n1065 GND.n1064 9.3005
R10261 GND.n6303 GND.n6302 9.3005
R10262 GND.n6304 GND.n1063 9.3005
R10263 GND.n6306 GND.n6305 9.3005
R10264 GND.n1059 GND.n1058 9.3005
R10265 GND.n6313 GND.n6312 9.3005
R10266 GND.n6314 GND.n1057 9.3005
R10267 GND.n6316 GND.n6315 9.3005
R10268 GND.n1053 GND.n1052 9.3005
R10269 GND.n6323 GND.n6322 9.3005
R10270 GND.n6324 GND.n1051 9.3005
R10271 GND.n6326 GND.n6325 9.3005
R10272 GND.n1047 GND.n1046 9.3005
R10273 GND.n6333 GND.n6332 9.3005
R10274 GND.n6334 GND.n1045 9.3005
R10275 GND.n6336 GND.n6335 9.3005
R10276 GND.n1041 GND.n1040 9.3005
R10277 GND.n6343 GND.n6342 9.3005
R10278 GND.n6344 GND.n1039 9.3005
R10279 GND.n6346 GND.n6345 9.3005
R10280 GND.n1035 GND.n1034 9.3005
R10281 GND.n6353 GND.n6352 9.3005
R10282 GND.n6354 GND.n1033 9.3005
R10283 GND.n6356 GND.n6355 9.3005
R10284 GND.n1029 GND.n1028 9.3005
R10285 GND.n6363 GND.n6362 9.3005
R10286 GND.n6364 GND.n1027 9.3005
R10287 GND.n6366 GND.n6365 9.3005
R10288 GND.n1023 GND.n1022 9.3005
R10289 GND.n6373 GND.n6372 9.3005
R10290 GND.n6374 GND.n1021 9.3005
R10291 GND.n6376 GND.n6375 9.3005
R10292 GND.n1017 GND.n1016 9.3005
R10293 GND.n6383 GND.n6382 9.3005
R10294 GND.n6384 GND.n1015 9.3005
R10295 GND.n6386 GND.n6385 9.3005
R10296 GND.n1011 GND.n1010 9.3005
R10297 GND.n6393 GND.n6392 9.3005
R10298 GND.n6394 GND.n1009 9.3005
R10299 GND.n6396 GND.n6395 9.3005
R10300 GND.n1005 GND.n1004 9.3005
R10301 GND.n6403 GND.n6402 9.3005
R10302 GND.n1071 GND.n1070 9.3005
R10303 GND.n523 GND.n522 9.3005
R10304 GND.n508 GND.n507 9.3005
R10305 GND.n517 GND.n516 9.3005
R10306 GND.n515 GND.n514 9.3005
R10307 GND.n500 GND.n499 9.3005
R10308 GND.n485 GND.n484 9.3005
R10309 GND.n494 GND.n493 9.3005
R10310 GND.n492 GND.n491 9.3005
R10311 GND.n479 GND.n478 9.3005
R10312 GND.n464 GND.n463 9.3005
R10313 GND.n473 GND.n472 9.3005
R10314 GND.n471 GND.n470 9.3005
R10315 GND.n456 GND.n455 9.3005
R10316 GND.n441 GND.n440 9.3005
R10317 GND.n450 GND.n449 9.3005
R10318 GND.n448 GND.n447 9.3005
R10319 GND.n435 GND.n434 9.3005
R10320 GND.n420 GND.n419 9.3005
R10321 GND.n429 GND.n428 9.3005
R10322 GND.n427 GND.n426 9.3005
R10323 GND.n412 GND.n411 9.3005
R10324 GND.n397 GND.n396 9.3005
R10325 GND.n406 GND.n405 9.3005
R10326 GND.n404 GND.n403 9.3005
R10327 GND.n391 GND.n390 9.3005
R10328 GND.n376 GND.n375 9.3005
R10329 GND.n385 GND.n384 9.3005
R10330 GND.n383 GND.n382 9.3005
R10331 GND.n368 GND.n367 9.3005
R10332 GND.n353 GND.n352 9.3005
R10333 GND.n362 GND.n361 9.3005
R10334 GND.n360 GND.n359 9.3005
R10335 GND.n347 GND.n346 9.3005
R10336 GND.n332 GND.n331 9.3005
R10337 GND.n341 GND.n340 9.3005
R10338 GND.n339 GND.n338 9.3005
R10339 GND.n324 GND.n323 9.3005
R10340 GND.n309 GND.n308 9.3005
R10341 GND.n318 GND.n317 9.3005
R10342 GND.n316 GND.n315 9.3005
R10343 GND.n304 GND.n303 9.3005
R10344 GND.n289 GND.n288 9.3005
R10345 GND.n298 GND.n297 9.3005
R10346 GND.n296 GND.n295 9.3005
R10347 GND.n281 GND.n280 9.3005
R10348 GND.n266 GND.n265 9.3005
R10349 GND.n275 GND.n274 9.3005
R10350 GND.n273 GND.n272 9.3005
R10351 GND.n4249 GND.n4248 9.3005
R10352 GND.n4250 GND.n4239 9.3005
R10353 GND.n4253 GND.n4238 9.3005
R10354 GND.n4254 GND.n4237 9.3005
R10355 GND.n4257 GND.n4236 9.3005
R10356 GND.n4258 GND.n4235 9.3005
R10357 GND.n4261 GND.n4234 9.3005
R10358 GND.n4262 GND.n4233 9.3005
R10359 GND.n4265 GND.n4232 9.3005
R10360 GND.n4268 GND.n4267 9.3005
R10361 GND.n4247 GND.n4244 9.3005
R10362 GND.n4246 GND.n4245 9.3005
R10363 GND.n4277 GND.n4102 9.3005
R10364 GND.n4279 GND.n4278 9.3005
R10365 GND.n4280 GND.n4101 9.3005
R10366 GND.n4284 GND.n4281 9.3005
R10367 GND.n4285 GND.n4100 9.3005
R10368 GND.n4303 GND.n4302 9.3005
R10369 GND.n4304 GND.n4099 9.3005
R10370 GND.n4306 GND.n4305 9.3005
R10371 GND.n4097 GND.n4096 9.3005
R10372 GND.n4318 GND.n4317 9.3005
R10373 GND.n4319 GND.n4095 9.3005
R10374 GND.n4321 GND.n4320 9.3005
R10375 GND.n4093 GND.n4092 9.3005
R10376 GND.n4333 GND.n4332 9.3005
R10377 GND.n4334 GND.n4091 9.3005
R10378 GND.n4347 GND.n4335 9.3005
R10379 GND.n4346 GND.n4336 9.3005
R10380 GND.n4345 GND.n4337 9.3005
R10381 GND.n4344 GND.n4338 9.3005
R10382 GND.n4342 GND.n4339 9.3005
R10383 GND.n4341 GND.n4340 9.3005
R10384 GND.n529 GND.n527 9.3005
R10385 GND.n4276 GND.n4103 9.3005
R10386 GND.n6858 GND.n6857 9.3005
R10387 GND.n530 GND.n528 9.3005
R10388 GND.n4450 GND.n4407 9.3005
R10389 GND.n4449 GND.n4408 9.3005
R10390 GND.n4448 GND.n4409 9.3005
R10391 GND.n4414 GND.n4410 9.3005
R10392 GND.n4438 GND.n4415 9.3005
R10393 GND.n4437 GND.n4416 9.3005
R10394 GND.n4436 GND.n4417 9.3005
R10395 GND.n4420 GND.n4418 9.3005
R10396 GND.n4426 GND.n4421 9.3005
R10397 GND.n4425 GND.n4422 9.3005
R10398 GND.n4424 GND.n4423 9.3005
R10399 GND.n793 GND.n792 9.3005
R10400 GND.n6621 GND.n6620 9.3005
R10401 GND.n6622 GND.n791 9.3005
R10402 GND.n6624 GND.n6623 9.3005
R10403 GND.n788 GND.n787 9.3005
R10404 GND.n6635 GND.n6634 9.3005
R10405 GND.n6636 GND.n786 9.3005
R10406 GND.n6639 GND.n6638 9.3005
R10407 GND.n6637 GND.n783 9.3005
R10408 GND.n6650 GND.n782 9.3005
R10409 GND.n6652 GND.n6651 9.3005
R10410 GND.n6671 GND.n760 9.3005
R10411 GND.n6670 GND.n763 9.3005
R10412 GND.n767 GND.n764 9.3005
R10413 GND.n768 GND.n765 9.3005
R10414 GND.n6663 GND.n769 9.3005
R10415 GND.n6662 GND.n770 9.3005
R10416 GND.n6661 GND.n771 9.3005
R10417 GND.n775 GND.n772 9.3005
R10418 GND.n6656 GND.n776 9.3005
R10419 GND.n6655 GND.n6654 9.3005
R10420 GND.n6653 GND.n779 9.3005
R10421 GND.n6673 GND.n6672 9.3005
R10422 GND.n6787 GND.n650 9.3005
R10423 GND.n6786 GND.n652 9.3005
R10424 GND.n657 GND.n653 9.3005
R10425 GND.n6781 GND.n658 9.3005
R10426 GND.n6780 GND.n659 9.3005
R10427 GND.n6779 GND.n660 9.3005
R10428 GND.n664 GND.n661 9.3005
R10429 GND.n6774 GND.n665 9.3005
R10430 GND.n6773 GND.n666 9.3005
R10431 GND.n6772 GND.n6771 9.3005
R10432 GND.n6770 GND.n667 9.3005
R10433 GND.n6769 GND.n6768 9.3005
R10434 GND.n673 GND.n672 9.3005
R10435 GND.n6763 GND.n677 9.3005
R10436 GND.n6762 GND.n678 9.3005
R10437 GND.n6761 GND.n679 9.3005
R10438 GND.n683 GND.n680 9.3005
R10439 GND.n6756 GND.n684 9.3005
R10440 GND.n6755 GND.n685 9.3005
R10441 GND.n6754 GND.n686 9.3005
R10442 GND.n693 GND.n687 9.3005
R10443 GND.n6749 GND.n6748 9.3005
R10444 GND.n6747 GND.n690 9.3005
R10445 GND.n6746 GND.n6745 9.3005
R10446 GND.n695 GND.n694 9.3005
R10447 GND.n6740 GND.n698 9.3005
R10448 GND.n6739 GND.n699 9.3005
R10449 GND.n6738 GND.n700 9.3005
R10450 GND.n704 GND.n701 9.3005
R10451 GND.n6733 GND.n705 9.3005
R10452 GND.n6732 GND.n706 9.3005
R10453 GND.n6731 GND.n707 9.3005
R10454 GND.n711 GND.n708 9.3005
R10455 GND.n6726 GND.n712 9.3005
R10456 GND.n6722 GND.n713 9.3005
R10457 GND.n6721 GND.n714 9.3005
R10458 GND.n718 GND.n715 9.3005
R10459 GND.n6716 GND.n719 9.3005
R10460 GND.n6715 GND.n720 9.3005
R10461 GND.n6714 GND.n721 9.3005
R10462 GND.n725 GND.n722 9.3005
R10463 GND.n6709 GND.n726 9.3005
R10464 GND.n6708 GND.n727 9.3005
R10465 GND.n6707 GND.n728 9.3005
R10466 GND.n732 GND.n729 9.3005
R10467 GND.n6702 GND.n733 9.3005
R10468 GND.n6698 GND.n734 9.3005
R10469 GND.n6697 GND.n735 9.3005
R10470 GND.n739 GND.n736 9.3005
R10471 GND.n6692 GND.n740 9.3005
R10472 GND.n6691 GND.n741 9.3005
R10473 GND.n6690 GND.n742 9.3005
R10474 GND.n746 GND.n743 9.3005
R10475 GND.n6685 GND.n747 9.3005
R10476 GND.n6684 GND.n748 9.3005
R10477 GND.n6683 GND.n749 9.3005
R10478 GND.n753 GND.n750 9.3005
R10479 GND.n6678 GND.n754 9.3005
R10480 GND.n6677 GND.n6676 9.3005
R10481 GND.n6675 GND.n757 9.3005
R10482 GND.n6789 GND.n6788 9.3005
R10483 GND.n4542 GND.n4541 9.3005
R10484 GND.n3939 GND.n3937 9.3005
R10485 GND.n4291 GND.n4290 9.3005
R10486 GND.n4294 GND.n4289 9.3005
R10487 GND.n4296 GND.n4295 9.3005
R10488 GND.n4297 GND.n3978 9.3005
R10489 GND.n4521 GND.n3979 9.3005
R10490 GND.n4520 GND.n3980 9.3005
R10491 GND.n4519 GND.n3981 9.3005
R10492 GND.n4312 GND.n3982 9.3005
R10493 GND.n4509 GND.n4000 9.3005
R10494 GND.n4508 GND.n4001 9.3005
R10495 GND.n4507 GND.n4002 9.3005
R10496 GND.n4327 GND.n4003 9.3005
R10497 GND.n4497 GND.n4021 9.3005
R10498 GND.n4496 GND.n4022 9.3005
R10499 GND.n4495 GND.n4023 9.3005
R10500 GND.n4354 GND.n4024 9.3005
R10501 GND.n4355 GND.n4049 9.3005
R10502 GND.n4472 GND.n4050 9.3005
R10503 GND.n4471 GND.n4051 9.3005
R10504 GND.n4470 GND.n4052 9.3005
R10505 GND.n4360 GND.n4053 9.3005
R10506 GND.n4460 GND.n4361 9.3005
R10507 GND.n4459 GND.n4366 9.3005
R10508 GND.n4458 GND.n4367 9.3005
R10509 GND.n4412 GND.n557 9.3005
R10510 GND.n6845 GND.n558 9.3005
R10511 GND.n6844 GND.n559 9.3005
R10512 GND.n6843 GND.n560 9.3005
R10513 GND.n4419 GND.n561 9.3005
R10514 GND.n6833 GND.n578 9.3005
R10515 GND.n6832 GND.n579 9.3005
R10516 GND.n6831 GND.n580 9.3005
R10517 GND.n795 GND.n581 9.3005
R10518 GND.n6821 GND.n598 9.3005
R10519 GND.n6820 GND.n599 9.3005
R10520 GND.n6819 GND.n600 9.3005
R10521 GND.n790 GND.n601 9.3005
R10522 GND.n6809 GND.n619 9.3005
R10523 GND.n6808 GND.n620 9.3005
R10524 GND.n6807 GND.n621 9.3005
R10525 GND.n785 GND.n622 9.3005
R10526 GND.n6797 GND.n640 9.3005
R10527 GND.n6796 GND.n641 9.3005
R10528 GND.n6795 GND.n642 9.3005
R10529 GND.n3938 GND.n3936 9.3005
R10530 GND.n4541 GND.n4540 9.3005
R10531 GND.n4539 GND.n3939 9.3005
R10532 GND.n4290 GND.n3941 9.3005
R10533 GND.n4289 GND.n4288 9.3005
R10534 GND.n4296 GND.n4286 9.3005
R10535 GND.n4298 GND.n4297 9.3005
R10536 GND.n4098 GND.n3979 9.3005
R10537 GND.n4310 GND.n3980 9.3005
R10538 GND.n4311 GND.n3981 9.3005
R10539 GND.n4313 GND.n4312 9.3005
R10540 GND.n4094 GND.n4000 9.3005
R10541 GND.n4325 GND.n4001 9.3005
R10542 GND.n4326 GND.n4002 9.3005
R10543 GND.n4328 GND.n4327 9.3005
R10544 GND.n4054 GND.n4021 9.3005
R10545 GND.n4351 GND.n4022 9.3005
R10546 GND.n4352 GND.n4023 9.3005
R10547 GND.n4354 GND.n4353 9.3005
R10548 GND.n4357 GND.n4355 9.3005
R10549 GND.n4358 GND.n4050 9.3005
R10550 GND.n4359 GND.n4051 9.3005
R10551 GND.n4466 GND.n4052 9.3005
R10552 GND.n4465 GND.n4360 9.3005
R10553 GND.n4464 GND.n4361 9.3005
R10554 GND.n4366 GND.n4362 9.3005
R10555 GND.n4411 GND.n4367 9.3005
R10556 GND.n4444 GND.n4412 9.3005
R10557 GND.n4443 GND.n558 9.3005
R10558 GND.n4442 GND.n559 9.3005
R10559 GND.n4413 GND.n560 9.3005
R10560 GND.n4432 GND.n4419 9.3005
R10561 GND.n4431 GND.n578 9.3005
R10562 GND.n4430 GND.n579 9.3005
R10563 GND.n794 GND.n580 9.3005
R10564 GND.n6614 GND.n795 9.3005
R10565 GND.n6615 GND.n598 9.3005
R10566 GND.n6616 GND.n599 9.3005
R10567 GND.n789 GND.n600 9.3005
R10568 GND.n6628 GND.n790 9.3005
R10569 GND.n6629 GND.n619 9.3005
R10570 GND.n6630 GND.n620 9.3005
R10571 GND.n784 GND.n621 9.3005
R10572 GND.n6643 GND.n785 9.3005
R10573 GND.n6644 GND.n640 9.3005
R10574 GND.n6646 GND.n641 9.3005
R10575 GND.n6645 GND.n642 9.3005
R10576 GND.n3940 GND.n3938 9.3005
R10577 GND.n4231 GND.n4138 9.3005
R10578 GND.n4230 GND.n4229 9.3005
R10579 GND.n4226 GND.n4139 9.3005
R10580 GND.n4223 GND.n4222 9.3005
R10581 GND.n4221 GND.n4140 9.3005
R10582 GND.n4220 GND.n4219 9.3005
R10583 GND.n4216 GND.n4141 9.3005
R10584 GND.n4213 GND.n4212 9.3005
R10585 GND.n4211 GND.n4142 9.3005
R10586 GND.n4210 GND.n4209 9.3005
R10587 GND.n4206 GND.n4143 9.3005
R10588 GND.n4203 GND.n4202 9.3005
R10589 GND.n4201 GND.n4144 9.3005
R10590 GND.n4200 GND.n4199 9.3005
R10591 GND.n4193 GND.n4145 9.3005
R10592 GND.n4190 GND.n4189 9.3005
R10593 GND.n4188 GND.n4146 9.3005
R10594 GND.n4187 GND.n4186 9.3005
R10595 GND.n4183 GND.n4147 9.3005
R10596 GND.n4180 GND.n4179 9.3005
R10597 GND.n4178 GND.n4148 9.3005
R10598 GND.n4177 GND.n4176 9.3005
R10599 GND.n4173 GND.n4149 9.3005
R10600 GND.n4170 GND.n4169 9.3005
R10601 GND.n4168 GND.n4150 9.3005
R10602 GND.n4167 GND.n4166 9.3005
R10603 GND.n4160 GND.n4151 9.3005
R10604 GND.n4157 GND.n4156 9.3005
R10605 GND.n4155 GND.n4153 9.3005
R10606 GND.n4154 GND.n3885 9.3005
R10607 GND.n4634 GND.n3884 9.3005
R10608 GND.n4580 GND.n3880 9.3005
R10609 GND.n4582 GND.n4581 9.3005
R10610 GND.n4585 GND.n4579 9.3005
R10611 GND.n4587 GND.n4578 9.3005
R10612 GND.n4589 GND.n4573 9.3005
R10613 GND.n4592 GND.n4572 9.3005
R10614 GND.n4593 GND.n4571 9.3005
R10615 GND.n4596 GND.n4570 9.3005
R10616 GND.n4597 GND.n4569 9.3005
R10617 GND.n4600 GND.n4568 9.3005
R10618 GND.n4601 GND.n4567 9.3005
R10619 GND.n4604 GND.n4566 9.3005
R10620 GND.n4605 GND.n4565 9.3005
R10621 GND.n4608 GND.n4564 9.3005
R10622 GND.n4610 GND.n4563 9.3005
R10623 GND.n4612 GND.n4558 9.3005
R10624 GND.n4615 GND.n4557 9.3005
R10625 GND.n4616 GND.n4556 9.3005
R10626 GND.n4619 GND.n4555 9.3005
R10627 GND.n4620 GND.n4554 9.3005
R10628 GND.n4623 GND.n4553 9.3005
R10629 GND.n4625 GND.n4552 9.3005
R10630 GND.n4626 GND.n4551 9.3005
R10631 GND.n4627 GND.n4550 9.3005
R10632 GND.n4628 GND.n4549 9.3005
R10633 GND.n4611 GND.n4560 9.3005
R10634 GND.n4588 GND.n4575 9.3005
R10635 GND.n4271 GND.n4270 9.3005
R10636 GND.n4546 GND.n3927 9.3005
R10637 GND.n3962 GND.n3928 9.3005
R10638 GND.n3965 GND.n3964 9.3005
R10639 GND.n3966 GND.n3961 9.3005
R10640 GND.n4527 GND.n3967 9.3005
R10641 GND.n4526 GND.n3968 9.3005
R10642 GND.n4525 GND.n3969 9.3005
R10643 GND.n3989 GND.n3970 9.3005
R10644 GND.n4515 GND.n3990 9.3005
R10645 GND.n4514 GND.n3991 9.3005
R10646 GND.n4513 GND.n3992 9.3005
R10647 GND.n4010 GND.n3993 9.3005
R10648 GND.n4503 GND.n4011 9.3005
R10649 GND.n4502 GND.n4012 9.3005
R10650 GND.n4501 GND.n4013 9.3005
R10651 GND.n4015 GND.n4014 9.3005
R10652 GND.n4491 GND.n542 9.3005
R10653 GND.n548 GND.n541 9.3005
R10654 GND.n6839 GND.n568 9.3005
R10655 GND.n6838 GND.n569 9.3005
R10656 GND.n6837 GND.n570 9.3005
R10657 GND.n588 GND.n571 9.3005
R10658 GND.n6827 GND.n589 9.3005
R10659 GND.n6826 GND.n590 9.3005
R10660 GND.n6825 GND.n591 9.3005
R10661 GND.n608 GND.n592 9.3005
R10662 GND.n6815 GND.n609 9.3005
R10663 GND.n6814 GND.n610 9.3005
R10664 GND.n6813 GND.n611 9.3005
R10665 GND.n629 GND.n612 9.3005
R10666 GND.n6803 GND.n630 9.3005
R10667 GND.n6802 GND.n631 9.3005
R10668 GND.n6801 GND.n632 9.3005
R10669 GND.n649 GND.n633 9.3005
R10670 GND.n6791 GND.n6790 9.3005
R10671 GND.n4548 GND.n4547 9.3005
R10672 GND.n6850 GND.n6849 9.3005
R10673 GND.n2736 GND.n2703 9.3005
R10674 GND.n2706 GND.n2704 9.3005
R10675 GND.n2730 GND.n2707 9.3005
R10676 GND.n2729 GND.n2708 9.3005
R10677 GND.n2728 GND.n2709 9.3005
R10678 GND.n2714 GND.n2710 9.3005
R10679 GND.n2724 GND.n2715 9.3005
R10680 GND.n2723 GND.n2716 9.3005
R10681 GND.n2722 GND.n2717 9.3005
R10682 GND.n2720 GND.n2719 9.3005
R10683 GND.n2718 GND.n2095 9.3005
R10684 GND.n2093 GND.n2092 9.3005
R10685 GND.n2828 GND.n2827 9.3005
R10686 GND.n2829 GND.n2091 9.3005
R10687 GND.n2834 GND.n2830 9.3005
R10688 GND.n2833 GND.n2832 9.3005
R10689 GND.n2831 GND.n2065 9.3005
R10690 GND.n2063 GND.n2062 9.3005
R10691 GND.n2914 GND.n2913 9.3005
R10692 GND.n2915 GND.n2061 9.3005
R10693 GND.n4885 GND.n2916 9.3005
R10694 GND.n4884 GND.n2917 9.3005
R10695 GND.n4883 GND.n2918 9.3005
R10696 GND.n2923 GND.n2919 9.3005
R10697 GND.n4877 GND.n2924 9.3005
R10698 GND.n4876 GND.n2925 9.3005
R10699 GND.n4875 GND.n2926 9.3005
R10700 GND.n2941 GND.n2927 9.3005
R10701 GND.n4863 GND.n2942 9.3005
R10702 GND.n4862 GND.n2943 9.3005
R10703 GND.n4861 GND.n2944 9.3005
R10704 GND.n3546 GND.n2945 9.3005
R10705 GND.n3547 GND.n3545 9.3005
R10706 GND.n3550 GND.n3549 9.3005
R10707 GND.n3548 GND.n3000 9.3005
R10708 GND.n4808 GND.n3001 9.3005
R10709 GND.n4807 GND.n3002 9.3005
R10710 GND.n4806 GND.n3003 9.3005
R10711 GND.n3041 GND.n3004 9.3005
R10712 GND.n3044 GND.n3043 9.3005
R10713 GND.n3045 GND.n3040 9.3005
R10714 GND.n4787 GND.n3046 9.3005
R10715 GND.n4786 GND.n3047 9.3005
R10716 GND.n4785 GND.n3048 9.3005
R10717 GND.n3085 GND.n3049 9.3005
R10718 GND.n3088 GND.n3087 9.3005
R10719 GND.n3089 GND.n3084 9.3005
R10720 GND.n4766 GND.n3090 9.3005
R10721 GND.n4765 GND.n3091 9.3005
R10722 GND.n4764 GND.n3092 9.3005
R10723 GND.n3135 GND.n3093 9.3005
R10724 GND.n3137 GND.n3136 9.3005
R10725 GND.n3141 GND.n3140 9.3005
R10726 GND.n3142 GND.n3134 9.3005
R10727 GND.n4739 GND.n3143 9.3005
R10728 GND.n4738 GND.n3144 9.3005
R10729 GND.n4737 GND.n3145 9.3005
R10730 GND.n3330 GND.n3146 9.3005
R10731 GND.n3332 GND.n3331 9.3005
R10732 GND.n3329 GND.n3328 9.3005
R10733 GND.n3337 GND.n3336 9.3005
R10734 GND.n3338 GND.n3327 9.3005
R10735 GND.n3340 GND.n3339 9.3005
R10736 GND.n3325 GND.n3324 9.3005
R10737 GND.n3741 GND.n3740 9.3005
R10738 GND.n3742 GND.n3323 9.3005
R10739 GND.n3747 GND.n3743 9.3005
R10740 GND.n3746 GND.n3745 9.3005
R10741 GND.n3744 GND.n3218 9.3005
R10742 GND.n4689 GND.n3219 9.3005
R10743 GND.n4688 GND.n3220 9.3005
R10744 GND.n4687 GND.n3221 9.3005
R10745 GND.n3236 GND.n3222 9.3005
R10746 GND.n4675 GND.n3237 9.3005
R10747 GND.n4674 GND.n3238 9.3005
R10748 GND.n4673 GND.n3239 9.3005
R10749 GND.n4114 GND.n3240 9.3005
R10750 GND.n4115 GND.n4113 9.3005
R10751 GND.n4119 GND.n4116 9.3005
R10752 GND.n4118 GND.n4117 9.3005
R10753 GND.n4109 GND.n4108 9.3005
R10754 GND.n4127 GND.n4126 9.3005
R10755 GND.n4128 GND.n4107 9.3005
R10756 GND.n4133 GND.n4129 9.3005
R10757 GND.n4132 GND.n4131 9.3005
R10758 GND.n4130 GND.n3947 9.3005
R10759 GND.n4534 GND.n3948 9.3005
R10760 GND.n4533 GND.n3949 9.3005
R10761 GND.n4532 GND.n3950 9.3005
R10762 GND.n4066 GND.n3951 9.3005
R10763 GND.n4067 GND.n4065 9.3005
R10764 GND.n4069 GND.n4068 9.3005
R10765 GND.n4063 GND.n4062 9.3005
R10766 GND.n4074 GND.n4073 9.3005
R10767 GND.n4075 GND.n4061 9.3005
R10768 GND.n4077 GND.n4076 9.3005
R10769 GND.n4059 GND.n4058 9.3005
R10770 GND.n4082 GND.n4081 9.3005
R10771 GND.n4083 GND.n4057 9.3005
R10772 GND.n4088 GND.n4084 9.3005
R10773 GND.n4087 GND.n4086 9.3005
R10774 GND.n4085 GND.n4036 9.3005
R10775 GND.n4401 GND.n4383 9.3005
R10776 GND.n4386 GND.n4384 9.3005
R10777 GND.n4397 GND.n4387 9.3005
R10778 GND.n4396 GND.n4388 9.3005
R10779 GND.n4395 GND.n4389 9.3005
R10780 GND.n4392 GND.n4391 9.3005
R10781 GND.n4390 GND.n799 9.3005
R10782 GND.n6609 GND.n800 9.3005
R10783 GND.n6608 GND.n801 9.3005
R10784 GND.n6607 GND.n802 9.3005
R10785 GND.n805 GND.n803 9.3005
R10786 GND.n6603 GND.n806 9.3005
R10787 GND.n6602 GND.n807 9.3005
R10788 GND.n6601 GND.n808 9.3005
R10789 GND.n811 GND.n809 9.3005
R10790 GND.n6597 GND.n812 9.3005
R10791 GND.n6596 GND.n813 9.3005
R10792 GND.n6595 GND.n814 9.3005
R10793 GND.n817 GND.n815 9.3005
R10794 GND.n6590 GND.n818 9.3005
R10795 GND.n6589 GND.n819 9.3005
R10796 GND.n6588 GND.n820 9.3005
R10797 GND.n826 GND.n821 9.3005
R10798 GND.n6582 GND.n827 9.3005
R10799 GND.n6581 GND.n828 9.3005
R10800 GND.n6580 GND.n829 9.3005
R10801 GND.n834 GND.n830 9.3005
R10802 GND.n6574 GND.n835 9.3005
R10803 GND.n6573 GND.n836 9.3005
R10804 GND.n6572 GND.n837 9.3005
R10805 GND.n842 GND.n838 9.3005
R10806 GND.n6566 GND.n843 9.3005
R10807 GND.n6565 GND.n844 9.3005
R10808 GND.n6564 GND.n845 9.3005
R10809 GND.n850 GND.n846 9.3005
R10810 GND.n6558 GND.n851 9.3005
R10811 GND.n6557 GND.n852 9.3005
R10812 GND.n6556 GND.n853 9.3005
R10813 GND.n858 GND.n854 9.3005
R10814 GND.n6550 GND.n859 9.3005
R10815 GND.n6549 GND.n860 9.3005
R10816 GND.n6548 GND.n861 9.3005
R10817 GND.n866 GND.n862 9.3005
R10818 GND.n6542 GND.n867 9.3005
R10819 GND.n6541 GND.n868 9.3005
R10820 GND.n6540 GND.n869 9.3005
R10821 GND.n874 GND.n870 9.3005
R10822 GND.n6534 GND.n875 9.3005
R10823 GND.n6533 GND.n876 9.3005
R10824 GND.n6532 GND.n877 9.3005
R10825 GND.n882 GND.n878 9.3005
R10826 GND.n6526 GND.n883 9.3005
R10827 GND.n6525 GND.n884 9.3005
R10828 GND.n6524 GND.n885 9.3005
R10829 GND.n890 GND.n886 9.3005
R10830 GND.n6518 GND.n891 9.3005
R10831 GND.n6517 GND.n892 9.3005
R10832 GND.n6516 GND.n893 9.3005
R10833 GND.n898 GND.n894 9.3005
R10834 GND.n6510 GND.n899 9.3005
R10835 GND.n6509 GND.n900 9.3005
R10836 GND.n6508 GND.n901 9.3005
R10837 GND.n906 GND.n902 9.3005
R10838 GND.n6502 GND.n907 9.3005
R10839 GND.n6501 GND.n908 9.3005
R10840 GND.n6500 GND.n909 9.3005
R10841 GND.n914 GND.n910 9.3005
R10842 GND.n6494 GND.n915 9.3005
R10843 GND.n6493 GND.n916 9.3005
R10844 GND.n6492 GND.n917 9.3005
R10845 GND.n922 GND.n918 9.3005
R10846 GND.n6486 GND.n923 9.3005
R10847 GND.n6485 GND.n924 9.3005
R10848 GND.n6484 GND.n925 9.3005
R10849 GND.n930 GND.n926 9.3005
R10850 GND.n6478 GND.n931 9.3005
R10851 GND.n6477 GND.n932 9.3005
R10852 GND.n6476 GND.n933 9.3005
R10853 GND.n938 GND.n934 9.3005
R10854 GND.n6470 GND.n939 9.3005
R10855 GND.n6469 GND.n940 9.3005
R10856 GND.n6468 GND.n941 9.3005
R10857 GND.n946 GND.n942 9.3005
R10858 GND.n6462 GND.n947 9.3005
R10859 GND.n6461 GND.n948 9.3005
R10860 GND.n6460 GND.n949 9.3005
R10861 GND.n954 GND.n950 9.3005
R10862 GND.n6454 GND.n955 9.3005
R10863 GND.n6453 GND.n956 9.3005
R10864 GND.n6452 GND.n957 9.3005
R10865 GND.n962 GND.n958 9.3005
R10866 GND.n6446 GND.n963 9.3005
R10867 GND.n6445 GND.n964 9.3005
R10868 GND.n6444 GND.n965 9.3005
R10869 GND.n970 GND.n966 9.3005
R10870 GND.n6438 GND.n971 9.3005
R10871 GND.n6437 GND.n972 9.3005
R10872 GND.n6436 GND.n973 9.3005
R10873 GND.n978 GND.n974 9.3005
R10874 GND.n6430 GND.n979 9.3005
R10875 GND.n6429 GND.n980 9.3005
R10876 GND.n6428 GND.n981 9.3005
R10877 GND.n986 GND.n982 9.3005
R10878 GND.n6422 GND.n987 9.3005
R10879 GND.n6421 GND.n988 9.3005
R10880 GND.n6420 GND.n989 9.3005
R10881 GND.n994 GND.n990 9.3005
R10882 GND.n6414 GND.n995 9.3005
R10883 GND.n6413 GND.n996 9.3005
R10884 GND.n6412 GND.n997 9.3005
R10885 GND.n1002 GND.n998 9.3005
R10886 GND.n6406 GND.n1003 9.3005
R10887 GND.n6405 GND.n6404 9.3005
R10888 GND.n2283 GND.n2280 9.3005
R10889 GND.n2497 GND.n2496 9.3005
R10890 GND.n2495 GND.n2285 9.3005
R10891 GND.n2494 GND.n2493 9.3005
R10892 GND.n2287 GND.n2286 9.3005
R10893 GND.n2487 GND.n2486 9.3005
R10894 GND.n2485 GND.n2289 9.3005
R10895 GND.n2484 GND.n2483 9.3005
R10896 GND.n2291 GND.n2290 9.3005
R10897 GND.n2477 GND.n2476 9.3005
R10898 GND.n2475 GND.n2293 9.3005
R10899 GND.n2474 GND.n2473 9.3005
R10900 GND.n2295 GND.n2294 9.3005
R10901 GND.n2467 GND.n2463 9.3005
R10902 GND.n2462 GND.n2297 9.3005
R10903 GND.n2461 GND.n2460 9.3005
R10904 GND.n2299 GND.n2298 9.3005
R10905 GND.n2454 GND.n2453 9.3005
R10906 GND.n2452 GND.n2301 9.3005
R10907 GND.n2451 GND.n2450 9.3005
R10908 GND.n2303 GND.n2302 9.3005
R10909 GND.n2444 GND.n2443 9.3005
R10910 GND.n2442 GND.n2305 9.3005
R10911 GND.n2441 GND.n2440 9.3005
R10912 GND.n2307 GND.n2306 9.3005
R10913 GND.n2434 GND.n2430 9.3005
R10914 GND.n2429 GND.n2309 9.3005
R10915 GND.n2428 GND.n2427 9.3005
R10916 GND.n2311 GND.n2310 9.3005
R10917 GND.n2421 GND.n2420 9.3005
R10918 GND.n2419 GND.n2313 9.3005
R10919 GND.n2418 GND.n2417 9.3005
R10920 GND.n2315 GND.n2314 9.3005
R10921 GND.n2411 GND.n2410 9.3005
R10922 GND.n2409 GND.n2317 9.3005
R10923 GND.n2408 GND.n2407 9.3005
R10924 GND.n2319 GND.n2318 9.3005
R10925 GND.n2397 GND.n2321 9.3005
R10926 GND.n2396 GND.n2395 9.3005
R10927 GND.n2323 GND.n2322 9.3005
R10928 GND.n2389 GND.n2388 9.3005
R10929 GND.n2387 GND.n2325 9.3005
R10930 GND.n2386 GND.n2385 9.3005
R10931 GND.n2327 GND.n2326 9.3005
R10932 GND.n2379 GND.n2378 9.3005
R10933 GND.n2377 GND.n2329 9.3005
R10934 GND.n2376 GND.n2375 9.3005
R10935 GND.n2331 GND.n2330 9.3005
R10936 GND.n2365 GND.n2333 9.3005
R10937 GND.n2364 GND.n2363 9.3005
R10938 GND.n2335 GND.n2334 9.3005
R10939 GND.n2357 GND.n2356 9.3005
R10940 GND.n2355 GND.n2337 9.3005
R10941 GND.n2354 GND.n2353 9.3005
R10942 GND.n2339 GND.n2338 9.3005
R10943 GND.n2347 GND.n2346 9.3005
R10944 GND.n2345 GND.n2342 9.3005
R10945 GND.n2344 GND.n2343 9.3005
R10946 GND.n2369 GND.n2366 9.3005
R10947 GND.n2401 GND.n2398 9.3005
R10948 GND.n2503 GND.n2502 9.3005
R10949 GND.n5131 GND.n1882 9.3005
R10950 GND.n5130 GND.n1883 9.3005
R10951 GND.n2260 GND.n1884 9.3005
R10952 GND.n2593 GND.n2592 9.3005
R10953 GND.n2594 GND.n2259 9.3005
R10954 GND.n2598 GND.n2595 9.3005
R10955 GND.n2597 GND.n2596 9.3005
R10956 GND.n2238 GND.n2237 9.3005
R10957 GND.n2617 GND.n2616 9.3005
R10958 GND.n2618 GND.n2236 9.3005
R10959 GND.n2622 GND.n2619 9.3005
R10960 GND.n2621 GND.n2620 9.3005
R10961 GND.n2204 GND.n2203 9.3005
R10962 GND.n2667 GND.n2666 9.3005
R10963 GND.n2668 GND.n2202 9.3005
R10964 GND.n2670 GND.n2669 9.3005
R10965 GND.n2671 GND.n2141 9.3005
R10966 GND.n2771 GND.n2768 9.3005
R10967 GND.n2770 GND.n2769 9.3005
R10968 GND.n2121 GND.n2120 9.3005
R10969 GND.n2791 GND.n2790 9.3005
R10970 GND.n2792 GND.n2119 9.3005
R10971 GND.n2796 GND.n2793 9.3005
R10972 GND.n2795 GND.n2794 9.3005
R10973 GND.n2100 GND.n2099 9.3005
R10974 GND.n2817 GND.n2816 9.3005
R10975 GND.n2818 GND.n2098 9.3005
R10976 GND.n2820 GND.n2819 9.3005
R10977 GND.n2076 GND.n2075 9.3005
R10978 GND.n2897 GND.n2896 9.3005
R10979 GND.n2898 GND.n2074 9.3005
R10980 GND.n2902 GND.n2899 9.3005
R10981 GND.n2901 GND.n2900 9.3005
R10982 GND.n1993 GND.n1992 9.3005
R10983 GND.n5054 GND.n5053 9.3005
R10984 GND.n5132 GND.n1881 9.3005
R10985 GND.n2767 GND.n2140 9.3005
R10986 GND.n1687 GND.n1686 9.3005
R10987 GND.n1692 GND.n1691 9.3005
R10988 GND.n5316 GND.n1693 9.3005
R10989 GND.n5315 GND.n1694 9.3005
R10990 GND.n5314 GND.n1695 9.3005
R10991 GND.n1700 GND.n1696 9.3005
R10992 GND.n5308 GND.n1701 9.3005
R10993 GND.n5307 GND.n1702 9.3005
R10994 GND.n5306 GND.n1703 9.3005
R10995 GND.n1708 GND.n1704 9.3005
R10996 GND.n5300 GND.n1709 9.3005
R10997 GND.n5299 GND.n1710 9.3005
R10998 GND.n5298 GND.n1711 9.3005
R10999 GND.n1716 GND.n1712 9.3005
R11000 GND.n5292 GND.n1717 9.3005
R11001 GND.n5291 GND.n1718 9.3005
R11002 GND.n5290 GND.n1719 9.3005
R11003 GND.n1724 GND.n1720 9.3005
R11004 GND.n5284 GND.n1725 9.3005
R11005 GND.n5283 GND.n1726 9.3005
R11006 GND.n5282 GND.n1727 9.3005
R11007 GND.n1732 GND.n1728 9.3005
R11008 GND.n5276 GND.n1733 9.3005
R11009 GND.n5275 GND.n1734 9.3005
R11010 GND.n5274 GND.n1735 9.3005
R11011 GND.n1740 GND.n1736 9.3005
R11012 GND.n5268 GND.n1741 9.3005
R11013 GND.n5267 GND.n1742 9.3005
R11014 GND.n5266 GND.n1743 9.3005
R11015 GND.n1748 GND.n1744 9.3005
R11016 GND.n5260 GND.n1749 9.3005
R11017 GND.n5259 GND.n1750 9.3005
R11018 GND.n5258 GND.n1751 9.3005
R11019 GND.n1756 GND.n1752 9.3005
R11020 GND.n5252 GND.n1757 9.3005
R11021 GND.n5251 GND.n1758 9.3005
R11022 GND.n5250 GND.n1759 9.3005
R11023 GND.n1764 GND.n1760 9.3005
R11024 GND.n5244 GND.n1765 9.3005
R11025 GND.n5243 GND.n1766 9.3005
R11026 GND.n5242 GND.n1767 9.3005
R11027 GND.n1772 GND.n1768 9.3005
R11028 GND.n5236 GND.n1773 9.3005
R11029 GND.n5235 GND.n1774 9.3005
R11030 GND.n5234 GND.n1775 9.3005
R11031 GND.n1780 GND.n1776 9.3005
R11032 GND.n5228 GND.n1781 9.3005
R11033 GND.n5227 GND.n1782 9.3005
R11034 GND.n5226 GND.n1783 9.3005
R11035 GND.n1788 GND.n1784 9.3005
R11036 GND.n5220 GND.n1789 9.3005
R11037 GND.n5219 GND.n1790 9.3005
R11038 GND.n5218 GND.n1791 9.3005
R11039 GND.n1796 GND.n1792 9.3005
R11040 GND.n5212 GND.n1797 9.3005
R11041 GND.n5211 GND.n1798 9.3005
R11042 GND.n5210 GND.n1799 9.3005
R11043 GND.n1804 GND.n1800 9.3005
R11044 GND.n5204 GND.n1805 9.3005
R11045 GND.n5203 GND.n1806 9.3005
R11046 GND.n5202 GND.n1807 9.3005
R11047 GND.n1812 GND.n1808 9.3005
R11048 GND.n5196 GND.n1813 9.3005
R11049 GND.n5195 GND.n1814 9.3005
R11050 GND.n5194 GND.n1815 9.3005
R11051 GND.n1820 GND.n1816 9.3005
R11052 GND.n5188 GND.n1821 9.3005
R11053 GND.n5187 GND.n1822 9.3005
R11054 GND.n5186 GND.n1823 9.3005
R11055 GND.n1828 GND.n1824 9.3005
R11056 GND.n5180 GND.n1829 9.3005
R11057 GND.n5179 GND.n1830 9.3005
R11058 GND.n5178 GND.n1831 9.3005
R11059 GND.n1836 GND.n1832 9.3005
R11060 GND.n5172 GND.n1837 9.3005
R11061 GND.n5171 GND.n1838 9.3005
R11062 GND.n5170 GND.n1839 9.3005
R11063 GND.n1844 GND.n1840 9.3005
R11064 GND.n5164 GND.n1845 9.3005
R11065 GND.n5163 GND.n1846 9.3005
R11066 GND.n5162 GND.n1847 9.3005
R11067 GND.n1852 GND.n1848 9.3005
R11068 GND.n5156 GND.n1853 9.3005
R11069 GND.n5155 GND.n1854 9.3005
R11070 GND.n5154 GND.n1855 9.3005
R11071 GND.n1860 GND.n1856 9.3005
R11072 GND.n5148 GND.n1861 9.3005
R11073 GND.n5147 GND.n1862 9.3005
R11074 GND.n5146 GND.n1863 9.3005
R11075 GND.n1868 GND.n1864 9.3005
R11076 GND.n5140 GND.n1869 9.3005
R11077 GND.n5139 GND.n1870 9.3005
R11078 GND.n5138 GND.n1871 9.3005
R11079 GND.n2554 GND.n1872 9.3005
R11080 GND.n2556 GND.n2555 9.3005
R11081 GND.n2553 GND.n2552 9.3005
R11082 GND.n2561 GND.n2560 9.3005
R11083 GND.n2562 GND.n2551 9.3005
R11084 GND.n2583 GND.n2563 9.3005
R11085 GND.n2582 GND.n2564 9.3005
R11086 GND.n2581 GND.n2565 9.3005
R11087 GND.n2568 GND.n2566 9.3005
R11088 GND.n2577 GND.n2569 9.3005
R11089 GND.n2576 GND.n2570 9.3005
R11090 GND.n2575 GND.n2571 9.3005
R11091 GND.n2573 GND.n2572 9.3005
R11092 GND.n2219 GND.n2218 9.3005
R11093 GND.n2640 GND.n2639 9.3005
R11094 GND.n2641 GND.n2217 9.3005
R11095 GND.n2658 GND.n2642 9.3005
R11096 GND.n2657 GND.n2643 9.3005
R11097 GND.n2656 GND.n2644 9.3005
R11098 GND.n5324 GND.n5323 9.3005
R11099 GND.n5327 GND.n1685 9.3005
R11100 GND.n1684 GND.n1680 9.3005
R11101 GND.n5334 GND.n1679 9.3005
R11102 GND.n5335 GND.n1678 9.3005
R11103 GND.n5336 GND.n1677 9.3005
R11104 GND.n1676 GND.n1672 9.3005
R11105 GND.n5342 GND.n1671 9.3005
R11106 GND.n5343 GND.n1670 9.3005
R11107 GND.n5344 GND.n1669 9.3005
R11108 GND.n1668 GND.n1664 9.3005
R11109 GND.n5350 GND.n1663 9.3005
R11110 GND.n5351 GND.n1662 9.3005
R11111 GND.n5352 GND.n1661 9.3005
R11112 GND.n1660 GND.n1656 9.3005
R11113 GND.n5358 GND.n1655 9.3005
R11114 GND.n5359 GND.n1654 9.3005
R11115 GND.n5360 GND.n1653 9.3005
R11116 GND.n1652 GND.n1648 9.3005
R11117 GND.n5366 GND.n1647 9.3005
R11118 GND.n5367 GND.n1646 9.3005
R11119 GND.n5368 GND.n1645 9.3005
R11120 GND.n1644 GND.n1640 9.3005
R11121 GND.n5374 GND.n1639 9.3005
R11122 GND.n5375 GND.n1638 9.3005
R11123 GND.n5376 GND.n1637 9.3005
R11124 GND.n1636 GND.n1632 9.3005
R11125 GND.n5382 GND.n1631 9.3005
R11126 GND.n5383 GND.n1630 9.3005
R11127 GND.n5384 GND.n1629 9.3005
R11128 GND.n1628 GND.n1624 9.3005
R11129 GND.n5390 GND.n1623 9.3005
R11130 GND.n5391 GND.n1622 9.3005
R11131 GND.n5392 GND.n1621 9.3005
R11132 GND.n1620 GND.n1616 9.3005
R11133 GND.n5398 GND.n1615 9.3005
R11134 GND.n5399 GND.n1614 9.3005
R11135 GND.n5400 GND.n1613 9.3005
R11136 GND.n1612 GND.n1608 9.3005
R11137 GND.n5406 GND.n1607 9.3005
R11138 GND.n5407 GND.n1606 9.3005
R11139 GND.n5408 GND.n1605 9.3005
R11140 GND.n1604 GND.n1600 9.3005
R11141 GND.n5414 GND.n1599 9.3005
R11142 GND.n5415 GND.n1598 9.3005
R11143 GND.n5416 GND.n1597 9.3005
R11144 GND.n5326 GND.n5325 9.3005
R11145 GND.n2686 GND.n2185 9.3005
R11146 GND.n2688 GND.n2687 9.3005
R11147 GND.n2689 GND.n2184 9.3005
R11148 GND.n2691 GND.n2690 9.3005
R11149 GND.n2132 GND.n2131 9.3005
R11150 GND.n2776 GND.n2775 9.3005
R11151 GND.n2777 GND.n2129 9.3005
R11152 GND.n2780 GND.n2779 9.3005
R11153 GND.n2778 GND.n2130 9.3005
R11154 GND.n2112 GND.n2111 9.3005
R11155 GND.n2801 GND.n2800 9.3005
R11156 GND.n2802 GND.n2109 9.3005
R11157 GND.n2808 GND.n2807 9.3005
R11158 GND.n2806 GND.n2110 9.3005
R11159 GND.n2805 GND.n2804 9.3005
R11160 GND.n2088 GND.n2086 9.3005
R11161 GND.n2889 GND.n2888 9.3005
R11162 GND.n2887 GND.n2087 9.3005
R11163 GND.n2886 GND.n2885 9.3005
R11164 GND.n2884 GND.n2089 9.3005
R11165 GND.n2883 GND.n2882 9.3005
R11166 GND.n2881 GND.n2840 9.3005
R11167 GND.n2880 GND.n2879 9.3005
R11168 GND.n2850 GND.n2849 9.3005
R11169 GND.n2853 GND.n2845 9.3005
R11170 GND.n2857 GND.n2856 9.3005
R11171 GND.n2858 GND.n2844 9.3005
R11172 GND.n2860 GND.n2859 9.3005
R11173 GND.n2863 GND.n2843 9.3005
R11174 GND.n2867 GND.n2866 9.3005
R11175 GND.n2868 GND.n2842 9.3005
R11176 GND.n2870 GND.n2869 9.3005
R11177 GND.n2875 GND.n2841 9.3005
R11178 GND.n2878 GND.n2877 9.3005
R11179 GND.n2848 GND.n2847 9.3005
R11180 GND.n5013 GND.n2029 9.3005
R11181 GND.n5015 GND.n5014 9.3005
R11182 GND.n5016 GND.n2028 9.3005
R11183 GND.n5018 GND.n5017 9.3005
R11184 GND.n5019 GND.n2022 9.3005
R11185 GND.n5021 GND.n5020 9.3005
R11186 GND.n5022 GND.n2021 9.3005
R11187 GND.n5024 GND.n5023 9.3005
R11188 GND.n5025 GND.n2017 9.3005
R11189 GND.n5027 GND.n5026 9.3005
R11190 GND.n5028 GND.n2016 9.3005
R11191 GND.n5030 GND.n5029 9.3005
R11192 GND.n5031 GND.n2012 9.3005
R11193 GND.n5033 GND.n5032 9.3005
R11194 GND.n5034 GND.n2011 9.3005
R11195 GND.n5036 GND.n5035 9.3005
R11196 GND.n5037 GND.n2008 9.3005
R11197 GND.n5038 GND.n2003 9.3005
R11198 GND.n5040 GND.n5039 9.3005
R11199 GND.n5041 GND.n2002 9.3005
R11200 GND.n5043 GND.n5042 9.3005
R11201 GND.n5044 GND.n1998 9.3005
R11202 GND.n5046 GND.n5045 9.3005
R11203 GND.n5047 GND.n1997 9.3005
R11204 GND.n5049 GND.n5048 9.3005
R11205 GND.n5050 GND.n1994 9.3005
R11206 GND.n5052 GND.n5051 9.3005
R11207 GND.n4893 GND.n4889 9.3005
R11208 GND.n5005 GND.n5004 9.3005
R11209 GND.n5003 GND.n4891 9.3005
R11210 GND.n5002 GND.n5001 9.3005
R11211 GND.n5000 GND.n4894 9.3005
R11212 GND.n4999 GND.n4998 9.3005
R11213 GND.n4997 GND.n4996 9.3005
R11214 GND.n4995 GND.n4903 9.3005
R11215 GND.n4994 GND.n4993 9.3005
R11216 GND.n4992 GND.n4908 9.3005
R11217 GND.n4991 GND.n4990 9.3005
R11218 GND.n4989 GND.n4909 9.3005
R11219 GND.n4988 GND.n4987 9.3005
R11220 GND.n4986 GND.n4916 9.3005
R11221 GND.n4985 GND.n4984 9.3005
R11222 GND.n4983 GND.n4917 9.3005
R11223 GND.n4982 GND.n4981 9.3005
R11224 GND.n4980 GND.n4924 9.3005
R11225 GND.n4979 GND.n4978 9.3005
R11226 GND.n4977 GND.n4925 9.3005
R11227 GND.n4976 GND.n4975 9.3005
R11228 GND.n4974 GND.n4935 9.3005
R11229 GND.n4973 GND.n4972 9.3005
R11230 GND.n4971 GND.n4936 9.3005
R11231 GND.n4970 GND.n4969 9.3005
R11232 GND.n4968 GND.n4943 9.3005
R11233 GND.n4967 GND.n4966 9.3005
R11234 GND.n4965 GND.n4944 9.3005
R11235 GND.n4964 GND.n4963 9.3005
R11236 GND.n4962 GND.n4951 9.3005
R11237 GND.n4961 GND.n4960 9.3005
R11238 GND.n4959 GND.n4952 9.3005
R11239 GND.n1894 GND.n1892 9.3005
R11240 GND.n5126 GND.n5125 9.3005
R11241 GND.n1895 GND.n1893 9.3005
R11242 GND.n5121 GND.n1900 9.3005
R11243 GND.n5120 GND.n1901 9.3005
R11244 GND.n5119 GND.n1902 9.3005
R11245 GND.n2244 GND.n1903 9.3005
R11246 GND.n5115 GND.n1908 9.3005
R11247 GND.n5114 GND.n1909 9.3005
R11248 GND.n5113 GND.n1910 9.3005
R11249 GND.n2232 GND.n1911 9.3005
R11250 GND.n5109 GND.n1916 9.3005
R11251 GND.n5108 GND.n1917 9.3005
R11252 GND.n5107 GND.n1918 9.3005
R11253 GND.n2212 GND.n1919 9.3005
R11254 GND.n5103 GND.n1924 9.3005
R11255 GND.n5102 GND.n1925 9.3005
R11256 GND.n5101 GND.n1926 9.3005
R11257 GND.n2153 GND.n1927 9.3005
R11258 GND.n5097 GND.n1932 9.3005
R11259 GND.n5096 GND.n1933 9.3005
R11260 GND.n5095 GND.n1934 9.3005
R11261 GND.n2168 GND.n1935 9.3005
R11262 GND.n5091 GND.n1940 9.3005
R11263 GND.n5090 GND.n1941 9.3005
R11264 GND.n5089 GND.n1942 9.3005
R11265 GND.n2181 GND.n1943 9.3005
R11266 GND.n5085 GND.n1948 9.3005
R11267 GND.n5084 GND.n1949 9.3005
R11268 GND.n5083 GND.n1950 9.3005
R11269 GND.n2127 GND.n1951 9.3005
R11270 GND.n5079 GND.n1956 9.3005
R11271 GND.n5078 GND.n1957 9.3005
R11272 GND.n5077 GND.n1958 9.3005
R11273 GND.n2106 GND.n1959 9.3005
R11274 GND.n5073 GND.n1964 9.3005
R11275 GND.n5072 GND.n1965 9.3005
R11276 GND.n5071 GND.n1966 9.3005
R11277 GND.n2082 GND.n1967 9.3005
R11278 GND.n5067 GND.n1972 9.3005
R11279 GND.n5066 GND.n1973 9.3005
R11280 GND.n5065 GND.n1974 9.3005
R11281 GND.n2069 GND.n1975 9.3005
R11282 GND.n5061 GND.n1980 9.3005
R11283 GND.n5060 GND.n1981 9.3005
R11284 GND.n5059 GND.n1982 9.3005
R11285 GND.n2506 GND.n2504 9.3005
R11286 GND.n1896 GND.n1894 9.3005
R11287 GND.n5125 GND.n5124 9.3005
R11288 GND.n5123 GND.n1895 9.3005
R11289 GND.n5122 GND.n5121 9.3005
R11290 GND.n5120 GND.n1899 9.3005
R11291 GND.n5119 GND.n5118 9.3005
R11292 GND.n5117 GND.n1903 9.3005
R11293 GND.n5116 GND.n5115 9.3005
R11294 GND.n5114 GND.n1907 9.3005
R11295 GND.n5113 GND.n5112 9.3005
R11296 GND.n5111 GND.n1911 9.3005
R11297 GND.n5110 GND.n5109 9.3005
R11298 GND.n5108 GND.n1915 9.3005
R11299 GND.n5107 GND.n5106 9.3005
R11300 GND.n5105 GND.n1919 9.3005
R11301 GND.n5104 GND.n5103 9.3005
R11302 GND.n5102 GND.n1923 9.3005
R11303 GND.n5101 GND.n5100 9.3005
R11304 GND.n5099 GND.n1927 9.3005
R11305 GND.n5098 GND.n5097 9.3005
R11306 GND.n5096 GND.n1931 9.3005
R11307 GND.n5095 GND.n5094 9.3005
R11308 GND.n5093 GND.n1935 9.3005
R11309 GND.n5092 GND.n5091 9.3005
R11310 GND.n5090 GND.n1939 9.3005
R11311 GND.n5089 GND.n5088 9.3005
R11312 GND.n5087 GND.n1943 9.3005
R11313 GND.n5086 GND.n5085 9.3005
R11314 GND.n5084 GND.n1947 9.3005
R11315 GND.n5083 GND.n5082 9.3005
R11316 GND.n5081 GND.n1951 9.3005
R11317 GND.n5080 GND.n5079 9.3005
R11318 GND.n5078 GND.n1955 9.3005
R11319 GND.n5077 GND.n5076 9.3005
R11320 GND.n5075 GND.n1959 9.3005
R11321 GND.n5074 GND.n5073 9.3005
R11322 GND.n5072 GND.n1963 9.3005
R11323 GND.n5071 GND.n5070 9.3005
R11324 GND.n5069 GND.n1967 9.3005
R11325 GND.n5068 GND.n5067 9.3005
R11326 GND.n5066 GND.n1971 9.3005
R11327 GND.n5065 GND.n5064 9.3005
R11328 GND.n5063 GND.n1975 9.3005
R11329 GND.n5062 GND.n5061 9.3005
R11330 GND.n5060 GND.n1979 9.3005
R11331 GND.n5059 GND.n5058 9.3005
R11332 GND.n2506 GND.n2505 9.3005
R11333 GND.n2530 GND.n2529 9.3005
R11334 GND.n2528 GND.n2271 9.3005
R11335 GND.n2527 GND.n2526 9.3005
R11336 GND.n2273 GND.n2272 9.3005
R11337 GND.n2520 GND.n2519 9.3005
R11338 GND.n2518 GND.n2275 9.3005
R11339 GND.n2517 GND.n2516 9.3005
R11340 GND.n2277 GND.n2276 9.3005
R11341 GND.n2510 GND.n2509 9.3005
R11342 GND.n2508 GND.n2279 9.3005
R11343 GND.n2269 GND.n2266 9.3005
R11344 GND.n2536 GND.n2535 9.3005
R11345 GND.n2542 GND.n2265 9.3005
R11346 GND.n2544 GND.n2543 9.3005
R11347 GND.n2545 GND.n2264 9.3005
R11348 GND.n2547 GND.n2546 9.3005
R11349 GND.n2251 GND.n2250 9.3005
R11350 GND.n2603 GND.n2602 9.3005
R11351 GND.n2604 GND.n2248 9.3005
R11352 GND.n2607 GND.n2606 9.3005
R11353 GND.n2605 GND.n2249 9.3005
R11354 GND.n2227 GND.n2226 9.3005
R11355 GND.n2627 GND.n2626 9.3005
R11356 GND.n2628 GND.n2224 9.3005
R11357 GND.n2633 GND.n2632 9.3005
R11358 GND.n2631 GND.n2225 9.3005
R11359 GND.n2630 GND.n2629 9.3005
R11360 GND.n2193 GND.n2192 9.3005
R11361 GND.n2676 GND.n2675 9.3005
R11362 GND.n2677 GND.n2190 9.3005
R11363 GND.n2679 GND.n2678 9.3005
R11364 GND.n2680 GND.n2189 9.3005
R11365 GND.n2682 GND.n2681 9.3005
R11366 GND.n2683 GND.n2186 9.3005
R11367 GND.n2538 GND.n2537 9.3005
R11368 GND.n2685 GND.n2684 9.3005
R11369 GND.n2712 GND.t16 8.87284
R11370 GND.n3532 GND.n3529 8.87284
R11371 GND.t96 GND.n3006 8.87284
R11372 GND.n3382 GND.n3381 8.87284
R11373 GND.n3643 GND.n3642 8.87284
R11374 GND.n3685 GND.n3361 8.87284
R11375 GND.n4713 GND.n3186 8.87284
R11376 GND.t170 GND.t152 8.87284
R11377 GND.n3829 GND.t226 8.87284
R11378 GND.t4 GND.n3995 8.87284
R11379 GND.n4960 GND.n4951 8.53383
R11380 GND.n4229 GND.n4138 8.53383
R11381 GND.n6678 GND.n6677 8.53383
R11382 GND.n2497 GND.n2283 8.53383
R11383 GND.n4888 GND.n2032 8.19036
R11384 GND.n3615 GND.n3382 8.19036
R11385 GND.n3643 GND.n3375 8.19036
R11386 GND.n3685 GND.n3684 8.19036
R11387 GND.n4714 GND.n4713 8.19036
R11388 GND.n4631 GND.n3923 8.19036
R11389 GND.n6859 GND.n6858 8.09467
R11390 GND.n2684 GND.n263 8.09467
R11391 GND.n5019 GND.n5018 7.95202
R11392 GND.n4588 GND.n4587 7.95202
R11393 GND.n6749 GND.n690 7.95202
R11394 GND.n2401 GND.n2319 7.95202
R11395 GND.n2955 GND.n2949 7.50787
R11396 GND.n3575 GND.n3387 7.50787
R11397 GND.n3651 GND.n3650 7.50787
R11398 GND.n3666 GND.n3123 7.50787
R11399 GND.n3320 GND.n3195 7.50787
R11400 GND.n3829 GND.n3823 7.50787
R11401 GND.n86 GND.n42 7.44662
R11402 GND.n350 GND.n306 7.44662
R11403 GND.n4804 GND.t195 6.82538
R11404 GND.n3620 GND.n3035 6.82538
R11405 GND.n3632 GND.n3053 6.82538
R11406 GND.n3699 GND.n3354 6.82538
R11407 GND.n4720 GND.n3175 6.82538
R11408 GND.t99 GND.n3192 6.82538
R11409 GND.n3839 GND.t103 6.82538
R11410 GND.t183 GND.n4670 6.82538
R11411 GND.n263 GND.n262 6.60521
R11412 GND.n6859 GND.n526 6.60521
R11413 GND.n2732 GND.t31 6.14289
R11414 GND.n4853 GND.n4852 6.14289
R11415 GND.n3553 GND.n3552 6.14289
R11416 GND.n4817 GND.t116 6.14289
R11417 GND.n3557 GND.n2989 6.14289
R11418 GND.n3656 GND.n3103 6.14289
R11419 GND.n3368 GND.n3106 6.14289
R11420 GND.n4699 GND.n3206 6.14289
R11421 GND.n4693 GND.n3212 6.14289
R11422 GND.n3824 GND.n3215 6.14289
R11423 GND.t103 GND.n3234 6.14289
R11424 GND.n4090 GND.t14 6.14289
R11425 GND.n4828 GND.n4827 5.62474
R11426 GND.n3804 GND.n3759 5.62474
R11427 GND.n3626 GND.n3037 5.4604
R11428 GND.n3628 GND.n3051 5.4604
R11429 GND.n4728 GND.n4727 5.4604
R11430 GND.n3709 GND.n3708 5.4604
R11431 GND.t93 GND.n3206 5.4604
R11432 GND.n4928 GND.n4924 5.23686
R11433 GND.n4199 GND.n4196 5.23686
R11434 GND.n6702 GND.n6701 5.23686
R11435 GND.n2467 GND.n2466 5.23686
R11436 GND.n238 GND.t27 5.18375
R11437 GND.n238 GND.t34 5.18375
R11438 GND.n240 GND.t59 5.18375
R11439 GND.n240 GND.t43 5.18375
R11440 GND.n194 GND.t57 5.18375
R11441 GND.n194 GND.t61 5.18375
R11442 GND.n196 GND.t80 5.18375
R11443 GND.n196 GND.t62 5.18375
R11444 GND.n150 GND.t29 5.18375
R11445 GND.n150 GND.t35 5.18375
R11446 GND.n152 GND.t60 5.18375
R11447 GND.n152 GND.t44 5.18375
R11448 GND.n106 GND.t70 5.18375
R11449 GND.n106 GND.t48 5.18375
R11450 GND.n108 GND.t54 5.18375
R11451 GND.n108 GND.t72 5.18375
R11452 GND.n62 GND.t67 5.18375
R11453 GND.n62 GND.t73 5.18375
R11454 GND.n64 GND.t40 5.18375
R11455 GND.n64 GND.t68 5.18375
R11456 GND.n19 GND.t23 5.18375
R11457 GND.n19 GND.t32 5.18375
R11458 GND.n21 GND.t81 5.18375
R11459 GND.n21 GND.t21 5.18375
R11460 GND.n504 GND.t85 5.18375
R11461 GND.n504 GND.t12 5.18375
R11462 GND.n502 GND.t83 5.18375
R11463 GND.n502 GND.t9 5.18375
R11464 GND.n460 GND.t25 5.18375
R11465 GND.n460 GND.t38 5.18375
R11466 GND.n458 GND.t15 5.18375
R11467 GND.n458 GND.t30 5.18375
R11468 GND.n416 GND.t86 5.18375
R11469 GND.n416 GND.t13 5.18375
R11470 GND.n414 GND.t84 5.18375
R11471 GND.n414 GND.t10 5.18375
R11472 GND.n372 GND.t75 5.18375
R11473 GND.n372 GND.t77 5.18375
R11474 GND.n370 GND.t49 5.18375
R11475 GND.n370 GND.t51 5.18375
R11476 GND.n328 GND.t74 5.18375
R11477 GND.n328 GND.t76 5.18375
R11478 GND.n326 GND.t79 5.18375
R11479 GND.n326 GND.t78 5.18375
R11480 GND.n285 GND.t36 5.18375
R11481 GND.n285 GND.t37 5.18375
R11482 GND.n283 GND.t45 5.18375
R11483 GND.n283 GND.t46 5.18375
R11484 GND.n3444 GND.n3418 5.11262
R11485 GND.n3433 GND.n3421 5.11262
R11486 GND.n3257 GND.n3256 5.11262
R11487 GND.n3264 GND.n3249 5.11262
R11488 GND.n262 GND.n261 4.94662
R11489 GND.n526 GND.n525 4.94662
R11490 GND.n218 GND.n217 4.88412
R11491 GND.n174 GND.n173 4.88412
R11492 GND.n130 GND.n129 4.88412
R11493 GND.n86 GND.n85 4.88412
R11494 GND.n482 GND.n481 4.88412
R11495 GND.n438 GND.n437 4.88412
R11496 GND.n394 GND.n393 4.88412
R11497 GND.n350 GND.n349 4.88412
R11498 GND.t41 GND.n2229 4.77792
R11499 GND.n3543 GND.n3542 4.77792
R11500 GND.n3576 GND.t96 4.77792
R11501 GND.n3642 GND.t2 4.77792
R11502 GND.n4762 GND.n4761 4.77792
R11503 GND.n3672 GND.n3120 4.77792
R11504 GND.t3 GND.n3361 4.77792
R11505 GND.n3749 GND.n3203 4.77792
R11506 GND.n4692 GND.n4691 4.77792
R11507 GND.t164 GND.n3226 4.77792
R11508 GND.n6611 GND.t6 4.77792
R11509 GND.n4043 GND.n546 4.74817
R11510 GND.n4477 GND.n545 4.74817
R11511 GND.n6853 GND.n539 4.74817
R11512 GND.n6851 GND.n540 4.74817
R11513 GND.n547 GND.n544 4.74817
R11514 GND.n4490 GND.n546 4.74817
R11515 GND.n4044 GND.n545 4.74817
R11516 GND.n4476 GND.n539 4.74817
R11517 GND.n6852 GND.n6851 4.74817
R11518 GND.n4454 GND.n544 4.74817
R11519 GND.n2646 GND.n2645 4.74817
R11520 GND.n2756 GND.n2161 4.74817
R11521 GND.n2754 GND.n2753 4.74817
R11522 GND.n2702 GND.n2701 4.74817
R11523 GND.n2738 GND.n2737 4.74817
R11524 GND.n4484 GND.n4483 4.74817
R11525 GND.n4374 GND.n4037 4.74817
R11526 GND.n4375 GND.n4373 4.74817
R11527 GND.n4382 GND.n4381 4.74817
R11528 GND.n4403 GND.n4402 4.74817
R11529 GND.n4485 GND.n4484 4.74817
R11530 GND.n4482 GND.n4037 4.74817
R11531 GND.n4376 GND.n4375 4.74817
R11532 GND.n4381 GND.n4380 4.74817
R11533 GND.n4404 GND.n4403 4.74817
R11534 GND.n2766 GND.n2765 4.74817
R11535 GND.n2171 GND.n2146 4.74817
R11536 GND.n2747 GND.n2145 4.74817
R11537 GND.n2177 GND.n2144 4.74817
R11538 GND.n2693 GND.n2143 4.74817
R11539 GND.n2766 GND.n2147 4.74817
R11540 GND.n2764 GND.n2146 4.74817
R11541 GND.n2172 GND.n2145 4.74817
R11542 GND.n2748 GND.n2144 4.74817
R11543 GND.n2176 GND.n2143 4.74817
R11544 GND.n2648 GND.n2646 4.74817
R11545 GND.n2647 GND.n2161 4.74817
R11546 GND.n2755 GND.n2754 4.74817
R11547 GND.n2701 GND.n2162 4.74817
R11548 GND.n2739 GND.n2738 4.74817
R11549 GND.n4996 GND.n4902 4.65505
R11550 GND.n4163 GND.n4150 4.65505
R11551 GND.n6725 GND.n6722 4.65505
R11552 GND.n2433 GND.n2307 4.65505
R11553 GND.n4635 GND.n3883 4.6132
R11554 GND.n4892 GND.n2031 4.6132
R11555 GND.n228 GND.n224 4.40546
R11556 GND.n251 GND.n247 4.40546
R11557 GND.n184 GND.n180 4.40546
R11558 GND.n207 GND.n203 4.40546
R11559 GND.n140 GND.n136 4.40546
R11560 GND.n163 GND.n159 4.40546
R11561 GND.n96 GND.n92 4.40546
R11562 GND.n119 GND.n115 4.40546
R11563 GND.n52 GND.n48 4.40546
R11564 GND.n75 GND.n71 4.40546
R11565 GND.n9 GND.n5 4.40546
R11566 GND.n32 GND.n28 4.40546
R11567 GND.n515 GND.n511 4.40546
R11568 GND.n492 GND.n488 4.40546
R11569 GND.n471 GND.n467 4.40546
R11570 GND.n448 GND.n444 4.40546
R11571 GND.n427 GND.n423 4.40546
R11572 GND.n404 GND.n400 4.40546
R11573 GND.n383 GND.n379 4.40546
R11574 GND.n360 GND.n356 4.40546
R11575 GND.n339 GND.n335 4.40546
R11576 GND.n316 GND.n312 4.40546
R11577 GND.n296 GND.n292 4.40546
R11578 GND.n273 GND.n269 4.40546
R11579 GND.n5136 GND.n1874 4.09543
R11580 GND.n4811 GND.t177 4.09543
R11581 GND.n4797 GND.n4796 4.09543
R11582 GND.n3735 GND.n3344 4.09543
R11583 GND.n3232 GND.t164 4.09543
R11584 GND.n4111 GND.t119 4.09543
R11585 GND.n6591 GND.n655 4.09543
R11586 GND.n262 GND.n218 3.65143
R11587 GND.n526 GND.n482 3.65143
R11588 GND.n237 GND.n219 3.49141
R11589 GND.n260 GND.n242 3.49141
R11590 GND.n193 GND.n175 3.49141
R11591 GND.n216 GND.n198 3.49141
R11592 GND.n149 GND.n131 3.49141
R11593 GND.n172 GND.n154 3.49141
R11594 GND.n105 GND.n87 3.49141
R11595 GND.n128 GND.n110 3.49141
R11596 GND.n61 GND.n43 3.49141
R11597 GND.n84 GND.n66 3.49141
R11598 GND.n18 GND.n0 3.49141
R11599 GND.n41 GND.n23 3.49141
R11600 GND.n524 GND.n506 3.49141
R11601 GND.n501 GND.n483 3.49141
R11602 GND.n480 GND.n462 3.49141
R11603 GND.n457 GND.n439 3.49141
R11604 GND.n436 GND.n418 3.49141
R11605 GND.n413 GND.n395 3.49141
R11606 GND.n392 GND.n374 3.49141
R11607 GND.n369 GND.n351 3.49141
R11608 GND.n348 GND.n330 3.49141
R11609 GND.n325 GND.n307 3.49141
R11610 GND.n305 GND.n287 3.49141
R11611 GND.n282 GND.n264 3.49141
R11612 GND.t22 GND.n2180 3.41294
R11613 GND.t223 GND.n4859 3.41294
R11614 GND.n4804 GND.n3006 3.41294
R11615 GND.n4776 GND.t1 3.41294
R11616 GND.n4768 GND.n3081 3.41294
R11617 GND.n4742 GND.n4741 3.41294
R11618 GND.n3692 GND.t0 3.41294
R11619 GND.n4707 GND.n3192 3.41294
R11620 GND.n4685 GND.n3224 3.41294
R11621 GND.n4480 GND.t8 3.41294
R11622 GND.n4803 GND.n3008 2.73045
R11623 GND.n4769 GND.n3079 2.73045
R11624 GND.n3662 GND.n3131 2.73045
R11625 GND.n3729 GND.n3728 2.73045
R11626 GND.n235 GND.n234 2.71565
R11627 GND.n258 GND.n257 2.71565
R11628 GND.n191 GND.n190 2.71565
R11629 GND.n214 GND.n213 2.71565
R11630 GND.n147 GND.n146 2.71565
R11631 GND.n170 GND.n169 2.71565
R11632 GND.n103 GND.n102 2.71565
R11633 GND.n126 GND.n125 2.71565
R11634 GND.n59 GND.n58 2.71565
R11635 GND.n82 GND.n81 2.71565
R11636 GND.n16 GND.n15 2.71565
R11637 GND.n39 GND.n38 2.71565
R11638 GND.n522 GND.n521 2.71565
R11639 GND.n499 GND.n498 2.71565
R11640 GND.n478 GND.n477 2.71565
R11641 GND.n455 GND.n454 2.71565
R11642 GND.n434 GND.n433 2.71565
R11643 GND.n411 GND.n410 2.71565
R11644 GND.n390 GND.n389 2.71565
R11645 GND.n367 GND.n366 2.71565
R11646 GND.n346 GND.n345 2.71565
R11647 GND.n323 GND.n322 2.71565
R11648 GND.n303 GND.n302 2.71565
R11649 GND.n280 GND.n279 2.71565
R11650 GND.n130 GND.n86 2.563
R11651 GND.n174 GND.n130 2.563
R11652 GND.n218 GND.n174 2.563
R11653 GND.n394 GND.n350 2.563
R11654 GND.n438 GND.n394 2.563
R11655 GND.n482 GND.n438 2.563
R11656 GND.n3274 GND.n3248 2.32777
R11657 GND.n6850 GND.n546 2.27742
R11658 GND.n6850 GND.n545 2.27742
R11659 GND.n6850 GND.n539 2.27742
R11660 GND.n6851 GND.n6850 2.27742
R11661 GND.n6850 GND.n544 2.27742
R11662 GND.n4484 GND.n543 2.27742
R11663 GND.n4037 GND.n543 2.27742
R11664 GND.n4375 GND.n543 2.27742
R11665 GND.n4381 GND.n543 2.27742
R11666 GND.n4403 GND.n543 2.27742
R11667 GND.n2767 GND.n2766 2.27742
R11668 GND.n2767 GND.n2146 2.27742
R11669 GND.n2767 GND.n2145 2.27742
R11670 GND.n2767 GND.n2144 2.27742
R11671 GND.n2767 GND.n2143 2.27742
R11672 GND.n2646 GND.n2142 2.27742
R11673 GND.n2161 GND.n2142 2.27742
R11674 GND.n2754 GND.n2142 2.27742
R11675 GND.n2701 GND.n2142 2.27742
R11676 GND.n2738 GND.n2142 2.27742
R11677 GND.n261 GND.n241 2.19016
R11678 GND.n241 GND.n239 2.19016
R11679 GND.n217 GND.n197 2.19016
R11680 GND.n197 GND.n195 2.19016
R11681 GND.n173 GND.n153 2.19016
R11682 GND.n153 GND.n151 2.19016
R11683 GND.n129 GND.n109 2.19016
R11684 GND.n109 GND.n107 2.19016
R11685 GND.n85 GND.n65 2.19016
R11686 GND.n65 GND.n63 2.19016
R11687 GND.n42 GND.n22 2.19016
R11688 GND.n22 GND.n20 2.19016
R11689 GND.n505 GND.n503 2.19016
R11690 GND.n525 GND.n505 2.19016
R11691 GND.n461 GND.n459 2.19016
R11692 GND.n481 GND.n461 2.19016
R11693 GND.n417 GND.n415 2.19016
R11694 GND.n437 GND.n417 2.19016
R11695 GND.n373 GND.n371 2.19016
R11696 GND.n393 GND.n373 2.19016
R11697 GND.n329 GND.n327 2.19016
R11698 GND.n349 GND.n329 2.19016
R11699 GND.n286 GND.n284 2.19016
R11700 GND.n306 GND.n286 2.19016
R11701 GND.t39 GND.n2660 2.04796
R11702 GND.n4865 GND.n2939 2.04796
R11703 GND.n3616 GND.n3026 2.04796
R11704 GND.n3376 GND.n3062 2.04796
R11705 GND.n4735 GND.n3148 2.04796
R11706 GND.n3736 GND.n3183 2.04796
R11707 GND.n4678 GND.n4677 2.04796
R11708 GND.t11 GND.n566 2.04796
R11709 GND.n231 GND.n221 1.93989
R11710 GND.n254 GND.n244 1.93989
R11711 GND.n187 GND.n177 1.93989
R11712 GND.n210 GND.n200 1.93989
R11713 GND.n143 GND.n133 1.93989
R11714 GND.n166 GND.n156 1.93989
R11715 GND.n99 GND.n89 1.93989
R11716 GND.n122 GND.n112 1.93989
R11717 GND.n55 GND.n45 1.93989
R11718 GND.n78 GND.n68 1.93989
R11719 GND.n12 GND.n2 1.93989
R11720 GND.n35 GND.n25 1.93989
R11721 GND.n4999 GND.n4902 1.93989
R11722 GND.n4166 GND.n4163 1.93989
R11723 GND.n6726 GND.n6725 1.93989
R11724 GND.n518 GND.n508 1.93989
R11725 GND.n495 GND.n485 1.93989
R11726 GND.n474 GND.n464 1.93989
R11727 GND.n451 GND.n441 1.93989
R11728 GND.n430 GND.n420 1.93989
R11729 GND.n407 GND.n397 1.93989
R11730 GND.n386 GND.n376 1.93989
R11731 GND.n363 GND.n353 1.93989
R11732 GND.n342 GND.n332 1.93989
R11733 GND.n319 GND.n309 1.93989
R11734 GND.n299 GND.n289 1.93989
R11735 GND.n276 GND.n266 1.93989
R11736 GND.n2434 GND.n2433 1.93989
R11737 GND.n2262 GND.t89 1.36548
R11738 GND.n2904 GND.t122 1.36548
R11739 GND.n3388 GND.n2997 1.36548
R11740 GND.n3652 GND.n3095 1.36548
R11741 GND.n4749 GND.n4748 1.36548
R11742 GND.t180 GND.n3319 1.36548
R11743 GND.t152 GND.n4692 1.36548
R11744 GND.t145 GND.n3944 1.36548
R11745 GND.n6641 GND.t109 1.36548
R11746 GND.n4978 GND.n4928 1.35808
R11747 GND.n4196 GND.n4144 1.35808
R11748 GND.n6701 GND.n6698 1.35808
R11749 GND.n2466 GND.n2295 1.35808
R11750 GND.n3872 GND.n3871 1.24928
R11751 GND.n3402 GND.n3401 1.24928
R11752 GND.n3478 GND.n3409 1.24928
R11753 GND.n4644 GND.n4643 1.24928
R11754 GND.n230 GND.n223 1.16414
R11755 GND.n253 GND.n246 1.16414
R11756 GND.n186 GND.n179 1.16414
R11757 GND.n209 GND.n202 1.16414
R11758 GND.n142 GND.n135 1.16414
R11759 GND.n165 GND.n158 1.16414
R11760 GND.n98 GND.n91 1.16414
R11761 GND.n121 GND.n114 1.16414
R11762 GND.n54 GND.n47 1.16414
R11763 GND.n77 GND.n70 1.16414
R11764 GND.n11 GND.n4 1.16414
R11765 GND.n34 GND.n27 1.16414
R11766 GND.n517 GND.n510 1.16414
R11767 GND.n494 GND.n487 1.16414
R11768 GND.n473 GND.n466 1.16414
R11769 GND.n450 GND.n443 1.16414
R11770 GND.n429 GND.n422 1.16414
R11771 GND.n406 GND.n399 1.16414
R11772 GND.n385 GND.n378 1.16414
R11773 GND.n362 GND.n355 1.16414
R11774 GND.n341 GND.n334 1.16414
R11775 GND.n318 GND.n311 1.16414
R11776 GND.n298 GND.n291 1.16414
R11777 GND.n275 GND.n268 1.16414
R11778 GND.n4879 GND.n2921 1.02423
R11779 GND.n4111 GND.n3282 1.02423
R11780 GND.n4889 GND.n2031 0.970197
R11781 GND.n4829 GND.n4828 0.970197
R11782 GND.n3800 GND.n3759 0.970197
R11783 GND.n4635 GND.n4634 0.970197
R11784 GND GND.n263 0.853393
R11785 GND GND.n6859 0.783912
R11786 GND.n3428 GND.n3426 0.716017
R11787 GND.n3272 GND.n3270 0.716017
R11788 GND.t20 GND.n2152 0.682988
R11789 GND.t186 GND.n2929 0.682988
R11790 GND.n4873 GND.n4872 0.682988
R11791 GND.n3523 GND.t106 0.682988
R11792 GND.n4852 GND.t205 0.682988
R11793 GND.t177 GND.n4810 0.682988
R11794 GND.n4790 GND.n4789 0.682988
R11795 GND.n4783 GND.n4782 0.682988
R11796 GND.t1 GND.n4775 0.682988
R11797 GND.n4734 GND.t0 0.682988
R11798 GND.n3698 GND.n3163 0.682988
R11799 GND.n4721 GND.n3172 0.682988
R11800 GND.n4671 GND.n3242 0.682988
R11801 GND.t24 GND.n4368 0.682988
R11802 GND.n3771 GND.n3770 0.460866
R11803 GND.n3813 GND.n3812 0.460866
R11804 GND.n4821 GND.n4820 0.460866
R11805 GND.n3013 GND.n2967 0.460866
R11806 GND.n6653 GND.n6652 0.447146
R11807 GND.n2537 GND.n2536 0.447146
R11808 GND.n1597 GND.n1592 0.441049
R11809 GND.n6285 GND.n1070 0.441049
R11810 GND.n6404 GND.n6403 0.441049
R11811 GND.n5325 GND.n5324 0.441049
R11812 GND.n6790 GND.n6789 0.434951
R11813 GND.n4549 GND.n4548 0.434951
R11814 GND.n5053 GND.n5052 0.434951
R11815 GND.n2344 GND.n1881 0.434951
R11816 GND.n6850 GND.n543 0.3925
R11817 GND.n2767 GND.n2142 0.3925
R11818 GND.n227 GND.n226 0.388379
R11819 GND.n250 GND.n249 0.388379
R11820 GND.n183 GND.n182 0.388379
R11821 GND.n206 GND.n205 0.388379
R11822 GND.n139 GND.n138 0.388379
R11823 GND.n162 GND.n161 0.388379
R11824 GND.n95 GND.n94 0.388379
R11825 GND.n118 GND.n117 0.388379
R11826 GND.n51 GND.n50 0.388379
R11827 GND.n74 GND.n73 0.388379
R11828 GND.n8 GND.n7 0.388379
R11829 GND.n31 GND.n30 0.388379
R11830 GND.n514 GND.n513 0.388379
R11831 GND.n491 GND.n490 0.388379
R11832 GND.n470 GND.n469 0.388379
R11833 GND.n447 GND.n446 0.388379
R11834 GND.n426 GND.n425 0.388379
R11835 GND.n403 GND.n402 0.388379
R11836 GND.n382 GND.n381 0.388379
R11837 GND.n359 GND.n358 0.388379
R11838 GND.n338 GND.n337 0.388379
R11839 GND.n315 GND.n314 0.388379
R11840 GND.n295 GND.n294 0.388379
R11841 GND.n272 GND.n271 0.388379
R11842 GND.n4636 GND.n3295 0.312695
R11843 GND.n3489 GND.n3404 0.312695
R11844 GND.n3405 GND.n3404 0.312695
R11845 GND.n4637 GND.n4636 0.312695
R11846 GND.n4246 GND.n4103 0.269198
R11847 GND.n2880 GND.n2878 0.269198
R11848 GND.n6674 GND.n6673 0.253549
R11849 GND.n2508 GND.n2507 0.253549
R11850 GND.n6675 GND.n6674 0.241354
R11851 GND.n4270 GND.n4269 0.241354
R11852 GND.n2507 GND.n2503 0.241354
R11853 GND.n4952 GND.n1983 0.241354
R11854 GND.n4580 GND.n3883 0.229039
R11855 GND.n3884 GND.n3883 0.229039
R11856 GND.n4892 GND.n2029 0.229039
R11857 GND.n4893 GND.n4892 0.229039
R11858 GND.n236 GND.n220 0.155672
R11859 GND.n229 GND.n220 0.155672
R11860 GND.n229 GND.n228 0.155672
R11861 GND.n259 GND.n243 0.155672
R11862 GND.n252 GND.n243 0.155672
R11863 GND.n252 GND.n251 0.155672
R11864 GND.n192 GND.n176 0.155672
R11865 GND.n185 GND.n176 0.155672
R11866 GND.n185 GND.n184 0.155672
R11867 GND.n215 GND.n199 0.155672
R11868 GND.n208 GND.n199 0.155672
R11869 GND.n208 GND.n207 0.155672
R11870 GND.n148 GND.n132 0.155672
R11871 GND.n141 GND.n132 0.155672
R11872 GND.n141 GND.n140 0.155672
R11873 GND.n171 GND.n155 0.155672
R11874 GND.n164 GND.n155 0.155672
R11875 GND.n164 GND.n163 0.155672
R11876 GND.n104 GND.n88 0.155672
R11877 GND.n97 GND.n88 0.155672
R11878 GND.n97 GND.n96 0.155672
R11879 GND.n127 GND.n111 0.155672
R11880 GND.n120 GND.n111 0.155672
R11881 GND.n120 GND.n119 0.155672
R11882 GND.n60 GND.n44 0.155672
R11883 GND.n53 GND.n44 0.155672
R11884 GND.n53 GND.n52 0.155672
R11885 GND.n83 GND.n67 0.155672
R11886 GND.n76 GND.n67 0.155672
R11887 GND.n76 GND.n75 0.155672
R11888 GND.n17 GND.n1 0.155672
R11889 GND.n10 GND.n1 0.155672
R11890 GND.n10 GND.n9 0.155672
R11891 GND.n40 GND.n24 0.155672
R11892 GND.n33 GND.n24 0.155672
R11893 GND.n33 GND.n32 0.155672
R11894 GND.n523 GND.n507 0.155672
R11895 GND.n516 GND.n507 0.155672
R11896 GND.n516 GND.n515 0.155672
R11897 GND.n500 GND.n484 0.155672
R11898 GND.n493 GND.n484 0.155672
R11899 GND.n493 GND.n492 0.155672
R11900 GND.n479 GND.n463 0.155672
R11901 GND.n472 GND.n463 0.155672
R11902 GND.n472 GND.n471 0.155672
R11903 GND.n456 GND.n440 0.155672
R11904 GND.n449 GND.n440 0.155672
R11905 GND.n449 GND.n448 0.155672
R11906 GND.n435 GND.n419 0.155672
R11907 GND.n428 GND.n419 0.155672
R11908 GND.n428 GND.n427 0.155672
R11909 GND.n412 GND.n396 0.155672
R11910 GND.n405 GND.n396 0.155672
R11911 GND.n405 GND.n404 0.155672
R11912 GND.n391 GND.n375 0.155672
R11913 GND.n384 GND.n375 0.155672
R11914 GND.n384 GND.n383 0.155672
R11915 GND.n368 GND.n352 0.155672
R11916 GND.n361 GND.n352 0.155672
R11917 GND.n361 GND.n360 0.155672
R11918 GND.n347 GND.n331 0.155672
R11919 GND.n340 GND.n331 0.155672
R11920 GND.n340 GND.n339 0.155672
R11921 GND.n324 GND.n308 0.155672
R11922 GND.n317 GND.n308 0.155672
R11923 GND.n317 GND.n316 0.155672
R11924 GND.n304 GND.n288 0.155672
R11925 GND.n297 GND.n288 0.155672
R11926 GND.n297 GND.n296 0.155672
R11927 GND.n281 GND.n265 0.155672
R11928 GND.n274 GND.n265 0.155672
R11929 GND.n274 GND.n273 0.155672
R11930 GND.n3771 GND.n3768 0.152939
R11931 GND.n3779 GND.n3768 0.152939
R11932 GND.n3780 GND.n3779 0.152939
R11933 GND.n3781 GND.n3780 0.152939
R11934 GND.n3781 GND.n3764 0.152939
R11935 GND.n3789 GND.n3764 0.152939
R11936 GND.n3790 GND.n3789 0.152939
R11937 GND.n3792 GND.n3790 0.152939
R11938 GND.n3792 GND.n3791 0.152939
R11939 GND.n3791 GND.n3760 0.152939
R11940 GND.n3801 GND.n3760 0.152939
R11941 GND.n3803 GND.n3801 0.152939
R11942 GND.n3803 GND.n3802 0.152939
R11943 GND.n3802 GND.n3754 0.152939
R11944 GND.n3812 GND.n3754 0.152939
R11945 GND.n4820 GND.n2985 0.152939
R11946 GND.n3384 GND.n2985 0.152939
R11947 GND.n3579 GND.n3384 0.152939
R11948 GND.n3580 GND.n3579 0.152939
R11949 GND.n3581 GND.n3580 0.152939
R11950 GND.n3582 GND.n3581 0.152939
R11951 GND.n3583 GND.n3582 0.152939
R11952 GND.n3586 GND.n3583 0.152939
R11953 GND.n3587 GND.n3586 0.152939
R11954 GND.n3588 GND.n3587 0.152939
R11955 GND.n3589 GND.n3588 0.152939
R11956 GND.n3590 GND.n3589 0.152939
R11957 GND.n3591 GND.n3590 0.152939
R11958 GND.n3592 GND.n3591 0.152939
R11959 GND.n3594 GND.n3592 0.152939
R11960 GND.n3596 GND.n3594 0.152939
R11961 GND.n3596 GND.n3595 0.152939
R11962 GND.n3595 GND.n3367 0.152939
R11963 GND.n3367 GND.n3365 0.152939
R11964 GND.n3679 GND.n3365 0.152939
R11965 GND.n3680 GND.n3679 0.152939
R11966 GND.n3681 GND.n3680 0.152939
R11967 GND.n3681 GND.n3352 0.152939
R11968 GND.n3702 GND.n3352 0.152939
R11969 GND.n3703 GND.n3702 0.152939
R11970 GND.n3705 GND.n3703 0.152939
R11971 GND.n3705 GND.n3704 0.152939
R11972 GND.n3704 GND.n3346 0.152939
R11973 GND.n3347 GND.n3346 0.152939
R11974 GND.n3348 GND.n3347 0.152939
R11975 GND.n3348 GND.n3315 0.152939
R11976 GND.n3752 GND.n3315 0.152939
R11977 GND.n3753 GND.n3752 0.152939
R11978 GND.n3813 GND.n3753 0.152939
R11979 GND.n2968 GND.n2967 0.152939
R11980 GND.n2969 GND.n2968 0.152939
R11981 GND.n2970 GND.n2969 0.152939
R11982 GND.n2971 GND.n2970 0.152939
R11983 GND.n2972 GND.n2971 0.152939
R11984 GND.n2973 GND.n2972 0.152939
R11985 GND.n2974 GND.n2973 0.152939
R11986 GND.n2975 GND.n2974 0.152939
R11987 GND.n2976 GND.n2975 0.152939
R11988 GND.n2977 GND.n2976 0.152939
R11989 GND.n2978 GND.n2977 0.152939
R11990 GND.n2981 GND.n2978 0.152939
R11991 GND.n2982 GND.n2981 0.152939
R11992 GND.n4822 GND.n2982 0.152939
R11993 GND.n4822 GND.n4821 0.152939
R11994 GND.n3013 GND.n3012 0.152939
R11995 GND.n3019 GND.n3012 0.152939
R11996 GND.n3020 GND.n3019 0.152939
R11997 GND.n3021 GND.n3020 0.152939
R11998 GND.n3022 GND.n3021 0.152939
R11999 GND.n3023 GND.n3022 0.152939
R12000 GND.n3066 GND.n3023 0.152939
R12001 GND.n3067 GND.n3066 0.152939
R12002 GND.n3072 GND.n3067 0.152939
R12003 GND.n3073 GND.n3072 0.152939
R12004 GND.n3074 GND.n3073 0.152939
R12005 GND.n3075 GND.n3074 0.152939
R12006 GND.n3076 GND.n3075 0.152939
R12007 GND.n3110 GND.n3076 0.152939
R12008 GND.n3113 GND.n3110 0.152939
R12009 GND.n3114 GND.n3113 0.152939
R12010 GND.n3115 GND.n3114 0.152939
R12011 GND.n3116 GND.n3115 0.152939
R12012 GND.n3117 GND.n3116 0.152939
R12013 GND.n3153 GND.n3117 0.152939
R12014 GND.n3156 GND.n3153 0.152939
R12015 GND.n3157 GND.n3156 0.152939
R12016 GND.n3158 GND.n3157 0.152939
R12017 GND.n3159 GND.n3158 0.152939
R12018 GND.n3160 GND.n3159 0.152939
R12019 GND.n3177 GND.n3160 0.152939
R12020 GND.n3178 GND.n3177 0.152939
R12021 GND.n3179 GND.n3178 0.152939
R12022 GND.n3180 GND.n3179 0.152939
R12023 GND.n3197 GND.n3180 0.152939
R12024 GND.n3198 GND.n3197 0.152939
R12025 GND.n3199 GND.n3198 0.152939
R12026 GND.n3200 GND.n3199 0.152939
R12027 GND.n3770 GND.n3200 0.152939
R12028 GND.n5423 GND.n1592 0.152939
R12029 GND.n5424 GND.n5423 0.152939
R12030 GND.n5425 GND.n5424 0.152939
R12031 GND.n5425 GND.n1586 0.152939
R12032 GND.n5433 GND.n1586 0.152939
R12033 GND.n5434 GND.n5433 0.152939
R12034 GND.n5435 GND.n5434 0.152939
R12035 GND.n5435 GND.n1580 0.152939
R12036 GND.n5443 GND.n1580 0.152939
R12037 GND.n5444 GND.n5443 0.152939
R12038 GND.n5445 GND.n5444 0.152939
R12039 GND.n5445 GND.n1574 0.152939
R12040 GND.n5453 GND.n1574 0.152939
R12041 GND.n5454 GND.n5453 0.152939
R12042 GND.n5455 GND.n5454 0.152939
R12043 GND.n5455 GND.n1568 0.152939
R12044 GND.n5463 GND.n1568 0.152939
R12045 GND.n5464 GND.n5463 0.152939
R12046 GND.n5465 GND.n5464 0.152939
R12047 GND.n5465 GND.n1562 0.152939
R12048 GND.n5473 GND.n1562 0.152939
R12049 GND.n5474 GND.n5473 0.152939
R12050 GND.n5475 GND.n5474 0.152939
R12051 GND.n5475 GND.n1556 0.152939
R12052 GND.n5483 GND.n1556 0.152939
R12053 GND.n5484 GND.n5483 0.152939
R12054 GND.n5485 GND.n5484 0.152939
R12055 GND.n5485 GND.n1550 0.152939
R12056 GND.n5493 GND.n1550 0.152939
R12057 GND.n5494 GND.n5493 0.152939
R12058 GND.n5495 GND.n5494 0.152939
R12059 GND.n5495 GND.n1544 0.152939
R12060 GND.n5503 GND.n1544 0.152939
R12061 GND.n5504 GND.n5503 0.152939
R12062 GND.n5505 GND.n5504 0.152939
R12063 GND.n5505 GND.n1538 0.152939
R12064 GND.n5513 GND.n1538 0.152939
R12065 GND.n5514 GND.n5513 0.152939
R12066 GND.n5515 GND.n5514 0.152939
R12067 GND.n5515 GND.n1532 0.152939
R12068 GND.n5523 GND.n1532 0.152939
R12069 GND.n5524 GND.n5523 0.152939
R12070 GND.n5525 GND.n5524 0.152939
R12071 GND.n5525 GND.n1526 0.152939
R12072 GND.n5533 GND.n1526 0.152939
R12073 GND.n5534 GND.n5533 0.152939
R12074 GND.n5535 GND.n5534 0.152939
R12075 GND.n5535 GND.n1520 0.152939
R12076 GND.n5543 GND.n1520 0.152939
R12077 GND.n5544 GND.n5543 0.152939
R12078 GND.n5545 GND.n5544 0.152939
R12079 GND.n5545 GND.n1514 0.152939
R12080 GND.n5553 GND.n1514 0.152939
R12081 GND.n5554 GND.n5553 0.152939
R12082 GND.n5555 GND.n5554 0.152939
R12083 GND.n5555 GND.n1508 0.152939
R12084 GND.n5563 GND.n1508 0.152939
R12085 GND.n5564 GND.n5563 0.152939
R12086 GND.n5565 GND.n5564 0.152939
R12087 GND.n5565 GND.n1502 0.152939
R12088 GND.n5573 GND.n1502 0.152939
R12089 GND.n5574 GND.n5573 0.152939
R12090 GND.n5575 GND.n5574 0.152939
R12091 GND.n5575 GND.n1496 0.152939
R12092 GND.n5583 GND.n1496 0.152939
R12093 GND.n5584 GND.n5583 0.152939
R12094 GND.n5585 GND.n5584 0.152939
R12095 GND.n5585 GND.n1490 0.152939
R12096 GND.n5593 GND.n1490 0.152939
R12097 GND.n5594 GND.n5593 0.152939
R12098 GND.n5595 GND.n5594 0.152939
R12099 GND.n5595 GND.n1484 0.152939
R12100 GND.n5603 GND.n1484 0.152939
R12101 GND.n5604 GND.n5603 0.152939
R12102 GND.n5605 GND.n5604 0.152939
R12103 GND.n5605 GND.n1478 0.152939
R12104 GND.n5613 GND.n1478 0.152939
R12105 GND.n5614 GND.n5613 0.152939
R12106 GND.n5615 GND.n5614 0.152939
R12107 GND.n5615 GND.n1472 0.152939
R12108 GND.n5623 GND.n1472 0.152939
R12109 GND.n5624 GND.n5623 0.152939
R12110 GND.n5625 GND.n5624 0.152939
R12111 GND.n5625 GND.n1466 0.152939
R12112 GND.n5633 GND.n1466 0.152939
R12113 GND.n5634 GND.n5633 0.152939
R12114 GND.n5635 GND.n5634 0.152939
R12115 GND.n5635 GND.n1460 0.152939
R12116 GND.n5643 GND.n1460 0.152939
R12117 GND.n5644 GND.n5643 0.152939
R12118 GND.n5645 GND.n5644 0.152939
R12119 GND.n5645 GND.n1454 0.152939
R12120 GND.n5653 GND.n1454 0.152939
R12121 GND.n5654 GND.n5653 0.152939
R12122 GND.n5655 GND.n5654 0.152939
R12123 GND.n5655 GND.n1448 0.152939
R12124 GND.n5663 GND.n1448 0.152939
R12125 GND.n5664 GND.n5663 0.152939
R12126 GND.n5665 GND.n5664 0.152939
R12127 GND.n5665 GND.n1442 0.152939
R12128 GND.n5673 GND.n1442 0.152939
R12129 GND.n5674 GND.n5673 0.152939
R12130 GND.n5675 GND.n5674 0.152939
R12131 GND.n5675 GND.n1436 0.152939
R12132 GND.n5683 GND.n1436 0.152939
R12133 GND.n5684 GND.n5683 0.152939
R12134 GND.n5685 GND.n5684 0.152939
R12135 GND.n5685 GND.n1430 0.152939
R12136 GND.n5693 GND.n1430 0.152939
R12137 GND.n5694 GND.n5693 0.152939
R12138 GND.n5695 GND.n5694 0.152939
R12139 GND.n5695 GND.n1424 0.152939
R12140 GND.n5703 GND.n1424 0.152939
R12141 GND.n5704 GND.n5703 0.152939
R12142 GND.n5705 GND.n5704 0.152939
R12143 GND.n5705 GND.n1418 0.152939
R12144 GND.n5713 GND.n1418 0.152939
R12145 GND.n5714 GND.n5713 0.152939
R12146 GND.n5715 GND.n5714 0.152939
R12147 GND.n5715 GND.n1412 0.152939
R12148 GND.n5723 GND.n1412 0.152939
R12149 GND.n5724 GND.n5723 0.152939
R12150 GND.n5725 GND.n5724 0.152939
R12151 GND.n5725 GND.n1406 0.152939
R12152 GND.n5733 GND.n1406 0.152939
R12153 GND.n5734 GND.n5733 0.152939
R12154 GND.n5735 GND.n5734 0.152939
R12155 GND.n5735 GND.n1400 0.152939
R12156 GND.n5743 GND.n1400 0.152939
R12157 GND.n5744 GND.n5743 0.152939
R12158 GND.n5745 GND.n5744 0.152939
R12159 GND.n5745 GND.n1394 0.152939
R12160 GND.n5753 GND.n1394 0.152939
R12161 GND.n5754 GND.n5753 0.152939
R12162 GND.n5755 GND.n5754 0.152939
R12163 GND.n5755 GND.n1388 0.152939
R12164 GND.n5763 GND.n1388 0.152939
R12165 GND.n5764 GND.n5763 0.152939
R12166 GND.n5765 GND.n5764 0.152939
R12167 GND.n5765 GND.n1382 0.152939
R12168 GND.n5773 GND.n1382 0.152939
R12169 GND.n5774 GND.n5773 0.152939
R12170 GND.n5775 GND.n5774 0.152939
R12171 GND.n5775 GND.n1376 0.152939
R12172 GND.n5783 GND.n1376 0.152939
R12173 GND.n5784 GND.n5783 0.152939
R12174 GND.n5785 GND.n5784 0.152939
R12175 GND.n5785 GND.n1370 0.152939
R12176 GND.n5793 GND.n1370 0.152939
R12177 GND.n5794 GND.n5793 0.152939
R12178 GND.n5795 GND.n5794 0.152939
R12179 GND.n5795 GND.n1364 0.152939
R12180 GND.n5803 GND.n1364 0.152939
R12181 GND.n5804 GND.n5803 0.152939
R12182 GND.n5805 GND.n5804 0.152939
R12183 GND.n5805 GND.n1358 0.152939
R12184 GND.n5813 GND.n1358 0.152939
R12185 GND.n5814 GND.n5813 0.152939
R12186 GND.n5815 GND.n5814 0.152939
R12187 GND.n5815 GND.n1352 0.152939
R12188 GND.n5823 GND.n1352 0.152939
R12189 GND.n5824 GND.n5823 0.152939
R12190 GND.n5825 GND.n5824 0.152939
R12191 GND.n5825 GND.n1346 0.152939
R12192 GND.n5833 GND.n1346 0.152939
R12193 GND.n5834 GND.n5833 0.152939
R12194 GND.n5835 GND.n5834 0.152939
R12195 GND.n5835 GND.n1340 0.152939
R12196 GND.n5843 GND.n1340 0.152939
R12197 GND.n5844 GND.n5843 0.152939
R12198 GND.n5845 GND.n5844 0.152939
R12199 GND.n5845 GND.n1334 0.152939
R12200 GND.n5853 GND.n1334 0.152939
R12201 GND.n5854 GND.n5853 0.152939
R12202 GND.n5855 GND.n5854 0.152939
R12203 GND.n5855 GND.n1328 0.152939
R12204 GND.n5863 GND.n1328 0.152939
R12205 GND.n5864 GND.n5863 0.152939
R12206 GND.n5865 GND.n5864 0.152939
R12207 GND.n5865 GND.n1322 0.152939
R12208 GND.n5873 GND.n1322 0.152939
R12209 GND.n5874 GND.n5873 0.152939
R12210 GND.n5875 GND.n5874 0.152939
R12211 GND.n5875 GND.n1316 0.152939
R12212 GND.n5883 GND.n1316 0.152939
R12213 GND.n5884 GND.n5883 0.152939
R12214 GND.n5885 GND.n5884 0.152939
R12215 GND.n5885 GND.n1310 0.152939
R12216 GND.n5893 GND.n1310 0.152939
R12217 GND.n5894 GND.n5893 0.152939
R12218 GND.n5895 GND.n5894 0.152939
R12219 GND.n5895 GND.n1304 0.152939
R12220 GND.n5903 GND.n1304 0.152939
R12221 GND.n5904 GND.n5903 0.152939
R12222 GND.n5905 GND.n5904 0.152939
R12223 GND.n5905 GND.n1298 0.152939
R12224 GND.n5913 GND.n1298 0.152939
R12225 GND.n5914 GND.n5913 0.152939
R12226 GND.n5915 GND.n5914 0.152939
R12227 GND.n5915 GND.n1292 0.152939
R12228 GND.n5923 GND.n1292 0.152939
R12229 GND.n5924 GND.n5923 0.152939
R12230 GND.n5925 GND.n5924 0.152939
R12231 GND.n5925 GND.n1286 0.152939
R12232 GND.n5933 GND.n1286 0.152939
R12233 GND.n5934 GND.n5933 0.152939
R12234 GND.n5935 GND.n5934 0.152939
R12235 GND.n5935 GND.n1280 0.152939
R12236 GND.n5943 GND.n1280 0.152939
R12237 GND.n5944 GND.n5943 0.152939
R12238 GND.n5945 GND.n5944 0.152939
R12239 GND.n5945 GND.n1274 0.152939
R12240 GND.n5953 GND.n1274 0.152939
R12241 GND.n5954 GND.n5953 0.152939
R12242 GND.n5955 GND.n5954 0.152939
R12243 GND.n5955 GND.n1268 0.152939
R12244 GND.n5963 GND.n1268 0.152939
R12245 GND.n5964 GND.n5963 0.152939
R12246 GND.n5965 GND.n5964 0.152939
R12247 GND.n5965 GND.n1262 0.152939
R12248 GND.n5973 GND.n1262 0.152939
R12249 GND.n5974 GND.n5973 0.152939
R12250 GND.n5975 GND.n5974 0.152939
R12251 GND.n5975 GND.n1256 0.152939
R12252 GND.n5983 GND.n1256 0.152939
R12253 GND.n5984 GND.n5983 0.152939
R12254 GND.n5985 GND.n5984 0.152939
R12255 GND.n5985 GND.n1250 0.152939
R12256 GND.n5993 GND.n1250 0.152939
R12257 GND.n5994 GND.n5993 0.152939
R12258 GND.n5995 GND.n5994 0.152939
R12259 GND.n5995 GND.n1244 0.152939
R12260 GND.n6003 GND.n1244 0.152939
R12261 GND.n6004 GND.n6003 0.152939
R12262 GND.n6005 GND.n6004 0.152939
R12263 GND.n6005 GND.n1238 0.152939
R12264 GND.n6013 GND.n1238 0.152939
R12265 GND.n6014 GND.n6013 0.152939
R12266 GND.n6015 GND.n6014 0.152939
R12267 GND.n6015 GND.n1232 0.152939
R12268 GND.n6023 GND.n1232 0.152939
R12269 GND.n6024 GND.n6023 0.152939
R12270 GND.n6025 GND.n6024 0.152939
R12271 GND.n6025 GND.n1226 0.152939
R12272 GND.n6033 GND.n1226 0.152939
R12273 GND.n6034 GND.n6033 0.152939
R12274 GND.n6035 GND.n6034 0.152939
R12275 GND.n6035 GND.n1220 0.152939
R12276 GND.n6043 GND.n1220 0.152939
R12277 GND.n6044 GND.n6043 0.152939
R12278 GND.n6045 GND.n6044 0.152939
R12279 GND.n6045 GND.n1214 0.152939
R12280 GND.n6053 GND.n1214 0.152939
R12281 GND.n6054 GND.n6053 0.152939
R12282 GND.n6055 GND.n6054 0.152939
R12283 GND.n6055 GND.n1208 0.152939
R12284 GND.n6063 GND.n1208 0.152939
R12285 GND.n6064 GND.n6063 0.152939
R12286 GND.n6065 GND.n6064 0.152939
R12287 GND.n6065 GND.n1202 0.152939
R12288 GND.n6073 GND.n1202 0.152939
R12289 GND.n6074 GND.n6073 0.152939
R12290 GND.n6075 GND.n6074 0.152939
R12291 GND.n6075 GND.n1196 0.152939
R12292 GND.n6083 GND.n1196 0.152939
R12293 GND.n6084 GND.n6083 0.152939
R12294 GND.n6085 GND.n6084 0.152939
R12295 GND.n6085 GND.n1190 0.152939
R12296 GND.n6093 GND.n1190 0.152939
R12297 GND.n6094 GND.n6093 0.152939
R12298 GND.n6095 GND.n6094 0.152939
R12299 GND.n6095 GND.n1184 0.152939
R12300 GND.n6103 GND.n1184 0.152939
R12301 GND.n6104 GND.n6103 0.152939
R12302 GND.n6105 GND.n6104 0.152939
R12303 GND.n6105 GND.n1178 0.152939
R12304 GND.n6113 GND.n1178 0.152939
R12305 GND.n6114 GND.n6113 0.152939
R12306 GND.n6115 GND.n6114 0.152939
R12307 GND.n6115 GND.n1172 0.152939
R12308 GND.n6123 GND.n1172 0.152939
R12309 GND.n6124 GND.n6123 0.152939
R12310 GND.n6125 GND.n6124 0.152939
R12311 GND.n6125 GND.n1166 0.152939
R12312 GND.n6133 GND.n1166 0.152939
R12313 GND.n6134 GND.n6133 0.152939
R12314 GND.n6135 GND.n6134 0.152939
R12315 GND.n6135 GND.n1160 0.152939
R12316 GND.n6143 GND.n1160 0.152939
R12317 GND.n6144 GND.n6143 0.152939
R12318 GND.n6145 GND.n6144 0.152939
R12319 GND.n6145 GND.n1154 0.152939
R12320 GND.n6153 GND.n1154 0.152939
R12321 GND.n6154 GND.n6153 0.152939
R12322 GND.n6155 GND.n6154 0.152939
R12323 GND.n6155 GND.n1148 0.152939
R12324 GND.n6163 GND.n1148 0.152939
R12325 GND.n6164 GND.n6163 0.152939
R12326 GND.n6165 GND.n6164 0.152939
R12327 GND.n6165 GND.n1142 0.152939
R12328 GND.n6173 GND.n1142 0.152939
R12329 GND.n6174 GND.n6173 0.152939
R12330 GND.n6175 GND.n6174 0.152939
R12331 GND.n6175 GND.n1136 0.152939
R12332 GND.n6183 GND.n1136 0.152939
R12333 GND.n6184 GND.n6183 0.152939
R12334 GND.n6185 GND.n6184 0.152939
R12335 GND.n6185 GND.n1130 0.152939
R12336 GND.n6193 GND.n1130 0.152939
R12337 GND.n6194 GND.n6193 0.152939
R12338 GND.n6195 GND.n6194 0.152939
R12339 GND.n6195 GND.n1124 0.152939
R12340 GND.n6203 GND.n1124 0.152939
R12341 GND.n6204 GND.n6203 0.152939
R12342 GND.n6205 GND.n6204 0.152939
R12343 GND.n6205 GND.n1118 0.152939
R12344 GND.n6213 GND.n1118 0.152939
R12345 GND.n6214 GND.n6213 0.152939
R12346 GND.n6215 GND.n6214 0.152939
R12347 GND.n6215 GND.n1112 0.152939
R12348 GND.n6223 GND.n1112 0.152939
R12349 GND.n6224 GND.n6223 0.152939
R12350 GND.n6225 GND.n6224 0.152939
R12351 GND.n6225 GND.n1106 0.152939
R12352 GND.n6233 GND.n1106 0.152939
R12353 GND.n6234 GND.n6233 0.152939
R12354 GND.n6235 GND.n6234 0.152939
R12355 GND.n6235 GND.n1100 0.152939
R12356 GND.n6243 GND.n1100 0.152939
R12357 GND.n6244 GND.n6243 0.152939
R12358 GND.n6245 GND.n6244 0.152939
R12359 GND.n6245 GND.n1094 0.152939
R12360 GND.n6253 GND.n1094 0.152939
R12361 GND.n6254 GND.n6253 0.152939
R12362 GND.n6255 GND.n6254 0.152939
R12363 GND.n6255 GND.n1088 0.152939
R12364 GND.n6263 GND.n1088 0.152939
R12365 GND.n6264 GND.n6263 0.152939
R12366 GND.n6265 GND.n6264 0.152939
R12367 GND.n6265 GND.n1082 0.152939
R12368 GND.n6273 GND.n1082 0.152939
R12369 GND.n6274 GND.n6273 0.152939
R12370 GND.n6275 GND.n6274 0.152939
R12371 GND.n6275 GND.n1076 0.152939
R12372 GND.n6283 GND.n1076 0.152939
R12373 GND.n6284 GND.n6283 0.152939
R12374 GND.n6285 GND.n6284 0.152939
R12375 GND.n6293 GND.n1070 0.152939
R12376 GND.n6294 GND.n6293 0.152939
R12377 GND.n6295 GND.n6294 0.152939
R12378 GND.n6295 GND.n1064 0.152939
R12379 GND.n6303 GND.n1064 0.152939
R12380 GND.n6304 GND.n6303 0.152939
R12381 GND.n6305 GND.n6304 0.152939
R12382 GND.n6305 GND.n1058 0.152939
R12383 GND.n6313 GND.n1058 0.152939
R12384 GND.n6314 GND.n6313 0.152939
R12385 GND.n6315 GND.n6314 0.152939
R12386 GND.n6315 GND.n1052 0.152939
R12387 GND.n6323 GND.n1052 0.152939
R12388 GND.n6324 GND.n6323 0.152939
R12389 GND.n6325 GND.n6324 0.152939
R12390 GND.n6325 GND.n1046 0.152939
R12391 GND.n6333 GND.n1046 0.152939
R12392 GND.n6334 GND.n6333 0.152939
R12393 GND.n6335 GND.n6334 0.152939
R12394 GND.n6335 GND.n1040 0.152939
R12395 GND.n6343 GND.n1040 0.152939
R12396 GND.n6344 GND.n6343 0.152939
R12397 GND.n6345 GND.n6344 0.152939
R12398 GND.n6345 GND.n1034 0.152939
R12399 GND.n6353 GND.n1034 0.152939
R12400 GND.n6354 GND.n6353 0.152939
R12401 GND.n6355 GND.n6354 0.152939
R12402 GND.n6355 GND.n1028 0.152939
R12403 GND.n6363 GND.n1028 0.152939
R12404 GND.n6364 GND.n6363 0.152939
R12405 GND.n6365 GND.n6364 0.152939
R12406 GND.n6365 GND.n1022 0.152939
R12407 GND.n6373 GND.n1022 0.152939
R12408 GND.n6374 GND.n6373 0.152939
R12409 GND.n6375 GND.n6374 0.152939
R12410 GND.n6375 GND.n1016 0.152939
R12411 GND.n6383 GND.n1016 0.152939
R12412 GND.n6384 GND.n6383 0.152939
R12413 GND.n6385 GND.n6384 0.152939
R12414 GND.n6385 GND.n1010 0.152939
R12415 GND.n6393 GND.n1010 0.152939
R12416 GND.n6394 GND.n6393 0.152939
R12417 GND.n6395 GND.n6394 0.152939
R12418 GND.n6395 GND.n1004 0.152939
R12419 GND.n6403 GND.n1004 0.152939
R12420 GND.n4386 GND.n4383 0.152939
R12421 GND.n4387 GND.n4386 0.152939
R12422 GND.n4388 GND.n4387 0.152939
R12423 GND.n4389 GND.n4388 0.152939
R12424 GND.n4391 GND.n4389 0.152939
R12425 GND.n4391 GND.n4390 0.152939
R12426 GND.n4390 GND.n800 0.152939
R12427 GND.n801 GND.n800 0.152939
R12428 GND.n802 GND.n801 0.152939
R12429 GND.n805 GND.n802 0.152939
R12430 GND.n806 GND.n805 0.152939
R12431 GND.n807 GND.n806 0.152939
R12432 GND.n808 GND.n807 0.152939
R12433 GND.n811 GND.n808 0.152939
R12434 GND.n812 GND.n811 0.152939
R12435 GND.n813 GND.n812 0.152939
R12436 GND.n814 GND.n813 0.152939
R12437 GND.n817 GND.n814 0.152939
R12438 GND.n818 GND.n817 0.152939
R12439 GND.n819 GND.n818 0.152939
R12440 GND.n820 GND.n819 0.152939
R12441 GND.n826 GND.n820 0.152939
R12442 GND.n827 GND.n826 0.152939
R12443 GND.n828 GND.n827 0.152939
R12444 GND.n829 GND.n828 0.152939
R12445 GND.n834 GND.n829 0.152939
R12446 GND.n835 GND.n834 0.152939
R12447 GND.n836 GND.n835 0.152939
R12448 GND.n837 GND.n836 0.152939
R12449 GND.n842 GND.n837 0.152939
R12450 GND.n843 GND.n842 0.152939
R12451 GND.n844 GND.n843 0.152939
R12452 GND.n845 GND.n844 0.152939
R12453 GND.n850 GND.n845 0.152939
R12454 GND.n851 GND.n850 0.152939
R12455 GND.n852 GND.n851 0.152939
R12456 GND.n853 GND.n852 0.152939
R12457 GND.n858 GND.n853 0.152939
R12458 GND.n859 GND.n858 0.152939
R12459 GND.n860 GND.n859 0.152939
R12460 GND.n861 GND.n860 0.152939
R12461 GND.n866 GND.n861 0.152939
R12462 GND.n867 GND.n866 0.152939
R12463 GND.n868 GND.n867 0.152939
R12464 GND.n869 GND.n868 0.152939
R12465 GND.n874 GND.n869 0.152939
R12466 GND.n875 GND.n874 0.152939
R12467 GND.n876 GND.n875 0.152939
R12468 GND.n877 GND.n876 0.152939
R12469 GND.n882 GND.n877 0.152939
R12470 GND.n883 GND.n882 0.152939
R12471 GND.n884 GND.n883 0.152939
R12472 GND.n885 GND.n884 0.152939
R12473 GND.n890 GND.n885 0.152939
R12474 GND.n891 GND.n890 0.152939
R12475 GND.n892 GND.n891 0.152939
R12476 GND.n893 GND.n892 0.152939
R12477 GND.n898 GND.n893 0.152939
R12478 GND.n899 GND.n898 0.152939
R12479 GND.n900 GND.n899 0.152939
R12480 GND.n901 GND.n900 0.152939
R12481 GND.n906 GND.n901 0.152939
R12482 GND.n907 GND.n906 0.152939
R12483 GND.n908 GND.n907 0.152939
R12484 GND.n909 GND.n908 0.152939
R12485 GND.n914 GND.n909 0.152939
R12486 GND.n915 GND.n914 0.152939
R12487 GND.n916 GND.n915 0.152939
R12488 GND.n917 GND.n916 0.152939
R12489 GND.n922 GND.n917 0.152939
R12490 GND.n923 GND.n922 0.152939
R12491 GND.n924 GND.n923 0.152939
R12492 GND.n925 GND.n924 0.152939
R12493 GND.n930 GND.n925 0.152939
R12494 GND.n931 GND.n930 0.152939
R12495 GND.n932 GND.n931 0.152939
R12496 GND.n933 GND.n932 0.152939
R12497 GND.n938 GND.n933 0.152939
R12498 GND.n939 GND.n938 0.152939
R12499 GND.n940 GND.n939 0.152939
R12500 GND.n941 GND.n940 0.152939
R12501 GND.n946 GND.n941 0.152939
R12502 GND.n947 GND.n946 0.152939
R12503 GND.n948 GND.n947 0.152939
R12504 GND.n949 GND.n948 0.152939
R12505 GND.n954 GND.n949 0.152939
R12506 GND.n955 GND.n954 0.152939
R12507 GND.n956 GND.n955 0.152939
R12508 GND.n957 GND.n956 0.152939
R12509 GND.n962 GND.n957 0.152939
R12510 GND.n963 GND.n962 0.152939
R12511 GND.n964 GND.n963 0.152939
R12512 GND.n965 GND.n964 0.152939
R12513 GND.n970 GND.n965 0.152939
R12514 GND.n971 GND.n970 0.152939
R12515 GND.n972 GND.n971 0.152939
R12516 GND.n973 GND.n972 0.152939
R12517 GND.n978 GND.n973 0.152939
R12518 GND.n979 GND.n978 0.152939
R12519 GND.n980 GND.n979 0.152939
R12520 GND.n981 GND.n980 0.152939
R12521 GND.n986 GND.n981 0.152939
R12522 GND.n987 GND.n986 0.152939
R12523 GND.n988 GND.n987 0.152939
R12524 GND.n989 GND.n988 0.152939
R12525 GND.n994 GND.n989 0.152939
R12526 GND.n995 GND.n994 0.152939
R12527 GND.n996 GND.n995 0.152939
R12528 GND.n997 GND.n996 0.152939
R12529 GND.n1002 GND.n997 0.152939
R12530 GND.n1003 GND.n1002 0.152939
R12531 GND.n6404 GND.n1003 0.152939
R12532 GND.n6850 GND.n541 0.152939
R12533 GND.n568 GND.n541 0.152939
R12534 GND.n569 GND.n568 0.152939
R12535 GND.n570 GND.n569 0.152939
R12536 GND.n588 GND.n570 0.152939
R12537 GND.n589 GND.n588 0.152939
R12538 GND.n590 GND.n589 0.152939
R12539 GND.n591 GND.n590 0.152939
R12540 GND.n608 GND.n591 0.152939
R12541 GND.n609 GND.n608 0.152939
R12542 GND.n610 GND.n609 0.152939
R12543 GND.n611 GND.n610 0.152939
R12544 GND.n629 GND.n611 0.152939
R12545 GND.n630 GND.n629 0.152939
R12546 GND.n631 GND.n630 0.152939
R12547 GND.n632 GND.n631 0.152939
R12548 GND.n649 GND.n632 0.152939
R12549 GND.n6790 GND.n649 0.152939
R12550 GND.n4103 GND.n4102 0.152939
R12551 GND.n4279 GND.n4102 0.152939
R12552 GND.n4280 GND.n4279 0.152939
R12553 GND.n4281 GND.n4280 0.152939
R12554 GND.n4281 GND.n4100 0.152939
R12555 GND.n4303 GND.n4100 0.152939
R12556 GND.n4304 GND.n4303 0.152939
R12557 GND.n4305 GND.n4304 0.152939
R12558 GND.n4305 GND.n4096 0.152939
R12559 GND.n4318 GND.n4096 0.152939
R12560 GND.n4319 GND.n4318 0.152939
R12561 GND.n4320 GND.n4319 0.152939
R12562 GND.n4320 GND.n4092 0.152939
R12563 GND.n4333 GND.n4092 0.152939
R12564 GND.n4334 GND.n4333 0.152939
R12565 GND.n4335 GND.n4334 0.152939
R12566 GND.n4336 GND.n4335 0.152939
R12567 GND.n4337 GND.n4336 0.152939
R12568 GND.n4338 GND.n4337 0.152939
R12569 GND.n4339 GND.n4338 0.152939
R12570 GND.n4340 GND.n4339 0.152939
R12571 GND.n4340 GND.n527 0.152939
R12572 GND.n4407 GND.n528 0.152939
R12573 GND.n4408 GND.n4407 0.152939
R12574 GND.n4409 GND.n4408 0.152939
R12575 GND.n4414 GND.n4409 0.152939
R12576 GND.n4415 GND.n4414 0.152939
R12577 GND.n4416 GND.n4415 0.152939
R12578 GND.n4417 GND.n4416 0.152939
R12579 GND.n4420 GND.n4417 0.152939
R12580 GND.n4421 GND.n4420 0.152939
R12581 GND.n4422 GND.n4421 0.152939
R12582 GND.n4423 GND.n4422 0.152939
R12583 GND.n4423 GND.n792 0.152939
R12584 GND.n6621 GND.n792 0.152939
R12585 GND.n6622 GND.n6621 0.152939
R12586 GND.n6623 GND.n6622 0.152939
R12587 GND.n6623 GND.n787 0.152939
R12588 GND.n6635 GND.n787 0.152939
R12589 GND.n6636 GND.n6635 0.152939
R12590 GND.n6638 GND.n6636 0.152939
R12591 GND.n6638 GND.n6637 0.152939
R12592 GND.n6637 GND.n782 0.152939
R12593 GND.n6652 GND.n782 0.152939
R12594 GND.n6673 GND.n760 0.152939
R12595 GND.n763 GND.n760 0.152939
R12596 GND.n767 GND.n763 0.152939
R12597 GND.n768 GND.n767 0.152939
R12598 GND.n769 GND.n768 0.152939
R12599 GND.n770 GND.n769 0.152939
R12600 GND.n771 GND.n770 0.152939
R12601 GND.n775 GND.n771 0.152939
R12602 GND.n776 GND.n775 0.152939
R12603 GND.n6654 GND.n776 0.152939
R12604 GND.n6654 GND.n6653 0.152939
R12605 GND.n6789 GND.n650 0.152939
R12606 GND.n652 GND.n650 0.152939
R12607 GND.n657 GND.n652 0.152939
R12608 GND.n658 GND.n657 0.152939
R12609 GND.n659 GND.n658 0.152939
R12610 GND.n660 GND.n659 0.152939
R12611 GND.n664 GND.n660 0.152939
R12612 GND.n665 GND.n664 0.152939
R12613 GND.n666 GND.n665 0.152939
R12614 GND.n6771 GND.n666 0.152939
R12615 GND.n6771 GND.n6770 0.152939
R12616 GND.n6770 GND.n6769 0.152939
R12617 GND.n6769 GND.n672 0.152939
R12618 GND.n677 GND.n672 0.152939
R12619 GND.n678 GND.n677 0.152939
R12620 GND.n679 GND.n678 0.152939
R12621 GND.n683 GND.n679 0.152939
R12622 GND.n684 GND.n683 0.152939
R12623 GND.n685 GND.n684 0.152939
R12624 GND.n686 GND.n685 0.152939
R12625 GND.n693 GND.n686 0.152939
R12626 GND.n6748 GND.n693 0.152939
R12627 GND.n6748 GND.n6747 0.152939
R12628 GND.n6747 GND.n6746 0.152939
R12629 GND.n6746 GND.n694 0.152939
R12630 GND.n698 GND.n694 0.152939
R12631 GND.n699 GND.n698 0.152939
R12632 GND.n700 GND.n699 0.152939
R12633 GND.n704 GND.n700 0.152939
R12634 GND.n705 GND.n704 0.152939
R12635 GND.n706 GND.n705 0.152939
R12636 GND.n707 GND.n706 0.152939
R12637 GND.n711 GND.n707 0.152939
R12638 GND.n712 GND.n711 0.152939
R12639 GND.n713 GND.n712 0.152939
R12640 GND.n714 GND.n713 0.152939
R12641 GND.n718 GND.n714 0.152939
R12642 GND.n719 GND.n718 0.152939
R12643 GND.n720 GND.n719 0.152939
R12644 GND.n721 GND.n720 0.152939
R12645 GND.n725 GND.n721 0.152939
R12646 GND.n726 GND.n725 0.152939
R12647 GND.n727 GND.n726 0.152939
R12648 GND.n728 GND.n727 0.152939
R12649 GND.n732 GND.n728 0.152939
R12650 GND.n733 GND.n732 0.152939
R12651 GND.n734 GND.n733 0.152939
R12652 GND.n735 GND.n734 0.152939
R12653 GND.n739 GND.n735 0.152939
R12654 GND.n740 GND.n739 0.152939
R12655 GND.n741 GND.n740 0.152939
R12656 GND.n742 GND.n741 0.152939
R12657 GND.n746 GND.n742 0.152939
R12658 GND.n747 GND.n746 0.152939
R12659 GND.n748 GND.n747 0.152939
R12660 GND.n749 GND.n748 0.152939
R12661 GND.n753 GND.n749 0.152939
R12662 GND.n754 GND.n753 0.152939
R12663 GND.n6676 GND.n754 0.152939
R12664 GND.n6676 GND.n6675 0.152939
R12665 GND.n4550 GND.n4549 0.152939
R12666 GND.n4551 GND.n4550 0.152939
R12667 GND.n4552 GND.n4551 0.152939
R12668 GND.n4553 GND.n4552 0.152939
R12669 GND.n4554 GND.n4553 0.152939
R12670 GND.n4555 GND.n4554 0.152939
R12671 GND.n4556 GND.n4555 0.152939
R12672 GND.n4557 GND.n4556 0.152939
R12673 GND.n4558 GND.n4557 0.152939
R12674 GND.n4560 GND.n4558 0.152939
R12675 GND.n4563 GND.n4560 0.152939
R12676 GND.n4564 GND.n4563 0.152939
R12677 GND.n4565 GND.n4564 0.152939
R12678 GND.n4566 GND.n4565 0.152939
R12679 GND.n4567 GND.n4566 0.152939
R12680 GND.n4568 GND.n4567 0.152939
R12681 GND.n4569 GND.n4568 0.152939
R12682 GND.n4570 GND.n4569 0.152939
R12683 GND.n4571 GND.n4570 0.152939
R12684 GND.n4572 GND.n4571 0.152939
R12685 GND.n4573 GND.n4572 0.152939
R12686 GND.n4575 GND.n4573 0.152939
R12687 GND.n4578 GND.n4575 0.152939
R12688 GND.n4579 GND.n4578 0.152939
R12689 GND.n4581 GND.n4579 0.152939
R12690 GND.n4581 GND.n4580 0.152939
R12691 GND.n4154 GND.n3884 0.152939
R12692 GND.n4155 GND.n4154 0.152939
R12693 GND.n4156 GND.n4155 0.152939
R12694 GND.n4156 GND.n4151 0.152939
R12695 GND.n4167 GND.n4151 0.152939
R12696 GND.n4168 GND.n4167 0.152939
R12697 GND.n4169 GND.n4168 0.152939
R12698 GND.n4169 GND.n4149 0.152939
R12699 GND.n4177 GND.n4149 0.152939
R12700 GND.n4178 GND.n4177 0.152939
R12701 GND.n4179 GND.n4178 0.152939
R12702 GND.n4179 GND.n4147 0.152939
R12703 GND.n4187 GND.n4147 0.152939
R12704 GND.n4188 GND.n4187 0.152939
R12705 GND.n4189 GND.n4188 0.152939
R12706 GND.n4189 GND.n4145 0.152939
R12707 GND.n4200 GND.n4145 0.152939
R12708 GND.n4201 GND.n4200 0.152939
R12709 GND.n4202 GND.n4201 0.152939
R12710 GND.n4202 GND.n4143 0.152939
R12711 GND.n4210 GND.n4143 0.152939
R12712 GND.n4211 GND.n4210 0.152939
R12713 GND.n4212 GND.n4211 0.152939
R12714 GND.n4212 GND.n4141 0.152939
R12715 GND.n4220 GND.n4141 0.152939
R12716 GND.n4221 GND.n4220 0.152939
R12717 GND.n4222 GND.n4221 0.152939
R12718 GND.n4222 GND.n4139 0.152939
R12719 GND.n4230 GND.n4139 0.152939
R12720 GND.n4231 GND.n4230 0.152939
R12721 GND.n4270 GND.n4231 0.152939
R12722 GND.n4548 GND.n3927 0.152939
R12723 GND.n3962 GND.n3927 0.152939
R12724 GND.n3965 GND.n3962 0.152939
R12725 GND.n3966 GND.n3965 0.152939
R12726 GND.n3967 GND.n3966 0.152939
R12727 GND.n3968 GND.n3967 0.152939
R12728 GND.n3969 GND.n3968 0.152939
R12729 GND.n3989 GND.n3969 0.152939
R12730 GND.n3990 GND.n3989 0.152939
R12731 GND.n3991 GND.n3990 0.152939
R12732 GND.n3992 GND.n3991 0.152939
R12733 GND.n4010 GND.n3992 0.152939
R12734 GND.n4011 GND.n4010 0.152939
R12735 GND.n4012 GND.n4011 0.152939
R12736 GND.n4013 GND.n4012 0.152939
R12737 GND.n4014 GND.n4013 0.152939
R12738 GND.n4014 GND.n542 0.152939
R12739 GND.n6850 GND.n542 0.152939
R12740 GND.n2706 GND.n2703 0.152939
R12741 GND.n2707 GND.n2706 0.152939
R12742 GND.n2708 GND.n2707 0.152939
R12743 GND.n2709 GND.n2708 0.152939
R12744 GND.n2714 GND.n2709 0.152939
R12745 GND.n2715 GND.n2714 0.152939
R12746 GND.n2716 GND.n2715 0.152939
R12747 GND.n2717 GND.n2716 0.152939
R12748 GND.n2719 GND.n2717 0.152939
R12749 GND.n2719 GND.n2718 0.152939
R12750 GND.n2718 GND.n2092 0.152939
R12751 GND.n2828 GND.n2092 0.152939
R12752 GND.n2829 GND.n2828 0.152939
R12753 GND.n2830 GND.n2829 0.152939
R12754 GND.n2832 GND.n2830 0.152939
R12755 GND.n2832 GND.n2831 0.152939
R12756 GND.n2831 GND.n2062 0.152939
R12757 GND.n2914 GND.n2062 0.152939
R12758 GND.n2915 GND.n2914 0.152939
R12759 GND.n2916 GND.n2915 0.152939
R12760 GND.n2917 GND.n2916 0.152939
R12761 GND.n2918 GND.n2917 0.152939
R12762 GND.n2923 GND.n2918 0.152939
R12763 GND.n2924 GND.n2923 0.152939
R12764 GND.n2925 GND.n2924 0.152939
R12765 GND.n2926 GND.n2925 0.152939
R12766 GND.n2941 GND.n2926 0.152939
R12767 GND.n2942 GND.n2941 0.152939
R12768 GND.n2943 GND.n2942 0.152939
R12769 GND.n2944 GND.n2943 0.152939
R12770 GND.n3546 GND.n2944 0.152939
R12771 GND.n3547 GND.n3546 0.152939
R12772 GND.n3549 GND.n3547 0.152939
R12773 GND.n3549 GND.n3548 0.152939
R12774 GND.n3548 GND.n3001 0.152939
R12775 GND.n3002 GND.n3001 0.152939
R12776 GND.n3003 GND.n3002 0.152939
R12777 GND.n3041 GND.n3003 0.152939
R12778 GND.n3044 GND.n3041 0.152939
R12779 GND.n3045 GND.n3044 0.152939
R12780 GND.n3046 GND.n3045 0.152939
R12781 GND.n3047 GND.n3046 0.152939
R12782 GND.n3048 GND.n3047 0.152939
R12783 GND.n3085 GND.n3048 0.152939
R12784 GND.n3088 GND.n3085 0.152939
R12785 GND.n3089 GND.n3088 0.152939
R12786 GND.n3090 GND.n3089 0.152939
R12787 GND.n3091 GND.n3090 0.152939
R12788 GND.n3092 GND.n3091 0.152939
R12789 GND.n3135 GND.n3092 0.152939
R12790 GND.n3136 GND.n3135 0.152939
R12791 GND.n3141 GND.n3136 0.152939
R12792 GND.n3142 GND.n3141 0.152939
R12793 GND.n3143 GND.n3142 0.152939
R12794 GND.n3144 GND.n3143 0.152939
R12795 GND.n3145 GND.n3144 0.152939
R12796 GND.n3330 GND.n3145 0.152939
R12797 GND.n3331 GND.n3330 0.152939
R12798 GND.n3331 GND.n3328 0.152939
R12799 GND.n3337 GND.n3328 0.152939
R12800 GND.n3338 GND.n3337 0.152939
R12801 GND.n3339 GND.n3338 0.152939
R12802 GND.n3339 GND.n3324 0.152939
R12803 GND.n3741 GND.n3324 0.152939
R12804 GND.n3742 GND.n3741 0.152939
R12805 GND.n3743 GND.n3742 0.152939
R12806 GND.n3745 GND.n3743 0.152939
R12807 GND.n3745 GND.n3744 0.152939
R12808 GND.n3744 GND.n3219 0.152939
R12809 GND.n3220 GND.n3219 0.152939
R12810 GND.n3221 GND.n3220 0.152939
R12811 GND.n3236 GND.n3221 0.152939
R12812 GND.n3237 GND.n3236 0.152939
R12813 GND.n3238 GND.n3237 0.152939
R12814 GND.n3239 GND.n3238 0.152939
R12815 GND.n4114 GND.n3239 0.152939
R12816 GND.n4115 GND.n4114 0.152939
R12817 GND.n4116 GND.n4115 0.152939
R12818 GND.n4117 GND.n4116 0.152939
R12819 GND.n4117 GND.n4108 0.152939
R12820 GND.n4127 GND.n4108 0.152939
R12821 GND.n4128 GND.n4127 0.152939
R12822 GND.n4129 GND.n4128 0.152939
R12823 GND.n4131 GND.n4129 0.152939
R12824 GND.n4131 GND.n4130 0.152939
R12825 GND.n4130 GND.n3948 0.152939
R12826 GND.n3949 GND.n3948 0.152939
R12827 GND.n3950 GND.n3949 0.152939
R12828 GND.n4066 GND.n3950 0.152939
R12829 GND.n4067 GND.n4066 0.152939
R12830 GND.n4068 GND.n4067 0.152939
R12831 GND.n4068 GND.n4062 0.152939
R12832 GND.n4074 GND.n4062 0.152939
R12833 GND.n4075 GND.n4074 0.152939
R12834 GND.n4076 GND.n4075 0.152939
R12835 GND.n4076 GND.n4058 0.152939
R12836 GND.n4082 GND.n4058 0.152939
R12837 GND.n4083 GND.n4082 0.152939
R12838 GND.n4084 GND.n4083 0.152939
R12839 GND.n4086 GND.n4084 0.152939
R12840 GND.n4086 GND.n4085 0.152939
R12841 GND.n2768 GND.n2767 0.152939
R12842 GND.n2769 GND.n2768 0.152939
R12843 GND.n2769 GND.n2120 0.152939
R12844 GND.n2791 GND.n2120 0.152939
R12845 GND.n2792 GND.n2791 0.152939
R12846 GND.n2793 GND.n2792 0.152939
R12847 GND.n2794 GND.n2793 0.152939
R12848 GND.n2794 GND.n2099 0.152939
R12849 GND.n2817 GND.n2099 0.152939
R12850 GND.n2818 GND.n2817 0.152939
R12851 GND.n2819 GND.n2818 0.152939
R12852 GND.n2819 GND.n2075 0.152939
R12853 GND.n2897 GND.n2075 0.152939
R12854 GND.n2898 GND.n2897 0.152939
R12855 GND.n2899 GND.n2898 0.152939
R12856 GND.n2900 GND.n2899 0.152939
R12857 GND.n2900 GND.n1993 0.152939
R12858 GND.n5053 GND.n1993 0.152939
R12859 GND.n2345 GND.n2344 0.152939
R12860 GND.n2346 GND.n2345 0.152939
R12861 GND.n2346 GND.n2338 0.152939
R12862 GND.n2354 GND.n2338 0.152939
R12863 GND.n2355 GND.n2354 0.152939
R12864 GND.n2356 GND.n2355 0.152939
R12865 GND.n2356 GND.n2334 0.152939
R12866 GND.n2364 GND.n2334 0.152939
R12867 GND.n2365 GND.n2364 0.152939
R12868 GND.n2366 GND.n2365 0.152939
R12869 GND.n2366 GND.n2330 0.152939
R12870 GND.n2376 GND.n2330 0.152939
R12871 GND.n2377 GND.n2376 0.152939
R12872 GND.n2378 GND.n2377 0.152939
R12873 GND.n2378 GND.n2326 0.152939
R12874 GND.n2386 GND.n2326 0.152939
R12875 GND.n2387 GND.n2386 0.152939
R12876 GND.n2388 GND.n2387 0.152939
R12877 GND.n2388 GND.n2322 0.152939
R12878 GND.n2396 GND.n2322 0.152939
R12879 GND.n2397 GND.n2396 0.152939
R12880 GND.n2398 GND.n2397 0.152939
R12881 GND.n2398 GND.n2318 0.152939
R12882 GND.n2408 GND.n2318 0.152939
R12883 GND.n2409 GND.n2408 0.152939
R12884 GND.n2410 GND.n2409 0.152939
R12885 GND.n2410 GND.n2314 0.152939
R12886 GND.n2418 GND.n2314 0.152939
R12887 GND.n2419 GND.n2418 0.152939
R12888 GND.n2420 GND.n2419 0.152939
R12889 GND.n2420 GND.n2310 0.152939
R12890 GND.n2428 GND.n2310 0.152939
R12891 GND.n2429 GND.n2428 0.152939
R12892 GND.n2430 GND.n2429 0.152939
R12893 GND.n2430 GND.n2306 0.152939
R12894 GND.n2441 GND.n2306 0.152939
R12895 GND.n2442 GND.n2441 0.152939
R12896 GND.n2443 GND.n2442 0.152939
R12897 GND.n2443 GND.n2302 0.152939
R12898 GND.n2451 GND.n2302 0.152939
R12899 GND.n2452 GND.n2451 0.152939
R12900 GND.n2453 GND.n2452 0.152939
R12901 GND.n2453 GND.n2298 0.152939
R12902 GND.n2461 GND.n2298 0.152939
R12903 GND.n2462 GND.n2461 0.152939
R12904 GND.n2463 GND.n2462 0.152939
R12905 GND.n2463 GND.n2294 0.152939
R12906 GND.n2474 GND.n2294 0.152939
R12907 GND.n2475 GND.n2474 0.152939
R12908 GND.n2476 GND.n2475 0.152939
R12909 GND.n2476 GND.n2290 0.152939
R12910 GND.n2484 GND.n2290 0.152939
R12911 GND.n2485 GND.n2484 0.152939
R12912 GND.n2486 GND.n2485 0.152939
R12913 GND.n2486 GND.n2286 0.152939
R12914 GND.n2494 GND.n2286 0.152939
R12915 GND.n2495 GND.n2494 0.152939
R12916 GND.n2496 GND.n2495 0.152939
R12917 GND.n2496 GND.n2280 0.152939
R12918 GND.n2503 GND.n2280 0.152939
R12919 GND.n1882 GND.n1881 0.152939
R12920 GND.n1883 GND.n1882 0.152939
R12921 GND.n2260 GND.n1883 0.152939
R12922 GND.n2593 GND.n2260 0.152939
R12923 GND.n2594 GND.n2593 0.152939
R12924 GND.n2595 GND.n2594 0.152939
R12925 GND.n2596 GND.n2595 0.152939
R12926 GND.n2596 GND.n2237 0.152939
R12927 GND.n2617 GND.n2237 0.152939
R12928 GND.n2618 GND.n2617 0.152939
R12929 GND.n2619 GND.n2618 0.152939
R12930 GND.n2620 GND.n2619 0.152939
R12931 GND.n2620 GND.n2203 0.152939
R12932 GND.n2667 GND.n2203 0.152939
R12933 GND.n2668 GND.n2667 0.152939
R12934 GND.n2669 GND.n2668 0.152939
R12935 GND.n2669 GND.n2141 0.152939
R12936 GND.n2767 GND.n2141 0.152939
R12937 GND.n5324 GND.n1686 0.152939
R12938 GND.n1692 GND.n1686 0.152939
R12939 GND.n1693 GND.n1692 0.152939
R12940 GND.n1694 GND.n1693 0.152939
R12941 GND.n1695 GND.n1694 0.152939
R12942 GND.n1700 GND.n1695 0.152939
R12943 GND.n1701 GND.n1700 0.152939
R12944 GND.n1702 GND.n1701 0.152939
R12945 GND.n1703 GND.n1702 0.152939
R12946 GND.n1708 GND.n1703 0.152939
R12947 GND.n1709 GND.n1708 0.152939
R12948 GND.n1710 GND.n1709 0.152939
R12949 GND.n1711 GND.n1710 0.152939
R12950 GND.n1716 GND.n1711 0.152939
R12951 GND.n1717 GND.n1716 0.152939
R12952 GND.n1718 GND.n1717 0.152939
R12953 GND.n1719 GND.n1718 0.152939
R12954 GND.n1724 GND.n1719 0.152939
R12955 GND.n1725 GND.n1724 0.152939
R12956 GND.n1726 GND.n1725 0.152939
R12957 GND.n1727 GND.n1726 0.152939
R12958 GND.n1732 GND.n1727 0.152939
R12959 GND.n1733 GND.n1732 0.152939
R12960 GND.n1734 GND.n1733 0.152939
R12961 GND.n1735 GND.n1734 0.152939
R12962 GND.n1740 GND.n1735 0.152939
R12963 GND.n1741 GND.n1740 0.152939
R12964 GND.n1742 GND.n1741 0.152939
R12965 GND.n1743 GND.n1742 0.152939
R12966 GND.n1748 GND.n1743 0.152939
R12967 GND.n1749 GND.n1748 0.152939
R12968 GND.n1750 GND.n1749 0.152939
R12969 GND.n1751 GND.n1750 0.152939
R12970 GND.n1756 GND.n1751 0.152939
R12971 GND.n1757 GND.n1756 0.152939
R12972 GND.n1758 GND.n1757 0.152939
R12973 GND.n1759 GND.n1758 0.152939
R12974 GND.n1764 GND.n1759 0.152939
R12975 GND.n1765 GND.n1764 0.152939
R12976 GND.n1766 GND.n1765 0.152939
R12977 GND.n1767 GND.n1766 0.152939
R12978 GND.n1772 GND.n1767 0.152939
R12979 GND.n1773 GND.n1772 0.152939
R12980 GND.n1774 GND.n1773 0.152939
R12981 GND.n1775 GND.n1774 0.152939
R12982 GND.n1780 GND.n1775 0.152939
R12983 GND.n1781 GND.n1780 0.152939
R12984 GND.n1782 GND.n1781 0.152939
R12985 GND.n1783 GND.n1782 0.152939
R12986 GND.n1788 GND.n1783 0.152939
R12987 GND.n1789 GND.n1788 0.152939
R12988 GND.n1790 GND.n1789 0.152939
R12989 GND.n1791 GND.n1790 0.152939
R12990 GND.n1796 GND.n1791 0.152939
R12991 GND.n1797 GND.n1796 0.152939
R12992 GND.n1798 GND.n1797 0.152939
R12993 GND.n1799 GND.n1798 0.152939
R12994 GND.n1804 GND.n1799 0.152939
R12995 GND.n1805 GND.n1804 0.152939
R12996 GND.n1806 GND.n1805 0.152939
R12997 GND.n1807 GND.n1806 0.152939
R12998 GND.n1812 GND.n1807 0.152939
R12999 GND.n1813 GND.n1812 0.152939
R13000 GND.n1814 GND.n1813 0.152939
R13001 GND.n1815 GND.n1814 0.152939
R13002 GND.n1820 GND.n1815 0.152939
R13003 GND.n1821 GND.n1820 0.152939
R13004 GND.n1822 GND.n1821 0.152939
R13005 GND.n1823 GND.n1822 0.152939
R13006 GND.n1828 GND.n1823 0.152939
R13007 GND.n1829 GND.n1828 0.152939
R13008 GND.n1830 GND.n1829 0.152939
R13009 GND.n1831 GND.n1830 0.152939
R13010 GND.n1836 GND.n1831 0.152939
R13011 GND.n1837 GND.n1836 0.152939
R13012 GND.n1838 GND.n1837 0.152939
R13013 GND.n1839 GND.n1838 0.152939
R13014 GND.n1844 GND.n1839 0.152939
R13015 GND.n1845 GND.n1844 0.152939
R13016 GND.n1846 GND.n1845 0.152939
R13017 GND.n1847 GND.n1846 0.152939
R13018 GND.n1852 GND.n1847 0.152939
R13019 GND.n1853 GND.n1852 0.152939
R13020 GND.n1854 GND.n1853 0.152939
R13021 GND.n1855 GND.n1854 0.152939
R13022 GND.n1860 GND.n1855 0.152939
R13023 GND.n1861 GND.n1860 0.152939
R13024 GND.n1862 GND.n1861 0.152939
R13025 GND.n1863 GND.n1862 0.152939
R13026 GND.n1868 GND.n1863 0.152939
R13027 GND.n1869 GND.n1868 0.152939
R13028 GND.n1870 GND.n1869 0.152939
R13029 GND.n1871 GND.n1870 0.152939
R13030 GND.n2554 GND.n1871 0.152939
R13031 GND.n2555 GND.n2554 0.152939
R13032 GND.n2555 GND.n2552 0.152939
R13033 GND.n2561 GND.n2552 0.152939
R13034 GND.n2562 GND.n2561 0.152939
R13035 GND.n2563 GND.n2562 0.152939
R13036 GND.n2564 GND.n2563 0.152939
R13037 GND.n2565 GND.n2564 0.152939
R13038 GND.n2568 GND.n2565 0.152939
R13039 GND.n2569 GND.n2568 0.152939
R13040 GND.n2570 GND.n2569 0.152939
R13041 GND.n2571 GND.n2570 0.152939
R13042 GND.n2572 GND.n2571 0.152939
R13043 GND.n2572 GND.n2218 0.152939
R13044 GND.n2640 GND.n2218 0.152939
R13045 GND.n2641 GND.n2640 0.152939
R13046 GND.n2642 GND.n2641 0.152939
R13047 GND.n2643 GND.n2642 0.152939
R13048 GND.n2644 GND.n2643 0.152939
R13049 GND.n1598 GND.n1597 0.152939
R13050 GND.n1599 GND.n1598 0.152939
R13051 GND.n1604 GND.n1599 0.152939
R13052 GND.n1605 GND.n1604 0.152939
R13053 GND.n1606 GND.n1605 0.152939
R13054 GND.n1607 GND.n1606 0.152939
R13055 GND.n1612 GND.n1607 0.152939
R13056 GND.n1613 GND.n1612 0.152939
R13057 GND.n1614 GND.n1613 0.152939
R13058 GND.n1615 GND.n1614 0.152939
R13059 GND.n1620 GND.n1615 0.152939
R13060 GND.n1621 GND.n1620 0.152939
R13061 GND.n1622 GND.n1621 0.152939
R13062 GND.n1623 GND.n1622 0.152939
R13063 GND.n1628 GND.n1623 0.152939
R13064 GND.n1629 GND.n1628 0.152939
R13065 GND.n1630 GND.n1629 0.152939
R13066 GND.n1631 GND.n1630 0.152939
R13067 GND.n1636 GND.n1631 0.152939
R13068 GND.n1637 GND.n1636 0.152939
R13069 GND.n1638 GND.n1637 0.152939
R13070 GND.n1639 GND.n1638 0.152939
R13071 GND.n1644 GND.n1639 0.152939
R13072 GND.n1645 GND.n1644 0.152939
R13073 GND.n1646 GND.n1645 0.152939
R13074 GND.n1647 GND.n1646 0.152939
R13075 GND.n1652 GND.n1647 0.152939
R13076 GND.n1653 GND.n1652 0.152939
R13077 GND.n1654 GND.n1653 0.152939
R13078 GND.n1655 GND.n1654 0.152939
R13079 GND.n1660 GND.n1655 0.152939
R13080 GND.n1661 GND.n1660 0.152939
R13081 GND.n1662 GND.n1661 0.152939
R13082 GND.n1663 GND.n1662 0.152939
R13083 GND.n1668 GND.n1663 0.152939
R13084 GND.n1669 GND.n1668 0.152939
R13085 GND.n1670 GND.n1669 0.152939
R13086 GND.n1671 GND.n1670 0.152939
R13087 GND.n1676 GND.n1671 0.152939
R13088 GND.n1677 GND.n1676 0.152939
R13089 GND.n1678 GND.n1677 0.152939
R13090 GND.n1679 GND.n1678 0.152939
R13091 GND.n1684 GND.n1679 0.152939
R13092 GND.n1685 GND.n1684 0.152939
R13093 GND.n5325 GND.n1685 0.152939
R13094 GND.n2688 GND.n2185 0.152939
R13095 GND.n2689 GND.n2688 0.152939
R13096 GND.n2690 GND.n2689 0.152939
R13097 GND.n2690 GND.n2131 0.152939
R13098 GND.n2776 GND.n2131 0.152939
R13099 GND.n2777 GND.n2776 0.152939
R13100 GND.n2779 GND.n2777 0.152939
R13101 GND.n2779 GND.n2778 0.152939
R13102 GND.n2778 GND.n2111 0.152939
R13103 GND.n2801 GND.n2111 0.152939
R13104 GND.n2802 GND.n2801 0.152939
R13105 GND.n2807 GND.n2802 0.152939
R13106 GND.n2807 GND.n2806 0.152939
R13107 GND.n2806 GND.n2805 0.152939
R13108 GND.n2805 GND.n2088 0.152939
R13109 GND.n2888 GND.n2088 0.152939
R13110 GND.n2888 GND.n2887 0.152939
R13111 GND.n2887 GND.n2886 0.152939
R13112 GND.n2886 GND.n2089 0.152939
R13113 GND.n2882 GND.n2089 0.152939
R13114 GND.n2882 GND.n2881 0.152939
R13115 GND.n2881 GND.n2880 0.152939
R13116 GND.n5052 GND.n1994 0.152939
R13117 GND.n5048 GND.n1994 0.152939
R13118 GND.n5048 GND.n5047 0.152939
R13119 GND.n5047 GND.n5046 0.152939
R13120 GND.n5046 GND.n1998 0.152939
R13121 GND.n5042 GND.n1998 0.152939
R13122 GND.n5042 GND.n5041 0.152939
R13123 GND.n5041 GND.n5040 0.152939
R13124 GND.n5040 GND.n2003 0.152939
R13125 GND.n2008 GND.n2003 0.152939
R13126 GND.n5035 GND.n2008 0.152939
R13127 GND.n5035 GND.n5034 0.152939
R13128 GND.n5034 GND.n5033 0.152939
R13129 GND.n5033 GND.n2012 0.152939
R13130 GND.n5029 GND.n2012 0.152939
R13131 GND.n5029 GND.n5028 0.152939
R13132 GND.n5028 GND.n5027 0.152939
R13133 GND.n5027 GND.n2017 0.152939
R13134 GND.n5023 GND.n2017 0.152939
R13135 GND.n5023 GND.n5022 0.152939
R13136 GND.n5022 GND.n5021 0.152939
R13137 GND.n5021 GND.n2022 0.152939
R13138 GND.n5017 GND.n2022 0.152939
R13139 GND.n5017 GND.n5016 0.152939
R13140 GND.n5016 GND.n5015 0.152939
R13141 GND.n5015 GND.n2029 0.152939
R13142 GND.n5004 GND.n4893 0.152939
R13143 GND.n5004 GND.n5003 0.152939
R13144 GND.n5003 GND.n5002 0.152939
R13145 GND.n5002 GND.n4894 0.152939
R13146 GND.n4998 GND.n4894 0.152939
R13147 GND.n4998 GND.n4997 0.152939
R13148 GND.n4997 GND.n4903 0.152939
R13149 GND.n4993 GND.n4903 0.152939
R13150 GND.n4993 GND.n4992 0.152939
R13151 GND.n4992 GND.n4991 0.152939
R13152 GND.n4991 GND.n4909 0.152939
R13153 GND.n4987 GND.n4909 0.152939
R13154 GND.n4987 GND.n4986 0.152939
R13155 GND.n4986 GND.n4985 0.152939
R13156 GND.n4985 GND.n4917 0.152939
R13157 GND.n4981 GND.n4917 0.152939
R13158 GND.n4981 GND.n4980 0.152939
R13159 GND.n4980 GND.n4979 0.152939
R13160 GND.n4979 GND.n4925 0.152939
R13161 GND.n4975 GND.n4925 0.152939
R13162 GND.n4975 GND.n4974 0.152939
R13163 GND.n4974 GND.n4973 0.152939
R13164 GND.n4973 GND.n4936 0.152939
R13165 GND.n4969 GND.n4936 0.152939
R13166 GND.n4969 GND.n4968 0.152939
R13167 GND.n4968 GND.n4967 0.152939
R13168 GND.n4967 GND.n4944 0.152939
R13169 GND.n4963 GND.n4944 0.152939
R13170 GND.n4963 GND.n4962 0.152939
R13171 GND.n4962 GND.n4961 0.152939
R13172 GND.n4961 GND.n4952 0.152939
R13173 GND.n2509 GND.n2508 0.152939
R13174 GND.n2509 GND.n2276 0.152939
R13175 GND.n2517 GND.n2276 0.152939
R13176 GND.n2518 GND.n2517 0.152939
R13177 GND.n2519 GND.n2518 0.152939
R13178 GND.n2519 GND.n2272 0.152939
R13179 GND.n2527 GND.n2272 0.152939
R13180 GND.n2528 GND.n2527 0.152939
R13181 GND.n2529 GND.n2528 0.152939
R13182 GND.n2529 GND.n2266 0.152939
R13183 GND.n2536 GND.n2266 0.152939
R13184 GND.n2537 GND.n2265 0.152939
R13185 GND.n2544 GND.n2265 0.152939
R13186 GND.n2545 GND.n2544 0.152939
R13187 GND.n2546 GND.n2545 0.152939
R13188 GND.n2546 GND.n2250 0.152939
R13189 GND.n2603 GND.n2250 0.152939
R13190 GND.n2604 GND.n2603 0.152939
R13191 GND.n2606 GND.n2604 0.152939
R13192 GND.n2606 GND.n2605 0.152939
R13193 GND.n2605 GND.n2226 0.152939
R13194 GND.n2627 GND.n2226 0.152939
R13195 GND.n2628 GND.n2627 0.152939
R13196 GND.n2632 GND.n2628 0.152939
R13197 GND.n2632 GND.n2631 0.152939
R13198 GND.n2631 GND.n2630 0.152939
R13199 GND.n2630 GND.n2192 0.152939
R13200 GND.n2676 GND.n2192 0.152939
R13201 GND.n2677 GND.n2676 0.152939
R13202 GND.n2678 GND.n2677 0.152939
R13203 GND.n2678 GND.n2189 0.152939
R13204 GND.n2682 GND.n2189 0.152939
R13205 GND.n2683 GND.n2682 0.152939
R13206 GND.n6858 GND.n527 0.145814
R13207 GND.n6858 GND.n528 0.145814
R13208 GND.n2684 GND.n2185 0.145814
R13209 GND.n2684 GND.n2683 0.145814
R13210 GND.n4383 GND.n543 0.0858659
R13211 GND.n2644 GND.n2142 0.0858659
R13212 GND.n4269 GND.n4268 0.0756008
R13213 GND.n2848 GND.n1983 0.0756008
R13214 GND.n2703 GND.n2142 0.0675732
R13215 GND.n4085 GND.n543 0.0675732
R13216 GND.n4269 GND.n3938 0.0436386
R13217 GND.n6674 GND.n642 0.0436386
R13218 GND.n2507 GND.n2506 0.0436386
R13219 GND.n5059 GND.n1983 0.0436386
R13220 GND.n4541 GND.n3938 0.0344674
R13221 GND.n4541 GND.n3939 0.0344674
R13222 GND.n4290 GND.n3939 0.0344674
R13223 GND.n4290 GND.n4289 0.0344674
R13224 GND.n4296 GND.n4289 0.0344674
R13225 GND.n4297 GND.n4296 0.0344674
R13226 GND.n4297 GND.n3979 0.0344674
R13227 GND.n3980 GND.n3979 0.0344674
R13228 GND.n3981 GND.n3980 0.0344674
R13229 GND.n4312 GND.n3981 0.0344674
R13230 GND.n4312 GND.n4000 0.0344674
R13231 GND.n4001 GND.n4000 0.0344674
R13232 GND.n4002 GND.n4001 0.0344674
R13233 GND.n4327 GND.n4002 0.0344674
R13234 GND.n4327 GND.n4021 0.0344674
R13235 GND.n4022 GND.n4021 0.0344674
R13236 GND.n4023 GND.n4022 0.0344674
R13237 GND.n4354 GND.n4023 0.0344674
R13238 GND.n4355 GND.n4354 0.0344674
R13239 GND.n4355 GND.n4050 0.0344674
R13240 GND.n4051 GND.n4050 0.0344674
R13241 GND.n4052 GND.n4051 0.0344674
R13242 GND.n4360 GND.n4052 0.0344674
R13243 GND.n4361 GND.n4360 0.0344674
R13244 GND.n4366 GND.n4361 0.0344674
R13245 GND.n4367 GND.n4366 0.0344674
R13246 GND.n4412 GND.n4367 0.0344674
R13247 GND.n4412 GND.n558 0.0344674
R13248 GND.n559 GND.n558 0.0344674
R13249 GND.n560 GND.n559 0.0344674
R13250 GND.n4419 GND.n560 0.0344674
R13251 GND.n4419 GND.n578 0.0344674
R13252 GND.n579 GND.n578 0.0344674
R13253 GND.n580 GND.n579 0.0344674
R13254 GND.n795 GND.n580 0.0344674
R13255 GND.n795 GND.n598 0.0344674
R13256 GND.n599 GND.n598 0.0344674
R13257 GND.n600 GND.n599 0.0344674
R13258 GND.n790 GND.n600 0.0344674
R13259 GND.n790 GND.n619 0.0344674
R13260 GND.n620 GND.n619 0.0344674
R13261 GND.n621 GND.n620 0.0344674
R13262 GND.n785 GND.n621 0.0344674
R13263 GND.n785 GND.n640 0.0344674
R13264 GND.n641 GND.n640 0.0344674
R13265 GND.n642 GND.n641 0.0344674
R13266 GND.n2506 GND.n1894 0.0344674
R13267 GND.n5125 GND.n1894 0.0344674
R13268 GND.n5125 GND.n1895 0.0344674
R13269 GND.n5121 GND.n1895 0.0344674
R13270 GND.n5121 GND.n5120 0.0344674
R13271 GND.n5120 GND.n5119 0.0344674
R13272 GND.n5119 GND.n1903 0.0344674
R13273 GND.n5115 GND.n1903 0.0344674
R13274 GND.n5115 GND.n5114 0.0344674
R13275 GND.n5114 GND.n5113 0.0344674
R13276 GND.n5113 GND.n1911 0.0344674
R13277 GND.n5109 GND.n1911 0.0344674
R13278 GND.n5109 GND.n5108 0.0344674
R13279 GND.n5108 GND.n5107 0.0344674
R13280 GND.n5107 GND.n1919 0.0344674
R13281 GND.n5103 GND.n1919 0.0344674
R13282 GND.n5103 GND.n5102 0.0344674
R13283 GND.n5102 GND.n5101 0.0344674
R13284 GND.n5101 GND.n1927 0.0344674
R13285 GND.n5097 GND.n1927 0.0344674
R13286 GND.n5097 GND.n5096 0.0344674
R13287 GND.n5096 GND.n5095 0.0344674
R13288 GND.n5095 GND.n1935 0.0344674
R13289 GND.n5091 GND.n1935 0.0344674
R13290 GND.n5091 GND.n5090 0.0344674
R13291 GND.n5090 GND.n5089 0.0344674
R13292 GND.n5089 GND.n1943 0.0344674
R13293 GND.n5085 GND.n1943 0.0344674
R13294 GND.n5085 GND.n5084 0.0344674
R13295 GND.n5084 GND.n5083 0.0344674
R13296 GND.n5083 GND.n1951 0.0344674
R13297 GND.n5079 GND.n1951 0.0344674
R13298 GND.n5079 GND.n5078 0.0344674
R13299 GND.n5078 GND.n5077 0.0344674
R13300 GND.n5077 GND.n1959 0.0344674
R13301 GND.n5073 GND.n1959 0.0344674
R13302 GND.n5073 GND.n5072 0.0344674
R13303 GND.n5072 GND.n5071 0.0344674
R13304 GND.n5071 GND.n1967 0.0344674
R13305 GND.n5067 GND.n1967 0.0344674
R13306 GND.n5067 GND.n5066 0.0344674
R13307 GND.n5066 GND.n5065 0.0344674
R13308 GND.n5065 GND.n1975 0.0344674
R13309 GND.n5061 GND.n1975 0.0344674
R13310 GND.n5061 GND.n5060 0.0344674
R13311 GND.n5060 GND.n5059 0.0344674
R13312 GND.n4268 GND.n4232 0.0105806
R13313 GND.n4233 GND.n4232 0.0105806
R13314 GND.n4234 GND.n4233 0.0105806
R13315 GND.n4235 GND.n4234 0.0105806
R13316 GND.n4236 GND.n4235 0.0105806
R13317 GND.n4237 GND.n4236 0.0105806
R13318 GND.n4238 GND.n4237 0.0105806
R13319 GND.n4239 GND.n4238 0.0105806
R13320 GND.n4248 GND.n4239 0.0105806
R13321 GND.n4248 GND.n4247 0.0105806
R13322 GND.n4247 GND.n4246 0.0105806
R13323 GND.n2849 GND.n2848 0.0105806
R13324 GND.n2849 GND.n2845 0.0105806
R13325 GND.n2857 GND.n2845 0.0105806
R13326 GND.n2858 GND.n2857 0.0105806
R13327 GND.n2859 GND.n2858 0.0105806
R13328 GND.n2859 GND.n2843 0.0105806
R13329 GND.n2867 GND.n2843 0.0105806
R13330 GND.n2868 GND.n2867 0.0105806
R13331 GND.n2869 GND.n2868 0.0105806
R13332 GND.n2869 GND.n2841 0.0105806
R13333 GND.n2878 GND.n2841 0.0105806
R13334 a_n10279_8682.t5 a_n10279_8682.n9 217.09
R13335 a_n10279_8682.t9 a_n10279_8682.n7 212.185
R13336 a_n10279_8682.t7 a_n10279_8682.n7 217.09
R13337 a_n10279_8682.t3 a_n10279_8682.n9 212.185
R13338 a_n10279_8682.n8 a_n10279_8682.t0 134.072
R13339 a_n10279_8682.n8 a_n10279_8682.t1 100.406
R13340 a_n10279_8682.n1 a_n10279_8682.t25 22.0743
R13341 a_n10279_8682.n1 a_n10279_8682.t29 22.0743
R13342 a_n10279_8682.n2 a_n10279_8682.n6 5.01366
R13343 a_n10279_8682.n2 a_n10279_8682.n5 5.47385
R13344 a_n10279_8682.n0 a_n10279_8682.n8 25.1399
R13345 a_n10279_8682.n0 a_n10279_8682.t4 31.6465
R13346 a_n10279_8682.n0 a_n10279_8682.t10 31.6465
R13347 a_n10279_8682.t8 a_n10279_8682.n6 31.6465
R13348 a_n10279_8682.t11 a_n10279_8682.n5 31.6465
R13349 a_n10279_8682.t27 a_n10279_8682.n1 31.1761
R13350 a_n10279_8682.t22 a_n10279_8682.n1 33.5758
R13351 a_n10279_8682.t18 a_n10279_8682.n1 22.0743
R13352 a_n10279_8682.t13 a_n10279_8682.n4 36.8915
R13353 a_n10279_8682.t26 a_n10279_8682.n1 31.1761
R13354 a_n10279_8682.t20 a_n10279_8682.n1 33.5758
R13355 a_n10279_8682.t12 a_n10279_8682.n1 22.0743
R13356 a_n10279_8682.t15 a_n10279_8682.n3 31.1753
R13357 a_n10279_8682.t21 a_n10279_8682.n1 33.5758
R13358 a_n10279_8682.n1 a_n10279_8682.n7 22.4048
R13359 a_n10279_8682.n9 a_n10279_8682.n1 20.7634
R13360 a_n10279_8682.n4 a_n10279_8682.t19 29.8492
R13361 a_n10279_8682.n1 a_n10279_8682.n2 8.59338
R13362 a_n10279_8682.n0 a_n10279_8682.t2 33.7664
R13363 a_n10279_8682.n0 a_n10279_8682.t14 33.7664
R13364 a_n10279_8682.n6 a_n10279_8682.t6 33.7664
R13365 a_n10279_8682.n5 a_n10279_8682.t24 33.7664
R13366 a_n10279_8682.n1 a_n10279_8682.t28 46.3402
R13367 a_n10279_8682.n1 a_n10279_8682.t17 46.0948
R13368 a_n10279_8682.n1 a_n10279_8682.t23 46.3402
R13369 a_n10279_8682.n3 a_n10279_8682.t16 46.3411
R13370 a_n10279_8682.n1 a_n10279_8682.n0 29.1959
R13371 a_n10279_8682.n1 a_n10279_8682.n3 18.002
R13372 a_n10279_8682.n4 a_n10279_8682.n1 16.0666
R13373 a_n4238_7449.n76 a_n4238_7449.n2 498.942
R13374 a_n4238_7449.n78 a_n4238_7449.n4 498.942
R13375 a_n4238_7449.n64 a_n4238_7449.n6 498.942
R13376 a_n4238_7449.n67 a_n4238_7449.n8 498.942
R13377 a_n4238_7449.n69 a_n4238_7449.n10 498.942
R13378 a_n4238_7449.n73 a_n4238_7449.n12 498.942
R13379 a_n4238_7449.n59 a_n4238_7449.n14 498.942
R13380 a_n4238_7449.n61 a_n4238_7449.n16 498.942
R13381 a_n4238_7449.n1 a_n4238_7449.n2 8.87206
R13382 a_n4238_7449.n76 a_n4238_7449.n20 585
R13383 a_n4238_7449.n36 a_n4238_7449.n35 585
R13384 a_n4238_7449.n3 a_n4238_7449.n4 8.87206
R13385 a_n4238_7449.n78 a_n4238_7449.n22 585
R13386 a_n4238_7449.n39 a_n4238_7449.n38 585
R13387 a_n4238_7449.n5 a_n4238_7449.n6 8.87206
R13388 a_n4238_7449.n64 a_n4238_7449.n24 585
R13389 a_n4238_7449.n42 a_n4238_7449.n41 585
R13390 a_n4238_7449.n7 a_n4238_7449.n8 8.87206
R13391 a_n4238_7449.n67 a_n4238_7449.n26 585
R13392 a_n4238_7449.n45 a_n4238_7449.n44 585
R13393 a_n4238_7449.n9 a_n4238_7449.n10 8.87206
R13394 a_n4238_7449.n69 a_n4238_7449.n28 585
R13395 a_n4238_7449.n48 a_n4238_7449.n47 585
R13396 a_n4238_7449.n11 a_n4238_7449.n12 8.87206
R13397 a_n4238_7449.n73 a_n4238_7449.n30 585
R13398 a_n4238_7449.n51 a_n4238_7449.n50 585
R13399 a_n4238_7449.n13 a_n4238_7449.n14 8.87206
R13400 a_n4238_7449.n59 a_n4238_7449.n32 585
R13401 a_n4238_7449.n54 a_n4238_7449.n53 585
R13402 a_n4238_7449.n15 a_n4238_7449.n16 8.87206
R13403 a_n4238_7449.n61 a_n4238_7449.n34 585
R13404 a_n4238_7449.n57 a_n4238_7449.n56 585
R13405 a_n4238_7449.n76 a_n4238_7449.n35 171.744
R13406 a_n4238_7449.n78 a_n4238_7449.n38 171.744
R13407 a_n4238_7449.n64 a_n4238_7449.n41 171.744
R13408 a_n4238_7449.n67 a_n4238_7449.n44 171.744
R13409 a_n4238_7449.n69 a_n4238_7449.n47 171.744
R13410 a_n4238_7449.n73 a_n4238_7449.n50 171.744
R13411 a_n4238_7449.n59 a_n4238_7449.n53 171.744
R13412 a_n4238_7449.n61 a_n4238_7449.n56 171.744
R13413 a_n4238_7449.n17 a_n4238_7449.n66 115.632
R13414 a_n4238_7449.n72 a_n4238_7449.n71 115.632
R13415 a_n4238_7449.t2 a_n4238_7449.n35 85.8723
R13416 a_n4238_7449.t4 a_n4238_7449.n38 85.8723
R13417 a_n4238_7449.t3 a_n4238_7449.n41 85.8723
R13418 a_n4238_7449.t1 a_n4238_7449.n44 85.8723
R13419 a_n4238_7449.t8 a_n4238_7449.n47 85.8723
R13420 a_n4238_7449.t5 a_n4238_7449.n50 85.8723
R13421 a_n4238_7449.t0 a_n4238_7449.n53 85.8723
R13422 a_n4238_7449.t9 a_n4238_7449.n56 85.8723
R13423 a_n4238_7449.n0 a_n4238_7449.n63 45.9506
R13424 a_n4238_7449.n80 a_n4238_7449.n77 41.5511
R13425 a_n4238_7449.n17 a_n4238_7449.n65 41.5511
R13426 a_n4238_7449.n63 a_n4238_7449.n60 41.5511
R13427 a_n4238_7449.n80 a_n4238_7449.n79 36.646
R13428 a_n4238_7449.n18 a_n4238_7449.n68 36.646
R13429 a_n4238_7449.n18 a_n4238_7449.n70 36.646
R13430 a_n4238_7449.n75 a_n4238_7449.n74 36.646
R13431 a_n4238_7449.n63 a_n4238_7449.n62 36.646
R13432 a_n4238_7449.n0 a_n4238_7449.n80 21.1212
R13433 a_n4238_7449.n37 a_n4238_7449.n36 5.21215
R13434 a_n4238_7449.n40 a_n4238_7449.n39 5.21215
R13435 a_n4238_7449.n43 a_n4238_7449.n42 5.21215
R13436 a_n4238_7449.n46 a_n4238_7449.n45 5.21215
R13437 a_n4238_7449.n49 a_n4238_7449.n48 5.21215
R13438 a_n4238_7449.n52 a_n4238_7449.n51 5.21215
R13439 a_n4238_7449.n55 a_n4238_7449.n54 5.21215
R13440 a_n4238_7449.n58 a_n4238_7449.n57 5.21215
R13441 a_n4238_7449.n20 a_n4238_7449.n36 12.8005
R13442 a_n4238_7449.n22 a_n4238_7449.n39 12.8005
R13443 a_n4238_7449.n24 a_n4238_7449.n42 12.8005
R13444 a_n4238_7449.n26 a_n4238_7449.n45 12.8005
R13445 a_n4238_7449.n28 a_n4238_7449.n48 12.8005
R13446 a_n4238_7449.n30 a_n4238_7449.n51 12.8005
R13447 a_n4238_7449.n32 a_n4238_7449.n54 12.8005
R13448 a_n4238_7449.n34 a_n4238_7449.n57 12.8005
R13449 a_n4238_7449.n66 a_n4238_7449.t11 9.70349
R13450 a_n4238_7449.n66 a_n4238_7449.t6 9.70349
R13451 a_n4238_7449.n71 a_n4238_7449.t10 9.70349
R13452 a_n4238_7449.n71 a_n4238_7449.t7 9.70349
R13453 a_n4238_7449.n58 a_n4238_7449.n33 1.35994
R13454 a_n4238_7449.n77 a_n4238_7449.n19 9.45567
R13455 a_n4238_7449.n79 a_n4238_7449.n21 9.45567
R13456 a_n4238_7449.n65 a_n4238_7449.n23 9.45567
R13457 a_n4238_7449.n68 a_n4238_7449.n25 9.45567
R13458 a_n4238_7449.n70 a_n4238_7449.n27 9.45567
R13459 a_n4238_7449.n74 a_n4238_7449.n29 9.45567
R13460 a_n4238_7449.n60 a_n4238_7449.n31 9.45567
R13461 a_n4238_7449.n62 a_n4238_7449.n33 9.45567
R13462 a_n4238_7449.n75 a_n4238_7449.n72 4.90567
R13463 a_n4238_7449.n18 a_n4238_7449.n17 4.90567
R13464 a_n4238_7449.n37 a_n4238_7449.t2 339.173
R13465 a_n4238_7449.n40 a_n4238_7449.t4 339.173
R13466 a_n4238_7449.n43 a_n4238_7449.t3 339.173
R13467 a_n4238_7449.n46 a_n4238_7449.t1 339.173
R13468 a_n4238_7449.n49 a_n4238_7449.t8 339.173
R13469 a_n4238_7449.n52 a_n4238_7449.t5 339.173
R13470 a_n4238_7449.n55 a_n4238_7449.t0 339.173
R13471 a_n4238_7449.n58 a_n4238_7449.t9 339.173
R13472 a_n4238_7449.n19 a_n4238_7449.n1 3.48794
R13473 a_n4238_7449.n21 a_n4238_7449.n3 3.48794
R13474 a_n4238_7449.n23 a_n4238_7449.n5 3.48794
R13475 a_n4238_7449.n25 a_n4238_7449.n7 3.48794
R13476 a_n4238_7449.n27 a_n4238_7449.n9 3.48794
R13477 a_n4238_7449.n29 a_n4238_7449.n11 3.48794
R13478 a_n4238_7449.n31 a_n4238_7449.n13 3.48794
R13479 a_n4238_7449.n33 a_n4238_7449.n15 3.48794
R13480 a_n4238_7449.t12 a_n4238_7449.n0 10.7089
R13481 a_n4238_7449.n0 a_n4238_7449.n75 10.589
R13482 a_n4238_7449.n34 a_n4238_7449.n15 3.73143
R13483 a_n4238_7449.n32 a_n4238_7449.n13 3.73143
R13484 a_n4238_7449.n30 a_n4238_7449.n11 3.73143
R13485 a_n4238_7449.n28 a_n4238_7449.n9 3.73143
R13486 a_n4238_7449.n26 a_n4238_7449.n7 3.73143
R13487 a_n4238_7449.n24 a_n4238_7449.n5 3.73143
R13488 a_n4238_7449.n22 a_n4238_7449.n3 3.73143
R13489 a_n4238_7449.n20 a_n4238_7449.n1 3.73143
R13490 a_n4238_7449.n72 a_n4238_7449.n18 6.15136
R13491 a_n4238_7449.n37 a_n4238_7449.n19 1.35994
R13492 a_n4238_7449.n40 a_n4238_7449.n21 1.35994
R13493 a_n4238_7449.n43 a_n4238_7449.n23 1.35994
R13494 a_n4238_7449.n46 a_n4238_7449.n25 1.35994
R13495 a_n4238_7449.n49 a_n4238_7449.n27 1.35994
R13496 a_n4238_7449.n52 a_n4238_7449.n29 1.35994
R13497 a_n4238_7449.n55 a_n4238_7449.n31 1.35994
R13498 a_n4238_7449.n77 a_n4238_7449.n2 9.00755
R13499 a_n4238_7449.n79 a_n4238_7449.n4 9.00755
R13500 a_n4238_7449.n65 a_n4238_7449.n6 9.00755
R13501 a_n4238_7449.n68 a_n4238_7449.n8 9.00755
R13502 a_n4238_7449.n70 a_n4238_7449.n10 9.00755
R13503 a_n4238_7449.n74 a_n4238_7449.n12 9.00755
R13504 a_n4238_7449.n60 a_n4238_7449.n14 9.00755
R13505 a_n4238_7449.n62 a_n4238_7449.n16 9.00755
R13506 a_n16148_7944.n41 a_n16148_7944.n21 195.792
R13507 a_n16148_7944.n42 a_n16148_7944.n41 187.833
R13508 a_n16148_7944.n5 a_n16148_7944.n15 6.99781
R13509 a_n16148_7944.n3 a_n16148_7944.n16 6.99781
R13510 a_n16148_7944.n4 a_n16148_7944.n3 5.13815
R13511 a_n16148_7944.n1 a_n16148_7944.n17 6.99781
R13512 a_n16148_7944.n11 a_n16148_7944.n12 6.99781
R13513 a_n16148_7944.n9 a_n16148_7944.n10 6.99781
R13514 a_n16148_7944.n7 a_n16148_7944.n8 6.99781
R13515 a_n16148_7944.n22 a_n16148_7944.t1 135.649
R13516 a_n16148_7944.n22 a_n16148_7944.t0 101.43
R13517 a_n16148_7944.n5 a_n16148_7944.n6 5.13815
R13518 a_n16148_7944.n1 a_n16148_7944.n2 5.13815
R13519 a_n16148_7944.n39 a_n16148_7944.n38 67.2291
R13520 a_n16148_7944.n36 a_n16148_7944.n35 67.2291
R13521 a_n16148_7944.n33 a_n16148_7944.n32 67.2291
R13522 a_n16148_7944.n30 a_n16148_7944.n29 67.2291
R13523 a_n16148_7944.n27 a_n16148_7944.n26 67.2291
R13524 a_n16148_7944.n24 a_n16148_7944.n23 67.2291
R13525 a_n16148_7944.n29 a_n16148_7944.t22 48.8458
R13526 a_n16148_7944.n26 a_n16148_7944.t19 48.8458
R13527 a_n16148_7944.n23 a_n16148_7944.t20 48.8458
R13528 a_n16148_7944.n38 a_n16148_7944.t27 48.8456
R13529 a_n16148_7944.n35 a_n16148_7944.t25 48.8456
R13530 a_n16148_7944.n32 a_n16148_7944.t26 48.8456
R13531 a_n16148_7944.n39 a_n16148_7944.n15 53.4479
R13532 a_n16148_7944.n37 a_n16148_7944.n4 67.3823
R13533 a_n16148_7944.n36 a_n16148_7944.n16 53.4479
R13534 a_n16148_7944.n33 a_n16148_7944.n17 53.4479
R13535 a_n16148_7944.n31 a_n16148_7944.n12 53.4479
R13536 a_n16148_7944.n18 a_n16148_7944.n31 67.3832
R13537 a_n16148_7944.n28 a_n16148_7944.n10 53.4479
R13538 a_n16148_7944.n19 a_n16148_7944.n28 67.3832
R13539 a_n16148_7944.n25 a_n16148_7944.n8 53.4479
R13540 a_n16148_7944.n20 a_n16148_7944.n25 67.3832
R13541 a_n16148_7944.n6 a_n16148_7944.n40 67.3823
R13542 a_n16148_7944.n2 a_n16148_7944.n34 67.3823
R13543 a_n16148_7944.n6 a_n16148_7944.t9 48.3479
R13544 a_n16148_7944.n40 a_n16148_7944.t18 17.1913
R13545 a_n16148_7944.n39 a_n16148_7944.t16 17.1913
R13546 a_n16148_7944.n4 a_n16148_7944.t28 48.3479
R13547 a_n16148_7944.n37 a_n16148_7944.t15 17.1913
R13548 a_n16148_7944.n36 a_n16148_7944.t11 17.1913
R13549 a_n16148_7944.n2 a_n16148_7944.t6 48.3479
R13550 a_n16148_7944.n34 a_n16148_7944.t17 17.1913
R13551 a_n16148_7944.n33 a_n16148_7944.t13 17.1913
R13552 a_n16148_7944.n30 a_n16148_7944.t24 17.1913
R13553 a_n16148_7944.n31 a_n16148_7944.t10 17.1913
R13554 a_n16148_7944.n18 a_n16148_7944.t14 48.3473
R13555 a_n16148_7944.n27 a_n16148_7944.t21 17.1913
R13556 a_n16148_7944.n28 a_n16148_7944.t29 17.1913
R13557 a_n16148_7944.n19 a_n16148_7944.t8 48.3473
R13558 a_n16148_7944.n24 a_n16148_7944.t23 17.1913
R13559 a_n16148_7944.n25 a_n16148_7944.t7 17.1913
R13560 a_n16148_7944.n20 a_n16148_7944.t12 48.3473
R13561 a_n16148_7944.n0 a_n16148_7944.n22 12.5597
R13562 a_n16148_7944.n41 a_n16148_7944.n0 11.4887
R13563 a_n16148_7944.n21 a_n16148_7944.t2 9.70349
R13564 a_n16148_7944.n21 a_n16148_7944.t4 9.70349
R13565 a_n16148_7944.n42 a_n16148_7944.t3 9.70349
R13566 a_n16148_7944.t5 a_n16148_7944.n42 9.70349
R13567 a_n16148_7944.n0 a_n16148_7944.n14 8.24786
R13568 a_n16148_7944.n13 a_n16148_7944.n1 6.7537
R13569 a_n16148_7944.n14 a_n16148_7944.n7 6.7537
R13570 a_n16148_7944.n40 a_n16148_7944.n15 53.4474
R13571 a_n16148_7944.n37 a_n16148_7944.n16 53.4474
R13572 a_n16148_7944.n34 a_n16148_7944.n17 53.4474
R13573 a_n16148_7944.n12 a_n16148_7944.n30 53.4474
R13574 a_n16148_7944.n10 a_n16148_7944.n27 53.4474
R13575 a_n16148_7944.n8 a_n16148_7944.n24 53.4474
R13576 a_n16148_7944.n0 a_n16148_7944.n13 11.4692
R13577 a_n16148_7944.n5 a_n16148_7944.n38 8.24659
R13578 a_n16148_7944.n1 a_n16148_7944.n32 8.24659
R13579 a_n16148_7944.n13 a_n16148_7944.n3 7.76726
R13580 a_n16148_7944.n11 a_n16148_7944.n18 7.76508
R13581 a_n16148_7944.n9 a_n16148_7944.n19 7.76508
R13582 a_n16148_7944.n7 a_n16148_7944.n20 7.76508
R13583 a_n16148_7944.n14 a_n16148_7944.n11 6.7537
R13584 a_n16148_7944.n13 a_n16148_7944.n5 6.7537
R13585 a_n16148_7944.n11 a_n16148_7944.n29 5.61943
R13586 a_n16148_7944.n9 a_n16148_7944.n26 5.61943
R13587 a_n16148_7944.n7 a_n16148_7944.n23 5.61943
R13588 a_n16148_7944.n3 a_n16148_7944.n35 5.61939
R13589 a_n16148_7944.n14 a_n16148_7944.n9 5.14007
R13590 VDD.n2728 VDD.n92 471.221
R13591 VDD.n2681 VDD.n90 471.221
R13592 VDD.n2559 VDD.n218 471.221
R13593 VDD.n2557 VDD.n220 471.221
R13594 VDD.n1517 VDD.n1516 471.221
R13595 VDD.n1553 VDD.n1080 471.221
R13596 VDD.n1324 VDD.n1226 471.221
R13597 VDD.n1322 VDD.n1228 471.221
R13598 VDD.n2199 VDD.n2049 351.221
R13599 VDD.n2477 VDD.n283 351.221
R13600 VDD.n2449 VDD.n2448 351.221
R13601 VDD.n2057 VDD.n1897 351.221
R13602 VDD.n1883 VDD.n541 351.221
R13603 VDD.n1853 VDD.n1852 351.221
R13604 VDD.n828 VDD.n765 351.221
R13605 VDD.n1591 VDD.n767 351.221
R13606 VDD.n2426 VDD.n2425 351.221
R13607 VDD.n2487 VDD.n275 351.221
R13608 VDD.n2048 VDD.n1898 351.221
R13609 VDD.n2201 VDD.n515 351.221
R13610 VDD.n1831 VDD.n1830 351.221
R13611 VDD.n1893 VDD.n533 351.221
R13612 VDD.n1038 VDD.n766 351.221
R13613 VDD.n1593 VDD.n763 351.221
R13614 VDD.n1900 VDD.t66 338.822
R13615 VDD.n295 VDD.t104 338.822
R13616 VDD.n2058 VDD.t56 338.822
R13617 VDD.n270 VDD.t95 338.822
R13618 VDD.n796 VDD.t45 338.822
R13619 VDD.n821 VDD.t79 338.822
R13620 VDD.n543 VDD.t87 338.822
R13621 VDD.n1800 VDD.t51 338.822
R13622 VDD.n1552 VDD.t0 304.31
R13623 VDD.t1 VDD.n219 304.31
R13624 VDD.t0 VDD.t36 292.241
R13625 VDD.t15 VDD.t1 292.241
R13626 VDD.t36 VDD.t29 245.26
R13627 VDD.t29 VDD.t31 245.26
R13628 VDD.t31 VDD.t18 245.26
R13629 VDD.t10 VDD.t4 245.26
R13630 VDD.t4 VDD.t6 245.26
R13631 VDD.t6 VDD.t15 245.26
R13632 VDD.n1271 VDD.t76 234.716
R13633 VDD.n1289 VDD.t85 234.716
R13634 VDD.n1308 VDD.t82 234.716
R13635 VDD.n233 VDD.t69 234.716
R13636 VDD.n247 VDD.t72 234.716
R13637 VDD.n261 VDD.t63 234.716
R13638 VDD.n136 VDD.t40 234.716
R13639 VDD.n122 VDD.t58 234.716
R13640 VDD.n104 VDD.t47 234.716
R13641 VDD.n1091 VDD.t98 234.716
R13642 VDD.n1062 VDD.t101 234.716
R13643 VDD.n1076 VDD.t91 234.716
R13644 VDD.n1901 VDD.t65 228.47
R13645 VDD.n296 VDD.t105 228.47
R13646 VDD.n2059 VDD.t55 228.47
R13647 VDD.n271 VDD.t96 228.47
R13648 VDD.n797 VDD.t44 228.47
R13649 VDD.n822 VDD.t78 228.47
R13650 VDD.n544 VDD.t88 228.47
R13651 VDD.n1801 VDD.t52 228.47
R13652 VDD.n1271 VDD.t73 225.686
R13653 VDD.n1289 VDD.t83 225.686
R13654 VDD.n1308 VDD.t80 225.686
R13655 VDD.n233 VDD.t67 225.686
R13656 VDD.n247 VDD.t70 225.686
R13657 VDD.n261 VDD.t60 225.686
R13658 VDD.n136 VDD.t38 225.686
R13659 VDD.n122 VDD.t57 225.686
R13660 VDD.n104 VDD.t46 225.686
R13661 VDD.n1091 VDD.t97 225.686
R13662 VDD.n1062 VDD.t100 225.686
R13663 VDD.n1076 VDD.t89 225.686
R13664 VDD.n1900 VDD.t64 225.288
R13665 VDD.n295 VDD.t103 225.288
R13666 VDD.n2058 VDD.t53 225.288
R13667 VDD.n270 VDD.t93 225.288
R13668 VDD.n796 VDD.t42 225.288
R13669 VDD.n821 VDD.t77 225.288
R13670 VDD.n543 VDD.t86 225.288
R13671 VDD.n1800 VDD.t49 225.288
R13672 VDD.n1832 VDD.n1831 185
R13673 VDD.n1831 VDD.n516 185
R13674 VDD.n1833 VDD.n539 185
R13675 VDD.n1888 VDD.n539 185
R13676 VDD.n1835 VDD.n1834 185
R13677 VDD.n1834 VDD.n537 185
R13678 VDD.n1836 VDD.n550 185
R13679 VDD.n1846 VDD.n550 185
R13680 VDD.n1837 VDD.n558 185
R13681 VDD.n558 VDD.n548 185
R13682 VDD.n1839 VDD.n1838 185
R13683 VDD.n1840 VDD.n1839 185
R13684 VDD.n1799 VDD.n557 185
R13685 VDD.n557 VDD.n554 185
R13686 VDD.n1798 VDD.n1797 185
R13687 VDD.n1797 VDD.n1796 185
R13688 VDD.n560 VDD.n559 185
R13689 VDD.n561 VDD.n560 185
R13690 VDD.n1789 VDD.n1788 185
R13691 VDD.n1790 VDD.n1789 185
R13692 VDD.n1787 VDD.n569 185
R13693 VDD.n937 VDD.n569 185
R13694 VDD.n1786 VDD.n1785 185
R13695 VDD.n1785 VDD.n1784 185
R13696 VDD.n571 VDD.n570 185
R13697 VDD.n572 VDD.n571 185
R13698 VDD.n1777 VDD.n1776 185
R13699 VDD.n1778 VDD.n1777 185
R13700 VDD.n1775 VDD.n581 185
R13701 VDD.n581 VDD.n578 185
R13702 VDD.n1774 VDD.n1773 185
R13703 VDD.n1773 VDD.n1772 185
R13704 VDD.n583 VDD.n582 185
R13705 VDD.n584 VDD.n583 185
R13706 VDD.n1765 VDD.n1764 185
R13707 VDD.n1766 VDD.n1765 185
R13708 VDD.n1763 VDD.n593 185
R13709 VDD.n593 VDD.n590 185
R13710 VDD.n1762 VDD.n1761 185
R13711 VDD.n1761 VDD.n1760 185
R13712 VDD.n595 VDD.n594 185
R13713 VDD.n596 VDD.n595 185
R13714 VDD.n1753 VDD.n1752 185
R13715 VDD.n1754 VDD.n1753 185
R13716 VDD.n1751 VDD.n605 185
R13717 VDD.n605 VDD.n602 185
R13718 VDD.n1750 VDD.n1749 185
R13719 VDD.n1749 VDD.n1748 185
R13720 VDD.n607 VDD.n606 185
R13721 VDD.n608 VDD.n607 185
R13722 VDD.n1741 VDD.n1740 185
R13723 VDD.n1742 VDD.n1741 185
R13724 VDD.n1739 VDD.n617 185
R13725 VDD.n617 VDD.n614 185
R13726 VDD.n1738 VDD.n1737 185
R13727 VDD.n1737 VDD.n1736 185
R13728 VDD.n619 VDD.n618 185
R13729 VDD.n620 VDD.n619 185
R13730 VDD.n1729 VDD.n1728 185
R13731 VDD.n1730 VDD.n1729 185
R13732 VDD.n1727 VDD.n628 185
R13733 VDD.n634 VDD.n628 185
R13734 VDD.n1726 VDD.n1725 185
R13735 VDD.n1725 VDD.n1724 185
R13736 VDD.n630 VDD.n629 185
R13737 VDD.n631 VDD.n630 185
R13738 VDD.n1717 VDD.n1716 185
R13739 VDD.n1718 VDD.n1717 185
R13740 VDD.n1715 VDD.n641 185
R13741 VDD.n641 VDD.n638 185
R13742 VDD.n1714 VDD.n1713 185
R13743 VDD.n1713 VDD.n1712 185
R13744 VDD.n643 VDD.n642 185
R13745 VDD.n644 VDD.n643 185
R13746 VDD.n1705 VDD.n1704 185
R13747 VDD.n1706 VDD.n1705 185
R13748 VDD.n1703 VDD.n653 185
R13749 VDD.n653 VDD.n650 185
R13750 VDD.n1702 VDD.n1701 185
R13751 VDD.n1701 VDD.n1700 185
R13752 VDD.n655 VDD.n654 185
R13753 VDD.n656 VDD.n655 185
R13754 VDD.n1693 VDD.n1692 185
R13755 VDD.n1694 VDD.n1693 185
R13756 VDD.n1691 VDD.n665 185
R13757 VDD.n665 VDD.n662 185
R13758 VDD.n1690 VDD.n1689 185
R13759 VDD.n1689 VDD.n1688 185
R13760 VDD.n667 VDD.n666 185
R13761 VDD.n675 VDD.n667 185
R13762 VDD.n1681 VDD.n1680 185
R13763 VDD.n1682 VDD.n1681 185
R13764 VDD.n1679 VDD.n676 185
R13765 VDD.n682 VDD.n676 185
R13766 VDD.n1678 VDD.n1677 185
R13767 VDD.n1677 VDD.n1676 185
R13768 VDD.n678 VDD.n677 185
R13769 VDD.n679 VDD.n678 185
R13770 VDD.n1669 VDD.n1668 185
R13771 VDD.n1670 VDD.n1669 185
R13772 VDD.n1667 VDD.n689 185
R13773 VDD.n689 VDD.n686 185
R13774 VDD.n1666 VDD.n1665 185
R13775 VDD.n1665 VDD.n1664 185
R13776 VDD.n691 VDD.n690 185
R13777 VDD.n692 VDD.n691 185
R13778 VDD.n1657 VDD.n1656 185
R13779 VDD.n1658 VDD.n1657 185
R13780 VDD.n1655 VDD.n701 185
R13781 VDD.n701 VDD.n698 185
R13782 VDD.n1654 VDD.n1653 185
R13783 VDD.n1653 VDD.n1652 185
R13784 VDD.n703 VDD.n702 185
R13785 VDD.n704 VDD.n703 185
R13786 VDD.n1645 VDD.n1644 185
R13787 VDD.n1646 VDD.n1645 185
R13788 VDD.n1643 VDD.n713 185
R13789 VDD.n713 VDD.n710 185
R13790 VDD.n1642 VDD.n1641 185
R13791 VDD.n1641 VDD.n1640 185
R13792 VDD.n715 VDD.n714 185
R13793 VDD.n716 VDD.n715 185
R13794 VDD.n1633 VDD.n1632 185
R13795 VDD.n1634 VDD.n1633 185
R13796 VDD.n1631 VDD.n725 185
R13797 VDD.n725 VDD.n722 185
R13798 VDD.n1630 VDD.n1629 185
R13799 VDD.n1629 VDD.n1628 185
R13800 VDD.n727 VDD.n726 185
R13801 VDD.n728 VDD.n727 185
R13802 VDD.n1621 VDD.n1620 185
R13803 VDD.n1622 VDD.n1621 185
R13804 VDD.n1619 VDD.n736 185
R13805 VDD.n742 VDD.n736 185
R13806 VDD.n1618 VDD.n1617 185
R13807 VDD.n1617 VDD.n1616 185
R13808 VDD.n738 VDD.n737 185
R13809 VDD.n739 VDD.n738 185
R13810 VDD.n1609 VDD.n1608 185
R13811 VDD.n1610 VDD.n1609 185
R13812 VDD.n1607 VDD.n749 185
R13813 VDD.n749 VDD.n746 185
R13814 VDD.n1606 VDD.n1605 185
R13815 VDD.n1605 VDD.n1604 185
R13816 VDD.n751 VDD.n750 185
R13817 VDD.n752 VDD.n751 185
R13818 VDD.n1597 VDD.n1596 185
R13819 VDD.n1598 VDD.n1597 185
R13820 VDD.n1595 VDD.n761 185
R13821 VDD.n761 VDD.n758 185
R13822 VDD.n1594 VDD.n1593 185
R13823 VDD.n1593 VDD.n1592 185
R13824 VDD.n763 VDD.n762 185
R13825 VDD.n780 VDD.n779 185
R13826 VDD.n782 VDD.n781 185
R13827 VDD.n784 VDD.n777 185
R13828 VDD.n787 VDD.n786 185
R13829 VDD.n788 VDD.n776 185
R13830 VDD.n790 VDD.n789 185
R13831 VDD.n792 VDD.n774 185
R13832 VDD.n1053 VDD.n1052 185
R13833 VDD.n1050 VDD.n775 185
R13834 VDD.n1049 VDD.n1048 185
R13835 VDD.n1047 VDD.n1046 185
R13836 VDD.n1045 VDD.n794 185
R13837 VDD.n1043 VDD.n1042 185
R13838 VDD.n1040 VDD.n795 185
R13839 VDD.n1039 VDD.n1038 185
R13840 VDD.n1893 VDD.n1892 185
R13841 VDD.n534 VDD.n532 185
R13842 VDD.n1804 VDD.n1803 185
R13843 VDD.n1806 VDD.n1805 185
R13844 VDD.n1808 VDD.n1807 185
R13845 VDD.n1810 VDD.n1809 185
R13846 VDD.n1812 VDD.n1811 185
R13847 VDD.n1814 VDD.n1813 185
R13848 VDD.n1816 VDD.n1815 185
R13849 VDD.n1818 VDD.n1817 185
R13850 VDD.n1820 VDD.n1819 185
R13851 VDD.n1822 VDD.n1821 185
R13852 VDD.n1824 VDD.n1823 185
R13853 VDD.n1826 VDD.n1825 185
R13854 VDD.n1828 VDD.n1827 185
R13855 VDD.n1830 VDD.n1829 185
R13856 VDD.n1891 VDD.n533 185
R13857 VDD.n533 VDD.n516 185
R13858 VDD.n1890 VDD.n1889 185
R13859 VDD.n1889 VDD.n1888 185
R13860 VDD.n536 VDD.n535 185
R13861 VDD.n537 VDD.n536 185
R13862 VDD.n798 VDD.n549 185
R13863 VDD.n1846 VDD.n549 185
R13864 VDD.n800 VDD.n799 185
R13865 VDD.n799 VDD.n548 185
R13866 VDD.n801 VDD.n556 185
R13867 VDD.n1840 VDD.n556 185
R13868 VDD.n803 VDD.n802 185
R13869 VDD.n802 VDD.n554 185
R13870 VDD.n804 VDD.n563 185
R13871 VDD.n1796 VDD.n563 185
R13872 VDD.n806 VDD.n805 185
R13873 VDD.n805 VDD.n561 185
R13874 VDD.n807 VDD.n568 185
R13875 VDD.n1790 VDD.n568 185
R13876 VDD.n939 VDD.n938 185
R13877 VDD.n938 VDD.n937 185
R13878 VDD.n940 VDD.n574 185
R13879 VDD.n1784 VDD.n574 185
R13880 VDD.n942 VDD.n941 185
R13881 VDD.n941 VDD.n572 185
R13882 VDD.n943 VDD.n580 185
R13883 VDD.n1778 VDD.n580 185
R13884 VDD.n945 VDD.n944 185
R13885 VDD.n944 VDD.n578 185
R13886 VDD.n946 VDD.n586 185
R13887 VDD.n1772 VDD.n586 185
R13888 VDD.n948 VDD.n947 185
R13889 VDD.n947 VDD.n584 185
R13890 VDD.n949 VDD.n592 185
R13891 VDD.n1766 VDD.n592 185
R13892 VDD.n951 VDD.n950 185
R13893 VDD.n950 VDD.n590 185
R13894 VDD.n952 VDD.n598 185
R13895 VDD.n1760 VDD.n598 185
R13896 VDD.n954 VDD.n953 185
R13897 VDD.n953 VDD.n596 185
R13898 VDD.n955 VDD.n604 185
R13899 VDD.n1754 VDD.n604 185
R13900 VDD.n957 VDD.n956 185
R13901 VDD.n956 VDD.n602 185
R13902 VDD.n958 VDD.n610 185
R13903 VDD.n1748 VDD.n610 185
R13904 VDD.n960 VDD.n959 185
R13905 VDD.n959 VDD.n608 185
R13906 VDD.n961 VDD.n616 185
R13907 VDD.n1742 VDD.n616 185
R13908 VDD.n963 VDD.n962 185
R13909 VDD.n962 VDD.n614 185
R13910 VDD.n964 VDD.n622 185
R13911 VDD.n1736 VDD.n622 185
R13912 VDD.n966 VDD.n965 185
R13913 VDD.n965 VDD.n620 185
R13914 VDD.n967 VDD.n627 185
R13915 VDD.n1730 VDD.n627 185
R13916 VDD.n969 VDD.n968 185
R13917 VDD.n968 VDD.n634 185
R13918 VDD.n970 VDD.n633 185
R13919 VDD.n1724 VDD.n633 185
R13920 VDD.n972 VDD.n971 185
R13921 VDD.n971 VDD.n631 185
R13922 VDD.n973 VDD.n640 185
R13923 VDD.n1718 VDD.n640 185
R13924 VDD.n975 VDD.n974 185
R13925 VDD.n974 VDD.n638 185
R13926 VDD.n976 VDD.n646 185
R13927 VDD.n1712 VDD.n646 185
R13928 VDD.n978 VDD.n977 185
R13929 VDD.n977 VDD.n644 185
R13930 VDD.n979 VDD.n652 185
R13931 VDD.n1706 VDD.n652 185
R13932 VDD.n981 VDD.n980 185
R13933 VDD.n980 VDD.n650 185
R13934 VDD.n982 VDD.n658 185
R13935 VDD.n1700 VDD.n658 185
R13936 VDD.n984 VDD.n983 185
R13937 VDD.n983 VDD.n656 185
R13938 VDD.n985 VDD.n664 185
R13939 VDD.n1694 VDD.n664 185
R13940 VDD.n987 VDD.n986 185
R13941 VDD.n986 VDD.n662 185
R13942 VDD.n988 VDD.n669 185
R13943 VDD.n1688 VDD.n669 185
R13944 VDD.n990 VDD.n989 185
R13945 VDD.n989 VDD.n675 185
R13946 VDD.n991 VDD.n674 185
R13947 VDD.n1682 VDD.n674 185
R13948 VDD.n993 VDD.n992 185
R13949 VDD.n992 VDD.n682 185
R13950 VDD.n994 VDD.n681 185
R13951 VDD.n1676 VDD.n681 185
R13952 VDD.n996 VDD.n995 185
R13953 VDD.n995 VDD.n679 185
R13954 VDD.n997 VDD.n688 185
R13955 VDD.n1670 VDD.n688 185
R13956 VDD.n999 VDD.n998 185
R13957 VDD.n998 VDD.n686 185
R13958 VDD.n1000 VDD.n694 185
R13959 VDD.n1664 VDD.n694 185
R13960 VDD.n1002 VDD.n1001 185
R13961 VDD.n1001 VDD.n692 185
R13962 VDD.n1003 VDD.n700 185
R13963 VDD.n1658 VDD.n700 185
R13964 VDD.n1005 VDD.n1004 185
R13965 VDD.n1004 VDD.n698 185
R13966 VDD.n1006 VDD.n706 185
R13967 VDD.n1652 VDD.n706 185
R13968 VDD.n1008 VDD.n1007 185
R13969 VDD.n1007 VDD.n704 185
R13970 VDD.n1009 VDD.n712 185
R13971 VDD.n1646 VDD.n712 185
R13972 VDD.n1011 VDD.n1010 185
R13973 VDD.n1010 VDD.n710 185
R13974 VDD.n1012 VDD.n718 185
R13975 VDD.n1640 VDD.n718 185
R13976 VDD.n1014 VDD.n1013 185
R13977 VDD.n1013 VDD.n716 185
R13978 VDD.n1015 VDD.n724 185
R13979 VDD.n1634 VDD.n724 185
R13980 VDD.n1017 VDD.n1016 185
R13981 VDD.n1016 VDD.n722 185
R13982 VDD.n1018 VDD.n730 185
R13983 VDD.n1628 VDD.n730 185
R13984 VDD.n1020 VDD.n1019 185
R13985 VDD.n1019 VDD.n728 185
R13986 VDD.n1021 VDD.n735 185
R13987 VDD.n1622 VDD.n735 185
R13988 VDD.n1023 VDD.n1022 185
R13989 VDD.n1022 VDD.n742 185
R13990 VDD.n1024 VDD.n741 185
R13991 VDD.n1616 VDD.n741 185
R13992 VDD.n1026 VDD.n1025 185
R13993 VDD.n1025 VDD.n739 185
R13994 VDD.n1027 VDD.n748 185
R13995 VDD.n1610 VDD.n748 185
R13996 VDD.n1029 VDD.n1028 185
R13997 VDD.n1028 VDD.n746 185
R13998 VDD.n1030 VDD.n754 185
R13999 VDD.n1604 VDD.n754 185
R14000 VDD.n1032 VDD.n1031 185
R14001 VDD.n1031 VDD.n752 185
R14002 VDD.n1033 VDD.n760 185
R14003 VDD.n1598 VDD.n760 185
R14004 VDD.n1035 VDD.n1034 185
R14005 VDD.n1034 VDD.n758 185
R14006 VDD.n1036 VDD.n766 185
R14007 VDD.n1592 VDD.n766 185
R14008 VDD.n2427 VDD.n2426 185
R14009 VDD.n2426 VDD.n280 185
R14010 VDD.n2428 VDD.n281 185
R14011 VDD.n2482 VDD.n281 185
R14012 VDD.n2430 VDD.n2429 185
R14013 VDD.n2429 VDD.n278 185
R14014 VDD.n2431 VDD.n301 185
R14015 VDD.n2441 VDD.n301 185
R14016 VDD.n2432 VDD.n309 185
R14017 VDD.n309 VDD.n299 185
R14018 VDD.n2434 VDD.n2433 185
R14019 VDD.n2435 VDD.n2434 185
R14020 VDD.n2407 VDD.n308 185
R14021 VDD.n308 VDD.n305 185
R14022 VDD.n2406 VDD.n2405 185
R14023 VDD.n2405 VDD.n2404 185
R14024 VDD.n311 VDD.n310 185
R14025 VDD.n312 VDD.n311 185
R14026 VDD.n2397 VDD.n2396 185
R14027 VDD.n2398 VDD.n2397 185
R14028 VDD.n2395 VDD.n320 185
R14029 VDD.n326 VDD.n320 185
R14030 VDD.n2394 VDD.n2393 185
R14031 VDD.n2393 VDD.n2392 185
R14032 VDD.n322 VDD.n321 185
R14033 VDD.n323 VDD.n322 185
R14034 VDD.n2385 VDD.n2384 185
R14035 VDD.n2386 VDD.n2385 185
R14036 VDD.n2383 VDD.n333 185
R14037 VDD.n333 VDD.n330 185
R14038 VDD.n2382 VDD.n2381 185
R14039 VDD.n2381 VDD.n2380 185
R14040 VDD.n335 VDD.n334 185
R14041 VDD.n336 VDD.n335 185
R14042 VDD.n2373 VDD.n2372 185
R14043 VDD.n2374 VDD.n2373 185
R14044 VDD.n2371 VDD.n345 185
R14045 VDD.n345 VDD.n342 185
R14046 VDD.n2370 VDD.n2369 185
R14047 VDD.n2369 VDD.n2368 185
R14048 VDD.n347 VDD.n346 185
R14049 VDD.n348 VDD.n347 185
R14050 VDD.n2361 VDD.n2360 185
R14051 VDD.n2362 VDD.n2361 185
R14052 VDD.n2359 VDD.n357 185
R14053 VDD.n357 VDD.n354 185
R14054 VDD.n2358 VDD.n2357 185
R14055 VDD.n2357 VDD.n2356 185
R14056 VDD.n359 VDD.n358 185
R14057 VDD.n360 VDD.n359 185
R14058 VDD.n2349 VDD.n2348 185
R14059 VDD.n2350 VDD.n2349 185
R14060 VDD.n2347 VDD.n369 185
R14061 VDD.n369 VDD.n366 185
R14062 VDD.n2346 VDD.n2345 185
R14063 VDD.n2345 VDD.n2344 185
R14064 VDD.n371 VDD.n370 185
R14065 VDD.n372 VDD.n371 185
R14066 VDD.n2337 VDD.n2336 185
R14067 VDD.n2338 VDD.n2337 185
R14068 VDD.n2335 VDD.n380 185
R14069 VDD.n385 VDD.n380 185
R14070 VDD.n2334 VDD.n2333 185
R14071 VDD.n2333 VDD.n2332 185
R14072 VDD.n382 VDD.n381 185
R14073 VDD.n392 VDD.n382 185
R14074 VDD.n2325 VDD.n2324 185
R14075 VDD.n2326 VDD.n2325 185
R14076 VDD.n2323 VDD.n393 185
R14077 VDD.n393 VDD.n389 185
R14078 VDD.n2322 VDD.n2321 185
R14079 VDD.n2321 VDD.n2320 185
R14080 VDD.n395 VDD.n394 185
R14081 VDD.n396 VDD.n395 185
R14082 VDD.n2313 VDD.n2312 185
R14083 VDD.n2314 VDD.n2313 185
R14084 VDD.n2311 VDD.n405 185
R14085 VDD.n405 VDD.n402 185
R14086 VDD.n2310 VDD.n2309 185
R14087 VDD.n2309 VDD.n2308 185
R14088 VDD.n407 VDD.n406 185
R14089 VDD.n408 VDD.n407 185
R14090 VDD.n2301 VDD.n2300 185
R14091 VDD.n2302 VDD.n2301 185
R14092 VDD.n2299 VDD.n417 185
R14093 VDD.n417 VDD.n414 185
R14094 VDD.n2298 VDD.n2297 185
R14095 VDD.n2297 VDD.n2296 185
R14096 VDD.n419 VDD.n418 185
R14097 VDD.n420 VDD.n419 185
R14098 VDD.n2289 VDD.n2288 185
R14099 VDD.n2290 VDD.n2289 185
R14100 VDD.n2287 VDD.n428 185
R14101 VDD.n434 VDD.n428 185
R14102 VDD.n2286 VDD.n2285 185
R14103 VDD.n2285 VDD.n2284 185
R14104 VDD.n430 VDD.n429 185
R14105 VDD.n431 VDD.n430 185
R14106 VDD.n2277 VDD.n2276 185
R14107 VDD.n2278 VDD.n2277 185
R14108 VDD.n2275 VDD.n441 185
R14109 VDD.n441 VDD.n438 185
R14110 VDD.n2274 VDD.n2273 185
R14111 VDD.n2273 VDD.n2272 185
R14112 VDD.n443 VDD.n442 185
R14113 VDD.n444 VDD.n443 185
R14114 VDD.n2265 VDD.n2264 185
R14115 VDD.n2266 VDD.n2265 185
R14116 VDD.n2263 VDD.n453 185
R14117 VDD.n453 VDD.n450 185
R14118 VDD.n2262 VDD.n2261 185
R14119 VDD.n2261 VDD.n2260 185
R14120 VDD.n455 VDD.n454 185
R14121 VDD.n456 VDD.n455 185
R14122 VDD.n2253 VDD.n2252 185
R14123 VDD.n2254 VDD.n2253 185
R14124 VDD.n2251 VDD.n465 185
R14125 VDD.n465 VDD.n462 185
R14126 VDD.n2250 VDD.n2249 185
R14127 VDD.n2249 VDD.n2248 185
R14128 VDD.n467 VDD.n466 185
R14129 VDD.n468 VDD.n467 185
R14130 VDD.n2241 VDD.n2240 185
R14131 VDD.n2242 VDD.n2241 185
R14132 VDD.n2239 VDD.n477 185
R14133 VDD.n477 VDD.n474 185
R14134 VDD.n2238 VDD.n2237 185
R14135 VDD.n2237 VDD.n2236 185
R14136 VDD.n479 VDD.n478 185
R14137 VDD.n480 VDD.n479 185
R14138 VDD.n2229 VDD.n2228 185
R14139 VDD.n2230 VDD.n2229 185
R14140 VDD.n2227 VDD.n488 185
R14141 VDD.n494 VDD.n488 185
R14142 VDD.n2226 VDD.n2225 185
R14143 VDD.n2225 VDD.n2224 185
R14144 VDD.n490 VDD.n489 185
R14145 VDD.n491 VDD.n490 185
R14146 VDD.n2217 VDD.n2216 185
R14147 VDD.n2218 VDD.n2217 185
R14148 VDD.n2215 VDD.n501 185
R14149 VDD.n501 VDD.n498 185
R14150 VDD.n2214 VDD.n2213 185
R14151 VDD.n2213 VDD.n2212 185
R14152 VDD.n503 VDD.n502 185
R14153 VDD.n504 VDD.n503 185
R14154 VDD.n2205 VDD.n2204 185
R14155 VDD.n2206 VDD.n2205 185
R14156 VDD.n2203 VDD.n513 185
R14157 VDD.n513 VDD.n510 185
R14158 VDD.n2202 VDD.n2201 185
R14159 VDD.n2201 VDD.n2200 185
R14160 VDD.n515 VDD.n514 185
R14161 VDD.n1911 VDD.n1909 185
R14162 VDD.n1914 VDD.n1913 185
R14163 VDD.n1915 VDD.n1908 185
R14164 VDD.n1917 VDD.n1916 185
R14165 VDD.n1919 VDD.n1907 185
R14166 VDD.n1922 VDD.n1921 185
R14167 VDD.n1923 VDD.n1906 185
R14168 VDD.n1925 VDD.n1924 185
R14169 VDD.n1927 VDD.n1905 185
R14170 VDD.n1930 VDD.n1929 185
R14171 VDD.n1931 VDD.n1904 185
R14172 VDD.n1933 VDD.n1932 185
R14173 VDD.n1935 VDD.n1903 185
R14174 VDD.n1938 VDD.n1937 185
R14175 VDD.n1939 VDD.n1898 185
R14176 VDD.n2487 VDD.n2486 185
R14177 VDD.n2489 VDD.n274 185
R14178 VDD.n2491 VDD.n2490 185
R14179 VDD.n2492 VDD.n269 185
R14180 VDD.n2494 VDD.n2493 185
R14181 VDD.n2496 VDD.n268 185
R14182 VDD.n2497 VDD.n265 185
R14183 VDD.n2500 VDD.n2499 185
R14184 VDD.n266 VDD.n264 185
R14185 VDD.n2414 VDD.n2413 185
R14186 VDD.n2416 VDD.n2415 185
R14187 VDD.n2418 VDD.n2410 185
R14188 VDD.n2420 VDD.n2419 185
R14189 VDD.n2421 VDD.n2409 185
R14190 VDD.n2423 VDD.n2422 185
R14191 VDD.n2425 VDD.n2408 185
R14192 VDD.n2485 VDD.n275 185
R14193 VDD.n280 VDD.n275 185
R14194 VDD.n2484 VDD.n2483 185
R14195 VDD.n2483 VDD.n2482 185
R14196 VDD.n277 VDD.n276 185
R14197 VDD.n278 VDD.n277 185
R14198 VDD.n1940 VDD.n300 185
R14199 VDD.n2441 VDD.n300 185
R14200 VDD.n1942 VDD.n1941 185
R14201 VDD.n1941 VDD.n299 185
R14202 VDD.n1943 VDD.n307 185
R14203 VDD.n2435 VDD.n307 185
R14204 VDD.n1945 VDD.n1944 185
R14205 VDD.n1944 VDD.n305 185
R14206 VDD.n1946 VDD.n314 185
R14207 VDD.n2404 VDD.n314 185
R14208 VDD.n1948 VDD.n1947 185
R14209 VDD.n1947 VDD.n312 185
R14210 VDD.n1949 VDD.n319 185
R14211 VDD.n2398 VDD.n319 185
R14212 VDD.n1951 VDD.n1950 185
R14213 VDD.n1950 VDD.n326 185
R14214 VDD.n1952 VDD.n325 185
R14215 VDD.n2392 VDD.n325 185
R14216 VDD.n1954 VDD.n1953 185
R14217 VDD.n1953 VDD.n323 185
R14218 VDD.n1955 VDD.n332 185
R14219 VDD.n2386 VDD.n332 185
R14220 VDD.n1957 VDD.n1956 185
R14221 VDD.n1956 VDD.n330 185
R14222 VDD.n1958 VDD.n338 185
R14223 VDD.n2380 VDD.n338 185
R14224 VDD.n1960 VDD.n1959 185
R14225 VDD.n1959 VDD.n336 185
R14226 VDD.n1961 VDD.n344 185
R14227 VDD.n2374 VDD.n344 185
R14228 VDD.n1963 VDD.n1962 185
R14229 VDD.n1962 VDD.n342 185
R14230 VDD.n1964 VDD.n350 185
R14231 VDD.n2368 VDD.n350 185
R14232 VDD.n1966 VDD.n1965 185
R14233 VDD.n1965 VDD.n348 185
R14234 VDD.n1967 VDD.n356 185
R14235 VDD.n2362 VDD.n356 185
R14236 VDD.n1969 VDD.n1968 185
R14237 VDD.n1968 VDD.n354 185
R14238 VDD.n1970 VDD.n362 185
R14239 VDD.n2356 VDD.n362 185
R14240 VDD.n1972 VDD.n1971 185
R14241 VDD.n1971 VDD.n360 185
R14242 VDD.n1973 VDD.n368 185
R14243 VDD.n2350 VDD.n368 185
R14244 VDD.n1975 VDD.n1974 185
R14245 VDD.n1974 VDD.n366 185
R14246 VDD.n1976 VDD.n374 185
R14247 VDD.n2344 VDD.n374 185
R14248 VDD.n1978 VDD.n1977 185
R14249 VDD.n1977 VDD.n372 185
R14250 VDD.n1979 VDD.n379 185
R14251 VDD.n2338 VDD.n379 185
R14252 VDD.n1981 VDD.n1980 185
R14253 VDD.n1980 VDD.n385 185
R14254 VDD.n1982 VDD.n384 185
R14255 VDD.n2332 VDD.n384 185
R14256 VDD.n1984 VDD.n1983 185
R14257 VDD.n1983 VDD.n392 185
R14258 VDD.n1985 VDD.n391 185
R14259 VDD.n2326 VDD.n391 185
R14260 VDD.n1987 VDD.n1986 185
R14261 VDD.n1986 VDD.n389 185
R14262 VDD.n1988 VDD.n398 185
R14263 VDD.n2320 VDD.n398 185
R14264 VDD.n1990 VDD.n1989 185
R14265 VDD.n1989 VDD.n396 185
R14266 VDD.n1991 VDD.n404 185
R14267 VDD.n2314 VDD.n404 185
R14268 VDD.n1993 VDD.n1992 185
R14269 VDD.n1992 VDD.n402 185
R14270 VDD.n1994 VDD.n410 185
R14271 VDD.n2308 VDD.n410 185
R14272 VDD.n1996 VDD.n1995 185
R14273 VDD.n1995 VDD.n408 185
R14274 VDD.n1997 VDD.n416 185
R14275 VDD.n2302 VDD.n416 185
R14276 VDD.n1999 VDD.n1998 185
R14277 VDD.n1998 VDD.n414 185
R14278 VDD.n2000 VDD.n422 185
R14279 VDD.n2296 VDD.n422 185
R14280 VDD.n2002 VDD.n2001 185
R14281 VDD.n2001 VDD.n420 185
R14282 VDD.n2003 VDD.n427 185
R14283 VDD.n2290 VDD.n427 185
R14284 VDD.n2005 VDD.n2004 185
R14285 VDD.n2004 VDD.n434 185
R14286 VDD.n2006 VDD.n433 185
R14287 VDD.n2284 VDD.n433 185
R14288 VDD.n2008 VDD.n2007 185
R14289 VDD.n2007 VDD.n431 185
R14290 VDD.n2009 VDD.n440 185
R14291 VDD.n2278 VDD.n440 185
R14292 VDD.n2011 VDD.n2010 185
R14293 VDD.n2010 VDD.n438 185
R14294 VDD.n2012 VDD.n446 185
R14295 VDD.n2272 VDD.n446 185
R14296 VDD.n2014 VDD.n2013 185
R14297 VDD.n2013 VDD.n444 185
R14298 VDD.n2015 VDD.n452 185
R14299 VDD.n2266 VDD.n452 185
R14300 VDD.n2017 VDD.n2016 185
R14301 VDD.n2016 VDD.n450 185
R14302 VDD.n2018 VDD.n458 185
R14303 VDD.n2260 VDD.n458 185
R14304 VDD.n2020 VDD.n2019 185
R14305 VDD.n2019 VDD.n456 185
R14306 VDD.n2021 VDD.n464 185
R14307 VDD.n2254 VDD.n464 185
R14308 VDD.n2023 VDD.n2022 185
R14309 VDD.n2022 VDD.n462 185
R14310 VDD.n2024 VDD.n470 185
R14311 VDD.n2248 VDD.n470 185
R14312 VDD.n2026 VDD.n2025 185
R14313 VDD.n2025 VDD.n468 185
R14314 VDD.n2027 VDD.n476 185
R14315 VDD.n2242 VDD.n476 185
R14316 VDD.n2029 VDD.n2028 185
R14317 VDD.n2028 VDD.n474 185
R14318 VDD.n2030 VDD.n482 185
R14319 VDD.n2236 VDD.n482 185
R14320 VDD.n2032 VDD.n2031 185
R14321 VDD.n2031 VDD.n480 185
R14322 VDD.n2033 VDD.n487 185
R14323 VDD.n2230 VDD.n487 185
R14324 VDD.n2035 VDD.n2034 185
R14325 VDD.n2034 VDD.n494 185
R14326 VDD.n2036 VDD.n493 185
R14327 VDD.n2224 VDD.n493 185
R14328 VDD.n2038 VDD.n2037 185
R14329 VDD.n2037 VDD.n491 185
R14330 VDD.n2039 VDD.n500 185
R14331 VDD.n2218 VDD.n500 185
R14332 VDD.n2041 VDD.n2040 185
R14333 VDD.n2040 VDD.n498 185
R14334 VDD.n2042 VDD.n506 185
R14335 VDD.n2212 VDD.n506 185
R14336 VDD.n2044 VDD.n2043 185
R14337 VDD.n2043 VDD.n504 185
R14338 VDD.n2045 VDD.n512 185
R14339 VDD.n2206 VDD.n512 185
R14340 VDD.n2046 VDD.n1899 185
R14341 VDD.n1899 VDD.n510 185
R14342 VDD.n2048 VDD.n2047 185
R14343 VDD.n2200 VDD.n2048 185
R14344 VDD.n1885 VDD.n541 185
R14345 VDD.n541 VDD.n516 185
R14346 VDD.n1887 VDD.n1886 185
R14347 VDD.n1888 VDD.n1887 185
R14348 VDD.n542 VDD.n540 185
R14349 VDD.n540 VDD.n537 185
R14350 VDD.n1845 VDD.n1844 185
R14351 VDD.n1846 VDD.n1845 185
R14352 VDD.n1843 VDD.n551 185
R14353 VDD.n551 VDD.n548 185
R14354 VDD.n1842 VDD.n1841 185
R14355 VDD.n1841 VDD.n1840 185
R14356 VDD.n553 VDD.n552 185
R14357 VDD.n554 VDD.n553 185
R14358 VDD.n1795 VDD.n1794 185
R14359 VDD.n1796 VDD.n1795 185
R14360 VDD.n1793 VDD.n564 185
R14361 VDD.n564 VDD.n561 185
R14362 VDD.n1792 VDD.n1791 185
R14363 VDD.n1791 VDD.n1790 185
R14364 VDD.n566 VDD.n565 185
R14365 VDD.n937 VDD.n566 185
R14366 VDD.n1783 VDD.n1782 185
R14367 VDD.n1784 VDD.n1783 185
R14368 VDD.n1781 VDD.n575 185
R14369 VDD.n575 VDD.n572 185
R14370 VDD.n1780 VDD.n1779 185
R14371 VDD.n1779 VDD.n1778 185
R14372 VDD.n577 VDD.n576 185
R14373 VDD.n578 VDD.n577 185
R14374 VDD.n1771 VDD.n1770 185
R14375 VDD.n1772 VDD.n1771 185
R14376 VDD.n1769 VDD.n587 185
R14377 VDD.n587 VDD.n584 185
R14378 VDD.n1768 VDD.n1767 185
R14379 VDD.n1767 VDD.n1766 185
R14380 VDD.n589 VDD.n588 185
R14381 VDD.n590 VDD.n589 185
R14382 VDD.n1759 VDD.n1758 185
R14383 VDD.n1760 VDD.n1759 185
R14384 VDD.n1757 VDD.n599 185
R14385 VDD.n599 VDD.n596 185
R14386 VDD.n1756 VDD.n1755 185
R14387 VDD.n1755 VDD.n1754 185
R14388 VDD.n601 VDD.n600 185
R14389 VDD.n602 VDD.n601 185
R14390 VDD.n1747 VDD.n1746 185
R14391 VDD.n1748 VDD.n1747 185
R14392 VDD.n1745 VDD.n611 185
R14393 VDD.n611 VDD.n608 185
R14394 VDD.n1744 VDD.n1743 185
R14395 VDD.n1743 VDD.n1742 185
R14396 VDD.n613 VDD.n612 185
R14397 VDD.n614 VDD.n613 185
R14398 VDD.n1735 VDD.n1734 185
R14399 VDD.n1736 VDD.n1735 185
R14400 VDD.n1733 VDD.n623 185
R14401 VDD.n623 VDD.n620 185
R14402 VDD.n1732 VDD.n1731 185
R14403 VDD.n1731 VDD.n1730 185
R14404 VDD.n625 VDD.n624 185
R14405 VDD.n634 VDD.n625 185
R14406 VDD.n1723 VDD.n1722 185
R14407 VDD.n1724 VDD.n1723 185
R14408 VDD.n1721 VDD.n635 185
R14409 VDD.n635 VDD.n631 185
R14410 VDD.n1720 VDD.n1719 185
R14411 VDD.n1719 VDD.n1718 185
R14412 VDD.n637 VDD.n636 185
R14413 VDD.n638 VDD.n637 185
R14414 VDD.n1711 VDD.n1710 185
R14415 VDD.n1712 VDD.n1711 185
R14416 VDD.n1709 VDD.n647 185
R14417 VDD.n647 VDD.n644 185
R14418 VDD.n1708 VDD.n1707 185
R14419 VDD.n1707 VDD.n1706 185
R14420 VDD.n649 VDD.n648 185
R14421 VDD.n650 VDD.n649 185
R14422 VDD.n1699 VDD.n1698 185
R14423 VDD.n1700 VDD.n1699 185
R14424 VDD.n1697 VDD.n659 185
R14425 VDD.n659 VDD.n656 185
R14426 VDD.n1696 VDD.n1695 185
R14427 VDD.n1695 VDD.n1694 185
R14428 VDD.n661 VDD.n660 185
R14429 VDD.n662 VDD.n661 185
R14430 VDD.n1687 VDD.n1686 185
R14431 VDD.n1688 VDD.n1687 185
R14432 VDD.n1685 VDD.n670 185
R14433 VDD.n675 VDD.n670 185
R14434 VDD.n1684 VDD.n1683 185
R14435 VDD.n1683 VDD.n1682 185
R14436 VDD.n672 VDD.n671 185
R14437 VDD.n682 VDD.n672 185
R14438 VDD.n1675 VDD.n1674 185
R14439 VDD.n1676 VDD.n1675 185
R14440 VDD.n1673 VDD.n683 185
R14441 VDD.n683 VDD.n679 185
R14442 VDD.n1672 VDD.n1671 185
R14443 VDD.n1671 VDD.n1670 185
R14444 VDD.n685 VDD.n684 185
R14445 VDD.n686 VDD.n685 185
R14446 VDD.n1663 VDD.n1662 185
R14447 VDD.n1664 VDD.n1663 185
R14448 VDD.n1661 VDD.n695 185
R14449 VDD.n695 VDD.n692 185
R14450 VDD.n1660 VDD.n1659 185
R14451 VDD.n1659 VDD.n1658 185
R14452 VDD.n697 VDD.n696 185
R14453 VDD.n698 VDD.n697 185
R14454 VDD.n1651 VDD.n1650 185
R14455 VDD.n1652 VDD.n1651 185
R14456 VDD.n1649 VDD.n707 185
R14457 VDD.n707 VDD.n704 185
R14458 VDD.n1648 VDD.n1647 185
R14459 VDD.n1647 VDD.n1646 185
R14460 VDD.n709 VDD.n708 185
R14461 VDD.n710 VDD.n709 185
R14462 VDD.n1639 VDD.n1638 185
R14463 VDD.n1640 VDD.n1639 185
R14464 VDD.n1637 VDD.n719 185
R14465 VDD.n719 VDD.n716 185
R14466 VDD.n1636 VDD.n1635 185
R14467 VDD.n1635 VDD.n1634 185
R14468 VDD.n721 VDD.n720 185
R14469 VDD.n722 VDD.n721 185
R14470 VDD.n1627 VDD.n1626 185
R14471 VDD.n1628 VDD.n1627 185
R14472 VDD.n1625 VDD.n731 185
R14473 VDD.n731 VDD.n728 185
R14474 VDD.n1624 VDD.n1623 185
R14475 VDD.n1623 VDD.n1622 185
R14476 VDD.n733 VDD.n732 185
R14477 VDD.n742 VDD.n733 185
R14478 VDD.n1615 VDD.n1614 185
R14479 VDD.n1616 VDD.n1615 185
R14480 VDD.n1613 VDD.n743 185
R14481 VDD.n743 VDD.n739 185
R14482 VDD.n1612 VDD.n1611 185
R14483 VDD.n1611 VDD.n1610 185
R14484 VDD.n745 VDD.n744 185
R14485 VDD.n746 VDD.n745 185
R14486 VDD.n1603 VDD.n1602 185
R14487 VDD.n1604 VDD.n1603 185
R14488 VDD.n1601 VDD.n755 185
R14489 VDD.n755 VDD.n752 185
R14490 VDD.n1600 VDD.n1599 185
R14491 VDD.n1599 VDD.n1598 185
R14492 VDD.n757 VDD.n756 185
R14493 VDD.n758 VDD.n757 185
R14494 VDD.n1591 VDD.n1590 185
R14495 VDD.n1592 VDD.n1591 185
R14496 VDD.n1589 VDD.n767 185
R14497 VDD.n1588 VDD.n1587 185
R14498 VDD.n1585 VDD.n768 185
R14499 VDD.n1585 VDD.n764 185
R14500 VDD.n1584 VDD.n1583 185
R14501 VDD.n1582 VDD.n1581 185
R14502 VDD.n1580 VDD.n770 185
R14503 VDD.n1578 VDD.n1577 185
R14504 VDD.n1576 VDD.n771 185
R14505 VDD.n812 VDD.n772 185
R14506 VDD.n814 VDD.n813 185
R14507 VDD.n816 VDD.n810 185
R14508 VDD.n819 VDD.n818 185
R14509 VDD.n820 VDD.n809 185
R14510 VDD.n825 VDD.n824 185
R14511 VDD.n827 VDD.n808 185
R14512 VDD.n829 VDD.n828 185
R14513 VDD.n828 VDD.n764 185
R14514 VDD.n1854 VDD.n1853 185
R14515 VDD.n1856 VDD.n1855 185
R14516 VDD.n1858 VDD.n1857 185
R14517 VDD.n1860 VDD.n1859 185
R14518 VDD.n1862 VDD.n1861 185
R14519 VDD.n1864 VDD.n1863 185
R14520 VDD.n1866 VDD.n1865 185
R14521 VDD.n1868 VDD.n1867 185
R14522 VDD.n1870 VDD.n1869 185
R14523 VDD.n1872 VDD.n1871 185
R14524 VDD.n1874 VDD.n1873 185
R14525 VDD.n1876 VDD.n1875 185
R14526 VDD.n1878 VDD.n1877 185
R14527 VDD.n1880 VDD.n1879 185
R14528 VDD.n1882 VDD.n1881 185
R14529 VDD.n1884 VDD.n1883 185
R14530 VDD.n1852 VDD.n1851 185
R14531 VDD.n1852 VDD.n516 185
R14532 VDD.n1850 VDD.n538 185
R14533 VDD.n1888 VDD.n538 185
R14534 VDD.n1849 VDD.n1848 185
R14535 VDD.n1848 VDD.n537 185
R14536 VDD.n1847 VDD.n546 185
R14537 VDD.n1847 VDD.n1846 185
R14538 VDD.n927 VDD.n547 185
R14539 VDD.n548 VDD.n547 185
R14540 VDD.n928 VDD.n555 185
R14541 VDD.n1840 VDD.n555 185
R14542 VDD.n930 VDD.n929 185
R14543 VDD.n929 VDD.n554 185
R14544 VDD.n931 VDD.n562 185
R14545 VDD.n1796 VDD.n562 185
R14546 VDD.n933 VDD.n932 185
R14547 VDD.n932 VDD.n561 185
R14548 VDD.n934 VDD.n567 185
R14549 VDD.n1790 VDD.n567 185
R14550 VDD.n936 VDD.n935 185
R14551 VDD.n937 VDD.n936 185
R14552 VDD.n926 VDD.n573 185
R14553 VDD.n1784 VDD.n573 185
R14554 VDD.n925 VDD.n924 185
R14555 VDD.n924 VDD.n572 185
R14556 VDD.n923 VDD.n579 185
R14557 VDD.n1778 VDD.n579 185
R14558 VDD.n922 VDD.n921 185
R14559 VDD.n921 VDD.n578 185
R14560 VDD.n920 VDD.n585 185
R14561 VDD.n1772 VDD.n585 185
R14562 VDD.n919 VDD.n918 185
R14563 VDD.n918 VDD.n584 185
R14564 VDD.n917 VDD.n591 185
R14565 VDD.n1766 VDD.n591 185
R14566 VDD.n916 VDD.n915 185
R14567 VDD.n915 VDD.n590 185
R14568 VDD.n914 VDD.n597 185
R14569 VDD.n1760 VDD.n597 185
R14570 VDD.n913 VDD.n912 185
R14571 VDD.n912 VDD.n596 185
R14572 VDD.n911 VDD.n603 185
R14573 VDD.n1754 VDD.n603 185
R14574 VDD.n910 VDD.n909 185
R14575 VDD.n909 VDD.n602 185
R14576 VDD.n908 VDD.n609 185
R14577 VDD.n1748 VDD.n609 185
R14578 VDD.n907 VDD.n906 185
R14579 VDD.n906 VDD.n608 185
R14580 VDD.n905 VDD.n615 185
R14581 VDD.n1742 VDD.n615 185
R14582 VDD.n904 VDD.n903 185
R14583 VDD.n903 VDD.n614 185
R14584 VDD.n902 VDD.n621 185
R14585 VDD.n1736 VDD.n621 185
R14586 VDD.n901 VDD.n900 185
R14587 VDD.n900 VDD.n620 185
R14588 VDD.n899 VDD.n626 185
R14589 VDD.n1730 VDD.n626 185
R14590 VDD.n898 VDD.n897 185
R14591 VDD.n897 VDD.n634 185
R14592 VDD.n896 VDD.n632 185
R14593 VDD.n1724 VDD.n632 185
R14594 VDD.n895 VDD.n894 185
R14595 VDD.n894 VDD.n631 185
R14596 VDD.n893 VDD.n639 185
R14597 VDD.n1718 VDD.n639 185
R14598 VDD.n892 VDD.n891 185
R14599 VDD.n891 VDD.n638 185
R14600 VDD.n890 VDD.n645 185
R14601 VDD.n1712 VDD.n645 185
R14602 VDD.n889 VDD.n888 185
R14603 VDD.n888 VDD.n644 185
R14604 VDD.n887 VDD.n651 185
R14605 VDD.n1706 VDD.n651 185
R14606 VDD.n886 VDD.n885 185
R14607 VDD.n885 VDD.n650 185
R14608 VDD.n884 VDD.n657 185
R14609 VDD.n1700 VDD.n657 185
R14610 VDD.n883 VDD.n882 185
R14611 VDD.n882 VDD.n656 185
R14612 VDD.n881 VDD.n663 185
R14613 VDD.n1694 VDD.n663 185
R14614 VDD.n880 VDD.n879 185
R14615 VDD.n879 VDD.n662 185
R14616 VDD.n878 VDD.n668 185
R14617 VDD.n1688 VDD.n668 185
R14618 VDD.n877 VDD.n876 185
R14619 VDD.n876 VDD.n675 185
R14620 VDD.n875 VDD.n673 185
R14621 VDD.n1682 VDD.n673 185
R14622 VDD.n874 VDD.n873 185
R14623 VDD.n873 VDD.n682 185
R14624 VDD.n872 VDD.n680 185
R14625 VDD.n1676 VDD.n680 185
R14626 VDD.n871 VDD.n870 185
R14627 VDD.n870 VDD.n679 185
R14628 VDD.n869 VDD.n687 185
R14629 VDD.n1670 VDD.n687 185
R14630 VDD.n868 VDD.n867 185
R14631 VDD.n867 VDD.n686 185
R14632 VDD.n866 VDD.n693 185
R14633 VDD.n1664 VDD.n693 185
R14634 VDD.n865 VDD.n864 185
R14635 VDD.n864 VDD.n692 185
R14636 VDD.n863 VDD.n699 185
R14637 VDD.n1658 VDD.n699 185
R14638 VDD.n862 VDD.n861 185
R14639 VDD.n861 VDD.n698 185
R14640 VDD.n860 VDD.n705 185
R14641 VDD.n1652 VDD.n705 185
R14642 VDD.n859 VDD.n858 185
R14643 VDD.n858 VDD.n704 185
R14644 VDD.n857 VDD.n711 185
R14645 VDD.n1646 VDD.n711 185
R14646 VDD.n856 VDD.n855 185
R14647 VDD.n855 VDD.n710 185
R14648 VDD.n854 VDD.n717 185
R14649 VDD.n1640 VDD.n717 185
R14650 VDD.n853 VDD.n852 185
R14651 VDD.n852 VDD.n716 185
R14652 VDD.n851 VDD.n723 185
R14653 VDD.n1634 VDD.n723 185
R14654 VDD.n850 VDD.n849 185
R14655 VDD.n849 VDD.n722 185
R14656 VDD.n848 VDD.n729 185
R14657 VDD.n1628 VDD.n729 185
R14658 VDD.n847 VDD.n846 185
R14659 VDD.n846 VDD.n728 185
R14660 VDD.n845 VDD.n734 185
R14661 VDD.n1622 VDD.n734 185
R14662 VDD.n844 VDD.n843 185
R14663 VDD.n843 VDD.n742 185
R14664 VDD.n842 VDD.n740 185
R14665 VDD.n1616 VDD.n740 185
R14666 VDD.n841 VDD.n840 185
R14667 VDD.n840 VDD.n739 185
R14668 VDD.n839 VDD.n747 185
R14669 VDD.n1610 VDD.n747 185
R14670 VDD.n838 VDD.n837 185
R14671 VDD.n837 VDD.n746 185
R14672 VDD.n836 VDD.n753 185
R14673 VDD.n1604 VDD.n753 185
R14674 VDD.n835 VDD.n834 185
R14675 VDD.n834 VDD.n752 185
R14676 VDD.n833 VDD.n759 185
R14677 VDD.n1598 VDD.n759 185
R14678 VDD.n832 VDD.n831 185
R14679 VDD.n831 VDD.n758 185
R14680 VDD.n830 VDD.n765 185
R14681 VDD.n1592 VDD.n765 185
R14682 VDD.n2728 VDD.n2727 185
R14683 VDD.n2729 VDD.n2728 185
R14684 VDD.n86 VDD.n85 185
R14685 VDD.n2730 VDD.n86 185
R14686 VDD.n2733 VDD.n2732 185
R14687 VDD.n2732 VDD.n2731 185
R14688 VDD.n2734 VDD.n80 185
R14689 VDD.n87 VDD.n80 185
R14690 VDD.n2736 VDD.n2735 185
R14691 VDD.n2737 VDD.n2736 185
R14692 VDD.n76 VDD.n75 185
R14693 VDD.n2738 VDD.n76 185
R14694 VDD.n2741 VDD.n2740 185
R14695 VDD.n2740 VDD.n2739 185
R14696 VDD.n2742 VDD.n70 185
R14697 VDD.n70 VDD.n69 185
R14698 VDD.n2744 VDD.n2743 185
R14699 VDD.n2745 VDD.n2744 185
R14700 VDD.n65 VDD.n64 185
R14701 VDD.n2746 VDD.n65 185
R14702 VDD.n2749 VDD.n2748 185
R14703 VDD.n2748 VDD.n2747 185
R14704 VDD.n2750 VDD.n59 185
R14705 VDD.n59 VDD.n58 185
R14706 VDD.n2752 VDD.n2751 185
R14707 VDD.n2753 VDD.n2752 185
R14708 VDD.n54 VDD.n53 185
R14709 VDD.n2754 VDD.n54 185
R14710 VDD.n2757 VDD.n2756 185
R14711 VDD.n2756 VDD.n2755 185
R14712 VDD.n2758 VDD.n48 185
R14713 VDD.n48 VDD.n47 185
R14714 VDD.n2760 VDD.n2759 185
R14715 VDD.n2761 VDD.n2760 185
R14716 VDD.n43 VDD.n42 185
R14717 VDD.n2762 VDD.n43 185
R14718 VDD.n2765 VDD.n2764 185
R14719 VDD.n2764 VDD.n2763 185
R14720 VDD.n2766 VDD.n38 185
R14721 VDD.n38 VDD.n37 185
R14722 VDD.n2768 VDD.n2767 185
R14723 VDD.n2769 VDD.n2768 185
R14724 VDD.n32 VDD.n30 185
R14725 VDD.n2770 VDD.n32 185
R14726 VDD.n2773 VDD.n2772 185
R14727 VDD.n2772 VDD.n2771 185
R14728 VDD.n31 VDD.n29 185
R14729 VDD.n33 VDD.n31 185
R14730 VDD.n2638 VDD.n2637 185
R14731 VDD.n2639 VDD.n2638 185
R14732 VDD.n163 VDD.n162 185
R14733 VDD.n162 VDD.n161 185
R14734 VDD.n2633 VDD.n2632 185
R14735 VDD.n2632 VDD.n2631 185
R14736 VDD.n166 VDD.n165 185
R14737 VDD.n167 VDD.n166 185
R14738 VDD.n2622 VDD.n2621 185
R14739 VDD.n2623 VDD.n2622 185
R14740 VDD.n175 VDD.n174 185
R14741 VDD.n174 VDD.n173 185
R14742 VDD.n2617 VDD.n2616 185
R14743 VDD.n2616 VDD.n2615 185
R14744 VDD.n178 VDD.n177 185
R14745 VDD.n179 VDD.n178 185
R14746 VDD.n2606 VDD.n2605 185
R14747 VDD.n2607 VDD.n2606 185
R14748 VDD.n187 VDD.n186 185
R14749 VDD.n186 VDD.n185 185
R14750 VDD.n2601 VDD.n2600 185
R14751 VDD.n2600 VDD.n2599 185
R14752 VDD.n190 VDD.n189 185
R14753 VDD.n191 VDD.n190 185
R14754 VDD.n2590 VDD.n2589 185
R14755 VDD.n2591 VDD.n2590 185
R14756 VDD.n199 VDD.n198 185
R14757 VDD.n198 VDD.n197 185
R14758 VDD.n2585 VDD.n2584 185
R14759 VDD.n2584 VDD.n2583 185
R14760 VDD.n202 VDD.n201 185
R14761 VDD.n203 VDD.n202 185
R14762 VDD.n2574 VDD.n2573 185
R14763 VDD.n2575 VDD.n2574 185
R14764 VDD.n210 VDD.n209 185
R14765 VDD.n2566 VDD.n209 185
R14766 VDD.n2569 VDD.n2568 185
R14767 VDD.n2568 VDD.n2567 185
R14768 VDD.n213 VDD.n212 185
R14769 VDD.n214 VDD.n213 185
R14770 VDD.n2557 VDD.n2556 185
R14771 VDD.n2558 VDD.n2557 185
R14772 VDD.n2551 VDD.n220 185
R14773 VDD.n2550 VDD.n2549 185
R14774 VDD.n2547 VDD.n224 185
R14775 VDD.n2547 VDD.n219 185
R14776 VDD.n2546 VDD.n2545 185
R14777 VDD.n2544 VDD.n2543 185
R14778 VDD.n2542 VDD.n229 185
R14779 VDD.n2540 VDD.n2539 185
R14780 VDD.n2538 VDD.n230 185
R14781 VDD.n2537 VDD.n2536 185
R14782 VDD.n2534 VDD.n237 185
R14783 VDD.n2532 VDD.n2531 185
R14784 VDD.n2530 VDD.n238 185
R14785 VDD.n2529 VDD.n2528 185
R14786 VDD.n2526 VDD.n242 185
R14787 VDD.n2524 VDD.n2523 185
R14788 VDD.n2522 VDD.n243 185
R14789 VDD.n2521 VDD.n2520 185
R14790 VDD.n2518 VDD.n250 185
R14791 VDD.n2516 VDD.n2515 185
R14792 VDD.n2514 VDD.n251 185
R14793 VDD.n2513 VDD.n2512 185
R14794 VDD.n2510 VDD.n256 185
R14795 VDD.n2508 VDD.n2507 185
R14796 VDD.n2506 VDD.n258 185
R14797 VDD.n2503 VDD.n218 185
R14798 VDD.n2681 VDD.n2680 185
R14799 VDD.n2683 VDD.n134 185
R14800 VDD.n2685 VDD.n2684 185
R14801 VDD.n2686 VDD.n129 185
R14802 VDD.n2688 VDD.n2687 185
R14803 VDD.n2690 VDD.n128 185
R14804 VDD.n2691 VDD.n125 185
R14805 VDD.n2694 VDD.n2693 185
R14806 VDD.n127 VDD.n121 185
R14807 VDD.n2698 VDD.n118 185
R14808 VDD.n2700 VDD.n2699 185
R14809 VDD.n2702 VDD.n116 185
R14810 VDD.n2704 VDD.n2703 185
R14811 VDD.n2705 VDD.n112 185
R14812 VDD.n2707 VDD.n2706 185
R14813 VDD.n2709 VDD.n109 185
R14814 VDD.n2711 VDD.n2710 185
R14815 VDD.n110 VDD.n103 185
R14816 VDD.n2715 VDD.n107 185
R14817 VDD.n2716 VDD.n99 185
R14818 VDD.n2718 VDD.n2717 185
R14819 VDD.n2720 VDD.n97 185
R14820 VDD.n2722 VDD.n2721 185
R14821 VDD.n2723 VDD.n95 185
R14822 VDD.n2724 VDD.n92 185
R14823 VDD.n92 VDD.n91 185
R14824 VDD.n2677 VDD.n90 185
R14825 VDD.n2729 VDD.n90 185
R14826 VDD.n2676 VDD.n89 185
R14827 VDD.n2730 VDD.n89 185
R14828 VDD.n2675 VDD.n88 185
R14829 VDD.n2731 VDD.n88 185
R14830 VDD.n142 VDD.n141 185
R14831 VDD.n141 VDD.n87 185
R14832 VDD.n2671 VDD.n79 185
R14833 VDD.n2737 VDD.n79 185
R14834 VDD.n2670 VDD.n78 185
R14835 VDD.n2738 VDD.n78 185
R14836 VDD.n2669 VDD.n77 185
R14837 VDD.n2739 VDD.n77 185
R14838 VDD.n145 VDD.n144 185
R14839 VDD.n144 VDD.n69 185
R14840 VDD.n2665 VDD.n68 185
R14841 VDD.n2745 VDD.n68 185
R14842 VDD.n2664 VDD.n67 185
R14843 VDD.n2746 VDD.n67 185
R14844 VDD.n2663 VDD.n66 185
R14845 VDD.n2747 VDD.n66 185
R14846 VDD.n148 VDD.n147 185
R14847 VDD.n147 VDD.n58 185
R14848 VDD.n2659 VDD.n57 185
R14849 VDD.n2753 VDD.n57 185
R14850 VDD.n2658 VDD.n56 185
R14851 VDD.n2754 VDD.n56 185
R14852 VDD.n2657 VDD.n55 185
R14853 VDD.n2755 VDD.n55 185
R14854 VDD.n151 VDD.n150 185
R14855 VDD.n150 VDD.n47 185
R14856 VDD.n2653 VDD.n46 185
R14857 VDD.n2761 VDD.n46 185
R14858 VDD.n2652 VDD.n45 185
R14859 VDD.n2762 VDD.n45 185
R14860 VDD.n2651 VDD.n44 185
R14861 VDD.n2763 VDD.n44 185
R14862 VDD.n154 VDD.n153 185
R14863 VDD.n153 VDD.n37 185
R14864 VDD.n2647 VDD.n36 185
R14865 VDD.n2769 VDD.n36 185
R14866 VDD.n2646 VDD.n35 185
R14867 VDD.n2770 VDD.n35 185
R14868 VDD.n2645 VDD.n34 185
R14869 VDD.n2771 VDD.n34 185
R14870 VDD.n160 VDD.n156 185
R14871 VDD.n160 VDD.n33 185
R14872 VDD.n2641 VDD.n2640 185
R14873 VDD.n2640 VDD.n2639 185
R14874 VDD.n159 VDD.n158 185
R14875 VDD.n161 VDD.n159 185
R14876 VDD.n2630 VDD.n2629 185
R14877 VDD.n2631 VDD.n2630 185
R14878 VDD.n169 VDD.n168 185
R14879 VDD.n168 VDD.n167 185
R14880 VDD.n2625 VDD.n2624 185
R14881 VDD.n2624 VDD.n2623 185
R14882 VDD.n172 VDD.n171 185
R14883 VDD.n173 VDD.n172 185
R14884 VDD.n2614 VDD.n2613 185
R14885 VDD.n2615 VDD.n2614 185
R14886 VDD.n181 VDD.n180 185
R14887 VDD.n180 VDD.n179 185
R14888 VDD.n2609 VDD.n2608 185
R14889 VDD.n2608 VDD.n2607 185
R14890 VDD.n184 VDD.n183 185
R14891 VDD.n185 VDD.n184 185
R14892 VDD.n2598 VDD.n2597 185
R14893 VDD.n2599 VDD.n2598 185
R14894 VDD.n193 VDD.n192 185
R14895 VDD.n192 VDD.n191 185
R14896 VDD.n2593 VDD.n2592 185
R14897 VDD.n2592 VDD.n2591 185
R14898 VDD.n196 VDD.n195 185
R14899 VDD.n197 VDD.n196 185
R14900 VDD.n2582 VDD.n2581 185
R14901 VDD.n2583 VDD.n2582 185
R14902 VDD.n205 VDD.n204 185
R14903 VDD.n204 VDD.n203 185
R14904 VDD.n2577 VDD.n2576 185
R14905 VDD.n2576 VDD.n2575 185
R14906 VDD.n208 VDD.n207 185
R14907 VDD.n2566 VDD.n208 185
R14908 VDD.n2565 VDD.n2564 185
R14909 VDD.n2567 VDD.n2565 185
R14910 VDD.n216 VDD.n215 185
R14911 VDD.n215 VDD.n214 185
R14912 VDD.n2560 VDD.n2559 185
R14913 VDD.n2559 VDD.n2558 185
R14914 VDD.n2197 VDD.n2049 185
R14915 VDD.n2196 VDD.n2195 185
R14916 VDD.n2193 VDD.n2050 185
R14917 VDD.n2193 VDD.n1896 185
R14918 VDD.n2192 VDD.n2191 185
R14919 VDD.n2190 VDD.n2189 185
R14920 VDD.n2188 VDD.n2052 185
R14921 VDD.n2186 VDD.n2185 185
R14922 VDD.n2184 VDD.n2053 185
R14923 VDD.n2183 VDD.n2182 185
R14924 VDD.n2180 VDD.n2054 185
R14925 VDD.n2178 VDD.n2177 185
R14926 VDD.n2176 VDD.n2055 185
R14927 VDD.n2175 VDD.n2174 185
R14928 VDD.n2172 VDD.n2056 185
R14929 VDD.n2170 VDD.n2169 185
R14930 VDD.n2168 VDD.n2057 185
R14931 VDD.n2057 VDD.n1896 185
R14932 VDD.n2450 VDD.n2449 185
R14933 VDD.n2451 VDD.n294 185
R14934 VDD.n2454 VDD.n2453 185
R14935 VDD.n2456 VDD.n292 185
R14936 VDD.n2458 VDD.n2457 185
R14937 VDD.n2459 VDD.n291 185
R14938 VDD.n2461 VDD.n2460 185
R14939 VDD.n2463 VDD.n290 185
R14940 VDD.n2465 VDD.n2464 185
R14941 VDD.n2467 VDD.n288 185
R14942 VDD.n2469 VDD.n2468 185
R14943 VDD.n2470 VDD.n287 185
R14944 VDD.n2472 VDD.n2471 185
R14945 VDD.n2474 VDD.n286 185
R14946 VDD.n2475 VDD.n285 185
R14947 VDD.n2478 VDD.n2477 185
R14948 VDD.n2448 VDD.n2446 185
R14949 VDD.n2448 VDD.n280 185
R14950 VDD.n2445 VDD.n279 185
R14951 VDD.n2482 VDD.n279 185
R14952 VDD.n2444 VDD.n2443 185
R14953 VDD.n2443 VDD.n278 185
R14954 VDD.n2442 VDD.n297 185
R14955 VDD.n2442 VDD.n2441 185
R14956 VDD.n2061 VDD.n298 185
R14957 VDD.n299 VDD.n298 185
R14958 VDD.n2062 VDD.n306 185
R14959 VDD.n2435 VDD.n306 185
R14960 VDD.n2064 VDD.n2063 185
R14961 VDD.n2063 VDD.n305 185
R14962 VDD.n2065 VDD.n313 185
R14963 VDD.n2404 VDD.n313 185
R14964 VDD.n2067 VDD.n2066 185
R14965 VDD.n2066 VDD.n312 185
R14966 VDD.n2068 VDD.n318 185
R14967 VDD.n2398 VDD.n318 185
R14968 VDD.n2070 VDD.n2069 185
R14969 VDD.n2069 VDD.n326 185
R14970 VDD.n2071 VDD.n324 185
R14971 VDD.n2392 VDD.n324 185
R14972 VDD.n2073 VDD.n2072 185
R14973 VDD.n2072 VDD.n323 185
R14974 VDD.n2074 VDD.n331 185
R14975 VDD.n2386 VDD.n331 185
R14976 VDD.n2076 VDD.n2075 185
R14977 VDD.n2075 VDD.n330 185
R14978 VDD.n2077 VDD.n337 185
R14979 VDD.n2380 VDD.n337 185
R14980 VDD.n2079 VDD.n2078 185
R14981 VDD.n2078 VDD.n336 185
R14982 VDD.n2080 VDD.n343 185
R14983 VDD.n2374 VDD.n343 185
R14984 VDD.n2082 VDD.n2081 185
R14985 VDD.n2081 VDD.n342 185
R14986 VDD.n2083 VDD.n349 185
R14987 VDD.n2368 VDD.n349 185
R14988 VDD.n2085 VDD.n2084 185
R14989 VDD.n2084 VDD.n348 185
R14990 VDD.n2086 VDD.n355 185
R14991 VDD.n2362 VDD.n355 185
R14992 VDD.n2088 VDD.n2087 185
R14993 VDD.n2087 VDD.n354 185
R14994 VDD.n2089 VDD.n361 185
R14995 VDD.n2356 VDD.n361 185
R14996 VDD.n2091 VDD.n2090 185
R14997 VDD.n2090 VDD.n360 185
R14998 VDD.n2092 VDD.n367 185
R14999 VDD.n2350 VDD.n367 185
R15000 VDD.n2094 VDD.n2093 185
R15001 VDD.n2093 VDD.n366 185
R15002 VDD.n2095 VDD.n373 185
R15003 VDD.n2344 VDD.n373 185
R15004 VDD.n2097 VDD.n2096 185
R15005 VDD.n2096 VDD.n372 185
R15006 VDD.n2098 VDD.n378 185
R15007 VDD.n2338 VDD.n378 185
R15008 VDD.n2100 VDD.n2099 185
R15009 VDD.n2099 VDD.n385 185
R15010 VDD.n2101 VDD.n383 185
R15011 VDD.n2332 VDD.n383 185
R15012 VDD.n2103 VDD.n2102 185
R15013 VDD.n2102 VDD.n392 185
R15014 VDD.n2104 VDD.n390 185
R15015 VDD.n2326 VDD.n390 185
R15016 VDD.n2106 VDD.n2105 185
R15017 VDD.n2105 VDD.n389 185
R15018 VDD.n2107 VDD.n397 185
R15019 VDD.n2320 VDD.n397 185
R15020 VDD.n2109 VDD.n2108 185
R15021 VDD.n2108 VDD.n396 185
R15022 VDD.n2110 VDD.n403 185
R15023 VDD.n2314 VDD.n403 185
R15024 VDD.n2112 VDD.n2111 185
R15025 VDD.n2111 VDD.n402 185
R15026 VDD.n2113 VDD.n409 185
R15027 VDD.n2308 VDD.n409 185
R15028 VDD.n2115 VDD.n2114 185
R15029 VDD.n2114 VDD.n408 185
R15030 VDD.n2116 VDD.n415 185
R15031 VDD.n2302 VDD.n415 185
R15032 VDD.n2118 VDD.n2117 185
R15033 VDD.n2117 VDD.n414 185
R15034 VDD.n2119 VDD.n421 185
R15035 VDD.n2296 VDD.n421 185
R15036 VDD.n2121 VDD.n2120 185
R15037 VDD.n2120 VDD.n420 185
R15038 VDD.n2122 VDD.n426 185
R15039 VDD.n2290 VDD.n426 185
R15040 VDD.n2124 VDD.n2123 185
R15041 VDD.n2123 VDD.n434 185
R15042 VDD.n2125 VDD.n432 185
R15043 VDD.n2284 VDD.n432 185
R15044 VDD.n2127 VDD.n2126 185
R15045 VDD.n2126 VDD.n431 185
R15046 VDD.n2128 VDD.n439 185
R15047 VDD.n2278 VDD.n439 185
R15048 VDD.n2130 VDD.n2129 185
R15049 VDD.n2129 VDD.n438 185
R15050 VDD.n2131 VDD.n445 185
R15051 VDD.n2272 VDD.n445 185
R15052 VDD.n2133 VDD.n2132 185
R15053 VDD.n2132 VDD.n444 185
R15054 VDD.n2134 VDD.n451 185
R15055 VDD.n2266 VDD.n451 185
R15056 VDD.n2136 VDD.n2135 185
R15057 VDD.n2135 VDD.n450 185
R15058 VDD.n2137 VDD.n457 185
R15059 VDD.n2260 VDD.n457 185
R15060 VDD.n2139 VDD.n2138 185
R15061 VDD.n2138 VDD.n456 185
R15062 VDD.n2140 VDD.n463 185
R15063 VDD.n2254 VDD.n463 185
R15064 VDD.n2142 VDD.n2141 185
R15065 VDD.n2141 VDD.n462 185
R15066 VDD.n2143 VDD.n469 185
R15067 VDD.n2248 VDD.n469 185
R15068 VDD.n2145 VDD.n2144 185
R15069 VDD.n2144 VDD.n468 185
R15070 VDD.n2146 VDD.n475 185
R15071 VDD.n2242 VDD.n475 185
R15072 VDD.n2148 VDD.n2147 185
R15073 VDD.n2147 VDD.n474 185
R15074 VDD.n2149 VDD.n481 185
R15075 VDD.n2236 VDD.n481 185
R15076 VDD.n2151 VDD.n2150 185
R15077 VDD.n2150 VDD.n480 185
R15078 VDD.n2152 VDD.n486 185
R15079 VDD.n2230 VDD.n486 185
R15080 VDD.n2154 VDD.n2153 185
R15081 VDD.n2153 VDD.n494 185
R15082 VDD.n2155 VDD.n492 185
R15083 VDD.n2224 VDD.n492 185
R15084 VDD.n2157 VDD.n2156 185
R15085 VDD.n2156 VDD.n491 185
R15086 VDD.n2158 VDD.n499 185
R15087 VDD.n2218 VDD.n499 185
R15088 VDD.n2160 VDD.n2159 185
R15089 VDD.n2159 VDD.n498 185
R15090 VDD.n2161 VDD.n505 185
R15091 VDD.n2212 VDD.n505 185
R15092 VDD.n2163 VDD.n2162 185
R15093 VDD.n2162 VDD.n504 185
R15094 VDD.n2164 VDD.n511 185
R15095 VDD.n2206 VDD.n511 185
R15096 VDD.n2166 VDD.n2165 185
R15097 VDD.n2165 VDD.n510 185
R15098 VDD.n2167 VDD.n1897 185
R15099 VDD.n2200 VDD.n1897 185
R15100 VDD.n2199 VDD.n2198 185
R15101 VDD.n2200 VDD.n2199 185
R15102 VDD.n509 VDD.n508 185
R15103 VDD.n510 VDD.n509 185
R15104 VDD.n2208 VDD.n2207 185
R15105 VDD.n2207 VDD.n2206 185
R15106 VDD.n2209 VDD.n507 185
R15107 VDD.n507 VDD.n504 185
R15108 VDD.n2211 VDD.n2210 185
R15109 VDD.n2212 VDD.n2211 185
R15110 VDD.n497 VDD.n496 185
R15111 VDD.n498 VDD.n497 185
R15112 VDD.n2220 VDD.n2219 185
R15113 VDD.n2219 VDD.n2218 185
R15114 VDD.n2221 VDD.n495 185
R15115 VDD.n495 VDD.n491 185
R15116 VDD.n2223 VDD.n2222 185
R15117 VDD.n2224 VDD.n2223 185
R15118 VDD.n485 VDD.n484 185
R15119 VDD.n494 VDD.n485 185
R15120 VDD.n2232 VDD.n2231 185
R15121 VDD.n2231 VDD.n2230 185
R15122 VDD.n2233 VDD.n483 185
R15123 VDD.n483 VDD.n480 185
R15124 VDD.n2235 VDD.n2234 185
R15125 VDD.n2236 VDD.n2235 185
R15126 VDD.n473 VDD.n472 185
R15127 VDD.n474 VDD.n473 185
R15128 VDD.n2244 VDD.n2243 185
R15129 VDD.n2243 VDD.n2242 185
R15130 VDD.n2245 VDD.n471 185
R15131 VDD.n471 VDD.n468 185
R15132 VDD.n2247 VDD.n2246 185
R15133 VDD.n2248 VDD.n2247 185
R15134 VDD.n461 VDD.n460 185
R15135 VDD.n462 VDD.n461 185
R15136 VDD.n2256 VDD.n2255 185
R15137 VDD.n2255 VDD.n2254 185
R15138 VDD.n2257 VDD.n459 185
R15139 VDD.n459 VDD.n456 185
R15140 VDD.n2259 VDD.n2258 185
R15141 VDD.n2260 VDD.n2259 185
R15142 VDD.n449 VDD.n448 185
R15143 VDD.n450 VDD.n449 185
R15144 VDD.n2268 VDD.n2267 185
R15145 VDD.n2267 VDD.n2266 185
R15146 VDD.n2269 VDD.n447 185
R15147 VDD.n447 VDD.n444 185
R15148 VDD.n2271 VDD.n2270 185
R15149 VDD.n2272 VDD.n2271 185
R15150 VDD.n437 VDD.n436 185
R15151 VDD.n438 VDD.n437 185
R15152 VDD.n2280 VDD.n2279 185
R15153 VDD.n2279 VDD.n2278 185
R15154 VDD.n2281 VDD.n435 185
R15155 VDD.n435 VDD.n431 185
R15156 VDD.n2283 VDD.n2282 185
R15157 VDD.n2284 VDD.n2283 185
R15158 VDD.n425 VDD.n424 185
R15159 VDD.n434 VDD.n425 185
R15160 VDD.n2292 VDD.n2291 185
R15161 VDD.n2291 VDD.n2290 185
R15162 VDD.n2293 VDD.n423 185
R15163 VDD.n423 VDD.n420 185
R15164 VDD.n2295 VDD.n2294 185
R15165 VDD.n2296 VDD.n2295 185
R15166 VDD.n413 VDD.n412 185
R15167 VDD.n414 VDD.n413 185
R15168 VDD.n2304 VDD.n2303 185
R15169 VDD.n2303 VDD.n2302 185
R15170 VDD.n2305 VDD.n411 185
R15171 VDD.n411 VDD.n408 185
R15172 VDD.n2307 VDD.n2306 185
R15173 VDD.n2308 VDD.n2307 185
R15174 VDD.n401 VDD.n400 185
R15175 VDD.n402 VDD.n401 185
R15176 VDD.n2316 VDD.n2315 185
R15177 VDD.n2315 VDD.n2314 185
R15178 VDD.n2317 VDD.n399 185
R15179 VDD.n399 VDD.n396 185
R15180 VDD.n2319 VDD.n2318 185
R15181 VDD.n2320 VDD.n2319 185
R15182 VDD.n388 VDD.n387 185
R15183 VDD.n389 VDD.n388 185
R15184 VDD.n2328 VDD.n2327 185
R15185 VDD.n2327 VDD.n2326 185
R15186 VDD.n2329 VDD.n386 185
R15187 VDD.n392 VDD.n386 185
R15188 VDD.n2331 VDD.n2330 185
R15189 VDD.n2332 VDD.n2331 185
R15190 VDD.n377 VDD.n376 185
R15191 VDD.n385 VDD.n377 185
R15192 VDD.n2340 VDD.n2339 185
R15193 VDD.n2339 VDD.n2338 185
R15194 VDD.n2341 VDD.n375 185
R15195 VDD.n375 VDD.n372 185
R15196 VDD.n2343 VDD.n2342 185
R15197 VDD.n2344 VDD.n2343 185
R15198 VDD.n365 VDD.n364 185
R15199 VDD.n366 VDD.n365 185
R15200 VDD.n2352 VDD.n2351 185
R15201 VDD.n2351 VDD.n2350 185
R15202 VDD.n2353 VDD.n363 185
R15203 VDD.n363 VDD.n360 185
R15204 VDD.n2355 VDD.n2354 185
R15205 VDD.n2356 VDD.n2355 185
R15206 VDD.n353 VDD.n352 185
R15207 VDD.n354 VDD.n353 185
R15208 VDD.n2364 VDD.n2363 185
R15209 VDD.n2363 VDD.n2362 185
R15210 VDD.n2365 VDD.n351 185
R15211 VDD.n351 VDD.n348 185
R15212 VDD.n2367 VDD.n2366 185
R15213 VDD.n2368 VDD.n2367 185
R15214 VDD.n341 VDD.n340 185
R15215 VDD.n342 VDD.n341 185
R15216 VDD.n2376 VDD.n2375 185
R15217 VDD.n2375 VDD.n2374 185
R15218 VDD.n2377 VDD.n339 185
R15219 VDD.n339 VDD.n336 185
R15220 VDD.n2379 VDD.n2378 185
R15221 VDD.n2380 VDD.n2379 185
R15222 VDD.n329 VDD.n328 185
R15223 VDD.n330 VDD.n329 185
R15224 VDD.n2388 VDD.n2387 185
R15225 VDD.n2387 VDD.n2386 185
R15226 VDD.n2389 VDD.n327 185
R15227 VDD.n327 VDD.n323 185
R15228 VDD.n2391 VDD.n2390 185
R15229 VDD.n2392 VDD.n2391 185
R15230 VDD.n317 VDD.n316 185
R15231 VDD.n326 VDD.n317 185
R15232 VDD.n2400 VDD.n2399 185
R15233 VDD.n2399 VDD.n2398 185
R15234 VDD.n2401 VDD.n315 185
R15235 VDD.n315 VDD.n312 185
R15236 VDD.n2403 VDD.n2402 185
R15237 VDD.n2404 VDD.n2403 185
R15238 VDD.n304 VDD.n303 185
R15239 VDD.n305 VDD.n304 185
R15240 VDD.n2437 VDD.n2436 185
R15241 VDD.n2436 VDD.n2435 185
R15242 VDD.n2438 VDD.n302 185
R15243 VDD.n302 VDD.n299 185
R15244 VDD.n2440 VDD.n2439 185
R15245 VDD.n2441 VDD.n2440 185
R15246 VDD.n284 VDD.n282 185
R15247 VDD.n282 VDD.n278 185
R15248 VDD.n2481 VDD.n2480 185
R15249 VDD.n2482 VDD.n2481 185
R15250 VDD.n2479 VDD.n283 185
R15251 VDD.n283 VDD.n280 185
R15252 VDD.n1554 VDD.n1553 185
R15253 VDD.n1553 VDD.n1552 185
R15254 VDD.n1079 VDD.n1074 185
R15255 VDD.n1558 VDD.n1073 185
R15256 VDD.n1559 VDD.n1072 185
R15257 VDD.n1560 VDD.n1071 185
R15258 VDD.n1548 VDD.n1069 185
R15259 VDD.n1564 VDD.n1068 185
R15260 VDD.n1565 VDD.n1067 185
R15261 VDD.n1566 VDD.n1066 185
R15262 VDD.n1545 VDD.n1064 185
R15263 VDD.n1570 VDD.n1061 185
R15264 VDD.n1571 VDD.n1060 185
R15265 VDD.n1572 VDD.n1059 185
R15266 VDD.n1542 VDD.n1058 185
R15267 VDD.n1541 VDD.n1540 185
R15268 VDD.n1088 VDD.n1087 185
R15269 VDD.n1536 VDD.n1535 185
R15270 VDD.n1534 VDD.n1533 185
R15271 VDD.n1532 VDD.n1531 185
R15272 VDD.n1530 VDD.n1090 185
R15273 VDD.n1526 VDD.n1525 185
R15274 VDD.n1524 VDD.n1523 185
R15275 VDD.n1522 VDD.n1096 185
R15276 VDD.n1095 VDD.n1094 185
R15277 VDD.n1518 VDD.n1517 185
R15278 VDD.n1105 VDD.n1080 185
R15279 VDD.n1081 VDD.n1080 185
R15280 VDD.n1507 VDD.n1506 185
R15281 VDD.n1508 VDD.n1507 185
R15282 VDD.n1104 VDD.n1103 185
R15283 VDD.n1509 VDD.n1103 185
R15284 VDD.n1501 VDD.n1500 185
R15285 VDD.n1500 VDD.n1102 185
R15286 VDD.n1499 VDD.n1107 185
R15287 VDD.n1499 VDD.n1498 185
R15288 VDD.n1118 VDD.n1108 185
R15289 VDD.n1109 VDD.n1108 185
R15290 VDD.n1489 VDD.n1488 185
R15291 VDD.n1490 VDD.n1489 185
R15292 VDD.n1117 VDD.n1116 185
R15293 VDD.n1116 VDD.n1115 185
R15294 VDD.n1483 VDD.n1482 185
R15295 VDD.n1482 VDD.n1481 185
R15296 VDD.n1121 VDD.n1120 185
R15297 VDD.n1122 VDD.n1121 185
R15298 VDD.n1472 VDD.n1471 185
R15299 VDD.n1473 VDD.n1472 185
R15300 VDD.n1130 VDD.n1129 185
R15301 VDD.n1129 VDD.n1128 185
R15302 VDD.n1467 VDD.n1466 185
R15303 VDD.n1466 VDD.n1465 185
R15304 VDD.n1133 VDD.n1132 185
R15305 VDD.n1456 VDD.n1133 185
R15306 VDD.n1455 VDD.n1454 185
R15307 VDD.n1457 VDD.n1455 185
R15308 VDD.n1141 VDD.n1140 185
R15309 VDD.n1140 VDD.n1139 185
R15310 VDD.n1450 VDD.n1449 185
R15311 VDD.n1449 VDD.n1448 185
R15312 VDD.n1144 VDD.n1143 185
R15313 VDD.n1145 VDD.n1144 185
R15314 VDD.n1439 VDD.n1438 185
R15315 VDD.n1440 VDD.n1439 185
R15316 VDD.n1152 VDD.n1151 185
R15317 VDD.n1157 VDD.n1151 185
R15318 VDD.n1434 VDD.n1433 185
R15319 VDD.n1433 VDD.n1432 185
R15320 VDD.n1155 VDD.n1154 185
R15321 VDD.n1156 VDD.n1155 185
R15322 VDD.n1411 VDD.n1410 185
R15323 VDD.n1412 VDD.n1411 185
R15324 VDD.n1165 VDD.n1164 185
R15325 VDD.n1164 VDD.n1163 185
R15326 VDD.n1406 VDD.n1405 185
R15327 VDD.n1405 VDD.n1404 185
R15328 VDD.n1168 VDD.n1167 185
R15329 VDD.n1169 VDD.n1168 185
R15330 VDD.n1395 VDD.n1394 185
R15331 VDD.n1396 VDD.n1395 185
R15332 VDD.n1177 VDD.n1176 185
R15333 VDD.n1176 VDD.n1175 185
R15334 VDD.n1390 VDD.n1389 185
R15335 VDD.n1389 VDD.n1388 185
R15336 VDD.n1180 VDD.n1179 185
R15337 VDD.n1181 VDD.n1180 185
R15338 VDD.n1379 VDD.n1378 185
R15339 VDD.n1380 VDD.n1379 185
R15340 VDD.n1189 VDD.n1188 185
R15341 VDD.n1188 VDD.n1187 185
R15342 VDD.n1374 VDD.n1373 185
R15343 VDD.n1373 VDD.n1372 185
R15344 VDD.n1192 VDD.n1191 185
R15345 VDD.n1193 VDD.n1192 185
R15346 VDD.n1363 VDD.n1362 185
R15347 VDD.n1364 VDD.n1363 185
R15348 VDD.n1201 VDD.n1200 185
R15349 VDD.n1200 VDD.n1199 185
R15350 VDD.n1358 VDD.n1357 185
R15351 VDD.n1357 VDD.n1356 185
R15352 VDD.n1204 VDD.n1203 185
R15353 VDD.n1205 VDD.n1204 185
R15354 VDD.n1347 VDD.n1346 185
R15355 VDD.n1348 VDD.n1347 185
R15356 VDD.n1213 VDD.n1212 185
R15357 VDD.n1212 VDD.n1211 185
R15358 VDD.n1342 VDD.n1341 185
R15359 VDD.n1341 VDD.n1340 185
R15360 VDD.n1216 VDD.n1215 185
R15361 VDD.n1331 VDD.n1216 185
R15362 VDD.n1330 VDD.n1329 185
R15363 VDD.n1332 VDD.n1330 185
R15364 VDD.n1224 VDD.n1223 185
R15365 VDD.n1223 VDD.n1222 185
R15366 VDD.n1325 VDD.n1324 185
R15367 VDD.n1324 VDD.n1323 185
R15368 VDD.n1318 VDD.n1228 185
R15369 VDD.n1317 VDD.n1231 185
R15370 VDD.n1316 VDD.n1232 185
R15371 VDD.n1232 VDD.n1227 185
R15372 VDD.n1235 VDD.n1233 185
R15373 VDD.n1312 VDD.n1237 185
R15374 VDD.n1311 VDD.n1238 185
R15375 VDD.n1310 VDD.n1307 185
R15376 VDD.n1305 VDD.n1239 185
R15377 VDD.n1303 VDD.n1302 185
R15378 VDD.n1242 VDD.n1241 185
R15379 VDD.n1298 VDD.n1246 185
R15380 VDD.n1297 VDD.n1247 185
R15381 VDD.n1296 VDD.n1249 185
R15382 VDD.n1252 VDD.n1250 185
R15383 VDD.n1292 VDD.n1254 185
R15384 VDD.n1291 VDD.n1288 185
R15385 VDD.n1286 VDD.n1255 185
R15386 VDD.n1285 VDD.n1284 185
R15387 VDD.n1260 VDD.n1257 185
R15388 VDD.n1280 VDD.n1261 185
R15389 VDD.n1279 VDD.n1263 185
R15390 VDD.n1278 VDD.n1264 185
R15391 VDD.n1267 VDD.n1265 185
R15392 VDD.n1274 VDD.n1269 185
R15393 VDD.n1270 VDD.n1226 185
R15394 VDD.n1516 VDD.n1515 185
R15395 VDD.n1516 VDD.n1081 185
R15396 VDD.n1098 VDD.n1097 185
R15397 VDD.n1508 VDD.n1097 185
R15398 VDD.n1511 VDD.n1510 185
R15399 VDD.n1510 VDD.n1509 185
R15400 VDD.n1101 VDD.n1100 185
R15401 VDD.n1102 VDD.n1101 185
R15402 VDD.n1497 VDD.n1496 185
R15403 VDD.n1498 VDD.n1497 185
R15404 VDD.n1111 VDD.n1110 185
R15405 VDD.n1110 VDD.n1109 185
R15406 VDD.n1492 VDD.n1491 185
R15407 VDD.n1491 VDD.n1490 185
R15408 VDD.n1114 VDD.n1113 185
R15409 VDD.n1115 VDD.n1114 185
R15410 VDD.n1480 VDD.n1479 185
R15411 VDD.n1481 VDD.n1480 185
R15412 VDD.n1124 VDD.n1123 185
R15413 VDD.n1123 VDD.n1122 185
R15414 VDD.n1475 VDD.n1474 185
R15415 VDD.n1474 VDD.n1473 185
R15416 VDD.n1127 VDD.n1126 185
R15417 VDD.n1128 VDD.n1127 185
R15418 VDD.n1464 VDD.n1463 185
R15419 VDD.n1465 VDD.n1464 185
R15420 VDD.n1135 VDD.n1134 185
R15421 VDD.n1456 VDD.n1134 185
R15422 VDD.n1459 VDD.n1458 185
R15423 VDD.n1458 VDD.n1457 185
R15424 VDD.n1138 VDD.n1137 185
R15425 VDD.n1139 VDD.n1138 185
R15426 VDD.n1447 VDD.n1446 185
R15427 VDD.n1448 VDD.n1447 185
R15428 VDD.n1147 VDD.n1146 185
R15429 VDD.n1146 VDD.n1145 185
R15430 VDD.n1442 VDD.n1441 185
R15431 VDD.n1441 VDD.n1440 185
R15432 VDD.n1150 VDD.n1149 185
R15433 VDD.n1157 VDD.n1150 185
R15434 VDD.n1431 VDD.n1430 185
R15435 VDD.n1432 VDD.n1431 185
R15436 VDD.n1159 VDD.n1158 185
R15437 VDD.n1158 VDD.n1156 185
R15438 VDD.n1414 VDD.n1413 185
R15439 VDD.n1413 VDD.n1412 185
R15440 VDD.n1162 VDD.n1161 185
R15441 VDD.n1163 VDD.n1162 185
R15442 VDD.n1403 VDD.n1402 185
R15443 VDD.n1404 VDD.n1403 185
R15444 VDD.n1171 VDD.n1170 185
R15445 VDD.n1170 VDD.n1169 185
R15446 VDD.n1398 VDD.n1397 185
R15447 VDD.n1397 VDD.n1396 185
R15448 VDD.n1174 VDD.n1173 185
R15449 VDD.n1175 VDD.n1174 185
R15450 VDD.n1387 VDD.n1386 185
R15451 VDD.n1388 VDD.n1387 185
R15452 VDD.n1183 VDD.n1182 185
R15453 VDD.n1182 VDD.n1181 185
R15454 VDD.n1382 VDD.n1381 185
R15455 VDD.n1381 VDD.n1380 185
R15456 VDD.n1186 VDD.n1185 185
R15457 VDD.n1187 VDD.n1186 185
R15458 VDD.n1371 VDD.n1370 185
R15459 VDD.n1372 VDD.n1371 185
R15460 VDD.n1195 VDD.n1194 185
R15461 VDD.n1194 VDD.n1193 185
R15462 VDD.n1366 VDD.n1365 185
R15463 VDD.n1365 VDD.n1364 185
R15464 VDD.n1198 VDD.n1197 185
R15465 VDD.n1199 VDD.n1198 185
R15466 VDD.n1355 VDD.n1354 185
R15467 VDD.n1356 VDD.n1355 185
R15468 VDD.n1207 VDD.n1206 185
R15469 VDD.n1206 VDD.n1205 185
R15470 VDD.n1350 VDD.n1349 185
R15471 VDD.n1349 VDD.n1348 185
R15472 VDD.n1210 VDD.n1209 185
R15473 VDD.n1211 VDD.n1210 185
R15474 VDD.n1339 VDD.n1338 185
R15475 VDD.n1340 VDD.n1339 185
R15476 VDD.n1218 VDD.n1217 185
R15477 VDD.n1331 VDD.n1217 185
R15478 VDD.n1334 VDD.n1333 185
R15479 VDD.n1333 VDD.n1332 185
R15480 VDD.n1221 VDD.n1220 185
R15481 VDD.n1222 VDD.n1221 185
R15482 VDD.n1322 VDD.n1321 185
R15483 VDD.n1323 VDD.n1322 185
R15484 VDD.n24 VDD.t137 173.494
R15485 VDD.n20 VDD.t109 173.494
R15486 VDD.n17 VDD.t134 173.494
R15487 VDD.n1423 VDD.t131 173.494
R15488 VDD.n1419 VDD.t135 173.494
R15489 VDD.n1416 VDD.t129 173.494
R15490 VDD.n1272 VDD.t75 171.493
R15491 VDD.n1290 VDD.t84 171.493
R15492 VDD.n1309 VDD.t81 171.493
R15493 VDD.n234 VDD.t68 171.493
R15494 VDD.n248 VDD.t71 171.493
R15495 VDD.n262 VDD.t62 171.493
R15496 VDD.n137 VDD.t41 171.493
R15497 VDD.n123 VDD.t59 171.493
R15498 VDD.n105 VDD.t48 171.493
R15499 VDD.n1092 VDD.t99 171.493
R15500 VDD.n1063 VDD.t102 171.493
R15501 VDD.n1077 VDD.t92 171.493
R15502 VDD.n25 VDD.t112 170.683
R15503 VDD.n21 VDD.t113 170.683
R15504 VDD.n18 VDD.t111 170.683
R15505 VDD.n1424 VDD.t120 170.683
R15506 VDD.n1420 VDD.t121 170.683
R15507 VDD.n1417 VDD.t118 170.683
R15508 VDD.n1896 VDD.n1895 156.466
R15509 VDD.n24 VDD.n23 155.131
R15510 VDD.n20 VDD.n19 155.131
R15511 VDD.n17 VDD.n16 155.131
R15512 VDD.n1423 VDD.n1422 155.131
R15513 VDD.n1419 VDD.n1418 155.131
R15514 VDD.n1416 VDD.n1415 155.131
R15515 VDD.n95 VDD.n92 146.341
R15516 VDD.n2721 VDD.n2720 146.341
R15517 VDD.n2718 VDD.n99 146.341
R15518 VDD.n110 VDD.n107 146.341
R15519 VDD.n2710 VDD.n2709 146.341
R15520 VDD.n2707 VDD.n112 146.341
R15521 VDD.n2703 VDD.n2702 146.341
R15522 VDD.n2700 VDD.n118 146.341
R15523 VDD.n2693 VDD.n127 146.341
R15524 VDD.n2691 VDD.n2690 146.341
R15525 VDD.n2688 VDD.n129 146.341
R15526 VDD.n2684 VDD.n2683 146.341
R15527 VDD.n2559 VDD.n215 146.341
R15528 VDD.n2565 VDD.n215 146.341
R15529 VDD.n2565 VDD.n208 146.341
R15530 VDD.n2576 VDD.n208 146.341
R15531 VDD.n2576 VDD.n204 146.341
R15532 VDD.n2582 VDD.n204 146.341
R15533 VDD.n2582 VDD.n196 146.341
R15534 VDD.n2592 VDD.n196 146.341
R15535 VDD.n2592 VDD.n192 146.341
R15536 VDD.n2598 VDD.n192 146.341
R15537 VDD.n2598 VDD.n184 146.341
R15538 VDD.n2608 VDD.n184 146.341
R15539 VDD.n2608 VDD.n180 146.341
R15540 VDD.n2614 VDD.n180 146.341
R15541 VDD.n2614 VDD.n172 146.341
R15542 VDD.n2624 VDD.n172 146.341
R15543 VDD.n2624 VDD.n168 146.341
R15544 VDD.n2630 VDD.n168 146.341
R15545 VDD.n2630 VDD.n159 146.341
R15546 VDD.n2640 VDD.n159 146.341
R15547 VDD.n2640 VDD.n160 146.341
R15548 VDD.n160 VDD.n34 146.341
R15549 VDD.n35 VDD.n34 146.341
R15550 VDD.n36 VDD.n35 146.341
R15551 VDD.n153 VDD.n36 146.341
R15552 VDD.n153 VDD.n44 146.341
R15553 VDD.n45 VDD.n44 146.341
R15554 VDD.n46 VDD.n45 146.341
R15555 VDD.n150 VDD.n46 146.341
R15556 VDD.n150 VDD.n55 146.341
R15557 VDD.n56 VDD.n55 146.341
R15558 VDD.n57 VDD.n56 146.341
R15559 VDD.n147 VDD.n57 146.341
R15560 VDD.n147 VDD.n66 146.341
R15561 VDD.n67 VDD.n66 146.341
R15562 VDD.n68 VDD.n67 146.341
R15563 VDD.n144 VDD.n68 146.341
R15564 VDD.n144 VDD.n77 146.341
R15565 VDD.n78 VDD.n77 146.341
R15566 VDD.n79 VDD.n78 146.341
R15567 VDD.n141 VDD.n79 146.341
R15568 VDD.n141 VDD.n88 146.341
R15569 VDD.n89 VDD.n88 146.341
R15570 VDD.n90 VDD.n89 146.341
R15571 VDD.n2549 VDD.n2547 146.341
R15572 VDD.n2547 VDD.n2546 146.341
R15573 VDD.n2543 VDD.n2542 146.341
R15574 VDD.n2540 VDD.n230 146.341
R15575 VDD.n2536 VDD.n2534 146.341
R15576 VDD.n2532 VDD.n238 146.341
R15577 VDD.n2528 VDD.n2526 146.341
R15578 VDD.n2524 VDD.n243 146.341
R15579 VDD.n2520 VDD.n2518 146.341
R15580 VDD.n2516 VDD.n251 146.341
R15581 VDD.n2512 VDD.n2510 146.341
R15582 VDD.n2508 VDD.n258 146.341
R15583 VDD.n2557 VDD.n213 146.341
R15584 VDD.n2568 VDD.n213 146.341
R15585 VDD.n2568 VDD.n209 146.341
R15586 VDD.n2574 VDD.n209 146.341
R15587 VDD.n2574 VDD.n202 146.341
R15588 VDD.n2584 VDD.n202 146.341
R15589 VDD.n2584 VDD.n198 146.341
R15590 VDD.n2590 VDD.n198 146.341
R15591 VDD.n2590 VDD.n190 146.341
R15592 VDD.n2600 VDD.n190 146.341
R15593 VDD.n2600 VDD.n186 146.341
R15594 VDD.n2606 VDD.n186 146.341
R15595 VDD.n2606 VDD.n178 146.341
R15596 VDD.n2616 VDD.n178 146.341
R15597 VDD.n2616 VDD.n174 146.341
R15598 VDD.n2622 VDD.n174 146.341
R15599 VDD.n2622 VDD.n166 146.341
R15600 VDD.n2632 VDD.n166 146.341
R15601 VDD.n2632 VDD.n162 146.341
R15602 VDD.n2638 VDD.n162 146.341
R15603 VDD.n2638 VDD.n31 146.341
R15604 VDD.n2772 VDD.n31 146.341
R15605 VDD.n2772 VDD.n32 146.341
R15606 VDD.n2768 VDD.n32 146.341
R15607 VDD.n2768 VDD.n38 146.341
R15608 VDD.n2764 VDD.n38 146.341
R15609 VDD.n2764 VDD.n43 146.341
R15610 VDD.n2760 VDD.n43 146.341
R15611 VDD.n2760 VDD.n48 146.341
R15612 VDD.n2756 VDD.n48 146.341
R15613 VDD.n2756 VDD.n54 146.341
R15614 VDD.n2752 VDD.n54 146.341
R15615 VDD.n2752 VDD.n59 146.341
R15616 VDD.n2748 VDD.n59 146.341
R15617 VDD.n2748 VDD.n65 146.341
R15618 VDD.n2744 VDD.n65 146.341
R15619 VDD.n2744 VDD.n70 146.341
R15620 VDD.n2740 VDD.n70 146.341
R15621 VDD.n2740 VDD.n76 146.341
R15622 VDD.n2736 VDD.n76 146.341
R15623 VDD.n2736 VDD.n80 146.341
R15624 VDD.n2732 VDD.n80 146.341
R15625 VDD.n2732 VDD.n86 146.341
R15626 VDD.n2728 VDD.n86 146.341
R15627 VDD.n1096 VDD.n1095 146.341
R15628 VDD.n1525 VDD.n1524 146.341
R15629 VDD.n1531 VDD.n1530 146.341
R15630 VDD.n1535 VDD.n1534 146.341
R15631 VDD.n1541 VDD.n1087 146.341
R15632 VDD.n1542 VDD.n1059 146.341
R15633 VDD.n1061 VDD.n1060 146.341
R15634 VDD.n1545 VDD.n1066 146.341
R15635 VDD.n1068 VDD.n1067 146.341
R15636 VDD.n1548 VDD.n1071 146.341
R15637 VDD.n1073 VDD.n1072 146.341
R15638 VDD.n1553 VDD.n1079 146.341
R15639 VDD.n1324 VDD.n1223 146.341
R15640 VDD.n1330 VDD.n1223 146.341
R15641 VDD.n1330 VDD.n1216 146.341
R15642 VDD.n1341 VDD.n1216 146.341
R15643 VDD.n1341 VDD.n1212 146.341
R15644 VDD.n1347 VDD.n1212 146.341
R15645 VDD.n1347 VDD.n1204 146.341
R15646 VDD.n1357 VDD.n1204 146.341
R15647 VDD.n1357 VDD.n1200 146.341
R15648 VDD.n1363 VDD.n1200 146.341
R15649 VDD.n1363 VDD.n1192 146.341
R15650 VDD.n1373 VDD.n1192 146.341
R15651 VDD.n1373 VDD.n1188 146.341
R15652 VDD.n1379 VDD.n1188 146.341
R15653 VDD.n1379 VDD.n1180 146.341
R15654 VDD.n1389 VDD.n1180 146.341
R15655 VDD.n1389 VDD.n1176 146.341
R15656 VDD.n1395 VDD.n1176 146.341
R15657 VDD.n1395 VDD.n1168 146.341
R15658 VDD.n1405 VDD.n1168 146.341
R15659 VDD.n1405 VDD.n1164 146.341
R15660 VDD.n1411 VDD.n1164 146.341
R15661 VDD.n1411 VDD.n1155 146.341
R15662 VDD.n1433 VDD.n1155 146.341
R15663 VDD.n1433 VDD.n1151 146.341
R15664 VDD.n1439 VDD.n1151 146.341
R15665 VDD.n1439 VDD.n1144 146.341
R15666 VDD.n1449 VDD.n1144 146.341
R15667 VDD.n1449 VDD.n1140 146.341
R15668 VDD.n1455 VDD.n1140 146.341
R15669 VDD.n1455 VDD.n1133 146.341
R15670 VDD.n1466 VDD.n1133 146.341
R15671 VDD.n1466 VDD.n1129 146.341
R15672 VDD.n1472 VDD.n1129 146.341
R15673 VDD.n1472 VDD.n1121 146.341
R15674 VDD.n1482 VDD.n1121 146.341
R15675 VDD.n1482 VDD.n1116 146.341
R15676 VDD.n1489 VDD.n1116 146.341
R15677 VDD.n1489 VDD.n1108 146.341
R15678 VDD.n1499 VDD.n1108 146.341
R15679 VDD.n1500 VDD.n1499 146.341
R15680 VDD.n1500 VDD.n1103 146.341
R15681 VDD.n1507 VDD.n1103 146.341
R15682 VDD.n1507 VDD.n1080 146.341
R15683 VDD.n1232 VDD.n1231 146.341
R15684 VDD.n1235 VDD.n1232 146.341
R15685 VDD.n1238 VDD.n1237 146.341
R15686 VDD.n1307 VDD.n1305 146.341
R15687 VDD.n1303 VDD.n1241 146.341
R15688 VDD.n1247 VDD.n1246 146.341
R15689 VDD.n1252 VDD.n1249 146.341
R15690 VDD.n1288 VDD.n1254 146.341
R15691 VDD.n1286 VDD.n1285 146.341
R15692 VDD.n1261 VDD.n1260 146.341
R15693 VDD.n1264 VDD.n1263 146.341
R15694 VDD.n1269 VDD.n1267 146.341
R15695 VDD.n1322 VDD.n1221 146.341
R15696 VDD.n1333 VDD.n1221 146.341
R15697 VDD.n1333 VDD.n1217 146.341
R15698 VDD.n1339 VDD.n1217 146.341
R15699 VDD.n1339 VDD.n1210 146.341
R15700 VDD.n1349 VDD.n1210 146.341
R15701 VDD.n1349 VDD.n1206 146.341
R15702 VDD.n1355 VDD.n1206 146.341
R15703 VDD.n1355 VDD.n1198 146.341
R15704 VDD.n1365 VDD.n1198 146.341
R15705 VDD.n1365 VDD.n1194 146.341
R15706 VDD.n1371 VDD.n1194 146.341
R15707 VDD.n1371 VDD.n1186 146.341
R15708 VDD.n1381 VDD.n1186 146.341
R15709 VDD.n1381 VDD.n1182 146.341
R15710 VDD.n1387 VDD.n1182 146.341
R15711 VDD.n1387 VDD.n1174 146.341
R15712 VDD.n1397 VDD.n1174 146.341
R15713 VDD.n1397 VDD.n1170 146.341
R15714 VDD.n1403 VDD.n1170 146.341
R15715 VDD.n1403 VDD.n1162 146.341
R15716 VDD.n1413 VDD.n1162 146.341
R15717 VDD.n1413 VDD.n1158 146.341
R15718 VDD.n1431 VDD.n1158 146.341
R15719 VDD.n1431 VDD.n1150 146.341
R15720 VDD.n1441 VDD.n1150 146.341
R15721 VDD.n1441 VDD.n1146 146.341
R15722 VDD.n1447 VDD.n1146 146.341
R15723 VDD.n1447 VDD.n1138 146.341
R15724 VDD.n1458 VDD.n1138 146.341
R15725 VDD.n1458 VDD.n1134 146.341
R15726 VDD.n1464 VDD.n1134 146.341
R15727 VDD.n1464 VDD.n1127 146.341
R15728 VDD.n1474 VDD.n1127 146.341
R15729 VDD.n1474 VDD.n1123 146.341
R15730 VDD.n1480 VDD.n1123 146.341
R15731 VDD.n1480 VDD.n1114 146.341
R15732 VDD.n1491 VDD.n1114 146.341
R15733 VDD.n1491 VDD.n1110 146.341
R15734 VDD.n1497 VDD.n1110 146.341
R15735 VDD.n1497 VDD.n1101 146.341
R15736 VDD.n1510 VDD.n1101 146.341
R15737 VDD.n1510 VDD.n1097 146.341
R15738 VDD.n1516 VDD.n1097 146.341
R15739 VDD.n9 VDD.n7 137.216
R15740 VDD.n2 VDD.n0 137.216
R15741 VDD.n9 VDD.n8 132.311
R15742 VDD.n11 VDD.n10 132.311
R15743 VDD.n13 VDD.n12 132.311
R15744 VDD.n6 VDD.n5 132.311
R15745 VDD.n4 VDD.n3 132.311
R15746 VDD.n2 VDD.n1 132.311
R15747 VDD.t18 VDD.n764 125.431
R15748 VDD.n267 VDD.t10 125.431
R15749 VDD.n1901 VDD.n1900 110.353
R15750 VDD.n296 VDD.n295 110.353
R15751 VDD.n2059 VDD.n2058 110.353
R15752 VDD.n271 VDD.n270 110.353
R15753 VDD.n797 VDD.n796 110.353
R15754 VDD.n822 VDD.n821 110.353
R15755 VDD.n544 VDD.n543 110.353
R15756 VDD.n1801 VDD.n1800 110.353
R15757 VDD.n2199 VDD.n509 99.5127
R15758 VDD.n2207 VDD.n509 99.5127
R15759 VDD.n2207 VDD.n507 99.5127
R15760 VDD.n2211 VDD.n507 99.5127
R15761 VDD.n2211 VDD.n497 99.5127
R15762 VDD.n2219 VDD.n497 99.5127
R15763 VDD.n2219 VDD.n495 99.5127
R15764 VDD.n2223 VDD.n495 99.5127
R15765 VDD.n2223 VDD.n485 99.5127
R15766 VDD.n2231 VDD.n485 99.5127
R15767 VDD.n2231 VDD.n483 99.5127
R15768 VDD.n2235 VDD.n483 99.5127
R15769 VDD.n2235 VDD.n473 99.5127
R15770 VDD.n2243 VDD.n473 99.5127
R15771 VDD.n2243 VDD.n471 99.5127
R15772 VDD.n2247 VDD.n471 99.5127
R15773 VDD.n2247 VDD.n461 99.5127
R15774 VDD.n2255 VDD.n461 99.5127
R15775 VDD.n2255 VDD.n459 99.5127
R15776 VDD.n2259 VDD.n459 99.5127
R15777 VDD.n2259 VDD.n449 99.5127
R15778 VDD.n2267 VDD.n449 99.5127
R15779 VDD.n2267 VDD.n447 99.5127
R15780 VDD.n2271 VDD.n447 99.5127
R15781 VDD.n2271 VDD.n437 99.5127
R15782 VDD.n2279 VDD.n437 99.5127
R15783 VDD.n2279 VDD.n435 99.5127
R15784 VDD.n2283 VDD.n435 99.5127
R15785 VDD.n2283 VDD.n425 99.5127
R15786 VDD.n2291 VDD.n425 99.5127
R15787 VDD.n2291 VDD.n423 99.5127
R15788 VDD.n2295 VDD.n423 99.5127
R15789 VDD.n2295 VDD.n413 99.5127
R15790 VDD.n2303 VDD.n413 99.5127
R15791 VDD.n2303 VDD.n411 99.5127
R15792 VDD.n2307 VDD.n411 99.5127
R15793 VDD.n2307 VDD.n401 99.5127
R15794 VDD.n2315 VDD.n401 99.5127
R15795 VDD.n2315 VDD.n399 99.5127
R15796 VDD.n2319 VDD.n399 99.5127
R15797 VDD.n2319 VDD.n388 99.5127
R15798 VDD.n2327 VDD.n388 99.5127
R15799 VDD.n2327 VDD.n386 99.5127
R15800 VDD.n2331 VDD.n386 99.5127
R15801 VDD.n2331 VDD.n377 99.5127
R15802 VDD.n2339 VDD.n377 99.5127
R15803 VDD.n2339 VDD.n375 99.5127
R15804 VDD.n2343 VDD.n375 99.5127
R15805 VDD.n2343 VDD.n365 99.5127
R15806 VDD.n2351 VDD.n365 99.5127
R15807 VDD.n2351 VDD.n363 99.5127
R15808 VDD.n2355 VDD.n363 99.5127
R15809 VDD.n2355 VDD.n353 99.5127
R15810 VDD.n2363 VDD.n353 99.5127
R15811 VDD.n2363 VDD.n351 99.5127
R15812 VDD.n2367 VDD.n351 99.5127
R15813 VDD.n2367 VDD.n341 99.5127
R15814 VDD.n2375 VDD.n341 99.5127
R15815 VDD.n2375 VDD.n339 99.5127
R15816 VDD.n2379 VDD.n339 99.5127
R15817 VDD.n2379 VDD.n329 99.5127
R15818 VDD.n2387 VDD.n329 99.5127
R15819 VDD.n2387 VDD.n327 99.5127
R15820 VDD.n2391 VDD.n327 99.5127
R15821 VDD.n2391 VDD.n317 99.5127
R15822 VDD.n2399 VDD.n317 99.5127
R15823 VDD.n2399 VDD.n315 99.5127
R15824 VDD.n2403 VDD.n315 99.5127
R15825 VDD.n2403 VDD.n304 99.5127
R15826 VDD.n2436 VDD.n304 99.5127
R15827 VDD.n2436 VDD.n302 99.5127
R15828 VDD.n2440 VDD.n302 99.5127
R15829 VDD.n2440 VDD.n282 99.5127
R15830 VDD.n2481 VDD.n282 99.5127
R15831 VDD.n2481 VDD.n283 99.5127
R15832 VDD.n2475 VDD.n2474 99.5127
R15833 VDD.n2472 VDD.n287 99.5127
R15834 VDD.n2468 VDD.n2467 99.5127
R15835 VDD.n2465 VDD.n2463 99.5127
R15836 VDD.n2461 VDD.n291 99.5127
R15837 VDD.n2457 VDD.n2456 99.5127
R15838 VDD.n2454 VDD.n294 99.5127
R15839 VDD.n2165 VDD.n1897 99.5127
R15840 VDD.n2165 VDD.n511 99.5127
R15841 VDD.n2162 VDD.n511 99.5127
R15842 VDD.n2162 VDD.n505 99.5127
R15843 VDD.n2159 VDD.n505 99.5127
R15844 VDD.n2159 VDD.n499 99.5127
R15845 VDD.n2156 VDD.n499 99.5127
R15846 VDD.n2156 VDD.n492 99.5127
R15847 VDD.n2153 VDD.n492 99.5127
R15848 VDD.n2153 VDD.n486 99.5127
R15849 VDD.n2150 VDD.n486 99.5127
R15850 VDD.n2150 VDD.n481 99.5127
R15851 VDD.n2147 VDD.n481 99.5127
R15852 VDD.n2147 VDD.n475 99.5127
R15853 VDD.n2144 VDD.n475 99.5127
R15854 VDD.n2144 VDD.n469 99.5127
R15855 VDD.n2141 VDD.n469 99.5127
R15856 VDD.n2141 VDD.n463 99.5127
R15857 VDD.n2138 VDD.n463 99.5127
R15858 VDD.n2138 VDD.n457 99.5127
R15859 VDD.n2135 VDD.n457 99.5127
R15860 VDD.n2135 VDD.n451 99.5127
R15861 VDD.n2132 VDD.n451 99.5127
R15862 VDD.n2132 VDD.n445 99.5127
R15863 VDD.n2129 VDD.n445 99.5127
R15864 VDD.n2129 VDD.n439 99.5127
R15865 VDD.n2126 VDD.n439 99.5127
R15866 VDD.n2126 VDD.n432 99.5127
R15867 VDD.n2123 VDD.n432 99.5127
R15868 VDD.n2123 VDD.n426 99.5127
R15869 VDD.n2120 VDD.n426 99.5127
R15870 VDD.n2120 VDD.n421 99.5127
R15871 VDD.n2117 VDD.n421 99.5127
R15872 VDD.n2117 VDD.n415 99.5127
R15873 VDD.n2114 VDD.n415 99.5127
R15874 VDD.n2114 VDD.n409 99.5127
R15875 VDD.n2111 VDD.n409 99.5127
R15876 VDD.n2111 VDD.n403 99.5127
R15877 VDD.n2108 VDD.n403 99.5127
R15878 VDD.n2108 VDD.n397 99.5127
R15879 VDD.n2105 VDD.n397 99.5127
R15880 VDD.n2105 VDD.n390 99.5127
R15881 VDD.n2102 VDD.n390 99.5127
R15882 VDD.n2102 VDD.n383 99.5127
R15883 VDD.n2099 VDD.n383 99.5127
R15884 VDD.n2099 VDD.n378 99.5127
R15885 VDD.n2096 VDD.n378 99.5127
R15886 VDD.n2096 VDD.n373 99.5127
R15887 VDD.n2093 VDD.n373 99.5127
R15888 VDD.n2093 VDD.n367 99.5127
R15889 VDD.n2090 VDD.n367 99.5127
R15890 VDD.n2090 VDD.n361 99.5127
R15891 VDD.n2087 VDD.n361 99.5127
R15892 VDD.n2087 VDD.n355 99.5127
R15893 VDD.n2084 VDD.n355 99.5127
R15894 VDD.n2084 VDD.n349 99.5127
R15895 VDD.n2081 VDD.n349 99.5127
R15896 VDD.n2081 VDD.n343 99.5127
R15897 VDD.n2078 VDD.n343 99.5127
R15898 VDD.n2078 VDD.n337 99.5127
R15899 VDD.n2075 VDD.n337 99.5127
R15900 VDD.n2075 VDD.n331 99.5127
R15901 VDD.n2072 VDD.n331 99.5127
R15902 VDD.n2072 VDD.n324 99.5127
R15903 VDD.n2069 VDD.n324 99.5127
R15904 VDD.n2069 VDD.n318 99.5127
R15905 VDD.n2066 VDD.n318 99.5127
R15906 VDD.n2066 VDD.n313 99.5127
R15907 VDD.n2063 VDD.n313 99.5127
R15908 VDD.n2063 VDD.n306 99.5127
R15909 VDD.n306 VDD.n298 99.5127
R15910 VDD.n2442 VDD.n298 99.5127
R15911 VDD.n2443 VDD.n2442 99.5127
R15912 VDD.n2443 VDD.n279 99.5127
R15913 VDD.n2448 VDD.n279 99.5127
R15914 VDD.n2195 VDD.n2193 99.5127
R15915 VDD.n2193 VDD.n2192 99.5127
R15916 VDD.n2189 VDD.n2188 99.5127
R15917 VDD.n2186 VDD.n2053 99.5127
R15918 VDD.n2182 VDD.n2180 99.5127
R15919 VDD.n2178 VDD.n2055 99.5127
R15920 VDD.n2174 VDD.n2172 99.5127
R15921 VDD.n2170 VDD.n2057 99.5127
R15922 VDD.n1881 VDD.n1880 99.5127
R15923 VDD.n1877 VDD.n1876 99.5127
R15924 VDD.n1873 VDD.n1872 99.5127
R15925 VDD.n1869 VDD.n1868 99.5127
R15926 VDD.n1865 VDD.n1864 99.5127
R15927 VDD.n1861 VDD.n1860 99.5127
R15928 VDD.n1857 VDD.n1856 99.5127
R15929 VDD.n831 VDD.n765 99.5127
R15930 VDD.n831 VDD.n759 99.5127
R15931 VDD.n834 VDD.n759 99.5127
R15932 VDD.n834 VDD.n753 99.5127
R15933 VDD.n837 VDD.n753 99.5127
R15934 VDD.n837 VDD.n747 99.5127
R15935 VDD.n840 VDD.n747 99.5127
R15936 VDD.n840 VDD.n740 99.5127
R15937 VDD.n843 VDD.n740 99.5127
R15938 VDD.n843 VDD.n734 99.5127
R15939 VDD.n846 VDD.n734 99.5127
R15940 VDD.n846 VDD.n729 99.5127
R15941 VDD.n849 VDD.n729 99.5127
R15942 VDD.n849 VDD.n723 99.5127
R15943 VDD.n852 VDD.n723 99.5127
R15944 VDD.n852 VDD.n717 99.5127
R15945 VDD.n855 VDD.n717 99.5127
R15946 VDD.n855 VDD.n711 99.5127
R15947 VDD.n858 VDD.n711 99.5127
R15948 VDD.n858 VDD.n705 99.5127
R15949 VDD.n861 VDD.n705 99.5127
R15950 VDD.n861 VDD.n699 99.5127
R15951 VDD.n864 VDD.n699 99.5127
R15952 VDD.n864 VDD.n693 99.5127
R15953 VDD.n867 VDD.n693 99.5127
R15954 VDD.n867 VDD.n687 99.5127
R15955 VDD.n870 VDD.n687 99.5127
R15956 VDD.n870 VDD.n680 99.5127
R15957 VDD.n873 VDD.n680 99.5127
R15958 VDD.n873 VDD.n673 99.5127
R15959 VDD.n876 VDD.n673 99.5127
R15960 VDD.n876 VDD.n668 99.5127
R15961 VDD.n879 VDD.n668 99.5127
R15962 VDD.n879 VDD.n663 99.5127
R15963 VDD.n882 VDD.n663 99.5127
R15964 VDD.n882 VDD.n657 99.5127
R15965 VDD.n885 VDD.n657 99.5127
R15966 VDD.n885 VDD.n651 99.5127
R15967 VDD.n888 VDD.n651 99.5127
R15968 VDD.n888 VDD.n645 99.5127
R15969 VDD.n891 VDD.n645 99.5127
R15970 VDD.n891 VDD.n639 99.5127
R15971 VDD.n894 VDD.n639 99.5127
R15972 VDD.n894 VDD.n632 99.5127
R15973 VDD.n897 VDD.n632 99.5127
R15974 VDD.n897 VDD.n626 99.5127
R15975 VDD.n900 VDD.n626 99.5127
R15976 VDD.n900 VDD.n621 99.5127
R15977 VDD.n903 VDD.n621 99.5127
R15978 VDD.n903 VDD.n615 99.5127
R15979 VDD.n906 VDD.n615 99.5127
R15980 VDD.n906 VDD.n609 99.5127
R15981 VDD.n909 VDD.n609 99.5127
R15982 VDD.n909 VDD.n603 99.5127
R15983 VDD.n912 VDD.n603 99.5127
R15984 VDD.n912 VDD.n597 99.5127
R15985 VDD.n915 VDD.n597 99.5127
R15986 VDD.n915 VDD.n591 99.5127
R15987 VDD.n918 VDD.n591 99.5127
R15988 VDD.n918 VDD.n585 99.5127
R15989 VDD.n921 VDD.n585 99.5127
R15990 VDD.n921 VDD.n579 99.5127
R15991 VDD.n924 VDD.n579 99.5127
R15992 VDD.n924 VDD.n573 99.5127
R15993 VDD.n936 VDD.n573 99.5127
R15994 VDD.n936 VDD.n567 99.5127
R15995 VDD.n932 VDD.n567 99.5127
R15996 VDD.n932 VDD.n562 99.5127
R15997 VDD.n929 VDD.n562 99.5127
R15998 VDD.n929 VDD.n555 99.5127
R15999 VDD.n555 VDD.n547 99.5127
R16000 VDD.n1847 VDD.n547 99.5127
R16001 VDD.n1848 VDD.n1847 99.5127
R16002 VDD.n1848 VDD.n538 99.5127
R16003 VDD.n1852 VDD.n538 99.5127
R16004 VDD.n1587 VDD.n1585 99.5127
R16005 VDD.n1585 VDD.n1584 99.5127
R16006 VDD.n1581 VDD.n1580 99.5127
R16007 VDD.n1578 VDD.n771 99.5127
R16008 VDD.n814 VDD.n812 99.5127
R16009 VDD.n818 VDD.n816 99.5127
R16010 VDD.n825 VDD.n809 99.5127
R16011 VDD.n828 VDD.n827 99.5127
R16012 VDD.n1591 VDD.n757 99.5127
R16013 VDD.n1599 VDD.n757 99.5127
R16014 VDD.n1599 VDD.n755 99.5127
R16015 VDD.n1603 VDD.n755 99.5127
R16016 VDD.n1603 VDD.n745 99.5127
R16017 VDD.n1611 VDD.n745 99.5127
R16018 VDD.n1611 VDD.n743 99.5127
R16019 VDD.n1615 VDD.n743 99.5127
R16020 VDD.n1615 VDD.n733 99.5127
R16021 VDD.n1623 VDD.n733 99.5127
R16022 VDD.n1623 VDD.n731 99.5127
R16023 VDD.n1627 VDD.n731 99.5127
R16024 VDD.n1627 VDD.n721 99.5127
R16025 VDD.n1635 VDD.n721 99.5127
R16026 VDD.n1635 VDD.n719 99.5127
R16027 VDD.n1639 VDD.n719 99.5127
R16028 VDD.n1639 VDD.n709 99.5127
R16029 VDD.n1647 VDD.n709 99.5127
R16030 VDD.n1647 VDD.n707 99.5127
R16031 VDD.n1651 VDD.n707 99.5127
R16032 VDD.n1651 VDD.n697 99.5127
R16033 VDD.n1659 VDD.n697 99.5127
R16034 VDD.n1659 VDD.n695 99.5127
R16035 VDD.n1663 VDD.n695 99.5127
R16036 VDD.n1663 VDD.n685 99.5127
R16037 VDD.n1671 VDD.n685 99.5127
R16038 VDD.n1671 VDD.n683 99.5127
R16039 VDD.n1675 VDD.n683 99.5127
R16040 VDD.n1675 VDD.n672 99.5127
R16041 VDD.n1683 VDD.n672 99.5127
R16042 VDD.n1683 VDD.n670 99.5127
R16043 VDD.n1687 VDD.n670 99.5127
R16044 VDD.n1687 VDD.n661 99.5127
R16045 VDD.n1695 VDD.n661 99.5127
R16046 VDD.n1695 VDD.n659 99.5127
R16047 VDD.n1699 VDD.n659 99.5127
R16048 VDD.n1699 VDD.n649 99.5127
R16049 VDD.n1707 VDD.n649 99.5127
R16050 VDD.n1707 VDD.n647 99.5127
R16051 VDD.n1711 VDD.n647 99.5127
R16052 VDD.n1711 VDD.n637 99.5127
R16053 VDD.n1719 VDD.n637 99.5127
R16054 VDD.n1719 VDD.n635 99.5127
R16055 VDD.n1723 VDD.n635 99.5127
R16056 VDD.n1723 VDD.n625 99.5127
R16057 VDD.n1731 VDD.n625 99.5127
R16058 VDD.n1731 VDD.n623 99.5127
R16059 VDD.n1735 VDD.n623 99.5127
R16060 VDD.n1735 VDD.n613 99.5127
R16061 VDD.n1743 VDD.n613 99.5127
R16062 VDD.n1743 VDD.n611 99.5127
R16063 VDD.n1747 VDD.n611 99.5127
R16064 VDD.n1747 VDD.n601 99.5127
R16065 VDD.n1755 VDD.n601 99.5127
R16066 VDD.n1755 VDD.n599 99.5127
R16067 VDD.n1759 VDD.n599 99.5127
R16068 VDD.n1759 VDD.n589 99.5127
R16069 VDD.n1767 VDD.n589 99.5127
R16070 VDD.n1767 VDD.n587 99.5127
R16071 VDD.n1771 VDD.n587 99.5127
R16072 VDD.n1771 VDD.n577 99.5127
R16073 VDD.n1779 VDD.n577 99.5127
R16074 VDD.n1779 VDD.n575 99.5127
R16075 VDD.n1783 VDD.n575 99.5127
R16076 VDD.n1783 VDD.n566 99.5127
R16077 VDD.n1791 VDD.n566 99.5127
R16078 VDD.n1791 VDD.n564 99.5127
R16079 VDD.n1795 VDD.n564 99.5127
R16080 VDD.n1795 VDD.n553 99.5127
R16081 VDD.n1841 VDD.n553 99.5127
R16082 VDD.n1841 VDD.n551 99.5127
R16083 VDD.n1845 VDD.n551 99.5127
R16084 VDD.n1845 VDD.n540 99.5127
R16085 VDD.n1887 VDD.n540 99.5127
R16086 VDD.n1887 VDD.n541 99.5127
R16087 VDD.n2423 VDD.n2409 99.5127
R16088 VDD.n2419 VDD.n2418 99.5127
R16089 VDD.n2416 VDD.n2413 99.5127
R16090 VDD.n2499 VDD.n266 99.5127
R16091 VDD.n2497 VDD.n2496 99.5127
R16092 VDD.n2494 VDD.n269 99.5127
R16093 VDD.n2490 VDD.n2489 99.5127
R16094 VDD.n2048 VDD.n1899 99.5127
R16095 VDD.n1899 VDD.n512 99.5127
R16096 VDD.n2043 VDD.n512 99.5127
R16097 VDD.n2043 VDD.n506 99.5127
R16098 VDD.n2040 VDD.n506 99.5127
R16099 VDD.n2040 VDD.n500 99.5127
R16100 VDD.n2037 VDD.n500 99.5127
R16101 VDD.n2037 VDD.n493 99.5127
R16102 VDD.n2034 VDD.n493 99.5127
R16103 VDD.n2034 VDD.n487 99.5127
R16104 VDD.n2031 VDD.n487 99.5127
R16105 VDD.n2031 VDD.n482 99.5127
R16106 VDD.n2028 VDD.n482 99.5127
R16107 VDD.n2028 VDD.n476 99.5127
R16108 VDD.n2025 VDD.n476 99.5127
R16109 VDD.n2025 VDD.n470 99.5127
R16110 VDD.n2022 VDD.n470 99.5127
R16111 VDD.n2022 VDD.n464 99.5127
R16112 VDD.n2019 VDD.n464 99.5127
R16113 VDD.n2019 VDD.n458 99.5127
R16114 VDD.n2016 VDD.n458 99.5127
R16115 VDD.n2016 VDD.n452 99.5127
R16116 VDD.n2013 VDD.n452 99.5127
R16117 VDD.n2013 VDD.n446 99.5127
R16118 VDD.n2010 VDD.n446 99.5127
R16119 VDD.n2010 VDD.n440 99.5127
R16120 VDD.n2007 VDD.n440 99.5127
R16121 VDD.n2007 VDD.n433 99.5127
R16122 VDD.n2004 VDD.n433 99.5127
R16123 VDD.n2004 VDD.n427 99.5127
R16124 VDD.n2001 VDD.n427 99.5127
R16125 VDD.n2001 VDD.n422 99.5127
R16126 VDD.n1998 VDD.n422 99.5127
R16127 VDD.n1998 VDD.n416 99.5127
R16128 VDD.n1995 VDD.n416 99.5127
R16129 VDD.n1995 VDD.n410 99.5127
R16130 VDD.n1992 VDD.n410 99.5127
R16131 VDD.n1992 VDD.n404 99.5127
R16132 VDD.n1989 VDD.n404 99.5127
R16133 VDD.n1989 VDD.n398 99.5127
R16134 VDD.n1986 VDD.n398 99.5127
R16135 VDD.n1986 VDD.n391 99.5127
R16136 VDD.n1983 VDD.n391 99.5127
R16137 VDD.n1983 VDD.n384 99.5127
R16138 VDD.n1980 VDD.n384 99.5127
R16139 VDD.n1980 VDD.n379 99.5127
R16140 VDD.n1977 VDD.n379 99.5127
R16141 VDD.n1977 VDD.n374 99.5127
R16142 VDD.n1974 VDD.n374 99.5127
R16143 VDD.n1974 VDD.n368 99.5127
R16144 VDD.n1971 VDD.n368 99.5127
R16145 VDD.n1971 VDD.n362 99.5127
R16146 VDD.n1968 VDD.n362 99.5127
R16147 VDD.n1968 VDD.n356 99.5127
R16148 VDD.n1965 VDD.n356 99.5127
R16149 VDD.n1965 VDD.n350 99.5127
R16150 VDD.n1962 VDD.n350 99.5127
R16151 VDD.n1962 VDD.n344 99.5127
R16152 VDD.n1959 VDD.n344 99.5127
R16153 VDD.n1959 VDD.n338 99.5127
R16154 VDD.n1956 VDD.n338 99.5127
R16155 VDD.n1956 VDD.n332 99.5127
R16156 VDD.n1953 VDD.n332 99.5127
R16157 VDD.n1953 VDD.n325 99.5127
R16158 VDD.n1950 VDD.n325 99.5127
R16159 VDD.n1950 VDD.n319 99.5127
R16160 VDD.n1947 VDD.n319 99.5127
R16161 VDD.n1947 VDD.n314 99.5127
R16162 VDD.n1944 VDD.n314 99.5127
R16163 VDD.n1944 VDD.n307 99.5127
R16164 VDD.n1941 VDD.n307 99.5127
R16165 VDD.n1941 VDD.n300 99.5127
R16166 VDD.n300 VDD.n277 99.5127
R16167 VDD.n2483 VDD.n277 99.5127
R16168 VDD.n2483 VDD.n275 99.5127
R16169 VDD.n1913 VDD.n1911 99.5127
R16170 VDD.n1917 VDD.n1908 99.5127
R16171 VDD.n1921 VDD.n1919 99.5127
R16172 VDD.n1925 VDD.n1906 99.5127
R16173 VDD.n1929 VDD.n1927 99.5127
R16174 VDD.n1933 VDD.n1904 99.5127
R16175 VDD.n1937 VDD.n1935 99.5127
R16176 VDD.n2201 VDD.n513 99.5127
R16177 VDD.n2205 VDD.n513 99.5127
R16178 VDD.n2205 VDD.n503 99.5127
R16179 VDD.n2213 VDD.n503 99.5127
R16180 VDD.n2213 VDD.n501 99.5127
R16181 VDD.n2217 VDD.n501 99.5127
R16182 VDD.n2217 VDD.n490 99.5127
R16183 VDD.n2225 VDD.n490 99.5127
R16184 VDD.n2225 VDD.n488 99.5127
R16185 VDD.n2229 VDD.n488 99.5127
R16186 VDD.n2229 VDD.n479 99.5127
R16187 VDD.n2237 VDD.n479 99.5127
R16188 VDD.n2237 VDD.n477 99.5127
R16189 VDD.n2241 VDD.n477 99.5127
R16190 VDD.n2241 VDD.n467 99.5127
R16191 VDD.n2249 VDD.n467 99.5127
R16192 VDD.n2249 VDD.n465 99.5127
R16193 VDD.n2253 VDD.n465 99.5127
R16194 VDD.n2253 VDD.n455 99.5127
R16195 VDD.n2261 VDD.n455 99.5127
R16196 VDD.n2261 VDD.n453 99.5127
R16197 VDD.n2265 VDD.n453 99.5127
R16198 VDD.n2265 VDD.n443 99.5127
R16199 VDD.n2273 VDD.n443 99.5127
R16200 VDD.n2273 VDD.n441 99.5127
R16201 VDD.n2277 VDD.n441 99.5127
R16202 VDD.n2277 VDD.n430 99.5127
R16203 VDD.n2285 VDD.n430 99.5127
R16204 VDD.n2285 VDD.n428 99.5127
R16205 VDD.n2289 VDD.n428 99.5127
R16206 VDD.n2289 VDD.n419 99.5127
R16207 VDD.n2297 VDD.n419 99.5127
R16208 VDD.n2297 VDD.n417 99.5127
R16209 VDD.n2301 VDD.n417 99.5127
R16210 VDD.n2301 VDD.n407 99.5127
R16211 VDD.n2309 VDD.n407 99.5127
R16212 VDD.n2309 VDD.n405 99.5127
R16213 VDD.n2313 VDD.n405 99.5127
R16214 VDD.n2313 VDD.n395 99.5127
R16215 VDD.n2321 VDD.n395 99.5127
R16216 VDD.n2321 VDD.n393 99.5127
R16217 VDD.n2325 VDD.n393 99.5127
R16218 VDD.n2325 VDD.n382 99.5127
R16219 VDD.n2333 VDD.n382 99.5127
R16220 VDD.n2333 VDD.n380 99.5127
R16221 VDD.n2337 VDD.n380 99.5127
R16222 VDD.n2337 VDD.n371 99.5127
R16223 VDD.n2345 VDD.n371 99.5127
R16224 VDD.n2345 VDD.n369 99.5127
R16225 VDD.n2349 VDD.n369 99.5127
R16226 VDD.n2349 VDD.n359 99.5127
R16227 VDD.n2357 VDD.n359 99.5127
R16228 VDD.n2357 VDD.n357 99.5127
R16229 VDD.n2361 VDD.n357 99.5127
R16230 VDD.n2361 VDD.n347 99.5127
R16231 VDD.n2369 VDD.n347 99.5127
R16232 VDD.n2369 VDD.n345 99.5127
R16233 VDD.n2373 VDD.n345 99.5127
R16234 VDD.n2373 VDD.n335 99.5127
R16235 VDD.n2381 VDD.n335 99.5127
R16236 VDD.n2381 VDD.n333 99.5127
R16237 VDD.n2385 VDD.n333 99.5127
R16238 VDD.n2385 VDD.n322 99.5127
R16239 VDD.n2393 VDD.n322 99.5127
R16240 VDD.n2393 VDD.n320 99.5127
R16241 VDD.n2397 VDD.n320 99.5127
R16242 VDD.n2397 VDD.n311 99.5127
R16243 VDD.n2405 VDD.n311 99.5127
R16244 VDD.n2405 VDD.n308 99.5127
R16245 VDD.n2434 VDD.n308 99.5127
R16246 VDD.n2434 VDD.n309 99.5127
R16247 VDD.n309 VDD.n301 99.5127
R16248 VDD.n2429 VDD.n301 99.5127
R16249 VDD.n2429 VDD.n281 99.5127
R16250 VDD.n2426 VDD.n281 99.5127
R16251 VDD.n1827 VDD.n1826 99.5127
R16252 VDD.n1823 VDD.n1822 99.5127
R16253 VDD.n1819 VDD.n1818 99.5127
R16254 VDD.n1815 VDD.n1814 99.5127
R16255 VDD.n1811 VDD.n1810 99.5127
R16256 VDD.n1807 VDD.n1806 99.5127
R16257 VDD.n1803 VDD.n532 99.5127
R16258 VDD.n1034 VDD.n766 99.5127
R16259 VDD.n1034 VDD.n760 99.5127
R16260 VDD.n1031 VDD.n760 99.5127
R16261 VDD.n1031 VDD.n754 99.5127
R16262 VDD.n1028 VDD.n754 99.5127
R16263 VDD.n1028 VDD.n748 99.5127
R16264 VDD.n1025 VDD.n748 99.5127
R16265 VDD.n1025 VDD.n741 99.5127
R16266 VDD.n1022 VDD.n741 99.5127
R16267 VDD.n1022 VDD.n735 99.5127
R16268 VDD.n1019 VDD.n735 99.5127
R16269 VDD.n1019 VDD.n730 99.5127
R16270 VDD.n1016 VDD.n730 99.5127
R16271 VDD.n1016 VDD.n724 99.5127
R16272 VDD.n1013 VDD.n724 99.5127
R16273 VDD.n1013 VDD.n718 99.5127
R16274 VDD.n1010 VDD.n718 99.5127
R16275 VDD.n1010 VDD.n712 99.5127
R16276 VDD.n1007 VDD.n712 99.5127
R16277 VDD.n1007 VDD.n706 99.5127
R16278 VDD.n1004 VDD.n706 99.5127
R16279 VDD.n1004 VDD.n700 99.5127
R16280 VDD.n1001 VDD.n700 99.5127
R16281 VDD.n1001 VDD.n694 99.5127
R16282 VDD.n998 VDD.n694 99.5127
R16283 VDD.n998 VDD.n688 99.5127
R16284 VDD.n995 VDD.n688 99.5127
R16285 VDD.n995 VDD.n681 99.5127
R16286 VDD.n992 VDD.n681 99.5127
R16287 VDD.n992 VDD.n674 99.5127
R16288 VDD.n989 VDD.n674 99.5127
R16289 VDD.n989 VDD.n669 99.5127
R16290 VDD.n986 VDD.n669 99.5127
R16291 VDD.n986 VDD.n664 99.5127
R16292 VDD.n983 VDD.n664 99.5127
R16293 VDD.n983 VDD.n658 99.5127
R16294 VDD.n980 VDD.n658 99.5127
R16295 VDD.n980 VDD.n652 99.5127
R16296 VDD.n977 VDD.n652 99.5127
R16297 VDD.n977 VDD.n646 99.5127
R16298 VDD.n974 VDD.n646 99.5127
R16299 VDD.n974 VDD.n640 99.5127
R16300 VDD.n971 VDD.n640 99.5127
R16301 VDD.n971 VDD.n633 99.5127
R16302 VDD.n968 VDD.n633 99.5127
R16303 VDD.n968 VDD.n627 99.5127
R16304 VDD.n965 VDD.n627 99.5127
R16305 VDD.n965 VDD.n622 99.5127
R16306 VDD.n962 VDD.n622 99.5127
R16307 VDD.n962 VDD.n616 99.5127
R16308 VDD.n959 VDD.n616 99.5127
R16309 VDD.n959 VDD.n610 99.5127
R16310 VDD.n956 VDD.n610 99.5127
R16311 VDD.n956 VDD.n604 99.5127
R16312 VDD.n953 VDD.n604 99.5127
R16313 VDD.n953 VDD.n598 99.5127
R16314 VDD.n950 VDD.n598 99.5127
R16315 VDD.n950 VDD.n592 99.5127
R16316 VDD.n947 VDD.n592 99.5127
R16317 VDD.n947 VDD.n586 99.5127
R16318 VDD.n944 VDD.n586 99.5127
R16319 VDD.n944 VDD.n580 99.5127
R16320 VDD.n941 VDD.n580 99.5127
R16321 VDD.n941 VDD.n574 99.5127
R16322 VDD.n938 VDD.n574 99.5127
R16323 VDD.n938 VDD.n568 99.5127
R16324 VDD.n805 VDD.n568 99.5127
R16325 VDD.n805 VDD.n563 99.5127
R16326 VDD.n802 VDD.n563 99.5127
R16327 VDD.n802 VDD.n556 99.5127
R16328 VDD.n799 VDD.n556 99.5127
R16329 VDD.n799 VDD.n549 99.5127
R16330 VDD.n549 VDD.n536 99.5127
R16331 VDD.n1889 VDD.n536 99.5127
R16332 VDD.n1889 VDD.n533 99.5127
R16333 VDD.n782 VDD.n779 99.5127
R16334 VDD.n786 VDD.n784 99.5127
R16335 VDD.n790 VDD.n776 99.5127
R16336 VDD.n1052 VDD.n792 99.5127
R16337 VDD.n1050 VDD.n1049 99.5127
R16338 VDD.n1046 VDD.n1045 99.5127
R16339 VDD.n1043 VDD.n795 99.5127
R16340 VDD.n1593 VDD.n761 99.5127
R16341 VDD.n1597 VDD.n761 99.5127
R16342 VDD.n1597 VDD.n751 99.5127
R16343 VDD.n1605 VDD.n751 99.5127
R16344 VDD.n1605 VDD.n749 99.5127
R16345 VDD.n1609 VDD.n749 99.5127
R16346 VDD.n1609 VDD.n738 99.5127
R16347 VDD.n1617 VDD.n738 99.5127
R16348 VDD.n1617 VDD.n736 99.5127
R16349 VDD.n1621 VDD.n736 99.5127
R16350 VDD.n1621 VDD.n727 99.5127
R16351 VDD.n1629 VDD.n727 99.5127
R16352 VDD.n1629 VDD.n725 99.5127
R16353 VDD.n1633 VDD.n725 99.5127
R16354 VDD.n1633 VDD.n715 99.5127
R16355 VDD.n1641 VDD.n715 99.5127
R16356 VDD.n1641 VDD.n713 99.5127
R16357 VDD.n1645 VDD.n713 99.5127
R16358 VDD.n1645 VDD.n703 99.5127
R16359 VDD.n1653 VDD.n703 99.5127
R16360 VDD.n1653 VDD.n701 99.5127
R16361 VDD.n1657 VDD.n701 99.5127
R16362 VDD.n1657 VDD.n691 99.5127
R16363 VDD.n1665 VDD.n691 99.5127
R16364 VDD.n1665 VDD.n689 99.5127
R16365 VDD.n1669 VDD.n689 99.5127
R16366 VDD.n1669 VDD.n678 99.5127
R16367 VDD.n1677 VDD.n678 99.5127
R16368 VDD.n1677 VDD.n676 99.5127
R16369 VDD.n1681 VDD.n676 99.5127
R16370 VDD.n1681 VDD.n667 99.5127
R16371 VDD.n1689 VDD.n667 99.5127
R16372 VDD.n1689 VDD.n665 99.5127
R16373 VDD.n1693 VDD.n665 99.5127
R16374 VDD.n1693 VDD.n655 99.5127
R16375 VDD.n1701 VDD.n655 99.5127
R16376 VDD.n1701 VDD.n653 99.5127
R16377 VDD.n1705 VDD.n653 99.5127
R16378 VDD.n1705 VDD.n643 99.5127
R16379 VDD.n1713 VDD.n643 99.5127
R16380 VDD.n1713 VDD.n641 99.5127
R16381 VDD.n1717 VDD.n641 99.5127
R16382 VDD.n1717 VDD.n630 99.5127
R16383 VDD.n1725 VDD.n630 99.5127
R16384 VDD.n1725 VDD.n628 99.5127
R16385 VDD.n1729 VDD.n628 99.5127
R16386 VDD.n1729 VDD.n619 99.5127
R16387 VDD.n1737 VDD.n619 99.5127
R16388 VDD.n1737 VDD.n617 99.5127
R16389 VDD.n1741 VDD.n617 99.5127
R16390 VDD.n1741 VDD.n607 99.5127
R16391 VDD.n1749 VDD.n607 99.5127
R16392 VDD.n1749 VDD.n605 99.5127
R16393 VDD.n1753 VDD.n605 99.5127
R16394 VDD.n1753 VDD.n595 99.5127
R16395 VDD.n1761 VDD.n595 99.5127
R16396 VDD.n1761 VDD.n593 99.5127
R16397 VDD.n1765 VDD.n593 99.5127
R16398 VDD.n1765 VDD.n583 99.5127
R16399 VDD.n1773 VDD.n583 99.5127
R16400 VDD.n1773 VDD.n581 99.5127
R16401 VDD.n1777 VDD.n581 99.5127
R16402 VDD.n1777 VDD.n571 99.5127
R16403 VDD.n1785 VDD.n571 99.5127
R16404 VDD.n1785 VDD.n569 99.5127
R16405 VDD.n1789 VDD.n569 99.5127
R16406 VDD.n1789 VDD.n560 99.5127
R16407 VDD.n1797 VDD.n560 99.5127
R16408 VDD.n1797 VDD.n557 99.5127
R16409 VDD.n1839 VDD.n557 99.5127
R16410 VDD.n1839 VDD.n558 99.5127
R16411 VDD.n558 VDD.n550 99.5127
R16412 VDD.n1834 VDD.n550 99.5127
R16413 VDD.n1834 VDD.n539 99.5127
R16414 VDD.n1831 VDD.n539 99.5127
R16415 VDD.n778 VDD.n764 72.8958
R16416 VDD.n783 VDD.n764 72.8958
R16417 VDD.n785 VDD.n764 72.8958
R16418 VDD.n791 VDD.n764 72.8958
R16419 VDD.n1051 VDD.n764 72.8958
R16420 VDD.n793 VDD.n764 72.8958
R16421 VDD.n1044 VDD.n764 72.8958
R16422 VDD.n1037 VDD.n764 72.8958
R16423 VDD.n1895 VDD.n1894 72.8958
R16424 VDD.n1895 VDD.n531 72.8958
R16425 VDD.n1895 VDD.n530 72.8958
R16426 VDD.n1895 VDD.n529 72.8958
R16427 VDD.n1895 VDD.n528 72.8958
R16428 VDD.n1895 VDD.n527 72.8958
R16429 VDD.n1895 VDD.n526 72.8958
R16430 VDD.n1895 VDD.n525 72.8958
R16431 VDD.n1910 VDD.n1896 72.8958
R16432 VDD.n1912 VDD.n1896 72.8958
R16433 VDD.n1918 VDD.n1896 72.8958
R16434 VDD.n1920 VDD.n1896 72.8958
R16435 VDD.n1926 VDD.n1896 72.8958
R16436 VDD.n1928 VDD.n1896 72.8958
R16437 VDD.n1934 VDD.n1896 72.8958
R16438 VDD.n1936 VDD.n1896 72.8958
R16439 VDD.n2488 VDD.n267 72.8958
R16440 VDD.n273 VDD.n267 72.8958
R16441 VDD.n2495 VDD.n267 72.8958
R16442 VDD.n2498 VDD.n267 72.8958
R16443 VDD.n2412 VDD.n267 72.8958
R16444 VDD.n2417 VDD.n267 72.8958
R16445 VDD.n2411 VDD.n267 72.8958
R16446 VDD.n2424 VDD.n267 72.8958
R16447 VDD.n1586 VDD.n764 72.8958
R16448 VDD.n769 VDD.n764 72.8958
R16449 VDD.n1579 VDD.n764 72.8958
R16450 VDD.n811 VDD.n764 72.8958
R16451 VDD.n815 VDD.n764 72.8958
R16452 VDD.n817 VDD.n764 72.8958
R16453 VDD.n826 VDD.n764 72.8958
R16454 VDD.n1895 VDD.n524 72.8958
R16455 VDD.n1895 VDD.n523 72.8958
R16456 VDD.n1895 VDD.n522 72.8958
R16457 VDD.n1895 VDD.n521 72.8958
R16458 VDD.n1895 VDD.n520 72.8958
R16459 VDD.n1895 VDD.n519 72.8958
R16460 VDD.n1895 VDD.n518 72.8958
R16461 VDD.n1895 VDD.n517 72.8958
R16462 VDD.n2194 VDD.n1896 72.8958
R16463 VDD.n2051 VDD.n1896 72.8958
R16464 VDD.n2187 VDD.n1896 72.8958
R16465 VDD.n2181 VDD.n1896 72.8958
R16466 VDD.n2179 VDD.n1896 72.8958
R16467 VDD.n2173 VDD.n1896 72.8958
R16468 VDD.n2171 VDD.n1896 72.8958
R16469 VDD.n2447 VDD.n267 72.8958
R16470 VDD.n2455 VDD.n267 72.8958
R16471 VDD.n293 VDD.n267 72.8958
R16472 VDD.n2462 VDD.n267 72.8958
R16473 VDD.n2466 VDD.n267 72.8958
R16474 VDD.n289 VDD.n267 72.8958
R16475 VDD.n2473 VDD.n267 72.8958
R16476 VDD.n2476 VDD.n267 72.8958
R16477 VDD.n2548 VDD.n219 66.2847
R16478 VDD.n225 VDD.n219 66.2847
R16479 VDD.n2541 VDD.n219 66.2847
R16480 VDD.n2535 VDD.n219 66.2847
R16481 VDD.n2533 VDD.n219 66.2847
R16482 VDD.n2527 VDD.n219 66.2847
R16483 VDD.n2525 VDD.n219 66.2847
R16484 VDD.n2519 VDD.n219 66.2847
R16485 VDD.n2517 VDD.n219 66.2847
R16486 VDD.n2511 VDD.n219 66.2847
R16487 VDD.n2509 VDD.n219 66.2847
R16488 VDD.n257 VDD.n219 66.2847
R16489 VDD.n2682 VDD.n91 66.2847
R16490 VDD.n135 VDD.n91 66.2847
R16491 VDD.n2689 VDD.n91 66.2847
R16492 VDD.n2692 VDD.n91 66.2847
R16493 VDD.n126 VDD.n91 66.2847
R16494 VDD.n2701 VDD.n91 66.2847
R16495 VDD.n117 VDD.n91 66.2847
R16496 VDD.n2708 VDD.n91 66.2847
R16497 VDD.n111 VDD.n91 66.2847
R16498 VDD.n106 VDD.n91 66.2847
R16499 VDD.n2719 VDD.n91 66.2847
R16500 VDD.n98 VDD.n91 66.2847
R16501 VDD.n1552 VDD.n1551 66.2847
R16502 VDD.n1552 VDD.n1550 66.2847
R16503 VDD.n1552 VDD.n1549 66.2847
R16504 VDD.n1552 VDD.n1547 66.2847
R16505 VDD.n1552 VDD.n1546 66.2847
R16506 VDD.n1552 VDD.n1544 66.2847
R16507 VDD.n1552 VDD.n1543 66.2847
R16508 VDD.n1552 VDD.n1086 66.2847
R16509 VDD.n1552 VDD.n1085 66.2847
R16510 VDD.n1552 VDD.n1084 66.2847
R16511 VDD.n1552 VDD.n1083 66.2847
R16512 VDD.n1552 VDD.n1082 66.2847
R16513 VDD.n1230 VDD.n1227 66.2847
R16514 VDD.n1236 VDD.n1227 66.2847
R16515 VDD.n1306 VDD.n1227 66.2847
R16516 VDD.n1304 VDD.n1227 66.2847
R16517 VDD.n1245 VDD.n1227 66.2847
R16518 VDD.n1248 VDD.n1227 66.2847
R16519 VDD.n1253 VDD.n1227 66.2847
R16520 VDD.n1287 VDD.n1227 66.2847
R16521 VDD.n1256 VDD.n1227 66.2847
R16522 VDD.n1262 VDD.n1227 66.2847
R16523 VDD.n1266 VDD.n1227 66.2847
R16524 VDD.n1268 VDD.n1227 66.2847
R16525 VDD.n1272 VDD.n1271 63.2247
R16526 VDD.n1290 VDD.n1289 63.2247
R16527 VDD.n1309 VDD.n1308 63.2247
R16528 VDD.n234 VDD.n233 63.2247
R16529 VDD.n248 VDD.n247 63.2247
R16530 VDD.n262 VDD.n261 63.2247
R16531 VDD.n137 VDD.n136 63.2247
R16532 VDD.n123 VDD.n122 63.2247
R16533 VDD.n105 VDD.n104 63.2247
R16534 VDD.n1092 VDD.n1091 63.2247
R16535 VDD.n1063 VDD.n1062 63.2247
R16536 VDD.n1077 VDD.n1076 63.2247
R16537 VDD.n2721 VDD.n98 52.4337
R16538 VDD.n2719 VDD.n2718 52.4337
R16539 VDD.n107 VDD.n106 52.4337
R16540 VDD.n2710 VDD.n111 52.4337
R16541 VDD.n2708 VDD.n2707 52.4337
R16542 VDD.n2703 VDD.n117 52.4337
R16543 VDD.n2701 VDD.n2700 52.4337
R16544 VDD.n127 VDD.n126 52.4337
R16545 VDD.n2692 VDD.n2691 52.4337
R16546 VDD.n2689 VDD.n2688 52.4337
R16547 VDD.n2684 VDD.n135 52.4337
R16548 VDD.n2682 VDD.n2681 52.4337
R16549 VDD.n2548 VDD.n220 52.4337
R16550 VDD.n2546 VDD.n225 52.4337
R16551 VDD.n2542 VDD.n2541 52.4337
R16552 VDD.n2535 VDD.n230 52.4337
R16553 VDD.n2534 VDD.n2533 52.4337
R16554 VDD.n2527 VDD.n238 52.4337
R16555 VDD.n2526 VDD.n2525 52.4337
R16556 VDD.n2519 VDD.n243 52.4337
R16557 VDD.n2518 VDD.n2517 52.4337
R16558 VDD.n2511 VDD.n251 52.4337
R16559 VDD.n2510 VDD.n2509 52.4337
R16560 VDD.n258 VDD.n257 52.4337
R16561 VDD.n2549 VDD.n2548 52.4337
R16562 VDD.n2543 VDD.n225 52.4337
R16563 VDD.n2541 VDD.n2540 52.4337
R16564 VDD.n2536 VDD.n2535 52.4337
R16565 VDD.n2533 VDD.n2532 52.4337
R16566 VDD.n2528 VDD.n2527 52.4337
R16567 VDD.n2525 VDD.n2524 52.4337
R16568 VDD.n2520 VDD.n2519 52.4337
R16569 VDD.n2517 VDD.n2516 52.4337
R16570 VDD.n2512 VDD.n2511 52.4337
R16571 VDD.n2509 VDD.n2508 52.4337
R16572 VDD.n257 VDD.n218 52.4337
R16573 VDD.n2683 VDD.n2682 52.4337
R16574 VDD.n135 VDD.n129 52.4337
R16575 VDD.n2690 VDD.n2689 52.4337
R16576 VDD.n2693 VDD.n2692 52.4337
R16577 VDD.n126 VDD.n118 52.4337
R16578 VDD.n2702 VDD.n2701 52.4337
R16579 VDD.n117 VDD.n112 52.4337
R16580 VDD.n2709 VDD.n2708 52.4337
R16581 VDD.n111 VDD.n110 52.4337
R16582 VDD.n106 VDD.n99 52.4337
R16583 VDD.n2720 VDD.n2719 52.4337
R16584 VDD.n98 VDD.n95 52.4337
R16585 VDD.n1517 VDD.n1082 52.4337
R16586 VDD.n1096 VDD.n1083 52.4337
R16587 VDD.n1525 VDD.n1084 52.4337
R16588 VDD.n1531 VDD.n1085 52.4337
R16589 VDD.n1535 VDD.n1086 52.4337
R16590 VDD.n1543 VDD.n1541 52.4337
R16591 VDD.n1544 VDD.n1059 52.4337
R16592 VDD.n1546 VDD.n1061 52.4337
R16593 VDD.n1547 VDD.n1066 52.4337
R16594 VDD.n1549 VDD.n1068 52.4337
R16595 VDD.n1550 VDD.n1071 52.4337
R16596 VDD.n1551 VDD.n1073 52.4337
R16597 VDD.n1551 VDD.n1079 52.4337
R16598 VDD.n1550 VDD.n1072 52.4337
R16599 VDD.n1549 VDD.n1548 52.4337
R16600 VDD.n1547 VDD.n1067 52.4337
R16601 VDD.n1546 VDD.n1545 52.4337
R16602 VDD.n1544 VDD.n1060 52.4337
R16603 VDD.n1543 VDD.n1542 52.4337
R16604 VDD.n1087 VDD.n1086 52.4337
R16605 VDD.n1534 VDD.n1085 52.4337
R16606 VDD.n1530 VDD.n1084 52.4337
R16607 VDD.n1524 VDD.n1083 52.4337
R16608 VDD.n1095 VDD.n1082 52.4337
R16609 VDD.n1230 VDD.n1228 52.4337
R16610 VDD.n1236 VDD.n1235 52.4337
R16611 VDD.n1306 VDD.n1238 52.4337
R16612 VDD.n1305 VDD.n1304 52.4337
R16613 VDD.n1245 VDD.n1241 52.4337
R16614 VDD.n1248 VDD.n1247 52.4337
R16615 VDD.n1253 VDD.n1252 52.4337
R16616 VDD.n1288 VDD.n1287 52.4337
R16617 VDD.n1285 VDD.n1256 52.4337
R16618 VDD.n1262 VDD.n1261 52.4337
R16619 VDD.n1266 VDD.n1264 52.4337
R16620 VDD.n1269 VDD.n1268 52.4337
R16621 VDD.n1231 VDD.n1230 52.4337
R16622 VDD.n1237 VDD.n1236 52.4337
R16623 VDD.n1307 VDD.n1306 52.4337
R16624 VDD.n1304 VDD.n1303 52.4337
R16625 VDD.n1246 VDD.n1245 52.4337
R16626 VDD.n1249 VDD.n1248 52.4337
R16627 VDD.n1254 VDD.n1253 52.4337
R16628 VDD.n1287 VDD.n1286 52.4337
R16629 VDD.n1260 VDD.n1256 52.4337
R16630 VDD.n1263 VDD.n1262 52.4337
R16631 VDD.n1267 VDD.n1266 52.4337
R16632 VDD.n1268 VDD.n1226 52.4337
R16633 VDD.n2476 VDD.n2475 39.2114
R16634 VDD.n2473 VDD.n2472 39.2114
R16635 VDD.n2468 VDD.n289 39.2114
R16636 VDD.n2466 VDD.n2465 39.2114
R16637 VDD.n2462 VDD.n2461 39.2114
R16638 VDD.n2457 VDD.n293 39.2114
R16639 VDD.n2455 VDD.n2454 39.2114
R16640 VDD.n2449 VDD.n2447 39.2114
R16641 VDD.n2194 VDD.n2049 39.2114
R16642 VDD.n2192 VDD.n2051 39.2114
R16643 VDD.n2188 VDD.n2187 39.2114
R16644 VDD.n2181 VDD.n2053 39.2114
R16645 VDD.n2180 VDD.n2179 39.2114
R16646 VDD.n2173 VDD.n2055 39.2114
R16647 VDD.n2172 VDD.n2171 39.2114
R16648 VDD.n1881 VDD.n517 39.2114
R16649 VDD.n1877 VDD.n518 39.2114
R16650 VDD.n1873 VDD.n519 39.2114
R16651 VDD.n1869 VDD.n520 39.2114
R16652 VDD.n1865 VDD.n521 39.2114
R16653 VDD.n1861 VDD.n522 39.2114
R16654 VDD.n1857 VDD.n523 39.2114
R16655 VDD.n1853 VDD.n524 39.2114
R16656 VDD.n1586 VDD.n767 39.2114
R16657 VDD.n1584 VDD.n769 39.2114
R16658 VDD.n1580 VDD.n1579 39.2114
R16659 VDD.n811 VDD.n771 39.2114
R16660 VDD.n815 VDD.n814 39.2114
R16661 VDD.n818 VDD.n817 39.2114
R16662 VDD.n826 VDD.n825 39.2114
R16663 VDD.n2424 VDD.n2423 39.2114
R16664 VDD.n2419 VDD.n2411 39.2114
R16665 VDD.n2417 VDD.n2416 39.2114
R16666 VDD.n2412 VDD.n266 39.2114
R16667 VDD.n2498 VDD.n2497 39.2114
R16668 VDD.n2495 VDD.n2494 39.2114
R16669 VDD.n2490 VDD.n273 39.2114
R16670 VDD.n2488 VDD.n2487 39.2114
R16671 VDD.n1910 VDD.n515 39.2114
R16672 VDD.n1913 VDD.n1912 39.2114
R16673 VDD.n1918 VDD.n1917 39.2114
R16674 VDD.n1921 VDD.n1920 39.2114
R16675 VDD.n1926 VDD.n1925 39.2114
R16676 VDD.n1929 VDD.n1928 39.2114
R16677 VDD.n1934 VDD.n1933 39.2114
R16678 VDD.n1937 VDD.n1936 39.2114
R16679 VDD.n1827 VDD.n525 39.2114
R16680 VDD.n1823 VDD.n526 39.2114
R16681 VDD.n1819 VDD.n527 39.2114
R16682 VDD.n1815 VDD.n528 39.2114
R16683 VDD.n1811 VDD.n529 39.2114
R16684 VDD.n1807 VDD.n530 39.2114
R16685 VDD.n1803 VDD.n531 39.2114
R16686 VDD.n1894 VDD.n1893 39.2114
R16687 VDD.n778 VDD.n763 39.2114
R16688 VDD.n783 VDD.n782 39.2114
R16689 VDD.n786 VDD.n785 39.2114
R16690 VDD.n791 VDD.n790 39.2114
R16691 VDD.n1052 VDD.n1051 39.2114
R16692 VDD.n1049 VDD.n793 39.2114
R16693 VDD.n1045 VDD.n1044 39.2114
R16694 VDD.n1037 VDD.n795 39.2114
R16695 VDD.n779 VDD.n778 39.2114
R16696 VDD.n784 VDD.n783 39.2114
R16697 VDD.n785 VDD.n776 39.2114
R16698 VDD.n792 VDD.n791 39.2114
R16699 VDD.n1051 VDD.n1050 39.2114
R16700 VDD.n1046 VDD.n793 39.2114
R16701 VDD.n1044 VDD.n1043 39.2114
R16702 VDD.n1038 VDD.n1037 39.2114
R16703 VDD.n1894 VDD.n532 39.2114
R16704 VDD.n1806 VDD.n531 39.2114
R16705 VDD.n1810 VDD.n530 39.2114
R16706 VDD.n1814 VDD.n529 39.2114
R16707 VDD.n1818 VDD.n528 39.2114
R16708 VDD.n1822 VDD.n527 39.2114
R16709 VDD.n1826 VDD.n526 39.2114
R16710 VDD.n1830 VDD.n525 39.2114
R16711 VDD.n1911 VDD.n1910 39.2114
R16712 VDD.n1912 VDD.n1908 39.2114
R16713 VDD.n1919 VDD.n1918 39.2114
R16714 VDD.n1920 VDD.n1906 39.2114
R16715 VDD.n1927 VDD.n1926 39.2114
R16716 VDD.n1928 VDD.n1904 39.2114
R16717 VDD.n1935 VDD.n1934 39.2114
R16718 VDD.n1936 VDD.n1898 39.2114
R16719 VDD.n2489 VDD.n2488 39.2114
R16720 VDD.n273 VDD.n269 39.2114
R16721 VDD.n2496 VDD.n2495 39.2114
R16722 VDD.n2499 VDD.n2498 39.2114
R16723 VDD.n2413 VDD.n2412 39.2114
R16724 VDD.n2418 VDD.n2417 39.2114
R16725 VDD.n2411 VDD.n2409 39.2114
R16726 VDD.n2425 VDD.n2424 39.2114
R16727 VDD.n1587 VDD.n1586 39.2114
R16728 VDD.n1581 VDD.n769 39.2114
R16729 VDD.n1579 VDD.n1578 39.2114
R16730 VDD.n812 VDD.n811 39.2114
R16731 VDD.n816 VDD.n815 39.2114
R16732 VDD.n817 VDD.n809 39.2114
R16733 VDD.n827 VDD.n826 39.2114
R16734 VDD.n1856 VDD.n524 39.2114
R16735 VDD.n1860 VDD.n523 39.2114
R16736 VDD.n1864 VDD.n522 39.2114
R16737 VDD.n1868 VDD.n521 39.2114
R16738 VDD.n1872 VDD.n520 39.2114
R16739 VDD.n1876 VDD.n519 39.2114
R16740 VDD.n1880 VDD.n518 39.2114
R16741 VDD.n1883 VDD.n517 39.2114
R16742 VDD.n2195 VDD.n2194 39.2114
R16743 VDD.n2189 VDD.n2051 39.2114
R16744 VDD.n2187 VDD.n2186 39.2114
R16745 VDD.n2182 VDD.n2181 39.2114
R16746 VDD.n2179 VDD.n2178 39.2114
R16747 VDD.n2174 VDD.n2173 39.2114
R16748 VDD.n2171 VDD.n2170 39.2114
R16749 VDD.n2447 VDD.n294 39.2114
R16750 VDD.n2456 VDD.n2455 39.2114
R16751 VDD.n293 VDD.n291 39.2114
R16752 VDD.n2463 VDD.n2462 39.2114
R16753 VDD.n2467 VDD.n2466 39.2114
R16754 VDD.n289 VDD.n287 39.2114
R16755 VDD.n2474 VDD.n2473 39.2114
R16756 VDD.n2477 VDD.n2476 39.2114
R16757 VDD.n2168 VDD.n2167 37.4639
R16758 VDD.n2450 VDD.n2446 37.4639
R16759 VDD.n2198 VDD.n2197 37.4639
R16760 VDD.n2479 VDD.n2478 37.4639
R16761 VDD.n2427 VDD.n2408 37.4639
R16762 VDD.n2486 VDD.n2485 37.4639
R16763 VDD.n2047 VDD.n1939 37.4639
R16764 VDD.n2202 VDD.n514 37.4639
R16765 VDD.n1590 VDD.n1589 37.4639
R16766 VDD.n1885 VDD.n1884 37.4639
R16767 VDD.n1854 VDD.n1851 37.4639
R16768 VDD.n830 VDD.n829 37.4639
R16769 VDD.n1832 VDD.n1829 37.4639
R16770 VDD.n1892 VDD.n1891 37.4639
R16771 VDD.n1039 VDD.n1036 37.4639
R16772 VDD.n1594 VDD.n762 37.4639
R16773 VDD.n1273 VDD.n1272 37.2369
R16774 VDD.n1291 VDD.n1290 37.2369
R16775 VDD.n1310 VDD.n1309 37.2369
R16776 VDD.n2539 VDD.n234 37.2369
R16777 VDD.n2522 VDD.n248 37.2369
R16778 VDD.n263 VDD.n262 37.2369
R16779 VDD.n138 VDD.n137 37.2369
R16780 VDD.n2698 VDD.n123 37.2369
R16781 VDD.n2715 VDD.n105 37.2369
R16782 VDD.n1532 VDD.n1092 37.2369
R16783 VDD.n1064 VDD.n1063 37.2369
R16784 VDD.n1078 VDD.n1077 37.2369
R16785 VDD.n1323 VDD.n1227 35.7764
R16786 VDD.n1552 VDD.n1081 35.7764
R16787 VDD.n2558 VDD.n219 35.7764
R16788 VDD.n2729 VDD.n91 35.7764
R16789 VDD.n1592 VDD.n764 30.6039
R16790 VDD.n1895 VDD.n516 30.6039
R16791 VDD.n2200 VDD.n1896 30.6039
R16792 VDD.n280 VDD.n267 30.6039
R16793 VDD.n1902 VDD.n1901 30.449
R16794 VDD.n2452 VDD.n296 30.449
R16795 VDD.n2060 VDD.n2059 30.449
R16796 VDD.n272 VDD.n271 30.449
R16797 VDD.n1041 VDD.n797 30.449
R16798 VDD.n823 VDD.n822 30.449
R16799 VDD.n545 VDD.n544 30.449
R16800 VDD.n1802 VDD.n1801 30.449
R16801 VDD.n1323 VDD.n1222 21.5522
R16802 VDD.n1332 VDD.n1222 21.5522
R16803 VDD.n1332 VDD.n1331 21.5522
R16804 VDD.n1340 VDD.n1211 21.5522
R16805 VDD.n1348 VDD.n1211 21.5522
R16806 VDD.n1348 VDD.n1205 21.5522
R16807 VDD.n1356 VDD.n1205 21.5522
R16808 VDD.n1356 VDD.n1199 21.5522
R16809 VDD.n1364 VDD.n1199 21.5522
R16810 VDD.n1364 VDD.n1193 21.5522
R16811 VDD.n1372 VDD.n1193 21.5522
R16812 VDD.n1380 VDD.n1187 21.5522
R16813 VDD.n1380 VDD.n1181 21.5522
R16814 VDD.n1388 VDD.n1181 21.5522
R16815 VDD.n1388 VDD.n1175 21.5522
R16816 VDD.n1396 VDD.n1175 21.5522
R16817 VDD.n1404 VDD.n1169 21.5522
R16818 VDD.n1404 VDD.n1163 21.5522
R16819 VDD.n1412 VDD.n1163 21.5522
R16820 VDD.n1412 VDD.n1156 21.5522
R16821 VDD.n1432 VDD.n1156 21.5522
R16822 VDD.n1432 VDD.n1157 21.5522
R16823 VDD.n1440 VDD.n1145 21.5522
R16824 VDD.n1448 VDD.n1145 21.5522
R16825 VDD.n1448 VDD.n1139 21.5522
R16826 VDD.n1457 VDD.n1139 21.5522
R16827 VDD.n1457 VDD.n1456 21.5522
R16828 VDD.n1465 VDD.n1128 21.5522
R16829 VDD.n1473 VDD.n1128 21.5522
R16830 VDD.n1473 VDD.n1122 21.5522
R16831 VDD.n1481 VDD.n1122 21.5522
R16832 VDD.n1481 VDD.n1115 21.5522
R16833 VDD.n1490 VDD.n1115 21.5522
R16834 VDD.n1490 VDD.n1109 21.5522
R16835 VDD.n1498 VDD.n1109 21.5522
R16836 VDD.n1509 VDD.n1102 21.5522
R16837 VDD.n1509 VDD.n1508 21.5522
R16838 VDD.n1508 VDD.n1081 21.5522
R16839 VDD.n2558 VDD.n214 21.5522
R16840 VDD.n2567 VDD.n214 21.5522
R16841 VDD.n2567 VDD.n2566 21.5522
R16842 VDD.n2575 VDD.n203 21.5522
R16843 VDD.n2583 VDD.n203 21.5522
R16844 VDD.n2583 VDD.n197 21.5522
R16845 VDD.n2591 VDD.n197 21.5522
R16846 VDD.n2591 VDD.n191 21.5522
R16847 VDD.n2599 VDD.n191 21.5522
R16848 VDD.n2599 VDD.n185 21.5522
R16849 VDD.n2607 VDD.n185 21.5522
R16850 VDD.n2615 VDD.n179 21.5522
R16851 VDD.n2615 VDD.n173 21.5522
R16852 VDD.n2623 VDD.n173 21.5522
R16853 VDD.n2623 VDD.n167 21.5522
R16854 VDD.n2631 VDD.n167 21.5522
R16855 VDD.n2639 VDD.n161 21.5522
R16856 VDD.n2639 VDD.n33 21.5522
R16857 VDD.n2771 VDD.n33 21.5522
R16858 VDD.n2771 VDD.n2770 21.5522
R16859 VDD.n2770 VDD.n2769 21.5522
R16860 VDD.n2769 VDD.n37 21.5522
R16861 VDD.n2763 VDD.n2762 21.5522
R16862 VDD.n2762 VDD.n2761 21.5522
R16863 VDD.n2761 VDD.n47 21.5522
R16864 VDD.n2755 VDD.n47 21.5522
R16865 VDD.n2755 VDD.n2754 21.5522
R16866 VDD.n2753 VDD.n58 21.5522
R16867 VDD.n2747 VDD.n58 21.5522
R16868 VDD.n2747 VDD.n2746 21.5522
R16869 VDD.n2746 VDD.n2745 21.5522
R16870 VDD.n2745 VDD.n69 21.5522
R16871 VDD.n2739 VDD.n69 21.5522
R16872 VDD.n2739 VDD.n2738 21.5522
R16873 VDD.n2738 VDD.n2737 21.5522
R16874 VDD.n2731 VDD.n87 21.5522
R16875 VDD.n2731 VDD.n2730 21.5522
R16876 VDD.n2730 VDD.n2729 21.5522
R16877 VDD.n1284 VDD.n1255 19.3944
R16878 VDD.n1284 VDD.n1257 19.3944
R16879 VDD.n1280 VDD.n1257 19.3944
R16880 VDD.n1280 VDD.n1279 19.3944
R16881 VDD.n1279 VDD.n1278 19.3944
R16882 VDD.n1278 VDD.n1265 19.3944
R16883 VDD.n1274 VDD.n1265 19.3944
R16884 VDD.n1302 VDD.n1239 19.3944
R16885 VDD.n1302 VDD.n1242 19.3944
R16886 VDD.n1298 VDD.n1242 19.3944
R16887 VDD.n1298 VDD.n1297 19.3944
R16888 VDD.n1297 VDD.n1296 19.3944
R16889 VDD.n1296 VDD.n1250 19.3944
R16890 VDD.n1292 VDD.n1250 19.3944
R16891 VDD.n1318 VDD.n1317 19.3944
R16892 VDD.n1317 VDD.n1316 19.3944
R16893 VDD.n1316 VDD.n1233 19.3944
R16894 VDD.n1312 VDD.n1233 19.3944
R16895 VDD.n1312 VDD.n1311 19.3944
R16896 VDD.n1325 VDD.n1224 19.3944
R16897 VDD.n1329 VDD.n1224 19.3944
R16898 VDD.n1329 VDD.n1215 19.3944
R16899 VDD.n1342 VDD.n1215 19.3944
R16900 VDD.n1342 VDD.n1213 19.3944
R16901 VDD.n1346 VDD.n1213 19.3944
R16902 VDD.n1346 VDD.n1203 19.3944
R16903 VDD.n1358 VDD.n1203 19.3944
R16904 VDD.n1358 VDD.n1201 19.3944
R16905 VDD.n1362 VDD.n1201 19.3944
R16906 VDD.n1362 VDD.n1191 19.3944
R16907 VDD.n1374 VDD.n1191 19.3944
R16908 VDD.n1374 VDD.n1189 19.3944
R16909 VDD.n1378 VDD.n1189 19.3944
R16910 VDD.n1378 VDD.n1179 19.3944
R16911 VDD.n1390 VDD.n1179 19.3944
R16912 VDD.n1390 VDD.n1177 19.3944
R16913 VDD.n1394 VDD.n1177 19.3944
R16914 VDD.n1394 VDD.n1167 19.3944
R16915 VDD.n1406 VDD.n1167 19.3944
R16916 VDD.n1406 VDD.n1165 19.3944
R16917 VDD.n1410 VDD.n1165 19.3944
R16918 VDD.n1410 VDD.n1154 19.3944
R16919 VDD.n1434 VDD.n1154 19.3944
R16920 VDD.n1434 VDD.n1152 19.3944
R16921 VDD.n1438 VDD.n1152 19.3944
R16922 VDD.n1438 VDD.n1143 19.3944
R16923 VDD.n1450 VDD.n1143 19.3944
R16924 VDD.n1450 VDD.n1141 19.3944
R16925 VDD.n1454 VDD.n1141 19.3944
R16926 VDD.n1454 VDD.n1132 19.3944
R16927 VDD.n1467 VDD.n1132 19.3944
R16928 VDD.n1467 VDD.n1130 19.3944
R16929 VDD.n1471 VDD.n1130 19.3944
R16930 VDD.n1471 VDD.n1120 19.3944
R16931 VDD.n1483 VDD.n1120 19.3944
R16932 VDD.n1483 VDD.n1117 19.3944
R16933 VDD.n1488 VDD.n1117 19.3944
R16934 VDD.n1488 VDD.n1118 19.3944
R16935 VDD.n1118 VDD.n1107 19.3944
R16936 VDD.n1501 VDD.n1107 19.3944
R16937 VDD.n1501 VDD.n1104 19.3944
R16938 VDD.n1506 VDD.n1104 19.3944
R16939 VDD.n1506 VDD.n1105 19.3944
R16940 VDD.n2551 VDD.n2550 19.3944
R16941 VDD.n2550 VDD.n224 19.3944
R16942 VDD.n2545 VDD.n224 19.3944
R16943 VDD.n2545 VDD.n2544 19.3944
R16944 VDD.n2544 VDD.n229 19.3944
R16945 VDD.n2538 VDD.n2537 19.3944
R16946 VDD.n2537 VDD.n237 19.3944
R16947 VDD.n2531 VDD.n237 19.3944
R16948 VDD.n2531 VDD.n2530 19.3944
R16949 VDD.n2530 VDD.n2529 19.3944
R16950 VDD.n2529 VDD.n242 19.3944
R16951 VDD.n2523 VDD.n242 19.3944
R16952 VDD.n2521 VDD.n250 19.3944
R16953 VDD.n2515 VDD.n250 19.3944
R16954 VDD.n2515 VDD.n2514 19.3944
R16955 VDD.n2514 VDD.n2513 19.3944
R16956 VDD.n2513 VDD.n256 19.3944
R16957 VDD.n2507 VDD.n256 19.3944
R16958 VDD.n2507 VDD.n2506 19.3944
R16959 VDD.n2556 VDD.n212 19.3944
R16960 VDD.n2569 VDD.n212 19.3944
R16961 VDD.n2569 VDD.n210 19.3944
R16962 VDD.n2573 VDD.n210 19.3944
R16963 VDD.n2573 VDD.n201 19.3944
R16964 VDD.n2585 VDD.n201 19.3944
R16965 VDD.n2585 VDD.n199 19.3944
R16966 VDD.n2589 VDD.n199 19.3944
R16967 VDD.n2589 VDD.n189 19.3944
R16968 VDD.n2601 VDD.n189 19.3944
R16969 VDD.n2601 VDD.n187 19.3944
R16970 VDD.n2605 VDD.n187 19.3944
R16971 VDD.n2605 VDD.n177 19.3944
R16972 VDD.n2617 VDD.n177 19.3944
R16973 VDD.n2617 VDD.n175 19.3944
R16974 VDD.n2621 VDD.n175 19.3944
R16975 VDD.n2621 VDD.n165 19.3944
R16976 VDD.n2633 VDD.n165 19.3944
R16977 VDD.n2633 VDD.n163 19.3944
R16978 VDD.n2637 VDD.n163 19.3944
R16979 VDD.n2637 VDD.n29 19.3944
R16980 VDD.n2773 VDD.n29 19.3944
R16981 VDD.n2773 VDD.n30 19.3944
R16982 VDD.n2767 VDD.n30 19.3944
R16983 VDD.n2767 VDD.n2766 19.3944
R16984 VDD.n2766 VDD.n2765 19.3944
R16985 VDD.n2765 VDD.n42 19.3944
R16986 VDD.n2759 VDD.n42 19.3944
R16987 VDD.n2759 VDD.n2758 19.3944
R16988 VDD.n2758 VDD.n2757 19.3944
R16989 VDD.n2757 VDD.n53 19.3944
R16990 VDD.n2751 VDD.n53 19.3944
R16991 VDD.n2751 VDD.n2750 19.3944
R16992 VDD.n2750 VDD.n2749 19.3944
R16993 VDD.n2749 VDD.n64 19.3944
R16994 VDD.n2743 VDD.n64 19.3944
R16995 VDD.n2743 VDD.n2742 19.3944
R16996 VDD.n2742 VDD.n2741 19.3944
R16997 VDD.n2741 VDD.n75 19.3944
R16998 VDD.n2735 VDD.n75 19.3944
R16999 VDD.n2735 VDD.n2734 19.3944
R17000 VDD.n2734 VDD.n2733 19.3944
R17001 VDD.n2733 VDD.n85 19.3944
R17002 VDD.n2727 VDD.n85 19.3944
R17003 VDD.n2694 VDD.n121 19.3944
R17004 VDD.n2694 VDD.n125 19.3944
R17005 VDD.n128 VDD.n125 19.3944
R17006 VDD.n2687 VDD.n128 19.3944
R17007 VDD.n2687 VDD.n2686 19.3944
R17008 VDD.n2686 VDD.n2685 19.3944
R17009 VDD.n2685 VDD.n134 19.3944
R17010 VDD.n2711 VDD.n103 19.3944
R17011 VDD.n2711 VDD.n109 19.3944
R17012 VDD.n2706 VDD.n109 19.3944
R17013 VDD.n2706 VDD.n2705 19.3944
R17014 VDD.n2705 VDD.n2704 19.3944
R17015 VDD.n2704 VDD.n116 19.3944
R17016 VDD.n2699 VDD.n116 19.3944
R17017 VDD.n2724 VDD.n2723 19.3944
R17018 VDD.n2723 VDD.n2722 19.3944
R17019 VDD.n2722 VDD.n97 19.3944
R17020 VDD.n2717 VDD.n97 19.3944
R17021 VDD.n2717 VDD.n2716 19.3944
R17022 VDD.n2560 VDD.n216 19.3944
R17023 VDD.n2564 VDD.n216 19.3944
R17024 VDD.n2564 VDD.n207 19.3944
R17025 VDD.n2577 VDD.n207 19.3944
R17026 VDD.n2577 VDD.n205 19.3944
R17027 VDD.n2581 VDD.n205 19.3944
R17028 VDD.n2581 VDD.n195 19.3944
R17029 VDD.n2593 VDD.n195 19.3944
R17030 VDD.n2593 VDD.n193 19.3944
R17031 VDD.n2597 VDD.n193 19.3944
R17032 VDD.n2597 VDD.n183 19.3944
R17033 VDD.n2609 VDD.n183 19.3944
R17034 VDD.n2609 VDD.n181 19.3944
R17035 VDD.n2613 VDD.n181 19.3944
R17036 VDD.n2613 VDD.n171 19.3944
R17037 VDD.n2625 VDD.n171 19.3944
R17038 VDD.n2625 VDD.n169 19.3944
R17039 VDD.n2629 VDD.n169 19.3944
R17040 VDD.n2629 VDD.n158 19.3944
R17041 VDD.n2641 VDD.n158 19.3944
R17042 VDD.n2641 VDD.n156 19.3944
R17043 VDD.n2645 VDD.n156 19.3944
R17044 VDD.n2646 VDD.n2645 19.3944
R17045 VDD.n2647 VDD.n2646 19.3944
R17046 VDD.n2647 VDD.n154 19.3944
R17047 VDD.n2651 VDD.n154 19.3944
R17048 VDD.n2652 VDD.n2651 19.3944
R17049 VDD.n2653 VDD.n2652 19.3944
R17050 VDD.n2653 VDD.n151 19.3944
R17051 VDD.n2657 VDD.n151 19.3944
R17052 VDD.n2658 VDD.n2657 19.3944
R17053 VDD.n2659 VDD.n2658 19.3944
R17054 VDD.n2659 VDD.n148 19.3944
R17055 VDD.n2663 VDD.n148 19.3944
R17056 VDD.n2664 VDD.n2663 19.3944
R17057 VDD.n2665 VDD.n2664 19.3944
R17058 VDD.n2665 VDD.n145 19.3944
R17059 VDD.n2669 VDD.n145 19.3944
R17060 VDD.n2670 VDD.n2669 19.3944
R17061 VDD.n2671 VDD.n2670 19.3944
R17062 VDD.n2671 VDD.n142 19.3944
R17063 VDD.n2675 VDD.n142 19.3944
R17064 VDD.n2676 VDD.n2675 19.3944
R17065 VDD.n2677 VDD.n2676 19.3944
R17066 VDD.n1518 VDD.n1094 19.3944
R17067 VDD.n1522 VDD.n1094 19.3944
R17068 VDD.n1523 VDD.n1522 19.3944
R17069 VDD.n1526 VDD.n1523 19.3944
R17070 VDD.n1526 VDD.n1090 19.3944
R17071 VDD.n1536 VDD.n1533 19.3944
R17072 VDD.n1536 VDD.n1088 19.3944
R17073 VDD.n1540 VDD.n1088 19.3944
R17074 VDD.n1540 VDD.n1058 19.3944
R17075 VDD.n1572 VDD.n1058 19.3944
R17076 VDD.n1572 VDD.n1571 19.3944
R17077 VDD.n1571 VDD.n1570 19.3944
R17078 VDD.n1566 VDD.n1565 19.3944
R17079 VDD.n1565 VDD.n1564 19.3944
R17080 VDD.n1564 VDD.n1069 19.3944
R17081 VDD.n1560 VDD.n1069 19.3944
R17082 VDD.n1560 VDD.n1559 19.3944
R17083 VDD.n1559 VDD.n1558 19.3944
R17084 VDD.n1558 VDD.n1074 19.3944
R17085 VDD.n1321 VDD.n1220 19.3944
R17086 VDD.n1334 VDD.n1220 19.3944
R17087 VDD.n1334 VDD.n1218 19.3944
R17088 VDD.n1338 VDD.n1218 19.3944
R17089 VDD.n1338 VDD.n1209 19.3944
R17090 VDD.n1350 VDD.n1209 19.3944
R17091 VDD.n1350 VDD.n1207 19.3944
R17092 VDD.n1354 VDD.n1207 19.3944
R17093 VDD.n1354 VDD.n1197 19.3944
R17094 VDD.n1366 VDD.n1197 19.3944
R17095 VDD.n1366 VDD.n1195 19.3944
R17096 VDD.n1370 VDD.n1195 19.3944
R17097 VDD.n1370 VDD.n1185 19.3944
R17098 VDD.n1382 VDD.n1185 19.3944
R17099 VDD.n1382 VDD.n1183 19.3944
R17100 VDD.n1386 VDD.n1183 19.3944
R17101 VDD.n1386 VDD.n1173 19.3944
R17102 VDD.n1398 VDD.n1173 19.3944
R17103 VDD.n1398 VDD.n1171 19.3944
R17104 VDD.n1402 VDD.n1171 19.3944
R17105 VDD.n1402 VDD.n1161 19.3944
R17106 VDD.n1414 VDD.n1161 19.3944
R17107 VDD.n1414 VDD.n1159 19.3944
R17108 VDD.n1430 VDD.n1159 19.3944
R17109 VDD.n1430 VDD.n1149 19.3944
R17110 VDD.n1442 VDD.n1149 19.3944
R17111 VDD.n1442 VDD.n1147 19.3944
R17112 VDD.n1446 VDD.n1147 19.3944
R17113 VDD.n1446 VDD.n1137 19.3944
R17114 VDD.n1459 VDD.n1137 19.3944
R17115 VDD.n1459 VDD.n1135 19.3944
R17116 VDD.n1463 VDD.n1135 19.3944
R17117 VDD.n1463 VDD.n1126 19.3944
R17118 VDD.n1475 VDD.n1126 19.3944
R17119 VDD.n1475 VDD.n1124 19.3944
R17120 VDD.n1479 VDD.n1124 19.3944
R17121 VDD.n1479 VDD.n1113 19.3944
R17122 VDD.n1492 VDD.n1113 19.3944
R17123 VDD.n1492 VDD.n1111 19.3944
R17124 VDD.n1496 VDD.n1111 19.3944
R17125 VDD.n1496 VDD.n1100 19.3944
R17126 VDD.n1511 VDD.n1100 19.3944
R17127 VDD.n1511 VDD.n1098 19.3944
R17128 VDD.n1515 VDD.n1098 19.3944
R17129 VDD.n1291 VDD.n1255 18.8126
R17130 VDD.n2522 VDD.n2521 18.8126
R17131 VDD.n2698 VDD.n121 18.8126
R17132 VDD.n1566 VDD.n1064 18.8126
R17133 VDD.t117 VDD.n1187 16.8108
R17134 VDD.n1456 VDD.t128 16.8108
R17135 VDD.t108 VDD.n179 16.8108
R17136 VDD.n2754 VDD.t110 16.8108
R17137 VDD.n1396 VDD.t114 15.9488
R17138 VDD.n1440 VDD.t106 15.9488
R17139 VDD.n2631 VDD.t122 15.9488
R17140 VDD.n2763 VDD.t125 15.9488
R17141 VDD.n23 VDD.t124 15.5531
R17142 VDD.n23 VDD.t130 15.5531
R17143 VDD.n19 VDD.t127 15.5531
R17144 VDD.n19 VDD.t132 15.5531
R17145 VDD.n16 VDD.t123 15.5531
R17146 VDD.n16 VDD.t126 15.5531
R17147 VDD.n1422 VDD.t116 15.5531
R17148 VDD.n1422 VDD.t136 15.5531
R17149 VDD.n1418 VDD.t119 15.5531
R17150 VDD.n1418 VDD.t107 15.5531
R17151 VDD.n1415 VDD.t115 15.5531
R17152 VDD.n1415 VDD.t133 15.5531
R17153 VDD.n1592 VDD.n758 14.6557
R17154 VDD.n1598 VDD.n758 14.6557
R17155 VDD.n1598 VDD.n752 14.6557
R17156 VDD.n1604 VDD.n752 14.6557
R17157 VDD.n1604 VDD.n746 14.6557
R17158 VDD.n1610 VDD.n746 14.6557
R17159 VDD.n1610 VDD.n739 14.6557
R17160 VDD.n1616 VDD.n739 14.6557
R17161 VDD.n1616 VDD.n742 14.6557
R17162 VDD.n1622 VDD.n728 14.6557
R17163 VDD.n1628 VDD.n728 14.6557
R17164 VDD.n1628 VDD.n722 14.6557
R17165 VDD.n1634 VDD.n722 14.6557
R17166 VDD.n1640 VDD.n716 14.6557
R17167 VDD.n1640 VDD.n710 14.6557
R17168 VDD.n1646 VDD.n710 14.6557
R17169 VDD.n1646 VDD.n704 14.6557
R17170 VDD.n1652 VDD.n704 14.6557
R17171 VDD.n1652 VDD.n698 14.6557
R17172 VDD.n1658 VDD.n698 14.6557
R17173 VDD.n1658 VDD.n692 14.6557
R17174 VDD.n1664 VDD.n692 14.6557
R17175 VDD.n1664 VDD.n686 14.6557
R17176 VDD.n1670 VDD.n686 14.6557
R17177 VDD.n1670 VDD.n679 14.6557
R17178 VDD.n1676 VDD.n679 14.6557
R17179 VDD.n1676 VDD.n682 14.6557
R17180 VDD.n1682 VDD.n675 14.6557
R17181 VDD.n1688 VDD.n662 14.6557
R17182 VDD.n1694 VDD.n662 14.6557
R17183 VDD.n1694 VDD.n656 14.6557
R17184 VDD.n1700 VDD.n656 14.6557
R17185 VDD.n1700 VDD.n650 14.6557
R17186 VDD.n1706 VDD.n650 14.6557
R17187 VDD.n1706 VDD.n644 14.6557
R17188 VDD.n1712 VDD.n644 14.6557
R17189 VDD.n1712 VDD.n638 14.6557
R17190 VDD.n1718 VDD.n638 14.6557
R17191 VDD.n1718 VDD.n631 14.6557
R17192 VDD.n1724 VDD.n631 14.6557
R17193 VDD.n1724 VDD.n634 14.6557
R17194 VDD.n1730 VDD.n620 14.6557
R17195 VDD.n1736 VDD.n620 14.6557
R17196 VDD.n1742 VDD.n614 14.6557
R17197 VDD.n1742 VDD.n608 14.6557
R17198 VDD.n1748 VDD.n608 14.6557
R17199 VDD.n1748 VDD.n602 14.6557
R17200 VDD.n1754 VDD.n602 14.6557
R17201 VDD.n1754 VDD.n596 14.6557
R17202 VDD.n1760 VDD.n596 14.6557
R17203 VDD.n1760 VDD.n590 14.6557
R17204 VDD.n1766 VDD.n590 14.6557
R17205 VDD.n1766 VDD.n584 14.6557
R17206 VDD.n1772 VDD.n584 14.6557
R17207 VDD.n1772 VDD.n578 14.6557
R17208 VDD.n1778 VDD.n578 14.6557
R17209 VDD.n1778 VDD.n572 14.6557
R17210 VDD.n1784 VDD.n572 14.6557
R17211 VDD.n1790 VDD.n561 14.6557
R17212 VDD.n1796 VDD.n561 14.6557
R17213 VDD.n1796 VDD.n554 14.6557
R17214 VDD.n1840 VDD.n554 14.6557
R17215 VDD.n1840 VDD.n548 14.6557
R17216 VDD.n1846 VDD.n548 14.6557
R17217 VDD.n1846 VDD.n537 14.6557
R17218 VDD.n1888 VDD.n537 14.6557
R17219 VDD.n1888 VDD.n516 14.6557
R17220 VDD.n2200 VDD.n510 14.6557
R17221 VDD.n2206 VDD.n510 14.6557
R17222 VDD.n2206 VDD.n504 14.6557
R17223 VDD.n2212 VDD.n504 14.6557
R17224 VDD.n2212 VDD.n498 14.6557
R17225 VDD.n2218 VDD.n498 14.6557
R17226 VDD.n2218 VDD.n491 14.6557
R17227 VDD.n2224 VDD.n491 14.6557
R17228 VDD.n2224 VDD.n494 14.6557
R17229 VDD.n2236 VDD.n480 14.6557
R17230 VDD.n2236 VDD.n474 14.6557
R17231 VDD.n2242 VDD.n474 14.6557
R17232 VDD.n2242 VDD.n468 14.6557
R17233 VDD.n2248 VDD.n468 14.6557
R17234 VDD.n2248 VDD.n462 14.6557
R17235 VDD.n2254 VDD.n462 14.6557
R17236 VDD.n2254 VDD.n456 14.6557
R17237 VDD.n2260 VDD.n456 14.6557
R17238 VDD.n2260 VDD.n450 14.6557
R17239 VDD.n2266 VDD.n450 14.6557
R17240 VDD.n2266 VDD.n444 14.6557
R17241 VDD.n2272 VDD.n444 14.6557
R17242 VDD.n2272 VDD.n438 14.6557
R17243 VDD.n2278 VDD.n438 14.6557
R17244 VDD.n2284 VDD.n431 14.6557
R17245 VDD.n2284 VDD.n434 14.6557
R17246 VDD.n2290 VDD.n420 14.6557
R17247 VDD.n2296 VDD.n420 14.6557
R17248 VDD.n2296 VDD.n414 14.6557
R17249 VDD.n2302 VDD.n414 14.6557
R17250 VDD.n2302 VDD.n408 14.6557
R17251 VDD.n2308 VDD.n408 14.6557
R17252 VDD.n2308 VDD.n402 14.6557
R17253 VDD.n2314 VDD.n402 14.6557
R17254 VDD.n2314 VDD.n396 14.6557
R17255 VDD.n2320 VDD.n396 14.6557
R17256 VDD.n2320 VDD.n389 14.6557
R17257 VDD.n2326 VDD.n389 14.6557
R17258 VDD.n2326 VDD.n392 14.6557
R17259 VDD.n2332 VDD.n385 14.6557
R17260 VDD.n2338 VDD.n372 14.6557
R17261 VDD.n2344 VDD.n372 14.6557
R17262 VDD.n2344 VDD.n366 14.6557
R17263 VDD.n2350 VDD.n366 14.6557
R17264 VDD.n2350 VDD.n360 14.6557
R17265 VDD.n2356 VDD.n360 14.6557
R17266 VDD.n2356 VDD.n354 14.6557
R17267 VDD.n2362 VDD.n354 14.6557
R17268 VDD.n2362 VDD.n348 14.6557
R17269 VDD.n2368 VDD.n348 14.6557
R17270 VDD.n2368 VDD.n342 14.6557
R17271 VDD.n2374 VDD.n342 14.6557
R17272 VDD.n2374 VDD.n336 14.6557
R17273 VDD.n2380 VDD.n336 14.6557
R17274 VDD.n2386 VDD.n330 14.6557
R17275 VDD.n2386 VDD.n323 14.6557
R17276 VDD.n2392 VDD.n323 14.6557
R17277 VDD.n2392 VDD.n326 14.6557
R17278 VDD.n2398 VDD.n312 14.6557
R17279 VDD.n2404 VDD.n312 14.6557
R17280 VDD.n2404 VDD.n305 14.6557
R17281 VDD.n2435 VDD.n305 14.6557
R17282 VDD.n2435 VDD.n299 14.6557
R17283 VDD.n2441 VDD.n299 14.6557
R17284 VDD.n2441 VDD.n278 14.6557
R17285 VDD.n2482 VDD.n278 14.6557
R17286 VDD.n2482 VDD.n280 14.6557
R17287 VDD.t8 VDD.n614 13.7936
R17288 VDD.n2278 VDD.t26 13.7936
R17289 VDD.n1310 VDD.n1239 13.3823
R17290 VDD.n2539 VDD.n2538 13.3823
R17291 VDD.n2715 VDD.n103 13.3823
R17292 VDD.n1533 VDD.n1532 13.3823
R17293 VDD.n1682 VDD.t12 12.716
R17294 VDD.n634 VDD.t17 12.716
R17295 VDD.n2290 VDD.t28 12.716
R17296 VDD.n385 VDD.t35 12.716
R17297 VDD.n1311 VDD.n1310 12.6066
R17298 VDD.n2539 VDD.n229 12.6066
R17299 VDD.n2716 VDD.n2715 12.6066
R17300 VDD.n1532 VDD.n1090 12.6066
R17301 VDD.n1622 VDD.t43 11.8539
R17302 VDD.n937 VDD.t50 11.8539
R17303 VDD.n2230 VDD.t54 11.8539
R17304 VDD.n326 VDD.t94 11.8539
R17305 VDD.n1784 VDD.t20 11.6384
R17306 VDD.t24 VDD.n480 11.6384
R17307 VDD.n2553 VDD.n222 11.3952
R17308 VDD.n2502 VDD.n2501 11.3952
R17309 VDD.n1575 VDD.n1574 11.3949
R17310 VDD.n1055 VDD.n1054 11.3949
R17311 VDD.n1331 VDD.t74 11.2074
R17312 VDD.t90 VDD.n1102 11.2074
R17313 VDD.n2566 VDD.t61 11.2074
R17314 VDD.n87 VDD.t39 11.2074
R17315 VDD.n2167 VDD.n2166 10.6151
R17316 VDD.n2166 VDD.n2164 10.6151
R17317 VDD.n2164 VDD.n2163 10.6151
R17318 VDD.n2163 VDD.n2161 10.6151
R17319 VDD.n2161 VDD.n2160 10.6151
R17320 VDD.n2160 VDD.n2158 10.6151
R17321 VDD.n2158 VDD.n2157 10.6151
R17322 VDD.n2157 VDD.n2155 10.6151
R17323 VDD.n2155 VDD.n2154 10.6151
R17324 VDD.n2154 VDD.n2152 10.6151
R17325 VDD.n2152 VDD.n2151 10.6151
R17326 VDD.n2151 VDD.n2149 10.6151
R17327 VDD.n2149 VDD.n2148 10.6151
R17328 VDD.n2148 VDD.n2146 10.6151
R17329 VDD.n2146 VDD.n2145 10.6151
R17330 VDD.n2145 VDD.n2143 10.6151
R17331 VDD.n2143 VDD.n2142 10.6151
R17332 VDD.n2142 VDD.n2140 10.6151
R17333 VDD.n2140 VDD.n2139 10.6151
R17334 VDD.n2139 VDD.n2137 10.6151
R17335 VDD.n2137 VDD.n2136 10.6151
R17336 VDD.n2136 VDD.n2134 10.6151
R17337 VDD.n2134 VDD.n2133 10.6151
R17338 VDD.n2133 VDD.n2131 10.6151
R17339 VDD.n2131 VDD.n2130 10.6151
R17340 VDD.n2130 VDD.n2128 10.6151
R17341 VDD.n2128 VDD.n2127 10.6151
R17342 VDD.n2127 VDD.n2125 10.6151
R17343 VDD.n2125 VDD.n2124 10.6151
R17344 VDD.n2124 VDD.n2122 10.6151
R17345 VDD.n2122 VDD.n2121 10.6151
R17346 VDD.n2121 VDD.n2119 10.6151
R17347 VDD.n2119 VDD.n2118 10.6151
R17348 VDD.n2118 VDD.n2116 10.6151
R17349 VDD.n2116 VDD.n2115 10.6151
R17350 VDD.n2115 VDD.n2113 10.6151
R17351 VDD.n2113 VDD.n2112 10.6151
R17352 VDD.n2112 VDD.n2110 10.6151
R17353 VDD.n2110 VDD.n2109 10.6151
R17354 VDD.n2109 VDD.n2107 10.6151
R17355 VDD.n2107 VDD.n2106 10.6151
R17356 VDD.n2106 VDD.n2104 10.6151
R17357 VDD.n2104 VDD.n2103 10.6151
R17358 VDD.n2103 VDD.n2101 10.6151
R17359 VDD.n2101 VDD.n2100 10.6151
R17360 VDD.n2100 VDD.n2098 10.6151
R17361 VDD.n2098 VDD.n2097 10.6151
R17362 VDD.n2097 VDD.n2095 10.6151
R17363 VDD.n2095 VDD.n2094 10.6151
R17364 VDD.n2094 VDD.n2092 10.6151
R17365 VDD.n2092 VDD.n2091 10.6151
R17366 VDD.n2091 VDD.n2089 10.6151
R17367 VDD.n2089 VDD.n2088 10.6151
R17368 VDD.n2088 VDD.n2086 10.6151
R17369 VDD.n2086 VDD.n2085 10.6151
R17370 VDD.n2085 VDD.n2083 10.6151
R17371 VDD.n2083 VDD.n2082 10.6151
R17372 VDD.n2082 VDD.n2080 10.6151
R17373 VDD.n2080 VDD.n2079 10.6151
R17374 VDD.n2079 VDD.n2077 10.6151
R17375 VDD.n2077 VDD.n2076 10.6151
R17376 VDD.n2076 VDD.n2074 10.6151
R17377 VDD.n2074 VDD.n2073 10.6151
R17378 VDD.n2073 VDD.n2071 10.6151
R17379 VDD.n2071 VDD.n2070 10.6151
R17380 VDD.n2070 VDD.n2068 10.6151
R17381 VDD.n2068 VDD.n2067 10.6151
R17382 VDD.n2067 VDD.n2065 10.6151
R17383 VDD.n2065 VDD.n2064 10.6151
R17384 VDD.n2064 VDD.n2062 10.6151
R17385 VDD.n2062 VDD.n2061 10.6151
R17386 VDD.n2061 VDD.n297 10.6151
R17387 VDD.n2444 VDD.n297 10.6151
R17388 VDD.n2445 VDD.n2444 10.6151
R17389 VDD.n2446 VDD.n2445 10.6151
R17390 VDD.n2197 VDD.n2196 10.6151
R17391 VDD.n2196 VDD.n2050 10.6151
R17392 VDD.n2191 VDD.n2050 10.6151
R17393 VDD.n2191 VDD.n2190 10.6151
R17394 VDD.n2190 VDD.n2052 10.6151
R17395 VDD.n2185 VDD.n2052 10.6151
R17396 VDD.n2185 VDD.n2184 10.6151
R17397 VDD.n2184 VDD.n2183 10.6151
R17398 VDD.n2183 VDD.n2054 10.6151
R17399 VDD.n2177 VDD.n2054 10.6151
R17400 VDD.n2177 VDD.n2176 10.6151
R17401 VDD.n2176 VDD.n2175 10.6151
R17402 VDD.n2175 VDD.n2056 10.6151
R17403 VDD.n2169 VDD.n2168 10.6151
R17404 VDD.n2198 VDD.n508 10.6151
R17405 VDD.n2208 VDD.n508 10.6151
R17406 VDD.n2209 VDD.n2208 10.6151
R17407 VDD.n2210 VDD.n2209 10.6151
R17408 VDD.n2210 VDD.n496 10.6151
R17409 VDD.n2220 VDD.n496 10.6151
R17410 VDD.n2221 VDD.n2220 10.6151
R17411 VDD.n2222 VDD.n2221 10.6151
R17412 VDD.n2222 VDD.n484 10.6151
R17413 VDD.n2232 VDD.n484 10.6151
R17414 VDD.n2233 VDD.n2232 10.6151
R17415 VDD.n2234 VDD.n2233 10.6151
R17416 VDD.n2234 VDD.n472 10.6151
R17417 VDD.n2244 VDD.n472 10.6151
R17418 VDD.n2245 VDD.n2244 10.6151
R17419 VDD.n2246 VDD.n2245 10.6151
R17420 VDD.n2246 VDD.n460 10.6151
R17421 VDD.n2256 VDD.n460 10.6151
R17422 VDD.n2257 VDD.n2256 10.6151
R17423 VDD.n2258 VDD.n2257 10.6151
R17424 VDD.n2258 VDD.n448 10.6151
R17425 VDD.n2268 VDD.n448 10.6151
R17426 VDD.n2269 VDD.n2268 10.6151
R17427 VDD.n2270 VDD.n2269 10.6151
R17428 VDD.n2270 VDD.n436 10.6151
R17429 VDD.n2280 VDD.n436 10.6151
R17430 VDD.n2281 VDD.n2280 10.6151
R17431 VDD.n2282 VDD.n2281 10.6151
R17432 VDD.n2282 VDD.n424 10.6151
R17433 VDD.n2292 VDD.n424 10.6151
R17434 VDD.n2293 VDD.n2292 10.6151
R17435 VDD.n2294 VDD.n2293 10.6151
R17436 VDD.n2294 VDD.n412 10.6151
R17437 VDD.n2304 VDD.n412 10.6151
R17438 VDD.n2305 VDD.n2304 10.6151
R17439 VDD.n2306 VDD.n2305 10.6151
R17440 VDD.n2306 VDD.n400 10.6151
R17441 VDD.n2316 VDD.n400 10.6151
R17442 VDD.n2317 VDD.n2316 10.6151
R17443 VDD.n2318 VDD.n2317 10.6151
R17444 VDD.n2318 VDD.n387 10.6151
R17445 VDD.n2328 VDD.n387 10.6151
R17446 VDD.n2329 VDD.n2328 10.6151
R17447 VDD.n2330 VDD.n2329 10.6151
R17448 VDD.n2330 VDD.n376 10.6151
R17449 VDD.n2340 VDD.n376 10.6151
R17450 VDD.n2341 VDD.n2340 10.6151
R17451 VDD.n2342 VDD.n2341 10.6151
R17452 VDD.n2342 VDD.n364 10.6151
R17453 VDD.n2352 VDD.n364 10.6151
R17454 VDD.n2353 VDD.n2352 10.6151
R17455 VDD.n2354 VDD.n2353 10.6151
R17456 VDD.n2354 VDD.n352 10.6151
R17457 VDD.n2364 VDD.n352 10.6151
R17458 VDD.n2365 VDD.n2364 10.6151
R17459 VDD.n2366 VDD.n2365 10.6151
R17460 VDD.n2366 VDD.n340 10.6151
R17461 VDD.n2376 VDD.n340 10.6151
R17462 VDD.n2377 VDD.n2376 10.6151
R17463 VDD.n2378 VDD.n2377 10.6151
R17464 VDD.n2378 VDD.n328 10.6151
R17465 VDD.n2388 VDD.n328 10.6151
R17466 VDD.n2389 VDD.n2388 10.6151
R17467 VDD.n2390 VDD.n2389 10.6151
R17468 VDD.n2390 VDD.n316 10.6151
R17469 VDD.n2400 VDD.n316 10.6151
R17470 VDD.n2401 VDD.n2400 10.6151
R17471 VDD.n2402 VDD.n2401 10.6151
R17472 VDD.n2402 VDD.n303 10.6151
R17473 VDD.n2437 VDD.n303 10.6151
R17474 VDD.n2438 VDD.n2437 10.6151
R17475 VDD.n2439 VDD.n2438 10.6151
R17476 VDD.n2439 VDD.n284 10.6151
R17477 VDD.n2480 VDD.n284 10.6151
R17478 VDD.n2480 VDD.n2479 10.6151
R17479 VDD.n2478 VDD.n285 10.6151
R17480 VDD.n286 VDD.n285 10.6151
R17481 VDD.n2471 VDD.n286 10.6151
R17482 VDD.n2471 VDD.n2470 10.6151
R17483 VDD.n2470 VDD.n2469 10.6151
R17484 VDD.n2469 VDD.n288 10.6151
R17485 VDD.n2464 VDD.n288 10.6151
R17486 VDD.n2460 VDD.n290 10.6151
R17487 VDD.n2460 VDD.n2459 10.6151
R17488 VDD.n2459 VDD.n2458 10.6151
R17489 VDD.n2458 VDD.n292 10.6151
R17490 VDD.n2453 VDD.n292 10.6151
R17491 VDD.n2451 VDD.n2450 10.6151
R17492 VDD.n2422 VDD.n2408 10.6151
R17493 VDD.n2422 VDD.n2421 10.6151
R17494 VDD.n2421 VDD.n2420 10.6151
R17495 VDD.n2420 VDD.n2410 10.6151
R17496 VDD.n2415 VDD.n2410 10.6151
R17497 VDD.n2415 VDD.n2414 10.6151
R17498 VDD.n2414 VDD.n264 10.6151
R17499 VDD.n2500 VDD.n265 10.6151
R17500 VDD.n268 VDD.n265 10.6151
R17501 VDD.n2493 VDD.n268 10.6151
R17502 VDD.n2493 VDD.n2492 10.6151
R17503 VDD.n2492 VDD.n2491 10.6151
R17504 VDD.n2486 VDD.n274 10.6151
R17505 VDD.n2047 VDD.n2046 10.6151
R17506 VDD.n2046 VDD.n2045 10.6151
R17507 VDD.n2045 VDD.n2044 10.6151
R17508 VDD.n2044 VDD.n2042 10.6151
R17509 VDD.n2042 VDD.n2041 10.6151
R17510 VDD.n2041 VDD.n2039 10.6151
R17511 VDD.n2039 VDD.n2038 10.6151
R17512 VDD.n2038 VDD.n2036 10.6151
R17513 VDD.n2036 VDD.n2035 10.6151
R17514 VDD.n2035 VDD.n2033 10.6151
R17515 VDD.n2033 VDD.n2032 10.6151
R17516 VDD.n2032 VDD.n2030 10.6151
R17517 VDD.n2030 VDD.n2029 10.6151
R17518 VDD.n2029 VDD.n2027 10.6151
R17519 VDD.n2027 VDD.n2026 10.6151
R17520 VDD.n2026 VDD.n2024 10.6151
R17521 VDD.n2024 VDD.n2023 10.6151
R17522 VDD.n2023 VDD.n2021 10.6151
R17523 VDD.n2021 VDD.n2020 10.6151
R17524 VDD.n2020 VDD.n2018 10.6151
R17525 VDD.n2018 VDD.n2017 10.6151
R17526 VDD.n2017 VDD.n2015 10.6151
R17527 VDD.n2015 VDD.n2014 10.6151
R17528 VDD.n2014 VDD.n2012 10.6151
R17529 VDD.n2012 VDD.n2011 10.6151
R17530 VDD.n2011 VDD.n2009 10.6151
R17531 VDD.n2009 VDD.n2008 10.6151
R17532 VDD.n2008 VDD.n2006 10.6151
R17533 VDD.n2006 VDD.n2005 10.6151
R17534 VDD.n2005 VDD.n2003 10.6151
R17535 VDD.n2003 VDD.n2002 10.6151
R17536 VDD.n2002 VDD.n2000 10.6151
R17537 VDD.n2000 VDD.n1999 10.6151
R17538 VDD.n1999 VDD.n1997 10.6151
R17539 VDD.n1997 VDD.n1996 10.6151
R17540 VDD.n1996 VDD.n1994 10.6151
R17541 VDD.n1994 VDD.n1993 10.6151
R17542 VDD.n1993 VDD.n1991 10.6151
R17543 VDD.n1991 VDD.n1990 10.6151
R17544 VDD.n1990 VDD.n1988 10.6151
R17545 VDD.n1988 VDD.n1987 10.6151
R17546 VDD.n1987 VDD.n1985 10.6151
R17547 VDD.n1985 VDD.n1984 10.6151
R17548 VDD.n1984 VDD.n1982 10.6151
R17549 VDD.n1982 VDD.n1981 10.6151
R17550 VDD.n1981 VDD.n1979 10.6151
R17551 VDD.n1979 VDD.n1978 10.6151
R17552 VDD.n1978 VDD.n1976 10.6151
R17553 VDD.n1976 VDD.n1975 10.6151
R17554 VDD.n1975 VDD.n1973 10.6151
R17555 VDD.n1973 VDD.n1972 10.6151
R17556 VDD.n1972 VDD.n1970 10.6151
R17557 VDD.n1970 VDD.n1969 10.6151
R17558 VDD.n1969 VDD.n1967 10.6151
R17559 VDD.n1967 VDD.n1966 10.6151
R17560 VDD.n1966 VDD.n1964 10.6151
R17561 VDD.n1964 VDD.n1963 10.6151
R17562 VDD.n1963 VDD.n1961 10.6151
R17563 VDD.n1961 VDD.n1960 10.6151
R17564 VDD.n1960 VDD.n1958 10.6151
R17565 VDD.n1958 VDD.n1957 10.6151
R17566 VDD.n1957 VDD.n1955 10.6151
R17567 VDD.n1955 VDD.n1954 10.6151
R17568 VDD.n1954 VDD.n1952 10.6151
R17569 VDD.n1952 VDD.n1951 10.6151
R17570 VDD.n1951 VDD.n1949 10.6151
R17571 VDD.n1949 VDD.n1948 10.6151
R17572 VDD.n1948 VDD.n1946 10.6151
R17573 VDD.n1946 VDD.n1945 10.6151
R17574 VDD.n1945 VDD.n1943 10.6151
R17575 VDD.n1943 VDD.n1942 10.6151
R17576 VDD.n1942 VDD.n1940 10.6151
R17577 VDD.n1940 VDD.n276 10.6151
R17578 VDD.n2484 VDD.n276 10.6151
R17579 VDD.n2485 VDD.n2484 10.6151
R17580 VDD.n1909 VDD.n514 10.6151
R17581 VDD.n1914 VDD.n1909 10.6151
R17582 VDD.n1915 VDD.n1914 10.6151
R17583 VDD.n1916 VDD.n1915 10.6151
R17584 VDD.n1916 VDD.n1907 10.6151
R17585 VDD.n1922 VDD.n1907 10.6151
R17586 VDD.n1923 VDD.n1922 10.6151
R17587 VDD.n1924 VDD.n1923 10.6151
R17588 VDD.n1924 VDD.n1905 10.6151
R17589 VDD.n1930 VDD.n1905 10.6151
R17590 VDD.n1931 VDD.n1930 10.6151
R17591 VDD.n1932 VDD.n1931 10.6151
R17592 VDD.n1932 VDD.n1903 10.6151
R17593 VDD.n1939 VDD.n1938 10.6151
R17594 VDD.n2203 VDD.n2202 10.6151
R17595 VDD.n2204 VDD.n2203 10.6151
R17596 VDD.n2204 VDD.n502 10.6151
R17597 VDD.n2214 VDD.n502 10.6151
R17598 VDD.n2215 VDD.n2214 10.6151
R17599 VDD.n2216 VDD.n2215 10.6151
R17600 VDD.n2216 VDD.n489 10.6151
R17601 VDD.n2226 VDD.n489 10.6151
R17602 VDD.n2227 VDD.n2226 10.6151
R17603 VDD.n2228 VDD.n2227 10.6151
R17604 VDD.n2228 VDD.n478 10.6151
R17605 VDD.n2238 VDD.n478 10.6151
R17606 VDD.n2239 VDD.n2238 10.6151
R17607 VDD.n2240 VDD.n2239 10.6151
R17608 VDD.n2240 VDD.n466 10.6151
R17609 VDD.n2250 VDD.n466 10.6151
R17610 VDD.n2251 VDD.n2250 10.6151
R17611 VDD.n2252 VDD.n2251 10.6151
R17612 VDD.n2252 VDD.n454 10.6151
R17613 VDD.n2262 VDD.n454 10.6151
R17614 VDD.n2263 VDD.n2262 10.6151
R17615 VDD.n2264 VDD.n2263 10.6151
R17616 VDD.n2264 VDD.n442 10.6151
R17617 VDD.n2274 VDD.n442 10.6151
R17618 VDD.n2275 VDD.n2274 10.6151
R17619 VDD.n2276 VDD.n2275 10.6151
R17620 VDD.n2276 VDD.n429 10.6151
R17621 VDD.n2286 VDD.n429 10.6151
R17622 VDD.n2287 VDD.n2286 10.6151
R17623 VDD.n2288 VDD.n2287 10.6151
R17624 VDD.n2288 VDD.n418 10.6151
R17625 VDD.n2298 VDD.n418 10.6151
R17626 VDD.n2299 VDD.n2298 10.6151
R17627 VDD.n2300 VDD.n2299 10.6151
R17628 VDD.n2300 VDD.n406 10.6151
R17629 VDD.n2310 VDD.n406 10.6151
R17630 VDD.n2311 VDD.n2310 10.6151
R17631 VDD.n2312 VDD.n2311 10.6151
R17632 VDD.n2312 VDD.n394 10.6151
R17633 VDD.n2322 VDD.n394 10.6151
R17634 VDD.n2323 VDD.n2322 10.6151
R17635 VDD.n2324 VDD.n2323 10.6151
R17636 VDD.n2324 VDD.n381 10.6151
R17637 VDD.n2334 VDD.n381 10.6151
R17638 VDD.n2335 VDD.n2334 10.6151
R17639 VDD.n2336 VDD.n2335 10.6151
R17640 VDD.n2336 VDD.n370 10.6151
R17641 VDD.n2346 VDD.n370 10.6151
R17642 VDD.n2347 VDD.n2346 10.6151
R17643 VDD.n2348 VDD.n2347 10.6151
R17644 VDD.n2348 VDD.n358 10.6151
R17645 VDD.n2358 VDD.n358 10.6151
R17646 VDD.n2359 VDD.n2358 10.6151
R17647 VDD.n2360 VDD.n2359 10.6151
R17648 VDD.n2360 VDD.n346 10.6151
R17649 VDD.n2370 VDD.n346 10.6151
R17650 VDD.n2371 VDD.n2370 10.6151
R17651 VDD.n2372 VDD.n2371 10.6151
R17652 VDD.n2372 VDD.n334 10.6151
R17653 VDD.n2382 VDD.n334 10.6151
R17654 VDD.n2383 VDD.n2382 10.6151
R17655 VDD.n2384 VDD.n2383 10.6151
R17656 VDD.n2384 VDD.n321 10.6151
R17657 VDD.n2394 VDD.n321 10.6151
R17658 VDD.n2395 VDD.n2394 10.6151
R17659 VDD.n2396 VDD.n2395 10.6151
R17660 VDD.n2396 VDD.n310 10.6151
R17661 VDD.n2406 VDD.n310 10.6151
R17662 VDD.n2407 VDD.n2406 10.6151
R17663 VDD.n2433 VDD.n2407 10.6151
R17664 VDD.n2433 VDD.n2432 10.6151
R17665 VDD.n2432 VDD.n2431 10.6151
R17666 VDD.n2431 VDD.n2430 10.6151
R17667 VDD.n2430 VDD.n2428 10.6151
R17668 VDD.n2428 VDD.n2427 10.6151
R17669 VDD.n1590 VDD.n756 10.6151
R17670 VDD.n1600 VDD.n756 10.6151
R17671 VDD.n1601 VDD.n1600 10.6151
R17672 VDD.n1602 VDD.n1601 10.6151
R17673 VDD.n1602 VDD.n744 10.6151
R17674 VDD.n1612 VDD.n744 10.6151
R17675 VDD.n1613 VDD.n1612 10.6151
R17676 VDD.n1614 VDD.n1613 10.6151
R17677 VDD.n1614 VDD.n732 10.6151
R17678 VDD.n1624 VDD.n732 10.6151
R17679 VDD.n1625 VDD.n1624 10.6151
R17680 VDD.n1626 VDD.n1625 10.6151
R17681 VDD.n1626 VDD.n720 10.6151
R17682 VDD.n1636 VDD.n720 10.6151
R17683 VDD.n1637 VDD.n1636 10.6151
R17684 VDD.n1638 VDD.n1637 10.6151
R17685 VDD.n1638 VDD.n708 10.6151
R17686 VDD.n1648 VDD.n708 10.6151
R17687 VDD.n1649 VDD.n1648 10.6151
R17688 VDD.n1650 VDD.n1649 10.6151
R17689 VDD.n1650 VDD.n696 10.6151
R17690 VDD.n1660 VDD.n696 10.6151
R17691 VDD.n1661 VDD.n1660 10.6151
R17692 VDD.n1662 VDD.n1661 10.6151
R17693 VDD.n1662 VDD.n684 10.6151
R17694 VDD.n1672 VDD.n684 10.6151
R17695 VDD.n1673 VDD.n1672 10.6151
R17696 VDD.n1674 VDD.n1673 10.6151
R17697 VDD.n1674 VDD.n671 10.6151
R17698 VDD.n1684 VDD.n671 10.6151
R17699 VDD.n1685 VDD.n1684 10.6151
R17700 VDD.n1686 VDD.n1685 10.6151
R17701 VDD.n1686 VDD.n660 10.6151
R17702 VDD.n1696 VDD.n660 10.6151
R17703 VDD.n1697 VDD.n1696 10.6151
R17704 VDD.n1698 VDD.n1697 10.6151
R17705 VDD.n1698 VDD.n648 10.6151
R17706 VDD.n1708 VDD.n648 10.6151
R17707 VDD.n1709 VDD.n1708 10.6151
R17708 VDD.n1710 VDD.n1709 10.6151
R17709 VDD.n1710 VDD.n636 10.6151
R17710 VDD.n1720 VDD.n636 10.6151
R17711 VDD.n1721 VDD.n1720 10.6151
R17712 VDD.n1722 VDD.n1721 10.6151
R17713 VDD.n1722 VDD.n624 10.6151
R17714 VDD.n1732 VDD.n624 10.6151
R17715 VDD.n1733 VDD.n1732 10.6151
R17716 VDD.n1734 VDD.n1733 10.6151
R17717 VDD.n1734 VDD.n612 10.6151
R17718 VDD.n1744 VDD.n612 10.6151
R17719 VDD.n1745 VDD.n1744 10.6151
R17720 VDD.n1746 VDD.n1745 10.6151
R17721 VDD.n1746 VDD.n600 10.6151
R17722 VDD.n1756 VDD.n600 10.6151
R17723 VDD.n1757 VDD.n1756 10.6151
R17724 VDD.n1758 VDD.n1757 10.6151
R17725 VDD.n1758 VDD.n588 10.6151
R17726 VDD.n1768 VDD.n588 10.6151
R17727 VDD.n1769 VDD.n1768 10.6151
R17728 VDD.n1770 VDD.n1769 10.6151
R17729 VDD.n1770 VDD.n576 10.6151
R17730 VDD.n1780 VDD.n576 10.6151
R17731 VDD.n1781 VDD.n1780 10.6151
R17732 VDD.n1782 VDD.n1781 10.6151
R17733 VDD.n1782 VDD.n565 10.6151
R17734 VDD.n1792 VDD.n565 10.6151
R17735 VDD.n1793 VDD.n1792 10.6151
R17736 VDD.n1794 VDD.n1793 10.6151
R17737 VDD.n1794 VDD.n552 10.6151
R17738 VDD.n1842 VDD.n552 10.6151
R17739 VDD.n1843 VDD.n1842 10.6151
R17740 VDD.n1844 VDD.n1843 10.6151
R17741 VDD.n1844 VDD.n542 10.6151
R17742 VDD.n1886 VDD.n542 10.6151
R17743 VDD.n1886 VDD.n1885 10.6151
R17744 VDD.n1884 VDD.n1882 10.6151
R17745 VDD.n1882 VDD.n1879 10.6151
R17746 VDD.n1879 VDD.n1878 10.6151
R17747 VDD.n1878 VDD.n1875 10.6151
R17748 VDD.n1875 VDD.n1874 10.6151
R17749 VDD.n1874 VDD.n1871 10.6151
R17750 VDD.n1871 VDD.n1870 10.6151
R17751 VDD.n1870 VDD.n1867 10.6151
R17752 VDD.n1867 VDD.n1866 10.6151
R17753 VDD.n1866 VDD.n1863 10.6151
R17754 VDD.n1863 VDD.n1862 10.6151
R17755 VDD.n1862 VDD.n1859 10.6151
R17756 VDD.n1859 VDD.n1858 10.6151
R17757 VDD.n1855 VDD.n1854 10.6151
R17758 VDD.n832 VDD.n830 10.6151
R17759 VDD.n833 VDD.n832 10.6151
R17760 VDD.n835 VDD.n833 10.6151
R17761 VDD.n836 VDD.n835 10.6151
R17762 VDD.n838 VDD.n836 10.6151
R17763 VDD.n839 VDD.n838 10.6151
R17764 VDD.n841 VDD.n839 10.6151
R17765 VDD.n842 VDD.n841 10.6151
R17766 VDD.n844 VDD.n842 10.6151
R17767 VDD.n845 VDD.n844 10.6151
R17768 VDD.n847 VDD.n845 10.6151
R17769 VDD.n848 VDD.n847 10.6151
R17770 VDD.n850 VDD.n848 10.6151
R17771 VDD.n851 VDD.n850 10.6151
R17772 VDD.n853 VDD.n851 10.6151
R17773 VDD.n854 VDD.n853 10.6151
R17774 VDD.n856 VDD.n854 10.6151
R17775 VDD.n857 VDD.n856 10.6151
R17776 VDD.n859 VDD.n857 10.6151
R17777 VDD.n860 VDD.n859 10.6151
R17778 VDD.n862 VDD.n860 10.6151
R17779 VDD.n863 VDD.n862 10.6151
R17780 VDD.n865 VDD.n863 10.6151
R17781 VDD.n866 VDD.n865 10.6151
R17782 VDD.n868 VDD.n866 10.6151
R17783 VDD.n869 VDD.n868 10.6151
R17784 VDD.n871 VDD.n869 10.6151
R17785 VDD.n872 VDD.n871 10.6151
R17786 VDD.n874 VDD.n872 10.6151
R17787 VDD.n875 VDD.n874 10.6151
R17788 VDD.n877 VDD.n875 10.6151
R17789 VDD.n878 VDD.n877 10.6151
R17790 VDD.n880 VDD.n878 10.6151
R17791 VDD.n881 VDD.n880 10.6151
R17792 VDD.n883 VDD.n881 10.6151
R17793 VDD.n884 VDD.n883 10.6151
R17794 VDD.n886 VDD.n884 10.6151
R17795 VDD.n887 VDD.n886 10.6151
R17796 VDD.n889 VDD.n887 10.6151
R17797 VDD.n890 VDD.n889 10.6151
R17798 VDD.n892 VDD.n890 10.6151
R17799 VDD.n893 VDD.n892 10.6151
R17800 VDD.n895 VDD.n893 10.6151
R17801 VDD.n896 VDD.n895 10.6151
R17802 VDD.n898 VDD.n896 10.6151
R17803 VDD.n899 VDD.n898 10.6151
R17804 VDD.n901 VDD.n899 10.6151
R17805 VDD.n902 VDD.n901 10.6151
R17806 VDD.n904 VDD.n902 10.6151
R17807 VDD.n905 VDD.n904 10.6151
R17808 VDD.n907 VDD.n905 10.6151
R17809 VDD.n908 VDD.n907 10.6151
R17810 VDD.n910 VDD.n908 10.6151
R17811 VDD.n911 VDD.n910 10.6151
R17812 VDD.n913 VDD.n911 10.6151
R17813 VDD.n914 VDD.n913 10.6151
R17814 VDD.n916 VDD.n914 10.6151
R17815 VDD.n917 VDD.n916 10.6151
R17816 VDD.n919 VDD.n917 10.6151
R17817 VDD.n920 VDD.n919 10.6151
R17818 VDD.n922 VDD.n920 10.6151
R17819 VDD.n923 VDD.n922 10.6151
R17820 VDD.n925 VDD.n923 10.6151
R17821 VDD.n926 VDD.n925 10.6151
R17822 VDD.n935 VDD.n926 10.6151
R17823 VDD.n935 VDD.n934 10.6151
R17824 VDD.n934 VDD.n933 10.6151
R17825 VDD.n933 VDD.n931 10.6151
R17826 VDD.n931 VDD.n930 10.6151
R17827 VDD.n930 VDD.n928 10.6151
R17828 VDD.n928 VDD.n927 10.6151
R17829 VDD.n927 VDD.n546 10.6151
R17830 VDD.n1849 VDD.n546 10.6151
R17831 VDD.n1850 VDD.n1849 10.6151
R17832 VDD.n1851 VDD.n1850 10.6151
R17833 VDD.n1589 VDD.n1588 10.6151
R17834 VDD.n1588 VDD.n768 10.6151
R17835 VDD.n1583 VDD.n768 10.6151
R17836 VDD.n1583 VDD.n1582 10.6151
R17837 VDD.n1582 VDD.n770 10.6151
R17838 VDD.n1577 VDD.n770 10.6151
R17839 VDD.n1577 VDD.n1576 10.6151
R17840 VDD.n813 VDD.n772 10.6151
R17841 VDD.n813 VDD.n810 10.6151
R17842 VDD.n819 VDD.n810 10.6151
R17843 VDD.n820 VDD.n819 10.6151
R17844 VDD.n824 VDD.n820 10.6151
R17845 VDD.n829 VDD.n808 10.6151
R17846 VDD.n1829 VDD.n1828 10.6151
R17847 VDD.n1828 VDD.n1825 10.6151
R17848 VDD.n1825 VDD.n1824 10.6151
R17849 VDD.n1824 VDD.n1821 10.6151
R17850 VDD.n1821 VDD.n1820 10.6151
R17851 VDD.n1820 VDD.n1817 10.6151
R17852 VDD.n1817 VDD.n1816 10.6151
R17853 VDD.n1816 VDD.n1813 10.6151
R17854 VDD.n1813 VDD.n1812 10.6151
R17855 VDD.n1812 VDD.n1809 10.6151
R17856 VDD.n1809 VDD.n1808 10.6151
R17857 VDD.n1808 VDD.n1805 10.6151
R17858 VDD.n1805 VDD.n1804 10.6151
R17859 VDD.n1892 VDD.n534 10.6151
R17860 VDD.n1036 VDD.n1035 10.6151
R17861 VDD.n1035 VDD.n1033 10.6151
R17862 VDD.n1033 VDD.n1032 10.6151
R17863 VDD.n1032 VDD.n1030 10.6151
R17864 VDD.n1030 VDD.n1029 10.6151
R17865 VDD.n1029 VDD.n1027 10.6151
R17866 VDD.n1027 VDD.n1026 10.6151
R17867 VDD.n1026 VDD.n1024 10.6151
R17868 VDD.n1024 VDD.n1023 10.6151
R17869 VDD.n1023 VDD.n1021 10.6151
R17870 VDD.n1021 VDD.n1020 10.6151
R17871 VDD.n1020 VDD.n1018 10.6151
R17872 VDD.n1018 VDD.n1017 10.6151
R17873 VDD.n1017 VDD.n1015 10.6151
R17874 VDD.n1015 VDD.n1014 10.6151
R17875 VDD.n1014 VDD.n1012 10.6151
R17876 VDD.n1012 VDD.n1011 10.6151
R17877 VDD.n1011 VDD.n1009 10.6151
R17878 VDD.n1009 VDD.n1008 10.6151
R17879 VDD.n1008 VDD.n1006 10.6151
R17880 VDD.n1006 VDD.n1005 10.6151
R17881 VDD.n1005 VDD.n1003 10.6151
R17882 VDD.n1003 VDD.n1002 10.6151
R17883 VDD.n1002 VDD.n1000 10.6151
R17884 VDD.n1000 VDD.n999 10.6151
R17885 VDD.n999 VDD.n997 10.6151
R17886 VDD.n997 VDD.n996 10.6151
R17887 VDD.n996 VDD.n994 10.6151
R17888 VDD.n994 VDD.n993 10.6151
R17889 VDD.n993 VDD.n991 10.6151
R17890 VDD.n991 VDD.n990 10.6151
R17891 VDD.n990 VDD.n988 10.6151
R17892 VDD.n988 VDD.n987 10.6151
R17893 VDD.n987 VDD.n985 10.6151
R17894 VDD.n985 VDD.n984 10.6151
R17895 VDD.n984 VDD.n982 10.6151
R17896 VDD.n982 VDD.n981 10.6151
R17897 VDD.n981 VDD.n979 10.6151
R17898 VDD.n979 VDD.n978 10.6151
R17899 VDD.n978 VDD.n976 10.6151
R17900 VDD.n976 VDD.n975 10.6151
R17901 VDD.n975 VDD.n973 10.6151
R17902 VDD.n973 VDD.n972 10.6151
R17903 VDD.n972 VDD.n970 10.6151
R17904 VDD.n970 VDD.n969 10.6151
R17905 VDD.n969 VDD.n967 10.6151
R17906 VDD.n967 VDD.n966 10.6151
R17907 VDD.n966 VDD.n964 10.6151
R17908 VDD.n964 VDD.n963 10.6151
R17909 VDD.n963 VDD.n961 10.6151
R17910 VDD.n961 VDD.n960 10.6151
R17911 VDD.n960 VDD.n958 10.6151
R17912 VDD.n958 VDD.n957 10.6151
R17913 VDD.n957 VDD.n955 10.6151
R17914 VDD.n955 VDD.n954 10.6151
R17915 VDD.n954 VDD.n952 10.6151
R17916 VDD.n952 VDD.n951 10.6151
R17917 VDD.n951 VDD.n949 10.6151
R17918 VDD.n949 VDD.n948 10.6151
R17919 VDD.n948 VDD.n946 10.6151
R17920 VDD.n946 VDD.n945 10.6151
R17921 VDD.n945 VDD.n943 10.6151
R17922 VDD.n943 VDD.n942 10.6151
R17923 VDD.n942 VDD.n940 10.6151
R17924 VDD.n940 VDD.n939 10.6151
R17925 VDD.n939 VDD.n807 10.6151
R17926 VDD.n807 VDD.n806 10.6151
R17927 VDD.n806 VDD.n804 10.6151
R17928 VDD.n804 VDD.n803 10.6151
R17929 VDD.n803 VDD.n801 10.6151
R17930 VDD.n801 VDD.n800 10.6151
R17931 VDD.n800 VDD.n798 10.6151
R17932 VDD.n798 VDD.n535 10.6151
R17933 VDD.n1890 VDD.n535 10.6151
R17934 VDD.n1891 VDD.n1890 10.6151
R17935 VDD.n780 VDD.n762 10.6151
R17936 VDD.n781 VDD.n780 10.6151
R17937 VDD.n781 VDD.n777 10.6151
R17938 VDD.n787 VDD.n777 10.6151
R17939 VDD.n788 VDD.n787 10.6151
R17940 VDD.n789 VDD.n788 10.6151
R17941 VDD.n789 VDD.n774 10.6151
R17942 VDD.n1053 VDD.n775 10.6151
R17943 VDD.n1048 VDD.n775 10.6151
R17944 VDD.n1048 VDD.n1047 10.6151
R17945 VDD.n1047 VDD.n794 10.6151
R17946 VDD.n1042 VDD.n794 10.6151
R17947 VDD.n1040 VDD.n1039 10.6151
R17948 VDD.n1595 VDD.n1594 10.6151
R17949 VDD.n1596 VDD.n1595 10.6151
R17950 VDD.n1596 VDD.n750 10.6151
R17951 VDD.n1606 VDD.n750 10.6151
R17952 VDD.n1607 VDD.n1606 10.6151
R17953 VDD.n1608 VDD.n1607 10.6151
R17954 VDD.n1608 VDD.n737 10.6151
R17955 VDD.n1618 VDD.n737 10.6151
R17956 VDD.n1619 VDD.n1618 10.6151
R17957 VDD.n1620 VDD.n1619 10.6151
R17958 VDD.n1620 VDD.n726 10.6151
R17959 VDD.n1630 VDD.n726 10.6151
R17960 VDD.n1631 VDD.n1630 10.6151
R17961 VDD.n1632 VDD.n1631 10.6151
R17962 VDD.n1632 VDD.n714 10.6151
R17963 VDD.n1642 VDD.n714 10.6151
R17964 VDD.n1643 VDD.n1642 10.6151
R17965 VDD.n1644 VDD.n1643 10.6151
R17966 VDD.n1644 VDD.n702 10.6151
R17967 VDD.n1654 VDD.n702 10.6151
R17968 VDD.n1655 VDD.n1654 10.6151
R17969 VDD.n1656 VDD.n1655 10.6151
R17970 VDD.n1656 VDD.n690 10.6151
R17971 VDD.n1666 VDD.n690 10.6151
R17972 VDD.n1667 VDD.n1666 10.6151
R17973 VDD.n1668 VDD.n1667 10.6151
R17974 VDD.n1668 VDD.n677 10.6151
R17975 VDD.n1678 VDD.n677 10.6151
R17976 VDD.n1679 VDD.n1678 10.6151
R17977 VDD.n1680 VDD.n1679 10.6151
R17978 VDD.n1680 VDD.n666 10.6151
R17979 VDD.n1690 VDD.n666 10.6151
R17980 VDD.n1691 VDD.n1690 10.6151
R17981 VDD.n1692 VDD.n1691 10.6151
R17982 VDD.n1692 VDD.n654 10.6151
R17983 VDD.n1702 VDD.n654 10.6151
R17984 VDD.n1703 VDD.n1702 10.6151
R17985 VDD.n1704 VDD.n1703 10.6151
R17986 VDD.n1704 VDD.n642 10.6151
R17987 VDD.n1714 VDD.n642 10.6151
R17988 VDD.n1715 VDD.n1714 10.6151
R17989 VDD.n1716 VDD.n1715 10.6151
R17990 VDD.n1716 VDD.n629 10.6151
R17991 VDD.n1726 VDD.n629 10.6151
R17992 VDD.n1727 VDD.n1726 10.6151
R17993 VDD.n1728 VDD.n1727 10.6151
R17994 VDD.n1728 VDD.n618 10.6151
R17995 VDD.n1738 VDD.n618 10.6151
R17996 VDD.n1739 VDD.n1738 10.6151
R17997 VDD.n1740 VDD.n1739 10.6151
R17998 VDD.n1740 VDD.n606 10.6151
R17999 VDD.n1750 VDD.n606 10.6151
R18000 VDD.n1751 VDD.n1750 10.6151
R18001 VDD.n1752 VDD.n1751 10.6151
R18002 VDD.n1752 VDD.n594 10.6151
R18003 VDD.n1762 VDD.n594 10.6151
R18004 VDD.n1763 VDD.n1762 10.6151
R18005 VDD.n1764 VDD.n1763 10.6151
R18006 VDD.n1764 VDD.n582 10.6151
R18007 VDD.n1774 VDD.n582 10.6151
R18008 VDD.n1775 VDD.n1774 10.6151
R18009 VDD.n1776 VDD.n1775 10.6151
R18010 VDD.n1776 VDD.n570 10.6151
R18011 VDD.n1786 VDD.n570 10.6151
R18012 VDD.n1787 VDD.n1786 10.6151
R18013 VDD.n1788 VDD.n1787 10.6151
R18014 VDD.n1788 VDD.n559 10.6151
R18015 VDD.n1798 VDD.n559 10.6151
R18016 VDD.n1799 VDD.n1798 10.6151
R18017 VDD.n1838 VDD.n1799 10.6151
R18018 VDD.n1838 VDD.n1837 10.6151
R18019 VDD.n1837 VDD.n1836 10.6151
R18020 VDD.n1836 VDD.n1835 10.6151
R18021 VDD.n1835 VDD.n1833 10.6151
R18022 VDD.n1833 VDD.n1832 10.6151
R18023 VDD.n1340 VDD.t74 10.3453
R18024 VDD.n1498 VDD.t90 10.3453
R18025 VDD.n2575 VDD.t61 10.3453
R18026 VDD.n2737 VDD.t39 10.3453
R18027 VDD.n1688 VDD.t13 9.91429
R18028 VDD.n392 VDD.t22 9.91429
R18029 VDD.n7 VDD.t7 9.70349
R18030 VDD.n7 VDD.t16 9.70349
R18031 VDD.n8 VDD.t11 9.70349
R18032 VDD.n8 VDD.t5 9.70349
R18033 VDD.n10 VDD.t23 9.70349
R18034 VDD.n10 VDD.t34 9.70349
R18035 VDD.n12 VDD.t25 9.70349
R18036 VDD.n12 VDD.t27 9.70349
R18037 VDD.n5 VDD.t9 9.70349
R18038 VDD.n5 VDD.t21 9.70349
R18039 VDD.n3 VDD.t3 9.70349
R18040 VDD.n3 VDD.t14 9.70349
R18041 VDD.n1 VDD.t32 9.70349
R18042 VDD.n1 VDD.t19 9.70349
R18043 VDD.n0 VDD.t37 9.70349
R18044 VDD.n0 VDD.t30 9.70349
R18045 VDD.n2562 VDD.n216 9.3005
R18046 VDD.n2564 VDD.n2563 9.3005
R18047 VDD.n207 VDD.n206 9.3005
R18048 VDD.n2578 VDD.n2577 9.3005
R18049 VDD.n2579 VDD.n205 9.3005
R18050 VDD.n2581 VDD.n2580 9.3005
R18051 VDD.n195 VDD.n194 9.3005
R18052 VDD.n2594 VDD.n2593 9.3005
R18053 VDD.n2595 VDD.n193 9.3005
R18054 VDD.n2597 VDD.n2596 9.3005
R18055 VDD.n183 VDD.n182 9.3005
R18056 VDD.n2610 VDD.n2609 9.3005
R18057 VDD.n2611 VDD.n181 9.3005
R18058 VDD.n2613 VDD.n2612 9.3005
R18059 VDD.n171 VDD.n170 9.3005
R18060 VDD.n2626 VDD.n2625 9.3005
R18061 VDD.n2627 VDD.n169 9.3005
R18062 VDD.n2629 VDD.n2628 9.3005
R18063 VDD.n158 VDD.n157 9.3005
R18064 VDD.n2642 VDD.n2641 9.3005
R18065 VDD.n2643 VDD.n156 9.3005
R18066 VDD.n2645 VDD.n2644 9.3005
R18067 VDD.n2646 VDD.n155 9.3005
R18068 VDD.n2648 VDD.n2647 9.3005
R18069 VDD.n2649 VDD.n154 9.3005
R18070 VDD.n2651 VDD.n2650 9.3005
R18071 VDD.n2652 VDD.n152 9.3005
R18072 VDD.n2654 VDD.n2653 9.3005
R18073 VDD.n2655 VDD.n151 9.3005
R18074 VDD.n2657 VDD.n2656 9.3005
R18075 VDD.n2658 VDD.n149 9.3005
R18076 VDD.n2660 VDD.n2659 9.3005
R18077 VDD.n2661 VDD.n148 9.3005
R18078 VDD.n2663 VDD.n2662 9.3005
R18079 VDD.n2664 VDD.n146 9.3005
R18080 VDD.n2666 VDD.n2665 9.3005
R18081 VDD.n2667 VDD.n145 9.3005
R18082 VDD.n2669 VDD.n2668 9.3005
R18083 VDD.n2670 VDD.n143 9.3005
R18084 VDD.n2672 VDD.n2671 9.3005
R18085 VDD.n2673 VDD.n142 9.3005
R18086 VDD.n2675 VDD.n2674 9.3005
R18087 VDD.n2676 VDD.n140 9.3005
R18088 VDD.n2678 VDD.n2677 9.3005
R18089 VDD.n2561 VDD.n2560 9.3005
R18090 VDD.n2723 VDD.n94 9.3005
R18091 VDD.n2722 VDD.n96 9.3005
R18092 VDD.n100 VDD.n97 9.3005
R18093 VDD.n2717 VDD.n101 9.3005
R18094 VDD.n2716 VDD.n102 9.3005
R18095 VDD.n2715 VDD.n2714 9.3005
R18096 VDD.n2713 VDD.n103 9.3005
R18097 VDD.n2712 VDD.n2711 9.3005
R18098 VDD.n109 VDD.n108 9.3005
R18099 VDD.n2706 VDD.n113 9.3005
R18100 VDD.n2705 VDD.n114 9.3005
R18101 VDD.n2704 VDD.n115 9.3005
R18102 VDD.n119 VDD.n116 9.3005
R18103 VDD.n2699 VDD.n120 9.3005
R18104 VDD.n2698 VDD.n2697 9.3005
R18105 VDD.n2696 VDD.n121 9.3005
R18106 VDD.n2695 VDD.n2694 9.3005
R18107 VDD.n125 VDD.n124 9.3005
R18108 VDD.n130 VDD.n128 9.3005
R18109 VDD.n2687 VDD.n131 9.3005
R18110 VDD.n2686 VDD.n132 9.3005
R18111 VDD.n2685 VDD.n133 9.3005
R18112 VDD.n139 VDD.n134 9.3005
R18113 VDD.n2680 VDD.n2679 9.3005
R18114 VDD.n2725 VDD.n2724 9.3005
R18115 VDD.n30 VDD.n28 9.3005
R18116 VDD.n2767 VDD.n39 9.3005
R18117 VDD.n2766 VDD.n40 9.3005
R18118 VDD.n2765 VDD.n41 9.3005
R18119 VDD.n49 VDD.n42 9.3005
R18120 VDD.n2759 VDD.n50 9.3005
R18121 VDD.n2758 VDD.n51 9.3005
R18122 VDD.n2757 VDD.n52 9.3005
R18123 VDD.n60 VDD.n53 9.3005
R18124 VDD.n2751 VDD.n61 9.3005
R18125 VDD.n2750 VDD.n62 9.3005
R18126 VDD.n2749 VDD.n63 9.3005
R18127 VDD.n71 VDD.n64 9.3005
R18128 VDD.n2743 VDD.n72 9.3005
R18129 VDD.n2742 VDD.n73 9.3005
R18130 VDD.n2741 VDD.n74 9.3005
R18131 VDD.n81 VDD.n75 9.3005
R18132 VDD.n2735 VDD.n82 9.3005
R18133 VDD.n2734 VDD.n83 9.3005
R18134 VDD.n2733 VDD.n84 9.3005
R18135 VDD.n93 VDD.n85 9.3005
R18136 VDD.n2727 VDD.n2726 9.3005
R18137 VDD.n2774 VDD.n2773 9.3005
R18138 VDD.n212 VDD.n211 9.3005
R18139 VDD.n2570 VDD.n2569 9.3005
R18140 VDD.n2571 VDD.n210 9.3005
R18141 VDD.n2573 VDD.n2572 9.3005
R18142 VDD.n201 VDD.n200 9.3005
R18143 VDD.n2586 VDD.n2585 9.3005
R18144 VDD.n2587 VDD.n199 9.3005
R18145 VDD.n2589 VDD.n2588 9.3005
R18146 VDD.n189 VDD.n188 9.3005
R18147 VDD.n2602 VDD.n2601 9.3005
R18148 VDD.n2603 VDD.n187 9.3005
R18149 VDD.n2605 VDD.n2604 9.3005
R18150 VDD.n177 VDD.n176 9.3005
R18151 VDD.n2618 VDD.n2617 9.3005
R18152 VDD.n2619 VDD.n175 9.3005
R18153 VDD.n2621 VDD.n2620 9.3005
R18154 VDD.n165 VDD.n164 9.3005
R18155 VDD.n2634 VDD.n2633 9.3005
R18156 VDD.n2635 VDD.n163 9.3005
R18157 VDD.n2637 VDD.n2636 9.3005
R18158 VDD.n29 VDD.n27 9.3005
R18159 VDD.n2556 VDD.n2555 9.3005
R18160 VDD.n2506 VDD.n2505 9.3005
R18161 VDD.n2507 VDD.n260 9.3005
R18162 VDD.n259 VDD.n256 9.3005
R18163 VDD.n2513 VDD.n255 9.3005
R18164 VDD.n2514 VDD.n254 9.3005
R18165 VDD.n2515 VDD.n253 9.3005
R18166 VDD.n252 VDD.n250 9.3005
R18167 VDD.n2521 VDD.n249 9.3005
R18168 VDD.n2522 VDD.n246 9.3005
R18169 VDD.n2523 VDD.n245 9.3005
R18170 VDD.n244 VDD.n242 9.3005
R18171 VDD.n2529 VDD.n221 9.3005
R18172 VDD.n2530 VDD.n241 9.3005
R18173 VDD.n2531 VDD.n240 9.3005
R18174 VDD.n239 VDD.n237 9.3005
R18175 VDD.n2537 VDD.n236 9.3005
R18176 VDD.n2538 VDD.n235 9.3005
R18177 VDD.n2539 VDD.n232 9.3005
R18178 VDD.n231 VDD.n229 9.3005
R18179 VDD.n2544 VDD.n228 9.3005
R18180 VDD.n2545 VDD.n227 9.3005
R18181 VDD.n226 VDD.n224 9.3005
R18182 VDD.n2550 VDD.n223 9.3005
R18183 VDD.n2552 VDD.n2551 9.3005
R18184 VDD.n2504 VDD.n2503 9.3005
R18185 VDD.n1428 VDD.n1159 9.3005
R18186 VDD.n1430 VDD.n1429 9.3005
R18187 VDD.n1149 VDD.n1148 9.3005
R18188 VDD.n1443 VDD.n1442 9.3005
R18189 VDD.n1444 VDD.n1147 9.3005
R18190 VDD.n1446 VDD.n1445 9.3005
R18191 VDD.n1137 VDD.n1136 9.3005
R18192 VDD.n1460 VDD.n1459 9.3005
R18193 VDD.n1461 VDD.n1135 9.3005
R18194 VDD.n1463 VDD.n1462 9.3005
R18195 VDD.n1126 VDD.n1125 9.3005
R18196 VDD.n1476 VDD.n1475 9.3005
R18197 VDD.n1477 VDD.n1124 9.3005
R18198 VDD.n1479 VDD.n1478 9.3005
R18199 VDD.n1113 VDD.n1112 9.3005
R18200 VDD.n1493 VDD.n1492 9.3005
R18201 VDD.n1494 VDD.n1111 9.3005
R18202 VDD.n1496 VDD.n1495 9.3005
R18203 VDD.n1100 VDD.n1099 9.3005
R18204 VDD.n1512 VDD.n1511 9.3005
R18205 VDD.n1513 VDD.n1098 9.3005
R18206 VDD.n1515 VDD.n1514 9.3005
R18207 VDD.n1520 VDD.n1094 9.3005
R18208 VDD.n1522 VDD.n1521 9.3005
R18209 VDD.n1523 VDD.n1093 9.3005
R18210 VDD.n1527 VDD.n1526 9.3005
R18211 VDD.n1528 VDD.n1090 9.3005
R18212 VDD.n1532 VDD.n1529 9.3005
R18213 VDD.n1533 VDD.n1089 9.3005
R18214 VDD.n1537 VDD.n1536 9.3005
R18215 VDD.n1538 VDD.n1088 9.3005
R18216 VDD.n1540 VDD.n1539 9.3005
R18217 VDD.n1058 VDD.n1056 9.3005
R18218 VDD.n1573 VDD.n1572 9.3005
R18219 VDD.n1571 VDD.n1057 9.3005
R18220 VDD.n1570 VDD.n1569 9.3005
R18221 VDD.n1568 VDD.n1064 9.3005
R18222 VDD.n1567 VDD.n1566 9.3005
R18223 VDD.n1565 VDD.n1065 9.3005
R18224 VDD.n1564 VDD.n1563 9.3005
R18225 VDD.n1562 VDD.n1069 9.3005
R18226 VDD.n1561 VDD.n1560 9.3005
R18227 VDD.n1559 VDD.n1070 9.3005
R18228 VDD.n1558 VDD.n1557 9.3005
R18229 VDD.n1556 VDD.n1074 9.3005
R18230 VDD.n1555 VDD.n1554 9.3005
R18231 VDD.n1519 VDD.n1518 9.3005
R18232 VDD.n1327 VDD.n1224 9.3005
R18233 VDD.n1329 VDD.n1328 9.3005
R18234 VDD.n1215 VDD.n1214 9.3005
R18235 VDD.n1343 VDD.n1342 9.3005
R18236 VDD.n1344 VDD.n1213 9.3005
R18237 VDD.n1346 VDD.n1345 9.3005
R18238 VDD.n1203 VDD.n1202 9.3005
R18239 VDD.n1359 VDD.n1358 9.3005
R18240 VDD.n1360 VDD.n1201 9.3005
R18241 VDD.n1362 VDD.n1361 9.3005
R18242 VDD.n1191 VDD.n1190 9.3005
R18243 VDD.n1375 VDD.n1374 9.3005
R18244 VDD.n1376 VDD.n1189 9.3005
R18245 VDD.n1378 VDD.n1377 9.3005
R18246 VDD.n1179 VDD.n1178 9.3005
R18247 VDD.n1391 VDD.n1390 9.3005
R18248 VDD.n1392 VDD.n1177 9.3005
R18249 VDD.n1394 VDD.n1393 9.3005
R18250 VDD.n1167 VDD.n1166 9.3005
R18251 VDD.n1407 VDD.n1406 9.3005
R18252 VDD.n1408 VDD.n1165 9.3005
R18253 VDD.n1410 VDD.n1409 9.3005
R18254 VDD.n1154 VDD.n1153 9.3005
R18255 VDD.n1435 VDD.n1434 9.3005
R18256 VDD.n1436 VDD.n1152 9.3005
R18257 VDD.n1438 VDD.n1437 9.3005
R18258 VDD.n1143 VDD.n1142 9.3005
R18259 VDD.n1451 VDD.n1450 9.3005
R18260 VDD.n1452 VDD.n1141 9.3005
R18261 VDD.n1454 VDD.n1453 9.3005
R18262 VDD.n1132 VDD.n1131 9.3005
R18263 VDD.n1468 VDD.n1467 9.3005
R18264 VDD.n1469 VDD.n1130 9.3005
R18265 VDD.n1471 VDD.n1470 9.3005
R18266 VDD.n1120 VDD.n1119 9.3005
R18267 VDD.n1484 VDD.n1483 9.3005
R18268 VDD.n1485 VDD.n1117 9.3005
R18269 VDD.n1488 VDD.n1487 9.3005
R18270 VDD.n1486 VDD.n1118 9.3005
R18271 VDD.n1107 VDD.n1106 9.3005
R18272 VDD.n1502 VDD.n1501 9.3005
R18273 VDD.n1503 VDD.n1104 9.3005
R18274 VDD.n1506 VDD.n1505 9.3005
R18275 VDD.n1504 VDD.n1105 9.3005
R18276 VDD.n1326 VDD.n1325 9.3005
R18277 VDD.n1275 VDD.n1274 9.3005
R18278 VDD.n1276 VDD.n1265 9.3005
R18279 VDD.n1278 VDD.n1277 9.3005
R18280 VDD.n1279 VDD.n1259 9.3005
R18281 VDD.n1281 VDD.n1280 9.3005
R18282 VDD.n1282 VDD.n1257 9.3005
R18283 VDD.n1284 VDD.n1283 9.3005
R18284 VDD.n1258 VDD.n1255 9.3005
R18285 VDD.n1291 VDD.n1251 9.3005
R18286 VDD.n1293 VDD.n1292 9.3005
R18287 VDD.n1294 VDD.n1250 9.3005
R18288 VDD.n1296 VDD.n1295 9.3005
R18289 VDD.n1297 VDD.n1244 9.3005
R18290 VDD.n1299 VDD.n1298 9.3005
R18291 VDD.n1300 VDD.n1242 9.3005
R18292 VDD.n1302 VDD.n1301 9.3005
R18293 VDD.n1243 VDD.n1239 9.3005
R18294 VDD.n1310 VDD.n1240 9.3005
R18295 VDD.n1311 VDD.n1234 9.3005
R18296 VDD.n1313 VDD.n1312 9.3005
R18297 VDD.n1314 VDD.n1233 9.3005
R18298 VDD.n1316 VDD.n1315 9.3005
R18299 VDD.n1317 VDD.n1229 9.3005
R18300 VDD.n1319 VDD.n1318 9.3005
R18301 VDD.n1270 VDD.n1225 9.3005
R18302 VDD.n1220 VDD.n1219 9.3005
R18303 VDD.n1335 VDD.n1334 9.3005
R18304 VDD.n1336 VDD.n1218 9.3005
R18305 VDD.n1338 VDD.n1337 9.3005
R18306 VDD.n1209 VDD.n1208 9.3005
R18307 VDD.n1351 VDD.n1350 9.3005
R18308 VDD.n1352 VDD.n1207 9.3005
R18309 VDD.n1354 VDD.n1353 9.3005
R18310 VDD.n1197 VDD.n1196 9.3005
R18311 VDD.n1367 VDD.n1366 9.3005
R18312 VDD.n1368 VDD.n1195 9.3005
R18313 VDD.n1370 VDD.n1369 9.3005
R18314 VDD.n1185 VDD.n1184 9.3005
R18315 VDD.n1383 VDD.n1382 9.3005
R18316 VDD.n1384 VDD.n1183 9.3005
R18317 VDD.n1386 VDD.n1385 9.3005
R18318 VDD.n1173 VDD.n1172 9.3005
R18319 VDD.n1399 VDD.n1398 9.3005
R18320 VDD.n1400 VDD.n1171 9.3005
R18321 VDD.n1402 VDD.n1401 9.3005
R18322 VDD.n1161 VDD.n1160 9.3005
R18323 VDD.n1321 VDD.n1320 9.3005
R18324 VDD.n1427 VDD.n1414 9.3005
R18325 VDD.n1634 VDD.t2 8.62119
R18326 VDD.t33 VDD.n330 8.62119
R18327 VDD.n15 VDD.n14 8.20441
R18328 VDD.n2775 VDD.n2774 8.15725
R18329 VDD.n1427 VDD.n1426 8.15725
R18330 VDD.n1292 VDD.n1291 7.17626
R18331 VDD.n2523 VDD.n2522 7.17626
R18332 VDD.n2699 VDD.n2698 7.17626
R18333 VDD.n1570 VDD.n1064 7.17626
R18334 VDD.n2060 VDD.n2056 6.86879
R18335 VDD.n2453 VDD.n2452 6.86879
R18336 VDD.n2491 VDD.n272 6.86879
R18337 VDD.n1903 VDD.n1902 6.86879
R18338 VDD.n1858 VDD.n545 6.86879
R18339 VDD.n824 VDD.n823 6.86879
R18340 VDD.n1804 VDD.n1802 6.86879
R18341 VDD.n1042 VDD.n1041 6.86879
R18342 VDD.n22 VDD.n18 6.70309
R18343 VDD.n1421 VDD.n1417 6.70309
R18344 VDD.n2775 VDD.n26 6.38454
R18345 VDD.n1426 VDD.n1425 6.38454
R18346 VDD.n11 VDD.n9 6.15136
R18347 VDD.n4 VDD.n2 6.15136
R18348 VDD.t2 VDD.n716 6.03498
R18349 VDD.n2380 VDD.t33 6.03498
R18350 VDD.t114 VDD.n1169 5.60395
R18351 VDD.n1157 VDD.t106 5.60395
R18352 VDD.t122 VDD.n161 5.60395
R18353 VDD.t125 VDD.n37 5.60395
R18354 VDD.n2464 VDD.n222 5.30782
R18355 VDD.n290 VDD.n222 5.30782
R18356 VDD.n2501 VDD.n264 5.30782
R18357 VDD.n2501 VDD.n2500 5.30782
R18358 VDD.n1576 VDD.n1575 5.30782
R18359 VDD.n1575 VDD.n772 5.30782
R18360 VDD.n1054 VDD.n774 5.30782
R18361 VDD.n1054 VDD.n1053 5.30782
R18362 VDD.n13 VDD.n11 4.90567
R18363 VDD.n6 VDD.n4 4.90567
R18364 VDD.n26 VDD.n25 4.88412
R18365 VDD.n22 VDD.n21 4.88412
R18366 VDD.n1425 VDD.n1424 4.88412
R18367 VDD.n1421 VDD.n1420 4.88412
R18368 VDD.n1273 VDD.n1270 4.84898
R18369 VDD.n2503 VDD.n263 4.84898
R18370 VDD.n2680 VDD.n138 4.84898
R18371 VDD.n1554 VDD.n1078 4.84898
R18372 VDD.n1372 VDD.t117 4.74188
R18373 VDD.n1465 VDD.t128 4.74188
R18374 VDD.n675 VDD.t13 4.74188
R18375 VDD.n2332 VDD.t22 4.74188
R18376 VDD.n2607 VDD.t108 4.74188
R18377 VDD.t110 VDD.n2753 4.74188
R18378 VDD.n221 VDD.n217 4.25965
R18379 VDD.n2554 VDD.n221 4.04623
R18380 VDD.n14 VDD.n13 3.76491
R18381 VDD.n14 VDD.n6 3.76491
R18382 VDD.n2169 VDD.n2060 3.74684
R18383 VDD.n2452 VDD.n2451 3.74684
R18384 VDD.n274 VDD.n272 3.74684
R18385 VDD.n1938 VDD.n1902 3.74684
R18386 VDD.n1855 VDD.n545 3.74684
R18387 VDD.n823 VDD.n808 3.74684
R18388 VDD.n1802 VDD.n534 3.74684
R18389 VDD.n1041 VDD.n1040 3.74684
R18390 VDD.n1574 VDD.n1573 3.70782
R18391 VDD.n1573 VDD.n1055 3.70782
R18392 VDD.n937 VDD.t20 3.01774
R18393 VDD.n2230 VDD.t24 3.01774
R18394 VDD.n25 VDD.n24 2.81084
R18395 VDD.n21 VDD.n20 2.81084
R18396 VDD.n18 VDD.n17 2.81084
R18397 VDD.n1424 VDD.n1423 2.81084
R18398 VDD.n1420 VDD.n1419 2.81084
R18399 VDD.n1417 VDD.n1416 2.81084
R18400 VDD.n742 VDD.t43 2.80222
R18401 VDD.n1790 VDD.t50 2.80222
R18402 VDD.n494 VDD.t54 2.80222
R18403 VDD.n2398 VDD.t94 2.80222
R18404 VDD.n1426 VDD.n15 2.29206
R18405 VDD VDD.n2775 2.28423
R18406 VDD.n682 VDD.t12 1.94016
R18407 VDD.n1730 VDD.t17 1.94016
R18408 VDD.n434 VDD.t28 1.94016
R18409 VDD.n2338 VDD.t35 1.94016
R18410 VDD.n26 VDD.n22 1.81947
R18411 VDD.n1425 VDD.n1421 1.81947
R18412 VDD.n1274 VDD.n1273 1.74595
R18413 VDD.n2506 VDD.n263 1.74595
R18414 VDD.n138 VDD.n134 1.74595
R18415 VDD.n1078 VDD.n1074 1.74595
R18416 VDD.n1736 VDD.t8 0.862569
R18417 VDD.t26 VDD.n431 0.862569
R18418 VDD.n1555 VDD.n1075 0.60111
R18419 VDD.n2679 VDD.n2678 0.491354
R18420 VDD.n2726 VDD.n2725 0.491354
R18421 VDD.n1326 VDD.n1225 0.491354
R18422 VDD.n1320 VDD.n1319 0.491354
R18423 VDD.n2555 VDD.n2554 0.404463
R18424 VDD.n1514 VDD.n773 0.404463
R18425 VDD.n1519 VDD.n773 0.387695
R18426 VDD.n2552 VDD.n223 0.305378
R18427 VDD.n226 VDD.n223 0.305378
R18428 VDD.n227 VDD.n226 0.305378
R18429 VDD.n228 VDD.n227 0.305378
R18430 VDD.n231 VDD.n228 0.305378
R18431 VDD.n232 VDD.n231 0.305378
R18432 VDD.n235 VDD.n232 0.305378
R18433 VDD.n236 VDD.n235 0.305378
R18434 VDD.n239 VDD.n236 0.305378
R18435 VDD.n240 VDD.n239 0.305378
R18436 VDD.n241 VDD.n240 0.305378
R18437 VDD.n241 VDD.n221 0.305378
R18438 VDD.n244 VDD.n221 0.305378
R18439 VDD.n245 VDD.n244 0.305378
R18440 VDD.n246 VDD.n245 0.305378
R18441 VDD.n249 VDD.n246 0.305378
R18442 VDD.n252 VDD.n249 0.305378
R18443 VDD.n253 VDD.n252 0.305378
R18444 VDD.n254 VDD.n253 0.305378
R18445 VDD.n255 VDD.n254 0.305378
R18446 VDD.n259 VDD.n255 0.305378
R18447 VDD.n260 VDD.n259 0.305378
R18448 VDD.n2505 VDD.n260 0.305378
R18449 VDD.n2505 VDD.n2504 0.305378
R18450 VDD.n1520 VDD.n1519 0.305378
R18451 VDD.n1521 VDD.n1520 0.305378
R18452 VDD.n1521 VDD.n1093 0.305378
R18453 VDD.n1527 VDD.n1093 0.305378
R18454 VDD.n1528 VDD.n1527 0.305378
R18455 VDD.n1529 VDD.n1528 0.305378
R18456 VDD.n1529 VDD.n1089 0.305378
R18457 VDD.n1537 VDD.n1089 0.305378
R18458 VDD.n1538 VDD.n1537 0.305378
R18459 VDD.n1539 VDD.n1538 0.305378
R18460 VDD.n1539 VDD.n1056 0.305378
R18461 VDD.n1573 VDD.n1056 0.305378
R18462 VDD.n1573 VDD.n1057 0.305378
R18463 VDD.n1569 VDD.n1057 0.305378
R18464 VDD.n1569 VDD.n1568 0.305378
R18465 VDD.n1568 VDD.n1567 0.305378
R18466 VDD.n1567 VDD.n1065 0.305378
R18467 VDD.n1563 VDD.n1065 0.305378
R18468 VDD.n1563 VDD.n1562 0.305378
R18469 VDD.n1562 VDD.n1561 0.305378
R18470 VDD.n1561 VDD.n1070 0.305378
R18471 VDD.n1557 VDD.n1070 0.305378
R18472 VDD.n1557 VDD.n1556 0.305378
R18473 VDD.n1556 VDD.n1555 0.305378
R18474 VDD.n2561 VDD.n217 0.191049
R18475 VDD.n1504 VDD.n1075 0.191049
R18476 VDD.n2562 VDD.n2561 0.152939
R18477 VDD.n2563 VDD.n2562 0.152939
R18478 VDD.n2563 VDD.n206 0.152939
R18479 VDD.n2578 VDD.n206 0.152939
R18480 VDD.n2579 VDD.n2578 0.152939
R18481 VDD.n2580 VDD.n2579 0.152939
R18482 VDD.n2580 VDD.n194 0.152939
R18483 VDD.n2594 VDD.n194 0.152939
R18484 VDD.n2595 VDD.n2594 0.152939
R18485 VDD.n2596 VDD.n2595 0.152939
R18486 VDD.n2596 VDD.n182 0.152939
R18487 VDD.n2610 VDD.n182 0.152939
R18488 VDD.n2611 VDD.n2610 0.152939
R18489 VDD.n2612 VDD.n2611 0.152939
R18490 VDD.n2612 VDD.n170 0.152939
R18491 VDD.n2626 VDD.n170 0.152939
R18492 VDD.n2627 VDD.n2626 0.152939
R18493 VDD.n2628 VDD.n2627 0.152939
R18494 VDD.n2628 VDD.n157 0.152939
R18495 VDD.n2642 VDD.n157 0.152939
R18496 VDD.n2643 VDD.n2642 0.152939
R18497 VDD.n2644 VDD.n2643 0.152939
R18498 VDD.n2644 VDD.n155 0.152939
R18499 VDD.n2648 VDD.n155 0.152939
R18500 VDD.n2649 VDD.n2648 0.152939
R18501 VDD.n2650 VDD.n2649 0.152939
R18502 VDD.n2650 VDD.n152 0.152939
R18503 VDD.n2654 VDD.n152 0.152939
R18504 VDD.n2655 VDD.n2654 0.152939
R18505 VDD.n2656 VDD.n2655 0.152939
R18506 VDD.n2656 VDD.n149 0.152939
R18507 VDD.n2660 VDD.n149 0.152939
R18508 VDD.n2661 VDD.n2660 0.152939
R18509 VDD.n2662 VDD.n2661 0.152939
R18510 VDD.n2662 VDD.n146 0.152939
R18511 VDD.n2666 VDD.n146 0.152939
R18512 VDD.n2667 VDD.n2666 0.152939
R18513 VDD.n2668 VDD.n2667 0.152939
R18514 VDD.n2668 VDD.n143 0.152939
R18515 VDD.n2672 VDD.n143 0.152939
R18516 VDD.n2673 VDD.n2672 0.152939
R18517 VDD.n2674 VDD.n2673 0.152939
R18518 VDD.n2674 VDD.n140 0.152939
R18519 VDD.n2678 VDD.n140 0.152939
R18520 VDD.n2725 VDD.n94 0.152939
R18521 VDD.n96 VDD.n94 0.152939
R18522 VDD.n100 VDD.n96 0.152939
R18523 VDD.n101 VDD.n100 0.152939
R18524 VDD.n102 VDD.n101 0.152939
R18525 VDD.n2714 VDD.n102 0.152939
R18526 VDD.n2714 VDD.n2713 0.152939
R18527 VDD.n2713 VDD.n2712 0.152939
R18528 VDD.n2712 VDD.n108 0.152939
R18529 VDD.n113 VDD.n108 0.152939
R18530 VDD.n114 VDD.n113 0.152939
R18531 VDD.n115 VDD.n114 0.152939
R18532 VDD.n119 VDD.n115 0.152939
R18533 VDD.n120 VDD.n119 0.152939
R18534 VDD.n2697 VDD.n120 0.152939
R18535 VDD.n2697 VDD.n2696 0.152939
R18536 VDD.n2696 VDD.n2695 0.152939
R18537 VDD.n2695 VDD.n124 0.152939
R18538 VDD.n130 VDD.n124 0.152939
R18539 VDD.n131 VDD.n130 0.152939
R18540 VDD.n132 VDD.n131 0.152939
R18541 VDD.n133 VDD.n132 0.152939
R18542 VDD.n139 VDD.n133 0.152939
R18543 VDD.n2679 VDD.n139 0.152939
R18544 VDD.n39 VDD.n28 0.152939
R18545 VDD.n40 VDD.n39 0.152939
R18546 VDD.n41 VDD.n40 0.152939
R18547 VDD.n49 VDD.n41 0.152939
R18548 VDD.n50 VDD.n49 0.152939
R18549 VDD.n51 VDD.n50 0.152939
R18550 VDD.n52 VDD.n51 0.152939
R18551 VDD.n60 VDD.n52 0.152939
R18552 VDD.n61 VDD.n60 0.152939
R18553 VDD.n62 VDD.n61 0.152939
R18554 VDD.n63 VDD.n62 0.152939
R18555 VDD.n71 VDD.n63 0.152939
R18556 VDD.n72 VDD.n71 0.152939
R18557 VDD.n73 VDD.n72 0.152939
R18558 VDD.n74 VDD.n73 0.152939
R18559 VDD.n81 VDD.n74 0.152939
R18560 VDD.n82 VDD.n81 0.152939
R18561 VDD.n83 VDD.n82 0.152939
R18562 VDD.n84 VDD.n83 0.152939
R18563 VDD.n93 VDD.n84 0.152939
R18564 VDD.n2726 VDD.n93 0.152939
R18565 VDD.n2555 VDD.n211 0.152939
R18566 VDD.n2570 VDD.n211 0.152939
R18567 VDD.n2571 VDD.n2570 0.152939
R18568 VDD.n2572 VDD.n2571 0.152939
R18569 VDD.n2572 VDD.n200 0.152939
R18570 VDD.n2586 VDD.n200 0.152939
R18571 VDD.n2587 VDD.n2586 0.152939
R18572 VDD.n2588 VDD.n2587 0.152939
R18573 VDD.n2588 VDD.n188 0.152939
R18574 VDD.n2602 VDD.n188 0.152939
R18575 VDD.n2603 VDD.n2602 0.152939
R18576 VDD.n2604 VDD.n2603 0.152939
R18577 VDD.n2604 VDD.n176 0.152939
R18578 VDD.n2618 VDD.n176 0.152939
R18579 VDD.n2619 VDD.n2618 0.152939
R18580 VDD.n2620 VDD.n2619 0.152939
R18581 VDD.n2620 VDD.n164 0.152939
R18582 VDD.n2634 VDD.n164 0.152939
R18583 VDD.n2635 VDD.n2634 0.152939
R18584 VDD.n2636 VDD.n2635 0.152939
R18585 VDD.n2636 VDD.n27 0.152939
R18586 VDD.n1429 VDD.n1428 0.152939
R18587 VDD.n1429 VDD.n1148 0.152939
R18588 VDD.n1443 VDD.n1148 0.152939
R18589 VDD.n1444 VDD.n1443 0.152939
R18590 VDD.n1445 VDD.n1444 0.152939
R18591 VDD.n1445 VDD.n1136 0.152939
R18592 VDD.n1460 VDD.n1136 0.152939
R18593 VDD.n1461 VDD.n1460 0.152939
R18594 VDD.n1462 VDD.n1461 0.152939
R18595 VDD.n1462 VDD.n1125 0.152939
R18596 VDD.n1476 VDD.n1125 0.152939
R18597 VDD.n1477 VDD.n1476 0.152939
R18598 VDD.n1478 VDD.n1477 0.152939
R18599 VDD.n1478 VDD.n1112 0.152939
R18600 VDD.n1493 VDD.n1112 0.152939
R18601 VDD.n1494 VDD.n1493 0.152939
R18602 VDD.n1495 VDD.n1494 0.152939
R18603 VDD.n1495 VDD.n1099 0.152939
R18604 VDD.n1512 VDD.n1099 0.152939
R18605 VDD.n1513 VDD.n1512 0.152939
R18606 VDD.n1514 VDD.n1513 0.152939
R18607 VDD.n1327 VDD.n1326 0.152939
R18608 VDD.n1328 VDD.n1327 0.152939
R18609 VDD.n1328 VDD.n1214 0.152939
R18610 VDD.n1343 VDD.n1214 0.152939
R18611 VDD.n1344 VDD.n1343 0.152939
R18612 VDD.n1345 VDD.n1344 0.152939
R18613 VDD.n1345 VDD.n1202 0.152939
R18614 VDD.n1359 VDD.n1202 0.152939
R18615 VDD.n1360 VDD.n1359 0.152939
R18616 VDD.n1361 VDD.n1360 0.152939
R18617 VDD.n1361 VDD.n1190 0.152939
R18618 VDD.n1375 VDD.n1190 0.152939
R18619 VDD.n1376 VDD.n1375 0.152939
R18620 VDD.n1377 VDD.n1376 0.152939
R18621 VDD.n1377 VDD.n1178 0.152939
R18622 VDD.n1391 VDD.n1178 0.152939
R18623 VDD.n1392 VDD.n1391 0.152939
R18624 VDD.n1393 VDD.n1392 0.152939
R18625 VDD.n1393 VDD.n1166 0.152939
R18626 VDD.n1407 VDD.n1166 0.152939
R18627 VDD.n1408 VDD.n1407 0.152939
R18628 VDD.n1409 VDD.n1408 0.152939
R18629 VDD.n1409 VDD.n1153 0.152939
R18630 VDD.n1435 VDD.n1153 0.152939
R18631 VDD.n1436 VDD.n1435 0.152939
R18632 VDD.n1437 VDD.n1436 0.152939
R18633 VDD.n1437 VDD.n1142 0.152939
R18634 VDD.n1451 VDD.n1142 0.152939
R18635 VDD.n1452 VDD.n1451 0.152939
R18636 VDD.n1453 VDD.n1452 0.152939
R18637 VDD.n1453 VDD.n1131 0.152939
R18638 VDD.n1468 VDD.n1131 0.152939
R18639 VDD.n1469 VDD.n1468 0.152939
R18640 VDD.n1470 VDD.n1469 0.152939
R18641 VDD.n1470 VDD.n1119 0.152939
R18642 VDD.n1484 VDD.n1119 0.152939
R18643 VDD.n1485 VDD.n1484 0.152939
R18644 VDD.n1487 VDD.n1485 0.152939
R18645 VDD.n1487 VDD.n1486 0.152939
R18646 VDD.n1486 VDD.n1106 0.152939
R18647 VDD.n1502 VDD.n1106 0.152939
R18648 VDD.n1503 VDD.n1502 0.152939
R18649 VDD.n1505 VDD.n1503 0.152939
R18650 VDD.n1505 VDD.n1504 0.152939
R18651 VDD.n1319 VDD.n1229 0.152939
R18652 VDD.n1315 VDD.n1229 0.152939
R18653 VDD.n1315 VDD.n1314 0.152939
R18654 VDD.n1314 VDD.n1313 0.152939
R18655 VDD.n1313 VDD.n1234 0.152939
R18656 VDD.n1240 VDD.n1234 0.152939
R18657 VDD.n1243 VDD.n1240 0.152939
R18658 VDD.n1301 VDD.n1243 0.152939
R18659 VDD.n1301 VDD.n1300 0.152939
R18660 VDD.n1300 VDD.n1299 0.152939
R18661 VDD.n1299 VDD.n1244 0.152939
R18662 VDD.n1295 VDD.n1244 0.152939
R18663 VDD.n1295 VDD.n1294 0.152939
R18664 VDD.n1294 VDD.n1293 0.152939
R18665 VDD.n1293 VDD.n1251 0.152939
R18666 VDD.n1258 VDD.n1251 0.152939
R18667 VDD.n1283 VDD.n1258 0.152939
R18668 VDD.n1283 VDD.n1282 0.152939
R18669 VDD.n1282 VDD.n1281 0.152939
R18670 VDD.n1281 VDD.n1259 0.152939
R18671 VDD.n1277 VDD.n1259 0.152939
R18672 VDD.n1277 VDD.n1276 0.152939
R18673 VDD.n1276 VDD.n1275 0.152939
R18674 VDD.n1275 VDD.n1225 0.152939
R18675 VDD.n1320 VDD.n1219 0.152939
R18676 VDD.n1335 VDD.n1219 0.152939
R18677 VDD.n1336 VDD.n1335 0.152939
R18678 VDD.n1337 VDD.n1336 0.152939
R18679 VDD.n1337 VDD.n1208 0.152939
R18680 VDD.n1351 VDD.n1208 0.152939
R18681 VDD.n1352 VDD.n1351 0.152939
R18682 VDD.n1353 VDD.n1352 0.152939
R18683 VDD.n1353 VDD.n1196 0.152939
R18684 VDD.n1367 VDD.n1196 0.152939
R18685 VDD.n1368 VDD.n1367 0.152939
R18686 VDD.n1369 VDD.n1368 0.152939
R18687 VDD.n1369 VDD.n1184 0.152939
R18688 VDD.n1383 VDD.n1184 0.152939
R18689 VDD.n1384 VDD.n1383 0.152939
R18690 VDD.n1385 VDD.n1384 0.152939
R18691 VDD.n1385 VDD.n1172 0.152939
R18692 VDD.n1399 VDD.n1172 0.152939
R18693 VDD.n1400 VDD.n1399 0.152939
R18694 VDD.n1401 VDD.n1400 0.152939
R18695 VDD.n1401 VDD.n1160 0.152939
R18696 VDD.n2774 VDD.n28 0.145814
R18697 VDD.n2774 VDD.n27 0.145814
R18698 VDD.n1428 VDD.n1427 0.145814
R18699 VDD.n1427 VDD.n1160 0.145814
R18700 VDD.n1075 VDD.n1055 0.0649893
R18701 VDD.n2502 VDD.n217 0.0646768
R18702 VDD.n2553 VDD.n2552 0.0492805
R18703 VDD.n2504 VDD.n2502 0.0492805
R18704 VDD VDD.n15 0.00833333
R18705 VDD.n1574 VDD.n773 0.0070625
R18706 VDD.n2554 VDD.n2553 0.00675
R18707 VP.n2 VP.t5 243.97
R18708 VP.n7 VP.t2 243.255
R18709 VP.n6 VP.n5 223.454
R18710 VP.n4 VP.n3 223.454
R18711 VP.n2 VP.n1 223.454
R18712 VP.n0 VP.t9 78.253
R18713 VP.n0 VP.t8 59.6292
R18714 VP.n5 VP.t0 19.8005
R18715 VP.n5 VP.t6 19.8005
R18716 VP.n3 VP.t7 19.8005
R18717 VP.n3 VP.t4 19.8005
R18718 VP.n1 VP.t1 19.8005
R18719 VP.n1 VP.t3 19.8005
R18720 VP VP.n8 15.4161
R18721 VP.n8 VP.n7 4.80222
R18722 VP.n8 VP.n0 0.972091
R18723 VP.n4 VP.n2 0.716017
R18724 VP.n6 VP.n4 0.716017
R18725 VP.n7 VP.n6 0.716017
R18726 VN.n2 VN.t0 243.97
R18727 VN.n7 VN.t5 243.255
R18728 VN.n2 VN.n1 223.454
R18729 VN.n4 VN.n3 223.454
R18730 VN.n6 VN.n5 223.454
R18731 VN.n0 VN.t9 78.0383
R18732 VN.n0 VN.t8 59.412
R18733 VN.n1 VN.t2 19.8005
R18734 VN.n1 VN.t4 19.8005
R18735 VN.n3 VN.t7 19.8005
R18736 VN.n3 VN.t6 19.8005
R18737 VN.n5 VN.t1 19.8005
R18738 VN.n5 VN.t3 19.8005
R18739 VN VN.n8 18.137
R18740 VN.n8 VN.n7 5.04791
R18741 VN.n8 VN.n0 1.188
R18742 VN.n7 VN.n6 0.716017
R18743 VN.n6 VN.n4 0.716017
R18744 VN.n4 VN.n2 0.716017
R18745 a_n1140_n227.n1 a_n1140_n227.t3 83.7273
R18746 a_n1140_n227.n1 a_n1140_n227.t1 83.7273
R18747 a_n1140_n227.n2 a_n1140_n227.t4 83.7273
R18748 a_n1140_n227.t2 a_n1140_n227.n2 83.7273
R18749 a_n1140_n227.n0 a_n1140_n227.n1 6.61795
R18750 a_n1140_n227.n2 a_n1140_n227.n0 4.86452
R18751 a_n1140_n227.t0 a_n1140_n227.n0 193.358
R18752 DIFFPAIR_BIAS.n0 DIFFPAIR_BIAS.t1 129.107
R18753 DIFFPAIR_BIAS.n1 DIFFPAIR_BIAS.t2 91.3632
R18754 DIFFPAIR_BIAS.n0 DIFFPAIR_BIAS.t0 69.4984
R18755 DIFFPAIR_BIAS.n1 DIFFPAIR_BIAS.n0 4.43723
R18756 DIFFPAIR_BIAS DIFFPAIR_BIAS.n1 2.19744
R18757 a_n10357_8879.n34 a_n10357_8879.n1 498.942
R18758 a_n10357_8879.n39 a_n10357_8879.n3 498.942
R18759 a_n10357_8879.n41 a_n10357_8879.n5 498.942
R18760 a_n10357_8879.n29 a_n10357_8879.n7 498.942
R18761 a_n10357_8879.n0 a_n10357_8879.n1 8.87206
R18762 a_n10357_8879.n34 a_n10357_8879.n10 585
R18763 a_n10357_8879.n18 a_n10357_8879.n17 585
R18764 a_n10357_8879.n2 a_n10357_8879.n3 8.87206
R18765 a_n10357_8879.n39 a_n10357_8879.n12 585
R18766 a_n10357_8879.n21 a_n10357_8879.n20 585
R18767 a_n10357_8879.n4 a_n10357_8879.n5 8.87206
R18768 a_n10357_8879.n41 a_n10357_8879.n14 585
R18769 a_n10357_8879.n24 a_n10357_8879.n23 585
R18770 a_n10357_8879.n6 a_n10357_8879.n7 8.87206
R18771 a_n10357_8879.n29 a_n10357_8879.n16 585
R18772 a_n10357_8879.n27 a_n10357_8879.n26 585
R18773 a_n10357_8879.n34 a_n10357_8879.n17 171.744
R18774 a_n10357_8879.n39 a_n10357_8879.n20 171.744
R18775 a_n10357_8879.n41 a_n10357_8879.n23 171.744
R18776 a_n10357_8879.n29 a_n10357_8879.n26 171.744
R18777 a_n10357_8879.n33 a_n10357_8879.n32 169.725
R18778 a_n10357_8879.n33 a_n10357_8879.n31 158.649
R18779 a_n10357_8879.n38 a_n10357_8879.n37 115.632
R18780 a_n10357_8879.n44 a_n10357_8879.n43 115.632
R18781 a_n10357_8879.t7 a_n10357_8879.n17 85.8723
R18782 a_n10357_8879.t6 a_n10357_8879.n20 85.8723
R18783 a_n10357_8879.t11 a_n10357_8879.n23 85.8723
R18784 a_n10357_8879.t9 a_n10357_8879.n26 85.8723
R18785 a_n10357_8879.n43 a_n10357_8879.n30 41.5511
R18786 a_n10357_8879.n36 a_n10357_8879.n35 36.646
R18787 a_n10357_8879.n8 a_n10357_8879.n40 36.646
R18788 a_n10357_8879.n8 a_n10357_8879.n42 36.646
R18789 a_n10357_8879.n19 a_n10357_8879.n18 5.21215
R18790 a_n10357_8879.n22 a_n10357_8879.n21 5.21215
R18791 a_n10357_8879.n25 a_n10357_8879.n24 5.21215
R18792 a_n10357_8879.n28 a_n10357_8879.n27 5.21215
R18793 a_n10357_8879.n10 a_n10357_8879.n18 12.8005
R18794 a_n10357_8879.n12 a_n10357_8879.n21 12.8005
R18795 a_n10357_8879.n14 a_n10357_8879.n24 12.8005
R18796 a_n10357_8879.n16 a_n10357_8879.n27 12.8005
R18797 a_n10357_8879.n37 a_n10357_8879.t4 9.70349
R18798 a_n10357_8879.n37 a_n10357_8879.t5 9.70349
R18799 a_n10357_8879.n31 a_n10357_8879.t2 9.70349
R18800 a_n10357_8879.n31 a_n10357_8879.t3 9.70349
R18801 a_n10357_8879.n32 a_n10357_8879.t0 9.70349
R18802 a_n10357_8879.n32 a_n10357_8879.t1 9.70349
R18803 a_n10357_8879.t10 a_n10357_8879.n44 9.70349
R18804 a_n10357_8879.n44 a_n10357_8879.t8 9.70349
R18805 a_n10357_8879.n28 a_n10357_8879.n15 1.35994
R18806 a_n10357_8879.n35 a_n10357_8879.n9 9.45567
R18807 a_n10357_8879.n40 a_n10357_8879.n11 9.45567
R18808 a_n10357_8879.n42 a_n10357_8879.n13 9.45567
R18809 a_n10357_8879.n30 a_n10357_8879.n15 9.45567
R18810 a_n10357_8879.n36 a_n10357_8879.n33 7.93369
R18811 a_n10357_8879.n8 a_n10357_8879.n38 4.90567
R18812 a_n10357_8879.n38 a_n10357_8879.n36 4.90567
R18813 a_n10357_8879.n19 a_n10357_8879.t7 339.173
R18814 a_n10357_8879.n22 a_n10357_8879.t6 339.173
R18815 a_n10357_8879.n25 a_n10357_8879.t11 339.173
R18816 a_n10357_8879.n28 a_n10357_8879.t9 339.173
R18817 a_n10357_8879.n9 a_n10357_8879.n0 3.48794
R18818 a_n10357_8879.n11 a_n10357_8879.n2 3.48794
R18819 a_n10357_8879.n13 a_n10357_8879.n4 3.48794
R18820 a_n10357_8879.n15 a_n10357_8879.n6 3.48794
R18821 a_n10357_8879.n16 a_n10357_8879.n6 3.73143
R18822 a_n10357_8879.n14 a_n10357_8879.n4 3.73143
R18823 a_n10357_8879.n12 a_n10357_8879.n2 3.73143
R18824 a_n10357_8879.n10 a_n10357_8879.n0 3.73143
R18825 a_n10357_8879.n43 a_n10357_8879.n8 6.15136
R18826 a_n10357_8879.n19 a_n10357_8879.n9 1.35994
R18827 a_n10357_8879.n22 a_n10357_8879.n11 1.35994
R18828 a_n10357_8879.n25 a_n10357_8879.n13 1.35994
R18829 a_n10357_8879.n35 a_n10357_8879.n1 9.00755
R18830 a_n10357_8879.n40 a_n10357_8879.n3 9.00755
R18831 a_n10357_8879.n42 a_n10357_8879.n5 9.00755
R18832 a_n10357_8879.n30 a_n10357_8879.n7 9.00755
C0 CS_BIAS VP 0.417694f
C1 VOUT VN 0.980676f
C2 CS_BIAS VN 0.428985f
C3 a_n819_n2194# VP 7.52e-19
C4 VP VN 10.512799f
C5 a_n819_n2194# VN 3.29e-19
C6 a_n11713_8879# VDD 1.68006f
C7 VP DIFFPAIR_BIAS 0.00716f
C8 a_n819_n2194# DIFFPAIR_BIAS 1.33318f
C9 VN DIFFPAIR_BIAS 0.010672f
C10 a_53_n2194# VP 8.59e-19
C11 VDD VOUT 26.3811f
C12 a_n819_n2194# a_53_n2194# 0.103039f
C13 a_53_n2194# VN 6.03e-19
C14 a_10485_8879# VDD 1.67952f
C15 VOUT CS_BIAS 35.456398f
C16 a_53_n2194# DIFFPAIR_BIAS 0.989992f
C17 VDD VN 0.106779f
C18 VOUT VP 4.68998f
C19 DIFFPAIR_BIAS GND 9.54093f
C20 VN GND 29.849329f
C21 VP GND 28.9007f
C22 CS_BIAS GND 0.138375p
C23 VOUT GND 80.3872f
C24 VDD GND 0.479968p
C25 a_53_n2194# GND 0.690734f
C26 a_n819_n2194# GND 1.04919f
C27 a_10485_8879# GND 0.677986f
C28 a_n11713_8879# GND 0.677986f
C29 a_n10357_8879.n0 GND 0.025792f
C30 a_n10357_8879.n1 GND 0.081937f
C31 a_n10357_8879.n2 GND 0.025792f
C32 a_n10357_8879.n3 GND 0.081937f
C33 a_n10357_8879.n4 GND 0.025792f
C34 a_n10357_8879.n5 GND 0.081937f
C35 a_n10357_8879.n6 GND 0.025792f
C36 a_n10357_8879.n7 GND 0.081937f
C37 a_n10357_8879.n8 GND 1.77328f
C38 a_n10357_8879.n9 GND 0.60694f
C39 a_n10357_8879.n10 GND 0.047043f
C40 a_n10357_8879.n11 GND 0.60694f
C41 a_n10357_8879.n12 GND 0.047043f
C42 a_n10357_8879.n13 GND 0.60694f
C43 a_n10357_8879.n14 GND 0.047043f
C44 a_n10357_8879.n15 GND 0.60694f
C45 a_n10357_8879.n16 GND 0.047043f
C46 a_n10357_8879.n17 GND 0.040506f
C47 a_n10357_8879.n18 GND 0.056192f
C48 a_n10357_8879.n19 GND 0.158184f
C49 a_n10357_8879.n20 GND 0.040506f
C50 a_n10357_8879.n21 GND 0.056192f
C51 a_n10357_8879.n22 GND 0.158184f
C52 a_n10357_8879.n23 GND 0.040506f
C53 a_n10357_8879.n24 GND 0.056192f
C54 a_n10357_8879.n25 GND 0.158184f
C55 a_n10357_8879.n26 GND 0.040506f
C56 a_n10357_8879.n27 GND 0.056192f
C57 a_n10357_8879.n28 GND 0.158184f
C58 a_n10357_8879.t9 GND 0.124293f
C59 a_n10357_8879.n29 GND 0.14217f
C60 a_n10357_8879.n30 GND 0.188098f
C61 a_n10357_8879.t2 GND 0.112567f
C62 a_n10357_8879.t3 GND 0.112567f
C63 a_n10357_8879.n31 GND 1.38835f
C64 a_n10357_8879.t0 GND 0.112567f
C65 a_n10357_8879.t1 GND 0.112567f
C66 a_n10357_8879.n32 GND 2.66378f
C67 a_n10357_8879.n33 GND 18.5849f
C68 a_n10357_8879.t7 GND 0.124293f
C69 a_n10357_8879.n34 GND 0.14217f
C70 a_n10357_8879.n35 GND 0.101555f
C71 a_n10357_8879.n36 GND 1.48627f
C72 a_n10357_8879.t4 GND 0.112567f
C73 a_n10357_8879.t5 GND 0.112567f
C74 a_n10357_8879.n37 GND 0.534939f
C75 a_n10357_8879.n38 GND 1.93072f
C76 a_n10357_8879.t6 GND 0.124293f
C77 a_n10357_8879.n39 GND 0.14217f
C78 a_n10357_8879.n40 GND 0.101555f
C79 a_n10357_8879.t11 GND 0.124293f
C80 a_n10357_8879.n41 GND 0.14217f
C81 a_n10357_8879.n42 GND 0.101555f
C82 a_n10357_8879.n43 GND 2.57726f
C83 a_n10357_8879.t8 GND 0.112567f
C84 a_n10357_8879.n44 GND 0.534939f
C85 a_n10357_8879.t10 GND 0.112567f
C86 a_n1140_n227.n0 GND 2.82523f
C87 a_n1140_n227.n1 GND 1.61528f
C88 a_n1140_n227.n2 GND 1.49303f
C89 a_n1140_n227.t4 GND 0.229329f
C90 a_n1140_n227.t3 GND 0.22933f
C91 a_n1140_n227.t1 GND 0.22933f
C92 a_n1140_n227.t0 GND 0.349146f
C93 a_n1140_n227.t2 GND 0.229329f
C94 VN.t8 GND 0.467313f
C95 VN.t9 GND 0.591597f
C96 VN.n0 GND 0.953702f
C97 VN.t0 GND 0.017019f
C98 VN.t2 GND 0.003039f
C99 VN.t4 GND 0.003039f
C100 VN.n1 GND 0.009856f
C101 VN.n2 GND 0.076517f
C102 VN.t7 GND 0.003039f
C103 VN.t6 GND 0.003039f
C104 VN.n3 GND 0.009856f
C105 VN.n4 GND 0.041354f
C106 VN.t1 GND 0.003039f
C107 VN.t3 GND 0.003039f
C108 VN.n5 GND 0.009856f
C109 VN.n6 GND 0.041354f
C110 VN.t5 GND 0.016916f
C111 VN.n7 GND 0.051252f
C112 VN.n8 GND 1.73904f
C113 VP.t8 GND 0.854597f
C114 VP.t9 GND 1.08301f
C115 VP.n0 GND 1.75127f
C116 VP.t5 GND 0.031033f
C117 VP.t1 GND 0.005542f
C118 VP.t3 GND 0.005542f
C119 VP.n1 GND 0.017973f
C120 VP.n2 GND 0.139525f
C121 VP.t7 GND 0.005542f
C122 VP.t4 GND 0.005542f
C123 VP.n3 GND 0.017973f
C124 VP.n4 GND 0.075408f
C125 VP.t0 GND 0.005542f
C126 VP.t6 GND 0.005542f
C127 VP.n5 GND 0.017973f
C128 VP.n6 GND 0.075408f
C129 VP.t2 GND 0.030845f
C130 VP.n7 GND 0.083704f
C131 VP.n8 GND 2.17023f
C132 VDD.t37 GND 0.009346f
C133 VDD.t30 GND 0.009346f
C134 VDD.n0 GND 0.056787f
C135 VDD.t32 GND 0.009346f
C136 VDD.t19 GND 0.009346f
C137 VDD.n1 GND 0.051072f
C138 VDD.n2 GND 0.326751f
C139 VDD.t3 GND 0.009346f
C140 VDD.t14 GND 0.009346f
C141 VDD.n3 GND 0.051072f
C142 VDD.n4 GND 0.172607f
C143 VDD.t9 GND 0.009346f
C144 VDD.t21 GND 0.009346f
C145 VDD.n5 GND 0.051072f
C146 VDD.n6 GND 0.145479f
C147 VDD.t7 GND 0.009346f
C148 VDD.t16 GND 0.009346f
C149 VDD.n7 GND 0.056787f
C150 VDD.t11 GND 0.009346f
C151 VDD.t5 GND 0.009346f
C152 VDD.n8 GND 0.051072f
C153 VDD.n9 GND 0.326751f
C154 VDD.t23 GND 0.009346f
C155 VDD.t34 GND 0.009346f
C156 VDD.n10 GND 0.051072f
C157 VDD.n11 GND 0.172607f
C158 VDD.t25 GND 0.009346f
C159 VDD.t27 GND 0.009346f
C160 VDD.n12 GND 0.051072f
C161 VDD.n13 GND 0.145479f
C162 VDD.n14 GND 0.10686f
C163 VDD.n15 GND 2.57896f
C164 VDD.t134 GND 0.036671f
C165 VDD.t123 GND 0.005831f
C166 VDD.t126 GND 0.005831f
C167 VDD.n16 GND 0.022552f
C168 VDD.n17 GND 0.173338f
C169 VDD.t111 GND 0.035481f
C170 VDD.n18 GND 0.092021f
C171 VDD.t109 GND 0.036671f
C172 VDD.t127 GND 0.005831f
C173 VDD.t132 GND 0.005831f
C174 VDD.n19 GND 0.022552f
C175 VDD.n20 GND 0.173338f
C176 VDD.t113 GND 0.035481f
C177 VDD.n21 GND 0.084902f
C178 VDD.n22 GND 0.064618f
C179 VDD.t137 GND 0.036671f
C180 VDD.t124 GND 0.005831f
C181 VDD.t130 GND 0.005831f
C182 VDD.n23 GND 0.022552f
C183 VDD.n24 GND 0.173338f
C184 VDD.t112 GND 0.035481f
C185 VDD.n25 GND 0.084902f
C186 VDD.n26 GND 0.123752f
C187 VDD.n27 GND 0.006908f
C188 VDD.n28 GND 0.006908f
C189 VDD.n29 GND 0.00558f
C190 VDD.n30 GND 0.00558f
C191 VDD.n31 GND 0.006932f
C192 VDD.n32 GND 0.006932f
C193 VDD.n33 GND 0.372649f
C194 VDD.n34 GND 0.006932f
C195 VDD.n35 GND 0.006932f
C196 VDD.n36 GND 0.006932f
C197 VDD.n37 GND 0.234769f
C198 VDD.n38 GND 0.006932f
C199 VDD.n39 GND 0.006932f
C200 VDD.n40 GND 0.006932f
C201 VDD.n41 GND 0.006932f
C202 VDD.n42 GND 0.00558f
C203 VDD.n43 GND 0.006932f
C204 VDD.t125 GND 0.186324f
C205 VDD.n44 GND 0.006932f
C206 VDD.n45 GND 0.006932f
C207 VDD.n46 GND 0.006932f
C208 VDD.n47 GND 0.372649f
C209 VDD.n48 GND 0.006932f
C210 VDD.n49 GND 0.006932f
C211 VDD.n50 GND 0.006932f
C212 VDD.n51 GND 0.006932f
C213 VDD.n52 GND 0.006932f
C214 VDD.n53 GND 0.00558f
C215 VDD.n54 GND 0.006932f
C216 VDD.n55 GND 0.006932f
C217 VDD.n56 GND 0.006932f
C218 VDD.n57 GND 0.006932f
C219 VDD.n58 GND 0.372649f
C220 VDD.n59 GND 0.006932f
C221 VDD.n60 GND 0.006932f
C222 VDD.n61 GND 0.006932f
C223 VDD.n62 GND 0.006932f
C224 VDD.n63 GND 0.006932f
C225 VDD.n64 GND 0.00558f
C226 VDD.n65 GND 0.006932f
C227 VDD.n66 GND 0.006932f
C228 VDD.n67 GND 0.006932f
C229 VDD.n68 GND 0.006932f
C230 VDD.n69 GND 0.372649f
C231 VDD.n70 GND 0.006932f
C232 VDD.n71 GND 0.006932f
C233 VDD.n72 GND 0.006932f
C234 VDD.n73 GND 0.006932f
C235 VDD.n74 GND 0.006932f
C236 VDD.n75 GND 0.00558f
C237 VDD.n76 GND 0.006932f
C238 VDD.n77 GND 0.006932f
C239 VDD.n78 GND 0.006932f
C240 VDD.n79 GND 0.006932f
C241 VDD.t39 GND 0.186324f
C242 VDD.n80 GND 0.006932f
C243 VDD.n81 GND 0.006932f
C244 VDD.n82 GND 0.006932f
C245 VDD.n83 GND 0.006932f
C246 VDD.n84 GND 0.006932f
C247 VDD.n85 GND 0.00558f
C248 VDD.n86 GND 0.006932f
C249 VDD.n87 GND 0.283213f
C250 VDD.n88 GND 0.006932f
C251 VDD.n89 GND 0.006932f
C252 VDD.n90 GND 0.016004f
C253 VDD.n91 GND 0.834733f
C254 VDD.n92 GND 0.016092f
C255 VDD.n93 GND 0.006932f
C256 VDD.n94 GND 0.006932f
C257 VDD.n95 GND 0.006932f
C258 VDD.n96 GND 0.006932f
C259 VDD.n97 GND 0.00558f
C260 VDD.n99 GND 0.006932f
C261 VDD.n100 GND 0.006932f
C262 VDD.n101 GND 0.006932f
C263 VDD.n102 GND 0.006932f
C264 VDD.n103 GND 0.004715f
C265 VDD.t48 GND 0.030733f
C266 VDD.t47 GND 0.039858f
C267 VDD.t46 GND 0.203294f
C268 VDD.n104 GND 0.050408f
C269 VDD.n105 GND 0.037394f
C270 VDD.n107 GND 0.006932f
C271 VDD.n108 GND 0.006932f
C272 VDD.n109 GND 0.00558f
C273 VDD.n110 GND 0.006932f
C274 VDD.n112 GND 0.006932f
C275 VDD.n113 GND 0.006932f
C276 VDD.n114 GND 0.006932f
C277 VDD.n115 GND 0.006932f
C278 VDD.n116 GND 0.00558f
C279 VDD.n118 GND 0.006932f
C280 VDD.n119 GND 0.006932f
C281 VDD.n120 GND 0.006932f
C282 VDD.n121 GND 0.005496f
C283 VDD.t59 GND 0.030733f
C284 VDD.t58 GND 0.039858f
C285 VDD.t57 GND 0.203294f
C286 VDD.n122 GND 0.050408f
C287 VDD.n123 GND 0.037394f
C288 VDD.n124 GND 0.006932f
C289 VDD.n125 GND 0.00558f
C290 VDD.n127 GND 0.006932f
C291 VDD.n128 GND 0.00558f
C292 VDD.n129 GND 0.006932f
C293 VDD.n130 GND 0.006932f
C294 VDD.n131 GND 0.006932f
C295 VDD.n132 GND 0.006932f
C296 VDD.n133 GND 0.006932f
C297 VDD.n134 GND 0.003041f
C298 VDD.t41 GND 0.030733f
C299 VDD.t40 GND 0.039858f
C300 VDD.t38 GND 0.203294f
C301 VDD.n136 GND 0.050408f
C302 VDD.n137 GND 0.037394f
C303 VDD.n138 GND 0.008593f
C304 VDD.n139 GND 0.006932f
C305 VDD.n140 GND 0.006932f
C306 VDD.n141 GND 0.006932f
C307 VDD.n142 GND 0.00558f
C308 VDD.n143 GND 0.006932f
C309 VDD.n144 GND 0.006932f
C310 VDD.n145 GND 0.00558f
C311 VDD.n146 GND 0.006932f
C312 VDD.n147 GND 0.006932f
C313 VDD.n148 GND 0.00558f
C314 VDD.n149 GND 0.006932f
C315 VDD.n150 GND 0.006932f
C316 VDD.n151 GND 0.00558f
C317 VDD.n152 GND 0.006932f
C318 VDD.n153 GND 0.006932f
C319 VDD.n154 GND 0.00558f
C320 VDD.n155 GND 0.006932f
C321 VDD.n156 GND 0.00558f
C322 VDD.n157 GND 0.006932f
C323 VDD.n158 GND 0.00558f
C324 VDD.n159 GND 0.006932f
C325 VDD.n160 GND 0.006932f
C326 VDD.n161 GND 0.234769f
C327 VDD.n162 GND 0.006932f
C328 VDD.n163 GND 0.00558f
C329 VDD.n164 GND 0.006932f
C330 VDD.n165 GND 0.00558f
C331 VDD.n166 GND 0.006932f
C332 VDD.n167 GND 0.372649f
C333 VDD.n168 GND 0.006932f
C334 VDD.n169 GND 0.00558f
C335 VDD.n170 GND 0.006932f
C336 VDD.n171 GND 0.00558f
C337 VDD.n172 GND 0.006932f
C338 VDD.n173 GND 0.372649f
C339 VDD.n174 GND 0.006932f
C340 VDD.n175 GND 0.00558f
C341 VDD.n176 GND 0.006932f
C342 VDD.n177 GND 0.00558f
C343 VDD.n178 GND 0.006932f
C344 VDD.n179 GND 0.331657f
C345 VDD.n180 GND 0.006932f
C346 VDD.n181 GND 0.00558f
C347 VDD.n182 GND 0.006932f
C348 VDD.n183 GND 0.00558f
C349 VDD.n184 GND 0.006932f
C350 VDD.n185 GND 0.372649f
C351 VDD.t108 GND 0.186324f
C352 VDD.n186 GND 0.006932f
C353 VDD.n187 GND 0.00558f
C354 VDD.n188 GND 0.006932f
C355 VDD.n189 GND 0.00558f
C356 VDD.n190 GND 0.006932f
C357 VDD.n191 GND 0.372649f
C358 VDD.n192 GND 0.006932f
C359 VDD.n193 GND 0.00558f
C360 VDD.n194 GND 0.006932f
C361 VDD.n195 GND 0.00558f
C362 VDD.n196 GND 0.006932f
C363 VDD.n197 GND 0.372649f
C364 VDD.n198 GND 0.006932f
C365 VDD.n199 GND 0.00558f
C366 VDD.n200 GND 0.006932f
C367 VDD.n201 GND 0.00558f
C368 VDD.n202 GND 0.006932f
C369 VDD.n203 GND 0.372649f
C370 VDD.n204 GND 0.006932f
C371 VDD.n205 GND 0.00558f
C372 VDD.n206 GND 0.006932f
C373 VDD.n207 GND 0.00558f
C374 VDD.n208 GND 0.006932f
C375 VDD.t61 GND 0.186324f
C376 VDD.n209 GND 0.006932f
C377 VDD.n210 GND 0.00558f
C378 VDD.n211 GND 0.006932f
C379 VDD.n212 GND 0.00558f
C380 VDD.n213 GND 0.006932f
C381 VDD.n214 GND 0.372649f
C382 VDD.n215 GND 0.006932f
C383 VDD.n216 GND 0.00558f
C384 VDD.n217 GND 0.029908f
C385 VDD.n218 GND 0.016092f
C386 VDD.n219 GND 2.9402f
C387 VDD.n220 GND 0.016092f
C388 VDD.n221 GND 0.050674f
C389 VDD.n222 GND 0.209537f
C390 VDD.n223 GND 0.003466f
C391 VDD.n224 GND 0.00558f
C392 VDD.n226 GND 0.003466f
C393 VDD.n227 GND 0.003466f
C394 VDD.n228 GND 0.003466f
C395 VDD.n229 GND 0.004603f
C396 VDD.n230 GND 0.006932f
C397 VDD.n231 GND 0.003466f
C398 VDD.n232 GND 0.003466f
C399 VDD.t68 GND 0.030733f
C400 VDD.t69 GND 0.039858f
C401 VDD.t67 GND 0.203294f
C402 VDD.n233 GND 0.050408f
C403 VDD.n234 GND 0.037394f
C404 VDD.n235 GND 0.003466f
C405 VDD.n236 GND 0.003466f
C406 VDD.n237 GND 0.00558f
C407 VDD.n238 GND 0.006932f
C408 VDD.n239 GND 0.003466f
C409 VDD.n240 GND 0.003466f
C410 VDD.n241 GND 0.003466f
C411 VDD.n242 GND 0.00558f
C412 VDD.n243 GND 0.006932f
C413 VDD.n244 GND 0.003466f
C414 VDD.n245 GND 0.003466f
C415 VDD.n246 GND 0.003466f
C416 VDD.t71 GND 0.030733f
C417 VDD.t72 GND 0.039858f
C418 VDD.t70 GND 0.203294f
C419 VDD.n247 GND 0.050408f
C420 VDD.n248 GND 0.037394f
C421 VDD.n249 GND 0.003466f
C422 VDD.n250 GND 0.00558f
C423 VDD.n251 GND 0.006932f
C424 VDD.n252 GND 0.003466f
C425 VDD.n253 GND 0.003466f
C426 VDD.n254 GND 0.003466f
C427 VDD.n255 GND 0.003466f
C428 VDD.n256 GND 0.00558f
C429 VDD.n258 GND 0.006932f
C430 VDD.n259 GND 0.003466f
C431 VDD.n260 GND 0.003466f
C432 VDD.t62 GND 0.030733f
C433 VDD.t63 GND 0.039858f
C434 VDD.t60 GND 0.203294f
C435 VDD.n261 GND 0.050408f
C436 VDD.n262 GND 0.037394f
C437 VDD.n263 GND 0.008593f
C438 VDD.n264 GND 0.003535f
C439 VDD.n265 GND 0.004714f
C440 VDD.n266 GND 0.004714f
C441 VDD.t1 GND 5.15746f
C442 VDD.t15 GND 4.64693f
C443 VDD.t6 GND 4.24074f
C444 VDD.t4 GND 4.24074f
C445 VDD.t10 GND 3.20478f
C446 VDD.n267 GND 1.34899f
C447 VDD.n268 GND 0.004714f
C448 VDD.n269 GND 0.004714f
C449 VDD.t96 GND 0.03345f
C450 VDD.t95 GND 0.055799f
C451 VDD.t93 GND 0.595646f
C452 VDD.n270 GND 0.093248f
C453 VDD.n271 GND 0.071157f
C454 VDD.n272 GND 0.006737f
C455 VDD.n274 GND 0.003189f
C456 VDD.n275 GND 0.011836f
C457 VDD.n276 GND 0.004714f
C458 VDD.n277 GND 0.004714f
C459 VDD.n278 GND 0.253401f
C460 VDD.n279 GND 0.004714f
C461 VDD.n280 GND 0.391281f
C462 VDD.n281 GND 0.004714f
C463 VDD.n282 GND 0.004714f
C464 VDD.n283 GND 0.011836f
C465 VDD.n284 GND 0.004714f
C466 VDD.n285 GND 0.004714f
C467 VDD.n286 GND 0.004714f
C468 VDD.n287 GND 0.004714f
C469 VDD.n288 GND 0.004714f
C470 VDD.n290 GND 0.003535f
C471 VDD.n291 GND 0.004714f
C472 VDD.n292 GND 0.004714f
C473 VDD.n294 GND 0.004714f
C474 VDD.t105 GND 0.03345f
C475 VDD.t104 GND 0.055799f
C476 VDD.t103 GND 0.595646f
C477 VDD.n295 GND 0.093248f
C478 VDD.n296 GND 0.071157f
C479 VDD.n297 GND 0.004714f
C480 VDD.n298 GND 0.004714f
C481 VDD.n299 GND 0.253401f
C482 VDD.n300 GND 0.004714f
C483 VDD.n301 GND 0.004714f
C484 VDD.n302 GND 0.004714f
C485 VDD.n303 GND 0.004714f
C486 VDD.n304 GND 0.004714f
C487 VDD.n305 GND 0.253401f
C488 VDD.n306 GND 0.004714f
C489 VDD.n307 GND 0.004714f
C490 VDD.n308 GND 0.004714f
C491 VDD.n309 GND 0.004714f
C492 VDD.n310 GND 0.004714f
C493 VDD.n311 GND 0.004714f
C494 VDD.n312 GND 0.253401f
C495 VDD.n313 GND 0.004714f
C496 VDD.n314 GND 0.004714f
C497 VDD.n315 GND 0.004714f
C498 VDD.n316 GND 0.004714f
C499 VDD.n317 GND 0.004714f
C500 VDD.t94 GND 0.126701f
C501 VDD.n318 GND 0.004714f
C502 VDD.n319 GND 0.004714f
C503 VDD.n320 GND 0.004714f
C504 VDD.n321 GND 0.004714f
C505 VDD.n322 GND 0.004714f
C506 VDD.n323 GND 0.253401f
C507 VDD.n324 GND 0.004714f
C508 VDD.n325 GND 0.004714f
C509 VDD.n326 GND 0.229179f
C510 VDD.n327 GND 0.004714f
C511 VDD.n328 GND 0.004714f
C512 VDD.n329 GND 0.004714f
C513 VDD.n330 GND 0.20123f
C514 VDD.n331 GND 0.004714f
C515 VDD.n332 GND 0.004714f
C516 VDD.n333 GND 0.004714f
C517 VDD.n334 GND 0.004714f
C518 VDD.n335 GND 0.004714f
C519 VDD.n336 GND 0.253401f
C520 VDD.n337 GND 0.004714f
C521 VDD.n338 GND 0.004714f
C522 VDD.t33 GND 0.126701f
C523 VDD.n339 GND 0.004714f
C524 VDD.n340 GND 0.004714f
C525 VDD.n341 GND 0.004714f
C526 VDD.n342 GND 0.253401f
C527 VDD.n343 GND 0.004714f
C528 VDD.n344 GND 0.004714f
C529 VDD.n345 GND 0.004714f
C530 VDD.n346 GND 0.004714f
C531 VDD.n347 GND 0.004714f
C532 VDD.n348 GND 0.253401f
C533 VDD.n349 GND 0.004714f
C534 VDD.n350 GND 0.004714f
C535 VDD.n351 GND 0.004714f
C536 VDD.n352 GND 0.004714f
C537 VDD.n353 GND 0.004714f
C538 VDD.n354 GND 0.253401f
C539 VDD.n355 GND 0.004714f
C540 VDD.n356 GND 0.004714f
C541 VDD.n357 GND 0.004714f
C542 VDD.n358 GND 0.004714f
C543 VDD.n359 GND 0.004714f
C544 VDD.n360 GND 0.253401f
C545 VDD.n361 GND 0.004714f
C546 VDD.n362 GND 0.004714f
C547 VDD.n363 GND 0.004714f
C548 VDD.n364 GND 0.004714f
C549 VDD.n365 GND 0.004714f
C550 VDD.n366 GND 0.253401f
C551 VDD.n367 GND 0.004714f
C552 VDD.n368 GND 0.004714f
C553 VDD.n369 GND 0.004714f
C554 VDD.n370 GND 0.004714f
C555 VDD.n371 GND 0.004714f
C556 VDD.n372 GND 0.253401f
C557 VDD.n373 GND 0.004714f
C558 VDD.n374 GND 0.004714f
C559 VDD.n375 GND 0.004714f
C560 VDD.n376 GND 0.004714f
C561 VDD.n377 GND 0.004714f
C562 VDD.t35 GND 0.126701f
C563 VDD.n378 GND 0.004714f
C564 VDD.n379 GND 0.004714f
C565 VDD.n380 GND 0.004714f
C566 VDD.n381 GND 0.004714f
C567 VDD.n382 GND 0.004714f
C568 VDD.t22 GND 0.126701f
C569 VDD.n383 GND 0.004714f
C570 VDD.n384 GND 0.004714f
C571 VDD.n385 GND 0.236632f
C572 VDD.n386 GND 0.004714f
C573 VDD.n387 GND 0.004714f
C574 VDD.n388 GND 0.004714f
C575 VDD.n389 GND 0.253401f
C576 VDD.n390 GND 0.004714f
C577 VDD.n391 GND 0.004714f
C578 VDD.n392 GND 0.21241f
C579 VDD.n393 GND 0.004714f
C580 VDD.n394 GND 0.004714f
C581 VDD.n395 GND 0.004714f
C582 VDD.n396 GND 0.253401f
C583 VDD.n397 GND 0.004714f
C584 VDD.n398 GND 0.004714f
C585 VDD.n399 GND 0.004714f
C586 VDD.n400 GND 0.004714f
C587 VDD.n401 GND 0.004714f
C588 VDD.n402 GND 0.253401f
C589 VDD.n403 GND 0.004714f
C590 VDD.n404 GND 0.004714f
C591 VDD.n405 GND 0.004714f
C592 VDD.n406 GND 0.004714f
C593 VDD.n407 GND 0.004714f
C594 VDD.n408 GND 0.253401f
C595 VDD.n409 GND 0.004714f
C596 VDD.n410 GND 0.004714f
C597 VDD.n411 GND 0.004714f
C598 VDD.n412 GND 0.004714f
C599 VDD.n413 GND 0.004714f
C600 VDD.n414 GND 0.253401f
C601 VDD.n415 GND 0.004714f
C602 VDD.n416 GND 0.004714f
C603 VDD.n417 GND 0.004714f
C604 VDD.n418 GND 0.004714f
C605 VDD.n419 GND 0.004714f
C606 VDD.n420 GND 0.253401f
C607 VDD.n421 GND 0.004714f
C608 VDD.n422 GND 0.004714f
C609 VDD.n423 GND 0.004714f
C610 VDD.n424 GND 0.004714f
C611 VDD.n425 GND 0.004714f
C612 VDD.t28 GND 0.126701f
C613 VDD.n426 GND 0.004714f
C614 VDD.n427 GND 0.004714f
C615 VDD.n428 GND 0.004714f
C616 VDD.n429 GND 0.004714f
C617 VDD.n430 GND 0.004714f
C618 VDD.n431 GND 0.134154f
C619 VDD.n432 GND 0.004714f
C620 VDD.n433 GND 0.004714f
C621 VDD.n434 GND 0.14347f
C622 VDD.n435 GND 0.004714f
C623 VDD.n436 GND 0.004714f
C624 VDD.n437 GND 0.004714f
C625 VDD.n438 GND 0.253401f
C626 VDD.n439 GND 0.004714f
C627 VDD.n440 GND 0.004714f
C628 VDD.t26 GND 0.126701f
C629 VDD.n441 GND 0.004714f
C630 VDD.n442 GND 0.004714f
C631 VDD.n443 GND 0.004714f
C632 VDD.n444 GND 0.253401f
C633 VDD.n445 GND 0.004714f
C634 VDD.n446 GND 0.004714f
C635 VDD.n447 GND 0.004714f
C636 VDD.n448 GND 0.004714f
C637 VDD.n449 GND 0.004714f
C638 VDD.n450 GND 0.253401f
C639 VDD.n451 GND 0.004714f
C640 VDD.n452 GND 0.004714f
C641 VDD.n453 GND 0.004714f
C642 VDD.n454 GND 0.004714f
C643 VDD.n455 GND 0.004714f
C644 VDD.n456 GND 0.253401f
C645 VDD.n457 GND 0.004714f
C646 VDD.n458 GND 0.004714f
C647 VDD.n459 GND 0.004714f
C648 VDD.n460 GND 0.004714f
C649 VDD.n461 GND 0.004714f
C650 VDD.n462 GND 0.253401f
C651 VDD.n463 GND 0.004714f
C652 VDD.n464 GND 0.004714f
C653 VDD.n465 GND 0.004714f
C654 VDD.n466 GND 0.004714f
C655 VDD.n467 GND 0.004714f
C656 VDD.n468 GND 0.253401f
C657 VDD.n469 GND 0.004714f
C658 VDD.n470 GND 0.004714f
C659 VDD.n471 GND 0.004714f
C660 VDD.n472 GND 0.004714f
C661 VDD.n473 GND 0.004714f
C662 VDD.n474 GND 0.253401f
C663 VDD.n475 GND 0.004714f
C664 VDD.n476 GND 0.004714f
C665 VDD.n477 GND 0.004714f
C666 VDD.n478 GND 0.004714f
C667 VDD.n479 GND 0.004714f
C668 VDD.n480 GND 0.227316f
C669 VDD.n481 GND 0.004714f
C670 VDD.n482 GND 0.004714f
C671 VDD.n483 GND 0.004714f
C672 VDD.n484 GND 0.004714f
C673 VDD.n485 GND 0.004714f
C674 VDD.t54 GND 0.126701f
C675 VDD.n486 GND 0.004714f
C676 VDD.n487 GND 0.004714f
C677 VDD.t24 GND 0.126701f
C678 VDD.n488 GND 0.004714f
C679 VDD.n489 GND 0.004714f
C680 VDD.n490 GND 0.004714f
C681 VDD.n491 GND 0.253401f
C682 VDD.n492 GND 0.004714f
C683 VDD.n493 GND 0.004714f
C684 VDD.n494 GND 0.150923f
C685 VDD.n495 GND 0.004714f
C686 VDD.n496 GND 0.004714f
C687 VDD.n497 GND 0.004714f
C688 VDD.n498 GND 0.253401f
C689 VDD.n499 GND 0.004714f
C690 VDD.n500 GND 0.004714f
C691 VDD.n501 GND 0.004714f
C692 VDD.n502 GND 0.004714f
C693 VDD.n503 GND 0.004714f
C694 VDD.n504 GND 0.253401f
C695 VDD.n505 GND 0.004714f
C696 VDD.n506 GND 0.004714f
C697 VDD.n507 GND 0.004714f
C698 VDD.n508 GND 0.004714f
C699 VDD.n509 GND 0.004714f
C700 VDD.n510 GND 0.253401f
C701 VDD.n511 GND 0.004714f
C702 VDD.n512 GND 0.004714f
C703 VDD.n513 GND 0.004714f
C704 VDD.n514 GND 0.012357f
C705 VDD.n515 GND 0.012357f
C706 VDD.n516 GND 0.391281f
C707 VDD.n532 GND 0.004714f
C708 VDD.n533 GND 0.011836f
C709 VDD.n534 GND 0.003189f
C710 VDD.n535 GND 0.004714f
C711 VDD.n536 GND 0.004714f
C712 VDD.n537 GND 0.253401f
C713 VDD.n538 GND 0.004714f
C714 VDD.n539 GND 0.004714f
C715 VDD.n540 GND 0.004714f
C716 VDD.n541 GND 0.011836f
C717 VDD.n542 GND 0.004714f
C718 VDD.t88 GND 0.03345f
C719 VDD.t87 GND 0.055799f
C720 VDD.t86 GND 0.595646f
C721 VDD.n543 GND 0.093248f
C722 VDD.n544 GND 0.071157f
C723 VDD.n545 GND 0.006737f
C724 VDD.n546 GND 0.004714f
C725 VDD.n547 GND 0.004714f
C726 VDD.n548 GND 0.253401f
C727 VDD.n549 GND 0.004714f
C728 VDD.n550 GND 0.004714f
C729 VDD.n551 GND 0.004714f
C730 VDD.n552 GND 0.004714f
C731 VDD.n553 GND 0.004714f
C732 VDD.n554 GND 0.253401f
C733 VDD.n555 GND 0.004714f
C734 VDD.n556 GND 0.004714f
C735 VDD.n557 GND 0.004714f
C736 VDD.n558 GND 0.004714f
C737 VDD.n559 GND 0.004714f
C738 VDD.n560 GND 0.004714f
C739 VDD.n561 GND 0.253401f
C740 VDD.n562 GND 0.004714f
C741 VDD.n563 GND 0.004714f
C742 VDD.n564 GND 0.004714f
C743 VDD.n565 GND 0.004714f
C744 VDD.n566 GND 0.004714f
C745 VDD.t50 GND 0.126701f
C746 VDD.n567 GND 0.004714f
C747 VDD.n568 GND 0.004714f
C748 VDD.n569 GND 0.004714f
C749 VDD.n570 GND 0.004714f
C750 VDD.n571 GND 0.004714f
C751 VDD.n572 GND 0.253401f
C752 VDD.n573 GND 0.004714f
C753 VDD.n574 GND 0.004714f
C754 VDD.t20 GND 0.126701f
C755 VDD.n575 GND 0.004714f
C756 VDD.n576 GND 0.004714f
C757 VDD.n577 GND 0.004714f
C758 VDD.n578 GND 0.253401f
C759 VDD.n579 GND 0.004714f
C760 VDD.n580 GND 0.004714f
C761 VDD.n581 GND 0.004714f
C762 VDD.n582 GND 0.004714f
C763 VDD.n583 GND 0.004714f
C764 VDD.n584 GND 0.253401f
C765 VDD.n585 GND 0.004714f
C766 VDD.n586 GND 0.004714f
C767 VDD.n587 GND 0.004714f
C768 VDD.n588 GND 0.004714f
C769 VDD.n589 GND 0.004714f
C770 VDD.n590 GND 0.253401f
C771 VDD.n591 GND 0.004714f
C772 VDD.n592 GND 0.004714f
C773 VDD.n593 GND 0.004714f
C774 VDD.n594 GND 0.004714f
C775 VDD.n595 GND 0.004714f
C776 VDD.n596 GND 0.253401f
C777 VDD.n597 GND 0.004714f
C778 VDD.n598 GND 0.004714f
C779 VDD.n599 GND 0.004714f
C780 VDD.n600 GND 0.004714f
C781 VDD.n601 GND 0.004714f
C782 VDD.n602 GND 0.253401f
C783 VDD.n603 GND 0.004714f
C784 VDD.n604 GND 0.004714f
C785 VDD.n605 GND 0.004714f
C786 VDD.n606 GND 0.004714f
C787 VDD.n607 GND 0.004714f
C788 VDD.n608 GND 0.253401f
C789 VDD.n609 GND 0.004714f
C790 VDD.n610 GND 0.004714f
C791 VDD.n611 GND 0.004714f
C792 VDD.n612 GND 0.004714f
C793 VDD.n613 GND 0.004714f
C794 VDD.n614 GND 0.245948f
C795 VDD.n615 GND 0.004714f
C796 VDD.n616 GND 0.004714f
C797 VDD.n617 GND 0.004714f
C798 VDD.n618 GND 0.004714f
C799 VDD.n619 GND 0.004714f
C800 VDD.n620 GND 0.253401f
C801 VDD.n621 GND 0.004714f
C802 VDD.n622 GND 0.004714f
C803 VDD.t8 GND 0.126701f
C804 VDD.n623 GND 0.004714f
C805 VDD.n624 GND 0.004714f
C806 VDD.n625 GND 0.004714f
C807 VDD.t17 GND 0.126701f
C808 VDD.n626 GND 0.004714f
C809 VDD.n627 GND 0.004714f
C810 VDD.n628 GND 0.004714f
C811 VDD.n629 GND 0.004714f
C812 VDD.n630 GND 0.004714f
C813 VDD.n631 GND 0.253401f
C814 VDD.n632 GND 0.004714f
C815 VDD.n633 GND 0.004714f
C816 VDD.n634 GND 0.236632f
C817 VDD.n635 GND 0.004714f
C818 VDD.n636 GND 0.004714f
C819 VDD.n637 GND 0.004714f
C820 VDD.n638 GND 0.253401f
C821 VDD.n639 GND 0.004714f
C822 VDD.n640 GND 0.004714f
C823 VDD.n641 GND 0.004714f
C824 VDD.n642 GND 0.004714f
C825 VDD.n643 GND 0.004714f
C826 VDD.n644 GND 0.253401f
C827 VDD.n645 GND 0.004714f
C828 VDD.n646 GND 0.004714f
C829 VDD.n647 GND 0.004714f
C830 VDD.n648 GND 0.004714f
C831 VDD.n649 GND 0.004714f
C832 VDD.n650 GND 0.253401f
C833 VDD.n651 GND 0.004714f
C834 VDD.n652 GND 0.004714f
C835 VDD.n653 GND 0.004714f
C836 VDD.n654 GND 0.004714f
C837 VDD.n655 GND 0.004714f
C838 VDD.n656 GND 0.253401f
C839 VDD.n657 GND 0.004714f
C840 VDD.n658 GND 0.004714f
C841 VDD.n659 GND 0.004714f
C842 VDD.n660 GND 0.004714f
C843 VDD.n661 GND 0.004714f
C844 VDD.n662 GND 0.253401f
C845 VDD.n663 GND 0.004714f
C846 VDD.n664 GND 0.004714f
C847 VDD.n665 GND 0.004714f
C848 VDD.n666 GND 0.004714f
C849 VDD.n667 GND 0.004714f
C850 VDD.t13 GND 0.126701f
C851 VDD.n668 GND 0.004714f
C852 VDD.n669 GND 0.004714f
C853 VDD.n670 GND 0.004714f
C854 VDD.n671 GND 0.004714f
C855 VDD.n672 GND 0.004714f
C856 VDD.t12 GND 0.126701f
C857 VDD.n673 GND 0.004714f
C858 VDD.n674 GND 0.004714f
C859 VDD.n675 GND 0.167692f
C860 VDD.n676 GND 0.004714f
C861 VDD.n677 GND 0.004714f
C862 VDD.n678 GND 0.004714f
C863 VDD.n679 GND 0.253401f
C864 VDD.n680 GND 0.004714f
C865 VDD.n681 GND 0.004714f
C866 VDD.n682 GND 0.14347f
C867 VDD.n683 GND 0.004714f
C868 VDD.n684 GND 0.004714f
C869 VDD.n685 GND 0.004714f
C870 VDD.n686 GND 0.253401f
C871 VDD.n687 GND 0.004714f
C872 VDD.n688 GND 0.004714f
C873 VDD.n689 GND 0.004714f
C874 VDD.n690 GND 0.004714f
C875 VDD.n691 GND 0.004714f
C876 VDD.n692 GND 0.253401f
C877 VDD.n693 GND 0.004714f
C878 VDD.n694 GND 0.004714f
C879 VDD.n695 GND 0.004714f
C880 VDD.n696 GND 0.004714f
C881 VDD.n697 GND 0.004714f
C882 VDD.n698 GND 0.253401f
C883 VDD.n699 GND 0.004714f
C884 VDD.n700 GND 0.004714f
C885 VDD.n701 GND 0.004714f
C886 VDD.n702 GND 0.004714f
C887 VDD.n703 GND 0.004714f
C888 VDD.n704 GND 0.253401f
C889 VDD.n705 GND 0.004714f
C890 VDD.n706 GND 0.004714f
C891 VDD.n707 GND 0.004714f
C892 VDD.n708 GND 0.004714f
C893 VDD.n709 GND 0.004714f
C894 VDD.n710 GND 0.253401f
C895 VDD.n711 GND 0.004714f
C896 VDD.n712 GND 0.004714f
C897 VDD.n713 GND 0.004714f
C898 VDD.n714 GND 0.004714f
C899 VDD.n715 GND 0.004714f
C900 VDD.n716 GND 0.178871f
C901 VDD.n717 GND 0.004714f
C902 VDD.n718 GND 0.004714f
C903 VDD.n719 GND 0.004714f
C904 VDD.n720 GND 0.004714f
C905 VDD.n721 GND 0.004714f
C906 VDD.n722 GND 0.253401f
C907 VDD.n723 GND 0.004714f
C908 VDD.n724 GND 0.004714f
C909 VDD.t2 GND 0.126701f
C910 VDD.n725 GND 0.004714f
C911 VDD.n726 GND 0.004714f
C912 VDD.n727 GND 0.004714f
C913 VDD.n728 GND 0.253401f
C914 VDD.n729 GND 0.004714f
C915 VDD.n730 GND 0.004714f
C916 VDD.n731 GND 0.004714f
C917 VDD.n732 GND 0.004714f
C918 VDD.n733 GND 0.004714f
C919 VDD.t43 GND 0.126701f
C920 VDD.n734 GND 0.004714f
C921 VDD.n735 GND 0.004714f
C922 VDD.n736 GND 0.004714f
C923 VDD.n737 GND 0.004714f
C924 VDD.n738 GND 0.004714f
C925 VDD.n739 GND 0.253401f
C926 VDD.n740 GND 0.004714f
C927 VDD.n741 GND 0.004714f
C928 VDD.n742 GND 0.150923f
C929 VDD.n743 GND 0.004714f
C930 VDD.n744 GND 0.004714f
C931 VDD.n745 GND 0.004714f
C932 VDD.n746 GND 0.253401f
C933 VDD.n747 GND 0.004714f
C934 VDD.n748 GND 0.004714f
C935 VDD.n749 GND 0.004714f
C936 VDD.n750 GND 0.004714f
C937 VDD.n751 GND 0.004714f
C938 VDD.n752 GND 0.253401f
C939 VDD.n753 GND 0.004714f
C940 VDD.n754 GND 0.004714f
C941 VDD.n755 GND 0.004714f
C942 VDD.n756 GND 0.004714f
C943 VDD.n757 GND 0.004714f
C944 VDD.n758 GND 0.253401f
C945 VDD.n759 GND 0.004714f
C946 VDD.n760 GND 0.004714f
C947 VDD.n761 GND 0.004714f
C948 VDD.n762 GND 0.012357f
C949 VDD.n763 GND 0.012357f
C950 VDD.n764 GND 1.34899f
C951 VDD.n765 GND 0.011836f
C952 VDD.n766 GND 0.011836f
C953 VDD.n767 GND 0.012357f
C954 VDD.n768 GND 0.004714f
C955 VDD.n770 GND 0.004714f
C956 VDD.n771 GND 0.004714f
C957 VDD.n772 GND 0.003535f
C958 VDD.n773 GND 0.010251f
C959 VDD.n774 GND 0.003535f
C960 VDD.n775 GND 0.004714f
C961 VDD.n776 GND 0.004714f
C962 VDD.n777 GND 0.004714f
C963 VDD.n779 GND 0.004714f
C964 VDD.n780 GND 0.004714f
C965 VDD.n781 GND 0.004714f
C966 VDD.n782 GND 0.004714f
C967 VDD.n784 GND 0.004714f
C968 VDD.n786 GND 0.004714f
C969 VDD.n787 GND 0.004714f
C970 VDD.n788 GND 0.004714f
C971 VDD.n789 GND 0.004714f
C972 VDD.n790 GND 0.004714f
C973 VDD.n792 GND 0.004714f
C974 VDD.n794 GND 0.004714f
C975 VDD.n795 GND 0.004714f
C976 VDD.t44 GND 0.03345f
C977 VDD.t45 GND 0.055799f
C978 VDD.t42 GND 0.595646f
C979 VDD.n796 GND 0.093248f
C980 VDD.n797 GND 0.071157f
C981 VDD.n798 GND 0.004714f
C982 VDD.n799 GND 0.004714f
C983 VDD.n800 GND 0.004714f
C984 VDD.n801 GND 0.004714f
C985 VDD.n802 GND 0.004714f
C986 VDD.n803 GND 0.004714f
C987 VDD.n804 GND 0.004714f
C988 VDD.n805 GND 0.004714f
C989 VDD.n806 GND 0.004714f
C990 VDD.n807 GND 0.004714f
C991 VDD.n808 GND 0.003189f
C992 VDD.n809 GND 0.004714f
C993 VDD.n810 GND 0.004714f
C994 VDD.n812 GND 0.004714f
C995 VDD.n813 GND 0.004714f
C996 VDD.n814 GND 0.004714f
C997 VDD.n816 GND 0.004714f
C998 VDD.n818 GND 0.004714f
C999 VDD.n819 GND 0.004714f
C1000 VDD.n820 GND 0.004714f
C1001 VDD.t78 GND 0.03345f
C1002 VDD.t79 GND 0.055799f
C1003 VDD.t77 GND 0.595646f
C1004 VDD.n821 GND 0.093248f
C1005 VDD.n822 GND 0.071157f
C1006 VDD.n823 GND 0.006737f
C1007 VDD.n824 GND 0.003882f
C1008 VDD.n825 GND 0.004714f
C1009 VDD.n827 GND 0.004714f
C1010 VDD.n828 GND 0.012357f
C1011 VDD.n829 GND 0.012357f
C1012 VDD.n830 GND 0.011836f
C1013 VDD.n831 GND 0.004714f
C1014 VDD.n832 GND 0.004714f
C1015 VDD.n833 GND 0.004714f
C1016 VDD.n834 GND 0.004714f
C1017 VDD.n835 GND 0.004714f
C1018 VDD.n836 GND 0.004714f
C1019 VDD.n837 GND 0.004714f
C1020 VDD.n838 GND 0.004714f
C1021 VDD.n839 GND 0.004714f
C1022 VDD.n840 GND 0.004714f
C1023 VDD.n841 GND 0.004714f
C1024 VDD.n842 GND 0.004714f
C1025 VDD.n843 GND 0.004714f
C1026 VDD.n844 GND 0.004714f
C1027 VDD.n845 GND 0.004714f
C1028 VDD.n846 GND 0.004714f
C1029 VDD.n847 GND 0.004714f
C1030 VDD.n848 GND 0.004714f
C1031 VDD.n849 GND 0.004714f
C1032 VDD.n850 GND 0.004714f
C1033 VDD.n851 GND 0.004714f
C1034 VDD.n852 GND 0.004714f
C1035 VDD.n853 GND 0.004714f
C1036 VDD.n854 GND 0.004714f
C1037 VDD.n855 GND 0.004714f
C1038 VDD.n856 GND 0.004714f
C1039 VDD.n857 GND 0.004714f
C1040 VDD.n858 GND 0.004714f
C1041 VDD.n859 GND 0.004714f
C1042 VDD.n860 GND 0.004714f
C1043 VDD.n861 GND 0.004714f
C1044 VDD.n862 GND 0.004714f
C1045 VDD.n863 GND 0.004714f
C1046 VDD.n864 GND 0.004714f
C1047 VDD.n865 GND 0.004714f
C1048 VDD.n866 GND 0.004714f
C1049 VDD.n867 GND 0.004714f
C1050 VDD.n868 GND 0.004714f
C1051 VDD.n869 GND 0.004714f
C1052 VDD.n870 GND 0.004714f
C1053 VDD.n871 GND 0.004714f
C1054 VDD.n872 GND 0.004714f
C1055 VDD.n873 GND 0.004714f
C1056 VDD.n874 GND 0.004714f
C1057 VDD.n875 GND 0.004714f
C1058 VDD.n876 GND 0.004714f
C1059 VDD.n877 GND 0.004714f
C1060 VDD.n878 GND 0.004714f
C1061 VDD.n879 GND 0.004714f
C1062 VDD.n880 GND 0.004714f
C1063 VDD.n881 GND 0.004714f
C1064 VDD.n882 GND 0.004714f
C1065 VDD.n883 GND 0.004714f
C1066 VDD.n884 GND 0.004714f
C1067 VDD.n885 GND 0.004714f
C1068 VDD.n886 GND 0.004714f
C1069 VDD.n887 GND 0.004714f
C1070 VDD.n888 GND 0.004714f
C1071 VDD.n889 GND 0.004714f
C1072 VDD.n890 GND 0.004714f
C1073 VDD.n891 GND 0.004714f
C1074 VDD.n892 GND 0.004714f
C1075 VDD.n893 GND 0.004714f
C1076 VDD.n894 GND 0.004714f
C1077 VDD.n895 GND 0.004714f
C1078 VDD.n896 GND 0.004714f
C1079 VDD.n897 GND 0.004714f
C1080 VDD.n898 GND 0.004714f
C1081 VDD.n899 GND 0.004714f
C1082 VDD.n900 GND 0.004714f
C1083 VDD.n901 GND 0.004714f
C1084 VDD.n902 GND 0.004714f
C1085 VDD.n903 GND 0.004714f
C1086 VDD.n904 GND 0.004714f
C1087 VDD.n905 GND 0.004714f
C1088 VDD.n906 GND 0.004714f
C1089 VDD.n907 GND 0.004714f
C1090 VDD.n908 GND 0.004714f
C1091 VDD.n909 GND 0.004714f
C1092 VDD.n910 GND 0.004714f
C1093 VDD.n911 GND 0.004714f
C1094 VDD.n912 GND 0.004714f
C1095 VDD.n913 GND 0.004714f
C1096 VDD.n914 GND 0.004714f
C1097 VDD.n915 GND 0.004714f
C1098 VDD.n916 GND 0.004714f
C1099 VDD.n917 GND 0.004714f
C1100 VDD.n918 GND 0.004714f
C1101 VDD.n919 GND 0.004714f
C1102 VDD.n920 GND 0.004714f
C1103 VDD.n921 GND 0.004714f
C1104 VDD.n922 GND 0.004714f
C1105 VDD.n923 GND 0.004714f
C1106 VDD.n924 GND 0.004714f
C1107 VDD.n925 GND 0.004714f
C1108 VDD.n926 GND 0.004714f
C1109 VDD.n927 GND 0.004714f
C1110 VDD.n928 GND 0.004714f
C1111 VDD.n929 GND 0.004714f
C1112 VDD.n930 GND 0.004714f
C1113 VDD.n931 GND 0.004714f
C1114 VDD.n932 GND 0.004714f
C1115 VDD.n933 GND 0.004714f
C1116 VDD.n934 GND 0.004714f
C1117 VDD.n935 GND 0.004714f
C1118 VDD.n936 GND 0.004714f
C1119 VDD.n937 GND 0.128564f
C1120 VDD.n938 GND 0.004714f
C1121 VDD.n939 GND 0.004714f
C1122 VDD.n940 GND 0.004714f
C1123 VDD.n941 GND 0.004714f
C1124 VDD.n942 GND 0.004714f
C1125 VDD.n943 GND 0.004714f
C1126 VDD.n944 GND 0.004714f
C1127 VDD.n945 GND 0.004714f
C1128 VDD.n946 GND 0.004714f
C1129 VDD.n947 GND 0.004714f
C1130 VDD.n948 GND 0.004714f
C1131 VDD.n949 GND 0.004714f
C1132 VDD.n950 GND 0.004714f
C1133 VDD.n951 GND 0.004714f
C1134 VDD.n952 GND 0.004714f
C1135 VDD.n953 GND 0.004714f
C1136 VDD.n954 GND 0.004714f
C1137 VDD.n955 GND 0.004714f
C1138 VDD.n956 GND 0.004714f
C1139 VDD.n957 GND 0.004714f
C1140 VDD.n958 GND 0.004714f
C1141 VDD.n959 GND 0.004714f
C1142 VDD.n960 GND 0.004714f
C1143 VDD.n961 GND 0.004714f
C1144 VDD.n962 GND 0.004714f
C1145 VDD.n963 GND 0.004714f
C1146 VDD.n964 GND 0.004714f
C1147 VDD.n965 GND 0.004714f
C1148 VDD.n966 GND 0.004714f
C1149 VDD.n967 GND 0.004714f
C1150 VDD.n968 GND 0.004714f
C1151 VDD.n969 GND 0.004714f
C1152 VDD.n970 GND 0.004714f
C1153 VDD.n971 GND 0.004714f
C1154 VDD.n972 GND 0.004714f
C1155 VDD.n973 GND 0.004714f
C1156 VDD.n974 GND 0.004714f
C1157 VDD.n975 GND 0.004714f
C1158 VDD.n976 GND 0.004714f
C1159 VDD.n977 GND 0.004714f
C1160 VDD.n978 GND 0.004714f
C1161 VDD.n979 GND 0.004714f
C1162 VDD.n980 GND 0.004714f
C1163 VDD.n981 GND 0.004714f
C1164 VDD.n982 GND 0.004714f
C1165 VDD.n983 GND 0.004714f
C1166 VDD.n984 GND 0.004714f
C1167 VDD.n985 GND 0.004714f
C1168 VDD.n986 GND 0.004714f
C1169 VDD.n987 GND 0.004714f
C1170 VDD.n988 GND 0.004714f
C1171 VDD.n989 GND 0.004714f
C1172 VDD.n990 GND 0.004714f
C1173 VDD.n991 GND 0.004714f
C1174 VDD.n992 GND 0.004714f
C1175 VDD.n993 GND 0.004714f
C1176 VDD.n994 GND 0.004714f
C1177 VDD.n995 GND 0.004714f
C1178 VDD.n996 GND 0.004714f
C1179 VDD.n997 GND 0.004714f
C1180 VDD.n998 GND 0.004714f
C1181 VDD.n999 GND 0.004714f
C1182 VDD.n1000 GND 0.004714f
C1183 VDD.n1001 GND 0.004714f
C1184 VDD.n1002 GND 0.004714f
C1185 VDD.n1003 GND 0.004714f
C1186 VDD.n1004 GND 0.004714f
C1187 VDD.n1005 GND 0.004714f
C1188 VDD.n1006 GND 0.004714f
C1189 VDD.n1007 GND 0.004714f
C1190 VDD.n1008 GND 0.004714f
C1191 VDD.n1009 GND 0.004714f
C1192 VDD.n1010 GND 0.004714f
C1193 VDD.n1011 GND 0.004714f
C1194 VDD.n1012 GND 0.004714f
C1195 VDD.n1013 GND 0.004714f
C1196 VDD.n1014 GND 0.004714f
C1197 VDD.n1015 GND 0.004714f
C1198 VDD.n1016 GND 0.004714f
C1199 VDD.n1017 GND 0.004714f
C1200 VDD.n1018 GND 0.004714f
C1201 VDD.n1019 GND 0.004714f
C1202 VDD.n1020 GND 0.004714f
C1203 VDD.n1021 GND 0.004714f
C1204 VDD.n1022 GND 0.004714f
C1205 VDD.n1023 GND 0.004714f
C1206 VDD.n1024 GND 0.004714f
C1207 VDD.n1025 GND 0.004714f
C1208 VDD.n1026 GND 0.004714f
C1209 VDD.n1027 GND 0.004714f
C1210 VDD.n1028 GND 0.004714f
C1211 VDD.n1029 GND 0.004714f
C1212 VDD.n1030 GND 0.004714f
C1213 VDD.n1031 GND 0.004714f
C1214 VDD.n1032 GND 0.004714f
C1215 VDD.n1033 GND 0.004714f
C1216 VDD.n1034 GND 0.004714f
C1217 VDD.n1035 GND 0.004714f
C1218 VDD.n1036 GND 0.011836f
C1219 VDD.n1038 GND 0.012357f
C1220 VDD.n1039 GND 0.012357f
C1221 VDD.n1040 GND 0.003189f
C1222 VDD.n1041 GND 0.006737f
C1223 VDD.n1042 GND 0.003882f
C1224 VDD.n1043 GND 0.004714f
C1225 VDD.n1045 GND 0.004714f
C1226 VDD.n1046 GND 0.004714f
C1227 VDD.n1047 GND 0.004714f
C1228 VDD.n1048 GND 0.004714f
C1229 VDD.n1049 GND 0.004714f
C1230 VDD.n1050 GND 0.004714f
C1231 VDD.n1052 GND 0.004714f
C1232 VDD.n1053 GND 0.003535f
C1233 VDD.n1054 GND 0.211802f
C1234 VDD.n1055 GND 2.09122f
C1235 VDD.n1056 GND 0.003466f
C1236 VDD.n1057 GND 0.003466f
C1237 VDD.n1058 GND 0.00558f
C1238 VDD.n1059 GND 0.006932f
C1239 VDD.n1060 GND 0.006932f
C1240 VDD.n1061 GND 0.006932f
C1241 VDD.t102 GND 0.030733f
C1242 VDD.t101 GND 0.039858f
C1243 VDD.t100 GND 0.203294f
C1244 VDD.n1062 GND 0.050408f
C1245 VDD.n1063 GND 0.037394f
C1246 VDD.n1064 GND 0.011382f
C1247 VDD.n1065 GND 0.003466f
C1248 VDD.n1066 GND 0.006932f
C1249 VDD.n1067 GND 0.006932f
C1250 VDD.n1068 GND 0.006932f
C1251 VDD.n1069 GND 0.00558f
C1252 VDD.n1070 GND 0.003466f
C1253 VDD.n1071 GND 0.006932f
C1254 VDD.n1072 GND 0.006932f
C1255 VDD.n1073 GND 0.006932f
C1256 VDD.n1074 GND 0.003041f
C1257 VDD.n1075 GND 0.009175f
C1258 VDD.t92 GND 0.030733f
C1259 VDD.t91 GND 0.039858f
C1260 VDD.t89 GND 0.203294f
C1261 VDD.n1076 GND 0.050408f
C1262 VDD.n1077 GND 0.037394f
C1263 VDD.n1078 GND 0.008593f
C1264 VDD.n1079 GND 0.006932f
C1265 VDD.n1080 GND 0.016004f
C1266 VDD.n1081 GND 0.495623f
C1267 VDD.n1087 GND 0.006932f
C1268 VDD.n1088 GND 0.00558f
C1269 VDD.n1089 GND 0.003466f
C1270 VDD.n1090 GND 0.004603f
C1271 VDD.t99 GND 0.030733f
C1272 VDD.t98 GND 0.039858f
C1273 VDD.t97 GND 0.203294f
C1274 VDD.n1091 GND 0.050408f
C1275 VDD.n1092 GND 0.037394f
C1276 VDD.n1093 GND 0.003466f
C1277 VDD.n1094 GND 0.00558f
C1278 VDD.n1095 GND 0.006932f
C1279 VDD.n1096 GND 0.006932f
C1280 VDD.n1097 GND 0.006932f
C1281 VDD.n1098 GND 0.00558f
C1282 VDD.n1099 GND 0.006932f
C1283 VDD.n1100 GND 0.00558f
C1284 VDD.n1101 GND 0.006932f
C1285 VDD.n1102 GND 0.283213f
C1286 VDD.n1103 GND 0.006932f
C1287 VDD.n1104 GND 0.00558f
C1288 VDD.n1105 GND 0.004631f
C1289 VDD.n1106 GND 0.006932f
C1290 VDD.n1107 GND 0.00558f
C1291 VDD.n1108 GND 0.006932f
C1292 VDD.n1109 GND 0.372649f
C1293 VDD.t90 GND 0.186324f
C1294 VDD.n1110 GND 0.006932f
C1295 VDD.n1111 GND 0.00558f
C1296 VDD.n1112 GND 0.006932f
C1297 VDD.n1113 GND 0.00558f
C1298 VDD.n1114 GND 0.006932f
C1299 VDD.n1115 GND 0.372649f
C1300 VDD.n1116 GND 0.006932f
C1301 VDD.n1117 GND 0.00558f
C1302 VDD.n1118 GND 0.00558f
C1303 VDD.n1119 GND 0.006932f
C1304 VDD.n1120 GND 0.00558f
C1305 VDD.n1121 GND 0.006932f
C1306 VDD.n1122 GND 0.372649f
C1307 VDD.n1123 GND 0.006932f
C1308 VDD.n1124 GND 0.00558f
C1309 VDD.n1125 GND 0.006932f
C1310 VDD.n1126 GND 0.00558f
C1311 VDD.n1127 GND 0.006932f
C1312 VDD.n1128 GND 0.372649f
C1313 VDD.n1129 GND 0.006932f
C1314 VDD.n1130 GND 0.00558f
C1315 VDD.n1131 GND 0.006932f
C1316 VDD.n1132 GND 0.00558f
C1317 VDD.n1133 GND 0.006932f
C1318 VDD.t128 GND 0.186324f
C1319 VDD.n1134 GND 0.006932f
C1320 VDD.n1135 GND 0.00558f
C1321 VDD.n1136 GND 0.006932f
C1322 VDD.n1137 GND 0.00558f
C1323 VDD.n1138 GND 0.006932f
C1324 VDD.n1139 GND 0.372649f
C1325 VDD.n1140 GND 0.006932f
C1326 VDD.n1141 GND 0.00558f
C1327 VDD.n1142 GND 0.006932f
C1328 VDD.n1143 GND 0.00558f
C1329 VDD.n1144 GND 0.006932f
C1330 VDD.n1145 GND 0.372649f
C1331 VDD.n1146 GND 0.006932f
C1332 VDD.n1147 GND 0.00558f
C1333 VDD.n1148 GND 0.006932f
C1334 VDD.n1149 GND 0.00558f
C1335 VDD.n1150 GND 0.006932f
C1336 VDD.t106 GND 0.186324f
C1337 VDD.n1151 GND 0.006932f
C1338 VDD.n1152 GND 0.00558f
C1339 VDD.n1153 GND 0.006932f
C1340 VDD.n1154 GND 0.00558f
C1341 VDD.n1155 GND 0.006932f
C1342 VDD.n1156 GND 0.372649f
C1343 VDD.n1157 GND 0.234769f
C1344 VDD.n1158 GND 0.006932f
C1345 VDD.n1159 GND 0.00558f
C1346 VDD.n1160 GND 0.006908f
C1347 VDD.n1161 GND 0.00558f
C1348 VDD.n1162 GND 0.006932f
C1349 VDD.n1163 GND 0.372649f
C1350 VDD.n1164 GND 0.006932f
C1351 VDD.n1165 GND 0.00558f
C1352 VDD.n1166 GND 0.006932f
C1353 VDD.n1167 GND 0.00558f
C1354 VDD.n1168 GND 0.006932f
C1355 VDD.n1169 GND 0.234769f
C1356 VDD.n1170 GND 0.006932f
C1357 VDD.n1171 GND 0.00558f
C1358 VDD.n1172 GND 0.006932f
C1359 VDD.n1173 GND 0.00558f
C1360 VDD.n1174 GND 0.006932f
C1361 VDD.n1175 GND 0.372649f
C1362 VDD.n1176 GND 0.006932f
C1363 VDD.n1177 GND 0.00558f
C1364 VDD.n1178 GND 0.006932f
C1365 VDD.n1179 GND 0.00558f
C1366 VDD.n1180 GND 0.006932f
C1367 VDD.n1181 GND 0.372649f
C1368 VDD.n1182 GND 0.006932f
C1369 VDD.n1183 GND 0.00558f
C1370 VDD.n1184 GND 0.006932f
C1371 VDD.n1185 GND 0.00558f
C1372 VDD.n1186 GND 0.006932f
C1373 VDD.n1187 GND 0.331657f
C1374 VDD.n1188 GND 0.006932f
C1375 VDD.n1189 GND 0.00558f
C1376 VDD.n1190 GND 0.006932f
C1377 VDD.n1191 GND 0.00558f
C1378 VDD.n1192 GND 0.006932f
C1379 VDD.n1193 GND 0.372649f
C1380 VDD.t117 GND 0.186324f
C1381 VDD.n1194 GND 0.006932f
C1382 VDD.n1195 GND 0.00558f
C1383 VDD.n1196 GND 0.006932f
C1384 VDD.n1197 GND 0.00558f
C1385 VDD.n1198 GND 0.006932f
C1386 VDD.n1199 GND 0.372649f
C1387 VDD.n1200 GND 0.006932f
C1388 VDD.n1201 GND 0.00558f
C1389 VDD.n1202 GND 0.006932f
C1390 VDD.n1203 GND 0.00558f
C1391 VDD.n1204 GND 0.006932f
C1392 VDD.n1205 GND 0.372649f
C1393 VDD.n1206 GND 0.006932f
C1394 VDD.n1207 GND 0.00558f
C1395 VDD.n1208 GND 0.006932f
C1396 VDD.n1209 GND 0.00558f
C1397 VDD.n1210 GND 0.006932f
C1398 VDD.n1211 GND 0.372649f
C1399 VDD.n1212 GND 0.006932f
C1400 VDD.n1213 GND 0.00558f
C1401 VDD.n1214 GND 0.006932f
C1402 VDD.n1215 GND 0.00558f
C1403 VDD.n1216 GND 0.006932f
C1404 VDD.t74 GND 0.186324f
C1405 VDD.n1217 GND 0.006932f
C1406 VDD.n1218 GND 0.00558f
C1407 VDD.n1219 GND 0.006932f
C1408 VDD.n1220 GND 0.00558f
C1409 VDD.n1221 GND 0.006932f
C1410 VDD.n1222 GND 0.372649f
C1411 VDD.n1223 GND 0.006932f
C1412 VDD.n1224 GND 0.00558f
C1413 VDD.n1225 GND 0.016092f
C1414 VDD.n1226 GND 0.016092f
C1415 VDD.n1227 GND 0.834733f
C1416 VDD.n1228 GND 0.016092f
C1417 VDD.n1229 GND 0.006932f
C1418 VDD.n1231 GND 0.006932f
C1419 VDD.n1232 GND 0.006932f
C1420 VDD.n1233 GND 0.00558f
C1421 VDD.n1234 GND 0.006932f
C1422 VDD.n1235 GND 0.006932f
C1423 VDD.n1237 GND 0.006932f
C1424 VDD.n1238 GND 0.006932f
C1425 VDD.n1239 GND 0.004715f
C1426 VDD.n1240 GND 0.006932f
C1427 VDD.n1241 GND 0.006932f
C1428 VDD.n1242 GND 0.00558f
C1429 VDD.n1243 GND 0.006932f
C1430 VDD.n1244 GND 0.006932f
C1431 VDD.n1246 GND 0.006932f
C1432 VDD.n1247 GND 0.006932f
C1433 VDD.n1249 GND 0.006932f
C1434 VDD.n1250 GND 0.00558f
C1435 VDD.n1251 GND 0.006932f
C1436 VDD.n1252 GND 0.006932f
C1437 VDD.n1254 GND 0.006932f
C1438 VDD.n1255 GND 0.005496f
C1439 VDD.n1257 GND 0.00558f
C1440 VDD.n1258 GND 0.006932f
C1441 VDD.n1259 GND 0.006932f
C1442 VDD.n1260 GND 0.006932f
C1443 VDD.n1261 GND 0.006932f
C1444 VDD.n1263 GND 0.006932f
C1445 VDD.n1264 GND 0.006932f
C1446 VDD.n1265 GND 0.00558f
C1447 VDD.n1267 GND 0.006932f
C1448 VDD.n1269 GND 0.006932f
C1449 VDD.n1270 GND 0.002539f
C1450 VDD.t75 GND 0.030733f
C1451 VDD.t76 GND 0.039858f
C1452 VDD.t73 GND 0.203294f
C1453 VDD.n1271 GND 0.050408f
C1454 VDD.n1272 GND 0.037394f
C1455 VDD.n1273 GND 0.008593f
C1456 VDD.n1274 GND 0.003041f
C1457 VDD.n1275 GND 0.006932f
C1458 VDD.n1276 GND 0.006932f
C1459 VDD.n1277 GND 0.006932f
C1460 VDD.n1278 GND 0.00558f
C1461 VDD.n1279 GND 0.00558f
C1462 VDD.n1280 GND 0.00558f
C1463 VDD.n1281 GND 0.006932f
C1464 VDD.n1282 GND 0.006932f
C1465 VDD.n1283 GND 0.006932f
C1466 VDD.n1284 GND 0.00558f
C1467 VDD.n1285 GND 0.006932f
C1468 VDD.n1286 GND 0.006932f
C1469 VDD.n1288 GND 0.006932f
C1470 VDD.t84 GND 0.030733f
C1471 VDD.t85 GND 0.039858f
C1472 VDD.t83 GND 0.203294f
C1473 VDD.n1289 GND 0.050408f
C1474 VDD.n1290 GND 0.037394f
C1475 VDD.n1291 GND 0.011382f
C1476 VDD.n1292 GND 0.003822f
C1477 VDD.n1293 GND 0.006932f
C1478 VDD.n1294 GND 0.006932f
C1479 VDD.n1295 GND 0.006932f
C1480 VDD.n1296 GND 0.00558f
C1481 VDD.n1297 GND 0.00558f
C1482 VDD.n1298 GND 0.00558f
C1483 VDD.n1299 GND 0.006932f
C1484 VDD.n1300 GND 0.006932f
C1485 VDD.n1301 GND 0.006932f
C1486 VDD.n1302 GND 0.00558f
C1487 VDD.n1303 GND 0.006932f
C1488 VDD.n1305 GND 0.006932f
C1489 VDD.n1307 GND 0.006932f
C1490 VDD.t81 GND 0.030733f
C1491 VDD.t82 GND 0.039858f
C1492 VDD.t80 GND 0.203294f
C1493 VDD.n1308 GND 0.050408f
C1494 VDD.n1309 GND 0.037394f
C1495 VDD.n1310 GND 0.011382f
C1496 VDD.n1311 GND 0.004603f
C1497 VDD.n1312 GND 0.00558f
C1498 VDD.n1313 GND 0.006932f
C1499 VDD.n1314 GND 0.006932f
C1500 VDD.n1315 GND 0.006932f
C1501 VDD.n1316 GND 0.00558f
C1502 VDD.n1317 GND 0.00558f
C1503 VDD.n1318 GND 0.004631f
C1504 VDD.n1319 GND 0.016092f
C1505 VDD.n1320 GND 0.016004f
C1506 VDD.n1321 GND 0.004631f
C1507 VDD.n1322 GND 0.016004f
C1508 VDD.n1323 GND 0.495623f
C1509 VDD.n1324 GND 0.016004f
C1510 VDD.n1325 GND 0.004631f
C1511 VDD.n1326 GND 0.016004f
C1512 VDD.n1327 GND 0.006932f
C1513 VDD.n1328 GND 0.006932f
C1514 VDD.n1329 GND 0.00558f
C1515 VDD.n1330 GND 0.006932f
C1516 VDD.n1331 GND 0.283213f
C1517 VDD.n1332 GND 0.372649f
C1518 VDD.n1333 GND 0.006932f
C1519 VDD.n1334 GND 0.00558f
C1520 VDD.n1335 GND 0.006932f
C1521 VDD.n1336 GND 0.006932f
C1522 VDD.n1337 GND 0.006932f
C1523 VDD.n1338 GND 0.00558f
C1524 VDD.n1339 GND 0.006932f
C1525 VDD.n1340 GND 0.27576f
C1526 VDD.n1341 GND 0.006932f
C1527 VDD.n1342 GND 0.00558f
C1528 VDD.n1343 GND 0.006932f
C1529 VDD.n1344 GND 0.006932f
C1530 VDD.n1345 GND 0.006932f
C1531 VDD.n1346 GND 0.00558f
C1532 VDD.n1347 GND 0.006932f
C1533 VDD.n1348 GND 0.372649f
C1534 VDD.n1349 GND 0.006932f
C1535 VDD.n1350 GND 0.00558f
C1536 VDD.n1351 GND 0.006932f
C1537 VDD.n1352 GND 0.006932f
C1538 VDD.n1353 GND 0.006932f
C1539 VDD.n1354 GND 0.00558f
C1540 VDD.n1355 GND 0.006932f
C1541 VDD.n1356 GND 0.372649f
C1542 VDD.n1357 GND 0.006932f
C1543 VDD.n1358 GND 0.00558f
C1544 VDD.n1359 GND 0.006932f
C1545 VDD.n1360 GND 0.006932f
C1546 VDD.n1361 GND 0.006932f
C1547 VDD.n1362 GND 0.00558f
C1548 VDD.n1363 GND 0.006932f
C1549 VDD.n1364 GND 0.372649f
C1550 VDD.n1365 GND 0.006932f
C1551 VDD.n1366 GND 0.00558f
C1552 VDD.n1367 GND 0.006932f
C1553 VDD.n1368 GND 0.006932f
C1554 VDD.n1369 GND 0.006932f
C1555 VDD.n1370 GND 0.00558f
C1556 VDD.n1371 GND 0.006932f
C1557 VDD.n1372 GND 0.227316f
C1558 VDD.n1373 GND 0.006932f
C1559 VDD.n1374 GND 0.00558f
C1560 VDD.n1375 GND 0.006932f
C1561 VDD.n1376 GND 0.006932f
C1562 VDD.n1377 GND 0.006932f
C1563 VDD.n1378 GND 0.00558f
C1564 VDD.n1379 GND 0.006932f
C1565 VDD.n1380 GND 0.372649f
C1566 VDD.n1381 GND 0.006932f
C1567 VDD.n1382 GND 0.00558f
C1568 VDD.n1383 GND 0.006932f
C1569 VDD.n1384 GND 0.006932f
C1570 VDD.n1385 GND 0.006932f
C1571 VDD.n1386 GND 0.00558f
C1572 VDD.n1387 GND 0.006932f
C1573 VDD.n1388 GND 0.372649f
C1574 VDD.n1389 GND 0.006932f
C1575 VDD.n1390 GND 0.00558f
C1576 VDD.n1391 GND 0.006932f
C1577 VDD.n1392 GND 0.006932f
C1578 VDD.n1393 GND 0.006932f
C1579 VDD.n1394 GND 0.00558f
C1580 VDD.n1395 GND 0.006932f
C1581 VDD.t114 GND 0.186324f
C1582 VDD.n1396 GND 0.324204f
C1583 VDD.n1397 GND 0.006932f
C1584 VDD.n1398 GND 0.00558f
C1585 VDD.n1399 GND 0.006932f
C1586 VDD.n1400 GND 0.006932f
C1587 VDD.n1401 GND 0.006932f
C1588 VDD.n1402 GND 0.00558f
C1589 VDD.n1403 GND 0.006932f
C1590 VDD.n1404 GND 0.372649f
C1591 VDD.n1405 GND 0.006932f
C1592 VDD.n1406 GND 0.00558f
C1593 VDD.n1407 GND 0.006932f
C1594 VDD.n1408 GND 0.006932f
C1595 VDD.n1409 GND 0.006932f
C1596 VDD.n1410 GND 0.00558f
C1597 VDD.n1411 GND 0.006932f
C1598 VDD.n1412 GND 0.372649f
C1599 VDD.n1413 GND 0.006932f
C1600 VDD.n1414 GND 0.00558f
C1601 VDD.t129 GND 0.036671f
C1602 VDD.t115 GND 0.005831f
C1603 VDD.t133 GND 0.005831f
C1604 VDD.n1415 GND 0.022552f
C1605 VDD.n1416 GND 0.173338f
C1606 VDD.t118 GND 0.035481f
C1607 VDD.n1417 GND 0.092021f
C1608 VDD.t135 GND 0.036671f
C1609 VDD.t119 GND 0.005831f
C1610 VDD.t107 GND 0.005831f
C1611 VDD.n1418 GND 0.022552f
C1612 VDD.n1419 GND 0.173338f
C1613 VDD.t121 GND 0.035481f
C1614 VDD.n1420 GND 0.084902f
C1615 VDD.n1421 GND 0.064618f
C1616 VDD.t131 GND 0.036671f
C1617 VDD.t116 GND 0.005831f
C1618 VDD.t136 GND 0.005831f
C1619 VDD.n1422 GND 0.022552f
C1620 VDD.n1423 GND 0.173338f
C1621 VDD.t120 GND 0.035481f
C1622 VDD.n1424 GND 0.084902f
C1623 VDD.n1425 GND 0.123752f
C1624 VDD.n1426 GND 2.7946f
C1625 VDD.n1427 GND 0.397993f
C1626 VDD.n1428 GND 0.006908f
C1627 VDD.n1429 GND 0.006932f
C1628 VDD.n1430 GND 0.00558f
C1629 VDD.n1431 GND 0.006932f
C1630 VDD.n1432 GND 0.372649f
C1631 VDD.n1433 GND 0.006932f
C1632 VDD.n1434 GND 0.00558f
C1633 VDD.n1435 GND 0.006932f
C1634 VDD.n1436 GND 0.006932f
C1635 VDD.n1437 GND 0.006932f
C1636 VDD.n1438 GND 0.00558f
C1637 VDD.n1439 GND 0.006932f
C1638 VDD.n1440 GND 0.324204f
C1639 VDD.n1441 GND 0.006932f
C1640 VDD.n1442 GND 0.00558f
C1641 VDD.n1443 GND 0.006932f
C1642 VDD.n1444 GND 0.006932f
C1643 VDD.n1445 GND 0.006932f
C1644 VDD.n1446 GND 0.00558f
C1645 VDD.n1447 GND 0.006932f
C1646 VDD.n1448 GND 0.372649f
C1647 VDD.n1449 GND 0.006932f
C1648 VDD.n1450 GND 0.00558f
C1649 VDD.n1451 GND 0.006932f
C1650 VDD.n1452 GND 0.006932f
C1651 VDD.n1453 GND 0.006932f
C1652 VDD.n1454 GND 0.00558f
C1653 VDD.n1455 GND 0.006932f
C1654 VDD.n1456 GND 0.331657f
C1655 VDD.n1457 GND 0.372649f
C1656 VDD.n1458 GND 0.006932f
C1657 VDD.n1459 GND 0.00558f
C1658 VDD.n1460 GND 0.006932f
C1659 VDD.n1461 GND 0.006932f
C1660 VDD.n1462 GND 0.006932f
C1661 VDD.n1463 GND 0.00558f
C1662 VDD.n1464 GND 0.006932f
C1663 VDD.n1465 GND 0.227316f
C1664 VDD.n1466 GND 0.006932f
C1665 VDD.n1467 GND 0.00558f
C1666 VDD.n1468 GND 0.006932f
C1667 VDD.n1469 GND 0.006932f
C1668 VDD.n1470 GND 0.006932f
C1669 VDD.n1471 GND 0.00558f
C1670 VDD.n1472 GND 0.006932f
C1671 VDD.n1473 GND 0.372649f
C1672 VDD.n1474 GND 0.006932f
C1673 VDD.n1475 GND 0.00558f
C1674 VDD.n1476 GND 0.006932f
C1675 VDD.n1477 GND 0.006932f
C1676 VDD.n1478 GND 0.006932f
C1677 VDD.n1479 GND 0.00558f
C1678 VDD.n1480 GND 0.006932f
C1679 VDD.n1481 GND 0.372649f
C1680 VDD.n1482 GND 0.006932f
C1681 VDD.n1483 GND 0.00558f
C1682 VDD.n1484 GND 0.006932f
C1683 VDD.n1485 GND 0.006932f
C1684 VDD.n1486 GND 0.006932f
C1685 VDD.n1487 GND 0.006932f
C1686 VDD.n1488 GND 0.00558f
C1687 VDD.n1489 GND 0.006932f
C1688 VDD.n1490 GND 0.372649f
C1689 VDD.n1491 GND 0.006932f
C1690 VDD.n1492 GND 0.00558f
C1691 VDD.n1493 GND 0.006932f
C1692 VDD.n1494 GND 0.006932f
C1693 VDD.n1495 GND 0.006932f
C1694 VDD.n1496 GND 0.00558f
C1695 VDD.n1497 GND 0.006932f
C1696 VDD.n1498 GND 0.27576f
C1697 VDD.n1499 GND 0.006932f
C1698 VDD.n1500 GND 0.006932f
C1699 VDD.n1501 GND 0.00558f
C1700 VDD.n1502 GND 0.006932f
C1701 VDD.n1503 GND 0.006932f
C1702 VDD.n1504 GND 0.007799f
C1703 VDD.n1505 GND 0.006932f
C1704 VDD.n1506 GND 0.00558f
C1705 VDD.n1507 GND 0.006932f
C1706 VDD.n1508 GND 0.372649f
C1707 VDD.n1509 GND 0.372649f
C1708 VDD.n1510 GND 0.006932f
C1709 VDD.n1511 GND 0.00558f
C1710 VDD.n1512 GND 0.006932f
C1711 VDD.n1513 GND 0.006932f
C1712 VDD.n1514 GND 0.011479f
C1713 VDD.n1515 GND 0.004631f
C1714 VDD.n1516 GND 0.016004f
C1715 VDD.n1517 GND 0.016092f
C1716 VDD.n1518 GND 0.004631f
C1717 VDD.n1519 GND 0.003934f
C1718 VDD.n1520 GND 0.003466f
C1719 VDD.n1521 GND 0.003466f
C1720 VDD.n1522 GND 0.00558f
C1721 VDD.n1523 GND 0.00558f
C1722 VDD.n1524 GND 0.006932f
C1723 VDD.n1525 GND 0.006932f
C1724 VDD.n1526 GND 0.00558f
C1725 VDD.n1527 GND 0.003466f
C1726 VDD.n1528 GND 0.003466f
C1727 VDD.n1529 GND 0.003466f
C1728 VDD.n1530 GND 0.006932f
C1729 VDD.n1531 GND 0.006932f
C1730 VDD.n1532 GND 0.011382f
C1731 VDD.n1533 GND 0.004715f
C1732 VDD.n1534 GND 0.006932f
C1733 VDD.n1535 GND 0.006932f
C1734 VDD.n1536 GND 0.00558f
C1735 VDD.n1537 GND 0.003466f
C1736 VDD.n1538 GND 0.003466f
C1737 VDD.n1539 GND 0.003466f
C1738 VDD.n1540 GND 0.00558f
C1739 VDD.n1541 GND 0.006932f
C1740 VDD.n1542 GND 0.006932f
C1741 VDD.n1545 GND 0.006932f
C1742 VDD.n1548 GND 0.006932f
C1743 VDD.t18 GND 3.20478f
C1744 VDD.t31 GND 4.24074f
C1745 VDD.t29 GND 4.24074f
C1746 VDD.t36 GND 4.64693f
C1747 VDD.t0 GND 5.15746f
C1748 VDD.n1552 GND 2.9402f
C1749 VDD.n1553 GND 0.016092f
C1750 VDD.n1554 GND 0.002539f
C1751 VDD.n1555 GND 0.005147f
C1752 VDD.n1556 GND 0.003466f
C1753 VDD.n1557 GND 0.003466f
C1754 VDD.n1558 GND 0.00558f
C1755 VDD.n1559 GND 0.00558f
C1756 VDD.n1560 GND 0.00558f
C1757 VDD.n1561 GND 0.003466f
C1758 VDD.n1562 GND 0.003466f
C1759 VDD.n1563 GND 0.003466f
C1760 VDD.n1564 GND 0.00558f
C1761 VDD.n1565 GND 0.00558f
C1762 VDD.n1566 GND 0.005496f
C1763 VDD.n1567 GND 0.003466f
C1764 VDD.n1568 GND 0.003466f
C1765 VDD.n1569 GND 0.003466f
C1766 VDD.n1570 GND 0.003822f
C1767 VDD.n1571 GND 0.00558f
C1768 VDD.n1572 GND 0.00558f
C1769 VDD.n1573 GND 0.045614f
C1770 VDD.n1574 GND 2.08151f
C1771 VDD.n1575 GND 0.211802f
C1772 VDD.n1576 GND 0.003535f
C1773 VDD.n1577 GND 0.004714f
C1774 VDD.n1578 GND 0.004714f
C1775 VDD.n1580 GND 0.004714f
C1776 VDD.n1581 GND 0.004714f
C1777 VDD.n1582 GND 0.004714f
C1778 VDD.n1583 GND 0.004714f
C1779 VDD.n1584 GND 0.004714f
C1780 VDD.n1585 GND 0.004714f
C1781 VDD.n1587 GND 0.004714f
C1782 VDD.n1588 GND 0.004714f
C1783 VDD.n1589 GND 0.012357f
C1784 VDD.n1590 GND 0.011836f
C1785 VDD.n1591 GND 0.011836f
C1786 VDD.n1592 GND 0.391281f
C1787 VDD.n1593 GND 0.011836f
C1788 VDD.n1594 GND 0.011836f
C1789 VDD.n1595 GND 0.004714f
C1790 VDD.n1596 GND 0.004714f
C1791 VDD.n1597 GND 0.004714f
C1792 VDD.n1598 GND 0.253401f
C1793 VDD.n1599 GND 0.004714f
C1794 VDD.n1600 GND 0.004714f
C1795 VDD.n1601 GND 0.004714f
C1796 VDD.n1602 GND 0.004714f
C1797 VDD.n1603 GND 0.004714f
C1798 VDD.n1604 GND 0.253401f
C1799 VDD.n1605 GND 0.004714f
C1800 VDD.n1606 GND 0.004714f
C1801 VDD.n1607 GND 0.004714f
C1802 VDD.n1608 GND 0.004714f
C1803 VDD.n1609 GND 0.004714f
C1804 VDD.n1610 GND 0.253401f
C1805 VDD.n1611 GND 0.004714f
C1806 VDD.n1612 GND 0.004714f
C1807 VDD.n1613 GND 0.004714f
C1808 VDD.n1614 GND 0.004714f
C1809 VDD.n1615 GND 0.004714f
C1810 VDD.n1616 GND 0.253401f
C1811 VDD.n1617 GND 0.004714f
C1812 VDD.n1618 GND 0.004714f
C1813 VDD.n1619 GND 0.004714f
C1814 VDD.n1620 GND 0.004714f
C1815 VDD.n1621 GND 0.004714f
C1816 VDD.n1622 GND 0.229179f
C1817 VDD.n1623 GND 0.004714f
C1818 VDD.n1624 GND 0.004714f
C1819 VDD.n1625 GND 0.004714f
C1820 VDD.n1626 GND 0.004714f
C1821 VDD.n1627 GND 0.004714f
C1822 VDD.n1628 GND 0.253401f
C1823 VDD.n1629 GND 0.004714f
C1824 VDD.n1630 GND 0.004714f
C1825 VDD.n1631 GND 0.004714f
C1826 VDD.n1632 GND 0.004714f
C1827 VDD.n1633 GND 0.004714f
C1828 VDD.n1634 GND 0.20123f
C1829 VDD.n1635 GND 0.004714f
C1830 VDD.n1636 GND 0.004714f
C1831 VDD.n1637 GND 0.004714f
C1832 VDD.n1638 GND 0.004714f
C1833 VDD.n1639 GND 0.004714f
C1834 VDD.n1640 GND 0.253401f
C1835 VDD.n1641 GND 0.004714f
C1836 VDD.n1642 GND 0.004714f
C1837 VDD.n1643 GND 0.004714f
C1838 VDD.n1644 GND 0.004714f
C1839 VDD.n1645 GND 0.004714f
C1840 VDD.n1646 GND 0.253401f
C1841 VDD.n1647 GND 0.004714f
C1842 VDD.n1648 GND 0.004714f
C1843 VDD.n1649 GND 0.004714f
C1844 VDD.n1650 GND 0.004714f
C1845 VDD.n1651 GND 0.004714f
C1846 VDD.n1652 GND 0.253401f
C1847 VDD.n1653 GND 0.004714f
C1848 VDD.n1654 GND 0.004714f
C1849 VDD.n1655 GND 0.004714f
C1850 VDD.n1656 GND 0.004714f
C1851 VDD.n1657 GND 0.004714f
C1852 VDD.n1658 GND 0.253401f
C1853 VDD.n1659 GND 0.004714f
C1854 VDD.n1660 GND 0.004714f
C1855 VDD.n1661 GND 0.004714f
C1856 VDD.n1662 GND 0.004714f
C1857 VDD.n1663 GND 0.004714f
C1858 VDD.n1664 GND 0.253401f
C1859 VDD.n1665 GND 0.004714f
C1860 VDD.n1666 GND 0.004714f
C1861 VDD.n1667 GND 0.004714f
C1862 VDD.n1668 GND 0.004714f
C1863 VDD.n1669 GND 0.004714f
C1864 VDD.n1670 GND 0.253401f
C1865 VDD.n1671 GND 0.004714f
C1866 VDD.n1672 GND 0.004714f
C1867 VDD.n1673 GND 0.004714f
C1868 VDD.n1674 GND 0.004714f
C1869 VDD.n1675 GND 0.004714f
C1870 VDD.n1676 GND 0.253401f
C1871 VDD.n1677 GND 0.004714f
C1872 VDD.n1678 GND 0.004714f
C1873 VDD.n1679 GND 0.004714f
C1874 VDD.n1680 GND 0.004714f
C1875 VDD.n1681 GND 0.004714f
C1876 VDD.n1682 GND 0.236632f
C1877 VDD.n1683 GND 0.004714f
C1878 VDD.n1684 GND 0.004714f
C1879 VDD.n1685 GND 0.004714f
C1880 VDD.n1686 GND 0.004714f
C1881 VDD.n1687 GND 0.004714f
C1882 VDD.n1688 GND 0.21241f
C1883 VDD.n1689 GND 0.004714f
C1884 VDD.n1690 GND 0.004714f
C1885 VDD.n1691 GND 0.004714f
C1886 VDD.n1692 GND 0.004714f
C1887 VDD.n1693 GND 0.004714f
C1888 VDD.n1694 GND 0.253401f
C1889 VDD.n1695 GND 0.004714f
C1890 VDD.n1696 GND 0.004714f
C1891 VDD.n1697 GND 0.004714f
C1892 VDD.n1698 GND 0.004714f
C1893 VDD.n1699 GND 0.004714f
C1894 VDD.n1700 GND 0.253401f
C1895 VDD.n1701 GND 0.004714f
C1896 VDD.n1702 GND 0.004714f
C1897 VDD.n1703 GND 0.004714f
C1898 VDD.n1704 GND 0.004714f
C1899 VDD.n1705 GND 0.004714f
C1900 VDD.n1706 GND 0.253401f
C1901 VDD.n1707 GND 0.004714f
C1902 VDD.n1708 GND 0.004714f
C1903 VDD.n1709 GND 0.004714f
C1904 VDD.n1710 GND 0.004714f
C1905 VDD.n1711 GND 0.004714f
C1906 VDD.n1712 GND 0.253401f
C1907 VDD.n1713 GND 0.004714f
C1908 VDD.n1714 GND 0.004714f
C1909 VDD.n1715 GND 0.004714f
C1910 VDD.n1716 GND 0.004714f
C1911 VDD.n1717 GND 0.004714f
C1912 VDD.n1718 GND 0.253401f
C1913 VDD.n1719 GND 0.004714f
C1914 VDD.n1720 GND 0.004714f
C1915 VDD.n1721 GND 0.004714f
C1916 VDD.n1722 GND 0.004714f
C1917 VDD.n1723 GND 0.004714f
C1918 VDD.n1724 GND 0.253401f
C1919 VDD.n1725 GND 0.004714f
C1920 VDD.n1726 GND 0.004714f
C1921 VDD.n1727 GND 0.004714f
C1922 VDD.n1728 GND 0.004714f
C1923 VDD.n1729 GND 0.004714f
C1924 VDD.n1730 GND 0.14347f
C1925 VDD.n1731 GND 0.004714f
C1926 VDD.n1732 GND 0.004714f
C1927 VDD.n1733 GND 0.004714f
C1928 VDD.n1734 GND 0.004714f
C1929 VDD.n1735 GND 0.004714f
C1930 VDD.n1736 GND 0.134154f
C1931 VDD.n1737 GND 0.004714f
C1932 VDD.n1738 GND 0.004714f
C1933 VDD.n1739 GND 0.004714f
C1934 VDD.n1740 GND 0.004714f
C1935 VDD.n1741 GND 0.004714f
C1936 VDD.n1742 GND 0.253401f
C1937 VDD.n1743 GND 0.004714f
C1938 VDD.n1744 GND 0.004714f
C1939 VDD.n1745 GND 0.004714f
C1940 VDD.n1746 GND 0.004714f
C1941 VDD.n1747 GND 0.004714f
C1942 VDD.n1748 GND 0.253401f
C1943 VDD.n1749 GND 0.004714f
C1944 VDD.n1750 GND 0.004714f
C1945 VDD.n1751 GND 0.004714f
C1946 VDD.n1752 GND 0.004714f
C1947 VDD.n1753 GND 0.004714f
C1948 VDD.n1754 GND 0.253401f
C1949 VDD.n1755 GND 0.004714f
C1950 VDD.n1756 GND 0.004714f
C1951 VDD.n1757 GND 0.004714f
C1952 VDD.n1758 GND 0.004714f
C1953 VDD.n1759 GND 0.004714f
C1954 VDD.n1760 GND 0.253401f
C1955 VDD.n1761 GND 0.004714f
C1956 VDD.n1762 GND 0.004714f
C1957 VDD.n1763 GND 0.004714f
C1958 VDD.n1764 GND 0.004714f
C1959 VDD.n1765 GND 0.004714f
C1960 VDD.n1766 GND 0.253401f
C1961 VDD.n1767 GND 0.004714f
C1962 VDD.n1768 GND 0.004714f
C1963 VDD.n1769 GND 0.004714f
C1964 VDD.n1770 GND 0.004714f
C1965 VDD.n1771 GND 0.004714f
C1966 VDD.n1772 GND 0.253401f
C1967 VDD.n1773 GND 0.004714f
C1968 VDD.n1774 GND 0.004714f
C1969 VDD.n1775 GND 0.004714f
C1970 VDD.n1776 GND 0.004714f
C1971 VDD.n1777 GND 0.004714f
C1972 VDD.n1778 GND 0.253401f
C1973 VDD.n1779 GND 0.004714f
C1974 VDD.n1780 GND 0.004714f
C1975 VDD.n1781 GND 0.004714f
C1976 VDD.n1782 GND 0.004714f
C1977 VDD.n1783 GND 0.004714f
C1978 VDD.n1784 GND 0.227316f
C1979 VDD.n1785 GND 0.004714f
C1980 VDD.n1786 GND 0.004714f
C1981 VDD.n1787 GND 0.004714f
C1982 VDD.n1788 GND 0.004714f
C1983 VDD.n1789 GND 0.004714f
C1984 VDD.n1790 GND 0.150923f
C1985 VDD.n1791 GND 0.004714f
C1986 VDD.n1792 GND 0.004714f
C1987 VDD.n1793 GND 0.004714f
C1988 VDD.n1794 GND 0.004714f
C1989 VDD.n1795 GND 0.004714f
C1990 VDD.n1796 GND 0.253401f
C1991 VDD.n1797 GND 0.004714f
C1992 VDD.n1798 GND 0.004714f
C1993 VDD.n1799 GND 0.004714f
C1994 VDD.t52 GND 0.03345f
C1995 VDD.t51 GND 0.055799f
C1996 VDD.t49 GND 0.595646f
C1997 VDD.n1800 GND 0.093248f
C1998 VDD.n1801 GND 0.071157f
C1999 VDD.n1802 GND 0.006737f
C2000 VDD.n1803 GND 0.004714f
C2001 VDD.n1804 GND 0.003882f
C2002 VDD.n1805 GND 0.004714f
C2003 VDD.n1806 GND 0.004714f
C2004 VDD.n1807 GND 0.004714f
C2005 VDD.n1808 GND 0.004714f
C2006 VDD.n1809 GND 0.004714f
C2007 VDD.n1810 GND 0.004714f
C2008 VDD.n1811 GND 0.004714f
C2009 VDD.n1812 GND 0.004714f
C2010 VDD.n1813 GND 0.004714f
C2011 VDD.n1814 GND 0.004714f
C2012 VDD.n1815 GND 0.004714f
C2013 VDD.n1816 GND 0.004714f
C2014 VDD.n1817 GND 0.004714f
C2015 VDD.n1818 GND 0.004714f
C2016 VDD.n1819 GND 0.004714f
C2017 VDD.n1820 GND 0.004714f
C2018 VDD.n1821 GND 0.004714f
C2019 VDD.n1822 GND 0.004714f
C2020 VDD.n1823 GND 0.004714f
C2021 VDD.n1824 GND 0.004714f
C2022 VDD.n1825 GND 0.004714f
C2023 VDD.n1826 GND 0.004714f
C2024 VDD.n1827 GND 0.004714f
C2025 VDD.n1828 GND 0.004714f
C2026 VDD.n1829 GND 0.012357f
C2027 VDD.n1830 GND 0.012357f
C2028 VDD.n1831 GND 0.011836f
C2029 VDD.n1832 GND 0.011836f
C2030 VDD.n1833 GND 0.004714f
C2031 VDD.n1834 GND 0.004714f
C2032 VDD.n1835 GND 0.004714f
C2033 VDD.n1836 GND 0.004714f
C2034 VDD.n1837 GND 0.004714f
C2035 VDD.n1838 GND 0.004714f
C2036 VDD.n1839 GND 0.004714f
C2037 VDD.n1840 GND 0.253401f
C2038 VDD.n1841 GND 0.004714f
C2039 VDD.n1842 GND 0.004714f
C2040 VDD.n1843 GND 0.004714f
C2041 VDD.n1844 GND 0.004714f
C2042 VDD.n1845 GND 0.004714f
C2043 VDD.n1846 GND 0.253401f
C2044 VDD.n1847 GND 0.004714f
C2045 VDD.n1848 GND 0.004714f
C2046 VDD.n1849 GND 0.004714f
C2047 VDD.n1850 GND 0.004714f
C2048 VDD.n1851 GND 0.012322f
C2049 VDD.n1852 GND 0.011836f
C2050 VDD.n1853 GND 0.012357f
C2051 VDD.n1854 GND 0.011872f
C2052 VDD.n1855 GND 0.003189f
C2053 VDD.n1856 GND 0.004714f
C2054 VDD.n1857 GND 0.004714f
C2055 VDD.n1858 GND 0.003882f
C2056 VDD.n1859 GND 0.004714f
C2057 VDD.n1860 GND 0.004714f
C2058 VDD.n1861 GND 0.004714f
C2059 VDD.n1862 GND 0.004714f
C2060 VDD.n1863 GND 0.004714f
C2061 VDD.n1864 GND 0.004714f
C2062 VDD.n1865 GND 0.004714f
C2063 VDD.n1866 GND 0.004714f
C2064 VDD.n1867 GND 0.004714f
C2065 VDD.n1868 GND 0.004714f
C2066 VDD.n1869 GND 0.004714f
C2067 VDD.n1870 GND 0.004714f
C2068 VDD.n1871 GND 0.004714f
C2069 VDD.n1872 GND 0.004714f
C2070 VDD.n1873 GND 0.004714f
C2071 VDD.n1874 GND 0.004714f
C2072 VDD.n1875 GND 0.004714f
C2073 VDD.n1876 GND 0.004714f
C2074 VDD.n1877 GND 0.004714f
C2075 VDD.n1878 GND 0.004714f
C2076 VDD.n1879 GND 0.004714f
C2077 VDD.n1880 GND 0.004714f
C2078 VDD.n1881 GND 0.004714f
C2079 VDD.n1882 GND 0.004714f
C2080 VDD.n1883 GND 0.012357f
C2081 VDD.n1884 GND 0.012357f
C2082 VDD.n1885 GND 0.011836f
C2083 VDD.n1886 GND 0.004714f
C2084 VDD.n1887 GND 0.004714f
C2085 VDD.n1888 GND 0.253401f
C2086 VDD.n1889 GND 0.004714f
C2087 VDD.n1890 GND 0.004714f
C2088 VDD.n1891 GND 0.012322f
C2089 VDD.n1892 GND 0.011872f
C2090 VDD.n1893 GND 0.012357f
C2091 VDD.n1895 GND 1.6173f
C2092 VDD.n1896 GND 1.6173f
C2093 VDD.n1897 GND 0.011836f
C2094 VDD.n1898 GND 0.012357f
C2095 VDD.n1899 GND 0.004714f
C2096 VDD.t65 GND 0.03345f
C2097 VDD.t66 GND 0.055799f
C2098 VDD.t64 GND 0.595646f
C2099 VDD.n1900 GND 0.093248f
C2100 VDD.n1901 GND 0.071157f
C2101 VDD.n1902 GND 0.006737f
C2102 VDD.n1903 GND 0.003882f
C2103 VDD.n1904 GND 0.004714f
C2104 VDD.n1905 GND 0.004714f
C2105 VDD.n1906 GND 0.004714f
C2106 VDD.n1907 GND 0.004714f
C2107 VDD.n1908 GND 0.004714f
C2108 VDD.n1909 GND 0.004714f
C2109 VDD.n1911 GND 0.004714f
C2110 VDD.n1913 GND 0.004714f
C2111 VDD.n1914 GND 0.004714f
C2112 VDD.n1915 GND 0.004714f
C2113 VDD.n1916 GND 0.004714f
C2114 VDD.n1917 GND 0.004714f
C2115 VDD.n1919 GND 0.004714f
C2116 VDD.n1921 GND 0.004714f
C2117 VDD.n1922 GND 0.004714f
C2118 VDD.n1923 GND 0.004714f
C2119 VDD.n1924 GND 0.004714f
C2120 VDD.n1925 GND 0.004714f
C2121 VDD.n1927 GND 0.004714f
C2122 VDD.n1929 GND 0.004714f
C2123 VDD.n1930 GND 0.004714f
C2124 VDD.n1931 GND 0.004714f
C2125 VDD.n1932 GND 0.004714f
C2126 VDD.n1933 GND 0.004714f
C2127 VDD.n1935 GND 0.004714f
C2128 VDD.n1937 GND 0.004714f
C2129 VDD.n1938 GND 0.003189f
C2130 VDD.n1939 GND 0.012357f
C2131 VDD.n1940 GND 0.004714f
C2132 VDD.n1941 GND 0.004714f
C2133 VDD.n1942 GND 0.004714f
C2134 VDD.n1943 GND 0.004714f
C2135 VDD.n1944 GND 0.004714f
C2136 VDD.n1945 GND 0.004714f
C2137 VDD.n1946 GND 0.004714f
C2138 VDD.n1947 GND 0.004714f
C2139 VDD.n1948 GND 0.004714f
C2140 VDD.n1949 GND 0.004714f
C2141 VDD.n1950 GND 0.004714f
C2142 VDD.n1951 GND 0.004714f
C2143 VDD.n1952 GND 0.004714f
C2144 VDD.n1953 GND 0.004714f
C2145 VDD.n1954 GND 0.004714f
C2146 VDD.n1955 GND 0.004714f
C2147 VDD.n1956 GND 0.004714f
C2148 VDD.n1957 GND 0.004714f
C2149 VDD.n1958 GND 0.004714f
C2150 VDD.n1959 GND 0.004714f
C2151 VDD.n1960 GND 0.004714f
C2152 VDD.n1961 GND 0.004714f
C2153 VDD.n1962 GND 0.004714f
C2154 VDD.n1963 GND 0.004714f
C2155 VDD.n1964 GND 0.004714f
C2156 VDD.n1965 GND 0.004714f
C2157 VDD.n1966 GND 0.004714f
C2158 VDD.n1967 GND 0.004714f
C2159 VDD.n1968 GND 0.004714f
C2160 VDD.n1969 GND 0.004714f
C2161 VDD.n1970 GND 0.004714f
C2162 VDD.n1971 GND 0.004714f
C2163 VDD.n1972 GND 0.004714f
C2164 VDD.n1973 GND 0.004714f
C2165 VDD.n1974 GND 0.004714f
C2166 VDD.n1975 GND 0.004714f
C2167 VDD.n1976 GND 0.004714f
C2168 VDD.n1977 GND 0.004714f
C2169 VDD.n1978 GND 0.004714f
C2170 VDD.n1979 GND 0.004714f
C2171 VDD.n1980 GND 0.004714f
C2172 VDD.n1981 GND 0.004714f
C2173 VDD.n1982 GND 0.004714f
C2174 VDD.n1983 GND 0.004714f
C2175 VDD.n1984 GND 0.004714f
C2176 VDD.n1985 GND 0.004714f
C2177 VDD.n1986 GND 0.004714f
C2178 VDD.n1987 GND 0.004714f
C2179 VDD.n1988 GND 0.004714f
C2180 VDD.n1989 GND 0.004714f
C2181 VDD.n1990 GND 0.004714f
C2182 VDD.n1991 GND 0.004714f
C2183 VDD.n1992 GND 0.004714f
C2184 VDD.n1993 GND 0.004714f
C2185 VDD.n1994 GND 0.004714f
C2186 VDD.n1995 GND 0.004714f
C2187 VDD.n1996 GND 0.004714f
C2188 VDD.n1997 GND 0.004714f
C2189 VDD.n1998 GND 0.004714f
C2190 VDD.n1999 GND 0.004714f
C2191 VDD.n2000 GND 0.004714f
C2192 VDD.n2001 GND 0.004714f
C2193 VDD.n2002 GND 0.004714f
C2194 VDD.n2003 GND 0.004714f
C2195 VDD.n2004 GND 0.004714f
C2196 VDD.n2005 GND 0.004714f
C2197 VDD.n2006 GND 0.004714f
C2198 VDD.n2007 GND 0.004714f
C2199 VDD.n2008 GND 0.004714f
C2200 VDD.n2009 GND 0.004714f
C2201 VDD.n2010 GND 0.004714f
C2202 VDD.n2011 GND 0.004714f
C2203 VDD.n2012 GND 0.004714f
C2204 VDD.n2013 GND 0.004714f
C2205 VDD.n2014 GND 0.004714f
C2206 VDD.n2015 GND 0.004714f
C2207 VDD.n2016 GND 0.004714f
C2208 VDD.n2017 GND 0.004714f
C2209 VDD.n2018 GND 0.004714f
C2210 VDD.n2019 GND 0.004714f
C2211 VDD.n2020 GND 0.004714f
C2212 VDD.n2021 GND 0.004714f
C2213 VDD.n2022 GND 0.004714f
C2214 VDD.n2023 GND 0.004714f
C2215 VDD.n2024 GND 0.004714f
C2216 VDD.n2025 GND 0.004714f
C2217 VDD.n2026 GND 0.004714f
C2218 VDD.n2027 GND 0.004714f
C2219 VDD.n2028 GND 0.004714f
C2220 VDD.n2029 GND 0.004714f
C2221 VDD.n2030 GND 0.004714f
C2222 VDD.n2031 GND 0.004714f
C2223 VDD.n2032 GND 0.004714f
C2224 VDD.n2033 GND 0.004714f
C2225 VDD.n2034 GND 0.004714f
C2226 VDD.n2035 GND 0.004714f
C2227 VDD.n2036 GND 0.004714f
C2228 VDD.n2037 GND 0.004714f
C2229 VDD.n2038 GND 0.004714f
C2230 VDD.n2039 GND 0.004714f
C2231 VDD.n2040 GND 0.004714f
C2232 VDD.n2041 GND 0.004714f
C2233 VDD.n2042 GND 0.004714f
C2234 VDD.n2043 GND 0.004714f
C2235 VDD.n2044 GND 0.004714f
C2236 VDD.n2045 GND 0.004714f
C2237 VDD.n2046 GND 0.004714f
C2238 VDD.n2047 GND 0.011836f
C2239 VDD.n2048 GND 0.011836f
C2240 VDD.n2049 GND 0.012357f
C2241 VDD.n2050 GND 0.004714f
C2242 VDD.n2052 GND 0.004714f
C2243 VDD.n2053 GND 0.004714f
C2244 VDD.n2054 GND 0.004714f
C2245 VDD.n2055 GND 0.004714f
C2246 VDD.n2056 GND 0.003882f
C2247 VDD.n2057 GND 0.012357f
C2248 VDD.t55 GND 0.03345f
C2249 VDD.t56 GND 0.055799f
C2250 VDD.t53 GND 0.595646f
C2251 VDD.n2058 GND 0.093248f
C2252 VDD.n2059 GND 0.071157f
C2253 VDD.n2060 GND 0.006737f
C2254 VDD.n2061 GND 0.004714f
C2255 VDD.n2062 GND 0.004714f
C2256 VDD.n2063 GND 0.004714f
C2257 VDD.n2064 GND 0.004714f
C2258 VDD.n2065 GND 0.004714f
C2259 VDD.n2066 GND 0.004714f
C2260 VDD.n2067 GND 0.004714f
C2261 VDD.n2068 GND 0.004714f
C2262 VDD.n2069 GND 0.004714f
C2263 VDD.n2070 GND 0.004714f
C2264 VDD.n2071 GND 0.004714f
C2265 VDD.n2072 GND 0.004714f
C2266 VDD.n2073 GND 0.004714f
C2267 VDD.n2074 GND 0.004714f
C2268 VDD.n2075 GND 0.004714f
C2269 VDD.n2076 GND 0.004714f
C2270 VDD.n2077 GND 0.004714f
C2271 VDD.n2078 GND 0.004714f
C2272 VDD.n2079 GND 0.004714f
C2273 VDD.n2080 GND 0.004714f
C2274 VDD.n2081 GND 0.004714f
C2275 VDD.n2082 GND 0.004714f
C2276 VDD.n2083 GND 0.004714f
C2277 VDD.n2084 GND 0.004714f
C2278 VDD.n2085 GND 0.004714f
C2279 VDD.n2086 GND 0.004714f
C2280 VDD.n2087 GND 0.004714f
C2281 VDD.n2088 GND 0.004714f
C2282 VDD.n2089 GND 0.004714f
C2283 VDD.n2090 GND 0.004714f
C2284 VDD.n2091 GND 0.004714f
C2285 VDD.n2092 GND 0.004714f
C2286 VDD.n2093 GND 0.004714f
C2287 VDD.n2094 GND 0.004714f
C2288 VDD.n2095 GND 0.004714f
C2289 VDD.n2096 GND 0.004714f
C2290 VDD.n2097 GND 0.004714f
C2291 VDD.n2098 GND 0.004714f
C2292 VDD.n2099 GND 0.004714f
C2293 VDD.n2100 GND 0.004714f
C2294 VDD.n2101 GND 0.004714f
C2295 VDD.n2102 GND 0.004714f
C2296 VDD.n2103 GND 0.004714f
C2297 VDD.n2104 GND 0.004714f
C2298 VDD.n2105 GND 0.004714f
C2299 VDD.n2106 GND 0.004714f
C2300 VDD.n2107 GND 0.004714f
C2301 VDD.n2108 GND 0.004714f
C2302 VDD.n2109 GND 0.004714f
C2303 VDD.n2110 GND 0.004714f
C2304 VDD.n2111 GND 0.004714f
C2305 VDD.n2112 GND 0.004714f
C2306 VDD.n2113 GND 0.004714f
C2307 VDD.n2114 GND 0.004714f
C2308 VDD.n2115 GND 0.004714f
C2309 VDD.n2116 GND 0.004714f
C2310 VDD.n2117 GND 0.004714f
C2311 VDD.n2118 GND 0.004714f
C2312 VDD.n2119 GND 0.004714f
C2313 VDD.n2120 GND 0.004714f
C2314 VDD.n2121 GND 0.004714f
C2315 VDD.n2122 GND 0.004714f
C2316 VDD.n2123 GND 0.004714f
C2317 VDD.n2124 GND 0.004714f
C2318 VDD.n2125 GND 0.004714f
C2319 VDD.n2126 GND 0.004714f
C2320 VDD.n2127 GND 0.004714f
C2321 VDD.n2128 GND 0.004714f
C2322 VDD.n2129 GND 0.004714f
C2323 VDD.n2130 GND 0.004714f
C2324 VDD.n2131 GND 0.004714f
C2325 VDD.n2132 GND 0.004714f
C2326 VDD.n2133 GND 0.004714f
C2327 VDD.n2134 GND 0.004714f
C2328 VDD.n2135 GND 0.004714f
C2329 VDD.n2136 GND 0.004714f
C2330 VDD.n2137 GND 0.004714f
C2331 VDD.n2138 GND 0.004714f
C2332 VDD.n2139 GND 0.004714f
C2333 VDD.n2140 GND 0.004714f
C2334 VDD.n2141 GND 0.004714f
C2335 VDD.n2142 GND 0.004714f
C2336 VDD.n2143 GND 0.004714f
C2337 VDD.n2144 GND 0.004714f
C2338 VDD.n2145 GND 0.004714f
C2339 VDD.n2146 GND 0.004714f
C2340 VDD.n2147 GND 0.004714f
C2341 VDD.n2148 GND 0.004714f
C2342 VDD.n2149 GND 0.004714f
C2343 VDD.n2150 GND 0.004714f
C2344 VDD.n2151 GND 0.004714f
C2345 VDD.n2152 GND 0.004714f
C2346 VDD.n2153 GND 0.004714f
C2347 VDD.n2154 GND 0.004714f
C2348 VDD.n2155 GND 0.004714f
C2349 VDD.n2156 GND 0.004714f
C2350 VDD.n2157 GND 0.004714f
C2351 VDD.n2158 GND 0.004714f
C2352 VDD.n2159 GND 0.004714f
C2353 VDD.n2160 GND 0.004714f
C2354 VDD.n2161 GND 0.004714f
C2355 VDD.n2162 GND 0.004714f
C2356 VDD.n2163 GND 0.004714f
C2357 VDD.n2164 GND 0.004714f
C2358 VDD.n2165 GND 0.004714f
C2359 VDD.n2166 GND 0.004714f
C2360 VDD.n2167 GND 0.011836f
C2361 VDD.n2168 GND 0.012357f
C2362 VDD.n2169 GND 0.003189f
C2363 VDD.n2170 GND 0.004714f
C2364 VDD.n2172 GND 0.004714f
C2365 VDD.n2174 GND 0.004714f
C2366 VDD.n2175 GND 0.004714f
C2367 VDD.n2176 GND 0.004714f
C2368 VDD.n2177 GND 0.004714f
C2369 VDD.n2178 GND 0.004714f
C2370 VDD.n2180 GND 0.004714f
C2371 VDD.n2182 GND 0.004714f
C2372 VDD.n2183 GND 0.004714f
C2373 VDD.n2184 GND 0.004714f
C2374 VDD.n2185 GND 0.004714f
C2375 VDD.n2186 GND 0.004714f
C2376 VDD.n2188 GND 0.004714f
C2377 VDD.n2189 GND 0.004714f
C2378 VDD.n2190 GND 0.004714f
C2379 VDD.n2191 GND 0.004714f
C2380 VDD.n2192 GND 0.004714f
C2381 VDD.n2193 GND 0.004714f
C2382 VDD.n2195 GND 0.004714f
C2383 VDD.n2196 GND 0.004714f
C2384 VDD.n2197 GND 0.012357f
C2385 VDD.n2198 GND 0.011836f
C2386 VDD.n2199 GND 0.011836f
C2387 VDD.n2200 GND 0.391281f
C2388 VDD.n2201 GND 0.011836f
C2389 VDD.n2202 GND 0.011836f
C2390 VDD.n2203 GND 0.004714f
C2391 VDD.n2204 GND 0.004714f
C2392 VDD.n2205 GND 0.004714f
C2393 VDD.n2206 GND 0.253401f
C2394 VDD.n2207 GND 0.004714f
C2395 VDD.n2208 GND 0.004714f
C2396 VDD.n2209 GND 0.004714f
C2397 VDD.n2210 GND 0.004714f
C2398 VDD.n2211 GND 0.004714f
C2399 VDD.n2212 GND 0.253401f
C2400 VDD.n2213 GND 0.004714f
C2401 VDD.n2214 GND 0.004714f
C2402 VDD.n2215 GND 0.004714f
C2403 VDD.n2216 GND 0.004714f
C2404 VDD.n2217 GND 0.004714f
C2405 VDD.n2218 GND 0.253401f
C2406 VDD.n2219 GND 0.004714f
C2407 VDD.n2220 GND 0.004714f
C2408 VDD.n2221 GND 0.004714f
C2409 VDD.n2222 GND 0.004714f
C2410 VDD.n2223 GND 0.004714f
C2411 VDD.n2224 GND 0.253401f
C2412 VDD.n2225 GND 0.004714f
C2413 VDD.n2226 GND 0.004714f
C2414 VDD.n2227 GND 0.004714f
C2415 VDD.n2228 GND 0.004714f
C2416 VDD.n2229 GND 0.004714f
C2417 VDD.n2230 GND 0.128564f
C2418 VDD.n2231 GND 0.004714f
C2419 VDD.n2232 GND 0.004714f
C2420 VDD.n2233 GND 0.004714f
C2421 VDD.n2234 GND 0.004714f
C2422 VDD.n2235 GND 0.004714f
C2423 VDD.n2236 GND 0.253401f
C2424 VDD.n2237 GND 0.004714f
C2425 VDD.n2238 GND 0.004714f
C2426 VDD.n2239 GND 0.004714f
C2427 VDD.n2240 GND 0.004714f
C2428 VDD.n2241 GND 0.004714f
C2429 VDD.n2242 GND 0.253401f
C2430 VDD.n2243 GND 0.004714f
C2431 VDD.n2244 GND 0.004714f
C2432 VDD.n2245 GND 0.004714f
C2433 VDD.n2246 GND 0.004714f
C2434 VDD.n2247 GND 0.004714f
C2435 VDD.n2248 GND 0.253401f
C2436 VDD.n2249 GND 0.004714f
C2437 VDD.n2250 GND 0.004714f
C2438 VDD.n2251 GND 0.004714f
C2439 VDD.n2252 GND 0.004714f
C2440 VDD.n2253 GND 0.004714f
C2441 VDD.n2254 GND 0.253401f
C2442 VDD.n2255 GND 0.004714f
C2443 VDD.n2256 GND 0.004714f
C2444 VDD.n2257 GND 0.004714f
C2445 VDD.n2258 GND 0.004714f
C2446 VDD.n2259 GND 0.004714f
C2447 VDD.n2260 GND 0.253401f
C2448 VDD.n2261 GND 0.004714f
C2449 VDD.n2262 GND 0.004714f
C2450 VDD.n2263 GND 0.004714f
C2451 VDD.n2264 GND 0.004714f
C2452 VDD.n2265 GND 0.004714f
C2453 VDD.n2266 GND 0.253401f
C2454 VDD.n2267 GND 0.004714f
C2455 VDD.n2268 GND 0.004714f
C2456 VDD.n2269 GND 0.004714f
C2457 VDD.n2270 GND 0.004714f
C2458 VDD.n2271 GND 0.004714f
C2459 VDD.n2272 GND 0.253401f
C2460 VDD.n2273 GND 0.004714f
C2461 VDD.n2274 GND 0.004714f
C2462 VDD.n2275 GND 0.004714f
C2463 VDD.n2276 GND 0.004714f
C2464 VDD.n2277 GND 0.004714f
C2465 VDD.n2278 GND 0.245948f
C2466 VDD.n2279 GND 0.004714f
C2467 VDD.n2280 GND 0.004714f
C2468 VDD.n2281 GND 0.004714f
C2469 VDD.n2282 GND 0.004714f
C2470 VDD.n2283 GND 0.004714f
C2471 VDD.n2284 GND 0.253401f
C2472 VDD.n2285 GND 0.004714f
C2473 VDD.n2286 GND 0.004714f
C2474 VDD.n2287 GND 0.004714f
C2475 VDD.n2288 GND 0.004714f
C2476 VDD.n2289 GND 0.004714f
C2477 VDD.n2290 GND 0.236632f
C2478 VDD.n2291 GND 0.004714f
C2479 VDD.n2292 GND 0.004714f
C2480 VDD.n2293 GND 0.004714f
C2481 VDD.n2294 GND 0.004714f
C2482 VDD.n2295 GND 0.004714f
C2483 VDD.n2296 GND 0.253401f
C2484 VDD.n2297 GND 0.004714f
C2485 VDD.n2298 GND 0.004714f
C2486 VDD.n2299 GND 0.004714f
C2487 VDD.n2300 GND 0.004714f
C2488 VDD.n2301 GND 0.004714f
C2489 VDD.n2302 GND 0.253401f
C2490 VDD.n2303 GND 0.004714f
C2491 VDD.n2304 GND 0.004714f
C2492 VDD.n2305 GND 0.004714f
C2493 VDD.n2306 GND 0.004714f
C2494 VDD.n2307 GND 0.004714f
C2495 VDD.n2308 GND 0.253401f
C2496 VDD.n2309 GND 0.004714f
C2497 VDD.n2310 GND 0.004714f
C2498 VDD.n2311 GND 0.004714f
C2499 VDD.n2312 GND 0.004714f
C2500 VDD.n2313 GND 0.004714f
C2501 VDD.n2314 GND 0.253401f
C2502 VDD.n2315 GND 0.004714f
C2503 VDD.n2316 GND 0.004714f
C2504 VDD.n2317 GND 0.004714f
C2505 VDD.n2318 GND 0.004714f
C2506 VDD.n2319 GND 0.004714f
C2507 VDD.n2320 GND 0.253401f
C2508 VDD.n2321 GND 0.004714f
C2509 VDD.n2322 GND 0.004714f
C2510 VDD.n2323 GND 0.004714f
C2511 VDD.n2324 GND 0.004714f
C2512 VDD.n2325 GND 0.004714f
C2513 VDD.n2326 GND 0.253401f
C2514 VDD.n2327 GND 0.004714f
C2515 VDD.n2328 GND 0.004714f
C2516 VDD.n2329 GND 0.004714f
C2517 VDD.n2330 GND 0.004714f
C2518 VDD.n2331 GND 0.004714f
C2519 VDD.n2332 GND 0.167692f
C2520 VDD.n2333 GND 0.004714f
C2521 VDD.n2334 GND 0.004714f
C2522 VDD.n2335 GND 0.004714f
C2523 VDD.n2336 GND 0.004714f
C2524 VDD.n2337 GND 0.004714f
C2525 VDD.n2338 GND 0.14347f
C2526 VDD.n2339 GND 0.004714f
C2527 VDD.n2340 GND 0.004714f
C2528 VDD.n2341 GND 0.004714f
C2529 VDD.n2342 GND 0.004714f
C2530 VDD.n2343 GND 0.004714f
C2531 VDD.n2344 GND 0.253401f
C2532 VDD.n2345 GND 0.004714f
C2533 VDD.n2346 GND 0.004714f
C2534 VDD.n2347 GND 0.004714f
C2535 VDD.n2348 GND 0.004714f
C2536 VDD.n2349 GND 0.004714f
C2537 VDD.n2350 GND 0.253401f
C2538 VDD.n2351 GND 0.004714f
C2539 VDD.n2352 GND 0.004714f
C2540 VDD.n2353 GND 0.004714f
C2541 VDD.n2354 GND 0.004714f
C2542 VDD.n2355 GND 0.004714f
C2543 VDD.n2356 GND 0.253401f
C2544 VDD.n2357 GND 0.004714f
C2545 VDD.n2358 GND 0.004714f
C2546 VDD.n2359 GND 0.004714f
C2547 VDD.n2360 GND 0.004714f
C2548 VDD.n2361 GND 0.004714f
C2549 VDD.n2362 GND 0.253401f
C2550 VDD.n2363 GND 0.004714f
C2551 VDD.n2364 GND 0.004714f
C2552 VDD.n2365 GND 0.004714f
C2553 VDD.n2366 GND 0.004714f
C2554 VDD.n2367 GND 0.004714f
C2555 VDD.n2368 GND 0.253401f
C2556 VDD.n2369 GND 0.004714f
C2557 VDD.n2370 GND 0.004714f
C2558 VDD.n2371 GND 0.004714f
C2559 VDD.n2372 GND 0.004714f
C2560 VDD.n2373 GND 0.004714f
C2561 VDD.n2374 GND 0.253401f
C2562 VDD.n2375 GND 0.004714f
C2563 VDD.n2376 GND 0.004714f
C2564 VDD.n2377 GND 0.004714f
C2565 VDD.n2378 GND 0.004714f
C2566 VDD.n2379 GND 0.004714f
C2567 VDD.n2380 GND 0.178871f
C2568 VDD.n2381 GND 0.004714f
C2569 VDD.n2382 GND 0.004714f
C2570 VDD.n2383 GND 0.004714f
C2571 VDD.n2384 GND 0.004714f
C2572 VDD.n2385 GND 0.004714f
C2573 VDD.n2386 GND 0.253401f
C2574 VDD.n2387 GND 0.004714f
C2575 VDD.n2388 GND 0.004714f
C2576 VDD.n2389 GND 0.004714f
C2577 VDD.n2390 GND 0.004714f
C2578 VDD.n2391 GND 0.004714f
C2579 VDD.n2392 GND 0.253401f
C2580 VDD.n2393 GND 0.004714f
C2581 VDD.n2394 GND 0.004714f
C2582 VDD.n2395 GND 0.004714f
C2583 VDD.n2396 GND 0.004714f
C2584 VDD.n2397 GND 0.004714f
C2585 VDD.n2398 GND 0.150923f
C2586 VDD.n2399 GND 0.004714f
C2587 VDD.n2400 GND 0.004714f
C2588 VDD.n2401 GND 0.004714f
C2589 VDD.n2402 GND 0.004714f
C2590 VDD.n2403 GND 0.004714f
C2591 VDD.n2404 GND 0.253401f
C2592 VDD.n2405 GND 0.004714f
C2593 VDD.n2406 GND 0.004714f
C2594 VDD.n2407 GND 0.004714f
C2595 VDD.n2408 GND 0.012357f
C2596 VDD.n2409 GND 0.004714f
C2597 VDD.n2410 GND 0.004714f
C2598 VDD.n2413 GND 0.004714f
C2599 VDD.n2414 GND 0.004714f
C2600 VDD.n2415 GND 0.004714f
C2601 VDD.n2416 GND 0.004714f
C2602 VDD.n2418 GND 0.004714f
C2603 VDD.n2419 GND 0.004714f
C2604 VDD.n2420 GND 0.004714f
C2605 VDD.n2421 GND 0.004714f
C2606 VDD.n2422 GND 0.004714f
C2607 VDD.n2423 GND 0.004714f
C2608 VDD.n2425 GND 0.012357f
C2609 VDD.n2426 GND 0.011836f
C2610 VDD.n2427 GND 0.011836f
C2611 VDD.n2428 GND 0.004714f
C2612 VDD.n2429 GND 0.004714f
C2613 VDD.n2430 GND 0.004714f
C2614 VDD.n2431 GND 0.004714f
C2615 VDD.n2432 GND 0.004714f
C2616 VDD.n2433 GND 0.004714f
C2617 VDD.n2434 GND 0.004714f
C2618 VDD.n2435 GND 0.253401f
C2619 VDD.n2436 GND 0.004714f
C2620 VDD.n2437 GND 0.004714f
C2621 VDD.n2438 GND 0.004714f
C2622 VDD.n2439 GND 0.004714f
C2623 VDD.n2440 GND 0.004714f
C2624 VDD.n2441 GND 0.253401f
C2625 VDD.n2442 GND 0.004714f
C2626 VDD.n2443 GND 0.004714f
C2627 VDD.n2444 GND 0.004714f
C2628 VDD.n2445 GND 0.004714f
C2629 VDD.n2446 GND 0.012322f
C2630 VDD.n2448 GND 0.011836f
C2631 VDD.n2449 GND 0.012357f
C2632 VDD.n2450 GND 0.011872f
C2633 VDD.n2451 GND 0.003189f
C2634 VDD.n2452 GND 0.006737f
C2635 VDD.n2453 GND 0.003882f
C2636 VDD.n2454 GND 0.004714f
C2637 VDD.n2456 GND 0.004714f
C2638 VDD.n2457 GND 0.004714f
C2639 VDD.n2458 GND 0.004714f
C2640 VDD.n2459 GND 0.004714f
C2641 VDD.n2460 GND 0.004714f
C2642 VDD.n2461 GND 0.004714f
C2643 VDD.n2463 GND 0.004714f
C2644 VDD.n2464 GND 0.003535f
C2645 VDD.n2465 GND 0.004714f
C2646 VDD.n2467 GND 0.004714f
C2647 VDD.n2468 GND 0.004714f
C2648 VDD.n2469 GND 0.004714f
C2649 VDD.n2470 GND 0.004714f
C2650 VDD.n2471 GND 0.004714f
C2651 VDD.n2472 GND 0.004714f
C2652 VDD.n2474 GND 0.004714f
C2653 VDD.n2475 GND 0.004714f
C2654 VDD.n2477 GND 0.012357f
C2655 VDD.n2478 GND 0.012357f
C2656 VDD.n2479 GND 0.011836f
C2657 VDD.n2480 GND 0.004714f
C2658 VDD.n2481 GND 0.004714f
C2659 VDD.n2482 GND 0.253401f
C2660 VDD.n2483 GND 0.004714f
C2661 VDD.n2484 GND 0.004714f
C2662 VDD.n2485 GND 0.012322f
C2663 VDD.n2486 GND 0.011872f
C2664 VDD.n2487 GND 0.012357f
C2665 VDD.n2489 GND 0.004714f
C2666 VDD.n2490 GND 0.004714f
C2667 VDD.n2491 GND 0.003882f
C2668 VDD.n2492 GND 0.004714f
C2669 VDD.n2493 GND 0.004714f
C2670 VDD.n2494 GND 0.004714f
C2671 VDD.n2496 GND 0.004714f
C2672 VDD.n2497 GND 0.004714f
C2673 VDD.n2499 GND 0.004714f
C2674 VDD.n2500 GND 0.003535f
C2675 VDD.n2501 GND 0.209537f
C2676 VDD.n2502 GND 2.07275f
C2677 VDD.n2503 GND 0.002539f
C2678 VDD.n2504 GND 0.00201f
C2679 VDD.n2505 GND 0.003466f
C2680 VDD.n2506 GND 0.003041f
C2681 VDD.n2507 GND 0.00558f
C2682 VDD.n2508 GND 0.006932f
C2683 VDD.n2510 GND 0.006932f
C2684 VDD.n2512 GND 0.006932f
C2685 VDD.n2513 GND 0.00558f
C2686 VDD.n2514 GND 0.00558f
C2687 VDD.n2515 GND 0.00558f
C2688 VDD.n2516 GND 0.006932f
C2689 VDD.n2518 GND 0.006932f
C2690 VDD.n2520 GND 0.006932f
C2691 VDD.n2521 GND 0.005496f
C2692 VDD.n2522 GND 0.011382f
C2693 VDD.n2523 GND 0.003822f
C2694 VDD.n2524 GND 0.006932f
C2695 VDD.n2526 GND 0.006932f
C2696 VDD.n2528 GND 0.006932f
C2697 VDD.n2529 GND 0.00558f
C2698 VDD.n2530 GND 0.00558f
C2699 VDD.n2531 GND 0.00558f
C2700 VDD.n2532 GND 0.006932f
C2701 VDD.n2534 GND 0.006932f
C2702 VDD.n2536 GND 0.006932f
C2703 VDD.n2537 GND 0.00558f
C2704 VDD.n2538 GND 0.004715f
C2705 VDD.n2539 GND 0.011382f
C2706 VDD.n2540 GND 0.006932f
C2707 VDD.n2542 GND 0.006932f
C2708 VDD.n2543 GND 0.006932f
C2709 VDD.n2544 GND 0.00558f
C2710 VDD.n2545 GND 0.00558f
C2711 VDD.n2546 GND 0.006932f
C2712 VDD.n2547 GND 0.006932f
C2713 VDD.n2549 GND 0.006932f
C2714 VDD.n2550 GND 0.00558f
C2715 VDD.n2551 GND 0.004631f
C2716 VDD.n2552 GND 0.00201f
C2717 VDD.n2553 GND 2.06314f
C2718 VDD.n2554 GND 0.030878f
C2719 VDD.n2555 GND 0.011479f
C2720 VDD.n2556 GND 0.004631f
C2721 VDD.n2557 GND 0.016004f
C2722 VDD.n2558 GND 0.495623f
C2723 VDD.n2559 GND 0.016004f
C2724 VDD.n2560 GND 0.004631f
C2725 VDD.n2561 GND 0.007799f
C2726 VDD.n2562 GND 0.006932f
C2727 VDD.n2563 GND 0.006932f
C2728 VDD.n2564 GND 0.00558f
C2729 VDD.n2565 GND 0.006932f
C2730 VDD.n2566 GND 0.283213f
C2731 VDD.n2567 GND 0.372649f
C2732 VDD.n2568 GND 0.006932f
C2733 VDD.n2569 GND 0.00558f
C2734 VDD.n2570 GND 0.006932f
C2735 VDD.n2571 GND 0.006932f
C2736 VDD.n2572 GND 0.006932f
C2737 VDD.n2573 GND 0.00558f
C2738 VDD.n2574 GND 0.006932f
C2739 VDD.n2575 GND 0.27576f
C2740 VDD.n2576 GND 0.006932f
C2741 VDD.n2577 GND 0.00558f
C2742 VDD.n2578 GND 0.006932f
C2743 VDD.n2579 GND 0.006932f
C2744 VDD.n2580 GND 0.006932f
C2745 VDD.n2581 GND 0.00558f
C2746 VDD.n2582 GND 0.006932f
C2747 VDD.n2583 GND 0.372649f
C2748 VDD.n2584 GND 0.006932f
C2749 VDD.n2585 GND 0.00558f
C2750 VDD.n2586 GND 0.006932f
C2751 VDD.n2587 GND 0.006932f
C2752 VDD.n2588 GND 0.006932f
C2753 VDD.n2589 GND 0.00558f
C2754 VDD.n2590 GND 0.006932f
C2755 VDD.n2591 GND 0.372649f
C2756 VDD.n2592 GND 0.006932f
C2757 VDD.n2593 GND 0.00558f
C2758 VDD.n2594 GND 0.006932f
C2759 VDD.n2595 GND 0.006932f
C2760 VDD.n2596 GND 0.006932f
C2761 VDD.n2597 GND 0.00558f
C2762 VDD.n2598 GND 0.006932f
C2763 VDD.n2599 GND 0.372649f
C2764 VDD.n2600 GND 0.006932f
C2765 VDD.n2601 GND 0.00558f
C2766 VDD.n2602 GND 0.006932f
C2767 VDD.n2603 GND 0.006932f
C2768 VDD.n2604 GND 0.006932f
C2769 VDD.n2605 GND 0.00558f
C2770 VDD.n2606 GND 0.006932f
C2771 VDD.n2607 GND 0.227316f
C2772 VDD.n2608 GND 0.006932f
C2773 VDD.n2609 GND 0.00558f
C2774 VDD.n2610 GND 0.006932f
C2775 VDD.n2611 GND 0.006932f
C2776 VDD.n2612 GND 0.006932f
C2777 VDD.n2613 GND 0.00558f
C2778 VDD.n2614 GND 0.006932f
C2779 VDD.n2615 GND 0.372649f
C2780 VDD.n2616 GND 0.006932f
C2781 VDD.n2617 GND 0.00558f
C2782 VDD.n2618 GND 0.006932f
C2783 VDD.n2619 GND 0.006932f
C2784 VDD.n2620 GND 0.006932f
C2785 VDD.n2621 GND 0.00558f
C2786 VDD.n2622 GND 0.006932f
C2787 VDD.n2623 GND 0.372649f
C2788 VDD.n2624 GND 0.006932f
C2789 VDD.n2625 GND 0.00558f
C2790 VDD.n2626 GND 0.006932f
C2791 VDD.n2627 GND 0.006932f
C2792 VDD.n2628 GND 0.006932f
C2793 VDD.n2629 GND 0.00558f
C2794 VDD.n2630 GND 0.006932f
C2795 VDD.t122 GND 0.186324f
C2796 VDD.n2631 GND 0.324204f
C2797 VDD.n2632 GND 0.006932f
C2798 VDD.n2633 GND 0.00558f
C2799 VDD.n2634 GND 0.006932f
C2800 VDD.n2635 GND 0.006932f
C2801 VDD.n2636 GND 0.006932f
C2802 VDD.n2637 GND 0.00558f
C2803 VDD.n2638 GND 0.006932f
C2804 VDD.n2639 GND 0.372649f
C2805 VDD.n2640 GND 0.006932f
C2806 VDD.n2641 GND 0.00558f
C2807 VDD.n2642 GND 0.006932f
C2808 VDD.n2643 GND 0.006932f
C2809 VDD.n2644 GND 0.006932f
C2810 VDD.n2645 GND 0.00558f
C2811 VDD.n2646 GND 0.00558f
C2812 VDD.n2647 GND 0.00558f
C2813 VDD.n2648 GND 0.006932f
C2814 VDD.n2649 GND 0.006932f
C2815 VDD.n2650 GND 0.006932f
C2816 VDD.n2651 GND 0.00558f
C2817 VDD.n2652 GND 0.00558f
C2818 VDD.n2653 GND 0.00558f
C2819 VDD.n2654 GND 0.006932f
C2820 VDD.n2655 GND 0.006932f
C2821 VDD.n2656 GND 0.006932f
C2822 VDD.n2657 GND 0.00558f
C2823 VDD.n2658 GND 0.00558f
C2824 VDD.n2659 GND 0.00558f
C2825 VDD.n2660 GND 0.006932f
C2826 VDD.n2661 GND 0.006932f
C2827 VDD.n2662 GND 0.006932f
C2828 VDD.n2663 GND 0.00558f
C2829 VDD.n2664 GND 0.00558f
C2830 VDD.n2665 GND 0.00558f
C2831 VDD.n2666 GND 0.006932f
C2832 VDD.n2667 GND 0.006932f
C2833 VDD.n2668 GND 0.006932f
C2834 VDD.n2669 GND 0.00558f
C2835 VDD.n2670 GND 0.00558f
C2836 VDD.n2671 GND 0.00558f
C2837 VDD.n2672 GND 0.006932f
C2838 VDD.n2673 GND 0.006932f
C2839 VDD.n2674 GND 0.006932f
C2840 VDD.n2675 GND 0.00558f
C2841 VDD.n2676 GND 0.00558f
C2842 VDD.n2677 GND 0.004631f
C2843 VDD.n2678 GND 0.016004f
C2844 VDD.n2679 GND 0.016092f
C2845 VDD.n2680 GND 0.002539f
C2846 VDD.n2681 GND 0.016092f
C2847 VDD.n2683 GND 0.006932f
C2848 VDD.n2684 GND 0.006932f
C2849 VDD.n2685 GND 0.00558f
C2850 VDD.n2686 GND 0.00558f
C2851 VDD.n2687 GND 0.00558f
C2852 VDD.n2688 GND 0.006932f
C2853 VDD.n2690 GND 0.006932f
C2854 VDD.n2691 GND 0.006932f
C2855 VDD.n2693 GND 0.006932f
C2856 VDD.n2694 GND 0.00558f
C2857 VDD.n2695 GND 0.006932f
C2858 VDD.n2696 GND 0.006932f
C2859 VDD.n2697 GND 0.006932f
C2860 VDD.n2698 GND 0.011382f
C2861 VDD.n2699 GND 0.003822f
C2862 VDD.n2700 GND 0.006932f
C2863 VDD.n2702 GND 0.006932f
C2864 VDD.n2703 GND 0.006932f
C2865 VDD.n2704 GND 0.00558f
C2866 VDD.n2705 GND 0.00558f
C2867 VDD.n2706 GND 0.00558f
C2868 VDD.n2707 GND 0.006932f
C2869 VDD.n2709 GND 0.006932f
C2870 VDD.n2710 GND 0.006932f
C2871 VDD.n2711 GND 0.00558f
C2872 VDD.n2712 GND 0.006932f
C2873 VDD.n2713 GND 0.006932f
C2874 VDD.n2714 GND 0.006932f
C2875 VDD.n2715 GND 0.011382f
C2876 VDD.n2716 GND 0.004603f
C2877 VDD.n2717 GND 0.00558f
C2878 VDD.n2718 GND 0.006932f
C2879 VDD.n2720 GND 0.006932f
C2880 VDD.n2721 GND 0.006932f
C2881 VDD.n2722 GND 0.00558f
C2882 VDD.n2723 GND 0.00558f
C2883 VDD.n2724 GND 0.004631f
C2884 VDD.n2725 GND 0.016092f
C2885 VDD.n2726 GND 0.016004f
C2886 VDD.n2727 GND 0.004631f
C2887 VDD.n2728 GND 0.016004f
C2888 VDD.n2729 GND 0.495623f
C2889 VDD.n2730 GND 0.372649f
C2890 VDD.n2731 GND 0.372649f
C2891 VDD.n2732 GND 0.006932f
C2892 VDD.n2733 GND 0.00558f
C2893 VDD.n2734 GND 0.00558f
C2894 VDD.n2735 GND 0.00558f
C2895 VDD.n2736 GND 0.006932f
C2896 VDD.n2737 GND 0.27576f
C2897 VDD.n2738 GND 0.372649f
C2898 VDD.n2739 GND 0.372649f
C2899 VDD.n2740 GND 0.006932f
C2900 VDD.n2741 GND 0.00558f
C2901 VDD.n2742 GND 0.00558f
C2902 VDD.n2743 GND 0.00558f
C2903 VDD.n2744 GND 0.006932f
C2904 VDD.n2745 GND 0.372649f
C2905 VDD.n2746 GND 0.372649f
C2906 VDD.n2747 GND 0.372649f
C2907 VDD.n2748 GND 0.006932f
C2908 VDD.n2749 GND 0.00558f
C2909 VDD.n2750 GND 0.00558f
C2910 VDD.n2751 GND 0.00558f
C2911 VDD.n2752 GND 0.006932f
C2912 VDD.n2753 GND 0.227316f
C2913 VDD.t110 GND 0.186324f
C2914 VDD.n2754 GND 0.331657f
C2915 VDD.n2755 GND 0.372649f
C2916 VDD.n2756 GND 0.006932f
C2917 VDD.n2757 GND 0.00558f
C2918 VDD.n2758 GND 0.00558f
C2919 VDD.n2759 GND 0.00558f
C2920 VDD.n2760 GND 0.006932f
C2921 VDD.n2761 GND 0.372649f
C2922 VDD.n2762 GND 0.372649f
C2923 VDD.n2763 GND 0.324204f
C2924 VDD.n2764 GND 0.006932f
C2925 VDD.n2765 GND 0.00558f
C2926 VDD.n2766 GND 0.00558f
C2927 VDD.n2767 GND 0.00558f
C2928 VDD.n2768 GND 0.006932f
C2929 VDD.n2769 GND 0.372649f
C2930 VDD.n2770 GND 0.372649f
C2931 VDD.n2771 GND 0.372649f
C2932 VDD.n2772 GND 0.006932f
C2933 VDD.n2773 GND 0.00558f
C2934 VDD.n2774 GND 0.397993f
C2935 VDD.n2775 GND 2.78768f
C2936 a_n16148_7944.n0 GND 27.9869f
C2937 a_n16148_7944.n1 GND 1.0753f
C2938 a_n16148_7944.n2 GND 0.332362f
C2939 a_n16148_7944.n3 GND 1.04582f
C2940 a_n16148_7944.n4 GND 0.332362f
C2941 a_n16148_7944.n5 GND 1.04582f
C2942 a_n16148_7944.n6 GND 0.332362f
C2943 a_n16148_7944.n7 GND 1.0753f
C2944 a_n16148_7944.n8 GND 0.165689f
C2945 a_n16148_7944.n9 GND 1.04582f
C2946 a_n16148_7944.n10 GND 0.165689f
C2947 a_n16148_7944.n11 GND 1.04582f
C2948 a_n16148_7944.n12 GND 0.165689f
C2949 a_n16148_7944.n13 GND 2.54525f
C2950 a_n16148_7944.n14 GND 2.82768f
C2951 a_n16148_7944.n15 GND 0.165689f
C2952 a_n16148_7944.n16 GND 0.165689f
C2953 a_n16148_7944.n17 GND 0.165689f
C2954 a_n16148_7944.n18 GND 0.332366f
C2955 a_n16148_7944.n19 GND 0.332366f
C2956 a_n16148_7944.n20 GND 0.332366f
C2957 a_n16148_7944.t3 GND 0.037883f
C2958 a_n16148_7944.t2 GND 0.037883f
C2959 a_n16148_7944.t4 GND 0.037883f
C2960 a_n16148_7944.n21 GND 1.18976f
C2961 a_n16148_7944.t0 GND 0.236474f
C2962 a_n16148_7944.t1 GND 0.455527f
C2963 a_n16148_7944.n22 GND 2.21683f
C2964 a_n16148_7944.t12 GND 0.837024f
C2965 a_n16148_7944.t7 GND 0.529129f
C2966 a_n16148_7944.t20 GND 0.842555f
C2967 a_n16148_7944.n23 GND 0.357638f
C2968 a_n16148_7944.t23 GND 0.529129f
C2969 a_n16148_7944.n24 GND 0.467446f
C2970 a_n16148_7944.n25 GND 0.467636f
C2971 a_n16148_7944.t8 GND 0.837024f
C2972 a_n16148_7944.t29 GND 0.529129f
C2973 a_n16148_7944.t19 GND 0.842555f
C2974 a_n16148_7944.n26 GND 0.357638f
C2975 a_n16148_7944.t21 GND 0.529129f
C2976 a_n16148_7944.n27 GND 0.467446f
C2977 a_n16148_7944.n28 GND 0.467636f
C2978 a_n16148_7944.t14 GND 0.837024f
C2979 a_n16148_7944.t10 GND 0.529129f
C2980 a_n16148_7944.t22 GND 0.842555f
C2981 a_n16148_7944.n29 GND 0.357638f
C2982 a_n16148_7944.t24 GND 0.529129f
C2983 a_n16148_7944.n30 GND 0.467446f
C2984 a_n16148_7944.n31 GND 0.467636f
C2985 a_n16148_7944.t6 GND 0.837027f
C2986 a_n16148_7944.t17 GND 0.529129f
C2987 a_n16148_7944.t26 GND 0.842553f
C2988 a_n16148_7944.n32 GND 0.357638f
C2989 a_n16148_7944.t13 GND 0.529129f
C2990 a_n16148_7944.n33 GND 0.467447f
C2991 a_n16148_7944.n34 GND 0.467636f
C2992 a_n16148_7944.t28 GND 0.837027f
C2993 a_n16148_7944.t15 GND 0.529129f
C2994 a_n16148_7944.t25 GND 0.842553f
C2995 a_n16148_7944.n35 GND 0.357638f
C2996 a_n16148_7944.t11 GND 0.529129f
C2997 a_n16148_7944.n36 GND 0.467447f
C2998 a_n16148_7944.n37 GND 0.467636f
C2999 a_n16148_7944.t9 GND 0.837027f
C3000 a_n16148_7944.t18 GND 0.529129f
C3001 a_n16148_7944.t27 GND 0.842553f
C3002 a_n16148_7944.n38 GND 0.357638f
C3003 a_n16148_7944.t16 GND 0.529129f
C3004 a_n16148_7944.n39 GND 0.467447f
C3005 a_n16148_7944.n40 GND 0.467636f
C3006 a_n16148_7944.n41 GND 9.21097f
C3007 a_n16148_7944.n42 GND 0.973476f
C3008 a_n16148_7944.t5 GND 0.037883f
C3009 a_n4238_7449.n0 GND 7.69508f
C3010 a_n4238_7449.n1 GND 0.010337f
C3011 a_n4238_7449.n2 GND 0.032837f
C3012 a_n4238_7449.n3 GND 0.010337f
C3013 a_n4238_7449.n4 GND 0.032837f
C3014 a_n4238_7449.n5 GND 0.010337f
C3015 a_n4238_7449.n6 GND 0.032837f
C3016 a_n4238_7449.n7 GND 0.010337f
C3017 a_n4238_7449.n8 GND 0.032837f
C3018 a_n4238_7449.n9 GND 0.010337f
C3019 a_n4238_7449.n10 GND 0.032837f
C3020 a_n4238_7449.n11 GND 0.010337f
C3021 a_n4238_7449.n12 GND 0.032837f
C3022 a_n4238_7449.n13 GND 0.010337f
C3023 a_n4238_7449.n14 GND 0.032837f
C3024 a_n4238_7449.n15 GND 0.010337f
C3025 a_n4238_7449.n16 GND 0.032837f
C3026 a_n4238_7449.n17 GND 1.03285f
C3027 a_n4238_7449.n18 GND 0.710651f
C3028 a_n4238_7449.n19 GND 0.243235f
C3029 a_n4238_7449.n20 GND 0.018853f
C3030 a_n4238_7449.n21 GND 0.243235f
C3031 a_n4238_7449.n22 GND 0.018853f
C3032 a_n4238_7449.n23 GND 0.243235f
C3033 a_n4238_7449.n24 GND 0.018853f
C3034 a_n4238_7449.n25 GND 0.243235f
C3035 a_n4238_7449.n26 GND 0.018853f
C3036 a_n4238_7449.n27 GND 0.243235f
C3037 a_n4238_7449.n28 GND 0.018853f
C3038 a_n4238_7449.n29 GND 0.243235f
C3039 a_n4238_7449.n30 GND 0.018853f
C3040 a_n4238_7449.n31 GND 0.243235f
C3041 a_n4238_7449.n32 GND 0.018853f
C3042 a_n4238_7449.n33 GND 0.243235f
C3043 a_n4238_7449.n34 GND 0.018853f
C3044 a_n4238_7449.t12 GND 36.6464f
C3045 a_n4238_7449.n35 GND 0.016233f
C3046 a_n4238_7449.n36 GND 0.022519f
C3047 a_n4238_7449.n37 GND 0.063393f
C3048 a_n4238_7449.n38 GND 0.016233f
C3049 a_n4238_7449.n39 GND 0.022519f
C3050 a_n4238_7449.n40 GND 0.063393f
C3051 a_n4238_7449.n41 GND 0.016233f
C3052 a_n4238_7449.n42 GND 0.022519f
C3053 a_n4238_7449.n43 GND 0.063393f
C3054 a_n4238_7449.n44 GND 0.016233f
C3055 a_n4238_7449.n45 GND 0.022519f
C3056 a_n4238_7449.n46 GND 0.063393f
C3057 a_n4238_7449.n47 GND 0.016233f
C3058 a_n4238_7449.n48 GND 0.022519f
C3059 a_n4238_7449.n49 GND 0.063393f
C3060 a_n4238_7449.n50 GND 0.016233f
C3061 a_n4238_7449.n51 GND 0.022519f
C3062 a_n4238_7449.n52 GND 0.063393f
C3063 a_n4238_7449.n53 GND 0.016233f
C3064 a_n4238_7449.n54 GND 0.022519f
C3065 a_n4238_7449.n55 GND 0.063393f
C3066 a_n4238_7449.n56 GND 0.016233f
C3067 a_n4238_7449.n57 GND 0.022519f
C3068 a_n4238_7449.n58 GND 0.063393f
C3069 a_n4238_7449.t0 GND 0.049811f
C3070 a_n4238_7449.n59 GND 0.056976f
C3071 a_n4238_7449.n60 GND 0.075381f
C3072 a_n4238_7449.t9 GND 0.049811f
C3073 a_n4238_7449.n61 GND 0.056976f
C3074 a_n4238_7449.n62 GND 0.040699f
C3075 a_n4238_7449.n63 GND 2.23514f
C3076 a_n4238_7449.t3 GND 0.049811f
C3077 a_n4238_7449.n64 GND 0.056976f
C3078 a_n4238_7449.n65 GND 0.075381f
C3079 a_n4238_7449.t11 GND 0.045112f
C3080 a_n4238_7449.t6 GND 0.045112f
C3081 a_n4238_7449.n66 GND 0.21438f
C3082 a_n4238_7449.t1 GND 0.049811f
C3083 a_n4238_7449.n67 GND 0.056976f
C3084 a_n4238_7449.n68 GND 0.040699f
C3085 a_n4238_7449.t8 GND 0.049811f
C3086 a_n4238_7449.n69 GND 0.056976f
C3087 a_n4238_7449.n70 GND 0.040699f
C3088 a_n4238_7449.t10 GND 0.045112f
C3089 a_n4238_7449.t7 GND 0.045112f
C3090 a_n4238_7449.n71 GND 0.21438f
C3091 a_n4238_7449.n72 GND 0.773746f
C3092 a_n4238_7449.t5 GND 0.049811f
C3093 a_n4238_7449.n73 GND 0.056976f
C3094 a_n4238_7449.n74 GND 0.040699f
C3095 a_n4238_7449.n75 GND 0.595631f
C3096 a_n4238_7449.t2 GND 0.049811f
C3097 a_n4238_7449.n76 GND 0.056976f
C3098 a_n4238_7449.n77 GND 0.075381f
C3099 a_n4238_7449.t4 GND 0.049811f
C3100 a_n4238_7449.n78 GND 0.056976f
C3101 a_n4238_7449.n79 GND 0.040699f
C3102 a_n4238_7449.n80 GND 1.65809f
C3103 a_n10279_8682.n0 GND 9.19557f
C3104 a_n10279_8682.n1 GND 21.2555f
C3105 a_n10279_8682.n2 GND 1.8253f
C3106 a_n10279_8682.t28 GND 2.52592f
C3107 a_n10279_8682.t23 GND 2.52592f
C3108 a_n10279_8682.n3 GND 0.762833f
C3109 a_n10279_8682.t17 GND 2.51319f
C3110 a_n10279_8682.n4 GND 0.409118f
C3111 a_n10279_8682.n5 GND 2.54647f
C3112 a_n10279_8682.n6 GND 2.38741f
C3113 a_n10279_8682.t14 GND 2.88729f
C3114 a_n10279_8682.t2 GND 2.88729f
C3115 a_n10279_8682.t12 GND 2.91585f
C3116 a_n10279_8682.t29 GND 2.91585f
C3117 a_n10279_8682.t18 GND 2.91585f
C3118 a_n10279_8682.t25 GND 2.91585f
C3119 a_n10279_8682.t4 GND 2.86779f
C3120 a_n10279_8682.t10 GND 2.86779f
C3121 a_n10279_8682.t7 GND 0.179302f
C3122 a_n10279_8682.t9 GND 0.165421f
C3123 a_n10279_8682.n7 GND 2.26879f
C3124 a_n10279_8682.t8 GND 2.86779f
C3125 a_n10279_8682.t6 GND 2.88729f
C3126 a_n10279_8682.t11 GND 2.86779f
C3127 a_n10279_8682.t24 GND 2.88729f
C3128 a_n10279_8682.t22 GND 2.87384f
C3129 a_n10279_8682.t27 GND 2.86544f
C3130 a_n10279_8682.t13 GND 2.91424f
C3131 a_n10279_8682.t19 GND 2.85286f
C3132 a_n10279_8682.t20 GND 2.87384f
C3133 a_n10279_8682.t26 GND 2.86544f
C3134 a_n10279_8682.t21 GND 2.87384f
C3135 a_n10279_8682.t15 GND 2.87158f
C3136 a_n10279_8682.t16 GND 2.53007f
C3137 a_n10279_8682.t0 GND 0.473749f
C3138 a_n10279_8682.t1 GND 0.256705f
C3139 a_n10279_8682.n8 GND 4.04772f
C3140 a_n10279_8682.t5 GND 0.179302f
C3141 a_n10279_8682.n9 GND 2.21155f
C3142 a_n10279_8682.t3 GND 0.165421f
C3143 VOUT.t18 GND 0.012118f
C3144 VOUT.t4 GND 0.012118f
C3145 VOUT.n0 GND 0.058644f
C3146 VOUT.t0 GND 0.012118f
C3147 VOUT.t81 GND 0.012118f
C3148 VOUT.n1 GND 0.05519f
C3149 VOUT.n2 GND 0.469419f
C3150 VOUT.t83 GND 0.012118f
C3151 VOUT.t2 GND 0.012118f
C3152 VOUT.n3 GND 0.058644f
C3153 VOUT.t8 GND 0.012118f
C3154 VOUT.t12 GND 0.012118f
C3155 VOUT.n4 GND 0.05519f
C3156 VOUT.n5 GND 0.453622f
C3157 VOUT.n6 GND 0.174057f
C3158 VOUT.t3 GND 0.012118f
C3159 VOUT.t19 GND 0.012118f
C3160 VOUT.n7 GND 0.058644f
C3161 VOUT.t7 GND 0.012118f
C3162 VOUT.t14 GND 0.012118f
C3163 VOUT.n8 GND 0.05519f
C3164 VOUT.n9 GND 0.453622f
C3165 VOUT.n10 GND 0.282489f
C3166 VOUT.n11 GND 10.3031f
C3167 VOUT.t84 GND 8.75049f
C3168 VOUT.t85 GND 5.76942f
C3169 VOUT.n12 GND 9.327339f
C3170 VOUT.n13 GND 2.27558f
C3171 VOUT.t10 GND 0.012118f
C3172 VOUT.t13 GND 0.012118f
C3173 VOUT.n14 GND 0.058644f
C3174 VOUT.t16 GND 0.012118f
C3175 VOUT.t1 GND 0.012118f
C3176 VOUT.n15 GND 0.05519f
C3177 VOUT.n16 GND 0.469419f
C3178 VOUT.t15 GND 0.012118f
C3179 VOUT.t17 GND 0.012118f
C3180 VOUT.n17 GND 0.058644f
C3181 VOUT.t6 GND 0.012118f
C3182 VOUT.t82 GND 0.012118f
C3183 VOUT.n18 GND 0.05519f
C3184 VOUT.n19 GND 0.453622f
C3185 VOUT.n20 GND 0.174057f
C3186 VOUT.t20 GND 0.012118f
C3187 VOUT.t11 GND 0.012118f
C3188 VOUT.n21 GND 0.058644f
C3189 VOUT.t5 GND 0.012118f
C3190 VOUT.t9 GND 0.012118f
C3191 VOUT.n22 GND 0.05519f
C3192 VOUT.n23 GND 0.453623f
C3193 VOUT.n24 GND 0.282489f
C3194 VOUT.n25 GND 13.4912f
C3195 VOUT.t68 GND 0.022149f
C3196 VOUT.t51 GND 0.022149f
C3197 VOUT.n26 GND 0.177597f
C3198 VOUT.t53 GND 0.022149f
C3199 VOUT.t38 GND 0.022149f
C3200 VOUT.n27 GND 0.172853f
C3201 VOUT.n28 GND 0.31842f
C3202 VOUT.t35 GND 0.022149f
C3203 VOUT.t71 GND 0.022149f
C3204 VOUT.n29 GND 0.172853f
C3205 VOUT.n30 GND 0.220124f
C3206 VOUT.t63 GND 0.022149f
C3207 VOUT.t23 GND 0.022149f
C3208 VOUT.n31 GND 0.177597f
C3209 VOUT.t80 GND 0.022149f
C3210 VOUT.t24 GND 0.022149f
C3211 VOUT.n32 GND 0.172853f
C3212 VOUT.n33 GND 0.31842f
C3213 VOUT.t22 GND 0.022149f
C3214 VOUT.t39 GND 0.022149f
C3215 VOUT.n34 GND 0.172853f
C3216 VOUT.n35 GND 0.195177f
C3217 VOUT.n36 GND 0.209054f
C3218 VOUT.t61 GND 0.022149f
C3219 VOUT.t76 GND 0.022149f
C3220 VOUT.n37 GND 0.177597f
C3221 VOUT.t78 GND 0.022149f
C3222 VOUT.t30 GND 0.022149f
C3223 VOUT.n38 GND 0.172853f
C3224 VOUT.n39 GND 0.31842f
C3225 VOUT.t40 GND 0.022149f
C3226 VOUT.t73 GND 0.022149f
C3227 VOUT.n40 GND 0.172853f
C3228 VOUT.n41 GND 0.195177f
C3229 VOUT.n42 GND 0.145815f
C3230 VOUT.t57 GND 0.022149f
C3231 VOUT.t42 GND 0.022149f
C3232 VOUT.n43 GND 0.177597f
C3233 VOUT.t41 GND 0.022149f
C3234 VOUT.t29 GND 0.022149f
C3235 VOUT.n44 GND 0.172853f
C3236 VOUT.n45 GND 0.31842f
C3237 VOUT.t31 GND 0.022149f
C3238 VOUT.t77 GND 0.022149f
C3239 VOUT.n46 GND 0.172853f
C3240 VOUT.n47 GND 0.195177f
C3241 VOUT.n48 GND 0.145815f
C3242 VOUT.t66 GND 0.022149f
C3243 VOUT.t48 GND 0.022149f
C3244 VOUT.n49 GND 0.177597f
C3245 VOUT.t49 GND 0.022149f
C3246 VOUT.t33 GND 0.022149f
C3247 VOUT.n50 GND 0.172853f
C3248 VOUT.n51 GND 0.31842f
C3249 VOUT.t34 GND 0.022149f
C3250 VOUT.t21 GND 0.022149f
C3251 VOUT.n52 GND 0.172853f
C3252 VOUT.n53 GND 0.195177f
C3253 VOUT.n54 GND 0.263161f
C3254 VOUT.n55 GND 11.6008f
C3255 VOUT.t59 GND 0.022149f
C3256 VOUT.t79 GND 0.022149f
C3257 VOUT.n56 GND 0.177597f
C3258 VOUT.t60 GND 0.022149f
C3259 VOUT.t72 GND 0.022149f
C3260 VOUT.n57 GND 0.172853f
C3261 VOUT.n58 GND 0.31842f
C3262 VOUT.t25 GND 0.022149f
C3263 VOUT.t43 GND 0.022149f
C3264 VOUT.n59 GND 0.172853f
C3265 VOUT.n60 GND 0.220124f
C3266 VOUT.t32 GND 0.022149f
C3267 VOUT.t56 GND 0.022149f
C3268 VOUT.n61 GND 0.177597f
C3269 VOUT.t47 GND 0.022149f
C3270 VOUT.t52 GND 0.022149f
C3271 VOUT.n62 GND 0.172853f
C3272 VOUT.n63 GND 0.31842f
C3273 VOUT.t62 GND 0.022149f
C3274 VOUT.t58 GND 0.022149f
C3275 VOUT.n64 GND 0.172853f
C3276 VOUT.n65 GND 0.195177f
C3277 VOUT.n66 GND 0.209054f
C3278 VOUT.t75 GND 0.022149f
C3279 VOUT.t74 GND 0.022149f
C3280 VOUT.n67 GND 0.177597f
C3281 VOUT.t27 GND 0.022149f
C3282 VOUT.t67 GND 0.022149f
C3283 VOUT.n68 GND 0.172853f
C3284 VOUT.n69 GND 0.31842f
C3285 VOUT.t70 GND 0.022149f
C3286 VOUT.t69 GND 0.022149f
C3287 VOUT.n70 GND 0.172853f
C3288 VOUT.n71 GND 0.195177f
C3289 VOUT.n72 GND 0.145815f
C3290 VOUT.t28 GND 0.022149f
C3291 VOUT.t26 GND 0.022149f
C3292 VOUT.n73 GND 0.177597f
C3293 VOUT.t65 GND 0.022149f
C3294 VOUT.t64 GND 0.022149f
C3295 VOUT.n74 GND 0.172853f
C3296 VOUT.n75 GND 0.31842f
C3297 VOUT.t46 GND 0.022149f
C3298 VOUT.t36 GND 0.022149f
C3299 VOUT.n76 GND 0.172853f
C3300 VOUT.n77 GND 0.195177f
C3301 VOUT.n78 GND 0.145815f
C3302 VOUT.t54 GND 0.022149f
C3303 VOUT.t55 GND 0.022149f
C3304 VOUT.n79 GND 0.177597f
C3305 VOUT.t50 GND 0.022149f
C3306 VOUT.t37 GND 0.022149f
C3307 VOUT.n80 GND 0.172853f
C3308 VOUT.n81 GND 0.31842f
C3309 VOUT.t45 GND 0.022149f
C3310 VOUT.t44 GND 0.022149f
C3311 VOUT.n82 GND 0.172853f
C3312 VOUT.n83 GND 0.195177f
C3313 VOUT.n84 GND 0.263161f
C3314 VOUT.n85 GND 8.76436f
C3315 VOUT.n86 GND 6.11559f
C3316 CS_BIAS.n0 GND 0.010508f
C3317 CS_BIAS.t83 GND 0.172127f
C3318 CS_BIAS.n1 GND 0.007113f
C3319 CS_BIAS.n2 GND 0.007971f
C3320 CS_BIAS.t79 GND 0.172127f
C3321 CS_BIAS.n3 GND 0.015368f
C3322 CS_BIAS.n4 GND 0.007971f
C3323 CS_BIAS.t71 GND 0.172127f
C3324 CS_BIAS.n5 GND 0.070158f
C3325 CS_BIAS.n6 GND 0.007933f
C3326 CS_BIAS.n7 GND 0.015759f
C3327 CS_BIAS.n8 GND 0.010508f
C3328 CS_BIAS.t16 GND 0.172127f
C3329 CS_BIAS.n9 GND 0.007113f
C3330 CS_BIAS.n10 GND 0.007971f
C3331 CS_BIAS.t0 GND 0.172127f
C3332 CS_BIAS.n11 GND 0.015368f
C3333 CS_BIAS.n12 GND 0.007971f
C3334 CS_BIAS.t20 GND 0.172127f
C3335 CS_BIAS.n13 GND 0.070158f
C3336 CS_BIAS.n14 GND 0.007971f
C3337 CS_BIAS.n15 GND 0.015759f
C3338 CS_BIAS.n16 GND 0.007971f
C3339 CS_BIAS.t2 GND 0.172127f
C3340 CS_BIAS.n17 GND 0.006602f
C3341 CS_BIAS.n18 GND 0.06794f
C3342 CS_BIAS.t22 GND 0.172127f
C3343 CS_BIAS.t4 GND 0.222799f
C3344 CS_BIAS.n19 GND 0.087264f
C3345 CS_BIAS.n20 GND 0.091464f
C3346 CS_BIAS.n21 GND 0.012008f
C3347 CS_BIAS.n22 GND 0.015368f
C3348 CS_BIAS.n23 GND 0.007971f
C3349 CS_BIAS.n24 GND 0.007971f
C3350 CS_BIAS.n25 GND 0.007971f
C3351 CS_BIAS.n26 GND 0.015985f
C3352 CS_BIAS.n27 GND 0.010841f
C3353 CS_BIAS.n28 GND 0.070158f
C3354 CS_BIAS.n29 GND 0.011425f
C3355 CS_BIAS.n30 GND 0.007971f
C3356 CS_BIAS.n31 GND 0.007971f
C3357 CS_BIAS.n32 GND 0.007971f
C3358 CS_BIAS.n33 GND 0.006438f
C3359 CS_BIAS.n34 GND 0.015759f
C3360 CS_BIAS.n35 GND 0.011425f
C3361 CS_BIAS.n36 GND 0.007971f
C3362 CS_BIAS.n37 GND 0.007971f
C3363 CS_BIAS.n38 GND 0.010841f
C3364 CS_BIAS.n39 GND 0.015985f
C3365 CS_BIAS.n40 GND 0.006602f
C3366 CS_BIAS.n41 GND 0.007971f
C3367 CS_BIAS.n42 GND 0.007971f
C3368 CS_BIAS.n43 GND 0.007971f
C3369 CS_BIAS.n44 GND 0.012008f
C3370 CS_BIAS.n45 GND 0.070158f
C3371 CS_BIAS.n46 GND 0.010257f
C3372 CS_BIAS.n47 GND 0.015989f
C3373 CS_BIAS.n48 GND 0.007971f
C3374 CS_BIAS.n49 GND 0.007971f
C3375 CS_BIAS.n50 GND 0.007971f
C3376 CS_BIAS.n51 GND 0.014853f
C3377 CS_BIAS.n52 GND 0.012592f
C3378 CS_BIAS.n53 GND 0.095669f
C3379 CS_BIAS.n54 GND 0.062155f
C3380 CS_BIAS.t17 GND 0.009386f
C3381 CS_BIAS.t1 GND 0.009386f
C3382 CS_BIAS.n55 GND 0.073253f
C3383 CS_BIAS.n56 GND 0.102116f
C3384 CS_BIAS.t21 GND 0.009386f
C3385 CS_BIAS.t3 GND 0.009386f
C3386 CS_BIAS.n57 GND 0.073253f
C3387 CS_BIAS.t23 GND 0.009386f
C3388 CS_BIAS.t5 GND 0.009386f
C3389 CS_BIAS.n58 GND 0.075229f
C3390 CS_BIAS.n59 GND 0.185343f
C3391 CS_BIAS.n60 GND 0.007971f
C3392 CS_BIAS.t74 GND 0.172127f
C3393 CS_BIAS.n61 GND 0.006602f
C3394 CS_BIAS.n62 GND 0.06794f
C3395 CS_BIAS.t65 GND 0.172127f
C3396 CS_BIAS.t51 GND 0.222799f
C3397 CS_BIAS.n63 GND 0.087264f
C3398 CS_BIAS.n64 GND 0.091464f
C3399 CS_BIAS.n65 GND 0.012008f
C3400 CS_BIAS.n66 GND 0.015368f
C3401 CS_BIAS.n67 GND 0.007971f
C3402 CS_BIAS.n68 GND 0.007971f
C3403 CS_BIAS.n69 GND 0.007971f
C3404 CS_BIAS.n70 GND 0.015985f
C3405 CS_BIAS.n71 GND 0.010841f
C3406 CS_BIAS.n72 GND 0.070158f
C3407 CS_BIAS.n73 GND 0.011425f
C3408 CS_BIAS.n74 GND 0.007971f
C3409 CS_BIAS.n75 GND 0.007933f
C3410 CS_BIAS.n76 GND 0.05762f
C3411 CS_BIAS.n77 GND 0.006438f
C3412 CS_BIAS.n78 GND 0.015759f
C3413 CS_BIAS.n79 GND 0.011425f
C3414 CS_BIAS.n80 GND 0.007971f
C3415 CS_BIAS.n81 GND 0.007971f
C3416 CS_BIAS.n82 GND 0.010841f
C3417 CS_BIAS.n83 GND 0.015985f
C3418 CS_BIAS.n84 GND 0.006602f
C3419 CS_BIAS.n85 GND 0.007971f
C3420 CS_BIAS.n86 GND 0.007971f
C3421 CS_BIAS.n87 GND 0.007971f
C3422 CS_BIAS.n88 GND 0.012008f
C3423 CS_BIAS.n89 GND 0.070158f
C3424 CS_BIAS.n90 GND 0.010257f
C3425 CS_BIAS.n91 GND 0.015989f
C3426 CS_BIAS.n92 GND 0.007971f
C3427 CS_BIAS.n93 GND 0.007971f
C3428 CS_BIAS.n94 GND 0.007971f
C3429 CS_BIAS.n95 GND 0.014853f
C3430 CS_BIAS.n96 GND 0.012592f
C3431 CS_BIAS.n97 GND 0.095669f
C3432 CS_BIAS.n98 GND 0.041095f
C3433 CS_BIAS.n99 GND 0.010508f
C3434 CS_BIAS.t43 GND 0.172127f
C3435 CS_BIAS.n100 GND 0.007113f
C3436 CS_BIAS.n101 GND 0.007971f
C3437 CS_BIAS.t26 GND 0.172127f
C3438 CS_BIAS.n102 GND 0.015368f
C3439 CS_BIAS.n103 GND 0.007971f
C3440 CS_BIAS.t81 GND 0.172127f
C3441 CS_BIAS.n104 GND 0.070158f
C3442 CS_BIAS.n105 GND 0.007971f
C3443 CS_BIAS.n106 GND 0.015759f
C3444 CS_BIAS.n107 GND 0.007971f
C3445 CS_BIAS.t25 GND 0.172127f
C3446 CS_BIAS.n108 GND 0.006602f
C3447 CS_BIAS.n109 GND 0.06794f
C3448 CS_BIAS.t80 GND 0.172127f
C3449 CS_BIAS.t73 GND 0.222799f
C3450 CS_BIAS.n110 GND 0.087264f
C3451 CS_BIAS.n111 GND 0.091464f
C3452 CS_BIAS.n112 GND 0.012008f
C3453 CS_BIAS.n113 GND 0.015368f
C3454 CS_BIAS.n114 GND 0.007971f
C3455 CS_BIAS.n115 GND 0.007971f
C3456 CS_BIAS.n116 GND 0.007971f
C3457 CS_BIAS.n117 GND 0.015985f
C3458 CS_BIAS.n118 GND 0.010841f
C3459 CS_BIAS.n119 GND 0.070158f
C3460 CS_BIAS.n120 GND 0.011425f
C3461 CS_BIAS.n121 GND 0.007971f
C3462 CS_BIAS.n122 GND 0.007971f
C3463 CS_BIAS.n123 GND 0.007971f
C3464 CS_BIAS.n124 GND 0.006438f
C3465 CS_BIAS.n125 GND 0.015759f
C3466 CS_BIAS.n126 GND 0.011425f
C3467 CS_BIAS.n127 GND 0.007971f
C3468 CS_BIAS.n128 GND 0.007971f
C3469 CS_BIAS.n129 GND 0.010841f
C3470 CS_BIAS.n130 GND 0.015985f
C3471 CS_BIAS.n131 GND 0.006602f
C3472 CS_BIAS.n132 GND 0.007971f
C3473 CS_BIAS.n133 GND 0.007971f
C3474 CS_BIAS.n134 GND 0.007971f
C3475 CS_BIAS.n135 GND 0.012008f
C3476 CS_BIAS.n136 GND 0.070158f
C3477 CS_BIAS.n137 GND 0.010257f
C3478 CS_BIAS.n138 GND 0.015989f
C3479 CS_BIAS.n139 GND 0.007971f
C3480 CS_BIAS.n140 GND 0.007971f
C3481 CS_BIAS.n141 GND 0.007971f
C3482 CS_BIAS.n142 GND 0.014853f
C3483 CS_BIAS.n143 GND 0.012592f
C3484 CS_BIAS.n144 GND 0.095669f
C3485 CS_BIAS.n145 GND 0.030371f
C3486 CS_BIAS.n146 GND 0.086423f
C3487 CS_BIAS.n147 GND 0.010508f
C3488 CS_BIAS.t45 GND 0.172127f
C3489 CS_BIAS.n148 GND 0.007113f
C3490 CS_BIAS.n149 GND 0.007971f
C3491 CS_BIAS.t57 GND 0.172127f
C3492 CS_BIAS.n150 GND 0.015368f
C3493 CS_BIAS.n151 GND 0.007971f
C3494 CS_BIAS.t55 GND 0.172127f
C3495 CS_BIAS.n152 GND 0.070158f
C3496 CS_BIAS.n153 GND 0.007971f
C3497 CS_BIAS.n154 GND 0.015759f
C3498 CS_BIAS.n155 GND 0.007971f
C3499 CS_BIAS.t34 GND 0.172127f
C3500 CS_BIAS.n156 GND 0.006602f
C3501 CS_BIAS.n157 GND 0.06794f
C3502 CS_BIAS.t32 GND 0.172127f
C3503 CS_BIAS.t49 GND 0.222799f
C3504 CS_BIAS.n158 GND 0.087264f
C3505 CS_BIAS.n159 GND 0.091464f
C3506 CS_BIAS.n160 GND 0.012008f
C3507 CS_BIAS.n161 GND 0.015368f
C3508 CS_BIAS.n162 GND 0.007971f
C3509 CS_BIAS.n163 GND 0.007971f
C3510 CS_BIAS.n164 GND 0.007971f
C3511 CS_BIAS.n165 GND 0.015985f
C3512 CS_BIAS.n166 GND 0.010841f
C3513 CS_BIAS.n167 GND 0.070158f
C3514 CS_BIAS.n168 GND 0.011425f
C3515 CS_BIAS.n169 GND 0.007971f
C3516 CS_BIAS.n170 GND 0.007971f
C3517 CS_BIAS.n171 GND 0.007971f
C3518 CS_BIAS.n172 GND 0.006438f
C3519 CS_BIAS.n173 GND 0.015759f
C3520 CS_BIAS.n174 GND 0.011425f
C3521 CS_BIAS.n175 GND 0.007971f
C3522 CS_BIAS.n176 GND 0.007971f
C3523 CS_BIAS.n177 GND 0.010841f
C3524 CS_BIAS.n178 GND 0.015985f
C3525 CS_BIAS.n179 GND 0.006602f
C3526 CS_BIAS.n180 GND 0.007971f
C3527 CS_BIAS.n181 GND 0.007971f
C3528 CS_BIAS.n182 GND 0.007971f
C3529 CS_BIAS.n183 GND 0.012008f
C3530 CS_BIAS.n184 GND 0.070158f
C3531 CS_BIAS.n185 GND 0.010257f
C3532 CS_BIAS.n186 GND 0.015989f
C3533 CS_BIAS.n187 GND 0.007971f
C3534 CS_BIAS.n188 GND 0.007971f
C3535 CS_BIAS.n189 GND 0.007971f
C3536 CS_BIAS.n190 GND 0.014853f
C3537 CS_BIAS.n191 GND 0.012592f
C3538 CS_BIAS.n192 GND 0.095669f
C3539 CS_BIAS.n193 GND 0.030371f
C3540 CS_BIAS.n194 GND 0.062469f
C3541 CS_BIAS.n195 GND 0.010508f
C3542 CS_BIAS.t78 GND 0.172127f
C3543 CS_BIAS.n196 GND 0.007113f
C3544 CS_BIAS.n197 GND 0.007971f
C3545 CS_BIAS.t30 GND 0.172127f
C3546 CS_BIAS.n198 GND 0.015368f
C3547 CS_BIAS.n199 GND 0.007971f
C3548 CS_BIAS.t31 GND 0.172127f
C3549 CS_BIAS.n200 GND 0.070158f
C3550 CS_BIAS.n201 GND 0.007971f
C3551 CS_BIAS.n202 GND 0.015759f
C3552 CS_BIAS.n203 GND 0.007971f
C3553 CS_BIAS.t35 GND 0.172127f
C3554 CS_BIAS.n204 GND 0.006602f
C3555 CS_BIAS.n205 GND 0.06794f
C3556 CS_BIAS.t33 GND 0.172127f
C3557 CS_BIAS.t56 GND 0.222799f
C3558 CS_BIAS.n206 GND 0.087264f
C3559 CS_BIAS.n207 GND 0.091464f
C3560 CS_BIAS.n208 GND 0.012008f
C3561 CS_BIAS.n209 GND 0.015368f
C3562 CS_BIAS.n210 GND 0.007971f
C3563 CS_BIAS.n211 GND 0.007971f
C3564 CS_BIAS.n212 GND 0.007971f
C3565 CS_BIAS.n213 GND 0.015985f
C3566 CS_BIAS.n214 GND 0.010841f
C3567 CS_BIAS.n215 GND 0.070158f
C3568 CS_BIAS.n216 GND 0.011425f
C3569 CS_BIAS.n217 GND 0.007971f
C3570 CS_BIAS.n218 GND 0.007971f
C3571 CS_BIAS.n219 GND 0.007971f
C3572 CS_BIAS.n220 GND 0.006438f
C3573 CS_BIAS.n221 GND 0.015759f
C3574 CS_BIAS.n222 GND 0.011425f
C3575 CS_BIAS.n223 GND 0.007971f
C3576 CS_BIAS.n224 GND 0.007971f
C3577 CS_BIAS.n225 GND 0.010841f
C3578 CS_BIAS.n226 GND 0.015985f
C3579 CS_BIAS.n227 GND 0.006602f
C3580 CS_BIAS.n228 GND 0.007971f
C3581 CS_BIAS.n229 GND 0.007971f
C3582 CS_BIAS.n230 GND 0.007971f
C3583 CS_BIAS.n231 GND 0.012008f
C3584 CS_BIAS.n232 GND 0.070158f
C3585 CS_BIAS.n233 GND 0.010257f
C3586 CS_BIAS.n234 GND 0.015989f
C3587 CS_BIAS.n235 GND 0.007971f
C3588 CS_BIAS.n236 GND 0.007971f
C3589 CS_BIAS.n237 GND 0.007971f
C3590 CS_BIAS.n238 GND 0.014853f
C3591 CS_BIAS.n239 GND 0.012592f
C3592 CS_BIAS.n240 GND 0.095669f
C3593 CS_BIAS.n241 GND 0.030371f
C3594 CS_BIAS.n242 GND 0.062469f
C3595 CS_BIAS.n243 GND 0.010508f
C3596 CS_BIAS.t40 GND 0.172127f
C3597 CS_BIAS.n244 GND 0.007113f
C3598 CS_BIAS.n245 GND 0.007971f
C3599 CS_BIAS.t61 GND 0.172127f
C3600 CS_BIAS.n246 GND 0.015368f
C3601 CS_BIAS.n247 GND 0.007971f
C3602 CS_BIAS.t60 GND 0.172127f
C3603 CS_BIAS.n248 GND 0.070158f
C3604 CS_BIAS.n249 GND 0.007971f
C3605 CS_BIAS.n250 GND 0.015759f
C3606 CS_BIAS.n251 GND 0.007971f
C3607 CS_BIAS.t67 GND 0.172127f
C3608 CS_BIAS.n252 GND 0.006602f
C3609 CS_BIAS.n253 GND 0.06794f
C3610 CS_BIAS.t66 GND 0.172127f
C3611 CS_BIAS.t82 GND 0.222799f
C3612 CS_BIAS.n254 GND 0.087264f
C3613 CS_BIAS.n255 GND 0.091464f
C3614 CS_BIAS.n256 GND 0.012008f
C3615 CS_BIAS.n257 GND 0.015368f
C3616 CS_BIAS.n258 GND 0.007971f
C3617 CS_BIAS.n259 GND 0.007971f
C3618 CS_BIAS.n260 GND 0.007971f
C3619 CS_BIAS.n261 GND 0.015985f
C3620 CS_BIAS.n262 GND 0.010841f
C3621 CS_BIAS.n263 GND 0.070158f
C3622 CS_BIAS.n264 GND 0.011425f
C3623 CS_BIAS.n265 GND 0.007971f
C3624 CS_BIAS.n266 GND 0.007971f
C3625 CS_BIAS.n267 GND 0.007971f
C3626 CS_BIAS.n268 GND 0.006438f
C3627 CS_BIAS.n269 GND 0.015759f
C3628 CS_BIAS.n270 GND 0.011425f
C3629 CS_BIAS.n271 GND 0.007971f
C3630 CS_BIAS.n272 GND 0.007971f
C3631 CS_BIAS.n273 GND 0.010841f
C3632 CS_BIAS.n274 GND 0.015985f
C3633 CS_BIAS.n275 GND 0.006602f
C3634 CS_BIAS.n276 GND 0.007971f
C3635 CS_BIAS.n277 GND 0.007971f
C3636 CS_BIAS.n278 GND 0.007971f
C3637 CS_BIAS.n279 GND 0.012008f
C3638 CS_BIAS.n280 GND 0.070158f
C3639 CS_BIAS.n281 GND 0.010257f
C3640 CS_BIAS.n282 GND 0.015989f
C3641 CS_BIAS.n283 GND 0.007971f
C3642 CS_BIAS.n284 GND 0.007971f
C3643 CS_BIAS.n285 GND 0.007971f
C3644 CS_BIAS.n286 GND 0.014853f
C3645 CS_BIAS.n287 GND 0.012592f
C3646 CS_BIAS.n288 GND 0.095669f
C3647 CS_BIAS.n289 GND 0.030371f
C3648 CS_BIAS.n290 GND 0.291216f
C3649 CS_BIAS.n291 GND 0.010508f
C3650 CS_BIAS.t54 GND 0.172127f
C3651 CS_BIAS.n292 GND 0.007113f
C3652 CS_BIAS.n293 GND 0.007971f
C3653 CS_BIAS.t47 GND 0.172127f
C3654 CS_BIAS.n294 GND 0.015368f
C3655 CS_BIAS.n295 GND 0.007971f
C3656 CS_BIAS.t50 GND 0.172127f
C3657 CS_BIAS.n296 GND 0.070158f
C3658 CS_BIAS.n297 GND 0.007933f
C3659 CS_BIAS.n298 GND 0.015759f
C3660 CS_BIAS.n299 GND 0.007971f
C3661 CS_BIAS.t46 GND 0.172127f
C3662 CS_BIAS.n300 GND 0.006602f
C3663 CS_BIAS.n301 GND 0.06794f
C3664 CS_BIAS.t29 GND 0.172127f
C3665 CS_BIAS.t24 GND 0.222799f
C3666 CS_BIAS.n302 GND 0.087264f
C3667 CS_BIAS.n303 GND 0.091464f
C3668 CS_BIAS.n304 GND 0.012008f
C3669 CS_BIAS.n305 GND 0.015368f
C3670 CS_BIAS.n306 GND 0.007971f
C3671 CS_BIAS.n307 GND 0.007971f
C3672 CS_BIAS.n308 GND 0.007971f
C3673 CS_BIAS.n309 GND 0.015985f
C3674 CS_BIAS.n310 GND 0.010841f
C3675 CS_BIAS.n311 GND 0.070158f
C3676 CS_BIAS.n312 GND 0.011425f
C3677 CS_BIAS.n313 GND 0.007971f
C3678 CS_BIAS.n314 GND 0.007933f
C3679 CS_BIAS.t19 GND 0.009386f
C3680 CS_BIAS.t15 GND 0.009386f
C3681 CS_BIAS.n315 GND 0.075229f
C3682 CS_BIAS.t11 GND 0.009386f
C3683 CS_BIAS.t7 GND 0.009386f
C3684 CS_BIAS.n316 GND 0.073253f
C3685 CS_BIAS.n317 GND 0.010508f
C3686 CS_BIAS.t8 GND 0.172127f
C3687 CS_BIAS.n318 GND 0.007113f
C3688 CS_BIAS.n319 GND 0.007971f
C3689 CS_BIAS.t12 GND 0.172127f
C3690 CS_BIAS.n320 GND 0.015368f
C3691 CS_BIAS.n321 GND 0.007971f
C3692 CS_BIAS.t6 GND 0.172127f
C3693 CS_BIAS.n322 GND 0.070158f
C3694 CS_BIAS.n323 GND 0.007971f
C3695 CS_BIAS.n324 GND 0.015759f
C3696 CS_BIAS.n325 GND 0.007971f
C3697 CS_BIAS.t10 GND 0.172127f
C3698 CS_BIAS.n326 GND 0.006602f
C3699 CS_BIAS.n327 GND 0.06794f
C3700 CS_BIAS.t14 GND 0.172127f
C3701 CS_BIAS.t18 GND 0.222799f
C3702 CS_BIAS.n328 GND 0.087264f
C3703 CS_BIAS.n329 GND 0.091464f
C3704 CS_BIAS.n330 GND 0.012008f
C3705 CS_BIAS.n331 GND 0.015368f
C3706 CS_BIAS.n332 GND 0.007971f
C3707 CS_BIAS.n333 GND 0.007971f
C3708 CS_BIAS.n334 GND 0.007971f
C3709 CS_BIAS.n335 GND 0.015985f
C3710 CS_BIAS.n336 GND 0.010841f
C3711 CS_BIAS.n337 GND 0.070158f
C3712 CS_BIAS.n338 GND 0.011425f
C3713 CS_BIAS.n339 GND 0.007971f
C3714 CS_BIAS.n340 GND 0.007971f
C3715 CS_BIAS.n341 GND 0.007971f
C3716 CS_BIAS.n342 GND 0.006438f
C3717 CS_BIAS.n343 GND 0.015759f
C3718 CS_BIAS.n344 GND 0.011425f
C3719 CS_BIAS.n345 GND 0.007971f
C3720 CS_BIAS.n346 GND 0.007971f
C3721 CS_BIAS.n347 GND 0.010841f
C3722 CS_BIAS.n348 GND 0.015985f
C3723 CS_BIAS.n349 GND 0.006602f
C3724 CS_BIAS.n350 GND 0.007971f
C3725 CS_BIAS.n351 GND 0.007971f
C3726 CS_BIAS.n352 GND 0.007971f
C3727 CS_BIAS.n353 GND 0.012008f
C3728 CS_BIAS.n354 GND 0.070158f
C3729 CS_BIAS.n355 GND 0.010257f
C3730 CS_BIAS.n356 GND 0.015989f
C3731 CS_BIAS.n357 GND 0.007971f
C3732 CS_BIAS.n358 GND 0.007971f
C3733 CS_BIAS.n359 GND 0.007971f
C3734 CS_BIAS.n360 GND 0.014853f
C3735 CS_BIAS.n361 GND 0.012592f
C3736 CS_BIAS.n362 GND 0.095669f
C3737 CS_BIAS.n363 GND 0.062155f
C3738 CS_BIAS.t13 GND 0.009386f
C3739 CS_BIAS.t9 GND 0.009386f
C3740 CS_BIAS.n364 GND 0.073253f
C3741 CS_BIAS.n365 GND 0.102116f
C3742 CS_BIAS.n366 GND 0.185343f
C3743 CS_BIAS.n367 GND 0.05762f
C3744 CS_BIAS.n368 GND 0.006438f
C3745 CS_BIAS.n369 GND 0.015759f
C3746 CS_BIAS.n370 GND 0.011425f
C3747 CS_BIAS.n371 GND 0.007971f
C3748 CS_BIAS.n372 GND 0.007971f
C3749 CS_BIAS.n373 GND 0.010841f
C3750 CS_BIAS.n374 GND 0.015985f
C3751 CS_BIAS.n375 GND 0.006602f
C3752 CS_BIAS.n376 GND 0.007971f
C3753 CS_BIAS.n377 GND 0.007971f
C3754 CS_BIAS.n378 GND 0.007971f
C3755 CS_BIAS.n379 GND 0.012008f
C3756 CS_BIAS.n380 GND 0.070158f
C3757 CS_BIAS.n381 GND 0.010257f
C3758 CS_BIAS.n382 GND 0.015989f
C3759 CS_BIAS.n383 GND 0.007971f
C3760 CS_BIAS.n384 GND 0.007971f
C3761 CS_BIAS.n385 GND 0.007971f
C3762 CS_BIAS.n386 GND 0.014853f
C3763 CS_BIAS.n387 GND 0.012592f
C3764 CS_BIAS.n388 GND 0.095669f
C3765 CS_BIAS.n389 GND 0.041095f
C3766 CS_BIAS.n390 GND 0.010508f
C3767 CS_BIAS.t77 GND 0.172127f
C3768 CS_BIAS.n391 GND 0.007113f
C3769 CS_BIAS.n392 GND 0.007971f
C3770 CS_BIAS.t68 GND 0.172127f
C3771 CS_BIAS.n393 GND 0.015368f
C3772 CS_BIAS.n394 GND 0.007971f
C3773 CS_BIAS.t72 GND 0.172127f
C3774 CS_BIAS.n395 GND 0.070158f
C3775 CS_BIAS.n396 GND 0.007971f
C3776 CS_BIAS.n397 GND 0.015759f
C3777 CS_BIAS.n398 GND 0.007971f
C3778 CS_BIAS.t62 GND 0.172127f
C3779 CS_BIAS.n399 GND 0.006602f
C3780 CS_BIAS.n400 GND 0.06794f
C3781 CS_BIAS.t48 GND 0.172127f
C3782 CS_BIAS.t44 GND 0.222799f
C3783 CS_BIAS.n401 GND 0.087264f
C3784 CS_BIAS.n402 GND 0.091464f
C3785 CS_BIAS.n403 GND 0.012008f
C3786 CS_BIAS.n404 GND 0.015368f
C3787 CS_BIAS.n405 GND 0.007971f
C3788 CS_BIAS.n406 GND 0.007971f
C3789 CS_BIAS.n407 GND 0.007971f
C3790 CS_BIAS.n408 GND 0.015985f
C3791 CS_BIAS.n409 GND 0.010841f
C3792 CS_BIAS.n410 GND 0.070158f
C3793 CS_BIAS.n411 GND 0.011425f
C3794 CS_BIAS.n412 GND 0.007971f
C3795 CS_BIAS.n413 GND 0.007971f
C3796 CS_BIAS.n414 GND 0.007971f
C3797 CS_BIAS.n415 GND 0.006438f
C3798 CS_BIAS.n416 GND 0.015759f
C3799 CS_BIAS.n417 GND 0.011425f
C3800 CS_BIAS.n418 GND 0.007971f
C3801 CS_BIAS.n419 GND 0.007971f
C3802 CS_BIAS.n420 GND 0.010841f
C3803 CS_BIAS.n421 GND 0.015985f
C3804 CS_BIAS.n422 GND 0.006602f
C3805 CS_BIAS.n423 GND 0.007971f
C3806 CS_BIAS.n424 GND 0.007971f
C3807 CS_BIAS.n425 GND 0.007971f
C3808 CS_BIAS.n426 GND 0.012008f
C3809 CS_BIAS.n427 GND 0.070158f
C3810 CS_BIAS.n428 GND 0.010257f
C3811 CS_BIAS.n429 GND 0.015989f
C3812 CS_BIAS.n430 GND 0.007971f
C3813 CS_BIAS.n431 GND 0.007971f
C3814 CS_BIAS.n432 GND 0.007971f
C3815 CS_BIAS.n433 GND 0.014853f
C3816 CS_BIAS.n434 GND 0.012592f
C3817 CS_BIAS.n435 GND 0.095669f
C3818 CS_BIAS.n436 GND 0.030371f
C3819 CS_BIAS.n437 GND 0.086423f
C3820 CS_BIAS.n438 GND 0.010508f
C3821 CS_BIAS.t59 GND 0.172127f
C3822 CS_BIAS.n439 GND 0.007113f
C3823 CS_BIAS.n440 GND 0.007971f
C3824 CS_BIAS.t58 GND 0.172127f
C3825 CS_BIAS.n441 GND 0.015368f
C3826 CS_BIAS.n442 GND 0.007971f
C3827 CS_BIAS.t39 GND 0.172127f
C3828 CS_BIAS.n443 GND 0.070158f
C3829 CS_BIAS.n444 GND 0.007971f
C3830 CS_BIAS.n445 GND 0.015759f
C3831 CS_BIAS.n446 GND 0.007971f
C3832 CS_BIAS.t37 GND 0.172127f
C3833 CS_BIAS.n447 GND 0.006602f
C3834 CS_BIAS.n448 GND 0.06794f
C3835 CS_BIAS.t53 GND 0.172127f
C3836 CS_BIAS.t52 GND 0.222799f
C3837 CS_BIAS.n449 GND 0.087264f
C3838 CS_BIAS.n450 GND 0.091464f
C3839 CS_BIAS.n451 GND 0.012008f
C3840 CS_BIAS.n452 GND 0.015368f
C3841 CS_BIAS.n453 GND 0.007971f
C3842 CS_BIAS.n454 GND 0.007971f
C3843 CS_BIAS.n455 GND 0.007971f
C3844 CS_BIAS.n456 GND 0.015985f
C3845 CS_BIAS.n457 GND 0.010841f
C3846 CS_BIAS.n458 GND 0.070158f
C3847 CS_BIAS.n459 GND 0.011425f
C3848 CS_BIAS.n460 GND 0.007971f
C3849 CS_BIAS.n461 GND 0.007971f
C3850 CS_BIAS.n462 GND 0.007971f
C3851 CS_BIAS.n463 GND 0.006438f
C3852 CS_BIAS.n464 GND 0.015759f
C3853 CS_BIAS.n465 GND 0.011425f
C3854 CS_BIAS.n466 GND 0.007971f
C3855 CS_BIAS.n467 GND 0.007971f
C3856 CS_BIAS.n468 GND 0.010841f
C3857 CS_BIAS.n469 GND 0.015985f
C3858 CS_BIAS.n470 GND 0.006602f
C3859 CS_BIAS.n471 GND 0.007971f
C3860 CS_BIAS.n472 GND 0.007971f
C3861 CS_BIAS.n473 GND 0.007971f
C3862 CS_BIAS.n474 GND 0.012008f
C3863 CS_BIAS.n475 GND 0.070158f
C3864 CS_BIAS.n476 GND 0.010257f
C3865 CS_BIAS.n477 GND 0.015989f
C3866 CS_BIAS.n478 GND 0.007971f
C3867 CS_BIAS.n479 GND 0.007971f
C3868 CS_BIAS.n480 GND 0.007971f
C3869 CS_BIAS.n481 GND 0.014853f
C3870 CS_BIAS.n482 GND 0.012592f
C3871 CS_BIAS.n483 GND 0.095669f
C3872 CS_BIAS.n484 GND 0.030371f
C3873 CS_BIAS.n485 GND 0.062469f
C3874 CS_BIAS.n486 GND 0.010508f
C3875 CS_BIAS.t38 GND 0.172127f
C3876 CS_BIAS.n487 GND 0.007113f
C3877 CS_BIAS.n488 GND 0.007971f
C3878 CS_BIAS.t36 GND 0.172127f
C3879 CS_BIAS.n489 GND 0.015368f
C3880 CS_BIAS.n490 GND 0.007971f
C3881 CS_BIAS.t42 GND 0.172127f
C3882 CS_BIAS.n491 GND 0.070158f
C3883 CS_BIAS.n492 GND 0.007971f
C3884 CS_BIAS.n493 GND 0.015759f
C3885 CS_BIAS.n494 GND 0.007971f
C3886 CS_BIAS.t41 GND 0.172127f
C3887 CS_BIAS.n495 GND 0.006602f
C3888 CS_BIAS.n496 GND 0.06794f
C3889 CS_BIAS.t64 GND 0.172127f
C3890 CS_BIAS.t63 GND 0.222799f
C3891 CS_BIAS.n497 GND 0.087264f
C3892 CS_BIAS.n498 GND 0.091464f
C3893 CS_BIAS.n499 GND 0.012008f
C3894 CS_BIAS.n500 GND 0.015368f
C3895 CS_BIAS.n501 GND 0.007971f
C3896 CS_BIAS.n502 GND 0.007971f
C3897 CS_BIAS.n503 GND 0.007971f
C3898 CS_BIAS.n504 GND 0.015985f
C3899 CS_BIAS.n505 GND 0.010841f
C3900 CS_BIAS.n506 GND 0.070158f
C3901 CS_BIAS.n507 GND 0.011425f
C3902 CS_BIAS.n508 GND 0.007971f
C3903 CS_BIAS.n509 GND 0.007971f
C3904 CS_BIAS.n510 GND 0.007971f
C3905 CS_BIAS.n511 GND 0.006438f
C3906 CS_BIAS.n512 GND 0.015759f
C3907 CS_BIAS.n513 GND 0.011425f
C3908 CS_BIAS.n514 GND 0.007971f
C3909 CS_BIAS.n515 GND 0.007971f
C3910 CS_BIAS.n516 GND 0.010841f
C3911 CS_BIAS.n517 GND 0.015985f
C3912 CS_BIAS.n518 GND 0.006602f
C3913 CS_BIAS.n519 GND 0.007971f
C3914 CS_BIAS.n520 GND 0.007971f
C3915 CS_BIAS.n521 GND 0.007971f
C3916 CS_BIAS.n522 GND 0.012008f
C3917 CS_BIAS.n523 GND 0.070158f
C3918 CS_BIAS.n524 GND 0.010257f
C3919 CS_BIAS.n525 GND 0.015989f
C3920 CS_BIAS.n526 GND 0.007971f
C3921 CS_BIAS.n527 GND 0.007971f
C3922 CS_BIAS.n528 GND 0.007971f
C3923 CS_BIAS.n529 GND 0.014853f
C3924 CS_BIAS.n530 GND 0.012592f
C3925 CS_BIAS.n531 GND 0.095669f
C3926 CS_BIAS.n532 GND 0.030371f
C3927 CS_BIAS.n533 GND 0.062469f
C3928 CS_BIAS.n534 GND 0.010508f
C3929 CS_BIAS.t69 GND 0.172127f
C3930 CS_BIAS.n535 GND 0.007113f
C3931 CS_BIAS.n536 GND 0.007971f
C3932 CS_BIAS.t70 GND 0.172127f
C3933 CS_BIAS.n537 GND 0.015368f
C3934 CS_BIAS.n538 GND 0.007971f
C3935 CS_BIAS.t75 GND 0.172127f
C3936 CS_BIAS.n539 GND 0.070158f
C3937 CS_BIAS.n540 GND 0.007971f
C3938 CS_BIAS.n541 GND 0.015759f
C3939 CS_BIAS.n542 GND 0.007971f
C3940 CS_BIAS.t76 GND 0.172127f
C3941 CS_BIAS.n543 GND 0.006602f
C3942 CS_BIAS.n544 GND 0.06794f
C3943 CS_BIAS.t28 GND 0.172127f
C3944 CS_BIAS.t27 GND 0.222799f
C3945 CS_BIAS.n545 GND 0.087264f
C3946 CS_BIAS.n546 GND 0.091464f
C3947 CS_BIAS.n547 GND 0.012008f
C3948 CS_BIAS.n548 GND 0.015368f
C3949 CS_BIAS.n549 GND 0.007971f
C3950 CS_BIAS.n550 GND 0.007971f
C3951 CS_BIAS.n551 GND 0.007971f
C3952 CS_BIAS.n552 GND 0.015985f
C3953 CS_BIAS.n553 GND 0.010841f
C3954 CS_BIAS.n554 GND 0.070158f
C3955 CS_BIAS.n555 GND 0.011425f
C3956 CS_BIAS.n556 GND 0.007971f
C3957 CS_BIAS.n557 GND 0.007971f
C3958 CS_BIAS.n558 GND 0.007971f
C3959 CS_BIAS.n559 GND 0.006438f
C3960 CS_BIAS.n560 GND 0.015759f
C3961 CS_BIAS.n561 GND 0.011425f
C3962 CS_BIAS.n562 GND 0.007971f
C3963 CS_BIAS.n563 GND 0.007971f
C3964 CS_BIAS.n564 GND 0.010841f
C3965 CS_BIAS.n565 GND 0.015985f
C3966 CS_BIAS.n566 GND 0.006602f
C3967 CS_BIAS.n567 GND 0.007971f
C3968 CS_BIAS.n568 GND 0.007971f
C3969 CS_BIAS.n569 GND 0.007971f
C3970 CS_BIAS.n570 GND 0.012008f
C3971 CS_BIAS.n571 GND 0.070158f
C3972 CS_BIAS.n572 GND 0.010257f
C3973 CS_BIAS.n573 GND 0.015989f
C3974 CS_BIAS.n574 GND 0.007971f
C3975 CS_BIAS.n575 GND 0.007971f
C3976 CS_BIAS.n576 GND 0.007971f
C3977 CS_BIAS.n577 GND 0.014853f
C3978 CS_BIAS.n578 GND 0.012592f
C3979 CS_BIAS.n579 GND 0.095669f
C3980 CS_BIAS.n580 GND 0.030371f
C3981 CS_BIAS.n581 GND 0.1276f
C3982 CS_BIAS.n582 GND 4.77864f
.ends

