* NGSPICE file created from diff_pair_sample_1589.ext - technology: sky130A

.subckt diff_pair_sample_1589 VTAIL VN VP B VDD2 VDD1
X0 B.t19 B.t17 B.t18 B.t11 sky130_fd_pr__nfet_01v8 ad=5.4873 pd=28.92 as=0 ps=0 w=14.07 l=3.71
X1 B.t16 B.t14 B.t15 B.t7 sky130_fd_pr__nfet_01v8 ad=5.4873 pd=28.92 as=0 ps=0 w=14.07 l=3.71
X2 VDD1.t5 VP.t0 VTAIL.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=5.4873 pd=28.92 as=2.32155 ps=14.4 w=14.07 l=3.71
X3 VDD2.t5 VN.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.32155 pd=14.4 as=5.4873 ps=28.92 w=14.07 l=3.71
X4 VTAIL.t6 VP.t1 VDD1.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=2.32155 pd=14.4 as=2.32155 ps=14.4 w=14.07 l=3.71
X5 VDD1.t3 VP.t2 VTAIL.t7 B.t0 sky130_fd_pr__nfet_01v8 ad=2.32155 pd=14.4 as=5.4873 ps=28.92 w=14.07 l=3.71
X6 VTAIL.t3 VN.t1 VDD2.t4 B.t5 sky130_fd_pr__nfet_01v8 ad=2.32155 pd=14.4 as=2.32155 ps=14.4 w=14.07 l=3.71
X7 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=5.4873 pd=28.92 as=0 ps=0 w=14.07 l=3.71
X8 VTAIL.t4 VN.t2 VDD2.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.32155 pd=14.4 as=2.32155 ps=14.4 w=14.07 l=3.71
X9 VDD2.t2 VN.t3 VTAIL.t11 B.t4 sky130_fd_pr__nfet_01v8 ad=2.32155 pd=14.4 as=5.4873 ps=28.92 w=14.07 l=3.71
X10 VTAIL.t8 VP.t3 VDD1.t2 B.t5 sky130_fd_pr__nfet_01v8 ad=2.32155 pd=14.4 as=2.32155 ps=14.4 w=14.07 l=3.71
X11 VDD2.t1 VN.t4 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=5.4873 pd=28.92 as=2.32155 ps=14.4 w=14.07 l=3.71
X12 VDD1.t1 VP.t4 VTAIL.t10 B.t2 sky130_fd_pr__nfet_01v8 ad=5.4873 pd=28.92 as=2.32155 ps=14.4 w=14.07 l=3.71
X13 VDD1.t0 VP.t5 VTAIL.t9 B.t4 sky130_fd_pr__nfet_01v8 ad=2.32155 pd=14.4 as=5.4873 ps=28.92 w=14.07 l=3.71
X14 VDD2.t0 VN.t5 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=5.4873 pd=28.92 as=2.32155 ps=14.4 w=14.07 l=3.71
X15 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=5.4873 pd=28.92 as=0 ps=0 w=14.07 l=3.71
R0 B.n979 B.n978 585
R1 B.n980 B.n979 585
R2 B.n365 B.n155 585
R3 B.n364 B.n363 585
R4 B.n362 B.n361 585
R5 B.n360 B.n359 585
R6 B.n358 B.n357 585
R7 B.n356 B.n355 585
R8 B.n354 B.n353 585
R9 B.n352 B.n351 585
R10 B.n350 B.n349 585
R11 B.n348 B.n347 585
R12 B.n346 B.n345 585
R13 B.n344 B.n343 585
R14 B.n342 B.n341 585
R15 B.n340 B.n339 585
R16 B.n338 B.n337 585
R17 B.n336 B.n335 585
R18 B.n334 B.n333 585
R19 B.n332 B.n331 585
R20 B.n330 B.n329 585
R21 B.n328 B.n327 585
R22 B.n326 B.n325 585
R23 B.n324 B.n323 585
R24 B.n322 B.n321 585
R25 B.n320 B.n319 585
R26 B.n318 B.n317 585
R27 B.n316 B.n315 585
R28 B.n314 B.n313 585
R29 B.n312 B.n311 585
R30 B.n310 B.n309 585
R31 B.n308 B.n307 585
R32 B.n306 B.n305 585
R33 B.n304 B.n303 585
R34 B.n302 B.n301 585
R35 B.n300 B.n299 585
R36 B.n298 B.n297 585
R37 B.n296 B.n295 585
R38 B.n294 B.n293 585
R39 B.n292 B.n291 585
R40 B.n290 B.n289 585
R41 B.n288 B.n287 585
R42 B.n286 B.n285 585
R43 B.n284 B.n283 585
R44 B.n282 B.n281 585
R45 B.n280 B.n279 585
R46 B.n278 B.n277 585
R47 B.n276 B.n275 585
R48 B.n274 B.n273 585
R49 B.n271 B.n270 585
R50 B.n269 B.n268 585
R51 B.n267 B.n266 585
R52 B.n265 B.n264 585
R53 B.n263 B.n262 585
R54 B.n261 B.n260 585
R55 B.n259 B.n258 585
R56 B.n257 B.n256 585
R57 B.n255 B.n254 585
R58 B.n253 B.n252 585
R59 B.n251 B.n250 585
R60 B.n249 B.n248 585
R61 B.n247 B.n246 585
R62 B.n245 B.n244 585
R63 B.n243 B.n242 585
R64 B.n241 B.n240 585
R65 B.n239 B.n238 585
R66 B.n237 B.n236 585
R67 B.n235 B.n234 585
R68 B.n233 B.n232 585
R69 B.n231 B.n230 585
R70 B.n229 B.n228 585
R71 B.n227 B.n226 585
R72 B.n225 B.n224 585
R73 B.n223 B.n222 585
R74 B.n221 B.n220 585
R75 B.n219 B.n218 585
R76 B.n217 B.n216 585
R77 B.n215 B.n214 585
R78 B.n213 B.n212 585
R79 B.n211 B.n210 585
R80 B.n209 B.n208 585
R81 B.n207 B.n206 585
R82 B.n205 B.n204 585
R83 B.n203 B.n202 585
R84 B.n201 B.n200 585
R85 B.n199 B.n198 585
R86 B.n197 B.n196 585
R87 B.n195 B.n194 585
R88 B.n193 B.n192 585
R89 B.n191 B.n190 585
R90 B.n189 B.n188 585
R91 B.n187 B.n186 585
R92 B.n185 B.n184 585
R93 B.n183 B.n182 585
R94 B.n181 B.n180 585
R95 B.n179 B.n178 585
R96 B.n177 B.n176 585
R97 B.n175 B.n174 585
R98 B.n173 B.n172 585
R99 B.n171 B.n170 585
R100 B.n169 B.n168 585
R101 B.n167 B.n166 585
R102 B.n165 B.n164 585
R103 B.n163 B.n162 585
R104 B.n103 B.n102 585
R105 B.n983 B.n982 585
R106 B.n977 B.n156 585
R107 B.n156 B.n100 585
R108 B.n976 B.n99 585
R109 B.n987 B.n99 585
R110 B.n975 B.n98 585
R111 B.n988 B.n98 585
R112 B.n974 B.n97 585
R113 B.n989 B.n97 585
R114 B.n973 B.n972 585
R115 B.n972 B.n93 585
R116 B.n971 B.n92 585
R117 B.n995 B.n92 585
R118 B.n970 B.n91 585
R119 B.n996 B.n91 585
R120 B.n969 B.n90 585
R121 B.n997 B.n90 585
R122 B.n968 B.n967 585
R123 B.n967 B.n86 585
R124 B.n966 B.n85 585
R125 B.n1003 B.n85 585
R126 B.n965 B.n84 585
R127 B.n1004 B.n84 585
R128 B.n964 B.n83 585
R129 B.n1005 B.n83 585
R130 B.n963 B.n962 585
R131 B.n962 B.n79 585
R132 B.n961 B.n78 585
R133 B.n1011 B.n78 585
R134 B.n960 B.n77 585
R135 B.n1012 B.n77 585
R136 B.n959 B.n76 585
R137 B.n1013 B.n76 585
R138 B.n958 B.n957 585
R139 B.n957 B.n72 585
R140 B.n956 B.n71 585
R141 B.n1019 B.n71 585
R142 B.n955 B.n70 585
R143 B.n1020 B.n70 585
R144 B.n954 B.n69 585
R145 B.n1021 B.n69 585
R146 B.n953 B.n952 585
R147 B.n952 B.n65 585
R148 B.n951 B.n64 585
R149 B.n1027 B.n64 585
R150 B.n950 B.n63 585
R151 B.n1028 B.n63 585
R152 B.n949 B.n62 585
R153 B.n1029 B.n62 585
R154 B.n948 B.n947 585
R155 B.n947 B.n61 585
R156 B.n946 B.n57 585
R157 B.n1035 B.n57 585
R158 B.n945 B.n56 585
R159 B.n1036 B.n56 585
R160 B.n944 B.n55 585
R161 B.n1037 B.n55 585
R162 B.n943 B.n942 585
R163 B.n942 B.n51 585
R164 B.n941 B.n50 585
R165 B.n1043 B.n50 585
R166 B.n940 B.n49 585
R167 B.n1044 B.n49 585
R168 B.n939 B.n48 585
R169 B.n1045 B.n48 585
R170 B.n938 B.n937 585
R171 B.n937 B.n44 585
R172 B.n936 B.n43 585
R173 B.n1051 B.n43 585
R174 B.n935 B.n42 585
R175 B.n1052 B.n42 585
R176 B.n934 B.n41 585
R177 B.n1053 B.n41 585
R178 B.n933 B.n932 585
R179 B.n932 B.n40 585
R180 B.n931 B.n36 585
R181 B.n1059 B.n36 585
R182 B.n930 B.n35 585
R183 B.n1060 B.n35 585
R184 B.n929 B.n34 585
R185 B.n1061 B.n34 585
R186 B.n928 B.n927 585
R187 B.n927 B.n30 585
R188 B.n926 B.n29 585
R189 B.n1067 B.n29 585
R190 B.n925 B.n28 585
R191 B.n1068 B.n28 585
R192 B.n924 B.n27 585
R193 B.n1069 B.n27 585
R194 B.n923 B.n922 585
R195 B.n922 B.n23 585
R196 B.n921 B.n22 585
R197 B.n1075 B.n22 585
R198 B.n920 B.n21 585
R199 B.n1076 B.n21 585
R200 B.n919 B.n20 585
R201 B.n1077 B.n20 585
R202 B.n918 B.n917 585
R203 B.n917 B.n16 585
R204 B.n916 B.n15 585
R205 B.n1083 B.n15 585
R206 B.n915 B.n14 585
R207 B.n1084 B.n14 585
R208 B.n914 B.n13 585
R209 B.n1085 B.n13 585
R210 B.n913 B.n912 585
R211 B.n912 B.n12 585
R212 B.n911 B.n910 585
R213 B.n911 B.n8 585
R214 B.n909 B.n7 585
R215 B.n1092 B.n7 585
R216 B.n908 B.n6 585
R217 B.n1093 B.n6 585
R218 B.n907 B.n5 585
R219 B.n1094 B.n5 585
R220 B.n906 B.n905 585
R221 B.n905 B.n4 585
R222 B.n904 B.n366 585
R223 B.n904 B.n903 585
R224 B.n894 B.n367 585
R225 B.n368 B.n367 585
R226 B.n896 B.n895 585
R227 B.n897 B.n896 585
R228 B.n893 B.n373 585
R229 B.n373 B.n372 585
R230 B.n892 B.n891 585
R231 B.n891 B.n890 585
R232 B.n375 B.n374 585
R233 B.n376 B.n375 585
R234 B.n883 B.n882 585
R235 B.n884 B.n883 585
R236 B.n881 B.n381 585
R237 B.n381 B.n380 585
R238 B.n880 B.n879 585
R239 B.n879 B.n878 585
R240 B.n383 B.n382 585
R241 B.n384 B.n383 585
R242 B.n871 B.n870 585
R243 B.n872 B.n871 585
R244 B.n869 B.n389 585
R245 B.n389 B.n388 585
R246 B.n868 B.n867 585
R247 B.n867 B.n866 585
R248 B.n391 B.n390 585
R249 B.n392 B.n391 585
R250 B.n859 B.n858 585
R251 B.n860 B.n859 585
R252 B.n857 B.n397 585
R253 B.n397 B.n396 585
R254 B.n856 B.n855 585
R255 B.n855 B.n854 585
R256 B.n399 B.n398 585
R257 B.n847 B.n399 585
R258 B.n846 B.n845 585
R259 B.n848 B.n846 585
R260 B.n844 B.n404 585
R261 B.n404 B.n403 585
R262 B.n843 B.n842 585
R263 B.n842 B.n841 585
R264 B.n406 B.n405 585
R265 B.n407 B.n406 585
R266 B.n834 B.n833 585
R267 B.n835 B.n834 585
R268 B.n832 B.n412 585
R269 B.n412 B.n411 585
R270 B.n831 B.n830 585
R271 B.n830 B.n829 585
R272 B.n414 B.n413 585
R273 B.n415 B.n414 585
R274 B.n822 B.n821 585
R275 B.n823 B.n822 585
R276 B.n820 B.n420 585
R277 B.n420 B.n419 585
R278 B.n819 B.n818 585
R279 B.n818 B.n817 585
R280 B.n422 B.n421 585
R281 B.n810 B.n422 585
R282 B.n809 B.n808 585
R283 B.n811 B.n809 585
R284 B.n807 B.n427 585
R285 B.n427 B.n426 585
R286 B.n806 B.n805 585
R287 B.n805 B.n804 585
R288 B.n429 B.n428 585
R289 B.n430 B.n429 585
R290 B.n797 B.n796 585
R291 B.n798 B.n797 585
R292 B.n795 B.n435 585
R293 B.n435 B.n434 585
R294 B.n794 B.n793 585
R295 B.n793 B.n792 585
R296 B.n437 B.n436 585
R297 B.n438 B.n437 585
R298 B.n785 B.n784 585
R299 B.n786 B.n785 585
R300 B.n783 B.n443 585
R301 B.n443 B.n442 585
R302 B.n782 B.n781 585
R303 B.n781 B.n780 585
R304 B.n445 B.n444 585
R305 B.n446 B.n445 585
R306 B.n773 B.n772 585
R307 B.n774 B.n773 585
R308 B.n771 B.n451 585
R309 B.n451 B.n450 585
R310 B.n770 B.n769 585
R311 B.n769 B.n768 585
R312 B.n453 B.n452 585
R313 B.n454 B.n453 585
R314 B.n761 B.n760 585
R315 B.n762 B.n761 585
R316 B.n759 B.n459 585
R317 B.n459 B.n458 585
R318 B.n758 B.n757 585
R319 B.n757 B.n756 585
R320 B.n461 B.n460 585
R321 B.n462 B.n461 585
R322 B.n749 B.n748 585
R323 B.n750 B.n749 585
R324 B.n747 B.n467 585
R325 B.n467 B.n466 585
R326 B.n746 B.n745 585
R327 B.n745 B.n744 585
R328 B.n469 B.n468 585
R329 B.n470 B.n469 585
R330 B.n740 B.n739 585
R331 B.n473 B.n472 585
R332 B.n736 B.n735 585
R333 B.n737 B.n736 585
R334 B.n734 B.n525 585
R335 B.n733 B.n732 585
R336 B.n731 B.n730 585
R337 B.n729 B.n728 585
R338 B.n727 B.n726 585
R339 B.n725 B.n724 585
R340 B.n723 B.n722 585
R341 B.n721 B.n720 585
R342 B.n719 B.n718 585
R343 B.n717 B.n716 585
R344 B.n715 B.n714 585
R345 B.n713 B.n712 585
R346 B.n711 B.n710 585
R347 B.n709 B.n708 585
R348 B.n707 B.n706 585
R349 B.n705 B.n704 585
R350 B.n703 B.n702 585
R351 B.n701 B.n700 585
R352 B.n699 B.n698 585
R353 B.n697 B.n696 585
R354 B.n695 B.n694 585
R355 B.n693 B.n692 585
R356 B.n691 B.n690 585
R357 B.n689 B.n688 585
R358 B.n687 B.n686 585
R359 B.n685 B.n684 585
R360 B.n683 B.n682 585
R361 B.n681 B.n680 585
R362 B.n679 B.n678 585
R363 B.n677 B.n676 585
R364 B.n675 B.n674 585
R365 B.n673 B.n672 585
R366 B.n671 B.n670 585
R367 B.n669 B.n668 585
R368 B.n667 B.n666 585
R369 B.n665 B.n664 585
R370 B.n663 B.n662 585
R371 B.n661 B.n660 585
R372 B.n659 B.n658 585
R373 B.n657 B.n656 585
R374 B.n655 B.n654 585
R375 B.n653 B.n652 585
R376 B.n651 B.n650 585
R377 B.n649 B.n648 585
R378 B.n647 B.n646 585
R379 B.n644 B.n643 585
R380 B.n642 B.n641 585
R381 B.n640 B.n639 585
R382 B.n638 B.n637 585
R383 B.n636 B.n635 585
R384 B.n634 B.n633 585
R385 B.n632 B.n631 585
R386 B.n630 B.n629 585
R387 B.n628 B.n627 585
R388 B.n626 B.n625 585
R389 B.n624 B.n623 585
R390 B.n622 B.n621 585
R391 B.n620 B.n619 585
R392 B.n618 B.n617 585
R393 B.n616 B.n615 585
R394 B.n614 B.n613 585
R395 B.n612 B.n611 585
R396 B.n610 B.n609 585
R397 B.n608 B.n607 585
R398 B.n606 B.n605 585
R399 B.n604 B.n603 585
R400 B.n602 B.n601 585
R401 B.n600 B.n599 585
R402 B.n598 B.n597 585
R403 B.n596 B.n595 585
R404 B.n594 B.n593 585
R405 B.n592 B.n591 585
R406 B.n590 B.n589 585
R407 B.n588 B.n587 585
R408 B.n586 B.n585 585
R409 B.n584 B.n583 585
R410 B.n582 B.n581 585
R411 B.n580 B.n579 585
R412 B.n578 B.n577 585
R413 B.n576 B.n575 585
R414 B.n574 B.n573 585
R415 B.n572 B.n571 585
R416 B.n570 B.n569 585
R417 B.n568 B.n567 585
R418 B.n566 B.n565 585
R419 B.n564 B.n563 585
R420 B.n562 B.n561 585
R421 B.n560 B.n559 585
R422 B.n558 B.n557 585
R423 B.n556 B.n555 585
R424 B.n554 B.n553 585
R425 B.n552 B.n551 585
R426 B.n550 B.n549 585
R427 B.n548 B.n547 585
R428 B.n546 B.n545 585
R429 B.n544 B.n543 585
R430 B.n542 B.n541 585
R431 B.n540 B.n539 585
R432 B.n538 B.n537 585
R433 B.n536 B.n535 585
R434 B.n534 B.n533 585
R435 B.n532 B.n531 585
R436 B.n741 B.n471 585
R437 B.n471 B.n470 585
R438 B.n743 B.n742 585
R439 B.n744 B.n743 585
R440 B.n465 B.n464 585
R441 B.n466 B.n465 585
R442 B.n752 B.n751 585
R443 B.n751 B.n750 585
R444 B.n753 B.n463 585
R445 B.n463 B.n462 585
R446 B.n755 B.n754 585
R447 B.n756 B.n755 585
R448 B.n457 B.n456 585
R449 B.n458 B.n457 585
R450 B.n764 B.n763 585
R451 B.n763 B.n762 585
R452 B.n765 B.n455 585
R453 B.n455 B.n454 585
R454 B.n767 B.n766 585
R455 B.n768 B.n767 585
R456 B.n449 B.n448 585
R457 B.n450 B.n449 585
R458 B.n776 B.n775 585
R459 B.n775 B.n774 585
R460 B.n777 B.n447 585
R461 B.n447 B.n446 585
R462 B.n779 B.n778 585
R463 B.n780 B.n779 585
R464 B.n441 B.n440 585
R465 B.n442 B.n441 585
R466 B.n788 B.n787 585
R467 B.n787 B.n786 585
R468 B.n789 B.n439 585
R469 B.n439 B.n438 585
R470 B.n791 B.n790 585
R471 B.n792 B.n791 585
R472 B.n433 B.n432 585
R473 B.n434 B.n433 585
R474 B.n800 B.n799 585
R475 B.n799 B.n798 585
R476 B.n801 B.n431 585
R477 B.n431 B.n430 585
R478 B.n803 B.n802 585
R479 B.n804 B.n803 585
R480 B.n425 B.n424 585
R481 B.n426 B.n425 585
R482 B.n813 B.n812 585
R483 B.n812 B.n811 585
R484 B.n814 B.n423 585
R485 B.n810 B.n423 585
R486 B.n816 B.n815 585
R487 B.n817 B.n816 585
R488 B.n418 B.n417 585
R489 B.n419 B.n418 585
R490 B.n825 B.n824 585
R491 B.n824 B.n823 585
R492 B.n826 B.n416 585
R493 B.n416 B.n415 585
R494 B.n828 B.n827 585
R495 B.n829 B.n828 585
R496 B.n410 B.n409 585
R497 B.n411 B.n410 585
R498 B.n837 B.n836 585
R499 B.n836 B.n835 585
R500 B.n838 B.n408 585
R501 B.n408 B.n407 585
R502 B.n840 B.n839 585
R503 B.n841 B.n840 585
R504 B.n402 B.n401 585
R505 B.n403 B.n402 585
R506 B.n850 B.n849 585
R507 B.n849 B.n848 585
R508 B.n851 B.n400 585
R509 B.n847 B.n400 585
R510 B.n853 B.n852 585
R511 B.n854 B.n853 585
R512 B.n395 B.n394 585
R513 B.n396 B.n395 585
R514 B.n862 B.n861 585
R515 B.n861 B.n860 585
R516 B.n863 B.n393 585
R517 B.n393 B.n392 585
R518 B.n865 B.n864 585
R519 B.n866 B.n865 585
R520 B.n387 B.n386 585
R521 B.n388 B.n387 585
R522 B.n874 B.n873 585
R523 B.n873 B.n872 585
R524 B.n875 B.n385 585
R525 B.n385 B.n384 585
R526 B.n877 B.n876 585
R527 B.n878 B.n877 585
R528 B.n379 B.n378 585
R529 B.n380 B.n379 585
R530 B.n886 B.n885 585
R531 B.n885 B.n884 585
R532 B.n887 B.n377 585
R533 B.n377 B.n376 585
R534 B.n889 B.n888 585
R535 B.n890 B.n889 585
R536 B.n371 B.n370 585
R537 B.n372 B.n371 585
R538 B.n899 B.n898 585
R539 B.n898 B.n897 585
R540 B.n900 B.n369 585
R541 B.n369 B.n368 585
R542 B.n902 B.n901 585
R543 B.n903 B.n902 585
R544 B.n3 B.n0 585
R545 B.n4 B.n3 585
R546 B.n1091 B.n1 585
R547 B.n1092 B.n1091 585
R548 B.n1090 B.n1089 585
R549 B.n1090 B.n8 585
R550 B.n1088 B.n9 585
R551 B.n12 B.n9 585
R552 B.n1087 B.n1086 585
R553 B.n1086 B.n1085 585
R554 B.n11 B.n10 585
R555 B.n1084 B.n11 585
R556 B.n1082 B.n1081 585
R557 B.n1083 B.n1082 585
R558 B.n1080 B.n17 585
R559 B.n17 B.n16 585
R560 B.n1079 B.n1078 585
R561 B.n1078 B.n1077 585
R562 B.n19 B.n18 585
R563 B.n1076 B.n19 585
R564 B.n1074 B.n1073 585
R565 B.n1075 B.n1074 585
R566 B.n1072 B.n24 585
R567 B.n24 B.n23 585
R568 B.n1071 B.n1070 585
R569 B.n1070 B.n1069 585
R570 B.n26 B.n25 585
R571 B.n1068 B.n26 585
R572 B.n1066 B.n1065 585
R573 B.n1067 B.n1066 585
R574 B.n1064 B.n31 585
R575 B.n31 B.n30 585
R576 B.n1063 B.n1062 585
R577 B.n1062 B.n1061 585
R578 B.n33 B.n32 585
R579 B.n1060 B.n33 585
R580 B.n1058 B.n1057 585
R581 B.n1059 B.n1058 585
R582 B.n1056 B.n37 585
R583 B.n40 B.n37 585
R584 B.n1055 B.n1054 585
R585 B.n1054 B.n1053 585
R586 B.n39 B.n38 585
R587 B.n1052 B.n39 585
R588 B.n1050 B.n1049 585
R589 B.n1051 B.n1050 585
R590 B.n1048 B.n45 585
R591 B.n45 B.n44 585
R592 B.n1047 B.n1046 585
R593 B.n1046 B.n1045 585
R594 B.n47 B.n46 585
R595 B.n1044 B.n47 585
R596 B.n1042 B.n1041 585
R597 B.n1043 B.n1042 585
R598 B.n1040 B.n52 585
R599 B.n52 B.n51 585
R600 B.n1039 B.n1038 585
R601 B.n1038 B.n1037 585
R602 B.n54 B.n53 585
R603 B.n1036 B.n54 585
R604 B.n1034 B.n1033 585
R605 B.n1035 B.n1034 585
R606 B.n1032 B.n58 585
R607 B.n61 B.n58 585
R608 B.n1031 B.n1030 585
R609 B.n1030 B.n1029 585
R610 B.n60 B.n59 585
R611 B.n1028 B.n60 585
R612 B.n1026 B.n1025 585
R613 B.n1027 B.n1026 585
R614 B.n1024 B.n66 585
R615 B.n66 B.n65 585
R616 B.n1023 B.n1022 585
R617 B.n1022 B.n1021 585
R618 B.n68 B.n67 585
R619 B.n1020 B.n68 585
R620 B.n1018 B.n1017 585
R621 B.n1019 B.n1018 585
R622 B.n1016 B.n73 585
R623 B.n73 B.n72 585
R624 B.n1015 B.n1014 585
R625 B.n1014 B.n1013 585
R626 B.n75 B.n74 585
R627 B.n1012 B.n75 585
R628 B.n1010 B.n1009 585
R629 B.n1011 B.n1010 585
R630 B.n1008 B.n80 585
R631 B.n80 B.n79 585
R632 B.n1007 B.n1006 585
R633 B.n1006 B.n1005 585
R634 B.n82 B.n81 585
R635 B.n1004 B.n82 585
R636 B.n1002 B.n1001 585
R637 B.n1003 B.n1002 585
R638 B.n1000 B.n87 585
R639 B.n87 B.n86 585
R640 B.n999 B.n998 585
R641 B.n998 B.n997 585
R642 B.n89 B.n88 585
R643 B.n996 B.n89 585
R644 B.n994 B.n993 585
R645 B.n995 B.n994 585
R646 B.n992 B.n94 585
R647 B.n94 B.n93 585
R648 B.n991 B.n990 585
R649 B.n990 B.n989 585
R650 B.n96 B.n95 585
R651 B.n988 B.n96 585
R652 B.n986 B.n985 585
R653 B.n987 B.n986 585
R654 B.n984 B.n101 585
R655 B.n101 B.n100 585
R656 B.n1095 B.n1094 585
R657 B.n1093 B.n2 585
R658 B.n982 B.n101 521.33
R659 B.n979 B.n156 521.33
R660 B.n531 B.n469 521.33
R661 B.n739 B.n471 521.33
R662 B.n157 B.t15 396.079
R663 B.n528 B.t13 396.079
R664 B.n159 B.t8 396.079
R665 B.n526 B.t19 396.079
R666 B.n158 B.t16 317.728
R667 B.n529 B.t12 317.728
R668 B.n160 B.t9 317.728
R669 B.n527 B.t18 317.728
R670 B.n159 B.t6 300.671
R671 B.n157 B.t14 300.671
R672 B.n528 B.t10 300.671
R673 B.n526 B.t17 300.671
R674 B.n980 B.n154 256.663
R675 B.n980 B.n153 256.663
R676 B.n980 B.n152 256.663
R677 B.n980 B.n151 256.663
R678 B.n980 B.n150 256.663
R679 B.n980 B.n149 256.663
R680 B.n980 B.n148 256.663
R681 B.n980 B.n147 256.663
R682 B.n980 B.n146 256.663
R683 B.n980 B.n145 256.663
R684 B.n980 B.n144 256.663
R685 B.n980 B.n143 256.663
R686 B.n980 B.n142 256.663
R687 B.n980 B.n141 256.663
R688 B.n980 B.n140 256.663
R689 B.n980 B.n139 256.663
R690 B.n980 B.n138 256.663
R691 B.n980 B.n137 256.663
R692 B.n980 B.n136 256.663
R693 B.n980 B.n135 256.663
R694 B.n980 B.n134 256.663
R695 B.n980 B.n133 256.663
R696 B.n980 B.n132 256.663
R697 B.n980 B.n131 256.663
R698 B.n980 B.n130 256.663
R699 B.n980 B.n129 256.663
R700 B.n980 B.n128 256.663
R701 B.n980 B.n127 256.663
R702 B.n980 B.n126 256.663
R703 B.n980 B.n125 256.663
R704 B.n980 B.n124 256.663
R705 B.n980 B.n123 256.663
R706 B.n980 B.n122 256.663
R707 B.n980 B.n121 256.663
R708 B.n980 B.n120 256.663
R709 B.n980 B.n119 256.663
R710 B.n980 B.n118 256.663
R711 B.n980 B.n117 256.663
R712 B.n980 B.n116 256.663
R713 B.n980 B.n115 256.663
R714 B.n980 B.n114 256.663
R715 B.n980 B.n113 256.663
R716 B.n980 B.n112 256.663
R717 B.n980 B.n111 256.663
R718 B.n980 B.n110 256.663
R719 B.n980 B.n109 256.663
R720 B.n980 B.n108 256.663
R721 B.n980 B.n107 256.663
R722 B.n980 B.n106 256.663
R723 B.n980 B.n105 256.663
R724 B.n980 B.n104 256.663
R725 B.n981 B.n980 256.663
R726 B.n738 B.n737 256.663
R727 B.n737 B.n474 256.663
R728 B.n737 B.n475 256.663
R729 B.n737 B.n476 256.663
R730 B.n737 B.n477 256.663
R731 B.n737 B.n478 256.663
R732 B.n737 B.n479 256.663
R733 B.n737 B.n480 256.663
R734 B.n737 B.n481 256.663
R735 B.n737 B.n482 256.663
R736 B.n737 B.n483 256.663
R737 B.n737 B.n484 256.663
R738 B.n737 B.n485 256.663
R739 B.n737 B.n486 256.663
R740 B.n737 B.n487 256.663
R741 B.n737 B.n488 256.663
R742 B.n737 B.n489 256.663
R743 B.n737 B.n490 256.663
R744 B.n737 B.n491 256.663
R745 B.n737 B.n492 256.663
R746 B.n737 B.n493 256.663
R747 B.n737 B.n494 256.663
R748 B.n737 B.n495 256.663
R749 B.n737 B.n496 256.663
R750 B.n737 B.n497 256.663
R751 B.n737 B.n498 256.663
R752 B.n737 B.n499 256.663
R753 B.n737 B.n500 256.663
R754 B.n737 B.n501 256.663
R755 B.n737 B.n502 256.663
R756 B.n737 B.n503 256.663
R757 B.n737 B.n504 256.663
R758 B.n737 B.n505 256.663
R759 B.n737 B.n506 256.663
R760 B.n737 B.n507 256.663
R761 B.n737 B.n508 256.663
R762 B.n737 B.n509 256.663
R763 B.n737 B.n510 256.663
R764 B.n737 B.n511 256.663
R765 B.n737 B.n512 256.663
R766 B.n737 B.n513 256.663
R767 B.n737 B.n514 256.663
R768 B.n737 B.n515 256.663
R769 B.n737 B.n516 256.663
R770 B.n737 B.n517 256.663
R771 B.n737 B.n518 256.663
R772 B.n737 B.n519 256.663
R773 B.n737 B.n520 256.663
R774 B.n737 B.n521 256.663
R775 B.n737 B.n522 256.663
R776 B.n737 B.n523 256.663
R777 B.n737 B.n524 256.663
R778 B.n1097 B.n1096 256.663
R779 B.n162 B.n103 163.367
R780 B.n166 B.n165 163.367
R781 B.n170 B.n169 163.367
R782 B.n174 B.n173 163.367
R783 B.n178 B.n177 163.367
R784 B.n182 B.n181 163.367
R785 B.n186 B.n185 163.367
R786 B.n190 B.n189 163.367
R787 B.n194 B.n193 163.367
R788 B.n198 B.n197 163.367
R789 B.n202 B.n201 163.367
R790 B.n206 B.n205 163.367
R791 B.n210 B.n209 163.367
R792 B.n214 B.n213 163.367
R793 B.n218 B.n217 163.367
R794 B.n222 B.n221 163.367
R795 B.n226 B.n225 163.367
R796 B.n230 B.n229 163.367
R797 B.n234 B.n233 163.367
R798 B.n238 B.n237 163.367
R799 B.n242 B.n241 163.367
R800 B.n246 B.n245 163.367
R801 B.n250 B.n249 163.367
R802 B.n254 B.n253 163.367
R803 B.n258 B.n257 163.367
R804 B.n262 B.n261 163.367
R805 B.n266 B.n265 163.367
R806 B.n270 B.n269 163.367
R807 B.n275 B.n274 163.367
R808 B.n279 B.n278 163.367
R809 B.n283 B.n282 163.367
R810 B.n287 B.n286 163.367
R811 B.n291 B.n290 163.367
R812 B.n295 B.n294 163.367
R813 B.n299 B.n298 163.367
R814 B.n303 B.n302 163.367
R815 B.n307 B.n306 163.367
R816 B.n311 B.n310 163.367
R817 B.n315 B.n314 163.367
R818 B.n319 B.n318 163.367
R819 B.n323 B.n322 163.367
R820 B.n327 B.n326 163.367
R821 B.n331 B.n330 163.367
R822 B.n335 B.n334 163.367
R823 B.n339 B.n338 163.367
R824 B.n343 B.n342 163.367
R825 B.n347 B.n346 163.367
R826 B.n351 B.n350 163.367
R827 B.n355 B.n354 163.367
R828 B.n359 B.n358 163.367
R829 B.n363 B.n362 163.367
R830 B.n979 B.n155 163.367
R831 B.n745 B.n469 163.367
R832 B.n745 B.n467 163.367
R833 B.n749 B.n467 163.367
R834 B.n749 B.n461 163.367
R835 B.n757 B.n461 163.367
R836 B.n757 B.n459 163.367
R837 B.n761 B.n459 163.367
R838 B.n761 B.n453 163.367
R839 B.n769 B.n453 163.367
R840 B.n769 B.n451 163.367
R841 B.n773 B.n451 163.367
R842 B.n773 B.n445 163.367
R843 B.n781 B.n445 163.367
R844 B.n781 B.n443 163.367
R845 B.n785 B.n443 163.367
R846 B.n785 B.n437 163.367
R847 B.n793 B.n437 163.367
R848 B.n793 B.n435 163.367
R849 B.n797 B.n435 163.367
R850 B.n797 B.n429 163.367
R851 B.n805 B.n429 163.367
R852 B.n805 B.n427 163.367
R853 B.n809 B.n427 163.367
R854 B.n809 B.n422 163.367
R855 B.n818 B.n422 163.367
R856 B.n818 B.n420 163.367
R857 B.n822 B.n420 163.367
R858 B.n822 B.n414 163.367
R859 B.n830 B.n414 163.367
R860 B.n830 B.n412 163.367
R861 B.n834 B.n412 163.367
R862 B.n834 B.n406 163.367
R863 B.n842 B.n406 163.367
R864 B.n842 B.n404 163.367
R865 B.n846 B.n404 163.367
R866 B.n846 B.n399 163.367
R867 B.n855 B.n399 163.367
R868 B.n855 B.n397 163.367
R869 B.n859 B.n397 163.367
R870 B.n859 B.n391 163.367
R871 B.n867 B.n391 163.367
R872 B.n867 B.n389 163.367
R873 B.n871 B.n389 163.367
R874 B.n871 B.n383 163.367
R875 B.n879 B.n383 163.367
R876 B.n879 B.n381 163.367
R877 B.n883 B.n381 163.367
R878 B.n883 B.n375 163.367
R879 B.n891 B.n375 163.367
R880 B.n891 B.n373 163.367
R881 B.n896 B.n373 163.367
R882 B.n896 B.n367 163.367
R883 B.n904 B.n367 163.367
R884 B.n905 B.n904 163.367
R885 B.n905 B.n5 163.367
R886 B.n6 B.n5 163.367
R887 B.n7 B.n6 163.367
R888 B.n911 B.n7 163.367
R889 B.n912 B.n911 163.367
R890 B.n912 B.n13 163.367
R891 B.n14 B.n13 163.367
R892 B.n15 B.n14 163.367
R893 B.n917 B.n15 163.367
R894 B.n917 B.n20 163.367
R895 B.n21 B.n20 163.367
R896 B.n22 B.n21 163.367
R897 B.n922 B.n22 163.367
R898 B.n922 B.n27 163.367
R899 B.n28 B.n27 163.367
R900 B.n29 B.n28 163.367
R901 B.n927 B.n29 163.367
R902 B.n927 B.n34 163.367
R903 B.n35 B.n34 163.367
R904 B.n36 B.n35 163.367
R905 B.n932 B.n36 163.367
R906 B.n932 B.n41 163.367
R907 B.n42 B.n41 163.367
R908 B.n43 B.n42 163.367
R909 B.n937 B.n43 163.367
R910 B.n937 B.n48 163.367
R911 B.n49 B.n48 163.367
R912 B.n50 B.n49 163.367
R913 B.n942 B.n50 163.367
R914 B.n942 B.n55 163.367
R915 B.n56 B.n55 163.367
R916 B.n57 B.n56 163.367
R917 B.n947 B.n57 163.367
R918 B.n947 B.n62 163.367
R919 B.n63 B.n62 163.367
R920 B.n64 B.n63 163.367
R921 B.n952 B.n64 163.367
R922 B.n952 B.n69 163.367
R923 B.n70 B.n69 163.367
R924 B.n71 B.n70 163.367
R925 B.n957 B.n71 163.367
R926 B.n957 B.n76 163.367
R927 B.n77 B.n76 163.367
R928 B.n78 B.n77 163.367
R929 B.n962 B.n78 163.367
R930 B.n962 B.n83 163.367
R931 B.n84 B.n83 163.367
R932 B.n85 B.n84 163.367
R933 B.n967 B.n85 163.367
R934 B.n967 B.n90 163.367
R935 B.n91 B.n90 163.367
R936 B.n92 B.n91 163.367
R937 B.n972 B.n92 163.367
R938 B.n972 B.n97 163.367
R939 B.n98 B.n97 163.367
R940 B.n99 B.n98 163.367
R941 B.n156 B.n99 163.367
R942 B.n736 B.n473 163.367
R943 B.n736 B.n525 163.367
R944 B.n732 B.n731 163.367
R945 B.n728 B.n727 163.367
R946 B.n724 B.n723 163.367
R947 B.n720 B.n719 163.367
R948 B.n716 B.n715 163.367
R949 B.n712 B.n711 163.367
R950 B.n708 B.n707 163.367
R951 B.n704 B.n703 163.367
R952 B.n700 B.n699 163.367
R953 B.n696 B.n695 163.367
R954 B.n692 B.n691 163.367
R955 B.n688 B.n687 163.367
R956 B.n684 B.n683 163.367
R957 B.n680 B.n679 163.367
R958 B.n676 B.n675 163.367
R959 B.n672 B.n671 163.367
R960 B.n668 B.n667 163.367
R961 B.n664 B.n663 163.367
R962 B.n660 B.n659 163.367
R963 B.n656 B.n655 163.367
R964 B.n652 B.n651 163.367
R965 B.n648 B.n647 163.367
R966 B.n643 B.n642 163.367
R967 B.n639 B.n638 163.367
R968 B.n635 B.n634 163.367
R969 B.n631 B.n630 163.367
R970 B.n627 B.n626 163.367
R971 B.n623 B.n622 163.367
R972 B.n619 B.n618 163.367
R973 B.n615 B.n614 163.367
R974 B.n611 B.n610 163.367
R975 B.n607 B.n606 163.367
R976 B.n603 B.n602 163.367
R977 B.n599 B.n598 163.367
R978 B.n595 B.n594 163.367
R979 B.n591 B.n590 163.367
R980 B.n587 B.n586 163.367
R981 B.n583 B.n582 163.367
R982 B.n579 B.n578 163.367
R983 B.n575 B.n574 163.367
R984 B.n571 B.n570 163.367
R985 B.n567 B.n566 163.367
R986 B.n563 B.n562 163.367
R987 B.n559 B.n558 163.367
R988 B.n555 B.n554 163.367
R989 B.n551 B.n550 163.367
R990 B.n547 B.n546 163.367
R991 B.n543 B.n542 163.367
R992 B.n539 B.n538 163.367
R993 B.n535 B.n534 163.367
R994 B.n743 B.n471 163.367
R995 B.n743 B.n465 163.367
R996 B.n751 B.n465 163.367
R997 B.n751 B.n463 163.367
R998 B.n755 B.n463 163.367
R999 B.n755 B.n457 163.367
R1000 B.n763 B.n457 163.367
R1001 B.n763 B.n455 163.367
R1002 B.n767 B.n455 163.367
R1003 B.n767 B.n449 163.367
R1004 B.n775 B.n449 163.367
R1005 B.n775 B.n447 163.367
R1006 B.n779 B.n447 163.367
R1007 B.n779 B.n441 163.367
R1008 B.n787 B.n441 163.367
R1009 B.n787 B.n439 163.367
R1010 B.n791 B.n439 163.367
R1011 B.n791 B.n433 163.367
R1012 B.n799 B.n433 163.367
R1013 B.n799 B.n431 163.367
R1014 B.n803 B.n431 163.367
R1015 B.n803 B.n425 163.367
R1016 B.n812 B.n425 163.367
R1017 B.n812 B.n423 163.367
R1018 B.n816 B.n423 163.367
R1019 B.n816 B.n418 163.367
R1020 B.n824 B.n418 163.367
R1021 B.n824 B.n416 163.367
R1022 B.n828 B.n416 163.367
R1023 B.n828 B.n410 163.367
R1024 B.n836 B.n410 163.367
R1025 B.n836 B.n408 163.367
R1026 B.n840 B.n408 163.367
R1027 B.n840 B.n402 163.367
R1028 B.n849 B.n402 163.367
R1029 B.n849 B.n400 163.367
R1030 B.n853 B.n400 163.367
R1031 B.n853 B.n395 163.367
R1032 B.n861 B.n395 163.367
R1033 B.n861 B.n393 163.367
R1034 B.n865 B.n393 163.367
R1035 B.n865 B.n387 163.367
R1036 B.n873 B.n387 163.367
R1037 B.n873 B.n385 163.367
R1038 B.n877 B.n385 163.367
R1039 B.n877 B.n379 163.367
R1040 B.n885 B.n379 163.367
R1041 B.n885 B.n377 163.367
R1042 B.n889 B.n377 163.367
R1043 B.n889 B.n371 163.367
R1044 B.n898 B.n371 163.367
R1045 B.n898 B.n369 163.367
R1046 B.n902 B.n369 163.367
R1047 B.n902 B.n3 163.367
R1048 B.n1095 B.n3 163.367
R1049 B.n1091 B.n2 163.367
R1050 B.n1091 B.n1090 163.367
R1051 B.n1090 B.n9 163.367
R1052 B.n1086 B.n9 163.367
R1053 B.n1086 B.n11 163.367
R1054 B.n1082 B.n11 163.367
R1055 B.n1082 B.n17 163.367
R1056 B.n1078 B.n17 163.367
R1057 B.n1078 B.n19 163.367
R1058 B.n1074 B.n19 163.367
R1059 B.n1074 B.n24 163.367
R1060 B.n1070 B.n24 163.367
R1061 B.n1070 B.n26 163.367
R1062 B.n1066 B.n26 163.367
R1063 B.n1066 B.n31 163.367
R1064 B.n1062 B.n31 163.367
R1065 B.n1062 B.n33 163.367
R1066 B.n1058 B.n33 163.367
R1067 B.n1058 B.n37 163.367
R1068 B.n1054 B.n37 163.367
R1069 B.n1054 B.n39 163.367
R1070 B.n1050 B.n39 163.367
R1071 B.n1050 B.n45 163.367
R1072 B.n1046 B.n45 163.367
R1073 B.n1046 B.n47 163.367
R1074 B.n1042 B.n47 163.367
R1075 B.n1042 B.n52 163.367
R1076 B.n1038 B.n52 163.367
R1077 B.n1038 B.n54 163.367
R1078 B.n1034 B.n54 163.367
R1079 B.n1034 B.n58 163.367
R1080 B.n1030 B.n58 163.367
R1081 B.n1030 B.n60 163.367
R1082 B.n1026 B.n60 163.367
R1083 B.n1026 B.n66 163.367
R1084 B.n1022 B.n66 163.367
R1085 B.n1022 B.n68 163.367
R1086 B.n1018 B.n68 163.367
R1087 B.n1018 B.n73 163.367
R1088 B.n1014 B.n73 163.367
R1089 B.n1014 B.n75 163.367
R1090 B.n1010 B.n75 163.367
R1091 B.n1010 B.n80 163.367
R1092 B.n1006 B.n80 163.367
R1093 B.n1006 B.n82 163.367
R1094 B.n1002 B.n82 163.367
R1095 B.n1002 B.n87 163.367
R1096 B.n998 B.n87 163.367
R1097 B.n998 B.n89 163.367
R1098 B.n994 B.n89 163.367
R1099 B.n994 B.n94 163.367
R1100 B.n990 B.n94 163.367
R1101 B.n990 B.n96 163.367
R1102 B.n986 B.n96 163.367
R1103 B.n986 B.n101 163.367
R1104 B.n160 B.n159 78.352
R1105 B.n158 B.n157 78.352
R1106 B.n529 B.n528 78.352
R1107 B.n527 B.n526 78.352
R1108 B.n737 B.n470 75.6273
R1109 B.n980 B.n100 75.6273
R1110 B.n982 B.n981 71.676
R1111 B.n162 B.n104 71.676
R1112 B.n166 B.n105 71.676
R1113 B.n170 B.n106 71.676
R1114 B.n174 B.n107 71.676
R1115 B.n178 B.n108 71.676
R1116 B.n182 B.n109 71.676
R1117 B.n186 B.n110 71.676
R1118 B.n190 B.n111 71.676
R1119 B.n194 B.n112 71.676
R1120 B.n198 B.n113 71.676
R1121 B.n202 B.n114 71.676
R1122 B.n206 B.n115 71.676
R1123 B.n210 B.n116 71.676
R1124 B.n214 B.n117 71.676
R1125 B.n218 B.n118 71.676
R1126 B.n222 B.n119 71.676
R1127 B.n226 B.n120 71.676
R1128 B.n230 B.n121 71.676
R1129 B.n234 B.n122 71.676
R1130 B.n238 B.n123 71.676
R1131 B.n242 B.n124 71.676
R1132 B.n246 B.n125 71.676
R1133 B.n250 B.n126 71.676
R1134 B.n254 B.n127 71.676
R1135 B.n258 B.n128 71.676
R1136 B.n262 B.n129 71.676
R1137 B.n266 B.n130 71.676
R1138 B.n270 B.n131 71.676
R1139 B.n275 B.n132 71.676
R1140 B.n279 B.n133 71.676
R1141 B.n283 B.n134 71.676
R1142 B.n287 B.n135 71.676
R1143 B.n291 B.n136 71.676
R1144 B.n295 B.n137 71.676
R1145 B.n299 B.n138 71.676
R1146 B.n303 B.n139 71.676
R1147 B.n307 B.n140 71.676
R1148 B.n311 B.n141 71.676
R1149 B.n315 B.n142 71.676
R1150 B.n319 B.n143 71.676
R1151 B.n323 B.n144 71.676
R1152 B.n327 B.n145 71.676
R1153 B.n331 B.n146 71.676
R1154 B.n335 B.n147 71.676
R1155 B.n339 B.n148 71.676
R1156 B.n343 B.n149 71.676
R1157 B.n347 B.n150 71.676
R1158 B.n351 B.n151 71.676
R1159 B.n355 B.n152 71.676
R1160 B.n359 B.n153 71.676
R1161 B.n363 B.n154 71.676
R1162 B.n155 B.n154 71.676
R1163 B.n362 B.n153 71.676
R1164 B.n358 B.n152 71.676
R1165 B.n354 B.n151 71.676
R1166 B.n350 B.n150 71.676
R1167 B.n346 B.n149 71.676
R1168 B.n342 B.n148 71.676
R1169 B.n338 B.n147 71.676
R1170 B.n334 B.n146 71.676
R1171 B.n330 B.n145 71.676
R1172 B.n326 B.n144 71.676
R1173 B.n322 B.n143 71.676
R1174 B.n318 B.n142 71.676
R1175 B.n314 B.n141 71.676
R1176 B.n310 B.n140 71.676
R1177 B.n306 B.n139 71.676
R1178 B.n302 B.n138 71.676
R1179 B.n298 B.n137 71.676
R1180 B.n294 B.n136 71.676
R1181 B.n290 B.n135 71.676
R1182 B.n286 B.n134 71.676
R1183 B.n282 B.n133 71.676
R1184 B.n278 B.n132 71.676
R1185 B.n274 B.n131 71.676
R1186 B.n269 B.n130 71.676
R1187 B.n265 B.n129 71.676
R1188 B.n261 B.n128 71.676
R1189 B.n257 B.n127 71.676
R1190 B.n253 B.n126 71.676
R1191 B.n249 B.n125 71.676
R1192 B.n245 B.n124 71.676
R1193 B.n241 B.n123 71.676
R1194 B.n237 B.n122 71.676
R1195 B.n233 B.n121 71.676
R1196 B.n229 B.n120 71.676
R1197 B.n225 B.n119 71.676
R1198 B.n221 B.n118 71.676
R1199 B.n217 B.n117 71.676
R1200 B.n213 B.n116 71.676
R1201 B.n209 B.n115 71.676
R1202 B.n205 B.n114 71.676
R1203 B.n201 B.n113 71.676
R1204 B.n197 B.n112 71.676
R1205 B.n193 B.n111 71.676
R1206 B.n189 B.n110 71.676
R1207 B.n185 B.n109 71.676
R1208 B.n181 B.n108 71.676
R1209 B.n177 B.n107 71.676
R1210 B.n173 B.n106 71.676
R1211 B.n169 B.n105 71.676
R1212 B.n165 B.n104 71.676
R1213 B.n981 B.n103 71.676
R1214 B.n739 B.n738 71.676
R1215 B.n525 B.n474 71.676
R1216 B.n731 B.n475 71.676
R1217 B.n727 B.n476 71.676
R1218 B.n723 B.n477 71.676
R1219 B.n719 B.n478 71.676
R1220 B.n715 B.n479 71.676
R1221 B.n711 B.n480 71.676
R1222 B.n707 B.n481 71.676
R1223 B.n703 B.n482 71.676
R1224 B.n699 B.n483 71.676
R1225 B.n695 B.n484 71.676
R1226 B.n691 B.n485 71.676
R1227 B.n687 B.n486 71.676
R1228 B.n683 B.n487 71.676
R1229 B.n679 B.n488 71.676
R1230 B.n675 B.n489 71.676
R1231 B.n671 B.n490 71.676
R1232 B.n667 B.n491 71.676
R1233 B.n663 B.n492 71.676
R1234 B.n659 B.n493 71.676
R1235 B.n655 B.n494 71.676
R1236 B.n651 B.n495 71.676
R1237 B.n647 B.n496 71.676
R1238 B.n642 B.n497 71.676
R1239 B.n638 B.n498 71.676
R1240 B.n634 B.n499 71.676
R1241 B.n630 B.n500 71.676
R1242 B.n626 B.n501 71.676
R1243 B.n622 B.n502 71.676
R1244 B.n618 B.n503 71.676
R1245 B.n614 B.n504 71.676
R1246 B.n610 B.n505 71.676
R1247 B.n606 B.n506 71.676
R1248 B.n602 B.n507 71.676
R1249 B.n598 B.n508 71.676
R1250 B.n594 B.n509 71.676
R1251 B.n590 B.n510 71.676
R1252 B.n586 B.n511 71.676
R1253 B.n582 B.n512 71.676
R1254 B.n578 B.n513 71.676
R1255 B.n574 B.n514 71.676
R1256 B.n570 B.n515 71.676
R1257 B.n566 B.n516 71.676
R1258 B.n562 B.n517 71.676
R1259 B.n558 B.n518 71.676
R1260 B.n554 B.n519 71.676
R1261 B.n550 B.n520 71.676
R1262 B.n546 B.n521 71.676
R1263 B.n542 B.n522 71.676
R1264 B.n538 B.n523 71.676
R1265 B.n534 B.n524 71.676
R1266 B.n738 B.n473 71.676
R1267 B.n732 B.n474 71.676
R1268 B.n728 B.n475 71.676
R1269 B.n724 B.n476 71.676
R1270 B.n720 B.n477 71.676
R1271 B.n716 B.n478 71.676
R1272 B.n712 B.n479 71.676
R1273 B.n708 B.n480 71.676
R1274 B.n704 B.n481 71.676
R1275 B.n700 B.n482 71.676
R1276 B.n696 B.n483 71.676
R1277 B.n692 B.n484 71.676
R1278 B.n688 B.n485 71.676
R1279 B.n684 B.n486 71.676
R1280 B.n680 B.n487 71.676
R1281 B.n676 B.n488 71.676
R1282 B.n672 B.n489 71.676
R1283 B.n668 B.n490 71.676
R1284 B.n664 B.n491 71.676
R1285 B.n660 B.n492 71.676
R1286 B.n656 B.n493 71.676
R1287 B.n652 B.n494 71.676
R1288 B.n648 B.n495 71.676
R1289 B.n643 B.n496 71.676
R1290 B.n639 B.n497 71.676
R1291 B.n635 B.n498 71.676
R1292 B.n631 B.n499 71.676
R1293 B.n627 B.n500 71.676
R1294 B.n623 B.n501 71.676
R1295 B.n619 B.n502 71.676
R1296 B.n615 B.n503 71.676
R1297 B.n611 B.n504 71.676
R1298 B.n607 B.n505 71.676
R1299 B.n603 B.n506 71.676
R1300 B.n599 B.n507 71.676
R1301 B.n595 B.n508 71.676
R1302 B.n591 B.n509 71.676
R1303 B.n587 B.n510 71.676
R1304 B.n583 B.n511 71.676
R1305 B.n579 B.n512 71.676
R1306 B.n575 B.n513 71.676
R1307 B.n571 B.n514 71.676
R1308 B.n567 B.n515 71.676
R1309 B.n563 B.n516 71.676
R1310 B.n559 B.n517 71.676
R1311 B.n555 B.n518 71.676
R1312 B.n551 B.n519 71.676
R1313 B.n547 B.n520 71.676
R1314 B.n543 B.n521 71.676
R1315 B.n539 B.n522 71.676
R1316 B.n535 B.n523 71.676
R1317 B.n531 B.n524 71.676
R1318 B.n1096 B.n1095 71.676
R1319 B.n1096 B.n2 71.676
R1320 B.n161 B.n160 59.5399
R1321 B.n272 B.n158 59.5399
R1322 B.n530 B.n529 59.5399
R1323 B.n645 B.n527 59.5399
R1324 B.n744 B.n470 38.6668
R1325 B.n744 B.n466 38.6668
R1326 B.n750 B.n466 38.6668
R1327 B.n750 B.n462 38.6668
R1328 B.n756 B.n462 38.6668
R1329 B.n756 B.n458 38.6668
R1330 B.n762 B.n458 38.6668
R1331 B.n762 B.n454 38.6668
R1332 B.n768 B.n454 38.6668
R1333 B.n774 B.n450 38.6668
R1334 B.n774 B.n446 38.6668
R1335 B.n780 B.n446 38.6668
R1336 B.n780 B.n442 38.6668
R1337 B.n786 B.n442 38.6668
R1338 B.n786 B.n438 38.6668
R1339 B.n792 B.n438 38.6668
R1340 B.n792 B.n434 38.6668
R1341 B.n798 B.n434 38.6668
R1342 B.n798 B.n430 38.6668
R1343 B.n804 B.n430 38.6668
R1344 B.n804 B.n426 38.6668
R1345 B.n811 B.n426 38.6668
R1346 B.n811 B.n810 38.6668
R1347 B.n817 B.n419 38.6668
R1348 B.n823 B.n419 38.6668
R1349 B.n823 B.n415 38.6668
R1350 B.n829 B.n415 38.6668
R1351 B.n829 B.n411 38.6668
R1352 B.n835 B.n411 38.6668
R1353 B.n835 B.n407 38.6668
R1354 B.n841 B.n407 38.6668
R1355 B.n841 B.n403 38.6668
R1356 B.n848 B.n403 38.6668
R1357 B.n848 B.n847 38.6668
R1358 B.n854 B.n396 38.6668
R1359 B.n860 B.n396 38.6668
R1360 B.n860 B.n392 38.6668
R1361 B.n866 B.n392 38.6668
R1362 B.n866 B.n388 38.6668
R1363 B.n872 B.n388 38.6668
R1364 B.n872 B.n384 38.6668
R1365 B.n878 B.n384 38.6668
R1366 B.n878 B.n380 38.6668
R1367 B.n884 B.n380 38.6668
R1368 B.n890 B.n376 38.6668
R1369 B.n890 B.n372 38.6668
R1370 B.n897 B.n372 38.6668
R1371 B.n897 B.n368 38.6668
R1372 B.n903 B.n368 38.6668
R1373 B.n903 B.n4 38.6668
R1374 B.n1094 B.n4 38.6668
R1375 B.n1094 B.n1093 38.6668
R1376 B.n1093 B.n1092 38.6668
R1377 B.n1092 B.n8 38.6668
R1378 B.n12 B.n8 38.6668
R1379 B.n1085 B.n12 38.6668
R1380 B.n1085 B.n1084 38.6668
R1381 B.n1084 B.n1083 38.6668
R1382 B.n1083 B.n16 38.6668
R1383 B.n1077 B.n1076 38.6668
R1384 B.n1076 B.n1075 38.6668
R1385 B.n1075 B.n23 38.6668
R1386 B.n1069 B.n23 38.6668
R1387 B.n1069 B.n1068 38.6668
R1388 B.n1068 B.n1067 38.6668
R1389 B.n1067 B.n30 38.6668
R1390 B.n1061 B.n30 38.6668
R1391 B.n1061 B.n1060 38.6668
R1392 B.n1060 B.n1059 38.6668
R1393 B.n1053 B.n40 38.6668
R1394 B.n1053 B.n1052 38.6668
R1395 B.n1052 B.n1051 38.6668
R1396 B.n1051 B.n44 38.6668
R1397 B.n1045 B.n44 38.6668
R1398 B.n1045 B.n1044 38.6668
R1399 B.n1044 B.n1043 38.6668
R1400 B.n1043 B.n51 38.6668
R1401 B.n1037 B.n51 38.6668
R1402 B.n1037 B.n1036 38.6668
R1403 B.n1036 B.n1035 38.6668
R1404 B.n1029 B.n61 38.6668
R1405 B.n1029 B.n1028 38.6668
R1406 B.n1028 B.n1027 38.6668
R1407 B.n1027 B.n65 38.6668
R1408 B.n1021 B.n65 38.6668
R1409 B.n1021 B.n1020 38.6668
R1410 B.n1020 B.n1019 38.6668
R1411 B.n1019 B.n72 38.6668
R1412 B.n1013 B.n72 38.6668
R1413 B.n1013 B.n1012 38.6668
R1414 B.n1012 B.n1011 38.6668
R1415 B.n1011 B.n79 38.6668
R1416 B.n1005 B.n79 38.6668
R1417 B.n1005 B.n1004 38.6668
R1418 B.n1003 B.n86 38.6668
R1419 B.n997 B.n86 38.6668
R1420 B.n997 B.n996 38.6668
R1421 B.n996 B.n995 38.6668
R1422 B.n995 B.n93 38.6668
R1423 B.n989 B.n93 38.6668
R1424 B.n989 B.n988 38.6668
R1425 B.n988 B.n987 38.6668
R1426 B.n987 B.n100 38.6668
R1427 B.n884 B.t4 36.961
R1428 B.n1077 B.t2 36.961
R1429 B.n854 B.t3 35.8237
R1430 B.n1059 B.t5 35.8237
R1431 B.t11 B.n450 34.6865
R1432 B.n1004 B.t7 34.6865
R1433 B.n741 B.n740 33.8737
R1434 B.n532 B.n468 33.8737
R1435 B.n978 B.n977 33.8737
R1436 B.n984 B.n983 33.8737
R1437 B.n817 B.t1 31.2747
R1438 B.n1035 B.t0 31.2747
R1439 B B.n1097 18.0485
R1440 B.n742 B.n741 10.6151
R1441 B.n742 B.n464 10.6151
R1442 B.n752 B.n464 10.6151
R1443 B.n753 B.n752 10.6151
R1444 B.n754 B.n753 10.6151
R1445 B.n754 B.n456 10.6151
R1446 B.n764 B.n456 10.6151
R1447 B.n765 B.n764 10.6151
R1448 B.n766 B.n765 10.6151
R1449 B.n766 B.n448 10.6151
R1450 B.n776 B.n448 10.6151
R1451 B.n777 B.n776 10.6151
R1452 B.n778 B.n777 10.6151
R1453 B.n778 B.n440 10.6151
R1454 B.n788 B.n440 10.6151
R1455 B.n789 B.n788 10.6151
R1456 B.n790 B.n789 10.6151
R1457 B.n790 B.n432 10.6151
R1458 B.n800 B.n432 10.6151
R1459 B.n801 B.n800 10.6151
R1460 B.n802 B.n801 10.6151
R1461 B.n802 B.n424 10.6151
R1462 B.n813 B.n424 10.6151
R1463 B.n814 B.n813 10.6151
R1464 B.n815 B.n814 10.6151
R1465 B.n815 B.n417 10.6151
R1466 B.n825 B.n417 10.6151
R1467 B.n826 B.n825 10.6151
R1468 B.n827 B.n826 10.6151
R1469 B.n827 B.n409 10.6151
R1470 B.n837 B.n409 10.6151
R1471 B.n838 B.n837 10.6151
R1472 B.n839 B.n838 10.6151
R1473 B.n839 B.n401 10.6151
R1474 B.n850 B.n401 10.6151
R1475 B.n851 B.n850 10.6151
R1476 B.n852 B.n851 10.6151
R1477 B.n852 B.n394 10.6151
R1478 B.n862 B.n394 10.6151
R1479 B.n863 B.n862 10.6151
R1480 B.n864 B.n863 10.6151
R1481 B.n864 B.n386 10.6151
R1482 B.n874 B.n386 10.6151
R1483 B.n875 B.n874 10.6151
R1484 B.n876 B.n875 10.6151
R1485 B.n876 B.n378 10.6151
R1486 B.n886 B.n378 10.6151
R1487 B.n887 B.n886 10.6151
R1488 B.n888 B.n887 10.6151
R1489 B.n888 B.n370 10.6151
R1490 B.n899 B.n370 10.6151
R1491 B.n900 B.n899 10.6151
R1492 B.n901 B.n900 10.6151
R1493 B.n901 B.n0 10.6151
R1494 B.n740 B.n472 10.6151
R1495 B.n735 B.n472 10.6151
R1496 B.n735 B.n734 10.6151
R1497 B.n734 B.n733 10.6151
R1498 B.n733 B.n730 10.6151
R1499 B.n730 B.n729 10.6151
R1500 B.n729 B.n726 10.6151
R1501 B.n726 B.n725 10.6151
R1502 B.n725 B.n722 10.6151
R1503 B.n722 B.n721 10.6151
R1504 B.n721 B.n718 10.6151
R1505 B.n718 B.n717 10.6151
R1506 B.n717 B.n714 10.6151
R1507 B.n714 B.n713 10.6151
R1508 B.n713 B.n710 10.6151
R1509 B.n710 B.n709 10.6151
R1510 B.n709 B.n706 10.6151
R1511 B.n706 B.n705 10.6151
R1512 B.n705 B.n702 10.6151
R1513 B.n702 B.n701 10.6151
R1514 B.n701 B.n698 10.6151
R1515 B.n698 B.n697 10.6151
R1516 B.n697 B.n694 10.6151
R1517 B.n694 B.n693 10.6151
R1518 B.n693 B.n690 10.6151
R1519 B.n690 B.n689 10.6151
R1520 B.n689 B.n686 10.6151
R1521 B.n686 B.n685 10.6151
R1522 B.n685 B.n682 10.6151
R1523 B.n682 B.n681 10.6151
R1524 B.n681 B.n678 10.6151
R1525 B.n678 B.n677 10.6151
R1526 B.n677 B.n674 10.6151
R1527 B.n674 B.n673 10.6151
R1528 B.n673 B.n670 10.6151
R1529 B.n670 B.n669 10.6151
R1530 B.n669 B.n666 10.6151
R1531 B.n666 B.n665 10.6151
R1532 B.n665 B.n662 10.6151
R1533 B.n662 B.n661 10.6151
R1534 B.n661 B.n658 10.6151
R1535 B.n658 B.n657 10.6151
R1536 B.n657 B.n654 10.6151
R1537 B.n654 B.n653 10.6151
R1538 B.n653 B.n650 10.6151
R1539 B.n650 B.n649 10.6151
R1540 B.n649 B.n646 10.6151
R1541 B.n644 B.n641 10.6151
R1542 B.n641 B.n640 10.6151
R1543 B.n640 B.n637 10.6151
R1544 B.n637 B.n636 10.6151
R1545 B.n636 B.n633 10.6151
R1546 B.n633 B.n632 10.6151
R1547 B.n632 B.n629 10.6151
R1548 B.n629 B.n628 10.6151
R1549 B.n625 B.n624 10.6151
R1550 B.n624 B.n621 10.6151
R1551 B.n621 B.n620 10.6151
R1552 B.n620 B.n617 10.6151
R1553 B.n617 B.n616 10.6151
R1554 B.n616 B.n613 10.6151
R1555 B.n613 B.n612 10.6151
R1556 B.n612 B.n609 10.6151
R1557 B.n609 B.n608 10.6151
R1558 B.n608 B.n605 10.6151
R1559 B.n605 B.n604 10.6151
R1560 B.n604 B.n601 10.6151
R1561 B.n601 B.n600 10.6151
R1562 B.n600 B.n597 10.6151
R1563 B.n597 B.n596 10.6151
R1564 B.n596 B.n593 10.6151
R1565 B.n593 B.n592 10.6151
R1566 B.n592 B.n589 10.6151
R1567 B.n589 B.n588 10.6151
R1568 B.n588 B.n585 10.6151
R1569 B.n585 B.n584 10.6151
R1570 B.n584 B.n581 10.6151
R1571 B.n581 B.n580 10.6151
R1572 B.n580 B.n577 10.6151
R1573 B.n577 B.n576 10.6151
R1574 B.n576 B.n573 10.6151
R1575 B.n573 B.n572 10.6151
R1576 B.n572 B.n569 10.6151
R1577 B.n569 B.n568 10.6151
R1578 B.n568 B.n565 10.6151
R1579 B.n565 B.n564 10.6151
R1580 B.n564 B.n561 10.6151
R1581 B.n561 B.n560 10.6151
R1582 B.n560 B.n557 10.6151
R1583 B.n557 B.n556 10.6151
R1584 B.n556 B.n553 10.6151
R1585 B.n553 B.n552 10.6151
R1586 B.n552 B.n549 10.6151
R1587 B.n549 B.n548 10.6151
R1588 B.n548 B.n545 10.6151
R1589 B.n545 B.n544 10.6151
R1590 B.n544 B.n541 10.6151
R1591 B.n541 B.n540 10.6151
R1592 B.n540 B.n537 10.6151
R1593 B.n537 B.n536 10.6151
R1594 B.n536 B.n533 10.6151
R1595 B.n533 B.n532 10.6151
R1596 B.n746 B.n468 10.6151
R1597 B.n747 B.n746 10.6151
R1598 B.n748 B.n747 10.6151
R1599 B.n748 B.n460 10.6151
R1600 B.n758 B.n460 10.6151
R1601 B.n759 B.n758 10.6151
R1602 B.n760 B.n759 10.6151
R1603 B.n760 B.n452 10.6151
R1604 B.n770 B.n452 10.6151
R1605 B.n771 B.n770 10.6151
R1606 B.n772 B.n771 10.6151
R1607 B.n772 B.n444 10.6151
R1608 B.n782 B.n444 10.6151
R1609 B.n783 B.n782 10.6151
R1610 B.n784 B.n783 10.6151
R1611 B.n784 B.n436 10.6151
R1612 B.n794 B.n436 10.6151
R1613 B.n795 B.n794 10.6151
R1614 B.n796 B.n795 10.6151
R1615 B.n796 B.n428 10.6151
R1616 B.n806 B.n428 10.6151
R1617 B.n807 B.n806 10.6151
R1618 B.n808 B.n807 10.6151
R1619 B.n808 B.n421 10.6151
R1620 B.n819 B.n421 10.6151
R1621 B.n820 B.n819 10.6151
R1622 B.n821 B.n820 10.6151
R1623 B.n821 B.n413 10.6151
R1624 B.n831 B.n413 10.6151
R1625 B.n832 B.n831 10.6151
R1626 B.n833 B.n832 10.6151
R1627 B.n833 B.n405 10.6151
R1628 B.n843 B.n405 10.6151
R1629 B.n844 B.n843 10.6151
R1630 B.n845 B.n844 10.6151
R1631 B.n845 B.n398 10.6151
R1632 B.n856 B.n398 10.6151
R1633 B.n857 B.n856 10.6151
R1634 B.n858 B.n857 10.6151
R1635 B.n858 B.n390 10.6151
R1636 B.n868 B.n390 10.6151
R1637 B.n869 B.n868 10.6151
R1638 B.n870 B.n869 10.6151
R1639 B.n870 B.n382 10.6151
R1640 B.n880 B.n382 10.6151
R1641 B.n881 B.n880 10.6151
R1642 B.n882 B.n881 10.6151
R1643 B.n882 B.n374 10.6151
R1644 B.n892 B.n374 10.6151
R1645 B.n893 B.n892 10.6151
R1646 B.n895 B.n893 10.6151
R1647 B.n895 B.n894 10.6151
R1648 B.n894 B.n366 10.6151
R1649 B.n906 B.n366 10.6151
R1650 B.n907 B.n906 10.6151
R1651 B.n908 B.n907 10.6151
R1652 B.n909 B.n908 10.6151
R1653 B.n910 B.n909 10.6151
R1654 B.n913 B.n910 10.6151
R1655 B.n914 B.n913 10.6151
R1656 B.n915 B.n914 10.6151
R1657 B.n916 B.n915 10.6151
R1658 B.n918 B.n916 10.6151
R1659 B.n919 B.n918 10.6151
R1660 B.n920 B.n919 10.6151
R1661 B.n921 B.n920 10.6151
R1662 B.n923 B.n921 10.6151
R1663 B.n924 B.n923 10.6151
R1664 B.n925 B.n924 10.6151
R1665 B.n926 B.n925 10.6151
R1666 B.n928 B.n926 10.6151
R1667 B.n929 B.n928 10.6151
R1668 B.n930 B.n929 10.6151
R1669 B.n931 B.n930 10.6151
R1670 B.n933 B.n931 10.6151
R1671 B.n934 B.n933 10.6151
R1672 B.n935 B.n934 10.6151
R1673 B.n936 B.n935 10.6151
R1674 B.n938 B.n936 10.6151
R1675 B.n939 B.n938 10.6151
R1676 B.n940 B.n939 10.6151
R1677 B.n941 B.n940 10.6151
R1678 B.n943 B.n941 10.6151
R1679 B.n944 B.n943 10.6151
R1680 B.n945 B.n944 10.6151
R1681 B.n946 B.n945 10.6151
R1682 B.n948 B.n946 10.6151
R1683 B.n949 B.n948 10.6151
R1684 B.n950 B.n949 10.6151
R1685 B.n951 B.n950 10.6151
R1686 B.n953 B.n951 10.6151
R1687 B.n954 B.n953 10.6151
R1688 B.n955 B.n954 10.6151
R1689 B.n956 B.n955 10.6151
R1690 B.n958 B.n956 10.6151
R1691 B.n959 B.n958 10.6151
R1692 B.n960 B.n959 10.6151
R1693 B.n961 B.n960 10.6151
R1694 B.n963 B.n961 10.6151
R1695 B.n964 B.n963 10.6151
R1696 B.n965 B.n964 10.6151
R1697 B.n966 B.n965 10.6151
R1698 B.n968 B.n966 10.6151
R1699 B.n969 B.n968 10.6151
R1700 B.n970 B.n969 10.6151
R1701 B.n971 B.n970 10.6151
R1702 B.n973 B.n971 10.6151
R1703 B.n974 B.n973 10.6151
R1704 B.n975 B.n974 10.6151
R1705 B.n976 B.n975 10.6151
R1706 B.n977 B.n976 10.6151
R1707 B.n1089 B.n1 10.6151
R1708 B.n1089 B.n1088 10.6151
R1709 B.n1088 B.n1087 10.6151
R1710 B.n1087 B.n10 10.6151
R1711 B.n1081 B.n10 10.6151
R1712 B.n1081 B.n1080 10.6151
R1713 B.n1080 B.n1079 10.6151
R1714 B.n1079 B.n18 10.6151
R1715 B.n1073 B.n18 10.6151
R1716 B.n1073 B.n1072 10.6151
R1717 B.n1072 B.n1071 10.6151
R1718 B.n1071 B.n25 10.6151
R1719 B.n1065 B.n25 10.6151
R1720 B.n1065 B.n1064 10.6151
R1721 B.n1064 B.n1063 10.6151
R1722 B.n1063 B.n32 10.6151
R1723 B.n1057 B.n32 10.6151
R1724 B.n1057 B.n1056 10.6151
R1725 B.n1056 B.n1055 10.6151
R1726 B.n1055 B.n38 10.6151
R1727 B.n1049 B.n38 10.6151
R1728 B.n1049 B.n1048 10.6151
R1729 B.n1048 B.n1047 10.6151
R1730 B.n1047 B.n46 10.6151
R1731 B.n1041 B.n46 10.6151
R1732 B.n1041 B.n1040 10.6151
R1733 B.n1040 B.n1039 10.6151
R1734 B.n1039 B.n53 10.6151
R1735 B.n1033 B.n53 10.6151
R1736 B.n1033 B.n1032 10.6151
R1737 B.n1032 B.n1031 10.6151
R1738 B.n1031 B.n59 10.6151
R1739 B.n1025 B.n59 10.6151
R1740 B.n1025 B.n1024 10.6151
R1741 B.n1024 B.n1023 10.6151
R1742 B.n1023 B.n67 10.6151
R1743 B.n1017 B.n67 10.6151
R1744 B.n1017 B.n1016 10.6151
R1745 B.n1016 B.n1015 10.6151
R1746 B.n1015 B.n74 10.6151
R1747 B.n1009 B.n74 10.6151
R1748 B.n1009 B.n1008 10.6151
R1749 B.n1008 B.n1007 10.6151
R1750 B.n1007 B.n81 10.6151
R1751 B.n1001 B.n81 10.6151
R1752 B.n1001 B.n1000 10.6151
R1753 B.n1000 B.n999 10.6151
R1754 B.n999 B.n88 10.6151
R1755 B.n993 B.n88 10.6151
R1756 B.n993 B.n992 10.6151
R1757 B.n992 B.n991 10.6151
R1758 B.n991 B.n95 10.6151
R1759 B.n985 B.n95 10.6151
R1760 B.n985 B.n984 10.6151
R1761 B.n983 B.n102 10.6151
R1762 B.n163 B.n102 10.6151
R1763 B.n164 B.n163 10.6151
R1764 B.n167 B.n164 10.6151
R1765 B.n168 B.n167 10.6151
R1766 B.n171 B.n168 10.6151
R1767 B.n172 B.n171 10.6151
R1768 B.n175 B.n172 10.6151
R1769 B.n176 B.n175 10.6151
R1770 B.n179 B.n176 10.6151
R1771 B.n180 B.n179 10.6151
R1772 B.n183 B.n180 10.6151
R1773 B.n184 B.n183 10.6151
R1774 B.n187 B.n184 10.6151
R1775 B.n188 B.n187 10.6151
R1776 B.n191 B.n188 10.6151
R1777 B.n192 B.n191 10.6151
R1778 B.n195 B.n192 10.6151
R1779 B.n196 B.n195 10.6151
R1780 B.n199 B.n196 10.6151
R1781 B.n200 B.n199 10.6151
R1782 B.n203 B.n200 10.6151
R1783 B.n204 B.n203 10.6151
R1784 B.n207 B.n204 10.6151
R1785 B.n208 B.n207 10.6151
R1786 B.n211 B.n208 10.6151
R1787 B.n212 B.n211 10.6151
R1788 B.n215 B.n212 10.6151
R1789 B.n216 B.n215 10.6151
R1790 B.n219 B.n216 10.6151
R1791 B.n220 B.n219 10.6151
R1792 B.n223 B.n220 10.6151
R1793 B.n224 B.n223 10.6151
R1794 B.n227 B.n224 10.6151
R1795 B.n228 B.n227 10.6151
R1796 B.n231 B.n228 10.6151
R1797 B.n232 B.n231 10.6151
R1798 B.n235 B.n232 10.6151
R1799 B.n236 B.n235 10.6151
R1800 B.n239 B.n236 10.6151
R1801 B.n240 B.n239 10.6151
R1802 B.n243 B.n240 10.6151
R1803 B.n244 B.n243 10.6151
R1804 B.n247 B.n244 10.6151
R1805 B.n248 B.n247 10.6151
R1806 B.n251 B.n248 10.6151
R1807 B.n252 B.n251 10.6151
R1808 B.n256 B.n255 10.6151
R1809 B.n259 B.n256 10.6151
R1810 B.n260 B.n259 10.6151
R1811 B.n263 B.n260 10.6151
R1812 B.n264 B.n263 10.6151
R1813 B.n267 B.n264 10.6151
R1814 B.n268 B.n267 10.6151
R1815 B.n271 B.n268 10.6151
R1816 B.n276 B.n273 10.6151
R1817 B.n277 B.n276 10.6151
R1818 B.n280 B.n277 10.6151
R1819 B.n281 B.n280 10.6151
R1820 B.n284 B.n281 10.6151
R1821 B.n285 B.n284 10.6151
R1822 B.n288 B.n285 10.6151
R1823 B.n289 B.n288 10.6151
R1824 B.n292 B.n289 10.6151
R1825 B.n293 B.n292 10.6151
R1826 B.n296 B.n293 10.6151
R1827 B.n297 B.n296 10.6151
R1828 B.n300 B.n297 10.6151
R1829 B.n301 B.n300 10.6151
R1830 B.n304 B.n301 10.6151
R1831 B.n305 B.n304 10.6151
R1832 B.n308 B.n305 10.6151
R1833 B.n309 B.n308 10.6151
R1834 B.n312 B.n309 10.6151
R1835 B.n313 B.n312 10.6151
R1836 B.n316 B.n313 10.6151
R1837 B.n317 B.n316 10.6151
R1838 B.n320 B.n317 10.6151
R1839 B.n321 B.n320 10.6151
R1840 B.n324 B.n321 10.6151
R1841 B.n325 B.n324 10.6151
R1842 B.n328 B.n325 10.6151
R1843 B.n329 B.n328 10.6151
R1844 B.n332 B.n329 10.6151
R1845 B.n333 B.n332 10.6151
R1846 B.n336 B.n333 10.6151
R1847 B.n337 B.n336 10.6151
R1848 B.n340 B.n337 10.6151
R1849 B.n341 B.n340 10.6151
R1850 B.n344 B.n341 10.6151
R1851 B.n345 B.n344 10.6151
R1852 B.n348 B.n345 10.6151
R1853 B.n349 B.n348 10.6151
R1854 B.n352 B.n349 10.6151
R1855 B.n353 B.n352 10.6151
R1856 B.n356 B.n353 10.6151
R1857 B.n357 B.n356 10.6151
R1858 B.n360 B.n357 10.6151
R1859 B.n361 B.n360 10.6151
R1860 B.n364 B.n361 10.6151
R1861 B.n365 B.n364 10.6151
R1862 B.n978 B.n365 10.6151
R1863 B.n1097 B.n0 8.11757
R1864 B.n1097 B.n1 8.11757
R1865 B.n810 B.t1 7.39259
R1866 B.n61 B.t0 7.39259
R1867 B.n645 B.n644 6.5566
R1868 B.n628 B.n530 6.5566
R1869 B.n255 B.n161 6.5566
R1870 B.n272 B.n271 6.5566
R1871 B.n646 B.n645 4.05904
R1872 B.n625 B.n530 4.05904
R1873 B.n252 B.n161 4.05904
R1874 B.n273 B.n272 4.05904
R1875 B.n768 B.t11 3.98086
R1876 B.t7 B.n1003 3.98086
R1877 B.n847 B.t3 2.84361
R1878 B.n40 B.t5 2.84361
R1879 B.t4 B.n376 1.70637
R1880 B.t2 B.n16 1.70637
R1881 VP.n16 VP.n13 161.3
R1882 VP.n18 VP.n17 161.3
R1883 VP.n19 VP.n12 161.3
R1884 VP.n21 VP.n20 161.3
R1885 VP.n22 VP.n11 161.3
R1886 VP.n24 VP.n23 161.3
R1887 VP.n25 VP.n10 161.3
R1888 VP.n27 VP.n26 161.3
R1889 VP.n56 VP.n55 161.3
R1890 VP.n54 VP.n1 161.3
R1891 VP.n53 VP.n52 161.3
R1892 VP.n51 VP.n2 161.3
R1893 VP.n50 VP.n49 161.3
R1894 VP.n48 VP.n3 161.3
R1895 VP.n47 VP.n46 161.3
R1896 VP.n45 VP.n4 161.3
R1897 VP.n44 VP.n43 161.3
R1898 VP.n42 VP.n5 161.3
R1899 VP.n41 VP.n40 161.3
R1900 VP.n39 VP.n6 161.3
R1901 VP.n38 VP.n37 161.3
R1902 VP.n36 VP.n7 161.3
R1903 VP.n35 VP.n34 161.3
R1904 VP.n33 VP.n8 161.3
R1905 VP.n32 VP.n31 161.3
R1906 VP.n15 VP.t4 124.061
R1907 VP.n43 VP.t1 91.3986
R1908 VP.n30 VP.t0 91.3986
R1909 VP.n0 VP.t5 91.3986
R1910 VP.n14 VP.t3 91.3986
R1911 VP.n9 VP.t2 91.3986
R1912 VP.n30 VP.n29 88.1101
R1913 VP.n57 VP.n0 88.1101
R1914 VP.n28 VP.n9 88.1101
R1915 VP.n29 VP.n28 54.613
R1916 VP.n15 VP.n14 50.4823
R1917 VP.n37 VP.n36 42.4359
R1918 VP.n49 VP.n2 42.4359
R1919 VP.n20 VP.n11 42.4359
R1920 VP.n37 VP.n6 38.5509
R1921 VP.n49 VP.n48 38.5509
R1922 VP.n20 VP.n19 38.5509
R1923 VP.n31 VP.n8 24.4675
R1924 VP.n35 VP.n8 24.4675
R1925 VP.n36 VP.n35 24.4675
R1926 VP.n41 VP.n6 24.4675
R1927 VP.n42 VP.n41 24.4675
R1928 VP.n43 VP.n42 24.4675
R1929 VP.n43 VP.n4 24.4675
R1930 VP.n47 VP.n4 24.4675
R1931 VP.n48 VP.n47 24.4675
R1932 VP.n53 VP.n2 24.4675
R1933 VP.n54 VP.n53 24.4675
R1934 VP.n55 VP.n54 24.4675
R1935 VP.n24 VP.n11 24.4675
R1936 VP.n25 VP.n24 24.4675
R1937 VP.n26 VP.n25 24.4675
R1938 VP.n14 VP.n13 24.4675
R1939 VP.n18 VP.n13 24.4675
R1940 VP.n19 VP.n18 24.4675
R1941 VP.n16 VP.n15 2.48381
R1942 VP.n31 VP.n30 1.95786
R1943 VP.n55 VP.n0 1.95786
R1944 VP.n26 VP.n9 1.95786
R1945 VP.n28 VP.n27 0.354971
R1946 VP.n32 VP.n29 0.354971
R1947 VP.n57 VP.n56 0.354971
R1948 VP VP.n57 0.26696
R1949 VP.n17 VP.n16 0.189894
R1950 VP.n17 VP.n12 0.189894
R1951 VP.n21 VP.n12 0.189894
R1952 VP.n22 VP.n21 0.189894
R1953 VP.n23 VP.n22 0.189894
R1954 VP.n23 VP.n10 0.189894
R1955 VP.n27 VP.n10 0.189894
R1956 VP.n33 VP.n32 0.189894
R1957 VP.n34 VP.n33 0.189894
R1958 VP.n34 VP.n7 0.189894
R1959 VP.n38 VP.n7 0.189894
R1960 VP.n39 VP.n38 0.189894
R1961 VP.n40 VP.n39 0.189894
R1962 VP.n40 VP.n5 0.189894
R1963 VP.n44 VP.n5 0.189894
R1964 VP.n45 VP.n44 0.189894
R1965 VP.n46 VP.n45 0.189894
R1966 VP.n46 VP.n3 0.189894
R1967 VP.n50 VP.n3 0.189894
R1968 VP.n51 VP.n50 0.189894
R1969 VP.n52 VP.n51 0.189894
R1970 VP.n52 VP.n1 0.189894
R1971 VP.n56 VP.n1 0.189894
R1972 VTAIL.n314 VTAIL.n242 289.615
R1973 VTAIL.n74 VTAIL.n2 289.615
R1974 VTAIL.n236 VTAIL.n164 289.615
R1975 VTAIL.n156 VTAIL.n84 289.615
R1976 VTAIL.n266 VTAIL.n265 185
R1977 VTAIL.n271 VTAIL.n270 185
R1978 VTAIL.n273 VTAIL.n272 185
R1979 VTAIL.n262 VTAIL.n261 185
R1980 VTAIL.n279 VTAIL.n278 185
R1981 VTAIL.n281 VTAIL.n280 185
R1982 VTAIL.n258 VTAIL.n257 185
R1983 VTAIL.n287 VTAIL.n286 185
R1984 VTAIL.n289 VTAIL.n288 185
R1985 VTAIL.n254 VTAIL.n253 185
R1986 VTAIL.n295 VTAIL.n294 185
R1987 VTAIL.n297 VTAIL.n296 185
R1988 VTAIL.n250 VTAIL.n249 185
R1989 VTAIL.n303 VTAIL.n302 185
R1990 VTAIL.n305 VTAIL.n304 185
R1991 VTAIL.n246 VTAIL.n245 185
R1992 VTAIL.n312 VTAIL.n311 185
R1993 VTAIL.n313 VTAIL.n244 185
R1994 VTAIL.n315 VTAIL.n314 185
R1995 VTAIL.n26 VTAIL.n25 185
R1996 VTAIL.n31 VTAIL.n30 185
R1997 VTAIL.n33 VTAIL.n32 185
R1998 VTAIL.n22 VTAIL.n21 185
R1999 VTAIL.n39 VTAIL.n38 185
R2000 VTAIL.n41 VTAIL.n40 185
R2001 VTAIL.n18 VTAIL.n17 185
R2002 VTAIL.n47 VTAIL.n46 185
R2003 VTAIL.n49 VTAIL.n48 185
R2004 VTAIL.n14 VTAIL.n13 185
R2005 VTAIL.n55 VTAIL.n54 185
R2006 VTAIL.n57 VTAIL.n56 185
R2007 VTAIL.n10 VTAIL.n9 185
R2008 VTAIL.n63 VTAIL.n62 185
R2009 VTAIL.n65 VTAIL.n64 185
R2010 VTAIL.n6 VTAIL.n5 185
R2011 VTAIL.n72 VTAIL.n71 185
R2012 VTAIL.n73 VTAIL.n4 185
R2013 VTAIL.n75 VTAIL.n74 185
R2014 VTAIL.n237 VTAIL.n236 185
R2015 VTAIL.n235 VTAIL.n166 185
R2016 VTAIL.n234 VTAIL.n233 185
R2017 VTAIL.n169 VTAIL.n167 185
R2018 VTAIL.n228 VTAIL.n227 185
R2019 VTAIL.n226 VTAIL.n225 185
R2020 VTAIL.n173 VTAIL.n172 185
R2021 VTAIL.n220 VTAIL.n219 185
R2022 VTAIL.n218 VTAIL.n217 185
R2023 VTAIL.n177 VTAIL.n176 185
R2024 VTAIL.n212 VTAIL.n211 185
R2025 VTAIL.n210 VTAIL.n209 185
R2026 VTAIL.n181 VTAIL.n180 185
R2027 VTAIL.n204 VTAIL.n203 185
R2028 VTAIL.n202 VTAIL.n201 185
R2029 VTAIL.n185 VTAIL.n184 185
R2030 VTAIL.n196 VTAIL.n195 185
R2031 VTAIL.n194 VTAIL.n193 185
R2032 VTAIL.n189 VTAIL.n188 185
R2033 VTAIL.n157 VTAIL.n156 185
R2034 VTAIL.n155 VTAIL.n86 185
R2035 VTAIL.n154 VTAIL.n153 185
R2036 VTAIL.n89 VTAIL.n87 185
R2037 VTAIL.n148 VTAIL.n147 185
R2038 VTAIL.n146 VTAIL.n145 185
R2039 VTAIL.n93 VTAIL.n92 185
R2040 VTAIL.n140 VTAIL.n139 185
R2041 VTAIL.n138 VTAIL.n137 185
R2042 VTAIL.n97 VTAIL.n96 185
R2043 VTAIL.n132 VTAIL.n131 185
R2044 VTAIL.n130 VTAIL.n129 185
R2045 VTAIL.n101 VTAIL.n100 185
R2046 VTAIL.n124 VTAIL.n123 185
R2047 VTAIL.n122 VTAIL.n121 185
R2048 VTAIL.n105 VTAIL.n104 185
R2049 VTAIL.n116 VTAIL.n115 185
R2050 VTAIL.n114 VTAIL.n113 185
R2051 VTAIL.n109 VTAIL.n108 185
R2052 VTAIL.n267 VTAIL.t0 147.659
R2053 VTAIL.n27 VTAIL.t9 147.659
R2054 VTAIL.n190 VTAIL.t7 147.659
R2055 VTAIL.n110 VTAIL.t11 147.659
R2056 VTAIL.n271 VTAIL.n265 104.615
R2057 VTAIL.n272 VTAIL.n271 104.615
R2058 VTAIL.n272 VTAIL.n261 104.615
R2059 VTAIL.n279 VTAIL.n261 104.615
R2060 VTAIL.n280 VTAIL.n279 104.615
R2061 VTAIL.n280 VTAIL.n257 104.615
R2062 VTAIL.n287 VTAIL.n257 104.615
R2063 VTAIL.n288 VTAIL.n287 104.615
R2064 VTAIL.n288 VTAIL.n253 104.615
R2065 VTAIL.n295 VTAIL.n253 104.615
R2066 VTAIL.n296 VTAIL.n295 104.615
R2067 VTAIL.n296 VTAIL.n249 104.615
R2068 VTAIL.n303 VTAIL.n249 104.615
R2069 VTAIL.n304 VTAIL.n303 104.615
R2070 VTAIL.n304 VTAIL.n245 104.615
R2071 VTAIL.n312 VTAIL.n245 104.615
R2072 VTAIL.n313 VTAIL.n312 104.615
R2073 VTAIL.n314 VTAIL.n313 104.615
R2074 VTAIL.n31 VTAIL.n25 104.615
R2075 VTAIL.n32 VTAIL.n31 104.615
R2076 VTAIL.n32 VTAIL.n21 104.615
R2077 VTAIL.n39 VTAIL.n21 104.615
R2078 VTAIL.n40 VTAIL.n39 104.615
R2079 VTAIL.n40 VTAIL.n17 104.615
R2080 VTAIL.n47 VTAIL.n17 104.615
R2081 VTAIL.n48 VTAIL.n47 104.615
R2082 VTAIL.n48 VTAIL.n13 104.615
R2083 VTAIL.n55 VTAIL.n13 104.615
R2084 VTAIL.n56 VTAIL.n55 104.615
R2085 VTAIL.n56 VTAIL.n9 104.615
R2086 VTAIL.n63 VTAIL.n9 104.615
R2087 VTAIL.n64 VTAIL.n63 104.615
R2088 VTAIL.n64 VTAIL.n5 104.615
R2089 VTAIL.n72 VTAIL.n5 104.615
R2090 VTAIL.n73 VTAIL.n72 104.615
R2091 VTAIL.n74 VTAIL.n73 104.615
R2092 VTAIL.n236 VTAIL.n235 104.615
R2093 VTAIL.n235 VTAIL.n234 104.615
R2094 VTAIL.n234 VTAIL.n167 104.615
R2095 VTAIL.n227 VTAIL.n167 104.615
R2096 VTAIL.n227 VTAIL.n226 104.615
R2097 VTAIL.n226 VTAIL.n172 104.615
R2098 VTAIL.n219 VTAIL.n172 104.615
R2099 VTAIL.n219 VTAIL.n218 104.615
R2100 VTAIL.n218 VTAIL.n176 104.615
R2101 VTAIL.n211 VTAIL.n176 104.615
R2102 VTAIL.n211 VTAIL.n210 104.615
R2103 VTAIL.n210 VTAIL.n180 104.615
R2104 VTAIL.n203 VTAIL.n180 104.615
R2105 VTAIL.n203 VTAIL.n202 104.615
R2106 VTAIL.n202 VTAIL.n184 104.615
R2107 VTAIL.n195 VTAIL.n184 104.615
R2108 VTAIL.n195 VTAIL.n194 104.615
R2109 VTAIL.n194 VTAIL.n188 104.615
R2110 VTAIL.n156 VTAIL.n155 104.615
R2111 VTAIL.n155 VTAIL.n154 104.615
R2112 VTAIL.n154 VTAIL.n87 104.615
R2113 VTAIL.n147 VTAIL.n87 104.615
R2114 VTAIL.n147 VTAIL.n146 104.615
R2115 VTAIL.n146 VTAIL.n92 104.615
R2116 VTAIL.n139 VTAIL.n92 104.615
R2117 VTAIL.n139 VTAIL.n138 104.615
R2118 VTAIL.n138 VTAIL.n96 104.615
R2119 VTAIL.n131 VTAIL.n96 104.615
R2120 VTAIL.n131 VTAIL.n130 104.615
R2121 VTAIL.n130 VTAIL.n100 104.615
R2122 VTAIL.n123 VTAIL.n100 104.615
R2123 VTAIL.n123 VTAIL.n122 104.615
R2124 VTAIL.n122 VTAIL.n104 104.615
R2125 VTAIL.n115 VTAIL.n104 104.615
R2126 VTAIL.n115 VTAIL.n114 104.615
R2127 VTAIL.n114 VTAIL.n108 104.615
R2128 VTAIL.t0 VTAIL.n265 52.3082
R2129 VTAIL.t9 VTAIL.n25 52.3082
R2130 VTAIL.t7 VTAIL.n188 52.3082
R2131 VTAIL.t11 VTAIL.n108 52.3082
R2132 VTAIL.n163 VTAIL.n162 47.2447
R2133 VTAIL.n83 VTAIL.n82 47.2447
R2134 VTAIL.n1 VTAIL.n0 47.2445
R2135 VTAIL.n81 VTAIL.n80 47.2445
R2136 VTAIL.n319 VTAIL.n318 35.0944
R2137 VTAIL.n79 VTAIL.n78 35.0944
R2138 VTAIL.n241 VTAIL.n240 35.0944
R2139 VTAIL.n161 VTAIL.n160 35.0944
R2140 VTAIL.n83 VTAIL.n81 31.4617
R2141 VTAIL.n319 VTAIL.n241 27.9789
R2142 VTAIL.n267 VTAIL.n266 15.6677
R2143 VTAIL.n27 VTAIL.n26 15.6677
R2144 VTAIL.n190 VTAIL.n189 15.6677
R2145 VTAIL.n110 VTAIL.n109 15.6677
R2146 VTAIL.n315 VTAIL.n244 13.1884
R2147 VTAIL.n75 VTAIL.n4 13.1884
R2148 VTAIL.n237 VTAIL.n166 13.1884
R2149 VTAIL.n157 VTAIL.n86 13.1884
R2150 VTAIL.n270 VTAIL.n269 12.8005
R2151 VTAIL.n311 VTAIL.n310 12.8005
R2152 VTAIL.n316 VTAIL.n242 12.8005
R2153 VTAIL.n30 VTAIL.n29 12.8005
R2154 VTAIL.n71 VTAIL.n70 12.8005
R2155 VTAIL.n76 VTAIL.n2 12.8005
R2156 VTAIL.n238 VTAIL.n164 12.8005
R2157 VTAIL.n233 VTAIL.n168 12.8005
R2158 VTAIL.n193 VTAIL.n192 12.8005
R2159 VTAIL.n158 VTAIL.n84 12.8005
R2160 VTAIL.n153 VTAIL.n88 12.8005
R2161 VTAIL.n113 VTAIL.n112 12.8005
R2162 VTAIL.n273 VTAIL.n264 12.0247
R2163 VTAIL.n309 VTAIL.n246 12.0247
R2164 VTAIL.n33 VTAIL.n24 12.0247
R2165 VTAIL.n69 VTAIL.n6 12.0247
R2166 VTAIL.n232 VTAIL.n169 12.0247
R2167 VTAIL.n196 VTAIL.n187 12.0247
R2168 VTAIL.n152 VTAIL.n89 12.0247
R2169 VTAIL.n116 VTAIL.n107 12.0247
R2170 VTAIL.n274 VTAIL.n262 11.249
R2171 VTAIL.n306 VTAIL.n305 11.249
R2172 VTAIL.n34 VTAIL.n22 11.249
R2173 VTAIL.n66 VTAIL.n65 11.249
R2174 VTAIL.n229 VTAIL.n228 11.249
R2175 VTAIL.n197 VTAIL.n185 11.249
R2176 VTAIL.n149 VTAIL.n148 11.249
R2177 VTAIL.n117 VTAIL.n105 11.249
R2178 VTAIL.n278 VTAIL.n277 10.4732
R2179 VTAIL.n302 VTAIL.n248 10.4732
R2180 VTAIL.n38 VTAIL.n37 10.4732
R2181 VTAIL.n62 VTAIL.n8 10.4732
R2182 VTAIL.n225 VTAIL.n171 10.4732
R2183 VTAIL.n201 VTAIL.n200 10.4732
R2184 VTAIL.n145 VTAIL.n91 10.4732
R2185 VTAIL.n121 VTAIL.n120 10.4732
R2186 VTAIL.n281 VTAIL.n260 9.69747
R2187 VTAIL.n301 VTAIL.n250 9.69747
R2188 VTAIL.n41 VTAIL.n20 9.69747
R2189 VTAIL.n61 VTAIL.n10 9.69747
R2190 VTAIL.n224 VTAIL.n173 9.69747
R2191 VTAIL.n204 VTAIL.n183 9.69747
R2192 VTAIL.n144 VTAIL.n93 9.69747
R2193 VTAIL.n124 VTAIL.n103 9.69747
R2194 VTAIL.n318 VTAIL.n317 9.45567
R2195 VTAIL.n78 VTAIL.n77 9.45567
R2196 VTAIL.n240 VTAIL.n239 9.45567
R2197 VTAIL.n160 VTAIL.n159 9.45567
R2198 VTAIL.n317 VTAIL.n316 9.3005
R2199 VTAIL.n256 VTAIL.n255 9.3005
R2200 VTAIL.n285 VTAIL.n284 9.3005
R2201 VTAIL.n283 VTAIL.n282 9.3005
R2202 VTAIL.n260 VTAIL.n259 9.3005
R2203 VTAIL.n277 VTAIL.n276 9.3005
R2204 VTAIL.n275 VTAIL.n274 9.3005
R2205 VTAIL.n264 VTAIL.n263 9.3005
R2206 VTAIL.n269 VTAIL.n268 9.3005
R2207 VTAIL.n291 VTAIL.n290 9.3005
R2208 VTAIL.n293 VTAIL.n292 9.3005
R2209 VTAIL.n252 VTAIL.n251 9.3005
R2210 VTAIL.n299 VTAIL.n298 9.3005
R2211 VTAIL.n301 VTAIL.n300 9.3005
R2212 VTAIL.n248 VTAIL.n247 9.3005
R2213 VTAIL.n307 VTAIL.n306 9.3005
R2214 VTAIL.n309 VTAIL.n308 9.3005
R2215 VTAIL.n310 VTAIL.n243 9.3005
R2216 VTAIL.n77 VTAIL.n76 9.3005
R2217 VTAIL.n16 VTAIL.n15 9.3005
R2218 VTAIL.n45 VTAIL.n44 9.3005
R2219 VTAIL.n43 VTAIL.n42 9.3005
R2220 VTAIL.n20 VTAIL.n19 9.3005
R2221 VTAIL.n37 VTAIL.n36 9.3005
R2222 VTAIL.n35 VTAIL.n34 9.3005
R2223 VTAIL.n24 VTAIL.n23 9.3005
R2224 VTAIL.n29 VTAIL.n28 9.3005
R2225 VTAIL.n51 VTAIL.n50 9.3005
R2226 VTAIL.n53 VTAIL.n52 9.3005
R2227 VTAIL.n12 VTAIL.n11 9.3005
R2228 VTAIL.n59 VTAIL.n58 9.3005
R2229 VTAIL.n61 VTAIL.n60 9.3005
R2230 VTAIL.n8 VTAIL.n7 9.3005
R2231 VTAIL.n67 VTAIL.n66 9.3005
R2232 VTAIL.n69 VTAIL.n68 9.3005
R2233 VTAIL.n70 VTAIL.n3 9.3005
R2234 VTAIL.n216 VTAIL.n215 9.3005
R2235 VTAIL.n175 VTAIL.n174 9.3005
R2236 VTAIL.n222 VTAIL.n221 9.3005
R2237 VTAIL.n224 VTAIL.n223 9.3005
R2238 VTAIL.n171 VTAIL.n170 9.3005
R2239 VTAIL.n230 VTAIL.n229 9.3005
R2240 VTAIL.n232 VTAIL.n231 9.3005
R2241 VTAIL.n168 VTAIL.n165 9.3005
R2242 VTAIL.n239 VTAIL.n238 9.3005
R2243 VTAIL.n214 VTAIL.n213 9.3005
R2244 VTAIL.n179 VTAIL.n178 9.3005
R2245 VTAIL.n208 VTAIL.n207 9.3005
R2246 VTAIL.n206 VTAIL.n205 9.3005
R2247 VTAIL.n183 VTAIL.n182 9.3005
R2248 VTAIL.n200 VTAIL.n199 9.3005
R2249 VTAIL.n198 VTAIL.n197 9.3005
R2250 VTAIL.n187 VTAIL.n186 9.3005
R2251 VTAIL.n192 VTAIL.n191 9.3005
R2252 VTAIL.n136 VTAIL.n135 9.3005
R2253 VTAIL.n95 VTAIL.n94 9.3005
R2254 VTAIL.n142 VTAIL.n141 9.3005
R2255 VTAIL.n144 VTAIL.n143 9.3005
R2256 VTAIL.n91 VTAIL.n90 9.3005
R2257 VTAIL.n150 VTAIL.n149 9.3005
R2258 VTAIL.n152 VTAIL.n151 9.3005
R2259 VTAIL.n88 VTAIL.n85 9.3005
R2260 VTAIL.n159 VTAIL.n158 9.3005
R2261 VTAIL.n134 VTAIL.n133 9.3005
R2262 VTAIL.n99 VTAIL.n98 9.3005
R2263 VTAIL.n128 VTAIL.n127 9.3005
R2264 VTAIL.n126 VTAIL.n125 9.3005
R2265 VTAIL.n103 VTAIL.n102 9.3005
R2266 VTAIL.n120 VTAIL.n119 9.3005
R2267 VTAIL.n118 VTAIL.n117 9.3005
R2268 VTAIL.n107 VTAIL.n106 9.3005
R2269 VTAIL.n112 VTAIL.n111 9.3005
R2270 VTAIL.n282 VTAIL.n258 8.92171
R2271 VTAIL.n298 VTAIL.n297 8.92171
R2272 VTAIL.n42 VTAIL.n18 8.92171
R2273 VTAIL.n58 VTAIL.n57 8.92171
R2274 VTAIL.n221 VTAIL.n220 8.92171
R2275 VTAIL.n205 VTAIL.n181 8.92171
R2276 VTAIL.n141 VTAIL.n140 8.92171
R2277 VTAIL.n125 VTAIL.n101 8.92171
R2278 VTAIL.n286 VTAIL.n285 8.14595
R2279 VTAIL.n294 VTAIL.n252 8.14595
R2280 VTAIL.n46 VTAIL.n45 8.14595
R2281 VTAIL.n54 VTAIL.n12 8.14595
R2282 VTAIL.n217 VTAIL.n175 8.14595
R2283 VTAIL.n209 VTAIL.n208 8.14595
R2284 VTAIL.n137 VTAIL.n95 8.14595
R2285 VTAIL.n129 VTAIL.n128 8.14595
R2286 VTAIL.n289 VTAIL.n256 7.3702
R2287 VTAIL.n293 VTAIL.n254 7.3702
R2288 VTAIL.n49 VTAIL.n16 7.3702
R2289 VTAIL.n53 VTAIL.n14 7.3702
R2290 VTAIL.n216 VTAIL.n177 7.3702
R2291 VTAIL.n212 VTAIL.n179 7.3702
R2292 VTAIL.n136 VTAIL.n97 7.3702
R2293 VTAIL.n132 VTAIL.n99 7.3702
R2294 VTAIL.n290 VTAIL.n289 6.59444
R2295 VTAIL.n290 VTAIL.n254 6.59444
R2296 VTAIL.n50 VTAIL.n49 6.59444
R2297 VTAIL.n50 VTAIL.n14 6.59444
R2298 VTAIL.n213 VTAIL.n177 6.59444
R2299 VTAIL.n213 VTAIL.n212 6.59444
R2300 VTAIL.n133 VTAIL.n97 6.59444
R2301 VTAIL.n133 VTAIL.n132 6.59444
R2302 VTAIL.n286 VTAIL.n256 5.81868
R2303 VTAIL.n294 VTAIL.n293 5.81868
R2304 VTAIL.n46 VTAIL.n16 5.81868
R2305 VTAIL.n54 VTAIL.n53 5.81868
R2306 VTAIL.n217 VTAIL.n216 5.81868
R2307 VTAIL.n209 VTAIL.n179 5.81868
R2308 VTAIL.n137 VTAIL.n136 5.81868
R2309 VTAIL.n129 VTAIL.n99 5.81868
R2310 VTAIL.n285 VTAIL.n258 5.04292
R2311 VTAIL.n297 VTAIL.n252 5.04292
R2312 VTAIL.n45 VTAIL.n18 5.04292
R2313 VTAIL.n57 VTAIL.n12 5.04292
R2314 VTAIL.n220 VTAIL.n175 5.04292
R2315 VTAIL.n208 VTAIL.n181 5.04292
R2316 VTAIL.n140 VTAIL.n95 5.04292
R2317 VTAIL.n128 VTAIL.n101 5.04292
R2318 VTAIL.n268 VTAIL.n267 4.38563
R2319 VTAIL.n28 VTAIL.n27 4.38563
R2320 VTAIL.n191 VTAIL.n190 4.38563
R2321 VTAIL.n111 VTAIL.n110 4.38563
R2322 VTAIL.n282 VTAIL.n281 4.26717
R2323 VTAIL.n298 VTAIL.n250 4.26717
R2324 VTAIL.n42 VTAIL.n41 4.26717
R2325 VTAIL.n58 VTAIL.n10 4.26717
R2326 VTAIL.n221 VTAIL.n173 4.26717
R2327 VTAIL.n205 VTAIL.n204 4.26717
R2328 VTAIL.n141 VTAIL.n93 4.26717
R2329 VTAIL.n125 VTAIL.n124 4.26717
R2330 VTAIL.n278 VTAIL.n260 3.49141
R2331 VTAIL.n302 VTAIL.n301 3.49141
R2332 VTAIL.n38 VTAIL.n20 3.49141
R2333 VTAIL.n62 VTAIL.n61 3.49141
R2334 VTAIL.n225 VTAIL.n224 3.49141
R2335 VTAIL.n201 VTAIL.n183 3.49141
R2336 VTAIL.n145 VTAIL.n144 3.49141
R2337 VTAIL.n121 VTAIL.n103 3.49141
R2338 VTAIL.n161 VTAIL.n83 3.48326
R2339 VTAIL.n241 VTAIL.n163 3.48326
R2340 VTAIL.n81 VTAIL.n79 3.48326
R2341 VTAIL.n277 VTAIL.n262 2.71565
R2342 VTAIL.n305 VTAIL.n248 2.71565
R2343 VTAIL.n37 VTAIL.n22 2.71565
R2344 VTAIL.n65 VTAIL.n8 2.71565
R2345 VTAIL.n228 VTAIL.n171 2.71565
R2346 VTAIL.n200 VTAIL.n185 2.71565
R2347 VTAIL.n148 VTAIL.n91 2.71565
R2348 VTAIL.n120 VTAIL.n105 2.71565
R2349 VTAIL VTAIL.n319 2.55438
R2350 VTAIL.n163 VTAIL.n161 2.21171
R2351 VTAIL.n79 VTAIL.n1 2.21171
R2352 VTAIL.n274 VTAIL.n273 1.93989
R2353 VTAIL.n306 VTAIL.n246 1.93989
R2354 VTAIL.n34 VTAIL.n33 1.93989
R2355 VTAIL.n66 VTAIL.n6 1.93989
R2356 VTAIL.n229 VTAIL.n169 1.93989
R2357 VTAIL.n197 VTAIL.n196 1.93989
R2358 VTAIL.n149 VTAIL.n89 1.93989
R2359 VTAIL.n117 VTAIL.n116 1.93989
R2360 VTAIL.n0 VTAIL.t2 1.40775
R2361 VTAIL.n0 VTAIL.t3 1.40775
R2362 VTAIL.n80 VTAIL.t5 1.40775
R2363 VTAIL.n80 VTAIL.t6 1.40775
R2364 VTAIL.n162 VTAIL.t10 1.40775
R2365 VTAIL.n162 VTAIL.t8 1.40775
R2366 VTAIL.n82 VTAIL.t1 1.40775
R2367 VTAIL.n82 VTAIL.t4 1.40775
R2368 VTAIL.n270 VTAIL.n264 1.16414
R2369 VTAIL.n311 VTAIL.n309 1.16414
R2370 VTAIL.n318 VTAIL.n242 1.16414
R2371 VTAIL.n30 VTAIL.n24 1.16414
R2372 VTAIL.n71 VTAIL.n69 1.16414
R2373 VTAIL.n78 VTAIL.n2 1.16414
R2374 VTAIL.n240 VTAIL.n164 1.16414
R2375 VTAIL.n233 VTAIL.n232 1.16414
R2376 VTAIL.n193 VTAIL.n187 1.16414
R2377 VTAIL.n160 VTAIL.n84 1.16414
R2378 VTAIL.n153 VTAIL.n152 1.16414
R2379 VTAIL.n113 VTAIL.n107 1.16414
R2380 VTAIL VTAIL.n1 0.929379
R2381 VTAIL.n269 VTAIL.n266 0.388379
R2382 VTAIL.n310 VTAIL.n244 0.388379
R2383 VTAIL.n316 VTAIL.n315 0.388379
R2384 VTAIL.n29 VTAIL.n26 0.388379
R2385 VTAIL.n70 VTAIL.n4 0.388379
R2386 VTAIL.n76 VTAIL.n75 0.388379
R2387 VTAIL.n238 VTAIL.n237 0.388379
R2388 VTAIL.n168 VTAIL.n166 0.388379
R2389 VTAIL.n192 VTAIL.n189 0.388379
R2390 VTAIL.n158 VTAIL.n157 0.388379
R2391 VTAIL.n88 VTAIL.n86 0.388379
R2392 VTAIL.n112 VTAIL.n109 0.388379
R2393 VTAIL.n268 VTAIL.n263 0.155672
R2394 VTAIL.n275 VTAIL.n263 0.155672
R2395 VTAIL.n276 VTAIL.n275 0.155672
R2396 VTAIL.n276 VTAIL.n259 0.155672
R2397 VTAIL.n283 VTAIL.n259 0.155672
R2398 VTAIL.n284 VTAIL.n283 0.155672
R2399 VTAIL.n284 VTAIL.n255 0.155672
R2400 VTAIL.n291 VTAIL.n255 0.155672
R2401 VTAIL.n292 VTAIL.n291 0.155672
R2402 VTAIL.n292 VTAIL.n251 0.155672
R2403 VTAIL.n299 VTAIL.n251 0.155672
R2404 VTAIL.n300 VTAIL.n299 0.155672
R2405 VTAIL.n300 VTAIL.n247 0.155672
R2406 VTAIL.n307 VTAIL.n247 0.155672
R2407 VTAIL.n308 VTAIL.n307 0.155672
R2408 VTAIL.n308 VTAIL.n243 0.155672
R2409 VTAIL.n317 VTAIL.n243 0.155672
R2410 VTAIL.n28 VTAIL.n23 0.155672
R2411 VTAIL.n35 VTAIL.n23 0.155672
R2412 VTAIL.n36 VTAIL.n35 0.155672
R2413 VTAIL.n36 VTAIL.n19 0.155672
R2414 VTAIL.n43 VTAIL.n19 0.155672
R2415 VTAIL.n44 VTAIL.n43 0.155672
R2416 VTAIL.n44 VTAIL.n15 0.155672
R2417 VTAIL.n51 VTAIL.n15 0.155672
R2418 VTAIL.n52 VTAIL.n51 0.155672
R2419 VTAIL.n52 VTAIL.n11 0.155672
R2420 VTAIL.n59 VTAIL.n11 0.155672
R2421 VTAIL.n60 VTAIL.n59 0.155672
R2422 VTAIL.n60 VTAIL.n7 0.155672
R2423 VTAIL.n67 VTAIL.n7 0.155672
R2424 VTAIL.n68 VTAIL.n67 0.155672
R2425 VTAIL.n68 VTAIL.n3 0.155672
R2426 VTAIL.n77 VTAIL.n3 0.155672
R2427 VTAIL.n239 VTAIL.n165 0.155672
R2428 VTAIL.n231 VTAIL.n165 0.155672
R2429 VTAIL.n231 VTAIL.n230 0.155672
R2430 VTAIL.n230 VTAIL.n170 0.155672
R2431 VTAIL.n223 VTAIL.n170 0.155672
R2432 VTAIL.n223 VTAIL.n222 0.155672
R2433 VTAIL.n222 VTAIL.n174 0.155672
R2434 VTAIL.n215 VTAIL.n174 0.155672
R2435 VTAIL.n215 VTAIL.n214 0.155672
R2436 VTAIL.n214 VTAIL.n178 0.155672
R2437 VTAIL.n207 VTAIL.n178 0.155672
R2438 VTAIL.n207 VTAIL.n206 0.155672
R2439 VTAIL.n206 VTAIL.n182 0.155672
R2440 VTAIL.n199 VTAIL.n182 0.155672
R2441 VTAIL.n199 VTAIL.n198 0.155672
R2442 VTAIL.n198 VTAIL.n186 0.155672
R2443 VTAIL.n191 VTAIL.n186 0.155672
R2444 VTAIL.n159 VTAIL.n85 0.155672
R2445 VTAIL.n151 VTAIL.n85 0.155672
R2446 VTAIL.n151 VTAIL.n150 0.155672
R2447 VTAIL.n150 VTAIL.n90 0.155672
R2448 VTAIL.n143 VTAIL.n90 0.155672
R2449 VTAIL.n143 VTAIL.n142 0.155672
R2450 VTAIL.n142 VTAIL.n94 0.155672
R2451 VTAIL.n135 VTAIL.n94 0.155672
R2452 VTAIL.n135 VTAIL.n134 0.155672
R2453 VTAIL.n134 VTAIL.n98 0.155672
R2454 VTAIL.n127 VTAIL.n98 0.155672
R2455 VTAIL.n127 VTAIL.n126 0.155672
R2456 VTAIL.n126 VTAIL.n102 0.155672
R2457 VTAIL.n119 VTAIL.n102 0.155672
R2458 VTAIL.n119 VTAIL.n118 0.155672
R2459 VTAIL.n118 VTAIL.n106 0.155672
R2460 VTAIL.n111 VTAIL.n106 0.155672
R2461 VDD1.n72 VDD1.n0 289.615
R2462 VDD1.n149 VDD1.n77 289.615
R2463 VDD1.n73 VDD1.n72 185
R2464 VDD1.n71 VDD1.n2 185
R2465 VDD1.n70 VDD1.n69 185
R2466 VDD1.n5 VDD1.n3 185
R2467 VDD1.n64 VDD1.n63 185
R2468 VDD1.n62 VDD1.n61 185
R2469 VDD1.n9 VDD1.n8 185
R2470 VDD1.n56 VDD1.n55 185
R2471 VDD1.n54 VDD1.n53 185
R2472 VDD1.n13 VDD1.n12 185
R2473 VDD1.n48 VDD1.n47 185
R2474 VDD1.n46 VDD1.n45 185
R2475 VDD1.n17 VDD1.n16 185
R2476 VDD1.n40 VDD1.n39 185
R2477 VDD1.n38 VDD1.n37 185
R2478 VDD1.n21 VDD1.n20 185
R2479 VDD1.n32 VDD1.n31 185
R2480 VDD1.n30 VDD1.n29 185
R2481 VDD1.n25 VDD1.n24 185
R2482 VDD1.n101 VDD1.n100 185
R2483 VDD1.n106 VDD1.n105 185
R2484 VDD1.n108 VDD1.n107 185
R2485 VDD1.n97 VDD1.n96 185
R2486 VDD1.n114 VDD1.n113 185
R2487 VDD1.n116 VDD1.n115 185
R2488 VDD1.n93 VDD1.n92 185
R2489 VDD1.n122 VDD1.n121 185
R2490 VDD1.n124 VDD1.n123 185
R2491 VDD1.n89 VDD1.n88 185
R2492 VDD1.n130 VDD1.n129 185
R2493 VDD1.n132 VDD1.n131 185
R2494 VDD1.n85 VDD1.n84 185
R2495 VDD1.n138 VDD1.n137 185
R2496 VDD1.n140 VDD1.n139 185
R2497 VDD1.n81 VDD1.n80 185
R2498 VDD1.n147 VDD1.n146 185
R2499 VDD1.n148 VDD1.n79 185
R2500 VDD1.n150 VDD1.n149 185
R2501 VDD1.n26 VDD1.t1 147.659
R2502 VDD1.n102 VDD1.t5 147.659
R2503 VDD1.n72 VDD1.n71 104.615
R2504 VDD1.n71 VDD1.n70 104.615
R2505 VDD1.n70 VDD1.n3 104.615
R2506 VDD1.n63 VDD1.n3 104.615
R2507 VDD1.n63 VDD1.n62 104.615
R2508 VDD1.n62 VDD1.n8 104.615
R2509 VDD1.n55 VDD1.n8 104.615
R2510 VDD1.n55 VDD1.n54 104.615
R2511 VDD1.n54 VDD1.n12 104.615
R2512 VDD1.n47 VDD1.n12 104.615
R2513 VDD1.n47 VDD1.n46 104.615
R2514 VDD1.n46 VDD1.n16 104.615
R2515 VDD1.n39 VDD1.n16 104.615
R2516 VDD1.n39 VDD1.n38 104.615
R2517 VDD1.n38 VDD1.n20 104.615
R2518 VDD1.n31 VDD1.n20 104.615
R2519 VDD1.n31 VDD1.n30 104.615
R2520 VDD1.n30 VDD1.n24 104.615
R2521 VDD1.n106 VDD1.n100 104.615
R2522 VDD1.n107 VDD1.n106 104.615
R2523 VDD1.n107 VDD1.n96 104.615
R2524 VDD1.n114 VDD1.n96 104.615
R2525 VDD1.n115 VDD1.n114 104.615
R2526 VDD1.n115 VDD1.n92 104.615
R2527 VDD1.n122 VDD1.n92 104.615
R2528 VDD1.n123 VDD1.n122 104.615
R2529 VDD1.n123 VDD1.n88 104.615
R2530 VDD1.n130 VDD1.n88 104.615
R2531 VDD1.n131 VDD1.n130 104.615
R2532 VDD1.n131 VDD1.n84 104.615
R2533 VDD1.n138 VDD1.n84 104.615
R2534 VDD1.n139 VDD1.n138 104.615
R2535 VDD1.n139 VDD1.n80 104.615
R2536 VDD1.n147 VDD1.n80 104.615
R2537 VDD1.n148 VDD1.n147 104.615
R2538 VDD1.n149 VDD1.n148 104.615
R2539 VDD1.n155 VDD1.n154 64.7387
R2540 VDD1.n157 VDD1.n156 63.9233
R2541 VDD1 VDD1.n76 54.4435
R2542 VDD1.n155 VDD1.n153 54.3299
R2543 VDD1.t1 VDD1.n24 52.3082
R2544 VDD1.t5 VDD1.n100 52.3082
R2545 VDD1.n157 VDD1.n155 49.488
R2546 VDD1.n26 VDD1.n25 15.6677
R2547 VDD1.n102 VDD1.n101 15.6677
R2548 VDD1.n73 VDD1.n2 13.1884
R2549 VDD1.n150 VDD1.n79 13.1884
R2550 VDD1.n74 VDD1.n0 12.8005
R2551 VDD1.n69 VDD1.n4 12.8005
R2552 VDD1.n29 VDD1.n28 12.8005
R2553 VDD1.n105 VDD1.n104 12.8005
R2554 VDD1.n146 VDD1.n145 12.8005
R2555 VDD1.n151 VDD1.n77 12.8005
R2556 VDD1.n68 VDD1.n5 12.0247
R2557 VDD1.n32 VDD1.n23 12.0247
R2558 VDD1.n108 VDD1.n99 12.0247
R2559 VDD1.n144 VDD1.n81 12.0247
R2560 VDD1.n65 VDD1.n64 11.249
R2561 VDD1.n33 VDD1.n21 11.249
R2562 VDD1.n109 VDD1.n97 11.249
R2563 VDD1.n141 VDD1.n140 11.249
R2564 VDD1.n61 VDD1.n7 10.4732
R2565 VDD1.n37 VDD1.n36 10.4732
R2566 VDD1.n113 VDD1.n112 10.4732
R2567 VDD1.n137 VDD1.n83 10.4732
R2568 VDD1.n60 VDD1.n9 9.69747
R2569 VDD1.n40 VDD1.n19 9.69747
R2570 VDD1.n116 VDD1.n95 9.69747
R2571 VDD1.n136 VDD1.n85 9.69747
R2572 VDD1.n76 VDD1.n75 9.45567
R2573 VDD1.n153 VDD1.n152 9.45567
R2574 VDD1.n52 VDD1.n51 9.3005
R2575 VDD1.n11 VDD1.n10 9.3005
R2576 VDD1.n58 VDD1.n57 9.3005
R2577 VDD1.n60 VDD1.n59 9.3005
R2578 VDD1.n7 VDD1.n6 9.3005
R2579 VDD1.n66 VDD1.n65 9.3005
R2580 VDD1.n68 VDD1.n67 9.3005
R2581 VDD1.n4 VDD1.n1 9.3005
R2582 VDD1.n75 VDD1.n74 9.3005
R2583 VDD1.n50 VDD1.n49 9.3005
R2584 VDD1.n15 VDD1.n14 9.3005
R2585 VDD1.n44 VDD1.n43 9.3005
R2586 VDD1.n42 VDD1.n41 9.3005
R2587 VDD1.n19 VDD1.n18 9.3005
R2588 VDD1.n36 VDD1.n35 9.3005
R2589 VDD1.n34 VDD1.n33 9.3005
R2590 VDD1.n23 VDD1.n22 9.3005
R2591 VDD1.n28 VDD1.n27 9.3005
R2592 VDD1.n152 VDD1.n151 9.3005
R2593 VDD1.n91 VDD1.n90 9.3005
R2594 VDD1.n120 VDD1.n119 9.3005
R2595 VDD1.n118 VDD1.n117 9.3005
R2596 VDD1.n95 VDD1.n94 9.3005
R2597 VDD1.n112 VDD1.n111 9.3005
R2598 VDD1.n110 VDD1.n109 9.3005
R2599 VDD1.n99 VDD1.n98 9.3005
R2600 VDD1.n104 VDD1.n103 9.3005
R2601 VDD1.n126 VDD1.n125 9.3005
R2602 VDD1.n128 VDD1.n127 9.3005
R2603 VDD1.n87 VDD1.n86 9.3005
R2604 VDD1.n134 VDD1.n133 9.3005
R2605 VDD1.n136 VDD1.n135 9.3005
R2606 VDD1.n83 VDD1.n82 9.3005
R2607 VDD1.n142 VDD1.n141 9.3005
R2608 VDD1.n144 VDD1.n143 9.3005
R2609 VDD1.n145 VDD1.n78 9.3005
R2610 VDD1.n57 VDD1.n56 8.92171
R2611 VDD1.n41 VDD1.n17 8.92171
R2612 VDD1.n117 VDD1.n93 8.92171
R2613 VDD1.n133 VDD1.n132 8.92171
R2614 VDD1.n53 VDD1.n11 8.14595
R2615 VDD1.n45 VDD1.n44 8.14595
R2616 VDD1.n121 VDD1.n120 8.14595
R2617 VDD1.n129 VDD1.n87 8.14595
R2618 VDD1.n52 VDD1.n13 7.3702
R2619 VDD1.n48 VDD1.n15 7.3702
R2620 VDD1.n124 VDD1.n91 7.3702
R2621 VDD1.n128 VDD1.n89 7.3702
R2622 VDD1.n49 VDD1.n13 6.59444
R2623 VDD1.n49 VDD1.n48 6.59444
R2624 VDD1.n125 VDD1.n124 6.59444
R2625 VDD1.n125 VDD1.n89 6.59444
R2626 VDD1.n53 VDD1.n52 5.81868
R2627 VDD1.n45 VDD1.n15 5.81868
R2628 VDD1.n121 VDD1.n91 5.81868
R2629 VDD1.n129 VDD1.n128 5.81868
R2630 VDD1.n56 VDD1.n11 5.04292
R2631 VDD1.n44 VDD1.n17 5.04292
R2632 VDD1.n120 VDD1.n93 5.04292
R2633 VDD1.n132 VDD1.n87 5.04292
R2634 VDD1.n27 VDD1.n26 4.38563
R2635 VDD1.n103 VDD1.n102 4.38563
R2636 VDD1.n57 VDD1.n9 4.26717
R2637 VDD1.n41 VDD1.n40 4.26717
R2638 VDD1.n117 VDD1.n116 4.26717
R2639 VDD1.n133 VDD1.n85 4.26717
R2640 VDD1.n61 VDD1.n60 3.49141
R2641 VDD1.n37 VDD1.n19 3.49141
R2642 VDD1.n113 VDD1.n95 3.49141
R2643 VDD1.n137 VDD1.n136 3.49141
R2644 VDD1.n64 VDD1.n7 2.71565
R2645 VDD1.n36 VDD1.n21 2.71565
R2646 VDD1.n112 VDD1.n97 2.71565
R2647 VDD1.n140 VDD1.n83 2.71565
R2648 VDD1.n65 VDD1.n5 1.93989
R2649 VDD1.n33 VDD1.n32 1.93989
R2650 VDD1.n109 VDD1.n108 1.93989
R2651 VDD1.n141 VDD1.n81 1.93989
R2652 VDD1.n156 VDD1.t2 1.40775
R2653 VDD1.n156 VDD1.t3 1.40775
R2654 VDD1.n154 VDD1.t4 1.40775
R2655 VDD1.n154 VDD1.t0 1.40775
R2656 VDD1.n76 VDD1.n0 1.16414
R2657 VDD1.n69 VDD1.n68 1.16414
R2658 VDD1.n29 VDD1.n23 1.16414
R2659 VDD1.n105 VDD1.n99 1.16414
R2660 VDD1.n146 VDD1.n144 1.16414
R2661 VDD1.n153 VDD1.n77 1.16414
R2662 VDD1 VDD1.n157 0.813
R2663 VDD1.n74 VDD1.n73 0.388379
R2664 VDD1.n4 VDD1.n2 0.388379
R2665 VDD1.n28 VDD1.n25 0.388379
R2666 VDD1.n104 VDD1.n101 0.388379
R2667 VDD1.n145 VDD1.n79 0.388379
R2668 VDD1.n151 VDD1.n150 0.388379
R2669 VDD1.n75 VDD1.n1 0.155672
R2670 VDD1.n67 VDD1.n1 0.155672
R2671 VDD1.n67 VDD1.n66 0.155672
R2672 VDD1.n66 VDD1.n6 0.155672
R2673 VDD1.n59 VDD1.n6 0.155672
R2674 VDD1.n59 VDD1.n58 0.155672
R2675 VDD1.n58 VDD1.n10 0.155672
R2676 VDD1.n51 VDD1.n10 0.155672
R2677 VDD1.n51 VDD1.n50 0.155672
R2678 VDD1.n50 VDD1.n14 0.155672
R2679 VDD1.n43 VDD1.n14 0.155672
R2680 VDD1.n43 VDD1.n42 0.155672
R2681 VDD1.n42 VDD1.n18 0.155672
R2682 VDD1.n35 VDD1.n18 0.155672
R2683 VDD1.n35 VDD1.n34 0.155672
R2684 VDD1.n34 VDD1.n22 0.155672
R2685 VDD1.n27 VDD1.n22 0.155672
R2686 VDD1.n103 VDD1.n98 0.155672
R2687 VDD1.n110 VDD1.n98 0.155672
R2688 VDD1.n111 VDD1.n110 0.155672
R2689 VDD1.n111 VDD1.n94 0.155672
R2690 VDD1.n118 VDD1.n94 0.155672
R2691 VDD1.n119 VDD1.n118 0.155672
R2692 VDD1.n119 VDD1.n90 0.155672
R2693 VDD1.n126 VDD1.n90 0.155672
R2694 VDD1.n127 VDD1.n126 0.155672
R2695 VDD1.n127 VDD1.n86 0.155672
R2696 VDD1.n134 VDD1.n86 0.155672
R2697 VDD1.n135 VDD1.n134 0.155672
R2698 VDD1.n135 VDD1.n82 0.155672
R2699 VDD1.n142 VDD1.n82 0.155672
R2700 VDD1.n143 VDD1.n142 0.155672
R2701 VDD1.n143 VDD1.n78 0.155672
R2702 VDD1.n152 VDD1.n78 0.155672
R2703 VN.n38 VN.n37 161.3
R2704 VN.n36 VN.n21 161.3
R2705 VN.n35 VN.n34 161.3
R2706 VN.n33 VN.n22 161.3
R2707 VN.n32 VN.n31 161.3
R2708 VN.n30 VN.n23 161.3
R2709 VN.n29 VN.n28 161.3
R2710 VN.n27 VN.n24 161.3
R2711 VN.n18 VN.n17 161.3
R2712 VN.n16 VN.n1 161.3
R2713 VN.n15 VN.n14 161.3
R2714 VN.n13 VN.n2 161.3
R2715 VN.n12 VN.n11 161.3
R2716 VN.n10 VN.n3 161.3
R2717 VN.n9 VN.n8 161.3
R2718 VN.n7 VN.n4 161.3
R2719 VN.n26 VN.t3 124.062
R2720 VN.n6 VN.t5 124.062
R2721 VN.n5 VN.t1 91.3986
R2722 VN.n0 VN.t0 91.3986
R2723 VN.n25 VN.t2 91.3986
R2724 VN.n20 VN.t4 91.3986
R2725 VN.n19 VN.n0 88.1101
R2726 VN.n39 VN.n20 88.1101
R2727 VN VN.n39 54.7783
R2728 VN.n6 VN.n5 50.4823
R2729 VN.n26 VN.n25 50.4823
R2730 VN.n11 VN.n2 42.4359
R2731 VN.n31 VN.n22 42.4359
R2732 VN.n11 VN.n10 38.5509
R2733 VN.n31 VN.n30 38.5509
R2734 VN.n5 VN.n4 24.4675
R2735 VN.n9 VN.n4 24.4675
R2736 VN.n10 VN.n9 24.4675
R2737 VN.n15 VN.n2 24.4675
R2738 VN.n16 VN.n15 24.4675
R2739 VN.n17 VN.n16 24.4675
R2740 VN.n30 VN.n29 24.4675
R2741 VN.n29 VN.n24 24.4675
R2742 VN.n25 VN.n24 24.4675
R2743 VN.n37 VN.n36 24.4675
R2744 VN.n36 VN.n35 24.4675
R2745 VN.n35 VN.n22 24.4675
R2746 VN.n7 VN.n6 2.48382
R2747 VN.n27 VN.n26 2.48382
R2748 VN.n17 VN.n0 1.95786
R2749 VN.n37 VN.n20 1.95786
R2750 VN.n39 VN.n38 0.354971
R2751 VN.n19 VN.n18 0.354971
R2752 VN VN.n19 0.26696
R2753 VN.n38 VN.n21 0.189894
R2754 VN.n34 VN.n21 0.189894
R2755 VN.n34 VN.n33 0.189894
R2756 VN.n33 VN.n32 0.189894
R2757 VN.n32 VN.n23 0.189894
R2758 VN.n28 VN.n23 0.189894
R2759 VN.n28 VN.n27 0.189894
R2760 VN.n8 VN.n7 0.189894
R2761 VN.n8 VN.n3 0.189894
R2762 VN.n12 VN.n3 0.189894
R2763 VN.n13 VN.n12 0.189894
R2764 VN.n14 VN.n13 0.189894
R2765 VN.n14 VN.n1 0.189894
R2766 VN.n18 VN.n1 0.189894
R2767 VDD2.n151 VDD2.n79 289.615
R2768 VDD2.n72 VDD2.n0 289.615
R2769 VDD2.n152 VDD2.n151 185
R2770 VDD2.n150 VDD2.n81 185
R2771 VDD2.n149 VDD2.n148 185
R2772 VDD2.n84 VDD2.n82 185
R2773 VDD2.n143 VDD2.n142 185
R2774 VDD2.n141 VDD2.n140 185
R2775 VDD2.n88 VDD2.n87 185
R2776 VDD2.n135 VDD2.n134 185
R2777 VDD2.n133 VDD2.n132 185
R2778 VDD2.n92 VDD2.n91 185
R2779 VDD2.n127 VDD2.n126 185
R2780 VDD2.n125 VDD2.n124 185
R2781 VDD2.n96 VDD2.n95 185
R2782 VDD2.n119 VDD2.n118 185
R2783 VDD2.n117 VDD2.n116 185
R2784 VDD2.n100 VDD2.n99 185
R2785 VDD2.n111 VDD2.n110 185
R2786 VDD2.n109 VDD2.n108 185
R2787 VDD2.n104 VDD2.n103 185
R2788 VDD2.n24 VDD2.n23 185
R2789 VDD2.n29 VDD2.n28 185
R2790 VDD2.n31 VDD2.n30 185
R2791 VDD2.n20 VDD2.n19 185
R2792 VDD2.n37 VDD2.n36 185
R2793 VDD2.n39 VDD2.n38 185
R2794 VDD2.n16 VDD2.n15 185
R2795 VDD2.n45 VDD2.n44 185
R2796 VDD2.n47 VDD2.n46 185
R2797 VDD2.n12 VDD2.n11 185
R2798 VDD2.n53 VDD2.n52 185
R2799 VDD2.n55 VDD2.n54 185
R2800 VDD2.n8 VDD2.n7 185
R2801 VDD2.n61 VDD2.n60 185
R2802 VDD2.n63 VDD2.n62 185
R2803 VDD2.n4 VDD2.n3 185
R2804 VDD2.n70 VDD2.n69 185
R2805 VDD2.n71 VDD2.n2 185
R2806 VDD2.n73 VDD2.n72 185
R2807 VDD2.n105 VDD2.t1 147.659
R2808 VDD2.n25 VDD2.t0 147.659
R2809 VDD2.n151 VDD2.n150 104.615
R2810 VDD2.n150 VDD2.n149 104.615
R2811 VDD2.n149 VDD2.n82 104.615
R2812 VDD2.n142 VDD2.n82 104.615
R2813 VDD2.n142 VDD2.n141 104.615
R2814 VDD2.n141 VDD2.n87 104.615
R2815 VDD2.n134 VDD2.n87 104.615
R2816 VDD2.n134 VDD2.n133 104.615
R2817 VDD2.n133 VDD2.n91 104.615
R2818 VDD2.n126 VDD2.n91 104.615
R2819 VDD2.n126 VDD2.n125 104.615
R2820 VDD2.n125 VDD2.n95 104.615
R2821 VDD2.n118 VDD2.n95 104.615
R2822 VDD2.n118 VDD2.n117 104.615
R2823 VDD2.n117 VDD2.n99 104.615
R2824 VDD2.n110 VDD2.n99 104.615
R2825 VDD2.n110 VDD2.n109 104.615
R2826 VDD2.n109 VDD2.n103 104.615
R2827 VDD2.n29 VDD2.n23 104.615
R2828 VDD2.n30 VDD2.n29 104.615
R2829 VDD2.n30 VDD2.n19 104.615
R2830 VDD2.n37 VDD2.n19 104.615
R2831 VDD2.n38 VDD2.n37 104.615
R2832 VDD2.n38 VDD2.n15 104.615
R2833 VDD2.n45 VDD2.n15 104.615
R2834 VDD2.n46 VDD2.n45 104.615
R2835 VDD2.n46 VDD2.n11 104.615
R2836 VDD2.n53 VDD2.n11 104.615
R2837 VDD2.n54 VDD2.n53 104.615
R2838 VDD2.n54 VDD2.n7 104.615
R2839 VDD2.n61 VDD2.n7 104.615
R2840 VDD2.n62 VDD2.n61 104.615
R2841 VDD2.n62 VDD2.n3 104.615
R2842 VDD2.n70 VDD2.n3 104.615
R2843 VDD2.n71 VDD2.n70 104.615
R2844 VDD2.n72 VDD2.n71 104.615
R2845 VDD2.n78 VDD2.n77 64.7387
R2846 VDD2 VDD2.n157 64.7358
R2847 VDD2.n78 VDD2.n76 54.3299
R2848 VDD2.t1 VDD2.n103 52.3082
R2849 VDD2.t0 VDD2.n23 52.3082
R2850 VDD2.n156 VDD2.n155 51.7732
R2851 VDD2.n156 VDD2.n78 47.1636
R2852 VDD2.n105 VDD2.n104 15.6677
R2853 VDD2.n25 VDD2.n24 15.6677
R2854 VDD2.n152 VDD2.n81 13.1884
R2855 VDD2.n73 VDD2.n2 13.1884
R2856 VDD2.n153 VDD2.n79 12.8005
R2857 VDD2.n148 VDD2.n83 12.8005
R2858 VDD2.n108 VDD2.n107 12.8005
R2859 VDD2.n28 VDD2.n27 12.8005
R2860 VDD2.n69 VDD2.n68 12.8005
R2861 VDD2.n74 VDD2.n0 12.8005
R2862 VDD2.n147 VDD2.n84 12.0247
R2863 VDD2.n111 VDD2.n102 12.0247
R2864 VDD2.n31 VDD2.n22 12.0247
R2865 VDD2.n67 VDD2.n4 12.0247
R2866 VDD2.n144 VDD2.n143 11.249
R2867 VDD2.n112 VDD2.n100 11.249
R2868 VDD2.n32 VDD2.n20 11.249
R2869 VDD2.n64 VDD2.n63 11.249
R2870 VDD2.n140 VDD2.n86 10.4732
R2871 VDD2.n116 VDD2.n115 10.4732
R2872 VDD2.n36 VDD2.n35 10.4732
R2873 VDD2.n60 VDD2.n6 10.4732
R2874 VDD2.n139 VDD2.n88 9.69747
R2875 VDD2.n119 VDD2.n98 9.69747
R2876 VDD2.n39 VDD2.n18 9.69747
R2877 VDD2.n59 VDD2.n8 9.69747
R2878 VDD2.n155 VDD2.n154 9.45567
R2879 VDD2.n76 VDD2.n75 9.45567
R2880 VDD2.n131 VDD2.n130 9.3005
R2881 VDD2.n90 VDD2.n89 9.3005
R2882 VDD2.n137 VDD2.n136 9.3005
R2883 VDD2.n139 VDD2.n138 9.3005
R2884 VDD2.n86 VDD2.n85 9.3005
R2885 VDD2.n145 VDD2.n144 9.3005
R2886 VDD2.n147 VDD2.n146 9.3005
R2887 VDD2.n83 VDD2.n80 9.3005
R2888 VDD2.n154 VDD2.n153 9.3005
R2889 VDD2.n129 VDD2.n128 9.3005
R2890 VDD2.n94 VDD2.n93 9.3005
R2891 VDD2.n123 VDD2.n122 9.3005
R2892 VDD2.n121 VDD2.n120 9.3005
R2893 VDD2.n98 VDD2.n97 9.3005
R2894 VDD2.n115 VDD2.n114 9.3005
R2895 VDD2.n113 VDD2.n112 9.3005
R2896 VDD2.n102 VDD2.n101 9.3005
R2897 VDD2.n107 VDD2.n106 9.3005
R2898 VDD2.n75 VDD2.n74 9.3005
R2899 VDD2.n14 VDD2.n13 9.3005
R2900 VDD2.n43 VDD2.n42 9.3005
R2901 VDD2.n41 VDD2.n40 9.3005
R2902 VDD2.n18 VDD2.n17 9.3005
R2903 VDD2.n35 VDD2.n34 9.3005
R2904 VDD2.n33 VDD2.n32 9.3005
R2905 VDD2.n22 VDD2.n21 9.3005
R2906 VDD2.n27 VDD2.n26 9.3005
R2907 VDD2.n49 VDD2.n48 9.3005
R2908 VDD2.n51 VDD2.n50 9.3005
R2909 VDD2.n10 VDD2.n9 9.3005
R2910 VDD2.n57 VDD2.n56 9.3005
R2911 VDD2.n59 VDD2.n58 9.3005
R2912 VDD2.n6 VDD2.n5 9.3005
R2913 VDD2.n65 VDD2.n64 9.3005
R2914 VDD2.n67 VDD2.n66 9.3005
R2915 VDD2.n68 VDD2.n1 9.3005
R2916 VDD2.n136 VDD2.n135 8.92171
R2917 VDD2.n120 VDD2.n96 8.92171
R2918 VDD2.n40 VDD2.n16 8.92171
R2919 VDD2.n56 VDD2.n55 8.92171
R2920 VDD2.n132 VDD2.n90 8.14595
R2921 VDD2.n124 VDD2.n123 8.14595
R2922 VDD2.n44 VDD2.n43 8.14595
R2923 VDD2.n52 VDD2.n10 8.14595
R2924 VDD2.n131 VDD2.n92 7.3702
R2925 VDD2.n127 VDD2.n94 7.3702
R2926 VDD2.n47 VDD2.n14 7.3702
R2927 VDD2.n51 VDD2.n12 7.3702
R2928 VDD2.n128 VDD2.n92 6.59444
R2929 VDD2.n128 VDD2.n127 6.59444
R2930 VDD2.n48 VDD2.n47 6.59444
R2931 VDD2.n48 VDD2.n12 6.59444
R2932 VDD2.n132 VDD2.n131 5.81868
R2933 VDD2.n124 VDD2.n94 5.81868
R2934 VDD2.n44 VDD2.n14 5.81868
R2935 VDD2.n52 VDD2.n51 5.81868
R2936 VDD2.n135 VDD2.n90 5.04292
R2937 VDD2.n123 VDD2.n96 5.04292
R2938 VDD2.n43 VDD2.n16 5.04292
R2939 VDD2.n55 VDD2.n10 5.04292
R2940 VDD2.n106 VDD2.n105 4.38563
R2941 VDD2.n26 VDD2.n25 4.38563
R2942 VDD2.n136 VDD2.n88 4.26717
R2943 VDD2.n120 VDD2.n119 4.26717
R2944 VDD2.n40 VDD2.n39 4.26717
R2945 VDD2.n56 VDD2.n8 4.26717
R2946 VDD2.n140 VDD2.n139 3.49141
R2947 VDD2.n116 VDD2.n98 3.49141
R2948 VDD2.n36 VDD2.n18 3.49141
R2949 VDD2.n60 VDD2.n59 3.49141
R2950 VDD2.n143 VDD2.n86 2.71565
R2951 VDD2.n115 VDD2.n100 2.71565
R2952 VDD2.n35 VDD2.n20 2.71565
R2953 VDD2.n63 VDD2.n6 2.71565
R2954 VDD2 VDD2.n156 2.67076
R2955 VDD2.n144 VDD2.n84 1.93989
R2956 VDD2.n112 VDD2.n111 1.93989
R2957 VDD2.n32 VDD2.n31 1.93989
R2958 VDD2.n64 VDD2.n4 1.93989
R2959 VDD2.n157 VDD2.t3 1.40775
R2960 VDD2.n157 VDD2.t2 1.40775
R2961 VDD2.n77 VDD2.t4 1.40775
R2962 VDD2.n77 VDD2.t5 1.40775
R2963 VDD2.n155 VDD2.n79 1.16414
R2964 VDD2.n148 VDD2.n147 1.16414
R2965 VDD2.n108 VDD2.n102 1.16414
R2966 VDD2.n28 VDD2.n22 1.16414
R2967 VDD2.n69 VDD2.n67 1.16414
R2968 VDD2.n76 VDD2.n0 1.16414
R2969 VDD2.n153 VDD2.n152 0.388379
R2970 VDD2.n83 VDD2.n81 0.388379
R2971 VDD2.n107 VDD2.n104 0.388379
R2972 VDD2.n27 VDD2.n24 0.388379
R2973 VDD2.n68 VDD2.n2 0.388379
R2974 VDD2.n74 VDD2.n73 0.388379
R2975 VDD2.n154 VDD2.n80 0.155672
R2976 VDD2.n146 VDD2.n80 0.155672
R2977 VDD2.n146 VDD2.n145 0.155672
R2978 VDD2.n145 VDD2.n85 0.155672
R2979 VDD2.n138 VDD2.n85 0.155672
R2980 VDD2.n138 VDD2.n137 0.155672
R2981 VDD2.n137 VDD2.n89 0.155672
R2982 VDD2.n130 VDD2.n89 0.155672
R2983 VDD2.n130 VDD2.n129 0.155672
R2984 VDD2.n129 VDD2.n93 0.155672
R2985 VDD2.n122 VDD2.n93 0.155672
R2986 VDD2.n122 VDD2.n121 0.155672
R2987 VDD2.n121 VDD2.n97 0.155672
R2988 VDD2.n114 VDD2.n97 0.155672
R2989 VDD2.n114 VDD2.n113 0.155672
R2990 VDD2.n113 VDD2.n101 0.155672
R2991 VDD2.n106 VDD2.n101 0.155672
R2992 VDD2.n26 VDD2.n21 0.155672
R2993 VDD2.n33 VDD2.n21 0.155672
R2994 VDD2.n34 VDD2.n33 0.155672
R2995 VDD2.n34 VDD2.n17 0.155672
R2996 VDD2.n41 VDD2.n17 0.155672
R2997 VDD2.n42 VDD2.n41 0.155672
R2998 VDD2.n42 VDD2.n13 0.155672
R2999 VDD2.n49 VDD2.n13 0.155672
R3000 VDD2.n50 VDD2.n49 0.155672
R3001 VDD2.n50 VDD2.n9 0.155672
R3002 VDD2.n57 VDD2.n9 0.155672
R3003 VDD2.n58 VDD2.n57 0.155672
R3004 VDD2.n58 VDD2.n5 0.155672
R3005 VDD2.n65 VDD2.n5 0.155672
R3006 VDD2.n66 VDD2.n65 0.155672
R3007 VDD2.n66 VDD2.n1 0.155672
R3008 VDD2.n75 VDD2.n1 0.155672
C0 VN VDD2 8.28767f
C1 VTAIL VDD2 8.84085f
C2 VP VDD2 0.552044f
C3 VDD1 VDD2 1.83911f
C4 VTAIL VN 8.61509f
C5 VP VN 8.391809f
C6 VDD1 VN 0.152089f
C7 VTAIL VP 8.629701f
C8 VTAIL VDD1 8.782001f
C9 VDD1 VP 8.68468f
C10 VDD2 B 7.18725f
C11 VDD1 B 7.378621f
C12 VTAIL B 9.357997f
C13 VN B 16.316711f
C14 VP B 15.018399f
C15 VDD2.n0 B 0.02854f
C16 VDD2.n1 B 0.021221f
C17 VDD2.n2 B 0.011739f
C18 VDD2.n3 B 0.026953f
C19 VDD2.n4 B 0.012074f
C20 VDD2.n5 B 0.021221f
C21 VDD2.n6 B 0.011403f
C22 VDD2.n7 B 0.026953f
C23 VDD2.n8 B 0.012074f
C24 VDD2.n9 B 0.021221f
C25 VDD2.n10 B 0.011403f
C26 VDD2.n11 B 0.026953f
C27 VDD2.n12 B 0.012074f
C28 VDD2.n13 B 0.021221f
C29 VDD2.n14 B 0.011403f
C30 VDD2.n15 B 0.026953f
C31 VDD2.n16 B 0.012074f
C32 VDD2.n17 B 0.021221f
C33 VDD2.n18 B 0.011403f
C34 VDD2.n19 B 0.026953f
C35 VDD2.n20 B 0.012074f
C36 VDD2.n21 B 0.021221f
C37 VDD2.n22 B 0.011403f
C38 VDD2.n23 B 0.020215f
C39 VDD2.n24 B 0.015922f
C40 VDD2.t0 B 0.044375f
C41 VDD2.n25 B 0.13346f
C42 VDD2.n26 B 1.29023f
C43 VDD2.n27 B 0.011403f
C44 VDD2.n28 B 0.012074f
C45 VDD2.n29 B 0.026953f
C46 VDD2.n30 B 0.026953f
C47 VDD2.n31 B 0.012074f
C48 VDD2.n32 B 0.011403f
C49 VDD2.n33 B 0.021221f
C50 VDD2.n34 B 0.021221f
C51 VDD2.n35 B 0.011403f
C52 VDD2.n36 B 0.012074f
C53 VDD2.n37 B 0.026953f
C54 VDD2.n38 B 0.026953f
C55 VDD2.n39 B 0.012074f
C56 VDD2.n40 B 0.011403f
C57 VDD2.n41 B 0.021221f
C58 VDD2.n42 B 0.021221f
C59 VDD2.n43 B 0.011403f
C60 VDD2.n44 B 0.012074f
C61 VDD2.n45 B 0.026953f
C62 VDD2.n46 B 0.026953f
C63 VDD2.n47 B 0.012074f
C64 VDD2.n48 B 0.011403f
C65 VDD2.n49 B 0.021221f
C66 VDD2.n50 B 0.021221f
C67 VDD2.n51 B 0.011403f
C68 VDD2.n52 B 0.012074f
C69 VDD2.n53 B 0.026953f
C70 VDD2.n54 B 0.026953f
C71 VDD2.n55 B 0.012074f
C72 VDD2.n56 B 0.011403f
C73 VDD2.n57 B 0.021221f
C74 VDD2.n58 B 0.021221f
C75 VDD2.n59 B 0.011403f
C76 VDD2.n60 B 0.012074f
C77 VDD2.n61 B 0.026953f
C78 VDD2.n62 B 0.026953f
C79 VDD2.n63 B 0.012074f
C80 VDD2.n64 B 0.011403f
C81 VDD2.n65 B 0.021221f
C82 VDD2.n66 B 0.021221f
C83 VDD2.n67 B 0.011403f
C84 VDD2.n68 B 0.011403f
C85 VDD2.n69 B 0.012074f
C86 VDD2.n70 B 0.026953f
C87 VDD2.n71 B 0.026953f
C88 VDD2.n72 B 0.05607f
C89 VDD2.n73 B 0.011739f
C90 VDD2.n74 B 0.011403f
C91 VDD2.n75 B 0.0534f
C92 VDD2.n76 B 0.056166f
C93 VDD2.t4 B 0.235948f
C94 VDD2.t5 B 0.235948f
C95 VDD2.n77 B 2.13477f
C96 VDD2.n78 B 2.78745f
C97 VDD2.n79 B 0.02854f
C98 VDD2.n80 B 0.021221f
C99 VDD2.n81 B 0.011739f
C100 VDD2.n82 B 0.026953f
C101 VDD2.n83 B 0.011403f
C102 VDD2.n84 B 0.012074f
C103 VDD2.n85 B 0.021221f
C104 VDD2.n86 B 0.011403f
C105 VDD2.n87 B 0.026953f
C106 VDD2.n88 B 0.012074f
C107 VDD2.n89 B 0.021221f
C108 VDD2.n90 B 0.011403f
C109 VDD2.n91 B 0.026953f
C110 VDD2.n92 B 0.012074f
C111 VDD2.n93 B 0.021221f
C112 VDD2.n94 B 0.011403f
C113 VDD2.n95 B 0.026953f
C114 VDD2.n96 B 0.012074f
C115 VDD2.n97 B 0.021221f
C116 VDD2.n98 B 0.011403f
C117 VDD2.n99 B 0.026953f
C118 VDD2.n100 B 0.012074f
C119 VDD2.n101 B 0.021221f
C120 VDD2.n102 B 0.011403f
C121 VDD2.n103 B 0.020215f
C122 VDD2.n104 B 0.015922f
C123 VDD2.t1 B 0.044375f
C124 VDD2.n105 B 0.13346f
C125 VDD2.n106 B 1.29023f
C126 VDD2.n107 B 0.011403f
C127 VDD2.n108 B 0.012074f
C128 VDD2.n109 B 0.026953f
C129 VDD2.n110 B 0.026953f
C130 VDD2.n111 B 0.012074f
C131 VDD2.n112 B 0.011403f
C132 VDD2.n113 B 0.021221f
C133 VDD2.n114 B 0.021221f
C134 VDD2.n115 B 0.011403f
C135 VDD2.n116 B 0.012074f
C136 VDD2.n117 B 0.026953f
C137 VDD2.n118 B 0.026953f
C138 VDD2.n119 B 0.012074f
C139 VDD2.n120 B 0.011403f
C140 VDD2.n121 B 0.021221f
C141 VDD2.n122 B 0.021221f
C142 VDD2.n123 B 0.011403f
C143 VDD2.n124 B 0.012074f
C144 VDD2.n125 B 0.026953f
C145 VDD2.n126 B 0.026953f
C146 VDD2.n127 B 0.012074f
C147 VDD2.n128 B 0.011403f
C148 VDD2.n129 B 0.021221f
C149 VDD2.n130 B 0.021221f
C150 VDD2.n131 B 0.011403f
C151 VDD2.n132 B 0.012074f
C152 VDD2.n133 B 0.026953f
C153 VDD2.n134 B 0.026953f
C154 VDD2.n135 B 0.012074f
C155 VDD2.n136 B 0.011403f
C156 VDD2.n137 B 0.021221f
C157 VDD2.n138 B 0.021221f
C158 VDD2.n139 B 0.011403f
C159 VDD2.n140 B 0.012074f
C160 VDD2.n141 B 0.026953f
C161 VDD2.n142 B 0.026953f
C162 VDD2.n143 B 0.012074f
C163 VDD2.n144 B 0.011403f
C164 VDD2.n145 B 0.021221f
C165 VDD2.n146 B 0.021221f
C166 VDD2.n147 B 0.011403f
C167 VDD2.n148 B 0.012074f
C168 VDD2.n149 B 0.026953f
C169 VDD2.n150 B 0.026953f
C170 VDD2.n151 B 0.05607f
C171 VDD2.n152 B 0.011739f
C172 VDD2.n153 B 0.011403f
C173 VDD2.n154 B 0.0534f
C174 VDD2.n155 B 0.04589f
C175 VDD2.n156 B 2.56871f
C176 VDD2.t3 B 0.235948f
C177 VDD2.t2 B 0.235948f
C178 VDD2.n157 B 2.13474f
C179 VN.t0 B 2.57553f
C180 VN.n0 B 0.961239f
C181 VN.n1 B 0.018033f
C182 VN.n2 B 0.035435f
C183 VN.n3 B 0.018033f
C184 VN.n4 B 0.033609f
C185 VN.t1 B 2.57553f
C186 VN.n5 B 0.969759f
C187 VN.t5 B 2.84878f
C188 VN.n6 B 0.92157f
C189 VN.n7 B 0.230121f
C190 VN.n8 B 0.018033f
C191 VN.n9 B 0.033609f
C192 VN.n10 B 0.036154f
C193 VN.n11 B 0.014671f
C194 VN.n12 B 0.018033f
C195 VN.n13 B 0.018033f
C196 VN.n14 B 0.018033f
C197 VN.n15 B 0.033609f
C198 VN.n16 B 0.033609f
C199 VN.n17 B 0.018344f
C200 VN.n18 B 0.029105f
C201 VN.n19 B 0.054963f
C202 VN.t4 B 2.57553f
C203 VN.n20 B 0.961239f
C204 VN.n21 B 0.018033f
C205 VN.n22 B 0.035435f
C206 VN.n23 B 0.018033f
C207 VN.n24 B 0.033609f
C208 VN.t3 B 2.84878f
C209 VN.t2 B 2.57553f
C210 VN.n25 B 0.969759f
C211 VN.n26 B 0.92157f
C212 VN.n27 B 0.230121f
C213 VN.n28 B 0.018033f
C214 VN.n29 B 0.033609f
C215 VN.n30 B 0.036154f
C216 VN.n31 B 0.014671f
C217 VN.n32 B 0.018033f
C218 VN.n33 B 0.018033f
C219 VN.n34 B 0.018033f
C220 VN.n35 B 0.033609f
C221 VN.n36 B 0.033609f
C222 VN.n37 B 0.018344f
C223 VN.n38 B 0.029105f
C224 VN.n39 B 1.17969f
C225 VDD1.n0 B 0.029074f
C226 VDD1.n1 B 0.021618f
C227 VDD1.n2 B 0.011958f
C228 VDD1.n3 B 0.027458f
C229 VDD1.n4 B 0.011617f
C230 VDD1.n5 B 0.0123f
C231 VDD1.n6 B 0.021618f
C232 VDD1.n7 B 0.011617f
C233 VDD1.n8 B 0.027458f
C234 VDD1.n9 B 0.0123f
C235 VDD1.n10 B 0.021618f
C236 VDD1.n11 B 0.011617f
C237 VDD1.n12 B 0.027458f
C238 VDD1.n13 B 0.0123f
C239 VDD1.n14 B 0.021618f
C240 VDD1.n15 B 0.011617f
C241 VDD1.n16 B 0.027458f
C242 VDD1.n17 B 0.0123f
C243 VDD1.n18 B 0.021618f
C244 VDD1.n19 B 0.011617f
C245 VDD1.n20 B 0.027458f
C246 VDD1.n21 B 0.0123f
C247 VDD1.n22 B 0.021618f
C248 VDD1.n23 B 0.011617f
C249 VDD1.n24 B 0.020593f
C250 VDD1.n25 B 0.01622f
C251 VDD1.t1 B 0.045206f
C252 VDD1.n26 B 0.135959f
C253 VDD1.n27 B 1.31438f
C254 VDD1.n28 B 0.011617f
C255 VDD1.n29 B 0.0123f
C256 VDD1.n30 B 0.027458f
C257 VDD1.n31 B 0.027458f
C258 VDD1.n32 B 0.0123f
C259 VDD1.n33 B 0.011617f
C260 VDD1.n34 B 0.021618f
C261 VDD1.n35 B 0.021618f
C262 VDD1.n36 B 0.011617f
C263 VDD1.n37 B 0.0123f
C264 VDD1.n38 B 0.027458f
C265 VDD1.n39 B 0.027458f
C266 VDD1.n40 B 0.0123f
C267 VDD1.n41 B 0.011617f
C268 VDD1.n42 B 0.021618f
C269 VDD1.n43 B 0.021618f
C270 VDD1.n44 B 0.011617f
C271 VDD1.n45 B 0.0123f
C272 VDD1.n46 B 0.027458f
C273 VDD1.n47 B 0.027458f
C274 VDD1.n48 B 0.0123f
C275 VDD1.n49 B 0.011617f
C276 VDD1.n50 B 0.021618f
C277 VDD1.n51 B 0.021618f
C278 VDD1.n52 B 0.011617f
C279 VDD1.n53 B 0.0123f
C280 VDD1.n54 B 0.027458f
C281 VDD1.n55 B 0.027458f
C282 VDD1.n56 B 0.0123f
C283 VDD1.n57 B 0.011617f
C284 VDD1.n58 B 0.021618f
C285 VDD1.n59 B 0.021618f
C286 VDD1.n60 B 0.011617f
C287 VDD1.n61 B 0.0123f
C288 VDD1.n62 B 0.027458f
C289 VDD1.n63 B 0.027458f
C290 VDD1.n64 B 0.0123f
C291 VDD1.n65 B 0.011617f
C292 VDD1.n66 B 0.021618f
C293 VDD1.n67 B 0.021618f
C294 VDD1.n68 B 0.011617f
C295 VDD1.n69 B 0.0123f
C296 VDD1.n70 B 0.027458f
C297 VDD1.n71 B 0.027458f
C298 VDD1.n72 B 0.05712f
C299 VDD1.n73 B 0.011958f
C300 VDD1.n74 B 0.011617f
C301 VDD1.n75 B 0.0544f
C302 VDD1.n76 B 0.058038f
C303 VDD1.n77 B 0.029074f
C304 VDD1.n78 B 0.021618f
C305 VDD1.n79 B 0.011958f
C306 VDD1.n80 B 0.027458f
C307 VDD1.n81 B 0.0123f
C308 VDD1.n82 B 0.021618f
C309 VDD1.n83 B 0.011617f
C310 VDD1.n84 B 0.027458f
C311 VDD1.n85 B 0.0123f
C312 VDD1.n86 B 0.021618f
C313 VDD1.n87 B 0.011617f
C314 VDD1.n88 B 0.027458f
C315 VDD1.n89 B 0.0123f
C316 VDD1.n90 B 0.021618f
C317 VDD1.n91 B 0.011617f
C318 VDD1.n92 B 0.027458f
C319 VDD1.n93 B 0.0123f
C320 VDD1.n94 B 0.021618f
C321 VDD1.n95 B 0.011617f
C322 VDD1.n96 B 0.027458f
C323 VDD1.n97 B 0.0123f
C324 VDD1.n98 B 0.021618f
C325 VDD1.n99 B 0.011617f
C326 VDD1.n100 B 0.020593f
C327 VDD1.n101 B 0.01622f
C328 VDD1.t5 B 0.045206f
C329 VDD1.n102 B 0.135959f
C330 VDD1.n103 B 1.31438f
C331 VDD1.n104 B 0.011617f
C332 VDD1.n105 B 0.0123f
C333 VDD1.n106 B 0.027458f
C334 VDD1.n107 B 0.027458f
C335 VDD1.n108 B 0.0123f
C336 VDD1.n109 B 0.011617f
C337 VDD1.n110 B 0.021618f
C338 VDD1.n111 B 0.021618f
C339 VDD1.n112 B 0.011617f
C340 VDD1.n113 B 0.0123f
C341 VDD1.n114 B 0.027458f
C342 VDD1.n115 B 0.027458f
C343 VDD1.n116 B 0.0123f
C344 VDD1.n117 B 0.011617f
C345 VDD1.n118 B 0.021618f
C346 VDD1.n119 B 0.021618f
C347 VDD1.n120 B 0.011617f
C348 VDD1.n121 B 0.0123f
C349 VDD1.n122 B 0.027458f
C350 VDD1.n123 B 0.027458f
C351 VDD1.n124 B 0.0123f
C352 VDD1.n125 B 0.011617f
C353 VDD1.n126 B 0.021618f
C354 VDD1.n127 B 0.021618f
C355 VDD1.n128 B 0.011617f
C356 VDD1.n129 B 0.0123f
C357 VDD1.n130 B 0.027458f
C358 VDD1.n131 B 0.027458f
C359 VDD1.n132 B 0.0123f
C360 VDD1.n133 B 0.011617f
C361 VDD1.n134 B 0.021618f
C362 VDD1.n135 B 0.021618f
C363 VDD1.n136 B 0.011617f
C364 VDD1.n137 B 0.0123f
C365 VDD1.n138 B 0.027458f
C366 VDD1.n139 B 0.027458f
C367 VDD1.n140 B 0.0123f
C368 VDD1.n141 B 0.011617f
C369 VDD1.n142 B 0.021618f
C370 VDD1.n143 B 0.021618f
C371 VDD1.n144 B 0.011617f
C372 VDD1.n145 B 0.011617f
C373 VDD1.n146 B 0.0123f
C374 VDD1.n147 B 0.027458f
C375 VDD1.n148 B 0.027458f
C376 VDD1.n149 B 0.05712f
C377 VDD1.n150 B 0.011958f
C378 VDD1.n151 B 0.011617f
C379 VDD1.n152 B 0.0544f
C380 VDD1.n153 B 0.057218f
C381 VDD1.t4 B 0.240365f
C382 VDD1.t0 B 0.240365f
C383 VDD1.n154 B 2.17474f
C384 VDD1.n155 B 2.97416f
C385 VDD1.t2 B 0.240365f
C386 VDD1.t3 B 0.240365f
C387 VDD1.n156 B 2.16866f
C388 VDD1.n157 B 2.81331f
C389 VTAIL.t2 B 0.264589f
C390 VTAIL.t3 B 0.264589f
C391 VTAIL.n0 B 2.32142f
C392 VTAIL.n1 B 0.465182f
C393 VTAIL.n2 B 0.032004f
C394 VTAIL.n3 B 0.023797f
C395 VTAIL.n4 B 0.013164f
C396 VTAIL.n5 B 0.030225f
C397 VTAIL.n6 B 0.01354f
C398 VTAIL.n7 B 0.023797f
C399 VTAIL.n8 B 0.012788f
C400 VTAIL.n9 B 0.030225f
C401 VTAIL.n10 B 0.01354f
C402 VTAIL.n11 B 0.023797f
C403 VTAIL.n12 B 0.012788f
C404 VTAIL.n13 B 0.030225f
C405 VTAIL.n14 B 0.01354f
C406 VTAIL.n15 B 0.023797f
C407 VTAIL.n16 B 0.012788f
C408 VTAIL.n17 B 0.030225f
C409 VTAIL.n18 B 0.01354f
C410 VTAIL.n19 B 0.023797f
C411 VTAIL.n20 B 0.012788f
C412 VTAIL.n21 B 0.030225f
C413 VTAIL.n22 B 0.01354f
C414 VTAIL.n23 B 0.023797f
C415 VTAIL.n24 B 0.012788f
C416 VTAIL.n25 B 0.022669f
C417 VTAIL.n26 B 0.017855f
C418 VTAIL.t9 B 0.049762f
C419 VTAIL.n27 B 0.149661f
C420 VTAIL.n28 B 1.44685f
C421 VTAIL.n29 B 0.012788f
C422 VTAIL.n30 B 0.01354f
C423 VTAIL.n31 B 0.030225f
C424 VTAIL.n32 B 0.030225f
C425 VTAIL.n33 B 0.01354f
C426 VTAIL.n34 B 0.012788f
C427 VTAIL.n35 B 0.023797f
C428 VTAIL.n36 B 0.023797f
C429 VTAIL.n37 B 0.012788f
C430 VTAIL.n38 B 0.01354f
C431 VTAIL.n39 B 0.030225f
C432 VTAIL.n40 B 0.030225f
C433 VTAIL.n41 B 0.01354f
C434 VTAIL.n42 B 0.012788f
C435 VTAIL.n43 B 0.023797f
C436 VTAIL.n44 B 0.023797f
C437 VTAIL.n45 B 0.012788f
C438 VTAIL.n46 B 0.01354f
C439 VTAIL.n47 B 0.030225f
C440 VTAIL.n48 B 0.030225f
C441 VTAIL.n49 B 0.01354f
C442 VTAIL.n50 B 0.012788f
C443 VTAIL.n51 B 0.023797f
C444 VTAIL.n52 B 0.023797f
C445 VTAIL.n53 B 0.012788f
C446 VTAIL.n54 B 0.01354f
C447 VTAIL.n55 B 0.030225f
C448 VTAIL.n56 B 0.030225f
C449 VTAIL.n57 B 0.01354f
C450 VTAIL.n58 B 0.012788f
C451 VTAIL.n59 B 0.023797f
C452 VTAIL.n60 B 0.023797f
C453 VTAIL.n61 B 0.012788f
C454 VTAIL.n62 B 0.01354f
C455 VTAIL.n63 B 0.030225f
C456 VTAIL.n64 B 0.030225f
C457 VTAIL.n65 B 0.01354f
C458 VTAIL.n66 B 0.012788f
C459 VTAIL.n67 B 0.023797f
C460 VTAIL.n68 B 0.023797f
C461 VTAIL.n69 B 0.012788f
C462 VTAIL.n70 B 0.012788f
C463 VTAIL.n71 B 0.01354f
C464 VTAIL.n72 B 0.030225f
C465 VTAIL.n73 B 0.030225f
C466 VTAIL.n74 B 0.062877f
C467 VTAIL.n75 B 0.013164f
C468 VTAIL.n76 B 0.012788f
C469 VTAIL.n77 B 0.059882f
C470 VTAIL.n78 B 0.035064f
C471 VTAIL.n79 B 0.459694f
C472 VTAIL.t5 B 0.264589f
C473 VTAIL.t6 B 0.264589f
C474 VTAIL.n80 B 2.32142f
C475 VTAIL.n81 B 2.2789f
C476 VTAIL.t1 B 0.264589f
C477 VTAIL.t4 B 0.264589f
C478 VTAIL.n82 B 2.32143f
C479 VTAIL.n83 B 2.27889f
C480 VTAIL.n84 B 0.032004f
C481 VTAIL.n85 B 0.023797f
C482 VTAIL.n86 B 0.013164f
C483 VTAIL.n87 B 0.030225f
C484 VTAIL.n88 B 0.012788f
C485 VTAIL.n89 B 0.01354f
C486 VTAIL.n90 B 0.023797f
C487 VTAIL.n91 B 0.012788f
C488 VTAIL.n92 B 0.030225f
C489 VTAIL.n93 B 0.01354f
C490 VTAIL.n94 B 0.023797f
C491 VTAIL.n95 B 0.012788f
C492 VTAIL.n96 B 0.030225f
C493 VTAIL.n97 B 0.01354f
C494 VTAIL.n98 B 0.023797f
C495 VTAIL.n99 B 0.012788f
C496 VTAIL.n100 B 0.030225f
C497 VTAIL.n101 B 0.01354f
C498 VTAIL.n102 B 0.023797f
C499 VTAIL.n103 B 0.012788f
C500 VTAIL.n104 B 0.030225f
C501 VTAIL.n105 B 0.01354f
C502 VTAIL.n106 B 0.023797f
C503 VTAIL.n107 B 0.012788f
C504 VTAIL.n108 B 0.022669f
C505 VTAIL.n109 B 0.017855f
C506 VTAIL.t11 B 0.049762f
C507 VTAIL.n110 B 0.149661f
C508 VTAIL.n111 B 1.44685f
C509 VTAIL.n112 B 0.012788f
C510 VTAIL.n113 B 0.01354f
C511 VTAIL.n114 B 0.030225f
C512 VTAIL.n115 B 0.030225f
C513 VTAIL.n116 B 0.01354f
C514 VTAIL.n117 B 0.012788f
C515 VTAIL.n118 B 0.023797f
C516 VTAIL.n119 B 0.023797f
C517 VTAIL.n120 B 0.012788f
C518 VTAIL.n121 B 0.01354f
C519 VTAIL.n122 B 0.030225f
C520 VTAIL.n123 B 0.030225f
C521 VTAIL.n124 B 0.01354f
C522 VTAIL.n125 B 0.012788f
C523 VTAIL.n126 B 0.023797f
C524 VTAIL.n127 B 0.023797f
C525 VTAIL.n128 B 0.012788f
C526 VTAIL.n129 B 0.01354f
C527 VTAIL.n130 B 0.030225f
C528 VTAIL.n131 B 0.030225f
C529 VTAIL.n132 B 0.01354f
C530 VTAIL.n133 B 0.012788f
C531 VTAIL.n134 B 0.023797f
C532 VTAIL.n135 B 0.023797f
C533 VTAIL.n136 B 0.012788f
C534 VTAIL.n137 B 0.01354f
C535 VTAIL.n138 B 0.030225f
C536 VTAIL.n139 B 0.030225f
C537 VTAIL.n140 B 0.01354f
C538 VTAIL.n141 B 0.012788f
C539 VTAIL.n142 B 0.023797f
C540 VTAIL.n143 B 0.023797f
C541 VTAIL.n144 B 0.012788f
C542 VTAIL.n145 B 0.01354f
C543 VTAIL.n146 B 0.030225f
C544 VTAIL.n147 B 0.030225f
C545 VTAIL.n148 B 0.01354f
C546 VTAIL.n149 B 0.012788f
C547 VTAIL.n150 B 0.023797f
C548 VTAIL.n151 B 0.023797f
C549 VTAIL.n152 B 0.012788f
C550 VTAIL.n153 B 0.01354f
C551 VTAIL.n154 B 0.030225f
C552 VTAIL.n155 B 0.030225f
C553 VTAIL.n156 B 0.062877f
C554 VTAIL.n157 B 0.013164f
C555 VTAIL.n158 B 0.012788f
C556 VTAIL.n159 B 0.059882f
C557 VTAIL.n160 B 0.035064f
C558 VTAIL.n161 B 0.459694f
C559 VTAIL.t10 B 0.264589f
C560 VTAIL.t8 B 0.264589f
C561 VTAIL.n162 B 2.32143f
C562 VTAIL.n163 B 0.661002f
C563 VTAIL.n164 B 0.032004f
C564 VTAIL.n165 B 0.023797f
C565 VTAIL.n166 B 0.013164f
C566 VTAIL.n167 B 0.030225f
C567 VTAIL.n168 B 0.012788f
C568 VTAIL.n169 B 0.01354f
C569 VTAIL.n170 B 0.023797f
C570 VTAIL.n171 B 0.012788f
C571 VTAIL.n172 B 0.030225f
C572 VTAIL.n173 B 0.01354f
C573 VTAIL.n174 B 0.023797f
C574 VTAIL.n175 B 0.012788f
C575 VTAIL.n176 B 0.030225f
C576 VTAIL.n177 B 0.01354f
C577 VTAIL.n178 B 0.023797f
C578 VTAIL.n179 B 0.012788f
C579 VTAIL.n180 B 0.030225f
C580 VTAIL.n181 B 0.01354f
C581 VTAIL.n182 B 0.023797f
C582 VTAIL.n183 B 0.012788f
C583 VTAIL.n184 B 0.030225f
C584 VTAIL.n185 B 0.01354f
C585 VTAIL.n186 B 0.023797f
C586 VTAIL.n187 B 0.012788f
C587 VTAIL.n188 B 0.022669f
C588 VTAIL.n189 B 0.017855f
C589 VTAIL.t7 B 0.049762f
C590 VTAIL.n190 B 0.149661f
C591 VTAIL.n191 B 1.44685f
C592 VTAIL.n192 B 0.012788f
C593 VTAIL.n193 B 0.01354f
C594 VTAIL.n194 B 0.030225f
C595 VTAIL.n195 B 0.030225f
C596 VTAIL.n196 B 0.01354f
C597 VTAIL.n197 B 0.012788f
C598 VTAIL.n198 B 0.023797f
C599 VTAIL.n199 B 0.023797f
C600 VTAIL.n200 B 0.012788f
C601 VTAIL.n201 B 0.01354f
C602 VTAIL.n202 B 0.030225f
C603 VTAIL.n203 B 0.030225f
C604 VTAIL.n204 B 0.01354f
C605 VTAIL.n205 B 0.012788f
C606 VTAIL.n206 B 0.023797f
C607 VTAIL.n207 B 0.023797f
C608 VTAIL.n208 B 0.012788f
C609 VTAIL.n209 B 0.01354f
C610 VTAIL.n210 B 0.030225f
C611 VTAIL.n211 B 0.030225f
C612 VTAIL.n212 B 0.01354f
C613 VTAIL.n213 B 0.012788f
C614 VTAIL.n214 B 0.023797f
C615 VTAIL.n215 B 0.023797f
C616 VTAIL.n216 B 0.012788f
C617 VTAIL.n217 B 0.01354f
C618 VTAIL.n218 B 0.030225f
C619 VTAIL.n219 B 0.030225f
C620 VTAIL.n220 B 0.01354f
C621 VTAIL.n221 B 0.012788f
C622 VTAIL.n222 B 0.023797f
C623 VTAIL.n223 B 0.023797f
C624 VTAIL.n224 B 0.012788f
C625 VTAIL.n225 B 0.01354f
C626 VTAIL.n226 B 0.030225f
C627 VTAIL.n227 B 0.030225f
C628 VTAIL.n228 B 0.01354f
C629 VTAIL.n229 B 0.012788f
C630 VTAIL.n230 B 0.023797f
C631 VTAIL.n231 B 0.023797f
C632 VTAIL.n232 B 0.012788f
C633 VTAIL.n233 B 0.01354f
C634 VTAIL.n234 B 0.030225f
C635 VTAIL.n235 B 0.030225f
C636 VTAIL.n236 B 0.062877f
C637 VTAIL.n237 B 0.013164f
C638 VTAIL.n238 B 0.012788f
C639 VTAIL.n239 B 0.059882f
C640 VTAIL.n240 B 0.035064f
C641 VTAIL.n241 B 1.81052f
C642 VTAIL.n242 B 0.032004f
C643 VTAIL.n243 B 0.023797f
C644 VTAIL.n244 B 0.013164f
C645 VTAIL.n245 B 0.030225f
C646 VTAIL.n246 B 0.01354f
C647 VTAIL.n247 B 0.023797f
C648 VTAIL.n248 B 0.012788f
C649 VTAIL.n249 B 0.030225f
C650 VTAIL.n250 B 0.01354f
C651 VTAIL.n251 B 0.023797f
C652 VTAIL.n252 B 0.012788f
C653 VTAIL.n253 B 0.030225f
C654 VTAIL.n254 B 0.01354f
C655 VTAIL.n255 B 0.023797f
C656 VTAIL.n256 B 0.012788f
C657 VTAIL.n257 B 0.030225f
C658 VTAIL.n258 B 0.01354f
C659 VTAIL.n259 B 0.023797f
C660 VTAIL.n260 B 0.012788f
C661 VTAIL.n261 B 0.030225f
C662 VTAIL.n262 B 0.01354f
C663 VTAIL.n263 B 0.023797f
C664 VTAIL.n264 B 0.012788f
C665 VTAIL.n265 B 0.022669f
C666 VTAIL.n266 B 0.017855f
C667 VTAIL.t0 B 0.049762f
C668 VTAIL.n267 B 0.149661f
C669 VTAIL.n268 B 1.44685f
C670 VTAIL.n269 B 0.012788f
C671 VTAIL.n270 B 0.01354f
C672 VTAIL.n271 B 0.030225f
C673 VTAIL.n272 B 0.030225f
C674 VTAIL.n273 B 0.01354f
C675 VTAIL.n274 B 0.012788f
C676 VTAIL.n275 B 0.023797f
C677 VTAIL.n276 B 0.023797f
C678 VTAIL.n277 B 0.012788f
C679 VTAIL.n278 B 0.01354f
C680 VTAIL.n279 B 0.030225f
C681 VTAIL.n280 B 0.030225f
C682 VTAIL.n281 B 0.01354f
C683 VTAIL.n282 B 0.012788f
C684 VTAIL.n283 B 0.023797f
C685 VTAIL.n284 B 0.023797f
C686 VTAIL.n285 B 0.012788f
C687 VTAIL.n286 B 0.01354f
C688 VTAIL.n287 B 0.030225f
C689 VTAIL.n288 B 0.030225f
C690 VTAIL.n289 B 0.01354f
C691 VTAIL.n290 B 0.012788f
C692 VTAIL.n291 B 0.023797f
C693 VTAIL.n292 B 0.023797f
C694 VTAIL.n293 B 0.012788f
C695 VTAIL.n294 B 0.01354f
C696 VTAIL.n295 B 0.030225f
C697 VTAIL.n296 B 0.030225f
C698 VTAIL.n297 B 0.01354f
C699 VTAIL.n298 B 0.012788f
C700 VTAIL.n299 B 0.023797f
C701 VTAIL.n300 B 0.023797f
C702 VTAIL.n301 B 0.012788f
C703 VTAIL.n302 B 0.01354f
C704 VTAIL.n303 B 0.030225f
C705 VTAIL.n304 B 0.030225f
C706 VTAIL.n305 B 0.01354f
C707 VTAIL.n306 B 0.012788f
C708 VTAIL.n307 B 0.023797f
C709 VTAIL.n308 B 0.023797f
C710 VTAIL.n309 B 0.012788f
C711 VTAIL.n310 B 0.012788f
C712 VTAIL.n311 B 0.01354f
C713 VTAIL.n312 B 0.030225f
C714 VTAIL.n313 B 0.030225f
C715 VTAIL.n314 B 0.062877f
C716 VTAIL.n315 B 0.013164f
C717 VTAIL.n316 B 0.012788f
C718 VTAIL.n317 B 0.059882f
C719 VTAIL.n318 B 0.035064f
C720 VTAIL.n319 B 1.7393f
C721 VP.t5 B 2.61887f
C722 VP.n0 B 0.977416f
C723 VP.n1 B 0.018337f
C724 VP.n2 B 0.036031f
C725 VP.n3 B 0.018337f
C726 VP.n4 B 0.034175f
C727 VP.n5 B 0.018337f
C728 VP.t1 B 2.61887f
C729 VP.n6 B 0.036762f
C730 VP.n7 B 0.018337f
C731 VP.n8 B 0.034175f
C732 VP.t2 B 2.61887f
C733 VP.n9 B 0.977416f
C734 VP.n10 B 0.018337f
C735 VP.n11 B 0.036031f
C736 VP.n12 B 0.018337f
C737 VP.n13 B 0.034175f
C738 VP.t4 B 2.89672f
C739 VP.t3 B 2.61887f
C740 VP.n14 B 0.986079f
C741 VP.n15 B 0.93708f
C742 VP.n16 B 0.233994f
C743 VP.n17 B 0.018337f
C744 VP.n18 B 0.034175f
C745 VP.n19 B 0.036762f
C746 VP.n20 B 0.014918f
C747 VP.n21 B 0.018337f
C748 VP.n22 B 0.018337f
C749 VP.n23 B 0.018337f
C750 VP.n24 B 0.034175f
C751 VP.n25 B 0.034175f
C752 VP.n26 B 0.018652f
C753 VP.n27 B 0.029595f
C754 VP.n28 B 1.19225f
C755 VP.n29 B 1.20432f
C756 VP.t0 B 2.61887f
C757 VP.n30 B 0.977416f
C758 VP.n31 B 0.018652f
C759 VP.n32 B 0.029595f
C760 VP.n33 B 0.018337f
C761 VP.n34 B 0.018337f
C762 VP.n35 B 0.034175f
C763 VP.n36 B 0.036031f
C764 VP.n37 B 0.014918f
C765 VP.n38 B 0.018337f
C766 VP.n39 B 0.018337f
C767 VP.n40 B 0.018337f
C768 VP.n41 B 0.034175f
C769 VP.n42 B 0.034175f
C770 VP.n43 B 0.928315f
C771 VP.n44 B 0.018337f
C772 VP.n45 B 0.018337f
C773 VP.n46 B 0.018337f
C774 VP.n47 B 0.034175f
C775 VP.n48 B 0.036762f
C776 VP.n49 B 0.014918f
C777 VP.n50 B 0.018337f
C778 VP.n51 B 0.018337f
C779 VP.n52 B 0.018337f
C780 VP.n53 B 0.034175f
C781 VP.n54 B 0.034175f
C782 VP.n55 B 0.018652f
C783 VP.n56 B 0.029595f
C784 VP.n57 B 0.055888f
.ends

