* NGSPICE file created from diff_pair_sample_0083.ext - technology: sky130A

.subckt diff_pair_sample_0083 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2512_n2740# sky130_fd_pr__pfet_01v8 ad=3.4554 pd=18.5 as=0 ps=0 w=8.86 l=2.24
X1 VDD1.t3 VP.t0 VTAIL.t7 w_n2512_n2740# sky130_fd_pr__pfet_01v8 ad=1.4619 pd=9.19 as=3.4554 ps=18.5 w=8.86 l=2.24
X2 B.t8 B.t6 B.t7 w_n2512_n2740# sky130_fd_pr__pfet_01v8 ad=3.4554 pd=18.5 as=0 ps=0 w=8.86 l=2.24
X3 VTAIL.t6 VP.t1 VDD1.t2 w_n2512_n2740# sky130_fd_pr__pfet_01v8 ad=3.4554 pd=18.5 as=1.4619 ps=9.19 w=8.86 l=2.24
X4 VTAIL.t3 VN.t0 VDD2.t3 w_n2512_n2740# sky130_fd_pr__pfet_01v8 ad=3.4554 pd=18.5 as=1.4619 ps=9.19 w=8.86 l=2.24
X5 VDD2.t2 VN.t1 VTAIL.t0 w_n2512_n2740# sky130_fd_pr__pfet_01v8 ad=1.4619 pd=9.19 as=3.4554 ps=18.5 w=8.86 l=2.24
X6 VTAIL.t5 VP.t2 VDD1.t1 w_n2512_n2740# sky130_fd_pr__pfet_01v8 ad=3.4554 pd=18.5 as=1.4619 ps=9.19 w=8.86 l=2.24
X7 VDD1.t0 VP.t3 VTAIL.t4 w_n2512_n2740# sky130_fd_pr__pfet_01v8 ad=1.4619 pd=9.19 as=3.4554 ps=18.5 w=8.86 l=2.24
X8 VTAIL.t1 VN.t2 VDD2.t1 w_n2512_n2740# sky130_fd_pr__pfet_01v8 ad=3.4554 pd=18.5 as=1.4619 ps=9.19 w=8.86 l=2.24
X9 VDD2.t0 VN.t3 VTAIL.t2 w_n2512_n2740# sky130_fd_pr__pfet_01v8 ad=1.4619 pd=9.19 as=3.4554 ps=18.5 w=8.86 l=2.24
X10 B.t5 B.t3 B.t4 w_n2512_n2740# sky130_fd_pr__pfet_01v8 ad=3.4554 pd=18.5 as=0 ps=0 w=8.86 l=2.24
X11 B.t2 B.t0 B.t1 w_n2512_n2740# sky130_fd_pr__pfet_01v8 ad=3.4554 pd=18.5 as=0 ps=0 w=8.86 l=2.24
R0 B.n400 B.n59 585
R1 B.n402 B.n401 585
R2 B.n403 B.n58 585
R3 B.n405 B.n404 585
R4 B.n406 B.n57 585
R5 B.n408 B.n407 585
R6 B.n409 B.n56 585
R7 B.n411 B.n410 585
R8 B.n412 B.n55 585
R9 B.n414 B.n413 585
R10 B.n415 B.n54 585
R11 B.n417 B.n416 585
R12 B.n418 B.n53 585
R13 B.n420 B.n419 585
R14 B.n421 B.n52 585
R15 B.n423 B.n422 585
R16 B.n424 B.n51 585
R17 B.n426 B.n425 585
R18 B.n427 B.n50 585
R19 B.n429 B.n428 585
R20 B.n430 B.n49 585
R21 B.n432 B.n431 585
R22 B.n433 B.n48 585
R23 B.n435 B.n434 585
R24 B.n436 B.n47 585
R25 B.n438 B.n437 585
R26 B.n439 B.n46 585
R27 B.n441 B.n440 585
R28 B.n442 B.n45 585
R29 B.n444 B.n443 585
R30 B.n445 B.n41 585
R31 B.n447 B.n446 585
R32 B.n448 B.n40 585
R33 B.n450 B.n449 585
R34 B.n451 B.n39 585
R35 B.n453 B.n452 585
R36 B.n454 B.n38 585
R37 B.n456 B.n455 585
R38 B.n457 B.n37 585
R39 B.n459 B.n458 585
R40 B.n460 B.n36 585
R41 B.n462 B.n461 585
R42 B.n464 B.n33 585
R43 B.n466 B.n465 585
R44 B.n467 B.n32 585
R45 B.n469 B.n468 585
R46 B.n470 B.n31 585
R47 B.n472 B.n471 585
R48 B.n473 B.n30 585
R49 B.n475 B.n474 585
R50 B.n476 B.n29 585
R51 B.n478 B.n477 585
R52 B.n479 B.n28 585
R53 B.n481 B.n480 585
R54 B.n482 B.n27 585
R55 B.n484 B.n483 585
R56 B.n485 B.n26 585
R57 B.n487 B.n486 585
R58 B.n488 B.n25 585
R59 B.n490 B.n489 585
R60 B.n491 B.n24 585
R61 B.n493 B.n492 585
R62 B.n494 B.n23 585
R63 B.n496 B.n495 585
R64 B.n497 B.n22 585
R65 B.n499 B.n498 585
R66 B.n500 B.n21 585
R67 B.n502 B.n501 585
R68 B.n503 B.n20 585
R69 B.n505 B.n504 585
R70 B.n506 B.n19 585
R71 B.n508 B.n507 585
R72 B.n509 B.n18 585
R73 B.n511 B.n510 585
R74 B.n399 B.n398 585
R75 B.n397 B.n60 585
R76 B.n396 B.n395 585
R77 B.n394 B.n61 585
R78 B.n393 B.n392 585
R79 B.n391 B.n62 585
R80 B.n390 B.n389 585
R81 B.n388 B.n63 585
R82 B.n387 B.n386 585
R83 B.n385 B.n64 585
R84 B.n384 B.n383 585
R85 B.n382 B.n65 585
R86 B.n381 B.n380 585
R87 B.n379 B.n66 585
R88 B.n378 B.n377 585
R89 B.n376 B.n67 585
R90 B.n375 B.n374 585
R91 B.n373 B.n68 585
R92 B.n372 B.n371 585
R93 B.n370 B.n69 585
R94 B.n369 B.n368 585
R95 B.n367 B.n70 585
R96 B.n366 B.n365 585
R97 B.n364 B.n71 585
R98 B.n363 B.n362 585
R99 B.n361 B.n72 585
R100 B.n360 B.n359 585
R101 B.n358 B.n73 585
R102 B.n357 B.n356 585
R103 B.n355 B.n74 585
R104 B.n354 B.n353 585
R105 B.n352 B.n75 585
R106 B.n351 B.n350 585
R107 B.n349 B.n76 585
R108 B.n348 B.n347 585
R109 B.n346 B.n77 585
R110 B.n345 B.n344 585
R111 B.n343 B.n78 585
R112 B.n342 B.n341 585
R113 B.n340 B.n79 585
R114 B.n339 B.n338 585
R115 B.n337 B.n80 585
R116 B.n336 B.n335 585
R117 B.n334 B.n81 585
R118 B.n333 B.n332 585
R119 B.n331 B.n82 585
R120 B.n330 B.n329 585
R121 B.n328 B.n83 585
R122 B.n327 B.n326 585
R123 B.n325 B.n84 585
R124 B.n324 B.n323 585
R125 B.n322 B.n85 585
R126 B.n321 B.n320 585
R127 B.n319 B.n86 585
R128 B.n318 B.n317 585
R129 B.n316 B.n87 585
R130 B.n315 B.n314 585
R131 B.n313 B.n88 585
R132 B.n312 B.n311 585
R133 B.n310 B.n89 585
R134 B.n309 B.n308 585
R135 B.n307 B.n90 585
R136 B.n306 B.n305 585
R137 B.n193 B.n132 585
R138 B.n195 B.n194 585
R139 B.n196 B.n131 585
R140 B.n198 B.n197 585
R141 B.n199 B.n130 585
R142 B.n201 B.n200 585
R143 B.n202 B.n129 585
R144 B.n204 B.n203 585
R145 B.n205 B.n128 585
R146 B.n207 B.n206 585
R147 B.n208 B.n127 585
R148 B.n210 B.n209 585
R149 B.n211 B.n126 585
R150 B.n213 B.n212 585
R151 B.n214 B.n125 585
R152 B.n216 B.n215 585
R153 B.n217 B.n124 585
R154 B.n219 B.n218 585
R155 B.n220 B.n123 585
R156 B.n222 B.n221 585
R157 B.n223 B.n122 585
R158 B.n225 B.n224 585
R159 B.n226 B.n121 585
R160 B.n228 B.n227 585
R161 B.n229 B.n120 585
R162 B.n231 B.n230 585
R163 B.n232 B.n119 585
R164 B.n234 B.n233 585
R165 B.n235 B.n118 585
R166 B.n237 B.n236 585
R167 B.n238 B.n117 585
R168 B.n240 B.n239 585
R169 B.n242 B.n114 585
R170 B.n244 B.n243 585
R171 B.n245 B.n113 585
R172 B.n247 B.n246 585
R173 B.n248 B.n112 585
R174 B.n250 B.n249 585
R175 B.n251 B.n111 585
R176 B.n253 B.n252 585
R177 B.n254 B.n110 585
R178 B.n256 B.n255 585
R179 B.n258 B.n257 585
R180 B.n259 B.n106 585
R181 B.n261 B.n260 585
R182 B.n262 B.n105 585
R183 B.n264 B.n263 585
R184 B.n265 B.n104 585
R185 B.n267 B.n266 585
R186 B.n268 B.n103 585
R187 B.n270 B.n269 585
R188 B.n271 B.n102 585
R189 B.n273 B.n272 585
R190 B.n274 B.n101 585
R191 B.n276 B.n275 585
R192 B.n277 B.n100 585
R193 B.n279 B.n278 585
R194 B.n280 B.n99 585
R195 B.n282 B.n281 585
R196 B.n283 B.n98 585
R197 B.n285 B.n284 585
R198 B.n286 B.n97 585
R199 B.n288 B.n287 585
R200 B.n289 B.n96 585
R201 B.n291 B.n290 585
R202 B.n292 B.n95 585
R203 B.n294 B.n293 585
R204 B.n295 B.n94 585
R205 B.n297 B.n296 585
R206 B.n298 B.n93 585
R207 B.n300 B.n299 585
R208 B.n301 B.n92 585
R209 B.n303 B.n302 585
R210 B.n304 B.n91 585
R211 B.n192 B.n191 585
R212 B.n190 B.n133 585
R213 B.n189 B.n188 585
R214 B.n187 B.n134 585
R215 B.n186 B.n185 585
R216 B.n184 B.n135 585
R217 B.n183 B.n182 585
R218 B.n181 B.n136 585
R219 B.n180 B.n179 585
R220 B.n178 B.n137 585
R221 B.n177 B.n176 585
R222 B.n175 B.n138 585
R223 B.n174 B.n173 585
R224 B.n172 B.n139 585
R225 B.n171 B.n170 585
R226 B.n169 B.n140 585
R227 B.n168 B.n167 585
R228 B.n166 B.n141 585
R229 B.n165 B.n164 585
R230 B.n163 B.n142 585
R231 B.n162 B.n161 585
R232 B.n160 B.n143 585
R233 B.n159 B.n158 585
R234 B.n157 B.n144 585
R235 B.n156 B.n155 585
R236 B.n154 B.n145 585
R237 B.n153 B.n152 585
R238 B.n151 B.n146 585
R239 B.n150 B.n149 585
R240 B.n148 B.n147 585
R241 B.n2 B.n0 585
R242 B.n557 B.n1 585
R243 B.n556 B.n555 585
R244 B.n554 B.n3 585
R245 B.n553 B.n552 585
R246 B.n551 B.n4 585
R247 B.n550 B.n549 585
R248 B.n548 B.n5 585
R249 B.n547 B.n546 585
R250 B.n545 B.n6 585
R251 B.n544 B.n543 585
R252 B.n542 B.n7 585
R253 B.n541 B.n540 585
R254 B.n539 B.n8 585
R255 B.n538 B.n537 585
R256 B.n536 B.n9 585
R257 B.n535 B.n534 585
R258 B.n533 B.n10 585
R259 B.n532 B.n531 585
R260 B.n530 B.n11 585
R261 B.n529 B.n528 585
R262 B.n527 B.n12 585
R263 B.n526 B.n525 585
R264 B.n524 B.n13 585
R265 B.n523 B.n522 585
R266 B.n521 B.n14 585
R267 B.n520 B.n519 585
R268 B.n518 B.n15 585
R269 B.n517 B.n516 585
R270 B.n515 B.n16 585
R271 B.n514 B.n513 585
R272 B.n512 B.n17 585
R273 B.n559 B.n558 585
R274 B.n191 B.n132 492.5
R275 B.n510 B.n17 492.5
R276 B.n305 B.n304 492.5
R277 B.n400 B.n399 492.5
R278 B.n107 B.t9 302.755
R279 B.n115 B.t0 302.755
R280 B.n34 B.t6 302.755
R281 B.n42 B.t3 302.755
R282 B.n191 B.n190 163.367
R283 B.n190 B.n189 163.367
R284 B.n189 B.n134 163.367
R285 B.n185 B.n134 163.367
R286 B.n185 B.n184 163.367
R287 B.n184 B.n183 163.367
R288 B.n183 B.n136 163.367
R289 B.n179 B.n136 163.367
R290 B.n179 B.n178 163.367
R291 B.n178 B.n177 163.367
R292 B.n177 B.n138 163.367
R293 B.n173 B.n138 163.367
R294 B.n173 B.n172 163.367
R295 B.n172 B.n171 163.367
R296 B.n171 B.n140 163.367
R297 B.n167 B.n140 163.367
R298 B.n167 B.n166 163.367
R299 B.n166 B.n165 163.367
R300 B.n165 B.n142 163.367
R301 B.n161 B.n142 163.367
R302 B.n161 B.n160 163.367
R303 B.n160 B.n159 163.367
R304 B.n159 B.n144 163.367
R305 B.n155 B.n144 163.367
R306 B.n155 B.n154 163.367
R307 B.n154 B.n153 163.367
R308 B.n153 B.n146 163.367
R309 B.n149 B.n146 163.367
R310 B.n149 B.n148 163.367
R311 B.n148 B.n2 163.367
R312 B.n558 B.n2 163.367
R313 B.n558 B.n557 163.367
R314 B.n557 B.n556 163.367
R315 B.n556 B.n3 163.367
R316 B.n552 B.n3 163.367
R317 B.n552 B.n551 163.367
R318 B.n551 B.n550 163.367
R319 B.n550 B.n5 163.367
R320 B.n546 B.n5 163.367
R321 B.n546 B.n545 163.367
R322 B.n545 B.n544 163.367
R323 B.n544 B.n7 163.367
R324 B.n540 B.n7 163.367
R325 B.n540 B.n539 163.367
R326 B.n539 B.n538 163.367
R327 B.n538 B.n9 163.367
R328 B.n534 B.n9 163.367
R329 B.n534 B.n533 163.367
R330 B.n533 B.n532 163.367
R331 B.n532 B.n11 163.367
R332 B.n528 B.n11 163.367
R333 B.n528 B.n527 163.367
R334 B.n527 B.n526 163.367
R335 B.n526 B.n13 163.367
R336 B.n522 B.n13 163.367
R337 B.n522 B.n521 163.367
R338 B.n521 B.n520 163.367
R339 B.n520 B.n15 163.367
R340 B.n516 B.n15 163.367
R341 B.n516 B.n515 163.367
R342 B.n515 B.n514 163.367
R343 B.n514 B.n17 163.367
R344 B.n195 B.n132 163.367
R345 B.n196 B.n195 163.367
R346 B.n197 B.n196 163.367
R347 B.n197 B.n130 163.367
R348 B.n201 B.n130 163.367
R349 B.n202 B.n201 163.367
R350 B.n203 B.n202 163.367
R351 B.n203 B.n128 163.367
R352 B.n207 B.n128 163.367
R353 B.n208 B.n207 163.367
R354 B.n209 B.n208 163.367
R355 B.n209 B.n126 163.367
R356 B.n213 B.n126 163.367
R357 B.n214 B.n213 163.367
R358 B.n215 B.n214 163.367
R359 B.n215 B.n124 163.367
R360 B.n219 B.n124 163.367
R361 B.n220 B.n219 163.367
R362 B.n221 B.n220 163.367
R363 B.n221 B.n122 163.367
R364 B.n225 B.n122 163.367
R365 B.n226 B.n225 163.367
R366 B.n227 B.n226 163.367
R367 B.n227 B.n120 163.367
R368 B.n231 B.n120 163.367
R369 B.n232 B.n231 163.367
R370 B.n233 B.n232 163.367
R371 B.n233 B.n118 163.367
R372 B.n237 B.n118 163.367
R373 B.n238 B.n237 163.367
R374 B.n239 B.n238 163.367
R375 B.n239 B.n114 163.367
R376 B.n244 B.n114 163.367
R377 B.n245 B.n244 163.367
R378 B.n246 B.n245 163.367
R379 B.n246 B.n112 163.367
R380 B.n250 B.n112 163.367
R381 B.n251 B.n250 163.367
R382 B.n252 B.n251 163.367
R383 B.n252 B.n110 163.367
R384 B.n256 B.n110 163.367
R385 B.n257 B.n256 163.367
R386 B.n257 B.n106 163.367
R387 B.n261 B.n106 163.367
R388 B.n262 B.n261 163.367
R389 B.n263 B.n262 163.367
R390 B.n263 B.n104 163.367
R391 B.n267 B.n104 163.367
R392 B.n268 B.n267 163.367
R393 B.n269 B.n268 163.367
R394 B.n269 B.n102 163.367
R395 B.n273 B.n102 163.367
R396 B.n274 B.n273 163.367
R397 B.n275 B.n274 163.367
R398 B.n275 B.n100 163.367
R399 B.n279 B.n100 163.367
R400 B.n280 B.n279 163.367
R401 B.n281 B.n280 163.367
R402 B.n281 B.n98 163.367
R403 B.n285 B.n98 163.367
R404 B.n286 B.n285 163.367
R405 B.n287 B.n286 163.367
R406 B.n287 B.n96 163.367
R407 B.n291 B.n96 163.367
R408 B.n292 B.n291 163.367
R409 B.n293 B.n292 163.367
R410 B.n293 B.n94 163.367
R411 B.n297 B.n94 163.367
R412 B.n298 B.n297 163.367
R413 B.n299 B.n298 163.367
R414 B.n299 B.n92 163.367
R415 B.n303 B.n92 163.367
R416 B.n304 B.n303 163.367
R417 B.n305 B.n90 163.367
R418 B.n309 B.n90 163.367
R419 B.n310 B.n309 163.367
R420 B.n311 B.n310 163.367
R421 B.n311 B.n88 163.367
R422 B.n315 B.n88 163.367
R423 B.n316 B.n315 163.367
R424 B.n317 B.n316 163.367
R425 B.n317 B.n86 163.367
R426 B.n321 B.n86 163.367
R427 B.n322 B.n321 163.367
R428 B.n323 B.n322 163.367
R429 B.n323 B.n84 163.367
R430 B.n327 B.n84 163.367
R431 B.n328 B.n327 163.367
R432 B.n329 B.n328 163.367
R433 B.n329 B.n82 163.367
R434 B.n333 B.n82 163.367
R435 B.n334 B.n333 163.367
R436 B.n335 B.n334 163.367
R437 B.n335 B.n80 163.367
R438 B.n339 B.n80 163.367
R439 B.n340 B.n339 163.367
R440 B.n341 B.n340 163.367
R441 B.n341 B.n78 163.367
R442 B.n345 B.n78 163.367
R443 B.n346 B.n345 163.367
R444 B.n347 B.n346 163.367
R445 B.n347 B.n76 163.367
R446 B.n351 B.n76 163.367
R447 B.n352 B.n351 163.367
R448 B.n353 B.n352 163.367
R449 B.n353 B.n74 163.367
R450 B.n357 B.n74 163.367
R451 B.n358 B.n357 163.367
R452 B.n359 B.n358 163.367
R453 B.n359 B.n72 163.367
R454 B.n363 B.n72 163.367
R455 B.n364 B.n363 163.367
R456 B.n365 B.n364 163.367
R457 B.n365 B.n70 163.367
R458 B.n369 B.n70 163.367
R459 B.n370 B.n369 163.367
R460 B.n371 B.n370 163.367
R461 B.n371 B.n68 163.367
R462 B.n375 B.n68 163.367
R463 B.n376 B.n375 163.367
R464 B.n377 B.n376 163.367
R465 B.n377 B.n66 163.367
R466 B.n381 B.n66 163.367
R467 B.n382 B.n381 163.367
R468 B.n383 B.n382 163.367
R469 B.n383 B.n64 163.367
R470 B.n387 B.n64 163.367
R471 B.n388 B.n387 163.367
R472 B.n389 B.n388 163.367
R473 B.n389 B.n62 163.367
R474 B.n393 B.n62 163.367
R475 B.n394 B.n393 163.367
R476 B.n395 B.n394 163.367
R477 B.n395 B.n60 163.367
R478 B.n399 B.n60 163.367
R479 B.n510 B.n509 163.367
R480 B.n509 B.n508 163.367
R481 B.n508 B.n19 163.367
R482 B.n504 B.n19 163.367
R483 B.n504 B.n503 163.367
R484 B.n503 B.n502 163.367
R485 B.n502 B.n21 163.367
R486 B.n498 B.n21 163.367
R487 B.n498 B.n497 163.367
R488 B.n497 B.n496 163.367
R489 B.n496 B.n23 163.367
R490 B.n492 B.n23 163.367
R491 B.n492 B.n491 163.367
R492 B.n491 B.n490 163.367
R493 B.n490 B.n25 163.367
R494 B.n486 B.n25 163.367
R495 B.n486 B.n485 163.367
R496 B.n485 B.n484 163.367
R497 B.n484 B.n27 163.367
R498 B.n480 B.n27 163.367
R499 B.n480 B.n479 163.367
R500 B.n479 B.n478 163.367
R501 B.n478 B.n29 163.367
R502 B.n474 B.n29 163.367
R503 B.n474 B.n473 163.367
R504 B.n473 B.n472 163.367
R505 B.n472 B.n31 163.367
R506 B.n468 B.n31 163.367
R507 B.n468 B.n467 163.367
R508 B.n467 B.n466 163.367
R509 B.n466 B.n33 163.367
R510 B.n461 B.n33 163.367
R511 B.n461 B.n460 163.367
R512 B.n460 B.n459 163.367
R513 B.n459 B.n37 163.367
R514 B.n455 B.n37 163.367
R515 B.n455 B.n454 163.367
R516 B.n454 B.n453 163.367
R517 B.n453 B.n39 163.367
R518 B.n449 B.n39 163.367
R519 B.n449 B.n448 163.367
R520 B.n448 B.n447 163.367
R521 B.n447 B.n41 163.367
R522 B.n443 B.n41 163.367
R523 B.n443 B.n442 163.367
R524 B.n442 B.n441 163.367
R525 B.n441 B.n46 163.367
R526 B.n437 B.n46 163.367
R527 B.n437 B.n436 163.367
R528 B.n436 B.n435 163.367
R529 B.n435 B.n48 163.367
R530 B.n431 B.n48 163.367
R531 B.n431 B.n430 163.367
R532 B.n430 B.n429 163.367
R533 B.n429 B.n50 163.367
R534 B.n425 B.n50 163.367
R535 B.n425 B.n424 163.367
R536 B.n424 B.n423 163.367
R537 B.n423 B.n52 163.367
R538 B.n419 B.n52 163.367
R539 B.n419 B.n418 163.367
R540 B.n418 B.n417 163.367
R541 B.n417 B.n54 163.367
R542 B.n413 B.n54 163.367
R543 B.n413 B.n412 163.367
R544 B.n412 B.n411 163.367
R545 B.n411 B.n56 163.367
R546 B.n407 B.n56 163.367
R547 B.n407 B.n406 163.367
R548 B.n406 B.n405 163.367
R549 B.n405 B.n58 163.367
R550 B.n401 B.n58 163.367
R551 B.n401 B.n400 163.367
R552 B.n107 B.t11 158.381
R553 B.n42 B.t4 158.381
R554 B.n115 B.t2 158.371
R555 B.n34 B.t7 158.371
R556 B.n108 B.t10 108.54
R557 B.n43 B.t5 108.54
R558 B.n116 B.t1 108.529
R559 B.n35 B.t8 108.529
R560 B.n109 B.n108 59.5399
R561 B.n241 B.n116 59.5399
R562 B.n463 B.n35 59.5399
R563 B.n44 B.n43 59.5399
R564 B.n108 B.n107 49.8429
R565 B.n116 B.n115 49.8429
R566 B.n35 B.n34 49.8429
R567 B.n43 B.n42 49.8429
R568 B.n512 B.n511 32.0005
R569 B.n398 B.n59 32.0005
R570 B.n306 B.n91 32.0005
R571 B.n193 B.n192 32.0005
R572 B B.n559 18.0485
R573 B.n511 B.n18 10.6151
R574 B.n507 B.n18 10.6151
R575 B.n507 B.n506 10.6151
R576 B.n506 B.n505 10.6151
R577 B.n505 B.n20 10.6151
R578 B.n501 B.n20 10.6151
R579 B.n501 B.n500 10.6151
R580 B.n500 B.n499 10.6151
R581 B.n499 B.n22 10.6151
R582 B.n495 B.n22 10.6151
R583 B.n495 B.n494 10.6151
R584 B.n494 B.n493 10.6151
R585 B.n493 B.n24 10.6151
R586 B.n489 B.n24 10.6151
R587 B.n489 B.n488 10.6151
R588 B.n488 B.n487 10.6151
R589 B.n487 B.n26 10.6151
R590 B.n483 B.n26 10.6151
R591 B.n483 B.n482 10.6151
R592 B.n482 B.n481 10.6151
R593 B.n481 B.n28 10.6151
R594 B.n477 B.n28 10.6151
R595 B.n477 B.n476 10.6151
R596 B.n476 B.n475 10.6151
R597 B.n475 B.n30 10.6151
R598 B.n471 B.n30 10.6151
R599 B.n471 B.n470 10.6151
R600 B.n470 B.n469 10.6151
R601 B.n469 B.n32 10.6151
R602 B.n465 B.n32 10.6151
R603 B.n465 B.n464 10.6151
R604 B.n462 B.n36 10.6151
R605 B.n458 B.n36 10.6151
R606 B.n458 B.n457 10.6151
R607 B.n457 B.n456 10.6151
R608 B.n456 B.n38 10.6151
R609 B.n452 B.n38 10.6151
R610 B.n452 B.n451 10.6151
R611 B.n451 B.n450 10.6151
R612 B.n450 B.n40 10.6151
R613 B.n446 B.n445 10.6151
R614 B.n445 B.n444 10.6151
R615 B.n444 B.n45 10.6151
R616 B.n440 B.n45 10.6151
R617 B.n440 B.n439 10.6151
R618 B.n439 B.n438 10.6151
R619 B.n438 B.n47 10.6151
R620 B.n434 B.n47 10.6151
R621 B.n434 B.n433 10.6151
R622 B.n433 B.n432 10.6151
R623 B.n432 B.n49 10.6151
R624 B.n428 B.n49 10.6151
R625 B.n428 B.n427 10.6151
R626 B.n427 B.n426 10.6151
R627 B.n426 B.n51 10.6151
R628 B.n422 B.n51 10.6151
R629 B.n422 B.n421 10.6151
R630 B.n421 B.n420 10.6151
R631 B.n420 B.n53 10.6151
R632 B.n416 B.n53 10.6151
R633 B.n416 B.n415 10.6151
R634 B.n415 B.n414 10.6151
R635 B.n414 B.n55 10.6151
R636 B.n410 B.n55 10.6151
R637 B.n410 B.n409 10.6151
R638 B.n409 B.n408 10.6151
R639 B.n408 B.n57 10.6151
R640 B.n404 B.n57 10.6151
R641 B.n404 B.n403 10.6151
R642 B.n403 B.n402 10.6151
R643 B.n402 B.n59 10.6151
R644 B.n307 B.n306 10.6151
R645 B.n308 B.n307 10.6151
R646 B.n308 B.n89 10.6151
R647 B.n312 B.n89 10.6151
R648 B.n313 B.n312 10.6151
R649 B.n314 B.n313 10.6151
R650 B.n314 B.n87 10.6151
R651 B.n318 B.n87 10.6151
R652 B.n319 B.n318 10.6151
R653 B.n320 B.n319 10.6151
R654 B.n320 B.n85 10.6151
R655 B.n324 B.n85 10.6151
R656 B.n325 B.n324 10.6151
R657 B.n326 B.n325 10.6151
R658 B.n326 B.n83 10.6151
R659 B.n330 B.n83 10.6151
R660 B.n331 B.n330 10.6151
R661 B.n332 B.n331 10.6151
R662 B.n332 B.n81 10.6151
R663 B.n336 B.n81 10.6151
R664 B.n337 B.n336 10.6151
R665 B.n338 B.n337 10.6151
R666 B.n338 B.n79 10.6151
R667 B.n342 B.n79 10.6151
R668 B.n343 B.n342 10.6151
R669 B.n344 B.n343 10.6151
R670 B.n344 B.n77 10.6151
R671 B.n348 B.n77 10.6151
R672 B.n349 B.n348 10.6151
R673 B.n350 B.n349 10.6151
R674 B.n350 B.n75 10.6151
R675 B.n354 B.n75 10.6151
R676 B.n355 B.n354 10.6151
R677 B.n356 B.n355 10.6151
R678 B.n356 B.n73 10.6151
R679 B.n360 B.n73 10.6151
R680 B.n361 B.n360 10.6151
R681 B.n362 B.n361 10.6151
R682 B.n362 B.n71 10.6151
R683 B.n366 B.n71 10.6151
R684 B.n367 B.n366 10.6151
R685 B.n368 B.n367 10.6151
R686 B.n368 B.n69 10.6151
R687 B.n372 B.n69 10.6151
R688 B.n373 B.n372 10.6151
R689 B.n374 B.n373 10.6151
R690 B.n374 B.n67 10.6151
R691 B.n378 B.n67 10.6151
R692 B.n379 B.n378 10.6151
R693 B.n380 B.n379 10.6151
R694 B.n380 B.n65 10.6151
R695 B.n384 B.n65 10.6151
R696 B.n385 B.n384 10.6151
R697 B.n386 B.n385 10.6151
R698 B.n386 B.n63 10.6151
R699 B.n390 B.n63 10.6151
R700 B.n391 B.n390 10.6151
R701 B.n392 B.n391 10.6151
R702 B.n392 B.n61 10.6151
R703 B.n396 B.n61 10.6151
R704 B.n397 B.n396 10.6151
R705 B.n398 B.n397 10.6151
R706 B.n194 B.n193 10.6151
R707 B.n194 B.n131 10.6151
R708 B.n198 B.n131 10.6151
R709 B.n199 B.n198 10.6151
R710 B.n200 B.n199 10.6151
R711 B.n200 B.n129 10.6151
R712 B.n204 B.n129 10.6151
R713 B.n205 B.n204 10.6151
R714 B.n206 B.n205 10.6151
R715 B.n206 B.n127 10.6151
R716 B.n210 B.n127 10.6151
R717 B.n211 B.n210 10.6151
R718 B.n212 B.n211 10.6151
R719 B.n212 B.n125 10.6151
R720 B.n216 B.n125 10.6151
R721 B.n217 B.n216 10.6151
R722 B.n218 B.n217 10.6151
R723 B.n218 B.n123 10.6151
R724 B.n222 B.n123 10.6151
R725 B.n223 B.n222 10.6151
R726 B.n224 B.n223 10.6151
R727 B.n224 B.n121 10.6151
R728 B.n228 B.n121 10.6151
R729 B.n229 B.n228 10.6151
R730 B.n230 B.n229 10.6151
R731 B.n230 B.n119 10.6151
R732 B.n234 B.n119 10.6151
R733 B.n235 B.n234 10.6151
R734 B.n236 B.n235 10.6151
R735 B.n236 B.n117 10.6151
R736 B.n240 B.n117 10.6151
R737 B.n243 B.n242 10.6151
R738 B.n243 B.n113 10.6151
R739 B.n247 B.n113 10.6151
R740 B.n248 B.n247 10.6151
R741 B.n249 B.n248 10.6151
R742 B.n249 B.n111 10.6151
R743 B.n253 B.n111 10.6151
R744 B.n254 B.n253 10.6151
R745 B.n255 B.n254 10.6151
R746 B.n259 B.n258 10.6151
R747 B.n260 B.n259 10.6151
R748 B.n260 B.n105 10.6151
R749 B.n264 B.n105 10.6151
R750 B.n265 B.n264 10.6151
R751 B.n266 B.n265 10.6151
R752 B.n266 B.n103 10.6151
R753 B.n270 B.n103 10.6151
R754 B.n271 B.n270 10.6151
R755 B.n272 B.n271 10.6151
R756 B.n272 B.n101 10.6151
R757 B.n276 B.n101 10.6151
R758 B.n277 B.n276 10.6151
R759 B.n278 B.n277 10.6151
R760 B.n278 B.n99 10.6151
R761 B.n282 B.n99 10.6151
R762 B.n283 B.n282 10.6151
R763 B.n284 B.n283 10.6151
R764 B.n284 B.n97 10.6151
R765 B.n288 B.n97 10.6151
R766 B.n289 B.n288 10.6151
R767 B.n290 B.n289 10.6151
R768 B.n290 B.n95 10.6151
R769 B.n294 B.n95 10.6151
R770 B.n295 B.n294 10.6151
R771 B.n296 B.n295 10.6151
R772 B.n296 B.n93 10.6151
R773 B.n300 B.n93 10.6151
R774 B.n301 B.n300 10.6151
R775 B.n302 B.n301 10.6151
R776 B.n302 B.n91 10.6151
R777 B.n192 B.n133 10.6151
R778 B.n188 B.n133 10.6151
R779 B.n188 B.n187 10.6151
R780 B.n187 B.n186 10.6151
R781 B.n186 B.n135 10.6151
R782 B.n182 B.n135 10.6151
R783 B.n182 B.n181 10.6151
R784 B.n181 B.n180 10.6151
R785 B.n180 B.n137 10.6151
R786 B.n176 B.n137 10.6151
R787 B.n176 B.n175 10.6151
R788 B.n175 B.n174 10.6151
R789 B.n174 B.n139 10.6151
R790 B.n170 B.n139 10.6151
R791 B.n170 B.n169 10.6151
R792 B.n169 B.n168 10.6151
R793 B.n168 B.n141 10.6151
R794 B.n164 B.n141 10.6151
R795 B.n164 B.n163 10.6151
R796 B.n163 B.n162 10.6151
R797 B.n162 B.n143 10.6151
R798 B.n158 B.n143 10.6151
R799 B.n158 B.n157 10.6151
R800 B.n157 B.n156 10.6151
R801 B.n156 B.n145 10.6151
R802 B.n152 B.n145 10.6151
R803 B.n152 B.n151 10.6151
R804 B.n151 B.n150 10.6151
R805 B.n150 B.n147 10.6151
R806 B.n147 B.n0 10.6151
R807 B.n555 B.n1 10.6151
R808 B.n555 B.n554 10.6151
R809 B.n554 B.n553 10.6151
R810 B.n553 B.n4 10.6151
R811 B.n549 B.n4 10.6151
R812 B.n549 B.n548 10.6151
R813 B.n548 B.n547 10.6151
R814 B.n547 B.n6 10.6151
R815 B.n543 B.n6 10.6151
R816 B.n543 B.n542 10.6151
R817 B.n542 B.n541 10.6151
R818 B.n541 B.n8 10.6151
R819 B.n537 B.n8 10.6151
R820 B.n537 B.n536 10.6151
R821 B.n536 B.n535 10.6151
R822 B.n535 B.n10 10.6151
R823 B.n531 B.n10 10.6151
R824 B.n531 B.n530 10.6151
R825 B.n530 B.n529 10.6151
R826 B.n529 B.n12 10.6151
R827 B.n525 B.n12 10.6151
R828 B.n525 B.n524 10.6151
R829 B.n524 B.n523 10.6151
R830 B.n523 B.n14 10.6151
R831 B.n519 B.n14 10.6151
R832 B.n519 B.n518 10.6151
R833 B.n518 B.n517 10.6151
R834 B.n517 B.n16 10.6151
R835 B.n513 B.n16 10.6151
R836 B.n513 B.n512 10.6151
R837 B.n464 B.n463 9.36635
R838 B.n446 B.n44 9.36635
R839 B.n241 B.n240 9.36635
R840 B.n258 B.n109 9.36635
R841 B.n559 B.n0 2.81026
R842 B.n559 B.n1 2.81026
R843 B.n463 B.n462 1.24928
R844 B.n44 B.n40 1.24928
R845 B.n242 B.n241 1.24928
R846 B.n255 B.n109 1.24928
R847 VP.n12 VP.n0 161.3
R848 VP.n11 VP.n10 161.3
R849 VP.n9 VP.n1 161.3
R850 VP.n8 VP.n7 161.3
R851 VP.n6 VP.n2 161.3
R852 VP.n3 VP.t2 131.358
R853 VP.n3 VP.t3 130.714
R854 VP.n5 VP.n4 96.8909
R855 VP.n14 VP.n13 96.8909
R856 VP.n5 VP.t1 95.3246
R857 VP.n13 VP.t0 95.3246
R858 VP.n4 VP.n3 48.4936
R859 VP.n7 VP.n1 40.577
R860 VP.n11 VP.n1 40.577
R861 VP.n7 VP.n6 24.5923
R862 VP.n12 VP.n11 24.5923
R863 VP.n6 VP.n5 14.0178
R864 VP.n13 VP.n12 14.0178
R865 VP.n4 VP.n2 0.278335
R866 VP.n14 VP.n0 0.278335
R867 VP.n8 VP.n2 0.189894
R868 VP.n9 VP.n8 0.189894
R869 VP.n10 VP.n9 0.189894
R870 VP.n10 VP.n0 0.189894
R871 VP VP.n14 0.153485
R872 VTAIL.n5 VTAIL.t5 66.0076
R873 VTAIL.n4 VTAIL.t0 66.0076
R874 VTAIL.n3 VTAIL.t3 66.0076
R875 VTAIL.n6 VTAIL.t4 66.0073
R876 VTAIL.n7 VTAIL.t2 66.0073
R877 VTAIL.n0 VTAIL.t1 66.0073
R878 VTAIL.n1 VTAIL.t7 66.0073
R879 VTAIL.n2 VTAIL.t6 66.0073
R880 VTAIL.n7 VTAIL.n6 22.2203
R881 VTAIL.n3 VTAIL.n2 22.2203
R882 VTAIL.n4 VTAIL.n3 2.21602
R883 VTAIL.n6 VTAIL.n5 2.21602
R884 VTAIL.n2 VTAIL.n1 2.21602
R885 VTAIL VTAIL.n0 1.16645
R886 VTAIL VTAIL.n7 1.05007
R887 VTAIL.n5 VTAIL.n4 0.470328
R888 VTAIL.n1 VTAIL.n0 0.470328
R889 VDD1 VDD1.n1 117.541
R890 VDD1 VDD1.n0 79.0757
R891 VDD1.n0 VDD1.t1 3.66924
R892 VDD1.n0 VDD1.t0 3.66924
R893 VDD1.n1 VDD1.t2 3.66924
R894 VDD1.n1 VDD1.t3 3.66924
R895 VN.n0 VN.t2 131.358
R896 VN.n1 VN.t1 131.358
R897 VN.n0 VN.t3 130.714
R898 VN.n1 VN.t0 130.714
R899 VN VN.n1 48.7724
R900 VN VN.n0 5.71558
R901 VDD2.n2 VDD2.n0 117.016
R902 VDD2.n2 VDD2.n1 79.0175
R903 VDD2.n1 VDD2.t3 3.66924
R904 VDD2.n1 VDD2.t2 3.66924
R905 VDD2.n0 VDD2.t1 3.66924
R906 VDD2.n0 VDD2.t0 3.66924
R907 VDD2 VDD2.n2 0.0586897
C0 VDD1 VP 3.71542f
C1 B VP 1.53968f
C2 VDD1 B 1.11497f
C3 w_n2512_n2740# VP 4.45335f
C4 VDD1 w_n2512_n2740# 1.29647f
C5 w_n2512_n2740# B 7.92307f
C6 VTAIL VP 3.4985f
C7 VDD1 VTAIL 4.58044f
C8 VDD2 VP 0.371561f
C9 VTAIL B 3.77052f
C10 VDD1 VDD2 0.941919f
C11 VDD2 B 1.1612f
C12 VN VP 5.34808f
C13 VTAIL w_n2512_n2740# 3.25682f
C14 VDD1 VN 0.148838f
C15 w_n2512_n2740# VDD2 1.34453f
C16 VN B 1.00699f
C17 w_n2512_n2740# VN 4.13133f
C18 VTAIL VDD2 4.63223f
C19 VTAIL VN 3.48439f
C20 VN VDD2 3.49335f
C21 VDD2 VSUBS 0.805649f
C22 VDD1 VSUBS 5.10271f
C23 VTAIL VSUBS 1.021157f
C24 VN VSUBS 5.198599f
C25 VP VSUBS 1.983693f
C26 B VSUBS 3.695606f
C27 w_n2512_n2740# VSUBS 85.2171f
C28 VDD2.t1 VSUBS 0.188468f
C29 VDD2.t0 VSUBS 0.188468f
C30 VDD2.n0 VSUBS 1.93931f
C31 VDD2.t3 VSUBS 0.188468f
C32 VDD2.t2 VSUBS 0.188468f
C33 VDD2.n1 VSUBS 1.38797f
C34 VDD2.n2 VSUBS 3.82088f
C35 VN.t2 VSUBS 2.32711f
C36 VN.t3 VSUBS 2.32241f
C37 VN.n0 VSUBS 1.52823f
C38 VN.t1 VSUBS 2.32711f
C39 VN.t0 VSUBS 2.32241f
C40 VN.n1 VSUBS 3.29928f
C41 VDD1.t1 VSUBS 0.19078f
C42 VDD1.t0 VSUBS 0.19078f
C43 VDD1.n0 VSUBS 1.40551f
C44 VDD1.t2 VSUBS 0.19078f
C45 VDD1.t3 VSUBS 0.19078f
C46 VDD1.n1 VSUBS 1.98622f
C47 VTAIL.t1 VSUBS 1.55513f
C48 VTAIL.n0 VSUBS 0.730253f
C49 VTAIL.t7 VSUBS 1.55513f
C50 VTAIL.n1 VSUBS 0.814109f
C51 VTAIL.t6 VSUBS 1.55513f
C52 VTAIL.n2 VSUBS 1.90063f
C53 VTAIL.t3 VSUBS 1.55514f
C54 VTAIL.n3 VSUBS 1.90062f
C55 VTAIL.t0 VSUBS 1.55514f
C56 VTAIL.n4 VSUBS 0.814104f
C57 VTAIL.t5 VSUBS 1.55514f
C58 VTAIL.n5 VSUBS 0.814104f
C59 VTAIL.t4 VSUBS 1.55513f
C60 VTAIL.n6 VSUBS 1.90063f
C61 VTAIL.t2 VSUBS 1.55513f
C62 VTAIL.n7 VSUBS 1.80748f
C63 VP.n0 VSUBS 0.052798f
C64 VP.t0 VSUBS 2.14372f
C65 VP.n1 VSUBS 0.032347f
C66 VP.n2 VSUBS 0.052798f
C67 VP.t1 VSUBS 2.14372f
C68 VP.t3 VSUBS 2.41535f
C69 VP.t2 VSUBS 2.42024f
C70 VP.n3 VSUBS 3.41039f
C71 VP.n4 VSUBS 2.02688f
C72 VP.n5 VSUBS 0.9017f
C73 VP.n6 VSUBS 0.058503f
C74 VP.n7 VSUBS 0.079179f
C75 VP.n8 VSUBS 0.04005f
C76 VP.n9 VSUBS 0.04005f
C77 VP.n10 VSUBS 0.04005f
C78 VP.n11 VSUBS 0.079179f
C79 VP.n12 VSUBS 0.058503f
C80 VP.n13 VSUBS 0.9017f
C81 VP.n14 VSUBS 0.056975f
C82 B.n0 VSUBS 0.004759f
C83 B.n1 VSUBS 0.004759f
C84 B.n2 VSUBS 0.007526f
C85 B.n3 VSUBS 0.007526f
C86 B.n4 VSUBS 0.007526f
C87 B.n5 VSUBS 0.007526f
C88 B.n6 VSUBS 0.007526f
C89 B.n7 VSUBS 0.007526f
C90 B.n8 VSUBS 0.007526f
C91 B.n9 VSUBS 0.007526f
C92 B.n10 VSUBS 0.007526f
C93 B.n11 VSUBS 0.007526f
C94 B.n12 VSUBS 0.007526f
C95 B.n13 VSUBS 0.007526f
C96 B.n14 VSUBS 0.007526f
C97 B.n15 VSUBS 0.007526f
C98 B.n16 VSUBS 0.007526f
C99 B.n17 VSUBS 0.017232f
C100 B.n18 VSUBS 0.007526f
C101 B.n19 VSUBS 0.007526f
C102 B.n20 VSUBS 0.007526f
C103 B.n21 VSUBS 0.007526f
C104 B.n22 VSUBS 0.007526f
C105 B.n23 VSUBS 0.007526f
C106 B.n24 VSUBS 0.007526f
C107 B.n25 VSUBS 0.007526f
C108 B.n26 VSUBS 0.007526f
C109 B.n27 VSUBS 0.007526f
C110 B.n28 VSUBS 0.007526f
C111 B.n29 VSUBS 0.007526f
C112 B.n30 VSUBS 0.007526f
C113 B.n31 VSUBS 0.007526f
C114 B.n32 VSUBS 0.007526f
C115 B.n33 VSUBS 0.007526f
C116 B.t8 VSUBS 0.298721f
C117 B.t7 VSUBS 0.319028f
C118 B.t6 VSUBS 0.980203f
C119 B.n34 VSUBS 0.164272f
C120 B.n35 VSUBS 0.07526f
C121 B.n36 VSUBS 0.007526f
C122 B.n37 VSUBS 0.007526f
C123 B.n38 VSUBS 0.007526f
C124 B.n39 VSUBS 0.007526f
C125 B.n40 VSUBS 0.004206f
C126 B.n41 VSUBS 0.007526f
C127 B.t5 VSUBS 0.298717f
C128 B.t4 VSUBS 0.319025f
C129 B.t3 VSUBS 0.980203f
C130 B.n42 VSUBS 0.164276f
C131 B.n43 VSUBS 0.075263f
C132 B.n44 VSUBS 0.017437f
C133 B.n45 VSUBS 0.007526f
C134 B.n46 VSUBS 0.007526f
C135 B.n47 VSUBS 0.007526f
C136 B.n48 VSUBS 0.007526f
C137 B.n49 VSUBS 0.007526f
C138 B.n50 VSUBS 0.007526f
C139 B.n51 VSUBS 0.007526f
C140 B.n52 VSUBS 0.007526f
C141 B.n53 VSUBS 0.007526f
C142 B.n54 VSUBS 0.007526f
C143 B.n55 VSUBS 0.007526f
C144 B.n56 VSUBS 0.007526f
C145 B.n57 VSUBS 0.007526f
C146 B.n58 VSUBS 0.007526f
C147 B.n59 VSUBS 0.016613f
C148 B.n60 VSUBS 0.007526f
C149 B.n61 VSUBS 0.007526f
C150 B.n62 VSUBS 0.007526f
C151 B.n63 VSUBS 0.007526f
C152 B.n64 VSUBS 0.007526f
C153 B.n65 VSUBS 0.007526f
C154 B.n66 VSUBS 0.007526f
C155 B.n67 VSUBS 0.007526f
C156 B.n68 VSUBS 0.007526f
C157 B.n69 VSUBS 0.007526f
C158 B.n70 VSUBS 0.007526f
C159 B.n71 VSUBS 0.007526f
C160 B.n72 VSUBS 0.007526f
C161 B.n73 VSUBS 0.007526f
C162 B.n74 VSUBS 0.007526f
C163 B.n75 VSUBS 0.007526f
C164 B.n76 VSUBS 0.007526f
C165 B.n77 VSUBS 0.007526f
C166 B.n78 VSUBS 0.007526f
C167 B.n79 VSUBS 0.007526f
C168 B.n80 VSUBS 0.007526f
C169 B.n81 VSUBS 0.007526f
C170 B.n82 VSUBS 0.007526f
C171 B.n83 VSUBS 0.007526f
C172 B.n84 VSUBS 0.007526f
C173 B.n85 VSUBS 0.007526f
C174 B.n86 VSUBS 0.007526f
C175 B.n87 VSUBS 0.007526f
C176 B.n88 VSUBS 0.007526f
C177 B.n89 VSUBS 0.007526f
C178 B.n90 VSUBS 0.007526f
C179 B.n91 VSUBS 0.01752f
C180 B.n92 VSUBS 0.007526f
C181 B.n93 VSUBS 0.007526f
C182 B.n94 VSUBS 0.007526f
C183 B.n95 VSUBS 0.007526f
C184 B.n96 VSUBS 0.007526f
C185 B.n97 VSUBS 0.007526f
C186 B.n98 VSUBS 0.007526f
C187 B.n99 VSUBS 0.007526f
C188 B.n100 VSUBS 0.007526f
C189 B.n101 VSUBS 0.007526f
C190 B.n102 VSUBS 0.007526f
C191 B.n103 VSUBS 0.007526f
C192 B.n104 VSUBS 0.007526f
C193 B.n105 VSUBS 0.007526f
C194 B.n106 VSUBS 0.007526f
C195 B.t10 VSUBS 0.298717f
C196 B.t11 VSUBS 0.319025f
C197 B.t9 VSUBS 0.980203f
C198 B.n107 VSUBS 0.164276f
C199 B.n108 VSUBS 0.075263f
C200 B.n109 VSUBS 0.017437f
C201 B.n110 VSUBS 0.007526f
C202 B.n111 VSUBS 0.007526f
C203 B.n112 VSUBS 0.007526f
C204 B.n113 VSUBS 0.007526f
C205 B.n114 VSUBS 0.007526f
C206 B.t1 VSUBS 0.298721f
C207 B.t2 VSUBS 0.319028f
C208 B.t0 VSUBS 0.980203f
C209 B.n115 VSUBS 0.164272f
C210 B.n116 VSUBS 0.07526f
C211 B.n117 VSUBS 0.007526f
C212 B.n118 VSUBS 0.007526f
C213 B.n119 VSUBS 0.007526f
C214 B.n120 VSUBS 0.007526f
C215 B.n121 VSUBS 0.007526f
C216 B.n122 VSUBS 0.007526f
C217 B.n123 VSUBS 0.007526f
C218 B.n124 VSUBS 0.007526f
C219 B.n125 VSUBS 0.007526f
C220 B.n126 VSUBS 0.007526f
C221 B.n127 VSUBS 0.007526f
C222 B.n128 VSUBS 0.007526f
C223 B.n129 VSUBS 0.007526f
C224 B.n130 VSUBS 0.007526f
C225 B.n131 VSUBS 0.007526f
C226 B.n132 VSUBS 0.01752f
C227 B.n133 VSUBS 0.007526f
C228 B.n134 VSUBS 0.007526f
C229 B.n135 VSUBS 0.007526f
C230 B.n136 VSUBS 0.007526f
C231 B.n137 VSUBS 0.007526f
C232 B.n138 VSUBS 0.007526f
C233 B.n139 VSUBS 0.007526f
C234 B.n140 VSUBS 0.007526f
C235 B.n141 VSUBS 0.007526f
C236 B.n142 VSUBS 0.007526f
C237 B.n143 VSUBS 0.007526f
C238 B.n144 VSUBS 0.007526f
C239 B.n145 VSUBS 0.007526f
C240 B.n146 VSUBS 0.007526f
C241 B.n147 VSUBS 0.007526f
C242 B.n148 VSUBS 0.007526f
C243 B.n149 VSUBS 0.007526f
C244 B.n150 VSUBS 0.007526f
C245 B.n151 VSUBS 0.007526f
C246 B.n152 VSUBS 0.007526f
C247 B.n153 VSUBS 0.007526f
C248 B.n154 VSUBS 0.007526f
C249 B.n155 VSUBS 0.007526f
C250 B.n156 VSUBS 0.007526f
C251 B.n157 VSUBS 0.007526f
C252 B.n158 VSUBS 0.007526f
C253 B.n159 VSUBS 0.007526f
C254 B.n160 VSUBS 0.007526f
C255 B.n161 VSUBS 0.007526f
C256 B.n162 VSUBS 0.007526f
C257 B.n163 VSUBS 0.007526f
C258 B.n164 VSUBS 0.007526f
C259 B.n165 VSUBS 0.007526f
C260 B.n166 VSUBS 0.007526f
C261 B.n167 VSUBS 0.007526f
C262 B.n168 VSUBS 0.007526f
C263 B.n169 VSUBS 0.007526f
C264 B.n170 VSUBS 0.007526f
C265 B.n171 VSUBS 0.007526f
C266 B.n172 VSUBS 0.007526f
C267 B.n173 VSUBS 0.007526f
C268 B.n174 VSUBS 0.007526f
C269 B.n175 VSUBS 0.007526f
C270 B.n176 VSUBS 0.007526f
C271 B.n177 VSUBS 0.007526f
C272 B.n178 VSUBS 0.007526f
C273 B.n179 VSUBS 0.007526f
C274 B.n180 VSUBS 0.007526f
C275 B.n181 VSUBS 0.007526f
C276 B.n182 VSUBS 0.007526f
C277 B.n183 VSUBS 0.007526f
C278 B.n184 VSUBS 0.007526f
C279 B.n185 VSUBS 0.007526f
C280 B.n186 VSUBS 0.007526f
C281 B.n187 VSUBS 0.007526f
C282 B.n188 VSUBS 0.007526f
C283 B.n189 VSUBS 0.007526f
C284 B.n190 VSUBS 0.007526f
C285 B.n191 VSUBS 0.017232f
C286 B.n192 VSUBS 0.017232f
C287 B.n193 VSUBS 0.01752f
C288 B.n194 VSUBS 0.007526f
C289 B.n195 VSUBS 0.007526f
C290 B.n196 VSUBS 0.007526f
C291 B.n197 VSUBS 0.007526f
C292 B.n198 VSUBS 0.007526f
C293 B.n199 VSUBS 0.007526f
C294 B.n200 VSUBS 0.007526f
C295 B.n201 VSUBS 0.007526f
C296 B.n202 VSUBS 0.007526f
C297 B.n203 VSUBS 0.007526f
C298 B.n204 VSUBS 0.007526f
C299 B.n205 VSUBS 0.007526f
C300 B.n206 VSUBS 0.007526f
C301 B.n207 VSUBS 0.007526f
C302 B.n208 VSUBS 0.007526f
C303 B.n209 VSUBS 0.007526f
C304 B.n210 VSUBS 0.007526f
C305 B.n211 VSUBS 0.007526f
C306 B.n212 VSUBS 0.007526f
C307 B.n213 VSUBS 0.007526f
C308 B.n214 VSUBS 0.007526f
C309 B.n215 VSUBS 0.007526f
C310 B.n216 VSUBS 0.007526f
C311 B.n217 VSUBS 0.007526f
C312 B.n218 VSUBS 0.007526f
C313 B.n219 VSUBS 0.007526f
C314 B.n220 VSUBS 0.007526f
C315 B.n221 VSUBS 0.007526f
C316 B.n222 VSUBS 0.007526f
C317 B.n223 VSUBS 0.007526f
C318 B.n224 VSUBS 0.007526f
C319 B.n225 VSUBS 0.007526f
C320 B.n226 VSUBS 0.007526f
C321 B.n227 VSUBS 0.007526f
C322 B.n228 VSUBS 0.007526f
C323 B.n229 VSUBS 0.007526f
C324 B.n230 VSUBS 0.007526f
C325 B.n231 VSUBS 0.007526f
C326 B.n232 VSUBS 0.007526f
C327 B.n233 VSUBS 0.007526f
C328 B.n234 VSUBS 0.007526f
C329 B.n235 VSUBS 0.007526f
C330 B.n236 VSUBS 0.007526f
C331 B.n237 VSUBS 0.007526f
C332 B.n238 VSUBS 0.007526f
C333 B.n239 VSUBS 0.007526f
C334 B.n240 VSUBS 0.007083f
C335 B.n241 VSUBS 0.017437f
C336 B.n242 VSUBS 0.004206f
C337 B.n243 VSUBS 0.007526f
C338 B.n244 VSUBS 0.007526f
C339 B.n245 VSUBS 0.007526f
C340 B.n246 VSUBS 0.007526f
C341 B.n247 VSUBS 0.007526f
C342 B.n248 VSUBS 0.007526f
C343 B.n249 VSUBS 0.007526f
C344 B.n250 VSUBS 0.007526f
C345 B.n251 VSUBS 0.007526f
C346 B.n252 VSUBS 0.007526f
C347 B.n253 VSUBS 0.007526f
C348 B.n254 VSUBS 0.007526f
C349 B.n255 VSUBS 0.004206f
C350 B.n256 VSUBS 0.007526f
C351 B.n257 VSUBS 0.007526f
C352 B.n258 VSUBS 0.007083f
C353 B.n259 VSUBS 0.007526f
C354 B.n260 VSUBS 0.007526f
C355 B.n261 VSUBS 0.007526f
C356 B.n262 VSUBS 0.007526f
C357 B.n263 VSUBS 0.007526f
C358 B.n264 VSUBS 0.007526f
C359 B.n265 VSUBS 0.007526f
C360 B.n266 VSUBS 0.007526f
C361 B.n267 VSUBS 0.007526f
C362 B.n268 VSUBS 0.007526f
C363 B.n269 VSUBS 0.007526f
C364 B.n270 VSUBS 0.007526f
C365 B.n271 VSUBS 0.007526f
C366 B.n272 VSUBS 0.007526f
C367 B.n273 VSUBS 0.007526f
C368 B.n274 VSUBS 0.007526f
C369 B.n275 VSUBS 0.007526f
C370 B.n276 VSUBS 0.007526f
C371 B.n277 VSUBS 0.007526f
C372 B.n278 VSUBS 0.007526f
C373 B.n279 VSUBS 0.007526f
C374 B.n280 VSUBS 0.007526f
C375 B.n281 VSUBS 0.007526f
C376 B.n282 VSUBS 0.007526f
C377 B.n283 VSUBS 0.007526f
C378 B.n284 VSUBS 0.007526f
C379 B.n285 VSUBS 0.007526f
C380 B.n286 VSUBS 0.007526f
C381 B.n287 VSUBS 0.007526f
C382 B.n288 VSUBS 0.007526f
C383 B.n289 VSUBS 0.007526f
C384 B.n290 VSUBS 0.007526f
C385 B.n291 VSUBS 0.007526f
C386 B.n292 VSUBS 0.007526f
C387 B.n293 VSUBS 0.007526f
C388 B.n294 VSUBS 0.007526f
C389 B.n295 VSUBS 0.007526f
C390 B.n296 VSUBS 0.007526f
C391 B.n297 VSUBS 0.007526f
C392 B.n298 VSUBS 0.007526f
C393 B.n299 VSUBS 0.007526f
C394 B.n300 VSUBS 0.007526f
C395 B.n301 VSUBS 0.007526f
C396 B.n302 VSUBS 0.007526f
C397 B.n303 VSUBS 0.007526f
C398 B.n304 VSUBS 0.01752f
C399 B.n305 VSUBS 0.017232f
C400 B.n306 VSUBS 0.017232f
C401 B.n307 VSUBS 0.007526f
C402 B.n308 VSUBS 0.007526f
C403 B.n309 VSUBS 0.007526f
C404 B.n310 VSUBS 0.007526f
C405 B.n311 VSUBS 0.007526f
C406 B.n312 VSUBS 0.007526f
C407 B.n313 VSUBS 0.007526f
C408 B.n314 VSUBS 0.007526f
C409 B.n315 VSUBS 0.007526f
C410 B.n316 VSUBS 0.007526f
C411 B.n317 VSUBS 0.007526f
C412 B.n318 VSUBS 0.007526f
C413 B.n319 VSUBS 0.007526f
C414 B.n320 VSUBS 0.007526f
C415 B.n321 VSUBS 0.007526f
C416 B.n322 VSUBS 0.007526f
C417 B.n323 VSUBS 0.007526f
C418 B.n324 VSUBS 0.007526f
C419 B.n325 VSUBS 0.007526f
C420 B.n326 VSUBS 0.007526f
C421 B.n327 VSUBS 0.007526f
C422 B.n328 VSUBS 0.007526f
C423 B.n329 VSUBS 0.007526f
C424 B.n330 VSUBS 0.007526f
C425 B.n331 VSUBS 0.007526f
C426 B.n332 VSUBS 0.007526f
C427 B.n333 VSUBS 0.007526f
C428 B.n334 VSUBS 0.007526f
C429 B.n335 VSUBS 0.007526f
C430 B.n336 VSUBS 0.007526f
C431 B.n337 VSUBS 0.007526f
C432 B.n338 VSUBS 0.007526f
C433 B.n339 VSUBS 0.007526f
C434 B.n340 VSUBS 0.007526f
C435 B.n341 VSUBS 0.007526f
C436 B.n342 VSUBS 0.007526f
C437 B.n343 VSUBS 0.007526f
C438 B.n344 VSUBS 0.007526f
C439 B.n345 VSUBS 0.007526f
C440 B.n346 VSUBS 0.007526f
C441 B.n347 VSUBS 0.007526f
C442 B.n348 VSUBS 0.007526f
C443 B.n349 VSUBS 0.007526f
C444 B.n350 VSUBS 0.007526f
C445 B.n351 VSUBS 0.007526f
C446 B.n352 VSUBS 0.007526f
C447 B.n353 VSUBS 0.007526f
C448 B.n354 VSUBS 0.007526f
C449 B.n355 VSUBS 0.007526f
C450 B.n356 VSUBS 0.007526f
C451 B.n357 VSUBS 0.007526f
C452 B.n358 VSUBS 0.007526f
C453 B.n359 VSUBS 0.007526f
C454 B.n360 VSUBS 0.007526f
C455 B.n361 VSUBS 0.007526f
C456 B.n362 VSUBS 0.007526f
C457 B.n363 VSUBS 0.007526f
C458 B.n364 VSUBS 0.007526f
C459 B.n365 VSUBS 0.007526f
C460 B.n366 VSUBS 0.007526f
C461 B.n367 VSUBS 0.007526f
C462 B.n368 VSUBS 0.007526f
C463 B.n369 VSUBS 0.007526f
C464 B.n370 VSUBS 0.007526f
C465 B.n371 VSUBS 0.007526f
C466 B.n372 VSUBS 0.007526f
C467 B.n373 VSUBS 0.007526f
C468 B.n374 VSUBS 0.007526f
C469 B.n375 VSUBS 0.007526f
C470 B.n376 VSUBS 0.007526f
C471 B.n377 VSUBS 0.007526f
C472 B.n378 VSUBS 0.007526f
C473 B.n379 VSUBS 0.007526f
C474 B.n380 VSUBS 0.007526f
C475 B.n381 VSUBS 0.007526f
C476 B.n382 VSUBS 0.007526f
C477 B.n383 VSUBS 0.007526f
C478 B.n384 VSUBS 0.007526f
C479 B.n385 VSUBS 0.007526f
C480 B.n386 VSUBS 0.007526f
C481 B.n387 VSUBS 0.007526f
C482 B.n388 VSUBS 0.007526f
C483 B.n389 VSUBS 0.007526f
C484 B.n390 VSUBS 0.007526f
C485 B.n391 VSUBS 0.007526f
C486 B.n392 VSUBS 0.007526f
C487 B.n393 VSUBS 0.007526f
C488 B.n394 VSUBS 0.007526f
C489 B.n395 VSUBS 0.007526f
C490 B.n396 VSUBS 0.007526f
C491 B.n397 VSUBS 0.007526f
C492 B.n398 VSUBS 0.01814f
C493 B.n399 VSUBS 0.017232f
C494 B.n400 VSUBS 0.01752f
C495 B.n401 VSUBS 0.007526f
C496 B.n402 VSUBS 0.007526f
C497 B.n403 VSUBS 0.007526f
C498 B.n404 VSUBS 0.007526f
C499 B.n405 VSUBS 0.007526f
C500 B.n406 VSUBS 0.007526f
C501 B.n407 VSUBS 0.007526f
C502 B.n408 VSUBS 0.007526f
C503 B.n409 VSUBS 0.007526f
C504 B.n410 VSUBS 0.007526f
C505 B.n411 VSUBS 0.007526f
C506 B.n412 VSUBS 0.007526f
C507 B.n413 VSUBS 0.007526f
C508 B.n414 VSUBS 0.007526f
C509 B.n415 VSUBS 0.007526f
C510 B.n416 VSUBS 0.007526f
C511 B.n417 VSUBS 0.007526f
C512 B.n418 VSUBS 0.007526f
C513 B.n419 VSUBS 0.007526f
C514 B.n420 VSUBS 0.007526f
C515 B.n421 VSUBS 0.007526f
C516 B.n422 VSUBS 0.007526f
C517 B.n423 VSUBS 0.007526f
C518 B.n424 VSUBS 0.007526f
C519 B.n425 VSUBS 0.007526f
C520 B.n426 VSUBS 0.007526f
C521 B.n427 VSUBS 0.007526f
C522 B.n428 VSUBS 0.007526f
C523 B.n429 VSUBS 0.007526f
C524 B.n430 VSUBS 0.007526f
C525 B.n431 VSUBS 0.007526f
C526 B.n432 VSUBS 0.007526f
C527 B.n433 VSUBS 0.007526f
C528 B.n434 VSUBS 0.007526f
C529 B.n435 VSUBS 0.007526f
C530 B.n436 VSUBS 0.007526f
C531 B.n437 VSUBS 0.007526f
C532 B.n438 VSUBS 0.007526f
C533 B.n439 VSUBS 0.007526f
C534 B.n440 VSUBS 0.007526f
C535 B.n441 VSUBS 0.007526f
C536 B.n442 VSUBS 0.007526f
C537 B.n443 VSUBS 0.007526f
C538 B.n444 VSUBS 0.007526f
C539 B.n445 VSUBS 0.007526f
C540 B.n446 VSUBS 0.007083f
C541 B.n447 VSUBS 0.007526f
C542 B.n448 VSUBS 0.007526f
C543 B.n449 VSUBS 0.007526f
C544 B.n450 VSUBS 0.007526f
C545 B.n451 VSUBS 0.007526f
C546 B.n452 VSUBS 0.007526f
C547 B.n453 VSUBS 0.007526f
C548 B.n454 VSUBS 0.007526f
C549 B.n455 VSUBS 0.007526f
C550 B.n456 VSUBS 0.007526f
C551 B.n457 VSUBS 0.007526f
C552 B.n458 VSUBS 0.007526f
C553 B.n459 VSUBS 0.007526f
C554 B.n460 VSUBS 0.007526f
C555 B.n461 VSUBS 0.007526f
C556 B.n462 VSUBS 0.004206f
C557 B.n463 VSUBS 0.017437f
C558 B.n464 VSUBS 0.007083f
C559 B.n465 VSUBS 0.007526f
C560 B.n466 VSUBS 0.007526f
C561 B.n467 VSUBS 0.007526f
C562 B.n468 VSUBS 0.007526f
C563 B.n469 VSUBS 0.007526f
C564 B.n470 VSUBS 0.007526f
C565 B.n471 VSUBS 0.007526f
C566 B.n472 VSUBS 0.007526f
C567 B.n473 VSUBS 0.007526f
C568 B.n474 VSUBS 0.007526f
C569 B.n475 VSUBS 0.007526f
C570 B.n476 VSUBS 0.007526f
C571 B.n477 VSUBS 0.007526f
C572 B.n478 VSUBS 0.007526f
C573 B.n479 VSUBS 0.007526f
C574 B.n480 VSUBS 0.007526f
C575 B.n481 VSUBS 0.007526f
C576 B.n482 VSUBS 0.007526f
C577 B.n483 VSUBS 0.007526f
C578 B.n484 VSUBS 0.007526f
C579 B.n485 VSUBS 0.007526f
C580 B.n486 VSUBS 0.007526f
C581 B.n487 VSUBS 0.007526f
C582 B.n488 VSUBS 0.007526f
C583 B.n489 VSUBS 0.007526f
C584 B.n490 VSUBS 0.007526f
C585 B.n491 VSUBS 0.007526f
C586 B.n492 VSUBS 0.007526f
C587 B.n493 VSUBS 0.007526f
C588 B.n494 VSUBS 0.007526f
C589 B.n495 VSUBS 0.007526f
C590 B.n496 VSUBS 0.007526f
C591 B.n497 VSUBS 0.007526f
C592 B.n498 VSUBS 0.007526f
C593 B.n499 VSUBS 0.007526f
C594 B.n500 VSUBS 0.007526f
C595 B.n501 VSUBS 0.007526f
C596 B.n502 VSUBS 0.007526f
C597 B.n503 VSUBS 0.007526f
C598 B.n504 VSUBS 0.007526f
C599 B.n505 VSUBS 0.007526f
C600 B.n506 VSUBS 0.007526f
C601 B.n507 VSUBS 0.007526f
C602 B.n508 VSUBS 0.007526f
C603 B.n509 VSUBS 0.007526f
C604 B.n510 VSUBS 0.01752f
C605 B.n511 VSUBS 0.01752f
C606 B.n512 VSUBS 0.017232f
C607 B.n513 VSUBS 0.007526f
C608 B.n514 VSUBS 0.007526f
C609 B.n515 VSUBS 0.007526f
C610 B.n516 VSUBS 0.007526f
C611 B.n517 VSUBS 0.007526f
C612 B.n518 VSUBS 0.007526f
C613 B.n519 VSUBS 0.007526f
C614 B.n520 VSUBS 0.007526f
C615 B.n521 VSUBS 0.007526f
C616 B.n522 VSUBS 0.007526f
C617 B.n523 VSUBS 0.007526f
C618 B.n524 VSUBS 0.007526f
C619 B.n525 VSUBS 0.007526f
C620 B.n526 VSUBS 0.007526f
C621 B.n527 VSUBS 0.007526f
C622 B.n528 VSUBS 0.007526f
C623 B.n529 VSUBS 0.007526f
C624 B.n530 VSUBS 0.007526f
C625 B.n531 VSUBS 0.007526f
C626 B.n532 VSUBS 0.007526f
C627 B.n533 VSUBS 0.007526f
C628 B.n534 VSUBS 0.007526f
C629 B.n535 VSUBS 0.007526f
C630 B.n536 VSUBS 0.007526f
C631 B.n537 VSUBS 0.007526f
C632 B.n538 VSUBS 0.007526f
C633 B.n539 VSUBS 0.007526f
C634 B.n540 VSUBS 0.007526f
C635 B.n541 VSUBS 0.007526f
C636 B.n542 VSUBS 0.007526f
C637 B.n543 VSUBS 0.007526f
C638 B.n544 VSUBS 0.007526f
C639 B.n545 VSUBS 0.007526f
C640 B.n546 VSUBS 0.007526f
C641 B.n547 VSUBS 0.007526f
C642 B.n548 VSUBS 0.007526f
C643 B.n549 VSUBS 0.007526f
C644 B.n550 VSUBS 0.007526f
C645 B.n551 VSUBS 0.007526f
C646 B.n552 VSUBS 0.007526f
C647 B.n553 VSUBS 0.007526f
C648 B.n554 VSUBS 0.007526f
C649 B.n555 VSUBS 0.007526f
C650 B.n556 VSUBS 0.007526f
C651 B.n557 VSUBS 0.007526f
C652 B.n558 VSUBS 0.007526f
C653 B.n559 VSUBS 0.017042f
.ends

