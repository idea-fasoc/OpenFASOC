* NGSPICE file created from diff_pair_sample_1222.ext - technology: sky130A

.subckt diff_pair_sample_1222 VTAIL VN VP B VDD2 VDD1
X0 B.t17 B.t15 B.t16 B.t9 sky130_fd_pr__nfet_01v8 ad=3.2799 pd=17.6 as=0 ps=0 w=8.41 l=2.68
X1 VTAIL.t7 VP.t0 VDD1.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=3.2799 pd=17.6 as=1.38765 ps=8.74 w=8.41 l=2.68
X2 VTAIL.t0 VN.t0 VDD2.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=3.2799 pd=17.6 as=1.38765 ps=8.74 w=8.41 l=2.68
X3 VTAIL.t6 VP.t1 VDD1.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=3.2799 pd=17.6 as=1.38765 ps=8.74 w=8.41 l=2.68
X4 VDD1.t3 VP.t2 VTAIL.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=1.38765 pd=8.74 as=3.2799 ps=17.6 w=8.41 l=2.68
X5 B.t14 B.t12 B.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=3.2799 pd=17.6 as=0 ps=0 w=8.41 l=2.68
X6 VDD2.t2 VN.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.38765 pd=8.74 as=3.2799 ps=17.6 w=8.41 l=2.68
X7 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=3.2799 pd=17.6 as=0 ps=0 w=8.41 l=2.68
X8 VDD2.t1 VN.t2 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.38765 pd=8.74 as=3.2799 ps=17.6 w=8.41 l=2.68
X9 VTAIL.t3 VN.t3 VDD2.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=3.2799 pd=17.6 as=1.38765 ps=8.74 w=8.41 l=2.68
X10 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=3.2799 pd=17.6 as=0 ps=0 w=8.41 l=2.68
X11 VDD1.t1 VP.t3 VTAIL.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=1.38765 pd=8.74 as=3.2799 ps=17.6 w=8.41 l=2.68
R0 B.n506 B.n505 585
R1 B.n508 B.n106 585
R2 B.n511 B.n510 585
R3 B.n512 B.n105 585
R4 B.n514 B.n513 585
R5 B.n516 B.n104 585
R6 B.n519 B.n518 585
R7 B.n520 B.n103 585
R8 B.n522 B.n521 585
R9 B.n524 B.n102 585
R10 B.n527 B.n526 585
R11 B.n528 B.n101 585
R12 B.n530 B.n529 585
R13 B.n532 B.n100 585
R14 B.n535 B.n534 585
R15 B.n536 B.n99 585
R16 B.n538 B.n537 585
R17 B.n540 B.n98 585
R18 B.n543 B.n542 585
R19 B.n544 B.n97 585
R20 B.n546 B.n545 585
R21 B.n548 B.n96 585
R22 B.n551 B.n550 585
R23 B.n552 B.n95 585
R24 B.n554 B.n553 585
R25 B.n556 B.n94 585
R26 B.n559 B.n558 585
R27 B.n560 B.n93 585
R28 B.n562 B.n561 585
R29 B.n564 B.n92 585
R30 B.n567 B.n566 585
R31 B.n569 B.n89 585
R32 B.n571 B.n570 585
R33 B.n573 B.n88 585
R34 B.n576 B.n575 585
R35 B.n577 B.n87 585
R36 B.n579 B.n578 585
R37 B.n581 B.n86 585
R38 B.n584 B.n583 585
R39 B.n585 B.n82 585
R40 B.n587 B.n586 585
R41 B.n589 B.n81 585
R42 B.n592 B.n591 585
R43 B.n593 B.n80 585
R44 B.n595 B.n594 585
R45 B.n597 B.n79 585
R46 B.n600 B.n599 585
R47 B.n601 B.n78 585
R48 B.n603 B.n602 585
R49 B.n605 B.n77 585
R50 B.n608 B.n607 585
R51 B.n609 B.n76 585
R52 B.n611 B.n610 585
R53 B.n613 B.n75 585
R54 B.n616 B.n615 585
R55 B.n617 B.n74 585
R56 B.n619 B.n618 585
R57 B.n621 B.n73 585
R58 B.n624 B.n623 585
R59 B.n625 B.n72 585
R60 B.n627 B.n626 585
R61 B.n629 B.n71 585
R62 B.n632 B.n631 585
R63 B.n633 B.n70 585
R64 B.n635 B.n634 585
R65 B.n637 B.n69 585
R66 B.n640 B.n639 585
R67 B.n641 B.n68 585
R68 B.n643 B.n642 585
R69 B.n645 B.n67 585
R70 B.n648 B.n647 585
R71 B.n649 B.n66 585
R72 B.n504 B.n64 585
R73 B.n652 B.n64 585
R74 B.n503 B.n63 585
R75 B.n653 B.n63 585
R76 B.n502 B.n62 585
R77 B.n654 B.n62 585
R78 B.n501 B.n500 585
R79 B.n500 B.n58 585
R80 B.n499 B.n57 585
R81 B.n660 B.n57 585
R82 B.n498 B.n56 585
R83 B.n661 B.n56 585
R84 B.n497 B.n55 585
R85 B.n662 B.n55 585
R86 B.n496 B.n495 585
R87 B.n495 B.n54 585
R88 B.n494 B.n50 585
R89 B.n668 B.n50 585
R90 B.n493 B.n49 585
R91 B.n669 B.n49 585
R92 B.n492 B.n48 585
R93 B.n670 B.n48 585
R94 B.n491 B.n490 585
R95 B.n490 B.n44 585
R96 B.n489 B.n43 585
R97 B.n676 B.n43 585
R98 B.n488 B.n42 585
R99 B.n677 B.n42 585
R100 B.n487 B.n41 585
R101 B.n678 B.n41 585
R102 B.n486 B.n485 585
R103 B.n485 B.n37 585
R104 B.n484 B.n36 585
R105 B.n684 B.n36 585
R106 B.n483 B.n35 585
R107 B.n685 B.n35 585
R108 B.n482 B.n34 585
R109 B.n686 B.n34 585
R110 B.n481 B.n480 585
R111 B.n480 B.n33 585
R112 B.n479 B.n29 585
R113 B.n692 B.n29 585
R114 B.n478 B.n28 585
R115 B.n693 B.n28 585
R116 B.n477 B.n27 585
R117 B.n694 B.n27 585
R118 B.n476 B.n475 585
R119 B.n475 B.n23 585
R120 B.n474 B.n22 585
R121 B.n700 B.n22 585
R122 B.n473 B.n21 585
R123 B.n701 B.n21 585
R124 B.n472 B.n20 585
R125 B.n702 B.n20 585
R126 B.n471 B.n470 585
R127 B.n470 B.n16 585
R128 B.n469 B.n15 585
R129 B.n708 B.n15 585
R130 B.n468 B.n14 585
R131 B.n709 B.n14 585
R132 B.n467 B.n13 585
R133 B.n710 B.n13 585
R134 B.n466 B.n465 585
R135 B.n465 B.n12 585
R136 B.n464 B.n463 585
R137 B.n464 B.n8 585
R138 B.n462 B.n7 585
R139 B.n717 B.n7 585
R140 B.n461 B.n6 585
R141 B.n718 B.n6 585
R142 B.n460 B.n5 585
R143 B.n719 B.n5 585
R144 B.n459 B.n458 585
R145 B.n458 B.n4 585
R146 B.n457 B.n107 585
R147 B.n457 B.n456 585
R148 B.n447 B.n108 585
R149 B.n109 B.n108 585
R150 B.n449 B.n448 585
R151 B.n450 B.n449 585
R152 B.n446 B.n114 585
R153 B.n114 B.n113 585
R154 B.n445 B.n444 585
R155 B.n444 B.n443 585
R156 B.n116 B.n115 585
R157 B.n117 B.n116 585
R158 B.n436 B.n435 585
R159 B.n437 B.n436 585
R160 B.n434 B.n122 585
R161 B.n122 B.n121 585
R162 B.n433 B.n432 585
R163 B.n432 B.n431 585
R164 B.n124 B.n123 585
R165 B.n125 B.n124 585
R166 B.n424 B.n423 585
R167 B.n425 B.n424 585
R168 B.n422 B.n130 585
R169 B.n130 B.n129 585
R170 B.n421 B.n420 585
R171 B.n420 B.n419 585
R172 B.n132 B.n131 585
R173 B.n412 B.n132 585
R174 B.n411 B.n410 585
R175 B.n413 B.n411 585
R176 B.n409 B.n137 585
R177 B.n137 B.n136 585
R178 B.n408 B.n407 585
R179 B.n407 B.n406 585
R180 B.n139 B.n138 585
R181 B.n140 B.n139 585
R182 B.n399 B.n398 585
R183 B.n400 B.n399 585
R184 B.n397 B.n145 585
R185 B.n145 B.n144 585
R186 B.n396 B.n395 585
R187 B.n395 B.n394 585
R188 B.n147 B.n146 585
R189 B.n148 B.n147 585
R190 B.n387 B.n386 585
R191 B.n388 B.n387 585
R192 B.n385 B.n153 585
R193 B.n153 B.n152 585
R194 B.n384 B.n383 585
R195 B.n383 B.n382 585
R196 B.n155 B.n154 585
R197 B.n375 B.n155 585
R198 B.n374 B.n373 585
R199 B.n376 B.n374 585
R200 B.n372 B.n160 585
R201 B.n160 B.n159 585
R202 B.n371 B.n370 585
R203 B.n370 B.n369 585
R204 B.n162 B.n161 585
R205 B.n163 B.n162 585
R206 B.n362 B.n361 585
R207 B.n363 B.n362 585
R208 B.n360 B.n168 585
R209 B.n168 B.n167 585
R210 B.n359 B.n358 585
R211 B.n358 B.n357 585
R212 B.n354 B.n172 585
R213 B.n353 B.n352 585
R214 B.n350 B.n173 585
R215 B.n350 B.n171 585
R216 B.n349 B.n348 585
R217 B.n347 B.n346 585
R218 B.n345 B.n175 585
R219 B.n343 B.n342 585
R220 B.n341 B.n176 585
R221 B.n340 B.n339 585
R222 B.n337 B.n177 585
R223 B.n335 B.n334 585
R224 B.n333 B.n178 585
R225 B.n332 B.n331 585
R226 B.n329 B.n179 585
R227 B.n327 B.n326 585
R228 B.n325 B.n180 585
R229 B.n324 B.n323 585
R230 B.n321 B.n181 585
R231 B.n319 B.n318 585
R232 B.n317 B.n182 585
R233 B.n316 B.n315 585
R234 B.n313 B.n183 585
R235 B.n311 B.n310 585
R236 B.n309 B.n184 585
R237 B.n308 B.n307 585
R238 B.n305 B.n185 585
R239 B.n303 B.n302 585
R240 B.n301 B.n186 585
R241 B.n300 B.n299 585
R242 B.n297 B.n187 585
R243 B.n295 B.n294 585
R244 B.n292 B.n188 585
R245 B.n291 B.n290 585
R246 B.n288 B.n191 585
R247 B.n286 B.n285 585
R248 B.n284 B.n192 585
R249 B.n283 B.n282 585
R250 B.n280 B.n193 585
R251 B.n278 B.n277 585
R252 B.n276 B.n194 585
R253 B.n275 B.n274 585
R254 B.n272 B.n271 585
R255 B.n270 B.n269 585
R256 B.n268 B.n199 585
R257 B.n266 B.n265 585
R258 B.n264 B.n200 585
R259 B.n263 B.n262 585
R260 B.n260 B.n201 585
R261 B.n258 B.n257 585
R262 B.n256 B.n202 585
R263 B.n255 B.n254 585
R264 B.n252 B.n203 585
R265 B.n250 B.n249 585
R266 B.n248 B.n204 585
R267 B.n247 B.n246 585
R268 B.n244 B.n205 585
R269 B.n242 B.n241 585
R270 B.n240 B.n206 585
R271 B.n239 B.n238 585
R272 B.n236 B.n207 585
R273 B.n234 B.n233 585
R274 B.n232 B.n208 585
R275 B.n231 B.n230 585
R276 B.n228 B.n209 585
R277 B.n226 B.n225 585
R278 B.n224 B.n210 585
R279 B.n223 B.n222 585
R280 B.n220 B.n211 585
R281 B.n218 B.n217 585
R282 B.n216 B.n212 585
R283 B.n215 B.n214 585
R284 B.n170 B.n169 585
R285 B.n171 B.n170 585
R286 B.n356 B.n355 585
R287 B.n357 B.n356 585
R288 B.n166 B.n165 585
R289 B.n167 B.n166 585
R290 B.n365 B.n364 585
R291 B.n364 B.n363 585
R292 B.n366 B.n164 585
R293 B.n164 B.n163 585
R294 B.n368 B.n367 585
R295 B.n369 B.n368 585
R296 B.n158 B.n157 585
R297 B.n159 B.n158 585
R298 B.n378 B.n377 585
R299 B.n377 B.n376 585
R300 B.n379 B.n156 585
R301 B.n375 B.n156 585
R302 B.n381 B.n380 585
R303 B.n382 B.n381 585
R304 B.n151 B.n150 585
R305 B.n152 B.n151 585
R306 B.n390 B.n389 585
R307 B.n389 B.n388 585
R308 B.n391 B.n149 585
R309 B.n149 B.n148 585
R310 B.n393 B.n392 585
R311 B.n394 B.n393 585
R312 B.n143 B.n142 585
R313 B.n144 B.n143 585
R314 B.n402 B.n401 585
R315 B.n401 B.n400 585
R316 B.n403 B.n141 585
R317 B.n141 B.n140 585
R318 B.n405 B.n404 585
R319 B.n406 B.n405 585
R320 B.n135 B.n134 585
R321 B.n136 B.n135 585
R322 B.n415 B.n414 585
R323 B.n414 B.n413 585
R324 B.n416 B.n133 585
R325 B.n412 B.n133 585
R326 B.n418 B.n417 585
R327 B.n419 B.n418 585
R328 B.n128 B.n127 585
R329 B.n129 B.n128 585
R330 B.n427 B.n426 585
R331 B.n426 B.n425 585
R332 B.n428 B.n126 585
R333 B.n126 B.n125 585
R334 B.n430 B.n429 585
R335 B.n431 B.n430 585
R336 B.n120 B.n119 585
R337 B.n121 B.n120 585
R338 B.n439 B.n438 585
R339 B.n438 B.n437 585
R340 B.n440 B.n118 585
R341 B.n118 B.n117 585
R342 B.n442 B.n441 585
R343 B.n443 B.n442 585
R344 B.n112 B.n111 585
R345 B.n113 B.n112 585
R346 B.n452 B.n451 585
R347 B.n451 B.n450 585
R348 B.n453 B.n110 585
R349 B.n110 B.n109 585
R350 B.n455 B.n454 585
R351 B.n456 B.n455 585
R352 B.n3 B.n0 585
R353 B.n4 B.n3 585
R354 B.n716 B.n1 585
R355 B.n717 B.n716 585
R356 B.n715 B.n714 585
R357 B.n715 B.n8 585
R358 B.n713 B.n9 585
R359 B.n12 B.n9 585
R360 B.n712 B.n711 585
R361 B.n711 B.n710 585
R362 B.n11 B.n10 585
R363 B.n709 B.n11 585
R364 B.n707 B.n706 585
R365 B.n708 B.n707 585
R366 B.n705 B.n17 585
R367 B.n17 B.n16 585
R368 B.n704 B.n703 585
R369 B.n703 B.n702 585
R370 B.n19 B.n18 585
R371 B.n701 B.n19 585
R372 B.n699 B.n698 585
R373 B.n700 B.n699 585
R374 B.n697 B.n24 585
R375 B.n24 B.n23 585
R376 B.n696 B.n695 585
R377 B.n695 B.n694 585
R378 B.n26 B.n25 585
R379 B.n693 B.n26 585
R380 B.n691 B.n690 585
R381 B.n692 B.n691 585
R382 B.n689 B.n30 585
R383 B.n33 B.n30 585
R384 B.n688 B.n687 585
R385 B.n687 B.n686 585
R386 B.n32 B.n31 585
R387 B.n685 B.n32 585
R388 B.n683 B.n682 585
R389 B.n684 B.n683 585
R390 B.n681 B.n38 585
R391 B.n38 B.n37 585
R392 B.n680 B.n679 585
R393 B.n679 B.n678 585
R394 B.n40 B.n39 585
R395 B.n677 B.n40 585
R396 B.n675 B.n674 585
R397 B.n676 B.n675 585
R398 B.n673 B.n45 585
R399 B.n45 B.n44 585
R400 B.n672 B.n671 585
R401 B.n671 B.n670 585
R402 B.n47 B.n46 585
R403 B.n669 B.n47 585
R404 B.n667 B.n666 585
R405 B.n668 B.n667 585
R406 B.n665 B.n51 585
R407 B.n54 B.n51 585
R408 B.n664 B.n663 585
R409 B.n663 B.n662 585
R410 B.n53 B.n52 585
R411 B.n661 B.n53 585
R412 B.n659 B.n658 585
R413 B.n660 B.n659 585
R414 B.n657 B.n59 585
R415 B.n59 B.n58 585
R416 B.n656 B.n655 585
R417 B.n655 B.n654 585
R418 B.n61 B.n60 585
R419 B.n653 B.n61 585
R420 B.n651 B.n650 585
R421 B.n652 B.n651 585
R422 B.n720 B.n719 585
R423 B.n718 B.n2 585
R424 B.n651 B.n66 502.111
R425 B.n506 B.n64 502.111
R426 B.n358 B.n170 502.111
R427 B.n356 B.n172 502.111
R428 B.n83 B.t8 283.791
R429 B.n90 B.t15 283.791
R430 B.n195 B.t4 283.791
R431 B.n189 B.t12 283.791
R432 B.n507 B.n65 256.663
R433 B.n509 B.n65 256.663
R434 B.n515 B.n65 256.663
R435 B.n517 B.n65 256.663
R436 B.n523 B.n65 256.663
R437 B.n525 B.n65 256.663
R438 B.n531 B.n65 256.663
R439 B.n533 B.n65 256.663
R440 B.n539 B.n65 256.663
R441 B.n541 B.n65 256.663
R442 B.n547 B.n65 256.663
R443 B.n549 B.n65 256.663
R444 B.n555 B.n65 256.663
R445 B.n557 B.n65 256.663
R446 B.n563 B.n65 256.663
R447 B.n565 B.n65 256.663
R448 B.n572 B.n65 256.663
R449 B.n574 B.n65 256.663
R450 B.n580 B.n65 256.663
R451 B.n582 B.n65 256.663
R452 B.n588 B.n65 256.663
R453 B.n590 B.n65 256.663
R454 B.n596 B.n65 256.663
R455 B.n598 B.n65 256.663
R456 B.n604 B.n65 256.663
R457 B.n606 B.n65 256.663
R458 B.n612 B.n65 256.663
R459 B.n614 B.n65 256.663
R460 B.n620 B.n65 256.663
R461 B.n622 B.n65 256.663
R462 B.n628 B.n65 256.663
R463 B.n630 B.n65 256.663
R464 B.n636 B.n65 256.663
R465 B.n638 B.n65 256.663
R466 B.n644 B.n65 256.663
R467 B.n646 B.n65 256.663
R468 B.n351 B.n171 256.663
R469 B.n174 B.n171 256.663
R470 B.n344 B.n171 256.663
R471 B.n338 B.n171 256.663
R472 B.n336 B.n171 256.663
R473 B.n330 B.n171 256.663
R474 B.n328 B.n171 256.663
R475 B.n322 B.n171 256.663
R476 B.n320 B.n171 256.663
R477 B.n314 B.n171 256.663
R478 B.n312 B.n171 256.663
R479 B.n306 B.n171 256.663
R480 B.n304 B.n171 256.663
R481 B.n298 B.n171 256.663
R482 B.n296 B.n171 256.663
R483 B.n289 B.n171 256.663
R484 B.n287 B.n171 256.663
R485 B.n281 B.n171 256.663
R486 B.n279 B.n171 256.663
R487 B.n273 B.n171 256.663
R488 B.n198 B.n171 256.663
R489 B.n267 B.n171 256.663
R490 B.n261 B.n171 256.663
R491 B.n259 B.n171 256.663
R492 B.n253 B.n171 256.663
R493 B.n251 B.n171 256.663
R494 B.n245 B.n171 256.663
R495 B.n243 B.n171 256.663
R496 B.n237 B.n171 256.663
R497 B.n235 B.n171 256.663
R498 B.n229 B.n171 256.663
R499 B.n227 B.n171 256.663
R500 B.n221 B.n171 256.663
R501 B.n219 B.n171 256.663
R502 B.n213 B.n171 256.663
R503 B.n722 B.n721 256.663
R504 B.n647 B.n645 163.367
R505 B.n643 B.n68 163.367
R506 B.n639 B.n637 163.367
R507 B.n635 B.n70 163.367
R508 B.n631 B.n629 163.367
R509 B.n627 B.n72 163.367
R510 B.n623 B.n621 163.367
R511 B.n619 B.n74 163.367
R512 B.n615 B.n613 163.367
R513 B.n611 B.n76 163.367
R514 B.n607 B.n605 163.367
R515 B.n603 B.n78 163.367
R516 B.n599 B.n597 163.367
R517 B.n595 B.n80 163.367
R518 B.n591 B.n589 163.367
R519 B.n587 B.n82 163.367
R520 B.n583 B.n581 163.367
R521 B.n579 B.n87 163.367
R522 B.n575 B.n573 163.367
R523 B.n571 B.n89 163.367
R524 B.n566 B.n564 163.367
R525 B.n562 B.n93 163.367
R526 B.n558 B.n556 163.367
R527 B.n554 B.n95 163.367
R528 B.n550 B.n548 163.367
R529 B.n546 B.n97 163.367
R530 B.n542 B.n540 163.367
R531 B.n538 B.n99 163.367
R532 B.n534 B.n532 163.367
R533 B.n530 B.n101 163.367
R534 B.n526 B.n524 163.367
R535 B.n522 B.n103 163.367
R536 B.n518 B.n516 163.367
R537 B.n514 B.n105 163.367
R538 B.n510 B.n508 163.367
R539 B.n358 B.n168 163.367
R540 B.n362 B.n168 163.367
R541 B.n362 B.n162 163.367
R542 B.n370 B.n162 163.367
R543 B.n370 B.n160 163.367
R544 B.n374 B.n160 163.367
R545 B.n374 B.n155 163.367
R546 B.n383 B.n155 163.367
R547 B.n383 B.n153 163.367
R548 B.n387 B.n153 163.367
R549 B.n387 B.n147 163.367
R550 B.n395 B.n147 163.367
R551 B.n395 B.n145 163.367
R552 B.n399 B.n145 163.367
R553 B.n399 B.n139 163.367
R554 B.n407 B.n139 163.367
R555 B.n407 B.n137 163.367
R556 B.n411 B.n137 163.367
R557 B.n411 B.n132 163.367
R558 B.n420 B.n132 163.367
R559 B.n420 B.n130 163.367
R560 B.n424 B.n130 163.367
R561 B.n424 B.n124 163.367
R562 B.n432 B.n124 163.367
R563 B.n432 B.n122 163.367
R564 B.n436 B.n122 163.367
R565 B.n436 B.n116 163.367
R566 B.n444 B.n116 163.367
R567 B.n444 B.n114 163.367
R568 B.n449 B.n114 163.367
R569 B.n449 B.n108 163.367
R570 B.n457 B.n108 163.367
R571 B.n458 B.n457 163.367
R572 B.n458 B.n5 163.367
R573 B.n6 B.n5 163.367
R574 B.n7 B.n6 163.367
R575 B.n464 B.n7 163.367
R576 B.n465 B.n464 163.367
R577 B.n465 B.n13 163.367
R578 B.n14 B.n13 163.367
R579 B.n15 B.n14 163.367
R580 B.n470 B.n15 163.367
R581 B.n470 B.n20 163.367
R582 B.n21 B.n20 163.367
R583 B.n22 B.n21 163.367
R584 B.n475 B.n22 163.367
R585 B.n475 B.n27 163.367
R586 B.n28 B.n27 163.367
R587 B.n29 B.n28 163.367
R588 B.n480 B.n29 163.367
R589 B.n480 B.n34 163.367
R590 B.n35 B.n34 163.367
R591 B.n36 B.n35 163.367
R592 B.n485 B.n36 163.367
R593 B.n485 B.n41 163.367
R594 B.n42 B.n41 163.367
R595 B.n43 B.n42 163.367
R596 B.n490 B.n43 163.367
R597 B.n490 B.n48 163.367
R598 B.n49 B.n48 163.367
R599 B.n50 B.n49 163.367
R600 B.n495 B.n50 163.367
R601 B.n495 B.n55 163.367
R602 B.n56 B.n55 163.367
R603 B.n57 B.n56 163.367
R604 B.n500 B.n57 163.367
R605 B.n500 B.n62 163.367
R606 B.n63 B.n62 163.367
R607 B.n64 B.n63 163.367
R608 B.n352 B.n350 163.367
R609 B.n350 B.n349 163.367
R610 B.n346 B.n345 163.367
R611 B.n343 B.n176 163.367
R612 B.n339 B.n337 163.367
R613 B.n335 B.n178 163.367
R614 B.n331 B.n329 163.367
R615 B.n327 B.n180 163.367
R616 B.n323 B.n321 163.367
R617 B.n319 B.n182 163.367
R618 B.n315 B.n313 163.367
R619 B.n311 B.n184 163.367
R620 B.n307 B.n305 163.367
R621 B.n303 B.n186 163.367
R622 B.n299 B.n297 163.367
R623 B.n295 B.n188 163.367
R624 B.n290 B.n288 163.367
R625 B.n286 B.n192 163.367
R626 B.n282 B.n280 163.367
R627 B.n278 B.n194 163.367
R628 B.n274 B.n272 163.367
R629 B.n269 B.n268 163.367
R630 B.n266 B.n200 163.367
R631 B.n262 B.n260 163.367
R632 B.n258 B.n202 163.367
R633 B.n254 B.n252 163.367
R634 B.n250 B.n204 163.367
R635 B.n246 B.n244 163.367
R636 B.n242 B.n206 163.367
R637 B.n238 B.n236 163.367
R638 B.n234 B.n208 163.367
R639 B.n230 B.n228 163.367
R640 B.n226 B.n210 163.367
R641 B.n222 B.n220 163.367
R642 B.n218 B.n212 163.367
R643 B.n214 B.n170 163.367
R644 B.n356 B.n166 163.367
R645 B.n364 B.n166 163.367
R646 B.n364 B.n164 163.367
R647 B.n368 B.n164 163.367
R648 B.n368 B.n158 163.367
R649 B.n377 B.n158 163.367
R650 B.n377 B.n156 163.367
R651 B.n381 B.n156 163.367
R652 B.n381 B.n151 163.367
R653 B.n389 B.n151 163.367
R654 B.n389 B.n149 163.367
R655 B.n393 B.n149 163.367
R656 B.n393 B.n143 163.367
R657 B.n401 B.n143 163.367
R658 B.n401 B.n141 163.367
R659 B.n405 B.n141 163.367
R660 B.n405 B.n135 163.367
R661 B.n414 B.n135 163.367
R662 B.n414 B.n133 163.367
R663 B.n418 B.n133 163.367
R664 B.n418 B.n128 163.367
R665 B.n426 B.n128 163.367
R666 B.n426 B.n126 163.367
R667 B.n430 B.n126 163.367
R668 B.n430 B.n120 163.367
R669 B.n438 B.n120 163.367
R670 B.n438 B.n118 163.367
R671 B.n442 B.n118 163.367
R672 B.n442 B.n112 163.367
R673 B.n451 B.n112 163.367
R674 B.n451 B.n110 163.367
R675 B.n455 B.n110 163.367
R676 B.n455 B.n3 163.367
R677 B.n720 B.n3 163.367
R678 B.n716 B.n2 163.367
R679 B.n716 B.n715 163.367
R680 B.n715 B.n9 163.367
R681 B.n711 B.n9 163.367
R682 B.n711 B.n11 163.367
R683 B.n707 B.n11 163.367
R684 B.n707 B.n17 163.367
R685 B.n703 B.n17 163.367
R686 B.n703 B.n19 163.367
R687 B.n699 B.n19 163.367
R688 B.n699 B.n24 163.367
R689 B.n695 B.n24 163.367
R690 B.n695 B.n26 163.367
R691 B.n691 B.n26 163.367
R692 B.n691 B.n30 163.367
R693 B.n687 B.n30 163.367
R694 B.n687 B.n32 163.367
R695 B.n683 B.n32 163.367
R696 B.n683 B.n38 163.367
R697 B.n679 B.n38 163.367
R698 B.n679 B.n40 163.367
R699 B.n675 B.n40 163.367
R700 B.n675 B.n45 163.367
R701 B.n671 B.n45 163.367
R702 B.n671 B.n47 163.367
R703 B.n667 B.n47 163.367
R704 B.n667 B.n51 163.367
R705 B.n663 B.n51 163.367
R706 B.n663 B.n53 163.367
R707 B.n659 B.n53 163.367
R708 B.n659 B.n59 163.367
R709 B.n655 B.n59 163.367
R710 B.n655 B.n61 163.367
R711 B.n651 B.n61 163.367
R712 B.n90 B.t16 131.714
R713 B.n195 B.t7 131.714
R714 B.n83 B.t10 131.703
R715 B.n189 B.t14 131.703
R716 B.n357 B.n171 108.513
R717 B.n652 B.n65 108.513
R718 B.n91 B.t17 73.3377
R719 B.n196 B.t6 73.3377
R720 B.n84 B.t11 73.328
R721 B.n190 B.t13 73.328
R722 B.n646 B.n66 71.676
R723 B.n645 B.n644 71.676
R724 B.n638 B.n68 71.676
R725 B.n637 B.n636 71.676
R726 B.n630 B.n70 71.676
R727 B.n629 B.n628 71.676
R728 B.n622 B.n72 71.676
R729 B.n621 B.n620 71.676
R730 B.n614 B.n74 71.676
R731 B.n613 B.n612 71.676
R732 B.n606 B.n76 71.676
R733 B.n605 B.n604 71.676
R734 B.n598 B.n78 71.676
R735 B.n597 B.n596 71.676
R736 B.n590 B.n80 71.676
R737 B.n589 B.n588 71.676
R738 B.n582 B.n82 71.676
R739 B.n581 B.n580 71.676
R740 B.n574 B.n87 71.676
R741 B.n573 B.n572 71.676
R742 B.n565 B.n89 71.676
R743 B.n564 B.n563 71.676
R744 B.n557 B.n93 71.676
R745 B.n556 B.n555 71.676
R746 B.n549 B.n95 71.676
R747 B.n548 B.n547 71.676
R748 B.n541 B.n97 71.676
R749 B.n540 B.n539 71.676
R750 B.n533 B.n99 71.676
R751 B.n532 B.n531 71.676
R752 B.n525 B.n101 71.676
R753 B.n524 B.n523 71.676
R754 B.n517 B.n103 71.676
R755 B.n516 B.n515 71.676
R756 B.n509 B.n105 71.676
R757 B.n508 B.n507 71.676
R758 B.n507 B.n506 71.676
R759 B.n510 B.n509 71.676
R760 B.n515 B.n514 71.676
R761 B.n518 B.n517 71.676
R762 B.n523 B.n522 71.676
R763 B.n526 B.n525 71.676
R764 B.n531 B.n530 71.676
R765 B.n534 B.n533 71.676
R766 B.n539 B.n538 71.676
R767 B.n542 B.n541 71.676
R768 B.n547 B.n546 71.676
R769 B.n550 B.n549 71.676
R770 B.n555 B.n554 71.676
R771 B.n558 B.n557 71.676
R772 B.n563 B.n562 71.676
R773 B.n566 B.n565 71.676
R774 B.n572 B.n571 71.676
R775 B.n575 B.n574 71.676
R776 B.n580 B.n579 71.676
R777 B.n583 B.n582 71.676
R778 B.n588 B.n587 71.676
R779 B.n591 B.n590 71.676
R780 B.n596 B.n595 71.676
R781 B.n599 B.n598 71.676
R782 B.n604 B.n603 71.676
R783 B.n607 B.n606 71.676
R784 B.n612 B.n611 71.676
R785 B.n615 B.n614 71.676
R786 B.n620 B.n619 71.676
R787 B.n623 B.n622 71.676
R788 B.n628 B.n627 71.676
R789 B.n631 B.n630 71.676
R790 B.n636 B.n635 71.676
R791 B.n639 B.n638 71.676
R792 B.n644 B.n643 71.676
R793 B.n647 B.n646 71.676
R794 B.n351 B.n172 71.676
R795 B.n349 B.n174 71.676
R796 B.n345 B.n344 71.676
R797 B.n338 B.n176 71.676
R798 B.n337 B.n336 71.676
R799 B.n330 B.n178 71.676
R800 B.n329 B.n328 71.676
R801 B.n322 B.n180 71.676
R802 B.n321 B.n320 71.676
R803 B.n314 B.n182 71.676
R804 B.n313 B.n312 71.676
R805 B.n306 B.n184 71.676
R806 B.n305 B.n304 71.676
R807 B.n298 B.n186 71.676
R808 B.n297 B.n296 71.676
R809 B.n289 B.n188 71.676
R810 B.n288 B.n287 71.676
R811 B.n281 B.n192 71.676
R812 B.n280 B.n279 71.676
R813 B.n273 B.n194 71.676
R814 B.n272 B.n198 71.676
R815 B.n268 B.n267 71.676
R816 B.n261 B.n200 71.676
R817 B.n260 B.n259 71.676
R818 B.n253 B.n202 71.676
R819 B.n252 B.n251 71.676
R820 B.n245 B.n204 71.676
R821 B.n244 B.n243 71.676
R822 B.n237 B.n206 71.676
R823 B.n236 B.n235 71.676
R824 B.n229 B.n208 71.676
R825 B.n228 B.n227 71.676
R826 B.n221 B.n210 71.676
R827 B.n220 B.n219 71.676
R828 B.n213 B.n212 71.676
R829 B.n352 B.n351 71.676
R830 B.n346 B.n174 71.676
R831 B.n344 B.n343 71.676
R832 B.n339 B.n338 71.676
R833 B.n336 B.n335 71.676
R834 B.n331 B.n330 71.676
R835 B.n328 B.n327 71.676
R836 B.n323 B.n322 71.676
R837 B.n320 B.n319 71.676
R838 B.n315 B.n314 71.676
R839 B.n312 B.n311 71.676
R840 B.n307 B.n306 71.676
R841 B.n304 B.n303 71.676
R842 B.n299 B.n298 71.676
R843 B.n296 B.n295 71.676
R844 B.n290 B.n289 71.676
R845 B.n287 B.n286 71.676
R846 B.n282 B.n281 71.676
R847 B.n279 B.n278 71.676
R848 B.n274 B.n273 71.676
R849 B.n269 B.n198 71.676
R850 B.n267 B.n266 71.676
R851 B.n262 B.n261 71.676
R852 B.n259 B.n258 71.676
R853 B.n254 B.n253 71.676
R854 B.n251 B.n250 71.676
R855 B.n246 B.n245 71.676
R856 B.n243 B.n242 71.676
R857 B.n238 B.n237 71.676
R858 B.n235 B.n234 71.676
R859 B.n230 B.n229 71.676
R860 B.n227 B.n226 71.676
R861 B.n222 B.n221 71.676
R862 B.n219 B.n218 71.676
R863 B.n214 B.n213 71.676
R864 B.n721 B.n720 71.676
R865 B.n721 B.n2 71.676
R866 B.n85 B.n84 59.5399
R867 B.n568 B.n91 59.5399
R868 B.n197 B.n196 59.5399
R869 B.n293 B.n190 59.5399
R870 B.n84 B.n83 58.3763
R871 B.n91 B.n90 58.3763
R872 B.n196 B.n195 58.3763
R873 B.n190 B.n189 58.3763
R874 B.n357 B.n167 54.6589
R875 B.n363 B.n167 54.6589
R876 B.n363 B.n163 54.6589
R877 B.n369 B.n163 54.6589
R878 B.n369 B.n159 54.6589
R879 B.n376 B.n159 54.6589
R880 B.n376 B.n375 54.6589
R881 B.n382 B.n152 54.6589
R882 B.n388 B.n152 54.6589
R883 B.n388 B.n148 54.6589
R884 B.n394 B.n148 54.6589
R885 B.n394 B.n144 54.6589
R886 B.n400 B.n144 54.6589
R887 B.n400 B.n140 54.6589
R888 B.n406 B.n140 54.6589
R889 B.n406 B.n136 54.6589
R890 B.n413 B.n136 54.6589
R891 B.n413 B.n412 54.6589
R892 B.n419 B.n129 54.6589
R893 B.n425 B.n129 54.6589
R894 B.n425 B.n125 54.6589
R895 B.n431 B.n125 54.6589
R896 B.n431 B.n121 54.6589
R897 B.n437 B.n121 54.6589
R898 B.n437 B.n117 54.6589
R899 B.n443 B.n117 54.6589
R900 B.n450 B.n113 54.6589
R901 B.n450 B.n109 54.6589
R902 B.n456 B.n109 54.6589
R903 B.n456 B.n4 54.6589
R904 B.n719 B.n4 54.6589
R905 B.n719 B.n718 54.6589
R906 B.n718 B.n717 54.6589
R907 B.n717 B.n8 54.6589
R908 B.n12 B.n8 54.6589
R909 B.n710 B.n12 54.6589
R910 B.n710 B.n709 54.6589
R911 B.n708 B.n16 54.6589
R912 B.n702 B.n16 54.6589
R913 B.n702 B.n701 54.6589
R914 B.n701 B.n700 54.6589
R915 B.n700 B.n23 54.6589
R916 B.n694 B.n23 54.6589
R917 B.n694 B.n693 54.6589
R918 B.n693 B.n692 54.6589
R919 B.n686 B.n33 54.6589
R920 B.n686 B.n685 54.6589
R921 B.n685 B.n684 54.6589
R922 B.n684 B.n37 54.6589
R923 B.n678 B.n37 54.6589
R924 B.n678 B.n677 54.6589
R925 B.n677 B.n676 54.6589
R926 B.n676 B.n44 54.6589
R927 B.n670 B.n44 54.6589
R928 B.n670 B.n669 54.6589
R929 B.n669 B.n668 54.6589
R930 B.n662 B.n54 54.6589
R931 B.n662 B.n661 54.6589
R932 B.n661 B.n660 54.6589
R933 B.n660 B.n58 54.6589
R934 B.n654 B.n58 54.6589
R935 B.n654 B.n653 54.6589
R936 B.n653 B.n652 54.6589
R937 B.n412 B.t0 33.7601
R938 B.n33 B.t1 33.7601
R939 B.n355 B.n354 32.6249
R940 B.n359 B.n169 32.6249
R941 B.n505 B.n504 32.6249
R942 B.n650 B.n649 32.6249
R943 B.n375 B.t5 30.5449
R944 B.n54 B.t9 30.5449
R945 B.t2 B.n113 28.9373
R946 B.n709 B.t3 28.9373
R947 B.n443 B.t2 25.7221
R948 B.t3 B.n708 25.7221
R949 B.n382 B.t5 24.1145
R950 B.n668 B.t9 24.1145
R951 B.n419 B.t0 20.8993
R952 B.n692 B.t1 20.8993
R953 B B.n722 18.0485
R954 B.n355 B.n165 10.6151
R955 B.n365 B.n165 10.6151
R956 B.n366 B.n365 10.6151
R957 B.n367 B.n366 10.6151
R958 B.n367 B.n157 10.6151
R959 B.n378 B.n157 10.6151
R960 B.n379 B.n378 10.6151
R961 B.n380 B.n379 10.6151
R962 B.n380 B.n150 10.6151
R963 B.n390 B.n150 10.6151
R964 B.n391 B.n390 10.6151
R965 B.n392 B.n391 10.6151
R966 B.n392 B.n142 10.6151
R967 B.n402 B.n142 10.6151
R968 B.n403 B.n402 10.6151
R969 B.n404 B.n403 10.6151
R970 B.n404 B.n134 10.6151
R971 B.n415 B.n134 10.6151
R972 B.n416 B.n415 10.6151
R973 B.n417 B.n416 10.6151
R974 B.n417 B.n127 10.6151
R975 B.n427 B.n127 10.6151
R976 B.n428 B.n427 10.6151
R977 B.n429 B.n428 10.6151
R978 B.n429 B.n119 10.6151
R979 B.n439 B.n119 10.6151
R980 B.n440 B.n439 10.6151
R981 B.n441 B.n440 10.6151
R982 B.n441 B.n111 10.6151
R983 B.n452 B.n111 10.6151
R984 B.n453 B.n452 10.6151
R985 B.n454 B.n453 10.6151
R986 B.n454 B.n0 10.6151
R987 B.n354 B.n353 10.6151
R988 B.n353 B.n173 10.6151
R989 B.n348 B.n173 10.6151
R990 B.n348 B.n347 10.6151
R991 B.n347 B.n175 10.6151
R992 B.n342 B.n175 10.6151
R993 B.n342 B.n341 10.6151
R994 B.n341 B.n340 10.6151
R995 B.n340 B.n177 10.6151
R996 B.n334 B.n177 10.6151
R997 B.n334 B.n333 10.6151
R998 B.n333 B.n332 10.6151
R999 B.n332 B.n179 10.6151
R1000 B.n326 B.n179 10.6151
R1001 B.n326 B.n325 10.6151
R1002 B.n325 B.n324 10.6151
R1003 B.n324 B.n181 10.6151
R1004 B.n318 B.n181 10.6151
R1005 B.n318 B.n317 10.6151
R1006 B.n317 B.n316 10.6151
R1007 B.n316 B.n183 10.6151
R1008 B.n310 B.n183 10.6151
R1009 B.n310 B.n309 10.6151
R1010 B.n309 B.n308 10.6151
R1011 B.n308 B.n185 10.6151
R1012 B.n302 B.n185 10.6151
R1013 B.n302 B.n301 10.6151
R1014 B.n301 B.n300 10.6151
R1015 B.n300 B.n187 10.6151
R1016 B.n294 B.n187 10.6151
R1017 B.n292 B.n291 10.6151
R1018 B.n291 B.n191 10.6151
R1019 B.n285 B.n191 10.6151
R1020 B.n285 B.n284 10.6151
R1021 B.n284 B.n283 10.6151
R1022 B.n283 B.n193 10.6151
R1023 B.n277 B.n193 10.6151
R1024 B.n277 B.n276 10.6151
R1025 B.n276 B.n275 10.6151
R1026 B.n271 B.n270 10.6151
R1027 B.n270 B.n199 10.6151
R1028 B.n265 B.n199 10.6151
R1029 B.n265 B.n264 10.6151
R1030 B.n264 B.n263 10.6151
R1031 B.n263 B.n201 10.6151
R1032 B.n257 B.n201 10.6151
R1033 B.n257 B.n256 10.6151
R1034 B.n256 B.n255 10.6151
R1035 B.n255 B.n203 10.6151
R1036 B.n249 B.n203 10.6151
R1037 B.n249 B.n248 10.6151
R1038 B.n248 B.n247 10.6151
R1039 B.n247 B.n205 10.6151
R1040 B.n241 B.n205 10.6151
R1041 B.n241 B.n240 10.6151
R1042 B.n240 B.n239 10.6151
R1043 B.n239 B.n207 10.6151
R1044 B.n233 B.n207 10.6151
R1045 B.n233 B.n232 10.6151
R1046 B.n232 B.n231 10.6151
R1047 B.n231 B.n209 10.6151
R1048 B.n225 B.n209 10.6151
R1049 B.n225 B.n224 10.6151
R1050 B.n224 B.n223 10.6151
R1051 B.n223 B.n211 10.6151
R1052 B.n217 B.n211 10.6151
R1053 B.n217 B.n216 10.6151
R1054 B.n216 B.n215 10.6151
R1055 B.n215 B.n169 10.6151
R1056 B.n360 B.n359 10.6151
R1057 B.n361 B.n360 10.6151
R1058 B.n361 B.n161 10.6151
R1059 B.n371 B.n161 10.6151
R1060 B.n372 B.n371 10.6151
R1061 B.n373 B.n372 10.6151
R1062 B.n373 B.n154 10.6151
R1063 B.n384 B.n154 10.6151
R1064 B.n385 B.n384 10.6151
R1065 B.n386 B.n385 10.6151
R1066 B.n386 B.n146 10.6151
R1067 B.n396 B.n146 10.6151
R1068 B.n397 B.n396 10.6151
R1069 B.n398 B.n397 10.6151
R1070 B.n398 B.n138 10.6151
R1071 B.n408 B.n138 10.6151
R1072 B.n409 B.n408 10.6151
R1073 B.n410 B.n409 10.6151
R1074 B.n410 B.n131 10.6151
R1075 B.n421 B.n131 10.6151
R1076 B.n422 B.n421 10.6151
R1077 B.n423 B.n422 10.6151
R1078 B.n423 B.n123 10.6151
R1079 B.n433 B.n123 10.6151
R1080 B.n434 B.n433 10.6151
R1081 B.n435 B.n434 10.6151
R1082 B.n435 B.n115 10.6151
R1083 B.n445 B.n115 10.6151
R1084 B.n446 B.n445 10.6151
R1085 B.n448 B.n446 10.6151
R1086 B.n448 B.n447 10.6151
R1087 B.n447 B.n107 10.6151
R1088 B.n459 B.n107 10.6151
R1089 B.n460 B.n459 10.6151
R1090 B.n461 B.n460 10.6151
R1091 B.n462 B.n461 10.6151
R1092 B.n463 B.n462 10.6151
R1093 B.n466 B.n463 10.6151
R1094 B.n467 B.n466 10.6151
R1095 B.n468 B.n467 10.6151
R1096 B.n469 B.n468 10.6151
R1097 B.n471 B.n469 10.6151
R1098 B.n472 B.n471 10.6151
R1099 B.n473 B.n472 10.6151
R1100 B.n474 B.n473 10.6151
R1101 B.n476 B.n474 10.6151
R1102 B.n477 B.n476 10.6151
R1103 B.n478 B.n477 10.6151
R1104 B.n479 B.n478 10.6151
R1105 B.n481 B.n479 10.6151
R1106 B.n482 B.n481 10.6151
R1107 B.n483 B.n482 10.6151
R1108 B.n484 B.n483 10.6151
R1109 B.n486 B.n484 10.6151
R1110 B.n487 B.n486 10.6151
R1111 B.n488 B.n487 10.6151
R1112 B.n489 B.n488 10.6151
R1113 B.n491 B.n489 10.6151
R1114 B.n492 B.n491 10.6151
R1115 B.n493 B.n492 10.6151
R1116 B.n494 B.n493 10.6151
R1117 B.n496 B.n494 10.6151
R1118 B.n497 B.n496 10.6151
R1119 B.n498 B.n497 10.6151
R1120 B.n499 B.n498 10.6151
R1121 B.n501 B.n499 10.6151
R1122 B.n502 B.n501 10.6151
R1123 B.n503 B.n502 10.6151
R1124 B.n504 B.n503 10.6151
R1125 B.n714 B.n1 10.6151
R1126 B.n714 B.n713 10.6151
R1127 B.n713 B.n712 10.6151
R1128 B.n712 B.n10 10.6151
R1129 B.n706 B.n10 10.6151
R1130 B.n706 B.n705 10.6151
R1131 B.n705 B.n704 10.6151
R1132 B.n704 B.n18 10.6151
R1133 B.n698 B.n18 10.6151
R1134 B.n698 B.n697 10.6151
R1135 B.n697 B.n696 10.6151
R1136 B.n696 B.n25 10.6151
R1137 B.n690 B.n25 10.6151
R1138 B.n690 B.n689 10.6151
R1139 B.n689 B.n688 10.6151
R1140 B.n688 B.n31 10.6151
R1141 B.n682 B.n31 10.6151
R1142 B.n682 B.n681 10.6151
R1143 B.n681 B.n680 10.6151
R1144 B.n680 B.n39 10.6151
R1145 B.n674 B.n39 10.6151
R1146 B.n674 B.n673 10.6151
R1147 B.n673 B.n672 10.6151
R1148 B.n672 B.n46 10.6151
R1149 B.n666 B.n46 10.6151
R1150 B.n666 B.n665 10.6151
R1151 B.n665 B.n664 10.6151
R1152 B.n664 B.n52 10.6151
R1153 B.n658 B.n52 10.6151
R1154 B.n658 B.n657 10.6151
R1155 B.n657 B.n656 10.6151
R1156 B.n656 B.n60 10.6151
R1157 B.n650 B.n60 10.6151
R1158 B.n649 B.n648 10.6151
R1159 B.n648 B.n67 10.6151
R1160 B.n642 B.n67 10.6151
R1161 B.n642 B.n641 10.6151
R1162 B.n641 B.n640 10.6151
R1163 B.n640 B.n69 10.6151
R1164 B.n634 B.n69 10.6151
R1165 B.n634 B.n633 10.6151
R1166 B.n633 B.n632 10.6151
R1167 B.n632 B.n71 10.6151
R1168 B.n626 B.n71 10.6151
R1169 B.n626 B.n625 10.6151
R1170 B.n625 B.n624 10.6151
R1171 B.n624 B.n73 10.6151
R1172 B.n618 B.n73 10.6151
R1173 B.n618 B.n617 10.6151
R1174 B.n617 B.n616 10.6151
R1175 B.n616 B.n75 10.6151
R1176 B.n610 B.n75 10.6151
R1177 B.n610 B.n609 10.6151
R1178 B.n609 B.n608 10.6151
R1179 B.n608 B.n77 10.6151
R1180 B.n602 B.n77 10.6151
R1181 B.n602 B.n601 10.6151
R1182 B.n601 B.n600 10.6151
R1183 B.n600 B.n79 10.6151
R1184 B.n594 B.n79 10.6151
R1185 B.n594 B.n593 10.6151
R1186 B.n593 B.n592 10.6151
R1187 B.n592 B.n81 10.6151
R1188 B.n586 B.n585 10.6151
R1189 B.n585 B.n584 10.6151
R1190 B.n584 B.n86 10.6151
R1191 B.n578 B.n86 10.6151
R1192 B.n578 B.n577 10.6151
R1193 B.n577 B.n576 10.6151
R1194 B.n576 B.n88 10.6151
R1195 B.n570 B.n88 10.6151
R1196 B.n570 B.n569 10.6151
R1197 B.n567 B.n92 10.6151
R1198 B.n561 B.n92 10.6151
R1199 B.n561 B.n560 10.6151
R1200 B.n560 B.n559 10.6151
R1201 B.n559 B.n94 10.6151
R1202 B.n553 B.n94 10.6151
R1203 B.n553 B.n552 10.6151
R1204 B.n552 B.n551 10.6151
R1205 B.n551 B.n96 10.6151
R1206 B.n545 B.n96 10.6151
R1207 B.n545 B.n544 10.6151
R1208 B.n544 B.n543 10.6151
R1209 B.n543 B.n98 10.6151
R1210 B.n537 B.n98 10.6151
R1211 B.n537 B.n536 10.6151
R1212 B.n536 B.n535 10.6151
R1213 B.n535 B.n100 10.6151
R1214 B.n529 B.n100 10.6151
R1215 B.n529 B.n528 10.6151
R1216 B.n528 B.n527 10.6151
R1217 B.n527 B.n102 10.6151
R1218 B.n521 B.n102 10.6151
R1219 B.n521 B.n520 10.6151
R1220 B.n520 B.n519 10.6151
R1221 B.n519 B.n104 10.6151
R1222 B.n513 B.n104 10.6151
R1223 B.n513 B.n512 10.6151
R1224 B.n512 B.n511 10.6151
R1225 B.n511 B.n106 10.6151
R1226 B.n505 B.n106 10.6151
R1227 B.n294 B.n293 9.36635
R1228 B.n271 B.n197 9.36635
R1229 B.n85 B.n81 9.36635
R1230 B.n568 B.n567 9.36635
R1231 B.n722 B.n0 8.11757
R1232 B.n722 B.n1 8.11757
R1233 B.n293 B.n292 1.24928
R1234 B.n275 B.n197 1.24928
R1235 B.n586 B.n85 1.24928
R1236 B.n569 B.n568 1.24928
R1237 VP.n16 VP.n0 161.3
R1238 VP.n15 VP.n14 161.3
R1239 VP.n13 VP.n1 161.3
R1240 VP.n12 VP.n11 161.3
R1241 VP.n10 VP.n2 161.3
R1242 VP.n9 VP.n8 161.3
R1243 VP.n7 VP.n3 161.3
R1244 VP.n6 VP.n5 110.511
R1245 VP.n18 VP.n17 110.511
R1246 VP.n4 VP.t1 109.444
R1247 VP.n4 VP.t3 108.578
R1248 VP.n5 VP.t0 75.6277
R1249 VP.n17 VP.t2 75.6277
R1250 VP.n6 VP.n4 47.4072
R1251 VP.n11 VP.n10 40.4934
R1252 VP.n11 VP.n1 40.4934
R1253 VP.n9 VP.n3 24.4675
R1254 VP.n10 VP.n9 24.4675
R1255 VP.n15 VP.n1 24.4675
R1256 VP.n16 VP.n15 24.4675
R1257 VP.n7 VP.n6 0.278367
R1258 VP.n18 VP.n0 0.278367
R1259 VP.n5 VP.n3 0.24517
R1260 VP.n17 VP.n16 0.24517
R1261 VP.n8 VP.n7 0.189894
R1262 VP.n8 VP.n2 0.189894
R1263 VP.n12 VP.n2 0.189894
R1264 VP.n13 VP.n12 0.189894
R1265 VP.n14 VP.n13 0.189894
R1266 VP.n14 VP.n0 0.189894
R1267 VP VP.n18 0.153454
R1268 VDD1 VDD1.n1 101.347
R1269 VDD1 VDD1.n0 62.1309
R1270 VDD1.n0 VDD1.t0 2.35484
R1271 VDD1.n0 VDD1.t1 2.35484
R1272 VDD1.n1 VDD1.t2 2.35484
R1273 VDD1.n1 VDD1.t3 2.35484
R1274 VTAIL.n5 VTAIL.t6 47.7483
R1275 VTAIL.n4 VTAIL.t2 47.7483
R1276 VTAIL.n3 VTAIL.t0 47.7483
R1277 VTAIL.n6 VTAIL.t4 47.7482
R1278 VTAIL.n7 VTAIL.t1 47.7481
R1279 VTAIL.n0 VTAIL.t3 47.7481
R1280 VTAIL.n1 VTAIL.t5 47.7481
R1281 VTAIL.n2 VTAIL.t7 47.7481
R1282 VTAIL.n7 VTAIL.n6 22.2117
R1283 VTAIL.n3 VTAIL.n2 22.2117
R1284 VTAIL.n4 VTAIL.n3 2.59533
R1285 VTAIL.n6 VTAIL.n5 2.59533
R1286 VTAIL.n2 VTAIL.n1 2.59533
R1287 VTAIL VTAIL.n0 1.3561
R1288 VTAIL VTAIL.n7 1.23972
R1289 VTAIL.n5 VTAIL.n4 0.470328
R1290 VTAIL.n1 VTAIL.n0 0.470328
R1291 VN.n0 VN.t3 109.444
R1292 VN.n1 VN.t2 109.444
R1293 VN.n0 VN.t1 108.578
R1294 VN.n1 VN.t0 108.578
R1295 VN VN.n1 47.6861
R1296 VN VN.n0 3.6823
R1297 VDD2.n2 VDD2.n0 100.822
R1298 VDD2.n2 VDD2.n1 62.0727
R1299 VDD2.n1 VDD2.t3 2.35484
R1300 VDD2.n1 VDD2.t1 2.35484
R1301 VDD2.n0 VDD2.t0 2.35484
R1302 VDD2.n0 VDD2.t2 2.35484
R1303 VDD2 VDD2.n2 0.0586897
C0 VDD1 VP 3.69491f
C1 VTAIL VDD1 4.57692f
C2 VN VDD2 3.44534f
C3 VDD2 VP 0.399232f
C4 VDD2 VTAIL 4.63166f
C5 VN VP 5.58775f
C6 VN VTAIL 3.52168f
C7 VDD2 VDD1 1.03886f
C8 VTAIL VP 3.53579f
C9 VN VDD1 0.148908f
C10 VDD2 B 3.539187f
C11 VDD1 B 7.37868f
C12 VTAIL B 7.966367f
C13 VN B 10.56686f
C14 VP B 8.868258f
C15 VDD2.t0 B 0.179417f
C16 VDD2.t2 B 0.179417f
C17 VDD2.n0 B 2.10704f
C18 VDD2.t3 B 0.179417f
C19 VDD2.t1 B 0.179417f
C20 VDD2.n1 B 1.54838f
C21 VDD2.n2 B 3.39538f
C22 VN.t3 B 1.81722f
C23 VN.t1 B 1.81139f
C24 VN.n0 B 1.15831f
C25 VN.t2 B 1.81722f
C26 VN.t0 B 1.81139f
C27 VN.n1 B 2.49858f
C28 VTAIL.t3 B 1.22593f
C29 VTAIL.n0 B 0.340479f
C30 VTAIL.t5 B 1.22593f
C31 VTAIL.n1 B 0.411212f
C32 VTAIL.t7 B 1.22593f
C33 VTAIL.n2 B 1.18694f
C34 VTAIL.t0 B 1.22593f
C35 VTAIL.n3 B 1.18693f
C36 VTAIL.t2 B 1.22593f
C37 VTAIL.n4 B 0.411206f
C38 VTAIL.t6 B 1.22593f
C39 VTAIL.n5 B 0.411206f
C40 VTAIL.t4 B 1.22593f
C41 VTAIL.n6 B 1.18693f
C42 VTAIL.t1 B 1.22593f
C43 VTAIL.n7 B 1.10956f
C44 VDD1.t0 B 0.183854f
C45 VDD1.t1 B 0.183854f
C46 VDD1.n0 B 1.58711f
C47 VDD1.t2 B 0.183854f
C48 VDD1.t3 B 0.183854f
C49 VDD1.n1 B 2.18535f
C50 VP.n0 B 0.035398f
C51 VP.t2 B 1.62867f
C52 VP.n1 B 0.053362f
C53 VP.n2 B 0.026849f
C54 VP.n3 B 0.02558f
C55 VP.t3 B 1.86033f
C56 VP.t1 B 1.86632f
C57 VP.n4 B 2.55178f
C58 VP.t0 B 1.62867f
C59 VP.n5 B 0.669167f
C60 VP.n6 B 1.36284f
C61 VP.n7 B 0.035398f
C62 VP.n8 B 0.026849f
C63 VP.n9 B 0.05004f
C64 VP.n10 B 0.053362f
C65 VP.n11 B 0.021705f
C66 VP.n12 B 0.026849f
C67 VP.n13 B 0.026849f
C68 VP.n14 B 0.026849f
C69 VP.n15 B 0.05004f
C70 VP.n16 B 0.02558f
C71 VP.n17 B 0.669167f
C72 VP.n18 B 0.050097f
.ends

