* NGSPICE file created from diff_pair_sample_1457.ext - technology: sky130A

.subckt diff_pair_sample_1457 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1938_n1318# sky130_fd_pr__pfet_01v8 ad=0.6825 pd=4.28 as=0 ps=0 w=1.75 l=2.09
X1 VDD2.t1 VN.t0 VTAIL.t2 w_n1938_n1318# sky130_fd_pr__pfet_01v8 ad=0.6825 pd=4.28 as=0.6825 ps=4.28 w=1.75 l=2.09
X2 B.t8 B.t6 B.t7 w_n1938_n1318# sky130_fd_pr__pfet_01v8 ad=0.6825 pd=4.28 as=0 ps=0 w=1.75 l=2.09
X3 VDD1.t1 VP.t0 VTAIL.t1 w_n1938_n1318# sky130_fd_pr__pfet_01v8 ad=0.6825 pd=4.28 as=0.6825 ps=4.28 w=1.75 l=2.09
X4 VDD1.t0 VP.t1 VTAIL.t0 w_n1938_n1318# sky130_fd_pr__pfet_01v8 ad=0.6825 pd=4.28 as=0.6825 ps=4.28 w=1.75 l=2.09
X5 VDD2.t0 VN.t1 VTAIL.t3 w_n1938_n1318# sky130_fd_pr__pfet_01v8 ad=0.6825 pd=4.28 as=0.6825 ps=4.28 w=1.75 l=2.09
X6 B.t5 B.t3 B.t4 w_n1938_n1318# sky130_fd_pr__pfet_01v8 ad=0.6825 pd=4.28 as=0 ps=0 w=1.75 l=2.09
X7 B.t2 B.t0 B.t1 w_n1938_n1318# sky130_fd_pr__pfet_01v8 ad=0.6825 pd=4.28 as=0 ps=0 w=1.75 l=2.09
R0 B.n170 B.n169 585
R1 B.n168 B.n57 585
R2 B.n167 B.n166 585
R3 B.n165 B.n58 585
R4 B.n164 B.n163 585
R5 B.n162 B.n59 585
R6 B.n161 B.n160 585
R7 B.n159 B.n60 585
R8 B.n158 B.n157 585
R9 B.n156 B.n61 585
R10 B.n155 B.n154 585
R11 B.n153 B.n62 585
R12 B.n152 B.n151 585
R13 B.n147 B.n63 585
R14 B.n146 B.n145 585
R15 B.n144 B.n64 585
R16 B.n143 B.n142 585
R17 B.n141 B.n65 585
R18 B.n140 B.n139 585
R19 B.n138 B.n66 585
R20 B.n137 B.n136 585
R21 B.n134 B.n67 585
R22 B.n133 B.n132 585
R23 B.n131 B.n70 585
R24 B.n130 B.n129 585
R25 B.n128 B.n71 585
R26 B.n127 B.n126 585
R27 B.n125 B.n72 585
R28 B.n124 B.n123 585
R29 B.n122 B.n73 585
R30 B.n121 B.n120 585
R31 B.n119 B.n74 585
R32 B.n118 B.n117 585
R33 B.n171 B.n56 585
R34 B.n173 B.n172 585
R35 B.n174 B.n55 585
R36 B.n176 B.n175 585
R37 B.n177 B.n54 585
R38 B.n179 B.n178 585
R39 B.n180 B.n53 585
R40 B.n182 B.n181 585
R41 B.n183 B.n52 585
R42 B.n185 B.n184 585
R43 B.n186 B.n51 585
R44 B.n188 B.n187 585
R45 B.n189 B.n50 585
R46 B.n191 B.n190 585
R47 B.n192 B.n49 585
R48 B.n194 B.n193 585
R49 B.n195 B.n48 585
R50 B.n197 B.n196 585
R51 B.n198 B.n47 585
R52 B.n200 B.n199 585
R53 B.n201 B.n46 585
R54 B.n203 B.n202 585
R55 B.n204 B.n45 585
R56 B.n206 B.n205 585
R57 B.n207 B.n44 585
R58 B.n209 B.n208 585
R59 B.n210 B.n43 585
R60 B.n212 B.n211 585
R61 B.n213 B.n42 585
R62 B.n215 B.n214 585
R63 B.n216 B.n41 585
R64 B.n218 B.n217 585
R65 B.n219 B.n40 585
R66 B.n221 B.n220 585
R67 B.n222 B.n39 585
R68 B.n224 B.n223 585
R69 B.n225 B.n38 585
R70 B.n227 B.n226 585
R71 B.n228 B.n37 585
R72 B.n230 B.n229 585
R73 B.n231 B.n36 585
R74 B.n233 B.n232 585
R75 B.n234 B.n35 585
R76 B.n236 B.n235 585
R77 B.n237 B.n34 585
R78 B.n239 B.n238 585
R79 B.n290 B.n13 585
R80 B.n289 B.n288 585
R81 B.n287 B.n14 585
R82 B.n286 B.n285 585
R83 B.n284 B.n15 585
R84 B.n283 B.n282 585
R85 B.n281 B.n16 585
R86 B.n280 B.n279 585
R87 B.n278 B.n17 585
R88 B.n277 B.n276 585
R89 B.n275 B.n18 585
R90 B.n274 B.n273 585
R91 B.n271 B.n19 585
R92 B.n270 B.n269 585
R93 B.n268 B.n22 585
R94 B.n267 B.n266 585
R95 B.n265 B.n23 585
R96 B.n264 B.n263 585
R97 B.n262 B.n24 585
R98 B.n261 B.n260 585
R99 B.n259 B.n25 585
R100 B.n257 B.n256 585
R101 B.n255 B.n28 585
R102 B.n254 B.n253 585
R103 B.n252 B.n29 585
R104 B.n251 B.n250 585
R105 B.n249 B.n30 585
R106 B.n248 B.n247 585
R107 B.n246 B.n31 585
R108 B.n245 B.n244 585
R109 B.n243 B.n32 585
R110 B.n242 B.n241 585
R111 B.n240 B.n33 585
R112 B.n292 B.n291 585
R113 B.n293 B.n12 585
R114 B.n295 B.n294 585
R115 B.n296 B.n11 585
R116 B.n298 B.n297 585
R117 B.n299 B.n10 585
R118 B.n301 B.n300 585
R119 B.n302 B.n9 585
R120 B.n304 B.n303 585
R121 B.n305 B.n8 585
R122 B.n307 B.n306 585
R123 B.n308 B.n7 585
R124 B.n310 B.n309 585
R125 B.n311 B.n6 585
R126 B.n313 B.n312 585
R127 B.n314 B.n5 585
R128 B.n316 B.n315 585
R129 B.n317 B.n4 585
R130 B.n319 B.n318 585
R131 B.n320 B.n3 585
R132 B.n322 B.n321 585
R133 B.n323 B.n0 585
R134 B.n2 B.n1 585
R135 B.n86 B.n85 585
R136 B.n88 B.n87 585
R137 B.n89 B.n84 585
R138 B.n91 B.n90 585
R139 B.n92 B.n83 585
R140 B.n94 B.n93 585
R141 B.n95 B.n82 585
R142 B.n97 B.n96 585
R143 B.n98 B.n81 585
R144 B.n100 B.n99 585
R145 B.n101 B.n80 585
R146 B.n103 B.n102 585
R147 B.n104 B.n79 585
R148 B.n106 B.n105 585
R149 B.n107 B.n78 585
R150 B.n109 B.n108 585
R151 B.n110 B.n77 585
R152 B.n112 B.n111 585
R153 B.n113 B.n76 585
R154 B.n115 B.n114 585
R155 B.n116 B.n75 585
R156 B.n118 B.n75 434.841
R157 B.n171 B.n170 434.841
R158 B.n238 B.n33 434.841
R159 B.n292 B.n13 434.841
R160 B.n148 B.t7 290.423
R161 B.n26 B.t11 290.423
R162 B.n68 B.t4 290.423
R163 B.n20 B.t2 290.423
R164 B.n325 B.n324 256.663
R165 B.n149 B.t8 243.489
R166 B.n27 B.t10 243.489
R167 B.n69 B.t5 243.488
R168 B.n21 B.t1 243.488
R169 B.n324 B.n323 235.042
R170 B.n324 B.n2 235.042
R171 B.n68 B.t3 227.302
R172 B.n148 B.t6 227.302
R173 B.n26 B.t9 227.302
R174 B.n20 B.t0 227.302
R175 B.n119 B.n118 163.367
R176 B.n120 B.n119 163.367
R177 B.n120 B.n73 163.367
R178 B.n124 B.n73 163.367
R179 B.n125 B.n124 163.367
R180 B.n126 B.n125 163.367
R181 B.n126 B.n71 163.367
R182 B.n130 B.n71 163.367
R183 B.n131 B.n130 163.367
R184 B.n132 B.n131 163.367
R185 B.n132 B.n67 163.367
R186 B.n137 B.n67 163.367
R187 B.n138 B.n137 163.367
R188 B.n139 B.n138 163.367
R189 B.n139 B.n65 163.367
R190 B.n143 B.n65 163.367
R191 B.n144 B.n143 163.367
R192 B.n145 B.n144 163.367
R193 B.n145 B.n63 163.367
R194 B.n152 B.n63 163.367
R195 B.n153 B.n152 163.367
R196 B.n154 B.n153 163.367
R197 B.n154 B.n61 163.367
R198 B.n158 B.n61 163.367
R199 B.n159 B.n158 163.367
R200 B.n160 B.n159 163.367
R201 B.n160 B.n59 163.367
R202 B.n164 B.n59 163.367
R203 B.n165 B.n164 163.367
R204 B.n166 B.n165 163.367
R205 B.n166 B.n57 163.367
R206 B.n170 B.n57 163.367
R207 B.n238 B.n237 163.367
R208 B.n237 B.n236 163.367
R209 B.n236 B.n35 163.367
R210 B.n232 B.n35 163.367
R211 B.n232 B.n231 163.367
R212 B.n231 B.n230 163.367
R213 B.n230 B.n37 163.367
R214 B.n226 B.n37 163.367
R215 B.n226 B.n225 163.367
R216 B.n225 B.n224 163.367
R217 B.n224 B.n39 163.367
R218 B.n220 B.n39 163.367
R219 B.n220 B.n219 163.367
R220 B.n219 B.n218 163.367
R221 B.n218 B.n41 163.367
R222 B.n214 B.n41 163.367
R223 B.n214 B.n213 163.367
R224 B.n213 B.n212 163.367
R225 B.n212 B.n43 163.367
R226 B.n208 B.n43 163.367
R227 B.n208 B.n207 163.367
R228 B.n207 B.n206 163.367
R229 B.n206 B.n45 163.367
R230 B.n202 B.n45 163.367
R231 B.n202 B.n201 163.367
R232 B.n201 B.n200 163.367
R233 B.n200 B.n47 163.367
R234 B.n196 B.n47 163.367
R235 B.n196 B.n195 163.367
R236 B.n195 B.n194 163.367
R237 B.n194 B.n49 163.367
R238 B.n190 B.n49 163.367
R239 B.n190 B.n189 163.367
R240 B.n189 B.n188 163.367
R241 B.n188 B.n51 163.367
R242 B.n184 B.n51 163.367
R243 B.n184 B.n183 163.367
R244 B.n183 B.n182 163.367
R245 B.n182 B.n53 163.367
R246 B.n178 B.n53 163.367
R247 B.n178 B.n177 163.367
R248 B.n177 B.n176 163.367
R249 B.n176 B.n55 163.367
R250 B.n172 B.n55 163.367
R251 B.n172 B.n171 163.367
R252 B.n288 B.n13 163.367
R253 B.n288 B.n287 163.367
R254 B.n287 B.n286 163.367
R255 B.n286 B.n15 163.367
R256 B.n282 B.n15 163.367
R257 B.n282 B.n281 163.367
R258 B.n281 B.n280 163.367
R259 B.n280 B.n17 163.367
R260 B.n276 B.n17 163.367
R261 B.n276 B.n275 163.367
R262 B.n275 B.n274 163.367
R263 B.n274 B.n19 163.367
R264 B.n269 B.n19 163.367
R265 B.n269 B.n268 163.367
R266 B.n268 B.n267 163.367
R267 B.n267 B.n23 163.367
R268 B.n263 B.n23 163.367
R269 B.n263 B.n262 163.367
R270 B.n262 B.n261 163.367
R271 B.n261 B.n25 163.367
R272 B.n256 B.n25 163.367
R273 B.n256 B.n255 163.367
R274 B.n255 B.n254 163.367
R275 B.n254 B.n29 163.367
R276 B.n250 B.n29 163.367
R277 B.n250 B.n249 163.367
R278 B.n249 B.n248 163.367
R279 B.n248 B.n31 163.367
R280 B.n244 B.n31 163.367
R281 B.n244 B.n243 163.367
R282 B.n243 B.n242 163.367
R283 B.n242 B.n33 163.367
R284 B.n293 B.n292 163.367
R285 B.n294 B.n293 163.367
R286 B.n294 B.n11 163.367
R287 B.n298 B.n11 163.367
R288 B.n299 B.n298 163.367
R289 B.n300 B.n299 163.367
R290 B.n300 B.n9 163.367
R291 B.n304 B.n9 163.367
R292 B.n305 B.n304 163.367
R293 B.n306 B.n305 163.367
R294 B.n306 B.n7 163.367
R295 B.n310 B.n7 163.367
R296 B.n311 B.n310 163.367
R297 B.n312 B.n311 163.367
R298 B.n312 B.n5 163.367
R299 B.n316 B.n5 163.367
R300 B.n317 B.n316 163.367
R301 B.n318 B.n317 163.367
R302 B.n318 B.n3 163.367
R303 B.n322 B.n3 163.367
R304 B.n323 B.n322 163.367
R305 B.n85 B.n2 163.367
R306 B.n88 B.n85 163.367
R307 B.n89 B.n88 163.367
R308 B.n90 B.n89 163.367
R309 B.n90 B.n83 163.367
R310 B.n94 B.n83 163.367
R311 B.n95 B.n94 163.367
R312 B.n96 B.n95 163.367
R313 B.n96 B.n81 163.367
R314 B.n100 B.n81 163.367
R315 B.n101 B.n100 163.367
R316 B.n102 B.n101 163.367
R317 B.n102 B.n79 163.367
R318 B.n106 B.n79 163.367
R319 B.n107 B.n106 163.367
R320 B.n108 B.n107 163.367
R321 B.n108 B.n77 163.367
R322 B.n112 B.n77 163.367
R323 B.n113 B.n112 163.367
R324 B.n114 B.n113 163.367
R325 B.n114 B.n75 163.367
R326 B.n135 B.n69 59.5399
R327 B.n150 B.n149 59.5399
R328 B.n258 B.n27 59.5399
R329 B.n272 B.n21 59.5399
R330 B.n69 B.n68 46.9338
R331 B.n149 B.n148 46.9338
R332 B.n27 B.n26 46.9338
R333 B.n21 B.n20 46.9338
R334 B.n169 B.n56 28.2542
R335 B.n291 B.n290 28.2542
R336 B.n240 B.n239 28.2542
R337 B.n117 B.n116 28.2542
R338 B B.n325 18.0485
R339 B.n291 B.n12 10.6151
R340 B.n295 B.n12 10.6151
R341 B.n296 B.n295 10.6151
R342 B.n297 B.n296 10.6151
R343 B.n297 B.n10 10.6151
R344 B.n301 B.n10 10.6151
R345 B.n302 B.n301 10.6151
R346 B.n303 B.n302 10.6151
R347 B.n303 B.n8 10.6151
R348 B.n307 B.n8 10.6151
R349 B.n308 B.n307 10.6151
R350 B.n309 B.n308 10.6151
R351 B.n309 B.n6 10.6151
R352 B.n313 B.n6 10.6151
R353 B.n314 B.n313 10.6151
R354 B.n315 B.n314 10.6151
R355 B.n315 B.n4 10.6151
R356 B.n319 B.n4 10.6151
R357 B.n320 B.n319 10.6151
R358 B.n321 B.n320 10.6151
R359 B.n321 B.n0 10.6151
R360 B.n290 B.n289 10.6151
R361 B.n289 B.n14 10.6151
R362 B.n285 B.n14 10.6151
R363 B.n285 B.n284 10.6151
R364 B.n284 B.n283 10.6151
R365 B.n283 B.n16 10.6151
R366 B.n279 B.n16 10.6151
R367 B.n279 B.n278 10.6151
R368 B.n278 B.n277 10.6151
R369 B.n277 B.n18 10.6151
R370 B.n273 B.n18 10.6151
R371 B.n271 B.n270 10.6151
R372 B.n270 B.n22 10.6151
R373 B.n266 B.n22 10.6151
R374 B.n266 B.n265 10.6151
R375 B.n265 B.n264 10.6151
R376 B.n264 B.n24 10.6151
R377 B.n260 B.n24 10.6151
R378 B.n260 B.n259 10.6151
R379 B.n257 B.n28 10.6151
R380 B.n253 B.n28 10.6151
R381 B.n253 B.n252 10.6151
R382 B.n252 B.n251 10.6151
R383 B.n251 B.n30 10.6151
R384 B.n247 B.n30 10.6151
R385 B.n247 B.n246 10.6151
R386 B.n246 B.n245 10.6151
R387 B.n245 B.n32 10.6151
R388 B.n241 B.n32 10.6151
R389 B.n241 B.n240 10.6151
R390 B.n239 B.n34 10.6151
R391 B.n235 B.n34 10.6151
R392 B.n235 B.n234 10.6151
R393 B.n234 B.n233 10.6151
R394 B.n233 B.n36 10.6151
R395 B.n229 B.n36 10.6151
R396 B.n229 B.n228 10.6151
R397 B.n228 B.n227 10.6151
R398 B.n227 B.n38 10.6151
R399 B.n223 B.n38 10.6151
R400 B.n223 B.n222 10.6151
R401 B.n222 B.n221 10.6151
R402 B.n221 B.n40 10.6151
R403 B.n217 B.n40 10.6151
R404 B.n217 B.n216 10.6151
R405 B.n216 B.n215 10.6151
R406 B.n215 B.n42 10.6151
R407 B.n211 B.n42 10.6151
R408 B.n211 B.n210 10.6151
R409 B.n210 B.n209 10.6151
R410 B.n209 B.n44 10.6151
R411 B.n205 B.n44 10.6151
R412 B.n205 B.n204 10.6151
R413 B.n204 B.n203 10.6151
R414 B.n203 B.n46 10.6151
R415 B.n199 B.n46 10.6151
R416 B.n199 B.n198 10.6151
R417 B.n198 B.n197 10.6151
R418 B.n197 B.n48 10.6151
R419 B.n193 B.n48 10.6151
R420 B.n193 B.n192 10.6151
R421 B.n192 B.n191 10.6151
R422 B.n191 B.n50 10.6151
R423 B.n187 B.n50 10.6151
R424 B.n187 B.n186 10.6151
R425 B.n186 B.n185 10.6151
R426 B.n185 B.n52 10.6151
R427 B.n181 B.n52 10.6151
R428 B.n181 B.n180 10.6151
R429 B.n180 B.n179 10.6151
R430 B.n179 B.n54 10.6151
R431 B.n175 B.n54 10.6151
R432 B.n175 B.n174 10.6151
R433 B.n174 B.n173 10.6151
R434 B.n173 B.n56 10.6151
R435 B.n86 B.n1 10.6151
R436 B.n87 B.n86 10.6151
R437 B.n87 B.n84 10.6151
R438 B.n91 B.n84 10.6151
R439 B.n92 B.n91 10.6151
R440 B.n93 B.n92 10.6151
R441 B.n93 B.n82 10.6151
R442 B.n97 B.n82 10.6151
R443 B.n98 B.n97 10.6151
R444 B.n99 B.n98 10.6151
R445 B.n99 B.n80 10.6151
R446 B.n103 B.n80 10.6151
R447 B.n104 B.n103 10.6151
R448 B.n105 B.n104 10.6151
R449 B.n105 B.n78 10.6151
R450 B.n109 B.n78 10.6151
R451 B.n110 B.n109 10.6151
R452 B.n111 B.n110 10.6151
R453 B.n111 B.n76 10.6151
R454 B.n115 B.n76 10.6151
R455 B.n116 B.n115 10.6151
R456 B.n117 B.n74 10.6151
R457 B.n121 B.n74 10.6151
R458 B.n122 B.n121 10.6151
R459 B.n123 B.n122 10.6151
R460 B.n123 B.n72 10.6151
R461 B.n127 B.n72 10.6151
R462 B.n128 B.n127 10.6151
R463 B.n129 B.n128 10.6151
R464 B.n129 B.n70 10.6151
R465 B.n133 B.n70 10.6151
R466 B.n134 B.n133 10.6151
R467 B.n136 B.n66 10.6151
R468 B.n140 B.n66 10.6151
R469 B.n141 B.n140 10.6151
R470 B.n142 B.n141 10.6151
R471 B.n142 B.n64 10.6151
R472 B.n146 B.n64 10.6151
R473 B.n147 B.n146 10.6151
R474 B.n151 B.n147 10.6151
R475 B.n155 B.n62 10.6151
R476 B.n156 B.n155 10.6151
R477 B.n157 B.n156 10.6151
R478 B.n157 B.n60 10.6151
R479 B.n161 B.n60 10.6151
R480 B.n162 B.n161 10.6151
R481 B.n163 B.n162 10.6151
R482 B.n163 B.n58 10.6151
R483 B.n167 B.n58 10.6151
R484 B.n168 B.n167 10.6151
R485 B.n169 B.n168 10.6151
R486 B.n325 B.n0 8.11757
R487 B.n325 B.n1 8.11757
R488 B.n272 B.n271 6.5566
R489 B.n259 B.n258 6.5566
R490 B.n136 B.n135 6.5566
R491 B.n151 B.n150 6.5566
R492 B.n273 B.n272 4.05904
R493 B.n258 B.n257 4.05904
R494 B.n135 B.n134 4.05904
R495 B.n150 B.n62 4.05904
R496 VN VN.t1 114.77
R497 VN VN.t0 79.2819
R498 VTAIL.n26 VTAIL.n24 756.745
R499 VTAIL.n2 VTAIL.n0 756.745
R500 VTAIL.n18 VTAIL.n16 756.745
R501 VTAIL.n10 VTAIL.n8 756.745
R502 VTAIL.n27 VTAIL.n26 585
R503 VTAIL.n3 VTAIL.n2 585
R504 VTAIL.n19 VTAIL.n18 585
R505 VTAIL.n11 VTAIL.n10 585
R506 VTAIL.t2 VTAIL.n25 415.613
R507 VTAIL.t1 VTAIL.n1 415.613
R508 VTAIL.t0 VTAIL.n17 415.613
R509 VTAIL.t3 VTAIL.n9 415.613
R510 VTAIL.n26 VTAIL.t2 85.8723
R511 VTAIL.n2 VTAIL.t1 85.8723
R512 VTAIL.n18 VTAIL.t0 85.8723
R513 VTAIL.n10 VTAIL.t3 85.8723
R514 VTAIL.n31 VTAIL.n30 33.5429
R515 VTAIL.n7 VTAIL.n6 33.5429
R516 VTAIL.n23 VTAIL.n22 33.5429
R517 VTAIL.n15 VTAIL.n14 33.5429
R518 VTAIL.n15 VTAIL.n7 18.0479
R519 VTAIL.n31 VTAIL.n23 15.9617
R520 VTAIL.n27 VTAIL.n25 14.9339
R521 VTAIL.n3 VTAIL.n1 14.9339
R522 VTAIL.n19 VTAIL.n17 14.9339
R523 VTAIL.n11 VTAIL.n9 14.9339
R524 VTAIL.n28 VTAIL.n24 12.8005
R525 VTAIL.n4 VTAIL.n0 12.8005
R526 VTAIL.n20 VTAIL.n16 12.8005
R527 VTAIL.n12 VTAIL.n8 12.8005
R528 VTAIL.n30 VTAIL.n29 9.45567
R529 VTAIL.n6 VTAIL.n5 9.45567
R530 VTAIL.n22 VTAIL.n21 9.45567
R531 VTAIL.n14 VTAIL.n13 9.45567
R532 VTAIL.n29 VTAIL.n28 9.3005
R533 VTAIL.n5 VTAIL.n4 9.3005
R534 VTAIL.n21 VTAIL.n20 9.3005
R535 VTAIL.n13 VTAIL.n12 9.3005
R536 VTAIL.n29 VTAIL.n25 5.44463
R537 VTAIL.n5 VTAIL.n1 5.44463
R538 VTAIL.n21 VTAIL.n17 5.44463
R539 VTAIL.n13 VTAIL.n9 5.44463
R540 VTAIL.n23 VTAIL.n15 1.51343
R541 VTAIL.n30 VTAIL.n24 1.16414
R542 VTAIL.n6 VTAIL.n0 1.16414
R543 VTAIL.n22 VTAIL.n16 1.16414
R544 VTAIL.n14 VTAIL.n8 1.16414
R545 VTAIL VTAIL.n7 1.05007
R546 VTAIL VTAIL.n31 0.463862
R547 VTAIL.n28 VTAIL.n27 0.388379
R548 VTAIL.n4 VTAIL.n3 0.388379
R549 VTAIL.n20 VTAIL.n19 0.388379
R550 VTAIL.n12 VTAIL.n11 0.388379
R551 VDD2.n9 VDD2.n7 756.745
R552 VDD2.n2 VDD2.n0 756.745
R553 VDD2.n10 VDD2.n9 585
R554 VDD2.n3 VDD2.n2 585
R555 VDD2.t1 VDD2.n1 415.613
R556 VDD2.t0 VDD2.n8 415.613
R557 VDD2.n9 VDD2.t0 85.8723
R558 VDD2.n2 VDD2.t1 85.8723
R559 VDD2.n14 VDD2.n6 79.5622
R560 VDD2.n14 VDD2.n13 50.2217
R561 VDD2.n10 VDD2.n8 14.9339
R562 VDD2.n3 VDD2.n1 14.9339
R563 VDD2.n11 VDD2.n7 12.8005
R564 VDD2.n4 VDD2.n0 12.8005
R565 VDD2.n13 VDD2.n12 9.45567
R566 VDD2.n6 VDD2.n5 9.45567
R567 VDD2.n12 VDD2.n11 9.3005
R568 VDD2.n5 VDD2.n4 9.3005
R569 VDD2.n12 VDD2.n8 5.44463
R570 VDD2.n5 VDD2.n1 5.44463
R571 VDD2.n13 VDD2.n7 1.16414
R572 VDD2.n6 VDD2.n0 1.16414
R573 VDD2 VDD2.n14 0.580241
R574 VDD2.n11 VDD2.n10 0.388379
R575 VDD2.n4 VDD2.n3 0.388379
R576 VP.n0 VP.t1 114.579
R577 VP.n0 VP.t0 79.0407
R578 VP VP.n0 0.241678
R579 VDD1.n2 VDD1.n0 756.745
R580 VDD1.n9 VDD1.n7 756.745
R581 VDD1.n3 VDD1.n2 585
R582 VDD1.n10 VDD1.n9 585
R583 VDD1.t1 VDD1.n8 415.613
R584 VDD1.t0 VDD1.n1 415.613
R585 VDD1.n2 VDD1.t0 85.8723
R586 VDD1.n9 VDD1.t1 85.8723
R587 VDD1 VDD1.n13 80.6086
R588 VDD1 VDD1.n6 50.8015
R589 VDD1.n3 VDD1.n1 14.9339
R590 VDD1.n10 VDD1.n8 14.9339
R591 VDD1.n4 VDD1.n0 12.8005
R592 VDD1.n11 VDD1.n7 12.8005
R593 VDD1.n6 VDD1.n5 9.45567
R594 VDD1.n13 VDD1.n12 9.45567
R595 VDD1.n5 VDD1.n4 9.3005
R596 VDD1.n12 VDD1.n11 9.3005
R597 VDD1.n5 VDD1.n1 5.44463
R598 VDD1.n12 VDD1.n8 5.44463
R599 VDD1.n6 VDD1.n0 1.16414
R600 VDD1.n13 VDD1.n7 1.16414
R601 VDD1.n4 VDD1.n3 0.388379
R602 VDD1.n11 VDD1.n10 0.388379
C0 VDD1 w_n1938_n1318# 0.997372f
C1 VTAIL VN 0.848638f
C2 VDD2 B 0.86138f
C3 VTAIL w_n1938_n1318# 1.22805f
C4 VDD1 B 0.835475f
C5 VTAIL B 1.14153f
C6 VDD2 VP 0.318181f
C7 VDD1 VP 0.768507f
C8 VTAIL VP 0.862778f
C9 VN w_n1938_n1318# 2.39812f
C10 VN B 0.805427f
C11 w_n1938_n1318# B 5.404089f
C12 VDD2 VDD1 0.612442f
C13 VN VP 3.32223f
C14 VTAIL VDD2 2.24473f
C15 VP w_n1938_n1318# 2.63844f
C16 VTAIL VDD1 2.19526f
C17 VP B 1.20658f
C18 VN VDD2 0.606429f
C19 VDD2 w_n1938_n1318# 1.01635f
C20 VN VDD1 0.154556f
C21 VDD2 VSUBS 0.496747f
C22 VDD1 VSUBS 2.003811f
C23 VTAIL VSUBS 0.32923f
C24 VN VSUBS 5.10471f
C25 VP VSUBS 1.050852f
C26 B VSUBS 2.512051f
C27 w_n1938_n1318# VSUBS 32.674698f
C28 VDD1.n0 VSUBS 0.017058f
C29 VDD1.n1 VSUBS 0.045276f
C30 VDD1.t0 VSUBS 0.043795f
C31 VDD1.n2 VSUBS 0.041663f
C32 VDD1.n3 VSUBS 0.011253f
C33 VDD1.n4 VSUBS 0.008964f
C34 VDD1.n5 VSUBS 0.095563f
C35 VDD1.n6 VSUBS 0.03571f
C36 VDD1.n7 VSUBS 0.017058f
C37 VDD1.n8 VSUBS 0.045276f
C38 VDD1.t1 VSUBS 0.043795f
C39 VDD1.n9 VSUBS 0.041663f
C40 VDD1.n10 VSUBS 0.011253f
C41 VDD1.n11 VSUBS 0.008964f
C42 VDD1.n12 VSUBS 0.095563f
C43 VDD1.n13 VSUBS 0.273743f
C44 VP.t1 VSUBS 1.52914f
C45 VP.t0 VSUBS 0.903056f
C46 VP.n0 VSUBS 3.36894f
C47 VDD2.n0 VSUBS 0.017549f
C48 VDD2.n1 VSUBS 0.046581f
C49 VDD2.t1 VSUBS 0.045057f
C50 VDD2.n2 VSUBS 0.042863f
C51 VDD2.n3 VSUBS 0.011577f
C52 VDD2.n4 VSUBS 0.009222f
C53 VDD2.n5 VSUBS 0.098316f
C54 VDD2.n6 VSUBS 0.257823f
C55 VDD2.n7 VSUBS 0.017549f
C56 VDD2.n8 VSUBS 0.046581f
C57 VDD2.t0 VSUBS 0.045057f
C58 VDD2.n9 VSUBS 0.042863f
C59 VDD2.n10 VSUBS 0.011577f
C60 VDD2.n11 VSUBS 0.009222f
C61 VDD2.n12 VSUBS 0.098316f
C62 VDD2.n13 VSUBS 0.035985f
C63 VDD2.n14 VSUBS 1.27364f
C64 VTAIL.n0 VSUBS 0.021833f
C65 VTAIL.n1 VSUBS 0.057952f
C66 VTAIL.t1 VSUBS 0.056056f
C67 VTAIL.n2 VSUBS 0.053327f
C68 VTAIL.n3 VSUBS 0.014403f
C69 VTAIL.n4 VSUBS 0.011473f
C70 VTAIL.n5 VSUBS 0.122316f
C71 VTAIL.n6 VSUBS 0.030042f
C72 VTAIL.n7 VSUBS 0.772484f
C73 VTAIL.n8 VSUBS 0.021833f
C74 VTAIL.n9 VSUBS 0.057952f
C75 VTAIL.t3 VSUBS 0.056056f
C76 VTAIL.n10 VSUBS 0.053327f
C77 VTAIL.n11 VSUBS 0.014403f
C78 VTAIL.n12 VSUBS 0.011473f
C79 VTAIL.n13 VSUBS 0.122316f
C80 VTAIL.n14 VSUBS 0.030042f
C81 VTAIL.n15 VSUBS 0.804363f
C82 VTAIL.n16 VSUBS 0.021833f
C83 VTAIL.n17 VSUBS 0.057952f
C84 VTAIL.t0 VSUBS 0.056056f
C85 VTAIL.n18 VSUBS 0.053327f
C86 VTAIL.n19 VSUBS 0.014403f
C87 VTAIL.n20 VSUBS 0.011473f
C88 VTAIL.n21 VSUBS 0.122316f
C89 VTAIL.n22 VSUBS 0.030042f
C90 VTAIL.n23 VSUBS 0.660833f
C91 VTAIL.n24 VSUBS 0.021833f
C92 VTAIL.n25 VSUBS 0.057952f
C93 VTAIL.t2 VSUBS 0.056056f
C94 VTAIL.n26 VSUBS 0.053327f
C95 VTAIL.n27 VSUBS 0.014403f
C96 VTAIL.n28 VSUBS 0.011473f
C97 VTAIL.n29 VSUBS 0.122316f
C98 VTAIL.n30 VSUBS 0.030042f
C99 VTAIL.n31 VSUBS 0.588624f
C100 VN.t0 VSUBS 0.861781f
C101 VN.t1 VSUBS 1.46817f
C102 B.n0 VSUBS 0.008508f
C103 B.n1 VSUBS 0.008508f
C104 B.n2 VSUBS 0.012583f
C105 B.n3 VSUBS 0.009642f
C106 B.n4 VSUBS 0.009642f
C107 B.n5 VSUBS 0.009642f
C108 B.n6 VSUBS 0.009642f
C109 B.n7 VSUBS 0.009642f
C110 B.n8 VSUBS 0.009642f
C111 B.n9 VSUBS 0.009642f
C112 B.n10 VSUBS 0.009642f
C113 B.n11 VSUBS 0.009642f
C114 B.n12 VSUBS 0.009642f
C115 B.n13 VSUBS 0.021283f
C116 B.n14 VSUBS 0.009642f
C117 B.n15 VSUBS 0.009642f
C118 B.n16 VSUBS 0.009642f
C119 B.n17 VSUBS 0.009642f
C120 B.n18 VSUBS 0.009642f
C121 B.n19 VSUBS 0.009642f
C122 B.t1 VSUBS 0.0408f
C123 B.t2 VSUBS 0.052053f
C124 B.t0 VSUBS 0.248616f
C125 B.n20 VSUBS 0.097902f
C126 B.n21 VSUBS 0.083387f
C127 B.n22 VSUBS 0.009642f
C128 B.n23 VSUBS 0.009642f
C129 B.n24 VSUBS 0.009642f
C130 B.n25 VSUBS 0.009642f
C131 B.t10 VSUBS 0.0408f
C132 B.t11 VSUBS 0.052053f
C133 B.t9 VSUBS 0.248616f
C134 B.n26 VSUBS 0.097902f
C135 B.n27 VSUBS 0.083387f
C136 B.n28 VSUBS 0.009642f
C137 B.n29 VSUBS 0.009642f
C138 B.n30 VSUBS 0.009642f
C139 B.n31 VSUBS 0.009642f
C140 B.n32 VSUBS 0.009642f
C141 B.n33 VSUBS 0.021283f
C142 B.n34 VSUBS 0.009642f
C143 B.n35 VSUBS 0.009642f
C144 B.n36 VSUBS 0.009642f
C145 B.n37 VSUBS 0.009642f
C146 B.n38 VSUBS 0.009642f
C147 B.n39 VSUBS 0.009642f
C148 B.n40 VSUBS 0.009642f
C149 B.n41 VSUBS 0.009642f
C150 B.n42 VSUBS 0.009642f
C151 B.n43 VSUBS 0.009642f
C152 B.n44 VSUBS 0.009642f
C153 B.n45 VSUBS 0.009642f
C154 B.n46 VSUBS 0.009642f
C155 B.n47 VSUBS 0.009642f
C156 B.n48 VSUBS 0.009642f
C157 B.n49 VSUBS 0.009642f
C158 B.n50 VSUBS 0.009642f
C159 B.n51 VSUBS 0.009642f
C160 B.n52 VSUBS 0.009642f
C161 B.n53 VSUBS 0.009642f
C162 B.n54 VSUBS 0.009642f
C163 B.n55 VSUBS 0.009642f
C164 B.n56 VSUBS 0.021155f
C165 B.n57 VSUBS 0.009642f
C166 B.n58 VSUBS 0.009642f
C167 B.n59 VSUBS 0.009642f
C168 B.n60 VSUBS 0.009642f
C169 B.n61 VSUBS 0.009642f
C170 B.n62 VSUBS 0.006664f
C171 B.n63 VSUBS 0.009642f
C172 B.n64 VSUBS 0.009642f
C173 B.n65 VSUBS 0.009642f
C174 B.n66 VSUBS 0.009642f
C175 B.n67 VSUBS 0.009642f
C176 B.t5 VSUBS 0.0408f
C177 B.t4 VSUBS 0.052053f
C178 B.t3 VSUBS 0.248616f
C179 B.n68 VSUBS 0.097902f
C180 B.n69 VSUBS 0.083387f
C181 B.n70 VSUBS 0.009642f
C182 B.n71 VSUBS 0.009642f
C183 B.n72 VSUBS 0.009642f
C184 B.n73 VSUBS 0.009642f
C185 B.n74 VSUBS 0.009642f
C186 B.n75 VSUBS 0.019838f
C187 B.n76 VSUBS 0.009642f
C188 B.n77 VSUBS 0.009642f
C189 B.n78 VSUBS 0.009642f
C190 B.n79 VSUBS 0.009642f
C191 B.n80 VSUBS 0.009642f
C192 B.n81 VSUBS 0.009642f
C193 B.n82 VSUBS 0.009642f
C194 B.n83 VSUBS 0.009642f
C195 B.n84 VSUBS 0.009642f
C196 B.n85 VSUBS 0.009642f
C197 B.n86 VSUBS 0.009642f
C198 B.n87 VSUBS 0.009642f
C199 B.n88 VSUBS 0.009642f
C200 B.n89 VSUBS 0.009642f
C201 B.n90 VSUBS 0.009642f
C202 B.n91 VSUBS 0.009642f
C203 B.n92 VSUBS 0.009642f
C204 B.n93 VSUBS 0.009642f
C205 B.n94 VSUBS 0.009642f
C206 B.n95 VSUBS 0.009642f
C207 B.n96 VSUBS 0.009642f
C208 B.n97 VSUBS 0.009642f
C209 B.n98 VSUBS 0.009642f
C210 B.n99 VSUBS 0.009642f
C211 B.n100 VSUBS 0.009642f
C212 B.n101 VSUBS 0.009642f
C213 B.n102 VSUBS 0.009642f
C214 B.n103 VSUBS 0.009642f
C215 B.n104 VSUBS 0.009642f
C216 B.n105 VSUBS 0.009642f
C217 B.n106 VSUBS 0.009642f
C218 B.n107 VSUBS 0.009642f
C219 B.n108 VSUBS 0.009642f
C220 B.n109 VSUBS 0.009642f
C221 B.n110 VSUBS 0.009642f
C222 B.n111 VSUBS 0.009642f
C223 B.n112 VSUBS 0.009642f
C224 B.n113 VSUBS 0.009642f
C225 B.n114 VSUBS 0.009642f
C226 B.n115 VSUBS 0.009642f
C227 B.n116 VSUBS 0.019838f
C228 B.n117 VSUBS 0.021283f
C229 B.n118 VSUBS 0.021283f
C230 B.n119 VSUBS 0.009642f
C231 B.n120 VSUBS 0.009642f
C232 B.n121 VSUBS 0.009642f
C233 B.n122 VSUBS 0.009642f
C234 B.n123 VSUBS 0.009642f
C235 B.n124 VSUBS 0.009642f
C236 B.n125 VSUBS 0.009642f
C237 B.n126 VSUBS 0.009642f
C238 B.n127 VSUBS 0.009642f
C239 B.n128 VSUBS 0.009642f
C240 B.n129 VSUBS 0.009642f
C241 B.n130 VSUBS 0.009642f
C242 B.n131 VSUBS 0.009642f
C243 B.n132 VSUBS 0.009642f
C244 B.n133 VSUBS 0.009642f
C245 B.n134 VSUBS 0.006664f
C246 B.n135 VSUBS 0.02234f
C247 B.n136 VSUBS 0.007799f
C248 B.n137 VSUBS 0.009642f
C249 B.n138 VSUBS 0.009642f
C250 B.n139 VSUBS 0.009642f
C251 B.n140 VSUBS 0.009642f
C252 B.n141 VSUBS 0.009642f
C253 B.n142 VSUBS 0.009642f
C254 B.n143 VSUBS 0.009642f
C255 B.n144 VSUBS 0.009642f
C256 B.n145 VSUBS 0.009642f
C257 B.n146 VSUBS 0.009642f
C258 B.n147 VSUBS 0.009642f
C259 B.t8 VSUBS 0.0408f
C260 B.t7 VSUBS 0.052053f
C261 B.t6 VSUBS 0.248616f
C262 B.n148 VSUBS 0.097902f
C263 B.n149 VSUBS 0.083387f
C264 B.n150 VSUBS 0.02234f
C265 B.n151 VSUBS 0.007799f
C266 B.n152 VSUBS 0.009642f
C267 B.n153 VSUBS 0.009642f
C268 B.n154 VSUBS 0.009642f
C269 B.n155 VSUBS 0.009642f
C270 B.n156 VSUBS 0.009642f
C271 B.n157 VSUBS 0.009642f
C272 B.n158 VSUBS 0.009642f
C273 B.n159 VSUBS 0.009642f
C274 B.n160 VSUBS 0.009642f
C275 B.n161 VSUBS 0.009642f
C276 B.n162 VSUBS 0.009642f
C277 B.n163 VSUBS 0.009642f
C278 B.n164 VSUBS 0.009642f
C279 B.n165 VSUBS 0.009642f
C280 B.n166 VSUBS 0.009642f
C281 B.n167 VSUBS 0.009642f
C282 B.n168 VSUBS 0.009642f
C283 B.n169 VSUBS 0.019966f
C284 B.n170 VSUBS 0.021283f
C285 B.n171 VSUBS 0.019838f
C286 B.n172 VSUBS 0.009642f
C287 B.n173 VSUBS 0.009642f
C288 B.n174 VSUBS 0.009642f
C289 B.n175 VSUBS 0.009642f
C290 B.n176 VSUBS 0.009642f
C291 B.n177 VSUBS 0.009642f
C292 B.n178 VSUBS 0.009642f
C293 B.n179 VSUBS 0.009642f
C294 B.n180 VSUBS 0.009642f
C295 B.n181 VSUBS 0.009642f
C296 B.n182 VSUBS 0.009642f
C297 B.n183 VSUBS 0.009642f
C298 B.n184 VSUBS 0.009642f
C299 B.n185 VSUBS 0.009642f
C300 B.n186 VSUBS 0.009642f
C301 B.n187 VSUBS 0.009642f
C302 B.n188 VSUBS 0.009642f
C303 B.n189 VSUBS 0.009642f
C304 B.n190 VSUBS 0.009642f
C305 B.n191 VSUBS 0.009642f
C306 B.n192 VSUBS 0.009642f
C307 B.n193 VSUBS 0.009642f
C308 B.n194 VSUBS 0.009642f
C309 B.n195 VSUBS 0.009642f
C310 B.n196 VSUBS 0.009642f
C311 B.n197 VSUBS 0.009642f
C312 B.n198 VSUBS 0.009642f
C313 B.n199 VSUBS 0.009642f
C314 B.n200 VSUBS 0.009642f
C315 B.n201 VSUBS 0.009642f
C316 B.n202 VSUBS 0.009642f
C317 B.n203 VSUBS 0.009642f
C318 B.n204 VSUBS 0.009642f
C319 B.n205 VSUBS 0.009642f
C320 B.n206 VSUBS 0.009642f
C321 B.n207 VSUBS 0.009642f
C322 B.n208 VSUBS 0.009642f
C323 B.n209 VSUBS 0.009642f
C324 B.n210 VSUBS 0.009642f
C325 B.n211 VSUBS 0.009642f
C326 B.n212 VSUBS 0.009642f
C327 B.n213 VSUBS 0.009642f
C328 B.n214 VSUBS 0.009642f
C329 B.n215 VSUBS 0.009642f
C330 B.n216 VSUBS 0.009642f
C331 B.n217 VSUBS 0.009642f
C332 B.n218 VSUBS 0.009642f
C333 B.n219 VSUBS 0.009642f
C334 B.n220 VSUBS 0.009642f
C335 B.n221 VSUBS 0.009642f
C336 B.n222 VSUBS 0.009642f
C337 B.n223 VSUBS 0.009642f
C338 B.n224 VSUBS 0.009642f
C339 B.n225 VSUBS 0.009642f
C340 B.n226 VSUBS 0.009642f
C341 B.n227 VSUBS 0.009642f
C342 B.n228 VSUBS 0.009642f
C343 B.n229 VSUBS 0.009642f
C344 B.n230 VSUBS 0.009642f
C345 B.n231 VSUBS 0.009642f
C346 B.n232 VSUBS 0.009642f
C347 B.n233 VSUBS 0.009642f
C348 B.n234 VSUBS 0.009642f
C349 B.n235 VSUBS 0.009642f
C350 B.n236 VSUBS 0.009642f
C351 B.n237 VSUBS 0.009642f
C352 B.n238 VSUBS 0.019838f
C353 B.n239 VSUBS 0.019838f
C354 B.n240 VSUBS 0.021283f
C355 B.n241 VSUBS 0.009642f
C356 B.n242 VSUBS 0.009642f
C357 B.n243 VSUBS 0.009642f
C358 B.n244 VSUBS 0.009642f
C359 B.n245 VSUBS 0.009642f
C360 B.n246 VSUBS 0.009642f
C361 B.n247 VSUBS 0.009642f
C362 B.n248 VSUBS 0.009642f
C363 B.n249 VSUBS 0.009642f
C364 B.n250 VSUBS 0.009642f
C365 B.n251 VSUBS 0.009642f
C366 B.n252 VSUBS 0.009642f
C367 B.n253 VSUBS 0.009642f
C368 B.n254 VSUBS 0.009642f
C369 B.n255 VSUBS 0.009642f
C370 B.n256 VSUBS 0.009642f
C371 B.n257 VSUBS 0.006664f
C372 B.n258 VSUBS 0.02234f
C373 B.n259 VSUBS 0.007799f
C374 B.n260 VSUBS 0.009642f
C375 B.n261 VSUBS 0.009642f
C376 B.n262 VSUBS 0.009642f
C377 B.n263 VSUBS 0.009642f
C378 B.n264 VSUBS 0.009642f
C379 B.n265 VSUBS 0.009642f
C380 B.n266 VSUBS 0.009642f
C381 B.n267 VSUBS 0.009642f
C382 B.n268 VSUBS 0.009642f
C383 B.n269 VSUBS 0.009642f
C384 B.n270 VSUBS 0.009642f
C385 B.n271 VSUBS 0.007799f
C386 B.n272 VSUBS 0.02234f
C387 B.n273 VSUBS 0.006664f
C388 B.n274 VSUBS 0.009642f
C389 B.n275 VSUBS 0.009642f
C390 B.n276 VSUBS 0.009642f
C391 B.n277 VSUBS 0.009642f
C392 B.n278 VSUBS 0.009642f
C393 B.n279 VSUBS 0.009642f
C394 B.n280 VSUBS 0.009642f
C395 B.n281 VSUBS 0.009642f
C396 B.n282 VSUBS 0.009642f
C397 B.n283 VSUBS 0.009642f
C398 B.n284 VSUBS 0.009642f
C399 B.n285 VSUBS 0.009642f
C400 B.n286 VSUBS 0.009642f
C401 B.n287 VSUBS 0.009642f
C402 B.n288 VSUBS 0.009642f
C403 B.n289 VSUBS 0.009642f
C404 B.n290 VSUBS 0.021283f
C405 B.n291 VSUBS 0.019838f
C406 B.n292 VSUBS 0.019838f
C407 B.n293 VSUBS 0.009642f
C408 B.n294 VSUBS 0.009642f
C409 B.n295 VSUBS 0.009642f
C410 B.n296 VSUBS 0.009642f
C411 B.n297 VSUBS 0.009642f
C412 B.n298 VSUBS 0.009642f
C413 B.n299 VSUBS 0.009642f
C414 B.n300 VSUBS 0.009642f
C415 B.n301 VSUBS 0.009642f
C416 B.n302 VSUBS 0.009642f
C417 B.n303 VSUBS 0.009642f
C418 B.n304 VSUBS 0.009642f
C419 B.n305 VSUBS 0.009642f
C420 B.n306 VSUBS 0.009642f
C421 B.n307 VSUBS 0.009642f
C422 B.n308 VSUBS 0.009642f
C423 B.n309 VSUBS 0.009642f
C424 B.n310 VSUBS 0.009642f
C425 B.n311 VSUBS 0.009642f
C426 B.n312 VSUBS 0.009642f
C427 B.n313 VSUBS 0.009642f
C428 B.n314 VSUBS 0.009642f
C429 B.n315 VSUBS 0.009642f
C430 B.n316 VSUBS 0.009642f
C431 B.n317 VSUBS 0.009642f
C432 B.n318 VSUBS 0.009642f
C433 B.n319 VSUBS 0.009642f
C434 B.n320 VSUBS 0.009642f
C435 B.n321 VSUBS 0.009642f
C436 B.n322 VSUBS 0.009642f
C437 B.n323 VSUBS 0.012583f
C438 B.n324 VSUBS 0.013403f
C439 B.n325 VSUBS 0.026654f
.ends

