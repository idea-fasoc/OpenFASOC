* NGSPICE file created from diff_pair_sample_1060.ext - technology: sky130A

.subckt diff_pair_sample_1060 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=1.3533 pd=7.72 as=1.3533 ps=7.72 w=3.47 l=0.88
X1 VDD1.t1 VP.t0 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=1.3533 pd=7.72 as=1.3533 ps=7.72 w=3.47 l=0.88
X2 VDD1.t0 VP.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.3533 pd=7.72 as=1.3533 ps=7.72 w=3.47 l=0.88
X3 VDD2.t0 VN.t1 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=1.3533 pd=7.72 as=1.3533 ps=7.72 w=3.47 l=0.88
X4 B.t15 B.t13 B.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=1.3533 pd=7.72 as=0 ps=0 w=3.47 l=0.88
X5 B.t12 B.t10 B.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=1.3533 pd=7.72 as=0 ps=0 w=3.47 l=0.88
X6 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=1.3533 pd=7.72 as=0 ps=0 w=3.47 l=0.88
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=1.3533 pd=7.72 as=0 ps=0 w=3.47 l=0.88
R0 VN VN.t0 335.274
R1 VN VN.t1 301.296
R2 VTAIL.n1 VTAIL.t1 64.1939
R3 VTAIL.n3 VTAIL.t2 64.1938
R4 VTAIL.n0 VTAIL.t0 64.1938
R5 VTAIL.n2 VTAIL.t3 64.1938
R6 VTAIL.n1 VTAIL.n0 17.4617
R7 VTAIL.n3 VTAIL.n2 16.4186
R8 VTAIL.n2 VTAIL.n1 0.991879
R9 VTAIL VTAIL.n0 0.789293
R10 VTAIL VTAIL.n3 0.203086
R11 VDD2.n0 VDD2.t0 109.626
R12 VDD2.n0 VDD2.t1 80.8726
R13 VDD2 VDD2.n0 0.319466
R14 B.n346 B.n345 585
R15 B.n347 B.n346 585
R16 B.n139 B.n53 585
R17 B.n138 B.n137 585
R18 B.n136 B.n135 585
R19 B.n134 B.n133 585
R20 B.n132 B.n131 585
R21 B.n130 B.n129 585
R22 B.n128 B.n127 585
R23 B.n126 B.n125 585
R24 B.n124 B.n123 585
R25 B.n122 B.n121 585
R26 B.n120 B.n119 585
R27 B.n118 B.n117 585
R28 B.n116 B.n115 585
R29 B.n114 B.n113 585
R30 B.n112 B.n111 585
R31 B.n110 B.n109 585
R32 B.n108 B.n107 585
R33 B.n106 B.n105 585
R34 B.n104 B.n103 585
R35 B.n102 B.n101 585
R36 B.n100 B.n99 585
R37 B.n98 B.n97 585
R38 B.n96 B.n95 585
R39 B.n94 B.n93 585
R40 B.n92 B.n91 585
R41 B.n89 B.n88 585
R42 B.n87 B.n86 585
R43 B.n85 B.n84 585
R44 B.n83 B.n82 585
R45 B.n81 B.n80 585
R46 B.n79 B.n78 585
R47 B.n77 B.n76 585
R48 B.n75 B.n74 585
R49 B.n73 B.n72 585
R50 B.n71 B.n70 585
R51 B.n69 B.n68 585
R52 B.n67 B.n66 585
R53 B.n65 B.n64 585
R54 B.n63 B.n62 585
R55 B.n61 B.n60 585
R56 B.n32 B.n31 585
R57 B.n350 B.n349 585
R58 B.n344 B.n54 585
R59 B.n54 B.n29 585
R60 B.n343 B.n28 585
R61 B.n354 B.n28 585
R62 B.n342 B.n27 585
R63 B.n355 B.n27 585
R64 B.n341 B.n26 585
R65 B.n356 B.n26 585
R66 B.n340 B.n339 585
R67 B.n339 B.n25 585
R68 B.n338 B.n21 585
R69 B.n362 B.n21 585
R70 B.n337 B.n20 585
R71 B.n363 B.n20 585
R72 B.n336 B.n19 585
R73 B.n364 B.n19 585
R74 B.n335 B.n334 585
R75 B.n334 B.n15 585
R76 B.n333 B.n14 585
R77 B.n370 B.n14 585
R78 B.n332 B.n13 585
R79 B.n371 B.n13 585
R80 B.n331 B.n12 585
R81 B.n372 B.n12 585
R82 B.n330 B.n329 585
R83 B.n329 B.n8 585
R84 B.n328 B.n7 585
R85 B.n378 B.n7 585
R86 B.n327 B.n6 585
R87 B.n379 B.n6 585
R88 B.n326 B.n5 585
R89 B.n380 B.n5 585
R90 B.n325 B.n324 585
R91 B.n324 B.n4 585
R92 B.n323 B.n140 585
R93 B.n323 B.n322 585
R94 B.n313 B.n141 585
R95 B.n142 B.n141 585
R96 B.n315 B.n314 585
R97 B.n316 B.n315 585
R98 B.n312 B.n147 585
R99 B.n147 B.n146 585
R100 B.n311 B.n310 585
R101 B.n310 B.n309 585
R102 B.n149 B.n148 585
R103 B.n150 B.n149 585
R104 B.n302 B.n301 585
R105 B.n303 B.n302 585
R106 B.n300 B.n155 585
R107 B.n155 B.n154 585
R108 B.n299 B.n298 585
R109 B.n298 B.n297 585
R110 B.n157 B.n156 585
R111 B.n290 B.n157 585
R112 B.n289 B.n288 585
R113 B.n291 B.n289 585
R114 B.n287 B.n162 585
R115 B.n162 B.n161 585
R116 B.n286 B.n285 585
R117 B.n285 B.n284 585
R118 B.n164 B.n163 585
R119 B.n165 B.n164 585
R120 B.n280 B.n279 585
R121 B.n168 B.n167 585
R122 B.n276 B.n275 585
R123 B.n277 B.n276 585
R124 B.n274 B.n189 585
R125 B.n273 B.n272 585
R126 B.n271 B.n270 585
R127 B.n269 B.n268 585
R128 B.n267 B.n266 585
R129 B.n265 B.n264 585
R130 B.n263 B.n262 585
R131 B.n261 B.n260 585
R132 B.n259 B.n258 585
R133 B.n257 B.n256 585
R134 B.n255 B.n254 585
R135 B.n253 B.n252 585
R136 B.n251 B.n250 585
R137 B.n249 B.n248 585
R138 B.n247 B.n246 585
R139 B.n245 B.n244 585
R140 B.n243 B.n242 585
R141 B.n241 B.n240 585
R142 B.n239 B.n238 585
R143 B.n237 B.n236 585
R144 B.n235 B.n234 585
R145 B.n233 B.n232 585
R146 B.n231 B.n230 585
R147 B.n228 B.n227 585
R148 B.n226 B.n225 585
R149 B.n224 B.n223 585
R150 B.n222 B.n221 585
R151 B.n220 B.n219 585
R152 B.n218 B.n217 585
R153 B.n216 B.n215 585
R154 B.n214 B.n213 585
R155 B.n212 B.n211 585
R156 B.n210 B.n209 585
R157 B.n208 B.n207 585
R158 B.n206 B.n205 585
R159 B.n204 B.n203 585
R160 B.n202 B.n201 585
R161 B.n200 B.n199 585
R162 B.n198 B.n197 585
R163 B.n196 B.n195 585
R164 B.n281 B.n166 585
R165 B.n166 B.n165 585
R166 B.n283 B.n282 585
R167 B.n284 B.n283 585
R168 B.n160 B.n159 585
R169 B.n161 B.n160 585
R170 B.n293 B.n292 585
R171 B.n292 B.n291 585
R172 B.n294 B.n158 585
R173 B.n290 B.n158 585
R174 B.n296 B.n295 585
R175 B.n297 B.n296 585
R176 B.n153 B.n152 585
R177 B.n154 B.n153 585
R178 B.n305 B.n304 585
R179 B.n304 B.n303 585
R180 B.n306 B.n151 585
R181 B.n151 B.n150 585
R182 B.n308 B.n307 585
R183 B.n309 B.n308 585
R184 B.n145 B.n144 585
R185 B.n146 B.n145 585
R186 B.n318 B.n317 585
R187 B.n317 B.n316 585
R188 B.n319 B.n143 585
R189 B.n143 B.n142 585
R190 B.n321 B.n320 585
R191 B.n322 B.n321 585
R192 B.n2 B.n0 585
R193 B.n4 B.n2 585
R194 B.n3 B.n1 585
R195 B.n379 B.n3 585
R196 B.n377 B.n376 585
R197 B.n378 B.n377 585
R198 B.n375 B.n9 585
R199 B.n9 B.n8 585
R200 B.n374 B.n373 585
R201 B.n373 B.n372 585
R202 B.n11 B.n10 585
R203 B.n371 B.n11 585
R204 B.n369 B.n368 585
R205 B.n370 B.n369 585
R206 B.n367 B.n16 585
R207 B.n16 B.n15 585
R208 B.n366 B.n365 585
R209 B.n365 B.n364 585
R210 B.n18 B.n17 585
R211 B.n363 B.n18 585
R212 B.n361 B.n360 585
R213 B.n362 B.n361 585
R214 B.n359 B.n22 585
R215 B.n25 B.n22 585
R216 B.n358 B.n357 585
R217 B.n357 B.n356 585
R218 B.n24 B.n23 585
R219 B.n355 B.n24 585
R220 B.n353 B.n352 585
R221 B.n354 B.n353 585
R222 B.n351 B.n30 585
R223 B.n30 B.n29 585
R224 B.n382 B.n381 585
R225 B.n381 B.n380 585
R226 B.n279 B.n166 516.524
R227 B.n349 B.n30 516.524
R228 B.n195 B.n164 516.524
R229 B.n346 B.n54 516.524
R230 B.n193 B.t2 297.067
R231 B.n190 B.t10 297.067
R232 B.n58 B.t13 297.067
R233 B.n55 B.t6 297.067
R234 B.n347 B.n52 256.663
R235 B.n347 B.n51 256.663
R236 B.n347 B.n50 256.663
R237 B.n347 B.n49 256.663
R238 B.n347 B.n48 256.663
R239 B.n347 B.n47 256.663
R240 B.n347 B.n46 256.663
R241 B.n347 B.n45 256.663
R242 B.n347 B.n44 256.663
R243 B.n347 B.n43 256.663
R244 B.n347 B.n42 256.663
R245 B.n347 B.n41 256.663
R246 B.n347 B.n40 256.663
R247 B.n347 B.n39 256.663
R248 B.n347 B.n38 256.663
R249 B.n347 B.n37 256.663
R250 B.n347 B.n36 256.663
R251 B.n347 B.n35 256.663
R252 B.n347 B.n34 256.663
R253 B.n347 B.n33 256.663
R254 B.n348 B.n347 256.663
R255 B.n278 B.n277 256.663
R256 B.n277 B.n169 256.663
R257 B.n277 B.n170 256.663
R258 B.n277 B.n171 256.663
R259 B.n277 B.n172 256.663
R260 B.n277 B.n173 256.663
R261 B.n277 B.n174 256.663
R262 B.n277 B.n175 256.663
R263 B.n277 B.n176 256.663
R264 B.n277 B.n177 256.663
R265 B.n277 B.n178 256.663
R266 B.n277 B.n179 256.663
R267 B.n277 B.n180 256.663
R268 B.n277 B.n181 256.663
R269 B.n277 B.n182 256.663
R270 B.n277 B.n183 256.663
R271 B.n277 B.n184 256.663
R272 B.n277 B.n185 256.663
R273 B.n277 B.n186 256.663
R274 B.n277 B.n187 256.663
R275 B.n277 B.n188 256.663
R276 B.n277 B.n165 174.445
R277 B.n347 B.n29 174.445
R278 B.n283 B.n166 163.367
R279 B.n283 B.n160 163.367
R280 B.n292 B.n160 163.367
R281 B.n292 B.n158 163.367
R282 B.n296 B.n158 163.367
R283 B.n296 B.n153 163.367
R284 B.n304 B.n153 163.367
R285 B.n304 B.n151 163.367
R286 B.n308 B.n151 163.367
R287 B.n308 B.n145 163.367
R288 B.n317 B.n145 163.367
R289 B.n317 B.n143 163.367
R290 B.n321 B.n143 163.367
R291 B.n321 B.n2 163.367
R292 B.n381 B.n2 163.367
R293 B.n381 B.n3 163.367
R294 B.n377 B.n3 163.367
R295 B.n377 B.n9 163.367
R296 B.n373 B.n9 163.367
R297 B.n373 B.n11 163.367
R298 B.n369 B.n11 163.367
R299 B.n369 B.n16 163.367
R300 B.n365 B.n16 163.367
R301 B.n365 B.n18 163.367
R302 B.n361 B.n18 163.367
R303 B.n361 B.n22 163.367
R304 B.n357 B.n22 163.367
R305 B.n357 B.n24 163.367
R306 B.n353 B.n24 163.367
R307 B.n353 B.n30 163.367
R308 B.n276 B.n168 163.367
R309 B.n276 B.n189 163.367
R310 B.n272 B.n271 163.367
R311 B.n268 B.n267 163.367
R312 B.n264 B.n263 163.367
R313 B.n260 B.n259 163.367
R314 B.n256 B.n255 163.367
R315 B.n252 B.n251 163.367
R316 B.n248 B.n247 163.367
R317 B.n244 B.n243 163.367
R318 B.n240 B.n239 163.367
R319 B.n236 B.n235 163.367
R320 B.n232 B.n231 163.367
R321 B.n227 B.n226 163.367
R322 B.n223 B.n222 163.367
R323 B.n219 B.n218 163.367
R324 B.n215 B.n214 163.367
R325 B.n211 B.n210 163.367
R326 B.n207 B.n206 163.367
R327 B.n203 B.n202 163.367
R328 B.n199 B.n198 163.367
R329 B.n285 B.n164 163.367
R330 B.n285 B.n162 163.367
R331 B.n289 B.n162 163.367
R332 B.n289 B.n157 163.367
R333 B.n298 B.n157 163.367
R334 B.n298 B.n155 163.367
R335 B.n302 B.n155 163.367
R336 B.n302 B.n149 163.367
R337 B.n310 B.n149 163.367
R338 B.n310 B.n147 163.367
R339 B.n315 B.n147 163.367
R340 B.n315 B.n141 163.367
R341 B.n323 B.n141 163.367
R342 B.n324 B.n323 163.367
R343 B.n324 B.n5 163.367
R344 B.n6 B.n5 163.367
R345 B.n7 B.n6 163.367
R346 B.n329 B.n7 163.367
R347 B.n329 B.n12 163.367
R348 B.n13 B.n12 163.367
R349 B.n14 B.n13 163.367
R350 B.n334 B.n14 163.367
R351 B.n334 B.n19 163.367
R352 B.n20 B.n19 163.367
R353 B.n21 B.n20 163.367
R354 B.n339 B.n21 163.367
R355 B.n339 B.n26 163.367
R356 B.n27 B.n26 163.367
R357 B.n28 B.n27 163.367
R358 B.n54 B.n28 163.367
R359 B.n60 B.n32 163.367
R360 B.n64 B.n63 163.367
R361 B.n68 B.n67 163.367
R362 B.n72 B.n71 163.367
R363 B.n76 B.n75 163.367
R364 B.n80 B.n79 163.367
R365 B.n84 B.n83 163.367
R366 B.n88 B.n87 163.367
R367 B.n93 B.n92 163.367
R368 B.n97 B.n96 163.367
R369 B.n101 B.n100 163.367
R370 B.n105 B.n104 163.367
R371 B.n109 B.n108 163.367
R372 B.n113 B.n112 163.367
R373 B.n117 B.n116 163.367
R374 B.n121 B.n120 163.367
R375 B.n125 B.n124 163.367
R376 B.n129 B.n128 163.367
R377 B.n133 B.n132 163.367
R378 B.n137 B.n136 163.367
R379 B.n346 B.n53 163.367
R380 B.n193 B.t5 97.4918
R381 B.n55 B.t8 97.4918
R382 B.n190 B.t12 97.489
R383 B.n58 B.t14 97.489
R384 B.n284 B.n165 85.3399
R385 B.n284 B.n161 85.3399
R386 B.n291 B.n161 85.3399
R387 B.n291 B.n290 85.3399
R388 B.n297 B.n154 85.3399
R389 B.n303 B.n154 85.3399
R390 B.n303 B.n150 85.3399
R391 B.n309 B.n150 85.3399
R392 B.n309 B.n146 85.3399
R393 B.n316 B.n146 85.3399
R394 B.n322 B.n142 85.3399
R395 B.n322 B.n4 85.3399
R396 B.n380 B.n4 85.3399
R397 B.n380 B.n379 85.3399
R398 B.n379 B.n378 85.3399
R399 B.n378 B.n8 85.3399
R400 B.n372 B.n371 85.3399
R401 B.n371 B.n370 85.3399
R402 B.n370 B.n15 85.3399
R403 B.n364 B.n15 85.3399
R404 B.n364 B.n363 85.3399
R405 B.n363 B.n362 85.3399
R406 B.n356 B.n25 85.3399
R407 B.n356 B.n355 85.3399
R408 B.n355 B.n354 85.3399
R409 B.n354 B.n29 85.3399
R410 B.n194 B.t4 74.0252
R411 B.n56 B.t9 74.0252
R412 B.n191 B.t11 74.0223
R413 B.n59 B.t15 74.0223
R414 B.n290 B.t3 72.79
R415 B.n25 B.t7 72.79
R416 B.n279 B.n278 71.676
R417 B.n189 B.n169 71.676
R418 B.n271 B.n170 71.676
R419 B.n267 B.n171 71.676
R420 B.n263 B.n172 71.676
R421 B.n259 B.n173 71.676
R422 B.n255 B.n174 71.676
R423 B.n251 B.n175 71.676
R424 B.n247 B.n176 71.676
R425 B.n243 B.n177 71.676
R426 B.n239 B.n178 71.676
R427 B.n235 B.n179 71.676
R428 B.n231 B.n180 71.676
R429 B.n226 B.n181 71.676
R430 B.n222 B.n182 71.676
R431 B.n218 B.n183 71.676
R432 B.n214 B.n184 71.676
R433 B.n210 B.n185 71.676
R434 B.n206 B.n186 71.676
R435 B.n202 B.n187 71.676
R436 B.n198 B.n188 71.676
R437 B.n349 B.n348 71.676
R438 B.n60 B.n33 71.676
R439 B.n64 B.n34 71.676
R440 B.n68 B.n35 71.676
R441 B.n72 B.n36 71.676
R442 B.n76 B.n37 71.676
R443 B.n80 B.n38 71.676
R444 B.n84 B.n39 71.676
R445 B.n88 B.n40 71.676
R446 B.n93 B.n41 71.676
R447 B.n97 B.n42 71.676
R448 B.n101 B.n43 71.676
R449 B.n105 B.n44 71.676
R450 B.n109 B.n45 71.676
R451 B.n113 B.n46 71.676
R452 B.n117 B.n47 71.676
R453 B.n121 B.n48 71.676
R454 B.n125 B.n49 71.676
R455 B.n129 B.n50 71.676
R456 B.n133 B.n51 71.676
R457 B.n137 B.n52 71.676
R458 B.n53 B.n52 71.676
R459 B.n136 B.n51 71.676
R460 B.n132 B.n50 71.676
R461 B.n128 B.n49 71.676
R462 B.n124 B.n48 71.676
R463 B.n120 B.n47 71.676
R464 B.n116 B.n46 71.676
R465 B.n112 B.n45 71.676
R466 B.n108 B.n44 71.676
R467 B.n104 B.n43 71.676
R468 B.n100 B.n42 71.676
R469 B.n96 B.n41 71.676
R470 B.n92 B.n40 71.676
R471 B.n87 B.n39 71.676
R472 B.n83 B.n38 71.676
R473 B.n79 B.n37 71.676
R474 B.n75 B.n36 71.676
R475 B.n71 B.n35 71.676
R476 B.n67 B.n34 71.676
R477 B.n63 B.n33 71.676
R478 B.n348 B.n32 71.676
R479 B.n278 B.n168 71.676
R480 B.n272 B.n169 71.676
R481 B.n268 B.n170 71.676
R482 B.n264 B.n171 71.676
R483 B.n260 B.n172 71.676
R484 B.n256 B.n173 71.676
R485 B.n252 B.n174 71.676
R486 B.n248 B.n175 71.676
R487 B.n244 B.n176 71.676
R488 B.n240 B.n177 71.676
R489 B.n236 B.n178 71.676
R490 B.n232 B.n179 71.676
R491 B.n227 B.n180 71.676
R492 B.n223 B.n181 71.676
R493 B.n219 B.n182 71.676
R494 B.n215 B.n183 71.676
R495 B.n211 B.n184 71.676
R496 B.n207 B.n185 71.676
R497 B.n203 B.n186 71.676
R498 B.n199 B.n187 71.676
R499 B.n195 B.n188 71.676
R500 B.n229 B.n194 59.5399
R501 B.n192 B.n191 59.5399
R502 B.n90 B.n59 59.5399
R503 B.n57 B.n56 59.5399
R504 B.n316 B.t0 52.7101
R505 B.n372 B.t1 52.7101
R506 B.n351 B.n350 33.5615
R507 B.n345 B.n344 33.5615
R508 B.n196 B.n163 33.5615
R509 B.n281 B.n280 33.5615
R510 B.t0 B.n142 32.6303
R511 B.t1 B.n8 32.6303
R512 B.n194 B.n193 23.4672
R513 B.n191 B.n190 23.4672
R514 B.n59 B.n58 23.4672
R515 B.n56 B.n55 23.4672
R516 B B.n382 18.0485
R517 B.n297 B.t3 12.5504
R518 B.n362 B.t7 12.5504
R519 B.n350 B.n31 10.6151
R520 B.n61 B.n31 10.6151
R521 B.n62 B.n61 10.6151
R522 B.n65 B.n62 10.6151
R523 B.n66 B.n65 10.6151
R524 B.n69 B.n66 10.6151
R525 B.n70 B.n69 10.6151
R526 B.n73 B.n70 10.6151
R527 B.n74 B.n73 10.6151
R528 B.n77 B.n74 10.6151
R529 B.n78 B.n77 10.6151
R530 B.n81 B.n78 10.6151
R531 B.n82 B.n81 10.6151
R532 B.n85 B.n82 10.6151
R533 B.n86 B.n85 10.6151
R534 B.n89 B.n86 10.6151
R535 B.n94 B.n91 10.6151
R536 B.n95 B.n94 10.6151
R537 B.n98 B.n95 10.6151
R538 B.n99 B.n98 10.6151
R539 B.n102 B.n99 10.6151
R540 B.n103 B.n102 10.6151
R541 B.n106 B.n103 10.6151
R542 B.n107 B.n106 10.6151
R543 B.n111 B.n110 10.6151
R544 B.n114 B.n111 10.6151
R545 B.n115 B.n114 10.6151
R546 B.n118 B.n115 10.6151
R547 B.n119 B.n118 10.6151
R548 B.n122 B.n119 10.6151
R549 B.n123 B.n122 10.6151
R550 B.n126 B.n123 10.6151
R551 B.n127 B.n126 10.6151
R552 B.n130 B.n127 10.6151
R553 B.n131 B.n130 10.6151
R554 B.n134 B.n131 10.6151
R555 B.n135 B.n134 10.6151
R556 B.n138 B.n135 10.6151
R557 B.n139 B.n138 10.6151
R558 B.n345 B.n139 10.6151
R559 B.n286 B.n163 10.6151
R560 B.n287 B.n286 10.6151
R561 B.n288 B.n287 10.6151
R562 B.n288 B.n156 10.6151
R563 B.n299 B.n156 10.6151
R564 B.n300 B.n299 10.6151
R565 B.n301 B.n300 10.6151
R566 B.n301 B.n148 10.6151
R567 B.n311 B.n148 10.6151
R568 B.n312 B.n311 10.6151
R569 B.n314 B.n312 10.6151
R570 B.n314 B.n313 10.6151
R571 B.n313 B.n140 10.6151
R572 B.n325 B.n140 10.6151
R573 B.n326 B.n325 10.6151
R574 B.n327 B.n326 10.6151
R575 B.n328 B.n327 10.6151
R576 B.n330 B.n328 10.6151
R577 B.n331 B.n330 10.6151
R578 B.n332 B.n331 10.6151
R579 B.n333 B.n332 10.6151
R580 B.n335 B.n333 10.6151
R581 B.n336 B.n335 10.6151
R582 B.n337 B.n336 10.6151
R583 B.n338 B.n337 10.6151
R584 B.n340 B.n338 10.6151
R585 B.n341 B.n340 10.6151
R586 B.n342 B.n341 10.6151
R587 B.n343 B.n342 10.6151
R588 B.n344 B.n343 10.6151
R589 B.n280 B.n167 10.6151
R590 B.n275 B.n167 10.6151
R591 B.n275 B.n274 10.6151
R592 B.n274 B.n273 10.6151
R593 B.n273 B.n270 10.6151
R594 B.n270 B.n269 10.6151
R595 B.n269 B.n266 10.6151
R596 B.n266 B.n265 10.6151
R597 B.n265 B.n262 10.6151
R598 B.n262 B.n261 10.6151
R599 B.n261 B.n258 10.6151
R600 B.n258 B.n257 10.6151
R601 B.n257 B.n254 10.6151
R602 B.n254 B.n253 10.6151
R603 B.n253 B.n250 10.6151
R604 B.n250 B.n249 10.6151
R605 B.n246 B.n245 10.6151
R606 B.n245 B.n242 10.6151
R607 B.n242 B.n241 10.6151
R608 B.n241 B.n238 10.6151
R609 B.n238 B.n237 10.6151
R610 B.n237 B.n234 10.6151
R611 B.n234 B.n233 10.6151
R612 B.n233 B.n230 10.6151
R613 B.n228 B.n225 10.6151
R614 B.n225 B.n224 10.6151
R615 B.n224 B.n221 10.6151
R616 B.n221 B.n220 10.6151
R617 B.n220 B.n217 10.6151
R618 B.n217 B.n216 10.6151
R619 B.n216 B.n213 10.6151
R620 B.n213 B.n212 10.6151
R621 B.n212 B.n209 10.6151
R622 B.n209 B.n208 10.6151
R623 B.n208 B.n205 10.6151
R624 B.n205 B.n204 10.6151
R625 B.n204 B.n201 10.6151
R626 B.n201 B.n200 10.6151
R627 B.n200 B.n197 10.6151
R628 B.n197 B.n196 10.6151
R629 B.n282 B.n281 10.6151
R630 B.n282 B.n159 10.6151
R631 B.n293 B.n159 10.6151
R632 B.n294 B.n293 10.6151
R633 B.n295 B.n294 10.6151
R634 B.n295 B.n152 10.6151
R635 B.n305 B.n152 10.6151
R636 B.n306 B.n305 10.6151
R637 B.n307 B.n306 10.6151
R638 B.n307 B.n144 10.6151
R639 B.n318 B.n144 10.6151
R640 B.n319 B.n318 10.6151
R641 B.n320 B.n319 10.6151
R642 B.n320 B.n0 10.6151
R643 B.n376 B.n1 10.6151
R644 B.n376 B.n375 10.6151
R645 B.n375 B.n374 10.6151
R646 B.n374 B.n10 10.6151
R647 B.n368 B.n10 10.6151
R648 B.n368 B.n367 10.6151
R649 B.n367 B.n366 10.6151
R650 B.n366 B.n17 10.6151
R651 B.n360 B.n17 10.6151
R652 B.n360 B.n359 10.6151
R653 B.n359 B.n358 10.6151
R654 B.n358 B.n23 10.6151
R655 B.n352 B.n23 10.6151
R656 B.n352 B.n351 10.6151
R657 B.n91 B.n90 7.18099
R658 B.n107 B.n57 7.18099
R659 B.n246 B.n192 7.18099
R660 B.n230 B.n229 7.18099
R661 B.n90 B.n89 3.43465
R662 B.n110 B.n57 3.43465
R663 B.n249 B.n192 3.43465
R664 B.n229 B.n228 3.43465
R665 B.n382 B.n0 2.81026
R666 B.n382 B.n1 2.81026
R667 VP.n0 VP.t0 334.892
R668 VP.n0 VP.t1 301.245
R669 VP VP.n0 0.0516364
R670 VDD1 VDD1.t0 110.412
R671 VDD1 VDD1.t1 81.1916
C0 VDD1 VTAIL 2.48294f
C1 VTAIL VP 0.768029f
C2 VTAIL VN 0.753793f
C3 VDD2 VDD1 0.477691f
C4 VDD2 VP 0.266293f
C5 VDD2 VN 0.791868f
C6 VDD2 VTAIL 2.52296f
C7 VDD1 VP 0.90314f
C8 VDD1 VN 0.153303f
C9 VP VN 3.06938f
C10 VDD2 B 2.259765f
C11 VDD1 B 3.83226f
C12 VTAIL B 3.050335f
C13 VN B 5.80172f
C14 VP B 3.558993f
C15 VDD1.t1 B 0.418399f
C16 VDD1.t0 B 0.60256f
C17 VP.t0 B 0.538229f
C18 VP.t1 B 0.427435f
C19 VP.n0 B 2.11746f
C20 VDD2.t0 B 0.602607f
C21 VDD2.t1 B 0.427621f
C22 VDD2.n0 B 1.42593f
C23 VTAIL.t0 B 0.458073f
C24 VTAIL.n0 B 0.811314f
C25 VTAIL.t1 B 0.458076f
C26 VTAIL.n1 B 0.823624f
C27 VTAIL.t3 B 0.458073f
C28 VTAIL.n2 B 0.760228f
C29 VTAIL.t2 B 0.458073f
C30 VTAIL.n3 B 0.712286f
C31 VN.t1 B 0.420452f
C32 VN.t0 B 0.532963f
.ends

