* NGSPICE file created from diff_pair_sample_0121.ext - technology: sky130A

.subckt diff_pair_sample_0121 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=0.42735 pd=2.92 as=1.0101 ps=5.96 w=2.59 l=0.3
X1 VDD2.t5 VN.t0 VTAIL.t11 B.t4 sky130_fd_pr__nfet_01v8 ad=1.0101 pd=5.96 as=0.42735 ps=2.92 w=2.59 l=0.3
X2 B.t19 B.t17 B.t18 B.t14 sky130_fd_pr__nfet_01v8 ad=1.0101 pd=5.96 as=0 ps=0 w=2.59 l=0.3
X3 VDD2.t4 VN.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.0101 pd=5.96 as=0.42735 ps=2.92 w=2.59 l=0.3
X4 VDD1.t4 VP.t1 VTAIL.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=1.0101 pd=5.96 as=0.42735 ps=2.92 w=2.59 l=0.3
X5 B.t16 B.t13 B.t15 B.t14 sky130_fd_pr__nfet_01v8 ad=1.0101 pd=5.96 as=0 ps=0 w=2.59 l=0.3
X6 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=1.0101 pd=5.96 as=0 ps=0 w=2.59 l=0.3
X7 VTAIL.t5 VP.t2 VDD1.t3 B.t5 sky130_fd_pr__nfet_01v8 ad=0.42735 pd=2.92 as=0.42735 ps=2.92 w=2.59 l=0.3
X8 VDD1.t2 VP.t3 VTAIL.t3 B.t4 sky130_fd_pr__nfet_01v8 ad=1.0101 pd=5.96 as=0.42735 ps=2.92 w=2.59 l=0.3
X9 VDD2.t3 VN.t2 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.42735 pd=2.92 as=1.0101 ps=5.96 w=2.59 l=0.3
X10 VDD2.t2 VN.t3 VTAIL.t10 B.t3 sky130_fd_pr__nfet_01v8 ad=0.42735 pd=2.92 as=1.0101 ps=5.96 w=2.59 l=0.3
X11 VTAIL.t7 VP.t4 VDD1.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=0.42735 pd=2.92 as=0.42735 ps=2.92 w=2.59 l=0.3
X12 VDD1.t0 VP.t5 VTAIL.t8 B.t3 sky130_fd_pr__nfet_01v8 ad=0.42735 pd=2.92 as=1.0101 ps=5.96 w=2.59 l=0.3
X13 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=1.0101 pd=5.96 as=0 ps=0 w=2.59 l=0.3
X14 VTAIL.t9 VN.t4 VDD2.t1 B.t5 sky130_fd_pr__nfet_01v8 ad=0.42735 pd=2.92 as=0.42735 ps=2.92 w=2.59 l=0.3
X15 VTAIL.t2 VN.t5 VDD2.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=0.42735 pd=2.92 as=0.42735 ps=2.92 w=2.59 l=0.3
R0 VP.n7 VP.t0 368.803
R1 VP.n5 VP.t3 368.803
R2 VP.n0 VP.t1 368.803
R3 VP.n2 VP.t5 368.803
R4 VP.n6 VP.t4 313.3
R5 VP.n1 VP.t2 313.3
R6 VP.n3 VP.n0 161.489
R7 VP.n8 VP.n7 161.3
R8 VP.n3 VP.n2 161.3
R9 VP.n5 VP.n4 161.3
R10 VP.n6 VP.n5 36.5157
R11 VP.n7 VP.n6 36.5157
R12 VP.n1 VP.n0 36.5157
R13 VP.n2 VP.n1 36.5157
R14 VP.n4 VP.n3 32.671
R15 VP.n8 VP.n4 0.189894
R16 VP VP.n8 0.0516364
R17 VTAIL.n50 VTAIL.n44 289.615
R18 VTAIL.n8 VTAIL.n2 289.615
R19 VTAIL.n38 VTAIL.n32 289.615
R20 VTAIL.n24 VTAIL.n18 289.615
R21 VTAIL.n49 VTAIL.n48 185
R22 VTAIL.n51 VTAIL.n50 185
R23 VTAIL.n7 VTAIL.n6 185
R24 VTAIL.n9 VTAIL.n8 185
R25 VTAIL.n39 VTAIL.n38 185
R26 VTAIL.n37 VTAIL.n36 185
R27 VTAIL.n25 VTAIL.n24 185
R28 VTAIL.n23 VTAIL.n22 185
R29 VTAIL.n47 VTAIL.t10 151.613
R30 VTAIL.n5 VTAIL.t6 151.613
R31 VTAIL.n35 VTAIL.t8 151.613
R32 VTAIL.n21 VTAIL.t1 151.613
R33 VTAIL.n50 VTAIL.n49 104.615
R34 VTAIL.n8 VTAIL.n7 104.615
R35 VTAIL.n38 VTAIL.n37 104.615
R36 VTAIL.n24 VTAIL.n23 104.615
R37 VTAIL.n31 VTAIL.n30 71.9653
R38 VTAIL.n17 VTAIL.n16 71.9653
R39 VTAIL.n1 VTAIL.n0 71.9652
R40 VTAIL.n15 VTAIL.n14 71.9652
R41 VTAIL.n49 VTAIL.t10 52.3082
R42 VTAIL.n7 VTAIL.t6 52.3082
R43 VTAIL.n37 VTAIL.t8 52.3082
R44 VTAIL.n23 VTAIL.t1 52.3082
R45 VTAIL.n55 VTAIL.n54 35.8702
R46 VTAIL.n13 VTAIL.n12 35.8702
R47 VTAIL.n43 VTAIL.n42 35.8702
R48 VTAIL.n29 VTAIL.n28 35.8702
R49 VTAIL.n17 VTAIL.n15 15.6858
R50 VTAIL.n48 VTAIL.n47 15.3979
R51 VTAIL.n6 VTAIL.n5 15.3979
R52 VTAIL.n36 VTAIL.n35 15.3979
R53 VTAIL.n22 VTAIL.n21 15.3979
R54 VTAIL.n55 VTAIL.n43 15.1427
R55 VTAIL.n51 VTAIL.n46 12.8005
R56 VTAIL.n9 VTAIL.n4 12.8005
R57 VTAIL.n39 VTAIL.n34 12.8005
R58 VTAIL.n25 VTAIL.n20 12.8005
R59 VTAIL.n52 VTAIL.n44 12.0247
R60 VTAIL.n10 VTAIL.n2 12.0247
R61 VTAIL.n40 VTAIL.n32 12.0247
R62 VTAIL.n26 VTAIL.n18 12.0247
R63 VTAIL.n54 VTAIL.n53 9.45567
R64 VTAIL.n12 VTAIL.n11 9.45567
R65 VTAIL.n42 VTAIL.n41 9.45567
R66 VTAIL.n28 VTAIL.n27 9.45567
R67 VTAIL.n53 VTAIL.n52 9.3005
R68 VTAIL.n46 VTAIL.n45 9.3005
R69 VTAIL.n11 VTAIL.n10 9.3005
R70 VTAIL.n4 VTAIL.n3 9.3005
R71 VTAIL.n41 VTAIL.n40 9.3005
R72 VTAIL.n34 VTAIL.n33 9.3005
R73 VTAIL.n27 VTAIL.n26 9.3005
R74 VTAIL.n20 VTAIL.n19 9.3005
R75 VTAIL.n0 VTAIL.t0 7.64529
R76 VTAIL.n0 VTAIL.t9 7.64529
R77 VTAIL.n14 VTAIL.t3 7.64529
R78 VTAIL.n14 VTAIL.t7 7.64529
R79 VTAIL.n30 VTAIL.t4 7.64529
R80 VTAIL.n30 VTAIL.t5 7.64529
R81 VTAIL.n16 VTAIL.t11 7.64529
R82 VTAIL.n16 VTAIL.t2 7.64529
R83 VTAIL.n47 VTAIL.n45 4.69785
R84 VTAIL.n5 VTAIL.n3 4.69785
R85 VTAIL.n35 VTAIL.n33 4.69785
R86 VTAIL.n21 VTAIL.n19 4.69785
R87 VTAIL.n54 VTAIL.n44 1.93989
R88 VTAIL.n12 VTAIL.n2 1.93989
R89 VTAIL.n42 VTAIL.n32 1.93989
R90 VTAIL.n28 VTAIL.n18 1.93989
R91 VTAIL.n52 VTAIL.n51 1.16414
R92 VTAIL.n10 VTAIL.n9 1.16414
R93 VTAIL.n40 VTAIL.n39 1.16414
R94 VTAIL.n26 VTAIL.n25 1.16414
R95 VTAIL.n31 VTAIL.n29 0.741879
R96 VTAIL.n13 VTAIL.n1 0.741879
R97 VTAIL.n29 VTAIL.n17 0.543603
R98 VTAIL.n43 VTAIL.n31 0.543603
R99 VTAIL.n15 VTAIL.n13 0.543603
R100 VTAIL.n48 VTAIL.n46 0.388379
R101 VTAIL.n6 VTAIL.n4 0.388379
R102 VTAIL.n36 VTAIL.n34 0.388379
R103 VTAIL.n22 VTAIL.n20 0.388379
R104 VTAIL VTAIL.n55 0.349638
R105 VTAIL VTAIL.n1 0.194466
R106 VTAIL.n53 VTAIL.n45 0.155672
R107 VTAIL.n11 VTAIL.n3 0.155672
R108 VTAIL.n41 VTAIL.n33 0.155672
R109 VTAIL.n27 VTAIL.n19 0.155672
R110 VDD1.n6 VDD1.n0 289.615
R111 VDD1.n17 VDD1.n11 289.615
R112 VDD1.n7 VDD1.n6 185
R113 VDD1.n5 VDD1.n4 185
R114 VDD1.n16 VDD1.n15 185
R115 VDD1.n18 VDD1.n17 185
R116 VDD1.n3 VDD1.t4 151.613
R117 VDD1.n14 VDD1.t2 151.613
R118 VDD1.n6 VDD1.n5 104.615
R119 VDD1.n17 VDD1.n16 104.615
R120 VDD1.n23 VDD1.n22 88.7245
R121 VDD1.n25 VDD1.n24 88.644
R122 VDD1 VDD1.n10 53.0145
R123 VDD1.n23 VDD1.n21 52.901
R124 VDD1.n5 VDD1.t4 52.3082
R125 VDD1.n16 VDD1.t2 52.3082
R126 VDD1.n25 VDD1.n23 28.5677
R127 VDD1.n4 VDD1.n3 15.3979
R128 VDD1.n15 VDD1.n14 15.3979
R129 VDD1.n7 VDD1.n2 12.8005
R130 VDD1.n18 VDD1.n13 12.8005
R131 VDD1.n8 VDD1.n0 12.0247
R132 VDD1.n19 VDD1.n11 12.0247
R133 VDD1.n10 VDD1.n9 9.45567
R134 VDD1.n21 VDD1.n20 9.45567
R135 VDD1.n9 VDD1.n8 9.3005
R136 VDD1.n2 VDD1.n1 9.3005
R137 VDD1.n20 VDD1.n19 9.3005
R138 VDD1.n13 VDD1.n12 9.3005
R139 VDD1.n24 VDD1.t3 7.64529
R140 VDD1.n24 VDD1.t0 7.64529
R141 VDD1.n22 VDD1.t1 7.64529
R142 VDD1.n22 VDD1.t5 7.64529
R143 VDD1.n3 VDD1.n1 4.69785
R144 VDD1.n14 VDD1.n12 4.69785
R145 VDD1.n10 VDD1.n0 1.93989
R146 VDD1.n21 VDD1.n11 1.93989
R147 VDD1.n8 VDD1.n7 1.16414
R148 VDD1.n19 VDD1.n18 1.16414
R149 VDD1.n4 VDD1.n2 0.388379
R150 VDD1.n15 VDD1.n13 0.388379
R151 VDD1.n9 VDD1.n1 0.155672
R152 VDD1.n20 VDD1.n12 0.155672
R153 VDD1 VDD1.n25 0.0780862
R154 B.n319 B.n318 585
R155 B.n320 B.n319 585
R156 B.n124 B.n50 585
R157 B.n123 B.n122 585
R158 B.n121 B.n120 585
R159 B.n119 B.n118 585
R160 B.n117 B.n116 585
R161 B.n115 B.n114 585
R162 B.n113 B.n112 585
R163 B.n111 B.n110 585
R164 B.n109 B.n108 585
R165 B.n107 B.n106 585
R166 B.n105 B.n104 585
R167 B.n103 B.n102 585
R168 B.n101 B.n100 585
R169 B.n98 B.n97 585
R170 B.n96 B.n95 585
R171 B.n94 B.n93 585
R172 B.n92 B.n91 585
R173 B.n90 B.n89 585
R174 B.n88 B.n87 585
R175 B.n86 B.n85 585
R176 B.n84 B.n83 585
R177 B.n82 B.n81 585
R178 B.n80 B.n79 585
R179 B.n78 B.n77 585
R180 B.n76 B.n75 585
R181 B.n74 B.n73 585
R182 B.n72 B.n71 585
R183 B.n70 B.n69 585
R184 B.n68 B.n67 585
R185 B.n66 B.n65 585
R186 B.n64 B.n63 585
R187 B.n62 B.n61 585
R188 B.n60 B.n59 585
R189 B.n58 B.n57 585
R190 B.n32 B.n31 585
R191 B.n323 B.n322 585
R192 B.n317 B.n51 585
R193 B.n51 B.n29 585
R194 B.n316 B.n28 585
R195 B.n327 B.n28 585
R196 B.n315 B.n27 585
R197 B.n328 B.n27 585
R198 B.n314 B.n26 585
R199 B.n329 B.n26 585
R200 B.n313 B.n312 585
R201 B.n312 B.n25 585
R202 B.n311 B.n21 585
R203 B.n335 B.n21 585
R204 B.n310 B.n20 585
R205 B.n336 B.n20 585
R206 B.n309 B.n19 585
R207 B.n337 B.n19 585
R208 B.n308 B.n307 585
R209 B.n307 B.n15 585
R210 B.n306 B.n14 585
R211 B.n343 B.n14 585
R212 B.n305 B.n13 585
R213 B.n344 B.n13 585
R214 B.n304 B.n12 585
R215 B.n345 B.n12 585
R216 B.n303 B.n302 585
R217 B.n302 B.n301 585
R218 B.n300 B.n299 585
R219 B.n300 B.n8 585
R220 B.n298 B.n7 585
R221 B.n352 B.n7 585
R222 B.n297 B.n6 585
R223 B.n353 B.n6 585
R224 B.n296 B.n5 585
R225 B.n354 B.n5 585
R226 B.n295 B.n294 585
R227 B.n294 B.n4 585
R228 B.n293 B.n125 585
R229 B.n293 B.n292 585
R230 B.n282 B.n126 585
R231 B.n285 B.n126 585
R232 B.n284 B.n283 585
R233 B.n286 B.n284 585
R234 B.n281 B.n131 585
R235 B.n131 B.n130 585
R236 B.n280 B.n279 585
R237 B.n279 B.n278 585
R238 B.n133 B.n132 585
R239 B.n134 B.n133 585
R240 B.n271 B.n270 585
R241 B.n272 B.n271 585
R242 B.n269 B.n139 585
R243 B.n139 B.n138 585
R244 B.n268 B.n267 585
R245 B.n267 B.n266 585
R246 B.n141 B.n140 585
R247 B.n259 B.n141 585
R248 B.n258 B.n257 585
R249 B.n260 B.n258 585
R250 B.n256 B.n146 585
R251 B.n146 B.n145 585
R252 B.n255 B.n254 585
R253 B.n254 B.n253 585
R254 B.n148 B.n147 585
R255 B.n149 B.n148 585
R256 B.n249 B.n248 585
R257 B.n152 B.n151 585
R258 B.n245 B.n244 585
R259 B.n246 B.n245 585
R260 B.n243 B.n170 585
R261 B.n242 B.n241 585
R262 B.n240 B.n239 585
R263 B.n238 B.n237 585
R264 B.n236 B.n235 585
R265 B.n234 B.n233 585
R266 B.n232 B.n231 585
R267 B.n230 B.n229 585
R268 B.n228 B.n227 585
R269 B.n226 B.n225 585
R270 B.n224 B.n223 585
R271 B.n221 B.n220 585
R272 B.n219 B.n218 585
R273 B.n217 B.n216 585
R274 B.n215 B.n214 585
R275 B.n213 B.n212 585
R276 B.n211 B.n210 585
R277 B.n209 B.n208 585
R278 B.n207 B.n206 585
R279 B.n205 B.n204 585
R280 B.n203 B.n202 585
R281 B.n201 B.n200 585
R282 B.n199 B.n198 585
R283 B.n197 B.n196 585
R284 B.n195 B.n194 585
R285 B.n193 B.n192 585
R286 B.n191 B.n190 585
R287 B.n189 B.n188 585
R288 B.n187 B.n186 585
R289 B.n185 B.n184 585
R290 B.n183 B.n182 585
R291 B.n181 B.n180 585
R292 B.n179 B.n178 585
R293 B.n177 B.n176 585
R294 B.n250 B.n150 585
R295 B.n150 B.n149 585
R296 B.n252 B.n251 585
R297 B.n253 B.n252 585
R298 B.n144 B.n143 585
R299 B.n145 B.n144 585
R300 B.n262 B.n261 585
R301 B.n261 B.n260 585
R302 B.n263 B.n142 585
R303 B.n259 B.n142 585
R304 B.n265 B.n264 585
R305 B.n266 B.n265 585
R306 B.n137 B.n136 585
R307 B.n138 B.n137 585
R308 B.n274 B.n273 585
R309 B.n273 B.n272 585
R310 B.n275 B.n135 585
R311 B.n135 B.n134 585
R312 B.n277 B.n276 585
R313 B.n278 B.n277 585
R314 B.n129 B.n128 585
R315 B.n130 B.n129 585
R316 B.n288 B.n287 585
R317 B.n287 B.n286 585
R318 B.n289 B.n127 585
R319 B.n285 B.n127 585
R320 B.n291 B.n290 585
R321 B.n292 B.n291 585
R322 B.n3 B.n0 585
R323 B.n4 B.n3 585
R324 B.n351 B.n1 585
R325 B.n352 B.n351 585
R326 B.n350 B.n349 585
R327 B.n350 B.n8 585
R328 B.n348 B.n9 585
R329 B.n301 B.n9 585
R330 B.n347 B.n346 585
R331 B.n346 B.n345 585
R332 B.n11 B.n10 585
R333 B.n344 B.n11 585
R334 B.n342 B.n341 585
R335 B.n343 B.n342 585
R336 B.n340 B.n16 585
R337 B.n16 B.n15 585
R338 B.n339 B.n338 585
R339 B.n338 B.n337 585
R340 B.n18 B.n17 585
R341 B.n336 B.n18 585
R342 B.n334 B.n333 585
R343 B.n335 B.n334 585
R344 B.n332 B.n22 585
R345 B.n25 B.n22 585
R346 B.n331 B.n330 585
R347 B.n330 B.n329 585
R348 B.n24 B.n23 585
R349 B.n328 B.n24 585
R350 B.n326 B.n325 585
R351 B.n327 B.n326 585
R352 B.n324 B.n30 585
R353 B.n30 B.n29 585
R354 B.n355 B.n354 585
R355 B.n353 B.n2 585
R356 B.n322 B.n30 540.549
R357 B.n319 B.n51 540.549
R358 B.n176 B.n148 540.549
R359 B.n248 B.n150 540.549
R360 B.n54 B.t10 424.33
R361 B.n52 B.t6 424.33
R362 B.n173 B.t13 424.33
R363 B.n171 B.t17 424.33
R364 B.n320 B.n49 256.663
R365 B.n320 B.n48 256.663
R366 B.n320 B.n47 256.663
R367 B.n320 B.n46 256.663
R368 B.n320 B.n45 256.663
R369 B.n320 B.n44 256.663
R370 B.n320 B.n43 256.663
R371 B.n320 B.n42 256.663
R372 B.n320 B.n41 256.663
R373 B.n320 B.n40 256.663
R374 B.n320 B.n39 256.663
R375 B.n320 B.n38 256.663
R376 B.n320 B.n37 256.663
R377 B.n320 B.n36 256.663
R378 B.n320 B.n35 256.663
R379 B.n320 B.n34 256.663
R380 B.n320 B.n33 256.663
R381 B.n321 B.n320 256.663
R382 B.n247 B.n246 256.663
R383 B.n246 B.n153 256.663
R384 B.n246 B.n154 256.663
R385 B.n246 B.n155 256.663
R386 B.n246 B.n156 256.663
R387 B.n246 B.n157 256.663
R388 B.n246 B.n158 256.663
R389 B.n246 B.n159 256.663
R390 B.n246 B.n160 256.663
R391 B.n246 B.n161 256.663
R392 B.n246 B.n162 256.663
R393 B.n246 B.n163 256.663
R394 B.n246 B.n164 256.663
R395 B.n246 B.n165 256.663
R396 B.n246 B.n166 256.663
R397 B.n246 B.n167 256.663
R398 B.n246 B.n168 256.663
R399 B.n246 B.n169 256.663
R400 B.n357 B.n356 256.663
R401 B.n246 B.n149 174.826
R402 B.n320 B.n29 174.826
R403 B.n57 B.n32 163.367
R404 B.n61 B.n60 163.367
R405 B.n65 B.n64 163.367
R406 B.n69 B.n68 163.367
R407 B.n73 B.n72 163.367
R408 B.n77 B.n76 163.367
R409 B.n81 B.n80 163.367
R410 B.n85 B.n84 163.367
R411 B.n89 B.n88 163.367
R412 B.n93 B.n92 163.367
R413 B.n97 B.n96 163.367
R414 B.n102 B.n101 163.367
R415 B.n106 B.n105 163.367
R416 B.n110 B.n109 163.367
R417 B.n114 B.n113 163.367
R418 B.n118 B.n117 163.367
R419 B.n122 B.n121 163.367
R420 B.n319 B.n50 163.367
R421 B.n254 B.n148 163.367
R422 B.n254 B.n146 163.367
R423 B.n258 B.n146 163.367
R424 B.n258 B.n141 163.367
R425 B.n267 B.n141 163.367
R426 B.n267 B.n139 163.367
R427 B.n271 B.n139 163.367
R428 B.n271 B.n133 163.367
R429 B.n279 B.n133 163.367
R430 B.n279 B.n131 163.367
R431 B.n284 B.n131 163.367
R432 B.n284 B.n126 163.367
R433 B.n293 B.n126 163.367
R434 B.n294 B.n293 163.367
R435 B.n294 B.n5 163.367
R436 B.n6 B.n5 163.367
R437 B.n7 B.n6 163.367
R438 B.n300 B.n7 163.367
R439 B.n302 B.n300 163.367
R440 B.n302 B.n12 163.367
R441 B.n13 B.n12 163.367
R442 B.n14 B.n13 163.367
R443 B.n307 B.n14 163.367
R444 B.n307 B.n19 163.367
R445 B.n20 B.n19 163.367
R446 B.n21 B.n20 163.367
R447 B.n312 B.n21 163.367
R448 B.n312 B.n26 163.367
R449 B.n27 B.n26 163.367
R450 B.n28 B.n27 163.367
R451 B.n51 B.n28 163.367
R452 B.n245 B.n152 163.367
R453 B.n245 B.n170 163.367
R454 B.n241 B.n240 163.367
R455 B.n237 B.n236 163.367
R456 B.n233 B.n232 163.367
R457 B.n229 B.n228 163.367
R458 B.n225 B.n224 163.367
R459 B.n220 B.n219 163.367
R460 B.n216 B.n215 163.367
R461 B.n212 B.n211 163.367
R462 B.n208 B.n207 163.367
R463 B.n204 B.n203 163.367
R464 B.n200 B.n199 163.367
R465 B.n196 B.n195 163.367
R466 B.n192 B.n191 163.367
R467 B.n188 B.n187 163.367
R468 B.n184 B.n183 163.367
R469 B.n180 B.n179 163.367
R470 B.n252 B.n150 163.367
R471 B.n252 B.n144 163.367
R472 B.n261 B.n144 163.367
R473 B.n261 B.n142 163.367
R474 B.n265 B.n142 163.367
R475 B.n265 B.n137 163.367
R476 B.n273 B.n137 163.367
R477 B.n273 B.n135 163.367
R478 B.n277 B.n135 163.367
R479 B.n277 B.n129 163.367
R480 B.n287 B.n129 163.367
R481 B.n287 B.n127 163.367
R482 B.n291 B.n127 163.367
R483 B.n291 B.n3 163.367
R484 B.n355 B.n3 163.367
R485 B.n351 B.n2 163.367
R486 B.n351 B.n350 163.367
R487 B.n350 B.n9 163.367
R488 B.n346 B.n9 163.367
R489 B.n346 B.n11 163.367
R490 B.n342 B.n11 163.367
R491 B.n342 B.n16 163.367
R492 B.n338 B.n16 163.367
R493 B.n338 B.n18 163.367
R494 B.n334 B.n18 163.367
R495 B.n334 B.n22 163.367
R496 B.n330 B.n22 163.367
R497 B.n330 B.n24 163.367
R498 B.n326 B.n24 163.367
R499 B.n326 B.n30 163.367
R500 B.n52 B.t8 136.662
R501 B.n173 B.t16 136.662
R502 B.n54 B.t11 136.662
R503 B.n171 B.t19 136.662
R504 B.n53 B.t9 124.445
R505 B.n174 B.t15 124.445
R506 B.n55 B.t12 124.445
R507 B.n172 B.t18 124.445
R508 B.n253 B.n149 95.1054
R509 B.n253 B.n145 95.1054
R510 B.n260 B.n145 95.1054
R511 B.n260 B.n259 95.1054
R512 B.n266 B.n138 95.1054
R513 B.n272 B.n138 95.1054
R514 B.n272 B.n134 95.1054
R515 B.n278 B.n134 95.1054
R516 B.n286 B.n130 95.1054
R517 B.n292 B.n4 95.1054
R518 B.n354 B.n4 95.1054
R519 B.n354 B.n353 95.1054
R520 B.n353 B.n352 95.1054
R521 B.n352 B.n8 95.1054
R522 B.n345 B.n344 95.1054
R523 B.n343 B.n15 95.1054
R524 B.n337 B.n15 95.1054
R525 B.n337 B.n336 95.1054
R526 B.n336 B.n335 95.1054
R527 B.n329 B.n25 95.1054
R528 B.n329 B.n328 95.1054
R529 B.n328 B.n327 95.1054
R530 B.n327 B.n29 95.1054
R531 B.n285 B.t1 92.3082
R532 B.n301 B.t0 92.3082
R533 B.t2 B.n285 83.9166
R534 B.n301 B.t5 83.9166
R535 B.n266 B.t14 75.525
R536 B.n335 B.t7 75.525
R537 B.n322 B.n321 71.676
R538 B.n57 B.n33 71.676
R539 B.n61 B.n34 71.676
R540 B.n65 B.n35 71.676
R541 B.n69 B.n36 71.676
R542 B.n73 B.n37 71.676
R543 B.n77 B.n38 71.676
R544 B.n81 B.n39 71.676
R545 B.n85 B.n40 71.676
R546 B.n89 B.n41 71.676
R547 B.n93 B.n42 71.676
R548 B.n97 B.n43 71.676
R549 B.n102 B.n44 71.676
R550 B.n106 B.n45 71.676
R551 B.n110 B.n46 71.676
R552 B.n114 B.n47 71.676
R553 B.n118 B.n48 71.676
R554 B.n122 B.n49 71.676
R555 B.n50 B.n49 71.676
R556 B.n121 B.n48 71.676
R557 B.n117 B.n47 71.676
R558 B.n113 B.n46 71.676
R559 B.n109 B.n45 71.676
R560 B.n105 B.n44 71.676
R561 B.n101 B.n43 71.676
R562 B.n96 B.n42 71.676
R563 B.n92 B.n41 71.676
R564 B.n88 B.n40 71.676
R565 B.n84 B.n39 71.676
R566 B.n80 B.n38 71.676
R567 B.n76 B.n37 71.676
R568 B.n72 B.n36 71.676
R569 B.n68 B.n35 71.676
R570 B.n64 B.n34 71.676
R571 B.n60 B.n33 71.676
R572 B.n321 B.n32 71.676
R573 B.n248 B.n247 71.676
R574 B.n170 B.n153 71.676
R575 B.n240 B.n154 71.676
R576 B.n236 B.n155 71.676
R577 B.n232 B.n156 71.676
R578 B.n228 B.n157 71.676
R579 B.n224 B.n158 71.676
R580 B.n219 B.n159 71.676
R581 B.n215 B.n160 71.676
R582 B.n211 B.n161 71.676
R583 B.n207 B.n162 71.676
R584 B.n203 B.n163 71.676
R585 B.n199 B.n164 71.676
R586 B.n195 B.n165 71.676
R587 B.n191 B.n166 71.676
R588 B.n187 B.n167 71.676
R589 B.n183 B.n168 71.676
R590 B.n179 B.n169 71.676
R591 B.n247 B.n152 71.676
R592 B.n241 B.n153 71.676
R593 B.n237 B.n154 71.676
R594 B.n233 B.n155 71.676
R595 B.n229 B.n156 71.676
R596 B.n225 B.n157 71.676
R597 B.n220 B.n158 71.676
R598 B.n216 B.n159 71.676
R599 B.n212 B.n160 71.676
R600 B.n208 B.n161 71.676
R601 B.n204 B.n162 71.676
R602 B.n200 B.n163 71.676
R603 B.n196 B.n164 71.676
R604 B.n192 B.n165 71.676
R605 B.n188 B.n166 71.676
R606 B.n184 B.n167 71.676
R607 B.n180 B.n168 71.676
R608 B.n176 B.n169 71.676
R609 B.n356 B.n355 71.676
R610 B.n356 B.n2 71.676
R611 B.t4 B.n130 69.9306
R612 B.n344 B.t3 69.9306
R613 B.n56 B.n55 59.5399
R614 B.n99 B.n53 59.5399
R615 B.n175 B.n174 59.5399
R616 B.n222 B.n172 59.5399
R617 B.n250 B.n249 35.1225
R618 B.n177 B.n147 35.1225
R619 B.n318 B.n317 35.1225
R620 B.n324 B.n323 35.1225
R621 B.n278 B.t4 25.1753
R622 B.t3 B.n343 25.1753
R623 B.n259 B.t14 19.5809
R624 B.n25 B.t7 19.5809
R625 B B.n357 18.0485
R626 B.n55 B.n54 12.2187
R627 B.n53 B.n52 12.2187
R628 B.n174 B.n173 12.2187
R629 B.n172 B.n171 12.2187
R630 B.n286 B.t2 11.1893
R631 B.n345 B.t5 11.1893
R632 B.n251 B.n250 10.6151
R633 B.n251 B.n143 10.6151
R634 B.n262 B.n143 10.6151
R635 B.n263 B.n262 10.6151
R636 B.n264 B.n263 10.6151
R637 B.n264 B.n136 10.6151
R638 B.n274 B.n136 10.6151
R639 B.n275 B.n274 10.6151
R640 B.n276 B.n275 10.6151
R641 B.n276 B.n128 10.6151
R642 B.n288 B.n128 10.6151
R643 B.n289 B.n288 10.6151
R644 B.n290 B.n289 10.6151
R645 B.n290 B.n0 10.6151
R646 B.n249 B.n151 10.6151
R647 B.n244 B.n151 10.6151
R648 B.n244 B.n243 10.6151
R649 B.n243 B.n242 10.6151
R650 B.n242 B.n239 10.6151
R651 B.n239 B.n238 10.6151
R652 B.n238 B.n235 10.6151
R653 B.n235 B.n234 10.6151
R654 B.n234 B.n231 10.6151
R655 B.n231 B.n230 10.6151
R656 B.n230 B.n227 10.6151
R657 B.n227 B.n226 10.6151
R658 B.n226 B.n223 10.6151
R659 B.n221 B.n218 10.6151
R660 B.n218 B.n217 10.6151
R661 B.n217 B.n214 10.6151
R662 B.n214 B.n213 10.6151
R663 B.n213 B.n210 10.6151
R664 B.n210 B.n209 10.6151
R665 B.n209 B.n206 10.6151
R666 B.n206 B.n205 10.6151
R667 B.n202 B.n201 10.6151
R668 B.n201 B.n198 10.6151
R669 B.n198 B.n197 10.6151
R670 B.n197 B.n194 10.6151
R671 B.n194 B.n193 10.6151
R672 B.n193 B.n190 10.6151
R673 B.n190 B.n189 10.6151
R674 B.n189 B.n186 10.6151
R675 B.n186 B.n185 10.6151
R676 B.n185 B.n182 10.6151
R677 B.n182 B.n181 10.6151
R678 B.n181 B.n178 10.6151
R679 B.n178 B.n177 10.6151
R680 B.n255 B.n147 10.6151
R681 B.n256 B.n255 10.6151
R682 B.n257 B.n256 10.6151
R683 B.n257 B.n140 10.6151
R684 B.n268 B.n140 10.6151
R685 B.n269 B.n268 10.6151
R686 B.n270 B.n269 10.6151
R687 B.n270 B.n132 10.6151
R688 B.n280 B.n132 10.6151
R689 B.n281 B.n280 10.6151
R690 B.n283 B.n281 10.6151
R691 B.n283 B.n282 10.6151
R692 B.n282 B.n125 10.6151
R693 B.n295 B.n125 10.6151
R694 B.n296 B.n295 10.6151
R695 B.n297 B.n296 10.6151
R696 B.n298 B.n297 10.6151
R697 B.n299 B.n298 10.6151
R698 B.n303 B.n299 10.6151
R699 B.n304 B.n303 10.6151
R700 B.n305 B.n304 10.6151
R701 B.n306 B.n305 10.6151
R702 B.n308 B.n306 10.6151
R703 B.n309 B.n308 10.6151
R704 B.n310 B.n309 10.6151
R705 B.n311 B.n310 10.6151
R706 B.n313 B.n311 10.6151
R707 B.n314 B.n313 10.6151
R708 B.n315 B.n314 10.6151
R709 B.n316 B.n315 10.6151
R710 B.n317 B.n316 10.6151
R711 B.n349 B.n1 10.6151
R712 B.n349 B.n348 10.6151
R713 B.n348 B.n347 10.6151
R714 B.n347 B.n10 10.6151
R715 B.n341 B.n10 10.6151
R716 B.n341 B.n340 10.6151
R717 B.n340 B.n339 10.6151
R718 B.n339 B.n17 10.6151
R719 B.n333 B.n17 10.6151
R720 B.n333 B.n332 10.6151
R721 B.n332 B.n331 10.6151
R722 B.n331 B.n23 10.6151
R723 B.n325 B.n23 10.6151
R724 B.n325 B.n324 10.6151
R725 B.n323 B.n31 10.6151
R726 B.n58 B.n31 10.6151
R727 B.n59 B.n58 10.6151
R728 B.n62 B.n59 10.6151
R729 B.n63 B.n62 10.6151
R730 B.n66 B.n63 10.6151
R731 B.n67 B.n66 10.6151
R732 B.n70 B.n67 10.6151
R733 B.n71 B.n70 10.6151
R734 B.n74 B.n71 10.6151
R735 B.n75 B.n74 10.6151
R736 B.n78 B.n75 10.6151
R737 B.n79 B.n78 10.6151
R738 B.n83 B.n82 10.6151
R739 B.n86 B.n83 10.6151
R740 B.n87 B.n86 10.6151
R741 B.n90 B.n87 10.6151
R742 B.n91 B.n90 10.6151
R743 B.n94 B.n91 10.6151
R744 B.n95 B.n94 10.6151
R745 B.n98 B.n95 10.6151
R746 B.n103 B.n100 10.6151
R747 B.n104 B.n103 10.6151
R748 B.n107 B.n104 10.6151
R749 B.n108 B.n107 10.6151
R750 B.n111 B.n108 10.6151
R751 B.n112 B.n111 10.6151
R752 B.n115 B.n112 10.6151
R753 B.n116 B.n115 10.6151
R754 B.n119 B.n116 10.6151
R755 B.n120 B.n119 10.6151
R756 B.n123 B.n120 10.6151
R757 B.n124 B.n123 10.6151
R758 B.n318 B.n124 10.6151
R759 B.n357 B.n0 8.11757
R760 B.n357 B.n1 8.11757
R761 B.n222 B.n221 6.5566
R762 B.n205 B.n175 6.5566
R763 B.n82 B.n56 6.5566
R764 B.n99 B.n98 6.5566
R765 B.n223 B.n222 4.05904
R766 B.n202 B.n175 4.05904
R767 B.n79 B.n56 4.05904
R768 B.n100 B.n99 4.05904
R769 B.n292 B.t1 2.7977
R770 B.t0 B.n8 2.7977
R771 VN.n2 VN.t3 368.803
R772 VN.n0 VN.t1 368.803
R773 VN.n6 VN.t0 368.803
R774 VN.n4 VN.t2 368.803
R775 VN.n1 VN.t4 313.3
R776 VN.n5 VN.t5 313.3
R777 VN.n7 VN.n4 161.489
R778 VN.n3 VN.n0 161.489
R779 VN.n3 VN.n2 161.3
R780 VN.n7 VN.n6 161.3
R781 VN.n1 VN.n0 36.5157
R782 VN.n2 VN.n1 36.5157
R783 VN.n6 VN.n5 36.5157
R784 VN.n5 VN.n4 36.5157
R785 VN VN.n7 33.0516
R786 VN VN.n3 0.0516364
R787 VDD2.n19 VDD2.n13 289.615
R788 VDD2.n6 VDD2.n0 289.615
R789 VDD2.n20 VDD2.n19 185
R790 VDD2.n18 VDD2.n17 185
R791 VDD2.n5 VDD2.n4 185
R792 VDD2.n7 VDD2.n6 185
R793 VDD2.n16 VDD2.t5 151.613
R794 VDD2.n3 VDD2.t4 151.613
R795 VDD2.n19 VDD2.n18 104.615
R796 VDD2.n6 VDD2.n5 104.615
R797 VDD2.n12 VDD2.n11 88.7245
R798 VDD2 VDD2.n25 88.7216
R799 VDD2.n12 VDD2.n10 52.901
R800 VDD2.n24 VDD2.n23 52.549
R801 VDD2.n18 VDD2.t5 52.3082
R802 VDD2.n5 VDD2.t4 52.3082
R803 VDD2.n24 VDD2.n12 27.7131
R804 VDD2.n17 VDD2.n16 15.3979
R805 VDD2.n4 VDD2.n3 15.3979
R806 VDD2.n20 VDD2.n15 12.8005
R807 VDD2.n7 VDD2.n2 12.8005
R808 VDD2.n21 VDD2.n13 12.0247
R809 VDD2.n8 VDD2.n0 12.0247
R810 VDD2.n23 VDD2.n22 9.45567
R811 VDD2.n10 VDD2.n9 9.45567
R812 VDD2.n22 VDD2.n21 9.3005
R813 VDD2.n15 VDD2.n14 9.3005
R814 VDD2.n9 VDD2.n8 9.3005
R815 VDD2.n2 VDD2.n1 9.3005
R816 VDD2.n25 VDD2.t0 7.64529
R817 VDD2.n25 VDD2.t3 7.64529
R818 VDD2.n11 VDD2.t1 7.64529
R819 VDD2.n11 VDD2.t2 7.64529
R820 VDD2.n16 VDD2.n14 4.69785
R821 VDD2.n3 VDD2.n1 4.69785
R822 VDD2.n23 VDD2.n13 1.93989
R823 VDD2.n10 VDD2.n0 1.93989
R824 VDD2.n21 VDD2.n20 1.16414
R825 VDD2.n8 VDD2.n7 1.16414
R826 VDD2 VDD2.n24 0.466017
R827 VDD2.n17 VDD2.n15 0.388379
R828 VDD2.n4 VDD2.n2 0.388379
R829 VDD2.n22 VDD2.n14 0.155672
R830 VDD2.n9 VDD2.n1 0.155672
C0 VN VTAIL 0.838226f
C1 VDD1 VP 0.942851f
C2 VDD2 VTAIL 4.29656f
C3 VDD2 VN 0.829413f
C4 VDD1 VTAIL 4.26031f
C5 VDD1 VN 0.153029f
C6 VTAIL VP 0.852474f
C7 VN VP 2.95235f
C8 VDD1 VDD2 0.566287f
C9 VDD2 VP 0.268193f
C10 VDD2 B 2.418909f
C11 VDD1 B 2.428163f
C12 VTAIL B 2.538773f
C13 VN B 4.887461f
C14 VP B 3.794935f
C15 VDD2.n0 B 0.031235f
C16 VDD2.n1 B 0.174666f
C17 VDD2.n2 B 0.011999f
C18 VDD2.t4 B 0.049864f
C19 VDD2.n3 B 0.080937f
C20 VDD2.n4 B 0.016054f
C21 VDD2.n5 B 0.021271f
C22 VDD2.n6 B 0.06113f
C23 VDD2.n7 B 0.012705f
C24 VDD2.n8 B 0.011999f
C25 VDD2.n9 B 0.057409f
C26 VDD2.n10 B 0.050211f
C27 VDD2.t1 B 0.045702f
C28 VDD2.t2 B 0.045702f
C29 VDD2.n11 B 0.325521f
C30 VDD2.n12 B 0.996968f
C31 VDD2.n13 B 0.031235f
C32 VDD2.n14 B 0.174666f
C33 VDD2.n15 B 0.011999f
C34 VDD2.t5 B 0.049864f
C35 VDD2.n16 B 0.080937f
C36 VDD2.n17 B 0.016054f
C37 VDD2.n18 B 0.021271f
C38 VDD2.n19 B 0.06113f
C39 VDD2.n20 B 0.012705f
C40 VDD2.n21 B 0.011999f
C41 VDD2.n22 B 0.057409f
C42 VDD2.n23 B 0.049725f
C43 VDD2.n24 B 1.05182f
C44 VDD2.t0 B 0.045702f
C45 VDD2.t3 B 0.045702f
C46 VDD2.n25 B 0.325508f
C47 VN.t1 B 0.092043f
C48 VN.n0 B 0.06272f
C49 VN.t4 B 0.083637f
C50 VN.n1 B 0.051756f
C51 VN.t3 B 0.092043f
C52 VN.n2 B 0.062662f
C53 VN.n3 B 0.078254f
C54 VN.t2 B 0.092043f
C55 VN.n4 B 0.06272f
C56 VN.t0 B 0.092043f
C57 VN.t5 B 0.083637f
C58 VN.n5 B 0.051756f
C59 VN.n6 B 0.062662f
C60 VN.n7 B 1.03354f
C61 VDD1.n0 B 0.030648f
C62 VDD1.n1 B 0.171379f
C63 VDD1.n2 B 0.011773f
C64 VDD1.t4 B 0.048926f
C65 VDD1.n3 B 0.079414f
C66 VDD1.n4 B 0.015752f
C67 VDD1.n5 B 0.020871f
C68 VDD1.n6 B 0.05998f
C69 VDD1.n7 B 0.012466f
C70 VDD1.n8 B 0.011773f
C71 VDD1.n9 B 0.056329f
C72 VDD1.n10 B 0.049477f
C73 VDD1.n11 B 0.030648f
C74 VDD1.n12 B 0.171379f
C75 VDD1.n13 B 0.011773f
C76 VDD1.t2 B 0.048926f
C77 VDD1.n14 B 0.079414f
C78 VDD1.n15 B 0.015752f
C79 VDD1.n16 B 0.020871f
C80 VDD1.n17 B 0.05998f
C81 VDD1.n18 B 0.012466f
C82 VDD1.n19 B 0.011773f
C83 VDD1.n20 B 0.056329f
C84 VDD1.n21 B 0.049266f
C85 VDD1.t1 B 0.044842f
C86 VDD1.t5 B 0.044842f
C87 VDD1.n22 B 0.319395f
C88 VDD1.n23 B 1.03513f
C89 VDD1.t3 B 0.044842f
C90 VDD1.t0 B 0.044842f
C91 VDD1.n24 B 0.319193f
C92 VDD1.n25 B 1.19359f
C93 VTAIL.t0 B 0.054808f
C94 VTAIL.t9 B 0.054808f
C95 VTAIL.n0 B 0.345079f
C96 VTAIL.n1 B 0.288878f
C97 VTAIL.n2 B 0.037459f
C98 VTAIL.n3 B 0.209469f
C99 VTAIL.n4 B 0.01439f
C100 VTAIL.t6 B 0.0598f
C101 VTAIL.n5 B 0.097064f
C102 VTAIL.n6 B 0.019253f
C103 VTAIL.n7 B 0.025509f
C104 VTAIL.n8 B 0.073311f
C105 VTAIL.n9 B 0.015236f
C106 VTAIL.n10 B 0.01439f
C107 VTAIL.n11 B 0.068849f
C108 VTAIL.n12 B 0.041191f
C109 VTAIL.n13 B 0.137639f
C110 VTAIL.t3 B 0.054808f
C111 VTAIL.t7 B 0.054808f
C112 VTAIL.n14 B 0.345079f
C113 VTAIL.n15 B 0.905176f
C114 VTAIL.t11 B 0.054808f
C115 VTAIL.t2 B 0.054808f
C116 VTAIL.n16 B 0.345081f
C117 VTAIL.n17 B 0.905174f
C118 VTAIL.n18 B 0.037459f
C119 VTAIL.n19 B 0.209469f
C120 VTAIL.n20 B 0.01439f
C121 VTAIL.t1 B 0.0598f
C122 VTAIL.n21 B 0.097064f
C123 VTAIL.n22 B 0.019253f
C124 VTAIL.n23 B 0.025509f
C125 VTAIL.n24 B 0.073311f
C126 VTAIL.n25 B 0.015236f
C127 VTAIL.n26 B 0.01439f
C128 VTAIL.n27 B 0.068849f
C129 VTAIL.n28 B 0.041191f
C130 VTAIL.n29 B 0.137639f
C131 VTAIL.t4 B 0.054808f
C132 VTAIL.t5 B 0.054808f
C133 VTAIL.n30 B 0.345081f
C134 VTAIL.n31 B 0.319002f
C135 VTAIL.n32 B 0.037459f
C136 VTAIL.n33 B 0.209469f
C137 VTAIL.n34 B 0.01439f
C138 VTAIL.t8 B 0.0598f
C139 VTAIL.n35 B 0.097064f
C140 VTAIL.n36 B 0.019253f
C141 VTAIL.n37 B 0.025509f
C142 VTAIL.n38 B 0.073311f
C143 VTAIL.n39 B 0.015236f
C144 VTAIL.n40 B 0.01439f
C145 VTAIL.n41 B 0.068849f
C146 VTAIL.n42 B 0.041191f
C147 VTAIL.n43 B 0.676947f
C148 VTAIL.n44 B 0.037459f
C149 VTAIL.n45 B 0.209469f
C150 VTAIL.n46 B 0.01439f
C151 VTAIL.t10 B 0.0598f
C152 VTAIL.n47 B 0.097064f
C153 VTAIL.n48 B 0.019253f
C154 VTAIL.n49 B 0.025509f
C155 VTAIL.n50 B 0.073311f
C156 VTAIL.n51 B 0.015236f
C157 VTAIL.n52 B 0.01439f
C158 VTAIL.n53 B 0.068849f
C159 VTAIL.n54 B 0.041191f
C160 VTAIL.n55 B 0.66021f
C161 VP.t1 B 0.093664f
C162 VP.n0 B 0.063825f
C163 VP.t2 B 0.08511f
C164 VP.n1 B 0.052667f
C165 VP.t5 B 0.093664f
C166 VP.n2 B 0.063766f
C167 VP.n3 B 1.02663f
C168 VP.n4 B 1.01748f
C169 VP.t4 B 0.08511f
C170 VP.t3 B 0.093664f
C171 VP.n5 B 0.063766f
C172 VP.n6 B 0.052667f
C173 VP.t0 B 0.093664f
C174 VP.n7 B 0.063766f
C175 VP.n8 B 0.029128f
.ends

