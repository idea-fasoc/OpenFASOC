* NGSPICE file created from diff_pair_sample_1559.ext - technology: sky130A

.subckt diff_pair_sample_1559 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t9 VN.t0 VTAIL.t10 w_n4786_n3892# sky130_fd_pr__pfet_01v8 ad=2.4123 pd=14.95 as=2.4123 ps=14.95 w=14.62 l=2.85
X1 B.t11 B.t9 B.t10 w_n4786_n3892# sky130_fd_pr__pfet_01v8 ad=5.7018 pd=30.02 as=0 ps=0 w=14.62 l=2.85
X2 VDD1.t9 VP.t0 VTAIL.t4 w_n4786_n3892# sky130_fd_pr__pfet_01v8 ad=2.4123 pd=14.95 as=2.4123 ps=14.95 w=14.62 l=2.85
X3 VTAIL.t12 VN.t1 VDD2.t8 w_n4786_n3892# sky130_fd_pr__pfet_01v8 ad=2.4123 pd=14.95 as=2.4123 ps=14.95 w=14.62 l=2.85
X4 VDD1.t8 VP.t1 VTAIL.t8 w_n4786_n3892# sky130_fd_pr__pfet_01v8 ad=5.7018 pd=30.02 as=2.4123 ps=14.95 w=14.62 l=2.85
X5 VDD1.t7 VP.t2 VTAIL.t7 w_n4786_n3892# sky130_fd_pr__pfet_01v8 ad=5.7018 pd=30.02 as=2.4123 ps=14.95 w=14.62 l=2.85
X6 VTAIL.t6 VP.t3 VDD1.t6 w_n4786_n3892# sky130_fd_pr__pfet_01v8 ad=2.4123 pd=14.95 as=2.4123 ps=14.95 w=14.62 l=2.85
X7 VTAIL.t11 VN.t2 VDD2.t7 w_n4786_n3892# sky130_fd_pr__pfet_01v8 ad=2.4123 pd=14.95 as=2.4123 ps=14.95 w=14.62 l=2.85
X8 VDD2.t6 VN.t3 VTAIL.t15 w_n4786_n3892# sky130_fd_pr__pfet_01v8 ad=2.4123 pd=14.95 as=5.7018 ps=30.02 w=14.62 l=2.85
X9 VDD2.t5 VN.t4 VTAIL.t14 w_n4786_n3892# sky130_fd_pr__pfet_01v8 ad=5.7018 pd=30.02 as=2.4123 ps=14.95 w=14.62 l=2.85
X10 VDD2.t4 VN.t5 VTAIL.t18 w_n4786_n3892# sky130_fd_pr__pfet_01v8 ad=5.7018 pd=30.02 as=2.4123 ps=14.95 w=14.62 l=2.85
X11 B.t8 B.t6 B.t7 w_n4786_n3892# sky130_fd_pr__pfet_01v8 ad=5.7018 pd=30.02 as=0 ps=0 w=14.62 l=2.85
X12 VTAIL.t5 VP.t4 VDD1.t5 w_n4786_n3892# sky130_fd_pr__pfet_01v8 ad=2.4123 pd=14.95 as=2.4123 ps=14.95 w=14.62 l=2.85
X13 VTAIL.t3 VP.t5 VDD1.t4 w_n4786_n3892# sky130_fd_pr__pfet_01v8 ad=2.4123 pd=14.95 as=2.4123 ps=14.95 w=14.62 l=2.85
X14 VDD1.t3 VP.t6 VTAIL.t9 w_n4786_n3892# sky130_fd_pr__pfet_01v8 ad=2.4123 pd=14.95 as=2.4123 ps=14.95 w=14.62 l=2.85
X15 VDD2.t3 VN.t6 VTAIL.t17 w_n4786_n3892# sky130_fd_pr__pfet_01v8 ad=2.4123 pd=14.95 as=2.4123 ps=14.95 w=14.62 l=2.85
X16 VDD2.t2 VN.t7 VTAIL.t19 w_n4786_n3892# sky130_fd_pr__pfet_01v8 ad=2.4123 pd=14.95 as=5.7018 ps=30.02 w=14.62 l=2.85
X17 B.t5 B.t3 B.t4 w_n4786_n3892# sky130_fd_pr__pfet_01v8 ad=5.7018 pd=30.02 as=0 ps=0 w=14.62 l=2.85
X18 VDD1.t2 VP.t7 VTAIL.t1 w_n4786_n3892# sky130_fd_pr__pfet_01v8 ad=2.4123 pd=14.95 as=5.7018 ps=30.02 w=14.62 l=2.85
X19 VTAIL.t2 VP.t8 VDD1.t1 w_n4786_n3892# sky130_fd_pr__pfet_01v8 ad=2.4123 pd=14.95 as=2.4123 ps=14.95 w=14.62 l=2.85
X20 VTAIL.t16 VN.t8 VDD2.t1 w_n4786_n3892# sky130_fd_pr__pfet_01v8 ad=2.4123 pd=14.95 as=2.4123 ps=14.95 w=14.62 l=2.85
X21 B.t2 B.t0 B.t1 w_n4786_n3892# sky130_fd_pr__pfet_01v8 ad=5.7018 pd=30.02 as=0 ps=0 w=14.62 l=2.85
X22 VTAIL.t13 VN.t9 VDD2.t0 w_n4786_n3892# sky130_fd_pr__pfet_01v8 ad=2.4123 pd=14.95 as=2.4123 ps=14.95 w=14.62 l=2.85
X23 VDD1.t0 VP.t9 VTAIL.t0 w_n4786_n3892# sky130_fd_pr__pfet_01v8 ad=2.4123 pd=14.95 as=5.7018 ps=30.02 w=14.62 l=2.85
R0 VN.n85 VN.n44 161.3
R1 VN.n84 VN.n83 161.3
R2 VN.n82 VN.n45 161.3
R3 VN.n81 VN.n80 161.3
R4 VN.n79 VN.n46 161.3
R5 VN.n78 VN.n77 161.3
R6 VN.n76 VN.n47 161.3
R7 VN.n75 VN.n74 161.3
R8 VN.n73 VN.n48 161.3
R9 VN.n72 VN.n71 161.3
R10 VN.n70 VN.n50 161.3
R11 VN.n69 VN.n68 161.3
R12 VN.n67 VN.n51 161.3
R13 VN.n65 VN.n64 161.3
R14 VN.n63 VN.n52 161.3
R15 VN.n62 VN.n61 161.3
R16 VN.n60 VN.n53 161.3
R17 VN.n59 VN.n58 161.3
R18 VN.n57 VN.n54 161.3
R19 VN.n41 VN.n0 161.3
R20 VN.n40 VN.n39 161.3
R21 VN.n38 VN.n1 161.3
R22 VN.n37 VN.n36 161.3
R23 VN.n35 VN.n2 161.3
R24 VN.n34 VN.n33 161.3
R25 VN.n32 VN.n3 161.3
R26 VN.n31 VN.n30 161.3
R27 VN.n28 VN.n4 161.3
R28 VN.n27 VN.n26 161.3
R29 VN.n25 VN.n5 161.3
R30 VN.n24 VN.n23 161.3
R31 VN.n22 VN.n6 161.3
R32 VN.n20 VN.n19 161.3
R33 VN.n18 VN.n7 161.3
R34 VN.n17 VN.n16 161.3
R35 VN.n15 VN.n8 161.3
R36 VN.n14 VN.n13 161.3
R37 VN.n12 VN.n9 161.3
R38 VN.n11 VN.t4 157.819
R39 VN.n56 VN.t3 157.819
R40 VN.n10 VN.t2 123.629
R41 VN.n21 VN.t0 123.629
R42 VN.n29 VN.t1 123.629
R43 VN.n42 VN.t7 123.629
R44 VN.n55 VN.t8 123.629
R45 VN.n66 VN.t6 123.629
R46 VN.n49 VN.t9 123.629
R47 VN.n86 VN.t5 123.629
R48 VN.n43 VN.n42 105.499
R49 VN.n87 VN.n86 105.499
R50 VN VN.n87 56.7482
R51 VN.n16 VN.n15 56.0773
R52 VN.n27 VN.n5 56.0773
R53 VN.n61 VN.n60 56.0773
R54 VN.n72 VN.n50 56.0773
R55 VN.n11 VN.n10 52.6217
R56 VN.n56 VN.n55 52.6217
R57 VN.n36 VN.n1 42.5146
R58 VN.n80 VN.n45 42.5146
R59 VN.n36 VN.n35 38.6395
R60 VN.n80 VN.n79 38.6395
R61 VN.n15 VN.n14 25.0767
R62 VN.n28 VN.n27 25.0767
R63 VN.n60 VN.n59 25.0767
R64 VN.n73 VN.n72 25.0767
R65 VN.n14 VN.n9 24.5923
R66 VN.n16 VN.n7 24.5923
R67 VN.n20 VN.n7 24.5923
R68 VN.n23 VN.n22 24.5923
R69 VN.n23 VN.n5 24.5923
R70 VN.n30 VN.n28 24.5923
R71 VN.n34 VN.n3 24.5923
R72 VN.n35 VN.n34 24.5923
R73 VN.n40 VN.n1 24.5923
R74 VN.n41 VN.n40 24.5923
R75 VN.n59 VN.n54 24.5923
R76 VN.n68 VN.n50 24.5923
R77 VN.n68 VN.n67 24.5923
R78 VN.n65 VN.n52 24.5923
R79 VN.n61 VN.n52 24.5923
R80 VN.n79 VN.n78 24.5923
R81 VN.n78 VN.n47 24.5923
R82 VN.n74 VN.n73 24.5923
R83 VN.n85 VN.n84 24.5923
R84 VN.n84 VN.n45 24.5923
R85 VN.n10 VN.n9 21.1495
R86 VN.n30 VN.n29 21.1495
R87 VN.n55 VN.n54 21.1495
R88 VN.n74 VN.n49 21.1495
R89 VN.n21 VN.n20 12.2964
R90 VN.n22 VN.n21 12.2964
R91 VN.n67 VN.n66 12.2964
R92 VN.n66 VN.n65 12.2964
R93 VN.n42 VN.n41 5.4107
R94 VN.n86 VN.n85 5.4107
R95 VN.n57 VN.n56 4.94439
R96 VN.n12 VN.n11 4.94439
R97 VN.n29 VN.n3 3.44336
R98 VN.n49 VN.n47 3.44336
R99 VN.n87 VN.n44 0.278335
R100 VN.n43 VN.n0 0.278335
R101 VN.n83 VN.n44 0.189894
R102 VN.n83 VN.n82 0.189894
R103 VN.n82 VN.n81 0.189894
R104 VN.n81 VN.n46 0.189894
R105 VN.n77 VN.n46 0.189894
R106 VN.n77 VN.n76 0.189894
R107 VN.n76 VN.n75 0.189894
R108 VN.n75 VN.n48 0.189894
R109 VN.n71 VN.n48 0.189894
R110 VN.n71 VN.n70 0.189894
R111 VN.n70 VN.n69 0.189894
R112 VN.n69 VN.n51 0.189894
R113 VN.n64 VN.n51 0.189894
R114 VN.n64 VN.n63 0.189894
R115 VN.n63 VN.n62 0.189894
R116 VN.n62 VN.n53 0.189894
R117 VN.n58 VN.n53 0.189894
R118 VN.n58 VN.n57 0.189894
R119 VN.n13 VN.n12 0.189894
R120 VN.n13 VN.n8 0.189894
R121 VN.n17 VN.n8 0.189894
R122 VN.n18 VN.n17 0.189894
R123 VN.n19 VN.n18 0.189894
R124 VN.n19 VN.n6 0.189894
R125 VN.n24 VN.n6 0.189894
R126 VN.n25 VN.n24 0.189894
R127 VN.n26 VN.n25 0.189894
R128 VN.n26 VN.n4 0.189894
R129 VN.n31 VN.n4 0.189894
R130 VN.n32 VN.n31 0.189894
R131 VN.n33 VN.n32 0.189894
R132 VN.n33 VN.n2 0.189894
R133 VN.n37 VN.n2 0.189894
R134 VN.n38 VN.n37 0.189894
R135 VN.n39 VN.n38 0.189894
R136 VN.n39 VN.n0 0.189894
R137 VN VN.n43 0.153485
R138 VTAIL.n11 VTAIL.t15 56.4926
R139 VTAIL.n16 VTAIL.t1 56.4925
R140 VTAIL.n17 VTAIL.t19 56.4923
R141 VTAIL.n2 VTAIL.t0 56.4923
R142 VTAIL.n15 VTAIL.n14 54.2692
R143 VTAIL.n13 VTAIL.n12 54.2692
R144 VTAIL.n10 VTAIL.n9 54.2692
R145 VTAIL.n8 VTAIL.n7 54.2692
R146 VTAIL.n19 VTAIL.n18 54.2692
R147 VTAIL.n1 VTAIL.n0 54.2692
R148 VTAIL.n4 VTAIL.n3 54.2692
R149 VTAIL.n6 VTAIL.n5 54.2692
R150 VTAIL.n8 VTAIL.n6 30.4531
R151 VTAIL.n17 VTAIL.n16 27.7117
R152 VTAIL.n10 VTAIL.n8 2.74188
R153 VTAIL.n11 VTAIL.n10 2.74188
R154 VTAIL.n15 VTAIL.n13 2.74188
R155 VTAIL.n16 VTAIL.n15 2.74188
R156 VTAIL.n6 VTAIL.n4 2.74188
R157 VTAIL.n4 VTAIL.n2 2.74188
R158 VTAIL.n19 VTAIL.n17 2.74188
R159 VTAIL.n18 VTAIL.t10 2.22382
R160 VTAIL.n18 VTAIL.t12 2.22382
R161 VTAIL.n0 VTAIL.t14 2.22382
R162 VTAIL.n0 VTAIL.t11 2.22382
R163 VTAIL.n3 VTAIL.t9 2.22382
R164 VTAIL.n3 VTAIL.t2 2.22382
R165 VTAIL.n5 VTAIL.t8 2.22382
R166 VTAIL.n5 VTAIL.t6 2.22382
R167 VTAIL.n14 VTAIL.t4 2.22382
R168 VTAIL.n14 VTAIL.t5 2.22382
R169 VTAIL.n12 VTAIL.t7 2.22382
R170 VTAIL.n12 VTAIL.t3 2.22382
R171 VTAIL.n9 VTAIL.t17 2.22382
R172 VTAIL.n9 VTAIL.t16 2.22382
R173 VTAIL.n7 VTAIL.t18 2.22382
R174 VTAIL.n7 VTAIL.t13 2.22382
R175 VTAIL VTAIL.n1 2.11472
R176 VTAIL.n13 VTAIL.n11 1.84102
R177 VTAIL.n2 VTAIL.n1 1.84102
R178 VTAIL VTAIL.n19 0.627655
R179 VDD2.n1 VDD2.t5 75.9125
R180 VDD2.n4 VDD2.t4 73.1714
R181 VDD2.n3 VDD2.n2 72.9487
R182 VDD2 VDD2.n7 72.9459
R183 VDD2.n6 VDD2.n5 70.948
R184 VDD2.n1 VDD2.n0 70.948
R185 VDD2.n4 VDD2.n3 49.3403
R186 VDD2.n6 VDD2.n4 2.74188
R187 VDD2.n7 VDD2.t1 2.22382
R188 VDD2.n7 VDD2.t6 2.22382
R189 VDD2.n5 VDD2.t0 2.22382
R190 VDD2.n5 VDD2.t3 2.22382
R191 VDD2.n2 VDD2.t8 2.22382
R192 VDD2.n2 VDD2.t2 2.22382
R193 VDD2.n0 VDD2.t7 2.22382
R194 VDD2.n0 VDD2.t9 2.22382
R195 VDD2 VDD2.n6 0.744035
R196 VDD2.n3 VDD2.n1 0.630499
R197 B.n700 B.n699 585
R198 B.n701 B.n92 585
R199 B.n703 B.n702 585
R200 B.n704 B.n91 585
R201 B.n706 B.n705 585
R202 B.n707 B.n90 585
R203 B.n709 B.n708 585
R204 B.n710 B.n89 585
R205 B.n712 B.n711 585
R206 B.n713 B.n88 585
R207 B.n715 B.n714 585
R208 B.n716 B.n87 585
R209 B.n718 B.n717 585
R210 B.n719 B.n86 585
R211 B.n721 B.n720 585
R212 B.n722 B.n85 585
R213 B.n724 B.n723 585
R214 B.n725 B.n84 585
R215 B.n727 B.n726 585
R216 B.n728 B.n83 585
R217 B.n730 B.n729 585
R218 B.n731 B.n82 585
R219 B.n733 B.n732 585
R220 B.n734 B.n81 585
R221 B.n736 B.n735 585
R222 B.n737 B.n80 585
R223 B.n739 B.n738 585
R224 B.n740 B.n79 585
R225 B.n742 B.n741 585
R226 B.n743 B.n78 585
R227 B.n745 B.n744 585
R228 B.n746 B.n77 585
R229 B.n748 B.n747 585
R230 B.n749 B.n76 585
R231 B.n751 B.n750 585
R232 B.n752 B.n75 585
R233 B.n754 B.n753 585
R234 B.n755 B.n74 585
R235 B.n757 B.n756 585
R236 B.n758 B.n73 585
R237 B.n760 B.n759 585
R238 B.n761 B.n72 585
R239 B.n763 B.n762 585
R240 B.n764 B.n71 585
R241 B.n766 B.n765 585
R242 B.n767 B.n70 585
R243 B.n769 B.n768 585
R244 B.n770 B.n69 585
R245 B.n772 B.n771 585
R246 B.n774 B.n66 585
R247 B.n776 B.n775 585
R248 B.n777 B.n65 585
R249 B.n779 B.n778 585
R250 B.n780 B.n64 585
R251 B.n782 B.n781 585
R252 B.n783 B.n63 585
R253 B.n785 B.n784 585
R254 B.n786 B.n59 585
R255 B.n788 B.n787 585
R256 B.n789 B.n58 585
R257 B.n791 B.n790 585
R258 B.n792 B.n57 585
R259 B.n794 B.n793 585
R260 B.n795 B.n56 585
R261 B.n797 B.n796 585
R262 B.n798 B.n55 585
R263 B.n800 B.n799 585
R264 B.n801 B.n54 585
R265 B.n803 B.n802 585
R266 B.n804 B.n53 585
R267 B.n806 B.n805 585
R268 B.n807 B.n52 585
R269 B.n809 B.n808 585
R270 B.n810 B.n51 585
R271 B.n812 B.n811 585
R272 B.n813 B.n50 585
R273 B.n815 B.n814 585
R274 B.n816 B.n49 585
R275 B.n818 B.n817 585
R276 B.n819 B.n48 585
R277 B.n821 B.n820 585
R278 B.n822 B.n47 585
R279 B.n824 B.n823 585
R280 B.n825 B.n46 585
R281 B.n827 B.n826 585
R282 B.n828 B.n45 585
R283 B.n830 B.n829 585
R284 B.n831 B.n44 585
R285 B.n833 B.n832 585
R286 B.n834 B.n43 585
R287 B.n836 B.n835 585
R288 B.n837 B.n42 585
R289 B.n839 B.n838 585
R290 B.n840 B.n41 585
R291 B.n842 B.n841 585
R292 B.n843 B.n40 585
R293 B.n845 B.n844 585
R294 B.n846 B.n39 585
R295 B.n848 B.n847 585
R296 B.n849 B.n38 585
R297 B.n851 B.n850 585
R298 B.n852 B.n37 585
R299 B.n854 B.n853 585
R300 B.n855 B.n36 585
R301 B.n857 B.n856 585
R302 B.n858 B.n35 585
R303 B.n860 B.n859 585
R304 B.n861 B.n34 585
R305 B.n698 B.n93 585
R306 B.n697 B.n696 585
R307 B.n695 B.n94 585
R308 B.n694 B.n693 585
R309 B.n692 B.n95 585
R310 B.n691 B.n690 585
R311 B.n689 B.n96 585
R312 B.n688 B.n687 585
R313 B.n686 B.n97 585
R314 B.n685 B.n684 585
R315 B.n683 B.n98 585
R316 B.n682 B.n681 585
R317 B.n680 B.n99 585
R318 B.n679 B.n678 585
R319 B.n677 B.n100 585
R320 B.n676 B.n675 585
R321 B.n674 B.n101 585
R322 B.n673 B.n672 585
R323 B.n671 B.n102 585
R324 B.n670 B.n669 585
R325 B.n668 B.n103 585
R326 B.n667 B.n666 585
R327 B.n665 B.n104 585
R328 B.n664 B.n663 585
R329 B.n662 B.n105 585
R330 B.n661 B.n660 585
R331 B.n659 B.n106 585
R332 B.n658 B.n657 585
R333 B.n656 B.n107 585
R334 B.n655 B.n654 585
R335 B.n653 B.n108 585
R336 B.n652 B.n651 585
R337 B.n650 B.n109 585
R338 B.n649 B.n648 585
R339 B.n647 B.n110 585
R340 B.n646 B.n645 585
R341 B.n644 B.n111 585
R342 B.n643 B.n642 585
R343 B.n641 B.n112 585
R344 B.n640 B.n639 585
R345 B.n638 B.n113 585
R346 B.n637 B.n636 585
R347 B.n635 B.n114 585
R348 B.n634 B.n633 585
R349 B.n632 B.n115 585
R350 B.n631 B.n630 585
R351 B.n629 B.n116 585
R352 B.n628 B.n627 585
R353 B.n626 B.n117 585
R354 B.n625 B.n624 585
R355 B.n623 B.n118 585
R356 B.n622 B.n621 585
R357 B.n620 B.n119 585
R358 B.n619 B.n618 585
R359 B.n617 B.n120 585
R360 B.n616 B.n615 585
R361 B.n614 B.n121 585
R362 B.n613 B.n612 585
R363 B.n611 B.n122 585
R364 B.n610 B.n609 585
R365 B.n608 B.n123 585
R366 B.n607 B.n606 585
R367 B.n605 B.n124 585
R368 B.n604 B.n603 585
R369 B.n602 B.n125 585
R370 B.n601 B.n600 585
R371 B.n599 B.n126 585
R372 B.n598 B.n597 585
R373 B.n596 B.n127 585
R374 B.n595 B.n594 585
R375 B.n593 B.n128 585
R376 B.n592 B.n591 585
R377 B.n590 B.n129 585
R378 B.n589 B.n588 585
R379 B.n587 B.n130 585
R380 B.n586 B.n585 585
R381 B.n584 B.n131 585
R382 B.n583 B.n582 585
R383 B.n581 B.n132 585
R384 B.n580 B.n579 585
R385 B.n578 B.n133 585
R386 B.n577 B.n576 585
R387 B.n575 B.n134 585
R388 B.n574 B.n573 585
R389 B.n572 B.n135 585
R390 B.n571 B.n570 585
R391 B.n569 B.n136 585
R392 B.n568 B.n567 585
R393 B.n566 B.n137 585
R394 B.n565 B.n564 585
R395 B.n563 B.n138 585
R396 B.n562 B.n561 585
R397 B.n560 B.n139 585
R398 B.n559 B.n558 585
R399 B.n557 B.n140 585
R400 B.n556 B.n555 585
R401 B.n554 B.n141 585
R402 B.n553 B.n552 585
R403 B.n551 B.n142 585
R404 B.n550 B.n549 585
R405 B.n548 B.n143 585
R406 B.n547 B.n546 585
R407 B.n545 B.n144 585
R408 B.n544 B.n543 585
R409 B.n542 B.n145 585
R410 B.n541 B.n540 585
R411 B.n539 B.n146 585
R412 B.n538 B.n537 585
R413 B.n536 B.n147 585
R414 B.n535 B.n534 585
R415 B.n533 B.n148 585
R416 B.n532 B.n531 585
R417 B.n530 B.n149 585
R418 B.n529 B.n528 585
R419 B.n527 B.n150 585
R420 B.n526 B.n525 585
R421 B.n524 B.n151 585
R422 B.n523 B.n522 585
R423 B.n521 B.n152 585
R424 B.n520 B.n519 585
R425 B.n518 B.n153 585
R426 B.n517 B.n516 585
R427 B.n515 B.n154 585
R428 B.n514 B.n513 585
R429 B.n512 B.n155 585
R430 B.n511 B.n510 585
R431 B.n509 B.n156 585
R432 B.n508 B.n507 585
R433 B.n506 B.n157 585
R434 B.n343 B.n342 585
R435 B.n344 B.n215 585
R436 B.n346 B.n345 585
R437 B.n347 B.n214 585
R438 B.n349 B.n348 585
R439 B.n350 B.n213 585
R440 B.n352 B.n351 585
R441 B.n353 B.n212 585
R442 B.n355 B.n354 585
R443 B.n356 B.n211 585
R444 B.n358 B.n357 585
R445 B.n359 B.n210 585
R446 B.n361 B.n360 585
R447 B.n362 B.n209 585
R448 B.n364 B.n363 585
R449 B.n365 B.n208 585
R450 B.n367 B.n366 585
R451 B.n368 B.n207 585
R452 B.n370 B.n369 585
R453 B.n371 B.n206 585
R454 B.n373 B.n372 585
R455 B.n374 B.n205 585
R456 B.n376 B.n375 585
R457 B.n377 B.n204 585
R458 B.n379 B.n378 585
R459 B.n380 B.n203 585
R460 B.n382 B.n381 585
R461 B.n383 B.n202 585
R462 B.n385 B.n384 585
R463 B.n386 B.n201 585
R464 B.n388 B.n387 585
R465 B.n389 B.n200 585
R466 B.n391 B.n390 585
R467 B.n392 B.n199 585
R468 B.n394 B.n393 585
R469 B.n395 B.n198 585
R470 B.n397 B.n396 585
R471 B.n398 B.n197 585
R472 B.n400 B.n399 585
R473 B.n401 B.n196 585
R474 B.n403 B.n402 585
R475 B.n404 B.n195 585
R476 B.n406 B.n405 585
R477 B.n407 B.n194 585
R478 B.n409 B.n408 585
R479 B.n410 B.n193 585
R480 B.n412 B.n411 585
R481 B.n413 B.n192 585
R482 B.n415 B.n414 585
R483 B.n417 B.n416 585
R484 B.n418 B.n188 585
R485 B.n420 B.n419 585
R486 B.n421 B.n187 585
R487 B.n423 B.n422 585
R488 B.n424 B.n186 585
R489 B.n426 B.n425 585
R490 B.n427 B.n185 585
R491 B.n429 B.n428 585
R492 B.n430 B.n182 585
R493 B.n433 B.n432 585
R494 B.n434 B.n181 585
R495 B.n436 B.n435 585
R496 B.n437 B.n180 585
R497 B.n439 B.n438 585
R498 B.n440 B.n179 585
R499 B.n442 B.n441 585
R500 B.n443 B.n178 585
R501 B.n445 B.n444 585
R502 B.n446 B.n177 585
R503 B.n448 B.n447 585
R504 B.n449 B.n176 585
R505 B.n451 B.n450 585
R506 B.n452 B.n175 585
R507 B.n454 B.n453 585
R508 B.n455 B.n174 585
R509 B.n457 B.n456 585
R510 B.n458 B.n173 585
R511 B.n460 B.n459 585
R512 B.n461 B.n172 585
R513 B.n463 B.n462 585
R514 B.n464 B.n171 585
R515 B.n466 B.n465 585
R516 B.n467 B.n170 585
R517 B.n469 B.n468 585
R518 B.n470 B.n169 585
R519 B.n472 B.n471 585
R520 B.n473 B.n168 585
R521 B.n475 B.n474 585
R522 B.n476 B.n167 585
R523 B.n478 B.n477 585
R524 B.n479 B.n166 585
R525 B.n481 B.n480 585
R526 B.n482 B.n165 585
R527 B.n484 B.n483 585
R528 B.n485 B.n164 585
R529 B.n487 B.n486 585
R530 B.n488 B.n163 585
R531 B.n490 B.n489 585
R532 B.n491 B.n162 585
R533 B.n493 B.n492 585
R534 B.n494 B.n161 585
R535 B.n496 B.n495 585
R536 B.n497 B.n160 585
R537 B.n499 B.n498 585
R538 B.n500 B.n159 585
R539 B.n502 B.n501 585
R540 B.n503 B.n158 585
R541 B.n505 B.n504 585
R542 B.n341 B.n216 585
R543 B.n340 B.n339 585
R544 B.n338 B.n217 585
R545 B.n337 B.n336 585
R546 B.n335 B.n218 585
R547 B.n334 B.n333 585
R548 B.n332 B.n219 585
R549 B.n331 B.n330 585
R550 B.n329 B.n220 585
R551 B.n328 B.n327 585
R552 B.n326 B.n221 585
R553 B.n325 B.n324 585
R554 B.n323 B.n222 585
R555 B.n322 B.n321 585
R556 B.n320 B.n223 585
R557 B.n319 B.n318 585
R558 B.n317 B.n224 585
R559 B.n316 B.n315 585
R560 B.n314 B.n225 585
R561 B.n313 B.n312 585
R562 B.n311 B.n226 585
R563 B.n310 B.n309 585
R564 B.n308 B.n227 585
R565 B.n307 B.n306 585
R566 B.n305 B.n228 585
R567 B.n304 B.n303 585
R568 B.n302 B.n229 585
R569 B.n301 B.n300 585
R570 B.n299 B.n230 585
R571 B.n298 B.n297 585
R572 B.n296 B.n231 585
R573 B.n295 B.n294 585
R574 B.n293 B.n232 585
R575 B.n292 B.n291 585
R576 B.n290 B.n233 585
R577 B.n289 B.n288 585
R578 B.n287 B.n234 585
R579 B.n286 B.n285 585
R580 B.n284 B.n235 585
R581 B.n283 B.n282 585
R582 B.n281 B.n236 585
R583 B.n280 B.n279 585
R584 B.n278 B.n237 585
R585 B.n277 B.n276 585
R586 B.n275 B.n238 585
R587 B.n274 B.n273 585
R588 B.n272 B.n239 585
R589 B.n271 B.n270 585
R590 B.n269 B.n240 585
R591 B.n268 B.n267 585
R592 B.n266 B.n241 585
R593 B.n265 B.n264 585
R594 B.n263 B.n242 585
R595 B.n262 B.n261 585
R596 B.n260 B.n243 585
R597 B.n259 B.n258 585
R598 B.n257 B.n244 585
R599 B.n256 B.n255 585
R600 B.n254 B.n245 585
R601 B.n253 B.n252 585
R602 B.n251 B.n246 585
R603 B.n250 B.n249 585
R604 B.n248 B.n247 585
R605 B.n2 B.n0 585
R606 B.n957 B.n1 585
R607 B.n956 B.n955 585
R608 B.n954 B.n3 585
R609 B.n953 B.n952 585
R610 B.n951 B.n4 585
R611 B.n950 B.n949 585
R612 B.n948 B.n5 585
R613 B.n947 B.n946 585
R614 B.n945 B.n6 585
R615 B.n944 B.n943 585
R616 B.n942 B.n7 585
R617 B.n941 B.n940 585
R618 B.n939 B.n8 585
R619 B.n938 B.n937 585
R620 B.n936 B.n9 585
R621 B.n935 B.n934 585
R622 B.n933 B.n10 585
R623 B.n932 B.n931 585
R624 B.n930 B.n11 585
R625 B.n929 B.n928 585
R626 B.n927 B.n12 585
R627 B.n926 B.n925 585
R628 B.n924 B.n13 585
R629 B.n923 B.n922 585
R630 B.n921 B.n14 585
R631 B.n920 B.n919 585
R632 B.n918 B.n15 585
R633 B.n917 B.n916 585
R634 B.n915 B.n16 585
R635 B.n914 B.n913 585
R636 B.n912 B.n17 585
R637 B.n911 B.n910 585
R638 B.n909 B.n18 585
R639 B.n908 B.n907 585
R640 B.n906 B.n19 585
R641 B.n905 B.n904 585
R642 B.n903 B.n20 585
R643 B.n902 B.n901 585
R644 B.n900 B.n21 585
R645 B.n899 B.n898 585
R646 B.n897 B.n22 585
R647 B.n896 B.n895 585
R648 B.n894 B.n23 585
R649 B.n893 B.n892 585
R650 B.n891 B.n24 585
R651 B.n890 B.n889 585
R652 B.n888 B.n25 585
R653 B.n887 B.n886 585
R654 B.n885 B.n26 585
R655 B.n884 B.n883 585
R656 B.n882 B.n27 585
R657 B.n881 B.n880 585
R658 B.n879 B.n28 585
R659 B.n878 B.n877 585
R660 B.n876 B.n29 585
R661 B.n875 B.n874 585
R662 B.n873 B.n30 585
R663 B.n872 B.n871 585
R664 B.n870 B.n31 585
R665 B.n869 B.n868 585
R666 B.n867 B.n32 585
R667 B.n866 B.n865 585
R668 B.n864 B.n33 585
R669 B.n863 B.n862 585
R670 B.n959 B.n958 585
R671 B.n343 B.n216 554.963
R672 B.n862 B.n861 554.963
R673 B.n506 B.n505 554.963
R674 B.n699 B.n698 554.963
R675 B.n183 B.t9 332.024
R676 B.n189 B.t6 332.024
R677 B.n60 B.t0 332.024
R678 B.n67 B.t3 332.024
R679 B.n183 B.t11 174.883
R680 B.n67 B.t4 174.883
R681 B.n189 B.t8 174.865
R682 B.n60 B.t1 174.865
R683 B.n339 B.n216 163.367
R684 B.n339 B.n338 163.367
R685 B.n338 B.n337 163.367
R686 B.n337 B.n218 163.367
R687 B.n333 B.n218 163.367
R688 B.n333 B.n332 163.367
R689 B.n332 B.n331 163.367
R690 B.n331 B.n220 163.367
R691 B.n327 B.n220 163.367
R692 B.n327 B.n326 163.367
R693 B.n326 B.n325 163.367
R694 B.n325 B.n222 163.367
R695 B.n321 B.n222 163.367
R696 B.n321 B.n320 163.367
R697 B.n320 B.n319 163.367
R698 B.n319 B.n224 163.367
R699 B.n315 B.n224 163.367
R700 B.n315 B.n314 163.367
R701 B.n314 B.n313 163.367
R702 B.n313 B.n226 163.367
R703 B.n309 B.n226 163.367
R704 B.n309 B.n308 163.367
R705 B.n308 B.n307 163.367
R706 B.n307 B.n228 163.367
R707 B.n303 B.n228 163.367
R708 B.n303 B.n302 163.367
R709 B.n302 B.n301 163.367
R710 B.n301 B.n230 163.367
R711 B.n297 B.n230 163.367
R712 B.n297 B.n296 163.367
R713 B.n296 B.n295 163.367
R714 B.n295 B.n232 163.367
R715 B.n291 B.n232 163.367
R716 B.n291 B.n290 163.367
R717 B.n290 B.n289 163.367
R718 B.n289 B.n234 163.367
R719 B.n285 B.n234 163.367
R720 B.n285 B.n284 163.367
R721 B.n284 B.n283 163.367
R722 B.n283 B.n236 163.367
R723 B.n279 B.n236 163.367
R724 B.n279 B.n278 163.367
R725 B.n278 B.n277 163.367
R726 B.n277 B.n238 163.367
R727 B.n273 B.n238 163.367
R728 B.n273 B.n272 163.367
R729 B.n272 B.n271 163.367
R730 B.n271 B.n240 163.367
R731 B.n267 B.n240 163.367
R732 B.n267 B.n266 163.367
R733 B.n266 B.n265 163.367
R734 B.n265 B.n242 163.367
R735 B.n261 B.n242 163.367
R736 B.n261 B.n260 163.367
R737 B.n260 B.n259 163.367
R738 B.n259 B.n244 163.367
R739 B.n255 B.n244 163.367
R740 B.n255 B.n254 163.367
R741 B.n254 B.n253 163.367
R742 B.n253 B.n246 163.367
R743 B.n249 B.n246 163.367
R744 B.n249 B.n248 163.367
R745 B.n248 B.n2 163.367
R746 B.n958 B.n2 163.367
R747 B.n958 B.n957 163.367
R748 B.n957 B.n956 163.367
R749 B.n956 B.n3 163.367
R750 B.n952 B.n3 163.367
R751 B.n952 B.n951 163.367
R752 B.n951 B.n950 163.367
R753 B.n950 B.n5 163.367
R754 B.n946 B.n5 163.367
R755 B.n946 B.n945 163.367
R756 B.n945 B.n944 163.367
R757 B.n944 B.n7 163.367
R758 B.n940 B.n7 163.367
R759 B.n940 B.n939 163.367
R760 B.n939 B.n938 163.367
R761 B.n938 B.n9 163.367
R762 B.n934 B.n9 163.367
R763 B.n934 B.n933 163.367
R764 B.n933 B.n932 163.367
R765 B.n932 B.n11 163.367
R766 B.n928 B.n11 163.367
R767 B.n928 B.n927 163.367
R768 B.n927 B.n926 163.367
R769 B.n926 B.n13 163.367
R770 B.n922 B.n13 163.367
R771 B.n922 B.n921 163.367
R772 B.n921 B.n920 163.367
R773 B.n920 B.n15 163.367
R774 B.n916 B.n15 163.367
R775 B.n916 B.n915 163.367
R776 B.n915 B.n914 163.367
R777 B.n914 B.n17 163.367
R778 B.n910 B.n17 163.367
R779 B.n910 B.n909 163.367
R780 B.n909 B.n908 163.367
R781 B.n908 B.n19 163.367
R782 B.n904 B.n19 163.367
R783 B.n904 B.n903 163.367
R784 B.n903 B.n902 163.367
R785 B.n902 B.n21 163.367
R786 B.n898 B.n21 163.367
R787 B.n898 B.n897 163.367
R788 B.n897 B.n896 163.367
R789 B.n896 B.n23 163.367
R790 B.n892 B.n23 163.367
R791 B.n892 B.n891 163.367
R792 B.n891 B.n890 163.367
R793 B.n890 B.n25 163.367
R794 B.n886 B.n25 163.367
R795 B.n886 B.n885 163.367
R796 B.n885 B.n884 163.367
R797 B.n884 B.n27 163.367
R798 B.n880 B.n27 163.367
R799 B.n880 B.n879 163.367
R800 B.n879 B.n878 163.367
R801 B.n878 B.n29 163.367
R802 B.n874 B.n29 163.367
R803 B.n874 B.n873 163.367
R804 B.n873 B.n872 163.367
R805 B.n872 B.n31 163.367
R806 B.n868 B.n31 163.367
R807 B.n868 B.n867 163.367
R808 B.n867 B.n866 163.367
R809 B.n866 B.n33 163.367
R810 B.n862 B.n33 163.367
R811 B.n344 B.n343 163.367
R812 B.n345 B.n344 163.367
R813 B.n345 B.n214 163.367
R814 B.n349 B.n214 163.367
R815 B.n350 B.n349 163.367
R816 B.n351 B.n350 163.367
R817 B.n351 B.n212 163.367
R818 B.n355 B.n212 163.367
R819 B.n356 B.n355 163.367
R820 B.n357 B.n356 163.367
R821 B.n357 B.n210 163.367
R822 B.n361 B.n210 163.367
R823 B.n362 B.n361 163.367
R824 B.n363 B.n362 163.367
R825 B.n363 B.n208 163.367
R826 B.n367 B.n208 163.367
R827 B.n368 B.n367 163.367
R828 B.n369 B.n368 163.367
R829 B.n369 B.n206 163.367
R830 B.n373 B.n206 163.367
R831 B.n374 B.n373 163.367
R832 B.n375 B.n374 163.367
R833 B.n375 B.n204 163.367
R834 B.n379 B.n204 163.367
R835 B.n380 B.n379 163.367
R836 B.n381 B.n380 163.367
R837 B.n381 B.n202 163.367
R838 B.n385 B.n202 163.367
R839 B.n386 B.n385 163.367
R840 B.n387 B.n386 163.367
R841 B.n387 B.n200 163.367
R842 B.n391 B.n200 163.367
R843 B.n392 B.n391 163.367
R844 B.n393 B.n392 163.367
R845 B.n393 B.n198 163.367
R846 B.n397 B.n198 163.367
R847 B.n398 B.n397 163.367
R848 B.n399 B.n398 163.367
R849 B.n399 B.n196 163.367
R850 B.n403 B.n196 163.367
R851 B.n404 B.n403 163.367
R852 B.n405 B.n404 163.367
R853 B.n405 B.n194 163.367
R854 B.n409 B.n194 163.367
R855 B.n410 B.n409 163.367
R856 B.n411 B.n410 163.367
R857 B.n411 B.n192 163.367
R858 B.n415 B.n192 163.367
R859 B.n416 B.n415 163.367
R860 B.n416 B.n188 163.367
R861 B.n420 B.n188 163.367
R862 B.n421 B.n420 163.367
R863 B.n422 B.n421 163.367
R864 B.n422 B.n186 163.367
R865 B.n426 B.n186 163.367
R866 B.n427 B.n426 163.367
R867 B.n428 B.n427 163.367
R868 B.n428 B.n182 163.367
R869 B.n433 B.n182 163.367
R870 B.n434 B.n433 163.367
R871 B.n435 B.n434 163.367
R872 B.n435 B.n180 163.367
R873 B.n439 B.n180 163.367
R874 B.n440 B.n439 163.367
R875 B.n441 B.n440 163.367
R876 B.n441 B.n178 163.367
R877 B.n445 B.n178 163.367
R878 B.n446 B.n445 163.367
R879 B.n447 B.n446 163.367
R880 B.n447 B.n176 163.367
R881 B.n451 B.n176 163.367
R882 B.n452 B.n451 163.367
R883 B.n453 B.n452 163.367
R884 B.n453 B.n174 163.367
R885 B.n457 B.n174 163.367
R886 B.n458 B.n457 163.367
R887 B.n459 B.n458 163.367
R888 B.n459 B.n172 163.367
R889 B.n463 B.n172 163.367
R890 B.n464 B.n463 163.367
R891 B.n465 B.n464 163.367
R892 B.n465 B.n170 163.367
R893 B.n469 B.n170 163.367
R894 B.n470 B.n469 163.367
R895 B.n471 B.n470 163.367
R896 B.n471 B.n168 163.367
R897 B.n475 B.n168 163.367
R898 B.n476 B.n475 163.367
R899 B.n477 B.n476 163.367
R900 B.n477 B.n166 163.367
R901 B.n481 B.n166 163.367
R902 B.n482 B.n481 163.367
R903 B.n483 B.n482 163.367
R904 B.n483 B.n164 163.367
R905 B.n487 B.n164 163.367
R906 B.n488 B.n487 163.367
R907 B.n489 B.n488 163.367
R908 B.n489 B.n162 163.367
R909 B.n493 B.n162 163.367
R910 B.n494 B.n493 163.367
R911 B.n495 B.n494 163.367
R912 B.n495 B.n160 163.367
R913 B.n499 B.n160 163.367
R914 B.n500 B.n499 163.367
R915 B.n501 B.n500 163.367
R916 B.n501 B.n158 163.367
R917 B.n505 B.n158 163.367
R918 B.n507 B.n506 163.367
R919 B.n507 B.n156 163.367
R920 B.n511 B.n156 163.367
R921 B.n512 B.n511 163.367
R922 B.n513 B.n512 163.367
R923 B.n513 B.n154 163.367
R924 B.n517 B.n154 163.367
R925 B.n518 B.n517 163.367
R926 B.n519 B.n518 163.367
R927 B.n519 B.n152 163.367
R928 B.n523 B.n152 163.367
R929 B.n524 B.n523 163.367
R930 B.n525 B.n524 163.367
R931 B.n525 B.n150 163.367
R932 B.n529 B.n150 163.367
R933 B.n530 B.n529 163.367
R934 B.n531 B.n530 163.367
R935 B.n531 B.n148 163.367
R936 B.n535 B.n148 163.367
R937 B.n536 B.n535 163.367
R938 B.n537 B.n536 163.367
R939 B.n537 B.n146 163.367
R940 B.n541 B.n146 163.367
R941 B.n542 B.n541 163.367
R942 B.n543 B.n542 163.367
R943 B.n543 B.n144 163.367
R944 B.n547 B.n144 163.367
R945 B.n548 B.n547 163.367
R946 B.n549 B.n548 163.367
R947 B.n549 B.n142 163.367
R948 B.n553 B.n142 163.367
R949 B.n554 B.n553 163.367
R950 B.n555 B.n554 163.367
R951 B.n555 B.n140 163.367
R952 B.n559 B.n140 163.367
R953 B.n560 B.n559 163.367
R954 B.n561 B.n560 163.367
R955 B.n561 B.n138 163.367
R956 B.n565 B.n138 163.367
R957 B.n566 B.n565 163.367
R958 B.n567 B.n566 163.367
R959 B.n567 B.n136 163.367
R960 B.n571 B.n136 163.367
R961 B.n572 B.n571 163.367
R962 B.n573 B.n572 163.367
R963 B.n573 B.n134 163.367
R964 B.n577 B.n134 163.367
R965 B.n578 B.n577 163.367
R966 B.n579 B.n578 163.367
R967 B.n579 B.n132 163.367
R968 B.n583 B.n132 163.367
R969 B.n584 B.n583 163.367
R970 B.n585 B.n584 163.367
R971 B.n585 B.n130 163.367
R972 B.n589 B.n130 163.367
R973 B.n590 B.n589 163.367
R974 B.n591 B.n590 163.367
R975 B.n591 B.n128 163.367
R976 B.n595 B.n128 163.367
R977 B.n596 B.n595 163.367
R978 B.n597 B.n596 163.367
R979 B.n597 B.n126 163.367
R980 B.n601 B.n126 163.367
R981 B.n602 B.n601 163.367
R982 B.n603 B.n602 163.367
R983 B.n603 B.n124 163.367
R984 B.n607 B.n124 163.367
R985 B.n608 B.n607 163.367
R986 B.n609 B.n608 163.367
R987 B.n609 B.n122 163.367
R988 B.n613 B.n122 163.367
R989 B.n614 B.n613 163.367
R990 B.n615 B.n614 163.367
R991 B.n615 B.n120 163.367
R992 B.n619 B.n120 163.367
R993 B.n620 B.n619 163.367
R994 B.n621 B.n620 163.367
R995 B.n621 B.n118 163.367
R996 B.n625 B.n118 163.367
R997 B.n626 B.n625 163.367
R998 B.n627 B.n626 163.367
R999 B.n627 B.n116 163.367
R1000 B.n631 B.n116 163.367
R1001 B.n632 B.n631 163.367
R1002 B.n633 B.n632 163.367
R1003 B.n633 B.n114 163.367
R1004 B.n637 B.n114 163.367
R1005 B.n638 B.n637 163.367
R1006 B.n639 B.n638 163.367
R1007 B.n639 B.n112 163.367
R1008 B.n643 B.n112 163.367
R1009 B.n644 B.n643 163.367
R1010 B.n645 B.n644 163.367
R1011 B.n645 B.n110 163.367
R1012 B.n649 B.n110 163.367
R1013 B.n650 B.n649 163.367
R1014 B.n651 B.n650 163.367
R1015 B.n651 B.n108 163.367
R1016 B.n655 B.n108 163.367
R1017 B.n656 B.n655 163.367
R1018 B.n657 B.n656 163.367
R1019 B.n657 B.n106 163.367
R1020 B.n661 B.n106 163.367
R1021 B.n662 B.n661 163.367
R1022 B.n663 B.n662 163.367
R1023 B.n663 B.n104 163.367
R1024 B.n667 B.n104 163.367
R1025 B.n668 B.n667 163.367
R1026 B.n669 B.n668 163.367
R1027 B.n669 B.n102 163.367
R1028 B.n673 B.n102 163.367
R1029 B.n674 B.n673 163.367
R1030 B.n675 B.n674 163.367
R1031 B.n675 B.n100 163.367
R1032 B.n679 B.n100 163.367
R1033 B.n680 B.n679 163.367
R1034 B.n681 B.n680 163.367
R1035 B.n681 B.n98 163.367
R1036 B.n685 B.n98 163.367
R1037 B.n686 B.n685 163.367
R1038 B.n687 B.n686 163.367
R1039 B.n687 B.n96 163.367
R1040 B.n691 B.n96 163.367
R1041 B.n692 B.n691 163.367
R1042 B.n693 B.n692 163.367
R1043 B.n693 B.n94 163.367
R1044 B.n697 B.n94 163.367
R1045 B.n698 B.n697 163.367
R1046 B.n861 B.n860 163.367
R1047 B.n860 B.n35 163.367
R1048 B.n856 B.n35 163.367
R1049 B.n856 B.n855 163.367
R1050 B.n855 B.n854 163.367
R1051 B.n854 B.n37 163.367
R1052 B.n850 B.n37 163.367
R1053 B.n850 B.n849 163.367
R1054 B.n849 B.n848 163.367
R1055 B.n848 B.n39 163.367
R1056 B.n844 B.n39 163.367
R1057 B.n844 B.n843 163.367
R1058 B.n843 B.n842 163.367
R1059 B.n842 B.n41 163.367
R1060 B.n838 B.n41 163.367
R1061 B.n838 B.n837 163.367
R1062 B.n837 B.n836 163.367
R1063 B.n836 B.n43 163.367
R1064 B.n832 B.n43 163.367
R1065 B.n832 B.n831 163.367
R1066 B.n831 B.n830 163.367
R1067 B.n830 B.n45 163.367
R1068 B.n826 B.n45 163.367
R1069 B.n826 B.n825 163.367
R1070 B.n825 B.n824 163.367
R1071 B.n824 B.n47 163.367
R1072 B.n820 B.n47 163.367
R1073 B.n820 B.n819 163.367
R1074 B.n819 B.n818 163.367
R1075 B.n818 B.n49 163.367
R1076 B.n814 B.n49 163.367
R1077 B.n814 B.n813 163.367
R1078 B.n813 B.n812 163.367
R1079 B.n812 B.n51 163.367
R1080 B.n808 B.n51 163.367
R1081 B.n808 B.n807 163.367
R1082 B.n807 B.n806 163.367
R1083 B.n806 B.n53 163.367
R1084 B.n802 B.n53 163.367
R1085 B.n802 B.n801 163.367
R1086 B.n801 B.n800 163.367
R1087 B.n800 B.n55 163.367
R1088 B.n796 B.n55 163.367
R1089 B.n796 B.n795 163.367
R1090 B.n795 B.n794 163.367
R1091 B.n794 B.n57 163.367
R1092 B.n790 B.n57 163.367
R1093 B.n790 B.n789 163.367
R1094 B.n789 B.n788 163.367
R1095 B.n788 B.n59 163.367
R1096 B.n784 B.n59 163.367
R1097 B.n784 B.n783 163.367
R1098 B.n783 B.n782 163.367
R1099 B.n782 B.n64 163.367
R1100 B.n778 B.n64 163.367
R1101 B.n778 B.n777 163.367
R1102 B.n777 B.n776 163.367
R1103 B.n776 B.n66 163.367
R1104 B.n771 B.n66 163.367
R1105 B.n771 B.n770 163.367
R1106 B.n770 B.n769 163.367
R1107 B.n769 B.n70 163.367
R1108 B.n765 B.n70 163.367
R1109 B.n765 B.n764 163.367
R1110 B.n764 B.n763 163.367
R1111 B.n763 B.n72 163.367
R1112 B.n759 B.n72 163.367
R1113 B.n759 B.n758 163.367
R1114 B.n758 B.n757 163.367
R1115 B.n757 B.n74 163.367
R1116 B.n753 B.n74 163.367
R1117 B.n753 B.n752 163.367
R1118 B.n752 B.n751 163.367
R1119 B.n751 B.n76 163.367
R1120 B.n747 B.n76 163.367
R1121 B.n747 B.n746 163.367
R1122 B.n746 B.n745 163.367
R1123 B.n745 B.n78 163.367
R1124 B.n741 B.n78 163.367
R1125 B.n741 B.n740 163.367
R1126 B.n740 B.n739 163.367
R1127 B.n739 B.n80 163.367
R1128 B.n735 B.n80 163.367
R1129 B.n735 B.n734 163.367
R1130 B.n734 B.n733 163.367
R1131 B.n733 B.n82 163.367
R1132 B.n729 B.n82 163.367
R1133 B.n729 B.n728 163.367
R1134 B.n728 B.n727 163.367
R1135 B.n727 B.n84 163.367
R1136 B.n723 B.n84 163.367
R1137 B.n723 B.n722 163.367
R1138 B.n722 B.n721 163.367
R1139 B.n721 B.n86 163.367
R1140 B.n717 B.n86 163.367
R1141 B.n717 B.n716 163.367
R1142 B.n716 B.n715 163.367
R1143 B.n715 B.n88 163.367
R1144 B.n711 B.n88 163.367
R1145 B.n711 B.n710 163.367
R1146 B.n710 B.n709 163.367
R1147 B.n709 B.n90 163.367
R1148 B.n705 B.n90 163.367
R1149 B.n705 B.n704 163.367
R1150 B.n704 B.n703 163.367
R1151 B.n703 B.n92 163.367
R1152 B.n699 B.n92 163.367
R1153 B.n184 B.t10 113.21
R1154 B.n68 B.t5 113.21
R1155 B.n190 B.t7 113.192
R1156 B.n61 B.t2 113.192
R1157 B.n184 B.n183 61.6732
R1158 B.n190 B.n189 61.6732
R1159 B.n61 B.n60 61.6732
R1160 B.n68 B.n67 61.6732
R1161 B.n431 B.n184 59.5399
R1162 B.n191 B.n190 59.5399
R1163 B.n62 B.n61 59.5399
R1164 B.n773 B.n68 59.5399
R1165 B.n700 B.n93 36.059
R1166 B.n863 B.n34 36.059
R1167 B.n504 B.n157 36.059
R1168 B.n342 B.n341 36.059
R1169 B B.n959 18.0485
R1170 B.n859 B.n34 10.6151
R1171 B.n859 B.n858 10.6151
R1172 B.n858 B.n857 10.6151
R1173 B.n857 B.n36 10.6151
R1174 B.n853 B.n36 10.6151
R1175 B.n853 B.n852 10.6151
R1176 B.n852 B.n851 10.6151
R1177 B.n851 B.n38 10.6151
R1178 B.n847 B.n38 10.6151
R1179 B.n847 B.n846 10.6151
R1180 B.n846 B.n845 10.6151
R1181 B.n845 B.n40 10.6151
R1182 B.n841 B.n40 10.6151
R1183 B.n841 B.n840 10.6151
R1184 B.n840 B.n839 10.6151
R1185 B.n839 B.n42 10.6151
R1186 B.n835 B.n42 10.6151
R1187 B.n835 B.n834 10.6151
R1188 B.n834 B.n833 10.6151
R1189 B.n833 B.n44 10.6151
R1190 B.n829 B.n44 10.6151
R1191 B.n829 B.n828 10.6151
R1192 B.n828 B.n827 10.6151
R1193 B.n827 B.n46 10.6151
R1194 B.n823 B.n46 10.6151
R1195 B.n823 B.n822 10.6151
R1196 B.n822 B.n821 10.6151
R1197 B.n821 B.n48 10.6151
R1198 B.n817 B.n48 10.6151
R1199 B.n817 B.n816 10.6151
R1200 B.n816 B.n815 10.6151
R1201 B.n815 B.n50 10.6151
R1202 B.n811 B.n50 10.6151
R1203 B.n811 B.n810 10.6151
R1204 B.n810 B.n809 10.6151
R1205 B.n809 B.n52 10.6151
R1206 B.n805 B.n52 10.6151
R1207 B.n805 B.n804 10.6151
R1208 B.n804 B.n803 10.6151
R1209 B.n803 B.n54 10.6151
R1210 B.n799 B.n54 10.6151
R1211 B.n799 B.n798 10.6151
R1212 B.n798 B.n797 10.6151
R1213 B.n797 B.n56 10.6151
R1214 B.n793 B.n56 10.6151
R1215 B.n793 B.n792 10.6151
R1216 B.n792 B.n791 10.6151
R1217 B.n791 B.n58 10.6151
R1218 B.n787 B.n786 10.6151
R1219 B.n786 B.n785 10.6151
R1220 B.n785 B.n63 10.6151
R1221 B.n781 B.n63 10.6151
R1222 B.n781 B.n780 10.6151
R1223 B.n780 B.n779 10.6151
R1224 B.n779 B.n65 10.6151
R1225 B.n775 B.n65 10.6151
R1226 B.n775 B.n774 10.6151
R1227 B.n772 B.n69 10.6151
R1228 B.n768 B.n69 10.6151
R1229 B.n768 B.n767 10.6151
R1230 B.n767 B.n766 10.6151
R1231 B.n766 B.n71 10.6151
R1232 B.n762 B.n71 10.6151
R1233 B.n762 B.n761 10.6151
R1234 B.n761 B.n760 10.6151
R1235 B.n760 B.n73 10.6151
R1236 B.n756 B.n73 10.6151
R1237 B.n756 B.n755 10.6151
R1238 B.n755 B.n754 10.6151
R1239 B.n754 B.n75 10.6151
R1240 B.n750 B.n75 10.6151
R1241 B.n750 B.n749 10.6151
R1242 B.n749 B.n748 10.6151
R1243 B.n748 B.n77 10.6151
R1244 B.n744 B.n77 10.6151
R1245 B.n744 B.n743 10.6151
R1246 B.n743 B.n742 10.6151
R1247 B.n742 B.n79 10.6151
R1248 B.n738 B.n79 10.6151
R1249 B.n738 B.n737 10.6151
R1250 B.n737 B.n736 10.6151
R1251 B.n736 B.n81 10.6151
R1252 B.n732 B.n81 10.6151
R1253 B.n732 B.n731 10.6151
R1254 B.n731 B.n730 10.6151
R1255 B.n730 B.n83 10.6151
R1256 B.n726 B.n83 10.6151
R1257 B.n726 B.n725 10.6151
R1258 B.n725 B.n724 10.6151
R1259 B.n724 B.n85 10.6151
R1260 B.n720 B.n85 10.6151
R1261 B.n720 B.n719 10.6151
R1262 B.n719 B.n718 10.6151
R1263 B.n718 B.n87 10.6151
R1264 B.n714 B.n87 10.6151
R1265 B.n714 B.n713 10.6151
R1266 B.n713 B.n712 10.6151
R1267 B.n712 B.n89 10.6151
R1268 B.n708 B.n89 10.6151
R1269 B.n708 B.n707 10.6151
R1270 B.n707 B.n706 10.6151
R1271 B.n706 B.n91 10.6151
R1272 B.n702 B.n91 10.6151
R1273 B.n702 B.n701 10.6151
R1274 B.n701 B.n700 10.6151
R1275 B.n508 B.n157 10.6151
R1276 B.n509 B.n508 10.6151
R1277 B.n510 B.n509 10.6151
R1278 B.n510 B.n155 10.6151
R1279 B.n514 B.n155 10.6151
R1280 B.n515 B.n514 10.6151
R1281 B.n516 B.n515 10.6151
R1282 B.n516 B.n153 10.6151
R1283 B.n520 B.n153 10.6151
R1284 B.n521 B.n520 10.6151
R1285 B.n522 B.n521 10.6151
R1286 B.n522 B.n151 10.6151
R1287 B.n526 B.n151 10.6151
R1288 B.n527 B.n526 10.6151
R1289 B.n528 B.n527 10.6151
R1290 B.n528 B.n149 10.6151
R1291 B.n532 B.n149 10.6151
R1292 B.n533 B.n532 10.6151
R1293 B.n534 B.n533 10.6151
R1294 B.n534 B.n147 10.6151
R1295 B.n538 B.n147 10.6151
R1296 B.n539 B.n538 10.6151
R1297 B.n540 B.n539 10.6151
R1298 B.n540 B.n145 10.6151
R1299 B.n544 B.n145 10.6151
R1300 B.n545 B.n544 10.6151
R1301 B.n546 B.n545 10.6151
R1302 B.n546 B.n143 10.6151
R1303 B.n550 B.n143 10.6151
R1304 B.n551 B.n550 10.6151
R1305 B.n552 B.n551 10.6151
R1306 B.n552 B.n141 10.6151
R1307 B.n556 B.n141 10.6151
R1308 B.n557 B.n556 10.6151
R1309 B.n558 B.n557 10.6151
R1310 B.n558 B.n139 10.6151
R1311 B.n562 B.n139 10.6151
R1312 B.n563 B.n562 10.6151
R1313 B.n564 B.n563 10.6151
R1314 B.n564 B.n137 10.6151
R1315 B.n568 B.n137 10.6151
R1316 B.n569 B.n568 10.6151
R1317 B.n570 B.n569 10.6151
R1318 B.n570 B.n135 10.6151
R1319 B.n574 B.n135 10.6151
R1320 B.n575 B.n574 10.6151
R1321 B.n576 B.n575 10.6151
R1322 B.n576 B.n133 10.6151
R1323 B.n580 B.n133 10.6151
R1324 B.n581 B.n580 10.6151
R1325 B.n582 B.n581 10.6151
R1326 B.n582 B.n131 10.6151
R1327 B.n586 B.n131 10.6151
R1328 B.n587 B.n586 10.6151
R1329 B.n588 B.n587 10.6151
R1330 B.n588 B.n129 10.6151
R1331 B.n592 B.n129 10.6151
R1332 B.n593 B.n592 10.6151
R1333 B.n594 B.n593 10.6151
R1334 B.n594 B.n127 10.6151
R1335 B.n598 B.n127 10.6151
R1336 B.n599 B.n598 10.6151
R1337 B.n600 B.n599 10.6151
R1338 B.n600 B.n125 10.6151
R1339 B.n604 B.n125 10.6151
R1340 B.n605 B.n604 10.6151
R1341 B.n606 B.n605 10.6151
R1342 B.n606 B.n123 10.6151
R1343 B.n610 B.n123 10.6151
R1344 B.n611 B.n610 10.6151
R1345 B.n612 B.n611 10.6151
R1346 B.n612 B.n121 10.6151
R1347 B.n616 B.n121 10.6151
R1348 B.n617 B.n616 10.6151
R1349 B.n618 B.n617 10.6151
R1350 B.n618 B.n119 10.6151
R1351 B.n622 B.n119 10.6151
R1352 B.n623 B.n622 10.6151
R1353 B.n624 B.n623 10.6151
R1354 B.n624 B.n117 10.6151
R1355 B.n628 B.n117 10.6151
R1356 B.n629 B.n628 10.6151
R1357 B.n630 B.n629 10.6151
R1358 B.n630 B.n115 10.6151
R1359 B.n634 B.n115 10.6151
R1360 B.n635 B.n634 10.6151
R1361 B.n636 B.n635 10.6151
R1362 B.n636 B.n113 10.6151
R1363 B.n640 B.n113 10.6151
R1364 B.n641 B.n640 10.6151
R1365 B.n642 B.n641 10.6151
R1366 B.n642 B.n111 10.6151
R1367 B.n646 B.n111 10.6151
R1368 B.n647 B.n646 10.6151
R1369 B.n648 B.n647 10.6151
R1370 B.n648 B.n109 10.6151
R1371 B.n652 B.n109 10.6151
R1372 B.n653 B.n652 10.6151
R1373 B.n654 B.n653 10.6151
R1374 B.n654 B.n107 10.6151
R1375 B.n658 B.n107 10.6151
R1376 B.n659 B.n658 10.6151
R1377 B.n660 B.n659 10.6151
R1378 B.n660 B.n105 10.6151
R1379 B.n664 B.n105 10.6151
R1380 B.n665 B.n664 10.6151
R1381 B.n666 B.n665 10.6151
R1382 B.n666 B.n103 10.6151
R1383 B.n670 B.n103 10.6151
R1384 B.n671 B.n670 10.6151
R1385 B.n672 B.n671 10.6151
R1386 B.n672 B.n101 10.6151
R1387 B.n676 B.n101 10.6151
R1388 B.n677 B.n676 10.6151
R1389 B.n678 B.n677 10.6151
R1390 B.n678 B.n99 10.6151
R1391 B.n682 B.n99 10.6151
R1392 B.n683 B.n682 10.6151
R1393 B.n684 B.n683 10.6151
R1394 B.n684 B.n97 10.6151
R1395 B.n688 B.n97 10.6151
R1396 B.n689 B.n688 10.6151
R1397 B.n690 B.n689 10.6151
R1398 B.n690 B.n95 10.6151
R1399 B.n694 B.n95 10.6151
R1400 B.n695 B.n694 10.6151
R1401 B.n696 B.n695 10.6151
R1402 B.n696 B.n93 10.6151
R1403 B.n342 B.n215 10.6151
R1404 B.n346 B.n215 10.6151
R1405 B.n347 B.n346 10.6151
R1406 B.n348 B.n347 10.6151
R1407 B.n348 B.n213 10.6151
R1408 B.n352 B.n213 10.6151
R1409 B.n353 B.n352 10.6151
R1410 B.n354 B.n353 10.6151
R1411 B.n354 B.n211 10.6151
R1412 B.n358 B.n211 10.6151
R1413 B.n359 B.n358 10.6151
R1414 B.n360 B.n359 10.6151
R1415 B.n360 B.n209 10.6151
R1416 B.n364 B.n209 10.6151
R1417 B.n365 B.n364 10.6151
R1418 B.n366 B.n365 10.6151
R1419 B.n366 B.n207 10.6151
R1420 B.n370 B.n207 10.6151
R1421 B.n371 B.n370 10.6151
R1422 B.n372 B.n371 10.6151
R1423 B.n372 B.n205 10.6151
R1424 B.n376 B.n205 10.6151
R1425 B.n377 B.n376 10.6151
R1426 B.n378 B.n377 10.6151
R1427 B.n378 B.n203 10.6151
R1428 B.n382 B.n203 10.6151
R1429 B.n383 B.n382 10.6151
R1430 B.n384 B.n383 10.6151
R1431 B.n384 B.n201 10.6151
R1432 B.n388 B.n201 10.6151
R1433 B.n389 B.n388 10.6151
R1434 B.n390 B.n389 10.6151
R1435 B.n390 B.n199 10.6151
R1436 B.n394 B.n199 10.6151
R1437 B.n395 B.n394 10.6151
R1438 B.n396 B.n395 10.6151
R1439 B.n396 B.n197 10.6151
R1440 B.n400 B.n197 10.6151
R1441 B.n401 B.n400 10.6151
R1442 B.n402 B.n401 10.6151
R1443 B.n402 B.n195 10.6151
R1444 B.n406 B.n195 10.6151
R1445 B.n407 B.n406 10.6151
R1446 B.n408 B.n407 10.6151
R1447 B.n408 B.n193 10.6151
R1448 B.n412 B.n193 10.6151
R1449 B.n413 B.n412 10.6151
R1450 B.n414 B.n413 10.6151
R1451 B.n418 B.n417 10.6151
R1452 B.n419 B.n418 10.6151
R1453 B.n419 B.n187 10.6151
R1454 B.n423 B.n187 10.6151
R1455 B.n424 B.n423 10.6151
R1456 B.n425 B.n424 10.6151
R1457 B.n425 B.n185 10.6151
R1458 B.n429 B.n185 10.6151
R1459 B.n430 B.n429 10.6151
R1460 B.n432 B.n181 10.6151
R1461 B.n436 B.n181 10.6151
R1462 B.n437 B.n436 10.6151
R1463 B.n438 B.n437 10.6151
R1464 B.n438 B.n179 10.6151
R1465 B.n442 B.n179 10.6151
R1466 B.n443 B.n442 10.6151
R1467 B.n444 B.n443 10.6151
R1468 B.n444 B.n177 10.6151
R1469 B.n448 B.n177 10.6151
R1470 B.n449 B.n448 10.6151
R1471 B.n450 B.n449 10.6151
R1472 B.n450 B.n175 10.6151
R1473 B.n454 B.n175 10.6151
R1474 B.n455 B.n454 10.6151
R1475 B.n456 B.n455 10.6151
R1476 B.n456 B.n173 10.6151
R1477 B.n460 B.n173 10.6151
R1478 B.n461 B.n460 10.6151
R1479 B.n462 B.n461 10.6151
R1480 B.n462 B.n171 10.6151
R1481 B.n466 B.n171 10.6151
R1482 B.n467 B.n466 10.6151
R1483 B.n468 B.n467 10.6151
R1484 B.n468 B.n169 10.6151
R1485 B.n472 B.n169 10.6151
R1486 B.n473 B.n472 10.6151
R1487 B.n474 B.n473 10.6151
R1488 B.n474 B.n167 10.6151
R1489 B.n478 B.n167 10.6151
R1490 B.n479 B.n478 10.6151
R1491 B.n480 B.n479 10.6151
R1492 B.n480 B.n165 10.6151
R1493 B.n484 B.n165 10.6151
R1494 B.n485 B.n484 10.6151
R1495 B.n486 B.n485 10.6151
R1496 B.n486 B.n163 10.6151
R1497 B.n490 B.n163 10.6151
R1498 B.n491 B.n490 10.6151
R1499 B.n492 B.n491 10.6151
R1500 B.n492 B.n161 10.6151
R1501 B.n496 B.n161 10.6151
R1502 B.n497 B.n496 10.6151
R1503 B.n498 B.n497 10.6151
R1504 B.n498 B.n159 10.6151
R1505 B.n502 B.n159 10.6151
R1506 B.n503 B.n502 10.6151
R1507 B.n504 B.n503 10.6151
R1508 B.n341 B.n340 10.6151
R1509 B.n340 B.n217 10.6151
R1510 B.n336 B.n217 10.6151
R1511 B.n336 B.n335 10.6151
R1512 B.n335 B.n334 10.6151
R1513 B.n334 B.n219 10.6151
R1514 B.n330 B.n219 10.6151
R1515 B.n330 B.n329 10.6151
R1516 B.n329 B.n328 10.6151
R1517 B.n328 B.n221 10.6151
R1518 B.n324 B.n221 10.6151
R1519 B.n324 B.n323 10.6151
R1520 B.n323 B.n322 10.6151
R1521 B.n322 B.n223 10.6151
R1522 B.n318 B.n223 10.6151
R1523 B.n318 B.n317 10.6151
R1524 B.n317 B.n316 10.6151
R1525 B.n316 B.n225 10.6151
R1526 B.n312 B.n225 10.6151
R1527 B.n312 B.n311 10.6151
R1528 B.n311 B.n310 10.6151
R1529 B.n310 B.n227 10.6151
R1530 B.n306 B.n227 10.6151
R1531 B.n306 B.n305 10.6151
R1532 B.n305 B.n304 10.6151
R1533 B.n304 B.n229 10.6151
R1534 B.n300 B.n229 10.6151
R1535 B.n300 B.n299 10.6151
R1536 B.n299 B.n298 10.6151
R1537 B.n298 B.n231 10.6151
R1538 B.n294 B.n231 10.6151
R1539 B.n294 B.n293 10.6151
R1540 B.n293 B.n292 10.6151
R1541 B.n292 B.n233 10.6151
R1542 B.n288 B.n233 10.6151
R1543 B.n288 B.n287 10.6151
R1544 B.n287 B.n286 10.6151
R1545 B.n286 B.n235 10.6151
R1546 B.n282 B.n235 10.6151
R1547 B.n282 B.n281 10.6151
R1548 B.n281 B.n280 10.6151
R1549 B.n280 B.n237 10.6151
R1550 B.n276 B.n237 10.6151
R1551 B.n276 B.n275 10.6151
R1552 B.n275 B.n274 10.6151
R1553 B.n274 B.n239 10.6151
R1554 B.n270 B.n239 10.6151
R1555 B.n270 B.n269 10.6151
R1556 B.n269 B.n268 10.6151
R1557 B.n268 B.n241 10.6151
R1558 B.n264 B.n241 10.6151
R1559 B.n264 B.n263 10.6151
R1560 B.n263 B.n262 10.6151
R1561 B.n262 B.n243 10.6151
R1562 B.n258 B.n243 10.6151
R1563 B.n258 B.n257 10.6151
R1564 B.n257 B.n256 10.6151
R1565 B.n256 B.n245 10.6151
R1566 B.n252 B.n245 10.6151
R1567 B.n252 B.n251 10.6151
R1568 B.n251 B.n250 10.6151
R1569 B.n250 B.n247 10.6151
R1570 B.n247 B.n0 10.6151
R1571 B.n955 B.n1 10.6151
R1572 B.n955 B.n954 10.6151
R1573 B.n954 B.n953 10.6151
R1574 B.n953 B.n4 10.6151
R1575 B.n949 B.n4 10.6151
R1576 B.n949 B.n948 10.6151
R1577 B.n948 B.n947 10.6151
R1578 B.n947 B.n6 10.6151
R1579 B.n943 B.n6 10.6151
R1580 B.n943 B.n942 10.6151
R1581 B.n942 B.n941 10.6151
R1582 B.n941 B.n8 10.6151
R1583 B.n937 B.n8 10.6151
R1584 B.n937 B.n936 10.6151
R1585 B.n936 B.n935 10.6151
R1586 B.n935 B.n10 10.6151
R1587 B.n931 B.n10 10.6151
R1588 B.n931 B.n930 10.6151
R1589 B.n930 B.n929 10.6151
R1590 B.n929 B.n12 10.6151
R1591 B.n925 B.n12 10.6151
R1592 B.n925 B.n924 10.6151
R1593 B.n924 B.n923 10.6151
R1594 B.n923 B.n14 10.6151
R1595 B.n919 B.n14 10.6151
R1596 B.n919 B.n918 10.6151
R1597 B.n918 B.n917 10.6151
R1598 B.n917 B.n16 10.6151
R1599 B.n913 B.n16 10.6151
R1600 B.n913 B.n912 10.6151
R1601 B.n912 B.n911 10.6151
R1602 B.n911 B.n18 10.6151
R1603 B.n907 B.n18 10.6151
R1604 B.n907 B.n906 10.6151
R1605 B.n906 B.n905 10.6151
R1606 B.n905 B.n20 10.6151
R1607 B.n901 B.n20 10.6151
R1608 B.n901 B.n900 10.6151
R1609 B.n900 B.n899 10.6151
R1610 B.n899 B.n22 10.6151
R1611 B.n895 B.n22 10.6151
R1612 B.n895 B.n894 10.6151
R1613 B.n894 B.n893 10.6151
R1614 B.n893 B.n24 10.6151
R1615 B.n889 B.n24 10.6151
R1616 B.n889 B.n888 10.6151
R1617 B.n888 B.n887 10.6151
R1618 B.n887 B.n26 10.6151
R1619 B.n883 B.n26 10.6151
R1620 B.n883 B.n882 10.6151
R1621 B.n882 B.n881 10.6151
R1622 B.n881 B.n28 10.6151
R1623 B.n877 B.n28 10.6151
R1624 B.n877 B.n876 10.6151
R1625 B.n876 B.n875 10.6151
R1626 B.n875 B.n30 10.6151
R1627 B.n871 B.n30 10.6151
R1628 B.n871 B.n870 10.6151
R1629 B.n870 B.n869 10.6151
R1630 B.n869 B.n32 10.6151
R1631 B.n865 B.n32 10.6151
R1632 B.n865 B.n864 10.6151
R1633 B.n864 B.n863 10.6151
R1634 B.n62 B.n58 9.36635
R1635 B.n773 B.n772 9.36635
R1636 B.n414 B.n191 9.36635
R1637 B.n432 B.n431 9.36635
R1638 B.n959 B.n0 2.81026
R1639 B.n959 B.n1 2.81026
R1640 B.n787 B.n62 1.24928
R1641 B.n774 B.n773 1.24928
R1642 B.n417 B.n191 1.24928
R1643 B.n431 B.n430 1.24928
R1644 VP.n26 VP.n23 161.3
R1645 VP.n28 VP.n27 161.3
R1646 VP.n29 VP.n22 161.3
R1647 VP.n31 VP.n30 161.3
R1648 VP.n32 VP.n21 161.3
R1649 VP.n34 VP.n33 161.3
R1650 VP.n36 VP.n20 161.3
R1651 VP.n38 VP.n37 161.3
R1652 VP.n39 VP.n19 161.3
R1653 VP.n41 VP.n40 161.3
R1654 VP.n42 VP.n18 161.3
R1655 VP.n45 VP.n44 161.3
R1656 VP.n46 VP.n17 161.3
R1657 VP.n48 VP.n47 161.3
R1658 VP.n49 VP.n16 161.3
R1659 VP.n51 VP.n50 161.3
R1660 VP.n52 VP.n15 161.3
R1661 VP.n54 VP.n53 161.3
R1662 VP.n55 VP.n14 161.3
R1663 VP.n100 VP.n0 161.3
R1664 VP.n99 VP.n98 161.3
R1665 VP.n97 VP.n1 161.3
R1666 VP.n96 VP.n95 161.3
R1667 VP.n94 VP.n2 161.3
R1668 VP.n93 VP.n92 161.3
R1669 VP.n91 VP.n3 161.3
R1670 VP.n90 VP.n89 161.3
R1671 VP.n87 VP.n4 161.3
R1672 VP.n86 VP.n85 161.3
R1673 VP.n84 VP.n5 161.3
R1674 VP.n83 VP.n82 161.3
R1675 VP.n81 VP.n6 161.3
R1676 VP.n79 VP.n78 161.3
R1677 VP.n77 VP.n7 161.3
R1678 VP.n76 VP.n75 161.3
R1679 VP.n74 VP.n8 161.3
R1680 VP.n73 VP.n72 161.3
R1681 VP.n71 VP.n9 161.3
R1682 VP.n70 VP.n69 161.3
R1683 VP.n67 VP.n10 161.3
R1684 VP.n66 VP.n65 161.3
R1685 VP.n64 VP.n11 161.3
R1686 VP.n63 VP.n62 161.3
R1687 VP.n61 VP.n12 161.3
R1688 VP.n60 VP.n59 161.3
R1689 VP.n25 VP.t2 157.819
R1690 VP.n13 VP.t1 123.629
R1691 VP.n68 VP.t3 123.629
R1692 VP.n80 VP.t6 123.629
R1693 VP.n88 VP.t8 123.629
R1694 VP.n101 VP.t9 123.629
R1695 VP.n56 VP.t7 123.629
R1696 VP.n43 VP.t4 123.629
R1697 VP.n35 VP.t0 123.629
R1698 VP.n24 VP.t5 123.629
R1699 VP.n58 VP.n13 105.499
R1700 VP.n102 VP.n101 105.499
R1701 VP.n57 VP.n56 105.499
R1702 VP.n58 VP.n57 56.4693
R1703 VP.n75 VP.n74 56.0773
R1704 VP.n86 VP.n5 56.0773
R1705 VP.n41 VP.n19 56.0773
R1706 VP.n30 VP.n29 56.0773
R1707 VP.n25 VP.n24 52.6217
R1708 VP.n62 VP.n11 42.5146
R1709 VP.n95 VP.n1 42.5146
R1710 VP.n50 VP.n15 42.5146
R1711 VP.n66 VP.n11 38.6395
R1712 VP.n95 VP.n94 38.6395
R1713 VP.n50 VP.n49 38.6395
R1714 VP.n74 VP.n73 25.0767
R1715 VP.n87 VP.n86 25.0767
R1716 VP.n42 VP.n41 25.0767
R1717 VP.n29 VP.n28 25.0767
R1718 VP.n61 VP.n60 24.5923
R1719 VP.n62 VP.n61 24.5923
R1720 VP.n67 VP.n66 24.5923
R1721 VP.n69 VP.n67 24.5923
R1722 VP.n73 VP.n9 24.5923
R1723 VP.n75 VP.n7 24.5923
R1724 VP.n79 VP.n7 24.5923
R1725 VP.n82 VP.n81 24.5923
R1726 VP.n82 VP.n5 24.5923
R1727 VP.n89 VP.n87 24.5923
R1728 VP.n93 VP.n3 24.5923
R1729 VP.n94 VP.n93 24.5923
R1730 VP.n99 VP.n1 24.5923
R1731 VP.n100 VP.n99 24.5923
R1732 VP.n54 VP.n15 24.5923
R1733 VP.n55 VP.n54 24.5923
R1734 VP.n44 VP.n42 24.5923
R1735 VP.n48 VP.n17 24.5923
R1736 VP.n49 VP.n48 24.5923
R1737 VP.n30 VP.n21 24.5923
R1738 VP.n34 VP.n21 24.5923
R1739 VP.n37 VP.n36 24.5923
R1740 VP.n37 VP.n19 24.5923
R1741 VP.n28 VP.n23 24.5923
R1742 VP.n68 VP.n9 21.1495
R1743 VP.n89 VP.n88 21.1495
R1744 VP.n44 VP.n43 21.1495
R1745 VP.n24 VP.n23 21.1495
R1746 VP.n80 VP.n79 12.2964
R1747 VP.n81 VP.n80 12.2964
R1748 VP.n35 VP.n34 12.2964
R1749 VP.n36 VP.n35 12.2964
R1750 VP.n60 VP.n13 5.4107
R1751 VP.n101 VP.n100 5.4107
R1752 VP.n56 VP.n55 5.4107
R1753 VP.n26 VP.n25 4.94439
R1754 VP.n69 VP.n68 3.44336
R1755 VP.n88 VP.n3 3.44336
R1756 VP.n43 VP.n17 3.44336
R1757 VP.n57 VP.n14 0.278335
R1758 VP.n59 VP.n58 0.278335
R1759 VP.n102 VP.n0 0.278335
R1760 VP.n27 VP.n26 0.189894
R1761 VP.n27 VP.n22 0.189894
R1762 VP.n31 VP.n22 0.189894
R1763 VP.n32 VP.n31 0.189894
R1764 VP.n33 VP.n32 0.189894
R1765 VP.n33 VP.n20 0.189894
R1766 VP.n38 VP.n20 0.189894
R1767 VP.n39 VP.n38 0.189894
R1768 VP.n40 VP.n39 0.189894
R1769 VP.n40 VP.n18 0.189894
R1770 VP.n45 VP.n18 0.189894
R1771 VP.n46 VP.n45 0.189894
R1772 VP.n47 VP.n46 0.189894
R1773 VP.n47 VP.n16 0.189894
R1774 VP.n51 VP.n16 0.189894
R1775 VP.n52 VP.n51 0.189894
R1776 VP.n53 VP.n52 0.189894
R1777 VP.n53 VP.n14 0.189894
R1778 VP.n59 VP.n12 0.189894
R1779 VP.n63 VP.n12 0.189894
R1780 VP.n64 VP.n63 0.189894
R1781 VP.n65 VP.n64 0.189894
R1782 VP.n65 VP.n10 0.189894
R1783 VP.n70 VP.n10 0.189894
R1784 VP.n71 VP.n70 0.189894
R1785 VP.n72 VP.n71 0.189894
R1786 VP.n72 VP.n8 0.189894
R1787 VP.n76 VP.n8 0.189894
R1788 VP.n77 VP.n76 0.189894
R1789 VP.n78 VP.n77 0.189894
R1790 VP.n78 VP.n6 0.189894
R1791 VP.n83 VP.n6 0.189894
R1792 VP.n84 VP.n83 0.189894
R1793 VP.n85 VP.n84 0.189894
R1794 VP.n85 VP.n4 0.189894
R1795 VP.n90 VP.n4 0.189894
R1796 VP.n91 VP.n90 0.189894
R1797 VP.n92 VP.n91 0.189894
R1798 VP.n92 VP.n2 0.189894
R1799 VP.n96 VP.n2 0.189894
R1800 VP.n97 VP.n96 0.189894
R1801 VP.n98 VP.n97 0.189894
R1802 VP.n98 VP.n0 0.189894
R1803 VP VP.n102 0.153485
R1804 VDD1.n1 VDD1.t7 75.9127
R1805 VDD1.n3 VDD1.t8 75.9125
R1806 VDD1.n5 VDD1.n4 72.9487
R1807 VDD1.n7 VDD1.n6 70.948
R1808 VDD1.n1 VDD1.n0 70.948
R1809 VDD1.n3 VDD1.n2 70.948
R1810 VDD1.n7 VDD1.n5 51.294
R1811 VDD1.n6 VDD1.t5 2.22382
R1812 VDD1.n6 VDD1.t2 2.22382
R1813 VDD1.n0 VDD1.t4 2.22382
R1814 VDD1.n0 VDD1.t9 2.22382
R1815 VDD1.n4 VDD1.t1 2.22382
R1816 VDD1.n4 VDD1.t0 2.22382
R1817 VDD1.n2 VDD1.t6 2.22382
R1818 VDD1.n2 VDD1.t3 2.22382
R1819 VDD1 VDD1.n7 1.99834
R1820 VDD1 VDD1.n1 0.744035
R1821 VDD1.n5 VDD1.n3 0.630499
C0 w_n4786_n3892# VDD2 3.21963f
C1 VP VDD1 13.574201f
C2 VTAIL VDD2 11.6712f
C3 VN VDD1 0.154145f
C4 VP B 2.43215f
C5 VN B 1.38168f
C6 VDD1 w_n4786_n3892# 3.06308f
C7 VTAIL VDD1 11.6189f
C8 VDD1 VDD2 2.33663f
C9 VP VN 9.24286f
C10 w_n4786_n3892# B 11.702f
C11 VTAIL B 4.42913f
C12 VDD2 B 2.91406f
C13 VP w_n4786_n3892# 10.9682f
C14 VP VTAIL 13.7631f
C15 VP VDD2 0.615878f
C16 VN w_n4786_n3892# 10.3443f
C17 VN VTAIL 13.7488f
C18 VN VDD2 13.1168f
C19 VDD1 B 2.78641f
C20 VTAIL w_n4786_n3892# 3.60357f
C21 VDD2 VSUBS 2.3242f
C22 VDD1 VSUBS 2.130326f
C23 VTAIL VSUBS 1.453109f
C24 VN VSUBS 8.16145f
C25 VP VSUBS 4.645203f
C26 B VSUBS 5.898821f
C27 w_n4786_n3892# VSUBS 0.228522p
C28 VDD1.t7 VSUBS 3.59076f
C29 VDD1.t4 VSUBS 0.339579f
C30 VDD1.t9 VSUBS 0.339579f
C31 VDD1.n0 VSUBS 2.73125f
C32 VDD1.n1 VSUBS 1.81751f
C33 VDD1.t8 VSUBS 3.59076f
C34 VDD1.t6 VSUBS 0.339579f
C35 VDD1.t3 VSUBS 0.339579f
C36 VDD1.n2 VSUBS 2.73125f
C37 VDD1.n3 VSUBS 1.80785f
C38 VDD1.t1 VSUBS 0.339579f
C39 VDD1.t0 VSUBS 0.339579f
C40 VDD1.n4 VSUBS 2.75966f
C41 VDD1.n5 VSUBS 4.24442f
C42 VDD1.t5 VSUBS 0.339579f
C43 VDD1.t2 VSUBS 0.339579f
C44 VDD1.n6 VSUBS 2.73125f
C45 VDD1.n7 VSUBS 4.419f
C46 VP.n0 VSUBS 0.036061f
C47 VP.t9 VSUBS 3.1213f
C48 VP.n1 VSUBS 0.05347f
C49 VP.n2 VSUBS 0.027354f
C50 VP.n3 VSUBS 0.029189f
C51 VP.n4 VSUBS 0.027354f
C52 VP.n5 VSUBS 0.046507f
C53 VP.n6 VSUBS 0.027354f
C54 VP.t6 VSUBS 3.1213f
C55 VP.n7 VSUBS 0.050725f
C56 VP.n8 VSUBS 0.027354f
C57 VP.n9 VSUBS 0.047219f
C58 VP.n10 VSUBS 0.027354f
C59 VP.n11 VSUBS 0.022233f
C60 VP.n12 VSUBS 0.027354f
C61 VP.t1 VSUBS 3.1213f
C62 VP.n13 VSUBS 1.18302f
C63 VP.n14 VSUBS 0.036061f
C64 VP.t7 VSUBS 3.1213f
C65 VP.n15 VSUBS 0.05347f
C66 VP.n16 VSUBS 0.027354f
C67 VP.n17 VSUBS 0.029189f
C68 VP.n18 VSUBS 0.027354f
C69 VP.n19 VSUBS 0.046507f
C70 VP.n20 VSUBS 0.027354f
C71 VP.t0 VSUBS 3.1213f
C72 VP.n21 VSUBS 0.050725f
C73 VP.n22 VSUBS 0.027354f
C74 VP.n23 VSUBS 0.047219f
C75 VP.t2 VSUBS 3.39737f
C76 VP.t5 VSUBS 3.1213f
C77 VP.n24 VSUBS 1.18338f
C78 VP.n25 VSUBS 1.1313f
C79 VP.n26 VSUBS 0.288475f
C80 VP.n27 VSUBS 0.027354f
C81 VP.n28 VSUBS 0.051199f
C82 VP.n29 VSUBS 0.032545f
C83 VP.n30 VSUBS 0.046507f
C84 VP.n31 VSUBS 0.027354f
C85 VP.n32 VSUBS 0.027354f
C86 VP.n33 VSUBS 0.027354f
C87 VP.n34 VSUBS 0.038204f
C88 VP.n35 VSUBS 1.08975f
C89 VP.n36 VSUBS 0.038204f
C90 VP.n37 VSUBS 0.050725f
C91 VP.n38 VSUBS 0.027354f
C92 VP.n39 VSUBS 0.027354f
C93 VP.n40 VSUBS 0.027354f
C94 VP.n41 VSUBS 0.032545f
C95 VP.n42 VSUBS 0.051199f
C96 VP.t4 VSUBS 3.1213f
C97 VP.n43 VSUBS 1.08975f
C98 VP.n44 VSUBS 0.047219f
C99 VP.n45 VSUBS 0.027354f
C100 VP.n46 VSUBS 0.027354f
C101 VP.n47 VSUBS 0.027354f
C102 VP.n48 VSUBS 0.050725f
C103 VP.n49 VSUBS 0.054549f
C104 VP.n50 VSUBS 0.022233f
C105 VP.n51 VSUBS 0.027354f
C106 VP.n52 VSUBS 0.027354f
C107 VP.n53 VSUBS 0.027354f
C108 VP.n54 VSUBS 0.050725f
C109 VP.n55 VSUBS 0.031193f
C110 VP.n56 VSUBS 1.18302f
C111 VP.n57 VSUBS 1.81707f
C112 VP.n58 VSUBS 1.83453f
C113 VP.n59 VSUBS 0.036061f
C114 VP.n60 VSUBS 0.031193f
C115 VP.n61 VSUBS 0.050725f
C116 VP.n62 VSUBS 0.05347f
C117 VP.n63 VSUBS 0.027354f
C118 VP.n64 VSUBS 0.027354f
C119 VP.n65 VSUBS 0.027354f
C120 VP.n66 VSUBS 0.054549f
C121 VP.n67 VSUBS 0.050725f
C122 VP.t3 VSUBS 3.1213f
C123 VP.n68 VSUBS 1.08975f
C124 VP.n69 VSUBS 0.029189f
C125 VP.n70 VSUBS 0.027354f
C126 VP.n71 VSUBS 0.027354f
C127 VP.n72 VSUBS 0.027354f
C128 VP.n73 VSUBS 0.051199f
C129 VP.n74 VSUBS 0.032545f
C130 VP.n75 VSUBS 0.046507f
C131 VP.n76 VSUBS 0.027354f
C132 VP.n77 VSUBS 0.027354f
C133 VP.n78 VSUBS 0.027354f
C134 VP.n79 VSUBS 0.038204f
C135 VP.n80 VSUBS 1.08975f
C136 VP.n81 VSUBS 0.038204f
C137 VP.n82 VSUBS 0.050725f
C138 VP.n83 VSUBS 0.027354f
C139 VP.n84 VSUBS 0.027354f
C140 VP.n85 VSUBS 0.027354f
C141 VP.n86 VSUBS 0.032545f
C142 VP.n87 VSUBS 0.051199f
C143 VP.t8 VSUBS 3.1213f
C144 VP.n88 VSUBS 1.08975f
C145 VP.n89 VSUBS 0.047219f
C146 VP.n90 VSUBS 0.027354f
C147 VP.n91 VSUBS 0.027354f
C148 VP.n92 VSUBS 0.027354f
C149 VP.n93 VSUBS 0.050725f
C150 VP.n94 VSUBS 0.054549f
C151 VP.n95 VSUBS 0.022233f
C152 VP.n96 VSUBS 0.027354f
C153 VP.n97 VSUBS 0.027354f
C154 VP.n98 VSUBS 0.027354f
C155 VP.n99 VSUBS 0.050725f
C156 VP.n100 VSUBS 0.031193f
C157 VP.n101 VSUBS 1.18302f
C158 VP.n102 VSUBS 0.049965f
C159 B.n0 VSUBS 0.005412f
C160 B.n1 VSUBS 0.005412f
C161 B.n2 VSUBS 0.008559f
C162 B.n3 VSUBS 0.008559f
C163 B.n4 VSUBS 0.008559f
C164 B.n5 VSUBS 0.008559f
C165 B.n6 VSUBS 0.008559f
C166 B.n7 VSUBS 0.008559f
C167 B.n8 VSUBS 0.008559f
C168 B.n9 VSUBS 0.008559f
C169 B.n10 VSUBS 0.008559f
C170 B.n11 VSUBS 0.008559f
C171 B.n12 VSUBS 0.008559f
C172 B.n13 VSUBS 0.008559f
C173 B.n14 VSUBS 0.008559f
C174 B.n15 VSUBS 0.008559f
C175 B.n16 VSUBS 0.008559f
C176 B.n17 VSUBS 0.008559f
C177 B.n18 VSUBS 0.008559f
C178 B.n19 VSUBS 0.008559f
C179 B.n20 VSUBS 0.008559f
C180 B.n21 VSUBS 0.008559f
C181 B.n22 VSUBS 0.008559f
C182 B.n23 VSUBS 0.008559f
C183 B.n24 VSUBS 0.008559f
C184 B.n25 VSUBS 0.008559f
C185 B.n26 VSUBS 0.008559f
C186 B.n27 VSUBS 0.008559f
C187 B.n28 VSUBS 0.008559f
C188 B.n29 VSUBS 0.008559f
C189 B.n30 VSUBS 0.008559f
C190 B.n31 VSUBS 0.008559f
C191 B.n32 VSUBS 0.008559f
C192 B.n33 VSUBS 0.008559f
C193 B.n34 VSUBS 0.021921f
C194 B.n35 VSUBS 0.008559f
C195 B.n36 VSUBS 0.008559f
C196 B.n37 VSUBS 0.008559f
C197 B.n38 VSUBS 0.008559f
C198 B.n39 VSUBS 0.008559f
C199 B.n40 VSUBS 0.008559f
C200 B.n41 VSUBS 0.008559f
C201 B.n42 VSUBS 0.008559f
C202 B.n43 VSUBS 0.008559f
C203 B.n44 VSUBS 0.008559f
C204 B.n45 VSUBS 0.008559f
C205 B.n46 VSUBS 0.008559f
C206 B.n47 VSUBS 0.008559f
C207 B.n48 VSUBS 0.008559f
C208 B.n49 VSUBS 0.008559f
C209 B.n50 VSUBS 0.008559f
C210 B.n51 VSUBS 0.008559f
C211 B.n52 VSUBS 0.008559f
C212 B.n53 VSUBS 0.008559f
C213 B.n54 VSUBS 0.008559f
C214 B.n55 VSUBS 0.008559f
C215 B.n56 VSUBS 0.008559f
C216 B.n57 VSUBS 0.008559f
C217 B.n58 VSUBS 0.008055f
C218 B.n59 VSUBS 0.008559f
C219 B.t2 VSUBS 0.593768f
C220 B.t1 VSUBS 0.620934f
C221 B.t0 VSUBS 2.3063f
C222 B.n60 VSUBS 0.340639f
C223 B.n61 VSUBS 0.089232f
C224 B.n62 VSUBS 0.019829f
C225 B.n63 VSUBS 0.008559f
C226 B.n64 VSUBS 0.008559f
C227 B.n65 VSUBS 0.008559f
C228 B.n66 VSUBS 0.008559f
C229 B.t5 VSUBS 0.593753f
C230 B.t4 VSUBS 0.620921f
C231 B.t3 VSUBS 2.3063f
C232 B.n67 VSUBS 0.340652f
C233 B.n68 VSUBS 0.089247f
C234 B.n69 VSUBS 0.008559f
C235 B.n70 VSUBS 0.008559f
C236 B.n71 VSUBS 0.008559f
C237 B.n72 VSUBS 0.008559f
C238 B.n73 VSUBS 0.008559f
C239 B.n74 VSUBS 0.008559f
C240 B.n75 VSUBS 0.008559f
C241 B.n76 VSUBS 0.008559f
C242 B.n77 VSUBS 0.008559f
C243 B.n78 VSUBS 0.008559f
C244 B.n79 VSUBS 0.008559f
C245 B.n80 VSUBS 0.008559f
C246 B.n81 VSUBS 0.008559f
C247 B.n82 VSUBS 0.008559f
C248 B.n83 VSUBS 0.008559f
C249 B.n84 VSUBS 0.008559f
C250 B.n85 VSUBS 0.008559f
C251 B.n86 VSUBS 0.008559f
C252 B.n87 VSUBS 0.008559f
C253 B.n88 VSUBS 0.008559f
C254 B.n89 VSUBS 0.008559f
C255 B.n90 VSUBS 0.008559f
C256 B.n91 VSUBS 0.008559f
C257 B.n92 VSUBS 0.008559f
C258 B.n93 VSUBS 0.021787f
C259 B.n94 VSUBS 0.008559f
C260 B.n95 VSUBS 0.008559f
C261 B.n96 VSUBS 0.008559f
C262 B.n97 VSUBS 0.008559f
C263 B.n98 VSUBS 0.008559f
C264 B.n99 VSUBS 0.008559f
C265 B.n100 VSUBS 0.008559f
C266 B.n101 VSUBS 0.008559f
C267 B.n102 VSUBS 0.008559f
C268 B.n103 VSUBS 0.008559f
C269 B.n104 VSUBS 0.008559f
C270 B.n105 VSUBS 0.008559f
C271 B.n106 VSUBS 0.008559f
C272 B.n107 VSUBS 0.008559f
C273 B.n108 VSUBS 0.008559f
C274 B.n109 VSUBS 0.008559f
C275 B.n110 VSUBS 0.008559f
C276 B.n111 VSUBS 0.008559f
C277 B.n112 VSUBS 0.008559f
C278 B.n113 VSUBS 0.008559f
C279 B.n114 VSUBS 0.008559f
C280 B.n115 VSUBS 0.008559f
C281 B.n116 VSUBS 0.008559f
C282 B.n117 VSUBS 0.008559f
C283 B.n118 VSUBS 0.008559f
C284 B.n119 VSUBS 0.008559f
C285 B.n120 VSUBS 0.008559f
C286 B.n121 VSUBS 0.008559f
C287 B.n122 VSUBS 0.008559f
C288 B.n123 VSUBS 0.008559f
C289 B.n124 VSUBS 0.008559f
C290 B.n125 VSUBS 0.008559f
C291 B.n126 VSUBS 0.008559f
C292 B.n127 VSUBS 0.008559f
C293 B.n128 VSUBS 0.008559f
C294 B.n129 VSUBS 0.008559f
C295 B.n130 VSUBS 0.008559f
C296 B.n131 VSUBS 0.008559f
C297 B.n132 VSUBS 0.008559f
C298 B.n133 VSUBS 0.008559f
C299 B.n134 VSUBS 0.008559f
C300 B.n135 VSUBS 0.008559f
C301 B.n136 VSUBS 0.008559f
C302 B.n137 VSUBS 0.008559f
C303 B.n138 VSUBS 0.008559f
C304 B.n139 VSUBS 0.008559f
C305 B.n140 VSUBS 0.008559f
C306 B.n141 VSUBS 0.008559f
C307 B.n142 VSUBS 0.008559f
C308 B.n143 VSUBS 0.008559f
C309 B.n144 VSUBS 0.008559f
C310 B.n145 VSUBS 0.008559f
C311 B.n146 VSUBS 0.008559f
C312 B.n147 VSUBS 0.008559f
C313 B.n148 VSUBS 0.008559f
C314 B.n149 VSUBS 0.008559f
C315 B.n150 VSUBS 0.008559f
C316 B.n151 VSUBS 0.008559f
C317 B.n152 VSUBS 0.008559f
C318 B.n153 VSUBS 0.008559f
C319 B.n154 VSUBS 0.008559f
C320 B.n155 VSUBS 0.008559f
C321 B.n156 VSUBS 0.008559f
C322 B.n157 VSUBS 0.020872f
C323 B.n158 VSUBS 0.008559f
C324 B.n159 VSUBS 0.008559f
C325 B.n160 VSUBS 0.008559f
C326 B.n161 VSUBS 0.008559f
C327 B.n162 VSUBS 0.008559f
C328 B.n163 VSUBS 0.008559f
C329 B.n164 VSUBS 0.008559f
C330 B.n165 VSUBS 0.008559f
C331 B.n166 VSUBS 0.008559f
C332 B.n167 VSUBS 0.008559f
C333 B.n168 VSUBS 0.008559f
C334 B.n169 VSUBS 0.008559f
C335 B.n170 VSUBS 0.008559f
C336 B.n171 VSUBS 0.008559f
C337 B.n172 VSUBS 0.008559f
C338 B.n173 VSUBS 0.008559f
C339 B.n174 VSUBS 0.008559f
C340 B.n175 VSUBS 0.008559f
C341 B.n176 VSUBS 0.008559f
C342 B.n177 VSUBS 0.008559f
C343 B.n178 VSUBS 0.008559f
C344 B.n179 VSUBS 0.008559f
C345 B.n180 VSUBS 0.008559f
C346 B.n181 VSUBS 0.008559f
C347 B.n182 VSUBS 0.008559f
C348 B.t10 VSUBS 0.593753f
C349 B.t11 VSUBS 0.620921f
C350 B.t9 VSUBS 2.3063f
C351 B.n183 VSUBS 0.340652f
C352 B.n184 VSUBS 0.089247f
C353 B.n185 VSUBS 0.008559f
C354 B.n186 VSUBS 0.008559f
C355 B.n187 VSUBS 0.008559f
C356 B.n188 VSUBS 0.008559f
C357 B.t7 VSUBS 0.593768f
C358 B.t8 VSUBS 0.620934f
C359 B.t6 VSUBS 2.3063f
C360 B.n189 VSUBS 0.340639f
C361 B.n190 VSUBS 0.089232f
C362 B.n191 VSUBS 0.019829f
C363 B.n192 VSUBS 0.008559f
C364 B.n193 VSUBS 0.008559f
C365 B.n194 VSUBS 0.008559f
C366 B.n195 VSUBS 0.008559f
C367 B.n196 VSUBS 0.008559f
C368 B.n197 VSUBS 0.008559f
C369 B.n198 VSUBS 0.008559f
C370 B.n199 VSUBS 0.008559f
C371 B.n200 VSUBS 0.008559f
C372 B.n201 VSUBS 0.008559f
C373 B.n202 VSUBS 0.008559f
C374 B.n203 VSUBS 0.008559f
C375 B.n204 VSUBS 0.008559f
C376 B.n205 VSUBS 0.008559f
C377 B.n206 VSUBS 0.008559f
C378 B.n207 VSUBS 0.008559f
C379 B.n208 VSUBS 0.008559f
C380 B.n209 VSUBS 0.008559f
C381 B.n210 VSUBS 0.008559f
C382 B.n211 VSUBS 0.008559f
C383 B.n212 VSUBS 0.008559f
C384 B.n213 VSUBS 0.008559f
C385 B.n214 VSUBS 0.008559f
C386 B.n215 VSUBS 0.008559f
C387 B.n216 VSUBS 0.020872f
C388 B.n217 VSUBS 0.008559f
C389 B.n218 VSUBS 0.008559f
C390 B.n219 VSUBS 0.008559f
C391 B.n220 VSUBS 0.008559f
C392 B.n221 VSUBS 0.008559f
C393 B.n222 VSUBS 0.008559f
C394 B.n223 VSUBS 0.008559f
C395 B.n224 VSUBS 0.008559f
C396 B.n225 VSUBS 0.008559f
C397 B.n226 VSUBS 0.008559f
C398 B.n227 VSUBS 0.008559f
C399 B.n228 VSUBS 0.008559f
C400 B.n229 VSUBS 0.008559f
C401 B.n230 VSUBS 0.008559f
C402 B.n231 VSUBS 0.008559f
C403 B.n232 VSUBS 0.008559f
C404 B.n233 VSUBS 0.008559f
C405 B.n234 VSUBS 0.008559f
C406 B.n235 VSUBS 0.008559f
C407 B.n236 VSUBS 0.008559f
C408 B.n237 VSUBS 0.008559f
C409 B.n238 VSUBS 0.008559f
C410 B.n239 VSUBS 0.008559f
C411 B.n240 VSUBS 0.008559f
C412 B.n241 VSUBS 0.008559f
C413 B.n242 VSUBS 0.008559f
C414 B.n243 VSUBS 0.008559f
C415 B.n244 VSUBS 0.008559f
C416 B.n245 VSUBS 0.008559f
C417 B.n246 VSUBS 0.008559f
C418 B.n247 VSUBS 0.008559f
C419 B.n248 VSUBS 0.008559f
C420 B.n249 VSUBS 0.008559f
C421 B.n250 VSUBS 0.008559f
C422 B.n251 VSUBS 0.008559f
C423 B.n252 VSUBS 0.008559f
C424 B.n253 VSUBS 0.008559f
C425 B.n254 VSUBS 0.008559f
C426 B.n255 VSUBS 0.008559f
C427 B.n256 VSUBS 0.008559f
C428 B.n257 VSUBS 0.008559f
C429 B.n258 VSUBS 0.008559f
C430 B.n259 VSUBS 0.008559f
C431 B.n260 VSUBS 0.008559f
C432 B.n261 VSUBS 0.008559f
C433 B.n262 VSUBS 0.008559f
C434 B.n263 VSUBS 0.008559f
C435 B.n264 VSUBS 0.008559f
C436 B.n265 VSUBS 0.008559f
C437 B.n266 VSUBS 0.008559f
C438 B.n267 VSUBS 0.008559f
C439 B.n268 VSUBS 0.008559f
C440 B.n269 VSUBS 0.008559f
C441 B.n270 VSUBS 0.008559f
C442 B.n271 VSUBS 0.008559f
C443 B.n272 VSUBS 0.008559f
C444 B.n273 VSUBS 0.008559f
C445 B.n274 VSUBS 0.008559f
C446 B.n275 VSUBS 0.008559f
C447 B.n276 VSUBS 0.008559f
C448 B.n277 VSUBS 0.008559f
C449 B.n278 VSUBS 0.008559f
C450 B.n279 VSUBS 0.008559f
C451 B.n280 VSUBS 0.008559f
C452 B.n281 VSUBS 0.008559f
C453 B.n282 VSUBS 0.008559f
C454 B.n283 VSUBS 0.008559f
C455 B.n284 VSUBS 0.008559f
C456 B.n285 VSUBS 0.008559f
C457 B.n286 VSUBS 0.008559f
C458 B.n287 VSUBS 0.008559f
C459 B.n288 VSUBS 0.008559f
C460 B.n289 VSUBS 0.008559f
C461 B.n290 VSUBS 0.008559f
C462 B.n291 VSUBS 0.008559f
C463 B.n292 VSUBS 0.008559f
C464 B.n293 VSUBS 0.008559f
C465 B.n294 VSUBS 0.008559f
C466 B.n295 VSUBS 0.008559f
C467 B.n296 VSUBS 0.008559f
C468 B.n297 VSUBS 0.008559f
C469 B.n298 VSUBS 0.008559f
C470 B.n299 VSUBS 0.008559f
C471 B.n300 VSUBS 0.008559f
C472 B.n301 VSUBS 0.008559f
C473 B.n302 VSUBS 0.008559f
C474 B.n303 VSUBS 0.008559f
C475 B.n304 VSUBS 0.008559f
C476 B.n305 VSUBS 0.008559f
C477 B.n306 VSUBS 0.008559f
C478 B.n307 VSUBS 0.008559f
C479 B.n308 VSUBS 0.008559f
C480 B.n309 VSUBS 0.008559f
C481 B.n310 VSUBS 0.008559f
C482 B.n311 VSUBS 0.008559f
C483 B.n312 VSUBS 0.008559f
C484 B.n313 VSUBS 0.008559f
C485 B.n314 VSUBS 0.008559f
C486 B.n315 VSUBS 0.008559f
C487 B.n316 VSUBS 0.008559f
C488 B.n317 VSUBS 0.008559f
C489 B.n318 VSUBS 0.008559f
C490 B.n319 VSUBS 0.008559f
C491 B.n320 VSUBS 0.008559f
C492 B.n321 VSUBS 0.008559f
C493 B.n322 VSUBS 0.008559f
C494 B.n323 VSUBS 0.008559f
C495 B.n324 VSUBS 0.008559f
C496 B.n325 VSUBS 0.008559f
C497 B.n326 VSUBS 0.008559f
C498 B.n327 VSUBS 0.008559f
C499 B.n328 VSUBS 0.008559f
C500 B.n329 VSUBS 0.008559f
C501 B.n330 VSUBS 0.008559f
C502 B.n331 VSUBS 0.008559f
C503 B.n332 VSUBS 0.008559f
C504 B.n333 VSUBS 0.008559f
C505 B.n334 VSUBS 0.008559f
C506 B.n335 VSUBS 0.008559f
C507 B.n336 VSUBS 0.008559f
C508 B.n337 VSUBS 0.008559f
C509 B.n338 VSUBS 0.008559f
C510 B.n339 VSUBS 0.008559f
C511 B.n340 VSUBS 0.008559f
C512 B.n341 VSUBS 0.020872f
C513 B.n342 VSUBS 0.021921f
C514 B.n343 VSUBS 0.021921f
C515 B.n344 VSUBS 0.008559f
C516 B.n345 VSUBS 0.008559f
C517 B.n346 VSUBS 0.008559f
C518 B.n347 VSUBS 0.008559f
C519 B.n348 VSUBS 0.008559f
C520 B.n349 VSUBS 0.008559f
C521 B.n350 VSUBS 0.008559f
C522 B.n351 VSUBS 0.008559f
C523 B.n352 VSUBS 0.008559f
C524 B.n353 VSUBS 0.008559f
C525 B.n354 VSUBS 0.008559f
C526 B.n355 VSUBS 0.008559f
C527 B.n356 VSUBS 0.008559f
C528 B.n357 VSUBS 0.008559f
C529 B.n358 VSUBS 0.008559f
C530 B.n359 VSUBS 0.008559f
C531 B.n360 VSUBS 0.008559f
C532 B.n361 VSUBS 0.008559f
C533 B.n362 VSUBS 0.008559f
C534 B.n363 VSUBS 0.008559f
C535 B.n364 VSUBS 0.008559f
C536 B.n365 VSUBS 0.008559f
C537 B.n366 VSUBS 0.008559f
C538 B.n367 VSUBS 0.008559f
C539 B.n368 VSUBS 0.008559f
C540 B.n369 VSUBS 0.008559f
C541 B.n370 VSUBS 0.008559f
C542 B.n371 VSUBS 0.008559f
C543 B.n372 VSUBS 0.008559f
C544 B.n373 VSUBS 0.008559f
C545 B.n374 VSUBS 0.008559f
C546 B.n375 VSUBS 0.008559f
C547 B.n376 VSUBS 0.008559f
C548 B.n377 VSUBS 0.008559f
C549 B.n378 VSUBS 0.008559f
C550 B.n379 VSUBS 0.008559f
C551 B.n380 VSUBS 0.008559f
C552 B.n381 VSUBS 0.008559f
C553 B.n382 VSUBS 0.008559f
C554 B.n383 VSUBS 0.008559f
C555 B.n384 VSUBS 0.008559f
C556 B.n385 VSUBS 0.008559f
C557 B.n386 VSUBS 0.008559f
C558 B.n387 VSUBS 0.008559f
C559 B.n388 VSUBS 0.008559f
C560 B.n389 VSUBS 0.008559f
C561 B.n390 VSUBS 0.008559f
C562 B.n391 VSUBS 0.008559f
C563 B.n392 VSUBS 0.008559f
C564 B.n393 VSUBS 0.008559f
C565 B.n394 VSUBS 0.008559f
C566 B.n395 VSUBS 0.008559f
C567 B.n396 VSUBS 0.008559f
C568 B.n397 VSUBS 0.008559f
C569 B.n398 VSUBS 0.008559f
C570 B.n399 VSUBS 0.008559f
C571 B.n400 VSUBS 0.008559f
C572 B.n401 VSUBS 0.008559f
C573 B.n402 VSUBS 0.008559f
C574 B.n403 VSUBS 0.008559f
C575 B.n404 VSUBS 0.008559f
C576 B.n405 VSUBS 0.008559f
C577 B.n406 VSUBS 0.008559f
C578 B.n407 VSUBS 0.008559f
C579 B.n408 VSUBS 0.008559f
C580 B.n409 VSUBS 0.008559f
C581 B.n410 VSUBS 0.008559f
C582 B.n411 VSUBS 0.008559f
C583 B.n412 VSUBS 0.008559f
C584 B.n413 VSUBS 0.008559f
C585 B.n414 VSUBS 0.008055f
C586 B.n415 VSUBS 0.008559f
C587 B.n416 VSUBS 0.008559f
C588 B.n417 VSUBS 0.004783f
C589 B.n418 VSUBS 0.008559f
C590 B.n419 VSUBS 0.008559f
C591 B.n420 VSUBS 0.008559f
C592 B.n421 VSUBS 0.008559f
C593 B.n422 VSUBS 0.008559f
C594 B.n423 VSUBS 0.008559f
C595 B.n424 VSUBS 0.008559f
C596 B.n425 VSUBS 0.008559f
C597 B.n426 VSUBS 0.008559f
C598 B.n427 VSUBS 0.008559f
C599 B.n428 VSUBS 0.008559f
C600 B.n429 VSUBS 0.008559f
C601 B.n430 VSUBS 0.004783f
C602 B.n431 VSUBS 0.019829f
C603 B.n432 VSUBS 0.008055f
C604 B.n433 VSUBS 0.008559f
C605 B.n434 VSUBS 0.008559f
C606 B.n435 VSUBS 0.008559f
C607 B.n436 VSUBS 0.008559f
C608 B.n437 VSUBS 0.008559f
C609 B.n438 VSUBS 0.008559f
C610 B.n439 VSUBS 0.008559f
C611 B.n440 VSUBS 0.008559f
C612 B.n441 VSUBS 0.008559f
C613 B.n442 VSUBS 0.008559f
C614 B.n443 VSUBS 0.008559f
C615 B.n444 VSUBS 0.008559f
C616 B.n445 VSUBS 0.008559f
C617 B.n446 VSUBS 0.008559f
C618 B.n447 VSUBS 0.008559f
C619 B.n448 VSUBS 0.008559f
C620 B.n449 VSUBS 0.008559f
C621 B.n450 VSUBS 0.008559f
C622 B.n451 VSUBS 0.008559f
C623 B.n452 VSUBS 0.008559f
C624 B.n453 VSUBS 0.008559f
C625 B.n454 VSUBS 0.008559f
C626 B.n455 VSUBS 0.008559f
C627 B.n456 VSUBS 0.008559f
C628 B.n457 VSUBS 0.008559f
C629 B.n458 VSUBS 0.008559f
C630 B.n459 VSUBS 0.008559f
C631 B.n460 VSUBS 0.008559f
C632 B.n461 VSUBS 0.008559f
C633 B.n462 VSUBS 0.008559f
C634 B.n463 VSUBS 0.008559f
C635 B.n464 VSUBS 0.008559f
C636 B.n465 VSUBS 0.008559f
C637 B.n466 VSUBS 0.008559f
C638 B.n467 VSUBS 0.008559f
C639 B.n468 VSUBS 0.008559f
C640 B.n469 VSUBS 0.008559f
C641 B.n470 VSUBS 0.008559f
C642 B.n471 VSUBS 0.008559f
C643 B.n472 VSUBS 0.008559f
C644 B.n473 VSUBS 0.008559f
C645 B.n474 VSUBS 0.008559f
C646 B.n475 VSUBS 0.008559f
C647 B.n476 VSUBS 0.008559f
C648 B.n477 VSUBS 0.008559f
C649 B.n478 VSUBS 0.008559f
C650 B.n479 VSUBS 0.008559f
C651 B.n480 VSUBS 0.008559f
C652 B.n481 VSUBS 0.008559f
C653 B.n482 VSUBS 0.008559f
C654 B.n483 VSUBS 0.008559f
C655 B.n484 VSUBS 0.008559f
C656 B.n485 VSUBS 0.008559f
C657 B.n486 VSUBS 0.008559f
C658 B.n487 VSUBS 0.008559f
C659 B.n488 VSUBS 0.008559f
C660 B.n489 VSUBS 0.008559f
C661 B.n490 VSUBS 0.008559f
C662 B.n491 VSUBS 0.008559f
C663 B.n492 VSUBS 0.008559f
C664 B.n493 VSUBS 0.008559f
C665 B.n494 VSUBS 0.008559f
C666 B.n495 VSUBS 0.008559f
C667 B.n496 VSUBS 0.008559f
C668 B.n497 VSUBS 0.008559f
C669 B.n498 VSUBS 0.008559f
C670 B.n499 VSUBS 0.008559f
C671 B.n500 VSUBS 0.008559f
C672 B.n501 VSUBS 0.008559f
C673 B.n502 VSUBS 0.008559f
C674 B.n503 VSUBS 0.008559f
C675 B.n504 VSUBS 0.021921f
C676 B.n505 VSUBS 0.021921f
C677 B.n506 VSUBS 0.020872f
C678 B.n507 VSUBS 0.008559f
C679 B.n508 VSUBS 0.008559f
C680 B.n509 VSUBS 0.008559f
C681 B.n510 VSUBS 0.008559f
C682 B.n511 VSUBS 0.008559f
C683 B.n512 VSUBS 0.008559f
C684 B.n513 VSUBS 0.008559f
C685 B.n514 VSUBS 0.008559f
C686 B.n515 VSUBS 0.008559f
C687 B.n516 VSUBS 0.008559f
C688 B.n517 VSUBS 0.008559f
C689 B.n518 VSUBS 0.008559f
C690 B.n519 VSUBS 0.008559f
C691 B.n520 VSUBS 0.008559f
C692 B.n521 VSUBS 0.008559f
C693 B.n522 VSUBS 0.008559f
C694 B.n523 VSUBS 0.008559f
C695 B.n524 VSUBS 0.008559f
C696 B.n525 VSUBS 0.008559f
C697 B.n526 VSUBS 0.008559f
C698 B.n527 VSUBS 0.008559f
C699 B.n528 VSUBS 0.008559f
C700 B.n529 VSUBS 0.008559f
C701 B.n530 VSUBS 0.008559f
C702 B.n531 VSUBS 0.008559f
C703 B.n532 VSUBS 0.008559f
C704 B.n533 VSUBS 0.008559f
C705 B.n534 VSUBS 0.008559f
C706 B.n535 VSUBS 0.008559f
C707 B.n536 VSUBS 0.008559f
C708 B.n537 VSUBS 0.008559f
C709 B.n538 VSUBS 0.008559f
C710 B.n539 VSUBS 0.008559f
C711 B.n540 VSUBS 0.008559f
C712 B.n541 VSUBS 0.008559f
C713 B.n542 VSUBS 0.008559f
C714 B.n543 VSUBS 0.008559f
C715 B.n544 VSUBS 0.008559f
C716 B.n545 VSUBS 0.008559f
C717 B.n546 VSUBS 0.008559f
C718 B.n547 VSUBS 0.008559f
C719 B.n548 VSUBS 0.008559f
C720 B.n549 VSUBS 0.008559f
C721 B.n550 VSUBS 0.008559f
C722 B.n551 VSUBS 0.008559f
C723 B.n552 VSUBS 0.008559f
C724 B.n553 VSUBS 0.008559f
C725 B.n554 VSUBS 0.008559f
C726 B.n555 VSUBS 0.008559f
C727 B.n556 VSUBS 0.008559f
C728 B.n557 VSUBS 0.008559f
C729 B.n558 VSUBS 0.008559f
C730 B.n559 VSUBS 0.008559f
C731 B.n560 VSUBS 0.008559f
C732 B.n561 VSUBS 0.008559f
C733 B.n562 VSUBS 0.008559f
C734 B.n563 VSUBS 0.008559f
C735 B.n564 VSUBS 0.008559f
C736 B.n565 VSUBS 0.008559f
C737 B.n566 VSUBS 0.008559f
C738 B.n567 VSUBS 0.008559f
C739 B.n568 VSUBS 0.008559f
C740 B.n569 VSUBS 0.008559f
C741 B.n570 VSUBS 0.008559f
C742 B.n571 VSUBS 0.008559f
C743 B.n572 VSUBS 0.008559f
C744 B.n573 VSUBS 0.008559f
C745 B.n574 VSUBS 0.008559f
C746 B.n575 VSUBS 0.008559f
C747 B.n576 VSUBS 0.008559f
C748 B.n577 VSUBS 0.008559f
C749 B.n578 VSUBS 0.008559f
C750 B.n579 VSUBS 0.008559f
C751 B.n580 VSUBS 0.008559f
C752 B.n581 VSUBS 0.008559f
C753 B.n582 VSUBS 0.008559f
C754 B.n583 VSUBS 0.008559f
C755 B.n584 VSUBS 0.008559f
C756 B.n585 VSUBS 0.008559f
C757 B.n586 VSUBS 0.008559f
C758 B.n587 VSUBS 0.008559f
C759 B.n588 VSUBS 0.008559f
C760 B.n589 VSUBS 0.008559f
C761 B.n590 VSUBS 0.008559f
C762 B.n591 VSUBS 0.008559f
C763 B.n592 VSUBS 0.008559f
C764 B.n593 VSUBS 0.008559f
C765 B.n594 VSUBS 0.008559f
C766 B.n595 VSUBS 0.008559f
C767 B.n596 VSUBS 0.008559f
C768 B.n597 VSUBS 0.008559f
C769 B.n598 VSUBS 0.008559f
C770 B.n599 VSUBS 0.008559f
C771 B.n600 VSUBS 0.008559f
C772 B.n601 VSUBS 0.008559f
C773 B.n602 VSUBS 0.008559f
C774 B.n603 VSUBS 0.008559f
C775 B.n604 VSUBS 0.008559f
C776 B.n605 VSUBS 0.008559f
C777 B.n606 VSUBS 0.008559f
C778 B.n607 VSUBS 0.008559f
C779 B.n608 VSUBS 0.008559f
C780 B.n609 VSUBS 0.008559f
C781 B.n610 VSUBS 0.008559f
C782 B.n611 VSUBS 0.008559f
C783 B.n612 VSUBS 0.008559f
C784 B.n613 VSUBS 0.008559f
C785 B.n614 VSUBS 0.008559f
C786 B.n615 VSUBS 0.008559f
C787 B.n616 VSUBS 0.008559f
C788 B.n617 VSUBS 0.008559f
C789 B.n618 VSUBS 0.008559f
C790 B.n619 VSUBS 0.008559f
C791 B.n620 VSUBS 0.008559f
C792 B.n621 VSUBS 0.008559f
C793 B.n622 VSUBS 0.008559f
C794 B.n623 VSUBS 0.008559f
C795 B.n624 VSUBS 0.008559f
C796 B.n625 VSUBS 0.008559f
C797 B.n626 VSUBS 0.008559f
C798 B.n627 VSUBS 0.008559f
C799 B.n628 VSUBS 0.008559f
C800 B.n629 VSUBS 0.008559f
C801 B.n630 VSUBS 0.008559f
C802 B.n631 VSUBS 0.008559f
C803 B.n632 VSUBS 0.008559f
C804 B.n633 VSUBS 0.008559f
C805 B.n634 VSUBS 0.008559f
C806 B.n635 VSUBS 0.008559f
C807 B.n636 VSUBS 0.008559f
C808 B.n637 VSUBS 0.008559f
C809 B.n638 VSUBS 0.008559f
C810 B.n639 VSUBS 0.008559f
C811 B.n640 VSUBS 0.008559f
C812 B.n641 VSUBS 0.008559f
C813 B.n642 VSUBS 0.008559f
C814 B.n643 VSUBS 0.008559f
C815 B.n644 VSUBS 0.008559f
C816 B.n645 VSUBS 0.008559f
C817 B.n646 VSUBS 0.008559f
C818 B.n647 VSUBS 0.008559f
C819 B.n648 VSUBS 0.008559f
C820 B.n649 VSUBS 0.008559f
C821 B.n650 VSUBS 0.008559f
C822 B.n651 VSUBS 0.008559f
C823 B.n652 VSUBS 0.008559f
C824 B.n653 VSUBS 0.008559f
C825 B.n654 VSUBS 0.008559f
C826 B.n655 VSUBS 0.008559f
C827 B.n656 VSUBS 0.008559f
C828 B.n657 VSUBS 0.008559f
C829 B.n658 VSUBS 0.008559f
C830 B.n659 VSUBS 0.008559f
C831 B.n660 VSUBS 0.008559f
C832 B.n661 VSUBS 0.008559f
C833 B.n662 VSUBS 0.008559f
C834 B.n663 VSUBS 0.008559f
C835 B.n664 VSUBS 0.008559f
C836 B.n665 VSUBS 0.008559f
C837 B.n666 VSUBS 0.008559f
C838 B.n667 VSUBS 0.008559f
C839 B.n668 VSUBS 0.008559f
C840 B.n669 VSUBS 0.008559f
C841 B.n670 VSUBS 0.008559f
C842 B.n671 VSUBS 0.008559f
C843 B.n672 VSUBS 0.008559f
C844 B.n673 VSUBS 0.008559f
C845 B.n674 VSUBS 0.008559f
C846 B.n675 VSUBS 0.008559f
C847 B.n676 VSUBS 0.008559f
C848 B.n677 VSUBS 0.008559f
C849 B.n678 VSUBS 0.008559f
C850 B.n679 VSUBS 0.008559f
C851 B.n680 VSUBS 0.008559f
C852 B.n681 VSUBS 0.008559f
C853 B.n682 VSUBS 0.008559f
C854 B.n683 VSUBS 0.008559f
C855 B.n684 VSUBS 0.008559f
C856 B.n685 VSUBS 0.008559f
C857 B.n686 VSUBS 0.008559f
C858 B.n687 VSUBS 0.008559f
C859 B.n688 VSUBS 0.008559f
C860 B.n689 VSUBS 0.008559f
C861 B.n690 VSUBS 0.008559f
C862 B.n691 VSUBS 0.008559f
C863 B.n692 VSUBS 0.008559f
C864 B.n693 VSUBS 0.008559f
C865 B.n694 VSUBS 0.008559f
C866 B.n695 VSUBS 0.008559f
C867 B.n696 VSUBS 0.008559f
C868 B.n697 VSUBS 0.008559f
C869 B.n698 VSUBS 0.020872f
C870 B.n699 VSUBS 0.021921f
C871 B.n700 VSUBS 0.021006f
C872 B.n701 VSUBS 0.008559f
C873 B.n702 VSUBS 0.008559f
C874 B.n703 VSUBS 0.008559f
C875 B.n704 VSUBS 0.008559f
C876 B.n705 VSUBS 0.008559f
C877 B.n706 VSUBS 0.008559f
C878 B.n707 VSUBS 0.008559f
C879 B.n708 VSUBS 0.008559f
C880 B.n709 VSUBS 0.008559f
C881 B.n710 VSUBS 0.008559f
C882 B.n711 VSUBS 0.008559f
C883 B.n712 VSUBS 0.008559f
C884 B.n713 VSUBS 0.008559f
C885 B.n714 VSUBS 0.008559f
C886 B.n715 VSUBS 0.008559f
C887 B.n716 VSUBS 0.008559f
C888 B.n717 VSUBS 0.008559f
C889 B.n718 VSUBS 0.008559f
C890 B.n719 VSUBS 0.008559f
C891 B.n720 VSUBS 0.008559f
C892 B.n721 VSUBS 0.008559f
C893 B.n722 VSUBS 0.008559f
C894 B.n723 VSUBS 0.008559f
C895 B.n724 VSUBS 0.008559f
C896 B.n725 VSUBS 0.008559f
C897 B.n726 VSUBS 0.008559f
C898 B.n727 VSUBS 0.008559f
C899 B.n728 VSUBS 0.008559f
C900 B.n729 VSUBS 0.008559f
C901 B.n730 VSUBS 0.008559f
C902 B.n731 VSUBS 0.008559f
C903 B.n732 VSUBS 0.008559f
C904 B.n733 VSUBS 0.008559f
C905 B.n734 VSUBS 0.008559f
C906 B.n735 VSUBS 0.008559f
C907 B.n736 VSUBS 0.008559f
C908 B.n737 VSUBS 0.008559f
C909 B.n738 VSUBS 0.008559f
C910 B.n739 VSUBS 0.008559f
C911 B.n740 VSUBS 0.008559f
C912 B.n741 VSUBS 0.008559f
C913 B.n742 VSUBS 0.008559f
C914 B.n743 VSUBS 0.008559f
C915 B.n744 VSUBS 0.008559f
C916 B.n745 VSUBS 0.008559f
C917 B.n746 VSUBS 0.008559f
C918 B.n747 VSUBS 0.008559f
C919 B.n748 VSUBS 0.008559f
C920 B.n749 VSUBS 0.008559f
C921 B.n750 VSUBS 0.008559f
C922 B.n751 VSUBS 0.008559f
C923 B.n752 VSUBS 0.008559f
C924 B.n753 VSUBS 0.008559f
C925 B.n754 VSUBS 0.008559f
C926 B.n755 VSUBS 0.008559f
C927 B.n756 VSUBS 0.008559f
C928 B.n757 VSUBS 0.008559f
C929 B.n758 VSUBS 0.008559f
C930 B.n759 VSUBS 0.008559f
C931 B.n760 VSUBS 0.008559f
C932 B.n761 VSUBS 0.008559f
C933 B.n762 VSUBS 0.008559f
C934 B.n763 VSUBS 0.008559f
C935 B.n764 VSUBS 0.008559f
C936 B.n765 VSUBS 0.008559f
C937 B.n766 VSUBS 0.008559f
C938 B.n767 VSUBS 0.008559f
C939 B.n768 VSUBS 0.008559f
C940 B.n769 VSUBS 0.008559f
C941 B.n770 VSUBS 0.008559f
C942 B.n771 VSUBS 0.008559f
C943 B.n772 VSUBS 0.008055f
C944 B.n773 VSUBS 0.019829f
C945 B.n774 VSUBS 0.004783f
C946 B.n775 VSUBS 0.008559f
C947 B.n776 VSUBS 0.008559f
C948 B.n777 VSUBS 0.008559f
C949 B.n778 VSUBS 0.008559f
C950 B.n779 VSUBS 0.008559f
C951 B.n780 VSUBS 0.008559f
C952 B.n781 VSUBS 0.008559f
C953 B.n782 VSUBS 0.008559f
C954 B.n783 VSUBS 0.008559f
C955 B.n784 VSUBS 0.008559f
C956 B.n785 VSUBS 0.008559f
C957 B.n786 VSUBS 0.008559f
C958 B.n787 VSUBS 0.004783f
C959 B.n788 VSUBS 0.008559f
C960 B.n789 VSUBS 0.008559f
C961 B.n790 VSUBS 0.008559f
C962 B.n791 VSUBS 0.008559f
C963 B.n792 VSUBS 0.008559f
C964 B.n793 VSUBS 0.008559f
C965 B.n794 VSUBS 0.008559f
C966 B.n795 VSUBS 0.008559f
C967 B.n796 VSUBS 0.008559f
C968 B.n797 VSUBS 0.008559f
C969 B.n798 VSUBS 0.008559f
C970 B.n799 VSUBS 0.008559f
C971 B.n800 VSUBS 0.008559f
C972 B.n801 VSUBS 0.008559f
C973 B.n802 VSUBS 0.008559f
C974 B.n803 VSUBS 0.008559f
C975 B.n804 VSUBS 0.008559f
C976 B.n805 VSUBS 0.008559f
C977 B.n806 VSUBS 0.008559f
C978 B.n807 VSUBS 0.008559f
C979 B.n808 VSUBS 0.008559f
C980 B.n809 VSUBS 0.008559f
C981 B.n810 VSUBS 0.008559f
C982 B.n811 VSUBS 0.008559f
C983 B.n812 VSUBS 0.008559f
C984 B.n813 VSUBS 0.008559f
C985 B.n814 VSUBS 0.008559f
C986 B.n815 VSUBS 0.008559f
C987 B.n816 VSUBS 0.008559f
C988 B.n817 VSUBS 0.008559f
C989 B.n818 VSUBS 0.008559f
C990 B.n819 VSUBS 0.008559f
C991 B.n820 VSUBS 0.008559f
C992 B.n821 VSUBS 0.008559f
C993 B.n822 VSUBS 0.008559f
C994 B.n823 VSUBS 0.008559f
C995 B.n824 VSUBS 0.008559f
C996 B.n825 VSUBS 0.008559f
C997 B.n826 VSUBS 0.008559f
C998 B.n827 VSUBS 0.008559f
C999 B.n828 VSUBS 0.008559f
C1000 B.n829 VSUBS 0.008559f
C1001 B.n830 VSUBS 0.008559f
C1002 B.n831 VSUBS 0.008559f
C1003 B.n832 VSUBS 0.008559f
C1004 B.n833 VSUBS 0.008559f
C1005 B.n834 VSUBS 0.008559f
C1006 B.n835 VSUBS 0.008559f
C1007 B.n836 VSUBS 0.008559f
C1008 B.n837 VSUBS 0.008559f
C1009 B.n838 VSUBS 0.008559f
C1010 B.n839 VSUBS 0.008559f
C1011 B.n840 VSUBS 0.008559f
C1012 B.n841 VSUBS 0.008559f
C1013 B.n842 VSUBS 0.008559f
C1014 B.n843 VSUBS 0.008559f
C1015 B.n844 VSUBS 0.008559f
C1016 B.n845 VSUBS 0.008559f
C1017 B.n846 VSUBS 0.008559f
C1018 B.n847 VSUBS 0.008559f
C1019 B.n848 VSUBS 0.008559f
C1020 B.n849 VSUBS 0.008559f
C1021 B.n850 VSUBS 0.008559f
C1022 B.n851 VSUBS 0.008559f
C1023 B.n852 VSUBS 0.008559f
C1024 B.n853 VSUBS 0.008559f
C1025 B.n854 VSUBS 0.008559f
C1026 B.n855 VSUBS 0.008559f
C1027 B.n856 VSUBS 0.008559f
C1028 B.n857 VSUBS 0.008559f
C1029 B.n858 VSUBS 0.008559f
C1030 B.n859 VSUBS 0.008559f
C1031 B.n860 VSUBS 0.008559f
C1032 B.n861 VSUBS 0.021921f
C1033 B.n862 VSUBS 0.020872f
C1034 B.n863 VSUBS 0.020872f
C1035 B.n864 VSUBS 0.008559f
C1036 B.n865 VSUBS 0.008559f
C1037 B.n866 VSUBS 0.008559f
C1038 B.n867 VSUBS 0.008559f
C1039 B.n868 VSUBS 0.008559f
C1040 B.n869 VSUBS 0.008559f
C1041 B.n870 VSUBS 0.008559f
C1042 B.n871 VSUBS 0.008559f
C1043 B.n872 VSUBS 0.008559f
C1044 B.n873 VSUBS 0.008559f
C1045 B.n874 VSUBS 0.008559f
C1046 B.n875 VSUBS 0.008559f
C1047 B.n876 VSUBS 0.008559f
C1048 B.n877 VSUBS 0.008559f
C1049 B.n878 VSUBS 0.008559f
C1050 B.n879 VSUBS 0.008559f
C1051 B.n880 VSUBS 0.008559f
C1052 B.n881 VSUBS 0.008559f
C1053 B.n882 VSUBS 0.008559f
C1054 B.n883 VSUBS 0.008559f
C1055 B.n884 VSUBS 0.008559f
C1056 B.n885 VSUBS 0.008559f
C1057 B.n886 VSUBS 0.008559f
C1058 B.n887 VSUBS 0.008559f
C1059 B.n888 VSUBS 0.008559f
C1060 B.n889 VSUBS 0.008559f
C1061 B.n890 VSUBS 0.008559f
C1062 B.n891 VSUBS 0.008559f
C1063 B.n892 VSUBS 0.008559f
C1064 B.n893 VSUBS 0.008559f
C1065 B.n894 VSUBS 0.008559f
C1066 B.n895 VSUBS 0.008559f
C1067 B.n896 VSUBS 0.008559f
C1068 B.n897 VSUBS 0.008559f
C1069 B.n898 VSUBS 0.008559f
C1070 B.n899 VSUBS 0.008559f
C1071 B.n900 VSUBS 0.008559f
C1072 B.n901 VSUBS 0.008559f
C1073 B.n902 VSUBS 0.008559f
C1074 B.n903 VSUBS 0.008559f
C1075 B.n904 VSUBS 0.008559f
C1076 B.n905 VSUBS 0.008559f
C1077 B.n906 VSUBS 0.008559f
C1078 B.n907 VSUBS 0.008559f
C1079 B.n908 VSUBS 0.008559f
C1080 B.n909 VSUBS 0.008559f
C1081 B.n910 VSUBS 0.008559f
C1082 B.n911 VSUBS 0.008559f
C1083 B.n912 VSUBS 0.008559f
C1084 B.n913 VSUBS 0.008559f
C1085 B.n914 VSUBS 0.008559f
C1086 B.n915 VSUBS 0.008559f
C1087 B.n916 VSUBS 0.008559f
C1088 B.n917 VSUBS 0.008559f
C1089 B.n918 VSUBS 0.008559f
C1090 B.n919 VSUBS 0.008559f
C1091 B.n920 VSUBS 0.008559f
C1092 B.n921 VSUBS 0.008559f
C1093 B.n922 VSUBS 0.008559f
C1094 B.n923 VSUBS 0.008559f
C1095 B.n924 VSUBS 0.008559f
C1096 B.n925 VSUBS 0.008559f
C1097 B.n926 VSUBS 0.008559f
C1098 B.n927 VSUBS 0.008559f
C1099 B.n928 VSUBS 0.008559f
C1100 B.n929 VSUBS 0.008559f
C1101 B.n930 VSUBS 0.008559f
C1102 B.n931 VSUBS 0.008559f
C1103 B.n932 VSUBS 0.008559f
C1104 B.n933 VSUBS 0.008559f
C1105 B.n934 VSUBS 0.008559f
C1106 B.n935 VSUBS 0.008559f
C1107 B.n936 VSUBS 0.008559f
C1108 B.n937 VSUBS 0.008559f
C1109 B.n938 VSUBS 0.008559f
C1110 B.n939 VSUBS 0.008559f
C1111 B.n940 VSUBS 0.008559f
C1112 B.n941 VSUBS 0.008559f
C1113 B.n942 VSUBS 0.008559f
C1114 B.n943 VSUBS 0.008559f
C1115 B.n944 VSUBS 0.008559f
C1116 B.n945 VSUBS 0.008559f
C1117 B.n946 VSUBS 0.008559f
C1118 B.n947 VSUBS 0.008559f
C1119 B.n948 VSUBS 0.008559f
C1120 B.n949 VSUBS 0.008559f
C1121 B.n950 VSUBS 0.008559f
C1122 B.n951 VSUBS 0.008559f
C1123 B.n952 VSUBS 0.008559f
C1124 B.n953 VSUBS 0.008559f
C1125 B.n954 VSUBS 0.008559f
C1126 B.n955 VSUBS 0.008559f
C1127 B.n956 VSUBS 0.008559f
C1128 B.n957 VSUBS 0.008559f
C1129 B.n958 VSUBS 0.008559f
C1130 B.n959 VSUBS 0.01938f
C1131 VDD2.t5 VSUBS 3.58089f
C1132 VDD2.t7 VSUBS 0.338646f
C1133 VDD2.t9 VSUBS 0.338646f
C1134 VDD2.n0 VSUBS 2.72375f
C1135 VDD2.n1 VSUBS 1.80289f
C1136 VDD2.t8 VSUBS 0.338646f
C1137 VDD2.t2 VSUBS 0.338646f
C1138 VDD2.n2 VSUBS 2.75208f
C1139 VDD2.n3 VSUBS 4.07613f
C1140 VDD2.t4 VSUBS 3.5468f
C1141 VDD2.n4 VSUBS 4.36708f
C1142 VDD2.t0 VSUBS 0.338646f
C1143 VDD2.t3 VSUBS 0.338646f
C1144 VDD2.n5 VSUBS 2.72375f
C1145 VDD2.n6 VSUBS 0.902253f
C1146 VDD2.t1 VSUBS 0.338646f
C1147 VDD2.t6 VSUBS 0.338646f
C1148 VDD2.n7 VSUBS 2.75203f
C1149 VTAIL.t14 VSUBS 0.326739f
C1150 VTAIL.t11 VSUBS 0.326739f
C1151 VTAIL.n0 VSUBS 2.45969f
C1152 VTAIL.n1 VSUBS 1.0432f
C1153 VTAIL.t0 VSUBS 3.23178f
C1154 VTAIL.n2 VSUBS 1.21937f
C1155 VTAIL.t9 VSUBS 0.326739f
C1156 VTAIL.t2 VSUBS 0.326739f
C1157 VTAIL.n3 VSUBS 2.45969f
C1158 VTAIL.n4 VSUBS 1.18245f
C1159 VTAIL.t8 VSUBS 0.326739f
C1160 VTAIL.t6 VSUBS 0.326739f
C1161 VTAIL.n5 VSUBS 2.45969f
C1162 VTAIL.n6 VSUBS 2.96497f
C1163 VTAIL.t18 VSUBS 0.326739f
C1164 VTAIL.t13 VSUBS 0.326739f
C1165 VTAIL.n7 VSUBS 2.4597f
C1166 VTAIL.n8 VSUBS 2.96497f
C1167 VTAIL.t17 VSUBS 0.326739f
C1168 VTAIL.t16 VSUBS 0.326739f
C1169 VTAIL.n9 VSUBS 2.4597f
C1170 VTAIL.n10 VSUBS 1.18244f
C1171 VTAIL.t15 VSUBS 3.23179f
C1172 VTAIL.n11 VSUBS 1.21936f
C1173 VTAIL.t7 VSUBS 0.326739f
C1174 VTAIL.t3 VSUBS 0.326739f
C1175 VTAIL.n12 VSUBS 2.4597f
C1176 VTAIL.n13 VSUBS 1.10034f
C1177 VTAIL.t4 VSUBS 0.326739f
C1178 VTAIL.t5 VSUBS 0.326739f
C1179 VTAIL.n14 VSUBS 2.4597f
C1180 VTAIL.n15 VSUBS 1.18244f
C1181 VTAIL.t1 VSUBS 3.23179f
C1182 VTAIL.n16 VSUBS 2.83416f
C1183 VTAIL.t19 VSUBS 3.23178f
C1184 VTAIL.n17 VSUBS 2.83417f
C1185 VTAIL.t10 VSUBS 0.326739f
C1186 VTAIL.t12 VSUBS 0.326739f
C1187 VTAIL.n18 VSUBS 2.45969f
C1188 VTAIL.n19 VSUBS 0.989778f
C1189 VN.n0 VSUBS 0.033367f
C1190 VN.t7 VSUBS 2.8881f
C1191 VN.n1 VSUBS 0.049475f
C1192 VN.n2 VSUBS 0.02531f
C1193 VN.n3 VSUBS 0.027009f
C1194 VN.n4 VSUBS 0.02531f
C1195 VN.n5 VSUBS 0.043033f
C1196 VN.n6 VSUBS 0.02531f
C1197 VN.t0 VSUBS 2.8881f
C1198 VN.n7 VSUBS 0.046936f
C1199 VN.n8 VSUBS 0.02531f
C1200 VN.n9 VSUBS 0.043692f
C1201 VN.t4 VSUBS 3.14354f
C1202 VN.t2 VSUBS 2.8881f
C1203 VN.n10 VSUBS 1.09497f
C1204 VN.n11 VSUBS 1.04678f
C1205 VN.n12 VSUBS 0.266922f
C1206 VN.n13 VSUBS 0.02531f
C1207 VN.n14 VSUBS 0.047374f
C1208 VN.n15 VSUBS 0.030113f
C1209 VN.n16 VSUBS 0.043033f
C1210 VN.n17 VSUBS 0.02531f
C1211 VN.n18 VSUBS 0.02531f
C1212 VN.n19 VSUBS 0.02531f
C1213 VN.n20 VSUBS 0.03535f
C1214 VN.n21 VSUBS 1.00833f
C1215 VN.n22 VSUBS 0.03535f
C1216 VN.n23 VSUBS 0.046936f
C1217 VN.n24 VSUBS 0.02531f
C1218 VN.n25 VSUBS 0.02531f
C1219 VN.n26 VSUBS 0.02531f
C1220 VN.n27 VSUBS 0.030113f
C1221 VN.n28 VSUBS 0.047374f
C1222 VN.t1 VSUBS 2.8881f
C1223 VN.n29 VSUBS 1.00833f
C1224 VN.n30 VSUBS 0.043692f
C1225 VN.n31 VSUBS 0.02531f
C1226 VN.n32 VSUBS 0.02531f
C1227 VN.n33 VSUBS 0.02531f
C1228 VN.n34 VSUBS 0.046936f
C1229 VN.n35 VSUBS 0.050473f
C1230 VN.n36 VSUBS 0.020572f
C1231 VN.n37 VSUBS 0.02531f
C1232 VN.n38 VSUBS 0.02531f
C1233 VN.n39 VSUBS 0.02531f
C1234 VN.n40 VSUBS 0.046936f
C1235 VN.n41 VSUBS 0.028862f
C1236 VN.n42 VSUBS 1.09464f
C1237 VN.n43 VSUBS 0.046232f
C1238 VN.n44 VSUBS 0.033367f
C1239 VN.t5 VSUBS 2.8881f
C1240 VN.n45 VSUBS 0.049475f
C1241 VN.n46 VSUBS 0.02531f
C1242 VN.n47 VSUBS 0.027009f
C1243 VN.n48 VSUBS 0.02531f
C1244 VN.t9 VSUBS 2.8881f
C1245 VN.n49 VSUBS 1.00833f
C1246 VN.n50 VSUBS 0.043033f
C1247 VN.n51 VSUBS 0.02531f
C1248 VN.t6 VSUBS 2.8881f
C1249 VN.n52 VSUBS 0.046936f
C1250 VN.n53 VSUBS 0.02531f
C1251 VN.n54 VSUBS 0.043692f
C1252 VN.t3 VSUBS 3.14354f
C1253 VN.t8 VSUBS 2.8881f
C1254 VN.n55 VSUBS 1.09497f
C1255 VN.n56 VSUBS 1.04678f
C1256 VN.n57 VSUBS 0.266922f
C1257 VN.n58 VSUBS 0.02531f
C1258 VN.n59 VSUBS 0.047374f
C1259 VN.n60 VSUBS 0.030113f
C1260 VN.n61 VSUBS 0.043033f
C1261 VN.n62 VSUBS 0.02531f
C1262 VN.n63 VSUBS 0.02531f
C1263 VN.n64 VSUBS 0.02531f
C1264 VN.n65 VSUBS 0.03535f
C1265 VN.n66 VSUBS 1.00833f
C1266 VN.n67 VSUBS 0.03535f
C1267 VN.n68 VSUBS 0.046936f
C1268 VN.n69 VSUBS 0.02531f
C1269 VN.n70 VSUBS 0.02531f
C1270 VN.n71 VSUBS 0.02531f
C1271 VN.n72 VSUBS 0.030113f
C1272 VN.n73 VSUBS 0.047374f
C1273 VN.n74 VSUBS 0.043692f
C1274 VN.n75 VSUBS 0.02531f
C1275 VN.n76 VSUBS 0.02531f
C1276 VN.n77 VSUBS 0.02531f
C1277 VN.n78 VSUBS 0.046936f
C1278 VN.n79 VSUBS 0.050473f
C1279 VN.n80 VSUBS 0.020572f
C1280 VN.n81 VSUBS 0.02531f
C1281 VN.n82 VSUBS 0.02531f
C1282 VN.n83 VSUBS 0.02531f
C1283 VN.n84 VSUBS 0.046936f
C1284 VN.n85 VSUBS 0.028862f
C1285 VN.n86 VSUBS 1.09464f
C1286 VN.n87 VSUBS 1.69467f
.ends

