* NGSPICE file created from diff_pair_sample_0311.ext - technology: sky130A

.subckt diff_pair_sample_0311 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t3 w_n1606_n3736# sky130_fd_pr__pfet_01v8 ad=5.3976 pd=28.46 as=5.3976 ps=28.46 w=13.84 l=1.26
X1 B.t11 B.t9 B.t10 w_n1606_n3736# sky130_fd_pr__pfet_01v8 ad=5.3976 pd=28.46 as=0 ps=0 w=13.84 l=1.26
X2 B.t8 B.t6 B.t7 w_n1606_n3736# sky130_fd_pr__pfet_01v8 ad=5.3976 pd=28.46 as=0 ps=0 w=13.84 l=1.26
X3 VDD2.t0 VN.t1 VTAIL.t2 w_n1606_n3736# sky130_fd_pr__pfet_01v8 ad=5.3976 pd=28.46 as=5.3976 ps=28.46 w=13.84 l=1.26
X4 VDD1.t1 VP.t0 VTAIL.t0 w_n1606_n3736# sky130_fd_pr__pfet_01v8 ad=5.3976 pd=28.46 as=5.3976 ps=28.46 w=13.84 l=1.26
X5 B.t5 B.t3 B.t4 w_n1606_n3736# sky130_fd_pr__pfet_01v8 ad=5.3976 pd=28.46 as=0 ps=0 w=13.84 l=1.26
X6 VDD1.t0 VP.t1 VTAIL.t1 w_n1606_n3736# sky130_fd_pr__pfet_01v8 ad=5.3976 pd=28.46 as=5.3976 ps=28.46 w=13.84 l=1.26
X7 B.t2 B.t0 B.t1 w_n1606_n3736# sky130_fd_pr__pfet_01v8 ad=5.3976 pd=28.46 as=0 ps=0 w=13.84 l=1.26
R0 VN VN.t1 419.281
R1 VN VN.t0 376.644
R2 VTAIL.n2 VTAIL.t1 56.0655
R3 VTAIL.n1 VTAIL.t2 56.0655
R4 VTAIL.n3 VTAIL.t3 56.0653
R5 VTAIL.n0 VTAIL.t0 56.0653
R6 VTAIL.n1 VTAIL.n0 27.0393
R7 VTAIL.n3 VTAIL.n2 25.6686
R8 VTAIL.n2 VTAIL.n1 1.15567
R9 VTAIL VTAIL.n0 0.87119
R10 VTAIL VTAIL.n3 0.284983
R11 VDD2.n0 VDD2.t1 111.076
R12 VDD2.n0 VDD2.t0 72.7443
R13 VDD2 VDD2.n0 0.401362
R14 B.n330 B.n85 585
R15 B.n329 B.n328 585
R16 B.n327 B.n86 585
R17 B.n326 B.n325 585
R18 B.n324 B.n87 585
R19 B.n323 B.n322 585
R20 B.n321 B.n88 585
R21 B.n320 B.n319 585
R22 B.n318 B.n89 585
R23 B.n317 B.n316 585
R24 B.n315 B.n90 585
R25 B.n314 B.n313 585
R26 B.n312 B.n91 585
R27 B.n311 B.n310 585
R28 B.n309 B.n92 585
R29 B.n308 B.n307 585
R30 B.n306 B.n93 585
R31 B.n305 B.n304 585
R32 B.n303 B.n94 585
R33 B.n302 B.n301 585
R34 B.n300 B.n95 585
R35 B.n299 B.n298 585
R36 B.n297 B.n96 585
R37 B.n296 B.n295 585
R38 B.n294 B.n97 585
R39 B.n293 B.n292 585
R40 B.n291 B.n98 585
R41 B.n290 B.n289 585
R42 B.n288 B.n99 585
R43 B.n287 B.n286 585
R44 B.n285 B.n100 585
R45 B.n284 B.n283 585
R46 B.n282 B.n101 585
R47 B.n281 B.n280 585
R48 B.n279 B.n102 585
R49 B.n278 B.n277 585
R50 B.n276 B.n103 585
R51 B.n275 B.n274 585
R52 B.n273 B.n104 585
R53 B.n272 B.n271 585
R54 B.n270 B.n105 585
R55 B.n269 B.n268 585
R56 B.n267 B.n106 585
R57 B.n266 B.n265 585
R58 B.n264 B.n107 585
R59 B.n263 B.n262 585
R60 B.n261 B.n108 585
R61 B.n260 B.n259 585
R62 B.n255 B.n109 585
R63 B.n254 B.n253 585
R64 B.n252 B.n110 585
R65 B.n251 B.n250 585
R66 B.n249 B.n111 585
R67 B.n248 B.n247 585
R68 B.n246 B.n112 585
R69 B.n245 B.n244 585
R70 B.n243 B.n113 585
R71 B.n241 B.n240 585
R72 B.n239 B.n116 585
R73 B.n238 B.n237 585
R74 B.n236 B.n117 585
R75 B.n235 B.n234 585
R76 B.n233 B.n118 585
R77 B.n232 B.n231 585
R78 B.n230 B.n119 585
R79 B.n229 B.n228 585
R80 B.n227 B.n120 585
R81 B.n226 B.n225 585
R82 B.n224 B.n121 585
R83 B.n223 B.n222 585
R84 B.n221 B.n122 585
R85 B.n220 B.n219 585
R86 B.n218 B.n123 585
R87 B.n217 B.n216 585
R88 B.n215 B.n124 585
R89 B.n214 B.n213 585
R90 B.n212 B.n125 585
R91 B.n211 B.n210 585
R92 B.n209 B.n126 585
R93 B.n208 B.n207 585
R94 B.n206 B.n127 585
R95 B.n205 B.n204 585
R96 B.n203 B.n128 585
R97 B.n202 B.n201 585
R98 B.n200 B.n129 585
R99 B.n199 B.n198 585
R100 B.n197 B.n130 585
R101 B.n196 B.n195 585
R102 B.n194 B.n131 585
R103 B.n193 B.n192 585
R104 B.n191 B.n132 585
R105 B.n190 B.n189 585
R106 B.n188 B.n133 585
R107 B.n187 B.n186 585
R108 B.n185 B.n134 585
R109 B.n184 B.n183 585
R110 B.n182 B.n135 585
R111 B.n181 B.n180 585
R112 B.n179 B.n136 585
R113 B.n178 B.n177 585
R114 B.n176 B.n137 585
R115 B.n175 B.n174 585
R116 B.n173 B.n138 585
R117 B.n172 B.n171 585
R118 B.n332 B.n331 585
R119 B.n333 B.n84 585
R120 B.n335 B.n334 585
R121 B.n336 B.n83 585
R122 B.n338 B.n337 585
R123 B.n339 B.n82 585
R124 B.n341 B.n340 585
R125 B.n342 B.n81 585
R126 B.n344 B.n343 585
R127 B.n345 B.n80 585
R128 B.n347 B.n346 585
R129 B.n348 B.n79 585
R130 B.n350 B.n349 585
R131 B.n351 B.n78 585
R132 B.n353 B.n352 585
R133 B.n354 B.n77 585
R134 B.n356 B.n355 585
R135 B.n357 B.n76 585
R136 B.n359 B.n358 585
R137 B.n360 B.n75 585
R138 B.n362 B.n361 585
R139 B.n363 B.n74 585
R140 B.n365 B.n364 585
R141 B.n366 B.n73 585
R142 B.n368 B.n367 585
R143 B.n369 B.n72 585
R144 B.n371 B.n370 585
R145 B.n372 B.n71 585
R146 B.n374 B.n373 585
R147 B.n375 B.n70 585
R148 B.n377 B.n376 585
R149 B.n378 B.n69 585
R150 B.n380 B.n379 585
R151 B.n381 B.n68 585
R152 B.n383 B.n382 585
R153 B.n384 B.n67 585
R154 B.n542 B.n541 585
R155 B.n540 B.n11 585
R156 B.n539 B.n538 585
R157 B.n537 B.n12 585
R158 B.n536 B.n535 585
R159 B.n534 B.n13 585
R160 B.n533 B.n532 585
R161 B.n531 B.n14 585
R162 B.n530 B.n529 585
R163 B.n528 B.n15 585
R164 B.n527 B.n526 585
R165 B.n525 B.n16 585
R166 B.n524 B.n523 585
R167 B.n522 B.n17 585
R168 B.n521 B.n520 585
R169 B.n519 B.n18 585
R170 B.n518 B.n517 585
R171 B.n516 B.n19 585
R172 B.n515 B.n514 585
R173 B.n513 B.n20 585
R174 B.n512 B.n511 585
R175 B.n510 B.n21 585
R176 B.n509 B.n508 585
R177 B.n507 B.n22 585
R178 B.n506 B.n505 585
R179 B.n504 B.n23 585
R180 B.n503 B.n502 585
R181 B.n501 B.n24 585
R182 B.n500 B.n499 585
R183 B.n498 B.n25 585
R184 B.n497 B.n496 585
R185 B.n495 B.n26 585
R186 B.n494 B.n493 585
R187 B.n492 B.n27 585
R188 B.n491 B.n490 585
R189 B.n489 B.n28 585
R190 B.n488 B.n487 585
R191 B.n486 B.n29 585
R192 B.n485 B.n484 585
R193 B.n483 B.n30 585
R194 B.n482 B.n481 585
R195 B.n480 B.n31 585
R196 B.n479 B.n478 585
R197 B.n477 B.n32 585
R198 B.n476 B.n475 585
R199 B.n474 B.n33 585
R200 B.n473 B.n472 585
R201 B.n471 B.n470 585
R202 B.n469 B.n37 585
R203 B.n468 B.n467 585
R204 B.n466 B.n38 585
R205 B.n465 B.n464 585
R206 B.n463 B.n39 585
R207 B.n462 B.n461 585
R208 B.n460 B.n40 585
R209 B.n459 B.n458 585
R210 B.n457 B.n41 585
R211 B.n455 B.n454 585
R212 B.n453 B.n44 585
R213 B.n452 B.n451 585
R214 B.n450 B.n45 585
R215 B.n449 B.n448 585
R216 B.n447 B.n46 585
R217 B.n446 B.n445 585
R218 B.n444 B.n47 585
R219 B.n443 B.n442 585
R220 B.n441 B.n48 585
R221 B.n440 B.n439 585
R222 B.n438 B.n49 585
R223 B.n437 B.n436 585
R224 B.n435 B.n50 585
R225 B.n434 B.n433 585
R226 B.n432 B.n51 585
R227 B.n431 B.n430 585
R228 B.n429 B.n52 585
R229 B.n428 B.n427 585
R230 B.n426 B.n53 585
R231 B.n425 B.n424 585
R232 B.n423 B.n54 585
R233 B.n422 B.n421 585
R234 B.n420 B.n55 585
R235 B.n419 B.n418 585
R236 B.n417 B.n56 585
R237 B.n416 B.n415 585
R238 B.n414 B.n57 585
R239 B.n413 B.n412 585
R240 B.n411 B.n58 585
R241 B.n410 B.n409 585
R242 B.n408 B.n59 585
R243 B.n407 B.n406 585
R244 B.n405 B.n60 585
R245 B.n404 B.n403 585
R246 B.n402 B.n61 585
R247 B.n401 B.n400 585
R248 B.n399 B.n62 585
R249 B.n398 B.n397 585
R250 B.n396 B.n63 585
R251 B.n395 B.n394 585
R252 B.n393 B.n64 585
R253 B.n392 B.n391 585
R254 B.n390 B.n65 585
R255 B.n389 B.n388 585
R256 B.n387 B.n66 585
R257 B.n386 B.n385 585
R258 B.n543 B.n10 585
R259 B.n545 B.n544 585
R260 B.n546 B.n9 585
R261 B.n548 B.n547 585
R262 B.n549 B.n8 585
R263 B.n551 B.n550 585
R264 B.n552 B.n7 585
R265 B.n554 B.n553 585
R266 B.n555 B.n6 585
R267 B.n557 B.n556 585
R268 B.n558 B.n5 585
R269 B.n560 B.n559 585
R270 B.n561 B.n4 585
R271 B.n563 B.n562 585
R272 B.n564 B.n3 585
R273 B.n566 B.n565 585
R274 B.n567 B.n0 585
R275 B.n2 B.n1 585
R276 B.n148 B.n147 585
R277 B.n149 B.n146 585
R278 B.n151 B.n150 585
R279 B.n152 B.n145 585
R280 B.n154 B.n153 585
R281 B.n155 B.n144 585
R282 B.n157 B.n156 585
R283 B.n158 B.n143 585
R284 B.n160 B.n159 585
R285 B.n161 B.n142 585
R286 B.n163 B.n162 585
R287 B.n164 B.n141 585
R288 B.n166 B.n165 585
R289 B.n167 B.n140 585
R290 B.n169 B.n168 585
R291 B.n170 B.n139 585
R292 B.n114 B.t0 469.137
R293 B.n256 B.t6 469.137
R294 B.n42 B.t3 469.137
R295 B.n34 B.t9 469.137
R296 B.n172 B.n139 463.671
R297 B.n332 B.n85 463.671
R298 B.n386 B.n67 463.671
R299 B.n543 B.n542 463.671
R300 B.n569 B.n568 256.663
R301 B.n568 B.n567 235.042
R302 B.n568 B.n2 235.042
R303 B.n173 B.n172 163.367
R304 B.n174 B.n173 163.367
R305 B.n174 B.n137 163.367
R306 B.n178 B.n137 163.367
R307 B.n179 B.n178 163.367
R308 B.n180 B.n179 163.367
R309 B.n180 B.n135 163.367
R310 B.n184 B.n135 163.367
R311 B.n185 B.n184 163.367
R312 B.n186 B.n185 163.367
R313 B.n186 B.n133 163.367
R314 B.n190 B.n133 163.367
R315 B.n191 B.n190 163.367
R316 B.n192 B.n191 163.367
R317 B.n192 B.n131 163.367
R318 B.n196 B.n131 163.367
R319 B.n197 B.n196 163.367
R320 B.n198 B.n197 163.367
R321 B.n198 B.n129 163.367
R322 B.n202 B.n129 163.367
R323 B.n203 B.n202 163.367
R324 B.n204 B.n203 163.367
R325 B.n204 B.n127 163.367
R326 B.n208 B.n127 163.367
R327 B.n209 B.n208 163.367
R328 B.n210 B.n209 163.367
R329 B.n210 B.n125 163.367
R330 B.n214 B.n125 163.367
R331 B.n215 B.n214 163.367
R332 B.n216 B.n215 163.367
R333 B.n216 B.n123 163.367
R334 B.n220 B.n123 163.367
R335 B.n221 B.n220 163.367
R336 B.n222 B.n221 163.367
R337 B.n222 B.n121 163.367
R338 B.n226 B.n121 163.367
R339 B.n227 B.n226 163.367
R340 B.n228 B.n227 163.367
R341 B.n228 B.n119 163.367
R342 B.n232 B.n119 163.367
R343 B.n233 B.n232 163.367
R344 B.n234 B.n233 163.367
R345 B.n234 B.n117 163.367
R346 B.n238 B.n117 163.367
R347 B.n239 B.n238 163.367
R348 B.n240 B.n239 163.367
R349 B.n240 B.n113 163.367
R350 B.n245 B.n113 163.367
R351 B.n246 B.n245 163.367
R352 B.n247 B.n246 163.367
R353 B.n247 B.n111 163.367
R354 B.n251 B.n111 163.367
R355 B.n252 B.n251 163.367
R356 B.n253 B.n252 163.367
R357 B.n253 B.n109 163.367
R358 B.n260 B.n109 163.367
R359 B.n261 B.n260 163.367
R360 B.n262 B.n261 163.367
R361 B.n262 B.n107 163.367
R362 B.n266 B.n107 163.367
R363 B.n267 B.n266 163.367
R364 B.n268 B.n267 163.367
R365 B.n268 B.n105 163.367
R366 B.n272 B.n105 163.367
R367 B.n273 B.n272 163.367
R368 B.n274 B.n273 163.367
R369 B.n274 B.n103 163.367
R370 B.n278 B.n103 163.367
R371 B.n279 B.n278 163.367
R372 B.n280 B.n279 163.367
R373 B.n280 B.n101 163.367
R374 B.n284 B.n101 163.367
R375 B.n285 B.n284 163.367
R376 B.n286 B.n285 163.367
R377 B.n286 B.n99 163.367
R378 B.n290 B.n99 163.367
R379 B.n291 B.n290 163.367
R380 B.n292 B.n291 163.367
R381 B.n292 B.n97 163.367
R382 B.n296 B.n97 163.367
R383 B.n297 B.n296 163.367
R384 B.n298 B.n297 163.367
R385 B.n298 B.n95 163.367
R386 B.n302 B.n95 163.367
R387 B.n303 B.n302 163.367
R388 B.n304 B.n303 163.367
R389 B.n304 B.n93 163.367
R390 B.n308 B.n93 163.367
R391 B.n309 B.n308 163.367
R392 B.n310 B.n309 163.367
R393 B.n310 B.n91 163.367
R394 B.n314 B.n91 163.367
R395 B.n315 B.n314 163.367
R396 B.n316 B.n315 163.367
R397 B.n316 B.n89 163.367
R398 B.n320 B.n89 163.367
R399 B.n321 B.n320 163.367
R400 B.n322 B.n321 163.367
R401 B.n322 B.n87 163.367
R402 B.n326 B.n87 163.367
R403 B.n327 B.n326 163.367
R404 B.n328 B.n327 163.367
R405 B.n328 B.n85 163.367
R406 B.n382 B.n67 163.367
R407 B.n382 B.n381 163.367
R408 B.n381 B.n380 163.367
R409 B.n380 B.n69 163.367
R410 B.n376 B.n69 163.367
R411 B.n376 B.n375 163.367
R412 B.n375 B.n374 163.367
R413 B.n374 B.n71 163.367
R414 B.n370 B.n71 163.367
R415 B.n370 B.n369 163.367
R416 B.n369 B.n368 163.367
R417 B.n368 B.n73 163.367
R418 B.n364 B.n73 163.367
R419 B.n364 B.n363 163.367
R420 B.n363 B.n362 163.367
R421 B.n362 B.n75 163.367
R422 B.n358 B.n75 163.367
R423 B.n358 B.n357 163.367
R424 B.n357 B.n356 163.367
R425 B.n356 B.n77 163.367
R426 B.n352 B.n77 163.367
R427 B.n352 B.n351 163.367
R428 B.n351 B.n350 163.367
R429 B.n350 B.n79 163.367
R430 B.n346 B.n79 163.367
R431 B.n346 B.n345 163.367
R432 B.n345 B.n344 163.367
R433 B.n344 B.n81 163.367
R434 B.n340 B.n81 163.367
R435 B.n340 B.n339 163.367
R436 B.n339 B.n338 163.367
R437 B.n338 B.n83 163.367
R438 B.n334 B.n83 163.367
R439 B.n334 B.n333 163.367
R440 B.n333 B.n332 163.367
R441 B.n542 B.n11 163.367
R442 B.n538 B.n11 163.367
R443 B.n538 B.n537 163.367
R444 B.n537 B.n536 163.367
R445 B.n536 B.n13 163.367
R446 B.n532 B.n13 163.367
R447 B.n532 B.n531 163.367
R448 B.n531 B.n530 163.367
R449 B.n530 B.n15 163.367
R450 B.n526 B.n15 163.367
R451 B.n526 B.n525 163.367
R452 B.n525 B.n524 163.367
R453 B.n524 B.n17 163.367
R454 B.n520 B.n17 163.367
R455 B.n520 B.n519 163.367
R456 B.n519 B.n518 163.367
R457 B.n518 B.n19 163.367
R458 B.n514 B.n19 163.367
R459 B.n514 B.n513 163.367
R460 B.n513 B.n512 163.367
R461 B.n512 B.n21 163.367
R462 B.n508 B.n21 163.367
R463 B.n508 B.n507 163.367
R464 B.n507 B.n506 163.367
R465 B.n506 B.n23 163.367
R466 B.n502 B.n23 163.367
R467 B.n502 B.n501 163.367
R468 B.n501 B.n500 163.367
R469 B.n500 B.n25 163.367
R470 B.n496 B.n25 163.367
R471 B.n496 B.n495 163.367
R472 B.n495 B.n494 163.367
R473 B.n494 B.n27 163.367
R474 B.n490 B.n27 163.367
R475 B.n490 B.n489 163.367
R476 B.n489 B.n488 163.367
R477 B.n488 B.n29 163.367
R478 B.n484 B.n29 163.367
R479 B.n484 B.n483 163.367
R480 B.n483 B.n482 163.367
R481 B.n482 B.n31 163.367
R482 B.n478 B.n31 163.367
R483 B.n478 B.n477 163.367
R484 B.n477 B.n476 163.367
R485 B.n476 B.n33 163.367
R486 B.n472 B.n33 163.367
R487 B.n472 B.n471 163.367
R488 B.n471 B.n37 163.367
R489 B.n467 B.n37 163.367
R490 B.n467 B.n466 163.367
R491 B.n466 B.n465 163.367
R492 B.n465 B.n39 163.367
R493 B.n461 B.n39 163.367
R494 B.n461 B.n460 163.367
R495 B.n460 B.n459 163.367
R496 B.n459 B.n41 163.367
R497 B.n454 B.n41 163.367
R498 B.n454 B.n453 163.367
R499 B.n453 B.n452 163.367
R500 B.n452 B.n45 163.367
R501 B.n448 B.n45 163.367
R502 B.n448 B.n447 163.367
R503 B.n447 B.n446 163.367
R504 B.n446 B.n47 163.367
R505 B.n442 B.n47 163.367
R506 B.n442 B.n441 163.367
R507 B.n441 B.n440 163.367
R508 B.n440 B.n49 163.367
R509 B.n436 B.n49 163.367
R510 B.n436 B.n435 163.367
R511 B.n435 B.n434 163.367
R512 B.n434 B.n51 163.367
R513 B.n430 B.n51 163.367
R514 B.n430 B.n429 163.367
R515 B.n429 B.n428 163.367
R516 B.n428 B.n53 163.367
R517 B.n424 B.n53 163.367
R518 B.n424 B.n423 163.367
R519 B.n423 B.n422 163.367
R520 B.n422 B.n55 163.367
R521 B.n418 B.n55 163.367
R522 B.n418 B.n417 163.367
R523 B.n417 B.n416 163.367
R524 B.n416 B.n57 163.367
R525 B.n412 B.n57 163.367
R526 B.n412 B.n411 163.367
R527 B.n411 B.n410 163.367
R528 B.n410 B.n59 163.367
R529 B.n406 B.n59 163.367
R530 B.n406 B.n405 163.367
R531 B.n405 B.n404 163.367
R532 B.n404 B.n61 163.367
R533 B.n400 B.n61 163.367
R534 B.n400 B.n399 163.367
R535 B.n399 B.n398 163.367
R536 B.n398 B.n63 163.367
R537 B.n394 B.n63 163.367
R538 B.n394 B.n393 163.367
R539 B.n393 B.n392 163.367
R540 B.n392 B.n65 163.367
R541 B.n388 B.n65 163.367
R542 B.n388 B.n387 163.367
R543 B.n387 B.n386 163.367
R544 B.n544 B.n543 163.367
R545 B.n544 B.n9 163.367
R546 B.n548 B.n9 163.367
R547 B.n549 B.n548 163.367
R548 B.n550 B.n549 163.367
R549 B.n550 B.n7 163.367
R550 B.n554 B.n7 163.367
R551 B.n555 B.n554 163.367
R552 B.n556 B.n555 163.367
R553 B.n556 B.n5 163.367
R554 B.n560 B.n5 163.367
R555 B.n561 B.n560 163.367
R556 B.n562 B.n561 163.367
R557 B.n562 B.n3 163.367
R558 B.n566 B.n3 163.367
R559 B.n567 B.n566 163.367
R560 B.n148 B.n2 163.367
R561 B.n149 B.n148 163.367
R562 B.n150 B.n149 163.367
R563 B.n150 B.n145 163.367
R564 B.n154 B.n145 163.367
R565 B.n155 B.n154 163.367
R566 B.n156 B.n155 163.367
R567 B.n156 B.n143 163.367
R568 B.n160 B.n143 163.367
R569 B.n161 B.n160 163.367
R570 B.n162 B.n161 163.367
R571 B.n162 B.n141 163.367
R572 B.n166 B.n141 163.367
R573 B.n167 B.n166 163.367
R574 B.n168 B.n167 163.367
R575 B.n168 B.n139 163.367
R576 B.n256 B.t7 142.232
R577 B.n42 B.t5 142.232
R578 B.n114 B.t1 142.215
R579 B.n34 B.t11 142.215
R580 B.n257 B.t8 111.397
R581 B.n43 B.t4 111.397
R582 B.n115 B.t2 111.379
R583 B.n35 B.t10 111.379
R584 B.n242 B.n115 59.5399
R585 B.n258 B.n257 59.5399
R586 B.n456 B.n43 59.5399
R587 B.n36 B.n35 59.5399
R588 B.n115 B.n114 30.8369
R589 B.n257 B.n256 30.8369
R590 B.n43 B.n42 30.8369
R591 B.n35 B.n34 30.8369
R592 B.n541 B.n10 30.1273
R593 B.n385 B.n384 30.1273
R594 B.n331 B.n330 30.1273
R595 B.n171 B.n170 30.1273
R596 B B.n569 18.0485
R597 B.n545 B.n10 10.6151
R598 B.n546 B.n545 10.6151
R599 B.n547 B.n546 10.6151
R600 B.n547 B.n8 10.6151
R601 B.n551 B.n8 10.6151
R602 B.n552 B.n551 10.6151
R603 B.n553 B.n552 10.6151
R604 B.n553 B.n6 10.6151
R605 B.n557 B.n6 10.6151
R606 B.n558 B.n557 10.6151
R607 B.n559 B.n558 10.6151
R608 B.n559 B.n4 10.6151
R609 B.n563 B.n4 10.6151
R610 B.n564 B.n563 10.6151
R611 B.n565 B.n564 10.6151
R612 B.n565 B.n0 10.6151
R613 B.n541 B.n540 10.6151
R614 B.n540 B.n539 10.6151
R615 B.n539 B.n12 10.6151
R616 B.n535 B.n12 10.6151
R617 B.n535 B.n534 10.6151
R618 B.n534 B.n533 10.6151
R619 B.n533 B.n14 10.6151
R620 B.n529 B.n14 10.6151
R621 B.n529 B.n528 10.6151
R622 B.n528 B.n527 10.6151
R623 B.n527 B.n16 10.6151
R624 B.n523 B.n16 10.6151
R625 B.n523 B.n522 10.6151
R626 B.n522 B.n521 10.6151
R627 B.n521 B.n18 10.6151
R628 B.n517 B.n18 10.6151
R629 B.n517 B.n516 10.6151
R630 B.n516 B.n515 10.6151
R631 B.n515 B.n20 10.6151
R632 B.n511 B.n20 10.6151
R633 B.n511 B.n510 10.6151
R634 B.n510 B.n509 10.6151
R635 B.n509 B.n22 10.6151
R636 B.n505 B.n22 10.6151
R637 B.n505 B.n504 10.6151
R638 B.n504 B.n503 10.6151
R639 B.n503 B.n24 10.6151
R640 B.n499 B.n24 10.6151
R641 B.n499 B.n498 10.6151
R642 B.n498 B.n497 10.6151
R643 B.n497 B.n26 10.6151
R644 B.n493 B.n26 10.6151
R645 B.n493 B.n492 10.6151
R646 B.n492 B.n491 10.6151
R647 B.n491 B.n28 10.6151
R648 B.n487 B.n28 10.6151
R649 B.n487 B.n486 10.6151
R650 B.n486 B.n485 10.6151
R651 B.n485 B.n30 10.6151
R652 B.n481 B.n30 10.6151
R653 B.n481 B.n480 10.6151
R654 B.n480 B.n479 10.6151
R655 B.n479 B.n32 10.6151
R656 B.n475 B.n32 10.6151
R657 B.n475 B.n474 10.6151
R658 B.n474 B.n473 10.6151
R659 B.n470 B.n469 10.6151
R660 B.n469 B.n468 10.6151
R661 B.n468 B.n38 10.6151
R662 B.n464 B.n38 10.6151
R663 B.n464 B.n463 10.6151
R664 B.n463 B.n462 10.6151
R665 B.n462 B.n40 10.6151
R666 B.n458 B.n40 10.6151
R667 B.n458 B.n457 10.6151
R668 B.n455 B.n44 10.6151
R669 B.n451 B.n44 10.6151
R670 B.n451 B.n450 10.6151
R671 B.n450 B.n449 10.6151
R672 B.n449 B.n46 10.6151
R673 B.n445 B.n46 10.6151
R674 B.n445 B.n444 10.6151
R675 B.n444 B.n443 10.6151
R676 B.n443 B.n48 10.6151
R677 B.n439 B.n48 10.6151
R678 B.n439 B.n438 10.6151
R679 B.n438 B.n437 10.6151
R680 B.n437 B.n50 10.6151
R681 B.n433 B.n50 10.6151
R682 B.n433 B.n432 10.6151
R683 B.n432 B.n431 10.6151
R684 B.n431 B.n52 10.6151
R685 B.n427 B.n52 10.6151
R686 B.n427 B.n426 10.6151
R687 B.n426 B.n425 10.6151
R688 B.n425 B.n54 10.6151
R689 B.n421 B.n54 10.6151
R690 B.n421 B.n420 10.6151
R691 B.n420 B.n419 10.6151
R692 B.n419 B.n56 10.6151
R693 B.n415 B.n56 10.6151
R694 B.n415 B.n414 10.6151
R695 B.n414 B.n413 10.6151
R696 B.n413 B.n58 10.6151
R697 B.n409 B.n58 10.6151
R698 B.n409 B.n408 10.6151
R699 B.n408 B.n407 10.6151
R700 B.n407 B.n60 10.6151
R701 B.n403 B.n60 10.6151
R702 B.n403 B.n402 10.6151
R703 B.n402 B.n401 10.6151
R704 B.n401 B.n62 10.6151
R705 B.n397 B.n62 10.6151
R706 B.n397 B.n396 10.6151
R707 B.n396 B.n395 10.6151
R708 B.n395 B.n64 10.6151
R709 B.n391 B.n64 10.6151
R710 B.n391 B.n390 10.6151
R711 B.n390 B.n389 10.6151
R712 B.n389 B.n66 10.6151
R713 B.n385 B.n66 10.6151
R714 B.n384 B.n383 10.6151
R715 B.n383 B.n68 10.6151
R716 B.n379 B.n68 10.6151
R717 B.n379 B.n378 10.6151
R718 B.n378 B.n377 10.6151
R719 B.n377 B.n70 10.6151
R720 B.n373 B.n70 10.6151
R721 B.n373 B.n372 10.6151
R722 B.n372 B.n371 10.6151
R723 B.n371 B.n72 10.6151
R724 B.n367 B.n72 10.6151
R725 B.n367 B.n366 10.6151
R726 B.n366 B.n365 10.6151
R727 B.n365 B.n74 10.6151
R728 B.n361 B.n74 10.6151
R729 B.n361 B.n360 10.6151
R730 B.n360 B.n359 10.6151
R731 B.n359 B.n76 10.6151
R732 B.n355 B.n76 10.6151
R733 B.n355 B.n354 10.6151
R734 B.n354 B.n353 10.6151
R735 B.n353 B.n78 10.6151
R736 B.n349 B.n78 10.6151
R737 B.n349 B.n348 10.6151
R738 B.n348 B.n347 10.6151
R739 B.n347 B.n80 10.6151
R740 B.n343 B.n80 10.6151
R741 B.n343 B.n342 10.6151
R742 B.n342 B.n341 10.6151
R743 B.n341 B.n82 10.6151
R744 B.n337 B.n82 10.6151
R745 B.n337 B.n336 10.6151
R746 B.n336 B.n335 10.6151
R747 B.n335 B.n84 10.6151
R748 B.n331 B.n84 10.6151
R749 B.n147 B.n1 10.6151
R750 B.n147 B.n146 10.6151
R751 B.n151 B.n146 10.6151
R752 B.n152 B.n151 10.6151
R753 B.n153 B.n152 10.6151
R754 B.n153 B.n144 10.6151
R755 B.n157 B.n144 10.6151
R756 B.n158 B.n157 10.6151
R757 B.n159 B.n158 10.6151
R758 B.n159 B.n142 10.6151
R759 B.n163 B.n142 10.6151
R760 B.n164 B.n163 10.6151
R761 B.n165 B.n164 10.6151
R762 B.n165 B.n140 10.6151
R763 B.n169 B.n140 10.6151
R764 B.n170 B.n169 10.6151
R765 B.n171 B.n138 10.6151
R766 B.n175 B.n138 10.6151
R767 B.n176 B.n175 10.6151
R768 B.n177 B.n176 10.6151
R769 B.n177 B.n136 10.6151
R770 B.n181 B.n136 10.6151
R771 B.n182 B.n181 10.6151
R772 B.n183 B.n182 10.6151
R773 B.n183 B.n134 10.6151
R774 B.n187 B.n134 10.6151
R775 B.n188 B.n187 10.6151
R776 B.n189 B.n188 10.6151
R777 B.n189 B.n132 10.6151
R778 B.n193 B.n132 10.6151
R779 B.n194 B.n193 10.6151
R780 B.n195 B.n194 10.6151
R781 B.n195 B.n130 10.6151
R782 B.n199 B.n130 10.6151
R783 B.n200 B.n199 10.6151
R784 B.n201 B.n200 10.6151
R785 B.n201 B.n128 10.6151
R786 B.n205 B.n128 10.6151
R787 B.n206 B.n205 10.6151
R788 B.n207 B.n206 10.6151
R789 B.n207 B.n126 10.6151
R790 B.n211 B.n126 10.6151
R791 B.n212 B.n211 10.6151
R792 B.n213 B.n212 10.6151
R793 B.n213 B.n124 10.6151
R794 B.n217 B.n124 10.6151
R795 B.n218 B.n217 10.6151
R796 B.n219 B.n218 10.6151
R797 B.n219 B.n122 10.6151
R798 B.n223 B.n122 10.6151
R799 B.n224 B.n223 10.6151
R800 B.n225 B.n224 10.6151
R801 B.n225 B.n120 10.6151
R802 B.n229 B.n120 10.6151
R803 B.n230 B.n229 10.6151
R804 B.n231 B.n230 10.6151
R805 B.n231 B.n118 10.6151
R806 B.n235 B.n118 10.6151
R807 B.n236 B.n235 10.6151
R808 B.n237 B.n236 10.6151
R809 B.n237 B.n116 10.6151
R810 B.n241 B.n116 10.6151
R811 B.n244 B.n243 10.6151
R812 B.n244 B.n112 10.6151
R813 B.n248 B.n112 10.6151
R814 B.n249 B.n248 10.6151
R815 B.n250 B.n249 10.6151
R816 B.n250 B.n110 10.6151
R817 B.n254 B.n110 10.6151
R818 B.n255 B.n254 10.6151
R819 B.n259 B.n255 10.6151
R820 B.n263 B.n108 10.6151
R821 B.n264 B.n263 10.6151
R822 B.n265 B.n264 10.6151
R823 B.n265 B.n106 10.6151
R824 B.n269 B.n106 10.6151
R825 B.n270 B.n269 10.6151
R826 B.n271 B.n270 10.6151
R827 B.n271 B.n104 10.6151
R828 B.n275 B.n104 10.6151
R829 B.n276 B.n275 10.6151
R830 B.n277 B.n276 10.6151
R831 B.n277 B.n102 10.6151
R832 B.n281 B.n102 10.6151
R833 B.n282 B.n281 10.6151
R834 B.n283 B.n282 10.6151
R835 B.n283 B.n100 10.6151
R836 B.n287 B.n100 10.6151
R837 B.n288 B.n287 10.6151
R838 B.n289 B.n288 10.6151
R839 B.n289 B.n98 10.6151
R840 B.n293 B.n98 10.6151
R841 B.n294 B.n293 10.6151
R842 B.n295 B.n294 10.6151
R843 B.n295 B.n96 10.6151
R844 B.n299 B.n96 10.6151
R845 B.n300 B.n299 10.6151
R846 B.n301 B.n300 10.6151
R847 B.n301 B.n94 10.6151
R848 B.n305 B.n94 10.6151
R849 B.n306 B.n305 10.6151
R850 B.n307 B.n306 10.6151
R851 B.n307 B.n92 10.6151
R852 B.n311 B.n92 10.6151
R853 B.n312 B.n311 10.6151
R854 B.n313 B.n312 10.6151
R855 B.n313 B.n90 10.6151
R856 B.n317 B.n90 10.6151
R857 B.n318 B.n317 10.6151
R858 B.n319 B.n318 10.6151
R859 B.n319 B.n88 10.6151
R860 B.n323 B.n88 10.6151
R861 B.n324 B.n323 10.6151
R862 B.n325 B.n324 10.6151
R863 B.n325 B.n86 10.6151
R864 B.n329 B.n86 10.6151
R865 B.n330 B.n329 10.6151
R866 B.n473 B.n36 9.36635
R867 B.n456 B.n455 9.36635
R868 B.n242 B.n241 9.36635
R869 B.n258 B.n108 9.36635
R870 B.n569 B.n0 8.11757
R871 B.n569 B.n1 8.11757
R872 B.n470 B.n36 1.24928
R873 B.n457 B.n456 1.24928
R874 B.n243 B.n242 1.24928
R875 B.n259 B.n258 1.24928
R876 VP.n0 VP.t1 418.995
R877 VP.n0 VP.t0 376.498
R878 VP VP.n0 0.146778
R879 VDD1 VDD1.t1 111.944
R880 VDD1 VDD1.t0 73.1451
C0 VDD1 VTAIL 5.71469f
C1 B VTAIL 3.38652f
C2 B VDD1 1.64929f
C3 VP w_n1606_n3736# 2.33767f
C4 VN w_n1606_n3736# 2.13598f
C5 VDD2 w_n1606_n3736# 1.77461f
C6 VP VN 5.16648f
C7 VP VDD2 0.277531f
C8 VDD2 VN 2.71976f
C9 w_n1606_n3736# VTAIL 3.10263f
C10 VDD1 w_n1606_n3736# 1.76438f
C11 VP VTAIL 2.2259f
C12 VP VDD1 2.84537f
C13 VN VTAIL 2.21138f
C14 VDD1 VN 0.147842f
C15 VDD2 VTAIL 5.75331f
C16 VDD2 VDD1 0.520122f
C17 B w_n1606_n3736# 7.87566f
C18 VP B 1.17358f
C19 B VN 0.847379f
C20 VDD2 B 1.66788f
C21 VDD2 VSUBS 0.846636f
C22 VDD1 VSUBS 4.294515f
C23 VTAIL VSUBS 0.907134f
C24 VN VSUBS 8.003619f
C25 VP VSUBS 1.355626f
C26 B VSUBS 3.060151f
C27 w_n1606_n3736# VSUBS 73.676895f
C28 VDD1.t0 VSUBS 2.28478f
C29 VDD1.t1 VSUBS 2.8735f
C30 VP.t1 VSUBS 3.32332f
C31 VP.t0 VSUBS 2.99564f
C32 VP.n0 VSUBS 6.13141f
C33 B.n0 VSUBS 0.005891f
C34 B.n1 VSUBS 0.005891f
C35 B.n2 VSUBS 0.008712f
C36 B.n3 VSUBS 0.006676f
C37 B.n4 VSUBS 0.006676f
C38 B.n5 VSUBS 0.006676f
C39 B.n6 VSUBS 0.006676f
C40 B.n7 VSUBS 0.006676f
C41 B.n8 VSUBS 0.006676f
C42 B.n9 VSUBS 0.006676f
C43 B.n10 VSUBS 0.014314f
C44 B.n11 VSUBS 0.006676f
C45 B.n12 VSUBS 0.006676f
C46 B.n13 VSUBS 0.006676f
C47 B.n14 VSUBS 0.006676f
C48 B.n15 VSUBS 0.006676f
C49 B.n16 VSUBS 0.006676f
C50 B.n17 VSUBS 0.006676f
C51 B.n18 VSUBS 0.006676f
C52 B.n19 VSUBS 0.006676f
C53 B.n20 VSUBS 0.006676f
C54 B.n21 VSUBS 0.006676f
C55 B.n22 VSUBS 0.006676f
C56 B.n23 VSUBS 0.006676f
C57 B.n24 VSUBS 0.006676f
C58 B.n25 VSUBS 0.006676f
C59 B.n26 VSUBS 0.006676f
C60 B.n27 VSUBS 0.006676f
C61 B.n28 VSUBS 0.006676f
C62 B.n29 VSUBS 0.006676f
C63 B.n30 VSUBS 0.006676f
C64 B.n31 VSUBS 0.006676f
C65 B.n32 VSUBS 0.006676f
C66 B.n33 VSUBS 0.006676f
C67 B.t10 VSUBS 0.436317f
C68 B.t11 VSUBS 0.447974f
C69 B.t9 VSUBS 0.710432f
C70 B.n34 VSUBS 0.184614f
C71 B.n35 VSUBS 0.063282f
C72 B.n36 VSUBS 0.015468f
C73 B.n37 VSUBS 0.006676f
C74 B.n38 VSUBS 0.006676f
C75 B.n39 VSUBS 0.006676f
C76 B.n40 VSUBS 0.006676f
C77 B.n41 VSUBS 0.006676f
C78 B.t4 VSUBS 0.436307f
C79 B.t5 VSUBS 0.447964f
C80 B.t3 VSUBS 0.710432f
C81 B.n42 VSUBS 0.184623f
C82 B.n43 VSUBS 0.063292f
C83 B.n44 VSUBS 0.006676f
C84 B.n45 VSUBS 0.006676f
C85 B.n46 VSUBS 0.006676f
C86 B.n47 VSUBS 0.006676f
C87 B.n48 VSUBS 0.006676f
C88 B.n49 VSUBS 0.006676f
C89 B.n50 VSUBS 0.006676f
C90 B.n51 VSUBS 0.006676f
C91 B.n52 VSUBS 0.006676f
C92 B.n53 VSUBS 0.006676f
C93 B.n54 VSUBS 0.006676f
C94 B.n55 VSUBS 0.006676f
C95 B.n56 VSUBS 0.006676f
C96 B.n57 VSUBS 0.006676f
C97 B.n58 VSUBS 0.006676f
C98 B.n59 VSUBS 0.006676f
C99 B.n60 VSUBS 0.006676f
C100 B.n61 VSUBS 0.006676f
C101 B.n62 VSUBS 0.006676f
C102 B.n63 VSUBS 0.006676f
C103 B.n64 VSUBS 0.006676f
C104 B.n65 VSUBS 0.006676f
C105 B.n66 VSUBS 0.006676f
C106 B.n67 VSUBS 0.014314f
C107 B.n68 VSUBS 0.006676f
C108 B.n69 VSUBS 0.006676f
C109 B.n70 VSUBS 0.006676f
C110 B.n71 VSUBS 0.006676f
C111 B.n72 VSUBS 0.006676f
C112 B.n73 VSUBS 0.006676f
C113 B.n74 VSUBS 0.006676f
C114 B.n75 VSUBS 0.006676f
C115 B.n76 VSUBS 0.006676f
C116 B.n77 VSUBS 0.006676f
C117 B.n78 VSUBS 0.006676f
C118 B.n79 VSUBS 0.006676f
C119 B.n80 VSUBS 0.006676f
C120 B.n81 VSUBS 0.006676f
C121 B.n82 VSUBS 0.006676f
C122 B.n83 VSUBS 0.006676f
C123 B.n84 VSUBS 0.006676f
C124 B.n85 VSUBS 0.015336f
C125 B.n86 VSUBS 0.006676f
C126 B.n87 VSUBS 0.006676f
C127 B.n88 VSUBS 0.006676f
C128 B.n89 VSUBS 0.006676f
C129 B.n90 VSUBS 0.006676f
C130 B.n91 VSUBS 0.006676f
C131 B.n92 VSUBS 0.006676f
C132 B.n93 VSUBS 0.006676f
C133 B.n94 VSUBS 0.006676f
C134 B.n95 VSUBS 0.006676f
C135 B.n96 VSUBS 0.006676f
C136 B.n97 VSUBS 0.006676f
C137 B.n98 VSUBS 0.006676f
C138 B.n99 VSUBS 0.006676f
C139 B.n100 VSUBS 0.006676f
C140 B.n101 VSUBS 0.006676f
C141 B.n102 VSUBS 0.006676f
C142 B.n103 VSUBS 0.006676f
C143 B.n104 VSUBS 0.006676f
C144 B.n105 VSUBS 0.006676f
C145 B.n106 VSUBS 0.006676f
C146 B.n107 VSUBS 0.006676f
C147 B.n108 VSUBS 0.006283f
C148 B.n109 VSUBS 0.006676f
C149 B.n110 VSUBS 0.006676f
C150 B.n111 VSUBS 0.006676f
C151 B.n112 VSUBS 0.006676f
C152 B.n113 VSUBS 0.006676f
C153 B.t2 VSUBS 0.436317f
C154 B.t1 VSUBS 0.447974f
C155 B.t0 VSUBS 0.710432f
C156 B.n114 VSUBS 0.184614f
C157 B.n115 VSUBS 0.063282f
C158 B.n116 VSUBS 0.006676f
C159 B.n117 VSUBS 0.006676f
C160 B.n118 VSUBS 0.006676f
C161 B.n119 VSUBS 0.006676f
C162 B.n120 VSUBS 0.006676f
C163 B.n121 VSUBS 0.006676f
C164 B.n122 VSUBS 0.006676f
C165 B.n123 VSUBS 0.006676f
C166 B.n124 VSUBS 0.006676f
C167 B.n125 VSUBS 0.006676f
C168 B.n126 VSUBS 0.006676f
C169 B.n127 VSUBS 0.006676f
C170 B.n128 VSUBS 0.006676f
C171 B.n129 VSUBS 0.006676f
C172 B.n130 VSUBS 0.006676f
C173 B.n131 VSUBS 0.006676f
C174 B.n132 VSUBS 0.006676f
C175 B.n133 VSUBS 0.006676f
C176 B.n134 VSUBS 0.006676f
C177 B.n135 VSUBS 0.006676f
C178 B.n136 VSUBS 0.006676f
C179 B.n137 VSUBS 0.006676f
C180 B.n138 VSUBS 0.006676f
C181 B.n139 VSUBS 0.014314f
C182 B.n140 VSUBS 0.006676f
C183 B.n141 VSUBS 0.006676f
C184 B.n142 VSUBS 0.006676f
C185 B.n143 VSUBS 0.006676f
C186 B.n144 VSUBS 0.006676f
C187 B.n145 VSUBS 0.006676f
C188 B.n146 VSUBS 0.006676f
C189 B.n147 VSUBS 0.006676f
C190 B.n148 VSUBS 0.006676f
C191 B.n149 VSUBS 0.006676f
C192 B.n150 VSUBS 0.006676f
C193 B.n151 VSUBS 0.006676f
C194 B.n152 VSUBS 0.006676f
C195 B.n153 VSUBS 0.006676f
C196 B.n154 VSUBS 0.006676f
C197 B.n155 VSUBS 0.006676f
C198 B.n156 VSUBS 0.006676f
C199 B.n157 VSUBS 0.006676f
C200 B.n158 VSUBS 0.006676f
C201 B.n159 VSUBS 0.006676f
C202 B.n160 VSUBS 0.006676f
C203 B.n161 VSUBS 0.006676f
C204 B.n162 VSUBS 0.006676f
C205 B.n163 VSUBS 0.006676f
C206 B.n164 VSUBS 0.006676f
C207 B.n165 VSUBS 0.006676f
C208 B.n166 VSUBS 0.006676f
C209 B.n167 VSUBS 0.006676f
C210 B.n168 VSUBS 0.006676f
C211 B.n169 VSUBS 0.006676f
C212 B.n170 VSUBS 0.014314f
C213 B.n171 VSUBS 0.015336f
C214 B.n172 VSUBS 0.015336f
C215 B.n173 VSUBS 0.006676f
C216 B.n174 VSUBS 0.006676f
C217 B.n175 VSUBS 0.006676f
C218 B.n176 VSUBS 0.006676f
C219 B.n177 VSUBS 0.006676f
C220 B.n178 VSUBS 0.006676f
C221 B.n179 VSUBS 0.006676f
C222 B.n180 VSUBS 0.006676f
C223 B.n181 VSUBS 0.006676f
C224 B.n182 VSUBS 0.006676f
C225 B.n183 VSUBS 0.006676f
C226 B.n184 VSUBS 0.006676f
C227 B.n185 VSUBS 0.006676f
C228 B.n186 VSUBS 0.006676f
C229 B.n187 VSUBS 0.006676f
C230 B.n188 VSUBS 0.006676f
C231 B.n189 VSUBS 0.006676f
C232 B.n190 VSUBS 0.006676f
C233 B.n191 VSUBS 0.006676f
C234 B.n192 VSUBS 0.006676f
C235 B.n193 VSUBS 0.006676f
C236 B.n194 VSUBS 0.006676f
C237 B.n195 VSUBS 0.006676f
C238 B.n196 VSUBS 0.006676f
C239 B.n197 VSUBS 0.006676f
C240 B.n198 VSUBS 0.006676f
C241 B.n199 VSUBS 0.006676f
C242 B.n200 VSUBS 0.006676f
C243 B.n201 VSUBS 0.006676f
C244 B.n202 VSUBS 0.006676f
C245 B.n203 VSUBS 0.006676f
C246 B.n204 VSUBS 0.006676f
C247 B.n205 VSUBS 0.006676f
C248 B.n206 VSUBS 0.006676f
C249 B.n207 VSUBS 0.006676f
C250 B.n208 VSUBS 0.006676f
C251 B.n209 VSUBS 0.006676f
C252 B.n210 VSUBS 0.006676f
C253 B.n211 VSUBS 0.006676f
C254 B.n212 VSUBS 0.006676f
C255 B.n213 VSUBS 0.006676f
C256 B.n214 VSUBS 0.006676f
C257 B.n215 VSUBS 0.006676f
C258 B.n216 VSUBS 0.006676f
C259 B.n217 VSUBS 0.006676f
C260 B.n218 VSUBS 0.006676f
C261 B.n219 VSUBS 0.006676f
C262 B.n220 VSUBS 0.006676f
C263 B.n221 VSUBS 0.006676f
C264 B.n222 VSUBS 0.006676f
C265 B.n223 VSUBS 0.006676f
C266 B.n224 VSUBS 0.006676f
C267 B.n225 VSUBS 0.006676f
C268 B.n226 VSUBS 0.006676f
C269 B.n227 VSUBS 0.006676f
C270 B.n228 VSUBS 0.006676f
C271 B.n229 VSUBS 0.006676f
C272 B.n230 VSUBS 0.006676f
C273 B.n231 VSUBS 0.006676f
C274 B.n232 VSUBS 0.006676f
C275 B.n233 VSUBS 0.006676f
C276 B.n234 VSUBS 0.006676f
C277 B.n235 VSUBS 0.006676f
C278 B.n236 VSUBS 0.006676f
C279 B.n237 VSUBS 0.006676f
C280 B.n238 VSUBS 0.006676f
C281 B.n239 VSUBS 0.006676f
C282 B.n240 VSUBS 0.006676f
C283 B.n241 VSUBS 0.006283f
C284 B.n242 VSUBS 0.015468f
C285 B.n243 VSUBS 0.003731f
C286 B.n244 VSUBS 0.006676f
C287 B.n245 VSUBS 0.006676f
C288 B.n246 VSUBS 0.006676f
C289 B.n247 VSUBS 0.006676f
C290 B.n248 VSUBS 0.006676f
C291 B.n249 VSUBS 0.006676f
C292 B.n250 VSUBS 0.006676f
C293 B.n251 VSUBS 0.006676f
C294 B.n252 VSUBS 0.006676f
C295 B.n253 VSUBS 0.006676f
C296 B.n254 VSUBS 0.006676f
C297 B.n255 VSUBS 0.006676f
C298 B.t8 VSUBS 0.436307f
C299 B.t7 VSUBS 0.447964f
C300 B.t6 VSUBS 0.710432f
C301 B.n256 VSUBS 0.184623f
C302 B.n257 VSUBS 0.063292f
C303 B.n258 VSUBS 0.015468f
C304 B.n259 VSUBS 0.003731f
C305 B.n260 VSUBS 0.006676f
C306 B.n261 VSUBS 0.006676f
C307 B.n262 VSUBS 0.006676f
C308 B.n263 VSUBS 0.006676f
C309 B.n264 VSUBS 0.006676f
C310 B.n265 VSUBS 0.006676f
C311 B.n266 VSUBS 0.006676f
C312 B.n267 VSUBS 0.006676f
C313 B.n268 VSUBS 0.006676f
C314 B.n269 VSUBS 0.006676f
C315 B.n270 VSUBS 0.006676f
C316 B.n271 VSUBS 0.006676f
C317 B.n272 VSUBS 0.006676f
C318 B.n273 VSUBS 0.006676f
C319 B.n274 VSUBS 0.006676f
C320 B.n275 VSUBS 0.006676f
C321 B.n276 VSUBS 0.006676f
C322 B.n277 VSUBS 0.006676f
C323 B.n278 VSUBS 0.006676f
C324 B.n279 VSUBS 0.006676f
C325 B.n280 VSUBS 0.006676f
C326 B.n281 VSUBS 0.006676f
C327 B.n282 VSUBS 0.006676f
C328 B.n283 VSUBS 0.006676f
C329 B.n284 VSUBS 0.006676f
C330 B.n285 VSUBS 0.006676f
C331 B.n286 VSUBS 0.006676f
C332 B.n287 VSUBS 0.006676f
C333 B.n288 VSUBS 0.006676f
C334 B.n289 VSUBS 0.006676f
C335 B.n290 VSUBS 0.006676f
C336 B.n291 VSUBS 0.006676f
C337 B.n292 VSUBS 0.006676f
C338 B.n293 VSUBS 0.006676f
C339 B.n294 VSUBS 0.006676f
C340 B.n295 VSUBS 0.006676f
C341 B.n296 VSUBS 0.006676f
C342 B.n297 VSUBS 0.006676f
C343 B.n298 VSUBS 0.006676f
C344 B.n299 VSUBS 0.006676f
C345 B.n300 VSUBS 0.006676f
C346 B.n301 VSUBS 0.006676f
C347 B.n302 VSUBS 0.006676f
C348 B.n303 VSUBS 0.006676f
C349 B.n304 VSUBS 0.006676f
C350 B.n305 VSUBS 0.006676f
C351 B.n306 VSUBS 0.006676f
C352 B.n307 VSUBS 0.006676f
C353 B.n308 VSUBS 0.006676f
C354 B.n309 VSUBS 0.006676f
C355 B.n310 VSUBS 0.006676f
C356 B.n311 VSUBS 0.006676f
C357 B.n312 VSUBS 0.006676f
C358 B.n313 VSUBS 0.006676f
C359 B.n314 VSUBS 0.006676f
C360 B.n315 VSUBS 0.006676f
C361 B.n316 VSUBS 0.006676f
C362 B.n317 VSUBS 0.006676f
C363 B.n318 VSUBS 0.006676f
C364 B.n319 VSUBS 0.006676f
C365 B.n320 VSUBS 0.006676f
C366 B.n321 VSUBS 0.006676f
C367 B.n322 VSUBS 0.006676f
C368 B.n323 VSUBS 0.006676f
C369 B.n324 VSUBS 0.006676f
C370 B.n325 VSUBS 0.006676f
C371 B.n326 VSUBS 0.006676f
C372 B.n327 VSUBS 0.006676f
C373 B.n328 VSUBS 0.006676f
C374 B.n329 VSUBS 0.006676f
C375 B.n330 VSUBS 0.014481f
C376 B.n331 VSUBS 0.015169f
C377 B.n332 VSUBS 0.014314f
C378 B.n333 VSUBS 0.006676f
C379 B.n334 VSUBS 0.006676f
C380 B.n335 VSUBS 0.006676f
C381 B.n336 VSUBS 0.006676f
C382 B.n337 VSUBS 0.006676f
C383 B.n338 VSUBS 0.006676f
C384 B.n339 VSUBS 0.006676f
C385 B.n340 VSUBS 0.006676f
C386 B.n341 VSUBS 0.006676f
C387 B.n342 VSUBS 0.006676f
C388 B.n343 VSUBS 0.006676f
C389 B.n344 VSUBS 0.006676f
C390 B.n345 VSUBS 0.006676f
C391 B.n346 VSUBS 0.006676f
C392 B.n347 VSUBS 0.006676f
C393 B.n348 VSUBS 0.006676f
C394 B.n349 VSUBS 0.006676f
C395 B.n350 VSUBS 0.006676f
C396 B.n351 VSUBS 0.006676f
C397 B.n352 VSUBS 0.006676f
C398 B.n353 VSUBS 0.006676f
C399 B.n354 VSUBS 0.006676f
C400 B.n355 VSUBS 0.006676f
C401 B.n356 VSUBS 0.006676f
C402 B.n357 VSUBS 0.006676f
C403 B.n358 VSUBS 0.006676f
C404 B.n359 VSUBS 0.006676f
C405 B.n360 VSUBS 0.006676f
C406 B.n361 VSUBS 0.006676f
C407 B.n362 VSUBS 0.006676f
C408 B.n363 VSUBS 0.006676f
C409 B.n364 VSUBS 0.006676f
C410 B.n365 VSUBS 0.006676f
C411 B.n366 VSUBS 0.006676f
C412 B.n367 VSUBS 0.006676f
C413 B.n368 VSUBS 0.006676f
C414 B.n369 VSUBS 0.006676f
C415 B.n370 VSUBS 0.006676f
C416 B.n371 VSUBS 0.006676f
C417 B.n372 VSUBS 0.006676f
C418 B.n373 VSUBS 0.006676f
C419 B.n374 VSUBS 0.006676f
C420 B.n375 VSUBS 0.006676f
C421 B.n376 VSUBS 0.006676f
C422 B.n377 VSUBS 0.006676f
C423 B.n378 VSUBS 0.006676f
C424 B.n379 VSUBS 0.006676f
C425 B.n380 VSUBS 0.006676f
C426 B.n381 VSUBS 0.006676f
C427 B.n382 VSUBS 0.006676f
C428 B.n383 VSUBS 0.006676f
C429 B.n384 VSUBS 0.014314f
C430 B.n385 VSUBS 0.015336f
C431 B.n386 VSUBS 0.015336f
C432 B.n387 VSUBS 0.006676f
C433 B.n388 VSUBS 0.006676f
C434 B.n389 VSUBS 0.006676f
C435 B.n390 VSUBS 0.006676f
C436 B.n391 VSUBS 0.006676f
C437 B.n392 VSUBS 0.006676f
C438 B.n393 VSUBS 0.006676f
C439 B.n394 VSUBS 0.006676f
C440 B.n395 VSUBS 0.006676f
C441 B.n396 VSUBS 0.006676f
C442 B.n397 VSUBS 0.006676f
C443 B.n398 VSUBS 0.006676f
C444 B.n399 VSUBS 0.006676f
C445 B.n400 VSUBS 0.006676f
C446 B.n401 VSUBS 0.006676f
C447 B.n402 VSUBS 0.006676f
C448 B.n403 VSUBS 0.006676f
C449 B.n404 VSUBS 0.006676f
C450 B.n405 VSUBS 0.006676f
C451 B.n406 VSUBS 0.006676f
C452 B.n407 VSUBS 0.006676f
C453 B.n408 VSUBS 0.006676f
C454 B.n409 VSUBS 0.006676f
C455 B.n410 VSUBS 0.006676f
C456 B.n411 VSUBS 0.006676f
C457 B.n412 VSUBS 0.006676f
C458 B.n413 VSUBS 0.006676f
C459 B.n414 VSUBS 0.006676f
C460 B.n415 VSUBS 0.006676f
C461 B.n416 VSUBS 0.006676f
C462 B.n417 VSUBS 0.006676f
C463 B.n418 VSUBS 0.006676f
C464 B.n419 VSUBS 0.006676f
C465 B.n420 VSUBS 0.006676f
C466 B.n421 VSUBS 0.006676f
C467 B.n422 VSUBS 0.006676f
C468 B.n423 VSUBS 0.006676f
C469 B.n424 VSUBS 0.006676f
C470 B.n425 VSUBS 0.006676f
C471 B.n426 VSUBS 0.006676f
C472 B.n427 VSUBS 0.006676f
C473 B.n428 VSUBS 0.006676f
C474 B.n429 VSUBS 0.006676f
C475 B.n430 VSUBS 0.006676f
C476 B.n431 VSUBS 0.006676f
C477 B.n432 VSUBS 0.006676f
C478 B.n433 VSUBS 0.006676f
C479 B.n434 VSUBS 0.006676f
C480 B.n435 VSUBS 0.006676f
C481 B.n436 VSUBS 0.006676f
C482 B.n437 VSUBS 0.006676f
C483 B.n438 VSUBS 0.006676f
C484 B.n439 VSUBS 0.006676f
C485 B.n440 VSUBS 0.006676f
C486 B.n441 VSUBS 0.006676f
C487 B.n442 VSUBS 0.006676f
C488 B.n443 VSUBS 0.006676f
C489 B.n444 VSUBS 0.006676f
C490 B.n445 VSUBS 0.006676f
C491 B.n446 VSUBS 0.006676f
C492 B.n447 VSUBS 0.006676f
C493 B.n448 VSUBS 0.006676f
C494 B.n449 VSUBS 0.006676f
C495 B.n450 VSUBS 0.006676f
C496 B.n451 VSUBS 0.006676f
C497 B.n452 VSUBS 0.006676f
C498 B.n453 VSUBS 0.006676f
C499 B.n454 VSUBS 0.006676f
C500 B.n455 VSUBS 0.006283f
C501 B.n456 VSUBS 0.015468f
C502 B.n457 VSUBS 0.003731f
C503 B.n458 VSUBS 0.006676f
C504 B.n459 VSUBS 0.006676f
C505 B.n460 VSUBS 0.006676f
C506 B.n461 VSUBS 0.006676f
C507 B.n462 VSUBS 0.006676f
C508 B.n463 VSUBS 0.006676f
C509 B.n464 VSUBS 0.006676f
C510 B.n465 VSUBS 0.006676f
C511 B.n466 VSUBS 0.006676f
C512 B.n467 VSUBS 0.006676f
C513 B.n468 VSUBS 0.006676f
C514 B.n469 VSUBS 0.006676f
C515 B.n470 VSUBS 0.003731f
C516 B.n471 VSUBS 0.006676f
C517 B.n472 VSUBS 0.006676f
C518 B.n473 VSUBS 0.006283f
C519 B.n474 VSUBS 0.006676f
C520 B.n475 VSUBS 0.006676f
C521 B.n476 VSUBS 0.006676f
C522 B.n477 VSUBS 0.006676f
C523 B.n478 VSUBS 0.006676f
C524 B.n479 VSUBS 0.006676f
C525 B.n480 VSUBS 0.006676f
C526 B.n481 VSUBS 0.006676f
C527 B.n482 VSUBS 0.006676f
C528 B.n483 VSUBS 0.006676f
C529 B.n484 VSUBS 0.006676f
C530 B.n485 VSUBS 0.006676f
C531 B.n486 VSUBS 0.006676f
C532 B.n487 VSUBS 0.006676f
C533 B.n488 VSUBS 0.006676f
C534 B.n489 VSUBS 0.006676f
C535 B.n490 VSUBS 0.006676f
C536 B.n491 VSUBS 0.006676f
C537 B.n492 VSUBS 0.006676f
C538 B.n493 VSUBS 0.006676f
C539 B.n494 VSUBS 0.006676f
C540 B.n495 VSUBS 0.006676f
C541 B.n496 VSUBS 0.006676f
C542 B.n497 VSUBS 0.006676f
C543 B.n498 VSUBS 0.006676f
C544 B.n499 VSUBS 0.006676f
C545 B.n500 VSUBS 0.006676f
C546 B.n501 VSUBS 0.006676f
C547 B.n502 VSUBS 0.006676f
C548 B.n503 VSUBS 0.006676f
C549 B.n504 VSUBS 0.006676f
C550 B.n505 VSUBS 0.006676f
C551 B.n506 VSUBS 0.006676f
C552 B.n507 VSUBS 0.006676f
C553 B.n508 VSUBS 0.006676f
C554 B.n509 VSUBS 0.006676f
C555 B.n510 VSUBS 0.006676f
C556 B.n511 VSUBS 0.006676f
C557 B.n512 VSUBS 0.006676f
C558 B.n513 VSUBS 0.006676f
C559 B.n514 VSUBS 0.006676f
C560 B.n515 VSUBS 0.006676f
C561 B.n516 VSUBS 0.006676f
C562 B.n517 VSUBS 0.006676f
C563 B.n518 VSUBS 0.006676f
C564 B.n519 VSUBS 0.006676f
C565 B.n520 VSUBS 0.006676f
C566 B.n521 VSUBS 0.006676f
C567 B.n522 VSUBS 0.006676f
C568 B.n523 VSUBS 0.006676f
C569 B.n524 VSUBS 0.006676f
C570 B.n525 VSUBS 0.006676f
C571 B.n526 VSUBS 0.006676f
C572 B.n527 VSUBS 0.006676f
C573 B.n528 VSUBS 0.006676f
C574 B.n529 VSUBS 0.006676f
C575 B.n530 VSUBS 0.006676f
C576 B.n531 VSUBS 0.006676f
C577 B.n532 VSUBS 0.006676f
C578 B.n533 VSUBS 0.006676f
C579 B.n534 VSUBS 0.006676f
C580 B.n535 VSUBS 0.006676f
C581 B.n536 VSUBS 0.006676f
C582 B.n537 VSUBS 0.006676f
C583 B.n538 VSUBS 0.006676f
C584 B.n539 VSUBS 0.006676f
C585 B.n540 VSUBS 0.006676f
C586 B.n541 VSUBS 0.015336f
C587 B.n542 VSUBS 0.015336f
C588 B.n543 VSUBS 0.014314f
C589 B.n544 VSUBS 0.006676f
C590 B.n545 VSUBS 0.006676f
C591 B.n546 VSUBS 0.006676f
C592 B.n547 VSUBS 0.006676f
C593 B.n548 VSUBS 0.006676f
C594 B.n549 VSUBS 0.006676f
C595 B.n550 VSUBS 0.006676f
C596 B.n551 VSUBS 0.006676f
C597 B.n552 VSUBS 0.006676f
C598 B.n553 VSUBS 0.006676f
C599 B.n554 VSUBS 0.006676f
C600 B.n555 VSUBS 0.006676f
C601 B.n556 VSUBS 0.006676f
C602 B.n557 VSUBS 0.006676f
C603 B.n558 VSUBS 0.006676f
C604 B.n559 VSUBS 0.006676f
C605 B.n560 VSUBS 0.006676f
C606 B.n561 VSUBS 0.006676f
C607 B.n562 VSUBS 0.006676f
C608 B.n563 VSUBS 0.006676f
C609 B.n564 VSUBS 0.006676f
C610 B.n565 VSUBS 0.006676f
C611 B.n566 VSUBS 0.006676f
C612 B.n567 VSUBS 0.008712f
C613 B.n568 VSUBS 0.009281f
C614 B.n569 VSUBS 0.018455f
C615 VDD2.t1 VSUBS 2.87088f
C616 VDD2.t0 VSUBS 2.30218f
C617 VDD2.n0 VSUBS 3.25536f
C618 VTAIL.t0 VSUBS 3.02553f
C619 VTAIL.n0 VSUBS 2.6111f
C620 VTAIL.t2 VSUBS 3.02555f
C621 VTAIL.n1 VSUBS 2.63708f
C622 VTAIL.t1 VSUBS 3.02555f
C623 VTAIL.n2 VSUBS 2.51182f
C624 VTAIL.t3 VSUBS 3.02553f
C625 VTAIL.n3 VSUBS 2.43227f
C626 VN.t0 VSUBS 2.90586f
C627 VN.t1 VSUBS 3.22834f
.ends

