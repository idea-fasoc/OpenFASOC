* NGSPICE file created from diff_pair_sample_0261.ext - technology: sky130A

.subckt diff_pair_sample_0261 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t14 VP.t0 VDD1.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=2.99145 pd=18.46 as=2.99145 ps=18.46 w=18.13 l=3.62
X1 VDD2.t7 VN.t0 VTAIL.t15 B.t21 sky130_fd_pr__nfet_01v8 ad=2.99145 pd=18.46 as=7.0707 ps=37.04 w=18.13 l=3.62
X2 VTAIL.t2 VN.t1 VDD2.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=7.0707 pd=37.04 as=2.99145 ps=18.46 w=18.13 l=3.62
X3 B.t20 B.t18 B.t19 B.t15 sky130_fd_pr__nfet_01v8 ad=7.0707 pd=37.04 as=0 ps=0 w=18.13 l=3.62
X4 VDD2.t5 VN.t2 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.99145 pd=18.46 as=2.99145 ps=18.46 w=18.13 l=3.62
X5 VTAIL.t13 VP.t1 VDD1.t4 B.t5 sky130_fd_pr__nfet_01v8 ad=2.99145 pd=18.46 as=2.99145 ps=18.46 w=18.13 l=3.62
X6 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=7.0707 pd=37.04 as=0 ps=0 w=18.13 l=3.62
X7 B.t13 B.t11 B.t12 B.t8 sky130_fd_pr__nfet_01v8 ad=7.0707 pd=37.04 as=0 ps=0 w=18.13 l=3.62
X8 VDD1.t3 VP.t2 VTAIL.t12 B.t0 sky130_fd_pr__nfet_01v8 ad=2.99145 pd=18.46 as=2.99145 ps=18.46 w=18.13 l=3.62
X9 VDD2.t4 VN.t3 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.99145 pd=18.46 as=2.99145 ps=18.46 w=18.13 l=3.62
X10 VTAIL.t5 VN.t4 VDD2.t3 B.t5 sky130_fd_pr__nfet_01v8 ad=2.99145 pd=18.46 as=2.99145 ps=18.46 w=18.13 l=3.62
X11 VDD1.t7 VP.t3 VTAIL.t11 B.t1 sky130_fd_pr__nfet_01v8 ad=2.99145 pd=18.46 as=2.99145 ps=18.46 w=18.13 l=3.62
X12 VTAIL.t10 VP.t4 VDD1.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=7.0707 pd=37.04 as=2.99145 ps=18.46 w=18.13 l=3.62
X13 VTAIL.t4 VN.t5 VDD2.t2 B.t4 sky130_fd_pr__nfet_01v8 ad=2.99145 pd=18.46 as=2.99145 ps=18.46 w=18.13 l=3.62
X14 VDD1.t2 VP.t5 VTAIL.t9 B.t21 sky130_fd_pr__nfet_01v8 ad=2.99145 pd=18.46 as=7.0707 ps=37.04 w=18.13 l=3.62
X15 VDD2.t1 VN.t6 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=2.99145 pd=18.46 as=7.0707 ps=37.04 w=18.13 l=3.62
X16 VTAIL.t3 VN.t7 VDD2.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=7.0707 pd=37.04 as=2.99145 ps=18.46 w=18.13 l=3.62
X17 VDD1.t1 VP.t6 VTAIL.t8 B.t6 sky130_fd_pr__nfet_01v8 ad=2.99145 pd=18.46 as=7.0707 ps=37.04 w=18.13 l=3.62
X18 B.t10 B.t7 B.t9 B.t8 sky130_fd_pr__nfet_01v8 ad=7.0707 pd=37.04 as=0 ps=0 w=18.13 l=3.62
X19 VTAIL.t7 VP.t7 VDD1.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=7.0707 pd=37.04 as=2.99145 ps=18.46 w=18.13 l=3.62
R0 VP.n24 VP.n21 161.3
R1 VP.n26 VP.n25 161.3
R2 VP.n27 VP.n20 161.3
R3 VP.n29 VP.n28 161.3
R4 VP.n30 VP.n19 161.3
R5 VP.n32 VP.n31 161.3
R6 VP.n33 VP.n18 161.3
R7 VP.n36 VP.n35 161.3
R8 VP.n37 VP.n17 161.3
R9 VP.n39 VP.n38 161.3
R10 VP.n40 VP.n16 161.3
R11 VP.n42 VP.n41 161.3
R12 VP.n43 VP.n15 161.3
R13 VP.n45 VP.n44 161.3
R14 VP.n46 VP.n14 161.3
R15 VP.n48 VP.n47 161.3
R16 VP.n89 VP.n88 161.3
R17 VP.n87 VP.n1 161.3
R18 VP.n86 VP.n85 161.3
R19 VP.n84 VP.n2 161.3
R20 VP.n83 VP.n82 161.3
R21 VP.n81 VP.n3 161.3
R22 VP.n80 VP.n79 161.3
R23 VP.n78 VP.n4 161.3
R24 VP.n77 VP.n76 161.3
R25 VP.n74 VP.n5 161.3
R26 VP.n73 VP.n72 161.3
R27 VP.n71 VP.n6 161.3
R28 VP.n70 VP.n69 161.3
R29 VP.n68 VP.n7 161.3
R30 VP.n67 VP.n66 161.3
R31 VP.n65 VP.n8 161.3
R32 VP.n64 VP.n63 161.3
R33 VP.n61 VP.n9 161.3
R34 VP.n60 VP.n59 161.3
R35 VP.n58 VP.n10 161.3
R36 VP.n57 VP.n56 161.3
R37 VP.n55 VP.n11 161.3
R38 VP.n54 VP.n53 161.3
R39 VP.n52 VP.n12 161.3
R40 VP.n23 VP.t4 153.856
R41 VP.n50 VP.t7 120.701
R42 VP.n62 VP.t3 120.701
R43 VP.n75 VP.t1 120.701
R44 VP.n0 VP.t6 120.701
R45 VP.n13 VP.t5 120.701
R46 VP.n34 VP.t0 120.701
R47 VP.n22 VP.t2 120.701
R48 VP.n51 VP.n50 81.504
R49 VP.n90 VP.n0 81.504
R50 VP.n49 VP.n13 81.504
R51 VP.n23 VP.n22 63.5476
R52 VP.n51 VP.n49 60.4084
R53 VP.n56 VP.n10 56.5193
R54 VP.n69 VP.n6 56.5193
R55 VP.n82 VP.n2 56.5193
R56 VP.n41 VP.n15 56.5193
R57 VP.n28 VP.n19 56.5193
R58 VP.n54 VP.n12 24.4675
R59 VP.n55 VP.n54 24.4675
R60 VP.n56 VP.n55 24.4675
R61 VP.n60 VP.n10 24.4675
R62 VP.n61 VP.n60 24.4675
R63 VP.n63 VP.n61 24.4675
R64 VP.n67 VP.n8 24.4675
R65 VP.n68 VP.n67 24.4675
R66 VP.n69 VP.n68 24.4675
R67 VP.n73 VP.n6 24.4675
R68 VP.n74 VP.n73 24.4675
R69 VP.n76 VP.n74 24.4675
R70 VP.n80 VP.n4 24.4675
R71 VP.n81 VP.n80 24.4675
R72 VP.n82 VP.n81 24.4675
R73 VP.n86 VP.n2 24.4675
R74 VP.n87 VP.n86 24.4675
R75 VP.n88 VP.n87 24.4675
R76 VP.n45 VP.n15 24.4675
R77 VP.n46 VP.n45 24.4675
R78 VP.n47 VP.n46 24.4675
R79 VP.n32 VP.n19 24.4675
R80 VP.n33 VP.n32 24.4675
R81 VP.n35 VP.n33 24.4675
R82 VP.n39 VP.n17 24.4675
R83 VP.n40 VP.n39 24.4675
R84 VP.n41 VP.n40 24.4675
R85 VP.n26 VP.n21 24.4675
R86 VP.n27 VP.n26 24.4675
R87 VP.n28 VP.n27 24.4675
R88 VP.n63 VP.n62 13.4574
R89 VP.n75 VP.n4 13.4574
R90 VP.n34 VP.n17 13.4574
R91 VP.n62 VP.n8 11.0107
R92 VP.n76 VP.n75 11.0107
R93 VP.n35 VP.n34 11.0107
R94 VP.n22 VP.n21 11.0107
R95 VP.n50 VP.n12 8.56395
R96 VP.n88 VP.n0 8.56395
R97 VP.n47 VP.n13 8.56395
R98 VP.n24 VP.n23 3.20385
R99 VP.n49 VP.n48 0.354971
R100 VP.n52 VP.n51 0.354971
R101 VP.n90 VP.n89 0.354971
R102 VP VP.n90 0.26696
R103 VP.n25 VP.n24 0.189894
R104 VP.n25 VP.n20 0.189894
R105 VP.n29 VP.n20 0.189894
R106 VP.n30 VP.n29 0.189894
R107 VP.n31 VP.n30 0.189894
R108 VP.n31 VP.n18 0.189894
R109 VP.n36 VP.n18 0.189894
R110 VP.n37 VP.n36 0.189894
R111 VP.n38 VP.n37 0.189894
R112 VP.n38 VP.n16 0.189894
R113 VP.n42 VP.n16 0.189894
R114 VP.n43 VP.n42 0.189894
R115 VP.n44 VP.n43 0.189894
R116 VP.n44 VP.n14 0.189894
R117 VP.n48 VP.n14 0.189894
R118 VP.n53 VP.n52 0.189894
R119 VP.n53 VP.n11 0.189894
R120 VP.n57 VP.n11 0.189894
R121 VP.n58 VP.n57 0.189894
R122 VP.n59 VP.n58 0.189894
R123 VP.n59 VP.n9 0.189894
R124 VP.n64 VP.n9 0.189894
R125 VP.n65 VP.n64 0.189894
R126 VP.n66 VP.n65 0.189894
R127 VP.n66 VP.n7 0.189894
R128 VP.n70 VP.n7 0.189894
R129 VP.n71 VP.n70 0.189894
R130 VP.n72 VP.n71 0.189894
R131 VP.n72 VP.n5 0.189894
R132 VP.n77 VP.n5 0.189894
R133 VP.n78 VP.n77 0.189894
R134 VP.n79 VP.n78 0.189894
R135 VP.n79 VP.n3 0.189894
R136 VP.n83 VP.n3 0.189894
R137 VP.n84 VP.n83 0.189894
R138 VP.n85 VP.n84 0.189894
R139 VP.n85 VP.n1 0.189894
R140 VP.n89 VP.n1 0.189894
R141 VDD1 VDD1.n0 60.2757
R142 VDD1.n3 VDD1.n2 60.162
R143 VDD1.n3 VDD1.n1 60.162
R144 VDD1.n5 VDD1.n4 58.5148
R145 VDD1.n5 VDD1.n3 55.2509
R146 VDD1 VDD1.n5 1.6449
R147 VDD1.n4 VDD1.t5 1.09261
R148 VDD1.n4 VDD1.t2 1.09261
R149 VDD1.n0 VDD1.t6 1.09261
R150 VDD1.n0 VDD1.t3 1.09261
R151 VDD1.n2 VDD1.t4 1.09261
R152 VDD1.n2 VDD1.t1 1.09261
R153 VDD1.n1 VDD1.t0 1.09261
R154 VDD1.n1 VDD1.t7 1.09261
R155 VTAIL.n818 VTAIL.n722 289.615
R156 VTAIL.n98 VTAIL.n2 289.615
R157 VTAIL.n200 VTAIL.n104 289.615
R158 VTAIL.n304 VTAIL.n208 289.615
R159 VTAIL.n716 VTAIL.n620 289.615
R160 VTAIL.n612 VTAIL.n516 289.615
R161 VTAIL.n510 VTAIL.n414 289.615
R162 VTAIL.n406 VTAIL.n310 289.615
R163 VTAIL.n754 VTAIL.n753 185
R164 VTAIL.n759 VTAIL.n758 185
R165 VTAIL.n761 VTAIL.n760 185
R166 VTAIL.n750 VTAIL.n749 185
R167 VTAIL.n767 VTAIL.n766 185
R168 VTAIL.n769 VTAIL.n768 185
R169 VTAIL.n746 VTAIL.n745 185
R170 VTAIL.n775 VTAIL.n774 185
R171 VTAIL.n777 VTAIL.n776 185
R172 VTAIL.n742 VTAIL.n741 185
R173 VTAIL.n783 VTAIL.n782 185
R174 VTAIL.n785 VTAIL.n784 185
R175 VTAIL.n738 VTAIL.n737 185
R176 VTAIL.n791 VTAIL.n790 185
R177 VTAIL.n793 VTAIL.n792 185
R178 VTAIL.n734 VTAIL.n733 185
R179 VTAIL.n800 VTAIL.n799 185
R180 VTAIL.n801 VTAIL.n732 185
R181 VTAIL.n803 VTAIL.n802 185
R182 VTAIL.n730 VTAIL.n729 185
R183 VTAIL.n809 VTAIL.n808 185
R184 VTAIL.n811 VTAIL.n810 185
R185 VTAIL.n726 VTAIL.n725 185
R186 VTAIL.n817 VTAIL.n816 185
R187 VTAIL.n819 VTAIL.n818 185
R188 VTAIL.n34 VTAIL.n33 185
R189 VTAIL.n39 VTAIL.n38 185
R190 VTAIL.n41 VTAIL.n40 185
R191 VTAIL.n30 VTAIL.n29 185
R192 VTAIL.n47 VTAIL.n46 185
R193 VTAIL.n49 VTAIL.n48 185
R194 VTAIL.n26 VTAIL.n25 185
R195 VTAIL.n55 VTAIL.n54 185
R196 VTAIL.n57 VTAIL.n56 185
R197 VTAIL.n22 VTAIL.n21 185
R198 VTAIL.n63 VTAIL.n62 185
R199 VTAIL.n65 VTAIL.n64 185
R200 VTAIL.n18 VTAIL.n17 185
R201 VTAIL.n71 VTAIL.n70 185
R202 VTAIL.n73 VTAIL.n72 185
R203 VTAIL.n14 VTAIL.n13 185
R204 VTAIL.n80 VTAIL.n79 185
R205 VTAIL.n81 VTAIL.n12 185
R206 VTAIL.n83 VTAIL.n82 185
R207 VTAIL.n10 VTAIL.n9 185
R208 VTAIL.n89 VTAIL.n88 185
R209 VTAIL.n91 VTAIL.n90 185
R210 VTAIL.n6 VTAIL.n5 185
R211 VTAIL.n97 VTAIL.n96 185
R212 VTAIL.n99 VTAIL.n98 185
R213 VTAIL.n136 VTAIL.n135 185
R214 VTAIL.n141 VTAIL.n140 185
R215 VTAIL.n143 VTAIL.n142 185
R216 VTAIL.n132 VTAIL.n131 185
R217 VTAIL.n149 VTAIL.n148 185
R218 VTAIL.n151 VTAIL.n150 185
R219 VTAIL.n128 VTAIL.n127 185
R220 VTAIL.n157 VTAIL.n156 185
R221 VTAIL.n159 VTAIL.n158 185
R222 VTAIL.n124 VTAIL.n123 185
R223 VTAIL.n165 VTAIL.n164 185
R224 VTAIL.n167 VTAIL.n166 185
R225 VTAIL.n120 VTAIL.n119 185
R226 VTAIL.n173 VTAIL.n172 185
R227 VTAIL.n175 VTAIL.n174 185
R228 VTAIL.n116 VTAIL.n115 185
R229 VTAIL.n182 VTAIL.n181 185
R230 VTAIL.n183 VTAIL.n114 185
R231 VTAIL.n185 VTAIL.n184 185
R232 VTAIL.n112 VTAIL.n111 185
R233 VTAIL.n191 VTAIL.n190 185
R234 VTAIL.n193 VTAIL.n192 185
R235 VTAIL.n108 VTAIL.n107 185
R236 VTAIL.n199 VTAIL.n198 185
R237 VTAIL.n201 VTAIL.n200 185
R238 VTAIL.n240 VTAIL.n239 185
R239 VTAIL.n245 VTAIL.n244 185
R240 VTAIL.n247 VTAIL.n246 185
R241 VTAIL.n236 VTAIL.n235 185
R242 VTAIL.n253 VTAIL.n252 185
R243 VTAIL.n255 VTAIL.n254 185
R244 VTAIL.n232 VTAIL.n231 185
R245 VTAIL.n261 VTAIL.n260 185
R246 VTAIL.n263 VTAIL.n262 185
R247 VTAIL.n228 VTAIL.n227 185
R248 VTAIL.n269 VTAIL.n268 185
R249 VTAIL.n271 VTAIL.n270 185
R250 VTAIL.n224 VTAIL.n223 185
R251 VTAIL.n277 VTAIL.n276 185
R252 VTAIL.n279 VTAIL.n278 185
R253 VTAIL.n220 VTAIL.n219 185
R254 VTAIL.n286 VTAIL.n285 185
R255 VTAIL.n287 VTAIL.n218 185
R256 VTAIL.n289 VTAIL.n288 185
R257 VTAIL.n216 VTAIL.n215 185
R258 VTAIL.n295 VTAIL.n294 185
R259 VTAIL.n297 VTAIL.n296 185
R260 VTAIL.n212 VTAIL.n211 185
R261 VTAIL.n303 VTAIL.n302 185
R262 VTAIL.n305 VTAIL.n304 185
R263 VTAIL.n717 VTAIL.n716 185
R264 VTAIL.n715 VTAIL.n714 185
R265 VTAIL.n624 VTAIL.n623 185
R266 VTAIL.n709 VTAIL.n708 185
R267 VTAIL.n707 VTAIL.n706 185
R268 VTAIL.n628 VTAIL.n627 185
R269 VTAIL.n701 VTAIL.n700 185
R270 VTAIL.n699 VTAIL.n630 185
R271 VTAIL.n698 VTAIL.n697 185
R272 VTAIL.n633 VTAIL.n631 185
R273 VTAIL.n692 VTAIL.n691 185
R274 VTAIL.n690 VTAIL.n689 185
R275 VTAIL.n637 VTAIL.n636 185
R276 VTAIL.n684 VTAIL.n683 185
R277 VTAIL.n682 VTAIL.n681 185
R278 VTAIL.n641 VTAIL.n640 185
R279 VTAIL.n676 VTAIL.n675 185
R280 VTAIL.n674 VTAIL.n673 185
R281 VTAIL.n645 VTAIL.n644 185
R282 VTAIL.n668 VTAIL.n667 185
R283 VTAIL.n666 VTAIL.n665 185
R284 VTAIL.n649 VTAIL.n648 185
R285 VTAIL.n660 VTAIL.n659 185
R286 VTAIL.n658 VTAIL.n657 185
R287 VTAIL.n653 VTAIL.n652 185
R288 VTAIL.n613 VTAIL.n612 185
R289 VTAIL.n611 VTAIL.n610 185
R290 VTAIL.n520 VTAIL.n519 185
R291 VTAIL.n605 VTAIL.n604 185
R292 VTAIL.n603 VTAIL.n602 185
R293 VTAIL.n524 VTAIL.n523 185
R294 VTAIL.n597 VTAIL.n596 185
R295 VTAIL.n595 VTAIL.n526 185
R296 VTAIL.n594 VTAIL.n593 185
R297 VTAIL.n529 VTAIL.n527 185
R298 VTAIL.n588 VTAIL.n587 185
R299 VTAIL.n586 VTAIL.n585 185
R300 VTAIL.n533 VTAIL.n532 185
R301 VTAIL.n580 VTAIL.n579 185
R302 VTAIL.n578 VTAIL.n577 185
R303 VTAIL.n537 VTAIL.n536 185
R304 VTAIL.n572 VTAIL.n571 185
R305 VTAIL.n570 VTAIL.n569 185
R306 VTAIL.n541 VTAIL.n540 185
R307 VTAIL.n564 VTAIL.n563 185
R308 VTAIL.n562 VTAIL.n561 185
R309 VTAIL.n545 VTAIL.n544 185
R310 VTAIL.n556 VTAIL.n555 185
R311 VTAIL.n554 VTAIL.n553 185
R312 VTAIL.n549 VTAIL.n548 185
R313 VTAIL.n511 VTAIL.n510 185
R314 VTAIL.n509 VTAIL.n508 185
R315 VTAIL.n418 VTAIL.n417 185
R316 VTAIL.n503 VTAIL.n502 185
R317 VTAIL.n501 VTAIL.n500 185
R318 VTAIL.n422 VTAIL.n421 185
R319 VTAIL.n495 VTAIL.n494 185
R320 VTAIL.n493 VTAIL.n424 185
R321 VTAIL.n492 VTAIL.n491 185
R322 VTAIL.n427 VTAIL.n425 185
R323 VTAIL.n486 VTAIL.n485 185
R324 VTAIL.n484 VTAIL.n483 185
R325 VTAIL.n431 VTAIL.n430 185
R326 VTAIL.n478 VTAIL.n477 185
R327 VTAIL.n476 VTAIL.n475 185
R328 VTAIL.n435 VTAIL.n434 185
R329 VTAIL.n470 VTAIL.n469 185
R330 VTAIL.n468 VTAIL.n467 185
R331 VTAIL.n439 VTAIL.n438 185
R332 VTAIL.n462 VTAIL.n461 185
R333 VTAIL.n460 VTAIL.n459 185
R334 VTAIL.n443 VTAIL.n442 185
R335 VTAIL.n454 VTAIL.n453 185
R336 VTAIL.n452 VTAIL.n451 185
R337 VTAIL.n447 VTAIL.n446 185
R338 VTAIL.n407 VTAIL.n406 185
R339 VTAIL.n405 VTAIL.n404 185
R340 VTAIL.n314 VTAIL.n313 185
R341 VTAIL.n399 VTAIL.n398 185
R342 VTAIL.n397 VTAIL.n396 185
R343 VTAIL.n318 VTAIL.n317 185
R344 VTAIL.n391 VTAIL.n390 185
R345 VTAIL.n389 VTAIL.n320 185
R346 VTAIL.n388 VTAIL.n387 185
R347 VTAIL.n323 VTAIL.n321 185
R348 VTAIL.n382 VTAIL.n381 185
R349 VTAIL.n380 VTAIL.n379 185
R350 VTAIL.n327 VTAIL.n326 185
R351 VTAIL.n374 VTAIL.n373 185
R352 VTAIL.n372 VTAIL.n371 185
R353 VTAIL.n331 VTAIL.n330 185
R354 VTAIL.n366 VTAIL.n365 185
R355 VTAIL.n364 VTAIL.n363 185
R356 VTAIL.n335 VTAIL.n334 185
R357 VTAIL.n358 VTAIL.n357 185
R358 VTAIL.n356 VTAIL.n355 185
R359 VTAIL.n339 VTAIL.n338 185
R360 VTAIL.n350 VTAIL.n349 185
R361 VTAIL.n348 VTAIL.n347 185
R362 VTAIL.n343 VTAIL.n342 185
R363 VTAIL.n755 VTAIL.t15 147.659
R364 VTAIL.n35 VTAIL.t3 147.659
R365 VTAIL.n137 VTAIL.t8 147.659
R366 VTAIL.n241 VTAIL.t7 147.659
R367 VTAIL.n654 VTAIL.t9 147.659
R368 VTAIL.n550 VTAIL.t10 147.659
R369 VTAIL.n448 VTAIL.t6 147.659
R370 VTAIL.n344 VTAIL.t2 147.659
R371 VTAIL.n759 VTAIL.n753 104.615
R372 VTAIL.n760 VTAIL.n759 104.615
R373 VTAIL.n760 VTAIL.n749 104.615
R374 VTAIL.n767 VTAIL.n749 104.615
R375 VTAIL.n768 VTAIL.n767 104.615
R376 VTAIL.n768 VTAIL.n745 104.615
R377 VTAIL.n775 VTAIL.n745 104.615
R378 VTAIL.n776 VTAIL.n775 104.615
R379 VTAIL.n776 VTAIL.n741 104.615
R380 VTAIL.n783 VTAIL.n741 104.615
R381 VTAIL.n784 VTAIL.n783 104.615
R382 VTAIL.n784 VTAIL.n737 104.615
R383 VTAIL.n791 VTAIL.n737 104.615
R384 VTAIL.n792 VTAIL.n791 104.615
R385 VTAIL.n792 VTAIL.n733 104.615
R386 VTAIL.n800 VTAIL.n733 104.615
R387 VTAIL.n801 VTAIL.n800 104.615
R388 VTAIL.n802 VTAIL.n801 104.615
R389 VTAIL.n802 VTAIL.n729 104.615
R390 VTAIL.n809 VTAIL.n729 104.615
R391 VTAIL.n810 VTAIL.n809 104.615
R392 VTAIL.n810 VTAIL.n725 104.615
R393 VTAIL.n817 VTAIL.n725 104.615
R394 VTAIL.n818 VTAIL.n817 104.615
R395 VTAIL.n39 VTAIL.n33 104.615
R396 VTAIL.n40 VTAIL.n39 104.615
R397 VTAIL.n40 VTAIL.n29 104.615
R398 VTAIL.n47 VTAIL.n29 104.615
R399 VTAIL.n48 VTAIL.n47 104.615
R400 VTAIL.n48 VTAIL.n25 104.615
R401 VTAIL.n55 VTAIL.n25 104.615
R402 VTAIL.n56 VTAIL.n55 104.615
R403 VTAIL.n56 VTAIL.n21 104.615
R404 VTAIL.n63 VTAIL.n21 104.615
R405 VTAIL.n64 VTAIL.n63 104.615
R406 VTAIL.n64 VTAIL.n17 104.615
R407 VTAIL.n71 VTAIL.n17 104.615
R408 VTAIL.n72 VTAIL.n71 104.615
R409 VTAIL.n72 VTAIL.n13 104.615
R410 VTAIL.n80 VTAIL.n13 104.615
R411 VTAIL.n81 VTAIL.n80 104.615
R412 VTAIL.n82 VTAIL.n81 104.615
R413 VTAIL.n82 VTAIL.n9 104.615
R414 VTAIL.n89 VTAIL.n9 104.615
R415 VTAIL.n90 VTAIL.n89 104.615
R416 VTAIL.n90 VTAIL.n5 104.615
R417 VTAIL.n97 VTAIL.n5 104.615
R418 VTAIL.n98 VTAIL.n97 104.615
R419 VTAIL.n141 VTAIL.n135 104.615
R420 VTAIL.n142 VTAIL.n141 104.615
R421 VTAIL.n142 VTAIL.n131 104.615
R422 VTAIL.n149 VTAIL.n131 104.615
R423 VTAIL.n150 VTAIL.n149 104.615
R424 VTAIL.n150 VTAIL.n127 104.615
R425 VTAIL.n157 VTAIL.n127 104.615
R426 VTAIL.n158 VTAIL.n157 104.615
R427 VTAIL.n158 VTAIL.n123 104.615
R428 VTAIL.n165 VTAIL.n123 104.615
R429 VTAIL.n166 VTAIL.n165 104.615
R430 VTAIL.n166 VTAIL.n119 104.615
R431 VTAIL.n173 VTAIL.n119 104.615
R432 VTAIL.n174 VTAIL.n173 104.615
R433 VTAIL.n174 VTAIL.n115 104.615
R434 VTAIL.n182 VTAIL.n115 104.615
R435 VTAIL.n183 VTAIL.n182 104.615
R436 VTAIL.n184 VTAIL.n183 104.615
R437 VTAIL.n184 VTAIL.n111 104.615
R438 VTAIL.n191 VTAIL.n111 104.615
R439 VTAIL.n192 VTAIL.n191 104.615
R440 VTAIL.n192 VTAIL.n107 104.615
R441 VTAIL.n199 VTAIL.n107 104.615
R442 VTAIL.n200 VTAIL.n199 104.615
R443 VTAIL.n245 VTAIL.n239 104.615
R444 VTAIL.n246 VTAIL.n245 104.615
R445 VTAIL.n246 VTAIL.n235 104.615
R446 VTAIL.n253 VTAIL.n235 104.615
R447 VTAIL.n254 VTAIL.n253 104.615
R448 VTAIL.n254 VTAIL.n231 104.615
R449 VTAIL.n261 VTAIL.n231 104.615
R450 VTAIL.n262 VTAIL.n261 104.615
R451 VTAIL.n262 VTAIL.n227 104.615
R452 VTAIL.n269 VTAIL.n227 104.615
R453 VTAIL.n270 VTAIL.n269 104.615
R454 VTAIL.n270 VTAIL.n223 104.615
R455 VTAIL.n277 VTAIL.n223 104.615
R456 VTAIL.n278 VTAIL.n277 104.615
R457 VTAIL.n278 VTAIL.n219 104.615
R458 VTAIL.n286 VTAIL.n219 104.615
R459 VTAIL.n287 VTAIL.n286 104.615
R460 VTAIL.n288 VTAIL.n287 104.615
R461 VTAIL.n288 VTAIL.n215 104.615
R462 VTAIL.n295 VTAIL.n215 104.615
R463 VTAIL.n296 VTAIL.n295 104.615
R464 VTAIL.n296 VTAIL.n211 104.615
R465 VTAIL.n303 VTAIL.n211 104.615
R466 VTAIL.n304 VTAIL.n303 104.615
R467 VTAIL.n716 VTAIL.n715 104.615
R468 VTAIL.n715 VTAIL.n623 104.615
R469 VTAIL.n708 VTAIL.n623 104.615
R470 VTAIL.n708 VTAIL.n707 104.615
R471 VTAIL.n707 VTAIL.n627 104.615
R472 VTAIL.n700 VTAIL.n627 104.615
R473 VTAIL.n700 VTAIL.n699 104.615
R474 VTAIL.n699 VTAIL.n698 104.615
R475 VTAIL.n698 VTAIL.n631 104.615
R476 VTAIL.n691 VTAIL.n631 104.615
R477 VTAIL.n691 VTAIL.n690 104.615
R478 VTAIL.n690 VTAIL.n636 104.615
R479 VTAIL.n683 VTAIL.n636 104.615
R480 VTAIL.n683 VTAIL.n682 104.615
R481 VTAIL.n682 VTAIL.n640 104.615
R482 VTAIL.n675 VTAIL.n640 104.615
R483 VTAIL.n675 VTAIL.n674 104.615
R484 VTAIL.n674 VTAIL.n644 104.615
R485 VTAIL.n667 VTAIL.n644 104.615
R486 VTAIL.n667 VTAIL.n666 104.615
R487 VTAIL.n666 VTAIL.n648 104.615
R488 VTAIL.n659 VTAIL.n648 104.615
R489 VTAIL.n659 VTAIL.n658 104.615
R490 VTAIL.n658 VTAIL.n652 104.615
R491 VTAIL.n612 VTAIL.n611 104.615
R492 VTAIL.n611 VTAIL.n519 104.615
R493 VTAIL.n604 VTAIL.n519 104.615
R494 VTAIL.n604 VTAIL.n603 104.615
R495 VTAIL.n603 VTAIL.n523 104.615
R496 VTAIL.n596 VTAIL.n523 104.615
R497 VTAIL.n596 VTAIL.n595 104.615
R498 VTAIL.n595 VTAIL.n594 104.615
R499 VTAIL.n594 VTAIL.n527 104.615
R500 VTAIL.n587 VTAIL.n527 104.615
R501 VTAIL.n587 VTAIL.n586 104.615
R502 VTAIL.n586 VTAIL.n532 104.615
R503 VTAIL.n579 VTAIL.n532 104.615
R504 VTAIL.n579 VTAIL.n578 104.615
R505 VTAIL.n578 VTAIL.n536 104.615
R506 VTAIL.n571 VTAIL.n536 104.615
R507 VTAIL.n571 VTAIL.n570 104.615
R508 VTAIL.n570 VTAIL.n540 104.615
R509 VTAIL.n563 VTAIL.n540 104.615
R510 VTAIL.n563 VTAIL.n562 104.615
R511 VTAIL.n562 VTAIL.n544 104.615
R512 VTAIL.n555 VTAIL.n544 104.615
R513 VTAIL.n555 VTAIL.n554 104.615
R514 VTAIL.n554 VTAIL.n548 104.615
R515 VTAIL.n510 VTAIL.n509 104.615
R516 VTAIL.n509 VTAIL.n417 104.615
R517 VTAIL.n502 VTAIL.n417 104.615
R518 VTAIL.n502 VTAIL.n501 104.615
R519 VTAIL.n501 VTAIL.n421 104.615
R520 VTAIL.n494 VTAIL.n421 104.615
R521 VTAIL.n494 VTAIL.n493 104.615
R522 VTAIL.n493 VTAIL.n492 104.615
R523 VTAIL.n492 VTAIL.n425 104.615
R524 VTAIL.n485 VTAIL.n425 104.615
R525 VTAIL.n485 VTAIL.n484 104.615
R526 VTAIL.n484 VTAIL.n430 104.615
R527 VTAIL.n477 VTAIL.n430 104.615
R528 VTAIL.n477 VTAIL.n476 104.615
R529 VTAIL.n476 VTAIL.n434 104.615
R530 VTAIL.n469 VTAIL.n434 104.615
R531 VTAIL.n469 VTAIL.n468 104.615
R532 VTAIL.n468 VTAIL.n438 104.615
R533 VTAIL.n461 VTAIL.n438 104.615
R534 VTAIL.n461 VTAIL.n460 104.615
R535 VTAIL.n460 VTAIL.n442 104.615
R536 VTAIL.n453 VTAIL.n442 104.615
R537 VTAIL.n453 VTAIL.n452 104.615
R538 VTAIL.n452 VTAIL.n446 104.615
R539 VTAIL.n406 VTAIL.n405 104.615
R540 VTAIL.n405 VTAIL.n313 104.615
R541 VTAIL.n398 VTAIL.n313 104.615
R542 VTAIL.n398 VTAIL.n397 104.615
R543 VTAIL.n397 VTAIL.n317 104.615
R544 VTAIL.n390 VTAIL.n317 104.615
R545 VTAIL.n390 VTAIL.n389 104.615
R546 VTAIL.n389 VTAIL.n388 104.615
R547 VTAIL.n388 VTAIL.n321 104.615
R548 VTAIL.n381 VTAIL.n321 104.615
R549 VTAIL.n381 VTAIL.n380 104.615
R550 VTAIL.n380 VTAIL.n326 104.615
R551 VTAIL.n373 VTAIL.n326 104.615
R552 VTAIL.n373 VTAIL.n372 104.615
R553 VTAIL.n372 VTAIL.n330 104.615
R554 VTAIL.n365 VTAIL.n330 104.615
R555 VTAIL.n365 VTAIL.n364 104.615
R556 VTAIL.n364 VTAIL.n334 104.615
R557 VTAIL.n357 VTAIL.n334 104.615
R558 VTAIL.n357 VTAIL.n356 104.615
R559 VTAIL.n356 VTAIL.n338 104.615
R560 VTAIL.n349 VTAIL.n338 104.615
R561 VTAIL.n349 VTAIL.n348 104.615
R562 VTAIL.n348 VTAIL.n342 104.615
R563 VTAIL.t15 VTAIL.n753 52.3082
R564 VTAIL.t3 VTAIL.n33 52.3082
R565 VTAIL.t8 VTAIL.n135 52.3082
R566 VTAIL.t7 VTAIL.n239 52.3082
R567 VTAIL.t9 VTAIL.n652 52.3082
R568 VTAIL.t10 VTAIL.n548 52.3082
R569 VTAIL.t6 VTAIL.n446 52.3082
R570 VTAIL.t2 VTAIL.n342 52.3082
R571 VTAIL.n619 VTAIL.n618 41.8362
R572 VTAIL.n413 VTAIL.n412 41.8362
R573 VTAIL.n1 VTAIL.n0 41.836
R574 VTAIL.n207 VTAIL.n206 41.836
R575 VTAIL.n823 VTAIL.n721 31.4014
R576 VTAIL.n411 VTAIL.n309 31.4014
R577 VTAIL.n823 VTAIL.n822 30.052
R578 VTAIL.n103 VTAIL.n102 30.052
R579 VTAIL.n205 VTAIL.n204 30.052
R580 VTAIL.n309 VTAIL.n308 30.052
R581 VTAIL.n721 VTAIL.n720 30.052
R582 VTAIL.n617 VTAIL.n616 30.052
R583 VTAIL.n515 VTAIL.n514 30.052
R584 VTAIL.n411 VTAIL.n410 30.052
R585 VTAIL.n755 VTAIL.n754 15.6677
R586 VTAIL.n35 VTAIL.n34 15.6677
R587 VTAIL.n137 VTAIL.n136 15.6677
R588 VTAIL.n241 VTAIL.n240 15.6677
R589 VTAIL.n654 VTAIL.n653 15.6677
R590 VTAIL.n550 VTAIL.n549 15.6677
R591 VTAIL.n448 VTAIL.n447 15.6677
R592 VTAIL.n344 VTAIL.n343 15.6677
R593 VTAIL.n803 VTAIL.n732 13.1884
R594 VTAIL.n83 VTAIL.n12 13.1884
R595 VTAIL.n185 VTAIL.n114 13.1884
R596 VTAIL.n289 VTAIL.n218 13.1884
R597 VTAIL.n701 VTAIL.n630 13.1884
R598 VTAIL.n597 VTAIL.n526 13.1884
R599 VTAIL.n495 VTAIL.n424 13.1884
R600 VTAIL.n391 VTAIL.n320 13.1884
R601 VTAIL.n758 VTAIL.n757 12.8005
R602 VTAIL.n799 VTAIL.n798 12.8005
R603 VTAIL.n804 VTAIL.n730 12.8005
R604 VTAIL.n38 VTAIL.n37 12.8005
R605 VTAIL.n79 VTAIL.n78 12.8005
R606 VTAIL.n84 VTAIL.n10 12.8005
R607 VTAIL.n140 VTAIL.n139 12.8005
R608 VTAIL.n181 VTAIL.n180 12.8005
R609 VTAIL.n186 VTAIL.n112 12.8005
R610 VTAIL.n244 VTAIL.n243 12.8005
R611 VTAIL.n285 VTAIL.n284 12.8005
R612 VTAIL.n290 VTAIL.n216 12.8005
R613 VTAIL.n702 VTAIL.n628 12.8005
R614 VTAIL.n697 VTAIL.n632 12.8005
R615 VTAIL.n657 VTAIL.n656 12.8005
R616 VTAIL.n598 VTAIL.n524 12.8005
R617 VTAIL.n593 VTAIL.n528 12.8005
R618 VTAIL.n553 VTAIL.n552 12.8005
R619 VTAIL.n496 VTAIL.n422 12.8005
R620 VTAIL.n491 VTAIL.n426 12.8005
R621 VTAIL.n451 VTAIL.n450 12.8005
R622 VTAIL.n392 VTAIL.n318 12.8005
R623 VTAIL.n387 VTAIL.n322 12.8005
R624 VTAIL.n347 VTAIL.n346 12.8005
R625 VTAIL.n761 VTAIL.n752 12.0247
R626 VTAIL.n797 VTAIL.n734 12.0247
R627 VTAIL.n808 VTAIL.n807 12.0247
R628 VTAIL.n41 VTAIL.n32 12.0247
R629 VTAIL.n77 VTAIL.n14 12.0247
R630 VTAIL.n88 VTAIL.n87 12.0247
R631 VTAIL.n143 VTAIL.n134 12.0247
R632 VTAIL.n179 VTAIL.n116 12.0247
R633 VTAIL.n190 VTAIL.n189 12.0247
R634 VTAIL.n247 VTAIL.n238 12.0247
R635 VTAIL.n283 VTAIL.n220 12.0247
R636 VTAIL.n294 VTAIL.n293 12.0247
R637 VTAIL.n706 VTAIL.n705 12.0247
R638 VTAIL.n696 VTAIL.n633 12.0247
R639 VTAIL.n660 VTAIL.n651 12.0247
R640 VTAIL.n602 VTAIL.n601 12.0247
R641 VTAIL.n592 VTAIL.n529 12.0247
R642 VTAIL.n556 VTAIL.n547 12.0247
R643 VTAIL.n500 VTAIL.n499 12.0247
R644 VTAIL.n490 VTAIL.n427 12.0247
R645 VTAIL.n454 VTAIL.n445 12.0247
R646 VTAIL.n396 VTAIL.n395 12.0247
R647 VTAIL.n386 VTAIL.n323 12.0247
R648 VTAIL.n350 VTAIL.n341 12.0247
R649 VTAIL.n762 VTAIL.n750 11.249
R650 VTAIL.n794 VTAIL.n793 11.249
R651 VTAIL.n811 VTAIL.n728 11.249
R652 VTAIL.n42 VTAIL.n30 11.249
R653 VTAIL.n74 VTAIL.n73 11.249
R654 VTAIL.n91 VTAIL.n8 11.249
R655 VTAIL.n144 VTAIL.n132 11.249
R656 VTAIL.n176 VTAIL.n175 11.249
R657 VTAIL.n193 VTAIL.n110 11.249
R658 VTAIL.n248 VTAIL.n236 11.249
R659 VTAIL.n280 VTAIL.n279 11.249
R660 VTAIL.n297 VTAIL.n214 11.249
R661 VTAIL.n709 VTAIL.n626 11.249
R662 VTAIL.n693 VTAIL.n692 11.249
R663 VTAIL.n661 VTAIL.n649 11.249
R664 VTAIL.n605 VTAIL.n522 11.249
R665 VTAIL.n589 VTAIL.n588 11.249
R666 VTAIL.n557 VTAIL.n545 11.249
R667 VTAIL.n503 VTAIL.n420 11.249
R668 VTAIL.n487 VTAIL.n486 11.249
R669 VTAIL.n455 VTAIL.n443 11.249
R670 VTAIL.n399 VTAIL.n316 11.249
R671 VTAIL.n383 VTAIL.n382 11.249
R672 VTAIL.n351 VTAIL.n339 11.249
R673 VTAIL.n766 VTAIL.n765 10.4732
R674 VTAIL.n790 VTAIL.n736 10.4732
R675 VTAIL.n812 VTAIL.n726 10.4732
R676 VTAIL.n46 VTAIL.n45 10.4732
R677 VTAIL.n70 VTAIL.n16 10.4732
R678 VTAIL.n92 VTAIL.n6 10.4732
R679 VTAIL.n148 VTAIL.n147 10.4732
R680 VTAIL.n172 VTAIL.n118 10.4732
R681 VTAIL.n194 VTAIL.n108 10.4732
R682 VTAIL.n252 VTAIL.n251 10.4732
R683 VTAIL.n276 VTAIL.n222 10.4732
R684 VTAIL.n298 VTAIL.n212 10.4732
R685 VTAIL.n710 VTAIL.n624 10.4732
R686 VTAIL.n689 VTAIL.n635 10.4732
R687 VTAIL.n665 VTAIL.n664 10.4732
R688 VTAIL.n606 VTAIL.n520 10.4732
R689 VTAIL.n585 VTAIL.n531 10.4732
R690 VTAIL.n561 VTAIL.n560 10.4732
R691 VTAIL.n504 VTAIL.n418 10.4732
R692 VTAIL.n483 VTAIL.n429 10.4732
R693 VTAIL.n459 VTAIL.n458 10.4732
R694 VTAIL.n400 VTAIL.n314 10.4732
R695 VTAIL.n379 VTAIL.n325 10.4732
R696 VTAIL.n355 VTAIL.n354 10.4732
R697 VTAIL.n769 VTAIL.n748 9.69747
R698 VTAIL.n789 VTAIL.n738 9.69747
R699 VTAIL.n816 VTAIL.n815 9.69747
R700 VTAIL.n49 VTAIL.n28 9.69747
R701 VTAIL.n69 VTAIL.n18 9.69747
R702 VTAIL.n96 VTAIL.n95 9.69747
R703 VTAIL.n151 VTAIL.n130 9.69747
R704 VTAIL.n171 VTAIL.n120 9.69747
R705 VTAIL.n198 VTAIL.n197 9.69747
R706 VTAIL.n255 VTAIL.n234 9.69747
R707 VTAIL.n275 VTAIL.n224 9.69747
R708 VTAIL.n302 VTAIL.n301 9.69747
R709 VTAIL.n714 VTAIL.n713 9.69747
R710 VTAIL.n688 VTAIL.n637 9.69747
R711 VTAIL.n668 VTAIL.n647 9.69747
R712 VTAIL.n610 VTAIL.n609 9.69747
R713 VTAIL.n584 VTAIL.n533 9.69747
R714 VTAIL.n564 VTAIL.n543 9.69747
R715 VTAIL.n508 VTAIL.n507 9.69747
R716 VTAIL.n482 VTAIL.n431 9.69747
R717 VTAIL.n462 VTAIL.n441 9.69747
R718 VTAIL.n404 VTAIL.n403 9.69747
R719 VTAIL.n378 VTAIL.n327 9.69747
R720 VTAIL.n358 VTAIL.n337 9.69747
R721 VTAIL.n822 VTAIL.n821 9.45567
R722 VTAIL.n102 VTAIL.n101 9.45567
R723 VTAIL.n204 VTAIL.n203 9.45567
R724 VTAIL.n308 VTAIL.n307 9.45567
R725 VTAIL.n720 VTAIL.n719 9.45567
R726 VTAIL.n616 VTAIL.n615 9.45567
R727 VTAIL.n514 VTAIL.n513 9.45567
R728 VTAIL.n410 VTAIL.n409 9.45567
R729 VTAIL.n821 VTAIL.n820 9.3005
R730 VTAIL.n724 VTAIL.n723 9.3005
R731 VTAIL.n815 VTAIL.n814 9.3005
R732 VTAIL.n813 VTAIL.n812 9.3005
R733 VTAIL.n728 VTAIL.n727 9.3005
R734 VTAIL.n807 VTAIL.n806 9.3005
R735 VTAIL.n805 VTAIL.n804 9.3005
R736 VTAIL.n744 VTAIL.n743 9.3005
R737 VTAIL.n773 VTAIL.n772 9.3005
R738 VTAIL.n771 VTAIL.n770 9.3005
R739 VTAIL.n748 VTAIL.n747 9.3005
R740 VTAIL.n765 VTAIL.n764 9.3005
R741 VTAIL.n763 VTAIL.n762 9.3005
R742 VTAIL.n752 VTAIL.n751 9.3005
R743 VTAIL.n757 VTAIL.n756 9.3005
R744 VTAIL.n779 VTAIL.n778 9.3005
R745 VTAIL.n781 VTAIL.n780 9.3005
R746 VTAIL.n740 VTAIL.n739 9.3005
R747 VTAIL.n787 VTAIL.n786 9.3005
R748 VTAIL.n789 VTAIL.n788 9.3005
R749 VTAIL.n736 VTAIL.n735 9.3005
R750 VTAIL.n795 VTAIL.n794 9.3005
R751 VTAIL.n797 VTAIL.n796 9.3005
R752 VTAIL.n798 VTAIL.n731 9.3005
R753 VTAIL.n101 VTAIL.n100 9.3005
R754 VTAIL.n4 VTAIL.n3 9.3005
R755 VTAIL.n95 VTAIL.n94 9.3005
R756 VTAIL.n93 VTAIL.n92 9.3005
R757 VTAIL.n8 VTAIL.n7 9.3005
R758 VTAIL.n87 VTAIL.n86 9.3005
R759 VTAIL.n85 VTAIL.n84 9.3005
R760 VTAIL.n24 VTAIL.n23 9.3005
R761 VTAIL.n53 VTAIL.n52 9.3005
R762 VTAIL.n51 VTAIL.n50 9.3005
R763 VTAIL.n28 VTAIL.n27 9.3005
R764 VTAIL.n45 VTAIL.n44 9.3005
R765 VTAIL.n43 VTAIL.n42 9.3005
R766 VTAIL.n32 VTAIL.n31 9.3005
R767 VTAIL.n37 VTAIL.n36 9.3005
R768 VTAIL.n59 VTAIL.n58 9.3005
R769 VTAIL.n61 VTAIL.n60 9.3005
R770 VTAIL.n20 VTAIL.n19 9.3005
R771 VTAIL.n67 VTAIL.n66 9.3005
R772 VTAIL.n69 VTAIL.n68 9.3005
R773 VTAIL.n16 VTAIL.n15 9.3005
R774 VTAIL.n75 VTAIL.n74 9.3005
R775 VTAIL.n77 VTAIL.n76 9.3005
R776 VTAIL.n78 VTAIL.n11 9.3005
R777 VTAIL.n203 VTAIL.n202 9.3005
R778 VTAIL.n106 VTAIL.n105 9.3005
R779 VTAIL.n197 VTAIL.n196 9.3005
R780 VTAIL.n195 VTAIL.n194 9.3005
R781 VTAIL.n110 VTAIL.n109 9.3005
R782 VTAIL.n189 VTAIL.n188 9.3005
R783 VTAIL.n187 VTAIL.n186 9.3005
R784 VTAIL.n126 VTAIL.n125 9.3005
R785 VTAIL.n155 VTAIL.n154 9.3005
R786 VTAIL.n153 VTAIL.n152 9.3005
R787 VTAIL.n130 VTAIL.n129 9.3005
R788 VTAIL.n147 VTAIL.n146 9.3005
R789 VTAIL.n145 VTAIL.n144 9.3005
R790 VTAIL.n134 VTAIL.n133 9.3005
R791 VTAIL.n139 VTAIL.n138 9.3005
R792 VTAIL.n161 VTAIL.n160 9.3005
R793 VTAIL.n163 VTAIL.n162 9.3005
R794 VTAIL.n122 VTAIL.n121 9.3005
R795 VTAIL.n169 VTAIL.n168 9.3005
R796 VTAIL.n171 VTAIL.n170 9.3005
R797 VTAIL.n118 VTAIL.n117 9.3005
R798 VTAIL.n177 VTAIL.n176 9.3005
R799 VTAIL.n179 VTAIL.n178 9.3005
R800 VTAIL.n180 VTAIL.n113 9.3005
R801 VTAIL.n307 VTAIL.n306 9.3005
R802 VTAIL.n210 VTAIL.n209 9.3005
R803 VTAIL.n301 VTAIL.n300 9.3005
R804 VTAIL.n299 VTAIL.n298 9.3005
R805 VTAIL.n214 VTAIL.n213 9.3005
R806 VTAIL.n293 VTAIL.n292 9.3005
R807 VTAIL.n291 VTAIL.n290 9.3005
R808 VTAIL.n230 VTAIL.n229 9.3005
R809 VTAIL.n259 VTAIL.n258 9.3005
R810 VTAIL.n257 VTAIL.n256 9.3005
R811 VTAIL.n234 VTAIL.n233 9.3005
R812 VTAIL.n251 VTAIL.n250 9.3005
R813 VTAIL.n249 VTAIL.n248 9.3005
R814 VTAIL.n238 VTAIL.n237 9.3005
R815 VTAIL.n243 VTAIL.n242 9.3005
R816 VTAIL.n265 VTAIL.n264 9.3005
R817 VTAIL.n267 VTAIL.n266 9.3005
R818 VTAIL.n226 VTAIL.n225 9.3005
R819 VTAIL.n273 VTAIL.n272 9.3005
R820 VTAIL.n275 VTAIL.n274 9.3005
R821 VTAIL.n222 VTAIL.n221 9.3005
R822 VTAIL.n281 VTAIL.n280 9.3005
R823 VTAIL.n283 VTAIL.n282 9.3005
R824 VTAIL.n284 VTAIL.n217 9.3005
R825 VTAIL.n680 VTAIL.n679 9.3005
R826 VTAIL.n639 VTAIL.n638 9.3005
R827 VTAIL.n686 VTAIL.n685 9.3005
R828 VTAIL.n688 VTAIL.n687 9.3005
R829 VTAIL.n635 VTAIL.n634 9.3005
R830 VTAIL.n694 VTAIL.n693 9.3005
R831 VTAIL.n696 VTAIL.n695 9.3005
R832 VTAIL.n632 VTAIL.n629 9.3005
R833 VTAIL.n719 VTAIL.n718 9.3005
R834 VTAIL.n622 VTAIL.n621 9.3005
R835 VTAIL.n713 VTAIL.n712 9.3005
R836 VTAIL.n711 VTAIL.n710 9.3005
R837 VTAIL.n626 VTAIL.n625 9.3005
R838 VTAIL.n705 VTAIL.n704 9.3005
R839 VTAIL.n703 VTAIL.n702 9.3005
R840 VTAIL.n678 VTAIL.n677 9.3005
R841 VTAIL.n643 VTAIL.n642 9.3005
R842 VTAIL.n672 VTAIL.n671 9.3005
R843 VTAIL.n670 VTAIL.n669 9.3005
R844 VTAIL.n647 VTAIL.n646 9.3005
R845 VTAIL.n664 VTAIL.n663 9.3005
R846 VTAIL.n662 VTAIL.n661 9.3005
R847 VTAIL.n651 VTAIL.n650 9.3005
R848 VTAIL.n656 VTAIL.n655 9.3005
R849 VTAIL.n576 VTAIL.n575 9.3005
R850 VTAIL.n535 VTAIL.n534 9.3005
R851 VTAIL.n582 VTAIL.n581 9.3005
R852 VTAIL.n584 VTAIL.n583 9.3005
R853 VTAIL.n531 VTAIL.n530 9.3005
R854 VTAIL.n590 VTAIL.n589 9.3005
R855 VTAIL.n592 VTAIL.n591 9.3005
R856 VTAIL.n528 VTAIL.n525 9.3005
R857 VTAIL.n615 VTAIL.n614 9.3005
R858 VTAIL.n518 VTAIL.n517 9.3005
R859 VTAIL.n609 VTAIL.n608 9.3005
R860 VTAIL.n607 VTAIL.n606 9.3005
R861 VTAIL.n522 VTAIL.n521 9.3005
R862 VTAIL.n601 VTAIL.n600 9.3005
R863 VTAIL.n599 VTAIL.n598 9.3005
R864 VTAIL.n574 VTAIL.n573 9.3005
R865 VTAIL.n539 VTAIL.n538 9.3005
R866 VTAIL.n568 VTAIL.n567 9.3005
R867 VTAIL.n566 VTAIL.n565 9.3005
R868 VTAIL.n543 VTAIL.n542 9.3005
R869 VTAIL.n560 VTAIL.n559 9.3005
R870 VTAIL.n558 VTAIL.n557 9.3005
R871 VTAIL.n547 VTAIL.n546 9.3005
R872 VTAIL.n552 VTAIL.n551 9.3005
R873 VTAIL.n474 VTAIL.n473 9.3005
R874 VTAIL.n433 VTAIL.n432 9.3005
R875 VTAIL.n480 VTAIL.n479 9.3005
R876 VTAIL.n482 VTAIL.n481 9.3005
R877 VTAIL.n429 VTAIL.n428 9.3005
R878 VTAIL.n488 VTAIL.n487 9.3005
R879 VTAIL.n490 VTAIL.n489 9.3005
R880 VTAIL.n426 VTAIL.n423 9.3005
R881 VTAIL.n513 VTAIL.n512 9.3005
R882 VTAIL.n416 VTAIL.n415 9.3005
R883 VTAIL.n507 VTAIL.n506 9.3005
R884 VTAIL.n505 VTAIL.n504 9.3005
R885 VTAIL.n420 VTAIL.n419 9.3005
R886 VTAIL.n499 VTAIL.n498 9.3005
R887 VTAIL.n497 VTAIL.n496 9.3005
R888 VTAIL.n472 VTAIL.n471 9.3005
R889 VTAIL.n437 VTAIL.n436 9.3005
R890 VTAIL.n466 VTAIL.n465 9.3005
R891 VTAIL.n464 VTAIL.n463 9.3005
R892 VTAIL.n441 VTAIL.n440 9.3005
R893 VTAIL.n458 VTAIL.n457 9.3005
R894 VTAIL.n456 VTAIL.n455 9.3005
R895 VTAIL.n445 VTAIL.n444 9.3005
R896 VTAIL.n450 VTAIL.n449 9.3005
R897 VTAIL.n370 VTAIL.n369 9.3005
R898 VTAIL.n329 VTAIL.n328 9.3005
R899 VTAIL.n376 VTAIL.n375 9.3005
R900 VTAIL.n378 VTAIL.n377 9.3005
R901 VTAIL.n325 VTAIL.n324 9.3005
R902 VTAIL.n384 VTAIL.n383 9.3005
R903 VTAIL.n386 VTAIL.n385 9.3005
R904 VTAIL.n322 VTAIL.n319 9.3005
R905 VTAIL.n409 VTAIL.n408 9.3005
R906 VTAIL.n312 VTAIL.n311 9.3005
R907 VTAIL.n403 VTAIL.n402 9.3005
R908 VTAIL.n401 VTAIL.n400 9.3005
R909 VTAIL.n316 VTAIL.n315 9.3005
R910 VTAIL.n395 VTAIL.n394 9.3005
R911 VTAIL.n393 VTAIL.n392 9.3005
R912 VTAIL.n368 VTAIL.n367 9.3005
R913 VTAIL.n333 VTAIL.n332 9.3005
R914 VTAIL.n362 VTAIL.n361 9.3005
R915 VTAIL.n360 VTAIL.n359 9.3005
R916 VTAIL.n337 VTAIL.n336 9.3005
R917 VTAIL.n354 VTAIL.n353 9.3005
R918 VTAIL.n352 VTAIL.n351 9.3005
R919 VTAIL.n341 VTAIL.n340 9.3005
R920 VTAIL.n346 VTAIL.n345 9.3005
R921 VTAIL.n770 VTAIL.n746 8.92171
R922 VTAIL.n786 VTAIL.n785 8.92171
R923 VTAIL.n819 VTAIL.n724 8.92171
R924 VTAIL.n50 VTAIL.n26 8.92171
R925 VTAIL.n66 VTAIL.n65 8.92171
R926 VTAIL.n99 VTAIL.n4 8.92171
R927 VTAIL.n152 VTAIL.n128 8.92171
R928 VTAIL.n168 VTAIL.n167 8.92171
R929 VTAIL.n201 VTAIL.n106 8.92171
R930 VTAIL.n256 VTAIL.n232 8.92171
R931 VTAIL.n272 VTAIL.n271 8.92171
R932 VTAIL.n305 VTAIL.n210 8.92171
R933 VTAIL.n717 VTAIL.n622 8.92171
R934 VTAIL.n685 VTAIL.n684 8.92171
R935 VTAIL.n669 VTAIL.n645 8.92171
R936 VTAIL.n613 VTAIL.n518 8.92171
R937 VTAIL.n581 VTAIL.n580 8.92171
R938 VTAIL.n565 VTAIL.n541 8.92171
R939 VTAIL.n511 VTAIL.n416 8.92171
R940 VTAIL.n479 VTAIL.n478 8.92171
R941 VTAIL.n463 VTAIL.n439 8.92171
R942 VTAIL.n407 VTAIL.n312 8.92171
R943 VTAIL.n375 VTAIL.n374 8.92171
R944 VTAIL.n359 VTAIL.n335 8.92171
R945 VTAIL.n774 VTAIL.n773 8.14595
R946 VTAIL.n782 VTAIL.n740 8.14595
R947 VTAIL.n820 VTAIL.n722 8.14595
R948 VTAIL.n54 VTAIL.n53 8.14595
R949 VTAIL.n62 VTAIL.n20 8.14595
R950 VTAIL.n100 VTAIL.n2 8.14595
R951 VTAIL.n156 VTAIL.n155 8.14595
R952 VTAIL.n164 VTAIL.n122 8.14595
R953 VTAIL.n202 VTAIL.n104 8.14595
R954 VTAIL.n260 VTAIL.n259 8.14595
R955 VTAIL.n268 VTAIL.n226 8.14595
R956 VTAIL.n306 VTAIL.n208 8.14595
R957 VTAIL.n718 VTAIL.n620 8.14595
R958 VTAIL.n681 VTAIL.n639 8.14595
R959 VTAIL.n673 VTAIL.n672 8.14595
R960 VTAIL.n614 VTAIL.n516 8.14595
R961 VTAIL.n577 VTAIL.n535 8.14595
R962 VTAIL.n569 VTAIL.n568 8.14595
R963 VTAIL.n512 VTAIL.n414 8.14595
R964 VTAIL.n475 VTAIL.n433 8.14595
R965 VTAIL.n467 VTAIL.n466 8.14595
R966 VTAIL.n408 VTAIL.n310 8.14595
R967 VTAIL.n371 VTAIL.n329 8.14595
R968 VTAIL.n363 VTAIL.n362 8.14595
R969 VTAIL.n777 VTAIL.n744 7.3702
R970 VTAIL.n781 VTAIL.n742 7.3702
R971 VTAIL.n57 VTAIL.n24 7.3702
R972 VTAIL.n61 VTAIL.n22 7.3702
R973 VTAIL.n159 VTAIL.n126 7.3702
R974 VTAIL.n163 VTAIL.n124 7.3702
R975 VTAIL.n263 VTAIL.n230 7.3702
R976 VTAIL.n267 VTAIL.n228 7.3702
R977 VTAIL.n680 VTAIL.n641 7.3702
R978 VTAIL.n676 VTAIL.n643 7.3702
R979 VTAIL.n576 VTAIL.n537 7.3702
R980 VTAIL.n572 VTAIL.n539 7.3702
R981 VTAIL.n474 VTAIL.n435 7.3702
R982 VTAIL.n470 VTAIL.n437 7.3702
R983 VTAIL.n370 VTAIL.n331 7.3702
R984 VTAIL.n366 VTAIL.n333 7.3702
R985 VTAIL.n778 VTAIL.n777 6.59444
R986 VTAIL.n778 VTAIL.n742 6.59444
R987 VTAIL.n58 VTAIL.n57 6.59444
R988 VTAIL.n58 VTAIL.n22 6.59444
R989 VTAIL.n160 VTAIL.n159 6.59444
R990 VTAIL.n160 VTAIL.n124 6.59444
R991 VTAIL.n264 VTAIL.n263 6.59444
R992 VTAIL.n264 VTAIL.n228 6.59444
R993 VTAIL.n677 VTAIL.n641 6.59444
R994 VTAIL.n677 VTAIL.n676 6.59444
R995 VTAIL.n573 VTAIL.n537 6.59444
R996 VTAIL.n573 VTAIL.n572 6.59444
R997 VTAIL.n471 VTAIL.n435 6.59444
R998 VTAIL.n471 VTAIL.n470 6.59444
R999 VTAIL.n367 VTAIL.n331 6.59444
R1000 VTAIL.n367 VTAIL.n366 6.59444
R1001 VTAIL.n774 VTAIL.n744 5.81868
R1002 VTAIL.n782 VTAIL.n781 5.81868
R1003 VTAIL.n822 VTAIL.n722 5.81868
R1004 VTAIL.n54 VTAIL.n24 5.81868
R1005 VTAIL.n62 VTAIL.n61 5.81868
R1006 VTAIL.n102 VTAIL.n2 5.81868
R1007 VTAIL.n156 VTAIL.n126 5.81868
R1008 VTAIL.n164 VTAIL.n163 5.81868
R1009 VTAIL.n204 VTAIL.n104 5.81868
R1010 VTAIL.n260 VTAIL.n230 5.81868
R1011 VTAIL.n268 VTAIL.n267 5.81868
R1012 VTAIL.n308 VTAIL.n208 5.81868
R1013 VTAIL.n720 VTAIL.n620 5.81868
R1014 VTAIL.n681 VTAIL.n680 5.81868
R1015 VTAIL.n673 VTAIL.n643 5.81868
R1016 VTAIL.n616 VTAIL.n516 5.81868
R1017 VTAIL.n577 VTAIL.n576 5.81868
R1018 VTAIL.n569 VTAIL.n539 5.81868
R1019 VTAIL.n514 VTAIL.n414 5.81868
R1020 VTAIL.n475 VTAIL.n474 5.81868
R1021 VTAIL.n467 VTAIL.n437 5.81868
R1022 VTAIL.n410 VTAIL.n310 5.81868
R1023 VTAIL.n371 VTAIL.n370 5.81868
R1024 VTAIL.n363 VTAIL.n333 5.81868
R1025 VTAIL.n773 VTAIL.n746 5.04292
R1026 VTAIL.n785 VTAIL.n740 5.04292
R1027 VTAIL.n820 VTAIL.n819 5.04292
R1028 VTAIL.n53 VTAIL.n26 5.04292
R1029 VTAIL.n65 VTAIL.n20 5.04292
R1030 VTAIL.n100 VTAIL.n99 5.04292
R1031 VTAIL.n155 VTAIL.n128 5.04292
R1032 VTAIL.n167 VTAIL.n122 5.04292
R1033 VTAIL.n202 VTAIL.n201 5.04292
R1034 VTAIL.n259 VTAIL.n232 5.04292
R1035 VTAIL.n271 VTAIL.n226 5.04292
R1036 VTAIL.n306 VTAIL.n305 5.04292
R1037 VTAIL.n718 VTAIL.n717 5.04292
R1038 VTAIL.n684 VTAIL.n639 5.04292
R1039 VTAIL.n672 VTAIL.n645 5.04292
R1040 VTAIL.n614 VTAIL.n613 5.04292
R1041 VTAIL.n580 VTAIL.n535 5.04292
R1042 VTAIL.n568 VTAIL.n541 5.04292
R1043 VTAIL.n512 VTAIL.n511 5.04292
R1044 VTAIL.n478 VTAIL.n433 5.04292
R1045 VTAIL.n466 VTAIL.n439 5.04292
R1046 VTAIL.n408 VTAIL.n407 5.04292
R1047 VTAIL.n374 VTAIL.n329 5.04292
R1048 VTAIL.n362 VTAIL.n335 5.04292
R1049 VTAIL.n756 VTAIL.n755 4.38563
R1050 VTAIL.n36 VTAIL.n35 4.38563
R1051 VTAIL.n138 VTAIL.n137 4.38563
R1052 VTAIL.n242 VTAIL.n241 4.38563
R1053 VTAIL.n655 VTAIL.n654 4.38563
R1054 VTAIL.n551 VTAIL.n550 4.38563
R1055 VTAIL.n449 VTAIL.n448 4.38563
R1056 VTAIL.n345 VTAIL.n344 4.38563
R1057 VTAIL.n770 VTAIL.n769 4.26717
R1058 VTAIL.n786 VTAIL.n738 4.26717
R1059 VTAIL.n816 VTAIL.n724 4.26717
R1060 VTAIL.n50 VTAIL.n49 4.26717
R1061 VTAIL.n66 VTAIL.n18 4.26717
R1062 VTAIL.n96 VTAIL.n4 4.26717
R1063 VTAIL.n152 VTAIL.n151 4.26717
R1064 VTAIL.n168 VTAIL.n120 4.26717
R1065 VTAIL.n198 VTAIL.n106 4.26717
R1066 VTAIL.n256 VTAIL.n255 4.26717
R1067 VTAIL.n272 VTAIL.n224 4.26717
R1068 VTAIL.n302 VTAIL.n210 4.26717
R1069 VTAIL.n714 VTAIL.n622 4.26717
R1070 VTAIL.n685 VTAIL.n637 4.26717
R1071 VTAIL.n669 VTAIL.n668 4.26717
R1072 VTAIL.n610 VTAIL.n518 4.26717
R1073 VTAIL.n581 VTAIL.n533 4.26717
R1074 VTAIL.n565 VTAIL.n564 4.26717
R1075 VTAIL.n508 VTAIL.n416 4.26717
R1076 VTAIL.n479 VTAIL.n431 4.26717
R1077 VTAIL.n463 VTAIL.n462 4.26717
R1078 VTAIL.n404 VTAIL.n312 4.26717
R1079 VTAIL.n375 VTAIL.n327 4.26717
R1080 VTAIL.n359 VTAIL.n358 4.26717
R1081 VTAIL.n766 VTAIL.n748 3.49141
R1082 VTAIL.n790 VTAIL.n789 3.49141
R1083 VTAIL.n815 VTAIL.n726 3.49141
R1084 VTAIL.n46 VTAIL.n28 3.49141
R1085 VTAIL.n70 VTAIL.n69 3.49141
R1086 VTAIL.n95 VTAIL.n6 3.49141
R1087 VTAIL.n148 VTAIL.n130 3.49141
R1088 VTAIL.n172 VTAIL.n171 3.49141
R1089 VTAIL.n197 VTAIL.n108 3.49141
R1090 VTAIL.n252 VTAIL.n234 3.49141
R1091 VTAIL.n276 VTAIL.n275 3.49141
R1092 VTAIL.n301 VTAIL.n212 3.49141
R1093 VTAIL.n713 VTAIL.n624 3.49141
R1094 VTAIL.n689 VTAIL.n688 3.49141
R1095 VTAIL.n665 VTAIL.n647 3.49141
R1096 VTAIL.n609 VTAIL.n520 3.49141
R1097 VTAIL.n585 VTAIL.n584 3.49141
R1098 VTAIL.n561 VTAIL.n543 3.49141
R1099 VTAIL.n507 VTAIL.n418 3.49141
R1100 VTAIL.n483 VTAIL.n482 3.49141
R1101 VTAIL.n459 VTAIL.n441 3.49141
R1102 VTAIL.n403 VTAIL.n314 3.49141
R1103 VTAIL.n379 VTAIL.n378 3.49141
R1104 VTAIL.n355 VTAIL.n337 3.49141
R1105 VTAIL.n413 VTAIL.n411 3.40567
R1106 VTAIL.n515 VTAIL.n413 3.40567
R1107 VTAIL.n619 VTAIL.n617 3.40567
R1108 VTAIL.n721 VTAIL.n619 3.40567
R1109 VTAIL.n309 VTAIL.n207 3.40567
R1110 VTAIL.n207 VTAIL.n205 3.40567
R1111 VTAIL.n103 VTAIL.n1 3.40567
R1112 VTAIL VTAIL.n823 3.34748
R1113 VTAIL.n765 VTAIL.n750 2.71565
R1114 VTAIL.n793 VTAIL.n736 2.71565
R1115 VTAIL.n812 VTAIL.n811 2.71565
R1116 VTAIL.n45 VTAIL.n30 2.71565
R1117 VTAIL.n73 VTAIL.n16 2.71565
R1118 VTAIL.n92 VTAIL.n91 2.71565
R1119 VTAIL.n147 VTAIL.n132 2.71565
R1120 VTAIL.n175 VTAIL.n118 2.71565
R1121 VTAIL.n194 VTAIL.n193 2.71565
R1122 VTAIL.n251 VTAIL.n236 2.71565
R1123 VTAIL.n279 VTAIL.n222 2.71565
R1124 VTAIL.n298 VTAIL.n297 2.71565
R1125 VTAIL.n710 VTAIL.n709 2.71565
R1126 VTAIL.n692 VTAIL.n635 2.71565
R1127 VTAIL.n664 VTAIL.n649 2.71565
R1128 VTAIL.n606 VTAIL.n605 2.71565
R1129 VTAIL.n588 VTAIL.n531 2.71565
R1130 VTAIL.n560 VTAIL.n545 2.71565
R1131 VTAIL.n504 VTAIL.n503 2.71565
R1132 VTAIL.n486 VTAIL.n429 2.71565
R1133 VTAIL.n458 VTAIL.n443 2.71565
R1134 VTAIL.n400 VTAIL.n399 2.71565
R1135 VTAIL.n382 VTAIL.n325 2.71565
R1136 VTAIL.n354 VTAIL.n339 2.71565
R1137 VTAIL.n762 VTAIL.n761 1.93989
R1138 VTAIL.n794 VTAIL.n734 1.93989
R1139 VTAIL.n808 VTAIL.n728 1.93989
R1140 VTAIL.n42 VTAIL.n41 1.93989
R1141 VTAIL.n74 VTAIL.n14 1.93989
R1142 VTAIL.n88 VTAIL.n8 1.93989
R1143 VTAIL.n144 VTAIL.n143 1.93989
R1144 VTAIL.n176 VTAIL.n116 1.93989
R1145 VTAIL.n190 VTAIL.n110 1.93989
R1146 VTAIL.n248 VTAIL.n247 1.93989
R1147 VTAIL.n280 VTAIL.n220 1.93989
R1148 VTAIL.n294 VTAIL.n214 1.93989
R1149 VTAIL.n706 VTAIL.n626 1.93989
R1150 VTAIL.n693 VTAIL.n633 1.93989
R1151 VTAIL.n661 VTAIL.n660 1.93989
R1152 VTAIL.n602 VTAIL.n522 1.93989
R1153 VTAIL.n589 VTAIL.n529 1.93989
R1154 VTAIL.n557 VTAIL.n556 1.93989
R1155 VTAIL.n500 VTAIL.n420 1.93989
R1156 VTAIL.n487 VTAIL.n427 1.93989
R1157 VTAIL.n455 VTAIL.n454 1.93989
R1158 VTAIL.n396 VTAIL.n316 1.93989
R1159 VTAIL.n383 VTAIL.n323 1.93989
R1160 VTAIL.n351 VTAIL.n350 1.93989
R1161 VTAIL.n758 VTAIL.n752 1.16414
R1162 VTAIL.n799 VTAIL.n797 1.16414
R1163 VTAIL.n807 VTAIL.n730 1.16414
R1164 VTAIL.n38 VTAIL.n32 1.16414
R1165 VTAIL.n79 VTAIL.n77 1.16414
R1166 VTAIL.n87 VTAIL.n10 1.16414
R1167 VTAIL.n140 VTAIL.n134 1.16414
R1168 VTAIL.n181 VTAIL.n179 1.16414
R1169 VTAIL.n189 VTAIL.n112 1.16414
R1170 VTAIL.n244 VTAIL.n238 1.16414
R1171 VTAIL.n285 VTAIL.n283 1.16414
R1172 VTAIL.n293 VTAIL.n216 1.16414
R1173 VTAIL.n705 VTAIL.n628 1.16414
R1174 VTAIL.n697 VTAIL.n696 1.16414
R1175 VTAIL.n657 VTAIL.n651 1.16414
R1176 VTAIL.n601 VTAIL.n524 1.16414
R1177 VTAIL.n593 VTAIL.n592 1.16414
R1178 VTAIL.n553 VTAIL.n547 1.16414
R1179 VTAIL.n499 VTAIL.n422 1.16414
R1180 VTAIL.n491 VTAIL.n490 1.16414
R1181 VTAIL.n451 VTAIL.n445 1.16414
R1182 VTAIL.n395 VTAIL.n318 1.16414
R1183 VTAIL.n387 VTAIL.n386 1.16414
R1184 VTAIL.n347 VTAIL.n341 1.16414
R1185 VTAIL.n0 VTAIL.t0 1.09261
R1186 VTAIL.n0 VTAIL.t4 1.09261
R1187 VTAIL.n206 VTAIL.t11 1.09261
R1188 VTAIL.n206 VTAIL.t13 1.09261
R1189 VTAIL.n618 VTAIL.t12 1.09261
R1190 VTAIL.n618 VTAIL.t14 1.09261
R1191 VTAIL.n412 VTAIL.t1 1.09261
R1192 VTAIL.n412 VTAIL.t5 1.09261
R1193 VTAIL.n617 VTAIL.n515 0.470328
R1194 VTAIL.n205 VTAIL.n103 0.470328
R1195 VTAIL.n757 VTAIL.n754 0.388379
R1196 VTAIL.n798 VTAIL.n732 0.388379
R1197 VTAIL.n804 VTAIL.n803 0.388379
R1198 VTAIL.n37 VTAIL.n34 0.388379
R1199 VTAIL.n78 VTAIL.n12 0.388379
R1200 VTAIL.n84 VTAIL.n83 0.388379
R1201 VTAIL.n139 VTAIL.n136 0.388379
R1202 VTAIL.n180 VTAIL.n114 0.388379
R1203 VTAIL.n186 VTAIL.n185 0.388379
R1204 VTAIL.n243 VTAIL.n240 0.388379
R1205 VTAIL.n284 VTAIL.n218 0.388379
R1206 VTAIL.n290 VTAIL.n289 0.388379
R1207 VTAIL.n702 VTAIL.n701 0.388379
R1208 VTAIL.n632 VTAIL.n630 0.388379
R1209 VTAIL.n656 VTAIL.n653 0.388379
R1210 VTAIL.n598 VTAIL.n597 0.388379
R1211 VTAIL.n528 VTAIL.n526 0.388379
R1212 VTAIL.n552 VTAIL.n549 0.388379
R1213 VTAIL.n496 VTAIL.n495 0.388379
R1214 VTAIL.n426 VTAIL.n424 0.388379
R1215 VTAIL.n450 VTAIL.n447 0.388379
R1216 VTAIL.n392 VTAIL.n391 0.388379
R1217 VTAIL.n322 VTAIL.n320 0.388379
R1218 VTAIL.n346 VTAIL.n343 0.388379
R1219 VTAIL.n756 VTAIL.n751 0.155672
R1220 VTAIL.n763 VTAIL.n751 0.155672
R1221 VTAIL.n764 VTAIL.n763 0.155672
R1222 VTAIL.n764 VTAIL.n747 0.155672
R1223 VTAIL.n771 VTAIL.n747 0.155672
R1224 VTAIL.n772 VTAIL.n771 0.155672
R1225 VTAIL.n772 VTAIL.n743 0.155672
R1226 VTAIL.n779 VTAIL.n743 0.155672
R1227 VTAIL.n780 VTAIL.n779 0.155672
R1228 VTAIL.n780 VTAIL.n739 0.155672
R1229 VTAIL.n787 VTAIL.n739 0.155672
R1230 VTAIL.n788 VTAIL.n787 0.155672
R1231 VTAIL.n788 VTAIL.n735 0.155672
R1232 VTAIL.n795 VTAIL.n735 0.155672
R1233 VTAIL.n796 VTAIL.n795 0.155672
R1234 VTAIL.n796 VTAIL.n731 0.155672
R1235 VTAIL.n805 VTAIL.n731 0.155672
R1236 VTAIL.n806 VTAIL.n805 0.155672
R1237 VTAIL.n806 VTAIL.n727 0.155672
R1238 VTAIL.n813 VTAIL.n727 0.155672
R1239 VTAIL.n814 VTAIL.n813 0.155672
R1240 VTAIL.n814 VTAIL.n723 0.155672
R1241 VTAIL.n821 VTAIL.n723 0.155672
R1242 VTAIL.n36 VTAIL.n31 0.155672
R1243 VTAIL.n43 VTAIL.n31 0.155672
R1244 VTAIL.n44 VTAIL.n43 0.155672
R1245 VTAIL.n44 VTAIL.n27 0.155672
R1246 VTAIL.n51 VTAIL.n27 0.155672
R1247 VTAIL.n52 VTAIL.n51 0.155672
R1248 VTAIL.n52 VTAIL.n23 0.155672
R1249 VTAIL.n59 VTAIL.n23 0.155672
R1250 VTAIL.n60 VTAIL.n59 0.155672
R1251 VTAIL.n60 VTAIL.n19 0.155672
R1252 VTAIL.n67 VTAIL.n19 0.155672
R1253 VTAIL.n68 VTAIL.n67 0.155672
R1254 VTAIL.n68 VTAIL.n15 0.155672
R1255 VTAIL.n75 VTAIL.n15 0.155672
R1256 VTAIL.n76 VTAIL.n75 0.155672
R1257 VTAIL.n76 VTAIL.n11 0.155672
R1258 VTAIL.n85 VTAIL.n11 0.155672
R1259 VTAIL.n86 VTAIL.n85 0.155672
R1260 VTAIL.n86 VTAIL.n7 0.155672
R1261 VTAIL.n93 VTAIL.n7 0.155672
R1262 VTAIL.n94 VTAIL.n93 0.155672
R1263 VTAIL.n94 VTAIL.n3 0.155672
R1264 VTAIL.n101 VTAIL.n3 0.155672
R1265 VTAIL.n138 VTAIL.n133 0.155672
R1266 VTAIL.n145 VTAIL.n133 0.155672
R1267 VTAIL.n146 VTAIL.n145 0.155672
R1268 VTAIL.n146 VTAIL.n129 0.155672
R1269 VTAIL.n153 VTAIL.n129 0.155672
R1270 VTAIL.n154 VTAIL.n153 0.155672
R1271 VTAIL.n154 VTAIL.n125 0.155672
R1272 VTAIL.n161 VTAIL.n125 0.155672
R1273 VTAIL.n162 VTAIL.n161 0.155672
R1274 VTAIL.n162 VTAIL.n121 0.155672
R1275 VTAIL.n169 VTAIL.n121 0.155672
R1276 VTAIL.n170 VTAIL.n169 0.155672
R1277 VTAIL.n170 VTAIL.n117 0.155672
R1278 VTAIL.n177 VTAIL.n117 0.155672
R1279 VTAIL.n178 VTAIL.n177 0.155672
R1280 VTAIL.n178 VTAIL.n113 0.155672
R1281 VTAIL.n187 VTAIL.n113 0.155672
R1282 VTAIL.n188 VTAIL.n187 0.155672
R1283 VTAIL.n188 VTAIL.n109 0.155672
R1284 VTAIL.n195 VTAIL.n109 0.155672
R1285 VTAIL.n196 VTAIL.n195 0.155672
R1286 VTAIL.n196 VTAIL.n105 0.155672
R1287 VTAIL.n203 VTAIL.n105 0.155672
R1288 VTAIL.n242 VTAIL.n237 0.155672
R1289 VTAIL.n249 VTAIL.n237 0.155672
R1290 VTAIL.n250 VTAIL.n249 0.155672
R1291 VTAIL.n250 VTAIL.n233 0.155672
R1292 VTAIL.n257 VTAIL.n233 0.155672
R1293 VTAIL.n258 VTAIL.n257 0.155672
R1294 VTAIL.n258 VTAIL.n229 0.155672
R1295 VTAIL.n265 VTAIL.n229 0.155672
R1296 VTAIL.n266 VTAIL.n265 0.155672
R1297 VTAIL.n266 VTAIL.n225 0.155672
R1298 VTAIL.n273 VTAIL.n225 0.155672
R1299 VTAIL.n274 VTAIL.n273 0.155672
R1300 VTAIL.n274 VTAIL.n221 0.155672
R1301 VTAIL.n281 VTAIL.n221 0.155672
R1302 VTAIL.n282 VTAIL.n281 0.155672
R1303 VTAIL.n282 VTAIL.n217 0.155672
R1304 VTAIL.n291 VTAIL.n217 0.155672
R1305 VTAIL.n292 VTAIL.n291 0.155672
R1306 VTAIL.n292 VTAIL.n213 0.155672
R1307 VTAIL.n299 VTAIL.n213 0.155672
R1308 VTAIL.n300 VTAIL.n299 0.155672
R1309 VTAIL.n300 VTAIL.n209 0.155672
R1310 VTAIL.n307 VTAIL.n209 0.155672
R1311 VTAIL.n719 VTAIL.n621 0.155672
R1312 VTAIL.n712 VTAIL.n621 0.155672
R1313 VTAIL.n712 VTAIL.n711 0.155672
R1314 VTAIL.n711 VTAIL.n625 0.155672
R1315 VTAIL.n704 VTAIL.n625 0.155672
R1316 VTAIL.n704 VTAIL.n703 0.155672
R1317 VTAIL.n703 VTAIL.n629 0.155672
R1318 VTAIL.n695 VTAIL.n629 0.155672
R1319 VTAIL.n695 VTAIL.n694 0.155672
R1320 VTAIL.n694 VTAIL.n634 0.155672
R1321 VTAIL.n687 VTAIL.n634 0.155672
R1322 VTAIL.n687 VTAIL.n686 0.155672
R1323 VTAIL.n686 VTAIL.n638 0.155672
R1324 VTAIL.n679 VTAIL.n638 0.155672
R1325 VTAIL.n679 VTAIL.n678 0.155672
R1326 VTAIL.n678 VTAIL.n642 0.155672
R1327 VTAIL.n671 VTAIL.n642 0.155672
R1328 VTAIL.n671 VTAIL.n670 0.155672
R1329 VTAIL.n670 VTAIL.n646 0.155672
R1330 VTAIL.n663 VTAIL.n646 0.155672
R1331 VTAIL.n663 VTAIL.n662 0.155672
R1332 VTAIL.n662 VTAIL.n650 0.155672
R1333 VTAIL.n655 VTAIL.n650 0.155672
R1334 VTAIL.n615 VTAIL.n517 0.155672
R1335 VTAIL.n608 VTAIL.n517 0.155672
R1336 VTAIL.n608 VTAIL.n607 0.155672
R1337 VTAIL.n607 VTAIL.n521 0.155672
R1338 VTAIL.n600 VTAIL.n521 0.155672
R1339 VTAIL.n600 VTAIL.n599 0.155672
R1340 VTAIL.n599 VTAIL.n525 0.155672
R1341 VTAIL.n591 VTAIL.n525 0.155672
R1342 VTAIL.n591 VTAIL.n590 0.155672
R1343 VTAIL.n590 VTAIL.n530 0.155672
R1344 VTAIL.n583 VTAIL.n530 0.155672
R1345 VTAIL.n583 VTAIL.n582 0.155672
R1346 VTAIL.n582 VTAIL.n534 0.155672
R1347 VTAIL.n575 VTAIL.n534 0.155672
R1348 VTAIL.n575 VTAIL.n574 0.155672
R1349 VTAIL.n574 VTAIL.n538 0.155672
R1350 VTAIL.n567 VTAIL.n538 0.155672
R1351 VTAIL.n567 VTAIL.n566 0.155672
R1352 VTAIL.n566 VTAIL.n542 0.155672
R1353 VTAIL.n559 VTAIL.n542 0.155672
R1354 VTAIL.n559 VTAIL.n558 0.155672
R1355 VTAIL.n558 VTAIL.n546 0.155672
R1356 VTAIL.n551 VTAIL.n546 0.155672
R1357 VTAIL.n513 VTAIL.n415 0.155672
R1358 VTAIL.n506 VTAIL.n415 0.155672
R1359 VTAIL.n506 VTAIL.n505 0.155672
R1360 VTAIL.n505 VTAIL.n419 0.155672
R1361 VTAIL.n498 VTAIL.n419 0.155672
R1362 VTAIL.n498 VTAIL.n497 0.155672
R1363 VTAIL.n497 VTAIL.n423 0.155672
R1364 VTAIL.n489 VTAIL.n423 0.155672
R1365 VTAIL.n489 VTAIL.n488 0.155672
R1366 VTAIL.n488 VTAIL.n428 0.155672
R1367 VTAIL.n481 VTAIL.n428 0.155672
R1368 VTAIL.n481 VTAIL.n480 0.155672
R1369 VTAIL.n480 VTAIL.n432 0.155672
R1370 VTAIL.n473 VTAIL.n432 0.155672
R1371 VTAIL.n473 VTAIL.n472 0.155672
R1372 VTAIL.n472 VTAIL.n436 0.155672
R1373 VTAIL.n465 VTAIL.n436 0.155672
R1374 VTAIL.n465 VTAIL.n464 0.155672
R1375 VTAIL.n464 VTAIL.n440 0.155672
R1376 VTAIL.n457 VTAIL.n440 0.155672
R1377 VTAIL.n457 VTAIL.n456 0.155672
R1378 VTAIL.n456 VTAIL.n444 0.155672
R1379 VTAIL.n449 VTAIL.n444 0.155672
R1380 VTAIL.n409 VTAIL.n311 0.155672
R1381 VTAIL.n402 VTAIL.n311 0.155672
R1382 VTAIL.n402 VTAIL.n401 0.155672
R1383 VTAIL.n401 VTAIL.n315 0.155672
R1384 VTAIL.n394 VTAIL.n315 0.155672
R1385 VTAIL.n394 VTAIL.n393 0.155672
R1386 VTAIL.n393 VTAIL.n319 0.155672
R1387 VTAIL.n385 VTAIL.n319 0.155672
R1388 VTAIL.n385 VTAIL.n384 0.155672
R1389 VTAIL.n384 VTAIL.n324 0.155672
R1390 VTAIL.n377 VTAIL.n324 0.155672
R1391 VTAIL.n377 VTAIL.n376 0.155672
R1392 VTAIL.n376 VTAIL.n328 0.155672
R1393 VTAIL.n369 VTAIL.n328 0.155672
R1394 VTAIL.n369 VTAIL.n368 0.155672
R1395 VTAIL.n368 VTAIL.n332 0.155672
R1396 VTAIL.n361 VTAIL.n332 0.155672
R1397 VTAIL.n361 VTAIL.n360 0.155672
R1398 VTAIL.n360 VTAIL.n336 0.155672
R1399 VTAIL.n353 VTAIL.n336 0.155672
R1400 VTAIL.n353 VTAIL.n352 0.155672
R1401 VTAIL.n352 VTAIL.n340 0.155672
R1402 VTAIL.n345 VTAIL.n340 0.155672
R1403 VTAIL VTAIL.n1 0.0586897
R1404 B.n929 B.n189 585
R1405 B.n189 B.n120 585
R1406 B.n931 B.n930 585
R1407 B.n933 B.n188 585
R1408 B.n936 B.n935 585
R1409 B.n937 B.n187 585
R1410 B.n939 B.n938 585
R1411 B.n941 B.n186 585
R1412 B.n944 B.n943 585
R1413 B.n945 B.n185 585
R1414 B.n947 B.n946 585
R1415 B.n949 B.n184 585
R1416 B.n952 B.n951 585
R1417 B.n953 B.n183 585
R1418 B.n955 B.n954 585
R1419 B.n957 B.n182 585
R1420 B.n960 B.n959 585
R1421 B.n961 B.n181 585
R1422 B.n963 B.n962 585
R1423 B.n965 B.n180 585
R1424 B.n968 B.n967 585
R1425 B.n969 B.n179 585
R1426 B.n971 B.n970 585
R1427 B.n973 B.n178 585
R1428 B.n976 B.n975 585
R1429 B.n977 B.n177 585
R1430 B.n979 B.n978 585
R1431 B.n981 B.n176 585
R1432 B.n984 B.n983 585
R1433 B.n985 B.n175 585
R1434 B.n987 B.n986 585
R1435 B.n989 B.n174 585
R1436 B.n992 B.n991 585
R1437 B.n993 B.n173 585
R1438 B.n995 B.n994 585
R1439 B.n997 B.n172 585
R1440 B.n1000 B.n999 585
R1441 B.n1001 B.n171 585
R1442 B.n1003 B.n1002 585
R1443 B.n1005 B.n170 585
R1444 B.n1008 B.n1007 585
R1445 B.n1009 B.n169 585
R1446 B.n1011 B.n1010 585
R1447 B.n1013 B.n168 585
R1448 B.n1016 B.n1015 585
R1449 B.n1017 B.n167 585
R1450 B.n1019 B.n1018 585
R1451 B.n1021 B.n166 585
R1452 B.n1024 B.n1023 585
R1453 B.n1025 B.n165 585
R1454 B.n1027 B.n1026 585
R1455 B.n1029 B.n164 585
R1456 B.n1032 B.n1031 585
R1457 B.n1033 B.n163 585
R1458 B.n1035 B.n1034 585
R1459 B.n1037 B.n162 585
R1460 B.n1040 B.n1039 585
R1461 B.n1041 B.n161 585
R1462 B.n1043 B.n1042 585
R1463 B.n1045 B.n160 585
R1464 B.n1048 B.n1047 585
R1465 B.n1050 B.n157 585
R1466 B.n1052 B.n1051 585
R1467 B.n1054 B.n156 585
R1468 B.n1057 B.n1056 585
R1469 B.n1058 B.n155 585
R1470 B.n1060 B.n1059 585
R1471 B.n1062 B.n154 585
R1472 B.n1065 B.n1064 585
R1473 B.n1066 B.n151 585
R1474 B.n1069 B.n1068 585
R1475 B.n1071 B.n150 585
R1476 B.n1074 B.n1073 585
R1477 B.n1075 B.n149 585
R1478 B.n1077 B.n1076 585
R1479 B.n1079 B.n148 585
R1480 B.n1082 B.n1081 585
R1481 B.n1083 B.n147 585
R1482 B.n1085 B.n1084 585
R1483 B.n1087 B.n146 585
R1484 B.n1090 B.n1089 585
R1485 B.n1091 B.n145 585
R1486 B.n1093 B.n1092 585
R1487 B.n1095 B.n144 585
R1488 B.n1098 B.n1097 585
R1489 B.n1099 B.n143 585
R1490 B.n1101 B.n1100 585
R1491 B.n1103 B.n142 585
R1492 B.n1106 B.n1105 585
R1493 B.n1107 B.n141 585
R1494 B.n1109 B.n1108 585
R1495 B.n1111 B.n140 585
R1496 B.n1114 B.n1113 585
R1497 B.n1115 B.n139 585
R1498 B.n1117 B.n1116 585
R1499 B.n1119 B.n138 585
R1500 B.n1122 B.n1121 585
R1501 B.n1123 B.n137 585
R1502 B.n1125 B.n1124 585
R1503 B.n1127 B.n136 585
R1504 B.n1130 B.n1129 585
R1505 B.n1131 B.n135 585
R1506 B.n1133 B.n1132 585
R1507 B.n1135 B.n134 585
R1508 B.n1138 B.n1137 585
R1509 B.n1139 B.n133 585
R1510 B.n1141 B.n1140 585
R1511 B.n1143 B.n132 585
R1512 B.n1146 B.n1145 585
R1513 B.n1147 B.n131 585
R1514 B.n1149 B.n1148 585
R1515 B.n1151 B.n130 585
R1516 B.n1154 B.n1153 585
R1517 B.n1155 B.n129 585
R1518 B.n1157 B.n1156 585
R1519 B.n1159 B.n128 585
R1520 B.n1162 B.n1161 585
R1521 B.n1163 B.n127 585
R1522 B.n1165 B.n1164 585
R1523 B.n1167 B.n126 585
R1524 B.n1170 B.n1169 585
R1525 B.n1171 B.n125 585
R1526 B.n1173 B.n1172 585
R1527 B.n1175 B.n124 585
R1528 B.n1178 B.n1177 585
R1529 B.n1179 B.n123 585
R1530 B.n1181 B.n1180 585
R1531 B.n1183 B.n122 585
R1532 B.n1186 B.n1185 585
R1533 B.n1187 B.n121 585
R1534 B.n928 B.n119 585
R1535 B.n1190 B.n119 585
R1536 B.n927 B.n118 585
R1537 B.n1191 B.n118 585
R1538 B.n926 B.n117 585
R1539 B.n1192 B.n117 585
R1540 B.n925 B.n924 585
R1541 B.n924 B.n113 585
R1542 B.n923 B.n112 585
R1543 B.n1198 B.n112 585
R1544 B.n922 B.n111 585
R1545 B.n1199 B.n111 585
R1546 B.n921 B.n110 585
R1547 B.n1200 B.n110 585
R1548 B.n920 B.n919 585
R1549 B.n919 B.n106 585
R1550 B.n918 B.n105 585
R1551 B.n1206 B.n105 585
R1552 B.n917 B.n104 585
R1553 B.n1207 B.n104 585
R1554 B.n916 B.n103 585
R1555 B.n1208 B.n103 585
R1556 B.n915 B.n914 585
R1557 B.n914 B.n99 585
R1558 B.n913 B.n98 585
R1559 B.n1214 B.n98 585
R1560 B.n912 B.n97 585
R1561 B.n1215 B.n97 585
R1562 B.n911 B.n96 585
R1563 B.n1216 B.n96 585
R1564 B.n910 B.n909 585
R1565 B.n909 B.n92 585
R1566 B.n908 B.n91 585
R1567 B.n1222 B.n91 585
R1568 B.n907 B.n90 585
R1569 B.n1223 B.n90 585
R1570 B.n906 B.n89 585
R1571 B.n1224 B.n89 585
R1572 B.n905 B.n904 585
R1573 B.n904 B.n85 585
R1574 B.n903 B.n84 585
R1575 B.n1230 B.n84 585
R1576 B.n902 B.n83 585
R1577 B.n1231 B.n83 585
R1578 B.n901 B.n82 585
R1579 B.n1232 B.n82 585
R1580 B.n900 B.n899 585
R1581 B.n899 B.n81 585
R1582 B.n898 B.n77 585
R1583 B.n1238 B.n77 585
R1584 B.n897 B.n76 585
R1585 B.n1239 B.n76 585
R1586 B.n896 B.n75 585
R1587 B.n1240 B.n75 585
R1588 B.n895 B.n894 585
R1589 B.n894 B.n71 585
R1590 B.n893 B.n70 585
R1591 B.n1246 B.n70 585
R1592 B.n892 B.n69 585
R1593 B.n1247 B.n69 585
R1594 B.n891 B.n68 585
R1595 B.n1248 B.n68 585
R1596 B.n890 B.n889 585
R1597 B.n889 B.n64 585
R1598 B.n888 B.n63 585
R1599 B.n1254 B.n63 585
R1600 B.n887 B.n62 585
R1601 B.n1255 B.n62 585
R1602 B.n886 B.n61 585
R1603 B.n1256 B.n61 585
R1604 B.n885 B.n884 585
R1605 B.n884 B.n60 585
R1606 B.n883 B.n56 585
R1607 B.n1262 B.n56 585
R1608 B.n882 B.n55 585
R1609 B.n1263 B.n55 585
R1610 B.n881 B.n54 585
R1611 B.n1264 B.n54 585
R1612 B.n880 B.n879 585
R1613 B.n879 B.n50 585
R1614 B.n878 B.n49 585
R1615 B.n1270 B.n49 585
R1616 B.n877 B.n48 585
R1617 B.n1271 B.n48 585
R1618 B.n876 B.n47 585
R1619 B.n1272 B.n47 585
R1620 B.n875 B.n874 585
R1621 B.n874 B.n43 585
R1622 B.n873 B.n42 585
R1623 B.n1278 B.n42 585
R1624 B.n872 B.n41 585
R1625 B.n1279 B.n41 585
R1626 B.n871 B.n40 585
R1627 B.n1280 B.n40 585
R1628 B.n870 B.n869 585
R1629 B.n869 B.n36 585
R1630 B.n868 B.n35 585
R1631 B.n1286 B.n35 585
R1632 B.n867 B.n34 585
R1633 B.n1287 B.n34 585
R1634 B.n866 B.n33 585
R1635 B.n1288 B.n33 585
R1636 B.n865 B.n864 585
R1637 B.n864 B.n29 585
R1638 B.n863 B.n28 585
R1639 B.n1294 B.n28 585
R1640 B.n862 B.n27 585
R1641 B.n1295 B.n27 585
R1642 B.n861 B.n26 585
R1643 B.n1296 B.n26 585
R1644 B.n860 B.n859 585
R1645 B.n859 B.n22 585
R1646 B.n858 B.n21 585
R1647 B.n1302 B.n21 585
R1648 B.n857 B.n20 585
R1649 B.n1303 B.n20 585
R1650 B.n856 B.n19 585
R1651 B.n1304 B.n19 585
R1652 B.n855 B.n854 585
R1653 B.n854 B.n15 585
R1654 B.n853 B.n14 585
R1655 B.n1310 B.n14 585
R1656 B.n852 B.n13 585
R1657 B.n1311 B.n13 585
R1658 B.n851 B.n12 585
R1659 B.n1312 B.n12 585
R1660 B.n850 B.n849 585
R1661 B.n849 B.n8 585
R1662 B.n848 B.n7 585
R1663 B.n1318 B.n7 585
R1664 B.n847 B.n6 585
R1665 B.n1319 B.n6 585
R1666 B.n846 B.n5 585
R1667 B.n1320 B.n5 585
R1668 B.n845 B.n844 585
R1669 B.n844 B.n4 585
R1670 B.n843 B.n190 585
R1671 B.n843 B.n842 585
R1672 B.n833 B.n191 585
R1673 B.n192 B.n191 585
R1674 B.n835 B.n834 585
R1675 B.n836 B.n835 585
R1676 B.n832 B.n197 585
R1677 B.n197 B.n196 585
R1678 B.n831 B.n830 585
R1679 B.n830 B.n829 585
R1680 B.n199 B.n198 585
R1681 B.n200 B.n199 585
R1682 B.n822 B.n821 585
R1683 B.n823 B.n822 585
R1684 B.n820 B.n205 585
R1685 B.n205 B.n204 585
R1686 B.n819 B.n818 585
R1687 B.n818 B.n817 585
R1688 B.n207 B.n206 585
R1689 B.n208 B.n207 585
R1690 B.n810 B.n809 585
R1691 B.n811 B.n810 585
R1692 B.n808 B.n213 585
R1693 B.n213 B.n212 585
R1694 B.n807 B.n806 585
R1695 B.n806 B.n805 585
R1696 B.n215 B.n214 585
R1697 B.n216 B.n215 585
R1698 B.n798 B.n797 585
R1699 B.n799 B.n798 585
R1700 B.n796 B.n221 585
R1701 B.n221 B.n220 585
R1702 B.n795 B.n794 585
R1703 B.n794 B.n793 585
R1704 B.n223 B.n222 585
R1705 B.n224 B.n223 585
R1706 B.n786 B.n785 585
R1707 B.n787 B.n786 585
R1708 B.n784 B.n229 585
R1709 B.n229 B.n228 585
R1710 B.n783 B.n782 585
R1711 B.n782 B.n781 585
R1712 B.n231 B.n230 585
R1713 B.n232 B.n231 585
R1714 B.n774 B.n773 585
R1715 B.n775 B.n774 585
R1716 B.n772 B.n237 585
R1717 B.n237 B.n236 585
R1718 B.n771 B.n770 585
R1719 B.n770 B.n769 585
R1720 B.n239 B.n238 585
R1721 B.n240 B.n239 585
R1722 B.n762 B.n761 585
R1723 B.n763 B.n762 585
R1724 B.n760 B.n245 585
R1725 B.n245 B.n244 585
R1726 B.n759 B.n758 585
R1727 B.n758 B.n757 585
R1728 B.n247 B.n246 585
R1729 B.n750 B.n247 585
R1730 B.n749 B.n748 585
R1731 B.n751 B.n749 585
R1732 B.n747 B.n252 585
R1733 B.n252 B.n251 585
R1734 B.n746 B.n745 585
R1735 B.n745 B.n744 585
R1736 B.n254 B.n253 585
R1737 B.n255 B.n254 585
R1738 B.n737 B.n736 585
R1739 B.n738 B.n737 585
R1740 B.n735 B.n260 585
R1741 B.n260 B.n259 585
R1742 B.n734 B.n733 585
R1743 B.n733 B.n732 585
R1744 B.n262 B.n261 585
R1745 B.n263 B.n262 585
R1746 B.n725 B.n724 585
R1747 B.n726 B.n725 585
R1748 B.n723 B.n268 585
R1749 B.n268 B.n267 585
R1750 B.n722 B.n721 585
R1751 B.n721 B.n720 585
R1752 B.n270 B.n269 585
R1753 B.n713 B.n270 585
R1754 B.n712 B.n711 585
R1755 B.n714 B.n712 585
R1756 B.n710 B.n275 585
R1757 B.n275 B.n274 585
R1758 B.n709 B.n708 585
R1759 B.n708 B.n707 585
R1760 B.n277 B.n276 585
R1761 B.n278 B.n277 585
R1762 B.n700 B.n699 585
R1763 B.n701 B.n700 585
R1764 B.n698 B.n283 585
R1765 B.n283 B.n282 585
R1766 B.n697 B.n696 585
R1767 B.n696 B.n695 585
R1768 B.n285 B.n284 585
R1769 B.n286 B.n285 585
R1770 B.n688 B.n687 585
R1771 B.n689 B.n688 585
R1772 B.n686 B.n291 585
R1773 B.n291 B.n290 585
R1774 B.n685 B.n684 585
R1775 B.n684 B.n683 585
R1776 B.n293 B.n292 585
R1777 B.n294 B.n293 585
R1778 B.n676 B.n675 585
R1779 B.n677 B.n676 585
R1780 B.n674 B.n299 585
R1781 B.n299 B.n298 585
R1782 B.n673 B.n672 585
R1783 B.n672 B.n671 585
R1784 B.n301 B.n300 585
R1785 B.n302 B.n301 585
R1786 B.n664 B.n663 585
R1787 B.n665 B.n664 585
R1788 B.n662 B.n307 585
R1789 B.n307 B.n306 585
R1790 B.n661 B.n660 585
R1791 B.n660 B.n659 585
R1792 B.n309 B.n308 585
R1793 B.n310 B.n309 585
R1794 B.n652 B.n651 585
R1795 B.n653 B.n652 585
R1796 B.n650 B.n315 585
R1797 B.n315 B.n314 585
R1798 B.n649 B.n648 585
R1799 B.n648 B.n647 585
R1800 B.n644 B.n319 585
R1801 B.n643 B.n642 585
R1802 B.n640 B.n320 585
R1803 B.n640 B.n318 585
R1804 B.n639 B.n638 585
R1805 B.n637 B.n636 585
R1806 B.n635 B.n322 585
R1807 B.n633 B.n632 585
R1808 B.n631 B.n323 585
R1809 B.n630 B.n629 585
R1810 B.n627 B.n324 585
R1811 B.n625 B.n624 585
R1812 B.n623 B.n325 585
R1813 B.n622 B.n621 585
R1814 B.n619 B.n326 585
R1815 B.n617 B.n616 585
R1816 B.n615 B.n327 585
R1817 B.n614 B.n613 585
R1818 B.n611 B.n328 585
R1819 B.n609 B.n608 585
R1820 B.n607 B.n329 585
R1821 B.n606 B.n605 585
R1822 B.n603 B.n330 585
R1823 B.n601 B.n600 585
R1824 B.n599 B.n331 585
R1825 B.n598 B.n597 585
R1826 B.n595 B.n332 585
R1827 B.n593 B.n592 585
R1828 B.n591 B.n333 585
R1829 B.n590 B.n589 585
R1830 B.n587 B.n334 585
R1831 B.n585 B.n584 585
R1832 B.n583 B.n335 585
R1833 B.n582 B.n581 585
R1834 B.n579 B.n336 585
R1835 B.n577 B.n576 585
R1836 B.n575 B.n337 585
R1837 B.n574 B.n573 585
R1838 B.n571 B.n338 585
R1839 B.n569 B.n568 585
R1840 B.n567 B.n339 585
R1841 B.n566 B.n565 585
R1842 B.n563 B.n340 585
R1843 B.n561 B.n560 585
R1844 B.n559 B.n341 585
R1845 B.n558 B.n557 585
R1846 B.n555 B.n342 585
R1847 B.n553 B.n552 585
R1848 B.n551 B.n343 585
R1849 B.n550 B.n549 585
R1850 B.n547 B.n344 585
R1851 B.n545 B.n544 585
R1852 B.n543 B.n345 585
R1853 B.n542 B.n541 585
R1854 B.n539 B.n346 585
R1855 B.n537 B.n536 585
R1856 B.n535 B.n347 585
R1857 B.n534 B.n533 585
R1858 B.n531 B.n348 585
R1859 B.n529 B.n528 585
R1860 B.n527 B.n349 585
R1861 B.n525 B.n524 585
R1862 B.n522 B.n352 585
R1863 B.n520 B.n519 585
R1864 B.n518 B.n353 585
R1865 B.n517 B.n516 585
R1866 B.n514 B.n354 585
R1867 B.n512 B.n511 585
R1868 B.n510 B.n355 585
R1869 B.n509 B.n508 585
R1870 B.n506 B.n505 585
R1871 B.n504 B.n503 585
R1872 B.n502 B.n360 585
R1873 B.n500 B.n499 585
R1874 B.n498 B.n361 585
R1875 B.n497 B.n496 585
R1876 B.n494 B.n362 585
R1877 B.n492 B.n491 585
R1878 B.n490 B.n363 585
R1879 B.n489 B.n488 585
R1880 B.n486 B.n364 585
R1881 B.n484 B.n483 585
R1882 B.n482 B.n365 585
R1883 B.n481 B.n480 585
R1884 B.n478 B.n366 585
R1885 B.n476 B.n475 585
R1886 B.n474 B.n367 585
R1887 B.n473 B.n472 585
R1888 B.n470 B.n368 585
R1889 B.n468 B.n467 585
R1890 B.n466 B.n369 585
R1891 B.n465 B.n464 585
R1892 B.n462 B.n370 585
R1893 B.n460 B.n459 585
R1894 B.n458 B.n371 585
R1895 B.n457 B.n456 585
R1896 B.n454 B.n372 585
R1897 B.n452 B.n451 585
R1898 B.n450 B.n373 585
R1899 B.n449 B.n448 585
R1900 B.n446 B.n374 585
R1901 B.n444 B.n443 585
R1902 B.n442 B.n375 585
R1903 B.n441 B.n440 585
R1904 B.n438 B.n376 585
R1905 B.n436 B.n435 585
R1906 B.n434 B.n377 585
R1907 B.n433 B.n432 585
R1908 B.n430 B.n378 585
R1909 B.n428 B.n427 585
R1910 B.n426 B.n379 585
R1911 B.n425 B.n424 585
R1912 B.n422 B.n380 585
R1913 B.n420 B.n419 585
R1914 B.n418 B.n381 585
R1915 B.n417 B.n416 585
R1916 B.n414 B.n382 585
R1917 B.n412 B.n411 585
R1918 B.n410 B.n383 585
R1919 B.n409 B.n408 585
R1920 B.n406 B.n384 585
R1921 B.n404 B.n403 585
R1922 B.n402 B.n385 585
R1923 B.n401 B.n400 585
R1924 B.n398 B.n386 585
R1925 B.n396 B.n395 585
R1926 B.n394 B.n387 585
R1927 B.n393 B.n392 585
R1928 B.n390 B.n388 585
R1929 B.n317 B.n316 585
R1930 B.n646 B.n645 585
R1931 B.n647 B.n646 585
R1932 B.n313 B.n312 585
R1933 B.n314 B.n313 585
R1934 B.n655 B.n654 585
R1935 B.n654 B.n653 585
R1936 B.n656 B.n311 585
R1937 B.n311 B.n310 585
R1938 B.n658 B.n657 585
R1939 B.n659 B.n658 585
R1940 B.n305 B.n304 585
R1941 B.n306 B.n305 585
R1942 B.n667 B.n666 585
R1943 B.n666 B.n665 585
R1944 B.n668 B.n303 585
R1945 B.n303 B.n302 585
R1946 B.n670 B.n669 585
R1947 B.n671 B.n670 585
R1948 B.n297 B.n296 585
R1949 B.n298 B.n297 585
R1950 B.n679 B.n678 585
R1951 B.n678 B.n677 585
R1952 B.n680 B.n295 585
R1953 B.n295 B.n294 585
R1954 B.n682 B.n681 585
R1955 B.n683 B.n682 585
R1956 B.n289 B.n288 585
R1957 B.n290 B.n289 585
R1958 B.n691 B.n690 585
R1959 B.n690 B.n689 585
R1960 B.n692 B.n287 585
R1961 B.n287 B.n286 585
R1962 B.n694 B.n693 585
R1963 B.n695 B.n694 585
R1964 B.n281 B.n280 585
R1965 B.n282 B.n281 585
R1966 B.n703 B.n702 585
R1967 B.n702 B.n701 585
R1968 B.n704 B.n279 585
R1969 B.n279 B.n278 585
R1970 B.n706 B.n705 585
R1971 B.n707 B.n706 585
R1972 B.n273 B.n272 585
R1973 B.n274 B.n273 585
R1974 B.n716 B.n715 585
R1975 B.n715 B.n714 585
R1976 B.n717 B.n271 585
R1977 B.n713 B.n271 585
R1978 B.n719 B.n718 585
R1979 B.n720 B.n719 585
R1980 B.n266 B.n265 585
R1981 B.n267 B.n266 585
R1982 B.n728 B.n727 585
R1983 B.n727 B.n726 585
R1984 B.n729 B.n264 585
R1985 B.n264 B.n263 585
R1986 B.n731 B.n730 585
R1987 B.n732 B.n731 585
R1988 B.n258 B.n257 585
R1989 B.n259 B.n258 585
R1990 B.n740 B.n739 585
R1991 B.n739 B.n738 585
R1992 B.n741 B.n256 585
R1993 B.n256 B.n255 585
R1994 B.n743 B.n742 585
R1995 B.n744 B.n743 585
R1996 B.n250 B.n249 585
R1997 B.n251 B.n250 585
R1998 B.n753 B.n752 585
R1999 B.n752 B.n751 585
R2000 B.n754 B.n248 585
R2001 B.n750 B.n248 585
R2002 B.n756 B.n755 585
R2003 B.n757 B.n756 585
R2004 B.n243 B.n242 585
R2005 B.n244 B.n243 585
R2006 B.n765 B.n764 585
R2007 B.n764 B.n763 585
R2008 B.n766 B.n241 585
R2009 B.n241 B.n240 585
R2010 B.n768 B.n767 585
R2011 B.n769 B.n768 585
R2012 B.n235 B.n234 585
R2013 B.n236 B.n235 585
R2014 B.n777 B.n776 585
R2015 B.n776 B.n775 585
R2016 B.n778 B.n233 585
R2017 B.n233 B.n232 585
R2018 B.n780 B.n779 585
R2019 B.n781 B.n780 585
R2020 B.n227 B.n226 585
R2021 B.n228 B.n227 585
R2022 B.n789 B.n788 585
R2023 B.n788 B.n787 585
R2024 B.n790 B.n225 585
R2025 B.n225 B.n224 585
R2026 B.n792 B.n791 585
R2027 B.n793 B.n792 585
R2028 B.n219 B.n218 585
R2029 B.n220 B.n219 585
R2030 B.n801 B.n800 585
R2031 B.n800 B.n799 585
R2032 B.n802 B.n217 585
R2033 B.n217 B.n216 585
R2034 B.n804 B.n803 585
R2035 B.n805 B.n804 585
R2036 B.n211 B.n210 585
R2037 B.n212 B.n211 585
R2038 B.n813 B.n812 585
R2039 B.n812 B.n811 585
R2040 B.n814 B.n209 585
R2041 B.n209 B.n208 585
R2042 B.n816 B.n815 585
R2043 B.n817 B.n816 585
R2044 B.n203 B.n202 585
R2045 B.n204 B.n203 585
R2046 B.n825 B.n824 585
R2047 B.n824 B.n823 585
R2048 B.n826 B.n201 585
R2049 B.n201 B.n200 585
R2050 B.n828 B.n827 585
R2051 B.n829 B.n828 585
R2052 B.n195 B.n194 585
R2053 B.n196 B.n195 585
R2054 B.n838 B.n837 585
R2055 B.n837 B.n836 585
R2056 B.n839 B.n193 585
R2057 B.n193 B.n192 585
R2058 B.n841 B.n840 585
R2059 B.n842 B.n841 585
R2060 B.n2 B.n0 585
R2061 B.n4 B.n2 585
R2062 B.n3 B.n1 585
R2063 B.n1319 B.n3 585
R2064 B.n1317 B.n1316 585
R2065 B.n1318 B.n1317 585
R2066 B.n1315 B.n9 585
R2067 B.n9 B.n8 585
R2068 B.n1314 B.n1313 585
R2069 B.n1313 B.n1312 585
R2070 B.n11 B.n10 585
R2071 B.n1311 B.n11 585
R2072 B.n1309 B.n1308 585
R2073 B.n1310 B.n1309 585
R2074 B.n1307 B.n16 585
R2075 B.n16 B.n15 585
R2076 B.n1306 B.n1305 585
R2077 B.n1305 B.n1304 585
R2078 B.n18 B.n17 585
R2079 B.n1303 B.n18 585
R2080 B.n1301 B.n1300 585
R2081 B.n1302 B.n1301 585
R2082 B.n1299 B.n23 585
R2083 B.n23 B.n22 585
R2084 B.n1298 B.n1297 585
R2085 B.n1297 B.n1296 585
R2086 B.n25 B.n24 585
R2087 B.n1295 B.n25 585
R2088 B.n1293 B.n1292 585
R2089 B.n1294 B.n1293 585
R2090 B.n1291 B.n30 585
R2091 B.n30 B.n29 585
R2092 B.n1290 B.n1289 585
R2093 B.n1289 B.n1288 585
R2094 B.n32 B.n31 585
R2095 B.n1287 B.n32 585
R2096 B.n1285 B.n1284 585
R2097 B.n1286 B.n1285 585
R2098 B.n1283 B.n37 585
R2099 B.n37 B.n36 585
R2100 B.n1282 B.n1281 585
R2101 B.n1281 B.n1280 585
R2102 B.n39 B.n38 585
R2103 B.n1279 B.n39 585
R2104 B.n1277 B.n1276 585
R2105 B.n1278 B.n1277 585
R2106 B.n1275 B.n44 585
R2107 B.n44 B.n43 585
R2108 B.n1274 B.n1273 585
R2109 B.n1273 B.n1272 585
R2110 B.n46 B.n45 585
R2111 B.n1271 B.n46 585
R2112 B.n1269 B.n1268 585
R2113 B.n1270 B.n1269 585
R2114 B.n1267 B.n51 585
R2115 B.n51 B.n50 585
R2116 B.n1266 B.n1265 585
R2117 B.n1265 B.n1264 585
R2118 B.n53 B.n52 585
R2119 B.n1263 B.n53 585
R2120 B.n1261 B.n1260 585
R2121 B.n1262 B.n1261 585
R2122 B.n1259 B.n57 585
R2123 B.n60 B.n57 585
R2124 B.n1258 B.n1257 585
R2125 B.n1257 B.n1256 585
R2126 B.n59 B.n58 585
R2127 B.n1255 B.n59 585
R2128 B.n1253 B.n1252 585
R2129 B.n1254 B.n1253 585
R2130 B.n1251 B.n65 585
R2131 B.n65 B.n64 585
R2132 B.n1250 B.n1249 585
R2133 B.n1249 B.n1248 585
R2134 B.n67 B.n66 585
R2135 B.n1247 B.n67 585
R2136 B.n1245 B.n1244 585
R2137 B.n1246 B.n1245 585
R2138 B.n1243 B.n72 585
R2139 B.n72 B.n71 585
R2140 B.n1242 B.n1241 585
R2141 B.n1241 B.n1240 585
R2142 B.n74 B.n73 585
R2143 B.n1239 B.n74 585
R2144 B.n1237 B.n1236 585
R2145 B.n1238 B.n1237 585
R2146 B.n1235 B.n78 585
R2147 B.n81 B.n78 585
R2148 B.n1234 B.n1233 585
R2149 B.n1233 B.n1232 585
R2150 B.n80 B.n79 585
R2151 B.n1231 B.n80 585
R2152 B.n1229 B.n1228 585
R2153 B.n1230 B.n1229 585
R2154 B.n1227 B.n86 585
R2155 B.n86 B.n85 585
R2156 B.n1226 B.n1225 585
R2157 B.n1225 B.n1224 585
R2158 B.n88 B.n87 585
R2159 B.n1223 B.n88 585
R2160 B.n1221 B.n1220 585
R2161 B.n1222 B.n1221 585
R2162 B.n1219 B.n93 585
R2163 B.n93 B.n92 585
R2164 B.n1218 B.n1217 585
R2165 B.n1217 B.n1216 585
R2166 B.n95 B.n94 585
R2167 B.n1215 B.n95 585
R2168 B.n1213 B.n1212 585
R2169 B.n1214 B.n1213 585
R2170 B.n1211 B.n100 585
R2171 B.n100 B.n99 585
R2172 B.n1210 B.n1209 585
R2173 B.n1209 B.n1208 585
R2174 B.n102 B.n101 585
R2175 B.n1207 B.n102 585
R2176 B.n1205 B.n1204 585
R2177 B.n1206 B.n1205 585
R2178 B.n1203 B.n107 585
R2179 B.n107 B.n106 585
R2180 B.n1202 B.n1201 585
R2181 B.n1201 B.n1200 585
R2182 B.n109 B.n108 585
R2183 B.n1199 B.n109 585
R2184 B.n1197 B.n1196 585
R2185 B.n1198 B.n1197 585
R2186 B.n1195 B.n114 585
R2187 B.n114 B.n113 585
R2188 B.n1194 B.n1193 585
R2189 B.n1193 B.n1192 585
R2190 B.n116 B.n115 585
R2191 B.n1191 B.n116 585
R2192 B.n1189 B.n1188 585
R2193 B.n1190 B.n1189 585
R2194 B.n1322 B.n1321 585
R2195 B.n1321 B.n1320 585
R2196 B.n646 B.n319 521.33
R2197 B.n1189 B.n121 521.33
R2198 B.n648 B.n317 521.33
R2199 B.n189 B.n119 521.33
R2200 B.n356 B.t17 464.219
R2201 B.n158 B.t12 464.219
R2202 B.n350 B.t20 464.219
R2203 B.n152 B.t9 464.219
R2204 B.n357 B.t16 387.613
R2205 B.n159 B.t13 387.613
R2206 B.n351 B.t19 387.613
R2207 B.n153 B.t10 387.613
R2208 B.n356 B.t14 329.899
R2209 B.n350 B.t18 329.899
R2210 B.n152 B.t7 329.899
R2211 B.n158 B.t11 329.899
R2212 B.n932 B.n120 256.663
R2213 B.n934 B.n120 256.663
R2214 B.n940 B.n120 256.663
R2215 B.n942 B.n120 256.663
R2216 B.n948 B.n120 256.663
R2217 B.n950 B.n120 256.663
R2218 B.n956 B.n120 256.663
R2219 B.n958 B.n120 256.663
R2220 B.n964 B.n120 256.663
R2221 B.n966 B.n120 256.663
R2222 B.n972 B.n120 256.663
R2223 B.n974 B.n120 256.663
R2224 B.n980 B.n120 256.663
R2225 B.n982 B.n120 256.663
R2226 B.n988 B.n120 256.663
R2227 B.n990 B.n120 256.663
R2228 B.n996 B.n120 256.663
R2229 B.n998 B.n120 256.663
R2230 B.n1004 B.n120 256.663
R2231 B.n1006 B.n120 256.663
R2232 B.n1012 B.n120 256.663
R2233 B.n1014 B.n120 256.663
R2234 B.n1020 B.n120 256.663
R2235 B.n1022 B.n120 256.663
R2236 B.n1028 B.n120 256.663
R2237 B.n1030 B.n120 256.663
R2238 B.n1036 B.n120 256.663
R2239 B.n1038 B.n120 256.663
R2240 B.n1044 B.n120 256.663
R2241 B.n1046 B.n120 256.663
R2242 B.n1053 B.n120 256.663
R2243 B.n1055 B.n120 256.663
R2244 B.n1061 B.n120 256.663
R2245 B.n1063 B.n120 256.663
R2246 B.n1070 B.n120 256.663
R2247 B.n1072 B.n120 256.663
R2248 B.n1078 B.n120 256.663
R2249 B.n1080 B.n120 256.663
R2250 B.n1086 B.n120 256.663
R2251 B.n1088 B.n120 256.663
R2252 B.n1094 B.n120 256.663
R2253 B.n1096 B.n120 256.663
R2254 B.n1102 B.n120 256.663
R2255 B.n1104 B.n120 256.663
R2256 B.n1110 B.n120 256.663
R2257 B.n1112 B.n120 256.663
R2258 B.n1118 B.n120 256.663
R2259 B.n1120 B.n120 256.663
R2260 B.n1126 B.n120 256.663
R2261 B.n1128 B.n120 256.663
R2262 B.n1134 B.n120 256.663
R2263 B.n1136 B.n120 256.663
R2264 B.n1142 B.n120 256.663
R2265 B.n1144 B.n120 256.663
R2266 B.n1150 B.n120 256.663
R2267 B.n1152 B.n120 256.663
R2268 B.n1158 B.n120 256.663
R2269 B.n1160 B.n120 256.663
R2270 B.n1166 B.n120 256.663
R2271 B.n1168 B.n120 256.663
R2272 B.n1174 B.n120 256.663
R2273 B.n1176 B.n120 256.663
R2274 B.n1182 B.n120 256.663
R2275 B.n1184 B.n120 256.663
R2276 B.n641 B.n318 256.663
R2277 B.n321 B.n318 256.663
R2278 B.n634 B.n318 256.663
R2279 B.n628 B.n318 256.663
R2280 B.n626 B.n318 256.663
R2281 B.n620 B.n318 256.663
R2282 B.n618 B.n318 256.663
R2283 B.n612 B.n318 256.663
R2284 B.n610 B.n318 256.663
R2285 B.n604 B.n318 256.663
R2286 B.n602 B.n318 256.663
R2287 B.n596 B.n318 256.663
R2288 B.n594 B.n318 256.663
R2289 B.n588 B.n318 256.663
R2290 B.n586 B.n318 256.663
R2291 B.n580 B.n318 256.663
R2292 B.n578 B.n318 256.663
R2293 B.n572 B.n318 256.663
R2294 B.n570 B.n318 256.663
R2295 B.n564 B.n318 256.663
R2296 B.n562 B.n318 256.663
R2297 B.n556 B.n318 256.663
R2298 B.n554 B.n318 256.663
R2299 B.n548 B.n318 256.663
R2300 B.n546 B.n318 256.663
R2301 B.n540 B.n318 256.663
R2302 B.n538 B.n318 256.663
R2303 B.n532 B.n318 256.663
R2304 B.n530 B.n318 256.663
R2305 B.n523 B.n318 256.663
R2306 B.n521 B.n318 256.663
R2307 B.n515 B.n318 256.663
R2308 B.n513 B.n318 256.663
R2309 B.n507 B.n318 256.663
R2310 B.n359 B.n318 256.663
R2311 B.n501 B.n318 256.663
R2312 B.n495 B.n318 256.663
R2313 B.n493 B.n318 256.663
R2314 B.n487 B.n318 256.663
R2315 B.n485 B.n318 256.663
R2316 B.n479 B.n318 256.663
R2317 B.n477 B.n318 256.663
R2318 B.n471 B.n318 256.663
R2319 B.n469 B.n318 256.663
R2320 B.n463 B.n318 256.663
R2321 B.n461 B.n318 256.663
R2322 B.n455 B.n318 256.663
R2323 B.n453 B.n318 256.663
R2324 B.n447 B.n318 256.663
R2325 B.n445 B.n318 256.663
R2326 B.n439 B.n318 256.663
R2327 B.n437 B.n318 256.663
R2328 B.n431 B.n318 256.663
R2329 B.n429 B.n318 256.663
R2330 B.n423 B.n318 256.663
R2331 B.n421 B.n318 256.663
R2332 B.n415 B.n318 256.663
R2333 B.n413 B.n318 256.663
R2334 B.n407 B.n318 256.663
R2335 B.n405 B.n318 256.663
R2336 B.n399 B.n318 256.663
R2337 B.n397 B.n318 256.663
R2338 B.n391 B.n318 256.663
R2339 B.n389 B.n318 256.663
R2340 B.n646 B.n313 163.367
R2341 B.n654 B.n313 163.367
R2342 B.n654 B.n311 163.367
R2343 B.n658 B.n311 163.367
R2344 B.n658 B.n305 163.367
R2345 B.n666 B.n305 163.367
R2346 B.n666 B.n303 163.367
R2347 B.n670 B.n303 163.367
R2348 B.n670 B.n297 163.367
R2349 B.n678 B.n297 163.367
R2350 B.n678 B.n295 163.367
R2351 B.n682 B.n295 163.367
R2352 B.n682 B.n289 163.367
R2353 B.n690 B.n289 163.367
R2354 B.n690 B.n287 163.367
R2355 B.n694 B.n287 163.367
R2356 B.n694 B.n281 163.367
R2357 B.n702 B.n281 163.367
R2358 B.n702 B.n279 163.367
R2359 B.n706 B.n279 163.367
R2360 B.n706 B.n273 163.367
R2361 B.n715 B.n273 163.367
R2362 B.n715 B.n271 163.367
R2363 B.n719 B.n271 163.367
R2364 B.n719 B.n266 163.367
R2365 B.n727 B.n266 163.367
R2366 B.n727 B.n264 163.367
R2367 B.n731 B.n264 163.367
R2368 B.n731 B.n258 163.367
R2369 B.n739 B.n258 163.367
R2370 B.n739 B.n256 163.367
R2371 B.n743 B.n256 163.367
R2372 B.n743 B.n250 163.367
R2373 B.n752 B.n250 163.367
R2374 B.n752 B.n248 163.367
R2375 B.n756 B.n248 163.367
R2376 B.n756 B.n243 163.367
R2377 B.n764 B.n243 163.367
R2378 B.n764 B.n241 163.367
R2379 B.n768 B.n241 163.367
R2380 B.n768 B.n235 163.367
R2381 B.n776 B.n235 163.367
R2382 B.n776 B.n233 163.367
R2383 B.n780 B.n233 163.367
R2384 B.n780 B.n227 163.367
R2385 B.n788 B.n227 163.367
R2386 B.n788 B.n225 163.367
R2387 B.n792 B.n225 163.367
R2388 B.n792 B.n219 163.367
R2389 B.n800 B.n219 163.367
R2390 B.n800 B.n217 163.367
R2391 B.n804 B.n217 163.367
R2392 B.n804 B.n211 163.367
R2393 B.n812 B.n211 163.367
R2394 B.n812 B.n209 163.367
R2395 B.n816 B.n209 163.367
R2396 B.n816 B.n203 163.367
R2397 B.n824 B.n203 163.367
R2398 B.n824 B.n201 163.367
R2399 B.n828 B.n201 163.367
R2400 B.n828 B.n195 163.367
R2401 B.n837 B.n195 163.367
R2402 B.n837 B.n193 163.367
R2403 B.n841 B.n193 163.367
R2404 B.n841 B.n2 163.367
R2405 B.n1321 B.n2 163.367
R2406 B.n1321 B.n3 163.367
R2407 B.n1317 B.n3 163.367
R2408 B.n1317 B.n9 163.367
R2409 B.n1313 B.n9 163.367
R2410 B.n1313 B.n11 163.367
R2411 B.n1309 B.n11 163.367
R2412 B.n1309 B.n16 163.367
R2413 B.n1305 B.n16 163.367
R2414 B.n1305 B.n18 163.367
R2415 B.n1301 B.n18 163.367
R2416 B.n1301 B.n23 163.367
R2417 B.n1297 B.n23 163.367
R2418 B.n1297 B.n25 163.367
R2419 B.n1293 B.n25 163.367
R2420 B.n1293 B.n30 163.367
R2421 B.n1289 B.n30 163.367
R2422 B.n1289 B.n32 163.367
R2423 B.n1285 B.n32 163.367
R2424 B.n1285 B.n37 163.367
R2425 B.n1281 B.n37 163.367
R2426 B.n1281 B.n39 163.367
R2427 B.n1277 B.n39 163.367
R2428 B.n1277 B.n44 163.367
R2429 B.n1273 B.n44 163.367
R2430 B.n1273 B.n46 163.367
R2431 B.n1269 B.n46 163.367
R2432 B.n1269 B.n51 163.367
R2433 B.n1265 B.n51 163.367
R2434 B.n1265 B.n53 163.367
R2435 B.n1261 B.n53 163.367
R2436 B.n1261 B.n57 163.367
R2437 B.n1257 B.n57 163.367
R2438 B.n1257 B.n59 163.367
R2439 B.n1253 B.n59 163.367
R2440 B.n1253 B.n65 163.367
R2441 B.n1249 B.n65 163.367
R2442 B.n1249 B.n67 163.367
R2443 B.n1245 B.n67 163.367
R2444 B.n1245 B.n72 163.367
R2445 B.n1241 B.n72 163.367
R2446 B.n1241 B.n74 163.367
R2447 B.n1237 B.n74 163.367
R2448 B.n1237 B.n78 163.367
R2449 B.n1233 B.n78 163.367
R2450 B.n1233 B.n80 163.367
R2451 B.n1229 B.n80 163.367
R2452 B.n1229 B.n86 163.367
R2453 B.n1225 B.n86 163.367
R2454 B.n1225 B.n88 163.367
R2455 B.n1221 B.n88 163.367
R2456 B.n1221 B.n93 163.367
R2457 B.n1217 B.n93 163.367
R2458 B.n1217 B.n95 163.367
R2459 B.n1213 B.n95 163.367
R2460 B.n1213 B.n100 163.367
R2461 B.n1209 B.n100 163.367
R2462 B.n1209 B.n102 163.367
R2463 B.n1205 B.n102 163.367
R2464 B.n1205 B.n107 163.367
R2465 B.n1201 B.n107 163.367
R2466 B.n1201 B.n109 163.367
R2467 B.n1197 B.n109 163.367
R2468 B.n1197 B.n114 163.367
R2469 B.n1193 B.n114 163.367
R2470 B.n1193 B.n116 163.367
R2471 B.n1189 B.n116 163.367
R2472 B.n642 B.n640 163.367
R2473 B.n640 B.n639 163.367
R2474 B.n636 B.n635 163.367
R2475 B.n633 B.n323 163.367
R2476 B.n629 B.n627 163.367
R2477 B.n625 B.n325 163.367
R2478 B.n621 B.n619 163.367
R2479 B.n617 B.n327 163.367
R2480 B.n613 B.n611 163.367
R2481 B.n609 B.n329 163.367
R2482 B.n605 B.n603 163.367
R2483 B.n601 B.n331 163.367
R2484 B.n597 B.n595 163.367
R2485 B.n593 B.n333 163.367
R2486 B.n589 B.n587 163.367
R2487 B.n585 B.n335 163.367
R2488 B.n581 B.n579 163.367
R2489 B.n577 B.n337 163.367
R2490 B.n573 B.n571 163.367
R2491 B.n569 B.n339 163.367
R2492 B.n565 B.n563 163.367
R2493 B.n561 B.n341 163.367
R2494 B.n557 B.n555 163.367
R2495 B.n553 B.n343 163.367
R2496 B.n549 B.n547 163.367
R2497 B.n545 B.n345 163.367
R2498 B.n541 B.n539 163.367
R2499 B.n537 B.n347 163.367
R2500 B.n533 B.n531 163.367
R2501 B.n529 B.n349 163.367
R2502 B.n524 B.n522 163.367
R2503 B.n520 B.n353 163.367
R2504 B.n516 B.n514 163.367
R2505 B.n512 B.n355 163.367
R2506 B.n508 B.n506 163.367
R2507 B.n503 B.n502 163.367
R2508 B.n500 B.n361 163.367
R2509 B.n496 B.n494 163.367
R2510 B.n492 B.n363 163.367
R2511 B.n488 B.n486 163.367
R2512 B.n484 B.n365 163.367
R2513 B.n480 B.n478 163.367
R2514 B.n476 B.n367 163.367
R2515 B.n472 B.n470 163.367
R2516 B.n468 B.n369 163.367
R2517 B.n464 B.n462 163.367
R2518 B.n460 B.n371 163.367
R2519 B.n456 B.n454 163.367
R2520 B.n452 B.n373 163.367
R2521 B.n448 B.n446 163.367
R2522 B.n444 B.n375 163.367
R2523 B.n440 B.n438 163.367
R2524 B.n436 B.n377 163.367
R2525 B.n432 B.n430 163.367
R2526 B.n428 B.n379 163.367
R2527 B.n424 B.n422 163.367
R2528 B.n420 B.n381 163.367
R2529 B.n416 B.n414 163.367
R2530 B.n412 B.n383 163.367
R2531 B.n408 B.n406 163.367
R2532 B.n404 B.n385 163.367
R2533 B.n400 B.n398 163.367
R2534 B.n396 B.n387 163.367
R2535 B.n392 B.n390 163.367
R2536 B.n648 B.n315 163.367
R2537 B.n652 B.n315 163.367
R2538 B.n652 B.n309 163.367
R2539 B.n660 B.n309 163.367
R2540 B.n660 B.n307 163.367
R2541 B.n664 B.n307 163.367
R2542 B.n664 B.n301 163.367
R2543 B.n672 B.n301 163.367
R2544 B.n672 B.n299 163.367
R2545 B.n676 B.n299 163.367
R2546 B.n676 B.n293 163.367
R2547 B.n684 B.n293 163.367
R2548 B.n684 B.n291 163.367
R2549 B.n688 B.n291 163.367
R2550 B.n688 B.n285 163.367
R2551 B.n696 B.n285 163.367
R2552 B.n696 B.n283 163.367
R2553 B.n700 B.n283 163.367
R2554 B.n700 B.n277 163.367
R2555 B.n708 B.n277 163.367
R2556 B.n708 B.n275 163.367
R2557 B.n712 B.n275 163.367
R2558 B.n712 B.n270 163.367
R2559 B.n721 B.n270 163.367
R2560 B.n721 B.n268 163.367
R2561 B.n725 B.n268 163.367
R2562 B.n725 B.n262 163.367
R2563 B.n733 B.n262 163.367
R2564 B.n733 B.n260 163.367
R2565 B.n737 B.n260 163.367
R2566 B.n737 B.n254 163.367
R2567 B.n745 B.n254 163.367
R2568 B.n745 B.n252 163.367
R2569 B.n749 B.n252 163.367
R2570 B.n749 B.n247 163.367
R2571 B.n758 B.n247 163.367
R2572 B.n758 B.n245 163.367
R2573 B.n762 B.n245 163.367
R2574 B.n762 B.n239 163.367
R2575 B.n770 B.n239 163.367
R2576 B.n770 B.n237 163.367
R2577 B.n774 B.n237 163.367
R2578 B.n774 B.n231 163.367
R2579 B.n782 B.n231 163.367
R2580 B.n782 B.n229 163.367
R2581 B.n786 B.n229 163.367
R2582 B.n786 B.n223 163.367
R2583 B.n794 B.n223 163.367
R2584 B.n794 B.n221 163.367
R2585 B.n798 B.n221 163.367
R2586 B.n798 B.n215 163.367
R2587 B.n806 B.n215 163.367
R2588 B.n806 B.n213 163.367
R2589 B.n810 B.n213 163.367
R2590 B.n810 B.n207 163.367
R2591 B.n818 B.n207 163.367
R2592 B.n818 B.n205 163.367
R2593 B.n822 B.n205 163.367
R2594 B.n822 B.n199 163.367
R2595 B.n830 B.n199 163.367
R2596 B.n830 B.n197 163.367
R2597 B.n835 B.n197 163.367
R2598 B.n835 B.n191 163.367
R2599 B.n843 B.n191 163.367
R2600 B.n844 B.n843 163.367
R2601 B.n844 B.n5 163.367
R2602 B.n6 B.n5 163.367
R2603 B.n7 B.n6 163.367
R2604 B.n849 B.n7 163.367
R2605 B.n849 B.n12 163.367
R2606 B.n13 B.n12 163.367
R2607 B.n14 B.n13 163.367
R2608 B.n854 B.n14 163.367
R2609 B.n854 B.n19 163.367
R2610 B.n20 B.n19 163.367
R2611 B.n21 B.n20 163.367
R2612 B.n859 B.n21 163.367
R2613 B.n859 B.n26 163.367
R2614 B.n27 B.n26 163.367
R2615 B.n28 B.n27 163.367
R2616 B.n864 B.n28 163.367
R2617 B.n864 B.n33 163.367
R2618 B.n34 B.n33 163.367
R2619 B.n35 B.n34 163.367
R2620 B.n869 B.n35 163.367
R2621 B.n869 B.n40 163.367
R2622 B.n41 B.n40 163.367
R2623 B.n42 B.n41 163.367
R2624 B.n874 B.n42 163.367
R2625 B.n874 B.n47 163.367
R2626 B.n48 B.n47 163.367
R2627 B.n49 B.n48 163.367
R2628 B.n879 B.n49 163.367
R2629 B.n879 B.n54 163.367
R2630 B.n55 B.n54 163.367
R2631 B.n56 B.n55 163.367
R2632 B.n884 B.n56 163.367
R2633 B.n884 B.n61 163.367
R2634 B.n62 B.n61 163.367
R2635 B.n63 B.n62 163.367
R2636 B.n889 B.n63 163.367
R2637 B.n889 B.n68 163.367
R2638 B.n69 B.n68 163.367
R2639 B.n70 B.n69 163.367
R2640 B.n894 B.n70 163.367
R2641 B.n894 B.n75 163.367
R2642 B.n76 B.n75 163.367
R2643 B.n77 B.n76 163.367
R2644 B.n899 B.n77 163.367
R2645 B.n899 B.n82 163.367
R2646 B.n83 B.n82 163.367
R2647 B.n84 B.n83 163.367
R2648 B.n904 B.n84 163.367
R2649 B.n904 B.n89 163.367
R2650 B.n90 B.n89 163.367
R2651 B.n91 B.n90 163.367
R2652 B.n909 B.n91 163.367
R2653 B.n909 B.n96 163.367
R2654 B.n97 B.n96 163.367
R2655 B.n98 B.n97 163.367
R2656 B.n914 B.n98 163.367
R2657 B.n914 B.n103 163.367
R2658 B.n104 B.n103 163.367
R2659 B.n105 B.n104 163.367
R2660 B.n919 B.n105 163.367
R2661 B.n919 B.n110 163.367
R2662 B.n111 B.n110 163.367
R2663 B.n112 B.n111 163.367
R2664 B.n924 B.n112 163.367
R2665 B.n924 B.n117 163.367
R2666 B.n118 B.n117 163.367
R2667 B.n119 B.n118 163.367
R2668 B.n1185 B.n1183 163.367
R2669 B.n1181 B.n123 163.367
R2670 B.n1177 B.n1175 163.367
R2671 B.n1173 B.n125 163.367
R2672 B.n1169 B.n1167 163.367
R2673 B.n1165 B.n127 163.367
R2674 B.n1161 B.n1159 163.367
R2675 B.n1157 B.n129 163.367
R2676 B.n1153 B.n1151 163.367
R2677 B.n1149 B.n131 163.367
R2678 B.n1145 B.n1143 163.367
R2679 B.n1141 B.n133 163.367
R2680 B.n1137 B.n1135 163.367
R2681 B.n1133 B.n135 163.367
R2682 B.n1129 B.n1127 163.367
R2683 B.n1125 B.n137 163.367
R2684 B.n1121 B.n1119 163.367
R2685 B.n1117 B.n139 163.367
R2686 B.n1113 B.n1111 163.367
R2687 B.n1109 B.n141 163.367
R2688 B.n1105 B.n1103 163.367
R2689 B.n1101 B.n143 163.367
R2690 B.n1097 B.n1095 163.367
R2691 B.n1093 B.n145 163.367
R2692 B.n1089 B.n1087 163.367
R2693 B.n1085 B.n147 163.367
R2694 B.n1081 B.n1079 163.367
R2695 B.n1077 B.n149 163.367
R2696 B.n1073 B.n1071 163.367
R2697 B.n1069 B.n151 163.367
R2698 B.n1064 B.n1062 163.367
R2699 B.n1060 B.n155 163.367
R2700 B.n1056 B.n1054 163.367
R2701 B.n1052 B.n157 163.367
R2702 B.n1047 B.n1045 163.367
R2703 B.n1043 B.n161 163.367
R2704 B.n1039 B.n1037 163.367
R2705 B.n1035 B.n163 163.367
R2706 B.n1031 B.n1029 163.367
R2707 B.n1027 B.n165 163.367
R2708 B.n1023 B.n1021 163.367
R2709 B.n1019 B.n167 163.367
R2710 B.n1015 B.n1013 163.367
R2711 B.n1011 B.n169 163.367
R2712 B.n1007 B.n1005 163.367
R2713 B.n1003 B.n171 163.367
R2714 B.n999 B.n997 163.367
R2715 B.n995 B.n173 163.367
R2716 B.n991 B.n989 163.367
R2717 B.n987 B.n175 163.367
R2718 B.n983 B.n981 163.367
R2719 B.n979 B.n177 163.367
R2720 B.n975 B.n973 163.367
R2721 B.n971 B.n179 163.367
R2722 B.n967 B.n965 163.367
R2723 B.n963 B.n181 163.367
R2724 B.n959 B.n957 163.367
R2725 B.n955 B.n183 163.367
R2726 B.n951 B.n949 163.367
R2727 B.n947 B.n185 163.367
R2728 B.n943 B.n941 163.367
R2729 B.n939 B.n187 163.367
R2730 B.n935 B.n933 163.367
R2731 B.n931 B.n189 163.367
R2732 B.n357 B.n356 76.6066
R2733 B.n351 B.n350 76.6066
R2734 B.n153 B.n152 76.6066
R2735 B.n159 B.n158 76.6066
R2736 B.n641 B.n319 71.676
R2737 B.n639 B.n321 71.676
R2738 B.n635 B.n634 71.676
R2739 B.n628 B.n323 71.676
R2740 B.n627 B.n626 71.676
R2741 B.n620 B.n325 71.676
R2742 B.n619 B.n618 71.676
R2743 B.n612 B.n327 71.676
R2744 B.n611 B.n610 71.676
R2745 B.n604 B.n329 71.676
R2746 B.n603 B.n602 71.676
R2747 B.n596 B.n331 71.676
R2748 B.n595 B.n594 71.676
R2749 B.n588 B.n333 71.676
R2750 B.n587 B.n586 71.676
R2751 B.n580 B.n335 71.676
R2752 B.n579 B.n578 71.676
R2753 B.n572 B.n337 71.676
R2754 B.n571 B.n570 71.676
R2755 B.n564 B.n339 71.676
R2756 B.n563 B.n562 71.676
R2757 B.n556 B.n341 71.676
R2758 B.n555 B.n554 71.676
R2759 B.n548 B.n343 71.676
R2760 B.n547 B.n546 71.676
R2761 B.n540 B.n345 71.676
R2762 B.n539 B.n538 71.676
R2763 B.n532 B.n347 71.676
R2764 B.n531 B.n530 71.676
R2765 B.n523 B.n349 71.676
R2766 B.n522 B.n521 71.676
R2767 B.n515 B.n353 71.676
R2768 B.n514 B.n513 71.676
R2769 B.n507 B.n355 71.676
R2770 B.n506 B.n359 71.676
R2771 B.n502 B.n501 71.676
R2772 B.n495 B.n361 71.676
R2773 B.n494 B.n493 71.676
R2774 B.n487 B.n363 71.676
R2775 B.n486 B.n485 71.676
R2776 B.n479 B.n365 71.676
R2777 B.n478 B.n477 71.676
R2778 B.n471 B.n367 71.676
R2779 B.n470 B.n469 71.676
R2780 B.n463 B.n369 71.676
R2781 B.n462 B.n461 71.676
R2782 B.n455 B.n371 71.676
R2783 B.n454 B.n453 71.676
R2784 B.n447 B.n373 71.676
R2785 B.n446 B.n445 71.676
R2786 B.n439 B.n375 71.676
R2787 B.n438 B.n437 71.676
R2788 B.n431 B.n377 71.676
R2789 B.n430 B.n429 71.676
R2790 B.n423 B.n379 71.676
R2791 B.n422 B.n421 71.676
R2792 B.n415 B.n381 71.676
R2793 B.n414 B.n413 71.676
R2794 B.n407 B.n383 71.676
R2795 B.n406 B.n405 71.676
R2796 B.n399 B.n385 71.676
R2797 B.n398 B.n397 71.676
R2798 B.n391 B.n387 71.676
R2799 B.n390 B.n389 71.676
R2800 B.n1184 B.n121 71.676
R2801 B.n1183 B.n1182 71.676
R2802 B.n1176 B.n123 71.676
R2803 B.n1175 B.n1174 71.676
R2804 B.n1168 B.n125 71.676
R2805 B.n1167 B.n1166 71.676
R2806 B.n1160 B.n127 71.676
R2807 B.n1159 B.n1158 71.676
R2808 B.n1152 B.n129 71.676
R2809 B.n1151 B.n1150 71.676
R2810 B.n1144 B.n131 71.676
R2811 B.n1143 B.n1142 71.676
R2812 B.n1136 B.n133 71.676
R2813 B.n1135 B.n1134 71.676
R2814 B.n1128 B.n135 71.676
R2815 B.n1127 B.n1126 71.676
R2816 B.n1120 B.n137 71.676
R2817 B.n1119 B.n1118 71.676
R2818 B.n1112 B.n139 71.676
R2819 B.n1111 B.n1110 71.676
R2820 B.n1104 B.n141 71.676
R2821 B.n1103 B.n1102 71.676
R2822 B.n1096 B.n143 71.676
R2823 B.n1095 B.n1094 71.676
R2824 B.n1088 B.n145 71.676
R2825 B.n1087 B.n1086 71.676
R2826 B.n1080 B.n147 71.676
R2827 B.n1079 B.n1078 71.676
R2828 B.n1072 B.n149 71.676
R2829 B.n1071 B.n1070 71.676
R2830 B.n1063 B.n151 71.676
R2831 B.n1062 B.n1061 71.676
R2832 B.n1055 B.n155 71.676
R2833 B.n1054 B.n1053 71.676
R2834 B.n1046 B.n157 71.676
R2835 B.n1045 B.n1044 71.676
R2836 B.n1038 B.n161 71.676
R2837 B.n1037 B.n1036 71.676
R2838 B.n1030 B.n163 71.676
R2839 B.n1029 B.n1028 71.676
R2840 B.n1022 B.n165 71.676
R2841 B.n1021 B.n1020 71.676
R2842 B.n1014 B.n167 71.676
R2843 B.n1013 B.n1012 71.676
R2844 B.n1006 B.n169 71.676
R2845 B.n1005 B.n1004 71.676
R2846 B.n998 B.n171 71.676
R2847 B.n997 B.n996 71.676
R2848 B.n990 B.n173 71.676
R2849 B.n989 B.n988 71.676
R2850 B.n982 B.n175 71.676
R2851 B.n981 B.n980 71.676
R2852 B.n974 B.n177 71.676
R2853 B.n973 B.n972 71.676
R2854 B.n966 B.n179 71.676
R2855 B.n965 B.n964 71.676
R2856 B.n958 B.n181 71.676
R2857 B.n957 B.n956 71.676
R2858 B.n950 B.n183 71.676
R2859 B.n949 B.n948 71.676
R2860 B.n942 B.n185 71.676
R2861 B.n941 B.n940 71.676
R2862 B.n934 B.n187 71.676
R2863 B.n933 B.n932 71.676
R2864 B.n932 B.n931 71.676
R2865 B.n935 B.n934 71.676
R2866 B.n940 B.n939 71.676
R2867 B.n943 B.n942 71.676
R2868 B.n948 B.n947 71.676
R2869 B.n951 B.n950 71.676
R2870 B.n956 B.n955 71.676
R2871 B.n959 B.n958 71.676
R2872 B.n964 B.n963 71.676
R2873 B.n967 B.n966 71.676
R2874 B.n972 B.n971 71.676
R2875 B.n975 B.n974 71.676
R2876 B.n980 B.n979 71.676
R2877 B.n983 B.n982 71.676
R2878 B.n988 B.n987 71.676
R2879 B.n991 B.n990 71.676
R2880 B.n996 B.n995 71.676
R2881 B.n999 B.n998 71.676
R2882 B.n1004 B.n1003 71.676
R2883 B.n1007 B.n1006 71.676
R2884 B.n1012 B.n1011 71.676
R2885 B.n1015 B.n1014 71.676
R2886 B.n1020 B.n1019 71.676
R2887 B.n1023 B.n1022 71.676
R2888 B.n1028 B.n1027 71.676
R2889 B.n1031 B.n1030 71.676
R2890 B.n1036 B.n1035 71.676
R2891 B.n1039 B.n1038 71.676
R2892 B.n1044 B.n1043 71.676
R2893 B.n1047 B.n1046 71.676
R2894 B.n1053 B.n1052 71.676
R2895 B.n1056 B.n1055 71.676
R2896 B.n1061 B.n1060 71.676
R2897 B.n1064 B.n1063 71.676
R2898 B.n1070 B.n1069 71.676
R2899 B.n1073 B.n1072 71.676
R2900 B.n1078 B.n1077 71.676
R2901 B.n1081 B.n1080 71.676
R2902 B.n1086 B.n1085 71.676
R2903 B.n1089 B.n1088 71.676
R2904 B.n1094 B.n1093 71.676
R2905 B.n1097 B.n1096 71.676
R2906 B.n1102 B.n1101 71.676
R2907 B.n1105 B.n1104 71.676
R2908 B.n1110 B.n1109 71.676
R2909 B.n1113 B.n1112 71.676
R2910 B.n1118 B.n1117 71.676
R2911 B.n1121 B.n1120 71.676
R2912 B.n1126 B.n1125 71.676
R2913 B.n1129 B.n1128 71.676
R2914 B.n1134 B.n1133 71.676
R2915 B.n1137 B.n1136 71.676
R2916 B.n1142 B.n1141 71.676
R2917 B.n1145 B.n1144 71.676
R2918 B.n1150 B.n1149 71.676
R2919 B.n1153 B.n1152 71.676
R2920 B.n1158 B.n1157 71.676
R2921 B.n1161 B.n1160 71.676
R2922 B.n1166 B.n1165 71.676
R2923 B.n1169 B.n1168 71.676
R2924 B.n1174 B.n1173 71.676
R2925 B.n1177 B.n1176 71.676
R2926 B.n1182 B.n1181 71.676
R2927 B.n1185 B.n1184 71.676
R2928 B.n642 B.n641 71.676
R2929 B.n636 B.n321 71.676
R2930 B.n634 B.n633 71.676
R2931 B.n629 B.n628 71.676
R2932 B.n626 B.n625 71.676
R2933 B.n621 B.n620 71.676
R2934 B.n618 B.n617 71.676
R2935 B.n613 B.n612 71.676
R2936 B.n610 B.n609 71.676
R2937 B.n605 B.n604 71.676
R2938 B.n602 B.n601 71.676
R2939 B.n597 B.n596 71.676
R2940 B.n594 B.n593 71.676
R2941 B.n589 B.n588 71.676
R2942 B.n586 B.n585 71.676
R2943 B.n581 B.n580 71.676
R2944 B.n578 B.n577 71.676
R2945 B.n573 B.n572 71.676
R2946 B.n570 B.n569 71.676
R2947 B.n565 B.n564 71.676
R2948 B.n562 B.n561 71.676
R2949 B.n557 B.n556 71.676
R2950 B.n554 B.n553 71.676
R2951 B.n549 B.n548 71.676
R2952 B.n546 B.n545 71.676
R2953 B.n541 B.n540 71.676
R2954 B.n538 B.n537 71.676
R2955 B.n533 B.n532 71.676
R2956 B.n530 B.n529 71.676
R2957 B.n524 B.n523 71.676
R2958 B.n521 B.n520 71.676
R2959 B.n516 B.n515 71.676
R2960 B.n513 B.n512 71.676
R2961 B.n508 B.n507 71.676
R2962 B.n503 B.n359 71.676
R2963 B.n501 B.n500 71.676
R2964 B.n496 B.n495 71.676
R2965 B.n493 B.n492 71.676
R2966 B.n488 B.n487 71.676
R2967 B.n485 B.n484 71.676
R2968 B.n480 B.n479 71.676
R2969 B.n477 B.n476 71.676
R2970 B.n472 B.n471 71.676
R2971 B.n469 B.n468 71.676
R2972 B.n464 B.n463 71.676
R2973 B.n461 B.n460 71.676
R2974 B.n456 B.n455 71.676
R2975 B.n453 B.n452 71.676
R2976 B.n448 B.n447 71.676
R2977 B.n445 B.n444 71.676
R2978 B.n440 B.n439 71.676
R2979 B.n437 B.n436 71.676
R2980 B.n432 B.n431 71.676
R2981 B.n429 B.n428 71.676
R2982 B.n424 B.n423 71.676
R2983 B.n421 B.n420 71.676
R2984 B.n416 B.n415 71.676
R2985 B.n413 B.n412 71.676
R2986 B.n408 B.n407 71.676
R2987 B.n405 B.n404 71.676
R2988 B.n400 B.n399 71.676
R2989 B.n397 B.n396 71.676
R2990 B.n392 B.n391 71.676
R2991 B.n389 B.n317 71.676
R2992 B.n647 B.n318 64.3885
R2993 B.n1190 B.n120 64.3885
R2994 B.n358 B.n357 59.5399
R2995 B.n526 B.n351 59.5399
R2996 B.n1067 B.n153 59.5399
R2997 B.n1049 B.n159 59.5399
R2998 B.n1188 B.n1187 33.8737
R2999 B.n929 B.n928 33.8737
R3000 B.n649 B.n316 33.8737
R3001 B.n645 B.n644 33.8737
R3002 B.n647 B.n314 31.9595
R3003 B.n653 B.n314 31.9595
R3004 B.n653 B.n310 31.9595
R3005 B.n659 B.n310 31.9595
R3006 B.n659 B.n306 31.9595
R3007 B.n665 B.n306 31.9595
R3008 B.n665 B.n302 31.9595
R3009 B.n671 B.n302 31.9595
R3010 B.n677 B.n298 31.9595
R3011 B.n677 B.n294 31.9595
R3012 B.n683 B.n294 31.9595
R3013 B.n683 B.n290 31.9595
R3014 B.n689 B.n290 31.9595
R3015 B.n689 B.n286 31.9595
R3016 B.n695 B.n286 31.9595
R3017 B.n695 B.n282 31.9595
R3018 B.n701 B.n282 31.9595
R3019 B.n701 B.n278 31.9595
R3020 B.n707 B.n278 31.9595
R3021 B.n707 B.n274 31.9595
R3022 B.n714 B.n274 31.9595
R3023 B.n714 B.n713 31.9595
R3024 B.n720 B.n267 31.9595
R3025 B.n726 B.n267 31.9595
R3026 B.n726 B.n263 31.9595
R3027 B.n732 B.n263 31.9595
R3028 B.n732 B.n259 31.9595
R3029 B.n738 B.n259 31.9595
R3030 B.n738 B.n255 31.9595
R3031 B.n744 B.n255 31.9595
R3032 B.n744 B.n251 31.9595
R3033 B.n751 B.n251 31.9595
R3034 B.n751 B.n750 31.9595
R3035 B.n757 B.n244 31.9595
R3036 B.n763 B.n244 31.9595
R3037 B.n763 B.n240 31.9595
R3038 B.n769 B.n240 31.9595
R3039 B.n769 B.n236 31.9595
R3040 B.n775 B.n236 31.9595
R3041 B.n775 B.n232 31.9595
R3042 B.n781 B.n232 31.9595
R3043 B.n781 B.n228 31.9595
R3044 B.n787 B.n228 31.9595
R3045 B.n793 B.n224 31.9595
R3046 B.n793 B.n220 31.9595
R3047 B.n799 B.n220 31.9595
R3048 B.n799 B.n216 31.9595
R3049 B.n805 B.n216 31.9595
R3050 B.n805 B.n212 31.9595
R3051 B.n811 B.n212 31.9595
R3052 B.n811 B.n208 31.9595
R3053 B.n817 B.n208 31.9595
R3054 B.n817 B.n204 31.9595
R3055 B.n823 B.n204 31.9595
R3056 B.n829 B.n200 31.9595
R3057 B.n829 B.n196 31.9595
R3058 B.n836 B.n196 31.9595
R3059 B.n836 B.n192 31.9595
R3060 B.n842 B.n192 31.9595
R3061 B.n842 B.n4 31.9595
R3062 B.n1320 B.n4 31.9595
R3063 B.n1320 B.n1319 31.9595
R3064 B.n1319 B.n1318 31.9595
R3065 B.n1318 B.n8 31.9595
R3066 B.n1312 B.n8 31.9595
R3067 B.n1312 B.n1311 31.9595
R3068 B.n1311 B.n1310 31.9595
R3069 B.n1310 B.n15 31.9595
R3070 B.n1304 B.n1303 31.9595
R3071 B.n1303 B.n1302 31.9595
R3072 B.n1302 B.n22 31.9595
R3073 B.n1296 B.n22 31.9595
R3074 B.n1296 B.n1295 31.9595
R3075 B.n1295 B.n1294 31.9595
R3076 B.n1294 B.n29 31.9595
R3077 B.n1288 B.n29 31.9595
R3078 B.n1288 B.n1287 31.9595
R3079 B.n1287 B.n1286 31.9595
R3080 B.n1286 B.n36 31.9595
R3081 B.n1280 B.n1279 31.9595
R3082 B.n1279 B.n1278 31.9595
R3083 B.n1278 B.n43 31.9595
R3084 B.n1272 B.n43 31.9595
R3085 B.n1272 B.n1271 31.9595
R3086 B.n1271 B.n1270 31.9595
R3087 B.n1270 B.n50 31.9595
R3088 B.n1264 B.n50 31.9595
R3089 B.n1264 B.n1263 31.9595
R3090 B.n1263 B.n1262 31.9595
R3091 B.n1256 B.n60 31.9595
R3092 B.n1256 B.n1255 31.9595
R3093 B.n1255 B.n1254 31.9595
R3094 B.n1254 B.n64 31.9595
R3095 B.n1248 B.n64 31.9595
R3096 B.n1248 B.n1247 31.9595
R3097 B.n1247 B.n1246 31.9595
R3098 B.n1246 B.n71 31.9595
R3099 B.n1240 B.n71 31.9595
R3100 B.n1240 B.n1239 31.9595
R3101 B.n1239 B.n1238 31.9595
R3102 B.n1232 B.n81 31.9595
R3103 B.n1232 B.n1231 31.9595
R3104 B.n1231 B.n1230 31.9595
R3105 B.n1230 B.n85 31.9595
R3106 B.n1224 B.n85 31.9595
R3107 B.n1224 B.n1223 31.9595
R3108 B.n1223 B.n1222 31.9595
R3109 B.n1222 B.n92 31.9595
R3110 B.n1216 B.n92 31.9595
R3111 B.n1216 B.n1215 31.9595
R3112 B.n1215 B.n1214 31.9595
R3113 B.n1214 B.n99 31.9595
R3114 B.n1208 B.n99 31.9595
R3115 B.n1208 B.n1207 31.9595
R3116 B.n1206 B.n106 31.9595
R3117 B.n1200 B.n106 31.9595
R3118 B.n1200 B.n1199 31.9595
R3119 B.n1199 B.n1198 31.9595
R3120 B.n1198 B.n113 31.9595
R3121 B.n1192 B.n113 31.9595
R3122 B.n1192 B.n1191 31.9595
R3123 B.n1191 B.n1190 31.9595
R3124 B.n787 B.t5 31.0195
R3125 B.n1280 B.t0 31.0195
R3126 B.n671 B.t15 29.1396
R3127 B.t8 B.n1206 29.1396
R3128 B.n713 B.t2 23.4998
R3129 B.n81 B.t21 23.4998
R3130 B.n757 B.t1 20.6798
R3131 B.n1262 B.t4 20.6798
R3132 B.n823 B.t6 18.7999
R3133 B.n1304 B.t3 18.7999
R3134 B B.n1322 18.0485
R3135 B.t6 B.n200 13.1601
R3136 B.t3 B.n15 13.1601
R3137 B.n750 B.t1 11.2801
R3138 B.n60 B.t4 11.2801
R3139 B.n1187 B.n1186 10.6151
R3140 B.n1186 B.n122 10.6151
R3141 B.n1180 B.n122 10.6151
R3142 B.n1180 B.n1179 10.6151
R3143 B.n1179 B.n1178 10.6151
R3144 B.n1178 B.n124 10.6151
R3145 B.n1172 B.n124 10.6151
R3146 B.n1172 B.n1171 10.6151
R3147 B.n1171 B.n1170 10.6151
R3148 B.n1170 B.n126 10.6151
R3149 B.n1164 B.n126 10.6151
R3150 B.n1164 B.n1163 10.6151
R3151 B.n1163 B.n1162 10.6151
R3152 B.n1162 B.n128 10.6151
R3153 B.n1156 B.n128 10.6151
R3154 B.n1156 B.n1155 10.6151
R3155 B.n1155 B.n1154 10.6151
R3156 B.n1154 B.n130 10.6151
R3157 B.n1148 B.n130 10.6151
R3158 B.n1148 B.n1147 10.6151
R3159 B.n1147 B.n1146 10.6151
R3160 B.n1146 B.n132 10.6151
R3161 B.n1140 B.n132 10.6151
R3162 B.n1140 B.n1139 10.6151
R3163 B.n1139 B.n1138 10.6151
R3164 B.n1138 B.n134 10.6151
R3165 B.n1132 B.n134 10.6151
R3166 B.n1132 B.n1131 10.6151
R3167 B.n1131 B.n1130 10.6151
R3168 B.n1130 B.n136 10.6151
R3169 B.n1124 B.n136 10.6151
R3170 B.n1124 B.n1123 10.6151
R3171 B.n1123 B.n1122 10.6151
R3172 B.n1122 B.n138 10.6151
R3173 B.n1116 B.n138 10.6151
R3174 B.n1116 B.n1115 10.6151
R3175 B.n1115 B.n1114 10.6151
R3176 B.n1114 B.n140 10.6151
R3177 B.n1108 B.n140 10.6151
R3178 B.n1108 B.n1107 10.6151
R3179 B.n1107 B.n1106 10.6151
R3180 B.n1106 B.n142 10.6151
R3181 B.n1100 B.n142 10.6151
R3182 B.n1100 B.n1099 10.6151
R3183 B.n1099 B.n1098 10.6151
R3184 B.n1098 B.n144 10.6151
R3185 B.n1092 B.n144 10.6151
R3186 B.n1092 B.n1091 10.6151
R3187 B.n1091 B.n1090 10.6151
R3188 B.n1090 B.n146 10.6151
R3189 B.n1084 B.n146 10.6151
R3190 B.n1084 B.n1083 10.6151
R3191 B.n1083 B.n1082 10.6151
R3192 B.n1082 B.n148 10.6151
R3193 B.n1076 B.n148 10.6151
R3194 B.n1076 B.n1075 10.6151
R3195 B.n1075 B.n1074 10.6151
R3196 B.n1074 B.n150 10.6151
R3197 B.n1068 B.n150 10.6151
R3198 B.n1066 B.n1065 10.6151
R3199 B.n1065 B.n154 10.6151
R3200 B.n1059 B.n154 10.6151
R3201 B.n1059 B.n1058 10.6151
R3202 B.n1058 B.n1057 10.6151
R3203 B.n1057 B.n156 10.6151
R3204 B.n1051 B.n156 10.6151
R3205 B.n1051 B.n1050 10.6151
R3206 B.n1048 B.n160 10.6151
R3207 B.n1042 B.n160 10.6151
R3208 B.n1042 B.n1041 10.6151
R3209 B.n1041 B.n1040 10.6151
R3210 B.n1040 B.n162 10.6151
R3211 B.n1034 B.n162 10.6151
R3212 B.n1034 B.n1033 10.6151
R3213 B.n1033 B.n1032 10.6151
R3214 B.n1032 B.n164 10.6151
R3215 B.n1026 B.n164 10.6151
R3216 B.n1026 B.n1025 10.6151
R3217 B.n1025 B.n1024 10.6151
R3218 B.n1024 B.n166 10.6151
R3219 B.n1018 B.n166 10.6151
R3220 B.n1018 B.n1017 10.6151
R3221 B.n1017 B.n1016 10.6151
R3222 B.n1016 B.n168 10.6151
R3223 B.n1010 B.n168 10.6151
R3224 B.n1010 B.n1009 10.6151
R3225 B.n1009 B.n1008 10.6151
R3226 B.n1008 B.n170 10.6151
R3227 B.n1002 B.n170 10.6151
R3228 B.n1002 B.n1001 10.6151
R3229 B.n1001 B.n1000 10.6151
R3230 B.n1000 B.n172 10.6151
R3231 B.n994 B.n172 10.6151
R3232 B.n994 B.n993 10.6151
R3233 B.n993 B.n992 10.6151
R3234 B.n992 B.n174 10.6151
R3235 B.n986 B.n174 10.6151
R3236 B.n986 B.n985 10.6151
R3237 B.n985 B.n984 10.6151
R3238 B.n984 B.n176 10.6151
R3239 B.n978 B.n176 10.6151
R3240 B.n978 B.n977 10.6151
R3241 B.n977 B.n976 10.6151
R3242 B.n976 B.n178 10.6151
R3243 B.n970 B.n178 10.6151
R3244 B.n970 B.n969 10.6151
R3245 B.n969 B.n968 10.6151
R3246 B.n968 B.n180 10.6151
R3247 B.n962 B.n180 10.6151
R3248 B.n962 B.n961 10.6151
R3249 B.n961 B.n960 10.6151
R3250 B.n960 B.n182 10.6151
R3251 B.n954 B.n182 10.6151
R3252 B.n954 B.n953 10.6151
R3253 B.n953 B.n952 10.6151
R3254 B.n952 B.n184 10.6151
R3255 B.n946 B.n184 10.6151
R3256 B.n946 B.n945 10.6151
R3257 B.n945 B.n944 10.6151
R3258 B.n944 B.n186 10.6151
R3259 B.n938 B.n186 10.6151
R3260 B.n938 B.n937 10.6151
R3261 B.n937 B.n936 10.6151
R3262 B.n936 B.n188 10.6151
R3263 B.n930 B.n188 10.6151
R3264 B.n930 B.n929 10.6151
R3265 B.n650 B.n649 10.6151
R3266 B.n651 B.n650 10.6151
R3267 B.n651 B.n308 10.6151
R3268 B.n661 B.n308 10.6151
R3269 B.n662 B.n661 10.6151
R3270 B.n663 B.n662 10.6151
R3271 B.n663 B.n300 10.6151
R3272 B.n673 B.n300 10.6151
R3273 B.n674 B.n673 10.6151
R3274 B.n675 B.n674 10.6151
R3275 B.n675 B.n292 10.6151
R3276 B.n685 B.n292 10.6151
R3277 B.n686 B.n685 10.6151
R3278 B.n687 B.n686 10.6151
R3279 B.n687 B.n284 10.6151
R3280 B.n697 B.n284 10.6151
R3281 B.n698 B.n697 10.6151
R3282 B.n699 B.n698 10.6151
R3283 B.n699 B.n276 10.6151
R3284 B.n709 B.n276 10.6151
R3285 B.n710 B.n709 10.6151
R3286 B.n711 B.n710 10.6151
R3287 B.n711 B.n269 10.6151
R3288 B.n722 B.n269 10.6151
R3289 B.n723 B.n722 10.6151
R3290 B.n724 B.n723 10.6151
R3291 B.n724 B.n261 10.6151
R3292 B.n734 B.n261 10.6151
R3293 B.n735 B.n734 10.6151
R3294 B.n736 B.n735 10.6151
R3295 B.n736 B.n253 10.6151
R3296 B.n746 B.n253 10.6151
R3297 B.n747 B.n746 10.6151
R3298 B.n748 B.n747 10.6151
R3299 B.n748 B.n246 10.6151
R3300 B.n759 B.n246 10.6151
R3301 B.n760 B.n759 10.6151
R3302 B.n761 B.n760 10.6151
R3303 B.n761 B.n238 10.6151
R3304 B.n771 B.n238 10.6151
R3305 B.n772 B.n771 10.6151
R3306 B.n773 B.n772 10.6151
R3307 B.n773 B.n230 10.6151
R3308 B.n783 B.n230 10.6151
R3309 B.n784 B.n783 10.6151
R3310 B.n785 B.n784 10.6151
R3311 B.n785 B.n222 10.6151
R3312 B.n795 B.n222 10.6151
R3313 B.n796 B.n795 10.6151
R3314 B.n797 B.n796 10.6151
R3315 B.n797 B.n214 10.6151
R3316 B.n807 B.n214 10.6151
R3317 B.n808 B.n807 10.6151
R3318 B.n809 B.n808 10.6151
R3319 B.n809 B.n206 10.6151
R3320 B.n819 B.n206 10.6151
R3321 B.n820 B.n819 10.6151
R3322 B.n821 B.n820 10.6151
R3323 B.n821 B.n198 10.6151
R3324 B.n831 B.n198 10.6151
R3325 B.n832 B.n831 10.6151
R3326 B.n834 B.n832 10.6151
R3327 B.n834 B.n833 10.6151
R3328 B.n833 B.n190 10.6151
R3329 B.n845 B.n190 10.6151
R3330 B.n846 B.n845 10.6151
R3331 B.n847 B.n846 10.6151
R3332 B.n848 B.n847 10.6151
R3333 B.n850 B.n848 10.6151
R3334 B.n851 B.n850 10.6151
R3335 B.n852 B.n851 10.6151
R3336 B.n853 B.n852 10.6151
R3337 B.n855 B.n853 10.6151
R3338 B.n856 B.n855 10.6151
R3339 B.n857 B.n856 10.6151
R3340 B.n858 B.n857 10.6151
R3341 B.n860 B.n858 10.6151
R3342 B.n861 B.n860 10.6151
R3343 B.n862 B.n861 10.6151
R3344 B.n863 B.n862 10.6151
R3345 B.n865 B.n863 10.6151
R3346 B.n866 B.n865 10.6151
R3347 B.n867 B.n866 10.6151
R3348 B.n868 B.n867 10.6151
R3349 B.n870 B.n868 10.6151
R3350 B.n871 B.n870 10.6151
R3351 B.n872 B.n871 10.6151
R3352 B.n873 B.n872 10.6151
R3353 B.n875 B.n873 10.6151
R3354 B.n876 B.n875 10.6151
R3355 B.n877 B.n876 10.6151
R3356 B.n878 B.n877 10.6151
R3357 B.n880 B.n878 10.6151
R3358 B.n881 B.n880 10.6151
R3359 B.n882 B.n881 10.6151
R3360 B.n883 B.n882 10.6151
R3361 B.n885 B.n883 10.6151
R3362 B.n886 B.n885 10.6151
R3363 B.n887 B.n886 10.6151
R3364 B.n888 B.n887 10.6151
R3365 B.n890 B.n888 10.6151
R3366 B.n891 B.n890 10.6151
R3367 B.n892 B.n891 10.6151
R3368 B.n893 B.n892 10.6151
R3369 B.n895 B.n893 10.6151
R3370 B.n896 B.n895 10.6151
R3371 B.n897 B.n896 10.6151
R3372 B.n898 B.n897 10.6151
R3373 B.n900 B.n898 10.6151
R3374 B.n901 B.n900 10.6151
R3375 B.n902 B.n901 10.6151
R3376 B.n903 B.n902 10.6151
R3377 B.n905 B.n903 10.6151
R3378 B.n906 B.n905 10.6151
R3379 B.n907 B.n906 10.6151
R3380 B.n908 B.n907 10.6151
R3381 B.n910 B.n908 10.6151
R3382 B.n911 B.n910 10.6151
R3383 B.n912 B.n911 10.6151
R3384 B.n913 B.n912 10.6151
R3385 B.n915 B.n913 10.6151
R3386 B.n916 B.n915 10.6151
R3387 B.n917 B.n916 10.6151
R3388 B.n918 B.n917 10.6151
R3389 B.n920 B.n918 10.6151
R3390 B.n921 B.n920 10.6151
R3391 B.n922 B.n921 10.6151
R3392 B.n923 B.n922 10.6151
R3393 B.n925 B.n923 10.6151
R3394 B.n926 B.n925 10.6151
R3395 B.n927 B.n926 10.6151
R3396 B.n928 B.n927 10.6151
R3397 B.n644 B.n643 10.6151
R3398 B.n643 B.n320 10.6151
R3399 B.n638 B.n320 10.6151
R3400 B.n638 B.n637 10.6151
R3401 B.n637 B.n322 10.6151
R3402 B.n632 B.n322 10.6151
R3403 B.n632 B.n631 10.6151
R3404 B.n631 B.n630 10.6151
R3405 B.n630 B.n324 10.6151
R3406 B.n624 B.n324 10.6151
R3407 B.n624 B.n623 10.6151
R3408 B.n623 B.n622 10.6151
R3409 B.n622 B.n326 10.6151
R3410 B.n616 B.n326 10.6151
R3411 B.n616 B.n615 10.6151
R3412 B.n615 B.n614 10.6151
R3413 B.n614 B.n328 10.6151
R3414 B.n608 B.n328 10.6151
R3415 B.n608 B.n607 10.6151
R3416 B.n607 B.n606 10.6151
R3417 B.n606 B.n330 10.6151
R3418 B.n600 B.n330 10.6151
R3419 B.n600 B.n599 10.6151
R3420 B.n599 B.n598 10.6151
R3421 B.n598 B.n332 10.6151
R3422 B.n592 B.n332 10.6151
R3423 B.n592 B.n591 10.6151
R3424 B.n591 B.n590 10.6151
R3425 B.n590 B.n334 10.6151
R3426 B.n584 B.n334 10.6151
R3427 B.n584 B.n583 10.6151
R3428 B.n583 B.n582 10.6151
R3429 B.n582 B.n336 10.6151
R3430 B.n576 B.n336 10.6151
R3431 B.n576 B.n575 10.6151
R3432 B.n575 B.n574 10.6151
R3433 B.n574 B.n338 10.6151
R3434 B.n568 B.n338 10.6151
R3435 B.n568 B.n567 10.6151
R3436 B.n567 B.n566 10.6151
R3437 B.n566 B.n340 10.6151
R3438 B.n560 B.n340 10.6151
R3439 B.n560 B.n559 10.6151
R3440 B.n559 B.n558 10.6151
R3441 B.n558 B.n342 10.6151
R3442 B.n552 B.n342 10.6151
R3443 B.n552 B.n551 10.6151
R3444 B.n551 B.n550 10.6151
R3445 B.n550 B.n344 10.6151
R3446 B.n544 B.n344 10.6151
R3447 B.n544 B.n543 10.6151
R3448 B.n543 B.n542 10.6151
R3449 B.n542 B.n346 10.6151
R3450 B.n536 B.n346 10.6151
R3451 B.n536 B.n535 10.6151
R3452 B.n535 B.n534 10.6151
R3453 B.n534 B.n348 10.6151
R3454 B.n528 B.n348 10.6151
R3455 B.n528 B.n527 10.6151
R3456 B.n525 B.n352 10.6151
R3457 B.n519 B.n352 10.6151
R3458 B.n519 B.n518 10.6151
R3459 B.n518 B.n517 10.6151
R3460 B.n517 B.n354 10.6151
R3461 B.n511 B.n354 10.6151
R3462 B.n511 B.n510 10.6151
R3463 B.n510 B.n509 10.6151
R3464 B.n505 B.n504 10.6151
R3465 B.n504 B.n360 10.6151
R3466 B.n499 B.n360 10.6151
R3467 B.n499 B.n498 10.6151
R3468 B.n498 B.n497 10.6151
R3469 B.n497 B.n362 10.6151
R3470 B.n491 B.n362 10.6151
R3471 B.n491 B.n490 10.6151
R3472 B.n490 B.n489 10.6151
R3473 B.n489 B.n364 10.6151
R3474 B.n483 B.n364 10.6151
R3475 B.n483 B.n482 10.6151
R3476 B.n482 B.n481 10.6151
R3477 B.n481 B.n366 10.6151
R3478 B.n475 B.n366 10.6151
R3479 B.n475 B.n474 10.6151
R3480 B.n474 B.n473 10.6151
R3481 B.n473 B.n368 10.6151
R3482 B.n467 B.n368 10.6151
R3483 B.n467 B.n466 10.6151
R3484 B.n466 B.n465 10.6151
R3485 B.n465 B.n370 10.6151
R3486 B.n459 B.n370 10.6151
R3487 B.n459 B.n458 10.6151
R3488 B.n458 B.n457 10.6151
R3489 B.n457 B.n372 10.6151
R3490 B.n451 B.n372 10.6151
R3491 B.n451 B.n450 10.6151
R3492 B.n450 B.n449 10.6151
R3493 B.n449 B.n374 10.6151
R3494 B.n443 B.n374 10.6151
R3495 B.n443 B.n442 10.6151
R3496 B.n442 B.n441 10.6151
R3497 B.n441 B.n376 10.6151
R3498 B.n435 B.n376 10.6151
R3499 B.n435 B.n434 10.6151
R3500 B.n434 B.n433 10.6151
R3501 B.n433 B.n378 10.6151
R3502 B.n427 B.n378 10.6151
R3503 B.n427 B.n426 10.6151
R3504 B.n426 B.n425 10.6151
R3505 B.n425 B.n380 10.6151
R3506 B.n419 B.n380 10.6151
R3507 B.n419 B.n418 10.6151
R3508 B.n418 B.n417 10.6151
R3509 B.n417 B.n382 10.6151
R3510 B.n411 B.n382 10.6151
R3511 B.n411 B.n410 10.6151
R3512 B.n410 B.n409 10.6151
R3513 B.n409 B.n384 10.6151
R3514 B.n403 B.n384 10.6151
R3515 B.n403 B.n402 10.6151
R3516 B.n402 B.n401 10.6151
R3517 B.n401 B.n386 10.6151
R3518 B.n395 B.n386 10.6151
R3519 B.n395 B.n394 10.6151
R3520 B.n394 B.n393 10.6151
R3521 B.n393 B.n388 10.6151
R3522 B.n388 B.n316 10.6151
R3523 B.n645 B.n312 10.6151
R3524 B.n655 B.n312 10.6151
R3525 B.n656 B.n655 10.6151
R3526 B.n657 B.n656 10.6151
R3527 B.n657 B.n304 10.6151
R3528 B.n667 B.n304 10.6151
R3529 B.n668 B.n667 10.6151
R3530 B.n669 B.n668 10.6151
R3531 B.n669 B.n296 10.6151
R3532 B.n679 B.n296 10.6151
R3533 B.n680 B.n679 10.6151
R3534 B.n681 B.n680 10.6151
R3535 B.n681 B.n288 10.6151
R3536 B.n691 B.n288 10.6151
R3537 B.n692 B.n691 10.6151
R3538 B.n693 B.n692 10.6151
R3539 B.n693 B.n280 10.6151
R3540 B.n703 B.n280 10.6151
R3541 B.n704 B.n703 10.6151
R3542 B.n705 B.n704 10.6151
R3543 B.n705 B.n272 10.6151
R3544 B.n716 B.n272 10.6151
R3545 B.n717 B.n716 10.6151
R3546 B.n718 B.n717 10.6151
R3547 B.n718 B.n265 10.6151
R3548 B.n728 B.n265 10.6151
R3549 B.n729 B.n728 10.6151
R3550 B.n730 B.n729 10.6151
R3551 B.n730 B.n257 10.6151
R3552 B.n740 B.n257 10.6151
R3553 B.n741 B.n740 10.6151
R3554 B.n742 B.n741 10.6151
R3555 B.n742 B.n249 10.6151
R3556 B.n753 B.n249 10.6151
R3557 B.n754 B.n753 10.6151
R3558 B.n755 B.n754 10.6151
R3559 B.n755 B.n242 10.6151
R3560 B.n765 B.n242 10.6151
R3561 B.n766 B.n765 10.6151
R3562 B.n767 B.n766 10.6151
R3563 B.n767 B.n234 10.6151
R3564 B.n777 B.n234 10.6151
R3565 B.n778 B.n777 10.6151
R3566 B.n779 B.n778 10.6151
R3567 B.n779 B.n226 10.6151
R3568 B.n789 B.n226 10.6151
R3569 B.n790 B.n789 10.6151
R3570 B.n791 B.n790 10.6151
R3571 B.n791 B.n218 10.6151
R3572 B.n801 B.n218 10.6151
R3573 B.n802 B.n801 10.6151
R3574 B.n803 B.n802 10.6151
R3575 B.n803 B.n210 10.6151
R3576 B.n813 B.n210 10.6151
R3577 B.n814 B.n813 10.6151
R3578 B.n815 B.n814 10.6151
R3579 B.n815 B.n202 10.6151
R3580 B.n825 B.n202 10.6151
R3581 B.n826 B.n825 10.6151
R3582 B.n827 B.n826 10.6151
R3583 B.n827 B.n194 10.6151
R3584 B.n838 B.n194 10.6151
R3585 B.n839 B.n838 10.6151
R3586 B.n840 B.n839 10.6151
R3587 B.n840 B.n0 10.6151
R3588 B.n1316 B.n1 10.6151
R3589 B.n1316 B.n1315 10.6151
R3590 B.n1315 B.n1314 10.6151
R3591 B.n1314 B.n10 10.6151
R3592 B.n1308 B.n10 10.6151
R3593 B.n1308 B.n1307 10.6151
R3594 B.n1307 B.n1306 10.6151
R3595 B.n1306 B.n17 10.6151
R3596 B.n1300 B.n17 10.6151
R3597 B.n1300 B.n1299 10.6151
R3598 B.n1299 B.n1298 10.6151
R3599 B.n1298 B.n24 10.6151
R3600 B.n1292 B.n24 10.6151
R3601 B.n1292 B.n1291 10.6151
R3602 B.n1291 B.n1290 10.6151
R3603 B.n1290 B.n31 10.6151
R3604 B.n1284 B.n31 10.6151
R3605 B.n1284 B.n1283 10.6151
R3606 B.n1283 B.n1282 10.6151
R3607 B.n1282 B.n38 10.6151
R3608 B.n1276 B.n38 10.6151
R3609 B.n1276 B.n1275 10.6151
R3610 B.n1275 B.n1274 10.6151
R3611 B.n1274 B.n45 10.6151
R3612 B.n1268 B.n45 10.6151
R3613 B.n1268 B.n1267 10.6151
R3614 B.n1267 B.n1266 10.6151
R3615 B.n1266 B.n52 10.6151
R3616 B.n1260 B.n52 10.6151
R3617 B.n1260 B.n1259 10.6151
R3618 B.n1259 B.n1258 10.6151
R3619 B.n1258 B.n58 10.6151
R3620 B.n1252 B.n58 10.6151
R3621 B.n1252 B.n1251 10.6151
R3622 B.n1251 B.n1250 10.6151
R3623 B.n1250 B.n66 10.6151
R3624 B.n1244 B.n66 10.6151
R3625 B.n1244 B.n1243 10.6151
R3626 B.n1243 B.n1242 10.6151
R3627 B.n1242 B.n73 10.6151
R3628 B.n1236 B.n73 10.6151
R3629 B.n1236 B.n1235 10.6151
R3630 B.n1235 B.n1234 10.6151
R3631 B.n1234 B.n79 10.6151
R3632 B.n1228 B.n79 10.6151
R3633 B.n1228 B.n1227 10.6151
R3634 B.n1227 B.n1226 10.6151
R3635 B.n1226 B.n87 10.6151
R3636 B.n1220 B.n87 10.6151
R3637 B.n1220 B.n1219 10.6151
R3638 B.n1219 B.n1218 10.6151
R3639 B.n1218 B.n94 10.6151
R3640 B.n1212 B.n94 10.6151
R3641 B.n1212 B.n1211 10.6151
R3642 B.n1211 B.n1210 10.6151
R3643 B.n1210 B.n101 10.6151
R3644 B.n1204 B.n101 10.6151
R3645 B.n1204 B.n1203 10.6151
R3646 B.n1203 B.n1202 10.6151
R3647 B.n1202 B.n108 10.6151
R3648 B.n1196 B.n108 10.6151
R3649 B.n1196 B.n1195 10.6151
R3650 B.n1195 B.n1194 10.6151
R3651 B.n1194 B.n115 10.6151
R3652 B.n1188 B.n115 10.6151
R3653 B.n720 B.t2 8.46023
R3654 B.n1238 B.t21 8.46023
R3655 B.n1067 B.n1066 6.5566
R3656 B.n1050 B.n1049 6.5566
R3657 B.n526 B.n525 6.5566
R3658 B.n509 B.n358 6.5566
R3659 B.n1068 B.n1067 4.05904
R3660 B.n1049 B.n1048 4.05904
R3661 B.n527 B.n526 4.05904
R3662 B.n505 B.n358 4.05904
R3663 B.t15 B.n298 2.82041
R3664 B.n1207 B.t8 2.82041
R3665 B.n1322 B.n0 2.81026
R3666 B.n1322 B.n1 2.81026
R3667 B.t5 B.n224 0.94047
R3668 B.t0 B.n36 0.94047
R3669 VN.n72 VN.n71 161.3
R3670 VN.n70 VN.n38 161.3
R3671 VN.n69 VN.n68 161.3
R3672 VN.n67 VN.n39 161.3
R3673 VN.n66 VN.n65 161.3
R3674 VN.n64 VN.n40 161.3
R3675 VN.n63 VN.n62 161.3
R3676 VN.n61 VN.n41 161.3
R3677 VN.n60 VN.n59 161.3
R3678 VN.n58 VN.n42 161.3
R3679 VN.n57 VN.n56 161.3
R3680 VN.n55 VN.n44 161.3
R3681 VN.n54 VN.n53 161.3
R3682 VN.n52 VN.n45 161.3
R3683 VN.n51 VN.n50 161.3
R3684 VN.n49 VN.n46 161.3
R3685 VN.n35 VN.n34 161.3
R3686 VN.n33 VN.n1 161.3
R3687 VN.n32 VN.n31 161.3
R3688 VN.n30 VN.n2 161.3
R3689 VN.n29 VN.n28 161.3
R3690 VN.n27 VN.n3 161.3
R3691 VN.n26 VN.n25 161.3
R3692 VN.n24 VN.n4 161.3
R3693 VN.n23 VN.n22 161.3
R3694 VN.n20 VN.n5 161.3
R3695 VN.n19 VN.n18 161.3
R3696 VN.n17 VN.n6 161.3
R3697 VN.n16 VN.n15 161.3
R3698 VN.n14 VN.n7 161.3
R3699 VN.n13 VN.n12 161.3
R3700 VN.n11 VN.n8 161.3
R3701 VN.n48 VN.t6 153.856
R3702 VN.n10 VN.t7 153.856
R3703 VN.n9 VN.t2 120.701
R3704 VN.n21 VN.t5 120.701
R3705 VN.n0 VN.t0 120.701
R3706 VN.n47 VN.t4 120.701
R3707 VN.n43 VN.t3 120.701
R3708 VN.n37 VN.t1 120.701
R3709 VN.n36 VN.n0 81.504
R3710 VN.n73 VN.n37 81.504
R3711 VN.n10 VN.n9 63.5476
R3712 VN.n48 VN.n47 63.5476
R3713 VN VN.n73 60.5738
R3714 VN.n15 VN.n6 56.5193
R3715 VN.n28 VN.n2 56.5193
R3716 VN.n53 VN.n44 56.5193
R3717 VN.n65 VN.n39 56.5193
R3718 VN.n13 VN.n8 24.4675
R3719 VN.n14 VN.n13 24.4675
R3720 VN.n15 VN.n14 24.4675
R3721 VN.n19 VN.n6 24.4675
R3722 VN.n20 VN.n19 24.4675
R3723 VN.n22 VN.n20 24.4675
R3724 VN.n26 VN.n4 24.4675
R3725 VN.n27 VN.n26 24.4675
R3726 VN.n28 VN.n27 24.4675
R3727 VN.n32 VN.n2 24.4675
R3728 VN.n33 VN.n32 24.4675
R3729 VN.n34 VN.n33 24.4675
R3730 VN.n53 VN.n52 24.4675
R3731 VN.n52 VN.n51 24.4675
R3732 VN.n51 VN.n46 24.4675
R3733 VN.n65 VN.n64 24.4675
R3734 VN.n64 VN.n63 24.4675
R3735 VN.n63 VN.n41 24.4675
R3736 VN.n59 VN.n58 24.4675
R3737 VN.n58 VN.n57 24.4675
R3738 VN.n57 VN.n44 24.4675
R3739 VN.n71 VN.n70 24.4675
R3740 VN.n70 VN.n69 24.4675
R3741 VN.n69 VN.n39 24.4675
R3742 VN.n21 VN.n4 13.4574
R3743 VN.n43 VN.n41 13.4574
R3744 VN.n9 VN.n8 11.0107
R3745 VN.n22 VN.n21 11.0107
R3746 VN.n47 VN.n46 11.0107
R3747 VN.n59 VN.n43 11.0107
R3748 VN.n34 VN.n0 8.56395
R3749 VN.n71 VN.n37 8.56395
R3750 VN.n11 VN.n10 3.20386
R3751 VN.n49 VN.n48 3.20386
R3752 VN.n73 VN.n72 0.354971
R3753 VN.n36 VN.n35 0.354971
R3754 VN VN.n36 0.26696
R3755 VN.n72 VN.n38 0.189894
R3756 VN.n68 VN.n38 0.189894
R3757 VN.n68 VN.n67 0.189894
R3758 VN.n67 VN.n66 0.189894
R3759 VN.n66 VN.n40 0.189894
R3760 VN.n62 VN.n40 0.189894
R3761 VN.n62 VN.n61 0.189894
R3762 VN.n61 VN.n60 0.189894
R3763 VN.n60 VN.n42 0.189894
R3764 VN.n56 VN.n42 0.189894
R3765 VN.n56 VN.n55 0.189894
R3766 VN.n55 VN.n54 0.189894
R3767 VN.n54 VN.n45 0.189894
R3768 VN.n50 VN.n45 0.189894
R3769 VN.n50 VN.n49 0.189894
R3770 VN.n12 VN.n11 0.189894
R3771 VN.n12 VN.n7 0.189894
R3772 VN.n16 VN.n7 0.189894
R3773 VN.n17 VN.n16 0.189894
R3774 VN.n18 VN.n17 0.189894
R3775 VN.n18 VN.n5 0.189894
R3776 VN.n23 VN.n5 0.189894
R3777 VN.n24 VN.n23 0.189894
R3778 VN.n25 VN.n24 0.189894
R3779 VN.n25 VN.n3 0.189894
R3780 VN.n29 VN.n3 0.189894
R3781 VN.n30 VN.n29 0.189894
R3782 VN.n31 VN.n30 0.189894
R3783 VN.n31 VN.n1 0.189894
R3784 VN.n35 VN.n1 0.189894
R3785 VDD2.n2 VDD2.n1 60.162
R3786 VDD2.n2 VDD2.n0 60.162
R3787 VDD2 VDD2.n5 60.1592
R3788 VDD2.n4 VDD2.n3 58.515
R3789 VDD2.n4 VDD2.n2 54.6679
R3790 VDD2 VDD2.n4 1.76128
R3791 VDD2.n5 VDD2.t3 1.09261
R3792 VDD2.n5 VDD2.t1 1.09261
R3793 VDD2.n3 VDD2.t6 1.09261
R3794 VDD2.n3 VDD2.t4 1.09261
R3795 VDD2.n1 VDD2.t2 1.09261
R3796 VDD2.n1 VDD2.t7 1.09261
R3797 VDD2.n0 VDD2.t0 1.09261
R3798 VDD2.n0 VDD2.t5 1.09261
C0 VDD2 VTAIL 10.2974f
C1 VDD1 VDD2 2.30735f
C2 VP VN 10.0453f
C3 VP VTAIL 14.110099f
C4 VN VTAIL 14.096f
C5 VP VDD1 14.119401f
C6 VP VDD2 0.628351f
C7 VDD1 VN 0.153714f
C8 VDD2 VN 13.6466f
C9 VDD1 VTAIL 10.2362f
C10 VDD2 B 6.877338f
C11 VDD1 B 7.421714f
C12 VTAIL B 14.888446f
C13 VN B 19.906519f
C14 VP B 18.506662f
C15 VDD2.t0 B 0.377159f
C16 VDD2.t5 B 0.377159f
C17 VDD2.n0 B 3.45153f
C18 VDD2.t2 B 0.377159f
C19 VDD2.t7 B 0.377159f
C20 VDD2.n1 B 3.45153f
C21 VDD2.n2 B 4.49236f
C22 VDD2.t6 B 0.377159f
C23 VDD2.t4 B 0.377159f
C24 VDD2.n3 B 3.43342f
C25 VDD2.n4 B 3.97038f
C26 VDD2.t3 B 0.377159f
C27 VDD2.t1 B 0.377159f
C28 VDD2.n5 B 3.45148f
C29 VN.t0 B 3.02892f
C30 VN.n0 B 1.10934f
C31 VN.n1 B 0.016777f
C32 VN.n2 B 0.026828f
C33 VN.n3 B 0.016777f
C34 VN.n4 B 0.02432f
C35 VN.n5 B 0.016777f
C36 VN.n6 B 0.024491f
C37 VN.n7 B 0.016777f
C38 VN.n8 B 0.022776f
C39 VN.t2 B 3.02892f
C40 VN.n9 B 1.10161f
C41 VN.t7 B 3.28143f
C42 VN.n10 B 1.0524f
C43 VN.n11 B 0.21014f
C44 VN.n12 B 0.016777f
C45 VN.n13 B 0.031267f
C46 VN.n14 B 0.031267f
C47 VN.n15 B 0.024491f
C48 VN.n16 B 0.016777f
C49 VN.n17 B 0.016777f
C50 VN.n18 B 0.016777f
C51 VN.n19 B 0.031267f
C52 VN.n20 B 0.031267f
C53 VN.t5 B 3.02892f
C54 VN.n21 B 1.04399f
C55 VN.n22 B 0.022776f
C56 VN.n23 B 0.016777f
C57 VN.n24 B 0.016777f
C58 VN.n25 B 0.016777f
C59 VN.n26 B 0.031267f
C60 VN.n27 B 0.031267f
C61 VN.n28 B 0.022153f
C62 VN.n29 B 0.016777f
C63 VN.n30 B 0.016777f
C64 VN.n31 B 0.016777f
C65 VN.n32 B 0.031267f
C66 VN.n33 B 0.031267f
C67 VN.n34 B 0.021232f
C68 VN.n35 B 0.027077f
C69 VN.n36 B 0.046882f
C70 VN.t1 B 3.02892f
C71 VN.n37 B 1.10934f
C72 VN.n38 B 0.016777f
C73 VN.n39 B 0.026828f
C74 VN.n40 B 0.016777f
C75 VN.n41 B 0.02432f
C76 VN.n42 B 0.016777f
C77 VN.t3 B 3.02892f
C78 VN.n43 B 1.04399f
C79 VN.n44 B 0.024491f
C80 VN.n45 B 0.016777f
C81 VN.n46 B 0.022776f
C82 VN.t6 B 3.28143f
C83 VN.t4 B 3.02892f
C84 VN.n47 B 1.10161f
C85 VN.n48 B 1.0524f
C86 VN.n49 B 0.21014f
C87 VN.n50 B 0.016777f
C88 VN.n51 B 0.031267f
C89 VN.n52 B 0.031267f
C90 VN.n53 B 0.024491f
C91 VN.n54 B 0.016777f
C92 VN.n55 B 0.016777f
C93 VN.n56 B 0.016777f
C94 VN.n57 B 0.031267f
C95 VN.n58 B 0.031267f
C96 VN.n59 B 0.022776f
C97 VN.n60 B 0.016777f
C98 VN.n61 B 0.016777f
C99 VN.n62 B 0.016777f
C100 VN.n63 B 0.031267f
C101 VN.n64 B 0.031267f
C102 VN.n65 B 0.022153f
C103 VN.n66 B 0.016777f
C104 VN.n67 B 0.016777f
C105 VN.n68 B 0.016777f
C106 VN.n69 B 0.031267f
C107 VN.n70 B 0.031267f
C108 VN.n71 B 0.021232f
C109 VN.n72 B 0.027077f
C110 VN.n73 B 1.25285f
C111 VTAIL.t0 B 0.272698f
C112 VTAIL.t4 B 0.272698f
C113 VTAIL.n0 B 2.41983f
C114 VTAIL.n1 B 0.409915f
C115 VTAIL.n2 B 0.025341f
C116 VTAIL.n3 B 0.019034f
C117 VTAIL.n4 B 0.010228f
C118 VTAIL.n5 B 0.024175f
C119 VTAIL.n6 B 0.01083f
C120 VTAIL.n7 B 0.019034f
C121 VTAIL.n8 B 0.010228f
C122 VTAIL.n9 B 0.024175f
C123 VTAIL.n10 B 0.01083f
C124 VTAIL.n11 B 0.019034f
C125 VTAIL.n12 B 0.010529f
C126 VTAIL.n13 B 0.024175f
C127 VTAIL.n14 B 0.01083f
C128 VTAIL.n15 B 0.019034f
C129 VTAIL.n16 B 0.010228f
C130 VTAIL.n17 B 0.024175f
C131 VTAIL.n18 B 0.01083f
C132 VTAIL.n19 B 0.019034f
C133 VTAIL.n20 B 0.010228f
C134 VTAIL.n21 B 0.024175f
C135 VTAIL.n22 B 0.01083f
C136 VTAIL.n23 B 0.019034f
C137 VTAIL.n24 B 0.010228f
C138 VTAIL.n25 B 0.024175f
C139 VTAIL.n26 B 0.01083f
C140 VTAIL.n27 B 0.019034f
C141 VTAIL.n28 B 0.010228f
C142 VTAIL.n29 B 0.024175f
C143 VTAIL.n30 B 0.01083f
C144 VTAIL.n31 B 0.019034f
C145 VTAIL.n32 B 0.010228f
C146 VTAIL.n33 B 0.018132f
C147 VTAIL.n34 B 0.014281f
C148 VTAIL.t3 B 0.040067f
C149 VTAIL.n35 B 0.139081f
C150 VTAIL.n36 B 1.51142f
C151 VTAIL.n37 B 0.010228f
C152 VTAIL.n38 B 0.01083f
C153 VTAIL.n39 B 0.024175f
C154 VTAIL.n40 B 0.024175f
C155 VTAIL.n41 B 0.01083f
C156 VTAIL.n42 B 0.010228f
C157 VTAIL.n43 B 0.019034f
C158 VTAIL.n44 B 0.019034f
C159 VTAIL.n45 B 0.010228f
C160 VTAIL.n46 B 0.01083f
C161 VTAIL.n47 B 0.024175f
C162 VTAIL.n48 B 0.024175f
C163 VTAIL.n49 B 0.01083f
C164 VTAIL.n50 B 0.010228f
C165 VTAIL.n51 B 0.019034f
C166 VTAIL.n52 B 0.019034f
C167 VTAIL.n53 B 0.010228f
C168 VTAIL.n54 B 0.01083f
C169 VTAIL.n55 B 0.024175f
C170 VTAIL.n56 B 0.024175f
C171 VTAIL.n57 B 0.01083f
C172 VTAIL.n58 B 0.010228f
C173 VTAIL.n59 B 0.019034f
C174 VTAIL.n60 B 0.019034f
C175 VTAIL.n61 B 0.010228f
C176 VTAIL.n62 B 0.01083f
C177 VTAIL.n63 B 0.024175f
C178 VTAIL.n64 B 0.024175f
C179 VTAIL.n65 B 0.01083f
C180 VTAIL.n66 B 0.010228f
C181 VTAIL.n67 B 0.019034f
C182 VTAIL.n68 B 0.019034f
C183 VTAIL.n69 B 0.010228f
C184 VTAIL.n70 B 0.01083f
C185 VTAIL.n71 B 0.024175f
C186 VTAIL.n72 B 0.024175f
C187 VTAIL.n73 B 0.01083f
C188 VTAIL.n74 B 0.010228f
C189 VTAIL.n75 B 0.019034f
C190 VTAIL.n76 B 0.019034f
C191 VTAIL.n77 B 0.010228f
C192 VTAIL.n78 B 0.010228f
C193 VTAIL.n79 B 0.01083f
C194 VTAIL.n80 B 0.024175f
C195 VTAIL.n81 B 0.024175f
C196 VTAIL.n82 B 0.024175f
C197 VTAIL.n83 B 0.010529f
C198 VTAIL.n84 B 0.010228f
C199 VTAIL.n85 B 0.019034f
C200 VTAIL.n86 B 0.019034f
C201 VTAIL.n87 B 0.010228f
C202 VTAIL.n88 B 0.01083f
C203 VTAIL.n89 B 0.024175f
C204 VTAIL.n90 B 0.024175f
C205 VTAIL.n91 B 0.01083f
C206 VTAIL.n92 B 0.010228f
C207 VTAIL.n93 B 0.019034f
C208 VTAIL.n94 B 0.019034f
C209 VTAIL.n95 B 0.010228f
C210 VTAIL.n96 B 0.01083f
C211 VTAIL.n97 B 0.024175f
C212 VTAIL.n98 B 0.049838f
C213 VTAIL.n99 B 0.01083f
C214 VTAIL.n100 B 0.010228f
C215 VTAIL.n101 B 0.041136f
C216 VTAIL.n102 B 0.027539f
C217 VTAIL.n103 B 0.252306f
C218 VTAIL.n104 B 0.025341f
C219 VTAIL.n105 B 0.019034f
C220 VTAIL.n106 B 0.010228f
C221 VTAIL.n107 B 0.024175f
C222 VTAIL.n108 B 0.01083f
C223 VTAIL.n109 B 0.019034f
C224 VTAIL.n110 B 0.010228f
C225 VTAIL.n111 B 0.024175f
C226 VTAIL.n112 B 0.01083f
C227 VTAIL.n113 B 0.019034f
C228 VTAIL.n114 B 0.010529f
C229 VTAIL.n115 B 0.024175f
C230 VTAIL.n116 B 0.01083f
C231 VTAIL.n117 B 0.019034f
C232 VTAIL.n118 B 0.010228f
C233 VTAIL.n119 B 0.024175f
C234 VTAIL.n120 B 0.01083f
C235 VTAIL.n121 B 0.019034f
C236 VTAIL.n122 B 0.010228f
C237 VTAIL.n123 B 0.024175f
C238 VTAIL.n124 B 0.01083f
C239 VTAIL.n125 B 0.019034f
C240 VTAIL.n126 B 0.010228f
C241 VTAIL.n127 B 0.024175f
C242 VTAIL.n128 B 0.01083f
C243 VTAIL.n129 B 0.019034f
C244 VTAIL.n130 B 0.010228f
C245 VTAIL.n131 B 0.024175f
C246 VTAIL.n132 B 0.01083f
C247 VTAIL.n133 B 0.019034f
C248 VTAIL.n134 B 0.010228f
C249 VTAIL.n135 B 0.018132f
C250 VTAIL.n136 B 0.014281f
C251 VTAIL.t8 B 0.040067f
C252 VTAIL.n137 B 0.139081f
C253 VTAIL.n138 B 1.51142f
C254 VTAIL.n139 B 0.010228f
C255 VTAIL.n140 B 0.01083f
C256 VTAIL.n141 B 0.024175f
C257 VTAIL.n142 B 0.024175f
C258 VTAIL.n143 B 0.01083f
C259 VTAIL.n144 B 0.010228f
C260 VTAIL.n145 B 0.019034f
C261 VTAIL.n146 B 0.019034f
C262 VTAIL.n147 B 0.010228f
C263 VTAIL.n148 B 0.01083f
C264 VTAIL.n149 B 0.024175f
C265 VTAIL.n150 B 0.024175f
C266 VTAIL.n151 B 0.01083f
C267 VTAIL.n152 B 0.010228f
C268 VTAIL.n153 B 0.019034f
C269 VTAIL.n154 B 0.019034f
C270 VTAIL.n155 B 0.010228f
C271 VTAIL.n156 B 0.01083f
C272 VTAIL.n157 B 0.024175f
C273 VTAIL.n158 B 0.024175f
C274 VTAIL.n159 B 0.01083f
C275 VTAIL.n160 B 0.010228f
C276 VTAIL.n161 B 0.019034f
C277 VTAIL.n162 B 0.019034f
C278 VTAIL.n163 B 0.010228f
C279 VTAIL.n164 B 0.01083f
C280 VTAIL.n165 B 0.024175f
C281 VTAIL.n166 B 0.024175f
C282 VTAIL.n167 B 0.01083f
C283 VTAIL.n168 B 0.010228f
C284 VTAIL.n169 B 0.019034f
C285 VTAIL.n170 B 0.019034f
C286 VTAIL.n171 B 0.010228f
C287 VTAIL.n172 B 0.01083f
C288 VTAIL.n173 B 0.024175f
C289 VTAIL.n174 B 0.024175f
C290 VTAIL.n175 B 0.01083f
C291 VTAIL.n176 B 0.010228f
C292 VTAIL.n177 B 0.019034f
C293 VTAIL.n178 B 0.019034f
C294 VTAIL.n179 B 0.010228f
C295 VTAIL.n180 B 0.010228f
C296 VTAIL.n181 B 0.01083f
C297 VTAIL.n182 B 0.024175f
C298 VTAIL.n183 B 0.024175f
C299 VTAIL.n184 B 0.024175f
C300 VTAIL.n185 B 0.010529f
C301 VTAIL.n186 B 0.010228f
C302 VTAIL.n187 B 0.019034f
C303 VTAIL.n188 B 0.019034f
C304 VTAIL.n189 B 0.010228f
C305 VTAIL.n190 B 0.01083f
C306 VTAIL.n191 B 0.024175f
C307 VTAIL.n192 B 0.024175f
C308 VTAIL.n193 B 0.01083f
C309 VTAIL.n194 B 0.010228f
C310 VTAIL.n195 B 0.019034f
C311 VTAIL.n196 B 0.019034f
C312 VTAIL.n197 B 0.010228f
C313 VTAIL.n198 B 0.01083f
C314 VTAIL.n199 B 0.024175f
C315 VTAIL.n200 B 0.049838f
C316 VTAIL.n201 B 0.01083f
C317 VTAIL.n202 B 0.010228f
C318 VTAIL.n203 B 0.041136f
C319 VTAIL.n204 B 0.027539f
C320 VTAIL.n205 B 0.252306f
C321 VTAIL.t11 B 0.272698f
C322 VTAIL.t13 B 0.272698f
C323 VTAIL.n206 B 2.41983f
C324 VTAIL.n207 B 0.615192f
C325 VTAIL.n208 B 0.025341f
C326 VTAIL.n209 B 0.019034f
C327 VTAIL.n210 B 0.010228f
C328 VTAIL.n211 B 0.024175f
C329 VTAIL.n212 B 0.01083f
C330 VTAIL.n213 B 0.019034f
C331 VTAIL.n214 B 0.010228f
C332 VTAIL.n215 B 0.024175f
C333 VTAIL.n216 B 0.01083f
C334 VTAIL.n217 B 0.019034f
C335 VTAIL.n218 B 0.010529f
C336 VTAIL.n219 B 0.024175f
C337 VTAIL.n220 B 0.01083f
C338 VTAIL.n221 B 0.019034f
C339 VTAIL.n222 B 0.010228f
C340 VTAIL.n223 B 0.024175f
C341 VTAIL.n224 B 0.01083f
C342 VTAIL.n225 B 0.019034f
C343 VTAIL.n226 B 0.010228f
C344 VTAIL.n227 B 0.024175f
C345 VTAIL.n228 B 0.01083f
C346 VTAIL.n229 B 0.019034f
C347 VTAIL.n230 B 0.010228f
C348 VTAIL.n231 B 0.024175f
C349 VTAIL.n232 B 0.01083f
C350 VTAIL.n233 B 0.019034f
C351 VTAIL.n234 B 0.010228f
C352 VTAIL.n235 B 0.024175f
C353 VTAIL.n236 B 0.01083f
C354 VTAIL.n237 B 0.019034f
C355 VTAIL.n238 B 0.010228f
C356 VTAIL.n239 B 0.018132f
C357 VTAIL.n240 B 0.014281f
C358 VTAIL.t7 B 0.040067f
C359 VTAIL.n241 B 0.139081f
C360 VTAIL.n242 B 1.51142f
C361 VTAIL.n243 B 0.010228f
C362 VTAIL.n244 B 0.01083f
C363 VTAIL.n245 B 0.024175f
C364 VTAIL.n246 B 0.024175f
C365 VTAIL.n247 B 0.01083f
C366 VTAIL.n248 B 0.010228f
C367 VTAIL.n249 B 0.019034f
C368 VTAIL.n250 B 0.019034f
C369 VTAIL.n251 B 0.010228f
C370 VTAIL.n252 B 0.01083f
C371 VTAIL.n253 B 0.024175f
C372 VTAIL.n254 B 0.024175f
C373 VTAIL.n255 B 0.01083f
C374 VTAIL.n256 B 0.010228f
C375 VTAIL.n257 B 0.019034f
C376 VTAIL.n258 B 0.019034f
C377 VTAIL.n259 B 0.010228f
C378 VTAIL.n260 B 0.01083f
C379 VTAIL.n261 B 0.024175f
C380 VTAIL.n262 B 0.024175f
C381 VTAIL.n263 B 0.01083f
C382 VTAIL.n264 B 0.010228f
C383 VTAIL.n265 B 0.019034f
C384 VTAIL.n266 B 0.019034f
C385 VTAIL.n267 B 0.010228f
C386 VTAIL.n268 B 0.01083f
C387 VTAIL.n269 B 0.024175f
C388 VTAIL.n270 B 0.024175f
C389 VTAIL.n271 B 0.01083f
C390 VTAIL.n272 B 0.010228f
C391 VTAIL.n273 B 0.019034f
C392 VTAIL.n274 B 0.019034f
C393 VTAIL.n275 B 0.010228f
C394 VTAIL.n276 B 0.01083f
C395 VTAIL.n277 B 0.024175f
C396 VTAIL.n278 B 0.024175f
C397 VTAIL.n279 B 0.01083f
C398 VTAIL.n280 B 0.010228f
C399 VTAIL.n281 B 0.019034f
C400 VTAIL.n282 B 0.019034f
C401 VTAIL.n283 B 0.010228f
C402 VTAIL.n284 B 0.010228f
C403 VTAIL.n285 B 0.01083f
C404 VTAIL.n286 B 0.024175f
C405 VTAIL.n287 B 0.024175f
C406 VTAIL.n288 B 0.024175f
C407 VTAIL.n289 B 0.010529f
C408 VTAIL.n290 B 0.010228f
C409 VTAIL.n291 B 0.019034f
C410 VTAIL.n292 B 0.019034f
C411 VTAIL.n293 B 0.010228f
C412 VTAIL.n294 B 0.01083f
C413 VTAIL.n295 B 0.024175f
C414 VTAIL.n296 B 0.024175f
C415 VTAIL.n297 B 0.01083f
C416 VTAIL.n298 B 0.010228f
C417 VTAIL.n299 B 0.019034f
C418 VTAIL.n300 B 0.019034f
C419 VTAIL.n301 B 0.010228f
C420 VTAIL.n302 B 0.01083f
C421 VTAIL.n303 B 0.024175f
C422 VTAIL.n304 B 0.049838f
C423 VTAIL.n305 B 0.01083f
C424 VTAIL.n306 B 0.010228f
C425 VTAIL.n307 B 0.041136f
C426 VTAIL.n308 B 0.027539f
C427 VTAIL.n309 B 1.64947f
C428 VTAIL.n310 B 0.025341f
C429 VTAIL.n311 B 0.019034f
C430 VTAIL.n312 B 0.010228f
C431 VTAIL.n313 B 0.024175f
C432 VTAIL.n314 B 0.01083f
C433 VTAIL.n315 B 0.019034f
C434 VTAIL.n316 B 0.010228f
C435 VTAIL.n317 B 0.024175f
C436 VTAIL.n318 B 0.01083f
C437 VTAIL.n319 B 0.019034f
C438 VTAIL.n320 B 0.010529f
C439 VTAIL.n321 B 0.024175f
C440 VTAIL.n322 B 0.010228f
C441 VTAIL.n323 B 0.01083f
C442 VTAIL.n324 B 0.019034f
C443 VTAIL.n325 B 0.010228f
C444 VTAIL.n326 B 0.024175f
C445 VTAIL.n327 B 0.01083f
C446 VTAIL.n328 B 0.019034f
C447 VTAIL.n329 B 0.010228f
C448 VTAIL.n330 B 0.024175f
C449 VTAIL.n331 B 0.01083f
C450 VTAIL.n332 B 0.019034f
C451 VTAIL.n333 B 0.010228f
C452 VTAIL.n334 B 0.024175f
C453 VTAIL.n335 B 0.01083f
C454 VTAIL.n336 B 0.019034f
C455 VTAIL.n337 B 0.010228f
C456 VTAIL.n338 B 0.024175f
C457 VTAIL.n339 B 0.01083f
C458 VTAIL.n340 B 0.019034f
C459 VTAIL.n341 B 0.010228f
C460 VTAIL.n342 B 0.018132f
C461 VTAIL.n343 B 0.014281f
C462 VTAIL.t2 B 0.040067f
C463 VTAIL.n344 B 0.139081f
C464 VTAIL.n345 B 1.51142f
C465 VTAIL.n346 B 0.010228f
C466 VTAIL.n347 B 0.01083f
C467 VTAIL.n348 B 0.024175f
C468 VTAIL.n349 B 0.024175f
C469 VTAIL.n350 B 0.01083f
C470 VTAIL.n351 B 0.010228f
C471 VTAIL.n352 B 0.019034f
C472 VTAIL.n353 B 0.019034f
C473 VTAIL.n354 B 0.010228f
C474 VTAIL.n355 B 0.01083f
C475 VTAIL.n356 B 0.024175f
C476 VTAIL.n357 B 0.024175f
C477 VTAIL.n358 B 0.01083f
C478 VTAIL.n359 B 0.010228f
C479 VTAIL.n360 B 0.019034f
C480 VTAIL.n361 B 0.019034f
C481 VTAIL.n362 B 0.010228f
C482 VTAIL.n363 B 0.01083f
C483 VTAIL.n364 B 0.024175f
C484 VTAIL.n365 B 0.024175f
C485 VTAIL.n366 B 0.01083f
C486 VTAIL.n367 B 0.010228f
C487 VTAIL.n368 B 0.019034f
C488 VTAIL.n369 B 0.019034f
C489 VTAIL.n370 B 0.010228f
C490 VTAIL.n371 B 0.01083f
C491 VTAIL.n372 B 0.024175f
C492 VTAIL.n373 B 0.024175f
C493 VTAIL.n374 B 0.01083f
C494 VTAIL.n375 B 0.010228f
C495 VTAIL.n376 B 0.019034f
C496 VTAIL.n377 B 0.019034f
C497 VTAIL.n378 B 0.010228f
C498 VTAIL.n379 B 0.01083f
C499 VTAIL.n380 B 0.024175f
C500 VTAIL.n381 B 0.024175f
C501 VTAIL.n382 B 0.01083f
C502 VTAIL.n383 B 0.010228f
C503 VTAIL.n384 B 0.019034f
C504 VTAIL.n385 B 0.019034f
C505 VTAIL.n386 B 0.010228f
C506 VTAIL.n387 B 0.01083f
C507 VTAIL.n388 B 0.024175f
C508 VTAIL.n389 B 0.024175f
C509 VTAIL.n390 B 0.024175f
C510 VTAIL.n391 B 0.010529f
C511 VTAIL.n392 B 0.010228f
C512 VTAIL.n393 B 0.019034f
C513 VTAIL.n394 B 0.019034f
C514 VTAIL.n395 B 0.010228f
C515 VTAIL.n396 B 0.01083f
C516 VTAIL.n397 B 0.024175f
C517 VTAIL.n398 B 0.024175f
C518 VTAIL.n399 B 0.01083f
C519 VTAIL.n400 B 0.010228f
C520 VTAIL.n401 B 0.019034f
C521 VTAIL.n402 B 0.019034f
C522 VTAIL.n403 B 0.010228f
C523 VTAIL.n404 B 0.01083f
C524 VTAIL.n405 B 0.024175f
C525 VTAIL.n406 B 0.049838f
C526 VTAIL.n407 B 0.01083f
C527 VTAIL.n408 B 0.010228f
C528 VTAIL.n409 B 0.041136f
C529 VTAIL.n410 B 0.027539f
C530 VTAIL.n411 B 1.64947f
C531 VTAIL.t1 B 0.272698f
C532 VTAIL.t5 B 0.272698f
C533 VTAIL.n412 B 2.41984f
C534 VTAIL.n413 B 0.61518f
C535 VTAIL.n414 B 0.025341f
C536 VTAIL.n415 B 0.019034f
C537 VTAIL.n416 B 0.010228f
C538 VTAIL.n417 B 0.024175f
C539 VTAIL.n418 B 0.01083f
C540 VTAIL.n419 B 0.019034f
C541 VTAIL.n420 B 0.010228f
C542 VTAIL.n421 B 0.024175f
C543 VTAIL.n422 B 0.01083f
C544 VTAIL.n423 B 0.019034f
C545 VTAIL.n424 B 0.010529f
C546 VTAIL.n425 B 0.024175f
C547 VTAIL.n426 B 0.010228f
C548 VTAIL.n427 B 0.01083f
C549 VTAIL.n428 B 0.019034f
C550 VTAIL.n429 B 0.010228f
C551 VTAIL.n430 B 0.024175f
C552 VTAIL.n431 B 0.01083f
C553 VTAIL.n432 B 0.019034f
C554 VTAIL.n433 B 0.010228f
C555 VTAIL.n434 B 0.024175f
C556 VTAIL.n435 B 0.01083f
C557 VTAIL.n436 B 0.019034f
C558 VTAIL.n437 B 0.010228f
C559 VTAIL.n438 B 0.024175f
C560 VTAIL.n439 B 0.01083f
C561 VTAIL.n440 B 0.019034f
C562 VTAIL.n441 B 0.010228f
C563 VTAIL.n442 B 0.024175f
C564 VTAIL.n443 B 0.01083f
C565 VTAIL.n444 B 0.019034f
C566 VTAIL.n445 B 0.010228f
C567 VTAIL.n446 B 0.018132f
C568 VTAIL.n447 B 0.014281f
C569 VTAIL.t6 B 0.040067f
C570 VTAIL.n448 B 0.139081f
C571 VTAIL.n449 B 1.51142f
C572 VTAIL.n450 B 0.010228f
C573 VTAIL.n451 B 0.01083f
C574 VTAIL.n452 B 0.024175f
C575 VTAIL.n453 B 0.024175f
C576 VTAIL.n454 B 0.01083f
C577 VTAIL.n455 B 0.010228f
C578 VTAIL.n456 B 0.019034f
C579 VTAIL.n457 B 0.019034f
C580 VTAIL.n458 B 0.010228f
C581 VTAIL.n459 B 0.01083f
C582 VTAIL.n460 B 0.024175f
C583 VTAIL.n461 B 0.024175f
C584 VTAIL.n462 B 0.01083f
C585 VTAIL.n463 B 0.010228f
C586 VTAIL.n464 B 0.019034f
C587 VTAIL.n465 B 0.019034f
C588 VTAIL.n466 B 0.010228f
C589 VTAIL.n467 B 0.01083f
C590 VTAIL.n468 B 0.024175f
C591 VTAIL.n469 B 0.024175f
C592 VTAIL.n470 B 0.01083f
C593 VTAIL.n471 B 0.010228f
C594 VTAIL.n472 B 0.019034f
C595 VTAIL.n473 B 0.019034f
C596 VTAIL.n474 B 0.010228f
C597 VTAIL.n475 B 0.01083f
C598 VTAIL.n476 B 0.024175f
C599 VTAIL.n477 B 0.024175f
C600 VTAIL.n478 B 0.01083f
C601 VTAIL.n479 B 0.010228f
C602 VTAIL.n480 B 0.019034f
C603 VTAIL.n481 B 0.019034f
C604 VTAIL.n482 B 0.010228f
C605 VTAIL.n483 B 0.01083f
C606 VTAIL.n484 B 0.024175f
C607 VTAIL.n485 B 0.024175f
C608 VTAIL.n486 B 0.01083f
C609 VTAIL.n487 B 0.010228f
C610 VTAIL.n488 B 0.019034f
C611 VTAIL.n489 B 0.019034f
C612 VTAIL.n490 B 0.010228f
C613 VTAIL.n491 B 0.01083f
C614 VTAIL.n492 B 0.024175f
C615 VTAIL.n493 B 0.024175f
C616 VTAIL.n494 B 0.024175f
C617 VTAIL.n495 B 0.010529f
C618 VTAIL.n496 B 0.010228f
C619 VTAIL.n497 B 0.019034f
C620 VTAIL.n498 B 0.019034f
C621 VTAIL.n499 B 0.010228f
C622 VTAIL.n500 B 0.01083f
C623 VTAIL.n501 B 0.024175f
C624 VTAIL.n502 B 0.024175f
C625 VTAIL.n503 B 0.01083f
C626 VTAIL.n504 B 0.010228f
C627 VTAIL.n505 B 0.019034f
C628 VTAIL.n506 B 0.019034f
C629 VTAIL.n507 B 0.010228f
C630 VTAIL.n508 B 0.01083f
C631 VTAIL.n509 B 0.024175f
C632 VTAIL.n510 B 0.049838f
C633 VTAIL.n511 B 0.01083f
C634 VTAIL.n512 B 0.010228f
C635 VTAIL.n513 B 0.041136f
C636 VTAIL.n514 B 0.027539f
C637 VTAIL.n515 B 0.252306f
C638 VTAIL.n516 B 0.025341f
C639 VTAIL.n517 B 0.019034f
C640 VTAIL.n518 B 0.010228f
C641 VTAIL.n519 B 0.024175f
C642 VTAIL.n520 B 0.01083f
C643 VTAIL.n521 B 0.019034f
C644 VTAIL.n522 B 0.010228f
C645 VTAIL.n523 B 0.024175f
C646 VTAIL.n524 B 0.01083f
C647 VTAIL.n525 B 0.019034f
C648 VTAIL.n526 B 0.010529f
C649 VTAIL.n527 B 0.024175f
C650 VTAIL.n528 B 0.010228f
C651 VTAIL.n529 B 0.01083f
C652 VTAIL.n530 B 0.019034f
C653 VTAIL.n531 B 0.010228f
C654 VTAIL.n532 B 0.024175f
C655 VTAIL.n533 B 0.01083f
C656 VTAIL.n534 B 0.019034f
C657 VTAIL.n535 B 0.010228f
C658 VTAIL.n536 B 0.024175f
C659 VTAIL.n537 B 0.01083f
C660 VTAIL.n538 B 0.019034f
C661 VTAIL.n539 B 0.010228f
C662 VTAIL.n540 B 0.024175f
C663 VTAIL.n541 B 0.01083f
C664 VTAIL.n542 B 0.019034f
C665 VTAIL.n543 B 0.010228f
C666 VTAIL.n544 B 0.024175f
C667 VTAIL.n545 B 0.01083f
C668 VTAIL.n546 B 0.019034f
C669 VTAIL.n547 B 0.010228f
C670 VTAIL.n548 B 0.018132f
C671 VTAIL.n549 B 0.014281f
C672 VTAIL.t10 B 0.040067f
C673 VTAIL.n550 B 0.139081f
C674 VTAIL.n551 B 1.51142f
C675 VTAIL.n552 B 0.010228f
C676 VTAIL.n553 B 0.01083f
C677 VTAIL.n554 B 0.024175f
C678 VTAIL.n555 B 0.024175f
C679 VTAIL.n556 B 0.01083f
C680 VTAIL.n557 B 0.010228f
C681 VTAIL.n558 B 0.019034f
C682 VTAIL.n559 B 0.019034f
C683 VTAIL.n560 B 0.010228f
C684 VTAIL.n561 B 0.01083f
C685 VTAIL.n562 B 0.024175f
C686 VTAIL.n563 B 0.024175f
C687 VTAIL.n564 B 0.01083f
C688 VTAIL.n565 B 0.010228f
C689 VTAIL.n566 B 0.019034f
C690 VTAIL.n567 B 0.019034f
C691 VTAIL.n568 B 0.010228f
C692 VTAIL.n569 B 0.01083f
C693 VTAIL.n570 B 0.024175f
C694 VTAIL.n571 B 0.024175f
C695 VTAIL.n572 B 0.01083f
C696 VTAIL.n573 B 0.010228f
C697 VTAIL.n574 B 0.019034f
C698 VTAIL.n575 B 0.019034f
C699 VTAIL.n576 B 0.010228f
C700 VTAIL.n577 B 0.01083f
C701 VTAIL.n578 B 0.024175f
C702 VTAIL.n579 B 0.024175f
C703 VTAIL.n580 B 0.01083f
C704 VTAIL.n581 B 0.010228f
C705 VTAIL.n582 B 0.019034f
C706 VTAIL.n583 B 0.019034f
C707 VTAIL.n584 B 0.010228f
C708 VTAIL.n585 B 0.01083f
C709 VTAIL.n586 B 0.024175f
C710 VTAIL.n587 B 0.024175f
C711 VTAIL.n588 B 0.01083f
C712 VTAIL.n589 B 0.010228f
C713 VTAIL.n590 B 0.019034f
C714 VTAIL.n591 B 0.019034f
C715 VTAIL.n592 B 0.010228f
C716 VTAIL.n593 B 0.01083f
C717 VTAIL.n594 B 0.024175f
C718 VTAIL.n595 B 0.024175f
C719 VTAIL.n596 B 0.024175f
C720 VTAIL.n597 B 0.010529f
C721 VTAIL.n598 B 0.010228f
C722 VTAIL.n599 B 0.019034f
C723 VTAIL.n600 B 0.019034f
C724 VTAIL.n601 B 0.010228f
C725 VTAIL.n602 B 0.01083f
C726 VTAIL.n603 B 0.024175f
C727 VTAIL.n604 B 0.024175f
C728 VTAIL.n605 B 0.01083f
C729 VTAIL.n606 B 0.010228f
C730 VTAIL.n607 B 0.019034f
C731 VTAIL.n608 B 0.019034f
C732 VTAIL.n609 B 0.010228f
C733 VTAIL.n610 B 0.01083f
C734 VTAIL.n611 B 0.024175f
C735 VTAIL.n612 B 0.049838f
C736 VTAIL.n613 B 0.01083f
C737 VTAIL.n614 B 0.010228f
C738 VTAIL.n615 B 0.041136f
C739 VTAIL.n616 B 0.027539f
C740 VTAIL.n617 B 0.252306f
C741 VTAIL.t12 B 0.272698f
C742 VTAIL.t14 B 0.272698f
C743 VTAIL.n618 B 2.41984f
C744 VTAIL.n619 B 0.61518f
C745 VTAIL.n620 B 0.025341f
C746 VTAIL.n621 B 0.019034f
C747 VTAIL.n622 B 0.010228f
C748 VTAIL.n623 B 0.024175f
C749 VTAIL.n624 B 0.01083f
C750 VTAIL.n625 B 0.019034f
C751 VTAIL.n626 B 0.010228f
C752 VTAIL.n627 B 0.024175f
C753 VTAIL.n628 B 0.01083f
C754 VTAIL.n629 B 0.019034f
C755 VTAIL.n630 B 0.010529f
C756 VTAIL.n631 B 0.024175f
C757 VTAIL.n632 B 0.010228f
C758 VTAIL.n633 B 0.01083f
C759 VTAIL.n634 B 0.019034f
C760 VTAIL.n635 B 0.010228f
C761 VTAIL.n636 B 0.024175f
C762 VTAIL.n637 B 0.01083f
C763 VTAIL.n638 B 0.019034f
C764 VTAIL.n639 B 0.010228f
C765 VTAIL.n640 B 0.024175f
C766 VTAIL.n641 B 0.01083f
C767 VTAIL.n642 B 0.019034f
C768 VTAIL.n643 B 0.010228f
C769 VTAIL.n644 B 0.024175f
C770 VTAIL.n645 B 0.01083f
C771 VTAIL.n646 B 0.019034f
C772 VTAIL.n647 B 0.010228f
C773 VTAIL.n648 B 0.024175f
C774 VTAIL.n649 B 0.01083f
C775 VTAIL.n650 B 0.019034f
C776 VTAIL.n651 B 0.010228f
C777 VTAIL.n652 B 0.018132f
C778 VTAIL.n653 B 0.014281f
C779 VTAIL.t9 B 0.040067f
C780 VTAIL.n654 B 0.139081f
C781 VTAIL.n655 B 1.51142f
C782 VTAIL.n656 B 0.010228f
C783 VTAIL.n657 B 0.01083f
C784 VTAIL.n658 B 0.024175f
C785 VTAIL.n659 B 0.024175f
C786 VTAIL.n660 B 0.01083f
C787 VTAIL.n661 B 0.010228f
C788 VTAIL.n662 B 0.019034f
C789 VTAIL.n663 B 0.019034f
C790 VTAIL.n664 B 0.010228f
C791 VTAIL.n665 B 0.01083f
C792 VTAIL.n666 B 0.024175f
C793 VTAIL.n667 B 0.024175f
C794 VTAIL.n668 B 0.01083f
C795 VTAIL.n669 B 0.010228f
C796 VTAIL.n670 B 0.019034f
C797 VTAIL.n671 B 0.019034f
C798 VTAIL.n672 B 0.010228f
C799 VTAIL.n673 B 0.01083f
C800 VTAIL.n674 B 0.024175f
C801 VTAIL.n675 B 0.024175f
C802 VTAIL.n676 B 0.01083f
C803 VTAIL.n677 B 0.010228f
C804 VTAIL.n678 B 0.019034f
C805 VTAIL.n679 B 0.019034f
C806 VTAIL.n680 B 0.010228f
C807 VTAIL.n681 B 0.01083f
C808 VTAIL.n682 B 0.024175f
C809 VTAIL.n683 B 0.024175f
C810 VTAIL.n684 B 0.01083f
C811 VTAIL.n685 B 0.010228f
C812 VTAIL.n686 B 0.019034f
C813 VTAIL.n687 B 0.019034f
C814 VTAIL.n688 B 0.010228f
C815 VTAIL.n689 B 0.01083f
C816 VTAIL.n690 B 0.024175f
C817 VTAIL.n691 B 0.024175f
C818 VTAIL.n692 B 0.01083f
C819 VTAIL.n693 B 0.010228f
C820 VTAIL.n694 B 0.019034f
C821 VTAIL.n695 B 0.019034f
C822 VTAIL.n696 B 0.010228f
C823 VTAIL.n697 B 0.01083f
C824 VTAIL.n698 B 0.024175f
C825 VTAIL.n699 B 0.024175f
C826 VTAIL.n700 B 0.024175f
C827 VTAIL.n701 B 0.010529f
C828 VTAIL.n702 B 0.010228f
C829 VTAIL.n703 B 0.019034f
C830 VTAIL.n704 B 0.019034f
C831 VTAIL.n705 B 0.010228f
C832 VTAIL.n706 B 0.01083f
C833 VTAIL.n707 B 0.024175f
C834 VTAIL.n708 B 0.024175f
C835 VTAIL.n709 B 0.01083f
C836 VTAIL.n710 B 0.010228f
C837 VTAIL.n711 B 0.019034f
C838 VTAIL.n712 B 0.019034f
C839 VTAIL.n713 B 0.010228f
C840 VTAIL.n714 B 0.01083f
C841 VTAIL.n715 B 0.024175f
C842 VTAIL.n716 B 0.049838f
C843 VTAIL.n717 B 0.01083f
C844 VTAIL.n718 B 0.010228f
C845 VTAIL.n719 B 0.041136f
C846 VTAIL.n720 B 0.027539f
C847 VTAIL.n721 B 1.64947f
C848 VTAIL.n722 B 0.025341f
C849 VTAIL.n723 B 0.019034f
C850 VTAIL.n724 B 0.010228f
C851 VTAIL.n725 B 0.024175f
C852 VTAIL.n726 B 0.01083f
C853 VTAIL.n727 B 0.019034f
C854 VTAIL.n728 B 0.010228f
C855 VTAIL.n729 B 0.024175f
C856 VTAIL.n730 B 0.01083f
C857 VTAIL.n731 B 0.019034f
C858 VTAIL.n732 B 0.010529f
C859 VTAIL.n733 B 0.024175f
C860 VTAIL.n734 B 0.01083f
C861 VTAIL.n735 B 0.019034f
C862 VTAIL.n736 B 0.010228f
C863 VTAIL.n737 B 0.024175f
C864 VTAIL.n738 B 0.01083f
C865 VTAIL.n739 B 0.019034f
C866 VTAIL.n740 B 0.010228f
C867 VTAIL.n741 B 0.024175f
C868 VTAIL.n742 B 0.01083f
C869 VTAIL.n743 B 0.019034f
C870 VTAIL.n744 B 0.010228f
C871 VTAIL.n745 B 0.024175f
C872 VTAIL.n746 B 0.01083f
C873 VTAIL.n747 B 0.019034f
C874 VTAIL.n748 B 0.010228f
C875 VTAIL.n749 B 0.024175f
C876 VTAIL.n750 B 0.01083f
C877 VTAIL.n751 B 0.019034f
C878 VTAIL.n752 B 0.010228f
C879 VTAIL.n753 B 0.018132f
C880 VTAIL.n754 B 0.014281f
C881 VTAIL.t15 B 0.040067f
C882 VTAIL.n755 B 0.139081f
C883 VTAIL.n756 B 1.51142f
C884 VTAIL.n757 B 0.010228f
C885 VTAIL.n758 B 0.01083f
C886 VTAIL.n759 B 0.024175f
C887 VTAIL.n760 B 0.024175f
C888 VTAIL.n761 B 0.01083f
C889 VTAIL.n762 B 0.010228f
C890 VTAIL.n763 B 0.019034f
C891 VTAIL.n764 B 0.019034f
C892 VTAIL.n765 B 0.010228f
C893 VTAIL.n766 B 0.01083f
C894 VTAIL.n767 B 0.024175f
C895 VTAIL.n768 B 0.024175f
C896 VTAIL.n769 B 0.01083f
C897 VTAIL.n770 B 0.010228f
C898 VTAIL.n771 B 0.019034f
C899 VTAIL.n772 B 0.019034f
C900 VTAIL.n773 B 0.010228f
C901 VTAIL.n774 B 0.01083f
C902 VTAIL.n775 B 0.024175f
C903 VTAIL.n776 B 0.024175f
C904 VTAIL.n777 B 0.01083f
C905 VTAIL.n778 B 0.010228f
C906 VTAIL.n779 B 0.019034f
C907 VTAIL.n780 B 0.019034f
C908 VTAIL.n781 B 0.010228f
C909 VTAIL.n782 B 0.01083f
C910 VTAIL.n783 B 0.024175f
C911 VTAIL.n784 B 0.024175f
C912 VTAIL.n785 B 0.01083f
C913 VTAIL.n786 B 0.010228f
C914 VTAIL.n787 B 0.019034f
C915 VTAIL.n788 B 0.019034f
C916 VTAIL.n789 B 0.010228f
C917 VTAIL.n790 B 0.01083f
C918 VTAIL.n791 B 0.024175f
C919 VTAIL.n792 B 0.024175f
C920 VTAIL.n793 B 0.01083f
C921 VTAIL.n794 B 0.010228f
C922 VTAIL.n795 B 0.019034f
C923 VTAIL.n796 B 0.019034f
C924 VTAIL.n797 B 0.010228f
C925 VTAIL.n798 B 0.010228f
C926 VTAIL.n799 B 0.01083f
C927 VTAIL.n800 B 0.024175f
C928 VTAIL.n801 B 0.024175f
C929 VTAIL.n802 B 0.024175f
C930 VTAIL.n803 B 0.010529f
C931 VTAIL.n804 B 0.010228f
C932 VTAIL.n805 B 0.019034f
C933 VTAIL.n806 B 0.019034f
C934 VTAIL.n807 B 0.010228f
C935 VTAIL.n808 B 0.01083f
C936 VTAIL.n809 B 0.024175f
C937 VTAIL.n810 B 0.024175f
C938 VTAIL.n811 B 0.01083f
C939 VTAIL.n812 B 0.010228f
C940 VTAIL.n813 B 0.019034f
C941 VTAIL.n814 B 0.019034f
C942 VTAIL.n815 B 0.010228f
C943 VTAIL.n816 B 0.01083f
C944 VTAIL.n817 B 0.024175f
C945 VTAIL.n818 B 0.049838f
C946 VTAIL.n819 B 0.01083f
C947 VTAIL.n820 B 0.010228f
C948 VTAIL.n821 B 0.041136f
C949 VTAIL.n822 B 0.027539f
C950 VTAIL.n823 B 1.6459f
C951 VDD1.t6 B 0.381502f
C952 VDD1.t3 B 0.381502f
C953 VDD1.n0 B 3.49278f
C954 VDD1.t0 B 0.381502f
C955 VDD1.t7 B 0.381502f
C956 VDD1.n1 B 3.49127f
C957 VDD1.t4 B 0.381502f
C958 VDD1.t1 B 0.381502f
C959 VDD1.n2 B 3.49127f
C960 VDD1.n3 B 4.59875f
C961 VDD1.t5 B 0.381502f
C962 VDD1.t2 B 0.381502f
C963 VDD1.n4 B 3.47294f
C964 VDD1.n5 B 4.0498f
C965 VP.t6 B 3.07101f
C966 VP.n0 B 1.12475f
C967 VP.n1 B 0.01701f
C968 VP.n2 B 0.027201f
C969 VP.n3 B 0.01701f
C970 VP.n4 B 0.024658f
C971 VP.n5 B 0.01701f
C972 VP.n6 B 0.024831f
C973 VP.n7 B 0.01701f
C974 VP.n8 B 0.023093f
C975 VP.n9 B 0.01701f
C976 VP.n10 B 0.022461f
C977 VP.n11 B 0.01701f
C978 VP.n12 B 0.021527f
C979 VP.t5 B 3.07101f
C980 VP.n13 B 1.12475f
C981 VP.n14 B 0.01701f
C982 VP.n15 B 0.027201f
C983 VP.n16 B 0.01701f
C984 VP.n17 B 0.024658f
C985 VP.n18 B 0.01701f
C986 VP.n19 B 0.024831f
C987 VP.n20 B 0.01701f
C988 VP.n21 B 0.023093f
C989 VP.t4 B 3.32703f
C990 VP.t2 B 3.07101f
C991 VP.n22 B 1.11692f
C992 VP.n23 B 1.06703f
C993 VP.n24 B 0.213061f
C994 VP.n25 B 0.01701f
C995 VP.n26 B 0.031702f
C996 VP.n27 B 0.031702f
C997 VP.n28 B 0.024831f
C998 VP.n29 B 0.01701f
C999 VP.n30 B 0.01701f
C1000 VP.n31 B 0.01701f
C1001 VP.n32 B 0.031702f
C1002 VP.n33 B 0.031702f
C1003 VP.t0 B 3.07101f
C1004 VP.n34 B 1.05849f
C1005 VP.n35 B 0.023093f
C1006 VP.n36 B 0.01701f
C1007 VP.n37 B 0.01701f
C1008 VP.n38 B 0.01701f
C1009 VP.n39 B 0.031702f
C1010 VP.n40 B 0.031702f
C1011 VP.n41 B 0.022461f
C1012 VP.n42 B 0.01701f
C1013 VP.n43 B 0.01701f
C1014 VP.n44 B 0.01701f
C1015 VP.n45 B 0.031702f
C1016 VP.n46 B 0.031702f
C1017 VP.n47 B 0.021527f
C1018 VP.n48 B 0.027453f
C1019 VP.n49 B 1.26371f
C1020 VP.t7 B 3.07101f
C1021 VP.n50 B 1.12475f
C1022 VP.n51 B 1.27383f
C1023 VP.n52 B 0.027453f
C1024 VP.n53 B 0.01701f
C1025 VP.n54 B 0.031702f
C1026 VP.n55 B 0.031702f
C1027 VP.n56 B 0.027201f
C1028 VP.n57 B 0.01701f
C1029 VP.n58 B 0.01701f
C1030 VP.n59 B 0.01701f
C1031 VP.n60 B 0.031702f
C1032 VP.n61 B 0.031702f
C1033 VP.t3 B 3.07101f
C1034 VP.n62 B 1.05849f
C1035 VP.n63 B 0.024658f
C1036 VP.n64 B 0.01701f
C1037 VP.n65 B 0.01701f
C1038 VP.n66 B 0.01701f
C1039 VP.n67 B 0.031702f
C1040 VP.n68 B 0.031702f
C1041 VP.n69 B 0.024831f
C1042 VP.n70 B 0.01701f
C1043 VP.n71 B 0.01701f
C1044 VP.n72 B 0.01701f
C1045 VP.n73 B 0.031702f
C1046 VP.n74 B 0.031702f
C1047 VP.t1 B 3.07101f
C1048 VP.n75 B 1.05849f
C1049 VP.n76 B 0.023093f
C1050 VP.n77 B 0.01701f
C1051 VP.n78 B 0.01701f
C1052 VP.n79 B 0.01701f
C1053 VP.n80 B 0.031702f
C1054 VP.n81 B 0.031702f
C1055 VP.n82 B 0.022461f
C1056 VP.n83 B 0.01701f
C1057 VP.n84 B 0.01701f
C1058 VP.n85 B 0.01701f
C1059 VP.n86 B 0.031702f
C1060 VP.n87 B 0.031702f
C1061 VP.n88 B 0.021527f
C1062 VP.n89 B 0.027453f
C1063 VP.n90 B 0.047533f
.ends

