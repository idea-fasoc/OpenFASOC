* NGSPICE file created from diff_pair_sample_1710.ext - technology: sky130A

.subckt diff_pair_sample_1710 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t3 VP.t0 VTAIL.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=3.2901 pd=20.27 as=7.7766 ps=40.66 w=19.94 l=0.83
X1 VTAIL.t6 VP.t1 VDD1.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=7.7766 pd=40.66 as=3.2901 ps=20.27 w=19.94 l=0.83
X2 VTAIL.t4 VP.t2 VDD1.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=7.7766 pd=40.66 as=3.2901 ps=20.27 w=19.94 l=0.83
X3 B.t17 B.t15 B.t16 B.t5 sky130_fd_pr__nfet_01v8 ad=7.7766 pd=40.66 as=0 ps=0 w=19.94 l=0.83
X4 VDD2.t3 VN.t0 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=3.2901 pd=20.27 as=7.7766 ps=40.66 w=19.94 l=0.83
X5 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=7.7766 pd=40.66 as=0 ps=0 w=19.94 l=0.83
X6 VTAIL.t0 VN.t1 VDD2.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=7.7766 pd=40.66 as=3.2901 ps=20.27 w=19.94 l=0.83
X7 VDD2.t1 VN.t2 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=3.2901 pd=20.27 as=7.7766 ps=40.66 w=19.94 l=0.83
X8 VDD1.t0 VP.t3 VTAIL.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=3.2901 pd=20.27 as=7.7766 ps=40.66 w=19.94 l=0.83
X9 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=7.7766 pd=40.66 as=0 ps=0 w=19.94 l=0.83
X10 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=7.7766 pd=40.66 as=0 ps=0 w=19.94 l=0.83
X11 VTAIL.t1 VN.t3 VDD2.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=7.7766 pd=40.66 as=3.2901 ps=20.27 w=19.94 l=0.83
R0 VP.n1 VP.t1 647.888
R1 VP.n1 VP.t0 647.837
R2 VP.n3 VP.t2 626.89
R3 VP.n5 VP.t3 626.89
R4 VP.n6 VP.n5 161.3
R5 VP.n4 VP.n0 161.3
R6 VP.n3 VP.n2 161.3
R7 VP.n2 VP.n1 91.5787
R8 VP.n4 VP.n3 24.1005
R9 VP.n5 VP.n4 24.1005
R10 VP.n2 VP.n0 0.189894
R11 VP.n6 VP.n0 0.189894
R12 VP VP.n6 0.0516364
R13 VTAIL.n6 VTAIL.t7 42.969
R14 VTAIL.n5 VTAIL.t6 42.969
R15 VTAIL.n4 VTAIL.t3 42.969
R16 VTAIL.n3 VTAIL.t0 42.969
R17 VTAIL.n7 VTAIL.t2 42.9688
R18 VTAIL.n0 VTAIL.t1 42.9688
R19 VTAIL.n1 VTAIL.t5 42.9688
R20 VTAIL.n2 VTAIL.t4 42.9688
R21 VTAIL.n7 VTAIL.n6 30.5565
R22 VTAIL.n3 VTAIL.n2 30.5565
R23 VTAIL.n4 VTAIL.n3 1.0005
R24 VTAIL.n6 VTAIL.n5 1.0005
R25 VTAIL.n2 VTAIL.n1 1.0005
R26 VTAIL VTAIL.n0 0.55869
R27 VTAIL.n5 VTAIL.n4 0.470328
R28 VTAIL.n1 VTAIL.n0 0.470328
R29 VTAIL VTAIL.n7 0.44231
R30 VDD1 VDD1.n1 103.085
R31 VDD1 VDD1.n0 58.713
R32 VDD1.n0 VDD1.t2 0.993479
R33 VDD1.n0 VDD1.t3 0.993479
R34 VDD1.n1 VDD1.t1 0.993479
R35 VDD1.n1 VDD1.t0 0.993479
R36 B.n71 B.t12 780.597
R37 B.n77 B.t8 780.597
R38 B.n187 B.t4 780.597
R39 B.n179 B.t15 780.597
R40 B.n579 B.n112 585
R41 B.n112 B.n37 585
R42 B.n581 B.n580 585
R43 B.n583 B.n111 585
R44 B.n586 B.n585 585
R45 B.n587 B.n110 585
R46 B.n589 B.n588 585
R47 B.n591 B.n109 585
R48 B.n594 B.n593 585
R49 B.n595 B.n108 585
R50 B.n597 B.n596 585
R51 B.n599 B.n107 585
R52 B.n602 B.n601 585
R53 B.n603 B.n106 585
R54 B.n605 B.n604 585
R55 B.n607 B.n105 585
R56 B.n610 B.n609 585
R57 B.n611 B.n104 585
R58 B.n613 B.n612 585
R59 B.n615 B.n103 585
R60 B.n618 B.n617 585
R61 B.n619 B.n102 585
R62 B.n621 B.n620 585
R63 B.n623 B.n101 585
R64 B.n626 B.n625 585
R65 B.n627 B.n100 585
R66 B.n629 B.n628 585
R67 B.n631 B.n99 585
R68 B.n634 B.n633 585
R69 B.n635 B.n98 585
R70 B.n637 B.n636 585
R71 B.n639 B.n97 585
R72 B.n642 B.n641 585
R73 B.n643 B.n96 585
R74 B.n645 B.n644 585
R75 B.n647 B.n95 585
R76 B.n650 B.n649 585
R77 B.n651 B.n94 585
R78 B.n653 B.n652 585
R79 B.n655 B.n93 585
R80 B.n658 B.n657 585
R81 B.n659 B.n92 585
R82 B.n661 B.n660 585
R83 B.n663 B.n91 585
R84 B.n666 B.n665 585
R85 B.n667 B.n90 585
R86 B.n669 B.n668 585
R87 B.n671 B.n89 585
R88 B.n674 B.n673 585
R89 B.n675 B.n88 585
R90 B.n677 B.n676 585
R91 B.n679 B.n87 585
R92 B.n682 B.n681 585
R93 B.n683 B.n86 585
R94 B.n685 B.n684 585
R95 B.n687 B.n85 585
R96 B.n690 B.n689 585
R97 B.n691 B.n84 585
R98 B.n693 B.n692 585
R99 B.n695 B.n83 585
R100 B.n698 B.n697 585
R101 B.n699 B.n82 585
R102 B.n701 B.n700 585
R103 B.n703 B.n81 585
R104 B.n705 B.n704 585
R105 B.n707 B.n706 585
R106 B.n710 B.n709 585
R107 B.n711 B.n76 585
R108 B.n713 B.n712 585
R109 B.n715 B.n75 585
R110 B.n718 B.n717 585
R111 B.n719 B.n74 585
R112 B.n721 B.n720 585
R113 B.n723 B.n73 585
R114 B.n726 B.n725 585
R115 B.n728 B.n70 585
R116 B.n730 B.n729 585
R117 B.n732 B.n69 585
R118 B.n735 B.n734 585
R119 B.n736 B.n68 585
R120 B.n738 B.n737 585
R121 B.n740 B.n67 585
R122 B.n743 B.n742 585
R123 B.n744 B.n66 585
R124 B.n746 B.n745 585
R125 B.n748 B.n65 585
R126 B.n751 B.n750 585
R127 B.n752 B.n64 585
R128 B.n754 B.n753 585
R129 B.n756 B.n63 585
R130 B.n759 B.n758 585
R131 B.n760 B.n62 585
R132 B.n762 B.n761 585
R133 B.n764 B.n61 585
R134 B.n767 B.n766 585
R135 B.n768 B.n60 585
R136 B.n770 B.n769 585
R137 B.n772 B.n59 585
R138 B.n775 B.n774 585
R139 B.n776 B.n58 585
R140 B.n778 B.n777 585
R141 B.n780 B.n57 585
R142 B.n783 B.n782 585
R143 B.n784 B.n56 585
R144 B.n786 B.n785 585
R145 B.n788 B.n55 585
R146 B.n791 B.n790 585
R147 B.n792 B.n54 585
R148 B.n794 B.n793 585
R149 B.n796 B.n53 585
R150 B.n799 B.n798 585
R151 B.n800 B.n52 585
R152 B.n802 B.n801 585
R153 B.n804 B.n51 585
R154 B.n807 B.n806 585
R155 B.n808 B.n50 585
R156 B.n810 B.n809 585
R157 B.n812 B.n49 585
R158 B.n815 B.n814 585
R159 B.n816 B.n48 585
R160 B.n818 B.n817 585
R161 B.n820 B.n47 585
R162 B.n823 B.n822 585
R163 B.n824 B.n46 585
R164 B.n826 B.n825 585
R165 B.n828 B.n45 585
R166 B.n831 B.n830 585
R167 B.n832 B.n44 585
R168 B.n834 B.n833 585
R169 B.n836 B.n43 585
R170 B.n839 B.n838 585
R171 B.n840 B.n42 585
R172 B.n842 B.n841 585
R173 B.n844 B.n41 585
R174 B.n847 B.n846 585
R175 B.n848 B.n40 585
R176 B.n850 B.n849 585
R177 B.n852 B.n39 585
R178 B.n855 B.n854 585
R179 B.n856 B.n38 585
R180 B.n578 B.n36 585
R181 B.n859 B.n36 585
R182 B.n577 B.n35 585
R183 B.n860 B.n35 585
R184 B.n576 B.n34 585
R185 B.n861 B.n34 585
R186 B.n575 B.n574 585
R187 B.n574 B.n30 585
R188 B.n573 B.n29 585
R189 B.n867 B.n29 585
R190 B.n572 B.n28 585
R191 B.n868 B.n28 585
R192 B.n571 B.n27 585
R193 B.n869 B.n27 585
R194 B.n570 B.n569 585
R195 B.n569 B.n23 585
R196 B.n568 B.n22 585
R197 B.n875 B.n22 585
R198 B.n567 B.n21 585
R199 B.n876 B.n21 585
R200 B.n566 B.n20 585
R201 B.n877 B.n20 585
R202 B.n565 B.n564 585
R203 B.n564 B.n19 585
R204 B.n563 B.n15 585
R205 B.n883 B.n15 585
R206 B.n562 B.n14 585
R207 B.n884 B.n14 585
R208 B.n561 B.n13 585
R209 B.n885 B.n13 585
R210 B.n560 B.n559 585
R211 B.n559 B.n12 585
R212 B.n558 B.n557 585
R213 B.n558 B.n8 585
R214 B.n556 B.n7 585
R215 B.n892 B.n7 585
R216 B.n555 B.n6 585
R217 B.n893 B.n6 585
R218 B.n554 B.n5 585
R219 B.n894 B.n5 585
R220 B.n553 B.n552 585
R221 B.n552 B.n4 585
R222 B.n551 B.n113 585
R223 B.n551 B.n550 585
R224 B.n540 B.n114 585
R225 B.n543 B.n114 585
R226 B.n542 B.n541 585
R227 B.n544 B.n542 585
R228 B.n539 B.n119 585
R229 B.n119 B.n118 585
R230 B.n538 B.n537 585
R231 B.n537 B.n536 585
R232 B.n121 B.n120 585
R233 B.n529 B.n121 585
R234 B.n528 B.n527 585
R235 B.n530 B.n528 585
R236 B.n526 B.n126 585
R237 B.n126 B.n125 585
R238 B.n525 B.n524 585
R239 B.n524 B.n523 585
R240 B.n128 B.n127 585
R241 B.n129 B.n128 585
R242 B.n516 B.n515 585
R243 B.n517 B.n516 585
R244 B.n514 B.n133 585
R245 B.n137 B.n133 585
R246 B.n513 B.n512 585
R247 B.n512 B.n511 585
R248 B.n135 B.n134 585
R249 B.n136 B.n135 585
R250 B.n504 B.n503 585
R251 B.n505 B.n504 585
R252 B.n502 B.n142 585
R253 B.n142 B.n141 585
R254 B.n501 B.n500 585
R255 B.n500 B.n499 585
R256 B.n496 B.n146 585
R257 B.n495 B.n494 585
R258 B.n492 B.n147 585
R259 B.n492 B.n145 585
R260 B.n491 B.n490 585
R261 B.n489 B.n488 585
R262 B.n487 B.n149 585
R263 B.n485 B.n484 585
R264 B.n483 B.n150 585
R265 B.n482 B.n481 585
R266 B.n479 B.n151 585
R267 B.n477 B.n476 585
R268 B.n475 B.n152 585
R269 B.n474 B.n473 585
R270 B.n471 B.n153 585
R271 B.n469 B.n468 585
R272 B.n467 B.n154 585
R273 B.n466 B.n465 585
R274 B.n463 B.n155 585
R275 B.n461 B.n460 585
R276 B.n459 B.n156 585
R277 B.n458 B.n457 585
R278 B.n455 B.n157 585
R279 B.n453 B.n452 585
R280 B.n451 B.n158 585
R281 B.n450 B.n449 585
R282 B.n447 B.n159 585
R283 B.n445 B.n444 585
R284 B.n443 B.n160 585
R285 B.n442 B.n441 585
R286 B.n439 B.n161 585
R287 B.n437 B.n436 585
R288 B.n435 B.n162 585
R289 B.n434 B.n433 585
R290 B.n431 B.n163 585
R291 B.n429 B.n428 585
R292 B.n427 B.n164 585
R293 B.n426 B.n425 585
R294 B.n423 B.n165 585
R295 B.n421 B.n420 585
R296 B.n419 B.n166 585
R297 B.n418 B.n417 585
R298 B.n415 B.n167 585
R299 B.n413 B.n412 585
R300 B.n411 B.n168 585
R301 B.n410 B.n409 585
R302 B.n407 B.n169 585
R303 B.n405 B.n404 585
R304 B.n403 B.n170 585
R305 B.n402 B.n401 585
R306 B.n399 B.n171 585
R307 B.n397 B.n396 585
R308 B.n395 B.n172 585
R309 B.n394 B.n393 585
R310 B.n391 B.n173 585
R311 B.n389 B.n388 585
R312 B.n387 B.n174 585
R313 B.n386 B.n385 585
R314 B.n383 B.n175 585
R315 B.n381 B.n380 585
R316 B.n379 B.n176 585
R317 B.n378 B.n377 585
R318 B.n375 B.n177 585
R319 B.n373 B.n372 585
R320 B.n371 B.n178 585
R321 B.n370 B.n369 585
R322 B.n367 B.n366 585
R323 B.n365 B.n364 585
R324 B.n363 B.n183 585
R325 B.n361 B.n360 585
R326 B.n359 B.n184 585
R327 B.n358 B.n357 585
R328 B.n355 B.n185 585
R329 B.n353 B.n352 585
R330 B.n351 B.n186 585
R331 B.n349 B.n348 585
R332 B.n346 B.n189 585
R333 B.n344 B.n343 585
R334 B.n342 B.n190 585
R335 B.n341 B.n340 585
R336 B.n338 B.n191 585
R337 B.n336 B.n335 585
R338 B.n334 B.n192 585
R339 B.n333 B.n332 585
R340 B.n330 B.n193 585
R341 B.n328 B.n327 585
R342 B.n326 B.n194 585
R343 B.n325 B.n324 585
R344 B.n322 B.n195 585
R345 B.n320 B.n319 585
R346 B.n318 B.n196 585
R347 B.n317 B.n316 585
R348 B.n314 B.n197 585
R349 B.n312 B.n311 585
R350 B.n310 B.n198 585
R351 B.n309 B.n308 585
R352 B.n306 B.n199 585
R353 B.n304 B.n303 585
R354 B.n302 B.n200 585
R355 B.n301 B.n300 585
R356 B.n298 B.n201 585
R357 B.n296 B.n295 585
R358 B.n294 B.n202 585
R359 B.n293 B.n292 585
R360 B.n290 B.n203 585
R361 B.n288 B.n287 585
R362 B.n286 B.n204 585
R363 B.n285 B.n284 585
R364 B.n282 B.n205 585
R365 B.n280 B.n279 585
R366 B.n278 B.n206 585
R367 B.n277 B.n276 585
R368 B.n274 B.n207 585
R369 B.n272 B.n271 585
R370 B.n270 B.n208 585
R371 B.n269 B.n268 585
R372 B.n266 B.n209 585
R373 B.n264 B.n263 585
R374 B.n262 B.n210 585
R375 B.n261 B.n260 585
R376 B.n258 B.n211 585
R377 B.n256 B.n255 585
R378 B.n254 B.n212 585
R379 B.n253 B.n252 585
R380 B.n250 B.n213 585
R381 B.n248 B.n247 585
R382 B.n246 B.n214 585
R383 B.n245 B.n244 585
R384 B.n242 B.n215 585
R385 B.n240 B.n239 585
R386 B.n238 B.n216 585
R387 B.n237 B.n236 585
R388 B.n234 B.n217 585
R389 B.n232 B.n231 585
R390 B.n230 B.n218 585
R391 B.n229 B.n228 585
R392 B.n226 B.n219 585
R393 B.n224 B.n223 585
R394 B.n222 B.n221 585
R395 B.n144 B.n143 585
R396 B.n498 B.n497 585
R397 B.n499 B.n498 585
R398 B.n140 B.n139 585
R399 B.n141 B.n140 585
R400 B.n507 B.n506 585
R401 B.n506 B.n505 585
R402 B.n508 B.n138 585
R403 B.n138 B.n136 585
R404 B.n510 B.n509 585
R405 B.n511 B.n510 585
R406 B.n132 B.n131 585
R407 B.n137 B.n132 585
R408 B.n519 B.n518 585
R409 B.n518 B.n517 585
R410 B.n520 B.n130 585
R411 B.n130 B.n129 585
R412 B.n522 B.n521 585
R413 B.n523 B.n522 585
R414 B.n124 B.n123 585
R415 B.n125 B.n124 585
R416 B.n532 B.n531 585
R417 B.n531 B.n530 585
R418 B.n533 B.n122 585
R419 B.n529 B.n122 585
R420 B.n535 B.n534 585
R421 B.n536 B.n535 585
R422 B.n117 B.n116 585
R423 B.n118 B.n117 585
R424 B.n546 B.n545 585
R425 B.n545 B.n544 585
R426 B.n547 B.n115 585
R427 B.n543 B.n115 585
R428 B.n549 B.n548 585
R429 B.n550 B.n549 585
R430 B.n3 B.n0 585
R431 B.n4 B.n3 585
R432 B.n891 B.n1 585
R433 B.n892 B.n891 585
R434 B.n890 B.n889 585
R435 B.n890 B.n8 585
R436 B.n888 B.n9 585
R437 B.n12 B.n9 585
R438 B.n887 B.n886 585
R439 B.n886 B.n885 585
R440 B.n11 B.n10 585
R441 B.n884 B.n11 585
R442 B.n882 B.n881 585
R443 B.n883 B.n882 585
R444 B.n880 B.n16 585
R445 B.n19 B.n16 585
R446 B.n879 B.n878 585
R447 B.n878 B.n877 585
R448 B.n18 B.n17 585
R449 B.n876 B.n18 585
R450 B.n874 B.n873 585
R451 B.n875 B.n874 585
R452 B.n872 B.n24 585
R453 B.n24 B.n23 585
R454 B.n871 B.n870 585
R455 B.n870 B.n869 585
R456 B.n26 B.n25 585
R457 B.n868 B.n26 585
R458 B.n866 B.n865 585
R459 B.n867 B.n866 585
R460 B.n864 B.n31 585
R461 B.n31 B.n30 585
R462 B.n863 B.n862 585
R463 B.n862 B.n861 585
R464 B.n33 B.n32 585
R465 B.n860 B.n33 585
R466 B.n858 B.n857 585
R467 B.n859 B.n858 585
R468 B.n895 B.n894 585
R469 B.n893 B.n2 585
R470 B.n858 B.n38 516.524
R471 B.n112 B.n36 516.524
R472 B.n500 B.n144 516.524
R473 B.n498 B.n146 516.524
R474 B.n582 B.n37 256.663
R475 B.n584 B.n37 256.663
R476 B.n590 B.n37 256.663
R477 B.n592 B.n37 256.663
R478 B.n598 B.n37 256.663
R479 B.n600 B.n37 256.663
R480 B.n606 B.n37 256.663
R481 B.n608 B.n37 256.663
R482 B.n614 B.n37 256.663
R483 B.n616 B.n37 256.663
R484 B.n622 B.n37 256.663
R485 B.n624 B.n37 256.663
R486 B.n630 B.n37 256.663
R487 B.n632 B.n37 256.663
R488 B.n638 B.n37 256.663
R489 B.n640 B.n37 256.663
R490 B.n646 B.n37 256.663
R491 B.n648 B.n37 256.663
R492 B.n654 B.n37 256.663
R493 B.n656 B.n37 256.663
R494 B.n662 B.n37 256.663
R495 B.n664 B.n37 256.663
R496 B.n670 B.n37 256.663
R497 B.n672 B.n37 256.663
R498 B.n678 B.n37 256.663
R499 B.n680 B.n37 256.663
R500 B.n686 B.n37 256.663
R501 B.n688 B.n37 256.663
R502 B.n694 B.n37 256.663
R503 B.n696 B.n37 256.663
R504 B.n702 B.n37 256.663
R505 B.n80 B.n37 256.663
R506 B.n708 B.n37 256.663
R507 B.n714 B.n37 256.663
R508 B.n716 B.n37 256.663
R509 B.n722 B.n37 256.663
R510 B.n724 B.n37 256.663
R511 B.n731 B.n37 256.663
R512 B.n733 B.n37 256.663
R513 B.n739 B.n37 256.663
R514 B.n741 B.n37 256.663
R515 B.n747 B.n37 256.663
R516 B.n749 B.n37 256.663
R517 B.n755 B.n37 256.663
R518 B.n757 B.n37 256.663
R519 B.n763 B.n37 256.663
R520 B.n765 B.n37 256.663
R521 B.n771 B.n37 256.663
R522 B.n773 B.n37 256.663
R523 B.n779 B.n37 256.663
R524 B.n781 B.n37 256.663
R525 B.n787 B.n37 256.663
R526 B.n789 B.n37 256.663
R527 B.n795 B.n37 256.663
R528 B.n797 B.n37 256.663
R529 B.n803 B.n37 256.663
R530 B.n805 B.n37 256.663
R531 B.n811 B.n37 256.663
R532 B.n813 B.n37 256.663
R533 B.n819 B.n37 256.663
R534 B.n821 B.n37 256.663
R535 B.n827 B.n37 256.663
R536 B.n829 B.n37 256.663
R537 B.n835 B.n37 256.663
R538 B.n837 B.n37 256.663
R539 B.n843 B.n37 256.663
R540 B.n845 B.n37 256.663
R541 B.n851 B.n37 256.663
R542 B.n853 B.n37 256.663
R543 B.n493 B.n145 256.663
R544 B.n148 B.n145 256.663
R545 B.n486 B.n145 256.663
R546 B.n480 B.n145 256.663
R547 B.n478 B.n145 256.663
R548 B.n472 B.n145 256.663
R549 B.n470 B.n145 256.663
R550 B.n464 B.n145 256.663
R551 B.n462 B.n145 256.663
R552 B.n456 B.n145 256.663
R553 B.n454 B.n145 256.663
R554 B.n448 B.n145 256.663
R555 B.n446 B.n145 256.663
R556 B.n440 B.n145 256.663
R557 B.n438 B.n145 256.663
R558 B.n432 B.n145 256.663
R559 B.n430 B.n145 256.663
R560 B.n424 B.n145 256.663
R561 B.n422 B.n145 256.663
R562 B.n416 B.n145 256.663
R563 B.n414 B.n145 256.663
R564 B.n408 B.n145 256.663
R565 B.n406 B.n145 256.663
R566 B.n400 B.n145 256.663
R567 B.n398 B.n145 256.663
R568 B.n392 B.n145 256.663
R569 B.n390 B.n145 256.663
R570 B.n384 B.n145 256.663
R571 B.n382 B.n145 256.663
R572 B.n376 B.n145 256.663
R573 B.n374 B.n145 256.663
R574 B.n368 B.n145 256.663
R575 B.n182 B.n145 256.663
R576 B.n362 B.n145 256.663
R577 B.n356 B.n145 256.663
R578 B.n354 B.n145 256.663
R579 B.n347 B.n145 256.663
R580 B.n345 B.n145 256.663
R581 B.n339 B.n145 256.663
R582 B.n337 B.n145 256.663
R583 B.n331 B.n145 256.663
R584 B.n329 B.n145 256.663
R585 B.n323 B.n145 256.663
R586 B.n321 B.n145 256.663
R587 B.n315 B.n145 256.663
R588 B.n313 B.n145 256.663
R589 B.n307 B.n145 256.663
R590 B.n305 B.n145 256.663
R591 B.n299 B.n145 256.663
R592 B.n297 B.n145 256.663
R593 B.n291 B.n145 256.663
R594 B.n289 B.n145 256.663
R595 B.n283 B.n145 256.663
R596 B.n281 B.n145 256.663
R597 B.n275 B.n145 256.663
R598 B.n273 B.n145 256.663
R599 B.n267 B.n145 256.663
R600 B.n265 B.n145 256.663
R601 B.n259 B.n145 256.663
R602 B.n257 B.n145 256.663
R603 B.n251 B.n145 256.663
R604 B.n249 B.n145 256.663
R605 B.n243 B.n145 256.663
R606 B.n241 B.n145 256.663
R607 B.n235 B.n145 256.663
R608 B.n233 B.n145 256.663
R609 B.n227 B.n145 256.663
R610 B.n225 B.n145 256.663
R611 B.n220 B.n145 256.663
R612 B.n897 B.n896 256.663
R613 B.n854 B.n852 163.367
R614 B.n850 B.n40 163.367
R615 B.n846 B.n844 163.367
R616 B.n842 B.n42 163.367
R617 B.n838 B.n836 163.367
R618 B.n834 B.n44 163.367
R619 B.n830 B.n828 163.367
R620 B.n826 B.n46 163.367
R621 B.n822 B.n820 163.367
R622 B.n818 B.n48 163.367
R623 B.n814 B.n812 163.367
R624 B.n810 B.n50 163.367
R625 B.n806 B.n804 163.367
R626 B.n802 B.n52 163.367
R627 B.n798 B.n796 163.367
R628 B.n794 B.n54 163.367
R629 B.n790 B.n788 163.367
R630 B.n786 B.n56 163.367
R631 B.n782 B.n780 163.367
R632 B.n778 B.n58 163.367
R633 B.n774 B.n772 163.367
R634 B.n770 B.n60 163.367
R635 B.n766 B.n764 163.367
R636 B.n762 B.n62 163.367
R637 B.n758 B.n756 163.367
R638 B.n754 B.n64 163.367
R639 B.n750 B.n748 163.367
R640 B.n746 B.n66 163.367
R641 B.n742 B.n740 163.367
R642 B.n738 B.n68 163.367
R643 B.n734 B.n732 163.367
R644 B.n730 B.n70 163.367
R645 B.n725 B.n723 163.367
R646 B.n721 B.n74 163.367
R647 B.n717 B.n715 163.367
R648 B.n713 B.n76 163.367
R649 B.n709 B.n707 163.367
R650 B.n704 B.n703 163.367
R651 B.n701 B.n82 163.367
R652 B.n697 B.n695 163.367
R653 B.n693 B.n84 163.367
R654 B.n689 B.n687 163.367
R655 B.n685 B.n86 163.367
R656 B.n681 B.n679 163.367
R657 B.n677 B.n88 163.367
R658 B.n673 B.n671 163.367
R659 B.n669 B.n90 163.367
R660 B.n665 B.n663 163.367
R661 B.n661 B.n92 163.367
R662 B.n657 B.n655 163.367
R663 B.n653 B.n94 163.367
R664 B.n649 B.n647 163.367
R665 B.n645 B.n96 163.367
R666 B.n641 B.n639 163.367
R667 B.n637 B.n98 163.367
R668 B.n633 B.n631 163.367
R669 B.n629 B.n100 163.367
R670 B.n625 B.n623 163.367
R671 B.n621 B.n102 163.367
R672 B.n617 B.n615 163.367
R673 B.n613 B.n104 163.367
R674 B.n609 B.n607 163.367
R675 B.n605 B.n106 163.367
R676 B.n601 B.n599 163.367
R677 B.n597 B.n108 163.367
R678 B.n593 B.n591 163.367
R679 B.n589 B.n110 163.367
R680 B.n585 B.n583 163.367
R681 B.n581 B.n112 163.367
R682 B.n500 B.n142 163.367
R683 B.n504 B.n142 163.367
R684 B.n504 B.n135 163.367
R685 B.n512 B.n135 163.367
R686 B.n512 B.n133 163.367
R687 B.n516 B.n133 163.367
R688 B.n516 B.n128 163.367
R689 B.n524 B.n128 163.367
R690 B.n524 B.n126 163.367
R691 B.n528 B.n126 163.367
R692 B.n528 B.n121 163.367
R693 B.n537 B.n121 163.367
R694 B.n537 B.n119 163.367
R695 B.n542 B.n119 163.367
R696 B.n542 B.n114 163.367
R697 B.n551 B.n114 163.367
R698 B.n552 B.n551 163.367
R699 B.n552 B.n5 163.367
R700 B.n6 B.n5 163.367
R701 B.n7 B.n6 163.367
R702 B.n558 B.n7 163.367
R703 B.n559 B.n558 163.367
R704 B.n559 B.n13 163.367
R705 B.n14 B.n13 163.367
R706 B.n15 B.n14 163.367
R707 B.n564 B.n15 163.367
R708 B.n564 B.n20 163.367
R709 B.n21 B.n20 163.367
R710 B.n22 B.n21 163.367
R711 B.n569 B.n22 163.367
R712 B.n569 B.n27 163.367
R713 B.n28 B.n27 163.367
R714 B.n29 B.n28 163.367
R715 B.n574 B.n29 163.367
R716 B.n574 B.n34 163.367
R717 B.n35 B.n34 163.367
R718 B.n36 B.n35 163.367
R719 B.n494 B.n492 163.367
R720 B.n492 B.n491 163.367
R721 B.n488 B.n487 163.367
R722 B.n485 B.n150 163.367
R723 B.n481 B.n479 163.367
R724 B.n477 B.n152 163.367
R725 B.n473 B.n471 163.367
R726 B.n469 B.n154 163.367
R727 B.n465 B.n463 163.367
R728 B.n461 B.n156 163.367
R729 B.n457 B.n455 163.367
R730 B.n453 B.n158 163.367
R731 B.n449 B.n447 163.367
R732 B.n445 B.n160 163.367
R733 B.n441 B.n439 163.367
R734 B.n437 B.n162 163.367
R735 B.n433 B.n431 163.367
R736 B.n429 B.n164 163.367
R737 B.n425 B.n423 163.367
R738 B.n421 B.n166 163.367
R739 B.n417 B.n415 163.367
R740 B.n413 B.n168 163.367
R741 B.n409 B.n407 163.367
R742 B.n405 B.n170 163.367
R743 B.n401 B.n399 163.367
R744 B.n397 B.n172 163.367
R745 B.n393 B.n391 163.367
R746 B.n389 B.n174 163.367
R747 B.n385 B.n383 163.367
R748 B.n381 B.n176 163.367
R749 B.n377 B.n375 163.367
R750 B.n373 B.n178 163.367
R751 B.n369 B.n367 163.367
R752 B.n364 B.n363 163.367
R753 B.n361 B.n184 163.367
R754 B.n357 B.n355 163.367
R755 B.n353 B.n186 163.367
R756 B.n348 B.n346 163.367
R757 B.n344 B.n190 163.367
R758 B.n340 B.n338 163.367
R759 B.n336 B.n192 163.367
R760 B.n332 B.n330 163.367
R761 B.n328 B.n194 163.367
R762 B.n324 B.n322 163.367
R763 B.n320 B.n196 163.367
R764 B.n316 B.n314 163.367
R765 B.n312 B.n198 163.367
R766 B.n308 B.n306 163.367
R767 B.n304 B.n200 163.367
R768 B.n300 B.n298 163.367
R769 B.n296 B.n202 163.367
R770 B.n292 B.n290 163.367
R771 B.n288 B.n204 163.367
R772 B.n284 B.n282 163.367
R773 B.n280 B.n206 163.367
R774 B.n276 B.n274 163.367
R775 B.n272 B.n208 163.367
R776 B.n268 B.n266 163.367
R777 B.n264 B.n210 163.367
R778 B.n260 B.n258 163.367
R779 B.n256 B.n212 163.367
R780 B.n252 B.n250 163.367
R781 B.n248 B.n214 163.367
R782 B.n244 B.n242 163.367
R783 B.n240 B.n216 163.367
R784 B.n236 B.n234 163.367
R785 B.n232 B.n218 163.367
R786 B.n228 B.n226 163.367
R787 B.n224 B.n221 163.367
R788 B.n498 B.n140 163.367
R789 B.n506 B.n140 163.367
R790 B.n506 B.n138 163.367
R791 B.n510 B.n138 163.367
R792 B.n510 B.n132 163.367
R793 B.n518 B.n132 163.367
R794 B.n518 B.n130 163.367
R795 B.n522 B.n130 163.367
R796 B.n522 B.n124 163.367
R797 B.n531 B.n124 163.367
R798 B.n531 B.n122 163.367
R799 B.n535 B.n122 163.367
R800 B.n535 B.n117 163.367
R801 B.n545 B.n117 163.367
R802 B.n545 B.n115 163.367
R803 B.n549 B.n115 163.367
R804 B.n549 B.n3 163.367
R805 B.n895 B.n3 163.367
R806 B.n891 B.n2 163.367
R807 B.n891 B.n890 163.367
R808 B.n890 B.n9 163.367
R809 B.n886 B.n9 163.367
R810 B.n886 B.n11 163.367
R811 B.n882 B.n11 163.367
R812 B.n882 B.n16 163.367
R813 B.n878 B.n16 163.367
R814 B.n878 B.n18 163.367
R815 B.n874 B.n18 163.367
R816 B.n874 B.n24 163.367
R817 B.n870 B.n24 163.367
R818 B.n870 B.n26 163.367
R819 B.n866 B.n26 163.367
R820 B.n866 B.n31 163.367
R821 B.n862 B.n31 163.367
R822 B.n862 B.n33 163.367
R823 B.n858 B.n33 163.367
R824 B.n77 B.t10 93.908
R825 B.n187 B.t7 93.908
R826 B.n71 B.t13 93.8813
R827 B.n179 B.t17 93.8813
R828 B.n853 B.n38 71.676
R829 B.n852 B.n851 71.676
R830 B.n845 B.n40 71.676
R831 B.n844 B.n843 71.676
R832 B.n837 B.n42 71.676
R833 B.n836 B.n835 71.676
R834 B.n829 B.n44 71.676
R835 B.n828 B.n827 71.676
R836 B.n821 B.n46 71.676
R837 B.n820 B.n819 71.676
R838 B.n813 B.n48 71.676
R839 B.n812 B.n811 71.676
R840 B.n805 B.n50 71.676
R841 B.n804 B.n803 71.676
R842 B.n797 B.n52 71.676
R843 B.n796 B.n795 71.676
R844 B.n789 B.n54 71.676
R845 B.n788 B.n787 71.676
R846 B.n781 B.n56 71.676
R847 B.n780 B.n779 71.676
R848 B.n773 B.n58 71.676
R849 B.n772 B.n771 71.676
R850 B.n765 B.n60 71.676
R851 B.n764 B.n763 71.676
R852 B.n757 B.n62 71.676
R853 B.n756 B.n755 71.676
R854 B.n749 B.n64 71.676
R855 B.n748 B.n747 71.676
R856 B.n741 B.n66 71.676
R857 B.n740 B.n739 71.676
R858 B.n733 B.n68 71.676
R859 B.n732 B.n731 71.676
R860 B.n724 B.n70 71.676
R861 B.n723 B.n722 71.676
R862 B.n716 B.n74 71.676
R863 B.n715 B.n714 71.676
R864 B.n708 B.n76 71.676
R865 B.n707 B.n80 71.676
R866 B.n703 B.n702 71.676
R867 B.n696 B.n82 71.676
R868 B.n695 B.n694 71.676
R869 B.n688 B.n84 71.676
R870 B.n687 B.n686 71.676
R871 B.n680 B.n86 71.676
R872 B.n679 B.n678 71.676
R873 B.n672 B.n88 71.676
R874 B.n671 B.n670 71.676
R875 B.n664 B.n90 71.676
R876 B.n663 B.n662 71.676
R877 B.n656 B.n92 71.676
R878 B.n655 B.n654 71.676
R879 B.n648 B.n94 71.676
R880 B.n647 B.n646 71.676
R881 B.n640 B.n96 71.676
R882 B.n639 B.n638 71.676
R883 B.n632 B.n98 71.676
R884 B.n631 B.n630 71.676
R885 B.n624 B.n100 71.676
R886 B.n623 B.n622 71.676
R887 B.n616 B.n102 71.676
R888 B.n615 B.n614 71.676
R889 B.n608 B.n104 71.676
R890 B.n607 B.n606 71.676
R891 B.n600 B.n106 71.676
R892 B.n599 B.n598 71.676
R893 B.n592 B.n108 71.676
R894 B.n591 B.n590 71.676
R895 B.n584 B.n110 71.676
R896 B.n583 B.n582 71.676
R897 B.n582 B.n581 71.676
R898 B.n585 B.n584 71.676
R899 B.n590 B.n589 71.676
R900 B.n593 B.n592 71.676
R901 B.n598 B.n597 71.676
R902 B.n601 B.n600 71.676
R903 B.n606 B.n605 71.676
R904 B.n609 B.n608 71.676
R905 B.n614 B.n613 71.676
R906 B.n617 B.n616 71.676
R907 B.n622 B.n621 71.676
R908 B.n625 B.n624 71.676
R909 B.n630 B.n629 71.676
R910 B.n633 B.n632 71.676
R911 B.n638 B.n637 71.676
R912 B.n641 B.n640 71.676
R913 B.n646 B.n645 71.676
R914 B.n649 B.n648 71.676
R915 B.n654 B.n653 71.676
R916 B.n657 B.n656 71.676
R917 B.n662 B.n661 71.676
R918 B.n665 B.n664 71.676
R919 B.n670 B.n669 71.676
R920 B.n673 B.n672 71.676
R921 B.n678 B.n677 71.676
R922 B.n681 B.n680 71.676
R923 B.n686 B.n685 71.676
R924 B.n689 B.n688 71.676
R925 B.n694 B.n693 71.676
R926 B.n697 B.n696 71.676
R927 B.n702 B.n701 71.676
R928 B.n704 B.n80 71.676
R929 B.n709 B.n708 71.676
R930 B.n714 B.n713 71.676
R931 B.n717 B.n716 71.676
R932 B.n722 B.n721 71.676
R933 B.n725 B.n724 71.676
R934 B.n731 B.n730 71.676
R935 B.n734 B.n733 71.676
R936 B.n739 B.n738 71.676
R937 B.n742 B.n741 71.676
R938 B.n747 B.n746 71.676
R939 B.n750 B.n749 71.676
R940 B.n755 B.n754 71.676
R941 B.n758 B.n757 71.676
R942 B.n763 B.n762 71.676
R943 B.n766 B.n765 71.676
R944 B.n771 B.n770 71.676
R945 B.n774 B.n773 71.676
R946 B.n779 B.n778 71.676
R947 B.n782 B.n781 71.676
R948 B.n787 B.n786 71.676
R949 B.n790 B.n789 71.676
R950 B.n795 B.n794 71.676
R951 B.n798 B.n797 71.676
R952 B.n803 B.n802 71.676
R953 B.n806 B.n805 71.676
R954 B.n811 B.n810 71.676
R955 B.n814 B.n813 71.676
R956 B.n819 B.n818 71.676
R957 B.n822 B.n821 71.676
R958 B.n827 B.n826 71.676
R959 B.n830 B.n829 71.676
R960 B.n835 B.n834 71.676
R961 B.n838 B.n837 71.676
R962 B.n843 B.n842 71.676
R963 B.n846 B.n845 71.676
R964 B.n851 B.n850 71.676
R965 B.n854 B.n853 71.676
R966 B.n493 B.n146 71.676
R967 B.n491 B.n148 71.676
R968 B.n487 B.n486 71.676
R969 B.n480 B.n150 71.676
R970 B.n479 B.n478 71.676
R971 B.n472 B.n152 71.676
R972 B.n471 B.n470 71.676
R973 B.n464 B.n154 71.676
R974 B.n463 B.n462 71.676
R975 B.n456 B.n156 71.676
R976 B.n455 B.n454 71.676
R977 B.n448 B.n158 71.676
R978 B.n447 B.n446 71.676
R979 B.n440 B.n160 71.676
R980 B.n439 B.n438 71.676
R981 B.n432 B.n162 71.676
R982 B.n431 B.n430 71.676
R983 B.n424 B.n164 71.676
R984 B.n423 B.n422 71.676
R985 B.n416 B.n166 71.676
R986 B.n415 B.n414 71.676
R987 B.n408 B.n168 71.676
R988 B.n407 B.n406 71.676
R989 B.n400 B.n170 71.676
R990 B.n399 B.n398 71.676
R991 B.n392 B.n172 71.676
R992 B.n391 B.n390 71.676
R993 B.n384 B.n174 71.676
R994 B.n383 B.n382 71.676
R995 B.n376 B.n176 71.676
R996 B.n375 B.n374 71.676
R997 B.n368 B.n178 71.676
R998 B.n367 B.n182 71.676
R999 B.n363 B.n362 71.676
R1000 B.n356 B.n184 71.676
R1001 B.n355 B.n354 71.676
R1002 B.n347 B.n186 71.676
R1003 B.n346 B.n345 71.676
R1004 B.n339 B.n190 71.676
R1005 B.n338 B.n337 71.676
R1006 B.n331 B.n192 71.676
R1007 B.n330 B.n329 71.676
R1008 B.n323 B.n194 71.676
R1009 B.n322 B.n321 71.676
R1010 B.n315 B.n196 71.676
R1011 B.n314 B.n313 71.676
R1012 B.n307 B.n198 71.676
R1013 B.n306 B.n305 71.676
R1014 B.n299 B.n200 71.676
R1015 B.n298 B.n297 71.676
R1016 B.n291 B.n202 71.676
R1017 B.n290 B.n289 71.676
R1018 B.n283 B.n204 71.676
R1019 B.n282 B.n281 71.676
R1020 B.n275 B.n206 71.676
R1021 B.n274 B.n273 71.676
R1022 B.n267 B.n208 71.676
R1023 B.n266 B.n265 71.676
R1024 B.n259 B.n210 71.676
R1025 B.n258 B.n257 71.676
R1026 B.n251 B.n212 71.676
R1027 B.n250 B.n249 71.676
R1028 B.n243 B.n214 71.676
R1029 B.n242 B.n241 71.676
R1030 B.n235 B.n216 71.676
R1031 B.n234 B.n233 71.676
R1032 B.n227 B.n218 71.676
R1033 B.n226 B.n225 71.676
R1034 B.n221 B.n220 71.676
R1035 B.n494 B.n493 71.676
R1036 B.n488 B.n148 71.676
R1037 B.n486 B.n485 71.676
R1038 B.n481 B.n480 71.676
R1039 B.n478 B.n477 71.676
R1040 B.n473 B.n472 71.676
R1041 B.n470 B.n469 71.676
R1042 B.n465 B.n464 71.676
R1043 B.n462 B.n461 71.676
R1044 B.n457 B.n456 71.676
R1045 B.n454 B.n453 71.676
R1046 B.n449 B.n448 71.676
R1047 B.n446 B.n445 71.676
R1048 B.n441 B.n440 71.676
R1049 B.n438 B.n437 71.676
R1050 B.n433 B.n432 71.676
R1051 B.n430 B.n429 71.676
R1052 B.n425 B.n424 71.676
R1053 B.n422 B.n421 71.676
R1054 B.n417 B.n416 71.676
R1055 B.n414 B.n413 71.676
R1056 B.n409 B.n408 71.676
R1057 B.n406 B.n405 71.676
R1058 B.n401 B.n400 71.676
R1059 B.n398 B.n397 71.676
R1060 B.n393 B.n392 71.676
R1061 B.n390 B.n389 71.676
R1062 B.n385 B.n384 71.676
R1063 B.n382 B.n381 71.676
R1064 B.n377 B.n376 71.676
R1065 B.n374 B.n373 71.676
R1066 B.n369 B.n368 71.676
R1067 B.n364 B.n182 71.676
R1068 B.n362 B.n361 71.676
R1069 B.n357 B.n356 71.676
R1070 B.n354 B.n353 71.676
R1071 B.n348 B.n347 71.676
R1072 B.n345 B.n344 71.676
R1073 B.n340 B.n339 71.676
R1074 B.n337 B.n336 71.676
R1075 B.n332 B.n331 71.676
R1076 B.n329 B.n328 71.676
R1077 B.n324 B.n323 71.676
R1078 B.n321 B.n320 71.676
R1079 B.n316 B.n315 71.676
R1080 B.n313 B.n312 71.676
R1081 B.n308 B.n307 71.676
R1082 B.n305 B.n304 71.676
R1083 B.n300 B.n299 71.676
R1084 B.n297 B.n296 71.676
R1085 B.n292 B.n291 71.676
R1086 B.n289 B.n288 71.676
R1087 B.n284 B.n283 71.676
R1088 B.n281 B.n280 71.676
R1089 B.n276 B.n275 71.676
R1090 B.n273 B.n272 71.676
R1091 B.n268 B.n267 71.676
R1092 B.n265 B.n264 71.676
R1093 B.n260 B.n259 71.676
R1094 B.n257 B.n256 71.676
R1095 B.n252 B.n251 71.676
R1096 B.n249 B.n248 71.676
R1097 B.n244 B.n243 71.676
R1098 B.n241 B.n240 71.676
R1099 B.n236 B.n235 71.676
R1100 B.n233 B.n232 71.676
R1101 B.n228 B.n227 71.676
R1102 B.n225 B.n224 71.676
R1103 B.n220 B.n144 71.676
R1104 B.n896 B.n895 71.676
R1105 B.n896 B.n2 71.676
R1106 B.n78 B.t11 71.411
R1107 B.n188 B.t6 71.411
R1108 B.n72 B.t14 71.3843
R1109 B.n180 B.t16 71.3843
R1110 B.n727 B.n72 59.5399
R1111 B.n79 B.n78 59.5399
R1112 B.n350 B.n188 59.5399
R1113 B.n181 B.n180 59.5399
R1114 B.n499 B.n145 49.2966
R1115 B.n859 B.n37 49.2966
R1116 B.n497 B.n496 33.5615
R1117 B.n501 B.n143 33.5615
R1118 B.n579 B.n578 33.5615
R1119 B.n857 B.n856 33.5615
R1120 B.n499 B.n141 29.6654
R1121 B.n505 B.n141 29.6654
R1122 B.n505 B.n136 29.6654
R1123 B.n511 B.n136 29.6654
R1124 B.n511 B.n137 29.6654
R1125 B.n517 B.n129 29.6654
R1126 B.n523 B.n129 29.6654
R1127 B.n523 B.n125 29.6654
R1128 B.n530 B.n125 29.6654
R1129 B.n530 B.n529 29.6654
R1130 B.n536 B.n118 29.6654
R1131 B.n544 B.n118 29.6654
R1132 B.n544 B.n543 29.6654
R1133 B.n550 B.n4 29.6654
R1134 B.n894 B.n4 29.6654
R1135 B.n894 B.n893 29.6654
R1136 B.n893 B.n892 29.6654
R1137 B.n892 B.n8 29.6654
R1138 B.n885 B.n12 29.6654
R1139 B.n885 B.n884 29.6654
R1140 B.n884 B.n883 29.6654
R1141 B.n877 B.n19 29.6654
R1142 B.n877 B.n876 29.6654
R1143 B.n876 B.n875 29.6654
R1144 B.n875 B.n23 29.6654
R1145 B.n869 B.n23 29.6654
R1146 B.n868 B.n867 29.6654
R1147 B.n867 B.n30 29.6654
R1148 B.n861 B.n30 29.6654
R1149 B.n861 B.n860 29.6654
R1150 B.n860 B.n859 29.6654
R1151 B.n517 B.t5 24.8666
R1152 B.n869 B.t9 24.8666
R1153 B.n550 B.t3 23.9942
R1154 B.t1 B.n8 23.9942
R1155 B.n529 B.t0 23.1217
R1156 B.n19 B.t2 23.1217
R1157 B.n72 B.n71 22.4975
R1158 B.n78 B.n77 22.4975
R1159 B.n188 B.n187 22.4975
R1160 B.n180 B.n179 22.4975
R1161 B B.n897 18.0485
R1162 B.n497 B.n139 10.6151
R1163 B.n507 B.n139 10.6151
R1164 B.n508 B.n507 10.6151
R1165 B.n509 B.n508 10.6151
R1166 B.n509 B.n131 10.6151
R1167 B.n519 B.n131 10.6151
R1168 B.n520 B.n519 10.6151
R1169 B.n521 B.n520 10.6151
R1170 B.n521 B.n123 10.6151
R1171 B.n532 B.n123 10.6151
R1172 B.n533 B.n532 10.6151
R1173 B.n534 B.n533 10.6151
R1174 B.n534 B.n116 10.6151
R1175 B.n546 B.n116 10.6151
R1176 B.n547 B.n546 10.6151
R1177 B.n548 B.n547 10.6151
R1178 B.n548 B.n0 10.6151
R1179 B.n496 B.n495 10.6151
R1180 B.n495 B.n147 10.6151
R1181 B.n490 B.n147 10.6151
R1182 B.n490 B.n489 10.6151
R1183 B.n489 B.n149 10.6151
R1184 B.n484 B.n149 10.6151
R1185 B.n484 B.n483 10.6151
R1186 B.n483 B.n482 10.6151
R1187 B.n482 B.n151 10.6151
R1188 B.n476 B.n151 10.6151
R1189 B.n476 B.n475 10.6151
R1190 B.n475 B.n474 10.6151
R1191 B.n474 B.n153 10.6151
R1192 B.n468 B.n153 10.6151
R1193 B.n468 B.n467 10.6151
R1194 B.n467 B.n466 10.6151
R1195 B.n466 B.n155 10.6151
R1196 B.n460 B.n155 10.6151
R1197 B.n460 B.n459 10.6151
R1198 B.n459 B.n458 10.6151
R1199 B.n458 B.n157 10.6151
R1200 B.n452 B.n157 10.6151
R1201 B.n452 B.n451 10.6151
R1202 B.n451 B.n450 10.6151
R1203 B.n450 B.n159 10.6151
R1204 B.n444 B.n159 10.6151
R1205 B.n444 B.n443 10.6151
R1206 B.n443 B.n442 10.6151
R1207 B.n442 B.n161 10.6151
R1208 B.n436 B.n161 10.6151
R1209 B.n436 B.n435 10.6151
R1210 B.n435 B.n434 10.6151
R1211 B.n434 B.n163 10.6151
R1212 B.n428 B.n163 10.6151
R1213 B.n428 B.n427 10.6151
R1214 B.n427 B.n426 10.6151
R1215 B.n426 B.n165 10.6151
R1216 B.n420 B.n165 10.6151
R1217 B.n420 B.n419 10.6151
R1218 B.n419 B.n418 10.6151
R1219 B.n418 B.n167 10.6151
R1220 B.n412 B.n167 10.6151
R1221 B.n412 B.n411 10.6151
R1222 B.n411 B.n410 10.6151
R1223 B.n410 B.n169 10.6151
R1224 B.n404 B.n169 10.6151
R1225 B.n404 B.n403 10.6151
R1226 B.n403 B.n402 10.6151
R1227 B.n402 B.n171 10.6151
R1228 B.n396 B.n171 10.6151
R1229 B.n396 B.n395 10.6151
R1230 B.n395 B.n394 10.6151
R1231 B.n394 B.n173 10.6151
R1232 B.n388 B.n173 10.6151
R1233 B.n388 B.n387 10.6151
R1234 B.n387 B.n386 10.6151
R1235 B.n386 B.n175 10.6151
R1236 B.n380 B.n175 10.6151
R1237 B.n380 B.n379 10.6151
R1238 B.n379 B.n378 10.6151
R1239 B.n378 B.n177 10.6151
R1240 B.n372 B.n177 10.6151
R1241 B.n372 B.n371 10.6151
R1242 B.n371 B.n370 10.6151
R1243 B.n366 B.n365 10.6151
R1244 B.n365 B.n183 10.6151
R1245 B.n360 B.n183 10.6151
R1246 B.n360 B.n359 10.6151
R1247 B.n359 B.n358 10.6151
R1248 B.n358 B.n185 10.6151
R1249 B.n352 B.n185 10.6151
R1250 B.n352 B.n351 10.6151
R1251 B.n349 B.n189 10.6151
R1252 B.n343 B.n189 10.6151
R1253 B.n343 B.n342 10.6151
R1254 B.n342 B.n341 10.6151
R1255 B.n341 B.n191 10.6151
R1256 B.n335 B.n191 10.6151
R1257 B.n335 B.n334 10.6151
R1258 B.n334 B.n333 10.6151
R1259 B.n333 B.n193 10.6151
R1260 B.n327 B.n193 10.6151
R1261 B.n327 B.n326 10.6151
R1262 B.n326 B.n325 10.6151
R1263 B.n325 B.n195 10.6151
R1264 B.n319 B.n195 10.6151
R1265 B.n319 B.n318 10.6151
R1266 B.n318 B.n317 10.6151
R1267 B.n317 B.n197 10.6151
R1268 B.n311 B.n197 10.6151
R1269 B.n311 B.n310 10.6151
R1270 B.n310 B.n309 10.6151
R1271 B.n309 B.n199 10.6151
R1272 B.n303 B.n199 10.6151
R1273 B.n303 B.n302 10.6151
R1274 B.n302 B.n301 10.6151
R1275 B.n301 B.n201 10.6151
R1276 B.n295 B.n201 10.6151
R1277 B.n295 B.n294 10.6151
R1278 B.n294 B.n293 10.6151
R1279 B.n293 B.n203 10.6151
R1280 B.n287 B.n203 10.6151
R1281 B.n287 B.n286 10.6151
R1282 B.n286 B.n285 10.6151
R1283 B.n285 B.n205 10.6151
R1284 B.n279 B.n205 10.6151
R1285 B.n279 B.n278 10.6151
R1286 B.n278 B.n277 10.6151
R1287 B.n277 B.n207 10.6151
R1288 B.n271 B.n207 10.6151
R1289 B.n271 B.n270 10.6151
R1290 B.n270 B.n269 10.6151
R1291 B.n269 B.n209 10.6151
R1292 B.n263 B.n209 10.6151
R1293 B.n263 B.n262 10.6151
R1294 B.n262 B.n261 10.6151
R1295 B.n261 B.n211 10.6151
R1296 B.n255 B.n211 10.6151
R1297 B.n255 B.n254 10.6151
R1298 B.n254 B.n253 10.6151
R1299 B.n253 B.n213 10.6151
R1300 B.n247 B.n213 10.6151
R1301 B.n247 B.n246 10.6151
R1302 B.n246 B.n245 10.6151
R1303 B.n245 B.n215 10.6151
R1304 B.n239 B.n215 10.6151
R1305 B.n239 B.n238 10.6151
R1306 B.n238 B.n237 10.6151
R1307 B.n237 B.n217 10.6151
R1308 B.n231 B.n217 10.6151
R1309 B.n231 B.n230 10.6151
R1310 B.n230 B.n229 10.6151
R1311 B.n229 B.n219 10.6151
R1312 B.n223 B.n219 10.6151
R1313 B.n223 B.n222 10.6151
R1314 B.n222 B.n143 10.6151
R1315 B.n502 B.n501 10.6151
R1316 B.n503 B.n502 10.6151
R1317 B.n503 B.n134 10.6151
R1318 B.n513 B.n134 10.6151
R1319 B.n514 B.n513 10.6151
R1320 B.n515 B.n514 10.6151
R1321 B.n515 B.n127 10.6151
R1322 B.n525 B.n127 10.6151
R1323 B.n526 B.n525 10.6151
R1324 B.n527 B.n526 10.6151
R1325 B.n527 B.n120 10.6151
R1326 B.n538 B.n120 10.6151
R1327 B.n539 B.n538 10.6151
R1328 B.n541 B.n539 10.6151
R1329 B.n541 B.n540 10.6151
R1330 B.n540 B.n113 10.6151
R1331 B.n553 B.n113 10.6151
R1332 B.n554 B.n553 10.6151
R1333 B.n555 B.n554 10.6151
R1334 B.n556 B.n555 10.6151
R1335 B.n557 B.n556 10.6151
R1336 B.n560 B.n557 10.6151
R1337 B.n561 B.n560 10.6151
R1338 B.n562 B.n561 10.6151
R1339 B.n563 B.n562 10.6151
R1340 B.n565 B.n563 10.6151
R1341 B.n566 B.n565 10.6151
R1342 B.n567 B.n566 10.6151
R1343 B.n568 B.n567 10.6151
R1344 B.n570 B.n568 10.6151
R1345 B.n571 B.n570 10.6151
R1346 B.n572 B.n571 10.6151
R1347 B.n573 B.n572 10.6151
R1348 B.n575 B.n573 10.6151
R1349 B.n576 B.n575 10.6151
R1350 B.n577 B.n576 10.6151
R1351 B.n578 B.n577 10.6151
R1352 B.n889 B.n1 10.6151
R1353 B.n889 B.n888 10.6151
R1354 B.n888 B.n887 10.6151
R1355 B.n887 B.n10 10.6151
R1356 B.n881 B.n10 10.6151
R1357 B.n881 B.n880 10.6151
R1358 B.n880 B.n879 10.6151
R1359 B.n879 B.n17 10.6151
R1360 B.n873 B.n17 10.6151
R1361 B.n873 B.n872 10.6151
R1362 B.n872 B.n871 10.6151
R1363 B.n871 B.n25 10.6151
R1364 B.n865 B.n25 10.6151
R1365 B.n865 B.n864 10.6151
R1366 B.n864 B.n863 10.6151
R1367 B.n863 B.n32 10.6151
R1368 B.n857 B.n32 10.6151
R1369 B.n856 B.n855 10.6151
R1370 B.n855 B.n39 10.6151
R1371 B.n849 B.n39 10.6151
R1372 B.n849 B.n848 10.6151
R1373 B.n848 B.n847 10.6151
R1374 B.n847 B.n41 10.6151
R1375 B.n841 B.n41 10.6151
R1376 B.n841 B.n840 10.6151
R1377 B.n840 B.n839 10.6151
R1378 B.n839 B.n43 10.6151
R1379 B.n833 B.n43 10.6151
R1380 B.n833 B.n832 10.6151
R1381 B.n832 B.n831 10.6151
R1382 B.n831 B.n45 10.6151
R1383 B.n825 B.n45 10.6151
R1384 B.n825 B.n824 10.6151
R1385 B.n824 B.n823 10.6151
R1386 B.n823 B.n47 10.6151
R1387 B.n817 B.n47 10.6151
R1388 B.n817 B.n816 10.6151
R1389 B.n816 B.n815 10.6151
R1390 B.n815 B.n49 10.6151
R1391 B.n809 B.n49 10.6151
R1392 B.n809 B.n808 10.6151
R1393 B.n808 B.n807 10.6151
R1394 B.n807 B.n51 10.6151
R1395 B.n801 B.n51 10.6151
R1396 B.n801 B.n800 10.6151
R1397 B.n800 B.n799 10.6151
R1398 B.n799 B.n53 10.6151
R1399 B.n793 B.n53 10.6151
R1400 B.n793 B.n792 10.6151
R1401 B.n792 B.n791 10.6151
R1402 B.n791 B.n55 10.6151
R1403 B.n785 B.n55 10.6151
R1404 B.n785 B.n784 10.6151
R1405 B.n784 B.n783 10.6151
R1406 B.n783 B.n57 10.6151
R1407 B.n777 B.n57 10.6151
R1408 B.n777 B.n776 10.6151
R1409 B.n776 B.n775 10.6151
R1410 B.n775 B.n59 10.6151
R1411 B.n769 B.n59 10.6151
R1412 B.n769 B.n768 10.6151
R1413 B.n768 B.n767 10.6151
R1414 B.n767 B.n61 10.6151
R1415 B.n761 B.n61 10.6151
R1416 B.n761 B.n760 10.6151
R1417 B.n760 B.n759 10.6151
R1418 B.n759 B.n63 10.6151
R1419 B.n753 B.n63 10.6151
R1420 B.n753 B.n752 10.6151
R1421 B.n752 B.n751 10.6151
R1422 B.n751 B.n65 10.6151
R1423 B.n745 B.n65 10.6151
R1424 B.n745 B.n744 10.6151
R1425 B.n744 B.n743 10.6151
R1426 B.n743 B.n67 10.6151
R1427 B.n737 B.n67 10.6151
R1428 B.n737 B.n736 10.6151
R1429 B.n736 B.n735 10.6151
R1430 B.n735 B.n69 10.6151
R1431 B.n729 B.n69 10.6151
R1432 B.n729 B.n728 10.6151
R1433 B.n726 B.n73 10.6151
R1434 B.n720 B.n73 10.6151
R1435 B.n720 B.n719 10.6151
R1436 B.n719 B.n718 10.6151
R1437 B.n718 B.n75 10.6151
R1438 B.n712 B.n75 10.6151
R1439 B.n712 B.n711 10.6151
R1440 B.n711 B.n710 10.6151
R1441 B.n706 B.n705 10.6151
R1442 B.n705 B.n81 10.6151
R1443 B.n700 B.n81 10.6151
R1444 B.n700 B.n699 10.6151
R1445 B.n699 B.n698 10.6151
R1446 B.n698 B.n83 10.6151
R1447 B.n692 B.n83 10.6151
R1448 B.n692 B.n691 10.6151
R1449 B.n691 B.n690 10.6151
R1450 B.n690 B.n85 10.6151
R1451 B.n684 B.n85 10.6151
R1452 B.n684 B.n683 10.6151
R1453 B.n683 B.n682 10.6151
R1454 B.n682 B.n87 10.6151
R1455 B.n676 B.n87 10.6151
R1456 B.n676 B.n675 10.6151
R1457 B.n675 B.n674 10.6151
R1458 B.n674 B.n89 10.6151
R1459 B.n668 B.n89 10.6151
R1460 B.n668 B.n667 10.6151
R1461 B.n667 B.n666 10.6151
R1462 B.n666 B.n91 10.6151
R1463 B.n660 B.n91 10.6151
R1464 B.n660 B.n659 10.6151
R1465 B.n659 B.n658 10.6151
R1466 B.n658 B.n93 10.6151
R1467 B.n652 B.n93 10.6151
R1468 B.n652 B.n651 10.6151
R1469 B.n651 B.n650 10.6151
R1470 B.n650 B.n95 10.6151
R1471 B.n644 B.n95 10.6151
R1472 B.n644 B.n643 10.6151
R1473 B.n643 B.n642 10.6151
R1474 B.n642 B.n97 10.6151
R1475 B.n636 B.n97 10.6151
R1476 B.n636 B.n635 10.6151
R1477 B.n635 B.n634 10.6151
R1478 B.n634 B.n99 10.6151
R1479 B.n628 B.n99 10.6151
R1480 B.n628 B.n627 10.6151
R1481 B.n627 B.n626 10.6151
R1482 B.n626 B.n101 10.6151
R1483 B.n620 B.n101 10.6151
R1484 B.n620 B.n619 10.6151
R1485 B.n619 B.n618 10.6151
R1486 B.n618 B.n103 10.6151
R1487 B.n612 B.n103 10.6151
R1488 B.n612 B.n611 10.6151
R1489 B.n611 B.n610 10.6151
R1490 B.n610 B.n105 10.6151
R1491 B.n604 B.n105 10.6151
R1492 B.n604 B.n603 10.6151
R1493 B.n603 B.n602 10.6151
R1494 B.n602 B.n107 10.6151
R1495 B.n596 B.n107 10.6151
R1496 B.n596 B.n595 10.6151
R1497 B.n595 B.n594 10.6151
R1498 B.n594 B.n109 10.6151
R1499 B.n588 B.n109 10.6151
R1500 B.n588 B.n587 10.6151
R1501 B.n587 B.n586 10.6151
R1502 B.n586 B.n111 10.6151
R1503 B.n580 B.n111 10.6151
R1504 B.n580 B.n579 10.6151
R1505 B.n897 B.n0 8.11757
R1506 B.n897 B.n1 8.11757
R1507 B.n366 B.n181 6.5566
R1508 B.n351 B.n350 6.5566
R1509 B.n727 B.n726 6.5566
R1510 B.n710 B.n79 6.5566
R1511 B.n536 B.t0 6.54422
R1512 B.n883 B.t2 6.54422
R1513 B.n543 B.t3 5.67173
R1514 B.n12 B.t1 5.67173
R1515 B.n137 B.t5 4.79923
R1516 B.t9 B.n868 4.79923
R1517 B.n370 B.n181 4.05904
R1518 B.n350 B.n349 4.05904
R1519 B.n728 B.n727 4.05904
R1520 B.n706 B.n79 4.05904
R1521 VN.n0 VN.t3 647.888
R1522 VN.n1 VN.t2 647.888
R1523 VN.n0 VN.t0 647.837
R1524 VN.n1 VN.t1 647.837
R1525 VN VN.n1 91.9594
R1526 VN VN.n0 44.7132
R1527 VDD2.n2 VDD2.n0 102.559
R1528 VDD2.n2 VDD2.n1 58.6548
R1529 VDD2.n1 VDD2.t2 0.993479
R1530 VDD2.n1 VDD2.t1 0.993479
R1531 VDD2.n0 VDD2.t0 0.993479
R1532 VDD2.n0 VDD2.t3 0.993479
R1533 VDD2 VDD2.n2 0.0586897
C0 VN VDD2 5.46536f
C1 VN VDD1 0.146874f
C2 VP VTAIL 4.78973f
C3 VDD2 VDD1 0.596448f
C4 VN VTAIL 4.77562f
C5 VDD2 VTAIL 9.66763f
C6 VN VP 6.38638f
C7 VDD2 VP 0.281151f
C8 VDD1 VTAIL 9.62528f
C9 VP VDD1 5.59935f
C10 VDD2 B 3.393764f
C11 VDD1 B 7.9737f
C12 VTAIL B 13.433409f
C13 VN B 9.40114f
C14 VP B 5.706526f
C15 VDD2.t0 B 0.439848f
C16 VDD2.t3 B 0.439848f
C17 VDD2.n0 B 4.952621f
C18 VDD2.t2 B 0.439848f
C19 VDD2.t1 B 0.439848f
C20 VDD2.n1 B 4.01883f
C21 VDD2.n2 B 4.3732f
C22 VN.t3 B 2.18343f
C23 VN.t0 B 2.18337f
C24 VN.n0 B 1.55812f
C25 VN.t2 B 2.18343f
C26 VN.t1 B 2.18337f
C27 VN.n1 B 2.79509f
C28 VDD1.t2 B 0.436884f
C29 VDD1.t3 B 0.436884f
C30 VDD1.n0 B 3.99209f
C31 VDD1.t1 B 0.436884f
C32 VDD1.t0 B 0.436884f
C33 VDD1.n1 B 4.94934f
C34 VTAIL.t1 B 2.77317f
C35 VTAIL.n0 B 0.272171f
C36 VTAIL.t5 B 2.77317f
C37 VTAIL.n1 B 0.294133f
C38 VTAIL.t4 B 2.77317f
C39 VTAIL.n2 B 1.38453f
C40 VTAIL.t0 B 2.77319f
C41 VTAIL.n3 B 1.38451f
C42 VTAIL.t3 B 2.77319f
C43 VTAIL.n4 B 0.294118f
C44 VTAIL.t6 B 2.77319f
C45 VTAIL.n5 B 0.294118f
C46 VTAIL.t7 B 2.77318f
C47 VTAIL.n6 B 1.38452f
C48 VTAIL.t2 B 2.77317f
C49 VTAIL.n7 B 1.35678f
C50 VP.n0 B 0.04647f
C51 VP.t0 B 2.20498f
C52 VP.t1 B 2.20505f
C53 VP.n1 B 2.80233f
C54 VP.n2 B 3.49759f
C55 VP.t2 B 2.17877f
C56 VP.n3 B 0.807497f
C57 VP.n4 B 0.010545f
C58 VP.t3 B 2.17877f
C59 VP.n5 B 0.807497f
C60 VP.n6 B 0.036013f
.ends

