* NGSPICE file created from diff_pair_sample_1459.ext - technology: sky130A

.subckt diff_pair_sample_1459 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t5 VN.t0 VTAIL.t8 w_n1610_n3668# sky130_fd_pr__pfet_01v8 ad=5.265 pd=27.78 as=2.2275 ps=13.83 w=13.5 l=0.47
X1 B.t11 B.t9 B.t10 w_n1610_n3668# sky130_fd_pr__pfet_01v8 ad=5.265 pd=27.78 as=0 ps=0 w=13.5 l=0.47
X2 VDD2.t4 VN.t1 VTAIL.t6 w_n1610_n3668# sky130_fd_pr__pfet_01v8 ad=5.265 pd=27.78 as=2.2275 ps=13.83 w=13.5 l=0.47
X3 VDD1.t5 VP.t0 VTAIL.t5 w_n1610_n3668# sky130_fd_pr__pfet_01v8 ad=5.265 pd=27.78 as=2.2275 ps=13.83 w=13.5 l=0.47
X4 VTAIL.t4 VP.t1 VDD1.t4 w_n1610_n3668# sky130_fd_pr__pfet_01v8 ad=2.2275 pd=13.83 as=2.2275 ps=13.83 w=13.5 l=0.47
X5 VDD2.t3 VN.t2 VTAIL.t10 w_n1610_n3668# sky130_fd_pr__pfet_01v8 ad=2.2275 pd=13.83 as=5.265 ps=27.78 w=13.5 l=0.47
X6 VDD2.t2 VN.t3 VTAIL.t11 w_n1610_n3668# sky130_fd_pr__pfet_01v8 ad=2.2275 pd=13.83 as=5.265 ps=27.78 w=13.5 l=0.47
X7 VTAIL.t7 VN.t4 VDD2.t1 w_n1610_n3668# sky130_fd_pr__pfet_01v8 ad=2.2275 pd=13.83 as=2.2275 ps=13.83 w=13.5 l=0.47
X8 B.t8 B.t6 B.t7 w_n1610_n3668# sky130_fd_pr__pfet_01v8 ad=5.265 pd=27.78 as=0 ps=0 w=13.5 l=0.47
X9 VDD1.t3 VP.t2 VTAIL.t3 w_n1610_n3668# sky130_fd_pr__pfet_01v8 ad=2.2275 pd=13.83 as=5.265 ps=27.78 w=13.5 l=0.47
X10 VTAIL.t0 VP.t3 VDD1.t2 w_n1610_n3668# sky130_fd_pr__pfet_01v8 ad=2.2275 pd=13.83 as=2.2275 ps=13.83 w=13.5 l=0.47
X11 B.t5 B.t3 B.t4 w_n1610_n3668# sky130_fd_pr__pfet_01v8 ad=5.265 pd=27.78 as=0 ps=0 w=13.5 l=0.47
X12 VDD1.t1 VP.t4 VTAIL.t2 w_n1610_n3668# sky130_fd_pr__pfet_01v8 ad=2.2275 pd=13.83 as=5.265 ps=27.78 w=13.5 l=0.47
X13 VTAIL.t9 VN.t5 VDD2.t0 w_n1610_n3668# sky130_fd_pr__pfet_01v8 ad=2.2275 pd=13.83 as=2.2275 ps=13.83 w=13.5 l=0.47
X14 VDD1.t0 VP.t5 VTAIL.t1 w_n1610_n3668# sky130_fd_pr__pfet_01v8 ad=5.265 pd=27.78 as=2.2275 ps=13.83 w=13.5 l=0.47
X15 B.t2 B.t0 B.t1 w_n1610_n3668# sky130_fd_pr__pfet_01v8 ad=5.265 pd=27.78 as=0 ps=0 w=13.5 l=0.47
R0 VN.n0 VN.t1 802.601
R1 VN.n4 VN.t3 802.601
R2 VN.n2 VN.t2 785.309
R3 VN.n6 VN.t0 785.309
R4 VN.n1 VN.t4 775.816
R5 VN.n5 VN.t5 775.816
R6 VN.n3 VN.n2 161.3
R7 VN.n7 VN.n6 161.3
R8 VN.n7 VN.n4 72.2473
R9 VN.n3 VN.n0 72.2473
R10 VN VN.n7 41.9645
R11 VN.n2 VN.n1 38.7066
R12 VN.n6 VN.n5 38.7066
R13 VN.n5 VN.n4 17.2717
R14 VN.n1 VN.n0 17.2717
R15 VN VN.n3 0.0516364
R16 VTAIL.n298 VTAIL.n230 756.745
R17 VTAIL.n70 VTAIL.n2 756.745
R18 VTAIL.n224 VTAIL.n156 756.745
R19 VTAIL.n148 VTAIL.n80 756.745
R20 VTAIL.n255 VTAIL.n254 585
R21 VTAIL.n257 VTAIL.n256 585
R22 VTAIL.n250 VTAIL.n249 585
R23 VTAIL.n263 VTAIL.n262 585
R24 VTAIL.n265 VTAIL.n264 585
R25 VTAIL.n246 VTAIL.n245 585
R26 VTAIL.n272 VTAIL.n271 585
R27 VTAIL.n273 VTAIL.n244 585
R28 VTAIL.n275 VTAIL.n274 585
R29 VTAIL.n242 VTAIL.n241 585
R30 VTAIL.n281 VTAIL.n280 585
R31 VTAIL.n283 VTAIL.n282 585
R32 VTAIL.n238 VTAIL.n237 585
R33 VTAIL.n289 VTAIL.n288 585
R34 VTAIL.n291 VTAIL.n290 585
R35 VTAIL.n234 VTAIL.n233 585
R36 VTAIL.n297 VTAIL.n296 585
R37 VTAIL.n299 VTAIL.n298 585
R38 VTAIL.n27 VTAIL.n26 585
R39 VTAIL.n29 VTAIL.n28 585
R40 VTAIL.n22 VTAIL.n21 585
R41 VTAIL.n35 VTAIL.n34 585
R42 VTAIL.n37 VTAIL.n36 585
R43 VTAIL.n18 VTAIL.n17 585
R44 VTAIL.n44 VTAIL.n43 585
R45 VTAIL.n45 VTAIL.n16 585
R46 VTAIL.n47 VTAIL.n46 585
R47 VTAIL.n14 VTAIL.n13 585
R48 VTAIL.n53 VTAIL.n52 585
R49 VTAIL.n55 VTAIL.n54 585
R50 VTAIL.n10 VTAIL.n9 585
R51 VTAIL.n61 VTAIL.n60 585
R52 VTAIL.n63 VTAIL.n62 585
R53 VTAIL.n6 VTAIL.n5 585
R54 VTAIL.n69 VTAIL.n68 585
R55 VTAIL.n71 VTAIL.n70 585
R56 VTAIL.n225 VTAIL.n224 585
R57 VTAIL.n223 VTAIL.n222 585
R58 VTAIL.n160 VTAIL.n159 585
R59 VTAIL.n217 VTAIL.n216 585
R60 VTAIL.n215 VTAIL.n214 585
R61 VTAIL.n164 VTAIL.n163 585
R62 VTAIL.n209 VTAIL.n208 585
R63 VTAIL.n207 VTAIL.n206 585
R64 VTAIL.n168 VTAIL.n167 585
R65 VTAIL.n172 VTAIL.n170 585
R66 VTAIL.n201 VTAIL.n200 585
R67 VTAIL.n199 VTAIL.n198 585
R68 VTAIL.n174 VTAIL.n173 585
R69 VTAIL.n193 VTAIL.n192 585
R70 VTAIL.n191 VTAIL.n190 585
R71 VTAIL.n178 VTAIL.n177 585
R72 VTAIL.n185 VTAIL.n184 585
R73 VTAIL.n183 VTAIL.n182 585
R74 VTAIL.n149 VTAIL.n148 585
R75 VTAIL.n147 VTAIL.n146 585
R76 VTAIL.n84 VTAIL.n83 585
R77 VTAIL.n141 VTAIL.n140 585
R78 VTAIL.n139 VTAIL.n138 585
R79 VTAIL.n88 VTAIL.n87 585
R80 VTAIL.n133 VTAIL.n132 585
R81 VTAIL.n131 VTAIL.n130 585
R82 VTAIL.n92 VTAIL.n91 585
R83 VTAIL.n96 VTAIL.n94 585
R84 VTAIL.n125 VTAIL.n124 585
R85 VTAIL.n123 VTAIL.n122 585
R86 VTAIL.n98 VTAIL.n97 585
R87 VTAIL.n117 VTAIL.n116 585
R88 VTAIL.n115 VTAIL.n114 585
R89 VTAIL.n102 VTAIL.n101 585
R90 VTAIL.n109 VTAIL.n108 585
R91 VTAIL.n107 VTAIL.n106 585
R92 VTAIL.n253 VTAIL.t10 329.036
R93 VTAIL.n25 VTAIL.t2 329.036
R94 VTAIL.n181 VTAIL.t3 329.036
R95 VTAIL.n105 VTAIL.t11 329.036
R96 VTAIL.n256 VTAIL.n255 171.744
R97 VTAIL.n256 VTAIL.n249 171.744
R98 VTAIL.n263 VTAIL.n249 171.744
R99 VTAIL.n264 VTAIL.n263 171.744
R100 VTAIL.n264 VTAIL.n245 171.744
R101 VTAIL.n272 VTAIL.n245 171.744
R102 VTAIL.n273 VTAIL.n272 171.744
R103 VTAIL.n274 VTAIL.n273 171.744
R104 VTAIL.n274 VTAIL.n241 171.744
R105 VTAIL.n281 VTAIL.n241 171.744
R106 VTAIL.n282 VTAIL.n281 171.744
R107 VTAIL.n282 VTAIL.n237 171.744
R108 VTAIL.n289 VTAIL.n237 171.744
R109 VTAIL.n290 VTAIL.n289 171.744
R110 VTAIL.n290 VTAIL.n233 171.744
R111 VTAIL.n297 VTAIL.n233 171.744
R112 VTAIL.n298 VTAIL.n297 171.744
R113 VTAIL.n28 VTAIL.n27 171.744
R114 VTAIL.n28 VTAIL.n21 171.744
R115 VTAIL.n35 VTAIL.n21 171.744
R116 VTAIL.n36 VTAIL.n35 171.744
R117 VTAIL.n36 VTAIL.n17 171.744
R118 VTAIL.n44 VTAIL.n17 171.744
R119 VTAIL.n45 VTAIL.n44 171.744
R120 VTAIL.n46 VTAIL.n45 171.744
R121 VTAIL.n46 VTAIL.n13 171.744
R122 VTAIL.n53 VTAIL.n13 171.744
R123 VTAIL.n54 VTAIL.n53 171.744
R124 VTAIL.n54 VTAIL.n9 171.744
R125 VTAIL.n61 VTAIL.n9 171.744
R126 VTAIL.n62 VTAIL.n61 171.744
R127 VTAIL.n62 VTAIL.n5 171.744
R128 VTAIL.n69 VTAIL.n5 171.744
R129 VTAIL.n70 VTAIL.n69 171.744
R130 VTAIL.n224 VTAIL.n223 171.744
R131 VTAIL.n223 VTAIL.n159 171.744
R132 VTAIL.n216 VTAIL.n159 171.744
R133 VTAIL.n216 VTAIL.n215 171.744
R134 VTAIL.n215 VTAIL.n163 171.744
R135 VTAIL.n208 VTAIL.n163 171.744
R136 VTAIL.n208 VTAIL.n207 171.744
R137 VTAIL.n207 VTAIL.n167 171.744
R138 VTAIL.n172 VTAIL.n167 171.744
R139 VTAIL.n200 VTAIL.n172 171.744
R140 VTAIL.n200 VTAIL.n199 171.744
R141 VTAIL.n199 VTAIL.n173 171.744
R142 VTAIL.n192 VTAIL.n173 171.744
R143 VTAIL.n192 VTAIL.n191 171.744
R144 VTAIL.n191 VTAIL.n177 171.744
R145 VTAIL.n184 VTAIL.n177 171.744
R146 VTAIL.n184 VTAIL.n183 171.744
R147 VTAIL.n148 VTAIL.n147 171.744
R148 VTAIL.n147 VTAIL.n83 171.744
R149 VTAIL.n140 VTAIL.n83 171.744
R150 VTAIL.n140 VTAIL.n139 171.744
R151 VTAIL.n139 VTAIL.n87 171.744
R152 VTAIL.n132 VTAIL.n87 171.744
R153 VTAIL.n132 VTAIL.n131 171.744
R154 VTAIL.n131 VTAIL.n91 171.744
R155 VTAIL.n96 VTAIL.n91 171.744
R156 VTAIL.n124 VTAIL.n96 171.744
R157 VTAIL.n124 VTAIL.n123 171.744
R158 VTAIL.n123 VTAIL.n97 171.744
R159 VTAIL.n116 VTAIL.n97 171.744
R160 VTAIL.n116 VTAIL.n115 171.744
R161 VTAIL.n115 VTAIL.n101 171.744
R162 VTAIL.n108 VTAIL.n101 171.744
R163 VTAIL.n108 VTAIL.n107 171.744
R164 VTAIL.n255 VTAIL.t10 85.8723
R165 VTAIL.n27 VTAIL.t2 85.8723
R166 VTAIL.n183 VTAIL.t3 85.8723
R167 VTAIL.n107 VTAIL.t11 85.8723
R168 VTAIL.n155 VTAIL.n154 54.4385
R169 VTAIL.n79 VTAIL.n78 54.4385
R170 VTAIL.n1 VTAIL.n0 54.4383
R171 VTAIL.n77 VTAIL.n76 54.4383
R172 VTAIL.n303 VTAIL.n302 31.0217
R173 VTAIL.n75 VTAIL.n74 31.0217
R174 VTAIL.n229 VTAIL.n228 31.0217
R175 VTAIL.n153 VTAIL.n152 31.0217
R176 VTAIL.n79 VTAIL.n77 25.3841
R177 VTAIL.n303 VTAIL.n229 24.6945
R178 VTAIL.n275 VTAIL.n242 13.1884
R179 VTAIL.n47 VTAIL.n14 13.1884
R180 VTAIL.n170 VTAIL.n168 13.1884
R181 VTAIL.n94 VTAIL.n92 13.1884
R182 VTAIL.n276 VTAIL.n244 12.8005
R183 VTAIL.n280 VTAIL.n279 12.8005
R184 VTAIL.n48 VTAIL.n16 12.8005
R185 VTAIL.n52 VTAIL.n51 12.8005
R186 VTAIL.n206 VTAIL.n205 12.8005
R187 VTAIL.n202 VTAIL.n201 12.8005
R188 VTAIL.n130 VTAIL.n129 12.8005
R189 VTAIL.n126 VTAIL.n125 12.8005
R190 VTAIL.n271 VTAIL.n270 12.0247
R191 VTAIL.n283 VTAIL.n240 12.0247
R192 VTAIL.n43 VTAIL.n42 12.0247
R193 VTAIL.n55 VTAIL.n12 12.0247
R194 VTAIL.n209 VTAIL.n166 12.0247
R195 VTAIL.n198 VTAIL.n171 12.0247
R196 VTAIL.n133 VTAIL.n90 12.0247
R197 VTAIL.n122 VTAIL.n95 12.0247
R198 VTAIL.n269 VTAIL.n246 11.249
R199 VTAIL.n284 VTAIL.n238 11.249
R200 VTAIL.n41 VTAIL.n18 11.249
R201 VTAIL.n56 VTAIL.n10 11.249
R202 VTAIL.n210 VTAIL.n164 11.249
R203 VTAIL.n197 VTAIL.n174 11.249
R204 VTAIL.n134 VTAIL.n88 11.249
R205 VTAIL.n121 VTAIL.n98 11.249
R206 VTAIL.n254 VTAIL.n253 10.7239
R207 VTAIL.n26 VTAIL.n25 10.7239
R208 VTAIL.n182 VTAIL.n181 10.7239
R209 VTAIL.n106 VTAIL.n105 10.7239
R210 VTAIL.n266 VTAIL.n265 10.4732
R211 VTAIL.n288 VTAIL.n287 10.4732
R212 VTAIL.n38 VTAIL.n37 10.4732
R213 VTAIL.n60 VTAIL.n59 10.4732
R214 VTAIL.n214 VTAIL.n213 10.4732
R215 VTAIL.n194 VTAIL.n193 10.4732
R216 VTAIL.n138 VTAIL.n137 10.4732
R217 VTAIL.n118 VTAIL.n117 10.4732
R218 VTAIL.n262 VTAIL.n248 9.69747
R219 VTAIL.n291 VTAIL.n236 9.69747
R220 VTAIL.n34 VTAIL.n20 9.69747
R221 VTAIL.n63 VTAIL.n8 9.69747
R222 VTAIL.n217 VTAIL.n162 9.69747
R223 VTAIL.n190 VTAIL.n176 9.69747
R224 VTAIL.n141 VTAIL.n86 9.69747
R225 VTAIL.n114 VTAIL.n100 9.69747
R226 VTAIL.n302 VTAIL.n301 9.45567
R227 VTAIL.n74 VTAIL.n73 9.45567
R228 VTAIL.n228 VTAIL.n227 9.45567
R229 VTAIL.n152 VTAIL.n151 9.45567
R230 VTAIL.n301 VTAIL.n300 9.3005
R231 VTAIL.n295 VTAIL.n294 9.3005
R232 VTAIL.n293 VTAIL.n292 9.3005
R233 VTAIL.n236 VTAIL.n235 9.3005
R234 VTAIL.n287 VTAIL.n286 9.3005
R235 VTAIL.n285 VTAIL.n284 9.3005
R236 VTAIL.n240 VTAIL.n239 9.3005
R237 VTAIL.n279 VTAIL.n278 9.3005
R238 VTAIL.n252 VTAIL.n251 9.3005
R239 VTAIL.n259 VTAIL.n258 9.3005
R240 VTAIL.n261 VTAIL.n260 9.3005
R241 VTAIL.n248 VTAIL.n247 9.3005
R242 VTAIL.n267 VTAIL.n266 9.3005
R243 VTAIL.n269 VTAIL.n268 9.3005
R244 VTAIL.n270 VTAIL.n243 9.3005
R245 VTAIL.n277 VTAIL.n276 9.3005
R246 VTAIL.n232 VTAIL.n231 9.3005
R247 VTAIL.n73 VTAIL.n72 9.3005
R248 VTAIL.n67 VTAIL.n66 9.3005
R249 VTAIL.n65 VTAIL.n64 9.3005
R250 VTAIL.n8 VTAIL.n7 9.3005
R251 VTAIL.n59 VTAIL.n58 9.3005
R252 VTAIL.n57 VTAIL.n56 9.3005
R253 VTAIL.n12 VTAIL.n11 9.3005
R254 VTAIL.n51 VTAIL.n50 9.3005
R255 VTAIL.n24 VTAIL.n23 9.3005
R256 VTAIL.n31 VTAIL.n30 9.3005
R257 VTAIL.n33 VTAIL.n32 9.3005
R258 VTAIL.n20 VTAIL.n19 9.3005
R259 VTAIL.n39 VTAIL.n38 9.3005
R260 VTAIL.n41 VTAIL.n40 9.3005
R261 VTAIL.n42 VTAIL.n15 9.3005
R262 VTAIL.n49 VTAIL.n48 9.3005
R263 VTAIL.n4 VTAIL.n3 9.3005
R264 VTAIL.n180 VTAIL.n179 9.3005
R265 VTAIL.n187 VTAIL.n186 9.3005
R266 VTAIL.n189 VTAIL.n188 9.3005
R267 VTAIL.n176 VTAIL.n175 9.3005
R268 VTAIL.n195 VTAIL.n194 9.3005
R269 VTAIL.n197 VTAIL.n196 9.3005
R270 VTAIL.n171 VTAIL.n169 9.3005
R271 VTAIL.n203 VTAIL.n202 9.3005
R272 VTAIL.n227 VTAIL.n226 9.3005
R273 VTAIL.n158 VTAIL.n157 9.3005
R274 VTAIL.n221 VTAIL.n220 9.3005
R275 VTAIL.n219 VTAIL.n218 9.3005
R276 VTAIL.n162 VTAIL.n161 9.3005
R277 VTAIL.n213 VTAIL.n212 9.3005
R278 VTAIL.n211 VTAIL.n210 9.3005
R279 VTAIL.n166 VTAIL.n165 9.3005
R280 VTAIL.n205 VTAIL.n204 9.3005
R281 VTAIL.n104 VTAIL.n103 9.3005
R282 VTAIL.n111 VTAIL.n110 9.3005
R283 VTAIL.n113 VTAIL.n112 9.3005
R284 VTAIL.n100 VTAIL.n99 9.3005
R285 VTAIL.n119 VTAIL.n118 9.3005
R286 VTAIL.n121 VTAIL.n120 9.3005
R287 VTAIL.n95 VTAIL.n93 9.3005
R288 VTAIL.n127 VTAIL.n126 9.3005
R289 VTAIL.n151 VTAIL.n150 9.3005
R290 VTAIL.n82 VTAIL.n81 9.3005
R291 VTAIL.n145 VTAIL.n144 9.3005
R292 VTAIL.n143 VTAIL.n142 9.3005
R293 VTAIL.n86 VTAIL.n85 9.3005
R294 VTAIL.n137 VTAIL.n136 9.3005
R295 VTAIL.n135 VTAIL.n134 9.3005
R296 VTAIL.n90 VTAIL.n89 9.3005
R297 VTAIL.n129 VTAIL.n128 9.3005
R298 VTAIL.n261 VTAIL.n250 8.92171
R299 VTAIL.n292 VTAIL.n234 8.92171
R300 VTAIL.n33 VTAIL.n22 8.92171
R301 VTAIL.n64 VTAIL.n6 8.92171
R302 VTAIL.n218 VTAIL.n160 8.92171
R303 VTAIL.n189 VTAIL.n178 8.92171
R304 VTAIL.n142 VTAIL.n84 8.92171
R305 VTAIL.n113 VTAIL.n102 8.92171
R306 VTAIL.n258 VTAIL.n257 8.14595
R307 VTAIL.n296 VTAIL.n295 8.14595
R308 VTAIL.n30 VTAIL.n29 8.14595
R309 VTAIL.n68 VTAIL.n67 8.14595
R310 VTAIL.n222 VTAIL.n221 8.14595
R311 VTAIL.n186 VTAIL.n185 8.14595
R312 VTAIL.n146 VTAIL.n145 8.14595
R313 VTAIL.n110 VTAIL.n109 8.14595
R314 VTAIL.n254 VTAIL.n252 7.3702
R315 VTAIL.n299 VTAIL.n232 7.3702
R316 VTAIL.n302 VTAIL.n230 7.3702
R317 VTAIL.n26 VTAIL.n24 7.3702
R318 VTAIL.n71 VTAIL.n4 7.3702
R319 VTAIL.n74 VTAIL.n2 7.3702
R320 VTAIL.n228 VTAIL.n156 7.3702
R321 VTAIL.n225 VTAIL.n158 7.3702
R322 VTAIL.n182 VTAIL.n180 7.3702
R323 VTAIL.n152 VTAIL.n80 7.3702
R324 VTAIL.n149 VTAIL.n82 7.3702
R325 VTAIL.n106 VTAIL.n104 7.3702
R326 VTAIL.n300 VTAIL.n299 6.59444
R327 VTAIL.n300 VTAIL.n230 6.59444
R328 VTAIL.n72 VTAIL.n71 6.59444
R329 VTAIL.n72 VTAIL.n2 6.59444
R330 VTAIL.n226 VTAIL.n156 6.59444
R331 VTAIL.n226 VTAIL.n225 6.59444
R332 VTAIL.n150 VTAIL.n80 6.59444
R333 VTAIL.n150 VTAIL.n149 6.59444
R334 VTAIL.n257 VTAIL.n252 5.81868
R335 VTAIL.n296 VTAIL.n232 5.81868
R336 VTAIL.n29 VTAIL.n24 5.81868
R337 VTAIL.n68 VTAIL.n4 5.81868
R338 VTAIL.n222 VTAIL.n158 5.81868
R339 VTAIL.n185 VTAIL.n180 5.81868
R340 VTAIL.n146 VTAIL.n82 5.81868
R341 VTAIL.n109 VTAIL.n104 5.81868
R342 VTAIL.n258 VTAIL.n250 5.04292
R343 VTAIL.n295 VTAIL.n234 5.04292
R344 VTAIL.n30 VTAIL.n22 5.04292
R345 VTAIL.n67 VTAIL.n6 5.04292
R346 VTAIL.n221 VTAIL.n160 5.04292
R347 VTAIL.n186 VTAIL.n178 5.04292
R348 VTAIL.n145 VTAIL.n84 5.04292
R349 VTAIL.n110 VTAIL.n102 5.04292
R350 VTAIL.n262 VTAIL.n261 4.26717
R351 VTAIL.n292 VTAIL.n291 4.26717
R352 VTAIL.n34 VTAIL.n33 4.26717
R353 VTAIL.n64 VTAIL.n63 4.26717
R354 VTAIL.n218 VTAIL.n217 4.26717
R355 VTAIL.n190 VTAIL.n189 4.26717
R356 VTAIL.n142 VTAIL.n141 4.26717
R357 VTAIL.n114 VTAIL.n113 4.26717
R358 VTAIL.n265 VTAIL.n248 3.49141
R359 VTAIL.n288 VTAIL.n236 3.49141
R360 VTAIL.n37 VTAIL.n20 3.49141
R361 VTAIL.n60 VTAIL.n8 3.49141
R362 VTAIL.n214 VTAIL.n162 3.49141
R363 VTAIL.n193 VTAIL.n176 3.49141
R364 VTAIL.n138 VTAIL.n86 3.49141
R365 VTAIL.n117 VTAIL.n100 3.49141
R366 VTAIL.n266 VTAIL.n246 2.71565
R367 VTAIL.n287 VTAIL.n238 2.71565
R368 VTAIL.n38 VTAIL.n18 2.71565
R369 VTAIL.n59 VTAIL.n10 2.71565
R370 VTAIL.n213 VTAIL.n164 2.71565
R371 VTAIL.n194 VTAIL.n174 2.71565
R372 VTAIL.n137 VTAIL.n88 2.71565
R373 VTAIL.n118 VTAIL.n98 2.71565
R374 VTAIL.n253 VTAIL.n251 2.41282
R375 VTAIL.n25 VTAIL.n23 2.41282
R376 VTAIL.n181 VTAIL.n179 2.41282
R377 VTAIL.n105 VTAIL.n103 2.41282
R378 VTAIL.n0 VTAIL.t6 2.40828
R379 VTAIL.n0 VTAIL.t7 2.40828
R380 VTAIL.n76 VTAIL.t5 2.40828
R381 VTAIL.n76 VTAIL.t0 2.40828
R382 VTAIL.n154 VTAIL.t1 2.40828
R383 VTAIL.n154 VTAIL.t4 2.40828
R384 VTAIL.n78 VTAIL.t8 2.40828
R385 VTAIL.n78 VTAIL.t9 2.40828
R386 VTAIL.n271 VTAIL.n269 1.93989
R387 VTAIL.n284 VTAIL.n283 1.93989
R388 VTAIL.n43 VTAIL.n41 1.93989
R389 VTAIL.n56 VTAIL.n55 1.93989
R390 VTAIL.n210 VTAIL.n209 1.93989
R391 VTAIL.n198 VTAIL.n197 1.93989
R392 VTAIL.n134 VTAIL.n133 1.93989
R393 VTAIL.n122 VTAIL.n121 1.93989
R394 VTAIL.n270 VTAIL.n244 1.16414
R395 VTAIL.n280 VTAIL.n240 1.16414
R396 VTAIL.n42 VTAIL.n16 1.16414
R397 VTAIL.n52 VTAIL.n12 1.16414
R398 VTAIL.n206 VTAIL.n166 1.16414
R399 VTAIL.n201 VTAIL.n171 1.16414
R400 VTAIL.n130 VTAIL.n90 1.16414
R401 VTAIL.n125 VTAIL.n95 1.16414
R402 VTAIL.n155 VTAIL.n153 0.815155
R403 VTAIL.n75 VTAIL.n1 0.815155
R404 VTAIL.n153 VTAIL.n79 0.690155
R405 VTAIL.n229 VTAIL.n155 0.690155
R406 VTAIL.n77 VTAIL.n75 0.690155
R407 VTAIL VTAIL.n303 0.459552
R408 VTAIL.n276 VTAIL.n275 0.388379
R409 VTAIL.n279 VTAIL.n242 0.388379
R410 VTAIL.n48 VTAIL.n47 0.388379
R411 VTAIL.n51 VTAIL.n14 0.388379
R412 VTAIL.n205 VTAIL.n168 0.388379
R413 VTAIL.n202 VTAIL.n170 0.388379
R414 VTAIL.n129 VTAIL.n92 0.388379
R415 VTAIL.n126 VTAIL.n94 0.388379
R416 VTAIL VTAIL.n1 0.231103
R417 VTAIL.n259 VTAIL.n251 0.155672
R418 VTAIL.n260 VTAIL.n259 0.155672
R419 VTAIL.n260 VTAIL.n247 0.155672
R420 VTAIL.n267 VTAIL.n247 0.155672
R421 VTAIL.n268 VTAIL.n267 0.155672
R422 VTAIL.n268 VTAIL.n243 0.155672
R423 VTAIL.n277 VTAIL.n243 0.155672
R424 VTAIL.n278 VTAIL.n277 0.155672
R425 VTAIL.n278 VTAIL.n239 0.155672
R426 VTAIL.n285 VTAIL.n239 0.155672
R427 VTAIL.n286 VTAIL.n285 0.155672
R428 VTAIL.n286 VTAIL.n235 0.155672
R429 VTAIL.n293 VTAIL.n235 0.155672
R430 VTAIL.n294 VTAIL.n293 0.155672
R431 VTAIL.n294 VTAIL.n231 0.155672
R432 VTAIL.n301 VTAIL.n231 0.155672
R433 VTAIL.n31 VTAIL.n23 0.155672
R434 VTAIL.n32 VTAIL.n31 0.155672
R435 VTAIL.n32 VTAIL.n19 0.155672
R436 VTAIL.n39 VTAIL.n19 0.155672
R437 VTAIL.n40 VTAIL.n39 0.155672
R438 VTAIL.n40 VTAIL.n15 0.155672
R439 VTAIL.n49 VTAIL.n15 0.155672
R440 VTAIL.n50 VTAIL.n49 0.155672
R441 VTAIL.n50 VTAIL.n11 0.155672
R442 VTAIL.n57 VTAIL.n11 0.155672
R443 VTAIL.n58 VTAIL.n57 0.155672
R444 VTAIL.n58 VTAIL.n7 0.155672
R445 VTAIL.n65 VTAIL.n7 0.155672
R446 VTAIL.n66 VTAIL.n65 0.155672
R447 VTAIL.n66 VTAIL.n3 0.155672
R448 VTAIL.n73 VTAIL.n3 0.155672
R449 VTAIL.n227 VTAIL.n157 0.155672
R450 VTAIL.n220 VTAIL.n157 0.155672
R451 VTAIL.n220 VTAIL.n219 0.155672
R452 VTAIL.n219 VTAIL.n161 0.155672
R453 VTAIL.n212 VTAIL.n161 0.155672
R454 VTAIL.n212 VTAIL.n211 0.155672
R455 VTAIL.n211 VTAIL.n165 0.155672
R456 VTAIL.n204 VTAIL.n165 0.155672
R457 VTAIL.n204 VTAIL.n203 0.155672
R458 VTAIL.n203 VTAIL.n169 0.155672
R459 VTAIL.n196 VTAIL.n169 0.155672
R460 VTAIL.n196 VTAIL.n195 0.155672
R461 VTAIL.n195 VTAIL.n175 0.155672
R462 VTAIL.n188 VTAIL.n175 0.155672
R463 VTAIL.n188 VTAIL.n187 0.155672
R464 VTAIL.n187 VTAIL.n179 0.155672
R465 VTAIL.n151 VTAIL.n81 0.155672
R466 VTAIL.n144 VTAIL.n81 0.155672
R467 VTAIL.n144 VTAIL.n143 0.155672
R468 VTAIL.n143 VTAIL.n85 0.155672
R469 VTAIL.n136 VTAIL.n85 0.155672
R470 VTAIL.n136 VTAIL.n135 0.155672
R471 VTAIL.n135 VTAIL.n89 0.155672
R472 VTAIL.n128 VTAIL.n89 0.155672
R473 VTAIL.n128 VTAIL.n127 0.155672
R474 VTAIL.n127 VTAIL.n93 0.155672
R475 VTAIL.n120 VTAIL.n93 0.155672
R476 VTAIL.n120 VTAIL.n119 0.155672
R477 VTAIL.n119 VTAIL.n99 0.155672
R478 VTAIL.n112 VTAIL.n99 0.155672
R479 VTAIL.n112 VTAIL.n111 0.155672
R480 VTAIL.n111 VTAIL.n103 0.155672
R481 VDD2.n143 VDD2.n75 756.745
R482 VDD2.n68 VDD2.n0 756.745
R483 VDD2.n144 VDD2.n143 585
R484 VDD2.n142 VDD2.n141 585
R485 VDD2.n79 VDD2.n78 585
R486 VDD2.n136 VDD2.n135 585
R487 VDD2.n134 VDD2.n133 585
R488 VDD2.n83 VDD2.n82 585
R489 VDD2.n128 VDD2.n127 585
R490 VDD2.n126 VDD2.n125 585
R491 VDD2.n87 VDD2.n86 585
R492 VDD2.n91 VDD2.n89 585
R493 VDD2.n120 VDD2.n119 585
R494 VDD2.n118 VDD2.n117 585
R495 VDD2.n93 VDD2.n92 585
R496 VDD2.n112 VDD2.n111 585
R497 VDD2.n110 VDD2.n109 585
R498 VDD2.n97 VDD2.n96 585
R499 VDD2.n104 VDD2.n103 585
R500 VDD2.n102 VDD2.n101 585
R501 VDD2.n25 VDD2.n24 585
R502 VDD2.n27 VDD2.n26 585
R503 VDD2.n20 VDD2.n19 585
R504 VDD2.n33 VDD2.n32 585
R505 VDD2.n35 VDD2.n34 585
R506 VDD2.n16 VDD2.n15 585
R507 VDD2.n42 VDD2.n41 585
R508 VDD2.n43 VDD2.n14 585
R509 VDD2.n45 VDD2.n44 585
R510 VDD2.n12 VDD2.n11 585
R511 VDD2.n51 VDD2.n50 585
R512 VDD2.n53 VDD2.n52 585
R513 VDD2.n8 VDD2.n7 585
R514 VDD2.n59 VDD2.n58 585
R515 VDD2.n61 VDD2.n60 585
R516 VDD2.n4 VDD2.n3 585
R517 VDD2.n67 VDD2.n66 585
R518 VDD2.n69 VDD2.n68 585
R519 VDD2.n100 VDD2.t5 329.036
R520 VDD2.n23 VDD2.t4 329.036
R521 VDD2.n143 VDD2.n142 171.744
R522 VDD2.n142 VDD2.n78 171.744
R523 VDD2.n135 VDD2.n78 171.744
R524 VDD2.n135 VDD2.n134 171.744
R525 VDD2.n134 VDD2.n82 171.744
R526 VDD2.n127 VDD2.n82 171.744
R527 VDD2.n127 VDD2.n126 171.744
R528 VDD2.n126 VDD2.n86 171.744
R529 VDD2.n91 VDD2.n86 171.744
R530 VDD2.n119 VDD2.n91 171.744
R531 VDD2.n119 VDD2.n118 171.744
R532 VDD2.n118 VDD2.n92 171.744
R533 VDD2.n111 VDD2.n92 171.744
R534 VDD2.n111 VDD2.n110 171.744
R535 VDD2.n110 VDD2.n96 171.744
R536 VDD2.n103 VDD2.n96 171.744
R537 VDD2.n103 VDD2.n102 171.744
R538 VDD2.n26 VDD2.n25 171.744
R539 VDD2.n26 VDD2.n19 171.744
R540 VDD2.n33 VDD2.n19 171.744
R541 VDD2.n34 VDD2.n33 171.744
R542 VDD2.n34 VDD2.n15 171.744
R543 VDD2.n42 VDD2.n15 171.744
R544 VDD2.n43 VDD2.n42 171.744
R545 VDD2.n44 VDD2.n43 171.744
R546 VDD2.n44 VDD2.n11 171.744
R547 VDD2.n51 VDD2.n11 171.744
R548 VDD2.n52 VDD2.n51 171.744
R549 VDD2.n52 VDD2.n7 171.744
R550 VDD2.n59 VDD2.n7 171.744
R551 VDD2.n60 VDD2.n59 171.744
R552 VDD2.n60 VDD2.n3 171.744
R553 VDD2.n67 VDD2.n3 171.744
R554 VDD2.n68 VDD2.n67 171.744
R555 VDD2.n102 VDD2.t5 85.8723
R556 VDD2.n25 VDD2.t4 85.8723
R557 VDD2.n74 VDD2.n73 71.2341
R558 VDD2 VDD2.n149 71.2313
R559 VDD2.n74 VDD2.n72 48.1624
R560 VDD2.n148 VDD2.n147 47.7005
R561 VDD2.n148 VDD2.n74 37.5946
R562 VDD2.n89 VDD2.n87 13.1884
R563 VDD2.n45 VDD2.n12 13.1884
R564 VDD2.n125 VDD2.n124 12.8005
R565 VDD2.n121 VDD2.n120 12.8005
R566 VDD2.n46 VDD2.n14 12.8005
R567 VDD2.n50 VDD2.n49 12.8005
R568 VDD2.n128 VDD2.n85 12.0247
R569 VDD2.n117 VDD2.n90 12.0247
R570 VDD2.n41 VDD2.n40 12.0247
R571 VDD2.n53 VDD2.n10 12.0247
R572 VDD2.n129 VDD2.n83 11.249
R573 VDD2.n116 VDD2.n93 11.249
R574 VDD2.n39 VDD2.n16 11.249
R575 VDD2.n54 VDD2.n8 11.249
R576 VDD2.n101 VDD2.n100 10.7239
R577 VDD2.n24 VDD2.n23 10.7239
R578 VDD2.n133 VDD2.n132 10.4732
R579 VDD2.n113 VDD2.n112 10.4732
R580 VDD2.n36 VDD2.n35 10.4732
R581 VDD2.n58 VDD2.n57 10.4732
R582 VDD2.n136 VDD2.n81 9.69747
R583 VDD2.n109 VDD2.n95 9.69747
R584 VDD2.n32 VDD2.n18 9.69747
R585 VDD2.n61 VDD2.n6 9.69747
R586 VDD2.n147 VDD2.n146 9.45567
R587 VDD2.n72 VDD2.n71 9.45567
R588 VDD2.n99 VDD2.n98 9.3005
R589 VDD2.n106 VDD2.n105 9.3005
R590 VDD2.n108 VDD2.n107 9.3005
R591 VDD2.n95 VDD2.n94 9.3005
R592 VDD2.n114 VDD2.n113 9.3005
R593 VDD2.n116 VDD2.n115 9.3005
R594 VDD2.n90 VDD2.n88 9.3005
R595 VDD2.n122 VDD2.n121 9.3005
R596 VDD2.n146 VDD2.n145 9.3005
R597 VDD2.n77 VDD2.n76 9.3005
R598 VDD2.n140 VDD2.n139 9.3005
R599 VDD2.n138 VDD2.n137 9.3005
R600 VDD2.n81 VDD2.n80 9.3005
R601 VDD2.n132 VDD2.n131 9.3005
R602 VDD2.n130 VDD2.n129 9.3005
R603 VDD2.n85 VDD2.n84 9.3005
R604 VDD2.n124 VDD2.n123 9.3005
R605 VDD2.n71 VDD2.n70 9.3005
R606 VDD2.n65 VDD2.n64 9.3005
R607 VDD2.n63 VDD2.n62 9.3005
R608 VDD2.n6 VDD2.n5 9.3005
R609 VDD2.n57 VDD2.n56 9.3005
R610 VDD2.n55 VDD2.n54 9.3005
R611 VDD2.n10 VDD2.n9 9.3005
R612 VDD2.n49 VDD2.n48 9.3005
R613 VDD2.n22 VDD2.n21 9.3005
R614 VDD2.n29 VDD2.n28 9.3005
R615 VDD2.n31 VDD2.n30 9.3005
R616 VDD2.n18 VDD2.n17 9.3005
R617 VDD2.n37 VDD2.n36 9.3005
R618 VDD2.n39 VDD2.n38 9.3005
R619 VDD2.n40 VDD2.n13 9.3005
R620 VDD2.n47 VDD2.n46 9.3005
R621 VDD2.n2 VDD2.n1 9.3005
R622 VDD2.n137 VDD2.n79 8.92171
R623 VDD2.n108 VDD2.n97 8.92171
R624 VDD2.n31 VDD2.n20 8.92171
R625 VDD2.n62 VDD2.n4 8.92171
R626 VDD2.n141 VDD2.n140 8.14595
R627 VDD2.n105 VDD2.n104 8.14595
R628 VDD2.n28 VDD2.n27 8.14595
R629 VDD2.n66 VDD2.n65 8.14595
R630 VDD2.n147 VDD2.n75 7.3702
R631 VDD2.n144 VDD2.n77 7.3702
R632 VDD2.n101 VDD2.n99 7.3702
R633 VDD2.n24 VDD2.n22 7.3702
R634 VDD2.n69 VDD2.n2 7.3702
R635 VDD2.n72 VDD2.n0 7.3702
R636 VDD2.n145 VDD2.n75 6.59444
R637 VDD2.n145 VDD2.n144 6.59444
R638 VDD2.n70 VDD2.n69 6.59444
R639 VDD2.n70 VDD2.n0 6.59444
R640 VDD2.n141 VDD2.n77 5.81868
R641 VDD2.n104 VDD2.n99 5.81868
R642 VDD2.n27 VDD2.n22 5.81868
R643 VDD2.n66 VDD2.n2 5.81868
R644 VDD2.n140 VDD2.n79 5.04292
R645 VDD2.n105 VDD2.n97 5.04292
R646 VDD2.n28 VDD2.n20 5.04292
R647 VDD2.n65 VDD2.n4 5.04292
R648 VDD2.n137 VDD2.n136 4.26717
R649 VDD2.n109 VDD2.n108 4.26717
R650 VDD2.n32 VDD2.n31 4.26717
R651 VDD2.n62 VDD2.n61 4.26717
R652 VDD2.n133 VDD2.n81 3.49141
R653 VDD2.n112 VDD2.n95 3.49141
R654 VDD2.n35 VDD2.n18 3.49141
R655 VDD2.n58 VDD2.n6 3.49141
R656 VDD2.n132 VDD2.n83 2.71565
R657 VDD2.n113 VDD2.n93 2.71565
R658 VDD2.n36 VDD2.n16 2.71565
R659 VDD2.n57 VDD2.n8 2.71565
R660 VDD2.n100 VDD2.n98 2.41282
R661 VDD2.n23 VDD2.n21 2.41282
R662 VDD2.n149 VDD2.t0 2.40828
R663 VDD2.n149 VDD2.t2 2.40828
R664 VDD2.n73 VDD2.t1 2.40828
R665 VDD2.n73 VDD2.t3 2.40828
R666 VDD2.n129 VDD2.n128 1.93989
R667 VDD2.n117 VDD2.n116 1.93989
R668 VDD2.n41 VDD2.n39 1.93989
R669 VDD2.n54 VDD2.n53 1.93989
R670 VDD2.n125 VDD2.n85 1.16414
R671 VDD2.n120 VDD2.n90 1.16414
R672 VDD2.n40 VDD2.n14 1.16414
R673 VDD2.n50 VDD2.n10 1.16414
R674 VDD2 VDD2.n148 0.575931
R675 VDD2.n124 VDD2.n87 0.388379
R676 VDD2.n121 VDD2.n89 0.388379
R677 VDD2.n46 VDD2.n45 0.388379
R678 VDD2.n49 VDD2.n12 0.388379
R679 VDD2.n146 VDD2.n76 0.155672
R680 VDD2.n139 VDD2.n76 0.155672
R681 VDD2.n139 VDD2.n138 0.155672
R682 VDD2.n138 VDD2.n80 0.155672
R683 VDD2.n131 VDD2.n80 0.155672
R684 VDD2.n131 VDD2.n130 0.155672
R685 VDD2.n130 VDD2.n84 0.155672
R686 VDD2.n123 VDD2.n84 0.155672
R687 VDD2.n123 VDD2.n122 0.155672
R688 VDD2.n122 VDD2.n88 0.155672
R689 VDD2.n115 VDD2.n88 0.155672
R690 VDD2.n115 VDD2.n114 0.155672
R691 VDD2.n114 VDD2.n94 0.155672
R692 VDD2.n107 VDD2.n94 0.155672
R693 VDD2.n107 VDD2.n106 0.155672
R694 VDD2.n106 VDD2.n98 0.155672
R695 VDD2.n29 VDD2.n21 0.155672
R696 VDD2.n30 VDD2.n29 0.155672
R697 VDD2.n30 VDD2.n17 0.155672
R698 VDD2.n37 VDD2.n17 0.155672
R699 VDD2.n38 VDD2.n37 0.155672
R700 VDD2.n38 VDD2.n13 0.155672
R701 VDD2.n47 VDD2.n13 0.155672
R702 VDD2.n48 VDD2.n47 0.155672
R703 VDD2.n48 VDD2.n9 0.155672
R704 VDD2.n55 VDD2.n9 0.155672
R705 VDD2.n56 VDD2.n55 0.155672
R706 VDD2.n56 VDD2.n5 0.155672
R707 VDD2.n63 VDD2.n5 0.155672
R708 VDD2.n64 VDD2.n63 0.155672
R709 VDD2.n64 VDD2.n1 0.155672
R710 VDD2.n71 VDD2.n1 0.155672
R711 B.n113 B.t6 899.412
R712 B.n253 B.t9 899.412
R713 B.n42 B.t3 899.412
R714 B.n34 B.t0 899.412
R715 B.n326 B.n325 585
R716 B.n324 B.n85 585
R717 B.n323 B.n322 585
R718 B.n321 B.n86 585
R719 B.n320 B.n319 585
R720 B.n318 B.n87 585
R721 B.n317 B.n316 585
R722 B.n315 B.n88 585
R723 B.n314 B.n313 585
R724 B.n312 B.n89 585
R725 B.n311 B.n310 585
R726 B.n309 B.n90 585
R727 B.n308 B.n307 585
R728 B.n306 B.n91 585
R729 B.n305 B.n304 585
R730 B.n303 B.n92 585
R731 B.n302 B.n301 585
R732 B.n300 B.n93 585
R733 B.n299 B.n298 585
R734 B.n297 B.n94 585
R735 B.n296 B.n295 585
R736 B.n294 B.n95 585
R737 B.n293 B.n292 585
R738 B.n291 B.n96 585
R739 B.n290 B.n289 585
R740 B.n288 B.n97 585
R741 B.n287 B.n286 585
R742 B.n285 B.n98 585
R743 B.n284 B.n283 585
R744 B.n282 B.n99 585
R745 B.n281 B.n280 585
R746 B.n279 B.n100 585
R747 B.n278 B.n277 585
R748 B.n276 B.n101 585
R749 B.n275 B.n274 585
R750 B.n273 B.n102 585
R751 B.n272 B.n271 585
R752 B.n270 B.n103 585
R753 B.n269 B.n268 585
R754 B.n267 B.n104 585
R755 B.n266 B.n265 585
R756 B.n264 B.n105 585
R757 B.n263 B.n262 585
R758 B.n261 B.n106 585
R759 B.n260 B.n259 585
R760 B.n258 B.n107 585
R761 B.n257 B.n256 585
R762 B.n252 B.n108 585
R763 B.n251 B.n250 585
R764 B.n249 B.n109 585
R765 B.n248 B.n247 585
R766 B.n246 B.n110 585
R767 B.n245 B.n244 585
R768 B.n243 B.n111 585
R769 B.n242 B.n241 585
R770 B.n240 B.n112 585
R771 B.n238 B.n237 585
R772 B.n236 B.n115 585
R773 B.n235 B.n234 585
R774 B.n233 B.n116 585
R775 B.n232 B.n231 585
R776 B.n230 B.n117 585
R777 B.n229 B.n228 585
R778 B.n227 B.n118 585
R779 B.n226 B.n225 585
R780 B.n224 B.n119 585
R781 B.n223 B.n222 585
R782 B.n221 B.n120 585
R783 B.n220 B.n219 585
R784 B.n218 B.n121 585
R785 B.n217 B.n216 585
R786 B.n215 B.n122 585
R787 B.n214 B.n213 585
R788 B.n212 B.n123 585
R789 B.n211 B.n210 585
R790 B.n209 B.n124 585
R791 B.n208 B.n207 585
R792 B.n206 B.n125 585
R793 B.n205 B.n204 585
R794 B.n203 B.n126 585
R795 B.n202 B.n201 585
R796 B.n200 B.n127 585
R797 B.n199 B.n198 585
R798 B.n197 B.n128 585
R799 B.n196 B.n195 585
R800 B.n194 B.n129 585
R801 B.n193 B.n192 585
R802 B.n191 B.n130 585
R803 B.n190 B.n189 585
R804 B.n188 B.n131 585
R805 B.n187 B.n186 585
R806 B.n185 B.n132 585
R807 B.n184 B.n183 585
R808 B.n182 B.n133 585
R809 B.n181 B.n180 585
R810 B.n179 B.n134 585
R811 B.n178 B.n177 585
R812 B.n176 B.n135 585
R813 B.n175 B.n174 585
R814 B.n173 B.n136 585
R815 B.n172 B.n171 585
R816 B.n170 B.n137 585
R817 B.n327 B.n84 585
R818 B.n329 B.n328 585
R819 B.n330 B.n83 585
R820 B.n332 B.n331 585
R821 B.n333 B.n82 585
R822 B.n335 B.n334 585
R823 B.n336 B.n81 585
R824 B.n338 B.n337 585
R825 B.n339 B.n80 585
R826 B.n341 B.n340 585
R827 B.n342 B.n79 585
R828 B.n344 B.n343 585
R829 B.n345 B.n78 585
R830 B.n347 B.n346 585
R831 B.n348 B.n77 585
R832 B.n350 B.n349 585
R833 B.n351 B.n76 585
R834 B.n353 B.n352 585
R835 B.n354 B.n75 585
R836 B.n356 B.n355 585
R837 B.n357 B.n74 585
R838 B.n359 B.n358 585
R839 B.n360 B.n73 585
R840 B.n362 B.n361 585
R841 B.n363 B.n72 585
R842 B.n365 B.n364 585
R843 B.n366 B.n71 585
R844 B.n368 B.n367 585
R845 B.n369 B.n70 585
R846 B.n371 B.n370 585
R847 B.n372 B.n69 585
R848 B.n374 B.n373 585
R849 B.n375 B.n68 585
R850 B.n377 B.n376 585
R851 B.n378 B.n67 585
R852 B.n380 B.n379 585
R853 B.n534 B.n533 585
R854 B.n532 B.n11 585
R855 B.n531 B.n530 585
R856 B.n529 B.n12 585
R857 B.n528 B.n527 585
R858 B.n526 B.n13 585
R859 B.n525 B.n524 585
R860 B.n523 B.n14 585
R861 B.n522 B.n521 585
R862 B.n520 B.n15 585
R863 B.n519 B.n518 585
R864 B.n517 B.n16 585
R865 B.n516 B.n515 585
R866 B.n514 B.n17 585
R867 B.n513 B.n512 585
R868 B.n511 B.n18 585
R869 B.n510 B.n509 585
R870 B.n508 B.n19 585
R871 B.n507 B.n506 585
R872 B.n505 B.n20 585
R873 B.n504 B.n503 585
R874 B.n502 B.n21 585
R875 B.n501 B.n500 585
R876 B.n499 B.n22 585
R877 B.n498 B.n497 585
R878 B.n496 B.n23 585
R879 B.n495 B.n494 585
R880 B.n493 B.n24 585
R881 B.n492 B.n491 585
R882 B.n490 B.n25 585
R883 B.n489 B.n488 585
R884 B.n487 B.n26 585
R885 B.n486 B.n485 585
R886 B.n484 B.n27 585
R887 B.n483 B.n482 585
R888 B.n481 B.n28 585
R889 B.n480 B.n479 585
R890 B.n478 B.n29 585
R891 B.n477 B.n476 585
R892 B.n475 B.n30 585
R893 B.n474 B.n473 585
R894 B.n472 B.n31 585
R895 B.n471 B.n470 585
R896 B.n469 B.n32 585
R897 B.n468 B.n467 585
R898 B.n466 B.n33 585
R899 B.n464 B.n463 585
R900 B.n462 B.n36 585
R901 B.n461 B.n460 585
R902 B.n459 B.n37 585
R903 B.n458 B.n457 585
R904 B.n456 B.n38 585
R905 B.n455 B.n454 585
R906 B.n453 B.n39 585
R907 B.n452 B.n451 585
R908 B.n450 B.n40 585
R909 B.n449 B.n448 585
R910 B.n447 B.n41 585
R911 B.n446 B.n445 585
R912 B.n444 B.n45 585
R913 B.n443 B.n442 585
R914 B.n441 B.n46 585
R915 B.n440 B.n439 585
R916 B.n438 B.n47 585
R917 B.n437 B.n436 585
R918 B.n435 B.n48 585
R919 B.n434 B.n433 585
R920 B.n432 B.n49 585
R921 B.n431 B.n430 585
R922 B.n429 B.n50 585
R923 B.n428 B.n427 585
R924 B.n426 B.n51 585
R925 B.n425 B.n424 585
R926 B.n423 B.n52 585
R927 B.n422 B.n421 585
R928 B.n420 B.n53 585
R929 B.n419 B.n418 585
R930 B.n417 B.n54 585
R931 B.n416 B.n415 585
R932 B.n414 B.n55 585
R933 B.n413 B.n412 585
R934 B.n411 B.n56 585
R935 B.n410 B.n409 585
R936 B.n408 B.n57 585
R937 B.n407 B.n406 585
R938 B.n405 B.n58 585
R939 B.n404 B.n403 585
R940 B.n402 B.n59 585
R941 B.n401 B.n400 585
R942 B.n399 B.n60 585
R943 B.n398 B.n397 585
R944 B.n396 B.n61 585
R945 B.n395 B.n394 585
R946 B.n393 B.n62 585
R947 B.n392 B.n391 585
R948 B.n390 B.n63 585
R949 B.n389 B.n388 585
R950 B.n387 B.n64 585
R951 B.n386 B.n385 585
R952 B.n384 B.n65 585
R953 B.n383 B.n382 585
R954 B.n381 B.n66 585
R955 B.n535 B.n10 585
R956 B.n537 B.n536 585
R957 B.n538 B.n9 585
R958 B.n540 B.n539 585
R959 B.n541 B.n8 585
R960 B.n543 B.n542 585
R961 B.n544 B.n7 585
R962 B.n546 B.n545 585
R963 B.n547 B.n6 585
R964 B.n549 B.n548 585
R965 B.n550 B.n5 585
R966 B.n552 B.n551 585
R967 B.n553 B.n4 585
R968 B.n555 B.n554 585
R969 B.n556 B.n3 585
R970 B.n558 B.n557 585
R971 B.n559 B.n0 585
R972 B.n2 B.n1 585
R973 B.n146 B.n145 585
R974 B.n148 B.n147 585
R975 B.n149 B.n144 585
R976 B.n151 B.n150 585
R977 B.n152 B.n143 585
R978 B.n154 B.n153 585
R979 B.n155 B.n142 585
R980 B.n157 B.n156 585
R981 B.n158 B.n141 585
R982 B.n160 B.n159 585
R983 B.n161 B.n140 585
R984 B.n163 B.n162 585
R985 B.n164 B.n139 585
R986 B.n166 B.n165 585
R987 B.n167 B.n138 585
R988 B.n169 B.n168 585
R989 B.n170 B.n169 473.281
R990 B.n325 B.n84 473.281
R991 B.n379 B.n66 473.281
R992 B.n535 B.n534 473.281
R993 B.n253 B.t10 418.255
R994 B.n42 B.t5 418.255
R995 B.n113 B.t7 418.255
R996 B.n34 B.t2 418.255
R997 B.n254 B.t11 402.74
R998 B.n43 B.t4 402.74
R999 B.n114 B.t8 402.74
R1000 B.n35 B.t1 402.74
R1001 B.n561 B.n560 256.663
R1002 B.n560 B.n559 235.042
R1003 B.n560 B.n2 235.042
R1004 B.n171 B.n170 163.367
R1005 B.n171 B.n136 163.367
R1006 B.n175 B.n136 163.367
R1007 B.n176 B.n175 163.367
R1008 B.n177 B.n176 163.367
R1009 B.n177 B.n134 163.367
R1010 B.n181 B.n134 163.367
R1011 B.n182 B.n181 163.367
R1012 B.n183 B.n182 163.367
R1013 B.n183 B.n132 163.367
R1014 B.n187 B.n132 163.367
R1015 B.n188 B.n187 163.367
R1016 B.n189 B.n188 163.367
R1017 B.n189 B.n130 163.367
R1018 B.n193 B.n130 163.367
R1019 B.n194 B.n193 163.367
R1020 B.n195 B.n194 163.367
R1021 B.n195 B.n128 163.367
R1022 B.n199 B.n128 163.367
R1023 B.n200 B.n199 163.367
R1024 B.n201 B.n200 163.367
R1025 B.n201 B.n126 163.367
R1026 B.n205 B.n126 163.367
R1027 B.n206 B.n205 163.367
R1028 B.n207 B.n206 163.367
R1029 B.n207 B.n124 163.367
R1030 B.n211 B.n124 163.367
R1031 B.n212 B.n211 163.367
R1032 B.n213 B.n212 163.367
R1033 B.n213 B.n122 163.367
R1034 B.n217 B.n122 163.367
R1035 B.n218 B.n217 163.367
R1036 B.n219 B.n218 163.367
R1037 B.n219 B.n120 163.367
R1038 B.n223 B.n120 163.367
R1039 B.n224 B.n223 163.367
R1040 B.n225 B.n224 163.367
R1041 B.n225 B.n118 163.367
R1042 B.n229 B.n118 163.367
R1043 B.n230 B.n229 163.367
R1044 B.n231 B.n230 163.367
R1045 B.n231 B.n116 163.367
R1046 B.n235 B.n116 163.367
R1047 B.n236 B.n235 163.367
R1048 B.n237 B.n236 163.367
R1049 B.n237 B.n112 163.367
R1050 B.n242 B.n112 163.367
R1051 B.n243 B.n242 163.367
R1052 B.n244 B.n243 163.367
R1053 B.n244 B.n110 163.367
R1054 B.n248 B.n110 163.367
R1055 B.n249 B.n248 163.367
R1056 B.n250 B.n249 163.367
R1057 B.n250 B.n108 163.367
R1058 B.n257 B.n108 163.367
R1059 B.n258 B.n257 163.367
R1060 B.n259 B.n258 163.367
R1061 B.n259 B.n106 163.367
R1062 B.n263 B.n106 163.367
R1063 B.n264 B.n263 163.367
R1064 B.n265 B.n264 163.367
R1065 B.n265 B.n104 163.367
R1066 B.n269 B.n104 163.367
R1067 B.n270 B.n269 163.367
R1068 B.n271 B.n270 163.367
R1069 B.n271 B.n102 163.367
R1070 B.n275 B.n102 163.367
R1071 B.n276 B.n275 163.367
R1072 B.n277 B.n276 163.367
R1073 B.n277 B.n100 163.367
R1074 B.n281 B.n100 163.367
R1075 B.n282 B.n281 163.367
R1076 B.n283 B.n282 163.367
R1077 B.n283 B.n98 163.367
R1078 B.n287 B.n98 163.367
R1079 B.n288 B.n287 163.367
R1080 B.n289 B.n288 163.367
R1081 B.n289 B.n96 163.367
R1082 B.n293 B.n96 163.367
R1083 B.n294 B.n293 163.367
R1084 B.n295 B.n294 163.367
R1085 B.n295 B.n94 163.367
R1086 B.n299 B.n94 163.367
R1087 B.n300 B.n299 163.367
R1088 B.n301 B.n300 163.367
R1089 B.n301 B.n92 163.367
R1090 B.n305 B.n92 163.367
R1091 B.n306 B.n305 163.367
R1092 B.n307 B.n306 163.367
R1093 B.n307 B.n90 163.367
R1094 B.n311 B.n90 163.367
R1095 B.n312 B.n311 163.367
R1096 B.n313 B.n312 163.367
R1097 B.n313 B.n88 163.367
R1098 B.n317 B.n88 163.367
R1099 B.n318 B.n317 163.367
R1100 B.n319 B.n318 163.367
R1101 B.n319 B.n86 163.367
R1102 B.n323 B.n86 163.367
R1103 B.n324 B.n323 163.367
R1104 B.n325 B.n324 163.367
R1105 B.n379 B.n378 163.367
R1106 B.n378 B.n377 163.367
R1107 B.n377 B.n68 163.367
R1108 B.n373 B.n68 163.367
R1109 B.n373 B.n372 163.367
R1110 B.n372 B.n371 163.367
R1111 B.n371 B.n70 163.367
R1112 B.n367 B.n70 163.367
R1113 B.n367 B.n366 163.367
R1114 B.n366 B.n365 163.367
R1115 B.n365 B.n72 163.367
R1116 B.n361 B.n72 163.367
R1117 B.n361 B.n360 163.367
R1118 B.n360 B.n359 163.367
R1119 B.n359 B.n74 163.367
R1120 B.n355 B.n74 163.367
R1121 B.n355 B.n354 163.367
R1122 B.n354 B.n353 163.367
R1123 B.n353 B.n76 163.367
R1124 B.n349 B.n76 163.367
R1125 B.n349 B.n348 163.367
R1126 B.n348 B.n347 163.367
R1127 B.n347 B.n78 163.367
R1128 B.n343 B.n78 163.367
R1129 B.n343 B.n342 163.367
R1130 B.n342 B.n341 163.367
R1131 B.n341 B.n80 163.367
R1132 B.n337 B.n80 163.367
R1133 B.n337 B.n336 163.367
R1134 B.n336 B.n335 163.367
R1135 B.n335 B.n82 163.367
R1136 B.n331 B.n82 163.367
R1137 B.n331 B.n330 163.367
R1138 B.n330 B.n329 163.367
R1139 B.n329 B.n84 163.367
R1140 B.n534 B.n11 163.367
R1141 B.n530 B.n11 163.367
R1142 B.n530 B.n529 163.367
R1143 B.n529 B.n528 163.367
R1144 B.n528 B.n13 163.367
R1145 B.n524 B.n13 163.367
R1146 B.n524 B.n523 163.367
R1147 B.n523 B.n522 163.367
R1148 B.n522 B.n15 163.367
R1149 B.n518 B.n15 163.367
R1150 B.n518 B.n517 163.367
R1151 B.n517 B.n516 163.367
R1152 B.n516 B.n17 163.367
R1153 B.n512 B.n17 163.367
R1154 B.n512 B.n511 163.367
R1155 B.n511 B.n510 163.367
R1156 B.n510 B.n19 163.367
R1157 B.n506 B.n19 163.367
R1158 B.n506 B.n505 163.367
R1159 B.n505 B.n504 163.367
R1160 B.n504 B.n21 163.367
R1161 B.n500 B.n21 163.367
R1162 B.n500 B.n499 163.367
R1163 B.n499 B.n498 163.367
R1164 B.n498 B.n23 163.367
R1165 B.n494 B.n23 163.367
R1166 B.n494 B.n493 163.367
R1167 B.n493 B.n492 163.367
R1168 B.n492 B.n25 163.367
R1169 B.n488 B.n25 163.367
R1170 B.n488 B.n487 163.367
R1171 B.n487 B.n486 163.367
R1172 B.n486 B.n27 163.367
R1173 B.n482 B.n27 163.367
R1174 B.n482 B.n481 163.367
R1175 B.n481 B.n480 163.367
R1176 B.n480 B.n29 163.367
R1177 B.n476 B.n29 163.367
R1178 B.n476 B.n475 163.367
R1179 B.n475 B.n474 163.367
R1180 B.n474 B.n31 163.367
R1181 B.n470 B.n31 163.367
R1182 B.n470 B.n469 163.367
R1183 B.n469 B.n468 163.367
R1184 B.n468 B.n33 163.367
R1185 B.n463 B.n33 163.367
R1186 B.n463 B.n462 163.367
R1187 B.n462 B.n461 163.367
R1188 B.n461 B.n37 163.367
R1189 B.n457 B.n37 163.367
R1190 B.n457 B.n456 163.367
R1191 B.n456 B.n455 163.367
R1192 B.n455 B.n39 163.367
R1193 B.n451 B.n39 163.367
R1194 B.n451 B.n450 163.367
R1195 B.n450 B.n449 163.367
R1196 B.n449 B.n41 163.367
R1197 B.n445 B.n41 163.367
R1198 B.n445 B.n444 163.367
R1199 B.n444 B.n443 163.367
R1200 B.n443 B.n46 163.367
R1201 B.n439 B.n46 163.367
R1202 B.n439 B.n438 163.367
R1203 B.n438 B.n437 163.367
R1204 B.n437 B.n48 163.367
R1205 B.n433 B.n48 163.367
R1206 B.n433 B.n432 163.367
R1207 B.n432 B.n431 163.367
R1208 B.n431 B.n50 163.367
R1209 B.n427 B.n50 163.367
R1210 B.n427 B.n426 163.367
R1211 B.n426 B.n425 163.367
R1212 B.n425 B.n52 163.367
R1213 B.n421 B.n52 163.367
R1214 B.n421 B.n420 163.367
R1215 B.n420 B.n419 163.367
R1216 B.n419 B.n54 163.367
R1217 B.n415 B.n54 163.367
R1218 B.n415 B.n414 163.367
R1219 B.n414 B.n413 163.367
R1220 B.n413 B.n56 163.367
R1221 B.n409 B.n56 163.367
R1222 B.n409 B.n408 163.367
R1223 B.n408 B.n407 163.367
R1224 B.n407 B.n58 163.367
R1225 B.n403 B.n58 163.367
R1226 B.n403 B.n402 163.367
R1227 B.n402 B.n401 163.367
R1228 B.n401 B.n60 163.367
R1229 B.n397 B.n60 163.367
R1230 B.n397 B.n396 163.367
R1231 B.n396 B.n395 163.367
R1232 B.n395 B.n62 163.367
R1233 B.n391 B.n62 163.367
R1234 B.n391 B.n390 163.367
R1235 B.n390 B.n389 163.367
R1236 B.n389 B.n64 163.367
R1237 B.n385 B.n64 163.367
R1238 B.n385 B.n384 163.367
R1239 B.n384 B.n383 163.367
R1240 B.n383 B.n66 163.367
R1241 B.n536 B.n535 163.367
R1242 B.n536 B.n9 163.367
R1243 B.n540 B.n9 163.367
R1244 B.n541 B.n540 163.367
R1245 B.n542 B.n541 163.367
R1246 B.n542 B.n7 163.367
R1247 B.n546 B.n7 163.367
R1248 B.n547 B.n546 163.367
R1249 B.n548 B.n547 163.367
R1250 B.n548 B.n5 163.367
R1251 B.n552 B.n5 163.367
R1252 B.n553 B.n552 163.367
R1253 B.n554 B.n553 163.367
R1254 B.n554 B.n3 163.367
R1255 B.n558 B.n3 163.367
R1256 B.n559 B.n558 163.367
R1257 B.n146 B.n2 163.367
R1258 B.n147 B.n146 163.367
R1259 B.n147 B.n144 163.367
R1260 B.n151 B.n144 163.367
R1261 B.n152 B.n151 163.367
R1262 B.n153 B.n152 163.367
R1263 B.n153 B.n142 163.367
R1264 B.n157 B.n142 163.367
R1265 B.n158 B.n157 163.367
R1266 B.n159 B.n158 163.367
R1267 B.n159 B.n140 163.367
R1268 B.n163 B.n140 163.367
R1269 B.n164 B.n163 163.367
R1270 B.n165 B.n164 163.367
R1271 B.n165 B.n138 163.367
R1272 B.n169 B.n138 163.367
R1273 B.n239 B.n114 59.5399
R1274 B.n255 B.n254 59.5399
R1275 B.n44 B.n43 59.5399
R1276 B.n465 B.n35 59.5399
R1277 B.n533 B.n10 30.7517
R1278 B.n381 B.n380 30.7517
R1279 B.n327 B.n326 30.7517
R1280 B.n168 B.n137 30.7517
R1281 B B.n561 18.0485
R1282 B.n114 B.n113 15.5157
R1283 B.n254 B.n253 15.5157
R1284 B.n43 B.n42 15.5157
R1285 B.n35 B.n34 15.5157
R1286 B.n537 B.n10 10.6151
R1287 B.n538 B.n537 10.6151
R1288 B.n539 B.n538 10.6151
R1289 B.n539 B.n8 10.6151
R1290 B.n543 B.n8 10.6151
R1291 B.n544 B.n543 10.6151
R1292 B.n545 B.n544 10.6151
R1293 B.n545 B.n6 10.6151
R1294 B.n549 B.n6 10.6151
R1295 B.n550 B.n549 10.6151
R1296 B.n551 B.n550 10.6151
R1297 B.n551 B.n4 10.6151
R1298 B.n555 B.n4 10.6151
R1299 B.n556 B.n555 10.6151
R1300 B.n557 B.n556 10.6151
R1301 B.n557 B.n0 10.6151
R1302 B.n533 B.n532 10.6151
R1303 B.n532 B.n531 10.6151
R1304 B.n531 B.n12 10.6151
R1305 B.n527 B.n12 10.6151
R1306 B.n527 B.n526 10.6151
R1307 B.n526 B.n525 10.6151
R1308 B.n525 B.n14 10.6151
R1309 B.n521 B.n14 10.6151
R1310 B.n521 B.n520 10.6151
R1311 B.n520 B.n519 10.6151
R1312 B.n519 B.n16 10.6151
R1313 B.n515 B.n16 10.6151
R1314 B.n515 B.n514 10.6151
R1315 B.n514 B.n513 10.6151
R1316 B.n513 B.n18 10.6151
R1317 B.n509 B.n18 10.6151
R1318 B.n509 B.n508 10.6151
R1319 B.n508 B.n507 10.6151
R1320 B.n507 B.n20 10.6151
R1321 B.n503 B.n20 10.6151
R1322 B.n503 B.n502 10.6151
R1323 B.n502 B.n501 10.6151
R1324 B.n501 B.n22 10.6151
R1325 B.n497 B.n22 10.6151
R1326 B.n497 B.n496 10.6151
R1327 B.n496 B.n495 10.6151
R1328 B.n495 B.n24 10.6151
R1329 B.n491 B.n24 10.6151
R1330 B.n491 B.n490 10.6151
R1331 B.n490 B.n489 10.6151
R1332 B.n489 B.n26 10.6151
R1333 B.n485 B.n26 10.6151
R1334 B.n485 B.n484 10.6151
R1335 B.n484 B.n483 10.6151
R1336 B.n483 B.n28 10.6151
R1337 B.n479 B.n28 10.6151
R1338 B.n479 B.n478 10.6151
R1339 B.n478 B.n477 10.6151
R1340 B.n477 B.n30 10.6151
R1341 B.n473 B.n30 10.6151
R1342 B.n473 B.n472 10.6151
R1343 B.n472 B.n471 10.6151
R1344 B.n471 B.n32 10.6151
R1345 B.n467 B.n32 10.6151
R1346 B.n467 B.n466 10.6151
R1347 B.n464 B.n36 10.6151
R1348 B.n460 B.n36 10.6151
R1349 B.n460 B.n459 10.6151
R1350 B.n459 B.n458 10.6151
R1351 B.n458 B.n38 10.6151
R1352 B.n454 B.n38 10.6151
R1353 B.n454 B.n453 10.6151
R1354 B.n453 B.n452 10.6151
R1355 B.n452 B.n40 10.6151
R1356 B.n448 B.n447 10.6151
R1357 B.n447 B.n446 10.6151
R1358 B.n446 B.n45 10.6151
R1359 B.n442 B.n45 10.6151
R1360 B.n442 B.n441 10.6151
R1361 B.n441 B.n440 10.6151
R1362 B.n440 B.n47 10.6151
R1363 B.n436 B.n47 10.6151
R1364 B.n436 B.n435 10.6151
R1365 B.n435 B.n434 10.6151
R1366 B.n434 B.n49 10.6151
R1367 B.n430 B.n49 10.6151
R1368 B.n430 B.n429 10.6151
R1369 B.n429 B.n428 10.6151
R1370 B.n428 B.n51 10.6151
R1371 B.n424 B.n51 10.6151
R1372 B.n424 B.n423 10.6151
R1373 B.n423 B.n422 10.6151
R1374 B.n422 B.n53 10.6151
R1375 B.n418 B.n53 10.6151
R1376 B.n418 B.n417 10.6151
R1377 B.n417 B.n416 10.6151
R1378 B.n416 B.n55 10.6151
R1379 B.n412 B.n55 10.6151
R1380 B.n412 B.n411 10.6151
R1381 B.n411 B.n410 10.6151
R1382 B.n410 B.n57 10.6151
R1383 B.n406 B.n57 10.6151
R1384 B.n406 B.n405 10.6151
R1385 B.n405 B.n404 10.6151
R1386 B.n404 B.n59 10.6151
R1387 B.n400 B.n59 10.6151
R1388 B.n400 B.n399 10.6151
R1389 B.n399 B.n398 10.6151
R1390 B.n398 B.n61 10.6151
R1391 B.n394 B.n61 10.6151
R1392 B.n394 B.n393 10.6151
R1393 B.n393 B.n392 10.6151
R1394 B.n392 B.n63 10.6151
R1395 B.n388 B.n63 10.6151
R1396 B.n388 B.n387 10.6151
R1397 B.n387 B.n386 10.6151
R1398 B.n386 B.n65 10.6151
R1399 B.n382 B.n65 10.6151
R1400 B.n382 B.n381 10.6151
R1401 B.n380 B.n67 10.6151
R1402 B.n376 B.n67 10.6151
R1403 B.n376 B.n375 10.6151
R1404 B.n375 B.n374 10.6151
R1405 B.n374 B.n69 10.6151
R1406 B.n370 B.n69 10.6151
R1407 B.n370 B.n369 10.6151
R1408 B.n369 B.n368 10.6151
R1409 B.n368 B.n71 10.6151
R1410 B.n364 B.n71 10.6151
R1411 B.n364 B.n363 10.6151
R1412 B.n363 B.n362 10.6151
R1413 B.n362 B.n73 10.6151
R1414 B.n358 B.n73 10.6151
R1415 B.n358 B.n357 10.6151
R1416 B.n357 B.n356 10.6151
R1417 B.n356 B.n75 10.6151
R1418 B.n352 B.n75 10.6151
R1419 B.n352 B.n351 10.6151
R1420 B.n351 B.n350 10.6151
R1421 B.n350 B.n77 10.6151
R1422 B.n346 B.n77 10.6151
R1423 B.n346 B.n345 10.6151
R1424 B.n345 B.n344 10.6151
R1425 B.n344 B.n79 10.6151
R1426 B.n340 B.n79 10.6151
R1427 B.n340 B.n339 10.6151
R1428 B.n339 B.n338 10.6151
R1429 B.n338 B.n81 10.6151
R1430 B.n334 B.n81 10.6151
R1431 B.n334 B.n333 10.6151
R1432 B.n333 B.n332 10.6151
R1433 B.n332 B.n83 10.6151
R1434 B.n328 B.n83 10.6151
R1435 B.n328 B.n327 10.6151
R1436 B.n145 B.n1 10.6151
R1437 B.n148 B.n145 10.6151
R1438 B.n149 B.n148 10.6151
R1439 B.n150 B.n149 10.6151
R1440 B.n150 B.n143 10.6151
R1441 B.n154 B.n143 10.6151
R1442 B.n155 B.n154 10.6151
R1443 B.n156 B.n155 10.6151
R1444 B.n156 B.n141 10.6151
R1445 B.n160 B.n141 10.6151
R1446 B.n161 B.n160 10.6151
R1447 B.n162 B.n161 10.6151
R1448 B.n162 B.n139 10.6151
R1449 B.n166 B.n139 10.6151
R1450 B.n167 B.n166 10.6151
R1451 B.n168 B.n167 10.6151
R1452 B.n172 B.n137 10.6151
R1453 B.n173 B.n172 10.6151
R1454 B.n174 B.n173 10.6151
R1455 B.n174 B.n135 10.6151
R1456 B.n178 B.n135 10.6151
R1457 B.n179 B.n178 10.6151
R1458 B.n180 B.n179 10.6151
R1459 B.n180 B.n133 10.6151
R1460 B.n184 B.n133 10.6151
R1461 B.n185 B.n184 10.6151
R1462 B.n186 B.n185 10.6151
R1463 B.n186 B.n131 10.6151
R1464 B.n190 B.n131 10.6151
R1465 B.n191 B.n190 10.6151
R1466 B.n192 B.n191 10.6151
R1467 B.n192 B.n129 10.6151
R1468 B.n196 B.n129 10.6151
R1469 B.n197 B.n196 10.6151
R1470 B.n198 B.n197 10.6151
R1471 B.n198 B.n127 10.6151
R1472 B.n202 B.n127 10.6151
R1473 B.n203 B.n202 10.6151
R1474 B.n204 B.n203 10.6151
R1475 B.n204 B.n125 10.6151
R1476 B.n208 B.n125 10.6151
R1477 B.n209 B.n208 10.6151
R1478 B.n210 B.n209 10.6151
R1479 B.n210 B.n123 10.6151
R1480 B.n214 B.n123 10.6151
R1481 B.n215 B.n214 10.6151
R1482 B.n216 B.n215 10.6151
R1483 B.n216 B.n121 10.6151
R1484 B.n220 B.n121 10.6151
R1485 B.n221 B.n220 10.6151
R1486 B.n222 B.n221 10.6151
R1487 B.n222 B.n119 10.6151
R1488 B.n226 B.n119 10.6151
R1489 B.n227 B.n226 10.6151
R1490 B.n228 B.n227 10.6151
R1491 B.n228 B.n117 10.6151
R1492 B.n232 B.n117 10.6151
R1493 B.n233 B.n232 10.6151
R1494 B.n234 B.n233 10.6151
R1495 B.n234 B.n115 10.6151
R1496 B.n238 B.n115 10.6151
R1497 B.n241 B.n240 10.6151
R1498 B.n241 B.n111 10.6151
R1499 B.n245 B.n111 10.6151
R1500 B.n246 B.n245 10.6151
R1501 B.n247 B.n246 10.6151
R1502 B.n247 B.n109 10.6151
R1503 B.n251 B.n109 10.6151
R1504 B.n252 B.n251 10.6151
R1505 B.n256 B.n252 10.6151
R1506 B.n260 B.n107 10.6151
R1507 B.n261 B.n260 10.6151
R1508 B.n262 B.n261 10.6151
R1509 B.n262 B.n105 10.6151
R1510 B.n266 B.n105 10.6151
R1511 B.n267 B.n266 10.6151
R1512 B.n268 B.n267 10.6151
R1513 B.n268 B.n103 10.6151
R1514 B.n272 B.n103 10.6151
R1515 B.n273 B.n272 10.6151
R1516 B.n274 B.n273 10.6151
R1517 B.n274 B.n101 10.6151
R1518 B.n278 B.n101 10.6151
R1519 B.n279 B.n278 10.6151
R1520 B.n280 B.n279 10.6151
R1521 B.n280 B.n99 10.6151
R1522 B.n284 B.n99 10.6151
R1523 B.n285 B.n284 10.6151
R1524 B.n286 B.n285 10.6151
R1525 B.n286 B.n97 10.6151
R1526 B.n290 B.n97 10.6151
R1527 B.n291 B.n290 10.6151
R1528 B.n292 B.n291 10.6151
R1529 B.n292 B.n95 10.6151
R1530 B.n296 B.n95 10.6151
R1531 B.n297 B.n296 10.6151
R1532 B.n298 B.n297 10.6151
R1533 B.n298 B.n93 10.6151
R1534 B.n302 B.n93 10.6151
R1535 B.n303 B.n302 10.6151
R1536 B.n304 B.n303 10.6151
R1537 B.n304 B.n91 10.6151
R1538 B.n308 B.n91 10.6151
R1539 B.n309 B.n308 10.6151
R1540 B.n310 B.n309 10.6151
R1541 B.n310 B.n89 10.6151
R1542 B.n314 B.n89 10.6151
R1543 B.n315 B.n314 10.6151
R1544 B.n316 B.n315 10.6151
R1545 B.n316 B.n87 10.6151
R1546 B.n320 B.n87 10.6151
R1547 B.n321 B.n320 10.6151
R1548 B.n322 B.n321 10.6151
R1549 B.n322 B.n85 10.6151
R1550 B.n326 B.n85 10.6151
R1551 B.n466 B.n465 9.36635
R1552 B.n448 B.n44 9.36635
R1553 B.n239 B.n238 9.36635
R1554 B.n255 B.n107 9.36635
R1555 B.n561 B.n0 8.11757
R1556 B.n561 B.n1 8.11757
R1557 B.n465 B.n464 1.24928
R1558 B.n44 B.n40 1.24928
R1559 B.n240 B.n239 1.24928
R1560 B.n256 B.n255 1.24928
R1561 VP.n1 VP.t5 802.601
R1562 VP.n8 VP.t4 785.309
R1563 VP.n6 VP.t0 785.309
R1564 VP.n3 VP.t2 785.309
R1565 VP.n7 VP.t3 775.816
R1566 VP.n2 VP.t1 775.816
R1567 VP.n9 VP.n8 161.3
R1568 VP.n4 VP.n3 161.3
R1569 VP.n7 VP.n0 161.3
R1570 VP.n6 VP.n5 161.3
R1571 VP.n4 VP.n1 72.2473
R1572 VP.n5 VP.n4 41.5838
R1573 VP.n7 VP.n6 38.7066
R1574 VP.n8 VP.n7 38.7066
R1575 VP.n3 VP.n2 38.7066
R1576 VP.n2 VP.n1 17.2717
R1577 VP.n5 VP.n0 0.189894
R1578 VP.n9 VP.n0 0.189894
R1579 VP VP.n9 0.0516364
R1580 VDD1.n68 VDD1.n0 756.745
R1581 VDD1.n141 VDD1.n73 756.745
R1582 VDD1.n69 VDD1.n68 585
R1583 VDD1.n67 VDD1.n66 585
R1584 VDD1.n4 VDD1.n3 585
R1585 VDD1.n61 VDD1.n60 585
R1586 VDD1.n59 VDD1.n58 585
R1587 VDD1.n8 VDD1.n7 585
R1588 VDD1.n53 VDD1.n52 585
R1589 VDD1.n51 VDD1.n50 585
R1590 VDD1.n12 VDD1.n11 585
R1591 VDD1.n16 VDD1.n14 585
R1592 VDD1.n45 VDD1.n44 585
R1593 VDD1.n43 VDD1.n42 585
R1594 VDD1.n18 VDD1.n17 585
R1595 VDD1.n37 VDD1.n36 585
R1596 VDD1.n35 VDD1.n34 585
R1597 VDD1.n22 VDD1.n21 585
R1598 VDD1.n29 VDD1.n28 585
R1599 VDD1.n27 VDD1.n26 585
R1600 VDD1.n98 VDD1.n97 585
R1601 VDD1.n100 VDD1.n99 585
R1602 VDD1.n93 VDD1.n92 585
R1603 VDD1.n106 VDD1.n105 585
R1604 VDD1.n108 VDD1.n107 585
R1605 VDD1.n89 VDD1.n88 585
R1606 VDD1.n115 VDD1.n114 585
R1607 VDD1.n116 VDD1.n87 585
R1608 VDD1.n118 VDD1.n117 585
R1609 VDD1.n85 VDD1.n84 585
R1610 VDD1.n124 VDD1.n123 585
R1611 VDD1.n126 VDD1.n125 585
R1612 VDD1.n81 VDD1.n80 585
R1613 VDD1.n132 VDD1.n131 585
R1614 VDD1.n134 VDD1.n133 585
R1615 VDD1.n77 VDD1.n76 585
R1616 VDD1.n140 VDD1.n139 585
R1617 VDD1.n142 VDD1.n141 585
R1618 VDD1.n25 VDD1.t0 329.036
R1619 VDD1.n96 VDD1.t5 329.036
R1620 VDD1.n68 VDD1.n67 171.744
R1621 VDD1.n67 VDD1.n3 171.744
R1622 VDD1.n60 VDD1.n3 171.744
R1623 VDD1.n60 VDD1.n59 171.744
R1624 VDD1.n59 VDD1.n7 171.744
R1625 VDD1.n52 VDD1.n7 171.744
R1626 VDD1.n52 VDD1.n51 171.744
R1627 VDD1.n51 VDD1.n11 171.744
R1628 VDD1.n16 VDD1.n11 171.744
R1629 VDD1.n44 VDD1.n16 171.744
R1630 VDD1.n44 VDD1.n43 171.744
R1631 VDD1.n43 VDD1.n17 171.744
R1632 VDD1.n36 VDD1.n17 171.744
R1633 VDD1.n36 VDD1.n35 171.744
R1634 VDD1.n35 VDD1.n21 171.744
R1635 VDD1.n28 VDD1.n21 171.744
R1636 VDD1.n28 VDD1.n27 171.744
R1637 VDD1.n99 VDD1.n98 171.744
R1638 VDD1.n99 VDD1.n92 171.744
R1639 VDD1.n106 VDD1.n92 171.744
R1640 VDD1.n107 VDD1.n106 171.744
R1641 VDD1.n107 VDD1.n88 171.744
R1642 VDD1.n115 VDD1.n88 171.744
R1643 VDD1.n116 VDD1.n115 171.744
R1644 VDD1.n117 VDD1.n116 171.744
R1645 VDD1.n117 VDD1.n84 171.744
R1646 VDD1.n124 VDD1.n84 171.744
R1647 VDD1.n125 VDD1.n124 171.744
R1648 VDD1.n125 VDD1.n80 171.744
R1649 VDD1.n132 VDD1.n80 171.744
R1650 VDD1.n133 VDD1.n132 171.744
R1651 VDD1.n133 VDD1.n76 171.744
R1652 VDD1.n140 VDD1.n76 171.744
R1653 VDD1.n141 VDD1.n140 171.744
R1654 VDD1.n27 VDD1.t0 85.8723
R1655 VDD1.n98 VDD1.t5 85.8723
R1656 VDD1.n147 VDD1.n146 71.2341
R1657 VDD1.n149 VDD1.n148 71.1171
R1658 VDD1 VDD1.n72 48.2759
R1659 VDD1.n147 VDD1.n145 48.1624
R1660 VDD1.n149 VDD1.n147 38.5224
R1661 VDD1.n14 VDD1.n12 13.1884
R1662 VDD1.n118 VDD1.n85 13.1884
R1663 VDD1.n50 VDD1.n49 12.8005
R1664 VDD1.n46 VDD1.n45 12.8005
R1665 VDD1.n119 VDD1.n87 12.8005
R1666 VDD1.n123 VDD1.n122 12.8005
R1667 VDD1.n53 VDD1.n10 12.0247
R1668 VDD1.n42 VDD1.n15 12.0247
R1669 VDD1.n114 VDD1.n113 12.0247
R1670 VDD1.n126 VDD1.n83 12.0247
R1671 VDD1.n54 VDD1.n8 11.249
R1672 VDD1.n41 VDD1.n18 11.249
R1673 VDD1.n112 VDD1.n89 11.249
R1674 VDD1.n127 VDD1.n81 11.249
R1675 VDD1.n26 VDD1.n25 10.7239
R1676 VDD1.n97 VDD1.n96 10.7239
R1677 VDD1.n58 VDD1.n57 10.4732
R1678 VDD1.n38 VDD1.n37 10.4732
R1679 VDD1.n109 VDD1.n108 10.4732
R1680 VDD1.n131 VDD1.n130 10.4732
R1681 VDD1.n61 VDD1.n6 9.69747
R1682 VDD1.n34 VDD1.n20 9.69747
R1683 VDD1.n105 VDD1.n91 9.69747
R1684 VDD1.n134 VDD1.n79 9.69747
R1685 VDD1.n72 VDD1.n71 9.45567
R1686 VDD1.n145 VDD1.n144 9.45567
R1687 VDD1.n24 VDD1.n23 9.3005
R1688 VDD1.n31 VDD1.n30 9.3005
R1689 VDD1.n33 VDD1.n32 9.3005
R1690 VDD1.n20 VDD1.n19 9.3005
R1691 VDD1.n39 VDD1.n38 9.3005
R1692 VDD1.n41 VDD1.n40 9.3005
R1693 VDD1.n15 VDD1.n13 9.3005
R1694 VDD1.n47 VDD1.n46 9.3005
R1695 VDD1.n71 VDD1.n70 9.3005
R1696 VDD1.n2 VDD1.n1 9.3005
R1697 VDD1.n65 VDD1.n64 9.3005
R1698 VDD1.n63 VDD1.n62 9.3005
R1699 VDD1.n6 VDD1.n5 9.3005
R1700 VDD1.n57 VDD1.n56 9.3005
R1701 VDD1.n55 VDD1.n54 9.3005
R1702 VDD1.n10 VDD1.n9 9.3005
R1703 VDD1.n49 VDD1.n48 9.3005
R1704 VDD1.n144 VDD1.n143 9.3005
R1705 VDD1.n138 VDD1.n137 9.3005
R1706 VDD1.n136 VDD1.n135 9.3005
R1707 VDD1.n79 VDD1.n78 9.3005
R1708 VDD1.n130 VDD1.n129 9.3005
R1709 VDD1.n128 VDD1.n127 9.3005
R1710 VDD1.n83 VDD1.n82 9.3005
R1711 VDD1.n122 VDD1.n121 9.3005
R1712 VDD1.n95 VDD1.n94 9.3005
R1713 VDD1.n102 VDD1.n101 9.3005
R1714 VDD1.n104 VDD1.n103 9.3005
R1715 VDD1.n91 VDD1.n90 9.3005
R1716 VDD1.n110 VDD1.n109 9.3005
R1717 VDD1.n112 VDD1.n111 9.3005
R1718 VDD1.n113 VDD1.n86 9.3005
R1719 VDD1.n120 VDD1.n119 9.3005
R1720 VDD1.n75 VDD1.n74 9.3005
R1721 VDD1.n62 VDD1.n4 8.92171
R1722 VDD1.n33 VDD1.n22 8.92171
R1723 VDD1.n104 VDD1.n93 8.92171
R1724 VDD1.n135 VDD1.n77 8.92171
R1725 VDD1.n66 VDD1.n65 8.14595
R1726 VDD1.n30 VDD1.n29 8.14595
R1727 VDD1.n101 VDD1.n100 8.14595
R1728 VDD1.n139 VDD1.n138 8.14595
R1729 VDD1.n72 VDD1.n0 7.3702
R1730 VDD1.n69 VDD1.n2 7.3702
R1731 VDD1.n26 VDD1.n24 7.3702
R1732 VDD1.n97 VDD1.n95 7.3702
R1733 VDD1.n142 VDD1.n75 7.3702
R1734 VDD1.n145 VDD1.n73 7.3702
R1735 VDD1.n70 VDD1.n0 6.59444
R1736 VDD1.n70 VDD1.n69 6.59444
R1737 VDD1.n143 VDD1.n142 6.59444
R1738 VDD1.n143 VDD1.n73 6.59444
R1739 VDD1.n66 VDD1.n2 5.81868
R1740 VDD1.n29 VDD1.n24 5.81868
R1741 VDD1.n100 VDD1.n95 5.81868
R1742 VDD1.n139 VDD1.n75 5.81868
R1743 VDD1.n65 VDD1.n4 5.04292
R1744 VDD1.n30 VDD1.n22 5.04292
R1745 VDD1.n101 VDD1.n93 5.04292
R1746 VDD1.n138 VDD1.n77 5.04292
R1747 VDD1.n62 VDD1.n61 4.26717
R1748 VDD1.n34 VDD1.n33 4.26717
R1749 VDD1.n105 VDD1.n104 4.26717
R1750 VDD1.n135 VDD1.n134 4.26717
R1751 VDD1.n58 VDD1.n6 3.49141
R1752 VDD1.n37 VDD1.n20 3.49141
R1753 VDD1.n108 VDD1.n91 3.49141
R1754 VDD1.n131 VDD1.n79 3.49141
R1755 VDD1.n57 VDD1.n8 2.71565
R1756 VDD1.n38 VDD1.n18 2.71565
R1757 VDD1.n109 VDD1.n89 2.71565
R1758 VDD1.n130 VDD1.n81 2.71565
R1759 VDD1.n25 VDD1.n23 2.41282
R1760 VDD1.n96 VDD1.n94 2.41282
R1761 VDD1.n148 VDD1.t4 2.40828
R1762 VDD1.n148 VDD1.t3 2.40828
R1763 VDD1.n146 VDD1.t2 2.40828
R1764 VDD1.n146 VDD1.t1 2.40828
R1765 VDD1.n54 VDD1.n53 1.93989
R1766 VDD1.n42 VDD1.n41 1.93989
R1767 VDD1.n114 VDD1.n112 1.93989
R1768 VDD1.n127 VDD1.n126 1.93989
R1769 VDD1.n50 VDD1.n10 1.16414
R1770 VDD1.n45 VDD1.n15 1.16414
R1771 VDD1.n113 VDD1.n87 1.16414
R1772 VDD1.n123 VDD1.n83 1.16414
R1773 VDD1.n49 VDD1.n12 0.388379
R1774 VDD1.n46 VDD1.n14 0.388379
R1775 VDD1.n119 VDD1.n118 0.388379
R1776 VDD1.n122 VDD1.n85 0.388379
R1777 VDD1.n71 VDD1.n1 0.155672
R1778 VDD1.n64 VDD1.n1 0.155672
R1779 VDD1.n64 VDD1.n63 0.155672
R1780 VDD1.n63 VDD1.n5 0.155672
R1781 VDD1.n56 VDD1.n5 0.155672
R1782 VDD1.n56 VDD1.n55 0.155672
R1783 VDD1.n55 VDD1.n9 0.155672
R1784 VDD1.n48 VDD1.n9 0.155672
R1785 VDD1.n48 VDD1.n47 0.155672
R1786 VDD1.n47 VDD1.n13 0.155672
R1787 VDD1.n40 VDD1.n13 0.155672
R1788 VDD1.n40 VDD1.n39 0.155672
R1789 VDD1.n39 VDD1.n19 0.155672
R1790 VDD1.n32 VDD1.n19 0.155672
R1791 VDD1.n32 VDD1.n31 0.155672
R1792 VDD1.n31 VDD1.n23 0.155672
R1793 VDD1.n102 VDD1.n94 0.155672
R1794 VDD1.n103 VDD1.n102 0.155672
R1795 VDD1.n103 VDD1.n90 0.155672
R1796 VDD1.n110 VDD1.n90 0.155672
R1797 VDD1.n111 VDD1.n110 0.155672
R1798 VDD1.n111 VDD1.n86 0.155672
R1799 VDD1.n120 VDD1.n86 0.155672
R1800 VDD1.n121 VDD1.n120 0.155672
R1801 VDD1.n121 VDD1.n82 0.155672
R1802 VDD1.n128 VDD1.n82 0.155672
R1803 VDD1.n129 VDD1.n128 0.155672
R1804 VDD1.n129 VDD1.n78 0.155672
R1805 VDD1.n136 VDD1.n78 0.155672
R1806 VDD1.n137 VDD1.n136 0.155672
R1807 VDD1.n137 VDD1.n74 0.155672
R1808 VDD1.n144 VDD1.n74 0.155672
R1809 VDD1 VDD1.n149 0.114724
C0 VN B 0.73386f
C1 VTAIL VDD1 12.8505f
C2 B w_n1610_n3668# 7.158121f
C3 VTAIL VDD2 12.8811f
C4 VP B 1.06075f
C5 VN w_n1610_n3668# 2.5508f
C6 VP VN 5.12849f
C7 B VDD1 1.59442f
C8 VP w_n1610_n3668# 2.75302f
C9 B VDD2 1.61812f
C10 VN VDD1 0.148091f
C11 w_n1610_n3668# VDD1 1.8571f
C12 VN VDD2 3.91427f
C13 w_n1610_n3668# VDD2 1.87419f
C14 VP VDD1 4.03949f
C15 VTAIL B 2.80292f
C16 VP VDD2 0.278764f
C17 VN VTAIL 3.46397f
C18 VTAIL w_n1610_n3668# 3.19941f
C19 VDD1 VDD2 0.629077f
C20 VP VTAIL 3.47873f
C21 VDD2 VSUBS 1.377155f
C22 VDD1 VSUBS 1.114574f
C23 VTAIL VSUBS 0.706795f
C24 VN VSUBS 4.56483f
C25 VP VSUBS 1.360397f
C26 B VSUBS 2.643589f
C27 w_n1610_n3668# VSUBS 72.5466f
C28 VDD1.n0 VSUBS 0.027724f
C29 VDD1.n1 VSUBS 0.025133f
C30 VDD1.n2 VSUBS 0.013505f
C31 VDD1.n3 VSUBS 0.031922f
C32 VDD1.n4 VSUBS 0.0143f
C33 VDD1.n5 VSUBS 0.025133f
C34 VDD1.n6 VSUBS 0.013505f
C35 VDD1.n7 VSUBS 0.031922f
C36 VDD1.n8 VSUBS 0.0143f
C37 VDD1.n9 VSUBS 0.025133f
C38 VDD1.n10 VSUBS 0.013505f
C39 VDD1.n11 VSUBS 0.031922f
C40 VDD1.n12 VSUBS 0.013903f
C41 VDD1.n13 VSUBS 0.025133f
C42 VDD1.n14 VSUBS 0.013903f
C43 VDD1.n15 VSUBS 0.013505f
C44 VDD1.n16 VSUBS 0.031922f
C45 VDD1.n17 VSUBS 0.031922f
C46 VDD1.n18 VSUBS 0.0143f
C47 VDD1.n19 VSUBS 0.025133f
C48 VDD1.n20 VSUBS 0.013505f
C49 VDD1.n21 VSUBS 0.031922f
C50 VDD1.n22 VSUBS 0.0143f
C51 VDD1.n23 VSUBS 1.40005f
C52 VDD1.n24 VSUBS 0.013505f
C53 VDD1.t0 VSUBS 0.068912f
C54 VDD1.n25 VSUBS 0.21498f
C55 VDD1.n26 VSUBS 0.024013f
C56 VDD1.n27 VSUBS 0.023941f
C57 VDD1.n28 VSUBS 0.031922f
C58 VDD1.n29 VSUBS 0.0143f
C59 VDD1.n30 VSUBS 0.013505f
C60 VDD1.n31 VSUBS 0.025133f
C61 VDD1.n32 VSUBS 0.025133f
C62 VDD1.n33 VSUBS 0.013505f
C63 VDD1.n34 VSUBS 0.0143f
C64 VDD1.n35 VSUBS 0.031922f
C65 VDD1.n36 VSUBS 0.031922f
C66 VDD1.n37 VSUBS 0.0143f
C67 VDD1.n38 VSUBS 0.013505f
C68 VDD1.n39 VSUBS 0.025133f
C69 VDD1.n40 VSUBS 0.025133f
C70 VDD1.n41 VSUBS 0.013505f
C71 VDD1.n42 VSUBS 0.0143f
C72 VDD1.n43 VSUBS 0.031922f
C73 VDD1.n44 VSUBS 0.031922f
C74 VDD1.n45 VSUBS 0.0143f
C75 VDD1.n46 VSUBS 0.013505f
C76 VDD1.n47 VSUBS 0.025133f
C77 VDD1.n48 VSUBS 0.025133f
C78 VDD1.n49 VSUBS 0.013505f
C79 VDD1.n50 VSUBS 0.0143f
C80 VDD1.n51 VSUBS 0.031922f
C81 VDD1.n52 VSUBS 0.031922f
C82 VDD1.n53 VSUBS 0.0143f
C83 VDD1.n54 VSUBS 0.013505f
C84 VDD1.n55 VSUBS 0.025133f
C85 VDD1.n56 VSUBS 0.025133f
C86 VDD1.n57 VSUBS 0.013505f
C87 VDD1.n58 VSUBS 0.0143f
C88 VDD1.n59 VSUBS 0.031922f
C89 VDD1.n60 VSUBS 0.031922f
C90 VDD1.n61 VSUBS 0.0143f
C91 VDD1.n62 VSUBS 0.013505f
C92 VDD1.n63 VSUBS 0.025133f
C93 VDD1.n64 VSUBS 0.025133f
C94 VDD1.n65 VSUBS 0.013505f
C95 VDD1.n66 VSUBS 0.0143f
C96 VDD1.n67 VSUBS 0.031922f
C97 VDD1.n68 VSUBS 0.077647f
C98 VDD1.n69 VSUBS 0.0143f
C99 VDD1.n70 VSUBS 0.013505f
C100 VDD1.n71 VSUBS 0.056033f
C101 VDD1.n72 VSUBS 0.057489f
C102 VDD1.n73 VSUBS 0.027724f
C103 VDD1.n74 VSUBS 0.025133f
C104 VDD1.n75 VSUBS 0.013505f
C105 VDD1.n76 VSUBS 0.031922f
C106 VDD1.n77 VSUBS 0.0143f
C107 VDD1.n78 VSUBS 0.025133f
C108 VDD1.n79 VSUBS 0.013505f
C109 VDD1.n80 VSUBS 0.031922f
C110 VDD1.n81 VSUBS 0.0143f
C111 VDD1.n82 VSUBS 0.025133f
C112 VDD1.n83 VSUBS 0.013505f
C113 VDD1.n84 VSUBS 0.031922f
C114 VDD1.n85 VSUBS 0.013903f
C115 VDD1.n86 VSUBS 0.025133f
C116 VDD1.n87 VSUBS 0.0143f
C117 VDD1.n88 VSUBS 0.031922f
C118 VDD1.n89 VSUBS 0.0143f
C119 VDD1.n90 VSUBS 0.025133f
C120 VDD1.n91 VSUBS 0.013505f
C121 VDD1.n92 VSUBS 0.031922f
C122 VDD1.n93 VSUBS 0.0143f
C123 VDD1.n94 VSUBS 1.40005f
C124 VDD1.n95 VSUBS 0.013505f
C125 VDD1.t5 VSUBS 0.068912f
C126 VDD1.n96 VSUBS 0.21498f
C127 VDD1.n97 VSUBS 0.024013f
C128 VDD1.n98 VSUBS 0.023941f
C129 VDD1.n99 VSUBS 0.031922f
C130 VDD1.n100 VSUBS 0.0143f
C131 VDD1.n101 VSUBS 0.013505f
C132 VDD1.n102 VSUBS 0.025133f
C133 VDD1.n103 VSUBS 0.025133f
C134 VDD1.n104 VSUBS 0.013505f
C135 VDD1.n105 VSUBS 0.0143f
C136 VDD1.n106 VSUBS 0.031922f
C137 VDD1.n107 VSUBS 0.031922f
C138 VDD1.n108 VSUBS 0.0143f
C139 VDD1.n109 VSUBS 0.013505f
C140 VDD1.n110 VSUBS 0.025133f
C141 VDD1.n111 VSUBS 0.025133f
C142 VDD1.n112 VSUBS 0.013505f
C143 VDD1.n113 VSUBS 0.013505f
C144 VDD1.n114 VSUBS 0.0143f
C145 VDD1.n115 VSUBS 0.031922f
C146 VDD1.n116 VSUBS 0.031922f
C147 VDD1.n117 VSUBS 0.031922f
C148 VDD1.n118 VSUBS 0.013903f
C149 VDD1.n119 VSUBS 0.013505f
C150 VDD1.n120 VSUBS 0.025133f
C151 VDD1.n121 VSUBS 0.025133f
C152 VDD1.n122 VSUBS 0.013505f
C153 VDD1.n123 VSUBS 0.0143f
C154 VDD1.n124 VSUBS 0.031922f
C155 VDD1.n125 VSUBS 0.031922f
C156 VDD1.n126 VSUBS 0.0143f
C157 VDD1.n127 VSUBS 0.013505f
C158 VDD1.n128 VSUBS 0.025133f
C159 VDD1.n129 VSUBS 0.025133f
C160 VDD1.n130 VSUBS 0.013505f
C161 VDD1.n131 VSUBS 0.0143f
C162 VDD1.n132 VSUBS 0.031922f
C163 VDD1.n133 VSUBS 0.031922f
C164 VDD1.n134 VSUBS 0.0143f
C165 VDD1.n135 VSUBS 0.013505f
C166 VDD1.n136 VSUBS 0.025133f
C167 VDD1.n137 VSUBS 0.025133f
C168 VDD1.n138 VSUBS 0.013505f
C169 VDD1.n139 VSUBS 0.0143f
C170 VDD1.n140 VSUBS 0.031922f
C171 VDD1.n141 VSUBS 0.077647f
C172 VDD1.n142 VSUBS 0.0143f
C173 VDD1.n143 VSUBS 0.013505f
C174 VDD1.n144 VSUBS 0.056033f
C175 VDD1.n145 VSUBS 0.057194f
C176 VDD1.t2 VSUBS 0.26812f
C177 VDD1.t1 VSUBS 0.26812f
C178 VDD1.n146 VSUBS 2.12839f
C179 VDD1.n147 VSUBS 2.20472f
C180 VDD1.t4 VSUBS 0.26812f
C181 VDD1.t3 VSUBS 0.26812f
C182 VDD1.n148 VSUBS 2.12745f
C183 VDD1.n149 VSUBS 2.59786f
C184 VP.n0 VSUBS 0.064578f
C185 VP.t0 VSUBS 1.17161f
C186 VP.t5 VSUBS 1.18151f
C187 VP.n1 VSUBS 0.450093f
C188 VP.t1 VSUBS 1.16616f
C189 VP.n2 VSUBS 0.470313f
C190 VP.t2 VSUBS 1.17161f
C191 VP.n3 VSUBS 0.459494f
C192 VP.n4 VSUBS 2.77282f
C193 VP.n5 VSUBS 2.67746f
C194 VP.n6 VSUBS 0.459494f
C195 VP.t3 VSUBS 1.16616f
C196 VP.n7 VSUBS 0.470313f
C197 VP.t4 VSUBS 1.17161f
C198 VP.n8 VSUBS 0.459494f
C199 VP.n9 VSUBS 0.050045f
C200 B.n0 VSUBS 0.006559f
C201 B.n1 VSUBS 0.006559f
C202 B.n2 VSUBS 0.009701f
C203 B.n3 VSUBS 0.007434f
C204 B.n4 VSUBS 0.007434f
C205 B.n5 VSUBS 0.007434f
C206 B.n6 VSUBS 0.007434f
C207 B.n7 VSUBS 0.007434f
C208 B.n8 VSUBS 0.007434f
C209 B.n9 VSUBS 0.007434f
C210 B.n10 VSUBS 0.016123f
C211 B.n11 VSUBS 0.007434f
C212 B.n12 VSUBS 0.007434f
C213 B.n13 VSUBS 0.007434f
C214 B.n14 VSUBS 0.007434f
C215 B.n15 VSUBS 0.007434f
C216 B.n16 VSUBS 0.007434f
C217 B.n17 VSUBS 0.007434f
C218 B.n18 VSUBS 0.007434f
C219 B.n19 VSUBS 0.007434f
C220 B.n20 VSUBS 0.007434f
C221 B.n21 VSUBS 0.007434f
C222 B.n22 VSUBS 0.007434f
C223 B.n23 VSUBS 0.007434f
C224 B.n24 VSUBS 0.007434f
C225 B.n25 VSUBS 0.007434f
C226 B.n26 VSUBS 0.007434f
C227 B.n27 VSUBS 0.007434f
C228 B.n28 VSUBS 0.007434f
C229 B.n29 VSUBS 0.007434f
C230 B.n30 VSUBS 0.007434f
C231 B.n31 VSUBS 0.007434f
C232 B.n32 VSUBS 0.007434f
C233 B.n33 VSUBS 0.007434f
C234 B.t1 VSUBS 0.260182f
C235 B.t2 VSUBS 0.270159f
C236 B.t0 VSUBS 0.269363f
C237 B.n34 VSUBS 0.340844f
C238 B.n35 VSUBS 0.279582f
C239 B.n36 VSUBS 0.007434f
C240 B.n37 VSUBS 0.007434f
C241 B.n38 VSUBS 0.007434f
C242 B.n39 VSUBS 0.007434f
C243 B.n40 VSUBS 0.004154f
C244 B.n41 VSUBS 0.007434f
C245 B.t4 VSUBS 0.260185f
C246 B.t5 VSUBS 0.270163f
C247 B.t3 VSUBS 0.269363f
C248 B.n42 VSUBS 0.340841f
C249 B.n43 VSUBS 0.279579f
C250 B.n44 VSUBS 0.017223f
C251 B.n45 VSUBS 0.007434f
C252 B.n46 VSUBS 0.007434f
C253 B.n47 VSUBS 0.007434f
C254 B.n48 VSUBS 0.007434f
C255 B.n49 VSUBS 0.007434f
C256 B.n50 VSUBS 0.007434f
C257 B.n51 VSUBS 0.007434f
C258 B.n52 VSUBS 0.007434f
C259 B.n53 VSUBS 0.007434f
C260 B.n54 VSUBS 0.007434f
C261 B.n55 VSUBS 0.007434f
C262 B.n56 VSUBS 0.007434f
C263 B.n57 VSUBS 0.007434f
C264 B.n58 VSUBS 0.007434f
C265 B.n59 VSUBS 0.007434f
C266 B.n60 VSUBS 0.007434f
C267 B.n61 VSUBS 0.007434f
C268 B.n62 VSUBS 0.007434f
C269 B.n63 VSUBS 0.007434f
C270 B.n64 VSUBS 0.007434f
C271 B.n65 VSUBS 0.007434f
C272 B.n66 VSUBS 0.017329f
C273 B.n67 VSUBS 0.007434f
C274 B.n68 VSUBS 0.007434f
C275 B.n69 VSUBS 0.007434f
C276 B.n70 VSUBS 0.007434f
C277 B.n71 VSUBS 0.007434f
C278 B.n72 VSUBS 0.007434f
C279 B.n73 VSUBS 0.007434f
C280 B.n74 VSUBS 0.007434f
C281 B.n75 VSUBS 0.007434f
C282 B.n76 VSUBS 0.007434f
C283 B.n77 VSUBS 0.007434f
C284 B.n78 VSUBS 0.007434f
C285 B.n79 VSUBS 0.007434f
C286 B.n80 VSUBS 0.007434f
C287 B.n81 VSUBS 0.007434f
C288 B.n82 VSUBS 0.007434f
C289 B.n83 VSUBS 0.007434f
C290 B.n84 VSUBS 0.016123f
C291 B.n85 VSUBS 0.007434f
C292 B.n86 VSUBS 0.007434f
C293 B.n87 VSUBS 0.007434f
C294 B.n88 VSUBS 0.007434f
C295 B.n89 VSUBS 0.007434f
C296 B.n90 VSUBS 0.007434f
C297 B.n91 VSUBS 0.007434f
C298 B.n92 VSUBS 0.007434f
C299 B.n93 VSUBS 0.007434f
C300 B.n94 VSUBS 0.007434f
C301 B.n95 VSUBS 0.007434f
C302 B.n96 VSUBS 0.007434f
C303 B.n97 VSUBS 0.007434f
C304 B.n98 VSUBS 0.007434f
C305 B.n99 VSUBS 0.007434f
C306 B.n100 VSUBS 0.007434f
C307 B.n101 VSUBS 0.007434f
C308 B.n102 VSUBS 0.007434f
C309 B.n103 VSUBS 0.007434f
C310 B.n104 VSUBS 0.007434f
C311 B.n105 VSUBS 0.007434f
C312 B.n106 VSUBS 0.007434f
C313 B.n107 VSUBS 0.006997f
C314 B.n108 VSUBS 0.007434f
C315 B.n109 VSUBS 0.007434f
C316 B.n110 VSUBS 0.007434f
C317 B.n111 VSUBS 0.007434f
C318 B.n112 VSUBS 0.007434f
C319 B.t8 VSUBS 0.260182f
C320 B.t7 VSUBS 0.270159f
C321 B.t6 VSUBS 0.269363f
C322 B.n113 VSUBS 0.340844f
C323 B.n114 VSUBS 0.279582f
C324 B.n115 VSUBS 0.007434f
C325 B.n116 VSUBS 0.007434f
C326 B.n117 VSUBS 0.007434f
C327 B.n118 VSUBS 0.007434f
C328 B.n119 VSUBS 0.007434f
C329 B.n120 VSUBS 0.007434f
C330 B.n121 VSUBS 0.007434f
C331 B.n122 VSUBS 0.007434f
C332 B.n123 VSUBS 0.007434f
C333 B.n124 VSUBS 0.007434f
C334 B.n125 VSUBS 0.007434f
C335 B.n126 VSUBS 0.007434f
C336 B.n127 VSUBS 0.007434f
C337 B.n128 VSUBS 0.007434f
C338 B.n129 VSUBS 0.007434f
C339 B.n130 VSUBS 0.007434f
C340 B.n131 VSUBS 0.007434f
C341 B.n132 VSUBS 0.007434f
C342 B.n133 VSUBS 0.007434f
C343 B.n134 VSUBS 0.007434f
C344 B.n135 VSUBS 0.007434f
C345 B.n136 VSUBS 0.007434f
C346 B.n137 VSUBS 0.017329f
C347 B.n138 VSUBS 0.007434f
C348 B.n139 VSUBS 0.007434f
C349 B.n140 VSUBS 0.007434f
C350 B.n141 VSUBS 0.007434f
C351 B.n142 VSUBS 0.007434f
C352 B.n143 VSUBS 0.007434f
C353 B.n144 VSUBS 0.007434f
C354 B.n145 VSUBS 0.007434f
C355 B.n146 VSUBS 0.007434f
C356 B.n147 VSUBS 0.007434f
C357 B.n148 VSUBS 0.007434f
C358 B.n149 VSUBS 0.007434f
C359 B.n150 VSUBS 0.007434f
C360 B.n151 VSUBS 0.007434f
C361 B.n152 VSUBS 0.007434f
C362 B.n153 VSUBS 0.007434f
C363 B.n154 VSUBS 0.007434f
C364 B.n155 VSUBS 0.007434f
C365 B.n156 VSUBS 0.007434f
C366 B.n157 VSUBS 0.007434f
C367 B.n158 VSUBS 0.007434f
C368 B.n159 VSUBS 0.007434f
C369 B.n160 VSUBS 0.007434f
C370 B.n161 VSUBS 0.007434f
C371 B.n162 VSUBS 0.007434f
C372 B.n163 VSUBS 0.007434f
C373 B.n164 VSUBS 0.007434f
C374 B.n165 VSUBS 0.007434f
C375 B.n166 VSUBS 0.007434f
C376 B.n167 VSUBS 0.007434f
C377 B.n168 VSUBS 0.016123f
C378 B.n169 VSUBS 0.016123f
C379 B.n170 VSUBS 0.017329f
C380 B.n171 VSUBS 0.007434f
C381 B.n172 VSUBS 0.007434f
C382 B.n173 VSUBS 0.007434f
C383 B.n174 VSUBS 0.007434f
C384 B.n175 VSUBS 0.007434f
C385 B.n176 VSUBS 0.007434f
C386 B.n177 VSUBS 0.007434f
C387 B.n178 VSUBS 0.007434f
C388 B.n179 VSUBS 0.007434f
C389 B.n180 VSUBS 0.007434f
C390 B.n181 VSUBS 0.007434f
C391 B.n182 VSUBS 0.007434f
C392 B.n183 VSUBS 0.007434f
C393 B.n184 VSUBS 0.007434f
C394 B.n185 VSUBS 0.007434f
C395 B.n186 VSUBS 0.007434f
C396 B.n187 VSUBS 0.007434f
C397 B.n188 VSUBS 0.007434f
C398 B.n189 VSUBS 0.007434f
C399 B.n190 VSUBS 0.007434f
C400 B.n191 VSUBS 0.007434f
C401 B.n192 VSUBS 0.007434f
C402 B.n193 VSUBS 0.007434f
C403 B.n194 VSUBS 0.007434f
C404 B.n195 VSUBS 0.007434f
C405 B.n196 VSUBS 0.007434f
C406 B.n197 VSUBS 0.007434f
C407 B.n198 VSUBS 0.007434f
C408 B.n199 VSUBS 0.007434f
C409 B.n200 VSUBS 0.007434f
C410 B.n201 VSUBS 0.007434f
C411 B.n202 VSUBS 0.007434f
C412 B.n203 VSUBS 0.007434f
C413 B.n204 VSUBS 0.007434f
C414 B.n205 VSUBS 0.007434f
C415 B.n206 VSUBS 0.007434f
C416 B.n207 VSUBS 0.007434f
C417 B.n208 VSUBS 0.007434f
C418 B.n209 VSUBS 0.007434f
C419 B.n210 VSUBS 0.007434f
C420 B.n211 VSUBS 0.007434f
C421 B.n212 VSUBS 0.007434f
C422 B.n213 VSUBS 0.007434f
C423 B.n214 VSUBS 0.007434f
C424 B.n215 VSUBS 0.007434f
C425 B.n216 VSUBS 0.007434f
C426 B.n217 VSUBS 0.007434f
C427 B.n218 VSUBS 0.007434f
C428 B.n219 VSUBS 0.007434f
C429 B.n220 VSUBS 0.007434f
C430 B.n221 VSUBS 0.007434f
C431 B.n222 VSUBS 0.007434f
C432 B.n223 VSUBS 0.007434f
C433 B.n224 VSUBS 0.007434f
C434 B.n225 VSUBS 0.007434f
C435 B.n226 VSUBS 0.007434f
C436 B.n227 VSUBS 0.007434f
C437 B.n228 VSUBS 0.007434f
C438 B.n229 VSUBS 0.007434f
C439 B.n230 VSUBS 0.007434f
C440 B.n231 VSUBS 0.007434f
C441 B.n232 VSUBS 0.007434f
C442 B.n233 VSUBS 0.007434f
C443 B.n234 VSUBS 0.007434f
C444 B.n235 VSUBS 0.007434f
C445 B.n236 VSUBS 0.007434f
C446 B.n237 VSUBS 0.007434f
C447 B.n238 VSUBS 0.006997f
C448 B.n239 VSUBS 0.017223f
C449 B.n240 VSUBS 0.004154f
C450 B.n241 VSUBS 0.007434f
C451 B.n242 VSUBS 0.007434f
C452 B.n243 VSUBS 0.007434f
C453 B.n244 VSUBS 0.007434f
C454 B.n245 VSUBS 0.007434f
C455 B.n246 VSUBS 0.007434f
C456 B.n247 VSUBS 0.007434f
C457 B.n248 VSUBS 0.007434f
C458 B.n249 VSUBS 0.007434f
C459 B.n250 VSUBS 0.007434f
C460 B.n251 VSUBS 0.007434f
C461 B.n252 VSUBS 0.007434f
C462 B.t11 VSUBS 0.260185f
C463 B.t10 VSUBS 0.270163f
C464 B.t9 VSUBS 0.269363f
C465 B.n253 VSUBS 0.340841f
C466 B.n254 VSUBS 0.279579f
C467 B.n255 VSUBS 0.017223f
C468 B.n256 VSUBS 0.004154f
C469 B.n257 VSUBS 0.007434f
C470 B.n258 VSUBS 0.007434f
C471 B.n259 VSUBS 0.007434f
C472 B.n260 VSUBS 0.007434f
C473 B.n261 VSUBS 0.007434f
C474 B.n262 VSUBS 0.007434f
C475 B.n263 VSUBS 0.007434f
C476 B.n264 VSUBS 0.007434f
C477 B.n265 VSUBS 0.007434f
C478 B.n266 VSUBS 0.007434f
C479 B.n267 VSUBS 0.007434f
C480 B.n268 VSUBS 0.007434f
C481 B.n269 VSUBS 0.007434f
C482 B.n270 VSUBS 0.007434f
C483 B.n271 VSUBS 0.007434f
C484 B.n272 VSUBS 0.007434f
C485 B.n273 VSUBS 0.007434f
C486 B.n274 VSUBS 0.007434f
C487 B.n275 VSUBS 0.007434f
C488 B.n276 VSUBS 0.007434f
C489 B.n277 VSUBS 0.007434f
C490 B.n278 VSUBS 0.007434f
C491 B.n279 VSUBS 0.007434f
C492 B.n280 VSUBS 0.007434f
C493 B.n281 VSUBS 0.007434f
C494 B.n282 VSUBS 0.007434f
C495 B.n283 VSUBS 0.007434f
C496 B.n284 VSUBS 0.007434f
C497 B.n285 VSUBS 0.007434f
C498 B.n286 VSUBS 0.007434f
C499 B.n287 VSUBS 0.007434f
C500 B.n288 VSUBS 0.007434f
C501 B.n289 VSUBS 0.007434f
C502 B.n290 VSUBS 0.007434f
C503 B.n291 VSUBS 0.007434f
C504 B.n292 VSUBS 0.007434f
C505 B.n293 VSUBS 0.007434f
C506 B.n294 VSUBS 0.007434f
C507 B.n295 VSUBS 0.007434f
C508 B.n296 VSUBS 0.007434f
C509 B.n297 VSUBS 0.007434f
C510 B.n298 VSUBS 0.007434f
C511 B.n299 VSUBS 0.007434f
C512 B.n300 VSUBS 0.007434f
C513 B.n301 VSUBS 0.007434f
C514 B.n302 VSUBS 0.007434f
C515 B.n303 VSUBS 0.007434f
C516 B.n304 VSUBS 0.007434f
C517 B.n305 VSUBS 0.007434f
C518 B.n306 VSUBS 0.007434f
C519 B.n307 VSUBS 0.007434f
C520 B.n308 VSUBS 0.007434f
C521 B.n309 VSUBS 0.007434f
C522 B.n310 VSUBS 0.007434f
C523 B.n311 VSUBS 0.007434f
C524 B.n312 VSUBS 0.007434f
C525 B.n313 VSUBS 0.007434f
C526 B.n314 VSUBS 0.007434f
C527 B.n315 VSUBS 0.007434f
C528 B.n316 VSUBS 0.007434f
C529 B.n317 VSUBS 0.007434f
C530 B.n318 VSUBS 0.007434f
C531 B.n319 VSUBS 0.007434f
C532 B.n320 VSUBS 0.007434f
C533 B.n321 VSUBS 0.007434f
C534 B.n322 VSUBS 0.007434f
C535 B.n323 VSUBS 0.007434f
C536 B.n324 VSUBS 0.007434f
C537 B.n325 VSUBS 0.017329f
C538 B.n326 VSUBS 0.016396f
C539 B.n327 VSUBS 0.017056f
C540 B.n328 VSUBS 0.007434f
C541 B.n329 VSUBS 0.007434f
C542 B.n330 VSUBS 0.007434f
C543 B.n331 VSUBS 0.007434f
C544 B.n332 VSUBS 0.007434f
C545 B.n333 VSUBS 0.007434f
C546 B.n334 VSUBS 0.007434f
C547 B.n335 VSUBS 0.007434f
C548 B.n336 VSUBS 0.007434f
C549 B.n337 VSUBS 0.007434f
C550 B.n338 VSUBS 0.007434f
C551 B.n339 VSUBS 0.007434f
C552 B.n340 VSUBS 0.007434f
C553 B.n341 VSUBS 0.007434f
C554 B.n342 VSUBS 0.007434f
C555 B.n343 VSUBS 0.007434f
C556 B.n344 VSUBS 0.007434f
C557 B.n345 VSUBS 0.007434f
C558 B.n346 VSUBS 0.007434f
C559 B.n347 VSUBS 0.007434f
C560 B.n348 VSUBS 0.007434f
C561 B.n349 VSUBS 0.007434f
C562 B.n350 VSUBS 0.007434f
C563 B.n351 VSUBS 0.007434f
C564 B.n352 VSUBS 0.007434f
C565 B.n353 VSUBS 0.007434f
C566 B.n354 VSUBS 0.007434f
C567 B.n355 VSUBS 0.007434f
C568 B.n356 VSUBS 0.007434f
C569 B.n357 VSUBS 0.007434f
C570 B.n358 VSUBS 0.007434f
C571 B.n359 VSUBS 0.007434f
C572 B.n360 VSUBS 0.007434f
C573 B.n361 VSUBS 0.007434f
C574 B.n362 VSUBS 0.007434f
C575 B.n363 VSUBS 0.007434f
C576 B.n364 VSUBS 0.007434f
C577 B.n365 VSUBS 0.007434f
C578 B.n366 VSUBS 0.007434f
C579 B.n367 VSUBS 0.007434f
C580 B.n368 VSUBS 0.007434f
C581 B.n369 VSUBS 0.007434f
C582 B.n370 VSUBS 0.007434f
C583 B.n371 VSUBS 0.007434f
C584 B.n372 VSUBS 0.007434f
C585 B.n373 VSUBS 0.007434f
C586 B.n374 VSUBS 0.007434f
C587 B.n375 VSUBS 0.007434f
C588 B.n376 VSUBS 0.007434f
C589 B.n377 VSUBS 0.007434f
C590 B.n378 VSUBS 0.007434f
C591 B.n379 VSUBS 0.016123f
C592 B.n380 VSUBS 0.016123f
C593 B.n381 VSUBS 0.017329f
C594 B.n382 VSUBS 0.007434f
C595 B.n383 VSUBS 0.007434f
C596 B.n384 VSUBS 0.007434f
C597 B.n385 VSUBS 0.007434f
C598 B.n386 VSUBS 0.007434f
C599 B.n387 VSUBS 0.007434f
C600 B.n388 VSUBS 0.007434f
C601 B.n389 VSUBS 0.007434f
C602 B.n390 VSUBS 0.007434f
C603 B.n391 VSUBS 0.007434f
C604 B.n392 VSUBS 0.007434f
C605 B.n393 VSUBS 0.007434f
C606 B.n394 VSUBS 0.007434f
C607 B.n395 VSUBS 0.007434f
C608 B.n396 VSUBS 0.007434f
C609 B.n397 VSUBS 0.007434f
C610 B.n398 VSUBS 0.007434f
C611 B.n399 VSUBS 0.007434f
C612 B.n400 VSUBS 0.007434f
C613 B.n401 VSUBS 0.007434f
C614 B.n402 VSUBS 0.007434f
C615 B.n403 VSUBS 0.007434f
C616 B.n404 VSUBS 0.007434f
C617 B.n405 VSUBS 0.007434f
C618 B.n406 VSUBS 0.007434f
C619 B.n407 VSUBS 0.007434f
C620 B.n408 VSUBS 0.007434f
C621 B.n409 VSUBS 0.007434f
C622 B.n410 VSUBS 0.007434f
C623 B.n411 VSUBS 0.007434f
C624 B.n412 VSUBS 0.007434f
C625 B.n413 VSUBS 0.007434f
C626 B.n414 VSUBS 0.007434f
C627 B.n415 VSUBS 0.007434f
C628 B.n416 VSUBS 0.007434f
C629 B.n417 VSUBS 0.007434f
C630 B.n418 VSUBS 0.007434f
C631 B.n419 VSUBS 0.007434f
C632 B.n420 VSUBS 0.007434f
C633 B.n421 VSUBS 0.007434f
C634 B.n422 VSUBS 0.007434f
C635 B.n423 VSUBS 0.007434f
C636 B.n424 VSUBS 0.007434f
C637 B.n425 VSUBS 0.007434f
C638 B.n426 VSUBS 0.007434f
C639 B.n427 VSUBS 0.007434f
C640 B.n428 VSUBS 0.007434f
C641 B.n429 VSUBS 0.007434f
C642 B.n430 VSUBS 0.007434f
C643 B.n431 VSUBS 0.007434f
C644 B.n432 VSUBS 0.007434f
C645 B.n433 VSUBS 0.007434f
C646 B.n434 VSUBS 0.007434f
C647 B.n435 VSUBS 0.007434f
C648 B.n436 VSUBS 0.007434f
C649 B.n437 VSUBS 0.007434f
C650 B.n438 VSUBS 0.007434f
C651 B.n439 VSUBS 0.007434f
C652 B.n440 VSUBS 0.007434f
C653 B.n441 VSUBS 0.007434f
C654 B.n442 VSUBS 0.007434f
C655 B.n443 VSUBS 0.007434f
C656 B.n444 VSUBS 0.007434f
C657 B.n445 VSUBS 0.007434f
C658 B.n446 VSUBS 0.007434f
C659 B.n447 VSUBS 0.007434f
C660 B.n448 VSUBS 0.006997f
C661 B.n449 VSUBS 0.007434f
C662 B.n450 VSUBS 0.007434f
C663 B.n451 VSUBS 0.007434f
C664 B.n452 VSUBS 0.007434f
C665 B.n453 VSUBS 0.007434f
C666 B.n454 VSUBS 0.007434f
C667 B.n455 VSUBS 0.007434f
C668 B.n456 VSUBS 0.007434f
C669 B.n457 VSUBS 0.007434f
C670 B.n458 VSUBS 0.007434f
C671 B.n459 VSUBS 0.007434f
C672 B.n460 VSUBS 0.007434f
C673 B.n461 VSUBS 0.007434f
C674 B.n462 VSUBS 0.007434f
C675 B.n463 VSUBS 0.007434f
C676 B.n464 VSUBS 0.004154f
C677 B.n465 VSUBS 0.017223f
C678 B.n466 VSUBS 0.006997f
C679 B.n467 VSUBS 0.007434f
C680 B.n468 VSUBS 0.007434f
C681 B.n469 VSUBS 0.007434f
C682 B.n470 VSUBS 0.007434f
C683 B.n471 VSUBS 0.007434f
C684 B.n472 VSUBS 0.007434f
C685 B.n473 VSUBS 0.007434f
C686 B.n474 VSUBS 0.007434f
C687 B.n475 VSUBS 0.007434f
C688 B.n476 VSUBS 0.007434f
C689 B.n477 VSUBS 0.007434f
C690 B.n478 VSUBS 0.007434f
C691 B.n479 VSUBS 0.007434f
C692 B.n480 VSUBS 0.007434f
C693 B.n481 VSUBS 0.007434f
C694 B.n482 VSUBS 0.007434f
C695 B.n483 VSUBS 0.007434f
C696 B.n484 VSUBS 0.007434f
C697 B.n485 VSUBS 0.007434f
C698 B.n486 VSUBS 0.007434f
C699 B.n487 VSUBS 0.007434f
C700 B.n488 VSUBS 0.007434f
C701 B.n489 VSUBS 0.007434f
C702 B.n490 VSUBS 0.007434f
C703 B.n491 VSUBS 0.007434f
C704 B.n492 VSUBS 0.007434f
C705 B.n493 VSUBS 0.007434f
C706 B.n494 VSUBS 0.007434f
C707 B.n495 VSUBS 0.007434f
C708 B.n496 VSUBS 0.007434f
C709 B.n497 VSUBS 0.007434f
C710 B.n498 VSUBS 0.007434f
C711 B.n499 VSUBS 0.007434f
C712 B.n500 VSUBS 0.007434f
C713 B.n501 VSUBS 0.007434f
C714 B.n502 VSUBS 0.007434f
C715 B.n503 VSUBS 0.007434f
C716 B.n504 VSUBS 0.007434f
C717 B.n505 VSUBS 0.007434f
C718 B.n506 VSUBS 0.007434f
C719 B.n507 VSUBS 0.007434f
C720 B.n508 VSUBS 0.007434f
C721 B.n509 VSUBS 0.007434f
C722 B.n510 VSUBS 0.007434f
C723 B.n511 VSUBS 0.007434f
C724 B.n512 VSUBS 0.007434f
C725 B.n513 VSUBS 0.007434f
C726 B.n514 VSUBS 0.007434f
C727 B.n515 VSUBS 0.007434f
C728 B.n516 VSUBS 0.007434f
C729 B.n517 VSUBS 0.007434f
C730 B.n518 VSUBS 0.007434f
C731 B.n519 VSUBS 0.007434f
C732 B.n520 VSUBS 0.007434f
C733 B.n521 VSUBS 0.007434f
C734 B.n522 VSUBS 0.007434f
C735 B.n523 VSUBS 0.007434f
C736 B.n524 VSUBS 0.007434f
C737 B.n525 VSUBS 0.007434f
C738 B.n526 VSUBS 0.007434f
C739 B.n527 VSUBS 0.007434f
C740 B.n528 VSUBS 0.007434f
C741 B.n529 VSUBS 0.007434f
C742 B.n530 VSUBS 0.007434f
C743 B.n531 VSUBS 0.007434f
C744 B.n532 VSUBS 0.007434f
C745 B.n533 VSUBS 0.017329f
C746 B.n534 VSUBS 0.017329f
C747 B.n535 VSUBS 0.016123f
C748 B.n536 VSUBS 0.007434f
C749 B.n537 VSUBS 0.007434f
C750 B.n538 VSUBS 0.007434f
C751 B.n539 VSUBS 0.007434f
C752 B.n540 VSUBS 0.007434f
C753 B.n541 VSUBS 0.007434f
C754 B.n542 VSUBS 0.007434f
C755 B.n543 VSUBS 0.007434f
C756 B.n544 VSUBS 0.007434f
C757 B.n545 VSUBS 0.007434f
C758 B.n546 VSUBS 0.007434f
C759 B.n547 VSUBS 0.007434f
C760 B.n548 VSUBS 0.007434f
C761 B.n549 VSUBS 0.007434f
C762 B.n550 VSUBS 0.007434f
C763 B.n551 VSUBS 0.007434f
C764 B.n552 VSUBS 0.007434f
C765 B.n553 VSUBS 0.007434f
C766 B.n554 VSUBS 0.007434f
C767 B.n555 VSUBS 0.007434f
C768 B.n556 VSUBS 0.007434f
C769 B.n557 VSUBS 0.007434f
C770 B.n558 VSUBS 0.007434f
C771 B.n559 VSUBS 0.009701f
C772 B.n560 VSUBS 0.010334f
C773 B.n561 VSUBS 0.020549f
C774 VDD2.n0 VSUBS 0.027712f
C775 VDD2.n1 VSUBS 0.025122f
C776 VDD2.n2 VSUBS 0.0135f
C777 VDD2.n3 VSUBS 0.031908f
C778 VDD2.n4 VSUBS 0.014294f
C779 VDD2.n5 VSUBS 0.025122f
C780 VDD2.n6 VSUBS 0.0135f
C781 VDD2.n7 VSUBS 0.031908f
C782 VDD2.n8 VSUBS 0.014294f
C783 VDD2.n9 VSUBS 0.025122f
C784 VDD2.n10 VSUBS 0.0135f
C785 VDD2.n11 VSUBS 0.031908f
C786 VDD2.n12 VSUBS 0.013897f
C787 VDD2.n13 VSUBS 0.025122f
C788 VDD2.n14 VSUBS 0.014294f
C789 VDD2.n15 VSUBS 0.031908f
C790 VDD2.n16 VSUBS 0.014294f
C791 VDD2.n17 VSUBS 0.025122f
C792 VDD2.n18 VSUBS 0.0135f
C793 VDD2.n19 VSUBS 0.031908f
C794 VDD2.n20 VSUBS 0.014294f
C795 VDD2.n21 VSUBS 1.39945f
C796 VDD2.n22 VSUBS 0.0135f
C797 VDD2.t4 VSUBS 0.068883f
C798 VDD2.n23 VSUBS 0.214888f
C799 VDD2.n24 VSUBS 0.024003f
C800 VDD2.n25 VSUBS 0.023931f
C801 VDD2.n26 VSUBS 0.031908f
C802 VDD2.n27 VSUBS 0.014294f
C803 VDD2.n28 VSUBS 0.0135f
C804 VDD2.n29 VSUBS 0.025122f
C805 VDD2.n30 VSUBS 0.025122f
C806 VDD2.n31 VSUBS 0.0135f
C807 VDD2.n32 VSUBS 0.014294f
C808 VDD2.n33 VSUBS 0.031908f
C809 VDD2.n34 VSUBS 0.031908f
C810 VDD2.n35 VSUBS 0.014294f
C811 VDD2.n36 VSUBS 0.0135f
C812 VDD2.n37 VSUBS 0.025122f
C813 VDD2.n38 VSUBS 0.025122f
C814 VDD2.n39 VSUBS 0.0135f
C815 VDD2.n40 VSUBS 0.0135f
C816 VDD2.n41 VSUBS 0.014294f
C817 VDD2.n42 VSUBS 0.031908f
C818 VDD2.n43 VSUBS 0.031908f
C819 VDD2.n44 VSUBS 0.031908f
C820 VDD2.n45 VSUBS 0.013897f
C821 VDD2.n46 VSUBS 0.0135f
C822 VDD2.n47 VSUBS 0.025122f
C823 VDD2.n48 VSUBS 0.025122f
C824 VDD2.n49 VSUBS 0.0135f
C825 VDD2.n50 VSUBS 0.014294f
C826 VDD2.n51 VSUBS 0.031908f
C827 VDD2.n52 VSUBS 0.031908f
C828 VDD2.n53 VSUBS 0.014294f
C829 VDD2.n54 VSUBS 0.0135f
C830 VDD2.n55 VSUBS 0.025122f
C831 VDD2.n56 VSUBS 0.025122f
C832 VDD2.n57 VSUBS 0.0135f
C833 VDD2.n58 VSUBS 0.014294f
C834 VDD2.n59 VSUBS 0.031908f
C835 VDD2.n60 VSUBS 0.031908f
C836 VDD2.n61 VSUBS 0.014294f
C837 VDD2.n62 VSUBS 0.0135f
C838 VDD2.n63 VSUBS 0.025122f
C839 VDD2.n64 VSUBS 0.025122f
C840 VDD2.n65 VSUBS 0.0135f
C841 VDD2.n66 VSUBS 0.014294f
C842 VDD2.n67 VSUBS 0.031908f
C843 VDD2.n68 VSUBS 0.077614f
C844 VDD2.n69 VSUBS 0.014294f
C845 VDD2.n70 VSUBS 0.0135f
C846 VDD2.n71 VSUBS 0.056009f
C847 VDD2.n72 VSUBS 0.05717f
C848 VDD2.t1 VSUBS 0.268006f
C849 VDD2.t3 VSUBS 0.268006f
C850 VDD2.n73 VSUBS 2.12748f
C851 VDD2.n74 VSUBS 2.13125f
C852 VDD2.n75 VSUBS 0.027712f
C853 VDD2.n76 VSUBS 0.025122f
C854 VDD2.n77 VSUBS 0.0135f
C855 VDD2.n78 VSUBS 0.031908f
C856 VDD2.n79 VSUBS 0.014294f
C857 VDD2.n80 VSUBS 0.025122f
C858 VDD2.n81 VSUBS 0.0135f
C859 VDD2.n82 VSUBS 0.031908f
C860 VDD2.n83 VSUBS 0.014294f
C861 VDD2.n84 VSUBS 0.025122f
C862 VDD2.n85 VSUBS 0.0135f
C863 VDD2.n86 VSUBS 0.031908f
C864 VDD2.n87 VSUBS 0.013897f
C865 VDD2.n88 VSUBS 0.025122f
C866 VDD2.n89 VSUBS 0.013897f
C867 VDD2.n90 VSUBS 0.0135f
C868 VDD2.n91 VSUBS 0.031908f
C869 VDD2.n92 VSUBS 0.031908f
C870 VDD2.n93 VSUBS 0.014294f
C871 VDD2.n94 VSUBS 0.025122f
C872 VDD2.n95 VSUBS 0.0135f
C873 VDD2.n96 VSUBS 0.031908f
C874 VDD2.n97 VSUBS 0.014294f
C875 VDD2.n98 VSUBS 1.39945f
C876 VDD2.n99 VSUBS 0.0135f
C877 VDD2.t5 VSUBS 0.068883f
C878 VDD2.n100 VSUBS 0.214888f
C879 VDD2.n101 VSUBS 0.024003f
C880 VDD2.n102 VSUBS 0.023931f
C881 VDD2.n103 VSUBS 0.031908f
C882 VDD2.n104 VSUBS 0.014294f
C883 VDD2.n105 VSUBS 0.0135f
C884 VDD2.n106 VSUBS 0.025122f
C885 VDD2.n107 VSUBS 0.025122f
C886 VDD2.n108 VSUBS 0.0135f
C887 VDD2.n109 VSUBS 0.014294f
C888 VDD2.n110 VSUBS 0.031908f
C889 VDD2.n111 VSUBS 0.031908f
C890 VDD2.n112 VSUBS 0.014294f
C891 VDD2.n113 VSUBS 0.0135f
C892 VDD2.n114 VSUBS 0.025122f
C893 VDD2.n115 VSUBS 0.025122f
C894 VDD2.n116 VSUBS 0.0135f
C895 VDD2.n117 VSUBS 0.014294f
C896 VDD2.n118 VSUBS 0.031908f
C897 VDD2.n119 VSUBS 0.031908f
C898 VDD2.n120 VSUBS 0.014294f
C899 VDD2.n121 VSUBS 0.0135f
C900 VDD2.n122 VSUBS 0.025122f
C901 VDD2.n123 VSUBS 0.025122f
C902 VDD2.n124 VSUBS 0.0135f
C903 VDD2.n125 VSUBS 0.014294f
C904 VDD2.n126 VSUBS 0.031908f
C905 VDD2.n127 VSUBS 0.031908f
C906 VDD2.n128 VSUBS 0.014294f
C907 VDD2.n129 VSUBS 0.0135f
C908 VDD2.n130 VSUBS 0.025122f
C909 VDD2.n131 VSUBS 0.025122f
C910 VDD2.n132 VSUBS 0.0135f
C911 VDD2.n133 VSUBS 0.014294f
C912 VDD2.n134 VSUBS 0.031908f
C913 VDD2.n135 VSUBS 0.031908f
C914 VDD2.n136 VSUBS 0.014294f
C915 VDD2.n137 VSUBS 0.0135f
C916 VDD2.n138 VSUBS 0.025122f
C917 VDD2.n139 VSUBS 0.025122f
C918 VDD2.n140 VSUBS 0.0135f
C919 VDD2.n141 VSUBS 0.014294f
C920 VDD2.n142 VSUBS 0.031908f
C921 VDD2.n143 VSUBS 0.077614f
C922 VDD2.n144 VSUBS 0.014294f
C923 VDD2.n145 VSUBS 0.0135f
C924 VDD2.n146 VSUBS 0.056009f
C925 VDD2.n147 VSUBS 0.056346f
C926 VDD2.n148 VSUBS 2.10759f
C927 VDD2.t0 VSUBS 0.268006f
C928 VDD2.t2 VSUBS 0.268006f
C929 VDD2.n149 VSUBS 2.12745f
C930 VTAIL.t6 VSUBS 0.326123f
C931 VTAIL.t7 VSUBS 0.326123f
C932 VTAIL.n0 VSUBS 2.40772f
C933 VTAIL.n1 VSUBS 0.834586f
C934 VTAIL.n2 VSUBS 0.033721f
C935 VTAIL.n3 VSUBS 0.03057f
C936 VTAIL.n4 VSUBS 0.016427f
C937 VTAIL.n5 VSUBS 0.038827f
C938 VTAIL.n6 VSUBS 0.017393f
C939 VTAIL.n7 VSUBS 0.03057f
C940 VTAIL.n8 VSUBS 0.016427f
C941 VTAIL.n9 VSUBS 0.038827f
C942 VTAIL.n10 VSUBS 0.017393f
C943 VTAIL.n11 VSUBS 0.03057f
C944 VTAIL.n12 VSUBS 0.016427f
C945 VTAIL.n13 VSUBS 0.038827f
C946 VTAIL.n14 VSUBS 0.01691f
C947 VTAIL.n15 VSUBS 0.03057f
C948 VTAIL.n16 VSUBS 0.017393f
C949 VTAIL.n17 VSUBS 0.038827f
C950 VTAIL.n18 VSUBS 0.017393f
C951 VTAIL.n19 VSUBS 0.03057f
C952 VTAIL.n20 VSUBS 0.016427f
C953 VTAIL.n21 VSUBS 0.038827f
C954 VTAIL.n22 VSUBS 0.017393f
C955 VTAIL.n23 VSUBS 1.70292f
C956 VTAIL.n24 VSUBS 0.016427f
C957 VTAIL.t2 VSUBS 0.08382f
C958 VTAIL.n25 VSUBS 0.261487f
C959 VTAIL.n26 VSUBS 0.029208f
C960 VTAIL.n27 VSUBS 0.02912f
C961 VTAIL.n28 VSUBS 0.038827f
C962 VTAIL.n29 VSUBS 0.017393f
C963 VTAIL.n30 VSUBS 0.016427f
C964 VTAIL.n31 VSUBS 0.03057f
C965 VTAIL.n32 VSUBS 0.03057f
C966 VTAIL.n33 VSUBS 0.016427f
C967 VTAIL.n34 VSUBS 0.017393f
C968 VTAIL.n35 VSUBS 0.038827f
C969 VTAIL.n36 VSUBS 0.038827f
C970 VTAIL.n37 VSUBS 0.017393f
C971 VTAIL.n38 VSUBS 0.016427f
C972 VTAIL.n39 VSUBS 0.03057f
C973 VTAIL.n40 VSUBS 0.03057f
C974 VTAIL.n41 VSUBS 0.016427f
C975 VTAIL.n42 VSUBS 0.016427f
C976 VTAIL.n43 VSUBS 0.017393f
C977 VTAIL.n44 VSUBS 0.038827f
C978 VTAIL.n45 VSUBS 0.038827f
C979 VTAIL.n46 VSUBS 0.038827f
C980 VTAIL.n47 VSUBS 0.01691f
C981 VTAIL.n48 VSUBS 0.016427f
C982 VTAIL.n49 VSUBS 0.03057f
C983 VTAIL.n50 VSUBS 0.03057f
C984 VTAIL.n51 VSUBS 0.016427f
C985 VTAIL.n52 VSUBS 0.017393f
C986 VTAIL.n53 VSUBS 0.038827f
C987 VTAIL.n54 VSUBS 0.038827f
C988 VTAIL.n55 VSUBS 0.017393f
C989 VTAIL.n56 VSUBS 0.016427f
C990 VTAIL.n57 VSUBS 0.03057f
C991 VTAIL.n58 VSUBS 0.03057f
C992 VTAIL.n59 VSUBS 0.016427f
C993 VTAIL.n60 VSUBS 0.017393f
C994 VTAIL.n61 VSUBS 0.038827f
C995 VTAIL.n62 VSUBS 0.038827f
C996 VTAIL.n63 VSUBS 0.017393f
C997 VTAIL.n64 VSUBS 0.016427f
C998 VTAIL.n65 VSUBS 0.03057f
C999 VTAIL.n66 VSUBS 0.03057f
C1000 VTAIL.n67 VSUBS 0.016427f
C1001 VTAIL.n68 VSUBS 0.017393f
C1002 VTAIL.n69 VSUBS 0.038827f
C1003 VTAIL.n70 VSUBS 0.094444f
C1004 VTAIL.n71 VSUBS 0.017393f
C1005 VTAIL.n72 VSUBS 0.016427f
C1006 VTAIL.n73 VSUBS 0.068155f
C1007 VTAIL.n74 VSUBS 0.047437f
C1008 VTAIL.n75 VSUBS 0.172875f
C1009 VTAIL.t5 VSUBS 0.326123f
C1010 VTAIL.t0 VSUBS 0.326123f
C1011 VTAIL.n76 VSUBS 2.40772f
C1012 VTAIL.n77 VSUBS 2.49705f
C1013 VTAIL.t8 VSUBS 0.326123f
C1014 VTAIL.t9 VSUBS 0.326123f
C1015 VTAIL.n78 VSUBS 2.40774f
C1016 VTAIL.n79 VSUBS 2.49703f
C1017 VTAIL.n80 VSUBS 0.033721f
C1018 VTAIL.n81 VSUBS 0.03057f
C1019 VTAIL.n82 VSUBS 0.016427f
C1020 VTAIL.n83 VSUBS 0.038827f
C1021 VTAIL.n84 VSUBS 0.017393f
C1022 VTAIL.n85 VSUBS 0.03057f
C1023 VTAIL.n86 VSUBS 0.016427f
C1024 VTAIL.n87 VSUBS 0.038827f
C1025 VTAIL.n88 VSUBS 0.017393f
C1026 VTAIL.n89 VSUBS 0.03057f
C1027 VTAIL.n90 VSUBS 0.016427f
C1028 VTAIL.n91 VSUBS 0.038827f
C1029 VTAIL.n92 VSUBS 0.01691f
C1030 VTAIL.n93 VSUBS 0.03057f
C1031 VTAIL.n94 VSUBS 0.01691f
C1032 VTAIL.n95 VSUBS 0.016427f
C1033 VTAIL.n96 VSUBS 0.038827f
C1034 VTAIL.n97 VSUBS 0.038827f
C1035 VTAIL.n98 VSUBS 0.017393f
C1036 VTAIL.n99 VSUBS 0.03057f
C1037 VTAIL.n100 VSUBS 0.016427f
C1038 VTAIL.n101 VSUBS 0.038827f
C1039 VTAIL.n102 VSUBS 0.017393f
C1040 VTAIL.n103 VSUBS 1.70292f
C1041 VTAIL.n104 VSUBS 0.016427f
C1042 VTAIL.t11 VSUBS 0.08382f
C1043 VTAIL.n105 VSUBS 0.261487f
C1044 VTAIL.n106 VSUBS 0.029208f
C1045 VTAIL.n107 VSUBS 0.02912f
C1046 VTAIL.n108 VSUBS 0.038827f
C1047 VTAIL.n109 VSUBS 0.017393f
C1048 VTAIL.n110 VSUBS 0.016427f
C1049 VTAIL.n111 VSUBS 0.03057f
C1050 VTAIL.n112 VSUBS 0.03057f
C1051 VTAIL.n113 VSUBS 0.016427f
C1052 VTAIL.n114 VSUBS 0.017393f
C1053 VTAIL.n115 VSUBS 0.038827f
C1054 VTAIL.n116 VSUBS 0.038827f
C1055 VTAIL.n117 VSUBS 0.017393f
C1056 VTAIL.n118 VSUBS 0.016427f
C1057 VTAIL.n119 VSUBS 0.03057f
C1058 VTAIL.n120 VSUBS 0.03057f
C1059 VTAIL.n121 VSUBS 0.016427f
C1060 VTAIL.n122 VSUBS 0.017393f
C1061 VTAIL.n123 VSUBS 0.038827f
C1062 VTAIL.n124 VSUBS 0.038827f
C1063 VTAIL.n125 VSUBS 0.017393f
C1064 VTAIL.n126 VSUBS 0.016427f
C1065 VTAIL.n127 VSUBS 0.03057f
C1066 VTAIL.n128 VSUBS 0.03057f
C1067 VTAIL.n129 VSUBS 0.016427f
C1068 VTAIL.n130 VSUBS 0.017393f
C1069 VTAIL.n131 VSUBS 0.038827f
C1070 VTAIL.n132 VSUBS 0.038827f
C1071 VTAIL.n133 VSUBS 0.017393f
C1072 VTAIL.n134 VSUBS 0.016427f
C1073 VTAIL.n135 VSUBS 0.03057f
C1074 VTAIL.n136 VSUBS 0.03057f
C1075 VTAIL.n137 VSUBS 0.016427f
C1076 VTAIL.n138 VSUBS 0.017393f
C1077 VTAIL.n139 VSUBS 0.038827f
C1078 VTAIL.n140 VSUBS 0.038827f
C1079 VTAIL.n141 VSUBS 0.017393f
C1080 VTAIL.n142 VSUBS 0.016427f
C1081 VTAIL.n143 VSUBS 0.03057f
C1082 VTAIL.n144 VSUBS 0.03057f
C1083 VTAIL.n145 VSUBS 0.016427f
C1084 VTAIL.n146 VSUBS 0.017393f
C1085 VTAIL.n147 VSUBS 0.038827f
C1086 VTAIL.n148 VSUBS 0.094444f
C1087 VTAIL.n149 VSUBS 0.017393f
C1088 VTAIL.n150 VSUBS 0.016427f
C1089 VTAIL.n151 VSUBS 0.068155f
C1090 VTAIL.n152 VSUBS 0.047437f
C1091 VTAIL.n153 VSUBS 0.172875f
C1092 VTAIL.t1 VSUBS 0.326123f
C1093 VTAIL.t4 VSUBS 0.326123f
C1094 VTAIL.n154 VSUBS 2.40774f
C1095 VTAIL.n155 VSUBS 0.879787f
C1096 VTAIL.n156 VSUBS 0.033721f
C1097 VTAIL.n157 VSUBS 0.03057f
C1098 VTAIL.n158 VSUBS 0.016427f
C1099 VTAIL.n159 VSUBS 0.038827f
C1100 VTAIL.n160 VSUBS 0.017393f
C1101 VTAIL.n161 VSUBS 0.03057f
C1102 VTAIL.n162 VSUBS 0.016427f
C1103 VTAIL.n163 VSUBS 0.038827f
C1104 VTAIL.n164 VSUBS 0.017393f
C1105 VTAIL.n165 VSUBS 0.03057f
C1106 VTAIL.n166 VSUBS 0.016427f
C1107 VTAIL.n167 VSUBS 0.038827f
C1108 VTAIL.n168 VSUBS 0.01691f
C1109 VTAIL.n169 VSUBS 0.03057f
C1110 VTAIL.n170 VSUBS 0.01691f
C1111 VTAIL.n171 VSUBS 0.016427f
C1112 VTAIL.n172 VSUBS 0.038827f
C1113 VTAIL.n173 VSUBS 0.038827f
C1114 VTAIL.n174 VSUBS 0.017393f
C1115 VTAIL.n175 VSUBS 0.03057f
C1116 VTAIL.n176 VSUBS 0.016427f
C1117 VTAIL.n177 VSUBS 0.038827f
C1118 VTAIL.n178 VSUBS 0.017393f
C1119 VTAIL.n179 VSUBS 1.70292f
C1120 VTAIL.n180 VSUBS 0.016427f
C1121 VTAIL.t3 VSUBS 0.08382f
C1122 VTAIL.n181 VSUBS 0.261487f
C1123 VTAIL.n182 VSUBS 0.029208f
C1124 VTAIL.n183 VSUBS 0.02912f
C1125 VTAIL.n184 VSUBS 0.038827f
C1126 VTAIL.n185 VSUBS 0.017393f
C1127 VTAIL.n186 VSUBS 0.016427f
C1128 VTAIL.n187 VSUBS 0.03057f
C1129 VTAIL.n188 VSUBS 0.03057f
C1130 VTAIL.n189 VSUBS 0.016427f
C1131 VTAIL.n190 VSUBS 0.017393f
C1132 VTAIL.n191 VSUBS 0.038827f
C1133 VTAIL.n192 VSUBS 0.038827f
C1134 VTAIL.n193 VSUBS 0.017393f
C1135 VTAIL.n194 VSUBS 0.016427f
C1136 VTAIL.n195 VSUBS 0.03057f
C1137 VTAIL.n196 VSUBS 0.03057f
C1138 VTAIL.n197 VSUBS 0.016427f
C1139 VTAIL.n198 VSUBS 0.017393f
C1140 VTAIL.n199 VSUBS 0.038827f
C1141 VTAIL.n200 VSUBS 0.038827f
C1142 VTAIL.n201 VSUBS 0.017393f
C1143 VTAIL.n202 VSUBS 0.016427f
C1144 VTAIL.n203 VSUBS 0.03057f
C1145 VTAIL.n204 VSUBS 0.03057f
C1146 VTAIL.n205 VSUBS 0.016427f
C1147 VTAIL.n206 VSUBS 0.017393f
C1148 VTAIL.n207 VSUBS 0.038827f
C1149 VTAIL.n208 VSUBS 0.038827f
C1150 VTAIL.n209 VSUBS 0.017393f
C1151 VTAIL.n210 VSUBS 0.016427f
C1152 VTAIL.n211 VSUBS 0.03057f
C1153 VTAIL.n212 VSUBS 0.03057f
C1154 VTAIL.n213 VSUBS 0.016427f
C1155 VTAIL.n214 VSUBS 0.017393f
C1156 VTAIL.n215 VSUBS 0.038827f
C1157 VTAIL.n216 VSUBS 0.038827f
C1158 VTAIL.n217 VSUBS 0.017393f
C1159 VTAIL.n218 VSUBS 0.016427f
C1160 VTAIL.n219 VSUBS 0.03057f
C1161 VTAIL.n220 VSUBS 0.03057f
C1162 VTAIL.n221 VSUBS 0.016427f
C1163 VTAIL.n222 VSUBS 0.017393f
C1164 VTAIL.n223 VSUBS 0.038827f
C1165 VTAIL.n224 VSUBS 0.094444f
C1166 VTAIL.n225 VSUBS 0.017393f
C1167 VTAIL.n226 VSUBS 0.016427f
C1168 VTAIL.n227 VSUBS 0.068155f
C1169 VTAIL.n228 VSUBS 0.047437f
C1170 VTAIL.n229 VSUBS 1.72219f
C1171 VTAIL.n230 VSUBS 0.033721f
C1172 VTAIL.n231 VSUBS 0.03057f
C1173 VTAIL.n232 VSUBS 0.016427f
C1174 VTAIL.n233 VSUBS 0.038827f
C1175 VTAIL.n234 VSUBS 0.017393f
C1176 VTAIL.n235 VSUBS 0.03057f
C1177 VTAIL.n236 VSUBS 0.016427f
C1178 VTAIL.n237 VSUBS 0.038827f
C1179 VTAIL.n238 VSUBS 0.017393f
C1180 VTAIL.n239 VSUBS 0.03057f
C1181 VTAIL.n240 VSUBS 0.016427f
C1182 VTAIL.n241 VSUBS 0.038827f
C1183 VTAIL.n242 VSUBS 0.01691f
C1184 VTAIL.n243 VSUBS 0.03057f
C1185 VTAIL.n244 VSUBS 0.017393f
C1186 VTAIL.n245 VSUBS 0.038827f
C1187 VTAIL.n246 VSUBS 0.017393f
C1188 VTAIL.n247 VSUBS 0.03057f
C1189 VTAIL.n248 VSUBS 0.016427f
C1190 VTAIL.n249 VSUBS 0.038827f
C1191 VTAIL.n250 VSUBS 0.017393f
C1192 VTAIL.n251 VSUBS 1.70292f
C1193 VTAIL.n252 VSUBS 0.016427f
C1194 VTAIL.t10 VSUBS 0.08382f
C1195 VTAIL.n253 VSUBS 0.261487f
C1196 VTAIL.n254 VSUBS 0.029208f
C1197 VTAIL.n255 VSUBS 0.02912f
C1198 VTAIL.n256 VSUBS 0.038827f
C1199 VTAIL.n257 VSUBS 0.017393f
C1200 VTAIL.n258 VSUBS 0.016427f
C1201 VTAIL.n259 VSUBS 0.03057f
C1202 VTAIL.n260 VSUBS 0.03057f
C1203 VTAIL.n261 VSUBS 0.016427f
C1204 VTAIL.n262 VSUBS 0.017393f
C1205 VTAIL.n263 VSUBS 0.038827f
C1206 VTAIL.n264 VSUBS 0.038827f
C1207 VTAIL.n265 VSUBS 0.017393f
C1208 VTAIL.n266 VSUBS 0.016427f
C1209 VTAIL.n267 VSUBS 0.03057f
C1210 VTAIL.n268 VSUBS 0.03057f
C1211 VTAIL.n269 VSUBS 0.016427f
C1212 VTAIL.n270 VSUBS 0.016427f
C1213 VTAIL.n271 VSUBS 0.017393f
C1214 VTAIL.n272 VSUBS 0.038827f
C1215 VTAIL.n273 VSUBS 0.038827f
C1216 VTAIL.n274 VSUBS 0.038827f
C1217 VTAIL.n275 VSUBS 0.01691f
C1218 VTAIL.n276 VSUBS 0.016427f
C1219 VTAIL.n277 VSUBS 0.03057f
C1220 VTAIL.n278 VSUBS 0.03057f
C1221 VTAIL.n279 VSUBS 0.016427f
C1222 VTAIL.n280 VSUBS 0.017393f
C1223 VTAIL.n281 VSUBS 0.038827f
C1224 VTAIL.n282 VSUBS 0.038827f
C1225 VTAIL.n283 VSUBS 0.017393f
C1226 VTAIL.n284 VSUBS 0.016427f
C1227 VTAIL.n285 VSUBS 0.03057f
C1228 VTAIL.n286 VSUBS 0.03057f
C1229 VTAIL.n287 VSUBS 0.016427f
C1230 VTAIL.n288 VSUBS 0.017393f
C1231 VTAIL.n289 VSUBS 0.038827f
C1232 VTAIL.n290 VSUBS 0.038827f
C1233 VTAIL.n291 VSUBS 0.017393f
C1234 VTAIL.n292 VSUBS 0.016427f
C1235 VTAIL.n293 VSUBS 0.03057f
C1236 VTAIL.n294 VSUBS 0.03057f
C1237 VTAIL.n295 VSUBS 0.016427f
C1238 VTAIL.n296 VSUBS 0.017393f
C1239 VTAIL.n297 VSUBS 0.038827f
C1240 VTAIL.n298 VSUBS 0.094444f
C1241 VTAIL.n299 VSUBS 0.017393f
C1242 VTAIL.n300 VSUBS 0.016427f
C1243 VTAIL.n301 VSUBS 0.068155f
C1244 VTAIL.n302 VSUBS 0.047437f
C1245 VTAIL.n303 VSUBS 1.69947f
C1246 VN.t1 VSUBS 1.1517f
C1247 VN.n0 VSUBS 0.438739f
C1248 VN.t4 VSUBS 1.13675f
C1249 VN.n1 VSUBS 0.458449f
C1250 VN.t2 VSUBS 1.14205f
C1251 VN.n2 VSUBS 0.447903f
C1252 VN.n3 VSUBS 0.196315f
C1253 VN.t3 VSUBS 1.1517f
C1254 VN.n4 VSUBS 0.438739f
C1255 VN.t0 VSUBS 1.14205f
C1256 VN.t5 VSUBS 1.13675f
C1257 VN.n5 VSUBS 0.458449f
C1258 VN.n6 VSUBS 0.447903f
C1259 VN.n7 VSUBS 2.74423f
.ends

