* NGSPICE file created from diff_pair_sample_0237.ext - technology: sky130A

.subckt diff_pair_sample_0237 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t10 B.t6 sky130_fd_pr__nfet_01v8 ad=1.848 pd=11.53 as=4.368 ps=23.18 w=11.2 l=1.59
X1 VTAIL.t14 VP.t1 VDD1.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=4.368 pd=23.18 as=1.848 ps=11.53 w=11.2 l=1.59
X2 B.t21 B.t19 B.t20 B.t13 sky130_fd_pr__nfet_01v8 ad=4.368 pd=23.18 as=0 ps=0 w=11.2 l=1.59
X3 B.t18 B.t16 B.t17 B.t9 sky130_fd_pr__nfet_01v8 ad=4.368 pd=23.18 as=0 ps=0 w=11.2 l=1.59
X4 VDD2.t7 VN.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.848 pd=11.53 as=1.848 ps=11.53 w=11.2 l=1.59
X5 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=4.368 pd=23.18 as=0 ps=0 w=11.2 l=1.59
X6 VTAIL.t3 VN.t1 VDD2.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=4.368 pd=23.18 as=1.848 ps=11.53 w=11.2 l=1.59
X7 VTAIL.t0 VN.t2 VDD2.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=4.368 pd=23.18 as=1.848 ps=11.53 w=11.2 l=1.59
X8 VDD1.t5 VP.t2 VTAIL.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=1.848 pd=11.53 as=1.848 ps=11.53 w=11.2 l=1.59
X9 VDD2.t4 VN.t3 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=1.848 pd=11.53 as=4.368 ps=23.18 w=11.2 l=1.59
X10 VDD2.t3 VN.t4 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.848 pd=11.53 as=1.848 ps=11.53 w=11.2 l=1.59
X11 VDD2.t2 VN.t5 VTAIL.t15 B.t7 sky130_fd_pr__nfet_01v8 ad=1.848 pd=11.53 as=4.368 ps=23.18 w=11.2 l=1.59
X12 VTAIL.t2 VN.t6 VDD2.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=1.848 pd=11.53 as=1.848 ps=11.53 w=11.2 l=1.59
X13 VDD1.t4 VP.t3 VTAIL.t12 B.t7 sky130_fd_pr__nfet_01v8 ad=1.848 pd=11.53 as=4.368 ps=23.18 w=11.2 l=1.59
X14 VTAIL.t11 VP.t4 VDD1.t3 B.t4 sky130_fd_pr__nfet_01v8 ad=1.848 pd=11.53 as=1.848 ps=11.53 w=11.2 l=1.59
X15 VDD1.t2 VP.t5 VTAIL.t9 B.t1 sky130_fd_pr__nfet_01v8 ad=1.848 pd=11.53 as=1.848 ps=11.53 w=11.2 l=1.59
X16 VTAIL.t8 VP.t6 VDD1.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=4.368 pd=23.18 as=1.848 ps=11.53 w=11.2 l=1.59
X17 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=4.368 pd=23.18 as=0 ps=0 w=11.2 l=1.59
X18 VTAIL.t7 VP.t7 VDD1.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=1.848 pd=11.53 as=1.848 ps=11.53 w=11.2 l=1.59
X19 VTAIL.t4 VN.t7 VDD2.t0 B.t4 sky130_fd_pr__nfet_01v8 ad=1.848 pd=11.53 as=1.848 ps=11.53 w=11.2 l=1.59
R0 VP.n10 VP.t6 201.624
R1 VP.n28 VP.n27 179.499
R2 VP.n50 VP.n49 179.499
R3 VP.n26 VP.n25 179.499
R4 VP.n28 VP.t1 169.762
R5 VP.n35 VP.t2 169.762
R6 VP.n42 VP.t7 169.762
R7 VP.n49 VP.t0 169.762
R8 VP.n25 VP.t3 169.762
R9 VP.n18 VP.t4 169.762
R10 VP.n11 VP.t5 169.762
R11 VP.n13 VP.n12 161.3
R12 VP.n14 VP.n9 161.3
R13 VP.n16 VP.n15 161.3
R14 VP.n17 VP.n8 161.3
R15 VP.n20 VP.n19 161.3
R16 VP.n21 VP.n7 161.3
R17 VP.n23 VP.n22 161.3
R18 VP.n24 VP.n6 161.3
R19 VP.n48 VP.n0 161.3
R20 VP.n47 VP.n46 161.3
R21 VP.n45 VP.n1 161.3
R22 VP.n44 VP.n43 161.3
R23 VP.n41 VP.n2 161.3
R24 VP.n40 VP.n39 161.3
R25 VP.n38 VP.n3 161.3
R26 VP.n37 VP.n36 161.3
R27 VP.n34 VP.n4 161.3
R28 VP.n33 VP.n32 161.3
R29 VP.n31 VP.n5 161.3
R30 VP.n30 VP.n29 161.3
R31 VP.n40 VP.n3 56.5617
R32 VP.n16 VP.n9 56.5617
R33 VP.n33 VP.n5 56.5617
R34 VP.n47 VP.n1 56.5617
R35 VP.n23 VP.n7 56.5617
R36 VP.n11 VP.n10 55.8951
R37 VP.n27 VP.n26 45.455
R38 VP.n29 VP.n5 24.5923
R39 VP.n34 VP.n33 24.5923
R40 VP.n36 VP.n3 24.5923
R41 VP.n41 VP.n40 24.5923
R42 VP.n43 VP.n1 24.5923
R43 VP.n48 VP.n47 24.5923
R44 VP.n24 VP.n23 24.5923
R45 VP.n17 VP.n16 24.5923
R46 VP.n19 VP.n7 24.5923
R47 VP.n12 VP.n9 24.5923
R48 VP.n13 VP.n10 18.12
R49 VP.n35 VP.n34 14.2638
R50 VP.n43 VP.n42 14.2638
R51 VP.n19 VP.n18 14.2638
R52 VP.n36 VP.n35 10.3291
R53 VP.n42 VP.n41 10.3291
R54 VP.n18 VP.n17 10.3291
R55 VP.n12 VP.n11 10.3291
R56 VP.n29 VP.n28 6.39438
R57 VP.n49 VP.n48 6.39438
R58 VP.n25 VP.n24 6.39438
R59 VP.n14 VP.n13 0.189894
R60 VP.n15 VP.n14 0.189894
R61 VP.n15 VP.n8 0.189894
R62 VP.n20 VP.n8 0.189894
R63 VP.n21 VP.n20 0.189894
R64 VP.n22 VP.n21 0.189894
R65 VP.n22 VP.n6 0.189894
R66 VP.n26 VP.n6 0.189894
R67 VP.n30 VP.n27 0.189894
R68 VP.n31 VP.n30 0.189894
R69 VP.n32 VP.n31 0.189894
R70 VP.n32 VP.n4 0.189894
R71 VP.n37 VP.n4 0.189894
R72 VP.n38 VP.n37 0.189894
R73 VP.n39 VP.n38 0.189894
R74 VP.n39 VP.n2 0.189894
R75 VP.n44 VP.n2 0.189894
R76 VP.n45 VP.n44 0.189894
R77 VP.n46 VP.n45 0.189894
R78 VP.n46 VP.n0 0.189894
R79 VP.n50 VP.n0 0.189894
R80 VP VP.n50 0.0516364
R81 VTAIL.n11 VTAIL.t8 50.4012
R82 VTAIL.n10 VTAIL.t6 50.4012
R83 VTAIL.n7 VTAIL.t0 50.4012
R84 VTAIL.n15 VTAIL.t15 50.4011
R85 VTAIL.n2 VTAIL.t3 50.4011
R86 VTAIL.n3 VTAIL.t10 50.4011
R87 VTAIL.n6 VTAIL.t14 50.4011
R88 VTAIL.n14 VTAIL.t12 50.4011
R89 VTAIL.n13 VTAIL.n12 48.6334
R90 VTAIL.n9 VTAIL.n8 48.6334
R91 VTAIL.n1 VTAIL.n0 48.6331
R92 VTAIL.n5 VTAIL.n4 48.6331
R93 VTAIL.n15 VTAIL.n14 23.6772
R94 VTAIL.n7 VTAIL.n6 23.6772
R95 VTAIL.n0 VTAIL.t1 1.76836
R96 VTAIL.n0 VTAIL.t4 1.76836
R97 VTAIL.n4 VTAIL.t13 1.76836
R98 VTAIL.n4 VTAIL.t7 1.76836
R99 VTAIL.n12 VTAIL.t9 1.76836
R100 VTAIL.n12 VTAIL.t11 1.76836
R101 VTAIL.n8 VTAIL.t5 1.76836
R102 VTAIL.n8 VTAIL.t2 1.76836
R103 VTAIL.n9 VTAIL.n7 1.65567
R104 VTAIL.n10 VTAIL.n9 1.65567
R105 VTAIL.n13 VTAIL.n11 1.65567
R106 VTAIL.n14 VTAIL.n13 1.65567
R107 VTAIL.n6 VTAIL.n5 1.65567
R108 VTAIL.n5 VTAIL.n3 1.65567
R109 VTAIL.n2 VTAIL.n1 1.65567
R110 VTAIL VTAIL.n15 1.59748
R111 VTAIL.n11 VTAIL.n10 0.470328
R112 VTAIL.n3 VTAIL.n2 0.470328
R113 VTAIL VTAIL.n1 0.0586897
R114 VDD1 VDD1.n0 66.1979
R115 VDD1.n3 VDD1.n2 66.0842
R116 VDD1.n3 VDD1.n1 66.0842
R117 VDD1.n5 VDD1.n4 65.312
R118 VDD1.n5 VDD1.n3 41.4018
R119 VDD1.n4 VDD1.t3 1.76836
R120 VDD1.n4 VDD1.t4 1.76836
R121 VDD1.n0 VDD1.t1 1.76836
R122 VDD1.n0 VDD1.t2 1.76836
R123 VDD1.n2 VDD1.t0 1.76836
R124 VDD1.n2 VDD1.t7 1.76836
R125 VDD1.n1 VDD1.t6 1.76836
R126 VDD1.n1 VDD1.t5 1.76836
R127 VDD1 VDD1.n5 0.769897
R128 B.n743 B.n742 585
R129 B.n289 B.n112 585
R130 B.n288 B.n287 585
R131 B.n286 B.n285 585
R132 B.n284 B.n283 585
R133 B.n282 B.n281 585
R134 B.n280 B.n279 585
R135 B.n278 B.n277 585
R136 B.n276 B.n275 585
R137 B.n274 B.n273 585
R138 B.n272 B.n271 585
R139 B.n270 B.n269 585
R140 B.n268 B.n267 585
R141 B.n266 B.n265 585
R142 B.n264 B.n263 585
R143 B.n262 B.n261 585
R144 B.n260 B.n259 585
R145 B.n258 B.n257 585
R146 B.n256 B.n255 585
R147 B.n254 B.n253 585
R148 B.n252 B.n251 585
R149 B.n250 B.n249 585
R150 B.n248 B.n247 585
R151 B.n246 B.n245 585
R152 B.n244 B.n243 585
R153 B.n242 B.n241 585
R154 B.n240 B.n239 585
R155 B.n238 B.n237 585
R156 B.n236 B.n235 585
R157 B.n234 B.n233 585
R158 B.n232 B.n231 585
R159 B.n230 B.n229 585
R160 B.n228 B.n227 585
R161 B.n226 B.n225 585
R162 B.n224 B.n223 585
R163 B.n222 B.n221 585
R164 B.n220 B.n219 585
R165 B.n218 B.n217 585
R166 B.n216 B.n215 585
R167 B.n213 B.n212 585
R168 B.n211 B.n210 585
R169 B.n209 B.n208 585
R170 B.n207 B.n206 585
R171 B.n205 B.n204 585
R172 B.n203 B.n202 585
R173 B.n201 B.n200 585
R174 B.n199 B.n198 585
R175 B.n197 B.n196 585
R176 B.n195 B.n194 585
R177 B.n192 B.n191 585
R178 B.n190 B.n189 585
R179 B.n188 B.n187 585
R180 B.n186 B.n185 585
R181 B.n184 B.n183 585
R182 B.n182 B.n181 585
R183 B.n180 B.n179 585
R184 B.n178 B.n177 585
R185 B.n176 B.n175 585
R186 B.n174 B.n173 585
R187 B.n172 B.n171 585
R188 B.n170 B.n169 585
R189 B.n168 B.n167 585
R190 B.n166 B.n165 585
R191 B.n164 B.n163 585
R192 B.n162 B.n161 585
R193 B.n160 B.n159 585
R194 B.n158 B.n157 585
R195 B.n156 B.n155 585
R196 B.n154 B.n153 585
R197 B.n152 B.n151 585
R198 B.n150 B.n149 585
R199 B.n148 B.n147 585
R200 B.n146 B.n145 585
R201 B.n144 B.n143 585
R202 B.n142 B.n141 585
R203 B.n140 B.n139 585
R204 B.n138 B.n137 585
R205 B.n136 B.n135 585
R206 B.n134 B.n133 585
R207 B.n132 B.n131 585
R208 B.n130 B.n129 585
R209 B.n128 B.n127 585
R210 B.n126 B.n125 585
R211 B.n124 B.n123 585
R212 B.n122 B.n121 585
R213 B.n120 B.n119 585
R214 B.n118 B.n117 585
R215 B.n67 B.n66 585
R216 B.n741 B.n68 585
R217 B.n746 B.n68 585
R218 B.n740 B.n739 585
R219 B.n739 B.n64 585
R220 B.n738 B.n63 585
R221 B.n752 B.n63 585
R222 B.n737 B.n62 585
R223 B.n753 B.n62 585
R224 B.n736 B.n61 585
R225 B.n754 B.n61 585
R226 B.n735 B.n734 585
R227 B.n734 B.n57 585
R228 B.n733 B.n56 585
R229 B.n760 B.n56 585
R230 B.n732 B.n55 585
R231 B.n761 B.n55 585
R232 B.n731 B.n54 585
R233 B.n762 B.n54 585
R234 B.n730 B.n729 585
R235 B.n729 B.n50 585
R236 B.n728 B.n49 585
R237 B.n768 B.n49 585
R238 B.n727 B.n48 585
R239 B.n769 B.n48 585
R240 B.n726 B.n47 585
R241 B.n770 B.n47 585
R242 B.n725 B.n724 585
R243 B.n724 B.n43 585
R244 B.n723 B.n42 585
R245 B.n776 B.n42 585
R246 B.n722 B.n41 585
R247 B.n777 B.n41 585
R248 B.n721 B.n40 585
R249 B.n778 B.n40 585
R250 B.n720 B.n719 585
R251 B.n719 B.n36 585
R252 B.n718 B.n35 585
R253 B.n784 B.n35 585
R254 B.n717 B.n34 585
R255 B.n785 B.n34 585
R256 B.n716 B.n33 585
R257 B.n786 B.n33 585
R258 B.n715 B.n714 585
R259 B.n714 B.n29 585
R260 B.n713 B.n28 585
R261 B.n792 B.n28 585
R262 B.n712 B.n27 585
R263 B.n793 B.n27 585
R264 B.n711 B.n26 585
R265 B.n794 B.n26 585
R266 B.n710 B.n709 585
R267 B.n709 B.n22 585
R268 B.n708 B.n21 585
R269 B.n800 B.n21 585
R270 B.n707 B.n20 585
R271 B.n801 B.n20 585
R272 B.n706 B.n19 585
R273 B.n802 B.n19 585
R274 B.n705 B.n704 585
R275 B.n704 B.n15 585
R276 B.n703 B.n14 585
R277 B.n808 B.n14 585
R278 B.n702 B.n13 585
R279 B.n809 B.n13 585
R280 B.n701 B.n12 585
R281 B.n810 B.n12 585
R282 B.n700 B.n699 585
R283 B.n699 B.n698 585
R284 B.n697 B.n696 585
R285 B.n697 B.n8 585
R286 B.n695 B.n7 585
R287 B.n817 B.n7 585
R288 B.n694 B.n6 585
R289 B.n818 B.n6 585
R290 B.n693 B.n5 585
R291 B.n819 B.n5 585
R292 B.n692 B.n691 585
R293 B.n691 B.n4 585
R294 B.n690 B.n290 585
R295 B.n690 B.n689 585
R296 B.n680 B.n291 585
R297 B.n292 B.n291 585
R298 B.n682 B.n681 585
R299 B.n683 B.n682 585
R300 B.n679 B.n297 585
R301 B.n297 B.n296 585
R302 B.n678 B.n677 585
R303 B.n677 B.n676 585
R304 B.n299 B.n298 585
R305 B.n300 B.n299 585
R306 B.n669 B.n668 585
R307 B.n670 B.n669 585
R308 B.n667 B.n305 585
R309 B.n305 B.n304 585
R310 B.n666 B.n665 585
R311 B.n665 B.n664 585
R312 B.n307 B.n306 585
R313 B.n308 B.n307 585
R314 B.n657 B.n656 585
R315 B.n658 B.n657 585
R316 B.n655 B.n313 585
R317 B.n313 B.n312 585
R318 B.n654 B.n653 585
R319 B.n653 B.n652 585
R320 B.n315 B.n314 585
R321 B.n316 B.n315 585
R322 B.n645 B.n644 585
R323 B.n646 B.n645 585
R324 B.n643 B.n321 585
R325 B.n321 B.n320 585
R326 B.n642 B.n641 585
R327 B.n641 B.n640 585
R328 B.n323 B.n322 585
R329 B.n324 B.n323 585
R330 B.n633 B.n632 585
R331 B.n634 B.n633 585
R332 B.n631 B.n328 585
R333 B.n332 B.n328 585
R334 B.n630 B.n629 585
R335 B.n629 B.n628 585
R336 B.n330 B.n329 585
R337 B.n331 B.n330 585
R338 B.n621 B.n620 585
R339 B.n622 B.n621 585
R340 B.n619 B.n337 585
R341 B.n337 B.n336 585
R342 B.n618 B.n617 585
R343 B.n617 B.n616 585
R344 B.n339 B.n338 585
R345 B.n340 B.n339 585
R346 B.n609 B.n608 585
R347 B.n610 B.n609 585
R348 B.n607 B.n345 585
R349 B.n345 B.n344 585
R350 B.n606 B.n605 585
R351 B.n605 B.n604 585
R352 B.n347 B.n346 585
R353 B.n348 B.n347 585
R354 B.n597 B.n596 585
R355 B.n598 B.n597 585
R356 B.n595 B.n353 585
R357 B.n353 B.n352 585
R358 B.n594 B.n593 585
R359 B.n593 B.n592 585
R360 B.n355 B.n354 585
R361 B.n356 B.n355 585
R362 B.n585 B.n584 585
R363 B.n586 B.n585 585
R364 B.n359 B.n358 585
R365 B.n412 B.n411 585
R366 B.n413 B.n409 585
R367 B.n409 B.n360 585
R368 B.n415 B.n414 585
R369 B.n417 B.n408 585
R370 B.n420 B.n419 585
R371 B.n421 B.n407 585
R372 B.n423 B.n422 585
R373 B.n425 B.n406 585
R374 B.n428 B.n427 585
R375 B.n429 B.n405 585
R376 B.n431 B.n430 585
R377 B.n433 B.n404 585
R378 B.n436 B.n435 585
R379 B.n437 B.n403 585
R380 B.n439 B.n438 585
R381 B.n441 B.n402 585
R382 B.n444 B.n443 585
R383 B.n445 B.n401 585
R384 B.n447 B.n446 585
R385 B.n449 B.n400 585
R386 B.n452 B.n451 585
R387 B.n453 B.n399 585
R388 B.n455 B.n454 585
R389 B.n457 B.n398 585
R390 B.n460 B.n459 585
R391 B.n461 B.n397 585
R392 B.n463 B.n462 585
R393 B.n465 B.n396 585
R394 B.n468 B.n467 585
R395 B.n469 B.n395 585
R396 B.n471 B.n470 585
R397 B.n473 B.n394 585
R398 B.n476 B.n475 585
R399 B.n477 B.n393 585
R400 B.n479 B.n478 585
R401 B.n481 B.n392 585
R402 B.n484 B.n483 585
R403 B.n485 B.n389 585
R404 B.n488 B.n487 585
R405 B.n490 B.n388 585
R406 B.n493 B.n492 585
R407 B.n494 B.n387 585
R408 B.n496 B.n495 585
R409 B.n498 B.n386 585
R410 B.n501 B.n500 585
R411 B.n502 B.n385 585
R412 B.n504 B.n503 585
R413 B.n506 B.n384 585
R414 B.n509 B.n508 585
R415 B.n510 B.n380 585
R416 B.n512 B.n511 585
R417 B.n514 B.n379 585
R418 B.n517 B.n516 585
R419 B.n518 B.n378 585
R420 B.n520 B.n519 585
R421 B.n522 B.n377 585
R422 B.n525 B.n524 585
R423 B.n526 B.n376 585
R424 B.n528 B.n527 585
R425 B.n530 B.n375 585
R426 B.n533 B.n532 585
R427 B.n534 B.n374 585
R428 B.n536 B.n535 585
R429 B.n538 B.n373 585
R430 B.n541 B.n540 585
R431 B.n542 B.n372 585
R432 B.n544 B.n543 585
R433 B.n546 B.n371 585
R434 B.n549 B.n548 585
R435 B.n550 B.n370 585
R436 B.n552 B.n551 585
R437 B.n554 B.n369 585
R438 B.n557 B.n556 585
R439 B.n558 B.n368 585
R440 B.n560 B.n559 585
R441 B.n562 B.n367 585
R442 B.n565 B.n564 585
R443 B.n566 B.n366 585
R444 B.n568 B.n567 585
R445 B.n570 B.n365 585
R446 B.n573 B.n572 585
R447 B.n574 B.n364 585
R448 B.n576 B.n575 585
R449 B.n578 B.n363 585
R450 B.n579 B.n362 585
R451 B.n582 B.n581 585
R452 B.n583 B.n361 585
R453 B.n361 B.n360 585
R454 B.n588 B.n587 585
R455 B.n587 B.n586 585
R456 B.n589 B.n357 585
R457 B.n357 B.n356 585
R458 B.n591 B.n590 585
R459 B.n592 B.n591 585
R460 B.n351 B.n350 585
R461 B.n352 B.n351 585
R462 B.n600 B.n599 585
R463 B.n599 B.n598 585
R464 B.n601 B.n349 585
R465 B.n349 B.n348 585
R466 B.n603 B.n602 585
R467 B.n604 B.n603 585
R468 B.n343 B.n342 585
R469 B.n344 B.n343 585
R470 B.n612 B.n611 585
R471 B.n611 B.n610 585
R472 B.n613 B.n341 585
R473 B.n341 B.n340 585
R474 B.n615 B.n614 585
R475 B.n616 B.n615 585
R476 B.n335 B.n334 585
R477 B.n336 B.n335 585
R478 B.n624 B.n623 585
R479 B.n623 B.n622 585
R480 B.n625 B.n333 585
R481 B.n333 B.n331 585
R482 B.n627 B.n626 585
R483 B.n628 B.n627 585
R484 B.n327 B.n326 585
R485 B.n332 B.n327 585
R486 B.n636 B.n635 585
R487 B.n635 B.n634 585
R488 B.n637 B.n325 585
R489 B.n325 B.n324 585
R490 B.n639 B.n638 585
R491 B.n640 B.n639 585
R492 B.n319 B.n318 585
R493 B.n320 B.n319 585
R494 B.n648 B.n647 585
R495 B.n647 B.n646 585
R496 B.n649 B.n317 585
R497 B.n317 B.n316 585
R498 B.n651 B.n650 585
R499 B.n652 B.n651 585
R500 B.n311 B.n310 585
R501 B.n312 B.n311 585
R502 B.n660 B.n659 585
R503 B.n659 B.n658 585
R504 B.n661 B.n309 585
R505 B.n309 B.n308 585
R506 B.n663 B.n662 585
R507 B.n664 B.n663 585
R508 B.n303 B.n302 585
R509 B.n304 B.n303 585
R510 B.n672 B.n671 585
R511 B.n671 B.n670 585
R512 B.n673 B.n301 585
R513 B.n301 B.n300 585
R514 B.n675 B.n674 585
R515 B.n676 B.n675 585
R516 B.n295 B.n294 585
R517 B.n296 B.n295 585
R518 B.n685 B.n684 585
R519 B.n684 B.n683 585
R520 B.n686 B.n293 585
R521 B.n293 B.n292 585
R522 B.n688 B.n687 585
R523 B.n689 B.n688 585
R524 B.n3 B.n0 585
R525 B.n4 B.n3 585
R526 B.n816 B.n1 585
R527 B.n817 B.n816 585
R528 B.n815 B.n814 585
R529 B.n815 B.n8 585
R530 B.n813 B.n9 585
R531 B.n698 B.n9 585
R532 B.n812 B.n811 585
R533 B.n811 B.n810 585
R534 B.n11 B.n10 585
R535 B.n809 B.n11 585
R536 B.n807 B.n806 585
R537 B.n808 B.n807 585
R538 B.n805 B.n16 585
R539 B.n16 B.n15 585
R540 B.n804 B.n803 585
R541 B.n803 B.n802 585
R542 B.n18 B.n17 585
R543 B.n801 B.n18 585
R544 B.n799 B.n798 585
R545 B.n800 B.n799 585
R546 B.n797 B.n23 585
R547 B.n23 B.n22 585
R548 B.n796 B.n795 585
R549 B.n795 B.n794 585
R550 B.n25 B.n24 585
R551 B.n793 B.n25 585
R552 B.n791 B.n790 585
R553 B.n792 B.n791 585
R554 B.n789 B.n30 585
R555 B.n30 B.n29 585
R556 B.n788 B.n787 585
R557 B.n787 B.n786 585
R558 B.n32 B.n31 585
R559 B.n785 B.n32 585
R560 B.n783 B.n782 585
R561 B.n784 B.n783 585
R562 B.n781 B.n37 585
R563 B.n37 B.n36 585
R564 B.n780 B.n779 585
R565 B.n779 B.n778 585
R566 B.n39 B.n38 585
R567 B.n777 B.n39 585
R568 B.n775 B.n774 585
R569 B.n776 B.n775 585
R570 B.n773 B.n44 585
R571 B.n44 B.n43 585
R572 B.n772 B.n771 585
R573 B.n771 B.n770 585
R574 B.n46 B.n45 585
R575 B.n769 B.n46 585
R576 B.n767 B.n766 585
R577 B.n768 B.n767 585
R578 B.n765 B.n51 585
R579 B.n51 B.n50 585
R580 B.n764 B.n763 585
R581 B.n763 B.n762 585
R582 B.n53 B.n52 585
R583 B.n761 B.n53 585
R584 B.n759 B.n758 585
R585 B.n760 B.n759 585
R586 B.n757 B.n58 585
R587 B.n58 B.n57 585
R588 B.n756 B.n755 585
R589 B.n755 B.n754 585
R590 B.n60 B.n59 585
R591 B.n753 B.n60 585
R592 B.n751 B.n750 585
R593 B.n752 B.n751 585
R594 B.n749 B.n65 585
R595 B.n65 B.n64 585
R596 B.n748 B.n747 585
R597 B.n747 B.n746 585
R598 B.n820 B.n819 585
R599 B.n818 B.n2 585
R600 B.n747 B.n67 482.89
R601 B.n743 B.n68 482.89
R602 B.n585 B.n361 482.89
R603 B.n587 B.n359 482.89
R604 B.n115 B.t19 375.522
R605 B.n113 B.t12 375.522
R606 B.n381 B.t8 375.522
R607 B.n390 B.t16 375.522
R608 B.n745 B.n744 256.663
R609 B.n745 B.n111 256.663
R610 B.n745 B.n110 256.663
R611 B.n745 B.n109 256.663
R612 B.n745 B.n108 256.663
R613 B.n745 B.n107 256.663
R614 B.n745 B.n106 256.663
R615 B.n745 B.n105 256.663
R616 B.n745 B.n104 256.663
R617 B.n745 B.n103 256.663
R618 B.n745 B.n102 256.663
R619 B.n745 B.n101 256.663
R620 B.n745 B.n100 256.663
R621 B.n745 B.n99 256.663
R622 B.n745 B.n98 256.663
R623 B.n745 B.n97 256.663
R624 B.n745 B.n96 256.663
R625 B.n745 B.n95 256.663
R626 B.n745 B.n94 256.663
R627 B.n745 B.n93 256.663
R628 B.n745 B.n92 256.663
R629 B.n745 B.n91 256.663
R630 B.n745 B.n90 256.663
R631 B.n745 B.n89 256.663
R632 B.n745 B.n88 256.663
R633 B.n745 B.n87 256.663
R634 B.n745 B.n86 256.663
R635 B.n745 B.n85 256.663
R636 B.n745 B.n84 256.663
R637 B.n745 B.n83 256.663
R638 B.n745 B.n82 256.663
R639 B.n745 B.n81 256.663
R640 B.n745 B.n80 256.663
R641 B.n745 B.n79 256.663
R642 B.n745 B.n78 256.663
R643 B.n745 B.n77 256.663
R644 B.n745 B.n76 256.663
R645 B.n745 B.n75 256.663
R646 B.n745 B.n74 256.663
R647 B.n745 B.n73 256.663
R648 B.n745 B.n72 256.663
R649 B.n745 B.n71 256.663
R650 B.n745 B.n70 256.663
R651 B.n745 B.n69 256.663
R652 B.n410 B.n360 256.663
R653 B.n416 B.n360 256.663
R654 B.n418 B.n360 256.663
R655 B.n424 B.n360 256.663
R656 B.n426 B.n360 256.663
R657 B.n432 B.n360 256.663
R658 B.n434 B.n360 256.663
R659 B.n440 B.n360 256.663
R660 B.n442 B.n360 256.663
R661 B.n448 B.n360 256.663
R662 B.n450 B.n360 256.663
R663 B.n456 B.n360 256.663
R664 B.n458 B.n360 256.663
R665 B.n464 B.n360 256.663
R666 B.n466 B.n360 256.663
R667 B.n472 B.n360 256.663
R668 B.n474 B.n360 256.663
R669 B.n480 B.n360 256.663
R670 B.n482 B.n360 256.663
R671 B.n489 B.n360 256.663
R672 B.n491 B.n360 256.663
R673 B.n497 B.n360 256.663
R674 B.n499 B.n360 256.663
R675 B.n505 B.n360 256.663
R676 B.n507 B.n360 256.663
R677 B.n513 B.n360 256.663
R678 B.n515 B.n360 256.663
R679 B.n521 B.n360 256.663
R680 B.n523 B.n360 256.663
R681 B.n529 B.n360 256.663
R682 B.n531 B.n360 256.663
R683 B.n537 B.n360 256.663
R684 B.n539 B.n360 256.663
R685 B.n545 B.n360 256.663
R686 B.n547 B.n360 256.663
R687 B.n553 B.n360 256.663
R688 B.n555 B.n360 256.663
R689 B.n561 B.n360 256.663
R690 B.n563 B.n360 256.663
R691 B.n569 B.n360 256.663
R692 B.n571 B.n360 256.663
R693 B.n577 B.n360 256.663
R694 B.n580 B.n360 256.663
R695 B.n822 B.n821 256.663
R696 B.n119 B.n118 163.367
R697 B.n123 B.n122 163.367
R698 B.n127 B.n126 163.367
R699 B.n131 B.n130 163.367
R700 B.n135 B.n134 163.367
R701 B.n139 B.n138 163.367
R702 B.n143 B.n142 163.367
R703 B.n147 B.n146 163.367
R704 B.n151 B.n150 163.367
R705 B.n155 B.n154 163.367
R706 B.n159 B.n158 163.367
R707 B.n163 B.n162 163.367
R708 B.n167 B.n166 163.367
R709 B.n171 B.n170 163.367
R710 B.n175 B.n174 163.367
R711 B.n179 B.n178 163.367
R712 B.n183 B.n182 163.367
R713 B.n187 B.n186 163.367
R714 B.n191 B.n190 163.367
R715 B.n196 B.n195 163.367
R716 B.n200 B.n199 163.367
R717 B.n204 B.n203 163.367
R718 B.n208 B.n207 163.367
R719 B.n212 B.n211 163.367
R720 B.n217 B.n216 163.367
R721 B.n221 B.n220 163.367
R722 B.n225 B.n224 163.367
R723 B.n229 B.n228 163.367
R724 B.n233 B.n232 163.367
R725 B.n237 B.n236 163.367
R726 B.n241 B.n240 163.367
R727 B.n245 B.n244 163.367
R728 B.n249 B.n248 163.367
R729 B.n253 B.n252 163.367
R730 B.n257 B.n256 163.367
R731 B.n261 B.n260 163.367
R732 B.n265 B.n264 163.367
R733 B.n269 B.n268 163.367
R734 B.n273 B.n272 163.367
R735 B.n277 B.n276 163.367
R736 B.n281 B.n280 163.367
R737 B.n285 B.n284 163.367
R738 B.n287 B.n112 163.367
R739 B.n585 B.n355 163.367
R740 B.n593 B.n355 163.367
R741 B.n593 B.n353 163.367
R742 B.n597 B.n353 163.367
R743 B.n597 B.n347 163.367
R744 B.n605 B.n347 163.367
R745 B.n605 B.n345 163.367
R746 B.n609 B.n345 163.367
R747 B.n609 B.n339 163.367
R748 B.n617 B.n339 163.367
R749 B.n617 B.n337 163.367
R750 B.n621 B.n337 163.367
R751 B.n621 B.n330 163.367
R752 B.n629 B.n330 163.367
R753 B.n629 B.n328 163.367
R754 B.n633 B.n328 163.367
R755 B.n633 B.n323 163.367
R756 B.n641 B.n323 163.367
R757 B.n641 B.n321 163.367
R758 B.n645 B.n321 163.367
R759 B.n645 B.n315 163.367
R760 B.n653 B.n315 163.367
R761 B.n653 B.n313 163.367
R762 B.n657 B.n313 163.367
R763 B.n657 B.n307 163.367
R764 B.n665 B.n307 163.367
R765 B.n665 B.n305 163.367
R766 B.n669 B.n305 163.367
R767 B.n669 B.n299 163.367
R768 B.n677 B.n299 163.367
R769 B.n677 B.n297 163.367
R770 B.n682 B.n297 163.367
R771 B.n682 B.n291 163.367
R772 B.n690 B.n291 163.367
R773 B.n691 B.n690 163.367
R774 B.n691 B.n5 163.367
R775 B.n6 B.n5 163.367
R776 B.n7 B.n6 163.367
R777 B.n697 B.n7 163.367
R778 B.n699 B.n697 163.367
R779 B.n699 B.n12 163.367
R780 B.n13 B.n12 163.367
R781 B.n14 B.n13 163.367
R782 B.n704 B.n14 163.367
R783 B.n704 B.n19 163.367
R784 B.n20 B.n19 163.367
R785 B.n21 B.n20 163.367
R786 B.n709 B.n21 163.367
R787 B.n709 B.n26 163.367
R788 B.n27 B.n26 163.367
R789 B.n28 B.n27 163.367
R790 B.n714 B.n28 163.367
R791 B.n714 B.n33 163.367
R792 B.n34 B.n33 163.367
R793 B.n35 B.n34 163.367
R794 B.n719 B.n35 163.367
R795 B.n719 B.n40 163.367
R796 B.n41 B.n40 163.367
R797 B.n42 B.n41 163.367
R798 B.n724 B.n42 163.367
R799 B.n724 B.n47 163.367
R800 B.n48 B.n47 163.367
R801 B.n49 B.n48 163.367
R802 B.n729 B.n49 163.367
R803 B.n729 B.n54 163.367
R804 B.n55 B.n54 163.367
R805 B.n56 B.n55 163.367
R806 B.n734 B.n56 163.367
R807 B.n734 B.n61 163.367
R808 B.n62 B.n61 163.367
R809 B.n63 B.n62 163.367
R810 B.n739 B.n63 163.367
R811 B.n739 B.n68 163.367
R812 B.n411 B.n409 163.367
R813 B.n415 B.n409 163.367
R814 B.n419 B.n417 163.367
R815 B.n423 B.n407 163.367
R816 B.n427 B.n425 163.367
R817 B.n431 B.n405 163.367
R818 B.n435 B.n433 163.367
R819 B.n439 B.n403 163.367
R820 B.n443 B.n441 163.367
R821 B.n447 B.n401 163.367
R822 B.n451 B.n449 163.367
R823 B.n455 B.n399 163.367
R824 B.n459 B.n457 163.367
R825 B.n463 B.n397 163.367
R826 B.n467 B.n465 163.367
R827 B.n471 B.n395 163.367
R828 B.n475 B.n473 163.367
R829 B.n479 B.n393 163.367
R830 B.n483 B.n481 163.367
R831 B.n488 B.n389 163.367
R832 B.n492 B.n490 163.367
R833 B.n496 B.n387 163.367
R834 B.n500 B.n498 163.367
R835 B.n504 B.n385 163.367
R836 B.n508 B.n506 163.367
R837 B.n512 B.n380 163.367
R838 B.n516 B.n514 163.367
R839 B.n520 B.n378 163.367
R840 B.n524 B.n522 163.367
R841 B.n528 B.n376 163.367
R842 B.n532 B.n530 163.367
R843 B.n536 B.n374 163.367
R844 B.n540 B.n538 163.367
R845 B.n544 B.n372 163.367
R846 B.n548 B.n546 163.367
R847 B.n552 B.n370 163.367
R848 B.n556 B.n554 163.367
R849 B.n560 B.n368 163.367
R850 B.n564 B.n562 163.367
R851 B.n568 B.n366 163.367
R852 B.n572 B.n570 163.367
R853 B.n576 B.n364 163.367
R854 B.n579 B.n578 163.367
R855 B.n581 B.n361 163.367
R856 B.n587 B.n357 163.367
R857 B.n591 B.n357 163.367
R858 B.n591 B.n351 163.367
R859 B.n599 B.n351 163.367
R860 B.n599 B.n349 163.367
R861 B.n603 B.n349 163.367
R862 B.n603 B.n343 163.367
R863 B.n611 B.n343 163.367
R864 B.n611 B.n341 163.367
R865 B.n615 B.n341 163.367
R866 B.n615 B.n335 163.367
R867 B.n623 B.n335 163.367
R868 B.n623 B.n333 163.367
R869 B.n627 B.n333 163.367
R870 B.n627 B.n327 163.367
R871 B.n635 B.n327 163.367
R872 B.n635 B.n325 163.367
R873 B.n639 B.n325 163.367
R874 B.n639 B.n319 163.367
R875 B.n647 B.n319 163.367
R876 B.n647 B.n317 163.367
R877 B.n651 B.n317 163.367
R878 B.n651 B.n311 163.367
R879 B.n659 B.n311 163.367
R880 B.n659 B.n309 163.367
R881 B.n663 B.n309 163.367
R882 B.n663 B.n303 163.367
R883 B.n671 B.n303 163.367
R884 B.n671 B.n301 163.367
R885 B.n675 B.n301 163.367
R886 B.n675 B.n295 163.367
R887 B.n684 B.n295 163.367
R888 B.n684 B.n293 163.367
R889 B.n688 B.n293 163.367
R890 B.n688 B.n3 163.367
R891 B.n820 B.n3 163.367
R892 B.n816 B.n2 163.367
R893 B.n816 B.n815 163.367
R894 B.n815 B.n9 163.367
R895 B.n811 B.n9 163.367
R896 B.n811 B.n11 163.367
R897 B.n807 B.n11 163.367
R898 B.n807 B.n16 163.367
R899 B.n803 B.n16 163.367
R900 B.n803 B.n18 163.367
R901 B.n799 B.n18 163.367
R902 B.n799 B.n23 163.367
R903 B.n795 B.n23 163.367
R904 B.n795 B.n25 163.367
R905 B.n791 B.n25 163.367
R906 B.n791 B.n30 163.367
R907 B.n787 B.n30 163.367
R908 B.n787 B.n32 163.367
R909 B.n783 B.n32 163.367
R910 B.n783 B.n37 163.367
R911 B.n779 B.n37 163.367
R912 B.n779 B.n39 163.367
R913 B.n775 B.n39 163.367
R914 B.n775 B.n44 163.367
R915 B.n771 B.n44 163.367
R916 B.n771 B.n46 163.367
R917 B.n767 B.n46 163.367
R918 B.n767 B.n51 163.367
R919 B.n763 B.n51 163.367
R920 B.n763 B.n53 163.367
R921 B.n759 B.n53 163.367
R922 B.n759 B.n58 163.367
R923 B.n755 B.n58 163.367
R924 B.n755 B.n60 163.367
R925 B.n751 B.n60 163.367
R926 B.n751 B.n65 163.367
R927 B.n747 B.n65 163.367
R928 B.n113 B.t14 111.349
R929 B.n381 B.t11 111.349
R930 B.n115 B.t20 111.335
R931 B.n390 B.t18 111.335
R932 B.n586 B.n360 75.4481
R933 B.n746 B.n745 75.4481
R934 B.n114 B.t15 74.1123
R935 B.n382 B.t10 74.1123
R936 B.n116 B.t21 74.0986
R937 B.n391 B.t17 74.0986
R938 B.n69 B.n67 71.676
R939 B.n119 B.n70 71.676
R940 B.n123 B.n71 71.676
R941 B.n127 B.n72 71.676
R942 B.n131 B.n73 71.676
R943 B.n135 B.n74 71.676
R944 B.n139 B.n75 71.676
R945 B.n143 B.n76 71.676
R946 B.n147 B.n77 71.676
R947 B.n151 B.n78 71.676
R948 B.n155 B.n79 71.676
R949 B.n159 B.n80 71.676
R950 B.n163 B.n81 71.676
R951 B.n167 B.n82 71.676
R952 B.n171 B.n83 71.676
R953 B.n175 B.n84 71.676
R954 B.n179 B.n85 71.676
R955 B.n183 B.n86 71.676
R956 B.n187 B.n87 71.676
R957 B.n191 B.n88 71.676
R958 B.n196 B.n89 71.676
R959 B.n200 B.n90 71.676
R960 B.n204 B.n91 71.676
R961 B.n208 B.n92 71.676
R962 B.n212 B.n93 71.676
R963 B.n217 B.n94 71.676
R964 B.n221 B.n95 71.676
R965 B.n225 B.n96 71.676
R966 B.n229 B.n97 71.676
R967 B.n233 B.n98 71.676
R968 B.n237 B.n99 71.676
R969 B.n241 B.n100 71.676
R970 B.n245 B.n101 71.676
R971 B.n249 B.n102 71.676
R972 B.n253 B.n103 71.676
R973 B.n257 B.n104 71.676
R974 B.n261 B.n105 71.676
R975 B.n265 B.n106 71.676
R976 B.n269 B.n107 71.676
R977 B.n273 B.n108 71.676
R978 B.n277 B.n109 71.676
R979 B.n281 B.n110 71.676
R980 B.n285 B.n111 71.676
R981 B.n744 B.n112 71.676
R982 B.n744 B.n743 71.676
R983 B.n287 B.n111 71.676
R984 B.n284 B.n110 71.676
R985 B.n280 B.n109 71.676
R986 B.n276 B.n108 71.676
R987 B.n272 B.n107 71.676
R988 B.n268 B.n106 71.676
R989 B.n264 B.n105 71.676
R990 B.n260 B.n104 71.676
R991 B.n256 B.n103 71.676
R992 B.n252 B.n102 71.676
R993 B.n248 B.n101 71.676
R994 B.n244 B.n100 71.676
R995 B.n240 B.n99 71.676
R996 B.n236 B.n98 71.676
R997 B.n232 B.n97 71.676
R998 B.n228 B.n96 71.676
R999 B.n224 B.n95 71.676
R1000 B.n220 B.n94 71.676
R1001 B.n216 B.n93 71.676
R1002 B.n211 B.n92 71.676
R1003 B.n207 B.n91 71.676
R1004 B.n203 B.n90 71.676
R1005 B.n199 B.n89 71.676
R1006 B.n195 B.n88 71.676
R1007 B.n190 B.n87 71.676
R1008 B.n186 B.n86 71.676
R1009 B.n182 B.n85 71.676
R1010 B.n178 B.n84 71.676
R1011 B.n174 B.n83 71.676
R1012 B.n170 B.n82 71.676
R1013 B.n166 B.n81 71.676
R1014 B.n162 B.n80 71.676
R1015 B.n158 B.n79 71.676
R1016 B.n154 B.n78 71.676
R1017 B.n150 B.n77 71.676
R1018 B.n146 B.n76 71.676
R1019 B.n142 B.n75 71.676
R1020 B.n138 B.n74 71.676
R1021 B.n134 B.n73 71.676
R1022 B.n130 B.n72 71.676
R1023 B.n126 B.n71 71.676
R1024 B.n122 B.n70 71.676
R1025 B.n118 B.n69 71.676
R1026 B.n410 B.n359 71.676
R1027 B.n416 B.n415 71.676
R1028 B.n419 B.n418 71.676
R1029 B.n424 B.n423 71.676
R1030 B.n427 B.n426 71.676
R1031 B.n432 B.n431 71.676
R1032 B.n435 B.n434 71.676
R1033 B.n440 B.n439 71.676
R1034 B.n443 B.n442 71.676
R1035 B.n448 B.n447 71.676
R1036 B.n451 B.n450 71.676
R1037 B.n456 B.n455 71.676
R1038 B.n459 B.n458 71.676
R1039 B.n464 B.n463 71.676
R1040 B.n467 B.n466 71.676
R1041 B.n472 B.n471 71.676
R1042 B.n475 B.n474 71.676
R1043 B.n480 B.n479 71.676
R1044 B.n483 B.n482 71.676
R1045 B.n489 B.n488 71.676
R1046 B.n492 B.n491 71.676
R1047 B.n497 B.n496 71.676
R1048 B.n500 B.n499 71.676
R1049 B.n505 B.n504 71.676
R1050 B.n508 B.n507 71.676
R1051 B.n513 B.n512 71.676
R1052 B.n516 B.n515 71.676
R1053 B.n521 B.n520 71.676
R1054 B.n524 B.n523 71.676
R1055 B.n529 B.n528 71.676
R1056 B.n532 B.n531 71.676
R1057 B.n537 B.n536 71.676
R1058 B.n540 B.n539 71.676
R1059 B.n545 B.n544 71.676
R1060 B.n548 B.n547 71.676
R1061 B.n553 B.n552 71.676
R1062 B.n556 B.n555 71.676
R1063 B.n561 B.n560 71.676
R1064 B.n564 B.n563 71.676
R1065 B.n569 B.n568 71.676
R1066 B.n572 B.n571 71.676
R1067 B.n577 B.n576 71.676
R1068 B.n580 B.n579 71.676
R1069 B.n411 B.n410 71.676
R1070 B.n417 B.n416 71.676
R1071 B.n418 B.n407 71.676
R1072 B.n425 B.n424 71.676
R1073 B.n426 B.n405 71.676
R1074 B.n433 B.n432 71.676
R1075 B.n434 B.n403 71.676
R1076 B.n441 B.n440 71.676
R1077 B.n442 B.n401 71.676
R1078 B.n449 B.n448 71.676
R1079 B.n450 B.n399 71.676
R1080 B.n457 B.n456 71.676
R1081 B.n458 B.n397 71.676
R1082 B.n465 B.n464 71.676
R1083 B.n466 B.n395 71.676
R1084 B.n473 B.n472 71.676
R1085 B.n474 B.n393 71.676
R1086 B.n481 B.n480 71.676
R1087 B.n482 B.n389 71.676
R1088 B.n490 B.n489 71.676
R1089 B.n491 B.n387 71.676
R1090 B.n498 B.n497 71.676
R1091 B.n499 B.n385 71.676
R1092 B.n506 B.n505 71.676
R1093 B.n507 B.n380 71.676
R1094 B.n514 B.n513 71.676
R1095 B.n515 B.n378 71.676
R1096 B.n522 B.n521 71.676
R1097 B.n523 B.n376 71.676
R1098 B.n530 B.n529 71.676
R1099 B.n531 B.n374 71.676
R1100 B.n538 B.n537 71.676
R1101 B.n539 B.n372 71.676
R1102 B.n546 B.n545 71.676
R1103 B.n547 B.n370 71.676
R1104 B.n554 B.n553 71.676
R1105 B.n555 B.n368 71.676
R1106 B.n562 B.n561 71.676
R1107 B.n563 B.n366 71.676
R1108 B.n570 B.n569 71.676
R1109 B.n571 B.n364 71.676
R1110 B.n578 B.n577 71.676
R1111 B.n581 B.n580 71.676
R1112 B.n821 B.n820 71.676
R1113 B.n821 B.n2 71.676
R1114 B.n193 B.n116 59.5399
R1115 B.n214 B.n114 59.5399
R1116 B.n383 B.n382 59.5399
R1117 B.n486 B.n391 59.5399
R1118 B.n586 B.n356 45.4026
R1119 B.n592 B.n356 45.4026
R1120 B.n592 B.n352 45.4026
R1121 B.n598 B.n352 45.4026
R1122 B.n598 B.n348 45.4026
R1123 B.n604 B.n348 45.4026
R1124 B.n610 B.n344 45.4026
R1125 B.n610 B.n340 45.4026
R1126 B.n616 B.n340 45.4026
R1127 B.n616 B.n336 45.4026
R1128 B.n622 B.n336 45.4026
R1129 B.n622 B.n331 45.4026
R1130 B.n628 B.n331 45.4026
R1131 B.n628 B.n332 45.4026
R1132 B.n634 B.n324 45.4026
R1133 B.n640 B.n324 45.4026
R1134 B.n640 B.n320 45.4026
R1135 B.n646 B.n320 45.4026
R1136 B.n652 B.n316 45.4026
R1137 B.n652 B.n312 45.4026
R1138 B.n658 B.n312 45.4026
R1139 B.n658 B.n308 45.4026
R1140 B.n664 B.n308 45.4026
R1141 B.n670 B.n304 45.4026
R1142 B.n670 B.n300 45.4026
R1143 B.n676 B.n300 45.4026
R1144 B.n676 B.n296 45.4026
R1145 B.n683 B.n296 45.4026
R1146 B.n689 B.n292 45.4026
R1147 B.n689 B.n4 45.4026
R1148 B.n819 B.n4 45.4026
R1149 B.n819 B.n818 45.4026
R1150 B.n818 B.n817 45.4026
R1151 B.n817 B.n8 45.4026
R1152 B.n698 B.n8 45.4026
R1153 B.n810 B.n809 45.4026
R1154 B.n809 B.n808 45.4026
R1155 B.n808 B.n15 45.4026
R1156 B.n802 B.n15 45.4026
R1157 B.n802 B.n801 45.4026
R1158 B.n800 B.n22 45.4026
R1159 B.n794 B.n22 45.4026
R1160 B.n794 B.n793 45.4026
R1161 B.n793 B.n792 45.4026
R1162 B.n792 B.n29 45.4026
R1163 B.n786 B.n785 45.4026
R1164 B.n785 B.n784 45.4026
R1165 B.n784 B.n36 45.4026
R1166 B.n778 B.n36 45.4026
R1167 B.n777 B.n776 45.4026
R1168 B.n776 B.n43 45.4026
R1169 B.n770 B.n43 45.4026
R1170 B.n770 B.n769 45.4026
R1171 B.n769 B.n768 45.4026
R1172 B.n768 B.n50 45.4026
R1173 B.n762 B.n50 45.4026
R1174 B.n762 B.n761 45.4026
R1175 B.n760 B.n57 45.4026
R1176 B.n754 B.n57 45.4026
R1177 B.n754 B.n753 45.4026
R1178 B.n753 B.n752 45.4026
R1179 B.n752 B.n64 45.4026
R1180 B.n746 B.n64 45.4026
R1181 B.t6 B.n292 42.0642
R1182 B.n698 B.t3 42.0642
R1183 B.n634 B.t0 39.3935
R1184 B.n778 B.t7 39.3935
R1185 B.n116 B.n115 37.2369
R1186 B.n114 B.n113 37.2369
R1187 B.n382 B.n381 37.2369
R1188 B.n391 B.n390 37.2369
R1189 B.n646 B.t5 35.3874
R1190 B.n786 B.t4 35.3874
R1191 B.t9 B.n344 32.7167
R1192 B.n761 B.t13 32.7167
R1193 B.n588 B.n358 31.3761
R1194 B.n584 B.n583 31.3761
R1195 B.n742 B.n741 31.3761
R1196 B.n748 B.n66 31.3761
R1197 B.t2 B.n304 26.04
R1198 B.n801 B.t1 26.04
R1199 B.n664 B.t2 19.3632
R1200 B.t1 B.n800 19.3632
R1201 B B.n822 18.0485
R1202 B.n604 B.t9 12.6864
R1203 B.t13 B.n760 12.6864
R1204 B.n589 B.n588 10.6151
R1205 B.n590 B.n589 10.6151
R1206 B.n590 B.n350 10.6151
R1207 B.n600 B.n350 10.6151
R1208 B.n601 B.n600 10.6151
R1209 B.n602 B.n601 10.6151
R1210 B.n602 B.n342 10.6151
R1211 B.n612 B.n342 10.6151
R1212 B.n613 B.n612 10.6151
R1213 B.n614 B.n613 10.6151
R1214 B.n614 B.n334 10.6151
R1215 B.n624 B.n334 10.6151
R1216 B.n625 B.n624 10.6151
R1217 B.n626 B.n625 10.6151
R1218 B.n626 B.n326 10.6151
R1219 B.n636 B.n326 10.6151
R1220 B.n637 B.n636 10.6151
R1221 B.n638 B.n637 10.6151
R1222 B.n638 B.n318 10.6151
R1223 B.n648 B.n318 10.6151
R1224 B.n649 B.n648 10.6151
R1225 B.n650 B.n649 10.6151
R1226 B.n650 B.n310 10.6151
R1227 B.n660 B.n310 10.6151
R1228 B.n661 B.n660 10.6151
R1229 B.n662 B.n661 10.6151
R1230 B.n662 B.n302 10.6151
R1231 B.n672 B.n302 10.6151
R1232 B.n673 B.n672 10.6151
R1233 B.n674 B.n673 10.6151
R1234 B.n674 B.n294 10.6151
R1235 B.n685 B.n294 10.6151
R1236 B.n686 B.n685 10.6151
R1237 B.n687 B.n686 10.6151
R1238 B.n687 B.n0 10.6151
R1239 B.n412 B.n358 10.6151
R1240 B.n413 B.n412 10.6151
R1241 B.n414 B.n413 10.6151
R1242 B.n414 B.n408 10.6151
R1243 B.n420 B.n408 10.6151
R1244 B.n421 B.n420 10.6151
R1245 B.n422 B.n421 10.6151
R1246 B.n422 B.n406 10.6151
R1247 B.n428 B.n406 10.6151
R1248 B.n429 B.n428 10.6151
R1249 B.n430 B.n429 10.6151
R1250 B.n430 B.n404 10.6151
R1251 B.n436 B.n404 10.6151
R1252 B.n437 B.n436 10.6151
R1253 B.n438 B.n437 10.6151
R1254 B.n438 B.n402 10.6151
R1255 B.n444 B.n402 10.6151
R1256 B.n445 B.n444 10.6151
R1257 B.n446 B.n445 10.6151
R1258 B.n446 B.n400 10.6151
R1259 B.n452 B.n400 10.6151
R1260 B.n453 B.n452 10.6151
R1261 B.n454 B.n453 10.6151
R1262 B.n454 B.n398 10.6151
R1263 B.n460 B.n398 10.6151
R1264 B.n461 B.n460 10.6151
R1265 B.n462 B.n461 10.6151
R1266 B.n462 B.n396 10.6151
R1267 B.n468 B.n396 10.6151
R1268 B.n469 B.n468 10.6151
R1269 B.n470 B.n469 10.6151
R1270 B.n470 B.n394 10.6151
R1271 B.n476 B.n394 10.6151
R1272 B.n477 B.n476 10.6151
R1273 B.n478 B.n477 10.6151
R1274 B.n478 B.n392 10.6151
R1275 B.n484 B.n392 10.6151
R1276 B.n485 B.n484 10.6151
R1277 B.n487 B.n388 10.6151
R1278 B.n493 B.n388 10.6151
R1279 B.n494 B.n493 10.6151
R1280 B.n495 B.n494 10.6151
R1281 B.n495 B.n386 10.6151
R1282 B.n501 B.n386 10.6151
R1283 B.n502 B.n501 10.6151
R1284 B.n503 B.n502 10.6151
R1285 B.n503 B.n384 10.6151
R1286 B.n510 B.n509 10.6151
R1287 B.n511 B.n510 10.6151
R1288 B.n511 B.n379 10.6151
R1289 B.n517 B.n379 10.6151
R1290 B.n518 B.n517 10.6151
R1291 B.n519 B.n518 10.6151
R1292 B.n519 B.n377 10.6151
R1293 B.n525 B.n377 10.6151
R1294 B.n526 B.n525 10.6151
R1295 B.n527 B.n526 10.6151
R1296 B.n527 B.n375 10.6151
R1297 B.n533 B.n375 10.6151
R1298 B.n534 B.n533 10.6151
R1299 B.n535 B.n534 10.6151
R1300 B.n535 B.n373 10.6151
R1301 B.n541 B.n373 10.6151
R1302 B.n542 B.n541 10.6151
R1303 B.n543 B.n542 10.6151
R1304 B.n543 B.n371 10.6151
R1305 B.n549 B.n371 10.6151
R1306 B.n550 B.n549 10.6151
R1307 B.n551 B.n550 10.6151
R1308 B.n551 B.n369 10.6151
R1309 B.n557 B.n369 10.6151
R1310 B.n558 B.n557 10.6151
R1311 B.n559 B.n558 10.6151
R1312 B.n559 B.n367 10.6151
R1313 B.n565 B.n367 10.6151
R1314 B.n566 B.n565 10.6151
R1315 B.n567 B.n566 10.6151
R1316 B.n567 B.n365 10.6151
R1317 B.n573 B.n365 10.6151
R1318 B.n574 B.n573 10.6151
R1319 B.n575 B.n574 10.6151
R1320 B.n575 B.n363 10.6151
R1321 B.n363 B.n362 10.6151
R1322 B.n582 B.n362 10.6151
R1323 B.n583 B.n582 10.6151
R1324 B.n584 B.n354 10.6151
R1325 B.n594 B.n354 10.6151
R1326 B.n595 B.n594 10.6151
R1327 B.n596 B.n595 10.6151
R1328 B.n596 B.n346 10.6151
R1329 B.n606 B.n346 10.6151
R1330 B.n607 B.n606 10.6151
R1331 B.n608 B.n607 10.6151
R1332 B.n608 B.n338 10.6151
R1333 B.n618 B.n338 10.6151
R1334 B.n619 B.n618 10.6151
R1335 B.n620 B.n619 10.6151
R1336 B.n620 B.n329 10.6151
R1337 B.n630 B.n329 10.6151
R1338 B.n631 B.n630 10.6151
R1339 B.n632 B.n631 10.6151
R1340 B.n632 B.n322 10.6151
R1341 B.n642 B.n322 10.6151
R1342 B.n643 B.n642 10.6151
R1343 B.n644 B.n643 10.6151
R1344 B.n644 B.n314 10.6151
R1345 B.n654 B.n314 10.6151
R1346 B.n655 B.n654 10.6151
R1347 B.n656 B.n655 10.6151
R1348 B.n656 B.n306 10.6151
R1349 B.n666 B.n306 10.6151
R1350 B.n667 B.n666 10.6151
R1351 B.n668 B.n667 10.6151
R1352 B.n668 B.n298 10.6151
R1353 B.n678 B.n298 10.6151
R1354 B.n679 B.n678 10.6151
R1355 B.n681 B.n679 10.6151
R1356 B.n681 B.n680 10.6151
R1357 B.n680 B.n290 10.6151
R1358 B.n692 B.n290 10.6151
R1359 B.n693 B.n692 10.6151
R1360 B.n694 B.n693 10.6151
R1361 B.n695 B.n694 10.6151
R1362 B.n696 B.n695 10.6151
R1363 B.n700 B.n696 10.6151
R1364 B.n701 B.n700 10.6151
R1365 B.n702 B.n701 10.6151
R1366 B.n703 B.n702 10.6151
R1367 B.n705 B.n703 10.6151
R1368 B.n706 B.n705 10.6151
R1369 B.n707 B.n706 10.6151
R1370 B.n708 B.n707 10.6151
R1371 B.n710 B.n708 10.6151
R1372 B.n711 B.n710 10.6151
R1373 B.n712 B.n711 10.6151
R1374 B.n713 B.n712 10.6151
R1375 B.n715 B.n713 10.6151
R1376 B.n716 B.n715 10.6151
R1377 B.n717 B.n716 10.6151
R1378 B.n718 B.n717 10.6151
R1379 B.n720 B.n718 10.6151
R1380 B.n721 B.n720 10.6151
R1381 B.n722 B.n721 10.6151
R1382 B.n723 B.n722 10.6151
R1383 B.n725 B.n723 10.6151
R1384 B.n726 B.n725 10.6151
R1385 B.n727 B.n726 10.6151
R1386 B.n728 B.n727 10.6151
R1387 B.n730 B.n728 10.6151
R1388 B.n731 B.n730 10.6151
R1389 B.n732 B.n731 10.6151
R1390 B.n733 B.n732 10.6151
R1391 B.n735 B.n733 10.6151
R1392 B.n736 B.n735 10.6151
R1393 B.n737 B.n736 10.6151
R1394 B.n738 B.n737 10.6151
R1395 B.n740 B.n738 10.6151
R1396 B.n741 B.n740 10.6151
R1397 B.n814 B.n1 10.6151
R1398 B.n814 B.n813 10.6151
R1399 B.n813 B.n812 10.6151
R1400 B.n812 B.n10 10.6151
R1401 B.n806 B.n10 10.6151
R1402 B.n806 B.n805 10.6151
R1403 B.n805 B.n804 10.6151
R1404 B.n804 B.n17 10.6151
R1405 B.n798 B.n17 10.6151
R1406 B.n798 B.n797 10.6151
R1407 B.n797 B.n796 10.6151
R1408 B.n796 B.n24 10.6151
R1409 B.n790 B.n24 10.6151
R1410 B.n790 B.n789 10.6151
R1411 B.n789 B.n788 10.6151
R1412 B.n788 B.n31 10.6151
R1413 B.n782 B.n31 10.6151
R1414 B.n782 B.n781 10.6151
R1415 B.n781 B.n780 10.6151
R1416 B.n780 B.n38 10.6151
R1417 B.n774 B.n38 10.6151
R1418 B.n774 B.n773 10.6151
R1419 B.n773 B.n772 10.6151
R1420 B.n772 B.n45 10.6151
R1421 B.n766 B.n45 10.6151
R1422 B.n766 B.n765 10.6151
R1423 B.n765 B.n764 10.6151
R1424 B.n764 B.n52 10.6151
R1425 B.n758 B.n52 10.6151
R1426 B.n758 B.n757 10.6151
R1427 B.n757 B.n756 10.6151
R1428 B.n756 B.n59 10.6151
R1429 B.n750 B.n59 10.6151
R1430 B.n750 B.n749 10.6151
R1431 B.n749 B.n748 10.6151
R1432 B.n117 B.n66 10.6151
R1433 B.n120 B.n117 10.6151
R1434 B.n121 B.n120 10.6151
R1435 B.n124 B.n121 10.6151
R1436 B.n125 B.n124 10.6151
R1437 B.n128 B.n125 10.6151
R1438 B.n129 B.n128 10.6151
R1439 B.n132 B.n129 10.6151
R1440 B.n133 B.n132 10.6151
R1441 B.n136 B.n133 10.6151
R1442 B.n137 B.n136 10.6151
R1443 B.n140 B.n137 10.6151
R1444 B.n141 B.n140 10.6151
R1445 B.n144 B.n141 10.6151
R1446 B.n145 B.n144 10.6151
R1447 B.n148 B.n145 10.6151
R1448 B.n149 B.n148 10.6151
R1449 B.n152 B.n149 10.6151
R1450 B.n153 B.n152 10.6151
R1451 B.n156 B.n153 10.6151
R1452 B.n157 B.n156 10.6151
R1453 B.n160 B.n157 10.6151
R1454 B.n161 B.n160 10.6151
R1455 B.n164 B.n161 10.6151
R1456 B.n165 B.n164 10.6151
R1457 B.n168 B.n165 10.6151
R1458 B.n169 B.n168 10.6151
R1459 B.n172 B.n169 10.6151
R1460 B.n173 B.n172 10.6151
R1461 B.n176 B.n173 10.6151
R1462 B.n177 B.n176 10.6151
R1463 B.n180 B.n177 10.6151
R1464 B.n181 B.n180 10.6151
R1465 B.n184 B.n181 10.6151
R1466 B.n185 B.n184 10.6151
R1467 B.n188 B.n185 10.6151
R1468 B.n189 B.n188 10.6151
R1469 B.n192 B.n189 10.6151
R1470 B.n197 B.n194 10.6151
R1471 B.n198 B.n197 10.6151
R1472 B.n201 B.n198 10.6151
R1473 B.n202 B.n201 10.6151
R1474 B.n205 B.n202 10.6151
R1475 B.n206 B.n205 10.6151
R1476 B.n209 B.n206 10.6151
R1477 B.n210 B.n209 10.6151
R1478 B.n213 B.n210 10.6151
R1479 B.n218 B.n215 10.6151
R1480 B.n219 B.n218 10.6151
R1481 B.n222 B.n219 10.6151
R1482 B.n223 B.n222 10.6151
R1483 B.n226 B.n223 10.6151
R1484 B.n227 B.n226 10.6151
R1485 B.n230 B.n227 10.6151
R1486 B.n231 B.n230 10.6151
R1487 B.n234 B.n231 10.6151
R1488 B.n235 B.n234 10.6151
R1489 B.n238 B.n235 10.6151
R1490 B.n239 B.n238 10.6151
R1491 B.n242 B.n239 10.6151
R1492 B.n243 B.n242 10.6151
R1493 B.n246 B.n243 10.6151
R1494 B.n247 B.n246 10.6151
R1495 B.n250 B.n247 10.6151
R1496 B.n251 B.n250 10.6151
R1497 B.n254 B.n251 10.6151
R1498 B.n255 B.n254 10.6151
R1499 B.n258 B.n255 10.6151
R1500 B.n259 B.n258 10.6151
R1501 B.n262 B.n259 10.6151
R1502 B.n263 B.n262 10.6151
R1503 B.n266 B.n263 10.6151
R1504 B.n267 B.n266 10.6151
R1505 B.n270 B.n267 10.6151
R1506 B.n271 B.n270 10.6151
R1507 B.n274 B.n271 10.6151
R1508 B.n275 B.n274 10.6151
R1509 B.n278 B.n275 10.6151
R1510 B.n279 B.n278 10.6151
R1511 B.n282 B.n279 10.6151
R1512 B.n283 B.n282 10.6151
R1513 B.n286 B.n283 10.6151
R1514 B.n288 B.n286 10.6151
R1515 B.n289 B.n288 10.6151
R1516 B.n742 B.n289 10.6151
R1517 B.t5 B.n316 10.0157
R1518 B.t4 B.n29 10.0157
R1519 B.n486 B.n485 9.36635
R1520 B.n509 B.n383 9.36635
R1521 B.n193 B.n192 9.36635
R1522 B.n215 B.n214 9.36635
R1523 B.n822 B.n0 8.11757
R1524 B.n822 B.n1 8.11757
R1525 B.n332 B.t0 6.0096
R1526 B.t7 B.n777 6.0096
R1527 B.n683 B.t6 3.33889
R1528 B.n810 B.t3 3.33889
R1529 B.n487 B.n486 1.24928
R1530 B.n384 B.n383 1.24928
R1531 B.n194 B.n193 1.24928
R1532 B.n214 B.n213 1.24928
R1533 VN.n4 VN.t1 201.624
R1534 VN.n25 VN.t3 201.624
R1535 VN.n20 VN.n19 179.499
R1536 VN.n41 VN.n40 179.499
R1537 VN.n5 VN.t0 169.762
R1538 VN.n12 VN.t7 169.762
R1539 VN.n19 VN.t5 169.762
R1540 VN.n26 VN.t6 169.762
R1541 VN.n33 VN.t4 169.762
R1542 VN.n40 VN.t2 169.762
R1543 VN.n39 VN.n21 161.3
R1544 VN.n38 VN.n37 161.3
R1545 VN.n36 VN.n22 161.3
R1546 VN.n35 VN.n34 161.3
R1547 VN.n32 VN.n23 161.3
R1548 VN.n31 VN.n30 161.3
R1549 VN.n29 VN.n24 161.3
R1550 VN.n28 VN.n27 161.3
R1551 VN.n18 VN.n0 161.3
R1552 VN.n17 VN.n16 161.3
R1553 VN.n15 VN.n1 161.3
R1554 VN.n14 VN.n13 161.3
R1555 VN.n11 VN.n2 161.3
R1556 VN.n10 VN.n9 161.3
R1557 VN.n8 VN.n3 161.3
R1558 VN.n7 VN.n6 161.3
R1559 VN.n10 VN.n3 56.5617
R1560 VN.n31 VN.n24 56.5617
R1561 VN.n17 VN.n1 56.5617
R1562 VN.n38 VN.n22 56.5617
R1563 VN.n5 VN.n4 55.8951
R1564 VN.n26 VN.n25 55.8951
R1565 VN VN.n41 45.8357
R1566 VN.n6 VN.n3 24.5923
R1567 VN.n11 VN.n10 24.5923
R1568 VN.n13 VN.n1 24.5923
R1569 VN.n18 VN.n17 24.5923
R1570 VN.n27 VN.n24 24.5923
R1571 VN.n34 VN.n22 24.5923
R1572 VN.n32 VN.n31 24.5923
R1573 VN.n39 VN.n38 24.5923
R1574 VN.n28 VN.n25 18.12
R1575 VN.n7 VN.n4 18.12
R1576 VN.n13 VN.n12 14.2638
R1577 VN.n34 VN.n33 14.2638
R1578 VN.n6 VN.n5 10.3291
R1579 VN.n12 VN.n11 10.3291
R1580 VN.n27 VN.n26 10.3291
R1581 VN.n33 VN.n32 10.3291
R1582 VN.n19 VN.n18 6.39438
R1583 VN.n40 VN.n39 6.39438
R1584 VN.n41 VN.n21 0.189894
R1585 VN.n37 VN.n21 0.189894
R1586 VN.n37 VN.n36 0.189894
R1587 VN.n36 VN.n35 0.189894
R1588 VN.n35 VN.n23 0.189894
R1589 VN.n30 VN.n23 0.189894
R1590 VN.n30 VN.n29 0.189894
R1591 VN.n29 VN.n28 0.189894
R1592 VN.n8 VN.n7 0.189894
R1593 VN.n9 VN.n8 0.189894
R1594 VN.n9 VN.n2 0.189894
R1595 VN.n14 VN.n2 0.189894
R1596 VN.n15 VN.n14 0.189894
R1597 VN.n16 VN.n15 0.189894
R1598 VN.n16 VN.n0 0.189894
R1599 VN.n20 VN.n0 0.189894
R1600 VN VN.n20 0.0516364
R1601 VDD2.n2 VDD2.n1 66.0842
R1602 VDD2.n2 VDD2.n0 66.0842
R1603 VDD2 VDD2.n5 66.0814
R1604 VDD2.n4 VDD2.n3 65.3122
R1605 VDD2.n4 VDD2.n2 40.8187
R1606 VDD2.n5 VDD2.t1 1.76836
R1607 VDD2.n5 VDD2.t4 1.76836
R1608 VDD2.n3 VDD2.t5 1.76836
R1609 VDD2.n3 VDD2.t3 1.76836
R1610 VDD2.n1 VDD2.t0 1.76836
R1611 VDD2.n1 VDD2.t2 1.76836
R1612 VDD2.n0 VDD2.t6 1.76836
R1613 VDD2.n0 VDD2.t7 1.76836
R1614 VDD2 VDD2.n4 0.886276
C0 VDD2 VP 0.4126f
C1 VDD1 VP 7.472681f
C2 VTAIL VN 7.31433f
C3 VTAIL VDD2 8.05912f
C4 VDD1 VTAIL 8.01148f
C5 VTAIL VP 7.32844f
C6 VDD2 VN 7.21127f
C7 VDD1 VN 0.150306f
C8 VN VP 6.27554f
C9 VDD1 VDD2 1.2552f
C10 VDD2 B 4.315382f
C11 VDD1 B 4.643737f
C12 VTAIL B 9.256275f
C13 VN B 11.621039f
C14 VP B 10.057056f
C15 VDD2.t6 B 0.220445f
C16 VDD2.t7 B 0.220445f
C17 VDD2.n0 B 1.96337f
C18 VDD2.t0 B 0.220445f
C19 VDD2.t2 B 0.220445f
C20 VDD2.n1 B 1.96337f
C21 VDD2.n2 B 2.62718f
C22 VDD2.t5 B 0.220445f
C23 VDD2.t3 B 0.220445f
C24 VDD2.n3 B 1.95861f
C25 VDD2.n4 B 2.52551f
C26 VDD2.t1 B 0.220445f
C27 VDD2.t4 B 0.220445f
C28 VDD2.n5 B 1.96334f
C29 VN.n0 B 0.030031f
C30 VN.t5 B 1.45412f
C31 VN.n1 B 0.037007f
C32 VN.n2 B 0.030031f
C33 VN.t7 B 1.45412f
C34 VN.n3 B 0.043654f
C35 VN.t1 B 1.55646f
C36 VN.n4 B 0.599792f
C37 VN.t0 B 1.45412f
C38 VN.n5 B 0.5829f
C39 VN.n6 B 0.039744f
C40 VN.n7 B 0.190353f
C41 VN.n8 B 0.030031f
C42 VN.n9 B 0.030031f
C43 VN.n10 B 0.043654f
C44 VN.n11 B 0.039744f
C45 VN.n12 B 0.527067f
C46 VN.n13 B 0.044142f
C47 VN.n14 B 0.030031f
C48 VN.n15 B 0.030031f
C49 VN.n16 B 0.030031f
C50 VN.n17 B 0.050301f
C51 VN.n18 B 0.035345f
C52 VN.n19 B 0.58798f
C53 VN.n20 B 0.030145f
C54 VN.n21 B 0.030031f
C55 VN.t2 B 1.45412f
C56 VN.n22 B 0.037007f
C57 VN.n23 B 0.030031f
C58 VN.t4 B 1.45412f
C59 VN.n24 B 0.043654f
C60 VN.t3 B 1.55646f
C61 VN.n25 B 0.599792f
C62 VN.t6 B 1.45412f
C63 VN.n26 B 0.5829f
C64 VN.n27 B 0.039744f
C65 VN.n28 B 0.190353f
C66 VN.n29 B 0.030031f
C67 VN.n30 B 0.030031f
C68 VN.n31 B 0.043654f
C69 VN.n32 B 0.039744f
C70 VN.n33 B 0.527067f
C71 VN.n34 B 0.044142f
C72 VN.n35 B 0.030031f
C73 VN.n36 B 0.030031f
C74 VN.n37 B 0.030031f
C75 VN.n38 B 0.050301f
C76 VN.n39 B 0.035345f
C77 VN.n40 B 0.58798f
C78 VN.n41 B 1.4359f
C79 VDD1.t1 B 0.221991f
C80 VDD1.t2 B 0.221991f
C81 VDD1.n0 B 1.97796f
C82 VDD1.t6 B 0.221991f
C83 VDD1.t5 B 0.221991f
C84 VDD1.n1 B 1.97715f
C85 VDD1.t0 B 0.221991f
C86 VDD1.t7 B 0.221991f
C87 VDD1.n2 B 1.97715f
C88 VDD1.n3 B 2.69851f
C89 VDD1.t3 B 0.221991f
C90 VDD1.t4 B 0.221991f
C91 VDD1.n4 B 1.97235f
C92 VDD1.n5 B 2.57357f
C93 VTAIL.t1 B 0.171947f
C94 VTAIL.t4 B 0.171947f
C95 VTAIL.n0 B 1.47486f
C96 VTAIL.n1 B 0.291531f
C97 VTAIL.t3 B 1.88165f
C98 VTAIL.n2 B 0.379454f
C99 VTAIL.t10 B 1.88165f
C100 VTAIL.n3 B 0.379454f
C101 VTAIL.t13 B 0.171947f
C102 VTAIL.t7 B 0.171947f
C103 VTAIL.n4 B 1.47486f
C104 VTAIL.n5 B 0.391504f
C105 VTAIL.t14 B 1.88165f
C106 VTAIL.n6 B 1.32198f
C107 VTAIL.t0 B 1.88166f
C108 VTAIL.n7 B 1.32197f
C109 VTAIL.t5 B 0.171947f
C110 VTAIL.t2 B 0.171947f
C111 VTAIL.n8 B 1.47486f
C112 VTAIL.n9 B 0.391499f
C113 VTAIL.t6 B 1.88166f
C114 VTAIL.n10 B 0.379442f
C115 VTAIL.t8 B 1.88166f
C116 VTAIL.n11 B 0.379442f
C117 VTAIL.t9 B 0.171947f
C118 VTAIL.t11 B 0.171947f
C119 VTAIL.n12 B 1.47486f
C120 VTAIL.n13 B 0.391499f
C121 VTAIL.t12 B 1.88165f
C122 VTAIL.n14 B 1.32198f
C123 VTAIL.t15 B 1.88165f
C124 VTAIL.n15 B 1.31834f
C125 VP.n0 B 0.030526f
C126 VP.t0 B 1.47809f
C127 VP.n1 B 0.037618f
C128 VP.n2 B 0.030526f
C129 VP.t7 B 1.47809f
C130 VP.n3 B 0.044374f
C131 VP.n4 B 0.030526f
C132 VP.t2 B 1.47809f
C133 VP.n5 B 0.051131f
C134 VP.n6 B 0.030526f
C135 VP.t3 B 1.47809f
C136 VP.n7 B 0.037618f
C137 VP.n8 B 0.030526f
C138 VP.t4 B 1.47809f
C139 VP.n9 B 0.044374f
C140 VP.t6 B 1.58211f
C141 VP.n10 B 0.60968f
C142 VP.t5 B 1.47809f
C143 VP.n11 B 0.592509f
C144 VP.n12 B 0.040399f
C145 VP.n13 B 0.193491f
C146 VP.n14 B 0.030526f
C147 VP.n15 B 0.030526f
C148 VP.n16 B 0.044374f
C149 VP.n17 B 0.040399f
C150 VP.n18 B 0.535756f
C151 VP.n19 B 0.04487f
C152 VP.n20 B 0.030526f
C153 VP.n21 B 0.030526f
C154 VP.n22 B 0.030526f
C155 VP.n23 B 0.051131f
C156 VP.n24 B 0.035928f
C157 VP.n25 B 0.597674f
C158 VP.n26 B 1.43962f
C159 VP.n27 B 1.46383f
C160 VP.t1 B 1.47809f
C161 VP.n28 B 0.597674f
C162 VP.n29 B 0.035928f
C163 VP.n30 B 0.030526f
C164 VP.n31 B 0.030526f
C165 VP.n32 B 0.030526f
C166 VP.n33 B 0.037618f
C167 VP.n34 B 0.04487f
C168 VP.n35 B 0.535756f
C169 VP.n36 B 0.040399f
C170 VP.n37 B 0.030526f
C171 VP.n38 B 0.030526f
C172 VP.n39 B 0.030526f
C173 VP.n40 B 0.044374f
C174 VP.n41 B 0.040399f
C175 VP.n42 B 0.535756f
C176 VP.n43 B 0.04487f
C177 VP.n44 B 0.030526f
C178 VP.n45 B 0.030526f
C179 VP.n46 B 0.030526f
C180 VP.n47 B 0.051131f
C181 VP.n48 B 0.035928f
C182 VP.n49 B 0.597674f
C183 VP.n50 B 0.030642f
.ends

