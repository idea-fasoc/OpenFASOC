* NGSPICE file created from diff_pair_sample_0492.ext - technology: sky130A

.subckt diff_pair_sample_0492 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n3242_n1470# sky130_fd_pr__pfet_01v8 ad=0.9789 pd=5.8 as=0 ps=0 w=2.51 l=2.51
X1 VTAIL.t11 VN.t0 VDD2.t1 w_n3242_n1470# sky130_fd_pr__pfet_01v8 ad=0.41415 pd=2.84 as=0.41415 ps=2.84 w=2.51 l=2.51
X2 VTAIL.t5 VP.t0 VDD1.t5 w_n3242_n1470# sky130_fd_pr__pfet_01v8 ad=0.41415 pd=2.84 as=0.41415 ps=2.84 w=2.51 l=2.51
X3 VDD1.t4 VP.t1 VTAIL.t4 w_n3242_n1470# sky130_fd_pr__pfet_01v8 ad=0.41415 pd=2.84 as=0.9789 ps=5.8 w=2.51 l=2.51
X4 VDD1.t3 VP.t2 VTAIL.t0 w_n3242_n1470# sky130_fd_pr__pfet_01v8 ad=0.41415 pd=2.84 as=0.9789 ps=5.8 w=2.51 l=2.51
X5 VDD1.t2 VP.t3 VTAIL.t1 w_n3242_n1470# sky130_fd_pr__pfet_01v8 ad=0.9789 pd=5.8 as=0.41415 ps=2.84 w=2.51 l=2.51
X6 B.t8 B.t6 B.t7 w_n3242_n1470# sky130_fd_pr__pfet_01v8 ad=0.9789 pd=5.8 as=0 ps=0 w=2.51 l=2.51
X7 VDD2.t0 VN.t1 VTAIL.t10 w_n3242_n1470# sky130_fd_pr__pfet_01v8 ad=0.41415 pd=2.84 as=0.9789 ps=5.8 w=2.51 l=2.51
X8 B.t5 B.t3 B.t4 w_n3242_n1470# sky130_fd_pr__pfet_01v8 ad=0.9789 pd=5.8 as=0 ps=0 w=2.51 l=2.51
X9 VDD2.t2 VN.t2 VTAIL.t9 w_n3242_n1470# sky130_fd_pr__pfet_01v8 ad=0.41415 pd=2.84 as=0.9789 ps=5.8 w=2.51 l=2.51
X10 VDD2.t5 VN.t3 VTAIL.t8 w_n3242_n1470# sky130_fd_pr__pfet_01v8 ad=0.9789 pd=5.8 as=0.41415 ps=2.84 w=2.51 l=2.51
X11 VTAIL.t7 VN.t4 VDD2.t4 w_n3242_n1470# sky130_fd_pr__pfet_01v8 ad=0.41415 pd=2.84 as=0.41415 ps=2.84 w=2.51 l=2.51
X12 VDD2.t3 VN.t5 VTAIL.t6 w_n3242_n1470# sky130_fd_pr__pfet_01v8 ad=0.9789 pd=5.8 as=0.41415 ps=2.84 w=2.51 l=2.51
X13 B.t2 B.t0 B.t1 w_n3242_n1470# sky130_fd_pr__pfet_01v8 ad=0.9789 pd=5.8 as=0 ps=0 w=2.51 l=2.51
X14 VTAIL.t2 VP.t4 VDD1.t1 w_n3242_n1470# sky130_fd_pr__pfet_01v8 ad=0.41415 pd=2.84 as=0.41415 ps=2.84 w=2.51 l=2.51
X15 VDD1.t0 VP.t5 VTAIL.t3 w_n3242_n1470# sky130_fd_pr__pfet_01v8 ad=0.9789 pd=5.8 as=0.41415 ps=2.84 w=2.51 l=2.51
R0 B.n247 B.n246 585
R1 B.n245 B.n88 585
R2 B.n244 B.n243 585
R3 B.n242 B.n89 585
R4 B.n241 B.n240 585
R5 B.n239 B.n90 585
R6 B.n238 B.n237 585
R7 B.n236 B.n91 585
R8 B.n235 B.n234 585
R9 B.n233 B.n92 585
R10 B.n232 B.n231 585
R11 B.n230 B.n93 585
R12 B.n229 B.n228 585
R13 B.n227 B.n94 585
R14 B.n226 B.n225 585
R15 B.n221 B.n95 585
R16 B.n220 B.n219 585
R17 B.n218 B.n96 585
R18 B.n217 B.n216 585
R19 B.n215 B.n97 585
R20 B.n214 B.n213 585
R21 B.n212 B.n98 585
R22 B.n211 B.n210 585
R23 B.n208 B.n99 585
R24 B.n207 B.n206 585
R25 B.n205 B.n102 585
R26 B.n204 B.n203 585
R27 B.n202 B.n103 585
R28 B.n201 B.n200 585
R29 B.n199 B.n104 585
R30 B.n198 B.n197 585
R31 B.n196 B.n105 585
R32 B.n195 B.n194 585
R33 B.n193 B.n106 585
R34 B.n192 B.n191 585
R35 B.n190 B.n107 585
R36 B.n189 B.n188 585
R37 B.n248 B.n87 585
R38 B.n250 B.n249 585
R39 B.n251 B.n86 585
R40 B.n253 B.n252 585
R41 B.n254 B.n85 585
R42 B.n256 B.n255 585
R43 B.n257 B.n84 585
R44 B.n259 B.n258 585
R45 B.n260 B.n83 585
R46 B.n262 B.n261 585
R47 B.n263 B.n82 585
R48 B.n265 B.n264 585
R49 B.n266 B.n81 585
R50 B.n268 B.n267 585
R51 B.n269 B.n80 585
R52 B.n271 B.n270 585
R53 B.n272 B.n79 585
R54 B.n274 B.n273 585
R55 B.n275 B.n78 585
R56 B.n277 B.n276 585
R57 B.n278 B.n77 585
R58 B.n280 B.n279 585
R59 B.n281 B.n76 585
R60 B.n283 B.n282 585
R61 B.n284 B.n75 585
R62 B.n286 B.n285 585
R63 B.n287 B.n74 585
R64 B.n289 B.n288 585
R65 B.n290 B.n73 585
R66 B.n292 B.n291 585
R67 B.n293 B.n72 585
R68 B.n295 B.n294 585
R69 B.n296 B.n71 585
R70 B.n298 B.n297 585
R71 B.n299 B.n70 585
R72 B.n301 B.n300 585
R73 B.n302 B.n69 585
R74 B.n304 B.n303 585
R75 B.n305 B.n68 585
R76 B.n307 B.n306 585
R77 B.n308 B.n67 585
R78 B.n310 B.n309 585
R79 B.n311 B.n66 585
R80 B.n313 B.n312 585
R81 B.n314 B.n65 585
R82 B.n316 B.n315 585
R83 B.n317 B.n64 585
R84 B.n319 B.n318 585
R85 B.n320 B.n63 585
R86 B.n322 B.n321 585
R87 B.n323 B.n62 585
R88 B.n325 B.n324 585
R89 B.n326 B.n61 585
R90 B.n328 B.n327 585
R91 B.n329 B.n60 585
R92 B.n331 B.n330 585
R93 B.n332 B.n59 585
R94 B.n334 B.n333 585
R95 B.n335 B.n58 585
R96 B.n337 B.n336 585
R97 B.n338 B.n57 585
R98 B.n340 B.n339 585
R99 B.n341 B.n56 585
R100 B.n343 B.n342 585
R101 B.n344 B.n55 585
R102 B.n346 B.n345 585
R103 B.n347 B.n54 585
R104 B.n349 B.n348 585
R105 B.n350 B.n53 585
R106 B.n352 B.n351 585
R107 B.n353 B.n52 585
R108 B.n355 B.n354 585
R109 B.n356 B.n51 585
R110 B.n358 B.n357 585
R111 B.n359 B.n50 585
R112 B.n361 B.n360 585
R113 B.n362 B.n49 585
R114 B.n364 B.n363 585
R115 B.n365 B.n48 585
R116 B.n367 B.n366 585
R117 B.n368 B.n47 585
R118 B.n370 B.n369 585
R119 B.n371 B.n46 585
R120 B.n373 B.n372 585
R121 B.n430 B.n429 585
R122 B.n428 B.n23 585
R123 B.n427 B.n426 585
R124 B.n425 B.n24 585
R125 B.n424 B.n423 585
R126 B.n422 B.n25 585
R127 B.n421 B.n420 585
R128 B.n419 B.n26 585
R129 B.n418 B.n417 585
R130 B.n416 B.n27 585
R131 B.n415 B.n414 585
R132 B.n413 B.n28 585
R133 B.n412 B.n411 585
R134 B.n410 B.n29 585
R135 B.n408 B.n407 585
R136 B.n406 B.n32 585
R137 B.n405 B.n404 585
R138 B.n403 B.n33 585
R139 B.n402 B.n401 585
R140 B.n400 B.n34 585
R141 B.n399 B.n398 585
R142 B.n397 B.n35 585
R143 B.n396 B.n395 585
R144 B.n394 B.n393 585
R145 B.n392 B.n39 585
R146 B.n391 B.n390 585
R147 B.n389 B.n40 585
R148 B.n388 B.n387 585
R149 B.n386 B.n41 585
R150 B.n385 B.n384 585
R151 B.n383 B.n42 585
R152 B.n382 B.n381 585
R153 B.n380 B.n43 585
R154 B.n379 B.n378 585
R155 B.n377 B.n44 585
R156 B.n376 B.n375 585
R157 B.n374 B.n45 585
R158 B.n431 B.n22 585
R159 B.n433 B.n432 585
R160 B.n434 B.n21 585
R161 B.n436 B.n435 585
R162 B.n437 B.n20 585
R163 B.n439 B.n438 585
R164 B.n440 B.n19 585
R165 B.n442 B.n441 585
R166 B.n443 B.n18 585
R167 B.n445 B.n444 585
R168 B.n446 B.n17 585
R169 B.n448 B.n447 585
R170 B.n449 B.n16 585
R171 B.n451 B.n450 585
R172 B.n452 B.n15 585
R173 B.n454 B.n453 585
R174 B.n455 B.n14 585
R175 B.n457 B.n456 585
R176 B.n458 B.n13 585
R177 B.n460 B.n459 585
R178 B.n461 B.n12 585
R179 B.n463 B.n462 585
R180 B.n464 B.n11 585
R181 B.n466 B.n465 585
R182 B.n467 B.n10 585
R183 B.n469 B.n468 585
R184 B.n470 B.n9 585
R185 B.n472 B.n471 585
R186 B.n473 B.n8 585
R187 B.n475 B.n474 585
R188 B.n476 B.n7 585
R189 B.n478 B.n477 585
R190 B.n479 B.n6 585
R191 B.n481 B.n480 585
R192 B.n482 B.n5 585
R193 B.n484 B.n483 585
R194 B.n485 B.n4 585
R195 B.n487 B.n486 585
R196 B.n488 B.n3 585
R197 B.n490 B.n489 585
R198 B.n491 B.n0 585
R199 B.n2 B.n1 585
R200 B.n129 B.n128 585
R201 B.n130 B.n127 585
R202 B.n132 B.n131 585
R203 B.n133 B.n126 585
R204 B.n135 B.n134 585
R205 B.n136 B.n125 585
R206 B.n138 B.n137 585
R207 B.n139 B.n124 585
R208 B.n141 B.n140 585
R209 B.n142 B.n123 585
R210 B.n144 B.n143 585
R211 B.n145 B.n122 585
R212 B.n147 B.n146 585
R213 B.n148 B.n121 585
R214 B.n150 B.n149 585
R215 B.n151 B.n120 585
R216 B.n153 B.n152 585
R217 B.n154 B.n119 585
R218 B.n156 B.n155 585
R219 B.n157 B.n118 585
R220 B.n159 B.n158 585
R221 B.n160 B.n117 585
R222 B.n162 B.n161 585
R223 B.n163 B.n116 585
R224 B.n165 B.n164 585
R225 B.n166 B.n115 585
R226 B.n168 B.n167 585
R227 B.n169 B.n114 585
R228 B.n171 B.n170 585
R229 B.n172 B.n113 585
R230 B.n174 B.n173 585
R231 B.n175 B.n112 585
R232 B.n177 B.n176 585
R233 B.n178 B.n111 585
R234 B.n180 B.n179 585
R235 B.n181 B.n110 585
R236 B.n183 B.n182 585
R237 B.n184 B.n109 585
R238 B.n186 B.n185 585
R239 B.n187 B.n108 585
R240 B.n188 B.n187 502.111
R241 B.n246 B.n87 502.111
R242 B.n372 B.n45 502.111
R243 B.n431 B.n430 502.111
R244 B.n222 B.t7 279.524
R245 B.n36 B.t2 279.524
R246 B.n100 B.t10 279.524
R247 B.n30 B.t5 279.524
R248 B.n493 B.n492 256.663
R249 B.n492 B.n491 235.042
R250 B.n492 B.n2 235.042
R251 B.n100 B.t9 232.007
R252 B.n222 B.t6 232.007
R253 B.n36 B.t0 232.007
R254 B.n30 B.t3 232.007
R255 B.n223 B.t8 224.446
R256 B.n37 B.t1 224.446
R257 B.n101 B.t11 224.446
R258 B.n31 B.t4 224.446
R259 B.n188 B.n107 163.367
R260 B.n192 B.n107 163.367
R261 B.n193 B.n192 163.367
R262 B.n194 B.n193 163.367
R263 B.n194 B.n105 163.367
R264 B.n198 B.n105 163.367
R265 B.n199 B.n198 163.367
R266 B.n200 B.n199 163.367
R267 B.n200 B.n103 163.367
R268 B.n204 B.n103 163.367
R269 B.n205 B.n204 163.367
R270 B.n206 B.n205 163.367
R271 B.n206 B.n99 163.367
R272 B.n211 B.n99 163.367
R273 B.n212 B.n211 163.367
R274 B.n213 B.n212 163.367
R275 B.n213 B.n97 163.367
R276 B.n217 B.n97 163.367
R277 B.n218 B.n217 163.367
R278 B.n219 B.n218 163.367
R279 B.n219 B.n95 163.367
R280 B.n226 B.n95 163.367
R281 B.n227 B.n226 163.367
R282 B.n228 B.n227 163.367
R283 B.n228 B.n93 163.367
R284 B.n232 B.n93 163.367
R285 B.n233 B.n232 163.367
R286 B.n234 B.n233 163.367
R287 B.n234 B.n91 163.367
R288 B.n238 B.n91 163.367
R289 B.n239 B.n238 163.367
R290 B.n240 B.n239 163.367
R291 B.n240 B.n89 163.367
R292 B.n244 B.n89 163.367
R293 B.n245 B.n244 163.367
R294 B.n246 B.n245 163.367
R295 B.n372 B.n371 163.367
R296 B.n371 B.n370 163.367
R297 B.n370 B.n47 163.367
R298 B.n366 B.n47 163.367
R299 B.n366 B.n365 163.367
R300 B.n365 B.n364 163.367
R301 B.n364 B.n49 163.367
R302 B.n360 B.n49 163.367
R303 B.n360 B.n359 163.367
R304 B.n359 B.n358 163.367
R305 B.n358 B.n51 163.367
R306 B.n354 B.n51 163.367
R307 B.n354 B.n353 163.367
R308 B.n353 B.n352 163.367
R309 B.n352 B.n53 163.367
R310 B.n348 B.n53 163.367
R311 B.n348 B.n347 163.367
R312 B.n347 B.n346 163.367
R313 B.n346 B.n55 163.367
R314 B.n342 B.n55 163.367
R315 B.n342 B.n341 163.367
R316 B.n341 B.n340 163.367
R317 B.n340 B.n57 163.367
R318 B.n336 B.n57 163.367
R319 B.n336 B.n335 163.367
R320 B.n335 B.n334 163.367
R321 B.n334 B.n59 163.367
R322 B.n330 B.n59 163.367
R323 B.n330 B.n329 163.367
R324 B.n329 B.n328 163.367
R325 B.n328 B.n61 163.367
R326 B.n324 B.n61 163.367
R327 B.n324 B.n323 163.367
R328 B.n323 B.n322 163.367
R329 B.n322 B.n63 163.367
R330 B.n318 B.n63 163.367
R331 B.n318 B.n317 163.367
R332 B.n317 B.n316 163.367
R333 B.n316 B.n65 163.367
R334 B.n312 B.n65 163.367
R335 B.n312 B.n311 163.367
R336 B.n311 B.n310 163.367
R337 B.n310 B.n67 163.367
R338 B.n306 B.n67 163.367
R339 B.n306 B.n305 163.367
R340 B.n305 B.n304 163.367
R341 B.n304 B.n69 163.367
R342 B.n300 B.n69 163.367
R343 B.n300 B.n299 163.367
R344 B.n299 B.n298 163.367
R345 B.n298 B.n71 163.367
R346 B.n294 B.n71 163.367
R347 B.n294 B.n293 163.367
R348 B.n293 B.n292 163.367
R349 B.n292 B.n73 163.367
R350 B.n288 B.n73 163.367
R351 B.n288 B.n287 163.367
R352 B.n287 B.n286 163.367
R353 B.n286 B.n75 163.367
R354 B.n282 B.n75 163.367
R355 B.n282 B.n281 163.367
R356 B.n281 B.n280 163.367
R357 B.n280 B.n77 163.367
R358 B.n276 B.n77 163.367
R359 B.n276 B.n275 163.367
R360 B.n275 B.n274 163.367
R361 B.n274 B.n79 163.367
R362 B.n270 B.n79 163.367
R363 B.n270 B.n269 163.367
R364 B.n269 B.n268 163.367
R365 B.n268 B.n81 163.367
R366 B.n264 B.n81 163.367
R367 B.n264 B.n263 163.367
R368 B.n263 B.n262 163.367
R369 B.n262 B.n83 163.367
R370 B.n258 B.n83 163.367
R371 B.n258 B.n257 163.367
R372 B.n257 B.n256 163.367
R373 B.n256 B.n85 163.367
R374 B.n252 B.n85 163.367
R375 B.n252 B.n251 163.367
R376 B.n251 B.n250 163.367
R377 B.n250 B.n87 163.367
R378 B.n430 B.n23 163.367
R379 B.n426 B.n23 163.367
R380 B.n426 B.n425 163.367
R381 B.n425 B.n424 163.367
R382 B.n424 B.n25 163.367
R383 B.n420 B.n25 163.367
R384 B.n420 B.n419 163.367
R385 B.n419 B.n418 163.367
R386 B.n418 B.n27 163.367
R387 B.n414 B.n27 163.367
R388 B.n414 B.n413 163.367
R389 B.n413 B.n412 163.367
R390 B.n412 B.n29 163.367
R391 B.n407 B.n29 163.367
R392 B.n407 B.n406 163.367
R393 B.n406 B.n405 163.367
R394 B.n405 B.n33 163.367
R395 B.n401 B.n33 163.367
R396 B.n401 B.n400 163.367
R397 B.n400 B.n399 163.367
R398 B.n399 B.n35 163.367
R399 B.n395 B.n35 163.367
R400 B.n395 B.n394 163.367
R401 B.n394 B.n39 163.367
R402 B.n390 B.n39 163.367
R403 B.n390 B.n389 163.367
R404 B.n389 B.n388 163.367
R405 B.n388 B.n41 163.367
R406 B.n384 B.n41 163.367
R407 B.n384 B.n383 163.367
R408 B.n383 B.n382 163.367
R409 B.n382 B.n43 163.367
R410 B.n378 B.n43 163.367
R411 B.n378 B.n377 163.367
R412 B.n377 B.n376 163.367
R413 B.n376 B.n45 163.367
R414 B.n432 B.n431 163.367
R415 B.n432 B.n21 163.367
R416 B.n436 B.n21 163.367
R417 B.n437 B.n436 163.367
R418 B.n438 B.n437 163.367
R419 B.n438 B.n19 163.367
R420 B.n442 B.n19 163.367
R421 B.n443 B.n442 163.367
R422 B.n444 B.n443 163.367
R423 B.n444 B.n17 163.367
R424 B.n448 B.n17 163.367
R425 B.n449 B.n448 163.367
R426 B.n450 B.n449 163.367
R427 B.n450 B.n15 163.367
R428 B.n454 B.n15 163.367
R429 B.n455 B.n454 163.367
R430 B.n456 B.n455 163.367
R431 B.n456 B.n13 163.367
R432 B.n460 B.n13 163.367
R433 B.n461 B.n460 163.367
R434 B.n462 B.n461 163.367
R435 B.n462 B.n11 163.367
R436 B.n466 B.n11 163.367
R437 B.n467 B.n466 163.367
R438 B.n468 B.n467 163.367
R439 B.n468 B.n9 163.367
R440 B.n472 B.n9 163.367
R441 B.n473 B.n472 163.367
R442 B.n474 B.n473 163.367
R443 B.n474 B.n7 163.367
R444 B.n478 B.n7 163.367
R445 B.n479 B.n478 163.367
R446 B.n480 B.n479 163.367
R447 B.n480 B.n5 163.367
R448 B.n484 B.n5 163.367
R449 B.n485 B.n484 163.367
R450 B.n486 B.n485 163.367
R451 B.n486 B.n3 163.367
R452 B.n490 B.n3 163.367
R453 B.n491 B.n490 163.367
R454 B.n128 B.n2 163.367
R455 B.n128 B.n127 163.367
R456 B.n132 B.n127 163.367
R457 B.n133 B.n132 163.367
R458 B.n134 B.n133 163.367
R459 B.n134 B.n125 163.367
R460 B.n138 B.n125 163.367
R461 B.n139 B.n138 163.367
R462 B.n140 B.n139 163.367
R463 B.n140 B.n123 163.367
R464 B.n144 B.n123 163.367
R465 B.n145 B.n144 163.367
R466 B.n146 B.n145 163.367
R467 B.n146 B.n121 163.367
R468 B.n150 B.n121 163.367
R469 B.n151 B.n150 163.367
R470 B.n152 B.n151 163.367
R471 B.n152 B.n119 163.367
R472 B.n156 B.n119 163.367
R473 B.n157 B.n156 163.367
R474 B.n158 B.n157 163.367
R475 B.n158 B.n117 163.367
R476 B.n162 B.n117 163.367
R477 B.n163 B.n162 163.367
R478 B.n164 B.n163 163.367
R479 B.n164 B.n115 163.367
R480 B.n168 B.n115 163.367
R481 B.n169 B.n168 163.367
R482 B.n170 B.n169 163.367
R483 B.n170 B.n113 163.367
R484 B.n174 B.n113 163.367
R485 B.n175 B.n174 163.367
R486 B.n176 B.n175 163.367
R487 B.n176 B.n111 163.367
R488 B.n180 B.n111 163.367
R489 B.n181 B.n180 163.367
R490 B.n182 B.n181 163.367
R491 B.n182 B.n109 163.367
R492 B.n186 B.n109 163.367
R493 B.n187 B.n186 163.367
R494 B.n209 B.n101 59.5399
R495 B.n224 B.n223 59.5399
R496 B.n38 B.n37 59.5399
R497 B.n409 B.n31 59.5399
R498 B.n101 B.n100 55.0793
R499 B.n223 B.n222 55.0793
R500 B.n37 B.n36 55.0793
R501 B.n31 B.n30 55.0793
R502 B.n429 B.n22 32.6249
R503 B.n374 B.n373 32.6249
R504 B.n248 B.n247 32.6249
R505 B.n189 B.n108 32.6249
R506 B B.n493 18.0485
R507 B.n433 B.n22 10.6151
R508 B.n434 B.n433 10.6151
R509 B.n435 B.n434 10.6151
R510 B.n435 B.n20 10.6151
R511 B.n439 B.n20 10.6151
R512 B.n440 B.n439 10.6151
R513 B.n441 B.n440 10.6151
R514 B.n441 B.n18 10.6151
R515 B.n445 B.n18 10.6151
R516 B.n446 B.n445 10.6151
R517 B.n447 B.n446 10.6151
R518 B.n447 B.n16 10.6151
R519 B.n451 B.n16 10.6151
R520 B.n452 B.n451 10.6151
R521 B.n453 B.n452 10.6151
R522 B.n453 B.n14 10.6151
R523 B.n457 B.n14 10.6151
R524 B.n458 B.n457 10.6151
R525 B.n459 B.n458 10.6151
R526 B.n459 B.n12 10.6151
R527 B.n463 B.n12 10.6151
R528 B.n464 B.n463 10.6151
R529 B.n465 B.n464 10.6151
R530 B.n465 B.n10 10.6151
R531 B.n469 B.n10 10.6151
R532 B.n470 B.n469 10.6151
R533 B.n471 B.n470 10.6151
R534 B.n471 B.n8 10.6151
R535 B.n475 B.n8 10.6151
R536 B.n476 B.n475 10.6151
R537 B.n477 B.n476 10.6151
R538 B.n477 B.n6 10.6151
R539 B.n481 B.n6 10.6151
R540 B.n482 B.n481 10.6151
R541 B.n483 B.n482 10.6151
R542 B.n483 B.n4 10.6151
R543 B.n487 B.n4 10.6151
R544 B.n488 B.n487 10.6151
R545 B.n489 B.n488 10.6151
R546 B.n489 B.n0 10.6151
R547 B.n429 B.n428 10.6151
R548 B.n428 B.n427 10.6151
R549 B.n427 B.n24 10.6151
R550 B.n423 B.n24 10.6151
R551 B.n423 B.n422 10.6151
R552 B.n422 B.n421 10.6151
R553 B.n421 B.n26 10.6151
R554 B.n417 B.n26 10.6151
R555 B.n417 B.n416 10.6151
R556 B.n416 B.n415 10.6151
R557 B.n415 B.n28 10.6151
R558 B.n411 B.n28 10.6151
R559 B.n411 B.n410 10.6151
R560 B.n408 B.n32 10.6151
R561 B.n404 B.n32 10.6151
R562 B.n404 B.n403 10.6151
R563 B.n403 B.n402 10.6151
R564 B.n402 B.n34 10.6151
R565 B.n398 B.n34 10.6151
R566 B.n398 B.n397 10.6151
R567 B.n397 B.n396 10.6151
R568 B.n393 B.n392 10.6151
R569 B.n392 B.n391 10.6151
R570 B.n391 B.n40 10.6151
R571 B.n387 B.n40 10.6151
R572 B.n387 B.n386 10.6151
R573 B.n386 B.n385 10.6151
R574 B.n385 B.n42 10.6151
R575 B.n381 B.n42 10.6151
R576 B.n381 B.n380 10.6151
R577 B.n380 B.n379 10.6151
R578 B.n379 B.n44 10.6151
R579 B.n375 B.n44 10.6151
R580 B.n375 B.n374 10.6151
R581 B.n373 B.n46 10.6151
R582 B.n369 B.n46 10.6151
R583 B.n369 B.n368 10.6151
R584 B.n368 B.n367 10.6151
R585 B.n367 B.n48 10.6151
R586 B.n363 B.n48 10.6151
R587 B.n363 B.n362 10.6151
R588 B.n362 B.n361 10.6151
R589 B.n361 B.n50 10.6151
R590 B.n357 B.n50 10.6151
R591 B.n357 B.n356 10.6151
R592 B.n356 B.n355 10.6151
R593 B.n355 B.n52 10.6151
R594 B.n351 B.n52 10.6151
R595 B.n351 B.n350 10.6151
R596 B.n350 B.n349 10.6151
R597 B.n349 B.n54 10.6151
R598 B.n345 B.n54 10.6151
R599 B.n345 B.n344 10.6151
R600 B.n344 B.n343 10.6151
R601 B.n343 B.n56 10.6151
R602 B.n339 B.n56 10.6151
R603 B.n339 B.n338 10.6151
R604 B.n338 B.n337 10.6151
R605 B.n337 B.n58 10.6151
R606 B.n333 B.n58 10.6151
R607 B.n333 B.n332 10.6151
R608 B.n332 B.n331 10.6151
R609 B.n331 B.n60 10.6151
R610 B.n327 B.n60 10.6151
R611 B.n327 B.n326 10.6151
R612 B.n326 B.n325 10.6151
R613 B.n325 B.n62 10.6151
R614 B.n321 B.n62 10.6151
R615 B.n321 B.n320 10.6151
R616 B.n320 B.n319 10.6151
R617 B.n319 B.n64 10.6151
R618 B.n315 B.n64 10.6151
R619 B.n315 B.n314 10.6151
R620 B.n314 B.n313 10.6151
R621 B.n313 B.n66 10.6151
R622 B.n309 B.n66 10.6151
R623 B.n309 B.n308 10.6151
R624 B.n308 B.n307 10.6151
R625 B.n307 B.n68 10.6151
R626 B.n303 B.n68 10.6151
R627 B.n303 B.n302 10.6151
R628 B.n302 B.n301 10.6151
R629 B.n301 B.n70 10.6151
R630 B.n297 B.n70 10.6151
R631 B.n297 B.n296 10.6151
R632 B.n296 B.n295 10.6151
R633 B.n295 B.n72 10.6151
R634 B.n291 B.n72 10.6151
R635 B.n291 B.n290 10.6151
R636 B.n290 B.n289 10.6151
R637 B.n289 B.n74 10.6151
R638 B.n285 B.n74 10.6151
R639 B.n285 B.n284 10.6151
R640 B.n284 B.n283 10.6151
R641 B.n283 B.n76 10.6151
R642 B.n279 B.n76 10.6151
R643 B.n279 B.n278 10.6151
R644 B.n278 B.n277 10.6151
R645 B.n277 B.n78 10.6151
R646 B.n273 B.n78 10.6151
R647 B.n273 B.n272 10.6151
R648 B.n272 B.n271 10.6151
R649 B.n271 B.n80 10.6151
R650 B.n267 B.n80 10.6151
R651 B.n267 B.n266 10.6151
R652 B.n266 B.n265 10.6151
R653 B.n265 B.n82 10.6151
R654 B.n261 B.n82 10.6151
R655 B.n261 B.n260 10.6151
R656 B.n260 B.n259 10.6151
R657 B.n259 B.n84 10.6151
R658 B.n255 B.n84 10.6151
R659 B.n255 B.n254 10.6151
R660 B.n254 B.n253 10.6151
R661 B.n253 B.n86 10.6151
R662 B.n249 B.n86 10.6151
R663 B.n249 B.n248 10.6151
R664 B.n129 B.n1 10.6151
R665 B.n130 B.n129 10.6151
R666 B.n131 B.n130 10.6151
R667 B.n131 B.n126 10.6151
R668 B.n135 B.n126 10.6151
R669 B.n136 B.n135 10.6151
R670 B.n137 B.n136 10.6151
R671 B.n137 B.n124 10.6151
R672 B.n141 B.n124 10.6151
R673 B.n142 B.n141 10.6151
R674 B.n143 B.n142 10.6151
R675 B.n143 B.n122 10.6151
R676 B.n147 B.n122 10.6151
R677 B.n148 B.n147 10.6151
R678 B.n149 B.n148 10.6151
R679 B.n149 B.n120 10.6151
R680 B.n153 B.n120 10.6151
R681 B.n154 B.n153 10.6151
R682 B.n155 B.n154 10.6151
R683 B.n155 B.n118 10.6151
R684 B.n159 B.n118 10.6151
R685 B.n160 B.n159 10.6151
R686 B.n161 B.n160 10.6151
R687 B.n161 B.n116 10.6151
R688 B.n165 B.n116 10.6151
R689 B.n166 B.n165 10.6151
R690 B.n167 B.n166 10.6151
R691 B.n167 B.n114 10.6151
R692 B.n171 B.n114 10.6151
R693 B.n172 B.n171 10.6151
R694 B.n173 B.n172 10.6151
R695 B.n173 B.n112 10.6151
R696 B.n177 B.n112 10.6151
R697 B.n178 B.n177 10.6151
R698 B.n179 B.n178 10.6151
R699 B.n179 B.n110 10.6151
R700 B.n183 B.n110 10.6151
R701 B.n184 B.n183 10.6151
R702 B.n185 B.n184 10.6151
R703 B.n185 B.n108 10.6151
R704 B.n190 B.n189 10.6151
R705 B.n191 B.n190 10.6151
R706 B.n191 B.n106 10.6151
R707 B.n195 B.n106 10.6151
R708 B.n196 B.n195 10.6151
R709 B.n197 B.n196 10.6151
R710 B.n197 B.n104 10.6151
R711 B.n201 B.n104 10.6151
R712 B.n202 B.n201 10.6151
R713 B.n203 B.n202 10.6151
R714 B.n203 B.n102 10.6151
R715 B.n207 B.n102 10.6151
R716 B.n208 B.n207 10.6151
R717 B.n210 B.n98 10.6151
R718 B.n214 B.n98 10.6151
R719 B.n215 B.n214 10.6151
R720 B.n216 B.n215 10.6151
R721 B.n216 B.n96 10.6151
R722 B.n220 B.n96 10.6151
R723 B.n221 B.n220 10.6151
R724 B.n225 B.n221 10.6151
R725 B.n229 B.n94 10.6151
R726 B.n230 B.n229 10.6151
R727 B.n231 B.n230 10.6151
R728 B.n231 B.n92 10.6151
R729 B.n235 B.n92 10.6151
R730 B.n236 B.n235 10.6151
R731 B.n237 B.n236 10.6151
R732 B.n237 B.n90 10.6151
R733 B.n241 B.n90 10.6151
R734 B.n242 B.n241 10.6151
R735 B.n243 B.n242 10.6151
R736 B.n243 B.n88 10.6151
R737 B.n247 B.n88 10.6151
R738 B.n493 B.n0 8.11757
R739 B.n493 B.n1 8.11757
R740 B.n409 B.n408 6.5566
R741 B.n396 B.n38 6.5566
R742 B.n210 B.n209 6.5566
R743 B.n225 B.n224 6.5566
R744 B.n410 B.n409 4.05904
R745 B.n393 B.n38 4.05904
R746 B.n209 B.n208 4.05904
R747 B.n224 B.n94 4.05904
R748 VN.n29 VN.n16 161.3
R749 VN.n28 VN.n27 161.3
R750 VN.n26 VN.n17 161.3
R751 VN.n25 VN.n24 161.3
R752 VN.n23 VN.n18 161.3
R753 VN.n22 VN.n21 161.3
R754 VN.n13 VN.n0 161.3
R755 VN.n12 VN.n11 161.3
R756 VN.n10 VN.n1 161.3
R757 VN.n9 VN.n8 161.3
R758 VN.n7 VN.n2 161.3
R759 VN.n6 VN.n5 161.3
R760 VN.n15 VN.n14 106.353
R761 VN.n31 VN.n30 106.353
R762 VN.n4 VN.n3 59.8676
R763 VN.n20 VN.n19 59.8676
R764 VN.n8 VN.n1 56.5193
R765 VN.n24 VN.n17 56.5193
R766 VN.n4 VN.t5 55.9455
R767 VN.n20 VN.t1 55.9455
R768 VN VN.n31 41.3239
R769 VN.n7 VN.n6 24.4675
R770 VN.n8 VN.n7 24.4675
R771 VN.n12 VN.n1 24.4675
R772 VN.n13 VN.n12 24.4675
R773 VN.n24 VN.n23 24.4675
R774 VN.n23 VN.n22 24.4675
R775 VN.n29 VN.n28 24.4675
R776 VN.n28 VN.n17 24.4675
R777 VN.n3 VN.t4 24.1005
R778 VN.n14 VN.t2 24.1005
R779 VN.n19 VN.t0 24.1005
R780 VN.n30 VN.t3 24.1005
R781 VN.n6 VN.n3 12.234
R782 VN.n22 VN.n19 12.234
R783 VN.n21 VN.n20 7.20192
R784 VN.n5 VN.n4 7.20192
R785 VN.n14 VN.n13 4.40456
R786 VN.n30 VN.n29 4.40456
R787 VN.n31 VN.n16 0.278367
R788 VN.n15 VN.n0 0.278367
R789 VN.n27 VN.n16 0.189894
R790 VN.n27 VN.n26 0.189894
R791 VN.n26 VN.n25 0.189894
R792 VN.n25 VN.n18 0.189894
R793 VN.n21 VN.n18 0.189894
R794 VN.n5 VN.n2 0.189894
R795 VN.n9 VN.n2 0.189894
R796 VN.n10 VN.n9 0.189894
R797 VN.n11 VN.n10 0.189894
R798 VN.n11 VN.n0 0.189894
R799 VN VN.n15 0.153454
R800 VDD2.n19 VDD2.n13 756.745
R801 VDD2.n6 VDD2.n0 756.745
R802 VDD2.n20 VDD2.n19 585
R803 VDD2.n18 VDD2.n17 585
R804 VDD2.n5 VDD2.n4 585
R805 VDD2.n7 VDD2.n6 585
R806 VDD2.n16 VDD2.t5 355.474
R807 VDD2.n3 VDD2.t3 355.474
R808 VDD2.n19 VDD2.n18 171.744
R809 VDD2.n6 VDD2.n5 171.744
R810 VDD2.n12 VDD2.n11 154.411
R811 VDD2 VDD2.n25 154.407
R812 VDD2.n18 VDD2.t5 85.8723
R813 VDD2.n5 VDD2.t3 85.8723
R814 VDD2.n12 VDD2.n10 52.7783
R815 VDD2.n24 VDD2.n23 50.9975
R816 VDD2.n24 VDD2.n12 33.836
R817 VDD2.n17 VDD2.n16 15.8418
R818 VDD2.n4 VDD2.n3 15.8418
R819 VDD2.n25 VDD2.t1 12.9507
R820 VDD2.n25 VDD2.t0 12.9507
R821 VDD2.n11 VDD2.t4 12.9507
R822 VDD2.n11 VDD2.t2 12.9507
R823 VDD2.n20 VDD2.n15 12.8005
R824 VDD2.n7 VDD2.n2 12.8005
R825 VDD2.n21 VDD2.n13 12.0247
R826 VDD2.n8 VDD2.n0 12.0247
R827 VDD2.n23 VDD2.n22 9.45567
R828 VDD2.n10 VDD2.n9 9.45567
R829 VDD2.n22 VDD2.n21 9.3005
R830 VDD2.n15 VDD2.n14 9.3005
R831 VDD2.n9 VDD2.n8 9.3005
R832 VDD2.n2 VDD2.n1 9.3005
R833 VDD2.n16 VDD2.n14 4.29255
R834 VDD2.n3 VDD2.n1 4.29255
R835 VDD2.n23 VDD2.n13 1.93989
R836 VDD2.n10 VDD2.n0 1.93989
R837 VDD2 VDD2.n24 1.8949
R838 VDD2.n21 VDD2.n20 1.16414
R839 VDD2.n8 VDD2.n7 1.16414
R840 VDD2.n17 VDD2.n15 0.388379
R841 VDD2.n4 VDD2.n2 0.388379
R842 VDD2.n22 VDD2.n14 0.155672
R843 VDD2.n9 VDD2.n1 0.155672
R844 VTAIL.n50 VTAIL.n44 756.745
R845 VTAIL.n8 VTAIL.n2 756.745
R846 VTAIL.n38 VTAIL.n32 756.745
R847 VTAIL.n24 VTAIL.n18 756.745
R848 VTAIL.n49 VTAIL.n48 585
R849 VTAIL.n51 VTAIL.n50 585
R850 VTAIL.n7 VTAIL.n6 585
R851 VTAIL.n9 VTAIL.n8 585
R852 VTAIL.n39 VTAIL.n38 585
R853 VTAIL.n37 VTAIL.n36 585
R854 VTAIL.n25 VTAIL.n24 585
R855 VTAIL.n23 VTAIL.n22 585
R856 VTAIL.n47 VTAIL.t9 355.474
R857 VTAIL.n5 VTAIL.t0 355.474
R858 VTAIL.n35 VTAIL.t4 355.474
R859 VTAIL.n21 VTAIL.t10 355.474
R860 VTAIL.n50 VTAIL.n49 171.744
R861 VTAIL.n8 VTAIL.n7 171.744
R862 VTAIL.n38 VTAIL.n37 171.744
R863 VTAIL.n24 VTAIL.n23 171.744
R864 VTAIL.n31 VTAIL.n30 137.174
R865 VTAIL.n17 VTAIL.n16 137.174
R866 VTAIL.n1 VTAIL.n0 137.174
R867 VTAIL.n15 VTAIL.n14 137.174
R868 VTAIL.n49 VTAIL.t9 85.8723
R869 VTAIL.n7 VTAIL.t0 85.8723
R870 VTAIL.n37 VTAIL.t4 85.8723
R871 VTAIL.n23 VTAIL.t10 85.8723
R872 VTAIL.n55 VTAIL.n54 34.3187
R873 VTAIL.n13 VTAIL.n12 34.3187
R874 VTAIL.n43 VTAIL.n42 34.3187
R875 VTAIL.n29 VTAIL.n28 34.3187
R876 VTAIL.n17 VTAIL.n15 19.4272
R877 VTAIL.n55 VTAIL.n43 16.9789
R878 VTAIL.n48 VTAIL.n47 15.8418
R879 VTAIL.n6 VTAIL.n5 15.8418
R880 VTAIL.n36 VTAIL.n35 15.8418
R881 VTAIL.n22 VTAIL.n21 15.8418
R882 VTAIL.n0 VTAIL.t6 12.9507
R883 VTAIL.n0 VTAIL.t7 12.9507
R884 VTAIL.n14 VTAIL.t3 12.9507
R885 VTAIL.n14 VTAIL.t5 12.9507
R886 VTAIL.n30 VTAIL.t1 12.9507
R887 VTAIL.n30 VTAIL.t2 12.9507
R888 VTAIL.n16 VTAIL.t8 12.9507
R889 VTAIL.n16 VTAIL.t11 12.9507
R890 VTAIL.n51 VTAIL.n46 12.8005
R891 VTAIL.n9 VTAIL.n4 12.8005
R892 VTAIL.n39 VTAIL.n34 12.8005
R893 VTAIL.n25 VTAIL.n20 12.8005
R894 VTAIL.n52 VTAIL.n44 12.0247
R895 VTAIL.n10 VTAIL.n2 12.0247
R896 VTAIL.n40 VTAIL.n32 12.0247
R897 VTAIL.n26 VTAIL.n18 12.0247
R898 VTAIL.n54 VTAIL.n53 9.45567
R899 VTAIL.n12 VTAIL.n11 9.45567
R900 VTAIL.n42 VTAIL.n41 9.45567
R901 VTAIL.n28 VTAIL.n27 9.45567
R902 VTAIL.n53 VTAIL.n52 9.3005
R903 VTAIL.n46 VTAIL.n45 9.3005
R904 VTAIL.n11 VTAIL.n10 9.3005
R905 VTAIL.n4 VTAIL.n3 9.3005
R906 VTAIL.n41 VTAIL.n40 9.3005
R907 VTAIL.n34 VTAIL.n33 9.3005
R908 VTAIL.n27 VTAIL.n26 9.3005
R909 VTAIL.n20 VTAIL.n19 9.3005
R910 VTAIL.n35 VTAIL.n33 4.29255
R911 VTAIL.n21 VTAIL.n19 4.29255
R912 VTAIL.n47 VTAIL.n45 4.29255
R913 VTAIL.n5 VTAIL.n3 4.29255
R914 VTAIL.n29 VTAIL.n17 2.44878
R915 VTAIL.n43 VTAIL.n31 2.44878
R916 VTAIL.n15 VTAIL.n13 2.44878
R917 VTAIL.n54 VTAIL.n44 1.93989
R918 VTAIL.n12 VTAIL.n2 1.93989
R919 VTAIL.n42 VTAIL.n32 1.93989
R920 VTAIL.n28 VTAIL.n18 1.93989
R921 VTAIL VTAIL.n55 1.77852
R922 VTAIL.n31 VTAIL.n29 1.69447
R923 VTAIL.n13 VTAIL.n1 1.69447
R924 VTAIL.n52 VTAIL.n51 1.16414
R925 VTAIL.n10 VTAIL.n9 1.16414
R926 VTAIL.n40 VTAIL.n39 1.16414
R927 VTAIL.n26 VTAIL.n25 1.16414
R928 VTAIL VTAIL.n1 0.670759
R929 VTAIL.n48 VTAIL.n46 0.388379
R930 VTAIL.n6 VTAIL.n4 0.388379
R931 VTAIL.n36 VTAIL.n34 0.388379
R932 VTAIL.n22 VTAIL.n20 0.388379
R933 VTAIL.n53 VTAIL.n45 0.155672
R934 VTAIL.n11 VTAIL.n3 0.155672
R935 VTAIL.n41 VTAIL.n33 0.155672
R936 VTAIL.n27 VTAIL.n19 0.155672
R937 VP.n13 VP.n12 161.3
R938 VP.n14 VP.n9 161.3
R939 VP.n16 VP.n15 161.3
R940 VP.n17 VP.n8 161.3
R941 VP.n19 VP.n18 161.3
R942 VP.n20 VP.n7 161.3
R943 VP.n42 VP.n0 161.3
R944 VP.n41 VP.n40 161.3
R945 VP.n39 VP.n1 161.3
R946 VP.n38 VP.n37 161.3
R947 VP.n36 VP.n2 161.3
R948 VP.n35 VP.n34 161.3
R949 VP.n33 VP.n32 161.3
R950 VP.n31 VP.n4 161.3
R951 VP.n30 VP.n29 161.3
R952 VP.n28 VP.n5 161.3
R953 VP.n27 VP.n26 161.3
R954 VP.n25 VP.n6 161.3
R955 VP.n24 VP.n23 106.353
R956 VP.n44 VP.n43 106.353
R957 VP.n22 VP.n21 106.353
R958 VP.n11 VP.n10 59.8676
R959 VP.n30 VP.n5 56.5193
R960 VP.n37 VP.n1 56.5193
R961 VP.n15 VP.n8 56.5193
R962 VP.n11 VP.t3 55.9455
R963 VP.n23 VP.n22 41.045
R964 VP.n26 VP.n25 24.4675
R965 VP.n26 VP.n5 24.4675
R966 VP.n31 VP.n30 24.4675
R967 VP.n32 VP.n31 24.4675
R968 VP.n36 VP.n35 24.4675
R969 VP.n37 VP.n36 24.4675
R970 VP.n41 VP.n1 24.4675
R971 VP.n42 VP.n41 24.4675
R972 VP.n19 VP.n8 24.4675
R973 VP.n20 VP.n19 24.4675
R974 VP.n14 VP.n13 24.4675
R975 VP.n15 VP.n14 24.4675
R976 VP.n24 VP.t5 24.1005
R977 VP.n3 VP.t0 24.1005
R978 VP.n43 VP.t2 24.1005
R979 VP.n21 VP.t1 24.1005
R980 VP.n10 VP.t4 24.1005
R981 VP.n32 VP.n3 12.234
R982 VP.n35 VP.n3 12.234
R983 VP.n13 VP.n10 12.234
R984 VP.n12 VP.n11 7.20192
R985 VP.n25 VP.n24 4.40456
R986 VP.n43 VP.n42 4.40456
R987 VP.n21 VP.n20 4.40456
R988 VP.n22 VP.n7 0.278367
R989 VP.n23 VP.n6 0.278367
R990 VP.n44 VP.n0 0.278367
R991 VP.n12 VP.n9 0.189894
R992 VP.n16 VP.n9 0.189894
R993 VP.n17 VP.n16 0.189894
R994 VP.n18 VP.n17 0.189894
R995 VP.n18 VP.n7 0.189894
R996 VP.n27 VP.n6 0.189894
R997 VP.n28 VP.n27 0.189894
R998 VP.n29 VP.n28 0.189894
R999 VP.n29 VP.n4 0.189894
R1000 VP.n33 VP.n4 0.189894
R1001 VP.n34 VP.n33 0.189894
R1002 VP.n34 VP.n2 0.189894
R1003 VP.n38 VP.n2 0.189894
R1004 VP.n39 VP.n38 0.189894
R1005 VP.n40 VP.n39 0.189894
R1006 VP.n40 VP.n0 0.189894
R1007 VP VP.n44 0.153454
R1008 VDD1.n6 VDD1.n0 756.745
R1009 VDD1.n17 VDD1.n11 756.745
R1010 VDD1.n7 VDD1.n6 585
R1011 VDD1.n5 VDD1.n4 585
R1012 VDD1.n16 VDD1.n15 585
R1013 VDD1.n18 VDD1.n17 585
R1014 VDD1.n3 VDD1.t2 355.474
R1015 VDD1.n14 VDD1.t0 355.474
R1016 VDD1.n6 VDD1.n5 171.744
R1017 VDD1.n17 VDD1.n16 171.744
R1018 VDD1.n23 VDD1.n22 154.411
R1019 VDD1.n25 VDD1.n24 153.853
R1020 VDD1.n5 VDD1.t2 85.8723
R1021 VDD1.n16 VDD1.t0 85.8723
R1022 VDD1 VDD1.n10 52.8919
R1023 VDD1.n23 VDD1.n21 52.7783
R1024 VDD1.n25 VDD1.n23 35.6431
R1025 VDD1.n4 VDD1.n3 15.8418
R1026 VDD1.n15 VDD1.n14 15.8418
R1027 VDD1.n24 VDD1.t1 12.9507
R1028 VDD1.n24 VDD1.t4 12.9507
R1029 VDD1.n22 VDD1.t5 12.9507
R1030 VDD1.n22 VDD1.t3 12.9507
R1031 VDD1.n7 VDD1.n2 12.8005
R1032 VDD1.n18 VDD1.n13 12.8005
R1033 VDD1.n8 VDD1.n0 12.0247
R1034 VDD1.n19 VDD1.n11 12.0247
R1035 VDD1.n10 VDD1.n9 9.45567
R1036 VDD1.n21 VDD1.n20 9.45567
R1037 VDD1.n9 VDD1.n8 9.3005
R1038 VDD1.n2 VDD1.n1 9.3005
R1039 VDD1.n20 VDD1.n19 9.3005
R1040 VDD1.n13 VDD1.n12 9.3005
R1041 VDD1.n3 VDD1.n1 4.29255
R1042 VDD1.n14 VDD1.n12 4.29255
R1043 VDD1.n10 VDD1.n0 1.93989
R1044 VDD1.n21 VDD1.n11 1.93989
R1045 VDD1.n8 VDD1.n7 1.16414
R1046 VDD1.n19 VDD1.n18 1.16414
R1047 VDD1 VDD1.n25 0.554379
R1048 VDD1.n4 VDD1.n2 0.388379
R1049 VDD1.n15 VDD1.n13 0.388379
R1050 VDD1.n9 VDD1.n1 0.155672
R1051 VDD1.n20 VDD1.n12 0.155672
C0 VP VN 5.09276f
C1 VDD2 w_n3242_n1470# 1.68762f
C2 VP VDD2 0.456548f
C3 VN VDD1 0.156391f
C4 B w_n3242_n1470# 6.92058f
C5 B VP 1.73328f
C6 VTAIL VN 2.47235f
C7 VDD2 VDD1 1.37135f
C8 B VDD1 1.31956f
C9 VTAIL VDD2 4.27896f
C10 VP w_n3242_n1470# 6.36572f
C11 B VTAIL 1.47006f
C12 VDD1 w_n3242_n1470# 1.60607f
C13 VP VDD1 1.99787f
C14 VTAIL w_n3242_n1470# 1.60484f
C15 VTAIL VP 2.4865f
C16 VDD2 VN 1.70027f
C17 B VN 1.03491f
C18 VTAIL VDD1 4.22655f
C19 B VDD2 1.39176f
C20 VN w_n3242_n1470# 5.95003f
C21 VDD2 VSUBS 1.052798f
C22 VDD1 VSUBS 1.313736f
C23 VTAIL VSUBS 0.534388f
C24 VN VSUBS 5.42229f
C25 VP VSUBS 2.302525f
C26 B VSUBS 3.526675f
C27 w_n3242_n1470# VSUBS 60.5735f
C28 VDD1.n0 VSUBS 0.016461f
C29 VDD1.n1 VSUBS 0.110492f
C30 VDD1.n2 VSUBS 0.008373f
C31 VDD1.t2 VSUBS 0.044228f
C32 VDD1.n3 VSUBS 0.051938f
C33 VDD1.n4 VSUBS 0.011669f
C34 VDD1.n5 VSUBS 0.014843f
C35 VDD1.n6 VSUBS 0.045663f
C36 VDD1.n7 VSUBS 0.008865f
C37 VDD1.n8 VSUBS 0.008373f
C38 VDD1.n9 VSUBS 0.038357f
C39 VDD1.n10 VSUBS 0.038204f
C40 VDD1.n11 VSUBS 0.016461f
C41 VDD1.n12 VSUBS 0.110492f
C42 VDD1.n13 VSUBS 0.008373f
C43 VDD1.t0 VSUBS 0.044228f
C44 VDD1.n14 VSUBS 0.051938f
C45 VDD1.n15 VSUBS 0.011669f
C46 VDD1.n16 VSUBS 0.014843f
C47 VDD1.n17 VSUBS 0.045663f
C48 VDD1.n18 VSUBS 0.008865f
C49 VDD1.n19 VSUBS 0.008373f
C50 VDD1.n20 VSUBS 0.038357f
C51 VDD1.n21 VSUBS 0.037757f
C52 VDD1.t5 VSUBS 0.030905f
C53 VDD1.t3 VSUBS 0.030905f
C54 VDD1.n22 VSUBS 0.152342f
C55 VDD1.n23 VSUBS 1.41856f
C56 VDD1.t1 VSUBS 0.030905f
C57 VDD1.t4 VSUBS 0.030905f
C58 VDD1.n24 VSUBS 0.151114f
C59 VDD1.n25 VSUBS 1.31503f
C60 VP.n0 VSUBS 0.062598f
C61 VP.t2 VSUBS 0.726979f
C62 VP.n1 VSUBS 0.079898f
C63 VP.n2 VSUBS 0.04748f
C64 VP.t0 VSUBS 0.726979f
C65 VP.n3 VSUBS 0.323125f
C66 VP.n4 VSUBS 0.04748f
C67 VP.n5 VSUBS 0.079898f
C68 VP.n6 VSUBS 0.062598f
C69 VP.t5 VSUBS 0.726979f
C70 VP.n7 VSUBS 0.062598f
C71 VP.t1 VSUBS 0.726979f
C72 VP.n8 VSUBS 0.079898f
C73 VP.n9 VSUBS 0.04748f
C74 VP.t4 VSUBS 0.726979f
C75 VP.n10 VSUBS 0.457082f
C76 VP.t3 VSUBS 1.07194f
C77 VP.n11 VSUBS 0.444197f
C78 VP.n12 VSUBS 0.453545f
C79 VP.n13 VSUBS 0.066647f
C80 VP.n14 VSUBS 0.088492f
C81 VP.n15 VSUBS 0.058728f
C82 VP.n16 VSUBS 0.04748f
C83 VP.n17 VSUBS 0.04748f
C84 VP.n18 VSUBS 0.04748f
C85 VP.n19 VSUBS 0.088492f
C86 VP.n20 VSUBS 0.052667f
C87 VP.n21 VSUBS 0.46258f
C88 VP.n22 VSUBS 1.94847f
C89 VP.n23 VSUBS 1.99005f
C90 VP.n24 VSUBS 0.46258f
C91 VP.n25 VSUBS 0.052667f
C92 VP.n26 VSUBS 0.088492f
C93 VP.n27 VSUBS 0.04748f
C94 VP.n28 VSUBS 0.04748f
C95 VP.n29 VSUBS 0.04748f
C96 VP.n30 VSUBS 0.058728f
C97 VP.n31 VSUBS 0.088492f
C98 VP.n32 VSUBS 0.066647f
C99 VP.n33 VSUBS 0.04748f
C100 VP.n34 VSUBS 0.04748f
C101 VP.n35 VSUBS 0.066647f
C102 VP.n36 VSUBS 0.088492f
C103 VP.n37 VSUBS 0.058728f
C104 VP.n38 VSUBS 0.04748f
C105 VP.n39 VSUBS 0.04748f
C106 VP.n40 VSUBS 0.04748f
C107 VP.n41 VSUBS 0.088492f
C108 VP.n42 VSUBS 0.052667f
C109 VP.n43 VSUBS 0.46258f
C110 VP.n44 VSUBS 0.081717f
C111 VTAIL.t6 VSUBS 0.064918f
C112 VTAIL.t7 VSUBS 0.064918f
C113 VTAIL.n0 VSUBS 0.271541f
C114 VTAIL.n1 VSUBS 0.63429f
C115 VTAIL.n2 VSUBS 0.034577f
C116 VTAIL.n3 VSUBS 0.232091f
C117 VTAIL.n4 VSUBS 0.017587f
C118 VTAIL.t0 VSUBS 0.092901f
C119 VTAIL.n5 VSUBS 0.109098f
C120 VTAIL.n6 VSUBS 0.024511f
C121 VTAIL.n7 VSUBS 0.031177f
C122 VTAIL.n8 VSUBS 0.095917f
C123 VTAIL.n9 VSUBS 0.018622f
C124 VTAIL.n10 VSUBS 0.017587f
C125 VTAIL.n11 VSUBS 0.08057f
C126 VTAIL.n12 VSUBS 0.048173f
C127 VTAIL.n13 VSUBS 0.467578f
C128 VTAIL.t3 VSUBS 0.064918f
C129 VTAIL.t5 VSUBS 0.064918f
C130 VTAIL.n14 VSUBS 0.271541f
C131 VTAIL.n15 VSUBS 1.83233f
C132 VTAIL.t8 VSUBS 0.064918f
C133 VTAIL.t11 VSUBS 0.064918f
C134 VTAIL.n16 VSUBS 0.271543f
C135 VTAIL.n17 VSUBS 1.83233f
C136 VTAIL.n18 VSUBS 0.034577f
C137 VTAIL.n19 VSUBS 0.232091f
C138 VTAIL.n20 VSUBS 0.017587f
C139 VTAIL.t10 VSUBS 0.092901f
C140 VTAIL.n21 VSUBS 0.109098f
C141 VTAIL.n22 VSUBS 0.024511f
C142 VTAIL.n23 VSUBS 0.031177f
C143 VTAIL.n24 VSUBS 0.095917f
C144 VTAIL.n25 VSUBS 0.018622f
C145 VTAIL.n26 VSUBS 0.017587f
C146 VTAIL.n27 VSUBS 0.08057f
C147 VTAIL.n28 VSUBS 0.048173f
C148 VTAIL.n29 VSUBS 0.467578f
C149 VTAIL.t1 VSUBS 0.064918f
C150 VTAIL.t2 VSUBS 0.064918f
C151 VTAIL.n30 VSUBS 0.271543f
C152 VTAIL.n31 VSUBS 0.821799f
C153 VTAIL.n32 VSUBS 0.034577f
C154 VTAIL.n33 VSUBS 0.232091f
C155 VTAIL.n34 VSUBS 0.017587f
C156 VTAIL.t4 VSUBS 0.092901f
C157 VTAIL.n35 VSUBS 0.109098f
C158 VTAIL.n36 VSUBS 0.024511f
C159 VTAIL.n37 VSUBS 0.031177f
C160 VTAIL.n38 VSUBS 0.095917f
C161 VTAIL.n39 VSUBS 0.018622f
C162 VTAIL.n40 VSUBS 0.017587f
C163 VTAIL.n41 VSUBS 0.08057f
C164 VTAIL.n42 VSUBS 0.048173f
C165 VTAIL.n43 VSUBS 1.21991f
C166 VTAIL.n44 VSUBS 0.034577f
C167 VTAIL.n45 VSUBS 0.232091f
C168 VTAIL.n46 VSUBS 0.017587f
C169 VTAIL.t9 VSUBS 0.092901f
C170 VTAIL.n47 VSUBS 0.109098f
C171 VTAIL.n48 VSUBS 0.024511f
C172 VTAIL.n49 VSUBS 0.031177f
C173 VTAIL.n50 VSUBS 0.095917f
C174 VTAIL.n51 VSUBS 0.018622f
C175 VTAIL.n52 VSUBS 0.017587f
C176 VTAIL.n53 VSUBS 0.08057f
C177 VTAIL.n54 VSUBS 0.048173f
C178 VTAIL.n55 VSUBS 1.14923f
C179 VDD2.n0 VSUBS 0.017087f
C180 VDD2.n1 VSUBS 0.114694f
C181 VDD2.n2 VSUBS 0.008691f
C182 VDD2.t3 VSUBS 0.04591f
C183 VDD2.n3 VSUBS 0.053914f
C184 VDD2.n4 VSUBS 0.012113f
C185 VDD2.n5 VSUBS 0.015407f
C186 VDD2.n6 VSUBS 0.0474f
C187 VDD2.n7 VSUBS 0.009202f
C188 VDD2.n8 VSUBS 0.008691f
C189 VDD2.n9 VSUBS 0.039816f
C190 VDD2.n10 VSUBS 0.039193f
C191 VDD2.t4 VSUBS 0.032081f
C192 VDD2.t2 VSUBS 0.032081f
C193 VDD2.n11 VSUBS 0.158136f
C194 VDD2.n12 VSUBS 1.40005f
C195 VDD2.n13 VSUBS 0.017087f
C196 VDD2.n14 VSUBS 0.114694f
C197 VDD2.n15 VSUBS 0.008691f
C198 VDD2.t5 VSUBS 0.04591f
C199 VDD2.n16 VSUBS 0.053914f
C200 VDD2.n17 VSUBS 0.012113f
C201 VDD2.n18 VSUBS 0.015407f
C202 VDD2.n19 VSUBS 0.0474f
C203 VDD2.n20 VSUBS 0.009202f
C204 VDD2.n21 VSUBS 0.008691f
C205 VDD2.n22 VSUBS 0.039816f
C206 VDD2.n23 VSUBS 0.034956f
C207 VDD2.n24 VSUBS 1.15651f
C208 VDD2.t1 VSUBS 0.032081f
C209 VDD2.t0 VSUBS 0.032081f
C210 VDD2.n25 VSUBS 0.158126f
C211 VN.n0 VSUBS 0.060521f
C212 VN.t2 VSUBS 0.702857f
C213 VN.n1 VSUBS 0.077247f
C214 VN.n2 VSUBS 0.045905f
C215 VN.t4 VSUBS 0.702857f
C216 VN.n3 VSUBS 0.441916f
C217 VN.t5 VSUBS 1.03637f
C218 VN.n4 VSUBS 0.429458f
C219 VN.n5 VSUBS 0.438496f
C220 VN.n6 VSUBS 0.064436f
C221 VN.n7 VSUBS 0.085555f
C222 VN.n8 VSUBS 0.05678f
C223 VN.n9 VSUBS 0.045905f
C224 VN.n10 VSUBS 0.045905f
C225 VN.n11 VSUBS 0.045905f
C226 VN.n12 VSUBS 0.085555f
C227 VN.n13 VSUBS 0.050919f
C228 VN.n14 VSUBS 0.447231f
C229 VN.n15 VSUBS 0.079005f
C230 VN.n16 VSUBS 0.060521f
C231 VN.t3 VSUBS 0.702857f
C232 VN.n17 VSUBS 0.077247f
C233 VN.n18 VSUBS 0.045905f
C234 VN.t0 VSUBS 0.702857f
C235 VN.n19 VSUBS 0.441916f
C236 VN.t1 VSUBS 1.03637f
C237 VN.n20 VSUBS 0.429458f
C238 VN.n21 VSUBS 0.438496f
C239 VN.n22 VSUBS 0.064436f
C240 VN.n23 VSUBS 0.085555f
C241 VN.n24 VSUBS 0.05678f
C242 VN.n25 VSUBS 0.045905f
C243 VN.n26 VSUBS 0.045905f
C244 VN.n27 VSUBS 0.045905f
C245 VN.n28 VSUBS 0.085555f
C246 VN.n29 VSUBS 0.050919f
C247 VN.n30 VSUBS 0.447231f
C248 VN.n31 VSUBS 1.90934f
C249 B.n0 VSUBS 0.007226f
C250 B.n1 VSUBS 0.007226f
C251 B.n2 VSUBS 0.010687f
C252 B.n3 VSUBS 0.008189f
C253 B.n4 VSUBS 0.008189f
C254 B.n5 VSUBS 0.008189f
C255 B.n6 VSUBS 0.008189f
C256 B.n7 VSUBS 0.008189f
C257 B.n8 VSUBS 0.008189f
C258 B.n9 VSUBS 0.008189f
C259 B.n10 VSUBS 0.008189f
C260 B.n11 VSUBS 0.008189f
C261 B.n12 VSUBS 0.008189f
C262 B.n13 VSUBS 0.008189f
C263 B.n14 VSUBS 0.008189f
C264 B.n15 VSUBS 0.008189f
C265 B.n16 VSUBS 0.008189f
C266 B.n17 VSUBS 0.008189f
C267 B.n18 VSUBS 0.008189f
C268 B.n19 VSUBS 0.008189f
C269 B.n20 VSUBS 0.008189f
C270 B.n21 VSUBS 0.008189f
C271 B.n22 VSUBS 0.018665f
C272 B.n23 VSUBS 0.008189f
C273 B.n24 VSUBS 0.008189f
C274 B.n25 VSUBS 0.008189f
C275 B.n26 VSUBS 0.008189f
C276 B.n27 VSUBS 0.008189f
C277 B.n28 VSUBS 0.008189f
C278 B.n29 VSUBS 0.008189f
C279 B.t4 VSUBS 0.045522f
C280 B.t5 VSUBS 0.06177f
C281 B.t3 VSUBS 0.36026f
C282 B.n30 VSUBS 0.109995f
C283 B.n31 VSUBS 0.094138f
C284 B.n32 VSUBS 0.008189f
C285 B.n33 VSUBS 0.008189f
C286 B.n34 VSUBS 0.008189f
C287 B.n35 VSUBS 0.008189f
C288 B.t1 VSUBS 0.045523f
C289 B.t2 VSUBS 0.06177f
C290 B.t0 VSUBS 0.36026f
C291 B.n36 VSUBS 0.109995f
C292 B.n37 VSUBS 0.094137f
C293 B.n38 VSUBS 0.018974f
C294 B.n39 VSUBS 0.008189f
C295 B.n40 VSUBS 0.008189f
C296 B.n41 VSUBS 0.008189f
C297 B.n42 VSUBS 0.008189f
C298 B.n43 VSUBS 0.008189f
C299 B.n44 VSUBS 0.008189f
C300 B.n45 VSUBS 0.019633f
C301 B.n46 VSUBS 0.008189f
C302 B.n47 VSUBS 0.008189f
C303 B.n48 VSUBS 0.008189f
C304 B.n49 VSUBS 0.008189f
C305 B.n50 VSUBS 0.008189f
C306 B.n51 VSUBS 0.008189f
C307 B.n52 VSUBS 0.008189f
C308 B.n53 VSUBS 0.008189f
C309 B.n54 VSUBS 0.008189f
C310 B.n55 VSUBS 0.008189f
C311 B.n56 VSUBS 0.008189f
C312 B.n57 VSUBS 0.008189f
C313 B.n58 VSUBS 0.008189f
C314 B.n59 VSUBS 0.008189f
C315 B.n60 VSUBS 0.008189f
C316 B.n61 VSUBS 0.008189f
C317 B.n62 VSUBS 0.008189f
C318 B.n63 VSUBS 0.008189f
C319 B.n64 VSUBS 0.008189f
C320 B.n65 VSUBS 0.008189f
C321 B.n66 VSUBS 0.008189f
C322 B.n67 VSUBS 0.008189f
C323 B.n68 VSUBS 0.008189f
C324 B.n69 VSUBS 0.008189f
C325 B.n70 VSUBS 0.008189f
C326 B.n71 VSUBS 0.008189f
C327 B.n72 VSUBS 0.008189f
C328 B.n73 VSUBS 0.008189f
C329 B.n74 VSUBS 0.008189f
C330 B.n75 VSUBS 0.008189f
C331 B.n76 VSUBS 0.008189f
C332 B.n77 VSUBS 0.008189f
C333 B.n78 VSUBS 0.008189f
C334 B.n79 VSUBS 0.008189f
C335 B.n80 VSUBS 0.008189f
C336 B.n81 VSUBS 0.008189f
C337 B.n82 VSUBS 0.008189f
C338 B.n83 VSUBS 0.008189f
C339 B.n84 VSUBS 0.008189f
C340 B.n85 VSUBS 0.008189f
C341 B.n86 VSUBS 0.008189f
C342 B.n87 VSUBS 0.018665f
C343 B.n88 VSUBS 0.008189f
C344 B.n89 VSUBS 0.008189f
C345 B.n90 VSUBS 0.008189f
C346 B.n91 VSUBS 0.008189f
C347 B.n92 VSUBS 0.008189f
C348 B.n93 VSUBS 0.008189f
C349 B.n94 VSUBS 0.00566f
C350 B.n95 VSUBS 0.008189f
C351 B.n96 VSUBS 0.008189f
C352 B.n97 VSUBS 0.008189f
C353 B.n98 VSUBS 0.008189f
C354 B.n99 VSUBS 0.008189f
C355 B.t11 VSUBS 0.045522f
C356 B.t10 VSUBS 0.06177f
C357 B.t9 VSUBS 0.36026f
C358 B.n100 VSUBS 0.109995f
C359 B.n101 VSUBS 0.094138f
C360 B.n102 VSUBS 0.008189f
C361 B.n103 VSUBS 0.008189f
C362 B.n104 VSUBS 0.008189f
C363 B.n105 VSUBS 0.008189f
C364 B.n106 VSUBS 0.008189f
C365 B.n107 VSUBS 0.008189f
C366 B.n108 VSUBS 0.018665f
C367 B.n109 VSUBS 0.008189f
C368 B.n110 VSUBS 0.008189f
C369 B.n111 VSUBS 0.008189f
C370 B.n112 VSUBS 0.008189f
C371 B.n113 VSUBS 0.008189f
C372 B.n114 VSUBS 0.008189f
C373 B.n115 VSUBS 0.008189f
C374 B.n116 VSUBS 0.008189f
C375 B.n117 VSUBS 0.008189f
C376 B.n118 VSUBS 0.008189f
C377 B.n119 VSUBS 0.008189f
C378 B.n120 VSUBS 0.008189f
C379 B.n121 VSUBS 0.008189f
C380 B.n122 VSUBS 0.008189f
C381 B.n123 VSUBS 0.008189f
C382 B.n124 VSUBS 0.008189f
C383 B.n125 VSUBS 0.008189f
C384 B.n126 VSUBS 0.008189f
C385 B.n127 VSUBS 0.008189f
C386 B.n128 VSUBS 0.008189f
C387 B.n129 VSUBS 0.008189f
C388 B.n130 VSUBS 0.008189f
C389 B.n131 VSUBS 0.008189f
C390 B.n132 VSUBS 0.008189f
C391 B.n133 VSUBS 0.008189f
C392 B.n134 VSUBS 0.008189f
C393 B.n135 VSUBS 0.008189f
C394 B.n136 VSUBS 0.008189f
C395 B.n137 VSUBS 0.008189f
C396 B.n138 VSUBS 0.008189f
C397 B.n139 VSUBS 0.008189f
C398 B.n140 VSUBS 0.008189f
C399 B.n141 VSUBS 0.008189f
C400 B.n142 VSUBS 0.008189f
C401 B.n143 VSUBS 0.008189f
C402 B.n144 VSUBS 0.008189f
C403 B.n145 VSUBS 0.008189f
C404 B.n146 VSUBS 0.008189f
C405 B.n147 VSUBS 0.008189f
C406 B.n148 VSUBS 0.008189f
C407 B.n149 VSUBS 0.008189f
C408 B.n150 VSUBS 0.008189f
C409 B.n151 VSUBS 0.008189f
C410 B.n152 VSUBS 0.008189f
C411 B.n153 VSUBS 0.008189f
C412 B.n154 VSUBS 0.008189f
C413 B.n155 VSUBS 0.008189f
C414 B.n156 VSUBS 0.008189f
C415 B.n157 VSUBS 0.008189f
C416 B.n158 VSUBS 0.008189f
C417 B.n159 VSUBS 0.008189f
C418 B.n160 VSUBS 0.008189f
C419 B.n161 VSUBS 0.008189f
C420 B.n162 VSUBS 0.008189f
C421 B.n163 VSUBS 0.008189f
C422 B.n164 VSUBS 0.008189f
C423 B.n165 VSUBS 0.008189f
C424 B.n166 VSUBS 0.008189f
C425 B.n167 VSUBS 0.008189f
C426 B.n168 VSUBS 0.008189f
C427 B.n169 VSUBS 0.008189f
C428 B.n170 VSUBS 0.008189f
C429 B.n171 VSUBS 0.008189f
C430 B.n172 VSUBS 0.008189f
C431 B.n173 VSUBS 0.008189f
C432 B.n174 VSUBS 0.008189f
C433 B.n175 VSUBS 0.008189f
C434 B.n176 VSUBS 0.008189f
C435 B.n177 VSUBS 0.008189f
C436 B.n178 VSUBS 0.008189f
C437 B.n179 VSUBS 0.008189f
C438 B.n180 VSUBS 0.008189f
C439 B.n181 VSUBS 0.008189f
C440 B.n182 VSUBS 0.008189f
C441 B.n183 VSUBS 0.008189f
C442 B.n184 VSUBS 0.008189f
C443 B.n185 VSUBS 0.008189f
C444 B.n186 VSUBS 0.008189f
C445 B.n187 VSUBS 0.018665f
C446 B.n188 VSUBS 0.019633f
C447 B.n189 VSUBS 0.019633f
C448 B.n190 VSUBS 0.008189f
C449 B.n191 VSUBS 0.008189f
C450 B.n192 VSUBS 0.008189f
C451 B.n193 VSUBS 0.008189f
C452 B.n194 VSUBS 0.008189f
C453 B.n195 VSUBS 0.008189f
C454 B.n196 VSUBS 0.008189f
C455 B.n197 VSUBS 0.008189f
C456 B.n198 VSUBS 0.008189f
C457 B.n199 VSUBS 0.008189f
C458 B.n200 VSUBS 0.008189f
C459 B.n201 VSUBS 0.008189f
C460 B.n202 VSUBS 0.008189f
C461 B.n203 VSUBS 0.008189f
C462 B.n204 VSUBS 0.008189f
C463 B.n205 VSUBS 0.008189f
C464 B.n206 VSUBS 0.008189f
C465 B.n207 VSUBS 0.008189f
C466 B.n208 VSUBS 0.00566f
C467 B.n209 VSUBS 0.018974f
C468 B.n210 VSUBS 0.006624f
C469 B.n211 VSUBS 0.008189f
C470 B.n212 VSUBS 0.008189f
C471 B.n213 VSUBS 0.008189f
C472 B.n214 VSUBS 0.008189f
C473 B.n215 VSUBS 0.008189f
C474 B.n216 VSUBS 0.008189f
C475 B.n217 VSUBS 0.008189f
C476 B.n218 VSUBS 0.008189f
C477 B.n219 VSUBS 0.008189f
C478 B.n220 VSUBS 0.008189f
C479 B.n221 VSUBS 0.008189f
C480 B.t8 VSUBS 0.045523f
C481 B.t7 VSUBS 0.06177f
C482 B.t6 VSUBS 0.36026f
C483 B.n222 VSUBS 0.109995f
C484 B.n223 VSUBS 0.094137f
C485 B.n224 VSUBS 0.018974f
C486 B.n225 VSUBS 0.006624f
C487 B.n226 VSUBS 0.008189f
C488 B.n227 VSUBS 0.008189f
C489 B.n228 VSUBS 0.008189f
C490 B.n229 VSUBS 0.008189f
C491 B.n230 VSUBS 0.008189f
C492 B.n231 VSUBS 0.008189f
C493 B.n232 VSUBS 0.008189f
C494 B.n233 VSUBS 0.008189f
C495 B.n234 VSUBS 0.008189f
C496 B.n235 VSUBS 0.008189f
C497 B.n236 VSUBS 0.008189f
C498 B.n237 VSUBS 0.008189f
C499 B.n238 VSUBS 0.008189f
C500 B.n239 VSUBS 0.008189f
C501 B.n240 VSUBS 0.008189f
C502 B.n241 VSUBS 0.008189f
C503 B.n242 VSUBS 0.008189f
C504 B.n243 VSUBS 0.008189f
C505 B.n244 VSUBS 0.008189f
C506 B.n245 VSUBS 0.008189f
C507 B.n246 VSUBS 0.019633f
C508 B.n247 VSUBS 0.018665f
C509 B.n248 VSUBS 0.019633f
C510 B.n249 VSUBS 0.008189f
C511 B.n250 VSUBS 0.008189f
C512 B.n251 VSUBS 0.008189f
C513 B.n252 VSUBS 0.008189f
C514 B.n253 VSUBS 0.008189f
C515 B.n254 VSUBS 0.008189f
C516 B.n255 VSUBS 0.008189f
C517 B.n256 VSUBS 0.008189f
C518 B.n257 VSUBS 0.008189f
C519 B.n258 VSUBS 0.008189f
C520 B.n259 VSUBS 0.008189f
C521 B.n260 VSUBS 0.008189f
C522 B.n261 VSUBS 0.008189f
C523 B.n262 VSUBS 0.008189f
C524 B.n263 VSUBS 0.008189f
C525 B.n264 VSUBS 0.008189f
C526 B.n265 VSUBS 0.008189f
C527 B.n266 VSUBS 0.008189f
C528 B.n267 VSUBS 0.008189f
C529 B.n268 VSUBS 0.008189f
C530 B.n269 VSUBS 0.008189f
C531 B.n270 VSUBS 0.008189f
C532 B.n271 VSUBS 0.008189f
C533 B.n272 VSUBS 0.008189f
C534 B.n273 VSUBS 0.008189f
C535 B.n274 VSUBS 0.008189f
C536 B.n275 VSUBS 0.008189f
C537 B.n276 VSUBS 0.008189f
C538 B.n277 VSUBS 0.008189f
C539 B.n278 VSUBS 0.008189f
C540 B.n279 VSUBS 0.008189f
C541 B.n280 VSUBS 0.008189f
C542 B.n281 VSUBS 0.008189f
C543 B.n282 VSUBS 0.008189f
C544 B.n283 VSUBS 0.008189f
C545 B.n284 VSUBS 0.008189f
C546 B.n285 VSUBS 0.008189f
C547 B.n286 VSUBS 0.008189f
C548 B.n287 VSUBS 0.008189f
C549 B.n288 VSUBS 0.008189f
C550 B.n289 VSUBS 0.008189f
C551 B.n290 VSUBS 0.008189f
C552 B.n291 VSUBS 0.008189f
C553 B.n292 VSUBS 0.008189f
C554 B.n293 VSUBS 0.008189f
C555 B.n294 VSUBS 0.008189f
C556 B.n295 VSUBS 0.008189f
C557 B.n296 VSUBS 0.008189f
C558 B.n297 VSUBS 0.008189f
C559 B.n298 VSUBS 0.008189f
C560 B.n299 VSUBS 0.008189f
C561 B.n300 VSUBS 0.008189f
C562 B.n301 VSUBS 0.008189f
C563 B.n302 VSUBS 0.008189f
C564 B.n303 VSUBS 0.008189f
C565 B.n304 VSUBS 0.008189f
C566 B.n305 VSUBS 0.008189f
C567 B.n306 VSUBS 0.008189f
C568 B.n307 VSUBS 0.008189f
C569 B.n308 VSUBS 0.008189f
C570 B.n309 VSUBS 0.008189f
C571 B.n310 VSUBS 0.008189f
C572 B.n311 VSUBS 0.008189f
C573 B.n312 VSUBS 0.008189f
C574 B.n313 VSUBS 0.008189f
C575 B.n314 VSUBS 0.008189f
C576 B.n315 VSUBS 0.008189f
C577 B.n316 VSUBS 0.008189f
C578 B.n317 VSUBS 0.008189f
C579 B.n318 VSUBS 0.008189f
C580 B.n319 VSUBS 0.008189f
C581 B.n320 VSUBS 0.008189f
C582 B.n321 VSUBS 0.008189f
C583 B.n322 VSUBS 0.008189f
C584 B.n323 VSUBS 0.008189f
C585 B.n324 VSUBS 0.008189f
C586 B.n325 VSUBS 0.008189f
C587 B.n326 VSUBS 0.008189f
C588 B.n327 VSUBS 0.008189f
C589 B.n328 VSUBS 0.008189f
C590 B.n329 VSUBS 0.008189f
C591 B.n330 VSUBS 0.008189f
C592 B.n331 VSUBS 0.008189f
C593 B.n332 VSUBS 0.008189f
C594 B.n333 VSUBS 0.008189f
C595 B.n334 VSUBS 0.008189f
C596 B.n335 VSUBS 0.008189f
C597 B.n336 VSUBS 0.008189f
C598 B.n337 VSUBS 0.008189f
C599 B.n338 VSUBS 0.008189f
C600 B.n339 VSUBS 0.008189f
C601 B.n340 VSUBS 0.008189f
C602 B.n341 VSUBS 0.008189f
C603 B.n342 VSUBS 0.008189f
C604 B.n343 VSUBS 0.008189f
C605 B.n344 VSUBS 0.008189f
C606 B.n345 VSUBS 0.008189f
C607 B.n346 VSUBS 0.008189f
C608 B.n347 VSUBS 0.008189f
C609 B.n348 VSUBS 0.008189f
C610 B.n349 VSUBS 0.008189f
C611 B.n350 VSUBS 0.008189f
C612 B.n351 VSUBS 0.008189f
C613 B.n352 VSUBS 0.008189f
C614 B.n353 VSUBS 0.008189f
C615 B.n354 VSUBS 0.008189f
C616 B.n355 VSUBS 0.008189f
C617 B.n356 VSUBS 0.008189f
C618 B.n357 VSUBS 0.008189f
C619 B.n358 VSUBS 0.008189f
C620 B.n359 VSUBS 0.008189f
C621 B.n360 VSUBS 0.008189f
C622 B.n361 VSUBS 0.008189f
C623 B.n362 VSUBS 0.008189f
C624 B.n363 VSUBS 0.008189f
C625 B.n364 VSUBS 0.008189f
C626 B.n365 VSUBS 0.008189f
C627 B.n366 VSUBS 0.008189f
C628 B.n367 VSUBS 0.008189f
C629 B.n368 VSUBS 0.008189f
C630 B.n369 VSUBS 0.008189f
C631 B.n370 VSUBS 0.008189f
C632 B.n371 VSUBS 0.008189f
C633 B.n372 VSUBS 0.018665f
C634 B.n373 VSUBS 0.018665f
C635 B.n374 VSUBS 0.019633f
C636 B.n375 VSUBS 0.008189f
C637 B.n376 VSUBS 0.008189f
C638 B.n377 VSUBS 0.008189f
C639 B.n378 VSUBS 0.008189f
C640 B.n379 VSUBS 0.008189f
C641 B.n380 VSUBS 0.008189f
C642 B.n381 VSUBS 0.008189f
C643 B.n382 VSUBS 0.008189f
C644 B.n383 VSUBS 0.008189f
C645 B.n384 VSUBS 0.008189f
C646 B.n385 VSUBS 0.008189f
C647 B.n386 VSUBS 0.008189f
C648 B.n387 VSUBS 0.008189f
C649 B.n388 VSUBS 0.008189f
C650 B.n389 VSUBS 0.008189f
C651 B.n390 VSUBS 0.008189f
C652 B.n391 VSUBS 0.008189f
C653 B.n392 VSUBS 0.008189f
C654 B.n393 VSUBS 0.00566f
C655 B.n394 VSUBS 0.008189f
C656 B.n395 VSUBS 0.008189f
C657 B.n396 VSUBS 0.006624f
C658 B.n397 VSUBS 0.008189f
C659 B.n398 VSUBS 0.008189f
C660 B.n399 VSUBS 0.008189f
C661 B.n400 VSUBS 0.008189f
C662 B.n401 VSUBS 0.008189f
C663 B.n402 VSUBS 0.008189f
C664 B.n403 VSUBS 0.008189f
C665 B.n404 VSUBS 0.008189f
C666 B.n405 VSUBS 0.008189f
C667 B.n406 VSUBS 0.008189f
C668 B.n407 VSUBS 0.008189f
C669 B.n408 VSUBS 0.006624f
C670 B.n409 VSUBS 0.018974f
C671 B.n410 VSUBS 0.00566f
C672 B.n411 VSUBS 0.008189f
C673 B.n412 VSUBS 0.008189f
C674 B.n413 VSUBS 0.008189f
C675 B.n414 VSUBS 0.008189f
C676 B.n415 VSUBS 0.008189f
C677 B.n416 VSUBS 0.008189f
C678 B.n417 VSUBS 0.008189f
C679 B.n418 VSUBS 0.008189f
C680 B.n419 VSUBS 0.008189f
C681 B.n420 VSUBS 0.008189f
C682 B.n421 VSUBS 0.008189f
C683 B.n422 VSUBS 0.008189f
C684 B.n423 VSUBS 0.008189f
C685 B.n424 VSUBS 0.008189f
C686 B.n425 VSUBS 0.008189f
C687 B.n426 VSUBS 0.008189f
C688 B.n427 VSUBS 0.008189f
C689 B.n428 VSUBS 0.008189f
C690 B.n429 VSUBS 0.019633f
C691 B.n430 VSUBS 0.019633f
C692 B.n431 VSUBS 0.018665f
C693 B.n432 VSUBS 0.008189f
C694 B.n433 VSUBS 0.008189f
C695 B.n434 VSUBS 0.008189f
C696 B.n435 VSUBS 0.008189f
C697 B.n436 VSUBS 0.008189f
C698 B.n437 VSUBS 0.008189f
C699 B.n438 VSUBS 0.008189f
C700 B.n439 VSUBS 0.008189f
C701 B.n440 VSUBS 0.008189f
C702 B.n441 VSUBS 0.008189f
C703 B.n442 VSUBS 0.008189f
C704 B.n443 VSUBS 0.008189f
C705 B.n444 VSUBS 0.008189f
C706 B.n445 VSUBS 0.008189f
C707 B.n446 VSUBS 0.008189f
C708 B.n447 VSUBS 0.008189f
C709 B.n448 VSUBS 0.008189f
C710 B.n449 VSUBS 0.008189f
C711 B.n450 VSUBS 0.008189f
C712 B.n451 VSUBS 0.008189f
C713 B.n452 VSUBS 0.008189f
C714 B.n453 VSUBS 0.008189f
C715 B.n454 VSUBS 0.008189f
C716 B.n455 VSUBS 0.008189f
C717 B.n456 VSUBS 0.008189f
C718 B.n457 VSUBS 0.008189f
C719 B.n458 VSUBS 0.008189f
C720 B.n459 VSUBS 0.008189f
C721 B.n460 VSUBS 0.008189f
C722 B.n461 VSUBS 0.008189f
C723 B.n462 VSUBS 0.008189f
C724 B.n463 VSUBS 0.008189f
C725 B.n464 VSUBS 0.008189f
C726 B.n465 VSUBS 0.008189f
C727 B.n466 VSUBS 0.008189f
C728 B.n467 VSUBS 0.008189f
C729 B.n468 VSUBS 0.008189f
C730 B.n469 VSUBS 0.008189f
C731 B.n470 VSUBS 0.008189f
C732 B.n471 VSUBS 0.008189f
C733 B.n472 VSUBS 0.008189f
C734 B.n473 VSUBS 0.008189f
C735 B.n474 VSUBS 0.008189f
C736 B.n475 VSUBS 0.008189f
C737 B.n476 VSUBS 0.008189f
C738 B.n477 VSUBS 0.008189f
C739 B.n478 VSUBS 0.008189f
C740 B.n479 VSUBS 0.008189f
C741 B.n480 VSUBS 0.008189f
C742 B.n481 VSUBS 0.008189f
C743 B.n482 VSUBS 0.008189f
C744 B.n483 VSUBS 0.008189f
C745 B.n484 VSUBS 0.008189f
C746 B.n485 VSUBS 0.008189f
C747 B.n486 VSUBS 0.008189f
C748 B.n487 VSUBS 0.008189f
C749 B.n488 VSUBS 0.008189f
C750 B.n489 VSUBS 0.008189f
C751 B.n490 VSUBS 0.008189f
C752 B.n491 VSUBS 0.010687f
C753 B.n492 VSUBS 0.011384f
C754 B.n493 VSUBS 0.022639f
.ends

