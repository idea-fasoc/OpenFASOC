* NGSPICE file created from diff_pair_sample_1723.ext - technology: sky130A

.subckt diff_pair_sample_1723 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t16 w_n2662_n4736# sky130_fd_pr__pfet_01v8 ad=3.1086 pd=19.17 as=7.3476 ps=38.46 w=18.84 l=1.08
X1 VTAIL.t7 VN.t0 VDD2.t9 w_n2662_n4736# sky130_fd_pr__pfet_01v8 ad=3.1086 pd=19.17 as=3.1086 ps=19.17 w=18.84 l=1.08
X2 VDD2.t8 VN.t1 VTAIL.t9 w_n2662_n4736# sky130_fd_pr__pfet_01v8 ad=7.3476 pd=38.46 as=3.1086 ps=19.17 w=18.84 l=1.08
X3 B.t11 B.t9 B.t10 w_n2662_n4736# sky130_fd_pr__pfet_01v8 ad=7.3476 pd=38.46 as=0 ps=0 w=18.84 l=1.08
X4 VTAIL.t11 VP.t1 VDD1.t8 w_n2662_n4736# sky130_fd_pr__pfet_01v8 ad=3.1086 pd=19.17 as=3.1086 ps=19.17 w=18.84 l=1.08
X5 VTAIL.t19 VP.t2 VDD1.t7 w_n2662_n4736# sky130_fd_pr__pfet_01v8 ad=3.1086 pd=19.17 as=3.1086 ps=19.17 w=18.84 l=1.08
X6 VTAIL.t10 VP.t3 VDD1.t6 w_n2662_n4736# sky130_fd_pr__pfet_01v8 ad=3.1086 pd=19.17 as=3.1086 ps=19.17 w=18.84 l=1.08
X7 VTAIL.t0 VN.t2 VDD2.t7 w_n2662_n4736# sky130_fd_pr__pfet_01v8 ad=3.1086 pd=19.17 as=3.1086 ps=19.17 w=18.84 l=1.08
X8 VDD1.t5 VP.t4 VTAIL.t15 w_n2662_n4736# sky130_fd_pr__pfet_01v8 ad=7.3476 pd=38.46 as=3.1086 ps=19.17 w=18.84 l=1.08
X9 VDD2.t6 VN.t3 VTAIL.t8 w_n2662_n4736# sky130_fd_pr__pfet_01v8 ad=3.1086 pd=19.17 as=3.1086 ps=19.17 w=18.84 l=1.08
X10 VTAIL.t1 VN.t4 VDD2.t5 w_n2662_n4736# sky130_fd_pr__pfet_01v8 ad=3.1086 pd=19.17 as=3.1086 ps=19.17 w=18.84 l=1.08
X11 VDD2.t4 VN.t5 VTAIL.t5 w_n2662_n4736# sky130_fd_pr__pfet_01v8 ad=3.1086 pd=19.17 as=7.3476 ps=38.46 w=18.84 l=1.08
X12 VTAIL.t2 VN.t6 VDD2.t3 w_n2662_n4736# sky130_fd_pr__pfet_01v8 ad=3.1086 pd=19.17 as=3.1086 ps=19.17 w=18.84 l=1.08
X13 VDD1.t4 VP.t5 VTAIL.t17 w_n2662_n4736# sky130_fd_pr__pfet_01v8 ad=3.1086 pd=19.17 as=3.1086 ps=19.17 w=18.84 l=1.08
X14 VTAIL.t13 VP.t6 VDD1.t3 w_n2662_n4736# sky130_fd_pr__pfet_01v8 ad=3.1086 pd=19.17 as=3.1086 ps=19.17 w=18.84 l=1.08
X15 B.t8 B.t6 B.t7 w_n2662_n4736# sky130_fd_pr__pfet_01v8 ad=7.3476 pd=38.46 as=0 ps=0 w=18.84 l=1.08
X16 VDD1.t2 VP.t7 VTAIL.t18 w_n2662_n4736# sky130_fd_pr__pfet_01v8 ad=7.3476 pd=38.46 as=3.1086 ps=19.17 w=18.84 l=1.08
X17 B.t5 B.t3 B.t4 w_n2662_n4736# sky130_fd_pr__pfet_01v8 ad=7.3476 pd=38.46 as=0 ps=0 w=18.84 l=1.08
X18 VDD2.t2 VN.t7 VTAIL.t3 w_n2662_n4736# sky130_fd_pr__pfet_01v8 ad=3.1086 pd=19.17 as=7.3476 ps=38.46 w=18.84 l=1.08
X19 VDD1.t1 VP.t8 VTAIL.t14 w_n2662_n4736# sky130_fd_pr__pfet_01v8 ad=3.1086 pd=19.17 as=7.3476 ps=38.46 w=18.84 l=1.08
X20 VDD2.t1 VN.t8 VTAIL.t4 w_n2662_n4736# sky130_fd_pr__pfet_01v8 ad=3.1086 pd=19.17 as=3.1086 ps=19.17 w=18.84 l=1.08
X21 VDD2.t0 VN.t9 VTAIL.t6 w_n2662_n4736# sky130_fd_pr__pfet_01v8 ad=7.3476 pd=38.46 as=3.1086 ps=19.17 w=18.84 l=1.08
X22 VDD1.t0 VP.t9 VTAIL.t12 w_n2662_n4736# sky130_fd_pr__pfet_01v8 ad=3.1086 pd=19.17 as=3.1086 ps=19.17 w=18.84 l=1.08
X23 B.t2 B.t0 B.t1 w_n2662_n4736# sky130_fd_pr__pfet_01v8 ad=7.3476 pd=38.46 as=0 ps=0 w=18.84 l=1.08
R0 VP.n10 VP.t7 477.848
R1 VP.n5 VP.t4 456.784
R2 VP.n41 VP.t8 456.784
R3 VP.n23 VP.t0 456.784
R4 VP.n34 VP.t9 420.411
R5 VP.n29 VP.t1 420.411
R6 VP.n1 VP.t2 420.411
R7 VP.n16 VP.t5 420.411
R8 VP.n7 VP.t3 420.411
R9 VP.n11 VP.t6 420.411
R10 VP.n13 VP.n12 161.3
R11 VP.n14 VP.n9 161.3
R12 VP.n16 VP.n15 161.3
R13 VP.n17 VP.n8 161.3
R14 VP.n19 VP.n18 161.3
R15 VP.n21 VP.n20 161.3
R16 VP.n22 VP.n6 161.3
R17 VP.n40 VP.n0 161.3
R18 VP.n39 VP.n38 161.3
R19 VP.n37 VP.n36 161.3
R20 VP.n35 VP.n2 161.3
R21 VP.n34 VP.n33 161.3
R22 VP.n32 VP.n3 161.3
R23 VP.n31 VP.n30 161.3
R24 VP.n28 VP.n4 161.3
R25 VP.n27 VP.n26 161.3
R26 VP.n24 VP.n23 80.6037
R27 VP.n42 VP.n41 80.6037
R28 VP.n25 VP.n5 80.6037
R29 VP.n30 VP.n3 56.5617
R30 VP.n36 VP.n35 56.5617
R31 VP.n18 VP.n17 56.5617
R32 VP.n12 VP.n9 56.5617
R33 VP.n25 VP.n24 50.134
R34 VP.n27 VP.n5 40.8975
R35 VP.n41 VP.n40 40.8975
R36 VP.n23 VP.n22 40.8975
R37 VP.n11 VP.n10 37.106
R38 VP.n28 VP.n27 29.4362
R39 VP.n40 VP.n39 29.4362
R40 VP.n22 VP.n21 29.4362
R41 VP.n13 VP.n10 28.8662
R42 VP.n34 VP.n3 24.5923
R43 VP.n35 VP.n34 24.5923
R44 VP.n16 VP.n9 24.5923
R45 VP.n17 VP.n16 24.5923
R46 VP.n30 VP.n29 20.1658
R47 VP.n36 VP.n1 20.1658
R48 VP.n18 VP.n7 20.1658
R49 VP.n12 VP.n11 20.1658
R50 VP.n29 VP.n28 4.42703
R51 VP.n39 VP.n1 4.42703
R52 VP.n21 VP.n7 4.42703
R53 VP.n24 VP.n6 0.285035
R54 VP.n26 VP.n25 0.285035
R55 VP.n42 VP.n0 0.285035
R56 VP.n14 VP.n13 0.189894
R57 VP.n15 VP.n14 0.189894
R58 VP.n15 VP.n8 0.189894
R59 VP.n19 VP.n8 0.189894
R60 VP.n20 VP.n19 0.189894
R61 VP.n20 VP.n6 0.189894
R62 VP.n26 VP.n4 0.189894
R63 VP.n31 VP.n4 0.189894
R64 VP.n32 VP.n31 0.189894
R65 VP.n33 VP.n32 0.189894
R66 VP.n33 VP.n2 0.189894
R67 VP.n37 VP.n2 0.189894
R68 VP.n38 VP.n37 0.189894
R69 VP.n38 VP.n0 0.189894
R70 VP VP.n42 0.146778
R71 VTAIL.n432 VTAIL.n332 756.745
R72 VTAIL.n102 VTAIL.n2 756.745
R73 VTAIL.n326 VTAIL.n226 756.745
R74 VTAIL.n216 VTAIL.n116 756.745
R75 VTAIL.n367 VTAIL.n366 585
R76 VTAIL.n364 VTAIL.n363 585
R77 VTAIL.n373 VTAIL.n372 585
R78 VTAIL.n375 VTAIL.n374 585
R79 VTAIL.n360 VTAIL.n359 585
R80 VTAIL.n381 VTAIL.n380 585
R81 VTAIL.n383 VTAIL.n382 585
R82 VTAIL.n356 VTAIL.n355 585
R83 VTAIL.n389 VTAIL.n388 585
R84 VTAIL.n391 VTAIL.n390 585
R85 VTAIL.n352 VTAIL.n351 585
R86 VTAIL.n397 VTAIL.n396 585
R87 VTAIL.n399 VTAIL.n398 585
R88 VTAIL.n348 VTAIL.n347 585
R89 VTAIL.n405 VTAIL.n404 585
R90 VTAIL.n408 VTAIL.n407 585
R91 VTAIL.n406 VTAIL.n344 585
R92 VTAIL.n413 VTAIL.n343 585
R93 VTAIL.n415 VTAIL.n414 585
R94 VTAIL.n417 VTAIL.n416 585
R95 VTAIL.n340 VTAIL.n339 585
R96 VTAIL.n423 VTAIL.n422 585
R97 VTAIL.n425 VTAIL.n424 585
R98 VTAIL.n336 VTAIL.n335 585
R99 VTAIL.n431 VTAIL.n430 585
R100 VTAIL.n433 VTAIL.n432 585
R101 VTAIL.n37 VTAIL.n36 585
R102 VTAIL.n34 VTAIL.n33 585
R103 VTAIL.n43 VTAIL.n42 585
R104 VTAIL.n45 VTAIL.n44 585
R105 VTAIL.n30 VTAIL.n29 585
R106 VTAIL.n51 VTAIL.n50 585
R107 VTAIL.n53 VTAIL.n52 585
R108 VTAIL.n26 VTAIL.n25 585
R109 VTAIL.n59 VTAIL.n58 585
R110 VTAIL.n61 VTAIL.n60 585
R111 VTAIL.n22 VTAIL.n21 585
R112 VTAIL.n67 VTAIL.n66 585
R113 VTAIL.n69 VTAIL.n68 585
R114 VTAIL.n18 VTAIL.n17 585
R115 VTAIL.n75 VTAIL.n74 585
R116 VTAIL.n78 VTAIL.n77 585
R117 VTAIL.n76 VTAIL.n14 585
R118 VTAIL.n83 VTAIL.n13 585
R119 VTAIL.n85 VTAIL.n84 585
R120 VTAIL.n87 VTAIL.n86 585
R121 VTAIL.n10 VTAIL.n9 585
R122 VTAIL.n93 VTAIL.n92 585
R123 VTAIL.n95 VTAIL.n94 585
R124 VTAIL.n6 VTAIL.n5 585
R125 VTAIL.n101 VTAIL.n100 585
R126 VTAIL.n103 VTAIL.n102 585
R127 VTAIL.n327 VTAIL.n326 585
R128 VTAIL.n325 VTAIL.n324 585
R129 VTAIL.n230 VTAIL.n229 585
R130 VTAIL.n319 VTAIL.n318 585
R131 VTAIL.n317 VTAIL.n316 585
R132 VTAIL.n234 VTAIL.n233 585
R133 VTAIL.n311 VTAIL.n310 585
R134 VTAIL.n309 VTAIL.n308 585
R135 VTAIL.n307 VTAIL.n237 585
R136 VTAIL.n241 VTAIL.n238 585
R137 VTAIL.n302 VTAIL.n301 585
R138 VTAIL.n300 VTAIL.n299 585
R139 VTAIL.n243 VTAIL.n242 585
R140 VTAIL.n294 VTAIL.n293 585
R141 VTAIL.n292 VTAIL.n291 585
R142 VTAIL.n247 VTAIL.n246 585
R143 VTAIL.n286 VTAIL.n285 585
R144 VTAIL.n284 VTAIL.n283 585
R145 VTAIL.n251 VTAIL.n250 585
R146 VTAIL.n278 VTAIL.n277 585
R147 VTAIL.n276 VTAIL.n275 585
R148 VTAIL.n255 VTAIL.n254 585
R149 VTAIL.n270 VTAIL.n269 585
R150 VTAIL.n268 VTAIL.n267 585
R151 VTAIL.n259 VTAIL.n258 585
R152 VTAIL.n262 VTAIL.n261 585
R153 VTAIL.n217 VTAIL.n216 585
R154 VTAIL.n215 VTAIL.n214 585
R155 VTAIL.n120 VTAIL.n119 585
R156 VTAIL.n209 VTAIL.n208 585
R157 VTAIL.n207 VTAIL.n206 585
R158 VTAIL.n124 VTAIL.n123 585
R159 VTAIL.n201 VTAIL.n200 585
R160 VTAIL.n199 VTAIL.n198 585
R161 VTAIL.n197 VTAIL.n127 585
R162 VTAIL.n131 VTAIL.n128 585
R163 VTAIL.n192 VTAIL.n191 585
R164 VTAIL.n190 VTAIL.n189 585
R165 VTAIL.n133 VTAIL.n132 585
R166 VTAIL.n184 VTAIL.n183 585
R167 VTAIL.n182 VTAIL.n181 585
R168 VTAIL.n137 VTAIL.n136 585
R169 VTAIL.n176 VTAIL.n175 585
R170 VTAIL.n174 VTAIL.n173 585
R171 VTAIL.n141 VTAIL.n140 585
R172 VTAIL.n168 VTAIL.n167 585
R173 VTAIL.n166 VTAIL.n165 585
R174 VTAIL.n145 VTAIL.n144 585
R175 VTAIL.n160 VTAIL.n159 585
R176 VTAIL.n158 VTAIL.n157 585
R177 VTAIL.n149 VTAIL.n148 585
R178 VTAIL.n152 VTAIL.n151 585
R179 VTAIL.t16 VTAIL.n260 327.466
R180 VTAIL.t5 VTAIL.n150 327.466
R181 VTAIL.t3 VTAIL.n365 327.466
R182 VTAIL.t14 VTAIL.n35 327.466
R183 VTAIL.n366 VTAIL.n363 171.744
R184 VTAIL.n373 VTAIL.n363 171.744
R185 VTAIL.n374 VTAIL.n373 171.744
R186 VTAIL.n374 VTAIL.n359 171.744
R187 VTAIL.n381 VTAIL.n359 171.744
R188 VTAIL.n382 VTAIL.n381 171.744
R189 VTAIL.n382 VTAIL.n355 171.744
R190 VTAIL.n389 VTAIL.n355 171.744
R191 VTAIL.n390 VTAIL.n389 171.744
R192 VTAIL.n390 VTAIL.n351 171.744
R193 VTAIL.n397 VTAIL.n351 171.744
R194 VTAIL.n398 VTAIL.n397 171.744
R195 VTAIL.n398 VTAIL.n347 171.744
R196 VTAIL.n405 VTAIL.n347 171.744
R197 VTAIL.n407 VTAIL.n405 171.744
R198 VTAIL.n407 VTAIL.n406 171.744
R199 VTAIL.n406 VTAIL.n343 171.744
R200 VTAIL.n415 VTAIL.n343 171.744
R201 VTAIL.n416 VTAIL.n415 171.744
R202 VTAIL.n416 VTAIL.n339 171.744
R203 VTAIL.n423 VTAIL.n339 171.744
R204 VTAIL.n424 VTAIL.n423 171.744
R205 VTAIL.n424 VTAIL.n335 171.744
R206 VTAIL.n431 VTAIL.n335 171.744
R207 VTAIL.n432 VTAIL.n431 171.744
R208 VTAIL.n36 VTAIL.n33 171.744
R209 VTAIL.n43 VTAIL.n33 171.744
R210 VTAIL.n44 VTAIL.n43 171.744
R211 VTAIL.n44 VTAIL.n29 171.744
R212 VTAIL.n51 VTAIL.n29 171.744
R213 VTAIL.n52 VTAIL.n51 171.744
R214 VTAIL.n52 VTAIL.n25 171.744
R215 VTAIL.n59 VTAIL.n25 171.744
R216 VTAIL.n60 VTAIL.n59 171.744
R217 VTAIL.n60 VTAIL.n21 171.744
R218 VTAIL.n67 VTAIL.n21 171.744
R219 VTAIL.n68 VTAIL.n67 171.744
R220 VTAIL.n68 VTAIL.n17 171.744
R221 VTAIL.n75 VTAIL.n17 171.744
R222 VTAIL.n77 VTAIL.n75 171.744
R223 VTAIL.n77 VTAIL.n76 171.744
R224 VTAIL.n76 VTAIL.n13 171.744
R225 VTAIL.n85 VTAIL.n13 171.744
R226 VTAIL.n86 VTAIL.n85 171.744
R227 VTAIL.n86 VTAIL.n9 171.744
R228 VTAIL.n93 VTAIL.n9 171.744
R229 VTAIL.n94 VTAIL.n93 171.744
R230 VTAIL.n94 VTAIL.n5 171.744
R231 VTAIL.n101 VTAIL.n5 171.744
R232 VTAIL.n102 VTAIL.n101 171.744
R233 VTAIL.n326 VTAIL.n325 171.744
R234 VTAIL.n325 VTAIL.n229 171.744
R235 VTAIL.n318 VTAIL.n229 171.744
R236 VTAIL.n318 VTAIL.n317 171.744
R237 VTAIL.n317 VTAIL.n233 171.744
R238 VTAIL.n310 VTAIL.n233 171.744
R239 VTAIL.n310 VTAIL.n309 171.744
R240 VTAIL.n309 VTAIL.n237 171.744
R241 VTAIL.n241 VTAIL.n237 171.744
R242 VTAIL.n301 VTAIL.n241 171.744
R243 VTAIL.n301 VTAIL.n300 171.744
R244 VTAIL.n300 VTAIL.n242 171.744
R245 VTAIL.n293 VTAIL.n242 171.744
R246 VTAIL.n293 VTAIL.n292 171.744
R247 VTAIL.n292 VTAIL.n246 171.744
R248 VTAIL.n285 VTAIL.n246 171.744
R249 VTAIL.n285 VTAIL.n284 171.744
R250 VTAIL.n284 VTAIL.n250 171.744
R251 VTAIL.n277 VTAIL.n250 171.744
R252 VTAIL.n277 VTAIL.n276 171.744
R253 VTAIL.n276 VTAIL.n254 171.744
R254 VTAIL.n269 VTAIL.n254 171.744
R255 VTAIL.n269 VTAIL.n268 171.744
R256 VTAIL.n268 VTAIL.n258 171.744
R257 VTAIL.n261 VTAIL.n258 171.744
R258 VTAIL.n216 VTAIL.n215 171.744
R259 VTAIL.n215 VTAIL.n119 171.744
R260 VTAIL.n208 VTAIL.n119 171.744
R261 VTAIL.n208 VTAIL.n207 171.744
R262 VTAIL.n207 VTAIL.n123 171.744
R263 VTAIL.n200 VTAIL.n123 171.744
R264 VTAIL.n200 VTAIL.n199 171.744
R265 VTAIL.n199 VTAIL.n127 171.744
R266 VTAIL.n131 VTAIL.n127 171.744
R267 VTAIL.n191 VTAIL.n131 171.744
R268 VTAIL.n191 VTAIL.n190 171.744
R269 VTAIL.n190 VTAIL.n132 171.744
R270 VTAIL.n183 VTAIL.n132 171.744
R271 VTAIL.n183 VTAIL.n182 171.744
R272 VTAIL.n182 VTAIL.n136 171.744
R273 VTAIL.n175 VTAIL.n136 171.744
R274 VTAIL.n175 VTAIL.n174 171.744
R275 VTAIL.n174 VTAIL.n140 171.744
R276 VTAIL.n167 VTAIL.n140 171.744
R277 VTAIL.n167 VTAIL.n166 171.744
R278 VTAIL.n166 VTAIL.n144 171.744
R279 VTAIL.n159 VTAIL.n144 171.744
R280 VTAIL.n159 VTAIL.n158 171.744
R281 VTAIL.n158 VTAIL.n148 171.744
R282 VTAIL.n151 VTAIL.n148 171.744
R283 VTAIL.n366 VTAIL.t3 85.8723
R284 VTAIL.n36 VTAIL.t14 85.8723
R285 VTAIL.n261 VTAIL.t16 85.8723
R286 VTAIL.n151 VTAIL.t5 85.8723
R287 VTAIL.n439 VTAIL.n438 49.3789
R288 VTAIL.n1 VTAIL.n0 49.3789
R289 VTAIL.n109 VTAIL.n108 49.3789
R290 VTAIL.n111 VTAIL.n110 49.3789
R291 VTAIL.n225 VTAIL.n224 49.3789
R292 VTAIL.n223 VTAIL.n222 49.3789
R293 VTAIL.n115 VTAIL.n114 49.3789
R294 VTAIL.n113 VTAIL.n112 49.3789
R295 VTAIL.n113 VTAIL.n111 31.0393
R296 VTAIL.n437 VTAIL.n436 29.8581
R297 VTAIL.n107 VTAIL.n106 29.8581
R298 VTAIL.n331 VTAIL.n330 29.8581
R299 VTAIL.n221 VTAIL.n220 29.8581
R300 VTAIL.n437 VTAIL.n331 29.8238
R301 VTAIL.n367 VTAIL.n365 16.3895
R302 VTAIL.n37 VTAIL.n35 16.3895
R303 VTAIL.n262 VTAIL.n260 16.3895
R304 VTAIL.n152 VTAIL.n150 16.3895
R305 VTAIL.n414 VTAIL.n413 13.1884
R306 VTAIL.n84 VTAIL.n83 13.1884
R307 VTAIL.n308 VTAIL.n307 13.1884
R308 VTAIL.n198 VTAIL.n197 13.1884
R309 VTAIL.n368 VTAIL.n364 12.8005
R310 VTAIL.n412 VTAIL.n344 12.8005
R311 VTAIL.n417 VTAIL.n342 12.8005
R312 VTAIL.n38 VTAIL.n34 12.8005
R313 VTAIL.n82 VTAIL.n14 12.8005
R314 VTAIL.n87 VTAIL.n12 12.8005
R315 VTAIL.n311 VTAIL.n236 12.8005
R316 VTAIL.n306 VTAIL.n238 12.8005
R317 VTAIL.n263 VTAIL.n259 12.8005
R318 VTAIL.n201 VTAIL.n126 12.8005
R319 VTAIL.n196 VTAIL.n128 12.8005
R320 VTAIL.n153 VTAIL.n149 12.8005
R321 VTAIL.n372 VTAIL.n371 12.0247
R322 VTAIL.n409 VTAIL.n408 12.0247
R323 VTAIL.n418 VTAIL.n340 12.0247
R324 VTAIL.n42 VTAIL.n41 12.0247
R325 VTAIL.n79 VTAIL.n78 12.0247
R326 VTAIL.n88 VTAIL.n10 12.0247
R327 VTAIL.n312 VTAIL.n234 12.0247
R328 VTAIL.n303 VTAIL.n302 12.0247
R329 VTAIL.n267 VTAIL.n266 12.0247
R330 VTAIL.n202 VTAIL.n124 12.0247
R331 VTAIL.n193 VTAIL.n192 12.0247
R332 VTAIL.n157 VTAIL.n156 12.0247
R333 VTAIL.n375 VTAIL.n362 11.249
R334 VTAIL.n404 VTAIL.n346 11.249
R335 VTAIL.n422 VTAIL.n421 11.249
R336 VTAIL.n45 VTAIL.n32 11.249
R337 VTAIL.n74 VTAIL.n16 11.249
R338 VTAIL.n92 VTAIL.n91 11.249
R339 VTAIL.n316 VTAIL.n315 11.249
R340 VTAIL.n299 VTAIL.n240 11.249
R341 VTAIL.n270 VTAIL.n257 11.249
R342 VTAIL.n206 VTAIL.n205 11.249
R343 VTAIL.n189 VTAIL.n130 11.249
R344 VTAIL.n160 VTAIL.n147 11.249
R345 VTAIL.n376 VTAIL.n360 10.4732
R346 VTAIL.n403 VTAIL.n348 10.4732
R347 VTAIL.n425 VTAIL.n338 10.4732
R348 VTAIL.n46 VTAIL.n30 10.4732
R349 VTAIL.n73 VTAIL.n18 10.4732
R350 VTAIL.n95 VTAIL.n8 10.4732
R351 VTAIL.n319 VTAIL.n232 10.4732
R352 VTAIL.n298 VTAIL.n243 10.4732
R353 VTAIL.n271 VTAIL.n255 10.4732
R354 VTAIL.n209 VTAIL.n122 10.4732
R355 VTAIL.n188 VTAIL.n133 10.4732
R356 VTAIL.n161 VTAIL.n145 10.4732
R357 VTAIL.n380 VTAIL.n379 9.69747
R358 VTAIL.n400 VTAIL.n399 9.69747
R359 VTAIL.n426 VTAIL.n336 9.69747
R360 VTAIL.n50 VTAIL.n49 9.69747
R361 VTAIL.n70 VTAIL.n69 9.69747
R362 VTAIL.n96 VTAIL.n6 9.69747
R363 VTAIL.n320 VTAIL.n230 9.69747
R364 VTAIL.n295 VTAIL.n294 9.69747
R365 VTAIL.n275 VTAIL.n274 9.69747
R366 VTAIL.n210 VTAIL.n120 9.69747
R367 VTAIL.n185 VTAIL.n184 9.69747
R368 VTAIL.n165 VTAIL.n164 9.69747
R369 VTAIL.n436 VTAIL.n435 9.45567
R370 VTAIL.n106 VTAIL.n105 9.45567
R371 VTAIL.n330 VTAIL.n329 9.45567
R372 VTAIL.n220 VTAIL.n219 9.45567
R373 VTAIL.n334 VTAIL.n333 9.3005
R374 VTAIL.n429 VTAIL.n428 9.3005
R375 VTAIL.n427 VTAIL.n426 9.3005
R376 VTAIL.n338 VTAIL.n337 9.3005
R377 VTAIL.n421 VTAIL.n420 9.3005
R378 VTAIL.n419 VTAIL.n418 9.3005
R379 VTAIL.n342 VTAIL.n341 9.3005
R380 VTAIL.n387 VTAIL.n386 9.3005
R381 VTAIL.n385 VTAIL.n384 9.3005
R382 VTAIL.n358 VTAIL.n357 9.3005
R383 VTAIL.n379 VTAIL.n378 9.3005
R384 VTAIL.n377 VTAIL.n376 9.3005
R385 VTAIL.n362 VTAIL.n361 9.3005
R386 VTAIL.n371 VTAIL.n370 9.3005
R387 VTAIL.n369 VTAIL.n368 9.3005
R388 VTAIL.n354 VTAIL.n353 9.3005
R389 VTAIL.n393 VTAIL.n392 9.3005
R390 VTAIL.n395 VTAIL.n394 9.3005
R391 VTAIL.n350 VTAIL.n349 9.3005
R392 VTAIL.n401 VTAIL.n400 9.3005
R393 VTAIL.n403 VTAIL.n402 9.3005
R394 VTAIL.n346 VTAIL.n345 9.3005
R395 VTAIL.n410 VTAIL.n409 9.3005
R396 VTAIL.n412 VTAIL.n411 9.3005
R397 VTAIL.n435 VTAIL.n434 9.3005
R398 VTAIL.n4 VTAIL.n3 9.3005
R399 VTAIL.n99 VTAIL.n98 9.3005
R400 VTAIL.n97 VTAIL.n96 9.3005
R401 VTAIL.n8 VTAIL.n7 9.3005
R402 VTAIL.n91 VTAIL.n90 9.3005
R403 VTAIL.n89 VTAIL.n88 9.3005
R404 VTAIL.n12 VTAIL.n11 9.3005
R405 VTAIL.n57 VTAIL.n56 9.3005
R406 VTAIL.n55 VTAIL.n54 9.3005
R407 VTAIL.n28 VTAIL.n27 9.3005
R408 VTAIL.n49 VTAIL.n48 9.3005
R409 VTAIL.n47 VTAIL.n46 9.3005
R410 VTAIL.n32 VTAIL.n31 9.3005
R411 VTAIL.n41 VTAIL.n40 9.3005
R412 VTAIL.n39 VTAIL.n38 9.3005
R413 VTAIL.n24 VTAIL.n23 9.3005
R414 VTAIL.n63 VTAIL.n62 9.3005
R415 VTAIL.n65 VTAIL.n64 9.3005
R416 VTAIL.n20 VTAIL.n19 9.3005
R417 VTAIL.n71 VTAIL.n70 9.3005
R418 VTAIL.n73 VTAIL.n72 9.3005
R419 VTAIL.n16 VTAIL.n15 9.3005
R420 VTAIL.n80 VTAIL.n79 9.3005
R421 VTAIL.n82 VTAIL.n81 9.3005
R422 VTAIL.n105 VTAIL.n104 9.3005
R423 VTAIL.n288 VTAIL.n287 9.3005
R424 VTAIL.n290 VTAIL.n289 9.3005
R425 VTAIL.n245 VTAIL.n244 9.3005
R426 VTAIL.n296 VTAIL.n295 9.3005
R427 VTAIL.n298 VTAIL.n297 9.3005
R428 VTAIL.n240 VTAIL.n239 9.3005
R429 VTAIL.n304 VTAIL.n303 9.3005
R430 VTAIL.n306 VTAIL.n305 9.3005
R431 VTAIL.n329 VTAIL.n328 9.3005
R432 VTAIL.n228 VTAIL.n227 9.3005
R433 VTAIL.n323 VTAIL.n322 9.3005
R434 VTAIL.n321 VTAIL.n320 9.3005
R435 VTAIL.n232 VTAIL.n231 9.3005
R436 VTAIL.n315 VTAIL.n314 9.3005
R437 VTAIL.n313 VTAIL.n312 9.3005
R438 VTAIL.n236 VTAIL.n235 9.3005
R439 VTAIL.n249 VTAIL.n248 9.3005
R440 VTAIL.n282 VTAIL.n281 9.3005
R441 VTAIL.n280 VTAIL.n279 9.3005
R442 VTAIL.n253 VTAIL.n252 9.3005
R443 VTAIL.n274 VTAIL.n273 9.3005
R444 VTAIL.n272 VTAIL.n271 9.3005
R445 VTAIL.n257 VTAIL.n256 9.3005
R446 VTAIL.n266 VTAIL.n265 9.3005
R447 VTAIL.n264 VTAIL.n263 9.3005
R448 VTAIL.n178 VTAIL.n177 9.3005
R449 VTAIL.n180 VTAIL.n179 9.3005
R450 VTAIL.n135 VTAIL.n134 9.3005
R451 VTAIL.n186 VTAIL.n185 9.3005
R452 VTAIL.n188 VTAIL.n187 9.3005
R453 VTAIL.n130 VTAIL.n129 9.3005
R454 VTAIL.n194 VTAIL.n193 9.3005
R455 VTAIL.n196 VTAIL.n195 9.3005
R456 VTAIL.n219 VTAIL.n218 9.3005
R457 VTAIL.n118 VTAIL.n117 9.3005
R458 VTAIL.n213 VTAIL.n212 9.3005
R459 VTAIL.n211 VTAIL.n210 9.3005
R460 VTAIL.n122 VTAIL.n121 9.3005
R461 VTAIL.n205 VTAIL.n204 9.3005
R462 VTAIL.n203 VTAIL.n202 9.3005
R463 VTAIL.n126 VTAIL.n125 9.3005
R464 VTAIL.n139 VTAIL.n138 9.3005
R465 VTAIL.n172 VTAIL.n171 9.3005
R466 VTAIL.n170 VTAIL.n169 9.3005
R467 VTAIL.n143 VTAIL.n142 9.3005
R468 VTAIL.n164 VTAIL.n163 9.3005
R469 VTAIL.n162 VTAIL.n161 9.3005
R470 VTAIL.n147 VTAIL.n146 9.3005
R471 VTAIL.n156 VTAIL.n155 9.3005
R472 VTAIL.n154 VTAIL.n153 9.3005
R473 VTAIL.n383 VTAIL.n358 8.92171
R474 VTAIL.n396 VTAIL.n350 8.92171
R475 VTAIL.n430 VTAIL.n429 8.92171
R476 VTAIL.n53 VTAIL.n28 8.92171
R477 VTAIL.n66 VTAIL.n20 8.92171
R478 VTAIL.n100 VTAIL.n99 8.92171
R479 VTAIL.n324 VTAIL.n323 8.92171
R480 VTAIL.n291 VTAIL.n245 8.92171
R481 VTAIL.n278 VTAIL.n253 8.92171
R482 VTAIL.n214 VTAIL.n213 8.92171
R483 VTAIL.n181 VTAIL.n135 8.92171
R484 VTAIL.n168 VTAIL.n143 8.92171
R485 VTAIL.n384 VTAIL.n356 8.14595
R486 VTAIL.n395 VTAIL.n352 8.14595
R487 VTAIL.n433 VTAIL.n334 8.14595
R488 VTAIL.n54 VTAIL.n26 8.14595
R489 VTAIL.n65 VTAIL.n22 8.14595
R490 VTAIL.n103 VTAIL.n4 8.14595
R491 VTAIL.n327 VTAIL.n228 8.14595
R492 VTAIL.n290 VTAIL.n247 8.14595
R493 VTAIL.n279 VTAIL.n251 8.14595
R494 VTAIL.n217 VTAIL.n118 8.14595
R495 VTAIL.n180 VTAIL.n137 8.14595
R496 VTAIL.n169 VTAIL.n141 8.14595
R497 VTAIL.n388 VTAIL.n387 7.3702
R498 VTAIL.n392 VTAIL.n391 7.3702
R499 VTAIL.n434 VTAIL.n332 7.3702
R500 VTAIL.n58 VTAIL.n57 7.3702
R501 VTAIL.n62 VTAIL.n61 7.3702
R502 VTAIL.n104 VTAIL.n2 7.3702
R503 VTAIL.n328 VTAIL.n226 7.3702
R504 VTAIL.n287 VTAIL.n286 7.3702
R505 VTAIL.n283 VTAIL.n282 7.3702
R506 VTAIL.n218 VTAIL.n116 7.3702
R507 VTAIL.n177 VTAIL.n176 7.3702
R508 VTAIL.n173 VTAIL.n172 7.3702
R509 VTAIL.n388 VTAIL.n354 6.59444
R510 VTAIL.n391 VTAIL.n354 6.59444
R511 VTAIL.n436 VTAIL.n332 6.59444
R512 VTAIL.n58 VTAIL.n24 6.59444
R513 VTAIL.n61 VTAIL.n24 6.59444
R514 VTAIL.n106 VTAIL.n2 6.59444
R515 VTAIL.n330 VTAIL.n226 6.59444
R516 VTAIL.n286 VTAIL.n249 6.59444
R517 VTAIL.n283 VTAIL.n249 6.59444
R518 VTAIL.n220 VTAIL.n116 6.59444
R519 VTAIL.n176 VTAIL.n139 6.59444
R520 VTAIL.n173 VTAIL.n139 6.59444
R521 VTAIL.n387 VTAIL.n356 5.81868
R522 VTAIL.n392 VTAIL.n352 5.81868
R523 VTAIL.n434 VTAIL.n433 5.81868
R524 VTAIL.n57 VTAIL.n26 5.81868
R525 VTAIL.n62 VTAIL.n22 5.81868
R526 VTAIL.n104 VTAIL.n103 5.81868
R527 VTAIL.n328 VTAIL.n327 5.81868
R528 VTAIL.n287 VTAIL.n247 5.81868
R529 VTAIL.n282 VTAIL.n251 5.81868
R530 VTAIL.n218 VTAIL.n217 5.81868
R531 VTAIL.n177 VTAIL.n137 5.81868
R532 VTAIL.n172 VTAIL.n141 5.81868
R533 VTAIL.n384 VTAIL.n383 5.04292
R534 VTAIL.n396 VTAIL.n395 5.04292
R535 VTAIL.n430 VTAIL.n334 5.04292
R536 VTAIL.n54 VTAIL.n53 5.04292
R537 VTAIL.n66 VTAIL.n65 5.04292
R538 VTAIL.n100 VTAIL.n4 5.04292
R539 VTAIL.n324 VTAIL.n228 5.04292
R540 VTAIL.n291 VTAIL.n290 5.04292
R541 VTAIL.n279 VTAIL.n278 5.04292
R542 VTAIL.n214 VTAIL.n118 5.04292
R543 VTAIL.n181 VTAIL.n180 5.04292
R544 VTAIL.n169 VTAIL.n168 5.04292
R545 VTAIL.n380 VTAIL.n358 4.26717
R546 VTAIL.n399 VTAIL.n350 4.26717
R547 VTAIL.n429 VTAIL.n336 4.26717
R548 VTAIL.n50 VTAIL.n28 4.26717
R549 VTAIL.n69 VTAIL.n20 4.26717
R550 VTAIL.n99 VTAIL.n6 4.26717
R551 VTAIL.n323 VTAIL.n230 4.26717
R552 VTAIL.n294 VTAIL.n245 4.26717
R553 VTAIL.n275 VTAIL.n253 4.26717
R554 VTAIL.n213 VTAIL.n120 4.26717
R555 VTAIL.n184 VTAIL.n135 4.26717
R556 VTAIL.n165 VTAIL.n143 4.26717
R557 VTAIL.n369 VTAIL.n365 3.70982
R558 VTAIL.n39 VTAIL.n35 3.70982
R559 VTAIL.n264 VTAIL.n260 3.70982
R560 VTAIL.n154 VTAIL.n150 3.70982
R561 VTAIL.n379 VTAIL.n360 3.49141
R562 VTAIL.n400 VTAIL.n348 3.49141
R563 VTAIL.n426 VTAIL.n425 3.49141
R564 VTAIL.n49 VTAIL.n30 3.49141
R565 VTAIL.n70 VTAIL.n18 3.49141
R566 VTAIL.n96 VTAIL.n95 3.49141
R567 VTAIL.n320 VTAIL.n319 3.49141
R568 VTAIL.n295 VTAIL.n243 3.49141
R569 VTAIL.n274 VTAIL.n255 3.49141
R570 VTAIL.n210 VTAIL.n209 3.49141
R571 VTAIL.n185 VTAIL.n133 3.49141
R572 VTAIL.n164 VTAIL.n145 3.49141
R573 VTAIL.n376 VTAIL.n375 2.71565
R574 VTAIL.n404 VTAIL.n403 2.71565
R575 VTAIL.n422 VTAIL.n338 2.71565
R576 VTAIL.n46 VTAIL.n45 2.71565
R577 VTAIL.n74 VTAIL.n73 2.71565
R578 VTAIL.n92 VTAIL.n8 2.71565
R579 VTAIL.n316 VTAIL.n232 2.71565
R580 VTAIL.n299 VTAIL.n298 2.71565
R581 VTAIL.n271 VTAIL.n270 2.71565
R582 VTAIL.n206 VTAIL.n122 2.71565
R583 VTAIL.n189 VTAIL.n188 2.71565
R584 VTAIL.n161 VTAIL.n160 2.71565
R585 VTAIL.n372 VTAIL.n362 1.93989
R586 VTAIL.n408 VTAIL.n346 1.93989
R587 VTAIL.n421 VTAIL.n340 1.93989
R588 VTAIL.n42 VTAIL.n32 1.93989
R589 VTAIL.n78 VTAIL.n16 1.93989
R590 VTAIL.n91 VTAIL.n10 1.93989
R591 VTAIL.n315 VTAIL.n234 1.93989
R592 VTAIL.n302 VTAIL.n240 1.93989
R593 VTAIL.n267 VTAIL.n257 1.93989
R594 VTAIL.n205 VTAIL.n124 1.93989
R595 VTAIL.n192 VTAIL.n130 1.93989
R596 VTAIL.n157 VTAIL.n147 1.93989
R597 VTAIL.n438 VTAIL.t4 1.72582
R598 VTAIL.n438 VTAIL.t0 1.72582
R599 VTAIL.n0 VTAIL.t6 1.72582
R600 VTAIL.n0 VTAIL.t1 1.72582
R601 VTAIL.n108 VTAIL.t12 1.72582
R602 VTAIL.n108 VTAIL.t19 1.72582
R603 VTAIL.n110 VTAIL.t15 1.72582
R604 VTAIL.n110 VTAIL.t11 1.72582
R605 VTAIL.n224 VTAIL.t17 1.72582
R606 VTAIL.n224 VTAIL.t10 1.72582
R607 VTAIL.n222 VTAIL.t18 1.72582
R608 VTAIL.n222 VTAIL.t13 1.72582
R609 VTAIL.n114 VTAIL.t8 1.72582
R610 VTAIL.n114 VTAIL.t2 1.72582
R611 VTAIL.n112 VTAIL.t9 1.72582
R612 VTAIL.n112 VTAIL.t7 1.72582
R613 VTAIL.n115 VTAIL.n113 1.21602
R614 VTAIL.n221 VTAIL.n115 1.21602
R615 VTAIL.n225 VTAIL.n223 1.21602
R616 VTAIL.n331 VTAIL.n225 1.21602
R617 VTAIL.n111 VTAIL.n109 1.21602
R618 VTAIL.n109 VTAIL.n107 1.21602
R619 VTAIL.n439 VTAIL.n437 1.21602
R620 VTAIL.n371 VTAIL.n364 1.16414
R621 VTAIL.n409 VTAIL.n344 1.16414
R622 VTAIL.n418 VTAIL.n417 1.16414
R623 VTAIL.n41 VTAIL.n34 1.16414
R624 VTAIL.n79 VTAIL.n14 1.16414
R625 VTAIL.n88 VTAIL.n87 1.16414
R626 VTAIL.n312 VTAIL.n311 1.16414
R627 VTAIL.n303 VTAIL.n238 1.16414
R628 VTAIL.n266 VTAIL.n259 1.16414
R629 VTAIL.n202 VTAIL.n201 1.16414
R630 VTAIL.n193 VTAIL.n128 1.16414
R631 VTAIL.n156 VTAIL.n149 1.16414
R632 VTAIL.n223 VTAIL.n221 1.07809
R633 VTAIL.n107 VTAIL.n1 1.07809
R634 VTAIL VTAIL.n1 0.970328
R635 VTAIL.n368 VTAIL.n367 0.388379
R636 VTAIL.n413 VTAIL.n412 0.388379
R637 VTAIL.n414 VTAIL.n342 0.388379
R638 VTAIL.n38 VTAIL.n37 0.388379
R639 VTAIL.n83 VTAIL.n82 0.388379
R640 VTAIL.n84 VTAIL.n12 0.388379
R641 VTAIL.n308 VTAIL.n236 0.388379
R642 VTAIL.n307 VTAIL.n306 0.388379
R643 VTAIL.n263 VTAIL.n262 0.388379
R644 VTAIL.n198 VTAIL.n126 0.388379
R645 VTAIL.n197 VTAIL.n196 0.388379
R646 VTAIL.n153 VTAIL.n152 0.388379
R647 VTAIL VTAIL.n439 0.24619
R648 VTAIL.n370 VTAIL.n369 0.155672
R649 VTAIL.n370 VTAIL.n361 0.155672
R650 VTAIL.n377 VTAIL.n361 0.155672
R651 VTAIL.n378 VTAIL.n377 0.155672
R652 VTAIL.n378 VTAIL.n357 0.155672
R653 VTAIL.n385 VTAIL.n357 0.155672
R654 VTAIL.n386 VTAIL.n385 0.155672
R655 VTAIL.n386 VTAIL.n353 0.155672
R656 VTAIL.n393 VTAIL.n353 0.155672
R657 VTAIL.n394 VTAIL.n393 0.155672
R658 VTAIL.n394 VTAIL.n349 0.155672
R659 VTAIL.n401 VTAIL.n349 0.155672
R660 VTAIL.n402 VTAIL.n401 0.155672
R661 VTAIL.n402 VTAIL.n345 0.155672
R662 VTAIL.n410 VTAIL.n345 0.155672
R663 VTAIL.n411 VTAIL.n410 0.155672
R664 VTAIL.n411 VTAIL.n341 0.155672
R665 VTAIL.n419 VTAIL.n341 0.155672
R666 VTAIL.n420 VTAIL.n419 0.155672
R667 VTAIL.n420 VTAIL.n337 0.155672
R668 VTAIL.n427 VTAIL.n337 0.155672
R669 VTAIL.n428 VTAIL.n427 0.155672
R670 VTAIL.n428 VTAIL.n333 0.155672
R671 VTAIL.n435 VTAIL.n333 0.155672
R672 VTAIL.n40 VTAIL.n39 0.155672
R673 VTAIL.n40 VTAIL.n31 0.155672
R674 VTAIL.n47 VTAIL.n31 0.155672
R675 VTAIL.n48 VTAIL.n47 0.155672
R676 VTAIL.n48 VTAIL.n27 0.155672
R677 VTAIL.n55 VTAIL.n27 0.155672
R678 VTAIL.n56 VTAIL.n55 0.155672
R679 VTAIL.n56 VTAIL.n23 0.155672
R680 VTAIL.n63 VTAIL.n23 0.155672
R681 VTAIL.n64 VTAIL.n63 0.155672
R682 VTAIL.n64 VTAIL.n19 0.155672
R683 VTAIL.n71 VTAIL.n19 0.155672
R684 VTAIL.n72 VTAIL.n71 0.155672
R685 VTAIL.n72 VTAIL.n15 0.155672
R686 VTAIL.n80 VTAIL.n15 0.155672
R687 VTAIL.n81 VTAIL.n80 0.155672
R688 VTAIL.n81 VTAIL.n11 0.155672
R689 VTAIL.n89 VTAIL.n11 0.155672
R690 VTAIL.n90 VTAIL.n89 0.155672
R691 VTAIL.n90 VTAIL.n7 0.155672
R692 VTAIL.n97 VTAIL.n7 0.155672
R693 VTAIL.n98 VTAIL.n97 0.155672
R694 VTAIL.n98 VTAIL.n3 0.155672
R695 VTAIL.n105 VTAIL.n3 0.155672
R696 VTAIL.n329 VTAIL.n227 0.155672
R697 VTAIL.n322 VTAIL.n227 0.155672
R698 VTAIL.n322 VTAIL.n321 0.155672
R699 VTAIL.n321 VTAIL.n231 0.155672
R700 VTAIL.n314 VTAIL.n231 0.155672
R701 VTAIL.n314 VTAIL.n313 0.155672
R702 VTAIL.n313 VTAIL.n235 0.155672
R703 VTAIL.n305 VTAIL.n235 0.155672
R704 VTAIL.n305 VTAIL.n304 0.155672
R705 VTAIL.n304 VTAIL.n239 0.155672
R706 VTAIL.n297 VTAIL.n239 0.155672
R707 VTAIL.n297 VTAIL.n296 0.155672
R708 VTAIL.n296 VTAIL.n244 0.155672
R709 VTAIL.n289 VTAIL.n244 0.155672
R710 VTAIL.n289 VTAIL.n288 0.155672
R711 VTAIL.n288 VTAIL.n248 0.155672
R712 VTAIL.n281 VTAIL.n248 0.155672
R713 VTAIL.n281 VTAIL.n280 0.155672
R714 VTAIL.n280 VTAIL.n252 0.155672
R715 VTAIL.n273 VTAIL.n252 0.155672
R716 VTAIL.n273 VTAIL.n272 0.155672
R717 VTAIL.n272 VTAIL.n256 0.155672
R718 VTAIL.n265 VTAIL.n256 0.155672
R719 VTAIL.n265 VTAIL.n264 0.155672
R720 VTAIL.n219 VTAIL.n117 0.155672
R721 VTAIL.n212 VTAIL.n117 0.155672
R722 VTAIL.n212 VTAIL.n211 0.155672
R723 VTAIL.n211 VTAIL.n121 0.155672
R724 VTAIL.n204 VTAIL.n121 0.155672
R725 VTAIL.n204 VTAIL.n203 0.155672
R726 VTAIL.n203 VTAIL.n125 0.155672
R727 VTAIL.n195 VTAIL.n125 0.155672
R728 VTAIL.n195 VTAIL.n194 0.155672
R729 VTAIL.n194 VTAIL.n129 0.155672
R730 VTAIL.n187 VTAIL.n129 0.155672
R731 VTAIL.n187 VTAIL.n186 0.155672
R732 VTAIL.n186 VTAIL.n134 0.155672
R733 VTAIL.n179 VTAIL.n134 0.155672
R734 VTAIL.n179 VTAIL.n178 0.155672
R735 VTAIL.n178 VTAIL.n138 0.155672
R736 VTAIL.n171 VTAIL.n138 0.155672
R737 VTAIL.n171 VTAIL.n170 0.155672
R738 VTAIL.n170 VTAIL.n142 0.155672
R739 VTAIL.n163 VTAIL.n142 0.155672
R740 VTAIL.n163 VTAIL.n162 0.155672
R741 VTAIL.n162 VTAIL.n146 0.155672
R742 VTAIL.n155 VTAIL.n146 0.155672
R743 VTAIL.n155 VTAIL.n154 0.155672
R744 VDD1.n100 VDD1.n0 756.745
R745 VDD1.n207 VDD1.n107 756.745
R746 VDD1.n101 VDD1.n100 585
R747 VDD1.n99 VDD1.n98 585
R748 VDD1.n4 VDD1.n3 585
R749 VDD1.n93 VDD1.n92 585
R750 VDD1.n91 VDD1.n90 585
R751 VDD1.n8 VDD1.n7 585
R752 VDD1.n85 VDD1.n84 585
R753 VDD1.n83 VDD1.n82 585
R754 VDD1.n81 VDD1.n11 585
R755 VDD1.n15 VDD1.n12 585
R756 VDD1.n76 VDD1.n75 585
R757 VDD1.n74 VDD1.n73 585
R758 VDD1.n17 VDD1.n16 585
R759 VDD1.n68 VDD1.n67 585
R760 VDD1.n66 VDD1.n65 585
R761 VDD1.n21 VDD1.n20 585
R762 VDD1.n60 VDD1.n59 585
R763 VDD1.n58 VDD1.n57 585
R764 VDD1.n25 VDD1.n24 585
R765 VDD1.n52 VDD1.n51 585
R766 VDD1.n50 VDD1.n49 585
R767 VDD1.n29 VDD1.n28 585
R768 VDD1.n44 VDD1.n43 585
R769 VDD1.n42 VDD1.n41 585
R770 VDD1.n33 VDD1.n32 585
R771 VDD1.n36 VDD1.n35 585
R772 VDD1.n142 VDD1.n141 585
R773 VDD1.n139 VDD1.n138 585
R774 VDD1.n148 VDD1.n147 585
R775 VDD1.n150 VDD1.n149 585
R776 VDD1.n135 VDD1.n134 585
R777 VDD1.n156 VDD1.n155 585
R778 VDD1.n158 VDD1.n157 585
R779 VDD1.n131 VDD1.n130 585
R780 VDD1.n164 VDD1.n163 585
R781 VDD1.n166 VDD1.n165 585
R782 VDD1.n127 VDD1.n126 585
R783 VDD1.n172 VDD1.n171 585
R784 VDD1.n174 VDD1.n173 585
R785 VDD1.n123 VDD1.n122 585
R786 VDD1.n180 VDD1.n179 585
R787 VDD1.n183 VDD1.n182 585
R788 VDD1.n181 VDD1.n119 585
R789 VDD1.n188 VDD1.n118 585
R790 VDD1.n190 VDD1.n189 585
R791 VDD1.n192 VDD1.n191 585
R792 VDD1.n115 VDD1.n114 585
R793 VDD1.n198 VDD1.n197 585
R794 VDD1.n200 VDD1.n199 585
R795 VDD1.n111 VDD1.n110 585
R796 VDD1.n206 VDD1.n205 585
R797 VDD1.n208 VDD1.n207 585
R798 VDD1.t2 VDD1.n34 327.466
R799 VDD1.t5 VDD1.n140 327.466
R800 VDD1.n100 VDD1.n99 171.744
R801 VDD1.n99 VDD1.n3 171.744
R802 VDD1.n92 VDD1.n3 171.744
R803 VDD1.n92 VDD1.n91 171.744
R804 VDD1.n91 VDD1.n7 171.744
R805 VDD1.n84 VDD1.n7 171.744
R806 VDD1.n84 VDD1.n83 171.744
R807 VDD1.n83 VDD1.n11 171.744
R808 VDD1.n15 VDD1.n11 171.744
R809 VDD1.n75 VDD1.n15 171.744
R810 VDD1.n75 VDD1.n74 171.744
R811 VDD1.n74 VDD1.n16 171.744
R812 VDD1.n67 VDD1.n16 171.744
R813 VDD1.n67 VDD1.n66 171.744
R814 VDD1.n66 VDD1.n20 171.744
R815 VDD1.n59 VDD1.n20 171.744
R816 VDD1.n59 VDD1.n58 171.744
R817 VDD1.n58 VDD1.n24 171.744
R818 VDD1.n51 VDD1.n24 171.744
R819 VDD1.n51 VDD1.n50 171.744
R820 VDD1.n50 VDD1.n28 171.744
R821 VDD1.n43 VDD1.n28 171.744
R822 VDD1.n43 VDD1.n42 171.744
R823 VDD1.n42 VDD1.n32 171.744
R824 VDD1.n35 VDD1.n32 171.744
R825 VDD1.n141 VDD1.n138 171.744
R826 VDD1.n148 VDD1.n138 171.744
R827 VDD1.n149 VDD1.n148 171.744
R828 VDD1.n149 VDD1.n134 171.744
R829 VDD1.n156 VDD1.n134 171.744
R830 VDD1.n157 VDD1.n156 171.744
R831 VDD1.n157 VDD1.n130 171.744
R832 VDD1.n164 VDD1.n130 171.744
R833 VDD1.n165 VDD1.n164 171.744
R834 VDD1.n165 VDD1.n126 171.744
R835 VDD1.n172 VDD1.n126 171.744
R836 VDD1.n173 VDD1.n172 171.744
R837 VDD1.n173 VDD1.n122 171.744
R838 VDD1.n180 VDD1.n122 171.744
R839 VDD1.n182 VDD1.n180 171.744
R840 VDD1.n182 VDD1.n181 171.744
R841 VDD1.n181 VDD1.n118 171.744
R842 VDD1.n190 VDD1.n118 171.744
R843 VDD1.n191 VDD1.n190 171.744
R844 VDD1.n191 VDD1.n114 171.744
R845 VDD1.n198 VDD1.n114 171.744
R846 VDD1.n199 VDD1.n198 171.744
R847 VDD1.n199 VDD1.n110 171.744
R848 VDD1.n206 VDD1.n110 171.744
R849 VDD1.n207 VDD1.n206 171.744
R850 VDD1.n35 VDD1.t2 85.8723
R851 VDD1.n141 VDD1.t5 85.8723
R852 VDD1.n215 VDD1.n214 66.9139
R853 VDD1.n106 VDD1.n105 66.0577
R854 VDD1.n213 VDD1.n212 66.0577
R855 VDD1.n217 VDD1.n216 66.0575
R856 VDD1.n106 VDD1.n104 47.7524
R857 VDD1.n213 VDD1.n211 47.7524
R858 VDD1.n217 VDD1.n215 46.9212
R859 VDD1.n36 VDD1.n34 16.3895
R860 VDD1.n142 VDD1.n140 16.3895
R861 VDD1.n82 VDD1.n81 13.1884
R862 VDD1.n189 VDD1.n188 13.1884
R863 VDD1.n85 VDD1.n10 12.8005
R864 VDD1.n80 VDD1.n12 12.8005
R865 VDD1.n37 VDD1.n33 12.8005
R866 VDD1.n143 VDD1.n139 12.8005
R867 VDD1.n187 VDD1.n119 12.8005
R868 VDD1.n192 VDD1.n117 12.8005
R869 VDD1.n86 VDD1.n8 12.0247
R870 VDD1.n77 VDD1.n76 12.0247
R871 VDD1.n41 VDD1.n40 12.0247
R872 VDD1.n147 VDD1.n146 12.0247
R873 VDD1.n184 VDD1.n183 12.0247
R874 VDD1.n193 VDD1.n115 12.0247
R875 VDD1.n90 VDD1.n89 11.249
R876 VDD1.n73 VDD1.n14 11.249
R877 VDD1.n44 VDD1.n31 11.249
R878 VDD1.n150 VDD1.n137 11.249
R879 VDD1.n179 VDD1.n121 11.249
R880 VDD1.n197 VDD1.n196 11.249
R881 VDD1.n93 VDD1.n6 10.4732
R882 VDD1.n72 VDD1.n17 10.4732
R883 VDD1.n45 VDD1.n29 10.4732
R884 VDD1.n151 VDD1.n135 10.4732
R885 VDD1.n178 VDD1.n123 10.4732
R886 VDD1.n200 VDD1.n113 10.4732
R887 VDD1.n94 VDD1.n4 9.69747
R888 VDD1.n69 VDD1.n68 9.69747
R889 VDD1.n49 VDD1.n48 9.69747
R890 VDD1.n155 VDD1.n154 9.69747
R891 VDD1.n175 VDD1.n174 9.69747
R892 VDD1.n201 VDD1.n111 9.69747
R893 VDD1.n104 VDD1.n103 9.45567
R894 VDD1.n211 VDD1.n210 9.45567
R895 VDD1.n62 VDD1.n61 9.3005
R896 VDD1.n64 VDD1.n63 9.3005
R897 VDD1.n19 VDD1.n18 9.3005
R898 VDD1.n70 VDD1.n69 9.3005
R899 VDD1.n72 VDD1.n71 9.3005
R900 VDD1.n14 VDD1.n13 9.3005
R901 VDD1.n78 VDD1.n77 9.3005
R902 VDD1.n80 VDD1.n79 9.3005
R903 VDD1.n103 VDD1.n102 9.3005
R904 VDD1.n2 VDD1.n1 9.3005
R905 VDD1.n97 VDD1.n96 9.3005
R906 VDD1.n95 VDD1.n94 9.3005
R907 VDD1.n6 VDD1.n5 9.3005
R908 VDD1.n89 VDD1.n88 9.3005
R909 VDD1.n87 VDD1.n86 9.3005
R910 VDD1.n10 VDD1.n9 9.3005
R911 VDD1.n23 VDD1.n22 9.3005
R912 VDD1.n56 VDD1.n55 9.3005
R913 VDD1.n54 VDD1.n53 9.3005
R914 VDD1.n27 VDD1.n26 9.3005
R915 VDD1.n48 VDD1.n47 9.3005
R916 VDD1.n46 VDD1.n45 9.3005
R917 VDD1.n31 VDD1.n30 9.3005
R918 VDD1.n40 VDD1.n39 9.3005
R919 VDD1.n38 VDD1.n37 9.3005
R920 VDD1.n109 VDD1.n108 9.3005
R921 VDD1.n204 VDD1.n203 9.3005
R922 VDD1.n202 VDD1.n201 9.3005
R923 VDD1.n113 VDD1.n112 9.3005
R924 VDD1.n196 VDD1.n195 9.3005
R925 VDD1.n194 VDD1.n193 9.3005
R926 VDD1.n117 VDD1.n116 9.3005
R927 VDD1.n162 VDD1.n161 9.3005
R928 VDD1.n160 VDD1.n159 9.3005
R929 VDD1.n133 VDD1.n132 9.3005
R930 VDD1.n154 VDD1.n153 9.3005
R931 VDD1.n152 VDD1.n151 9.3005
R932 VDD1.n137 VDD1.n136 9.3005
R933 VDD1.n146 VDD1.n145 9.3005
R934 VDD1.n144 VDD1.n143 9.3005
R935 VDD1.n129 VDD1.n128 9.3005
R936 VDD1.n168 VDD1.n167 9.3005
R937 VDD1.n170 VDD1.n169 9.3005
R938 VDD1.n125 VDD1.n124 9.3005
R939 VDD1.n176 VDD1.n175 9.3005
R940 VDD1.n178 VDD1.n177 9.3005
R941 VDD1.n121 VDD1.n120 9.3005
R942 VDD1.n185 VDD1.n184 9.3005
R943 VDD1.n187 VDD1.n186 9.3005
R944 VDD1.n210 VDD1.n209 9.3005
R945 VDD1.n98 VDD1.n97 8.92171
R946 VDD1.n65 VDD1.n19 8.92171
R947 VDD1.n52 VDD1.n27 8.92171
R948 VDD1.n158 VDD1.n133 8.92171
R949 VDD1.n171 VDD1.n125 8.92171
R950 VDD1.n205 VDD1.n204 8.92171
R951 VDD1.n101 VDD1.n2 8.14595
R952 VDD1.n64 VDD1.n21 8.14595
R953 VDD1.n53 VDD1.n25 8.14595
R954 VDD1.n159 VDD1.n131 8.14595
R955 VDD1.n170 VDD1.n127 8.14595
R956 VDD1.n208 VDD1.n109 8.14595
R957 VDD1.n102 VDD1.n0 7.3702
R958 VDD1.n61 VDD1.n60 7.3702
R959 VDD1.n57 VDD1.n56 7.3702
R960 VDD1.n163 VDD1.n162 7.3702
R961 VDD1.n167 VDD1.n166 7.3702
R962 VDD1.n209 VDD1.n107 7.3702
R963 VDD1.n104 VDD1.n0 6.59444
R964 VDD1.n60 VDD1.n23 6.59444
R965 VDD1.n57 VDD1.n23 6.59444
R966 VDD1.n163 VDD1.n129 6.59444
R967 VDD1.n166 VDD1.n129 6.59444
R968 VDD1.n211 VDD1.n107 6.59444
R969 VDD1.n102 VDD1.n101 5.81868
R970 VDD1.n61 VDD1.n21 5.81868
R971 VDD1.n56 VDD1.n25 5.81868
R972 VDD1.n162 VDD1.n131 5.81868
R973 VDD1.n167 VDD1.n127 5.81868
R974 VDD1.n209 VDD1.n208 5.81868
R975 VDD1.n98 VDD1.n2 5.04292
R976 VDD1.n65 VDD1.n64 5.04292
R977 VDD1.n53 VDD1.n52 5.04292
R978 VDD1.n159 VDD1.n158 5.04292
R979 VDD1.n171 VDD1.n170 5.04292
R980 VDD1.n205 VDD1.n109 5.04292
R981 VDD1.n97 VDD1.n4 4.26717
R982 VDD1.n68 VDD1.n19 4.26717
R983 VDD1.n49 VDD1.n27 4.26717
R984 VDD1.n155 VDD1.n133 4.26717
R985 VDD1.n174 VDD1.n125 4.26717
R986 VDD1.n204 VDD1.n111 4.26717
R987 VDD1.n38 VDD1.n34 3.70982
R988 VDD1.n144 VDD1.n140 3.70982
R989 VDD1.n94 VDD1.n93 3.49141
R990 VDD1.n69 VDD1.n17 3.49141
R991 VDD1.n48 VDD1.n29 3.49141
R992 VDD1.n154 VDD1.n135 3.49141
R993 VDD1.n175 VDD1.n123 3.49141
R994 VDD1.n201 VDD1.n200 3.49141
R995 VDD1.n90 VDD1.n6 2.71565
R996 VDD1.n73 VDD1.n72 2.71565
R997 VDD1.n45 VDD1.n44 2.71565
R998 VDD1.n151 VDD1.n150 2.71565
R999 VDD1.n179 VDD1.n178 2.71565
R1000 VDD1.n197 VDD1.n113 2.71565
R1001 VDD1.n89 VDD1.n8 1.93989
R1002 VDD1.n76 VDD1.n14 1.93989
R1003 VDD1.n41 VDD1.n31 1.93989
R1004 VDD1.n147 VDD1.n137 1.93989
R1005 VDD1.n183 VDD1.n121 1.93989
R1006 VDD1.n196 VDD1.n115 1.93989
R1007 VDD1.n216 VDD1.t6 1.72582
R1008 VDD1.n216 VDD1.t9 1.72582
R1009 VDD1.n105 VDD1.t3 1.72582
R1010 VDD1.n105 VDD1.t4 1.72582
R1011 VDD1.n214 VDD1.t7 1.72582
R1012 VDD1.n214 VDD1.t1 1.72582
R1013 VDD1.n212 VDD1.t8 1.72582
R1014 VDD1.n212 VDD1.t0 1.72582
R1015 VDD1.n86 VDD1.n85 1.16414
R1016 VDD1.n77 VDD1.n12 1.16414
R1017 VDD1.n40 VDD1.n33 1.16414
R1018 VDD1.n146 VDD1.n139 1.16414
R1019 VDD1.n184 VDD1.n119 1.16414
R1020 VDD1.n193 VDD1.n192 1.16414
R1021 VDD1 VDD1.n217 0.853948
R1022 VDD1.n82 VDD1.n10 0.388379
R1023 VDD1.n81 VDD1.n80 0.388379
R1024 VDD1.n37 VDD1.n36 0.388379
R1025 VDD1.n143 VDD1.n142 0.388379
R1026 VDD1.n188 VDD1.n187 0.388379
R1027 VDD1.n189 VDD1.n117 0.388379
R1028 VDD1 VDD1.n106 0.362569
R1029 VDD1.n215 VDD1.n213 0.249033
R1030 VDD1.n103 VDD1.n1 0.155672
R1031 VDD1.n96 VDD1.n1 0.155672
R1032 VDD1.n96 VDD1.n95 0.155672
R1033 VDD1.n95 VDD1.n5 0.155672
R1034 VDD1.n88 VDD1.n5 0.155672
R1035 VDD1.n88 VDD1.n87 0.155672
R1036 VDD1.n87 VDD1.n9 0.155672
R1037 VDD1.n79 VDD1.n9 0.155672
R1038 VDD1.n79 VDD1.n78 0.155672
R1039 VDD1.n78 VDD1.n13 0.155672
R1040 VDD1.n71 VDD1.n13 0.155672
R1041 VDD1.n71 VDD1.n70 0.155672
R1042 VDD1.n70 VDD1.n18 0.155672
R1043 VDD1.n63 VDD1.n18 0.155672
R1044 VDD1.n63 VDD1.n62 0.155672
R1045 VDD1.n62 VDD1.n22 0.155672
R1046 VDD1.n55 VDD1.n22 0.155672
R1047 VDD1.n55 VDD1.n54 0.155672
R1048 VDD1.n54 VDD1.n26 0.155672
R1049 VDD1.n47 VDD1.n26 0.155672
R1050 VDD1.n47 VDD1.n46 0.155672
R1051 VDD1.n46 VDD1.n30 0.155672
R1052 VDD1.n39 VDD1.n30 0.155672
R1053 VDD1.n39 VDD1.n38 0.155672
R1054 VDD1.n145 VDD1.n144 0.155672
R1055 VDD1.n145 VDD1.n136 0.155672
R1056 VDD1.n152 VDD1.n136 0.155672
R1057 VDD1.n153 VDD1.n152 0.155672
R1058 VDD1.n153 VDD1.n132 0.155672
R1059 VDD1.n160 VDD1.n132 0.155672
R1060 VDD1.n161 VDD1.n160 0.155672
R1061 VDD1.n161 VDD1.n128 0.155672
R1062 VDD1.n168 VDD1.n128 0.155672
R1063 VDD1.n169 VDD1.n168 0.155672
R1064 VDD1.n169 VDD1.n124 0.155672
R1065 VDD1.n176 VDD1.n124 0.155672
R1066 VDD1.n177 VDD1.n176 0.155672
R1067 VDD1.n177 VDD1.n120 0.155672
R1068 VDD1.n185 VDD1.n120 0.155672
R1069 VDD1.n186 VDD1.n185 0.155672
R1070 VDD1.n186 VDD1.n116 0.155672
R1071 VDD1.n194 VDD1.n116 0.155672
R1072 VDD1.n195 VDD1.n194 0.155672
R1073 VDD1.n195 VDD1.n112 0.155672
R1074 VDD1.n202 VDD1.n112 0.155672
R1075 VDD1.n203 VDD1.n202 0.155672
R1076 VDD1.n203 VDD1.n108 0.155672
R1077 VDD1.n210 VDD1.n108 0.155672
R1078 VN.n4 VN.t9 477.848
R1079 VN.n23 VN.t5 477.848
R1080 VN.n17 VN.t7 456.784
R1081 VN.n36 VN.t1 456.784
R1082 VN.n10 VN.t8 420.411
R1083 VN.n5 VN.t4 420.411
R1084 VN.n1 VN.t2 420.411
R1085 VN.n29 VN.t3 420.411
R1086 VN.n24 VN.t6 420.411
R1087 VN.n20 VN.t0 420.411
R1088 VN.n35 VN.n19 161.3
R1089 VN.n34 VN.n33 161.3
R1090 VN.n32 VN.n31 161.3
R1091 VN.n30 VN.n21 161.3
R1092 VN.n29 VN.n28 161.3
R1093 VN.n27 VN.n22 161.3
R1094 VN.n26 VN.n25 161.3
R1095 VN.n16 VN.n0 161.3
R1096 VN.n15 VN.n14 161.3
R1097 VN.n13 VN.n12 161.3
R1098 VN.n11 VN.n2 161.3
R1099 VN.n10 VN.n9 161.3
R1100 VN.n8 VN.n3 161.3
R1101 VN.n7 VN.n6 161.3
R1102 VN.n37 VN.n36 80.6037
R1103 VN.n18 VN.n17 80.6037
R1104 VN.n6 VN.n3 56.5617
R1105 VN.n12 VN.n11 56.5617
R1106 VN.n25 VN.n22 56.5617
R1107 VN.n31 VN.n30 56.5617
R1108 VN VN.n37 50.4195
R1109 VN.n17 VN.n16 40.8975
R1110 VN.n36 VN.n35 40.8975
R1111 VN.n5 VN.n4 37.106
R1112 VN.n24 VN.n23 37.106
R1113 VN.n16 VN.n15 29.4362
R1114 VN.n35 VN.n34 29.4362
R1115 VN.n26 VN.n23 28.8662
R1116 VN.n7 VN.n4 28.8662
R1117 VN.n10 VN.n3 24.5923
R1118 VN.n11 VN.n10 24.5923
R1119 VN.n30 VN.n29 24.5923
R1120 VN.n29 VN.n22 24.5923
R1121 VN.n6 VN.n5 20.1658
R1122 VN.n12 VN.n1 20.1658
R1123 VN.n25 VN.n24 20.1658
R1124 VN.n31 VN.n20 20.1658
R1125 VN.n15 VN.n1 4.42703
R1126 VN.n34 VN.n20 4.42703
R1127 VN.n37 VN.n19 0.285035
R1128 VN.n18 VN.n0 0.285035
R1129 VN.n33 VN.n19 0.189894
R1130 VN.n33 VN.n32 0.189894
R1131 VN.n32 VN.n21 0.189894
R1132 VN.n28 VN.n21 0.189894
R1133 VN.n28 VN.n27 0.189894
R1134 VN.n27 VN.n26 0.189894
R1135 VN.n8 VN.n7 0.189894
R1136 VN.n9 VN.n8 0.189894
R1137 VN.n9 VN.n2 0.189894
R1138 VN.n13 VN.n2 0.189894
R1139 VN.n14 VN.n13 0.189894
R1140 VN.n14 VN.n0 0.189894
R1141 VN VN.n18 0.146778
R1142 VDD2.n209 VDD2.n109 756.745
R1143 VDD2.n100 VDD2.n0 756.745
R1144 VDD2.n210 VDD2.n209 585
R1145 VDD2.n208 VDD2.n207 585
R1146 VDD2.n113 VDD2.n112 585
R1147 VDD2.n202 VDD2.n201 585
R1148 VDD2.n200 VDD2.n199 585
R1149 VDD2.n117 VDD2.n116 585
R1150 VDD2.n194 VDD2.n193 585
R1151 VDD2.n192 VDD2.n191 585
R1152 VDD2.n190 VDD2.n120 585
R1153 VDD2.n124 VDD2.n121 585
R1154 VDD2.n185 VDD2.n184 585
R1155 VDD2.n183 VDD2.n182 585
R1156 VDD2.n126 VDD2.n125 585
R1157 VDD2.n177 VDD2.n176 585
R1158 VDD2.n175 VDD2.n174 585
R1159 VDD2.n130 VDD2.n129 585
R1160 VDD2.n169 VDD2.n168 585
R1161 VDD2.n167 VDD2.n166 585
R1162 VDD2.n134 VDD2.n133 585
R1163 VDD2.n161 VDD2.n160 585
R1164 VDD2.n159 VDD2.n158 585
R1165 VDD2.n138 VDD2.n137 585
R1166 VDD2.n153 VDD2.n152 585
R1167 VDD2.n151 VDD2.n150 585
R1168 VDD2.n142 VDD2.n141 585
R1169 VDD2.n145 VDD2.n144 585
R1170 VDD2.n35 VDD2.n34 585
R1171 VDD2.n32 VDD2.n31 585
R1172 VDD2.n41 VDD2.n40 585
R1173 VDD2.n43 VDD2.n42 585
R1174 VDD2.n28 VDD2.n27 585
R1175 VDD2.n49 VDD2.n48 585
R1176 VDD2.n51 VDD2.n50 585
R1177 VDD2.n24 VDD2.n23 585
R1178 VDD2.n57 VDD2.n56 585
R1179 VDD2.n59 VDD2.n58 585
R1180 VDD2.n20 VDD2.n19 585
R1181 VDD2.n65 VDD2.n64 585
R1182 VDD2.n67 VDD2.n66 585
R1183 VDD2.n16 VDD2.n15 585
R1184 VDD2.n73 VDD2.n72 585
R1185 VDD2.n76 VDD2.n75 585
R1186 VDD2.n74 VDD2.n12 585
R1187 VDD2.n81 VDD2.n11 585
R1188 VDD2.n83 VDD2.n82 585
R1189 VDD2.n85 VDD2.n84 585
R1190 VDD2.n8 VDD2.n7 585
R1191 VDD2.n91 VDD2.n90 585
R1192 VDD2.n93 VDD2.n92 585
R1193 VDD2.n4 VDD2.n3 585
R1194 VDD2.n99 VDD2.n98 585
R1195 VDD2.n101 VDD2.n100 585
R1196 VDD2.t8 VDD2.n143 327.466
R1197 VDD2.t0 VDD2.n33 327.466
R1198 VDD2.n209 VDD2.n208 171.744
R1199 VDD2.n208 VDD2.n112 171.744
R1200 VDD2.n201 VDD2.n112 171.744
R1201 VDD2.n201 VDD2.n200 171.744
R1202 VDD2.n200 VDD2.n116 171.744
R1203 VDD2.n193 VDD2.n116 171.744
R1204 VDD2.n193 VDD2.n192 171.744
R1205 VDD2.n192 VDD2.n120 171.744
R1206 VDD2.n124 VDD2.n120 171.744
R1207 VDD2.n184 VDD2.n124 171.744
R1208 VDD2.n184 VDD2.n183 171.744
R1209 VDD2.n183 VDD2.n125 171.744
R1210 VDD2.n176 VDD2.n125 171.744
R1211 VDD2.n176 VDD2.n175 171.744
R1212 VDD2.n175 VDD2.n129 171.744
R1213 VDD2.n168 VDD2.n129 171.744
R1214 VDD2.n168 VDD2.n167 171.744
R1215 VDD2.n167 VDD2.n133 171.744
R1216 VDD2.n160 VDD2.n133 171.744
R1217 VDD2.n160 VDD2.n159 171.744
R1218 VDD2.n159 VDD2.n137 171.744
R1219 VDD2.n152 VDD2.n137 171.744
R1220 VDD2.n152 VDD2.n151 171.744
R1221 VDD2.n151 VDD2.n141 171.744
R1222 VDD2.n144 VDD2.n141 171.744
R1223 VDD2.n34 VDD2.n31 171.744
R1224 VDD2.n41 VDD2.n31 171.744
R1225 VDD2.n42 VDD2.n41 171.744
R1226 VDD2.n42 VDD2.n27 171.744
R1227 VDD2.n49 VDD2.n27 171.744
R1228 VDD2.n50 VDD2.n49 171.744
R1229 VDD2.n50 VDD2.n23 171.744
R1230 VDD2.n57 VDD2.n23 171.744
R1231 VDD2.n58 VDD2.n57 171.744
R1232 VDD2.n58 VDD2.n19 171.744
R1233 VDD2.n65 VDD2.n19 171.744
R1234 VDD2.n66 VDD2.n65 171.744
R1235 VDD2.n66 VDD2.n15 171.744
R1236 VDD2.n73 VDD2.n15 171.744
R1237 VDD2.n75 VDD2.n73 171.744
R1238 VDD2.n75 VDD2.n74 171.744
R1239 VDD2.n74 VDD2.n11 171.744
R1240 VDD2.n83 VDD2.n11 171.744
R1241 VDD2.n84 VDD2.n83 171.744
R1242 VDD2.n84 VDD2.n7 171.744
R1243 VDD2.n91 VDD2.n7 171.744
R1244 VDD2.n92 VDD2.n91 171.744
R1245 VDD2.n92 VDD2.n3 171.744
R1246 VDD2.n99 VDD2.n3 171.744
R1247 VDD2.n100 VDD2.n99 171.744
R1248 VDD2.n144 VDD2.t8 85.8723
R1249 VDD2.n34 VDD2.t0 85.8723
R1250 VDD2.n108 VDD2.n107 66.9139
R1251 VDD2 VDD2.n217 66.9109
R1252 VDD2.n216 VDD2.n215 66.0577
R1253 VDD2.n106 VDD2.n105 66.0577
R1254 VDD2.n106 VDD2.n104 47.7524
R1255 VDD2.n214 VDD2.n213 46.5369
R1256 VDD2.n214 VDD2.n108 45.7304
R1257 VDD2.n145 VDD2.n143 16.3895
R1258 VDD2.n35 VDD2.n33 16.3895
R1259 VDD2.n191 VDD2.n190 13.1884
R1260 VDD2.n82 VDD2.n81 13.1884
R1261 VDD2.n194 VDD2.n119 12.8005
R1262 VDD2.n189 VDD2.n121 12.8005
R1263 VDD2.n146 VDD2.n142 12.8005
R1264 VDD2.n36 VDD2.n32 12.8005
R1265 VDD2.n80 VDD2.n12 12.8005
R1266 VDD2.n85 VDD2.n10 12.8005
R1267 VDD2.n195 VDD2.n117 12.0247
R1268 VDD2.n186 VDD2.n185 12.0247
R1269 VDD2.n150 VDD2.n149 12.0247
R1270 VDD2.n40 VDD2.n39 12.0247
R1271 VDD2.n77 VDD2.n76 12.0247
R1272 VDD2.n86 VDD2.n8 12.0247
R1273 VDD2.n199 VDD2.n198 11.249
R1274 VDD2.n182 VDD2.n123 11.249
R1275 VDD2.n153 VDD2.n140 11.249
R1276 VDD2.n43 VDD2.n30 11.249
R1277 VDD2.n72 VDD2.n14 11.249
R1278 VDD2.n90 VDD2.n89 11.249
R1279 VDD2.n202 VDD2.n115 10.4732
R1280 VDD2.n181 VDD2.n126 10.4732
R1281 VDD2.n154 VDD2.n138 10.4732
R1282 VDD2.n44 VDD2.n28 10.4732
R1283 VDD2.n71 VDD2.n16 10.4732
R1284 VDD2.n93 VDD2.n6 10.4732
R1285 VDD2.n203 VDD2.n113 9.69747
R1286 VDD2.n178 VDD2.n177 9.69747
R1287 VDD2.n158 VDD2.n157 9.69747
R1288 VDD2.n48 VDD2.n47 9.69747
R1289 VDD2.n68 VDD2.n67 9.69747
R1290 VDD2.n94 VDD2.n4 9.69747
R1291 VDD2.n213 VDD2.n212 9.45567
R1292 VDD2.n104 VDD2.n103 9.45567
R1293 VDD2.n171 VDD2.n170 9.3005
R1294 VDD2.n173 VDD2.n172 9.3005
R1295 VDD2.n128 VDD2.n127 9.3005
R1296 VDD2.n179 VDD2.n178 9.3005
R1297 VDD2.n181 VDD2.n180 9.3005
R1298 VDD2.n123 VDD2.n122 9.3005
R1299 VDD2.n187 VDD2.n186 9.3005
R1300 VDD2.n189 VDD2.n188 9.3005
R1301 VDD2.n212 VDD2.n211 9.3005
R1302 VDD2.n111 VDD2.n110 9.3005
R1303 VDD2.n206 VDD2.n205 9.3005
R1304 VDD2.n204 VDD2.n203 9.3005
R1305 VDD2.n115 VDD2.n114 9.3005
R1306 VDD2.n198 VDD2.n197 9.3005
R1307 VDD2.n196 VDD2.n195 9.3005
R1308 VDD2.n119 VDD2.n118 9.3005
R1309 VDD2.n132 VDD2.n131 9.3005
R1310 VDD2.n165 VDD2.n164 9.3005
R1311 VDD2.n163 VDD2.n162 9.3005
R1312 VDD2.n136 VDD2.n135 9.3005
R1313 VDD2.n157 VDD2.n156 9.3005
R1314 VDD2.n155 VDD2.n154 9.3005
R1315 VDD2.n140 VDD2.n139 9.3005
R1316 VDD2.n149 VDD2.n148 9.3005
R1317 VDD2.n147 VDD2.n146 9.3005
R1318 VDD2.n2 VDD2.n1 9.3005
R1319 VDD2.n97 VDD2.n96 9.3005
R1320 VDD2.n95 VDD2.n94 9.3005
R1321 VDD2.n6 VDD2.n5 9.3005
R1322 VDD2.n89 VDD2.n88 9.3005
R1323 VDD2.n87 VDD2.n86 9.3005
R1324 VDD2.n10 VDD2.n9 9.3005
R1325 VDD2.n55 VDD2.n54 9.3005
R1326 VDD2.n53 VDD2.n52 9.3005
R1327 VDD2.n26 VDD2.n25 9.3005
R1328 VDD2.n47 VDD2.n46 9.3005
R1329 VDD2.n45 VDD2.n44 9.3005
R1330 VDD2.n30 VDD2.n29 9.3005
R1331 VDD2.n39 VDD2.n38 9.3005
R1332 VDD2.n37 VDD2.n36 9.3005
R1333 VDD2.n22 VDD2.n21 9.3005
R1334 VDD2.n61 VDD2.n60 9.3005
R1335 VDD2.n63 VDD2.n62 9.3005
R1336 VDD2.n18 VDD2.n17 9.3005
R1337 VDD2.n69 VDD2.n68 9.3005
R1338 VDD2.n71 VDD2.n70 9.3005
R1339 VDD2.n14 VDD2.n13 9.3005
R1340 VDD2.n78 VDD2.n77 9.3005
R1341 VDD2.n80 VDD2.n79 9.3005
R1342 VDD2.n103 VDD2.n102 9.3005
R1343 VDD2.n207 VDD2.n206 8.92171
R1344 VDD2.n174 VDD2.n128 8.92171
R1345 VDD2.n161 VDD2.n136 8.92171
R1346 VDD2.n51 VDD2.n26 8.92171
R1347 VDD2.n64 VDD2.n18 8.92171
R1348 VDD2.n98 VDD2.n97 8.92171
R1349 VDD2.n210 VDD2.n111 8.14595
R1350 VDD2.n173 VDD2.n130 8.14595
R1351 VDD2.n162 VDD2.n134 8.14595
R1352 VDD2.n52 VDD2.n24 8.14595
R1353 VDD2.n63 VDD2.n20 8.14595
R1354 VDD2.n101 VDD2.n2 8.14595
R1355 VDD2.n211 VDD2.n109 7.3702
R1356 VDD2.n170 VDD2.n169 7.3702
R1357 VDD2.n166 VDD2.n165 7.3702
R1358 VDD2.n56 VDD2.n55 7.3702
R1359 VDD2.n60 VDD2.n59 7.3702
R1360 VDD2.n102 VDD2.n0 7.3702
R1361 VDD2.n213 VDD2.n109 6.59444
R1362 VDD2.n169 VDD2.n132 6.59444
R1363 VDD2.n166 VDD2.n132 6.59444
R1364 VDD2.n56 VDD2.n22 6.59444
R1365 VDD2.n59 VDD2.n22 6.59444
R1366 VDD2.n104 VDD2.n0 6.59444
R1367 VDD2.n211 VDD2.n210 5.81868
R1368 VDD2.n170 VDD2.n130 5.81868
R1369 VDD2.n165 VDD2.n134 5.81868
R1370 VDD2.n55 VDD2.n24 5.81868
R1371 VDD2.n60 VDD2.n20 5.81868
R1372 VDD2.n102 VDD2.n101 5.81868
R1373 VDD2.n207 VDD2.n111 5.04292
R1374 VDD2.n174 VDD2.n173 5.04292
R1375 VDD2.n162 VDD2.n161 5.04292
R1376 VDD2.n52 VDD2.n51 5.04292
R1377 VDD2.n64 VDD2.n63 5.04292
R1378 VDD2.n98 VDD2.n2 5.04292
R1379 VDD2.n206 VDD2.n113 4.26717
R1380 VDD2.n177 VDD2.n128 4.26717
R1381 VDD2.n158 VDD2.n136 4.26717
R1382 VDD2.n48 VDD2.n26 4.26717
R1383 VDD2.n67 VDD2.n18 4.26717
R1384 VDD2.n97 VDD2.n4 4.26717
R1385 VDD2.n147 VDD2.n143 3.70982
R1386 VDD2.n37 VDD2.n33 3.70982
R1387 VDD2.n203 VDD2.n202 3.49141
R1388 VDD2.n178 VDD2.n126 3.49141
R1389 VDD2.n157 VDD2.n138 3.49141
R1390 VDD2.n47 VDD2.n28 3.49141
R1391 VDD2.n68 VDD2.n16 3.49141
R1392 VDD2.n94 VDD2.n93 3.49141
R1393 VDD2.n199 VDD2.n115 2.71565
R1394 VDD2.n182 VDD2.n181 2.71565
R1395 VDD2.n154 VDD2.n153 2.71565
R1396 VDD2.n44 VDD2.n43 2.71565
R1397 VDD2.n72 VDD2.n71 2.71565
R1398 VDD2.n90 VDD2.n6 2.71565
R1399 VDD2.n198 VDD2.n117 1.93989
R1400 VDD2.n185 VDD2.n123 1.93989
R1401 VDD2.n150 VDD2.n140 1.93989
R1402 VDD2.n40 VDD2.n30 1.93989
R1403 VDD2.n76 VDD2.n14 1.93989
R1404 VDD2.n89 VDD2.n8 1.93989
R1405 VDD2.n217 VDD2.t3 1.72582
R1406 VDD2.n217 VDD2.t4 1.72582
R1407 VDD2.n215 VDD2.t9 1.72582
R1408 VDD2.n215 VDD2.t6 1.72582
R1409 VDD2.n107 VDD2.t7 1.72582
R1410 VDD2.n107 VDD2.t2 1.72582
R1411 VDD2.n105 VDD2.t5 1.72582
R1412 VDD2.n105 VDD2.t1 1.72582
R1413 VDD2.n216 VDD2.n214 1.21602
R1414 VDD2.n195 VDD2.n194 1.16414
R1415 VDD2.n186 VDD2.n121 1.16414
R1416 VDD2.n149 VDD2.n142 1.16414
R1417 VDD2.n39 VDD2.n32 1.16414
R1418 VDD2.n77 VDD2.n12 1.16414
R1419 VDD2.n86 VDD2.n85 1.16414
R1420 VDD2.n191 VDD2.n119 0.388379
R1421 VDD2.n190 VDD2.n189 0.388379
R1422 VDD2.n146 VDD2.n145 0.388379
R1423 VDD2.n36 VDD2.n35 0.388379
R1424 VDD2.n81 VDD2.n80 0.388379
R1425 VDD2.n82 VDD2.n10 0.388379
R1426 VDD2 VDD2.n216 0.362569
R1427 VDD2.n108 VDD2.n106 0.249033
R1428 VDD2.n212 VDD2.n110 0.155672
R1429 VDD2.n205 VDD2.n110 0.155672
R1430 VDD2.n205 VDD2.n204 0.155672
R1431 VDD2.n204 VDD2.n114 0.155672
R1432 VDD2.n197 VDD2.n114 0.155672
R1433 VDD2.n197 VDD2.n196 0.155672
R1434 VDD2.n196 VDD2.n118 0.155672
R1435 VDD2.n188 VDD2.n118 0.155672
R1436 VDD2.n188 VDD2.n187 0.155672
R1437 VDD2.n187 VDD2.n122 0.155672
R1438 VDD2.n180 VDD2.n122 0.155672
R1439 VDD2.n180 VDD2.n179 0.155672
R1440 VDD2.n179 VDD2.n127 0.155672
R1441 VDD2.n172 VDD2.n127 0.155672
R1442 VDD2.n172 VDD2.n171 0.155672
R1443 VDD2.n171 VDD2.n131 0.155672
R1444 VDD2.n164 VDD2.n131 0.155672
R1445 VDD2.n164 VDD2.n163 0.155672
R1446 VDD2.n163 VDD2.n135 0.155672
R1447 VDD2.n156 VDD2.n135 0.155672
R1448 VDD2.n156 VDD2.n155 0.155672
R1449 VDD2.n155 VDD2.n139 0.155672
R1450 VDD2.n148 VDD2.n139 0.155672
R1451 VDD2.n148 VDD2.n147 0.155672
R1452 VDD2.n38 VDD2.n37 0.155672
R1453 VDD2.n38 VDD2.n29 0.155672
R1454 VDD2.n45 VDD2.n29 0.155672
R1455 VDD2.n46 VDD2.n45 0.155672
R1456 VDD2.n46 VDD2.n25 0.155672
R1457 VDD2.n53 VDD2.n25 0.155672
R1458 VDD2.n54 VDD2.n53 0.155672
R1459 VDD2.n54 VDD2.n21 0.155672
R1460 VDD2.n61 VDD2.n21 0.155672
R1461 VDD2.n62 VDD2.n61 0.155672
R1462 VDD2.n62 VDD2.n17 0.155672
R1463 VDD2.n69 VDD2.n17 0.155672
R1464 VDD2.n70 VDD2.n69 0.155672
R1465 VDD2.n70 VDD2.n13 0.155672
R1466 VDD2.n78 VDD2.n13 0.155672
R1467 VDD2.n79 VDD2.n78 0.155672
R1468 VDD2.n79 VDD2.n9 0.155672
R1469 VDD2.n87 VDD2.n9 0.155672
R1470 VDD2.n88 VDD2.n87 0.155672
R1471 VDD2.n88 VDD2.n5 0.155672
R1472 VDD2.n95 VDD2.n5 0.155672
R1473 VDD2.n96 VDD2.n95 0.155672
R1474 VDD2.n96 VDD2.n1 0.155672
R1475 VDD2.n103 VDD2.n1 0.155672
R1476 B.n154 B.t0 623.851
R1477 B.n162 B.t3 623.851
R1478 B.n50 B.t6 623.851
R1479 B.n56 B.t9 623.851
R1480 B.n560 B.n89 585
R1481 B.n562 B.n561 585
R1482 B.n563 B.n88 585
R1483 B.n565 B.n564 585
R1484 B.n566 B.n87 585
R1485 B.n568 B.n567 585
R1486 B.n569 B.n86 585
R1487 B.n571 B.n570 585
R1488 B.n572 B.n85 585
R1489 B.n574 B.n573 585
R1490 B.n575 B.n84 585
R1491 B.n577 B.n576 585
R1492 B.n578 B.n83 585
R1493 B.n580 B.n579 585
R1494 B.n581 B.n82 585
R1495 B.n583 B.n582 585
R1496 B.n584 B.n81 585
R1497 B.n586 B.n585 585
R1498 B.n587 B.n80 585
R1499 B.n589 B.n588 585
R1500 B.n590 B.n79 585
R1501 B.n592 B.n591 585
R1502 B.n593 B.n78 585
R1503 B.n595 B.n594 585
R1504 B.n596 B.n77 585
R1505 B.n598 B.n597 585
R1506 B.n599 B.n76 585
R1507 B.n601 B.n600 585
R1508 B.n602 B.n75 585
R1509 B.n604 B.n603 585
R1510 B.n605 B.n74 585
R1511 B.n607 B.n606 585
R1512 B.n608 B.n73 585
R1513 B.n610 B.n609 585
R1514 B.n611 B.n72 585
R1515 B.n613 B.n612 585
R1516 B.n614 B.n71 585
R1517 B.n616 B.n615 585
R1518 B.n617 B.n70 585
R1519 B.n619 B.n618 585
R1520 B.n620 B.n69 585
R1521 B.n622 B.n621 585
R1522 B.n623 B.n68 585
R1523 B.n625 B.n624 585
R1524 B.n626 B.n67 585
R1525 B.n628 B.n627 585
R1526 B.n629 B.n66 585
R1527 B.n631 B.n630 585
R1528 B.n632 B.n65 585
R1529 B.n634 B.n633 585
R1530 B.n635 B.n64 585
R1531 B.n637 B.n636 585
R1532 B.n638 B.n63 585
R1533 B.n640 B.n639 585
R1534 B.n641 B.n62 585
R1535 B.n643 B.n642 585
R1536 B.n644 B.n61 585
R1537 B.n646 B.n645 585
R1538 B.n647 B.n60 585
R1539 B.n649 B.n648 585
R1540 B.n650 B.n59 585
R1541 B.n652 B.n651 585
R1542 B.n654 B.n653 585
R1543 B.n655 B.n55 585
R1544 B.n657 B.n656 585
R1545 B.n658 B.n54 585
R1546 B.n660 B.n659 585
R1547 B.n661 B.n53 585
R1548 B.n663 B.n662 585
R1549 B.n664 B.n52 585
R1550 B.n666 B.n665 585
R1551 B.n668 B.n49 585
R1552 B.n670 B.n669 585
R1553 B.n671 B.n48 585
R1554 B.n673 B.n672 585
R1555 B.n674 B.n47 585
R1556 B.n676 B.n675 585
R1557 B.n677 B.n46 585
R1558 B.n679 B.n678 585
R1559 B.n680 B.n45 585
R1560 B.n682 B.n681 585
R1561 B.n683 B.n44 585
R1562 B.n685 B.n684 585
R1563 B.n686 B.n43 585
R1564 B.n688 B.n687 585
R1565 B.n689 B.n42 585
R1566 B.n691 B.n690 585
R1567 B.n692 B.n41 585
R1568 B.n694 B.n693 585
R1569 B.n695 B.n40 585
R1570 B.n697 B.n696 585
R1571 B.n698 B.n39 585
R1572 B.n700 B.n699 585
R1573 B.n701 B.n38 585
R1574 B.n703 B.n702 585
R1575 B.n704 B.n37 585
R1576 B.n706 B.n705 585
R1577 B.n707 B.n36 585
R1578 B.n709 B.n708 585
R1579 B.n710 B.n35 585
R1580 B.n712 B.n711 585
R1581 B.n713 B.n34 585
R1582 B.n715 B.n714 585
R1583 B.n716 B.n33 585
R1584 B.n718 B.n717 585
R1585 B.n719 B.n32 585
R1586 B.n721 B.n720 585
R1587 B.n722 B.n31 585
R1588 B.n724 B.n723 585
R1589 B.n725 B.n30 585
R1590 B.n727 B.n726 585
R1591 B.n728 B.n29 585
R1592 B.n730 B.n729 585
R1593 B.n731 B.n28 585
R1594 B.n733 B.n732 585
R1595 B.n734 B.n27 585
R1596 B.n736 B.n735 585
R1597 B.n737 B.n26 585
R1598 B.n739 B.n738 585
R1599 B.n740 B.n25 585
R1600 B.n742 B.n741 585
R1601 B.n743 B.n24 585
R1602 B.n745 B.n744 585
R1603 B.n746 B.n23 585
R1604 B.n748 B.n747 585
R1605 B.n749 B.n22 585
R1606 B.n751 B.n750 585
R1607 B.n752 B.n21 585
R1608 B.n754 B.n753 585
R1609 B.n755 B.n20 585
R1610 B.n757 B.n756 585
R1611 B.n758 B.n19 585
R1612 B.n760 B.n759 585
R1613 B.n559 B.n558 585
R1614 B.n557 B.n90 585
R1615 B.n556 B.n555 585
R1616 B.n554 B.n91 585
R1617 B.n553 B.n552 585
R1618 B.n551 B.n92 585
R1619 B.n550 B.n549 585
R1620 B.n548 B.n93 585
R1621 B.n547 B.n546 585
R1622 B.n545 B.n94 585
R1623 B.n544 B.n543 585
R1624 B.n542 B.n95 585
R1625 B.n541 B.n540 585
R1626 B.n539 B.n96 585
R1627 B.n538 B.n537 585
R1628 B.n536 B.n97 585
R1629 B.n535 B.n534 585
R1630 B.n533 B.n98 585
R1631 B.n532 B.n531 585
R1632 B.n530 B.n99 585
R1633 B.n529 B.n528 585
R1634 B.n527 B.n100 585
R1635 B.n526 B.n525 585
R1636 B.n524 B.n101 585
R1637 B.n523 B.n522 585
R1638 B.n521 B.n102 585
R1639 B.n520 B.n519 585
R1640 B.n518 B.n103 585
R1641 B.n517 B.n516 585
R1642 B.n515 B.n104 585
R1643 B.n514 B.n513 585
R1644 B.n512 B.n105 585
R1645 B.n511 B.n510 585
R1646 B.n509 B.n106 585
R1647 B.n508 B.n507 585
R1648 B.n506 B.n107 585
R1649 B.n505 B.n504 585
R1650 B.n503 B.n108 585
R1651 B.n502 B.n501 585
R1652 B.n500 B.n109 585
R1653 B.n499 B.n498 585
R1654 B.n497 B.n110 585
R1655 B.n496 B.n495 585
R1656 B.n494 B.n111 585
R1657 B.n493 B.n492 585
R1658 B.n491 B.n112 585
R1659 B.n490 B.n489 585
R1660 B.n488 B.n113 585
R1661 B.n487 B.n486 585
R1662 B.n485 B.n114 585
R1663 B.n484 B.n483 585
R1664 B.n482 B.n115 585
R1665 B.n481 B.n480 585
R1666 B.n479 B.n116 585
R1667 B.n478 B.n477 585
R1668 B.n476 B.n117 585
R1669 B.n475 B.n474 585
R1670 B.n473 B.n118 585
R1671 B.n472 B.n471 585
R1672 B.n470 B.n119 585
R1673 B.n469 B.n468 585
R1674 B.n467 B.n120 585
R1675 B.n466 B.n465 585
R1676 B.n464 B.n121 585
R1677 B.n463 B.n462 585
R1678 B.n461 B.n122 585
R1679 B.n460 B.n459 585
R1680 B.n259 B.n258 585
R1681 B.n260 B.n193 585
R1682 B.n262 B.n261 585
R1683 B.n263 B.n192 585
R1684 B.n265 B.n264 585
R1685 B.n266 B.n191 585
R1686 B.n268 B.n267 585
R1687 B.n269 B.n190 585
R1688 B.n271 B.n270 585
R1689 B.n272 B.n189 585
R1690 B.n274 B.n273 585
R1691 B.n275 B.n188 585
R1692 B.n277 B.n276 585
R1693 B.n278 B.n187 585
R1694 B.n280 B.n279 585
R1695 B.n281 B.n186 585
R1696 B.n283 B.n282 585
R1697 B.n284 B.n185 585
R1698 B.n286 B.n285 585
R1699 B.n287 B.n184 585
R1700 B.n289 B.n288 585
R1701 B.n290 B.n183 585
R1702 B.n292 B.n291 585
R1703 B.n293 B.n182 585
R1704 B.n295 B.n294 585
R1705 B.n296 B.n181 585
R1706 B.n298 B.n297 585
R1707 B.n299 B.n180 585
R1708 B.n301 B.n300 585
R1709 B.n302 B.n179 585
R1710 B.n304 B.n303 585
R1711 B.n305 B.n178 585
R1712 B.n307 B.n306 585
R1713 B.n308 B.n177 585
R1714 B.n310 B.n309 585
R1715 B.n311 B.n176 585
R1716 B.n313 B.n312 585
R1717 B.n314 B.n175 585
R1718 B.n316 B.n315 585
R1719 B.n317 B.n174 585
R1720 B.n319 B.n318 585
R1721 B.n320 B.n173 585
R1722 B.n322 B.n321 585
R1723 B.n323 B.n172 585
R1724 B.n325 B.n324 585
R1725 B.n326 B.n171 585
R1726 B.n328 B.n327 585
R1727 B.n329 B.n170 585
R1728 B.n331 B.n330 585
R1729 B.n332 B.n169 585
R1730 B.n334 B.n333 585
R1731 B.n335 B.n168 585
R1732 B.n337 B.n336 585
R1733 B.n338 B.n167 585
R1734 B.n340 B.n339 585
R1735 B.n341 B.n166 585
R1736 B.n343 B.n342 585
R1737 B.n344 B.n165 585
R1738 B.n346 B.n345 585
R1739 B.n347 B.n164 585
R1740 B.n349 B.n348 585
R1741 B.n350 B.n161 585
R1742 B.n353 B.n352 585
R1743 B.n354 B.n160 585
R1744 B.n356 B.n355 585
R1745 B.n357 B.n159 585
R1746 B.n359 B.n358 585
R1747 B.n360 B.n158 585
R1748 B.n362 B.n361 585
R1749 B.n363 B.n157 585
R1750 B.n365 B.n364 585
R1751 B.n367 B.n366 585
R1752 B.n368 B.n153 585
R1753 B.n370 B.n369 585
R1754 B.n371 B.n152 585
R1755 B.n373 B.n372 585
R1756 B.n374 B.n151 585
R1757 B.n376 B.n375 585
R1758 B.n377 B.n150 585
R1759 B.n379 B.n378 585
R1760 B.n380 B.n149 585
R1761 B.n382 B.n381 585
R1762 B.n383 B.n148 585
R1763 B.n385 B.n384 585
R1764 B.n386 B.n147 585
R1765 B.n388 B.n387 585
R1766 B.n389 B.n146 585
R1767 B.n391 B.n390 585
R1768 B.n392 B.n145 585
R1769 B.n394 B.n393 585
R1770 B.n395 B.n144 585
R1771 B.n397 B.n396 585
R1772 B.n398 B.n143 585
R1773 B.n400 B.n399 585
R1774 B.n401 B.n142 585
R1775 B.n403 B.n402 585
R1776 B.n404 B.n141 585
R1777 B.n406 B.n405 585
R1778 B.n407 B.n140 585
R1779 B.n409 B.n408 585
R1780 B.n410 B.n139 585
R1781 B.n412 B.n411 585
R1782 B.n413 B.n138 585
R1783 B.n415 B.n414 585
R1784 B.n416 B.n137 585
R1785 B.n418 B.n417 585
R1786 B.n419 B.n136 585
R1787 B.n421 B.n420 585
R1788 B.n422 B.n135 585
R1789 B.n424 B.n423 585
R1790 B.n425 B.n134 585
R1791 B.n427 B.n426 585
R1792 B.n428 B.n133 585
R1793 B.n430 B.n429 585
R1794 B.n431 B.n132 585
R1795 B.n433 B.n432 585
R1796 B.n434 B.n131 585
R1797 B.n436 B.n435 585
R1798 B.n437 B.n130 585
R1799 B.n439 B.n438 585
R1800 B.n440 B.n129 585
R1801 B.n442 B.n441 585
R1802 B.n443 B.n128 585
R1803 B.n445 B.n444 585
R1804 B.n446 B.n127 585
R1805 B.n448 B.n447 585
R1806 B.n449 B.n126 585
R1807 B.n451 B.n450 585
R1808 B.n452 B.n125 585
R1809 B.n454 B.n453 585
R1810 B.n455 B.n124 585
R1811 B.n457 B.n456 585
R1812 B.n458 B.n123 585
R1813 B.n257 B.n194 585
R1814 B.n256 B.n255 585
R1815 B.n254 B.n195 585
R1816 B.n253 B.n252 585
R1817 B.n251 B.n196 585
R1818 B.n250 B.n249 585
R1819 B.n248 B.n197 585
R1820 B.n247 B.n246 585
R1821 B.n245 B.n198 585
R1822 B.n244 B.n243 585
R1823 B.n242 B.n199 585
R1824 B.n241 B.n240 585
R1825 B.n239 B.n200 585
R1826 B.n238 B.n237 585
R1827 B.n236 B.n201 585
R1828 B.n235 B.n234 585
R1829 B.n233 B.n202 585
R1830 B.n232 B.n231 585
R1831 B.n230 B.n203 585
R1832 B.n229 B.n228 585
R1833 B.n227 B.n204 585
R1834 B.n226 B.n225 585
R1835 B.n224 B.n205 585
R1836 B.n223 B.n222 585
R1837 B.n221 B.n206 585
R1838 B.n220 B.n219 585
R1839 B.n218 B.n207 585
R1840 B.n217 B.n216 585
R1841 B.n215 B.n208 585
R1842 B.n214 B.n213 585
R1843 B.n212 B.n209 585
R1844 B.n211 B.n210 585
R1845 B.n2 B.n0 585
R1846 B.n809 B.n1 585
R1847 B.n808 B.n807 585
R1848 B.n806 B.n3 585
R1849 B.n805 B.n804 585
R1850 B.n803 B.n4 585
R1851 B.n802 B.n801 585
R1852 B.n800 B.n5 585
R1853 B.n799 B.n798 585
R1854 B.n797 B.n6 585
R1855 B.n796 B.n795 585
R1856 B.n794 B.n7 585
R1857 B.n793 B.n792 585
R1858 B.n791 B.n8 585
R1859 B.n790 B.n789 585
R1860 B.n788 B.n9 585
R1861 B.n787 B.n786 585
R1862 B.n785 B.n10 585
R1863 B.n784 B.n783 585
R1864 B.n782 B.n11 585
R1865 B.n781 B.n780 585
R1866 B.n779 B.n12 585
R1867 B.n778 B.n777 585
R1868 B.n776 B.n13 585
R1869 B.n775 B.n774 585
R1870 B.n773 B.n14 585
R1871 B.n772 B.n771 585
R1872 B.n770 B.n15 585
R1873 B.n769 B.n768 585
R1874 B.n767 B.n16 585
R1875 B.n766 B.n765 585
R1876 B.n764 B.n17 585
R1877 B.n763 B.n762 585
R1878 B.n761 B.n18 585
R1879 B.n811 B.n810 585
R1880 B.n154 B.t2 526.131
R1881 B.n56 B.t10 526.131
R1882 B.n162 B.t5 526.131
R1883 B.n50 B.t7 526.131
R1884 B.n258 B.n257 502.111
R1885 B.n761 B.n760 502.111
R1886 B.n460 B.n123 502.111
R1887 B.n558 B.n89 502.111
R1888 B.n155 B.t1 498.786
R1889 B.n57 B.t11 498.786
R1890 B.n163 B.t4 498.786
R1891 B.n51 B.t8 498.786
R1892 B.n257 B.n256 163.367
R1893 B.n256 B.n195 163.367
R1894 B.n252 B.n195 163.367
R1895 B.n252 B.n251 163.367
R1896 B.n251 B.n250 163.367
R1897 B.n250 B.n197 163.367
R1898 B.n246 B.n197 163.367
R1899 B.n246 B.n245 163.367
R1900 B.n245 B.n244 163.367
R1901 B.n244 B.n199 163.367
R1902 B.n240 B.n199 163.367
R1903 B.n240 B.n239 163.367
R1904 B.n239 B.n238 163.367
R1905 B.n238 B.n201 163.367
R1906 B.n234 B.n201 163.367
R1907 B.n234 B.n233 163.367
R1908 B.n233 B.n232 163.367
R1909 B.n232 B.n203 163.367
R1910 B.n228 B.n203 163.367
R1911 B.n228 B.n227 163.367
R1912 B.n227 B.n226 163.367
R1913 B.n226 B.n205 163.367
R1914 B.n222 B.n205 163.367
R1915 B.n222 B.n221 163.367
R1916 B.n221 B.n220 163.367
R1917 B.n220 B.n207 163.367
R1918 B.n216 B.n207 163.367
R1919 B.n216 B.n215 163.367
R1920 B.n215 B.n214 163.367
R1921 B.n214 B.n209 163.367
R1922 B.n210 B.n209 163.367
R1923 B.n210 B.n2 163.367
R1924 B.n810 B.n2 163.367
R1925 B.n810 B.n809 163.367
R1926 B.n809 B.n808 163.367
R1927 B.n808 B.n3 163.367
R1928 B.n804 B.n3 163.367
R1929 B.n804 B.n803 163.367
R1930 B.n803 B.n802 163.367
R1931 B.n802 B.n5 163.367
R1932 B.n798 B.n5 163.367
R1933 B.n798 B.n797 163.367
R1934 B.n797 B.n796 163.367
R1935 B.n796 B.n7 163.367
R1936 B.n792 B.n7 163.367
R1937 B.n792 B.n791 163.367
R1938 B.n791 B.n790 163.367
R1939 B.n790 B.n9 163.367
R1940 B.n786 B.n9 163.367
R1941 B.n786 B.n785 163.367
R1942 B.n785 B.n784 163.367
R1943 B.n784 B.n11 163.367
R1944 B.n780 B.n11 163.367
R1945 B.n780 B.n779 163.367
R1946 B.n779 B.n778 163.367
R1947 B.n778 B.n13 163.367
R1948 B.n774 B.n13 163.367
R1949 B.n774 B.n773 163.367
R1950 B.n773 B.n772 163.367
R1951 B.n772 B.n15 163.367
R1952 B.n768 B.n15 163.367
R1953 B.n768 B.n767 163.367
R1954 B.n767 B.n766 163.367
R1955 B.n766 B.n17 163.367
R1956 B.n762 B.n17 163.367
R1957 B.n762 B.n761 163.367
R1958 B.n258 B.n193 163.367
R1959 B.n262 B.n193 163.367
R1960 B.n263 B.n262 163.367
R1961 B.n264 B.n263 163.367
R1962 B.n264 B.n191 163.367
R1963 B.n268 B.n191 163.367
R1964 B.n269 B.n268 163.367
R1965 B.n270 B.n269 163.367
R1966 B.n270 B.n189 163.367
R1967 B.n274 B.n189 163.367
R1968 B.n275 B.n274 163.367
R1969 B.n276 B.n275 163.367
R1970 B.n276 B.n187 163.367
R1971 B.n280 B.n187 163.367
R1972 B.n281 B.n280 163.367
R1973 B.n282 B.n281 163.367
R1974 B.n282 B.n185 163.367
R1975 B.n286 B.n185 163.367
R1976 B.n287 B.n286 163.367
R1977 B.n288 B.n287 163.367
R1978 B.n288 B.n183 163.367
R1979 B.n292 B.n183 163.367
R1980 B.n293 B.n292 163.367
R1981 B.n294 B.n293 163.367
R1982 B.n294 B.n181 163.367
R1983 B.n298 B.n181 163.367
R1984 B.n299 B.n298 163.367
R1985 B.n300 B.n299 163.367
R1986 B.n300 B.n179 163.367
R1987 B.n304 B.n179 163.367
R1988 B.n305 B.n304 163.367
R1989 B.n306 B.n305 163.367
R1990 B.n306 B.n177 163.367
R1991 B.n310 B.n177 163.367
R1992 B.n311 B.n310 163.367
R1993 B.n312 B.n311 163.367
R1994 B.n312 B.n175 163.367
R1995 B.n316 B.n175 163.367
R1996 B.n317 B.n316 163.367
R1997 B.n318 B.n317 163.367
R1998 B.n318 B.n173 163.367
R1999 B.n322 B.n173 163.367
R2000 B.n323 B.n322 163.367
R2001 B.n324 B.n323 163.367
R2002 B.n324 B.n171 163.367
R2003 B.n328 B.n171 163.367
R2004 B.n329 B.n328 163.367
R2005 B.n330 B.n329 163.367
R2006 B.n330 B.n169 163.367
R2007 B.n334 B.n169 163.367
R2008 B.n335 B.n334 163.367
R2009 B.n336 B.n335 163.367
R2010 B.n336 B.n167 163.367
R2011 B.n340 B.n167 163.367
R2012 B.n341 B.n340 163.367
R2013 B.n342 B.n341 163.367
R2014 B.n342 B.n165 163.367
R2015 B.n346 B.n165 163.367
R2016 B.n347 B.n346 163.367
R2017 B.n348 B.n347 163.367
R2018 B.n348 B.n161 163.367
R2019 B.n353 B.n161 163.367
R2020 B.n354 B.n353 163.367
R2021 B.n355 B.n354 163.367
R2022 B.n355 B.n159 163.367
R2023 B.n359 B.n159 163.367
R2024 B.n360 B.n359 163.367
R2025 B.n361 B.n360 163.367
R2026 B.n361 B.n157 163.367
R2027 B.n365 B.n157 163.367
R2028 B.n366 B.n365 163.367
R2029 B.n366 B.n153 163.367
R2030 B.n370 B.n153 163.367
R2031 B.n371 B.n370 163.367
R2032 B.n372 B.n371 163.367
R2033 B.n372 B.n151 163.367
R2034 B.n376 B.n151 163.367
R2035 B.n377 B.n376 163.367
R2036 B.n378 B.n377 163.367
R2037 B.n378 B.n149 163.367
R2038 B.n382 B.n149 163.367
R2039 B.n383 B.n382 163.367
R2040 B.n384 B.n383 163.367
R2041 B.n384 B.n147 163.367
R2042 B.n388 B.n147 163.367
R2043 B.n389 B.n388 163.367
R2044 B.n390 B.n389 163.367
R2045 B.n390 B.n145 163.367
R2046 B.n394 B.n145 163.367
R2047 B.n395 B.n394 163.367
R2048 B.n396 B.n395 163.367
R2049 B.n396 B.n143 163.367
R2050 B.n400 B.n143 163.367
R2051 B.n401 B.n400 163.367
R2052 B.n402 B.n401 163.367
R2053 B.n402 B.n141 163.367
R2054 B.n406 B.n141 163.367
R2055 B.n407 B.n406 163.367
R2056 B.n408 B.n407 163.367
R2057 B.n408 B.n139 163.367
R2058 B.n412 B.n139 163.367
R2059 B.n413 B.n412 163.367
R2060 B.n414 B.n413 163.367
R2061 B.n414 B.n137 163.367
R2062 B.n418 B.n137 163.367
R2063 B.n419 B.n418 163.367
R2064 B.n420 B.n419 163.367
R2065 B.n420 B.n135 163.367
R2066 B.n424 B.n135 163.367
R2067 B.n425 B.n424 163.367
R2068 B.n426 B.n425 163.367
R2069 B.n426 B.n133 163.367
R2070 B.n430 B.n133 163.367
R2071 B.n431 B.n430 163.367
R2072 B.n432 B.n431 163.367
R2073 B.n432 B.n131 163.367
R2074 B.n436 B.n131 163.367
R2075 B.n437 B.n436 163.367
R2076 B.n438 B.n437 163.367
R2077 B.n438 B.n129 163.367
R2078 B.n442 B.n129 163.367
R2079 B.n443 B.n442 163.367
R2080 B.n444 B.n443 163.367
R2081 B.n444 B.n127 163.367
R2082 B.n448 B.n127 163.367
R2083 B.n449 B.n448 163.367
R2084 B.n450 B.n449 163.367
R2085 B.n450 B.n125 163.367
R2086 B.n454 B.n125 163.367
R2087 B.n455 B.n454 163.367
R2088 B.n456 B.n455 163.367
R2089 B.n456 B.n123 163.367
R2090 B.n461 B.n460 163.367
R2091 B.n462 B.n461 163.367
R2092 B.n462 B.n121 163.367
R2093 B.n466 B.n121 163.367
R2094 B.n467 B.n466 163.367
R2095 B.n468 B.n467 163.367
R2096 B.n468 B.n119 163.367
R2097 B.n472 B.n119 163.367
R2098 B.n473 B.n472 163.367
R2099 B.n474 B.n473 163.367
R2100 B.n474 B.n117 163.367
R2101 B.n478 B.n117 163.367
R2102 B.n479 B.n478 163.367
R2103 B.n480 B.n479 163.367
R2104 B.n480 B.n115 163.367
R2105 B.n484 B.n115 163.367
R2106 B.n485 B.n484 163.367
R2107 B.n486 B.n485 163.367
R2108 B.n486 B.n113 163.367
R2109 B.n490 B.n113 163.367
R2110 B.n491 B.n490 163.367
R2111 B.n492 B.n491 163.367
R2112 B.n492 B.n111 163.367
R2113 B.n496 B.n111 163.367
R2114 B.n497 B.n496 163.367
R2115 B.n498 B.n497 163.367
R2116 B.n498 B.n109 163.367
R2117 B.n502 B.n109 163.367
R2118 B.n503 B.n502 163.367
R2119 B.n504 B.n503 163.367
R2120 B.n504 B.n107 163.367
R2121 B.n508 B.n107 163.367
R2122 B.n509 B.n508 163.367
R2123 B.n510 B.n509 163.367
R2124 B.n510 B.n105 163.367
R2125 B.n514 B.n105 163.367
R2126 B.n515 B.n514 163.367
R2127 B.n516 B.n515 163.367
R2128 B.n516 B.n103 163.367
R2129 B.n520 B.n103 163.367
R2130 B.n521 B.n520 163.367
R2131 B.n522 B.n521 163.367
R2132 B.n522 B.n101 163.367
R2133 B.n526 B.n101 163.367
R2134 B.n527 B.n526 163.367
R2135 B.n528 B.n527 163.367
R2136 B.n528 B.n99 163.367
R2137 B.n532 B.n99 163.367
R2138 B.n533 B.n532 163.367
R2139 B.n534 B.n533 163.367
R2140 B.n534 B.n97 163.367
R2141 B.n538 B.n97 163.367
R2142 B.n539 B.n538 163.367
R2143 B.n540 B.n539 163.367
R2144 B.n540 B.n95 163.367
R2145 B.n544 B.n95 163.367
R2146 B.n545 B.n544 163.367
R2147 B.n546 B.n545 163.367
R2148 B.n546 B.n93 163.367
R2149 B.n550 B.n93 163.367
R2150 B.n551 B.n550 163.367
R2151 B.n552 B.n551 163.367
R2152 B.n552 B.n91 163.367
R2153 B.n556 B.n91 163.367
R2154 B.n557 B.n556 163.367
R2155 B.n558 B.n557 163.367
R2156 B.n760 B.n19 163.367
R2157 B.n756 B.n19 163.367
R2158 B.n756 B.n755 163.367
R2159 B.n755 B.n754 163.367
R2160 B.n754 B.n21 163.367
R2161 B.n750 B.n21 163.367
R2162 B.n750 B.n749 163.367
R2163 B.n749 B.n748 163.367
R2164 B.n748 B.n23 163.367
R2165 B.n744 B.n23 163.367
R2166 B.n744 B.n743 163.367
R2167 B.n743 B.n742 163.367
R2168 B.n742 B.n25 163.367
R2169 B.n738 B.n25 163.367
R2170 B.n738 B.n737 163.367
R2171 B.n737 B.n736 163.367
R2172 B.n736 B.n27 163.367
R2173 B.n732 B.n27 163.367
R2174 B.n732 B.n731 163.367
R2175 B.n731 B.n730 163.367
R2176 B.n730 B.n29 163.367
R2177 B.n726 B.n29 163.367
R2178 B.n726 B.n725 163.367
R2179 B.n725 B.n724 163.367
R2180 B.n724 B.n31 163.367
R2181 B.n720 B.n31 163.367
R2182 B.n720 B.n719 163.367
R2183 B.n719 B.n718 163.367
R2184 B.n718 B.n33 163.367
R2185 B.n714 B.n33 163.367
R2186 B.n714 B.n713 163.367
R2187 B.n713 B.n712 163.367
R2188 B.n712 B.n35 163.367
R2189 B.n708 B.n35 163.367
R2190 B.n708 B.n707 163.367
R2191 B.n707 B.n706 163.367
R2192 B.n706 B.n37 163.367
R2193 B.n702 B.n37 163.367
R2194 B.n702 B.n701 163.367
R2195 B.n701 B.n700 163.367
R2196 B.n700 B.n39 163.367
R2197 B.n696 B.n39 163.367
R2198 B.n696 B.n695 163.367
R2199 B.n695 B.n694 163.367
R2200 B.n694 B.n41 163.367
R2201 B.n690 B.n41 163.367
R2202 B.n690 B.n689 163.367
R2203 B.n689 B.n688 163.367
R2204 B.n688 B.n43 163.367
R2205 B.n684 B.n43 163.367
R2206 B.n684 B.n683 163.367
R2207 B.n683 B.n682 163.367
R2208 B.n682 B.n45 163.367
R2209 B.n678 B.n45 163.367
R2210 B.n678 B.n677 163.367
R2211 B.n677 B.n676 163.367
R2212 B.n676 B.n47 163.367
R2213 B.n672 B.n47 163.367
R2214 B.n672 B.n671 163.367
R2215 B.n671 B.n670 163.367
R2216 B.n670 B.n49 163.367
R2217 B.n665 B.n49 163.367
R2218 B.n665 B.n664 163.367
R2219 B.n664 B.n663 163.367
R2220 B.n663 B.n53 163.367
R2221 B.n659 B.n53 163.367
R2222 B.n659 B.n658 163.367
R2223 B.n658 B.n657 163.367
R2224 B.n657 B.n55 163.367
R2225 B.n653 B.n55 163.367
R2226 B.n653 B.n652 163.367
R2227 B.n652 B.n59 163.367
R2228 B.n648 B.n59 163.367
R2229 B.n648 B.n647 163.367
R2230 B.n647 B.n646 163.367
R2231 B.n646 B.n61 163.367
R2232 B.n642 B.n61 163.367
R2233 B.n642 B.n641 163.367
R2234 B.n641 B.n640 163.367
R2235 B.n640 B.n63 163.367
R2236 B.n636 B.n63 163.367
R2237 B.n636 B.n635 163.367
R2238 B.n635 B.n634 163.367
R2239 B.n634 B.n65 163.367
R2240 B.n630 B.n65 163.367
R2241 B.n630 B.n629 163.367
R2242 B.n629 B.n628 163.367
R2243 B.n628 B.n67 163.367
R2244 B.n624 B.n67 163.367
R2245 B.n624 B.n623 163.367
R2246 B.n623 B.n622 163.367
R2247 B.n622 B.n69 163.367
R2248 B.n618 B.n69 163.367
R2249 B.n618 B.n617 163.367
R2250 B.n617 B.n616 163.367
R2251 B.n616 B.n71 163.367
R2252 B.n612 B.n71 163.367
R2253 B.n612 B.n611 163.367
R2254 B.n611 B.n610 163.367
R2255 B.n610 B.n73 163.367
R2256 B.n606 B.n73 163.367
R2257 B.n606 B.n605 163.367
R2258 B.n605 B.n604 163.367
R2259 B.n604 B.n75 163.367
R2260 B.n600 B.n75 163.367
R2261 B.n600 B.n599 163.367
R2262 B.n599 B.n598 163.367
R2263 B.n598 B.n77 163.367
R2264 B.n594 B.n77 163.367
R2265 B.n594 B.n593 163.367
R2266 B.n593 B.n592 163.367
R2267 B.n592 B.n79 163.367
R2268 B.n588 B.n79 163.367
R2269 B.n588 B.n587 163.367
R2270 B.n587 B.n586 163.367
R2271 B.n586 B.n81 163.367
R2272 B.n582 B.n81 163.367
R2273 B.n582 B.n581 163.367
R2274 B.n581 B.n580 163.367
R2275 B.n580 B.n83 163.367
R2276 B.n576 B.n83 163.367
R2277 B.n576 B.n575 163.367
R2278 B.n575 B.n574 163.367
R2279 B.n574 B.n85 163.367
R2280 B.n570 B.n85 163.367
R2281 B.n570 B.n569 163.367
R2282 B.n569 B.n568 163.367
R2283 B.n568 B.n87 163.367
R2284 B.n564 B.n87 163.367
R2285 B.n564 B.n563 163.367
R2286 B.n563 B.n562 163.367
R2287 B.n562 B.n89 163.367
R2288 B.n156 B.n155 59.5399
R2289 B.n351 B.n163 59.5399
R2290 B.n667 B.n51 59.5399
R2291 B.n58 B.n57 59.5399
R2292 B.n759 B.n18 32.6249
R2293 B.n560 B.n559 32.6249
R2294 B.n459 B.n458 32.6249
R2295 B.n259 B.n194 32.6249
R2296 B.n155 B.n154 27.346
R2297 B.n163 B.n162 27.346
R2298 B.n51 B.n50 27.346
R2299 B.n57 B.n56 27.346
R2300 B B.n811 18.0485
R2301 B.n759 B.n758 10.6151
R2302 B.n758 B.n757 10.6151
R2303 B.n757 B.n20 10.6151
R2304 B.n753 B.n20 10.6151
R2305 B.n753 B.n752 10.6151
R2306 B.n752 B.n751 10.6151
R2307 B.n751 B.n22 10.6151
R2308 B.n747 B.n22 10.6151
R2309 B.n747 B.n746 10.6151
R2310 B.n746 B.n745 10.6151
R2311 B.n745 B.n24 10.6151
R2312 B.n741 B.n24 10.6151
R2313 B.n741 B.n740 10.6151
R2314 B.n740 B.n739 10.6151
R2315 B.n739 B.n26 10.6151
R2316 B.n735 B.n26 10.6151
R2317 B.n735 B.n734 10.6151
R2318 B.n734 B.n733 10.6151
R2319 B.n733 B.n28 10.6151
R2320 B.n729 B.n28 10.6151
R2321 B.n729 B.n728 10.6151
R2322 B.n728 B.n727 10.6151
R2323 B.n727 B.n30 10.6151
R2324 B.n723 B.n30 10.6151
R2325 B.n723 B.n722 10.6151
R2326 B.n722 B.n721 10.6151
R2327 B.n721 B.n32 10.6151
R2328 B.n717 B.n32 10.6151
R2329 B.n717 B.n716 10.6151
R2330 B.n716 B.n715 10.6151
R2331 B.n715 B.n34 10.6151
R2332 B.n711 B.n34 10.6151
R2333 B.n711 B.n710 10.6151
R2334 B.n710 B.n709 10.6151
R2335 B.n709 B.n36 10.6151
R2336 B.n705 B.n36 10.6151
R2337 B.n705 B.n704 10.6151
R2338 B.n704 B.n703 10.6151
R2339 B.n703 B.n38 10.6151
R2340 B.n699 B.n38 10.6151
R2341 B.n699 B.n698 10.6151
R2342 B.n698 B.n697 10.6151
R2343 B.n697 B.n40 10.6151
R2344 B.n693 B.n40 10.6151
R2345 B.n693 B.n692 10.6151
R2346 B.n692 B.n691 10.6151
R2347 B.n691 B.n42 10.6151
R2348 B.n687 B.n42 10.6151
R2349 B.n687 B.n686 10.6151
R2350 B.n686 B.n685 10.6151
R2351 B.n685 B.n44 10.6151
R2352 B.n681 B.n44 10.6151
R2353 B.n681 B.n680 10.6151
R2354 B.n680 B.n679 10.6151
R2355 B.n679 B.n46 10.6151
R2356 B.n675 B.n46 10.6151
R2357 B.n675 B.n674 10.6151
R2358 B.n674 B.n673 10.6151
R2359 B.n673 B.n48 10.6151
R2360 B.n669 B.n48 10.6151
R2361 B.n669 B.n668 10.6151
R2362 B.n666 B.n52 10.6151
R2363 B.n662 B.n52 10.6151
R2364 B.n662 B.n661 10.6151
R2365 B.n661 B.n660 10.6151
R2366 B.n660 B.n54 10.6151
R2367 B.n656 B.n54 10.6151
R2368 B.n656 B.n655 10.6151
R2369 B.n655 B.n654 10.6151
R2370 B.n651 B.n650 10.6151
R2371 B.n650 B.n649 10.6151
R2372 B.n649 B.n60 10.6151
R2373 B.n645 B.n60 10.6151
R2374 B.n645 B.n644 10.6151
R2375 B.n644 B.n643 10.6151
R2376 B.n643 B.n62 10.6151
R2377 B.n639 B.n62 10.6151
R2378 B.n639 B.n638 10.6151
R2379 B.n638 B.n637 10.6151
R2380 B.n637 B.n64 10.6151
R2381 B.n633 B.n64 10.6151
R2382 B.n633 B.n632 10.6151
R2383 B.n632 B.n631 10.6151
R2384 B.n631 B.n66 10.6151
R2385 B.n627 B.n66 10.6151
R2386 B.n627 B.n626 10.6151
R2387 B.n626 B.n625 10.6151
R2388 B.n625 B.n68 10.6151
R2389 B.n621 B.n68 10.6151
R2390 B.n621 B.n620 10.6151
R2391 B.n620 B.n619 10.6151
R2392 B.n619 B.n70 10.6151
R2393 B.n615 B.n70 10.6151
R2394 B.n615 B.n614 10.6151
R2395 B.n614 B.n613 10.6151
R2396 B.n613 B.n72 10.6151
R2397 B.n609 B.n72 10.6151
R2398 B.n609 B.n608 10.6151
R2399 B.n608 B.n607 10.6151
R2400 B.n607 B.n74 10.6151
R2401 B.n603 B.n74 10.6151
R2402 B.n603 B.n602 10.6151
R2403 B.n602 B.n601 10.6151
R2404 B.n601 B.n76 10.6151
R2405 B.n597 B.n76 10.6151
R2406 B.n597 B.n596 10.6151
R2407 B.n596 B.n595 10.6151
R2408 B.n595 B.n78 10.6151
R2409 B.n591 B.n78 10.6151
R2410 B.n591 B.n590 10.6151
R2411 B.n590 B.n589 10.6151
R2412 B.n589 B.n80 10.6151
R2413 B.n585 B.n80 10.6151
R2414 B.n585 B.n584 10.6151
R2415 B.n584 B.n583 10.6151
R2416 B.n583 B.n82 10.6151
R2417 B.n579 B.n82 10.6151
R2418 B.n579 B.n578 10.6151
R2419 B.n578 B.n577 10.6151
R2420 B.n577 B.n84 10.6151
R2421 B.n573 B.n84 10.6151
R2422 B.n573 B.n572 10.6151
R2423 B.n572 B.n571 10.6151
R2424 B.n571 B.n86 10.6151
R2425 B.n567 B.n86 10.6151
R2426 B.n567 B.n566 10.6151
R2427 B.n566 B.n565 10.6151
R2428 B.n565 B.n88 10.6151
R2429 B.n561 B.n88 10.6151
R2430 B.n561 B.n560 10.6151
R2431 B.n459 B.n122 10.6151
R2432 B.n463 B.n122 10.6151
R2433 B.n464 B.n463 10.6151
R2434 B.n465 B.n464 10.6151
R2435 B.n465 B.n120 10.6151
R2436 B.n469 B.n120 10.6151
R2437 B.n470 B.n469 10.6151
R2438 B.n471 B.n470 10.6151
R2439 B.n471 B.n118 10.6151
R2440 B.n475 B.n118 10.6151
R2441 B.n476 B.n475 10.6151
R2442 B.n477 B.n476 10.6151
R2443 B.n477 B.n116 10.6151
R2444 B.n481 B.n116 10.6151
R2445 B.n482 B.n481 10.6151
R2446 B.n483 B.n482 10.6151
R2447 B.n483 B.n114 10.6151
R2448 B.n487 B.n114 10.6151
R2449 B.n488 B.n487 10.6151
R2450 B.n489 B.n488 10.6151
R2451 B.n489 B.n112 10.6151
R2452 B.n493 B.n112 10.6151
R2453 B.n494 B.n493 10.6151
R2454 B.n495 B.n494 10.6151
R2455 B.n495 B.n110 10.6151
R2456 B.n499 B.n110 10.6151
R2457 B.n500 B.n499 10.6151
R2458 B.n501 B.n500 10.6151
R2459 B.n501 B.n108 10.6151
R2460 B.n505 B.n108 10.6151
R2461 B.n506 B.n505 10.6151
R2462 B.n507 B.n506 10.6151
R2463 B.n507 B.n106 10.6151
R2464 B.n511 B.n106 10.6151
R2465 B.n512 B.n511 10.6151
R2466 B.n513 B.n512 10.6151
R2467 B.n513 B.n104 10.6151
R2468 B.n517 B.n104 10.6151
R2469 B.n518 B.n517 10.6151
R2470 B.n519 B.n518 10.6151
R2471 B.n519 B.n102 10.6151
R2472 B.n523 B.n102 10.6151
R2473 B.n524 B.n523 10.6151
R2474 B.n525 B.n524 10.6151
R2475 B.n525 B.n100 10.6151
R2476 B.n529 B.n100 10.6151
R2477 B.n530 B.n529 10.6151
R2478 B.n531 B.n530 10.6151
R2479 B.n531 B.n98 10.6151
R2480 B.n535 B.n98 10.6151
R2481 B.n536 B.n535 10.6151
R2482 B.n537 B.n536 10.6151
R2483 B.n537 B.n96 10.6151
R2484 B.n541 B.n96 10.6151
R2485 B.n542 B.n541 10.6151
R2486 B.n543 B.n542 10.6151
R2487 B.n543 B.n94 10.6151
R2488 B.n547 B.n94 10.6151
R2489 B.n548 B.n547 10.6151
R2490 B.n549 B.n548 10.6151
R2491 B.n549 B.n92 10.6151
R2492 B.n553 B.n92 10.6151
R2493 B.n554 B.n553 10.6151
R2494 B.n555 B.n554 10.6151
R2495 B.n555 B.n90 10.6151
R2496 B.n559 B.n90 10.6151
R2497 B.n260 B.n259 10.6151
R2498 B.n261 B.n260 10.6151
R2499 B.n261 B.n192 10.6151
R2500 B.n265 B.n192 10.6151
R2501 B.n266 B.n265 10.6151
R2502 B.n267 B.n266 10.6151
R2503 B.n267 B.n190 10.6151
R2504 B.n271 B.n190 10.6151
R2505 B.n272 B.n271 10.6151
R2506 B.n273 B.n272 10.6151
R2507 B.n273 B.n188 10.6151
R2508 B.n277 B.n188 10.6151
R2509 B.n278 B.n277 10.6151
R2510 B.n279 B.n278 10.6151
R2511 B.n279 B.n186 10.6151
R2512 B.n283 B.n186 10.6151
R2513 B.n284 B.n283 10.6151
R2514 B.n285 B.n284 10.6151
R2515 B.n285 B.n184 10.6151
R2516 B.n289 B.n184 10.6151
R2517 B.n290 B.n289 10.6151
R2518 B.n291 B.n290 10.6151
R2519 B.n291 B.n182 10.6151
R2520 B.n295 B.n182 10.6151
R2521 B.n296 B.n295 10.6151
R2522 B.n297 B.n296 10.6151
R2523 B.n297 B.n180 10.6151
R2524 B.n301 B.n180 10.6151
R2525 B.n302 B.n301 10.6151
R2526 B.n303 B.n302 10.6151
R2527 B.n303 B.n178 10.6151
R2528 B.n307 B.n178 10.6151
R2529 B.n308 B.n307 10.6151
R2530 B.n309 B.n308 10.6151
R2531 B.n309 B.n176 10.6151
R2532 B.n313 B.n176 10.6151
R2533 B.n314 B.n313 10.6151
R2534 B.n315 B.n314 10.6151
R2535 B.n315 B.n174 10.6151
R2536 B.n319 B.n174 10.6151
R2537 B.n320 B.n319 10.6151
R2538 B.n321 B.n320 10.6151
R2539 B.n321 B.n172 10.6151
R2540 B.n325 B.n172 10.6151
R2541 B.n326 B.n325 10.6151
R2542 B.n327 B.n326 10.6151
R2543 B.n327 B.n170 10.6151
R2544 B.n331 B.n170 10.6151
R2545 B.n332 B.n331 10.6151
R2546 B.n333 B.n332 10.6151
R2547 B.n333 B.n168 10.6151
R2548 B.n337 B.n168 10.6151
R2549 B.n338 B.n337 10.6151
R2550 B.n339 B.n338 10.6151
R2551 B.n339 B.n166 10.6151
R2552 B.n343 B.n166 10.6151
R2553 B.n344 B.n343 10.6151
R2554 B.n345 B.n344 10.6151
R2555 B.n345 B.n164 10.6151
R2556 B.n349 B.n164 10.6151
R2557 B.n350 B.n349 10.6151
R2558 B.n352 B.n160 10.6151
R2559 B.n356 B.n160 10.6151
R2560 B.n357 B.n356 10.6151
R2561 B.n358 B.n357 10.6151
R2562 B.n358 B.n158 10.6151
R2563 B.n362 B.n158 10.6151
R2564 B.n363 B.n362 10.6151
R2565 B.n364 B.n363 10.6151
R2566 B.n368 B.n367 10.6151
R2567 B.n369 B.n368 10.6151
R2568 B.n369 B.n152 10.6151
R2569 B.n373 B.n152 10.6151
R2570 B.n374 B.n373 10.6151
R2571 B.n375 B.n374 10.6151
R2572 B.n375 B.n150 10.6151
R2573 B.n379 B.n150 10.6151
R2574 B.n380 B.n379 10.6151
R2575 B.n381 B.n380 10.6151
R2576 B.n381 B.n148 10.6151
R2577 B.n385 B.n148 10.6151
R2578 B.n386 B.n385 10.6151
R2579 B.n387 B.n386 10.6151
R2580 B.n387 B.n146 10.6151
R2581 B.n391 B.n146 10.6151
R2582 B.n392 B.n391 10.6151
R2583 B.n393 B.n392 10.6151
R2584 B.n393 B.n144 10.6151
R2585 B.n397 B.n144 10.6151
R2586 B.n398 B.n397 10.6151
R2587 B.n399 B.n398 10.6151
R2588 B.n399 B.n142 10.6151
R2589 B.n403 B.n142 10.6151
R2590 B.n404 B.n403 10.6151
R2591 B.n405 B.n404 10.6151
R2592 B.n405 B.n140 10.6151
R2593 B.n409 B.n140 10.6151
R2594 B.n410 B.n409 10.6151
R2595 B.n411 B.n410 10.6151
R2596 B.n411 B.n138 10.6151
R2597 B.n415 B.n138 10.6151
R2598 B.n416 B.n415 10.6151
R2599 B.n417 B.n416 10.6151
R2600 B.n417 B.n136 10.6151
R2601 B.n421 B.n136 10.6151
R2602 B.n422 B.n421 10.6151
R2603 B.n423 B.n422 10.6151
R2604 B.n423 B.n134 10.6151
R2605 B.n427 B.n134 10.6151
R2606 B.n428 B.n427 10.6151
R2607 B.n429 B.n428 10.6151
R2608 B.n429 B.n132 10.6151
R2609 B.n433 B.n132 10.6151
R2610 B.n434 B.n433 10.6151
R2611 B.n435 B.n434 10.6151
R2612 B.n435 B.n130 10.6151
R2613 B.n439 B.n130 10.6151
R2614 B.n440 B.n439 10.6151
R2615 B.n441 B.n440 10.6151
R2616 B.n441 B.n128 10.6151
R2617 B.n445 B.n128 10.6151
R2618 B.n446 B.n445 10.6151
R2619 B.n447 B.n446 10.6151
R2620 B.n447 B.n126 10.6151
R2621 B.n451 B.n126 10.6151
R2622 B.n452 B.n451 10.6151
R2623 B.n453 B.n452 10.6151
R2624 B.n453 B.n124 10.6151
R2625 B.n457 B.n124 10.6151
R2626 B.n458 B.n457 10.6151
R2627 B.n255 B.n194 10.6151
R2628 B.n255 B.n254 10.6151
R2629 B.n254 B.n253 10.6151
R2630 B.n253 B.n196 10.6151
R2631 B.n249 B.n196 10.6151
R2632 B.n249 B.n248 10.6151
R2633 B.n248 B.n247 10.6151
R2634 B.n247 B.n198 10.6151
R2635 B.n243 B.n198 10.6151
R2636 B.n243 B.n242 10.6151
R2637 B.n242 B.n241 10.6151
R2638 B.n241 B.n200 10.6151
R2639 B.n237 B.n200 10.6151
R2640 B.n237 B.n236 10.6151
R2641 B.n236 B.n235 10.6151
R2642 B.n235 B.n202 10.6151
R2643 B.n231 B.n202 10.6151
R2644 B.n231 B.n230 10.6151
R2645 B.n230 B.n229 10.6151
R2646 B.n229 B.n204 10.6151
R2647 B.n225 B.n204 10.6151
R2648 B.n225 B.n224 10.6151
R2649 B.n224 B.n223 10.6151
R2650 B.n223 B.n206 10.6151
R2651 B.n219 B.n206 10.6151
R2652 B.n219 B.n218 10.6151
R2653 B.n218 B.n217 10.6151
R2654 B.n217 B.n208 10.6151
R2655 B.n213 B.n208 10.6151
R2656 B.n213 B.n212 10.6151
R2657 B.n212 B.n211 10.6151
R2658 B.n211 B.n0 10.6151
R2659 B.n807 B.n1 10.6151
R2660 B.n807 B.n806 10.6151
R2661 B.n806 B.n805 10.6151
R2662 B.n805 B.n4 10.6151
R2663 B.n801 B.n4 10.6151
R2664 B.n801 B.n800 10.6151
R2665 B.n800 B.n799 10.6151
R2666 B.n799 B.n6 10.6151
R2667 B.n795 B.n6 10.6151
R2668 B.n795 B.n794 10.6151
R2669 B.n794 B.n793 10.6151
R2670 B.n793 B.n8 10.6151
R2671 B.n789 B.n8 10.6151
R2672 B.n789 B.n788 10.6151
R2673 B.n788 B.n787 10.6151
R2674 B.n787 B.n10 10.6151
R2675 B.n783 B.n10 10.6151
R2676 B.n783 B.n782 10.6151
R2677 B.n782 B.n781 10.6151
R2678 B.n781 B.n12 10.6151
R2679 B.n777 B.n12 10.6151
R2680 B.n777 B.n776 10.6151
R2681 B.n776 B.n775 10.6151
R2682 B.n775 B.n14 10.6151
R2683 B.n771 B.n14 10.6151
R2684 B.n771 B.n770 10.6151
R2685 B.n770 B.n769 10.6151
R2686 B.n769 B.n16 10.6151
R2687 B.n765 B.n16 10.6151
R2688 B.n765 B.n764 10.6151
R2689 B.n764 B.n763 10.6151
R2690 B.n763 B.n18 10.6151
R2691 B.n667 B.n666 6.5566
R2692 B.n654 B.n58 6.5566
R2693 B.n352 B.n351 6.5566
R2694 B.n364 B.n156 6.5566
R2695 B.n668 B.n667 4.05904
R2696 B.n651 B.n58 4.05904
R2697 B.n351 B.n350 4.05904
R2698 B.n367 B.n156 4.05904
R2699 B.n811 B.n0 2.81026
R2700 B.n811 B.n1 2.81026
C0 w_n2662_n4736# B 9.90836f
C1 VN VP 7.42269f
C2 w_n2662_n4736# VP 5.69842f
C3 B VDD1 2.37706f
C4 VN VTAIL 12.3646f
C5 VP VDD1 12.857599f
C6 B VDD2 2.43593f
C7 w_n2662_n4736# VTAIL 4.06939f
C8 VP VDD2 0.39117f
C9 VTAIL VDD1 17.124401f
C10 w_n2662_n4736# VN 5.35654f
C11 VTAIL VDD2 17.1593f
C12 VN VDD1 0.150254f
C13 w_n2662_n4736# VDD1 2.69834f
C14 VN VDD2 12.6231f
C15 w_n2662_n4736# VDD2 2.76287f
C16 B VP 1.54557f
C17 VDD1 VDD2 1.21383f
C18 VTAIL B 4.27967f
C19 VTAIL VP 12.3793f
C20 VN B 0.97905f
C21 VDD2 VSUBS 1.829646f
C22 VDD1 VSUBS 1.520869f
C23 VTAIL VSUBS 1.126457f
C24 VN VSUBS 5.8437f
C25 VP VSUBS 2.570634f
C26 B VSUBS 4.061087f
C27 w_n2662_n4736# VSUBS 0.154066p
C28 B.n0 VSUBS 0.005405f
C29 B.n1 VSUBS 0.005405f
C30 B.n2 VSUBS 0.008548f
C31 B.n3 VSUBS 0.008548f
C32 B.n4 VSUBS 0.008548f
C33 B.n5 VSUBS 0.008548f
C34 B.n6 VSUBS 0.008548f
C35 B.n7 VSUBS 0.008548f
C36 B.n8 VSUBS 0.008548f
C37 B.n9 VSUBS 0.008548f
C38 B.n10 VSUBS 0.008548f
C39 B.n11 VSUBS 0.008548f
C40 B.n12 VSUBS 0.008548f
C41 B.n13 VSUBS 0.008548f
C42 B.n14 VSUBS 0.008548f
C43 B.n15 VSUBS 0.008548f
C44 B.n16 VSUBS 0.008548f
C45 B.n17 VSUBS 0.008548f
C46 B.n18 VSUBS 0.01953f
C47 B.n19 VSUBS 0.008548f
C48 B.n20 VSUBS 0.008548f
C49 B.n21 VSUBS 0.008548f
C50 B.n22 VSUBS 0.008548f
C51 B.n23 VSUBS 0.008548f
C52 B.n24 VSUBS 0.008548f
C53 B.n25 VSUBS 0.008548f
C54 B.n26 VSUBS 0.008548f
C55 B.n27 VSUBS 0.008548f
C56 B.n28 VSUBS 0.008548f
C57 B.n29 VSUBS 0.008548f
C58 B.n30 VSUBS 0.008548f
C59 B.n31 VSUBS 0.008548f
C60 B.n32 VSUBS 0.008548f
C61 B.n33 VSUBS 0.008548f
C62 B.n34 VSUBS 0.008548f
C63 B.n35 VSUBS 0.008548f
C64 B.n36 VSUBS 0.008548f
C65 B.n37 VSUBS 0.008548f
C66 B.n38 VSUBS 0.008548f
C67 B.n39 VSUBS 0.008548f
C68 B.n40 VSUBS 0.008548f
C69 B.n41 VSUBS 0.008548f
C70 B.n42 VSUBS 0.008548f
C71 B.n43 VSUBS 0.008548f
C72 B.n44 VSUBS 0.008548f
C73 B.n45 VSUBS 0.008548f
C74 B.n46 VSUBS 0.008548f
C75 B.n47 VSUBS 0.008548f
C76 B.n48 VSUBS 0.008548f
C77 B.n49 VSUBS 0.008548f
C78 B.t8 VSUBS 0.453535f
C79 B.t7 VSUBS 0.474001f
C80 B.t6 VSUBS 1.02784f
C81 B.n50 VSUBS 0.614026f
C82 B.n51 VSUBS 0.405945f
C83 B.n52 VSUBS 0.008548f
C84 B.n53 VSUBS 0.008548f
C85 B.n54 VSUBS 0.008548f
C86 B.n55 VSUBS 0.008548f
C87 B.t11 VSUBS 0.45354f
C88 B.t10 VSUBS 0.474005f
C89 B.t9 VSUBS 1.02784f
C90 B.n56 VSUBS 0.614022f
C91 B.n57 VSUBS 0.405941f
C92 B.n58 VSUBS 0.019804f
C93 B.n59 VSUBS 0.008548f
C94 B.n60 VSUBS 0.008548f
C95 B.n61 VSUBS 0.008548f
C96 B.n62 VSUBS 0.008548f
C97 B.n63 VSUBS 0.008548f
C98 B.n64 VSUBS 0.008548f
C99 B.n65 VSUBS 0.008548f
C100 B.n66 VSUBS 0.008548f
C101 B.n67 VSUBS 0.008548f
C102 B.n68 VSUBS 0.008548f
C103 B.n69 VSUBS 0.008548f
C104 B.n70 VSUBS 0.008548f
C105 B.n71 VSUBS 0.008548f
C106 B.n72 VSUBS 0.008548f
C107 B.n73 VSUBS 0.008548f
C108 B.n74 VSUBS 0.008548f
C109 B.n75 VSUBS 0.008548f
C110 B.n76 VSUBS 0.008548f
C111 B.n77 VSUBS 0.008548f
C112 B.n78 VSUBS 0.008548f
C113 B.n79 VSUBS 0.008548f
C114 B.n80 VSUBS 0.008548f
C115 B.n81 VSUBS 0.008548f
C116 B.n82 VSUBS 0.008548f
C117 B.n83 VSUBS 0.008548f
C118 B.n84 VSUBS 0.008548f
C119 B.n85 VSUBS 0.008548f
C120 B.n86 VSUBS 0.008548f
C121 B.n87 VSUBS 0.008548f
C122 B.n88 VSUBS 0.008548f
C123 B.n89 VSUBS 0.020443f
C124 B.n90 VSUBS 0.008548f
C125 B.n91 VSUBS 0.008548f
C126 B.n92 VSUBS 0.008548f
C127 B.n93 VSUBS 0.008548f
C128 B.n94 VSUBS 0.008548f
C129 B.n95 VSUBS 0.008548f
C130 B.n96 VSUBS 0.008548f
C131 B.n97 VSUBS 0.008548f
C132 B.n98 VSUBS 0.008548f
C133 B.n99 VSUBS 0.008548f
C134 B.n100 VSUBS 0.008548f
C135 B.n101 VSUBS 0.008548f
C136 B.n102 VSUBS 0.008548f
C137 B.n103 VSUBS 0.008548f
C138 B.n104 VSUBS 0.008548f
C139 B.n105 VSUBS 0.008548f
C140 B.n106 VSUBS 0.008548f
C141 B.n107 VSUBS 0.008548f
C142 B.n108 VSUBS 0.008548f
C143 B.n109 VSUBS 0.008548f
C144 B.n110 VSUBS 0.008548f
C145 B.n111 VSUBS 0.008548f
C146 B.n112 VSUBS 0.008548f
C147 B.n113 VSUBS 0.008548f
C148 B.n114 VSUBS 0.008548f
C149 B.n115 VSUBS 0.008548f
C150 B.n116 VSUBS 0.008548f
C151 B.n117 VSUBS 0.008548f
C152 B.n118 VSUBS 0.008548f
C153 B.n119 VSUBS 0.008548f
C154 B.n120 VSUBS 0.008548f
C155 B.n121 VSUBS 0.008548f
C156 B.n122 VSUBS 0.008548f
C157 B.n123 VSUBS 0.020443f
C158 B.n124 VSUBS 0.008548f
C159 B.n125 VSUBS 0.008548f
C160 B.n126 VSUBS 0.008548f
C161 B.n127 VSUBS 0.008548f
C162 B.n128 VSUBS 0.008548f
C163 B.n129 VSUBS 0.008548f
C164 B.n130 VSUBS 0.008548f
C165 B.n131 VSUBS 0.008548f
C166 B.n132 VSUBS 0.008548f
C167 B.n133 VSUBS 0.008548f
C168 B.n134 VSUBS 0.008548f
C169 B.n135 VSUBS 0.008548f
C170 B.n136 VSUBS 0.008548f
C171 B.n137 VSUBS 0.008548f
C172 B.n138 VSUBS 0.008548f
C173 B.n139 VSUBS 0.008548f
C174 B.n140 VSUBS 0.008548f
C175 B.n141 VSUBS 0.008548f
C176 B.n142 VSUBS 0.008548f
C177 B.n143 VSUBS 0.008548f
C178 B.n144 VSUBS 0.008548f
C179 B.n145 VSUBS 0.008548f
C180 B.n146 VSUBS 0.008548f
C181 B.n147 VSUBS 0.008548f
C182 B.n148 VSUBS 0.008548f
C183 B.n149 VSUBS 0.008548f
C184 B.n150 VSUBS 0.008548f
C185 B.n151 VSUBS 0.008548f
C186 B.n152 VSUBS 0.008548f
C187 B.n153 VSUBS 0.008548f
C188 B.t1 VSUBS 0.45354f
C189 B.t2 VSUBS 0.474005f
C190 B.t0 VSUBS 1.02784f
C191 B.n154 VSUBS 0.614022f
C192 B.n155 VSUBS 0.405941f
C193 B.n156 VSUBS 0.019804f
C194 B.n157 VSUBS 0.008548f
C195 B.n158 VSUBS 0.008548f
C196 B.n159 VSUBS 0.008548f
C197 B.n160 VSUBS 0.008548f
C198 B.n161 VSUBS 0.008548f
C199 B.t4 VSUBS 0.453535f
C200 B.t5 VSUBS 0.474001f
C201 B.t3 VSUBS 1.02784f
C202 B.n162 VSUBS 0.614026f
C203 B.n163 VSUBS 0.405945f
C204 B.n164 VSUBS 0.008548f
C205 B.n165 VSUBS 0.008548f
C206 B.n166 VSUBS 0.008548f
C207 B.n167 VSUBS 0.008548f
C208 B.n168 VSUBS 0.008548f
C209 B.n169 VSUBS 0.008548f
C210 B.n170 VSUBS 0.008548f
C211 B.n171 VSUBS 0.008548f
C212 B.n172 VSUBS 0.008548f
C213 B.n173 VSUBS 0.008548f
C214 B.n174 VSUBS 0.008548f
C215 B.n175 VSUBS 0.008548f
C216 B.n176 VSUBS 0.008548f
C217 B.n177 VSUBS 0.008548f
C218 B.n178 VSUBS 0.008548f
C219 B.n179 VSUBS 0.008548f
C220 B.n180 VSUBS 0.008548f
C221 B.n181 VSUBS 0.008548f
C222 B.n182 VSUBS 0.008548f
C223 B.n183 VSUBS 0.008548f
C224 B.n184 VSUBS 0.008548f
C225 B.n185 VSUBS 0.008548f
C226 B.n186 VSUBS 0.008548f
C227 B.n187 VSUBS 0.008548f
C228 B.n188 VSUBS 0.008548f
C229 B.n189 VSUBS 0.008548f
C230 B.n190 VSUBS 0.008548f
C231 B.n191 VSUBS 0.008548f
C232 B.n192 VSUBS 0.008548f
C233 B.n193 VSUBS 0.008548f
C234 B.n194 VSUBS 0.01953f
C235 B.n195 VSUBS 0.008548f
C236 B.n196 VSUBS 0.008548f
C237 B.n197 VSUBS 0.008548f
C238 B.n198 VSUBS 0.008548f
C239 B.n199 VSUBS 0.008548f
C240 B.n200 VSUBS 0.008548f
C241 B.n201 VSUBS 0.008548f
C242 B.n202 VSUBS 0.008548f
C243 B.n203 VSUBS 0.008548f
C244 B.n204 VSUBS 0.008548f
C245 B.n205 VSUBS 0.008548f
C246 B.n206 VSUBS 0.008548f
C247 B.n207 VSUBS 0.008548f
C248 B.n208 VSUBS 0.008548f
C249 B.n209 VSUBS 0.008548f
C250 B.n210 VSUBS 0.008548f
C251 B.n211 VSUBS 0.008548f
C252 B.n212 VSUBS 0.008548f
C253 B.n213 VSUBS 0.008548f
C254 B.n214 VSUBS 0.008548f
C255 B.n215 VSUBS 0.008548f
C256 B.n216 VSUBS 0.008548f
C257 B.n217 VSUBS 0.008548f
C258 B.n218 VSUBS 0.008548f
C259 B.n219 VSUBS 0.008548f
C260 B.n220 VSUBS 0.008548f
C261 B.n221 VSUBS 0.008548f
C262 B.n222 VSUBS 0.008548f
C263 B.n223 VSUBS 0.008548f
C264 B.n224 VSUBS 0.008548f
C265 B.n225 VSUBS 0.008548f
C266 B.n226 VSUBS 0.008548f
C267 B.n227 VSUBS 0.008548f
C268 B.n228 VSUBS 0.008548f
C269 B.n229 VSUBS 0.008548f
C270 B.n230 VSUBS 0.008548f
C271 B.n231 VSUBS 0.008548f
C272 B.n232 VSUBS 0.008548f
C273 B.n233 VSUBS 0.008548f
C274 B.n234 VSUBS 0.008548f
C275 B.n235 VSUBS 0.008548f
C276 B.n236 VSUBS 0.008548f
C277 B.n237 VSUBS 0.008548f
C278 B.n238 VSUBS 0.008548f
C279 B.n239 VSUBS 0.008548f
C280 B.n240 VSUBS 0.008548f
C281 B.n241 VSUBS 0.008548f
C282 B.n242 VSUBS 0.008548f
C283 B.n243 VSUBS 0.008548f
C284 B.n244 VSUBS 0.008548f
C285 B.n245 VSUBS 0.008548f
C286 B.n246 VSUBS 0.008548f
C287 B.n247 VSUBS 0.008548f
C288 B.n248 VSUBS 0.008548f
C289 B.n249 VSUBS 0.008548f
C290 B.n250 VSUBS 0.008548f
C291 B.n251 VSUBS 0.008548f
C292 B.n252 VSUBS 0.008548f
C293 B.n253 VSUBS 0.008548f
C294 B.n254 VSUBS 0.008548f
C295 B.n255 VSUBS 0.008548f
C296 B.n256 VSUBS 0.008548f
C297 B.n257 VSUBS 0.01953f
C298 B.n258 VSUBS 0.020443f
C299 B.n259 VSUBS 0.020443f
C300 B.n260 VSUBS 0.008548f
C301 B.n261 VSUBS 0.008548f
C302 B.n262 VSUBS 0.008548f
C303 B.n263 VSUBS 0.008548f
C304 B.n264 VSUBS 0.008548f
C305 B.n265 VSUBS 0.008548f
C306 B.n266 VSUBS 0.008548f
C307 B.n267 VSUBS 0.008548f
C308 B.n268 VSUBS 0.008548f
C309 B.n269 VSUBS 0.008548f
C310 B.n270 VSUBS 0.008548f
C311 B.n271 VSUBS 0.008548f
C312 B.n272 VSUBS 0.008548f
C313 B.n273 VSUBS 0.008548f
C314 B.n274 VSUBS 0.008548f
C315 B.n275 VSUBS 0.008548f
C316 B.n276 VSUBS 0.008548f
C317 B.n277 VSUBS 0.008548f
C318 B.n278 VSUBS 0.008548f
C319 B.n279 VSUBS 0.008548f
C320 B.n280 VSUBS 0.008548f
C321 B.n281 VSUBS 0.008548f
C322 B.n282 VSUBS 0.008548f
C323 B.n283 VSUBS 0.008548f
C324 B.n284 VSUBS 0.008548f
C325 B.n285 VSUBS 0.008548f
C326 B.n286 VSUBS 0.008548f
C327 B.n287 VSUBS 0.008548f
C328 B.n288 VSUBS 0.008548f
C329 B.n289 VSUBS 0.008548f
C330 B.n290 VSUBS 0.008548f
C331 B.n291 VSUBS 0.008548f
C332 B.n292 VSUBS 0.008548f
C333 B.n293 VSUBS 0.008548f
C334 B.n294 VSUBS 0.008548f
C335 B.n295 VSUBS 0.008548f
C336 B.n296 VSUBS 0.008548f
C337 B.n297 VSUBS 0.008548f
C338 B.n298 VSUBS 0.008548f
C339 B.n299 VSUBS 0.008548f
C340 B.n300 VSUBS 0.008548f
C341 B.n301 VSUBS 0.008548f
C342 B.n302 VSUBS 0.008548f
C343 B.n303 VSUBS 0.008548f
C344 B.n304 VSUBS 0.008548f
C345 B.n305 VSUBS 0.008548f
C346 B.n306 VSUBS 0.008548f
C347 B.n307 VSUBS 0.008548f
C348 B.n308 VSUBS 0.008548f
C349 B.n309 VSUBS 0.008548f
C350 B.n310 VSUBS 0.008548f
C351 B.n311 VSUBS 0.008548f
C352 B.n312 VSUBS 0.008548f
C353 B.n313 VSUBS 0.008548f
C354 B.n314 VSUBS 0.008548f
C355 B.n315 VSUBS 0.008548f
C356 B.n316 VSUBS 0.008548f
C357 B.n317 VSUBS 0.008548f
C358 B.n318 VSUBS 0.008548f
C359 B.n319 VSUBS 0.008548f
C360 B.n320 VSUBS 0.008548f
C361 B.n321 VSUBS 0.008548f
C362 B.n322 VSUBS 0.008548f
C363 B.n323 VSUBS 0.008548f
C364 B.n324 VSUBS 0.008548f
C365 B.n325 VSUBS 0.008548f
C366 B.n326 VSUBS 0.008548f
C367 B.n327 VSUBS 0.008548f
C368 B.n328 VSUBS 0.008548f
C369 B.n329 VSUBS 0.008548f
C370 B.n330 VSUBS 0.008548f
C371 B.n331 VSUBS 0.008548f
C372 B.n332 VSUBS 0.008548f
C373 B.n333 VSUBS 0.008548f
C374 B.n334 VSUBS 0.008548f
C375 B.n335 VSUBS 0.008548f
C376 B.n336 VSUBS 0.008548f
C377 B.n337 VSUBS 0.008548f
C378 B.n338 VSUBS 0.008548f
C379 B.n339 VSUBS 0.008548f
C380 B.n340 VSUBS 0.008548f
C381 B.n341 VSUBS 0.008548f
C382 B.n342 VSUBS 0.008548f
C383 B.n343 VSUBS 0.008548f
C384 B.n344 VSUBS 0.008548f
C385 B.n345 VSUBS 0.008548f
C386 B.n346 VSUBS 0.008548f
C387 B.n347 VSUBS 0.008548f
C388 B.n348 VSUBS 0.008548f
C389 B.n349 VSUBS 0.008548f
C390 B.n350 VSUBS 0.005908f
C391 B.n351 VSUBS 0.019804f
C392 B.n352 VSUBS 0.006914f
C393 B.n353 VSUBS 0.008548f
C394 B.n354 VSUBS 0.008548f
C395 B.n355 VSUBS 0.008548f
C396 B.n356 VSUBS 0.008548f
C397 B.n357 VSUBS 0.008548f
C398 B.n358 VSUBS 0.008548f
C399 B.n359 VSUBS 0.008548f
C400 B.n360 VSUBS 0.008548f
C401 B.n361 VSUBS 0.008548f
C402 B.n362 VSUBS 0.008548f
C403 B.n363 VSUBS 0.008548f
C404 B.n364 VSUBS 0.006914f
C405 B.n365 VSUBS 0.008548f
C406 B.n366 VSUBS 0.008548f
C407 B.n367 VSUBS 0.005908f
C408 B.n368 VSUBS 0.008548f
C409 B.n369 VSUBS 0.008548f
C410 B.n370 VSUBS 0.008548f
C411 B.n371 VSUBS 0.008548f
C412 B.n372 VSUBS 0.008548f
C413 B.n373 VSUBS 0.008548f
C414 B.n374 VSUBS 0.008548f
C415 B.n375 VSUBS 0.008548f
C416 B.n376 VSUBS 0.008548f
C417 B.n377 VSUBS 0.008548f
C418 B.n378 VSUBS 0.008548f
C419 B.n379 VSUBS 0.008548f
C420 B.n380 VSUBS 0.008548f
C421 B.n381 VSUBS 0.008548f
C422 B.n382 VSUBS 0.008548f
C423 B.n383 VSUBS 0.008548f
C424 B.n384 VSUBS 0.008548f
C425 B.n385 VSUBS 0.008548f
C426 B.n386 VSUBS 0.008548f
C427 B.n387 VSUBS 0.008548f
C428 B.n388 VSUBS 0.008548f
C429 B.n389 VSUBS 0.008548f
C430 B.n390 VSUBS 0.008548f
C431 B.n391 VSUBS 0.008548f
C432 B.n392 VSUBS 0.008548f
C433 B.n393 VSUBS 0.008548f
C434 B.n394 VSUBS 0.008548f
C435 B.n395 VSUBS 0.008548f
C436 B.n396 VSUBS 0.008548f
C437 B.n397 VSUBS 0.008548f
C438 B.n398 VSUBS 0.008548f
C439 B.n399 VSUBS 0.008548f
C440 B.n400 VSUBS 0.008548f
C441 B.n401 VSUBS 0.008548f
C442 B.n402 VSUBS 0.008548f
C443 B.n403 VSUBS 0.008548f
C444 B.n404 VSUBS 0.008548f
C445 B.n405 VSUBS 0.008548f
C446 B.n406 VSUBS 0.008548f
C447 B.n407 VSUBS 0.008548f
C448 B.n408 VSUBS 0.008548f
C449 B.n409 VSUBS 0.008548f
C450 B.n410 VSUBS 0.008548f
C451 B.n411 VSUBS 0.008548f
C452 B.n412 VSUBS 0.008548f
C453 B.n413 VSUBS 0.008548f
C454 B.n414 VSUBS 0.008548f
C455 B.n415 VSUBS 0.008548f
C456 B.n416 VSUBS 0.008548f
C457 B.n417 VSUBS 0.008548f
C458 B.n418 VSUBS 0.008548f
C459 B.n419 VSUBS 0.008548f
C460 B.n420 VSUBS 0.008548f
C461 B.n421 VSUBS 0.008548f
C462 B.n422 VSUBS 0.008548f
C463 B.n423 VSUBS 0.008548f
C464 B.n424 VSUBS 0.008548f
C465 B.n425 VSUBS 0.008548f
C466 B.n426 VSUBS 0.008548f
C467 B.n427 VSUBS 0.008548f
C468 B.n428 VSUBS 0.008548f
C469 B.n429 VSUBS 0.008548f
C470 B.n430 VSUBS 0.008548f
C471 B.n431 VSUBS 0.008548f
C472 B.n432 VSUBS 0.008548f
C473 B.n433 VSUBS 0.008548f
C474 B.n434 VSUBS 0.008548f
C475 B.n435 VSUBS 0.008548f
C476 B.n436 VSUBS 0.008548f
C477 B.n437 VSUBS 0.008548f
C478 B.n438 VSUBS 0.008548f
C479 B.n439 VSUBS 0.008548f
C480 B.n440 VSUBS 0.008548f
C481 B.n441 VSUBS 0.008548f
C482 B.n442 VSUBS 0.008548f
C483 B.n443 VSUBS 0.008548f
C484 B.n444 VSUBS 0.008548f
C485 B.n445 VSUBS 0.008548f
C486 B.n446 VSUBS 0.008548f
C487 B.n447 VSUBS 0.008548f
C488 B.n448 VSUBS 0.008548f
C489 B.n449 VSUBS 0.008548f
C490 B.n450 VSUBS 0.008548f
C491 B.n451 VSUBS 0.008548f
C492 B.n452 VSUBS 0.008548f
C493 B.n453 VSUBS 0.008548f
C494 B.n454 VSUBS 0.008548f
C495 B.n455 VSUBS 0.008548f
C496 B.n456 VSUBS 0.008548f
C497 B.n457 VSUBS 0.008548f
C498 B.n458 VSUBS 0.020443f
C499 B.n459 VSUBS 0.01953f
C500 B.n460 VSUBS 0.01953f
C501 B.n461 VSUBS 0.008548f
C502 B.n462 VSUBS 0.008548f
C503 B.n463 VSUBS 0.008548f
C504 B.n464 VSUBS 0.008548f
C505 B.n465 VSUBS 0.008548f
C506 B.n466 VSUBS 0.008548f
C507 B.n467 VSUBS 0.008548f
C508 B.n468 VSUBS 0.008548f
C509 B.n469 VSUBS 0.008548f
C510 B.n470 VSUBS 0.008548f
C511 B.n471 VSUBS 0.008548f
C512 B.n472 VSUBS 0.008548f
C513 B.n473 VSUBS 0.008548f
C514 B.n474 VSUBS 0.008548f
C515 B.n475 VSUBS 0.008548f
C516 B.n476 VSUBS 0.008548f
C517 B.n477 VSUBS 0.008548f
C518 B.n478 VSUBS 0.008548f
C519 B.n479 VSUBS 0.008548f
C520 B.n480 VSUBS 0.008548f
C521 B.n481 VSUBS 0.008548f
C522 B.n482 VSUBS 0.008548f
C523 B.n483 VSUBS 0.008548f
C524 B.n484 VSUBS 0.008548f
C525 B.n485 VSUBS 0.008548f
C526 B.n486 VSUBS 0.008548f
C527 B.n487 VSUBS 0.008548f
C528 B.n488 VSUBS 0.008548f
C529 B.n489 VSUBS 0.008548f
C530 B.n490 VSUBS 0.008548f
C531 B.n491 VSUBS 0.008548f
C532 B.n492 VSUBS 0.008548f
C533 B.n493 VSUBS 0.008548f
C534 B.n494 VSUBS 0.008548f
C535 B.n495 VSUBS 0.008548f
C536 B.n496 VSUBS 0.008548f
C537 B.n497 VSUBS 0.008548f
C538 B.n498 VSUBS 0.008548f
C539 B.n499 VSUBS 0.008548f
C540 B.n500 VSUBS 0.008548f
C541 B.n501 VSUBS 0.008548f
C542 B.n502 VSUBS 0.008548f
C543 B.n503 VSUBS 0.008548f
C544 B.n504 VSUBS 0.008548f
C545 B.n505 VSUBS 0.008548f
C546 B.n506 VSUBS 0.008548f
C547 B.n507 VSUBS 0.008548f
C548 B.n508 VSUBS 0.008548f
C549 B.n509 VSUBS 0.008548f
C550 B.n510 VSUBS 0.008548f
C551 B.n511 VSUBS 0.008548f
C552 B.n512 VSUBS 0.008548f
C553 B.n513 VSUBS 0.008548f
C554 B.n514 VSUBS 0.008548f
C555 B.n515 VSUBS 0.008548f
C556 B.n516 VSUBS 0.008548f
C557 B.n517 VSUBS 0.008548f
C558 B.n518 VSUBS 0.008548f
C559 B.n519 VSUBS 0.008548f
C560 B.n520 VSUBS 0.008548f
C561 B.n521 VSUBS 0.008548f
C562 B.n522 VSUBS 0.008548f
C563 B.n523 VSUBS 0.008548f
C564 B.n524 VSUBS 0.008548f
C565 B.n525 VSUBS 0.008548f
C566 B.n526 VSUBS 0.008548f
C567 B.n527 VSUBS 0.008548f
C568 B.n528 VSUBS 0.008548f
C569 B.n529 VSUBS 0.008548f
C570 B.n530 VSUBS 0.008548f
C571 B.n531 VSUBS 0.008548f
C572 B.n532 VSUBS 0.008548f
C573 B.n533 VSUBS 0.008548f
C574 B.n534 VSUBS 0.008548f
C575 B.n535 VSUBS 0.008548f
C576 B.n536 VSUBS 0.008548f
C577 B.n537 VSUBS 0.008548f
C578 B.n538 VSUBS 0.008548f
C579 B.n539 VSUBS 0.008548f
C580 B.n540 VSUBS 0.008548f
C581 B.n541 VSUBS 0.008548f
C582 B.n542 VSUBS 0.008548f
C583 B.n543 VSUBS 0.008548f
C584 B.n544 VSUBS 0.008548f
C585 B.n545 VSUBS 0.008548f
C586 B.n546 VSUBS 0.008548f
C587 B.n547 VSUBS 0.008548f
C588 B.n548 VSUBS 0.008548f
C589 B.n549 VSUBS 0.008548f
C590 B.n550 VSUBS 0.008548f
C591 B.n551 VSUBS 0.008548f
C592 B.n552 VSUBS 0.008548f
C593 B.n553 VSUBS 0.008548f
C594 B.n554 VSUBS 0.008548f
C595 B.n555 VSUBS 0.008548f
C596 B.n556 VSUBS 0.008548f
C597 B.n557 VSUBS 0.008548f
C598 B.n558 VSUBS 0.01953f
C599 B.n559 VSUBS 0.020541f
C600 B.n560 VSUBS 0.019432f
C601 B.n561 VSUBS 0.008548f
C602 B.n562 VSUBS 0.008548f
C603 B.n563 VSUBS 0.008548f
C604 B.n564 VSUBS 0.008548f
C605 B.n565 VSUBS 0.008548f
C606 B.n566 VSUBS 0.008548f
C607 B.n567 VSUBS 0.008548f
C608 B.n568 VSUBS 0.008548f
C609 B.n569 VSUBS 0.008548f
C610 B.n570 VSUBS 0.008548f
C611 B.n571 VSUBS 0.008548f
C612 B.n572 VSUBS 0.008548f
C613 B.n573 VSUBS 0.008548f
C614 B.n574 VSUBS 0.008548f
C615 B.n575 VSUBS 0.008548f
C616 B.n576 VSUBS 0.008548f
C617 B.n577 VSUBS 0.008548f
C618 B.n578 VSUBS 0.008548f
C619 B.n579 VSUBS 0.008548f
C620 B.n580 VSUBS 0.008548f
C621 B.n581 VSUBS 0.008548f
C622 B.n582 VSUBS 0.008548f
C623 B.n583 VSUBS 0.008548f
C624 B.n584 VSUBS 0.008548f
C625 B.n585 VSUBS 0.008548f
C626 B.n586 VSUBS 0.008548f
C627 B.n587 VSUBS 0.008548f
C628 B.n588 VSUBS 0.008548f
C629 B.n589 VSUBS 0.008548f
C630 B.n590 VSUBS 0.008548f
C631 B.n591 VSUBS 0.008548f
C632 B.n592 VSUBS 0.008548f
C633 B.n593 VSUBS 0.008548f
C634 B.n594 VSUBS 0.008548f
C635 B.n595 VSUBS 0.008548f
C636 B.n596 VSUBS 0.008548f
C637 B.n597 VSUBS 0.008548f
C638 B.n598 VSUBS 0.008548f
C639 B.n599 VSUBS 0.008548f
C640 B.n600 VSUBS 0.008548f
C641 B.n601 VSUBS 0.008548f
C642 B.n602 VSUBS 0.008548f
C643 B.n603 VSUBS 0.008548f
C644 B.n604 VSUBS 0.008548f
C645 B.n605 VSUBS 0.008548f
C646 B.n606 VSUBS 0.008548f
C647 B.n607 VSUBS 0.008548f
C648 B.n608 VSUBS 0.008548f
C649 B.n609 VSUBS 0.008548f
C650 B.n610 VSUBS 0.008548f
C651 B.n611 VSUBS 0.008548f
C652 B.n612 VSUBS 0.008548f
C653 B.n613 VSUBS 0.008548f
C654 B.n614 VSUBS 0.008548f
C655 B.n615 VSUBS 0.008548f
C656 B.n616 VSUBS 0.008548f
C657 B.n617 VSUBS 0.008548f
C658 B.n618 VSUBS 0.008548f
C659 B.n619 VSUBS 0.008548f
C660 B.n620 VSUBS 0.008548f
C661 B.n621 VSUBS 0.008548f
C662 B.n622 VSUBS 0.008548f
C663 B.n623 VSUBS 0.008548f
C664 B.n624 VSUBS 0.008548f
C665 B.n625 VSUBS 0.008548f
C666 B.n626 VSUBS 0.008548f
C667 B.n627 VSUBS 0.008548f
C668 B.n628 VSUBS 0.008548f
C669 B.n629 VSUBS 0.008548f
C670 B.n630 VSUBS 0.008548f
C671 B.n631 VSUBS 0.008548f
C672 B.n632 VSUBS 0.008548f
C673 B.n633 VSUBS 0.008548f
C674 B.n634 VSUBS 0.008548f
C675 B.n635 VSUBS 0.008548f
C676 B.n636 VSUBS 0.008548f
C677 B.n637 VSUBS 0.008548f
C678 B.n638 VSUBS 0.008548f
C679 B.n639 VSUBS 0.008548f
C680 B.n640 VSUBS 0.008548f
C681 B.n641 VSUBS 0.008548f
C682 B.n642 VSUBS 0.008548f
C683 B.n643 VSUBS 0.008548f
C684 B.n644 VSUBS 0.008548f
C685 B.n645 VSUBS 0.008548f
C686 B.n646 VSUBS 0.008548f
C687 B.n647 VSUBS 0.008548f
C688 B.n648 VSUBS 0.008548f
C689 B.n649 VSUBS 0.008548f
C690 B.n650 VSUBS 0.008548f
C691 B.n651 VSUBS 0.005908f
C692 B.n652 VSUBS 0.008548f
C693 B.n653 VSUBS 0.008548f
C694 B.n654 VSUBS 0.006914f
C695 B.n655 VSUBS 0.008548f
C696 B.n656 VSUBS 0.008548f
C697 B.n657 VSUBS 0.008548f
C698 B.n658 VSUBS 0.008548f
C699 B.n659 VSUBS 0.008548f
C700 B.n660 VSUBS 0.008548f
C701 B.n661 VSUBS 0.008548f
C702 B.n662 VSUBS 0.008548f
C703 B.n663 VSUBS 0.008548f
C704 B.n664 VSUBS 0.008548f
C705 B.n665 VSUBS 0.008548f
C706 B.n666 VSUBS 0.006914f
C707 B.n667 VSUBS 0.019804f
C708 B.n668 VSUBS 0.005908f
C709 B.n669 VSUBS 0.008548f
C710 B.n670 VSUBS 0.008548f
C711 B.n671 VSUBS 0.008548f
C712 B.n672 VSUBS 0.008548f
C713 B.n673 VSUBS 0.008548f
C714 B.n674 VSUBS 0.008548f
C715 B.n675 VSUBS 0.008548f
C716 B.n676 VSUBS 0.008548f
C717 B.n677 VSUBS 0.008548f
C718 B.n678 VSUBS 0.008548f
C719 B.n679 VSUBS 0.008548f
C720 B.n680 VSUBS 0.008548f
C721 B.n681 VSUBS 0.008548f
C722 B.n682 VSUBS 0.008548f
C723 B.n683 VSUBS 0.008548f
C724 B.n684 VSUBS 0.008548f
C725 B.n685 VSUBS 0.008548f
C726 B.n686 VSUBS 0.008548f
C727 B.n687 VSUBS 0.008548f
C728 B.n688 VSUBS 0.008548f
C729 B.n689 VSUBS 0.008548f
C730 B.n690 VSUBS 0.008548f
C731 B.n691 VSUBS 0.008548f
C732 B.n692 VSUBS 0.008548f
C733 B.n693 VSUBS 0.008548f
C734 B.n694 VSUBS 0.008548f
C735 B.n695 VSUBS 0.008548f
C736 B.n696 VSUBS 0.008548f
C737 B.n697 VSUBS 0.008548f
C738 B.n698 VSUBS 0.008548f
C739 B.n699 VSUBS 0.008548f
C740 B.n700 VSUBS 0.008548f
C741 B.n701 VSUBS 0.008548f
C742 B.n702 VSUBS 0.008548f
C743 B.n703 VSUBS 0.008548f
C744 B.n704 VSUBS 0.008548f
C745 B.n705 VSUBS 0.008548f
C746 B.n706 VSUBS 0.008548f
C747 B.n707 VSUBS 0.008548f
C748 B.n708 VSUBS 0.008548f
C749 B.n709 VSUBS 0.008548f
C750 B.n710 VSUBS 0.008548f
C751 B.n711 VSUBS 0.008548f
C752 B.n712 VSUBS 0.008548f
C753 B.n713 VSUBS 0.008548f
C754 B.n714 VSUBS 0.008548f
C755 B.n715 VSUBS 0.008548f
C756 B.n716 VSUBS 0.008548f
C757 B.n717 VSUBS 0.008548f
C758 B.n718 VSUBS 0.008548f
C759 B.n719 VSUBS 0.008548f
C760 B.n720 VSUBS 0.008548f
C761 B.n721 VSUBS 0.008548f
C762 B.n722 VSUBS 0.008548f
C763 B.n723 VSUBS 0.008548f
C764 B.n724 VSUBS 0.008548f
C765 B.n725 VSUBS 0.008548f
C766 B.n726 VSUBS 0.008548f
C767 B.n727 VSUBS 0.008548f
C768 B.n728 VSUBS 0.008548f
C769 B.n729 VSUBS 0.008548f
C770 B.n730 VSUBS 0.008548f
C771 B.n731 VSUBS 0.008548f
C772 B.n732 VSUBS 0.008548f
C773 B.n733 VSUBS 0.008548f
C774 B.n734 VSUBS 0.008548f
C775 B.n735 VSUBS 0.008548f
C776 B.n736 VSUBS 0.008548f
C777 B.n737 VSUBS 0.008548f
C778 B.n738 VSUBS 0.008548f
C779 B.n739 VSUBS 0.008548f
C780 B.n740 VSUBS 0.008548f
C781 B.n741 VSUBS 0.008548f
C782 B.n742 VSUBS 0.008548f
C783 B.n743 VSUBS 0.008548f
C784 B.n744 VSUBS 0.008548f
C785 B.n745 VSUBS 0.008548f
C786 B.n746 VSUBS 0.008548f
C787 B.n747 VSUBS 0.008548f
C788 B.n748 VSUBS 0.008548f
C789 B.n749 VSUBS 0.008548f
C790 B.n750 VSUBS 0.008548f
C791 B.n751 VSUBS 0.008548f
C792 B.n752 VSUBS 0.008548f
C793 B.n753 VSUBS 0.008548f
C794 B.n754 VSUBS 0.008548f
C795 B.n755 VSUBS 0.008548f
C796 B.n756 VSUBS 0.008548f
C797 B.n757 VSUBS 0.008548f
C798 B.n758 VSUBS 0.008548f
C799 B.n759 VSUBS 0.020443f
C800 B.n760 VSUBS 0.020443f
C801 B.n761 VSUBS 0.01953f
C802 B.n762 VSUBS 0.008548f
C803 B.n763 VSUBS 0.008548f
C804 B.n764 VSUBS 0.008548f
C805 B.n765 VSUBS 0.008548f
C806 B.n766 VSUBS 0.008548f
C807 B.n767 VSUBS 0.008548f
C808 B.n768 VSUBS 0.008548f
C809 B.n769 VSUBS 0.008548f
C810 B.n770 VSUBS 0.008548f
C811 B.n771 VSUBS 0.008548f
C812 B.n772 VSUBS 0.008548f
C813 B.n773 VSUBS 0.008548f
C814 B.n774 VSUBS 0.008548f
C815 B.n775 VSUBS 0.008548f
C816 B.n776 VSUBS 0.008548f
C817 B.n777 VSUBS 0.008548f
C818 B.n778 VSUBS 0.008548f
C819 B.n779 VSUBS 0.008548f
C820 B.n780 VSUBS 0.008548f
C821 B.n781 VSUBS 0.008548f
C822 B.n782 VSUBS 0.008548f
C823 B.n783 VSUBS 0.008548f
C824 B.n784 VSUBS 0.008548f
C825 B.n785 VSUBS 0.008548f
C826 B.n786 VSUBS 0.008548f
C827 B.n787 VSUBS 0.008548f
C828 B.n788 VSUBS 0.008548f
C829 B.n789 VSUBS 0.008548f
C830 B.n790 VSUBS 0.008548f
C831 B.n791 VSUBS 0.008548f
C832 B.n792 VSUBS 0.008548f
C833 B.n793 VSUBS 0.008548f
C834 B.n794 VSUBS 0.008548f
C835 B.n795 VSUBS 0.008548f
C836 B.n796 VSUBS 0.008548f
C837 B.n797 VSUBS 0.008548f
C838 B.n798 VSUBS 0.008548f
C839 B.n799 VSUBS 0.008548f
C840 B.n800 VSUBS 0.008548f
C841 B.n801 VSUBS 0.008548f
C842 B.n802 VSUBS 0.008548f
C843 B.n803 VSUBS 0.008548f
C844 B.n804 VSUBS 0.008548f
C845 B.n805 VSUBS 0.008548f
C846 B.n806 VSUBS 0.008548f
C847 B.n807 VSUBS 0.008548f
C848 B.n808 VSUBS 0.008548f
C849 B.n809 VSUBS 0.008548f
C850 B.n810 VSUBS 0.008548f
C851 B.n811 VSUBS 0.019355f
C852 VDD2.n0 VSUBS 0.028657f
C853 VDD2.n1 VSUBS 0.027017f
C854 VDD2.n2 VSUBS 0.014518f
C855 VDD2.n3 VSUBS 0.034315f
C856 VDD2.n4 VSUBS 0.015372f
C857 VDD2.n5 VSUBS 0.027017f
C858 VDD2.n6 VSUBS 0.014518f
C859 VDD2.n7 VSUBS 0.034315f
C860 VDD2.n8 VSUBS 0.015372f
C861 VDD2.n9 VSUBS 0.027017f
C862 VDD2.n10 VSUBS 0.014518f
C863 VDD2.n11 VSUBS 0.034315f
C864 VDD2.n12 VSUBS 0.015372f
C865 VDD2.n13 VSUBS 0.027017f
C866 VDD2.n14 VSUBS 0.014518f
C867 VDD2.n15 VSUBS 0.034315f
C868 VDD2.n16 VSUBS 0.015372f
C869 VDD2.n17 VSUBS 0.027017f
C870 VDD2.n18 VSUBS 0.014518f
C871 VDD2.n19 VSUBS 0.034315f
C872 VDD2.n20 VSUBS 0.015372f
C873 VDD2.n21 VSUBS 0.027017f
C874 VDD2.n22 VSUBS 0.014518f
C875 VDD2.n23 VSUBS 0.034315f
C876 VDD2.n24 VSUBS 0.015372f
C877 VDD2.n25 VSUBS 0.027017f
C878 VDD2.n26 VSUBS 0.014518f
C879 VDD2.n27 VSUBS 0.034315f
C880 VDD2.n28 VSUBS 0.015372f
C881 VDD2.n29 VSUBS 0.027017f
C882 VDD2.n30 VSUBS 0.014518f
C883 VDD2.n31 VSUBS 0.034315f
C884 VDD2.n32 VSUBS 0.015372f
C885 VDD2.n33 VSUBS 0.22105f
C886 VDD2.t0 VSUBS 0.07372f
C887 VDD2.n34 VSUBS 0.025736f
C888 VDD2.n35 VSUBS 0.02183f
C889 VDD2.n36 VSUBS 0.014518f
C890 VDD2.n37 VSUBS 2.19609f
C891 VDD2.n38 VSUBS 0.027017f
C892 VDD2.n39 VSUBS 0.014518f
C893 VDD2.n40 VSUBS 0.015372f
C894 VDD2.n41 VSUBS 0.034315f
C895 VDD2.n42 VSUBS 0.034315f
C896 VDD2.n43 VSUBS 0.015372f
C897 VDD2.n44 VSUBS 0.014518f
C898 VDD2.n45 VSUBS 0.027017f
C899 VDD2.n46 VSUBS 0.027017f
C900 VDD2.n47 VSUBS 0.014518f
C901 VDD2.n48 VSUBS 0.015372f
C902 VDD2.n49 VSUBS 0.034315f
C903 VDD2.n50 VSUBS 0.034315f
C904 VDD2.n51 VSUBS 0.015372f
C905 VDD2.n52 VSUBS 0.014518f
C906 VDD2.n53 VSUBS 0.027017f
C907 VDD2.n54 VSUBS 0.027017f
C908 VDD2.n55 VSUBS 0.014518f
C909 VDD2.n56 VSUBS 0.015372f
C910 VDD2.n57 VSUBS 0.034315f
C911 VDD2.n58 VSUBS 0.034315f
C912 VDD2.n59 VSUBS 0.015372f
C913 VDD2.n60 VSUBS 0.014518f
C914 VDD2.n61 VSUBS 0.027017f
C915 VDD2.n62 VSUBS 0.027017f
C916 VDD2.n63 VSUBS 0.014518f
C917 VDD2.n64 VSUBS 0.015372f
C918 VDD2.n65 VSUBS 0.034315f
C919 VDD2.n66 VSUBS 0.034315f
C920 VDD2.n67 VSUBS 0.015372f
C921 VDD2.n68 VSUBS 0.014518f
C922 VDD2.n69 VSUBS 0.027017f
C923 VDD2.n70 VSUBS 0.027017f
C924 VDD2.n71 VSUBS 0.014518f
C925 VDD2.n72 VSUBS 0.015372f
C926 VDD2.n73 VSUBS 0.034315f
C927 VDD2.n74 VSUBS 0.034315f
C928 VDD2.n75 VSUBS 0.034315f
C929 VDD2.n76 VSUBS 0.015372f
C930 VDD2.n77 VSUBS 0.014518f
C931 VDD2.n78 VSUBS 0.027017f
C932 VDD2.n79 VSUBS 0.027017f
C933 VDD2.n80 VSUBS 0.014518f
C934 VDD2.n81 VSUBS 0.014945f
C935 VDD2.n82 VSUBS 0.014945f
C936 VDD2.n83 VSUBS 0.034315f
C937 VDD2.n84 VSUBS 0.034315f
C938 VDD2.n85 VSUBS 0.015372f
C939 VDD2.n86 VSUBS 0.014518f
C940 VDD2.n87 VSUBS 0.027017f
C941 VDD2.n88 VSUBS 0.027017f
C942 VDD2.n89 VSUBS 0.014518f
C943 VDD2.n90 VSUBS 0.015372f
C944 VDD2.n91 VSUBS 0.034315f
C945 VDD2.n92 VSUBS 0.034315f
C946 VDD2.n93 VSUBS 0.015372f
C947 VDD2.n94 VSUBS 0.014518f
C948 VDD2.n95 VSUBS 0.027017f
C949 VDD2.n96 VSUBS 0.027017f
C950 VDD2.n97 VSUBS 0.014518f
C951 VDD2.n98 VSUBS 0.015372f
C952 VDD2.n99 VSUBS 0.034315f
C953 VDD2.n100 VSUBS 0.079568f
C954 VDD2.n101 VSUBS 0.015372f
C955 VDD2.n102 VSUBS 0.014518f
C956 VDD2.n103 VSUBS 0.05802f
C957 VDD2.n104 VSUBS 0.062364f
C958 VDD2.t5 VSUBS 0.402232f
C959 VDD2.t1 VSUBS 0.402232f
C960 VDD2.n105 VSUBS 3.34635f
C961 VDD2.n106 VSUBS 0.831029f
C962 VDD2.t7 VSUBS 0.402232f
C963 VDD2.t2 VSUBS 0.402232f
C964 VDD2.n107 VSUBS 3.35584f
C965 VDD2.n108 VSUBS 3.05841f
C966 VDD2.n109 VSUBS 0.028657f
C967 VDD2.n110 VSUBS 0.027017f
C968 VDD2.n111 VSUBS 0.014518f
C969 VDD2.n112 VSUBS 0.034315f
C970 VDD2.n113 VSUBS 0.015372f
C971 VDD2.n114 VSUBS 0.027017f
C972 VDD2.n115 VSUBS 0.014518f
C973 VDD2.n116 VSUBS 0.034315f
C974 VDD2.n117 VSUBS 0.015372f
C975 VDD2.n118 VSUBS 0.027017f
C976 VDD2.n119 VSUBS 0.014518f
C977 VDD2.n120 VSUBS 0.034315f
C978 VDD2.n121 VSUBS 0.015372f
C979 VDD2.n122 VSUBS 0.027017f
C980 VDD2.n123 VSUBS 0.014518f
C981 VDD2.n124 VSUBS 0.034315f
C982 VDD2.n125 VSUBS 0.034315f
C983 VDD2.n126 VSUBS 0.015372f
C984 VDD2.n127 VSUBS 0.027017f
C985 VDD2.n128 VSUBS 0.014518f
C986 VDD2.n129 VSUBS 0.034315f
C987 VDD2.n130 VSUBS 0.015372f
C988 VDD2.n131 VSUBS 0.027017f
C989 VDD2.n132 VSUBS 0.014518f
C990 VDD2.n133 VSUBS 0.034315f
C991 VDD2.n134 VSUBS 0.015372f
C992 VDD2.n135 VSUBS 0.027017f
C993 VDD2.n136 VSUBS 0.014518f
C994 VDD2.n137 VSUBS 0.034315f
C995 VDD2.n138 VSUBS 0.015372f
C996 VDD2.n139 VSUBS 0.027017f
C997 VDD2.n140 VSUBS 0.014518f
C998 VDD2.n141 VSUBS 0.034315f
C999 VDD2.n142 VSUBS 0.015372f
C1000 VDD2.n143 VSUBS 0.22105f
C1001 VDD2.t8 VSUBS 0.07372f
C1002 VDD2.n144 VSUBS 0.025736f
C1003 VDD2.n145 VSUBS 0.02183f
C1004 VDD2.n146 VSUBS 0.014518f
C1005 VDD2.n147 VSUBS 2.19609f
C1006 VDD2.n148 VSUBS 0.027017f
C1007 VDD2.n149 VSUBS 0.014518f
C1008 VDD2.n150 VSUBS 0.015372f
C1009 VDD2.n151 VSUBS 0.034315f
C1010 VDD2.n152 VSUBS 0.034315f
C1011 VDD2.n153 VSUBS 0.015372f
C1012 VDD2.n154 VSUBS 0.014518f
C1013 VDD2.n155 VSUBS 0.027017f
C1014 VDD2.n156 VSUBS 0.027017f
C1015 VDD2.n157 VSUBS 0.014518f
C1016 VDD2.n158 VSUBS 0.015372f
C1017 VDD2.n159 VSUBS 0.034315f
C1018 VDD2.n160 VSUBS 0.034315f
C1019 VDD2.n161 VSUBS 0.015372f
C1020 VDD2.n162 VSUBS 0.014518f
C1021 VDD2.n163 VSUBS 0.027017f
C1022 VDD2.n164 VSUBS 0.027017f
C1023 VDD2.n165 VSUBS 0.014518f
C1024 VDD2.n166 VSUBS 0.015372f
C1025 VDD2.n167 VSUBS 0.034315f
C1026 VDD2.n168 VSUBS 0.034315f
C1027 VDD2.n169 VSUBS 0.015372f
C1028 VDD2.n170 VSUBS 0.014518f
C1029 VDD2.n171 VSUBS 0.027017f
C1030 VDD2.n172 VSUBS 0.027017f
C1031 VDD2.n173 VSUBS 0.014518f
C1032 VDD2.n174 VSUBS 0.015372f
C1033 VDD2.n175 VSUBS 0.034315f
C1034 VDD2.n176 VSUBS 0.034315f
C1035 VDD2.n177 VSUBS 0.015372f
C1036 VDD2.n178 VSUBS 0.014518f
C1037 VDD2.n179 VSUBS 0.027017f
C1038 VDD2.n180 VSUBS 0.027017f
C1039 VDD2.n181 VSUBS 0.014518f
C1040 VDD2.n182 VSUBS 0.015372f
C1041 VDD2.n183 VSUBS 0.034315f
C1042 VDD2.n184 VSUBS 0.034315f
C1043 VDD2.n185 VSUBS 0.015372f
C1044 VDD2.n186 VSUBS 0.014518f
C1045 VDD2.n187 VSUBS 0.027017f
C1046 VDD2.n188 VSUBS 0.027017f
C1047 VDD2.n189 VSUBS 0.014518f
C1048 VDD2.n190 VSUBS 0.014945f
C1049 VDD2.n191 VSUBS 0.014945f
C1050 VDD2.n192 VSUBS 0.034315f
C1051 VDD2.n193 VSUBS 0.034315f
C1052 VDD2.n194 VSUBS 0.015372f
C1053 VDD2.n195 VSUBS 0.014518f
C1054 VDD2.n196 VSUBS 0.027017f
C1055 VDD2.n197 VSUBS 0.027017f
C1056 VDD2.n198 VSUBS 0.014518f
C1057 VDD2.n199 VSUBS 0.015372f
C1058 VDD2.n200 VSUBS 0.034315f
C1059 VDD2.n201 VSUBS 0.034315f
C1060 VDD2.n202 VSUBS 0.015372f
C1061 VDD2.n203 VSUBS 0.014518f
C1062 VDD2.n204 VSUBS 0.027017f
C1063 VDD2.n205 VSUBS 0.027017f
C1064 VDD2.n206 VSUBS 0.014518f
C1065 VDD2.n207 VSUBS 0.015372f
C1066 VDD2.n208 VSUBS 0.034315f
C1067 VDD2.n209 VSUBS 0.079568f
C1068 VDD2.n210 VSUBS 0.015372f
C1069 VDD2.n211 VSUBS 0.014518f
C1070 VDD2.n212 VSUBS 0.05802f
C1071 VDD2.n213 VSUBS 0.058411f
C1072 VDD2.n214 VSUBS 3.05143f
C1073 VDD2.t9 VSUBS 0.402232f
C1074 VDD2.t6 VSUBS 0.402232f
C1075 VDD2.n215 VSUBS 3.34636f
C1076 VDD2.n216 VSUBS 0.687029f
C1077 VDD2.t3 VSUBS 0.402232f
C1078 VDD2.t4 VSUBS 0.402232f
C1079 VDD2.n217 VSUBS 3.35579f
C1080 VN.n0 VSUBS 0.054319f
C1081 VN.t2 VSUBS 2.28018f
C1082 VN.n1 VSUBS 0.811018f
C1083 VN.n2 VSUBS 0.040708f
C1084 VN.t8 VSUBS 2.28018f
C1085 VN.n3 VSUBS 0.054107f
C1086 VN.t9 VSUBS 2.38618f
C1087 VN.n4 VSUBS 0.867132f
C1088 VN.t4 VSUBS 2.28018f
C1089 VN.n5 VSUBS 0.868685f
C1090 VN.n6 VSUBS 0.057535f
C1091 VN.n7 VSUBS 0.207182f
C1092 VN.n8 VSUBS 0.040708f
C1093 VN.n9 VSUBS 0.040708f
C1094 VN.n10 VSUBS 0.84924f
C1095 VN.n11 VSUBS 0.054107f
C1096 VN.n12 VSUBS 0.057535f
C1097 VN.n13 VSUBS 0.040708f
C1098 VN.n14 VSUBS 0.040708f
C1099 VN.n15 VSUBS 0.049836f
C1100 VN.n16 VSUBS 0.0354f
C1101 VN.t7 VSUBS 2.34713f
C1102 VN.n17 VSUBS 0.876738f
C1103 VN.n18 VSUBS 0.038124f
C1104 VN.n19 VSUBS 0.054319f
C1105 VN.t0 VSUBS 2.28018f
C1106 VN.n20 VSUBS 0.811018f
C1107 VN.n21 VSUBS 0.040708f
C1108 VN.t3 VSUBS 2.28018f
C1109 VN.n22 VSUBS 0.054107f
C1110 VN.t5 VSUBS 2.38618f
C1111 VN.n23 VSUBS 0.867132f
C1112 VN.t6 VSUBS 2.28018f
C1113 VN.n24 VSUBS 0.868685f
C1114 VN.n25 VSUBS 0.057535f
C1115 VN.n26 VSUBS 0.207182f
C1116 VN.n27 VSUBS 0.040708f
C1117 VN.n28 VSUBS 0.040708f
C1118 VN.n29 VSUBS 0.84924f
C1119 VN.n30 VSUBS 0.054107f
C1120 VN.n31 VSUBS 0.057535f
C1121 VN.n32 VSUBS 0.040708f
C1122 VN.n33 VSUBS 0.040708f
C1123 VN.n34 VSUBS 0.049836f
C1124 VN.n35 VSUBS 0.0354f
C1125 VN.t1 VSUBS 2.34713f
C1126 VN.n36 VSUBS 0.876738f
C1127 VN.n37 VSUBS 2.2587f
C1128 VDD1.n0 VSUBS 0.028657f
C1129 VDD1.n1 VSUBS 0.027018f
C1130 VDD1.n2 VSUBS 0.014518f
C1131 VDD1.n3 VSUBS 0.034315f
C1132 VDD1.n4 VSUBS 0.015372f
C1133 VDD1.n5 VSUBS 0.027018f
C1134 VDD1.n6 VSUBS 0.014518f
C1135 VDD1.n7 VSUBS 0.034315f
C1136 VDD1.n8 VSUBS 0.015372f
C1137 VDD1.n9 VSUBS 0.027018f
C1138 VDD1.n10 VSUBS 0.014518f
C1139 VDD1.n11 VSUBS 0.034315f
C1140 VDD1.n12 VSUBS 0.015372f
C1141 VDD1.n13 VSUBS 0.027018f
C1142 VDD1.n14 VSUBS 0.014518f
C1143 VDD1.n15 VSUBS 0.034315f
C1144 VDD1.n16 VSUBS 0.034315f
C1145 VDD1.n17 VSUBS 0.015372f
C1146 VDD1.n18 VSUBS 0.027018f
C1147 VDD1.n19 VSUBS 0.014518f
C1148 VDD1.n20 VSUBS 0.034315f
C1149 VDD1.n21 VSUBS 0.015372f
C1150 VDD1.n22 VSUBS 0.027018f
C1151 VDD1.n23 VSUBS 0.014518f
C1152 VDD1.n24 VSUBS 0.034315f
C1153 VDD1.n25 VSUBS 0.015372f
C1154 VDD1.n26 VSUBS 0.027018f
C1155 VDD1.n27 VSUBS 0.014518f
C1156 VDD1.n28 VSUBS 0.034315f
C1157 VDD1.n29 VSUBS 0.015372f
C1158 VDD1.n30 VSUBS 0.027018f
C1159 VDD1.n31 VSUBS 0.014518f
C1160 VDD1.n32 VSUBS 0.034315f
C1161 VDD1.n33 VSUBS 0.015372f
C1162 VDD1.n34 VSUBS 0.221051f
C1163 VDD1.t2 VSUBS 0.07372f
C1164 VDD1.n35 VSUBS 0.025737f
C1165 VDD1.n36 VSUBS 0.02183f
C1166 VDD1.n37 VSUBS 0.014518f
C1167 VDD1.n38 VSUBS 2.1961f
C1168 VDD1.n39 VSUBS 0.027018f
C1169 VDD1.n40 VSUBS 0.014518f
C1170 VDD1.n41 VSUBS 0.015372f
C1171 VDD1.n42 VSUBS 0.034315f
C1172 VDD1.n43 VSUBS 0.034315f
C1173 VDD1.n44 VSUBS 0.015372f
C1174 VDD1.n45 VSUBS 0.014518f
C1175 VDD1.n46 VSUBS 0.027018f
C1176 VDD1.n47 VSUBS 0.027018f
C1177 VDD1.n48 VSUBS 0.014518f
C1178 VDD1.n49 VSUBS 0.015372f
C1179 VDD1.n50 VSUBS 0.034315f
C1180 VDD1.n51 VSUBS 0.034315f
C1181 VDD1.n52 VSUBS 0.015372f
C1182 VDD1.n53 VSUBS 0.014518f
C1183 VDD1.n54 VSUBS 0.027018f
C1184 VDD1.n55 VSUBS 0.027018f
C1185 VDD1.n56 VSUBS 0.014518f
C1186 VDD1.n57 VSUBS 0.015372f
C1187 VDD1.n58 VSUBS 0.034315f
C1188 VDD1.n59 VSUBS 0.034315f
C1189 VDD1.n60 VSUBS 0.015372f
C1190 VDD1.n61 VSUBS 0.014518f
C1191 VDD1.n62 VSUBS 0.027018f
C1192 VDD1.n63 VSUBS 0.027018f
C1193 VDD1.n64 VSUBS 0.014518f
C1194 VDD1.n65 VSUBS 0.015372f
C1195 VDD1.n66 VSUBS 0.034315f
C1196 VDD1.n67 VSUBS 0.034315f
C1197 VDD1.n68 VSUBS 0.015372f
C1198 VDD1.n69 VSUBS 0.014518f
C1199 VDD1.n70 VSUBS 0.027018f
C1200 VDD1.n71 VSUBS 0.027018f
C1201 VDD1.n72 VSUBS 0.014518f
C1202 VDD1.n73 VSUBS 0.015372f
C1203 VDD1.n74 VSUBS 0.034315f
C1204 VDD1.n75 VSUBS 0.034315f
C1205 VDD1.n76 VSUBS 0.015372f
C1206 VDD1.n77 VSUBS 0.014518f
C1207 VDD1.n78 VSUBS 0.027018f
C1208 VDD1.n79 VSUBS 0.027018f
C1209 VDD1.n80 VSUBS 0.014518f
C1210 VDD1.n81 VSUBS 0.014945f
C1211 VDD1.n82 VSUBS 0.014945f
C1212 VDD1.n83 VSUBS 0.034315f
C1213 VDD1.n84 VSUBS 0.034315f
C1214 VDD1.n85 VSUBS 0.015372f
C1215 VDD1.n86 VSUBS 0.014518f
C1216 VDD1.n87 VSUBS 0.027018f
C1217 VDD1.n88 VSUBS 0.027018f
C1218 VDD1.n89 VSUBS 0.014518f
C1219 VDD1.n90 VSUBS 0.015372f
C1220 VDD1.n91 VSUBS 0.034315f
C1221 VDD1.n92 VSUBS 0.034315f
C1222 VDD1.n93 VSUBS 0.015372f
C1223 VDD1.n94 VSUBS 0.014518f
C1224 VDD1.n95 VSUBS 0.027018f
C1225 VDD1.n96 VSUBS 0.027018f
C1226 VDD1.n97 VSUBS 0.014518f
C1227 VDD1.n98 VSUBS 0.015372f
C1228 VDD1.n99 VSUBS 0.034315f
C1229 VDD1.n100 VSUBS 0.079568f
C1230 VDD1.n101 VSUBS 0.015372f
C1231 VDD1.n102 VSUBS 0.014518f
C1232 VDD1.n103 VSUBS 0.058021f
C1233 VDD1.n104 VSUBS 0.062364f
C1234 VDD1.t3 VSUBS 0.402235f
C1235 VDD1.t4 VSUBS 0.402235f
C1236 VDD1.n105 VSUBS 3.34638f
C1237 VDD1.n106 VSUBS 0.838388f
C1238 VDD1.n107 VSUBS 0.028657f
C1239 VDD1.n108 VSUBS 0.027018f
C1240 VDD1.n109 VSUBS 0.014518f
C1241 VDD1.n110 VSUBS 0.034315f
C1242 VDD1.n111 VSUBS 0.015372f
C1243 VDD1.n112 VSUBS 0.027018f
C1244 VDD1.n113 VSUBS 0.014518f
C1245 VDD1.n114 VSUBS 0.034315f
C1246 VDD1.n115 VSUBS 0.015372f
C1247 VDD1.n116 VSUBS 0.027018f
C1248 VDD1.n117 VSUBS 0.014518f
C1249 VDD1.n118 VSUBS 0.034315f
C1250 VDD1.n119 VSUBS 0.015372f
C1251 VDD1.n120 VSUBS 0.027018f
C1252 VDD1.n121 VSUBS 0.014518f
C1253 VDD1.n122 VSUBS 0.034315f
C1254 VDD1.n123 VSUBS 0.015372f
C1255 VDD1.n124 VSUBS 0.027018f
C1256 VDD1.n125 VSUBS 0.014518f
C1257 VDD1.n126 VSUBS 0.034315f
C1258 VDD1.n127 VSUBS 0.015372f
C1259 VDD1.n128 VSUBS 0.027018f
C1260 VDD1.n129 VSUBS 0.014518f
C1261 VDD1.n130 VSUBS 0.034315f
C1262 VDD1.n131 VSUBS 0.015372f
C1263 VDD1.n132 VSUBS 0.027018f
C1264 VDD1.n133 VSUBS 0.014518f
C1265 VDD1.n134 VSUBS 0.034315f
C1266 VDD1.n135 VSUBS 0.015372f
C1267 VDD1.n136 VSUBS 0.027018f
C1268 VDD1.n137 VSUBS 0.014518f
C1269 VDD1.n138 VSUBS 0.034315f
C1270 VDD1.n139 VSUBS 0.015372f
C1271 VDD1.n140 VSUBS 0.221051f
C1272 VDD1.t5 VSUBS 0.07372f
C1273 VDD1.n141 VSUBS 0.025737f
C1274 VDD1.n142 VSUBS 0.02183f
C1275 VDD1.n143 VSUBS 0.014518f
C1276 VDD1.n144 VSUBS 2.19611f
C1277 VDD1.n145 VSUBS 0.027018f
C1278 VDD1.n146 VSUBS 0.014518f
C1279 VDD1.n147 VSUBS 0.015372f
C1280 VDD1.n148 VSUBS 0.034315f
C1281 VDD1.n149 VSUBS 0.034315f
C1282 VDD1.n150 VSUBS 0.015372f
C1283 VDD1.n151 VSUBS 0.014518f
C1284 VDD1.n152 VSUBS 0.027018f
C1285 VDD1.n153 VSUBS 0.027018f
C1286 VDD1.n154 VSUBS 0.014518f
C1287 VDD1.n155 VSUBS 0.015372f
C1288 VDD1.n156 VSUBS 0.034315f
C1289 VDD1.n157 VSUBS 0.034315f
C1290 VDD1.n158 VSUBS 0.015372f
C1291 VDD1.n159 VSUBS 0.014518f
C1292 VDD1.n160 VSUBS 0.027018f
C1293 VDD1.n161 VSUBS 0.027018f
C1294 VDD1.n162 VSUBS 0.014518f
C1295 VDD1.n163 VSUBS 0.015372f
C1296 VDD1.n164 VSUBS 0.034315f
C1297 VDD1.n165 VSUBS 0.034315f
C1298 VDD1.n166 VSUBS 0.015372f
C1299 VDD1.n167 VSUBS 0.014518f
C1300 VDD1.n168 VSUBS 0.027018f
C1301 VDD1.n169 VSUBS 0.027018f
C1302 VDD1.n170 VSUBS 0.014518f
C1303 VDD1.n171 VSUBS 0.015372f
C1304 VDD1.n172 VSUBS 0.034315f
C1305 VDD1.n173 VSUBS 0.034315f
C1306 VDD1.n174 VSUBS 0.015372f
C1307 VDD1.n175 VSUBS 0.014518f
C1308 VDD1.n176 VSUBS 0.027018f
C1309 VDD1.n177 VSUBS 0.027018f
C1310 VDD1.n178 VSUBS 0.014518f
C1311 VDD1.n179 VSUBS 0.015372f
C1312 VDD1.n180 VSUBS 0.034315f
C1313 VDD1.n181 VSUBS 0.034315f
C1314 VDD1.n182 VSUBS 0.034315f
C1315 VDD1.n183 VSUBS 0.015372f
C1316 VDD1.n184 VSUBS 0.014518f
C1317 VDD1.n185 VSUBS 0.027018f
C1318 VDD1.n186 VSUBS 0.027018f
C1319 VDD1.n187 VSUBS 0.014518f
C1320 VDD1.n188 VSUBS 0.014945f
C1321 VDD1.n189 VSUBS 0.014945f
C1322 VDD1.n190 VSUBS 0.034315f
C1323 VDD1.n191 VSUBS 0.034315f
C1324 VDD1.n192 VSUBS 0.015372f
C1325 VDD1.n193 VSUBS 0.014518f
C1326 VDD1.n194 VSUBS 0.027018f
C1327 VDD1.n195 VSUBS 0.027018f
C1328 VDD1.n196 VSUBS 0.014518f
C1329 VDD1.n197 VSUBS 0.015372f
C1330 VDD1.n198 VSUBS 0.034315f
C1331 VDD1.n199 VSUBS 0.034315f
C1332 VDD1.n200 VSUBS 0.015372f
C1333 VDD1.n201 VSUBS 0.014518f
C1334 VDD1.n202 VSUBS 0.027018f
C1335 VDD1.n203 VSUBS 0.027018f
C1336 VDD1.n204 VSUBS 0.014518f
C1337 VDD1.n205 VSUBS 0.015372f
C1338 VDD1.n206 VSUBS 0.034315f
C1339 VDD1.n207 VSUBS 0.079568f
C1340 VDD1.n208 VSUBS 0.015372f
C1341 VDD1.n209 VSUBS 0.014518f
C1342 VDD1.n210 VSUBS 0.058021f
C1343 VDD1.n211 VSUBS 0.062364f
C1344 VDD1.t8 VSUBS 0.402235f
C1345 VDD1.t0 VSUBS 0.402235f
C1346 VDD1.n212 VSUBS 3.34637f
C1347 VDD1.n213 VSUBS 0.831034f
C1348 VDD1.t7 VSUBS 0.402235f
C1349 VDD1.t1 VSUBS 0.402235f
C1350 VDD1.n214 VSUBS 3.35586f
C1351 VDD1.n215 VSUBS 3.15393f
C1352 VDD1.t6 VSUBS 0.402235f
C1353 VDD1.t9 VSUBS 0.402235f
C1354 VDD1.n216 VSUBS 3.34636f
C1355 VDD1.n217 VSUBS 3.64114f
C1356 VTAIL.t6 VSUBS 0.405461f
C1357 VTAIL.t1 VSUBS 0.405461f
C1358 VTAIL.n0 VSUBS 3.1878f
C1359 VTAIL.n1 VSUBS 0.882179f
C1360 VTAIL.n2 VSUBS 0.028887f
C1361 VTAIL.n3 VSUBS 0.027234f
C1362 VTAIL.n4 VSUBS 0.014634f
C1363 VTAIL.n5 VSUBS 0.034591f
C1364 VTAIL.n6 VSUBS 0.015495f
C1365 VTAIL.n7 VSUBS 0.027234f
C1366 VTAIL.n8 VSUBS 0.014634f
C1367 VTAIL.n9 VSUBS 0.034591f
C1368 VTAIL.n10 VSUBS 0.015495f
C1369 VTAIL.n11 VSUBS 0.027234f
C1370 VTAIL.n12 VSUBS 0.014634f
C1371 VTAIL.n13 VSUBS 0.034591f
C1372 VTAIL.n14 VSUBS 0.015495f
C1373 VTAIL.n15 VSUBS 0.027234f
C1374 VTAIL.n16 VSUBS 0.014634f
C1375 VTAIL.n17 VSUBS 0.034591f
C1376 VTAIL.n18 VSUBS 0.015495f
C1377 VTAIL.n19 VSUBS 0.027234f
C1378 VTAIL.n20 VSUBS 0.014634f
C1379 VTAIL.n21 VSUBS 0.034591f
C1380 VTAIL.n22 VSUBS 0.015495f
C1381 VTAIL.n23 VSUBS 0.027234f
C1382 VTAIL.n24 VSUBS 0.014634f
C1383 VTAIL.n25 VSUBS 0.034591f
C1384 VTAIL.n26 VSUBS 0.015495f
C1385 VTAIL.n27 VSUBS 0.027234f
C1386 VTAIL.n28 VSUBS 0.014634f
C1387 VTAIL.n29 VSUBS 0.034591f
C1388 VTAIL.n30 VSUBS 0.015495f
C1389 VTAIL.n31 VSUBS 0.027234f
C1390 VTAIL.n32 VSUBS 0.014634f
C1391 VTAIL.n33 VSUBS 0.034591f
C1392 VTAIL.n34 VSUBS 0.015495f
C1393 VTAIL.n35 VSUBS 0.222824f
C1394 VTAIL.t14 VSUBS 0.074312f
C1395 VTAIL.n36 VSUBS 0.025943f
C1396 VTAIL.n37 VSUBS 0.022005f
C1397 VTAIL.n38 VSUBS 0.014634f
C1398 VTAIL.n39 VSUBS 2.21372f
C1399 VTAIL.n40 VSUBS 0.027234f
C1400 VTAIL.n41 VSUBS 0.014634f
C1401 VTAIL.n42 VSUBS 0.015495f
C1402 VTAIL.n43 VSUBS 0.034591f
C1403 VTAIL.n44 VSUBS 0.034591f
C1404 VTAIL.n45 VSUBS 0.015495f
C1405 VTAIL.n46 VSUBS 0.014634f
C1406 VTAIL.n47 VSUBS 0.027234f
C1407 VTAIL.n48 VSUBS 0.027234f
C1408 VTAIL.n49 VSUBS 0.014634f
C1409 VTAIL.n50 VSUBS 0.015495f
C1410 VTAIL.n51 VSUBS 0.034591f
C1411 VTAIL.n52 VSUBS 0.034591f
C1412 VTAIL.n53 VSUBS 0.015495f
C1413 VTAIL.n54 VSUBS 0.014634f
C1414 VTAIL.n55 VSUBS 0.027234f
C1415 VTAIL.n56 VSUBS 0.027234f
C1416 VTAIL.n57 VSUBS 0.014634f
C1417 VTAIL.n58 VSUBS 0.015495f
C1418 VTAIL.n59 VSUBS 0.034591f
C1419 VTAIL.n60 VSUBS 0.034591f
C1420 VTAIL.n61 VSUBS 0.015495f
C1421 VTAIL.n62 VSUBS 0.014634f
C1422 VTAIL.n63 VSUBS 0.027234f
C1423 VTAIL.n64 VSUBS 0.027234f
C1424 VTAIL.n65 VSUBS 0.014634f
C1425 VTAIL.n66 VSUBS 0.015495f
C1426 VTAIL.n67 VSUBS 0.034591f
C1427 VTAIL.n68 VSUBS 0.034591f
C1428 VTAIL.n69 VSUBS 0.015495f
C1429 VTAIL.n70 VSUBS 0.014634f
C1430 VTAIL.n71 VSUBS 0.027234f
C1431 VTAIL.n72 VSUBS 0.027234f
C1432 VTAIL.n73 VSUBS 0.014634f
C1433 VTAIL.n74 VSUBS 0.015495f
C1434 VTAIL.n75 VSUBS 0.034591f
C1435 VTAIL.n76 VSUBS 0.034591f
C1436 VTAIL.n77 VSUBS 0.034591f
C1437 VTAIL.n78 VSUBS 0.015495f
C1438 VTAIL.n79 VSUBS 0.014634f
C1439 VTAIL.n80 VSUBS 0.027234f
C1440 VTAIL.n81 VSUBS 0.027234f
C1441 VTAIL.n82 VSUBS 0.014634f
C1442 VTAIL.n83 VSUBS 0.015065f
C1443 VTAIL.n84 VSUBS 0.015065f
C1444 VTAIL.n85 VSUBS 0.034591f
C1445 VTAIL.n86 VSUBS 0.034591f
C1446 VTAIL.n87 VSUBS 0.015495f
C1447 VTAIL.n88 VSUBS 0.014634f
C1448 VTAIL.n89 VSUBS 0.027234f
C1449 VTAIL.n90 VSUBS 0.027234f
C1450 VTAIL.n91 VSUBS 0.014634f
C1451 VTAIL.n92 VSUBS 0.015495f
C1452 VTAIL.n93 VSUBS 0.034591f
C1453 VTAIL.n94 VSUBS 0.034591f
C1454 VTAIL.n95 VSUBS 0.015495f
C1455 VTAIL.n96 VSUBS 0.014634f
C1456 VTAIL.n97 VSUBS 0.027234f
C1457 VTAIL.n98 VSUBS 0.027234f
C1458 VTAIL.n99 VSUBS 0.014634f
C1459 VTAIL.n100 VSUBS 0.015495f
C1460 VTAIL.n101 VSUBS 0.034591f
C1461 VTAIL.n102 VSUBS 0.080206f
C1462 VTAIL.n103 VSUBS 0.015495f
C1463 VTAIL.n104 VSUBS 0.014634f
C1464 VTAIL.n105 VSUBS 0.058486f
C1465 VTAIL.n106 VSUBS 0.040036f
C1466 VTAIL.n107 VSUBS 0.221976f
C1467 VTAIL.t12 VSUBS 0.405461f
C1468 VTAIL.t19 VSUBS 0.405461f
C1469 VTAIL.n108 VSUBS 3.1878f
C1470 VTAIL.n109 VSUBS 0.915844f
C1471 VTAIL.t15 VSUBS 0.405461f
C1472 VTAIL.t11 VSUBS 0.405461f
C1473 VTAIL.n110 VSUBS 3.1878f
C1474 VTAIL.n111 VSUBS 2.81771f
C1475 VTAIL.t9 VSUBS 0.405461f
C1476 VTAIL.t7 VSUBS 0.405461f
C1477 VTAIL.n112 VSUBS 3.18781f
C1478 VTAIL.n113 VSUBS 2.8177f
C1479 VTAIL.t8 VSUBS 0.405461f
C1480 VTAIL.t2 VSUBS 0.405461f
C1481 VTAIL.n114 VSUBS 3.18781f
C1482 VTAIL.n115 VSUBS 0.915832f
C1483 VTAIL.n116 VSUBS 0.028887f
C1484 VTAIL.n117 VSUBS 0.027234f
C1485 VTAIL.n118 VSUBS 0.014634f
C1486 VTAIL.n119 VSUBS 0.034591f
C1487 VTAIL.n120 VSUBS 0.015495f
C1488 VTAIL.n121 VSUBS 0.027234f
C1489 VTAIL.n122 VSUBS 0.014634f
C1490 VTAIL.n123 VSUBS 0.034591f
C1491 VTAIL.n124 VSUBS 0.015495f
C1492 VTAIL.n125 VSUBS 0.027234f
C1493 VTAIL.n126 VSUBS 0.014634f
C1494 VTAIL.n127 VSUBS 0.034591f
C1495 VTAIL.n128 VSUBS 0.015495f
C1496 VTAIL.n129 VSUBS 0.027234f
C1497 VTAIL.n130 VSUBS 0.014634f
C1498 VTAIL.n131 VSUBS 0.034591f
C1499 VTAIL.n132 VSUBS 0.034591f
C1500 VTAIL.n133 VSUBS 0.015495f
C1501 VTAIL.n134 VSUBS 0.027234f
C1502 VTAIL.n135 VSUBS 0.014634f
C1503 VTAIL.n136 VSUBS 0.034591f
C1504 VTAIL.n137 VSUBS 0.015495f
C1505 VTAIL.n138 VSUBS 0.027234f
C1506 VTAIL.n139 VSUBS 0.014634f
C1507 VTAIL.n140 VSUBS 0.034591f
C1508 VTAIL.n141 VSUBS 0.015495f
C1509 VTAIL.n142 VSUBS 0.027234f
C1510 VTAIL.n143 VSUBS 0.014634f
C1511 VTAIL.n144 VSUBS 0.034591f
C1512 VTAIL.n145 VSUBS 0.015495f
C1513 VTAIL.n146 VSUBS 0.027234f
C1514 VTAIL.n147 VSUBS 0.014634f
C1515 VTAIL.n148 VSUBS 0.034591f
C1516 VTAIL.n149 VSUBS 0.015495f
C1517 VTAIL.n150 VSUBS 0.222824f
C1518 VTAIL.t5 VSUBS 0.074312f
C1519 VTAIL.n151 VSUBS 0.025943f
C1520 VTAIL.n152 VSUBS 0.022005f
C1521 VTAIL.n153 VSUBS 0.014634f
C1522 VTAIL.n154 VSUBS 2.21372f
C1523 VTAIL.n155 VSUBS 0.027234f
C1524 VTAIL.n156 VSUBS 0.014634f
C1525 VTAIL.n157 VSUBS 0.015495f
C1526 VTAIL.n158 VSUBS 0.034591f
C1527 VTAIL.n159 VSUBS 0.034591f
C1528 VTAIL.n160 VSUBS 0.015495f
C1529 VTAIL.n161 VSUBS 0.014634f
C1530 VTAIL.n162 VSUBS 0.027234f
C1531 VTAIL.n163 VSUBS 0.027234f
C1532 VTAIL.n164 VSUBS 0.014634f
C1533 VTAIL.n165 VSUBS 0.015495f
C1534 VTAIL.n166 VSUBS 0.034591f
C1535 VTAIL.n167 VSUBS 0.034591f
C1536 VTAIL.n168 VSUBS 0.015495f
C1537 VTAIL.n169 VSUBS 0.014634f
C1538 VTAIL.n170 VSUBS 0.027234f
C1539 VTAIL.n171 VSUBS 0.027234f
C1540 VTAIL.n172 VSUBS 0.014634f
C1541 VTAIL.n173 VSUBS 0.015495f
C1542 VTAIL.n174 VSUBS 0.034591f
C1543 VTAIL.n175 VSUBS 0.034591f
C1544 VTAIL.n176 VSUBS 0.015495f
C1545 VTAIL.n177 VSUBS 0.014634f
C1546 VTAIL.n178 VSUBS 0.027234f
C1547 VTAIL.n179 VSUBS 0.027234f
C1548 VTAIL.n180 VSUBS 0.014634f
C1549 VTAIL.n181 VSUBS 0.015495f
C1550 VTAIL.n182 VSUBS 0.034591f
C1551 VTAIL.n183 VSUBS 0.034591f
C1552 VTAIL.n184 VSUBS 0.015495f
C1553 VTAIL.n185 VSUBS 0.014634f
C1554 VTAIL.n186 VSUBS 0.027234f
C1555 VTAIL.n187 VSUBS 0.027234f
C1556 VTAIL.n188 VSUBS 0.014634f
C1557 VTAIL.n189 VSUBS 0.015495f
C1558 VTAIL.n190 VSUBS 0.034591f
C1559 VTAIL.n191 VSUBS 0.034591f
C1560 VTAIL.n192 VSUBS 0.015495f
C1561 VTAIL.n193 VSUBS 0.014634f
C1562 VTAIL.n194 VSUBS 0.027234f
C1563 VTAIL.n195 VSUBS 0.027234f
C1564 VTAIL.n196 VSUBS 0.014634f
C1565 VTAIL.n197 VSUBS 0.015065f
C1566 VTAIL.n198 VSUBS 0.015065f
C1567 VTAIL.n199 VSUBS 0.034591f
C1568 VTAIL.n200 VSUBS 0.034591f
C1569 VTAIL.n201 VSUBS 0.015495f
C1570 VTAIL.n202 VSUBS 0.014634f
C1571 VTAIL.n203 VSUBS 0.027234f
C1572 VTAIL.n204 VSUBS 0.027234f
C1573 VTAIL.n205 VSUBS 0.014634f
C1574 VTAIL.n206 VSUBS 0.015495f
C1575 VTAIL.n207 VSUBS 0.034591f
C1576 VTAIL.n208 VSUBS 0.034591f
C1577 VTAIL.n209 VSUBS 0.015495f
C1578 VTAIL.n210 VSUBS 0.014634f
C1579 VTAIL.n211 VSUBS 0.027234f
C1580 VTAIL.n212 VSUBS 0.027234f
C1581 VTAIL.n213 VSUBS 0.014634f
C1582 VTAIL.n214 VSUBS 0.015495f
C1583 VTAIL.n215 VSUBS 0.034591f
C1584 VTAIL.n216 VSUBS 0.080206f
C1585 VTAIL.n217 VSUBS 0.015495f
C1586 VTAIL.n218 VSUBS 0.014634f
C1587 VTAIL.n219 VSUBS 0.058486f
C1588 VTAIL.n220 VSUBS 0.040036f
C1589 VTAIL.n221 VSUBS 0.221976f
C1590 VTAIL.t18 VSUBS 0.405461f
C1591 VTAIL.t13 VSUBS 0.405461f
C1592 VTAIL.n222 VSUBS 3.18781f
C1593 VTAIL.n223 VSUBS 0.903728f
C1594 VTAIL.t17 VSUBS 0.405461f
C1595 VTAIL.t10 VSUBS 0.405461f
C1596 VTAIL.n224 VSUBS 3.18781f
C1597 VTAIL.n225 VSUBS 0.915832f
C1598 VTAIL.n226 VSUBS 0.028887f
C1599 VTAIL.n227 VSUBS 0.027234f
C1600 VTAIL.n228 VSUBS 0.014634f
C1601 VTAIL.n229 VSUBS 0.034591f
C1602 VTAIL.n230 VSUBS 0.015495f
C1603 VTAIL.n231 VSUBS 0.027234f
C1604 VTAIL.n232 VSUBS 0.014634f
C1605 VTAIL.n233 VSUBS 0.034591f
C1606 VTAIL.n234 VSUBS 0.015495f
C1607 VTAIL.n235 VSUBS 0.027234f
C1608 VTAIL.n236 VSUBS 0.014634f
C1609 VTAIL.n237 VSUBS 0.034591f
C1610 VTAIL.n238 VSUBS 0.015495f
C1611 VTAIL.n239 VSUBS 0.027234f
C1612 VTAIL.n240 VSUBS 0.014634f
C1613 VTAIL.n241 VSUBS 0.034591f
C1614 VTAIL.n242 VSUBS 0.034591f
C1615 VTAIL.n243 VSUBS 0.015495f
C1616 VTAIL.n244 VSUBS 0.027234f
C1617 VTAIL.n245 VSUBS 0.014634f
C1618 VTAIL.n246 VSUBS 0.034591f
C1619 VTAIL.n247 VSUBS 0.015495f
C1620 VTAIL.n248 VSUBS 0.027234f
C1621 VTAIL.n249 VSUBS 0.014634f
C1622 VTAIL.n250 VSUBS 0.034591f
C1623 VTAIL.n251 VSUBS 0.015495f
C1624 VTAIL.n252 VSUBS 0.027234f
C1625 VTAIL.n253 VSUBS 0.014634f
C1626 VTAIL.n254 VSUBS 0.034591f
C1627 VTAIL.n255 VSUBS 0.015495f
C1628 VTAIL.n256 VSUBS 0.027234f
C1629 VTAIL.n257 VSUBS 0.014634f
C1630 VTAIL.n258 VSUBS 0.034591f
C1631 VTAIL.n259 VSUBS 0.015495f
C1632 VTAIL.n260 VSUBS 0.222824f
C1633 VTAIL.t16 VSUBS 0.074312f
C1634 VTAIL.n261 VSUBS 0.025943f
C1635 VTAIL.n262 VSUBS 0.022005f
C1636 VTAIL.n263 VSUBS 0.014634f
C1637 VTAIL.n264 VSUBS 2.21372f
C1638 VTAIL.n265 VSUBS 0.027234f
C1639 VTAIL.n266 VSUBS 0.014634f
C1640 VTAIL.n267 VSUBS 0.015495f
C1641 VTAIL.n268 VSUBS 0.034591f
C1642 VTAIL.n269 VSUBS 0.034591f
C1643 VTAIL.n270 VSUBS 0.015495f
C1644 VTAIL.n271 VSUBS 0.014634f
C1645 VTAIL.n272 VSUBS 0.027234f
C1646 VTAIL.n273 VSUBS 0.027234f
C1647 VTAIL.n274 VSUBS 0.014634f
C1648 VTAIL.n275 VSUBS 0.015495f
C1649 VTAIL.n276 VSUBS 0.034591f
C1650 VTAIL.n277 VSUBS 0.034591f
C1651 VTAIL.n278 VSUBS 0.015495f
C1652 VTAIL.n279 VSUBS 0.014634f
C1653 VTAIL.n280 VSUBS 0.027234f
C1654 VTAIL.n281 VSUBS 0.027234f
C1655 VTAIL.n282 VSUBS 0.014634f
C1656 VTAIL.n283 VSUBS 0.015495f
C1657 VTAIL.n284 VSUBS 0.034591f
C1658 VTAIL.n285 VSUBS 0.034591f
C1659 VTAIL.n286 VSUBS 0.015495f
C1660 VTAIL.n287 VSUBS 0.014634f
C1661 VTAIL.n288 VSUBS 0.027234f
C1662 VTAIL.n289 VSUBS 0.027234f
C1663 VTAIL.n290 VSUBS 0.014634f
C1664 VTAIL.n291 VSUBS 0.015495f
C1665 VTAIL.n292 VSUBS 0.034591f
C1666 VTAIL.n293 VSUBS 0.034591f
C1667 VTAIL.n294 VSUBS 0.015495f
C1668 VTAIL.n295 VSUBS 0.014634f
C1669 VTAIL.n296 VSUBS 0.027234f
C1670 VTAIL.n297 VSUBS 0.027234f
C1671 VTAIL.n298 VSUBS 0.014634f
C1672 VTAIL.n299 VSUBS 0.015495f
C1673 VTAIL.n300 VSUBS 0.034591f
C1674 VTAIL.n301 VSUBS 0.034591f
C1675 VTAIL.n302 VSUBS 0.015495f
C1676 VTAIL.n303 VSUBS 0.014634f
C1677 VTAIL.n304 VSUBS 0.027234f
C1678 VTAIL.n305 VSUBS 0.027234f
C1679 VTAIL.n306 VSUBS 0.014634f
C1680 VTAIL.n307 VSUBS 0.015065f
C1681 VTAIL.n308 VSUBS 0.015065f
C1682 VTAIL.n309 VSUBS 0.034591f
C1683 VTAIL.n310 VSUBS 0.034591f
C1684 VTAIL.n311 VSUBS 0.015495f
C1685 VTAIL.n312 VSUBS 0.014634f
C1686 VTAIL.n313 VSUBS 0.027234f
C1687 VTAIL.n314 VSUBS 0.027234f
C1688 VTAIL.n315 VSUBS 0.014634f
C1689 VTAIL.n316 VSUBS 0.015495f
C1690 VTAIL.n317 VSUBS 0.034591f
C1691 VTAIL.n318 VSUBS 0.034591f
C1692 VTAIL.n319 VSUBS 0.015495f
C1693 VTAIL.n320 VSUBS 0.014634f
C1694 VTAIL.n321 VSUBS 0.027234f
C1695 VTAIL.n322 VSUBS 0.027234f
C1696 VTAIL.n323 VSUBS 0.014634f
C1697 VTAIL.n324 VSUBS 0.015495f
C1698 VTAIL.n325 VSUBS 0.034591f
C1699 VTAIL.n326 VSUBS 0.080206f
C1700 VTAIL.n327 VSUBS 0.015495f
C1701 VTAIL.n328 VSUBS 0.014634f
C1702 VTAIL.n329 VSUBS 0.058486f
C1703 VTAIL.n330 VSUBS 0.040036f
C1704 VTAIL.n331 VSUBS 2.02928f
C1705 VTAIL.n332 VSUBS 0.028887f
C1706 VTAIL.n333 VSUBS 0.027234f
C1707 VTAIL.n334 VSUBS 0.014634f
C1708 VTAIL.n335 VSUBS 0.034591f
C1709 VTAIL.n336 VSUBS 0.015495f
C1710 VTAIL.n337 VSUBS 0.027234f
C1711 VTAIL.n338 VSUBS 0.014634f
C1712 VTAIL.n339 VSUBS 0.034591f
C1713 VTAIL.n340 VSUBS 0.015495f
C1714 VTAIL.n341 VSUBS 0.027234f
C1715 VTAIL.n342 VSUBS 0.014634f
C1716 VTAIL.n343 VSUBS 0.034591f
C1717 VTAIL.n344 VSUBS 0.015495f
C1718 VTAIL.n345 VSUBS 0.027234f
C1719 VTAIL.n346 VSUBS 0.014634f
C1720 VTAIL.n347 VSUBS 0.034591f
C1721 VTAIL.n348 VSUBS 0.015495f
C1722 VTAIL.n349 VSUBS 0.027234f
C1723 VTAIL.n350 VSUBS 0.014634f
C1724 VTAIL.n351 VSUBS 0.034591f
C1725 VTAIL.n352 VSUBS 0.015495f
C1726 VTAIL.n353 VSUBS 0.027234f
C1727 VTAIL.n354 VSUBS 0.014634f
C1728 VTAIL.n355 VSUBS 0.034591f
C1729 VTAIL.n356 VSUBS 0.015495f
C1730 VTAIL.n357 VSUBS 0.027234f
C1731 VTAIL.n358 VSUBS 0.014634f
C1732 VTAIL.n359 VSUBS 0.034591f
C1733 VTAIL.n360 VSUBS 0.015495f
C1734 VTAIL.n361 VSUBS 0.027234f
C1735 VTAIL.n362 VSUBS 0.014634f
C1736 VTAIL.n363 VSUBS 0.034591f
C1737 VTAIL.n364 VSUBS 0.015495f
C1738 VTAIL.n365 VSUBS 0.222824f
C1739 VTAIL.t3 VSUBS 0.074312f
C1740 VTAIL.n366 VSUBS 0.025943f
C1741 VTAIL.n367 VSUBS 0.022005f
C1742 VTAIL.n368 VSUBS 0.014634f
C1743 VTAIL.n369 VSUBS 2.21372f
C1744 VTAIL.n370 VSUBS 0.027234f
C1745 VTAIL.n371 VSUBS 0.014634f
C1746 VTAIL.n372 VSUBS 0.015495f
C1747 VTAIL.n373 VSUBS 0.034591f
C1748 VTAIL.n374 VSUBS 0.034591f
C1749 VTAIL.n375 VSUBS 0.015495f
C1750 VTAIL.n376 VSUBS 0.014634f
C1751 VTAIL.n377 VSUBS 0.027234f
C1752 VTAIL.n378 VSUBS 0.027234f
C1753 VTAIL.n379 VSUBS 0.014634f
C1754 VTAIL.n380 VSUBS 0.015495f
C1755 VTAIL.n381 VSUBS 0.034591f
C1756 VTAIL.n382 VSUBS 0.034591f
C1757 VTAIL.n383 VSUBS 0.015495f
C1758 VTAIL.n384 VSUBS 0.014634f
C1759 VTAIL.n385 VSUBS 0.027234f
C1760 VTAIL.n386 VSUBS 0.027234f
C1761 VTAIL.n387 VSUBS 0.014634f
C1762 VTAIL.n388 VSUBS 0.015495f
C1763 VTAIL.n389 VSUBS 0.034591f
C1764 VTAIL.n390 VSUBS 0.034591f
C1765 VTAIL.n391 VSUBS 0.015495f
C1766 VTAIL.n392 VSUBS 0.014634f
C1767 VTAIL.n393 VSUBS 0.027234f
C1768 VTAIL.n394 VSUBS 0.027234f
C1769 VTAIL.n395 VSUBS 0.014634f
C1770 VTAIL.n396 VSUBS 0.015495f
C1771 VTAIL.n397 VSUBS 0.034591f
C1772 VTAIL.n398 VSUBS 0.034591f
C1773 VTAIL.n399 VSUBS 0.015495f
C1774 VTAIL.n400 VSUBS 0.014634f
C1775 VTAIL.n401 VSUBS 0.027234f
C1776 VTAIL.n402 VSUBS 0.027234f
C1777 VTAIL.n403 VSUBS 0.014634f
C1778 VTAIL.n404 VSUBS 0.015495f
C1779 VTAIL.n405 VSUBS 0.034591f
C1780 VTAIL.n406 VSUBS 0.034591f
C1781 VTAIL.n407 VSUBS 0.034591f
C1782 VTAIL.n408 VSUBS 0.015495f
C1783 VTAIL.n409 VSUBS 0.014634f
C1784 VTAIL.n410 VSUBS 0.027234f
C1785 VTAIL.n411 VSUBS 0.027234f
C1786 VTAIL.n412 VSUBS 0.014634f
C1787 VTAIL.n413 VSUBS 0.015065f
C1788 VTAIL.n414 VSUBS 0.015065f
C1789 VTAIL.n415 VSUBS 0.034591f
C1790 VTAIL.n416 VSUBS 0.034591f
C1791 VTAIL.n417 VSUBS 0.015495f
C1792 VTAIL.n418 VSUBS 0.014634f
C1793 VTAIL.n419 VSUBS 0.027234f
C1794 VTAIL.n420 VSUBS 0.027234f
C1795 VTAIL.n421 VSUBS 0.014634f
C1796 VTAIL.n422 VSUBS 0.015495f
C1797 VTAIL.n423 VSUBS 0.034591f
C1798 VTAIL.n424 VSUBS 0.034591f
C1799 VTAIL.n425 VSUBS 0.015495f
C1800 VTAIL.n426 VSUBS 0.014634f
C1801 VTAIL.n427 VSUBS 0.027234f
C1802 VTAIL.n428 VSUBS 0.027234f
C1803 VTAIL.n429 VSUBS 0.014634f
C1804 VTAIL.n430 VSUBS 0.015495f
C1805 VTAIL.n431 VSUBS 0.034591f
C1806 VTAIL.n432 VSUBS 0.080206f
C1807 VTAIL.n433 VSUBS 0.015495f
C1808 VTAIL.n434 VSUBS 0.014634f
C1809 VTAIL.n435 VSUBS 0.058486f
C1810 VTAIL.n436 VSUBS 0.040036f
C1811 VTAIL.n437 VSUBS 2.02928f
C1812 VTAIL.t4 VSUBS 0.405461f
C1813 VTAIL.t0 VSUBS 0.405461f
C1814 VTAIL.n438 VSUBS 3.1878f
C1815 VTAIL.n439 VSUBS 0.830737f
C1816 VP.n0 VSUBS 0.055265f
C1817 VP.t2 VSUBS 2.31989f
C1818 VP.n1 VSUBS 0.825141f
C1819 VP.n2 VSUBS 0.041417f
C1820 VP.t9 VSUBS 2.31989f
C1821 VP.n3 VSUBS 0.055049f
C1822 VP.n4 VSUBS 0.041417f
C1823 VP.t1 VSUBS 2.31989f
C1824 VP.t4 VSUBS 2.388f
C1825 VP.n5 VSUBS 0.892005f
C1826 VP.n6 VSUBS 0.055265f
C1827 VP.t0 VSUBS 2.388f
C1828 VP.t3 VSUBS 2.31989f
C1829 VP.n7 VSUBS 0.825141f
C1830 VP.n8 VSUBS 0.041417f
C1831 VP.t5 VSUBS 2.31989f
C1832 VP.n9 VSUBS 0.055049f
C1833 VP.t7 VSUBS 2.42773f
C1834 VP.n10 VSUBS 0.882231f
C1835 VP.t6 VSUBS 2.31989f
C1836 VP.n11 VSUBS 0.883811f
C1837 VP.n12 VSUBS 0.058537f
C1838 VP.n13 VSUBS 0.21079f
C1839 VP.n14 VSUBS 0.041417f
C1840 VP.n15 VSUBS 0.041417f
C1841 VP.n16 VSUBS 0.864028f
C1842 VP.n17 VSUBS 0.055049f
C1843 VP.n18 VSUBS 0.058537f
C1844 VP.n19 VSUBS 0.041417f
C1845 VP.n20 VSUBS 0.041417f
C1846 VP.n21 VSUBS 0.050704f
C1847 VP.n22 VSUBS 0.036016f
C1848 VP.n23 VSUBS 0.892005f
C1849 VP.n24 VSUBS 2.27546f
C1850 VP.n25 VSUBS 2.30524f
C1851 VP.n26 VSUBS 0.055265f
C1852 VP.n27 VSUBS 0.036016f
C1853 VP.n28 VSUBS 0.050704f
C1854 VP.n29 VSUBS 0.825141f
C1855 VP.n30 VSUBS 0.058537f
C1856 VP.n31 VSUBS 0.041417f
C1857 VP.n32 VSUBS 0.041417f
C1858 VP.n33 VSUBS 0.041417f
C1859 VP.n34 VSUBS 0.864028f
C1860 VP.n35 VSUBS 0.055049f
C1861 VP.n36 VSUBS 0.058537f
C1862 VP.n37 VSUBS 0.041417f
C1863 VP.n38 VSUBS 0.041417f
C1864 VP.n39 VSUBS 0.050704f
C1865 VP.n40 VSUBS 0.036016f
C1866 VP.t8 VSUBS 2.388f
C1867 VP.n41 VSUBS 0.892005f
C1868 VP.n42 VSUBS 0.038788f
.ends

