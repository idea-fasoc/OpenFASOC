* NGSPICE file created from diff_pair_sample_1407.ext - technology: sky130A

.subckt diff_pair_sample_1407 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t7 VN.t0 VTAIL.t10 w_n4230_n2876# sky130_fd_pr__pfet_01v8 ad=1.5741 pd=9.87 as=1.5741 ps=9.87 w=9.54 l=2.93
X1 VTAIL.t1 VP.t0 VDD1.t7 w_n4230_n2876# sky130_fd_pr__pfet_01v8 ad=3.7206 pd=19.86 as=1.5741 ps=9.87 w=9.54 l=2.93
X2 B.t11 B.t9 B.t10 w_n4230_n2876# sky130_fd_pr__pfet_01v8 ad=3.7206 pd=19.86 as=0 ps=0 w=9.54 l=2.93
X3 VDD2.t6 VN.t1 VTAIL.t14 w_n4230_n2876# sky130_fd_pr__pfet_01v8 ad=1.5741 pd=9.87 as=3.7206 ps=19.86 w=9.54 l=2.93
X4 VDD1.t6 VP.t1 VTAIL.t3 w_n4230_n2876# sky130_fd_pr__pfet_01v8 ad=1.5741 pd=9.87 as=1.5741 ps=9.87 w=9.54 l=2.93
X5 VDD2.t5 VN.t2 VTAIL.t11 w_n4230_n2876# sky130_fd_pr__pfet_01v8 ad=1.5741 pd=9.87 as=1.5741 ps=9.87 w=9.54 l=2.93
X6 VTAIL.t15 VN.t3 VDD2.t4 w_n4230_n2876# sky130_fd_pr__pfet_01v8 ad=3.7206 pd=19.86 as=1.5741 ps=9.87 w=9.54 l=2.93
X7 VDD2.t3 VN.t4 VTAIL.t13 w_n4230_n2876# sky130_fd_pr__pfet_01v8 ad=1.5741 pd=9.87 as=3.7206 ps=19.86 w=9.54 l=2.93
X8 VTAIL.t8 VN.t5 VDD2.t2 w_n4230_n2876# sky130_fd_pr__pfet_01v8 ad=3.7206 pd=19.86 as=1.5741 ps=9.87 w=9.54 l=2.93
X9 VDD1.t5 VP.t2 VTAIL.t5 w_n4230_n2876# sky130_fd_pr__pfet_01v8 ad=1.5741 pd=9.87 as=1.5741 ps=9.87 w=9.54 l=2.93
X10 B.t8 B.t6 B.t7 w_n4230_n2876# sky130_fd_pr__pfet_01v8 ad=3.7206 pd=19.86 as=0 ps=0 w=9.54 l=2.93
X11 VTAIL.t7 VP.t3 VDD1.t4 w_n4230_n2876# sky130_fd_pr__pfet_01v8 ad=1.5741 pd=9.87 as=1.5741 ps=9.87 w=9.54 l=2.93
X12 VTAIL.t0 VP.t4 VDD1.t3 w_n4230_n2876# sky130_fd_pr__pfet_01v8 ad=1.5741 pd=9.87 as=1.5741 ps=9.87 w=9.54 l=2.93
X13 B.t5 B.t3 B.t4 w_n4230_n2876# sky130_fd_pr__pfet_01v8 ad=3.7206 pd=19.86 as=0 ps=0 w=9.54 l=2.93
X14 VTAIL.t9 VN.t6 VDD2.t1 w_n4230_n2876# sky130_fd_pr__pfet_01v8 ad=1.5741 pd=9.87 as=1.5741 ps=9.87 w=9.54 l=2.93
X15 VTAIL.t12 VN.t7 VDD2.t0 w_n4230_n2876# sky130_fd_pr__pfet_01v8 ad=1.5741 pd=9.87 as=1.5741 ps=9.87 w=9.54 l=2.93
X16 VDD1.t2 VP.t5 VTAIL.t2 w_n4230_n2876# sky130_fd_pr__pfet_01v8 ad=1.5741 pd=9.87 as=3.7206 ps=19.86 w=9.54 l=2.93
X17 B.t2 B.t0 B.t1 w_n4230_n2876# sky130_fd_pr__pfet_01v8 ad=3.7206 pd=19.86 as=0 ps=0 w=9.54 l=2.93
X18 VTAIL.t6 VP.t6 VDD1.t1 w_n4230_n2876# sky130_fd_pr__pfet_01v8 ad=3.7206 pd=19.86 as=1.5741 ps=9.87 w=9.54 l=2.93
X19 VDD1.t0 VP.t7 VTAIL.t4 w_n4230_n2876# sky130_fd_pr__pfet_01v8 ad=1.5741 pd=9.87 as=3.7206 ps=19.86 w=9.54 l=2.93
R0 VN.n60 VN.n59 161.3
R1 VN.n58 VN.n32 161.3
R2 VN.n57 VN.n56 161.3
R3 VN.n55 VN.n33 161.3
R4 VN.n54 VN.n53 161.3
R5 VN.n52 VN.n34 161.3
R6 VN.n50 VN.n49 161.3
R7 VN.n48 VN.n35 161.3
R8 VN.n47 VN.n46 161.3
R9 VN.n45 VN.n36 161.3
R10 VN.n44 VN.n43 161.3
R11 VN.n42 VN.n37 161.3
R12 VN.n41 VN.n40 161.3
R13 VN.n29 VN.n28 161.3
R14 VN.n27 VN.n1 161.3
R15 VN.n26 VN.n25 161.3
R16 VN.n24 VN.n2 161.3
R17 VN.n23 VN.n22 161.3
R18 VN.n21 VN.n3 161.3
R19 VN.n19 VN.n18 161.3
R20 VN.n17 VN.n4 161.3
R21 VN.n16 VN.n15 161.3
R22 VN.n14 VN.n5 161.3
R23 VN.n13 VN.n12 161.3
R24 VN.n11 VN.n6 161.3
R25 VN.n10 VN.n9 161.3
R26 VN.n38 VN.t4 110.206
R27 VN.n7 VN.t5 110.206
R28 VN.n8 VN.t0 78.4694
R29 VN.n20 VN.t6 78.4694
R30 VN.n0 VN.t1 78.4694
R31 VN.n39 VN.t7 78.4694
R32 VN.n51 VN.t2 78.4694
R33 VN.n31 VN.t3 78.4694
R34 VN.n30 VN.n0 71.0639
R35 VN.n61 VN.n31 71.0639
R36 VN.n8 VN.n7 67.4245
R37 VN.n39 VN.n38 67.4245
R38 VN.n26 VN.n2 56.5617
R39 VN.n57 VN.n33 56.5617
R40 VN VN.n61 50.8315
R41 VN.n14 VN.n13 40.577
R42 VN.n15 VN.n14 40.577
R43 VN.n45 VN.n44 40.577
R44 VN.n46 VN.n45 40.577
R45 VN.n9 VN.n6 24.5923
R46 VN.n13 VN.n6 24.5923
R47 VN.n15 VN.n4 24.5923
R48 VN.n19 VN.n4 24.5923
R49 VN.n22 VN.n21 24.5923
R50 VN.n22 VN.n2 24.5923
R51 VN.n27 VN.n26 24.5923
R52 VN.n28 VN.n27 24.5923
R53 VN.n44 VN.n37 24.5923
R54 VN.n40 VN.n37 24.5923
R55 VN.n53 VN.n33 24.5923
R56 VN.n53 VN.n52 24.5923
R57 VN.n50 VN.n35 24.5923
R58 VN.n46 VN.n35 24.5923
R59 VN.n59 VN.n58 24.5923
R60 VN.n58 VN.n57 24.5923
R61 VN.n28 VN.n0 19.1821
R62 VN.n59 VN.n31 19.1821
R63 VN.n21 VN.n20 18.1985
R64 VN.n52 VN.n51 18.1985
R65 VN.n9 VN.n8 6.39438
R66 VN.n20 VN.n19 6.39438
R67 VN.n40 VN.n39 6.39438
R68 VN.n51 VN.n50 6.39438
R69 VN.n10 VN.n7 5.60224
R70 VN.n41 VN.n38 5.60224
R71 VN.n61 VN.n60 0.354861
R72 VN.n30 VN.n29 0.354861
R73 VN VN.n30 0.267071
R74 VN.n60 VN.n32 0.189894
R75 VN.n56 VN.n32 0.189894
R76 VN.n56 VN.n55 0.189894
R77 VN.n55 VN.n54 0.189894
R78 VN.n54 VN.n34 0.189894
R79 VN.n49 VN.n34 0.189894
R80 VN.n49 VN.n48 0.189894
R81 VN.n48 VN.n47 0.189894
R82 VN.n47 VN.n36 0.189894
R83 VN.n43 VN.n36 0.189894
R84 VN.n43 VN.n42 0.189894
R85 VN.n42 VN.n41 0.189894
R86 VN.n11 VN.n10 0.189894
R87 VN.n12 VN.n11 0.189894
R88 VN.n12 VN.n5 0.189894
R89 VN.n16 VN.n5 0.189894
R90 VN.n17 VN.n16 0.189894
R91 VN.n18 VN.n17 0.189894
R92 VN.n18 VN.n3 0.189894
R93 VN.n23 VN.n3 0.189894
R94 VN.n24 VN.n23 0.189894
R95 VN.n25 VN.n24 0.189894
R96 VN.n25 VN.n1 0.189894
R97 VN.n29 VN.n1 0.189894
R98 VTAIL.n11 VTAIL.t1 63.3851
R99 VTAIL.n10 VTAIL.t13 63.3851
R100 VTAIL.n7 VTAIL.t15 63.3851
R101 VTAIL.n15 VTAIL.t14 63.385
R102 VTAIL.n2 VTAIL.t8 63.385
R103 VTAIL.n3 VTAIL.t4 63.385
R104 VTAIL.n6 VTAIL.t6 63.385
R105 VTAIL.n14 VTAIL.t2 63.385
R106 VTAIL.n13 VTAIL.n12 59.978
R107 VTAIL.n9 VTAIL.n8 59.978
R108 VTAIL.n1 VTAIL.n0 59.9777
R109 VTAIL.n5 VTAIL.n4 59.9777
R110 VTAIL.n15 VTAIL.n14 23.4014
R111 VTAIL.n7 VTAIL.n6 23.4014
R112 VTAIL.n0 VTAIL.t10 3.40773
R113 VTAIL.n0 VTAIL.t9 3.40773
R114 VTAIL.n4 VTAIL.t5 3.40773
R115 VTAIL.n4 VTAIL.t0 3.40773
R116 VTAIL.n12 VTAIL.t3 3.40773
R117 VTAIL.n12 VTAIL.t7 3.40773
R118 VTAIL.n8 VTAIL.t11 3.40773
R119 VTAIL.n8 VTAIL.t12 3.40773
R120 VTAIL.n9 VTAIL.n7 2.81084
R121 VTAIL.n10 VTAIL.n9 2.81084
R122 VTAIL.n13 VTAIL.n11 2.81084
R123 VTAIL.n14 VTAIL.n13 2.81084
R124 VTAIL.n6 VTAIL.n5 2.81084
R125 VTAIL.n5 VTAIL.n3 2.81084
R126 VTAIL.n2 VTAIL.n1 2.81084
R127 VTAIL VTAIL.n15 2.75266
R128 VTAIL.n11 VTAIL.n10 0.470328
R129 VTAIL.n3 VTAIL.n2 0.470328
R130 VTAIL VTAIL.n1 0.0586897
R131 VDD2.n2 VDD2.n1 78.0063
R132 VDD2.n2 VDD2.n0 78.0063
R133 VDD2 VDD2.n5 78.0035
R134 VDD2.n4 VDD2.n3 76.6568
R135 VDD2.n4 VDD2.n2 44.586
R136 VDD2.n5 VDD2.t0 3.40773
R137 VDD2.n5 VDD2.t3 3.40773
R138 VDD2.n3 VDD2.t4 3.40773
R139 VDD2.n3 VDD2.t5 3.40773
R140 VDD2.n1 VDD2.t1 3.40773
R141 VDD2.n1 VDD2.t6 3.40773
R142 VDD2.n0 VDD2.t2 3.40773
R143 VDD2.n0 VDD2.t7 3.40773
R144 VDD2 VDD2.n4 1.46386
R145 VP.n21 VP.n20 161.3
R146 VP.n22 VP.n17 161.3
R147 VP.n24 VP.n23 161.3
R148 VP.n25 VP.n16 161.3
R149 VP.n27 VP.n26 161.3
R150 VP.n28 VP.n15 161.3
R151 VP.n30 VP.n29 161.3
R152 VP.n32 VP.n14 161.3
R153 VP.n34 VP.n33 161.3
R154 VP.n35 VP.n13 161.3
R155 VP.n37 VP.n36 161.3
R156 VP.n38 VP.n12 161.3
R157 VP.n40 VP.n39 161.3
R158 VP.n73 VP.n72 161.3
R159 VP.n71 VP.n1 161.3
R160 VP.n70 VP.n69 161.3
R161 VP.n68 VP.n2 161.3
R162 VP.n67 VP.n66 161.3
R163 VP.n65 VP.n3 161.3
R164 VP.n63 VP.n62 161.3
R165 VP.n61 VP.n4 161.3
R166 VP.n60 VP.n59 161.3
R167 VP.n58 VP.n5 161.3
R168 VP.n57 VP.n56 161.3
R169 VP.n55 VP.n6 161.3
R170 VP.n54 VP.n53 161.3
R171 VP.n51 VP.n7 161.3
R172 VP.n50 VP.n49 161.3
R173 VP.n48 VP.n8 161.3
R174 VP.n47 VP.n46 161.3
R175 VP.n45 VP.n9 161.3
R176 VP.n44 VP.n43 161.3
R177 VP.n18 VP.t0 110.206
R178 VP.n10 VP.t6 78.4694
R179 VP.n52 VP.t2 78.4694
R180 VP.n64 VP.t4 78.4694
R181 VP.n0 VP.t7 78.4694
R182 VP.n11 VP.t5 78.4694
R183 VP.n31 VP.t3 78.4694
R184 VP.n19 VP.t1 78.4694
R185 VP.n42 VP.n10 71.0639
R186 VP.n74 VP.n0 71.0639
R187 VP.n41 VP.n11 71.0639
R188 VP.n19 VP.n18 67.4245
R189 VP.n46 VP.n8 56.5617
R190 VP.n37 VP.n13 56.5617
R191 VP.n70 VP.n2 56.5617
R192 VP.n42 VP.n41 50.6662
R193 VP.n58 VP.n57 40.577
R194 VP.n59 VP.n58 40.577
R195 VP.n26 VP.n25 40.577
R196 VP.n25 VP.n24 40.577
R197 VP.n45 VP.n44 24.5923
R198 VP.n46 VP.n45 24.5923
R199 VP.n50 VP.n8 24.5923
R200 VP.n51 VP.n50 24.5923
R201 VP.n53 VP.n6 24.5923
R202 VP.n57 VP.n6 24.5923
R203 VP.n59 VP.n4 24.5923
R204 VP.n63 VP.n4 24.5923
R205 VP.n66 VP.n65 24.5923
R206 VP.n66 VP.n2 24.5923
R207 VP.n71 VP.n70 24.5923
R208 VP.n72 VP.n71 24.5923
R209 VP.n38 VP.n37 24.5923
R210 VP.n39 VP.n38 24.5923
R211 VP.n26 VP.n15 24.5923
R212 VP.n30 VP.n15 24.5923
R213 VP.n33 VP.n32 24.5923
R214 VP.n33 VP.n13 24.5923
R215 VP.n20 VP.n17 24.5923
R216 VP.n24 VP.n17 24.5923
R217 VP.n44 VP.n10 19.1821
R218 VP.n72 VP.n0 19.1821
R219 VP.n39 VP.n11 19.1821
R220 VP.n52 VP.n51 18.1985
R221 VP.n65 VP.n64 18.1985
R222 VP.n32 VP.n31 18.1985
R223 VP.n53 VP.n52 6.39438
R224 VP.n64 VP.n63 6.39438
R225 VP.n31 VP.n30 6.39438
R226 VP.n20 VP.n19 6.39438
R227 VP.n21 VP.n18 5.6022
R228 VP.n41 VP.n40 0.354861
R229 VP.n43 VP.n42 0.354861
R230 VP.n74 VP.n73 0.354861
R231 VP VP.n74 0.267071
R232 VP.n22 VP.n21 0.189894
R233 VP.n23 VP.n22 0.189894
R234 VP.n23 VP.n16 0.189894
R235 VP.n27 VP.n16 0.189894
R236 VP.n28 VP.n27 0.189894
R237 VP.n29 VP.n28 0.189894
R238 VP.n29 VP.n14 0.189894
R239 VP.n34 VP.n14 0.189894
R240 VP.n35 VP.n34 0.189894
R241 VP.n36 VP.n35 0.189894
R242 VP.n36 VP.n12 0.189894
R243 VP.n40 VP.n12 0.189894
R244 VP.n43 VP.n9 0.189894
R245 VP.n47 VP.n9 0.189894
R246 VP.n48 VP.n47 0.189894
R247 VP.n49 VP.n48 0.189894
R248 VP.n49 VP.n7 0.189894
R249 VP.n54 VP.n7 0.189894
R250 VP.n55 VP.n54 0.189894
R251 VP.n56 VP.n55 0.189894
R252 VP.n56 VP.n5 0.189894
R253 VP.n60 VP.n5 0.189894
R254 VP.n61 VP.n60 0.189894
R255 VP.n62 VP.n61 0.189894
R256 VP.n62 VP.n3 0.189894
R257 VP.n67 VP.n3 0.189894
R258 VP.n68 VP.n67 0.189894
R259 VP.n69 VP.n68 0.189894
R260 VP.n69 VP.n1 0.189894
R261 VP.n73 VP.n1 0.189894
R262 VDD1 VDD1.n0 78.1201
R263 VDD1.n3 VDD1.n2 78.0063
R264 VDD1.n3 VDD1.n1 78.0063
R265 VDD1.n5 VDD1.n4 76.6566
R266 VDD1.n5 VDD1.n3 45.169
R267 VDD1.n4 VDD1.t4 3.40773
R268 VDD1.n4 VDD1.t2 3.40773
R269 VDD1.n0 VDD1.t7 3.40773
R270 VDD1.n0 VDD1.t6 3.40773
R271 VDD1.n2 VDD1.t3 3.40773
R272 VDD1.n2 VDD1.t0 3.40773
R273 VDD1.n1 VDD1.t1 3.40773
R274 VDD1.n1 VDD1.t5 3.40773
R275 VDD1 VDD1.n5 1.34748
R276 B.n572 B.n73 585
R277 B.n574 B.n573 585
R278 B.n575 B.n72 585
R279 B.n577 B.n576 585
R280 B.n578 B.n71 585
R281 B.n580 B.n579 585
R282 B.n581 B.n70 585
R283 B.n583 B.n582 585
R284 B.n584 B.n69 585
R285 B.n586 B.n585 585
R286 B.n587 B.n68 585
R287 B.n589 B.n588 585
R288 B.n590 B.n67 585
R289 B.n592 B.n591 585
R290 B.n593 B.n66 585
R291 B.n595 B.n594 585
R292 B.n596 B.n65 585
R293 B.n598 B.n597 585
R294 B.n599 B.n64 585
R295 B.n601 B.n600 585
R296 B.n602 B.n63 585
R297 B.n604 B.n603 585
R298 B.n605 B.n62 585
R299 B.n607 B.n606 585
R300 B.n608 B.n61 585
R301 B.n610 B.n609 585
R302 B.n611 B.n60 585
R303 B.n613 B.n612 585
R304 B.n614 B.n59 585
R305 B.n616 B.n615 585
R306 B.n617 B.n58 585
R307 B.n619 B.n618 585
R308 B.n620 B.n57 585
R309 B.n622 B.n621 585
R310 B.n624 B.n623 585
R311 B.n625 B.n53 585
R312 B.n627 B.n626 585
R313 B.n628 B.n52 585
R314 B.n630 B.n629 585
R315 B.n631 B.n51 585
R316 B.n633 B.n632 585
R317 B.n634 B.n50 585
R318 B.n636 B.n635 585
R319 B.n637 B.n47 585
R320 B.n640 B.n639 585
R321 B.n641 B.n46 585
R322 B.n643 B.n642 585
R323 B.n644 B.n45 585
R324 B.n646 B.n645 585
R325 B.n647 B.n44 585
R326 B.n649 B.n648 585
R327 B.n650 B.n43 585
R328 B.n652 B.n651 585
R329 B.n653 B.n42 585
R330 B.n655 B.n654 585
R331 B.n656 B.n41 585
R332 B.n658 B.n657 585
R333 B.n659 B.n40 585
R334 B.n661 B.n660 585
R335 B.n662 B.n39 585
R336 B.n664 B.n663 585
R337 B.n665 B.n38 585
R338 B.n667 B.n666 585
R339 B.n668 B.n37 585
R340 B.n670 B.n669 585
R341 B.n671 B.n36 585
R342 B.n673 B.n672 585
R343 B.n674 B.n35 585
R344 B.n676 B.n675 585
R345 B.n677 B.n34 585
R346 B.n679 B.n678 585
R347 B.n680 B.n33 585
R348 B.n682 B.n681 585
R349 B.n683 B.n32 585
R350 B.n685 B.n684 585
R351 B.n686 B.n31 585
R352 B.n688 B.n687 585
R353 B.n689 B.n30 585
R354 B.n571 B.n570 585
R355 B.n569 B.n74 585
R356 B.n568 B.n567 585
R357 B.n566 B.n75 585
R358 B.n565 B.n564 585
R359 B.n563 B.n76 585
R360 B.n562 B.n561 585
R361 B.n560 B.n77 585
R362 B.n559 B.n558 585
R363 B.n557 B.n78 585
R364 B.n556 B.n555 585
R365 B.n554 B.n79 585
R366 B.n553 B.n552 585
R367 B.n551 B.n80 585
R368 B.n550 B.n549 585
R369 B.n548 B.n81 585
R370 B.n547 B.n546 585
R371 B.n545 B.n82 585
R372 B.n544 B.n543 585
R373 B.n542 B.n83 585
R374 B.n541 B.n540 585
R375 B.n539 B.n84 585
R376 B.n538 B.n537 585
R377 B.n536 B.n85 585
R378 B.n535 B.n534 585
R379 B.n533 B.n86 585
R380 B.n532 B.n531 585
R381 B.n530 B.n87 585
R382 B.n529 B.n528 585
R383 B.n527 B.n88 585
R384 B.n526 B.n525 585
R385 B.n524 B.n89 585
R386 B.n523 B.n522 585
R387 B.n521 B.n90 585
R388 B.n520 B.n519 585
R389 B.n518 B.n91 585
R390 B.n517 B.n516 585
R391 B.n515 B.n92 585
R392 B.n514 B.n513 585
R393 B.n512 B.n93 585
R394 B.n511 B.n510 585
R395 B.n509 B.n94 585
R396 B.n508 B.n507 585
R397 B.n506 B.n95 585
R398 B.n505 B.n504 585
R399 B.n503 B.n96 585
R400 B.n502 B.n501 585
R401 B.n500 B.n97 585
R402 B.n499 B.n498 585
R403 B.n497 B.n98 585
R404 B.n496 B.n495 585
R405 B.n494 B.n99 585
R406 B.n493 B.n492 585
R407 B.n491 B.n100 585
R408 B.n490 B.n489 585
R409 B.n488 B.n101 585
R410 B.n487 B.n486 585
R411 B.n485 B.n102 585
R412 B.n484 B.n483 585
R413 B.n482 B.n103 585
R414 B.n481 B.n480 585
R415 B.n479 B.n104 585
R416 B.n478 B.n477 585
R417 B.n476 B.n105 585
R418 B.n475 B.n474 585
R419 B.n473 B.n106 585
R420 B.n472 B.n471 585
R421 B.n470 B.n107 585
R422 B.n469 B.n468 585
R423 B.n467 B.n108 585
R424 B.n466 B.n465 585
R425 B.n464 B.n109 585
R426 B.n463 B.n462 585
R427 B.n461 B.n110 585
R428 B.n460 B.n459 585
R429 B.n458 B.n111 585
R430 B.n457 B.n456 585
R431 B.n455 B.n112 585
R432 B.n454 B.n453 585
R433 B.n452 B.n113 585
R434 B.n451 B.n450 585
R435 B.n449 B.n114 585
R436 B.n448 B.n447 585
R437 B.n446 B.n115 585
R438 B.n445 B.n444 585
R439 B.n443 B.n116 585
R440 B.n442 B.n441 585
R441 B.n440 B.n117 585
R442 B.n439 B.n438 585
R443 B.n437 B.n118 585
R444 B.n436 B.n435 585
R445 B.n434 B.n119 585
R446 B.n433 B.n432 585
R447 B.n431 B.n120 585
R448 B.n430 B.n429 585
R449 B.n428 B.n121 585
R450 B.n427 B.n426 585
R451 B.n425 B.n122 585
R452 B.n424 B.n423 585
R453 B.n422 B.n123 585
R454 B.n421 B.n420 585
R455 B.n419 B.n124 585
R456 B.n418 B.n417 585
R457 B.n416 B.n125 585
R458 B.n415 B.n414 585
R459 B.n413 B.n126 585
R460 B.n412 B.n411 585
R461 B.n410 B.n127 585
R462 B.n409 B.n408 585
R463 B.n407 B.n128 585
R464 B.n406 B.n405 585
R465 B.n404 B.n129 585
R466 B.n403 B.n402 585
R467 B.n284 B.n173 585
R468 B.n286 B.n285 585
R469 B.n287 B.n172 585
R470 B.n289 B.n288 585
R471 B.n290 B.n171 585
R472 B.n292 B.n291 585
R473 B.n293 B.n170 585
R474 B.n295 B.n294 585
R475 B.n296 B.n169 585
R476 B.n298 B.n297 585
R477 B.n299 B.n168 585
R478 B.n301 B.n300 585
R479 B.n302 B.n167 585
R480 B.n304 B.n303 585
R481 B.n305 B.n166 585
R482 B.n307 B.n306 585
R483 B.n308 B.n165 585
R484 B.n310 B.n309 585
R485 B.n311 B.n164 585
R486 B.n313 B.n312 585
R487 B.n314 B.n163 585
R488 B.n316 B.n315 585
R489 B.n317 B.n162 585
R490 B.n319 B.n318 585
R491 B.n320 B.n161 585
R492 B.n322 B.n321 585
R493 B.n323 B.n160 585
R494 B.n325 B.n324 585
R495 B.n326 B.n159 585
R496 B.n328 B.n327 585
R497 B.n329 B.n158 585
R498 B.n331 B.n330 585
R499 B.n332 B.n157 585
R500 B.n334 B.n333 585
R501 B.n336 B.n335 585
R502 B.n337 B.n153 585
R503 B.n339 B.n338 585
R504 B.n340 B.n152 585
R505 B.n342 B.n341 585
R506 B.n343 B.n151 585
R507 B.n345 B.n344 585
R508 B.n346 B.n150 585
R509 B.n348 B.n347 585
R510 B.n349 B.n147 585
R511 B.n352 B.n351 585
R512 B.n353 B.n146 585
R513 B.n355 B.n354 585
R514 B.n356 B.n145 585
R515 B.n358 B.n357 585
R516 B.n359 B.n144 585
R517 B.n361 B.n360 585
R518 B.n362 B.n143 585
R519 B.n364 B.n363 585
R520 B.n365 B.n142 585
R521 B.n367 B.n366 585
R522 B.n368 B.n141 585
R523 B.n370 B.n369 585
R524 B.n371 B.n140 585
R525 B.n373 B.n372 585
R526 B.n374 B.n139 585
R527 B.n376 B.n375 585
R528 B.n377 B.n138 585
R529 B.n379 B.n378 585
R530 B.n380 B.n137 585
R531 B.n382 B.n381 585
R532 B.n383 B.n136 585
R533 B.n385 B.n384 585
R534 B.n386 B.n135 585
R535 B.n388 B.n387 585
R536 B.n389 B.n134 585
R537 B.n391 B.n390 585
R538 B.n392 B.n133 585
R539 B.n394 B.n393 585
R540 B.n395 B.n132 585
R541 B.n397 B.n396 585
R542 B.n398 B.n131 585
R543 B.n400 B.n399 585
R544 B.n401 B.n130 585
R545 B.n283 B.n282 585
R546 B.n281 B.n174 585
R547 B.n280 B.n279 585
R548 B.n278 B.n175 585
R549 B.n277 B.n276 585
R550 B.n275 B.n176 585
R551 B.n274 B.n273 585
R552 B.n272 B.n177 585
R553 B.n271 B.n270 585
R554 B.n269 B.n178 585
R555 B.n268 B.n267 585
R556 B.n266 B.n179 585
R557 B.n265 B.n264 585
R558 B.n263 B.n180 585
R559 B.n262 B.n261 585
R560 B.n260 B.n181 585
R561 B.n259 B.n258 585
R562 B.n257 B.n182 585
R563 B.n256 B.n255 585
R564 B.n254 B.n183 585
R565 B.n253 B.n252 585
R566 B.n251 B.n184 585
R567 B.n250 B.n249 585
R568 B.n248 B.n185 585
R569 B.n247 B.n246 585
R570 B.n245 B.n186 585
R571 B.n244 B.n243 585
R572 B.n242 B.n187 585
R573 B.n241 B.n240 585
R574 B.n239 B.n188 585
R575 B.n238 B.n237 585
R576 B.n236 B.n189 585
R577 B.n235 B.n234 585
R578 B.n233 B.n190 585
R579 B.n232 B.n231 585
R580 B.n230 B.n191 585
R581 B.n229 B.n228 585
R582 B.n227 B.n192 585
R583 B.n226 B.n225 585
R584 B.n224 B.n193 585
R585 B.n223 B.n222 585
R586 B.n221 B.n194 585
R587 B.n220 B.n219 585
R588 B.n218 B.n195 585
R589 B.n217 B.n216 585
R590 B.n215 B.n196 585
R591 B.n214 B.n213 585
R592 B.n212 B.n197 585
R593 B.n211 B.n210 585
R594 B.n209 B.n198 585
R595 B.n208 B.n207 585
R596 B.n206 B.n199 585
R597 B.n205 B.n204 585
R598 B.n203 B.n200 585
R599 B.n202 B.n201 585
R600 B.n2 B.n0 585
R601 B.n773 B.n1 585
R602 B.n772 B.n771 585
R603 B.n770 B.n3 585
R604 B.n769 B.n768 585
R605 B.n767 B.n4 585
R606 B.n766 B.n765 585
R607 B.n764 B.n5 585
R608 B.n763 B.n762 585
R609 B.n761 B.n6 585
R610 B.n760 B.n759 585
R611 B.n758 B.n7 585
R612 B.n757 B.n756 585
R613 B.n755 B.n8 585
R614 B.n754 B.n753 585
R615 B.n752 B.n9 585
R616 B.n751 B.n750 585
R617 B.n749 B.n10 585
R618 B.n748 B.n747 585
R619 B.n746 B.n11 585
R620 B.n745 B.n744 585
R621 B.n743 B.n12 585
R622 B.n742 B.n741 585
R623 B.n740 B.n13 585
R624 B.n739 B.n738 585
R625 B.n737 B.n14 585
R626 B.n736 B.n735 585
R627 B.n734 B.n15 585
R628 B.n733 B.n732 585
R629 B.n731 B.n16 585
R630 B.n730 B.n729 585
R631 B.n728 B.n17 585
R632 B.n727 B.n726 585
R633 B.n725 B.n18 585
R634 B.n724 B.n723 585
R635 B.n722 B.n19 585
R636 B.n721 B.n720 585
R637 B.n719 B.n20 585
R638 B.n718 B.n717 585
R639 B.n716 B.n21 585
R640 B.n715 B.n714 585
R641 B.n713 B.n22 585
R642 B.n712 B.n711 585
R643 B.n710 B.n23 585
R644 B.n709 B.n708 585
R645 B.n707 B.n24 585
R646 B.n706 B.n705 585
R647 B.n704 B.n25 585
R648 B.n703 B.n702 585
R649 B.n701 B.n26 585
R650 B.n700 B.n699 585
R651 B.n698 B.n27 585
R652 B.n697 B.n696 585
R653 B.n695 B.n28 585
R654 B.n694 B.n693 585
R655 B.n692 B.n29 585
R656 B.n691 B.n690 585
R657 B.n775 B.n774 585
R658 B.n282 B.n173 535.745
R659 B.n690 B.n689 535.745
R660 B.n402 B.n401 535.745
R661 B.n570 B.n73 535.745
R662 B.n148 B.t0 286.966
R663 B.n154 B.t6 286.966
R664 B.n48 B.t3 286.966
R665 B.n54 B.t9 286.966
R666 B.n148 B.t2 171.458
R667 B.n54 B.t10 171.458
R668 B.n154 B.t8 171.447
R669 B.n48 B.t4 171.447
R670 B.n282 B.n281 163.367
R671 B.n281 B.n280 163.367
R672 B.n280 B.n175 163.367
R673 B.n276 B.n175 163.367
R674 B.n276 B.n275 163.367
R675 B.n275 B.n274 163.367
R676 B.n274 B.n177 163.367
R677 B.n270 B.n177 163.367
R678 B.n270 B.n269 163.367
R679 B.n269 B.n268 163.367
R680 B.n268 B.n179 163.367
R681 B.n264 B.n179 163.367
R682 B.n264 B.n263 163.367
R683 B.n263 B.n262 163.367
R684 B.n262 B.n181 163.367
R685 B.n258 B.n181 163.367
R686 B.n258 B.n257 163.367
R687 B.n257 B.n256 163.367
R688 B.n256 B.n183 163.367
R689 B.n252 B.n183 163.367
R690 B.n252 B.n251 163.367
R691 B.n251 B.n250 163.367
R692 B.n250 B.n185 163.367
R693 B.n246 B.n185 163.367
R694 B.n246 B.n245 163.367
R695 B.n245 B.n244 163.367
R696 B.n244 B.n187 163.367
R697 B.n240 B.n187 163.367
R698 B.n240 B.n239 163.367
R699 B.n239 B.n238 163.367
R700 B.n238 B.n189 163.367
R701 B.n234 B.n189 163.367
R702 B.n234 B.n233 163.367
R703 B.n233 B.n232 163.367
R704 B.n232 B.n191 163.367
R705 B.n228 B.n191 163.367
R706 B.n228 B.n227 163.367
R707 B.n227 B.n226 163.367
R708 B.n226 B.n193 163.367
R709 B.n222 B.n193 163.367
R710 B.n222 B.n221 163.367
R711 B.n221 B.n220 163.367
R712 B.n220 B.n195 163.367
R713 B.n216 B.n195 163.367
R714 B.n216 B.n215 163.367
R715 B.n215 B.n214 163.367
R716 B.n214 B.n197 163.367
R717 B.n210 B.n197 163.367
R718 B.n210 B.n209 163.367
R719 B.n209 B.n208 163.367
R720 B.n208 B.n199 163.367
R721 B.n204 B.n199 163.367
R722 B.n204 B.n203 163.367
R723 B.n203 B.n202 163.367
R724 B.n202 B.n2 163.367
R725 B.n774 B.n2 163.367
R726 B.n774 B.n773 163.367
R727 B.n773 B.n772 163.367
R728 B.n772 B.n3 163.367
R729 B.n768 B.n3 163.367
R730 B.n768 B.n767 163.367
R731 B.n767 B.n766 163.367
R732 B.n766 B.n5 163.367
R733 B.n762 B.n5 163.367
R734 B.n762 B.n761 163.367
R735 B.n761 B.n760 163.367
R736 B.n760 B.n7 163.367
R737 B.n756 B.n7 163.367
R738 B.n756 B.n755 163.367
R739 B.n755 B.n754 163.367
R740 B.n754 B.n9 163.367
R741 B.n750 B.n9 163.367
R742 B.n750 B.n749 163.367
R743 B.n749 B.n748 163.367
R744 B.n748 B.n11 163.367
R745 B.n744 B.n11 163.367
R746 B.n744 B.n743 163.367
R747 B.n743 B.n742 163.367
R748 B.n742 B.n13 163.367
R749 B.n738 B.n13 163.367
R750 B.n738 B.n737 163.367
R751 B.n737 B.n736 163.367
R752 B.n736 B.n15 163.367
R753 B.n732 B.n15 163.367
R754 B.n732 B.n731 163.367
R755 B.n731 B.n730 163.367
R756 B.n730 B.n17 163.367
R757 B.n726 B.n17 163.367
R758 B.n726 B.n725 163.367
R759 B.n725 B.n724 163.367
R760 B.n724 B.n19 163.367
R761 B.n720 B.n19 163.367
R762 B.n720 B.n719 163.367
R763 B.n719 B.n718 163.367
R764 B.n718 B.n21 163.367
R765 B.n714 B.n21 163.367
R766 B.n714 B.n713 163.367
R767 B.n713 B.n712 163.367
R768 B.n712 B.n23 163.367
R769 B.n708 B.n23 163.367
R770 B.n708 B.n707 163.367
R771 B.n707 B.n706 163.367
R772 B.n706 B.n25 163.367
R773 B.n702 B.n25 163.367
R774 B.n702 B.n701 163.367
R775 B.n701 B.n700 163.367
R776 B.n700 B.n27 163.367
R777 B.n696 B.n27 163.367
R778 B.n696 B.n695 163.367
R779 B.n695 B.n694 163.367
R780 B.n694 B.n29 163.367
R781 B.n690 B.n29 163.367
R782 B.n286 B.n173 163.367
R783 B.n287 B.n286 163.367
R784 B.n288 B.n287 163.367
R785 B.n288 B.n171 163.367
R786 B.n292 B.n171 163.367
R787 B.n293 B.n292 163.367
R788 B.n294 B.n293 163.367
R789 B.n294 B.n169 163.367
R790 B.n298 B.n169 163.367
R791 B.n299 B.n298 163.367
R792 B.n300 B.n299 163.367
R793 B.n300 B.n167 163.367
R794 B.n304 B.n167 163.367
R795 B.n305 B.n304 163.367
R796 B.n306 B.n305 163.367
R797 B.n306 B.n165 163.367
R798 B.n310 B.n165 163.367
R799 B.n311 B.n310 163.367
R800 B.n312 B.n311 163.367
R801 B.n312 B.n163 163.367
R802 B.n316 B.n163 163.367
R803 B.n317 B.n316 163.367
R804 B.n318 B.n317 163.367
R805 B.n318 B.n161 163.367
R806 B.n322 B.n161 163.367
R807 B.n323 B.n322 163.367
R808 B.n324 B.n323 163.367
R809 B.n324 B.n159 163.367
R810 B.n328 B.n159 163.367
R811 B.n329 B.n328 163.367
R812 B.n330 B.n329 163.367
R813 B.n330 B.n157 163.367
R814 B.n334 B.n157 163.367
R815 B.n335 B.n334 163.367
R816 B.n335 B.n153 163.367
R817 B.n339 B.n153 163.367
R818 B.n340 B.n339 163.367
R819 B.n341 B.n340 163.367
R820 B.n341 B.n151 163.367
R821 B.n345 B.n151 163.367
R822 B.n346 B.n345 163.367
R823 B.n347 B.n346 163.367
R824 B.n347 B.n147 163.367
R825 B.n352 B.n147 163.367
R826 B.n353 B.n352 163.367
R827 B.n354 B.n353 163.367
R828 B.n354 B.n145 163.367
R829 B.n358 B.n145 163.367
R830 B.n359 B.n358 163.367
R831 B.n360 B.n359 163.367
R832 B.n360 B.n143 163.367
R833 B.n364 B.n143 163.367
R834 B.n365 B.n364 163.367
R835 B.n366 B.n365 163.367
R836 B.n366 B.n141 163.367
R837 B.n370 B.n141 163.367
R838 B.n371 B.n370 163.367
R839 B.n372 B.n371 163.367
R840 B.n372 B.n139 163.367
R841 B.n376 B.n139 163.367
R842 B.n377 B.n376 163.367
R843 B.n378 B.n377 163.367
R844 B.n378 B.n137 163.367
R845 B.n382 B.n137 163.367
R846 B.n383 B.n382 163.367
R847 B.n384 B.n383 163.367
R848 B.n384 B.n135 163.367
R849 B.n388 B.n135 163.367
R850 B.n389 B.n388 163.367
R851 B.n390 B.n389 163.367
R852 B.n390 B.n133 163.367
R853 B.n394 B.n133 163.367
R854 B.n395 B.n394 163.367
R855 B.n396 B.n395 163.367
R856 B.n396 B.n131 163.367
R857 B.n400 B.n131 163.367
R858 B.n401 B.n400 163.367
R859 B.n402 B.n129 163.367
R860 B.n406 B.n129 163.367
R861 B.n407 B.n406 163.367
R862 B.n408 B.n407 163.367
R863 B.n408 B.n127 163.367
R864 B.n412 B.n127 163.367
R865 B.n413 B.n412 163.367
R866 B.n414 B.n413 163.367
R867 B.n414 B.n125 163.367
R868 B.n418 B.n125 163.367
R869 B.n419 B.n418 163.367
R870 B.n420 B.n419 163.367
R871 B.n420 B.n123 163.367
R872 B.n424 B.n123 163.367
R873 B.n425 B.n424 163.367
R874 B.n426 B.n425 163.367
R875 B.n426 B.n121 163.367
R876 B.n430 B.n121 163.367
R877 B.n431 B.n430 163.367
R878 B.n432 B.n431 163.367
R879 B.n432 B.n119 163.367
R880 B.n436 B.n119 163.367
R881 B.n437 B.n436 163.367
R882 B.n438 B.n437 163.367
R883 B.n438 B.n117 163.367
R884 B.n442 B.n117 163.367
R885 B.n443 B.n442 163.367
R886 B.n444 B.n443 163.367
R887 B.n444 B.n115 163.367
R888 B.n448 B.n115 163.367
R889 B.n449 B.n448 163.367
R890 B.n450 B.n449 163.367
R891 B.n450 B.n113 163.367
R892 B.n454 B.n113 163.367
R893 B.n455 B.n454 163.367
R894 B.n456 B.n455 163.367
R895 B.n456 B.n111 163.367
R896 B.n460 B.n111 163.367
R897 B.n461 B.n460 163.367
R898 B.n462 B.n461 163.367
R899 B.n462 B.n109 163.367
R900 B.n466 B.n109 163.367
R901 B.n467 B.n466 163.367
R902 B.n468 B.n467 163.367
R903 B.n468 B.n107 163.367
R904 B.n472 B.n107 163.367
R905 B.n473 B.n472 163.367
R906 B.n474 B.n473 163.367
R907 B.n474 B.n105 163.367
R908 B.n478 B.n105 163.367
R909 B.n479 B.n478 163.367
R910 B.n480 B.n479 163.367
R911 B.n480 B.n103 163.367
R912 B.n484 B.n103 163.367
R913 B.n485 B.n484 163.367
R914 B.n486 B.n485 163.367
R915 B.n486 B.n101 163.367
R916 B.n490 B.n101 163.367
R917 B.n491 B.n490 163.367
R918 B.n492 B.n491 163.367
R919 B.n492 B.n99 163.367
R920 B.n496 B.n99 163.367
R921 B.n497 B.n496 163.367
R922 B.n498 B.n497 163.367
R923 B.n498 B.n97 163.367
R924 B.n502 B.n97 163.367
R925 B.n503 B.n502 163.367
R926 B.n504 B.n503 163.367
R927 B.n504 B.n95 163.367
R928 B.n508 B.n95 163.367
R929 B.n509 B.n508 163.367
R930 B.n510 B.n509 163.367
R931 B.n510 B.n93 163.367
R932 B.n514 B.n93 163.367
R933 B.n515 B.n514 163.367
R934 B.n516 B.n515 163.367
R935 B.n516 B.n91 163.367
R936 B.n520 B.n91 163.367
R937 B.n521 B.n520 163.367
R938 B.n522 B.n521 163.367
R939 B.n522 B.n89 163.367
R940 B.n526 B.n89 163.367
R941 B.n527 B.n526 163.367
R942 B.n528 B.n527 163.367
R943 B.n528 B.n87 163.367
R944 B.n532 B.n87 163.367
R945 B.n533 B.n532 163.367
R946 B.n534 B.n533 163.367
R947 B.n534 B.n85 163.367
R948 B.n538 B.n85 163.367
R949 B.n539 B.n538 163.367
R950 B.n540 B.n539 163.367
R951 B.n540 B.n83 163.367
R952 B.n544 B.n83 163.367
R953 B.n545 B.n544 163.367
R954 B.n546 B.n545 163.367
R955 B.n546 B.n81 163.367
R956 B.n550 B.n81 163.367
R957 B.n551 B.n550 163.367
R958 B.n552 B.n551 163.367
R959 B.n552 B.n79 163.367
R960 B.n556 B.n79 163.367
R961 B.n557 B.n556 163.367
R962 B.n558 B.n557 163.367
R963 B.n558 B.n77 163.367
R964 B.n562 B.n77 163.367
R965 B.n563 B.n562 163.367
R966 B.n564 B.n563 163.367
R967 B.n564 B.n75 163.367
R968 B.n568 B.n75 163.367
R969 B.n569 B.n568 163.367
R970 B.n570 B.n569 163.367
R971 B.n689 B.n688 163.367
R972 B.n688 B.n31 163.367
R973 B.n684 B.n31 163.367
R974 B.n684 B.n683 163.367
R975 B.n683 B.n682 163.367
R976 B.n682 B.n33 163.367
R977 B.n678 B.n33 163.367
R978 B.n678 B.n677 163.367
R979 B.n677 B.n676 163.367
R980 B.n676 B.n35 163.367
R981 B.n672 B.n35 163.367
R982 B.n672 B.n671 163.367
R983 B.n671 B.n670 163.367
R984 B.n670 B.n37 163.367
R985 B.n666 B.n37 163.367
R986 B.n666 B.n665 163.367
R987 B.n665 B.n664 163.367
R988 B.n664 B.n39 163.367
R989 B.n660 B.n39 163.367
R990 B.n660 B.n659 163.367
R991 B.n659 B.n658 163.367
R992 B.n658 B.n41 163.367
R993 B.n654 B.n41 163.367
R994 B.n654 B.n653 163.367
R995 B.n653 B.n652 163.367
R996 B.n652 B.n43 163.367
R997 B.n648 B.n43 163.367
R998 B.n648 B.n647 163.367
R999 B.n647 B.n646 163.367
R1000 B.n646 B.n45 163.367
R1001 B.n642 B.n45 163.367
R1002 B.n642 B.n641 163.367
R1003 B.n641 B.n640 163.367
R1004 B.n640 B.n47 163.367
R1005 B.n635 B.n47 163.367
R1006 B.n635 B.n634 163.367
R1007 B.n634 B.n633 163.367
R1008 B.n633 B.n51 163.367
R1009 B.n629 B.n51 163.367
R1010 B.n629 B.n628 163.367
R1011 B.n628 B.n627 163.367
R1012 B.n627 B.n53 163.367
R1013 B.n623 B.n53 163.367
R1014 B.n623 B.n622 163.367
R1015 B.n622 B.n57 163.367
R1016 B.n618 B.n57 163.367
R1017 B.n618 B.n617 163.367
R1018 B.n617 B.n616 163.367
R1019 B.n616 B.n59 163.367
R1020 B.n612 B.n59 163.367
R1021 B.n612 B.n611 163.367
R1022 B.n611 B.n610 163.367
R1023 B.n610 B.n61 163.367
R1024 B.n606 B.n61 163.367
R1025 B.n606 B.n605 163.367
R1026 B.n605 B.n604 163.367
R1027 B.n604 B.n63 163.367
R1028 B.n600 B.n63 163.367
R1029 B.n600 B.n599 163.367
R1030 B.n599 B.n598 163.367
R1031 B.n598 B.n65 163.367
R1032 B.n594 B.n65 163.367
R1033 B.n594 B.n593 163.367
R1034 B.n593 B.n592 163.367
R1035 B.n592 B.n67 163.367
R1036 B.n588 B.n67 163.367
R1037 B.n588 B.n587 163.367
R1038 B.n587 B.n586 163.367
R1039 B.n586 B.n69 163.367
R1040 B.n582 B.n69 163.367
R1041 B.n582 B.n581 163.367
R1042 B.n581 B.n580 163.367
R1043 B.n580 B.n71 163.367
R1044 B.n576 B.n71 163.367
R1045 B.n576 B.n575 163.367
R1046 B.n575 B.n574 163.367
R1047 B.n574 B.n73 163.367
R1048 B.n149 B.t1 108.234
R1049 B.n55 B.t11 108.234
R1050 B.n155 B.t7 108.224
R1051 B.n49 B.t5 108.224
R1052 B.n149 B.n148 63.2247
R1053 B.n155 B.n154 63.2247
R1054 B.n49 B.n48 63.2247
R1055 B.n55 B.n54 63.2247
R1056 B.n350 B.n149 59.5399
R1057 B.n156 B.n155 59.5399
R1058 B.n638 B.n49 59.5399
R1059 B.n56 B.n55 59.5399
R1060 B.n691 B.n30 34.8103
R1061 B.n572 B.n571 34.8103
R1062 B.n403 B.n130 34.8103
R1063 B.n284 B.n283 34.8103
R1064 B B.n775 18.0485
R1065 B.n687 B.n30 10.6151
R1066 B.n687 B.n686 10.6151
R1067 B.n686 B.n685 10.6151
R1068 B.n685 B.n32 10.6151
R1069 B.n681 B.n32 10.6151
R1070 B.n681 B.n680 10.6151
R1071 B.n680 B.n679 10.6151
R1072 B.n679 B.n34 10.6151
R1073 B.n675 B.n34 10.6151
R1074 B.n675 B.n674 10.6151
R1075 B.n674 B.n673 10.6151
R1076 B.n673 B.n36 10.6151
R1077 B.n669 B.n36 10.6151
R1078 B.n669 B.n668 10.6151
R1079 B.n668 B.n667 10.6151
R1080 B.n667 B.n38 10.6151
R1081 B.n663 B.n38 10.6151
R1082 B.n663 B.n662 10.6151
R1083 B.n662 B.n661 10.6151
R1084 B.n661 B.n40 10.6151
R1085 B.n657 B.n40 10.6151
R1086 B.n657 B.n656 10.6151
R1087 B.n656 B.n655 10.6151
R1088 B.n655 B.n42 10.6151
R1089 B.n651 B.n42 10.6151
R1090 B.n651 B.n650 10.6151
R1091 B.n650 B.n649 10.6151
R1092 B.n649 B.n44 10.6151
R1093 B.n645 B.n44 10.6151
R1094 B.n645 B.n644 10.6151
R1095 B.n644 B.n643 10.6151
R1096 B.n643 B.n46 10.6151
R1097 B.n639 B.n46 10.6151
R1098 B.n637 B.n636 10.6151
R1099 B.n636 B.n50 10.6151
R1100 B.n632 B.n50 10.6151
R1101 B.n632 B.n631 10.6151
R1102 B.n631 B.n630 10.6151
R1103 B.n630 B.n52 10.6151
R1104 B.n626 B.n52 10.6151
R1105 B.n626 B.n625 10.6151
R1106 B.n625 B.n624 10.6151
R1107 B.n621 B.n620 10.6151
R1108 B.n620 B.n619 10.6151
R1109 B.n619 B.n58 10.6151
R1110 B.n615 B.n58 10.6151
R1111 B.n615 B.n614 10.6151
R1112 B.n614 B.n613 10.6151
R1113 B.n613 B.n60 10.6151
R1114 B.n609 B.n60 10.6151
R1115 B.n609 B.n608 10.6151
R1116 B.n608 B.n607 10.6151
R1117 B.n607 B.n62 10.6151
R1118 B.n603 B.n62 10.6151
R1119 B.n603 B.n602 10.6151
R1120 B.n602 B.n601 10.6151
R1121 B.n601 B.n64 10.6151
R1122 B.n597 B.n64 10.6151
R1123 B.n597 B.n596 10.6151
R1124 B.n596 B.n595 10.6151
R1125 B.n595 B.n66 10.6151
R1126 B.n591 B.n66 10.6151
R1127 B.n591 B.n590 10.6151
R1128 B.n590 B.n589 10.6151
R1129 B.n589 B.n68 10.6151
R1130 B.n585 B.n68 10.6151
R1131 B.n585 B.n584 10.6151
R1132 B.n584 B.n583 10.6151
R1133 B.n583 B.n70 10.6151
R1134 B.n579 B.n70 10.6151
R1135 B.n579 B.n578 10.6151
R1136 B.n578 B.n577 10.6151
R1137 B.n577 B.n72 10.6151
R1138 B.n573 B.n72 10.6151
R1139 B.n573 B.n572 10.6151
R1140 B.n404 B.n403 10.6151
R1141 B.n405 B.n404 10.6151
R1142 B.n405 B.n128 10.6151
R1143 B.n409 B.n128 10.6151
R1144 B.n410 B.n409 10.6151
R1145 B.n411 B.n410 10.6151
R1146 B.n411 B.n126 10.6151
R1147 B.n415 B.n126 10.6151
R1148 B.n416 B.n415 10.6151
R1149 B.n417 B.n416 10.6151
R1150 B.n417 B.n124 10.6151
R1151 B.n421 B.n124 10.6151
R1152 B.n422 B.n421 10.6151
R1153 B.n423 B.n422 10.6151
R1154 B.n423 B.n122 10.6151
R1155 B.n427 B.n122 10.6151
R1156 B.n428 B.n427 10.6151
R1157 B.n429 B.n428 10.6151
R1158 B.n429 B.n120 10.6151
R1159 B.n433 B.n120 10.6151
R1160 B.n434 B.n433 10.6151
R1161 B.n435 B.n434 10.6151
R1162 B.n435 B.n118 10.6151
R1163 B.n439 B.n118 10.6151
R1164 B.n440 B.n439 10.6151
R1165 B.n441 B.n440 10.6151
R1166 B.n441 B.n116 10.6151
R1167 B.n445 B.n116 10.6151
R1168 B.n446 B.n445 10.6151
R1169 B.n447 B.n446 10.6151
R1170 B.n447 B.n114 10.6151
R1171 B.n451 B.n114 10.6151
R1172 B.n452 B.n451 10.6151
R1173 B.n453 B.n452 10.6151
R1174 B.n453 B.n112 10.6151
R1175 B.n457 B.n112 10.6151
R1176 B.n458 B.n457 10.6151
R1177 B.n459 B.n458 10.6151
R1178 B.n459 B.n110 10.6151
R1179 B.n463 B.n110 10.6151
R1180 B.n464 B.n463 10.6151
R1181 B.n465 B.n464 10.6151
R1182 B.n465 B.n108 10.6151
R1183 B.n469 B.n108 10.6151
R1184 B.n470 B.n469 10.6151
R1185 B.n471 B.n470 10.6151
R1186 B.n471 B.n106 10.6151
R1187 B.n475 B.n106 10.6151
R1188 B.n476 B.n475 10.6151
R1189 B.n477 B.n476 10.6151
R1190 B.n477 B.n104 10.6151
R1191 B.n481 B.n104 10.6151
R1192 B.n482 B.n481 10.6151
R1193 B.n483 B.n482 10.6151
R1194 B.n483 B.n102 10.6151
R1195 B.n487 B.n102 10.6151
R1196 B.n488 B.n487 10.6151
R1197 B.n489 B.n488 10.6151
R1198 B.n489 B.n100 10.6151
R1199 B.n493 B.n100 10.6151
R1200 B.n494 B.n493 10.6151
R1201 B.n495 B.n494 10.6151
R1202 B.n495 B.n98 10.6151
R1203 B.n499 B.n98 10.6151
R1204 B.n500 B.n499 10.6151
R1205 B.n501 B.n500 10.6151
R1206 B.n501 B.n96 10.6151
R1207 B.n505 B.n96 10.6151
R1208 B.n506 B.n505 10.6151
R1209 B.n507 B.n506 10.6151
R1210 B.n507 B.n94 10.6151
R1211 B.n511 B.n94 10.6151
R1212 B.n512 B.n511 10.6151
R1213 B.n513 B.n512 10.6151
R1214 B.n513 B.n92 10.6151
R1215 B.n517 B.n92 10.6151
R1216 B.n518 B.n517 10.6151
R1217 B.n519 B.n518 10.6151
R1218 B.n519 B.n90 10.6151
R1219 B.n523 B.n90 10.6151
R1220 B.n524 B.n523 10.6151
R1221 B.n525 B.n524 10.6151
R1222 B.n525 B.n88 10.6151
R1223 B.n529 B.n88 10.6151
R1224 B.n530 B.n529 10.6151
R1225 B.n531 B.n530 10.6151
R1226 B.n531 B.n86 10.6151
R1227 B.n535 B.n86 10.6151
R1228 B.n536 B.n535 10.6151
R1229 B.n537 B.n536 10.6151
R1230 B.n537 B.n84 10.6151
R1231 B.n541 B.n84 10.6151
R1232 B.n542 B.n541 10.6151
R1233 B.n543 B.n542 10.6151
R1234 B.n543 B.n82 10.6151
R1235 B.n547 B.n82 10.6151
R1236 B.n548 B.n547 10.6151
R1237 B.n549 B.n548 10.6151
R1238 B.n549 B.n80 10.6151
R1239 B.n553 B.n80 10.6151
R1240 B.n554 B.n553 10.6151
R1241 B.n555 B.n554 10.6151
R1242 B.n555 B.n78 10.6151
R1243 B.n559 B.n78 10.6151
R1244 B.n560 B.n559 10.6151
R1245 B.n561 B.n560 10.6151
R1246 B.n561 B.n76 10.6151
R1247 B.n565 B.n76 10.6151
R1248 B.n566 B.n565 10.6151
R1249 B.n567 B.n566 10.6151
R1250 B.n567 B.n74 10.6151
R1251 B.n571 B.n74 10.6151
R1252 B.n285 B.n284 10.6151
R1253 B.n285 B.n172 10.6151
R1254 B.n289 B.n172 10.6151
R1255 B.n290 B.n289 10.6151
R1256 B.n291 B.n290 10.6151
R1257 B.n291 B.n170 10.6151
R1258 B.n295 B.n170 10.6151
R1259 B.n296 B.n295 10.6151
R1260 B.n297 B.n296 10.6151
R1261 B.n297 B.n168 10.6151
R1262 B.n301 B.n168 10.6151
R1263 B.n302 B.n301 10.6151
R1264 B.n303 B.n302 10.6151
R1265 B.n303 B.n166 10.6151
R1266 B.n307 B.n166 10.6151
R1267 B.n308 B.n307 10.6151
R1268 B.n309 B.n308 10.6151
R1269 B.n309 B.n164 10.6151
R1270 B.n313 B.n164 10.6151
R1271 B.n314 B.n313 10.6151
R1272 B.n315 B.n314 10.6151
R1273 B.n315 B.n162 10.6151
R1274 B.n319 B.n162 10.6151
R1275 B.n320 B.n319 10.6151
R1276 B.n321 B.n320 10.6151
R1277 B.n321 B.n160 10.6151
R1278 B.n325 B.n160 10.6151
R1279 B.n326 B.n325 10.6151
R1280 B.n327 B.n326 10.6151
R1281 B.n327 B.n158 10.6151
R1282 B.n331 B.n158 10.6151
R1283 B.n332 B.n331 10.6151
R1284 B.n333 B.n332 10.6151
R1285 B.n337 B.n336 10.6151
R1286 B.n338 B.n337 10.6151
R1287 B.n338 B.n152 10.6151
R1288 B.n342 B.n152 10.6151
R1289 B.n343 B.n342 10.6151
R1290 B.n344 B.n343 10.6151
R1291 B.n344 B.n150 10.6151
R1292 B.n348 B.n150 10.6151
R1293 B.n349 B.n348 10.6151
R1294 B.n351 B.n146 10.6151
R1295 B.n355 B.n146 10.6151
R1296 B.n356 B.n355 10.6151
R1297 B.n357 B.n356 10.6151
R1298 B.n357 B.n144 10.6151
R1299 B.n361 B.n144 10.6151
R1300 B.n362 B.n361 10.6151
R1301 B.n363 B.n362 10.6151
R1302 B.n363 B.n142 10.6151
R1303 B.n367 B.n142 10.6151
R1304 B.n368 B.n367 10.6151
R1305 B.n369 B.n368 10.6151
R1306 B.n369 B.n140 10.6151
R1307 B.n373 B.n140 10.6151
R1308 B.n374 B.n373 10.6151
R1309 B.n375 B.n374 10.6151
R1310 B.n375 B.n138 10.6151
R1311 B.n379 B.n138 10.6151
R1312 B.n380 B.n379 10.6151
R1313 B.n381 B.n380 10.6151
R1314 B.n381 B.n136 10.6151
R1315 B.n385 B.n136 10.6151
R1316 B.n386 B.n385 10.6151
R1317 B.n387 B.n386 10.6151
R1318 B.n387 B.n134 10.6151
R1319 B.n391 B.n134 10.6151
R1320 B.n392 B.n391 10.6151
R1321 B.n393 B.n392 10.6151
R1322 B.n393 B.n132 10.6151
R1323 B.n397 B.n132 10.6151
R1324 B.n398 B.n397 10.6151
R1325 B.n399 B.n398 10.6151
R1326 B.n399 B.n130 10.6151
R1327 B.n283 B.n174 10.6151
R1328 B.n279 B.n174 10.6151
R1329 B.n279 B.n278 10.6151
R1330 B.n278 B.n277 10.6151
R1331 B.n277 B.n176 10.6151
R1332 B.n273 B.n176 10.6151
R1333 B.n273 B.n272 10.6151
R1334 B.n272 B.n271 10.6151
R1335 B.n271 B.n178 10.6151
R1336 B.n267 B.n178 10.6151
R1337 B.n267 B.n266 10.6151
R1338 B.n266 B.n265 10.6151
R1339 B.n265 B.n180 10.6151
R1340 B.n261 B.n180 10.6151
R1341 B.n261 B.n260 10.6151
R1342 B.n260 B.n259 10.6151
R1343 B.n259 B.n182 10.6151
R1344 B.n255 B.n182 10.6151
R1345 B.n255 B.n254 10.6151
R1346 B.n254 B.n253 10.6151
R1347 B.n253 B.n184 10.6151
R1348 B.n249 B.n184 10.6151
R1349 B.n249 B.n248 10.6151
R1350 B.n248 B.n247 10.6151
R1351 B.n247 B.n186 10.6151
R1352 B.n243 B.n186 10.6151
R1353 B.n243 B.n242 10.6151
R1354 B.n242 B.n241 10.6151
R1355 B.n241 B.n188 10.6151
R1356 B.n237 B.n188 10.6151
R1357 B.n237 B.n236 10.6151
R1358 B.n236 B.n235 10.6151
R1359 B.n235 B.n190 10.6151
R1360 B.n231 B.n190 10.6151
R1361 B.n231 B.n230 10.6151
R1362 B.n230 B.n229 10.6151
R1363 B.n229 B.n192 10.6151
R1364 B.n225 B.n192 10.6151
R1365 B.n225 B.n224 10.6151
R1366 B.n224 B.n223 10.6151
R1367 B.n223 B.n194 10.6151
R1368 B.n219 B.n194 10.6151
R1369 B.n219 B.n218 10.6151
R1370 B.n218 B.n217 10.6151
R1371 B.n217 B.n196 10.6151
R1372 B.n213 B.n196 10.6151
R1373 B.n213 B.n212 10.6151
R1374 B.n212 B.n211 10.6151
R1375 B.n211 B.n198 10.6151
R1376 B.n207 B.n198 10.6151
R1377 B.n207 B.n206 10.6151
R1378 B.n206 B.n205 10.6151
R1379 B.n205 B.n200 10.6151
R1380 B.n201 B.n200 10.6151
R1381 B.n201 B.n0 10.6151
R1382 B.n771 B.n1 10.6151
R1383 B.n771 B.n770 10.6151
R1384 B.n770 B.n769 10.6151
R1385 B.n769 B.n4 10.6151
R1386 B.n765 B.n4 10.6151
R1387 B.n765 B.n764 10.6151
R1388 B.n764 B.n763 10.6151
R1389 B.n763 B.n6 10.6151
R1390 B.n759 B.n6 10.6151
R1391 B.n759 B.n758 10.6151
R1392 B.n758 B.n757 10.6151
R1393 B.n757 B.n8 10.6151
R1394 B.n753 B.n8 10.6151
R1395 B.n753 B.n752 10.6151
R1396 B.n752 B.n751 10.6151
R1397 B.n751 B.n10 10.6151
R1398 B.n747 B.n10 10.6151
R1399 B.n747 B.n746 10.6151
R1400 B.n746 B.n745 10.6151
R1401 B.n745 B.n12 10.6151
R1402 B.n741 B.n12 10.6151
R1403 B.n741 B.n740 10.6151
R1404 B.n740 B.n739 10.6151
R1405 B.n739 B.n14 10.6151
R1406 B.n735 B.n14 10.6151
R1407 B.n735 B.n734 10.6151
R1408 B.n734 B.n733 10.6151
R1409 B.n733 B.n16 10.6151
R1410 B.n729 B.n16 10.6151
R1411 B.n729 B.n728 10.6151
R1412 B.n728 B.n727 10.6151
R1413 B.n727 B.n18 10.6151
R1414 B.n723 B.n18 10.6151
R1415 B.n723 B.n722 10.6151
R1416 B.n722 B.n721 10.6151
R1417 B.n721 B.n20 10.6151
R1418 B.n717 B.n20 10.6151
R1419 B.n717 B.n716 10.6151
R1420 B.n716 B.n715 10.6151
R1421 B.n715 B.n22 10.6151
R1422 B.n711 B.n22 10.6151
R1423 B.n711 B.n710 10.6151
R1424 B.n710 B.n709 10.6151
R1425 B.n709 B.n24 10.6151
R1426 B.n705 B.n24 10.6151
R1427 B.n705 B.n704 10.6151
R1428 B.n704 B.n703 10.6151
R1429 B.n703 B.n26 10.6151
R1430 B.n699 B.n26 10.6151
R1431 B.n699 B.n698 10.6151
R1432 B.n698 B.n697 10.6151
R1433 B.n697 B.n28 10.6151
R1434 B.n693 B.n28 10.6151
R1435 B.n693 B.n692 10.6151
R1436 B.n692 B.n691 10.6151
R1437 B.n639 B.n638 9.36635
R1438 B.n621 B.n56 9.36635
R1439 B.n333 B.n156 9.36635
R1440 B.n351 B.n350 9.36635
R1441 B.n775 B.n0 2.81026
R1442 B.n775 B.n1 2.81026
R1443 B.n638 B.n637 1.24928
R1444 B.n624 B.n56 1.24928
R1445 B.n336 B.n156 1.24928
R1446 B.n350 B.n349 1.24928
C0 VDD1 B 1.68309f
C1 B VP 2.20111f
C2 w_n4230_n2876# VDD2 2.12651f
C3 VDD1 VTAIL 7.39086f
C4 VTAIL VP 7.798299f
C5 VDD1 VN 0.152774f
C6 VN VP 7.60816f
C7 B w_n4230_n2876# 9.93134f
C8 VTAIL w_n4230_n2876# 3.68363f
C9 w_n4230_n2876# VN 8.65261f
C10 B VDD2 1.7895f
C11 VTAIL VDD2 7.447491f
C12 VDD1 VP 7.55566f
C13 VN VDD2 7.154759f
C14 B VTAIL 4.30706f
C15 VDD1 w_n4230_n2876# 1.99796f
C16 w_n4230_n2876# VP 9.20272f
C17 B VN 1.27717f
C18 VTAIL VN 7.78419f
C19 VDD1 VDD2 1.9501f
C20 VDD2 VP 0.555236f
C21 VDD2 VSUBS 1.929609f
C22 VDD1 VSUBS 2.50709f
C23 VTAIL VSUBS 1.290141f
C24 VN VSUBS 7.13358f
C25 VP VSUBS 3.848366f
C26 B VSUBS 5.165455f
C27 w_n4230_n2876# VSUBS 0.150402p
C28 B.n0 VSUBS 0.005084f
C29 B.n1 VSUBS 0.005084f
C30 B.n2 VSUBS 0.008039f
C31 B.n3 VSUBS 0.008039f
C32 B.n4 VSUBS 0.008039f
C33 B.n5 VSUBS 0.008039f
C34 B.n6 VSUBS 0.008039f
C35 B.n7 VSUBS 0.008039f
C36 B.n8 VSUBS 0.008039f
C37 B.n9 VSUBS 0.008039f
C38 B.n10 VSUBS 0.008039f
C39 B.n11 VSUBS 0.008039f
C40 B.n12 VSUBS 0.008039f
C41 B.n13 VSUBS 0.008039f
C42 B.n14 VSUBS 0.008039f
C43 B.n15 VSUBS 0.008039f
C44 B.n16 VSUBS 0.008039f
C45 B.n17 VSUBS 0.008039f
C46 B.n18 VSUBS 0.008039f
C47 B.n19 VSUBS 0.008039f
C48 B.n20 VSUBS 0.008039f
C49 B.n21 VSUBS 0.008039f
C50 B.n22 VSUBS 0.008039f
C51 B.n23 VSUBS 0.008039f
C52 B.n24 VSUBS 0.008039f
C53 B.n25 VSUBS 0.008039f
C54 B.n26 VSUBS 0.008039f
C55 B.n27 VSUBS 0.008039f
C56 B.n28 VSUBS 0.008039f
C57 B.n29 VSUBS 0.008039f
C58 B.n30 VSUBS 0.019963f
C59 B.n31 VSUBS 0.008039f
C60 B.n32 VSUBS 0.008039f
C61 B.n33 VSUBS 0.008039f
C62 B.n34 VSUBS 0.008039f
C63 B.n35 VSUBS 0.008039f
C64 B.n36 VSUBS 0.008039f
C65 B.n37 VSUBS 0.008039f
C66 B.n38 VSUBS 0.008039f
C67 B.n39 VSUBS 0.008039f
C68 B.n40 VSUBS 0.008039f
C69 B.n41 VSUBS 0.008039f
C70 B.n42 VSUBS 0.008039f
C71 B.n43 VSUBS 0.008039f
C72 B.n44 VSUBS 0.008039f
C73 B.n45 VSUBS 0.008039f
C74 B.n46 VSUBS 0.008039f
C75 B.n47 VSUBS 0.008039f
C76 B.t5 VSUBS 0.347232f
C77 B.t4 VSUBS 0.373899f
C78 B.t3 VSUBS 1.49304f
C79 B.n48 VSUBS 0.201956f
C80 B.n49 VSUBS 0.083779f
C81 B.n50 VSUBS 0.008039f
C82 B.n51 VSUBS 0.008039f
C83 B.n52 VSUBS 0.008039f
C84 B.n53 VSUBS 0.008039f
C85 B.t11 VSUBS 0.347228f
C86 B.t10 VSUBS 0.373894f
C87 B.t9 VSUBS 1.49304f
C88 B.n54 VSUBS 0.201961f
C89 B.n55 VSUBS 0.083783f
C90 B.n56 VSUBS 0.018626f
C91 B.n57 VSUBS 0.008039f
C92 B.n58 VSUBS 0.008039f
C93 B.n59 VSUBS 0.008039f
C94 B.n60 VSUBS 0.008039f
C95 B.n61 VSUBS 0.008039f
C96 B.n62 VSUBS 0.008039f
C97 B.n63 VSUBS 0.008039f
C98 B.n64 VSUBS 0.008039f
C99 B.n65 VSUBS 0.008039f
C100 B.n66 VSUBS 0.008039f
C101 B.n67 VSUBS 0.008039f
C102 B.n68 VSUBS 0.008039f
C103 B.n69 VSUBS 0.008039f
C104 B.n70 VSUBS 0.008039f
C105 B.n71 VSUBS 0.008039f
C106 B.n72 VSUBS 0.008039f
C107 B.n73 VSUBS 0.019963f
C108 B.n74 VSUBS 0.008039f
C109 B.n75 VSUBS 0.008039f
C110 B.n76 VSUBS 0.008039f
C111 B.n77 VSUBS 0.008039f
C112 B.n78 VSUBS 0.008039f
C113 B.n79 VSUBS 0.008039f
C114 B.n80 VSUBS 0.008039f
C115 B.n81 VSUBS 0.008039f
C116 B.n82 VSUBS 0.008039f
C117 B.n83 VSUBS 0.008039f
C118 B.n84 VSUBS 0.008039f
C119 B.n85 VSUBS 0.008039f
C120 B.n86 VSUBS 0.008039f
C121 B.n87 VSUBS 0.008039f
C122 B.n88 VSUBS 0.008039f
C123 B.n89 VSUBS 0.008039f
C124 B.n90 VSUBS 0.008039f
C125 B.n91 VSUBS 0.008039f
C126 B.n92 VSUBS 0.008039f
C127 B.n93 VSUBS 0.008039f
C128 B.n94 VSUBS 0.008039f
C129 B.n95 VSUBS 0.008039f
C130 B.n96 VSUBS 0.008039f
C131 B.n97 VSUBS 0.008039f
C132 B.n98 VSUBS 0.008039f
C133 B.n99 VSUBS 0.008039f
C134 B.n100 VSUBS 0.008039f
C135 B.n101 VSUBS 0.008039f
C136 B.n102 VSUBS 0.008039f
C137 B.n103 VSUBS 0.008039f
C138 B.n104 VSUBS 0.008039f
C139 B.n105 VSUBS 0.008039f
C140 B.n106 VSUBS 0.008039f
C141 B.n107 VSUBS 0.008039f
C142 B.n108 VSUBS 0.008039f
C143 B.n109 VSUBS 0.008039f
C144 B.n110 VSUBS 0.008039f
C145 B.n111 VSUBS 0.008039f
C146 B.n112 VSUBS 0.008039f
C147 B.n113 VSUBS 0.008039f
C148 B.n114 VSUBS 0.008039f
C149 B.n115 VSUBS 0.008039f
C150 B.n116 VSUBS 0.008039f
C151 B.n117 VSUBS 0.008039f
C152 B.n118 VSUBS 0.008039f
C153 B.n119 VSUBS 0.008039f
C154 B.n120 VSUBS 0.008039f
C155 B.n121 VSUBS 0.008039f
C156 B.n122 VSUBS 0.008039f
C157 B.n123 VSUBS 0.008039f
C158 B.n124 VSUBS 0.008039f
C159 B.n125 VSUBS 0.008039f
C160 B.n126 VSUBS 0.008039f
C161 B.n127 VSUBS 0.008039f
C162 B.n128 VSUBS 0.008039f
C163 B.n129 VSUBS 0.008039f
C164 B.n130 VSUBS 0.019963f
C165 B.n131 VSUBS 0.008039f
C166 B.n132 VSUBS 0.008039f
C167 B.n133 VSUBS 0.008039f
C168 B.n134 VSUBS 0.008039f
C169 B.n135 VSUBS 0.008039f
C170 B.n136 VSUBS 0.008039f
C171 B.n137 VSUBS 0.008039f
C172 B.n138 VSUBS 0.008039f
C173 B.n139 VSUBS 0.008039f
C174 B.n140 VSUBS 0.008039f
C175 B.n141 VSUBS 0.008039f
C176 B.n142 VSUBS 0.008039f
C177 B.n143 VSUBS 0.008039f
C178 B.n144 VSUBS 0.008039f
C179 B.n145 VSUBS 0.008039f
C180 B.n146 VSUBS 0.008039f
C181 B.n147 VSUBS 0.008039f
C182 B.t1 VSUBS 0.347228f
C183 B.t2 VSUBS 0.373894f
C184 B.t0 VSUBS 1.49304f
C185 B.n148 VSUBS 0.201961f
C186 B.n149 VSUBS 0.083783f
C187 B.n150 VSUBS 0.008039f
C188 B.n151 VSUBS 0.008039f
C189 B.n152 VSUBS 0.008039f
C190 B.n153 VSUBS 0.008039f
C191 B.t7 VSUBS 0.347232f
C192 B.t8 VSUBS 0.373899f
C193 B.t6 VSUBS 1.49304f
C194 B.n154 VSUBS 0.201956f
C195 B.n155 VSUBS 0.083779f
C196 B.n156 VSUBS 0.018626f
C197 B.n157 VSUBS 0.008039f
C198 B.n158 VSUBS 0.008039f
C199 B.n159 VSUBS 0.008039f
C200 B.n160 VSUBS 0.008039f
C201 B.n161 VSUBS 0.008039f
C202 B.n162 VSUBS 0.008039f
C203 B.n163 VSUBS 0.008039f
C204 B.n164 VSUBS 0.008039f
C205 B.n165 VSUBS 0.008039f
C206 B.n166 VSUBS 0.008039f
C207 B.n167 VSUBS 0.008039f
C208 B.n168 VSUBS 0.008039f
C209 B.n169 VSUBS 0.008039f
C210 B.n170 VSUBS 0.008039f
C211 B.n171 VSUBS 0.008039f
C212 B.n172 VSUBS 0.008039f
C213 B.n173 VSUBS 0.019963f
C214 B.n174 VSUBS 0.008039f
C215 B.n175 VSUBS 0.008039f
C216 B.n176 VSUBS 0.008039f
C217 B.n177 VSUBS 0.008039f
C218 B.n178 VSUBS 0.008039f
C219 B.n179 VSUBS 0.008039f
C220 B.n180 VSUBS 0.008039f
C221 B.n181 VSUBS 0.008039f
C222 B.n182 VSUBS 0.008039f
C223 B.n183 VSUBS 0.008039f
C224 B.n184 VSUBS 0.008039f
C225 B.n185 VSUBS 0.008039f
C226 B.n186 VSUBS 0.008039f
C227 B.n187 VSUBS 0.008039f
C228 B.n188 VSUBS 0.008039f
C229 B.n189 VSUBS 0.008039f
C230 B.n190 VSUBS 0.008039f
C231 B.n191 VSUBS 0.008039f
C232 B.n192 VSUBS 0.008039f
C233 B.n193 VSUBS 0.008039f
C234 B.n194 VSUBS 0.008039f
C235 B.n195 VSUBS 0.008039f
C236 B.n196 VSUBS 0.008039f
C237 B.n197 VSUBS 0.008039f
C238 B.n198 VSUBS 0.008039f
C239 B.n199 VSUBS 0.008039f
C240 B.n200 VSUBS 0.008039f
C241 B.n201 VSUBS 0.008039f
C242 B.n202 VSUBS 0.008039f
C243 B.n203 VSUBS 0.008039f
C244 B.n204 VSUBS 0.008039f
C245 B.n205 VSUBS 0.008039f
C246 B.n206 VSUBS 0.008039f
C247 B.n207 VSUBS 0.008039f
C248 B.n208 VSUBS 0.008039f
C249 B.n209 VSUBS 0.008039f
C250 B.n210 VSUBS 0.008039f
C251 B.n211 VSUBS 0.008039f
C252 B.n212 VSUBS 0.008039f
C253 B.n213 VSUBS 0.008039f
C254 B.n214 VSUBS 0.008039f
C255 B.n215 VSUBS 0.008039f
C256 B.n216 VSUBS 0.008039f
C257 B.n217 VSUBS 0.008039f
C258 B.n218 VSUBS 0.008039f
C259 B.n219 VSUBS 0.008039f
C260 B.n220 VSUBS 0.008039f
C261 B.n221 VSUBS 0.008039f
C262 B.n222 VSUBS 0.008039f
C263 B.n223 VSUBS 0.008039f
C264 B.n224 VSUBS 0.008039f
C265 B.n225 VSUBS 0.008039f
C266 B.n226 VSUBS 0.008039f
C267 B.n227 VSUBS 0.008039f
C268 B.n228 VSUBS 0.008039f
C269 B.n229 VSUBS 0.008039f
C270 B.n230 VSUBS 0.008039f
C271 B.n231 VSUBS 0.008039f
C272 B.n232 VSUBS 0.008039f
C273 B.n233 VSUBS 0.008039f
C274 B.n234 VSUBS 0.008039f
C275 B.n235 VSUBS 0.008039f
C276 B.n236 VSUBS 0.008039f
C277 B.n237 VSUBS 0.008039f
C278 B.n238 VSUBS 0.008039f
C279 B.n239 VSUBS 0.008039f
C280 B.n240 VSUBS 0.008039f
C281 B.n241 VSUBS 0.008039f
C282 B.n242 VSUBS 0.008039f
C283 B.n243 VSUBS 0.008039f
C284 B.n244 VSUBS 0.008039f
C285 B.n245 VSUBS 0.008039f
C286 B.n246 VSUBS 0.008039f
C287 B.n247 VSUBS 0.008039f
C288 B.n248 VSUBS 0.008039f
C289 B.n249 VSUBS 0.008039f
C290 B.n250 VSUBS 0.008039f
C291 B.n251 VSUBS 0.008039f
C292 B.n252 VSUBS 0.008039f
C293 B.n253 VSUBS 0.008039f
C294 B.n254 VSUBS 0.008039f
C295 B.n255 VSUBS 0.008039f
C296 B.n256 VSUBS 0.008039f
C297 B.n257 VSUBS 0.008039f
C298 B.n258 VSUBS 0.008039f
C299 B.n259 VSUBS 0.008039f
C300 B.n260 VSUBS 0.008039f
C301 B.n261 VSUBS 0.008039f
C302 B.n262 VSUBS 0.008039f
C303 B.n263 VSUBS 0.008039f
C304 B.n264 VSUBS 0.008039f
C305 B.n265 VSUBS 0.008039f
C306 B.n266 VSUBS 0.008039f
C307 B.n267 VSUBS 0.008039f
C308 B.n268 VSUBS 0.008039f
C309 B.n269 VSUBS 0.008039f
C310 B.n270 VSUBS 0.008039f
C311 B.n271 VSUBS 0.008039f
C312 B.n272 VSUBS 0.008039f
C313 B.n273 VSUBS 0.008039f
C314 B.n274 VSUBS 0.008039f
C315 B.n275 VSUBS 0.008039f
C316 B.n276 VSUBS 0.008039f
C317 B.n277 VSUBS 0.008039f
C318 B.n278 VSUBS 0.008039f
C319 B.n279 VSUBS 0.008039f
C320 B.n280 VSUBS 0.008039f
C321 B.n281 VSUBS 0.008039f
C322 B.n282 VSUBS 0.019289f
C323 B.n283 VSUBS 0.019289f
C324 B.n284 VSUBS 0.019963f
C325 B.n285 VSUBS 0.008039f
C326 B.n286 VSUBS 0.008039f
C327 B.n287 VSUBS 0.008039f
C328 B.n288 VSUBS 0.008039f
C329 B.n289 VSUBS 0.008039f
C330 B.n290 VSUBS 0.008039f
C331 B.n291 VSUBS 0.008039f
C332 B.n292 VSUBS 0.008039f
C333 B.n293 VSUBS 0.008039f
C334 B.n294 VSUBS 0.008039f
C335 B.n295 VSUBS 0.008039f
C336 B.n296 VSUBS 0.008039f
C337 B.n297 VSUBS 0.008039f
C338 B.n298 VSUBS 0.008039f
C339 B.n299 VSUBS 0.008039f
C340 B.n300 VSUBS 0.008039f
C341 B.n301 VSUBS 0.008039f
C342 B.n302 VSUBS 0.008039f
C343 B.n303 VSUBS 0.008039f
C344 B.n304 VSUBS 0.008039f
C345 B.n305 VSUBS 0.008039f
C346 B.n306 VSUBS 0.008039f
C347 B.n307 VSUBS 0.008039f
C348 B.n308 VSUBS 0.008039f
C349 B.n309 VSUBS 0.008039f
C350 B.n310 VSUBS 0.008039f
C351 B.n311 VSUBS 0.008039f
C352 B.n312 VSUBS 0.008039f
C353 B.n313 VSUBS 0.008039f
C354 B.n314 VSUBS 0.008039f
C355 B.n315 VSUBS 0.008039f
C356 B.n316 VSUBS 0.008039f
C357 B.n317 VSUBS 0.008039f
C358 B.n318 VSUBS 0.008039f
C359 B.n319 VSUBS 0.008039f
C360 B.n320 VSUBS 0.008039f
C361 B.n321 VSUBS 0.008039f
C362 B.n322 VSUBS 0.008039f
C363 B.n323 VSUBS 0.008039f
C364 B.n324 VSUBS 0.008039f
C365 B.n325 VSUBS 0.008039f
C366 B.n326 VSUBS 0.008039f
C367 B.n327 VSUBS 0.008039f
C368 B.n328 VSUBS 0.008039f
C369 B.n329 VSUBS 0.008039f
C370 B.n330 VSUBS 0.008039f
C371 B.n331 VSUBS 0.008039f
C372 B.n332 VSUBS 0.008039f
C373 B.n333 VSUBS 0.007567f
C374 B.n334 VSUBS 0.008039f
C375 B.n335 VSUBS 0.008039f
C376 B.n336 VSUBS 0.004493f
C377 B.n337 VSUBS 0.008039f
C378 B.n338 VSUBS 0.008039f
C379 B.n339 VSUBS 0.008039f
C380 B.n340 VSUBS 0.008039f
C381 B.n341 VSUBS 0.008039f
C382 B.n342 VSUBS 0.008039f
C383 B.n343 VSUBS 0.008039f
C384 B.n344 VSUBS 0.008039f
C385 B.n345 VSUBS 0.008039f
C386 B.n346 VSUBS 0.008039f
C387 B.n347 VSUBS 0.008039f
C388 B.n348 VSUBS 0.008039f
C389 B.n349 VSUBS 0.004493f
C390 B.n350 VSUBS 0.018626f
C391 B.n351 VSUBS 0.007567f
C392 B.n352 VSUBS 0.008039f
C393 B.n353 VSUBS 0.008039f
C394 B.n354 VSUBS 0.008039f
C395 B.n355 VSUBS 0.008039f
C396 B.n356 VSUBS 0.008039f
C397 B.n357 VSUBS 0.008039f
C398 B.n358 VSUBS 0.008039f
C399 B.n359 VSUBS 0.008039f
C400 B.n360 VSUBS 0.008039f
C401 B.n361 VSUBS 0.008039f
C402 B.n362 VSUBS 0.008039f
C403 B.n363 VSUBS 0.008039f
C404 B.n364 VSUBS 0.008039f
C405 B.n365 VSUBS 0.008039f
C406 B.n366 VSUBS 0.008039f
C407 B.n367 VSUBS 0.008039f
C408 B.n368 VSUBS 0.008039f
C409 B.n369 VSUBS 0.008039f
C410 B.n370 VSUBS 0.008039f
C411 B.n371 VSUBS 0.008039f
C412 B.n372 VSUBS 0.008039f
C413 B.n373 VSUBS 0.008039f
C414 B.n374 VSUBS 0.008039f
C415 B.n375 VSUBS 0.008039f
C416 B.n376 VSUBS 0.008039f
C417 B.n377 VSUBS 0.008039f
C418 B.n378 VSUBS 0.008039f
C419 B.n379 VSUBS 0.008039f
C420 B.n380 VSUBS 0.008039f
C421 B.n381 VSUBS 0.008039f
C422 B.n382 VSUBS 0.008039f
C423 B.n383 VSUBS 0.008039f
C424 B.n384 VSUBS 0.008039f
C425 B.n385 VSUBS 0.008039f
C426 B.n386 VSUBS 0.008039f
C427 B.n387 VSUBS 0.008039f
C428 B.n388 VSUBS 0.008039f
C429 B.n389 VSUBS 0.008039f
C430 B.n390 VSUBS 0.008039f
C431 B.n391 VSUBS 0.008039f
C432 B.n392 VSUBS 0.008039f
C433 B.n393 VSUBS 0.008039f
C434 B.n394 VSUBS 0.008039f
C435 B.n395 VSUBS 0.008039f
C436 B.n396 VSUBS 0.008039f
C437 B.n397 VSUBS 0.008039f
C438 B.n398 VSUBS 0.008039f
C439 B.n399 VSUBS 0.008039f
C440 B.n400 VSUBS 0.008039f
C441 B.n401 VSUBS 0.019963f
C442 B.n402 VSUBS 0.019289f
C443 B.n403 VSUBS 0.019289f
C444 B.n404 VSUBS 0.008039f
C445 B.n405 VSUBS 0.008039f
C446 B.n406 VSUBS 0.008039f
C447 B.n407 VSUBS 0.008039f
C448 B.n408 VSUBS 0.008039f
C449 B.n409 VSUBS 0.008039f
C450 B.n410 VSUBS 0.008039f
C451 B.n411 VSUBS 0.008039f
C452 B.n412 VSUBS 0.008039f
C453 B.n413 VSUBS 0.008039f
C454 B.n414 VSUBS 0.008039f
C455 B.n415 VSUBS 0.008039f
C456 B.n416 VSUBS 0.008039f
C457 B.n417 VSUBS 0.008039f
C458 B.n418 VSUBS 0.008039f
C459 B.n419 VSUBS 0.008039f
C460 B.n420 VSUBS 0.008039f
C461 B.n421 VSUBS 0.008039f
C462 B.n422 VSUBS 0.008039f
C463 B.n423 VSUBS 0.008039f
C464 B.n424 VSUBS 0.008039f
C465 B.n425 VSUBS 0.008039f
C466 B.n426 VSUBS 0.008039f
C467 B.n427 VSUBS 0.008039f
C468 B.n428 VSUBS 0.008039f
C469 B.n429 VSUBS 0.008039f
C470 B.n430 VSUBS 0.008039f
C471 B.n431 VSUBS 0.008039f
C472 B.n432 VSUBS 0.008039f
C473 B.n433 VSUBS 0.008039f
C474 B.n434 VSUBS 0.008039f
C475 B.n435 VSUBS 0.008039f
C476 B.n436 VSUBS 0.008039f
C477 B.n437 VSUBS 0.008039f
C478 B.n438 VSUBS 0.008039f
C479 B.n439 VSUBS 0.008039f
C480 B.n440 VSUBS 0.008039f
C481 B.n441 VSUBS 0.008039f
C482 B.n442 VSUBS 0.008039f
C483 B.n443 VSUBS 0.008039f
C484 B.n444 VSUBS 0.008039f
C485 B.n445 VSUBS 0.008039f
C486 B.n446 VSUBS 0.008039f
C487 B.n447 VSUBS 0.008039f
C488 B.n448 VSUBS 0.008039f
C489 B.n449 VSUBS 0.008039f
C490 B.n450 VSUBS 0.008039f
C491 B.n451 VSUBS 0.008039f
C492 B.n452 VSUBS 0.008039f
C493 B.n453 VSUBS 0.008039f
C494 B.n454 VSUBS 0.008039f
C495 B.n455 VSUBS 0.008039f
C496 B.n456 VSUBS 0.008039f
C497 B.n457 VSUBS 0.008039f
C498 B.n458 VSUBS 0.008039f
C499 B.n459 VSUBS 0.008039f
C500 B.n460 VSUBS 0.008039f
C501 B.n461 VSUBS 0.008039f
C502 B.n462 VSUBS 0.008039f
C503 B.n463 VSUBS 0.008039f
C504 B.n464 VSUBS 0.008039f
C505 B.n465 VSUBS 0.008039f
C506 B.n466 VSUBS 0.008039f
C507 B.n467 VSUBS 0.008039f
C508 B.n468 VSUBS 0.008039f
C509 B.n469 VSUBS 0.008039f
C510 B.n470 VSUBS 0.008039f
C511 B.n471 VSUBS 0.008039f
C512 B.n472 VSUBS 0.008039f
C513 B.n473 VSUBS 0.008039f
C514 B.n474 VSUBS 0.008039f
C515 B.n475 VSUBS 0.008039f
C516 B.n476 VSUBS 0.008039f
C517 B.n477 VSUBS 0.008039f
C518 B.n478 VSUBS 0.008039f
C519 B.n479 VSUBS 0.008039f
C520 B.n480 VSUBS 0.008039f
C521 B.n481 VSUBS 0.008039f
C522 B.n482 VSUBS 0.008039f
C523 B.n483 VSUBS 0.008039f
C524 B.n484 VSUBS 0.008039f
C525 B.n485 VSUBS 0.008039f
C526 B.n486 VSUBS 0.008039f
C527 B.n487 VSUBS 0.008039f
C528 B.n488 VSUBS 0.008039f
C529 B.n489 VSUBS 0.008039f
C530 B.n490 VSUBS 0.008039f
C531 B.n491 VSUBS 0.008039f
C532 B.n492 VSUBS 0.008039f
C533 B.n493 VSUBS 0.008039f
C534 B.n494 VSUBS 0.008039f
C535 B.n495 VSUBS 0.008039f
C536 B.n496 VSUBS 0.008039f
C537 B.n497 VSUBS 0.008039f
C538 B.n498 VSUBS 0.008039f
C539 B.n499 VSUBS 0.008039f
C540 B.n500 VSUBS 0.008039f
C541 B.n501 VSUBS 0.008039f
C542 B.n502 VSUBS 0.008039f
C543 B.n503 VSUBS 0.008039f
C544 B.n504 VSUBS 0.008039f
C545 B.n505 VSUBS 0.008039f
C546 B.n506 VSUBS 0.008039f
C547 B.n507 VSUBS 0.008039f
C548 B.n508 VSUBS 0.008039f
C549 B.n509 VSUBS 0.008039f
C550 B.n510 VSUBS 0.008039f
C551 B.n511 VSUBS 0.008039f
C552 B.n512 VSUBS 0.008039f
C553 B.n513 VSUBS 0.008039f
C554 B.n514 VSUBS 0.008039f
C555 B.n515 VSUBS 0.008039f
C556 B.n516 VSUBS 0.008039f
C557 B.n517 VSUBS 0.008039f
C558 B.n518 VSUBS 0.008039f
C559 B.n519 VSUBS 0.008039f
C560 B.n520 VSUBS 0.008039f
C561 B.n521 VSUBS 0.008039f
C562 B.n522 VSUBS 0.008039f
C563 B.n523 VSUBS 0.008039f
C564 B.n524 VSUBS 0.008039f
C565 B.n525 VSUBS 0.008039f
C566 B.n526 VSUBS 0.008039f
C567 B.n527 VSUBS 0.008039f
C568 B.n528 VSUBS 0.008039f
C569 B.n529 VSUBS 0.008039f
C570 B.n530 VSUBS 0.008039f
C571 B.n531 VSUBS 0.008039f
C572 B.n532 VSUBS 0.008039f
C573 B.n533 VSUBS 0.008039f
C574 B.n534 VSUBS 0.008039f
C575 B.n535 VSUBS 0.008039f
C576 B.n536 VSUBS 0.008039f
C577 B.n537 VSUBS 0.008039f
C578 B.n538 VSUBS 0.008039f
C579 B.n539 VSUBS 0.008039f
C580 B.n540 VSUBS 0.008039f
C581 B.n541 VSUBS 0.008039f
C582 B.n542 VSUBS 0.008039f
C583 B.n543 VSUBS 0.008039f
C584 B.n544 VSUBS 0.008039f
C585 B.n545 VSUBS 0.008039f
C586 B.n546 VSUBS 0.008039f
C587 B.n547 VSUBS 0.008039f
C588 B.n548 VSUBS 0.008039f
C589 B.n549 VSUBS 0.008039f
C590 B.n550 VSUBS 0.008039f
C591 B.n551 VSUBS 0.008039f
C592 B.n552 VSUBS 0.008039f
C593 B.n553 VSUBS 0.008039f
C594 B.n554 VSUBS 0.008039f
C595 B.n555 VSUBS 0.008039f
C596 B.n556 VSUBS 0.008039f
C597 B.n557 VSUBS 0.008039f
C598 B.n558 VSUBS 0.008039f
C599 B.n559 VSUBS 0.008039f
C600 B.n560 VSUBS 0.008039f
C601 B.n561 VSUBS 0.008039f
C602 B.n562 VSUBS 0.008039f
C603 B.n563 VSUBS 0.008039f
C604 B.n564 VSUBS 0.008039f
C605 B.n565 VSUBS 0.008039f
C606 B.n566 VSUBS 0.008039f
C607 B.n567 VSUBS 0.008039f
C608 B.n568 VSUBS 0.008039f
C609 B.n569 VSUBS 0.008039f
C610 B.n570 VSUBS 0.019289f
C611 B.n571 VSUBS 0.02018f
C612 B.n572 VSUBS 0.019071f
C613 B.n573 VSUBS 0.008039f
C614 B.n574 VSUBS 0.008039f
C615 B.n575 VSUBS 0.008039f
C616 B.n576 VSUBS 0.008039f
C617 B.n577 VSUBS 0.008039f
C618 B.n578 VSUBS 0.008039f
C619 B.n579 VSUBS 0.008039f
C620 B.n580 VSUBS 0.008039f
C621 B.n581 VSUBS 0.008039f
C622 B.n582 VSUBS 0.008039f
C623 B.n583 VSUBS 0.008039f
C624 B.n584 VSUBS 0.008039f
C625 B.n585 VSUBS 0.008039f
C626 B.n586 VSUBS 0.008039f
C627 B.n587 VSUBS 0.008039f
C628 B.n588 VSUBS 0.008039f
C629 B.n589 VSUBS 0.008039f
C630 B.n590 VSUBS 0.008039f
C631 B.n591 VSUBS 0.008039f
C632 B.n592 VSUBS 0.008039f
C633 B.n593 VSUBS 0.008039f
C634 B.n594 VSUBS 0.008039f
C635 B.n595 VSUBS 0.008039f
C636 B.n596 VSUBS 0.008039f
C637 B.n597 VSUBS 0.008039f
C638 B.n598 VSUBS 0.008039f
C639 B.n599 VSUBS 0.008039f
C640 B.n600 VSUBS 0.008039f
C641 B.n601 VSUBS 0.008039f
C642 B.n602 VSUBS 0.008039f
C643 B.n603 VSUBS 0.008039f
C644 B.n604 VSUBS 0.008039f
C645 B.n605 VSUBS 0.008039f
C646 B.n606 VSUBS 0.008039f
C647 B.n607 VSUBS 0.008039f
C648 B.n608 VSUBS 0.008039f
C649 B.n609 VSUBS 0.008039f
C650 B.n610 VSUBS 0.008039f
C651 B.n611 VSUBS 0.008039f
C652 B.n612 VSUBS 0.008039f
C653 B.n613 VSUBS 0.008039f
C654 B.n614 VSUBS 0.008039f
C655 B.n615 VSUBS 0.008039f
C656 B.n616 VSUBS 0.008039f
C657 B.n617 VSUBS 0.008039f
C658 B.n618 VSUBS 0.008039f
C659 B.n619 VSUBS 0.008039f
C660 B.n620 VSUBS 0.008039f
C661 B.n621 VSUBS 0.007567f
C662 B.n622 VSUBS 0.008039f
C663 B.n623 VSUBS 0.008039f
C664 B.n624 VSUBS 0.004493f
C665 B.n625 VSUBS 0.008039f
C666 B.n626 VSUBS 0.008039f
C667 B.n627 VSUBS 0.008039f
C668 B.n628 VSUBS 0.008039f
C669 B.n629 VSUBS 0.008039f
C670 B.n630 VSUBS 0.008039f
C671 B.n631 VSUBS 0.008039f
C672 B.n632 VSUBS 0.008039f
C673 B.n633 VSUBS 0.008039f
C674 B.n634 VSUBS 0.008039f
C675 B.n635 VSUBS 0.008039f
C676 B.n636 VSUBS 0.008039f
C677 B.n637 VSUBS 0.004493f
C678 B.n638 VSUBS 0.018626f
C679 B.n639 VSUBS 0.007567f
C680 B.n640 VSUBS 0.008039f
C681 B.n641 VSUBS 0.008039f
C682 B.n642 VSUBS 0.008039f
C683 B.n643 VSUBS 0.008039f
C684 B.n644 VSUBS 0.008039f
C685 B.n645 VSUBS 0.008039f
C686 B.n646 VSUBS 0.008039f
C687 B.n647 VSUBS 0.008039f
C688 B.n648 VSUBS 0.008039f
C689 B.n649 VSUBS 0.008039f
C690 B.n650 VSUBS 0.008039f
C691 B.n651 VSUBS 0.008039f
C692 B.n652 VSUBS 0.008039f
C693 B.n653 VSUBS 0.008039f
C694 B.n654 VSUBS 0.008039f
C695 B.n655 VSUBS 0.008039f
C696 B.n656 VSUBS 0.008039f
C697 B.n657 VSUBS 0.008039f
C698 B.n658 VSUBS 0.008039f
C699 B.n659 VSUBS 0.008039f
C700 B.n660 VSUBS 0.008039f
C701 B.n661 VSUBS 0.008039f
C702 B.n662 VSUBS 0.008039f
C703 B.n663 VSUBS 0.008039f
C704 B.n664 VSUBS 0.008039f
C705 B.n665 VSUBS 0.008039f
C706 B.n666 VSUBS 0.008039f
C707 B.n667 VSUBS 0.008039f
C708 B.n668 VSUBS 0.008039f
C709 B.n669 VSUBS 0.008039f
C710 B.n670 VSUBS 0.008039f
C711 B.n671 VSUBS 0.008039f
C712 B.n672 VSUBS 0.008039f
C713 B.n673 VSUBS 0.008039f
C714 B.n674 VSUBS 0.008039f
C715 B.n675 VSUBS 0.008039f
C716 B.n676 VSUBS 0.008039f
C717 B.n677 VSUBS 0.008039f
C718 B.n678 VSUBS 0.008039f
C719 B.n679 VSUBS 0.008039f
C720 B.n680 VSUBS 0.008039f
C721 B.n681 VSUBS 0.008039f
C722 B.n682 VSUBS 0.008039f
C723 B.n683 VSUBS 0.008039f
C724 B.n684 VSUBS 0.008039f
C725 B.n685 VSUBS 0.008039f
C726 B.n686 VSUBS 0.008039f
C727 B.n687 VSUBS 0.008039f
C728 B.n688 VSUBS 0.008039f
C729 B.n689 VSUBS 0.019963f
C730 B.n690 VSUBS 0.019289f
C731 B.n691 VSUBS 0.019289f
C732 B.n692 VSUBS 0.008039f
C733 B.n693 VSUBS 0.008039f
C734 B.n694 VSUBS 0.008039f
C735 B.n695 VSUBS 0.008039f
C736 B.n696 VSUBS 0.008039f
C737 B.n697 VSUBS 0.008039f
C738 B.n698 VSUBS 0.008039f
C739 B.n699 VSUBS 0.008039f
C740 B.n700 VSUBS 0.008039f
C741 B.n701 VSUBS 0.008039f
C742 B.n702 VSUBS 0.008039f
C743 B.n703 VSUBS 0.008039f
C744 B.n704 VSUBS 0.008039f
C745 B.n705 VSUBS 0.008039f
C746 B.n706 VSUBS 0.008039f
C747 B.n707 VSUBS 0.008039f
C748 B.n708 VSUBS 0.008039f
C749 B.n709 VSUBS 0.008039f
C750 B.n710 VSUBS 0.008039f
C751 B.n711 VSUBS 0.008039f
C752 B.n712 VSUBS 0.008039f
C753 B.n713 VSUBS 0.008039f
C754 B.n714 VSUBS 0.008039f
C755 B.n715 VSUBS 0.008039f
C756 B.n716 VSUBS 0.008039f
C757 B.n717 VSUBS 0.008039f
C758 B.n718 VSUBS 0.008039f
C759 B.n719 VSUBS 0.008039f
C760 B.n720 VSUBS 0.008039f
C761 B.n721 VSUBS 0.008039f
C762 B.n722 VSUBS 0.008039f
C763 B.n723 VSUBS 0.008039f
C764 B.n724 VSUBS 0.008039f
C765 B.n725 VSUBS 0.008039f
C766 B.n726 VSUBS 0.008039f
C767 B.n727 VSUBS 0.008039f
C768 B.n728 VSUBS 0.008039f
C769 B.n729 VSUBS 0.008039f
C770 B.n730 VSUBS 0.008039f
C771 B.n731 VSUBS 0.008039f
C772 B.n732 VSUBS 0.008039f
C773 B.n733 VSUBS 0.008039f
C774 B.n734 VSUBS 0.008039f
C775 B.n735 VSUBS 0.008039f
C776 B.n736 VSUBS 0.008039f
C777 B.n737 VSUBS 0.008039f
C778 B.n738 VSUBS 0.008039f
C779 B.n739 VSUBS 0.008039f
C780 B.n740 VSUBS 0.008039f
C781 B.n741 VSUBS 0.008039f
C782 B.n742 VSUBS 0.008039f
C783 B.n743 VSUBS 0.008039f
C784 B.n744 VSUBS 0.008039f
C785 B.n745 VSUBS 0.008039f
C786 B.n746 VSUBS 0.008039f
C787 B.n747 VSUBS 0.008039f
C788 B.n748 VSUBS 0.008039f
C789 B.n749 VSUBS 0.008039f
C790 B.n750 VSUBS 0.008039f
C791 B.n751 VSUBS 0.008039f
C792 B.n752 VSUBS 0.008039f
C793 B.n753 VSUBS 0.008039f
C794 B.n754 VSUBS 0.008039f
C795 B.n755 VSUBS 0.008039f
C796 B.n756 VSUBS 0.008039f
C797 B.n757 VSUBS 0.008039f
C798 B.n758 VSUBS 0.008039f
C799 B.n759 VSUBS 0.008039f
C800 B.n760 VSUBS 0.008039f
C801 B.n761 VSUBS 0.008039f
C802 B.n762 VSUBS 0.008039f
C803 B.n763 VSUBS 0.008039f
C804 B.n764 VSUBS 0.008039f
C805 B.n765 VSUBS 0.008039f
C806 B.n766 VSUBS 0.008039f
C807 B.n767 VSUBS 0.008039f
C808 B.n768 VSUBS 0.008039f
C809 B.n769 VSUBS 0.008039f
C810 B.n770 VSUBS 0.008039f
C811 B.n771 VSUBS 0.008039f
C812 B.n772 VSUBS 0.008039f
C813 B.n773 VSUBS 0.008039f
C814 B.n774 VSUBS 0.008039f
C815 B.n775 VSUBS 0.018204f
C816 VDD1.t7 VSUBS 0.186026f
C817 VDD1.t6 VSUBS 0.186026f
C818 VDD1.n0 VSUBS 1.40317f
C819 VDD1.t1 VSUBS 0.186026f
C820 VDD1.t5 VSUBS 0.186026f
C821 VDD1.n1 VSUBS 1.40189f
C822 VDD1.t3 VSUBS 0.186026f
C823 VDD1.t0 VSUBS 0.186026f
C824 VDD1.n2 VSUBS 1.40189f
C825 VDD1.n3 VSUBS 3.8025f
C826 VDD1.t4 VSUBS 0.186026f
C827 VDD1.t2 VSUBS 0.186026f
C828 VDD1.n4 VSUBS 1.38829f
C829 VDD1.n5 VSUBS 3.11118f
C830 VP.t7 VSUBS 2.44966f
C831 VP.n0 VSUBS 0.998389f
C832 VP.n1 VSUBS 0.032404f
C833 VP.n2 VSUBS 0.048f
C834 VP.n3 VSUBS 0.032404f
C835 VP.t4 VSUBS 2.44966f
C836 VP.n4 VSUBS 0.06009f
C837 VP.n5 VSUBS 0.032404f
C838 VP.n6 VSUBS 0.06009f
C839 VP.n7 VSUBS 0.032404f
C840 VP.t2 VSUBS 2.44966f
C841 VP.n8 VSUBS 0.048f
C842 VP.n9 VSUBS 0.032404f
C843 VP.t6 VSUBS 2.44966f
C844 VP.n10 VSUBS 0.998389f
C845 VP.t5 VSUBS 2.44966f
C846 VP.n11 VSUBS 0.998389f
C847 VP.n12 VSUBS 0.032404f
C848 VP.n13 VSUBS 0.048f
C849 VP.n14 VSUBS 0.032404f
C850 VP.t3 VSUBS 2.44966f
C851 VP.n15 VSUBS 0.06009f
C852 VP.n16 VSUBS 0.032404f
C853 VP.n17 VSUBS 0.06009f
C854 VP.t0 VSUBS 2.76254f
C855 VP.n18 VSUBS 0.938843f
C856 VP.t1 VSUBS 2.44966f
C857 VP.n19 VSUBS 0.969869f
C858 VP.n20 VSUBS 0.038138f
C859 VP.n21 VSUBS 0.348123f
C860 VP.n22 VSUBS 0.032404f
C861 VP.n23 VSUBS 0.032404f
C862 VP.n24 VSUBS 0.064063f
C863 VP.n25 VSUBS 0.026171f
C864 VP.n26 VSUBS 0.064063f
C865 VP.n27 VSUBS 0.032404f
C866 VP.n28 VSUBS 0.032404f
C867 VP.n29 VSUBS 0.032404f
C868 VP.n30 VSUBS 0.038138f
C869 VP.n31 VSUBS 0.875782f
C870 VP.n32 VSUBS 0.052377f
C871 VP.n33 VSUBS 0.06009f
C872 VP.n34 VSUBS 0.032404f
C873 VP.n35 VSUBS 0.032404f
C874 VP.n36 VSUBS 0.032404f
C875 VP.n37 VSUBS 0.046207f
C876 VP.n38 VSUBS 0.06009f
C877 VP.n39 VSUBS 0.053563f
C878 VP.n40 VSUBS 0.052291f
C879 VP.n41 VSUBS 1.86612f
C880 VP.n42 VSUBS 1.88918f
C881 VP.n43 VSUBS 0.052291f
C882 VP.n44 VSUBS 0.053563f
C883 VP.n45 VSUBS 0.06009f
C884 VP.n46 VSUBS 0.046207f
C885 VP.n47 VSUBS 0.032404f
C886 VP.n48 VSUBS 0.032404f
C887 VP.n49 VSUBS 0.032404f
C888 VP.n50 VSUBS 0.06009f
C889 VP.n51 VSUBS 0.052377f
C890 VP.n52 VSUBS 0.875782f
C891 VP.n53 VSUBS 0.038138f
C892 VP.n54 VSUBS 0.032404f
C893 VP.n55 VSUBS 0.032404f
C894 VP.n56 VSUBS 0.032404f
C895 VP.n57 VSUBS 0.064063f
C896 VP.n58 VSUBS 0.026171f
C897 VP.n59 VSUBS 0.064063f
C898 VP.n60 VSUBS 0.032404f
C899 VP.n61 VSUBS 0.032404f
C900 VP.n62 VSUBS 0.032404f
C901 VP.n63 VSUBS 0.038138f
C902 VP.n64 VSUBS 0.875782f
C903 VP.n65 VSUBS 0.052377f
C904 VP.n66 VSUBS 0.06009f
C905 VP.n67 VSUBS 0.032404f
C906 VP.n68 VSUBS 0.032404f
C907 VP.n69 VSUBS 0.032404f
C908 VP.n70 VSUBS 0.046207f
C909 VP.n71 VSUBS 0.06009f
C910 VP.n72 VSUBS 0.053563f
C911 VP.n73 VSUBS 0.052291f
C912 VP.n74 VSUBS 0.067928f
C913 VDD2.t2 VSUBS 0.208375f
C914 VDD2.t7 VSUBS 0.208375f
C915 VDD2.n0 VSUBS 1.57031f
C916 VDD2.t1 VSUBS 0.208375f
C917 VDD2.t6 VSUBS 0.208375f
C918 VDD2.n1 VSUBS 1.57031f
C919 VDD2.n2 VSUBS 4.20187f
C920 VDD2.t4 VSUBS 0.208375f
C921 VDD2.t5 VSUBS 0.208375f
C922 VDD2.n3 VSUBS 1.55508f
C923 VDD2.n4 VSUBS 3.45068f
C924 VDD2.t0 VSUBS 0.208375f
C925 VDD2.t3 VSUBS 0.208375f
C926 VDD2.n5 VSUBS 1.57026f
C927 VTAIL.t10 VSUBS 0.200019f
C928 VTAIL.t9 VSUBS 0.200019f
C929 VTAIL.n0 VSUBS 1.36119f
C930 VTAIL.n1 VSUBS 0.818703f
C931 VTAIL.t8 VSUBS 1.81495f
C932 VTAIL.n2 VSUBS 0.945641f
C933 VTAIL.t4 VSUBS 1.81495f
C934 VTAIL.n3 VSUBS 0.945641f
C935 VTAIL.t5 VSUBS 0.200019f
C936 VTAIL.t0 VSUBS 0.200019f
C937 VTAIL.n4 VSUBS 1.36119f
C938 VTAIL.n5 VSUBS 1.05399f
C939 VTAIL.t6 VSUBS 1.81495f
C940 VTAIL.n6 VSUBS 2.20924f
C941 VTAIL.t15 VSUBS 1.81496f
C942 VTAIL.n7 VSUBS 2.20922f
C943 VTAIL.t11 VSUBS 0.200019f
C944 VTAIL.t12 VSUBS 0.200019f
C945 VTAIL.n8 VSUBS 1.3612f
C946 VTAIL.n9 VSUBS 1.05398f
C947 VTAIL.t13 VSUBS 1.81496f
C948 VTAIL.n10 VSUBS 0.945628f
C949 VTAIL.t1 VSUBS 1.81496f
C950 VTAIL.n11 VSUBS 0.945628f
C951 VTAIL.t3 VSUBS 0.200019f
C952 VTAIL.t7 VSUBS 0.200019f
C953 VTAIL.n12 VSUBS 1.3612f
C954 VTAIL.n13 VSUBS 1.05398f
C955 VTAIL.t2 VSUBS 1.81495f
C956 VTAIL.n14 VSUBS 2.20924f
C957 VTAIL.t14 VSUBS 1.81495f
C958 VTAIL.n15 VSUBS 2.20426f
C959 VN.t1 VSUBS 2.22596f
C960 VN.n0 VSUBS 0.907217f
C961 VN.n1 VSUBS 0.029445f
C962 VN.n2 VSUBS 0.043617f
C963 VN.n3 VSUBS 0.029445f
C964 VN.t6 VSUBS 2.22596f
C965 VN.n4 VSUBS 0.054602f
C966 VN.n5 VSUBS 0.029445f
C967 VN.n6 VSUBS 0.054602f
C968 VN.t5 VSUBS 2.51027f
C969 VN.n7 VSUBS 0.853107f
C970 VN.t0 VSUBS 2.22596f
C971 VN.n8 VSUBS 0.881301f
C972 VN.n9 VSUBS 0.034655f
C973 VN.n10 VSUBS 0.316332f
C974 VN.n11 VSUBS 0.029445f
C975 VN.n12 VSUBS 0.029445f
C976 VN.n13 VSUBS 0.058213f
C977 VN.n14 VSUBS 0.023781f
C978 VN.n15 VSUBS 0.058213f
C979 VN.n16 VSUBS 0.029445f
C980 VN.n17 VSUBS 0.029445f
C981 VN.n18 VSUBS 0.029445f
C982 VN.n19 VSUBS 0.034655f
C983 VN.n20 VSUBS 0.795807f
C984 VN.n21 VSUBS 0.047594f
C985 VN.n22 VSUBS 0.054602f
C986 VN.n23 VSUBS 0.029445f
C987 VN.n24 VSUBS 0.029445f
C988 VN.n25 VSUBS 0.029445f
C989 VN.n26 VSUBS 0.041988f
C990 VN.n27 VSUBS 0.054602f
C991 VN.n28 VSUBS 0.048672f
C992 VN.n29 VSUBS 0.047516f
C993 VN.n30 VSUBS 0.061725f
C994 VN.t3 VSUBS 2.22596f
C995 VN.n31 VSUBS 0.907217f
C996 VN.n32 VSUBS 0.029445f
C997 VN.n33 VSUBS 0.043617f
C998 VN.n34 VSUBS 0.029445f
C999 VN.t2 VSUBS 2.22596f
C1000 VN.n35 VSUBS 0.054602f
C1001 VN.n36 VSUBS 0.029445f
C1002 VN.n37 VSUBS 0.054602f
C1003 VN.t4 VSUBS 2.51027f
C1004 VN.n38 VSUBS 0.853107f
C1005 VN.t7 VSUBS 2.22596f
C1006 VN.n39 VSUBS 0.881301f
C1007 VN.n40 VSUBS 0.034655f
C1008 VN.n41 VSUBS 0.316332f
C1009 VN.n42 VSUBS 0.029445f
C1010 VN.n43 VSUBS 0.029445f
C1011 VN.n44 VSUBS 0.058213f
C1012 VN.n45 VSUBS 0.023781f
C1013 VN.n46 VSUBS 0.058213f
C1014 VN.n47 VSUBS 0.029445f
C1015 VN.n48 VSUBS 0.029445f
C1016 VN.n49 VSUBS 0.029445f
C1017 VN.n50 VSUBS 0.034655f
C1018 VN.n51 VSUBS 0.795807f
C1019 VN.n52 VSUBS 0.047594f
C1020 VN.n53 VSUBS 0.054602f
C1021 VN.n54 VSUBS 0.029445f
C1022 VN.n55 VSUBS 0.029445f
C1023 VN.n56 VSUBS 0.029445f
C1024 VN.n57 VSUBS 0.041988f
C1025 VN.n58 VSUBS 0.054602f
C1026 VN.n59 VSUBS 0.048672f
C1027 VN.n60 VSUBS 0.047516f
C1028 VN.n61 VSUBS 1.70771f
.ends

