* NGSPICE file created from diff_pair_sample_1794.ext - technology: sky130A

.subckt diff_pair_sample_1794 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t19 VP.t0 VDD1.t9 B.t1 sky130_fd_pr__nfet_01v8 ad=2.8941 pd=17.87 as=2.8941 ps=17.87 w=17.54 l=2.83
X1 VTAIL.t2 VN.t0 VDD2.t9 B.t2 sky130_fd_pr__nfet_01v8 ad=2.8941 pd=17.87 as=2.8941 ps=17.87 w=17.54 l=2.83
X2 B.t23 B.t21 B.t22 B.t11 sky130_fd_pr__nfet_01v8 ad=6.8406 pd=35.86 as=0 ps=0 w=17.54 l=2.83
X3 VDD2.t8 VN.t1 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=2.8941 pd=17.87 as=2.8941 ps=17.87 w=17.54 l=2.83
X4 VDD2.t7 VN.t2 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=6.8406 pd=35.86 as=2.8941 ps=17.87 w=17.54 l=2.83
X5 VDD1.t8 VP.t1 VTAIL.t18 B.t6 sky130_fd_pr__nfet_01v8 ad=2.8941 pd=17.87 as=2.8941 ps=17.87 w=17.54 l=2.83
X6 VDD1.t5 VP.t2 VTAIL.t17 B.t5 sky130_fd_pr__nfet_01v8 ad=2.8941 pd=17.87 as=6.8406 ps=35.86 w=17.54 l=2.83
X7 VTAIL.t3 VN.t3 VDD2.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=2.8941 pd=17.87 as=2.8941 ps=17.87 w=17.54 l=2.83
X8 VTAIL.t4 VN.t4 VDD2.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=2.8941 pd=17.87 as=2.8941 ps=17.87 w=17.54 l=2.83
X9 VTAIL.t16 VP.t3 VDD1.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=2.8941 pd=17.87 as=2.8941 ps=17.87 w=17.54 l=2.83
X10 B.t20 B.t18 B.t19 B.t15 sky130_fd_pr__nfet_01v8 ad=6.8406 pd=35.86 as=0 ps=0 w=17.54 l=2.83
X11 VTAIL.t15 VP.t4 VDD1.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=2.8941 pd=17.87 as=2.8941 ps=17.87 w=17.54 l=2.83
X12 VTAIL.t1 VN.t5 VDD2.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=2.8941 pd=17.87 as=2.8941 ps=17.87 w=17.54 l=2.83
X13 VDD2.t3 VN.t6 VTAIL.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=2.8941 pd=17.87 as=2.8941 ps=17.87 w=17.54 l=2.83
X14 VDD2.t2 VN.t7 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=2.8941 pd=17.87 as=6.8406 ps=35.86 w=17.54 l=2.83
X15 VDD1.t6 VP.t5 VTAIL.t14 B.t9 sky130_fd_pr__nfet_01v8 ad=6.8406 pd=35.86 as=2.8941 ps=17.87 w=17.54 l=2.83
X16 VDD1.t1 VP.t6 VTAIL.t13 B.t7 sky130_fd_pr__nfet_01v8 ad=2.8941 pd=17.87 as=6.8406 ps=35.86 w=17.54 l=2.83
X17 VDD2.t1 VN.t8 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.8941 pd=17.87 as=6.8406 ps=35.86 w=17.54 l=2.83
X18 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=6.8406 pd=35.86 as=0 ps=0 w=17.54 l=2.83
X19 VDD1.t0 VP.t7 VTAIL.t12 B.t8 sky130_fd_pr__nfet_01v8 ad=2.8941 pd=17.87 as=2.8941 ps=17.87 w=17.54 l=2.83
X20 VTAIL.t11 VP.t8 VDD1.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=2.8941 pd=17.87 as=2.8941 ps=17.87 w=17.54 l=2.83
X21 VDD1.t2 VP.t9 VTAIL.t10 B.t0 sky130_fd_pr__nfet_01v8 ad=6.8406 pd=35.86 as=2.8941 ps=17.87 w=17.54 l=2.83
X22 VDD2.t0 VN.t9 VTAIL.t9 B.t9 sky130_fd_pr__nfet_01v8 ad=6.8406 pd=35.86 as=2.8941 ps=17.87 w=17.54 l=2.83
X23 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=6.8406 pd=35.86 as=0 ps=0 w=17.54 l=2.83
R0 VP.n25 VP.t9 182.843
R1 VP.n26 VP.n23 161.3
R2 VP.n28 VP.n27 161.3
R3 VP.n29 VP.n22 161.3
R4 VP.n31 VP.n30 161.3
R5 VP.n32 VP.n21 161.3
R6 VP.n34 VP.n33 161.3
R7 VP.n36 VP.n20 161.3
R8 VP.n38 VP.n37 161.3
R9 VP.n39 VP.n19 161.3
R10 VP.n41 VP.n40 161.3
R11 VP.n42 VP.n18 161.3
R12 VP.n45 VP.n44 161.3
R13 VP.n46 VP.n17 161.3
R14 VP.n48 VP.n47 161.3
R15 VP.n49 VP.n16 161.3
R16 VP.n51 VP.n50 161.3
R17 VP.n52 VP.n15 161.3
R18 VP.n54 VP.n53 161.3
R19 VP.n55 VP.n14 161.3
R20 VP.n100 VP.n0 161.3
R21 VP.n99 VP.n98 161.3
R22 VP.n97 VP.n1 161.3
R23 VP.n96 VP.n95 161.3
R24 VP.n94 VP.n2 161.3
R25 VP.n93 VP.n92 161.3
R26 VP.n91 VP.n3 161.3
R27 VP.n90 VP.n89 161.3
R28 VP.n87 VP.n4 161.3
R29 VP.n86 VP.n85 161.3
R30 VP.n84 VP.n5 161.3
R31 VP.n83 VP.n82 161.3
R32 VP.n81 VP.n6 161.3
R33 VP.n79 VP.n78 161.3
R34 VP.n77 VP.n7 161.3
R35 VP.n76 VP.n75 161.3
R36 VP.n74 VP.n8 161.3
R37 VP.n73 VP.n72 161.3
R38 VP.n71 VP.n9 161.3
R39 VP.n70 VP.n69 161.3
R40 VP.n67 VP.n10 161.3
R41 VP.n66 VP.n65 161.3
R42 VP.n64 VP.n11 161.3
R43 VP.n63 VP.n62 161.3
R44 VP.n61 VP.n12 161.3
R45 VP.n60 VP.n59 161.3
R46 VP.n13 VP.t5 149.369
R47 VP.n68 VP.t8 149.369
R48 VP.n80 VP.t7 149.369
R49 VP.n88 VP.t3 149.369
R50 VP.n101 VP.t2 149.369
R51 VP.n56 VP.t6 149.369
R52 VP.n43 VP.t0 149.369
R53 VP.n35 VP.t1 149.369
R54 VP.n24 VP.t4 149.369
R55 VP.n58 VP.n13 107.466
R56 VP.n102 VP.n101 107.466
R57 VP.n57 VP.n56 107.466
R58 VP.n58 VP.n57 58.5375
R59 VP.n75 VP.n74 56.5617
R60 VP.n86 VP.n5 56.5617
R61 VP.n41 VP.n19 56.5617
R62 VP.n30 VP.n29 56.5617
R63 VP.n25 VP.n24 53.6463
R64 VP.n66 VP.n11 41.5458
R65 VP.n95 VP.n94 41.5458
R66 VP.n50 VP.n49 41.5458
R67 VP.n62 VP.n11 39.6083
R68 VP.n95 VP.n1 39.6083
R69 VP.n50 VP.n15 39.6083
R70 VP.n61 VP.n60 24.5923
R71 VP.n62 VP.n61 24.5923
R72 VP.n67 VP.n66 24.5923
R73 VP.n69 VP.n67 24.5923
R74 VP.n73 VP.n9 24.5923
R75 VP.n74 VP.n73 24.5923
R76 VP.n75 VP.n7 24.5923
R77 VP.n79 VP.n7 24.5923
R78 VP.n82 VP.n81 24.5923
R79 VP.n82 VP.n5 24.5923
R80 VP.n87 VP.n86 24.5923
R81 VP.n89 VP.n87 24.5923
R82 VP.n93 VP.n3 24.5923
R83 VP.n94 VP.n93 24.5923
R84 VP.n99 VP.n1 24.5923
R85 VP.n100 VP.n99 24.5923
R86 VP.n54 VP.n15 24.5923
R87 VP.n55 VP.n54 24.5923
R88 VP.n42 VP.n41 24.5923
R89 VP.n44 VP.n42 24.5923
R90 VP.n48 VP.n17 24.5923
R91 VP.n49 VP.n48 24.5923
R92 VP.n30 VP.n21 24.5923
R93 VP.n34 VP.n21 24.5923
R94 VP.n37 VP.n36 24.5923
R95 VP.n37 VP.n19 24.5923
R96 VP.n28 VP.n23 24.5923
R97 VP.n29 VP.n28 24.5923
R98 VP.n68 VP.n9 20.1658
R99 VP.n89 VP.n88 20.1658
R100 VP.n44 VP.n43 20.1658
R101 VP.n24 VP.n23 20.1658
R102 VP.n80 VP.n79 12.2964
R103 VP.n81 VP.n80 12.2964
R104 VP.n35 VP.n34 12.2964
R105 VP.n36 VP.n35 12.2964
R106 VP.n26 VP.n25 5.0289
R107 VP.n69 VP.n68 4.42703
R108 VP.n88 VP.n3 4.42703
R109 VP.n43 VP.n17 4.42703
R110 VP.n60 VP.n13 3.44336
R111 VP.n101 VP.n100 3.44336
R112 VP.n56 VP.n55 3.44336
R113 VP.n57 VP.n14 0.278335
R114 VP.n59 VP.n58 0.278335
R115 VP.n102 VP.n0 0.278335
R116 VP.n27 VP.n26 0.189894
R117 VP.n27 VP.n22 0.189894
R118 VP.n31 VP.n22 0.189894
R119 VP.n32 VP.n31 0.189894
R120 VP.n33 VP.n32 0.189894
R121 VP.n33 VP.n20 0.189894
R122 VP.n38 VP.n20 0.189894
R123 VP.n39 VP.n38 0.189894
R124 VP.n40 VP.n39 0.189894
R125 VP.n40 VP.n18 0.189894
R126 VP.n45 VP.n18 0.189894
R127 VP.n46 VP.n45 0.189894
R128 VP.n47 VP.n46 0.189894
R129 VP.n47 VP.n16 0.189894
R130 VP.n51 VP.n16 0.189894
R131 VP.n52 VP.n51 0.189894
R132 VP.n53 VP.n52 0.189894
R133 VP.n53 VP.n14 0.189894
R134 VP.n59 VP.n12 0.189894
R135 VP.n63 VP.n12 0.189894
R136 VP.n64 VP.n63 0.189894
R137 VP.n65 VP.n64 0.189894
R138 VP.n65 VP.n10 0.189894
R139 VP.n70 VP.n10 0.189894
R140 VP.n71 VP.n70 0.189894
R141 VP.n72 VP.n71 0.189894
R142 VP.n72 VP.n8 0.189894
R143 VP.n76 VP.n8 0.189894
R144 VP.n77 VP.n76 0.189894
R145 VP.n78 VP.n77 0.189894
R146 VP.n78 VP.n6 0.189894
R147 VP.n83 VP.n6 0.189894
R148 VP.n84 VP.n83 0.189894
R149 VP.n85 VP.n84 0.189894
R150 VP.n85 VP.n4 0.189894
R151 VP.n90 VP.n4 0.189894
R152 VP.n91 VP.n90 0.189894
R153 VP.n92 VP.n91 0.189894
R154 VP.n92 VP.n2 0.189894
R155 VP.n96 VP.n2 0.189894
R156 VP.n97 VP.n96 0.189894
R157 VP.n98 VP.n97 0.189894
R158 VP.n98 VP.n0 0.189894
R159 VP VP.n102 0.153485
R160 VDD1.n92 VDD1.n0 289.615
R161 VDD1.n191 VDD1.n99 289.615
R162 VDD1.n93 VDD1.n92 185
R163 VDD1.n91 VDD1.n90 185
R164 VDD1.n4 VDD1.n3 185
R165 VDD1.n85 VDD1.n84 185
R166 VDD1.n83 VDD1.n82 185
R167 VDD1.n8 VDD1.n7 185
R168 VDD1.n12 VDD1.n10 185
R169 VDD1.n77 VDD1.n76 185
R170 VDD1.n75 VDD1.n74 185
R171 VDD1.n14 VDD1.n13 185
R172 VDD1.n69 VDD1.n68 185
R173 VDD1.n67 VDD1.n66 185
R174 VDD1.n18 VDD1.n17 185
R175 VDD1.n61 VDD1.n60 185
R176 VDD1.n59 VDD1.n58 185
R177 VDD1.n22 VDD1.n21 185
R178 VDD1.n53 VDD1.n52 185
R179 VDD1.n51 VDD1.n50 185
R180 VDD1.n26 VDD1.n25 185
R181 VDD1.n45 VDD1.n44 185
R182 VDD1.n43 VDD1.n42 185
R183 VDD1.n30 VDD1.n29 185
R184 VDD1.n37 VDD1.n36 185
R185 VDD1.n35 VDD1.n34 185
R186 VDD1.n132 VDD1.n131 185
R187 VDD1.n134 VDD1.n133 185
R188 VDD1.n127 VDD1.n126 185
R189 VDD1.n140 VDD1.n139 185
R190 VDD1.n142 VDD1.n141 185
R191 VDD1.n123 VDD1.n122 185
R192 VDD1.n148 VDD1.n147 185
R193 VDD1.n150 VDD1.n149 185
R194 VDD1.n119 VDD1.n118 185
R195 VDD1.n156 VDD1.n155 185
R196 VDD1.n158 VDD1.n157 185
R197 VDD1.n115 VDD1.n114 185
R198 VDD1.n164 VDD1.n163 185
R199 VDD1.n166 VDD1.n165 185
R200 VDD1.n111 VDD1.n110 185
R201 VDD1.n173 VDD1.n172 185
R202 VDD1.n174 VDD1.n109 185
R203 VDD1.n176 VDD1.n175 185
R204 VDD1.n107 VDD1.n106 185
R205 VDD1.n182 VDD1.n181 185
R206 VDD1.n184 VDD1.n183 185
R207 VDD1.n103 VDD1.n102 185
R208 VDD1.n190 VDD1.n189 185
R209 VDD1.n192 VDD1.n191 185
R210 VDD1.n33 VDD1.t2 147.659
R211 VDD1.n130 VDD1.t6 147.659
R212 VDD1.n92 VDD1.n91 104.615
R213 VDD1.n91 VDD1.n3 104.615
R214 VDD1.n84 VDD1.n3 104.615
R215 VDD1.n84 VDD1.n83 104.615
R216 VDD1.n83 VDD1.n7 104.615
R217 VDD1.n12 VDD1.n7 104.615
R218 VDD1.n76 VDD1.n12 104.615
R219 VDD1.n76 VDD1.n75 104.615
R220 VDD1.n75 VDD1.n13 104.615
R221 VDD1.n68 VDD1.n13 104.615
R222 VDD1.n68 VDD1.n67 104.615
R223 VDD1.n67 VDD1.n17 104.615
R224 VDD1.n60 VDD1.n17 104.615
R225 VDD1.n60 VDD1.n59 104.615
R226 VDD1.n59 VDD1.n21 104.615
R227 VDD1.n52 VDD1.n21 104.615
R228 VDD1.n52 VDD1.n51 104.615
R229 VDD1.n51 VDD1.n25 104.615
R230 VDD1.n44 VDD1.n25 104.615
R231 VDD1.n44 VDD1.n43 104.615
R232 VDD1.n43 VDD1.n29 104.615
R233 VDD1.n36 VDD1.n29 104.615
R234 VDD1.n36 VDD1.n35 104.615
R235 VDD1.n133 VDD1.n132 104.615
R236 VDD1.n133 VDD1.n126 104.615
R237 VDD1.n140 VDD1.n126 104.615
R238 VDD1.n141 VDD1.n140 104.615
R239 VDD1.n141 VDD1.n122 104.615
R240 VDD1.n148 VDD1.n122 104.615
R241 VDD1.n149 VDD1.n148 104.615
R242 VDD1.n149 VDD1.n118 104.615
R243 VDD1.n156 VDD1.n118 104.615
R244 VDD1.n157 VDD1.n156 104.615
R245 VDD1.n157 VDD1.n114 104.615
R246 VDD1.n164 VDD1.n114 104.615
R247 VDD1.n165 VDD1.n164 104.615
R248 VDD1.n165 VDD1.n110 104.615
R249 VDD1.n173 VDD1.n110 104.615
R250 VDD1.n174 VDD1.n173 104.615
R251 VDD1.n175 VDD1.n174 104.615
R252 VDD1.n175 VDD1.n106 104.615
R253 VDD1.n182 VDD1.n106 104.615
R254 VDD1.n183 VDD1.n182 104.615
R255 VDD1.n183 VDD1.n102 104.615
R256 VDD1.n190 VDD1.n102 104.615
R257 VDD1.n191 VDD1.n190 104.615
R258 VDD1.n199 VDD1.n198 63.0576
R259 VDD1.n98 VDD1.n97 61.07
R260 VDD1.n197 VDD1.n196 61.0699
R261 VDD1.n201 VDD1.n200 61.0698
R262 VDD1.n201 VDD1.n199 53.7207
R263 VDD1.n35 VDD1.t2 52.3082
R264 VDD1.n132 VDD1.t6 52.3082
R265 VDD1.n98 VDD1.n96 51.9762
R266 VDD1.n197 VDD1.n195 51.9762
R267 VDD1.n34 VDD1.n33 15.6677
R268 VDD1.n131 VDD1.n130 15.6677
R269 VDD1.n10 VDD1.n8 13.1884
R270 VDD1.n176 VDD1.n107 13.1884
R271 VDD1.n82 VDD1.n81 12.8005
R272 VDD1.n78 VDD1.n77 12.8005
R273 VDD1.n37 VDD1.n32 12.8005
R274 VDD1.n134 VDD1.n129 12.8005
R275 VDD1.n177 VDD1.n109 12.8005
R276 VDD1.n181 VDD1.n180 12.8005
R277 VDD1.n85 VDD1.n6 12.0247
R278 VDD1.n74 VDD1.n11 12.0247
R279 VDD1.n38 VDD1.n30 12.0247
R280 VDD1.n135 VDD1.n127 12.0247
R281 VDD1.n172 VDD1.n171 12.0247
R282 VDD1.n184 VDD1.n105 12.0247
R283 VDD1.n86 VDD1.n4 11.249
R284 VDD1.n73 VDD1.n14 11.249
R285 VDD1.n42 VDD1.n41 11.249
R286 VDD1.n139 VDD1.n138 11.249
R287 VDD1.n170 VDD1.n111 11.249
R288 VDD1.n185 VDD1.n103 11.249
R289 VDD1.n90 VDD1.n89 10.4732
R290 VDD1.n70 VDD1.n69 10.4732
R291 VDD1.n45 VDD1.n28 10.4732
R292 VDD1.n142 VDD1.n125 10.4732
R293 VDD1.n167 VDD1.n166 10.4732
R294 VDD1.n189 VDD1.n188 10.4732
R295 VDD1.n93 VDD1.n2 9.69747
R296 VDD1.n66 VDD1.n16 9.69747
R297 VDD1.n46 VDD1.n26 9.69747
R298 VDD1.n143 VDD1.n123 9.69747
R299 VDD1.n163 VDD1.n113 9.69747
R300 VDD1.n192 VDD1.n101 9.69747
R301 VDD1.n96 VDD1.n95 9.45567
R302 VDD1.n195 VDD1.n194 9.45567
R303 VDD1.n20 VDD1.n19 9.3005
R304 VDD1.n63 VDD1.n62 9.3005
R305 VDD1.n65 VDD1.n64 9.3005
R306 VDD1.n16 VDD1.n15 9.3005
R307 VDD1.n71 VDD1.n70 9.3005
R308 VDD1.n73 VDD1.n72 9.3005
R309 VDD1.n11 VDD1.n9 9.3005
R310 VDD1.n79 VDD1.n78 9.3005
R311 VDD1.n95 VDD1.n94 9.3005
R312 VDD1.n2 VDD1.n1 9.3005
R313 VDD1.n89 VDD1.n88 9.3005
R314 VDD1.n87 VDD1.n86 9.3005
R315 VDD1.n6 VDD1.n5 9.3005
R316 VDD1.n81 VDD1.n80 9.3005
R317 VDD1.n57 VDD1.n56 9.3005
R318 VDD1.n55 VDD1.n54 9.3005
R319 VDD1.n24 VDD1.n23 9.3005
R320 VDD1.n49 VDD1.n48 9.3005
R321 VDD1.n47 VDD1.n46 9.3005
R322 VDD1.n28 VDD1.n27 9.3005
R323 VDD1.n41 VDD1.n40 9.3005
R324 VDD1.n39 VDD1.n38 9.3005
R325 VDD1.n32 VDD1.n31 9.3005
R326 VDD1.n194 VDD1.n193 9.3005
R327 VDD1.n101 VDD1.n100 9.3005
R328 VDD1.n188 VDD1.n187 9.3005
R329 VDD1.n186 VDD1.n185 9.3005
R330 VDD1.n105 VDD1.n104 9.3005
R331 VDD1.n180 VDD1.n179 9.3005
R332 VDD1.n152 VDD1.n151 9.3005
R333 VDD1.n121 VDD1.n120 9.3005
R334 VDD1.n146 VDD1.n145 9.3005
R335 VDD1.n144 VDD1.n143 9.3005
R336 VDD1.n125 VDD1.n124 9.3005
R337 VDD1.n138 VDD1.n137 9.3005
R338 VDD1.n136 VDD1.n135 9.3005
R339 VDD1.n129 VDD1.n128 9.3005
R340 VDD1.n154 VDD1.n153 9.3005
R341 VDD1.n117 VDD1.n116 9.3005
R342 VDD1.n160 VDD1.n159 9.3005
R343 VDD1.n162 VDD1.n161 9.3005
R344 VDD1.n113 VDD1.n112 9.3005
R345 VDD1.n168 VDD1.n167 9.3005
R346 VDD1.n170 VDD1.n169 9.3005
R347 VDD1.n171 VDD1.n108 9.3005
R348 VDD1.n178 VDD1.n177 9.3005
R349 VDD1.n94 VDD1.n0 8.92171
R350 VDD1.n65 VDD1.n18 8.92171
R351 VDD1.n50 VDD1.n49 8.92171
R352 VDD1.n147 VDD1.n146 8.92171
R353 VDD1.n162 VDD1.n115 8.92171
R354 VDD1.n193 VDD1.n99 8.92171
R355 VDD1.n62 VDD1.n61 8.14595
R356 VDD1.n53 VDD1.n24 8.14595
R357 VDD1.n150 VDD1.n121 8.14595
R358 VDD1.n159 VDD1.n158 8.14595
R359 VDD1.n58 VDD1.n20 7.3702
R360 VDD1.n54 VDD1.n22 7.3702
R361 VDD1.n151 VDD1.n119 7.3702
R362 VDD1.n155 VDD1.n117 7.3702
R363 VDD1.n58 VDD1.n57 6.59444
R364 VDD1.n57 VDD1.n22 6.59444
R365 VDD1.n154 VDD1.n119 6.59444
R366 VDD1.n155 VDD1.n154 6.59444
R367 VDD1.n61 VDD1.n20 5.81868
R368 VDD1.n54 VDD1.n53 5.81868
R369 VDD1.n151 VDD1.n150 5.81868
R370 VDD1.n158 VDD1.n117 5.81868
R371 VDD1.n96 VDD1.n0 5.04292
R372 VDD1.n62 VDD1.n18 5.04292
R373 VDD1.n50 VDD1.n24 5.04292
R374 VDD1.n147 VDD1.n121 5.04292
R375 VDD1.n159 VDD1.n115 5.04292
R376 VDD1.n195 VDD1.n99 5.04292
R377 VDD1.n33 VDD1.n31 4.38563
R378 VDD1.n130 VDD1.n128 4.38563
R379 VDD1.n94 VDD1.n93 4.26717
R380 VDD1.n66 VDD1.n65 4.26717
R381 VDD1.n49 VDD1.n26 4.26717
R382 VDD1.n146 VDD1.n123 4.26717
R383 VDD1.n163 VDD1.n162 4.26717
R384 VDD1.n193 VDD1.n192 4.26717
R385 VDD1.n90 VDD1.n2 3.49141
R386 VDD1.n69 VDD1.n16 3.49141
R387 VDD1.n46 VDD1.n45 3.49141
R388 VDD1.n143 VDD1.n142 3.49141
R389 VDD1.n166 VDD1.n113 3.49141
R390 VDD1.n189 VDD1.n101 3.49141
R391 VDD1.n89 VDD1.n4 2.71565
R392 VDD1.n70 VDD1.n14 2.71565
R393 VDD1.n42 VDD1.n28 2.71565
R394 VDD1.n139 VDD1.n125 2.71565
R395 VDD1.n167 VDD1.n111 2.71565
R396 VDD1.n188 VDD1.n103 2.71565
R397 VDD1 VDD1.n201 1.98541
R398 VDD1.n86 VDD1.n85 1.93989
R399 VDD1.n74 VDD1.n73 1.93989
R400 VDD1.n41 VDD1.n30 1.93989
R401 VDD1.n138 VDD1.n127 1.93989
R402 VDD1.n172 VDD1.n170 1.93989
R403 VDD1.n185 VDD1.n184 1.93989
R404 VDD1.n82 VDD1.n6 1.16414
R405 VDD1.n77 VDD1.n11 1.16414
R406 VDD1.n38 VDD1.n37 1.16414
R407 VDD1.n135 VDD1.n134 1.16414
R408 VDD1.n171 VDD1.n109 1.16414
R409 VDD1.n181 VDD1.n105 1.16414
R410 VDD1.n200 VDD1.t9 1.12935
R411 VDD1.n200 VDD1.t1 1.12935
R412 VDD1.n97 VDD1.t7 1.12935
R413 VDD1.n97 VDD1.t8 1.12935
R414 VDD1.n198 VDD1.t4 1.12935
R415 VDD1.n198 VDD1.t5 1.12935
R416 VDD1.n196 VDD1.t3 1.12935
R417 VDD1.n196 VDD1.t0 1.12935
R418 VDD1 VDD1.n98 0.739724
R419 VDD1.n199 VDD1.n197 0.626188
R420 VDD1.n81 VDD1.n8 0.388379
R421 VDD1.n78 VDD1.n10 0.388379
R422 VDD1.n34 VDD1.n32 0.388379
R423 VDD1.n131 VDD1.n129 0.388379
R424 VDD1.n177 VDD1.n176 0.388379
R425 VDD1.n180 VDD1.n107 0.388379
R426 VDD1.n95 VDD1.n1 0.155672
R427 VDD1.n88 VDD1.n1 0.155672
R428 VDD1.n88 VDD1.n87 0.155672
R429 VDD1.n87 VDD1.n5 0.155672
R430 VDD1.n80 VDD1.n5 0.155672
R431 VDD1.n80 VDD1.n79 0.155672
R432 VDD1.n79 VDD1.n9 0.155672
R433 VDD1.n72 VDD1.n9 0.155672
R434 VDD1.n72 VDD1.n71 0.155672
R435 VDD1.n71 VDD1.n15 0.155672
R436 VDD1.n64 VDD1.n15 0.155672
R437 VDD1.n64 VDD1.n63 0.155672
R438 VDD1.n63 VDD1.n19 0.155672
R439 VDD1.n56 VDD1.n19 0.155672
R440 VDD1.n56 VDD1.n55 0.155672
R441 VDD1.n55 VDD1.n23 0.155672
R442 VDD1.n48 VDD1.n23 0.155672
R443 VDD1.n48 VDD1.n47 0.155672
R444 VDD1.n47 VDD1.n27 0.155672
R445 VDD1.n40 VDD1.n27 0.155672
R446 VDD1.n40 VDD1.n39 0.155672
R447 VDD1.n39 VDD1.n31 0.155672
R448 VDD1.n136 VDD1.n128 0.155672
R449 VDD1.n137 VDD1.n136 0.155672
R450 VDD1.n137 VDD1.n124 0.155672
R451 VDD1.n144 VDD1.n124 0.155672
R452 VDD1.n145 VDD1.n144 0.155672
R453 VDD1.n145 VDD1.n120 0.155672
R454 VDD1.n152 VDD1.n120 0.155672
R455 VDD1.n153 VDD1.n152 0.155672
R456 VDD1.n153 VDD1.n116 0.155672
R457 VDD1.n160 VDD1.n116 0.155672
R458 VDD1.n161 VDD1.n160 0.155672
R459 VDD1.n161 VDD1.n112 0.155672
R460 VDD1.n168 VDD1.n112 0.155672
R461 VDD1.n169 VDD1.n168 0.155672
R462 VDD1.n169 VDD1.n108 0.155672
R463 VDD1.n178 VDD1.n108 0.155672
R464 VDD1.n179 VDD1.n178 0.155672
R465 VDD1.n179 VDD1.n104 0.155672
R466 VDD1.n186 VDD1.n104 0.155672
R467 VDD1.n187 VDD1.n186 0.155672
R468 VDD1.n187 VDD1.n100 0.155672
R469 VDD1.n194 VDD1.n100 0.155672
R470 VTAIL.n400 VTAIL.n308 289.615
R471 VTAIL.n94 VTAIL.n2 289.615
R472 VTAIL.n302 VTAIL.n210 289.615
R473 VTAIL.n200 VTAIL.n108 289.615
R474 VTAIL.n341 VTAIL.n340 185
R475 VTAIL.n343 VTAIL.n342 185
R476 VTAIL.n336 VTAIL.n335 185
R477 VTAIL.n349 VTAIL.n348 185
R478 VTAIL.n351 VTAIL.n350 185
R479 VTAIL.n332 VTAIL.n331 185
R480 VTAIL.n357 VTAIL.n356 185
R481 VTAIL.n359 VTAIL.n358 185
R482 VTAIL.n328 VTAIL.n327 185
R483 VTAIL.n365 VTAIL.n364 185
R484 VTAIL.n367 VTAIL.n366 185
R485 VTAIL.n324 VTAIL.n323 185
R486 VTAIL.n373 VTAIL.n372 185
R487 VTAIL.n375 VTAIL.n374 185
R488 VTAIL.n320 VTAIL.n319 185
R489 VTAIL.n382 VTAIL.n381 185
R490 VTAIL.n383 VTAIL.n318 185
R491 VTAIL.n385 VTAIL.n384 185
R492 VTAIL.n316 VTAIL.n315 185
R493 VTAIL.n391 VTAIL.n390 185
R494 VTAIL.n393 VTAIL.n392 185
R495 VTAIL.n312 VTAIL.n311 185
R496 VTAIL.n399 VTAIL.n398 185
R497 VTAIL.n401 VTAIL.n400 185
R498 VTAIL.n35 VTAIL.n34 185
R499 VTAIL.n37 VTAIL.n36 185
R500 VTAIL.n30 VTAIL.n29 185
R501 VTAIL.n43 VTAIL.n42 185
R502 VTAIL.n45 VTAIL.n44 185
R503 VTAIL.n26 VTAIL.n25 185
R504 VTAIL.n51 VTAIL.n50 185
R505 VTAIL.n53 VTAIL.n52 185
R506 VTAIL.n22 VTAIL.n21 185
R507 VTAIL.n59 VTAIL.n58 185
R508 VTAIL.n61 VTAIL.n60 185
R509 VTAIL.n18 VTAIL.n17 185
R510 VTAIL.n67 VTAIL.n66 185
R511 VTAIL.n69 VTAIL.n68 185
R512 VTAIL.n14 VTAIL.n13 185
R513 VTAIL.n76 VTAIL.n75 185
R514 VTAIL.n77 VTAIL.n12 185
R515 VTAIL.n79 VTAIL.n78 185
R516 VTAIL.n10 VTAIL.n9 185
R517 VTAIL.n85 VTAIL.n84 185
R518 VTAIL.n87 VTAIL.n86 185
R519 VTAIL.n6 VTAIL.n5 185
R520 VTAIL.n93 VTAIL.n92 185
R521 VTAIL.n95 VTAIL.n94 185
R522 VTAIL.n303 VTAIL.n302 185
R523 VTAIL.n301 VTAIL.n300 185
R524 VTAIL.n214 VTAIL.n213 185
R525 VTAIL.n295 VTAIL.n294 185
R526 VTAIL.n293 VTAIL.n292 185
R527 VTAIL.n218 VTAIL.n217 185
R528 VTAIL.n222 VTAIL.n220 185
R529 VTAIL.n287 VTAIL.n286 185
R530 VTAIL.n285 VTAIL.n284 185
R531 VTAIL.n224 VTAIL.n223 185
R532 VTAIL.n279 VTAIL.n278 185
R533 VTAIL.n277 VTAIL.n276 185
R534 VTAIL.n228 VTAIL.n227 185
R535 VTAIL.n271 VTAIL.n270 185
R536 VTAIL.n269 VTAIL.n268 185
R537 VTAIL.n232 VTAIL.n231 185
R538 VTAIL.n263 VTAIL.n262 185
R539 VTAIL.n261 VTAIL.n260 185
R540 VTAIL.n236 VTAIL.n235 185
R541 VTAIL.n255 VTAIL.n254 185
R542 VTAIL.n253 VTAIL.n252 185
R543 VTAIL.n240 VTAIL.n239 185
R544 VTAIL.n247 VTAIL.n246 185
R545 VTAIL.n245 VTAIL.n244 185
R546 VTAIL.n201 VTAIL.n200 185
R547 VTAIL.n199 VTAIL.n198 185
R548 VTAIL.n112 VTAIL.n111 185
R549 VTAIL.n193 VTAIL.n192 185
R550 VTAIL.n191 VTAIL.n190 185
R551 VTAIL.n116 VTAIL.n115 185
R552 VTAIL.n120 VTAIL.n118 185
R553 VTAIL.n185 VTAIL.n184 185
R554 VTAIL.n183 VTAIL.n182 185
R555 VTAIL.n122 VTAIL.n121 185
R556 VTAIL.n177 VTAIL.n176 185
R557 VTAIL.n175 VTAIL.n174 185
R558 VTAIL.n126 VTAIL.n125 185
R559 VTAIL.n169 VTAIL.n168 185
R560 VTAIL.n167 VTAIL.n166 185
R561 VTAIL.n130 VTAIL.n129 185
R562 VTAIL.n161 VTAIL.n160 185
R563 VTAIL.n159 VTAIL.n158 185
R564 VTAIL.n134 VTAIL.n133 185
R565 VTAIL.n153 VTAIL.n152 185
R566 VTAIL.n151 VTAIL.n150 185
R567 VTAIL.n138 VTAIL.n137 185
R568 VTAIL.n145 VTAIL.n144 185
R569 VTAIL.n143 VTAIL.n142 185
R570 VTAIL.n339 VTAIL.t7 147.659
R571 VTAIL.n33 VTAIL.t17 147.659
R572 VTAIL.n243 VTAIL.t13 147.659
R573 VTAIL.n141 VTAIL.t5 147.659
R574 VTAIL.n342 VTAIL.n341 104.615
R575 VTAIL.n342 VTAIL.n335 104.615
R576 VTAIL.n349 VTAIL.n335 104.615
R577 VTAIL.n350 VTAIL.n349 104.615
R578 VTAIL.n350 VTAIL.n331 104.615
R579 VTAIL.n357 VTAIL.n331 104.615
R580 VTAIL.n358 VTAIL.n357 104.615
R581 VTAIL.n358 VTAIL.n327 104.615
R582 VTAIL.n365 VTAIL.n327 104.615
R583 VTAIL.n366 VTAIL.n365 104.615
R584 VTAIL.n366 VTAIL.n323 104.615
R585 VTAIL.n373 VTAIL.n323 104.615
R586 VTAIL.n374 VTAIL.n373 104.615
R587 VTAIL.n374 VTAIL.n319 104.615
R588 VTAIL.n382 VTAIL.n319 104.615
R589 VTAIL.n383 VTAIL.n382 104.615
R590 VTAIL.n384 VTAIL.n383 104.615
R591 VTAIL.n384 VTAIL.n315 104.615
R592 VTAIL.n391 VTAIL.n315 104.615
R593 VTAIL.n392 VTAIL.n391 104.615
R594 VTAIL.n392 VTAIL.n311 104.615
R595 VTAIL.n399 VTAIL.n311 104.615
R596 VTAIL.n400 VTAIL.n399 104.615
R597 VTAIL.n36 VTAIL.n35 104.615
R598 VTAIL.n36 VTAIL.n29 104.615
R599 VTAIL.n43 VTAIL.n29 104.615
R600 VTAIL.n44 VTAIL.n43 104.615
R601 VTAIL.n44 VTAIL.n25 104.615
R602 VTAIL.n51 VTAIL.n25 104.615
R603 VTAIL.n52 VTAIL.n51 104.615
R604 VTAIL.n52 VTAIL.n21 104.615
R605 VTAIL.n59 VTAIL.n21 104.615
R606 VTAIL.n60 VTAIL.n59 104.615
R607 VTAIL.n60 VTAIL.n17 104.615
R608 VTAIL.n67 VTAIL.n17 104.615
R609 VTAIL.n68 VTAIL.n67 104.615
R610 VTAIL.n68 VTAIL.n13 104.615
R611 VTAIL.n76 VTAIL.n13 104.615
R612 VTAIL.n77 VTAIL.n76 104.615
R613 VTAIL.n78 VTAIL.n77 104.615
R614 VTAIL.n78 VTAIL.n9 104.615
R615 VTAIL.n85 VTAIL.n9 104.615
R616 VTAIL.n86 VTAIL.n85 104.615
R617 VTAIL.n86 VTAIL.n5 104.615
R618 VTAIL.n93 VTAIL.n5 104.615
R619 VTAIL.n94 VTAIL.n93 104.615
R620 VTAIL.n302 VTAIL.n301 104.615
R621 VTAIL.n301 VTAIL.n213 104.615
R622 VTAIL.n294 VTAIL.n213 104.615
R623 VTAIL.n294 VTAIL.n293 104.615
R624 VTAIL.n293 VTAIL.n217 104.615
R625 VTAIL.n222 VTAIL.n217 104.615
R626 VTAIL.n286 VTAIL.n222 104.615
R627 VTAIL.n286 VTAIL.n285 104.615
R628 VTAIL.n285 VTAIL.n223 104.615
R629 VTAIL.n278 VTAIL.n223 104.615
R630 VTAIL.n278 VTAIL.n277 104.615
R631 VTAIL.n277 VTAIL.n227 104.615
R632 VTAIL.n270 VTAIL.n227 104.615
R633 VTAIL.n270 VTAIL.n269 104.615
R634 VTAIL.n269 VTAIL.n231 104.615
R635 VTAIL.n262 VTAIL.n231 104.615
R636 VTAIL.n262 VTAIL.n261 104.615
R637 VTAIL.n261 VTAIL.n235 104.615
R638 VTAIL.n254 VTAIL.n235 104.615
R639 VTAIL.n254 VTAIL.n253 104.615
R640 VTAIL.n253 VTAIL.n239 104.615
R641 VTAIL.n246 VTAIL.n239 104.615
R642 VTAIL.n246 VTAIL.n245 104.615
R643 VTAIL.n200 VTAIL.n199 104.615
R644 VTAIL.n199 VTAIL.n111 104.615
R645 VTAIL.n192 VTAIL.n111 104.615
R646 VTAIL.n192 VTAIL.n191 104.615
R647 VTAIL.n191 VTAIL.n115 104.615
R648 VTAIL.n120 VTAIL.n115 104.615
R649 VTAIL.n184 VTAIL.n120 104.615
R650 VTAIL.n184 VTAIL.n183 104.615
R651 VTAIL.n183 VTAIL.n121 104.615
R652 VTAIL.n176 VTAIL.n121 104.615
R653 VTAIL.n176 VTAIL.n175 104.615
R654 VTAIL.n175 VTAIL.n125 104.615
R655 VTAIL.n168 VTAIL.n125 104.615
R656 VTAIL.n168 VTAIL.n167 104.615
R657 VTAIL.n167 VTAIL.n129 104.615
R658 VTAIL.n160 VTAIL.n129 104.615
R659 VTAIL.n160 VTAIL.n159 104.615
R660 VTAIL.n159 VTAIL.n133 104.615
R661 VTAIL.n152 VTAIL.n133 104.615
R662 VTAIL.n152 VTAIL.n151 104.615
R663 VTAIL.n151 VTAIL.n137 104.615
R664 VTAIL.n144 VTAIL.n137 104.615
R665 VTAIL.n144 VTAIL.n143 104.615
R666 VTAIL.n341 VTAIL.t7 52.3082
R667 VTAIL.n35 VTAIL.t17 52.3082
R668 VTAIL.n245 VTAIL.t13 52.3082
R669 VTAIL.n143 VTAIL.t5 52.3082
R670 VTAIL.n209 VTAIL.n208 44.3912
R671 VTAIL.n207 VTAIL.n206 44.3912
R672 VTAIL.n107 VTAIL.n106 44.3912
R673 VTAIL.n105 VTAIL.n104 44.3912
R674 VTAIL.n407 VTAIL.n406 44.3911
R675 VTAIL.n1 VTAIL.n0 44.3911
R676 VTAIL.n101 VTAIL.n100 44.3911
R677 VTAIL.n103 VTAIL.n102 44.3911
R678 VTAIL.n105 VTAIL.n103 32.9358
R679 VTAIL.n405 VTAIL.n404 32.5732
R680 VTAIL.n99 VTAIL.n98 32.5732
R681 VTAIL.n307 VTAIL.n306 32.5732
R682 VTAIL.n205 VTAIL.n204 32.5732
R683 VTAIL.n405 VTAIL.n307 30.2117
R684 VTAIL.n340 VTAIL.n339 15.6677
R685 VTAIL.n34 VTAIL.n33 15.6677
R686 VTAIL.n244 VTAIL.n243 15.6677
R687 VTAIL.n142 VTAIL.n141 15.6677
R688 VTAIL.n385 VTAIL.n316 13.1884
R689 VTAIL.n79 VTAIL.n10 13.1884
R690 VTAIL.n220 VTAIL.n218 13.1884
R691 VTAIL.n118 VTAIL.n116 13.1884
R692 VTAIL.n343 VTAIL.n338 12.8005
R693 VTAIL.n386 VTAIL.n318 12.8005
R694 VTAIL.n390 VTAIL.n389 12.8005
R695 VTAIL.n37 VTAIL.n32 12.8005
R696 VTAIL.n80 VTAIL.n12 12.8005
R697 VTAIL.n84 VTAIL.n83 12.8005
R698 VTAIL.n292 VTAIL.n291 12.8005
R699 VTAIL.n288 VTAIL.n287 12.8005
R700 VTAIL.n247 VTAIL.n242 12.8005
R701 VTAIL.n190 VTAIL.n189 12.8005
R702 VTAIL.n186 VTAIL.n185 12.8005
R703 VTAIL.n145 VTAIL.n140 12.8005
R704 VTAIL.n344 VTAIL.n336 12.0247
R705 VTAIL.n381 VTAIL.n380 12.0247
R706 VTAIL.n393 VTAIL.n314 12.0247
R707 VTAIL.n38 VTAIL.n30 12.0247
R708 VTAIL.n75 VTAIL.n74 12.0247
R709 VTAIL.n87 VTAIL.n8 12.0247
R710 VTAIL.n295 VTAIL.n216 12.0247
R711 VTAIL.n284 VTAIL.n221 12.0247
R712 VTAIL.n248 VTAIL.n240 12.0247
R713 VTAIL.n193 VTAIL.n114 12.0247
R714 VTAIL.n182 VTAIL.n119 12.0247
R715 VTAIL.n146 VTAIL.n138 12.0247
R716 VTAIL.n348 VTAIL.n347 11.249
R717 VTAIL.n379 VTAIL.n320 11.249
R718 VTAIL.n394 VTAIL.n312 11.249
R719 VTAIL.n42 VTAIL.n41 11.249
R720 VTAIL.n73 VTAIL.n14 11.249
R721 VTAIL.n88 VTAIL.n6 11.249
R722 VTAIL.n296 VTAIL.n214 11.249
R723 VTAIL.n283 VTAIL.n224 11.249
R724 VTAIL.n252 VTAIL.n251 11.249
R725 VTAIL.n194 VTAIL.n112 11.249
R726 VTAIL.n181 VTAIL.n122 11.249
R727 VTAIL.n150 VTAIL.n149 11.249
R728 VTAIL.n351 VTAIL.n334 10.4732
R729 VTAIL.n376 VTAIL.n375 10.4732
R730 VTAIL.n398 VTAIL.n397 10.4732
R731 VTAIL.n45 VTAIL.n28 10.4732
R732 VTAIL.n70 VTAIL.n69 10.4732
R733 VTAIL.n92 VTAIL.n91 10.4732
R734 VTAIL.n300 VTAIL.n299 10.4732
R735 VTAIL.n280 VTAIL.n279 10.4732
R736 VTAIL.n255 VTAIL.n238 10.4732
R737 VTAIL.n198 VTAIL.n197 10.4732
R738 VTAIL.n178 VTAIL.n177 10.4732
R739 VTAIL.n153 VTAIL.n136 10.4732
R740 VTAIL.n352 VTAIL.n332 9.69747
R741 VTAIL.n372 VTAIL.n322 9.69747
R742 VTAIL.n401 VTAIL.n310 9.69747
R743 VTAIL.n46 VTAIL.n26 9.69747
R744 VTAIL.n66 VTAIL.n16 9.69747
R745 VTAIL.n95 VTAIL.n4 9.69747
R746 VTAIL.n303 VTAIL.n212 9.69747
R747 VTAIL.n276 VTAIL.n226 9.69747
R748 VTAIL.n256 VTAIL.n236 9.69747
R749 VTAIL.n201 VTAIL.n110 9.69747
R750 VTAIL.n174 VTAIL.n124 9.69747
R751 VTAIL.n154 VTAIL.n134 9.69747
R752 VTAIL.n404 VTAIL.n403 9.45567
R753 VTAIL.n98 VTAIL.n97 9.45567
R754 VTAIL.n306 VTAIL.n305 9.45567
R755 VTAIL.n204 VTAIL.n203 9.45567
R756 VTAIL.n403 VTAIL.n402 9.3005
R757 VTAIL.n310 VTAIL.n309 9.3005
R758 VTAIL.n397 VTAIL.n396 9.3005
R759 VTAIL.n395 VTAIL.n394 9.3005
R760 VTAIL.n314 VTAIL.n313 9.3005
R761 VTAIL.n389 VTAIL.n388 9.3005
R762 VTAIL.n361 VTAIL.n360 9.3005
R763 VTAIL.n330 VTAIL.n329 9.3005
R764 VTAIL.n355 VTAIL.n354 9.3005
R765 VTAIL.n353 VTAIL.n352 9.3005
R766 VTAIL.n334 VTAIL.n333 9.3005
R767 VTAIL.n347 VTAIL.n346 9.3005
R768 VTAIL.n345 VTAIL.n344 9.3005
R769 VTAIL.n338 VTAIL.n337 9.3005
R770 VTAIL.n363 VTAIL.n362 9.3005
R771 VTAIL.n326 VTAIL.n325 9.3005
R772 VTAIL.n369 VTAIL.n368 9.3005
R773 VTAIL.n371 VTAIL.n370 9.3005
R774 VTAIL.n322 VTAIL.n321 9.3005
R775 VTAIL.n377 VTAIL.n376 9.3005
R776 VTAIL.n379 VTAIL.n378 9.3005
R777 VTAIL.n380 VTAIL.n317 9.3005
R778 VTAIL.n387 VTAIL.n386 9.3005
R779 VTAIL.n97 VTAIL.n96 9.3005
R780 VTAIL.n4 VTAIL.n3 9.3005
R781 VTAIL.n91 VTAIL.n90 9.3005
R782 VTAIL.n89 VTAIL.n88 9.3005
R783 VTAIL.n8 VTAIL.n7 9.3005
R784 VTAIL.n83 VTAIL.n82 9.3005
R785 VTAIL.n55 VTAIL.n54 9.3005
R786 VTAIL.n24 VTAIL.n23 9.3005
R787 VTAIL.n49 VTAIL.n48 9.3005
R788 VTAIL.n47 VTAIL.n46 9.3005
R789 VTAIL.n28 VTAIL.n27 9.3005
R790 VTAIL.n41 VTAIL.n40 9.3005
R791 VTAIL.n39 VTAIL.n38 9.3005
R792 VTAIL.n32 VTAIL.n31 9.3005
R793 VTAIL.n57 VTAIL.n56 9.3005
R794 VTAIL.n20 VTAIL.n19 9.3005
R795 VTAIL.n63 VTAIL.n62 9.3005
R796 VTAIL.n65 VTAIL.n64 9.3005
R797 VTAIL.n16 VTAIL.n15 9.3005
R798 VTAIL.n71 VTAIL.n70 9.3005
R799 VTAIL.n73 VTAIL.n72 9.3005
R800 VTAIL.n74 VTAIL.n11 9.3005
R801 VTAIL.n81 VTAIL.n80 9.3005
R802 VTAIL.n230 VTAIL.n229 9.3005
R803 VTAIL.n273 VTAIL.n272 9.3005
R804 VTAIL.n275 VTAIL.n274 9.3005
R805 VTAIL.n226 VTAIL.n225 9.3005
R806 VTAIL.n281 VTAIL.n280 9.3005
R807 VTAIL.n283 VTAIL.n282 9.3005
R808 VTAIL.n221 VTAIL.n219 9.3005
R809 VTAIL.n289 VTAIL.n288 9.3005
R810 VTAIL.n305 VTAIL.n304 9.3005
R811 VTAIL.n212 VTAIL.n211 9.3005
R812 VTAIL.n299 VTAIL.n298 9.3005
R813 VTAIL.n297 VTAIL.n296 9.3005
R814 VTAIL.n216 VTAIL.n215 9.3005
R815 VTAIL.n291 VTAIL.n290 9.3005
R816 VTAIL.n267 VTAIL.n266 9.3005
R817 VTAIL.n265 VTAIL.n264 9.3005
R818 VTAIL.n234 VTAIL.n233 9.3005
R819 VTAIL.n259 VTAIL.n258 9.3005
R820 VTAIL.n257 VTAIL.n256 9.3005
R821 VTAIL.n238 VTAIL.n237 9.3005
R822 VTAIL.n251 VTAIL.n250 9.3005
R823 VTAIL.n249 VTAIL.n248 9.3005
R824 VTAIL.n242 VTAIL.n241 9.3005
R825 VTAIL.n128 VTAIL.n127 9.3005
R826 VTAIL.n171 VTAIL.n170 9.3005
R827 VTAIL.n173 VTAIL.n172 9.3005
R828 VTAIL.n124 VTAIL.n123 9.3005
R829 VTAIL.n179 VTAIL.n178 9.3005
R830 VTAIL.n181 VTAIL.n180 9.3005
R831 VTAIL.n119 VTAIL.n117 9.3005
R832 VTAIL.n187 VTAIL.n186 9.3005
R833 VTAIL.n203 VTAIL.n202 9.3005
R834 VTAIL.n110 VTAIL.n109 9.3005
R835 VTAIL.n197 VTAIL.n196 9.3005
R836 VTAIL.n195 VTAIL.n194 9.3005
R837 VTAIL.n114 VTAIL.n113 9.3005
R838 VTAIL.n189 VTAIL.n188 9.3005
R839 VTAIL.n165 VTAIL.n164 9.3005
R840 VTAIL.n163 VTAIL.n162 9.3005
R841 VTAIL.n132 VTAIL.n131 9.3005
R842 VTAIL.n157 VTAIL.n156 9.3005
R843 VTAIL.n155 VTAIL.n154 9.3005
R844 VTAIL.n136 VTAIL.n135 9.3005
R845 VTAIL.n149 VTAIL.n148 9.3005
R846 VTAIL.n147 VTAIL.n146 9.3005
R847 VTAIL.n140 VTAIL.n139 9.3005
R848 VTAIL.n356 VTAIL.n355 8.92171
R849 VTAIL.n371 VTAIL.n324 8.92171
R850 VTAIL.n402 VTAIL.n308 8.92171
R851 VTAIL.n50 VTAIL.n49 8.92171
R852 VTAIL.n65 VTAIL.n18 8.92171
R853 VTAIL.n96 VTAIL.n2 8.92171
R854 VTAIL.n304 VTAIL.n210 8.92171
R855 VTAIL.n275 VTAIL.n228 8.92171
R856 VTAIL.n260 VTAIL.n259 8.92171
R857 VTAIL.n202 VTAIL.n108 8.92171
R858 VTAIL.n173 VTAIL.n126 8.92171
R859 VTAIL.n158 VTAIL.n157 8.92171
R860 VTAIL.n359 VTAIL.n330 8.14595
R861 VTAIL.n368 VTAIL.n367 8.14595
R862 VTAIL.n53 VTAIL.n24 8.14595
R863 VTAIL.n62 VTAIL.n61 8.14595
R864 VTAIL.n272 VTAIL.n271 8.14595
R865 VTAIL.n263 VTAIL.n234 8.14595
R866 VTAIL.n170 VTAIL.n169 8.14595
R867 VTAIL.n161 VTAIL.n132 8.14595
R868 VTAIL.n360 VTAIL.n328 7.3702
R869 VTAIL.n364 VTAIL.n326 7.3702
R870 VTAIL.n54 VTAIL.n22 7.3702
R871 VTAIL.n58 VTAIL.n20 7.3702
R872 VTAIL.n268 VTAIL.n230 7.3702
R873 VTAIL.n264 VTAIL.n232 7.3702
R874 VTAIL.n166 VTAIL.n128 7.3702
R875 VTAIL.n162 VTAIL.n130 7.3702
R876 VTAIL.n363 VTAIL.n328 6.59444
R877 VTAIL.n364 VTAIL.n363 6.59444
R878 VTAIL.n57 VTAIL.n22 6.59444
R879 VTAIL.n58 VTAIL.n57 6.59444
R880 VTAIL.n268 VTAIL.n267 6.59444
R881 VTAIL.n267 VTAIL.n232 6.59444
R882 VTAIL.n166 VTAIL.n165 6.59444
R883 VTAIL.n165 VTAIL.n130 6.59444
R884 VTAIL.n360 VTAIL.n359 5.81868
R885 VTAIL.n367 VTAIL.n326 5.81868
R886 VTAIL.n54 VTAIL.n53 5.81868
R887 VTAIL.n61 VTAIL.n20 5.81868
R888 VTAIL.n271 VTAIL.n230 5.81868
R889 VTAIL.n264 VTAIL.n263 5.81868
R890 VTAIL.n169 VTAIL.n128 5.81868
R891 VTAIL.n162 VTAIL.n161 5.81868
R892 VTAIL.n356 VTAIL.n330 5.04292
R893 VTAIL.n368 VTAIL.n324 5.04292
R894 VTAIL.n404 VTAIL.n308 5.04292
R895 VTAIL.n50 VTAIL.n24 5.04292
R896 VTAIL.n62 VTAIL.n18 5.04292
R897 VTAIL.n98 VTAIL.n2 5.04292
R898 VTAIL.n306 VTAIL.n210 5.04292
R899 VTAIL.n272 VTAIL.n228 5.04292
R900 VTAIL.n260 VTAIL.n234 5.04292
R901 VTAIL.n204 VTAIL.n108 5.04292
R902 VTAIL.n170 VTAIL.n126 5.04292
R903 VTAIL.n158 VTAIL.n132 5.04292
R904 VTAIL.n339 VTAIL.n337 4.38563
R905 VTAIL.n33 VTAIL.n31 4.38563
R906 VTAIL.n243 VTAIL.n241 4.38563
R907 VTAIL.n141 VTAIL.n139 4.38563
R908 VTAIL.n355 VTAIL.n332 4.26717
R909 VTAIL.n372 VTAIL.n371 4.26717
R910 VTAIL.n402 VTAIL.n401 4.26717
R911 VTAIL.n49 VTAIL.n26 4.26717
R912 VTAIL.n66 VTAIL.n65 4.26717
R913 VTAIL.n96 VTAIL.n95 4.26717
R914 VTAIL.n304 VTAIL.n303 4.26717
R915 VTAIL.n276 VTAIL.n275 4.26717
R916 VTAIL.n259 VTAIL.n236 4.26717
R917 VTAIL.n202 VTAIL.n201 4.26717
R918 VTAIL.n174 VTAIL.n173 4.26717
R919 VTAIL.n157 VTAIL.n134 4.26717
R920 VTAIL.n352 VTAIL.n351 3.49141
R921 VTAIL.n375 VTAIL.n322 3.49141
R922 VTAIL.n398 VTAIL.n310 3.49141
R923 VTAIL.n46 VTAIL.n45 3.49141
R924 VTAIL.n69 VTAIL.n16 3.49141
R925 VTAIL.n92 VTAIL.n4 3.49141
R926 VTAIL.n300 VTAIL.n212 3.49141
R927 VTAIL.n279 VTAIL.n226 3.49141
R928 VTAIL.n256 VTAIL.n255 3.49141
R929 VTAIL.n198 VTAIL.n110 3.49141
R930 VTAIL.n177 VTAIL.n124 3.49141
R931 VTAIL.n154 VTAIL.n153 3.49141
R932 VTAIL.n107 VTAIL.n105 2.72464
R933 VTAIL.n205 VTAIL.n107 2.72464
R934 VTAIL.n209 VTAIL.n207 2.72464
R935 VTAIL.n307 VTAIL.n209 2.72464
R936 VTAIL.n103 VTAIL.n101 2.72464
R937 VTAIL.n101 VTAIL.n99 2.72464
R938 VTAIL.n407 VTAIL.n405 2.72464
R939 VTAIL.n348 VTAIL.n334 2.71565
R940 VTAIL.n376 VTAIL.n320 2.71565
R941 VTAIL.n397 VTAIL.n312 2.71565
R942 VTAIL.n42 VTAIL.n28 2.71565
R943 VTAIL.n70 VTAIL.n14 2.71565
R944 VTAIL.n91 VTAIL.n6 2.71565
R945 VTAIL.n299 VTAIL.n214 2.71565
R946 VTAIL.n280 VTAIL.n224 2.71565
R947 VTAIL.n252 VTAIL.n238 2.71565
R948 VTAIL.n197 VTAIL.n112 2.71565
R949 VTAIL.n178 VTAIL.n122 2.71565
R950 VTAIL.n150 VTAIL.n136 2.71565
R951 VTAIL VTAIL.n1 2.10179
R952 VTAIL.n347 VTAIL.n336 1.93989
R953 VTAIL.n381 VTAIL.n379 1.93989
R954 VTAIL.n394 VTAIL.n393 1.93989
R955 VTAIL.n41 VTAIL.n30 1.93989
R956 VTAIL.n75 VTAIL.n73 1.93989
R957 VTAIL.n88 VTAIL.n87 1.93989
R958 VTAIL.n296 VTAIL.n295 1.93989
R959 VTAIL.n284 VTAIL.n283 1.93989
R960 VTAIL.n251 VTAIL.n240 1.93989
R961 VTAIL.n194 VTAIL.n193 1.93989
R962 VTAIL.n182 VTAIL.n181 1.93989
R963 VTAIL.n149 VTAIL.n138 1.93989
R964 VTAIL.n207 VTAIL.n205 1.8324
R965 VTAIL.n99 VTAIL.n1 1.8324
R966 VTAIL.n344 VTAIL.n343 1.16414
R967 VTAIL.n380 VTAIL.n318 1.16414
R968 VTAIL.n390 VTAIL.n314 1.16414
R969 VTAIL.n38 VTAIL.n37 1.16414
R970 VTAIL.n74 VTAIL.n12 1.16414
R971 VTAIL.n84 VTAIL.n8 1.16414
R972 VTAIL.n292 VTAIL.n216 1.16414
R973 VTAIL.n287 VTAIL.n221 1.16414
R974 VTAIL.n248 VTAIL.n247 1.16414
R975 VTAIL.n190 VTAIL.n114 1.16414
R976 VTAIL.n185 VTAIL.n119 1.16414
R977 VTAIL.n146 VTAIL.n145 1.16414
R978 VTAIL.n406 VTAIL.t6 1.12935
R979 VTAIL.n406 VTAIL.t1 1.12935
R980 VTAIL.n0 VTAIL.t0 1.12935
R981 VTAIL.n0 VTAIL.t3 1.12935
R982 VTAIL.n100 VTAIL.t12 1.12935
R983 VTAIL.n100 VTAIL.t16 1.12935
R984 VTAIL.n102 VTAIL.t14 1.12935
R985 VTAIL.n102 VTAIL.t11 1.12935
R986 VTAIL.n208 VTAIL.t18 1.12935
R987 VTAIL.n208 VTAIL.t19 1.12935
R988 VTAIL.n206 VTAIL.t10 1.12935
R989 VTAIL.n206 VTAIL.t15 1.12935
R990 VTAIL.n106 VTAIL.t8 1.12935
R991 VTAIL.n106 VTAIL.t4 1.12935
R992 VTAIL.n104 VTAIL.t9 1.12935
R993 VTAIL.n104 VTAIL.t2 1.12935
R994 VTAIL VTAIL.n407 0.623345
R995 VTAIL.n340 VTAIL.n338 0.388379
R996 VTAIL.n386 VTAIL.n385 0.388379
R997 VTAIL.n389 VTAIL.n316 0.388379
R998 VTAIL.n34 VTAIL.n32 0.388379
R999 VTAIL.n80 VTAIL.n79 0.388379
R1000 VTAIL.n83 VTAIL.n10 0.388379
R1001 VTAIL.n291 VTAIL.n218 0.388379
R1002 VTAIL.n288 VTAIL.n220 0.388379
R1003 VTAIL.n244 VTAIL.n242 0.388379
R1004 VTAIL.n189 VTAIL.n116 0.388379
R1005 VTAIL.n186 VTAIL.n118 0.388379
R1006 VTAIL.n142 VTAIL.n140 0.388379
R1007 VTAIL.n345 VTAIL.n337 0.155672
R1008 VTAIL.n346 VTAIL.n345 0.155672
R1009 VTAIL.n346 VTAIL.n333 0.155672
R1010 VTAIL.n353 VTAIL.n333 0.155672
R1011 VTAIL.n354 VTAIL.n353 0.155672
R1012 VTAIL.n354 VTAIL.n329 0.155672
R1013 VTAIL.n361 VTAIL.n329 0.155672
R1014 VTAIL.n362 VTAIL.n361 0.155672
R1015 VTAIL.n362 VTAIL.n325 0.155672
R1016 VTAIL.n369 VTAIL.n325 0.155672
R1017 VTAIL.n370 VTAIL.n369 0.155672
R1018 VTAIL.n370 VTAIL.n321 0.155672
R1019 VTAIL.n377 VTAIL.n321 0.155672
R1020 VTAIL.n378 VTAIL.n377 0.155672
R1021 VTAIL.n378 VTAIL.n317 0.155672
R1022 VTAIL.n387 VTAIL.n317 0.155672
R1023 VTAIL.n388 VTAIL.n387 0.155672
R1024 VTAIL.n388 VTAIL.n313 0.155672
R1025 VTAIL.n395 VTAIL.n313 0.155672
R1026 VTAIL.n396 VTAIL.n395 0.155672
R1027 VTAIL.n396 VTAIL.n309 0.155672
R1028 VTAIL.n403 VTAIL.n309 0.155672
R1029 VTAIL.n39 VTAIL.n31 0.155672
R1030 VTAIL.n40 VTAIL.n39 0.155672
R1031 VTAIL.n40 VTAIL.n27 0.155672
R1032 VTAIL.n47 VTAIL.n27 0.155672
R1033 VTAIL.n48 VTAIL.n47 0.155672
R1034 VTAIL.n48 VTAIL.n23 0.155672
R1035 VTAIL.n55 VTAIL.n23 0.155672
R1036 VTAIL.n56 VTAIL.n55 0.155672
R1037 VTAIL.n56 VTAIL.n19 0.155672
R1038 VTAIL.n63 VTAIL.n19 0.155672
R1039 VTAIL.n64 VTAIL.n63 0.155672
R1040 VTAIL.n64 VTAIL.n15 0.155672
R1041 VTAIL.n71 VTAIL.n15 0.155672
R1042 VTAIL.n72 VTAIL.n71 0.155672
R1043 VTAIL.n72 VTAIL.n11 0.155672
R1044 VTAIL.n81 VTAIL.n11 0.155672
R1045 VTAIL.n82 VTAIL.n81 0.155672
R1046 VTAIL.n82 VTAIL.n7 0.155672
R1047 VTAIL.n89 VTAIL.n7 0.155672
R1048 VTAIL.n90 VTAIL.n89 0.155672
R1049 VTAIL.n90 VTAIL.n3 0.155672
R1050 VTAIL.n97 VTAIL.n3 0.155672
R1051 VTAIL.n305 VTAIL.n211 0.155672
R1052 VTAIL.n298 VTAIL.n211 0.155672
R1053 VTAIL.n298 VTAIL.n297 0.155672
R1054 VTAIL.n297 VTAIL.n215 0.155672
R1055 VTAIL.n290 VTAIL.n215 0.155672
R1056 VTAIL.n290 VTAIL.n289 0.155672
R1057 VTAIL.n289 VTAIL.n219 0.155672
R1058 VTAIL.n282 VTAIL.n219 0.155672
R1059 VTAIL.n282 VTAIL.n281 0.155672
R1060 VTAIL.n281 VTAIL.n225 0.155672
R1061 VTAIL.n274 VTAIL.n225 0.155672
R1062 VTAIL.n274 VTAIL.n273 0.155672
R1063 VTAIL.n273 VTAIL.n229 0.155672
R1064 VTAIL.n266 VTAIL.n229 0.155672
R1065 VTAIL.n266 VTAIL.n265 0.155672
R1066 VTAIL.n265 VTAIL.n233 0.155672
R1067 VTAIL.n258 VTAIL.n233 0.155672
R1068 VTAIL.n258 VTAIL.n257 0.155672
R1069 VTAIL.n257 VTAIL.n237 0.155672
R1070 VTAIL.n250 VTAIL.n237 0.155672
R1071 VTAIL.n250 VTAIL.n249 0.155672
R1072 VTAIL.n249 VTAIL.n241 0.155672
R1073 VTAIL.n203 VTAIL.n109 0.155672
R1074 VTAIL.n196 VTAIL.n109 0.155672
R1075 VTAIL.n196 VTAIL.n195 0.155672
R1076 VTAIL.n195 VTAIL.n113 0.155672
R1077 VTAIL.n188 VTAIL.n113 0.155672
R1078 VTAIL.n188 VTAIL.n187 0.155672
R1079 VTAIL.n187 VTAIL.n117 0.155672
R1080 VTAIL.n180 VTAIL.n117 0.155672
R1081 VTAIL.n180 VTAIL.n179 0.155672
R1082 VTAIL.n179 VTAIL.n123 0.155672
R1083 VTAIL.n172 VTAIL.n123 0.155672
R1084 VTAIL.n172 VTAIL.n171 0.155672
R1085 VTAIL.n171 VTAIL.n127 0.155672
R1086 VTAIL.n164 VTAIL.n127 0.155672
R1087 VTAIL.n164 VTAIL.n163 0.155672
R1088 VTAIL.n163 VTAIL.n131 0.155672
R1089 VTAIL.n156 VTAIL.n131 0.155672
R1090 VTAIL.n156 VTAIL.n155 0.155672
R1091 VTAIL.n155 VTAIL.n135 0.155672
R1092 VTAIL.n148 VTAIL.n135 0.155672
R1093 VTAIL.n148 VTAIL.n147 0.155672
R1094 VTAIL.n147 VTAIL.n139 0.155672
R1095 B.n1150 B.n1149 585
R1096 B.n1151 B.n1150 585
R1097 B.n431 B.n180 585
R1098 B.n430 B.n429 585
R1099 B.n428 B.n427 585
R1100 B.n426 B.n425 585
R1101 B.n424 B.n423 585
R1102 B.n422 B.n421 585
R1103 B.n420 B.n419 585
R1104 B.n418 B.n417 585
R1105 B.n416 B.n415 585
R1106 B.n414 B.n413 585
R1107 B.n412 B.n411 585
R1108 B.n410 B.n409 585
R1109 B.n408 B.n407 585
R1110 B.n406 B.n405 585
R1111 B.n404 B.n403 585
R1112 B.n402 B.n401 585
R1113 B.n400 B.n399 585
R1114 B.n398 B.n397 585
R1115 B.n396 B.n395 585
R1116 B.n394 B.n393 585
R1117 B.n392 B.n391 585
R1118 B.n390 B.n389 585
R1119 B.n388 B.n387 585
R1120 B.n386 B.n385 585
R1121 B.n384 B.n383 585
R1122 B.n382 B.n381 585
R1123 B.n380 B.n379 585
R1124 B.n378 B.n377 585
R1125 B.n376 B.n375 585
R1126 B.n374 B.n373 585
R1127 B.n372 B.n371 585
R1128 B.n370 B.n369 585
R1129 B.n368 B.n367 585
R1130 B.n366 B.n365 585
R1131 B.n364 B.n363 585
R1132 B.n362 B.n361 585
R1133 B.n360 B.n359 585
R1134 B.n358 B.n357 585
R1135 B.n356 B.n355 585
R1136 B.n354 B.n353 585
R1137 B.n352 B.n351 585
R1138 B.n350 B.n349 585
R1139 B.n348 B.n347 585
R1140 B.n346 B.n345 585
R1141 B.n344 B.n343 585
R1142 B.n342 B.n341 585
R1143 B.n340 B.n339 585
R1144 B.n338 B.n337 585
R1145 B.n336 B.n335 585
R1146 B.n334 B.n333 585
R1147 B.n332 B.n331 585
R1148 B.n330 B.n329 585
R1149 B.n328 B.n327 585
R1150 B.n326 B.n325 585
R1151 B.n324 B.n323 585
R1152 B.n322 B.n321 585
R1153 B.n320 B.n319 585
R1154 B.n317 B.n316 585
R1155 B.n315 B.n314 585
R1156 B.n313 B.n312 585
R1157 B.n311 B.n310 585
R1158 B.n309 B.n308 585
R1159 B.n307 B.n306 585
R1160 B.n305 B.n304 585
R1161 B.n303 B.n302 585
R1162 B.n301 B.n300 585
R1163 B.n299 B.n298 585
R1164 B.n297 B.n296 585
R1165 B.n295 B.n294 585
R1166 B.n293 B.n292 585
R1167 B.n291 B.n290 585
R1168 B.n289 B.n288 585
R1169 B.n287 B.n286 585
R1170 B.n285 B.n284 585
R1171 B.n283 B.n282 585
R1172 B.n281 B.n280 585
R1173 B.n279 B.n278 585
R1174 B.n277 B.n276 585
R1175 B.n275 B.n274 585
R1176 B.n273 B.n272 585
R1177 B.n271 B.n270 585
R1178 B.n269 B.n268 585
R1179 B.n267 B.n266 585
R1180 B.n265 B.n264 585
R1181 B.n263 B.n262 585
R1182 B.n261 B.n260 585
R1183 B.n259 B.n258 585
R1184 B.n257 B.n256 585
R1185 B.n255 B.n254 585
R1186 B.n253 B.n252 585
R1187 B.n251 B.n250 585
R1188 B.n249 B.n248 585
R1189 B.n247 B.n246 585
R1190 B.n245 B.n244 585
R1191 B.n243 B.n242 585
R1192 B.n241 B.n240 585
R1193 B.n239 B.n238 585
R1194 B.n237 B.n236 585
R1195 B.n235 B.n234 585
R1196 B.n233 B.n232 585
R1197 B.n231 B.n230 585
R1198 B.n229 B.n228 585
R1199 B.n227 B.n226 585
R1200 B.n225 B.n224 585
R1201 B.n223 B.n222 585
R1202 B.n221 B.n220 585
R1203 B.n219 B.n218 585
R1204 B.n217 B.n216 585
R1205 B.n215 B.n214 585
R1206 B.n213 B.n212 585
R1207 B.n211 B.n210 585
R1208 B.n209 B.n208 585
R1209 B.n207 B.n206 585
R1210 B.n205 B.n204 585
R1211 B.n203 B.n202 585
R1212 B.n201 B.n200 585
R1213 B.n199 B.n198 585
R1214 B.n197 B.n196 585
R1215 B.n195 B.n194 585
R1216 B.n193 B.n192 585
R1217 B.n191 B.n190 585
R1218 B.n189 B.n188 585
R1219 B.n187 B.n186 585
R1220 B.n116 B.n115 585
R1221 B.n1148 B.n117 585
R1222 B.n1152 B.n117 585
R1223 B.n1147 B.n1146 585
R1224 B.n1146 B.n113 585
R1225 B.n1145 B.n112 585
R1226 B.n1158 B.n112 585
R1227 B.n1144 B.n111 585
R1228 B.n1159 B.n111 585
R1229 B.n1143 B.n110 585
R1230 B.n1160 B.n110 585
R1231 B.n1142 B.n1141 585
R1232 B.n1141 B.n106 585
R1233 B.n1140 B.n105 585
R1234 B.n1166 B.n105 585
R1235 B.n1139 B.n104 585
R1236 B.n1167 B.n104 585
R1237 B.n1138 B.n103 585
R1238 B.n1168 B.n103 585
R1239 B.n1137 B.n1136 585
R1240 B.n1136 B.n99 585
R1241 B.n1135 B.n98 585
R1242 B.n1174 B.n98 585
R1243 B.n1134 B.n97 585
R1244 B.n1175 B.n97 585
R1245 B.n1133 B.n96 585
R1246 B.n1176 B.n96 585
R1247 B.n1132 B.n1131 585
R1248 B.n1131 B.n92 585
R1249 B.n1130 B.n91 585
R1250 B.n1182 B.n91 585
R1251 B.n1129 B.n90 585
R1252 B.n1183 B.n90 585
R1253 B.n1128 B.n89 585
R1254 B.n1184 B.n89 585
R1255 B.n1127 B.n1126 585
R1256 B.n1126 B.n85 585
R1257 B.n1125 B.n84 585
R1258 B.n1190 B.n84 585
R1259 B.n1124 B.n83 585
R1260 B.n1191 B.n83 585
R1261 B.n1123 B.n82 585
R1262 B.n1192 B.n82 585
R1263 B.n1122 B.n1121 585
R1264 B.n1121 B.n78 585
R1265 B.n1120 B.n77 585
R1266 B.n1198 B.n77 585
R1267 B.n1119 B.n76 585
R1268 B.n1199 B.n76 585
R1269 B.n1118 B.n75 585
R1270 B.n1200 B.n75 585
R1271 B.n1117 B.n1116 585
R1272 B.n1116 B.n71 585
R1273 B.n1115 B.n70 585
R1274 B.n1206 B.n70 585
R1275 B.n1114 B.n69 585
R1276 B.n1207 B.n69 585
R1277 B.n1113 B.n68 585
R1278 B.n1208 B.n68 585
R1279 B.n1112 B.n1111 585
R1280 B.n1111 B.n67 585
R1281 B.n1110 B.n63 585
R1282 B.n1214 B.n63 585
R1283 B.n1109 B.n62 585
R1284 B.n1215 B.n62 585
R1285 B.n1108 B.n61 585
R1286 B.n1216 B.n61 585
R1287 B.n1107 B.n1106 585
R1288 B.n1106 B.n57 585
R1289 B.n1105 B.n56 585
R1290 B.n1222 B.n56 585
R1291 B.n1104 B.n55 585
R1292 B.n1223 B.n55 585
R1293 B.n1103 B.n54 585
R1294 B.n1224 B.n54 585
R1295 B.n1102 B.n1101 585
R1296 B.n1101 B.n50 585
R1297 B.n1100 B.n49 585
R1298 B.n1230 B.n49 585
R1299 B.n1099 B.n48 585
R1300 B.n1231 B.n48 585
R1301 B.n1098 B.n47 585
R1302 B.n1232 B.n47 585
R1303 B.n1097 B.n1096 585
R1304 B.n1096 B.n43 585
R1305 B.n1095 B.n42 585
R1306 B.n1238 B.n42 585
R1307 B.n1094 B.n41 585
R1308 B.n1239 B.n41 585
R1309 B.n1093 B.n40 585
R1310 B.n1240 B.n40 585
R1311 B.n1092 B.n1091 585
R1312 B.n1091 B.n36 585
R1313 B.n1090 B.n35 585
R1314 B.n1246 B.n35 585
R1315 B.n1089 B.n34 585
R1316 B.n1247 B.n34 585
R1317 B.n1088 B.n33 585
R1318 B.n1248 B.n33 585
R1319 B.n1087 B.n1086 585
R1320 B.n1086 B.n29 585
R1321 B.n1085 B.n28 585
R1322 B.n1254 B.n28 585
R1323 B.n1084 B.n27 585
R1324 B.n1255 B.n27 585
R1325 B.n1083 B.n26 585
R1326 B.n1256 B.n26 585
R1327 B.n1082 B.n1081 585
R1328 B.n1081 B.n22 585
R1329 B.n1080 B.n21 585
R1330 B.n1262 B.n21 585
R1331 B.n1079 B.n20 585
R1332 B.n1263 B.n20 585
R1333 B.n1078 B.n19 585
R1334 B.n1264 B.n19 585
R1335 B.n1077 B.n1076 585
R1336 B.n1076 B.n18 585
R1337 B.n1075 B.n14 585
R1338 B.n1270 B.n14 585
R1339 B.n1074 B.n13 585
R1340 B.n1271 B.n13 585
R1341 B.n1073 B.n12 585
R1342 B.n1272 B.n12 585
R1343 B.n1072 B.n1071 585
R1344 B.n1071 B.n8 585
R1345 B.n1070 B.n7 585
R1346 B.n1278 B.n7 585
R1347 B.n1069 B.n6 585
R1348 B.n1279 B.n6 585
R1349 B.n1068 B.n5 585
R1350 B.n1280 B.n5 585
R1351 B.n1067 B.n1066 585
R1352 B.n1066 B.n4 585
R1353 B.n1065 B.n432 585
R1354 B.n1065 B.n1064 585
R1355 B.n1055 B.n433 585
R1356 B.n434 B.n433 585
R1357 B.n1057 B.n1056 585
R1358 B.n1058 B.n1057 585
R1359 B.n1054 B.n439 585
R1360 B.n439 B.n438 585
R1361 B.n1053 B.n1052 585
R1362 B.n1052 B.n1051 585
R1363 B.n441 B.n440 585
R1364 B.n1044 B.n441 585
R1365 B.n1043 B.n1042 585
R1366 B.n1045 B.n1043 585
R1367 B.n1041 B.n446 585
R1368 B.n446 B.n445 585
R1369 B.n1040 B.n1039 585
R1370 B.n1039 B.n1038 585
R1371 B.n448 B.n447 585
R1372 B.n449 B.n448 585
R1373 B.n1031 B.n1030 585
R1374 B.n1032 B.n1031 585
R1375 B.n1029 B.n454 585
R1376 B.n454 B.n453 585
R1377 B.n1028 B.n1027 585
R1378 B.n1027 B.n1026 585
R1379 B.n456 B.n455 585
R1380 B.n457 B.n456 585
R1381 B.n1019 B.n1018 585
R1382 B.n1020 B.n1019 585
R1383 B.n1017 B.n462 585
R1384 B.n462 B.n461 585
R1385 B.n1016 B.n1015 585
R1386 B.n1015 B.n1014 585
R1387 B.n464 B.n463 585
R1388 B.n465 B.n464 585
R1389 B.n1007 B.n1006 585
R1390 B.n1008 B.n1007 585
R1391 B.n1005 B.n470 585
R1392 B.n470 B.n469 585
R1393 B.n1004 B.n1003 585
R1394 B.n1003 B.n1002 585
R1395 B.n472 B.n471 585
R1396 B.n473 B.n472 585
R1397 B.n995 B.n994 585
R1398 B.n996 B.n995 585
R1399 B.n993 B.n477 585
R1400 B.n481 B.n477 585
R1401 B.n992 B.n991 585
R1402 B.n991 B.n990 585
R1403 B.n479 B.n478 585
R1404 B.n480 B.n479 585
R1405 B.n983 B.n982 585
R1406 B.n984 B.n983 585
R1407 B.n981 B.n486 585
R1408 B.n486 B.n485 585
R1409 B.n980 B.n979 585
R1410 B.n979 B.n978 585
R1411 B.n488 B.n487 585
R1412 B.n489 B.n488 585
R1413 B.n971 B.n970 585
R1414 B.n972 B.n971 585
R1415 B.n969 B.n494 585
R1416 B.n494 B.n493 585
R1417 B.n968 B.n967 585
R1418 B.n967 B.n966 585
R1419 B.n496 B.n495 585
R1420 B.n959 B.n496 585
R1421 B.n958 B.n957 585
R1422 B.n960 B.n958 585
R1423 B.n956 B.n501 585
R1424 B.n501 B.n500 585
R1425 B.n955 B.n954 585
R1426 B.n954 B.n953 585
R1427 B.n503 B.n502 585
R1428 B.n504 B.n503 585
R1429 B.n946 B.n945 585
R1430 B.n947 B.n946 585
R1431 B.n944 B.n509 585
R1432 B.n509 B.n508 585
R1433 B.n943 B.n942 585
R1434 B.n942 B.n941 585
R1435 B.n511 B.n510 585
R1436 B.n512 B.n511 585
R1437 B.n934 B.n933 585
R1438 B.n935 B.n934 585
R1439 B.n932 B.n517 585
R1440 B.n517 B.n516 585
R1441 B.n931 B.n930 585
R1442 B.n930 B.n929 585
R1443 B.n519 B.n518 585
R1444 B.n520 B.n519 585
R1445 B.n922 B.n921 585
R1446 B.n923 B.n922 585
R1447 B.n920 B.n525 585
R1448 B.n525 B.n524 585
R1449 B.n919 B.n918 585
R1450 B.n918 B.n917 585
R1451 B.n527 B.n526 585
R1452 B.n528 B.n527 585
R1453 B.n910 B.n909 585
R1454 B.n911 B.n910 585
R1455 B.n908 B.n533 585
R1456 B.n533 B.n532 585
R1457 B.n907 B.n906 585
R1458 B.n906 B.n905 585
R1459 B.n535 B.n534 585
R1460 B.n536 B.n535 585
R1461 B.n898 B.n897 585
R1462 B.n899 B.n898 585
R1463 B.n896 B.n541 585
R1464 B.n541 B.n540 585
R1465 B.n895 B.n894 585
R1466 B.n894 B.n893 585
R1467 B.n543 B.n542 585
R1468 B.n544 B.n543 585
R1469 B.n886 B.n885 585
R1470 B.n887 B.n886 585
R1471 B.n884 B.n549 585
R1472 B.n549 B.n548 585
R1473 B.n883 B.n882 585
R1474 B.n882 B.n881 585
R1475 B.n551 B.n550 585
R1476 B.n552 B.n551 585
R1477 B.n874 B.n873 585
R1478 B.n875 B.n874 585
R1479 B.n555 B.n554 585
R1480 B.n624 B.n622 585
R1481 B.n625 B.n621 585
R1482 B.n625 B.n556 585
R1483 B.n628 B.n627 585
R1484 B.n629 B.n620 585
R1485 B.n631 B.n630 585
R1486 B.n633 B.n619 585
R1487 B.n636 B.n635 585
R1488 B.n637 B.n618 585
R1489 B.n639 B.n638 585
R1490 B.n641 B.n617 585
R1491 B.n644 B.n643 585
R1492 B.n645 B.n616 585
R1493 B.n647 B.n646 585
R1494 B.n649 B.n615 585
R1495 B.n652 B.n651 585
R1496 B.n653 B.n614 585
R1497 B.n655 B.n654 585
R1498 B.n657 B.n613 585
R1499 B.n660 B.n659 585
R1500 B.n661 B.n612 585
R1501 B.n663 B.n662 585
R1502 B.n665 B.n611 585
R1503 B.n668 B.n667 585
R1504 B.n669 B.n610 585
R1505 B.n671 B.n670 585
R1506 B.n673 B.n609 585
R1507 B.n676 B.n675 585
R1508 B.n677 B.n608 585
R1509 B.n679 B.n678 585
R1510 B.n681 B.n607 585
R1511 B.n684 B.n683 585
R1512 B.n685 B.n606 585
R1513 B.n687 B.n686 585
R1514 B.n689 B.n605 585
R1515 B.n692 B.n691 585
R1516 B.n693 B.n604 585
R1517 B.n695 B.n694 585
R1518 B.n697 B.n603 585
R1519 B.n700 B.n699 585
R1520 B.n701 B.n602 585
R1521 B.n703 B.n702 585
R1522 B.n705 B.n601 585
R1523 B.n708 B.n707 585
R1524 B.n709 B.n600 585
R1525 B.n711 B.n710 585
R1526 B.n713 B.n599 585
R1527 B.n716 B.n715 585
R1528 B.n717 B.n598 585
R1529 B.n719 B.n718 585
R1530 B.n721 B.n597 585
R1531 B.n724 B.n723 585
R1532 B.n725 B.n596 585
R1533 B.n727 B.n726 585
R1534 B.n729 B.n595 585
R1535 B.n732 B.n731 585
R1536 B.n733 B.n594 585
R1537 B.n738 B.n737 585
R1538 B.n740 B.n593 585
R1539 B.n743 B.n742 585
R1540 B.n744 B.n592 585
R1541 B.n746 B.n745 585
R1542 B.n748 B.n591 585
R1543 B.n751 B.n750 585
R1544 B.n752 B.n590 585
R1545 B.n754 B.n753 585
R1546 B.n756 B.n589 585
R1547 B.n759 B.n758 585
R1548 B.n760 B.n585 585
R1549 B.n762 B.n761 585
R1550 B.n764 B.n584 585
R1551 B.n767 B.n766 585
R1552 B.n768 B.n583 585
R1553 B.n770 B.n769 585
R1554 B.n772 B.n582 585
R1555 B.n775 B.n774 585
R1556 B.n776 B.n581 585
R1557 B.n778 B.n777 585
R1558 B.n780 B.n580 585
R1559 B.n783 B.n782 585
R1560 B.n784 B.n579 585
R1561 B.n786 B.n785 585
R1562 B.n788 B.n578 585
R1563 B.n791 B.n790 585
R1564 B.n792 B.n577 585
R1565 B.n794 B.n793 585
R1566 B.n796 B.n576 585
R1567 B.n799 B.n798 585
R1568 B.n800 B.n575 585
R1569 B.n802 B.n801 585
R1570 B.n804 B.n574 585
R1571 B.n807 B.n806 585
R1572 B.n808 B.n573 585
R1573 B.n810 B.n809 585
R1574 B.n812 B.n572 585
R1575 B.n815 B.n814 585
R1576 B.n816 B.n571 585
R1577 B.n818 B.n817 585
R1578 B.n820 B.n570 585
R1579 B.n823 B.n822 585
R1580 B.n824 B.n569 585
R1581 B.n826 B.n825 585
R1582 B.n828 B.n568 585
R1583 B.n831 B.n830 585
R1584 B.n832 B.n567 585
R1585 B.n834 B.n833 585
R1586 B.n836 B.n566 585
R1587 B.n839 B.n838 585
R1588 B.n840 B.n565 585
R1589 B.n842 B.n841 585
R1590 B.n844 B.n564 585
R1591 B.n847 B.n846 585
R1592 B.n848 B.n563 585
R1593 B.n850 B.n849 585
R1594 B.n852 B.n562 585
R1595 B.n855 B.n854 585
R1596 B.n856 B.n561 585
R1597 B.n858 B.n857 585
R1598 B.n860 B.n560 585
R1599 B.n863 B.n862 585
R1600 B.n864 B.n559 585
R1601 B.n866 B.n865 585
R1602 B.n868 B.n558 585
R1603 B.n871 B.n870 585
R1604 B.n872 B.n557 585
R1605 B.n877 B.n876 585
R1606 B.n876 B.n875 585
R1607 B.n878 B.n553 585
R1608 B.n553 B.n552 585
R1609 B.n880 B.n879 585
R1610 B.n881 B.n880 585
R1611 B.n547 B.n546 585
R1612 B.n548 B.n547 585
R1613 B.n889 B.n888 585
R1614 B.n888 B.n887 585
R1615 B.n890 B.n545 585
R1616 B.n545 B.n544 585
R1617 B.n892 B.n891 585
R1618 B.n893 B.n892 585
R1619 B.n539 B.n538 585
R1620 B.n540 B.n539 585
R1621 B.n901 B.n900 585
R1622 B.n900 B.n899 585
R1623 B.n902 B.n537 585
R1624 B.n537 B.n536 585
R1625 B.n904 B.n903 585
R1626 B.n905 B.n904 585
R1627 B.n531 B.n530 585
R1628 B.n532 B.n531 585
R1629 B.n913 B.n912 585
R1630 B.n912 B.n911 585
R1631 B.n914 B.n529 585
R1632 B.n529 B.n528 585
R1633 B.n916 B.n915 585
R1634 B.n917 B.n916 585
R1635 B.n523 B.n522 585
R1636 B.n524 B.n523 585
R1637 B.n925 B.n924 585
R1638 B.n924 B.n923 585
R1639 B.n926 B.n521 585
R1640 B.n521 B.n520 585
R1641 B.n928 B.n927 585
R1642 B.n929 B.n928 585
R1643 B.n515 B.n514 585
R1644 B.n516 B.n515 585
R1645 B.n937 B.n936 585
R1646 B.n936 B.n935 585
R1647 B.n938 B.n513 585
R1648 B.n513 B.n512 585
R1649 B.n940 B.n939 585
R1650 B.n941 B.n940 585
R1651 B.n507 B.n506 585
R1652 B.n508 B.n507 585
R1653 B.n949 B.n948 585
R1654 B.n948 B.n947 585
R1655 B.n950 B.n505 585
R1656 B.n505 B.n504 585
R1657 B.n952 B.n951 585
R1658 B.n953 B.n952 585
R1659 B.n499 B.n498 585
R1660 B.n500 B.n499 585
R1661 B.n962 B.n961 585
R1662 B.n961 B.n960 585
R1663 B.n963 B.n497 585
R1664 B.n959 B.n497 585
R1665 B.n965 B.n964 585
R1666 B.n966 B.n965 585
R1667 B.n492 B.n491 585
R1668 B.n493 B.n492 585
R1669 B.n974 B.n973 585
R1670 B.n973 B.n972 585
R1671 B.n975 B.n490 585
R1672 B.n490 B.n489 585
R1673 B.n977 B.n976 585
R1674 B.n978 B.n977 585
R1675 B.n484 B.n483 585
R1676 B.n485 B.n484 585
R1677 B.n986 B.n985 585
R1678 B.n985 B.n984 585
R1679 B.n987 B.n482 585
R1680 B.n482 B.n480 585
R1681 B.n989 B.n988 585
R1682 B.n990 B.n989 585
R1683 B.n476 B.n475 585
R1684 B.n481 B.n476 585
R1685 B.n998 B.n997 585
R1686 B.n997 B.n996 585
R1687 B.n999 B.n474 585
R1688 B.n474 B.n473 585
R1689 B.n1001 B.n1000 585
R1690 B.n1002 B.n1001 585
R1691 B.n468 B.n467 585
R1692 B.n469 B.n468 585
R1693 B.n1010 B.n1009 585
R1694 B.n1009 B.n1008 585
R1695 B.n1011 B.n466 585
R1696 B.n466 B.n465 585
R1697 B.n1013 B.n1012 585
R1698 B.n1014 B.n1013 585
R1699 B.n460 B.n459 585
R1700 B.n461 B.n460 585
R1701 B.n1022 B.n1021 585
R1702 B.n1021 B.n1020 585
R1703 B.n1023 B.n458 585
R1704 B.n458 B.n457 585
R1705 B.n1025 B.n1024 585
R1706 B.n1026 B.n1025 585
R1707 B.n452 B.n451 585
R1708 B.n453 B.n452 585
R1709 B.n1034 B.n1033 585
R1710 B.n1033 B.n1032 585
R1711 B.n1035 B.n450 585
R1712 B.n450 B.n449 585
R1713 B.n1037 B.n1036 585
R1714 B.n1038 B.n1037 585
R1715 B.n444 B.n443 585
R1716 B.n445 B.n444 585
R1717 B.n1047 B.n1046 585
R1718 B.n1046 B.n1045 585
R1719 B.n1048 B.n442 585
R1720 B.n1044 B.n442 585
R1721 B.n1050 B.n1049 585
R1722 B.n1051 B.n1050 585
R1723 B.n437 B.n436 585
R1724 B.n438 B.n437 585
R1725 B.n1060 B.n1059 585
R1726 B.n1059 B.n1058 585
R1727 B.n1061 B.n435 585
R1728 B.n435 B.n434 585
R1729 B.n1063 B.n1062 585
R1730 B.n1064 B.n1063 585
R1731 B.n2 B.n0 585
R1732 B.n4 B.n2 585
R1733 B.n3 B.n1 585
R1734 B.n1279 B.n3 585
R1735 B.n1277 B.n1276 585
R1736 B.n1278 B.n1277 585
R1737 B.n1275 B.n9 585
R1738 B.n9 B.n8 585
R1739 B.n1274 B.n1273 585
R1740 B.n1273 B.n1272 585
R1741 B.n11 B.n10 585
R1742 B.n1271 B.n11 585
R1743 B.n1269 B.n1268 585
R1744 B.n1270 B.n1269 585
R1745 B.n1267 B.n15 585
R1746 B.n18 B.n15 585
R1747 B.n1266 B.n1265 585
R1748 B.n1265 B.n1264 585
R1749 B.n17 B.n16 585
R1750 B.n1263 B.n17 585
R1751 B.n1261 B.n1260 585
R1752 B.n1262 B.n1261 585
R1753 B.n1259 B.n23 585
R1754 B.n23 B.n22 585
R1755 B.n1258 B.n1257 585
R1756 B.n1257 B.n1256 585
R1757 B.n25 B.n24 585
R1758 B.n1255 B.n25 585
R1759 B.n1253 B.n1252 585
R1760 B.n1254 B.n1253 585
R1761 B.n1251 B.n30 585
R1762 B.n30 B.n29 585
R1763 B.n1250 B.n1249 585
R1764 B.n1249 B.n1248 585
R1765 B.n32 B.n31 585
R1766 B.n1247 B.n32 585
R1767 B.n1245 B.n1244 585
R1768 B.n1246 B.n1245 585
R1769 B.n1243 B.n37 585
R1770 B.n37 B.n36 585
R1771 B.n1242 B.n1241 585
R1772 B.n1241 B.n1240 585
R1773 B.n39 B.n38 585
R1774 B.n1239 B.n39 585
R1775 B.n1237 B.n1236 585
R1776 B.n1238 B.n1237 585
R1777 B.n1235 B.n44 585
R1778 B.n44 B.n43 585
R1779 B.n1234 B.n1233 585
R1780 B.n1233 B.n1232 585
R1781 B.n46 B.n45 585
R1782 B.n1231 B.n46 585
R1783 B.n1229 B.n1228 585
R1784 B.n1230 B.n1229 585
R1785 B.n1227 B.n51 585
R1786 B.n51 B.n50 585
R1787 B.n1226 B.n1225 585
R1788 B.n1225 B.n1224 585
R1789 B.n53 B.n52 585
R1790 B.n1223 B.n53 585
R1791 B.n1221 B.n1220 585
R1792 B.n1222 B.n1221 585
R1793 B.n1219 B.n58 585
R1794 B.n58 B.n57 585
R1795 B.n1218 B.n1217 585
R1796 B.n1217 B.n1216 585
R1797 B.n60 B.n59 585
R1798 B.n1215 B.n60 585
R1799 B.n1213 B.n1212 585
R1800 B.n1214 B.n1213 585
R1801 B.n1211 B.n64 585
R1802 B.n67 B.n64 585
R1803 B.n1210 B.n1209 585
R1804 B.n1209 B.n1208 585
R1805 B.n66 B.n65 585
R1806 B.n1207 B.n66 585
R1807 B.n1205 B.n1204 585
R1808 B.n1206 B.n1205 585
R1809 B.n1203 B.n72 585
R1810 B.n72 B.n71 585
R1811 B.n1202 B.n1201 585
R1812 B.n1201 B.n1200 585
R1813 B.n74 B.n73 585
R1814 B.n1199 B.n74 585
R1815 B.n1197 B.n1196 585
R1816 B.n1198 B.n1197 585
R1817 B.n1195 B.n79 585
R1818 B.n79 B.n78 585
R1819 B.n1194 B.n1193 585
R1820 B.n1193 B.n1192 585
R1821 B.n81 B.n80 585
R1822 B.n1191 B.n81 585
R1823 B.n1189 B.n1188 585
R1824 B.n1190 B.n1189 585
R1825 B.n1187 B.n86 585
R1826 B.n86 B.n85 585
R1827 B.n1186 B.n1185 585
R1828 B.n1185 B.n1184 585
R1829 B.n88 B.n87 585
R1830 B.n1183 B.n88 585
R1831 B.n1181 B.n1180 585
R1832 B.n1182 B.n1181 585
R1833 B.n1179 B.n93 585
R1834 B.n93 B.n92 585
R1835 B.n1178 B.n1177 585
R1836 B.n1177 B.n1176 585
R1837 B.n95 B.n94 585
R1838 B.n1175 B.n95 585
R1839 B.n1173 B.n1172 585
R1840 B.n1174 B.n1173 585
R1841 B.n1171 B.n100 585
R1842 B.n100 B.n99 585
R1843 B.n1170 B.n1169 585
R1844 B.n1169 B.n1168 585
R1845 B.n102 B.n101 585
R1846 B.n1167 B.n102 585
R1847 B.n1165 B.n1164 585
R1848 B.n1166 B.n1165 585
R1849 B.n1163 B.n107 585
R1850 B.n107 B.n106 585
R1851 B.n1162 B.n1161 585
R1852 B.n1161 B.n1160 585
R1853 B.n109 B.n108 585
R1854 B.n1159 B.n109 585
R1855 B.n1157 B.n1156 585
R1856 B.n1158 B.n1157 585
R1857 B.n1155 B.n114 585
R1858 B.n114 B.n113 585
R1859 B.n1154 B.n1153 585
R1860 B.n1153 B.n1152 585
R1861 B.n1282 B.n1281 585
R1862 B.n1281 B.n1280 585
R1863 B.n876 B.n555 511.721
R1864 B.n1153 B.n116 511.721
R1865 B.n874 B.n557 511.721
R1866 B.n1150 B.n117 511.721
R1867 B.n586 B.t13 438.932
R1868 B.n734 B.t23 438.932
R1869 B.n183 B.t16 438.932
R1870 B.n181 B.t19 438.932
R1871 B.n587 B.t12 377.647
R1872 B.n182 B.t20 377.647
R1873 B.n735 B.t22 377.647
R1874 B.n184 B.t17 377.647
R1875 B.n586 B.t10 357.738
R1876 B.n734 B.t21 357.738
R1877 B.n183 B.t14 357.738
R1878 B.n181 B.t18 357.738
R1879 B.n1151 B.n179 256.663
R1880 B.n1151 B.n178 256.663
R1881 B.n1151 B.n177 256.663
R1882 B.n1151 B.n176 256.663
R1883 B.n1151 B.n175 256.663
R1884 B.n1151 B.n174 256.663
R1885 B.n1151 B.n173 256.663
R1886 B.n1151 B.n172 256.663
R1887 B.n1151 B.n171 256.663
R1888 B.n1151 B.n170 256.663
R1889 B.n1151 B.n169 256.663
R1890 B.n1151 B.n168 256.663
R1891 B.n1151 B.n167 256.663
R1892 B.n1151 B.n166 256.663
R1893 B.n1151 B.n165 256.663
R1894 B.n1151 B.n164 256.663
R1895 B.n1151 B.n163 256.663
R1896 B.n1151 B.n162 256.663
R1897 B.n1151 B.n161 256.663
R1898 B.n1151 B.n160 256.663
R1899 B.n1151 B.n159 256.663
R1900 B.n1151 B.n158 256.663
R1901 B.n1151 B.n157 256.663
R1902 B.n1151 B.n156 256.663
R1903 B.n1151 B.n155 256.663
R1904 B.n1151 B.n154 256.663
R1905 B.n1151 B.n153 256.663
R1906 B.n1151 B.n152 256.663
R1907 B.n1151 B.n151 256.663
R1908 B.n1151 B.n150 256.663
R1909 B.n1151 B.n149 256.663
R1910 B.n1151 B.n148 256.663
R1911 B.n1151 B.n147 256.663
R1912 B.n1151 B.n146 256.663
R1913 B.n1151 B.n145 256.663
R1914 B.n1151 B.n144 256.663
R1915 B.n1151 B.n143 256.663
R1916 B.n1151 B.n142 256.663
R1917 B.n1151 B.n141 256.663
R1918 B.n1151 B.n140 256.663
R1919 B.n1151 B.n139 256.663
R1920 B.n1151 B.n138 256.663
R1921 B.n1151 B.n137 256.663
R1922 B.n1151 B.n136 256.663
R1923 B.n1151 B.n135 256.663
R1924 B.n1151 B.n134 256.663
R1925 B.n1151 B.n133 256.663
R1926 B.n1151 B.n132 256.663
R1927 B.n1151 B.n131 256.663
R1928 B.n1151 B.n130 256.663
R1929 B.n1151 B.n129 256.663
R1930 B.n1151 B.n128 256.663
R1931 B.n1151 B.n127 256.663
R1932 B.n1151 B.n126 256.663
R1933 B.n1151 B.n125 256.663
R1934 B.n1151 B.n124 256.663
R1935 B.n1151 B.n123 256.663
R1936 B.n1151 B.n122 256.663
R1937 B.n1151 B.n121 256.663
R1938 B.n1151 B.n120 256.663
R1939 B.n1151 B.n119 256.663
R1940 B.n1151 B.n118 256.663
R1941 B.n623 B.n556 256.663
R1942 B.n626 B.n556 256.663
R1943 B.n632 B.n556 256.663
R1944 B.n634 B.n556 256.663
R1945 B.n640 B.n556 256.663
R1946 B.n642 B.n556 256.663
R1947 B.n648 B.n556 256.663
R1948 B.n650 B.n556 256.663
R1949 B.n656 B.n556 256.663
R1950 B.n658 B.n556 256.663
R1951 B.n664 B.n556 256.663
R1952 B.n666 B.n556 256.663
R1953 B.n672 B.n556 256.663
R1954 B.n674 B.n556 256.663
R1955 B.n680 B.n556 256.663
R1956 B.n682 B.n556 256.663
R1957 B.n688 B.n556 256.663
R1958 B.n690 B.n556 256.663
R1959 B.n696 B.n556 256.663
R1960 B.n698 B.n556 256.663
R1961 B.n704 B.n556 256.663
R1962 B.n706 B.n556 256.663
R1963 B.n712 B.n556 256.663
R1964 B.n714 B.n556 256.663
R1965 B.n720 B.n556 256.663
R1966 B.n722 B.n556 256.663
R1967 B.n728 B.n556 256.663
R1968 B.n730 B.n556 256.663
R1969 B.n739 B.n556 256.663
R1970 B.n741 B.n556 256.663
R1971 B.n747 B.n556 256.663
R1972 B.n749 B.n556 256.663
R1973 B.n755 B.n556 256.663
R1974 B.n757 B.n556 256.663
R1975 B.n763 B.n556 256.663
R1976 B.n765 B.n556 256.663
R1977 B.n771 B.n556 256.663
R1978 B.n773 B.n556 256.663
R1979 B.n779 B.n556 256.663
R1980 B.n781 B.n556 256.663
R1981 B.n787 B.n556 256.663
R1982 B.n789 B.n556 256.663
R1983 B.n795 B.n556 256.663
R1984 B.n797 B.n556 256.663
R1985 B.n803 B.n556 256.663
R1986 B.n805 B.n556 256.663
R1987 B.n811 B.n556 256.663
R1988 B.n813 B.n556 256.663
R1989 B.n819 B.n556 256.663
R1990 B.n821 B.n556 256.663
R1991 B.n827 B.n556 256.663
R1992 B.n829 B.n556 256.663
R1993 B.n835 B.n556 256.663
R1994 B.n837 B.n556 256.663
R1995 B.n843 B.n556 256.663
R1996 B.n845 B.n556 256.663
R1997 B.n851 B.n556 256.663
R1998 B.n853 B.n556 256.663
R1999 B.n859 B.n556 256.663
R2000 B.n861 B.n556 256.663
R2001 B.n867 B.n556 256.663
R2002 B.n869 B.n556 256.663
R2003 B.n876 B.n553 163.367
R2004 B.n880 B.n553 163.367
R2005 B.n880 B.n547 163.367
R2006 B.n888 B.n547 163.367
R2007 B.n888 B.n545 163.367
R2008 B.n892 B.n545 163.367
R2009 B.n892 B.n539 163.367
R2010 B.n900 B.n539 163.367
R2011 B.n900 B.n537 163.367
R2012 B.n904 B.n537 163.367
R2013 B.n904 B.n531 163.367
R2014 B.n912 B.n531 163.367
R2015 B.n912 B.n529 163.367
R2016 B.n916 B.n529 163.367
R2017 B.n916 B.n523 163.367
R2018 B.n924 B.n523 163.367
R2019 B.n924 B.n521 163.367
R2020 B.n928 B.n521 163.367
R2021 B.n928 B.n515 163.367
R2022 B.n936 B.n515 163.367
R2023 B.n936 B.n513 163.367
R2024 B.n940 B.n513 163.367
R2025 B.n940 B.n507 163.367
R2026 B.n948 B.n507 163.367
R2027 B.n948 B.n505 163.367
R2028 B.n952 B.n505 163.367
R2029 B.n952 B.n499 163.367
R2030 B.n961 B.n499 163.367
R2031 B.n961 B.n497 163.367
R2032 B.n965 B.n497 163.367
R2033 B.n965 B.n492 163.367
R2034 B.n973 B.n492 163.367
R2035 B.n973 B.n490 163.367
R2036 B.n977 B.n490 163.367
R2037 B.n977 B.n484 163.367
R2038 B.n985 B.n484 163.367
R2039 B.n985 B.n482 163.367
R2040 B.n989 B.n482 163.367
R2041 B.n989 B.n476 163.367
R2042 B.n997 B.n476 163.367
R2043 B.n997 B.n474 163.367
R2044 B.n1001 B.n474 163.367
R2045 B.n1001 B.n468 163.367
R2046 B.n1009 B.n468 163.367
R2047 B.n1009 B.n466 163.367
R2048 B.n1013 B.n466 163.367
R2049 B.n1013 B.n460 163.367
R2050 B.n1021 B.n460 163.367
R2051 B.n1021 B.n458 163.367
R2052 B.n1025 B.n458 163.367
R2053 B.n1025 B.n452 163.367
R2054 B.n1033 B.n452 163.367
R2055 B.n1033 B.n450 163.367
R2056 B.n1037 B.n450 163.367
R2057 B.n1037 B.n444 163.367
R2058 B.n1046 B.n444 163.367
R2059 B.n1046 B.n442 163.367
R2060 B.n1050 B.n442 163.367
R2061 B.n1050 B.n437 163.367
R2062 B.n1059 B.n437 163.367
R2063 B.n1059 B.n435 163.367
R2064 B.n1063 B.n435 163.367
R2065 B.n1063 B.n2 163.367
R2066 B.n1281 B.n2 163.367
R2067 B.n1281 B.n3 163.367
R2068 B.n1277 B.n3 163.367
R2069 B.n1277 B.n9 163.367
R2070 B.n1273 B.n9 163.367
R2071 B.n1273 B.n11 163.367
R2072 B.n1269 B.n11 163.367
R2073 B.n1269 B.n15 163.367
R2074 B.n1265 B.n15 163.367
R2075 B.n1265 B.n17 163.367
R2076 B.n1261 B.n17 163.367
R2077 B.n1261 B.n23 163.367
R2078 B.n1257 B.n23 163.367
R2079 B.n1257 B.n25 163.367
R2080 B.n1253 B.n25 163.367
R2081 B.n1253 B.n30 163.367
R2082 B.n1249 B.n30 163.367
R2083 B.n1249 B.n32 163.367
R2084 B.n1245 B.n32 163.367
R2085 B.n1245 B.n37 163.367
R2086 B.n1241 B.n37 163.367
R2087 B.n1241 B.n39 163.367
R2088 B.n1237 B.n39 163.367
R2089 B.n1237 B.n44 163.367
R2090 B.n1233 B.n44 163.367
R2091 B.n1233 B.n46 163.367
R2092 B.n1229 B.n46 163.367
R2093 B.n1229 B.n51 163.367
R2094 B.n1225 B.n51 163.367
R2095 B.n1225 B.n53 163.367
R2096 B.n1221 B.n53 163.367
R2097 B.n1221 B.n58 163.367
R2098 B.n1217 B.n58 163.367
R2099 B.n1217 B.n60 163.367
R2100 B.n1213 B.n60 163.367
R2101 B.n1213 B.n64 163.367
R2102 B.n1209 B.n64 163.367
R2103 B.n1209 B.n66 163.367
R2104 B.n1205 B.n66 163.367
R2105 B.n1205 B.n72 163.367
R2106 B.n1201 B.n72 163.367
R2107 B.n1201 B.n74 163.367
R2108 B.n1197 B.n74 163.367
R2109 B.n1197 B.n79 163.367
R2110 B.n1193 B.n79 163.367
R2111 B.n1193 B.n81 163.367
R2112 B.n1189 B.n81 163.367
R2113 B.n1189 B.n86 163.367
R2114 B.n1185 B.n86 163.367
R2115 B.n1185 B.n88 163.367
R2116 B.n1181 B.n88 163.367
R2117 B.n1181 B.n93 163.367
R2118 B.n1177 B.n93 163.367
R2119 B.n1177 B.n95 163.367
R2120 B.n1173 B.n95 163.367
R2121 B.n1173 B.n100 163.367
R2122 B.n1169 B.n100 163.367
R2123 B.n1169 B.n102 163.367
R2124 B.n1165 B.n102 163.367
R2125 B.n1165 B.n107 163.367
R2126 B.n1161 B.n107 163.367
R2127 B.n1161 B.n109 163.367
R2128 B.n1157 B.n109 163.367
R2129 B.n1157 B.n114 163.367
R2130 B.n1153 B.n114 163.367
R2131 B.n625 B.n624 163.367
R2132 B.n627 B.n625 163.367
R2133 B.n631 B.n620 163.367
R2134 B.n635 B.n633 163.367
R2135 B.n639 B.n618 163.367
R2136 B.n643 B.n641 163.367
R2137 B.n647 B.n616 163.367
R2138 B.n651 B.n649 163.367
R2139 B.n655 B.n614 163.367
R2140 B.n659 B.n657 163.367
R2141 B.n663 B.n612 163.367
R2142 B.n667 B.n665 163.367
R2143 B.n671 B.n610 163.367
R2144 B.n675 B.n673 163.367
R2145 B.n679 B.n608 163.367
R2146 B.n683 B.n681 163.367
R2147 B.n687 B.n606 163.367
R2148 B.n691 B.n689 163.367
R2149 B.n695 B.n604 163.367
R2150 B.n699 B.n697 163.367
R2151 B.n703 B.n602 163.367
R2152 B.n707 B.n705 163.367
R2153 B.n711 B.n600 163.367
R2154 B.n715 B.n713 163.367
R2155 B.n719 B.n598 163.367
R2156 B.n723 B.n721 163.367
R2157 B.n727 B.n596 163.367
R2158 B.n731 B.n729 163.367
R2159 B.n738 B.n594 163.367
R2160 B.n742 B.n740 163.367
R2161 B.n746 B.n592 163.367
R2162 B.n750 B.n748 163.367
R2163 B.n754 B.n590 163.367
R2164 B.n758 B.n756 163.367
R2165 B.n762 B.n585 163.367
R2166 B.n766 B.n764 163.367
R2167 B.n770 B.n583 163.367
R2168 B.n774 B.n772 163.367
R2169 B.n778 B.n581 163.367
R2170 B.n782 B.n780 163.367
R2171 B.n786 B.n579 163.367
R2172 B.n790 B.n788 163.367
R2173 B.n794 B.n577 163.367
R2174 B.n798 B.n796 163.367
R2175 B.n802 B.n575 163.367
R2176 B.n806 B.n804 163.367
R2177 B.n810 B.n573 163.367
R2178 B.n814 B.n812 163.367
R2179 B.n818 B.n571 163.367
R2180 B.n822 B.n820 163.367
R2181 B.n826 B.n569 163.367
R2182 B.n830 B.n828 163.367
R2183 B.n834 B.n567 163.367
R2184 B.n838 B.n836 163.367
R2185 B.n842 B.n565 163.367
R2186 B.n846 B.n844 163.367
R2187 B.n850 B.n563 163.367
R2188 B.n854 B.n852 163.367
R2189 B.n858 B.n561 163.367
R2190 B.n862 B.n860 163.367
R2191 B.n866 B.n559 163.367
R2192 B.n870 B.n868 163.367
R2193 B.n874 B.n551 163.367
R2194 B.n882 B.n551 163.367
R2195 B.n882 B.n549 163.367
R2196 B.n886 B.n549 163.367
R2197 B.n886 B.n543 163.367
R2198 B.n894 B.n543 163.367
R2199 B.n894 B.n541 163.367
R2200 B.n898 B.n541 163.367
R2201 B.n898 B.n535 163.367
R2202 B.n906 B.n535 163.367
R2203 B.n906 B.n533 163.367
R2204 B.n910 B.n533 163.367
R2205 B.n910 B.n527 163.367
R2206 B.n918 B.n527 163.367
R2207 B.n918 B.n525 163.367
R2208 B.n922 B.n525 163.367
R2209 B.n922 B.n519 163.367
R2210 B.n930 B.n519 163.367
R2211 B.n930 B.n517 163.367
R2212 B.n934 B.n517 163.367
R2213 B.n934 B.n511 163.367
R2214 B.n942 B.n511 163.367
R2215 B.n942 B.n509 163.367
R2216 B.n946 B.n509 163.367
R2217 B.n946 B.n503 163.367
R2218 B.n954 B.n503 163.367
R2219 B.n954 B.n501 163.367
R2220 B.n958 B.n501 163.367
R2221 B.n958 B.n496 163.367
R2222 B.n967 B.n496 163.367
R2223 B.n967 B.n494 163.367
R2224 B.n971 B.n494 163.367
R2225 B.n971 B.n488 163.367
R2226 B.n979 B.n488 163.367
R2227 B.n979 B.n486 163.367
R2228 B.n983 B.n486 163.367
R2229 B.n983 B.n479 163.367
R2230 B.n991 B.n479 163.367
R2231 B.n991 B.n477 163.367
R2232 B.n995 B.n477 163.367
R2233 B.n995 B.n472 163.367
R2234 B.n1003 B.n472 163.367
R2235 B.n1003 B.n470 163.367
R2236 B.n1007 B.n470 163.367
R2237 B.n1007 B.n464 163.367
R2238 B.n1015 B.n464 163.367
R2239 B.n1015 B.n462 163.367
R2240 B.n1019 B.n462 163.367
R2241 B.n1019 B.n456 163.367
R2242 B.n1027 B.n456 163.367
R2243 B.n1027 B.n454 163.367
R2244 B.n1031 B.n454 163.367
R2245 B.n1031 B.n448 163.367
R2246 B.n1039 B.n448 163.367
R2247 B.n1039 B.n446 163.367
R2248 B.n1043 B.n446 163.367
R2249 B.n1043 B.n441 163.367
R2250 B.n1052 B.n441 163.367
R2251 B.n1052 B.n439 163.367
R2252 B.n1057 B.n439 163.367
R2253 B.n1057 B.n433 163.367
R2254 B.n1065 B.n433 163.367
R2255 B.n1066 B.n1065 163.367
R2256 B.n1066 B.n5 163.367
R2257 B.n6 B.n5 163.367
R2258 B.n7 B.n6 163.367
R2259 B.n1071 B.n7 163.367
R2260 B.n1071 B.n12 163.367
R2261 B.n13 B.n12 163.367
R2262 B.n14 B.n13 163.367
R2263 B.n1076 B.n14 163.367
R2264 B.n1076 B.n19 163.367
R2265 B.n20 B.n19 163.367
R2266 B.n21 B.n20 163.367
R2267 B.n1081 B.n21 163.367
R2268 B.n1081 B.n26 163.367
R2269 B.n27 B.n26 163.367
R2270 B.n28 B.n27 163.367
R2271 B.n1086 B.n28 163.367
R2272 B.n1086 B.n33 163.367
R2273 B.n34 B.n33 163.367
R2274 B.n35 B.n34 163.367
R2275 B.n1091 B.n35 163.367
R2276 B.n1091 B.n40 163.367
R2277 B.n41 B.n40 163.367
R2278 B.n42 B.n41 163.367
R2279 B.n1096 B.n42 163.367
R2280 B.n1096 B.n47 163.367
R2281 B.n48 B.n47 163.367
R2282 B.n49 B.n48 163.367
R2283 B.n1101 B.n49 163.367
R2284 B.n1101 B.n54 163.367
R2285 B.n55 B.n54 163.367
R2286 B.n56 B.n55 163.367
R2287 B.n1106 B.n56 163.367
R2288 B.n1106 B.n61 163.367
R2289 B.n62 B.n61 163.367
R2290 B.n63 B.n62 163.367
R2291 B.n1111 B.n63 163.367
R2292 B.n1111 B.n68 163.367
R2293 B.n69 B.n68 163.367
R2294 B.n70 B.n69 163.367
R2295 B.n1116 B.n70 163.367
R2296 B.n1116 B.n75 163.367
R2297 B.n76 B.n75 163.367
R2298 B.n77 B.n76 163.367
R2299 B.n1121 B.n77 163.367
R2300 B.n1121 B.n82 163.367
R2301 B.n83 B.n82 163.367
R2302 B.n84 B.n83 163.367
R2303 B.n1126 B.n84 163.367
R2304 B.n1126 B.n89 163.367
R2305 B.n90 B.n89 163.367
R2306 B.n91 B.n90 163.367
R2307 B.n1131 B.n91 163.367
R2308 B.n1131 B.n96 163.367
R2309 B.n97 B.n96 163.367
R2310 B.n98 B.n97 163.367
R2311 B.n1136 B.n98 163.367
R2312 B.n1136 B.n103 163.367
R2313 B.n104 B.n103 163.367
R2314 B.n105 B.n104 163.367
R2315 B.n1141 B.n105 163.367
R2316 B.n1141 B.n110 163.367
R2317 B.n111 B.n110 163.367
R2318 B.n112 B.n111 163.367
R2319 B.n1146 B.n112 163.367
R2320 B.n1146 B.n117 163.367
R2321 B.n188 B.n187 163.367
R2322 B.n192 B.n191 163.367
R2323 B.n196 B.n195 163.367
R2324 B.n200 B.n199 163.367
R2325 B.n204 B.n203 163.367
R2326 B.n208 B.n207 163.367
R2327 B.n212 B.n211 163.367
R2328 B.n216 B.n215 163.367
R2329 B.n220 B.n219 163.367
R2330 B.n224 B.n223 163.367
R2331 B.n228 B.n227 163.367
R2332 B.n232 B.n231 163.367
R2333 B.n236 B.n235 163.367
R2334 B.n240 B.n239 163.367
R2335 B.n244 B.n243 163.367
R2336 B.n248 B.n247 163.367
R2337 B.n252 B.n251 163.367
R2338 B.n256 B.n255 163.367
R2339 B.n260 B.n259 163.367
R2340 B.n264 B.n263 163.367
R2341 B.n268 B.n267 163.367
R2342 B.n272 B.n271 163.367
R2343 B.n276 B.n275 163.367
R2344 B.n280 B.n279 163.367
R2345 B.n284 B.n283 163.367
R2346 B.n288 B.n287 163.367
R2347 B.n292 B.n291 163.367
R2348 B.n296 B.n295 163.367
R2349 B.n300 B.n299 163.367
R2350 B.n304 B.n303 163.367
R2351 B.n308 B.n307 163.367
R2352 B.n312 B.n311 163.367
R2353 B.n316 B.n315 163.367
R2354 B.n321 B.n320 163.367
R2355 B.n325 B.n324 163.367
R2356 B.n329 B.n328 163.367
R2357 B.n333 B.n332 163.367
R2358 B.n337 B.n336 163.367
R2359 B.n341 B.n340 163.367
R2360 B.n345 B.n344 163.367
R2361 B.n349 B.n348 163.367
R2362 B.n353 B.n352 163.367
R2363 B.n357 B.n356 163.367
R2364 B.n361 B.n360 163.367
R2365 B.n365 B.n364 163.367
R2366 B.n369 B.n368 163.367
R2367 B.n373 B.n372 163.367
R2368 B.n377 B.n376 163.367
R2369 B.n381 B.n380 163.367
R2370 B.n385 B.n384 163.367
R2371 B.n389 B.n388 163.367
R2372 B.n393 B.n392 163.367
R2373 B.n397 B.n396 163.367
R2374 B.n401 B.n400 163.367
R2375 B.n405 B.n404 163.367
R2376 B.n409 B.n408 163.367
R2377 B.n413 B.n412 163.367
R2378 B.n417 B.n416 163.367
R2379 B.n421 B.n420 163.367
R2380 B.n425 B.n424 163.367
R2381 B.n429 B.n428 163.367
R2382 B.n1150 B.n180 163.367
R2383 B.n623 B.n555 71.676
R2384 B.n627 B.n626 71.676
R2385 B.n632 B.n631 71.676
R2386 B.n635 B.n634 71.676
R2387 B.n640 B.n639 71.676
R2388 B.n643 B.n642 71.676
R2389 B.n648 B.n647 71.676
R2390 B.n651 B.n650 71.676
R2391 B.n656 B.n655 71.676
R2392 B.n659 B.n658 71.676
R2393 B.n664 B.n663 71.676
R2394 B.n667 B.n666 71.676
R2395 B.n672 B.n671 71.676
R2396 B.n675 B.n674 71.676
R2397 B.n680 B.n679 71.676
R2398 B.n683 B.n682 71.676
R2399 B.n688 B.n687 71.676
R2400 B.n691 B.n690 71.676
R2401 B.n696 B.n695 71.676
R2402 B.n699 B.n698 71.676
R2403 B.n704 B.n703 71.676
R2404 B.n707 B.n706 71.676
R2405 B.n712 B.n711 71.676
R2406 B.n715 B.n714 71.676
R2407 B.n720 B.n719 71.676
R2408 B.n723 B.n722 71.676
R2409 B.n728 B.n727 71.676
R2410 B.n731 B.n730 71.676
R2411 B.n739 B.n738 71.676
R2412 B.n742 B.n741 71.676
R2413 B.n747 B.n746 71.676
R2414 B.n750 B.n749 71.676
R2415 B.n755 B.n754 71.676
R2416 B.n758 B.n757 71.676
R2417 B.n763 B.n762 71.676
R2418 B.n766 B.n765 71.676
R2419 B.n771 B.n770 71.676
R2420 B.n774 B.n773 71.676
R2421 B.n779 B.n778 71.676
R2422 B.n782 B.n781 71.676
R2423 B.n787 B.n786 71.676
R2424 B.n790 B.n789 71.676
R2425 B.n795 B.n794 71.676
R2426 B.n798 B.n797 71.676
R2427 B.n803 B.n802 71.676
R2428 B.n806 B.n805 71.676
R2429 B.n811 B.n810 71.676
R2430 B.n814 B.n813 71.676
R2431 B.n819 B.n818 71.676
R2432 B.n822 B.n821 71.676
R2433 B.n827 B.n826 71.676
R2434 B.n830 B.n829 71.676
R2435 B.n835 B.n834 71.676
R2436 B.n838 B.n837 71.676
R2437 B.n843 B.n842 71.676
R2438 B.n846 B.n845 71.676
R2439 B.n851 B.n850 71.676
R2440 B.n854 B.n853 71.676
R2441 B.n859 B.n858 71.676
R2442 B.n862 B.n861 71.676
R2443 B.n867 B.n866 71.676
R2444 B.n870 B.n869 71.676
R2445 B.n118 B.n116 71.676
R2446 B.n188 B.n119 71.676
R2447 B.n192 B.n120 71.676
R2448 B.n196 B.n121 71.676
R2449 B.n200 B.n122 71.676
R2450 B.n204 B.n123 71.676
R2451 B.n208 B.n124 71.676
R2452 B.n212 B.n125 71.676
R2453 B.n216 B.n126 71.676
R2454 B.n220 B.n127 71.676
R2455 B.n224 B.n128 71.676
R2456 B.n228 B.n129 71.676
R2457 B.n232 B.n130 71.676
R2458 B.n236 B.n131 71.676
R2459 B.n240 B.n132 71.676
R2460 B.n244 B.n133 71.676
R2461 B.n248 B.n134 71.676
R2462 B.n252 B.n135 71.676
R2463 B.n256 B.n136 71.676
R2464 B.n260 B.n137 71.676
R2465 B.n264 B.n138 71.676
R2466 B.n268 B.n139 71.676
R2467 B.n272 B.n140 71.676
R2468 B.n276 B.n141 71.676
R2469 B.n280 B.n142 71.676
R2470 B.n284 B.n143 71.676
R2471 B.n288 B.n144 71.676
R2472 B.n292 B.n145 71.676
R2473 B.n296 B.n146 71.676
R2474 B.n300 B.n147 71.676
R2475 B.n304 B.n148 71.676
R2476 B.n308 B.n149 71.676
R2477 B.n312 B.n150 71.676
R2478 B.n316 B.n151 71.676
R2479 B.n321 B.n152 71.676
R2480 B.n325 B.n153 71.676
R2481 B.n329 B.n154 71.676
R2482 B.n333 B.n155 71.676
R2483 B.n337 B.n156 71.676
R2484 B.n341 B.n157 71.676
R2485 B.n345 B.n158 71.676
R2486 B.n349 B.n159 71.676
R2487 B.n353 B.n160 71.676
R2488 B.n357 B.n161 71.676
R2489 B.n361 B.n162 71.676
R2490 B.n365 B.n163 71.676
R2491 B.n369 B.n164 71.676
R2492 B.n373 B.n165 71.676
R2493 B.n377 B.n166 71.676
R2494 B.n381 B.n167 71.676
R2495 B.n385 B.n168 71.676
R2496 B.n389 B.n169 71.676
R2497 B.n393 B.n170 71.676
R2498 B.n397 B.n171 71.676
R2499 B.n401 B.n172 71.676
R2500 B.n405 B.n173 71.676
R2501 B.n409 B.n174 71.676
R2502 B.n413 B.n175 71.676
R2503 B.n417 B.n176 71.676
R2504 B.n421 B.n177 71.676
R2505 B.n425 B.n178 71.676
R2506 B.n429 B.n179 71.676
R2507 B.n180 B.n179 71.676
R2508 B.n428 B.n178 71.676
R2509 B.n424 B.n177 71.676
R2510 B.n420 B.n176 71.676
R2511 B.n416 B.n175 71.676
R2512 B.n412 B.n174 71.676
R2513 B.n408 B.n173 71.676
R2514 B.n404 B.n172 71.676
R2515 B.n400 B.n171 71.676
R2516 B.n396 B.n170 71.676
R2517 B.n392 B.n169 71.676
R2518 B.n388 B.n168 71.676
R2519 B.n384 B.n167 71.676
R2520 B.n380 B.n166 71.676
R2521 B.n376 B.n165 71.676
R2522 B.n372 B.n164 71.676
R2523 B.n368 B.n163 71.676
R2524 B.n364 B.n162 71.676
R2525 B.n360 B.n161 71.676
R2526 B.n356 B.n160 71.676
R2527 B.n352 B.n159 71.676
R2528 B.n348 B.n158 71.676
R2529 B.n344 B.n157 71.676
R2530 B.n340 B.n156 71.676
R2531 B.n336 B.n155 71.676
R2532 B.n332 B.n154 71.676
R2533 B.n328 B.n153 71.676
R2534 B.n324 B.n152 71.676
R2535 B.n320 B.n151 71.676
R2536 B.n315 B.n150 71.676
R2537 B.n311 B.n149 71.676
R2538 B.n307 B.n148 71.676
R2539 B.n303 B.n147 71.676
R2540 B.n299 B.n146 71.676
R2541 B.n295 B.n145 71.676
R2542 B.n291 B.n144 71.676
R2543 B.n287 B.n143 71.676
R2544 B.n283 B.n142 71.676
R2545 B.n279 B.n141 71.676
R2546 B.n275 B.n140 71.676
R2547 B.n271 B.n139 71.676
R2548 B.n267 B.n138 71.676
R2549 B.n263 B.n137 71.676
R2550 B.n259 B.n136 71.676
R2551 B.n255 B.n135 71.676
R2552 B.n251 B.n134 71.676
R2553 B.n247 B.n133 71.676
R2554 B.n243 B.n132 71.676
R2555 B.n239 B.n131 71.676
R2556 B.n235 B.n130 71.676
R2557 B.n231 B.n129 71.676
R2558 B.n227 B.n128 71.676
R2559 B.n223 B.n127 71.676
R2560 B.n219 B.n126 71.676
R2561 B.n215 B.n125 71.676
R2562 B.n211 B.n124 71.676
R2563 B.n207 B.n123 71.676
R2564 B.n203 B.n122 71.676
R2565 B.n199 B.n121 71.676
R2566 B.n195 B.n120 71.676
R2567 B.n191 B.n119 71.676
R2568 B.n187 B.n118 71.676
R2569 B.n624 B.n623 71.676
R2570 B.n626 B.n620 71.676
R2571 B.n633 B.n632 71.676
R2572 B.n634 B.n618 71.676
R2573 B.n641 B.n640 71.676
R2574 B.n642 B.n616 71.676
R2575 B.n649 B.n648 71.676
R2576 B.n650 B.n614 71.676
R2577 B.n657 B.n656 71.676
R2578 B.n658 B.n612 71.676
R2579 B.n665 B.n664 71.676
R2580 B.n666 B.n610 71.676
R2581 B.n673 B.n672 71.676
R2582 B.n674 B.n608 71.676
R2583 B.n681 B.n680 71.676
R2584 B.n682 B.n606 71.676
R2585 B.n689 B.n688 71.676
R2586 B.n690 B.n604 71.676
R2587 B.n697 B.n696 71.676
R2588 B.n698 B.n602 71.676
R2589 B.n705 B.n704 71.676
R2590 B.n706 B.n600 71.676
R2591 B.n713 B.n712 71.676
R2592 B.n714 B.n598 71.676
R2593 B.n721 B.n720 71.676
R2594 B.n722 B.n596 71.676
R2595 B.n729 B.n728 71.676
R2596 B.n730 B.n594 71.676
R2597 B.n740 B.n739 71.676
R2598 B.n741 B.n592 71.676
R2599 B.n748 B.n747 71.676
R2600 B.n749 B.n590 71.676
R2601 B.n756 B.n755 71.676
R2602 B.n757 B.n585 71.676
R2603 B.n764 B.n763 71.676
R2604 B.n765 B.n583 71.676
R2605 B.n772 B.n771 71.676
R2606 B.n773 B.n581 71.676
R2607 B.n780 B.n779 71.676
R2608 B.n781 B.n579 71.676
R2609 B.n788 B.n787 71.676
R2610 B.n789 B.n577 71.676
R2611 B.n796 B.n795 71.676
R2612 B.n797 B.n575 71.676
R2613 B.n804 B.n803 71.676
R2614 B.n805 B.n573 71.676
R2615 B.n812 B.n811 71.676
R2616 B.n813 B.n571 71.676
R2617 B.n820 B.n819 71.676
R2618 B.n821 B.n569 71.676
R2619 B.n828 B.n827 71.676
R2620 B.n829 B.n567 71.676
R2621 B.n836 B.n835 71.676
R2622 B.n837 B.n565 71.676
R2623 B.n844 B.n843 71.676
R2624 B.n845 B.n563 71.676
R2625 B.n852 B.n851 71.676
R2626 B.n853 B.n561 71.676
R2627 B.n860 B.n859 71.676
R2628 B.n861 B.n559 71.676
R2629 B.n868 B.n867 71.676
R2630 B.n869 B.n557 71.676
R2631 B.n587 B.n586 61.2853
R2632 B.n735 B.n734 61.2853
R2633 B.n184 B.n183 61.2853
R2634 B.n182 B.n181 61.2853
R2635 B.n588 B.n587 59.5399
R2636 B.n736 B.n735 59.5399
R2637 B.n185 B.n184 59.5399
R2638 B.n318 B.n182 59.5399
R2639 B.n875 B.n556 55.4465
R2640 B.n1152 B.n1151 55.4465
R2641 B.n1154 B.n115 33.2493
R2642 B.n1149 B.n1148 33.2493
R2643 B.n873 B.n872 33.2493
R2644 B.n877 B.n554 33.2493
R2645 B.n875 B.n552 32.7859
R2646 B.n881 B.n552 32.7859
R2647 B.n881 B.n548 32.7859
R2648 B.n887 B.n548 32.7859
R2649 B.n887 B.n544 32.7859
R2650 B.n893 B.n544 32.7859
R2651 B.n893 B.n540 32.7859
R2652 B.n899 B.n540 32.7859
R2653 B.n905 B.n536 32.7859
R2654 B.n905 B.n532 32.7859
R2655 B.n911 B.n532 32.7859
R2656 B.n911 B.n528 32.7859
R2657 B.n917 B.n528 32.7859
R2658 B.n917 B.n524 32.7859
R2659 B.n923 B.n524 32.7859
R2660 B.n923 B.n520 32.7859
R2661 B.n929 B.n520 32.7859
R2662 B.n929 B.n516 32.7859
R2663 B.n935 B.n516 32.7859
R2664 B.n941 B.n512 32.7859
R2665 B.n941 B.n508 32.7859
R2666 B.n947 B.n508 32.7859
R2667 B.n947 B.n504 32.7859
R2668 B.n953 B.n504 32.7859
R2669 B.n953 B.n500 32.7859
R2670 B.n960 B.n500 32.7859
R2671 B.n960 B.n959 32.7859
R2672 B.n966 B.n493 32.7859
R2673 B.n972 B.n493 32.7859
R2674 B.n972 B.n489 32.7859
R2675 B.n978 B.n489 32.7859
R2676 B.n978 B.n485 32.7859
R2677 B.n984 B.n485 32.7859
R2678 B.n984 B.n480 32.7859
R2679 B.n990 B.n480 32.7859
R2680 B.n990 B.n481 32.7859
R2681 B.n996 B.n473 32.7859
R2682 B.n1002 B.n473 32.7859
R2683 B.n1002 B.n469 32.7859
R2684 B.n1008 B.n469 32.7859
R2685 B.n1008 B.n465 32.7859
R2686 B.n1014 B.n465 32.7859
R2687 B.n1014 B.n461 32.7859
R2688 B.n1020 B.n461 32.7859
R2689 B.n1026 B.n457 32.7859
R2690 B.n1026 B.n453 32.7859
R2691 B.n1032 B.n453 32.7859
R2692 B.n1032 B.n449 32.7859
R2693 B.n1038 B.n449 32.7859
R2694 B.n1038 B.n445 32.7859
R2695 B.n1045 B.n445 32.7859
R2696 B.n1045 B.n1044 32.7859
R2697 B.n1051 B.n438 32.7859
R2698 B.n1058 B.n438 32.7859
R2699 B.n1058 B.n434 32.7859
R2700 B.n1064 B.n434 32.7859
R2701 B.n1064 B.n4 32.7859
R2702 B.n1280 B.n4 32.7859
R2703 B.n1280 B.n1279 32.7859
R2704 B.n1279 B.n1278 32.7859
R2705 B.n1278 B.n8 32.7859
R2706 B.n1272 B.n8 32.7859
R2707 B.n1272 B.n1271 32.7859
R2708 B.n1271 B.n1270 32.7859
R2709 B.n1264 B.n18 32.7859
R2710 B.n1264 B.n1263 32.7859
R2711 B.n1263 B.n1262 32.7859
R2712 B.n1262 B.n22 32.7859
R2713 B.n1256 B.n22 32.7859
R2714 B.n1256 B.n1255 32.7859
R2715 B.n1255 B.n1254 32.7859
R2716 B.n1254 B.n29 32.7859
R2717 B.n1248 B.n1247 32.7859
R2718 B.n1247 B.n1246 32.7859
R2719 B.n1246 B.n36 32.7859
R2720 B.n1240 B.n36 32.7859
R2721 B.n1240 B.n1239 32.7859
R2722 B.n1239 B.n1238 32.7859
R2723 B.n1238 B.n43 32.7859
R2724 B.n1232 B.n43 32.7859
R2725 B.n1231 B.n1230 32.7859
R2726 B.n1230 B.n50 32.7859
R2727 B.n1224 B.n50 32.7859
R2728 B.n1224 B.n1223 32.7859
R2729 B.n1223 B.n1222 32.7859
R2730 B.n1222 B.n57 32.7859
R2731 B.n1216 B.n57 32.7859
R2732 B.n1216 B.n1215 32.7859
R2733 B.n1215 B.n1214 32.7859
R2734 B.n1208 B.n67 32.7859
R2735 B.n1208 B.n1207 32.7859
R2736 B.n1207 B.n1206 32.7859
R2737 B.n1206 B.n71 32.7859
R2738 B.n1200 B.n71 32.7859
R2739 B.n1200 B.n1199 32.7859
R2740 B.n1199 B.n1198 32.7859
R2741 B.n1198 B.n78 32.7859
R2742 B.n1192 B.n1191 32.7859
R2743 B.n1191 B.n1190 32.7859
R2744 B.n1190 B.n85 32.7859
R2745 B.n1184 B.n85 32.7859
R2746 B.n1184 B.n1183 32.7859
R2747 B.n1183 B.n1182 32.7859
R2748 B.n1182 B.n92 32.7859
R2749 B.n1176 B.n92 32.7859
R2750 B.n1176 B.n1175 32.7859
R2751 B.n1175 B.n1174 32.7859
R2752 B.n1174 B.n99 32.7859
R2753 B.n1168 B.n1167 32.7859
R2754 B.n1167 B.n1166 32.7859
R2755 B.n1166 B.n106 32.7859
R2756 B.n1160 B.n106 32.7859
R2757 B.n1160 B.n1159 32.7859
R2758 B.n1159 B.n1158 32.7859
R2759 B.n1158 B.n113 32.7859
R2760 B.n1152 B.n113 32.7859
R2761 B.t11 B.n536 30.3753
R2762 B.t15 B.n99 30.3753
R2763 B.n959 B.t2 28.4467
R2764 B.n67 B.t1 28.4467
R2765 B.n996 B.t8 27.4824
R2766 B.n1232 B.t6 27.4824
R2767 B.n1044 B.t5 24.5896
R2768 B.n18 B.t0 24.5896
R2769 B.n935 B.t9 18.8039
R2770 B.n1192 B.t7 18.8039
R2771 B B.n1282 18.0485
R2772 B.t4 B.n457 17.8396
R2773 B.t3 B.n29 17.8396
R2774 B.n1020 B.t4 14.9468
R2775 B.n1248 B.t3 14.9468
R2776 B.t9 B.n512 13.9825
R2777 B.t7 B.n78 13.9825
R2778 B.n186 B.n115 10.6151
R2779 B.n189 B.n186 10.6151
R2780 B.n190 B.n189 10.6151
R2781 B.n193 B.n190 10.6151
R2782 B.n194 B.n193 10.6151
R2783 B.n197 B.n194 10.6151
R2784 B.n198 B.n197 10.6151
R2785 B.n201 B.n198 10.6151
R2786 B.n202 B.n201 10.6151
R2787 B.n205 B.n202 10.6151
R2788 B.n206 B.n205 10.6151
R2789 B.n209 B.n206 10.6151
R2790 B.n210 B.n209 10.6151
R2791 B.n213 B.n210 10.6151
R2792 B.n214 B.n213 10.6151
R2793 B.n217 B.n214 10.6151
R2794 B.n218 B.n217 10.6151
R2795 B.n221 B.n218 10.6151
R2796 B.n222 B.n221 10.6151
R2797 B.n225 B.n222 10.6151
R2798 B.n226 B.n225 10.6151
R2799 B.n229 B.n226 10.6151
R2800 B.n230 B.n229 10.6151
R2801 B.n233 B.n230 10.6151
R2802 B.n234 B.n233 10.6151
R2803 B.n237 B.n234 10.6151
R2804 B.n238 B.n237 10.6151
R2805 B.n241 B.n238 10.6151
R2806 B.n242 B.n241 10.6151
R2807 B.n245 B.n242 10.6151
R2808 B.n246 B.n245 10.6151
R2809 B.n249 B.n246 10.6151
R2810 B.n250 B.n249 10.6151
R2811 B.n253 B.n250 10.6151
R2812 B.n254 B.n253 10.6151
R2813 B.n257 B.n254 10.6151
R2814 B.n258 B.n257 10.6151
R2815 B.n261 B.n258 10.6151
R2816 B.n262 B.n261 10.6151
R2817 B.n265 B.n262 10.6151
R2818 B.n266 B.n265 10.6151
R2819 B.n269 B.n266 10.6151
R2820 B.n270 B.n269 10.6151
R2821 B.n273 B.n270 10.6151
R2822 B.n274 B.n273 10.6151
R2823 B.n277 B.n274 10.6151
R2824 B.n278 B.n277 10.6151
R2825 B.n281 B.n278 10.6151
R2826 B.n282 B.n281 10.6151
R2827 B.n285 B.n282 10.6151
R2828 B.n286 B.n285 10.6151
R2829 B.n289 B.n286 10.6151
R2830 B.n290 B.n289 10.6151
R2831 B.n293 B.n290 10.6151
R2832 B.n294 B.n293 10.6151
R2833 B.n297 B.n294 10.6151
R2834 B.n298 B.n297 10.6151
R2835 B.n302 B.n301 10.6151
R2836 B.n305 B.n302 10.6151
R2837 B.n306 B.n305 10.6151
R2838 B.n309 B.n306 10.6151
R2839 B.n310 B.n309 10.6151
R2840 B.n313 B.n310 10.6151
R2841 B.n314 B.n313 10.6151
R2842 B.n317 B.n314 10.6151
R2843 B.n322 B.n319 10.6151
R2844 B.n323 B.n322 10.6151
R2845 B.n326 B.n323 10.6151
R2846 B.n327 B.n326 10.6151
R2847 B.n330 B.n327 10.6151
R2848 B.n331 B.n330 10.6151
R2849 B.n334 B.n331 10.6151
R2850 B.n335 B.n334 10.6151
R2851 B.n338 B.n335 10.6151
R2852 B.n339 B.n338 10.6151
R2853 B.n342 B.n339 10.6151
R2854 B.n343 B.n342 10.6151
R2855 B.n346 B.n343 10.6151
R2856 B.n347 B.n346 10.6151
R2857 B.n350 B.n347 10.6151
R2858 B.n351 B.n350 10.6151
R2859 B.n354 B.n351 10.6151
R2860 B.n355 B.n354 10.6151
R2861 B.n358 B.n355 10.6151
R2862 B.n359 B.n358 10.6151
R2863 B.n362 B.n359 10.6151
R2864 B.n363 B.n362 10.6151
R2865 B.n366 B.n363 10.6151
R2866 B.n367 B.n366 10.6151
R2867 B.n370 B.n367 10.6151
R2868 B.n371 B.n370 10.6151
R2869 B.n374 B.n371 10.6151
R2870 B.n375 B.n374 10.6151
R2871 B.n378 B.n375 10.6151
R2872 B.n379 B.n378 10.6151
R2873 B.n382 B.n379 10.6151
R2874 B.n383 B.n382 10.6151
R2875 B.n386 B.n383 10.6151
R2876 B.n387 B.n386 10.6151
R2877 B.n390 B.n387 10.6151
R2878 B.n391 B.n390 10.6151
R2879 B.n394 B.n391 10.6151
R2880 B.n395 B.n394 10.6151
R2881 B.n398 B.n395 10.6151
R2882 B.n399 B.n398 10.6151
R2883 B.n402 B.n399 10.6151
R2884 B.n403 B.n402 10.6151
R2885 B.n406 B.n403 10.6151
R2886 B.n407 B.n406 10.6151
R2887 B.n410 B.n407 10.6151
R2888 B.n411 B.n410 10.6151
R2889 B.n414 B.n411 10.6151
R2890 B.n415 B.n414 10.6151
R2891 B.n418 B.n415 10.6151
R2892 B.n419 B.n418 10.6151
R2893 B.n422 B.n419 10.6151
R2894 B.n423 B.n422 10.6151
R2895 B.n426 B.n423 10.6151
R2896 B.n427 B.n426 10.6151
R2897 B.n430 B.n427 10.6151
R2898 B.n431 B.n430 10.6151
R2899 B.n1149 B.n431 10.6151
R2900 B.n873 B.n550 10.6151
R2901 B.n883 B.n550 10.6151
R2902 B.n884 B.n883 10.6151
R2903 B.n885 B.n884 10.6151
R2904 B.n885 B.n542 10.6151
R2905 B.n895 B.n542 10.6151
R2906 B.n896 B.n895 10.6151
R2907 B.n897 B.n896 10.6151
R2908 B.n897 B.n534 10.6151
R2909 B.n907 B.n534 10.6151
R2910 B.n908 B.n907 10.6151
R2911 B.n909 B.n908 10.6151
R2912 B.n909 B.n526 10.6151
R2913 B.n919 B.n526 10.6151
R2914 B.n920 B.n919 10.6151
R2915 B.n921 B.n920 10.6151
R2916 B.n921 B.n518 10.6151
R2917 B.n931 B.n518 10.6151
R2918 B.n932 B.n931 10.6151
R2919 B.n933 B.n932 10.6151
R2920 B.n933 B.n510 10.6151
R2921 B.n943 B.n510 10.6151
R2922 B.n944 B.n943 10.6151
R2923 B.n945 B.n944 10.6151
R2924 B.n945 B.n502 10.6151
R2925 B.n955 B.n502 10.6151
R2926 B.n956 B.n955 10.6151
R2927 B.n957 B.n956 10.6151
R2928 B.n957 B.n495 10.6151
R2929 B.n968 B.n495 10.6151
R2930 B.n969 B.n968 10.6151
R2931 B.n970 B.n969 10.6151
R2932 B.n970 B.n487 10.6151
R2933 B.n980 B.n487 10.6151
R2934 B.n981 B.n980 10.6151
R2935 B.n982 B.n981 10.6151
R2936 B.n982 B.n478 10.6151
R2937 B.n992 B.n478 10.6151
R2938 B.n993 B.n992 10.6151
R2939 B.n994 B.n993 10.6151
R2940 B.n994 B.n471 10.6151
R2941 B.n1004 B.n471 10.6151
R2942 B.n1005 B.n1004 10.6151
R2943 B.n1006 B.n1005 10.6151
R2944 B.n1006 B.n463 10.6151
R2945 B.n1016 B.n463 10.6151
R2946 B.n1017 B.n1016 10.6151
R2947 B.n1018 B.n1017 10.6151
R2948 B.n1018 B.n455 10.6151
R2949 B.n1028 B.n455 10.6151
R2950 B.n1029 B.n1028 10.6151
R2951 B.n1030 B.n1029 10.6151
R2952 B.n1030 B.n447 10.6151
R2953 B.n1040 B.n447 10.6151
R2954 B.n1041 B.n1040 10.6151
R2955 B.n1042 B.n1041 10.6151
R2956 B.n1042 B.n440 10.6151
R2957 B.n1053 B.n440 10.6151
R2958 B.n1054 B.n1053 10.6151
R2959 B.n1056 B.n1054 10.6151
R2960 B.n1056 B.n1055 10.6151
R2961 B.n1055 B.n432 10.6151
R2962 B.n1067 B.n432 10.6151
R2963 B.n1068 B.n1067 10.6151
R2964 B.n1069 B.n1068 10.6151
R2965 B.n1070 B.n1069 10.6151
R2966 B.n1072 B.n1070 10.6151
R2967 B.n1073 B.n1072 10.6151
R2968 B.n1074 B.n1073 10.6151
R2969 B.n1075 B.n1074 10.6151
R2970 B.n1077 B.n1075 10.6151
R2971 B.n1078 B.n1077 10.6151
R2972 B.n1079 B.n1078 10.6151
R2973 B.n1080 B.n1079 10.6151
R2974 B.n1082 B.n1080 10.6151
R2975 B.n1083 B.n1082 10.6151
R2976 B.n1084 B.n1083 10.6151
R2977 B.n1085 B.n1084 10.6151
R2978 B.n1087 B.n1085 10.6151
R2979 B.n1088 B.n1087 10.6151
R2980 B.n1089 B.n1088 10.6151
R2981 B.n1090 B.n1089 10.6151
R2982 B.n1092 B.n1090 10.6151
R2983 B.n1093 B.n1092 10.6151
R2984 B.n1094 B.n1093 10.6151
R2985 B.n1095 B.n1094 10.6151
R2986 B.n1097 B.n1095 10.6151
R2987 B.n1098 B.n1097 10.6151
R2988 B.n1099 B.n1098 10.6151
R2989 B.n1100 B.n1099 10.6151
R2990 B.n1102 B.n1100 10.6151
R2991 B.n1103 B.n1102 10.6151
R2992 B.n1104 B.n1103 10.6151
R2993 B.n1105 B.n1104 10.6151
R2994 B.n1107 B.n1105 10.6151
R2995 B.n1108 B.n1107 10.6151
R2996 B.n1109 B.n1108 10.6151
R2997 B.n1110 B.n1109 10.6151
R2998 B.n1112 B.n1110 10.6151
R2999 B.n1113 B.n1112 10.6151
R3000 B.n1114 B.n1113 10.6151
R3001 B.n1115 B.n1114 10.6151
R3002 B.n1117 B.n1115 10.6151
R3003 B.n1118 B.n1117 10.6151
R3004 B.n1119 B.n1118 10.6151
R3005 B.n1120 B.n1119 10.6151
R3006 B.n1122 B.n1120 10.6151
R3007 B.n1123 B.n1122 10.6151
R3008 B.n1124 B.n1123 10.6151
R3009 B.n1125 B.n1124 10.6151
R3010 B.n1127 B.n1125 10.6151
R3011 B.n1128 B.n1127 10.6151
R3012 B.n1129 B.n1128 10.6151
R3013 B.n1130 B.n1129 10.6151
R3014 B.n1132 B.n1130 10.6151
R3015 B.n1133 B.n1132 10.6151
R3016 B.n1134 B.n1133 10.6151
R3017 B.n1135 B.n1134 10.6151
R3018 B.n1137 B.n1135 10.6151
R3019 B.n1138 B.n1137 10.6151
R3020 B.n1139 B.n1138 10.6151
R3021 B.n1140 B.n1139 10.6151
R3022 B.n1142 B.n1140 10.6151
R3023 B.n1143 B.n1142 10.6151
R3024 B.n1144 B.n1143 10.6151
R3025 B.n1145 B.n1144 10.6151
R3026 B.n1147 B.n1145 10.6151
R3027 B.n1148 B.n1147 10.6151
R3028 B.n622 B.n554 10.6151
R3029 B.n622 B.n621 10.6151
R3030 B.n628 B.n621 10.6151
R3031 B.n629 B.n628 10.6151
R3032 B.n630 B.n629 10.6151
R3033 B.n630 B.n619 10.6151
R3034 B.n636 B.n619 10.6151
R3035 B.n637 B.n636 10.6151
R3036 B.n638 B.n637 10.6151
R3037 B.n638 B.n617 10.6151
R3038 B.n644 B.n617 10.6151
R3039 B.n645 B.n644 10.6151
R3040 B.n646 B.n645 10.6151
R3041 B.n646 B.n615 10.6151
R3042 B.n652 B.n615 10.6151
R3043 B.n653 B.n652 10.6151
R3044 B.n654 B.n653 10.6151
R3045 B.n654 B.n613 10.6151
R3046 B.n660 B.n613 10.6151
R3047 B.n661 B.n660 10.6151
R3048 B.n662 B.n661 10.6151
R3049 B.n662 B.n611 10.6151
R3050 B.n668 B.n611 10.6151
R3051 B.n669 B.n668 10.6151
R3052 B.n670 B.n669 10.6151
R3053 B.n670 B.n609 10.6151
R3054 B.n676 B.n609 10.6151
R3055 B.n677 B.n676 10.6151
R3056 B.n678 B.n677 10.6151
R3057 B.n678 B.n607 10.6151
R3058 B.n684 B.n607 10.6151
R3059 B.n685 B.n684 10.6151
R3060 B.n686 B.n685 10.6151
R3061 B.n686 B.n605 10.6151
R3062 B.n692 B.n605 10.6151
R3063 B.n693 B.n692 10.6151
R3064 B.n694 B.n693 10.6151
R3065 B.n694 B.n603 10.6151
R3066 B.n700 B.n603 10.6151
R3067 B.n701 B.n700 10.6151
R3068 B.n702 B.n701 10.6151
R3069 B.n702 B.n601 10.6151
R3070 B.n708 B.n601 10.6151
R3071 B.n709 B.n708 10.6151
R3072 B.n710 B.n709 10.6151
R3073 B.n710 B.n599 10.6151
R3074 B.n716 B.n599 10.6151
R3075 B.n717 B.n716 10.6151
R3076 B.n718 B.n717 10.6151
R3077 B.n718 B.n597 10.6151
R3078 B.n724 B.n597 10.6151
R3079 B.n725 B.n724 10.6151
R3080 B.n726 B.n725 10.6151
R3081 B.n726 B.n595 10.6151
R3082 B.n732 B.n595 10.6151
R3083 B.n733 B.n732 10.6151
R3084 B.n737 B.n733 10.6151
R3085 B.n743 B.n593 10.6151
R3086 B.n744 B.n743 10.6151
R3087 B.n745 B.n744 10.6151
R3088 B.n745 B.n591 10.6151
R3089 B.n751 B.n591 10.6151
R3090 B.n752 B.n751 10.6151
R3091 B.n753 B.n752 10.6151
R3092 B.n753 B.n589 10.6151
R3093 B.n760 B.n759 10.6151
R3094 B.n761 B.n760 10.6151
R3095 B.n761 B.n584 10.6151
R3096 B.n767 B.n584 10.6151
R3097 B.n768 B.n767 10.6151
R3098 B.n769 B.n768 10.6151
R3099 B.n769 B.n582 10.6151
R3100 B.n775 B.n582 10.6151
R3101 B.n776 B.n775 10.6151
R3102 B.n777 B.n776 10.6151
R3103 B.n777 B.n580 10.6151
R3104 B.n783 B.n580 10.6151
R3105 B.n784 B.n783 10.6151
R3106 B.n785 B.n784 10.6151
R3107 B.n785 B.n578 10.6151
R3108 B.n791 B.n578 10.6151
R3109 B.n792 B.n791 10.6151
R3110 B.n793 B.n792 10.6151
R3111 B.n793 B.n576 10.6151
R3112 B.n799 B.n576 10.6151
R3113 B.n800 B.n799 10.6151
R3114 B.n801 B.n800 10.6151
R3115 B.n801 B.n574 10.6151
R3116 B.n807 B.n574 10.6151
R3117 B.n808 B.n807 10.6151
R3118 B.n809 B.n808 10.6151
R3119 B.n809 B.n572 10.6151
R3120 B.n815 B.n572 10.6151
R3121 B.n816 B.n815 10.6151
R3122 B.n817 B.n816 10.6151
R3123 B.n817 B.n570 10.6151
R3124 B.n823 B.n570 10.6151
R3125 B.n824 B.n823 10.6151
R3126 B.n825 B.n824 10.6151
R3127 B.n825 B.n568 10.6151
R3128 B.n831 B.n568 10.6151
R3129 B.n832 B.n831 10.6151
R3130 B.n833 B.n832 10.6151
R3131 B.n833 B.n566 10.6151
R3132 B.n839 B.n566 10.6151
R3133 B.n840 B.n839 10.6151
R3134 B.n841 B.n840 10.6151
R3135 B.n841 B.n564 10.6151
R3136 B.n847 B.n564 10.6151
R3137 B.n848 B.n847 10.6151
R3138 B.n849 B.n848 10.6151
R3139 B.n849 B.n562 10.6151
R3140 B.n855 B.n562 10.6151
R3141 B.n856 B.n855 10.6151
R3142 B.n857 B.n856 10.6151
R3143 B.n857 B.n560 10.6151
R3144 B.n863 B.n560 10.6151
R3145 B.n864 B.n863 10.6151
R3146 B.n865 B.n864 10.6151
R3147 B.n865 B.n558 10.6151
R3148 B.n871 B.n558 10.6151
R3149 B.n872 B.n871 10.6151
R3150 B.n878 B.n877 10.6151
R3151 B.n879 B.n878 10.6151
R3152 B.n879 B.n546 10.6151
R3153 B.n889 B.n546 10.6151
R3154 B.n890 B.n889 10.6151
R3155 B.n891 B.n890 10.6151
R3156 B.n891 B.n538 10.6151
R3157 B.n901 B.n538 10.6151
R3158 B.n902 B.n901 10.6151
R3159 B.n903 B.n902 10.6151
R3160 B.n903 B.n530 10.6151
R3161 B.n913 B.n530 10.6151
R3162 B.n914 B.n913 10.6151
R3163 B.n915 B.n914 10.6151
R3164 B.n915 B.n522 10.6151
R3165 B.n925 B.n522 10.6151
R3166 B.n926 B.n925 10.6151
R3167 B.n927 B.n926 10.6151
R3168 B.n927 B.n514 10.6151
R3169 B.n937 B.n514 10.6151
R3170 B.n938 B.n937 10.6151
R3171 B.n939 B.n938 10.6151
R3172 B.n939 B.n506 10.6151
R3173 B.n949 B.n506 10.6151
R3174 B.n950 B.n949 10.6151
R3175 B.n951 B.n950 10.6151
R3176 B.n951 B.n498 10.6151
R3177 B.n962 B.n498 10.6151
R3178 B.n963 B.n962 10.6151
R3179 B.n964 B.n963 10.6151
R3180 B.n964 B.n491 10.6151
R3181 B.n974 B.n491 10.6151
R3182 B.n975 B.n974 10.6151
R3183 B.n976 B.n975 10.6151
R3184 B.n976 B.n483 10.6151
R3185 B.n986 B.n483 10.6151
R3186 B.n987 B.n986 10.6151
R3187 B.n988 B.n987 10.6151
R3188 B.n988 B.n475 10.6151
R3189 B.n998 B.n475 10.6151
R3190 B.n999 B.n998 10.6151
R3191 B.n1000 B.n999 10.6151
R3192 B.n1000 B.n467 10.6151
R3193 B.n1010 B.n467 10.6151
R3194 B.n1011 B.n1010 10.6151
R3195 B.n1012 B.n1011 10.6151
R3196 B.n1012 B.n459 10.6151
R3197 B.n1022 B.n459 10.6151
R3198 B.n1023 B.n1022 10.6151
R3199 B.n1024 B.n1023 10.6151
R3200 B.n1024 B.n451 10.6151
R3201 B.n1034 B.n451 10.6151
R3202 B.n1035 B.n1034 10.6151
R3203 B.n1036 B.n1035 10.6151
R3204 B.n1036 B.n443 10.6151
R3205 B.n1047 B.n443 10.6151
R3206 B.n1048 B.n1047 10.6151
R3207 B.n1049 B.n1048 10.6151
R3208 B.n1049 B.n436 10.6151
R3209 B.n1060 B.n436 10.6151
R3210 B.n1061 B.n1060 10.6151
R3211 B.n1062 B.n1061 10.6151
R3212 B.n1062 B.n0 10.6151
R3213 B.n1276 B.n1 10.6151
R3214 B.n1276 B.n1275 10.6151
R3215 B.n1275 B.n1274 10.6151
R3216 B.n1274 B.n10 10.6151
R3217 B.n1268 B.n10 10.6151
R3218 B.n1268 B.n1267 10.6151
R3219 B.n1267 B.n1266 10.6151
R3220 B.n1266 B.n16 10.6151
R3221 B.n1260 B.n16 10.6151
R3222 B.n1260 B.n1259 10.6151
R3223 B.n1259 B.n1258 10.6151
R3224 B.n1258 B.n24 10.6151
R3225 B.n1252 B.n24 10.6151
R3226 B.n1252 B.n1251 10.6151
R3227 B.n1251 B.n1250 10.6151
R3228 B.n1250 B.n31 10.6151
R3229 B.n1244 B.n31 10.6151
R3230 B.n1244 B.n1243 10.6151
R3231 B.n1243 B.n1242 10.6151
R3232 B.n1242 B.n38 10.6151
R3233 B.n1236 B.n38 10.6151
R3234 B.n1236 B.n1235 10.6151
R3235 B.n1235 B.n1234 10.6151
R3236 B.n1234 B.n45 10.6151
R3237 B.n1228 B.n45 10.6151
R3238 B.n1228 B.n1227 10.6151
R3239 B.n1227 B.n1226 10.6151
R3240 B.n1226 B.n52 10.6151
R3241 B.n1220 B.n52 10.6151
R3242 B.n1220 B.n1219 10.6151
R3243 B.n1219 B.n1218 10.6151
R3244 B.n1218 B.n59 10.6151
R3245 B.n1212 B.n59 10.6151
R3246 B.n1212 B.n1211 10.6151
R3247 B.n1211 B.n1210 10.6151
R3248 B.n1210 B.n65 10.6151
R3249 B.n1204 B.n65 10.6151
R3250 B.n1204 B.n1203 10.6151
R3251 B.n1203 B.n1202 10.6151
R3252 B.n1202 B.n73 10.6151
R3253 B.n1196 B.n73 10.6151
R3254 B.n1196 B.n1195 10.6151
R3255 B.n1195 B.n1194 10.6151
R3256 B.n1194 B.n80 10.6151
R3257 B.n1188 B.n80 10.6151
R3258 B.n1188 B.n1187 10.6151
R3259 B.n1187 B.n1186 10.6151
R3260 B.n1186 B.n87 10.6151
R3261 B.n1180 B.n87 10.6151
R3262 B.n1180 B.n1179 10.6151
R3263 B.n1179 B.n1178 10.6151
R3264 B.n1178 B.n94 10.6151
R3265 B.n1172 B.n94 10.6151
R3266 B.n1172 B.n1171 10.6151
R3267 B.n1171 B.n1170 10.6151
R3268 B.n1170 B.n101 10.6151
R3269 B.n1164 B.n101 10.6151
R3270 B.n1164 B.n1163 10.6151
R3271 B.n1163 B.n1162 10.6151
R3272 B.n1162 B.n108 10.6151
R3273 B.n1156 B.n108 10.6151
R3274 B.n1156 B.n1155 10.6151
R3275 B.n1155 B.n1154 10.6151
R3276 B.n1051 B.t5 8.19686
R3277 B.n1270 B.t0 8.19686
R3278 B.n301 B.n185 6.5566
R3279 B.n318 B.n317 6.5566
R3280 B.n736 B.n593 6.5566
R3281 B.n589 B.n588 6.5566
R3282 B.n481 B.t8 5.30403
R3283 B.t6 B.n1231 5.30403
R3284 B.n966 B.t2 4.33975
R3285 B.n1214 B.t1 4.33975
R3286 B.n298 B.n185 4.05904
R3287 B.n319 B.n318 4.05904
R3288 B.n737 B.n736 4.05904
R3289 B.n759 B.n588 4.05904
R3290 B.n1282 B.n0 2.81026
R3291 B.n1282 B.n1 2.81026
R3292 B.n899 B.t11 2.41119
R3293 B.n1168 B.t15 2.41119
R3294 VN.n11 VN.t2 182.843
R3295 VN.n56 VN.t8 182.843
R3296 VN.n85 VN.n44 161.3
R3297 VN.n84 VN.n83 161.3
R3298 VN.n82 VN.n45 161.3
R3299 VN.n81 VN.n80 161.3
R3300 VN.n79 VN.n46 161.3
R3301 VN.n78 VN.n77 161.3
R3302 VN.n76 VN.n47 161.3
R3303 VN.n75 VN.n74 161.3
R3304 VN.n73 VN.n48 161.3
R3305 VN.n72 VN.n71 161.3
R3306 VN.n70 VN.n50 161.3
R3307 VN.n69 VN.n68 161.3
R3308 VN.n67 VN.n51 161.3
R3309 VN.n65 VN.n64 161.3
R3310 VN.n63 VN.n52 161.3
R3311 VN.n62 VN.n61 161.3
R3312 VN.n60 VN.n53 161.3
R3313 VN.n59 VN.n58 161.3
R3314 VN.n57 VN.n54 161.3
R3315 VN.n41 VN.n0 161.3
R3316 VN.n40 VN.n39 161.3
R3317 VN.n38 VN.n1 161.3
R3318 VN.n37 VN.n36 161.3
R3319 VN.n35 VN.n2 161.3
R3320 VN.n34 VN.n33 161.3
R3321 VN.n32 VN.n3 161.3
R3322 VN.n31 VN.n30 161.3
R3323 VN.n28 VN.n4 161.3
R3324 VN.n27 VN.n26 161.3
R3325 VN.n25 VN.n5 161.3
R3326 VN.n24 VN.n23 161.3
R3327 VN.n22 VN.n6 161.3
R3328 VN.n20 VN.n19 161.3
R3329 VN.n18 VN.n7 161.3
R3330 VN.n17 VN.n16 161.3
R3331 VN.n15 VN.n8 161.3
R3332 VN.n14 VN.n13 161.3
R3333 VN.n12 VN.n9 161.3
R3334 VN.n10 VN.t3 149.369
R3335 VN.n21 VN.t1 149.369
R3336 VN.n29 VN.t5 149.369
R3337 VN.n42 VN.t7 149.369
R3338 VN.n55 VN.t4 149.369
R3339 VN.n66 VN.t6 149.369
R3340 VN.n49 VN.t0 149.369
R3341 VN.n86 VN.t9 149.369
R3342 VN.n43 VN.n42 107.466
R3343 VN.n87 VN.n86 107.466
R3344 VN VN.n87 58.8164
R3345 VN.n16 VN.n15 56.5617
R3346 VN.n27 VN.n5 56.5617
R3347 VN.n61 VN.n60 56.5617
R3348 VN.n72 VN.n50 56.5617
R3349 VN.n11 VN.n10 53.6463
R3350 VN.n56 VN.n55 53.6463
R3351 VN.n36 VN.n35 41.5458
R3352 VN.n80 VN.n79 41.5458
R3353 VN.n36 VN.n1 39.6083
R3354 VN.n80 VN.n45 39.6083
R3355 VN.n14 VN.n9 24.5923
R3356 VN.n15 VN.n14 24.5923
R3357 VN.n16 VN.n7 24.5923
R3358 VN.n20 VN.n7 24.5923
R3359 VN.n23 VN.n22 24.5923
R3360 VN.n23 VN.n5 24.5923
R3361 VN.n28 VN.n27 24.5923
R3362 VN.n30 VN.n28 24.5923
R3363 VN.n34 VN.n3 24.5923
R3364 VN.n35 VN.n34 24.5923
R3365 VN.n40 VN.n1 24.5923
R3366 VN.n41 VN.n40 24.5923
R3367 VN.n60 VN.n59 24.5923
R3368 VN.n59 VN.n54 24.5923
R3369 VN.n68 VN.n50 24.5923
R3370 VN.n68 VN.n67 24.5923
R3371 VN.n65 VN.n52 24.5923
R3372 VN.n61 VN.n52 24.5923
R3373 VN.n79 VN.n78 24.5923
R3374 VN.n78 VN.n47 24.5923
R3375 VN.n74 VN.n73 24.5923
R3376 VN.n73 VN.n72 24.5923
R3377 VN.n85 VN.n84 24.5923
R3378 VN.n84 VN.n45 24.5923
R3379 VN.n10 VN.n9 20.1658
R3380 VN.n30 VN.n29 20.1658
R3381 VN.n55 VN.n54 20.1658
R3382 VN.n74 VN.n49 20.1658
R3383 VN.n21 VN.n20 12.2964
R3384 VN.n22 VN.n21 12.2964
R3385 VN.n67 VN.n66 12.2964
R3386 VN.n66 VN.n65 12.2964
R3387 VN.n57 VN.n56 5.0289
R3388 VN.n12 VN.n11 5.0289
R3389 VN.n29 VN.n3 4.42703
R3390 VN.n49 VN.n47 4.42703
R3391 VN.n42 VN.n41 3.44336
R3392 VN.n86 VN.n85 3.44336
R3393 VN.n87 VN.n44 0.278335
R3394 VN.n43 VN.n0 0.278335
R3395 VN.n83 VN.n44 0.189894
R3396 VN.n83 VN.n82 0.189894
R3397 VN.n82 VN.n81 0.189894
R3398 VN.n81 VN.n46 0.189894
R3399 VN.n77 VN.n46 0.189894
R3400 VN.n77 VN.n76 0.189894
R3401 VN.n76 VN.n75 0.189894
R3402 VN.n75 VN.n48 0.189894
R3403 VN.n71 VN.n48 0.189894
R3404 VN.n71 VN.n70 0.189894
R3405 VN.n70 VN.n69 0.189894
R3406 VN.n69 VN.n51 0.189894
R3407 VN.n64 VN.n51 0.189894
R3408 VN.n64 VN.n63 0.189894
R3409 VN.n63 VN.n62 0.189894
R3410 VN.n62 VN.n53 0.189894
R3411 VN.n58 VN.n53 0.189894
R3412 VN.n58 VN.n57 0.189894
R3413 VN.n13 VN.n12 0.189894
R3414 VN.n13 VN.n8 0.189894
R3415 VN.n17 VN.n8 0.189894
R3416 VN.n18 VN.n17 0.189894
R3417 VN.n19 VN.n18 0.189894
R3418 VN.n19 VN.n6 0.189894
R3419 VN.n24 VN.n6 0.189894
R3420 VN.n25 VN.n24 0.189894
R3421 VN.n26 VN.n25 0.189894
R3422 VN.n26 VN.n4 0.189894
R3423 VN.n31 VN.n4 0.189894
R3424 VN.n32 VN.n31 0.189894
R3425 VN.n33 VN.n32 0.189894
R3426 VN.n33 VN.n2 0.189894
R3427 VN.n37 VN.n2 0.189894
R3428 VN.n38 VN.n37 0.189894
R3429 VN.n39 VN.n38 0.189894
R3430 VN.n39 VN.n0 0.189894
R3431 VN VN.n43 0.153485
R3432 VDD2.n193 VDD2.n101 289.615
R3433 VDD2.n92 VDD2.n0 289.615
R3434 VDD2.n194 VDD2.n193 185
R3435 VDD2.n192 VDD2.n191 185
R3436 VDD2.n105 VDD2.n104 185
R3437 VDD2.n186 VDD2.n185 185
R3438 VDD2.n184 VDD2.n183 185
R3439 VDD2.n109 VDD2.n108 185
R3440 VDD2.n113 VDD2.n111 185
R3441 VDD2.n178 VDD2.n177 185
R3442 VDD2.n176 VDD2.n175 185
R3443 VDD2.n115 VDD2.n114 185
R3444 VDD2.n170 VDD2.n169 185
R3445 VDD2.n168 VDD2.n167 185
R3446 VDD2.n119 VDD2.n118 185
R3447 VDD2.n162 VDD2.n161 185
R3448 VDD2.n160 VDD2.n159 185
R3449 VDD2.n123 VDD2.n122 185
R3450 VDD2.n154 VDD2.n153 185
R3451 VDD2.n152 VDD2.n151 185
R3452 VDD2.n127 VDD2.n126 185
R3453 VDD2.n146 VDD2.n145 185
R3454 VDD2.n144 VDD2.n143 185
R3455 VDD2.n131 VDD2.n130 185
R3456 VDD2.n138 VDD2.n137 185
R3457 VDD2.n136 VDD2.n135 185
R3458 VDD2.n33 VDD2.n32 185
R3459 VDD2.n35 VDD2.n34 185
R3460 VDD2.n28 VDD2.n27 185
R3461 VDD2.n41 VDD2.n40 185
R3462 VDD2.n43 VDD2.n42 185
R3463 VDD2.n24 VDD2.n23 185
R3464 VDD2.n49 VDD2.n48 185
R3465 VDD2.n51 VDD2.n50 185
R3466 VDD2.n20 VDD2.n19 185
R3467 VDD2.n57 VDD2.n56 185
R3468 VDD2.n59 VDD2.n58 185
R3469 VDD2.n16 VDD2.n15 185
R3470 VDD2.n65 VDD2.n64 185
R3471 VDD2.n67 VDD2.n66 185
R3472 VDD2.n12 VDD2.n11 185
R3473 VDD2.n74 VDD2.n73 185
R3474 VDD2.n75 VDD2.n10 185
R3475 VDD2.n77 VDD2.n76 185
R3476 VDD2.n8 VDD2.n7 185
R3477 VDD2.n83 VDD2.n82 185
R3478 VDD2.n85 VDD2.n84 185
R3479 VDD2.n4 VDD2.n3 185
R3480 VDD2.n91 VDD2.n90 185
R3481 VDD2.n93 VDD2.n92 185
R3482 VDD2.n134 VDD2.t0 147.659
R3483 VDD2.n31 VDD2.t7 147.659
R3484 VDD2.n193 VDD2.n192 104.615
R3485 VDD2.n192 VDD2.n104 104.615
R3486 VDD2.n185 VDD2.n104 104.615
R3487 VDD2.n185 VDD2.n184 104.615
R3488 VDD2.n184 VDD2.n108 104.615
R3489 VDD2.n113 VDD2.n108 104.615
R3490 VDD2.n177 VDD2.n113 104.615
R3491 VDD2.n177 VDD2.n176 104.615
R3492 VDD2.n176 VDD2.n114 104.615
R3493 VDD2.n169 VDD2.n114 104.615
R3494 VDD2.n169 VDD2.n168 104.615
R3495 VDD2.n168 VDD2.n118 104.615
R3496 VDD2.n161 VDD2.n118 104.615
R3497 VDD2.n161 VDD2.n160 104.615
R3498 VDD2.n160 VDD2.n122 104.615
R3499 VDD2.n153 VDD2.n122 104.615
R3500 VDD2.n153 VDD2.n152 104.615
R3501 VDD2.n152 VDD2.n126 104.615
R3502 VDD2.n145 VDD2.n126 104.615
R3503 VDD2.n145 VDD2.n144 104.615
R3504 VDD2.n144 VDD2.n130 104.615
R3505 VDD2.n137 VDD2.n130 104.615
R3506 VDD2.n137 VDD2.n136 104.615
R3507 VDD2.n34 VDD2.n33 104.615
R3508 VDD2.n34 VDD2.n27 104.615
R3509 VDD2.n41 VDD2.n27 104.615
R3510 VDD2.n42 VDD2.n41 104.615
R3511 VDD2.n42 VDD2.n23 104.615
R3512 VDD2.n49 VDD2.n23 104.615
R3513 VDD2.n50 VDD2.n49 104.615
R3514 VDD2.n50 VDD2.n19 104.615
R3515 VDD2.n57 VDD2.n19 104.615
R3516 VDD2.n58 VDD2.n57 104.615
R3517 VDD2.n58 VDD2.n15 104.615
R3518 VDD2.n65 VDD2.n15 104.615
R3519 VDD2.n66 VDD2.n65 104.615
R3520 VDD2.n66 VDD2.n11 104.615
R3521 VDD2.n74 VDD2.n11 104.615
R3522 VDD2.n75 VDD2.n74 104.615
R3523 VDD2.n76 VDD2.n75 104.615
R3524 VDD2.n76 VDD2.n7 104.615
R3525 VDD2.n83 VDD2.n7 104.615
R3526 VDD2.n84 VDD2.n83 104.615
R3527 VDD2.n84 VDD2.n3 104.615
R3528 VDD2.n91 VDD2.n3 104.615
R3529 VDD2.n92 VDD2.n91 104.615
R3530 VDD2.n100 VDD2.n99 63.0576
R3531 VDD2 VDD2.n201 63.0548
R3532 VDD2.n200 VDD2.n199 61.07
R3533 VDD2.n98 VDD2.n97 61.0699
R3534 VDD2.n136 VDD2.t0 52.3082
R3535 VDD2.n33 VDD2.t7 52.3082
R3536 VDD2.n98 VDD2.n96 51.9762
R3537 VDD2.n198 VDD2.n100 51.7756
R3538 VDD2.n198 VDD2.n197 49.252
R3539 VDD2.n135 VDD2.n134 15.6677
R3540 VDD2.n32 VDD2.n31 15.6677
R3541 VDD2.n111 VDD2.n109 13.1884
R3542 VDD2.n77 VDD2.n8 13.1884
R3543 VDD2.n183 VDD2.n182 12.8005
R3544 VDD2.n179 VDD2.n178 12.8005
R3545 VDD2.n138 VDD2.n133 12.8005
R3546 VDD2.n35 VDD2.n30 12.8005
R3547 VDD2.n78 VDD2.n10 12.8005
R3548 VDD2.n82 VDD2.n81 12.8005
R3549 VDD2.n186 VDD2.n107 12.0247
R3550 VDD2.n175 VDD2.n112 12.0247
R3551 VDD2.n139 VDD2.n131 12.0247
R3552 VDD2.n36 VDD2.n28 12.0247
R3553 VDD2.n73 VDD2.n72 12.0247
R3554 VDD2.n85 VDD2.n6 12.0247
R3555 VDD2.n187 VDD2.n105 11.249
R3556 VDD2.n174 VDD2.n115 11.249
R3557 VDD2.n143 VDD2.n142 11.249
R3558 VDD2.n40 VDD2.n39 11.249
R3559 VDD2.n71 VDD2.n12 11.249
R3560 VDD2.n86 VDD2.n4 11.249
R3561 VDD2.n191 VDD2.n190 10.4732
R3562 VDD2.n171 VDD2.n170 10.4732
R3563 VDD2.n146 VDD2.n129 10.4732
R3564 VDD2.n43 VDD2.n26 10.4732
R3565 VDD2.n68 VDD2.n67 10.4732
R3566 VDD2.n90 VDD2.n89 10.4732
R3567 VDD2.n194 VDD2.n103 9.69747
R3568 VDD2.n167 VDD2.n117 9.69747
R3569 VDD2.n147 VDD2.n127 9.69747
R3570 VDD2.n44 VDD2.n24 9.69747
R3571 VDD2.n64 VDD2.n14 9.69747
R3572 VDD2.n93 VDD2.n2 9.69747
R3573 VDD2.n197 VDD2.n196 9.45567
R3574 VDD2.n96 VDD2.n95 9.45567
R3575 VDD2.n121 VDD2.n120 9.3005
R3576 VDD2.n164 VDD2.n163 9.3005
R3577 VDD2.n166 VDD2.n165 9.3005
R3578 VDD2.n117 VDD2.n116 9.3005
R3579 VDD2.n172 VDD2.n171 9.3005
R3580 VDD2.n174 VDD2.n173 9.3005
R3581 VDD2.n112 VDD2.n110 9.3005
R3582 VDD2.n180 VDD2.n179 9.3005
R3583 VDD2.n196 VDD2.n195 9.3005
R3584 VDD2.n103 VDD2.n102 9.3005
R3585 VDD2.n190 VDD2.n189 9.3005
R3586 VDD2.n188 VDD2.n187 9.3005
R3587 VDD2.n107 VDD2.n106 9.3005
R3588 VDD2.n182 VDD2.n181 9.3005
R3589 VDD2.n158 VDD2.n157 9.3005
R3590 VDD2.n156 VDD2.n155 9.3005
R3591 VDD2.n125 VDD2.n124 9.3005
R3592 VDD2.n150 VDD2.n149 9.3005
R3593 VDD2.n148 VDD2.n147 9.3005
R3594 VDD2.n129 VDD2.n128 9.3005
R3595 VDD2.n142 VDD2.n141 9.3005
R3596 VDD2.n140 VDD2.n139 9.3005
R3597 VDD2.n133 VDD2.n132 9.3005
R3598 VDD2.n95 VDD2.n94 9.3005
R3599 VDD2.n2 VDD2.n1 9.3005
R3600 VDD2.n89 VDD2.n88 9.3005
R3601 VDD2.n87 VDD2.n86 9.3005
R3602 VDD2.n6 VDD2.n5 9.3005
R3603 VDD2.n81 VDD2.n80 9.3005
R3604 VDD2.n53 VDD2.n52 9.3005
R3605 VDD2.n22 VDD2.n21 9.3005
R3606 VDD2.n47 VDD2.n46 9.3005
R3607 VDD2.n45 VDD2.n44 9.3005
R3608 VDD2.n26 VDD2.n25 9.3005
R3609 VDD2.n39 VDD2.n38 9.3005
R3610 VDD2.n37 VDD2.n36 9.3005
R3611 VDD2.n30 VDD2.n29 9.3005
R3612 VDD2.n55 VDD2.n54 9.3005
R3613 VDD2.n18 VDD2.n17 9.3005
R3614 VDD2.n61 VDD2.n60 9.3005
R3615 VDD2.n63 VDD2.n62 9.3005
R3616 VDD2.n14 VDD2.n13 9.3005
R3617 VDD2.n69 VDD2.n68 9.3005
R3618 VDD2.n71 VDD2.n70 9.3005
R3619 VDD2.n72 VDD2.n9 9.3005
R3620 VDD2.n79 VDD2.n78 9.3005
R3621 VDD2.n195 VDD2.n101 8.92171
R3622 VDD2.n166 VDD2.n119 8.92171
R3623 VDD2.n151 VDD2.n150 8.92171
R3624 VDD2.n48 VDD2.n47 8.92171
R3625 VDD2.n63 VDD2.n16 8.92171
R3626 VDD2.n94 VDD2.n0 8.92171
R3627 VDD2.n163 VDD2.n162 8.14595
R3628 VDD2.n154 VDD2.n125 8.14595
R3629 VDD2.n51 VDD2.n22 8.14595
R3630 VDD2.n60 VDD2.n59 8.14595
R3631 VDD2.n159 VDD2.n121 7.3702
R3632 VDD2.n155 VDD2.n123 7.3702
R3633 VDD2.n52 VDD2.n20 7.3702
R3634 VDD2.n56 VDD2.n18 7.3702
R3635 VDD2.n159 VDD2.n158 6.59444
R3636 VDD2.n158 VDD2.n123 6.59444
R3637 VDD2.n55 VDD2.n20 6.59444
R3638 VDD2.n56 VDD2.n55 6.59444
R3639 VDD2.n162 VDD2.n121 5.81868
R3640 VDD2.n155 VDD2.n154 5.81868
R3641 VDD2.n52 VDD2.n51 5.81868
R3642 VDD2.n59 VDD2.n18 5.81868
R3643 VDD2.n197 VDD2.n101 5.04292
R3644 VDD2.n163 VDD2.n119 5.04292
R3645 VDD2.n151 VDD2.n125 5.04292
R3646 VDD2.n48 VDD2.n22 5.04292
R3647 VDD2.n60 VDD2.n16 5.04292
R3648 VDD2.n96 VDD2.n0 5.04292
R3649 VDD2.n134 VDD2.n132 4.38563
R3650 VDD2.n31 VDD2.n29 4.38563
R3651 VDD2.n195 VDD2.n194 4.26717
R3652 VDD2.n167 VDD2.n166 4.26717
R3653 VDD2.n150 VDD2.n127 4.26717
R3654 VDD2.n47 VDD2.n24 4.26717
R3655 VDD2.n64 VDD2.n63 4.26717
R3656 VDD2.n94 VDD2.n93 4.26717
R3657 VDD2.n191 VDD2.n103 3.49141
R3658 VDD2.n170 VDD2.n117 3.49141
R3659 VDD2.n147 VDD2.n146 3.49141
R3660 VDD2.n44 VDD2.n43 3.49141
R3661 VDD2.n67 VDD2.n14 3.49141
R3662 VDD2.n90 VDD2.n2 3.49141
R3663 VDD2.n200 VDD2.n198 2.72464
R3664 VDD2.n190 VDD2.n105 2.71565
R3665 VDD2.n171 VDD2.n115 2.71565
R3666 VDD2.n143 VDD2.n129 2.71565
R3667 VDD2.n40 VDD2.n26 2.71565
R3668 VDD2.n68 VDD2.n12 2.71565
R3669 VDD2.n89 VDD2.n4 2.71565
R3670 VDD2.n187 VDD2.n186 1.93989
R3671 VDD2.n175 VDD2.n174 1.93989
R3672 VDD2.n142 VDD2.n131 1.93989
R3673 VDD2.n39 VDD2.n28 1.93989
R3674 VDD2.n73 VDD2.n71 1.93989
R3675 VDD2.n86 VDD2.n85 1.93989
R3676 VDD2.n183 VDD2.n107 1.16414
R3677 VDD2.n178 VDD2.n112 1.16414
R3678 VDD2.n139 VDD2.n138 1.16414
R3679 VDD2.n36 VDD2.n35 1.16414
R3680 VDD2.n72 VDD2.n10 1.16414
R3681 VDD2.n82 VDD2.n6 1.16414
R3682 VDD2.n201 VDD2.t5 1.12935
R3683 VDD2.n201 VDD2.t1 1.12935
R3684 VDD2.n199 VDD2.t9 1.12935
R3685 VDD2.n199 VDD2.t3 1.12935
R3686 VDD2.n99 VDD2.t4 1.12935
R3687 VDD2.n99 VDD2.t2 1.12935
R3688 VDD2.n97 VDD2.t6 1.12935
R3689 VDD2.n97 VDD2.t8 1.12935
R3690 VDD2 VDD2.n200 0.739724
R3691 VDD2.n100 VDD2.n98 0.626188
R3692 VDD2.n182 VDD2.n109 0.388379
R3693 VDD2.n179 VDD2.n111 0.388379
R3694 VDD2.n135 VDD2.n133 0.388379
R3695 VDD2.n32 VDD2.n30 0.388379
R3696 VDD2.n78 VDD2.n77 0.388379
R3697 VDD2.n81 VDD2.n8 0.388379
R3698 VDD2.n196 VDD2.n102 0.155672
R3699 VDD2.n189 VDD2.n102 0.155672
R3700 VDD2.n189 VDD2.n188 0.155672
R3701 VDD2.n188 VDD2.n106 0.155672
R3702 VDD2.n181 VDD2.n106 0.155672
R3703 VDD2.n181 VDD2.n180 0.155672
R3704 VDD2.n180 VDD2.n110 0.155672
R3705 VDD2.n173 VDD2.n110 0.155672
R3706 VDD2.n173 VDD2.n172 0.155672
R3707 VDD2.n172 VDD2.n116 0.155672
R3708 VDD2.n165 VDD2.n116 0.155672
R3709 VDD2.n165 VDD2.n164 0.155672
R3710 VDD2.n164 VDD2.n120 0.155672
R3711 VDD2.n157 VDD2.n120 0.155672
R3712 VDD2.n157 VDD2.n156 0.155672
R3713 VDD2.n156 VDD2.n124 0.155672
R3714 VDD2.n149 VDD2.n124 0.155672
R3715 VDD2.n149 VDD2.n148 0.155672
R3716 VDD2.n148 VDD2.n128 0.155672
R3717 VDD2.n141 VDD2.n128 0.155672
R3718 VDD2.n141 VDD2.n140 0.155672
R3719 VDD2.n140 VDD2.n132 0.155672
R3720 VDD2.n37 VDD2.n29 0.155672
R3721 VDD2.n38 VDD2.n37 0.155672
R3722 VDD2.n38 VDD2.n25 0.155672
R3723 VDD2.n45 VDD2.n25 0.155672
R3724 VDD2.n46 VDD2.n45 0.155672
R3725 VDD2.n46 VDD2.n21 0.155672
R3726 VDD2.n53 VDD2.n21 0.155672
R3727 VDD2.n54 VDD2.n53 0.155672
R3728 VDD2.n54 VDD2.n17 0.155672
R3729 VDD2.n61 VDD2.n17 0.155672
R3730 VDD2.n62 VDD2.n61 0.155672
R3731 VDD2.n62 VDD2.n13 0.155672
R3732 VDD2.n69 VDD2.n13 0.155672
R3733 VDD2.n70 VDD2.n69 0.155672
R3734 VDD2.n70 VDD2.n9 0.155672
R3735 VDD2.n79 VDD2.n9 0.155672
R3736 VDD2.n80 VDD2.n79 0.155672
R3737 VDD2.n80 VDD2.n5 0.155672
R3738 VDD2.n87 VDD2.n5 0.155672
R3739 VDD2.n88 VDD2.n87 0.155672
R3740 VDD2.n88 VDD2.n1 0.155672
R3741 VDD2.n95 VDD2.n1 0.155672
C0 VDD1 VP 16.0665f
C1 VTAIL VN 16.1027f
C2 VDD1 VN 0.154099f
C3 VTAIL VDD2 12.9592f
C4 VDD1 VDD2 2.32391f
C5 VTAIL VDD1 12.907701f
C6 VP VN 9.7558f
C7 VP VDD2 0.613546f
C8 VN VDD2 15.6118f
C9 VTAIL VP 16.117f
C10 VDD2 B 8.44562f
C11 VDD1 B 8.425789f
C12 VTAIL B 10.604574f
C13 VN B 19.67078f
C14 VP B 18.140017f
C15 VDD2.n0 B 0.032822f
C16 VDD2.n1 B 0.023578f
C17 VDD2.n2 B 0.01267f
C18 VDD2.n3 B 0.029946f
C19 VDD2.n4 B 0.013415f
C20 VDD2.n5 B 0.023578f
C21 VDD2.n6 B 0.01267f
C22 VDD2.n7 B 0.029946f
C23 VDD2.n8 B 0.013042f
C24 VDD2.n9 B 0.023578f
C25 VDD2.n10 B 0.013415f
C26 VDD2.n11 B 0.029946f
C27 VDD2.n12 B 0.013415f
C28 VDD2.n13 B 0.023578f
C29 VDD2.n14 B 0.01267f
C30 VDD2.n15 B 0.029946f
C31 VDD2.n16 B 0.013415f
C32 VDD2.n17 B 0.023578f
C33 VDD2.n18 B 0.01267f
C34 VDD2.n19 B 0.029946f
C35 VDD2.n20 B 0.013415f
C36 VDD2.n21 B 0.023578f
C37 VDD2.n22 B 0.01267f
C38 VDD2.n23 B 0.029946f
C39 VDD2.n24 B 0.013415f
C40 VDD2.n25 B 0.023578f
C41 VDD2.n26 B 0.01267f
C42 VDD2.n27 B 0.029946f
C43 VDD2.n28 B 0.013415f
C44 VDD2.n29 B 1.80846f
C45 VDD2.n30 B 0.01267f
C46 VDD2.t7 B 0.049583f
C47 VDD2.n31 B 0.168794f
C48 VDD2.n32 B 0.01769f
C49 VDD2.n33 B 0.02246f
C50 VDD2.n34 B 0.029946f
C51 VDD2.n35 B 0.013415f
C52 VDD2.n36 B 0.01267f
C53 VDD2.n37 B 0.023578f
C54 VDD2.n38 B 0.023578f
C55 VDD2.n39 B 0.01267f
C56 VDD2.n40 B 0.013415f
C57 VDD2.n41 B 0.029946f
C58 VDD2.n42 B 0.029946f
C59 VDD2.n43 B 0.013415f
C60 VDD2.n44 B 0.01267f
C61 VDD2.n45 B 0.023578f
C62 VDD2.n46 B 0.023578f
C63 VDD2.n47 B 0.01267f
C64 VDD2.n48 B 0.013415f
C65 VDD2.n49 B 0.029946f
C66 VDD2.n50 B 0.029946f
C67 VDD2.n51 B 0.013415f
C68 VDD2.n52 B 0.01267f
C69 VDD2.n53 B 0.023578f
C70 VDD2.n54 B 0.023578f
C71 VDD2.n55 B 0.01267f
C72 VDD2.n56 B 0.013415f
C73 VDD2.n57 B 0.029946f
C74 VDD2.n58 B 0.029946f
C75 VDD2.n59 B 0.013415f
C76 VDD2.n60 B 0.01267f
C77 VDD2.n61 B 0.023578f
C78 VDD2.n62 B 0.023578f
C79 VDD2.n63 B 0.01267f
C80 VDD2.n64 B 0.013415f
C81 VDD2.n65 B 0.029946f
C82 VDD2.n66 B 0.029946f
C83 VDD2.n67 B 0.013415f
C84 VDD2.n68 B 0.01267f
C85 VDD2.n69 B 0.023578f
C86 VDD2.n70 B 0.023578f
C87 VDD2.n71 B 0.01267f
C88 VDD2.n72 B 0.01267f
C89 VDD2.n73 B 0.013415f
C90 VDD2.n74 B 0.029946f
C91 VDD2.n75 B 0.029946f
C92 VDD2.n76 B 0.029946f
C93 VDD2.n77 B 0.013042f
C94 VDD2.n78 B 0.01267f
C95 VDD2.n79 B 0.023578f
C96 VDD2.n80 B 0.023578f
C97 VDD2.n81 B 0.01267f
C98 VDD2.n82 B 0.013415f
C99 VDD2.n83 B 0.029946f
C100 VDD2.n84 B 0.029946f
C101 VDD2.n85 B 0.013415f
C102 VDD2.n86 B 0.01267f
C103 VDD2.n87 B 0.023578f
C104 VDD2.n88 B 0.023578f
C105 VDD2.n89 B 0.01267f
C106 VDD2.n90 B 0.013415f
C107 VDD2.n91 B 0.029946f
C108 VDD2.n92 B 0.064266f
C109 VDD2.n93 B 0.013415f
C110 VDD2.n94 B 0.01267f
C111 VDD2.n95 B 0.055143f
C112 VDD2.n96 B 0.065442f
C113 VDD2.t6 B 0.326801f
C114 VDD2.t8 B 0.326801f
C115 VDD2.n97 B 2.97429f
C116 VDD2.n98 B 0.690125f
C117 VDD2.t4 B 0.326801f
C118 VDD2.t2 B 0.326801f
C119 VDD2.n99 B 2.99203f
C120 VDD2.n100 B 3.18143f
C121 VDD2.n101 B 0.032822f
C122 VDD2.n102 B 0.023578f
C123 VDD2.n103 B 0.01267f
C124 VDD2.n104 B 0.029946f
C125 VDD2.n105 B 0.013415f
C126 VDD2.n106 B 0.023578f
C127 VDD2.n107 B 0.01267f
C128 VDD2.n108 B 0.029946f
C129 VDD2.n109 B 0.013042f
C130 VDD2.n110 B 0.023578f
C131 VDD2.n111 B 0.013042f
C132 VDD2.n112 B 0.01267f
C133 VDD2.n113 B 0.029946f
C134 VDD2.n114 B 0.029946f
C135 VDD2.n115 B 0.013415f
C136 VDD2.n116 B 0.023578f
C137 VDD2.n117 B 0.01267f
C138 VDD2.n118 B 0.029946f
C139 VDD2.n119 B 0.013415f
C140 VDD2.n120 B 0.023578f
C141 VDD2.n121 B 0.01267f
C142 VDD2.n122 B 0.029946f
C143 VDD2.n123 B 0.013415f
C144 VDD2.n124 B 0.023578f
C145 VDD2.n125 B 0.01267f
C146 VDD2.n126 B 0.029946f
C147 VDD2.n127 B 0.013415f
C148 VDD2.n128 B 0.023578f
C149 VDD2.n129 B 0.01267f
C150 VDD2.n130 B 0.029946f
C151 VDD2.n131 B 0.013415f
C152 VDD2.n132 B 1.80846f
C153 VDD2.n133 B 0.01267f
C154 VDD2.t0 B 0.049583f
C155 VDD2.n134 B 0.168794f
C156 VDD2.n135 B 0.01769f
C157 VDD2.n136 B 0.02246f
C158 VDD2.n137 B 0.029946f
C159 VDD2.n138 B 0.013415f
C160 VDD2.n139 B 0.01267f
C161 VDD2.n140 B 0.023578f
C162 VDD2.n141 B 0.023578f
C163 VDD2.n142 B 0.01267f
C164 VDD2.n143 B 0.013415f
C165 VDD2.n144 B 0.029946f
C166 VDD2.n145 B 0.029946f
C167 VDD2.n146 B 0.013415f
C168 VDD2.n147 B 0.01267f
C169 VDD2.n148 B 0.023578f
C170 VDD2.n149 B 0.023578f
C171 VDD2.n150 B 0.01267f
C172 VDD2.n151 B 0.013415f
C173 VDD2.n152 B 0.029946f
C174 VDD2.n153 B 0.029946f
C175 VDD2.n154 B 0.013415f
C176 VDD2.n155 B 0.01267f
C177 VDD2.n156 B 0.023578f
C178 VDD2.n157 B 0.023578f
C179 VDD2.n158 B 0.01267f
C180 VDD2.n159 B 0.013415f
C181 VDD2.n160 B 0.029946f
C182 VDD2.n161 B 0.029946f
C183 VDD2.n162 B 0.013415f
C184 VDD2.n163 B 0.01267f
C185 VDD2.n164 B 0.023578f
C186 VDD2.n165 B 0.023578f
C187 VDD2.n166 B 0.01267f
C188 VDD2.n167 B 0.013415f
C189 VDD2.n168 B 0.029946f
C190 VDD2.n169 B 0.029946f
C191 VDD2.n170 B 0.013415f
C192 VDD2.n171 B 0.01267f
C193 VDD2.n172 B 0.023578f
C194 VDD2.n173 B 0.023578f
C195 VDD2.n174 B 0.01267f
C196 VDD2.n175 B 0.013415f
C197 VDD2.n176 B 0.029946f
C198 VDD2.n177 B 0.029946f
C199 VDD2.n178 B 0.013415f
C200 VDD2.n179 B 0.01267f
C201 VDD2.n180 B 0.023578f
C202 VDD2.n181 B 0.023578f
C203 VDD2.n182 B 0.01267f
C204 VDD2.n183 B 0.013415f
C205 VDD2.n184 B 0.029946f
C206 VDD2.n185 B 0.029946f
C207 VDD2.n186 B 0.013415f
C208 VDD2.n187 B 0.01267f
C209 VDD2.n188 B 0.023578f
C210 VDD2.n189 B 0.023578f
C211 VDD2.n190 B 0.01267f
C212 VDD2.n191 B 0.013415f
C213 VDD2.n192 B 0.029946f
C214 VDD2.n193 B 0.064266f
C215 VDD2.n194 B 0.013415f
C216 VDD2.n195 B 0.01267f
C217 VDD2.n196 B 0.055143f
C218 VDD2.n197 B 0.052196f
C219 VDD2.n198 B 3.20889f
C220 VDD2.t9 B 0.326801f
C221 VDD2.t3 B 0.326801f
C222 VDD2.n199 B 2.97429f
C223 VDD2.n200 B 0.458385f
C224 VDD2.t5 B 0.326801f
C225 VDD2.t1 B 0.326801f
C226 VDD2.n201 B 2.99199f
C227 VN.n0 B 0.025647f
C228 VN.t7 B 2.65483f
C229 VN.n1 B 0.038642f
C230 VN.n2 B 0.019454f
C231 VN.n3 B 0.021472f
C232 VN.n4 B 0.019454f
C233 VN.n5 B 0.032586f
C234 VN.n6 B 0.019454f
C235 VN.t1 B 2.65483f
C236 VN.n7 B 0.036076f
C237 VN.n8 B 0.019454f
C238 VN.n9 B 0.03287f
C239 VN.t2 B 2.84704f
C240 VN.t3 B 2.65483f
C241 VN.n10 B 0.985498f
C242 VN.n11 B 0.950884f
C243 VN.n12 B 0.204802f
C244 VN.n13 B 0.019454f
C245 VN.n14 B 0.036076f
C246 VN.n15 B 0.023974f
C247 VN.n16 B 0.032586f
C248 VN.n17 B 0.019454f
C249 VN.n18 B 0.019454f
C250 VN.n19 B 0.019454f
C251 VN.n20 B 0.027171f
C252 VN.n21 B 0.919896f
C253 VN.n22 B 0.027171f
C254 VN.n23 B 0.036076f
C255 VN.n24 B 0.019454f
C256 VN.n25 B 0.019454f
C257 VN.n26 B 0.019454f
C258 VN.n27 B 0.023974f
C259 VN.n28 B 0.036076f
C260 VN.t5 B 2.65483f
C261 VN.n29 B 0.919896f
C262 VN.n30 B 0.03287f
C263 VN.n31 B 0.019454f
C264 VN.n32 B 0.019454f
C265 VN.n33 B 0.019454f
C266 VN.n34 B 0.036076f
C267 VN.n35 B 0.038256f
C268 VN.n36 B 0.015737f
C269 VN.n37 B 0.019454f
C270 VN.n38 B 0.019454f
C271 VN.n39 B 0.019454f
C272 VN.n40 B 0.036076f
C273 VN.n41 B 0.02076f
C274 VN.n42 B 0.983681f
C275 VN.n43 B 0.036265f
C276 VN.n44 B 0.025647f
C277 VN.t9 B 2.65483f
C278 VN.n45 B 0.038642f
C279 VN.n46 B 0.019454f
C280 VN.n47 B 0.021472f
C281 VN.n48 B 0.019454f
C282 VN.t0 B 2.65483f
C283 VN.n49 B 0.919896f
C284 VN.n50 B 0.032586f
C285 VN.n51 B 0.019454f
C286 VN.t6 B 2.65483f
C287 VN.n52 B 0.036076f
C288 VN.n53 B 0.019454f
C289 VN.n54 B 0.03287f
C290 VN.t8 B 2.84704f
C291 VN.t4 B 2.65483f
C292 VN.n55 B 0.985498f
C293 VN.n56 B 0.950884f
C294 VN.n57 B 0.204802f
C295 VN.n58 B 0.019454f
C296 VN.n59 B 0.036076f
C297 VN.n60 B 0.023974f
C298 VN.n61 B 0.032586f
C299 VN.n62 B 0.019454f
C300 VN.n63 B 0.019454f
C301 VN.n64 B 0.019454f
C302 VN.n65 B 0.027171f
C303 VN.n66 B 0.919896f
C304 VN.n67 B 0.027171f
C305 VN.n68 B 0.036076f
C306 VN.n69 B 0.019454f
C307 VN.n70 B 0.019454f
C308 VN.n71 B 0.019454f
C309 VN.n72 B 0.023974f
C310 VN.n73 B 0.036076f
C311 VN.n74 B 0.03287f
C312 VN.n75 B 0.019454f
C313 VN.n76 B 0.019454f
C314 VN.n77 B 0.019454f
C315 VN.n78 B 0.036076f
C316 VN.n79 B 0.038256f
C317 VN.n80 B 0.015737f
C318 VN.n81 B 0.019454f
C319 VN.n82 B 0.019454f
C320 VN.n83 B 0.019454f
C321 VN.n84 B 0.036076f
C322 VN.n85 B 0.02076f
C323 VN.n86 B 0.983681f
C324 VN.n87 B 1.36864f
C325 VTAIL.t0 B 0.330614f
C326 VTAIL.t3 B 0.330614f
C327 VTAIL.n0 B 2.93646f
C328 VTAIL.n1 B 0.539952f
C329 VTAIL.n2 B 0.033205f
C330 VTAIL.n3 B 0.023853f
C331 VTAIL.n4 B 0.012817f
C332 VTAIL.n5 B 0.030296f
C333 VTAIL.n6 B 0.013571f
C334 VTAIL.n7 B 0.023853f
C335 VTAIL.n8 B 0.012817f
C336 VTAIL.n9 B 0.030296f
C337 VTAIL.n10 B 0.013194f
C338 VTAIL.n11 B 0.023853f
C339 VTAIL.n12 B 0.013571f
C340 VTAIL.n13 B 0.030296f
C341 VTAIL.n14 B 0.013571f
C342 VTAIL.n15 B 0.023853f
C343 VTAIL.n16 B 0.012817f
C344 VTAIL.n17 B 0.030296f
C345 VTAIL.n18 B 0.013571f
C346 VTAIL.n19 B 0.023853f
C347 VTAIL.n20 B 0.012817f
C348 VTAIL.n21 B 0.030296f
C349 VTAIL.n22 B 0.013571f
C350 VTAIL.n23 B 0.023853f
C351 VTAIL.n24 B 0.012817f
C352 VTAIL.n25 B 0.030296f
C353 VTAIL.n26 B 0.013571f
C354 VTAIL.n27 B 0.023853f
C355 VTAIL.n28 B 0.012817f
C356 VTAIL.n29 B 0.030296f
C357 VTAIL.n30 B 0.013571f
C358 VTAIL.n31 B 1.82956f
C359 VTAIL.n32 B 0.012817f
C360 VTAIL.t17 B 0.050162f
C361 VTAIL.n33 B 0.170763f
C362 VTAIL.n34 B 0.017897f
C363 VTAIL.n35 B 0.022722f
C364 VTAIL.n36 B 0.030296f
C365 VTAIL.n37 B 0.013571f
C366 VTAIL.n38 B 0.012817f
C367 VTAIL.n39 B 0.023853f
C368 VTAIL.n40 B 0.023853f
C369 VTAIL.n41 B 0.012817f
C370 VTAIL.n42 B 0.013571f
C371 VTAIL.n43 B 0.030296f
C372 VTAIL.n44 B 0.030296f
C373 VTAIL.n45 B 0.013571f
C374 VTAIL.n46 B 0.012817f
C375 VTAIL.n47 B 0.023853f
C376 VTAIL.n48 B 0.023853f
C377 VTAIL.n49 B 0.012817f
C378 VTAIL.n50 B 0.013571f
C379 VTAIL.n51 B 0.030296f
C380 VTAIL.n52 B 0.030296f
C381 VTAIL.n53 B 0.013571f
C382 VTAIL.n54 B 0.012817f
C383 VTAIL.n55 B 0.023853f
C384 VTAIL.n56 B 0.023853f
C385 VTAIL.n57 B 0.012817f
C386 VTAIL.n58 B 0.013571f
C387 VTAIL.n59 B 0.030296f
C388 VTAIL.n60 B 0.030296f
C389 VTAIL.n61 B 0.013571f
C390 VTAIL.n62 B 0.012817f
C391 VTAIL.n63 B 0.023853f
C392 VTAIL.n64 B 0.023853f
C393 VTAIL.n65 B 0.012817f
C394 VTAIL.n66 B 0.013571f
C395 VTAIL.n67 B 0.030296f
C396 VTAIL.n68 B 0.030296f
C397 VTAIL.n69 B 0.013571f
C398 VTAIL.n70 B 0.012817f
C399 VTAIL.n71 B 0.023853f
C400 VTAIL.n72 B 0.023853f
C401 VTAIL.n73 B 0.012817f
C402 VTAIL.n74 B 0.012817f
C403 VTAIL.n75 B 0.013571f
C404 VTAIL.n76 B 0.030296f
C405 VTAIL.n77 B 0.030296f
C406 VTAIL.n78 B 0.030296f
C407 VTAIL.n79 B 0.013194f
C408 VTAIL.n80 B 0.012817f
C409 VTAIL.n81 B 0.023853f
C410 VTAIL.n82 B 0.023853f
C411 VTAIL.n83 B 0.012817f
C412 VTAIL.n84 B 0.013571f
C413 VTAIL.n85 B 0.030296f
C414 VTAIL.n86 B 0.030296f
C415 VTAIL.n87 B 0.013571f
C416 VTAIL.n88 B 0.012817f
C417 VTAIL.n89 B 0.023853f
C418 VTAIL.n90 B 0.023853f
C419 VTAIL.n91 B 0.012817f
C420 VTAIL.n92 B 0.013571f
C421 VTAIL.n93 B 0.030296f
C422 VTAIL.n94 B 0.065016f
C423 VTAIL.n95 B 0.013571f
C424 VTAIL.n96 B 0.012817f
C425 VTAIL.n97 B 0.055786f
C426 VTAIL.n98 B 0.03634f
C427 VTAIL.n99 B 0.370911f
C428 VTAIL.t12 B 0.330614f
C429 VTAIL.t16 B 0.330614f
C430 VTAIL.n100 B 2.93646f
C431 VTAIL.n101 B 0.656399f
C432 VTAIL.t14 B 0.330614f
C433 VTAIL.t11 B 0.330614f
C434 VTAIL.n102 B 2.93646f
C435 VTAIL.n103 B 2.35194f
C436 VTAIL.t9 B 0.330614f
C437 VTAIL.t2 B 0.330614f
C438 VTAIL.n104 B 2.93648f
C439 VTAIL.n105 B 2.35193f
C440 VTAIL.t8 B 0.330614f
C441 VTAIL.t4 B 0.330614f
C442 VTAIL.n106 B 2.93648f
C443 VTAIL.n107 B 0.656386f
C444 VTAIL.n108 B 0.033205f
C445 VTAIL.n109 B 0.023853f
C446 VTAIL.n110 B 0.012817f
C447 VTAIL.n111 B 0.030296f
C448 VTAIL.n112 B 0.013571f
C449 VTAIL.n113 B 0.023853f
C450 VTAIL.n114 B 0.012817f
C451 VTAIL.n115 B 0.030296f
C452 VTAIL.n116 B 0.013194f
C453 VTAIL.n117 B 0.023853f
C454 VTAIL.n118 B 0.013194f
C455 VTAIL.n119 B 0.012817f
C456 VTAIL.n120 B 0.030296f
C457 VTAIL.n121 B 0.030296f
C458 VTAIL.n122 B 0.013571f
C459 VTAIL.n123 B 0.023853f
C460 VTAIL.n124 B 0.012817f
C461 VTAIL.n125 B 0.030296f
C462 VTAIL.n126 B 0.013571f
C463 VTAIL.n127 B 0.023853f
C464 VTAIL.n128 B 0.012817f
C465 VTAIL.n129 B 0.030296f
C466 VTAIL.n130 B 0.013571f
C467 VTAIL.n131 B 0.023853f
C468 VTAIL.n132 B 0.012817f
C469 VTAIL.n133 B 0.030296f
C470 VTAIL.n134 B 0.013571f
C471 VTAIL.n135 B 0.023853f
C472 VTAIL.n136 B 0.012817f
C473 VTAIL.n137 B 0.030296f
C474 VTAIL.n138 B 0.013571f
C475 VTAIL.n139 B 1.82956f
C476 VTAIL.n140 B 0.012817f
C477 VTAIL.t5 B 0.050162f
C478 VTAIL.n141 B 0.170763f
C479 VTAIL.n142 B 0.017897f
C480 VTAIL.n143 B 0.022722f
C481 VTAIL.n144 B 0.030296f
C482 VTAIL.n145 B 0.013571f
C483 VTAIL.n146 B 0.012817f
C484 VTAIL.n147 B 0.023853f
C485 VTAIL.n148 B 0.023853f
C486 VTAIL.n149 B 0.012817f
C487 VTAIL.n150 B 0.013571f
C488 VTAIL.n151 B 0.030296f
C489 VTAIL.n152 B 0.030296f
C490 VTAIL.n153 B 0.013571f
C491 VTAIL.n154 B 0.012817f
C492 VTAIL.n155 B 0.023853f
C493 VTAIL.n156 B 0.023853f
C494 VTAIL.n157 B 0.012817f
C495 VTAIL.n158 B 0.013571f
C496 VTAIL.n159 B 0.030296f
C497 VTAIL.n160 B 0.030296f
C498 VTAIL.n161 B 0.013571f
C499 VTAIL.n162 B 0.012817f
C500 VTAIL.n163 B 0.023853f
C501 VTAIL.n164 B 0.023853f
C502 VTAIL.n165 B 0.012817f
C503 VTAIL.n166 B 0.013571f
C504 VTAIL.n167 B 0.030296f
C505 VTAIL.n168 B 0.030296f
C506 VTAIL.n169 B 0.013571f
C507 VTAIL.n170 B 0.012817f
C508 VTAIL.n171 B 0.023853f
C509 VTAIL.n172 B 0.023853f
C510 VTAIL.n173 B 0.012817f
C511 VTAIL.n174 B 0.013571f
C512 VTAIL.n175 B 0.030296f
C513 VTAIL.n176 B 0.030296f
C514 VTAIL.n177 B 0.013571f
C515 VTAIL.n178 B 0.012817f
C516 VTAIL.n179 B 0.023853f
C517 VTAIL.n180 B 0.023853f
C518 VTAIL.n181 B 0.012817f
C519 VTAIL.n182 B 0.013571f
C520 VTAIL.n183 B 0.030296f
C521 VTAIL.n184 B 0.030296f
C522 VTAIL.n185 B 0.013571f
C523 VTAIL.n186 B 0.012817f
C524 VTAIL.n187 B 0.023853f
C525 VTAIL.n188 B 0.023853f
C526 VTAIL.n189 B 0.012817f
C527 VTAIL.n190 B 0.013571f
C528 VTAIL.n191 B 0.030296f
C529 VTAIL.n192 B 0.030296f
C530 VTAIL.n193 B 0.013571f
C531 VTAIL.n194 B 0.012817f
C532 VTAIL.n195 B 0.023853f
C533 VTAIL.n196 B 0.023853f
C534 VTAIL.n197 B 0.012817f
C535 VTAIL.n198 B 0.013571f
C536 VTAIL.n199 B 0.030296f
C537 VTAIL.n200 B 0.065016f
C538 VTAIL.n201 B 0.013571f
C539 VTAIL.n202 B 0.012817f
C540 VTAIL.n203 B 0.055786f
C541 VTAIL.n204 B 0.03634f
C542 VTAIL.n205 B 0.370911f
C543 VTAIL.t10 B 0.330614f
C544 VTAIL.t15 B 0.330614f
C545 VTAIL.n206 B 2.93648f
C546 VTAIL.n207 B 0.587809f
C547 VTAIL.t18 B 0.330614f
C548 VTAIL.t19 B 0.330614f
C549 VTAIL.n208 B 2.93648f
C550 VTAIL.n209 B 0.656386f
C551 VTAIL.n210 B 0.033205f
C552 VTAIL.n211 B 0.023853f
C553 VTAIL.n212 B 0.012817f
C554 VTAIL.n213 B 0.030296f
C555 VTAIL.n214 B 0.013571f
C556 VTAIL.n215 B 0.023853f
C557 VTAIL.n216 B 0.012817f
C558 VTAIL.n217 B 0.030296f
C559 VTAIL.n218 B 0.013194f
C560 VTAIL.n219 B 0.023853f
C561 VTAIL.n220 B 0.013194f
C562 VTAIL.n221 B 0.012817f
C563 VTAIL.n222 B 0.030296f
C564 VTAIL.n223 B 0.030296f
C565 VTAIL.n224 B 0.013571f
C566 VTAIL.n225 B 0.023853f
C567 VTAIL.n226 B 0.012817f
C568 VTAIL.n227 B 0.030296f
C569 VTAIL.n228 B 0.013571f
C570 VTAIL.n229 B 0.023853f
C571 VTAIL.n230 B 0.012817f
C572 VTAIL.n231 B 0.030296f
C573 VTAIL.n232 B 0.013571f
C574 VTAIL.n233 B 0.023853f
C575 VTAIL.n234 B 0.012817f
C576 VTAIL.n235 B 0.030296f
C577 VTAIL.n236 B 0.013571f
C578 VTAIL.n237 B 0.023853f
C579 VTAIL.n238 B 0.012817f
C580 VTAIL.n239 B 0.030296f
C581 VTAIL.n240 B 0.013571f
C582 VTAIL.n241 B 1.82956f
C583 VTAIL.n242 B 0.012817f
C584 VTAIL.t13 B 0.050162f
C585 VTAIL.n243 B 0.170763f
C586 VTAIL.n244 B 0.017897f
C587 VTAIL.n245 B 0.022722f
C588 VTAIL.n246 B 0.030296f
C589 VTAIL.n247 B 0.013571f
C590 VTAIL.n248 B 0.012817f
C591 VTAIL.n249 B 0.023853f
C592 VTAIL.n250 B 0.023853f
C593 VTAIL.n251 B 0.012817f
C594 VTAIL.n252 B 0.013571f
C595 VTAIL.n253 B 0.030296f
C596 VTAIL.n254 B 0.030296f
C597 VTAIL.n255 B 0.013571f
C598 VTAIL.n256 B 0.012817f
C599 VTAIL.n257 B 0.023853f
C600 VTAIL.n258 B 0.023853f
C601 VTAIL.n259 B 0.012817f
C602 VTAIL.n260 B 0.013571f
C603 VTAIL.n261 B 0.030296f
C604 VTAIL.n262 B 0.030296f
C605 VTAIL.n263 B 0.013571f
C606 VTAIL.n264 B 0.012817f
C607 VTAIL.n265 B 0.023853f
C608 VTAIL.n266 B 0.023853f
C609 VTAIL.n267 B 0.012817f
C610 VTAIL.n268 B 0.013571f
C611 VTAIL.n269 B 0.030296f
C612 VTAIL.n270 B 0.030296f
C613 VTAIL.n271 B 0.013571f
C614 VTAIL.n272 B 0.012817f
C615 VTAIL.n273 B 0.023853f
C616 VTAIL.n274 B 0.023853f
C617 VTAIL.n275 B 0.012817f
C618 VTAIL.n276 B 0.013571f
C619 VTAIL.n277 B 0.030296f
C620 VTAIL.n278 B 0.030296f
C621 VTAIL.n279 B 0.013571f
C622 VTAIL.n280 B 0.012817f
C623 VTAIL.n281 B 0.023853f
C624 VTAIL.n282 B 0.023853f
C625 VTAIL.n283 B 0.012817f
C626 VTAIL.n284 B 0.013571f
C627 VTAIL.n285 B 0.030296f
C628 VTAIL.n286 B 0.030296f
C629 VTAIL.n287 B 0.013571f
C630 VTAIL.n288 B 0.012817f
C631 VTAIL.n289 B 0.023853f
C632 VTAIL.n290 B 0.023853f
C633 VTAIL.n291 B 0.012817f
C634 VTAIL.n292 B 0.013571f
C635 VTAIL.n293 B 0.030296f
C636 VTAIL.n294 B 0.030296f
C637 VTAIL.n295 B 0.013571f
C638 VTAIL.n296 B 0.012817f
C639 VTAIL.n297 B 0.023853f
C640 VTAIL.n298 B 0.023853f
C641 VTAIL.n299 B 0.012817f
C642 VTAIL.n300 B 0.013571f
C643 VTAIL.n301 B 0.030296f
C644 VTAIL.n302 B 0.065016f
C645 VTAIL.n303 B 0.013571f
C646 VTAIL.n304 B 0.012817f
C647 VTAIL.n305 B 0.055786f
C648 VTAIL.n306 B 0.03634f
C649 VTAIL.n307 B 1.92566f
C650 VTAIL.n308 B 0.033205f
C651 VTAIL.n309 B 0.023853f
C652 VTAIL.n310 B 0.012817f
C653 VTAIL.n311 B 0.030296f
C654 VTAIL.n312 B 0.013571f
C655 VTAIL.n313 B 0.023853f
C656 VTAIL.n314 B 0.012817f
C657 VTAIL.n315 B 0.030296f
C658 VTAIL.n316 B 0.013194f
C659 VTAIL.n317 B 0.023853f
C660 VTAIL.n318 B 0.013571f
C661 VTAIL.n319 B 0.030296f
C662 VTAIL.n320 B 0.013571f
C663 VTAIL.n321 B 0.023853f
C664 VTAIL.n322 B 0.012817f
C665 VTAIL.n323 B 0.030296f
C666 VTAIL.n324 B 0.013571f
C667 VTAIL.n325 B 0.023853f
C668 VTAIL.n326 B 0.012817f
C669 VTAIL.n327 B 0.030296f
C670 VTAIL.n328 B 0.013571f
C671 VTAIL.n329 B 0.023853f
C672 VTAIL.n330 B 0.012817f
C673 VTAIL.n331 B 0.030296f
C674 VTAIL.n332 B 0.013571f
C675 VTAIL.n333 B 0.023853f
C676 VTAIL.n334 B 0.012817f
C677 VTAIL.n335 B 0.030296f
C678 VTAIL.n336 B 0.013571f
C679 VTAIL.n337 B 1.82956f
C680 VTAIL.n338 B 0.012817f
C681 VTAIL.t7 B 0.050162f
C682 VTAIL.n339 B 0.170763f
C683 VTAIL.n340 B 0.017897f
C684 VTAIL.n341 B 0.022722f
C685 VTAIL.n342 B 0.030296f
C686 VTAIL.n343 B 0.013571f
C687 VTAIL.n344 B 0.012817f
C688 VTAIL.n345 B 0.023853f
C689 VTAIL.n346 B 0.023853f
C690 VTAIL.n347 B 0.012817f
C691 VTAIL.n348 B 0.013571f
C692 VTAIL.n349 B 0.030296f
C693 VTAIL.n350 B 0.030296f
C694 VTAIL.n351 B 0.013571f
C695 VTAIL.n352 B 0.012817f
C696 VTAIL.n353 B 0.023853f
C697 VTAIL.n354 B 0.023853f
C698 VTAIL.n355 B 0.012817f
C699 VTAIL.n356 B 0.013571f
C700 VTAIL.n357 B 0.030296f
C701 VTAIL.n358 B 0.030296f
C702 VTAIL.n359 B 0.013571f
C703 VTAIL.n360 B 0.012817f
C704 VTAIL.n361 B 0.023853f
C705 VTAIL.n362 B 0.023853f
C706 VTAIL.n363 B 0.012817f
C707 VTAIL.n364 B 0.013571f
C708 VTAIL.n365 B 0.030296f
C709 VTAIL.n366 B 0.030296f
C710 VTAIL.n367 B 0.013571f
C711 VTAIL.n368 B 0.012817f
C712 VTAIL.n369 B 0.023853f
C713 VTAIL.n370 B 0.023853f
C714 VTAIL.n371 B 0.012817f
C715 VTAIL.n372 B 0.013571f
C716 VTAIL.n373 B 0.030296f
C717 VTAIL.n374 B 0.030296f
C718 VTAIL.n375 B 0.013571f
C719 VTAIL.n376 B 0.012817f
C720 VTAIL.n377 B 0.023853f
C721 VTAIL.n378 B 0.023853f
C722 VTAIL.n379 B 0.012817f
C723 VTAIL.n380 B 0.012817f
C724 VTAIL.n381 B 0.013571f
C725 VTAIL.n382 B 0.030296f
C726 VTAIL.n383 B 0.030296f
C727 VTAIL.n384 B 0.030296f
C728 VTAIL.n385 B 0.013194f
C729 VTAIL.n386 B 0.012817f
C730 VTAIL.n387 B 0.023853f
C731 VTAIL.n388 B 0.023853f
C732 VTAIL.n389 B 0.012817f
C733 VTAIL.n390 B 0.013571f
C734 VTAIL.n391 B 0.030296f
C735 VTAIL.n392 B 0.030296f
C736 VTAIL.n393 B 0.013571f
C737 VTAIL.n394 B 0.012817f
C738 VTAIL.n395 B 0.023853f
C739 VTAIL.n396 B 0.023853f
C740 VTAIL.n397 B 0.012817f
C741 VTAIL.n398 B 0.013571f
C742 VTAIL.n399 B 0.030296f
C743 VTAIL.n400 B 0.065016f
C744 VTAIL.n401 B 0.013571f
C745 VTAIL.n402 B 0.012817f
C746 VTAIL.n403 B 0.055786f
C747 VTAIL.n404 B 0.03634f
C748 VTAIL.n405 B 1.92566f
C749 VTAIL.t6 B 0.330614f
C750 VTAIL.t1 B 0.330614f
C751 VTAIL.n406 B 2.93646f
C752 VTAIL.n407 B 0.494896f
C753 VDD1.n0 B 0.033154f
C754 VDD1.n1 B 0.023816f
C755 VDD1.n2 B 0.012798f
C756 VDD1.n3 B 0.030249f
C757 VDD1.n4 B 0.01355f
C758 VDD1.n5 B 0.023816f
C759 VDD1.n6 B 0.012798f
C760 VDD1.n7 B 0.030249f
C761 VDD1.n8 B 0.013174f
C762 VDD1.n9 B 0.023816f
C763 VDD1.n10 B 0.013174f
C764 VDD1.n11 B 0.012798f
C765 VDD1.n12 B 0.030249f
C766 VDD1.n13 B 0.030249f
C767 VDD1.n14 B 0.01355f
C768 VDD1.n15 B 0.023816f
C769 VDD1.n16 B 0.012798f
C770 VDD1.n17 B 0.030249f
C771 VDD1.n18 B 0.01355f
C772 VDD1.n19 B 0.023816f
C773 VDD1.n20 B 0.012798f
C774 VDD1.n21 B 0.030249f
C775 VDD1.n22 B 0.01355f
C776 VDD1.n23 B 0.023816f
C777 VDD1.n24 B 0.012798f
C778 VDD1.n25 B 0.030249f
C779 VDD1.n26 B 0.01355f
C780 VDD1.n27 B 0.023816f
C781 VDD1.n28 B 0.012798f
C782 VDD1.n29 B 0.030249f
C783 VDD1.n30 B 0.01355f
C784 VDD1.n31 B 1.82672f
C785 VDD1.n32 B 0.012798f
C786 VDD1.t2 B 0.050084f
C787 VDD1.n33 B 0.170498f
C788 VDD1.n34 B 0.017869f
C789 VDD1.n35 B 0.022687f
C790 VDD1.n36 B 0.030249f
C791 VDD1.n37 B 0.01355f
C792 VDD1.n38 B 0.012798f
C793 VDD1.n39 B 0.023816f
C794 VDD1.n40 B 0.023816f
C795 VDD1.n41 B 0.012798f
C796 VDD1.n42 B 0.01355f
C797 VDD1.n43 B 0.030249f
C798 VDD1.n44 B 0.030249f
C799 VDD1.n45 B 0.01355f
C800 VDD1.n46 B 0.012798f
C801 VDD1.n47 B 0.023816f
C802 VDD1.n48 B 0.023816f
C803 VDD1.n49 B 0.012798f
C804 VDD1.n50 B 0.01355f
C805 VDD1.n51 B 0.030249f
C806 VDD1.n52 B 0.030249f
C807 VDD1.n53 B 0.01355f
C808 VDD1.n54 B 0.012798f
C809 VDD1.n55 B 0.023816f
C810 VDD1.n56 B 0.023816f
C811 VDD1.n57 B 0.012798f
C812 VDD1.n58 B 0.01355f
C813 VDD1.n59 B 0.030249f
C814 VDD1.n60 B 0.030249f
C815 VDD1.n61 B 0.01355f
C816 VDD1.n62 B 0.012798f
C817 VDD1.n63 B 0.023816f
C818 VDD1.n64 B 0.023816f
C819 VDD1.n65 B 0.012798f
C820 VDD1.n66 B 0.01355f
C821 VDD1.n67 B 0.030249f
C822 VDD1.n68 B 0.030249f
C823 VDD1.n69 B 0.01355f
C824 VDD1.n70 B 0.012798f
C825 VDD1.n71 B 0.023816f
C826 VDD1.n72 B 0.023816f
C827 VDD1.n73 B 0.012798f
C828 VDD1.n74 B 0.01355f
C829 VDD1.n75 B 0.030249f
C830 VDD1.n76 B 0.030249f
C831 VDD1.n77 B 0.01355f
C832 VDD1.n78 B 0.012798f
C833 VDD1.n79 B 0.023816f
C834 VDD1.n80 B 0.023816f
C835 VDD1.n81 B 0.012798f
C836 VDD1.n82 B 0.01355f
C837 VDD1.n83 B 0.030249f
C838 VDD1.n84 B 0.030249f
C839 VDD1.n85 B 0.01355f
C840 VDD1.n86 B 0.012798f
C841 VDD1.n87 B 0.023816f
C842 VDD1.n88 B 0.023816f
C843 VDD1.n89 B 0.012798f
C844 VDD1.n90 B 0.01355f
C845 VDD1.n91 B 0.030249f
C846 VDD1.n92 B 0.064915f
C847 VDD1.n93 B 0.01355f
C848 VDD1.n94 B 0.012798f
C849 VDD1.n95 B 0.0557f
C850 VDD1.n96 B 0.066103f
C851 VDD1.t7 B 0.330102f
C852 VDD1.t8 B 0.330102f
C853 VDD1.n97 B 3.00433f
C854 VDD1.n98 B 0.704915f
C855 VDD1.n99 B 0.033154f
C856 VDD1.n100 B 0.023816f
C857 VDD1.n101 B 0.012798f
C858 VDD1.n102 B 0.030249f
C859 VDD1.n103 B 0.01355f
C860 VDD1.n104 B 0.023816f
C861 VDD1.n105 B 0.012798f
C862 VDD1.n106 B 0.030249f
C863 VDD1.n107 B 0.013174f
C864 VDD1.n108 B 0.023816f
C865 VDD1.n109 B 0.01355f
C866 VDD1.n110 B 0.030249f
C867 VDD1.n111 B 0.01355f
C868 VDD1.n112 B 0.023816f
C869 VDD1.n113 B 0.012798f
C870 VDD1.n114 B 0.030249f
C871 VDD1.n115 B 0.01355f
C872 VDD1.n116 B 0.023816f
C873 VDD1.n117 B 0.012798f
C874 VDD1.n118 B 0.030249f
C875 VDD1.n119 B 0.01355f
C876 VDD1.n120 B 0.023816f
C877 VDD1.n121 B 0.012798f
C878 VDD1.n122 B 0.030249f
C879 VDD1.n123 B 0.01355f
C880 VDD1.n124 B 0.023816f
C881 VDD1.n125 B 0.012798f
C882 VDD1.n126 B 0.030249f
C883 VDD1.n127 B 0.01355f
C884 VDD1.n128 B 1.82672f
C885 VDD1.n129 B 0.012798f
C886 VDD1.t6 B 0.050084f
C887 VDD1.n130 B 0.170498f
C888 VDD1.n131 B 0.017869f
C889 VDD1.n132 B 0.022687f
C890 VDD1.n133 B 0.030249f
C891 VDD1.n134 B 0.01355f
C892 VDD1.n135 B 0.012798f
C893 VDD1.n136 B 0.023816f
C894 VDD1.n137 B 0.023816f
C895 VDD1.n138 B 0.012798f
C896 VDD1.n139 B 0.01355f
C897 VDD1.n140 B 0.030249f
C898 VDD1.n141 B 0.030249f
C899 VDD1.n142 B 0.01355f
C900 VDD1.n143 B 0.012798f
C901 VDD1.n144 B 0.023816f
C902 VDD1.n145 B 0.023816f
C903 VDD1.n146 B 0.012798f
C904 VDD1.n147 B 0.01355f
C905 VDD1.n148 B 0.030249f
C906 VDD1.n149 B 0.030249f
C907 VDD1.n150 B 0.01355f
C908 VDD1.n151 B 0.012798f
C909 VDD1.n152 B 0.023816f
C910 VDD1.n153 B 0.023816f
C911 VDD1.n154 B 0.012798f
C912 VDD1.n155 B 0.01355f
C913 VDD1.n156 B 0.030249f
C914 VDD1.n157 B 0.030249f
C915 VDD1.n158 B 0.01355f
C916 VDD1.n159 B 0.012798f
C917 VDD1.n160 B 0.023816f
C918 VDD1.n161 B 0.023816f
C919 VDD1.n162 B 0.012798f
C920 VDD1.n163 B 0.01355f
C921 VDD1.n164 B 0.030249f
C922 VDD1.n165 B 0.030249f
C923 VDD1.n166 B 0.01355f
C924 VDD1.n167 B 0.012798f
C925 VDD1.n168 B 0.023816f
C926 VDD1.n169 B 0.023816f
C927 VDD1.n170 B 0.012798f
C928 VDD1.n171 B 0.012798f
C929 VDD1.n172 B 0.01355f
C930 VDD1.n173 B 0.030249f
C931 VDD1.n174 B 0.030249f
C932 VDD1.n175 B 0.030249f
C933 VDD1.n176 B 0.013174f
C934 VDD1.n177 B 0.012798f
C935 VDD1.n178 B 0.023816f
C936 VDD1.n179 B 0.023816f
C937 VDD1.n180 B 0.012798f
C938 VDD1.n181 B 0.01355f
C939 VDD1.n182 B 0.030249f
C940 VDD1.n183 B 0.030249f
C941 VDD1.n184 B 0.01355f
C942 VDD1.n185 B 0.012798f
C943 VDD1.n186 B 0.023816f
C944 VDD1.n187 B 0.023816f
C945 VDD1.n188 B 0.012798f
C946 VDD1.n189 B 0.01355f
C947 VDD1.n190 B 0.030249f
C948 VDD1.n191 B 0.064915f
C949 VDD1.n192 B 0.01355f
C950 VDD1.n193 B 0.012798f
C951 VDD1.n194 B 0.0557f
C952 VDD1.n195 B 0.066103f
C953 VDD1.t3 B 0.330102f
C954 VDD1.t0 B 0.330102f
C955 VDD1.n196 B 3.00432f
C956 VDD1.n197 B 0.697094f
C957 VDD1.t4 B 0.330102f
C958 VDD1.t5 B 0.330102f
C959 VDD1.n198 B 3.02225f
C960 VDD1.n199 B 3.34194f
C961 VDD1.t9 B 0.330102f
C962 VDD1.t1 B 0.330102f
C963 VDD1.n200 B 3.00432f
C964 VDD1.n201 B 3.51381f
C965 VP.n0 B 0.025973f
C966 VP.t2 B 2.68859f
C967 VP.n1 B 0.039133f
C968 VP.n2 B 0.019701f
C969 VP.n3 B 0.021745f
C970 VP.n4 B 0.019701f
C971 VP.n5 B 0.033f
C972 VP.n6 B 0.019701f
C973 VP.t7 B 2.68859f
C974 VP.n7 B 0.036535f
C975 VP.n8 B 0.019701f
C976 VP.n9 B 0.033288f
C977 VP.n10 B 0.019701f
C978 VP.n11 B 0.015937f
C979 VP.n12 B 0.019701f
C980 VP.t5 B 2.68859f
C981 VP.n13 B 0.996189f
C982 VP.n14 B 0.025973f
C983 VP.t6 B 2.68859f
C984 VP.n15 B 0.039133f
C985 VP.n16 B 0.019701f
C986 VP.n17 B 0.021745f
C987 VP.n18 B 0.019701f
C988 VP.n19 B 0.033f
C989 VP.n20 B 0.019701f
C990 VP.t1 B 2.68859f
C991 VP.n21 B 0.036535f
C992 VP.n22 B 0.019701f
C993 VP.n23 B 0.033288f
C994 VP.t9 B 2.88324f
C995 VP.t4 B 2.68859f
C996 VP.n24 B 0.99803f
C997 VP.n25 B 0.962975f
C998 VP.n26 B 0.207406f
C999 VP.n27 B 0.019701f
C1000 VP.n28 B 0.036535f
C1001 VP.n29 B 0.024279f
C1002 VP.n30 B 0.033f
C1003 VP.n31 B 0.019701f
C1004 VP.n32 B 0.019701f
C1005 VP.n33 B 0.019701f
C1006 VP.n34 B 0.027517f
C1007 VP.n35 B 0.931593f
C1008 VP.n36 B 0.027517f
C1009 VP.n37 B 0.036535f
C1010 VP.n38 B 0.019701f
C1011 VP.n39 B 0.019701f
C1012 VP.n40 B 0.019701f
C1013 VP.n41 B 0.024279f
C1014 VP.n42 B 0.036535f
C1015 VP.t0 B 2.68859f
C1016 VP.n43 B 0.931593f
C1017 VP.n44 B 0.033288f
C1018 VP.n45 B 0.019701f
C1019 VP.n46 B 0.019701f
C1020 VP.n47 B 0.019701f
C1021 VP.n48 B 0.036535f
C1022 VP.n49 B 0.038743f
C1023 VP.n50 B 0.015937f
C1024 VP.n51 B 0.019701f
C1025 VP.n52 B 0.019701f
C1026 VP.n53 B 0.019701f
C1027 VP.n54 B 0.036535f
C1028 VP.n55 B 0.021024f
C1029 VP.n56 B 0.996189f
C1030 VP.n57 B 1.3757f
C1031 VP.n58 B 1.38784f
C1032 VP.n59 B 0.025973f
C1033 VP.n60 B 0.021024f
C1034 VP.n61 B 0.036535f
C1035 VP.n62 B 0.039133f
C1036 VP.n63 B 0.019701f
C1037 VP.n64 B 0.019701f
C1038 VP.n65 B 0.019701f
C1039 VP.n66 B 0.038743f
C1040 VP.n67 B 0.036535f
C1041 VP.t8 B 2.68859f
C1042 VP.n68 B 0.931593f
C1043 VP.n69 B 0.021745f
C1044 VP.n70 B 0.019701f
C1045 VP.n71 B 0.019701f
C1046 VP.n72 B 0.019701f
C1047 VP.n73 B 0.036535f
C1048 VP.n74 B 0.024279f
C1049 VP.n75 B 0.033f
C1050 VP.n76 B 0.019701f
C1051 VP.n77 B 0.019701f
C1052 VP.n78 B 0.019701f
C1053 VP.n79 B 0.027517f
C1054 VP.n80 B 0.931593f
C1055 VP.n81 B 0.027517f
C1056 VP.n82 B 0.036535f
C1057 VP.n83 B 0.019701f
C1058 VP.n84 B 0.019701f
C1059 VP.n85 B 0.019701f
C1060 VP.n86 B 0.024279f
C1061 VP.n87 B 0.036535f
C1062 VP.t3 B 2.68859f
C1063 VP.n88 B 0.931593f
C1064 VP.n89 B 0.033288f
C1065 VP.n90 B 0.019701f
C1066 VP.n91 B 0.019701f
C1067 VP.n92 B 0.019701f
C1068 VP.n93 B 0.036535f
C1069 VP.n94 B 0.038743f
C1070 VP.n95 B 0.015937f
C1071 VP.n96 B 0.019701f
C1072 VP.n97 B 0.019701f
C1073 VP.n98 B 0.019701f
C1074 VP.n99 B 0.036535f
C1075 VP.n100 B 0.021024f
C1076 VP.n101 B 0.996189f
C1077 VP.n102 B 0.036726f
.ends

