* NGSPICE file created from diff_pair_sample_1707.ext - technology: sky130A

.subckt diff_pair_sample_1707 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VN.t0 VDD2.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=2.09715 pd=13.04 as=2.09715 ps=13.04 w=12.71 l=3.95
X1 VTAIL.t14 VN.t1 VDD2.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=2.09715 pd=13.04 as=2.09715 ps=13.04 w=12.71 l=3.95
X2 VTAIL.t0 VP.t0 VDD1.t7 B.t0 sky130_fd_pr__nfet_01v8 ad=2.09715 pd=13.04 as=2.09715 ps=13.04 w=12.71 l=3.95
X3 VTAIL.t2 VP.t1 VDD1.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=2.09715 pd=13.04 as=2.09715 ps=13.04 w=12.71 l=3.95
X4 B.t21 B.t19 B.t20 B.t16 sky130_fd_pr__nfet_01v8 ad=4.9569 pd=26.2 as=0 ps=0 w=12.71 l=3.95
X5 VTAIL.t13 VN.t2 VDD2.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=4.9569 pd=26.2 as=2.09715 ps=13.04 w=12.71 l=3.95
X6 VDD1.t5 VP.t2 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=2.09715 pd=13.04 as=4.9569 ps=26.2 w=12.71 l=3.95
X7 VDD2.t2 VN.t3 VTAIL.t12 B.t6 sky130_fd_pr__nfet_01v8 ad=2.09715 pd=13.04 as=4.9569 ps=26.2 w=12.71 l=3.95
X8 VDD1.t4 VP.t3 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.09715 pd=13.04 as=2.09715 ps=13.04 w=12.71 l=3.95
X9 B.t18 B.t15 B.t17 B.t16 sky130_fd_pr__nfet_01v8 ad=4.9569 pd=26.2 as=0 ps=0 w=12.71 l=3.95
X10 VTAIL.t7 VP.t4 VDD1.t3 B.t7 sky130_fd_pr__nfet_01v8 ad=4.9569 pd=26.2 as=2.09715 ps=13.04 w=12.71 l=3.95
X11 VTAIL.t3 VP.t5 VDD1.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=4.9569 pd=26.2 as=2.09715 ps=13.04 w=12.71 l=3.95
X12 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=4.9569 pd=26.2 as=0 ps=0 w=12.71 l=3.95
X13 VTAIL.t11 VN.t4 VDD2.t1 B.t7 sky130_fd_pr__nfet_01v8 ad=4.9569 pd=26.2 as=2.09715 ps=13.04 w=12.71 l=3.95
X14 VDD2.t0 VN.t5 VTAIL.t10 B.t4 sky130_fd_pr__nfet_01v8 ad=2.09715 pd=13.04 as=4.9569 ps=26.2 w=12.71 l=3.95
X15 VDD1.t1 VP.t6 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.09715 pd=13.04 as=2.09715 ps=13.04 w=12.71 l=3.95
X16 VDD2.t7 VN.t6 VTAIL.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=2.09715 pd=13.04 as=2.09715 ps=13.04 w=12.71 l=3.95
X17 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=4.9569 pd=26.2 as=0 ps=0 w=12.71 l=3.95
X18 VDD1.t0 VP.t7 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=2.09715 pd=13.04 as=4.9569 ps=26.2 w=12.71 l=3.95
X19 VDD2.t6 VN.t7 VTAIL.t8 B.t1 sky130_fd_pr__nfet_01v8 ad=2.09715 pd=13.04 as=2.09715 ps=13.04 w=12.71 l=3.95
R0 VN.n75 VN.n39 161.3
R1 VN.n74 VN.n73 161.3
R2 VN.n72 VN.n40 161.3
R3 VN.n71 VN.n70 161.3
R4 VN.n69 VN.n41 161.3
R5 VN.n68 VN.n67 161.3
R6 VN.n66 VN.n42 161.3
R7 VN.n65 VN.n64 161.3
R8 VN.n62 VN.n43 161.3
R9 VN.n61 VN.n60 161.3
R10 VN.n59 VN.n44 161.3
R11 VN.n58 VN.n57 161.3
R12 VN.n56 VN.n45 161.3
R13 VN.n55 VN.n54 161.3
R14 VN.n53 VN.n46 161.3
R15 VN.n52 VN.n51 161.3
R16 VN.n50 VN.n47 161.3
R17 VN.n36 VN.n0 161.3
R18 VN.n35 VN.n34 161.3
R19 VN.n33 VN.n1 161.3
R20 VN.n32 VN.n31 161.3
R21 VN.n30 VN.n2 161.3
R22 VN.n29 VN.n28 161.3
R23 VN.n27 VN.n3 161.3
R24 VN.n26 VN.n25 161.3
R25 VN.n23 VN.n4 161.3
R26 VN.n22 VN.n21 161.3
R27 VN.n20 VN.n5 161.3
R28 VN.n19 VN.n18 161.3
R29 VN.n17 VN.n6 161.3
R30 VN.n16 VN.n15 161.3
R31 VN.n14 VN.n7 161.3
R32 VN.n13 VN.n12 161.3
R33 VN.n11 VN.n8 161.3
R34 VN.n9 VN.t4 109.796
R35 VN.n48 VN.t5 109.796
R36 VN.n10 VN.t7 77.5476
R37 VN.n24 VN.t1 77.5476
R38 VN.n37 VN.t3 77.5476
R39 VN.n49 VN.t0 77.5476
R40 VN.n63 VN.t6 77.5476
R41 VN.n76 VN.t2 77.5476
R42 VN.n10 VN.n9 68.2271
R43 VN.n49 VN.n48 68.2271
R44 VN.n38 VN.n37 61.6295
R45 VN.n77 VN.n76 61.6295
R46 VN VN.n77 58.0269
R47 VN.n31 VN.n30 56.5193
R48 VN.n70 VN.n69 56.5193
R49 VN.n17 VN.n16 40.4934
R50 VN.n18 VN.n17 40.4934
R51 VN.n56 VN.n55 40.4934
R52 VN.n57 VN.n56 40.4934
R53 VN.n12 VN.n11 24.4675
R54 VN.n12 VN.n7 24.4675
R55 VN.n16 VN.n7 24.4675
R56 VN.n18 VN.n5 24.4675
R57 VN.n22 VN.n5 24.4675
R58 VN.n23 VN.n22 24.4675
R59 VN.n25 VN.n3 24.4675
R60 VN.n29 VN.n3 24.4675
R61 VN.n30 VN.n29 24.4675
R62 VN.n31 VN.n1 24.4675
R63 VN.n35 VN.n1 24.4675
R64 VN.n36 VN.n35 24.4675
R65 VN.n55 VN.n46 24.4675
R66 VN.n51 VN.n46 24.4675
R67 VN.n51 VN.n50 24.4675
R68 VN.n69 VN.n68 24.4675
R69 VN.n68 VN.n42 24.4675
R70 VN.n64 VN.n42 24.4675
R71 VN.n62 VN.n61 24.4675
R72 VN.n61 VN.n44 24.4675
R73 VN.n57 VN.n44 24.4675
R74 VN.n75 VN.n74 24.4675
R75 VN.n74 VN.n40 24.4675
R76 VN.n70 VN.n40 24.4675
R77 VN.n37 VN.n36 20.5528
R78 VN.n76 VN.n75 20.5528
R79 VN.n25 VN.n24 17.6167
R80 VN.n64 VN.n63 17.6167
R81 VN.n11 VN.n10 6.85126
R82 VN.n24 VN.n23 6.85126
R83 VN.n50 VN.n49 6.85126
R84 VN.n63 VN.n62 6.85126
R85 VN.n48 VN.n47 2.67497
R86 VN.n9 VN.n8 2.67497
R87 VN.n77 VN.n39 0.417535
R88 VN.n38 VN.n0 0.417535
R89 VN VN.n38 0.394291
R90 VN.n73 VN.n39 0.189894
R91 VN.n73 VN.n72 0.189894
R92 VN.n72 VN.n71 0.189894
R93 VN.n71 VN.n41 0.189894
R94 VN.n67 VN.n41 0.189894
R95 VN.n67 VN.n66 0.189894
R96 VN.n66 VN.n65 0.189894
R97 VN.n65 VN.n43 0.189894
R98 VN.n60 VN.n43 0.189894
R99 VN.n60 VN.n59 0.189894
R100 VN.n59 VN.n58 0.189894
R101 VN.n58 VN.n45 0.189894
R102 VN.n54 VN.n45 0.189894
R103 VN.n54 VN.n53 0.189894
R104 VN.n53 VN.n52 0.189894
R105 VN.n52 VN.n47 0.189894
R106 VN.n13 VN.n8 0.189894
R107 VN.n14 VN.n13 0.189894
R108 VN.n15 VN.n14 0.189894
R109 VN.n15 VN.n6 0.189894
R110 VN.n19 VN.n6 0.189894
R111 VN.n20 VN.n19 0.189894
R112 VN.n21 VN.n20 0.189894
R113 VN.n21 VN.n4 0.189894
R114 VN.n26 VN.n4 0.189894
R115 VN.n27 VN.n26 0.189894
R116 VN.n28 VN.n27 0.189894
R117 VN.n28 VN.n2 0.189894
R118 VN.n32 VN.n2 0.189894
R119 VN.n33 VN.n32 0.189894
R120 VN.n34 VN.n33 0.189894
R121 VN.n34 VN.n0 0.189894
R122 VDD2.n2 VDD2.n1 67.4575
R123 VDD2.n2 VDD2.n0 67.4575
R124 VDD2 VDD2.n5 67.4547
R125 VDD2.n4 VDD2.n3 65.669
R126 VDD2.n4 VDD2.n2 51.2756
R127 VDD2 VDD2.n4 1.90352
R128 VDD2.n5 VDD2.t5 1.55833
R129 VDD2.n5 VDD2.t0 1.55833
R130 VDD2.n3 VDD2.t3 1.55833
R131 VDD2.n3 VDD2.t7 1.55833
R132 VDD2.n1 VDD2.t4 1.55833
R133 VDD2.n1 VDD2.t2 1.55833
R134 VDD2.n0 VDD2.t1 1.55833
R135 VDD2.n0 VDD2.t6 1.55833
R136 VTAIL.n566 VTAIL.n565 289.615
R137 VTAIL.n70 VTAIL.n69 289.615
R138 VTAIL.n140 VTAIL.n139 289.615
R139 VTAIL.n212 VTAIL.n211 289.615
R140 VTAIL.n496 VTAIL.n495 289.615
R141 VTAIL.n424 VTAIL.n423 289.615
R142 VTAIL.n354 VTAIL.n353 289.615
R143 VTAIL.n282 VTAIL.n281 289.615
R144 VTAIL.n520 VTAIL.n519 185
R145 VTAIL.n525 VTAIL.n524 185
R146 VTAIL.n527 VTAIL.n526 185
R147 VTAIL.n516 VTAIL.n515 185
R148 VTAIL.n533 VTAIL.n532 185
R149 VTAIL.n535 VTAIL.n534 185
R150 VTAIL.n512 VTAIL.n511 185
R151 VTAIL.n541 VTAIL.n540 185
R152 VTAIL.n543 VTAIL.n542 185
R153 VTAIL.n508 VTAIL.n507 185
R154 VTAIL.n549 VTAIL.n548 185
R155 VTAIL.n551 VTAIL.n550 185
R156 VTAIL.n504 VTAIL.n503 185
R157 VTAIL.n557 VTAIL.n556 185
R158 VTAIL.n559 VTAIL.n558 185
R159 VTAIL.n500 VTAIL.n499 185
R160 VTAIL.n565 VTAIL.n564 185
R161 VTAIL.n24 VTAIL.n23 185
R162 VTAIL.n29 VTAIL.n28 185
R163 VTAIL.n31 VTAIL.n30 185
R164 VTAIL.n20 VTAIL.n19 185
R165 VTAIL.n37 VTAIL.n36 185
R166 VTAIL.n39 VTAIL.n38 185
R167 VTAIL.n16 VTAIL.n15 185
R168 VTAIL.n45 VTAIL.n44 185
R169 VTAIL.n47 VTAIL.n46 185
R170 VTAIL.n12 VTAIL.n11 185
R171 VTAIL.n53 VTAIL.n52 185
R172 VTAIL.n55 VTAIL.n54 185
R173 VTAIL.n8 VTAIL.n7 185
R174 VTAIL.n61 VTAIL.n60 185
R175 VTAIL.n63 VTAIL.n62 185
R176 VTAIL.n4 VTAIL.n3 185
R177 VTAIL.n69 VTAIL.n68 185
R178 VTAIL.n94 VTAIL.n93 185
R179 VTAIL.n99 VTAIL.n98 185
R180 VTAIL.n101 VTAIL.n100 185
R181 VTAIL.n90 VTAIL.n89 185
R182 VTAIL.n107 VTAIL.n106 185
R183 VTAIL.n109 VTAIL.n108 185
R184 VTAIL.n86 VTAIL.n85 185
R185 VTAIL.n115 VTAIL.n114 185
R186 VTAIL.n117 VTAIL.n116 185
R187 VTAIL.n82 VTAIL.n81 185
R188 VTAIL.n123 VTAIL.n122 185
R189 VTAIL.n125 VTAIL.n124 185
R190 VTAIL.n78 VTAIL.n77 185
R191 VTAIL.n131 VTAIL.n130 185
R192 VTAIL.n133 VTAIL.n132 185
R193 VTAIL.n74 VTAIL.n73 185
R194 VTAIL.n139 VTAIL.n138 185
R195 VTAIL.n166 VTAIL.n165 185
R196 VTAIL.n171 VTAIL.n170 185
R197 VTAIL.n173 VTAIL.n172 185
R198 VTAIL.n162 VTAIL.n161 185
R199 VTAIL.n179 VTAIL.n178 185
R200 VTAIL.n181 VTAIL.n180 185
R201 VTAIL.n158 VTAIL.n157 185
R202 VTAIL.n187 VTAIL.n186 185
R203 VTAIL.n189 VTAIL.n188 185
R204 VTAIL.n154 VTAIL.n153 185
R205 VTAIL.n195 VTAIL.n194 185
R206 VTAIL.n197 VTAIL.n196 185
R207 VTAIL.n150 VTAIL.n149 185
R208 VTAIL.n203 VTAIL.n202 185
R209 VTAIL.n205 VTAIL.n204 185
R210 VTAIL.n146 VTAIL.n145 185
R211 VTAIL.n211 VTAIL.n210 185
R212 VTAIL.n495 VTAIL.n494 185
R213 VTAIL.n430 VTAIL.n429 185
R214 VTAIL.n489 VTAIL.n488 185
R215 VTAIL.n487 VTAIL.n486 185
R216 VTAIL.n434 VTAIL.n433 185
R217 VTAIL.n481 VTAIL.n480 185
R218 VTAIL.n479 VTAIL.n478 185
R219 VTAIL.n438 VTAIL.n437 185
R220 VTAIL.n473 VTAIL.n472 185
R221 VTAIL.n471 VTAIL.n470 185
R222 VTAIL.n442 VTAIL.n441 185
R223 VTAIL.n465 VTAIL.n464 185
R224 VTAIL.n463 VTAIL.n462 185
R225 VTAIL.n446 VTAIL.n445 185
R226 VTAIL.n457 VTAIL.n456 185
R227 VTAIL.n455 VTAIL.n454 185
R228 VTAIL.n450 VTAIL.n449 185
R229 VTAIL.n423 VTAIL.n422 185
R230 VTAIL.n358 VTAIL.n357 185
R231 VTAIL.n417 VTAIL.n416 185
R232 VTAIL.n415 VTAIL.n414 185
R233 VTAIL.n362 VTAIL.n361 185
R234 VTAIL.n409 VTAIL.n408 185
R235 VTAIL.n407 VTAIL.n406 185
R236 VTAIL.n366 VTAIL.n365 185
R237 VTAIL.n401 VTAIL.n400 185
R238 VTAIL.n399 VTAIL.n398 185
R239 VTAIL.n370 VTAIL.n369 185
R240 VTAIL.n393 VTAIL.n392 185
R241 VTAIL.n391 VTAIL.n390 185
R242 VTAIL.n374 VTAIL.n373 185
R243 VTAIL.n385 VTAIL.n384 185
R244 VTAIL.n383 VTAIL.n382 185
R245 VTAIL.n378 VTAIL.n377 185
R246 VTAIL.n353 VTAIL.n352 185
R247 VTAIL.n288 VTAIL.n287 185
R248 VTAIL.n347 VTAIL.n346 185
R249 VTAIL.n345 VTAIL.n344 185
R250 VTAIL.n292 VTAIL.n291 185
R251 VTAIL.n339 VTAIL.n338 185
R252 VTAIL.n337 VTAIL.n336 185
R253 VTAIL.n296 VTAIL.n295 185
R254 VTAIL.n331 VTAIL.n330 185
R255 VTAIL.n329 VTAIL.n328 185
R256 VTAIL.n300 VTAIL.n299 185
R257 VTAIL.n323 VTAIL.n322 185
R258 VTAIL.n321 VTAIL.n320 185
R259 VTAIL.n304 VTAIL.n303 185
R260 VTAIL.n315 VTAIL.n314 185
R261 VTAIL.n313 VTAIL.n312 185
R262 VTAIL.n308 VTAIL.n307 185
R263 VTAIL.n281 VTAIL.n280 185
R264 VTAIL.n216 VTAIL.n215 185
R265 VTAIL.n275 VTAIL.n274 185
R266 VTAIL.n273 VTAIL.n272 185
R267 VTAIL.n220 VTAIL.n219 185
R268 VTAIL.n267 VTAIL.n266 185
R269 VTAIL.n265 VTAIL.n264 185
R270 VTAIL.n224 VTAIL.n223 185
R271 VTAIL.n259 VTAIL.n258 185
R272 VTAIL.n257 VTAIL.n256 185
R273 VTAIL.n228 VTAIL.n227 185
R274 VTAIL.n251 VTAIL.n250 185
R275 VTAIL.n249 VTAIL.n248 185
R276 VTAIL.n232 VTAIL.n231 185
R277 VTAIL.n243 VTAIL.n242 185
R278 VTAIL.n241 VTAIL.n240 185
R279 VTAIL.n236 VTAIL.n235 185
R280 VTAIL.n521 VTAIL.t12 147.659
R281 VTAIL.n25 VTAIL.t11 147.659
R282 VTAIL.n95 VTAIL.t4 147.659
R283 VTAIL.n167 VTAIL.t3 147.659
R284 VTAIL.n451 VTAIL.t6 147.659
R285 VTAIL.n379 VTAIL.t7 147.659
R286 VTAIL.n309 VTAIL.t10 147.659
R287 VTAIL.n237 VTAIL.t13 147.659
R288 VTAIL.n525 VTAIL.n519 104.615
R289 VTAIL.n526 VTAIL.n525 104.615
R290 VTAIL.n526 VTAIL.n515 104.615
R291 VTAIL.n533 VTAIL.n515 104.615
R292 VTAIL.n534 VTAIL.n533 104.615
R293 VTAIL.n534 VTAIL.n511 104.615
R294 VTAIL.n541 VTAIL.n511 104.615
R295 VTAIL.n542 VTAIL.n541 104.615
R296 VTAIL.n542 VTAIL.n507 104.615
R297 VTAIL.n549 VTAIL.n507 104.615
R298 VTAIL.n550 VTAIL.n549 104.615
R299 VTAIL.n550 VTAIL.n503 104.615
R300 VTAIL.n557 VTAIL.n503 104.615
R301 VTAIL.n558 VTAIL.n557 104.615
R302 VTAIL.n558 VTAIL.n499 104.615
R303 VTAIL.n565 VTAIL.n499 104.615
R304 VTAIL.n29 VTAIL.n23 104.615
R305 VTAIL.n30 VTAIL.n29 104.615
R306 VTAIL.n30 VTAIL.n19 104.615
R307 VTAIL.n37 VTAIL.n19 104.615
R308 VTAIL.n38 VTAIL.n37 104.615
R309 VTAIL.n38 VTAIL.n15 104.615
R310 VTAIL.n45 VTAIL.n15 104.615
R311 VTAIL.n46 VTAIL.n45 104.615
R312 VTAIL.n46 VTAIL.n11 104.615
R313 VTAIL.n53 VTAIL.n11 104.615
R314 VTAIL.n54 VTAIL.n53 104.615
R315 VTAIL.n54 VTAIL.n7 104.615
R316 VTAIL.n61 VTAIL.n7 104.615
R317 VTAIL.n62 VTAIL.n61 104.615
R318 VTAIL.n62 VTAIL.n3 104.615
R319 VTAIL.n69 VTAIL.n3 104.615
R320 VTAIL.n99 VTAIL.n93 104.615
R321 VTAIL.n100 VTAIL.n99 104.615
R322 VTAIL.n100 VTAIL.n89 104.615
R323 VTAIL.n107 VTAIL.n89 104.615
R324 VTAIL.n108 VTAIL.n107 104.615
R325 VTAIL.n108 VTAIL.n85 104.615
R326 VTAIL.n115 VTAIL.n85 104.615
R327 VTAIL.n116 VTAIL.n115 104.615
R328 VTAIL.n116 VTAIL.n81 104.615
R329 VTAIL.n123 VTAIL.n81 104.615
R330 VTAIL.n124 VTAIL.n123 104.615
R331 VTAIL.n124 VTAIL.n77 104.615
R332 VTAIL.n131 VTAIL.n77 104.615
R333 VTAIL.n132 VTAIL.n131 104.615
R334 VTAIL.n132 VTAIL.n73 104.615
R335 VTAIL.n139 VTAIL.n73 104.615
R336 VTAIL.n171 VTAIL.n165 104.615
R337 VTAIL.n172 VTAIL.n171 104.615
R338 VTAIL.n172 VTAIL.n161 104.615
R339 VTAIL.n179 VTAIL.n161 104.615
R340 VTAIL.n180 VTAIL.n179 104.615
R341 VTAIL.n180 VTAIL.n157 104.615
R342 VTAIL.n187 VTAIL.n157 104.615
R343 VTAIL.n188 VTAIL.n187 104.615
R344 VTAIL.n188 VTAIL.n153 104.615
R345 VTAIL.n195 VTAIL.n153 104.615
R346 VTAIL.n196 VTAIL.n195 104.615
R347 VTAIL.n196 VTAIL.n149 104.615
R348 VTAIL.n203 VTAIL.n149 104.615
R349 VTAIL.n204 VTAIL.n203 104.615
R350 VTAIL.n204 VTAIL.n145 104.615
R351 VTAIL.n211 VTAIL.n145 104.615
R352 VTAIL.n495 VTAIL.n429 104.615
R353 VTAIL.n488 VTAIL.n429 104.615
R354 VTAIL.n488 VTAIL.n487 104.615
R355 VTAIL.n487 VTAIL.n433 104.615
R356 VTAIL.n480 VTAIL.n433 104.615
R357 VTAIL.n480 VTAIL.n479 104.615
R358 VTAIL.n479 VTAIL.n437 104.615
R359 VTAIL.n472 VTAIL.n437 104.615
R360 VTAIL.n472 VTAIL.n471 104.615
R361 VTAIL.n471 VTAIL.n441 104.615
R362 VTAIL.n464 VTAIL.n441 104.615
R363 VTAIL.n464 VTAIL.n463 104.615
R364 VTAIL.n463 VTAIL.n445 104.615
R365 VTAIL.n456 VTAIL.n445 104.615
R366 VTAIL.n456 VTAIL.n455 104.615
R367 VTAIL.n455 VTAIL.n449 104.615
R368 VTAIL.n423 VTAIL.n357 104.615
R369 VTAIL.n416 VTAIL.n357 104.615
R370 VTAIL.n416 VTAIL.n415 104.615
R371 VTAIL.n415 VTAIL.n361 104.615
R372 VTAIL.n408 VTAIL.n361 104.615
R373 VTAIL.n408 VTAIL.n407 104.615
R374 VTAIL.n407 VTAIL.n365 104.615
R375 VTAIL.n400 VTAIL.n365 104.615
R376 VTAIL.n400 VTAIL.n399 104.615
R377 VTAIL.n399 VTAIL.n369 104.615
R378 VTAIL.n392 VTAIL.n369 104.615
R379 VTAIL.n392 VTAIL.n391 104.615
R380 VTAIL.n391 VTAIL.n373 104.615
R381 VTAIL.n384 VTAIL.n373 104.615
R382 VTAIL.n384 VTAIL.n383 104.615
R383 VTAIL.n383 VTAIL.n377 104.615
R384 VTAIL.n353 VTAIL.n287 104.615
R385 VTAIL.n346 VTAIL.n287 104.615
R386 VTAIL.n346 VTAIL.n345 104.615
R387 VTAIL.n345 VTAIL.n291 104.615
R388 VTAIL.n338 VTAIL.n291 104.615
R389 VTAIL.n338 VTAIL.n337 104.615
R390 VTAIL.n337 VTAIL.n295 104.615
R391 VTAIL.n330 VTAIL.n295 104.615
R392 VTAIL.n330 VTAIL.n329 104.615
R393 VTAIL.n329 VTAIL.n299 104.615
R394 VTAIL.n322 VTAIL.n299 104.615
R395 VTAIL.n322 VTAIL.n321 104.615
R396 VTAIL.n321 VTAIL.n303 104.615
R397 VTAIL.n314 VTAIL.n303 104.615
R398 VTAIL.n314 VTAIL.n313 104.615
R399 VTAIL.n313 VTAIL.n307 104.615
R400 VTAIL.n281 VTAIL.n215 104.615
R401 VTAIL.n274 VTAIL.n215 104.615
R402 VTAIL.n274 VTAIL.n273 104.615
R403 VTAIL.n273 VTAIL.n219 104.615
R404 VTAIL.n266 VTAIL.n219 104.615
R405 VTAIL.n266 VTAIL.n265 104.615
R406 VTAIL.n265 VTAIL.n223 104.615
R407 VTAIL.n258 VTAIL.n223 104.615
R408 VTAIL.n258 VTAIL.n257 104.615
R409 VTAIL.n257 VTAIL.n227 104.615
R410 VTAIL.n250 VTAIL.n227 104.615
R411 VTAIL.n250 VTAIL.n249 104.615
R412 VTAIL.n249 VTAIL.n231 104.615
R413 VTAIL.n242 VTAIL.n231 104.615
R414 VTAIL.n242 VTAIL.n241 104.615
R415 VTAIL.n241 VTAIL.n235 104.615
R416 VTAIL.t12 VTAIL.n519 52.3082
R417 VTAIL.t11 VTAIL.n23 52.3082
R418 VTAIL.t4 VTAIL.n93 52.3082
R419 VTAIL.t3 VTAIL.n165 52.3082
R420 VTAIL.t6 VTAIL.n449 52.3082
R421 VTAIL.t7 VTAIL.n377 52.3082
R422 VTAIL.t10 VTAIL.n307 52.3082
R423 VTAIL.t13 VTAIL.n235 52.3082
R424 VTAIL.n427 VTAIL.n426 48.9902
R425 VTAIL.n285 VTAIL.n284 48.9902
R426 VTAIL.n1 VTAIL.n0 48.9893
R427 VTAIL.n143 VTAIL.n142 48.9893
R428 VTAIL.n567 VTAIL.n566 36.2581
R429 VTAIL.n71 VTAIL.n70 36.2581
R430 VTAIL.n141 VTAIL.n140 36.2581
R431 VTAIL.n213 VTAIL.n212 36.2581
R432 VTAIL.n497 VTAIL.n496 36.2581
R433 VTAIL.n425 VTAIL.n424 36.2581
R434 VTAIL.n355 VTAIL.n354 36.2581
R435 VTAIL.n283 VTAIL.n282 36.2581
R436 VTAIL.n567 VTAIL.n497 27.0134
R437 VTAIL.n283 VTAIL.n213 27.0134
R438 VTAIL.n521 VTAIL.n520 15.6677
R439 VTAIL.n25 VTAIL.n24 15.6677
R440 VTAIL.n95 VTAIL.n94 15.6677
R441 VTAIL.n167 VTAIL.n166 15.6677
R442 VTAIL.n451 VTAIL.n450 15.6677
R443 VTAIL.n379 VTAIL.n378 15.6677
R444 VTAIL.n309 VTAIL.n308 15.6677
R445 VTAIL.n237 VTAIL.n236 15.6677
R446 VTAIL.n524 VTAIL.n523 12.8005
R447 VTAIL.n564 VTAIL.n498 12.8005
R448 VTAIL.n28 VTAIL.n27 12.8005
R449 VTAIL.n68 VTAIL.n2 12.8005
R450 VTAIL.n98 VTAIL.n97 12.8005
R451 VTAIL.n138 VTAIL.n72 12.8005
R452 VTAIL.n170 VTAIL.n169 12.8005
R453 VTAIL.n210 VTAIL.n144 12.8005
R454 VTAIL.n494 VTAIL.n428 12.8005
R455 VTAIL.n454 VTAIL.n453 12.8005
R456 VTAIL.n422 VTAIL.n356 12.8005
R457 VTAIL.n382 VTAIL.n381 12.8005
R458 VTAIL.n352 VTAIL.n286 12.8005
R459 VTAIL.n312 VTAIL.n311 12.8005
R460 VTAIL.n280 VTAIL.n214 12.8005
R461 VTAIL.n240 VTAIL.n239 12.8005
R462 VTAIL.n527 VTAIL.n518 12.0247
R463 VTAIL.n563 VTAIL.n500 12.0247
R464 VTAIL.n31 VTAIL.n22 12.0247
R465 VTAIL.n67 VTAIL.n4 12.0247
R466 VTAIL.n101 VTAIL.n92 12.0247
R467 VTAIL.n137 VTAIL.n74 12.0247
R468 VTAIL.n173 VTAIL.n164 12.0247
R469 VTAIL.n209 VTAIL.n146 12.0247
R470 VTAIL.n493 VTAIL.n430 12.0247
R471 VTAIL.n457 VTAIL.n448 12.0247
R472 VTAIL.n421 VTAIL.n358 12.0247
R473 VTAIL.n385 VTAIL.n376 12.0247
R474 VTAIL.n351 VTAIL.n288 12.0247
R475 VTAIL.n315 VTAIL.n306 12.0247
R476 VTAIL.n279 VTAIL.n216 12.0247
R477 VTAIL.n243 VTAIL.n234 12.0247
R478 VTAIL.n528 VTAIL.n516 11.249
R479 VTAIL.n560 VTAIL.n559 11.249
R480 VTAIL.n32 VTAIL.n20 11.249
R481 VTAIL.n64 VTAIL.n63 11.249
R482 VTAIL.n102 VTAIL.n90 11.249
R483 VTAIL.n134 VTAIL.n133 11.249
R484 VTAIL.n174 VTAIL.n162 11.249
R485 VTAIL.n206 VTAIL.n205 11.249
R486 VTAIL.n490 VTAIL.n489 11.249
R487 VTAIL.n458 VTAIL.n446 11.249
R488 VTAIL.n418 VTAIL.n417 11.249
R489 VTAIL.n386 VTAIL.n374 11.249
R490 VTAIL.n348 VTAIL.n347 11.249
R491 VTAIL.n316 VTAIL.n304 11.249
R492 VTAIL.n276 VTAIL.n275 11.249
R493 VTAIL.n244 VTAIL.n232 11.249
R494 VTAIL.n532 VTAIL.n531 10.4732
R495 VTAIL.n556 VTAIL.n502 10.4732
R496 VTAIL.n36 VTAIL.n35 10.4732
R497 VTAIL.n60 VTAIL.n6 10.4732
R498 VTAIL.n106 VTAIL.n105 10.4732
R499 VTAIL.n130 VTAIL.n76 10.4732
R500 VTAIL.n178 VTAIL.n177 10.4732
R501 VTAIL.n202 VTAIL.n148 10.4732
R502 VTAIL.n486 VTAIL.n432 10.4732
R503 VTAIL.n462 VTAIL.n461 10.4732
R504 VTAIL.n414 VTAIL.n360 10.4732
R505 VTAIL.n390 VTAIL.n389 10.4732
R506 VTAIL.n344 VTAIL.n290 10.4732
R507 VTAIL.n320 VTAIL.n319 10.4732
R508 VTAIL.n272 VTAIL.n218 10.4732
R509 VTAIL.n248 VTAIL.n247 10.4732
R510 VTAIL.n535 VTAIL.n514 9.69747
R511 VTAIL.n555 VTAIL.n504 9.69747
R512 VTAIL.n39 VTAIL.n18 9.69747
R513 VTAIL.n59 VTAIL.n8 9.69747
R514 VTAIL.n109 VTAIL.n88 9.69747
R515 VTAIL.n129 VTAIL.n78 9.69747
R516 VTAIL.n181 VTAIL.n160 9.69747
R517 VTAIL.n201 VTAIL.n150 9.69747
R518 VTAIL.n485 VTAIL.n434 9.69747
R519 VTAIL.n465 VTAIL.n444 9.69747
R520 VTAIL.n413 VTAIL.n362 9.69747
R521 VTAIL.n393 VTAIL.n372 9.69747
R522 VTAIL.n343 VTAIL.n292 9.69747
R523 VTAIL.n323 VTAIL.n302 9.69747
R524 VTAIL.n271 VTAIL.n220 9.69747
R525 VTAIL.n251 VTAIL.n230 9.69747
R526 VTAIL.n562 VTAIL.n498 9.45567
R527 VTAIL.n66 VTAIL.n2 9.45567
R528 VTAIL.n136 VTAIL.n72 9.45567
R529 VTAIL.n208 VTAIL.n144 9.45567
R530 VTAIL.n492 VTAIL.n428 9.45567
R531 VTAIL.n420 VTAIL.n356 9.45567
R532 VTAIL.n350 VTAIL.n286 9.45567
R533 VTAIL.n278 VTAIL.n214 9.45567
R534 VTAIL.n545 VTAIL.n544 9.3005
R535 VTAIL.n547 VTAIL.n546 9.3005
R536 VTAIL.n506 VTAIL.n505 9.3005
R537 VTAIL.n553 VTAIL.n552 9.3005
R538 VTAIL.n555 VTAIL.n554 9.3005
R539 VTAIL.n502 VTAIL.n501 9.3005
R540 VTAIL.n561 VTAIL.n560 9.3005
R541 VTAIL.n563 VTAIL.n562 9.3005
R542 VTAIL.n539 VTAIL.n538 9.3005
R543 VTAIL.n537 VTAIL.n536 9.3005
R544 VTAIL.n514 VTAIL.n513 9.3005
R545 VTAIL.n531 VTAIL.n530 9.3005
R546 VTAIL.n529 VTAIL.n528 9.3005
R547 VTAIL.n518 VTAIL.n517 9.3005
R548 VTAIL.n523 VTAIL.n522 9.3005
R549 VTAIL.n510 VTAIL.n509 9.3005
R550 VTAIL.n49 VTAIL.n48 9.3005
R551 VTAIL.n51 VTAIL.n50 9.3005
R552 VTAIL.n10 VTAIL.n9 9.3005
R553 VTAIL.n57 VTAIL.n56 9.3005
R554 VTAIL.n59 VTAIL.n58 9.3005
R555 VTAIL.n6 VTAIL.n5 9.3005
R556 VTAIL.n65 VTAIL.n64 9.3005
R557 VTAIL.n67 VTAIL.n66 9.3005
R558 VTAIL.n43 VTAIL.n42 9.3005
R559 VTAIL.n41 VTAIL.n40 9.3005
R560 VTAIL.n18 VTAIL.n17 9.3005
R561 VTAIL.n35 VTAIL.n34 9.3005
R562 VTAIL.n33 VTAIL.n32 9.3005
R563 VTAIL.n22 VTAIL.n21 9.3005
R564 VTAIL.n27 VTAIL.n26 9.3005
R565 VTAIL.n14 VTAIL.n13 9.3005
R566 VTAIL.n119 VTAIL.n118 9.3005
R567 VTAIL.n121 VTAIL.n120 9.3005
R568 VTAIL.n80 VTAIL.n79 9.3005
R569 VTAIL.n127 VTAIL.n126 9.3005
R570 VTAIL.n129 VTAIL.n128 9.3005
R571 VTAIL.n76 VTAIL.n75 9.3005
R572 VTAIL.n135 VTAIL.n134 9.3005
R573 VTAIL.n137 VTAIL.n136 9.3005
R574 VTAIL.n113 VTAIL.n112 9.3005
R575 VTAIL.n111 VTAIL.n110 9.3005
R576 VTAIL.n88 VTAIL.n87 9.3005
R577 VTAIL.n105 VTAIL.n104 9.3005
R578 VTAIL.n103 VTAIL.n102 9.3005
R579 VTAIL.n92 VTAIL.n91 9.3005
R580 VTAIL.n97 VTAIL.n96 9.3005
R581 VTAIL.n84 VTAIL.n83 9.3005
R582 VTAIL.n191 VTAIL.n190 9.3005
R583 VTAIL.n193 VTAIL.n192 9.3005
R584 VTAIL.n152 VTAIL.n151 9.3005
R585 VTAIL.n199 VTAIL.n198 9.3005
R586 VTAIL.n201 VTAIL.n200 9.3005
R587 VTAIL.n148 VTAIL.n147 9.3005
R588 VTAIL.n207 VTAIL.n206 9.3005
R589 VTAIL.n209 VTAIL.n208 9.3005
R590 VTAIL.n185 VTAIL.n184 9.3005
R591 VTAIL.n183 VTAIL.n182 9.3005
R592 VTAIL.n160 VTAIL.n159 9.3005
R593 VTAIL.n177 VTAIL.n176 9.3005
R594 VTAIL.n175 VTAIL.n174 9.3005
R595 VTAIL.n164 VTAIL.n163 9.3005
R596 VTAIL.n169 VTAIL.n168 9.3005
R597 VTAIL.n156 VTAIL.n155 9.3005
R598 VTAIL.n493 VTAIL.n492 9.3005
R599 VTAIL.n491 VTAIL.n490 9.3005
R600 VTAIL.n432 VTAIL.n431 9.3005
R601 VTAIL.n485 VTAIL.n484 9.3005
R602 VTAIL.n483 VTAIL.n482 9.3005
R603 VTAIL.n436 VTAIL.n435 9.3005
R604 VTAIL.n477 VTAIL.n476 9.3005
R605 VTAIL.n475 VTAIL.n474 9.3005
R606 VTAIL.n440 VTAIL.n439 9.3005
R607 VTAIL.n469 VTAIL.n468 9.3005
R608 VTAIL.n467 VTAIL.n466 9.3005
R609 VTAIL.n444 VTAIL.n443 9.3005
R610 VTAIL.n461 VTAIL.n460 9.3005
R611 VTAIL.n459 VTAIL.n458 9.3005
R612 VTAIL.n448 VTAIL.n447 9.3005
R613 VTAIL.n453 VTAIL.n452 9.3005
R614 VTAIL.n405 VTAIL.n404 9.3005
R615 VTAIL.n364 VTAIL.n363 9.3005
R616 VTAIL.n411 VTAIL.n410 9.3005
R617 VTAIL.n413 VTAIL.n412 9.3005
R618 VTAIL.n360 VTAIL.n359 9.3005
R619 VTAIL.n419 VTAIL.n418 9.3005
R620 VTAIL.n421 VTAIL.n420 9.3005
R621 VTAIL.n403 VTAIL.n402 9.3005
R622 VTAIL.n368 VTAIL.n367 9.3005
R623 VTAIL.n397 VTAIL.n396 9.3005
R624 VTAIL.n395 VTAIL.n394 9.3005
R625 VTAIL.n372 VTAIL.n371 9.3005
R626 VTAIL.n389 VTAIL.n388 9.3005
R627 VTAIL.n387 VTAIL.n386 9.3005
R628 VTAIL.n376 VTAIL.n375 9.3005
R629 VTAIL.n381 VTAIL.n380 9.3005
R630 VTAIL.n335 VTAIL.n334 9.3005
R631 VTAIL.n294 VTAIL.n293 9.3005
R632 VTAIL.n341 VTAIL.n340 9.3005
R633 VTAIL.n343 VTAIL.n342 9.3005
R634 VTAIL.n290 VTAIL.n289 9.3005
R635 VTAIL.n349 VTAIL.n348 9.3005
R636 VTAIL.n351 VTAIL.n350 9.3005
R637 VTAIL.n333 VTAIL.n332 9.3005
R638 VTAIL.n298 VTAIL.n297 9.3005
R639 VTAIL.n327 VTAIL.n326 9.3005
R640 VTAIL.n325 VTAIL.n324 9.3005
R641 VTAIL.n302 VTAIL.n301 9.3005
R642 VTAIL.n319 VTAIL.n318 9.3005
R643 VTAIL.n317 VTAIL.n316 9.3005
R644 VTAIL.n306 VTAIL.n305 9.3005
R645 VTAIL.n311 VTAIL.n310 9.3005
R646 VTAIL.n263 VTAIL.n262 9.3005
R647 VTAIL.n222 VTAIL.n221 9.3005
R648 VTAIL.n269 VTAIL.n268 9.3005
R649 VTAIL.n271 VTAIL.n270 9.3005
R650 VTAIL.n218 VTAIL.n217 9.3005
R651 VTAIL.n277 VTAIL.n276 9.3005
R652 VTAIL.n279 VTAIL.n278 9.3005
R653 VTAIL.n261 VTAIL.n260 9.3005
R654 VTAIL.n226 VTAIL.n225 9.3005
R655 VTAIL.n255 VTAIL.n254 9.3005
R656 VTAIL.n253 VTAIL.n252 9.3005
R657 VTAIL.n230 VTAIL.n229 9.3005
R658 VTAIL.n247 VTAIL.n246 9.3005
R659 VTAIL.n245 VTAIL.n244 9.3005
R660 VTAIL.n234 VTAIL.n233 9.3005
R661 VTAIL.n239 VTAIL.n238 9.3005
R662 VTAIL.n536 VTAIL.n512 8.92171
R663 VTAIL.n552 VTAIL.n551 8.92171
R664 VTAIL.n40 VTAIL.n16 8.92171
R665 VTAIL.n56 VTAIL.n55 8.92171
R666 VTAIL.n110 VTAIL.n86 8.92171
R667 VTAIL.n126 VTAIL.n125 8.92171
R668 VTAIL.n182 VTAIL.n158 8.92171
R669 VTAIL.n198 VTAIL.n197 8.92171
R670 VTAIL.n482 VTAIL.n481 8.92171
R671 VTAIL.n466 VTAIL.n442 8.92171
R672 VTAIL.n410 VTAIL.n409 8.92171
R673 VTAIL.n394 VTAIL.n370 8.92171
R674 VTAIL.n340 VTAIL.n339 8.92171
R675 VTAIL.n324 VTAIL.n300 8.92171
R676 VTAIL.n268 VTAIL.n267 8.92171
R677 VTAIL.n252 VTAIL.n228 8.92171
R678 VTAIL.n540 VTAIL.n539 8.14595
R679 VTAIL.n548 VTAIL.n506 8.14595
R680 VTAIL.n44 VTAIL.n43 8.14595
R681 VTAIL.n52 VTAIL.n10 8.14595
R682 VTAIL.n114 VTAIL.n113 8.14595
R683 VTAIL.n122 VTAIL.n80 8.14595
R684 VTAIL.n186 VTAIL.n185 8.14595
R685 VTAIL.n194 VTAIL.n152 8.14595
R686 VTAIL.n478 VTAIL.n436 8.14595
R687 VTAIL.n470 VTAIL.n469 8.14595
R688 VTAIL.n406 VTAIL.n364 8.14595
R689 VTAIL.n398 VTAIL.n397 8.14595
R690 VTAIL.n336 VTAIL.n294 8.14595
R691 VTAIL.n328 VTAIL.n327 8.14595
R692 VTAIL.n264 VTAIL.n222 8.14595
R693 VTAIL.n256 VTAIL.n255 8.14595
R694 VTAIL.n543 VTAIL.n510 7.3702
R695 VTAIL.n547 VTAIL.n508 7.3702
R696 VTAIL.n47 VTAIL.n14 7.3702
R697 VTAIL.n51 VTAIL.n12 7.3702
R698 VTAIL.n117 VTAIL.n84 7.3702
R699 VTAIL.n121 VTAIL.n82 7.3702
R700 VTAIL.n189 VTAIL.n156 7.3702
R701 VTAIL.n193 VTAIL.n154 7.3702
R702 VTAIL.n477 VTAIL.n438 7.3702
R703 VTAIL.n473 VTAIL.n440 7.3702
R704 VTAIL.n405 VTAIL.n366 7.3702
R705 VTAIL.n401 VTAIL.n368 7.3702
R706 VTAIL.n335 VTAIL.n296 7.3702
R707 VTAIL.n331 VTAIL.n298 7.3702
R708 VTAIL.n263 VTAIL.n224 7.3702
R709 VTAIL.n259 VTAIL.n226 7.3702
R710 VTAIL.n544 VTAIL.n543 6.59444
R711 VTAIL.n544 VTAIL.n508 6.59444
R712 VTAIL.n48 VTAIL.n47 6.59444
R713 VTAIL.n48 VTAIL.n12 6.59444
R714 VTAIL.n118 VTAIL.n117 6.59444
R715 VTAIL.n118 VTAIL.n82 6.59444
R716 VTAIL.n190 VTAIL.n189 6.59444
R717 VTAIL.n190 VTAIL.n154 6.59444
R718 VTAIL.n474 VTAIL.n438 6.59444
R719 VTAIL.n474 VTAIL.n473 6.59444
R720 VTAIL.n402 VTAIL.n366 6.59444
R721 VTAIL.n402 VTAIL.n401 6.59444
R722 VTAIL.n332 VTAIL.n296 6.59444
R723 VTAIL.n332 VTAIL.n331 6.59444
R724 VTAIL.n260 VTAIL.n224 6.59444
R725 VTAIL.n260 VTAIL.n259 6.59444
R726 VTAIL.n540 VTAIL.n510 5.81868
R727 VTAIL.n548 VTAIL.n547 5.81868
R728 VTAIL.n44 VTAIL.n14 5.81868
R729 VTAIL.n52 VTAIL.n51 5.81868
R730 VTAIL.n114 VTAIL.n84 5.81868
R731 VTAIL.n122 VTAIL.n121 5.81868
R732 VTAIL.n186 VTAIL.n156 5.81868
R733 VTAIL.n194 VTAIL.n193 5.81868
R734 VTAIL.n478 VTAIL.n477 5.81868
R735 VTAIL.n470 VTAIL.n440 5.81868
R736 VTAIL.n406 VTAIL.n405 5.81868
R737 VTAIL.n398 VTAIL.n368 5.81868
R738 VTAIL.n336 VTAIL.n335 5.81868
R739 VTAIL.n328 VTAIL.n298 5.81868
R740 VTAIL.n264 VTAIL.n263 5.81868
R741 VTAIL.n256 VTAIL.n226 5.81868
R742 VTAIL.n539 VTAIL.n512 5.04292
R743 VTAIL.n551 VTAIL.n506 5.04292
R744 VTAIL.n43 VTAIL.n16 5.04292
R745 VTAIL.n55 VTAIL.n10 5.04292
R746 VTAIL.n113 VTAIL.n86 5.04292
R747 VTAIL.n125 VTAIL.n80 5.04292
R748 VTAIL.n185 VTAIL.n158 5.04292
R749 VTAIL.n197 VTAIL.n152 5.04292
R750 VTAIL.n481 VTAIL.n436 5.04292
R751 VTAIL.n469 VTAIL.n442 5.04292
R752 VTAIL.n409 VTAIL.n364 5.04292
R753 VTAIL.n397 VTAIL.n370 5.04292
R754 VTAIL.n339 VTAIL.n294 5.04292
R755 VTAIL.n327 VTAIL.n300 5.04292
R756 VTAIL.n267 VTAIL.n222 5.04292
R757 VTAIL.n255 VTAIL.n228 5.04292
R758 VTAIL.n522 VTAIL.n521 4.38563
R759 VTAIL.n26 VTAIL.n25 4.38563
R760 VTAIL.n96 VTAIL.n95 4.38563
R761 VTAIL.n168 VTAIL.n167 4.38563
R762 VTAIL.n452 VTAIL.n451 4.38563
R763 VTAIL.n380 VTAIL.n379 4.38563
R764 VTAIL.n310 VTAIL.n309 4.38563
R765 VTAIL.n238 VTAIL.n237 4.38563
R766 VTAIL.n536 VTAIL.n535 4.26717
R767 VTAIL.n552 VTAIL.n504 4.26717
R768 VTAIL.n40 VTAIL.n39 4.26717
R769 VTAIL.n56 VTAIL.n8 4.26717
R770 VTAIL.n110 VTAIL.n109 4.26717
R771 VTAIL.n126 VTAIL.n78 4.26717
R772 VTAIL.n182 VTAIL.n181 4.26717
R773 VTAIL.n198 VTAIL.n150 4.26717
R774 VTAIL.n482 VTAIL.n434 4.26717
R775 VTAIL.n466 VTAIL.n465 4.26717
R776 VTAIL.n410 VTAIL.n362 4.26717
R777 VTAIL.n394 VTAIL.n393 4.26717
R778 VTAIL.n340 VTAIL.n292 4.26717
R779 VTAIL.n324 VTAIL.n323 4.26717
R780 VTAIL.n268 VTAIL.n220 4.26717
R781 VTAIL.n252 VTAIL.n251 4.26717
R782 VTAIL.n285 VTAIL.n283 3.69016
R783 VTAIL.n355 VTAIL.n285 3.69016
R784 VTAIL.n427 VTAIL.n425 3.69016
R785 VTAIL.n497 VTAIL.n427 3.69016
R786 VTAIL.n213 VTAIL.n143 3.69016
R787 VTAIL.n143 VTAIL.n141 3.69016
R788 VTAIL.n71 VTAIL.n1 3.69016
R789 VTAIL VTAIL.n567 3.63197
R790 VTAIL.n532 VTAIL.n514 3.49141
R791 VTAIL.n556 VTAIL.n555 3.49141
R792 VTAIL.n36 VTAIL.n18 3.49141
R793 VTAIL.n60 VTAIL.n59 3.49141
R794 VTAIL.n106 VTAIL.n88 3.49141
R795 VTAIL.n130 VTAIL.n129 3.49141
R796 VTAIL.n178 VTAIL.n160 3.49141
R797 VTAIL.n202 VTAIL.n201 3.49141
R798 VTAIL.n486 VTAIL.n485 3.49141
R799 VTAIL.n462 VTAIL.n444 3.49141
R800 VTAIL.n414 VTAIL.n413 3.49141
R801 VTAIL.n390 VTAIL.n372 3.49141
R802 VTAIL.n344 VTAIL.n343 3.49141
R803 VTAIL.n320 VTAIL.n302 3.49141
R804 VTAIL.n272 VTAIL.n271 3.49141
R805 VTAIL.n248 VTAIL.n230 3.49141
R806 VTAIL.n531 VTAIL.n516 2.71565
R807 VTAIL.n559 VTAIL.n502 2.71565
R808 VTAIL.n35 VTAIL.n20 2.71565
R809 VTAIL.n63 VTAIL.n6 2.71565
R810 VTAIL.n105 VTAIL.n90 2.71565
R811 VTAIL.n133 VTAIL.n76 2.71565
R812 VTAIL.n177 VTAIL.n162 2.71565
R813 VTAIL.n205 VTAIL.n148 2.71565
R814 VTAIL.n489 VTAIL.n432 2.71565
R815 VTAIL.n461 VTAIL.n446 2.71565
R816 VTAIL.n417 VTAIL.n360 2.71565
R817 VTAIL.n389 VTAIL.n374 2.71565
R818 VTAIL.n347 VTAIL.n290 2.71565
R819 VTAIL.n319 VTAIL.n304 2.71565
R820 VTAIL.n275 VTAIL.n218 2.71565
R821 VTAIL.n247 VTAIL.n232 2.71565
R822 VTAIL.n528 VTAIL.n527 1.93989
R823 VTAIL.n560 VTAIL.n500 1.93989
R824 VTAIL.n32 VTAIL.n31 1.93989
R825 VTAIL.n64 VTAIL.n4 1.93989
R826 VTAIL.n102 VTAIL.n101 1.93989
R827 VTAIL.n134 VTAIL.n74 1.93989
R828 VTAIL.n174 VTAIL.n173 1.93989
R829 VTAIL.n206 VTAIL.n146 1.93989
R830 VTAIL.n490 VTAIL.n430 1.93989
R831 VTAIL.n458 VTAIL.n457 1.93989
R832 VTAIL.n418 VTAIL.n358 1.93989
R833 VTAIL.n386 VTAIL.n385 1.93989
R834 VTAIL.n348 VTAIL.n288 1.93989
R835 VTAIL.n316 VTAIL.n315 1.93989
R836 VTAIL.n276 VTAIL.n216 1.93989
R837 VTAIL.n244 VTAIL.n243 1.93989
R838 VTAIL.n0 VTAIL.t8 1.55833
R839 VTAIL.n0 VTAIL.t14 1.55833
R840 VTAIL.n142 VTAIL.t5 1.55833
R841 VTAIL.n142 VTAIL.t0 1.55833
R842 VTAIL.n426 VTAIL.t1 1.55833
R843 VTAIL.n426 VTAIL.t2 1.55833
R844 VTAIL.n284 VTAIL.t9 1.55833
R845 VTAIL.n284 VTAIL.t15 1.55833
R846 VTAIL.n524 VTAIL.n518 1.16414
R847 VTAIL.n564 VTAIL.n563 1.16414
R848 VTAIL.n28 VTAIL.n22 1.16414
R849 VTAIL.n68 VTAIL.n67 1.16414
R850 VTAIL.n98 VTAIL.n92 1.16414
R851 VTAIL.n138 VTAIL.n137 1.16414
R852 VTAIL.n170 VTAIL.n164 1.16414
R853 VTAIL.n210 VTAIL.n209 1.16414
R854 VTAIL.n494 VTAIL.n493 1.16414
R855 VTAIL.n454 VTAIL.n448 1.16414
R856 VTAIL.n422 VTAIL.n421 1.16414
R857 VTAIL.n382 VTAIL.n376 1.16414
R858 VTAIL.n352 VTAIL.n351 1.16414
R859 VTAIL.n312 VTAIL.n306 1.16414
R860 VTAIL.n280 VTAIL.n279 1.16414
R861 VTAIL.n240 VTAIL.n234 1.16414
R862 VTAIL.n425 VTAIL.n355 0.470328
R863 VTAIL.n141 VTAIL.n71 0.470328
R864 VTAIL.n523 VTAIL.n520 0.388379
R865 VTAIL.n566 VTAIL.n498 0.388379
R866 VTAIL.n27 VTAIL.n24 0.388379
R867 VTAIL.n70 VTAIL.n2 0.388379
R868 VTAIL.n97 VTAIL.n94 0.388379
R869 VTAIL.n140 VTAIL.n72 0.388379
R870 VTAIL.n169 VTAIL.n166 0.388379
R871 VTAIL.n212 VTAIL.n144 0.388379
R872 VTAIL.n496 VTAIL.n428 0.388379
R873 VTAIL.n453 VTAIL.n450 0.388379
R874 VTAIL.n424 VTAIL.n356 0.388379
R875 VTAIL.n381 VTAIL.n378 0.388379
R876 VTAIL.n354 VTAIL.n286 0.388379
R877 VTAIL.n311 VTAIL.n308 0.388379
R878 VTAIL.n282 VTAIL.n214 0.388379
R879 VTAIL.n239 VTAIL.n236 0.388379
R880 VTAIL.n522 VTAIL.n517 0.155672
R881 VTAIL.n529 VTAIL.n517 0.155672
R882 VTAIL.n530 VTAIL.n529 0.155672
R883 VTAIL.n530 VTAIL.n513 0.155672
R884 VTAIL.n537 VTAIL.n513 0.155672
R885 VTAIL.n538 VTAIL.n537 0.155672
R886 VTAIL.n538 VTAIL.n509 0.155672
R887 VTAIL.n545 VTAIL.n509 0.155672
R888 VTAIL.n546 VTAIL.n545 0.155672
R889 VTAIL.n546 VTAIL.n505 0.155672
R890 VTAIL.n553 VTAIL.n505 0.155672
R891 VTAIL.n554 VTAIL.n553 0.155672
R892 VTAIL.n554 VTAIL.n501 0.155672
R893 VTAIL.n561 VTAIL.n501 0.155672
R894 VTAIL.n562 VTAIL.n561 0.155672
R895 VTAIL.n26 VTAIL.n21 0.155672
R896 VTAIL.n33 VTAIL.n21 0.155672
R897 VTAIL.n34 VTAIL.n33 0.155672
R898 VTAIL.n34 VTAIL.n17 0.155672
R899 VTAIL.n41 VTAIL.n17 0.155672
R900 VTAIL.n42 VTAIL.n41 0.155672
R901 VTAIL.n42 VTAIL.n13 0.155672
R902 VTAIL.n49 VTAIL.n13 0.155672
R903 VTAIL.n50 VTAIL.n49 0.155672
R904 VTAIL.n50 VTAIL.n9 0.155672
R905 VTAIL.n57 VTAIL.n9 0.155672
R906 VTAIL.n58 VTAIL.n57 0.155672
R907 VTAIL.n58 VTAIL.n5 0.155672
R908 VTAIL.n65 VTAIL.n5 0.155672
R909 VTAIL.n66 VTAIL.n65 0.155672
R910 VTAIL.n96 VTAIL.n91 0.155672
R911 VTAIL.n103 VTAIL.n91 0.155672
R912 VTAIL.n104 VTAIL.n103 0.155672
R913 VTAIL.n104 VTAIL.n87 0.155672
R914 VTAIL.n111 VTAIL.n87 0.155672
R915 VTAIL.n112 VTAIL.n111 0.155672
R916 VTAIL.n112 VTAIL.n83 0.155672
R917 VTAIL.n119 VTAIL.n83 0.155672
R918 VTAIL.n120 VTAIL.n119 0.155672
R919 VTAIL.n120 VTAIL.n79 0.155672
R920 VTAIL.n127 VTAIL.n79 0.155672
R921 VTAIL.n128 VTAIL.n127 0.155672
R922 VTAIL.n128 VTAIL.n75 0.155672
R923 VTAIL.n135 VTAIL.n75 0.155672
R924 VTAIL.n136 VTAIL.n135 0.155672
R925 VTAIL.n168 VTAIL.n163 0.155672
R926 VTAIL.n175 VTAIL.n163 0.155672
R927 VTAIL.n176 VTAIL.n175 0.155672
R928 VTAIL.n176 VTAIL.n159 0.155672
R929 VTAIL.n183 VTAIL.n159 0.155672
R930 VTAIL.n184 VTAIL.n183 0.155672
R931 VTAIL.n184 VTAIL.n155 0.155672
R932 VTAIL.n191 VTAIL.n155 0.155672
R933 VTAIL.n192 VTAIL.n191 0.155672
R934 VTAIL.n192 VTAIL.n151 0.155672
R935 VTAIL.n199 VTAIL.n151 0.155672
R936 VTAIL.n200 VTAIL.n199 0.155672
R937 VTAIL.n200 VTAIL.n147 0.155672
R938 VTAIL.n207 VTAIL.n147 0.155672
R939 VTAIL.n208 VTAIL.n207 0.155672
R940 VTAIL.n492 VTAIL.n491 0.155672
R941 VTAIL.n491 VTAIL.n431 0.155672
R942 VTAIL.n484 VTAIL.n431 0.155672
R943 VTAIL.n484 VTAIL.n483 0.155672
R944 VTAIL.n483 VTAIL.n435 0.155672
R945 VTAIL.n476 VTAIL.n435 0.155672
R946 VTAIL.n476 VTAIL.n475 0.155672
R947 VTAIL.n475 VTAIL.n439 0.155672
R948 VTAIL.n468 VTAIL.n439 0.155672
R949 VTAIL.n468 VTAIL.n467 0.155672
R950 VTAIL.n467 VTAIL.n443 0.155672
R951 VTAIL.n460 VTAIL.n443 0.155672
R952 VTAIL.n460 VTAIL.n459 0.155672
R953 VTAIL.n459 VTAIL.n447 0.155672
R954 VTAIL.n452 VTAIL.n447 0.155672
R955 VTAIL.n420 VTAIL.n419 0.155672
R956 VTAIL.n419 VTAIL.n359 0.155672
R957 VTAIL.n412 VTAIL.n359 0.155672
R958 VTAIL.n412 VTAIL.n411 0.155672
R959 VTAIL.n411 VTAIL.n363 0.155672
R960 VTAIL.n404 VTAIL.n363 0.155672
R961 VTAIL.n404 VTAIL.n403 0.155672
R962 VTAIL.n403 VTAIL.n367 0.155672
R963 VTAIL.n396 VTAIL.n367 0.155672
R964 VTAIL.n396 VTAIL.n395 0.155672
R965 VTAIL.n395 VTAIL.n371 0.155672
R966 VTAIL.n388 VTAIL.n371 0.155672
R967 VTAIL.n388 VTAIL.n387 0.155672
R968 VTAIL.n387 VTAIL.n375 0.155672
R969 VTAIL.n380 VTAIL.n375 0.155672
R970 VTAIL.n350 VTAIL.n349 0.155672
R971 VTAIL.n349 VTAIL.n289 0.155672
R972 VTAIL.n342 VTAIL.n289 0.155672
R973 VTAIL.n342 VTAIL.n341 0.155672
R974 VTAIL.n341 VTAIL.n293 0.155672
R975 VTAIL.n334 VTAIL.n293 0.155672
R976 VTAIL.n334 VTAIL.n333 0.155672
R977 VTAIL.n333 VTAIL.n297 0.155672
R978 VTAIL.n326 VTAIL.n297 0.155672
R979 VTAIL.n326 VTAIL.n325 0.155672
R980 VTAIL.n325 VTAIL.n301 0.155672
R981 VTAIL.n318 VTAIL.n301 0.155672
R982 VTAIL.n318 VTAIL.n317 0.155672
R983 VTAIL.n317 VTAIL.n305 0.155672
R984 VTAIL.n310 VTAIL.n305 0.155672
R985 VTAIL.n278 VTAIL.n277 0.155672
R986 VTAIL.n277 VTAIL.n217 0.155672
R987 VTAIL.n270 VTAIL.n217 0.155672
R988 VTAIL.n270 VTAIL.n269 0.155672
R989 VTAIL.n269 VTAIL.n221 0.155672
R990 VTAIL.n262 VTAIL.n221 0.155672
R991 VTAIL.n262 VTAIL.n261 0.155672
R992 VTAIL.n261 VTAIL.n225 0.155672
R993 VTAIL.n254 VTAIL.n225 0.155672
R994 VTAIL.n254 VTAIL.n253 0.155672
R995 VTAIL.n253 VTAIL.n229 0.155672
R996 VTAIL.n246 VTAIL.n229 0.155672
R997 VTAIL.n246 VTAIL.n245 0.155672
R998 VTAIL.n245 VTAIL.n233 0.155672
R999 VTAIL.n238 VTAIL.n233 0.155672
R1000 VTAIL VTAIL.n1 0.0586897
R1001 B.n1064 B.n1063 585
R1002 B.n1065 B.n1064 585
R1003 B.n372 B.n178 585
R1004 B.n371 B.n370 585
R1005 B.n369 B.n368 585
R1006 B.n367 B.n366 585
R1007 B.n365 B.n364 585
R1008 B.n363 B.n362 585
R1009 B.n361 B.n360 585
R1010 B.n359 B.n358 585
R1011 B.n357 B.n356 585
R1012 B.n355 B.n354 585
R1013 B.n353 B.n352 585
R1014 B.n351 B.n350 585
R1015 B.n349 B.n348 585
R1016 B.n347 B.n346 585
R1017 B.n345 B.n344 585
R1018 B.n343 B.n342 585
R1019 B.n341 B.n340 585
R1020 B.n339 B.n338 585
R1021 B.n337 B.n336 585
R1022 B.n335 B.n334 585
R1023 B.n333 B.n332 585
R1024 B.n331 B.n330 585
R1025 B.n329 B.n328 585
R1026 B.n327 B.n326 585
R1027 B.n325 B.n324 585
R1028 B.n323 B.n322 585
R1029 B.n321 B.n320 585
R1030 B.n319 B.n318 585
R1031 B.n317 B.n316 585
R1032 B.n315 B.n314 585
R1033 B.n313 B.n312 585
R1034 B.n311 B.n310 585
R1035 B.n309 B.n308 585
R1036 B.n307 B.n306 585
R1037 B.n305 B.n304 585
R1038 B.n303 B.n302 585
R1039 B.n301 B.n300 585
R1040 B.n299 B.n298 585
R1041 B.n297 B.n296 585
R1042 B.n295 B.n294 585
R1043 B.n293 B.n292 585
R1044 B.n291 B.n290 585
R1045 B.n289 B.n288 585
R1046 B.n286 B.n285 585
R1047 B.n284 B.n283 585
R1048 B.n282 B.n281 585
R1049 B.n280 B.n279 585
R1050 B.n278 B.n277 585
R1051 B.n276 B.n275 585
R1052 B.n274 B.n273 585
R1053 B.n272 B.n271 585
R1054 B.n270 B.n269 585
R1055 B.n268 B.n267 585
R1056 B.n266 B.n265 585
R1057 B.n264 B.n263 585
R1058 B.n262 B.n261 585
R1059 B.n260 B.n259 585
R1060 B.n258 B.n257 585
R1061 B.n256 B.n255 585
R1062 B.n254 B.n253 585
R1063 B.n252 B.n251 585
R1064 B.n250 B.n249 585
R1065 B.n248 B.n247 585
R1066 B.n246 B.n245 585
R1067 B.n244 B.n243 585
R1068 B.n242 B.n241 585
R1069 B.n240 B.n239 585
R1070 B.n238 B.n237 585
R1071 B.n236 B.n235 585
R1072 B.n234 B.n233 585
R1073 B.n232 B.n231 585
R1074 B.n230 B.n229 585
R1075 B.n228 B.n227 585
R1076 B.n226 B.n225 585
R1077 B.n224 B.n223 585
R1078 B.n222 B.n221 585
R1079 B.n220 B.n219 585
R1080 B.n218 B.n217 585
R1081 B.n216 B.n215 585
R1082 B.n214 B.n213 585
R1083 B.n212 B.n211 585
R1084 B.n210 B.n209 585
R1085 B.n208 B.n207 585
R1086 B.n206 B.n205 585
R1087 B.n204 B.n203 585
R1088 B.n202 B.n201 585
R1089 B.n200 B.n199 585
R1090 B.n198 B.n197 585
R1091 B.n196 B.n195 585
R1092 B.n194 B.n193 585
R1093 B.n192 B.n191 585
R1094 B.n190 B.n189 585
R1095 B.n188 B.n187 585
R1096 B.n186 B.n185 585
R1097 B.n130 B.n129 585
R1098 B.n1068 B.n1067 585
R1099 B.n1062 B.n179 585
R1100 B.n179 B.n127 585
R1101 B.n1061 B.n126 585
R1102 B.n1072 B.n126 585
R1103 B.n1060 B.n125 585
R1104 B.n1073 B.n125 585
R1105 B.n1059 B.n124 585
R1106 B.n1074 B.n124 585
R1107 B.n1058 B.n1057 585
R1108 B.n1057 B.n120 585
R1109 B.n1056 B.n119 585
R1110 B.n1080 B.n119 585
R1111 B.n1055 B.n118 585
R1112 B.n1081 B.n118 585
R1113 B.n1054 B.n117 585
R1114 B.n1082 B.n117 585
R1115 B.n1053 B.n1052 585
R1116 B.n1052 B.n113 585
R1117 B.n1051 B.n112 585
R1118 B.n1088 B.n112 585
R1119 B.n1050 B.n111 585
R1120 B.n1089 B.n111 585
R1121 B.n1049 B.n110 585
R1122 B.n1090 B.n110 585
R1123 B.n1048 B.n1047 585
R1124 B.n1047 B.n106 585
R1125 B.n1046 B.n105 585
R1126 B.n1096 B.n105 585
R1127 B.n1045 B.n104 585
R1128 B.n1097 B.n104 585
R1129 B.n1044 B.n103 585
R1130 B.n1098 B.n103 585
R1131 B.n1043 B.n1042 585
R1132 B.n1042 B.n99 585
R1133 B.n1041 B.n98 585
R1134 B.n1104 B.n98 585
R1135 B.n1040 B.n97 585
R1136 B.n1105 B.n97 585
R1137 B.n1039 B.n96 585
R1138 B.n1106 B.n96 585
R1139 B.n1038 B.n1037 585
R1140 B.n1037 B.n92 585
R1141 B.n1036 B.n91 585
R1142 B.n1112 B.n91 585
R1143 B.n1035 B.n90 585
R1144 B.n1113 B.n90 585
R1145 B.n1034 B.n89 585
R1146 B.n1114 B.n89 585
R1147 B.n1033 B.n1032 585
R1148 B.n1032 B.n85 585
R1149 B.n1031 B.n84 585
R1150 B.n1120 B.n84 585
R1151 B.n1030 B.n83 585
R1152 B.n1121 B.n83 585
R1153 B.n1029 B.n82 585
R1154 B.n1122 B.n82 585
R1155 B.n1028 B.n1027 585
R1156 B.n1027 B.n78 585
R1157 B.n1026 B.n77 585
R1158 B.n1128 B.n77 585
R1159 B.n1025 B.n76 585
R1160 B.n1129 B.n76 585
R1161 B.n1024 B.n75 585
R1162 B.n1130 B.n75 585
R1163 B.n1023 B.n1022 585
R1164 B.n1022 B.n71 585
R1165 B.n1021 B.n70 585
R1166 B.n1136 B.n70 585
R1167 B.n1020 B.n69 585
R1168 B.n1137 B.n69 585
R1169 B.n1019 B.n68 585
R1170 B.n1138 B.n68 585
R1171 B.n1018 B.n1017 585
R1172 B.n1017 B.n64 585
R1173 B.n1016 B.n63 585
R1174 B.n1144 B.n63 585
R1175 B.n1015 B.n62 585
R1176 B.n1145 B.n62 585
R1177 B.n1014 B.n61 585
R1178 B.n1146 B.n61 585
R1179 B.n1013 B.n1012 585
R1180 B.n1012 B.n57 585
R1181 B.n1011 B.n56 585
R1182 B.n1152 B.n56 585
R1183 B.n1010 B.n55 585
R1184 B.n1153 B.n55 585
R1185 B.n1009 B.n54 585
R1186 B.n1154 B.n54 585
R1187 B.n1008 B.n1007 585
R1188 B.n1007 B.n50 585
R1189 B.n1006 B.n49 585
R1190 B.n1160 B.n49 585
R1191 B.n1005 B.n48 585
R1192 B.n1161 B.n48 585
R1193 B.n1004 B.n47 585
R1194 B.n1162 B.n47 585
R1195 B.n1003 B.n1002 585
R1196 B.n1002 B.n43 585
R1197 B.n1001 B.n42 585
R1198 B.n1168 B.n42 585
R1199 B.n1000 B.n41 585
R1200 B.n1169 B.n41 585
R1201 B.n999 B.n40 585
R1202 B.n1170 B.n40 585
R1203 B.n998 B.n997 585
R1204 B.n997 B.n36 585
R1205 B.n996 B.n35 585
R1206 B.n1176 B.n35 585
R1207 B.n995 B.n34 585
R1208 B.n1177 B.n34 585
R1209 B.n994 B.n33 585
R1210 B.n1178 B.n33 585
R1211 B.n993 B.n992 585
R1212 B.n992 B.n29 585
R1213 B.n991 B.n28 585
R1214 B.n1184 B.n28 585
R1215 B.n990 B.n27 585
R1216 B.n1185 B.n27 585
R1217 B.n989 B.n26 585
R1218 B.n1186 B.n26 585
R1219 B.n988 B.n987 585
R1220 B.n987 B.n22 585
R1221 B.n986 B.n21 585
R1222 B.n1192 B.n21 585
R1223 B.n985 B.n20 585
R1224 B.n1193 B.n20 585
R1225 B.n984 B.n19 585
R1226 B.n1194 B.n19 585
R1227 B.n983 B.n982 585
R1228 B.n982 B.n15 585
R1229 B.n981 B.n14 585
R1230 B.n1200 B.n14 585
R1231 B.n980 B.n13 585
R1232 B.n1201 B.n13 585
R1233 B.n979 B.n12 585
R1234 B.n1202 B.n12 585
R1235 B.n978 B.n977 585
R1236 B.n977 B.n8 585
R1237 B.n976 B.n7 585
R1238 B.n1208 B.n7 585
R1239 B.n975 B.n6 585
R1240 B.n1209 B.n6 585
R1241 B.n974 B.n5 585
R1242 B.n1210 B.n5 585
R1243 B.n973 B.n972 585
R1244 B.n972 B.n4 585
R1245 B.n971 B.n373 585
R1246 B.n971 B.n970 585
R1247 B.n961 B.n374 585
R1248 B.n375 B.n374 585
R1249 B.n963 B.n962 585
R1250 B.n964 B.n963 585
R1251 B.n960 B.n380 585
R1252 B.n380 B.n379 585
R1253 B.n959 B.n958 585
R1254 B.n958 B.n957 585
R1255 B.n382 B.n381 585
R1256 B.n383 B.n382 585
R1257 B.n950 B.n949 585
R1258 B.n951 B.n950 585
R1259 B.n948 B.n388 585
R1260 B.n388 B.n387 585
R1261 B.n947 B.n946 585
R1262 B.n946 B.n945 585
R1263 B.n390 B.n389 585
R1264 B.n391 B.n390 585
R1265 B.n938 B.n937 585
R1266 B.n939 B.n938 585
R1267 B.n936 B.n396 585
R1268 B.n396 B.n395 585
R1269 B.n935 B.n934 585
R1270 B.n934 B.n933 585
R1271 B.n398 B.n397 585
R1272 B.n399 B.n398 585
R1273 B.n926 B.n925 585
R1274 B.n927 B.n926 585
R1275 B.n924 B.n404 585
R1276 B.n404 B.n403 585
R1277 B.n923 B.n922 585
R1278 B.n922 B.n921 585
R1279 B.n406 B.n405 585
R1280 B.n407 B.n406 585
R1281 B.n914 B.n913 585
R1282 B.n915 B.n914 585
R1283 B.n912 B.n411 585
R1284 B.n415 B.n411 585
R1285 B.n911 B.n910 585
R1286 B.n910 B.n909 585
R1287 B.n413 B.n412 585
R1288 B.n414 B.n413 585
R1289 B.n902 B.n901 585
R1290 B.n903 B.n902 585
R1291 B.n900 B.n420 585
R1292 B.n420 B.n419 585
R1293 B.n899 B.n898 585
R1294 B.n898 B.n897 585
R1295 B.n422 B.n421 585
R1296 B.n423 B.n422 585
R1297 B.n890 B.n889 585
R1298 B.n891 B.n890 585
R1299 B.n888 B.n428 585
R1300 B.n428 B.n427 585
R1301 B.n887 B.n886 585
R1302 B.n886 B.n885 585
R1303 B.n430 B.n429 585
R1304 B.n431 B.n430 585
R1305 B.n878 B.n877 585
R1306 B.n879 B.n878 585
R1307 B.n876 B.n436 585
R1308 B.n436 B.n435 585
R1309 B.n875 B.n874 585
R1310 B.n874 B.n873 585
R1311 B.n438 B.n437 585
R1312 B.n439 B.n438 585
R1313 B.n866 B.n865 585
R1314 B.n867 B.n866 585
R1315 B.n864 B.n444 585
R1316 B.n444 B.n443 585
R1317 B.n863 B.n862 585
R1318 B.n862 B.n861 585
R1319 B.n446 B.n445 585
R1320 B.n447 B.n446 585
R1321 B.n854 B.n853 585
R1322 B.n855 B.n854 585
R1323 B.n852 B.n452 585
R1324 B.n452 B.n451 585
R1325 B.n851 B.n850 585
R1326 B.n850 B.n849 585
R1327 B.n454 B.n453 585
R1328 B.n455 B.n454 585
R1329 B.n842 B.n841 585
R1330 B.n843 B.n842 585
R1331 B.n840 B.n460 585
R1332 B.n460 B.n459 585
R1333 B.n839 B.n838 585
R1334 B.n838 B.n837 585
R1335 B.n462 B.n461 585
R1336 B.n463 B.n462 585
R1337 B.n830 B.n829 585
R1338 B.n831 B.n830 585
R1339 B.n828 B.n468 585
R1340 B.n468 B.n467 585
R1341 B.n827 B.n826 585
R1342 B.n826 B.n825 585
R1343 B.n470 B.n469 585
R1344 B.n471 B.n470 585
R1345 B.n818 B.n817 585
R1346 B.n819 B.n818 585
R1347 B.n816 B.n476 585
R1348 B.n476 B.n475 585
R1349 B.n815 B.n814 585
R1350 B.n814 B.n813 585
R1351 B.n478 B.n477 585
R1352 B.n479 B.n478 585
R1353 B.n806 B.n805 585
R1354 B.n807 B.n806 585
R1355 B.n804 B.n484 585
R1356 B.n484 B.n483 585
R1357 B.n803 B.n802 585
R1358 B.n802 B.n801 585
R1359 B.n486 B.n485 585
R1360 B.n487 B.n486 585
R1361 B.n794 B.n793 585
R1362 B.n795 B.n794 585
R1363 B.n792 B.n492 585
R1364 B.n492 B.n491 585
R1365 B.n791 B.n790 585
R1366 B.n790 B.n789 585
R1367 B.n494 B.n493 585
R1368 B.n495 B.n494 585
R1369 B.n782 B.n781 585
R1370 B.n783 B.n782 585
R1371 B.n780 B.n500 585
R1372 B.n500 B.n499 585
R1373 B.n779 B.n778 585
R1374 B.n778 B.n777 585
R1375 B.n502 B.n501 585
R1376 B.n503 B.n502 585
R1377 B.n770 B.n769 585
R1378 B.n771 B.n770 585
R1379 B.n768 B.n508 585
R1380 B.n508 B.n507 585
R1381 B.n767 B.n766 585
R1382 B.n766 B.n765 585
R1383 B.n510 B.n509 585
R1384 B.n511 B.n510 585
R1385 B.n761 B.n760 585
R1386 B.n514 B.n513 585
R1387 B.n757 B.n756 585
R1388 B.n758 B.n757 585
R1389 B.n755 B.n562 585
R1390 B.n754 B.n753 585
R1391 B.n752 B.n751 585
R1392 B.n750 B.n749 585
R1393 B.n748 B.n747 585
R1394 B.n746 B.n745 585
R1395 B.n744 B.n743 585
R1396 B.n742 B.n741 585
R1397 B.n740 B.n739 585
R1398 B.n738 B.n737 585
R1399 B.n736 B.n735 585
R1400 B.n734 B.n733 585
R1401 B.n732 B.n731 585
R1402 B.n730 B.n729 585
R1403 B.n728 B.n727 585
R1404 B.n726 B.n725 585
R1405 B.n724 B.n723 585
R1406 B.n722 B.n721 585
R1407 B.n720 B.n719 585
R1408 B.n718 B.n717 585
R1409 B.n716 B.n715 585
R1410 B.n714 B.n713 585
R1411 B.n712 B.n711 585
R1412 B.n710 B.n709 585
R1413 B.n708 B.n707 585
R1414 B.n706 B.n705 585
R1415 B.n704 B.n703 585
R1416 B.n702 B.n701 585
R1417 B.n700 B.n699 585
R1418 B.n698 B.n697 585
R1419 B.n696 B.n695 585
R1420 B.n694 B.n693 585
R1421 B.n692 B.n691 585
R1422 B.n690 B.n689 585
R1423 B.n688 B.n687 585
R1424 B.n686 B.n685 585
R1425 B.n684 B.n683 585
R1426 B.n682 B.n681 585
R1427 B.n680 B.n679 585
R1428 B.n678 B.n677 585
R1429 B.n676 B.n675 585
R1430 B.n673 B.n672 585
R1431 B.n671 B.n670 585
R1432 B.n669 B.n668 585
R1433 B.n667 B.n666 585
R1434 B.n665 B.n664 585
R1435 B.n663 B.n662 585
R1436 B.n661 B.n660 585
R1437 B.n659 B.n658 585
R1438 B.n657 B.n656 585
R1439 B.n655 B.n654 585
R1440 B.n653 B.n652 585
R1441 B.n651 B.n650 585
R1442 B.n649 B.n648 585
R1443 B.n647 B.n646 585
R1444 B.n645 B.n644 585
R1445 B.n643 B.n642 585
R1446 B.n641 B.n640 585
R1447 B.n639 B.n638 585
R1448 B.n637 B.n636 585
R1449 B.n635 B.n634 585
R1450 B.n633 B.n632 585
R1451 B.n631 B.n630 585
R1452 B.n629 B.n628 585
R1453 B.n627 B.n626 585
R1454 B.n625 B.n624 585
R1455 B.n623 B.n622 585
R1456 B.n621 B.n620 585
R1457 B.n619 B.n618 585
R1458 B.n617 B.n616 585
R1459 B.n615 B.n614 585
R1460 B.n613 B.n612 585
R1461 B.n611 B.n610 585
R1462 B.n609 B.n608 585
R1463 B.n607 B.n606 585
R1464 B.n605 B.n604 585
R1465 B.n603 B.n602 585
R1466 B.n601 B.n600 585
R1467 B.n599 B.n598 585
R1468 B.n597 B.n596 585
R1469 B.n595 B.n594 585
R1470 B.n593 B.n592 585
R1471 B.n591 B.n590 585
R1472 B.n589 B.n588 585
R1473 B.n587 B.n586 585
R1474 B.n585 B.n584 585
R1475 B.n583 B.n582 585
R1476 B.n581 B.n580 585
R1477 B.n579 B.n578 585
R1478 B.n577 B.n576 585
R1479 B.n575 B.n574 585
R1480 B.n573 B.n572 585
R1481 B.n571 B.n570 585
R1482 B.n569 B.n568 585
R1483 B.n762 B.n512 585
R1484 B.n512 B.n511 585
R1485 B.n764 B.n763 585
R1486 B.n765 B.n764 585
R1487 B.n506 B.n505 585
R1488 B.n507 B.n506 585
R1489 B.n773 B.n772 585
R1490 B.n772 B.n771 585
R1491 B.n774 B.n504 585
R1492 B.n504 B.n503 585
R1493 B.n776 B.n775 585
R1494 B.n777 B.n776 585
R1495 B.n498 B.n497 585
R1496 B.n499 B.n498 585
R1497 B.n785 B.n784 585
R1498 B.n784 B.n783 585
R1499 B.n786 B.n496 585
R1500 B.n496 B.n495 585
R1501 B.n788 B.n787 585
R1502 B.n789 B.n788 585
R1503 B.n490 B.n489 585
R1504 B.n491 B.n490 585
R1505 B.n797 B.n796 585
R1506 B.n796 B.n795 585
R1507 B.n798 B.n488 585
R1508 B.n488 B.n487 585
R1509 B.n800 B.n799 585
R1510 B.n801 B.n800 585
R1511 B.n482 B.n481 585
R1512 B.n483 B.n482 585
R1513 B.n809 B.n808 585
R1514 B.n808 B.n807 585
R1515 B.n810 B.n480 585
R1516 B.n480 B.n479 585
R1517 B.n812 B.n811 585
R1518 B.n813 B.n812 585
R1519 B.n474 B.n473 585
R1520 B.n475 B.n474 585
R1521 B.n821 B.n820 585
R1522 B.n820 B.n819 585
R1523 B.n822 B.n472 585
R1524 B.n472 B.n471 585
R1525 B.n824 B.n823 585
R1526 B.n825 B.n824 585
R1527 B.n466 B.n465 585
R1528 B.n467 B.n466 585
R1529 B.n833 B.n832 585
R1530 B.n832 B.n831 585
R1531 B.n834 B.n464 585
R1532 B.n464 B.n463 585
R1533 B.n836 B.n835 585
R1534 B.n837 B.n836 585
R1535 B.n458 B.n457 585
R1536 B.n459 B.n458 585
R1537 B.n845 B.n844 585
R1538 B.n844 B.n843 585
R1539 B.n846 B.n456 585
R1540 B.n456 B.n455 585
R1541 B.n848 B.n847 585
R1542 B.n849 B.n848 585
R1543 B.n450 B.n449 585
R1544 B.n451 B.n450 585
R1545 B.n857 B.n856 585
R1546 B.n856 B.n855 585
R1547 B.n858 B.n448 585
R1548 B.n448 B.n447 585
R1549 B.n860 B.n859 585
R1550 B.n861 B.n860 585
R1551 B.n442 B.n441 585
R1552 B.n443 B.n442 585
R1553 B.n869 B.n868 585
R1554 B.n868 B.n867 585
R1555 B.n870 B.n440 585
R1556 B.n440 B.n439 585
R1557 B.n872 B.n871 585
R1558 B.n873 B.n872 585
R1559 B.n434 B.n433 585
R1560 B.n435 B.n434 585
R1561 B.n881 B.n880 585
R1562 B.n880 B.n879 585
R1563 B.n882 B.n432 585
R1564 B.n432 B.n431 585
R1565 B.n884 B.n883 585
R1566 B.n885 B.n884 585
R1567 B.n426 B.n425 585
R1568 B.n427 B.n426 585
R1569 B.n893 B.n892 585
R1570 B.n892 B.n891 585
R1571 B.n894 B.n424 585
R1572 B.n424 B.n423 585
R1573 B.n896 B.n895 585
R1574 B.n897 B.n896 585
R1575 B.n418 B.n417 585
R1576 B.n419 B.n418 585
R1577 B.n905 B.n904 585
R1578 B.n904 B.n903 585
R1579 B.n906 B.n416 585
R1580 B.n416 B.n414 585
R1581 B.n908 B.n907 585
R1582 B.n909 B.n908 585
R1583 B.n410 B.n409 585
R1584 B.n415 B.n410 585
R1585 B.n917 B.n916 585
R1586 B.n916 B.n915 585
R1587 B.n918 B.n408 585
R1588 B.n408 B.n407 585
R1589 B.n920 B.n919 585
R1590 B.n921 B.n920 585
R1591 B.n402 B.n401 585
R1592 B.n403 B.n402 585
R1593 B.n929 B.n928 585
R1594 B.n928 B.n927 585
R1595 B.n930 B.n400 585
R1596 B.n400 B.n399 585
R1597 B.n932 B.n931 585
R1598 B.n933 B.n932 585
R1599 B.n394 B.n393 585
R1600 B.n395 B.n394 585
R1601 B.n941 B.n940 585
R1602 B.n940 B.n939 585
R1603 B.n942 B.n392 585
R1604 B.n392 B.n391 585
R1605 B.n944 B.n943 585
R1606 B.n945 B.n944 585
R1607 B.n386 B.n385 585
R1608 B.n387 B.n386 585
R1609 B.n953 B.n952 585
R1610 B.n952 B.n951 585
R1611 B.n954 B.n384 585
R1612 B.n384 B.n383 585
R1613 B.n956 B.n955 585
R1614 B.n957 B.n956 585
R1615 B.n378 B.n377 585
R1616 B.n379 B.n378 585
R1617 B.n966 B.n965 585
R1618 B.n965 B.n964 585
R1619 B.n967 B.n376 585
R1620 B.n376 B.n375 585
R1621 B.n969 B.n968 585
R1622 B.n970 B.n969 585
R1623 B.n2 B.n0 585
R1624 B.n4 B.n2 585
R1625 B.n3 B.n1 585
R1626 B.n1209 B.n3 585
R1627 B.n1207 B.n1206 585
R1628 B.n1208 B.n1207 585
R1629 B.n1205 B.n9 585
R1630 B.n9 B.n8 585
R1631 B.n1204 B.n1203 585
R1632 B.n1203 B.n1202 585
R1633 B.n11 B.n10 585
R1634 B.n1201 B.n11 585
R1635 B.n1199 B.n1198 585
R1636 B.n1200 B.n1199 585
R1637 B.n1197 B.n16 585
R1638 B.n16 B.n15 585
R1639 B.n1196 B.n1195 585
R1640 B.n1195 B.n1194 585
R1641 B.n18 B.n17 585
R1642 B.n1193 B.n18 585
R1643 B.n1191 B.n1190 585
R1644 B.n1192 B.n1191 585
R1645 B.n1189 B.n23 585
R1646 B.n23 B.n22 585
R1647 B.n1188 B.n1187 585
R1648 B.n1187 B.n1186 585
R1649 B.n25 B.n24 585
R1650 B.n1185 B.n25 585
R1651 B.n1183 B.n1182 585
R1652 B.n1184 B.n1183 585
R1653 B.n1181 B.n30 585
R1654 B.n30 B.n29 585
R1655 B.n1180 B.n1179 585
R1656 B.n1179 B.n1178 585
R1657 B.n32 B.n31 585
R1658 B.n1177 B.n32 585
R1659 B.n1175 B.n1174 585
R1660 B.n1176 B.n1175 585
R1661 B.n1173 B.n37 585
R1662 B.n37 B.n36 585
R1663 B.n1172 B.n1171 585
R1664 B.n1171 B.n1170 585
R1665 B.n39 B.n38 585
R1666 B.n1169 B.n39 585
R1667 B.n1167 B.n1166 585
R1668 B.n1168 B.n1167 585
R1669 B.n1165 B.n44 585
R1670 B.n44 B.n43 585
R1671 B.n1164 B.n1163 585
R1672 B.n1163 B.n1162 585
R1673 B.n46 B.n45 585
R1674 B.n1161 B.n46 585
R1675 B.n1159 B.n1158 585
R1676 B.n1160 B.n1159 585
R1677 B.n1157 B.n51 585
R1678 B.n51 B.n50 585
R1679 B.n1156 B.n1155 585
R1680 B.n1155 B.n1154 585
R1681 B.n53 B.n52 585
R1682 B.n1153 B.n53 585
R1683 B.n1151 B.n1150 585
R1684 B.n1152 B.n1151 585
R1685 B.n1149 B.n58 585
R1686 B.n58 B.n57 585
R1687 B.n1148 B.n1147 585
R1688 B.n1147 B.n1146 585
R1689 B.n60 B.n59 585
R1690 B.n1145 B.n60 585
R1691 B.n1143 B.n1142 585
R1692 B.n1144 B.n1143 585
R1693 B.n1141 B.n65 585
R1694 B.n65 B.n64 585
R1695 B.n1140 B.n1139 585
R1696 B.n1139 B.n1138 585
R1697 B.n67 B.n66 585
R1698 B.n1137 B.n67 585
R1699 B.n1135 B.n1134 585
R1700 B.n1136 B.n1135 585
R1701 B.n1133 B.n72 585
R1702 B.n72 B.n71 585
R1703 B.n1132 B.n1131 585
R1704 B.n1131 B.n1130 585
R1705 B.n74 B.n73 585
R1706 B.n1129 B.n74 585
R1707 B.n1127 B.n1126 585
R1708 B.n1128 B.n1127 585
R1709 B.n1125 B.n79 585
R1710 B.n79 B.n78 585
R1711 B.n1124 B.n1123 585
R1712 B.n1123 B.n1122 585
R1713 B.n81 B.n80 585
R1714 B.n1121 B.n81 585
R1715 B.n1119 B.n1118 585
R1716 B.n1120 B.n1119 585
R1717 B.n1117 B.n86 585
R1718 B.n86 B.n85 585
R1719 B.n1116 B.n1115 585
R1720 B.n1115 B.n1114 585
R1721 B.n88 B.n87 585
R1722 B.n1113 B.n88 585
R1723 B.n1111 B.n1110 585
R1724 B.n1112 B.n1111 585
R1725 B.n1109 B.n93 585
R1726 B.n93 B.n92 585
R1727 B.n1108 B.n1107 585
R1728 B.n1107 B.n1106 585
R1729 B.n95 B.n94 585
R1730 B.n1105 B.n95 585
R1731 B.n1103 B.n1102 585
R1732 B.n1104 B.n1103 585
R1733 B.n1101 B.n100 585
R1734 B.n100 B.n99 585
R1735 B.n1100 B.n1099 585
R1736 B.n1099 B.n1098 585
R1737 B.n102 B.n101 585
R1738 B.n1097 B.n102 585
R1739 B.n1095 B.n1094 585
R1740 B.n1096 B.n1095 585
R1741 B.n1093 B.n107 585
R1742 B.n107 B.n106 585
R1743 B.n1092 B.n1091 585
R1744 B.n1091 B.n1090 585
R1745 B.n109 B.n108 585
R1746 B.n1089 B.n109 585
R1747 B.n1087 B.n1086 585
R1748 B.n1088 B.n1087 585
R1749 B.n1085 B.n114 585
R1750 B.n114 B.n113 585
R1751 B.n1084 B.n1083 585
R1752 B.n1083 B.n1082 585
R1753 B.n116 B.n115 585
R1754 B.n1081 B.n116 585
R1755 B.n1079 B.n1078 585
R1756 B.n1080 B.n1079 585
R1757 B.n1077 B.n121 585
R1758 B.n121 B.n120 585
R1759 B.n1076 B.n1075 585
R1760 B.n1075 B.n1074 585
R1761 B.n123 B.n122 585
R1762 B.n1073 B.n123 585
R1763 B.n1071 B.n1070 585
R1764 B.n1072 B.n1071 585
R1765 B.n1069 B.n128 585
R1766 B.n128 B.n127 585
R1767 B.n1212 B.n1211 585
R1768 B.n1211 B.n1210 585
R1769 B.n760 B.n512 506.916
R1770 B.n1067 B.n128 506.916
R1771 B.n568 B.n510 506.916
R1772 B.n1064 B.n179 506.916
R1773 B.n565 B.t14 377.308
R1774 B.n180 B.t17 377.308
R1775 B.n563 B.t11 377.308
R1776 B.n182 B.t20 377.308
R1777 B.n566 B.t13 294.303
R1778 B.n181 B.t18 294.303
R1779 B.n564 B.t10 294.303
R1780 B.n183 B.t21 294.303
R1781 B.n565 B.t12 287.003
R1782 B.n563 B.t8 287.003
R1783 B.n182 B.t19 287.003
R1784 B.n180 B.t15 287.003
R1785 B.n1065 B.n177 256.663
R1786 B.n1065 B.n176 256.663
R1787 B.n1065 B.n175 256.663
R1788 B.n1065 B.n174 256.663
R1789 B.n1065 B.n173 256.663
R1790 B.n1065 B.n172 256.663
R1791 B.n1065 B.n171 256.663
R1792 B.n1065 B.n170 256.663
R1793 B.n1065 B.n169 256.663
R1794 B.n1065 B.n168 256.663
R1795 B.n1065 B.n167 256.663
R1796 B.n1065 B.n166 256.663
R1797 B.n1065 B.n165 256.663
R1798 B.n1065 B.n164 256.663
R1799 B.n1065 B.n163 256.663
R1800 B.n1065 B.n162 256.663
R1801 B.n1065 B.n161 256.663
R1802 B.n1065 B.n160 256.663
R1803 B.n1065 B.n159 256.663
R1804 B.n1065 B.n158 256.663
R1805 B.n1065 B.n157 256.663
R1806 B.n1065 B.n156 256.663
R1807 B.n1065 B.n155 256.663
R1808 B.n1065 B.n154 256.663
R1809 B.n1065 B.n153 256.663
R1810 B.n1065 B.n152 256.663
R1811 B.n1065 B.n151 256.663
R1812 B.n1065 B.n150 256.663
R1813 B.n1065 B.n149 256.663
R1814 B.n1065 B.n148 256.663
R1815 B.n1065 B.n147 256.663
R1816 B.n1065 B.n146 256.663
R1817 B.n1065 B.n145 256.663
R1818 B.n1065 B.n144 256.663
R1819 B.n1065 B.n143 256.663
R1820 B.n1065 B.n142 256.663
R1821 B.n1065 B.n141 256.663
R1822 B.n1065 B.n140 256.663
R1823 B.n1065 B.n139 256.663
R1824 B.n1065 B.n138 256.663
R1825 B.n1065 B.n137 256.663
R1826 B.n1065 B.n136 256.663
R1827 B.n1065 B.n135 256.663
R1828 B.n1065 B.n134 256.663
R1829 B.n1065 B.n133 256.663
R1830 B.n1065 B.n132 256.663
R1831 B.n1065 B.n131 256.663
R1832 B.n1066 B.n1065 256.663
R1833 B.n759 B.n758 256.663
R1834 B.n758 B.n515 256.663
R1835 B.n758 B.n516 256.663
R1836 B.n758 B.n517 256.663
R1837 B.n758 B.n518 256.663
R1838 B.n758 B.n519 256.663
R1839 B.n758 B.n520 256.663
R1840 B.n758 B.n521 256.663
R1841 B.n758 B.n522 256.663
R1842 B.n758 B.n523 256.663
R1843 B.n758 B.n524 256.663
R1844 B.n758 B.n525 256.663
R1845 B.n758 B.n526 256.663
R1846 B.n758 B.n527 256.663
R1847 B.n758 B.n528 256.663
R1848 B.n758 B.n529 256.663
R1849 B.n758 B.n530 256.663
R1850 B.n758 B.n531 256.663
R1851 B.n758 B.n532 256.663
R1852 B.n758 B.n533 256.663
R1853 B.n758 B.n534 256.663
R1854 B.n758 B.n535 256.663
R1855 B.n758 B.n536 256.663
R1856 B.n758 B.n537 256.663
R1857 B.n758 B.n538 256.663
R1858 B.n758 B.n539 256.663
R1859 B.n758 B.n540 256.663
R1860 B.n758 B.n541 256.663
R1861 B.n758 B.n542 256.663
R1862 B.n758 B.n543 256.663
R1863 B.n758 B.n544 256.663
R1864 B.n758 B.n545 256.663
R1865 B.n758 B.n546 256.663
R1866 B.n758 B.n547 256.663
R1867 B.n758 B.n548 256.663
R1868 B.n758 B.n549 256.663
R1869 B.n758 B.n550 256.663
R1870 B.n758 B.n551 256.663
R1871 B.n758 B.n552 256.663
R1872 B.n758 B.n553 256.663
R1873 B.n758 B.n554 256.663
R1874 B.n758 B.n555 256.663
R1875 B.n758 B.n556 256.663
R1876 B.n758 B.n557 256.663
R1877 B.n758 B.n558 256.663
R1878 B.n758 B.n559 256.663
R1879 B.n758 B.n560 256.663
R1880 B.n758 B.n561 256.663
R1881 B.n764 B.n512 163.367
R1882 B.n764 B.n506 163.367
R1883 B.n772 B.n506 163.367
R1884 B.n772 B.n504 163.367
R1885 B.n776 B.n504 163.367
R1886 B.n776 B.n498 163.367
R1887 B.n784 B.n498 163.367
R1888 B.n784 B.n496 163.367
R1889 B.n788 B.n496 163.367
R1890 B.n788 B.n490 163.367
R1891 B.n796 B.n490 163.367
R1892 B.n796 B.n488 163.367
R1893 B.n800 B.n488 163.367
R1894 B.n800 B.n482 163.367
R1895 B.n808 B.n482 163.367
R1896 B.n808 B.n480 163.367
R1897 B.n812 B.n480 163.367
R1898 B.n812 B.n474 163.367
R1899 B.n820 B.n474 163.367
R1900 B.n820 B.n472 163.367
R1901 B.n824 B.n472 163.367
R1902 B.n824 B.n466 163.367
R1903 B.n832 B.n466 163.367
R1904 B.n832 B.n464 163.367
R1905 B.n836 B.n464 163.367
R1906 B.n836 B.n458 163.367
R1907 B.n844 B.n458 163.367
R1908 B.n844 B.n456 163.367
R1909 B.n848 B.n456 163.367
R1910 B.n848 B.n450 163.367
R1911 B.n856 B.n450 163.367
R1912 B.n856 B.n448 163.367
R1913 B.n860 B.n448 163.367
R1914 B.n860 B.n442 163.367
R1915 B.n868 B.n442 163.367
R1916 B.n868 B.n440 163.367
R1917 B.n872 B.n440 163.367
R1918 B.n872 B.n434 163.367
R1919 B.n880 B.n434 163.367
R1920 B.n880 B.n432 163.367
R1921 B.n884 B.n432 163.367
R1922 B.n884 B.n426 163.367
R1923 B.n892 B.n426 163.367
R1924 B.n892 B.n424 163.367
R1925 B.n896 B.n424 163.367
R1926 B.n896 B.n418 163.367
R1927 B.n904 B.n418 163.367
R1928 B.n904 B.n416 163.367
R1929 B.n908 B.n416 163.367
R1930 B.n908 B.n410 163.367
R1931 B.n916 B.n410 163.367
R1932 B.n916 B.n408 163.367
R1933 B.n920 B.n408 163.367
R1934 B.n920 B.n402 163.367
R1935 B.n928 B.n402 163.367
R1936 B.n928 B.n400 163.367
R1937 B.n932 B.n400 163.367
R1938 B.n932 B.n394 163.367
R1939 B.n940 B.n394 163.367
R1940 B.n940 B.n392 163.367
R1941 B.n944 B.n392 163.367
R1942 B.n944 B.n386 163.367
R1943 B.n952 B.n386 163.367
R1944 B.n952 B.n384 163.367
R1945 B.n956 B.n384 163.367
R1946 B.n956 B.n378 163.367
R1947 B.n965 B.n378 163.367
R1948 B.n965 B.n376 163.367
R1949 B.n969 B.n376 163.367
R1950 B.n969 B.n2 163.367
R1951 B.n1211 B.n2 163.367
R1952 B.n1211 B.n3 163.367
R1953 B.n1207 B.n3 163.367
R1954 B.n1207 B.n9 163.367
R1955 B.n1203 B.n9 163.367
R1956 B.n1203 B.n11 163.367
R1957 B.n1199 B.n11 163.367
R1958 B.n1199 B.n16 163.367
R1959 B.n1195 B.n16 163.367
R1960 B.n1195 B.n18 163.367
R1961 B.n1191 B.n18 163.367
R1962 B.n1191 B.n23 163.367
R1963 B.n1187 B.n23 163.367
R1964 B.n1187 B.n25 163.367
R1965 B.n1183 B.n25 163.367
R1966 B.n1183 B.n30 163.367
R1967 B.n1179 B.n30 163.367
R1968 B.n1179 B.n32 163.367
R1969 B.n1175 B.n32 163.367
R1970 B.n1175 B.n37 163.367
R1971 B.n1171 B.n37 163.367
R1972 B.n1171 B.n39 163.367
R1973 B.n1167 B.n39 163.367
R1974 B.n1167 B.n44 163.367
R1975 B.n1163 B.n44 163.367
R1976 B.n1163 B.n46 163.367
R1977 B.n1159 B.n46 163.367
R1978 B.n1159 B.n51 163.367
R1979 B.n1155 B.n51 163.367
R1980 B.n1155 B.n53 163.367
R1981 B.n1151 B.n53 163.367
R1982 B.n1151 B.n58 163.367
R1983 B.n1147 B.n58 163.367
R1984 B.n1147 B.n60 163.367
R1985 B.n1143 B.n60 163.367
R1986 B.n1143 B.n65 163.367
R1987 B.n1139 B.n65 163.367
R1988 B.n1139 B.n67 163.367
R1989 B.n1135 B.n67 163.367
R1990 B.n1135 B.n72 163.367
R1991 B.n1131 B.n72 163.367
R1992 B.n1131 B.n74 163.367
R1993 B.n1127 B.n74 163.367
R1994 B.n1127 B.n79 163.367
R1995 B.n1123 B.n79 163.367
R1996 B.n1123 B.n81 163.367
R1997 B.n1119 B.n81 163.367
R1998 B.n1119 B.n86 163.367
R1999 B.n1115 B.n86 163.367
R2000 B.n1115 B.n88 163.367
R2001 B.n1111 B.n88 163.367
R2002 B.n1111 B.n93 163.367
R2003 B.n1107 B.n93 163.367
R2004 B.n1107 B.n95 163.367
R2005 B.n1103 B.n95 163.367
R2006 B.n1103 B.n100 163.367
R2007 B.n1099 B.n100 163.367
R2008 B.n1099 B.n102 163.367
R2009 B.n1095 B.n102 163.367
R2010 B.n1095 B.n107 163.367
R2011 B.n1091 B.n107 163.367
R2012 B.n1091 B.n109 163.367
R2013 B.n1087 B.n109 163.367
R2014 B.n1087 B.n114 163.367
R2015 B.n1083 B.n114 163.367
R2016 B.n1083 B.n116 163.367
R2017 B.n1079 B.n116 163.367
R2018 B.n1079 B.n121 163.367
R2019 B.n1075 B.n121 163.367
R2020 B.n1075 B.n123 163.367
R2021 B.n1071 B.n123 163.367
R2022 B.n1071 B.n128 163.367
R2023 B.n757 B.n514 163.367
R2024 B.n757 B.n562 163.367
R2025 B.n753 B.n752 163.367
R2026 B.n749 B.n748 163.367
R2027 B.n745 B.n744 163.367
R2028 B.n741 B.n740 163.367
R2029 B.n737 B.n736 163.367
R2030 B.n733 B.n732 163.367
R2031 B.n729 B.n728 163.367
R2032 B.n725 B.n724 163.367
R2033 B.n721 B.n720 163.367
R2034 B.n717 B.n716 163.367
R2035 B.n713 B.n712 163.367
R2036 B.n709 B.n708 163.367
R2037 B.n705 B.n704 163.367
R2038 B.n701 B.n700 163.367
R2039 B.n697 B.n696 163.367
R2040 B.n693 B.n692 163.367
R2041 B.n689 B.n688 163.367
R2042 B.n685 B.n684 163.367
R2043 B.n681 B.n680 163.367
R2044 B.n677 B.n676 163.367
R2045 B.n672 B.n671 163.367
R2046 B.n668 B.n667 163.367
R2047 B.n664 B.n663 163.367
R2048 B.n660 B.n659 163.367
R2049 B.n656 B.n655 163.367
R2050 B.n652 B.n651 163.367
R2051 B.n648 B.n647 163.367
R2052 B.n644 B.n643 163.367
R2053 B.n640 B.n639 163.367
R2054 B.n636 B.n635 163.367
R2055 B.n632 B.n631 163.367
R2056 B.n628 B.n627 163.367
R2057 B.n624 B.n623 163.367
R2058 B.n620 B.n619 163.367
R2059 B.n616 B.n615 163.367
R2060 B.n612 B.n611 163.367
R2061 B.n608 B.n607 163.367
R2062 B.n604 B.n603 163.367
R2063 B.n600 B.n599 163.367
R2064 B.n596 B.n595 163.367
R2065 B.n592 B.n591 163.367
R2066 B.n588 B.n587 163.367
R2067 B.n584 B.n583 163.367
R2068 B.n580 B.n579 163.367
R2069 B.n576 B.n575 163.367
R2070 B.n572 B.n571 163.367
R2071 B.n766 B.n510 163.367
R2072 B.n766 B.n508 163.367
R2073 B.n770 B.n508 163.367
R2074 B.n770 B.n502 163.367
R2075 B.n778 B.n502 163.367
R2076 B.n778 B.n500 163.367
R2077 B.n782 B.n500 163.367
R2078 B.n782 B.n494 163.367
R2079 B.n790 B.n494 163.367
R2080 B.n790 B.n492 163.367
R2081 B.n794 B.n492 163.367
R2082 B.n794 B.n486 163.367
R2083 B.n802 B.n486 163.367
R2084 B.n802 B.n484 163.367
R2085 B.n806 B.n484 163.367
R2086 B.n806 B.n478 163.367
R2087 B.n814 B.n478 163.367
R2088 B.n814 B.n476 163.367
R2089 B.n818 B.n476 163.367
R2090 B.n818 B.n470 163.367
R2091 B.n826 B.n470 163.367
R2092 B.n826 B.n468 163.367
R2093 B.n830 B.n468 163.367
R2094 B.n830 B.n462 163.367
R2095 B.n838 B.n462 163.367
R2096 B.n838 B.n460 163.367
R2097 B.n842 B.n460 163.367
R2098 B.n842 B.n454 163.367
R2099 B.n850 B.n454 163.367
R2100 B.n850 B.n452 163.367
R2101 B.n854 B.n452 163.367
R2102 B.n854 B.n446 163.367
R2103 B.n862 B.n446 163.367
R2104 B.n862 B.n444 163.367
R2105 B.n866 B.n444 163.367
R2106 B.n866 B.n438 163.367
R2107 B.n874 B.n438 163.367
R2108 B.n874 B.n436 163.367
R2109 B.n878 B.n436 163.367
R2110 B.n878 B.n430 163.367
R2111 B.n886 B.n430 163.367
R2112 B.n886 B.n428 163.367
R2113 B.n890 B.n428 163.367
R2114 B.n890 B.n422 163.367
R2115 B.n898 B.n422 163.367
R2116 B.n898 B.n420 163.367
R2117 B.n902 B.n420 163.367
R2118 B.n902 B.n413 163.367
R2119 B.n910 B.n413 163.367
R2120 B.n910 B.n411 163.367
R2121 B.n914 B.n411 163.367
R2122 B.n914 B.n406 163.367
R2123 B.n922 B.n406 163.367
R2124 B.n922 B.n404 163.367
R2125 B.n926 B.n404 163.367
R2126 B.n926 B.n398 163.367
R2127 B.n934 B.n398 163.367
R2128 B.n934 B.n396 163.367
R2129 B.n938 B.n396 163.367
R2130 B.n938 B.n390 163.367
R2131 B.n946 B.n390 163.367
R2132 B.n946 B.n388 163.367
R2133 B.n950 B.n388 163.367
R2134 B.n950 B.n382 163.367
R2135 B.n958 B.n382 163.367
R2136 B.n958 B.n380 163.367
R2137 B.n963 B.n380 163.367
R2138 B.n963 B.n374 163.367
R2139 B.n971 B.n374 163.367
R2140 B.n972 B.n971 163.367
R2141 B.n972 B.n5 163.367
R2142 B.n6 B.n5 163.367
R2143 B.n7 B.n6 163.367
R2144 B.n977 B.n7 163.367
R2145 B.n977 B.n12 163.367
R2146 B.n13 B.n12 163.367
R2147 B.n14 B.n13 163.367
R2148 B.n982 B.n14 163.367
R2149 B.n982 B.n19 163.367
R2150 B.n20 B.n19 163.367
R2151 B.n21 B.n20 163.367
R2152 B.n987 B.n21 163.367
R2153 B.n987 B.n26 163.367
R2154 B.n27 B.n26 163.367
R2155 B.n28 B.n27 163.367
R2156 B.n992 B.n28 163.367
R2157 B.n992 B.n33 163.367
R2158 B.n34 B.n33 163.367
R2159 B.n35 B.n34 163.367
R2160 B.n997 B.n35 163.367
R2161 B.n997 B.n40 163.367
R2162 B.n41 B.n40 163.367
R2163 B.n42 B.n41 163.367
R2164 B.n1002 B.n42 163.367
R2165 B.n1002 B.n47 163.367
R2166 B.n48 B.n47 163.367
R2167 B.n49 B.n48 163.367
R2168 B.n1007 B.n49 163.367
R2169 B.n1007 B.n54 163.367
R2170 B.n55 B.n54 163.367
R2171 B.n56 B.n55 163.367
R2172 B.n1012 B.n56 163.367
R2173 B.n1012 B.n61 163.367
R2174 B.n62 B.n61 163.367
R2175 B.n63 B.n62 163.367
R2176 B.n1017 B.n63 163.367
R2177 B.n1017 B.n68 163.367
R2178 B.n69 B.n68 163.367
R2179 B.n70 B.n69 163.367
R2180 B.n1022 B.n70 163.367
R2181 B.n1022 B.n75 163.367
R2182 B.n76 B.n75 163.367
R2183 B.n77 B.n76 163.367
R2184 B.n1027 B.n77 163.367
R2185 B.n1027 B.n82 163.367
R2186 B.n83 B.n82 163.367
R2187 B.n84 B.n83 163.367
R2188 B.n1032 B.n84 163.367
R2189 B.n1032 B.n89 163.367
R2190 B.n90 B.n89 163.367
R2191 B.n91 B.n90 163.367
R2192 B.n1037 B.n91 163.367
R2193 B.n1037 B.n96 163.367
R2194 B.n97 B.n96 163.367
R2195 B.n98 B.n97 163.367
R2196 B.n1042 B.n98 163.367
R2197 B.n1042 B.n103 163.367
R2198 B.n104 B.n103 163.367
R2199 B.n105 B.n104 163.367
R2200 B.n1047 B.n105 163.367
R2201 B.n1047 B.n110 163.367
R2202 B.n111 B.n110 163.367
R2203 B.n112 B.n111 163.367
R2204 B.n1052 B.n112 163.367
R2205 B.n1052 B.n117 163.367
R2206 B.n118 B.n117 163.367
R2207 B.n119 B.n118 163.367
R2208 B.n1057 B.n119 163.367
R2209 B.n1057 B.n124 163.367
R2210 B.n125 B.n124 163.367
R2211 B.n126 B.n125 163.367
R2212 B.n179 B.n126 163.367
R2213 B.n185 B.n130 163.367
R2214 B.n189 B.n188 163.367
R2215 B.n193 B.n192 163.367
R2216 B.n197 B.n196 163.367
R2217 B.n201 B.n200 163.367
R2218 B.n205 B.n204 163.367
R2219 B.n209 B.n208 163.367
R2220 B.n213 B.n212 163.367
R2221 B.n217 B.n216 163.367
R2222 B.n221 B.n220 163.367
R2223 B.n225 B.n224 163.367
R2224 B.n229 B.n228 163.367
R2225 B.n233 B.n232 163.367
R2226 B.n237 B.n236 163.367
R2227 B.n241 B.n240 163.367
R2228 B.n245 B.n244 163.367
R2229 B.n249 B.n248 163.367
R2230 B.n253 B.n252 163.367
R2231 B.n257 B.n256 163.367
R2232 B.n261 B.n260 163.367
R2233 B.n265 B.n264 163.367
R2234 B.n269 B.n268 163.367
R2235 B.n273 B.n272 163.367
R2236 B.n277 B.n276 163.367
R2237 B.n281 B.n280 163.367
R2238 B.n285 B.n284 163.367
R2239 B.n290 B.n289 163.367
R2240 B.n294 B.n293 163.367
R2241 B.n298 B.n297 163.367
R2242 B.n302 B.n301 163.367
R2243 B.n306 B.n305 163.367
R2244 B.n310 B.n309 163.367
R2245 B.n314 B.n313 163.367
R2246 B.n318 B.n317 163.367
R2247 B.n322 B.n321 163.367
R2248 B.n326 B.n325 163.367
R2249 B.n330 B.n329 163.367
R2250 B.n334 B.n333 163.367
R2251 B.n338 B.n337 163.367
R2252 B.n342 B.n341 163.367
R2253 B.n346 B.n345 163.367
R2254 B.n350 B.n349 163.367
R2255 B.n354 B.n353 163.367
R2256 B.n358 B.n357 163.367
R2257 B.n362 B.n361 163.367
R2258 B.n366 B.n365 163.367
R2259 B.n370 B.n369 163.367
R2260 B.n1064 B.n178 163.367
R2261 B.n566 B.n565 83.0066
R2262 B.n564 B.n563 83.0066
R2263 B.n183 B.n182 83.0066
R2264 B.n181 B.n180 83.0066
R2265 B.n758 B.n511 77.6763
R2266 B.n1065 B.n127 77.6763
R2267 B.n760 B.n759 71.676
R2268 B.n562 B.n515 71.676
R2269 B.n752 B.n516 71.676
R2270 B.n748 B.n517 71.676
R2271 B.n744 B.n518 71.676
R2272 B.n740 B.n519 71.676
R2273 B.n736 B.n520 71.676
R2274 B.n732 B.n521 71.676
R2275 B.n728 B.n522 71.676
R2276 B.n724 B.n523 71.676
R2277 B.n720 B.n524 71.676
R2278 B.n716 B.n525 71.676
R2279 B.n712 B.n526 71.676
R2280 B.n708 B.n527 71.676
R2281 B.n704 B.n528 71.676
R2282 B.n700 B.n529 71.676
R2283 B.n696 B.n530 71.676
R2284 B.n692 B.n531 71.676
R2285 B.n688 B.n532 71.676
R2286 B.n684 B.n533 71.676
R2287 B.n680 B.n534 71.676
R2288 B.n676 B.n535 71.676
R2289 B.n671 B.n536 71.676
R2290 B.n667 B.n537 71.676
R2291 B.n663 B.n538 71.676
R2292 B.n659 B.n539 71.676
R2293 B.n655 B.n540 71.676
R2294 B.n651 B.n541 71.676
R2295 B.n647 B.n542 71.676
R2296 B.n643 B.n543 71.676
R2297 B.n639 B.n544 71.676
R2298 B.n635 B.n545 71.676
R2299 B.n631 B.n546 71.676
R2300 B.n627 B.n547 71.676
R2301 B.n623 B.n548 71.676
R2302 B.n619 B.n549 71.676
R2303 B.n615 B.n550 71.676
R2304 B.n611 B.n551 71.676
R2305 B.n607 B.n552 71.676
R2306 B.n603 B.n553 71.676
R2307 B.n599 B.n554 71.676
R2308 B.n595 B.n555 71.676
R2309 B.n591 B.n556 71.676
R2310 B.n587 B.n557 71.676
R2311 B.n583 B.n558 71.676
R2312 B.n579 B.n559 71.676
R2313 B.n575 B.n560 71.676
R2314 B.n571 B.n561 71.676
R2315 B.n1067 B.n1066 71.676
R2316 B.n185 B.n131 71.676
R2317 B.n189 B.n132 71.676
R2318 B.n193 B.n133 71.676
R2319 B.n197 B.n134 71.676
R2320 B.n201 B.n135 71.676
R2321 B.n205 B.n136 71.676
R2322 B.n209 B.n137 71.676
R2323 B.n213 B.n138 71.676
R2324 B.n217 B.n139 71.676
R2325 B.n221 B.n140 71.676
R2326 B.n225 B.n141 71.676
R2327 B.n229 B.n142 71.676
R2328 B.n233 B.n143 71.676
R2329 B.n237 B.n144 71.676
R2330 B.n241 B.n145 71.676
R2331 B.n245 B.n146 71.676
R2332 B.n249 B.n147 71.676
R2333 B.n253 B.n148 71.676
R2334 B.n257 B.n149 71.676
R2335 B.n261 B.n150 71.676
R2336 B.n265 B.n151 71.676
R2337 B.n269 B.n152 71.676
R2338 B.n273 B.n153 71.676
R2339 B.n277 B.n154 71.676
R2340 B.n281 B.n155 71.676
R2341 B.n285 B.n156 71.676
R2342 B.n290 B.n157 71.676
R2343 B.n294 B.n158 71.676
R2344 B.n298 B.n159 71.676
R2345 B.n302 B.n160 71.676
R2346 B.n306 B.n161 71.676
R2347 B.n310 B.n162 71.676
R2348 B.n314 B.n163 71.676
R2349 B.n318 B.n164 71.676
R2350 B.n322 B.n165 71.676
R2351 B.n326 B.n166 71.676
R2352 B.n330 B.n167 71.676
R2353 B.n334 B.n168 71.676
R2354 B.n338 B.n169 71.676
R2355 B.n342 B.n170 71.676
R2356 B.n346 B.n171 71.676
R2357 B.n350 B.n172 71.676
R2358 B.n354 B.n173 71.676
R2359 B.n358 B.n174 71.676
R2360 B.n362 B.n175 71.676
R2361 B.n366 B.n176 71.676
R2362 B.n370 B.n177 71.676
R2363 B.n178 B.n177 71.676
R2364 B.n369 B.n176 71.676
R2365 B.n365 B.n175 71.676
R2366 B.n361 B.n174 71.676
R2367 B.n357 B.n173 71.676
R2368 B.n353 B.n172 71.676
R2369 B.n349 B.n171 71.676
R2370 B.n345 B.n170 71.676
R2371 B.n341 B.n169 71.676
R2372 B.n337 B.n168 71.676
R2373 B.n333 B.n167 71.676
R2374 B.n329 B.n166 71.676
R2375 B.n325 B.n165 71.676
R2376 B.n321 B.n164 71.676
R2377 B.n317 B.n163 71.676
R2378 B.n313 B.n162 71.676
R2379 B.n309 B.n161 71.676
R2380 B.n305 B.n160 71.676
R2381 B.n301 B.n159 71.676
R2382 B.n297 B.n158 71.676
R2383 B.n293 B.n157 71.676
R2384 B.n289 B.n156 71.676
R2385 B.n284 B.n155 71.676
R2386 B.n280 B.n154 71.676
R2387 B.n276 B.n153 71.676
R2388 B.n272 B.n152 71.676
R2389 B.n268 B.n151 71.676
R2390 B.n264 B.n150 71.676
R2391 B.n260 B.n149 71.676
R2392 B.n256 B.n148 71.676
R2393 B.n252 B.n147 71.676
R2394 B.n248 B.n146 71.676
R2395 B.n244 B.n145 71.676
R2396 B.n240 B.n144 71.676
R2397 B.n236 B.n143 71.676
R2398 B.n232 B.n142 71.676
R2399 B.n228 B.n141 71.676
R2400 B.n224 B.n140 71.676
R2401 B.n220 B.n139 71.676
R2402 B.n216 B.n138 71.676
R2403 B.n212 B.n137 71.676
R2404 B.n208 B.n136 71.676
R2405 B.n204 B.n135 71.676
R2406 B.n200 B.n134 71.676
R2407 B.n196 B.n133 71.676
R2408 B.n192 B.n132 71.676
R2409 B.n188 B.n131 71.676
R2410 B.n1066 B.n130 71.676
R2411 B.n759 B.n514 71.676
R2412 B.n753 B.n515 71.676
R2413 B.n749 B.n516 71.676
R2414 B.n745 B.n517 71.676
R2415 B.n741 B.n518 71.676
R2416 B.n737 B.n519 71.676
R2417 B.n733 B.n520 71.676
R2418 B.n729 B.n521 71.676
R2419 B.n725 B.n522 71.676
R2420 B.n721 B.n523 71.676
R2421 B.n717 B.n524 71.676
R2422 B.n713 B.n525 71.676
R2423 B.n709 B.n526 71.676
R2424 B.n705 B.n527 71.676
R2425 B.n701 B.n528 71.676
R2426 B.n697 B.n529 71.676
R2427 B.n693 B.n530 71.676
R2428 B.n689 B.n531 71.676
R2429 B.n685 B.n532 71.676
R2430 B.n681 B.n533 71.676
R2431 B.n677 B.n534 71.676
R2432 B.n672 B.n535 71.676
R2433 B.n668 B.n536 71.676
R2434 B.n664 B.n537 71.676
R2435 B.n660 B.n538 71.676
R2436 B.n656 B.n539 71.676
R2437 B.n652 B.n540 71.676
R2438 B.n648 B.n541 71.676
R2439 B.n644 B.n542 71.676
R2440 B.n640 B.n543 71.676
R2441 B.n636 B.n544 71.676
R2442 B.n632 B.n545 71.676
R2443 B.n628 B.n546 71.676
R2444 B.n624 B.n547 71.676
R2445 B.n620 B.n548 71.676
R2446 B.n616 B.n549 71.676
R2447 B.n612 B.n550 71.676
R2448 B.n608 B.n551 71.676
R2449 B.n604 B.n552 71.676
R2450 B.n600 B.n553 71.676
R2451 B.n596 B.n554 71.676
R2452 B.n592 B.n555 71.676
R2453 B.n588 B.n556 71.676
R2454 B.n584 B.n557 71.676
R2455 B.n580 B.n558 71.676
R2456 B.n576 B.n559 71.676
R2457 B.n572 B.n560 71.676
R2458 B.n568 B.n561 71.676
R2459 B.n567 B.n566 59.5399
R2460 B.n674 B.n564 59.5399
R2461 B.n184 B.n183 59.5399
R2462 B.n287 B.n181 59.5399
R2463 B.n765 B.n511 41.5907
R2464 B.n765 B.n507 41.5907
R2465 B.n771 B.n507 41.5907
R2466 B.n771 B.n503 41.5907
R2467 B.n777 B.n503 41.5907
R2468 B.n777 B.n499 41.5907
R2469 B.n783 B.n499 41.5907
R2470 B.n783 B.n495 41.5907
R2471 B.n789 B.n495 41.5907
R2472 B.n795 B.n491 41.5907
R2473 B.n795 B.n487 41.5907
R2474 B.n801 B.n487 41.5907
R2475 B.n801 B.n483 41.5907
R2476 B.n807 B.n483 41.5907
R2477 B.n807 B.n479 41.5907
R2478 B.n813 B.n479 41.5907
R2479 B.n813 B.n475 41.5907
R2480 B.n819 B.n475 41.5907
R2481 B.n819 B.n471 41.5907
R2482 B.n825 B.n471 41.5907
R2483 B.n825 B.n467 41.5907
R2484 B.n831 B.n467 41.5907
R2485 B.n831 B.n463 41.5907
R2486 B.n837 B.n463 41.5907
R2487 B.n843 B.n459 41.5907
R2488 B.n843 B.n455 41.5907
R2489 B.n849 B.n455 41.5907
R2490 B.n849 B.n451 41.5907
R2491 B.n855 B.n451 41.5907
R2492 B.n855 B.n447 41.5907
R2493 B.n861 B.n447 41.5907
R2494 B.n861 B.n443 41.5907
R2495 B.n867 B.n443 41.5907
R2496 B.n867 B.n439 41.5907
R2497 B.n873 B.n439 41.5907
R2498 B.n879 B.n435 41.5907
R2499 B.n879 B.n431 41.5907
R2500 B.n885 B.n431 41.5907
R2501 B.n885 B.n427 41.5907
R2502 B.n891 B.n427 41.5907
R2503 B.n891 B.n423 41.5907
R2504 B.n897 B.n423 41.5907
R2505 B.n897 B.n419 41.5907
R2506 B.n903 B.n419 41.5907
R2507 B.n903 B.n414 41.5907
R2508 B.n909 B.n414 41.5907
R2509 B.n909 B.n415 41.5907
R2510 B.n915 B.n407 41.5907
R2511 B.n921 B.n407 41.5907
R2512 B.n921 B.n403 41.5907
R2513 B.n927 B.n403 41.5907
R2514 B.n927 B.n399 41.5907
R2515 B.n933 B.n399 41.5907
R2516 B.n933 B.n395 41.5907
R2517 B.n939 B.n395 41.5907
R2518 B.n939 B.n391 41.5907
R2519 B.n945 B.n391 41.5907
R2520 B.n945 B.n387 41.5907
R2521 B.n951 B.n387 41.5907
R2522 B.n957 B.n383 41.5907
R2523 B.n957 B.n379 41.5907
R2524 B.n964 B.n379 41.5907
R2525 B.n964 B.n375 41.5907
R2526 B.n970 B.n375 41.5907
R2527 B.n970 B.n4 41.5907
R2528 B.n1210 B.n4 41.5907
R2529 B.n1210 B.n1209 41.5907
R2530 B.n1209 B.n1208 41.5907
R2531 B.n1208 B.n8 41.5907
R2532 B.n1202 B.n8 41.5907
R2533 B.n1202 B.n1201 41.5907
R2534 B.n1201 B.n1200 41.5907
R2535 B.n1200 B.n15 41.5907
R2536 B.n1194 B.n1193 41.5907
R2537 B.n1193 B.n1192 41.5907
R2538 B.n1192 B.n22 41.5907
R2539 B.n1186 B.n22 41.5907
R2540 B.n1186 B.n1185 41.5907
R2541 B.n1185 B.n1184 41.5907
R2542 B.n1184 B.n29 41.5907
R2543 B.n1178 B.n29 41.5907
R2544 B.n1178 B.n1177 41.5907
R2545 B.n1177 B.n1176 41.5907
R2546 B.n1176 B.n36 41.5907
R2547 B.n1170 B.n36 41.5907
R2548 B.n1169 B.n1168 41.5907
R2549 B.n1168 B.n43 41.5907
R2550 B.n1162 B.n43 41.5907
R2551 B.n1162 B.n1161 41.5907
R2552 B.n1161 B.n1160 41.5907
R2553 B.n1160 B.n50 41.5907
R2554 B.n1154 B.n50 41.5907
R2555 B.n1154 B.n1153 41.5907
R2556 B.n1153 B.n1152 41.5907
R2557 B.n1152 B.n57 41.5907
R2558 B.n1146 B.n57 41.5907
R2559 B.n1146 B.n1145 41.5907
R2560 B.n1144 B.n64 41.5907
R2561 B.n1138 B.n64 41.5907
R2562 B.n1138 B.n1137 41.5907
R2563 B.n1137 B.n1136 41.5907
R2564 B.n1136 B.n71 41.5907
R2565 B.n1130 B.n71 41.5907
R2566 B.n1130 B.n1129 41.5907
R2567 B.n1129 B.n1128 41.5907
R2568 B.n1128 B.n78 41.5907
R2569 B.n1122 B.n78 41.5907
R2570 B.n1122 B.n1121 41.5907
R2571 B.n1120 B.n85 41.5907
R2572 B.n1114 B.n85 41.5907
R2573 B.n1114 B.n1113 41.5907
R2574 B.n1113 B.n1112 41.5907
R2575 B.n1112 B.n92 41.5907
R2576 B.n1106 B.n92 41.5907
R2577 B.n1106 B.n1105 41.5907
R2578 B.n1105 B.n1104 41.5907
R2579 B.n1104 B.n99 41.5907
R2580 B.n1098 B.n99 41.5907
R2581 B.n1098 B.n1097 41.5907
R2582 B.n1097 B.n1096 41.5907
R2583 B.n1096 B.n106 41.5907
R2584 B.n1090 B.n106 41.5907
R2585 B.n1090 B.n1089 41.5907
R2586 B.n1088 B.n113 41.5907
R2587 B.n1082 B.n113 41.5907
R2588 B.n1082 B.n1081 41.5907
R2589 B.n1081 B.n1080 41.5907
R2590 B.n1080 B.n120 41.5907
R2591 B.n1074 B.n120 41.5907
R2592 B.n1074 B.n1073 41.5907
R2593 B.n1073 B.n1072 41.5907
R2594 B.n1072 B.n127 41.5907
R2595 B.n873 B.t5 38.5326
R2596 B.t2 B.n1144 38.5326
R2597 B.t4 B.n383 37.3094
R2598 B.t7 B.n15 37.3094
R2599 B.n1069 B.n1068 32.9371
R2600 B.n1063 B.n1062 32.9371
R2601 B.n569 B.n509 32.9371
R2602 B.n762 B.n761 32.9371
R2603 B.t3 B.n459 27.5234
R2604 B.n1121 B.t6 27.5234
R2605 B.n789 B.t9 22.6305
R2606 B.t16 B.n1088 22.6305
R2607 B.n415 B.t0 21.4072
R2608 B.t1 B.n1169 21.4072
R2609 B.n915 B.t0 20.184
R2610 B.n1170 B.t1 20.184
R2611 B.t9 B.n491 18.9607
R2612 B.n1089 B.t16 18.9607
R2613 B B.n1212 18.0485
R2614 B.n837 B.t3 14.0678
R2615 B.t6 B.n1120 14.0678
R2616 B.n1068 B.n129 10.6151
R2617 B.n186 B.n129 10.6151
R2618 B.n187 B.n186 10.6151
R2619 B.n190 B.n187 10.6151
R2620 B.n191 B.n190 10.6151
R2621 B.n194 B.n191 10.6151
R2622 B.n195 B.n194 10.6151
R2623 B.n198 B.n195 10.6151
R2624 B.n199 B.n198 10.6151
R2625 B.n202 B.n199 10.6151
R2626 B.n203 B.n202 10.6151
R2627 B.n206 B.n203 10.6151
R2628 B.n207 B.n206 10.6151
R2629 B.n210 B.n207 10.6151
R2630 B.n211 B.n210 10.6151
R2631 B.n214 B.n211 10.6151
R2632 B.n215 B.n214 10.6151
R2633 B.n218 B.n215 10.6151
R2634 B.n219 B.n218 10.6151
R2635 B.n222 B.n219 10.6151
R2636 B.n223 B.n222 10.6151
R2637 B.n226 B.n223 10.6151
R2638 B.n227 B.n226 10.6151
R2639 B.n230 B.n227 10.6151
R2640 B.n231 B.n230 10.6151
R2641 B.n234 B.n231 10.6151
R2642 B.n235 B.n234 10.6151
R2643 B.n238 B.n235 10.6151
R2644 B.n239 B.n238 10.6151
R2645 B.n242 B.n239 10.6151
R2646 B.n243 B.n242 10.6151
R2647 B.n246 B.n243 10.6151
R2648 B.n247 B.n246 10.6151
R2649 B.n250 B.n247 10.6151
R2650 B.n251 B.n250 10.6151
R2651 B.n254 B.n251 10.6151
R2652 B.n255 B.n254 10.6151
R2653 B.n258 B.n255 10.6151
R2654 B.n259 B.n258 10.6151
R2655 B.n262 B.n259 10.6151
R2656 B.n263 B.n262 10.6151
R2657 B.n266 B.n263 10.6151
R2658 B.n267 B.n266 10.6151
R2659 B.n271 B.n270 10.6151
R2660 B.n274 B.n271 10.6151
R2661 B.n275 B.n274 10.6151
R2662 B.n278 B.n275 10.6151
R2663 B.n279 B.n278 10.6151
R2664 B.n282 B.n279 10.6151
R2665 B.n283 B.n282 10.6151
R2666 B.n286 B.n283 10.6151
R2667 B.n291 B.n288 10.6151
R2668 B.n292 B.n291 10.6151
R2669 B.n295 B.n292 10.6151
R2670 B.n296 B.n295 10.6151
R2671 B.n299 B.n296 10.6151
R2672 B.n300 B.n299 10.6151
R2673 B.n303 B.n300 10.6151
R2674 B.n304 B.n303 10.6151
R2675 B.n307 B.n304 10.6151
R2676 B.n308 B.n307 10.6151
R2677 B.n311 B.n308 10.6151
R2678 B.n312 B.n311 10.6151
R2679 B.n315 B.n312 10.6151
R2680 B.n316 B.n315 10.6151
R2681 B.n319 B.n316 10.6151
R2682 B.n320 B.n319 10.6151
R2683 B.n323 B.n320 10.6151
R2684 B.n324 B.n323 10.6151
R2685 B.n327 B.n324 10.6151
R2686 B.n328 B.n327 10.6151
R2687 B.n331 B.n328 10.6151
R2688 B.n332 B.n331 10.6151
R2689 B.n335 B.n332 10.6151
R2690 B.n336 B.n335 10.6151
R2691 B.n339 B.n336 10.6151
R2692 B.n340 B.n339 10.6151
R2693 B.n343 B.n340 10.6151
R2694 B.n344 B.n343 10.6151
R2695 B.n347 B.n344 10.6151
R2696 B.n348 B.n347 10.6151
R2697 B.n351 B.n348 10.6151
R2698 B.n352 B.n351 10.6151
R2699 B.n355 B.n352 10.6151
R2700 B.n356 B.n355 10.6151
R2701 B.n359 B.n356 10.6151
R2702 B.n360 B.n359 10.6151
R2703 B.n363 B.n360 10.6151
R2704 B.n364 B.n363 10.6151
R2705 B.n367 B.n364 10.6151
R2706 B.n368 B.n367 10.6151
R2707 B.n371 B.n368 10.6151
R2708 B.n372 B.n371 10.6151
R2709 B.n1063 B.n372 10.6151
R2710 B.n767 B.n509 10.6151
R2711 B.n768 B.n767 10.6151
R2712 B.n769 B.n768 10.6151
R2713 B.n769 B.n501 10.6151
R2714 B.n779 B.n501 10.6151
R2715 B.n780 B.n779 10.6151
R2716 B.n781 B.n780 10.6151
R2717 B.n781 B.n493 10.6151
R2718 B.n791 B.n493 10.6151
R2719 B.n792 B.n791 10.6151
R2720 B.n793 B.n792 10.6151
R2721 B.n793 B.n485 10.6151
R2722 B.n803 B.n485 10.6151
R2723 B.n804 B.n803 10.6151
R2724 B.n805 B.n804 10.6151
R2725 B.n805 B.n477 10.6151
R2726 B.n815 B.n477 10.6151
R2727 B.n816 B.n815 10.6151
R2728 B.n817 B.n816 10.6151
R2729 B.n817 B.n469 10.6151
R2730 B.n827 B.n469 10.6151
R2731 B.n828 B.n827 10.6151
R2732 B.n829 B.n828 10.6151
R2733 B.n829 B.n461 10.6151
R2734 B.n839 B.n461 10.6151
R2735 B.n840 B.n839 10.6151
R2736 B.n841 B.n840 10.6151
R2737 B.n841 B.n453 10.6151
R2738 B.n851 B.n453 10.6151
R2739 B.n852 B.n851 10.6151
R2740 B.n853 B.n852 10.6151
R2741 B.n853 B.n445 10.6151
R2742 B.n863 B.n445 10.6151
R2743 B.n864 B.n863 10.6151
R2744 B.n865 B.n864 10.6151
R2745 B.n865 B.n437 10.6151
R2746 B.n875 B.n437 10.6151
R2747 B.n876 B.n875 10.6151
R2748 B.n877 B.n876 10.6151
R2749 B.n877 B.n429 10.6151
R2750 B.n887 B.n429 10.6151
R2751 B.n888 B.n887 10.6151
R2752 B.n889 B.n888 10.6151
R2753 B.n889 B.n421 10.6151
R2754 B.n899 B.n421 10.6151
R2755 B.n900 B.n899 10.6151
R2756 B.n901 B.n900 10.6151
R2757 B.n901 B.n412 10.6151
R2758 B.n911 B.n412 10.6151
R2759 B.n912 B.n911 10.6151
R2760 B.n913 B.n912 10.6151
R2761 B.n913 B.n405 10.6151
R2762 B.n923 B.n405 10.6151
R2763 B.n924 B.n923 10.6151
R2764 B.n925 B.n924 10.6151
R2765 B.n925 B.n397 10.6151
R2766 B.n935 B.n397 10.6151
R2767 B.n936 B.n935 10.6151
R2768 B.n937 B.n936 10.6151
R2769 B.n937 B.n389 10.6151
R2770 B.n947 B.n389 10.6151
R2771 B.n948 B.n947 10.6151
R2772 B.n949 B.n948 10.6151
R2773 B.n949 B.n381 10.6151
R2774 B.n959 B.n381 10.6151
R2775 B.n960 B.n959 10.6151
R2776 B.n962 B.n960 10.6151
R2777 B.n962 B.n961 10.6151
R2778 B.n961 B.n373 10.6151
R2779 B.n973 B.n373 10.6151
R2780 B.n974 B.n973 10.6151
R2781 B.n975 B.n974 10.6151
R2782 B.n976 B.n975 10.6151
R2783 B.n978 B.n976 10.6151
R2784 B.n979 B.n978 10.6151
R2785 B.n980 B.n979 10.6151
R2786 B.n981 B.n980 10.6151
R2787 B.n983 B.n981 10.6151
R2788 B.n984 B.n983 10.6151
R2789 B.n985 B.n984 10.6151
R2790 B.n986 B.n985 10.6151
R2791 B.n988 B.n986 10.6151
R2792 B.n989 B.n988 10.6151
R2793 B.n990 B.n989 10.6151
R2794 B.n991 B.n990 10.6151
R2795 B.n993 B.n991 10.6151
R2796 B.n994 B.n993 10.6151
R2797 B.n995 B.n994 10.6151
R2798 B.n996 B.n995 10.6151
R2799 B.n998 B.n996 10.6151
R2800 B.n999 B.n998 10.6151
R2801 B.n1000 B.n999 10.6151
R2802 B.n1001 B.n1000 10.6151
R2803 B.n1003 B.n1001 10.6151
R2804 B.n1004 B.n1003 10.6151
R2805 B.n1005 B.n1004 10.6151
R2806 B.n1006 B.n1005 10.6151
R2807 B.n1008 B.n1006 10.6151
R2808 B.n1009 B.n1008 10.6151
R2809 B.n1010 B.n1009 10.6151
R2810 B.n1011 B.n1010 10.6151
R2811 B.n1013 B.n1011 10.6151
R2812 B.n1014 B.n1013 10.6151
R2813 B.n1015 B.n1014 10.6151
R2814 B.n1016 B.n1015 10.6151
R2815 B.n1018 B.n1016 10.6151
R2816 B.n1019 B.n1018 10.6151
R2817 B.n1020 B.n1019 10.6151
R2818 B.n1021 B.n1020 10.6151
R2819 B.n1023 B.n1021 10.6151
R2820 B.n1024 B.n1023 10.6151
R2821 B.n1025 B.n1024 10.6151
R2822 B.n1026 B.n1025 10.6151
R2823 B.n1028 B.n1026 10.6151
R2824 B.n1029 B.n1028 10.6151
R2825 B.n1030 B.n1029 10.6151
R2826 B.n1031 B.n1030 10.6151
R2827 B.n1033 B.n1031 10.6151
R2828 B.n1034 B.n1033 10.6151
R2829 B.n1035 B.n1034 10.6151
R2830 B.n1036 B.n1035 10.6151
R2831 B.n1038 B.n1036 10.6151
R2832 B.n1039 B.n1038 10.6151
R2833 B.n1040 B.n1039 10.6151
R2834 B.n1041 B.n1040 10.6151
R2835 B.n1043 B.n1041 10.6151
R2836 B.n1044 B.n1043 10.6151
R2837 B.n1045 B.n1044 10.6151
R2838 B.n1046 B.n1045 10.6151
R2839 B.n1048 B.n1046 10.6151
R2840 B.n1049 B.n1048 10.6151
R2841 B.n1050 B.n1049 10.6151
R2842 B.n1051 B.n1050 10.6151
R2843 B.n1053 B.n1051 10.6151
R2844 B.n1054 B.n1053 10.6151
R2845 B.n1055 B.n1054 10.6151
R2846 B.n1056 B.n1055 10.6151
R2847 B.n1058 B.n1056 10.6151
R2848 B.n1059 B.n1058 10.6151
R2849 B.n1060 B.n1059 10.6151
R2850 B.n1061 B.n1060 10.6151
R2851 B.n1062 B.n1061 10.6151
R2852 B.n761 B.n513 10.6151
R2853 B.n756 B.n513 10.6151
R2854 B.n756 B.n755 10.6151
R2855 B.n755 B.n754 10.6151
R2856 B.n754 B.n751 10.6151
R2857 B.n751 B.n750 10.6151
R2858 B.n750 B.n747 10.6151
R2859 B.n747 B.n746 10.6151
R2860 B.n746 B.n743 10.6151
R2861 B.n743 B.n742 10.6151
R2862 B.n742 B.n739 10.6151
R2863 B.n739 B.n738 10.6151
R2864 B.n738 B.n735 10.6151
R2865 B.n735 B.n734 10.6151
R2866 B.n734 B.n731 10.6151
R2867 B.n731 B.n730 10.6151
R2868 B.n730 B.n727 10.6151
R2869 B.n727 B.n726 10.6151
R2870 B.n726 B.n723 10.6151
R2871 B.n723 B.n722 10.6151
R2872 B.n722 B.n719 10.6151
R2873 B.n719 B.n718 10.6151
R2874 B.n718 B.n715 10.6151
R2875 B.n715 B.n714 10.6151
R2876 B.n714 B.n711 10.6151
R2877 B.n711 B.n710 10.6151
R2878 B.n710 B.n707 10.6151
R2879 B.n707 B.n706 10.6151
R2880 B.n706 B.n703 10.6151
R2881 B.n703 B.n702 10.6151
R2882 B.n702 B.n699 10.6151
R2883 B.n699 B.n698 10.6151
R2884 B.n698 B.n695 10.6151
R2885 B.n695 B.n694 10.6151
R2886 B.n694 B.n691 10.6151
R2887 B.n691 B.n690 10.6151
R2888 B.n690 B.n687 10.6151
R2889 B.n687 B.n686 10.6151
R2890 B.n686 B.n683 10.6151
R2891 B.n683 B.n682 10.6151
R2892 B.n682 B.n679 10.6151
R2893 B.n679 B.n678 10.6151
R2894 B.n678 B.n675 10.6151
R2895 B.n673 B.n670 10.6151
R2896 B.n670 B.n669 10.6151
R2897 B.n669 B.n666 10.6151
R2898 B.n666 B.n665 10.6151
R2899 B.n665 B.n662 10.6151
R2900 B.n662 B.n661 10.6151
R2901 B.n661 B.n658 10.6151
R2902 B.n658 B.n657 10.6151
R2903 B.n654 B.n653 10.6151
R2904 B.n653 B.n650 10.6151
R2905 B.n650 B.n649 10.6151
R2906 B.n649 B.n646 10.6151
R2907 B.n646 B.n645 10.6151
R2908 B.n645 B.n642 10.6151
R2909 B.n642 B.n641 10.6151
R2910 B.n641 B.n638 10.6151
R2911 B.n638 B.n637 10.6151
R2912 B.n637 B.n634 10.6151
R2913 B.n634 B.n633 10.6151
R2914 B.n633 B.n630 10.6151
R2915 B.n630 B.n629 10.6151
R2916 B.n629 B.n626 10.6151
R2917 B.n626 B.n625 10.6151
R2918 B.n625 B.n622 10.6151
R2919 B.n622 B.n621 10.6151
R2920 B.n621 B.n618 10.6151
R2921 B.n618 B.n617 10.6151
R2922 B.n617 B.n614 10.6151
R2923 B.n614 B.n613 10.6151
R2924 B.n613 B.n610 10.6151
R2925 B.n610 B.n609 10.6151
R2926 B.n609 B.n606 10.6151
R2927 B.n606 B.n605 10.6151
R2928 B.n605 B.n602 10.6151
R2929 B.n602 B.n601 10.6151
R2930 B.n601 B.n598 10.6151
R2931 B.n598 B.n597 10.6151
R2932 B.n597 B.n594 10.6151
R2933 B.n594 B.n593 10.6151
R2934 B.n593 B.n590 10.6151
R2935 B.n590 B.n589 10.6151
R2936 B.n589 B.n586 10.6151
R2937 B.n586 B.n585 10.6151
R2938 B.n585 B.n582 10.6151
R2939 B.n582 B.n581 10.6151
R2940 B.n581 B.n578 10.6151
R2941 B.n578 B.n577 10.6151
R2942 B.n577 B.n574 10.6151
R2943 B.n574 B.n573 10.6151
R2944 B.n573 B.n570 10.6151
R2945 B.n570 B.n569 10.6151
R2946 B.n763 B.n762 10.6151
R2947 B.n763 B.n505 10.6151
R2948 B.n773 B.n505 10.6151
R2949 B.n774 B.n773 10.6151
R2950 B.n775 B.n774 10.6151
R2951 B.n775 B.n497 10.6151
R2952 B.n785 B.n497 10.6151
R2953 B.n786 B.n785 10.6151
R2954 B.n787 B.n786 10.6151
R2955 B.n787 B.n489 10.6151
R2956 B.n797 B.n489 10.6151
R2957 B.n798 B.n797 10.6151
R2958 B.n799 B.n798 10.6151
R2959 B.n799 B.n481 10.6151
R2960 B.n809 B.n481 10.6151
R2961 B.n810 B.n809 10.6151
R2962 B.n811 B.n810 10.6151
R2963 B.n811 B.n473 10.6151
R2964 B.n821 B.n473 10.6151
R2965 B.n822 B.n821 10.6151
R2966 B.n823 B.n822 10.6151
R2967 B.n823 B.n465 10.6151
R2968 B.n833 B.n465 10.6151
R2969 B.n834 B.n833 10.6151
R2970 B.n835 B.n834 10.6151
R2971 B.n835 B.n457 10.6151
R2972 B.n845 B.n457 10.6151
R2973 B.n846 B.n845 10.6151
R2974 B.n847 B.n846 10.6151
R2975 B.n847 B.n449 10.6151
R2976 B.n857 B.n449 10.6151
R2977 B.n858 B.n857 10.6151
R2978 B.n859 B.n858 10.6151
R2979 B.n859 B.n441 10.6151
R2980 B.n869 B.n441 10.6151
R2981 B.n870 B.n869 10.6151
R2982 B.n871 B.n870 10.6151
R2983 B.n871 B.n433 10.6151
R2984 B.n881 B.n433 10.6151
R2985 B.n882 B.n881 10.6151
R2986 B.n883 B.n882 10.6151
R2987 B.n883 B.n425 10.6151
R2988 B.n893 B.n425 10.6151
R2989 B.n894 B.n893 10.6151
R2990 B.n895 B.n894 10.6151
R2991 B.n895 B.n417 10.6151
R2992 B.n905 B.n417 10.6151
R2993 B.n906 B.n905 10.6151
R2994 B.n907 B.n906 10.6151
R2995 B.n907 B.n409 10.6151
R2996 B.n917 B.n409 10.6151
R2997 B.n918 B.n917 10.6151
R2998 B.n919 B.n918 10.6151
R2999 B.n919 B.n401 10.6151
R3000 B.n929 B.n401 10.6151
R3001 B.n930 B.n929 10.6151
R3002 B.n931 B.n930 10.6151
R3003 B.n931 B.n393 10.6151
R3004 B.n941 B.n393 10.6151
R3005 B.n942 B.n941 10.6151
R3006 B.n943 B.n942 10.6151
R3007 B.n943 B.n385 10.6151
R3008 B.n953 B.n385 10.6151
R3009 B.n954 B.n953 10.6151
R3010 B.n955 B.n954 10.6151
R3011 B.n955 B.n377 10.6151
R3012 B.n966 B.n377 10.6151
R3013 B.n967 B.n966 10.6151
R3014 B.n968 B.n967 10.6151
R3015 B.n968 B.n0 10.6151
R3016 B.n1206 B.n1 10.6151
R3017 B.n1206 B.n1205 10.6151
R3018 B.n1205 B.n1204 10.6151
R3019 B.n1204 B.n10 10.6151
R3020 B.n1198 B.n10 10.6151
R3021 B.n1198 B.n1197 10.6151
R3022 B.n1197 B.n1196 10.6151
R3023 B.n1196 B.n17 10.6151
R3024 B.n1190 B.n17 10.6151
R3025 B.n1190 B.n1189 10.6151
R3026 B.n1189 B.n1188 10.6151
R3027 B.n1188 B.n24 10.6151
R3028 B.n1182 B.n24 10.6151
R3029 B.n1182 B.n1181 10.6151
R3030 B.n1181 B.n1180 10.6151
R3031 B.n1180 B.n31 10.6151
R3032 B.n1174 B.n31 10.6151
R3033 B.n1174 B.n1173 10.6151
R3034 B.n1173 B.n1172 10.6151
R3035 B.n1172 B.n38 10.6151
R3036 B.n1166 B.n38 10.6151
R3037 B.n1166 B.n1165 10.6151
R3038 B.n1165 B.n1164 10.6151
R3039 B.n1164 B.n45 10.6151
R3040 B.n1158 B.n45 10.6151
R3041 B.n1158 B.n1157 10.6151
R3042 B.n1157 B.n1156 10.6151
R3043 B.n1156 B.n52 10.6151
R3044 B.n1150 B.n52 10.6151
R3045 B.n1150 B.n1149 10.6151
R3046 B.n1149 B.n1148 10.6151
R3047 B.n1148 B.n59 10.6151
R3048 B.n1142 B.n59 10.6151
R3049 B.n1142 B.n1141 10.6151
R3050 B.n1141 B.n1140 10.6151
R3051 B.n1140 B.n66 10.6151
R3052 B.n1134 B.n66 10.6151
R3053 B.n1134 B.n1133 10.6151
R3054 B.n1133 B.n1132 10.6151
R3055 B.n1132 B.n73 10.6151
R3056 B.n1126 B.n73 10.6151
R3057 B.n1126 B.n1125 10.6151
R3058 B.n1125 B.n1124 10.6151
R3059 B.n1124 B.n80 10.6151
R3060 B.n1118 B.n80 10.6151
R3061 B.n1118 B.n1117 10.6151
R3062 B.n1117 B.n1116 10.6151
R3063 B.n1116 B.n87 10.6151
R3064 B.n1110 B.n87 10.6151
R3065 B.n1110 B.n1109 10.6151
R3066 B.n1109 B.n1108 10.6151
R3067 B.n1108 B.n94 10.6151
R3068 B.n1102 B.n94 10.6151
R3069 B.n1102 B.n1101 10.6151
R3070 B.n1101 B.n1100 10.6151
R3071 B.n1100 B.n101 10.6151
R3072 B.n1094 B.n101 10.6151
R3073 B.n1094 B.n1093 10.6151
R3074 B.n1093 B.n1092 10.6151
R3075 B.n1092 B.n108 10.6151
R3076 B.n1086 B.n108 10.6151
R3077 B.n1086 B.n1085 10.6151
R3078 B.n1085 B.n1084 10.6151
R3079 B.n1084 B.n115 10.6151
R3080 B.n1078 B.n115 10.6151
R3081 B.n1078 B.n1077 10.6151
R3082 B.n1077 B.n1076 10.6151
R3083 B.n1076 B.n122 10.6151
R3084 B.n1070 B.n122 10.6151
R3085 B.n1070 B.n1069 10.6151
R3086 B.n270 B.n184 6.5566
R3087 B.n287 B.n286 6.5566
R3088 B.n674 B.n673 6.5566
R3089 B.n657 B.n567 6.5566
R3090 B.n951 B.t4 4.28185
R3091 B.n1194 B.t7 4.28185
R3092 B.n267 B.n184 4.05904
R3093 B.n288 B.n287 4.05904
R3094 B.n675 B.n674 4.05904
R3095 B.n654 B.n567 4.05904
R3096 B.t5 B.n435 3.0586
R3097 B.n1145 B.t2 3.0586
R3098 B.n1212 B.n0 2.81026
R3099 B.n1212 B.n1 2.81026
R3100 VP.n24 VP.n21 161.3
R3101 VP.n26 VP.n25 161.3
R3102 VP.n27 VP.n20 161.3
R3103 VP.n29 VP.n28 161.3
R3104 VP.n30 VP.n19 161.3
R3105 VP.n32 VP.n31 161.3
R3106 VP.n33 VP.n18 161.3
R3107 VP.n35 VP.n34 161.3
R3108 VP.n36 VP.n17 161.3
R3109 VP.n39 VP.n38 161.3
R3110 VP.n40 VP.n16 161.3
R3111 VP.n42 VP.n41 161.3
R3112 VP.n43 VP.n15 161.3
R3113 VP.n45 VP.n44 161.3
R3114 VP.n46 VP.n14 161.3
R3115 VP.n48 VP.n47 161.3
R3116 VP.n49 VP.n13 161.3
R3117 VP.n92 VP.n0 161.3
R3118 VP.n91 VP.n90 161.3
R3119 VP.n89 VP.n1 161.3
R3120 VP.n88 VP.n87 161.3
R3121 VP.n86 VP.n2 161.3
R3122 VP.n85 VP.n84 161.3
R3123 VP.n83 VP.n3 161.3
R3124 VP.n82 VP.n81 161.3
R3125 VP.n79 VP.n4 161.3
R3126 VP.n78 VP.n77 161.3
R3127 VP.n76 VP.n5 161.3
R3128 VP.n75 VP.n74 161.3
R3129 VP.n73 VP.n6 161.3
R3130 VP.n72 VP.n71 161.3
R3131 VP.n70 VP.n7 161.3
R3132 VP.n69 VP.n68 161.3
R3133 VP.n67 VP.n8 161.3
R3134 VP.n65 VP.n64 161.3
R3135 VP.n63 VP.n9 161.3
R3136 VP.n62 VP.n61 161.3
R3137 VP.n60 VP.n10 161.3
R3138 VP.n59 VP.n58 161.3
R3139 VP.n57 VP.n11 161.3
R3140 VP.n56 VP.n55 161.3
R3141 VP.n54 VP.n12 161.3
R3142 VP.n22 VP.t4 109.796
R3143 VP.n53 VP.t5 77.5476
R3144 VP.n66 VP.t3 77.5476
R3145 VP.n80 VP.t0 77.5476
R3146 VP.n93 VP.t7 77.5476
R3147 VP.n50 VP.t2 77.5476
R3148 VP.n37 VP.t1 77.5476
R3149 VP.n23 VP.t6 77.5476
R3150 VP.n23 VP.n22 68.2271
R3151 VP.n53 VP.n52 61.6295
R3152 VP.n94 VP.n93 61.6295
R3153 VP.n51 VP.n50 61.6295
R3154 VP.n52 VP.n51 57.9888
R3155 VP.n60 VP.n59 56.5193
R3156 VP.n87 VP.n86 56.5193
R3157 VP.n44 VP.n43 56.5193
R3158 VP.n73 VP.n72 40.4934
R3159 VP.n74 VP.n73 40.4934
R3160 VP.n31 VP.n30 40.4934
R3161 VP.n30 VP.n29 40.4934
R3162 VP.n55 VP.n54 24.4675
R3163 VP.n55 VP.n11 24.4675
R3164 VP.n59 VP.n11 24.4675
R3165 VP.n61 VP.n60 24.4675
R3166 VP.n61 VP.n9 24.4675
R3167 VP.n65 VP.n9 24.4675
R3168 VP.n68 VP.n67 24.4675
R3169 VP.n68 VP.n7 24.4675
R3170 VP.n72 VP.n7 24.4675
R3171 VP.n74 VP.n5 24.4675
R3172 VP.n78 VP.n5 24.4675
R3173 VP.n79 VP.n78 24.4675
R3174 VP.n81 VP.n3 24.4675
R3175 VP.n85 VP.n3 24.4675
R3176 VP.n86 VP.n85 24.4675
R3177 VP.n87 VP.n1 24.4675
R3178 VP.n91 VP.n1 24.4675
R3179 VP.n92 VP.n91 24.4675
R3180 VP.n44 VP.n14 24.4675
R3181 VP.n48 VP.n14 24.4675
R3182 VP.n49 VP.n48 24.4675
R3183 VP.n31 VP.n18 24.4675
R3184 VP.n35 VP.n18 24.4675
R3185 VP.n36 VP.n35 24.4675
R3186 VP.n38 VP.n16 24.4675
R3187 VP.n42 VP.n16 24.4675
R3188 VP.n43 VP.n42 24.4675
R3189 VP.n25 VP.n24 24.4675
R3190 VP.n25 VP.n20 24.4675
R3191 VP.n29 VP.n20 24.4675
R3192 VP.n54 VP.n53 20.5528
R3193 VP.n93 VP.n92 20.5528
R3194 VP.n50 VP.n49 20.5528
R3195 VP.n66 VP.n65 17.6167
R3196 VP.n81 VP.n80 17.6167
R3197 VP.n38 VP.n37 17.6167
R3198 VP.n67 VP.n66 6.85126
R3199 VP.n80 VP.n79 6.85126
R3200 VP.n37 VP.n36 6.85126
R3201 VP.n24 VP.n23 6.85126
R3202 VP.n22 VP.n21 2.67494
R3203 VP.n51 VP.n13 0.417535
R3204 VP.n52 VP.n12 0.417535
R3205 VP.n94 VP.n0 0.417535
R3206 VP VP.n94 0.394291
R3207 VP.n26 VP.n21 0.189894
R3208 VP.n27 VP.n26 0.189894
R3209 VP.n28 VP.n27 0.189894
R3210 VP.n28 VP.n19 0.189894
R3211 VP.n32 VP.n19 0.189894
R3212 VP.n33 VP.n32 0.189894
R3213 VP.n34 VP.n33 0.189894
R3214 VP.n34 VP.n17 0.189894
R3215 VP.n39 VP.n17 0.189894
R3216 VP.n40 VP.n39 0.189894
R3217 VP.n41 VP.n40 0.189894
R3218 VP.n41 VP.n15 0.189894
R3219 VP.n45 VP.n15 0.189894
R3220 VP.n46 VP.n45 0.189894
R3221 VP.n47 VP.n46 0.189894
R3222 VP.n47 VP.n13 0.189894
R3223 VP.n56 VP.n12 0.189894
R3224 VP.n57 VP.n56 0.189894
R3225 VP.n58 VP.n57 0.189894
R3226 VP.n58 VP.n10 0.189894
R3227 VP.n62 VP.n10 0.189894
R3228 VP.n63 VP.n62 0.189894
R3229 VP.n64 VP.n63 0.189894
R3230 VP.n64 VP.n8 0.189894
R3231 VP.n69 VP.n8 0.189894
R3232 VP.n70 VP.n69 0.189894
R3233 VP.n71 VP.n70 0.189894
R3234 VP.n71 VP.n6 0.189894
R3235 VP.n75 VP.n6 0.189894
R3236 VP.n76 VP.n75 0.189894
R3237 VP.n77 VP.n76 0.189894
R3238 VP.n77 VP.n4 0.189894
R3239 VP.n82 VP.n4 0.189894
R3240 VP.n83 VP.n82 0.189894
R3241 VP.n84 VP.n83 0.189894
R3242 VP.n84 VP.n2 0.189894
R3243 VP.n88 VP.n2 0.189894
R3244 VP.n89 VP.n88 0.189894
R3245 VP.n90 VP.n89 0.189894
R3246 VP.n90 VP.n0 0.189894
R3247 VDD1 VDD1.n0 67.5721
R3248 VDD1.n3 VDD1.n2 67.4575
R3249 VDD1.n3 VDD1.n1 67.4575
R3250 VDD1.n5 VDD1.n4 65.668
R3251 VDD1.n5 VDD1.n3 51.8587
R3252 VDD1 VDD1.n5 1.78714
R3253 VDD1.n4 VDD1.t6 1.55833
R3254 VDD1.n4 VDD1.t5 1.55833
R3255 VDD1.n0 VDD1.t3 1.55833
R3256 VDD1.n0 VDD1.t1 1.55833
R3257 VDD1.n2 VDD1.t7 1.55833
R3258 VDD1.n2 VDD1.t0 1.55833
R3259 VDD1.n1 VDD1.t2 1.55833
R3260 VDD1.n1 VDD1.t4 1.55833
C0 VDD2 VP 0.663478f
C1 VN VTAIL 10.6476f
C2 VP VN 9.44842f
C3 VP VTAIL 10.6617f
C4 VDD1 VDD2 2.47962f
C5 VDD1 VN 0.154322f
C6 VDD2 VN 9.82425f
C7 VDD1 VTAIL 8.893041f
C8 VDD1 VP 10.3313f
C9 VDD2 VTAIL 8.95651f
C10 VDD2 B 6.80772f
C11 VDD1 B 7.38995f
C12 VTAIL B 11.810697f
C13 VN B 20.79114f
C14 VP B 19.45867f
C15 VDD1.t3 B 0.277218f
C16 VDD1.t1 B 0.277218f
C17 VDD1.n0 B 2.51054f
C18 VDD1.t2 B 0.277218f
C19 VDD1.t4 B 0.277218f
C20 VDD1.n1 B 2.50909f
C21 VDD1.t7 B 0.277218f
C22 VDD1.t0 B 0.277218f
C23 VDD1.n2 B 2.50909f
C24 VDD1.n3 B 4.57002f
C25 VDD1.t6 B 0.277218f
C26 VDD1.t5 B 0.277218f
C27 VDD1.n4 B 2.49007f
C28 VDD1.n5 B 3.85932f
C29 VP.n0 B 0.031961f
C30 VP.t7 B 2.32796f
C31 VP.n1 B 0.031668f
C32 VP.n2 B 0.016992f
C33 VP.n3 B 0.031668f
C34 VP.n4 B 0.016992f
C35 VP.t0 B 2.32796f
C36 VP.n5 B 0.031668f
C37 VP.n6 B 0.016992f
C38 VP.n7 B 0.031668f
C39 VP.n8 B 0.016992f
C40 VP.t3 B 2.32796f
C41 VP.n9 B 0.031668f
C42 VP.n10 B 0.016992f
C43 VP.n11 B 0.031668f
C44 VP.n12 B 0.031961f
C45 VP.t5 B 2.32796f
C46 VP.n13 B 0.031961f
C47 VP.t2 B 2.32796f
C48 VP.n14 B 0.031668f
C49 VP.n15 B 0.016992f
C50 VP.n16 B 0.031668f
C51 VP.n17 B 0.016992f
C52 VP.t1 B 2.32796f
C53 VP.n18 B 0.031668f
C54 VP.n19 B 0.016992f
C55 VP.n20 B 0.031668f
C56 VP.n21 B 0.225959f
C57 VP.t6 B 2.32796f
C58 VP.t4 B 2.60596f
C59 VP.n22 B 0.829274f
C60 VP.n23 B 0.871073f
C61 VP.n24 B 0.020411f
C62 VP.n25 B 0.031668f
C63 VP.n26 B 0.016992f
C64 VP.n27 B 0.016992f
C65 VP.n28 B 0.016992f
C66 VP.n29 B 0.033771f
C67 VP.n30 B 0.013736f
C68 VP.n31 B 0.033771f
C69 VP.n32 B 0.016992f
C70 VP.n33 B 0.016992f
C71 VP.n34 B 0.016992f
C72 VP.n35 B 0.031668f
C73 VP.n36 B 0.020411f
C74 VP.n37 B 0.812519f
C75 VP.n38 B 0.02729f
C76 VP.n39 B 0.016992f
C77 VP.n40 B 0.016992f
C78 VP.n41 B 0.016992f
C79 VP.n42 B 0.031668f
C80 VP.n43 B 0.026225f
C81 VP.n44 B 0.023384f
C82 VP.n45 B 0.016992f
C83 VP.n46 B 0.016992f
C84 VP.n47 B 0.016992f
C85 VP.n48 B 0.031668f
C86 VP.n49 B 0.029166f
C87 VP.n50 B 0.887101f
C88 VP.n51 B 1.21064f
C89 VP.n52 B 1.22117f
C90 VP.n53 B 0.887101f
C91 VP.n54 B 0.029166f
C92 VP.n55 B 0.031668f
C93 VP.n56 B 0.016992f
C94 VP.n57 B 0.016992f
C95 VP.n58 B 0.016992f
C96 VP.n59 B 0.023384f
C97 VP.n60 B 0.026225f
C98 VP.n61 B 0.031668f
C99 VP.n62 B 0.016992f
C100 VP.n63 B 0.016992f
C101 VP.n64 B 0.016992f
C102 VP.n65 B 0.02729f
C103 VP.n66 B 0.812519f
C104 VP.n67 B 0.020411f
C105 VP.n68 B 0.031668f
C106 VP.n69 B 0.016992f
C107 VP.n70 B 0.016992f
C108 VP.n71 B 0.016992f
C109 VP.n72 B 0.033771f
C110 VP.n73 B 0.013736f
C111 VP.n74 B 0.033771f
C112 VP.n75 B 0.016992f
C113 VP.n76 B 0.016992f
C114 VP.n77 B 0.016992f
C115 VP.n78 B 0.031668f
C116 VP.n79 B 0.020411f
C117 VP.n80 B 0.812519f
C118 VP.n81 B 0.02729f
C119 VP.n82 B 0.016992f
C120 VP.n83 B 0.016992f
C121 VP.n84 B 0.016992f
C122 VP.n85 B 0.031668f
C123 VP.n86 B 0.026225f
C124 VP.n87 B 0.023384f
C125 VP.n88 B 0.016992f
C126 VP.n89 B 0.016992f
C127 VP.n90 B 0.016992f
C128 VP.n91 B 0.031668f
C129 VP.n92 B 0.029166f
C130 VP.n93 B 0.887101f
C131 VP.n94 B 0.053691f
C132 VTAIL.t8 B 0.207228f
C133 VTAIL.t14 B 0.207228f
C134 VTAIL.n0 B 1.80729f
C135 VTAIL.n1 B 0.438142f
C136 VTAIL.n2 B 0.011647f
C137 VTAIL.n3 B 0.026206f
C138 VTAIL.n4 B 0.011739f
C139 VTAIL.n5 B 0.020632f
C140 VTAIL.n6 B 0.011087f
C141 VTAIL.n7 B 0.026206f
C142 VTAIL.n8 B 0.011739f
C143 VTAIL.n9 B 0.020632f
C144 VTAIL.n10 B 0.011087f
C145 VTAIL.n11 B 0.026206f
C146 VTAIL.n12 B 0.011739f
C147 VTAIL.n13 B 0.020632f
C148 VTAIL.n14 B 0.011087f
C149 VTAIL.n15 B 0.026206f
C150 VTAIL.n16 B 0.011739f
C151 VTAIL.n17 B 0.020632f
C152 VTAIL.n18 B 0.011087f
C153 VTAIL.n19 B 0.026206f
C154 VTAIL.n20 B 0.011739f
C155 VTAIL.n21 B 0.020632f
C156 VTAIL.n22 B 0.011087f
C157 VTAIL.n23 B 0.019654f
C158 VTAIL.n24 B 0.01548f
C159 VTAIL.t11 B 0.043048f
C160 VTAIL.n25 B 0.122723f
C161 VTAIL.n26 B 1.12583f
C162 VTAIL.n27 B 0.011087f
C163 VTAIL.n28 B 0.011739f
C164 VTAIL.n29 B 0.026206f
C165 VTAIL.n30 B 0.026206f
C166 VTAIL.n31 B 0.011739f
C167 VTAIL.n32 B 0.011087f
C168 VTAIL.n33 B 0.020632f
C169 VTAIL.n34 B 0.020632f
C170 VTAIL.n35 B 0.011087f
C171 VTAIL.n36 B 0.011739f
C172 VTAIL.n37 B 0.026206f
C173 VTAIL.n38 B 0.026206f
C174 VTAIL.n39 B 0.011739f
C175 VTAIL.n40 B 0.011087f
C176 VTAIL.n41 B 0.020632f
C177 VTAIL.n42 B 0.020632f
C178 VTAIL.n43 B 0.011087f
C179 VTAIL.n44 B 0.011739f
C180 VTAIL.n45 B 0.026206f
C181 VTAIL.n46 B 0.026206f
C182 VTAIL.n47 B 0.011739f
C183 VTAIL.n48 B 0.011087f
C184 VTAIL.n49 B 0.020632f
C185 VTAIL.n50 B 0.020632f
C186 VTAIL.n51 B 0.011087f
C187 VTAIL.n52 B 0.011739f
C188 VTAIL.n53 B 0.026206f
C189 VTAIL.n54 B 0.026206f
C190 VTAIL.n55 B 0.011739f
C191 VTAIL.n56 B 0.011087f
C192 VTAIL.n57 B 0.020632f
C193 VTAIL.n58 B 0.020632f
C194 VTAIL.n59 B 0.011087f
C195 VTAIL.n60 B 0.011739f
C196 VTAIL.n61 B 0.026206f
C197 VTAIL.n62 B 0.026206f
C198 VTAIL.n63 B 0.011739f
C199 VTAIL.n64 B 0.011087f
C200 VTAIL.n65 B 0.020632f
C201 VTAIL.n66 B 0.054173f
C202 VTAIL.n67 B 0.011087f
C203 VTAIL.n68 B 0.011739f
C204 VTAIL.n69 B 0.054515f
C205 VTAIL.n70 B 0.046233f
C206 VTAIL.n71 B 0.297503f
C207 VTAIL.n72 B 0.011647f
C208 VTAIL.n73 B 0.026206f
C209 VTAIL.n74 B 0.011739f
C210 VTAIL.n75 B 0.020632f
C211 VTAIL.n76 B 0.011087f
C212 VTAIL.n77 B 0.026206f
C213 VTAIL.n78 B 0.011739f
C214 VTAIL.n79 B 0.020632f
C215 VTAIL.n80 B 0.011087f
C216 VTAIL.n81 B 0.026206f
C217 VTAIL.n82 B 0.011739f
C218 VTAIL.n83 B 0.020632f
C219 VTAIL.n84 B 0.011087f
C220 VTAIL.n85 B 0.026206f
C221 VTAIL.n86 B 0.011739f
C222 VTAIL.n87 B 0.020632f
C223 VTAIL.n88 B 0.011087f
C224 VTAIL.n89 B 0.026206f
C225 VTAIL.n90 B 0.011739f
C226 VTAIL.n91 B 0.020632f
C227 VTAIL.n92 B 0.011087f
C228 VTAIL.n93 B 0.019654f
C229 VTAIL.n94 B 0.01548f
C230 VTAIL.t4 B 0.043048f
C231 VTAIL.n95 B 0.122723f
C232 VTAIL.n96 B 1.12583f
C233 VTAIL.n97 B 0.011087f
C234 VTAIL.n98 B 0.011739f
C235 VTAIL.n99 B 0.026206f
C236 VTAIL.n100 B 0.026206f
C237 VTAIL.n101 B 0.011739f
C238 VTAIL.n102 B 0.011087f
C239 VTAIL.n103 B 0.020632f
C240 VTAIL.n104 B 0.020632f
C241 VTAIL.n105 B 0.011087f
C242 VTAIL.n106 B 0.011739f
C243 VTAIL.n107 B 0.026206f
C244 VTAIL.n108 B 0.026206f
C245 VTAIL.n109 B 0.011739f
C246 VTAIL.n110 B 0.011087f
C247 VTAIL.n111 B 0.020632f
C248 VTAIL.n112 B 0.020632f
C249 VTAIL.n113 B 0.011087f
C250 VTAIL.n114 B 0.011739f
C251 VTAIL.n115 B 0.026206f
C252 VTAIL.n116 B 0.026206f
C253 VTAIL.n117 B 0.011739f
C254 VTAIL.n118 B 0.011087f
C255 VTAIL.n119 B 0.020632f
C256 VTAIL.n120 B 0.020632f
C257 VTAIL.n121 B 0.011087f
C258 VTAIL.n122 B 0.011739f
C259 VTAIL.n123 B 0.026206f
C260 VTAIL.n124 B 0.026206f
C261 VTAIL.n125 B 0.011739f
C262 VTAIL.n126 B 0.011087f
C263 VTAIL.n127 B 0.020632f
C264 VTAIL.n128 B 0.020632f
C265 VTAIL.n129 B 0.011087f
C266 VTAIL.n130 B 0.011739f
C267 VTAIL.n131 B 0.026206f
C268 VTAIL.n132 B 0.026206f
C269 VTAIL.n133 B 0.011739f
C270 VTAIL.n134 B 0.011087f
C271 VTAIL.n135 B 0.020632f
C272 VTAIL.n136 B 0.054173f
C273 VTAIL.n137 B 0.011087f
C274 VTAIL.n138 B 0.011739f
C275 VTAIL.n139 B 0.054515f
C276 VTAIL.n140 B 0.046233f
C277 VTAIL.n141 B 0.297503f
C278 VTAIL.t5 B 0.207228f
C279 VTAIL.t0 B 0.207228f
C280 VTAIL.n142 B 1.80729f
C281 VTAIL.n143 B 0.67957f
C282 VTAIL.n144 B 0.011647f
C283 VTAIL.n145 B 0.026206f
C284 VTAIL.n146 B 0.011739f
C285 VTAIL.n147 B 0.020632f
C286 VTAIL.n148 B 0.011087f
C287 VTAIL.n149 B 0.026206f
C288 VTAIL.n150 B 0.011739f
C289 VTAIL.n151 B 0.020632f
C290 VTAIL.n152 B 0.011087f
C291 VTAIL.n153 B 0.026206f
C292 VTAIL.n154 B 0.011739f
C293 VTAIL.n155 B 0.020632f
C294 VTAIL.n156 B 0.011087f
C295 VTAIL.n157 B 0.026206f
C296 VTAIL.n158 B 0.011739f
C297 VTAIL.n159 B 0.020632f
C298 VTAIL.n160 B 0.011087f
C299 VTAIL.n161 B 0.026206f
C300 VTAIL.n162 B 0.011739f
C301 VTAIL.n163 B 0.020632f
C302 VTAIL.n164 B 0.011087f
C303 VTAIL.n165 B 0.019654f
C304 VTAIL.n166 B 0.01548f
C305 VTAIL.t3 B 0.043048f
C306 VTAIL.n167 B 0.122723f
C307 VTAIL.n168 B 1.12583f
C308 VTAIL.n169 B 0.011087f
C309 VTAIL.n170 B 0.011739f
C310 VTAIL.n171 B 0.026206f
C311 VTAIL.n172 B 0.026206f
C312 VTAIL.n173 B 0.011739f
C313 VTAIL.n174 B 0.011087f
C314 VTAIL.n175 B 0.020632f
C315 VTAIL.n176 B 0.020632f
C316 VTAIL.n177 B 0.011087f
C317 VTAIL.n178 B 0.011739f
C318 VTAIL.n179 B 0.026206f
C319 VTAIL.n180 B 0.026206f
C320 VTAIL.n181 B 0.011739f
C321 VTAIL.n182 B 0.011087f
C322 VTAIL.n183 B 0.020632f
C323 VTAIL.n184 B 0.020632f
C324 VTAIL.n185 B 0.011087f
C325 VTAIL.n186 B 0.011739f
C326 VTAIL.n187 B 0.026206f
C327 VTAIL.n188 B 0.026206f
C328 VTAIL.n189 B 0.011739f
C329 VTAIL.n190 B 0.011087f
C330 VTAIL.n191 B 0.020632f
C331 VTAIL.n192 B 0.020632f
C332 VTAIL.n193 B 0.011087f
C333 VTAIL.n194 B 0.011739f
C334 VTAIL.n195 B 0.026206f
C335 VTAIL.n196 B 0.026206f
C336 VTAIL.n197 B 0.011739f
C337 VTAIL.n198 B 0.011087f
C338 VTAIL.n199 B 0.020632f
C339 VTAIL.n200 B 0.020632f
C340 VTAIL.n201 B 0.011087f
C341 VTAIL.n202 B 0.011739f
C342 VTAIL.n203 B 0.026206f
C343 VTAIL.n204 B 0.026206f
C344 VTAIL.n205 B 0.011739f
C345 VTAIL.n206 B 0.011087f
C346 VTAIL.n207 B 0.020632f
C347 VTAIL.n208 B 0.054173f
C348 VTAIL.n209 B 0.011087f
C349 VTAIL.n210 B 0.011739f
C350 VTAIL.n211 B 0.054515f
C351 VTAIL.n212 B 0.046233f
C352 VTAIL.n213 B 1.52027f
C353 VTAIL.n214 B 0.011647f
C354 VTAIL.n215 B 0.026206f
C355 VTAIL.n216 B 0.011739f
C356 VTAIL.n217 B 0.020632f
C357 VTAIL.n218 B 0.011087f
C358 VTAIL.n219 B 0.026206f
C359 VTAIL.n220 B 0.011739f
C360 VTAIL.n221 B 0.020632f
C361 VTAIL.n222 B 0.011087f
C362 VTAIL.n223 B 0.026206f
C363 VTAIL.n224 B 0.011739f
C364 VTAIL.n225 B 0.020632f
C365 VTAIL.n226 B 0.011087f
C366 VTAIL.n227 B 0.026206f
C367 VTAIL.n228 B 0.011739f
C368 VTAIL.n229 B 0.020632f
C369 VTAIL.n230 B 0.011087f
C370 VTAIL.n231 B 0.026206f
C371 VTAIL.n232 B 0.011739f
C372 VTAIL.n233 B 0.020632f
C373 VTAIL.n234 B 0.011087f
C374 VTAIL.n235 B 0.019654f
C375 VTAIL.n236 B 0.01548f
C376 VTAIL.t13 B 0.043048f
C377 VTAIL.n237 B 0.122723f
C378 VTAIL.n238 B 1.12583f
C379 VTAIL.n239 B 0.011087f
C380 VTAIL.n240 B 0.011739f
C381 VTAIL.n241 B 0.026206f
C382 VTAIL.n242 B 0.026206f
C383 VTAIL.n243 B 0.011739f
C384 VTAIL.n244 B 0.011087f
C385 VTAIL.n245 B 0.020632f
C386 VTAIL.n246 B 0.020632f
C387 VTAIL.n247 B 0.011087f
C388 VTAIL.n248 B 0.011739f
C389 VTAIL.n249 B 0.026206f
C390 VTAIL.n250 B 0.026206f
C391 VTAIL.n251 B 0.011739f
C392 VTAIL.n252 B 0.011087f
C393 VTAIL.n253 B 0.020632f
C394 VTAIL.n254 B 0.020632f
C395 VTAIL.n255 B 0.011087f
C396 VTAIL.n256 B 0.011739f
C397 VTAIL.n257 B 0.026206f
C398 VTAIL.n258 B 0.026206f
C399 VTAIL.n259 B 0.011739f
C400 VTAIL.n260 B 0.011087f
C401 VTAIL.n261 B 0.020632f
C402 VTAIL.n262 B 0.020632f
C403 VTAIL.n263 B 0.011087f
C404 VTAIL.n264 B 0.011739f
C405 VTAIL.n265 B 0.026206f
C406 VTAIL.n266 B 0.026206f
C407 VTAIL.n267 B 0.011739f
C408 VTAIL.n268 B 0.011087f
C409 VTAIL.n269 B 0.020632f
C410 VTAIL.n270 B 0.020632f
C411 VTAIL.n271 B 0.011087f
C412 VTAIL.n272 B 0.011739f
C413 VTAIL.n273 B 0.026206f
C414 VTAIL.n274 B 0.026206f
C415 VTAIL.n275 B 0.011739f
C416 VTAIL.n276 B 0.011087f
C417 VTAIL.n277 B 0.020632f
C418 VTAIL.n278 B 0.054173f
C419 VTAIL.n279 B 0.011087f
C420 VTAIL.n280 B 0.011739f
C421 VTAIL.n281 B 0.054515f
C422 VTAIL.n282 B 0.046233f
C423 VTAIL.n283 B 1.52027f
C424 VTAIL.t9 B 0.207228f
C425 VTAIL.t15 B 0.207228f
C426 VTAIL.n284 B 1.80728f
C427 VTAIL.n285 B 0.679575f
C428 VTAIL.n286 B 0.011647f
C429 VTAIL.n287 B 0.026206f
C430 VTAIL.n288 B 0.011739f
C431 VTAIL.n289 B 0.020632f
C432 VTAIL.n290 B 0.011087f
C433 VTAIL.n291 B 0.026206f
C434 VTAIL.n292 B 0.011739f
C435 VTAIL.n293 B 0.020632f
C436 VTAIL.n294 B 0.011087f
C437 VTAIL.n295 B 0.026206f
C438 VTAIL.n296 B 0.011739f
C439 VTAIL.n297 B 0.020632f
C440 VTAIL.n298 B 0.011087f
C441 VTAIL.n299 B 0.026206f
C442 VTAIL.n300 B 0.011739f
C443 VTAIL.n301 B 0.020632f
C444 VTAIL.n302 B 0.011087f
C445 VTAIL.n303 B 0.026206f
C446 VTAIL.n304 B 0.011739f
C447 VTAIL.n305 B 0.020632f
C448 VTAIL.n306 B 0.011087f
C449 VTAIL.n307 B 0.019654f
C450 VTAIL.n308 B 0.01548f
C451 VTAIL.t10 B 0.043048f
C452 VTAIL.n309 B 0.122723f
C453 VTAIL.n310 B 1.12583f
C454 VTAIL.n311 B 0.011087f
C455 VTAIL.n312 B 0.011739f
C456 VTAIL.n313 B 0.026206f
C457 VTAIL.n314 B 0.026206f
C458 VTAIL.n315 B 0.011739f
C459 VTAIL.n316 B 0.011087f
C460 VTAIL.n317 B 0.020632f
C461 VTAIL.n318 B 0.020632f
C462 VTAIL.n319 B 0.011087f
C463 VTAIL.n320 B 0.011739f
C464 VTAIL.n321 B 0.026206f
C465 VTAIL.n322 B 0.026206f
C466 VTAIL.n323 B 0.011739f
C467 VTAIL.n324 B 0.011087f
C468 VTAIL.n325 B 0.020632f
C469 VTAIL.n326 B 0.020632f
C470 VTAIL.n327 B 0.011087f
C471 VTAIL.n328 B 0.011739f
C472 VTAIL.n329 B 0.026206f
C473 VTAIL.n330 B 0.026206f
C474 VTAIL.n331 B 0.011739f
C475 VTAIL.n332 B 0.011087f
C476 VTAIL.n333 B 0.020632f
C477 VTAIL.n334 B 0.020632f
C478 VTAIL.n335 B 0.011087f
C479 VTAIL.n336 B 0.011739f
C480 VTAIL.n337 B 0.026206f
C481 VTAIL.n338 B 0.026206f
C482 VTAIL.n339 B 0.011739f
C483 VTAIL.n340 B 0.011087f
C484 VTAIL.n341 B 0.020632f
C485 VTAIL.n342 B 0.020632f
C486 VTAIL.n343 B 0.011087f
C487 VTAIL.n344 B 0.011739f
C488 VTAIL.n345 B 0.026206f
C489 VTAIL.n346 B 0.026206f
C490 VTAIL.n347 B 0.011739f
C491 VTAIL.n348 B 0.011087f
C492 VTAIL.n349 B 0.020632f
C493 VTAIL.n350 B 0.054173f
C494 VTAIL.n351 B 0.011087f
C495 VTAIL.n352 B 0.011739f
C496 VTAIL.n353 B 0.054515f
C497 VTAIL.n354 B 0.046233f
C498 VTAIL.n355 B 0.297503f
C499 VTAIL.n356 B 0.011647f
C500 VTAIL.n357 B 0.026206f
C501 VTAIL.n358 B 0.011739f
C502 VTAIL.n359 B 0.020632f
C503 VTAIL.n360 B 0.011087f
C504 VTAIL.n361 B 0.026206f
C505 VTAIL.n362 B 0.011739f
C506 VTAIL.n363 B 0.020632f
C507 VTAIL.n364 B 0.011087f
C508 VTAIL.n365 B 0.026206f
C509 VTAIL.n366 B 0.011739f
C510 VTAIL.n367 B 0.020632f
C511 VTAIL.n368 B 0.011087f
C512 VTAIL.n369 B 0.026206f
C513 VTAIL.n370 B 0.011739f
C514 VTAIL.n371 B 0.020632f
C515 VTAIL.n372 B 0.011087f
C516 VTAIL.n373 B 0.026206f
C517 VTAIL.n374 B 0.011739f
C518 VTAIL.n375 B 0.020632f
C519 VTAIL.n376 B 0.011087f
C520 VTAIL.n377 B 0.019654f
C521 VTAIL.n378 B 0.01548f
C522 VTAIL.t7 B 0.043048f
C523 VTAIL.n379 B 0.122723f
C524 VTAIL.n380 B 1.12583f
C525 VTAIL.n381 B 0.011087f
C526 VTAIL.n382 B 0.011739f
C527 VTAIL.n383 B 0.026206f
C528 VTAIL.n384 B 0.026206f
C529 VTAIL.n385 B 0.011739f
C530 VTAIL.n386 B 0.011087f
C531 VTAIL.n387 B 0.020632f
C532 VTAIL.n388 B 0.020632f
C533 VTAIL.n389 B 0.011087f
C534 VTAIL.n390 B 0.011739f
C535 VTAIL.n391 B 0.026206f
C536 VTAIL.n392 B 0.026206f
C537 VTAIL.n393 B 0.011739f
C538 VTAIL.n394 B 0.011087f
C539 VTAIL.n395 B 0.020632f
C540 VTAIL.n396 B 0.020632f
C541 VTAIL.n397 B 0.011087f
C542 VTAIL.n398 B 0.011739f
C543 VTAIL.n399 B 0.026206f
C544 VTAIL.n400 B 0.026206f
C545 VTAIL.n401 B 0.011739f
C546 VTAIL.n402 B 0.011087f
C547 VTAIL.n403 B 0.020632f
C548 VTAIL.n404 B 0.020632f
C549 VTAIL.n405 B 0.011087f
C550 VTAIL.n406 B 0.011739f
C551 VTAIL.n407 B 0.026206f
C552 VTAIL.n408 B 0.026206f
C553 VTAIL.n409 B 0.011739f
C554 VTAIL.n410 B 0.011087f
C555 VTAIL.n411 B 0.020632f
C556 VTAIL.n412 B 0.020632f
C557 VTAIL.n413 B 0.011087f
C558 VTAIL.n414 B 0.011739f
C559 VTAIL.n415 B 0.026206f
C560 VTAIL.n416 B 0.026206f
C561 VTAIL.n417 B 0.011739f
C562 VTAIL.n418 B 0.011087f
C563 VTAIL.n419 B 0.020632f
C564 VTAIL.n420 B 0.054173f
C565 VTAIL.n421 B 0.011087f
C566 VTAIL.n422 B 0.011739f
C567 VTAIL.n423 B 0.054515f
C568 VTAIL.n424 B 0.046233f
C569 VTAIL.n425 B 0.297503f
C570 VTAIL.t1 B 0.207228f
C571 VTAIL.t2 B 0.207228f
C572 VTAIL.n426 B 1.80728f
C573 VTAIL.n427 B 0.679575f
C574 VTAIL.n428 B 0.011647f
C575 VTAIL.n429 B 0.026206f
C576 VTAIL.n430 B 0.011739f
C577 VTAIL.n431 B 0.020632f
C578 VTAIL.n432 B 0.011087f
C579 VTAIL.n433 B 0.026206f
C580 VTAIL.n434 B 0.011739f
C581 VTAIL.n435 B 0.020632f
C582 VTAIL.n436 B 0.011087f
C583 VTAIL.n437 B 0.026206f
C584 VTAIL.n438 B 0.011739f
C585 VTAIL.n439 B 0.020632f
C586 VTAIL.n440 B 0.011087f
C587 VTAIL.n441 B 0.026206f
C588 VTAIL.n442 B 0.011739f
C589 VTAIL.n443 B 0.020632f
C590 VTAIL.n444 B 0.011087f
C591 VTAIL.n445 B 0.026206f
C592 VTAIL.n446 B 0.011739f
C593 VTAIL.n447 B 0.020632f
C594 VTAIL.n448 B 0.011087f
C595 VTAIL.n449 B 0.019654f
C596 VTAIL.n450 B 0.01548f
C597 VTAIL.t6 B 0.043048f
C598 VTAIL.n451 B 0.122723f
C599 VTAIL.n452 B 1.12583f
C600 VTAIL.n453 B 0.011087f
C601 VTAIL.n454 B 0.011739f
C602 VTAIL.n455 B 0.026206f
C603 VTAIL.n456 B 0.026206f
C604 VTAIL.n457 B 0.011739f
C605 VTAIL.n458 B 0.011087f
C606 VTAIL.n459 B 0.020632f
C607 VTAIL.n460 B 0.020632f
C608 VTAIL.n461 B 0.011087f
C609 VTAIL.n462 B 0.011739f
C610 VTAIL.n463 B 0.026206f
C611 VTAIL.n464 B 0.026206f
C612 VTAIL.n465 B 0.011739f
C613 VTAIL.n466 B 0.011087f
C614 VTAIL.n467 B 0.020632f
C615 VTAIL.n468 B 0.020632f
C616 VTAIL.n469 B 0.011087f
C617 VTAIL.n470 B 0.011739f
C618 VTAIL.n471 B 0.026206f
C619 VTAIL.n472 B 0.026206f
C620 VTAIL.n473 B 0.011739f
C621 VTAIL.n474 B 0.011087f
C622 VTAIL.n475 B 0.020632f
C623 VTAIL.n476 B 0.020632f
C624 VTAIL.n477 B 0.011087f
C625 VTAIL.n478 B 0.011739f
C626 VTAIL.n479 B 0.026206f
C627 VTAIL.n480 B 0.026206f
C628 VTAIL.n481 B 0.011739f
C629 VTAIL.n482 B 0.011087f
C630 VTAIL.n483 B 0.020632f
C631 VTAIL.n484 B 0.020632f
C632 VTAIL.n485 B 0.011087f
C633 VTAIL.n486 B 0.011739f
C634 VTAIL.n487 B 0.026206f
C635 VTAIL.n488 B 0.026206f
C636 VTAIL.n489 B 0.011739f
C637 VTAIL.n490 B 0.011087f
C638 VTAIL.n491 B 0.020632f
C639 VTAIL.n492 B 0.054173f
C640 VTAIL.n493 B 0.011087f
C641 VTAIL.n494 B 0.011739f
C642 VTAIL.n495 B 0.054515f
C643 VTAIL.n496 B 0.046233f
C644 VTAIL.n497 B 1.52027f
C645 VTAIL.n498 B 0.011647f
C646 VTAIL.n499 B 0.026206f
C647 VTAIL.n500 B 0.011739f
C648 VTAIL.n501 B 0.020632f
C649 VTAIL.n502 B 0.011087f
C650 VTAIL.n503 B 0.026206f
C651 VTAIL.n504 B 0.011739f
C652 VTAIL.n505 B 0.020632f
C653 VTAIL.n506 B 0.011087f
C654 VTAIL.n507 B 0.026206f
C655 VTAIL.n508 B 0.011739f
C656 VTAIL.n509 B 0.020632f
C657 VTAIL.n510 B 0.011087f
C658 VTAIL.n511 B 0.026206f
C659 VTAIL.n512 B 0.011739f
C660 VTAIL.n513 B 0.020632f
C661 VTAIL.n514 B 0.011087f
C662 VTAIL.n515 B 0.026206f
C663 VTAIL.n516 B 0.011739f
C664 VTAIL.n517 B 0.020632f
C665 VTAIL.n518 B 0.011087f
C666 VTAIL.n519 B 0.019654f
C667 VTAIL.n520 B 0.01548f
C668 VTAIL.t12 B 0.043048f
C669 VTAIL.n521 B 0.122723f
C670 VTAIL.n522 B 1.12583f
C671 VTAIL.n523 B 0.011087f
C672 VTAIL.n524 B 0.011739f
C673 VTAIL.n525 B 0.026206f
C674 VTAIL.n526 B 0.026206f
C675 VTAIL.n527 B 0.011739f
C676 VTAIL.n528 B 0.011087f
C677 VTAIL.n529 B 0.020632f
C678 VTAIL.n530 B 0.020632f
C679 VTAIL.n531 B 0.011087f
C680 VTAIL.n532 B 0.011739f
C681 VTAIL.n533 B 0.026206f
C682 VTAIL.n534 B 0.026206f
C683 VTAIL.n535 B 0.011739f
C684 VTAIL.n536 B 0.011087f
C685 VTAIL.n537 B 0.020632f
C686 VTAIL.n538 B 0.020632f
C687 VTAIL.n539 B 0.011087f
C688 VTAIL.n540 B 0.011739f
C689 VTAIL.n541 B 0.026206f
C690 VTAIL.n542 B 0.026206f
C691 VTAIL.n543 B 0.011739f
C692 VTAIL.n544 B 0.011087f
C693 VTAIL.n545 B 0.020632f
C694 VTAIL.n546 B 0.020632f
C695 VTAIL.n547 B 0.011087f
C696 VTAIL.n548 B 0.011739f
C697 VTAIL.n549 B 0.026206f
C698 VTAIL.n550 B 0.026206f
C699 VTAIL.n551 B 0.011739f
C700 VTAIL.n552 B 0.011087f
C701 VTAIL.n553 B 0.020632f
C702 VTAIL.n554 B 0.020632f
C703 VTAIL.n555 B 0.011087f
C704 VTAIL.n556 B 0.011739f
C705 VTAIL.n557 B 0.026206f
C706 VTAIL.n558 B 0.026206f
C707 VTAIL.n559 B 0.011739f
C708 VTAIL.n560 B 0.011087f
C709 VTAIL.n561 B 0.020632f
C710 VTAIL.n562 B 0.054173f
C711 VTAIL.n563 B 0.011087f
C712 VTAIL.n564 B 0.011739f
C713 VTAIL.n565 B 0.054515f
C714 VTAIL.n566 B 0.046233f
C715 VTAIL.n567 B 1.5164f
C716 VDD2.t1 B 0.273392f
C717 VDD2.t6 B 0.273392f
C718 VDD2.n0 B 2.47447f
C719 VDD2.t4 B 0.273392f
C720 VDD2.t2 B 0.273392f
C721 VDD2.n1 B 2.47447f
C722 VDD2.n2 B 4.45103f
C723 VDD2.t3 B 0.273392f
C724 VDD2.t7 B 0.273392f
C725 VDD2.n3 B 2.45571f
C726 VDD2.n4 B 3.77166f
C727 VDD2.t5 B 0.273392f
C728 VDD2.t0 B 0.273392f
C729 VDD2.n5 B 2.47442f
C730 VN.n0 B 0.031306f
C731 VN.t3 B 2.28022f
C732 VN.n1 B 0.031019f
C733 VN.n2 B 0.016643f
C734 VN.n3 B 0.031019f
C735 VN.n4 B 0.016643f
C736 VN.t1 B 2.28022f
C737 VN.n5 B 0.031019f
C738 VN.n6 B 0.016643f
C739 VN.n7 B 0.031019f
C740 VN.n8 B 0.221324f
C741 VN.t7 B 2.28022f
C742 VN.t4 B 2.55252f
C743 VN.n9 B 0.812266f
C744 VN.n10 B 0.853211f
C745 VN.n11 B 0.019993f
C746 VN.n12 B 0.031019f
C747 VN.n13 B 0.016643f
C748 VN.n14 B 0.016643f
C749 VN.n15 B 0.016643f
C750 VN.n16 B 0.033078f
C751 VN.n17 B 0.013454f
C752 VN.n18 B 0.033078f
C753 VN.n19 B 0.016643f
C754 VN.n20 B 0.016643f
C755 VN.n21 B 0.016643f
C756 VN.n22 B 0.031019f
C757 VN.n23 B 0.019993f
C758 VN.n24 B 0.795857f
C759 VN.n25 B 0.026731f
C760 VN.n26 B 0.016643f
C761 VN.n27 B 0.016643f
C762 VN.n28 B 0.016643f
C763 VN.n29 B 0.031019f
C764 VN.n30 B 0.025687f
C765 VN.n31 B 0.022905f
C766 VN.n32 B 0.016643f
C767 VN.n33 B 0.016643f
C768 VN.n34 B 0.016643f
C769 VN.n35 B 0.031019f
C770 VN.n36 B 0.028568f
C771 VN.n37 B 0.86891f
C772 VN.n38 B 0.05259f
C773 VN.n39 B 0.031306f
C774 VN.t2 B 2.28022f
C775 VN.n40 B 0.031019f
C776 VN.n41 B 0.016643f
C777 VN.n42 B 0.031019f
C778 VN.n43 B 0.016643f
C779 VN.t6 B 2.28022f
C780 VN.n44 B 0.031019f
C781 VN.n45 B 0.016643f
C782 VN.n46 B 0.031019f
C783 VN.n47 B 0.221324f
C784 VN.t0 B 2.28022f
C785 VN.t5 B 2.55252f
C786 VN.n48 B 0.812266f
C787 VN.n49 B 0.853211f
C788 VN.n50 B 0.019993f
C789 VN.n51 B 0.031019f
C790 VN.n52 B 0.016643f
C791 VN.n53 B 0.016643f
C792 VN.n54 B 0.016643f
C793 VN.n55 B 0.033078f
C794 VN.n56 B 0.013454f
C795 VN.n57 B 0.033078f
C796 VN.n58 B 0.016643f
C797 VN.n59 B 0.016643f
C798 VN.n60 B 0.016643f
C799 VN.n61 B 0.031019f
C800 VN.n62 B 0.019993f
C801 VN.n63 B 0.795857f
C802 VN.n64 B 0.026731f
C803 VN.n65 B 0.016643f
C804 VN.n66 B 0.016643f
C805 VN.n67 B 0.016643f
C806 VN.n68 B 0.031019f
C807 VN.n69 B 0.025687f
C808 VN.n70 B 0.022905f
C809 VN.n71 B 0.016643f
C810 VN.n72 B 0.016643f
C811 VN.n73 B 0.016643f
C812 VN.n74 B 0.031019f
C813 VN.n75 B 0.028568f
C814 VN.n76 B 0.86891f
C815 VN.n77 B 1.18971f
.ends

