* NGSPICE file created from diff_pair_sample_1506.ext - technology: sky130A

.subckt diff_pair_sample_1506 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2478_n3236# sky130_fd_pr__pfet_01v8 ad=4.4226 pd=23.46 as=0 ps=0 w=11.34 l=3.44
X1 VDD1.t1 VP.t0 VTAIL.t2 w_n2478_n3236# sky130_fd_pr__pfet_01v8 ad=4.4226 pd=23.46 as=4.4226 ps=23.46 w=11.34 l=3.44
X2 VDD1.t0 VP.t1 VTAIL.t1 w_n2478_n3236# sky130_fd_pr__pfet_01v8 ad=4.4226 pd=23.46 as=4.4226 ps=23.46 w=11.34 l=3.44
X3 B.t8 B.t6 B.t7 w_n2478_n3236# sky130_fd_pr__pfet_01v8 ad=4.4226 pd=23.46 as=0 ps=0 w=11.34 l=3.44
X4 VDD2.t1 VN.t0 VTAIL.t3 w_n2478_n3236# sky130_fd_pr__pfet_01v8 ad=4.4226 pd=23.46 as=4.4226 ps=23.46 w=11.34 l=3.44
X5 B.t5 B.t3 B.t4 w_n2478_n3236# sky130_fd_pr__pfet_01v8 ad=4.4226 pd=23.46 as=0 ps=0 w=11.34 l=3.44
X6 B.t2 B.t0 B.t1 w_n2478_n3236# sky130_fd_pr__pfet_01v8 ad=4.4226 pd=23.46 as=0 ps=0 w=11.34 l=3.44
X7 VDD2.t0 VN.t1 VTAIL.t0 w_n2478_n3236# sky130_fd_pr__pfet_01v8 ad=4.4226 pd=23.46 as=4.4226 ps=23.46 w=11.34 l=3.44
R0 B.n338 B.n337 585
R1 B.n336 B.n97 585
R2 B.n335 B.n334 585
R3 B.n333 B.n98 585
R4 B.n332 B.n331 585
R5 B.n330 B.n99 585
R6 B.n329 B.n328 585
R7 B.n327 B.n100 585
R8 B.n326 B.n325 585
R9 B.n324 B.n101 585
R10 B.n323 B.n322 585
R11 B.n321 B.n102 585
R12 B.n320 B.n319 585
R13 B.n318 B.n103 585
R14 B.n317 B.n316 585
R15 B.n315 B.n104 585
R16 B.n314 B.n313 585
R17 B.n312 B.n105 585
R18 B.n311 B.n310 585
R19 B.n309 B.n106 585
R20 B.n308 B.n307 585
R21 B.n306 B.n107 585
R22 B.n305 B.n304 585
R23 B.n303 B.n108 585
R24 B.n302 B.n301 585
R25 B.n300 B.n109 585
R26 B.n299 B.n298 585
R27 B.n297 B.n110 585
R28 B.n296 B.n295 585
R29 B.n294 B.n111 585
R30 B.n293 B.n292 585
R31 B.n291 B.n112 585
R32 B.n290 B.n289 585
R33 B.n288 B.n113 585
R34 B.n287 B.n286 585
R35 B.n285 B.n114 585
R36 B.n284 B.n283 585
R37 B.n282 B.n115 585
R38 B.n281 B.n280 585
R39 B.n279 B.n116 585
R40 B.n278 B.n277 585
R41 B.n273 B.n117 585
R42 B.n272 B.n271 585
R43 B.n270 B.n118 585
R44 B.n269 B.n268 585
R45 B.n267 B.n119 585
R46 B.n266 B.n265 585
R47 B.n264 B.n120 585
R48 B.n263 B.n262 585
R49 B.n260 B.n121 585
R50 B.n259 B.n258 585
R51 B.n257 B.n124 585
R52 B.n256 B.n255 585
R53 B.n254 B.n125 585
R54 B.n253 B.n252 585
R55 B.n251 B.n126 585
R56 B.n250 B.n249 585
R57 B.n248 B.n127 585
R58 B.n247 B.n246 585
R59 B.n245 B.n128 585
R60 B.n244 B.n243 585
R61 B.n242 B.n129 585
R62 B.n241 B.n240 585
R63 B.n239 B.n130 585
R64 B.n238 B.n237 585
R65 B.n236 B.n131 585
R66 B.n235 B.n234 585
R67 B.n233 B.n132 585
R68 B.n232 B.n231 585
R69 B.n230 B.n133 585
R70 B.n229 B.n228 585
R71 B.n227 B.n134 585
R72 B.n226 B.n225 585
R73 B.n224 B.n135 585
R74 B.n223 B.n222 585
R75 B.n221 B.n136 585
R76 B.n220 B.n219 585
R77 B.n218 B.n137 585
R78 B.n217 B.n216 585
R79 B.n215 B.n138 585
R80 B.n214 B.n213 585
R81 B.n212 B.n139 585
R82 B.n211 B.n210 585
R83 B.n209 B.n140 585
R84 B.n208 B.n207 585
R85 B.n206 B.n141 585
R86 B.n205 B.n204 585
R87 B.n203 B.n142 585
R88 B.n202 B.n201 585
R89 B.n339 B.n96 585
R90 B.n341 B.n340 585
R91 B.n342 B.n95 585
R92 B.n344 B.n343 585
R93 B.n345 B.n94 585
R94 B.n347 B.n346 585
R95 B.n348 B.n93 585
R96 B.n350 B.n349 585
R97 B.n351 B.n92 585
R98 B.n353 B.n352 585
R99 B.n354 B.n91 585
R100 B.n356 B.n355 585
R101 B.n357 B.n90 585
R102 B.n359 B.n358 585
R103 B.n360 B.n89 585
R104 B.n362 B.n361 585
R105 B.n363 B.n88 585
R106 B.n365 B.n364 585
R107 B.n366 B.n87 585
R108 B.n368 B.n367 585
R109 B.n369 B.n86 585
R110 B.n371 B.n370 585
R111 B.n372 B.n85 585
R112 B.n374 B.n373 585
R113 B.n375 B.n84 585
R114 B.n377 B.n376 585
R115 B.n378 B.n83 585
R116 B.n380 B.n379 585
R117 B.n381 B.n82 585
R118 B.n383 B.n382 585
R119 B.n384 B.n81 585
R120 B.n386 B.n385 585
R121 B.n387 B.n80 585
R122 B.n389 B.n388 585
R123 B.n390 B.n79 585
R124 B.n392 B.n391 585
R125 B.n393 B.n78 585
R126 B.n395 B.n394 585
R127 B.n396 B.n77 585
R128 B.n398 B.n397 585
R129 B.n399 B.n76 585
R130 B.n401 B.n400 585
R131 B.n402 B.n75 585
R132 B.n404 B.n403 585
R133 B.n405 B.n74 585
R134 B.n407 B.n406 585
R135 B.n408 B.n73 585
R136 B.n410 B.n409 585
R137 B.n411 B.n72 585
R138 B.n413 B.n412 585
R139 B.n414 B.n71 585
R140 B.n416 B.n415 585
R141 B.n417 B.n70 585
R142 B.n419 B.n418 585
R143 B.n420 B.n69 585
R144 B.n422 B.n421 585
R145 B.n423 B.n68 585
R146 B.n425 B.n424 585
R147 B.n426 B.n67 585
R148 B.n428 B.n427 585
R149 B.n429 B.n66 585
R150 B.n431 B.n430 585
R151 B.n566 B.n17 585
R152 B.n565 B.n564 585
R153 B.n563 B.n18 585
R154 B.n562 B.n561 585
R155 B.n560 B.n19 585
R156 B.n559 B.n558 585
R157 B.n557 B.n20 585
R158 B.n556 B.n555 585
R159 B.n554 B.n21 585
R160 B.n553 B.n552 585
R161 B.n551 B.n22 585
R162 B.n550 B.n549 585
R163 B.n548 B.n23 585
R164 B.n547 B.n546 585
R165 B.n545 B.n24 585
R166 B.n544 B.n543 585
R167 B.n542 B.n25 585
R168 B.n541 B.n540 585
R169 B.n539 B.n26 585
R170 B.n538 B.n537 585
R171 B.n536 B.n27 585
R172 B.n535 B.n534 585
R173 B.n533 B.n28 585
R174 B.n532 B.n531 585
R175 B.n530 B.n29 585
R176 B.n529 B.n528 585
R177 B.n527 B.n30 585
R178 B.n526 B.n525 585
R179 B.n524 B.n31 585
R180 B.n523 B.n522 585
R181 B.n521 B.n32 585
R182 B.n520 B.n519 585
R183 B.n518 B.n33 585
R184 B.n517 B.n516 585
R185 B.n515 B.n34 585
R186 B.n514 B.n513 585
R187 B.n512 B.n35 585
R188 B.n511 B.n510 585
R189 B.n509 B.n36 585
R190 B.n508 B.n507 585
R191 B.n505 B.n37 585
R192 B.n504 B.n503 585
R193 B.n502 B.n40 585
R194 B.n501 B.n500 585
R195 B.n499 B.n41 585
R196 B.n498 B.n497 585
R197 B.n496 B.n42 585
R198 B.n495 B.n494 585
R199 B.n493 B.n43 585
R200 B.n491 B.n490 585
R201 B.n489 B.n46 585
R202 B.n488 B.n487 585
R203 B.n486 B.n47 585
R204 B.n485 B.n484 585
R205 B.n483 B.n48 585
R206 B.n482 B.n481 585
R207 B.n480 B.n49 585
R208 B.n479 B.n478 585
R209 B.n477 B.n50 585
R210 B.n476 B.n475 585
R211 B.n474 B.n51 585
R212 B.n473 B.n472 585
R213 B.n471 B.n52 585
R214 B.n470 B.n469 585
R215 B.n468 B.n53 585
R216 B.n467 B.n466 585
R217 B.n465 B.n54 585
R218 B.n464 B.n463 585
R219 B.n462 B.n55 585
R220 B.n461 B.n460 585
R221 B.n459 B.n56 585
R222 B.n458 B.n457 585
R223 B.n456 B.n57 585
R224 B.n455 B.n454 585
R225 B.n453 B.n58 585
R226 B.n452 B.n451 585
R227 B.n450 B.n59 585
R228 B.n449 B.n448 585
R229 B.n447 B.n60 585
R230 B.n446 B.n445 585
R231 B.n444 B.n61 585
R232 B.n443 B.n442 585
R233 B.n441 B.n62 585
R234 B.n440 B.n439 585
R235 B.n438 B.n63 585
R236 B.n437 B.n436 585
R237 B.n435 B.n64 585
R238 B.n434 B.n433 585
R239 B.n432 B.n65 585
R240 B.n568 B.n567 585
R241 B.n569 B.n16 585
R242 B.n571 B.n570 585
R243 B.n572 B.n15 585
R244 B.n574 B.n573 585
R245 B.n575 B.n14 585
R246 B.n577 B.n576 585
R247 B.n578 B.n13 585
R248 B.n580 B.n579 585
R249 B.n581 B.n12 585
R250 B.n583 B.n582 585
R251 B.n584 B.n11 585
R252 B.n586 B.n585 585
R253 B.n587 B.n10 585
R254 B.n589 B.n588 585
R255 B.n590 B.n9 585
R256 B.n592 B.n591 585
R257 B.n593 B.n8 585
R258 B.n595 B.n594 585
R259 B.n596 B.n7 585
R260 B.n598 B.n597 585
R261 B.n599 B.n6 585
R262 B.n601 B.n600 585
R263 B.n602 B.n5 585
R264 B.n604 B.n603 585
R265 B.n605 B.n4 585
R266 B.n607 B.n606 585
R267 B.n608 B.n3 585
R268 B.n610 B.n609 585
R269 B.n611 B.n0 585
R270 B.n2 B.n1 585
R271 B.n158 B.n157 585
R272 B.n160 B.n159 585
R273 B.n161 B.n156 585
R274 B.n163 B.n162 585
R275 B.n164 B.n155 585
R276 B.n166 B.n165 585
R277 B.n167 B.n154 585
R278 B.n169 B.n168 585
R279 B.n170 B.n153 585
R280 B.n172 B.n171 585
R281 B.n173 B.n152 585
R282 B.n175 B.n174 585
R283 B.n176 B.n151 585
R284 B.n178 B.n177 585
R285 B.n179 B.n150 585
R286 B.n181 B.n180 585
R287 B.n182 B.n149 585
R288 B.n184 B.n183 585
R289 B.n185 B.n148 585
R290 B.n187 B.n186 585
R291 B.n188 B.n147 585
R292 B.n190 B.n189 585
R293 B.n191 B.n146 585
R294 B.n193 B.n192 585
R295 B.n194 B.n145 585
R296 B.n196 B.n195 585
R297 B.n197 B.n144 585
R298 B.n199 B.n198 585
R299 B.n200 B.n143 585
R300 B.n202 B.n143 458.866
R301 B.n339 B.n338 458.866
R302 B.n430 B.n65 458.866
R303 B.n568 B.n17 458.866
R304 B.n274 B.t1 436.788
R305 B.n44 B.t8 436.788
R306 B.n122 B.t10 436.788
R307 B.n38 B.t5 436.788
R308 B.n275 B.t2 363.673
R309 B.n45 B.t7 363.673
R310 B.n123 B.t11 363.673
R311 B.n39 B.t4 363.673
R312 B.n122 B.t9 288.486
R313 B.n274 B.t0 288.486
R314 B.n44 B.t6 288.486
R315 B.n38 B.t3 288.486
R316 B.n613 B.n612 256.663
R317 B.n612 B.n611 235.042
R318 B.n612 B.n2 235.042
R319 B.n203 B.n202 163.367
R320 B.n204 B.n203 163.367
R321 B.n204 B.n141 163.367
R322 B.n208 B.n141 163.367
R323 B.n209 B.n208 163.367
R324 B.n210 B.n209 163.367
R325 B.n210 B.n139 163.367
R326 B.n214 B.n139 163.367
R327 B.n215 B.n214 163.367
R328 B.n216 B.n215 163.367
R329 B.n216 B.n137 163.367
R330 B.n220 B.n137 163.367
R331 B.n221 B.n220 163.367
R332 B.n222 B.n221 163.367
R333 B.n222 B.n135 163.367
R334 B.n226 B.n135 163.367
R335 B.n227 B.n226 163.367
R336 B.n228 B.n227 163.367
R337 B.n228 B.n133 163.367
R338 B.n232 B.n133 163.367
R339 B.n233 B.n232 163.367
R340 B.n234 B.n233 163.367
R341 B.n234 B.n131 163.367
R342 B.n238 B.n131 163.367
R343 B.n239 B.n238 163.367
R344 B.n240 B.n239 163.367
R345 B.n240 B.n129 163.367
R346 B.n244 B.n129 163.367
R347 B.n245 B.n244 163.367
R348 B.n246 B.n245 163.367
R349 B.n246 B.n127 163.367
R350 B.n250 B.n127 163.367
R351 B.n251 B.n250 163.367
R352 B.n252 B.n251 163.367
R353 B.n252 B.n125 163.367
R354 B.n256 B.n125 163.367
R355 B.n257 B.n256 163.367
R356 B.n258 B.n257 163.367
R357 B.n258 B.n121 163.367
R358 B.n263 B.n121 163.367
R359 B.n264 B.n263 163.367
R360 B.n265 B.n264 163.367
R361 B.n265 B.n119 163.367
R362 B.n269 B.n119 163.367
R363 B.n270 B.n269 163.367
R364 B.n271 B.n270 163.367
R365 B.n271 B.n117 163.367
R366 B.n278 B.n117 163.367
R367 B.n279 B.n278 163.367
R368 B.n280 B.n279 163.367
R369 B.n280 B.n115 163.367
R370 B.n284 B.n115 163.367
R371 B.n285 B.n284 163.367
R372 B.n286 B.n285 163.367
R373 B.n286 B.n113 163.367
R374 B.n290 B.n113 163.367
R375 B.n291 B.n290 163.367
R376 B.n292 B.n291 163.367
R377 B.n292 B.n111 163.367
R378 B.n296 B.n111 163.367
R379 B.n297 B.n296 163.367
R380 B.n298 B.n297 163.367
R381 B.n298 B.n109 163.367
R382 B.n302 B.n109 163.367
R383 B.n303 B.n302 163.367
R384 B.n304 B.n303 163.367
R385 B.n304 B.n107 163.367
R386 B.n308 B.n107 163.367
R387 B.n309 B.n308 163.367
R388 B.n310 B.n309 163.367
R389 B.n310 B.n105 163.367
R390 B.n314 B.n105 163.367
R391 B.n315 B.n314 163.367
R392 B.n316 B.n315 163.367
R393 B.n316 B.n103 163.367
R394 B.n320 B.n103 163.367
R395 B.n321 B.n320 163.367
R396 B.n322 B.n321 163.367
R397 B.n322 B.n101 163.367
R398 B.n326 B.n101 163.367
R399 B.n327 B.n326 163.367
R400 B.n328 B.n327 163.367
R401 B.n328 B.n99 163.367
R402 B.n332 B.n99 163.367
R403 B.n333 B.n332 163.367
R404 B.n334 B.n333 163.367
R405 B.n334 B.n97 163.367
R406 B.n338 B.n97 163.367
R407 B.n430 B.n429 163.367
R408 B.n429 B.n428 163.367
R409 B.n428 B.n67 163.367
R410 B.n424 B.n67 163.367
R411 B.n424 B.n423 163.367
R412 B.n423 B.n422 163.367
R413 B.n422 B.n69 163.367
R414 B.n418 B.n69 163.367
R415 B.n418 B.n417 163.367
R416 B.n417 B.n416 163.367
R417 B.n416 B.n71 163.367
R418 B.n412 B.n71 163.367
R419 B.n412 B.n411 163.367
R420 B.n411 B.n410 163.367
R421 B.n410 B.n73 163.367
R422 B.n406 B.n73 163.367
R423 B.n406 B.n405 163.367
R424 B.n405 B.n404 163.367
R425 B.n404 B.n75 163.367
R426 B.n400 B.n75 163.367
R427 B.n400 B.n399 163.367
R428 B.n399 B.n398 163.367
R429 B.n398 B.n77 163.367
R430 B.n394 B.n77 163.367
R431 B.n394 B.n393 163.367
R432 B.n393 B.n392 163.367
R433 B.n392 B.n79 163.367
R434 B.n388 B.n79 163.367
R435 B.n388 B.n387 163.367
R436 B.n387 B.n386 163.367
R437 B.n386 B.n81 163.367
R438 B.n382 B.n81 163.367
R439 B.n382 B.n381 163.367
R440 B.n381 B.n380 163.367
R441 B.n380 B.n83 163.367
R442 B.n376 B.n83 163.367
R443 B.n376 B.n375 163.367
R444 B.n375 B.n374 163.367
R445 B.n374 B.n85 163.367
R446 B.n370 B.n85 163.367
R447 B.n370 B.n369 163.367
R448 B.n369 B.n368 163.367
R449 B.n368 B.n87 163.367
R450 B.n364 B.n87 163.367
R451 B.n364 B.n363 163.367
R452 B.n363 B.n362 163.367
R453 B.n362 B.n89 163.367
R454 B.n358 B.n89 163.367
R455 B.n358 B.n357 163.367
R456 B.n357 B.n356 163.367
R457 B.n356 B.n91 163.367
R458 B.n352 B.n91 163.367
R459 B.n352 B.n351 163.367
R460 B.n351 B.n350 163.367
R461 B.n350 B.n93 163.367
R462 B.n346 B.n93 163.367
R463 B.n346 B.n345 163.367
R464 B.n345 B.n344 163.367
R465 B.n344 B.n95 163.367
R466 B.n340 B.n95 163.367
R467 B.n340 B.n339 163.367
R468 B.n564 B.n17 163.367
R469 B.n564 B.n563 163.367
R470 B.n563 B.n562 163.367
R471 B.n562 B.n19 163.367
R472 B.n558 B.n19 163.367
R473 B.n558 B.n557 163.367
R474 B.n557 B.n556 163.367
R475 B.n556 B.n21 163.367
R476 B.n552 B.n21 163.367
R477 B.n552 B.n551 163.367
R478 B.n551 B.n550 163.367
R479 B.n550 B.n23 163.367
R480 B.n546 B.n23 163.367
R481 B.n546 B.n545 163.367
R482 B.n545 B.n544 163.367
R483 B.n544 B.n25 163.367
R484 B.n540 B.n25 163.367
R485 B.n540 B.n539 163.367
R486 B.n539 B.n538 163.367
R487 B.n538 B.n27 163.367
R488 B.n534 B.n27 163.367
R489 B.n534 B.n533 163.367
R490 B.n533 B.n532 163.367
R491 B.n532 B.n29 163.367
R492 B.n528 B.n29 163.367
R493 B.n528 B.n527 163.367
R494 B.n527 B.n526 163.367
R495 B.n526 B.n31 163.367
R496 B.n522 B.n31 163.367
R497 B.n522 B.n521 163.367
R498 B.n521 B.n520 163.367
R499 B.n520 B.n33 163.367
R500 B.n516 B.n33 163.367
R501 B.n516 B.n515 163.367
R502 B.n515 B.n514 163.367
R503 B.n514 B.n35 163.367
R504 B.n510 B.n35 163.367
R505 B.n510 B.n509 163.367
R506 B.n509 B.n508 163.367
R507 B.n508 B.n37 163.367
R508 B.n503 B.n37 163.367
R509 B.n503 B.n502 163.367
R510 B.n502 B.n501 163.367
R511 B.n501 B.n41 163.367
R512 B.n497 B.n41 163.367
R513 B.n497 B.n496 163.367
R514 B.n496 B.n495 163.367
R515 B.n495 B.n43 163.367
R516 B.n490 B.n43 163.367
R517 B.n490 B.n489 163.367
R518 B.n489 B.n488 163.367
R519 B.n488 B.n47 163.367
R520 B.n484 B.n47 163.367
R521 B.n484 B.n483 163.367
R522 B.n483 B.n482 163.367
R523 B.n482 B.n49 163.367
R524 B.n478 B.n49 163.367
R525 B.n478 B.n477 163.367
R526 B.n477 B.n476 163.367
R527 B.n476 B.n51 163.367
R528 B.n472 B.n51 163.367
R529 B.n472 B.n471 163.367
R530 B.n471 B.n470 163.367
R531 B.n470 B.n53 163.367
R532 B.n466 B.n53 163.367
R533 B.n466 B.n465 163.367
R534 B.n465 B.n464 163.367
R535 B.n464 B.n55 163.367
R536 B.n460 B.n55 163.367
R537 B.n460 B.n459 163.367
R538 B.n459 B.n458 163.367
R539 B.n458 B.n57 163.367
R540 B.n454 B.n57 163.367
R541 B.n454 B.n453 163.367
R542 B.n453 B.n452 163.367
R543 B.n452 B.n59 163.367
R544 B.n448 B.n59 163.367
R545 B.n448 B.n447 163.367
R546 B.n447 B.n446 163.367
R547 B.n446 B.n61 163.367
R548 B.n442 B.n61 163.367
R549 B.n442 B.n441 163.367
R550 B.n441 B.n440 163.367
R551 B.n440 B.n63 163.367
R552 B.n436 B.n63 163.367
R553 B.n436 B.n435 163.367
R554 B.n435 B.n434 163.367
R555 B.n434 B.n65 163.367
R556 B.n569 B.n568 163.367
R557 B.n570 B.n569 163.367
R558 B.n570 B.n15 163.367
R559 B.n574 B.n15 163.367
R560 B.n575 B.n574 163.367
R561 B.n576 B.n575 163.367
R562 B.n576 B.n13 163.367
R563 B.n580 B.n13 163.367
R564 B.n581 B.n580 163.367
R565 B.n582 B.n581 163.367
R566 B.n582 B.n11 163.367
R567 B.n586 B.n11 163.367
R568 B.n587 B.n586 163.367
R569 B.n588 B.n587 163.367
R570 B.n588 B.n9 163.367
R571 B.n592 B.n9 163.367
R572 B.n593 B.n592 163.367
R573 B.n594 B.n593 163.367
R574 B.n594 B.n7 163.367
R575 B.n598 B.n7 163.367
R576 B.n599 B.n598 163.367
R577 B.n600 B.n599 163.367
R578 B.n600 B.n5 163.367
R579 B.n604 B.n5 163.367
R580 B.n605 B.n604 163.367
R581 B.n606 B.n605 163.367
R582 B.n606 B.n3 163.367
R583 B.n610 B.n3 163.367
R584 B.n611 B.n610 163.367
R585 B.n157 B.n2 163.367
R586 B.n160 B.n157 163.367
R587 B.n161 B.n160 163.367
R588 B.n162 B.n161 163.367
R589 B.n162 B.n155 163.367
R590 B.n166 B.n155 163.367
R591 B.n167 B.n166 163.367
R592 B.n168 B.n167 163.367
R593 B.n168 B.n153 163.367
R594 B.n172 B.n153 163.367
R595 B.n173 B.n172 163.367
R596 B.n174 B.n173 163.367
R597 B.n174 B.n151 163.367
R598 B.n178 B.n151 163.367
R599 B.n179 B.n178 163.367
R600 B.n180 B.n179 163.367
R601 B.n180 B.n149 163.367
R602 B.n184 B.n149 163.367
R603 B.n185 B.n184 163.367
R604 B.n186 B.n185 163.367
R605 B.n186 B.n147 163.367
R606 B.n190 B.n147 163.367
R607 B.n191 B.n190 163.367
R608 B.n192 B.n191 163.367
R609 B.n192 B.n145 163.367
R610 B.n196 B.n145 163.367
R611 B.n197 B.n196 163.367
R612 B.n198 B.n197 163.367
R613 B.n198 B.n143 163.367
R614 B.n123 B.n122 73.1157
R615 B.n275 B.n274 73.1157
R616 B.n45 B.n44 73.1157
R617 B.n39 B.n38 73.1157
R618 B.n261 B.n123 59.5399
R619 B.n276 B.n275 59.5399
R620 B.n492 B.n45 59.5399
R621 B.n506 B.n39 59.5399
R622 B.n567 B.n566 29.8151
R623 B.n432 B.n431 29.8151
R624 B.n201 B.n200 29.8151
R625 B.n337 B.n96 29.8151
R626 B B.n613 18.0485
R627 B.n567 B.n16 10.6151
R628 B.n571 B.n16 10.6151
R629 B.n572 B.n571 10.6151
R630 B.n573 B.n572 10.6151
R631 B.n573 B.n14 10.6151
R632 B.n577 B.n14 10.6151
R633 B.n578 B.n577 10.6151
R634 B.n579 B.n578 10.6151
R635 B.n579 B.n12 10.6151
R636 B.n583 B.n12 10.6151
R637 B.n584 B.n583 10.6151
R638 B.n585 B.n584 10.6151
R639 B.n585 B.n10 10.6151
R640 B.n589 B.n10 10.6151
R641 B.n590 B.n589 10.6151
R642 B.n591 B.n590 10.6151
R643 B.n591 B.n8 10.6151
R644 B.n595 B.n8 10.6151
R645 B.n596 B.n595 10.6151
R646 B.n597 B.n596 10.6151
R647 B.n597 B.n6 10.6151
R648 B.n601 B.n6 10.6151
R649 B.n602 B.n601 10.6151
R650 B.n603 B.n602 10.6151
R651 B.n603 B.n4 10.6151
R652 B.n607 B.n4 10.6151
R653 B.n608 B.n607 10.6151
R654 B.n609 B.n608 10.6151
R655 B.n609 B.n0 10.6151
R656 B.n566 B.n565 10.6151
R657 B.n565 B.n18 10.6151
R658 B.n561 B.n18 10.6151
R659 B.n561 B.n560 10.6151
R660 B.n560 B.n559 10.6151
R661 B.n559 B.n20 10.6151
R662 B.n555 B.n20 10.6151
R663 B.n555 B.n554 10.6151
R664 B.n554 B.n553 10.6151
R665 B.n553 B.n22 10.6151
R666 B.n549 B.n22 10.6151
R667 B.n549 B.n548 10.6151
R668 B.n548 B.n547 10.6151
R669 B.n547 B.n24 10.6151
R670 B.n543 B.n24 10.6151
R671 B.n543 B.n542 10.6151
R672 B.n542 B.n541 10.6151
R673 B.n541 B.n26 10.6151
R674 B.n537 B.n26 10.6151
R675 B.n537 B.n536 10.6151
R676 B.n536 B.n535 10.6151
R677 B.n535 B.n28 10.6151
R678 B.n531 B.n28 10.6151
R679 B.n531 B.n530 10.6151
R680 B.n530 B.n529 10.6151
R681 B.n529 B.n30 10.6151
R682 B.n525 B.n30 10.6151
R683 B.n525 B.n524 10.6151
R684 B.n524 B.n523 10.6151
R685 B.n523 B.n32 10.6151
R686 B.n519 B.n32 10.6151
R687 B.n519 B.n518 10.6151
R688 B.n518 B.n517 10.6151
R689 B.n517 B.n34 10.6151
R690 B.n513 B.n34 10.6151
R691 B.n513 B.n512 10.6151
R692 B.n512 B.n511 10.6151
R693 B.n511 B.n36 10.6151
R694 B.n507 B.n36 10.6151
R695 B.n505 B.n504 10.6151
R696 B.n504 B.n40 10.6151
R697 B.n500 B.n40 10.6151
R698 B.n500 B.n499 10.6151
R699 B.n499 B.n498 10.6151
R700 B.n498 B.n42 10.6151
R701 B.n494 B.n42 10.6151
R702 B.n494 B.n493 10.6151
R703 B.n491 B.n46 10.6151
R704 B.n487 B.n46 10.6151
R705 B.n487 B.n486 10.6151
R706 B.n486 B.n485 10.6151
R707 B.n485 B.n48 10.6151
R708 B.n481 B.n48 10.6151
R709 B.n481 B.n480 10.6151
R710 B.n480 B.n479 10.6151
R711 B.n479 B.n50 10.6151
R712 B.n475 B.n50 10.6151
R713 B.n475 B.n474 10.6151
R714 B.n474 B.n473 10.6151
R715 B.n473 B.n52 10.6151
R716 B.n469 B.n52 10.6151
R717 B.n469 B.n468 10.6151
R718 B.n468 B.n467 10.6151
R719 B.n467 B.n54 10.6151
R720 B.n463 B.n54 10.6151
R721 B.n463 B.n462 10.6151
R722 B.n462 B.n461 10.6151
R723 B.n461 B.n56 10.6151
R724 B.n457 B.n56 10.6151
R725 B.n457 B.n456 10.6151
R726 B.n456 B.n455 10.6151
R727 B.n455 B.n58 10.6151
R728 B.n451 B.n58 10.6151
R729 B.n451 B.n450 10.6151
R730 B.n450 B.n449 10.6151
R731 B.n449 B.n60 10.6151
R732 B.n445 B.n60 10.6151
R733 B.n445 B.n444 10.6151
R734 B.n444 B.n443 10.6151
R735 B.n443 B.n62 10.6151
R736 B.n439 B.n62 10.6151
R737 B.n439 B.n438 10.6151
R738 B.n438 B.n437 10.6151
R739 B.n437 B.n64 10.6151
R740 B.n433 B.n64 10.6151
R741 B.n433 B.n432 10.6151
R742 B.n431 B.n66 10.6151
R743 B.n427 B.n66 10.6151
R744 B.n427 B.n426 10.6151
R745 B.n426 B.n425 10.6151
R746 B.n425 B.n68 10.6151
R747 B.n421 B.n68 10.6151
R748 B.n421 B.n420 10.6151
R749 B.n420 B.n419 10.6151
R750 B.n419 B.n70 10.6151
R751 B.n415 B.n70 10.6151
R752 B.n415 B.n414 10.6151
R753 B.n414 B.n413 10.6151
R754 B.n413 B.n72 10.6151
R755 B.n409 B.n72 10.6151
R756 B.n409 B.n408 10.6151
R757 B.n408 B.n407 10.6151
R758 B.n407 B.n74 10.6151
R759 B.n403 B.n74 10.6151
R760 B.n403 B.n402 10.6151
R761 B.n402 B.n401 10.6151
R762 B.n401 B.n76 10.6151
R763 B.n397 B.n76 10.6151
R764 B.n397 B.n396 10.6151
R765 B.n396 B.n395 10.6151
R766 B.n395 B.n78 10.6151
R767 B.n391 B.n78 10.6151
R768 B.n391 B.n390 10.6151
R769 B.n390 B.n389 10.6151
R770 B.n389 B.n80 10.6151
R771 B.n385 B.n80 10.6151
R772 B.n385 B.n384 10.6151
R773 B.n384 B.n383 10.6151
R774 B.n383 B.n82 10.6151
R775 B.n379 B.n82 10.6151
R776 B.n379 B.n378 10.6151
R777 B.n378 B.n377 10.6151
R778 B.n377 B.n84 10.6151
R779 B.n373 B.n84 10.6151
R780 B.n373 B.n372 10.6151
R781 B.n372 B.n371 10.6151
R782 B.n371 B.n86 10.6151
R783 B.n367 B.n86 10.6151
R784 B.n367 B.n366 10.6151
R785 B.n366 B.n365 10.6151
R786 B.n365 B.n88 10.6151
R787 B.n361 B.n88 10.6151
R788 B.n361 B.n360 10.6151
R789 B.n360 B.n359 10.6151
R790 B.n359 B.n90 10.6151
R791 B.n355 B.n90 10.6151
R792 B.n355 B.n354 10.6151
R793 B.n354 B.n353 10.6151
R794 B.n353 B.n92 10.6151
R795 B.n349 B.n92 10.6151
R796 B.n349 B.n348 10.6151
R797 B.n348 B.n347 10.6151
R798 B.n347 B.n94 10.6151
R799 B.n343 B.n94 10.6151
R800 B.n343 B.n342 10.6151
R801 B.n342 B.n341 10.6151
R802 B.n341 B.n96 10.6151
R803 B.n158 B.n1 10.6151
R804 B.n159 B.n158 10.6151
R805 B.n159 B.n156 10.6151
R806 B.n163 B.n156 10.6151
R807 B.n164 B.n163 10.6151
R808 B.n165 B.n164 10.6151
R809 B.n165 B.n154 10.6151
R810 B.n169 B.n154 10.6151
R811 B.n170 B.n169 10.6151
R812 B.n171 B.n170 10.6151
R813 B.n171 B.n152 10.6151
R814 B.n175 B.n152 10.6151
R815 B.n176 B.n175 10.6151
R816 B.n177 B.n176 10.6151
R817 B.n177 B.n150 10.6151
R818 B.n181 B.n150 10.6151
R819 B.n182 B.n181 10.6151
R820 B.n183 B.n182 10.6151
R821 B.n183 B.n148 10.6151
R822 B.n187 B.n148 10.6151
R823 B.n188 B.n187 10.6151
R824 B.n189 B.n188 10.6151
R825 B.n189 B.n146 10.6151
R826 B.n193 B.n146 10.6151
R827 B.n194 B.n193 10.6151
R828 B.n195 B.n194 10.6151
R829 B.n195 B.n144 10.6151
R830 B.n199 B.n144 10.6151
R831 B.n200 B.n199 10.6151
R832 B.n201 B.n142 10.6151
R833 B.n205 B.n142 10.6151
R834 B.n206 B.n205 10.6151
R835 B.n207 B.n206 10.6151
R836 B.n207 B.n140 10.6151
R837 B.n211 B.n140 10.6151
R838 B.n212 B.n211 10.6151
R839 B.n213 B.n212 10.6151
R840 B.n213 B.n138 10.6151
R841 B.n217 B.n138 10.6151
R842 B.n218 B.n217 10.6151
R843 B.n219 B.n218 10.6151
R844 B.n219 B.n136 10.6151
R845 B.n223 B.n136 10.6151
R846 B.n224 B.n223 10.6151
R847 B.n225 B.n224 10.6151
R848 B.n225 B.n134 10.6151
R849 B.n229 B.n134 10.6151
R850 B.n230 B.n229 10.6151
R851 B.n231 B.n230 10.6151
R852 B.n231 B.n132 10.6151
R853 B.n235 B.n132 10.6151
R854 B.n236 B.n235 10.6151
R855 B.n237 B.n236 10.6151
R856 B.n237 B.n130 10.6151
R857 B.n241 B.n130 10.6151
R858 B.n242 B.n241 10.6151
R859 B.n243 B.n242 10.6151
R860 B.n243 B.n128 10.6151
R861 B.n247 B.n128 10.6151
R862 B.n248 B.n247 10.6151
R863 B.n249 B.n248 10.6151
R864 B.n249 B.n126 10.6151
R865 B.n253 B.n126 10.6151
R866 B.n254 B.n253 10.6151
R867 B.n255 B.n254 10.6151
R868 B.n255 B.n124 10.6151
R869 B.n259 B.n124 10.6151
R870 B.n260 B.n259 10.6151
R871 B.n262 B.n120 10.6151
R872 B.n266 B.n120 10.6151
R873 B.n267 B.n266 10.6151
R874 B.n268 B.n267 10.6151
R875 B.n268 B.n118 10.6151
R876 B.n272 B.n118 10.6151
R877 B.n273 B.n272 10.6151
R878 B.n277 B.n273 10.6151
R879 B.n281 B.n116 10.6151
R880 B.n282 B.n281 10.6151
R881 B.n283 B.n282 10.6151
R882 B.n283 B.n114 10.6151
R883 B.n287 B.n114 10.6151
R884 B.n288 B.n287 10.6151
R885 B.n289 B.n288 10.6151
R886 B.n289 B.n112 10.6151
R887 B.n293 B.n112 10.6151
R888 B.n294 B.n293 10.6151
R889 B.n295 B.n294 10.6151
R890 B.n295 B.n110 10.6151
R891 B.n299 B.n110 10.6151
R892 B.n300 B.n299 10.6151
R893 B.n301 B.n300 10.6151
R894 B.n301 B.n108 10.6151
R895 B.n305 B.n108 10.6151
R896 B.n306 B.n305 10.6151
R897 B.n307 B.n306 10.6151
R898 B.n307 B.n106 10.6151
R899 B.n311 B.n106 10.6151
R900 B.n312 B.n311 10.6151
R901 B.n313 B.n312 10.6151
R902 B.n313 B.n104 10.6151
R903 B.n317 B.n104 10.6151
R904 B.n318 B.n317 10.6151
R905 B.n319 B.n318 10.6151
R906 B.n319 B.n102 10.6151
R907 B.n323 B.n102 10.6151
R908 B.n324 B.n323 10.6151
R909 B.n325 B.n324 10.6151
R910 B.n325 B.n100 10.6151
R911 B.n329 B.n100 10.6151
R912 B.n330 B.n329 10.6151
R913 B.n331 B.n330 10.6151
R914 B.n331 B.n98 10.6151
R915 B.n335 B.n98 10.6151
R916 B.n336 B.n335 10.6151
R917 B.n337 B.n336 10.6151
R918 B.n613 B.n0 8.11757
R919 B.n613 B.n1 8.11757
R920 B.n506 B.n505 6.5566
R921 B.n493 B.n492 6.5566
R922 B.n262 B.n261 6.5566
R923 B.n277 B.n276 6.5566
R924 B.n507 B.n506 4.05904
R925 B.n492 B.n491 4.05904
R926 B.n261 B.n260 4.05904
R927 B.n276 B.n116 4.05904
R928 VP.n0 VP.t0 164.675
R929 VP.n0 VP.t1 118.293
R930 VP VP.n0 0.526373
R931 VTAIL.n242 VTAIL.n186 756.745
R932 VTAIL.n56 VTAIL.n0 756.745
R933 VTAIL.n180 VTAIL.n124 756.745
R934 VTAIL.n118 VTAIL.n62 756.745
R935 VTAIL.n207 VTAIL.n206 585
R936 VTAIL.n209 VTAIL.n208 585
R937 VTAIL.n202 VTAIL.n201 585
R938 VTAIL.n215 VTAIL.n214 585
R939 VTAIL.n217 VTAIL.n216 585
R940 VTAIL.n198 VTAIL.n197 585
R941 VTAIL.n224 VTAIL.n223 585
R942 VTAIL.n225 VTAIL.n196 585
R943 VTAIL.n227 VTAIL.n226 585
R944 VTAIL.n194 VTAIL.n193 585
R945 VTAIL.n233 VTAIL.n232 585
R946 VTAIL.n235 VTAIL.n234 585
R947 VTAIL.n190 VTAIL.n189 585
R948 VTAIL.n241 VTAIL.n240 585
R949 VTAIL.n243 VTAIL.n242 585
R950 VTAIL.n21 VTAIL.n20 585
R951 VTAIL.n23 VTAIL.n22 585
R952 VTAIL.n16 VTAIL.n15 585
R953 VTAIL.n29 VTAIL.n28 585
R954 VTAIL.n31 VTAIL.n30 585
R955 VTAIL.n12 VTAIL.n11 585
R956 VTAIL.n38 VTAIL.n37 585
R957 VTAIL.n39 VTAIL.n10 585
R958 VTAIL.n41 VTAIL.n40 585
R959 VTAIL.n8 VTAIL.n7 585
R960 VTAIL.n47 VTAIL.n46 585
R961 VTAIL.n49 VTAIL.n48 585
R962 VTAIL.n4 VTAIL.n3 585
R963 VTAIL.n55 VTAIL.n54 585
R964 VTAIL.n57 VTAIL.n56 585
R965 VTAIL.n181 VTAIL.n180 585
R966 VTAIL.n179 VTAIL.n178 585
R967 VTAIL.n128 VTAIL.n127 585
R968 VTAIL.n173 VTAIL.n172 585
R969 VTAIL.n171 VTAIL.n170 585
R970 VTAIL.n132 VTAIL.n131 585
R971 VTAIL.n136 VTAIL.n134 585
R972 VTAIL.n165 VTAIL.n164 585
R973 VTAIL.n163 VTAIL.n162 585
R974 VTAIL.n138 VTAIL.n137 585
R975 VTAIL.n157 VTAIL.n156 585
R976 VTAIL.n155 VTAIL.n154 585
R977 VTAIL.n142 VTAIL.n141 585
R978 VTAIL.n149 VTAIL.n148 585
R979 VTAIL.n147 VTAIL.n146 585
R980 VTAIL.n119 VTAIL.n118 585
R981 VTAIL.n117 VTAIL.n116 585
R982 VTAIL.n66 VTAIL.n65 585
R983 VTAIL.n111 VTAIL.n110 585
R984 VTAIL.n109 VTAIL.n108 585
R985 VTAIL.n70 VTAIL.n69 585
R986 VTAIL.n74 VTAIL.n72 585
R987 VTAIL.n103 VTAIL.n102 585
R988 VTAIL.n101 VTAIL.n100 585
R989 VTAIL.n76 VTAIL.n75 585
R990 VTAIL.n95 VTAIL.n94 585
R991 VTAIL.n93 VTAIL.n92 585
R992 VTAIL.n80 VTAIL.n79 585
R993 VTAIL.n87 VTAIL.n86 585
R994 VTAIL.n85 VTAIL.n84 585
R995 VTAIL.n205 VTAIL.t0 329.036
R996 VTAIL.n19 VTAIL.t1 329.036
R997 VTAIL.n145 VTAIL.t2 329.036
R998 VTAIL.n83 VTAIL.t3 329.036
R999 VTAIL.n208 VTAIL.n207 171.744
R1000 VTAIL.n208 VTAIL.n201 171.744
R1001 VTAIL.n215 VTAIL.n201 171.744
R1002 VTAIL.n216 VTAIL.n215 171.744
R1003 VTAIL.n216 VTAIL.n197 171.744
R1004 VTAIL.n224 VTAIL.n197 171.744
R1005 VTAIL.n225 VTAIL.n224 171.744
R1006 VTAIL.n226 VTAIL.n225 171.744
R1007 VTAIL.n226 VTAIL.n193 171.744
R1008 VTAIL.n233 VTAIL.n193 171.744
R1009 VTAIL.n234 VTAIL.n233 171.744
R1010 VTAIL.n234 VTAIL.n189 171.744
R1011 VTAIL.n241 VTAIL.n189 171.744
R1012 VTAIL.n242 VTAIL.n241 171.744
R1013 VTAIL.n22 VTAIL.n21 171.744
R1014 VTAIL.n22 VTAIL.n15 171.744
R1015 VTAIL.n29 VTAIL.n15 171.744
R1016 VTAIL.n30 VTAIL.n29 171.744
R1017 VTAIL.n30 VTAIL.n11 171.744
R1018 VTAIL.n38 VTAIL.n11 171.744
R1019 VTAIL.n39 VTAIL.n38 171.744
R1020 VTAIL.n40 VTAIL.n39 171.744
R1021 VTAIL.n40 VTAIL.n7 171.744
R1022 VTAIL.n47 VTAIL.n7 171.744
R1023 VTAIL.n48 VTAIL.n47 171.744
R1024 VTAIL.n48 VTAIL.n3 171.744
R1025 VTAIL.n55 VTAIL.n3 171.744
R1026 VTAIL.n56 VTAIL.n55 171.744
R1027 VTAIL.n180 VTAIL.n179 171.744
R1028 VTAIL.n179 VTAIL.n127 171.744
R1029 VTAIL.n172 VTAIL.n127 171.744
R1030 VTAIL.n172 VTAIL.n171 171.744
R1031 VTAIL.n171 VTAIL.n131 171.744
R1032 VTAIL.n136 VTAIL.n131 171.744
R1033 VTAIL.n164 VTAIL.n136 171.744
R1034 VTAIL.n164 VTAIL.n163 171.744
R1035 VTAIL.n163 VTAIL.n137 171.744
R1036 VTAIL.n156 VTAIL.n137 171.744
R1037 VTAIL.n156 VTAIL.n155 171.744
R1038 VTAIL.n155 VTAIL.n141 171.744
R1039 VTAIL.n148 VTAIL.n141 171.744
R1040 VTAIL.n148 VTAIL.n147 171.744
R1041 VTAIL.n118 VTAIL.n117 171.744
R1042 VTAIL.n117 VTAIL.n65 171.744
R1043 VTAIL.n110 VTAIL.n65 171.744
R1044 VTAIL.n110 VTAIL.n109 171.744
R1045 VTAIL.n109 VTAIL.n69 171.744
R1046 VTAIL.n74 VTAIL.n69 171.744
R1047 VTAIL.n102 VTAIL.n74 171.744
R1048 VTAIL.n102 VTAIL.n101 171.744
R1049 VTAIL.n101 VTAIL.n75 171.744
R1050 VTAIL.n94 VTAIL.n75 171.744
R1051 VTAIL.n94 VTAIL.n93 171.744
R1052 VTAIL.n93 VTAIL.n79 171.744
R1053 VTAIL.n86 VTAIL.n79 171.744
R1054 VTAIL.n86 VTAIL.n85 171.744
R1055 VTAIL.n207 VTAIL.t0 85.8723
R1056 VTAIL.n21 VTAIL.t1 85.8723
R1057 VTAIL.n147 VTAIL.t2 85.8723
R1058 VTAIL.n85 VTAIL.t3 85.8723
R1059 VTAIL.n247 VTAIL.n246 31.0217
R1060 VTAIL.n61 VTAIL.n60 31.0217
R1061 VTAIL.n185 VTAIL.n184 31.0217
R1062 VTAIL.n123 VTAIL.n122 31.0217
R1063 VTAIL.n123 VTAIL.n61 28.6427
R1064 VTAIL.n247 VTAIL.n185 25.3927
R1065 VTAIL.n227 VTAIL.n194 13.1884
R1066 VTAIL.n41 VTAIL.n8 13.1884
R1067 VTAIL.n134 VTAIL.n132 13.1884
R1068 VTAIL.n72 VTAIL.n70 13.1884
R1069 VTAIL.n228 VTAIL.n196 12.8005
R1070 VTAIL.n232 VTAIL.n231 12.8005
R1071 VTAIL.n42 VTAIL.n10 12.8005
R1072 VTAIL.n46 VTAIL.n45 12.8005
R1073 VTAIL.n170 VTAIL.n169 12.8005
R1074 VTAIL.n166 VTAIL.n165 12.8005
R1075 VTAIL.n108 VTAIL.n107 12.8005
R1076 VTAIL.n104 VTAIL.n103 12.8005
R1077 VTAIL.n223 VTAIL.n222 12.0247
R1078 VTAIL.n235 VTAIL.n192 12.0247
R1079 VTAIL.n37 VTAIL.n36 12.0247
R1080 VTAIL.n49 VTAIL.n6 12.0247
R1081 VTAIL.n173 VTAIL.n130 12.0247
R1082 VTAIL.n162 VTAIL.n135 12.0247
R1083 VTAIL.n111 VTAIL.n68 12.0247
R1084 VTAIL.n100 VTAIL.n73 12.0247
R1085 VTAIL.n221 VTAIL.n198 11.249
R1086 VTAIL.n236 VTAIL.n190 11.249
R1087 VTAIL.n35 VTAIL.n12 11.249
R1088 VTAIL.n50 VTAIL.n4 11.249
R1089 VTAIL.n174 VTAIL.n128 11.249
R1090 VTAIL.n161 VTAIL.n138 11.249
R1091 VTAIL.n112 VTAIL.n66 11.249
R1092 VTAIL.n99 VTAIL.n76 11.249
R1093 VTAIL.n206 VTAIL.n205 10.7239
R1094 VTAIL.n20 VTAIL.n19 10.7239
R1095 VTAIL.n146 VTAIL.n145 10.7239
R1096 VTAIL.n84 VTAIL.n83 10.7239
R1097 VTAIL.n218 VTAIL.n217 10.4732
R1098 VTAIL.n240 VTAIL.n239 10.4732
R1099 VTAIL.n32 VTAIL.n31 10.4732
R1100 VTAIL.n54 VTAIL.n53 10.4732
R1101 VTAIL.n178 VTAIL.n177 10.4732
R1102 VTAIL.n158 VTAIL.n157 10.4732
R1103 VTAIL.n116 VTAIL.n115 10.4732
R1104 VTAIL.n96 VTAIL.n95 10.4732
R1105 VTAIL.n214 VTAIL.n200 9.69747
R1106 VTAIL.n243 VTAIL.n188 9.69747
R1107 VTAIL.n28 VTAIL.n14 9.69747
R1108 VTAIL.n57 VTAIL.n2 9.69747
R1109 VTAIL.n181 VTAIL.n126 9.69747
R1110 VTAIL.n154 VTAIL.n140 9.69747
R1111 VTAIL.n119 VTAIL.n64 9.69747
R1112 VTAIL.n92 VTAIL.n78 9.69747
R1113 VTAIL.n246 VTAIL.n245 9.45567
R1114 VTAIL.n60 VTAIL.n59 9.45567
R1115 VTAIL.n184 VTAIL.n183 9.45567
R1116 VTAIL.n122 VTAIL.n121 9.45567
R1117 VTAIL.n245 VTAIL.n244 9.3005
R1118 VTAIL.n188 VTAIL.n187 9.3005
R1119 VTAIL.n239 VTAIL.n238 9.3005
R1120 VTAIL.n237 VTAIL.n236 9.3005
R1121 VTAIL.n192 VTAIL.n191 9.3005
R1122 VTAIL.n231 VTAIL.n230 9.3005
R1123 VTAIL.n204 VTAIL.n203 9.3005
R1124 VTAIL.n211 VTAIL.n210 9.3005
R1125 VTAIL.n213 VTAIL.n212 9.3005
R1126 VTAIL.n200 VTAIL.n199 9.3005
R1127 VTAIL.n219 VTAIL.n218 9.3005
R1128 VTAIL.n221 VTAIL.n220 9.3005
R1129 VTAIL.n222 VTAIL.n195 9.3005
R1130 VTAIL.n229 VTAIL.n228 9.3005
R1131 VTAIL.n59 VTAIL.n58 9.3005
R1132 VTAIL.n2 VTAIL.n1 9.3005
R1133 VTAIL.n53 VTAIL.n52 9.3005
R1134 VTAIL.n51 VTAIL.n50 9.3005
R1135 VTAIL.n6 VTAIL.n5 9.3005
R1136 VTAIL.n45 VTAIL.n44 9.3005
R1137 VTAIL.n18 VTAIL.n17 9.3005
R1138 VTAIL.n25 VTAIL.n24 9.3005
R1139 VTAIL.n27 VTAIL.n26 9.3005
R1140 VTAIL.n14 VTAIL.n13 9.3005
R1141 VTAIL.n33 VTAIL.n32 9.3005
R1142 VTAIL.n35 VTAIL.n34 9.3005
R1143 VTAIL.n36 VTAIL.n9 9.3005
R1144 VTAIL.n43 VTAIL.n42 9.3005
R1145 VTAIL.n144 VTAIL.n143 9.3005
R1146 VTAIL.n151 VTAIL.n150 9.3005
R1147 VTAIL.n153 VTAIL.n152 9.3005
R1148 VTAIL.n140 VTAIL.n139 9.3005
R1149 VTAIL.n159 VTAIL.n158 9.3005
R1150 VTAIL.n161 VTAIL.n160 9.3005
R1151 VTAIL.n135 VTAIL.n133 9.3005
R1152 VTAIL.n167 VTAIL.n166 9.3005
R1153 VTAIL.n183 VTAIL.n182 9.3005
R1154 VTAIL.n126 VTAIL.n125 9.3005
R1155 VTAIL.n177 VTAIL.n176 9.3005
R1156 VTAIL.n175 VTAIL.n174 9.3005
R1157 VTAIL.n130 VTAIL.n129 9.3005
R1158 VTAIL.n169 VTAIL.n168 9.3005
R1159 VTAIL.n82 VTAIL.n81 9.3005
R1160 VTAIL.n89 VTAIL.n88 9.3005
R1161 VTAIL.n91 VTAIL.n90 9.3005
R1162 VTAIL.n78 VTAIL.n77 9.3005
R1163 VTAIL.n97 VTAIL.n96 9.3005
R1164 VTAIL.n99 VTAIL.n98 9.3005
R1165 VTAIL.n73 VTAIL.n71 9.3005
R1166 VTAIL.n105 VTAIL.n104 9.3005
R1167 VTAIL.n121 VTAIL.n120 9.3005
R1168 VTAIL.n64 VTAIL.n63 9.3005
R1169 VTAIL.n115 VTAIL.n114 9.3005
R1170 VTAIL.n113 VTAIL.n112 9.3005
R1171 VTAIL.n68 VTAIL.n67 9.3005
R1172 VTAIL.n107 VTAIL.n106 9.3005
R1173 VTAIL.n213 VTAIL.n202 8.92171
R1174 VTAIL.n244 VTAIL.n186 8.92171
R1175 VTAIL.n27 VTAIL.n16 8.92171
R1176 VTAIL.n58 VTAIL.n0 8.92171
R1177 VTAIL.n182 VTAIL.n124 8.92171
R1178 VTAIL.n153 VTAIL.n142 8.92171
R1179 VTAIL.n120 VTAIL.n62 8.92171
R1180 VTAIL.n91 VTAIL.n80 8.92171
R1181 VTAIL.n210 VTAIL.n209 8.14595
R1182 VTAIL.n24 VTAIL.n23 8.14595
R1183 VTAIL.n150 VTAIL.n149 8.14595
R1184 VTAIL.n88 VTAIL.n87 8.14595
R1185 VTAIL.n206 VTAIL.n204 7.3702
R1186 VTAIL.n20 VTAIL.n18 7.3702
R1187 VTAIL.n146 VTAIL.n144 7.3702
R1188 VTAIL.n84 VTAIL.n82 7.3702
R1189 VTAIL.n209 VTAIL.n204 5.81868
R1190 VTAIL.n23 VTAIL.n18 5.81868
R1191 VTAIL.n149 VTAIL.n144 5.81868
R1192 VTAIL.n87 VTAIL.n82 5.81868
R1193 VTAIL.n210 VTAIL.n202 5.04292
R1194 VTAIL.n246 VTAIL.n186 5.04292
R1195 VTAIL.n24 VTAIL.n16 5.04292
R1196 VTAIL.n60 VTAIL.n0 5.04292
R1197 VTAIL.n184 VTAIL.n124 5.04292
R1198 VTAIL.n150 VTAIL.n142 5.04292
R1199 VTAIL.n122 VTAIL.n62 5.04292
R1200 VTAIL.n88 VTAIL.n80 5.04292
R1201 VTAIL.n214 VTAIL.n213 4.26717
R1202 VTAIL.n244 VTAIL.n243 4.26717
R1203 VTAIL.n28 VTAIL.n27 4.26717
R1204 VTAIL.n58 VTAIL.n57 4.26717
R1205 VTAIL.n182 VTAIL.n181 4.26717
R1206 VTAIL.n154 VTAIL.n153 4.26717
R1207 VTAIL.n120 VTAIL.n119 4.26717
R1208 VTAIL.n92 VTAIL.n91 4.26717
R1209 VTAIL.n217 VTAIL.n200 3.49141
R1210 VTAIL.n240 VTAIL.n188 3.49141
R1211 VTAIL.n31 VTAIL.n14 3.49141
R1212 VTAIL.n54 VTAIL.n2 3.49141
R1213 VTAIL.n178 VTAIL.n126 3.49141
R1214 VTAIL.n157 VTAIL.n140 3.49141
R1215 VTAIL.n116 VTAIL.n64 3.49141
R1216 VTAIL.n95 VTAIL.n78 3.49141
R1217 VTAIL.n218 VTAIL.n198 2.71565
R1218 VTAIL.n239 VTAIL.n190 2.71565
R1219 VTAIL.n32 VTAIL.n12 2.71565
R1220 VTAIL.n53 VTAIL.n4 2.71565
R1221 VTAIL.n177 VTAIL.n128 2.71565
R1222 VTAIL.n158 VTAIL.n138 2.71565
R1223 VTAIL.n115 VTAIL.n66 2.71565
R1224 VTAIL.n96 VTAIL.n76 2.71565
R1225 VTAIL.n205 VTAIL.n203 2.41282
R1226 VTAIL.n19 VTAIL.n17 2.41282
R1227 VTAIL.n145 VTAIL.n143 2.41282
R1228 VTAIL.n83 VTAIL.n81 2.41282
R1229 VTAIL.n185 VTAIL.n123 2.09533
R1230 VTAIL.n223 VTAIL.n221 1.93989
R1231 VTAIL.n236 VTAIL.n235 1.93989
R1232 VTAIL.n37 VTAIL.n35 1.93989
R1233 VTAIL.n50 VTAIL.n49 1.93989
R1234 VTAIL.n174 VTAIL.n173 1.93989
R1235 VTAIL.n162 VTAIL.n161 1.93989
R1236 VTAIL.n112 VTAIL.n111 1.93989
R1237 VTAIL.n100 VTAIL.n99 1.93989
R1238 VTAIL VTAIL.n61 1.34102
R1239 VTAIL.n222 VTAIL.n196 1.16414
R1240 VTAIL.n232 VTAIL.n192 1.16414
R1241 VTAIL.n36 VTAIL.n10 1.16414
R1242 VTAIL.n46 VTAIL.n6 1.16414
R1243 VTAIL.n170 VTAIL.n130 1.16414
R1244 VTAIL.n165 VTAIL.n135 1.16414
R1245 VTAIL.n108 VTAIL.n68 1.16414
R1246 VTAIL.n103 VTAIL.n73 1.16414
R1247 VTAIL VTAIL.n247 0.75481
R1248 VTAIL.n228 VTAIL.n227 0.388379
R1249 VTAIL.n231 VTAIL.n194 0.388379
R1250 VTAIL.n42 VTAIL.n41 0.388379
R1251 VTAIL.n45 VTAIL.n8 0.388379
R1252 VTAIL.n169 VTAIL.n132 0.388379
R1253 VTAIL.n166 VTAIL.n134 0.388379
R1254 VTAIL.n107 VTAIL.n70 0.388379
R1255 VTAIL.n104 VTAIL.n72 0.388379
R1256 VTAIL.n211 VTAIL.n203 0.155672
R1257 VTAIL.n212 VTAIL.n211 0.155672
R1258 VTAIL.n212 VTAIL.n199 0.155672
R1259 VTAIL.n219 VTAIL.n199 0.155672
R1260 VTAIL.n220 VTAIL.n219 0.155672
R1261 VTAIL.n220 VTAIL.n195 0.155672
R1262 VTAIL.n229 VTAIL.n195 0.155672
R1263 VTAIL.n230 VTAIL.n229 0.155672
R1264 VTAIL.n230 VTAIL.n191 0.155672
R1265 VTAIL.n237 VTAIL.n191 0.155672
R1266 VTAIL.n238 VTAIL.n237 0.155672
R1267 VTAIL.n238 VTAIL.n187 0.155672
R1268 VTAIL.n245 VTAIL.n187 0.155672
R1269 VTAIL.n25 VTAIL.n17 0.155672
R1270 VTAIL.n26 VTAIL.n25 0.155672
R1271 VTAIL.n26 VTAIL.n13 0.155672
R1272 VTAIL.n33 VTAIL.n13 0.155672
R1273 VTAIL.n34 VTAIL.n33 0.155672
R1274 VTAIL.n34 VTAIL.n9 0.155672
R1275 VTAIL.n43 VTAIL.n9 0.155672
R1276 VTAIL.n44 VTAIL.n43 0.155672
R1277 VTAIL.n44 VTAIL.n5 0.155672
R1278 VTAIL.n51 VTAIL.n5 0.155672
R1279 VTAIL.n52 VTAIL.n51 0.155672
R1280 VTAIL.n52 VTAIL.n1 0.155672
R1281 VTAIL.n59 VTAIL.n1 0.155672
R1282 VTAIL.n183 VTAIL.n125 0.155672
R1283 VTAIL.n176 VTAIL.n125 0.155672
R1284 VTAIL.n176 VTAIL.n175 0.155672
R1285 VTAIL.n175 VTAIL.n129 0.155672
R1286 VTAIL.n168 VTAIL.n129 0.155672
R1287 VTAIL.n168 VTAIL.n167 0.155672
R1288 VTAIL.n167 VTAIL.n133 0.155672
R1289 VTAIL.n160 VTAIL.n133 0.155672
R1290 VTAIL.n160 VTAIL.n159 0.155672
R1291 VTAIL.n159 VTAIL.n139 0.155672
R1292 VTAIL.n152 VTAIL.n139 0.155672
R1293 VTAIL.n152 VTAIL.n151 0.155672
R1294 VTAIL.n151 VTAIL.n143 0.155672
R1295 VTAIL.n121 VTAIL.n63 0.155672
R1296 VTAIL.n114 VTAIL.n63 0.155672
R1297 VTAIL.n114 VTAIL.n113 0.155672
R1298 VTAIL.n113 VTAIL.n67 0.155672
R1299 VTAIL.n106 VTAIL.n67 0.155672
R1300 VTAIL.n106 VTAIL.n105 0.155672
R1301 VTAIL.n105 VTAIL.n71 0.155672
R1302 VTAIL.n98 VTAIL.n71 0.155672
R1303 VTAIL.n98 VTAIL.n97 0.155672
R1304 VTAIL.n97 VTAIL.n77 0.155672
R1305 VTAIL.n90 VTAIL.n77 0.155672
R1306 VTAIL.n90 VTAIL.n89 0.155672
R1307 VTAIL.n89 VTAIL.n81 0.155672
R1308 VDD1.n56 VDD1.n0 756.745
R1309 VDD1.n117 VDD1.n61 756.745
R1310 VDD1.n57 VDD1.n56 585
R1311 VDD1.n55 VDD1.n54 585
R1312 VDD1.n4 VDD1.n3 585
R1313 VDD1.n49 VDD1.n48 585
R1314 VDD1.n47 VDD1.n46 585
R1315 VDD1.n8 VDD1.n7 585
R1316 VDD1.n12 VDD1.n10 585
R1317 VDD1.n41 VDD1.n40 585
R1318 VDD1.n39 VDD1.n38 585
R1319 VDD1.n14 VDD1.n13 585
R1320 VDD1.n33 VDD1.n32 585
R1321 VDD1.n31 VDD1.n30 585
R1322 VDD1.n18 VDD1.n17 585
R1323 VDD1.n25 VDD1.n24 585
R1324 VDD1.n23 VDD1.n22 585
R1325 VDD1.n82 VDD1.n81 585
R1326 VDD1.n84 VDD1.n83 585
R1327 VDD1.n77 VDD1.n76 585
R1328 VDD1.n90 VDD1.n89 585
R1329 VDD1.n92 VDD1.n91 585
R1330 VDD1.n73 VDD1.n72 585
R1331 VDD1.n99 VDD1.n98 585
R1332 VDD1.n100 VDD1.n71 585
R1333 VDD1.n102 VDD1.n101 585
R1334 VDD1.n69 VDD1.n68 585
R1335 VDD1.n108 VDD1.n107 585
R1336 VDD1.n110 VDD1.n109 585
R1337 VDD1.n65 VDD1.n64 585
R1338 VDD1.n116 VDD1.n115 585
R1339 VDD1.n118 VDD1.n117 585
R1340 VDD1.n21 VDD1.t1 329.036
R1341 VDD1.n80 VDD1.t0 329.036
R1342 VDD1.n56 VDD1.n55 171.744
R1343 VDD1.n55 VDD1.n3 171.744
R1344 VDD1.n48 VDD1.n3 171.744
R1345 VDD1.n48 VDD1.n47 171.744
R1346 VDD1.n47 VDD1.n7 171.744
R1347 VDD1.n12 VDD1.n7 171.744
R1348 VDD1.n40 VDD1.n12 171.744
R1349 VDD1.n40 VDD1.n39 171.744
R1350 VDD1.n39 VDD1.n13 171.744
R1351 VDD1.n32 VDD1.n13 171.744
R1352 VDD1.n32 VDD1.n31 171.744
R1353 VDD1.n31 VDD1.n17 171.744
R1354 VDD1.n24 VDD1.n17 171.744
R1355 VDD1.n24 VDD1.n23 171.744
R1356 VDD1.n83 VDD1.n82 171.744
R1357 VDD1.n83 VDD1.n76 171.744
R1358 VDD1.n90 VDD1.n76 171.744
R1359 VDD1.n91 VDD1.n90 171.744
R1360 VDD1.n91 VDD1.n72 171.744
R1361 VDD1.n99 VDD1.n72 171.744
R1362 VDD1.n100 VDD1.n99 171.744
R1363 VDD1.n101 VDD1.n100 171.744
R1364 VDD1.n101 VDD1.n68 171.744
R1365 VDD1.n108 VDD1.n68 171.744
R1366 VDD1.n109 VDD1.n108 171.744
R1367 VDD1.n109 VDD1.n64 171.744
R1368 VDD1.n116 VDD1.n64 171.744
R1369 VDD1.n117 VDD1.n116 171.744
R1370 VDD1 VDD1.n121 88.9731
R1371 VDD1.n23 VDD1.t1 85.8723
R1372 VDD1.n82 VDD1.t0 85.8723
R1373 VDD1 VDD1.n60 48.5712
R1374 VDD1.n10 VDD1.n8 13.1884
R1375 VDD1.n102 VDD1.n69 13.1884
R1376 VDD1.n46 VDD1.n45 12.8005
R1377 VDD1.n42 VDD1.n41 12.8005
R1378 VDD1.n103 VDD1.n71 12.8005
R1379 VDD1.n107 VDD1.n106 12.8005
R1380 VDD1.n49 VDD1.n6 12.0247
R1381 VDD1.n38 VDD1.n11 12.0247
R1382 VDD1.n98 VDD1.n97 12.0247
R1383 VDD1.n110 VDD1.n67 12.0247
R1384 VDD1.n50 VDD1.n4 11.249
R1385 VDD1.n37 VDD1.n14 11.249
R1386 VDD1.n96 VDD1.n73 11.249
R1387 VDD1.n111 VDD1.n65 11.249
R1388 VDD1.n22 VDD1.n21 10.7239
R1389 VDD1.n81 VDD1.n80 10.7239
R1390 VDD1.n54 VDD1.n53 10.4732
R1391 VDD1.n34 VDD1.n33 10.4732
R1392 VDD1.n93 VDD1.n92 10.4732
R1393 VDD1.n115 VDD1.n114 10.4732
R1394 VDD1.n57 VDD1.n2 9.69747
R1395 VDD1.n30 VDD1.n16 9.69747
R1396 VDD1.n89 VDD1.n75 9.69747
R1397 VDD1.n118 VDD1.n63 9.69747
R1398 VDD1.n60 VDD1.n59 9.45567
R1399 VDD1.n121 VDD1.n120 9.45567
R1400 VDD1.n20 VDD1.n19 9.3005
R1401 VDD1.n27 VDD1.n26 9.3005
R1402 VDD1.n29 VDD1.n28 9.3005
R1403 VDD1.n16 VDD1.n15 9.3005
R1404 VDD1.n35 VDD1.n34 9.3005
R1405 VDD1.n37 VDD1.n36 9.3005
R1406 VDD1.n11 VDD1.n9 9.3005
R1407 VDD1.n43 VDD1.n42 9.3005
R1408 VDD1.n59 VDD1.n58 9.3005
R1409 VDD1.n2 VDD1.n1 9.3005
R1410 VDD1.n53 VDD1.n52 9.3005
R1411 VDD1.n51 VDD1.n50 9.3005
R1412 VDD1.n6 VDD1.n5 9.3005
R1413 VDD1.n45 VDD1.n44 9.3005
R1414 VDD1.n120 VDD1.n119 9.3005
R1415 VDD1.n63 VDD1.n62 9.3005
R1416 VDD1.n114 VDD1.n113 9.3005
R1417 VDD1.n112 VDD1.n111 9.3005
R1418 VDD1.n67 VDD1.n66 9.3005
R1419 VDD1.n106 VDD1.n105 9.3005
R1420 VDD1.n79 VDD1.n78 9.3005
R1421 VDD1.n86 VDD1.n85 9.3005
R1422 VDD1.n88 VDD1.n87 9.3005
R1423 VDD1.n75 VDD1.n74 9.3005
R1424 VDD1.n94 VDD1.n93 9.3005
R1425 VDD1.n96 VDD1.n95 9.3005
R1426 VDD1.n97 VDD1.n70 9.3005
R1427 VDD1.n104 VDD1.n103 9.3005
R1428 VDD1.n58 VDD1.n0 8.92171
R1429 VDD1.n29 VDD1.n18 8.92171
R1430 VDD1.n88 VDD1.n77 8.92171
R1431 VDD1.n119 VDD1.n61 8.92171
R1432 VDD1.n26 VDD1.n25 8.14595
R1433 VDD1.n85 VDD1.n84 8.14595
R1434 VDD1.n22 VDD1.n20 7.3702
R1435 VDD1.n81 VDD1.n79 7.3702
R1436 VDD1.n25 VDD1.n20 5.81868
R1437 VDD1.n84 VDD1.n79 5.81868
R1438 VDD1.n60 VDD1.n0 5.04292
R1439 VDD1.n26 VDD1.n18 5.04292
R1440 VDD1.n85 VDD1.n77 5.04292
R1441 VDD1.n121 VDD1.n61 5.04292
R1442 VDD1.n58 VDD1.n57 4.26717
R1443 VDD1.n30 VDD1.n29 4.26717
R1444 VDD1.n89 VDD1.n88 4.26717
R1445 VDD1.n119 VDD1.n118 4.26717
R1446 VDD1.n54 VDD1.n2 3.49141
R1447 VDD1.n33 VDD1.n16 3.49141
R1448 VDD1.n92 VDD1.n75 3.49141
R1449 VDD1.n115 VDD1.n63 3.49141
R1450 VDD1.n53 VDD1.n4 2.71565
R1451 VDD1.n34 VDD1.n14 2.71565
R1452 VDD1.n93 VDD1.n73 2.71565
R1453 VDD1.n114 VDD1.n65 2.71565
R1454 VDD1.n21 VDD1.n19 2.41282
R1455 VDD1.n80 VDD1.n78 2.41282
R1456 VDD1.n50 VDD1.n49 1.93989
R1457 VDD1.n38 VDD1.n37 1.93989
R1458 VDD1.n98 VDD1.n96 1.93989
R1459 VDD1.n111 VDD1.n110 1.93989
R1460 VDD1.n46 VDD1.n6 1.16414
R1461 VDD1.n41 VDD1.n11 1.16414
R1462 VDD1.n97 VDD1.n71 1.16414
R1463 VDD1.n107 VDD1.n67 1.16414
R1464 VDD1.n45 VDD1.n8 0.388379
R1465 VDD1.n42 VDD1.n10 0.388379
R1466 VDD1.n103 VDD1.n102 0.388379
R1467 VDD1.n106 VDD1.n69 0.388379
R1468 VDD1.n59 VDD1.n1 0.155672
R1469 VDD1.n52 VDD1.n1 0.155672
R1470 VDD1.n52 VDD1.n51 0.155672
R1471 VDD1.n51 VDD1.n5 0.155672
R1472 VDD1.n44 VDD1.n5 0.155672
R1473 VDD1.n44 VDD1.n43 0.155672
R1474 VDD1.n43 VDD1.n9 0.155672
R1475 VDD1.n36 VDD1.n9 0.155672
R1476 VDD1.n36 VDD1.n35 0.155672
R1477 VDD1.n35 VDD1.n15 0.155672
R1478 VDD1.n28 VDD1.n15 0.155672
R1479 VDD1.n28 VDD1.n27 0.155672
R1480 VDD1.n27 VDD1.n19 0.155672
R1481 VDD1.n86 VDD1.n78 0.155672
R1482 VDD1.n87 VDD1.n86 0.155672
R1483 VDD1.n87 VDD1.n74 0.155672
R1484 VDD1.n94 VDD1.n74 0.155672
R1485 VDD1.n95 VDD1.n94 0.155672
R1486 VDD1.n95 VDD1.n70 0.155672
R1487 VDD1.n104 VDD1.n70 0.155672
R1488 VDD1.n105 VDD1.n104 0.155672
R1489 VDD1.n105 VDD1.n66 0.155672
R1490 VDD1.n112 VDD1.n66 0.155672
R1491 VDD1.n113 VDD1.n112 0.155672
R1492 VDD1.n113 VDD1.n62 0.155672
R1493 VDD1.n120 VDD1.n62 0.155672
R1494 VN VN.t0 164.583
R1495 VN VN.t1 118.817
R1496 VDD2.n117 VDD2.n61 756.745
R1497 VDD2.n56 VDD2.n0 756.745
R1498 VDD2.n118 VDD2.n117 585
R1499 VDD2.n116 VDD2.n115 585
R1500 VDD2.n65 VDD2.n64 585
R1501 VDD2.n110 VDD2.n109 585
R1502 VDD2.n108 VDD2.n107 585
R1503 VDD2.n69 VDD2.n68 585
R1504 VDD2.n73 VDD2.n71 585
R1505 VDD2.n102 VDD2.n101 585
R1506 VDD2.n100 VDD2.n99 585
R1507 VDD2.n75 VDD2.n74 585
R1508 VDD2.n94 VDD2.n93 585
R1509 VDD2.n92 VDD2.n91 585
R1510 VDD2.n79 VDD2.n78 585
R1511 VDD2.n86 VDD2.n85 585
R1512 VDD2.n84 VDD2.n83 585
R1513 VDD2.n21 VDD2.n20 585
R1514 VDD2.n23 VDD2.n22 585
R1515 VDD2.n16 VDD2.n15 585
R1516 VDD2.n29 VDD2.n28 585
R1517 VDD2.n31 VDD2.n30 585
R1518 VDD2.n12 VDD2.n11 585
R1519 VDD2.n38 VDD2.n37 585
R1520 VDD2.n39 VDD2.n10 585
R1521 VDD2.n41 VDD2.n40 585
R1522 VDD2.n8 VDD2.n7 585
R1523 VDD2.n47 VDD2.n46 585
R1524 VDD2.n49 VDD2.n48 585
R1525 VDD2.n4 VDD2.n3 585
R1526 VDD2.n55 VDD2.n54 585
R1527 VDD2.n57 VDD2.n56 585
R1528 VDD2.n82 VDD2.t1 329.036
R1529 VDD2.n19 VDD2.t0 329.036
R1530 VDD2.n117 VDD2.n116 171.744
R1531 VDD2.n116 VDD2.n64 171.744
R1532 VDD2.n109 VDD2.n64 171.744
R1533 VDD2.n109 VDD2.n108 171.744
R1534 VDD2.n108 VDD2.n68 171.744
R1535 VDD2.n73 VDD2.n68 171.744
R1536 VDD2.n101 VDD2.n73 171.744
R1537 VDD2.n101 VDD2.n100 171.744
R1538 VDD2.n100 VDD2.n74 171.744
R1539 VDD2.n93 VDD2.n74 171.744
R1540 VDD2.n93 VDD2.n92 171.744
R1541 VDD2.n92 VDD2.n78 171.744
R1542 VDD2.n85 VDD2.n78 171.744
R1543 VDD2.n85 VDD2.n84 171.744
R1544 VDD2.n22 VDD2.n21 171.744
R1545 VDD2.n22 VDD2.n15 171.744
R1546 VDD2.n29 VDD2.n15 171.744
R1547 VDD2.n30 VDD2.n29 171.744
R1548 VDD2.n30 VDD2.n11 171.744
R1549 VDD2.n38 VDD2.n11 171.744
R1550 VDD2.n39 VDD2.n38 171.744
R1551 VDD2.n40 VDD2.n39 171.744
R1552 VDD2.n40 VDD2.n7 171.744
R1553 VDD2.n47 VDD2.n7 171.744
R1554 VDD2.n48 VDD2.n47 171.744
R1555 VDD2.n48 VDD2.n3 171.744
R1556 VDD2.n55 VDD2.n3 171.744
R1557 VDD2.n56 VDD2.n55 171.744
R1558 VDD2.n122 VDD2.n60 87.6358
R1559 VDD2.n84 VDD2.t1 85.8723
R1560 VDD2.n21 VDD2.t0 85.8723
R1561 VDD2.n122 VDD2.n121 47.7005
R1562 VDD2.n71 VDD2.n69 13.1884
R1563 VDD2.n41 VDD2.n8 13.1884
R1564 VDD2.n107 VDD2.n106 12.8005
R1565 VDD2.n103 VDD2.n102 12.8005
R1566 VDD2.n42 VDD2.n10 12.8005
R1567 VDD2.n46 VDD2.n45 12.8005
R1568 VDD2.n110 VDD2.n67 12.0247
R1569 VDD2.n99 VDD2.n72 12.0247
R1570 VDD2.n37 VDD2.n36 12.0247
R1571 VDD2.n49 VDD2.n6 12.0247
R1572 VDD2.n111 VDD2.n65 11.249
R1573 VDD2.n98 VDD2.n75 11.249
R1574 VDD2.n35 VDD2.n12 11.249
R1575 VDD2.n50 VDD2.n4 11.249
R1576 VDD2.n83 VDD2.n82 10.7239
R1577 VDD2.n20 VDD2.n19 10.7239
R1578 VDD2.n115 VDD2.n114 10.4732
R1579 VDD2.n95 VDD2.n94 10.4732
R1580 VDD2.n32 VDD2.n31 10.4732
R1581 VDD2.n54 VDD2.n53 10.4732
R1582 VDD2.n118 VDD2.n63 9.69747
R1583 VDD2.n91 VDD2.n77 9.69747
R1584 VDD2.n28 VDD2.n14 9.69747
R1585 VDD2.n57 VDD2.n2 9.69747
R1586 VDD2.n121 VDD2.n120 9.45567
R1587 VDD2.n60 VDD2.n59 9.45567
R1588 VDD2.n81 VDD2.n80 9.3005
R1589 VDD2.n88 VDD2.n87 9.3005
R1590 VDD2.n90 VDD2.n89 9.3005
R1591 VDD2.n77 VDD2.n76 9.3005
R1592 VDD2.n96 VDD2.n95 9.3005
R1593 VDD2.n98 VDD2.n97 9.3005
R1594 VDD2.n72 VDD2.n70 9.3005
R1595 VDD2.n104 VDD2.n103 9.3005
R1596 VDD2.n120 VDD2.n119 9.3005
R1597 VDD2.n63 VDD2.n62 9.3005
R1598 VDD2.n114 VDD2.n113 9.3005
R1599 VDD2.n112 VDD2.n111 9.3005
R1600 VDD2.n67 VDD2.n66 9.3005
R1601 VDD2.n106 VDD2.n105 9.3005
R1602 VDD2.n59 VDD2.n58 9.3005
R1603 VDD2.n2 VDD2.n1 9.3005
R1604 VDD2.n53 VDD2.n52 9.3005
R1605 VDD2.n51 VDD2.n50 9.3005
R1606 VDD2.n6 VDD2.n5 9.3005
R1607 VDD2.n45 VDD2.n44 9.3005
R1608 VDD2.n18 VDD2.n17 9.3005
R1609 VDD2.n25 VDD2.n24 9.3005
R1610 VDD2.n27 VDD2.n26 9.3005
R1611 VDD2.n14 VDD2.n13 9.3005
R1612 VDD2.n33 VDD2.n32 9.3005
R1613 VDD2.n35 VDD2.n34 9.3005
R1614 VDD2.n36 VDD2.n9 9.3005
R1615 VDD2.n43 VDD2.n42 9.3005
R1616 VDD2.n119 VDD2.n61 8.92171
R1617 VDD2.n90 VDD2.n79 8.92171
R1618 VDD2.n27 VDD2.n16 8.92171
R1619 VDD2.n58 VDD2.n0 8.92171
R1620 VDD2.n87 VDD2.n86 8.14595
R1621 VDD2.n24 VDD2.n23 8.14595
R1622 VDD2.n83 VDD2.n81 7.3702
R1623 VDD2.n20 VDD2.n18 7.3702
R1624 VDD2.n86 VDD2.n81 5.81868
R1625 VDD2.n23 VDD2.n18 5.81868
R1626 VDD2.n121 VDD2.n61 5.04292
R1627 VDD2.n87 VDD2.n79 5.04292
R1628 VDD2.n24 VDD2.n16 5.04292
R1629 VDD2.n60 VDD2.n0 5.04292
R1630 VDD2.n119 VDD2.n118 4.26717
R1631 VDD2.n91 VDD2.n90 4.26717
R1632 VDD2.n28 VDD2.n27 4.26717
R1633 VDD2.n58 VDD2.n57 4.26717
R1634 VDD2.n115 VDD2.n63 3.49141
R1635 VDD2.n94 VDD2.n77 3.49141
R1636 VDD2.n31 VDD2.n14 3.49141
R1637 VDD2.n54 VDD2.n2 3.49141
R1638 VDD2.n114 VDD2.n65 2.71565
R1639 VDD2.n95 VDD2.n75 2.71565
R1640 VDD2.n32 VDD2.n12 2.71565
R1641 VDD2.n53 VDD2.n4 2.71565
R1642 VDD2.n82 VDD2.n80 2.41282
R1643 VDD2.n19 VDD2.n17 2.41282
R1644 VDD2.n111 VDD2.n110 1.93989
R1645 VDD2.n99 VDD2.n98 1.93989
R1646 VDD2.n37 VDD2.n35 1.93989
R1647 VDD2.n50 VDD2.n49 1.93989
R1648 VDD2.n107 VDD2.n67 1.16414
R1649 VDD2.n102 VDD2.n72 1.16414
R1650 VDD2.n36 VDD2.n10 1.16414
R1651 VDD2.n46 VDD2.n6 1.16414
R1652 VDD2 VDD2.n122 0.87119
R1653 VDD2.n106 VDD2.n69 0.388379
R1654 VDD2.n103 VDD2.n71 0.388379
R1655 VDD2.n42 VDD2.n41 0.388379
R1656 VDD2.n45 VDD2.n8 0.388379
R1657 VDD2.n120 VDD2.n62 0.155672
R1658 VDD2.n113 VDD2.n62 0.155672
R1659 VDD2.n113 VDD2.n112 0.155672
R1660 VDD2.n112 VDD2.n66 0.155672
R1661 VDD2.n105 VDD2.n66 0.155672
R1662 VDD2.n105 VDD2.n104 0.155672
R1663 VDD2.n104 VDD2.n70 0.155672
R1664 VDD2.n97 VDD2.n70 0.155672
R1665 VDD2.n97 VDD2.n96 0.155672
R1666 VDD2.n96 VDD2.n76 0.155672
R1667 VDD2.n89 VDD2.n76 0.155672
R1668 VDD2.n89 VDD2.n88 0.155672
R1669 VDD2.n88 VDD2.n80 0.155672
R1670 VDD2.n25 VDD2.n17 0.155672
R1671 VDD2.n26 VDD2.n25 0.155672
R1672 VDD2.n26 VDD2.n13 0.155672
R1673 VDD2.n33 VDD2.n13 0.155672
R1674 VDD2.n34 VDD2.n33 0.155672
R1675 VDD2.n34 VDD2.n9 0.155672
R1676 VDD2.n43 VDD2.n9 0.155672
R1677 VDD2.n44 VDD2.n43 0.155672
R1678 VDD2.n44 VDD2.n5 0.155672
R1679 VDD2.n51 VDD2.n5 0.155672
R1680 VDD2.n52 VDD2.n51 0.155672
R1681 VDD2.n52 VDD2.n1 0.155672
R1682 VDD2.n59 VDD2.n1 0.155672
C0 w_n2478_n3236# VN 3.48624f
C1 w_n2478_n3236# VDD1 1.83098f
C2 VP VTAIL 2.50825f
C3 w_n2478_n3236# VTAIL 2.67563f
C4 VP w_n2478_n3236# 3.8037f
C5 VDD2 B 1.80149f
C6 VDD2 VN 2.74254f
C7 VDD2 VDD1 0.777116f
C8 B VN 1.18783f
C9 B VDD1 1.76392f
C10 VN VDD1 0.148842f
C11 VDD2 VTAIL 5.1168f
C12 VP VDD2 0.368652f
C13 B VTAIL 3.81477f
C14 VP B 1.71312f
C15 VN VTAIL 2.49403f
C16 VDD1 VTAIL 5.05971f
C17 VP VN 5.72389f
C18 VP VDD1 2.96025f
C19 VDD2 w_n2478_n3236# 1.86728f
C20 w_n2478_n3236# B 9.53133f
C21 VDD2 VSUBS 0.935153f
C22 VDD1 VSUBS 3.89082f
C23 VTAIL VSUBS 1.064528f
C24 VN VSUBS 7.95964f
C25 VP VSUBS 1.915307f
C26 B VSUBS 4.468689f
C27 w_n2478_n3236# VSUBS 98.8127f
C28 VDD2.n0 VSUBS 0.021379f
C29 VDD2.n1 VSUBS 0.020318f
C30 VDD2.n2 VSUBS 0.010918f
C31 VDD2.n3 VSUBS 0.025806f
C32 VDD2.n4 VSUBS 0.01156f
C33 VDD2.n5 VSUBS 0.020318f
C34 VDD2.n6 VSUBS 0.010918f
C35 VDD2.n7 VSUBS 0.025806f
C36 VDD2.n8 VSUBS 0.011239f
C37 VDD2.n9 VSUBS 0.020318f
C38 VDD2.n10 VSUBS 0.01156f
C39 VDD2.n11 VSUBS 0.025806f
C40 VDD2.n12 VSUBS 0.01156f
C41 VDD2.n13 VSUBS 0.020318f
C42 VDD2.n14 VSUBS 0.010918f
C43 VDD2.n15 VSUBS 0.025806f
C44 VDD2.n16 VSUBS 0.01156f
C45 VDD2.n17 VSUBS 0.939527f
C46 VDD2.n18 VSUBS 0.010918f
C47 VDD2.t0 VSUBS 0.055566f
C48 VDD2.n19 VSUBS 0.153954f
C49 VDD2.n20 VSUBS 0.019413f
C50 VDD2.n21 VSUBS 0.019355f
C51 VDD2.n22 VSUBS 0.025806f
C52 VDD2.n23 VSUBS 0.01156f
C53 VDD2.n24 VSUBS 0.010918f
C54 VDD2.n25 VSUBS 0.020318f
C55 VDD2.n26 VSUBS 0.020318f
C56 VDD2.n27 VSUBS 0.010918f
C57 VDD2.n28 VSUBS 0.01156f
C58 VDD2.n29 VSUBS 0.025806f
C59 VDD2.n30 VSUBS 0.025806f
C60 VDD2.n31 VSUBS 0.01156f
C61 VDD2.n32 VSUBS 0.010918f
C62 VDD2.n33 VSUBS 0.020318f
C63 VDD2.n34 VSUBS 0.020318f
C64 VDD2.n35 VSUBS 0.010918f
C65 VDD2.n36 VSUBS 0.010918f
C66 VDD2.n37 VSUBS 0.01156f
C67 VDD2.n38 VSUBS 0.025806f
C68 VDD2.n39 VSUBS 0.025806f
C69 VDD2.n40 VSUBS 0.025806f
C70 VDD2.n41 VSUBS 0.011239f
C71 VDD2.n42 VSUBS 0.010918f
C72 VDD2.n43 VSUBS 0.020318f
C73 VDD2.n44 VSUBS 0.020318f
C74 VDD2.n45 VSUBS 0.010918f
C75 VDD2.n46 VSUBS 0.01156f
C76 VDD2.n47 VSUBS 0.025806f
C77 VDD2.n48 VSUBS 0.025806f
C78 VDD2.n49 VSUBS 0.01156f
C79 VDD2.n50 VSUBS 0.010918f
C80 VDD2.n51 VSUBS 0.020318f
C81 VDD2.n52 VSUBS 0.020318f
C82 VDD2.n53 VSUBS 0.010918f
C83 VDD2.n54 VSUBS 0.01156f
C84 VDD2.n55 VSUBS 0.025806f
C85 VDD2.n56 VSUBS 0.059251f
C86 VDD2.n57 VSUBS 0.01156f
C87 VDD2.n58 VSUBS 0.010918f
C88 VDD2.n59 VSUBS 0.045299f
C89 VDD2.n60 VSUBS 0.628846f
C90 VDD2.n61 VSUBS 0.021379f
C91 VDD2.n62 VSUBS 0.020318f
C92 VDD2.n63 VSUBS 0.010918f
C93 VDD2.n64 VSUBS 0.025806f
C94 VDD2.n65 VSUBS 0.01156f
C95 VDD2.n66 VSUBS 0.020318f
C96 VDD2.n67 VSUBS 0.010918f
C97 VDD2.n68 VSUBS 0.025806f
C98 VDD2.n69 VSUBS 0.011239f
C99 VDD2.n70 VSUBS 0.020318f
C100 VDD2.n71 VSUBS 0.011239f
C101 VDD2.n72 VSUBS 0.010918f
C102 VDD2.n73 VSUBS 0.025806f
C103 VDD2.n74 VSUBS 0.025806f
C104 VDD2.n75 VSUBS 0.01156f
C105 VDD2.n76 VSUBS 0.020318f
C106 VDD2.n77 VSUBS 0.010918f
C107 VDD2.n78 VSUBS 0.025806f
C108 VDD2.n79 VSUBS 0.01156f
C109 VDD2.n80 VSUBS 0.939527f
C110 VDD2.n81 VSUBS 0.010918f
C111 VDD2.t1 VSUBS 0.055566f
C112 VDD2.n82 VSUBS 0.153954f
C113 VDD2.n83 VSUBS 0.019413f
C114 VDD2.n84 VSUBS 0.019355f
C115 VDD2.n85 VSUBS 0.025806f
C116 VDD2.n86 VSUBS 0.01156f
C117 VDD2.n87 VSUBS 0.010918f
C118 VDD2.n88 VSUBS 0.020318f
C119 VDD2.n89 VSUBS 0.020318f
C120 VDD2.n90 VSUBS 0.010918f
C121 VDD2.n91 VSUBS 0.01156f
C122 VDD2.n92 VSUBS 0.025806f
C123 VDD2.n93 VSUBS 0.025806f
C124 VDD2.n94 VSUBS 0.01156f
C125 VDD2.n95 VSUBS 0.010918f
C126 VDD2.n96 VSUBS 0.020318f
C127 VDD2.n97 VSUBS 0.020318f
C128 VDD2.n98 VSUBS 0.010918f
C129 VDD2.n99 VSUBS 0.01156f
C130 VDD2.n100 VSUBS 0.025806f
C131 VDD2.n101 VSUBS 0.025806f
C132 VDD2.n102 VSUBS 0.01156f
C133 VDD2.n103 VSUBS 0.010918f
C134 VDD2.n104 VSUBS 0.020318f
C135 VDD2.n105 VSUBS 0.020318f
C136 VDD2.n106 VSUBS 0.010918f
C137 VDD2.n107 VSUBS 0.01156f
C138 VDD2.n108 VSUBS 0.025806f
C139 VDD2.n109 VSUBS 0.025806f
C140 VDD2.n110 VSUBS 0.01156f
C141 VDD2.n111 VSUBS 0.010918f
C142 VDD2.n112 VSUBS 0.020318f
C143 VDD2.n113 VSUBS 0.020318f
C144 VDD2.n114 VSUBS 0.010918f
C145 VDD2.n115 VSUBS 0.01156f
C146 VDD2.n116 VSUBS 0.025806f
C147 VDD2.n117 VSUBS 0.059251f
C148 VDD2.n118 VSUBS 0.01156f
C149 VDD2.n119 VSUBS 0.010918f
C150 VDD2.n120 VSUBS 0.045299f
C151 VDD2.n121 VSUBS 0.043644f
C152 VDD2.n122 VSUBS 2.54937f
C153 VN.t1 VSUBS 4.18089f
C154 VN.t0 VSUBS 5.01663f
C155 VDD1.n0 VSUBS 0.02199f
C156 VDD1.n1 VSUBS 0.020898f
C157 VDD1.n2 VSUBS 0.01123f
C158 VDD1.n3 VSUBS 0.026543f
C159 VDD1.n4 VSUBS 0.011891f
C160 VDD1.n5 VSUBS 0.020898f
C161 VDD1.n6 VSUBS 0.01123f
C162 VDD1.n7 VSUBS 0.026543f
C163 VDD1.n8 VSUBS 0.01156f
C164 VDD1.n9 VSUBS 0.020898f
C165 VDD1.n10 VSUBS 0.01156f
C166 VDD1.n11 VSUBS 0.01123f
C167 VDD1.n12 VSUBS 0.026543f
C168 VDD1.n13 VSUBS 0.026543f
C169 VDD1.n14 VSUBS 0.011891f
C170 VDD1.n15 VSUBS 0.020898f
C171 VDD1.n16 VSUBS 0.01123f
C172 VDD1.n17 VSUBS 0.026543f
C173 VDD1.n18 VSUBS 0.011891f
C174 VDD1.n19 VSUBS 0.966365f
C175 VDD1.n20 VSUBS 0.01123f
C176 VDD1.t1 VSUBS 0.057153f
C177 VDD1.n21 VSUBS 0.158352f
C178 VDD1.n22 VSUBS 0.019967f
C179 VDD1.n23 VSUBS 0.019907f
C180 VDD1.n24 VSUBS 0.026543f
C181 VDD1.n25 VSUBS 0.011891f
C182 VDD1.n26 VSUBS 0.01123f
C183 VDD1.n27 VSUBS 0.020898f
C184 VDD1.n28 VSUBS 0.020898f
C185 VDD1.n29 VSUBS 0.01123f
C186 VDD1.n30 VSUBS 0.011891f
C187 VDD1.n31 VSUBS 0.026543f
C188 VDD1.n32 VSUBS 0.026543f
C189 VDD1.n33 VSUBS 0.011891f
C190 VDD1.n34 VSUBS 0.01123f
C191 VDD1.n35 VSUBS 0.020898f
C192 VDD1.n36 VSUBS 0.020898f
C193 VDD1.n37 VSUBS 0.01123f
C194 VDD1.n38 VSUBS 0.011891f
C195 VDD1.n39 VSUBS 0.026543f
C196 VDD1.n40 VSUBS 0.026543f
C197 VDD1.n41 VSUBS 0.011891f
C198 VDD1.n42 VSUBS 0.01123f
C199 VDD1.n43 VSUBS 0.020898f
C200 VDD1.n44 VSUBS 0.020898f
C201 VDD1.n45 VSUBS 0.01123f
C202 VDD1.n46 VSUBS 0.011891f
C203 VDD1.n47 VSUBS 0.026543f
C204 VDD1.n48 VSUBS 0.026543f
C205 VDD1.n49 VSUBS 0.011891f
C206 VDD1.n50 VSUBS 0.01123f
C207 VDD1.n51 VSUBS 0.020898f
C208 VDD1.n52 VSUBS 0.020898f
C209 VDD1.n53 VSUBS 0.01123f
C210 VDD1.n54 VSUBS 0.011891f
C211 VDD1.n55 VSUBS 0.026543f
C212 VDD1.n56 VSUBS 0.060943f
C213 VDD1.n57 VSUBS 0.011891f
C214 VDD1.n58 VSUBS 0.01123f
C215 VDD1.n59 VSUBS 0.046593f
C216 VDD1.n60 VSUBS 0.046646f
C217 VDD1.n61 VSUBS 0.02199f
C218 VDD1.n62 VSUBS 0.020898f
C219 VDD1.n63 VSUBS 0.01123f
C220 VDD1.n64 VSUBS 0.026543f
C221 VDD1.n65 VSUBS 0.011891f
C222 VDD1.n66 VSUBS 0.020898f
C223 VDD1.n67 VSUBS 0.01123f
C224 VDD1.n68 VSUBS 0.026543f
C225 VDD1.n69 VSUBS 0.01156f
C226 VDD1.n70 VSUBS 0.020898f
C227 VDD1.n71 VSUBS 0.011891f
C228 VDD1.n72 VSUBS 0.026543f
C229 VDD1.n73 VSUBS 0.011891f
C230 VDD1.n74 VSUBS 0.020898f
C231 VDD1.n75 VSUBS 0.01123f
C232 VDD1.n76 VSUBS 0.026543f
C233 VDD1.n77 VSUBS 0.011891f
C234 VDD1.n78 VSUBS 0.966366f
C235 VDD1.n79 VSUBS 0.01123f
C236 VDD1.t0 VSUBS 0.057153f
C237 VDD1.n80 VSUBS 0.158352f
C238 VDD1.n81 VSUBS 0.019967f
C239 VDD1.n82 VSUBS 0.019907f
C240 VDD1.n83 VSUBS 0.026543f
C241 VDD1.n84 VSUBS 0.011891f
C242 VDD1.n85 VSUBS 0.01123f
C243 VDD1.n86 VSUBS 0.020898f
C244 VDD1.n87 VSUBS 0.020898f
C245 VDD1.n88 VSUBS 0.01123f
C246 VDD1.n89 VSUBS 0.011891f
C247 VDD1.n90 VSUBS 0.026543f
C248 VDD1.n91 VSUBS 0.026543f
C249 VDD1.n92 VSUBS 0.011891f
C250 VDD1.n93 VSUBS 0.01123f
C251 VDD1.n94 VSUBS 0.020898f
C252 VDD1.n95 VSUBS 0.020898f
C253 VDD1.n96 VSUBS 0.01123f
C254 VDD1.n97 VSUBS 0.01123f
C255 VDD1.n98 VSUBS 0.011891f
C256 VDD1.n99 VSUBS 0.026543f
C257 VDD1.n100 VSUBS 0.026543f
C258 VDD1.n101 VSUBS 0.026543f
C259 VDD1.n102 VSUBS 0.01156f
C260 VDD1.n103 VSUBS 0.01123f
C261 VDD1.n104 VSUBS 0.020898f
C262 VDD1.n105 VSUBS 0.020898f
C263 VDD1.n106 VSUBS 0.01123f
C264 VDD1.n107 VSUBS 0.011891f
C265 VDD1.n108 VSUBS 0.026543f
C266 VDD1.n109 VSUBS 0.026543f
C267 VDD1.n110 VSUBS 0.011891f
C268 VDD1.n111 VSUBS 0.01123f
C269 VDD1.n112 VSUBS 0.020898f
C270 VDD1.n113 VSUBS 0.020898f
C271 VDD1.n114 VSUBS 0.01123f
C272 VDD1.n115 VSUBS 0.011891f
C273 VDD1.n116 VSUBS 0.026543f
C274 VDD1.n117 VSUBS 0.060943f
C275 VDD1.n118 VSUBS 0.011891f
C276 VDD1.n119 VSUBS 0.01123f
C277 VDD1.n120 VSUBS 0.046593f
C278 VDD1.n121 VSUBS 0.694117f
C279 VTAIL.n0 VSUBS 0.031991f
C280 VTAIL.n1 VSUBS 0.030403f
C281 VTAIL.n2 VSUBS 0.016337f
C282 VTAIL.n3 VSUBS 0.038616f
C283 VTAIL.n4 VSUBS 0.017298f
C284 VTAIL.n5 VSUBS 0.030403f
C285 VTAIL.n6 VSUBS 0.016337f
C286 VTAIL.n7 VSUBS 0.038616f
C287 VTAIL.n8 VSUBS 0.016818f
C288 VTAIL.n9 VSUBS 0.030403f
C289 VTAIL.n10 VSUBS 0.017298f
C290 VTAIL.n11 VSUBS 0.038616f
C291 VTAIL.n12 VSUBS 0.017298f
C292 VTAIL.n13 VSUBS 0.030403f
C293 VTAIL.n14 VSUBS 0.016337f
C294 VTAIL.n15 VSUBS 0.038616f
C295 VTAIL.n16 VSUBS 0.017298f
C296 VTAIL.n17 VSUBS 1.40588f
C297 VTAIL.n18 VSUBS 0.016337f
C298 VTAIL.t1 VSUBS 0.083147f
C299 VTAIL.n19 VSUBS 0.230373f
C300 VTAIL.n20 VSUBS 0.029049f
C301 VTAIL.n21 VSUBS 0.028962f
C302 VTAIL.n22 VSUBS 0.038616f
C303 VTAIL.n23 VSUBS 0.017298f
C304 VTAIL.n24 VSUBS 0.016337f
C305 VTAIL.n25 VSUBS 0.030403f
C306 VTAIL.n26 VSUBS 0.030403f
C307 VTAIL.n27 VSUBS 0.016337f
C308 VTAIL.n28 VSUBS 0.017298f
C309 VTAIL.n29 VSUBS 0.038616f
C310 VTAIL.n30 VSUBS 0.038616f
C311 VTAIL.n31 VSUBS 0.017298f
C312 VTAIL.n32 VSUBS 0.016337f
C313 VTAIL.n33 VSUBS 0.030403f
C314 VTAIL.n34 VSUBS 0.030403f
C315 VTAIL.n35 VSUBS 0.016337f
C316 VTAIL.n36 VSUBS 0.016337f
C317 VTAIL.n37 VSUBS 0.017298f
C318 VTAIL.n38 VSUBS 0.038616f
C319 VTAIL.n39 VSUBS 0.038616f
C320 VTAIL.n40 VSUBS 0.038616f
C321 VTAIL.n41 VSUBS 0.016818f
C322 VTAIL.n42 VSUBS 0.016337f
C323 VTAIL.n43 VSUBS 0.030403f
C324 VTAIL.n44 VSUBS 0.030403f
C325 VTAIL.n45 VSUBS 0.016337f
C326 VTAIL.n46 VSUBS 0.017298f
C327 VTAIL.n47 VSUBS 0.038616f
C328 VTAIL.n48 VSUBS 0.038616f
C329 VTAIL.n49 VSUBS 0.017298f
C330 VTAIL.n50 VSUBS 0.016337f
C331 VTAIL.n51 VSUBS 0.030403f
C332 VTAIL.n52 VSUBS 0.030403f
C333 VTAIL.n53 VSUBS 0.016337f
C334 VTAIL.n54 VSUBS 0.017298f
C335 VTAIL.n55 VSUBS 0.038616f
C336 VTAIL.n56 VSUBS 0.088661f
C337 VTAIL.n57 VSUBS 0.017298f
C338 VTAIL.n58 VSUBS 0.016337f
C339 VTAIL.n59 VSUBS 0.067784f
C340 VTAIL.n60 VSUBS 0.044295f
C341 VTAIL.n61 VSUBS 2.16337f
C342 VTAIL.n62 VSUBS 0.031991f
C343 VTAIL.n63 VSUBS 0.030403f
C344 VTAIL.n64 VSUBS 0.016337f
C345 VTAIL.n65 VSUBS 0.038616f
C346 VTAIL.n66 VSUBS 0.017298f
C347 VTAIL.n67 VSUBS 0.030403f
C348 VTAIL.n68 VSUBS 0.016337f
C349 VTAIL.n69 VSUBS 0.038616f
C350 VTAIL.n70 VSUBS 0.016818f
C351 VTAIL.n71 VSUBS 0.030403f
C352 VTAIL.n72 VSUBS 0.016818f
C353 VTAIL.n73 VSUBS 0.016337f
C354 VTAIL.n74 VSUBS 0.038616f
C355 VTAIL.n75 VSUBS 0.038616f
C356 VTAIL.n76 VSUBS 0.017298f
C357 VTAIL.n77 VSUBS 0.030403f
C358 VTAIL.n78 VSUBS 0.016337f
C359 VTAIL.n79 VSUBS 0.038616f
C360 VTAIL.n80 VSUBS 0.017298f
C361 VTAIL.n81 VSUBS 1.40588f
C362 VTAIL.n82 VSUBS 0.016337f
C363 VTAIL.t3 VSUBS 0.083147f
C364 VTAIL.n83 VSUBS 0.230373f
C365 VTAIL.n84 VSUBS 0.029049f
C366 VTAIL.n85 VSUBS 0.028962f
C367 VTAIL.n86 VSUBS 0.038616f
C368 VTAIL.n87 VSUBS 0.017298f
C369 VTAIL.n88 VSUBS 0.016337f
C370 VTAIL.n89 VSUBS 0.030403f
C371 VTAIL.n90 VSUBS 0.030403f
C372 VTAIL.n91 VSUBS 0.016337f
C373 VTAIL.n92 VSUBS 0.017298f
C374 VTAIL.n93 VSUBS 0.038616f
C375 VTAIL.n94 VSUBS 0.038616f
C376 VTAIL.n95 VSUBS 0.017298f
C377 VTAIL.n96 VSUBS 0.016337f
C378 VTAIL.n97 VSUBS 0.030403f
C379 VTAIL.n98 VSUBS 0.030403f
C380 VTAIL.n99 VSUBS 0.016337f
C381 VTAIL.n100 VSUBS 0.017298f
C382 VTAIL.n101 VSUBS 0.038616f
C383 VTAIL.n102 VSUBS 0.038616f
C384 VTAIL.n103 VSUBS 0.017298f
C385 VTAIL.n104 VSUBS 0.016337f
C386 VTAIL.n105 VSUBS 0.030403f
C387 VTAIL.n106 VSUBS 0.030403f
C388 VTAIL.n107 VSUBS 0.016337f
C389 VTAIL.n108 VSUBS 0.017298f
C390 VTAIL.n109 VSUBS 0.038616f
C391 VTAIL.n110 VSUBS 0.038616f
C392 VTAIL.n111 VSUBS 0.017298f
C393 VTAIL.n112 VSUBS 0.016337f
C394 VTAIL.n113 VSUBS 0.030403f
C395 VTAIL.n114 VSUBS 0.030403f
C396 VTAIL.n115 VSUBS 0.016337f
C397 VTAIL.n116 VSUBS 0.017298f
C398 VTAIL.n117 VSUBS 0.038616f
C399 VTAIL.n118 VSUBS 0.088661f
C400 VTAIL.n119 VSUBS 0.017298f
C401 VTAIL.n120 VSUBS 0.016337f
C402 VTAIL.n121 VSUBS 0.067784f
C403 VTAIL.n122 VSUBS 0.044295f
C404 VTAIL.n123 VSUBS 2.23726f
C405 VTAIL.n124 VSUBS 0.031991f
C406 VTAIL.n125 VSUBS 0.030403f
C407 VTAIL.n126 VSUBS 0.016337f
C408 VTAIL.n127 VSUBS 0.038616f
C409 VTAIL.n128 VSUBS 0.017298f
C410 VTAIL.n129 VSUBS 0.030403f
C411 VTAIL.n130 VSUBS 0.016337f
C412 VTAIL.n131 VSUBS 0.038616f
C413 VTAIL.n132 VSUBS 0.016818f
C414 VTAIL.n133 VSUBS 0.030403f
C415 VTAIL.n134 VSUBS 0.016818f
C416 VTAIL.n135 VSUBS 0.016337f
C417 VTAIL.n136 VSUBS 0.038616f
C418 VTAIL.n137 VSUBS 0.038616f
C419 VTAIL.n138 VSUBS 0.017298f
C420 VTAIL.n139 VSUBS 0.030403f
C421 VTAIL.n140 VSUBS 0.016337f
C422 VTAIL.n141 VSUBS 0.038616f
C423 VTAIL.n142 VSUBS 0.017298f
C424 VTAIL.n143 VSUBS 1.40588f
C425 VTAIL.n144 VSUBS 0.016337f
C426 VTAIL.t2 VSUBS 0.083147f
C427 VTAIL.n145 VSUBS 0.230373f
C428 VTAIL.n146 VSUBS 0.029049f
C429 VTAIL.n147 VSUBS 0.028962f
C430 VTAIL.n148 VSUBS 0.038616f
C431 VTAIL.n149 VSUBS 0.017298f
C432 VTAIL.n150 VSUBS 0.016337f
C433 VTAIL.n151 VSUBS 0.030403f
C434 VTAIL.n152 VSUBS 0.030403f
C435 VTAIL.n153 VSUBS 0.016337f
C436 VTAIL.n154 VSUBS 0.017298f
C437 VTAIL.n155 VSUBS 0.038616f
C438 VTAIL.n156 VSUBS 0.038616f
C439 VTAIL.n157 VSUBS 0.017298f
C440 VTAIL.n158 VSUBS 0.016337f
C441 VTAIL.n159 VSUBS 0.030403f
C442 VTAIL.n160 VSUBS 0.030403f
C443 VTAIL.n161 VSUBS 0.016337f
C444 VTAIL.n162 VSUBS 0.017298f
C445 VTAIL.n163 VSUBS 0.038616f
C446 VTAIL.n164 VSUBS 0.038616f
C447 VTAIL.n165 VSUBS 0.017298f
C448 VTAIL.n166 VSUBS 0.016337f
C449 VTAIL.n167 VSUBS 0.030403f
C450 VTAIL.n168 VSUBS 0.030403f
C451 VTAIL.n169 VSUBS 0.016337f
C452 VTAIL.n170 VSUBS 0.017298f
C453 VTAIL.n171 VSUBS 0.038616f
C454 VTAIL.n172 VSUBS 0.038616f
C455 VTAIL.n173 VSUBS 0.017298f
C456 VTAIL.n174 VSUBS 0.016337f
C457 VTAIL.n175 VSUBS 0.030403f
C458 VTAIL.n176 VSUBS 0.030403f
C459 VTAIL.n177 VSUBS 0.016337f
C460 VTAIL.n178 VSUBS 0.017298f
C461 VTAIL.n179 VSUBS 0.038616f
C462 VTAIL.n180 VSUBS 0.088661f
C463 VTAIL.n181 VSUBS 0.017298f
C464 VTAIL.n182 VSUBS 0.016337f
C465 VTAIL.n183 VSUBS 0.067784f
C466 VTAIL.n184 VSUBS 0.044295f
C467 VTAIL.n185 VSUBS 1.91887f
C468 VTAIL.n186 VSUBS 0.031991f
C469 VTAIL.n187 VSUBS 0.030403f
C470 VTAIL.n188 VSUBS 0.016337f
C471 VTAIL.n189 VSUBS 0.038616f
C472 VTAIL.n190 VSUBS 0.017298f
C473 VTAIL.n191 VSUBS 0.030403f
C474 VTAIL.n192 VSUBS 0.016337f
C475 VTAIL.n193 VSUBS 0.038616f
C476 VTAIL.n194 VSUBS 0.016818f
C477 VTAIL.n195 VSUBS 0.030403f
C478 VTAIL.n196 VSUBS 0.017298f
C479 VTAIL.n197 VSUBS 0.038616f
C480 VTAIL.n198 VSUBS 0.017298f
C481 VTAIL.n199 VSUBS 0.030403f
C482 VTAIL.n200 VSUBS 0.016337f
C483 VTAIL.n201 VSUBS 0.038616f
C484 VTAIL.n202 VSUBS 0.017298f
C485 VTAIL.n203 VSUBS 1.40588f
C486 VTAIL.n204 VSUBS 0.016337f
C487 VTAIL.t0 VSUBS 0.083147f
C488 VTAIL.n205 VSUBS 0.230373f
C489 VTAIL.n206 VSUBS 0.029049f
C490 VTAIL.n207 VSUBS 0.028962f
C491 VTAIL.n208 VSUBS 0.038616f
C492 VTAIL.n209 VSUBS 0.017298f
C493 VTAIL.n210 VSUBS 0.016337f
C494 VTAIL.n211 VSUBS 0.030403f
C495 VTAIL.n212 VSUBS 0.030403f
C496 VTAIL.n213 VSUBS 0.016337f
C497 VTAIL.n214 VSUBS 0.017298f
C498 VTAIL.n215 VSUBS 0.038616f
C499 VTAIL.n216 VSUBS 0.038616f
C500 VTAIL.n217 VSUBS 0.017298f
C501 VTAIL.n218 VSUBS 0.016337f
C502 VTAIL.n219 VSUBS 0.030403f
C503 VTAIL.n220 VSUBS 0.030403f
C504 VTAIL.n221 VSUBS 0.016337f
C505 VTAIL.n222 VSUBS 0.016337f
C506 VTAIL.n223 VSUBS 0.017298f
C507 VTAIL.n224 VSUBS 0.038616f
C508 VTAIL.n225 VSUBS 0.038616f
C509 VTAIL.n226 VSUBS 0.038616f
C510 VTAIL.n227 VSUBS 0.016818f
C511 VTAIL.n228 VSUBS 0.016337f
C512 VTAIL.n229 VSUBS 0.030403f
C513 VTAIL.n230 VSUBS 0.030403f
C514 VTAIL.n231 VSUBS 0.016337f
C515 VTAIL.n232 VSUBS 0.017298f
C516 VTAIL.n233 VSUBS 0.038616f
C517 VTAIL.n234 VSUBS 0.038616f
C518 VTAIL.n235 VSUBS 0.017298f
C519 VTAIL.n236 VSUBS 0.016337f
C520 VTAIL.n237 VSUBS 0.030403f
C521 VTAIL.n238 VSUBS 0.030403f
C522 VTAIL.n239 VSUBS 0.016337f
C523 VTAIL.n240 VSUBS 0.017298f
C524 VTAIL.n241 VSUBS 0.038616f
C525 VTAIL.n242 VSUBS 0.088661f
C526 VTAIL.n243 VSUBS 0.017298f
C527 VTAIL.n244 VSUBS 0.016337f
C528 VTAIL.n245 VSUBS 0.067784f
C529 VTAIL.n246 VSUBS 0.044295f
C530 VTAIL.n247 VSUBS 1.78755f
C531 VP.t0 VSUBS 5.243279f
C532 VP.t1 VSUBS 4.36387f
C533 VP.n0 VSUBS 5.2607f
C534 B.n0 VSUBS 0.005164f
C535 B.n1 VSUBS 0.005164f
C536 B.n2 VSUBS 0.007637f
C537 B.n3 VSUBS 0.005852f
C538 B.n4 VSUBS 0.005852f
C539 B.n5 VSUBS 0.005852f
C540 B.n6 VSUBS 0.005852f
C541 B.n7 VSUBS 0.005852f
C542 B.n8 VSUBS 0.005852f
C543 B.n9 VSUBS 0.005852f
C544 B.n10 VSUBS 0.005852f
C545 B.n11 VSUBS 0.005852f
C546 B.n12 VSUBS 0.005852f
C547 B.n13 VSUBS 0.005852f
C548 B.n14 VSUBS 0.005852f
C549 B.n15 VSUBS 0.005852f
C550 B.n16 VSUBS 0.005852f
C551 B.n17 VSUBS 0.013159f
C552 B.n18 VSUBS 0.005852f
C553 B.n19 VSUBS 0.005852f
C554 B.n20 VSUBS 0.005852f
C555 B.n21 VSUBS 0.005852f
C556 B.n22 VSUBS 0.005852f
C557 B.n23 VSUBS 0.005852f
C558 B.n24 VSUBS 0.005852f
C559 B.n25 VSUBS 0.005852f
C560 B.n26 VSUBS 0.005852f
C561 B.n27 VSUBS 0.005852f
C562 B.n28 VSUBS 0.005852f
C563 B.n29 VSUBS 0.005852f
C564 B.n30 VSUBS 0.005852f
C565 B.n31 VSUBS 0.005852f
C566 B.n32 VSUBS 0.005852f
C567 B.n33 VSUBS 0.005852f
C568 B.n34 VSUBS 0.005852f
C569 B.n35 VSUBS 0.005852f
C570 B.n36 VSUBS 0.005852f
C571 B.n37 VSUBS 0.005852f
C572 B.t4 VSUBS 0.164154f
C573 B.t5 VSUBS 0.197201f
C574 B.t3 VSUBS 1.51687f
C575 B.n38 VSUBS 0.315848f
C576 B.n39 VSUBS 0.205766f
C577 B.n40 VSUBS 0.005852f
C578 B.n41 VSUBS 0.005852f
C579 B.n42 VSUBS 0.005852f
C580 B.n43 VSUBS 0.005852f
C581 B.t7 VSUBS 0.164156f
C582 B.t8 VSUBS 0.197203f
C583 B.t6 VSUBS 1.51687f
C584 B.n44 VSUBS 0.315846f
C585 B.n45 VSUBS 0.205763f
C586 B.n46 VSUBS 0.005852f
C587 B.n47 VSUBS 0.005852f
C588 B.n48 VSUBS 0.005852f
C589 B.n49 VSUBS 0.005852f
C590 B.n50 VSUBS 0.005852f
C591 B.n51 VSUBS 0.005852f
C592 B.n52 VSUBS 0.005852f
C593 B.n53 VSUBS 0.005852f
C594 B.n54 VSUBS 0.005852f
C595 B.n55 VSUBS 0.005852f
C596 B.n56 VSUBS 0.005852f
C597 B.n57 VSUBS 0.005852f
C598 B.n58 VSUBS 0.005852f
C599 B.n59 VSUBS 0.005852f
C600 B.n60 VSUBS 0.005852f
C601 B.n61 VSUBS 0.005852f
C602 B.n62 VSUBS 0.005852f
C603 B.n63 VSUBS 0.005852f
C604 B.n64 VSUBS 0.005852f
C605 B.n65 VSUBS 0.013159f
C606 B.n66 VSUBS 0.005852f
C607 B.n67 VSUBS 0.005852f
C608 B.n68 VSUBS 0.005852f
C609 B.n69 VSUBS 0.005852f
C610 B.n70 VSUBS 0.005852f
C611 B.n71 VSUBS 0.005852f
C612 B.n72 VSUBS 0.005852f
C613 B.n73 VSUBS 0.005852f
C614 B.n74 VSUBS 0.005852f
C615 B.n75 VSUBS 0.005852f
C616 B.n76 VSUBS 0.005852f
C617 B.n77 VSUBS 0.005852f
C618 B.n78 VSUBS 0.005852f
C619 B.n79 VSUBS 0.005852f
C620 B.n80 VSUBS 0.005852f
C621 B.n81 VSUBS 0.005852f
C622 B.n82 VSUBS 0.005852f
C623 B.n83 VSUBS 0.005852f
C624 B.n84 VSUBS 0.005852f
C625 B.n85 VSUBS 0.005852f
C626 B.n86 VSUBS 0.005852f
C627 B.n87 VSUBS 0.005852f
C628 B.n88 VSUBS 0.005852f
C629 B.n89 VSUBS 0.005852f
C630 B.n90 VSUBS 0.005852f
C631 B.n91 VSUBS 0.005852f
C632 B.n92 VSUBS 0.005852f
C633 B.n93 VSUBS 0.005852f
C634 B.n94 VSUBS 0.005852f
C635 B.n95 VSUBS 0.005852f
C636 B.n96 VSUBS 0.013417f
C637 B.n97 VSUBS 0.005852f
C638 B.n98 VSUBS 0.005852f
C639 B.n99 VSUBS 0.005852f
C640 B.n100 VSUBS 0.005852f
C641 B.n101 VSUBS 0.005852f
C642 B.n102 VSUBS 0.005852f
C643 B.n103 VSUBS 0.005852f
C644 B.n104 VSUBS 0.005852f
C645 B.n105 VSUBS 0.005852f
C646 B.n106 VSUBS 0.005852f
C647 B.n107 VSUBS 0.005852f
C648 B.n108 VSUBS 0.005852f
C649 B.n109 VSUBS 0.005852f
C650 B.n110 VSUBS 0.005852f
C651 B.n111 VSUBS 0.005852f
C652 B.n112 VSUBS 0.005852f
C653 B.n113 VSUBS 0.005852f
C654 B.n114 VSUBS 0.005852f
C655 B.n115 VSUBS 0.005852f
C656 B.n116 VSUBS 0.004045f
C657 B.n117 VSUBS 0.005852f
C658 B.n118 VSUBS 0.005852f
C659 B.n119 VSUBS 0.005852f
C660 B.n120 VSUBS 0.005852f
C661 B.n121 VSUBS 0.005852f
C662 B.t11 VSUBS 0.164154f
C663 B.t10 VSUBS 0.197201f
C664 B.t9 VSUBS 1.51687f
C665 B.n122 VSUBS 0.315848f
C666 B.n123 VSUBS 0.205766f
C667 B.n124 VSUBS 0.005852f
C668 B.n125 VSUBS 0.005852f
C669 B.n126 VSUBS 0.005852f
C670 B.n127 VSUBS 0.005852f
C671 B.n128 VSUBS 0.005852f
C672 B.n129 VSUBS 0.005852f
C673 B.n130 VSUBS 0.005852f
C674 B.n131 VSUBS 0.005852f
C675 B.n132 VSUBS 0.005852f
C676 B.n133 VSUBS 0.005852f
C677 B.n134 VSUBS 0.005852f
C678 B.n135 VSUBS 0.005852f
C679 B.n136 VSUBS 0.005852f
C680 B.n137 VSUBS 0.005852f
C681 B.n138 VSUBS 0.005852f
C682 B.n139 VSUBS 0.005852f
C683 B.n140 VSUBS 0.005852f
C684 B.n141 VSUBS 0.005852f
C685 B.n142 VSUBS 0.005852f
C686 B.n143 VSUBS 0.01266f
C687 B.n144 VSUBS 0.005852f
C688 B.n145 VSUBS 0.005852f
C689 B.n146 VSUBS 0.005852f
C690 B.n147 VSUBS 0.005852f
C691 B.n148 VSUBS 0.005852f
C692 B.n149 VSUBS 0.005852f
C693 B.n150 VSUBS 0.005852f
C694 B.n151 VSUBS 0.005852f
C695 B.n152 VSUBS 0.005852f
C696 B.n153 VSUBS 0.005852f
C697 B.n154 VSUBS 0.005852f
C698 B.n155 VSUBS 0.005852f
C699 B.n156 VSUBS 0.005852f
C700 B.n157 VSUBS 0.005852f
C701 B.n158 VSUBS 0.005852f
C702 B.n159 VSUBS 0.005852f
C703 B.n160 VSUBS 0.005852f
C704 B.n161 VSUBS 0.005852f
C705 B.n162 VSUBS 0.005852f
C706 B.n163 VSUBS 0.005852f
C707 B.n164 VSUBS 0.005852f
C708 B.n165 VSUBS 0.005852f
C709 B.n166 VSUBS 0.005852f
C710 B.n167 VSUBS 0.005852f
C711 B.n168 VSUBS 0.005852f
C712 B.n169 VSUBS 0.005852f
C713 B.n170 VSUBS 0.005852f
C714 B.n171 VSUBS 0.005852f
C715 B.n172 VSUBS 0.005852f
C716 B.n173 VSUBS 0.005852f
C717 B.n174 VSUBS 0.005852f
C718 B.n175 VSUBS 0.005852f
C719 B.n176 VSUBS 0.005852f
C720 B.n177 VSUBS 0.005852f
C721 B.n178 VSUBS 0.005852f
C722 B.n179 VSUBS 0.005852f
C723 B.n180 VSUBS 0.005852f
C724 B.n181 VSUBS 0.005852f
C725 B.n182 VSUBS 0.005852f
C726 B.n183 VSUBS 0.005852f
C727 B.n184 VSUBS 0.005852f
C728 B.n185 VSUBS 0.005852f
C729 B.n186 VSUBS 0.005852f
C730 B.n187 VSUBS 0.005852f
C731 B.n188 VSUBS 0.005852f
C732 B.n189 VSUBS 0.005852f
C733 B.n190 VSUBS 0.005852f
C734 B.n191 VSUBS 0.005852f
C735 B.n192 VSUBS 0.005852f
C736 B.n193 VSUBS 0.005852f
C737 B.n194 VSUBS 0.005852f
C738 B.n195 VSUBS 0.005852f
C739 B.n196 VSUBS 0.005852f
C740 B.n197 VSUBS 0.005852f
C741 B.n198 VSUBS 0.005852f
C742 B.n199 VSUBS 0.005852f
C743 B.n200 VSUBS 0.01266f
C744 B.n201 VSUBS 0.013159f
C745 B.n202 VSUBS 0.013159f
C746 B.n203 VSUBS 0.005852f
C747 B.n204 VSUBS 0.005852f
C748 B.n205 VSUBS 0.005852f
C749 B.n206 VSUBS 0.005852f
C750 B.n207 VSUBS 0.005852f
C751 B.n208 VSUBS 0.005852f
C752 B.n209 VSUBS 0.005852f
C753 B.n210 VSUBS 0.005852f
C754 B.n211 VSUBS 0.005852f
C755 B.n212 VSUBS 0.005852f
C756 B.n213 VSUBS 0.005852f
C757 B.n214 VSUBS 0.005852f
C758 B.n215 VSUBS 0.005852f
C759 B.n216 VSUBS 0.005852f
C760 B.n217 VSUBS 0.005852f
C761 B.n218 VSUBS 0.005852f
C762 B.n219 VSUBS 0.005852f
C763 B.n220 VSUBS 0.005852f
C764 B.n221 VSUBS 0.005852f
C765 B.n222 VSUBS 0.005852f
C766 B.n223 VSUBS 0.005852f
C767 B.n224 VSUBS 0.005852f
C768 B.n225 VSUBS 0.005852f
C769 B.n226 VSUBS 0.005852f
C770 B.n227 VSUBS 0.005852f
C771 B.n228 VSUBS 0.005852f
C772 B.n229 VSUBS 0.005852f
C773 B.n230 VSUBS 0.005852f
C774 B.n231 VSUBS 0.005852f
C775 B.n232 VSUBS 0.005852f
C776 B.n233 VSUBS 0.005852f
C777 B.n234 VSUBS 0.005852f
C778 B.n235 VSUBS 0.005852f
C779 B.n236 VSUBS 0.005852f
C780 B.n237 VSUBS 0.005852f
C781 B.n238 VSUBS 0.005852f
C782 B.n239 VSUBS 0.005852f
C783 B.n240 VSUBS 0.005852f
C784 B.n241 VSUBS 0.005852f
C785 B.n242 VSUBS 0.005852f
C786 B.n243 VSUBS 0.005852f
C787 B.n244 VSUBS 0.005852f
C788 B.n245 VSUBS 0.005852f
C789 B.n246 VSUBS 0.005852f
C790 B.n247 VSUBS 0.005852f
C791 B.n248 VSUBS 0.005852f
C792 B.n249 VSUBS 0.005852f
C793 B.n250 VSUBS 0.005852f
C794 B.n251 VSUBS 0.005852f
C795 B.n252 VSUBS 0.005852f
C796 B.n253 VSUBS 0.005852f
C797 B.n254 VSUBS 0.005852f
C798 B.n255 VSUBS 0.005852f
C799 B.n256 VSUBS 0.005852f
C800 B.n257 VSUBS 0.005852f
C801 B.n258 VSUBS 0.005852f
C802 B.n259 VSUBS 0.005852f
C803 B.n260 VSUBS 0.004045f
C804 B.n261 VSUBS 0.013559f
C805 B.n262 VSUBS 0.004733f
C806 B.n263 VSUBS 0.005852f
C807 B.n264 VSUBS 0.005852f
C808 B.n265 VSUBS 0.005852f
C809 B.n266 VSUBS 0.005852f
C810 B.n267 VSUBS 0.005852f
C811 B.n268 VSUBS 0.005852f
C812 B.n269 VSUBS 0.005852f
C813 B.n270 VSUBS 0.005852f
C814 B.n271 VSUBS 0.005852f
C815 B.n272 VSUBS 0.005852f
C816 B.n273 VSUBS 0.005852f
C817 B.t2 VSUBS 0.164156f
C818 B.t1 VSUBS 0.197203f
C819 B.t0 VSUBS 1.51687f
C820 B.n274 VSUBS 0.315846f
C821 B.n275 VSUBS 0.205763f
C822 B.n276 VSUBS 0.013559f
C823 B.n277 VSUBS 0.004733f
C824 B.n278 VSUBS 0.005852f
C825 B.n279 VSUBS 0.005852f
C826 B.n280 VSUBS 0.005852f
C827 B.n281 VSUBS 0.005852f
C828 B.n282 VSUBS 0.005852f
C829 B.n283 VSUBS 0.005852f
C830 B.n284 VSUBS 0.005852f
C831 B.n285 VSUBS 0.005852f
C832 B.n286 VSUBS 0.005852f
C833 B.n287 VSUBS 0.005852f
C834 B.n288 VSUBS 0.005852f
C835 B.n289 VSUBS 0.005852f
C836 B.n290 VSUBS 0.005852f
C837 B.n291 VSUBS 0.005852f
C838 B.n292 VSUBS 0.005852f
C839 B.n293 VSUBS 0.005852f
C840 B.n294 VSUBS 0.005852f
C841 B.n295 VSUBS 0.005852f
C842 B.n296 VSUBS 0.005852f
C843 B.n297 VSUBS 0.005852f
C844 B.n298 VSUBS 0.005852f
C845 B.n299 VSUBS 0.005852f
C846 B.n300 VSUBS 0.005852f
C847 B.n301 VSUBS 0.005852f
C848 B.n302 VSUBS 0.005852f
C849 B.n303 VSUBS 0.005852f
C850 B.n304 VSUBS 0.005852f
C851 B.n305 VSUBS 0.005852f
C852 B.n306 VSUBS 0.005852f
C853 B.n307 VSUBS 0.005852f
C854 B.n308 VSUBS 0.005852f
C855 B.n309 VSUBS 0.005852f
C856 B.n310 VSUBS 0.005852f
C857 B.n311 VSUBS 0.005852f
C858 B.n312 VSUBS 0.005852f
C859 B.n313 VSUBS 0.005852f
C860 B.n314 VSUBS 0.005852f
C861 B.n315 VSUBS 0.005852f
C862 B.n316 VSUBS 0.005852f
C863 B.n317 VSUBS 0.005852f
C864 B.n318 VSUBS 0.005852f
C865 B.n319 VSUBS 0.005852f
C866 B.n320 VSUBS 0.005852f
C867 B.n321 VSUBS 0.005852f
C868 B.n322 VSUBS 0.005852f
C869 B.n323 VSUBS 0.005852f
C870 B.n324 VSUBS 0.005852f
C871 B.n325 VSUBS 0.005852f
C872 B.n326 VSUBS 0.005852f
C873 B.n327 VSUBS 0.005852f
C874 B.n328 VSUBS 0.005852f
C875 B.n329 VSUBS 0.005852f
C876 B.n330 VSUBS 0.005852f
C877 B.n331 VSUBS 0.005852f
C878 B.n332 VSUBS 0.005852f
C879 B.n333 VSUBS 0.005852f
C880 B.n334 VSUBS 0.005852f
C881 B.n335 VSUBS 0.005852f
C882 B.n336 VSUBS 0.005852f
C883 B.n337 VSUBS 0.012401f
C884 B.n338 VSUBS 0.013159f
C885 B.n339 VSUBS 0.01266f
C886 B.n340 VSUBS 0.005852f
C887 B.n341 VSUBS 0.005852f
C888 B.n342 VSUBS 0.005852f
C889 B.n343 VSUBS 0.005852f
C890 B.n344 VSUBS 0.005852f
C891 B.n345 VSUBS 0.005852f
C892 B.n346 VSUBS 0.005852f
C893 B.n347 VSUBS 0.005852f
C894 B.n348 VSUBS 0.005852f
C895 B.n349 VSUBS 0.005852f
C896 B.n350 VSUBS 0.005852f
C897 B.n351 VSUBS 0.005852f
C898 B.n352 VSUBS 0.005852f
C899 B.n353 VSUBS 0.005852f
C900 B.n354 VSUBS 0.005852f
C901 B.n355 VSUBS 0.005852f
C902 B.n356 VSUBS 0.005852f
C903 B.n357 VSUBS 0.005852f
C904 B.n358 VSUBS 0.005852f
C905 B.n359 VSUBS 0.005852f
C906 B.n360 VSUBS 0.005852f
C907 B.n361 VSUBS 0.005852f
C908 B.n362 VSUBS 0.005852f
C909 B.n363 VSUBS 0.005852f
C910 B.n364 VSUBS 0.005852f
C911 B.n365 VSUBS 0.005852f
C912 B.n366 VSUBS 0.005852f
C913 B.n367 VSUBS 0.005852f
C914 B.n368 VSUBS 0.005852f
C915 B.n369 VSUBS 0.005852f
C916 B.n370 VSUBS 0.005852f
C917 B.n371 VSUBS 0.005852f
C918 B.n372 VSUBS 0.005852f
C919 B.n373 VSUBS 0.005852f
C920 B.n374 VSUBS 0.005852f
C921 B.n375 VSUBS 0.005852f
C922 B.n376 VSUBS 0.005852f
C923 B.n377 VSUBS 0.005852f
C924 B.n378 VSUBS 0.005852f
C925 B.n379 VSUBS 0.005852f
C926 B.n380 VSUBS 0.005852f
C927 B.n381 VSUBS 0.005852f
C928 B.n382 VSUBS 0.005852f
C929 B.n383 VSUBS 0.005852f
C930 B.n384 VSUBS 0.005852f
C931 B.n385 VSUBS 0.005852f
C932 B.n386 VSUBS 0.005852f
C933 B.n387 VSUBS 0.005852f
C934 B.n388 VSUBS 0.005852f
C935 B.n389 VSUBS 0.005852f
C936 B.n390 VSUBS 0.005852f
C937 B.n391 VSUBS 0.005852f
C938 B.n392 VSUBS 0.005852f
C939 B.n393 VSUBS 0.005852f
C940 B.n394 VSUBS 0.005852f
C941 B.n395 VSUBS 0.005852f
C942 B.n396 VSUBS 0.005852f
C943 B.n397 VSUBS 0.005852f
C944 B.n398 VSUBS 0.005852f
C945 B.n399 VSUBS 0.005852f
C946 B.n400 VSUBS 0.005852f
C947 B.n401 VSUBS 0.005852f
C948 B.n402 VSUBS 0.005852f
C949 B.n403 VSUBS 0.005852f
C950 B.n404 VSUBS 0.005852f
C951 B.n405 VSUBS 0.005852f
C952 B.n406 VSUBS 0.005852f
C953 B.n407 VSUBS 0.005852f
C954 B.n408 VSUBS 0.005852f
C955 B.n409 VSUBS 0.005852f
C956 B.n410 VSUBS 0.005852f
C957 B.n411 VSUBS 0.005852f
C958 B.n412 VSUBS 0.005852f
C959 B.n413 VSUBS 0.005852f
C960 B.n414 VSUBS 0.005852f
C961 B.n415 VSUBS 0.005852f
C962 B.n416 VSUBS 0.005852f
C963 B.n417 VSUBS 0.005852f
C964 B.n418 VSUBS 0.005852f
C965 B.n419 VSUBS 0.005852f
C966 B.n420 VSUBS 0.005852f
C967 B.n421 VSUBS 0.005852f
C968 B.n422 VSUBS 0.005852f
C969 B.n423 VSUBS 0.005852f
C970 B.n424 VSUBS 0.005852f
C971 B.n425 VSUBS 0.005852f
C972 B.n426 VSUBS 0.005852f
C973 B.n427 VSUBS 0.005852f
C974 B.n428 VSUBS 0.005852f
C975 B.n429 VSUBS 0.005852f
C976 B.n430 VSUBS 0.01266f
C977 B.n431 VSUBS 0.01266f
C978 B.n432 VSUBS 0.013159f
C979 B.n433 VSUBS 0.005852f
C980 B.n434 VSUBS 0.005852f
C981 B.n435 VSUBS 0.005852f
C982 B.n436 VSUBS 0.005852f
C983 B.n437 VSUBS 0.005852f
C984 B.n438 VSUBS 0.005852f
C985 B.n439 VSUBS 0.005852f
C986 B.n440 VSUBS 0.005852f
C987 B.n441 VSUBS 0.005852f
C988 B.n442 VSUBS 0.005852f
C989 B.n443 VSUBS 0.005852f
C990 B.n444 VSUBS 0.005852f
C991 B.n445 VSUBS 0.005852f
C992 B.n446 VSUBS 0.005852f
C993 B.n447 VSUBS 0.005852f
C994 B.n448 VSUBS 0.005852f
C995 B.n449 VSUBS 0.005852f
C996 B.n450 VSUBS 0.005852f
C997 B.n451 VSUBS 0.005852f
C998 B.n452 VSUBS 0.005852f
C999 B.n453 VSUBS 0.005852f
C1000 B.n454 VSUBS 0.005852f
C1001 B.n455 VSUBS 0.005852f
C1002 B.n456 VSUBS 0.005852f
C1003 B.n457 VSUBS 0.005852f
C1004 B.n458 VSUBS 0.005852f
C1005 B.n459 VSUBS 0.005852f
C1006 B.n460 VSUBS 0.005852f
C1007 B.n461 VSUBS 0.005852f
C1008 B.n462 VSUBS 0.005852f
C1009 B.n463 VSUBS 0.005852f
C1010 B.n464 VSUBS 0.005852f
C1011 B.n465 VSUBS 0.005852f
C1012 B.n466 VSUBS 0.005852f
C1013 B.n467 VSUBS 0.005852f
C1014 B.n468 VSUBS 0.005852f
C1015 B.n469 VSUBS 0.005852f
C1016 B.n470 VSUBS 0.005852f
C1017 B.n471 VSUBS 0.005852f
C1018 B.n472 VSUBS 0.005852f
C1019 B.n473 VSUBS 0.005852f
C1020 B.n474 VSUBS 0.005852f
C1021 B.n475 VSUBS 0.005852f
C1022 B.n476 VSUBS 0.005852f
C1023 B.n477 VSUBS 0.005852f
C1024 B.n478 VSUBS 0.005852f
C1025 B.n479 VSUBS 0.005852f
C1026 B.n480 VSUBS 0.005852f
C1027 B.n481 VSUBS 0.005852f
C1028 B.n482 VSUBS 0.005852f
C1029 B.n483 VSUBS 0.005852f
C1030 B.n484 VSUBS 0.005852f
C1031 B.n485 VSUBS 0.005852f
C1032 B.n486 VSUBS 0.005852f
C1033 B.n487 VSUBS 0.005852f
C1034 B.n488 VSUBS 0.005852f
C1035 B.n489 VSUBS 0.005852f
C1036 B.n490 VSUBS 0.005852f
C1037 B.n491 VSUBS 0.004045f
C1038 B.n492 VSUBS 0.013559f
C1039 B.n493 VSUBS 0.004733f
C1040 B.n494 VSUBS 0.005852f
C1041 B.n495 VSUBS 0.005852f
C1042 B.n496 VSUBS 0.005852f
C1043 B.n497 VSUBS 0.005852f
C1044 B.n498 VSUBS 0.005852f
C1045 B.n499 VSUBS 0.005852f
C1046 B.n500 VSUBS 0.005852f
C1047 B.n501 VSUBS 0.005852f
C1048 B.n502 VSUBS 0.005852f
C1049 B.n503 VSUBS 0.005852f
C1050 B.n504 VSUBS 0.005852f
C1051 B.n505 VSUBS 0.004733f
C1052 B.n506 VSUBS 0.013559f
C1053 B.n507 VSUBS 0.004045f
C1054 B.n508 VSUBS 0.005852f
C1055 B.n509 VSUBS 0.005852f
C1056 B.n510 VSUBS 0.005852f
C1057 B.n511 VSUBS 0.005852f
C1058 B.n512 VSUBS 0.005852f
C1059 B.n513 VSUBS 0.005852f
C1060 B.n514 VSUBS 0.005852f
C1061 B.n515 VSUBS 0.005852f
C1062 B.n516 VSUBS 0.005852f
C1063 B.n517 VSUBS 0.005852f
C1064 B.n518 VSUBS 0.005852f
C1065 B.n519 VSUBS 0.005852f
C1066 B.n520 VSUBS 0.005852f
C1067 B.n521 VSUBS 0.005852f
C1068 B.n522 VSUBS 0.005852f
C1069 B.n523 VSUBS 0.005852f
C1070 B.n524 VSUBS 0.005852f
C1071 B.n525 VSUBS 0.005852f
C1072 B.n526 VSUBS 0.005852f
C1073 B.n527 VSUBS 0.005852f
C1074 B.n528 VSUBS 0.005852f
C1075 B.n529 VSUBS 0.005852f
C1076 B.n530 VSUBS 0.005852f
C1077 B.n531 VSUBS 0.005852f
C1078 B.n532 VSUBS 0.005852f
C1079 B.n533 VSUBS 0.005852f
C1080 B.n534 VSUBS 0.005852f
C1081 B.n535 VSUBS 0.005852f
C1082 B.n536 VSUBS 0.005852f
C1083 B.n537 VSUBS 0.005852f
C1084 B.n538 VSUBS 0.005852f
C1085 B.n539 VSUBS 0.005852f
C1086 B.n540 VSUBS 0.005852f
C1087 B.n541 VSUBS 0.005852f
C1088 B.n542 VSUBS 0.005852f
C1089 B.n543 VSUBS 0.005852f
C1090 B.n544 VSUBS 0.005852f
C1091 B.n545 VSUBS 0.005852f
C1092 B.n546 VSUBS 0.005852f
C1093 B.n547 VSUBS 0.005852f
C1094 B.n548 VSUBS 0.005852f
C1095 B.n549 VSUBS 0.005852f
C1096 B.n550 VSUBS 0.005852f
C1097 B.n551 VSUBS 0.005852f
C1098 B.n552 VSUBS 0.005852f
C1099 B.n553 VSUBS 0.005852f
C1100 B.n554 VSUBS 0.005852f
C1101 B.n555 VSUBS 0.005852f
C1102 B.n556 VSUBS 0.005852f
C1103 B.n557 VSUBS 0.005852f
C1104 B.n558 VSUBS 0.005852f
C1105 B.n559 VSUBS 0.005852f
C1106 B.n560 VSUBS 0.005852f
C1107 B.n561 VSUBS 0.005852f
C1108 B.n562 VSUBS 0.005852f
C1109 B.n563 VSUBS 0.005852f
C1110 B.n564 VSUBS 0.005852f
C1111 B.n565 VSUBS 0.005852f
C1112 B.n566 VSUBS 0.013159f
C1113 B.n567 VSUBS 0.01266f
C1114 B.n568 VSUBS 0.01266f
C1115 B.n569 VSUBS 0.005852f
C1116 B.n570 VSUBS 0.005852f
C1117 B.n571 VSUBS 0.005852f
C1118 B.n572 VSUBS 0.005852f
C1119 B.n573 VSUBS 0.005852f
C1120 B.n574 VSUBS 0.005852f
C1121 B.n575 VSUBS 0.005852f
C1122 B.n576 VSUBS 0.005852f
C1123 B.n577 VSUBS 0.005852f
C1124 B.n578 VSUBS 0.005852f
C1125 B.n579 VSUBS 0.005852f
C1126 B.n580 VSUBS 0.005852f
C1127 B.n581 VSUBS 0.005852f
C1128 B.n582 VSUBS 0.005852f
C1129 B.n583 VSUBS 0.005852f
C1130 B.n584 VSUBS 0.005852f
C1131 B.n585 VSUBS 0.005852f
C1132 B.n586 VSUBS 0.005852f
C1133 B.n587 VSUBS 0.005852f
C1134 B.n588 VSUBS 0.005852f
C1135 B.n589 VSUBS 0.005852f
C1136 B.n590 VSUBS 0.005852f
C1137 B.n591 VSUBS 0.005852f
C1138 B.n592 VSUBS 0.005852f
C1139 B.n593 VSUBS 0.005852f
C1140 B.n594 VSUBS 0.005852f
C1141 B.n595 VSUBS 0.005852f
C1142 B.n596 VSUBS 0.005852f
C1143 B.n597 VSUBS 0.005852f
C1144 B.n598 VSUBS 0.005852f
C1145 B.n599 VSUBS 0.005852f
C1146 B.n600 VSUBS 0.005852f
C1147 B.n601 VSUBS 0.005852f
C1148 B.n602 VSUBS 0.005852f
C1149 B.n603 VSUBS 0.005852f
C1150 B.n604 VSUBS 0.005852f
C1151 B.n605 VSUBS 0.005852f
C1152 B.n606 VSUBS 0.005852f
C1153 B.n607 VSUBS 0.005852f
C1154 B.n608 VSUBS 0.005852f
C1155 B.n609 VSUBS 0.005852f
C1156 B.n610 VSUBS 0.005852f
C1157 B.n611 VSUBS 0.007637f
C1158 B.n612 VSUBS 0.008135f
C1159 B.n613 VSUBS 0.016177f
.ends

