* NGSPICE file created from diff_pair_sample_1098.ext - technology: sky130A

.subckt diff_pair_sample_1098 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t9 B.t2 sky130_fd_pr__nfet_01v8 ad=1.089 pd=6.93 as=2.574 ps=13.98 w=6.6 l=0.85
X1 VDD1.t4 VP.t1 VTAIL.t7 B.t5 sky130_fd_pr__nfet_01v8 ad=2.574 pd=13.98 as=1.089 ps=6.93 w=6.6 l=0.85
X2 B.t19 B.t17 B.t18 B.t11 sky130_fd_pr__nfet_01v8 ad=2.574 pd=13.98 as=0 ps=0 w=6.6 l=0.85
X3 B.t16 B.t14 B.t15 B.t7 sky130_fd_pr__nfet_01v8 ad=2.574 pd=13.98 as=0 ps=0 w=6.6 l=0.85
X4 VDD2.t5 VN.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.574 pd=13.98 as=1.089 ps=6.93 w=6.6 l=0.85
X5 VDD2.t4 VN.t1 VTAIL.t11 B.t5 sky130_fd_pr__nfet_01v8 ad=2.574 pd=13.98 as=1.089 ps=6.93 w=6.6 l=0.85
X6 VTAIL.t4 VN.t2 VDD2.t3 B.t4 sky130_fd_pr__nfet_01v8 ad=1.089 pd=6.93 as=1.089 ps=6.93 w=6.6 l=0.85
X7 VDD1.t3 VP.t2 VTAIL.t10 B.t3 sky130_fd_pr__nfet_01v8 ad=1.089 pd=6.93 as=2.574 ps=13.98 w=6.6 l=0.85
X8 VTAIL.t5 VP.t3 VDD1.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=1.089 pd=6.93 as=1.089 ps=6.93 w=6.6 l=0.85
X9 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=2.574 pd=13.98 as=0 ps=0 w=6.6 l=0.85
X10 VTAIL.t1 VN.t3 VDD2.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=1.089 pd=6.93 as=1.089 ps=6.93 w=6.6 l=0.85
X11 VDD2.t1 VN.t4 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.089 pd=6.93 as=2.574 ps=13.98 w=6.6 l=0.85
X12 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=2.574 pd=13.98 as=0 ps=0 w=6.6 l=0.85
X13 VDD2.t0 VN.t5 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.089 pd=6.93 as=2.574 ps=13.98 w=6.6 l=0.85
X14 VTAIL.t8 VP.t4 VDD1.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=1.089 pd=6.93 as=1.089 ps=6.93 w=6.6 l=0.85
X15 VDD1.t0 VP.t5 VTAIL.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=2.574 pd=13.98 as=1.089 ps=6.93 w=6.6 l=0.85
R0 VP.n5 VP.t5 248.974
R1 VP.n12 VP.t1 233.345
R2 VP.n19 VP.t2 233.345
R3 VP.n9 VP.t0 233.345
R4 VP.n1 VP.t4 187.13
R5 VP.n4 VP.t3 187.13
R6 VP.n20 VP.n19 161.3
R7 VP.n7 VP.n6 161.3
R8 VP.n8 VP.n3 161.3
R9 VP.n10 VP.n9 161.3
R10 VP.n18 VP.n0 161.3
R11 VP.n17 VP.n16 161.3
R12 VP.n15 VP.n14 161.3
R13 VP.n13 VP.n2 161.3
R14 VP.n12 VP.n11 161.3
R15 VP.n14 VP.n13 56.0773
R16 VP.n18 VP.n17 56.0773
R17 VP.n8 VP.n7 56.0773
R18 VP.n6 VP.n5 43.8087
R19 VP.n5 VP.n4 42.8016
R20 VP.n11 VP.n10 37.6596
R21 VP.n14 VP.n1 12.2964
R22 VP.n17 VP.n1 12.2964
R23 VP.n7 VP.n4 12.2964
R24 VP.n13 VP.n12 0.730803
R25 VP.n19 VP.n18 0.730803
R26 VP.n9 VP.n8 0.730803
R27 VP.n6 VP.n3 0.189894
R28 VP.n10 VP.n3 0.189894
R29 VP.n11 VP.n2 0.189894
R30 VP.n15 VP.n2 0.189894
R31 VP.n16 VP.n15 0.189894
R32 VP.n16 VP.n0 0.189894
R33 VP.n20 VP.n0 0.189894
R34 VP VP.n20 0.0516364
R35 VTAIL.n146 VTAIL.n116 289.615
R36 VTAIL.n32 VTAIL.n2 289.615
R37 VTAIL.n110 VTAIL.n80 289.615
R38 VTAIL.n72 VTAIL.n42 289.615
R39 VTAIL.n129 VTAIL.n128 185
R40 VTAIL.n131 VTAIL.n130 185
R41 VTAIL.n124 VTAIL.n123 185
R42 VTAIL.n137 VTAIL.n136 185
R43 VTAIL.n139 VTAIL.n138 185
R44 VTAIL.n120 VTAIL.n119 185
R45 VTAIL.n145 VTAIL.n144 185
R46 VTAIL.n147 VTAIL.n146 185
R47 VTAIL.n15 VTAIL.n14 185
R48 VTAIL.n17 VTAIL.n16 185
R49 VTAIL.n10 VTAIL.n9 185
R50 VTAIL.n23 VTAIL.n22 185
R51 VTAIL.n25 VTAIL.n24 185
R52 VTAIL.n6 VTAIL.n5 185
R53 VTAIL.n31 VTAIL.n30 185
R54 VTAIL.n33 VTAIL.n32 185
R55 VTAIL.n111 VTAIL.n110 185
R56 VTAIL.n109 VTAIL.n108 185
R57 VTAIL.n84 VTAIL.n83 185
R58 VTAIL.n103 VTAIL.n102 185
R59 VTAIL.n101 VTAIL.n100 185
R60 VTAIL.n88 VTAIL.n87 185
R61 VTAIL.n95 VTAIL.n94 185
R62 VTAIL.n93 VTAIL.n92 185
R63 VTAIL.n73 VTAIL.n72 185
R64 VTAIL.n71 VTAIL.n70 185
R65 VTAIL.n46 VTAIL.n45 185
R66 VTAIL.n65 VTAIL.n64 185
R67 VTAIL.n63 VTAIL.n62 185
R68 VTAIL.n50 VTAIL.n49 185
R69 VTAIL.n57 VTAIL.n56 185
R70 VTAIL.n55 VTAIL.n54 185
R71 VTAIL.n127 VTAIL.t2 147.659
R72 VTAIL.n13 VTAIL.t10 147.659
R73 VTAIL.n91 VTAIL.t9 147.659
R74 VTAIL.n53 VTAIL.t3 147.659
R75 VTAIL.n130 VTAIL.n129 104.615
R76 VTAIL.n130 VTAIL.n123 104.615
R77 VTAIL.n137 VTAIL.n123 104.615
R78 VTAIL.n138 VTAIL.n137 104.615
R79 VTAIL.n138 VTAIL.n119 104.615
R80 VTAIL.n145 VTAIL.n119 104.615
R81 VTAIL.n146 VTAIL.n145 104.615
R82 VTAIL.n16 VTAIL.n15 104.615
R83 VTAIL.n16 VTAIL.n9 104.615
R84 VTAIL.n23 VTAIL.n9 104.615
R85 VTAIL.n24 VTAIL.n23 104.615
R86 VTAIL.n24 VTAIL.n5 104.615
R87 VTAIL.n31 VTAIL.n5 104.615
R88 VTAIL.n32 VTAIL.n31 104.615
R89 VTAIL.n110 VTAIL.n109 104.615
R90 VTAIL.n109 VTAIL.n83 104.615
R91 VTAIL.n102 VTAIL.n83 104.615
R92 VTAIL.n102 VTAIL.n101 104.615
R93 VTAIL.n101 VTAIL.n87 104.615
R94 VTAIL.n94 VTAIL.n87 104.615
R95 VTAIL.n94 VTAIL.n93 104.615
R96 VTAIL.n72 VTAIL.n71 104.615
R97 VTAIL.n71 VTAIL.n45 104.615
R98 VTAIL.n64 VTAIL.n45 104.615
R99 VTAIL.n64 VTAIL.n63 104.615
R100 VTAIL.n63 VTAIL.n49 104.615
R101 VTAIL.n56 VTAIL.n49 104.615
R102 VTAIL.n56 VTAIL.n55 104.615
R103 VTAIL.n129 VTAIL.t2 52.3082
R104 VTAIL.n15 VTAIL.t10 52.3082
R105 VTAIL.n93 VTAIL.t9 52.3082
R106 VTAIL.n55 VTAIL.t3 52.3082
R107 VTAIL.n79 VTAIL.n78 47.0681
R108 VTAIL.n41 VTAIL.n40 47.0681
R109 VTAIL.n1 VTAIL.n0 47.0679
R110 VTAIL.n39 VTAIL.n38 47.0679
R111 VTAIL.n151 VTAIL.n150 29.8581
R112 VTAIL.n37 VTAIL.n36 29.8581
R113 VTAIL.n115 VTAIL.n114 29.8581
R114 VTAIL.n77 VTAIL.n76 29.8581
R115 VTAIL.n41 VTAIL.n39 20.091
R116 VTAIL.n151 VTAIL.n115 19.0738
R117 VTAIL.n128 VTAIL.n127 15.6676
R118 VTAIL.n14 VTAIL.n13 15.6676
R119 VTAIL.n92 VTAIL.n91 15.6676
R120 VTAIL.n54 VTAIL.n53 15.6676
R121 VTAIL.n131 VTAIL.n126 12.8005
R122 VTAIL.n17 VTAIL.n12 12.8005
R123 VTAIL.n95 VTAIL.n90 12.8005
R124 VTAIL.n57 VTAIL.n52 12.8005
R125 VTAIL.n132 VTAIL.n124 12.0247
R126 VTAIL.n18 VTAIL.n10 12.0247
R127 VTAIL.n96 VTAIL.n88 12.0247
R128 VTAIL.n58 VTAIL.n50 12.0247
R129 VTAIL.n136 VTAIL.n135 11.249
R130 VTAIL.n22 VTAIL.n21 11.249
R131 VTAIL.n100 VTAIL.n99 11.249
R132 VTAIL.n62 VTAIL.n61 11.249
R133 VTAIL.n139 VTAIL.n122 10.4732
R134 VTAIL.n25 VTAIL.n8 10.4732
R135 VTAIL.n103 VTAIL.n86 10.4732
R136 VTAIL.n65 VTAIL.n48 10.4732
R137 VTAIL.n140 VTAIL.n120 9.69747
R138 VTAIL.n26 VTAIL.n6 9.69747
R139 VTAIL.n104 VTAIL.n84 9.69747
R140 VTAIL.n66 VTAIL.n46 9.69747
R141 VTAIL.n150 VTAIL.n149 9.45567
R142 VTAIL.n36 VTAIL.n35 9.45567
R143 VTAIL.n114 VTAIL.n113 9.45567
R144 VTAIL.n76 VTAIL.n75 9.45567
R145 VTAIL.n118 VTAIL.n117 9.3005
R146 VTAIL.n143 VTAIL.n142 9.3005
R147 VTAIL.n141 VTAIL.n140 9.3005
R148 VTAIL.n122 VTAIL.n121 9.3005
R149 VTAIL.n135 VTAIL.n134 9.3005
R150 VTAIL.n133 VTAIL.n132 9.3005
R151 VTAIL.n126 VTAIL.n125 9.3005
R152 VTAIL.n149 VTAIL.n148 9.3005
R153 VTAIL.n4 VTAIL.n3 9.3005
R154 VTAIL.n29 VTAIL.n28 9.3005
R155 VTAIL.n27 VTAIL.n26 9.3005
R156 VTAIL.n8 VTAIL.n7 9.3005
R157 VTAIL.n21 VTAIL.n20 9.3005
R158 VTAIL.n19 VTAIL.n18 9.3005
R159 VTAIL.n12 VTAIL.n11 9.3005
R160 VTAIL.n35 VTAIL.n34 9.3005
R161 VTAIL.n113 VTAIL.n112 9.3005
R162 VTAIL.n82 VTAIL.n81 9.3005
R163 VTAIL.n107 VTAIL.n106 9.3005
R164 VTAIL.n105 VTAIL.n104 9.3005
R165 VTAIL.n86 VTAIL.n85 9.3005
R166 VTAIL.n99 VTAIL.n98 9.3005
R167 VTAIL.n97 VTAIL.n96 9.3005
R168 VTAIL.n90 VTAIL.n89 9.3005
R169 VTAIL.n75 VTAIL.n74 9.3005
R170 VTAIL.n44 VTAIL.n43 9.3005
R171 VTAIL.n69 VTAIL.n68 9.3005
R172 VTAIL.n67 VTAIL.n66 9.3005
R173 VTAIL.n48 VTAIL.n47 9.3005
R174 VTAIL.n61 VTAIL.n60 9.3005
R175 VTAIL.n59 VTAIL.n58 9.3005
R176 VTAIL.n52 VTAIL.n51 9.3005
R177 VTAIL.n144 VTAIL.n143 8.92171
R178 VTAIL.n30 VTAIL.n29 8.92171
R179 VTAIL.n108 VTAIL.n107 8.92171
R180 VTAIL.n70 VTAIL.n69 8.92171
R181 VTAIL.n147 VTAIL.n118 8.14595
R182 VTAIL.n33 VTAIL.n4 8.14595
R183 VTAIL.n111 VTAIL.n82 8.14595
R184 VTAIL.n73 VTAIL.n44 8.14595
R185 VTAIL.n148 VTAIL.n116 7.3702
R186 VTAIL.n34 VTAIL.n2 7.3702
R187 VTAIL.n112 VTAIL.n80 7.3702
R188 VTAIL.n74 VTAIL.n42 7.3702
R189 VTAIL.n150 VTAIL.n116 6.59444
R190 VTAIL.n36 VTAIL.n2 6.59444
R191 VTAIL.n114 VTAIL.n80 6.59444
R192 VTAIL.n76 VTAIL.n42 6.59444
R193 VTAIL.n148 VTAIL.n147 5.81868
R194 VTAIL.n34 VTAIL.n33 5.81868
R195 VTAIL.n112 VTAIL.n111 5.81868
R196 VTAIL.n74 VTAIL.n73 5.81868
R197 VTAIL.n144 VTAIL.n118 5.04292
R198 VTAIL.n30 VTAIL.n4 5.04292
R199 VTAIL.n108 VTAIL.n82 5.04292
R200 VTAIL.n70 VTAIL.n44 5.04292
R201 VTAIL.n127 VTAIL.n125 4.38571
R202 VTAIL.n13 VTAIL.n11 4.38571
R203 VTAIL.n91 VTAIL.n89 4.38571
R204 VTAIL.n53 VTAIL.n51 4.38571
R205 VTAIL.n143 VTAIL.n120 4.26717
R206 VTAIL.n29 VTAIL.n6 4.26717
R207 VTAIL.n107 VTAIL.n84 4.26717
R208 VTAIL.n69 VTAIL.n46 4.26717
R209 VTAIL.n140 VTAIL.n139 3.49141
R210 VTAIL.n26 VTAIL.n25 3.49141
R211 VTAIL.n104 VTAIL.n103 3.49141
R212 VTAIL.n66 VTAIL.n65 3.49141
R213 VTAIL.n0 VTAIL.t0 3.0005
R214 VTAIL.n0 VTAIL.t1 3.0005
R215 VTAIL.n38 VTAIL.t7 3.0005
R216 VTAIL.n38 VTAIL.t8 3.0005
R217 VTAIL.n78 VTAIL.t6 3.0005
R218 VTAIL.n78 VTAIL.t5 3.0005
R219 VTAIL.n40 VTAIL.t11 3.0005
R220 VTAIL.n40 VTAIL.t4 3.0005
R221 VTAIL.n136 VTAIL.n122 2.71565
R222 VTAIL.n22 VTAIL.n8 2.71565
R223 VTAIL.n100 VTAIL.n86 2.71565
R224 VTAIL.n62 VTAIL.n48 2.71565
R225 VTAIL.n135 VTAIL.n124 1.93989
R226 VTAIL.n21 VTAIL.n10 1.93989
R227 VTAIL.n99 VTAIL.n88 1.93989
R228 VTAIL.n61 VTAIL.n50 1.93989
R229 VTAIL.n132 VTAIL.n131 1.16414
R230 VTAIL.n18 VTAIL.n17 1.16414
R231 VTAIL.n96 VTAIL.n95 1.16414
R232 VTAIL.n58 VTAIL.n57 1.16414
R233 VTAIL.n77 VTAIL.n41 1.01774
R234 VTAIL.n115 VTAIL.n79 1.01774
R235 VTAIL.n39 VTAIL.n37 1.01774
R236 VTAIL.n79 VTAIL.n77 0.978948
R237 VTAIL.n37 VTAIL.n1 0.978948
R238 VTAIL VTAIL.n151 0.705241
R239 VTAIL.n128 VTAIL.n126 0.388379
R240 VTAIL.n14 VTAIL.n12 0.388379
R241 VTAIL.n92 VTAIL.n90 0.388379
R242 VTAIL.n54 VTAIL.n52 0.388379
R243 VTAIL VTAIL.n1 0.313
R244 VTAIL.n133 VTAIL.n125 0.155672
R245 VTAIL.n134 VTAIL.n133 0.155672
R246 VTAIL.n134 VTAIL.n121 0.155672
R247 VTAIL.n141 VTAIL.n121 0.155672
R248 VTAIL.n142 VTAIL.n141 0.155672
R249 VTAIL.n142 VTAIL.n117 0.155672
R250 VTAIL.n149 VTAIL.n117 0.155672
R251 VTAIL.n19 VTAIL.n11 0.155672
R252 VTAIL.n20 VTAIL.n19 0.155672
R253 VTAIL.n20 VTAIL.n7 0.155672
R254 VTAIL.n27 VTAIL.n7 0.155672
R255 VTAIL.n28 VTAIL.n27 0.155672
R256 VTAIL.n28 VTAIL.n3 0.155672
R257 VTAIL.n35 VTAIL.n3 0.155672
R258 VTAIL.n113 VTAIL.n81 0.155672
R259 VTAIL.n106 VTAIL.n81 0.155672
R260 VTAIL.n106 VTAIL.n105 0.155672
R261 VTAIL.n105 VTAIL.n85 0.155672
R262 VTAIL.n98 VTAIL.n85 0.155672
R263 VTAIL.n98 VTAIL.n97 0.155672
R264 VTAIL.n97 VTAIL.n89 0.155672
R265 VTAIL.n75 VTAIL.n43 0.155672
R266 VTAIL.n68 VTAIL.n43 0.155672
R267 VTAIL.n68 VTAIL.n67 0.155672
R268 VTAIL.n67 VTAIL.n47 0.155672
R269 VTAIL.n60 VTAIL.n47 0.155672
R270 VTAIL.n60 VTAIL.n59 0.155672
R271 VTAIL.n59 VTAIL.n51 0.155672
R272 VDD1.n30 VDD1.n0 289.615
R273 VDD1.n65 VDD1.n35 289.615
R274 VDD1.n31 VDD1.n30 185
R275 VDD1.n29 VDD1.n28 185
R276 VDD1.n4 VDD1.n3 185
R277 VDD1.n23 VDD1.n22 185
R278 VDD1.n21 VDD1.n20 185
R279 VDD1.n8 VDD1.n7 185
R280 VDD1.n15 VDD1.n14 185
R281 VDD1.n13 VDD1.n12 185
R282 VDD1.n48 VDD1.n47 185
R283 VDD1.n50 VDD1.n49 185
R284 VDD1.n43 VDD1.n42 185
R285 VDD1.n56 VDD1.n55 185
R286 VDD1.n58 VDD1.n57 185
R287 VDD1.n39 VDD1.n38 185
R288 VDD1.n64 VDD1.n63 185
R289 VDD1.n66 VDD1.n65 185
R290 VDD1.n11 VDD1.t0 147.659
R291 VDD1.n46 VDD1.t4 147.659
R292 VDD1.n30 VDD1.n29 104.615
R293 VDD1.n29 VDD1.n3 104.615
R294 VDD1.n22 VDD1.n3 104.615
R295 VDD1.n22 VDD1.n21 104.615
R296 VDD1.n21 VDD1.n7 104.615
R297 VDD1.n14 VDD1.n7 104.615
R298 VDD1.n14 VDD1.n13 104.615
R299 VDD1.n49 VDD1.n48 104.615
R300 VDD1.n49 VDD1.n42 104.615
R301 VDD1.n56 VDD1.n42 104.615
R302 VDD1.n57 VDD1.n56 104.615
R303 VDD1.n57 VDD1.n38 104.615
R304 VDD1.n64 VDD1.n38 104.615
R305 VDD1.n65 VDD1.n64 104.615
R306 VDD1.n71 VDD1.n70 63.9457
R307 VDD1.n73 VDD1.n72 63.7467
R308 VDD1.n13 VDD1.t0 52.3082
R309 VDD1.n48 VDD1.t4 52.3082
R310 VDD1 VDD1.n34 47.358
R311 VDD1.n71 VDD1.n69 47.2444
R312 VDD1.n73 VDD1.n71 33.8026
R313 VDD1.n12 VDD1.n11 15.6676
R314 VDD1.n47 VDD1.n46 15.6676
R315 VDD1.n15 VDD1.n10 12.8005
R316 VDD1.n50 VDD1.n45 12.8005
R317 VDD1.n16 VDD1.n8 12.0247
R318 VDD1.n51 VDD1.n43 12.0247
R319 VDD1.n20 VDD1.n19 11.249
R320 VDD1.n55 VDD1.n54 11.249
R321 VDD1.n23 VDD1.n6 10.4732
R322 VDD1.n58 VDD1.n41 10.4732
R323 VDD1.n24 VDD1.n4 9.69747
R324 VDD1.n59 VDD1.n39 9.69747
R325 VDD1.n34 VDD1.n33 9.45567
R326 VDD1.n69 VDD1.n68 9.45567
R327 VDD1.n33 VDD1.n32 9.3005
R328 VDD1.n2 VDD1.n1 9.3005
R329 VDD1.n27 VDD1.n26 9.3005
R330 VDD1.n25 VDD1.n24 9.3005
R331 VDD1.n6 VDD1.n5 9.3005
R332 VDD1.n19 VDD1.n18 9.3005
R333 VDD1.n17 VDD1.n16 9.3005
R334 VDD1.n10 VDD1.n9 9.3005
R335 VDD1.n37 VDD1.n36 9.3005
R336 VDD1.n62 VDD1.n61 9.3005
R337 VDD1.n60 VDD1.n59 9.3005
R338 VDD1.n41 VDD1.n40 9.3005
R339 VDD1.n54 VDD1.n53 9.3005
R340 VDD1.n52 VDD1.n51 9.3005
R341 VDD1.n45 VDD1.n44 9.3005
R342 VDD1.n68 VDD1.n67 9.3005
R343 VDD1.n28 VDD1.n27 8.92171
R344 VDD1.n63 VDD1.n62 8.92171
R345 VDD1.n31 VDD1.n2 8.14595
R346 VDD1.n66 VDD1.n37 8.14595
R347 VDD1.n32 VDD1.n0 7.3702
R348 VDD1.n67 VDD1.n35 7.3702
R349 VDD1.n34 VDD1.n0 6.59444
R350 VDD1.n69 VDD1.n35 6.59444
R351 VDD1.n32 VDD1.n31 5.81868
R352 VDD1.n67 VDD1.n66 5.81868
R353 VDD1.n28 VDD1.n2 5.04292
R354 VDD1.n63 VDD1.n37 5.04292
R355 VDD1.n11 VDD1.n9 4.38571
R356 VDD1.n46 VDD1.n44 4.38571
R357 VDD1.n27 VDD1.n4 4.26717
R358 VDD1.n62 VDD1.n39 4.26717
R359 VDD1.n24 VDD1.n23 3.49141
R360 VDD1.n59 VDD1.n58 3.49141
R361 VDD1.n72 VDD1.t2 3.0005
R362 VDD1.n72 VDD1.t5 3.0005
R363 VDD1.n70 VDD1.t1 3.0005
R364 VDD1.n70 VDD1.t3 3.0005
R365 VDD1.n20 VDD1.n6 2.71565
R366 VDD1.n55 VDD1.n41 2.71565
R367 VDD1.n19 VDD1.n8 1.93989
R368 VDD1.n54 VDD1.n43 1.93989
R369 VDD1.n16 VDD1.n15 1.16414
R370 VDD1.n51 VDD1.n50 1.16414
R371 VDD1.n12 VDD1.n10 0.388379
R372 VDD1.n47 VDD1.n45 0.388379
R373 VDD1 VDD1.n73 0.196621
R374 VDD1.n33 VDD1.n1 0.155672
R375 VDD1.n26 VDD1.n1 0.155672
R376 VDD1.n26 VDD1.n25 0.155672
R377 VDD1.n25 VDD1.n5 0.155672
R378 VDD1.n18 VDD1.n5 0.155672
R379 VDD1.n18 VDD1.n17 0.155672
R380 VDD1.n17 VDD1.n9 0.155672
R381 VDD1.n52 VDD1.n44 0.155672
R382 VDD1.n53 VDD1.n52 0.155672
R383 VDD1.n53 VDD1.n40 0.155672
R384 VDD1.n60 VDD1.n40 0.155672
R385 VDD1.n61 VDD1.n60 0.155672
R386 VDD1.n61 VDD1.n36 0.155672
R387 VDD1.n68 VDD1.n36 0.155672
R388 B.n374 B.n373 585
R389 B.n374 B.n43 585
R390 B.n377 B.n376 585
R391 B.n378 B.n78 585
R392 B.n380 B.n379 585
R393 B.n382 B.n77 585
R394 B.n385 B.n384 585
R395 B.n386 B.n76 585
R396 B.n388 B.n387 585
R397 B.n390 B.n75 585
R398 B.n393 B.n392 585
R399 B.n394 B.n74 585
R400 B.n396 B.n395 585
R401 B.n398 B.n73 585
R402 B.n401 B.n400 585
R403 B.n402 B.n72 585
R404 B.n404 B.n403 585
R405 B.n406 B.n71 585
R406 B.n409 B.n408 585
R407 B.n410 B.n70 585
R408 B.n412 B.n411 585
R409 B.n414 B.n69 585
R410 B.n417 B.n416 585
R411 B.n418 B.n68 585
R412 B.n420 B.n419 585
R413 B.n422 B.n67 585
R414 B.n425 B.n424 585
R415 B.n427 B.n64 585
R416 B.n429 B.n428 585
R417 B.n431 B.n63 585
R418 B.n434 B.n433 585
R419 B.n435 B.n62 585
R420 B.n437 B.n436 585
R421 B.n439 B.n61 585
R422 B.n441 B.n440 585
R423 B.n443 B.n442 585
R424 B.n446 B.n445 585
R425 B.n447 B.n56 585
R426 B.n449 B.n448 585
R427 B.n451 B.n55 585
R428 B.n454 B.n453 585
R429 B.n455 B.n54 585
R430 B.n457 B.n456 585
R431 B.n459 B.n53 585
R432 B.n462 B.n461 585
R433 B.n463 B.n52 585
R434 B.n465 B.n464 585
R435 B.n467 B.n51 585
R436 B.n470 B.n469 585
R437 B.n471 B.n50 585
R438 B.n473 B.n472 585
R439 B.n475 B.n49 585
R440 B.n478 B.n477 585
R441 B.n479 B.n48 585
R442 B.n481 B.n480 585
R443 B.n483 B.n47 585
R444 B.n486 B.n485 585
R445 B.n487 B.n46 585
R446 B.n489 B.n488 585
R447 B.n491 B.n45 585
R448 B.n494 B.n493 585
R449 B.n495 B.n44 585
R450 B.n372 B.n42 585
R451 B.n498 B.n42 585
R452 B.n371 B.n41 585
R453 B.n499 B.n41 585
R454 B.n370 B.n40 585
R455 B.n500 B.n40 585
R456 B.n369 B.n368 585
R457 B.n368 B.n36 585
R458 B.n367 B.n35 585
R459 B.n506 B.n35 585
R460 B.n366 B.n34 585
R461 B.n507 B.n34 585
R462 B.n365 B.n33 585
R463 B.n508 B.n33 585
R464 B.n364 B.n363 585
R465 B.n363 B.n29 585
R466 B.n362 B.n28 585
R467 B.n514 B.n28 585
R468 B.n361 B.n27 585
R469 B.n515 B.n27 585
R470 B.n360 B.n26 585
R471 B.n516 B.n26 585
R472 B.n359 B.n358 585
R473 B.n358 B.n25 585
R474 B.n357 B.n21 585
R475 B.n522 B.n21 585
R476 B.n356 B.n20 585
R477 B.n523 B.n20 585
R478 B.n355 B.n19 585
R479 B.n524 B.n19 585
R480 B.n354 B.n353 585
R481 B.n353 B.n18 585
R482 B.n352 B.n14 585
R483 B.n530 B.n14 585
R484 B.n351 B.n13 585
R485 B.n531 B.n13 585
R486 B.n350 B.n12 585
R487 B.n532 B.n12 585
R488 B.n349 B.n348 585
R489 B.n348 B.n8 585
R490 B.n347 B.n7 585
R491 B.n538 B.n7 585
R492 B.n346 B.n6 585
R493 B.n539 B.n6 585
R494 B.n345 B.n5 585
R495 B.n540 B.n5 585
R496 B.n344 B.n343 585
R497 B.n343 B.n4 585
R498 B.n342 B.n79 585
R499 B.n342 B.n341 585
R500 B.n332 B.n80 585
R501 B.n81 B.n80 585
R502 B.n334 B.n333 585
R503 B.n335 B.n334 585
R504 B.n331 B.n86 585
R505 B.n86 B.n85 585
R506 B.n330 B.n329 585
R507 B.n329 B.n328 585
R508 B.n88 B.n87 585
R509 B.n321 B.n88 585
R510 B.n320 B.n319 585
R511 B.n322 B.n320 585
R512 B.n318 B.n93 585
R513 B.n93 B.n92 585
R514 B.n317 B.n316 585
R515 B.n316 B.n315 585
R516 B.n95 B.n94 585
R517 B.n308 B.n95 585
R518 B.n307 B.n306 585
R519 B.n309 B.n307 585
R520 B.n305 B.n100 585
R521 B.n100 B.n99 585
R522 B.n304 B.n303 585
R523 B.n303 B.n302 585
R524 B.n102 B.n101 585
R525 B.n103 B.n102 585
R526 B.n295 B.n294 585
R527 B.n296 B.n295 585
R528 B.n293 B.n107 585
R529 B.n111 B.n107 585
R530 B.n292 B.n291 585
R531 B.n291 B.n290 585
R532 B.n109 B.n108 585
R533 B.n110 B.n109 585
R534 B.n283 B.n282 585
R535 B.n284 B.n283 585
R536 B.n281 B.n116 585
R537 B.n116 B.n115 585
R538 B.n280 B.n279 585
R539 B.n279 B.n278 585
R540 B.n275 B.n120 585
R541 B.n274 B.n273 585
R542 B.n271 B.n121 585
R543 B.n271 B.n119 585
R544 B.n270 B.n269 585
R545 B.n268 B.n267 585
R546 B.n266 B.n123 585
R547 B.n264 B.n263 585
R548 B.n262 B.n124 585
R549 B.n261 B.n260 585
R550 B.n258 B.n125 585
R551 B.n256 B.n255 585
R552 B.n254 B.n126 585
R553 B.n253 B.n252 585
R554 B.n250 B.n127 585
R555 B.n248 B.n247 585
R556 B.n246 B.n128 585
R557 B.n245 B.n244 585
R558 B.n242 B.n129 585
R559 B.n240 B.n239 585
R560 B.n238 B.n130 585
R561 B.n237 B.n236 585
R562 B.n234 B.n131 585
R563 B.n232 B.n231 585
R564 B.n230 B.n132 585
R565 B.n229 B.n228 585
R566 B.n226 B.n133 585
R567 B.n224 B.n223 585
R568 B.n222 B.n134 585
R569 B.n221 B.n220 585
R570 B.n218 B.n138 585
R571 B.n216 B.n215 585
R572 B.n214 B.n139 585
R573 B.n213 B.n212 585
R574 B.n210 B.n140 585
R575 B.n208 B.n207 585
R576 B.n205 B.n141 585
R577 B.n204 B.n203 585
R578 B.n201 B.n144 585
R579 B.n199 B.n198 585
R580 B.n197 B.n145 585
R581 B.n196 B.n195 585
R582 B.n193 B.n146 585
R583 B.n191 B.n190 585
R584 B.n189 B.n147 585
R585 B.n188 B.n187 585
R586 B.n185 B.n148 585
R587 B.n183 B.n182 585
R588 B.n181 B.n149 585
R589 B.n180 B.n179 585
R590 B.n177 B.n150 585
R591 B.n175 B.n174 585
R592 B.n173 B.n151 585
R593 B.n172 B.n171 585
R594 B.n169 B.n152 585
R595 B.n167 B.n166 585
R596 B.n165 B.n153 585
R597 B.n164 B.n163 585
R598 B.n161 B.n154 585
R599 B.n159 B.n158 585
R600 B.n157 B.n156 585
R601 B.n118 B.n117 585
R602 B.n277 B.n276 585
R603 B.n278 B.n277 585
R604 B.n114 B.n113 585
R605 B.n115 B.n114 585
R606 B.n286 B.n285 585
R607 B.n285 B.n284 585
R608 B.n287 B.n112 585
R609 B.n112 B.n110 585
R610 B.n289 B.n288 585
R611 B.n290 B.n289 585
R612 B.n106 B.n105 585
R613 B.n111 B.n106 585
R614 B.n298 B.n297 585
R615 B.n297 B.n296 585
R616 B.n299 B.n104 585
R617 B.n104 B.n103 585
R618 B.n301 B.n300 585
R619 B.n302 B.n301 585
R620 B.n98 B.n97 585
R621 B.n99 B.n98 585
R622 B.n311 B.n310 585
R623 B.n310 B.n309 585
R624 B.n312 B.n96 585
R625 B.n308 B.n96 585
R626 B.n314 B.n313 585
R627 B.n315 B.n314 585
R628 B.n91 B.n90 585
R629 B.n92 B.n91 585
R630 B.n324 B.n323 585
R631 B.n323 B.n322 585
R632 B.n325 B.n89 585
R633 B.n321 B.n89 585
R634 B.n327 B.n326 585
R635 B.n328 B.n327 585
R636 B.n84 B.n83 585
R637 B.n85 B.n84 585
R638 B.n337 B.n336 585
R639 B.n336 B.n335 585
R640 B.n338 B.n82 585
R641 B.n82 B.n81 585
R642 B.n340 B.n339 585
R643 B.n341 B.n340 585
R644 B.n2 B.n0 585
R645 B.n4 B.n2 585
R646 B.n3 B.n1 585
R647 B.n539 B.n3 585
R648 B.n537 B.n536 585
R649 B.n538 B.n537 585
R650 B.n535 B.n9 585
R651 B.n9 B.n8 585
R652 B.n534 B.n533 585
R653 B.n533 B.n532 585
R654 B.n11 B.n10 585
R655 B.n531 B.n11 585
R656 B.n529 B.n528 585
R657 B.n530 B.n529 585
R658 B.n527 B.n15 585
R659 B.n18 B.n15 585
R660 B.n526 B.n525 585
R661 B.n525 B.n524 585
R662 B.n17 B.n16 585
R663 B.n523 B.n17 585
R664 B.n521 B.n520 585
R665 B.n522 B.n521 585
R666 B.n519 B.n22 585
R667 B.n25 B.n22 585
R668 B.n518 B.n517 585
R669 B.n517 B.n516 585
R670 B.n24 B.n23 585
R671 B.n515 B.n24 585
R672 B.n513 B.n512 585
R673 B.n514 B.n513 585
R674 B.n511 B.n30 585
R675 B.n30 B.n29 585
R676 B.n510 B.n509 585
R677 B.n509 B.n508 585
R678 B.n32 B.n31 585
R679 B.n507 B.n32 585
R680 B.n505 B.n504 585
R681 B.n506 B.n505 585
R682 B.n503 B.n37 585
R683 B.n37 B.n36 585
R684 B.n502 B.n501 585
R685 B.n501 B.n500 585
R686 B.n39 B.n38 585
R687 B.n499 B.n39 585
R688 B.n497 B.n496 585
R689 B.n498 B.n497 585
R690 B.n542 B.n541 585
R691 B.n541 B.n540 585
R692 B.n277 B.n120 502.111
R693 B.n497 B.n44 502.111
R694 B.n279 B.n118 502.111
R695 B.n374 B.n42 502.111
R696 B.n142 B.t14 388.918
R697 B.n135 B.t6 388.918
R698 B.n57 B.t10 388.918
R699 B.n65 B.t17 388.918
R700 B.n375 B.n43 256.663
R701 B.n381 B.n43 256.663
R702 B.n383 B.n43 256.663
R703 B.n389 B.n43 256.663
R704 B.n391 B.n43 256.663
R705 B.n397 B.n43 256.663
R706 B.n399 B.n43 256.663
R707 B.n405 B.n43 256.663
R708 B.n407 B.n43 256.663
R709 B.n413 B.n43 256.663
R710 B.n415 B.n43 256.663
R711 B.n421 B.n43 256.663
R712 B.n423 B.n43 256.663
R713 B.n430 B.n43 256.663
R714 B.n432 B.n43 256.663
R715 B.n438 B.n43 256.663
R716 B.n60 B.n43 256.663
R717 B.n444 B.n43 256.663
R718 B.n450 B.n43 256.663
R719 B.n452 B.n43 256.663
R720 B.n458 B.n43 256.663
R721 B.n460 B.n43 256.663
R722 B.n466 B.n43 256.663
R723 B.n468 B.n43 256.663
R724 B.n474 B.n43 256.663
R725 B.n476 B.n43 256.663
R726 B.n482 B.n43 256.663
R727 B.n484 B.n43 256.663
R728 B.n490 B.n43 256.663
R729 B.n492 B.n43 256.663
R730 B.n272 B.n119 256.663
R731 B.n122 B.n119 256.663
R732 B.n265 B.n119 256.663
R733 B.n259 B.n119 256.663
R734 B.n257 B.n119 256.663
R735 B.n251 B.n119 256.663
R736 B.n249 B.n119 256.663
R737 B.n243 B.n119 256.663
R738 B.n241 B.n119 256.663
R739 B.n235 B.n119 256.663
R740 B.n233 B.n119 256.663
R741 B.n227 B.n119 256.663
R742 B.n225 B.n119 256.663
R743 B.n219 B.n119 256.663
R744 B.n217 B.n119 256.663
R745 B.n211 B.n119 256.663
R746 B.n209 B.n119 256.663
R747 B.n202 B.n119 256.663
R748 B.n200 B.n119 256.663
R749 B.n194 B.n119 256.663
R750 B.n192 B.n119 256.663
R751 B.n186 B.n119 256.663
R752 B.n184 B.n119 256.663
R753 B.n178 B.n119 256.663
R754 B.n176 B.n119 256.663
R755 B.n170 B.n119 256.663
R756 B.n168 B.n119 256.663
R757 B.n162 B.n119 256.663
R758 B.n160 B.n119 256.663
R759 B.n155 B.n119 256.663
R760 B.n142 B.t16 211.999
R761 B.n65 B.t18 211.999
R762 B.n135 B.t9 211.999
R763 B.n57 B.t12 211.999
R764 B.n143 B.t15 189.113
R765 B.n66 B.t19 189.113
R766 B.n136 B.t8 189.113
R767 B.n58 B.t13 189.113
R768 B.n277 B.n114 163.367
R769 B.n285 B.n114 163.367
R770 B.n285 B.n112 163.367
R771 B.n289 B.n112 163.367
R772 B.n289 B.n106 163.367
R773 B.n297 B.n106 163.367
R774 B.n297 B.n104 163.367
R775 B.n301 B.n104 163.367
R776 B.n301 B.n98 163.367
R777 B.n310 B.n98 163.367
R778 B.n310 B.n96 163.367
R779 B.n314 B.n96 163.367
R780 B.n314 B.n91 163.367
R781 B.n323 B.n91 163.367
R782 B.n323 B.n89 163.367
R783 B.n327 B.n89 163.367
R784 B.n327 B.n84 163.367
R785 B.n336 B.n84 163.367
R786 B.n336 B.n82 163.367
R787 B.n340 B.n82 163.367
R788 B.n340 B.n2 163.367
R789 B.n541 B.n2 163.367
R790 B.n541 B.n3 163.367
R791 B.n537 B.n3 163.367
R792 B.n537 B.n9 163.367
R793 B.n533 B.n9 163.367
R794 B.n533 B.n11 163.367
R795 B.n529 B.n11 163.367
R796 B.n529 B.n15 163.367
R797 B.n525 B.n15 163.367
R798 B.n525 B.n17 163.367
R799 B.n521 B.n17 163.367
R800 B.n521 B.n22 163.367
R801 B.n517 B.n22 163.367
R802 B.n517 B.n24 163.367
R803 B.n513 B.n24 163.367
R804 B.n513 B.n30 163.367
R805 B.n509 B.n30 163.367
R806 B.n509 B.n32 163.367
R807 B.n505 B.n32 163.367
R808 B.n505 B.n37 163.367
R809 B.n501 B.n37 163.367
R810 B.n501 B.n39 163.367
R811 B.n497 B.n39 163.367
R812 B.n273 B.n271 163.367
R813 B.n271 B.n270 163.367
R814 B.n267 B.n266 163.367
R815 B.n264 B.n124 163.367
R816 B.n260 B.n258 163.367
R817 B.n256 B.n126 163.367
R818 B.n252 B.n250 163.367
R819 B.n248 B.n128 163.367
R820 B.n244 B.n242 163.367
R821 B.n240 B.n130 163.367
R822 B.n236 B.n234 163.367
R823 B.n232 B.n132 163.367
R824 B.n228 B.n226 163.367
R825 B.n224 B.n134 163.367
R826 B.n220 B.n218 163.367
R827 B.n216 B.n139 163.367
R828 B.n212 B.n210 163.367
R829 B.n208 B.n141 163.367
R830 B.n203 B.n201 163.367
R831 B.n199 B.n145 163.367
R832 B.n195 B.n193 163.367
R833 B.n191 B.n147 163.367
R834 B.n187 B.n185 163.367
R835 B.n183 B.n149 163.367
R836 B.n179 B.n177 163.367
R837 B.n175 B.n151 163.367
R838 B.n171 B.n169 163.367
R839 B.n167 B.n153 163.367
R840 B.n163 B.n161 163.367
R841 B.n159 B.n156 163.367
R842 B.n279 B.n116 163.367
R843 B.n283 B.n116 163.367
R844 B.n283 B.n109 163.367
R845 B.n291 B.n109 163.367
R846 B.n291 B.n107 163.367
R847 B.n295 B.n107 163.367
R848 B.n295 B.n102 163.367
R849 B.n303 B.n102 163.367
R850 B.n303 B.n100 163.367
R851 B.n307 B.n100 163.367
R852 B.n307 B.n95 163.367
R853 B.n316 B.n95 163.367
R854 B.n316 B.n93 163.367
R855 B.n320 B.n93 163.367
R856 B.n320 B.n88 163.367
R857 B.n329 B.n88 163.367
R858 B.n329 B.n86 163.367
R859 B.n334 B.n86 163.367
R860 B.n334 B.n80 163.367
R861 B.n342 B.n80 163.367
R862 B.n343 B.n342 163.367
R863 B.n343 B.n5 163.367
R864 B.n6 B.n5 163.367
R865 B.n7 B.n6 163.367
R866 B.n348 B.n7 163.367
R867 B.n348 B.n12 163.367
R868 B.n13 B.n12 163.367
R869 B.n14 B.n13 163.367
R870 B.n353 B.n14 163.367
R871 B.n353 B.n19 163.367
R872 B.n20 B.n19 163.367
R873 B.n21 B.n20 163.367
R874 B.n358 B.n21 163.367
R875 B.n358 B.n26 163.367
R876 B.n27 B.n26 163.367
R877 B.n28 B.n27 163.367
R878 B.n363 B.n28 163.367
R879 B.n363 B.n33 163.367
R880 B.n34 B.n33 163.367
R881 B.n35 B.n34 163.367
R882 B.n368 B.n35 163.367
R883 B.n368 B.n40 163.367
R884 B.n41 B.n40 163.367
R885 B.n42 B.n41 163.367
R886 B.n493 B.n491 163.367
R887 B.n489 B.n46 163.367
R888 B.n485 B.n483 163.367
R889 B.n481 B.n48 163.367
R890 B.n477 B.n475 163.367
R891 B.n473 B.n50 163.367
R892 B.n469 B.n467 163.367
R893 B.n465 B.n52 163.367
R894 B.n461 B.n459 163.367
R895 B.n457 B.n54 163.367
R896 B.n453 B.n451 163.367
R897 B.n449 B.n56 163.367
R898 B.n445 B.n443 163.367
R899 B.n440 B.n439 163.367
R900 B.n437 B.n62 163.367
R901 B.n433 B.n431 163.367
R902 B.n429 B.n64 163.367
R903 B.n424 B.n422 163.367
R904 B.n420 B.n68 163.367
R905 B.n416 B.n414 163.367
R906 B.n412 B.n70 163.367
R907 B.n408 B.n406 163.367
R908 B.n404 B.n72 163.367
R909 B.n400 B.n398 163.367
R910 B.n396 B.n74 163.367
R911 B.n392 B.n390 163.367
R912 B.n388 B.n76 163.367
R913 B.n384 B.n382 163.367
R914 B.n380 B.n78 163.367
R915 B.n376 B.n374 163.367
R916 B.n278 B.n119 113.938
R917 B.n498 B.n43 113.938
R918 B.n272 B.n120 71.676
R919 B.n270 B.n122 71.676
R920 B.n266 B.n265 71.676
R921 B.n259 B.n124 71.676
R922 B.n258 B.n257 71.676
R923 B.n251 B.n126 71.676
R924 B.n250 B.n249 71.676
R925 B.n243 B.n128 71.676
R926 B.n242 B.n241 71.676
R927 B.n235 B.n130 71.676
R928 B.n234 B.n233 71.676
R929 B.n227 B.n132 71.676
R930 B.n226 B.n225 71.676
R931 B.n219 B.n134 71.676
R932 B.n218 B.n217 71.676
R933 B.n211 B.n139 71.676
R934 B.n210 B.n209 71.676
R935 B.n202 B.n141 71.676
R936 B.n201 B.n200 71.676
R937 B.n194 B.n145 71.676
R938 B.n193 B.n192 71.676
R939 B.n186 B.n147 71.676
R940 B.n185 B.n184 71.676
R941 B.n178 B.n149 71.676
R942 B.n177 B.n176 71.676
R943 B.n170 B.n151 71.676
R944 B.n169 B.n168 71.676
R945 B.n162 B.n153 71.676
R946 B.n161 B.n160 71.676
R947 B.n156 B.n155 71.676
R948 B.n492 B.n44 71.676
R949 B.n491 B.n490 71.676
R950 B.n484 B.n46 71.676
R951 B.n483 B.n482 71.676
R952 B.n476 B.n48 71.676
R953 B.n475 B.n474 71.676
R954 B.n468 B.n50 71.676
R955 B.n467 B.n466 71.676
R956 B.n460 B.n52 71.676
R957 B.n459 B.n458 71.676
R958 B.n452 B.n54 71.676
R959 B.n451 B.n450 71.676
R960 B.n444 B.n56 71.676
R961 B.n443 B.n60 71.676
R962 B.n439 B.n438 71.676
R963 B.n432 B.n62 71.676
R964 B.n431 B.n430 71.676
R965 B.n423 B.n64 71.676
R966 B.n422 B.n421 71.676
R967 B.n415 B.n68 71.676
R968 B.n414 B.n413 71.676
R969 B.n407 B.n70 71.676
R970 B.n406 B.n405 71.676
R971 B.n399 B.n72 71.676
R972 B.n398 B.n397 71.676
R973 B.n391 B.n74 71.676
R974 B.n390 B.n389 71.676
R975 B.n383 B.n76 71.676
R976 B.n382 B.n381 71.676
R977 B.n375 B.n78 71.676
R978 B.n376 B.n375 71.676
R979 B.n381 B.n380 71.676
R980 B.n384 B.n383 71.676
R981 B.n389 B.n388 71.676
R982 B.n392 B.n391 71.676
R983 B.n397 B.n396 71.676
R984 B.n400 B.n399 71.676
R985 B.n405 B.n404 71.676
R986 B.n408 B.n407 71.676
R987 B.n413 B.n412 71.676
R988 B.n416 B.n415 71.676
R989 B.n421 B.n420 71.676
R990 B.n424 B.n423 71.676
R991 B.n430 B.n429 71.676
R992 B.n433 B.n432 71.676
R993 B.n438 B.n437 71.676
R994 B.n440 B.n60 71.676
R995 B.n445 B.n444 71.676
R996 B.n450 B.n449 71.676
R997 B.n453 B.n452 71.676
R998 B.n458 B.n457 71.676
R999 B.n461 B.n460 71.676
R1000 B.n466 B.n465 71.676
R1001 B.n469 B.n468 71.676
R1002 B.n474 B.n473 71.676
R1003 B.n477 B.n476 71.676
R1004 B.n482 B.n481 71.676
R1005 B.n485 B.n484 71.676
R1006 B.n490 B.n489 71.676
R1007 B.n493 B.n492 71.676
R1008 B.n273 B.n272 71.676
R1009 B.n267 B.n122 71.676
R1010 B.n265 B.n264 71.676
R1011 B.n260 B.n259 71.676
R1012 B.n257 B.n256 71.676
R1013 B.n252 B.n251 71.676
R1014 B.n249 B.n248 71.676
R1015 B.n244 B.n243 71.676
R1016 B.n241 B.n240 71.676
R1017 B.n236 B.n235 71.676
R1018 B.n233 B.n232 71.676
R1019 B.n228 B.n227 71.676
R1020 B.n225 B.n224 71.676
R1021 B.n220 B.n219 71.676
R1022 B.n217 B.n216 71.676
R1023 B.n212 B.n211 71.676
R1024 B.n209 B.n208 71.676
R1025 B.n203 B.n202 71.676
R1026 B.n200 B.n199 71.676
R1027 B.n195 B.n194 71.676
R1028 B.n192 B.n191 71.676
R1029 B.n187 B.n186 71.676
R1030 B.n184 B.n183 71.676
R1031 B.n179 B.n178 71.676
R1032 B.n176 B.n175 71.676
R1033 B.n171 B.n170 71.676
R1034 B.n168 B.n167 71.676
R1035 B.n163 B.n162 71.676
R1036 B.n160 B.n159 71.676
R1037 B.n155 B.n118 71.676
R1038 B.n278 B.n115 62.99
R1039 B.n284 B.n115 62.99
R1040 B.n284 B.n110 62.99
R1041 B.n290 B.n110 62.99
R1042 B.n290 B.n111 62.99
R1043 B.n296 B.n103 62.99
R1044 B.n302 B.n103 62.99
R1045 B.n302 B.n99 62.99
R1046 B.n309 B.n99 62.99
R1047 B.n309 B.n308 62.99
R1048 B.n315 B.n92 62.99
R1049 B.n322 B.n92 62.99
R1050 B.n322 B.n321 62.99
R1051 B.n328 B.n85 62.99
R1052 B.n335 B.n85 62.99
R1053 B.n341 B.n81 62.99
R1054 B.n341 B.n4 62.99
R1055 B.n540 B.n4 62.99
R1056 B.n540 B.n539 62.99
R1057 B.n539 B.n538 62.99
R1058 B.n538 B.n8 62.99
R1059 B.n532 B.n531 62.99
R1060 B.n531 B.n530 62.99
R1061 B.n524 B.n18 62.99
R1062 B.n524 B.n523 62.99
R1063 B.n523 B.n522 62.99
R1064 B.n516 B.n25 62.99
R1065 B.n516 B.n515 62.99
R1066 B.n515 B.n514 62.99
R1067 B.n514 B.n29 62.99
R1068 B.n508 B.n29 62.99
R1069 B.n507 B.n506 62.99
R1070 B.n506 B.n36 62.99
R1071 B.n500 B.n36 62.99
R1072 B.n500 B.n499 62.99
R1073 B.n499 B.n498 62.99
R1074 B.n296 B.t7 60.211
R1075 B.n508 B.t11 60.211
R1076 B.n206 B.n143 59.5399
R1077 B.n137 B.n136 59.5399
R1078 B.n59 B.n58 59.5399
R1079 B.n426 B.n66 59.5399
R1080 B.n328 B.t4 50.9479
R1081 B.n530 B.t1 50.9479
R1082 B.n308 B.t5 45.39
R1083 B.n25 B.t2 45.39
R1084 B.n335 B.t3 41.6847
R1085 B.n532 B.t0 41.6847
R1086 B.n496 B.n495 32.6249
R1087 B.n373 B.n372 32.6249
R1088 B.n280 B.n117 32.6249
R1089 B.n276 B.n275 32.6249
R1090 B.n143 B.n142 22.8853
R1091 B.n136 B.n135 22.8853
R1092 B.n58 B.n57 22.8853
R1093 B.n66 B.n65 22.8853
R1094 B.t3 B.n81 21.3058
R1095 B.t0 B.n8 21.3058
R1096 B B.n542 18.0485
R1097 B.n315 B.t5 17.6005
R1098 B.n522 B.t2 17.6005
R1099 B.n321 B.t4 12.0426
R1100 B.n18 B.t1 12.0426
R1101 B.n495 B.n494 10.6151
R1102 B.n494 B.n45 10.6151
R1103 B.n488 B.n45 10.6151
R1104 B.n488 B.n487 10.6151
R1105 B.n487 B.n486 10.6151
R1106 B.n486 B.n47 10.6151
R1107 B.n480 B.n47 10.6151
R1108 B.n480 B.n479 10.6151
R1109 B.n479 B.n478 10.6151
R1110 B.n478 B.n49 10.6151
R1111 B.n472 B.n49 10.6151
R1112 B.n472 B.n471 10.6151
R1113 B.n471 B.n470 10.6151
R1114 B.n470 B.n51 10.6151
R1115 B.n464 B.n51 10.6151
R1116 B.n464 B.n463 10.6151
R1117 B.n463 B.n462 10.6151
R1118 B.n462 B.n53 10.6151
R1119 B.n456 B.n53 10.6151
R1120 B.n456 B.n455 10.6151
R1121 B.n455 B.n454 10.6151
R1122 B.n454 B.n55 10.6151
R1123 B.n448 B.n55 10.6151
R1124 B.n448 B.n447 10.6151
R1125 B.n447 B.n446 10.6151
R1126 B.n442 B.n441 10.6151
R1127 B.n441 B.n61 10.6151
R1128 B.n436 B.n61 10.6151
R1129 B.n436 B.n435 10.6151
R1130 B.n435 B.n434 10.6151
R1131 B.n434 B.n63 10.6151
R1132 B.n428 B.n63 10.6151
R1133 B.n428 B.n427 10.6151
R1134 B.n425 B.n67 10.6151
R1135 B.n419 B.n67 10.6151
R1136 B.n419 B.n418 10.6151
R1137 B.n418 B.n417 10.6151
R1138 B.n417 B.n69 10.6151
R1139 B.n411 B.n69 10.6151
R1140 B.n411 B.n410 10.6151
R1141 B.n410 B.n409 10.6151
R1142 B.n409 B.n71 10.6151
R1143 B.n403 B.n71 10.6151
R1144 B.n403 B.n402 10.6151
R1145 B.n402 B.n401 10.6151
R1146 B.n401 B.n73 10.6151
R1147 B.n395 B.n73 10.6151
R1148 B.n395 B.n394 10.6151
R1149 B.n394 B.n393 10.6151
R1150 B.n393 B.n75 10.6151
R1151 B.n387 B.n75 10.6151
R1152 B.n387 B.n386 10.6151
R1153 B.n386 B.n385 10.6151
R1154 B.n385 B.n77 10.6151
R1155 B.n379 B.n77 10.6151
R1156 B.n379 B.n378 10.6151
R1157 B.n378 B.n377 10.6151
R1158 B.n377 B.n373 10.6151
R1159 B.n281 B.n280 10.6151
R1160 B.n282 B.n281 10.6151
R1161 B.n282 B.n108 10.6151
R1162 B.n292 B.n108 10.6151
R1163 B.n293 B.n292 10.6151
R1164 B.n294 B.n293 10.6151
R1165 B.n294 B.n101 10.6151
R1166 B.n304 B.n101 10.6151
R1167 B.n305 B.n304 10.6151
R1168 B.n306 B.n305 10.6151
R1169 B.n306 B.n94 10.6151
R1170 B.n317 B.n94 10.6151
R1171 B.n318 B.n317 10.6151
R1172 B.n319 B.n318 10.6151
R1173 B.n319 B.n87 10.6151
R1174 B.n330 B.n87 10.6151
R1175 B.n331 B.n330 10.6151
R1176 B.n333 B.n331 10.6151
R1177 B.n333 B.n332 10.6151
R1178 B.n332 B.n79 10.6151
R1179 B.n344 B.n79 10.6151
R1180 B.n345 B.n344 10.6151
R1181 B.n346 B.n345 10.6151
R1182 B.n347 B.n346 10.6151
R1183 B.n349 B.n347 10.6151
R1184 B.n350 B.n349 10.6151
R1185 B.n351 B.n350 10.6151
R1186 B.n352 B.n351 10.6151
R1187 B.n354 B.n352 10.6151
R1188 B.n355 B.n354 10.6151
R1189 B.n356 B.n355 10.6151
R1190 B.n357 B.n356 10.6151
R1191 B.n359 B.n357 10.6151
R1192 B.n360 B.n359 10.6151
R1193 B.n361 B.n360 10.6151
R1194 B.n362 B.n361 10.6151
R1195 B.n364 B.n362 10.6151
R1196 B.n365 B.n364 10.6151
R1197 B.n366 B.n365 10.6151
R1198 B.n367 B.n366 10.6151
R1199 B.n369 B.n367 10.6151
R1200 B.n370 B.n369 10.6151
R1201 B.n371 B.n370 10.6151
R1202 B.n372 B.n371 10.6151
R1203 B.n275 B.n274 10.6151
R1204 B.n274 B.n121 10.6151
R1205 B.n269 B.n121 10.6151
R1206 B.n269 B.n268 10.6151
R1207 B.n268 B.n123 10.6151
R1208 B.n263 B.n123 10.6151
R1209 B.n263 B.n262 10.6151
R1210 B.n262 B.n261 10.6151
R1211 B.n261 B.n125 10.6151
R1212 B.n255 B.n125 10.6151
R1213 B.n255 B.n254 10.6151
R1214 B.n254 B.n253 10.6151
R1215 B.n253 B.n127 10.6151
R1216 B.n247 B.n127 10.6151
R1217 B.n247 B.n246 10.6151
R1218 B.n246 B.n245 10.6151
R1219 B.n245 B.n129 10.6151
R1220 B.n239 B.n129 10.6151
R1221 B.n239 B.n238 10.6151
R1222 B.n238 B.n237 10.6151
R1223 B.n237 B.n131 10.6151
R1224 B.n231 B.n131 10.6151
R1225 B.n231 B.n230 10.6151
R1226 B.n230 B.n229 10.6151
R1227 B.n229 B.n133 10.6151
R1228 B.n223 B.n222 10.6151
R1229 B.n222 B.n221 10.6151
R1230 B.n221 B.n138 10.6151
R1231 B.n215 B.n138 10.6151
R1232 B.n215 B.n214 10.6151
R1233 B.n214 B.n213 10.6151
R1234 B.n213 B.n140 10.6151
R1235 B.n207 B.n140 10.6151
R1236 B.n205 B.n204 10.6151
R1237 B.n204 B.n144 10.6151
R1238 B.n198 B.n144 10.6151
R1239 B.n198 B.n197 10.6151
R1240 B.n197 B.n196 10.6151
R1241 B.n196 B.n146 10.6151
R1242 B.n190 B.n146 10.6151
R1243 B.n190 B.n189 10.6151
R1244 B.n189 B.n188 10.6151
R1245 B.n188 B.n148 10.6151
R1246 B.n182 B.n148 10.6151
R1247 B.n182 B.n181 10.6151
R1248 B.n181 B.n180 10.6151
R1249 B.n180 B.n150 10.6151
R1250 B.n174 B.n150 10.6151
R1251 B.n174 B.n173 10.6151
R1252 B.n173 B.n172 10.6151
R1253 B.n172 B.n152 10.6151
R1254 B.n166 B.n152 10.6151
R1255 B.n166 B.n165 10.6151
R1256 B.n165 B.n164 10.6151
R1257 B.n164 B.n154 10.6151
R1258 B.n158 B.n154 10.6151
R1259 B.n158 B.n157 10.6151
R1260 B.n157 B.n117 10.6151
R1261 B.n276 B.n113 10.6151
R1262 B.n286 B.n113 10.6151
R1263 B.n287 B.n286 10.6151
R1264 B.n288 B.n287 10.6151
R1265 B.n288 B.n105 10.6151
R1266 B.n298 B.n105 10.6151
R1267 B.n299 B.n298 10.6151
R1268 B.n300 B.n299 10.6151
R1269 B.n300 B.n97 10.6151
R1270 B.n311 B.n97 10.6151
R1271 B.n312 B.n311 10.6151
R1272 B.n313 B.n312 10.6151
R1273 B.n313 B.n90 10.6151
R1274 B.n324 B.n90 10.6151
R1275 B.n325 B.n324 10.6151
R1276 B.n326 B.n325 10.6151
R1277 B.n326 B.n83 10.6151
R1278 B.n337 B.n83 10.6151
R1279 B.n338 B.n337 10.6151
R1280 B.n339 B.n338 10.6151
R1281 B.n339 B.n0 10.6151
R1282 B.n536 B.n1 10.6151
R1283 B.n536 B.n535 10.6151
R1284 B.n535 B.n534 10.6151
R1285 B.n534 B.n10 10.6151
R1286 B.n528 B.n10 10.6151
R1287 B.n528 B.n527 10.6151
R1288 B.n527 B.n526 10.6151
R1289 B.n526 B.n16 10.6151
R1290 B.n520 B.n16 10.6151
R1291 B.n520 B.n519 10.6151
R1292 B.n519 B.n518 10.6151
R1293 B.n518 B.n23 10.6151
R1294 B.n512 B.n23 10.6151
R1295 B.n512 B.n511 10.6151
R1296 B.n511 B.n510 10.6151
R1297 B.n510 B.n31 10.6151
R1298 B.n504 B.n31 10.6151
R1299 B.n504 B.n503 10.6151
R1300 B.n503 B.n502 10.6151
R1301 B.n502 B.n38 10.6151
R1302 B.n496 B.n38 10.6151
R1303 B.n442 B.n59 6.5566
R1304 B.n427 B.n426 6.5566
R1305 B.n223 B.n137 6.5566
R1306 B.n207 B.n206 6.5566
R1307 B.n446 B.n59 4.05904
R1308 B.n426 B.n425 4.05904
R1309 B.n137 B.n133 4.05904
R1310 B.n206 B.n205 4.05904
R1311 B.n542 B.n0 2.81026
R1312 B.n542 B.n1 2.81026
R1313 B.n111 B.t7 2.77945
R1314 B.t11 B.n507 2.77945
R1315 VN.n2 VN.t0 248.974
R1316 VN.n10 VN.t5 248.974
R1317 VN.n6 VN.t4 233.345
R1318 VN.n14 VN.t1 233.345
R1319 VN.n1 VN.t3 187.13
R1320 VN.n9 VN.t2 187.13
R1321 VN.n7 VN.n6 161.3
R1322 VN.n15 VN.n14 161.3
R1323 VN.n13 VN.n8 161.3
R1324 VN.n12 VN.n11 161.3
R1325 VN.n5 VN.n0 161.3
R1326 VN.n4 VN.n3 161.3
R1327 VN.n5 VN.n4 56.0773
R1328 VN.n13 VN.n12 56.0773
R1329 VN.n11 VN.n10 43.8087
R1330 VN.n3 VN.n2 43.8087
R1331 VN.n2 VN.n1 42.8016
R1332 VN.n10 VN.n9 42.8016
R1333 VN VN.n15 38.0403
R1334 VN.n4 VN.n1 12.2964
R1335 VN.n12 VN.n9 12.2964
R1336 VN.n6 VN.n5 0.730803
R1337 VN.n14 VN.n13 0.730803
R1338 VN.n15 VN.n8 0.189894
R1339 VN.n11 VN.n8 0.189894
R1340 VN.n3 VN.n0 0.189894
R1341 VN.n7 VN.n0 0.189894
R1342 VN VN.n7 0.0516364
R1343 VDD2.n67 VDD2.n37 289.615
R1344 VDD2.n30 VDD2.n0 289.615
R1345 VDD2.n68 VDD2.n67 185
R1346 VDD2.n66 VDD2.n65 185
R1347 VDD2.n41 VDD2.n40 185
R1348 VDD2.n60 VDD2.n59 185
R1349 VDD2.n58 VDD2.n57 185
R1350 VDD2.n45 VDD2.n44 185
R1351 VDD2.n52 VDD2.n51 185
R1352 VDD2.n50 VDD2.n49 185
R1353 VDD2.n13 VDD2.n12 185
R1354 VDD2.n15 VDD2.n14 185
R1355 VDD2.n8 VDD2.n7 185
R1356 VDD2.n21 VDD2.n20 185
R1357 VDD2.n23 VDD2.n22 185
R1358 VDD2.n4 VDD2.n3 185
R1359 VDD2.n29 VDD2.n28 185
R1360 VDD2.n31 VDD2.n30 185
R1361 VDD2.n48 VDD2.t4 147.659
R1362 VDD2.n11 VDD2.t5 147.659
R1363 VDD2.n67 VDD2.n66 104.615
R1364 VDD2.n66 VDD2.n40 104.615
R1365 VDD2.n59 VDD2.n40 104.615
R1366 VDD2.n59 VDD2.n58 104.615
R1367 VDD2.n58 VDD2.n44 104.615
R1368 VDD2.n51 VDD2.n44 104.615
R1369 VDD2.n51 VDD2.n50 104.615
R1370 VDD2.n14 VDD2.n13 104.615
R1371 VDD2.n14 VDD2.n7 104.615
R1372 VDD2.n21 VDD2.n7 104.615
R1373 VDD2.n22 VDD2.n21 104.615
R1374 VDD2.n22 VDD2.n3 104.615
R1375 VDD2.n29 VDD2.n3 104.615
R1376 VDD2.n30 VDD2.n29 104.615
R1377 VDD2.n36 VDD2.n35 63.9457
R1378 VDD2 VDD2.n73 63.9428
R1379 VDD2.n50 VDD2.t4 52.3082
R1380 VDD2.n13 VDD2.t5 52.3082
R1381 VDD2.n36 VDD2.n34 47.2444
R1382 VDD2.n72 VDD2.n71 46.5369
R1383 VDD2.n72 VDD2.n36 32.711
R1384 VDD2.n49 VDD2.n48 15.6676
R1385 VDD2.n12 VDD2.n11 15.6676
R1386 VDD2.n52 VDD2.n47 12.8005
R1387 VDD2.n15 VDD2.n10 12.8005
R1388 VDD2.n53 VDD2.n45 12.0247
R1389 VDD2.n16 VDD2.n8 12.0247
R1390 VDD2.n57 VDD2.n56 11.249
R1391 VDD2.n20 VDD2.n19 11.249
R1392 VDD2.n60 VDD2.n43 10.4732
R1393 VDD2.n23 VDD2.n6 10.4732
R1394 VDD2.n61 VDD2.n41 9.69747
R1395 VDD2.n24 VDD2.n4 9.69747
R1396 VDD2.n71 VDD2.n70 9.45567
R1397 VDD2.n34 VDD2.n33 9.45567
R1398 VDD2.n70 VDD2.n69 9.3005
R1399 VDD2.n39 VDD2.n38 9.3005
R1400 VDD2.n64 VDD2.n63 9.3005
R1401 VDD2.n62 VDD2.n61 9.3005
R1402 VDD2.n43 VDD2.n42 9.3005
R1403 VDD2.n56 VDD2.n55 9.3005
R1404 VDD2.n54 VDD2.n53 9.3005
R1405 VDD2.n47 VDD2.n46 9.3005
R1406 VDD2.n2 VDD2.n1 9.3005
R1407 VDD2.n27 VDD2.n26 9.3005
R1408 VDD2.n25 VDD2.n24 9.3005
R1409 VDD2.n6 VDD2.n5 9.3005
R1410 VDD2.n19 VDD2.n18 9.3005
R1411 VDD2.n17 VDD2.n16 9.3005
R1412 VDD2.n10 VDD2.n9 9.3005
R1413 VDD2.n33 VDD2.n32 9.3005
R1414 VDD2.n65 VDD2.n64 8.92171
R1415 VDD2.n28 VDD2.n27 8.92171
R1416 VDD2.n68 VDD2.n39 8.14595
R1417 VDD2.n31 VDD2.n2 8.14595
R1418 VDD2.n69 VDD2.n37 7.3702
R1419 VDD2.n32 VDD2.n0 7.3702
R1420 VDD2.n71 VDD2.n37 6.59444
R1421 VDD2.n34 VDD2.n0 6.59444
R1422 VDD2.n69 VDD2.n68 5.81868
R1423 VDD2.n32 VDD2.n31 5.81868
R1424 VDD2.n65 VDD2.n39 5.04292
R1425 VDD2.n28 VDD2.n2 5.04292
R1426 VDD2.n48 VDD2.n46 4.38571
R1427 VDD2.n11 VDD2.n9 4.38571
R1428 VDD2.n64 VDD2.n41 4.26717
R1429 VDD2.n27 VDD2.n4 4.26717
R1430 VDD2.n61 VDD2.n60 3.49141
R1431 VDD2.n24 VDD2.n23 3.49141
R1432 VDD2.n73 VDD2.t3 3.0005
R1433 VDD2.n73 VDD2.t0 3.0005
R1434 VDD2.n35 VDD2.t2 3.0005
R1435 VDD2.n35 VDD2.t1 3.0005
R1436 VDD2.n57 VDD2.n43 2.71565
R1437 VDD2.n20 VDD2.n6 2.71565
R1438 VDD2.n56 VDD2.n45 1.93989
R1439 VDD2.n19 VDD2.n8 1.93989
R1440 VDD2.n53 VDD2.n52 1.16414
R1441 VDD2.n16 VDD2.n15 1.16414
R1442 VDD2 VDD2.n72 0.821621
R1443 VDD2.n49 VDD2.n47 0.388379
R1444 VDD2.n12 VDD2.n10 0.388379
R1445 VDD2.n70 VDD2.n38 0.155672
R1446 VDD2.n63 VDD2.n38 0.155672
R1447 VDD2.n63 VDD2.n62 0.155672
R1448 VDD2.n62 VDD2.n42 0.155672
R1449 VDD2.n55 VDD2.n42 0.155672
R1450 VDD2.n55 VDD2.n54 0.155672
R1451 VDD2.n54 VDD2.n46 0.155672
R1452 VDD2.n17 VDD2.n9 0.155672
R1453 VDD2.n18 VDD2.n17 0.155672
R1454 VDD2.n18 VDD2.n5 0.155672
R1455 VDD2.n25 VDD2.n5 0.155672
R1456 VDD2.n26 VDD2.n25 0.155672
R1457 VDD2.n26 VDD2.n1 0.155672
R1458 VDD2.n33 VDD2.n1 0.155672
C0 VDD1 VP 2.92432f
C1 VTAIL VP 2.78436f
C2 VDD1 VN 0.148721f
C3 VTAIL VN 2.77001f
C4 VDD1 VDD2 0.764176f
C5 VTAIL VDD2 6.03347f
C6 VP VN 4.22573f
C7 VDD2 VP 0.309877f
C8 VDD2 VN 2.76573f
C9 VTAIL VDD1 5.99507f
C10 VDD2 B 3.640864f
C11 VDD1 B 3.66671f
C12 VTAIL B 4.379722f
C13 VN B 7.4177f
C14 VP B 5.774481f
C15 VDD2.n0 B 0.030933f
C16 VDD2.n1 B 0.022886f
C17 VDD2.n2 B 0.012298f
C18 VDD2.n3 B 0.029068f
C19 VDD2.n4 B 0.013021f
C20 VDD2.n5 B 0.022886f
C21 VDD2.n6 B 0.012298f
C22 VDD2.n7 B 0.029068f
C23 VDD2.n8 B 0.013021f
C24 VDD2.n9 B 0.607753f
C25 VDD2.n10 B 0.012298f
C26 VDD2.t5 B 0.047335f
C27 VDD2.n11 B 0.101201f
C28 VDD2.n12 B 0.017171f
C29 VDD2.n13 B 0.021801f
C30 VDD2.n14 B 0.029068f
C31 VDD2.n15 B 0.013021f
C32 VDD2.n16 B 0.012298f
C33 VDD2.n17 B 0.022886f
C34 VDD2.n18 B 0.022886f
C35 VDD2.n19 B 0.012298f
C36 VDD2.n20 B 0.013021f
C37 VDD2.n21 B 0.029068f
C38 VDD2.n22 B 0.029068f
C39 VDD2.n23 B 0.013021f
C40 VDD2.n24 B 0.012298f
C41 VDD2.n25 B 0.022886f
C42 VDD2.n26 B 0.022886f
C43 VDD2.n27 B 0.012298f
C44 VDD2.n28 B 0.013021f
C45 VDD2.n29 B 0.029068f
C46 VDD2.n30 B 0.060743f
C47 VDD2.n31 B 0.013021f
C48 VDD2.n32 B 0.012298f
C49 VDD2.n33 B 0.049148f
C50 VDD2.n34 B 0.0509f
C51 VDD2.t2 B 0.119363f
C52 VDD2.t1 B 0.119363f
C53 VDD2.n35 B 1.0063f
C54 VDD2.n36 B 1.45901f
C55 VDD2.n37 B 0.030933f
C56 VDD2.n38 B 0.022886f
C57 VDD2.n39 B 0.012298f
C58 VDD2.n40 B 0.029068f
C59 VDD2.n41 B 0.013021f
C60 VDD2.n42 B 0.022886f
C61 VDD2.n43 B 0.012298f
C62 VDD2.n44 B 0.029068f
C63 VDD2.n45 B 0.013021f
C64 VDD2.n46 B 0.607753f
C65 VDD2.n47 B 0.012298f
C66 VDD2.t4 B 0.047335f
C67 VDD2.n48 B 0.101201f
C68 VDD2.n49 B 0.017171f
C69 VDD2.n50 B 0.021801f
C70 VDD2.n51 B 0.029068f
C71 VDD2.n52 B 0.013021f
C72 VDD2.n53 B 0.012298f
C73 VDD2.n54 B 0.022886f
C74 VDD2.n55 B 0.022886f
C75 VDD2.n56 B 0.012298f
C76 VDD2.n57 B 0.013021f
C77 VDD2.n58 B 0.029068f
C78 VDD2.n59 B 0.029068f
C79 VDD2.n60 B 0.013021f
C80 VDD2.n61 B 0.012298f
C81 VDD2.n62 B 0.022886f
C82 VDD2.n63 B 0.022886f
C83 VDD2.n64 B 0.012298f
C84 VDD2.n65 B 0.013021f
C85 VDD2.n66 B 0.029068f
C86 VDD2.n67 B 0.060743f
C87 VDD2.n68 B 0.013021f
C88 VDD2.n69 B 0.012298f
C89 VDD2.n70 B 0.049148f
C90 VDD2.n71 B 0.049479f
C91 VDD2.n72 B 1.51446f
C92 VDD2.t3 B 0.119363f
C93 VDD2.t0 B 0.119363f
C94 VDD2.n73 B 1.00628f
C95 VN.n0 B 0.044037f
C96 VN.t3 B 0.657376f
C97 VN.n1 B 0.310154f
C98 VN.t0 B 0.734798f
C99 VN.n2 B 0.32164f
C100 VN.n3 B 0.180977f
C101 VN.n4 B 0.054715f
C102 VN.n5 B 0.013513f
C103 VN.t4 B 0.714372f
C104 VN.n6 B 0.312024f
C105 VN.n7 B 0.034127f
C106 VN.n8 B 0.044037f
C107 VN.t2 B 0.657376f
C108 VN.n9 B 0.310154f
C109 VN.t5 B 0.734798f
C110 VN.n10 B 0.32164f
C111 VN.n11 B 0.180977f
C112 VN.n12 B 0.054715f
C113 VN.n13 B 0.013513f
C114 VN.t1 B 0.714372f
C115 VN.n14 B 0.312024f
C116 VN.n15 B 1.53348f
C117 VDD1.n0 B 0.030987f
C118 VDD1.n1 B 0.022926f
C119 VDD1.n2 B 0.012319f
C120 VDD1.n3 B 0.029119f
C121 VDD1.n4 B 0.013044f
C122 VDD1.n5 B 0.022926f
C123 VDD1.n6 B 0.012319f
C124 VDD1.n7 B 0.029119f
C125 VDD1.n8 B 0.013044f
C126 VDD1.n9 B 0.608811f
C127 VDD1.n10 B 0.012319f
C128 VDD1.t0 B 0.047417f
C129 VDD1.n11 B 0.101377f
C130 VDD1.n12 B 0.017201f
C131 VDD1.n13 B 0.021839f
C132 VDD1.n14 B 0.029119f
C133 VDD1.n15 B 0.013044f
C134 VDD1.n16 B 0.012319f
C135 VDD1.n17 B 0.022926f
C136 VDD1.n18 B 0.022926f
C137 VDD1.n19 B 0.012319f
C138 VDD1.n20 B 0.013044f
C139 VDD1.n21 B 0.029119f
C140 VDD1.n22 B 0.029119f
C141 VDD1.n23 B 0.013044f
C142 VDD1.n24 B 0.012319f
C143 VDD1.n25 B 0.022926f
C144 VDD1.n26 B 0.022926f
C145 VDD1.n27 B 0.012319f
C146 VDD1.n28 B 0.013044f
C147 VDD1.n29 B 0.029119f
C148 VDD1.n30 B 0.060849f
C149 VDD1.n31 B 0.013044f
C150 VDD1.n32 B 0.012319f
C151 VDD1.n33 B 0.049234f
C152 VDD1.n34 B 0.051345f
C153 VDD1.n35 B 0.030987f
C154 VDD1.n36 B 0.022926f
C155 VDD1.n37 B 0.012319f
C156 VDD1.n38 B 0.029119f
C157 VDD1.n39 B 0.013044f
C158 VDD1.n40 B 0.022926f
C159 VDD1.n41 B 0.012319f
C160 VDD1.n42 B 0.029119f
C161 VDD1.n43 B 0.013044f
C162 VDD1.n44 B 0.608811f
C163 VDD1.n45 B 0.012319f
C164 VDD1.t4 B 0.047417f
C165 VDD1.n46 B 0.101377f
C166 VDD1.n47 B 0.017201f
C167 VDD1.n48 B 0.021839f
C168 VDD1.n49 B 0.029119f
C169 VDD1.n50 B 0.013044f
C170 VDD1.n51 B 0.012319f
C171 VDD1.n52 B 0.022926f
C172 VDD1.n53 B 0.022926f
C173 VDD1.n54 B 0.012319f
C174 VDD1.n55 B 0.013044f
C175 VDD1.n56 B 0.029119f
C176 VDD1.n57 B 0.029119f
C177 VDD1.n58 B 0.013044f
C178 VDD1.n59 B 0.012319f
C179 VDD1.n60 B 0.022926f
C180 VDD1.n61 B 0.022926f
C181 VDD1.n62 B 0.012319f
C182 VDD1.n63 B 0.013044f
C183 VDD1.n64 B 0.029119f
C184 VDD1.n65 B 0.060849f
C185 VDD1.n66 B 0.013044f
C186 VDD1.n67 B 0.012319f
C187 VDD1.n68 B 0.049234f
C188 VDD1.n69 B 0.050988f
C189 VDD1.t1 B 0.119571f
C190 VDD1.t3 B 0.119571f
C191 VDD1.n70 B 1.00805f
C192 VDD1.n71 B 1.53319f
C193 VDD1.t2 B 0.119571f
C194 VDD1.t5 B 0.119571f
C195 VDD1.n72 B 1.00715f
C196 VDD1.n73 B 1.71527f
C197 VTAIL.t0 B 0.132786f
C198 VTAIL.t1 B 0.132786f
C199 VTAIL.n0 B 1.04584f
C200 VTAIL.n1 B 0.353731f
C201 VTAIL.n2 B 0.034412f
C202 VTAIL.n3 B 0.02546f
C203 VTAIL.n4 B 0.013681f
C204 VTAIL.n5 B 0.032337f
C205 VTAIL.n6 B 0.014486f
C206 VTAIL.n7 B 0.02546f
C207 VTAIL.n8 B 0.013681f
C208 VTAIL.n9 B 0.032337f
C209 VTAIL.n10 B 0.014486f
C210 VTAIL.n11 B 0.6761f
C211 VTAIL.n12 B 0.013681f
C212 VTAIL.t10 B 0.052658f
C213 VTAIL.n13 B 0.112581f
C214 VTAIL.n14 B 0.019102f
C215 VTAIL.n15 B 0.024253f
C216 VTAIL.n16 B 0.032337f
C217 VTAIL.n17 B 0.014486f
C218 VTAIL.n18 B 0.013681f
C219 VTAIL.n19 B 0.02546f
C220 VTAIL.n20 B 0.02546f
C221 VTAIL.n21 B 0.013681f
C222 VTAIL.n22 B 0.014486f
C223 VTAIL.n23 B 0.032337f
C224 VTAIL.n24 B 0.032337f
C225 VTAIL.n25 B 0.014486f
C226 VTAIL.n26 B 0.013681f
C227 VTAIL.n27 B 0.02546f
C228 VTAIL.n28 B 0.02546f
C229 VTAIL.n29 B 0.013681f
C230 VTAIL.n30 B 0.014486f
C231 VTAIL.n31 B 0.032337f
C232 VTAIL.n32 B 0.067574f
C233 VTAIL.n33 B 0.014486f
C234 VTAIL.n34 B 0.013681f
C235 VTAIL.n35 B 0.054676f
C236 VTAIL.n36 B 0.037428f
C237 VTAIL.n37 B 0.183115f
C238 VTAIL.t7 B 0.132786f
C239 VTAIL.t8 B 0.132786f
C240 VTAIL.n38 B 1.04584f
C241 VTAIL.n39 B 1.31079f
C242 VTAIL.t11 B 0.132786f
C243 VTAIL.t4 B 0.132786f
C244 VTAIL.n40 B 1.04584f
C245 VTAIL.n41 B 1.31078f
C246 VTAIL.n42 B 0.034412f
C247 VTAIL.n43 B 0.02546f
C248 VTAIL.n44 B 0.013681f
C249 VTAIL.n45 B 0.032337f
C250 VTAIL.n46 B 0.014486f
C251 VTAIL.n47 B 0.02546f
C252 VTAIL.n48 B 0.013681f
C253 VTAIL.n49 B 0.032337f
C254 VTAIL.n50 B 0.014486f
C255 VTAIL.n51 B 0.6761f
C256 VTAIL.n52 B 0.013681f
C257 VTAIL.t3 B 0.052658f
C258 VTAIL.n53 B 0.112581f
C259 VTAIL.n54 B 0.019102f
C260 VTAIL.n55 B 0.024253f
C261 VTAIL.n56 B 0.032337f
C262 VTAIL.n57 B 0.014486f
C263 VTAIL.n58 B 0.013681f
C264 VTAIL.n59 B 0.02546f
C265 VTAIL.n60 B 0.02546f
C266 VTAIL.n61 B 0.013681f
C267 VTAIL.n62 B 0.014486f
C268 VTAIL.n63 B 0.032337f
C269 VTAIL.n64 B 0.032337f
C270 VTAIL.n65 B 0.014486f
C271 VTAIL.n66 B 0.013681f
C272 VTAIL.n67 B 0.02546f
C273 VTAIL.n68 B 0.02546f
C274 VTAIL.n69 B 0.013681f
C275 VTAIL.n70 B 0.014486f
C276 VTAIL.n71 B 0.032337f
C277 VTAIL.n72 B 0.067574f
C278 VTAIL.n73 B 0.014486f
C279 VTAIL.n74 B 0.013681f
C280 VTAIL.n75 B 0.054676f
C281 VTAIL.n76 B 0.037428f
C282 VTAIL.n77 B 0.183115f
C283 VTAIL.t6 B 0.132786f
C284 VTAIL.t5 B 0.132786f
C285 VTAIL.n78 B 1.04584f
C286 VTAIL.n79 B 0.411539f
C287 VTAIL.n80 B 0.034412f
C288 VTAIL.n81 B 0.02546f
C289 VTAIL.n82 B 0.013681f
C290 VTAIL.n83 B 0.032337f
C291 VTAIL.n84 B 0.014486f
C292 VTAIL.n85 B 0.02546f
C293 VTAIL.n86 B 0.013681f
C294 VTAIL.n87 B 0.032337f
C295 VTAIL.n88 B 0.014486f
C296 VTAIL.n89 B 0.6761f
C297 VTAIL.n90 B 0.013681f
C298 VTAIL.t9 B 0.052658f
C299 VTAIL.n91 B 0.112581f
C300 VTAIL.n92 B 0.019102f
C301 VTAIL.n93 B 0.024253f
C302 VTAIL.n94 B 0.032337f
C303 VTAIL.n95 B 0.014486f
C304 VTAIL.n96 B 0.013681f
C305 VTAIL.n97 B 0.02546f
C306 VTAIL.n98 B 0.02546f
C307 VTAIL.n99 B 0.013681f
C308 VTAIL.n100 B 0.014486f
C309 VTAIL.n101 B 0.032337f
C310 VTAIL.n102 B 0.032337f
C311 VTAIL.n103 B 0.014486f
C312 VTAIL.n104 B 0.013681f
C313 VTAIL.n105 B 0.02546f
C314 VTAIL.n106 B 0.02546f
C315 VTAIL.n107 B 0.013681f
C316 VTAIL.n108 B 0.014486f
C317 VTAIL.n109 B 0.032337f
C318 VTAIL.n110 B 0.067574f
C319 VTAIL.n111 B 0.014486f
C320 VTAIL.n112 B 0.013681f
C321 VTAIL.n113 B 0.054676f
C322 VTAIL.n114 B 0.037428f
C323 VTAIL.n115 B 0.998904f
C324 VTAIL.n116 B 0.034412f
C325 VTAIL.n117 B 0.02546f
C326 VTAIL.n118 B 0.013681f
C327 VTAIL.n119 B 0.032337f
C328 VTAIL.n120 B 0.014486f
C329 VTAIL.n121 B 0.02546f
C330 VTAIL.n122 B 0.013681f
C331 VTAIL.n123 B 0.032337f
C332 VTAIL.n124 B 0.014486f
C333 VTAIL.n125 B 0.6761f
C334 VTAIL.n126 B 0.013681f
C335 VTAIL.t2 B 0.052658f
C336 VTAIL.n127 B 0.112581f
C337 VTAIL.n128 B 0.019102f
C338 VTAIL.n129 B 0.024253f
C339 VTAIL.n130 B 0.032337f
C340 VTAIL.n131 B 0.014486f
C341 VTAIL.n132 B 0.013681f
C342 VTAIL.n133 B 0.02546f
C343 VTAIL.n134 B 0.02546f
C344 VTAIL.n135 B 0.013681f
C345 VTAIL.n136 B 0.014486f
C346 VTAIL.n137 B 0.032337f
C347 VTAIL.n138 B 0.032337f
C348 VTAIL.n139 B 0.014486f
C349 VTAIL.n140 B 0.013681f
C350 VTAIL.n141 B 0.02546f
C351 VTAIL.n142 B 0.02546f
C352 VTAIL.n143 B 0.013681f
C353 VTAIL.n144 B 0.014486f
C354 VTAIL.n145 B 0.032337f
C355 VTAIL.n146 B 0.067574f
C356 VTAIL.n147 B 0.014486f
C357 VTAIL.n148 B 0.013681f
C358 VTAIL.n149 B 0.054676f
C359 VTAIL.n150 B 0.037428f
C360 VTAIL.n151 B 0.973267f
C361 VP.n0 B 0.044769f
C362 VP.t4 B 0.668305f
C363 VP.n1 B 0.275603f
C364 VP.n2 B 0.044769f
C365 VP.n3 B 0.044769f
C366 VP.t0 B 0.726249f
C367 VP.t3 B 0.668305f
C368 VP.n4 B 0.31531f
C369 VP.t5 B 0.747014f
C370 VP.n5 B 0.326987f
C371 VP.n6 B 0.183986f
C372 VP.n7 B 0.055624f
C373 VP.n8 B 0.013738f
C374 VP.n9 B 0.317211f
C375 VP.n10 B 1.52938f
C376 VP.n11 B 1.57223f
C377 VP.t1 B 0.726249f
C378 VP.n12 B 0.317211f
C379 VP.n13 B 0.013738f
C380 VP.n14 B 0.055624f
C381 VP.n15 B 0.044769f
C382 VP.n16 B 0.044769f
C383 VP.n17 B 0.055624f
C384 VP.n18 B 0.013738f
C385 VP.t2 B 0.726249f
C386 VP.n19 B 0.317211f
C387 VP.n20 B 0.034694f
.ends

