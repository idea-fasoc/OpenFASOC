* NGSPICE file created from diff_pair_sample_0466.ext - technology: sky130A

.subckt diff_pair_sample_0466 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2422_n3948# sky130_fd_pr__pfet_01v8 ad=5.811 pd=30.58 as=0 ps=0 w=14.9 l=3.3
X1 VDD2.t1 VN.t0 VTAIL.t3 w_n2422_n3948# sky130_fd_pr__pfet_01v8 ad=5.811 pd=30.58 as=5.811 ps=30.58 w=14.9 l=3.3
X2 B.t8 B.t6 B.t7 w_n2422_n3948# sky130_fd_pr__pfet_01v8 ad=5.811 pd=30.58 as=0 ps=0 w=14.9 l=3.3
X3 VDD1.t1 VP.t0 VTAIL.t0 w_n2422_n3948# sky130_fd_pr__pfet_01v8 ad=5.811 pd=30.58 as=5.811 ps=30.58 w=14.9 l=3.3
X4 B.t5 B.t3 B.t4 w_n2422_n3948# sky130_fd_pr__pfet_01v8 ad=5.811 pd=30.58 as=0 ps=0 w=14.9 l=3.3
X5 VDD2.t0 VN.t1 VTAIL.t2 w_n2422_n3948# sky130_fd_pr__pfet_01v8 ad=5.811 pd=30.58 as=5.811 ps=30.58 w=14.9 l=3.3
X6 VDD1.t0 VP.t1 VTAIL.t1 w_n2422_n3948# sky130_fd_pr__pfet_01v8 ad=5.811 pd=30.58 as=5.811 ps=30.58 w=14.9 l=3.3
X7 B.t2 B.t0 B.t1 w_n2422_n3948# sky130_fd_pr__pfet_01v8 ad=5.811 pd=30.58 as=0 ps=0 w=14.9 l=3.3
R0 B.n388 B.n387 585
R1 B.n386 B.n107 585
R2 B.n385 B.n384 585
R3 B.n383 B.n108 585
R4 B.n382 B.n381 585
R5 B.n380 B.n109 585
R6 B.n379 B.n378 585
R7 B.n377 B.n110 585
R8 B.n376 B.n375 585
R9 B.n374 B.n111 585
R10 B.n373 B.n372 585
R11 B.n371 B.n112 585
R12 B.n370 B.n369 585
R13 B.n368 B.n113 585
R14 B.n367 B.n366 585
R15 B.n365 B.n114 585
R16 B.n364 B.n363 585
R17 B.n362 B.n115 585
R18 B.n361 B.n360 585
R19 B.n359 B.n116 585
R20 B.n358 B.n357 585
R21 B.n356 B.n117 585
R22 B.n355 B.n354 585
R23 B.n353 B.n118 585
R24 B.n352 B.n351 585
R25 B.n350 B.n119 585
R26 B.n349 B.n348 585
R27 B.n347 B.n120 585
R28 B.n346 B.n345 585
R29 B.n344 B.n121 585
R30 B.n343 B.n342 585
R31 B.n341 B.n122 585
R32 B.n340 B.n339 585
R33 B.n338 B.n123 585
R34 B.n337 B.n336 585
R35 B.n335 B.n124 585
R36 B.n334 B.n333 585
R37 B.n332 B.n125 585
R38 B.n331 B.n330 585
R39 B.n329 B.n126 585
R40 B.n328 B.n327 585
R41 B.n326 B.n127 585
R42 B.n325 B.n324 585
R43 B.n323 B.n128 585
R44 B.n322 B.n321 585
R45 B.n320 B.n129 585
R46 B.n319 B.n318 585
R47 B.n317 B.n130 585
R48 B.n316 B.n315 585
R49 B.n314 B.n131 585
R50 B.n313 B.n312 585
R51 B.n308 B.n132 585
R52 B.n307 B.n306 585
R53 B.n305 B.n133 585
R54 B.n304 B.n303 585
R55 B.n302 B.n134 585
R56 B.n301 B.n300 585
R57 B.n299 B.n135 585
R58 B.n298 B.n297 585
R59 B.n296 B.n136 585
R60 B.n294 B.n293 585
R61 B.n292 B.n139 585
R62 B.n291 B.n290 585
R63 B.n289 B.n140 585
R64 B.n288 B.n287 585
R65 B.n286 B.n141 585
R66 B.n285 B.n284 585
R67 B.n283 B.n142 585
R68 B.n282 B.n281 585
R69 B.n280 B.n143 585
R70 B.n279 B.n278 585
R71 B.n277 B.n144 585
R72 B.n276 B.n275 585
R73 B.n274 B.n145 585
R74 B.n273 B.n272 585
R75 B.n271 B.n146 585
R76 B.n270 B.n269 585
R77 B.n268 B.n147 585
R78 B.n267 B.n266 585
R79 B.n265 B.n148 585
R80 B.n264 B.n263 585
R81 B.n262 B.n149 585
R82 B.n261 B.n260 585
R83 B.n259 B.n150 585
R84 B.n258 B.n257 585
R85 B.n256 B.n151 585
R86 B.n255 B.n254 585
R87 B.n253 B.n152 585
R88 B.n252 B.n251 585
R89 B.n250 B.n153 585
R90 B.n249 B.n248 585
R91 B.n247 B.n154 585
R92 B.n246 B.n245 585
R93 B.n244 B.n155 585
R94 B.n243 B.n242 585
R95 B.n241 B.n156 585
R96 B.n240 B.n239 585
R97 B.n238 B.n157 585
R98 B.n237 B.n236 585
R99 B.n235 B.n158 585
R100 B.n234 B.n233 585
R101 B.n232 B.n159 585
R102 B.n231 B.n230 585
R103 B.n229 B.n160 585
R104 B.n228 B.n227 585
R105 B.n226 B.n161 585
R106 B.n225 B.n224 585
R107 B.n223 B.n162 585
R108 B.n222 B.n221 585
R109 B.n220 B.n163 585
R110 B.n389 B.n106 585
R111 B.n391 B.n390 585
R112 B.n392 B.n105 585
R113 B.n394 B.n393 585
R114 B.n395 B.n104 585
R115 B.n397 B.n396 585
R116 B.n398 B.n103 585
R117 B.n400 B.n399 585
R118 B.n401 B.n102 585
R119 B.n403 B.n402 585
R120 B.n404 B.n101 585
R121 B.n406 B.n405 585
R122 B.n407 B.n100 585
R123 B.n409 B.n408 585
R124 B.n410 B.n99 585
R125 B.n412 B.n411 585
R126 B.n413 B.n98 585
R127 B.n415 B.n414 585
R128 B.n416 B.n97 585
R129 B.n418 B.n417 585
R130 B.n419 B.n96 585
R131 B.n421 B.n420 585
R132 B.n422 B.n95 585
R133 B.n424 B.n423 585
R134 B.n425 B.n94 585
R135 B.n427 B.n426 585
R136 B.n428 B.n93 585
R137 B.n430 B.n429 585
R138 B.n431 B.n92 585
R139 B.n433 B.n432 585
R140 B.n434 B.n91 585
R141 B.n436 B.n435 585
R142 B.n437 B.n90 585
R143 B.n439 B.n438 585
R144 B.n440 B.n89 585
R145 B.n442 B.n441 585
R146 B.n443 B.n88 585
R147 B.n445 B.n444 585
R148 B.n446 B.n87 585
R149 B.n448 B.n447 585
R150 B.n449 B.n86 585
R151 B.n451 B.n450 585
R152 B.n452 B.n85 585
R153 B.n454 B.n453 585
R154 B.n455 B.n84 585
R155 B.n457 B.n456 585
R156 B.n458 B.n83 585
R157 B.n460 B.n459 585
R158 B.n461 B.n82 585
R159 B.n463 B.n462 585
R160 B.n464 B.n81 585
R161 B.n466 B.n465 585
R162 B.n467 B.n80 585
R163 B.n469 B.n468 585
R164 B.n470 B.n79 585
R165 B.n472 B.n471 585
R166 B.n473 B.n78 585
R167 B.n475 B.n474 585
R168 B.n476 B.n77 585
R169 B.n478 B.n477 585
R170 B.n644 B.n643 585
R171 B.n642 B.n17 585
R172 B.n641 B.n640 585
R173 B.n639 B.n18 585
R174 B.n638 B.n637 585
R175 B.n636 B.n19 585
R176 B.n635 B.n634 585
R177 B.n633 B.n20 585
R178 B.n632 B.n631 585
R179 B.n630 B.n21 585
R180 B.n629 B.n628 585
R181 B.n627 B.n22 585
R182 B.n626 B.n625 585
R183 B.n624 B.n23 585
R184 B.n623 B.n622 585
R185 B.n621 B.n24 585
R186 B.n620 B.n619 585
R187 B.n618 B.n25 585
R188 B.n617 B.n616 585
R189 B.n615 B.n26 585
R190 B.n614 B.n613 585
R191 B.n612 B.n27 585
R192 B.n611 B.n610 585
R193 B.n609 B.n28 585
R194 B.n608 B.n607 585
R195 B.n606 B.n29 585
R196 B.n605 B.n604 585
R197 B.n603 B.n30 585
R198 B.n602 B.n601 585
R199 B.n600 B.n31 585
R200 B.n599 B.n598 585
R201 B.n597 B.n32 585
R202 B.n596 B.n595 585
R203 B.n594 B.n33 585
R204 B.n593 B.n592 585
R205 B.n591 B.n34 585
R206 B.n590 B.n589 585
R207 B.n588 B.n35 585
R208 B.n587 B.n586 585
R209 B.n585 B.n36 585
R210 B.n584 B.n583 585
R211 B.n582 B.n37 585
R212 B.n581 B.n580 585
R213 B.n579 B.n38 585
R214 B.n578 B.n577 585
R215 B.n576 B.n39 585
R216 B.n575 B.n574 585
R217 B.n573 B.n40 585
R218 B.n572 B.n571 585
R219 B.n570 B.n41 585
R220 B.n568 B.n567 585
R221 B.n566 B.n44 585
R222 B.n565 B.n564 585
R223 B.n563 B.n45 585
R224 B.n562 B.n561 585
R225 B.n560 B.n46 585
R226 B.n559 B.n558 585
R227 B.n557 B.n47 585
R228 B.n556 B.n555 585
R229 B.n554 B.n48 585
R230 B.n553 B.n552 585
R231 B.n551 B.n49 585
R232 B.n550 B.n549 585
R233 B.n548 B.n53 585
R234 B.n547 B.n546 585
R235 B.n545 B.n54 585
R236 B.n544 B.n543 585
R237 B.n542 B.n55 585
R238 B.n541 B.n540 585
R239 B.n539 B.n56 585
R240 B.n538 B.n537 585
R241 B.n536 B.n57 585
R242 B.n535 B.n534 585
R243 B.n533 B.n58 585
R244 B.n532 B.n531 585
R245 B.n530 B.n59 585
R246 B.n529 B.n528 585
R247 B.n527 B.n60 585
R248 B.n526 B.n525 585
R249 B.n524 B.n61 585
R250 B.n523 B.n522 585
R251 B.n521 B.n62 585
R252 B.n520 B.n519 585
R253 B.n518 B.n63 585
R254 B.n517 B.n516 585
R255 B.n515 B.n64 585
R256 B.n514 B.n513 585
R257 B.n512 B.n65 585
R258 B.n511 B.n510 585
R259 B.n509 B.n66 585
R260 B.n508 B.n507 585
R261 B.n506 B.n67 585
R262 B.n505 B.n504 585
R263 B.n503 B.n68 585
R264 B.n502 B.n501 585
R265 B.n500 B.n69 585
R266 B.n499 B.n498 585
R267 B.n497 B.n70 585
R268 B.n496 B.n495 585
R269 B.n494 B.n71 585
R270 B.n493 B.n492 585
R271 B.n491 B.n72 585
R272 B.n490 B.n489 585
R273 B.n488 B.n73 585
R274 B.n487 B.n486 585
R275 B.n485 B.n74 585
R276 B.n484 B.n483 585
R277 B.n482 B.n75 585
R278 B.n481 B.n480 585
R279 B.n479 B.n76 585
R280 B.n645 B.n16 585
R281 B.n647 B.n646 585
R282 B.n648 B.n15 585
R283 B.n650 B.n649 585
R284 B.n651 B.n14 585
R285 B.n653 B.n652 585
R286 B.n654 B.n13 585
R287 B.n656 B.n655 585
R288 B.n657 B.n12 585
R289 B.n659 B.n658 585
R290 B.n660 B.n11 585
R291 B.n662 B.n661 585
R292 B.n663 B.n10 585
R293 B.n665 B.n664 585
R294 B.n666 B.n9 585
R295 B.n668 B.n667 585
R296 B.n669 B.n8 585
R297 B.n671 B.n670 585
R298 B.n672 B.n7 585
R299 B.n674 B.n673 585
R300 B.n675 B.n6 585
R301 B.n677 B.n676 585
R302 B.n678 B.n5 585
R303 B.n680 B.n679 585
R304 B.n681 B.n4 585
R305 B.n683 B.n682 585
R306 B.n684 B.n3 585
R307 B.n686 B.n685 585
R308 B.n687 B.n0 585
R309 B.n2 B.n1 585
R310 B.n178 B.n177 585
R311 B.n180 B.n179 585
R312 B.n181 B.n176 585
R313 B.n183 B.n182 585
R314 B.n184 B.n175 585
R315 B.n186 B.n185 585
R316 B.n187 B.n174 585
R317 B.n189 B.n188 585
R318 B.n190 B.n173 585
R319 B.n192 B.n191 585
R320 B.n193 B.n172 585
R321 B.n195 B.n194 585
R322 B.n196 B.n171 585
R323 B.n198 B.n197 585
R324 B.n199 B.n170 585
R325 B.n201 B.n200 585
R326 B.n202 B.n169 585
R327 B.n204 B.n203 585
R328 B.n205 B.n168 585
R329 B.n207 B.n206 585
R330 B.n208 B.n167 585
R331 B.n210 B.n209 585
R332 B.n211 B.n166 585
R333 B.n213 B.n212 585
R334 B.n214 B.n165 585
R335 B.n216 B.n215 585
R336 B.n217 B.n164 585
R337 B.n219 B.n218 585
R338 B.n309 B.t10 498.411
R339 B.n50 B.t5 498.411
R340 B.n137 B.t7 498.411
R341 B.n42 B.t2 498.411
R342 B.n220 B.n219 482.89
R343 B.n387 B.n106 482.89
R344 B.n477 B.n76 482.89
R345 B.n645 B.n644 482.89
R346 B.n310 B.t11 428.012
R347 B.n51 B.t4 428.012
R348 B.n138 B.t8 428.012
R349 B.n43 B.t1 428.012
R350 B.n137 B.t6 317.721
R351 B.n309 B.t9 317.721
R352 B.n50 B.t3 317.721
R353 B.n42 B.t0 317.721
R354 B.n689 B.n688 256.663
R355 B.n688 B.n687 235.042
R356 B.n688 B.n2 235.042
R357 B.n221 B.n220 163.367
R358 B.n221 B.n162 163.367
R359 B.n225 B.n162 163.367
R360 B.n226 B.n225 163.367
R361 B.n227 B.n226 163.367
R362 B.n227 B.n160 163.367
R363 B.n231 B.n160 163.367
R364 B.n232 B.n231 163.367
R365 B.n233 B.n232 163.367
R366 B.n233 B.n158 163.367
R367 B.n237 B.n158 163.367
R368 B.n238 B.n237 163.367
R369 B.n239 B.n238 163.367
R370 B.n239 B.n156 163.367
R371 B.n243 B.n156 163.367
R372 B.n244 B.n243 163.367
R373 B.n245 B.n244 163.367
R374 B.n245 B.n154 163.367
R375 B.n249 B.n154 163.367
R376 B.n250 B.n249 163.367
R377 B.n251 B.n250 163.367
R378 B.n251 B.n152 163.367
R379 B.n255 B.n152 163.367
R380 B.n256 B.n255 163.367
R381 B.n257 B.n256 163.367
R382 B.n257 B.n150 163.367
R383 B.n261 B.n150 163.367
R384 B.n262 B.n261 163.367
R385 B.n263 B.n262 163.367
R386 B.n263 B.n148 163.367
R387 B.n267 B.n148 163.367
R388 B.n268 B.n267 163.367
R389 B.n269 B.n268 163.367
R390 B.n269 B.n146 163.367
R391 B.n273 B.n146 163.367
R392 B.n274 B.n273 163.367
R393 B.n275 B.n274 163.367
R394 B.n275 B.n144 163.367
R395 B.n279 B.n144 163.367
R396 B.n280 B.n279 163.367
R397 B.n281 B.n280 163.367
R398 B.n281 B.n142 163.367
R399 B.n285 B.n142 163.367
R400 B.n286 B.n285 163.367
R401 B.n287 B.n286 163.367
R402 B.n287 B.n140 163.367
R403 B.n291 B.n140 163.367
R404 B.n292 B.n291 163.367
R405 B.n293 B.n292 163.367
R406 B.n293 B.n136 163.367
R407 B.n298 B.n136 163.367
R408 B.n299 B.n298 163.367
R409 B.n300 B.n299 163.367
R410 B.n300 B.n134 163.367
R411 B.n304 B.n134 163.367
R412 B.n305 B.n304 163.367
R413 B.n306 B.n305 163.367
R414 B.n306 B.n132 163.367
R415 B.n313 B.n132 163.367
R416 B.n314 B.n313 163.367
R417 B.n315 B.n314 163.367
R418 B.n315 B.n130 163.367
R419 B.n319 B.n130 163.367
R420 B.n320 B.n319 163.367
R421 B.n321 B.n320 163.367
R422 B.n321 B.n128 163.367
R423 B.n325 B.n128 163.367
R424 B.n326 B.n325 163.367
R425 B.n327 B.n326 163.367
R426 B.n327 B.n126 163.367
R427 B.n331 B.n126 163.367
R428 B.n332 B.n331 163.367
R429 B.n333 B.n332 163.367
R430 B.n333 B.n124 163.367
R431 B.n337 B.n124 163.367
R432 B.n338 B.n337 163.367
R433 B.n339 B.n338 163.367
R434 B.n339 B.n122 163.367
R435 B.n343 B.n122 163.367
R436 B.n344 B.n343 163.367
R437 B.n345 B.n344 163.367
R438 B.n345 B.n120 163.367
R439 B.n349 B.n120 163.367
R440 B.n350 B.n349 163.367
R441 B.n351 B.n350 163.367
R442 B.n351 B.n118 163.367
R443 B.n355 B.n118 163.367
R444 B.n356 B.n355 163.367
R445 B.n357 B.n356 163.367
R446 B.n357 B.n116 163.367
R447 B.n361 B.n116 163.367
R448 B.n362 B.n361 163.367
R449 B.n363 B.n362 163.367
R450 B.n363 B.n114 163.367
R451 B.n367 B.n114 163.367
R452 B.n368 B.n367 163.367
R453 B.n369 B.n368 163.367
R454 B.n369 B.n112 163.367
R455 B.n373 B.n112 163.367
R456 B.n374 B.n373 163.367
R457 B.n375 B.n374 163.367
R458 B.n375 B.n110 163.367
R459 B.n379 B.n110 163.367
R460 B.n380 B.n379 163.367
R461 B.n381 B.n380 163.367
R462 B.n381 B.n108 163.367
R463 B.n385 B.n108 163.367
R464 B.n386 B.n385 163.367
R465 B.n387 B.n386 163.367
R466 B.n477 B.n476 163.367
R467 B.n476 B.n475 163.367
R468 B.n475 B.n78 163.367
R469 B.n471 B.n78 163.367
R470 B.n471 B.n470 163.367
R471 B.n470 B.n469 163.367
R472 B.n469 B.n80 163.367
R473 B.n465 B.n80 163.367
R474 B.n465 B.n464 163.367
R475 B.n464 B.n463 163.367
R476 B.n463 B.n82 163.367
R477 B.n459 B.n82 163.367
R478 B.n459 B.n458 163.367
R479 B.n458 B.n457 163.367
R480 B.n457 B.n84 163.367
R481 B.n453 B.n84 163.367
R482 B.n453 B.n452 163.367
R483 B.n452 B.n451 163.367
R484 B.n451 B.n86 163.367
R485 B.n447 B.n86 163.367
R486 B.n447 B.n446 163.367
R487 B.n446 B.n445 163.367
R488 B.n445 B.n88 163.367
R489 B.n441 B.n88 163.367
R490 B.n441 B.n440 163.367
R491 B.n440 B.n439 163.367
R492 B.n439 B.n90 163.367
R493 B.n435 B.n90 163.367
R494 B.n435 B.n434 163.367
R495 B.n434 B.n433 163.367
R496 B.n433 B.n92 163.367
R497 B.n429 B.n92 163.367
R498 B.n429 B.n428 163.367
R499 B.n428 B.n427 163.367
R500 B.n427 B.n94 163.367
R501 B.n423 B.n94 163.367
R502 B.n423 B.n422 163.367
R503 B.n422 B.n421 163.367
R504 B.n421 B.n96 163.367
R505 B.n417 B.n96 163.367
R506 B.n417 B.n416 163.367
R507 B.n416 B.n415 163.367
R508 B.n415 B.n98 163.367
R509 B.n411 B.n98 163.367
R510 B.n411 B.n410 163.367
R511 B.n410 B.n409 163.367
R512 B.n409 B.n100 163.367
R513 B.n405 B.n100 163.367
R514 B.n405 B.n404 163.367
R515 B.n404 B.n403 163.367
R516 B.n403 B.n102 163.367
R517 B.n399 B.n102 163.367
R518 B.n399 B.n398 163.367
R519 B.n398 B.n397 163.367
R520 B.n397 B.n104 163.367
R521 B.n393 B.n104 163.367
R522 B.n393 B.n392 163.367
R523 B.n392 B.n391 163.367
R524 B.n391 B.n106 163.367
R525 B.n644 B.n17 163.367
R526 B.n640 B.n17 163.367
R527 B.n640 B.n639 163.367
R528 B.n639 B.n638 163.367
R529 B.n638 B.n19 163.367
R530 B.n634 B.n19 163.367
R531 B.n634 B.n633 163.367
R532 B.n633 B.n632 163.367
R533 B.n632 B.n21 163.367
R534 B.n628 B.n21 163.367
R535 B.n628 B.n627 163.367
R536 B.n627 B.n626 163.367
R537 B.n626 B.n23 163.367
R538 B.n622 B.n23 163.367
R539 B.n622 B.n621 163.367
R540 B.n621 B.n620 163.367
R541 B.n620 B.n25 163.367
R542 B.n616 B.n25 163.367
R543 B.n616 B.n615 163.367
R544 B.n615 B.n614 163.367
R545 B.n614 B.n27 163.367
R546 B.n610 B.n27 163.367
R547 B.n610 B.n609 163.367
R548 B.n609 B.n608 163.367
R549 B.n608 B.n29 163.367
R550 B.n604 B.n29 163.367
R551 B.n604 B.n603 163.367
R552 B.n603 B.n602 163.367
R553 B.n602 B.n31 163.367
R554 B.n598 B.n31 163.367
R555 B.n598 B.n597 163.367
R556 B.n597 B.n596 163.367
R557 B.n596 B.n33 163.367
R558 B.n592 B.n33 163.367
R559 B.n592 B.n591 163.367
R560 B.n591 B.n590 163.367
R561 B.n590 B.n35 163.367
R562 B.n586 B.n35 163.367
R563 B.n586 B.n585 163.367
R564 B.n585 B.n584 163.367
R565 B.n584 B.n37 163.367
R566 B.n580 B.n37 163.367
R567 B.n580 B.n579 163.367
R568 B.n579 B.n578 163.367
R569 B.n578 B.n39 163.367
R570 B.n574 B.n39 163.367
R571 B.n574 B.n573 163.367
R572 B.n573 B.n572 163.367
R573 B.n572 B.n41 163.367
R574 B.n567 B.n41 163.367
R575 B.n567 B.n566 163.367
R576 B.n566 B.n565 163.367
R577 B.n565 B.n45 163.367
R578 B.n561 B.n45 163.367
R579 B.n561 B.n560 163.367
R580 B.n560 B.n559 163.367
R581 B.n559 B.n47 163.367
R582 B.n555 B.n47 163.367
R583 B.n555 B.n554 163.367
R584 B.n554 B.n553 163.367
R585 B.n553 B.n49 163.367
R586 B.n549 B.n49 163.367
R587 B.n549 B.n548 163.367
R588 B.n548 B.n547 163.367
R589 B.n547 B.n54 163.367
R590 B.n543 B.n54 163.367
R591 B.n543 B.n542 163.367
R592 B.n542 B.n541 163.367
R593 B.n541 B.n56 163.367
R594 B.n537 B.n56 163.367
R595 B.n537 B.n536 163.367
R596 B.n536 B.n535 163.367
R597 B.n535 B.n58 163.367
R598 B.n531 B.n58 163.367
R599 B.n531 B.n530 163.367
R600 B.n530 B.n529 163.367
R601 B.n529 B.n60 163.367
R602 B.n525 B.n60 163.367
R603 B.n525 B.n524 163.367
R604 B.n524 B.n523 163.367
R605 B.n523 B.n62 163.367
R606 B.n519 B.n62 163.367
R607 B.n519 B.n518 163.367
R608 B.n518 B.n517 163.367
R609 B.n517 B.n64 163.367
R610 B.n513 B.n64 163.367
R611 B.n513 B.n512 163.367
R612 B.n512 B.n511 163.367
R613 B.n511 B.n66 163.367
R614 B.n507 B.n66 163.367
R615 B.n507 B.n506 163.367
R616 B.n506 B.n505 163.367
R617 B.n505 B.n68 163.367
R618 B.n501 B.n68 163.367
R619 B.n501 B.n500 163.367
R620 B.n500 B.n499 163.367
R621 B.n499 B.n70 163.367
R622 B.n495 B.n70 163.367
R623 B.n495 B.n494 163.367
R624 B.n494 B.n493 163.367
R625 B.n493 B.n72 163.367
R626 B.n489 B.n72 163.367
R627 B.n489 B.n488 163.367
R628 B.n488 B.n487 163.367
R629 B.n487 B.n74 163.367
R630 B.n483 B.n74 163.367
R631 B.n483 B.n482 163.367
R632 B.n482 B.n481 163.367
R633 B.n481 B.n76 163.367
R634 B.n646 B.n645 163.367
R635 B.n646 B.n15 163.367
R636 B.n650 B.n15 163.367
R637 B.n651 B.n650 163.367
R638 B.n652 B.n651 163.367
R639 B.n652 B.n13 163.367
R640 B.n656 B.n13 163.367
R641 B.n657 B.n656 163.367
R642 B.n658 B.n657 163.367
R643 B.n658 B.n11 163.367
R644 B.n662 B.n11 163.367
R645 B.n663 B.n662 163.367
R646 B.n664 B.n663 163.367
R647 B.n664 B.n9 163.367
R648 B.n668 B.n9 163.367
R649 B.n669 B.n668 163.367
R650 B.n670 B.n669 163.367
R651 B.n670 B.n7 163.367
R652 B.n674 B.n7 163.367
R653 B.n675 B.n674 163.367
R654 B.n676 B.n675 163.367
R655 B.n676 B.n5 163.367
R656 B.n680 B.n5 163.367
R657 B.n681 B.n680 163.367
R658 B.n682 B.n681 163.367
R659 B.n682 B.n3 163.367
R660 B.n686 B.n3 163.367
R661 B.n687 B.n686 163.367
R662 B.n178 B.n2 163.367
R663 B.n179 B.n178 163.367
R664 B.n179 B.n176 163.367
R665 B.n183 B.n176 163.367
R666 B.n184 B.n183 163.367
R667 B.n185 B.n184 163.367
R668 B.n185 B.n174 163.367
R669 B.n189 B.n174 163.367
R670 B.n190 B.n189 163.367
R671 B.n191 B.n190 163.367
R672 B.n191 B.n172 163.367
R673 B.n195 B.n172 163.367
R674 B.n196 B.n195 163.367
R675 B.n197 B.n196 163.367
R676 B.n197 B.n170 163.367
R677 B.n201 B.n170 163.367
R678 B.n202 B.n201 163.367
R679 B.n203 B.n202 163.367
R680 B.n203 B.n168 163.367
R681 B.n207 B.n168 163.367
R682 B.n208 B.n207 163.367
R683 B.n209 B.n208 163.367
R684 B.n209 B.n166 163.367
R685 B.n213 B.n166 163.367
R686 B.n214 B.n213 163.367
R687 B.n215 B.n214 163.367
R688 B.n215 B.n164 163.367
R689 B.n219 B.n164 163.367
R690 B.n138 B.n137 70.4005
R691 B.n310 B.n309 70.4005
R692 B.n51 B.n50 70.4005
R693 B.n43 B.n42 70.4005
R694 B.n295 B.n138 59.5399
R695 B.n311 B.n310 59.5399
R696 B.n52 B.n51 59.5399
R697 B.n569 B.n43 59.5399
R698 B.n643 B.n16 31.3761
R699 B.n479 B.n478 31.3761
R700 B.n389 B.n388 31.3761
R701 B.n218 B.n163 31.3761
R702 B B.n689 18.0485
R703 B.n647 B.n16 10.6151
R704 B.n648 B.n647 10.6151
R705 B.n649 B.n648 10.6151
R706 B.n649 B.n14 10.6151
R707 B.n653 B.n14 10.6151
R708 B.n654 B.n653 10.6151
R709 B.n655 B.n654 10.6151
R710 B.n655 B.n12 10.6151
R711 B.n659 B.n12 10.6151
R712 B.n660 B.n659 10.6151
R713 B.n661 B.n660 10.6151
R714 B.n661 B.n10 10.6151
R715 B.n665 B.n10 10.6151
R716 B.n666 B.n665 10.6151
R717 B.n667 B.n666 10.6151
R718 B.n667 B.n8 10.6151
R719 B.n671 B.n8 10.6151
R720 B.n672 B.n671 10.6151
R721 B.n673 B.n672 10.6151
R722 B.n673 B.n6 10.6151
R723 B.n677 B.n6 10.6151
R724 B.n678 B.n677 10.6151
R725 B.n679 B.n678 10.6151
R726 B.n679 B.n4 10.6151
R727 B.n683 B.n4 10.6151
R728 B.n684 B.n683 10.6151
R729 B.n685 B.n684 10.6151
R730 B.n685 B.n0 10.6151
R731 B.n643 B.n642 10.6151
R732 B.n642 B.n641 10.6151
R733 B.n641 B.n18 10.6151
R734 B.n637 B.n18 10.6151
R735 B.n637 B.n636 10.6151
R736 B.n636 B.n635 10.6151
R737 B.n635 B.n20 10.6151
R738 B.n631 B.n20 10.6151
R739 B.n631 B.n630 10.6151
R740 B.n630 B.n629 10.6151
R741 B.n629 B.n22 10.6151
R742 B.n625 B.n22 10.6151
R743 B.n625 B.n624 10.6151
R744 B.n624 B.n623 10.6151
R745 B.n623 B.n24 10.6151
R746 B.n619 B.n24 10.6151
R747 B.n619 B.n618 10.6151
R748 B.n618 B.n617 10.6151
R749 B.n617 B.n26 10.6151
R750 B.n613 B.n26 10.6151
R751 B.n613 B.n612 10.6151
R752 B.n612 B.n611 10.6151
R753 B.n611 B.n28 10.6151
R754 B.n607 B.n28 10.6151
R755 B.n607 B.n606 10.6151
R756 B.n606 B.n605 10.6151
R757 B.n605 B.n30 10.6151
R758 B.n601 B.n30 10.6151
R759 B.n601 B.n600 10.6151
R760 B.n600 B.n599 10.6151
R761 B.n599 B.n32 10.6151
R762 B.n595 B.n32 10.6151
R763 B.n595 B.n594 10.6151
R764 B.n594 B.n593 10.6151
R765 B.n593 B.n34 10.6151
R766 B.n589 B.n34 10.6151
R767 B.n589 B.n588 10.6151
R768 B.n588 B.n587 10.6151
R769 B.n587 B.n36 10.6151
R770 B.n583 B.n36 10.6151
R771 B.n583 B.n582 10.6151
R772 B.n582 B.n581 10.6151
R773 B.n581 B.n38 10.6151
R774 B.n577 B.n38 10.6151
R775 B.n577 B.n576 10.6151
R776 B.n576 B.n575 10.6151
R777 B.n575 B.n40 10.6151
R778 B.n571 B.n40 10.6151
R779 B.n571 B.n570 10.6151
R780 B.n568 B.n44 10.6151
R781 B.n564 B.n44 10.6151
R782 B.n564 B.n563 10.6151
R783 B.n563 B.n562 10.6151
R784 B.n562 B.n46 10.6151
R785 B.n558 B.n46 10.6151
R786 B.n558 B.n557 10.6151
R787 B.n557 B.n556 10.6151
R788 B.n556 B.n48 10.6151
R789 B.n552 B.n551 10.6151
R790 B.n551 B.n550 10.6151
R791 B.n550 B.n53 10.6151
R792 B.n546 B.n53 10.6151
R793 B.n546 B.n545 10.6151
R794 B.n545 B.n544 10.6151
R795 B.n544 B.n55 10.6151
R796 B.n540 B.n55 10.6151
R797 B.n540 B.n539 10.6151
R798 B.n539 B.n538 10.6151
R799 B.n538 B.n57 10.6151
R800 B.n534 B.n57 10.6151
R801 B.n534 B.n533 10.6151
R802 B.n533 B.n532 10.6151
R803 B.n532 B.n59 10.6151
R804 B.n528 B.n59 10.6151
R805 B.n528 B.n527 10.6151
R806 B.n527 B.n526 10.6151
R807 B.n526 B.n61 10.6151
R808 B.n522 B.n61 10.6151
R809 B.n522 B.n521 10.6151
R810 B.n521 B.n520 10.6151
R811 B.n520 B.n63 10.6151
R812 B.n516 B.n63 10.6151
R813 B.n516 B.n515 10.6151
R814 B.n515 B.n514 10.6151
R815 B.n514 B.n65 10.6151
R816 B.n510 B.n65 10.6151
R817 B.n510 B.n509 10.6151
R818 B.n509 B.n508 10.6151
R819 B.n508 B.n67 10.6151
R820 B.n504 B.n67 10.6151
R821 B.n504 B.n503 10.6151
R822 B.n503 B.n502 10.6151
R823 B.n502 B.n69 10.6151
R824 B.n498 B.n69 10.6151
R825 B.n498 B.n497 10.6151
R826 B.n497 B.n496 10.6151
R827 B.n496 B.n71 10.6151
R828 B.n492 B.n71 10.6151
R829 B.n492 B.n491 10.6151
R830 B.n491 B.n490 10.6151
R831 B.n490 B.n73 10.6151
R832 B.n486 B.n73 10.6151
R833 B.n486 B.n485 10.6151
R834 B.n485 B.n484 10.6151
R835 B.n484 B.n75 10.6151
R836 B.n480 B.n75 10.6151
R837 B.n480 B.n479 10.6151
R838 B.n478 B.n77 10.6151
R839 B.n474 B.n77 10.6151
R840 B.n474 B.n473 10.6151
R841 B.n473 B.n472 10.6151
R842 B.n472 B.n79 10.6151
R843 B.n468 B.n79 10.6151
R844 B.n468 B.n467 10.6151
R845 B.n467 B.n466 10.6151
R846 B.n466 B.n81 10.6151
R847 B.n462 B.n81 10.6151
R848 B.n462 B.n461 10.6151
R849 B.n461 B.n460 10.6151
R850 B.n460 B.n83 10.6151
R851 B.n456 B.n83 10.6151
R852 B.n456 B.n455 10.6151
R853 B.n455 B.n454 10.6151
R854 B.n454 B.n85 10.6151
R855 B.n450 B.n85 10.6151
R856 B.n450 B.n449 10.6151
R857 B.n449 B.n448 10.6151
R858 B.n448 B.n87 10.6151
R859 B.n444 B.n87 10.6151
R860 B.n444 B.n443 10.6151
R861 B.n443 B.n442 10.6151
R862 B.n442 B.n89 10.6151
R863 B.n438 B.n89 10.6151
R864 B.n438 B.n437 10.6151
R865 B.n437 B.n436 10.6151
R866 B.n436 B.n91 10.6151
R867 B.n432 B.n91 10.6151
R868 B.n432 B.n431 10.6151
R869 B.n431 B.n430 10.6151
R870 B.n430 B.n93 10.6151
R871 B.n426 B.n93 10.6151
R872 B.n426 B.n425 10.6151
R873 B.n425 B.n424 10.6151
R874 B.n424 B.n95 10.6151
R875 B.n420 B.n95 10.6151
R876 B.n420 B.n419 10.6151
R877 B.n419 B.n418 10.6151
R878 B.n418 B.n97 10.6151
R879 B.n414 B.n97 10.6151
R880 B.n414 B.n413 10.6151
R881 B.n413 B.n412 10.6151
R882 B.n412 B.n99 10.6151
R883 B.n408 B.n99 10.6151
R884 B.n408 B.n407 10.6151
R885 B.n407 B.n406 10.6151
R886 B.n406 B.n101 10.6151
R887 B.n402 B.n101 10.6151
R888 B.n402 B.n401 10.6151
R889 B.n401 B.n400 10.6151
R890 B.n400 B.n103 10.6151
R891 B.n396 B.n103 10.6151
R892 B.n396 B.n395 10.6151
R893 B.n395 B.n394 10.6151
R894 B.n394 B.n105 10.6151
R895 B.n390 B.n105 10.6151
R896 B.n390 B.n389 10.6151
R897 B.n177 B.n1 10.6151
R898 B.n180 B.n177 10.6151
R899 B.n181 B.n180 10.6151
R900 B.n182 B.n181 10.6151
R901 B.n182 B.n175 10.6151
R902 B.n186 B.n175 10.6151
R903 B.n187 B.n186 10.6151
R904 B.n188 B.n187 10.6151
R905 B.n188 B.n173 10.6151
R906 B.n192 B.n173 10.6151
R907 B.n193 B.n192 10.6151
R908 B.n194 B.n193 10.6151
R909 B.n194 B.n171 10.6151
R910 B.n198 B.n171 10.6151
R911 B.n199 B.n198 10.6151
R912 B.n200 B.n199 10.6151
R913 B.n200 B.n169 10.6151
R914 B.n204 B.n169 10.6151
R915 B.n205 B.n204 10.6151
R916 B.n206 B.n205 10.6151
R917 B.n206 B.n167 10.6151
R918 B.n210 B.n167 10.6151
R919 B.n211 B.n210 10.6151
R920 B.n212 B.n211 10.6151
R921 B.n212 B.n165 10.6151
R922 B.n216 B.n165 10.6151
R923 B.n217 B.n216 10.6151
R924 B.n218 B.n217 10.6151
R925 B.n222 B.n163 10.6151
R926 B.n223 B.n222 10.6151
R927 B.n224 B.n223 10.6151
R928 B.n224 B.n161 10.6151
R929 B.n228 B.n161 10.6151
R930 B.n229 B.n228 10.6151
R931 B.n230 B.n229 10.6151
R932 B.n230 B.n159 10.6151
R933 B.n234 B.n159 10.6151
R934 B.n235 B.n234 10.6151
R935 B.n236 B.n235 10.6151
R936 B.n236 B.n157 10.6151
R937 B.n240 B.n157 10.6151
R938 B.n241 B.n240 10.6151
R939 B.n242 B.n241 10.6151
R940 B.n242 B.n155 10.6151
R941 B.n246 B.n155 10.6151
R942 B.n247 B.n246 10.6151
R943 B.n248 B.n247 10.6151
R944 B.n248 B.n153 10.6151
R945 B.n252 B.n153 10.6151
R946 B.n253 B.n252 10.6151
R947 B.n254 B.n253 10.6151
R948 B.n254 B.n151 10.6151
R949 B.n258 B.n151 10.6151
R950 B.n259 B.n258 10.6151
R951 B.n260 B.n259 10.6151
R952 B.n260 B.n149 10.6151
R953 B.n264 B.n149 10.6151
R954 B.n265 B.n264 10.6151
R955 B.n266 B.n265 10.6151
R956 B.n266 B.n147 10.6151
R957 B.n270 B.n147 10.6151
R958 B.n271 B.n270 10.6151
R959 B.n272 B.n271 10.6151
R960 B.n272 B.n145 10.6151
R961 B.n276 B.n145 10.6151
R962 B.n277 B.n276 10.6151
R963 B.n278 B.n277 10.6151
R964 B.n278 B.n143 10.6151
R965 B.n282 B.n143 10.6151
R966 B.n283 B.n282 10.6151
R967 B.n284 B.n283 10.6151
R968 B.n284 B.n141 10.6151
R969 B.n288 B.n141 10.6151
R970 B.n289 B.n288 10.6151
R971 B.n290 B.n289 10.6151
R972 B.n290 B.n139 10.6151
R973 B.n294 B.n139 10.6151
R974 B.n297 B.n296 10.6151
R975 B.n297 B.n135 10.6151
R976 B.n301 B.n135 10.6151
R977 B.n302 B.n301 10.6151
R978 B.n303 B.n302 10.6151
R979 B.n303 B.n133 10.6151
R980 B.n307 B.n133 10.6151
R981 B.n308 B.n307 10.6151
R982 B.n312 B.n308 10.6151
R983 B.n316 B.n131 10.6151
R984 B.n317 B.n316 10.6151
R985 B.n318 B.n317 10.6151
R986 B.n318 B.n129 10.6151
R987 B.n322 B.n129 10.6151
R988 B.n323 B.n322 10.6151
R989 B.n324 B.n323 10.6151
R990 B.n324 B.n127 10.6151
R991 B.n328 B.n127 10.6151
R992 B.n329 B.n328 10.6151
R993 B.n330 B.n329 10.6151
R994 B.n330 B.n125 10.6151
R995 B.n334 B.n125 10.6151
R996 B.n335 B.n334 10.6151
R997 B.n336 B.n335 10.6151
R998 B.n336 B.n123 10.6151
R999 B.n340 B.n123 10.6151
R1000 B.n341 B.n340 10.6151
R1001 B.n342 B.n341 10.6151
R1002 B.n342 B.n121 10.6151
R1003 B.n346 B.n121 10.6151
R1004 B.n347 B.n346 10.6151
R1005 B.n348 B.n347 10.6151
R1006 B.n348 B.n119 10.6151
R1007 B.n352 B.n119 10.6151
R1008 B.n353 B.n352 10.6151
R1009 B.n354 B.n353 10.6151
R1010 B.n354 B.n117 10.6151
R1011 B.n358 B.n117 10.6151
R1012 B.n359 B.n358 10.6151
R1013 B.n360 B.n359 10.6151
R1014 B.n360 B.n115 10.6151
R1015 B.n364 B.n115 10.6151
R1016 B.n365 B.n364 10.6151
R1017 B.n366 B.n365 10.6151
R1018 B.n366 B.n113 10.6151
R1019 B.n370 B.n113 10.6151
R1020 B.n371 B.n370 10.6151
R1021 B.n372 B.n371 10.6151
R1022 B.n372 B.n111 10.6151
R1023 B.n376 B.n111 10.6151
R1024 B.n377 B.n376 10.6151
R1025 B.n378 B.n377 10.6151
R1026 B.n378 B.n109 10.6151
R1027 B.n382 B.n109 10.6151
R1028 B.n383 B.n382 10.6151
R1029 B.n384 B.n383 10.6151
R1030 B.n384 B.n107 10.6151
R1031 B.n388 B.n107 10.6151
R1032 B.n570 B.n569 9.36635
R1033 B.n552 B.n52 9.36635
R1034 B.n295 B.n294 9.36635
R1035 B.n311 B.n131 9.36635
R1036 B.n689 B.n0 8.11757
R1037 B.n689 B.n1 8.11757
R1038 B.n569 B.n568 1.24928
R1039 B.n52 B.n48 1.24928
R1040 B.n296 B.n295 1.24928
R1041 B.n312 B.n311 1.24928
R1042 VN VN.t1 196.279
R1043 VN VN.t0 148.188
R1044 VTAIL.n322 VTAIL.n246 756.745
R1045 VTAIL.n76 VTAIL.n0 756.745
R1046 VTAIL.n240 VTAIL.n164 756.745
R1047 VTAIL.n158 VTAIL.n82 756.745
R1048 VTAIL.n273 VTAIL.n272 585
R1049 VTAIL.n270 VTAIL.n269 585
R1050 VTAIL.n279 VTAIL.n278 585
R1051 VTAIL.n281 VTAIL.n280 585
R1052 VTAIL.n266 VTAIL.n265 585
R1053 VTAIL.n287 VTAIL.n286 585
R1054 VTAIL.n290 VTAIL.n289 585
R1055 VTAIL.n288 VTAIL.n262 585
R1056 VTAIL.n295 VTAIL.n261 585
R1057 VTAIL.n297 VTAIL.n296 585
R1058 VTAIL.n299 VTAIL.n298 585
R1059 VTAIL.n258 VTAIL.n257 585
R1060 VTAIL.n305 VTAIL.n304 585
R1061 VTAIL.n307 VTAIL.n306 585
R1062 VTAIL.n254 VTAIL.n253 585
R1063 VTAIL.n313 VTAIL.n312 585
R1064 VTAIL.n315 VTAIL.n314 585
R1065 VTAIL.n250 VTAIL.n249 585
R1066 VTAIL.n321 VTAIL.n320 585
R1067 VTAIL.n323 VTAIL.n322 585
R1068 VTAIL.n27 VTAIL.n26 585
R1069 VTAIL.n24 VTAIL.n23 585
R1070 VTAIL.n33 VTAIL.n32 585
R1071 VTAIL.n35 VTAIL.n34 585
R1072 VTAIL.n20 VTAIL.n19 585
R1073 VTAIL.n41 VTAIL.n40 585
R1074 VTAIL.n44 VTAIL.n43 585
R1075 VTAIL.n42 VTAIL.n16 585
R1076 VTAIL.n49 VTAIL.n15 585
R1077 VTAIL.n51 VTAIL.n50 585
R1078 VTAIL.n53 VTAIL.n52 585
R1079 VTAIL.n12 VTAIL.n11 585
R1080 VTAIL.n59 VTAIL.n58 585
R1081 VTAIL.n61 VTAIL.n60 585
R1082 VTAIL.n8 VTAIL.n7 585
R1083 VTAIL.n67 VTAIL.n66 585
R1084 VTAIL.n69 VTAIL.n68 585
R1085 VTAIL.n4 VTAIL.n3 585
R1086 VTAIL.n75 VTAIL.n74 585
R1087 VTAIL.n77 VTAIL.n76 585
R1088 VTAIL.n241 VTAIL.n240 585
R1089 VTAIL.n239 VTAIL.n238 585
R1090 VTAIL.n168 VTAIL.n167 585
R1091 VTAIL.n233 VTAIL.n232 585
R1092 VTAIL.n231 VTAIL.n230 585
R1093 VTAIL.n172 VTAIL.n171 585
R1094 VTAIL.n225 VTAIL.n224 585
R1095 VTAIL.n223 VTAIL.n222 585
R1096 VTAIL.n176 VTAIL.n175 585
R1097 VTAIL.n217 VTAIL.n216 585
R1098 VTAIL.n215 VTAIL.n214 585
R1099 VTAIL.n213 VTAIL.n179 585
R1100 VTAIL.n183 VTAIL.n180 585
R1101 VTAIL.n208 VTAIL.n207 585
R1102 VTAIL.n206 VTAIL.n205 585
R1103 VTAIL.n185 VTAIL.n184 585
R1104 VTAIL.n200 VTAIL.n199 585
R1105 VTAIL.n198 VTAIL.n197 585
R1106 VTAIL.n189 VTAIL.n188 585
R1107 VTAIL.n192 VTAIL.n191 585
R1108 VTAIL.n159 VTAIL.n158 585
R1109 VTAIL.n157 VTAIL.n156 585
R1110 VTAIL.n86 VTAIL.n85 585
R1111 VTAIL.n151 VTAIL.n150 585
R1112 VTAIL.n149 VTAIL.n148 585
R1113 VTAIL.n90 VTAIL.n89 585
R1114 VTAIL.n143 VTAIL.n142 585
R1115 VTAIL.n141 VTAIL.n140 585
R1116 VTAIL.n94 VTAIL.n93 585
R1117 VTAIL.n135 VTAIL.n134 585
R1118 VTAIL.n133 VTAIL.n132 585
R1119 VTAIL.n131 VTAIL.n97 585
R1120 VTAIL.n101 VTAIL.n98 585
R1121 VTAIL.n126 VTAIL.n125 585
R1122 VTAIL.n124 VTAIL.n123 585
R1123 VTAIL.n103 VTAIL.n102 585
R1124 VTAIL.n118 VTAIL.n117 585
R1125 VTAIL.n116 VTAIL.n115 585
R1126 VTAIL.n107 VTAIL.n106 585
R1127 VTAIL.n110 VTAIL.n109 585
R1128 VTAIL.t3 VTAIL.n271 329.036
R1129 VTAIL.t1 VTAIL.n25 329.036
R1130 VTAIL.t0 VTAIL.n190 329.036
R1131 VTAIL.t2 VTAIL.n108 329.036
R1132 VTAIL.n272 VTAIL.n269 171.744
R1133 VTAIL.n279 VTAIL.n269 171.744
R1134 VTAIL.n280 VTAIL.n279 171.744
R1135 VTAIL.n280 VTAIL.n265 171.744
R1136 VTAIL.n287 VTAIL.n265 171.744
R1137 VTAIL.n289 VTAIL.n287 171.744
R1138 VTAIL.n289 VTAIL.n288 171.744
R1139 VTAIL.n288 VTAIL.n261 171.744
R1140 VTAIL.n297 VTAIL.n261 171.744
R1141 VTAIL.n298 VTAIL.n297 171.744
R1142 VTAIL.n298 VTAIL.n257 171.744
R1143 VTAIL.n305 VTAIL.n257 171.744
R1144 VTAIL.n306 VTAIL.n305 171.744
R1145 VTAIL.n306 VTAIL.n253 171.744
R1146 VTAIL.n313 VTAIL.n253 171.744
R1147 VTAIL.n314 VTAIL.n313 171.744
R1148 VTAIL.n314 VTAIL.n249 171.744
R1149 VTAIL.n321 VTAIL.n249 171.744
R1150 VTAIL.n322 VTAIL.n321 171.744
R1151 VTAIL.n26 VTAIL.n23 171.744
R1152 VTAIL.n33 VTAIL.n23 171.744
R1153 VTAIL.n34 VTAIL.n33 171.744
R1154 VTAIL.n34 VTAIL.n19 171.744
R1155 VTAIL.n41 VTAIL.n19 171.744
R1156 VTAIL.n43 VTAIL.n41 171.744
R1157 VTAIL.n43 VTAIL.n42 171.744
R1158 VTAIL.n42 VTAIL.n15 171.744
R1159 VTAIL.n51 VTAIL.n15 171.744
R1160 VTAIL.n52 VTAIL.n51 171.744
R1161 VTAIL.n52 VTAIL.n11 171.744
R1162 VTAIL.n59 VTAIL.n11 171.744
R1163 VTAIL.n60 VTAIL.n59 171.744
R1164 VTAIL.n60 VTAIL.n7 171.744
R1165 VTAIL.n67 VTAIL.n7 171.744
R1166 VTAIL.n68 VTAIL.n67 171.744
R1167 VTAIL.n68 VTAIL.n3 171.744
R1168 VTAIL.n75 VTAIL.n3 171.744
R1169 VTAIL.n76 VTAIL.n75 171.744
R1170 VTAIL.n240 VTAIL.n239 171.744
R1171 VTAIL.n239 VTAIL.n167 171.744
R1172 VTAIL.n232 VTAIL.n167 171.744
R1173 VTAIL.n232 VTAIL.n231 171.744
R1174 VTAIL.n231 VTAIL.n171 171.744
R1175 VTAIL.n224 VTAIL.n171 171.744
R1176 VTAIL.n224 VTAIL.n223 171.744
R1177 VTAIL.n223 VTAIL.n175 171.744
R1178 VTAIL.n216 VTAIL.n175 171.744
R1179 VTAIL.n216 VTAIL.n215 171.744
R1180 VTAIL.n215 VTAIL.n179 171.744
R1181 VTAIL.n183 VTAIL.n179 171.744
R1182 VTAIL.n207 VTAIL.n183 171.744
R1183 VTAIL.n207 VTAIL.n206 171.744
R1184 VTAIL.n206 VTAIL.n184 171.744
R1185 VTAIL.n199 VTAIL.n184 171.744
R1186 VTAIL.n199 VTAIL.n198 171.744
R1187 VTAIL.n198 VTAIL.n188 171.744
R1188 VTAIL.n191 VTAIL.n188 171.744
R1189 VTAIL.n158 VTAIL.n157 171.744
R1190 VTAIL.n157 VTAIL.n85 171.744
R1191 VTAIL.n150 VTAIL.n85 171.744
R1192 VTAIL.n150 VTAIL.n149 171.744
R1193 VTAIL.n149 VTAIL.n89 171.744
R1194 VTAIL.n142 VTAIL.n89 171.744
R1195 VTAIL.n142 VTAIL.n141 171.744
R1196 VTAIL.n141 VTAIL.n93 171.744
R1197 VTAIL.n134 VTAIL.n93 171.744
R1198 VTAIL.n134 VTAIL.n133 171.744
R1199 VTAIL.n133 VTAIL.n97 171.744
R1200 VTAIL.n101 VTAIL.n97 171.744
R1201 VTAIL.n125 VTAIL.n101 171.744
R1202 VTAIL.n125 VTAIL.n124 171.744
R1203 VTAIL.n124 VTAIL.n102 171.744
R1204 VTAIL.n117 VTAIL.n102 171.744
R1205 VTAIL.n117 VTAIL.n116 171.744
R1206 VTAIL.n116 VTAIL.n106 171.744
R1207 VTAIL.n109 VTAIL.n106 171.744
R1208 VTAIL.n272 VTAIL.t3 85.8723
R1209 VTAIL.n26 VTAIL.t1 85.8723
R1210 VTAIL.n191 VTAIL.t0 85.8723
R1211 VTAIL.n109 VTAIL.t2 85.8723
R1212 VTAIL.n163 VTAIL.n81 31.4703
R1213 VTAIL.n327 VTAIL.n326 30.246
R1214 VTAIL.n81 VTAIL.n80 30.246
R1215 VTAIL.n245 VTAIL.n244 30.246
R1216 VTAIL.n163 VTAIL.n162 30.246
R1217 VTAIL.n327 VTAIL.n245 28.341
R1218 VTAIL.n296 VTAIL.n295 13.1884
R1219 VTAIL.n50 VTAIL.n49 13.1884
R1220 VTAIL.n214 VTAIL.n213 13.1884
R1221 VTAIL.n132 VTAIL.n131 13.1884
R1222 VTAIL.n294 VTAIL.n262 12.8005
R1223 VTAIL.n299 VTAIL.n260 12.8005
R1224 VTAIL.n48 VTAIL.n16 12.8005
R1225 VTAIL.n53 VTAIL.n14 12.8005
R1226 VTAIL.n217 VTAIL.n178 12.8005
R1227 VTAIL.n212 VTAIL.n180 12.8005
R1228 VTAIL.n135 VTAIL.n96 12.8005
R1229 VTAIL.n130 VTAIL.n98 12.8005
R1230 VTAIL.n291 VTAIL.n290 12.0247
R1231 VTAIL.n300 VTAIL.n258 12.0247
R1232 VTAIL.n45 VTAIL.n44 12.0247
R1233 VTAIL.n54 VTAIL.n12 12.0247
R1234 VTAIL.n218 VTAIL.n176 12.0247
R1235 VTAIL.n209 VTAIL.n208 12.0247
R1236 VTAIL.n136 VTAIL.n94 12.0247
R1237 VTAIL.n127 VTAIL.n126 12.0247
R1238 VTAIL.n286 VTAIL.n264 11.249
R1239 VTAIL.n304 VTAIL.n303 11.249
R1240 VTAIL.n40 VTAIL.n18 11.249
R1241 VTAIL.n58 VTAIL.n57 11.249
R1242 VTAIL.n222 VTAIL.n221 11.249
R1243 VTAIL.n205 VTAIL.n182 11.249
R1244 VTAIL.n140 VTAIL.n139 11.249
R1245 VTAIL.n123 VTAIL.n100 11.249
R1246 VTAIL.n273 VTAIL.n271 10.7239
R1247 VTAIL.n27 VTAIL.n25 10.7239
R1248 VTAIL.n192 VTAIL.n190 10.7239
R1249 VTAIL.n110 VTAIL.n108 10.7239
R1250 VTAIL.n285 VTAIL.n266 10.4732
R1251 VTAIL.n307 VTAIL.n256 10.4732
R1252 VTAIL.n39 VTAIL.n20 10.4732
R1253 VTAIL.n61 VTAIL.n10 10.4732
R1254 VTAIL.n225 VTAIL.n174 10.4732
R1255 VTAIL.n204 VTAIL.n185 10.4732
R1256 VTAIL.n143 VTAIL.n92 10.4732
R1257 VTAIL.n122 VTAIL.n103 10.4732
R1258 VTAIL.n282 VTAIL.n281 9.69747
R1259 VTAIL.n308 VTAIL.n254 9.69747
R1260 VTAIL.n36 VTAIL.n35 9.69747
R1261 VTAIL.n62 VTAIL.n8 9.69747
R1262 VTAIL.n226 VTAIL.n172 9.69747
R1263 VTAIL.n201 VTAIL.n200 9.69747
R1264 VTAIL.n144 VTAIL.n90 9.69747
R1265 VTAIL.n119 VTAIL.n118 9.69747
R1266 VTAIL.n326 VTAIL.n325 9.45567
R1267 VTAIL.n80 VTAIL.n79 9.45567
R1268 VTAIL.n244 VTAIL.n243 9.45567
R1269 VTAIL.n162 VTAIL.n161 9.45567
R1270 VTAIL.n319 VTAIL.n318 9.3005
R1271 VTAIL.n248 VTAIL.n247 9.3005
R1272 VTAIL.n325 VTAIL.n324 9.3005
R1273 VTAIL.n252 VTAIL.n251 9.3005
R1274 VTAIL.n311 VTAIL.n310 9.3005
R1275 VTAIL.n309 VTAIL.n308 9.3005
R1276 VTAIL.n256 VTAIL.n255 9.3005
R1277 VTAIL.n303 VTAIL.n302 9.3005
R1278 VTAIL.n301 VTAIL.n300 9.3005
R1279 VTAIL.n260 VTAIL.n259 9.3005
R1280 VTAIL.n275 VTAIL.n274 9.3005
R1281 VTAIL.n277 VTAIL.n276 9.3005
R1282 VTAIL.n268 VTAIL.n267 9.3005
R1283 VTAIL.n283 VTAIL.n282 9.3005
R1284 VTAIL.n285 VTAIL.n284 9.3005
R1285 VTAIL.n264 VTAIL.n263 9.3005
R1286 VTAIL.n292 VTAIL.n291 9.3005
R1287 VTAIL.n294 VTAIL.n293 9.3005
R1288 VTAIL.n317 VTAIL.n316 9.3005
R1289 VTAIL.n73 VTAIL.n72 9.3005
R1290 VTAIL.n2 VTAIL.n1 9.3005
R1291 VTAIL.n79 VTAIL.n78 9.3005
R1292 VTAIL.n6 VTAIL.n5 9.3005
R1293 VTAIL.n65 VTAIL.n64 9.3005
R1294 VTAIL.n63 VTAIL.n62 9.3005
R1295 VTAIL.n10 VTAIL.n9 9.3005
R1296 VTAIL.n57 VTAIL.n56 9.3005
R1297 VTAIL.n55 VTAIL.n54 9.3005
R1298 VTAIL.n14 VTAIL.n13 9.3005
R1299 VTAIL.n29 VTAIL.n28 9.3005
R1300 VTAIL.n31 VTAIL.n30 9.3005
R1301 VTAIL.n22 VTAIL.n21 9.3005
R1302 VTAIL.n37 VTAIL.n36 9.3005
R1303 VTAIL.n39 VTAIL.n38 9.3005
R1304 VTAIL.n18 VTAIL.n17 9.3005
R1305 VTAIL.n46 VTAIL.n45 9.3005
R1306 VTAIL.n48 VTAIL.n47 9.3005
R1307 VTAIL.n71 VTAIL.n70 9.3005
R1308 VTAIL.n166 VTAIL.n165 9.3005
R1309 VTAIL.n237 VTAIL.n236 9.3005
R1310 VTAIL.n235 VTAIL.n234 9.3005
R1311 VTAIL.n170 VTAIL.n169 9.3005
R1312 VTAIL.n229 VTAIL.n228 9.3005
R1313 VTAIL.n227 VTAIL.n226 9.3005
R1314 VTAIL.n174 VTAIL.n173 9.3005
R1315 VTAIL.n221 VTAIL.n220 9.3005
R1316 VTAIL.n219 VTAIL.n218 9.3005
R1317 VTAIL.n178 VTAIL.n177 9.3005
R1318 VTAIL.n212 VTAIL.n211 9.3005
R1319 VTAIL.n210 VTAIL.n209 9.3005
R1320 VTAIL.n182 VTAIL.n181 9.3005
R1321 VTAIL.n204 VTAIL.n203 9.3005
R1322 VTAIL.n202 VTAIL.n201 9.3005
R1323 VTAIL.n187 VTAIL.n186 9.3005
R1324 VTAIL.n196 VTAIL.n195 9.3005
R1325 VTAIL.n194 VTAIL.n193 9.3005
R1326 VTAIL.n243 VTAIL.n242 9.3005
R1327 VTAIL.n112 VTAIL.n111 9.3005
R1328 VTAIL.n114 VTAIL.n113 9.3005
R1329 VTAIL.n105 VTAIL.n104 9.3005
R1330 VTAIL.n120 VTAIL.n119 9.3005
R1331 VTAIL.n122 VTAIL.n121 9.3005
R1332 VTAIL.n100 VTAIL.n99 9.3005
R1333 VTAIL.n128 VTAIL.n127 9.3005
R1334 VTAIL.n130 VTAIL.n129 9.3005
R1335 VTAIL.n84 VTAIL.n83 9.3005
R1336 VTAIL.n161 VTAIL.n160 9.3005
R1337 VTAIL.n155 VTAIL.n154 9.3005
R1338 VTAIL.n153 VTAIL.n152 9.3005
R1339 VTAIL.n88 VTAIL.n87 9.3005
R1340 VTAIL.n147 VTAIL.n146 9.3005
R1341 VTAIL.n145 VTAIL.n144 9.3005
R1342 VTAIL.n92 VTAIL.n91 9.3005
R1343 VTAIL.n139 VTAIL.n138 9.3005
R1344 VTAIL.n137 VTAIL.n136 9.3005
R1345 VTAIL.n96 VTAIL.n95 9.3005
R1346 VTAIL.n278 VTAIL.n268 8.92171
R1347 VTAIL.n312 VTAIL.n311 8.92171
R1348 VTAIL.n326 VTAIL.n246 8.92171
R1349 VTAIL.n32 VTAIL.n22 8.92171
R1350 VTAIL.n66 VTAIL.n65 8.92171
R1351 VTAIL.n80 VTAIL.n0 8.92171
R1352 VTAIL.n244 VTAIL.n164 8.92171
R1353 VTAIL.n230 VTAIL.n229 8.92171
R1354 VTAIL.n197 VTAIL.n187 8.92171
R1355 VTAIL.n162 VTAIL.n82 8.92171
R1356 VTAIL.n148 VTAIL.n147 8.92171
R1357 VTAIL.n115 VTAIL.n105 8.92171
R1358 VTAIL.n277 VTAIL.n270 8.14595
R1359 VTAIL.n315 VTAIL.n252 8.14595
R1360 VTAIL.n324 VTAIL.n323 8.14595
R1361 VTAIL.n31 VTAIL.n24 8.14595
R1362 VTAIL.n69 VTAIL.n6 8.14595
R1363 VTAIL.n78 VTAIL.n77 8.14595
R1364 VTAIL.n242 VTAIL.n241 8.14595
R1365 VTAIL.n233 VTAIL.n170 8.14595
R1366 VTAIL.n196 VTAIL.n189 8.14595
R1367 VTAIL.n160 VTAIL.n159 8.14595
R1368 VTAIL.n151 VTAIL.n88 8.14595
R1369 VTAIL.n114 VTAIL.n107 8.14595
R1370 VTAIL.n274 VTAIL.n273 7.3702
R1371 VTAIL.n316 VTAIL.n250 7.3702
R1372 VTAIL.n320 VTAIL.n248 7.3702
R1373 VTAIL.n28 VTAIL.n27 7.3702
R1374 VTAIL.n70 VTAIL.n4 7.3702
R1375 VTAIL.n74 VTAIL.n2 7.3702
R1376 VTAIL.n238 VTAIL.n166 7.3702
R1377 VTAIL.n234 VTAIL.n168 7.3702
R1378 VTAIL.n193 VTAIL.n192 7.3702
R1379 VTAIL.n156 VTAIL.n84 7.3702
R1380 VTAIL.n152 VTAIL.n86 7.3702
R1381 VTAIL.n111 VTAIL.n110 7.3702
R1382 VTAIL.n319 VTAIL.n250 6.59444
R1383 VTAIL.n320 VTAIL.n319 6.59444
R1384 VTAIL.n73 VTAIL.n4 6.59444
R1385 VTAIL.n74 VTAIL.n73 6.59444
R1386 VTAIL.n238 VTAIL.n237 6.59444
R1387 VTAIL.n237 VTAIL.n168 6.59444
R1388 VTAIL.n156 VTAIL.n155 6.59444
R1389 VTAIL.n155 VTAIL.n86 6.59444
R1390 VTAIL.n274 VTAIL.n270 5.81868
R1391 VTAIL.n316 VTAIL.n315 5.81868
R1392 VTAIL.n323 VTAIL.n248 5.81868
R1393 VTAIL.n28 VTAIL.n24 5.81868
R1394 VTAIL.n70 VTAIL.n69 5.81868
R1395 VTAIL.n77 VTAIL.n2 5.81868
R1396 VTAIL.n241 VTAIL.n166 5.81868
R1397 VTAIL.n234 VTAIL.n233 5.81868
R1398 VTAIL.n193 VTAIL.n189 5.81868
R1399 VTAIL.n159 VTAIL.n84 5.81868
R1400 VTAIL.n152 VTAIL.n151 5.81868
R1401 VTAIL.n111 VTAIL.n107 5.81868
R1402 VTAIL.n278 VTAIL.n277 5.04292
R1403 VTAIL.n312 VTAIL.n252 5.04292
R1404 VTAIL.n324 VTAIL.n246 5.04292
R1405 VTAIL.n32 VTAIL.n31 5.04292
R1406 VTAIL.n66 VTAIL.n6 5.04292
R1407 VTAIL.n78 VTAIL.n0 5.04292
R1408 VTAIL.n242 VTAIL.n164 5.04292
R1409 VTAIL.n230 VTAIL.n170 5.04292
R1410 VTAIL.n197 VTAIL.n196 5.04292
R1411 VTAIL.n160 VTAIL.n82 5.04292
R1412 VTAIL.n148 VTAIL.n88 5.04292
R1413 VTAIL.n115 VTAIL.n114 5.04292
R1414 VTAIL.n281 VTAIL.n268 4.26717
R1415 VTAIL.n311 VTAIL.n254 4.26717
R1416 VTAIL.n35 VTAIL.n22 4.26717
R1417 VTAIL.n65 VTAIL.n8 4.26717
R1418 VTAIL.n229 VTAIL.n172 4.26717
R1419 VTAIL.n200 VTAIL.n187 4.26717
R1420 VTAIL.n147 VTAIL.n90 4.26717
R1421 VTAIL.n118 VTAIL.n105 4.26717
R1422 VTAIL.n282 VTAIL.n266 3.49141
R1423 VTAIL.n308 VTAIL.n307 3.49141
R1424 VTAIL.n36 VTAIL.n20 3.49141
R1425 VTAIL.n62 VTAIL.n61 3.49141
R1426 VTAIL.n226 VTAIL.n225 3.49141
R1427 VTAIL.n201 VTAIL.n185 3.49141
R1428 VTAIL.n144 VTAIL.n143 3.49141
R1429 VTAIL.n119 VTAIL.n103 3.49141
R1430 VTAIL.n286 VTAIL.n285 2.71565
R1431 VTAIL.n304 VTAIL.n256 2.71565
R1432 VTAIL.n40 VTAIL.n39 2.71565
R1433 VTAIL.n58 VTAIL.n10 2.71565
R1434 VTAIL.n222 VTAIL.n174 2.71565
R1435 VTAIL.n205 VTAIL.n204 2.71565
R1436 VTAIL.n140 VTAIL.n92 2.71565
R1437 VTAIL.n123 VTAIL.n122 2.71565
R1438 VTAIL.n194 VTAIL.n190 2.41282
R1439 VTAIL.n112 VTAIL.n108 2.41282
R1440 VTAIL.n275 VTAIL.n271 2.41282
R1441 VTAIL.n29 VTAIL.n25 2.41282
R1442 VTAIL.n245 VTAIL.n163 2.03498
R1443 VTAIL.n290 VTAIL.n264 1.93989
R1444 VTAIL.n303 VTAIL.n258 1.93989
R1445 VTAIL.n44 VTAIL.n18 1.93989
R1446 VTAIL.n57 VTAIL.n12 1.93989
R1447 VTAIL.n221 VTAIL.n176 1.93989
R1448 VTAIL.n208 VTAIL.n182 1.93989
R1449 VTAIL.n139 VTAIL.n94 1.93989
R1450 VTAIL.n126 VTAIL.n100 1.93989
R1451 VTAIL VTAIL.n81 1.31084
R1452 VTAIL.n291 VTAIL.n262 1.16414
R1453 VTAIL.n300 VTAIL.n299 1.16414
R1454 VTAIL.n45 VTAIL.n16 1.16414
R1455 VTAIL.n54 VTAIL.n53 1.16414
R1456 VTAIL.n218 VTAIL.n217 1.16414
R1457 VTAIL.n209 VTAIL.n180 1.16414
R1458 VTAIL.n136 VTAIL.n135 1.16414
R1459 VTAIL.n127 VTAIL.n98 1.16414
R1460 VTAIL VTAIL.n327 0.724638
R1461 VTAIL.n295 VTAIL.n294 0.388379
R1462 VTAIL.n296 VTAIL.n260 0.388379
R1463 VTAIL.n49 VTAIL.n48 0.388379
R1464 VTAIL.n50 VTAIL.n14 0.388379
R1465 VTAIL.n214 VTAIL.n178 0.388379
R1466 VTAIL.n213 VTAIL.n212 0.388379
R1467 VTAIL.n132 VTAIL.n96 0.388379
R1468 VTAIL.n131 VTAIL.n130 0.388379
R1469 VTAIL.n276 VTAIL.n275 0.155672
R1470 VTAIL.n276 VTAIL.n267 0.155672
R1471 VTAIL.n283 VTAIL.n267 0.155672
R1472 VTAIL.n284 VTAIL.n283 0.155672
R1473 VTAIL.n284 VTAIL.n263 0.155672
R1474 VTAIL.n292 VTAIL.n263 0.155672
R1475 VTAIL.n293 VTAIL.n292 0.155672
R1476 VTAIL.n293 VTAIL.n259 0.155672
R1477 VTAIL.n301 VTAIL.n259 0.155672
R1478 VTAIL.n302 VTAIL.n301 0.155672
R1479 VTAIL.n302 VTAIL.n255 0.155672
R1480 VTAIL.n309 VTAIL.n255 0.155672
R1481 VTAIL.n310 VTAIL.n309 0.155672
R1482 VTAIL.n310 VTAIL.n251 0.155672
R1483 VTAIL.n317 VTAIL.n251 0.155672
R1484 VTAIL.n318 VTAIL.n317 0.155672
R1485 VTAIL.n318 VTAIL.n247 0.155672
R1486 VTAIL.n325 VTAIL.n247 0.155672
R1487 VTAIL.n30 VTAIL.n29 0.155672
R1488 VTAIL.n30 VTAIL.n21 0.155672
R1489 VTAIL.n37 VTAIL.n21 0.155672
R1490 VTAIL.n38 VTAIL.n37 0.155672
R1491 VTAIL.n38 VTAIL.n17 0.155672
R1492 VTAIL.n46 VTAIL.n17 0.155672
R1493 VTAIL.n47 VTAIL.n46 0.155672
R1494 VTAIL.n47 VTAIL.n13 0.155672
R1495 VTAIL.n55 VTAIL.n13 0.155672
R1496 VTAIL.n56 VTAIL.n55 0.155672
R1497 VTAIL.n56 VTAIL.n9 0.155672
R1498 VTAIL.n63 VTAIL.n9 0.155672
R1499 VTAIL.n64 VTAIL.n63 0.155672
R1500 VTAIL.n64 VTAIL.n5 0.155672
R1501 VTAIL.n71 VTAIL.n5 0.155672
R1502 VTAIL.n72 VTAIL.n71 0.155672
R1503 VTAIL.n72 VTAIL.n1 0.155672
R1504 VTAIL.n79 VTAIL.n1 0.155672
R1505 VTAIL.n243 VTAIL.n165 0.155672
R1506 VTAIL.n236 VTAIL.n165 0.155672
R1507 VTAIL.n236 VTAIL.n235 0.155672
R1508 VTAIL.n235 VTAIL.n169 0.155672
R1509 VTAIL.n228 VTAIL.n169 0.155672
R1510 VTAIL.n228 VTAIL.n227 0.155672
R1511 VTAIL.n227 VTAIL.n173 0.155672
R1512 VTAIL.n220 VTAIL.n173 0.155672
R1513 VTAIL.n220 VTAIL.n219 0.155672
R1514 VTAIL.n219 VTAIL.n177 0.155672
R1515 VTAIL.n211 VTAIL.n177 0.155672
R1516 VTAIL.n211 VTAIL.n210 0.155672
R1517 VTAIL.n210 VTAIL.n181 0.155672
R1518 VTAIL.n203 VTAIL.n181 0.155672
R1519 VTAIL.n203 VTAIL.n202 0.155672
R1520 VTAIL.n202 VTAIL.n186 0.155672
R1521 VTAIL.n195 VTAIL.n186 0.155672
R1522 VTAIL.n195 VTAIL.n194 0.155672
R1523 VTAIL.n161 VTAIL.n83 0.155672
R1524 VTAIL.n154 VTAIL.n83 0.155672
R1525 VTAIL.n154 VTAIL.n153 0.155672
R1526 VTAIL.n153 VTAIL.n87 0.155672
R1527 VTAIL.n146 VTAIL.n87 0.155672
R1528 VTAIL.n146 VTAIL.n145 0.155672
R1529 VTAIL.n145 VTAIL.n91 0.155672
R1530 VTAIL.n138 VTAIL.n91 0.155672
R1531 VTAIL.n138 VTAIL.n137 0.155672
R1532 VTAIL.n137 VTAIL.n95 0.155672
R1533 VTAIL.n129 VTAIL.n95 0.155672
R1534 VTAIL.n129 VTAIL.n128 0.155672
R1535 VTAIL.n128 VTAIL.n99 0.155672
R1536 VTAIL.n121 VTAIL.n99 0.155672
R1537 VTAIL.n121 VTAIL.n120 0.155672
R1538 VTAIL.n120 VTAIL.n104 0.155672
R1539 VTAIL.n113 VTAIL.n104 0.155672
R1540 VTAIL.n113 VTAIL.n112 0.155672
R1541 VDD2.n157 VDD2.n81 756.745
R1542 VDD2.n76 VDD2.n0 756.745
R1543 VDD2.n158 VDD2.n157 585
R1544 VDD2.n156 VDD2.n155 585
R1545 VDD2.n85 VDD2.n84 585
R1546 VDD2.n150 VDD2.n149 585
R1547 VDD2.n148 VDD2.n147 585
R1548 VDD2.n89 VDD2.n88 585
R1549 VDD2.n142 VDD2.n141 585
R1550 VDD2.n140 VDD2.n139 585
R1551 VDD2.n93 VDD2.n92 585
R1552 VDD2.n134 VDD2.n133 585
R1553 VDD2.n132 VDD2.n131 585
R1554 VDD2.n130 VDD2.n96 585
R1555 VDD2.n100 VDD2.n97 585
R1556 VDD2.n125 VDD2.n124 585
R1557 VDD2.n123 VDD2.n122 585
R1558 VDD2.n102 VDD2.n101 585
R1559 VDD2.n117 VDD2.n116 585
R1560 VDD2.n115 VDD2.n114 585
R1561 VDD2.n106 VDD2.n105 585
R1562 VDD2.n109 VDD2.n108 585
R1563 VDD2.n27 VDD2.n26 585
R1564 VDD2.n24 VDD2.n23 585
R1565 VDD2.n33 VDD2.n32 585
R1566 VDD2.n35 VDD2.n34 585
R1567 VDD2.n20 VDD2.n19 585
R1568 VDD2.n41 VDD2.n40 585
R1569 VDD2.n44 VDD2.n43 585
R1570 VDD2.n42 VDD2.n16 585
R1571 VDD2.n49 VDD2.n15 585
R1572 VDD2.n51 VDD2.n50 585
R1573 VDD2.n53 VDD2.n52 585
R1574 VDD2.n12 VDD2.n11 585
R1575 VDD2.n59 VDD2.n58 585
R1576 VDD2.n61 VDD2.n60 585
R1577 VDD2.n8 VDD2.n7 585
R1578 VDD2.n67 VDD2.n66 585
R1579 VDD2.n69 VDD2.n68 585
R1580 VDD2.n4 VDD2.n3 585
R1581 VDD2.n75 VDD2.n74 585
R1582 VDD2.n77 VDD2.n76 585
R1583 VDD2.t0 VDD2.n107 329.036
R1584 VDD2.t1 VDD2.n25 329.036
R1585 VDD2.n157 VDD2.n156 171.744
R1586 VDD2.n156 VDD2.n84 171.744
R1587 VDD2.n149 VDD2.n84 171.744
R1588 VDD2.n149 VDD2.n148 171.744
R1589 VDD2.n148 VDD2.n88 171.744
R1590 VDD2.n141 VDD2.n88 171.744
R1591 VDD2.n141 VDD2.n140 171.744
R1592 VDD2.n140 VDD2.n92 171.744
R1593 VDD2.n133 VDD2.n92 171.744
R1594 VDD2.n133 VDD2.n132 171.744
R1595 VDD2.n132 VDD2.n96 171.744
R1596 VDD2.n100 VDD2.n96 171.744
R1597 VDD2.n124 VDD2.n100 171.744
R1598 VDD2.n124 VDD2.n123 171.744
R1599 VDD2.n123 VDD2.n101 171.744
R1600 VDD2.n116 VDD2.n101 171.744
R1601 VDD2.n116 VDD2.n115 171.744
R1602 VDD2.n115 VDD2.n105 171.744
R1603 VDD2.n108 VDD2.n105 171.744
R1604 VDD2.n26 VDD2.n23 171.744
R1605 VDD2.n33 VDD2.n23 171.744
R1606 VDD2.n34 VDD2.n33 171.744
R1607 VDD2.n34 VDD2.n19 171.744
R1608 VDD2.n41 VDD2.n19 171.744
R1609 VDD2.n43 VDD2.n41 171.744
R1610 VDD2.n43 VDD2.n42 171.744
R1611 VDD2.n42 VDD2.n15 171.744
R1612 VDD2.n51 VDD2.n15 171.744
R1613 VDD2.n52 VDD2.n51 171.744
R1614 VDD2.n52 VDD2.n11 171.744
R1615 VDD2.n59 VDD2.n11 171.744
R1616 VDD2.n60 VDD2.n59 171.744
R1617 VDD2.n60 VDD2.n7 171.744
R1618 VDD2.n67 VDD2.n7 171.744
R1619 VDD2.n68 VDD2.n67 171.744
R1620 VDD2.n68 VDD2.n3 171.744
R1621 VDD2.n75 VDD2.n3 171.744
R1622 VDD2.n76 VDD2.n75 171.744
R1623 VDD2.n162 VDD2.n80 89.6876
R1624 VDD2.n108 VDD2.t0 85.8723
R1625 VDD2.n26 VDD2.t1 85.8723
R1626 VDD2.n162 VDD2.n161 46.9247
R1627 VDD2.n131 VDD2.n130 13.1884
R1628 VDD2.n50 VDD2.n49 13.1884
R1629 VDD2.n134 VDD2.n95 12.8005
R1630 VDD2.n129 VDD2.n97 12.8005
R1631 VDD2.n48 VDD2.n16 12.8005
R1632 VDD2.n53 VDD2.n14 12.8005
R1633 VDD2.n135 VDD2.n93 12.0247
R1634 VDD2.n126 VDD2.n125 12.0247
R1635 VDD2.n45 VDD2.n44 12.0247
R1636 VDD2.n54 VDD2.n12 12.0247
R1637 VDD2.n139 VDD2.n138 11.249
R1638 VDD2.n122 VDD2.n99 11.249
R1639 VDD2.n40 VDD2.n18 11.249
R1640 VDD2.n58 VDD2.n57 11.249
R1641 VDD2.n109 VDD2.n107 10.7239
R1642 VDD2.n27 VDD2.n25 10.7239
R1643 VDD2.n142 VDD2.n91 10.4732
R1644 VDD2.n121 VDD2.n102 10.4732
R1645 VDD2.n39 VDD2.n20 10.4732
R1646 VDD2.n61 VDD2.n10 10.4732
R1647 VDD2.n143 VDD2.n89 9.69747
R1648 VDD2.n118 VDD2.n117 9.69747
R1649 VDD2.n36 VDD2.n35 9.69747
R1650 VDD2.n62 VDD2.n8 9.69747
R1651 VDD2.n161 VDD2.n160 9.45567
R1652 VDD2.n80 VDD2.n79 9.45567
R1653 VDD2.n83 VDD2.n82 9.3005
R1654 VDD2.n154 VDD2.n153 9.3005
R1655 VDD2.n152 VDD2.n151 9.3005
R1656 VDD2.n87 VDD2.n86 9.3005
R1657 VDD2.n146 VDD2.n145 9.3005
R1658 VDD2.n144 VDD2.n143 9.3005
R1659 VDD2.n91 VDD2.n90 9.3005
R1660 VDD2.n138 VDD2.n137 9.3005
R1661 VDD2.n136 VDD2.n135 9.3005
R1662 VDD2.n95 VDD2.n94 9.3005
R1663 VDD2.n129 VDD2.n128 9.3005
R1664 VDD2.n127 VDD2.n126 9.3005
R1665 VDD2.n99 VDD2.n98 9.3005
R1666 VDD2.n121 VDD2.n120 9.3005
R1667 VDD2.n119 VDD2.n118 9.3005
R1668 VDD2.n104 VDD2.n103 9.3005
R1669 VDD2.n113 VDD2.n112 9.3005
R1670 VDD2.n111 VDD2.n110 9.3005
R1671 VDD2.n160 VDD2.n159 9.3005
R1672 VDD2.n73 VDD2.n72 9.3005
R1673 VDD2.n2 VDD2.n1 9.3005
R1674 VDD2.n79 VDD2.n78 9.3005
R1675 VDD2.n6 VDD2.n5 9.3005
R1676 VDD2.n65 VDD2.n64 9.3005
R1677 VDD2.n63 VDD2.n62 9.3005
R1678 VDD2.n10 VDD2.n9 9.3005
R1679 VDD2.n57 VDD2.n56 9.3005
R1680 VDD2.n55 VDD2.n54 9.3005
R1681 VDD2.n14 VDD2.n13 9.3005
R1682 VDD2.n29 VDD2.n28 9.3005
R1683 VDD2.n31 VDD2.n30 9.3005
R1684 VDD2.n22 VDD2.n21 9.3005
R1685 VDD2.n37 VDD2.n36 9.3005
R1686 VDD2.n39 VDD2.n38 9.3005
R1687 VDD2.n18 VDD2.n17 9.3005
R1688 VDD2.n46 VDD2.n45 9.3005
R1689 VDD2.n48 VDD2.n47 9.3005
R1690 VDD2.n71 VDD2.n70 9.3005
R1691 VDD2.n161 VDD2.n81 8.92171
R1692 VDD2.n147 VDD2.n146 8.92171
R1693 VDD2.n114 VDD2.n104 8.92171
R1694 VDD2.n32 VDD2.n22 8.92171
R1695 VDD2.n66 VDD2.n65 8.92171
R1696 VDD2.n80 VDD2.n0 8.92171
R1697 VDD2.n159 VDD2.n158 8.14595
R1698 VDD2.n150 VDD2.n87 8.14595
R1699 VDD2.n113 VDD2.n106 8.14595
R1700 VDD2.n31 VDD2.n24 8.14595
R1701 VDD2.n69 VDD2.n6 8.14595
R1702 VDD2.n78 VDD2.n77 8.14595
R1703 VDD2.n155 VDD2.n83 7.3702
R1704 VDD2.n151 VDD2.n85 7.3702
R1705 VDD2.n110 VDD2.n109 7.3702
R1706 VDD2.n28 VDD2.n27 7.3702
R1707 VDD2.n70 VDD2.n4 7.3702
R1708 VDD2.n74 VDD2.n2 7.3702
R1709 VDD2.n155 VDD2.n154 6.59444
R1710 VDD2.n154 VDD2.n85 6.59444
R1711 VDD2.n73 VDD2.n4 6.59444
R1712 VDD2.n74 VDD2.n73 6.59444
R1713 VDD2.n158 VDD2.n83 5.81868
R1714 VDD2.n151 VDD2.n150 5.81868
R1715 VDD2.n110 VDD2.n106 5.81868
R1716 VDD2.n28 VDD2.n24 5.81868
R1717 VDD2.n70 VDD2.n69 5.81868
R1718 VDD2.n77 VDD2.n2 5.81868
R1719 VDD2.n159 VDD2.n81 5.04292
R1720 VDD2.n147 VDD2.n87 5.04292
R1721 VDD2.n114 VDD2.n113 5.04292
R1722 VDD2.n32 VDD2.n31 5.04292
R1723 VDD2.n66 VDD2.n6 5.04292
R1724 VDD2.n78 VDD2.n0 5.04292
R1725 VDD2.n146 VDD2.n89 4.26717
R1726 VDD2.n117 VDD2.n104 4.26717
R1727 VDD2.n35 VDD2.n22 4.26717
R1728 VDD2.n65 VDD2.n8 4.26717
R1729 VDD2.n143 VDD2.n142 3.49141
R1730 VDD2.n118 VDD2.n102 3.49141
R1731 VDD2.n36 VDD2.n20 3.49141
R1732 VDD2.n62 VDD2.n61 3.49141
R1733 VDD2.n139 VDD2.n91 2.71565
R1734 VDD2.n122 VDD2.n121 2.71565
R1735 VDD2.n40 VDD2.n39 2.71565
R1736 VDD2.n58 VDD2.n10 2.71565
R1737 VDD2.n111 VDD2.n107 2.41282
R1738 VDD2.n29 VDD2.n25 2.41282
R1739 VDD2.n138 VDD2.n93 1.93989
R1740 VDD2.n125 VDD2.n99 1.93989
R1741 VDD2.n44 VDD2.n18 1.93989
R1742 VDD2.n57 VDD2.n12 1.93989
R1743 VDD2.n135 VDD2.n134 1.16414
R1744 VDD2.n126 VDD2.n97 1.16414
R1745 VDD2.n45 VDD2.n16 1.16414
R1746 VDD2.n54 VDD2.n53 1.16414
R1747 VDD2 VDD2.n162 0.841017
R1748 VDD2.n131 VDD2.n95 0.388379
R1749 VDD2.n130 VDD2.n129 0.388379
R1750 VDD2.n49 VDD2.n48 0.388379
R1751 VDD2.n50 VDD2.n14 0.388379
R1752 VDD2.n160 VDD2.n82 0.155672
R1753 VDD2.n153 VDD2.n82 0.155672
R1754 VDD2.n153 VDD2.n152 0.155672
R1755 VDD2.n152 VDD2.n86 0.155672
R1756 VDD2.n145 VDD2.n86 0.155672
R1757 VDD2.n145 VDD2.n144 0.155672
R1758 VDD2.n144 VDD2.n90 0.155672
R1759 VDD2.n137 VDD2.n90 0.155672
R1760 VDD2.n137 VDD2.n136 0.155672
R1761 VDD2.n136 VDD2.n94 0.155672
R1762 VDD2.n128 VDD2.n94 0.155672
R1763 VDD2.n128 VDD2.n127 0.155672
R1764 VDD2.n127 VDD2.n98 0.155672
R1765 VDD2.n120 VDD2.n98 0.155672
R1766 VDD2.n120 VDD2.n119 0.155672
R1767 VDD2.n119 VDD2.n103 0.155672
R1768 VDD2.n112 VDD2.n103 0.155672
R1769 VDD2.n112 VDD2.n111 0.155672
R1770 VDD2.n30 VDD2.n29 0.155672
R1771 VDD2.n30 VDD2.n21 0.155672
R1772 VDD2.n37 VDD2.n21 0.155672
R1773 VDD2.n38 VDD2.n37 0.155672
R1774 VDD2.n38 VDD2.n17 0.155672
R1775 VDD2.n46 VDD2.n17 0.155672
R1776 VDD2.n47 VDD2.n46 0.155672
R1777 VDD2.n47 VDD2.n13 0.155672
R1778 VDD2.n55 VDD2.n13 0.155672
R1779 VDD2.n56 VDD2.n55 0.155672
R1780 VDD2.n56 VDD2.n9 0.155672
R1781 VDD2.n63 VDD2.n9 0.155672
R1782 VDD2.n64 VDD2.n63 0.155672
R1783 VDD2.n64 VDD2.n5 0.155672
R1784 VDD2.n71 VDD2.n5 0.155672
R1785 VDD2.n72 VDD2.n71 0.155672
R1786 VDD2.n72 VDD2.n1 0.155672
R1787 VDD2.n79 VDD2.n1 0.155672
R1788 VP.n0 VP.t0 196.37
R1789 VP.n0 VP.t1 147.661
R1790 VP VP.n0 0.526373
R1791 VDD1.n76 VDD1.n0 756.745
R1792 VDD1.n157 VDD1.n81 756.745
R1793 VDD1.n77 VDD1.n76 585
R1794 VDD1.n75 VDD1.n74 585
R1795 VDD1.n4 VDD1.n3 585
R1796 VDD1.n69 VDD1.n68 585
R1797 VDD1.n67 VDD1.n66 585
R1798 VDD1.n8 VDD1.n7 585
R1799 VDD1.n61 VDD1.n60 585
R1800 VDD1.n59 VDD1.n58 585
R1801 VDD1.n12 VDD1.n11 585
R1802 VDD1.n53 VDD1.n52 585
R1803 VDD1.n51 VDD1.n50 585
R1804 VDD1.n49 VDD1.n15 585
R1805 VDD1.n19 VDD1.n16 585
R1806 VDD1.n44 VDD1.n43 585
R1807 VDD1.n42 VDD1.n41 585
R1808 VDD1.n21 VDD1.n20 585
R1809 VDD1.n36 VDD1.n35 585
R1810 VDD1.n34 VDD1.n33 585
R1811 VDD1.n25 VDD1.n24 585
R1812 VDD1.n28 VDD1.n27 585
R1813 VDD1.n108 VDD1.n107 585
R1814 VDD1.n105 VDD1.n104 585
R1815 VDD1.n114 VDD1.n113 585
R1816 VDD1.n116 VDD1.n115 585
R1817 VDD1.n101 VDD1.n100 585
R1818 VDD1.n122 VDD1.n121 585
R1819 VDD1.n125 VDD1.n124 585
R1820 VDD1.n123 VDD1.n97 585
R1821 VDD1.n130 VDD1.n96 585
R1822 VDD1.n132 VDD1.n131 585
R1823 VDD1.n134 VDD1.n133 585
R1824 VDD1.n93 VDD1.n92 585
R1825 VDD1.n140 VDD1.n139 585
R1826 VDD1.n142 VDD1.n141 585
R1827 VDD1.n89 VDD1.n88 585
R1828 VDD1.n148 VDD1.n147 585
R1829 VDD1.n150 VDD1.n149 585
R1830 VDD1.n85 VDD1.n84 585
R1831 VDD1.n156 VDD1.n155 585
R1832 VDD1.n158 VDD1.n157 585
R1833 VDD1.t1 VDD1.n26 329.036
R1834 VDD1.t0 VDD1.n106 329.036
R1835 VDD1.n76 VDD1.n75 171.744
R1836 VDD1.n75 VDD1.n3 171.744
R1837 VDD1.n68 VDD1.n3 171.744
R1838 VDD1.n68 VDD1.n67 171.744
R1839 VDD1.n67 VDD1.n7 171.744
R1840 VDD1.n60 VDD1.n7 171.744
R1841 VDD1.n60 VDD1.n59 171.744
R1842 VDD1.n59 VDD1.n11 171.744
R1843 VDD1.n52 VDD1.n11 171.744
R1844 VDD1.n52 VDD1.n51 171.744
R1845 VDD1.n51 VDD1.n15 171.744
R1846 VDD1.n19 VDD1.n15 171.744
R1847 VDD1.n43 VDD1.n19 171.744
R1848 VDD1.n43 VDD1.n42 171.744
R1849 VDD1.n42 VDD1.n20 171.744
R1850 VDD1.n35 VDD1.n20 171.744
R1851 VDD1.n35 VDD1.n34 171.744
R1852 VDD1.n34 VDD1.n24 171.744
R1853 VDD1.n27 VDD1.n24 171.744
R1854 VDD1.n107 VDD1.n104 171.744
R1855 VDD1.n114 VDD1.n104 171.744
R1856 VDD1.n115 VDD1.n114 171.744
R1857 VDD1.n115 VDD1.n100 171.744
R1858 VDD1.n122 VDD1.n100 171.744
R1859 VDD1.n124 VDD1.n122 171.744
R1860 VDD1.n124 VDD1.n123 171.744
R1861 VDD1.n123 VDD1.n96 171.744
R1862 VDD1.n132 VDD1.n96 171.744
R1863 VDD1.n133 VDD1.n132 171.744
R1864 VDD1.n133 VDD1.n92 171.744
R1865 VDD1.n140 VDD1.n92 171.744
R1866 VDD1.n141 VDD1.n140 171.744
R1867 VDD1.n141 VDD1.n88 171.744
R1868 VDD1.n148 VDD1.n88 171.744
R1869 VDD1.n149 VDD1.n148 171.744
R1870 VDD1.n149 VDD1.n84 171.744
R1871 VDD1.n156 VDD1.n84 171.744
R1872 VDD1.n157 VDD1.n156 171.744
R1873 VDD1 VDD1.n161 90.9948
R1874 VDD1.n27 VDD1.t1 85.8723
R1875 VDD1.n107 VDD1.t0 85.8723
R1876 VDD1 VDD1.n80 47.7653
R1877 VDD1.n50 VDD1.n49 13.1884
R1878 VDD1.n131 VDD1.n130 13.1884
R1879 VDD1.n53 VDD1.n14 12.8005
R1880 VDD1.n48 VDD1.n16 12.8005
R1881 VDD1.n129 VDD1.n97 12.8005
R1882 VDD1.n134 VDD1.n95 12.8005
R1883 VDD1.n54 VDD1.n12 12.0247
R1884 VDD1.n45 VDD1.n44 12.0247
R1885 VDD1.n126 VDD1.n125 12.0247
R1886 VDD1.n135 VDD1.n93 12.0247
R1887 VDD1.n58 VDD1.n57 11.249
R1888 VDD1.n41 VDD1.n18 11.249
R1889 VDD1.n121 VDD1.n99 11.249
R1890 VDD1.n139 VDD1.n138 11.249
R1891 VDD1.n28 VDD1.n26 10.7239
R1892 VDD1.n108 VDD1.n106 10.7239
R1893 VDD1.n61 VDD1.n10 10.4732
R1894 VDD1.n40 VDD1.n21 10.4732
R1895 VDD1.n120 VDD1.n101 10.4732
R1896 VDD1.n142 VDD1.n91 10.4732
R1897 VDD1.n62 VDD1.n8 9.69747
R1898 VDD1.n37 VDD1.n36 9.69747
R1899 VDD1.n117 VDD1.n116 9.69747
R1900 VDD1.n143 VDD1.n89 9.69747
R1901 VDD1.n80 VDD1.n79 9.45567
R1902 VDD1.n161 VDD1.n160 9.45567
R1903 VDD1.n2 VDD1.n1 9.3005
R1904 VDD1.n73 VDD1.n72 9.3005
R1905 VDD1.n71 VDD1.n70 9.3005
R1906 VDD1.n6 VDD1.n5 9.3005
R1907 VDD1.n65 VDD1.n64 9.3005
R1908 VDD1.n63 VDD1.n62 9.3005
R1909 VDD1.n10 VDD1.n9 9.3005
R1910 VDD1.n57 VDD1.n56 9.3005
R1911 VDD1.n55 VDD1.n54 9.3005
R1912 VDD1.n14 VDD1.n13 9.3005
R1913 VDD1.n48 VDD1.n47 9.3005
R1914 VDD1.n46 VDD1.n45 9.3005
R1915 VDD1.n18 VDD1.n17 9.3005
R1916 VDD1.n40 VDD1.n39 9.3005
R1917 VDD1.n38 VDD1.n37 9.3005
R1918 VDD1.n23 VDD1.n22 9.3005
R1919 VDD1.n32 VDD1.n31 9.3005
R1920 VDD1.n30 VDD1.n29 9.3005
R1921 VDD1.n79 VDD1.n78 9.3005
R1922 VDD1.n154 VDD1.n153 9.3005
R1923 VDD1.n83 VDD1.n82 9.3005
R1924 VDD1.n160 VDD1.n159 9.3005
R1925 VDD1.n87 VDD1.n86 9.3005
R1926 VDD1.n146 VDD1.n145 9.3005
R1927 VDD1.n144 VDD1.n143 9.3005
R1928 VDD1.n91 VDD1.n90 9.3005
R1929 VDD1.n138 VDD1.n137 9.3005
R1930 VDD1.n136 VDD1.n135 9.3005
R1931 VDD1.n95 VDD1.n94 9.3005
R1932 VDD1.n110 VDD1.n109 9.3005
R1933 VDD1.n112 VDD1.n111 9.3005
R1934 VDD1.n103 VDD1.n102 9.3005
R1935 VDD1.n118 VDD1.n117 9.3005
R1936 VDD1.n120 VDD1.n119 9.3005
R1937 VDD1.n99 VDD1.n98 9.3005
R1938 VDD1.n127 VDD1.n126 9.3005
R1939 VDD1.n129 VDD1.n128 9.3005
R1940 VDD1.n152 VDD1.n151 9.3005
R1941 VDD1.n80 VDD1.n0 8.92171
R1942 VDD1.n66 VDD1.n65 8.92171
R1943 VDD1.n33 VDD1.n23 8.92171
R1944 VDD1.n113 VDD1.n103 8.92171
R1945 VDD1.n147 VDD1.n146 8.92171
R1946 VDD1.n161 VDD1.n81 8.92171
R1947 VDD1.n78 VDD1.n77 8.14595
R1948 VDD1.n69 VDD1.n6 8.14595
R1949 VDD1.n32 VDD1.n25 8.14595
R1950 VDD1.n112 VDD1.n105 8.14595
R1951 VDD1.n150 VDD1.n87 8.14595
R1952 VDD1.n159 VDD1.n158 8.14595
R1953 VDD1.n74 VDD1.n2 7.3702
R1954 VDD1.n70 VDD1.n4 7.3702
R1955 VDD1.n29 VDD1.n28 7.3702
R1956 VDD1.n109 VDD1.n108 7.3702
R1957 VDD1.n151 VDD1.n85 7.3702
R1958 VDD1.n155 VDD1.n83 7.3702
R1959 VDD1.n74 VDD1.n73 6.59444
R1960 VDD1.n73 VDD1.n4 6.59444
R1961 VDD1.n154 VDD1.n85 6.59444
R1962 VDD1.n155 VDD1.n154 6.59444
R1963 VDD1.n77 VDD1.n2 5.81868
R1964 VDD1.n70 VDD1.n69 5.81868
R1965 VDD1.n29 VDD1.n25 5.81868
R1966 VDD1.n109 VDD1.n105 5.81868
R1967 VDD1.n151 VDD1.n150 5.81868
R1968 VDD1.n158 VDD1.n83 5.81868
R1969 VDD1.n78 VDD1.n0 5.04292
R1970 VDD1.n66 VDD1.n6 5.04292
R1971 VDD1.n33 VDD1.n32 5.04292
R1972 VDD1.n113 VDD1.n112 5.04292
R1973 VDD1.n147 VDD1.n87 5.04292
R1974 VDD1.n159 VDD1.n81 5.04292
R1975 VDD1.n65 VDD1.n8 4.26717
R1976 VDD1.n36 VDD1.n23 4.26717
R1977 VDD1.n116 VDD1.n103 4.26717
R1978 VDD1.n146 VDD1.n89 4.26717
R1979 VDD1.n62 VDD1.n61 3.49141
R1980 VDD1.n37 VDD1.n21 3.49141
R1981 VDD1.n117 VDD1.n101 3.49141
R1982 VDD1.n143 VDD1.n142 3.49141
R1983 VDD1.n58 VDD1.n10 2.71565
R1984 VDD1.n41 VDD1.n40 2.71565
R1985 VDD1.n121 VDD1.n120 2.71565
R1986 VDD1.n139 VDD1.n91 2.71565
R1987 VDD1.n30 VDD1.n26 2.41282
R1988 VDD1.n110 VDD1.n106 2.41282
R1989 VDD1.n57 VDD1.n12 1.93989
R1990 VDD1.n44 VDD1.n18 1.93989
R1991 VDD1.n125 VDD1.n99 1.93989
R1992 VDD1.n138 VDD1.n93 1.93989
R1993 VDD1.n54 VDD1.n53 1.16414
R1994 VDD1.n45 VDD1.n16 1.16414
R1995 VDD1.n126 VDD1.n97 1.16414
R1996 VDD1.n135 VDD1.n134 1.16414
R1997 VDD1.n50 VDD1.n14 0.388379
R1998 VDD1.n49 VDD1.n48 0.388379
R1999 VDD1.n130 VDD1.n129 0.388379
R2000 VDD1.n131 VDD1.n95 0.388379
R2001 VDD1.n79 VDD1.n1 0.155672
R2002 VDD1.n72 VDD1.n1 0.155672
R2003 VDD1.n72 VDD1.n71 0.155672
R2004 VDD1.n71 VDD1.n5 0.155672
R2005 VDD1.n64 VDD1.n5 0.155672
R2006 VDD1.n64 VDD1.n63 0.155672
R2007 VDD1.n63 VDD1.n9 0.155672
R2008 VDD1.n56 VDD1.n9 0.155672
R2009 VDD1.n56 VDD1.n55 0.155672
R2010 VDD1.n55 VDD1.n13 0.155672
R2011 VDD1.n47 VDD1.n13 0.155672
R2012 VDD1.n47 VDD1.n46 0.155672
R2013 VDD1.n46 VDD1.n17 0.155672
R2014 VDD1.n39 VDD1.n17 0.155672
R2015 VDD1.n39 VDD1.n38 0.155672
R2016 VDD1.n38 VDD1.n22 0.155672
R2017 VDD1.n31 VDD1.n22 0.155672
R2018 VDD1.n31 VDD1.n30 0.155672
R2019 VDD1.n111 VDD1.n110 0.155672
R2020 VDD1.n111 VDD1.n102 0.155672
R2021 VDD1.n118 VDD1.n102 0.155672
R2022 VDD1.n119 VDD1.n118 0.155672
R2023 VDD1.n119 VDD1.n98 0.155672
R2024 VDD1.n127 VDD1.n98 0.155672
R2025 VDD1.n128 VDD1.n127 0.155672
R2026 VDD1.n128 VDD1.n94 0.155672
R2027 VDD1.n136 VDD1.n94 0.155672
R2028 VDD1.n137 VDD1.n136 0.155672
R2029 VDD1.n137 VDD1.n90 0.155672
R2030 VDD1.n144 VDD1.n90 0.155672
R2031 VDD1.n145 VDD1.n144 0.155672
R2032 VDD1.n145 VDD1.n86 0.155672
R2033 VDD1.n152 VDD1.n86 0.155672
R2034 VDD1.n153 VDD1.n152 0.155672
R2035 VDD1.n153 VDD1.n82 0.155672
R2036 VDD1.n160 VDD1.n82 0.155672
C0 VTAIL VDD1 5.9316f
C1 VP w_n2422_n3948# 3.77869f
C2 VP VTAIL 3.09857f
C3 VDD2 VN 3.50625f
C4 VDD2 w_n2422_n3948# 2.09386f
C5 VDD2 VTAIL 5.987f
C6 VDD1 B 2.03124f
C7 VN w_n2422_n3948# 3.46866f
C8 VN VTAIL 3.08429f
C9 VP B 1.71851f
C10 w_n2422_n3948# VTAIL 3.1553f
C11 VP VDD1 3.71782f
C12 VDD2 B 2.06755f
C13 VDD2 VDD1 0.760206f
C14 VN B 1.206f
C15 VN VDD1 0.148778f
C16 VDD2 VP 0.362997f
C17 w_n2422_n3948# B 10.378099f
C18 VTAIL B 4.59813f
C19 w_n2422_n3948# VDD1 2.0593f
C20 VN VP 6.31976f
C21 VDD2 VSUBS 1.101308f
C22 VDD1 VSUBS 5.42906f
C23 VTAIL VSUBS 1.191426f
C24 VN VSUBS 8.633201f
C25 VP VSUBS 1.998757f
C26 B VSUBS 4.668555f
C27 w_n2422_n3948# VSUBS 0.117273p
C28 VDD1.n0 VSUBS 0.032338f
C29 VDD1.n1 VSUBS 0.028873f
C30 VDD1.n2 VSUBS 0.015515f
C31 VDD1.n3 VSUBS 0.036672f
C32 VDD1.n4 VSUBS 0.016428f
C33 VDD1.n5 VSUBS 0.028873f
C34 VDD1.n6 VSUBS 0.015515f
C35 VDD1.n7 VSUBS 0.036672f
C36 VDD1.n8 VSUBS 0.016428f
C37 VDD1.n9 VSUBS 0.028873f
C38 VDD1.n10 VSUBS 0.015515f
C39 VDD1.n11 VSUBS 0.036672f
C40 VDD1.n12 VSUBS 0.016428f
C41 VDD1.n13 VSUBS 0.028873f
C42 VDD1.n14 VSUBS 0.015515f
C43 VDD1.n15 VSUBS 0.036672f
C44 VDD1.n16 VSUBS 0.016428f
C45 VDD1.n17 VSUBS 0.028873f
C46 VDD1.n18 VSUBS 0.015515f
C47 VDD1.n19 VSUBS 0.036672f
C48 VDD1.n20 VSUBS 0.036672f
C49 VDD1.n21 VSUBS 0.016428f
C50 VDD1.n22 VSUBS 0.028873f
C51 VDD1.n23 VSUBS 0.015515f
C52 VDD1.n24 VSUBS 0.036672f
C53 VDD1.n25 VSUBS 0.016428f
C54 VDD1.n26 VSUBS 0.265245f
C55 VDD1.t1 VSUBS 0.079303f
C56 VDD1.n27 VSUBS 0.027504f
C57 VDD1.n28 VSUBS 0.027586f
C58 VDD1.n29 VSUBS 0.015515f
C59 VDD1.n30 VSUBS 1.78548f
C60 VDD1.n31 VSUBS 0.028873f
C61 VDD1.n32 VSUBS 0.015515f
C62 VDD1.n33 VSUBS 0.016428f
C63 VDD1.n34 VSUBS 0.036672f
C64 VDD1.n35 VSUBS 0.036672f
C65 VDD1.n36 VSUBS 0.016428f
C66 VDD1.n37 VSUBS 0.015515f
C67 VDD1.n38 VSUBS 0.028873f
C68 VDD1.n39 VSUBS 0.028873f
C69 VDD1.n40 VSUBS 0.015515f
C70 VDD1.n41 VSUBS 0.016428f
C71 VDD1.n42 VSUBS 0.036672f
C72 VDD1.n43 VSUBS 0.036672f
C73 VDD1.n44 VSUBS 0.016428f
C74 VDD1.n45 VSUBS 0.015515f
C75 VDD1.n46 VSUBS 0.028873f
C76 VDD1.n47 VSUBS 0.028873f
C77 VDD1.n48 VSUBS 0.015515f
C78 VDD1.n49 VSUBS 0.015971f
C79 VDD1.n50 VSUBS 0.015971f
C80 VDD1.n51 VSUBS 0.036672f
C81 VDD1.n52 VSUBS 0.036672f
C82 VDD1.n53 VSUBS 0.016428f
C83 VDD1.n54 VSUBS 0.015515f
C84 VDD1.n55 VSUBS 0.028873f
C85 VDD1.n56 VSUBS 0.028873f
C86 VDD1.n57 VSUBS 0.015515f
C87 VDD1.n58 VSUBS 0.016428f
C88 VDD1.n59 VSUBS 0.036672f
C89 VDD1.n60 VSUBS 0.036672f
C90 VDD1.n61 VSUBS 0.016428f
C91 VDD1.n62 VSUBS 0.015515f
C92 VDD1.n63 VSUBS 0.028873f
C93 VDD1.n64 VSUBS 0.028873f
C94 VDD1.n65 VSUBS 0.015515f
C95 VDD1.n66 VSUBS 0.016428f
C96 VDD1.n67 VSUBS 0.036672f
C97 VDD1.n68 VSUBS 0.036672f
C98 VDD1.n69 VSUBS 0.016428f
C99 VDD1.n70 VSUBS 0.015515f
C100 VDD1.n71 VSUBS 0.028873f
C101 VDD1.n72 VSUBS 0.028873f
C102 VDD1.n73 VSUBS 0.015515f
C103 VDD1.n74 VSUBS 0.016428f
C104 VDD1.n75 VSUBS 0.036672f
C105 VDD1.n76 VSUBS 0.090868f
C106 VDD1.n77 VSUBS 0.016428f
C107 VDD1.n78 VSUBS 0.015515f
C108 VDD1.n79 VSUBS 0.062793f
C109 VDD1.n80 VSUBS 0.067949f
C110 VDD1.n81 VSUBS 0.032338f
C111 VDD1.n82 VSUBS 0.028873f
C112 VDD1.n83 VSUBS 0.015515f
C113 VDD1.n84 VSUBS 0.036672f
C114 VDD1.n85 VSUBS 0.016428f
C115 VDD1.n86 VSUBS 0.028873f
C116 VDD1.n87 VSUBS 0.015515f
C117 VDD1.n88 VSUBS 0.036672f
C118 VDD1.n89 VSUBS 0.016428f
C119 VDD1.n90 VSUBS 0.028873f
C120 VDD1.n91 VSUBS 0.015515f
C121 VDD1.n92 VSUBS 0.036672f
C122 VDD1.n93 VSUBS 0.016428f
C123 VDD1.n94 VSUBS 0.028873f
C124 VDD1.n95 VSUBS 0.015515f
C125 VDD1.n96 VSUBS 0.036672f
C126 VDD1.n97 VSUBS 0.016428f
C127 VDD1.n98 VSUBS 0.028873f
C128 VDD1.n99 VSUBS 0.015515f
C129 VDD1.n100 VSUBS 0.036672f
C130 VDD1.n101 VSUBS 0.016428f
C131 VDD1.n102 VSUBS 0.028873f
C132 VDD1.n103 VSUBS 0.015515f
C133 VDD1.n104 VSUBS 0.036672f
C134 VDD1.n105 VSUBS 0.016428f
C135 VDD1.n106 VSUBS 0.265245f
C136 VDD1.t0 VSUBS 0.079302f
C137 VDD1.n107 VSUBS 0.027504f
C138 VDD1.n108 VSUBS 0.027586f
C139 VDD1.n109 VSUBS 0.015515f
C140 VDD1.n110 VSUBS 1.78548f
C141 VDD1.n111 VSUBS 0.028873f
C142 VDD1.n112 VSUBS 0.015515f
C143 VDD1.n113 VSUBS 0.016428f
C144 VDD1.n114 VSUBS 0.036672f
C145 VDD1.n115 VSUBS 0.036672f
C146 VDD1.n116 VSUBS 0.016428f
C147 VDD1.n117 VSUBS 0.015515f
C148 VDD1.n118 VSUBS 0.028873f
C149 VDD1.n119 VSUBS 0.028873f
C150 VDD1.n120 VSUBS 0.015515f
C151 VDD1.n121 VSUBS 0.016428f
C152 VDD1.n122 VSUBS 0.036672f
C153 VDD1.n123 VSUBS 0.036672f
C154 VDD1.n124 VSUBS 0.036672f
C155 VDD1.n125 VSUBS 0.016428f
C156 VDD1.n126 VSUBS 0.015515f
C157 VDD1.n127 VSUBS 0.028873f
C158 VDD1.n128 VSUBS 0.028873f
C159 VDD1.n129 VSUBS 0.015515f
C160 VDD1.n130 VSUBS 0.015971f
C161 VDD1.n131 VSUBS 0.015971f
C162 VDD1.n132 VSUBS 0.036672f
C163 VDD1.n133 VSUBS 0.036672f
C164 VDD1.n134 VSUBS 0.016428f
C165 VDD1.n135 VSUBS 0.015515f
C166 VDD1.n136 VSUBS 0.028873f
C167 VDD1.n137 VSUBS 0.028873f
C168 VDD1.n138 VSUBS 0.015515f
C169 VDD1.n139 VSUBS 0.016428f
C170 VDD1.n140 VSUBS 0.036672f
C171 VDD1.n141 VSUBS 0.036672f
C172 VDD1.n142 VSUBS 0.016428f
C173 VDD1.n143 VSUBS 0.015515f
C174 VDD1.n144 VSUBS 0.028873f
C175 VDD1.n145 VSUBS 0.028873f
C176 VDD1.n146 VSUBS 0.015515f
C177 VDD1.n147 VSUBS 0.016428f
C178 VDD1.n148 VSUBS 0.036672f
C179 VDD1.n149 VSUBS 0.036672f
C180 VDD1.n150 VSUBS 0.016428f
C181 VDD1.n151 VSUBS 0.015515f
C182 VDD1.n152 VSUBS 0.028873f
C183 VDD1.n153 VSUBS 0.028873f
C184 VDD1.n154 VSUBS 0.015515f
C185 VDD1.n155 VSUBS 0.016428f
C186 VDD1.n156 VSUBS 0.036672f
C187 VDD1.n157 VSUBS 0.090868f
C188 VDD1.n158 VSUBS 0.016428f
C189 VDD1.n159 VSUBS 0.015515f
C190 VDD1.n160 VSUBS 0.062793f
C191 VDD1.n161 VSUBS 1.11564f
C192 VP.t0 VSUBS 5.89339f
C193 VP.t1 VSUBS 5.05415f
C194 VP.n0 VSUBS 5.83386f
C195 VDD2.n0 VSUBS 0.032592f
C196 VDD2.n1 VSUBS 0.029099f
C197 VDD2.n2 VSUBS 0.015637f
C198 VDD2.n3 VSUBS 0.036959f
C199 VDD2.n4 VSUBS 0.016556f
C200 VDD2.n5 VSUBS 0.029099f
C201 VDD2.n6 VSUBS 0.015637f
C202 VDD2.n7 VSUBS 0.036959f
C203 VDD2.n8 VSUBS 0.016556f
C204 VDD2.n9 VSUBS 0.029099f
C205 VDD2.n10 VSUBS 0.015637f
C206 VDD2.n11 VSUBS 0.036959f
C207 VDD2.n12 VSUBS 0.016556f
C208 VDD2.n13 VSUBS 0.029099f
C209 VDD2.n14 VSUBS 0.015637f
C210 VDD2.n15 VSUBS 0.036959f
C211 VDD2.n16 VSUBS 0.016556f
C212 VDD2.n17 VSUBS 0.029099f
C213 VDD2.n18 VSUBS 0.015637f
C214 VDD2.n19 VSUBS 0.036959f
C215 VDD2.n20 VSUBS 0.016556f
C216 VDD2.n21 VSUBS 0.029099f
C217 VDD2.n22 VSUBS 0.015637f
C218 VDD2.n23 VSUBS 0.036959f
C219 VDD2.n24 VSUBS 0.016556f
C220 VDD2.n25 VSUBS 0.267326f
C221 VDD2.t1 VSUBS 0.079925f
C222 VDD2.n26 VSUBS 0.027719f
C223 VDD2.n27 VSUBS 0.027803f
C224 VDD2.n28 VSUBS 0.015637f
C225 VDD2.n29 VSUBS 1.79949f
C226 VDD2.n30 VSUBS 0.029099f
C227 VDD2.n31 VSUBS 0.015637f
C228 VDD2.n32 VSUBS 0.016556f
C229 VDD2.n33 VSUBS 0.036959f
C230 VDD2.n34 VSUBS 0.036959f
C231 VDD2.n35 VSUBS 0.016556f
C232 VDD2.n36 VSUBS 0.015637f
C233 VDD2.n37 VSUBS 0.029099f
C234 VDD2.n38 VSUBS 0.029099f
C235 VDD2.n39 VSUBS 0.015637f
C236 VDD2.n40 VSUBS 0.016556f
C237 VDD2.n41 VSUBS 0.036959f
C238 VDD2.n42 VSUBS 0.036959f
C239 VDD2.n43 VSUBS 0.036959f
C240 VDD2.n44 VSUBS 0.016556f
C241 VDD2.n45 VSUBS 0.015637f
C242 VDD2.n46 VSUBS 0.029099f
C243 VDD2.n47 VSUBS 0.029099f
C244 VDD2.n48 VSUBS 0.015637f
C245 VDD2.n49 VSUBS 0.016096f
C246 VDD2.n50 VSUBS 0.016096f
C247 VDD2.n51 VSUBS 0.036959f
C248 VDD2.n52 VSUBS 0.036959f
C249 VDD2.n53 VSUBS 0.016556f
C250 VDD2.n54 VSUBS 0.015637f
C251 VDD2.n55 VSUBS 0.029099f
C252 VDD2.n56 VSUBS 0.029099f
C253 VDD2.n57 VSUBS 0.015637f
C254 VDD2.n58 VSUBS 0.016556f
C255 VDD2.n59 VSUBS 0.036959f
C256 VDD2.n60 VSUBS 0.036959f
C257 VDD2.n61 VSUBS 0.016556f
C258 VDD2.n62 VSUBS 0.015637f
C259 VDD2.n63 VSUBS 0.029099f
C260 VDD2.n64 VSUBS 0.029099f
C261 VDD2.n65 VSUBS 0.015637f
C262 VDD2.n66 VSUBS 0.016556f
C263 VDD2.n67 VSUBS 0.036959f
C264 VDD2.n68 VSUBS 0.036959f
C265 VDD2.n69 VSUBS 0.016556f
C266 VDD2.n70 VSUBS 0.015637f
C267 VDD2.n71 VSUBS 0.029099f
C268 VDD2.n72 VSUBS 0.029099f
C269 VDD2.n73 VSUBS 0.015637f
C270 VDD2.n74 VSUBS 0.016556f
C271 VDD2.n75 VSUBS 0.036959f
C272 VDD2.n76 VSUBS 0.091581f
C273 VDD2.n77 VSUBS 0.016556f
C274 VDD2.n78 VSUBS 0.015637f
C275 VDD2.n79 VSUBS 0.063286f
C276 VDD2.n80 VSUBS 1.05579f
C277 VDD2.n81 VSUBS 0.032592f
C278 VDD2.n82 VSUBS 0.029099f
C279 VDD2.n83 VSUBS 0.015637f
C280 VDD2.n84 VSUBS 0.036959f
C281 VDD2.n85 VSUBS 0.016556f
C282 VDD2.n86 VSUBS 0.029099f
C283 VDD2.n87 VSUBS 0.015637f
C284 VDD2.n88 VSUBS 0.036959f
C285 VDD2.n89 VSUBS 0.016556f
C286 VDD2.n90 VSUBS 0.029099f
C287 VDD2.n91 VSUBS 0.015637f
C288 VDD2.n92 VSUBS 0.036959f
C289 VDD2.n93 VSUBS 0.016556f
C290 VDD2.n94 VSUBS 0.029099f
C291 VDD2.n95 VSUBS 0.015637f
C292 VDD2.n96 VSUBS 0.036959f
C293 VDD2.n97 VSUBS 0.016556f
C294 VDD2.n98 VSUBS 0.029099f
C295 VDD2.n99 VSUBS 0.015637f
C296 VDD2.n100 VSUBS 0.036959f
C297 VDD2.n101 VSUBS 0.036959f
C298 VDD2.n102 VSUBS 0.016556f
C299 VDD2.n103 VSUBS 0.029099f
C300 VDD2.n104 VSUBS 0.015637f
C301 VDD2.n105 VSUBS 0.036959f
C302 VDD2.n106 VSUBS 0.016556f
C303 VDD2.n107 VSUBS 0.267326f
C304 VDD2.t0 VSUBS 0.079925f
C305 VDD2.n108 VSUBS 0.027719f
C306 VDD2.n109 VSUBS 0.027803f
C307 VDD2.n110 VSUBS 0.015637f
C308 VDD2.n111 VSUBS 1.79949f
C309 VDD2.n112 VSUBS 0.029099f
C310 VDD2.n113 VSUBS 0.015637f
C311 VDD2.n114 VSUBS 0.016556f
C312 VDD2.n115 VSUBS 0.036959f
C313 VDD2.n116 VSUBS 0.036959f
C314 VDD2.n117 VSUBS 0.016556f
C315 VDD2.n118 VSUBS 0.015637f
C316 VDD2.n119 VSUBS 0.029099f
C317 VDD2.n120 VSUBS 0.029099f
C318 VDD2.n121 VSUBS 0.015637f
C319 VDD2.n122 VSUBS 0.016556f
C320 VDD2.n123 VSUBS 0.036959f
C321 VDD2.n124 VSUBS 0.036959f
C322 VDD2.n125 VSUBS 0.016556f
C323 VDD2.n126 VSUBS 0.015637f
C324 VDD2.n127 VSUBS 0.029099f
C325 VDD2.n128 VSUBS 0.029099f
C326 VDD2.n129 VSUBS 0.015637f
C327 VDD2.n130 VSUBS 0.016096f
C328 VDD2.n131 VSUBS 0.016096f
C329 VDD2.n132 VSUBS 0.036959f
C330 VDD2.n133 VSUBS 0.036959f
C331 VDD2.n134 VSUBS 0.016556f
C332 VDD2.n135 VSUBS 0.015637f
C333 VDD2.n136 VSUBS 0.029099f
C334 VDD2.n137 VSUBS 0.029099f
C335 VDD2.n138 VSUBS 0.015637f
C336 VDD2.n139 VSUBS 0.016556f
C337 VDD2.n140 VSUBS 0.036959f
C338 VDD2.n141 VSUBS 0.036959f
C339 VDD2.n142 VSUBS 0.016556f
C340 VDD2.n143 VSUBS 0.015637f
C341 VDD2.n144 VSUBS 0.029099f
C342 VDD2.n145 VSUBS 0.029099f
C343 VDD2.n146 VSUBS 0.015637f
C344 VDD2.n147 VSUBS 0.016556f
C345 VDD2.n148 VSUBS 0.036959f
C346 VDD2.n149 VSUBS 0.036959f
C347 VDD2.n150 VSUBS 0.016556f
C348 VDD2.n151 VSUBS 0.015637f
C349 VDD2.n152 VSUBS 0.029099f
C350 VDD2.n153 VSUBS 0.029099f
C351 VDD2.n154 VSUBS 0.015637f
C352 VDD2.n155 VSUBS 0.016556f
C353 VDD2.n156 VSUBS 0.036959f
C354 VDD2.n157 VSUBS 0.091581f
C355 VDD2.n158 VSUBS 0.016556f
C356 VDD2.n159 VSUBS 0.015637f
C357 VDD2.n160 VSUBS 0.063286f
C358 VDD2.n161 VSUBS 0.066149f
C359 VDD2.n162 VSUBS 4.0309f
C360 VTAIL.n0 VSUBS 0.03267f
C361 VTAIL.n1 VSUBS 0.029168f
C362 VTAIL.n2 VSUBS 0.015674f
C363 VTAIL.n3 VSUBS 0.037047f
C364 VTAIL.n4 VSUBS 0.016596f
C365 VTAIL.n5 VSUBS 0.029168f
C366 VTAIL.n6 VSUBS 0.015674f
C367 VTAIL.n7 VSUBS 0.037047f
C368 VTAIL.n8 VSUBS 0.016596f
C369 VTAIL.n9 VSUBS 0.029168f
C370 VTAIL.n10 VSUBS 0.015674f
C371 VTAIL.n11 VSUBS 0.037047f
C372 VTAIL.n12 VSUBS 0.016596f
C373 VTAIL.n13 VSUBS 0.029168f
C374 VTAIL.n14 VSUBS 0.015674f
C375 VTAIL.n15 VSUBS 0.037047f
C376 VTAIL.n16 VSUBS 0.016596f
C377 VTAIL.n17 VSUBS 0.029168f
C378 VTAIL.n18 VSUBS 0.015674f
C379 VTAIL.n19 VSUBS 0.037047f
C380 VTAIL.n20 VSUBS 0.016596f
C381 VTAIL.n21 VSUBS 0.029168f
C382 VTAIL.n22 VSUBS 0.015674f
C383 VTAIL.n23 VSUBS 0.037047f
C384 VTAIL.n24 VSUBS 0.016596f
C385 VTAIL.n25 VSUBS 0.267963f
C386 VTAIL.t1 VSUBS 0.080115f
C387 VTAIL.n26 VSUBS 0.027786f
C388 VTAIL.n27 VSUBS 0.027869f
C389 VTAIL.n28 VSUBS 0.015674f
C390 VTAIL.n29 VSUBS 1.80378f
C391 VTAIL.n30 VSUBS 0.029168f
C392 VTAIL.n31 VSUBS 0.015674f
C393 VTAIL.n32 VSUBS 0.016596f
C394 VTAIL.n33 VSUBS 0.037047f
C395 VTAIL.n34 VSUBS 0.037047f
C396 VTAIL.n35 VSUBS 0.016596f
C397 VTAIL.n36 VSUBS 0.015674f
C398 VTAIL.n37 VSUBS 0.029168f
C399 VTAIL.n38 VSUBS 0.029168f
C400 VTAIL.n39 VSUBS 0.015674f
C401 VTAIL.n40 VSUBS 0.016596f
C402 VTAIL.n41 VSUBS 0.037047f
C403 VTAIL.n42 VSUBS 0.037047f
C404 VTAIL.n43 VSUBS 0.037047f
C405 VTAIL.n44 VSUBS 0.016596f
C406 VTAIL.n45 VSUBS 0.015674f
C407 VTAIL.n46 VSUBS 0.029168f
C408 VTAIL.n47 VSUBS 0.029168f
C409 VTAIL.n48 VSUBS 0.015674f
C410 VTAIL.n49 VSUBS 0.016135f
C411 VTAIL.n50 VSUBS 0.016135f
C412 VTAIL.n51 VSUBS 0.037047f
C413 VTAIL.n52 VSUBS 0.037047f
C414 VTAIL.n53 VSUBS 0.016596f
C415 VTAIL.n54 VSUBS 0.015674f
C416 VTAIL.n55 VSUBS 0.029168f
C417 VTAIL.n56 VSUBS 0.029168f
C418 VTAIL.n57 VSUBS 0.015674f
C419 VTAIL.n58 VSUBS 0.016596f
C420 VTAIL.n59 VSUBS 0.037047f
C421 VTAIL.n60 VSUBS 0.037047f
C422 VTAIL.n61 VSUBS 0.016596f
C423 VTAIL.n62 VSUBS 0.015674f
C424 VTAIL.n63 VSUBS 0.029168f
C425 VTAIL.n64 VSUBS 0.029168f
C426 VTAIL.n65 VSUBS 0.015674f
C427 VTAIL.n66 VSUBS 0.016596f
C428 VTAIL.n67 VSUBS 0.037047f
C429 VTAIL.n68 VSUBS 0.037047f
C430 VTAIL.n69 VSUBS 0.016596f
C431 VTAIL.n70 VSUBS 0.015674f
C432 VTAIL.n71 VSUBS 0.029168f
C433 VTAIL.n72 VSUBS 0.029168f
C434 VTAIL.n73 VSUBS 0.015674f
C435 VTAIL.n74 VSUBS 0.016596f
C436 VTAIL.n75 VSUBS 0.037047f
C437 VTAIL.n76 VSUBS 0.091799f
C438 VTAIL.n77 VSUBS 0.016596f
C439 VTAIL.n78 VSUBS 0.015674f
C440 VTAIL.n79 VSUBS 0.063437f
C441 VTAIL.n80 VSUBS 0.046133f
C442 VTAIL.n81 VSUBS 2.33752f
C443 VTAIL.n82 VSUBS 0.03267f
C444 VTAIL.n83 VSUBS 0.029168f
C445 VTAIL.n84 VSUBS 0.015674f
C446 VTAIL.n85 VSUBS 0.037047f
C447 VTAIL.n86 VSUBS 0.016596f
C448 VTAIL.n87 VSUBS 0.029168f
C449 VTAIL.n88 VSUBS 0.015674f
C450 VTAIL.n89 VSUBS 0.037047f
C451 VTAIL.n90 VSUBS 0.016596f
C452 VTAIL.n91 VSUBS 0.029168f
C453 VTAIL.n92 VSUBS 0.015674f
C454 VTAIL.n93 VSUBS 0.037047f
C455 VTAIL.n94 VSUBS 0.016596f
C456 VTAIL.n95 VSUBS 0.029168f
C457 VTAIL.n96 VSUBS 0.015674f
C458 VTAIL.n97 VSUBS 0.037047f
C459 VTAIL.n98 VSUBS 0.016596f
C460 VTAIL.n99 VSUBS 0.029168f
C461 VTAIL.n100 VSUBS 0.015674f
C462 VTAIL.n101 VSUBS 0.037047f
C463 VTAIL.n102 VSUBS 0.037047f
C464 VTAIL.n103 VSUBS 0.016596f
C465 VTAIL.n104 VSUBS 0.029168f
C466 VTAIL.n105 VSUBS 0.015674f
C467 VTAIL.n106 VSUBS 0.037047f
C468 VTAIL.n107 VSUBS 0.016596f
C469 VTAIL.n108 VSUBS 0.267963f
C470 VTAIL.t2 VSUBS 0.080115f
C471 VTAIL.n109 VSUBS 0.027786f
C472 VTAIL.n110 VSUBS 0.027869f
C473 VTAIL.n111 VSUBS 0.015674f
C474 VTAIL.n112 VSUBS 1.80378f
C475 VTAIL.n113 VSUBS 0.029168f
C476 VTAIL.n114 VSUBS 0.015674f
C477 VTAIL.n115 VSUBS 0.016596f
C478 VTAIL.n116 VSUBS 0.037047f
C479 VTAIL.n117 VSUBS 0.037047f
C480 VTAIL.n118 VSUBS 0.016596f
C481 VTAIL.n119 VSUBS 0.015674f
C482 VTAIL.n120 VSUBS 0.029168f
C483 VTAIL.n121 VSUBS 0.029168f
C484 VTAIL.n122 VSUBS 0.015674f
C485 VTAIL.n123 VSUBS 0.016596f
C486 VTAIL.n124 VSUBS 0.037047f
C487 VTAIL.n125 VSUBS 0.037047f
C488 VTAIL.n126 VSUBS 0.016596f
C489 VTAIL.n127 VSUBS 0.015674f
C490 VTAIL.n128 VSUBS 0.029168f
C491 VTAIL.n129 VSUBS 0.029168f
C492 VTAIL.n130 VSUBS 0.015674f
C493 VTAIL.n131 VSUBS 0.016135f
C494 VTAIL.n132 VSUBS 0.016135f
C495 VTAIL.n133 VSUBS 0.037047f
C496 VTAIL.n134 VSUBS 0.037047f
C497 VTAIL.n135 VSUBS 0.016596f
C498 VTAIL.n136 VSUBS 0.015674f
C499 VTAIL.n137 VSUBS 0.029168f
C500 VTAIL.n138 VSUBS 0.029168f
C501 VTAIL.n139 VSUBS 0.015674f
C502 VTAIL.n140 VSUBS 0.016596f
C503 VTAIL.n141 VSUBS 0.037047f
C504 VTAIL.n142 VSUBS 0.037047f
C505 VTAIL.n143 VSUBS 0.016596f
C506 VTAIL.n144 VSUBS 0.015674f
C507 VTAIL.n145 VSUBS 0.029168f
C508 VTAIL.n146 VSUBS 0.029168f
C509 VTAIL.n147 VSUBS 0.015674f
C510 VTAIL.n148 VSUBS 0.016596f
C511 VTAIL.n149 VSUBS 0.037047f
C512 VTAIL.n150 VSUBS 0.037047f
C513 VTAIL.n151 VSUBS 0.016596f
C514 VTAIL.n152 VSUBS 0.015674f
C515 VTAIL.n153 VSUBS 0.029168f
C516 VTAIL.n154 VSUBS 0.029168f
C517 VTAIL.n155 VSUBS 0.015674f
C518 VTAIL.n156 VSUBS 0.016596f
C519 VTAIL.n157 VSUBS 0.037047f
C520 VTAIL.n158 VSUBS 0.091799f
C521 VTAIL.n159 VSUBS 0.016596f
C522 VTAIL.n160 VSUBS 0.015674f
C523 VTAIL.n161 VSUBS 0.063437f
C524 VTAIL.n162 VSUBS 0.046133f
C525 VTAIL.n163 VSUBS 2.40558f
C526 VTAIL.n164 VSUBS 0.03267f
C527 VTAIL.n165 VSUBS 0.029168f
C528 VTAIL.n166 VSUBS 0.015674f
C529 VTAIL.n167 VSUBS 0.037047f
C530 VTAIL.n168 VSUBS 0.016596f
C531 VTAIL.n169 VSUBS 0.029168f
C532 VTAIL.n170 VSUBS 0.015674f
C533 VTAIL.n171 VSUBS 0.037047f
C534 VTAIL.n172 VSUBS 0.016596f
C535 VTAIL.n173 VSUBS 0.029168f
C536 VTAIL.n174 VSUBS 0.015674f
C537 VTAIL.n175 VSUBS 0.037047f
C538 VTAIL.n176 VSUBS 0.016596f
C539 VTAIL.n177 VSUBS 0.029168f
C540 VTAIL.n178 VSUBS 0.015674f
C541 VTAIL.n179 VSUBS 0.037047f
C542 VTAIL.n180 VSUBS 0.016596f
C543 VTAIL.n181 VSUBS 0.029168f
C544 VTAIL.n182 VSUBS 0.015674f
C545 VTAIL.n183 VSUBS 0.037047f
C546 VTAIL.n184 VSUBS 0.037047f
C547 VTAIL.n185 VSUBS 0.016596f
C548 VTAIL.n186 VSUBS 0.029168f
C549 VTAIL.n187 VSUBS 0.015674f
C550 VTAIL.n188 VSUBS 0.037047f
C551 VTAIL.n189 VSUBS 0.016596f
C552 VTAIL.n190 VSUBS 0.267963f
C553 VTAIL.t0 VSUBS 0.080115f
C554 VTAIL.n191 VSUBS 0.027786f
C555 VTAIL.n192 VSUBS 0.027869f
C556 VTAIL.n193 VSUBS 0.015674f
C557 VTAIL.n194 VSUBS 1.80378f
C558 VTAIL.n195 VSUBS 0.029168f
C559 VTAIL.n196 VSUBS 0.015674f
C560 VTAIL.n197 VSUBS 0.016596f
C561 VTAIL.n198 VSUBS 0.037047f
C562 VTAIL.n199 VSUBS 0.037047f
C563 VTAIL.n200 VSUBS 0.016596f
C564 VTAIL.n201 VSUBS 0.015674f
C565 VTAIL.n202 VSUBS 0.029168f
C566 VTAIL.n203 VSUBS 0.029168f
C567 VTAIL.n204 VSUBS 0.015674f
C568 VTAIL.n205 VSUBS 0.016596f
C569 VTAIL.n206 VSUBS 0.037047f
C570 VTAIL.n207 VSUBS 0.037047f
C571 VTAIL.n208 VSUBS 0.016596f
C572 VTAIL.n209 VSUBS 0.015674f
C573 VTAIL.n210 VSUBS 0.029168f
C574 VTAIL.n211 VSUBS 0.029168f
C575 VTAIL.n212 VSUBS 0.015674f
C576 VTAIL.n213 VSUBS 0.016135f
C577 VTAIL.n214 VSUBS 0.016135f
C578 VTAIL.n215 VSUBS 0.037047f
C579 VTAIL.n216 VSUBS 0.037047f
C580 VTAIL.n217 VSUBS 0.016596f
C581 VTAIL.n218 VSUBS 0.015674f
C582 VTAIL.n219 VSUBS 0.029168f
C583 VTAIL.n220 VSUBS 0.029168f
C584 VTAIL.n221 VSUBS 0.015674f
C585 VTAIL.n222 VSUBS 0.016596f
C586 VTAIL.n223 VSUBS 0.037047f
C587 VTAIL.n224 VSUBS 0.037047f
C588 VTAIL.n225 VSUBS 0.016596f
C589 VTAIL.n226 VSUBS 0.015674f
C590 VTAIL.n227 VSUBS 0.029168f
C591 VTAIL.n228 VSUBS 0.029168f
C592 VTAIL.n229 VSUBS 0.015674f
C593 VTAIL.n230 VSUBS 0.016596f
C594 VTAIL.n231 VSUBS 0.037047f
C595 VTAIL.n232 VSUBS 0.037047f
C596 VTAIL.n233 VSUBS 0.016596f
C597 VTAIL.n234 VSUBS 0.015674f
C598 VTAIL.n235 VSUBS 0.029168f
C599 VTAIL.n236 VSUBS 0.029168f
C600 VTAIL.n237 VSUBS 0.015674f
C601 VTAIL.n238 VSUBS 0.016596f
C602 VTAIL.n239 VSUBS 0.037047f
C603 VTAIL.n240 VSUBS 0.091799f
C604 VTAIL.n241 VSUBS 0.016596f
C605 VTAIL.n242 VSUBS 0.015674f
C606 VTAIL.n243 VSUBS 0.063437f
C607 VTAIL.n244 VSUBS 0.046133f
C608 VTAIL.n245 VSUBS 2.11147f
C609 VTAIL.n246 VSUBS 0.03267f
C610 VTAIL.n247 VSUBS 0.029168f
C611 VTAIL.n248 VSUBS 0.015674f
C612 VTAIL.n249 VSUBS 0.037047f
C613 VTAIL.n250 VSUBS 0.016596f
C614 VTAIL.n251 VSUBS 0.029168f
C615 VTAIL.n252 VSUBS 0.015674f
C616 VTAIL.n253 VSUBS 0.037047f
C617 VTAIL.n254 VSUBS 0.016596f
C618 VTAIL.n255 VSUBS 0.029168f
C619 VTAIL.n256 VSUBS 0.015674f
C620 VTAIL.n257 VSUBS 0.037047f
C621 VTAIL.n258 VSUBS 0.016596f
C622 VTAIL.n259 VSUBS 0.029168f
C623 VTAIL.n260 VSUBS 0.015674f
C624 VTAIL.n261 VSUBS 0.037047f
C625 VTAIL.n262 VSUBS 0.016596f
C626 VTAIL.n263 VSUBS 0.029168f
C627 VTAIL.n264 VSUBS 0.015674f
C628 VTAIL.n265 VSUBS 0.037047f
C629 VTAIL.n266 VSUBS 0.016596f
C630 VTAIL.n267 VSUBS 0.029168f
C631 VTAIL.n268 VSUBS 0.015674f
C632 VTAIL.n269 VSUBS 0.037047f
C633 VTAIL.n270 VSUBS 0.016596f
C634 VTAIL.n271 VSUBS 0.267963f
C635 VTAIL.t3 VSUBS 0.080115f
C636 VTAIL.n272 VSUBS 0.027786f
C637 VTAIL.n273 VSUBS 0.027869f
C638 VTAIL.n274 VSUBS 0.015674f
C639 VTAIL.n275 VSUBS 1.80378f
C640 VTAIL.n276 VSUBS 0.029168f
C641 VTAIL.n277 VSUBS 0.015674f
C642 VTAIL.n278 VSUBS 0.016596f
C643 VTAIL.n279 VSUBS 0.037047f
C644 VTAIL.n280 VSUBS 0.037047f
C645 VTAIL.n281 VSUBS 0.016596f
C646 VTAIL.n282 VSUBS 0.015674f
C647 VTAIL.n283 VSUBS 0.029168f
C648 VTAIL.n284 VSUBS 0.029168f
C649 VTAIL.n285 VSUBS 0.015674f
C650 VTAIL.n286 VSUBS 0.016596f
C651 VTAIL.n287 VSUBS 0.037047f
C652 VTAIL.n288 VSUBS 0.037047f
C653 VTAIL.n289 VSUBS 0.037047f
C654 VTAIL.n290 VSUBS 0.016596f
C655 VTAIL.n291 VSUBS 0.015674f
C656 VTAIL.n292 VSUBS 0.029168f
C657 VTAIL.n293 VSUBS 0.029168f
C658 VTAIL.n294 VSUBS 0.015674f
C659 VTAIL.n295 VSUBS 0.016135f
C660 VTAIL.n296 VSUBS 0.016135f
C661 VTAIL.n297 VSUBS 0.037047f
C662 VTAIL.n298 VSUBS 0.037047f
C663 VTAIL.n299 VSUBS 0.016596f
C664 VTAIL.n300 VSUBS 0.015674f
C665 VTAIL.n301 VSUBS 0.029168f
C666 VTAIL.n302 VSUBS 0.029168f
C667 VTAIL.n303 VSUBS 0.015674f
C668 VTAIL.n304 VSUBS 0.016596f
C669 VTAIL.n305 VSUBS 0.037047f
C670 VTAIL.n306 VSUBS 0.037047f
C671 VTAIL.n307 VSUBS 0.016596f
C672 VTAIL.n308 VSUBS 0.015674f
C673 VTAIL.n309 VSUBS 0.029168f
C674 VTAIL.n310 VSUBS 0.029168f
C675 VTAIL.n311 VSUBS 0.015674f
C676 VTAIL.n312 VSUBS 0.016596f
C677 VTAIL.n313 VSUBS 0.037047f
C678 VTAIL.n314 VSUBS 0.037047f
C679 VTAIL.n315 VSUBS 0.016596f
C680 VTAIL.n316 VSUBS 0.015674f
C681 VTAIL.n317 VSUBS 0.029168f
C682 VTAIL.n318 VSUBS 0.029168f
C683 VTAIL.n319 VSUBS 0.015674f
C684 VTAIL.n320 VSUBS 0.016596f
C685 VTAIL.n321 VSUBS 0.037047f
C686 VTAIL.n322 VSUBS 0.091799f
C687 VTAIL.n323 VSUBS 0.016596f
C688 VTAIL.n324 VSUBS 0.015674f
C689 VTAIL.n325 VSUBS 0.063437f
C690 VTAIL.n326 VSUBS 0.046133f
C691 VTAIL.n327 VSUBS 1.98831f
C692 VN.t0 VSUBS 4.89627f
C693 VN.t1 VSUBS 5.70271f
C694 B.n0 VSUBS 0.006047f
C695 B.n1 VSUBS 0.006047f
C696 B.n2 VSUBS 0.008943f
C697 B.n3 VSUBS 0.006853f
C698 B.n4 VSUBS 0.006853f
C699 B.n5 VSUBS 0.006853f
C700 B.n6 VSUBS 0.006853f
C701 B.n7 VSUBS 0.006853f
C702 B.n8 VSUBS 0.006853f
C703 B.n9 VSUBS 0.006853f
C704 B.n10 VSUBS 0.006853f
C705 B.n11 VSUBS 0.006853f
C706 B.n12 VSUBS 0.006853f
C707 B.n13 VSUBS 0.006853f
C708 B.n14 VSUBS 0.006853f
C709 B.n15 VSUBS 0.006853f
C710 B.n16 VSUBS 0.015199f
C711 B.n17 VSUBS 0.006853f
C712 B.n18 VSUBS 0.006853f
C713 B.n19 VSUBS 0.006853f
C714 B.n20 VSUBS 0.006853f
C715 B.n21 VSUBS 0.006853f
C716 B.n22 VSUBS 0.006853f
C717 B.n23 VSUBS 0.006853f
C718 B.n24 VSUBS 0.006853f
C719 B.n25 VSUBS 0.006853f
C720 B.n26 VSUBS 0.006853f
C721 B.n27 VSUBS 0.006853f
C722 B.n28 VSUBS 0.006853f
C723 B.n29 VSUBS 0.006853f
C724 B.n30 VSUBS 0.006853f
C725 B.n31 VSUBS 0.006853f
C726 B.n32 VSUBS 0.006853f
C727 B.n33 VSUBS 0.006853f
C728 B.n34 VSUBS 0.006853f
C729 B.n35 VSUBS 0.006853f
C730 B.n36 VSUBS 0.006853f
C731 B.n37 VSUBS 0.006853f
C732 B.n38 VSUBS 0.006853f
C733 B.n39 VSUBS 0.006853f
C734 B.n40 VSUBS 0.006853f
C735 B.n41 VSUBS 0.006853f
C736 B.t1 VSUBS 0.271617f
C737 B.t2 VSUBS 0.310774f
C738 B.t0 VSUBS 2.19837f
C739 B.n42 VSUBS 0.491667f
C740 B.n43 VSUBS 0.286995f
C741 B.n44 VSUBS 0.006853f
C742 B.n45 VSUBS 0.006853f
C743 B.n46 VSUBS 0.006853f
C744 B.n47 VSUBS 0.006853f
C745 B.n48 VSUBS 0.00383f
C746 B.n49 VSUBS 0.006853f
C747 B.t4 VSUBS 0.27162f
C748 B.t5 VSUBS 0.310777f
C749 B.t3 VSUBS 2.19837f
C750 B.n50 VSUBS 0.491665f
C751 B.n51 VSUBS 0.286992f
C752 B.n52 VSUBS 0.015877f
C753 B.n53 VSUBS 0.006853f
C754 B.n54 VSUBS 0.006853f
C755 B.n55 VSUBS 0.006853f
C756 B.n56 VSUBS 0.006853f
C757 B.n57 VSUBS 0.006853f
C758 B.n58 VSUBS 0.006853f
C759 B.n59 VSUBS 0.006853f
C760 B.n60 VSUBS 0.006853f
C761 B.n61 VSUBS 0.006853f
C762 B.n62 VSUBS 0.006853f
C763 B.n63 VSUBS 0.006853f
C764 B.n64 VSUBS 0.006853f
C765 B.n65 VSUBS 0.006853f
C766 B.n66 VSUBS 0.006853f
C767 B.n67 VSUBS 0.006853f
C768 B.n68 VSUBS 0.006853f
C769 B.n69 VSUBS 0.006853f
C770 B.n70 VSUBS 0.006853f
C771 B.n71 VSUBS 0.006853f
C772 B.n72 VSUBS 0.006853f
C773 B.n73 VSUBS 0.006853f
C774 B.n74 VSUBS 0.006853f
C775 B.n75 VSUBS 0.006853f
C776 B.n76 VSUBS 0.016042f
C777 B.n77 VSUBS 0.006853f
C778 B.n78 VSUBS 0.006853f
C779 B.n79 VSUBS 0.006853f
C780 B.n80 VSUBS 0.006853f
C781 B.n81 VSUBS 0.006853f
C782 B.n82 VSUBS 0.006853f
C783 B.n83 VSUBS 0.006853f
C784 B.n84 VSUBS 0.006853f
C785 B.n85 VSUBS 0.006853f
C786 B.n86 VSUBS 0.006853f
C787 B.n87 VSUBS 0.006853f
C788 B.n88 VSUBS 0.006853f
C789 B.n89 VSUBS 0.006853f
C790 B.n90 VSUBS 0.006853f
C791 B.n91 VSUBS 0.006853f
C792 B.n92 VSUBS 0.006853f
C793 B.n93 VSUBS 0.006853f
C794 B.n94 VSUBS 0.006853f
C795 B.n95 VSUBS 0.006853f
C796 B.n96 VSUBS 0.006853f
C797 B.n97 VSUBS 0.006853f
C798 B.n98 VSUBS 0.006853f
C799 B.n99 VSUBS 0.006853f
C800 B.n100 VSUBS 0.006853f
C801 B.n101 VSUBS 0.006853f
C802 B.n102 VSUBS 0.006853f
C803 B.n103 VSUBS 0.006853f
C804 B.n104 VSUBS 0.006853f
C805 B.n105 VSUBS 0.006853f
C806 B.n106 VSUBS 0.015199f
C807 B.n107 VSUBS 0.006853f
C808 B.n108 VSUBS 0.006853f
C809 B.n109 VSUBS 0.006853f
C810 B.n110 VSUBS 0.006853f
C811 B.n111 VSUBS 0.006853f
C812 B.n112 VSUBS 0.006853f
C813 B.n113 VSUBS 0.006853f
C814 B.n114 VSUBS 0.006853f
C815 B.n115 VSUBS 0.006853f
C816 B.n116 VSUBS 0.006853f
C817 B.n117 VSUBS 0.006853f
C818 B.n118 VSUBS 0.006853f
C819 B.n119 VSUBS 0.006853f
C820 B.n120 VSUBS 0.006853f
C821 B.n121 VSUBS 0.006853f
C822 B.n122 VSUBS 0.006853f
C823 B.n123 VSUBS 0.006853f
C824 B.n124 VSUBS 0.006853f
C825 B.n125 VSUBS 0.006853f
C826 B.n126 VSUBS 0.006853f
C827 B.n127 VSUBS 0.006853f
C828 B.n128 VSUBS 0.006853f
C829 B.n129 VSUBS 0.006853f
C830 B.n130 VSUBS 0.006853f
C831 B.n131 VSUBS 0.00645f
C832 B.n132 VSUBS 0.006853f
C833 B.n133 VSUBS 0.006853f
C834 B.n134 VSUBS 0.006853f
C835 B.n135 VSUBS 0.006853f
C836 B.n136 VSUBS 0.006853f
C837 B.t8 VSUBS 0.271617f
C838 B.t7 VSUBS 0.310774f
C839 B.t6 VSUBS 2.19837f
C840 B.n137 VSUBS 0.491667f
C841 B.n138 VSUBS 0.286995f
C842 B.n139 VSUBS 0.006853f
C843 B.n140 VSUBS 0.006853f
C844 B.n141 VSUBS 0.006853f
C845 B.n142 VSUBS 0.006853f
C846 B.n143 VSUBS 0.006853f
C847 B.n144 VSUBS 0.006853f
C848 B.n145 VSUBS 0.006853f
C849 B.n146 VSUBS 0.006853f
C850 B.n147 VSUBS 0.006853f
C851 B.n148 VSUBS 0.006853f
C852 B.n149 VSUBS 0.006853f
C853 B.n150 VSUBS 0.006853f
C854 B.n151 VSUBS 0.006853f
C855 B.n152 VSUBS 0.006853f
C856 B.n153 VSUBS 0.006853f
C857 B.n154 VSUBS 0.006853f
C858 B.n155 VSUBS 0.006853f
C859 B.n156 VSUBS 0.006853f
C860 B.n157 VSUBS 0.006853f
C861 B.n158 VSUBS 0.006853f
C862 B.n159 VSUBS 0.006853f
C863 B.n160 VSUBS 0.006853f
C864 B.n161 VSUBS 0.006853f
C865 B.n162 VSUBS 0.006853f
C866 B.n163 VSUBS 0.016042f
C867 B.n164 VSUBS 0.006853f
C868 B.n165 VSUBS 0.006853f
C869 B.n166 VSUBS 0.006853f
C870 B.n167 VSUBS 0.006853f
C871 B.n168 VSUBS 0.006853f
C872 B.n169 VSUBS 0.006853f
C873 B.n170 VSUBS 0.006853f
C874 B.n171 VSUBS 0.006853f
C875 B.n172 VSUBS 0.006853f
C876 B.n173 VSUBS 0.006853f
C877 B.n174 VSUBS 0.006853f
C878 B.n175 VSUBS 0.006853f
C879 B.n176 VSUBS 0.006853f
C880 B.n177 VSUBS 0.006853f
C881 B.n178 VSUBS 0.006853f
C882 B.n179 VSUBS 0.006853f
C883 B.n180 VSUBS 0.006853f
C884 B.n181 VSUBS 0.006853f
C885 B.n182 VSUBS 0.006853f
C886 B.n183 VSUBS 0.006853f
C887 B.n184 VSUBS 0.006853f
C888 B.n185 VSUBS 0.006853f
C889 B.n186 VSUBS 0.006853f
C890 B.n187 VSUBS 0.006853f
C891 B.n188 VSUBS 0.006853f
C892 B.n189 VSUBS 0.006853f
C893 B.n190 VSUBS 0.006853f
C894 B.n191 VSUBS 0.006853f
C895 B.n192 VSUBS 0.006853f
C896 B.n193 VSUBS 0.006853f
C897 B.n194 VSUBS 0.006853f
C898 B.n195 VSUBS 0.006853f
C899 B.n196 VSUBS 0.006853f
C900 B.n197 VSUBS 0.006853f
C901 B.n198 VSUBS 0.006853f
C902 B.n199 VSUBS 0.006853f
C903 B.n200 VSUBS 0.006853f
C904 B.n201 VSUBS 0.006853f
C905 B.n202 VSUBS 0.006853f
C906 B.n203 VSUBS 0.006853f
C907 B.n204 VSUBS 0.006853f
C908 B.n205 VSUBS 0.006853f
C909 B.n206 VSUBS 0.006853f
C910 B.n207 VSUBS 0.006853f
C911 B.n208 VSUBS 0.006853f
C912 B.n209 VSUBS 0.006853f
C913 B.n210 VSUBS 0.006853f
C914 B.n211 VSUBS 0.006853f
C915 B.n212 VSUBS 0.006853f
C916 B.n213 VSUBS 0.006853f
C917 B.n214 VSUBS 0.006853f
C918 B.n215 VSUBS 0.006853f
C919 B.n216 VSUBS 0.006853f
C920 B.n217 VSUBS 0.006853f
C921 B.n218 VSUBS 0.015199f
C922 B.n219 VSUBS 0.015199f
C923 B.n220 VSUBS 0.016042f
C924 B.n221 VSUBS 0.006853f
C925 B.n222 VSUBS 0.006853f
C926 B.n223 VSUBS 0.006853f
C927 B.n224 VSUBS 0.006853f
C928 B.n225 VSUBS 0.006853f
C929 B.n226 VSUBS 0.006853f
C930 B.n227 VSUBS 0.006853f
C931 B.n228 VSUBS 0.006853f
C932 B.n229 VSUBS 0.006853f
C933 B.n230 VSUBS 0.006853f
C934 B.n231 VSUBS 0.006853f
C935 B.n232 VSUBS 0.006853f
C936 B.n233 VSUBS 0.006853f
C937 B.n234 VSUBS 0.006853f
C938 B.n235 VSUBS 0.006853f
C939 B.n236 VSUBS 0.006853f
C940 B.n237 VSUBS 0.006853f
C941 B.n238 VSUBS 0.006853f
C942 B.n239 VSUBS 0.006853f
C943 B.n240 VSUBS 0.006853f
C944 B.n241 VSUBS 0.006853f
C945 B.n242 VSUBS 0.006853f
C946 B.n243 VSUBS 0.006853f
C947 B.n244 VSUBS 0.006853f
C948 B.n245 VSUBS 0.006853f
C949 B.n246 VSUBS 0.006853f
C950 B.n247 VSUBS 0.006853f
C951 B.n248 VSUBS 0.006853f
C952 B.n249 VSUBS 0.006853f
C953 B.n250 VSUBS 0.006853f
C954 B.n251 VSUBS 0.006853f
C955 B.n252 VSUBS 0.006853f
C956 B.n253 VSUBS 0.006853f
C957 B.n254 VSUBS 0.006853f
C958 B.n255 VSUBS 0.006853f
C959 B.n256 VSUBS 0.006853f
C960 B.n257 VSUBS 0.006853f
C961 B.n258 VSUBS 0.006853f
C962 B.n259 VSUBS 0.006853f
C963 B.n260 VSUBS 0.006853f
C964 B.n261 VSUBS 0.006853f
C965 B.n262 VSUBS 0.006853f
C966 B.n263 VSUBS 0.006853f
C967 B.n264 VSUBS 0.006853f
C968 B.n265 VSUBS 0.006853f
C969 B.n266 VSUBS 0.006853f
C970 B.n267 VSUBS 0.006853f
C971 B.n268 VSUBS 0.006853f
C972 B.n269 VSUBS 0.006853f
C973 B.n270 VSUBS 0.006853f
C974 B.n271 VSUBS 0.006853f
C975 B.n272 VSUBS 0.006853f
C976 B.n273 VSUBS 0.006853f
C977 B.n274 VSUBS 0.006853f
C978 B.n275 VSUBS 0.006853f
C979 B.n276 VSUBS 0.006853f
C980 B.n277 VSUBS 0.006853f
C981 B.n278 VSUBS 0.006853f
C982 B.n279 VSUBS 0.006853f
C983 B.n280 VSUBS 0.006853f
C984 B.n281 VSUBS 0.006853f
C985 B.n282 VSUBS 0.006853f
C986 B.n283 VSUBS 0.006853f
C987 B.n284 VSUBS 0.006853f
C988 B.n285 VSUBS 0.006853f
C989 B.n286 VSUBS 0.006853f
C990 B.n287 VSUBS 0.006853f
C991 B.n288 VSUBS 0.006853f
C992 B.n289 VSUBS 0.006853f
C993 B.n290 VSUBS 0.006853f
C994 B.n291 VSUBS 0.006853f
C995 B.n292 VSUBS 0.006853f
C996 B.n293 VSUBS 0.006853f
C997 B.n294 VSUBS 0.00645f
C998 B.n295 VSUBS 0.015877f
C999 B.n296 VSUBS 0.00383f
C1000 B.n297 VSUBS 0.006853f
C1001 B.n298 VSUBS 0.006853f
C1002 B.n299 VSUBS 0.006853f
C1003 B.n300 VSUBS 0.006853f
C1004 B.n301 VSUBS 0.006853f
C1005 B.n302 VSUBS 0.006853f
C1006 B.n303 VSUBS 0.006853f
C1007 B.n304 VSUBS 0.006853f
C1008 B.n305 VSUBS 0.006853f
C1009 B.n306 VSUBS 0.006853f
C1010 B.n307 VSUBS 0.006853f
C1011 B.n308 VSUBS 0.006853f
C1012 B.t11 VSUBS 0.27162f
C1013 B.t10 VSUBS 0.310777f
C1014 B.t9 VSUBS 2.19837f
C1015 B.n309 VSUBS 0.491665f
C1016 B.n310 VSUBS 0.286992f
C1017 B.n311 VSUBS 0.015877f
C1018 B.n312 VSUBS 0.00383f
C1019 B.n313 VSUBS 0.006853f
C1020 B.n314 VSUBS 0.006853f
C1021 B.n315 VSUBS 0.006853f
C1022 B.n316 VSUBS 0.006853f
C1023 B.n317 VSUBS 0.006853f
C1024 B.n318 VSUBS 0.006853f
C1025 B.n319 VSUBS 0.006853f
C1026 B.n320 VSUBS 0.006853f
C1027 B.n321 VSUBS 0.006853f
C1028 B.n322 VSUBS 0.006853f
C1029 B.n323 VSUBS 0.006853f
C1030 B.n324 VSUBS 0.006853f
C1031 B.n325 VSUBS 0.006853f
C1032 B.n326 VSUBS 0.006853f
C1033 B.n327 VSUBS 0.006853f
C1034 B.n328 VSUBS 0.006853f
C1035 B.n329 VSUBS 0.006853f
C1036 B.n330 VSUBS 0.006853f
C1037 B.n331 VSUBS 0.006853f
C1038 B.n332 VSUBS 0.006853f
C1039 B.n333 VSUBS 0.006853f
C1040 B.n334 VSUBS 0.006853f
C1041 B.n335 VSUBS 0.006853f
C1042 B.n336 VSUBS 0.006853f
C1043 B.n337 VSUBS 0.006853f
C1044 B.n338 VSUBS 0.006853f
C1045 B.n339 VSUBS 0.006853f
C1046 B.n340 VSUBS 0.006853f
C1047 B.n341 VSUBS 0.006853f
C1048 B.n342 VSUBS 0.006853f
C1049 B.n343 VSUBS 0.006853f
C1050 B.n344 VSUBS 0.006853f
C1051 B.n345 VSUBS 0.006853f
C1052 B.n346 VSUBS 0.006853f
C1053 B.n347 VSUBS 0.006853f
C1054 B.n348 VSUBS 0.006853f
C1055 B.n349 VSUBS 0.006853f
C1056 B.n350 VSUBS 0.006853f
C1057 B.n351 VSUBS 0.006853f
C1058 B.n352 VSUBS 0.006853f
C1059 B.n353 VSUBS 0.006853f
C1060 B.n354 VSUBS 0.006853f
C1061 B.n355 VSUBS 0.006853f
C1062 B.n356 VSUBS 0.006853f
C1063 B.n357 VSUBS 0.006853f
C1064 B.n358 VSUBS 0.006853f
C1065 B.n359 VSUBS 0.006853f
C1066 B.n360 VSUBS 0.006853f
C1067 B.n361 VSUBS 0.006853f
C1068 B.n362 VSUBS 0.006853f
C1069 B.n363 VSUBS 0.006853f
C1070 B.n364 VSUBS 0.006853f
C1071 B.n365 VSUBS 0.006853f
C1072 B.n366 VSUBS 0.006853f
C1073 B.n367 VSUBS 0.006853f
C1074 B.n368 VSUBS 0.006853f
C1075 B.n369 VSUBS 0.006853f
C1076 B.n370 VSUBS 0.006853f
C1077 B.n371 VSUBS 0.006853f
C1078 B.n372 VSUBS 0.006853f
C1079 B.n373 VSUBS 0.006853f
C1080 B.n374 VSUBS 0.006853f
C1081 B.n375 VSUBS 0.006853f
C1082 B.n376 VSUBS 0.006853f
C1083 B.n377 VSUBS 0.006853f
C1084 B.n378 VSUBS 0.006853f
C1085 B.n379 VSUBS 0.006853f
C1086 B.n380 VSUBS 0.006853f
C1087 B.n381 VSUBS 0.006853f
C1088 B.n382 VSUBS 0.006853f
C1089 B.n383 VSUBS 0.006853f
C1090 B.n384 VSUBS 0.006853f
C1091 B.n385 VSUBS 0.006853f
C1092 B.n386 VSUBS 0.006853f
C1093 B.n387 VSUBS 0.016042f
C1094 B.n388 VSUBS 0.015199f
C1095 B.n389 VSUBS 0.016042f
C1096 B.n390 VSUBS 0.006853f
C1097 B.n391 VSUBS 0.006853f
C1098 B.n392 VSUBS 0.006853f
C1099 B.n393 VSUBS 0.006853f
C1100 B.n394 VSUBS 0.006853f
C1101 B.n395 VSUBS 0.006853f
C1102 B.n396 VSUBS 0.006853f
C1103 B.n397 VSUBS 0.006853f
C1104 B.n398 VSUBS 0.006853f
C1105 B.n399 VSUBS 0.006853f
C1106 B.n400 VSUBS 0.006853f
C1107 B.n401 VSUBS 0.006853f
C1108 B.n402 VSUBS 0.006853f
C1109 B.n403 VSUBS 0.006853f
C1110 B.n404 VSUBS 0.006853f
C1111 B.n405 VSUBS 0.006853f
C1112 B.n406 VSUBS 0.006853f
C1113 B.n407 VSUBS 0.006853f
C1114 B.n408 VSUBS 0.006853f
C1115 B.n409 VSUBS 0.006853f
C1116 B.n410 VSUBS 0.006853f
C1117 B.n411 VSUBS 0.006853f
C1118 B.n412 VSUBS 0.006853f
C1119 B.n413 VSUBS 0.006853f
C1120 B.n414 VSUBS 0.006853f
C1121 B.n415 VSUBS 0.006853f
C1122 B.n416 VSUBS 0.006853f
C1123 B.n417 VSUBS 0.006853f
C1124 B.n418 VSUBS 0.006853f
C1125 B.n419 VSUBS 0.006853f
C1126 B.n420 VSUBS 0.006853f
C1127 B.n421 VSUBS 0.006853f
C1128 B.n422 VSUBS 0.006853f
C1129 B.n423 VSUBS 0.006853f
C1130 B.n424 VSUBS 0.006853f
C1131 B.n425 VSUBS 0.006853f
C1132 B.n426 VSUBS 0.006853f
C1133 B.n427 VSUBS 0.006853f
C1134 B.n428 VSUBS 0.006853f
C1135 B.n429 VSUBS 0.006853f
C1136 B.n430 VSUBS 0.006853f
C1137 B.n431 VSUBS 0.006853f
C1138 B.n432 VSUBS 0.006853f
C1139 B.n433 VSUBS 0.006853f
C1140 B.n434 VSUBS 0.006853f
C1141 B.n435 VSUBS 0.006853f
C1142 B.n436 VSUBS 0.006853f
C1143 B.n437 VSUBS 0.006853f
C1144 B.n438 VSUBS 0.006853f
C1145 B.n439 VSUBS 0.006853f
C1146 B.n440 VSUBS 0.006853f
C1147 B.n441 VSUBS 0.006853f
C1148 B.n442 VSUBS 0.006853f
C1149 B.n443 VSUBS 0.006853f
C1150 B.n444 VSUBS 0.006853f
C1151 B.n445 VSUBS 0.006853f
C1152 B.n446 VSUBS 0.006853f
C1153 B.n447 VSUBS 0.006853f
C1154 B.n448 VSUBS 0.006853f
C1155 B.n449 VSUBS 0.006853f
C1156 B.n450 VSUBS 0.006853f
C1157 B.n451 VSUBS 0.006853f
C1158 B.n452 VSUBS 0.006853f
C1159 B.n453 VSUBS 0.006853f
C1160 B.n454 VSUBS 0.006853f
C1161 B.n455 VSUBS 0.006853f
C1162 B.n456 VSUBS 0.006853f
C1163 B.n457 VSUBS 0.006853f
C1164 B.n458 VSUBS 0.006853f
C1165 B.n459 VSUBS 0.006853f
C1166 B.n460 VSUBS 0.006853f
C1167 B.n461 VSUBS 0.006853f
C1168 B.n462 VSUBS 0.006853f
C1169 B.n463 VSUBS 0.006853f
C1170 B.n464 VSUBS 0.006853f
C1171 B.n465 VSUBS 0.006853f
C1172 B.n466 VSUBS 0.006853f
C1173 B.n467 VSUBS 0.006853f
C1174 B.n468 VSUBS 0.006853f
C1175 B.n469 VSUBS 0.006853f
C1176 B.n470 VSUBS 0.006853f
C1177 B.n471 VSUBS 0.006853f
C1178 B.n472 VSUBS 0.006853f
C1179 B.n473 VSUBS 0.006853f
C1180 B.n474 VSUBS 0.006853f
C1181 B.n475 VSUBS 0.006853f
C1182 B.n476 VSUBS 0.006853f
C1183 B.n477 VSUBS 0.015199f
C1184 B.n478 VSUBS 0.015199f
C1185 B.n479 VSUBS 0.016042f
C1186 B.n480 VSUBS 0.006853f
C1187 B.n481 VSUBS 0.006853f
C1188 B.n482 VSUBS 0.006853f
C1189 B.n483 VSUBS 0.006853f
C1190 B.n484 VSUBS 0.006853f
C1191 B.n485 VSUBS 0.006853f
C1192 B.n486 VSUBS 0.006853f
C1193 B.n487 VSUBS 0.006853f
C1194 B.n488 VSUBS 0.006853f
C1195 B.n489 VSUBS 0.006853f
C1196 B.n490 VSUBS 0.006853f
C1197 B.n491 VSUBS 0.006853f
C1198 B.n492 VSUBS 0.006853f
C1199 B.n493 VSUBS 0.006853f
C1200 B.n494 VSUBS 0.006853f
C1201 B.n495 VSUBS 0.006853f
C1202 B.n496 VSUBS 0.006853f
C1203 B.n497 VSUBS 0.006853f
C1204 B.n498 VSUBS 0.006853f
C1205 B.n499 VSUBS 0.006853f
C1206 B.n500 VSUBS 0.006853f
C1207 B.n501 VSUBS 0.006853f
C1208 B.n502 VSUBS 0.006853f
C1209 B.n503 VSUBS 0.006853f
C1210 B.n504 VSUBS 0.006853f
C1211 B.n505 VSUBS 0.006853f
C1212 B.n506 VSUBS 0.006853f
C1213 B.n507 VSUBS 0.006853f
C1214 B.n508 VSUBS 0.006853f
C1215 B.n509 VSUBS 0.006853f
C1216 B.n510 VSUBS 0.006853f
C1217 B.n511 VSUBS 0.006853f
C1218 B.n512 VSUBS 0.006853f
C1219 B.n513 VSUBS 0.006853f
C1220 B.n514 VSUBS 0.006853f
C1221 B.n515 VSUBS 0.006853f
C1222 B.n516 VSUBS 0.006853f
C1223 B.n517 VSUBS 0.006853f
C1224 B.n518 VSUBS 0.006853f
C1225 B.n519 VSUBS 0.006853f
C1226 B.n520 VSUBS 0.006853f
C1227 B.n521 VSUBS 0.006853f
C1228 B.n522 VSUBS 0.006853f
C1229 B.n523 VSUBS 0.006853f
C1230 B.n524 VSUBS 0.006853f
C1231 B.n525 VSUBS 0.006853f
C1232 B.n526 VSUBS 0.006853f
C1233 B.n527 VSUBS 0.006853f
C1234 B.n528 VSUBS 0.006853f
C1235 B.n529 VSUBS 0.006853f
C1236 B.n530 VSUBS 0.006853f
C1237 B.n531 VSUBS 0.006853f
C1238 B.n532 VSUBS 0.006853f
C1239 B.n533 VSUBS 0.006853f
C1240 B.n534 VSUBS 0.006853f
C1241 B.n535 VSUBS 0.006853f
C1242 B.n536 VSUBS 0.006853f
C1243 B.n537 VSUBS 0.006853f
C1244 B.n538 VSUBS 0.006853f
C1245 B.n539 VSUBS 0.006853f
C1246 B.n540 VSUBS 0.006853f
C1247 B.n541 VSUBS 0.006853f
C1248 B.n542 VSUBS 0.006853f
C1249 B.n543 VSUBS 0.006853f
C1250 B.n544 VSUBS 0.006853f
C1251 B.n545 VSUBS 0.006853f
C1252 B.n546 VSUBS 0.006853f
C1253 B.n547 VSUBS 0.006853f
C1254 B.n548 VSUBS 0.006853f
C1255 B.n549 VSUBS 0.006853f
C1256 B.n550 VSUBS 0.006853f
C1257 B.n551 VSUBS 0.006853f
C1258 B.n552 VSUBS 0.00645f
C1259 B.n553 VSUBS 0.006853f
C1260 B.n554 VSUBS 0.006853f
C1261 B.n555 VSUBS 0.006853f
C1262 B.n556 VSUBS 0.006853f
C1263 B.n557 VSUBS 0.006853f
C1264 B.n558 VSUBS 0.006853f
C1265 B.n559 VSUBS 0.006853f
C1266 B.n560 VSUBS 0.006853f
C1267 B.n561 VSUBS 0.006853f
C1268 B.n562 VSUBS 0.006853f
C1269 B.n563 VSUBS 0.006853f
C1270 B.n564 VSUBS 0.006853f
C1271 B.n565 VSUBS 0.006853f
C1272 B.n566 VSUBS 0.006853f
C1273 B.n567 VSUBS 0.006853f
C1274 B.n568 VSUBS 0.00383f
C1275 B.n569 VSUBS 0.015877f
C1276 B.n570 VSUBS 0.00645f
C1277 B.n571 VSUBS 0.006853f
C1278 B.n572 VSUBS 0.006853f
C1279 B.n573 VSUBS 0.006853f
C1280 B.n574 VSUBS 0.006853f
C1281 B.n575 VSUBS 0.006853f
C1282 B.n576 VSUBS 0.006853f
C1283 B.n577 VSUBS 0.006853f
C1284 B.n578 VSUBS 0.006853f
C1285 B.n579 VSUBS 0.006853f
C1286 B.n580 VSUBS 0.006853f
C1287 B.n581 VSUBS 0.006853f
C1288 B.n582 VSUBS 0.006853f
C1289 B.n583 VSUBS 0.006853f
C1290 B.n584 VSUBS 0.006853f
C1291 B.n585 VSUBS 0.006853f
C1292 B.n586 VSUBS 0.006853f
C1293 B.n587 VSUBS 0.006853f
C1294 B.n588 VSUBS 0.006853f
C1295 B.n589 VSUBS 0.006853f
C1296 B.n590 VSUBS 0.006853f
C1297 B.n591 VSUBS 0.006853f
C1298 B.n592 VSUBS 0.006853f
C1299 B.n593 VSUBS 0.006853f
C1300 B.n594 VSUBS 0.006853f
C1301 B.n595 VSUBS 0.006853f
C1302 B.n596 VSUBS 0.006853f
C1303 B.n597 VSUBS 0.006853f
C1304 B.n598 VSUBS 0.006853f
C1305 B.n599 VSUBS 0.006853f
C1306 B.n600 VSUBS 0.006853f
C1307 B.n601 VSUBS 0.006853f
C1308 B.n602 VSUBS 0.006853f
C1309 B.n603 VSUBS 0.006853f
C1310 B.n604 VSUBS 0.006853f
C1311 B.n605 VSUBS 0.006853f
C1312 B.n606 VSUBS 0.006853f
C1313 B.n607 VSUBS 0.006853f
C1314 B.n608 VSUBS 0.006853f
C1315 B.n609 VSUBS 0.006853f
C1316 B.n610 VSUBS 0.006853f
C1317 B.n611 VSUBS 0.006853f
C1318 B.n612 VSUBS 0.006853f
C1319 B.n613 VSUBS 0.006853f
C1320 B.n614 VSUBS 0.006853f
C1321 B.n615 VSUBS 0.006853f
C1322 B.n616 VSUBS 0.006853f
C1323 B.n617 VSUBS 0.006853f
C1324 B.n618 VSUBS 0.006853f
C1325 B.n619 VSUBS 0.006853f
C1326 B.n620 VSUBS 0.006853f
C1327 B.n621 VSUBS 0.006853f
C1328 B.n622 VSUBS 0.006853f
C1329 B.n623 VSUBS 0.006853f
C1330 B.n624 VSUBS 0.006853f
C1331 B.n625 VSUBS 0.006853f
C1332 B.n626 VSUBS 0.006853f
C1333 B.n627 VSUBS 0.006853f
C1334 B.n628 VSUBS 0.006853f
C1335 B.n629 VSUBS 0.006853f
C1336 B.n630 VSUBS 0.006853f
C1337 B.n631 VSUBS 0.006853f
C1338 B.n632 VSUBS 0.006853f
C1339 B.n633 VSUBS 0.006853f
C1340 B.n634 VSUBS 0.006853f
C1341 B.n635 VSUBS 0.006853f
C1342 B.n636 VSUBS 0.006853f
C1343 B.n637 VSUBS 0.006853f
C1344 B.n638 VSUBS 0.006853f
C1345 B.n639 VSUBS 0.006853f
C1346 B.n640 VSUBS 0.006853f
C1347 B.n641 VSUBS 0.006853f
C1348 B.n642 VSUBS 0.006853f
C1349 B.n643 VSUBS 0.016042f
C1350 B.n644 VSUBS 0.016042f
C1351 B.n645 VSUBS 0.015199f
C1352 B.n646 VSUBS 0.006853f
C1353 B.n647 VSUBS 0.006853f
C1354 B.n648 VSUBS 0.006853f
C1355 B.n649 VSUBS 0.006853f
C1356 B.n650 VSUBS 0.006853f
C1357 B.n651 VSUBS 0.006853f
C1358 B.n652 VSUBS 0.006853f
C1359 B.n653 VSUBS 0.006853f
C1360 B.n654 VSUBS 0.006853f
C1361 B.n655 VSUBS 0.006853f
C1362 B.n656 VSUBS 0.006853f
C1363 B.n657 VSUBS 0.006853f
C1364 B.n658 VSUBS 0.006853f
C1365 B.n659 VSUBS 0.006853f
C1366 B.n660 VSUBS 0.006853f
C1367 B.n661 VSUBS 0.006853f
C1368 B.n662 VSUBS 0.006853f
C1369 B.n663 VSUBS 0.006853f
C1370 B.n664 VSUBS 0.006853f
C1371 B.n665 VSUBS 0.006853f
C1372 B.n666 VSUBS 0.006853f
C1373 B.n667 VSUBS 0.006853f
C1374 B.n668 VSUBS 0.006853f
C1375 B.n669 VSUBS 0.006853f
C1376 B.n670 VSUBS 0.006853f
C1377 B.n671 VSUBS 0.006853f
C1378 B.n672 VSUBS 0.006853f
C1379 B.n673 VSUBS 0.006853f
C1380 B.n674 VSUBS 0.006853f
C1381 B.n675 VSUBS 0.006853f
C1382 B.n676 VSUBS 0.006853f
C1383 B.n677 VSUBS 0.006853f
C1384 B.n678 VSUBS 0.006853f
C1385 B.n679 VSUBS 0.006853f
C1386 B.n680 VSUBS 0.006853f
C1387 B.n681 VSUBS 0.006853f
C1388 B.n682 VSUBS 0.006853f
C1389 B.n683 VSUBS 0.006853f
C1390 B.n684 VSUBS 0.006853f
C1391 B.n685 VSUBS 0.006853f
C1392 B.n686 VSUBS 0.006853f
C1393 B.n687 VSUBS 0.008943f
C1394 B.n688 VSUBS 0.009526f
C1395 B.n689 VSUBS 0.018944f
.ends

