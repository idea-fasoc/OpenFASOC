* NGSPICE file created from diff_pair_sample_1045.ext - technology: sky130A

.subckt diff_pair_sample_1045 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2938_n2308# sky130_fd_pr__pfet_01v8 ad=2.613 pd=14.18 as=0 ps=0 w=6.7 l=2.95
X1 B.t8 B.t6 B.t7 w_n2938_n2308# sky130_fd_pr__pfet_01v8 ad=2.613 pd=14.18 as=0 ps=0 w=6.7 l=2.95
X2 B.t5 B.t3 B.t4 w_n2938_n2308# sky130_fd_pr__pfet_01v8 ad=2.613 pd=14.18 as=0 ps=0 w=6.7 l=2.95
X3 B.t2 B.t0 B.t1 w_n2938_n2308# sky130_fd_pr__pfet_01v8 ad=2.613 pd=14.18 as=0 ps=0 w=6.7 l=2.95
X4 VDD2.t3 VN.t0 VTAIL.t5 w_n2938_n2308# sky130_fd_pr__pfet_01v8 ad=1.1055 pd=7.03 as=2.613 ps=14.18 w=6.7 l=2.95
X5 VTAIL.t6 VN.t1 VDD2.t2 w_n2938_n2308# sky130_fd_pr__pfet_01v8 ad=2.613 pd=14.18 as=1.1055 ps=7.03 w=6.7 l=2.95
X6 VTAIL.t7 VN.t2 VDD2.t1 w_n2938_n2308# sky130_fd_pr__pfet_01v8 ad=2.613 pd=14.18 as=1.1055 ps=7.03 w=6.7 l=2.95
X7 VDD1.t3 VP.t0 VTAIL.t3 w_n2938_n2308# sky130_fd_pr__pfet_01v8 ad=1.1055 pd=7.03 as=2.613 ps=14.18 w=6.7 l=2.95
X8 VDD1.t2 VP.t1 VTAIL.t1 w_n2938_n2308# sky130_fd_pr__pfet_01v8 ad=1.1055 pd=7.03 as=2.613 ps=14.18 w=6.7 l=2.95
X9 VTAIL.t2 VP.t2 VDD1.t1 w_n2938_n2308# sky130_fd_pr__pfet_01v8 ad=2.613 pd=14.18 as=1.1055 ps=7.03 w=6.7 l=2.95
X10 VDD2.t0 VN.t3 VTAIL.t4 w_n2938_n2308# sky130_fd_pr__pfet_01v8 ad=1.1055 pd=7.03 as=2.613 ps=14.18 w=6.7 l=2.95
X11 VTAIL.t0 VP.t3 VDD1.t0 w_n2938_n2308# sky130_fd_pr__pfet_01v8 ad=2.613 pd=14.18 as=1.1055 ps=7.03 w=6.7 l=2.95
R0 B.n409 B.n56 585
R1 B.n411 B.n410 585
R2 B.n412 B.n55 585
R3 B.n414 B.n413 585
R4 B.n415 B.n54 585
R5 B.n417 B.n416 585
R6 B.n418 B.n53 585
R7 B.n420 B.n419 585
R8 B.n421 B.n52 585
R9 B.n423 B.n422 585
R10 B.n424 B.n51 585
R11 B.n426 B.n425 585
R12 B.n427 B.n50 585
R13 B.n429 B.n428 585
R14 B.n430 B.n49 585
R15 B.n432 B.n431 585
R16 B.n433 B.n48 585
R17 B.n435 B.n434 585
R18 B.n436 B.n47 585
R19 B.n438 B.n437 585
R20 B.n439 B.n46 585
R21 B.n441 B.n440 585
R22 B.n442 B.n45 585
R23 B.n444 B.n443 585
R24 B.n445 B.n41 585
R25 B.n447 B.n446 585
R26 B.n448 B.n40 585
R27 B.n450 B.n449 585
R28 B.n451 B.n39 585
R29 B.n453 B.n452 585
R30 B.n454 B.n38 585
R31 B.n456 B.n455 585
R32 B.n457 B.n37 585
R33 B.n459 B.n458 585
R34 B.n460 B.n36 585
R35 B.n462 B.n461 585
R36 B.n464 B.n33 585
R37 B.n466 B.n465 585
R38 B.n467 B.n32 585
R39 B.n469 B.n468 585
R40 B.n470 B.n31 585
R41 B.n472 B.n471 585
R42 B.n473 B.n30 585
R43 B.n475 B.n474 585
R44 B.n476 B.n29 585
R45 B.n478 B.n477 585
R46 B.n479 B.n28 585
R47 B.n481 B.n480 585
R48 B.n482 B.n27 585
R49 B.n484 B.n483 585
R50 B.n485 B.n26 585
R51 B.n487 B.n486 585
R52 B.n488 B.n25 585
R53 B.n490 B.n489 585
R54 B.n491 B.n24 585
R55 B.n493 B.n492 585
R56 B.n494 B.n23 585
R57 B.n496 B.n495 585
R58 B.n497 B.n22 585
R59 B.n499 B.n498 585
R60 B.n500 B.n21 585
R61 B.n502 B.n501 585
R62 B.n408 B.n407 585
R63 B.n406 B.n57 585
R64 B.n405 B.n404 585
R65 B.n403 B.n58 585
R66 B.n402 B.n401 585
R67 B.n400 B.n59 585
R68 B.n399 B.n398 585
R69 B.n397 B.n60 585
R70 B.n396 B.n395 585
R71 B.n394 B.n61 585
R72 B.n393 B.n392 585
R73 B.n391 B.n62 585
R74 B.n390 B.n389 585
R75 B.n388 B.n63 585
R76 B.n387 B.n386 585
R77 B.n385 B.n64 585
R78 B.n384 B.n383 585
R79 B.n382 B.n65 585
R80 B.n381 B.n380 585
R81 B.n379 B.n66 585
R82 B.n378 B.n377 585
R83 B.n376 B.n67 585
R84 B.n375 B.n374 585
R85 B.n373 B.n68 585
R86 B.n372 B.n371 585
R87 B.n370 B.n69 585
R88 B.n369 B.n368 585
R89 B.n367 B.n70 585
R90 B.n366 B.n365 585
R91 B.n364 B.n71 585
R92 B.n363 B.n362 585
R93 B.n361 B.n72 585
R94 B.n360 B.n359 585
R95 B.n358 B.n73 585
R96 B.n357 B.n356 585
R97 B.n355 B.n74 585
R98 B.n354 B.n353 585
R99 B.n352 B.n75 585
R100 B.n351 B.n350 585
R101 B.n349 B.n76 585
R102 B.n348 B.n347 585
R103 B.n346 B.n77 585
R104 B.n345 B.n344 585
R105 B.n343 B.n78 585
R106 B.n342 B.n341 585
R107 B.n340 B.n79 585
R108 B.n339 B.n338 585
R109 B.n337 B.n80 585
R110 B.n336 B.n335 585
R111 B.n334 B.n81 585
R112 B.n333 B.n332 585
R113 B.n331 B.n82 585
R114 B.n330 B.n329 585
R115 B.n328 B.n83 585
R116 B.n327 B.n326 585
R117 B.n325 B.n84 585
R118 B.n324 B.n323 585
R119 B.n322 B.n85 585
R120 B.n321 B.n320 585
R121 B.n319 B.n86 585
R122 B.n318 B.n317 585
R123 B.n316 B.n87 585
R124 B.n315 B.n314 585
R125 B.n313 B.n88 585
R126 B.n312 B.n311 585
R127 B.n310 B.n89 585
R128 B.n309 B.n308 585
R129 B.n307 B.n90 585
R130 B.n306 B.n305 585
R131 B.n304 B.n91 585
R132 B.n303 B.n302 585
R133 B.n301 B.n92 585
R134 B.n300 B.n299 585
R135 B.n298 B.n93 585
R136 B.n297 B.n296 585
R137 B.n202 B.n129 585
R138 B.n204 B.n203 585
R139 B.n205 B.n128 585
R140 B.n207 B.n206 585
R141 B.n208 B.n127 585
R142 B.n210 B.n209 585
R143 B.n211 B.n126 585
R144 B.n213 B.n212 585
R145 B.n214 B.n125 585
R146 B.n216 B.n215 585
R147 B.n217 B.n124 585
R148 B.n219 B.n218 585
R149 B.n220 B.n123 585
R150 B.n222 B.n221 585
R151 B.n223 B.n122 585
R152 B.n225 B.n224 585
R153 B.n226 B.n121 585
R154 B.n228 B.n227 585
R155 B.n229 B.n120 585
R156 B.n231 B.n230 585
R157 B.n232 B.n119 585
R158 B.n234 B.n233 585
R159 B.n235 B.n118 585
R160 B.n237 B.n236 585
R161 B.n238 B.n117 585
R162 B.n240 B.n239 585
R163 B.n242 B.n114 585
R164 B.n244 B.n243 585
R165 B.n245 B.n113 585
R166 B.n247 B.n246 585
R167 B.n248 B.n112 585
R168 B.n250 B.n249 585
R169 B.n251 B.n111 585
R170 B.n253 B.n252 585
R171 B.n254 B.n110 585
R172 B.n256 B.n255 585
R173 B.n258 B.n257 585
R174 B.n259 B.n106 585
R175 B.n261 B.n260 585
R176 B.n262 B.n105 585
R177 B.n264 B.n263 585
R178 B.n265 B.n104 585
R179 B.n267 B.n266 585
R180 B.n268 B.n103 585
R181 B.n270 B.n269 585
R182 B.n271 B.n102 585
R183 B.n273 B.n272 585
R184 B.n274 B.n101 585
R185 B.n276 B.n275 585
R186 B.n277 B.n100 585
R187 B.n279 B.n278 585
R188 B.n280 B.n99 585
R189 B.n282 B.n281 585
R190 B.n283 B.n98 585
R191 B.n285 B.n284 585
R192 B.n286 B.n97 585
R193 B.n288 B.n287 585
R194 B.n289 B.n96 585
R195 B.n291 B.n290 585
R196 B.n292 B.n95 585
R197 B.n294 B.n293 585
R198 B.n295 B.n94 585
R199 B.n201 B.n200 585
R200 B.n199 B.n130 585
R201 B.n198 B.n197 585
R202 B.n196 B.n131 585
R203 B.n195 B.n194 585
R204 B.n193 B.n132 585
R205 B.n192 B.n191 585
R206 B.n190 B.n133 585
R207 B.n189 B.n188 585
R208 B.n187 B.n134 585
R209 B.n186 B.n185 585
R210 B.n184 B.n135 585
R211 B.n183 B.n182 585
R212 B.n181 B.n136 585
R213 B.n180 B.n179 585
R214 B.n178 B.n137 585
R215 B.n177 B.n176 585
R216 B.n175 B.n138 585
R217 B.n174 B.n173 585
R218 B.n172 B.n139 585
R219 B.n171 B.n170 585
R220 B.n169 B.n140 585
R221 B.n168 B.n167 585
R222 B.n166 B.n141 585
R223 B.n165 B.n164 585
R224 B.n163 B.n142 585
R225 B.n162 B.n161 585
R226 B.n160 B.n143 585
R227 B.n159 B.n158 585
R228 B.n157 B.n144 585
R229 B.n156 B.n155 585
R230 B.n154 B.n145 585
R231 B.n153 B.n152 585
R232 B.n151 B.n146 585
R233 B.n150 B.n149 585
R234 B.n148 B.n147 585
R235 B.n2 B.n0 585
R236 B.n557 B.n1 585
R237 B.n556 B.n555 585
R238 B.n554 B.n3 585
R239 B.n553 B.n552 585
R240 B.n551 B.n4 585
R241 B.n550 B.n549 585
R242 B.n548 B.n5 585
R243 B.n547 B.n546 585
R244 B.n545 B.n6 585
R245 B.n544 B.n543 585
R246 B.n542 B.n7 585
R247 B.n541 B.n540 585
R248 B.n539 B.n8 585
R249 B.n538 B.n537 585
R250 B.n536 B.n9 585
R251 B.n535 B.n534 585
R252 B.n533 B.n10 585
R253 B.n532 B.n531 585
R254 B.n530 B.n11 585
R255 B.n529 B.n528 585
R256 B.n527 B.n12 585
R257 B.n526 B.n525 585
R258 B.n524 B.n13 585
R259 B.n523 B.n522 585
R260 B.n521 B.n14 585
R261 B.n520 B.n519 585
R262 B.n518 B.n15 585
R263 B.n517 B.n516 585
R264 B.n515 B.n16 585
R265 B.n514 B.n513 585
R266 B.n512 B.n17 585
R267 B.n511 B.n510 585
R268 B.n509 B.n18 585
R269 B.n508 B.n507 585
R270 B.n506 B.n19 585
R271 B.n505 B.n504 585
R272 B.n503 B.n20 585
R273 B.n559 B.n558 585
R274 B.n202 B.n201 478.086
R275 B.n503 B.n502 478.086
R276 B.n297 B.n94 478.086
R277 B.n407 B.n56 478.086
R278 B.n107 B.t5 344.187
R279 B.n42 B.t1 344.187
R280 B.n115 B.t8 344.187
R281 B.n34 B.t10 344.187
R282 B.n108 B.t4 280.575
R283 B.n43 B.t2 280.575
R284 B.n116 B.t7 280.575
R285 B.n35 B.t11 280.575
R286 B.n107 B.t3 263.257
R287 B.n115 B.t6 263.257
R288 B.n34 B.t9 263.257
R289 B.n42 B.t0 263.257
R290 B.n201 B.n130 163.367
R291 B.n197 B.n130 163.367
R292 B.n197 B.n196 163.367
R293 B.n196 B.n195 163.367
R294 B.n195 B.n132 163.367
R295 B.n191 B.n132 163.367
R296 B.n191 B.n190 163.367
R297 B.n190 B.n189 163.367
R298 B.n189 B.n134 163.367
R299 B.n185 B.n134 163.367
R300 B.n185 B.n184 163.367
R301 B.n184 B.n183 163.367
R302 B.n183 B.n136 163.367
R303 B.n179 B.n136 163.367
R304 B.n179 B.n178 163.367
R305 B.n178 B.n177 163.367
R306 B.n177 B.n138 163.367
R307 B.n173 B.n138 163.367
R308 B.n173 B.n172 163.367
R309 B.n172 B.n171 163.367
R310 B.n171 B.n140 163.367
R311 B.n167 B.n140 163.367
R312 B.n167 B.n166 163.367
R313 B.n166 B.n165 163.367
R314 B.n165 B.n142 163.367
R315 B.n161 B.n142 163.367
R316 B.n161 B.n160 163.367
R317 B.n160 B.n159 163.367
R318 B.n159 B.n144 163.367
R319 B.n155 B.n144 163.367
R320 B.n155 B.n154 163.367
R321 B.n154 B.n153 163.367
R322 B.n153 B.n146 163.367
R323 B.n149 B.n146 163.367
R324 B.n149 B.n148 163.367
R325 B.n148 B.n2 163.367
R326 B.n558 B.n2 163.367
R327 B.n558 B.n557 163.367
R328 B.n557 B.n556 163.367
R329 B.n556 B.n3 163.367
R330 B.n552 B.n3 163.367
R331 B.n552 B.n551 163.367
R332 B.n551 B.n550 163.367
R333 B.n550 B.n5 163.367
R334 B.n546 B.n5 163.367
R335 B.n546 B.n545 163.367
R336 B.n545 B.n544 163.367
R337 B.n544 B.n7 163.367
R338 B.n540 B.n7 163.367
R339 B.n540 B.n539 163.367
R340 B.n539 B.n538 163.367
R341 B.n538 B.n9 163.367
R342 B.n534 B.n9 163.367
R343 B.n534 B.n533 163.367
R344 B.n533 B.n532 163.367
R345 B.n532 B.n11 163.367
R346 B.n528 B.n11 163.367
R347 B.n528 B.n527 163.367
R348 B.n527 B.n526 163.367
R349 B.n526 B.n13 163.367
R350 B.n522 B.n13 163.367
R351 B.n522 B.n521 163.367
R352 B.n521 B.n520 163.367
R353 B.n520 B.n15 163.367
R354 B.n516 B.n15 163.367
R355 B.n516 B.n515 163.367
R356 B.n515 B.n514 163.367
R357 B.n514 B.n17 163.367
R358 B.n510 B.n17 163.367
R359 B.n510 B.n509 163.367
R360 B.n509 B.n508 163.367
R361 B.n508 B.n19 163.367
R362 B.n504 B.n19 163.367
R363 B.n504 B.n503 163.367
R364 B.n203 B.n202 163.367
R365 B.n203 B.n128 163.367
R366 B.n207 B.n128 163.367
R367 B.n208 B.n207 163.367
R368 B.n209 B.n208 163.367
R369 B.n209 B.n126 163.367
R370 B.n213 B.n126 163.367
R371 B.n214 B.n213 163.367
R372 B.n215 B.n214 163.367
R373 B.n215 B.n124 163.367
R374 B.n219 B.n124 163.367
R375 B.n220 B.n219 163.367
R376 B.n221 B.n220 163.367
R377 B.n221 B.n122 163.367
R378 B.n225 B.n122 163.367
R379 B.n226 B.n225 163.367
R380 B.n227 B.n226 163.367
R381 B.n227 B.n120 163.367
R382 B.n231 B.n120 163.367
R383 B.n232 B.n231 163.367
R384 B.n233 B.n232 163.367
R385 B.n233 B.n118 163.367
R386 B.n237 B.n118 163.367
R387 B.n238 B.n237 163.367
R388 B.n239 B.n238 163.367
R389 B.n239 B.n114 163.367
R390 B.n244 B.n114 163.367
R391 B.n245 B.n244 163.367
R392 B.n246 B.n245 163.367
R393 B.n246 B.n112 163.367
R394 B.n250 B.n112 163.367
R395 B.n251 B.n250 163.367
R396 B.n252 B.n251 163.367
R397 B.n252 B.n110 163.367
R398 B.n256 B.n110 163.367
R399 B.n257 B.n256 163.367
R400 B.n257 B.n106 163.367
R401 B.n261 B.n106 163.367
R402 B.n262 B.n261 163.367
R403 B.n263 B.n262 163.367
R404 B.n263 B.n104 163.367
R405 B.n267 B.n104 163.367
R406 B.n268 B.n267 163.367
R407 B.n269 B.n268 163.367
R408 B.n269 B.n102 163.367
R409 B.n273 B.n102 163.367
R410 B.n274 B.n273 163.367
R411 B.n275 B.n274 163.367
R412 B.n275 B.n100 163.367
R413 B.n279 B.n100 163.367
R414 B.n280 B.n279 163.367
R415 B.n281 B.n280 163.367
R416 B.n281 B.n98 163.367
R417 B.n285 B.n98 163.367
R418 B.n286 B.n285 163.367
R419 B.n287 B.n286 163.367
R420 B.n287 B.n96 163.367
R421 B.n291 B.n96 163.367
R422 B.n292 B.n291 163.367
R423 B.n293 B.n292 163.367
R424 B.n293 B.n94 163.367
R425 B.n298 B.n297 163.367
R426 B.n299 B.n298 163.367
R427 B.n299 B.n92 163.367
R428 B.n303 B.n92 163.367
R429 B.n304 B.n303 163.367
R430 B.n305 B.n304 163.367
R431 B.n305 B.n90 163.367
R432 B.n309 B.n90 163.367
R433 B.n310 B.n309 163.367
R434 B.n311 B.n310 163.367
R435 B.n311 B.n88 163.367
R436 B.n315 B.n88 163.367
R437 B.n316 B.n315 163.367
R438 B.n317 B.n316 163.367
R439 B.n317 B.n86 163.367
R440 B.n321 B.n86 163.367
R441 B.n322 B.n321 163.367
R442 B.n323 B.n322 163.367
R443 B.n323 B.n84 163.367
R444 B.n327 B.n84 163.367
R445 B.n328 B.n327 163.367
R446 B.n329 B.n328 163.367
R447 B.n329 B.n82 163.367
R448 B.n333 B.n82 163.367
R449 B.n334 B.n333 163.367
R450 B.n335 B.n334 163.367
R451 B.n335 B.n80 163.367
R452 B.n339 B.n80 163.367
R453 B.n340 B.n339 163.367
R454 B.n341 B.n340 163.367
R455 B.n341 B.n78 163.367
R456 B.n345 B.n78 163.367
R457 B.n346 B.n345 163.367
R458 B.n347 B.n346 163.367
R459 B.n347 B.n76 163.367
R460 B.n351 B.n76 163.367
R461 B.n352 B.n351 163.367
R462 B.n353 B.n352 163.367
R463 B.n353 B.n74 163.367
R464 B.n357 B.n74 163.367
R465 B.n358 B.n357 163.367
R466 B.n359 B.n358 163.367
R467 B.n359 B.n72 163.367
R468 B.n363 B.n72 163.367
R469 B.n364 B.n363 163.367
R470 B.n365 B.n364 163.367
R471 B.n365 B.n70 163.367
R472 B.n369 B.n70 163.367
R473 B.n370 B.n369 163.367
R474 B.n371 B.n370 163.367
R475 B.n371 B.n68 163.367
R476 B.n375 B.n68 163.367
R477 B.n376 B.n375 163.367
R478 B.n377 B.n376 163.367
R479 B.n377 B.n66 163.367
R480 B.n381 B.n66 163.367
R481 B.n382 B.n381 163.367
R482 B.n383 B.n382 163.367
R483 B.n383 B.n64 163.367
R484 B.n387 B.n64 163.367
R485 B.n388 B.n387 163.367
R486 B.n389 B.n388 163.367
R487 B.n389 B.n62 163.367
R488 B.n393 B.n62 163.367
R489 B.n394 B.n393 163.367
R490 B.n395 B.n394 163.367
R491 B.n395 B.n60 163.367
R492 B.n399 B.n60 163.367
R493 B.n400 B.n399 163.367
R494 B.n401 B.n400 163.367
R495 B.n401 B.n58 163.367
R496 B.n405 B.n58 163.367
R497 B.n406 B.n405 163.367
R498 B.n407 B.n406 163.367
R499 B.n502 B.n21 163.367
R500 B.n498 B.n21 163.367
R501 B.n498 B.n497 163.367
R502 B.n497 B.n496 163.367
R503 B.n496 B.n23 163.367
R504 B.n492 B.n23 163.367
R505 B.n492 B.n491 163.367
R506 B.n491 B.n490 163.367
R507 B.n490 B.n25 163.367
R508 B.n486 B.n25 163.367
R509 B.n486 B.n485 163.367
R510 B.n485 B.n484 163.367
R511 B.n484 B.n27 163.367
R512 B.n480 B.n27 163.367
R513 B.n480 B.n479 163.367
R514 B.n479 B.n478 163.367
R515 B.n478 B.n29 163.367
R516 B.n474 B.n29 163.367
R517 B.n474 B.n473 163.367
R518 B.n473 B.n472 163.367
R519 B.n472 B.n31 163.367
R520 B.n468 B.n31 163.367
R521 B.n468 B.n467 163.367
R522 B.n467 B.n466 163.367
R523 B.n466 B.n33 163.367
R524 B.n461 B.n33 163.367
R525 B.n461 B.n460 163.367
R526 B.n460 B.n459 163.367
R527 B.n459 B.n37 163.367
R528 B.n455 B.n37 163.367
R529 B.n455 B.n454 163.367
R530 B.n454 B.n453 163.367
R531 B.n453 B.n39 163.367
R532 B.n449 B.n39 163.367
R533 B.n449 B.n448 163.367
R534 B.n448 B.n447 163.367
R535 B.n447 B.n41 163.367
R536 B.n443 B.n41 163.367
R537 B.n443 B.n442 163.367
R538 B.n442 B.n441 163.367
R539 B.n441 B.n46 163.367
R540 B.n437 B.n46 163.367
R541 B.n437 B.n436 163.367
R542 B.n436 B.n435 163.367
R543 B.n435 B.n48 163.367
R544 B.n431 B.n48 163.367
R545 B.n431 B.n430 163.367
R546 B.n430 B.n429 163.367
R547 B.n429 B.n50 163.367
R548 B.n425 B.n50 163.367
R549 B.n425 B.n424 163.367
R550 B.n424 B.n423 163.367
R551 B.n423 B.n52 163.367
R552 B.n419 B.n52 163.367
R553 B.n419 B.n418 163.367
R554 B.n418 B.n417 163.367
R555 B.n417 B.n54 163.367
R556 B.n413 B.n54 163.367
R557 B.n413 B.n412 163.367
R558 B.n412 B.n411 163.367
R559 B.n411 B.n56 163.367
R560 B.n108 B.n107 63.6126
R561 B.n116 B.n115 63.6126
R562 B.n35 B.n34 63.6126
R563 B.n43 B.n42 63.6126
R564 B.n109 B.n108 59.5399
R565 B.n241 B.n116 59.5399
R566 B.n463 B.n35 59.5399
R567 B.n44 B.n43 59.5399
R568 B.n501 B.n20 31.0639
R569 B.n409 B.n408 31.0639
R570 B.n296 B.n295 31.0639
R571 B.n200 B.n129 31.0639
R572 B B.n559 18.0485
R573 B.n501 B.n500 10.6151
R574 B.n500 B.n499 10.6151
R575 B.n499 B.n22 10.6151
R576 B.n495 B.n22 10.6151
R577 B.n495 B.n494 10.6151
R578 B.n494 B.n493 10.6151
R579 B.n493 B.n24 10.6151
R580 B.n489 B.n24 10.6151
R581 B.n489 B.n488 10.6151
R582 B.n488 B.n487 10.6151
R583 B.n487 B.n26 10.6151
R584 B.n483 B.n26 10.6151
R585 B.n483 B.n482 10.6151
R586 B.n482 B.n481 10.6151
R587 B.n481 B.n28 10.6151
R588 B.n477 B.n28 10.6151
R589 B.n477 B.n476 10.6151
R590 B.n476 B.n475 10.6151
R591 B.n475 B.n30 10.6151
R592 B.n471 B.n30 10.6151
R593 B.n471 B.n470 10.6151
R594 B.n470 B.n469 10.6151
R595 B.n469 B.n32 10.6151
R596 B.n465 B.n32 10.6151
R597 B.n465 B.n464 10.6151
R598 B.n462 B.n36 10.6151
R599 B.n458 B.n36 10.6151
R600 B.n458 B.n457 10.6151
R601 B.n457 B.n456 10.6151
R602 B.n456 B.n38 10.6151
R603 B.n452 B.n38 10.6151
R604 B.n452 B.n451 10.6151
R605 B.n451 B.n450 10.6151
R606 B.n450 B.n40 10.6151
R607 B.n446 B.n445 10.6151
R608 B.n445 B.n444 10.6151
R609 B.n444 B.n45 10.6151
R610 B.n440 B.n45 10.6151
R611 B.n440 B.n439 10.6151
R612 B.n439 B.n438 10.6151
R613 B.n438 B.n47 10.6151
R614 B.n434 B.n47 10.6151
R615 B.n434 B.n433 10.6151
R616 B.n433 B.n432 10.6151
R617 B.n432 B.n49 10.6151
R618 B.n428 B.n49 10.6151
R619 B.n428 B.n427 10.6151
R620 B.n427 B.n426 10.6151
R621 B.n426 B.n51 10.6151
R622 B.n422 B.n51 10.6151
R623 B.n422 B.n421 10.6151
R624 B.n421 B.n420 10.6151
R625 B.n420 B.n53 10.6151
R626 B.n416 B.n53 10.6151
R627 B.n416 B.n415 10.6151
R628 B.n415 B.n414 10.6151
R629 B.n414 B.n55 10.6151
R630 B.n410 B.n55 10.6151
R631 B.n410 B.n409 10.6151
R632 B.n296 B.n93 10.6151
R633 B.n300 B.n93 10.6151
R634 B.n301 B.n300 10.6151
R635 B.n302 B.n301 10.6151
R636 B.n302 B.n91 10.6151
R637 B.n306 B.n91 10.6151
R638 B.n307 B.n306 10.6151
R639 B.n308 B.n307 10.6151
R640 B.n308 B.n89 10.6151
R641 B.n312 B.n89 10.6151
R642 B.n313 B.n312 10.6151
R643 B.n314 B.n313 10.6151
R644 B.n314 B.n87 10.6151
R645 B.n318 B.n87 10.6151
R646 B.n319 B.n318 10.6151
R647 B.n320 B.n319 10.6151
R648 B.n320 B.n85 10.6151
R649 B.n324 B.n85 10.6151
R650 B.n325 B.n324 10.6151
R651 B.n326 B.n325 10.6151
R652 B.n326 B.n83 10.6151
R653 B.n330 B.n83 10.6151
R654 B.n331 B.n330 10.6151
R655 B.n332 B.n331 10.6151
R656 B.n332 B.n81 10.6151
R657 B.n336 B.n81 10.6151
R658 B.n337 B.n336 10.6151
R659 B.n338 B.n337 10.6151
R660 B.n338 B.n79 10.6151
R661 B.n342 B.n79 10.6151
R662 B.n343 B.n342 10.6151
R663 B.n344 B.n343 10.6151
R664 B.n344 B.n77 10.6151
R665 B.n348 B.n77 10.6151
R666 B.n349 B.n348 10.6151
R667 B.n350 B.n349 10.6151
R668 B.n350 B.n75 10.6151
R669 B.n354 B.n75 10.6151
R670 B.n355 B.n354 10.6151
R671 B.n356 B.n355 10.6151
R672 B.n356 B.n73 10.6151
R673 B.n360 B.n73 10.6151
R674 B.n361 B.n360 10.6151
R675 B.n362 B.n361 10.6151
R676 B.n362 B.n71 10.6151
R677 B.n366 B.n71 10.6151
R678 B.n367 B.n366 10.6151
R679 B.n368 B.n367 10.6151
R680 B.n368 B.n69 10.6151
R681 B.n372 B.n69 10.6151
R682 B.n373 B.n372 10.6151
R683 B.n374 B.n373 10.6151
R684 B.n374 B.n67 10.6151
R685 B.n378 B.n67 10.6151
R686 B.n379 B.n378 10.6151
R687 B.n380 B.n379 10.6151
R688 B.n380 B.n65 10.6151
R689 B.n384 B.n65 10.6151
R690 B.n385 B.n384 10.6151
R691 B.n386 B.n385 10.6151
R692 B.n386 B.n63 10.6151
R693 B.n390 B.n63 10.6151
R694 B.n391 B.n390 10.6151
R695 B.n392 B.n391 10.6151
R696 B.n392 B.n61 10.6151
R697 B.n396 B.n61 10.6151
R698 B.n397 B.n396 10.6151
R699 B.n398 B.n397 10.6151
R700 B.n398 B.n59 10.6151
R701 B.n402 B.n59 10.6151
R702 B.n403 B.n402 10.6151
R703 B.n404 B.n403 10.6151
R704 B.n404 B.n57 10.6151
R705 B.n408 B.n57 10.6151
R706 B.n204 B.n129 10.6151
R707 B.n205 B.n204 10.6151
R708 B.n206 B.n205 10.6151
R709 B.n206 B.n127 10.6151
R710 B.n210 B.n127 10.6151
R711 B.n211 B.n210 10.6151
R712 B.n212 B.n211 10.6151
R713 B.n212 B.n125 10.6151
R714 B.n216 B.n125 10.6151
R715 B.n217 B.n216 10.6151
R716 B.n218 B.n217 10.6151
R717 B.n218 B.n123 10.6151
R718 B.n222 B.n123 10.6151
R719 B.n223 B.n222 10.6151
R720 B.n224 B.n223 10.6151
R721 B.n224 B.n121 10.6151
R722 B.n228 B.n121 10.6151
R723 B.n229 B.n228 10.6151
R724 B.n230 B.n229 10.6151
R725 B.n230 B.n119 10.6151
R726 B.n234 B.n119 10.6151
R727 B.n235 B.n234 10.6151
R728 B.n236 B.n235 10.6151
R729 B.n236 B.n117 10.6151
R730 B.n240 B.n117 10.6151
R731 B.n243 B.n242 10.6151
R732 B.n243 B.n113 10.6151
R733 B.n247 B.n113 10.6151
R734 B.n248 B.n247 10.6151
R735 B.n249 B.n248 10.6151
R736 B.n249 B.n111 10.6151
R737 B.n253 B.n111 10.6151
R738 B.n254 B.n253 10.6151
R739 B.n255 B.n254 10.6151
R740 B.n259 B.n258 10.6151
R741 B.n260 B.n259 10.6151
R742 B.n260 B.n105 10.6151
R743 B.n264 B.n105 10.6151
R744 B.n265 B.n264 10.6151
R745 B.n266 B.n265 10.6151
R746 B.n266 B.n103 10.6151
R747 B.n270 B.n103 10.6151
R748 B.n271 B.n270 10.6151
R749 B.n272 B.n271 10.6151
R750 B.n272 B.n101 10.6151
R751 B.n276 B.n101 10.6151
R752 B.n277 B.n276 10.6151
R753 B.n278 B.n277 10.6151
R754 B.n278 B.n99 10.6151
R755 B.n282 B.n99 10.6151
R756 B.n283 B.n282 10.6151
R757 B.n284 B.n283 10.6151
R758 B.n284 B.n97 10.6151
R759 B.n288 B.n97 10.6151
R760 B.n289 B.n288 10.6151
R761 B.n290 B.n289 10.6151
R762 B.n290 B.n95 10.6151
R763 B.n294 B.n95 10.6151
R764 B.n295 B.n294 10.6151
R765 B.n200 B.n199 10.6151
R766 B.n199 B.n198 10.6151
R767 B.n198 B.n131 10.6151
R768 B.n194 B.n131 10.6151
R769 B.n194 B.n193 10.6151
R770 B.n193 B.n192 10.6151
R771 B.n192 B.n133 10.6151
R772 B.n188 B.n133 10.6151
R773 B.n188 B.n187 10.6151
R774 B.n187 B.n186 10.6151
R775 B.n186 B.n135 10.6151
R776 B.n182 B.n135 10.6151
R777 B.n182 B.n181 10.6151
R778 B.n181 B.n180 10.6151
R779 B.n180 B.n137 10.6151
R780 B.n176 B.n137 10.6151
R781 B.n176 B.n175 10.6151
R782 B.n175 B.n174 10.6151
R783 B.n174 B.n139 10.6151
R784 B.n170 B.n139 10.6151
R785 B.n170 B.n169 10.6151
R786 B.n169 B.n168 10.6151
R787 B.n168 B.n141 10.6151
R788 B.n164 B.n141 10.6151
R789 B.n164 B.n163 10.6151
R790 B.n163 B.n162 10.6151
R791 B.n162 B.n143 10.6151
R792 B.n158 B.n143 10.6151
R793 B.n158 B.n157 10.6151
R794 B.n157 B.n156 10.6151
R795 B.n156 B.n145 10.6151
R796 B.n152 B.n145 10.6151
R797 B.n152 B.n151 10.6151
R798 B.n151 B.n150 10.6151
R799 B.n150 B.n147 10.6151
R800 B.n147 B.n0 10.6151
R801 B.n555 B.n1 10.6151
R802 B.n555 B.n554 10.6151
R803 B.n554 B.n553 10.6151
R804 B.n553 B.n4 10.6151
R805 B.n549 B.n4 10.6151
R806 B.n549 B.n548 10.6151
R807 B.n548 B.n547 10.6151
R808 B.n547 B.n6 10.6151
R809 B.n543 B.n6 10.6151
R810 B.n543 B.n542 10.6151
R811 B.n542 B.n541 10.6151
R812 B.n541 B.n8 10.6151
R813 B.n537 B.n8 10.6151
R814 B.n537 B.n536 10.6151
R815 B.n536 B.n535 10.6151
R816 B.n535 B.n10 10.6151
R817 B.n531 B.n10 10.6151
R818 B.n531 B.n530 10.6151
R819 B.n530 B.n529 10.6151
R820 B.n529 B.n12 10.6151
R821 B.n525 B.n12 10.6151
R822 B.n525 B.n524 10.6151
R823 B.n524 B.n523 10.6151
R824 B.n523 B.n14 10.6151
R825 B.n519 B.n14 10.6151
R826 B.n519 B.n518 10.6151
R827 B.n518 B.n517 10.6151
R828 B.n517 B.n16 10.6151
R829 B.n513 B.n16 10.6151
R830 B.n513 B.n512 10.6151
R831 B.n512 B.n511 10.6151
R832 B.n511 B.n18 10.6151
R833 B.n507 B.n18 10.6151
R834 B.n507 B.n506 10.6151
R835 B.n506 B.n505 10.6151
R836 B.n505 B.n20 10.6151
R837 B.n464 B.n463 9.36635
R838 B.n446 B.n44 9.36635
R839 B.n241 B.n240 9.36635
R840 B.n258 B.n109 9.36635
R841 B.n559 B.n0 2.81026
R842 B.n559 B.n1 2.81026
R843 B.n463 B.n462 1.24928
R844 B.n44 B.n40 1.24928
R845 B.n242 B.n241 1.24928
R846 B.n255 B.n109 1.24928
R847 VN.n0 VN.t2 89.1887
R848 VN.n1 VN.t0 89.1887
R849 VN.n0 VN.t3 88.2078
R850 VN.n1 VN.t1 88.2078
R851 VN VN.n1 46.6308
R852 VN VN.n0 3.08916
R853 VTAIL.n282 VTAIL.n252 756.745
R854 VTAIL.n30 VTAIL.n0 756.745
R855 VTAIL.n66 VTAIL.n36 756.745
R856 VTAIL.n102 VTAIL.n72 756.745
R857 VTAIL.n246 VTAIL.n216 756.745
R858 VTAIL.n210 VTAIL.n180 756.745
R859 VTAIL.n174 VTAIL.n144 756.745
R860 VTAIL.n138 VTAIL.n108 756.745
R861 VTAIL.n265 VTAIL.n264 585
R862 VTAIL.n267 VTAIL.n266 585
R863 VTAIL.n260 VTAIL.n259 585
R864 VTAIL.n273 VTAIL.n272 585
R865 VTAIL.n275 VTAIL.n274 585
R866 VTAIL.n256 VTAIL.n255 585
R867 VTAIL.n281 VTAIL.n280 585
R868 VTAIL.n283 VTAIL.n282 585
R869 VTAIL.n13 VTAIL.n12 585
R870 VTAIL.n15 VTAIL.n14 585
R871 VTAIL.n8 VTAIL.n7 585
R872 VTAIL.n21 VTAIL.n20 585
R873 VTAIL.n23 VTAIL.n22 585
R874 VTAIL.n4 VTAIL.n3 585
R875 VTAIL.n29 VTAIL.n28 585
R876 VTAIL.n31 VTAIL.n30 585
R877 VTAIL.n49 VTAIL.n48 585
R878 VTAIL.n51 VTAIL.n50 585
R879 VTAIL.n44 VTAIL.n43 585
R880 VTAIL.n57 VTAIL.n56 585
R881 VTAIL.n59 VTAIL.n58 585
R882 VTAIL.n40 VTAIL.n39 585
R883 VTAIL.n65 VTAIL.n64 585
R884 VTAIL.n67 VTAIL.n66 585
R885 VTAIL.n85 VTAIL.n84 585
R886 VTAIL.n87 VTAIL.n86 585
R887 VTAIL.n80 VTAIL.n79 585
R888 VTAIL.n93 VTAIL.n92 585
R889 VTAIL.n95 VTAIL.n94 585
R890 VTAIL.n76 VTAIL.n75 585
R891 VTAIL.n101 VTAIL.n100 585
R892 VTAIL.n103 VTAIL.n102 585
R893 VTAIL.n247 VTAIL.n246 585
R894 VTAIL.n245 VTAIL.n244 585
R895 VTAIL.n220 VTAIL.n219 585
R896 VTAIL.n239 VTAIL.n238 585
R897 VTAIL.n237 VTAIL.n236 585
R898 VTAIL.n224 VTAIL.n223 585
R899 VTAIL.n231 VTAIL.n230 585
R900 VTAIL.n229 VTAIL.n228 585
R901 VTAIL.n211 VTAIL.n210 585
R902 VTAIL.n209 VTAIL.n208 585
R903 VTAIL.n184 VTAIL.n183 585
R904 VTAIL.n203 VTAIL.n202 585
R905 VTAIL.n201 VTAIL.n200 585
R906 VTAIL.n188 VTAIL.n187 585
R907 VTAIL.n195 VTAIL.n194 585
R908 VTAIL.n193 VTAIL.n192 585
R909 VTAIL.n175 VTAIL.n174 585
R910 VTAIL.n173 VTAIL.n172 585
R911 VTAIL.n148 VTAIL.n147 585
R912 VTAIL.n167 VTAIL.n166 585
R913 VTAIL.n165 VTAIL.n164 585
R914 VTAIL.n152 VTAIL.n151 585
R915 VTAIL.n159 VTAIL.n158 585
R916 VTAIL.n157 VTAIL.n156 585
R917 VTAIL.n139 VTAIL.n138 585
R918 VTAIL.n137 VTAIL.n136 585
R919 VTAIL.n112 VTAIL.n111 585
R920 VTAIL.n131 VTAIL.n130 585
R921 VTAIL.n129 VTAIL.n128 585
R922 VTAIL.n116 VTAIL.n115 585
R923 VTAIL.n123 VTAIL.n122 585
R924 VTAIL.n121 VTAIL.n120 585
R925 VTAIL.n263 VTAIL.t4 327.514
R926 VTAIL.n11 VTAIL.t7 327.514
R927 VTAIL.n47 VTAIL.t3 327.514
R928 VTAIL.n83 VTAIL.t0 327.514
R929 VTAIL.n227 VTAIL.t1 327.514
R930 VTAIL.n191 VTAIL.t2 327.514
R931 VTAIL.n155 VTAIL.t5 327.514
R932 VTAIL.n119 VTAIL.t6 327.514
R933 VTAIL.n266 VTAIL.n265 171.744
R934 VTAIL.n266 VTAIL.n259 171.744
R935 VTAIL.n273 VTAIL.n259 171.744
R936 VTAIL.n274 VTAIL.n273 171.744
R937 VTAIL.n274 VTAIL.n255 171.744
R938 VTAIL.n281 VTAIL.n255 171.744
R939 VTAIL.n282 VTAIL.n281 171.744
R940 VTAIL.n14 VTAIL.n13 171.744
R941 VTAIL.n14 VTAIL.n7 171.744
R942 VTAIL.n21 VTAIL.n7 171.744
R943 VTAIL.n22 VTAIL.n21 171.744
R944 VTAIL.n22 VTAIL.n3 171.744
R945 VTAIL.n29 VTAIL.n3 171.744
R946 VTAIL.n30 VTAIL.n29 171.744
R947 VTAIL.n50 VTAIL.n49 171.744
R948 VTAIL.n50 VTAIL.n43 171.744
R949 VTAIL.n57 VTAIL.n43 171.744
R950 VTAIL.n58 VTAIL.n57 171.744
R951 VTAIL.n58 VTAIL.n39 171.744
R952 VTAIL.n65 VTAIL.n39 171.744
R953 VTAIL.n66 VTAIL.n65 171.744
R954 VTAIL.n86 VTAIL.n85 171.744
R955 VTAIL.n86 VTAIL.n79 171.744
R956 VTAIL.n93 VTAIL.n79 171.744
R957 VTAIL.n94 VTAIL.n93 171.744
R958 VTAIL.n94 VTAIL.n75 171.744
R959 VTAIL.n101 VTAIL.n75 171.744
R960 VTAIL.n102 VTAIL.n101 171.744
R961 VTAIL.n246 VTAIL.n245 171.744
R962 VTAIL.n245 VTAIL.n219 171.744
R963 VTAIL.n238 VTAIL.n219 171.744
R964 VTAIL.n238 VTAIL.n237 171.744
R965 VTAIL.n237 VTAIL.n223 171.744
R966 VTAIL.n230 VTAIL.n223 171.744
R967 VTAIL.n230 VTAIL.n229 171.744
R968 VTAIL.n210 VTAIL.n209 171.744
R969 VTAIL.n209 VTAIL.n183 171.744
R970 VTAIL.n202 VTAIL.n183 171.744
R971 VTAIL.n202 VTAIL.n201 171.744
R972 VTAIL.n201 VTAIL.n187 171.744
R973 VTAIL.n194 VTAIL.n187 171.744
R974 VTAIL.n194 VTAIL.n193 171.744
R975 VTAIL.n174 VTAIL.n173 171.744
R976 VTAIL.n173 VTAIL.n147 171.744
R977 VTAIL.n166 VTAIL.n147 171.744
R978 VTAIL.n166 VTAIL.n165 171.744
R979 VTAIL.n165 VTAIL.n151 171.744
R980 VTAIL.n158 VTAIL.n151 171.744
R981 VTAIL.n158 VTAIL.n157 171.744
R982 VTAIL.n138 VTAIL.n137 171.744
R983 VTAIL.n137 VTAIL.n111 171.744
R984 VTAIL.n130 VTAIL.n111 171.744
R985 VTAIL.n130 VTAIL.n129 171.744
R986 VTAIL.n129 VTAIL.n115 171.744
R987 VTAIL.n122 VTAIL.n115 171.744
R988 VTAIL.n122 VTAIL.n121 171.744
R989 VTAIL.n265 VTAIL.t4 85.8723
R990 VTAIL.n13 VTAIL.t7 85.8723
R991 VTAIL.n49 VTAIL.t3 85.8723
R992 VTAIL.n85 VTAIL.t0 85.8723
R993 VTAIL.n229 VTAIL.t1 85.8723
R994 VTAIL.n193 VTAIL.t2 85.8723
R995 VTAIL.n157 VTAIL.t5 85.8723
R996 VTAIL.n121 VTAIL.t6 85.8723
R997 VTAIL.n287 VTAIL.n286 31.7975
R998 VTAIL.n35 VTAIL.n34 31.7975
R999 VTAIL.n71 VTAIL.n70 31.7975
R1000 VTAIL.n107 VTAIL.n106 31.7975
R1001 VTAIL.n251 VTAIL.n250 31.7975
R1002 VTAIL.n215 VTAIL.n214 31.7975
R1003 VTAIL.n179 VTAIL.n178 31.7975
R1004 VTAIL.n143 VTAIL.n142 31.7975
R1005 VTAIL.n287 VTAIL.n251 20.9703
R1006 VTAIL.n143 VTAIL.n107 20.9703
R1007 VTAIL.n264 VTAIL.n263 16.3884
R1008 VTAIL.n12 VTAIL.n11 16.3884
R1009 VTAIL.n48 VTAIL.n47 16.3884
R1010 VTAIL.n84 VTAIL.n83 16.3884
R1011 VTAIL.n228 VTAIL.n227 16.3884
R1012 VTAIL.n192 VTAIL.n191 16.3884
R1013 VTAIL.n156 VTAIL.n155 16.3884
R1014 VTAIL.n120 VTAIL.n119 16.3884
R1015 VTAIL.n267 VTAIL.n262 12.8005
R1016 VTAIL.n15 VTAIL.n10 12.8005
R1017 VTAIL.n51 VTAIL.n46 12.8005
R1018 VTAIL.n87 VTAIL.n82 12.8005
R1019 VTAIL.n231 VTAIL.n226 12.8005
R1020 VTAIL.n195 VTAIL.n190 12.8005
R1021 VTAIL.n159 VTAIL.n154 12.8005
R1022 VTAIL.n123 VTAIL.n118 12.8005
R1023 VTAIL.n268 VTAIL.n260 12.0247
R1024 VTAIL.n16 VTAIL.n8 12.0247
R1025 VTAIL.n52 VTAIL.n44 12.0247
R1026 VTAIL.n88 VTAIL.n80 12.0247
R1027 VTAIL.n232 VTAIL.n224 12.0247
R1028 VTAIL.n196 VTAIL.n188 12.0247
R1029 VTAIL.n160 VTAIL.n152 12.0247
R1030 VTAIL.n124 VTAIL.n116 12.0247
R1031 VTAIL.n272 VTAIL.n271 11.249
R1032 VTAIL.n20 VTAIL.n19 11.249
R1033 VTAIL.n56 VTAIL.n55 11.249
R1034 VTAIL.n92 VTAIL.n91 11.249
R1035 VTAIL.n236 VTAIL.n235 11.249
R1036 VTAIL.n200 VTAIL.n199 11.249
R1037 VTAIL.n164 VTAIL.n163 11.249
R1038 VTAIL.n128 VTAIL.n127 11.249
R1039 VTAIL.n275 VTAIL.n258 10.4732
R1040 VTAIL.n23 VTAIL.n6 10.4732
R1041 VTAIL.n59 VTAIL.n42 10.4732
R1042 VTAIL.n95 VTAIL.n78 10.4732
R1043 VTAIL.n239 VTAIL.n222 10.4732
R1044 VTAIL.n203 VTAIL.n186 10.4732
R1045 VTAIL.n167 VTAIL.n150 10.4732
R1046 VTAIL.n131 VTAIL.n114 10.4732
R1047 VTAIL.n276 VTAIL.n256 9.69747
R1048 VTAIL.n24 VTAIL.n4 9.69747
R1049 VTAIL.n60 VTAIL.n40 9.69747
R1050 VTAIL.n96 VTAIL.n76 9.69747
R1051 VTAIL.n240 VTAIL.n220 9.69747
R1052 VTAIL.n204 VTAIL.n184 9.69747
R1053 VTAIL.n168 VTAIL.n148 9.69747
R1054 VTAIL.n132 VTAIL.n112 9.69747
R1055 VTAIL.n286 VTAIL.n285 9.45567
R1056 VTAIL.n34 VTAIL.n33 9.45567
R1057 VTAIL.n70 VTAIL.n69 9.45567
R1058 VTAIL.n106 VTAIL.n105 9.45567
R1059 VTAIL.n250 VTAIL.n249 9.45567
R1060 VTAIL.n214 VTAIL.n213 9.45567
R1061 VTAIL.n178 VTAIL.n177 9.45567
R1062 VTAIL.n142 VTAIL.n141 9.45567
R1063 VTAIL.n254 VTAIL.n253 9.3005
R1064 VTAIL.n279 VTAIL.n278 9.3005
R1065 VTAIL.n277 VTAIL.n276 9.3005
R1066 VTAIL.n258 VTAIL.n257 9.3005
R1067 VTAIL.n271 VTAIL.n270 9.3005
R1068 VTAIL.n269 VTAIL.n268 9.3005
R1069 VTAIL.n262 VTAIL.n261 9.3005
R1070 VTAIL.n285 VTAIL.n284 9.3005
R1071 VTAIL.n2 VTAIL.n1 9.3005
R1072 VTAIL.n27 VTAIL.n26 9.3005
R1073 VTAIL.n25 VTAIL.n24 9.3005
R1074 VTAIL.n6 VTAIL.n5 9.3005
R1075 VTAIL.n19 VTAIL.n18 9.3005
R1076 VTAIL.n17 VTAIL.n16 9.3005
R1077 VTAIL.n10 VTAIL.n9 9.3005
R1078 VTAIL.n33 VTAIL.n32 9.3005
R1079 VTAIL.n38 VTAIL.n37 9.3005
R1080 VTAIL.n63 VTAIL.n62 9.3005
R1081 VTAIL.n61 VTAIL.n60 9.3005
R1082 VTAIL.n42 VTAIL.n41 9.3005
R1083 VTAIL.n55 VTAIL.n54 9.3005
R1084 VTAIL.n53 VTAIL.n52 9.3005
R1085 VTAIL.n46 VTAIL.n45 9.3005
R1086 VTAIL.n69 VTAIL.n68 9.3005
R1087 VTAIL.n74 VTAIL.n73 9.3005
R1088 VTAIL.n99 VTAIL.n98 9.3005
R1089 VTAIL.n97 VTAIL.n96 9.3005
R1090 VTAIL.n78 VTAIL.n77 9.3005
R1091 VTAIL.n91 VTAIL.n90 9.3005
R1092 VTAIL.n89 VTAIL.n88 9.3005
R1093 VTAIL.n82 VTAIL.n81 9.3005
R1094 VTAIL.n105 VTAIL.n104 9.3005
R1095 VTAIL.n249 VTAIL.n248 9.3005
R1096 VTAIL.n218 VTAIL.n217 9.3005
R1097 VTAIL.n243 VTAIL.n242 9.3005
R1098 VTAIL.n241 VTAIL.n240 9.3005
R1099 VTAIL.n222 VTAIL.n221 9.3005
R1100 VTAIL.n235 VTAIL.n234 9.3005
R1101 VTAIL.n233 VTAIL.n232 9.3005
R1102 VTAIL.n226 VTAIL.n225 9.3005
R1103 VTAIL.n213 VTAIL.n212 9.3005
R1104 VTAIL.n182 VTAIL.n181 9.3005
R1105 VTAIL.n207 VTAIL.n206 9.3005
R1106 VTAIL.n205 VTAIL.n204 9.3005
R1107 VTAIL.n186 VTAIL.n185 9.3005
R1108 VTAIL.n199 VTAIL.n198 9.3005
R1109 VTAIL.n197 VTAIL.n196 9.3005
R1110 VTAIL.n190 VTAIL.n189 9.3005
R1111 VTAIL.n177 VTAIL.n176 9.3005
R1112 VTAIL.n146 VTAIL.n145 9.3005
R1113 VTAIL.n171 VTAIL.n170 9.3005
R1114 VTAIL.n169 VTAIL.n168 9.3005
R1115 VTAIL.n150 VTAIL.n149 9.3005
R1116 VTAIL.n163 VTAIL.n162 9.3005
R1117 VTAIL.n161 VTAIL.n160 9.3005
R1118 VTAIL.n154 VTAIL.n153 9.3005
R1119 VTAIL.n141 VTAIL.n140 9.3005
R1120 VTAIL.n110 VTAIL.n109 9.3005
R1121 VTAIL.n135 VTAIL.n134 9.3005
R1122 VTAIL.n133 VTAIL.n132 9.3005
R1123 VTAIL.n114 VTAIL.n113 9.3005
R1124 VTAIL.n127 VTAIL.n126 9.3005
R1125 VTAIL.n125 VTAIL.n124 9.3005
R1126 VTAIL.n118 VTAIL.n117 9.3005
R1127 VTAIL.n280 VTAIL.n279 8.92171
R1128 VTAIL.n28 VTAIL.n27 8.92171
R1129 VTAIL.n64 VTAIL.n63 8.92171
R1130 VTAIL.n100 VTAIL.n99 8.92171
R1131 VTAIL.n244 VTAIL.n243 8.92171
R1132 VTAIL.n208 VTAIL.n207 8.92171
R1133 VTAIL.n172 VTAIL.n171 8.92171
R1134 VTAIL.n136 VTAIL.n135 8.92171
R1135 VTAIL.n283 VTAIL.n254 8.14595
R1136 VTAIL.n31 VTAIL.n2 8.14595
R1137 VTAIL.n67 VTAIL.n38 8.14595
R1138 VTAIL.n103 VTAIL.n74 8.14595
R1139 VTAIL.n247 VTAIL.n218 8.14595
R1140 VTAIL.n211 VTAIL.n182 8.14595
R1141 VTAIL.n175 VTAIL.n146 8.14595
R1142 VTAIL.n139 VTAIL.n110 8.14595
R1143 VTAIL.n284 VTAIL.n252 7.3702
R1144 VTAIL.n32 VTAIL.n0 7.3702
R1145 VTAIL.n68 VTAIL.n36 7.3702
R1146 VTAIL.n104 VTAIL.n72 7.3702
R1147 VTAIL.n248 VTAIL.n216 7.3702
R1148 VTAIL.n212 VTAIL.n180 7.3702
R1149 VTAIL.n176 VTAIL.n144 7.3702
R1150 VTAIL.n140 VTAIL.n108 7.3702
R1151 VTAIL.n286 VTAIL.n252 6.59444
R1152 VTAIL.n34 VTAIL.n0 6.59444
R1153 VTAIL.n70 VTAIL.n36 6.59444
R1154 VTAIL.n106 VTAIL.n72 6.59444
R1155 VTAIL.n250 VTAIL.n216 6.59444
R1156 VTAIL.n214 VTAIL.n180 6.59444
R1157 VTAIL.n178 VTAIL.n144 6.59444
R1158 VTAIL.n142 VTAIL.n108 6.59444
R1159 VTAIL.n284 VTAIL.n283 5.81868
R1160 VTAIL.n32 VTAIL.n31 5.81868
R1161 VTAIL.n68 VTAIL.n67 5.81868
R1162 VTAIL.n104 VTAIL.n103 5.81868
R1163 VTAIL.n248 VTAIL.n247 5.81868
R1164 VTAIL.n212 VTAIL.n211 5.81868
R1165 VTAIL.n176 VTAIL.n175 5.81868
R1166 VTAIL.n140 VTAIL.n139 5.81868
R1167 VTAIL.n280 VTAIL.n254 5.04292
R1168 VTAIL.n28 VTAIL.n2 5.04292
R1169 VTAIL.n64 VTAIL.n38 5.04292
R1170 VTAIL.n100 VTAIL.n74 5.04292
R1171 VTAIL.n244 VTAIL.n218 5.04292
R1172 VTAIL.n208 VTAIL.n182 5.04292
R1173 VTAIL.n172 VTAIL.n146 5.04292
R1174 VTAIL.n136 VTAIL.n110 5.04292
R1175 VTAIL.n279 VTAIL.n256 4.26717
R1176 VTAIL.n27 VTAIL.n4 4.26717
R1177 VTAIL.n63 VTAIL.n40 4.26717
R1178 VTAIL.n99 VTAIL.n76 4.26717
R1179 VTAIL.n243 VTAIL.n220 4.26717
R1180 VTAIL.n207 VTAIL.n184 4.26717
R1181 VTAIL.n171 VTAIL.n148 4.26717
R1182 VTAIL.n135 VTAIL.n112 4.26717
R1183 VTAIL.n263 VTAIL.n261 3.71088
R1184 VTAIL.n11 VTAIL.n9 3.71088
R1185 VTAIL.n47 VTAIL.n45 3.71088
R1186 VTAIL.n83 VTAIL.n81 3.71088
R1187 VTAIL.n227 VTAIL.n225 3.71088
R1188 VTAIL.n191 VTAIL.n189 3.71088
R1189 VTAIL.n155 VTAIL.n153 3.71088
R1190 VTAIL.n119 VTAIL.n117 3.71088
R1191 VTAIL.n276 VTAIL.n275 3.49141
R1192 VTAIL.n24 VTAIL.n23 3.49141
R1193 VTAIL.n60 VTAIL.n59 3.49141
R1194 VTAIL.n96 VTAIL.n95 3.49141
R1195 VTAIL.n240 VTAIL.n239 3.49141
R1196 VTAIL.n204 VTAIL.n203 3.49141
R1197 VTAIL.n168 VTAIL.n167 3.49141
R1198 VTAIL.n132 VTAIL.n131 3.49141
R1199 VTAIL.n179 VTAIL.n143 2.82809
R1200 VTAIL.n251 VTAIL.n215 2.82809
R1201 VTAIL.n107 VTAIL.n71 2.82809
R1202 VTAIL.n272 VTAIL.n258 2.71565
R1203 VTAIL.n20 VTAIL.n6 2.71565
R1204 VTAIL.n56 VTAIL.n42 2.71565
R1205 VTAIL.n92 VTAIL.n78 2.71565
R1206 VTAIL.n236 VTAIL.n222 2.71565
R1207 VTAIL.n200 VTAIL.n186 2.71565
R1208 VTAIL.n164 VTAIL.n150 2.71565
R1209 VTAIL.n128 VTAIL.n114 2.71565
R1210 VTAIL.n271 VTAIL.n260 1.93989
R1211 VTAIL.n19 VTAIL.n8 1.93989
R1212 VTAIL.n55 VTAIL.n44 1.93989
R1213 VTAIL.n91 VTAIL.n80 1.93989
R1214 VTAIL.n235 VTAIL.n224 1.93989
R1215 VTAIL.n199 VTAIL.n188 1.93989
R1216 VTAIL.n163 VTAIL.n152 1.93989
R1217 VTAIL.n127 VTAIL.n116 1.93989
R1218 VTAIL VTAIL.n35 1.47248
R1219 VTAIL VTAIL.n287 1.3561
R1220 VTAIL.n268 VTAIL.n267 1.16414
R1221 VTAIL.n16 VTAIL.n15 1.16414
R1222 VTAIL.n52 VTAIL.n51 1.16414
R1223 VTAIL.n88 VTAIL.n87 1.16414
R1224 VTAIL.n232 VTAIL.n231 1.16414
R1225 VTAIL.n196 VTAIL.n195 1.16414
R1226 VTAIL.n160 VTAIL.n159 1.16414
R1227 VTAIL.n124 VTAIL.n123 1.16414
R1228 VTAIL.n215 VTAIL.n179 0.470328
R1229 VTAIL.n71 VTAIL.n35 0.470328
R1230 VTAIL.n264 VTAIL.n262 0.388379
R1231 VTAIL.n12 VTAIL.n10 0.388379
R1232 VTAIL.n48 VTAIL.n46 0.388379
R1233 VTAIL.n84 VTAIL.n82 0.388379
R1234 VTAIL.n228 VTAIL.n226 0.388379
R1235 VTAIL.n192 VTAIL.n190 0.388379
R1236 VTAIL.n156 VTAIL.n154 0.388379
R1237 VTAIL.n120 VTAIL.n118 0.388379
R1238 VTAIL.n269 VTAIL.n261 0.155672
R1239 VTAIL.n270 VTAIL.n269 0.155672
R1240 VTAIL.n270 VTAIL.n257 0.155672
R1241 VTAIL.n277 VTAIL.n257 0.155672
R1242 VTAIL.n278 VTAIL.n277 0.155672
R1243 VTAIL.n278 VTAIL.n253 0.155672
R1244 VTAIL.n285 VTAIL.n253 0.155672
R1245 VTAIL.n17 VTAIL.n9 0.155672
R1246 VTAIL.n18 VTAIL.n17 0.155672
R1247 VTAIL.n18 VTAIL.n5 0.155672
R1248 VTAIL.n25 VTAIL.n5 0.155672
R1249 VTAIL.n26 VTAIL.n25 0.155672
R1250 VTAIL.n26 VTAIL.n1 0.155672
R1251 VTAIL.n33 VTAIL.n1 0.155672
R1252 VTAIL.n53 VTAIL.n45 0.155672
R1253 VTAIL.n54 VTAIL.n53 0.155672
R1254 VTAIL.n54 VTAIL.n41 0.155672
R1255 VTAIL.n61 VTAIL.n41 0.155672
R1256 VTAIL.n62 VTAIL.n61 0.155672
R1257 VTAIL.n62 VTAIL.n37 0.155672
R1258 VTAIL.n69 VTAIL.n37 0.155672
R1259 VTAIL.n89 VTAIL.n81 0.155672
R1260 VTAIL.n90 VTAIL.n89 0.155672
R1261 VTAIL.n90 VTAIL.n77 0.155672
R1262 VTAIL.n97 VTAIL.n77 0.155672
R1263 VTAIL.n98 VTAIL.n97 0.155672
R1264 VTAIL.n98 VTAIL.n73 0.155672
R1265 VTAIL.n105 VTAIL.n73 0.155672
R1266 VTAIL.n249 VTAIL.n217 0.155672
R1267 VTAIL.n242 VTAIL.n217 0.155672
R1268 VTAIL.n242 VTAIL.n241 0.155672
R1269 VTAIL.n241 VTAIL.n221 0.155672
R1270 VTAIL.n234 VTAIL.n221 0.155672
R1271 VTAIL.n234 VTAIL.n233 0.155672
R1272 VTAIL.n233 VTAIL.n225 0.155672
R1273 VTAIL.n213 VTAIL.n181 0.155672
R1274 VTAIL.n206 VTAIL.n181 0.155672
R1275 VTAIL.n206 VTAIL.n205 0.155672
R1276 VTAIL.n205 VTAIL.n185 0.155672
R1277 VTAIL.n198 VTAIL.n185 0.155672
R1278 VTAIL.n198 VTAIL.n197 0.155672
R1279 VTAIL.n197 VTAIL.n189 0.155672
R1280 VTAIL.n177 VTAIL.n145 0.155672
R1281 VTAIL.n170 VTAIL.n145 0.155672
R1282 VTAIL.n170 VTAIL.n169 0.155672
R1283 VTAIL.n169 VTAIL.n149 0.155672
R1284 VTAIL.n162 VTAIL.n149 0.155672
R1285 VTAIL.n162 VTAIL.n161 0.155672
R1286 VTAIL.n161 VTAIL.n153 0.155672
R1287 VTAIL.n141 VTAIL.n109 0.155672
R1288 VTAIL.n134 VTAIL.n109 0.155672
R1289 VTAIL.n134 VTAIL.n133 0.155672
R1290 VTAIL.n133 VTAIL.n113 0.155672
R1291 VTAIL.n126 VTAIL.n113 0.155672
R1292 VTAIL.n126 VTAIL.n125 0.155672
R1293 VTAIL.n125 VTAIL.n117 0.155672
R1294 VDD2.n2 VDD2.n0 125.984
R1295 VDD2.n2 VDD2.n1 88.0109
R1296 VDD2.n1 VDD2.t2 4.85199
R1297 VDD2.n1 VDD2.t3 4.85199
R1298 VDD2.n0 VDD2.t1 4.85199
R1299 VDD2.n0 VDD2.t0 4.85199
R1300 VDD2 VDD2.n2 0.0586897
R1301 VP.n15 VP.n14 161.3
R1302 VP.n13 VP.n1 161.3
R1303 VP.n12 VP.n11 161.3
R1304 VP.n10 VP.n2 161.3
R1305 VP.n9 VP.n8 161.3
R1306 VP.n7 VP.n3 161.3
R1307 VP.n4 VP.t2 89.1885
R1308 VP.n4 VP.t1 88.2078
R1309 VP.n6 VP.n5 71.0639
R1310 VP.n16 VP.n0 71.0639
R1311 VP.n12 VP.n2 56.5617
R1312 VP.n6 VP.t3 54.7361
R1313 VP.n0 VP.t0 54.7361
R1314 VP.n5 VP.n4 46.4656
R1315 VP.n8 VP.n7 24.5923
R1316 VP.n8 VP.n2 24.5923
R1317 VP.n13 VP.n12 24.5923
R1318 VP.n14 VP.n13 24.5923
R1319 VP.n7 VP.n6 19.1821
R1320 VP.n14 VP.n0 19.1821
R1321 VP.n5 VP.n3 0.354861
R1322 VP.n16 VP.n15 0.354861
R1323 VP VP.n16 0.267071
R1324 VP.n9 VP.n3 0.189894
R1325 VP.n10 VP.n9 0.189894
R1326 VP.n11 VP.n10 0.189894
R1327 VP.n11 VP.n1 0.189894
R1328 VP.n15 VP.n1 0.189894
R1329 VDD1 VDD1.n1 126.51
R1330 VDD1 VDD1.n0 88.0691
R1331 VDD1.n0 VDD1.t1 4.85199
R1332 VDD1.n0 VDD1.t2 4.85199
R1333 VDD1.n1 VDD1.t0 4.85199
R1334 VDD1.n1 VDD1.t3 4.85199
C0 w_n2938_n2308# VP 5.32171f
C1 VTAIL B 3.32082f
C2 VN VP 5.46084f
C3 w_n2938_n2308# VDD2 1.44369f
C4 VN VDD2 2.85069f
C5 VDD1 VP 3.11712f
C6 VDD1 VDD2 1.11047f
C7 VN w_n2938_n2308# 4.94313f
C8 VP VTAIL 3.19211f
C9 VP B 1.7449f
C10 VTAIL VDD2 4.33188f
C11 VDD1 w_n2938_n2308# 1.37981f
C12 VDD2 B 1.23849f
C13 VDD1 VN 0.149791f
C14 w_n2938_n2308# VTAIL 2.80417f
C15 w_n2938_n2308# B 8.196031f
C16 VN VTAIL 3.17801f
C17 VN B 1.11504f
C18 VDD1 VTAIL 4.27532f
C19 VP VDD2 0.417051f
C20 VDD1 B 1.18053f
C21 VDD2 VSUBS 0.877988f
C22 VDD1 VSUBS 5.28826f
C23 VTAIL VSUBS 0.754112f
C24 VN VSUBS 5.4992f
C25 VP VSUBS 2.1551f
C26 B VSUBS 4.130918f
C27 w_n2938_n2308# VSUBS 84.438095f
C28 VDD1.t1 VSUBS 0.148886f
C29 VDD1.t2 VSUBS 0.148886f
C30 VDD1.n0 VSUBS 1.01576f
C31 VDD1.t0 VSUBS 0.148886f
C32 VDD1.t3 VSUBS 0.148886f
C33 VDD1.n1 VSUBS 1.53468f
C34 VP.t0 VSUBS 2.05201f
C35 VP.n0 VSUBS 0.903908f
C36 VP.n1 VSUBS 0.038986f
C37 VP.n2 VSUBS 0.056672f
C38 VP.n3 VSUBS 0.062912f
C39 VP.t3 VSUBS 2.05201f
C40 VP.t2 VSUBS 2.44872f
C41 VP.t1 VSUBS 2.43766f
C42 VP.n4 VSUBS 3.5145f
C43 VP.n5 VSUBS 1.96307f
C44 VP.n6 VSUBS 0.903908f
C45 VP.n7 VSUBS 0.064443f
C46 VP.n8 VSUBS 0.072295f
C47 VP.n9 VSUBS 0.038986f
C48 VP.n10 VSUBS 0.038986f
C49 VP.n11 VSUBS 0.038986f
C50 VP.n12 VSUBS 0.056672f
C51 VP.n13 VSUBS 0.072295f
C52 VP.n14 VSUBS 0.064443f
C53 VP.n15 VSUBS 0.062912f
C54 VP.n16 VSUBS 0.081992f
C55 VDD2.t1 VSUBS 0.146924f
C56 VDD2.t0 VSUBS 0.146924f
C57 VDD2.n0 VSUBS 1.49282f
C58 VDD2.t2 VSUBS 0.146924f
C59 VDD2.t3 VSUBS 0.146924f
C60 VDD2.n1 VSUBS 1.00189f
C61 VDD2.n2 VSUBS 3.85878f
C62 VTAIL.n0 VSUBS 0.030141f
C63 VTAIL.n1 VSUBS 0.027325f
C64 VTAIL.n2 VSUBS 0.014683f
C65 VTAIL.n3 VSUBS 0.034706f
C66 VTAIL.n4 VSUBS 0.015547f
C67 VTAIL.n5 VSUBS 0.027325f
C68 VTAIL.n6 VSUBS 0.014683f
C69 VTAIL.n7 VSUBS 0.034706f
C70 VTAIL.n8 VSUBS 0.015547f
C71 VTAIL.n9 VSUBS 0.714202f
C72 VTAIL.n10 VSUBS 0.014683f
C73 VTAIL.t7 VSUBS 0.074218f
C74 VTAIL.n11 VSUBS 0.126188f
C75 VTAIL.n12 VSUBS 0.022074f
C76 VTAIL.n13 VSUBS 0.026029f
C77 VTAIL.n14 VSUBS 0.034706f
C78 VTAIL.n15 VSUBS 0.015547f
C79 VTAIL.n16 VSUBS 0.014683f
C80 VTAIL.n17 VSUBS 0.027325f
C81 VTAIL.n18 VSUBS 0.027325f
C82 VTAIL.n19 VSUBS 0.014683f
C83 VTAIL.n20 VSUBS 0.015547f
C84 VTAIL.n21 VSUBS 0.034706f
C85 VTAIL.n22 VSUBS 0.034706f
C86 VTAIL.n23 VSUBS 0.015547f
C87 VTAIL.n24 VSUBS 0.014683f
C88 VTAIL.n25 VSUBS 0.027325f
C89 VTAIL.n26 VSUBS 0.027325f
C90 VTAIL.n27 VSUBS 0.014683f
C91 VTAIL.n28 VSUBS 0.015547f
C92 VTAIL.n29 VSUBS 0.034706f
C93 VTAIL.n30 VSUBS 0.084418f
C94 VTAIL.n31 VSUBS 0.015547f
C95 VTAIL.n32 VSUBS 0.014683f
C96 VTAIL.n33 VSUBS 0.062413f
C97 VTAIL.n34 VSUBS 0.042448f
C98 VTAIL.n35 VSUBS 0.193885f
C99 VTAIL.n36 VSUBS 0.030141f
C100 VTAIL.n37 VSUBS 0.027325f
C101 VTAIL.n38 VSUBS 0.014683f
C102 VTAIL.n39 VSUBS 0.034706f
C103 VTAIL.n40 VSUBS 0.015547f
C104 VTAIL.n41 VSUBS 0.027325f
C105 VTAIL.n42 VSUBS 0.014683f
C106 VTAIL.n43 VSUBS 0.034706f
C107 VTAIL.n44 VSUBS 0.015547f
C108 VTAIL.n45 VSUBS 0.714202f
C109 VTAIL.n46 VSUBS 0.014683f
C110 VTAIL.t3 VSUBS 0.074218f
C111 VTAIL.n47 VSUBS 0.126188f
C112 VTAIL.n48 VSUBS 0.022074f
C113 VTAIL.n49 VSUBS 0.026029f
C114 VTAIL.n50 VSUBS 0.034706f
C115 VTAIL.n51 VSUBS 0.015547f
C116 VTAIL.n52 VSUBS 0.014683f
C117 VTAIL.n53 VSUBS 0.027325f
C118 VTAIL.n54 VSUBS 0.027325f
C119 VTAIL.n55 VSUBS 0.014683f
C120 VTAIL.n56 VSUBS 0.015547f
C121 VTAIL.n57 VSUBS 0.034706f
C122 VTAIL.n58 VSUBS 0.034706f
C123 VTAIL.n59 VSUBS 0.015547f
C124 VTAIL.n60 VSUBS 0.014683f
C125 VTAIL.n61 VSUBS 0.027325f
C126 VTAIL.n62 VSUBS 0.027325f
C127 VTAIL.n63 VSUBS 0.014683f
C128 VTAIL.n64 VSUBS 0.015547f
C129 VTAIL.n65 VSUBS 0.034706f
C130 VTAIL.n66 VSUBS 0.084418f
C131 VTAIL.n67 VSUBS 0.015547f
C132 VTAIL.n68 VSUBS 0.014683f
C133 VTAIL.n69 VSUBS 0.062413f
C134 VTAIL.n70 VSUBS 0.042448f
C135 VTAIL.n71 VSUBS 0.313241f
C136 VTAIL.n72 VSUBS 0.030141f
C137 VTAIL.n73 VSUBS 0.027325f
C138 VTAIL.n74 VSUBS 0.014683f
C139 VTAIL.n75 VSUBS 0.034706f
C140 VTAIL.n76 VSUBS 0.015547f
C141 VTAIL.n77 VSUBS 0.027325f
C142 VTAIL.n78 VSUBS 0.014683f
C143 VTAIL.n79 VSUBS 0.034706f
C144 VTAIL.n80 VSUBS 0.015547f
C145 VTAIL.n81 VSUBS 0.714202f
C146 VTAIL.n82 VSUBS 0.014683f
C147 VTAIL.t0 VSUBS 0.074218f
C148 VTAIL.n83 VSUBS 0.126188f
C149 VTAIL.n84 VSUBS 0.022074f
C150 VTAIL.n85 VSUBS 0.026029f
C151 VTAIL.n86 VSUBS 0.034706f
C152 VTAIL.n87 VSUBS 0.015547f
C153 VTAIL.n88 VSUBS 0.014683f
C154 VTAIL.n89 VSUBS 0.027325f
C155 VTAIL.n90 VSUBS 0.027325f
C156 VTAIL.n91 VSUBS 0.014683f
C157 VTAIL.n92 VSUBS 0.015547f
C158 VTAIL.n93 VSUBS 0.034706f
C159 VTAIL.n94 VSUBS 0.034706f
C160 VTAIL.n95 VSUBS 0.015547f
C161 VTAIL.n96 VSUBS 0.014683f
C162 VTAIL.n97 VSUBS 0.027325f
C163 VTAIL.n98 VSUBS 0.027325f
C164 VTAIL.n99 VSUBS 0.014683f
C165 VTAIL.n100 VSUBS 0.015547f
C166 VTAIL.n101 VSUBS 0.034706f
C167 VTAIL.n102 VSUBS 0.084418f
C168 VTAIL.n103 VSUBS 0.015547f
C169 VTAIL.n104 VSUBS 0.014683f
C170 VTAIL.n105 VSUBS 0.062413f
C171 VTAIL.n106 VSUBS 0.042448f
C172 VTAIL.n107 VSUBS 1.40055f
C173 VTAIL.n108 VSUBS 0.030141f
C174 VTAIL.n109 VSUBS 0.027325f
C175 VTAIL.n110 VSUBS 0.014683f
C176 VTAIL.n111 VSUBS 0.034706f
C177 VTAIL.n112 VSUBS 0.015547f
C178 VTAIL.n113 VSUBS 0.027325f
C179 VTAIL.n114 VSUBS 0.014683f
C180 VTAIL.n115 VSUBS 0.034706f
C181 VTAIL.n116 VSUBS 0.015547f
C182 VTAIL.n117 VSUBS 0.714202f
C183 VTAIL.n118 VSUBS 0.014683f
C184 VTAIL.t6 VSUBS 0.074218f
C185 VTAIL.n119 VSUBS 0.126188f
C186 VTAIL.n120 VSUBS 0.022074f
C187 VTAIL.n121 VSUBS 0.026029f
C188 VTAIL.n122 VSUBS 0.034706f
C189 VTAIL.n123 VSUBS 0.015547f
C190 VTAIL.n124 VSUBS 0.014683f
C191 VTAIL.n125 VSUBS 0.027325f
C192 VTAIL.n126 VSUBS 0.027325f
C193 VTAIL.n127 VSUBS 0.014683f
C194 VTAIL.n128 VSUBS 0.015547f
C195 VTAIL.n129 VSUBS 0.034706f
C196 VTAIL.n130 VSUBS 0.034706f
C197 VTAIL.n131 VSUBS 0.015547f
C198 VTAIL.n132 VSUBS 0.014683f
C199 VTAIL.n133 VSUBS 0.027325f
C200 VTAIL.n134 VSUBS 0.027325f
C201 VTAIL.n135 VSUBS 0.014683f
C202 VTAIL.n136 VSUBS 0.015547f
C203 VTAIL.n137 VSUBS 0.034706f
C204 VTAIL.n138 VSUBS 0.084418f
C205 VTAIL.n139 VSUBS 0.015547f
C206 VTAIL.n140 VSUBS 0.014683f
C207 VTAIL.n141 VSUBS 0.062413f
C208 VTAIL.n142 VSUBS 0.042448f
C209 VTAIL.n143 VSUBS 1.40055f
C210 VTAIL.n144 VSUBS 0.030141f
C211 VTAIL.n145 VSUBS 0.027325f
C212 VTAIL.n146 VSUBS 0.014683f
C213 VTAIL.n147 VSUBS 0.034706f
C214 VTAIL.n148 VSUBS 0.015547f
C215 VTAIL.n149 VSUBS 0.027325f
C216 VTAIL.n150 VSUBS 0.014683f
C217 VTAIL.n151 VSUBS 0.034706f
C218 VTAIL.n152 VSUBS 0.015547f
C219 VTAIL.n153 VSUBS 0.714202f
C220 VTAIL.n154 VSUBS 0.014683f
C221 VTAIL.t5 VSUBS 0.074218f
C222 VTAIL.n155 VSUBS 0.126188f
C223 VTAIL.n156 VSUBS 0.022074f
C224 VTAIL.n157 VSUBS 0.026029f
C225 VTAIL.n158 VSUBS 0.034706f
C226 VTAIL.n159 VSUBS 0.015547f
C227 VTAIL.n160 VSUBS 0.014683f
C228 VTAIL.n161 VSUBS 0.027325f
C229 VTAIL.n162 VSUBS 0.027325f
C230 VTAIL.n163 VSUBS 0.014683f
C231 VTAIL.n164 VSUBS 0.015547f
C232 VTAIL.n165 VSUBS 0.034706f
C233 VTAIL.n166 VSUBS 0.034706f
C234 VTAIL.n167 VSUBS 0.015547f
C235 VTAIL.n168 VSUBS 0.014683f
C236 VTAIL.n169 VSUBS 0.027325f
C237 VTAIL.n170 VSUBS 0.027325f
C238 VTAIL.n171 VSUBS 0.014683f
C239 VTAIL.n172 VSUBS 0.015547f
C240 VTAIL.n173 VSUBS 0.034706f
C241 VTAIL.n174 VSUBS 0.084418f
C242 VTAIL.n175 VSUBS 0.015547f
C243 VTAIL.n176 VSUBS 0.014683f
C244 VTAIL.n177 VSUBS 0.062413f
C245 VTAIL.n178 VSUBS 0.042448f
C246 VTAIL.n179 VSUBS 0.313241f
C247 VTAIL.n180 VSUBS 0.030141f
C248 VTAIL.n181 VSUBS 0.027325f
C249 VTAIL.n182 VSUBS 0.014683f
C250 VTAIL.n183 VSUBS 0.034706f
C251 VTAIL.n184 VSUBS 0.015547f
C252 VTAIL.n185 VSUBS 0.027325f
C253 VTAIL.n186 VSUBS 0.014683f
C254 VTAIL.n187 VSUBS 0.034706f
C255 VTAIL.n188 VSUBS 0.015547f
C256 VTAIL.n189 VSUBS 0.714202f
C257 VTAIL.n190 VSUBS 0.014683f
C258 VTAIL.t2 VSUBS 0.074218f
C259 VTAIL.n191 VSUBS 0.126188f
C260 VTAIL.n192 VSUBS 0.022074f
C261 VTAIL.n193 VSUBS 0.026029f
C262 VTAIL.n194 VSUBS 0.034706f
C263 VTAIL.n195 VSUBS 0.015547f
C264 VTAIL.n196 VSUBS 0.014683f
C265 VTAIL.n197 VSUBS 0.027325f
C266 VTAIL.n198 VSUBS 0.027325f
C267 VTAIL.n199 VSUBS 0.014683f
C268 VTAIL.n200 VSUBS 0.015547f
C269 VTAIL.n201 VSUBS 0.034706f
C270 VTAIL.n202 VSUBS 0.034706f
C271 VTAIL.n203 VSUBS 0.015547f
C272 VTAIL.n204 VSUBS 0.014683f
C273 VTAIL.n205 VSUBS 0.027325f
C274 VTAIL.n206 VSUBS 0.027325f
C275 VTAIL.n207 VSUBS 0.014683f
C276 VTAIL.n208 VSUBS 0.015547f
C277 VTAIL.n209 VSUBS 0.034706f
C278 VTAIL.n210 VSUBS 0.084418f
C279 VTAIL.n211 VSUBS 0.015547f
C280 VTAIL.n212 VSUBS 0.014683f
C281 VTAIL.n213 VSUBS 0.062413f
C282 VTAIL.n214 VSUBS 0.042448f
C283 VTAIL.n215 VSUBS 0.313241f
C284 VTAIL.n216 VSUBS 0.030141f
C285 VTAIL.n217 VSUBS 0.027325f
C286 VTAIL.n218 VSUBS 0.014683f
C287 VTAIL.n219 VSUBS 0.034706f
C288 VTAIL.n220 VSUBS 0.015547f
C289 VTAIL.n221 VSUBS 0.027325f
C290 VTAIL.n222 VSUBS 0.014683f
C291 VTAIL.n223 VSUBS 0.034706f
C292 VTAIL.n224 VSUBS 0.015547f
C293 VTAIL.n225 VSUBS 0.714202f
C294 VTAIL.n226 VSUBS 0.014683f
C295 VTAIL.t1 VSUBS 0.074218f
C296 VTAIL.n227 VSUBS 0.126188f
C297 VTAIL.n228 VSUBS 0.022074f
C298 VTAIL.n229 VSUBS 0.026029f
C299 VTAIL.n230 VSUBS 0.034706f
C300 VTAIL.n231 VSUBS 0.015547f
C301 VTAIL.n232 VSUBS 0.014683f
C302 VTAIL.n233 VSUBS 0.027325f
C303 VTAIL.n234 VSUBS 0.027325f
C304 VTAIL.n235 VSUBS 0.014683f
C305 VTAIL.n236 VSUBS 0.015547f
C306 VTAIL.n237 VSUBS 0.034706f
C307 VTAIL.n238 VSUBS 0.034706f
C308 VTAIL.n239 VSUBS 0.015547f
C309 VTAIL.n240 VSUBS 0.014683f
C310 VTAIL.n241 VSUBS 0.027325f
C311 VTAIL.n242 VSUBS 0.027325f
C312 VTAIL.n243 VSUBS 0.014683f
C313 VTAIL.n244 VSUBS 0.015547f
C314 VTAIL.n245 VSUBS 0.034706f
C315 VTAIL.n246 VSUBS 0.084418f
C316 VTAIL.n247 VSUBS 0.015547f
C317 VTAIL.n248 VSUBS 0.014683f
C318 VTAIL.n249 VSUBS 0.062413f
C319 VTAIL.n250 VSUBS 0.042448f
C320 VTAIL.n251 VSUBS 1.40055f
C321 VTAIL.n252 VSUBS 0.030141f
C322 VTAIL.n253 VSUBS 0.027325f
C323 VTAIL.n254 VSUBS 0.014683f
C324 VTAIL.n255 VSUBS 0.034706f
C325 VTAIL.n256 VSUBS 0.015547f
C326 VTAIL.n257 VSUBS 0.027325f
C327 VTAIL.n258 VSUBS 0.014683f
C328 VTAIL.n259 VSUBS 0.034706f
C329 VTAIL.n260 VSUBS 0.015547f
C330 VTAIL.n261 VSUBS 0.714202f
C331 VTAIL.n262 VSUBS 0.014683f
C332 VTAIL.t4 VSUBS 0.074218f
C333 VTAIL.n263 VSUBS 0.126188f
C334 VTAIL.n264 VSUBS 0.022074f
C335 VTAIL.n265 VSUBS 0.026029f
C336 VTAIL.n266 VSUBS 0.034706f
C337 VTAIL.n267 VSUBS 0.015547f
C338 VTAIL.n268 VSUBS 0.014683f
C339 VTAIL.n269 VSUBS 0.027325f
C340 VTAIL.n270 VSUBS 0.027325f
C341 VTAIL.n271 VSUBS 0.014683f
C342 VTAIL.n272 VSUBS 0.015547f
C343 VTAIL.n273 VSUBS 0.034706f
C344 VTAIL.n274 VSUBS 0.034706f
C345 VTAIL.n275 VSUBS 0.015547f
C346 VTAIL.n276 VSUBS 0.014683f
C347 VTAIL.n277 VSUBS 0.027325f
C348 VTAIL.n278 VSUBS 0.027325f
C349 VTAIL.n279 VSUBS 0.014683f
C350 VTAIL.n280 VSUBS 0.015547f
C351 VTAIL.n281 VSUBS 0.034706f
C352 VTAIL.n282 VSUBS 0.084418f
C353 VTAIL.n283 VSUBS 0.015547f
C354 VTAIL.n284 VSUBS 0.014683f
C355 VTAIL.n285 VSUBS 0.062413f
C356 VTAIL.n286 VSUBS 0.042448f
C357 VTAIL.n287 VSUBS 1.27095f
C358 VN.t3 VSUBS 2.34461f
C359 VN.t2 VSUBS 2.35526f
C360 VN.n0 VSUBS 1.44108f
C361 VN.t0 VSUBS 2.35526f
C362 VN.t1 VSUBS 2.34461f
C363 VN.n1 VSUBS 3.39594f
C364 B.n0 VSUBS 0.00495f
C365 B.n1 VSUBS 0.00495f
C366 B.n2 VSUBS 0.007828f
C367 B.n3 VSUBS 0.007828f
C368 B.n4 VSUBS 0.007828f
C369 B.n5 VSUBS 0.007828f
C370 B.n6 VSUBS 0.007828f
C371 B.n7 VSUBS 0.007828f
C372 B.n8 VSUBS 0.007828f
C373 B.n9 VSUBS 0.007828f
C374 B.n10 VSUBS 0.007828f
C375 B.n11 VSUBS 0.007828f
C376 B.n12 VSUBS 0.007828f
C377 B.n13 VSUBS 0.007828f
C378 B.n14 VSUBS 0.007828f
C379 B.n15 VSUBS 0.007828f
C380 B.n16 VSUBS 0.007828f
C381 B.n17 VSUBS 0.007828f
C382 B.n18 VSUBS 0.007828f
C383 B.n19 VSUBS 0.007828f
C384 B.n20 VSUBS 0.017076f
C385 B.n21 VSUBS 0.007828f
C386 B.n22 VSUBS 0.007828f
C387 B.n23 VSUBS 0.007828f
C388 B.n24 VSUBS 0.007828f
C389 B.n25 VSUBS 0.007828f
C390 B.n26 VSUBS 0.007828f
C391 B.n27 VSUBS 0.007828f
C392 B.n28 VSUBS 0.007828f
C393 B.n29 VSUBS 0.007828f
C394 B.n30 VSUBS 0.007828f
C395 B.n31 VSUBS 0.007828f
C396 B.n32 VSUBS 0.007828f
C397 B.n33 VSUBS 0.007828f
C398 B.t11 VSUBS 0.114119f
C399 B.t10 VSUBS 0.147326f
C400 B.t9 VSUBS 1.04655f
C401 B.n34 VSUBS 0.246366f
C402 B.n35 VSUBS 0.190834f
C403 B.n36 VSUBS 0.007828f
C404 B.n37 VSUBS 0.007828f
C405 B.n38 VSUBS 0.007828f
C406 B.n39 VSUBS 0.007828f
C407 B.n40 VSUBS 0.004375f
C408 B.n41 VSUBS 0.007828f
C409 B.t2 VSUBS 0.114122f
C410 B.t1 VSUBS 0.147327f
C411 B.t0 VSUBS 1.04655f
C412 B.n42 VSUBS 0.246365f
C413 B.n43 VSUBS 0.190832f
C414 B.n44 VSUBS 0.018137f
C415 B.n45 VSUBS 0.007828f
C416 B.n46 VSUBS 0.007828f
C417 B.n47 VSUBS 0.007828f
C418 B.n48 VSUBS 0.007828f
C419 B.n49 VSUBS 0.007828f
C420 B.n50 VSUBS 0.007828f
C421 B.n51 VSUBS 0.007828f
C422 B.n52 VSUBS 0.007828f
C423 B.n53 VSUBS 0.007828f
C424 B.n54 VSUBS 0.007828f
C425 B.n55 VSUBS 0.007828f
C426 B.n56 VSUBS 0.018381f
C427 B.n57 VSUBS 0.007828f
C428 B.n58 VSUBS 0.007828f
C429 B.n59 VSUBS 0.007828f
C430 B.n60 VSUBS 0.007828f
C431 B.n61 VSUBS 0.007828f
C432 B.n62 VSUBS 0.007828f
C433 B.n63 VSUBS 0.007828f
C434 B.n64 VSUBS 0.007828f
C435 B.n65 VSUBS 0.007828f
C436 B.n66 VSUBS 0.007828f
C437 B.n67 VSUBS 0.007828f
C438 B.n68 VSUBS 0.007828f
C439 B.n69 VSUBS 0.007828f
C440 B.n70 VSUBS 0.007828f
C441 B.n71 VSUBS 0.007828f
C442 B.n72 VSUBS 0.007828f
C443 B.n73 VSUBS 0.007828f
C444 B.n74 VSUBS 0.007828f
C445 B.n75 VSUBS 0.007828f
C446 B.n76 VSUBS 0.007828f
C447 B.n77 VSUBS 0.007828f
C448 B.n78 VSUBS 0.007828f
C449 B.n79 VSUBS 0.007828f
C450 B.n80 VSUBS 0.007828f
C451 B.n81 VSUBS 0.007828f
C452 B.n82 VSUBS 0.007828f
C453 B.n83 VSUBS 0.007828f
C454 B.n84 VSUBS 0.007828f
C455 B.n85 VSUBS 0.007828f
C456 B.n86 VSUBS 0.007828f
C457 B.n87 VSUBS 0.007828f
C458 B.n88 VSUBS 0.007828f
C459 B.n89 VSUBS 0.007828f
C460 B.n90 VSUBS 0.007828f
C461 B.n91 VSUBS 0.007828f
C462 B.n92 VSUBS 0.007828f
C463 B.n93 VSUBS 0.007828f
C464 B.n94 VSUBS 0.018381f
C465 B.n95 VSUBS 0.007828f
C466 B.n96 VSUBS 0.007828f
C467 B.n97 VSUBS 0.007828f
C468 B.n98 VSUBS 0.007828f
C469 B.n99 VSUBS 0.007828f
C470 B.n100 VSUBS 0.007828f
C471 B.n101 VSUBS 0.007828f
C472 B.n102 VSUBS 0.007828f
C473 B.n103 VSUBS 0.007828f
C474 B.n104 VSUBS 0.007828f
C475 B.n105 VSUBS 0.007828f
C476 B.n106 VSUBS 0.007828f
C477 B.t4 VSUBS 0.114122f
C478 B.t5 VSUBS 0.147327f
C479 B.t3 VSUBS 1.04655f
C480 B.n107 VSUBS 0.246365f
C481 B.n108 VSUBS 0.190832f
C482 B.n109 VSUBS 0.018137f
C483 B.n110 VSUBS 0.007828f
C484 B.n111 VSUBS 0.007828f
C485 B.n112 VSUBS 0.007828f
C486 B.n113 VSUBS 0.007828f
C487 B.n114 VSUBS 0.007828f
C488 B.t7 VSUBS 0.114119f
C489 B.t8 VSUBS 0.147326f
C490 B.t6 VSUBS 1.04655f
C491 B.n115 VSUBS 0.246366f
C492 B.n116 VSUBS 0.190834f
C493 B.n117 VSUBS 0.007828f
C494 B.n118 VSUBS 0.007828f
C495 B.n119 VSUBS 0.007828f
C496 B.n120 VSUBS 0.007828f
C497 B.n121 VSUBS 0.007828f
C498 B.n122 VSUBS 0.007828f
C499 B.n123 VSUBS 0.007828f
C500 B.n124 VSUBS 0.007828f
C501 B.n125 VSUBS 0.007828f
C502 B.n126 VSUBS 0.007828f
C503 B.n127 VSUBS 0.007828f
C504 B.n128 VSUBS 0.007828f
C505 B.n129 VSUBS 0.018381f
C506 B.n130 VSUBS 0.007828f
C507 B.n131 VSUBS 0.007828f
C508 B.n132 VSUBS 0.007828f
C509 B.n133 VSUBS 0.007828f
C510 B.n134 VSUBS 0.007828f
C511 B.n135 VSUBS 0.007828f
C512 B.n136 VSUBS 0.007828f
C513 B.n137 VSUBS 0.007828f
C514 B.n138 VSUBS 0.007828f
C515 B.n139 VSUBS 0.007828f
C516 B.n140 VSUBS 0.007828f
C517 B.n141 VSUBS 0.007828f
C518 B.n142 VSUBS 0.007828f
C519 B.n143 VSUBS 0.007828f
C520 B.n144 VSUBS 0.007828f
C521 B.n145 VSUBS 0.007828f
C522 B.n146 VSUBS 0.007828f
C523 B.n147 VSUBS 0.007828f
C524 B.n148 VSUBS 0.007828f
C525 B.n149 VSUBS 0.007828f
C526 B.n150 VSUBS 0.007828f
C527 B.n151 VSUBS 0.007828f
C528 B.n152 VSUBS 0.007828f
C529 B.n153 VSUBS 0.007828f
C530 B.n154 VSUBS 0.007828f
C531 B.n155 VSUBS 0.007828f
C532 B.n156 VSUBS 0.007828f
C533 B.n157 VSUBS 0.007828f
C534 B.n158 VSUBS 0.007828f
C535 B.n159 VSUBS 0.007828f
C536 B.n160 VSUBS 0.007828f
C537 B.n161 VSUBS 0.007828f
C538 B.n162 VSUBS 0.007828f
C539 B.n163 VSUBS 0.007828f
C540 B.n164 VSUBS 0.007828f
C541 B.n165 VSUBS 0.007828f
C542 B.n166 VSUBS 0.007828f
C543 B.n167 VSUBS 0.007828f
C544 B.n168 VSUBS 0.007828f
C545 B.n169 VSUBS 0.007828f
C546 B.n170 VSUBS 0.007828f
C547 B.n171 VSUBS 0.007828f
C548 B.n172 VSUBS 0.007828f
C549 B.n173 VSUBS 0.007828f
C550 B.n174 VSUBS 0.007828f
C551 B.n175 VSUBS 0.007828f
C552 B.n176 VSUBS 0.007828f
C553 B.n177 VSUBS 0.007828f
C554 B.n178 VSUBS 0.007828f
C555 B.n179 VSUBS 0.007828f
C556 B.n180 VSUBS 0.007828f
C557 B.n181 VSUBS 0.007828f
C558 B.n182 VSUBS 0.007828f
C559 B.n183 VSUBS 0.007828f
C560 B.n184 VSUBS 0.007828f
C561 B.n185 VSUBS 0.007828f
C562 B.n186 VSUBS 0.007828f
C563 B.n187 VSUBS 0.007828f
C564 B.n188 VSUBS 0.007828f
C565 B.n189 VSUBS 0.007828f
C566 B.n190 VSUBS 0.007828f
C567 B.n191 VSUBS 0.007828f
C568 B.n192 VSUBS 0.007828f
C569 B.n193 VSUBS 0.007828f
C570 B.n194 VSUBS 0.007828f
C571 B.n195 VSUBS 0.007828f
C572 B.n196 VSUBS 0.007828f
C573 B.n197 VSUBS 0.007828f
C574 B.n198 VSUBS 0.007828f
C575 B.n199 VSUBS 0.007828f
C576 B.n200 VSUBS 0.017076f
C577 B.n201 VSUBS 0.017076f
C578 B.n202 VSUBS 0.018381f
C579 B.n203 VSUBS 0.007828f
C580 B.n204 VSUBS 0.007828f
C581 B.n205 VSUBS 0.007828f
C582 B.n206 VSUBS 0.007828f
C583 B.n207 VSUBS 0.007828f
C584 B.n208 VSUBS 0.007828f
C585 B.n209 VSUBS 0.007828f
C586 B.n210 VSUBS 0.007828f
C587 B.n211 VSUBS 0.007828f
C588 B.n212 VSUBS 0.007828f
C589 B.n213 VSUBS 0.007828f
C590 B.n214 VSUBS 0.007828f
C591 B.n215 VSUBS 0.007828f
C592 B.n216 VSUBS 0.007828f
C593 B.n217 VSUBS 0.007828f
C594 B.n218 VSUBS 0.007828f
C595 B.n219 VSUBS 0.007828f
C596 B.n220 VSUBS 0.007828f
C597 B.n221 VSUBS 0.007828f
C598 B.n222 VSUBS 0.007828f
C599 B.n223 VSUBS 0.007828f
C600 B.n224 VSUBS 0.007828f
C601 B.n225 VSUBS 0.007828f
C602 B.n226 VSUBS 0.007828f
C603 B.n227 VSUBS 0.007828f
C604 B.n228 VSUBS 0.007828f
C605 B.n229 VSUBS 0.007828f
C606 B.n230 VSUBS 0.007828f
C607 B.n231 VSUBS 0.007828f
C608 B.n232 VSUBS 0.007828f
C609 B.n233 VSUBS 0.007828f
C610 B.n234 VSUBS 0.007828f
C611 B.n235 VSUBS 0.007828f
C612 B.n236 VSUBS 0.007828f
C613 B.n237 VSUBS 0.007828f
C614 B.n238 VSUBS 0.007828f
C615 B.n239 VSUBS 0.007828f
C616 B.n240 VSUBS 0.007368f
C617 B.n241 VSUBS 0.018137f
C618 B.n242 VSUBS 0.004375f
C619 B.n243 VSUBS 0.007828f
C620 B.n244 VSUBS 0.007828f
C621 B.n245 VSUBS 0.007828f
C622 B.n246 VSUBS 0.007828f
C623 B.n247 VSUBS 0.007828f
C624 B.n248 VSUBS 0.007828f
C625 B.n249 VSUBS 0.007828f
C626 B.n250 VSUBS 0.007828f
C627 B.n251 VSUBS 0.007828f
C628 B.n252 VSUBS 0.007828f
C629 B.n253 VSUBS 0.007828f
C630 B.n254 VSUBS 0.007828f
C631 B.n255 VSUBS 0.004375f
C632 B.n256 VSUBS 0.007828f
C633 B.n257 VSUBS 0.007828f
C634 B.n258 VSUBS 0.007368f
C635 B.n259 VSUBS 0.007828f
C636 B.n260 VSUBS 0.007828f
C637 B.n261 VSUBS 0.007828f
C638 B.n262 VSUBS 0.007828f
C639 B.n263 VSUBS 0.007828f
C640 B.n264 VSUBS 0.007828f
C641 B.n265 VSUBS 0.007828f
C642 B.n266 VSUBS 0.007828f
C643 B.n267 VSUBS 0.007828f
C644 B.n268 VSUBS 0.007828f
C645 B.n269 VSUBS 0.007828f
C646 B.n270 VSUBS 0.007828f
C647 B.n271 VSUBS 0.007828f
C648 B.n272 VSUBS 0.007828f
C649 B.n273 VSUBS 0.007828f
C650 B.n274 VSUBS 0.007828f
C651 B.n275 VSUBS 0.007828f
C652 B.n276 VSUBS 0.007828f
C653 B.n277 VSUBS 0.007828f
C654 B.n278 VSUBS 0.007828f
C655 B.n279 VSUBS 0.007828f
C656 B.n280 VSUBS 0.007828f
C657 B.n281 VSUBS 0.007828f
C658 B.n282 VSUBS 0.007828f
C659 B.n283 VSUBS 0.007828f
C660 B.n284 VSUBS 0.007828f
C661 B.n285 VSUBS 0.007828f
C662 B.n286 VSUBS 0.007828f
C663 B.n287 VSUBS 0.007828f
C664 B.n288 VSUBS 0.007828f
C665 B.n289 VSUBS 0.007828f
C666 B.n290 VSUBS 0.007828f
C667 B.n291 VSUBS 0.007828f
C668 B.n292 VSUBS 0.007828f
C669 B.n293 VSUBS 0.007828f
C670 B.n294 VSUBS 0.007828f
C671 B.n295 VSUBS 0.018381f
C672 B.n296 VSUBS 0.017076f
C673 B.n297 VSUBS 0.017076f
C674 B.n298 VSUBS 0.007828f
C675 B.n299 VSUBS 0.007828f
C676 B.n300 VSUBS 0.007828f
C677 B.n301 VSUBS 0.007828f
C678 B.n302 VSUBS 0.007828f
C679 B.n303 VSUBS 0.007828f
C680 B.n304 VSUBS 0.007828f
C681 B.n305 VSUBS 0.007828f
C682 B.n306 VSUBS 0.007828f
C683 B.n307 VSUBS 0.007828f
C684 B.n308 VSUBS 0.007828f
C685 B.n309 VSUBS 0.007828f
C686 B.n310 VSUBS 0.007828f
C687 B.n311 VSUBS 0.007828f
C688 B.n312 VSUBS 0.007828f
C689 B.n313 VSUBS 0.007828f
C690 B.n314 VSUBS 0.007828f
C691 B.n315 VSUBS 0.007828f
C692 B.n316 VSUBS 0.007828f
C693 B.n317 VSUBS 0.007828f
C694 B.n318 VSUBS 0.007828f
C695 B.n319 VSUBS 0.007828f
C696 B.n320 VSUBS 0.007828f
C697 B.n321 VSUBS 0.007828f
C698 B.n322 VSUBS 0.007828f
C699 B.n323 VSUBS 0.007828f
C700 B.n324 VSUBS 0.007828f
C701 B.n325 VSUBS 0.007828f
C702 B.n326 VSUBS 0.007828f
C703 B.n327 VSUBS 0.007828f
C704 B.n328 VSUBS 0.007828f
C705 B.n329 VSUBS 0.007828f
C706 B.n330 VSUBS 0.007828f
C707 B.n331 VSUBS 0.007828f
C708 B.n332 VSUBS 0.007828f
C709 B.n333 VSUBS 0.007828f
C710 B.n334 VSUBS 0.007828f
C711 B.n335 VSUBS 0.007828f
C712 B.n336 VSUBS 0.007828f
C713 B.n337 VSUBS 0.007828f
C714 B.n338 VSUBS 0.007828f
C715 B.n339 VSUBS 0.007828f
C716 B.n340 VSUBS 0.007828f
C717 B.n341 VSUBS 0.007828f
C718 B.n342 VSUBS 0.007828f
C719 B.n343 VSUBS 0.007828f
C720 B.n344 VSUBS 0.007828f
C721 B.n345 VSUBS 0.007828f
C722 B.n346 VSUBS 0.007828f
C723 B.n347 VSUBS 0.007828f
C724 B.n348 VSUBS 0.007828f
C725 B.n349 VSUBS 0.007828f
C726 B.n350 VSUBS 0.007828f
C727 B.n351 VSUBS 0.007828f
C728 B.n352 VSUBS 0.007828f
C729 B.n353 VSUBS 0.007828f
C730 B.n354 VSUBS 0.007828f
C731 B.n355 VSUBS 0.007828f
C732 B.n356 VSUBS 0.007828f
C733 B.n357 VSUBS 0.007828f
C734 B.n358 VSUBS 0.007828f
C735 B.n359 VSUBS 0.007828f
C736 B.n360 VSUBS 0.007828f
C737 B.n361 VSUBS 0.007828f
C738 B.n362 VSUBS 0.007828f
C739 B.n363 VSUBS 0.007828f
C740 B.n364 VSUBS 0.007828f
C741 B.n365 VSUBS 0.007828f
C742 B.n366 VSUBS 0.007828f
C743 B.n367 VSUBS 0.007828f
C744 B.n368 VSUBS 0.007828f
C745 B.n369 VSUBS 0.007828f
C746 B.n370 VSUBS 0.007828f
C747 B.n371 VSUBS 0.007828f
C748 B.n372 VSUBS 0.007828f
C749 B.n373 VSUBS 0.007828f
C750 B.n374 VSUBS 0.007828f
C751 B.n375 VSUBS 0.007828f
C752 B.n376 VSUBS 0.007828f
C753 B.n377 VSUBS 0.007828f
C754 B.n378 VSUBS 0.007828f
C755 B.n379 VSUBS 0.007828f
C756 B.n380 VSUBS 0.007828f
C757 B.n381 VSUBS 0.007828f
C758 B.n382 VSUBS 0.007828f
C759 B.n383 VSUBS 0.007828f
C760 B.n384 VSUBS 0.007828f
C761 B.n385 VSUBS 0.007828f
C762 B.n386 VSUBS 0.007828f
C763 B.n387 VSUBS 0.007828f
C764 B.n388 VSUBS 0.007828f
C765 B.n389 VSUBS 0.007828f
C766 B.n390 VSUBS 0.007828f
C767 B.n391 VSUBS 0.007828f
C768 B.n392 VSUBS 0.007828f
C769 B.n393 VSUBS 0.007828f
C770 B.n394 VSUBS 0.007828f
C771 B.n395 VSUBS 0.007828f
C772 B.n396 VSUBS 0.007828f
C773 B.n397 VSUBS 0.007828f
C774 B.n398 VSUBS 0.007828f
C775 B.n399 VSUBS 0.007828f
C776 B.n400 VSUBS 0.007828f
C777 B.n401 VSUBS 0.007828f
C778 B.n402 VSUBS 0.007828f
C779 B.n403 VSUBS 0.007828f
C780 B.n404 VSUBS 0.007828f
C781 B.n405 VSUBS 0.007828f
C782 B.n406 VSUBS 0.007828f
C783 B.n407 VSUBS 0.017076f
C784 B.n408 VSUBS 0.018049f
C785 B.n409 VSUBS 0.017409f
C786 B.n410 VSUBS 0.007828f
C787 B.n411 VSUBS 0.007828f
C788 B.n412 VSUBS 0.007828f
C789 B.n413 VSUBS 0.007828f
C790 B.n414 VSUBS 0.007828f
C791 B.n415 VSUBS 0.007828f
C792 B.n416 VSUBS 0.007828f
C793 B.n417 VSUBS 0.007828f
C794 B.n418 VSUBS 0.007828f
C795 B.n419 VSUBS 0.007828f
C796 B.n420 VSUBS 0.007828f
C797 B.n421 VSUBS 0.007828f
C798 B.n422 VSUBS 0.007828f
C799 B.n423 VSUBS 0.007828f
C800 B.n424 VSUBS 0.007828f
C801 B.n425 VSUBS 0.007828f
C802 B.n426 VSUBS 0.007828f
C803 B.n427 VSUBS 0.007828f
C804 B.n428 VSUBS 0.007828f
C805 B.n429 VSUBS 0.007828f
C806 B.n430 VSUBS 0.007828f
C807 B.n431 VSUBS 0.007828f
C808 B.n432 VSUBS 0.007828f
C809 B.n433 VSUBS 0.007828f
C810 B.n434 VSUBS 0.007828f
C811 B.n435 VSUBS 0.007828f
C812 B.n436 VSUBS 0.007828f
C813 B.n437 VSUBS 0.007828f
C814 B.n438 VSUBS 0.007828f
C815 B.n439 VSUBS 0.007828f
C816 B.n440 VSUBS 0.007828f
C817 B.n441 VSUBS 0.007828f
C818 B.n442 VSUBS 0.007828f
C819 B.n443 VSUBS 0.007828f
C820 B.n444 VSUBS 0.007828f
C821 B.n445 VSUBS 0.007828f
C822 B.n446 VSUBS 0.007368f
C823 B.n447 VSUBS 0.007828f
C824 B.n448 VSUBS 0.007828f
C825 B.n449 VSUBS 0.007828f
C826 B.n450 VSUBS 0.007828f
C827 B.n451 VSUBS 0.007828f
C828 B.n452 VSUBS 0.007828f
C829 B.n453 VSUBS 0.007828f
C830 B.n454 VSUBS 0.007828f
C831 B.n455 VSUBS 0.007828f
C832 B.n456 VSUBS 0.007828f
C833 B.n457 VSUBS 0.007828f
C834 B.n458 VSUBS 0.007828f
C835 B.n459 VSUBS 0.007828f
C836 B.n460 VSUBS 0.007828f
C837 B.n461 VSUBS 0.007828f
C838 B.n462 VSUBS 0.004375f
C839 B.n463 VSUBS 0.018137f
C840 B.n464 VSUBS 0.007368f
C841 B.n465 VSUBS 0.007828f
C842 B.n466 VSUBS 0.007828f
C843 B.n467 VSUBS 0.007828f
C844 B.n468 VSUBS 0.007828f
C845 B.n469 VSUBS 0.007828f
C846 B.n470 VSUBS 0.007828f
C847 B.n471 VSUBS 0.007828f
C848 B.n472 VSUBS 0.007828f
C849 B.n473 VSUBS 0.007828f
C850 B.n474 VSUBS 0.007828f
C851 B.n475 VSUBS 0.007828f
C852 B.n476 VSUBS 0.007828f
C853 B.n477 VSUBS 0.007828f
C854 B.n478 VSUBS 0.007828f
C855 B.n479 VSUBS 0.007828f
C856 B.n480 VSUBS 0.007828f
C857 B.n481 VSUBS 0.007828f
C858 B.n482 VSUBS 0.007828f
C859 B.n483 VSUBS 0.007828f
C860 B.n484 VSUBS 0.007828f
C861 B.n485 VSUBS 0.007828f
C862 B.n486 VSUBS 0.007828f
C863 B.n487 VSUBS 0.007828f
C864 B.n488 VSUBS 0.007828f
C865 B.n489 VSUBS 0.007828f
C866 B.n490 VSUBS 0.007828f
C867 B.n491 VSUBS 0.007828f
C868 B.n492 VSUBS 0.007828f
C869 B.n493 VSUBS 0.007828f
C870 B.n494 VSUBS 0.007828f
C871 B.n495 VSUBS 0.007828f
C872 B.n496 VSUBS 0.007828f
C873 B.n497 VSUBS 0.007828f
C874 B.n498 VSUBS 0.007828f
C875 B.n499 VSUBS 0.007828f
C876 B.n500 VSUBS 0.007828f
C877 B.n501 VSUBS 0.018381f
C878 B.n502 VSUBS 0.018381f
C879 B.n503 VSUBS 0.017076f
C880 B.n504 VSUBS 0.007828f
C881 B.n505 VSUBS 0.007828f
C882 B.n506 VSUBS 0.007828f
C883 B.n507 VSUBS 0.007828f
C884 B.n508 VSUBS 0.007828f
C885 B.n509 VSUBS 0.007828f
C886 B.n510 VSUBS 0.007828f
C887 B.n511 VSUBS 0.007828f
C888 B.n512 VSUBS 0.007828f
C889 B.n513 VSUBS 0.007828f
C890 B.n514 VSUBS 0.007828f
C891 B.n515 VSUBS 0.007828f
C892 B.n516 VSUBS 0.007828f
C893 B.n517 VSUBS 0.007828f
C894 B.n518 VSUBS 0.007828f
C895 B.n519 VSUBS 0.007828f
C896 B.n520 VSUBS 0.007828f
C897 B.n521 VSUBS 0.007828f
C898 B.n522 VSUBS 0.007828f
C899 B.n523 VSUBS 0.007828f
C900 B.n524 VSUBS 0.007828f
C901 B.n525 VSUBS 0.007828f
C902 B.n526 VSUBS 0.007828f
C903 B.n527 VSUBS 0.007828f
C904 B.n528 VSUBS 0.007828f
C905 B.n529 VSUBS 0.007828f
C906 B.n530 VSUBS 0.007828f
C907 B.n531 VSUBS 0.007828f
C908 B.n532 VSUBS 0.007828f
C909 B.n533 VSUBS 0.007828f
C910 B.n534 VSUBS 0.007828f
C911 B.n535 VSUBS 0.007828f
C912 B.n536 VSUBS 0.007828f
C913 B.n537 VSUBS 0.007828f
C914 B.n538 VSUBS 0.007828f
C915 B.n539 VSUBS 0.007828f
C916 B.n540 VSUBS 0.007828f
C917 B.n541 VSUBS 0.007828f
C918 B.n542 VSUBS 0.007828f
C919 B.n543 VSUBS 0.007828f
C920 B.n544 VSUBS 0.007828f
C921 B.n545 VSUBS 0.007828f
C922 B.n546 VSUBS 0.007828f
C923 B.n547 VSUBS 0.007828f
C924 B.n548 VSUBS 0.007828f
C925 B.n549 VSUBS 0.007828f
C926 B.n550 VSUBS 0.007828f
C927 B.n551 VSUBS 0.007828f
C928 B.n552 VSUBS 0.007828f
C929 B.n553 VSUBS 0.007828f
C930 B.n554 VSUBS 0.007828f
C931 B.n555 VSUBS 0.007828f
C932 B.n556 VSUBS 0.007828f
C933 B.n557 VSUBS 0.007828f
C934 B.n558 VSUBS 0.007828f
C935 B.n559 VSUBS 0.017726f
.ends

