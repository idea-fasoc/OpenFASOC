* NGSPICE file created from opamp_sample_0007.ext - technology: sky130A

.subckt opamp_sample_0007 GND VOUT VDD VN VP CS_BIAS DIFFPAIR_BIAS
X0 a_n8335_8538.t6 a_n8335_8538.t5 a_n8413_8735.t15 VDD.t100 sky130_fd_pr__pfet_01v8 ad=0.46035 pd=3.12 as=0.46035 ps=3.12 w=2.79 l=4.28
X1 GND.t156 GND.t154 GND.t155 GND.t73 sky130_fd_pr__nfet_01v8 ad=1.3104 pd=7.5 as=0 ps=0 w=3.36 l=6.01
X2 GND.t153 GND.t151 VP.t1 GND.t152 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X3 VDD.t117 a_n8335_8538.t18 a_n5434_7417.t11 VDD.t116 sky130_fd_pr__pfet_01v8 ad=0.46035 pd=3.12 as=0.46035 ps=3.12 w=2.79 l=4.28
X4 GND.t150 GND.t148 GND.t149 GND.t63 sky130_fd_pr__nfet_01v8 ad=0.936 pd=5.58 as=0 ps=0 w=2.4 l=3.51
X5 a_n8335_8538.t16 a_n8335_8538.t15 a_n8413_8735.t14 VDD.t96 sky130_fd_pr__pfet_01v8 ad=1.0881 pd=6.36 as=0.46035 ps=3.12 w=2.79 l=4.28
X6 VDD.t115 a_n8335_8538.t19 a_n8413_8735.t4 VDD.t114 sky130_fd_pr__pfet_01v8 ad=0.46035 pd=3.12 as=1.0881 ps=6.36 w=2.79 l=4.28
X7 VDD.t70 VDD.t68 VDD.t69 VDD.t45 sky130_fd_pr__pfet_01v8 ad=1.9812 pd=10.94 as=0 ps=0 w=5.08 l=3.15
X8 VDD.t67 VDD.t65 VDD.t66 VDD.t45 sky130_fd_pr__pfet_01v8 ad=1.9812 pd=10.94 as=0 ps=0 w=5.08 l=3.15
X9 GND.t32 CS_BIAS.t16 VOUT.t39 GND.t12 sky130_fd_pr__nfet_01v8 ad=0.936 pd=5.58 as=0.396 ps=2.73 w=2.4 l=3.51
X10 VOUT.t46 a_n5434_7417.t0 sky130_fd_pr__cap_mim_m3_1 l=9.91 w=17.88
X11 VOUT.t38 CS_BIAS.t17 GND.t34 GND.t19 sky130_fd_pr__nfet_01v8 ad=0.396 pd=2.73 as=0.396 ps=2.73 w=2.4 l=3.51
X12 a_n8413_8735.t13 a_n8335_8538.t13 a_n8335_8538.t14 VDD.t101 sky130_fd_pr__pfet_01v8 ad=0.46035 pd=3.12 as=0.46035 ps=3.12 w=2.79 l=4.28
X13 a_n8413_8735.t12 a_n8335_8538.t11 a_n8335_8538.t12 VDD.t87 sky130_fd_pr__pfet_01v8 ad=0.46035 pd=3.12 as=1.0881 ps=6.36 w=2.79 l=4.28
X14 VOUT.t47 a_n5434_7417.t0 sky130_fd_pr__cap_mim_m3_1 l=9.91 w=17.88
X15 GND.t147 GND.t145 GND.t146 GND.t52 sky130_fd_pr__nfet_01v8 ad=0.936 pd=5.58 as=0 ps=0 w=2.4 l=3.51
X16 a_n8335_8538.t4 a_n8335_8538.t3 a_n8413_8735.t11 VDD.t90 sky130_fd_pr__pfet_01v8 ad=0.46035 pd=3.12 as=0.46035 ps=3.12 w=2.79 l=4.28
X17 a_n8335_8538.t8 a_n8335_8538.t7 a_n8413_8735.t10 VDD.t97 sky130_fd_pr__pfet_01v8 ad=1.0881 pd=6.36 as=0.46035 ps=3.12 w=2.79 l=4.28
X18 GND.t14 CS_BIAS.t18 VOUT.t37 GND.t5 sky130_fd_pr__nfet_01v8 ad=0.936 pd=5.58 as=0.396 ps=2.73 w=2.4 l=3.51
X19 a_n8413_8735.t9 a_n8335_8538.t1 a_n8335_8538.t2 VDD.t93 sky130_fd_pr__pfet_01v8 ad=0.46035 pd=3.12 as=0.46035 ps=3.12 w=2.79 l=4.28
X20 VDD.t64 VDD.t62 VDD.t63 VDD.t59 sky130_fd_pr__pfet_01v8 ad=1.0881 pd=6.36 as=0 ps=0 w=2.79 l=4.28
X21 GND.t42 CS_BIAS.t19 VOUT.t36 GND.t0 sky130_fd_pr__nfet_01v8 ad=0.396 pd=2.73 as=0.396 ps=2.73 w=2.4 l=3.51
X22 VDD.t61 VDD.t58 VDD.t60 VDD.t59 sky130_fd_pr__pfet_01v8 ad=1.0881 pd=6.36 as=0 ps=0 w=2.79 l=4.28
X23 VDD.t57 VDD.t55 VDD.t56 VDD.t49 sky130_fd_pr__pfet_01v8 ad=1.0881 pd=6.36 as=0 ps=0 w=2.79 l=4.28
X24 VOUT.t35 CS_BIAS.t20 GND.t40 GND.t21 sky130_fd_pr__nfet_01v8 ad=0.396 pd=2.73 as=0.936 ps=5.58 w=2.4 l=3.51
X25 CS_BIAS.t15 CS_BIAS.t14 GND.t38 GND.t2 sky130_fd_pr__nfet_01v8 ad=0.396 pd=2.73 as=0.936 ps=5.58 w=2.4 l=3.51
X26 GND.t144 GND.t142 GND.t143 GND.t63 sky130_fd_pr__nfet_01v8 ad=0.936 pd=5.58 as=0 ps=0 w=2.4 l=3.51
X27 GND.t46 CS_BIAS.t21 VOUT.t34 GND.t12 sky130_fd_pr__nfet_01v8 ad=0.936 pd=5.58 as=0.396 ps=2.73 w=2.4 l=3.51
X28 VOUT.t33 CS_BIAS.t22 GND.t165 GND.t9 sky130_fd_pr__nfet_01v8 ad=0.396 pd=2.73 as=0.396 ps=2.73 w=2.4 l=3.51
X29 GND.t7 CS_BIAS.t23 VOUT.t32 GND.t5 sky130_fd_pr__nfet_01v8 ad=0.936 pd=5.58 as=0.396 ps=2.73 w=2.4 l=3.51
X30 GND.t141 GND.t139 GND.t140 GND.t48 sky130_fd_pr__nfet_01v8 ad=1.3104 pd=7.5 as=0 ps=0 w=3.36 l=6.01
X31 GND.t138 GND.t136 GND.t137 GND.t59 sky130_fd_pr__nfet_01v8 ad=0.936 pd=5.58 as=0 ps=0 w=2.4 l=3.51
X32 VDD.t54 VDD.t52 VDD.t53 VDD.t4 sky130_fd_pr__pfet_01v8 ad=1.0881 pd=6.36 as=0 ps=0 w=2.79 l=4.28
X33 GND.t135 GND.t133 GND.t134 GND.t77 sky130_fd_pr__nfet_01v8 ad=0.936 pd=5.58 as=0 ps=0 w=2.4 l=3.51
X34 VDD.t105 a_n8335_8538.t20 a_n8413_8735.t0 VDD.t104 sky130_fd_pr__pfet_01v8 ad=0.46035 pd=3.12 as=0.46035 ps=3.12 w=2.79 l=4.28
X35 GND.t41 CS_BIAS.t24 VOUT.t31 GND.t15 sky130_fd_pr__nfet_01v8 ad=0.396 pd=2.73 as=0.396 ps=2.73 w=2.4 l=3.51
X36 a_n8335_8538.t17 VP.t2 a_n1578_n2628.t6 GND.t164 sky130_fd_pr__nfet_01v8 ad=1.3104 pd=7.5 as=1.3104 ps=7.5 w=3.36 l=6.01
X37 GND.t132 GND.t130 GND.t131 GND.t63 sky130_fd_pr__nfet_01v8 ad=0.936 pd=5.58 as=0 ps=0 w=2.4 l=3.51
X38 GND.t17 CS_BIAS.t12 CS_BIAS.t13 GND.t12 sky130_fd_pr__nfet_01v8 ad=0.936 pd=5.58 as=0.396 ps=2.73 w=2.4 l=3.51
X39 GND.t39 CS_BIAS.t25 VOUT.t30 GND.t0 sky130_fd_pr__nfet_01v8 ad=0.396 pd=2.73 as=0.396 ps=2.73 w=2.4 l=3.51
X40 VDD.t51 VDD.t48 VDD.t50 VDD.t49 sky130_fd_pr__pfet_01v8 ad=1.0881 pd=6.36 as=0 ps=0 w=2.79 l=4.28
X41 GND.t129 GND.t127 GND.t128 GND.t77 sky130_fd_pr__nfet_01v8 ad=0.936 pd=5.58 as=0 ps=0 w=2.4 l=3.51
X42 GND.t29 CS_BIAS.t26 VOUT.t29 GND.t12 sky130_fd_pr__nfet_01v8 ad=0.936 pd=5.58 as=0.396 ps=2.73 w=2.4 l=3.51
X43 VDD.t47 VDD.t44 VDD.t46 VDD.t45 sky130_fd_pr__pfet_01v8 ad=1.9812 pd=10.94 as=0 ps=0 w=5.08 l=3.15
X44 VOUT.t28 CS_BIAS.t27 GND.t169 GND.t9 sky130_fd_pr__nfet_01v8 ad=0.396 pd=2.73 as=0.396 ps=2.73 w=2.4 l=3.51
X45 VOUT.t27 CS_BIAS.t28 GND.t24 GND.t9 sky130_fd_pr__nfet_01v8 ad=0.396 pd=2.73 as=0.396 ps=2.73 w=2.4 l=3.51
X46 GND.t167 CS_BIAS.t29 VOUT.t26 GND.t0 sky130_fd_pr__nfet_01v8 ad=0.396 pd=2.73 as=0.396 ps=2.73 w=2.4 l=3.51
X47 VDD.t113 a_n8335_8538.t21 a_n5434_7417.t10 VDD.t112 sky130_fd_pr__pfet_01v8 ad=0.46035 pd=3.12 as=1.0881 ps=6.36 w=2.79 l=4.28
X48 VOUT.t25 CS_BIAS.t30 GND.t168 GND.t19 sky130_fd_pr__nfet_01v8 ad=0.396 pd=2.73 as=0.396 ps=2.73 w=2.4 l=3.51
X49 a_n8413_8735.t7 a_n8335_8538.t22 VDD.t111 VDD.t110 sky130_fd_pr__pfet_01v8 ad=1.0881 pd=6.36 as=0.46035 ps=3.12 w=2.79 l=4.28
X50 VOUT.t24 CS_BIAS.t31 GND.t11 GND.t2 sky130_fd_pr__nfet_01v8 ad=0.396 pd=2.73 as=0.936 ps=5.58 w=2.4 l=3.51
X51 VDD.t109 a_n8335_8538.t23 a_n5434_7417.t9 VDD.t108 sky130_fd_pr__pfet_01v8 ad=0.46035 pd=3.12 as=1.0881 ps=6.36 w=2.79 l=4.28
X52 a_n5434_7417.t8 a_n8335_8538.t24 VDD.t107 VDD.t106 sky130_fd_pr__pfet_01v8 ad=0.46035 pd=3.12 as=0.46035 ps=3.12 w=2.79 l=4.28
X53 GND.t126 GND.t124 GND.t125 GND.t77 sky130_fd_pr__nfet_01v8 ad=0.936 pd=5.58 as=0 ps=0 w=2.4 l=3.51
X54 GND.t25 CS_BIAS.t32 VOUT.t23 GND.t15 sky130_fd_pr__nfet_01v8 ad=0.396 pd=2.73 as=0.396 ps=2.73 w=2.4 l=3.51
X55 VP.t0 GND.t121 GND.t123 GND.t122 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X56 VOUT.t41 a_n12120_6849.t10 VDD.t2 VDD.t0 sky130_fd_pr__pfet_01v8 ad=1.9812 pd=10.94 as=1.9812 ps=10.94 w=5.08 l=3.15
X57 VOUT.t43 a_n12120_6849.t11 VDD.t74 VDD.t0 sky130_fd_pr__pfet_01v8 ad=1.9812 pd=10.94 as=1.9812 ps=10.94 w=5.08 l=3.15
X58 VOUT.t48 a_n5434_7417.t0 sky130_fd_pr__cap_mim_m3_1 l=9.91 w=17.88
X59 GND.t120 GND.t118 GND.t119 GND.t52 sky130_fd_pr__nfet_01v8 ad=0.936 pd=5.58 as=0 ps=0 w=2.4 l=3.51
X60 GND.t6 CS_BIAS.t10 CS_BIAS.t11 GND.t5 sky130_fd_pr__nfet_01v8 ad=0.936 pd=5.58 as=0.396 ps=2.73 w=2.4 l=3.51
X61 GND.t117 GND.t115 GND.t116 GND.t59 sky130_fd_pr__nfet_01v8 ad=0.936 pd=5.58 as=0 ps=0 w=2.4 l=3.51
X62 VDD.t103 a_n8335_8538.t25 a_n5434_7417.t7 VDD.t102 sky130_fd_pr__pfet_01v8 ad=0.46035 pd=3.12 as=0.46035 ps=3.12 w=2.79 l=4.28
X63 VDD.t43 VDD.t41 VDD.t42 VDD.t16 sky130_fd_pr__pfet_01v8 ad=1.9812 pd=10.94 as=0 ps=0 w=5.08 l=3.15
X64 VDD.t40 VDD.t38 VDD.t39 VDD.t16 sky130_fd_pr__pfet_01v8 ad=1.9812 pd=10.94 as=0 ps=0 w=5.08 l=3.15
X65 VDD.t37 VDD.t35 VDD.t36 VDD.t20 sky130_fd_pr__pfet_01v8 ad=1.0881 pd=6.36 as=0 ps=0 w=2.79 l=4.28
X66 a_n12120_6849.t9 a_n8335_8538.t26 a_n5434_7417.t12 VDD.t101 sky130_fd_pr__pfet_01v8 ad=0.46035 pd=3.12 as=0.46035 ps=3.12 w=2.79 l=4.28
X67 a_n12120_6849.t1 VN.t2 a_n1578_n2628.t4 GND.t164 sky130_fd_pr__nfet_01v8 ad=1.3104 pd=7.5 as=1.3104 ps=7.5 w=3.36 l=6.01
X68 a_n5434_7417.t1 a_n8335_8538.t27 a_n12120_6849.t8 VDD.t100 sky130_fd_pr__pfet_01v8 ad=0.46035 pd=3.12 as=0.46035 ps=3.12 w=2.79 l=4.28
X69 GND.t166 CS_BIAS.t33 VOUT.t22 GND.t0 sky130_fd_pr__nfet_01v8 ad=0.396 pd=2.73 as=0.396 ps=2.73 w=2.4 l=3.51
X70 GND.t114 GND.t112 GND.t113 GND.t63 sky130_fd_pr__nfet_01v8 ad=0.936 pd=5.58 as=0 ps=0 w=2.4 l=3.51
X71 a_n5434_7417.t6 a_n8335_8538.t28 VDD.t99 VDD.t98 sky130_fd_pr__pfet_01v8 ad=1.0881 pd=6.36 as=0.46035 ps=3.12 w=2.79 l=4.28
X72 a_n12120_6849.t0 VN.t3 a_n1578_n2628.t0 GND.t4 sky130_fd_pr__nfet_01v8 ad=1.3104 pd=7.5 as=1.3104 ps=7.5 w=3.36 l=6.01
X73 GND.t111 GND.t109 GND.t110 GND.t52 sky130_fd_pr__nfet_01v8 ad=0.936 pd=5.58 as=0 ps=0 w=2.4 l=3.51
X74 a_n12120_6849.t7 a_n8335_8538.t29 a_n5434_7417.t15 VDD.t82 sky130_fd_pr__pfet_01v8 ad=0.46035 pd=3.12 as=1.0881 ps=6.36 w=2.79 l=4.28
X75 VDD.t34 VDD.t32 VDD.t33 VDD.t12 sky130_fd_pr__pfet_01v8 ad=1.9812 pd=10.94 as=0 ps=0 w=5.08 l=3.15
X76 VDD.t31 VDD.t29 VDD.t30 VDD.t12 sky130_fd_pr__pfet_01v8 ad=1.9812 pd=10.94 as=0 ps=0 w=5.08 l=3.15
X77 VOUT.t21 CS_BIAS.t34 GND.t3 GND.t2 sky130_fd_pr__nfet_01v8 ad=0.396 pd=2.73 as=0.936 ps=5.58 w=2.4 l=3.51
X78 VOUT.t20 CS_BIAS.t35 GND.t22 GND.t21 sky130_fd_pr__nfet_01v8 ad=0.396 pd=2.73 as=0.936 ps=5.58 w=2.4 l=3.51
X79 VOUT.t45 a_n12120_6849.t12 VDD.t77 VDD.t72 sky130_fd_pr__pfet_01v8 ad=1.9812 pd=10.94 as=1.9812 ps=10.94 w=5.08 l=3.15
X80 VOUT.t44 a_n12120_6849.t13 VDD.t76 VDD.t72 sky130_fd_pr__pfet_01v8 ad=1.9812 pd=10.94 as=1.9812 ps=10.94 w=5.08 l=3.15
X81 GND.t108 GND.t106 GND.t107 GND.t77 sky130_fd_pr__nfet_01v8 ad=0.936 pd=5.58 as=0 ps=0 w=2.4 l=3.51
X82 a_n5434_7417.t13 a_n8335_8538.t30 a_n12120_6849.t6 VDD.t97 sky130_fd_pr__pfet_01v8 ad=1.0881 pd=6.36 as=0.46035 ps=3.12 w=2.79 l=4.28
X83 GND.t105 GND.t103 GND.t104 GND.t77 sky130_fd_pr__nfet_01v8 ad=0.936 pd=5.58 as=0 ps=0 w=2.4 l=3.51
X84 a_n1578_n2628.t3 DIFFPAIR_BIAS.t6 a_n2838_n2628.t2 GND.t159 sky130_fd_pr__nfet_01v8 ad=1.7862 pd=9.94 as=1.7862 ps=9.94 w=4.58 l=5.91
X85 a_n9553_8735# a_n9553_8735# a_n9553_8735# VDD.t75 sky130_fd_pr__pfet_01v8 ad=1.0881 pd=6.36 as=2.1762 ps=12.72 w=2.79 l=4.28
X86 VDD.t28 VDD.t26 VDD.t27 VDD.t8 sky130_fd_pr__pfet_01v8 ad=1.9812 pd=10.94 as=0 ps=0 w=5.08 l=3.15
X87 VDD.t25 VDD.t23 VDD.t24 VDD.t8 sky130_fd_pr__pfet_01v8 ad=1.9812 pd=10.94 as=0 ps=0 w=5.08 l=3.15
X88 VOUT.t19 CS_BIAS.t36 GND.t18 GND.t2 sky130_fd_pr__nfet_01v8 ad=0.396 pd=2.73 as=0.936 ps=5.58 w=2.4 l=3.51
X89 GND.t102 GND.t100 GND.t101 GND.t52 sky130_fd_pr__nfet_01v8 ad=0.936 pd=5.58 as=0 ps=0 w=2.4 l=3.51
X90 GND.t99 GND.t97 GND.t98 GND.t63 sky130_fd_pr__nfet_01v8 ad=0.936 pd=5.58 as=0 ps=0 w=2.4 l=3.51
X91 VDD.t22 VDD.t19 VDD.t21 VDD.t20 sky130_fd_pr__pfet_01v8 ad=1.0881 pd=6.36 as=0 ps=0 w=2.79 l=4.28
X92 GND.t96 GND.t94 GND.t95 GND.t59 sky130_fd_pr__nfet_01v8 ad=0.936 pd=5.58 as=0 ps=0 w=2.4 l=3.51
X93 a_n5434_7417.t2 a_n8335_8538.t31 a_n12120_6849.t5 VDD.t96 sky130_fd_pr__pfet_01v8 ad=1.0881 pd=6.36 as=0.46035 ps=3.12 w=2.79 l=4.28
X94 GND.t163 CS_BIAS.t37 VOUT.t18 GND.t0 sky130_fd_pr__nfet_01v8 ad=0.396 pd=2.73 as=0.396 ps=2.73 w=2.4 l=3.51
X95 VN.t1 GND.t91 GND.t93 GND.t92 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X96 VOUT.t40 a_n12120_6849.t14 VDD.t1 VDD.t0 sky130_fd_pr__pfet_01v8 ad=1.9812 pd=10.94 as=1.9812 ps=10.94 w=5.08 l=3.15
X97 VDD.t95 a_n8335_8538.t32 a_n8413_8735.t5 VDD.t94 sky130_fd_pr__pfet_01v8 ad=0.46035 pd=3.12 as=0.46035 ps=3.12 w=2.79 l=4.28
X98 GND.t1 CS_BIAS.t8 CS_BIAS.t9 GND.t0 sky130_fd_pr__nfet_01v8 ad=0.396 pd=2.73 as=0.396 ps=2.73 w=2.4 l=3.51
X99 GND.t90 GND.t87 GND.t89 GND.t88 sky130_fd_pr__nfet_01v8 ad=1.7862 pd=9.94 as=0 ps=0 w=4.58 l=5.91
X100 VOUT.t17 CS_BIAS.t38 GND.t170 GND.t9 sky130_fd_pr__nfet_01v8 ad=0.396 pd=2.73 as=0.396 ps=2.73 w=2.4 l=3.51
X101 VOUT.t16 CS_BIAS.t39 GND.t173 GND.t21 sky130_fd_pr__nfet_01v8 ad=0.396 pd=2.73 as=0.936 ps=5.58 w=2.4 l=3.51
X102 VDD.t18 VDD.t15 VDD.t17 VDD.t16 sky130_fd_pr__pfet_01v8 ad=1.9812 pd=10.94 as=0 ps=0 w=5.08 l=3.15
X103 a_n8335_8538.t0 VP.t3 a_n1578_n2628.t5 GND.t4 sky130_fd_pr__nfet_01v8 ad=1.3104 pd=7.5 as=1.3104 ps=7.5 w=3.36 l=6.01
X104 a_n12120_6849.t4 a_n8335_8538.t33 a_n5434_7417.t16 VDD.t93 sky130_fd_pr__pfet_01v8 ad=0.46035 pd=3.12 as=0.46035 ps=3.12 w=2.79 l=4.28
X105 GND.t35 CS_BIAS.t40 VOUT.t15 GND.t5 sky130_fd_pr__nfet_01v8 ad=0.936 pd=5.58 as=0.396 ps=2.73 w=2.4 l=3.51
X106 a_8541_8735# a_8541_8735# a_8541_8735# VDD.t71 sky130_fd_pr__pfet_01v8 ad=1.0881 pd=6.36 as=2.1762 ps=12.72 w=2.79 l=4.28
X107 DIFFPAIR_BIAS.t1 DIFFPAIR_BIAS.t0 a_n4284_n2628.t2 GND.t162 sky130_fd_pr__nfet_01v8 ad=1.7862 pd=9.94 as=1.7862 ps=9.94 w=4.58 l=5.91
X108 VOUT.t14 CS_BIAS.t41 GND.t36 GND.t9 sky130_fd_pr__nfet_01v8 ad=0.396 pd=2.73 as=0.396 ps=2.73 w=2.4 l=3.51
X109 a_n8413_8735.t3 a_n8335_8538.t34 VDD.t92 VDD.t91 sky130_fd_pr__pfet_01v8 ad=0.46035 pd=3.12 as=0.46035 ps=3.12 w=2.79 l=4.28
X110 GND.t16 CS_BIAS.t42 VOUT.t13 GND.t15 sky130_fd_pr__nfet_01v8 ad=0.396 pd=2.73 as=0.396 ps=2.73 w=2.4 l=3.51
X111 a_n5434_7417.t14 a_n8335_8538.t35 a_n12120_6849.t3 VDD.t90 sky130_fd_pr__pfet_01v8 ad=0.46035 pd=3.12 as=0.46035 ps=3.12 w=2.79 l=4.28
X112 VDD.t14 VDD.t11 VDD.t13 VDD.t12 sky130_fd_pr__pfet_01v8 ad=1.9812 pd=10.94 as=0 ps=0 w=5.08 l=3.15
X113 VOUT.t12 CS_BIAS.t43 GND.t28 GND.t19 sky130_fd_pr__nfet_01v8 ad=0.396 pd=2.73 as=0.396 ps=2.73 w=2.4 l=3.51
X114 DIFFPAIR_BIAS.t3 DIFFPAIR_BIAS.t2 a_n4284_n2628.t1 GND.t161 sky130_fd_pr__nfet_01v8 ad=1.7862 pd=9.94 as=1.7862 ps=9.94 w=4.58 l=5.91
X115 VOUT.t11 CS_BIAS.t44 GND.t31 GND.t21 sky130_fd_pr__nfet_01v8 ad=0.396 pd=2.73 as=0.936 ps=5.58 w=2.4 l=3.51
X116 GND.t13 CS_BIAS.t45 VOUT.t10 GND.t12 sky130_fd_pr__nfet_01v8 ad=0.936 pd=5.58 as=0.396 ps=2.73 w=2.4 l=3.51
X117 VDD.t89 a_n8335_8538.t36 a_n8413_8735.t2 VDD.t88 sky130_fd_pr__pfet_01v8 ad=0.46035 pd=3.12 as=1.0881 ps=6.36 w=2.79 l=4.28
X118 VOUT.t42 a_n12120_6849.t15 VDD.t73 VDD.t72 sky130_fd_pr__pfet_01v8 ad=1.9812 pd=10.94 as=1.9812 ps=10.94 w=5.08 l=3.15
X119 a_n12120_6849.t2 a_n8335_8538.t37 a_n5434_7417.t3 VDD.t87 sky130_fd_pr__pfet_01v8 ad=0.46035 pd=3.12 as=1.0881 ps=6.36 w=2.79 l=4.28
X120 GND.t86 GND.t84 GND.t85 GND.t59 sky130_fd_pr__nfet_01v8 ad=0.936 pd=5.58 as=0 ps=0 w=2.4 l=3.51
X121 GND.t83 GND.t80 GND.t82 GND.t81 sky130_fd_pr__nfet_01v8 ad=1.7862 pd=9.94 as=0 ps=0 w=4.58 l=5.91
X122 VDD.t10 VDD.t7 VDD.t9 VDD.t8 sky130_fd_pr__pfet_01v8 ad=1.9812 pd=10.94 as=0 ps=0 w=5.08 l=3.15
X123 VOUT.t49 a_n5434_7417.t0 sky130_fd_pr__cap_mim_m3_1 l=9.91 w=17.88
X124 GND.t26 CS_BIAS.t46 VOUT.t9 GND.t5 sky130_fd_pr__nfet_01v8 ad=0.936 pd=5.58 as=0.396 ps=2.73 w=2.4 l=3.51
X125 VOUT.t8 CS_BIAS.t47 GND.t8 GND.t2 sky130_fd_pr__nfet_01v8 ad=0.396 pd=2.73 as=0.936 ps=5.58 w=2.4 l=3.51
X126 GND.t43 CS_BIAS.t48 VOUT.t7 GND.t15 sky130_fd_pr__nfet_01v8 ad=0.396 pd=2.73 as=0.396 ps=2.73 w=2.4 l=3.51
X127 GND.t23 CS_BIAS.t49 VOUT.t6 GND.t15 sky130_fd_pr__nfet_01v8 ad=0.396 pd=2.73 as=0.396 ps=2.73 w=2.4 l=3.51
X128 GND.t79 GND.t76 GND.t78 GND.t77 sky130_fd_pr__nfet_01v8 ad=0.936 pd=5.58 as=0 ps=0 w=2.4 l=3.51
X129 GND.t27 CS_BIAS.t50 VOUT.t5 GND.t5 sky130_fd_pr__nfet_01v8 ad=0.936 pd=5.58 as=0.396 ps=2.73 w=2.4 l=3.51
X130 GND.t75 GND.t72 GND.t74 GND.t73 sky130_fd_pr__nfet_01v8 ad=1.3104 pd=7.5 as=0 ps=0 w=3.36 l=6.01
X131 GND.t171 CS_BIAS.t51 VOUT.t4 GND.t12 sky130_fd_pr__nfet_01v8 ad=0.936 pd=5.58 as=0.396 ps=2.73 w=2.4 l=3.51
X132 GND.t71 GND.t69 VN.t0 GND.t70 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X133 a_n5434_7417.t5 a_n8335_8538.t38 VDD.t86 VDD.t85 sky130_fd_pr__pfet_01v8 ad=1.0881 pd=6.36 as=0.46035 ps=3.12 w=2.79 l=4.28
X134 a_n1578_n2628.t2 DIFFPAIR_BIAS.t7 a_n2838_n2628.t1 GND.t158 sky130_fd_pr__nfet_01v8 ad=1.7862 pd=9.94 as=1.7862 ps=9.94 w=4.58 l=5.91
X135 VOUT.t3 CS_BIAS.t52 GND.t30 GND.t19 sky130_fd_pr__nfet_01v8 ad=0.396 pd=2.73 as=0.396 ps=2.73 w=2.4 l=3.51
X136 CS_BIAS.t7 CS_BIAS.t6 GND.t10 GND.t9 sky130_fd_pr__nfet_01v8 ad=0.396 pd=2.73 as=0.396 ps=2.73 w=2.4 l=3.51
X137 GND.t68 GND.t66 GND.t67 GND.t59 sky130_fd_pr__nfet_01v8 ad=0.936 pd=5.58 as=0 ps=0 w=2.4 l=3.51
X138 CS_BIAS.t5 CS_BIAS.t4 GND.t33 GND.t19 sky130_fd_pr__nfet_01v8 ad=0.396 pd=2.73 as=0.396 ps=2.73 w=2.4 l=3.51
X139 CS_BIAS.t3 CS_BIAS.t2 GND.t44 GND.t21 sky130_fd_pr__nfet_01v8 ad=0.396 pd=2.73 as=0.936 ps=5.58 w=2.4 l=3.51
X140 GND.t65 GND.t62 GND.t64 GND.t63 sky130_fd_pr__nfet_01v8 ad=0.936 pd=5.58 as=0 ps=0 w=2.4 l=3.51
X141 a_n8413_8735.t1 a_n8335_8538.t39 VDD.t84 VDD.t83 sky130_fd_pr__pfet_01v8 ad=1.0881 pd=6.36 as=0.46035 ps=3.12 w=2.79 l=4.28
X142 a_n1578_n2628.t1 DIFFPAIR_BIAS.t8 a_n2838_n2628.t0 GND.t157 sky130_fd_pr__nfet_01v8 ad=1.7862 pd=9.94 as=1.7862 ps=9.94 w=4.58 l=5.91
X143 GND.t61 GND.t58 GND.t60 GND.t59 sky130_fd_pr__nfet_01v8 ad=0.936 pd=5.58 as=0 ps=0 w=2.4 l=3.51
X144 VOUT.t2 CS_BIAS.t53 GND.t45 GND.t2 sky130_fd_pr__nfet_01v8 ad=0.396 pd=2.73 as=0.936 ps=5.58 w=2.4 l=3.51
X145 GND.t57 GND.t55 GND.t56 GND.t52 sky130_fd_pr__nfet_01v8 ad=0.936 pd=5.58 as=0 ps=0 w=2.4 l=3.51
X146 GND.t54 GND.t51 GND.t53 GND.t52 sky130_fd_pr__nfet_01v8 ad=0.936 pd=5.58 as=0 ps=0 w=2.4 l=3.51
X147 VOUT.t1 CS_BIAS.t54 GND.t20 GND.t19 sky130_fd_pr__nfet_01v8 ad=0.396 pd=2.73 as=0.396 ps=2.73 w=2.4 l=3.51
X148 a_n8413_8735.t8 a_n8335_8538.t9 a_n8335_8538.t10 VDD.t82 sky130_fd_pr__pfet_01v8 ad=0.46035 pd=3.12 as=1.0881 ps=6.36 w=2.79 l=4.28
X149 GND.t50 GND.t47 GND.t49 GND.t48 sky130_fd_pr__nfet_01v8 ad=1.3104 pd=7.5 as=0 ps=0 w=3.36 l=6.01
X150 DIFFPAIR_BIAS.t5 DIFFPAIR_BIAS.t4 a_n4284_n2628.t0 GND.t160 sky130_fd_pr__nfet_01v8 ad=1.7862 pd=9.94 as=1.7862 ps=9.94 w=4.58 l=5.91
X151 GND.t37 CS_BIAS.t0 CS_BIAS.t1 GND.t15 sky130_fd_pr__nfet_01v8 ad=0.396 pd=2.73 as=0.396 ps=2.73 w=2.4 l=3.51
X152 VOUT.t0 CS_BIAS.t55 GND.t172 GND.t21 sky130_fd_pr__nfet_01v8 ad=0.396 pd=2.73 as=0.936 ps=5.58 w=2.4 l=3.51
X153 VDD.t6 VDD.t3 VDD.t5 VDD.t4 sky130_fd_pr__pfet_01v8 ad=1.0881 pd=6.36 as=0 ps=0 w=2.79 l=4.28
X154 a_n5434_7417.t4 a_n8335_8538.t40 VDD.t81 VDD.t80 sky130_fd_pr__pfet_01v8 ad=0.46035 pd=3.12 as=0.46035 ps=3.12 w=2.79 l=4.28
X155 a_n8413_8735.t6 a_n8335_8538.t41 VDD.t79 VDD.t78 sky130_fd_pr__pfet_01v8 ad=0.46035 pd=3.12 as=0.46035 ps=3.12 w=2.79 l=4.28
R0 a_n8335_8538.n8 a_n8335_8538.t16 137.597
R1 a_n8335_8538.n7 a_n8335_8538.t10 137.597
R2 a_n8335_8538.n7 a_n8335_8538.t8 133.624
R3 a_n8335_8538.n8 a_n8335_8538.t12 133.624
R4 a_n8335_8538.n7 a_n8335_8538.t14 121.974
R5 a_n8335_8538.t4 a_n8335_8538.n8 121.974
R6 a_n8335_8538.n10 a_n8335_8538.t17 164.629
R7 a_n8335_8538.n10 a_n8335_8538.t0 128.333
R8 a_n8335_8538.n0 a_n8335_8538.n10 25.3229
R9 a_n8335_8538.n6 a_n8335_8538.n5 4.17479
R10 a_n8335_8538.n4 a_n8335_8538.n3 4.17479
R11 a_n8335_8538.n0 a_n8335_8538.t31 47.7962
R12 a_n8335_8538.n0 a_n8335_8538.t33 45.3884
R13 a_n8335_8538.n0 a_n8335_8538.t35 50.0379
R14 a_n8335_8538.n0 a_n8335_8538.t37 48.5131
R15 a_n8335_8538.n0 a_n8335_8538.t7 47.7962
R16 a_n8335_8538.n0 a_n8335_8538.t13 45.4802
R17 a_n8335_8538.n0 a_n8335_8538.t5 49.8889
R18 a_n8335_8538.n0 a_n8335_8538.t9 48.5131
R19 a_n8335_8538.n5 a_n8335_8538.t15 47.7962
R20 a_n8335_8538.n6 a_n8335_8538.t1 45.1247
R21 a_n8335_8538.n6 a_n8335_8538.t3 50.5896
R22 a_n8335_8538.n5 a_n8335_8538.t11 48.5131
R23 a_n8335_8538.n3 a_n8335_8538.t30 47.7962
R24 a_n8335_8538.n4 a_n8335_8538.t26 45.1247
R25 a_n8335_8538.n4 a_n8335_8538.t27 50.5896
R26 a_n8335_8538.n3 a_n8335_8538.t29 48.5131
R27 a_n8335_8538.n2 a_n8335_8538.t39 47.7962
R28 a_n8335_8538.n2 a_n8335_8538.t20 50.055
R29 a_n8335_8538.n2 a_n8335_8538.t41 45.3153
R30 a_n8335_8538.n2 a_n8335_8538.t19 48.5131
R31 a_n8335_8538.n2 a_n8335_8538.t22 47.7962
R32 a_n8335_8538.n2 a_n8335_8538.t32 45.6221
R33 a_n8335_8538.n2 a_n8335_8538.t34 45.9309
R34 a_n8335_8538.n2 a_n8335_8538.t36 51.2945
R35 a_n8335_8538.n2 a_n8335_8538.t38 47.7962
R36 a_n8335_8538.n2 a_n8335_8538.t18 46.1614
R37 a_n8335_8538.n2 a_n8335_8538.t40 45.6975
R38 a_n8335_8538.n2 a_n8335_8538.t23 51.3208
R39 a_n8335_8538.n2 a_n8335_8538.t28 47.7962
R40 a_n8335_8538.n2 a_n8335_8538.t25 45.9354
R41 a_n8335_8538.n2 a_n8335_8538.t24 48.9242
R42 a_n8335_8538.n2 a_n8335_8538.t21 48.4558
R43 a_n8335_8538.n9 a_n8335_8538.n0 29.1706
R44 a_n8335_8538.n2 a_n8335_8538.n1 24.3765
R45 a_n8335_8538.n9 a_n8335_8538.n2 22.144
R46 a_n8335_8538.n0 a_n8335_8538.n1 15.5174
R47 a_n8335_8538.n3 a_n8335_8538.n9 15.5022
R48 a_n8335_8538.n1 a_n8335_8538.n5 13.0591
R49 a_n8335_8538.t14 a_n8335_8538.t6 11.651
R50 a_n8335_8538.t2 a_n8335_8538.t4 11.651
R51 a_n8335_8538.n5 a_n8335_8538.n3 7.67445
R52 a_n8335_8538.n8 a_n8335_8538.n1 18.934
R53 a_n8335_8538.n9 a_n8335_8538.n7 17.5048
R54 a_n8413_8735.n12 a_n8413_8735.n11 142.626
R55 a_n8413_8735.n3 a_n8413_8735.n1 140.024
R56 a_n8413_8735.n3 a_n8413_8735.n2 138.653
R57 a_n8413_8735.n11 a_n8413_8735.n10 138.651
R58 a_n8413_8735.n5 a_n8413_8735.t7 137.597
R59 a_n8413_8735.n8 a_n8413_8735.t4 133.624
R60 a_n8413_8735.n0 a_n8413_8735.t1 133.624
R61 a_n8413_8735.n0 a_n8413_8735.t2 133.624
R62 a_n8413_8735.n7 a_n8413_8735.n6 121.974
R63 a_n8413_8735.n5 a_n8413_8735.n4 121.974
R64 a_n8413_8735.n9 a_n8413_8735.n3 31.9198
R65 a_n8413_8735.n11 a_n8413_8735.n9 18.4285
R66 a_n8413_8735.n10 a_n8413_8735.t11 11.651
R67 a_n8413_8735.n10 a_n8413_8735.t12 11.651
R68 a_n8413_8735.n6 a_n8413_8735.t0 11.651
R69 a_n8413_8735.n6 a_n8413_8735.t6 11.651
R70 a_n8413_8735.n4 a_n8413_8735.t5 11.651
R71 a_n8413_8735.n4 a_n8413_8735.t3 11.651
R72 a_n8413_8735.n2 a_n8413_8735.t15 11.651
R73 a_n8413_8735.n2 a_n8413_8735.t8 11.651
R74 a_n8413_8735.n1 a_n8413_8735.t10 11.651
R75 a_n8413_8735.n1 a_n8413_8735.t13 11.651
R76 a_n8413_8735.t14 a_n8413_8735.n12 11.651
R77 a_n8413_8735.n12 a_n8413_8735.t9 11.651
R78 a_n8413_8735.n9 a_n8413_8735.n8 7.46817
R79 a_n8413_8735.n7 a_n8413_8735.n0 4.99188
R80 a_n8413_8735.n0 a_n8413_8735.n5 3.97464
R81 a_n8413_8735.n8 a_n8413_8735.n7 3.97464
R82 VDD.n2679 VDD.n59 447.805
R83 VDD.n2951 VDD.n2768 447.805
R84 VDD.n2860 VDD.n2770 447.805
R85 VDD.n2683 VDD.n61 447.805
R86 VDD.n1333 VDD.n973 447.805
R87 VDD.n1336 VDD.n1335 447.805
R88 VDD.n1207 VDD.n1050 447.805
R89 VDD.n1209 VDD.n1048 447.805
R90 VDD.n2566 VDD.n141 289.757
R91 VDD.n2541 VDD.n156 289.757
R92 VDD.n2218 VDD.n2217 289.757
R93 VDD.n2245 VDD.n417 289.757
R94 VDD.n1908 VDD.n440 289.757
R95 VDD.n1880 VDD.n1879 289.757
R96 VDD.n1539 VDD.n1538 289.757
R97 VDD.n1566 VDD.n721 289.757
R98 VDD.n2519 VDD.n2518 289.757
R99 VDD.n2576 VDD.n133 289.757
R100 VDD.n2082 VDD.n1923 289.757
R101 VDD.n2249 VDD.n421 289.757
R102 VDD.n1865 VDD.n1864 289.757
R103 VDD.n1833 VDD.n432 289.757
R104 VDD.n933 VDD.n737 289.757
R105 VDD.n791 VDD.n717 289.757
R106 VDD.n745 VDD.t71 254.689
R107 VDD.n2681 VDD.t75 254.689
R108 VDD.n1052 VDD.t65 247.615
R109 VDD.n1069 VDD.t68 247.615
R110 VDD.n1086 VDD.t44 247.615
R111 VDD.n1338 VDD.t38 247.615
R112 VDD.n776 VDD.t41 247.615
R113 VDD.n750 VDD.t15 247.615
R114 VDD.n2862 VDD.t29 247.615
R115 VDD.n2822 VDD.t32 247.615
R116 VDD.n2805 VDD.t11 247.615
R117 VDD.n115 VDD.t23 247.615
R118 VDD.n2655 VDD.t7 247.615
R119 VDD.n64 VDD.t26 247.615
R120 VDD.n806 VDD.t22 231.37
R121 VDD.n461 VDD.t56 231.37
R122 VDD.n1403 VDD.t37 231.37
R123 VDD.n443 VDD.t50 231.37
R124 VDD.n1924 VDD.t64 231.37
R125 VDD.n151 VDD.t5 231.37
R126 VDD.n2085 VDD.t61 231.37
R127 VDD.n128 VDD.t53 231.37
R128 VDD.n806 VDD.t19 225.387
R129 VDD.n461 VDD.t55 225.387
R130 VDD.n1403 VDD.t35 225.387
R131 VDD.n443 VDD.t48 225.387
R132 VDD.n1924 VDD.t62 225.387
R133 VDD.n151 VDD.t3 225.387
R134 VDD.n2085 VDD.t58 225.387
R135 VDD.n128 VDD.t52 225.387
R136 VDD.t71 VDD.t98 222.656
R137 VDD.t114 VDD.t75 222.656
R138 VDD.n1052 VDD.t67 188.109
R139 VDD.n1069 VDD.t70 188.109
R140 VDD.n1086 VDD.t47 188.109
R141 VDD.n1338 VDD.t39 188.109
R142 VDD.n776 VDD.t42 188.109
R143 VDD.n750 VDD.t17 188.109
R144 VDD.n2862 VDD.t30 188.109
R145 VDD.n2822 VDD.t33 188.109
R146 VDD.n2805 VDD.t13 188.109
R147 VDD.n115 VDD.t25 188.109
R148 VDD.n2655 VDD.t10 188.109
R149 VDD.n64 VDD.t28 188.109
R150 VDD.n2520 VDD.n2519 185
R151 VDD.n2519 VDD.n138 185
R152 VDD.n2521 VDD.n139 185
R153 VDD.n2571 VDD.n139 185
R154 VDD.n2523 VDD.n2522 185
R155 VDD.n2522 VDD.n136 185
R156 VDD.n2524 VDD.n161 185
R157 VDD.n2534 VDD.n161 185
R158 VDD.n2525 VDD.n169 185
R159 VDD.n169 VDD.n159 185
R160 VDD.n2527 VDD.n2526 185
R161 VDD.n2528 VDD.n2527 185
R162 VDD.n2503 VDD.n168 185
R163 VDD.n168 VDD.n165 185
R164 VDD.n2502 VDD.n2501 185
R165 VDD.n2501 VDD.n2500 185
R166 VDD.n171 VDD.n170 185
R167 VDD.n180 VDD.n171 185
R168 VDD.n2493 VDD.n2492 185
R169 VDD.n2494 VDD.n2493 185
R170 VDD.n2491 VDD.n181 185
R171 VDD.n181 VDD.n177 185
R172 VDD.n2490 VDD.n2489 185
R173 VDD.n2489 VDD.n2488 185
R174 VDD.n183 VDD.n182 185
R175 VDD.n184 VDD.n183 185
R176 VDD.n2481 VDD.n2480 185
R177 VDD.n2482 VDD.n2481 185
R178 VDD.n2479 VDD.n193 185
R179 VDD.n193 VDD.n190 185
R180 VDD.n2478 VDD.n2477 185
R181 VDD.n2477 VDD.n2476 185
R182 VDD.n195 VDD.n194 185
R183 VDD.n196 VDD.n195 185
R184 VDD.n2469 VDD.n2468 185
R185 VDD.n2470 VDD.n2469 185
R186 VDD.n2467 VDD.n205 185
R187 VDD.n205 VDD.n202 185
R188 VDD.n2466 VDD.n2465 185
R189 VDD.n2465 VDD.n2464 185
R190 VDD.n207 VDD.n206 185
R191 VDD.n208 VDD.n207 185
R192 VDD.n2457 VDD.n2456 185
R193 VDD.n2458 VDD.n2457 185
R194 VDD.n2455 VDD.n216 185
R195 VDD.n222 VDD.n216 185
R196 VDD.n2454 VDD.n2453 185
R197 VDD.n2453 VDD.n2452 185
R198 VDD.n218 VDD.n217 185
R199 VDD.n219 VDD.n218 185
R200 VDD.n2445 VDD.n2444 185
R201 VDD.n2446 VDD.n2445 185
R202 VDD.n2443 VDD.n229 185
R203 VDD.n229 VDD.n226 185
R204 VDD.n2442 VDD.n2441 185
R205 VDD.n2441 VDD.n2440 185
R206 VDD.n231 VDD.n230 185
R207 VDD.n232 VDD.n231 185
R208 VDD.n2433 VDD.n2432 185
R209 VDD.n2434 VDD.n2433 185
R210 VDD.n2431 VDD.n241 185
R211 VDD.n241 VDD.n238 185
R212 VDD.n2430 VDD.n2429 185
R213 VDD.n2429 VDD.n2428 185
R214 VDD.n243 VDD.n242 185
R215 VDD.n244 VDD.n243 185
R216 VDD.n2421 VDD.n2420 185
R217 VDD.n2422 VDD.n2421 185
R218 VDD.n2419 VDD.n253 185
R219 VDD.n253 VDD.n250 185
R220 VDD.n2418 VDD.n2417 185
R221 VDD.n2417 VDD.n2416 185
R222 VDD.n255 VDD.n254 185
R223 VDD.n256 VDD.n255 185
R224 VDD.n2409 VDD.n2408 185
R225 VDD.n2410 VDD.n2409 185
R226 VDD.n2407 VDD.n265 185
R227 VDD.n265 VDD.n262 185
R228 VDD.n2406 VDD.n2405 185
R229 VDD.n2405 VDD.n2404 185
R230 VDD.n267 VDD.n266 185
R231 VDD.n268 VDD.n267 185
R232 VDD.n2397 VDD.n2396 185
R233 VDD.n2398 VDD.n2397 185
R234 VDD.n2395 VDD.n277 185
R235 VDD.n277 VDD.n274 185
R236 VDD.n2394 VDD.n2393 185
R237 VDD.n2393 VDD.n2392 185
R238 VDD.n279 VDD.n278 185
R239 VDD.n280 VDD.n279 185
R240 VDD.n2385 VDD.n2384 185
R241 VDD.n2386 VDD.n2385 185
R242 VDD.n2383 VDD.n289 185
R243 VDD.n289 VDD.n286 185
R244 VDD.n2382 VDD.n2381 185
R245 VDD.n2381 VDD.n2380 185
R246 VDD.n291 VDD.n290 185
R247 VDD.n292 VDD.n291 185
R248 VDD.n2373 VDD.n2372 185
R249 VDD.n2374 VDD.n2373 185
R250 VDD.n2371 VDD.n301 185
R251 VDD.n301 VDD.n298 185
R252 VDD.n2370 VDD.n2369 185
R253 VDD.n2369 VDD.n2368 185
R254 VDD.n303 VDD.n302 185
R255 VDD.n312 VDD.n303 185
R256 VDD.n2361 VDD.n2360 185
R257 VDD.n2362 VDD.n2361 185
R258 VDD.n2359 VDD.n313 185
R259 VDD.n313 VDD.n309 185
R260 VDD.n2358 VDD.n2357 185
R261 VDD.n2357 VDD.n2356 185
R262 VDD.n315 VDD.n314 185
R263 VDD.n324 VDD.n315 185
R264 VDD.n2349 VDD.n2348 185
R265 VDD.n2350 VDD.n2349 185
R266 VDD.n2347 VDD.n325 185
R267 VDD.n325 VDD.n321 185
R268 VDD.n2346 VDD.n2345 185
R269 VDD.n2345 VDD.n2344 185
R270 VDD.n327 VDD.n326 185
R271 VDD.n328 VDD.n327 185
R272 VDD.n2337 VDD.n2336 185
R273 VDD.n2338 VDD.n2337 185
R274 VDD.n2335 VDD.n337 185
R275 VDD.n337 VDD.n334 185
R276 VDD.n2334 VDD.n2333 185
R277 VDD.n2333 VDD.n2332 185
R278 VDD.n339 VDD.n338 185
R279 VDD.n340 VDD.n339 185
R280 VDD.n2325 VDD.n2324 185
R281 VDD.n2326 VDD.n2325 185
R282 VDD.n2323 VDD.n348 185
R283 VDD.n354 VDD.n348 185
R284 VDD.n2322 VDD.n2321 185
R285 VDD.n2321 VDD.n2320 185
R286 VDD.n350 VDD.n349 185
R287 VDD.n351 VDD.n350 185
R288 VDD.n2313 VDD.n2312 185
R289 VDD.n2314 VDD.n2313 185
R290 VDD.n2311 VDD.n360 185
R291 VDD.n366 VDD.n360 185
R292 VDD.n2310 VDD.n2309 185
R293 VDD.n2309 VDD.n2308 185
R294 VDD.n362 VDD.n361 185
R295 VDD.n363 VDD.n362 185
R296 VDD.n2301 VDD.n2300 185
R297 VDD.n2302 VDD.n2301 185
R298 VDD.n2299 VDD.n373 185
R299 VDD.n373 VDD.n370 185
R300 VDD.n2298 VDD.n2297 185
R301 VDD.n2297 VDD.n2296 185
R302 VDD.n375 VDD.n374 185
R303 VDD.n376 VDD.n375 185
R304 VDD.n2289 VDD.n2288 185
R305 VDD.n2290 VDD.n2289 185
R306 VDD.n2287 VDD.n385 185
R307 VDD.n385 VDD.n382 185
R308 VDD.n2286 VDD.n2285 185
R309 VDD.n2285 VDD.n2284 185
R310 VDD.n387 VDD.n386 185
R311 VDD.n388 VDD.n387 185
R312 VDD.n2277 VDD.n2276 185
R313 VDD.n2278 VDD.n2277 185
R314 VDD.n2275 VDD.n397 185
R315 VDD.n397 VDD.n394 185
R316 VDD.n2274 VDD.n2273 185
R317 VDD.n2273 VDD.n2272 185
R318 VDD.n399 VDD.n398 185
R319 VDD.n400 VDD.n399 185
R320 VDD.n2265 VDD.n2264 185
R321 VDD.n2266 VDD.n2265 185
R322 VDD.n2263 VDD.n409 185
R323 VDD.n409 VDD.n406 185
R324 VDD.n2262 VDD.n2261 185
R325 VDD.n2261 VDD.n2260 185
R326 VDD.n411 VDD.n410 185
R327 VDD.n412 VDD.n411 185
R328 VDD.n2253 VDD.n2252 185
R329 VDD.n2254 VDD.n2253 185
R330 VDD.n2251 VDD.n421 185
R331 VDD.n421 VDD.n418 185
R332 VDD.n2250 VDD.n2249 185
R333 VDD.n423 VDD.n422 185
R334 VDD.n1927 VDD.n1926 185
R335 VDD.n1929 VDD.n1928 185
R336 VDD.n1931 VDD.n1930 185
R337 VDD.n1933 VDD.n1932 185
R338 VDD.n1935 VDD.n1934 185
R339 VDD.n1937 VDD.n1936 185
R340 VDD.n1939 VDD.n1938 185
R341 VDD.n1941 VDD.n1940 185
R342 VDD.n1943 VDD.n1942 185
R343 VDD.n1945 VDD.n1944 185
R344 VDD.n1947 VDD.n1946 185
R345 VDD.n1949 VDD.n1922 185
R346 VDD.n2082 VDD.n2081 185
R347 VDD.n2247 VDD.n2082 185
R348 VDD.n2576 VDD.n2575 185
R349 VDD.n2578 VDD.n132 185
R350 VDD.n2580 VDD.n2579 185
R351 VDD.n2581 VDD.n127 185
R352 VDD.n2583 VDD.n2582 185
R353 VDD.n2585 VDD.n126 185
R354 VDD.n2586 VDD.n123 185
R355 VDD.n2589 VDD.n2588 185
R356 VDD.n124 VDD.n122 185
R357 VDD.n2510 VDD.n2507 185
R358 VDD.n2512 VDD.n2511 185
R359 VDD.n2513 VDD.n2506 185
R360 VDD.n2515 VDD.n2514 185
R361 VDD.n2517 VDD.n2505 185
R362 VDD.n2518 VDD.n2504 185
R363 VDD.n2518 VDD.n125 185
R364 VDD.n2574 VDD.n133 185
R365 VDD.n138 VDD.n133 185
R366 VDD.n2573 VDD.n2572 185
R367 VDD.n2572 VDD.n2571 185
R368 VDD.n135 VDD.n134 185
R369 VDD.n136 VDD.n135 185
R370 VDD.n1950 VDD.n160 185
R371 VDD.n2534 VDD.n160 185
R372 VDD.n1952 VDD.n1951 185
R373 VDD.n1951 VDD.n159 185
R374 VDD.n1953 VDD.n167 185
R375 VDD.n2528 VDD.n167 185
R376 VDD.n1955 VDD.n1954 185
R377 VDD.n1954 VDD.n165 185
R378 VDD.n1956 VDD.n173 185
R379 VDD.n2500 VDD.n173 185
R380 VDD.n1958 VDD.n1957 185
R381 VDD.n1957 VDD.n180 185
R382 VDD.n1959 VDD.n179 185
R383 VDD.n2494 VDD.n179 185
R384 VDD.n1961 VDD.n1960 185
R385 VDD.n1960 VDD.n177 185
R386 VDD.n1962 VDD.n186 185
R387 VDD.n2488 VDD.n186 185
R388 VDD.n1964 VDD.n1963 185
R389 VDD.n1963 VDD.n184 185
R390 VDD.n1965 VDD.n192 185
R391 VDD.n2482 VDD.n192 185
R392 VDD.n1967 VDD.n1966 185
R393 VDD.n1966 VDD.n190 185
R394 VDD.n1968 VDD.n198 185
R395 VDD.n2476 VDD.n198 185
R396 VDD.n1970 VDD.n1969 185
R397 VDD.n1969 VDD.n196 185
R398 VDD.n1971 VDD.n204 185
R399 VDD.n2470 VDD.n204 185
R400 VDD.n1973 VDD.n1972 185
R401 VDD.n1972 VDD.n202 185
R402 VDD.n1974 VDD.n210 185
R403 VDD.n2464 VDD.n210 185
R404 VDD.n1976 VDD.n1975 185
R405 VDD.n1975 VDD.n208 185
R406 VDD.n1977 VDD.n215 185
R407 VDD.n2458 VDD.n215 185
R408 VDD.n1979 VDD.n1978 185
R409 VDD.n1978 VDD.n222 185
R410 VDD.n1980 VDD.n221 185
R411 VDD.n2452 VDD.n221 185
R412 VDD.n1982 VDD.n1981 185
R413 VDD.n1981 VDD.n219 185
R414 VDD.n1983 VDD.n228 185
R415 VDD.n2446 VDD.n228 185
R416 VDD.n1985 VDD.n1984 185
R417 VDD.n1984 VDD.n226 185
R418 VDD.n1986 VDD.n234 185
R419 VDD.n2440 VDD.n234 185
R420 VDD.n1988 VDD.n1987 185
R421 VDD.n1987 VDD.n232 185
R422 VDD.n1989 VDD.n240 185
R423 VDD.n2434 VDD.n240 185
R424 VDD.n1991 VDD.n1990 185
R425 VDD.n1990 VDD.n238 185
R426 VDD.n1992 VDD.n246 185
R427 VDD.n2428 VDD.n246 185
R428 VDD.n1994 VDD.n1993 185
R429 VDD.n1993 VDD.n244 185
R430 VDD.n1995 VDD.n252 185
R431 VDD.n2422 VDD.n252 185
R432 VDD.n1997 VDD.n1996 185
R433 VDD.n1996 VDD.n250 185
R434 VDD.n1998 VDD.n258 185
R435 VDD.n2416 VDD.n258 185
R436 VDD.n2000 VDD.n1999 185
R437 VDD.n1999 VDD.n256 185
R438 VDD.n2001 VDD.n264 185
R439 VDD.n2410 VDD.n264 185
R440 VDD.n2003 VDD.n2002 185
R441 VDD.n2002 VDD.n262 185
R442 VDD.n2004 VDD.n270 185
R443 VDD.n2404 VDD.n270 185
R444 VDD.n2006 VDD.n2005 185
R445 VDD.n2005 VDD.n268 185
R446 VDD.n2007 VDD.n276 185
R447 VDD.n2398 VDD.n276 185
R448 VDD.n2009 VDD.n2008 185
R449 VDD.n2008 VDD.n274 185
R450 VDD.n2010 VDD.n282 185
R451 VDD.n2392 VDD.n282 185
R452 VDD.n2012 VDD.n2011 185
R453 VDD.n2011 VDD.n280 185
R454 VDD.n2013 VDD.n288 185
R455 VDD.n2386 VDD.n288 185
R456 VDD.n2015 VDD.n2014 185
R457 VDD.n2014 VDD.n286 185
R458 VDD.n2016 VDD.n294 185
R459 VDD.n2380 VDD.n294 185
R460 VDD.n2018 VDD.n2017 185
R461 VDD.n2017 VDD.n292 185
R462 VDD.n2019 VDD.n300 185
R463 VDD.n2374 VDD.n300 185
R464 VDD.n2021 VDD.n2020 185
R465 VDD.n2020 VDD.n298 185
R466 VDD.n2022 VDD.n305 185
R467 VDD.n2368 VDD.n305 185
R468 VDD.n2024 VDD.n2023 185
R469 VDD.n2023 VDD.n312 185
R470 VDD.n2025 VDD.n311 185
R471 VDD.n2362 VDD.n311 185
R472 VDD.n2027 VDD.n2026 185
R473 VDD.n2026 VDD.n309 185
R474 VDD.n2028 VDD.n317 185
R475 VDD.n2356 VDD.n317 185
R476 VDD.n2030 VDD.n2029 185
R477 VDD.n2029 VDD.n324 185
R478 VDD.n2031 VDD.n323 185
R479 VDD.n2350 VDD.n323 185
R480 VDD.n2033 VDD.n2032 185
R481 VDD.n2032 VDD.n321 185
R482 VDD.n2034 VDD.n330 185
R483 VDD.n2344 VDD.n330 185
R484 VDD.n2036 VDD.n2035 185
R485 VDD.n2035 VDD.n328 185
R486 VDD.n2037 VDD.n336 185
R487 VDD.n2338 VDD.n336 185
R488 VDD.n2039 VDD.n2038 185
R489 VDD.n2038 VDD.n334 185
R490 VDD.n2040 VDD.n342 185
R491 VDD.n2332 VDD.n342 185
R492 VDD.n2042 VDD.n2041 185
R493 VDD.n2041 VDD.n340 185
R494 VDD.n2043 VDD.n347 185
R495 VDD.n2326 VDD.n347 185
R496 VDD.n2045 VDD.n2044 185
R497 VDD.n2044 VDD.n354 185
R498 VDD.n2046 VDD.n353 185
R499 VDD.n2320 VDD.n353 185
R500 VDD.n2048 VDD.n2047 185
R501 VDD.n2047 VDD.n351 185
R502 VDD.n2049 VDD.n359 185
R503 VDD.n2314 VDD.n359 185
R504 VDD.n2051 VDD.n2050 185
R505 VDD.n2050 VDD.n366 185
R506 VDD.n2052 VDD.n365 185
R507 VDD.n2308 VDD.n365 185
R508 VDD.n2054 VDD.n2053 185
R509 VDD.n2053 VDD.n363 185
R510 VDD.n2055 VDD.n372 185
R511 VDD.n2302 VDD.n372 185
R512 VDD.n2057 VDD.n2056 185
R513 VDD.n2056 VDD.n370 185
R514 VDD.n2058 VDD.n378 185
R515 VDD.n2296 VDD.n378 185
R516 VDD.n2060 VDD.n2059 185
R517 VDD.n2059 VDD.n376 185
R518 VDD.n2061 VDD.n384 185
R519 VDD.n2290 VDD.n384 185
R520 VDD.n2063 VDD.n2062 185
R521 VDD.n2062 VDD.n382 185
R522 VDD.n2064 VDD.n390 185
R523 VDD.n2284 VDD.n390 185
R524 VDD.n2066 VDD.n2065 185
R525 VDD.n2065 VDD.n388 185
R526 VDD.n2067 VDD.n396 185
R527 VDD.n2278 VDD.n396 185
R528 VDD.n2069 VDD.n2068 185
R529 VDD.n2068 VDD.n394 185
R530 VDD.n2070 VDD.n402 185
R531 VDD.n2272 VDD.n402 185
R532 VDD.n2072 VDD.n2071 185
R533 VDD.n2071 VDD.n400 185
R534 VDD.n2073 VDD.n408 185
R535 VDD.n2266 VDD.n408 185
R536 VDD.n2075 VDD.n2074 185
R537 VDD.n2074 VDD.n406 185
R538 VDD.n2076 VDD.n414 185
R539 VDD.n2260 VDD.n414 185
R540 VDD.n2078 VDD.n2077 185
R541 VDD.n2077 VDD.n412 185
R542 VDD.n2079 VDD.n420 185
R543 VDD.n2254 VDD.n420 185
R544 VDD.n2080 VDD.n1923 185
R545 VDD.n1923 VDD.n418 185
R546 VDD.n442 VDD.n440 185
R547 VDD.n440 VDD.n424 185
R548 VDD.n1876 VDD.n1875 185
R549 VDD.n1877 VDD.n1876 185
R550 VDD.n1874 VDD.n452 185
R551 VDD.n452 VDD.n449 185
R552 VDD.n1873 VDD.n1872 185
R553 VDD.n1872 VDD.n1871 185
R554 VDD.n454 VDD.n453 185
R555 VDD.n455 VDD.n454 185
R556 VDD.n1824 VDD.n1823 185
R557 VDD.n1825 VDD.n1824 185
R558 VDD.n1822 VDD.n468 185
R559 VDD.n468 VDD.n465 185
R560 VDD.n1821 VDD.n1820 185
R561 VDD.n1820 VDD.n1819 185
R562 VDD.n470 VDD.n469 185
R563 VDD.n480 VDD.n470 185
R564 VDD.n1810 VDD.n1809 185
R565 VDD.n1811 VDD.n1810 185
R566 VDD.n1808 VDD.n481 185
R567 VDD.n481 VDD.n477 185
R568 VDD.n1807 VDD.n1806 185
R569 VDD.n1806 VDD.n1805 185
R570 VDD.n483 VDD.n482 185
R571 VDD.n484 VDD.n483 185
R572 VDD.n1798 VDD.n1797 185
R573 VDD.n1799 VDD.n1798 185
R574 VDD.n1796 VDD.n493 185
R575 VDD.n493 VDD.n490 185
R576 VDD.n1795 VDD.n1794 185
R577 VDD.n1794 VDD.n1793 185
R578 VDD.n495 VDD.n494 185
R579 VDD.n496 VDD.n495 185
R580 VDD.n1786 VDD.n1785 185
R581 VDD.n1787 VDD.n1786 185
R582 VDD.n1784 VDD.n505 185
R583 VDD.n505 VDD.n502 185
R584 VDD.n1783 VDD.n1782 185
R585 VDD.n1782 VDD.n1781 185
R586 VDD.n507 VDD.n506 185
R587 VDD.n508 VDD.n507 185
R588 VDD.n1774 VDD.n1773 185
R589 VDD.n1775 VDD.n1774 185
R590 VDD.n1772 VDD.n517 185
R591 VDD.n517 VDD.n514 185
R592 VDD.n1771 VDD.n1770 185
R593 VDD.n1770 VDD.n1769 185
R594 VDD.n519 VDD.n518 185
R595 VDD.n520 VDD.n519 185
R596 VDD.n1762 VDD.n1761 185
R597 VDD.n1763 VDD.n1762 185
R598 VDD.n1760 VDD.n529 185
R599 VDD.n529 VDD.n526 185
R600 VDD.n1759 VDD.n1758 185
R601 VDD.n1758 VDD.n1757 185
R602 VDD.n531 VDD.n530 185
R603 VDD.n532 VDD.n531 185
R604 VDD.n1750 VDD.n1749 185
R605 VDD.n1751 VDD.n1750 185
R606 VDD.n1748 VDD.n541 185
R607 VDD.n541 VDD.n538 185
R608 VDD.n1747 VDD.n1746 185
R609 VDD.n1746 VDD.n1745 185
R610 VDD.n543 VDD.n542 185
R611 VDD.n544 VDD.n543 185
R612 VDD.n1738 VDD.n1737 185
R613 VDD.n1739 VDD.n1738 185
R614 VDD.n1736 VDD.n553 185
R615 VDD.n553 VDD.n550 185
R616 VDD.n1735 VDD.n1734 185
R617 VDD.n1734 VDD.n1733 185
R618 VDD.n555 VDD.n554 185
R619 VDD.n556 VDD.n555 185
R620 VDD.n1726 VDD.n1725 185
R621 VDD.n1727 VDD.n1726 185
R622 VDD.n1724 VDD.n565 185
R623 VDD.n565 VDD.n562 185
R624 VDD.n1723 VDD.n1722 185
R625 VDD.n1722 VDD.n1721 185
R626 VDD.n567 VDD.n566 185
R627 VDD.n568 VDD.n567 185
R628 VDD.n1714 VDD.n1713 185
R629 VDD.n1715 VDD.n1714 185
R630 VDD.n1712 VDD.n577 185
R631 VDD.n577 VDD.n574 185
R632 VDD.n1711 VDD.n1710 185
R633 VDD.n1710 VDD.n1709 185
R634 VDD.n579 VDD.n578 185
R635 VDD.n580 VDD.n579 185
R636 VDD.n1702 VDD.n1701 185
R637 VDD.n1703 VDD.n1702 185
R638 VDD.n1700 VDD.n589 185
R639 VDD.n589 VDD.n586 185
R640 VDD.n1699 VDD.n1698 185
R641 VDD.n1698 VDD.n1697 185
R642 VDD.n591 VDD.n590 185
R643 VDD.n600 VDD.n591 185
R644 VDD.n1690 VDD.n1689 185
R645 VDD.n1691 VDD.n1690 185
R646 VDD.n1688 VDD.n601 185
R647 VDD.n601 VDD.n597 185
R648 VDD.n1687 VDD.n1686 185
R649 VDD.n1686 VDD.n1685 185
R650 VDD.n603 VDD.n602 185
R651 VDD.n612 VDD.n603 185
R652 VDD.n1678 VDD.n1677 185
R653 VDD.n1679 VDD.n1678 185
R654 VDD.n1676 VDD.n613 185
R655 VDD.n613 VDD.n609 185
R656 VDD.n1675 VDD.n1674 185
R657 VDD.n1674 VDD.n1673 185
R658 VDD.n615 VDD.n614 185
R659 VDD.n616 VDD.n615 185
R660 VDD.n1666 VDD.n1665 185
R661 VDD.n1667 VDD.n1666 185
R662 VDD.n1664 VDD.n625 185
R663 VDD.n625 VDD.n622 185
R664 VDD.n1663 VDD.n1662 185
R665 VDD.n1662 VDD.n1661 185
R666 VDD.n627 VDD.n626 185
R667 VDD.n628 VDD.n627 185
R668 VDD.n1654 VDD.n1653 185
R669 VDD.n1655 VDD.n1654 185
R670 VDD.n1652 VDD.n637 185
R671 VDD.n637 VDD.n634 185
R672 VDD.n1651 VDD.n1650 185
R673 VDD.n1650 VDD.n1649 185
R674 VDD.n639 VDD.n638 185
R675 VDD.n640 VDD.n639 185
R676 VDD.n1642 VDD.n1641 185
R677 VDD.n1643 VDD.n1642 185
R678 VDD.n1640 VDD.n648 185
R679 VDD.n654 VDD.n648 185
R680 VDD.n1639 VDD.n1638 185
R681 VDD.n1638 VDD.n1637 185
R682 VDD.n650 VDD.n649 185
R683 VDD.n651 VDD.n650 185
R684 VDD.n1630 VDD.n1629 185
R685 VDD.n1631 VDD.n1630 185
R686 VDD.n1628 VDD.n661 185
R687 VDD.n661 VDD.n658 185
R688 VDD.n1627 VDD.n1626 185
R689 VDD.n1626 VDD.n1625 185
R690 VDD.n663 VDD.n662 185
R691 VDD.n664 VDD.n663 185
R692 VDD.n1618 VDD.n1617 185
R693 VDD.n1619 VDD.n1618 185
R694 VDD.n1616 VDD.n673 185
R695 VDD.n673 VDD.n670 185
R696 VDD.n1615 VDD.n1614 185
R697 VDD.n1614 VDD.n1613 185
R698 VDD.n675 VDD.n674 185
R699 VDD.n676 VDD.n675 185
R700 VDD.n1606 VDD.n1605 185
R701 VDD.n1607 VDD.n1606 185
R702 VDD.n1604 VDD.n685 185
R703 VDD.n685 VDD.n682 185
R704 VDD.n1603 VDD.n1602 185
R705 VDD.n1602 VDD.n1601 185
R706 VDD.n687 VDD.n686 185
R707 VDD.n688 VDD.n687 185
R708 VDD.n1594 VDD.n1593 185
R709 VDD.n1595 VDD.n1594 185
R710 VDD.n1592 VDD.n697 185
R711 VDD.n697 VDD.n694 185
R712 VDD.n1591 VDD.n1590 185
R713 VDD.n1590 VDD.n1589 185
R714 VDD.n699 VDD.n698 185
R715 VDD.n700 VDD.n699 185
R716 VDD.n1582 VDD.n1581 185
R717 VDD.n1583 VDD.n1582 185
R718 VDD.n1580 VDD.n709 185
R719 VDD.n709 VDD.n706 185
R720 VDD.n1579 VDD.n1578 185
R721 VDD.n1578 VDD.n1577 185
R722 VDD.n711 VDD.n710 185
R723 VDD.n712 VDD.n711 185
R724 VDD.n1570 VDD.n1569 185
R725 VDD.n1571 VDD.n1570 185
R726 VDD.n1568 VDD.n721 185
R727 VDD.n721 VDD.n718 185
R728 VDD.n1567 VDD.n1566 185
R729 VDD.n723 VDD.n722 185
R730 VDD.n1563 VDD.n1562 185
R731 VDD.n1564 VDD.n1563 185
R732 VDD.n1561 VDD.n738 185
R733 VDD.n1560 VDD.n1559 185
R734 VDD.n1558 VDD.n1557 185
R735 VDD.n1556 VDD.n1555 185
R736 VDD.n1554 VDD.n1553 185
R737 VDD.n1552 VDD.n1551 185
R738 VDD.n1550 VDD.n1549 185
R739 VDD.n1548 VDD.n1547 185
R740 VDD.n1546 VDD.n1545 185
R741 VDD.n1544 VDD.n1543 185
R742 VDD.n1542 VDD.n1541 185
R743 VDD.n1540 VDD.n1539 185
R744 VDD.n1881 VDD.n1880 185
R745 VDD.n1883 VDD.n1882 185
R746 VDD.n1885 VDD.n1884 185
R747 VDD.n1887 VDD.n1886 185
R748 VDD.n1889 VDD.n1888 185
R749 VDD.n1891 VDD.n1890 185
R750 VDD.n1893 VDD.n1892 185
R751 VDD.n1895 VDD.n1894 185
R752 VDD.n1897 VDD.n1896 185
R753 VDD.n1899 VDD.n1898 185
R754 VDD.n1901 VDD.n1900 185
R755 VDD.n1903 VDD.n1902 185
R756 VDD.n1905 VDD.n1904 185
R757 VDD.n1906 VDD.n441 185
R758 VDD.n1908 VDD.n1907 185
R759 VDD.n1909 VDD.n1908 185
R760 VDD.n1879 VDD.n446 185
R761 VDD.n1879 VDD.n424 185
R762 VDD.n1878 VDD.n448 185
R763 VDD.n1878 VDD.n1877 185
R764 VDD.n1406 VDD.n447 185
R765 VDD.n449 VDD.n447 185
R766 VDD.n1407 VDD.n456 185
R767 VDD.n1871 VDD.n456 185
R768 VDD.n1409 VDD.n1408 185
R769 VDD.n1408 VDD.n455 185
R770 VDD.n1410 VDD.n466 185
R771 VDD.n1825 VDD.n466 185
R772 VDD.n1412 VDD.n1411 185
R773 VDD.n1411 VDD.n465 185
R774 VDD.n1413 VDD.n471 185
R775 VDD.n1819 VDD.n471 185
R776 VDD.n1415 VDD.n1414 185
R777 VDD.n1414 VDD.n480 185
R778 VDD.n1416 VDD.n478 185
R779 VDD.n1811 VDD.n478 185
R780 VDD.n1418 VDD.n1417 185
R781 VDD.n1417 VDD.n477 185
R782 VDD.n1419 VDD.n485 185
R783 VDD.n1805 VDD.n485 185
R784 VDD.n1421 VDD.n1420 185
R785 VDD.n1420 VDD.n484 185
R786 VDD.n1422 VDD.n491 185
R787 VDD.n1799 VDD.n491 185
R788 VDD.n1424 VDD.n1423 185
R789 VDD.n1423 VDD.n490 185
R790 VDD.n1425 VDD.n497 185
R791 VDD.n1793 VDD.n497 185
R792 VDD.n1427 VDD.n1426 185
R793 VDD.n1426 VDD.n496 185
R794 VDD.n1428 VDD.n503 185
R795 VDD.n1787 VDD.n503 185
R796 VDD.n1430 VDD.n1429 185
R797 VDD.n1429 VDD.n502 185
R798 VDD.n1431 VDD.n509 185
R799 VDD.n1781 VDD.n509 185
R800 VDD.n1433 VDD.n1432 185
R801 VDD.n1432 VDD.n508 185
R802 VDD.n1434 VDD.n515 185
R803 VDD.n1775 VDD.n515 185
R804 VDD.n1436 VDD.n1435 185
R805 VDD.n1435 VDD.n514 185
R806 VDD.n1437 VDD.n521 185
R807 VDD.n1769 VDD.n521 185
R808 VDD.n1439 VDD.n1438 185
R809 VDD.n1438 VDD.n520 185
R810 VDD.n1440 VDD.n527 185
R811 VDD.n1763 VDD.n527 185
R812 VDD.n1442 VDD.n1441 185
R813 VDD.n1441 VDD.n526 185
R814 VDD.n1443 VDD.n533 185
R815 VDD.n1757 VDD.n533 185
R816 VDD.n1445 VDD.n1444 185
R817 VDD.n1444 VDD.n532 185
R818 VDD.n1446 VDD.n539 185
R819 VDD.n1751 VDD.n539 185
R820 VDD.n1448 VDD.n1447 185
R821 VDD.n1447 VDD.n538 185
R822 VDD.n1449 VDD.n545 185
R823 VDD.n1745 VDD.n545 185
R824 VDD.n1451 VDD.n1450 185
R825 VDD.n1450 VDD.n544 185
R826 VDD.n1452 VDD.n551 185
R827 VDD.n1739 VDD.n551 185
R828 VDD.n1454 VDD.n1453 185
R829 VDD.n1453 VDD.n550 185
R830 VDD.n1455 VDD.n557 185
R831 VDD.n1733 VDD.n557 185
R832 VDD.n1457 VDD.n1456 185
R833 VDD.n1456 VDD.n556 185
R834 VDD.n1458 VDD.n563 185
R835 VDD.n1727 VDD.n563 185
R836 VDD.n1460 VDD.n1459 185
R837 VDD.n1459 VDD.n562 185
R838 VDD.n1461 VDD.n569 185
R839 VDD.n1721 VDD.n569 185
R840 VDD.n1463 VDD.n1462 185
R841 VDD.n1462 VDD.n568 185
R842 VDD.n1464 VDD.n575 185
R843 VDD.n1715 VDD.n575 185
R844 VDD.n1466 VDD.n1465 185
R845 VDD.n1465 VDD.n574 185
R846 VDD.n1467 VDD.n581 185
R847 VDD.n1709 VDD.n581 185
R848 VDD.n1469 VDD.n1468 185
R849 VDD.n1468 VDD.n580 185
R850 VDD.n1470 VDD.n587 185
R851 VDD.n1703 VDD.n587 185
R852 VDD.n1472 VDD.n1471 185
R853 VDD.n1471 VDD.n586 185
R854 VDD.n1473 VDD.n592 185
R855 VDD.n1697 VDD.n592 185
R856 VDD.n1475 VDD.n1474 185
R857 VDD.n1474 VDD.n600 185
R858 VDD.n1476 VDD.n598 185
R859 VDD.n1691 VDD.n598 185
R860 VDD.n1478 VDD.n1477 185
R861 VDD.n1477 VDD.n597 185
R862 VDD.n1479 VDD.n604 185
R863 VDD.n1685 VDD.n604 185
R864 VDD.n1481 VDD.n1480 185
R865 VDD.n1480 VDD.n612 185
R866 VDD.n1482 VDD.n610 185
R867 VDD.n1679 VDD.n610 185
R868 VDD.n1484 VDD.n1483 185
R869 VDD.n1483 VDD.n609 185
R870 VDD.n1485 VDD.n617 185
R871 VDD.n1673 VDD.n617 185
R872 VDD.n1487 VDD.n1486 185
R873 VDD.n1486 VDD.n616 185
R874 VDD.n1488 VDD.n623 185
R875 VDD.n1667 VDD.n623 185
R876 VDD.n1490 VDD.n1489 185
R877 VDD.n1489 VDD.n622 185
R878 VDD.n1491 VDD.n629 185
R879 VDD.n1661 VDD.n629 185
R880 VDD.n1493 VDD.n1492 185
R881 VDD.n1492 VDD.n628 185
R882 VDD.n1494 VDD.n635 185
R883 VDD.n1655 VDD.n635 185
R884 VDD.n1496 VDD.n1495 185
R885 VDD.n1495 VDD.n634 185
R886 VDD.n1497 VDD.n641 185
R887 VDD.n1649 VDD.n641 185
R888 VDD.n1499 VDD.n1498 185
R889 VDD.n1498 VDD.n640 185
R890 VDD.n1500 VDD.n646 185
R891 VDD.n1643 VDD.n646 185
R892 VDD.n1502 VDD.n1501 185
R893 VDD.n1501 VDD.n654 185
R894 VDD.n1503 VDD.n652 185
R895 VDD.n1637 VDD.n652 185
R896 VDD.n1505 VDD.n1504 185
R897 VDD.n1504 VDD.n651 185
R898 VDD.n1506 VDD.n659 185
R899 VDD.n1631 VDD.n659 185
R900 VDD.n1508 VDD.n1507 185
R901 VDD.n1507 VDD.n658 185
R902 VDD.n1509 VDD.n665 185
R903 VDD.n1625 VDD.n665 185
R904 VDD.n1511 VDD.n1510 185
R905 VDD.n1510 VDD.n664 185
R906 VDD.n1512 VDD.n671 185
R907 VDD.n1619 VDD.n671 185
R908 VDD.n1514 VDD.n1513 185
R909 VDD.n1513 VDD.n670 185
R910 VDD.n1515 VDD.n677 185
R911 VDD.n1613 VDD.n677 185
R912 VDD.n1517 VDD.n1516 185
R913 VDD.n1516 VDD.n676 185
R914 VDD.n1518 VDD.n683 185
R915 VDD.n1607 VDD.n683 185
R916 VDD.n1520 VDD.n1519 185
R917 VDD.n1519 VDD.n682 185
R918 VDD.n1521 VDD.n689 185
R919 VDD.n1601 VDD.n689 185
R920 VDD.n1523 VDD.n1522 185
R921 VDD.n1522 VDD.n688 185
R922 VDD.n1524 VDD.n695 185
R923 VDD.n1595 VDD.n695 185
R924 VDD.n1526 VDD.n1525 185
R925 VDD.n1525 VDD.n694 185
R926 VDD.n1527 VDD.n701 185
R927 VDD.n1589 VDD.n701 185
R928 VDD.n1529 VDD.n1528 185
R929 VDD.n1528 VDD.n700 185
R930 VDD.n1530 VDD.n707 185
R931 VDD.n1583 VDD.n707 185
R932 VDD.n1532 VDD.n1531 185
R933 VDD.n1531 VDD.n706 185
R934 VDD.n1533 VDD.n713 185
R935 VDD.n1577 VDD.n713 185
R936 VDD.n1535 VDD.n1534 185
R937 VDD.n1534 VDD.n712 185
R938 VDD.n1536 VDD.n719 185
R939 VDD.n1571 VDD.n719 185
R940 VDD.n1538 VDD.n1537 185
R941 VDD.n1538 VDD.n718 185
R942 VDD.n2568 VDD.n141 185
R943 VDD.n141 VDD.n138 185
R944 VDD.n2570 VDD.n2569 185
R945 VDD.n2571 VDD.n2570 185
R946 VDD.n142 VDD.n140 185
R947 VDD.n140 VDD.n136 185
R948 VDD.n2533 VDD.n2532 185
R949 VDD.n2534 VDD.n2533 185
R950 VDD.n2531 VDD.n162 185
R951 VDD.n162 VDD.n159 185
R952 VDD.n2530 VDD.n2529 185
R953 VDD.n2529 VDD.n2528 185
R954 VDD.n164 VDD.n163 185
R955 VDD.n165 VDD.n164 185
R956 VDD.n2499 VDD.n2498 185
R957 VDD.n2500 VDD.n2499 185
R958 VDD.n2497 VDD.n174 185
R959 VDD.n180 VDD.n174 185
R960 VDD.n2496 VDD.n2495 185
R961 VDD.n2495 VDD.n2494 185
R962 VDD.n176 VDD.n175 185
R963 VDD.n177 VDD.n176 185
R964 VDD.n2487 VDD.n2486 185
R965 VDD.n2488 VDD.n2487 185
R966 VDD.n2485 VDD.n187 185
R967 VDD.n187 VDD.n184 185
R968 VDD.n2484 VDD.n2483 185
R969 VDD.n2483 VDD.n2482 185
R970 VDD.n189 VDD.n188 185
R971 VDD.n190 VDD.n189 185
R972 VDD.n2475 VDD.n2474 185
R973 VDD.n2476 VDD.n2475 185
R974 VDD.n2473 VDD.n199 185
R975 VDD.n199 VDD.n196 185
R976 VDD.n2472 VDD.n2471 185
R977 VDD.n2471 VDD.n2470 185
R978 VDD.n201 VDD.n200 185
R979 VDD.n202 VDD.n201 185
R980 VDD.n2463 VDD.n2462 185
R981 VDD.n2464 VDD.n2463 185
R982 VDD.n2461 VDD.n211 185
R983 VDD.n211 VDD.n208 185
R984 VDD.n2460 VDD.n2459 185
R985 VDD.n2459 VDD.n2458 185
R986 VDD.n213 VDD.n212 185
R987 VDD.n222 VDD.n213 185
R988 VDD.n2451 VDD.n2450 185
R989 VDD.n2452 VDD.n2451 185
R990 VDD.n2449 VDD.n223 185
R991 VDD.n223 VDD.n219 185
R992 VDD.n2448 VDD.n2447 185
R993 VDD.n2447 VDD.n2446 185
R994 VDD.n225 VDD.n224 185
R995 VDD.n226 VDD.n225 185
R996 VDD.n2439 VDD.n2438 185
R997 VDD.n2440 VDD.n2439 185
R998 VDD.n2437 VDD.n235 185
R999 VDD.n235 VDD.n232 185
R1000 VDD.n2436 VDD.n2435 185
R1001 VDD.n2435 VDD.n2434 185
R1002 VDD.n237 VDD.n236 185
R1003 VDD.n238 VDD.n237 185
R1004 VDD.n2427 VDD.n2426 185
R1005 VDD.n2428 VDD.n2427 185
R1006 VDD.n2425 VDD.n247 185
R1007 VDD.n247 VDD.n244 185
R1008 VDD.n2424 VDD.n2423 185
R1009 VDD.n2423 VDD.n2422 185
R1010 VDD.n249 VDD.n248 185
R1011 VDD.n250 VDD.n249 185
R1012 VDD.n2415 VDD.n2414 185
R1013 VDD.n2416 VDD.n2415 185
R1014 VDD.n2413 VDD.n259 185
R1015 VDD.n259 VDD.n256 185
R1016 VDD.n2412 VDD.n2411 185
R1017 VDD.n2411 VDD.n2410 185
R1018 VDD.n261 VDD.n260 185
R1019 VDD.n262 VDD.n261 185
R1020 VDD.n2403 VDD.n2402 185
R1021 VDD.n2404 VDD.n2403 185
R1022 VDD.n2401 VDD.n271 185
R1023 VDD.n271 VDD.n268 185
R1024 VDD.n2400 VDD.n2399 185
R1025 VDD.n2399 VDD.n2398 185
R1026 VDD.n273 VDD.n272 185
R1027 VDD.n274 VDD.n273 185
R1028 VDD.n2391 VDD.n2390 185
R1029 VDD.n2392 VDD.n2391 185
R1030 VDD.n2389 VDD.n283 185
R1031 VDD.n283 VDD.n280 185
R1032 VDD.n2388 VDD.n2387 185
R1033 VDD.n2387 VDD.n2386 185
R1034 VDD.n285 VDD.n284 185
R1035 VDD.n286 VDD.n285 185
R1036 VDD.n2379 VDD.n2378 185
R1037 VDD.n2380 VDD.n2379 185
R1038 VDD.n2377 VDD.n295 185
R1039 VDD.n295 VDD.n292 185
R1040 VDD.n2376 VDD.n2375 185
R1041 VDD.n2375 VDD.n2374 185
R1042 VDD.n297 VDD.n296 185
R1043 VDD.n298 VDD.n297 185
R1044 VDD.n2367 VDD.n2366 185
R1045 VDD.n2368 VDD.n2367 185
R1046 VDD.n2365 VDD.n306 185
R1047 VDD.n312 VDD.n306 185
R1048 VDD.n2364 VDD.n2363 185
R1049 VDD.n2363 VDD.n2362 185
R1050 VDD.n308 VDD.n307 185
R1051 VDD.n309 VDD.n308 185
R1052 VDD.n2355 VDD.n2354 185
R1053 VDD.n2356 VDD.n2355 185
R1054 VDD.n2353 VDD.n318 185
R1055 VDD.n324 VDD.n318 185
R1056 VDD.n2352 VDD.n2351 185
R1057 VDD.n2351 VDD.n2350 185
R1058 VDD.n320 VDD.n319 185
R1059 VDD.n321 VDD.n320 185
R1060 VDD.n2343 VDD.n2342 185
R1061 VDD.n2344 VDD.n2343 185
R1062 VDD.n2341 VDD.n331 185
R1063 VDD.n331 VDD.n328 185
R1064 VDD.n2340 VDD.n2339 185
R1065 VDD.n2339 VDD.n2338 185
R1066 VDD.n333 VDD.n332 185
R1067 VDD.n334 VDD.n333 185
R1068 VDD.n2331 VDD.n2330 185
R1069 VDD.n2332 VDD.n2331 185
R1070 VDD.n2329 VDD.n343 185
R1071 VDD.n343 VDD.n340 185
R1072 VDD.n2328 VDD.n2327 185
R1073 VDD.n2327 VDD.n2326 185
R1074 VDD.n345 VDD.n344 185
R1075 VDD.n354 VDD.n345 185
R1076 VDD.n2319 VDD.n2318 185
R1077 VDD.n2320 VDD.n2319 185
R1078 VDD.n2317 VDD.n355 185
R1079 VDD.n355 VDD.n351 185
R1080 VDD.n2316 VDD.n2315 185
R1081 VDD.n2315 VDD.n2314 185
R1082 VDD.n357 VDD.n356 185
R1083 VDD.n366 VDD.n357 185
R1084 VDD.n2307 VDD.n2306 185
R1085 VDD.n2308 VDD.n2307 185
R1086 VDD.n2305 VDD.n367 185
R1087 VDD.n367 VDD.n363 185
R1088 VDD.n2304 VDD.n2303 185
R1089 VDD.n2303 VDD.n2302 185
R1090 VDD.n369 VDD.n368 185
R1091 VDD.n370 VDD.n369 185
R1092 VDD.n2295 VDD.n2294 185
R1093 VDD.n2296 VDD.n2295 185
R1094 VDD.n2293 VDD.n379 185
R1095 VDD.n379 VDD.n376 185
R1096 VDD.n2292 VDD.n2291 185
R1097 VDD.n2291 VDD.n2290 185
R1098 VDD.n381 VDD.n380 185
R1099 VDD.n382 VDD.n381 185
R1100 VDD.n2283 VDD.n2282 185
R1101 VDD.n2284 VDD.n2283 185
R1102 VDD.n2281 VDD.n391 185
R1103 VDD.n391 VDD.n388 185
R1104 VDD.n2280 VDD.n2279 185
R1105 VDD.n2279 VDD.n2278 185
R1106 VDD.n393 VDD.n392 185
R1107 VDD.n394 VDD.n393 185
R1108 VDD.n2271 VDD.n2270 185
R1109 VDD.n2272 VDD.n2271 185
R1110 VDD.n2269 VDD.n403 185
R1111 VDD.n403 VDD.n400 185
R1112 VDD.n2268 VDD.n2267 185
R1113 VDD.n2267 VDD.n2266 185
R1114 VDD.n405 VDD.n404 185
R1115 VDD.n406 VDD.n405 185
R1116 VDD.n2259 VDD.n2258 185
R1117 VDD.n2260 VDD.n2259 185
R1118 VDD.n2257 VDD.n415 185
R1119 VDD.n415 VDD.n412 185
R1120 VDD.n2256 VDD.n2255 185
R1121 VDD.n2255 VDD.n2254 185
R1122 VDD.n417 VDD.n416 185
R1123 VDD.n418 VDD.n417 185
R1124 VDD.n2245 VDD.n2244 185
R1125 VDD.n2243 VDD.n2084 185
R1126 VDD.n2242 VDD.n2083 185
R1127 VDD.n2247 VDD.n2083 185
R1128 VDD.n2241 VDD.n2240 185
R1129 VDD.n2239 VDD.n2238 185
R1130 VDD.n2237 VDD.n2236 185
R1131 VDD.n2235 VDD.n2234 185
R1132 VDD.n2233 VDD.n2232 185
R1133 VDD.n2231 VDD.n2230 185
R1134 VDD.n2229 VDD.n2228 185
R1135 VDD.n2227 VDD.n2226 185
R1136 VDD.n2225 VDD.n2224 185
R1137 VDD.n2223 VDD.n2222 185
R1138 VDD.n2221 VDD.n2220 185
R1139 VDD.n2219 VDD.n2218 185
R1140 VDD.n2541 VDD.n2540 185
R1141 VDD.n2543 VDD.n155 185
R1142 VDD.n2545 VDD.n2544 185
R1143 VDD.n2546 VDD.n150 185
R1144 VDD.n2548 VDD.n2547 185
R1145 VDD.n2550 VDD.n148 185
R1146 VDD.n2552 VDD.n2551 185
R1147 VDD.n2554 VDD.n147 185
R1148 VDD.n2556 VDD.n2555 185
R1149 VDD.n2558 VDD.n145 185
R1150 VDD.n2560 VDD.n2559 185
R1151 VDD.n2561 VDD.n144 185
R1152 VDD.n2563 VDD.n2562 185
R1153 VDD.n2565 VDD.n143 185
R1154 VDD.n2567 VDD.n2566 185
R1155 VDD.n2566 VDD.n125 185
R1156 VDD.n2539 VDD.n156 185
R1157 VDD.n156 VDD.n138 185
R1158 VDD.n2538 VDD.n137 185
R1159 VDD.n2571 VDD.n137 185
R1160 VDD.n2537 VDD.n2536 185
R1161 VDD.n2536 VDD.n136 185
R1162 VDD.n2535 VDD.n157 185
R1163 VDD.n2535 VDD.n2534 185
R1164 VDD.n2088 VDD.n158 185
R1165 VDD.n159 VDD.n158 185
R1166 VDD.n2089 VDD.n166 185
R1167 VDD.n2528 VDD.n166 185
R1168 VDD.n2091 VDD.n2090 185
R1169 VDD.n2090 VDD.n165 185
R1170 VDD.n2092 VDD.n172 185
R1171 VDD.n2500 VDD.n172 185
R1172 VDD.n2094 VDD.n2093 185
R1173 VDD.n2093 VDD.n180 185
R1174 VDD.n2095 VDD.n178 185
R1175 VDD.n2494 VDD.n178 185
R1176 VDD.n2097 VDD.n2096 185
R1177 VDD.n2096 VDD.n177 185
R1178 VDD.n2098 VDD.n185 185
R1179 VDD.n2488 VDD.n185 185
R1180 VDD.n2100 VDD.n2099 185
R1181 VDD.n2099 VDD.n184 185
R1182 VDD.n2101 VDD.n191 185
R1183 VDD.n2482 VDD.n191 185
R1184 VDD.n2103 VDD.n2102 185
R1185 VDD.n2102 VDD.n190 185
R1186 VDD.n2104 VDD.n197 185
R1187 VDD.n2476 VDD.n197 185
R1188 VDD.n2106 VDD.n2105 185
R1189 VDD.n2105 VDD.n196 185
R1190 VDD.n2107 VDD.n203 185
R1191 VDD.n2470 VDD.n203 185
R1192 VDD.n2109 VDD.n2108 185
R1193 VDD.n2108 VDD.n202 185
R1194 VDD.n2110 VDD.n209 185
R1195 VDD.n2464 VDD.n209 185
R1196 VDD.n2112 VDD.n2111 185
R1197 VDD.n2111 VDD.n208 185
R1198 VDD.n2113 VDD.n214 185
R1199 VDD.n2458 VDD.n214 185
R1200 VDD.n2115 VDD.n2114 185
R1201 VDD.n2114 VDD.n222 185
R1202 VDD.n2116 VDD.n220 185
R1203 VDD.n2452 VDD.n220 185
R1204 VDD.n2118 VDD.n2117 185
R1205 VDD.n2117 VDD.n219 185
R1206 VDD.n2119 VDD.n227 185
R1207 VDD.n2446 VDD.n227 185
R1208 VDD.n2121 VDD.n2120 185
R1209 VDD.n2120 VDD.n226 185
R1210 VDD.n2122 VDD.n233 185
R1211 VDD.n2440 VDD.n233 185
R1212 VDD.n2124 VDD.n2123 185
R1213 VDD.n2123 VDD.n232 185
R1214 VDD.n2125 VDD.n239 185
R1215 VDD.n2434 VDD.n239 185
R1216 VDD.n2127 VDD.n2126 185
R1217 VDD.n2126 VDD.n238 185
R1218 VDD.n2128 VDD.n245 185
R1219 VDD.n2428 VDD.n245 185
R1220 VDD.n2130 VDD.n2129 185
R1221 VDD.n2129 VDD.n244 185
R1222 VDD.n2131 VDD.n251 185
R1223 VDD.n2422 VDD.n251 185
R1224 VDD.n2133 VDD.n2132 185
R1225 VDD.n2132 VDD.n250 185
R1226 VDD.n2134 VDD.n257 185
R1227 VDD.n2416 VDD.n257 185
R1228 VDD.n2136 VDD.n2135 185
R1229 VDD.n2135 VDD.n256 185
R1230 VDD.n2137 VDD.n263 185
R1231 VDD.n2410 VDD.n263 185
R1232 VDD.n2139 VDD.n2138 185
R1233 VDD.n2138 VDD.n262 185
R1234 VDD.n2140 VDD.n269 185
R1235 VDD.n2404 VDD.n269 185
R1236 VDD.n2142 VDD.n2141 185
R1237 VDD.n2141 VDD.n268 185
R1238 VDD.n2143 VDD.n275 185
R1239 VDD.n2398 VDD.n275 185
R1240 VDD.n2145 VDD.n2144 185
R1241 VDD.n2144 VDD.n274 185
R1242 VDD.n2146 VDD.n281 185
R1243 VDD.n2392 VDD.n281 185
R1244 VDD.n2148 VDD.n2147 185
R1245 VDD.n2147 VDD.n280 185
R1246 VDD.n2149 VDD.n287 185
R1247 VDD.n2386 VDD.n287 185
R1248 VDD.n2151 VDD.n2150 185
R1249 VDD.n2150 VDD.n286 185
R1250 VDD.n2152 VDD.n293 185
R1251 VDD.n2380 VDD.n293 185
R1252 VDD.n2154 VDD.n2153 185
R1253 VDD.n2153 VDD.n292 185
R1254 VDD.n2155 VDD.n299 185
R1255 VDD.n2374 VDD.n299 185
R1256 VDD.n2157 VDD.n2156 185
R1257 VDD.n2156 VDD.n298 185
R1258 VDD.n2158 VDD.n304 185
R1259 VDD.n2368 VDD.n304 185
R1260 VDD.n2160 VDD.n2159 185
R1261 VDD.n2159 VDD.n312 185
R1262 VDD.n2161 VDD.n310 185
R1263 VDD.n2362 VDD.n310 185
R1264 VDD.n2163 VDD.n2162 185
R1265 VDD.n2162 VDD.n309 185
R1266 VDD.n2164 VDD.n316 185
R1267 VDD.n2356 VDD.n316 185
R1268 VDD.n2166 VDD.n2165 185
R1269 VDD.n2165 VDD.n324 185
R1270 VDD.n2167 VDD.n322 185
R1271 VDD.n2350 VDD.n322 185
R1272 VDD.n2169 VDD.n2168 185
R1273 VDD.n2168 VDD.n321 185
R1274 VDD.n2170 VDD.n329 185
R1275 VDD.n2344 VDD.n329 185
R1276 VDD.n2172 VDD.n2171 185
R1277 VDD.n2171 VDD.n328 185
R1278 VDD.n2173 VDD.n335 185
R1279 VDD.n2338 VDD.n335 185
R1280 VDD.n2175 VDD.n2174 185
R1281 VDD.n2174 VDD.n334 185
R1282 VDD.n2176 VDD.n341 185
R1283 VDD.n2332 VDD.n341 185
R1284 VDD.n2178 VDD.n2177 185
R1285 VDD.n2177 VDD.n340 185
R1286 VDD.n2179 VDD.n346 185
R1287 VDD.n2326 VDD.n346 185
R1288 VDD.n2181 VDD.n2180 185
R1289 VDD.n2180 VDD.n354 185
R1290 VDD.n2182 VDD.n352 185
R1291 VDD.n2320 VDD.n352 185
R1292 VDD.n2184 VDD.n2183 185
R1293 VDD.n2183 VDD.n351 185
R1294 VDD.n2185 VDD.n358 185
R1295 VDD.n2314 VDD.n358 185
R1296 VDD.n2187 VDD.n2186 185
R1297 VDD.n2186 VDD.n366 185
R1298 VDD.n2188 VDD.n364 185
R1299 VDD.n2308 VDD.n364 185
R1300 VDD.n2190 VDD.n2189 185
R1301 VDD.n2189 VDD.n363 185
R1302 VDD.n2191 VDD.n371 185
R1303 VDD.n2302 VDD.n371 185
R1304 VDD.n2193 VDD.n2192 185
R1305 VDD.n2192 VDD.n370 185
R1306 VDD.n2194 VDD.n377 185
R1307 VDD.n2296 VDD.n377 185
R1308 VDD.n2196 VDD.n2195 185
R1309 VDD.n2195 VDD.n376 185
R1310 VDD.n2197 VDD.n383 185
R1311 VDD.n2290 VDD.n383 185
R1312 VDD.n2199 VDD.n2198 185
R1313 VDD.n2198 VDD.n382 185
R1314 VDD.n2200 VDD.n389 185
R1315 VDD.n2284 VDD.n389 185
R1316 VDD.n2202 VDD.n2201 185
R1317 VDD.n2201 VDD.n388 185
R1318 VDD.n2203 VDD.n395 185
R1319 VDD.n2278 VDD.n395 185
R1320 VDD.n2205 VDD.n2204 185
R1321 VDD.n2204 VDD.n394 185
R1322 VDD.n2206 VDD.n401 185
R1323 VDD.n2272 VDD.n401 185
R1324 VDD.n2208 VDD.n2207 185
R1325 VDD.n2207 VDD.n400 185
R1326 VDD.n2209 VDD.n407 185
R1327 VDD.n2266 VDD.n407 185
R1328 VDD.n2211 VDD.n2210 185
R1329 VDD.n2210 VDD.n406 185
R1330 VDD.n2212 VDD.n413 185
R1331 VDD.n2260 VDD.n413 185
R1332 VDD.n2214 VDD.n2213 185
R1333 VDD.n2213 VDD.n412 185
R1334 VDD.n2215 VDD.n419 185
R1335 VDD.n2254 VDD.n419 185
R1336 VDD.n2217 VDD.n2216 185
R1337 VDD.n2217 VDD.n418 185
R1338 VDD.n1333 VDD.n1332 185
R1339 VDD.n1334 VDD.n1333 185
R1340 VDD.n974 VDD.n972 185
R1341 VDD.n972 VDD.n971 185
R1342 VDD.n1311 VDD.n1310 185
R1343 VDD.n1310 VDD.n1309 185
R1344 VDD.n977 VDD.n976 185
R1345 VDD.n978 VDD.n977 185
R1346 VDD.n1298 VDD.n1297 185
R1347 VDD.n1299 VDD.n1298 185
R1348 VDD.n987 VDD.n986 185
R1349 VDD.n986 VDD.n985 185
R1350 VDD.n1293 VDD.n1292 185
R1351 VDD.n1292 VDD.n1291 185
R1352 VDD.n990 VDD.n989 185
R1353 VDD.n991 VDD.n990 185
R1354 VDD.n1282 VDD.n1281 185
R1355 VDD.n1283 VDD.n1282 185
R1356 VDD.n999 VDD.n998 185
R1357 VDD.n998 VDD.n997 185
R1358 VDD.n1277 VDD.n1276 185
R1359 VDD.n1276 VDD.n1275 185
R1360 VDD.n1002 VDD.n1001 185
R1361 VDD.n1003 VDD.n1002 185
R1362 VDD.n1266 VDD.n1265 185
R1363 VDD.n1267 VDD.n1266 185
R1364 VDD.n1010 VDD.n1009 185
R1365 VDD.n1009 VDD.t72 185
R1366 VDD.n1258 VDD.n1257 185
R1367 VDD.n1257 VDD.n1256 185
R1368 VDD.n1013 VDD.n1012 185
R1369 VDD.n1014 VDD.n1013 185
R1370 VDD.n1247 VDD.n1246 185
R1371 VDD.n1248 VDD.n1247 185
R1372 VDD.n1022 VDD.n1021 185
R1373 VDD.n1021 VDD.n1020 185
R1374 VDD.n1242 VDD.n1241 185
R1375 VDD.n1241 VDD.n1240 185
R1376 VDD.n1025 VDD.n1024 185
R1377 VDD.n1026 VDD.n1025 185
R1378 VDD.n1231 VDD.n1230 185
R1379 VDD.n1232 VDD.n1231 185
R1380 VDD.n1034 VDD.n1033 185
R1381 VDD.n1033 VDD.n1032 185
R1382 VDD.n1226 VDD.n1225 185
R1383 VDD.n1225 VDD.n1224 185
R1384 VDD.n1037 VDD.n1036 185
R1385 VDD.n1044 VDD.n1037 185
R1386 VDD.n1215 VDD.n1214 185
R1387 VDD.n1216 VDD.n1215 185
R1388 VDD.n1046 VDD.n1045 185
R1389 VDD.n1045 VDD.n1043 185
R1390 VDD.n1210 VDD.n1209 185
R1391 VDD.n1209 VDD.n1208 185
R1392 VDD.n1099 VDD.n1048 185
R1393 VDD.n1103 VDD.n1101 185
R1394 VDD.n1104 VDD.n1098 185
R1395 VDD.n1104 VDD.n1049 185
R1396 VDD.n1107 VDD.n1106 185
R1397 VDD.n1096 VDD.n1095 185
R1398 VDD.n1112 VDD.n1111 185
R1399 VDD.n1114 VDD.n1094 185
R1400 VDD.n1117 VDD.n1116 185
R1401 VDD.n1092 VDD.n1091 185
R1402 VDD.n1122 VDD.n1121 185
R1403 VDD.n1124 VDD.n1090 185
R1404 VDD.n1127 VDD.n1126 185
R1405 VDD.n1088 VDD.n1085 185
R1406 VDD.n1132 VDD.n1131 185
R1407 VDD.n1134 VDD.n1084 185
R1408 VDD.n1137 VDD.n1136 185
R1409 VDD.n1082 VDD.n1081 185
R1410 VDD.n1142 VDD.n1141 185
R1411 VDD.n1144 VDD.n1080 185
R1412 VDD.n1147 VDD.n1146 185
R1413 VDD.n1078 VDD.n1077 185
R1414 VDD.n1153 VDD.n1152 185
R1415 VDD.n1155 VDD.n1076 185
R1416 VDD.n1156 VDD.n1073 185
R1417 VDD.n1159 VDD.n1158 185
R1418 VDD.n1075 VDD.n1071 185
R1419 VDD.n1163 VDD.n1067 185
R1420 VDD.n1165 VDD.n1164 185
R1421 VDD.n1167 VDD.n1066 185
R1422 VDD.n1170 VDD.n1169 185
R1423 VDD.n1064 VDD.n1063 185
R1424 VDD.n1175 VDD.n1174 185
R1425 VDD.n1177 VDD.n1062 185
R1426 VDD.n1180 VDD.n1179 185
R1427 VDD.n1060 VDD.n1059 185
R1428 VDD.n1185 VDD.n1184 185
R1429 VDD.n1187 VDD.n1058 185
R1430 VDD.n1190 VDD.n1189 185
R1431 VDD.n1056 VDD.n1055 185
R1432 VDD.n1196 VDD.n1195 185
R1433 VDD.n1198 VDD.n1054 185
R1434 VDD.n1201 VDD.n1200 185
R1435 VDD.n1203 VDD.n1050 185
R1436 VDD.n1337 VDD.n1336 185
R1437 VDD.n1341 VDD.n967 185
R1438 VDD.n966 VDD.n963 185
R1439 VDD.n1345 VDD.n962 185
R1440 VDD.n1346 VDD.n961 185
R1441 VDD.n1347 VDD.n959 185
R1442 VDD.n958 VDD.n952 185
R1443 VDD.n956 VDD.n955 185
R1444 VDD.n954 VDD.n790 185
R1445 VDD.n1351 VDD.n787 185
R1446 VDD.n1353 VDD.n1352 185
R1447 VDD.n1355 VDD.n785 185
R1448 VDD.n1357 VDD.n1356 185
R1449 VDD.n1358 VDD.n780 185
R1450 VDD.n1360 VDD.n1359 185
R1451 VDD.n1362 VDD.n778 185
R1452 VDD.n1364 VDD.n1363 185
R1453 VDD.n1365 VDD.n771 185
R1454 VDD.n1367 VDD.n1366 185
R1455 VDD.n1369 VDD.n769 185
R1456 VDD.n1371 VDD.n1370 185
R1457 VDD.n1372 VDD.n764 185
R1458 VDD.n1374 VDD.n1373 185
R1459 VDD.n1376 VDD.n762 185
R1460 VDD.n1378 VDD.n1377 185
R1461 VDD.n1379 VDD.n758 185
R1462 VDD.n1381 VDD.n1380 185
R1463 VDD.n1383 VDD.n755 185
R1464 VDD.n1385 VDD.n1384 185
R1465 VDD.n756 VDD.n749 185
R1466 VDD.n1389 VDD.n753 185
R1467 VDD.n1390 VDD.n747 185
R1468 VDD.n1392 VDD.n1391 185
R1469 VDD.n1394 VDD.n746 185
R1470 VDD.n1396 VDD.n1395 185
R1471 VDD.n1398 VDD.n742 185
R1472 VDD.n1400 VDD.n1399 185
R1473 VDD.n1317 VDD.n743 185
R1474 VDD.n1322 VDD.n1321 185
R1475 VDD.n1324 VDD.n1316 185
R1476 VDD.n1325 VDD.n1315 185
R1477 VDD.n1328 VDD.n1327 185
R1478 VDD.n1329 VDD.n973 185
R1479 VDD.n973 VDD.n745 185
R1480 VDD.n1335 VDD.n970 185
R1481 VDD.n1335 VDD.n1334 185
R1482 VDD.n981 VDD.n969 185
R1483 VDD.n971 VDD.n969 185
R1484 VDD.n1308 VDD.n1307 185
R1485 VDD.n1309 VDD.n1308 185
R1486 VDD.n980 VDD.n979 185
R1487 VDD.n979 VDD.n978 185
R1488 VDD.n1301 VDD.n1300 185
R1489 VDD.n1300 VDD.n1299 185
R1490 VDD.n984 VDD.n983 185
R1491 VDD.n985 VDD.n984 185
R1492 VDD.n1290 VDD.n1289 185
R1493 VDD.n1291 VDD.n1290 185
R1494 VDD.n993 VDD.n992 185
R1495 VDD.n992 VDD.n991 185
R1496 VDD.n1285 VDD.n1284 185
R1497 VDD.n1284 VDD.n1283 185
R1498 VDD.n996 VDD.n995 185
R1499 VDD.n997 VDD.n996 185
R1500 VDD.n1274 VDD.n1273 185
R1501 VDD.n1275 VDD.n1274 185
R1502 VDD.n1005 VDD.n1004 185
R1503 VDD.n1004 VDD.n1003 185
R1504 VDD.n1269 VDD.n1268 185
R1505 VDD.n1268 VDD.n1267 185
R1506 VDD.n1008 VDD.n1007 185
R1507 VDD.t72 VDD.n1008 185
R1508 VDD.n1255 VDD.n1254 185
R1509 VDD.n1256 VDD.n1255 185
R1510 VDD.n1016 VDD.n1015 185
R1511 VDD.n1015 VDD.n1014 185
R1512 VDD.n1250 VDD.n1249 185
R1513 VDD.n1249 VDD.n1248 185
R1514 VDD.n1019 VDD.n1018 185
R1515 VDD.n1020 VDD.n1019 185
R1516 VDD.n1239 VDD.n1238 185
R1517 VDD.n1240 VDD.n1239 185
R1518 VDD.n1028 VDD.n1027 185
R1519 VDD.n1027 VDD.n1026 185
R1520 VDD.n1234 VDD.n1233 185
R1521 VDD.n1233 VDD.n1232 185
R1522 VDD.n1031 VDD.n1030 185
R1523 VDD.n1032 VDD.n1031 185
R1524 VDD.n1223 VDD.n1222 185
R1525 VDD.n1224 VDD.n1223 185
R1526 VDD.n1039 VDD.n1038 185
R1527 VDD.n1044 VDD.n1038 185
R1528 VDD.n1218 VDD.n1217 185
R1529 VDD.n1217 VDD.n1216 185
R1530 VDD.n1042 VDD.n1041 185
R1531 VDD.n1043 VDD.n1042 185
R1532 VDD.n1207 VDD.n1206 185
R1533 VDD.n1208 VDD.n1207 185
R1534 VDD.n2679 VDD.n2678 185
R1535 VDD.n2677 VDD.n88 185
R1536 VDD.n2676 VDD.n87 185
R1537 VDD.n2681 VDD.n87 185
R1538 VDD.n2675 VDD.n2674 185
R1539 VDD.n2673 VDD.n2672 185
R1540 VDD.n2671 VDD.n2670 185
R1541 VDD.n2669 VDD.n2668 185
R1542 VDD.n2667 VDD.n2666 185
R1543 VDD.n2665 VDD.n2664 185
R1544 VDD.n2663 VDD.n2662 185
R1545 VDD.n2661 VDD.n2660 185
R1546 VDD.n2659 VDD.n2658 185
R1547 VDD.n2657 VDD.n101 185
R1548 VDD.n100 VDD.n99 185
R1549 VDD.n2651 VDD.n2650 185
R1550 VDD.n2649 VDD.n2648 185
R1551 VDD.n2647 VDD.n2646 185
R1552 VDD.n2645 VDD.n2644 185
R1553 VDD.n2643 VDD.n2642 185
R1554 VDD.n2641 VDD.n2640 185
R1555 VDD.n2639 VDD.n2638 185
R1556 VDD.n2637 VDD.n2636 185
R1557 VDD.n2635 VDD.n2634 185
R1558 VDD.n2633 VDD.n2632 185
R1559 VDD.n2631 VDD.n2630 185
R1560 VDD.n2629 VDD.n2628 185
R1561 VDD.n2627 VDD.n2626 185
R1562 VDD.n2625 VDD.n2624 185
R1563 VDD.n2618 VDD.n114 185
R1564 VDD.n2620 VDD.n2619 185
R1565 VDD.n2617 VDD.n2616 185
R1566 VDD.n2615 VDD.n2614 185
R1567 VDD.n2613 VDD.n2612 185
R1568 VDD.n2611 VDD.n2610 185
R1569 VDD.n2590 VDD.n120 185
R1570 VDD.n2592 VDD.n2591 185
R1571 VDD.n2606 VDD.n2593 185
R1572 VDD.n2605 VDD.n2604 185
R1573 VDD.n2603 VDD.n2602 185
R1574 VDD.n2601 VDD.n2600 185
R1575 VDD.n2599 VDD.n2598 185
R1576 VDD.n2597 VDD.n67 185
R1577 VDD.n2684 VDD.n2683 185
R1578 VDD.n2861 VDD.n2860 185
R1579 VDD.n2866 VDD.n2865 185
R1580 VDD.n2868 VDD.n2867 185
R1581 VDD.n2870 VDD.n2869 185
R1582 VDD.n2872 VDD.n2871 185
R1583 VDD.n2874 VDD.n2873 185
R1584 VDD.n2876 VDD.n2875 185
R1585 VDD.n2878 VDD.n2877 185
R1586 VDD.n2880 VDD.n2879 185
R1587 VDD.n2882 VDD.n2881 185
R1588 VDD.n2884 VDD.n2883 185
R1589 VDD.n2886 VDD.n2885 185
R1590 VDD.n2888 VDD.n2887 185
R1591 VDD.n2891 VDD.n2890 185
R1592 VDD.n2889 VDD.n2821 185
R1593 VDD.n2896 VDD.n2895 185
R1594 VDD.n2898 VDD.n2897 185
R1595 VDD.n2900 VDD.n2899 185
R1596 VDD.n2902 VDD.n2901 185
R1597 VDD.n2904 VDD.n2903 185
R1598 VDD.n2906 VDD.n2905 185
R1599 VDD.n2908 VDD.n2907 185
R1600 VDD.n2910 VDD.n2909 185
R1601 VDD.n2912 VDD.n2911 185
R1602 VDD.n2914 VDD.n2913 185
R1603 VDD.n2916 VDD.n2915 185
R1604 VDD.n2918 VDD.n2917 185
R1605 VDD.n2920 VDD.n2919 185
R1606 VDD.n2922 VDD.n2921 185
R1607 VDD.n2807 VDD.n2804 185
R1608 VDD.n2926 VDD.n2808 185
R1609 VDD.n2928 VDD.n2927 185
R1610 VDD.n2930 VDD.n2929 185
R1611 VDD.n2932 VDD.n2931 185
R1612 VDD.n2934 VDD.n2933 185
R1613 VDD.n2936 VDD.n2935 185
R1614 VDD.n2938 VDD.n2937 185
R1615 VDD.n2940 VDD.n2939 185
R1616 VDD.n2942 VDD.n2941 185
R1617 VDD.n2945 VDD.n2944 185
R1618 VDD.n2943 VDD.n2795 185
R1619 VDD.n2949 VDD.n2792 185
R1620 VDD.n2951 VDD.n2950 185
R1621 VDD.n2952 VDD.n2951 185
R1622 VDD.n2857 VDD.n2770 185
R1623 VDD.n2953 VDD.n2770 185
R1624 VDD.n2856 VDD.n2769 185
R1625 VDD.n2954 VDD.n2769 185
R1626 VDD.n2855 VDD.n2854 185
R1627 VDD.n2854 VDD.n2761 185
R1628 VDD.n2837 VDD.n2760 185
R1629 VDD.n2960 VDD.n2760 185
R1630 VDD.n2850 VDD.n2759 185
R1631 VDD.n2961 VDD.n2759 185
R1632 VDD.n2849 VDD.n2758 185
R1633 VDD.n2962 VDD.n2758 185
R1634 VDD.n2848 VDD.n2847 185
R1635 VDD.n2847 VDD.n2750 185
R1636 VDD.n2839 VDD.n2749 185
R1637 VDD.n2968 VDD.n2749 185
R1638 VDD.n2843 VDD.n2748 185
R1639 VDD.n2969 VDD.n2748 185
R1640 VDD.n2842 VDD.n2747 185
R1641 VDD.n2970 VDD.n2747 185
R1642 VDD.n2739 VDD.n2738 185
R1643 VDD.n2740 VDD.n2739 185
R1644 VDD.n2978 VDD.n2977 185
R1645 VDD.n2977 VDD.n2976 185
R1646 VDD.n2979 VDD.n25 185
R1647 VDD.n25 VDD.n23 185
R1648 VDD.n2981 VDD.n2980 185
R1649 VDD.t0 VDD.n2981 185
R1650 VDD.n26 VDD.n24 185
R1651 VDD.n24 VDD.n22 185
R1652 VDD.n2732 VDD.n2731 185
R1653 VDD.n2731 VDD.n2730 185
R1654 VDD.n29 VDD.n28 185
R1655 VDD.n30 VDD.n29 185
R1656 VDD.n2721 VDD.n2720 185
R1657 VDD.n2722 VDD.n2721 185
R1658 VDD.n38 VDD.n37 185
R1659 VDD.n37 VDD.n36 185
R1660 VDD.n2716 VDD.n2715 185
R1661 VDD.n2715 VDD.n2714 185
R1662 VDD.n41 VDD.n40 185
R1663 VDD.n42 VDD.n41 185
R1664 VDD.n2705 VDD.n2704 185
R1665 VDD.n2706 VDD.n2705 185
R1666 VDD.n50 VDD.n49 185
R1667 VDD.n49 VDD.n48 185
R1668 VDD.n2700 VDD.n2699 185
R1669 VDD.n2699 VDD.n2698 185
R1670 VDD.n53 VDD.n52 185
R1671 VDD.n54 VDD.n53 185
R1672 VDD.n2689 VDD.n2688 185
R1673 VDD.n2690 VDD.n2689 185
R1674 VDD.n62 VDD.n61 185
R1675 VDD.n61 VDD.n60 185
R1676 VDD.n59 VDD.n58 185
R1677 VDD.n60 VDD.n59 185
R1678 VDD.n2692 VDD.n2691 185
R1679 VDD.n2691 VDD.n2690 185
R1680 VDD.n56 VDD.n55 185
R1681 VDD.n55 VDD.n54 185
R1682 VDD.n2697 VDD.n2696 185
R1683 VDD.n2698 VDD.n2697 185
R1684 VDD.n47 VDD.n46 185
R1685 VDD.n48 VDD.n47 185
R1686 VDD.n2708 VDD.n2707 185
R1687 VDD.n2707 VDD.n2706 185
R1688 VDD.n44 VDD.n43 185
R1689 VDD.n43 VDD.n42 185
R1690 VDD.n2713 VDD.n2712 185
R1691 VDD.n2714 VDD.n2713 185
R1692 VDD.n35 VDD.n34 185
R1693 VDD.n36 VDD.n35 185
R1694 VDD.n2724 VDD.n2723 185
R1695 VDD.n2723 VDD.n2722 185
R1696 VDD.n32 VDD.n31 185
R1697 VDD.n31 VDD.n30 185
R1698 VDD.n2729 VDD.n2728 185
R1699 VDD.n2730 VDD.n2729 185
R1700 VDD.n20 VDD.n18 185
R1701 VDD.n22 VDD.n20 185
R1702 VDD.n2983 VDD.n2982 185
R1703 VDD.n2982 VDD.t0 185
R1704 VDD.n21 VDD.n19 185
R1705 VDD.n23 VDD.n21 185
R1706 VDD.n2975 VDD.n2974 185
R1707 VDD.n2976 VDD.n2975 185
R1708 VDD.n2973 VDD.n2741 185
R1709 VDD.n2741 VDD.n2740 185
R1710 VDD.n2972 VDD.n2971 185
R1711 VDD.n2971 VDD.n2970 185
R1712 VDD.n2746 VDD.n2745 185
R1713 VDD.n2969 VDD.n2746 185
R1714 VDD.n2967 VDD.n2966 185
R1715 VDD.n2968 VDD.n2967 185
R1716 VDD.n2965 VDD.n2751 185
R1717 VDD.n2751 VDD.n2750 185
R1718 VDD.n2964 VDD.n2963 185
R1719 VDD.n2963 VDD.n2962 185
R1720 VDD.n2757 VDD.n2756 185
R1721 VDD.n2961 VDD.n2757 185
R1722 VDD.n2959 VDD.n2958 185
R1723 VDD.n2960 VDD.n2959 185
R1724 VDD.n2957 VDD.n2762 185
R1725 VDD.n2762 VDD.n2761 185
R1726 VDD.n2956 VDD.n2955 185
R1727 VDD.n2955 VDD.n2954 185
R1728 VDD.n2768 VDD.n2767 185
R1729 VDD.n2953 VDD.n2768 185
R1730 VDD.n1866 VDD.n1865 185
R1731 VDD.n1865 VDD.n424 185
R1732 VDD.n1867 VDD.n451 185
R1733 VDD.n1877 VDD.n451 185
R1734 VDD.n1868 VDD.n459 185
R1735 VDD.n459 VDD.n449 185
R1736 VDD.n1870 VDD.n1869 185
R1737 VDD.n1871 VDD.n1870 185
R1738 VDD.n460 VDD.n458 185
R1739 VDD.n458 VDD.n455 185
R1740 VDD.n1815 VDD.n467 185
R1741 VDD.n1825 VDD.n467 185
R1742 VDD.n1816 VDD.n474 185
R1743 VDD.n474 VDD.n465 185
R1744 VDD.n1818 VDD.n1817 185
R1745 VDD.n1819 VDD.n1818 185
R1746 VDD.n1814 VDD.n473 185
R1747 VDD.n480 VDD.n473 185
R1748 VDD.n1813 VDD.n1812 185
R1749 VDD.n1812 VDD.n1811 185
R1750 VDD.n476 VDD.n475 185
R1751 VDD.n477 VDD.n476 185
R1752 VDD.n1804 VDD.n1803 185
R1753 VDD.n1805 VDD.n1804 185
R1754 VDD.n1802 VDD.n487 185
R1755 VDD.n487 VDD.n484 185
R1756 VDD.n1801 VDD.n1800 185
R1757 VDD.n1800 VDD.n1799 185
R1758 VDD.n489 VDD.n488 185
R1759 VDD.n490 VDD.n489 185
R1760 VDD.n1792 VDD.n1791 185
R1761 VDD.n1793 VDD.n1792 185
R1762 VDD.n1790 VDD.n499 185
R1763 VDD.n499 VDD.n496 185
R1764 VDD.n1789 VDD.n1788 185
R1765 VDD.n1788 VDD.n1787 185
R1766 VDD.n501 VDD.n500 185
R1767 VDD.n502 VDD.n501 185
R1768 VDD.n1780 VDD.n1779 185
R1769 VDD.n1781 VDD.n1780 185
R1770 VDD.n1778 VDD.n511 185
R1771 VDD.n511 VDD.n508 185
R1772 VDD.n1777 VDD.n1776 185
R1773 VDD.n1776 VDD.n1775 185
R1774 VDD.n513 VDD.n512 185
R1775 VDD.n514 VDD.n513 185
R1776 VDD.n1768 VDD.n1767 185
R1777 VDD.n1769 VDD.n1768 185
R1778 VDD.n1766 VDD.n523 185
R1779 VDD.n523 VDD.n520 185
R1780 VDD.n1765 VDD.n1764 185
R1781 VDD.n1764 VDD.n1763 185
R1782 VDD.n525 VDD.n524 185
R1783 VDD.n526 VDD.n525 185
R1784 VDD.n1756 VDD.n1755 185
R1785 VDD.n1757 VDD.n1756 185
R1786 VDD.n1754 VDD.n535 185
R1787 VDD.n535 VDD.n532 185
R1788 VDD.n1753 VDD.n1752 185
R1789 VDD.n1752 VDD.n1751 185
R1790 VDD.n537 VDD.n536 185
R1791 VDD.n538 VDD.n537 185
R1792 VDD.n1744 VDD.n1743 185
R1793 VDD.n1745 VDD.n1744 185
R1794 VDD.n1742 VDD.n547 185
R1795 VDD.n547 VDD.n544 185
R1796 VDD.n1741 VDD.n1740 185
R1797 VDD.n1740 VDD.n1739 185
R1798 VDD.n549 VDD.n548 185
R1799 VDD.n550 VDD.n549 185
R1800 VDD.n1732 VDD.n1731 185
R1801 VDD.n1733 VDD.n1732 185
R1802 VDD.n1730 VDD.n559 185
R1803 VDD.n559 VDD.n556 185
R1804 VDD.n1729 VDD.n1728 185
R1805 VDD.n1728 VDD.n1727 185
R1806 VDD.n561 VDD.n560 185
R1807 VDD.n562 VDD.n561 185
R1808 VDD.n1720 VDD.n1719 185
R1809 VDD.n1721 VDD.n1720 185
R1810 VDD.n1718 VDD.n571 185
R1811 VDD.n571 VDD.n568 185
R1812 VDD.n1717 VDD.n1716 185
R1813 VDD.n1716 VDD.n1715 185
R1814 VDD.n573 VDD.n572 185
R1815 VDD.n574 VDD.n573 185
R1816 VDD.n1708 VDD.n1707 185
R1817 VDD.n1709 VDD.n1708 185
R1818 VDD.n1706 VDD.n583 185
R1819 VDD.n583 VDD.n580 185
R1820 VDD.n1705 VDD.n1704 185
R1821 VDD.n1704 VDD.n1703 185
R1822 VDD.n585 VDD.n584 185
R1823 VDD.n586 VDD.n585 185
R1824 VDD.n1696 VDD.n1695 185
R1825 VDD.n1697 VDD.n1696 185
R1826 VDD.n1694 VDD.n594 185
R1827 VDD.n600 VDD.n594 185
R1828 VDD.n1693 VDD.n1692 185
R1829 VDD.n1692 VDD.n1691 185
R1830 VDD.n596 VDD.n595 185
R1831 VDD.n597 VDD.n596 185
R1832 VDD.n1684 VDD.n1683 185
R1833 VDD.n1685 VDD.n1684 185
R1834 VDD.n1682 VDD.n606 185
R1835 VDD.n612 VDD.n606 185
R1836 VDD.n1681 VDD.n1680 185
R1837 VDD.n1680 VDD.n1679 185
R1838 VDD.n608 VDD.n607 185
R1839 VDD.n609 VDD.n608 185
R1840 VDD.n1672 VDD.n1671 185
R1841 VDD.n1673 VDD.n1672 185
R1842 VDD.n1670 VDD.n619 185
R1843 VDD.n619 VDD.n616 185
R1844 VDD.n1669 VDD.n1668 185
R1845 VDD.n1668 VDD.n1667 185
R1846 VDD.n621 VDD.n620 185
R1847 VDD.n622 VDD.n621 185
R1848 VDD.n1660 VDD.n1659 185
R1849 VDD.n1661 VDD.n1660 185
R1850 VDD.n1658 VDD.n631 185
R1851 VDD.n631 VDD.n628 185
R1852 VDD.n1657 VDD.n1656 185
R1853 VDD.n1656 VDD.n1655 185
R1854 VDD.n633 VDD.n632 185
R1855 VDD.n634 VDD.n633 185
R1856 VDD.n1648 VDD.n1647 185
R1857 VDD.n1649 VDD.n1648 185
R1858 VDD.n1646 VDD.n643 185
R1859 VDD.n643 VDD.n640 185
R1860 VDD.n1645 VDD.n1644 185
R1861 VDD.n1644 VDD.n1643 185
R1862 VDD.n645 VDD.n644 185
R1863 VDD.n654 VDD.n645 185
R1864 VDD.n1636 VDD.n1635 185
R1865 VDD.n1637 VDD.n1636 185
R1866 VDD.n1634 VDD.n655 185
R1867 VDD.n655 VDD.n651 185
R1868 VDD.n1633 VDD.n1632 185
R1869 VDD.n1632 VDD.n1631 185
R1870 VDD.n657 VDD.n656 185
R1871 VDD.n658 VDD.n657 185
R1872 VDD.n1624 VDD.n1623 185
R1873 VDD.n1625 VDD.n1624 185
R1874 VDD.n1622 VDD.n667 185
R1875 VDD.n667 VDD.n664 185
R1876 VDD.n1621 VDD.n1620 185
R1877 VDD.n1620 VDD.n1619 185
R1878 VDD.n669 VDD.n668 185
R1879 VDD.n670 VDD.n669 185
R1880 VDD.n1612 VDD.n1611 185
R1881 VDD.n1613 VDD.n1612 185
R1882 VDD.n1610 VDD.n679 185
R1883 VDD.n679 VDD.n676 185
R1884 VDD.n1609 VDD.n1608 185
R1885 VDD.n1608 VDD.n1607 185
R1886 VDD.n681 VDD.n680 185
R1887 VDD.n682 VDD.n681 185
R1888 VDD.n1600 VDD.n1599 185
R1889 VDD.n1601 VDD.n1600 185
R1890 VDD.n1598 VDD.n691 185
R1891 VDD.n691 VDD.n688 185
R1892 VDD.n1597 VDD.n1596 185
R1893 VDD.n1596 VDD.n1595 185
R1894 VDD.n693 VDD.n692 185
R1895 VDD.n694 VDD.n693 185
R1896 VDD.n1588 VDD.n1587 185
R1897 VDD.n1589 VDD.n1588 185
R1898 VDD.n1586 VDD.n703 185
R1899 VDD.n703 VDD.n700 185
R1900 VDD.n1585 VDD.n1584 185
R1901 VDD.n1584 VDD.n1583 185
R1902 VDD.n705 VDD.n704 185
R1903 VDD.n706 VDD.n705 185
R1904 VDD.n1576 VDD.n1575 185
R1905 VDD.n1577 VDD.n1576 185
R1906 VDD.n1574 VDD.n715 185
R1907 VDD.n715 VDD.n712 185
R1908 VDD.n1573 VDD.n1572 185
R1909 VDD.n1572 VDD.n1571 185
R1910 VDD.n717 VDD.n716 185
R1911 VDD.n718 VDD.n717 185
R1912 VDD.n1835 VDD.n432 185
R1913 VDD.n1909 VDD.n432 185
R1914 VDD.n1837 VDD.n1836 185
R1915 VDD.n1840 VDD.n1839 185
R1916 VDD.n1842 VDD.n1841 185
R1917 VDD.n1844 VDD.n1843 185
R1918 VDD.n1846 VDD.n1845 185
R1919 VDD.n1848 VDD.n1847 185
R1920 VDD.n1850 VDD.n1849 185
R1921 VDD.n1852 VDD.n1851 185
R1922 VDD.n1854 VDD.n1853 185
R1923 VDD.n1856 VDD.n1855 185
R1924 VDD.n1858 VDD.n1857 185
R1925 VDD.n1860 VDD.n1859 185
R1926 VDD.n1862 VDD.n1861 185
R1927 VDD.n1864 VDD.n1863 185
R1928 VDD.n1834 VDD.n1833 185
R1929 VDD.n1833 VDD.n424 185
R1930 VDD.n1832 VDD.n450 185
R1931 VDD.n1877 VDD.n450 185
R1932 VDD.n1831 VDD.n1830 185
R1933 VDD.n1830 VDD.n449 185
R1934 VDD.n1829 VDD.n457 185
R1935 VDD.n1871 VDD.n457 185
R1936 VDD.n1828 VDD.n1827 185
R1937 VDD.n1827 VDD.n455 185
R1938 VDD.n1826 VDD.n463 185
R1939 VDD.n1826 VDD.n1825 185
R1940 VDD.n808 VDD.n464 185
R1941 VDD.n465 VDD.n464 185
R1942 VDD.n809 VDD.n472 185
R1943 VDD.n1819 VDD.n472 185
R1944 VDD.n811 VDD.n810 185
R1945 VDD.n810 VDD.n480 185
R1946 VDD.n812 VDD.n479 185
R1947 VDD.n1811 VDD.n479 185
R1948 VDD.n814 VDD.n813 185
R1949 VDD.n813 VDD.n477 185
R1950 VDD.n815 VDD.n486 185
R1951 VDD.n1805 VDD.n486 185
R1952 VDD.n817 VDD.n816 185
R1953 VDD.n816 VDD.n484 185
R1954 VDD.n818 VDD.n492 185
R1955 VDD.n1799 VDD.n492 185
R1956 VDD.n820 VDD.n819 185
R1957 VDD.n819 VDD.n490 185
R1958 VDD.n821 VDD.n498 185
R1959 VDD.n1793 VDD.n498 185
R1960 VDD.n823 VDD.n822 185
R1961 VDD.n822 VDD.n496 185
R1962 VDD.n824 VDD.n504 185
R1963 VDD.n1787 VDD.n504 185
R1964 VDD.n826 VDD.n825 185
R1965 VDD.n825 VDD.n502 185
R1966 VDD.n827 VDD.n510 185
R1967 VDD.n1781 VDD.n510 185
R1968 VDD.n829 VDD.n828 185
R1969 VDD.n828 VDD.n508 185
R1970 VDD.n830 VDD.n516 185
R1971 VDD.n1775 VDD.n516 185
R1972 VDD.n832 VDD.n831 185
R1973 VDD.n831 VDD.n514 185
R1974 VDD.n833 VDD.n522 185
R1975 VDD.n1769 VDD.n522 185
R1976 VDD.n835 VDD.n834 185
R1977 VDD.n834 VDD.n520 185
R1978 VDD.n836 VDD.n528 185
R1979 VDD.n1763 VDD.n528 185
R1980 VDD.n838 VDD.n837 185
R1981 VDD.n837 VDD.n526 185
R1982 VDD.n839 VDD.n534 185
R1983 VDD.n1757 VDD.n534 185
R1984 VDD.n841 VDD.n840 185
R1985 VDD.n840 VDD.n532 185
R1986 VDD.n842 VDD.n540 185
R1987 VDD.n1751 VDD.n540 185
R1988 VDD.n844 VDD.n843 185
R1989 VDD.n843 VDD.n538 185
R1990 VDD.n845 VDD.n546 185
R1991 VDD.n1745 VDD.n546 185
R1992 VDD.n847 VDD.n846 185
R1993 VDD.n846 VDD.n544 185
R1994 VDD.n848 VDD.n552 185
R1995 VDD.n1739 VDD.n552 185
R1996 VDD.n850 VDD.n849 185
R1997 VDD.n849 VDD.n550 185
R1998 VDD.n851 VDD.n558 185
R1999 VDD.n1733 VDD.n558 185
R2000 VDD.n853 VDD.n852 185
R2001 VDD.n852 VDD.n556 185
R2002 VDD.n854 VDD.n564 185
R2003 VDD.n1727 VDD.n564 185
R2004 VDD.n856 VDD.n855 185
R2005 VDD.n855 VDD.n562 185
R2006 VDD.n857 VDD.n570 185
R2007 VDD.n1721 VDD.n570 185
R2008 VDD.n859 VDD.n858 185
R2009 VDD.n858 VDD.n568 185
R2010 VDD.n860 VDD.n576 185
R2011 VDD.n1715 VDD.n576 185
R2012 VDD.n862 VDD.n861 185
R2013 VDD.n861 VDD.n574 185
R2014 VDD.n863 VDD.n582 185
R2015 VDD.n1709 VDD.n582 185
R2016 VDD.n865 VDD.n864 185
R2017 VDD.n864 VDD.n580 185
R2018 VDD.n866 VDD.n588 185
R2019 VDD.n1703 VDD.n588 185
R2020 VDD.n868 VDD.n867 185
R2021 VDD.n867 VDD.n586 185
R2022 VDD.n869 VDD.n593 185
R2023 VDD.n1697 VDD.n593 185
R2024 VDD.n871 VDD.n870 185
R2025 VDD.n870 VDD.n600 185
R2026 VDD.n872 VDD.n599 185
R2027 VDD.n1691 VDD.n599 185
R2028 VDD.n874 VDD.n873 185
R2029 VDD.n873 VDD.n597 185
R2030 VDD.n875 VDD.n605 185
R2031 VDD.n1685 VDD.n605 185
R2032 VDD.n877 VDD.n876 185
R2033 VDD.n876 VDD.n612 185
R2034 VDD.n878 VDD.n611 185
R2035 VDD.n1679 VDD.n611 185
R2036 VDD.n880 VDD.n879 185
R2037 VDD.n879 VDD.n609 185
R2038 VDD.n881 VDD.n618 185
R2039 VDD.n1673 VDD.n618 185
R2040 VDD.n883 VDD.n882 185
R2041 VDD.n882 VDD.n616 185
R2042 VDD.n884 VDD.n624 185
R2043 VDD.n1667 VDD.n624 185
R2044 VDD.n886 VDD.n885 185
R2045 VDD.n885 VDD.n622 185
R2046 VDD.n887 VDD.n630 185
R2047 VDD.n1661 VDD.n630 185
R2048 VDD.n889 VDD.n888 185
R2049 VDD.n888 VDD.n628 185
R2050 VDD.n890 VDD.n636 185
R2051 VDD.n1655 VDD.n636 185
R2052 VDD.n892 VDD.n891 185
R2053 VDD.n891 VDD.n634 185
R2054 VDD.n893 VDD.n642 185
R2055 VDD.n1649 VDD.n642 185
R2056 VDD.n895 VDD.n894 185
R2057 VDD.n894 VDD.n640 185
R2058 VDD.n896 VDD.n647 185
R2059 VDD.n1643 VDD.n647 185
R2060 VDD.n898 VDD.n897 185
R2061 VDD.n897 VDD.n654 185
R2062 VDD.n899 VDD.n653 185
R2063 VDD.n1637 VDD.n653 185
R2064 VDD.n901 VDD.n900 185
R2065 VDD.n900 VDD.n651 185
R2066 VDD.n902 VDD.n660 185
R2067 VDD.n1631 VDD.n660 185
R2068 VDD.n904 VDD.n903 185
R2069 VDD.n903 VDD.n658 185
R2070 VDD.n905 VDD.n666 185
R2071 VDD.n1625 VDD.n666 185
R2072 VDD.n907 VDD.n906 185
R2073 VDD.n906 VDD.n664 185
R2074 VDD.n908 VDD.n672 185
R2075 VDD.n1619 VDD.n672 185
R2076 VDD.n910 VDD.n909 185
R2077 VDD.n909 VDD.n670 185
R2078 VDD.n911 VDD.n678 185
R2079 VDD.n1613 VDD.n678 185
R2080 VDD.n913 VDD.n912 185
R2081 VDD.n912 VDD.n676 185
R2082 VDD.n914 VDD.n684 185
R2083 VDD.n1607 VDD.n684 185
R2084 VDD.n916 VDD.n915 185
R2085 VDD.n915 VDD.n682 185
R2086 VDD.n917 VDD.n690 185
R2087 VDD.n1601 VDD.n690 185
R2088 VDD.n919 VDD.n918 185
R2089 VDD.n918 VDD.n688 185
R2090 VDD.n920 VDD.n696 185
R2091 VDD.n1595 VDD.n696 185
R2092 VDD.n922 VDD.n921 185
R2093 VDD.n921 VDD.n694 185
R2094 VDD.n923 VDD.n702 185
R2095 VDD.n1589 VDD.n702 185
R2096 VDD.n925 VDD.n924 185
R2097 VDD.n924 VDD.n700 185
R2098 VDD.n926 VDD.n708 185
R2099 VDD.n1583 VDD.n708 185
R2100 VDD.n928 VDD.n927 185
R2101 VDD.n927 VDD.n706 185
R2102 VDD.n929 VDD.n714 185
R2103 VDD.n1577 VDD.n714 185
R2104 VDD.n931 VDD.n930 185
R2105 VDD.n930 VDD.n712 185
R2106 VDD.n932 VDD.n720 185
R2107 VDD.n1571 VDD.n720 185
R2108 VDD.n934 VDD.n933 185
R2109 VDD.n933 VDD.n718 185
R2110 VDD.n792 VDD.n791 185
R2111 VDD.n794 VDD.n793 185
R2112 VDD.n796 VDD.n795 185
R2113 VDD.n798 VDD.n797 185
R2114 VDD.n800 VDD.n799 185
R2115 VDD.n802 VDD.n801 185
R2116 VDD.n804 VDD.n803 185
R2117 VDD.n949 VDD.n805 185
R2118 VDD.n948 VDD.n947 185
R2119 VDD.n946 VDD.n945 185
R2120 VDD.n944 VDD.n943 185
R2121 VDD.n942 VDD.n941 185
R2122 VDD.n940 VDD.n939 185
R2123 VDD.n937 VDD.n936 185
R2124 VDD.n935 VDD.n737 185
R2125 VDD.n1564 VDD.n737 185
R2126 VDD.t98 VDD.t102 180.078
R2127 VDD.t78 VDD.t114 180.078
R2128 VDD.n2691 VDD.n59 146.341
R2129 VDD.n2691 VDD.n55 146.341
R2130 VDD.n2697 VDD.n55 146.341
R2131 VDD.n2697 VDD.n47 146.341
R2132 VDD.n2707 VDD.n47 146.341
R2133 VDD.n2707 VDD.n43 146.341
R2134 VDD.n2713 VDD.n43 146.341
R2135 VDD.n2713 VDD.n35 146.341
R2136 VDD.n2723 VDD.n35 146.341
R2137 VDD.n2723 VDD.n31 146.341
R2138 VDD.n2729 VDD.n31 146.341
R2139 VDD.n2729 VDD.n20 146.341
R2140 VDD.n2982 VDD.n20 146.341
R2141 VDD.n2982 VDD.n21 146.341
R2142 VDD.n2975 VDD.n21 146.341
R2143 VDD.n2975 VDD.n2741 146.341
R2144 VDD.n2971 VDD.n2741 146.341
R2145 VDD.n2971 VDD.n2746 146.341
R2146 VDD.n2967 VDD.n2746 146.341
R2147 VDD.n2967 VDD.n2751 146.341
R2148 VDD.n2963 VDD.n2751 146.341
R2149 VDD.n2963 VDD.n2757 146.341
R2150 VDD.n2959 VDD.n2757 146.341
R2151 VDD.n2959 VDD.n2762 146.341
R2152 VDD.n2955 VDD.n2762 146.341
R2153 VDD.n2955 VDD.n2768 146.341
R2154 VDD.n2951 VDD.n2792 146.341
R2155 VDD.n2944 VDD.n2943 146.341
R2156 VDD.n2941 VDD.n2940 146.341
R2157 VDD.n2937 VDD.n2936 146.341
R2158 VDD.n2933 VDD.n2932 146.341
R2159 VDD.n2929 VDD.n2928 146.341
R2160 VDD.n2808 VDD.n2807 146.341
R2161 VDD.n2921 VDD.n2920 146.341
R2162 VDD.n2917 VDD.n2916 146.341
R2163 VDD.n2913 VDD.n2912 146.341
R2164 VDD.n2909 VDD.n2908 146.341
R2165 VDD.n2905 VDD.n2904 146.341
R2166 VDD.n2901 VDD.n2900 146.341
R2167 VDD.n2897 VDD.n2896 146.341
R2168 VDD.n2890 VDD.n2889 146.341
R2169 VDD.n2887 VDD.n2886 146.341
R2170 VDD.n2883 VDD.n2882 146.341
R2171 VDD.n2879 VDD.n2878 146.341
R2172 VDD.n2875 VDD.n2874 146.341
R2173 VDD.n2871 VDD.n2870 146.341
R2174 VDD.n2867 VDD.n2866 146.341
R2175 VDD.n2689 VDD.n61 146.341
R2176 VDD.n2689 VDD.n53 146.341
R2177 VDD.n2699 VDD.n53 146.341
R2178 VDD.n2699 VDD.n49 146.341
R2179 VDD.n2705 VDD.n49 146.341
R2180 VDD.n2705 VDD.n41 146.341
R2181 VDD.n2715 VDD.n41 146.341
R2182 VDD.n2715 VDD.n37 146.341
R2183 VDD.n2721 VDD.n37 146.341
R2184 VDD.n2721 VDD.n29 146.341
R2185 VDD.n2731 VDD.n29 146.341
R2186 VDD.n2731 VDD.n24 146.341
R2187 VDD.n2981 VDD.n24 146.341
R2188 VDD.n2981 VDD.n25 146.341
R2189 VDD.n2977 VDD.n25 146.341
R2190 VDD.n2977 VDD.n2739 146.341
R2191 VDD.n2747 VDD.n2739 146.341
R2192 VDD.n2748 VDD.n2747 146.341
R2193 VDD.n2749 VDD.n2748 146.341
R2194 VDD.n2847 VDD.n2749 146.341
R2195 VDD.n2847 VDD.n2758 146.341
R2196 VDD.n2759 VDD.n2758 146.341
R2197 VDD.n2760 VDD.n2759 146.341
R2198 VDD.n2854 VDD.n2760 146.341
R2199 VDD.n2854 VDD.n2769 146.341
R2200 VDD.n2770 VDD.n2769 146.341
R2201 VDD.n88 VDD.n87 146.341
R2202 VDD.n2674 VDD.n87 146.341
R2203 VDD.n2672 VDD.n2671 146.341
R2204 VDD.n2668 VDD.n2667 146.341
R2205 VDD.n2664 VDD.n2663 146.341
R2206 VDD.n2660 VDD.n2659 146.341
R2207 VDD.n101 VDD.n100 146.341
R2208 VDD.n2650 VDD.n2649 146.341
R2209 VDD.n2646 VDD.n2645 146.341
R2210 VDD.n2642 VDD.n2641 146.341
R2211 VDD.n2638 VDD.n2637 146.341
R2212 VDD.n2634 VDD.n2633 146.341
R2213 VDD.n2630 VDD.n2629 146.341
R2214 VDD.n2626 VDD.n2625 146.341
R2215 VDD.n2619 VDD.n2618 146.341
R2216 VDD.n2616 VDD.n2615 146.341
R2217 VDD.n2612 VDD.n2611 146.341
R2218 VDD.n2591 VDD.n2590 146.341
R2219 VDD.n2604 VDD.n2593 146.341
R2220 VDD.n2602 VDD.n2601 146.341
R2221 VDD.n2598 VDD.n67 146.341
R2222 VDD.n1327 VDD.n973 146.341
R2223 VDD.n1325 VDD.n1324 146.341
R2224 VDD.n1322 VDD.n1317 146.341
R2225 VDD.n1399 VDD.n1398 146.341
R2226 VDD.n1396 VDD.n1394 146.341
R2227 VDD.n1392 VDD.n747 146.341
R2228 VDD.n756 VDD.n753 146.341
R2229 VDD.n1384 VDD.n1383 146.341
R2230 VDD.n1381 VDD.n758 146.341
R2231 VDD.n1377 VDD.n1376 146.341
R2232 VDD.n1374 VDD.n764 146.341
R2233 VDD.n1370 VDD.n1369 146.341
R2234 VDD.n1367 VDD.n771 146.341
R2235 VDD.n1363 VDD.n1362 146.341
R2236 VDD.n1360 VDD.n780 146.341
R2237 VDD.n1356 VDD.n1355 146.341
R2238 VDD.n1353 VDD.n787 146.341
R2239 VDD.n956 VDD.n954 146.341
R2240 VDD.n959 VDD.n958 146.341
R2241 VDD.n962 VDD.n961 146.341
R2242 VDD.n967 VDD.n966 146.341
R2243 VDD.n1207 VDD.n1042 146.341
R2244 VDD.n1217 VDD.n1042 146.341
R2245 VDD.n1217 VDD.n1038 146.341
R2246 VDD.n1223 VDD.n1038 146.341
R2247 VDD.n1223 VDD.n1031 146.341
R2248 VDD.n1233 VDD.n1031 146.341
R2249 VDD.n1233 VDD.n1027 146.341
R2250 VDD.n1239 VDD.n1027 146.341
R2251 VDD.n1239 VDD.n1019 146.341
R2252 VDD.n1249 VDD.n1019 146.341
R2253 VDD.n1249 VDD.n1015 146.341
R2254 VDD.n1255 VDD.n1015 146.341
R2255 VDD.n1255 VDD.n1008 146.341
R2256 VDD.n1268 VDD.n1008 146.341
R2257 VDD.n1268 VDD.n1004 146.341
R2258 VDD.n1274 VDD.n1004 146.341
R2259 VDD.n1274 VDD.n996 146.341
R2260 VDD.n1284 VDD.n996 146.341
R2261 VDD.n1284 VDD.n992 146.341
R2262 VDD.n1290 VDD.n992 146.341
R2263 VDD.n1290 VDD.n984 146.341
R2264 VDD.n1300 VDD.n984 146.341
R2265 VDD.n1300 VDD.n979 146.341
R2266 VDD.n1308 VDD.n979 146.341
R2267 VDD.n1308 VDD.n969 146.341
R2268 VDD.n1335 VDD.n969 146.341
R2269 VDD.n1104 VDD.n1103 146.341
R2270 VDD.n1106 VDD.n1104 146.341
R2271 VDD.n1112 VDD.n1095 146.341
R2272 VDD.n1116 VDD.n1114 146.341
R2273 VDD.n1122 VDD.n1091 146.341
R2274 VDD.n1126 VDD.n1124 146.341
R2275 VDD.n1132 VDD.n1085 146.341
R2276 VDD.n1136 VDD.n1134 146.341
R2277 VDD.n1142 VDD.n1081 146.341
R2278 VDD.n1146 VDD.n1144 146.341
R2279 VDD.n1153 VDD.n1077 146.341
R2280 VDD.n1156 VDD.n1155 146.341
R2281 VDD.n1158 VDD.n1075 146.341
R2282 VDD.n1165 VDD.n1067 146.341
R2283 VDD.n1169 VDD.n1167 146.341
R2284 VDD.n1175 VDD.n1063 146.341
R2285 VDD.n1179 VDD.n1177 146.341
R2286 VDD.n1185 VDD.n1059 146.341
R2287 VDD.n1189 VDD.n1187 146.341
R2288 VDD.n1196 VDD.n1055 146.341
R2289 VDD.n1200 VDD.n1198 146.341
R2290 VDD.n1209 VDD.n1045 146.341
R2291 VDD.n1215 VDD.n1045 146.341
R2292 VDD.n1215 VDD.n1037 146.341
R2293 VDD.n1225 VDD.n1037 146.341
R2294 VDD.n1225 VDD.n1033 146.341
R2295 VDD.n1231 VDD.n1033 146.341
R2296 VDD.n1231 VDD.n1025 146.341
R2297 VDD.n1241 VDD.n1025 146.341
R2298 VDD.n1241 VDD.n1021 146.341
R2299 VDD.n1247 VDD.n1021 146.341
R2300 VDD.n1247 VDD.n1013 146.341
R2301 VDD.n1257 VDD.n1013 146.341
R2302 VDD.n1257 VDD.n1009 146.341
R2303 VDD.n1266 VDD.n1009 146.341
R2304 VDD.n1266 VDD.n1002 146.341
R2305 VDD.n1276 VDD.n1002 146.341
R2306 VDD.n1276 VDD.n998 146.341
R2307 VDD.n1282 VDD.n998 146.341
R2308 VDD.n1282 VDD.n990 146.341
R2309 VDD.n1292 VDD.n990 146.341
R2310 VDD.n1292 VDD.n986 146.341
R2311 VDD.n1298 VDD.n986 146.341
R2312 VDD.n1298 VDD.n977 146.341
R2313 VDD.n1310 VDD.n977 146.341
R2314 VDD.n1310 VDD.n972 146.341
R2315 VDD.n1333 VDD.n972 146.341
R2316 VDD.n9 VDD.n7 142.626
R2317 VDD.n2 VDD.n0 142.626
R2318 VDD.n807 VDD.t21 141.964
R2319 VDD.n462 VDD.t57 141.964
R2320 VDD.n1404 VDD.t36 141.964
R2321 VDD.n444 VDD.t51 141.964
R2322 VDD.n1925 VDD.t63 141.964
R2323 VDD.n152 VDD.t6 141.964
R2324 VDD.n2086 VDD.t60 141.964
R2325 VDD.n129 VDD.t54 141.964
R2326 VDD.n2247 VDD.n1909 141.798
R2327 VDD.n9 VDD.n8 138.653
R2328 VDD.n11 VDD.n10 138.653
R2329 VDD.n13 VDD.n12 138.653
R2330 VDD.n6 VDD.n5 138.653
R2331 VDD.n4 VDD.n3 138.653
R2332 VDD.n2 VDD.n1 138.653
R2333 VDD.n1053 VDD.t66 120.618
R2334 VDD.n1070 VDD.t69 120.618
R2335 VDD.n1087 VDD.t46 120.618
R2336 VDD.n1339 VDD.t40 120.618
R2337 VDD.n777 VDD.t43 120.618
R2338 VDD.n751 VDD.t18 120.618
R2339 VDD.n2863 VDD.t31 120.618
R2340 VDD.n2823 VDD.t34 120.618
R2341 VDD.n2806 VDD.t14 120.618
R2342 VDD.n116 VDD.t24 120.618
R2343 VDD.n2656 VDD.t9 120.618
R2344 VDD.n65 VDD.t27 120.618
R2345 VDD.n1260 VDD.t76 102.752
R2346 VDD.n2985 VDD.t2 101.252
R2347 VDD.n1261 VDD.t73 99.6472
R2348 VDD.n1260 VDD.t77 99.6472
R2349 VDD.n2566 VDD.n2565 99.5127
R2350 VDD.n2563 VDD.n144 99.5127
R2351 VDD.n2559 VDD.n2558 99.5127
R2352 VDD.n2556 VDD.n147 99.5127
R2353 VDD.n2551 VDD.n2550 99.5127
R2354 VDD.n2548 VDD.n150 99.5127
R2355 VDD.n2544 VDD.n2543 99.5127
R2356 VDD.n2217 VDD.n419 99.5127
R2357 VDD.n2213 VDD.n419 99.5127
R2358 VDD.n2213 VDD.n413 99.5127
R2359 VDD.n2210 VDD.n413 99.5127
R2360 VDD.n2210 VDD.n407 99.5127
R2361 VDD.n2207 VDD.n407 99.5127
R2362 VDD.n2207 VDD.n401 99.5127
R2363 VDD.n2204 VDD.n401 99.5127
R2364 VDD.n2204 VDD.n395 99.5127
R2365 VDD.n2201 VDD.n395 99.5127
R2366 VDD.n2201 VDD.n389 99.5127
R2367 VDD.n2198 VDD.n389 99.5127
R2368 VDD.n2198 VDD.n383 99.5127
R2369 VDD.n2195 VDD.n383 99.5127
R2370 VDD.n2195 VDD.n377 99.5127
R2371 VDD.n2192 VDD.n377 99.5127
R2372 VDD.n2192 VDD.n371 99.5127
R2373 VDD.n2189 VDD.n371 99.5127
R2374 VDD.n2189 VDD.n364 99.5127
R2375 VDD.n2186 VDD.n364 99.5127
R2376 VDD.n2186 VDD.n358 99.5127
R2377 VDD.n2183 VDD.n358 99.5127
R2378 VDD.n2183 VDD.n352 99.5127
R2379 VDD.n2180 VDD.n352 99.5127
R2380 VDD.n2180 VDD.n346 99.5127
R2381 VDD.n2177 VDD.n346 99.5127
R2382 VDD.n2177 VDD.n341 99.5127
R2383 VDD.n2174 VDD.n341 99.5127
R2384 VDD.n2174 VDD.n335 99.5127
R2385 VDD.n2171 VDD.n335 99.5127
R2386 VDD.n2171 VDD.n329 99.5127
R2387 VDD.n2168 VDD.n329 99.5127
R2388 VDD.n2168 VDD.n322 99.5127
R2389 VDD.n2165 VDD.n322 99.5127
R2390 VDD.n2165 VDD.n316 99.5127
R2391 VDD.n2162 VDD.n316 99.5127
R2392 VDD.n2162 VDD.n310 99.5127
R2393 VDD.n2159 VDD.n310 99.5127
R2394 VDD.n2159 VDD.n304 99.5127
R2395 VDD.n2156 VDD.n304 99.5127
R2396 VDD.n2156 VDD.n299 99.5127
R2397 VDD.n2153 VDD.n299 99.5127
R2398 VDD.n2153 VDD.n293 99.5127
R2399 VDD.n2150 VDD.n293 99.5127
R2400 VDD.n2150 VDD.n287 99.5127
R2401 VDD.n2147 VDD.n287 99.5127
R2402 VDD.n2147 VDD.n281 99.5127
R2403 VDD.n2144 VDD.n281 99.5127
R2404 VDD.n2144 VDD.n275 99.5127
R2405 VDD.n2141 VDD.n275 99.5127
R2406 VDD.n2141 VDD.n269 99.5127
R2407 VDD.n2138 VDD.n269 99.5127
R2408 VDD.n2138 VDD.n263 99.5127
R2409 VDD.n2135 VDD.n263 99.5127
R2410 VDD.n2135 VDD.n257 99.5127
R2411 VDD.n2132 VDD.n257 99.5127
R2412 VDD.n2132 VDD.n251 99.5127
R2413 VDD.n2129 VDD.n251 99.5127
R2414 VDD.n2129 VDD.n245 99.5127
R2415 VDD.n2126 VDD.n245 99.5127
R2416 VDD.n2126 VDD.n239 99.5127
R2417 VDD.n2123 VDD.n239 99.5127
R2418 VDD.n2123 VDD.n233 99.5127
R2419 VDD.n2120 VDD.n233 99.5127
R2420 VDD.n2120 VDD.n227 99.5127
R2421 VDD.n2117 VDD.n227 99.5127
R2422 VDD.n2117 VDD.n220 99.5127
R2423 VDD.n2114 VDD.n220 99.5127
R2424 VDD.n2114 VDD.n214 99.5127
R2425 VDD.n2111 VDD.n214 99.5127
R2426 VDD.n2111 VDD.n209 99.5127
R2427 VDD.n2108 VDD.n209 99.5127
R2428 VDD.n2108 VDD.n203 99.5127
R2429 VDD.n2105 VDD.n203 99.5127
R2430 VDD.n2105 VDD.n197 99.5127
R2431 VDD.n2102 VDD.n197 99.5127
R2432 VDD.n2102 VDD.n191 99.5127
R2433 VDD.n2099 VDD.n191 99.5127
R2434 VDD.n2099 VDD.n185 99.5127
R2435 VDD.n2096 VDD.n185 99.5127
R2436 VDD.n2096 VDD.n178 99.5127
R2437 VDD.n2093 VDD.n178 99.5127
R2438 VDD.n2093 VDD.n172 99.5127
R2439 VDD.n2090 VDD.n172 99.5127
R2440 VDD.n2090 VDD.n166 99.5127
R2441 VDD.n166 VDD.n158 99.5127
R2442 VDD.n2535 VDD.n158 99.5127
R2443 VDD.n2536 VDD.n2535 99.5127
R2444 VDD.n2536 VDD.n137 99.5127
R2445 VDD.n156 VDD.n137 99.5127
R2446 VDD.n2084 VDD.n2083 99.5127
R2447 VDD.n2240 VDD.n2083 99.5127
R2448 VDD.n2238 VDD.n2237 99.5127
R2449 VDD.n2234 VDD.n2233 99.5127
R2450 VDD.n2230 VDD.n2229 99.5127
R2451 VDD.n2226 VDD.n2225 99.5127
R2452 VDD.n2222 VDD.n2221 99.5127
R2453 VDD.n2255 VDD.n417 99.5127
R2454 VDD.n2255 VDD.n415 99.5127
R2455 VDD.n2259 VDD.n415 99.5127
R2456 VDD.n2259 VDD.n405 99.5127
R2457 VDD.n2267 VDD.n405 99.5127
R2458 VDD.n2267 VDD.n403 99.5127
R2459 VDD.n2271 VDD.n403 99.5127
R2460 VDD.n2271 VDD.n393 99.5127
R2461 VDD.n2279 VDD.n393 99.5127
R2462 VDD.n2279 VDD.n391 99.5127
R2463 VDD.n2283 VDD.n391 99.5127
R2464 VDD.n2283 VDD.n381 99.5127
R2465 VDD.n2291 VDD.n381 99.5127
R2466 VDD.n2291 VDD.n379 99.5127
R2467 VDD.n2295 VDD.n379 99.5127
R2468 VDD.n2295 VDD.n369 99.5127
R2469 VDD.n2303 VDD.n369 99.5127
R2470 VDD.n2303 VDD.n367 99.5127
R2471 VDD.n2307 VDD.n367 99.5127
R2472 VDD.n2307 VDD.n357 99.5127
R2473 VDD.n2315 VDD.n357 99.5127
R2474 VDD.n2315 VDD.n355 99.5127
R2475 VDD.n2319 VDD.n355 99.5127
R2476 VDD.n2319 VDD.n345 99.5127
R2477 VDD.n2327 VDD.n345 99.5127
R2478 VDD.n2327 VDD.n343 99.5127
R2479 VDD.n2331 VDD.n343 99.5127
R2480 VDD.n2331 VDD.n333 99.5127
R2481 VDD.n2339 VDD.n333 99.5127
R2482 VDD.n2339 VDD.n331 99.5127
R2483 VDD.n2343 VDD.n331 99.5127
R2484 VDD.n2343 VDD.n320 99.5127
R2485 VDD.n2351 VDD.n320 99.5127
R2486 VDD.n2351 VDD.n318 99.5127
R2487 VDD.n2355 VDD.n318 99.5127
R2488 VDD.n2355 VDD.n308 99.5127
R2489 VDD.n2363 VDD.n308 99.5127
R2490 VDD.n2363 VDD.n306 99.5127
R2491 VDD.n2367 VDD.n306 99.5127
R2492 VDD.n2367 VDD.n297 99.5127
R2493 VDD.n2375 VDD.n297 99.5127
R2494 VDD.n2375 VDD.n295 99.5127
R2495 VDD.n2379 VDD.n295 99.5127
R2496 VDD.n2379 VDD.n285 99.5127
R2497 VDD.n2387 VDD.n285 99.5127
R2498 VDD.n2387 VDD.n283 99.5127
R2499 VDD.n2391 VDD.n283 99.5127
R2500 VDD.n2391 VDD.n273 99.5127
R2501 VDD.n2399 VDD.n273 99.5127
R2502 VDD.n2399 VDD.n271 99.5127
R2503 VDD.n2403 VDD.n271 99.5127
R2504 VDD.n2403 VDD.n261 99.5127
R2505 VDD.n2411 VDD.n261 99.5127
R2506 VDD.n2411 VDD.n259 99.5127
R2507 VDD.n2415 VDD.n259 99.5127
R2508 VDD.n2415 VDD.n249 99.5127
R2509 VDD.n2423 VDD.n249 99.5127
R2510 VDD.n2423 VDD.n247 99.5127
R2511 VDD.n2427 VDD.n247 99.5127
R2512 VDD.n2427 VDD.n237 99.5127
R2513 VDD.n2435 VDD.n237 99.5127
R2514 VDD.n2435 VDD.n235 99.5127
R2515 VDD.n2439 VDD.n235 99.5127
R2516 VDD.n2439 VDD.n225 99.5127
R2517 VDD.n2447 VDD.n225 99.5127
R2518 VDD.n2447 VDD.n223 99.5127
R2519 VDD.n2451 VDD.n223 99.5127
R2520 VDD.n2451 VDD.n213 99.5127
R2521 VDD.n2459 VDD.n213 99.5127
R2522 VDD.n2459 VDD.n211 99.5127
R2523 VDD.n2463 VDD.n211 99.5127
R2524 VDD.n2463 VDD.n201 99.5127
R2525 VDD.n2471 VDD.n201 99.5127
R2526 VDD.n2471 VDD.n199 99.5127
R2527 VDD.n2475 VDD.n199 99.5127
R2528 VDD.n2475 VDD.n189 99.5127
R2529 VDD.n2483 VDD.n189 99.5127
R2530 VDD.n2483 VDD.n187 99.5127
R2531 VDD.n2487 VDD.n187 99.5127
R2532 VDD.n2487 VDD.n176 99.5127
R2533 VDD.n2495 VDD.n176 99.5127
R2534 VDD.n2495 VDD.n174 99.5127
R2535 VDD.n2499 VDD.n174 99.5127
R2536 VDD.n2499 VDD.n164 99.5127
R2537 VDD.n2529 VDD.n164 99.5127
R2538 VDD.n2529 VDD.n162 99.5127
R2539 VDD.n2533 VDD.n162 99.5127
R2540 VDD.n2533 VDD.n140 99.5127
R2541 VDD.n2570 VDD.n140 99.5127
R2542 VDD.n2570 VDD.n141 99.5127
R2543 VDD.n1908 VDD.n441 99.5127
R2544 VDD.n1904 VDD.n1903 99.5127
R2545 VDD.n1900 VDD.n1899 99.5127
R2546 VDD.n1896 VDD.n1895 99.5127
R2547 VDD.n1892 VDD.n1891 99.5127
R2548 VDD.n1888 VDD.n1887 99.5127
R2549 VDD.n1884 VDD.n1883 99.5127
R2550 VDD.n1538 VDD.n719 99.5127
R2551 VDD.n1534 VDD.n719 99.5127
R2552 VDD.n1534 VDD.n713 99.5127
R2553 VDD.n1531 VDD.n713 99.5127
R2554 VDD.n1531 VDD.n707 99.5127
R2555 VDD.n1528 VDD.n707 99.5127
R2556 VDD.n1528 VDD.n701 99.5127
R2557 VDD.n1525 VDD.n701 99.5127
R2558 VDD.n1525 VDD.n695 99.5127
R2559 VDD.n1522 VDD.n695 99.5127
R2560 VDD.n1522 VDD.n689 99.5127
R2561 VDD.n1519 VDD.n689 99.5127
R2562 VDD.n1519 VDD.n683 99.5127
R2563 VDD.n1516 VDD.n683 99.5127
R2564 VDD.n1516 VDD.n677 99.5127
R2565 VDD.n1513 VDD.n677 99.5127
R2566 VDD.n1513 VDD.n671 99.5127
R2567 VDD.n1510 VDD.n671 99.5127
R2568 VDD.n1510 VDD.n665 99.5127
R2569 VDD.n1507 VDD.n665 99.5127
R2570 VDD.n1507 VDD.n659 99.5127
R2571 VDD.n1504 VDD.n659 99.5127
R2572 VDD.n1504 VDD.n652 99.5127
R2573 VDD.n1501 VDD.n652 99.5127
R2574 VDD.n1501 VDD.n646 99.5127
R2575 VDD.n1498 VDD.n646 99.5127
R2576 VDD.n1498 VDD.n641 99.5127
R2577 VDD.n1495 VDD.n641 99.5127
R2578 VDD.n1495 VDD.n635 99.5127
R2579 VDD.n1492 VDD.n635 99.5127
R2580 VDD.n1492 VDD.n629 99.5127
R2581 VDD.n1489 VDD.n629 99.5127
R2582 VDD.n1489 VDD.n623 99.5127
R2583 VDD.n1486 VDD.n623 99.5127
R2584 VDD.n1486 VDD.n617 99.5127
R2585 VDD.n1483 VDD.n617 99.5127
R2586 VDD.n1483 VDD.n610 99.5127
R2587 VDD.n1480 VDD.n610 99.5127
R2588 VDD.n1480 VDD.n604 99.5127
R2589 VDD.n1477 VDD.n604 99.5127
R2590 VDD.n1477 VDD.n598 99.5127
R2591 VDD.n1474 VDD.n598 99.5127
R2592 VDD.n1474 VDD.n592 99.5127
R2593 VDD.n1471 VDD.n592 99.5127
R2594 VDD.n1471 VDD.n587 99.5127
R2595 VDD.n1468 VDD.n587 99.5127
R2596 VDD.n1468 VDD.n581 99.5127
R2597 VDD.n1465 VDD.n581 99.5127
R2598 VDD.n1465 VDD.n575 99.5127
R2599 VDD.n1462 VDD.n575 99.5127
R2600 VDD.n1462 VDD.n569 99.5127
R2601 VDD.n1459 VDD.n569 99.5127
R2602 VDD.n1459 VDD.n563 99.5127
R2603 VDD.n1456 VDD.n563 99.5127
R2604 VDD.n1456 VDD.n557 99.5127
R2605 VDD.n1453 VDD.n557 99.5127
R2606 VDD.n1453 VDD.n551 99.5127
R2607 VDD.n1450 VDD.n551 99.5127
R2608 VDD.n1450 VDD.n545 99.5127
R2609 VDD.n1447 VDD.n545 99.5127
R2610 VDD.n1447 VDD.n539 99.5127
R2611 VDD.n1444 VDD.n539 99.5127
R2612 VDD.n1444 VDD.n533 99.5127
R2613 VDD.n1441 VDD.n533 99.5127
R2614 VDD.n1441 VDD.n527 99.5127
R2615 VDD.n1438 VDD.n527 99.5127
R2616 VDD.n1438 VDD.n521 99.5127
R2617 VDD.n1435 VDD.n521 99.5127
R2618 VDD.n1435 VDD.n515 99.5127
R2619 VDD.n1432 VDD.n515 99.5127
R2620 VDD.n1432 VDD.n509 99.5127
R2621 VDD.n1429 VDD.n509 99.5127
R2622 VDD.n1429 VDD.n503 99.5127
R2623 VDD.n1426 VDD.n503 99.5127
R2624 VDD.n1426 VDD.n497 99.5127
R2625 VDD.n1423 VDD.n497 99.5127
R2626 VDD.n1423 VDD.n491 99.5127
R2627 VDD.n1420 VDD.n491 99.5127
R2628 VDD.n1420 VDD.n485 99.5127
R2629 VDD.n1417 VDD.n485 99.5127
R2630 VDD.n1417 VDD.n478 99.5127
R2631 VDD.n1414 VDD.n478 99.5127
R2632 VDD.n1414 VDD.n471 99.5127
R2633 VDD.n1411 VDD.n471 99.5127
R2634 VDD.n1411 VDD.n466 99.5127
R2635 VDD.n1408 VDD.n466 99.5127
R2636 VDD.n1408 VDD.n456 99.5127
R2637 VDD.n456 VDD.n447 99.5127
R2638 VDD.n1878 VDD.n447 99.5127
R2639 VDD.n1879 VDD.n1878 99.5127
R2640 VDD.n1563 VDD.n723 99.5127
R2641 VDD.n1563 VDD.n738 99.5127
R2642 VDD.n1559 VDD.n1558 99.5127
R2643 VDD.n1555 VDD.n1554 99.5127
R2644 VDD.n1551 VDD.n1550 99.5127
R2645 VDD.n1547 VDD.n1546 99.5127
R2646 VDD.n1543 VDD.n1542 99.5127
R2647 VDD.n1570 VDD.n721 99.5127
R2648 VDD.n1570 VDD.n711 99.5127
R2649 VDD.n1578 VDD.n711 99.5127
R2650 VDD.n1578 VDD.n709 99.5127
R2651 VDD.n1582 VDD.n709 99.5127
R2652 VDD.n1582 VDD.n699 99.5127
R2653 VDD.n1590 VDD.n699 99.5127
R2654 VDD.n1590 VDD.n697 99.5127
R2655 VDD.n1594 VDD.n697 99.5127
R2656 VDD.n1594 VDD.n687 99.5127
R2657 VDD.n1602 VDD.n687 99.5127
R2658 VDD.n1602 VDD.n685 99.5127
R2659 VDD.n1606 VDD.n685 99.5127
R2660 VDD.n1606 VDD.n675 99.5127
R2661 VDD.n1614 VDD.n675 99.5127
R2662 VDD.n1614 VDD.n673 99.5127
R2663 VDD.n1618 VDD.n673 99.5127
R2664 VDD.n1618 VDD.n663 99.5127
R2665 VDD.n1626 VDD.n663 99.5127
R2666 VDD.n1626 VDD.n661 99.5127
R2667 VDD.n1630 VDD.n661 99.5127
R2668 VDD.n1630 VDD.n650 99.5127
R2669 VDD.n1638 VDD.n650 99.5127
R2670 VDD.n1638 VDD.n648 99.5127
R2671 VDD.n1642 VDD.n648 99.5127
R2672 VDD.n1642 VDD.n639 99.5127
R2673 VDD.n1650 VDD.n639 99.5127
R2674 VDD.n1650 VDD.n637 99.5127
R2675 VDD.n1654 VDD.n637 99.5127
R2676 VDD.n1654 VDD.n627 99.5127
R2677 VDD.n1662 VDD.n627 99.5127
R2678 VDD.n1662 VDD.n625 99.5127
R2679 VDD.n1666 VDD.n625 99.5127
R2680 VDD.n1666 VDD.n615 99.5127
R2681 VDD.n1674 VDD.n615 99.5127
R2682 VDD.n1674 VDD.n613 99.5127
R2683 VDD.n1678 VDD.n613 99.5127
R2684 VDD.n1678 VDD.n603 99.5127
R2685 VDD.n1686 VDD.n603 99.5127
R2686 VDD.n1686 VDD.n601 99.5127
R2687 VDD.n1690 VDD.n601 99.5127
R2688 VDD.n1690 VDD.n591 99.5127
R2689 VDD.n1698 VDD.n591 99.5127
R2690 VDD.n1698 VDD.n589 99.5127
R2691 VDD.n1702 VDD.n589 99.5127
R2692 VDD.n1702 VDD.n579 99.5127
R2693 VDD.n1710 VDD.n579 99.5127
R2694 VDD.n1710 VDD.n577 99.5127
R2695 VDD.n1714 VDD.n577 99.5127
R2696 VDD.n1714 VDD.n567 99.5127
R2697 VDD.n1722 VDD.n567 99.5127
R2698 VDD.n1722 VDD.n565 99.5127
R2699 VDD.n1726 VDD.n565 99.5127
R2700 VDD.n1726 VDD.n555 99.5127
R2701 VDD.n1734 VDD.n555 99.5127
R2702 VDD.n1734 VDD.n553 99.5127
R2703 VDD.n1738 VDD.n553 99.5127
R2704 VDD.n1738 VDD.n543 99.5127
R2705 VDD.n1746 VDD.n543 99.5127
R2706 VDD.n1746 VDD.n541 99.5127
R2707 VDD.n1750 VDD.n541 99.5127
R2708 VDD.n1750 VDD.n531 99.5127
R2709 VDD.n1758 VDD.n531 99.5127
R2710 VDD.n1758 VDD.n529 99.5127
R2711 VDD.n1762 VDD.n529 99.5127
R2712 VDD.n1762 VDD.n519 99.5127
R2713 VDD.n1770 VDD.n519 99.5127
R2714 VDD.n1770 VDD.n517 99.5127
R2715 VDD.n1774 VDD.n517 99.5127
R2716 VDD.n1774 VDD.n507 99.5127
R2717 VDD.n1782 VDD.n507 99.5127
R2718 VDD.n1782 VDD.n505 99.5127
R2719 VDD.n1786 VDD.n505 99.5127
R2720 VDD.n1786 VDD.n495 99.5127
R2721 VDD.n1794 VDD.n495 99.5127
R2722 VDD.n1794 VDD.n493 99.5127
R2723 VDD.n1798 VDD.n493 99.5127
R2724 VDD.n1798 VDD.n483 99.5127
R2725 VDD.n1806 VDD.n483 99.5127
R2726 VDD.n1806 VDD.n481 99.5127
R2727 VDD.n1810 VDD.n481 99.5127
R2728 VDD.n1810 VDD.n470 99.5127
R2729 VDD.n1820 VDD.n470 99.5127
R2730 VDD.n1820 VDD.n468 99.5127
R2731 VDD.n1824 VDD.n468 99.5127
R2732 VDD.n1824 VDD.n454 99.5127
R2733 VDD.n1872 VDD.n454 99.5127
R2734 VDD.n1872 VDD.n452 99.5127
R2735 VDD.n1876 VDD.n452 99.5127
R2736 VDD.n1876 VDD.n440 99.5127
R2737 VDD.n2518 VDD.n2517 99.5127
R2738 VDD.n2515 VDD.n2506 99.5127
R2739 VDD.n2511 VDD.n2510 99.5127
R2740 VDD.n2588 VDD.n124 99.5127
R2741 VDD.n2586 VDD.n2585 99.5127
R2742 VDD.n2583 VDD.n127 99.5127
R2743 VDD.n2579 VDD.n2578 99.5127
R2744 VDD.n1923 VDD.n420 99.5127
R2745 VDD.n2077 VDD.n420 99.5127
R2746 VDD.n2077 VDD.n414 99.5127
R2747 VDD.n2074 VDD.n414 99.5127
R2748 VDD.n2074 VDD.n408 99.5127
R2749 VDD.n2071 VDD.n408 99.5127
R2750 VDD.n2071 VDD.n402 99.5127
R2751 VDD.n2068 VDD.n402 99.5127
R2752 VDD.n2068 VDD.n396 99.5127
R2753 VDD.n2065 VDD.n396 99.5127
R2754 VDD.n2065 VDD.n390 99.5127
R2755 VDD.n2062 VDD.n390 99.5127
R2756 VDD.n2062 VDD.n384 99.5127
R2757 VDD.n2059 VDD.n384 99.5127
R2758 VDD.n2059 VDD.n378 99.5127
R2759 VDD.n2056 VDD.n378 99.5127
R2760 VDD.n2056 VDD.n372 99.5127
R2761 VDD.n2053 VDD.n372 99.5127
R2762 VDD.n2053 VDD.n365 99.5127
R2763 VDD.n2050 VDD.n365 99.5127
R2764 VDD.n2050 VDD.n359 99.5127
R2765 VDD.n2047 VDD.n359 99.5127
R2766 VDD.n2047 VDD.n353 99.5127
R2767 VDD.n2044 VDD.n353 99.5127
R2768 VDD.n2044 VDD.n347 99.5127
R2769 VDD.n2041 VDD.n347 99.5127
R2770 VDD.n2041 VDD.n342 99.5127
R2771 VDD.n2038 VDD.n342 99.5127
R2772 VDD.n2038 VDD.n336 99.5127
R2773 VDD.n2035 VDD.n336 99.5127
R2774 VDD.n2035 VDD.n330 99.5127
R2775 VDD.n2032 VDD.n330 99.5127
R2776 VDD.n2032 VDD.n323 99.5127
R2777 VDD.n2029 VDD.n323 99.5127
R2778 VDD.n2029 VDD.n317 99.5127
R2779 VDD.n2026 VDD.n317 99.5127
R2780 VDD.n2026 VDD.n311 99.5127
R2781 VDD.n2023 VDD.n311 99.5127
R2782 VDD.n2023 VDD.n305 99.5127
R2783 VDD.n2020 VDD.n305 99.5127
R2784 VDD.n2020 VDD.n300 99.5127
R2785 VDD.n2017 VDD.n300 99.5127
R2786 VDD.n2017 VDD.n294 99.5127
R2787 VDD.n2014 VDD.n294 99.5127
R2788 VDD.n2014 VDD.n288 99.5127
R2789 VDD.n2011 VDD.n288 99.5127
R2790 VDD.n2011 VDD.n282 99.5127
R2791 VDD.n2008 VDD.n282 99.5127
R2792 VDD.n2008 VDD.n276 99.5127
R2793 VDD.n2005 VDD.n276 99.5127
R2794 VDD.n2005 VDD.n270 99.5127
R2795 VDD.n2002 VDD.n270 99.5127
R2796 VDD.n2002 VDD.n264 99.5127
R2797 VDD.n1999 VDD.n264 99.5127
R2798 VDD.n1999 VDD.n258 99.5127
R2799 VDD.n1996 VDD.n258 99.5127
R2800 VDD.n1996 VDD.n252 99.5127
R2801 VDD.n1993 VDD.n252 99.5127
R2802 VDD.n1993 VDD.n246 99.5127
R2803 VDD.n1990 VDD.n246 99.5127
R2804 VDD.n1990 VDD.n240 99.5127
R2805 VDD.n1987 VDD.n240 99.5127
R2806 VDD.n1987 VDD.n234 99.5127
R2807 VDD.n1984 VDD.n234 99.5127
R2808 VDD.n1984 VDD.n228 99.5127
R2809 VDD.n1981 VDD.n228 99.5127
R2810 VDD.n1981 VDD.n221 99.5127
R2811 VDD.n1978 VDD.n221 99.5127
R2812 VDD.n1978 VDD.n215 99.5127
R2813 VDD.n1975 VDD.n215 99.5127
R2814 VDD.n1975 VDD.n210 99.5127
R2815 VDD.n1972 VDD.n210 99.5127
R2816 VDD.n1972 VDD.n204 99.5127
R2817 VDD.n1969 VDD.n204 99.5127
R2818 VDD.n1969 VDD.n198 99.5127
R2819 VDD.n1966 VDD.n198 99.5127
R2820 VDD.n1966 VDD.n192 99.5127
R2821 VDD.n1963 VDD.n192 99.5127
R2822 VDD.n1963 VDD.n186 99.5127
R2823 VDD.n1960 VDD.n186 99.5127
R2824 VDD.n1960 VDD.n179 99.5127
R2825 VDD.n1957 VDD.n179 99.5127
R2826 VDD.n1957 VDD.n173 99.5127
R2827 VDD.n1954 VDD.n173 99.5127
R2828 VDD.n1954 VDD.n167 99.5127
R2829 VDD.n1951 VDD.n167 99.5127
R2830 VDD.n1951 VDD.n160 99.5127
R2831 VDD.n160 VDD.n135 99.5127
R2832 VDD.n2572 VDD.n135 99.5127
R2833 VDD.n2572 VDD.n133 99.5127
R2834 VDD.n1926 VDD.n423 99.5127
R2835 VDD.n1930 VDD.n1929 99.5127
R2836 VDD.n1934 VDD.n1933 99.5127
R2837 VDD.n1938 VDD.n1937 99.5127
R2838 VDD.n1942 VDD.n1941 99.5127
R2839 VDD.n1946 VDD.n1945 99.5127
R2840 VDD.n2082 VDD.n1922 99.5127
R2841 VDD.n2253 VDD.n421 99.5127
R2842 VDD.n2253 VDD.n411 99.5127
R2843 VDD.n2261 VDD.n411 99.5127
R2844 VDD.n2261 VDD.n409 99.5127
R2845 VDD.n2265 VDD.n409 99.5127
R2846 VDD.n2265 VDD.n399 99.5127
R2847 VDD.n2273 VDD.n399 99.5127
R2848 VDD.n2273 VDD.n397 99.5127
R2849 VDD.n2277 VDD.n397 99.5127
R2850 VDD.n2277 VDD.n387 99.5127
R2851 VDD.n2285 VDD.n387 99.5127
R2852 VDD.n2285 VDD.n385 99.5127
R2853 VDD.n2289 VDD.n385 99.5127
R2854 VDD.n2289 VDD.n375 99.5127
R2855 VDD.n2297 VDD.n375 99.5127
R2856 VDD.n2297 VDD.n373 99.5127
R2857 VDD.n2301 VDD.n373 99.5127
R2858 VDD.n2301 VDD.n362 99.5127
R2859 VDD.n2309 VDD.n362 99.5127
R2860 VDD.n2309 VDD.n360 99.5127
R2861 VDD.n2313 VDD.n360 99.5127
R2862 VDD.n2313 VDD.n350 99.5127
R2863 VDD.n2321 VDD.n350 99.5127
R2864 VDD.n2321 VDD.n348 99.5127
R2865 VDD.n2325 VDD.n348 99.5127
R2866 VDD.n2325 VDD.n339 99.5127
R2867 VDD.n2333 VDD.n339 99.5127
R2868 VDD.n2333 VDD.n337 99.5127
R2869 VDD.n2337 VDD.n337 99.5127
R2870 VDD.n2337 VDD.n327 99.5127
R2871 VDD.n2345 VDD.n327 99.5127
R2872 VDD.n2345 VDD.n325 99.5127
R2873 VDD.n2349 VDD.n325 99.5127
R2874 VDD.n2349 VDD.n315 99.5127
R2875 VDD.n2357 VDD.n315 99.5127
R2876 VDD.n2357 VDD.n313 99.5127
R2877 VDD.n2361 VDD.n313 99.5127
R2878 VDD.n2361 VDD.n303 99.5127
R2879 VDD.n2369 VDD.n303 99.5127
R2880 VDD.n2369 VDD.n301 99.5127
R2881 VDD.n2373 VDD.n301 99.5127
R2882 VDD.n2373 VDD.n291 99.5127
R2883 VDD.n2381 VDD.n291 99.5127
R2884 VDD.n2381 VDD.n289 99.5127
R2885 VDD.n2385 VDD.n289 99.5127
R2886 VDD.n2385 VDD.n279 99.5127
R2887 VDD.n2393 VDD.n279 99.5127
R2888 VDD.n2393 VDD.n277 99.5127
R2889 VDD.n2397 VDD.n277 99.5127
R2890 VDD.n2397 VDD.n267 99.5127
R2891 VDD.n2405 VDD.n267 99.5127
R2892 VDD.n2405 VDD.n265 99.5127
R2893 VDD.n2409 VDD.n265 99.5127
R2894 VDD.n2409 VDD.n255 99.5127
R2895 VDD.n2417 VDD.n255 99.5127
R2896 VDD.n2417 VDD.n253 99.5127
R2897 VDD.n2421 VDD.n253 99.5127
R2898 VDD.n2421 VDD.n243 99.5127
R2899 VDD.n2429 VDD.n243 99.5127
R2900 VDD.n2429 VDD.n241 99.5127
R2901 VDD.n2433 VDD.n241 99.5127
R2902 VDD.n2433 VDD.n231 99.5127
R2903 VDD.n2441 VDD.n231 99.5127
R2904 VDD.n2441 VDD.n229 99.5127
R2905 VDD.n2445 VDD.n229 99.5127
R2906 VDD.n2445 VDD.n218 99.5127
R2907 VDD.n2453 VDD.n218 99.5127
R2908 VDD.n2453 VDD.n216 99.5127
R2909 VDD.n2457 VDD.n216 99.5127
R2910 VDD.n2457 VDD.n207 99.5127
R2911 VDD.n2465 VDD.n207 99.5127
R2912 VDD.n2465 VDD.n205 99.5127
R2913 VDD.n2469 VDD.n205 99.5127
R2914 VDD.n2469 VDD.n195 99.5127
R2915 VDD.n2477 VDD.n195 99.5127
R2916 VDD.n2477 VDD.n193 99.5127
R2917 VDD.n2481 VDD.n193 99.5127
R2918 VDD.n2481 VDD.n183 99.5127
R2919 VDD.n2489 VDD.n183 99.5127
R2920 VDD.n2489 VDD.n181 99.5127
R2921 VDD.n2493 VDD.n181 99.5127
R2922 VDD.n2493 VDD.n171 99.5127
R2923 VDD.n2501 VDD.n171 99.5127
R2924 VDD.n2501 VDD.n168 99.5127
R2925 VDD.n2527 VDD.n168 99.5127
R2926 VDD.n2527 VDD.n169 99.5127
R2927 VDD.n169 VDD.n161 99.5127
R2928 VDD.n2522 VDD.n161 99.5127
R2929 VDD.n2522 VDD.n139 99.5127
R2930 VDD.n2519 VDD.n139 99.5127
R2931 VDD.n1861 VDD.n1860 99.5127
R2932 VDD.n1857 VDD.n1856 99.5127
R2933 VDD.n1853 VDD.n1852 99.5127
R2934 VDD.n1849 VDD.n1848 99.5127
R2935 VDD.n1845 VDD.n1844 99.5127
R2936 VDD.n1841 VDD.n1840 99.5127
R2937 VDD.n1836 VDD.n432 99.5127
R2938 VDD.n933 VDD.n720 99.5127
R2939 VDD.n930 VDD.n720 99.5127
R2940 VDD.n930 VDD.n714 99.5127
R2941 VDD.n927 VDD.n714 99.5127
R2942 VDD.n927 VDD.n708 99.5127
R2943 VDD.n924 VDD.n708 99.5127
R2944 VDD.n924 VDD.n702 99.5127
R2945 VDD.n921 VDD.n702 99.5127
R2946 VDD.n921 VDD.n696 99.5127
R2947 VDD.n918 VDD.n696 99.5127
R2948 VDD.n918 VDD.n690 99.5127
R2949 VDD.n915 VDD.n690 99.5127
R2950 VDD.n915 VDD.n684 99.5127
R2951 VDD.n912 VDD.n684 99.5127
R2952 VDD.n912 VDD.n678 99.5127
R2953 VDD.n909 VDD.n678 99.5127
R2954 VDD.n909 VDD.n672 99.5127
R2955 VDD.n906 VDD.n672 99.5127
R2956 VDD.n906 VDD.n666 99.5127
R2957 VDD.n903 VDD.n666 99.5127
R2958 VDD.n903 VDD.n660 99.5127
R2959 VDD.n900 VDD.n660 99.5127
R2960 VDD.n900 VDD.n653 99.5127
R2961 VDD.n897 VDD.n653 99.5127
R2962 VDD.n897 VDD.n647 99.5127
R2963 VDD.n894 VDD.n647 99.5127
R2964 VDD.n894 VDD.n642 99.5127
R2965 VDD.n891 VDD.n642 99.5127
R2966 VDD.n891 VDD.n636 99.5127
R2967 VDD.n888 VDD.n636 99.5127
R2968 VDD.n888 VDD.n630 99.5127
R2969 VDD.n885 VDD.n630 99.5127
R2970 VDD.n885 VDD.n624 99.5127
R2971 VDD.n882 VDD.n624 99.5127
R2972 VDD.n882 VDD.n618 99.5127
R2973 VDD.n879 VDD.n618 99.5127
R2974 VDD.n879 VDD.n611 99.5127
R2975 VDD.n876 VDD.n611 99.5127
R2976 VDD.n876 VDD.n605 99.5127
R2977 VDD.n873 VDD.n605 99.5127
R2978 VDD.n873 VDD.n599 99.5127
R2979 VDD.n870 VDD.n599 99.5127
R2980 VDD.n870 VDD.n593 99.5127
R2981 VDD.n867 VDD.n593 99.5127
R2982 VDD.n867 VDD.n588 99.5127
R2983 VDD.n864 VDD.n588 99.5127
R2984 VDD.n864 VDD.n582 99.5127
R2985 VDD.n861 VDD.n582 99.5127
R2986 VDD.n861 VDD.n576 99.5127
R2987 VDD.n858 VDD.n576 99.5127
R2988 VDD.n858 VDD.n570 99.5127
R2989 VDD.n855 VDD.n570 99.5127
R2990 VDD.n855 VDD.n564 99.5127
R2991 VDD.n852 VDD.n564 99.5127
R2992 VDD.n852 VDD.n558 99.5127
R2993 VDD.n849 VDD.n558 99.5127
R2994 VDD.n849 VDD.n552 99.5127
R2995 VDD.n846 VDD.n552 99.5127
R2996 VDD.n846 VDD.n546 99.5127
R2997 VDD.n843 VDD.n546 99.5127
R2998 VDD.n843 VDD.n540 99.5127
R2999 VDD.n840 VDD.n540 99.5127
R3000 VDD.n840 VDD.n534 99.5127
R3001 VDD.n837 VDD.n534 99.5127
R3002 VDD.n837 VDD.n528 99.5127
R3003 VDD.n834 VDD.n528 99.5127
R3004 VDD.n834 VDD.n522 99.5127
R3005 VDD.n831 VDD.n522 99.5127
R3006 VDD.n831 VDD.n516 99.5127
R3007 VDD.n828 VDD.n516 99.5127
R3008 VDD.n828 VDD.n510 99.5127
R3009 VDD.n825 VDD.n510 99.5127
R3010 VDD.n825 VDD.n504 99.5127
R3011 VDD.n822 VDD.n504 99.5127
R3012 VDD.n822 VDD.n498 99.5127
R3013 VDD.n819 VDD.n498 99.5127
R3014 VDD.n819 VDD.n492 99.5127
R3015 VDD.n816 VDD.n492 99.5127
R3016 VDD.n816 VDD.n486 99.5127
R3017 VDD.n813 VDD.n486 99.5127
R3018 VDD.n813 VDD.n479 99.5127
R3019 VDD.n810 VDD.n479 99.5127
R3020 VDD.n810 VDD.n472 99.5127
R3021 VDD.n472 VDD.n464 99.5127
R3022 VDD.n1826 VDD.n464 99.5127
R3023 VDD.n1827 VDD.n1826 99.5127
R3024 VDD.n1827 VDD.n457 99.5127
R3025 VDD.n1830 VDD.n457 99.5127
R3026 VDD.n1830 VDD.n450 99.5127
R3027 VDD.n1833 VDD.n450 99.5127
R3028 VDD.n795 VDD.n794 99.5127
R3029 VDD.n799 VDD.n798 99.5127
R3030 VDD.n803 VDD.n802 99.5127
R3031 VDD.n947 VDD.n805 99.5127
R3032 VDD.n945 VDD.n944 99.5127
R3033 VDD.n941 VDD.n940 99.5127
R3034 VDD.n936 VDD.n737 99.5127
R3035 VDD.n1572 VDD.n717 99.5127
R3036 VDD.n1572 VDD.n715 99.5127
R3037 VDD.n1576 VDD.n715 99.5127
R3038 VDD.n1576 VDD.n705 99.5127
R3039 VDD.n1584 VDD.n705 99.5127
R3040 VDD.n1584 VDD.n703 99.5127
R3041 VDD.n1588 VDD.n703 99.5127
R3042 VDD.n1588 VDD.n693 99.5127
R3043 VDD.n1596 VDD.n693 99.5127
R3044 VDD.n1596 VDD.n691 99.5127
R3045 VDD.n1600 VDD.n691 99.5127
R3046 VDD.n1600 VDD.n681 99.5127
R3047 VDD.n1608 VDD.n681 99.5127
R3048 VDD.n1608 VDD.n679 99.5127
R3049 VDD.n1612 VDD.n679 99.5127
R3050 VDD.n1612 VDD.n669 99.5127
R3051 VDD.n1620 VDD.n669 99.5127
R3052 VDD.n1620 VDD.n667 99.5127
R3053 VDD.n1624 VDD.n667 99.5127
R3054 VDD.n1624 VDD.n657 99.5127
R3055 VDD.n1632 VDD.n657 99.5127
R3056 VDD.n1632 VDD.n655 99.5127
R3057 VDD.n1636 VDD.n655 99.5127
R3058 VDD.n1636 VDD.n645 99.5127
R3059 VDD.n1644 VDD.n645 99.5127
R3060 VDD.n1644 VDD.n643 99.5127
R3061 VDD.n1648 VDD.n643 99.5127
R3062 VDD.n1648 VDD.n633 99.5127
R3063 VDD.n1656 VDD.n633 99.5127
R3064 VDD.n1656 VDD.n631 99.5127
R3065 VDD.n1660 VDD.n631 99.5127
R3066 VDD.n1660 VDD.n621 99.5127
R3067 VDD.n1668 VDD.n621 99.5127
R3068 VDD.n1668 VDD.n619 99.5127
R3069 VDD.n1672 VDD.n619 99.5127
R3070 VDD.n1672 VDD.n608 99.5127
R3071 VDD.n1680 VDD.n608 99.5127
R3072 VDD.n1680 VDD.n606 99.5127
R3073 VDD.n1684 VDD.n606 99.5127
R3074 VDD.n1684 VDD.n596 99.5127
R3075 VDD.n1692 VDD.n596 99.5127
R3076 VDD.n1692 VDD.n594 99.5127
R3077 VDD.n1696 VDD.n594 99.5127
R3078 VDD.n1696 VDD.n585 99.5127
R3079 VDD.n1704 VDD.n585 99.5127
R3080 VDD.n1704 VDD.n583 99.5127
R3081 VDD.n1708 VDD.n583 99.5127
R3082 VDD.n1708 VDD.n573 99.5127
R3083 VDD.n1716 VDD.n573 99.5127
R3084 VDD.n1716 VDD.n571 99.5127
R3085 VDD.n1720 VDD.n571 99.5127
R3086 VDD.n1720 VDD.n561 99.5127
R3087 VDD.n1728 VDD.n561 99.5127
R3088 VDD.n1728 VDD.n559 99.5127
R3089 VDD.n1732 VDD.n559 99.5127
R3090 VDD.n1732 VDD.n549 99.5127
R3091 VDD.n1740 VDD.n549 99.5127
R3092 VDD.n1740 VDD.n547 99.5127
R3093 VDD.n1744 VDD.n547 99.5127
R3094 VDD.n1744 VDD.n537 99.5127
R3095 VDD.n1752 VDD.n537 99.5127
R3096 VDD.n1752 VDD.n535 99.5127
R3097 VDD.n1756 VDD.n535 99.5127
R3098 VDD.n1756 VDD.n525 99.5127
R3099 VDD.n1764 VDD.n525 99.5127
R3100 VDD.n1764 VDD.n523 99.5127
R3101 VDD.n1768 VDD.n523 99.5127
R3102 VDD.n1768 VDD.n513 99.5127
R3103 VDD.n1776 VDD.n513 99.5127
R3104 VDD.n1776 VDD.n511 99.5127
R3105 VDD.n1780 VDD.n511 99.5127
R3106 VDD.n1780 VDD.n501 99.5127
R3107 VDD.n1788 VDD.n501 99.5127
R3108 VDD.n1788 VDD.n499 99.5127
R3109 VDD.n1792 VDD.n499 99.5127
R3110 VDD.n1792 VDD.n489 99.5127
R3111 VDD.n1800 VDD.n489 99.5127
R3112 VDD.n1800 VDD.n487 99.5127
R3113 VDD.n1804 VDD.n487 99.5127
R3114 VDD.n1804 VDD.n476 99.5127
R3115 VDD.n1812 VDD.n476 99.5127
R3116 VDD.n1812 VDD.n473 99.5127
R3117 VDD.n1818 VDD.n473 99.5127
R3118 VDD.n1818 VDD.n474 99.5127
R3119 VDD.n474 VDD.n467 99.5127
R3120 VDD.n467 VDD.n458 99.5127
R3121 VDD.n1870 VDD.n458 99.5127
R3122 VDD.n1870 VDD.n459 99.5127
R3123 VDD.n459 VDD.n451 99.5127
R3124 VDD.n1865 VDD.n451 99.5127
R3125 VDD.n2986 VDD.t1 98.1472
R3126 VDD.n2985 VDD.t74 98.1472
R3127 VDD.n807 VDD.n806 89.4066
R3128 VDD.n462 VDD.n461 89.4066
R3129 VDD.n1404 VDD.n1403 89.4066
R3130 VDD.n444 VDD.n443 89.4066
R3131 VDD.n1925 VDD.n1924 89.4066
R3132 VDD.n152 VDD.n151 89.4066
R3133 VDD.n2086 VDD.n2085 89.4066
R3134 VDD.n129 VDD.n128 89.4066
R3135 VDD.n2248 VDD.n2247 72.8958
R3136 VDD.n2247 VDD.n1916 72.8958
R3137 VDD.n2247 VDD.n1917 72.8958
R3138 VDD.n2247 VDD.n1918 72.8958
R3139 VDD.n2247 VDD.n1919 72.8958
R3140 VDD.n2247 VDD.n1920 72.8958
R3141 VDD.n2247 VDD.n1921 72.8958
R3142 VDD.n2577 VDD.n125 72.8958
R3143 VDD.n131 VDD.n125 72.8958
R3144 VDD.n2584 VDD.n125 72.8958
R3145 VDD.n2587 VDD.n125 72.8958
R3146 VDD.n2509 VDD.n125 72.8958
R3147 VDD.n2508 VDD.n125 72.8958
R3148 VDD.n2516 VDD.n125 72.8958
R3149 VDD.n1565 VDD.n1564 72.8958
R3150 VDD.n1564 VDD.n724 72.8958
R3151 VDD.n1564 VDD.n725 72.8958
R3152 VDD.n1564 VDD.n726 72.8958
R3153 VDD.n1564 VDD.n727 72.8958
R3154 VDD.n1564 VDD.n728 72.8958
R3155 VDD.n1564 VDD.n729 72.8958
R3156 VDD.n1909 VDD.n433 72.8958
R3157 VDD.n1909 VDD.n434 72.8958
R3158 VDD.n1909 VDD.n435 72.8958
R3159 VDD.n1909 VDD.n436 72.8958
R3160 VDD.n1909 VDD.n437 72.8958
R3161 VDD.n1909 VDD.n438 72.8958
R3162 VDD.n1909 VDD.n439 72.8958
R3163 VDD.n2247 VDD.n2246 72.8958
R3164 VDD.n2247 VDD.n1910 72.8958
R3165 VDD.n2247 VDD.n1911 72.8958
R3166 VDD.n2247 VDD.n1912 72.8958
R3167 VDD.n2247 VDD.n1913 72.8958
R3168 VDD.n2247 VDD.n1914 72.8958
R3169 VDD.n2247 VDD.n1915 72.8958
R3170 VDD.n2542 VDD.n125 72.8958
R3171 VDD.n154 VDD.n125 72.8958
R3172 VDD.n2549 VDD.n125 72.8958
R3173 VDD.n149 VDD.n125 72.8958
R3174 VDD.n2557 VDD.n125 72.8958
R3175 VDD.n146 VDD.n125 72.8958
R3176 VDD.n2564 VDD.n125 72.8958
R3177 VDD.n1909 VDD.n431 72.8958
R3178 VDD.n1909 VDD.n430 72.8958
R3179 VDD.n1909 VDD.n429 72.8958
R3180 VDD.n1909 VDD.n428 72.8958
R3181 VDD.n1909 VDD.n427 72.8958
R3182 VDD.n1909 VDD.n426 72.8958
R3183 VDD.n1909 VDD.n425 72.8958
R3184 VDD.n1564 VDD.n730 72.8958
R3185 VDD.n1564 VDD.n731 72.8958
R3186 VDD.n1564 VDD.n732 72.8958
R3187 VDD.n1564 VDD.n733 72.8958
R3188 VDD.n1564 VDD.n734 72.8958
R3189 VDD.n1564 VDD.n735 72.8958
R3190 VDD.n1564 VDD.n736 72.8958
R3191 VDD.n1053 VDD.n1052 67.4914
R3192 VDD.n1070 VDD.n1069 67.4914
R3193 VDD.n1087 VDD.n1086 67.4914
R3194 VDD.n1339 VDD.n1338 67.4914
R3195 VDD.n777 VDD.n776 67.4914
R3196 VDD.n751 VDD.n750 67.4914
R3197 VDD.n2863 VDD.n2862 67.4914
R3198 VDD.n2823 VDD.n2822 67.4914
R3199 VDD.n2806 VDD.n2805 67.4914
R3200 VDD.n116 VDD.n115 67.4914
R3201 VDD.n2656 VDD.n2655 67.4914
R3202 VDD.n65 VDD.n64 67.4914
R3203 VDD.n1102 VDD.n1049 66.2847
R3204 VDD.n1105 VDD.n1049 66.2847
R3205 VDD.n1113 VDD.n1049 66.2847
R3206 VDD.n1115 VDD.n1049 66.2847
R3207 VDD.n1123 VDD.n1049 66.2847
R3208 VDD.n1125 VDD.n1049 66.2847
R3209 VDD.n1133 VDD.n1049 66.2847
R3210 VDD.n1135 VDD.n1049 66.2847
R3211 VDD.n1143 VDD.n1049 66.2847
R3212 VDD.n1145 VDD.n1049 66.2847
R3213 VDD.n1154 VDD.n1049 66.2847
R3214 VDD.n1157 VDD.n1049 66.2847
R3215 VDD.n1074 VDD.n1049 66.2847
R3216 VDD.n1166 VDD.n1049 66.2847
R3217 VDD.n1168 VDD.n1049 66.2847
R3218 VDD.n1176 VDD.n1049 66.2847
R3219 VDD.n1178 VDD.n1049 66.2847
R3220 VDD.n1186 VDD.n1049 66.2847
R3221 VDD.n1188 VDD.n1049 66.2847
R3222 VDD.n1197 VDD.n1049 66.2847
R3223 VDD.n1199 VDD.n1049 66.2847
R3224 VDD.n968 VDD.n745 66.2847
R3225 VDD.n965 VDD.n745 66.2847
R3226 VDD.n960 VDD.n745 66.2847
R3227 VDD.n957 VDD.n745 66.2847
R3228 VDD.n953 VDD.n745 66.2847
R3229 VDD.n1354 VDD.n745 66.2847
R3230 VDD.n786 VDD.n745 66.2847
R3231 VDD.n1361 VDD.n745 66.2847
R3232 VDD.n779 VDD.n745 66.2847
R3233 VDD.n1368 VDD.n745 66.2847
R3234 VDD.n770 VDD.n745 66.2847
R3235 VDD.n1375 VDD.n745 66.2847
R3236 VDD.n763 VDD.n745 66.2847
R3237 VDD.n1382 VDD.n745 66.2847
R3238 VDD.n757 VDD.n745 66.2847
R3239 VDD.n752 VDD.n745 66.2847
R3240 VDD.n1393 VDD.n745 66.2847
R3241 VDD.n1397 VDD.n745 66.2847
R3242 VDD.n745 VDD.n744 66.2847
R3243 VDD.n1323 VDD.n745 66.2847
R3244 VDD.n1326 VDD.n745 66.2847
R3245 VDD.n2681 VDD.n2680 66.2847
R3246 VDD.n2681 VDD.n68 66.2847
R3247 VDD.n2681 VDD.n69 66.2847
R3248 VDD.n2681 VDD.n70 66.2847
R3249 VDD.n2681 VDD.n71 66.2847
R3250 VDD.n2681 VDD.n72 66.2847
R3251 VDD.n2681 VDD.n73 66.2847
R3252 VDD.n2681 VDD.n74 66.2847
R3253 VDD.n2681 VDD.n75 66.2847
R3254 VDD.n2681 VDD.n76 66.2847
R3255 VDD.n2681 VDD.n77 66.2847
R3256 VDD.n2681 VDD.n78 66.2847
R3257 VDD.n2681 VDD.n79 66.2847
R3258 VDD.n2681 VDD.n80 66.2847
R3259 VDD.n2681 VDD.n81 66.2847
R3260 VDD.n2681 VDD.n82 66.2847
R3261 VDD.n2681 VDD.n83 66.2847
R3262 VDD.n2681 VDD.n84 66.2847
R3263 VDD.n2681 VDD.n85 66.2847
R3264 VDD.n2681 VDD.n86 66.2847
R3265 VDD.n2682 VDD.n2681 66.2847
R3266 VDD.n2952 VDD.n2771 66.2847
R3267 VDD.n2952 VDD.n2772 66.2847
R3268 VDD.n2952 VDD.n2773 66.2847
R3269 VDD.n2952 VDD.n2774 66.2847
R3270 VDD.n2952 VDD.n2775 66.2847
R3271 VDD.n2952 VDD.n2776 66.2847
R3272 VDD.n2952 VDD.n2777 66.2847
R3273 VDD.n2952 VDD.n2778 66.2847
R3274 VDD.n2952 VDD.n2779 66.2847
R3275 VDD.n2952 VDD.n2780 66.2847
R3276 VDD.n2952 VDD.n2781 66.2847
R3277 VDD.n2952 VDD.n2782 66.2847
R3278 VDD.n2952 VDD.n2783 66.2847
R3279 VDD.n2952 VDD.n2784 66.2847
R3280 VDD.n2952 VDD.n2785 66.2847
R3281 VDD.n2952 VDD.n2786 66.2847
R3282 VDD.n2952 VDD.n2787 66.2847
R3283 VDD.n2952 VDD.n2788 66.2847
R3284 VDD.n2952 VDD.n2789 66.2847
R3285 VDD.n2952 VDD.n2790 66.2847
R3286 VDD.n2952 VDD.n2791 66.2847
R3287 VDD.n2943 VDD.n2791 52.4337
R3288 VDD.n2941 VDD.n2790 52.4337
R3289 VDD.n2937 VDD.n2789 52.4337
R3290 VDD.n2933 VDD.n2788 52.4337
R3291 VDD.n2929 VDD.n2787 52.4337
R3292 VDD.n2808 VDD.n2786 52.4337
R3293 VDD.n2921 VDD.n2785 52.4337
R3294 VDD.n2917 VDD.n2784 52.4337
R3295 VDD.n2913 VDD.n2783 52.4337
R3296 VDD.n2909 VDD.n2782 52.4337
R3297 VDD.n2905 VDD.n2781 52.4337
R3298 VDD.n2901 VDD.n2780 52.4337
R3299 VDD.n2897 VDD.n2779 52.4337
R3300 VDD.n2889 VDD.n2778 52.4337
R3301 VDD.n2887 VDD.n2777 52.4337
R3302 VDD.n2883 VDD.n2776 52.4337
R3303 VDD.n2879 VDD.n2775 52.4337
R3304 VDD.n2875 VDD.n2774 52.4337
R3305 VDD.n2871 VDD.n2773 52.4337
R3306 VDD.n2867 VDD.n2772 52.4337
R3307 VDD.n2860 VDD.n2771 52.4337
R3308 VDD.n2680 VDD.n2679 52.4337
R3309 VDD.n2674 VDD.n68 52.4337
R3310 VDD.n2671 VDD.n69 52.4337
R3311 VDD.n2667 VDD.n70 52.4337
R3312 VDD.n2663 VDD.n71 52.4337
R3313 VDD.n2659 VDD.n72 52.4337
R3314 VDD.n100 VDD.n73 52.4337
R3315 VDD.n2649 VDD.n74 52.4337
R3316 VDD.n2645 VDD.n75 52.4337
R3317 VDD.n2641 VDD.n76 52.4337
R3318 VDD.n2637 VDD.n77 52.4337
R3319 VDD.n2633 VDD.n78 52.4337
R3320 VDD.n2629 VDD.n79 52.4337
R3321 VDD.n2625 VDD.n80 52.4337
R3322 VDD.n2619 VDD.n81 52.4337
R3323 VDD.n2615 VDD.n82 52.4337
R3324 VDD.n2611 VDD.n83 52.4337
R3325 VDD.n2591 VDD.n84 52.4337
R3326 VDD.n2604 VDD.n85 52.4337
R3327 VDD.n2601 VDD.n86 52.4337
R3328 VDD.n2682 VDD.n67 52.4337
R3329 VDD.n1326 VDD.n1325 52.4337
R3330 VDD.n1323 VDD.n1322 52.4337
R3331 VDD.n1399 VDD.n744 52.4337
R3332 VDD.n1397 VDD.n1396 52.4337
R3333 VDD.n1393 VDD.n1392 52.4337
R3334 VDD.n753 VDD.n752 52.4337
R3335 VDD.n1384 VDD.n757 52.4337
R3336 VDD.n1382 VDD.n1381 52.4337
R3337 VDD.n1377 VDD.n763 52.4337
R3338 VDD.n1375 VDD.n1374 52.4337
R3339 VDD.n1370 VDD.n770 52.4337
R3340 VDD.n1368 VDD.n1367 52.4337
R3341 VDD.n1363 VDD.n779 52.4337
R3342 VDD.n1361 VDD.n1360 52.4337
R3343 VDD.n1356 VDD.n786 52.4337
R3344 VDD.n1354 VDD.n1353 52.4337
R3345 VDD.n954 VDD.n953 52.4337
R3346 VDD.n958 VDD.n957 52.4337
R3347 VDD.n961 VDD.n960 52.4337
R3348 VDD.n966 VDD.n965 52.4337
R3349 VDD.n1336 VDD.n968 52.4337
R3350 VDD.n1102 VDD.n1048 52.4337
R3351 VDD.n1106 VDD.n1105 52.4337
R3352 VDD.n1113 VDD.n1112 52.4337
R3353 VDD.n1116 VDD.n1115 52.4337
R3354 VDD.n1123 VDD.n1122 52.4337
R3355 VDD.n1126 VDD.n1125 52.4337
R3356 VDD.n1133 VDD.n1132 52.4337
R3357 VDD.n1136 VDD.n1135 52.4337
R3358 VDD.n1143 VDD.n1142 52.4337
R3359 VDD.n1146 VDD.n1145 52.4337
R3360 VDD.n1154 VDD.n1153 52.4337
R3361 VDD.n1157 VDD.n1156 52.4337
R3362 VDD.n1075 VDD.n1074 52.4337
R3363 VDD.n1166 VDD.n1165 52.4337
R3364 VDD.n1169 VDD.n1168 52.4337
R3365 VDD.n1176 VDD.n1175 52.4337
R3366 VDD.n1179 VDD.n1178 52.4337
R3367 VDD.n1186 VDD.n1185 52.4337
R3368 VDD.n1189 VDD.n1188 52.4337
R3369 VDD.n1197 VDD.n1196 52.4337
R3370 VDD.n1200 VDD.n1199 52.4337
R3371 VDD.n1103 VDD.n1102 52.4337
R3372 VDD.n1105 VDD.n1095 52.4337
R3373 VDD.n1114 VDD.n1113 52.4337
R3374 VDD.n1115 VDD.n1091 52.4337
R3375 VDD.n1124 VDD.n1123 52.4337
R3376 VDD.n1125 VDD.n1085 52.4337
R3377 VDD.n1134 VDD.n1133 52.4337
R3378 VDD.n1135 VDD.n1081 52.4337
R3379 VDD.n1144 VDD.n1143 52.4337
R3380 VDD.n1145 VDD.n1077 52.4337
R3381 VDD.n1155 VDD.n1154 52.4337
R3382 VDD.n1158 VDD.n1157 52.4337
R3383 VDD.n1074 VDD.n1067 52.4337
R3384 VDD.n1167 VDD.n1166 52.4337
R3385 VDD.n1168 VDD.n1063 52.4337
R3386 VDD.n1177 VDD.n1176 52.4337
R3387 VDD.n1178 VDD.n1059 52.4337
R3388 VDD.n1187 VDD.n1186 52.4337
R3389 VDD.n1188 VDD.n1055 52.4337
R3390 VDD.n1198 VDD.n1197 52.4337
R3391 VDD.n1199 VDD.n1050 52.4337
R3392 VDD.n968 VDD.n967 52.4337
R3393 VDD.n965 VDD.n962 52.4337
R3394 VDD.n960 VDD.n959 52.4337
R3395 VDD.n957 VDD.n956 52.4337
R3396 VDD.n953 VDD.n787 52.4337
R3397 VDD.n1355 VDD.n1354 52.4337
R3398 VDD.n786 VDD.n780 52.4337
R3399 VDD.n1362 VDD.n1361 52.4337
R3400 VDD.n779 VDD.n771 52.4337
R3401 VDD.n1369 VDD.n1368 52.4337
R3402 VDD.n770 VDD.n764 52.4337
R3403 VDD.n1376 VDD.n1375 52.4337
R3404 VDD.n763 VDD.n758 52.4337
R3405 VDD.n1383 VDD.n1382 52.4337
R3406 VDD.n757 VDD.n756 52.4337
R3407 VDD.n752 VDD.n747 52.4337
R3408 VDD.n1394 VDD.n1393 52.4337
R3409 VDD.n1398 VDD.n1397 52.4337
R3410 VDD.n1317 VDD.n744 52.4337
R3411 VDD.n1324 VDD.n1323 52.4337
R3412 VDD.n1327 VDD.n1326 52.4337
R3413 VDD.n2680 VDD.n88 52.4337
R3414 VDD.n2672 VDD.n68 52.4337
R3415 VDD.n2668 VDD.n69 52.4337
R3416 VDD.n2664 VDD.n70 52.4337
R3417 VDD.n2660 VDD.n71 52.4337
R3418 VDD.n101 VDD.n72 52.4337
R3419 VDD.n2650 VDD.n73 52.4337
R3420 VDD.n2646 VDD.n74 52.4337
R3421 VDD.n2642 VDD.n75 52.4337
R3422 VDD.n2638 VDD.n76 52.4337
R3423 VDD.n2634 VDD.n77 52.4337
R3424 VDD.n2630 VDD.n78 52.4337
R3425 VDD.n2626 VDD.n79 52.4337
R3426 VDD.n2618 VDD.n80 52.4337
R3427 VDD.n2616 VDD.n81 52.4337
R3428 VDD.n2612 VDD.n82 52.4337
R3429 VDD.n2590 VDD.n83 52.4337
R3430 VDD.n2593 VDD.n84 52.4337
R3431 VDD.n2602 VDD.n85 52.4337
R3432 VDD.n2598 VDD.n86 52.4337
R3433 VDD.n2683 VDD.n2682 52.4337
R3434 VDD.n2866 VDD.n2771 52.4337
R3435 VDD.n2870 VDD.n2772 52.4337
R3436 VDD.n2874 VDD.n2773 52.4337
R3437 VDD.n2878 VDD.n2774 52.4337
R3438 VDD.n2882 VDD.n2775 52.4337
R3439 VDD.n2886 VDD.n2776 52.4337
R3440 VDD.n2890 VDD.n2777 52.4337
R3441 VDD.n2896 VDD.n2778 52.4337
R3442 VDD.n2900 VDD.n2779 52.4337
R3443 VDD.n2904 VDD.n2780 52.4337
R3444 VDD.n2908 VDD.n2781 52.4337
R3445 VDD.n2912 VDD.n2782 52.4337
R3446 VDD.n2916 VDD.n2783 52.4337
R3447 VDD.n2920 VDD.n2784 52.4337
R3448 VDD.n2807 VDD.n2785 52.4337
R3449 VDD.n2928 VDD.n2786 52.4337
R3450 VDD.n2932 VDD.n2787 52.4337
R3451 VDD.n2936 VDD.n2788 52.4337
R3452 VDD.n2940 VDD.n2789 52.4337
R3453 VDD.n2944 VDD.n2790 52.4337
R3454 VDD.n2792 VDD.n2791 52.4337
R3455 VDD.n1564 VDD.t102 50.3911
R3456 VDD.n125 VDD.t78 50.3911
R3457 VDD.n2564 VDD.n2563 39.2114
R3458 VDD.n2559 VDD.n146 39.2114
R3459 VDD.n2557 VDD.n2556 39.2114
R3460 VDD.n2551 VDD.n149 39.2114
R3461 VDD.n2549 VDD.n2548 39.2114
R3462 VDD.n2544 VDD.n154 39.2114
R3463 VDD.n2542 VDD.n2541 39.2114
R3464 VDD.n2246 VDD.n2245 39.2114
R3465 VDD.n2240 VDD.n1910 39.2114
R3466 VDD.n2237 VDD.n1911 39.2114
R3467 VDD.n2233 VDD.n1912 39.2114
R3468 VDD.n2229 VDD.n1913 39.2114
R3469 VDD.n2225 VDD.n1914 39.2114
R3470 VDD.n2221 VDD.n1915 39.2114
R3471 VDD.n1904 VDD.n439 39.2114
R3472 VDD.n1900 VDD.n438 39.2114
R3473 VDD.n1896 VDD.n437 39.2114
R3474 VDD.n1892 VDD.n436 39.2114
R3475 VDD.n1888 VDD.n435 39.2114
R3476 VDD.n1884 VDD.n434 39.2114
R3477 VDD.n1880 VDD.n433 39.2114
R3478 VDD.n1566 VDD.n1565 39.2114
R3479 VDD.n738 VDD.n724 39.2114
R3480 VDD.n1558 VDD.n725 39.2114
R3481 VDD.n1554 VDD.n726 39.2114
R3482 VDD.n1550 VDD.n727 39.2114
R3483 VDD.n1546 VDD.n728 39.2114
R3484 VDD.n1542 VDD.n729 39.2114
R3485 VDD.n2516 VDD.n2515 39.2114
R3486 VDD.n2511 VDD.n2508 39.2114
R3487 VDD.n2509 VDD.n124 39.2114
R3488 VDD.n2587 VDD.n2586 39.2114
R3489 VDD.n2584 VDD.n2583 39.2114
R3490 VDD.n2579 VDD.n131 39.2114
R3491 VDD.n2577 VDD.n2576 39.2114
R3492 VDD.n2249 VDD.n2248 39.2114
R3493 VDD.n1926 VDD.n1916 39.2114
R3494 VDD.n1930 VDD.n1917 39.2114
R3495 VDD.n1934 VDD.n1918 39.2114
R3496 VDD.n1938 VDD.n1919 39.2114
R3497 VDD.n1942 VDD.n1920 39.2114
R3498 VDD.n1946 VDD.n1921 39.2114
R3499 VDD.n2248 VDD.n423 39.2114
R3500 VDD.n1929 VDD.n1916 39.2114
R3501 VDD.n1933 VDD.n1917 39.2114
R3502 VDD.n1937 VDD.n1918 39.2114
R3503 VDD.n1941 VDD.n1919 39.2114
R3504 VDD.n1945 VDD.n1920 39.2114
R3505 VDD.n1922 VDD.n1921 39.2114
R3506 VDD.n2578 VDD.n2577 39.2114
R3507 VDD.n131 VDD.n127 39.2114
R3508 VDD.n2585 VDD.n2584 39.2114
R3509 VDD.n2588 VDD.n2587 39.2114
R3510 VDD.n2510 VDD.n2509 39.2114
R3511 VDD.n2508 VDD.n2506 39.2114
R3512 VDD.n2517 VDD.n2516 39.2114
R3513 VDD.n1565 VDD.n723 39.2114
R3514 VDD.n1559 VDD.n724 39.2114
R3515 VDD.n1555 VDD.n725 39.2114
R3516 VDD.n1551 VDD.n726 39.2114
R3517 VDD.n1547 VDD.n727 39.2114
R3518 VDD.n1543 VDD.n728 39.2114
R3519 VDD.n1539 VDD.n729 39.2114
R3520 VDD.n1883 VDD.n433 39.2114
R3521 VDD.n1887 VDD.n434 39.2114
R3522 VDD.n1891 VDD.n435 39.2114
R3523 VDD.n1895 VDD.n436 39.2114
R3524 VDD.n1899 VDD.n437 39.2114
R3525 VDD.n1903 VDD.n438 39.2114
R3526 VDD.n441 VDD.n439 39.2114
R3527 VDD.n2246 VDD.n2084 39.2114
R3528 VDD.n2238 VDD.n1910 39.2114
R3529 VDD.n2234 VDD.n1911 39.2114
R3530 VDD.n2230 VDD.n1912 39.2114
R3531 VDD.n2226 VDD.n1913 39.2114
R3532 VDD.n2222 VDD.n1914 39.2114
R3533 VDD.n2218 VDD.n1915 39.2114
R3534 VDD.n2543 VDD.n2542 39.2114
R3535 VDD.n154 VDD.n150 39.2114
R3536 VDD.n2550 VDD.n2549 39.2114
R3537 VDD.n149 VDD.n147 39.2114
R3538 VDD.n2558 VDD.n2557 39.2114
R3539 VDD.n146 VDD.n144 39.2114
R3540 VDD.n2565 VDD.n2564 39.2114
R3541 VDD.n1864 VDD.n425 39.2114
R3542 VDD.n1860 VDD.n426 39.2114
R3543 VDD.n1856 VDD.n427 39.2114
R3544 VDD.n1852 VDD.n428 39.2114
R3545 VDD.n1848 VDD.n429 39.2114
R3546 VDD.n1844 VDD.n430 39.2114
R3547 VDD.n1840 VDD.n431 39.2114
R3548 VDD.n791 VDD.n730 39.2114
R3549 VDD.n795 VDD.n731 39.2114
R3550 VDD.n799 VDD.n732 39.2114
R3551 VDD.n803 VDD.n733 39.2114
R3552 VDD.n947 VDD.n734 39.2114
R3553 VDD.n944 VDD.n735 39.2114
R3554 VDD.n940 VDD.n736 39.2114
R3555 VDD.n1836 VDD.n431 39.2114
R3556 VDD.n1841 VDD.n430 39.2114
R3557 VDD.n1845 VDD.n429 39.2114
R3558 VDD.n1849 VDD.n428 39.2114
R3559 VDD.n1853 VDD.n427 39.2114
R3560 VDD.n1857 VDD.n426 39.2114
R3561 VDD.n1861 VDD.n425 39.2114
R3562 VDD.n794 VDD.n730 39.2114
R3563 VDD.n798 VDD.n731 39.2114
R3564 VDD.n802 VDD.n732 39.2114
R3565 VDD.n805 VDD.n733 39.2114
R3566 VDD.n945 VDD.n734 39.2114
R3567 VDD.n941 VDD.n735 39.2114
R3568 VDD.n936 VDD.n736 39.2114
R3569 VDD.n1202 VDD.n1053 37.2369
R3570 VDD.n1164 VDD.n1070 37.2369
R3571 VDD.n1088 VDD.n1087 37.2369
R3572 VDD.n1340 VDD.n1339 37.2369
R3573 VDD.n778 VDD.n777 37.2369
R3574 VDD.n1389 VDD.n751 37.2369
R3575 VDD.n2864 VDD.n2863 37.2369
R3576 VDD.n2895 VDD.n2823 37.2369
R3577 VDD.n2926 VDD.n2806 37.2369
R3578 VDD.n2624 VDD.n116 37.2369
R3579 VDD.n2657 VDD.n2656 37.2369
R3580 VDD.n66 VDD.n65 37.2369
R3581 VDD.n1907 VDD.n442 30.9078
R3582 VDD.n1881 VDD.n446 30.9078
R3583 VDD.n1540 VDD.n1537 30.9078
R3584 VDD.n1568 VDD.n1567 30.9078
R3585 VDD.n2219 VDD.n2216 30.9078
R3586 VDD.n2540 VDD.n2539 30.9078
R3587 VDD.n2244 VDD.n416 30.9078
R3588 VDD.n2568 VDD.n2567 30.9078
R3589 VDD.n2520 VDD.n2504 30.9078
R3590 VDD.n2575 VDD.n2574 30.9078
R3591 VDD.n2081 VDD.n2080 30.9078
R3592 VDD.n2251 VDD.n2250 30.9078
R3593 VDD.n792 VDD.n716 30.9078
R3594 VDD.n1866 VDD.n1863 30.9078
R3595 VDD.n1835 VDD.n1834 30.9078
R3596 VDD.n935 VDD.n934 30.9078
R3597 VDD.n938 VDD.n807 30.449
R3598 VDD.n1838 VDD.n462 30.449
R3599 VDD.n1405 VDD.n1404 30.449
R3600 VDD.n445 VDD.n444 30.449
R3601 VDD.n1948 VDD.n1925 30.449
R3602 VDD.n153 VDD.n152 30.449
R3603 VDD.n2087 VDD.n2086 30.449
R3604 VDD.n130 VDD.n129 30.449
R3605 VDD.n1208 VDD.n1049 30.0786
R3606 VDD.n1334 VDD.n745 30.0786
R3607 VDD.n2681 VDD.n60 30.0786
R3608 VDD.n2953 VDD.n2952 30.0786
R3609 VDD.n1564 VDD.n718 23.8286
R3610 VDD.n1909 VDD.n424 23.8286
R3611 VDD.n2247 VDD.n418 23.8286
R3612 VDD.n138 VDD.n125 23.8286
R3613 VDD.n1208 VDD.n1043 19.5317
R3614 VDD.n1216 VDD.n1043 19.5317
R3615 VDD.n1216 VDD.n1044 19.5317
R3616 VDD.n1224 VDD.n1032 19.5317
R3617 VDD.n1232 VDD.n1032 19.5317
R3618 VDD.n1232 VDD.n1026 19.5317
R3619 VDD.n1240 VDD.n1026 19.5317
R3620 VDD.n1240 VDD.n1020 19.5317
R3621 VDD.n1248 VDD.n1020 19.5317
R3622 VDD.n1248 VDD.n1014 19.5317
R3623 VDD.n1256 VDD.n1014 19.5317
R3624 VDD.n1256 VDD.t72 19.5317
R3625 VDD.n1267 VDD.t72 19.5317
R3626 VDD.n1267 VDD.n1003 19.5317
R3627 VDD.n1275 VDD.n1003 19.5317
R3628 VDD.n1275 VDD.n997 19.5317
R3629 VDD.n1283 VDD.n997 19.5317
R3630 VDD.n1283 VDD.n991 19.5317
R3631 VDD.n1291 VDD.n991 19.5317
R3632 VDD.n1291 VDD.n985 19.5317
R3633 VDD.n1299 VDD.n985 19.5317
R3634 VDD.n1309 VDD.n978 19.5317
R3635 VDD.n1309 VDD.n971 19.5317
R3636 VDD.n1334 VDD.n971 19.5317
R3637 VDD.n2690 VDD.n60 19.5317
R3638 VDD.n2690 VDD.n54 19.5317
R3639 VDD.n2698 VDD.n54 19.5317
R3640 VDD.n2706 VDD.n48 19.5317
R3641 VDD.n2706 VDD.n42 19.5317
R3642 VDD.n2714 VDD.n42 19.5317
R3643 VDD.n2714 VDD.n36 19.5317
R3644 VDD.n2722 VDD.n36 19.5317
R3645 VDD.n2722 VDD.n30 19.5317
R3646 VDD.n2730 VDD.n30 19.5317
R3647 VDD.n2730 VDD.n22 19.5317
R3648 VDD.t0 VDD.n22 19.5317
R3649 VDD.t0 VDD.n23 19.5317
R3650 VDD.n2976 VDD.n23 19.5317
R3651 VDD.n2976 VDD.n2740 19.5317
R3652 VDD.n2970 VDD.n2740 19.5317
R3653 VDD.n2970 VDD.n2969 19.5317
R3654 VDD.n2969 VDD.n2968 19.5317
R3655 VDD.n2968 VDD.n2750 19.5317
R3656 VDD.n2962 VDD.n2750 19.5317
R3657 VDD.n2962 VDD.n2961 19.5317
R3658 VDD.n2960 VDD.n2761 19.5317
R3659 VDD.n2954 VDD.n2761 19.5317
R3660 VDD.n2954 VDD.n2953 19.5317
R3661 VDD.n1206 VDD.n1041 19.3944
R3662 VDD.n1218 VDD.n1041 19.3944
R3663 VDD.n1218 VDD.n1039 19.3944
R3664 VDD.n1222 VDD.n1039 19.3944
R3665 VDD.n1222 VDD.n1030 19.3944
R3666 VDD.n1234 VDD.n1030 19.3944
R3667 VDD.n1234 VDD.n1028 19.3944
R3668 VDD.n1238 VDD.n1028 19.3944
R3669 VDD.n1238 VDD.n1018 19.3944
R3670 VDD.n1250 VDD.n1018 19.3944
R3671 VDD.n1250 VDD.n1016 19.3944
R3672 VDD.n1254 VDD.n1016 19.3944
R3673 VDD.n1254 VDD.n1007 19.3944
R3674 VDD.n1269 VDD.n1007 19.3944
R3675 VDD.n1269 VDD.n1005 19.3944
R3676 VDD.n1273 VDD.n1005 19.3944
R3677 VDD.n1273 VDD.n995 19.3944
R3678 VDD.n1285 VDD.n995 19.3944
R3679 VDD.n1285 VDD.n993 19.3944
R3680 VDD.n1289 VDD.n993 19.3944
R3681 VDD.n1289 VDD.n983 19.3944
R3682 VDD.n1301 VDD.n983 19.3944
R3683 VDD.n1301 VDD.n980 19.3944
R3684 VDD.n1307 VDD.n980 19.3944
R3685 VDD.n1307 VDD.n981 19.3944
R3686 VDD.n981 VDD.n970 19.3944
R3687 VDD.n1170 VDD.n1066 19.3944
R3688 VDD.n1170 VDD.n1064 19.3944
R3689 VDD.n1174 VDD.n1064 19.3944
R3690 VDD.n1174 VDD.n1062 19.3944
R3691 VDD.n1180 VDD.n1062 19.3944
R3692 VDD.n1180 VDD.n1060 19.3944
R3693 VDD.n1184 VDD.n1060 19.3944
R3694 VDD.n1184 VDD.n1058 19.3944
R3695 VDD.n1190 VDD.n1058 19.3944
R3696 VDD.n1190 VDD.n1056 19.3944
R3697 VDD.n1195 VDD.n1056 19.3944
R3698 VDD.n1195 VDD.n1054 19.3944
R3699 VDD.n1201 VDD.n1054 19.3944
R3700 VDD.n1131 VDD.n1084 19.3944
R3701 VDD.n1137 VDD.n1084 19.3944
R3702 VDD.n1137 VDD.n1082 19.3944
R3703 VDD.n1141 VDD.n1082 19.3944
R3704 VDD.n1141 VDD.n1080 19.3944
R3705 VDD.n1147 VDD.n1080 19.3944
R3706 VDD.n1147 VDD.n1078 19.3944
R3707 VDD.n1152 VDD.n1078 19.3944
R3708 VDD.n1152 VDD.n1076 19.3944
R3709 VDD.n1076 VDD.n1073 19.3944
R3710 VDD.n1159 VDD.n1073 19.3944
R3711 VDD.n1159 VDD.n1071 19.3944
R3712 VDD.n1163 VDD.n1071 19.3944
R3713 VDD.n1101 VDD.n1099 19.3944
R3714 VDD.n1101 VDD.n1098 19.3944
R3715 VDD.n1107 VDD.n1098 19.3944
R3716 VDD.n1107 VDD.n1096 19.3944
R3717 VDD.n1111 VDD.n1096 19.3944
R3718 VDD.n1111 VDD.n1094 19.3944
R3719 VDD.n1117 VDD.n1094 19.3944
R3720 VDD.n1117 VDD.n1092 19.3944
R3721 VDD.n1121 VDD.n1092 19.3944
R3722 VDD.n1121 VDD.n1090 19.3944
R3723 VDD.n1127 VDD.n1090 19.3944
R3724 VDD.n1210 VDD.n1046 19.3944
R3725 VDD.n1214 VDD.n1046 19.3944
R3726 VDD.n1214 VDD.n1036 19.3944
R3727 VDD.n1226 VDD.n1036 19.3944
R3728 VDD.n1226 VDD.n1034 19.3944
R3729 VDD.n1230 VDD.n1034 19.3944
R3730 VDD.n1230 VDD.n1024 19.3944
R3731 VDD.n1242 VDD.n1024 19.3944
R3732 VDD.n1242 VDD.n1022 19.3944
R3733 VDD.n1246 VDD.n1022 19.3944
R3734 VDD.n1246 VDD.n1012 19.3944
R3735 VDD.n1258 VDD.n1012 19.3944
R3736 VDD.n1258 VDD.n1010 19.3944
R3737 VDD.n1265 VDD.n1010 19.3944
R3738 VDD.n1265 VDD.n1001 19.3944
R3739 VDD.n1277 VDD.n1001 19.3944
R3740 VDD.n1277 VDD.n999 19.3944
R3741 VDD.n1281 VDD.n999 19.3944
R3742 VDD.n1281 VDD.n989 19.3944
R3743 VDD.n1293 VDD.n989 19.3944
R3744 VDD.n1293 VDD.n987 19.3944
R3745 VDD.n1297 VDD.n987 19.3944
R3746 VDD.n1297 VDD.n976 19.3944
R3747 VDD.n1311 VDD.n976 19.3944
R3748 VDD.n1311 VDD.n974 19.3944
R3749 VDD.n1332 VDD.n974 19.3944
R3750 VDD.n1359 VDD.n1358 19.3944
R3751 VDD.n1358 VDD.n1357 19.3944
R3752 VDD.n1357 VDD.n785 19.3944
R3753 VDD.n1352 VDD.n785 19.3944
R3754 VDD.n1352 VDD.n1351 19.3944
R3755 VDD.n955 VDD.n790 19.3944
R3756 VDD.n1347 VDD.n952 19.3944
R3757 VDD.n1347 VDD.n1346 19.3944
R3758 VDD.n1346 VDD.n1345 19.3944
R3759 VDD.n1345 VDD.n963 19.3944
R3760 VDD.n1341 VDD.n963 19.3944
R3761 VDD.n1385 VDD.n749 19.3944
R3762 VDD.n1385 VDD.n755 19.3944
R3763 VDD.n1380 VDD.n755 19.3944
R3764 VDD.n1380 VDD.n1379 19.3944
R3765 VDD.n1379 VDD.n1378 19.3944
R3766 VDD.n1378 VDD.n762 19.3944
R3767 VDD.n1373 VDD.n762 19.3944
R3768 VDD.n1373 VDD.n1372 19.3944
R3769 VDD.n1372 VDD.n1371 19.3944
R3770 VDD.n1371 VDD.n769 19.3944
R3771 VDD.n1366 VDD.n769 19.3944
R3772 VDD.n1366 VDD.n1365 19.3944
R3773 VDD.n1365 VDD.n1364 19.3944
R3774 VDD.n1329 VDD.n1328 19.3944
R3775 VDD.n1328 VDD.n1315 19.3944
R3776 VDD.n1316 VDD.n1315 19.3944
R3777 VDD.n1321 VDD.n1316 19.3944
R3778 VDD.n1321 VDD.n743 19.3944
R3779 VDD.n1400 VDD.n743 19.3944
R3780 VDD.n1395 VDD.n742 19.3944
R3781 VDD.n1391 VDD.n746 19.3944
R3782 VDD.n1391 VDD.n1390 19.3944
R3783 VDD.n2688 VDD.n62 19.3944
R3784 VDD.n2688 VDD.n52 19.3944
R3785 VDD.n2700 VDD.n52 19.3944
R3786 VDD.n2700 VDD.n50 19.3944
R3787 VDD.n2704 VDD.n50 19.3944
R3788 VDD.n2704 VDD.n40 19.3944
R3789 VDD.n2716 VDD.n40 19.3944
R3790 VDD.n2716 VDD.n38 19.3944
R3791 VDD.n2720 VDD.n38 19.3944
R3792 VDD.n2720 VDD.n28 19.3944
R3793 VDD.n2732 VDD.n28 19.3944
R3794 VDD.n2732 VDD.n26 19.3944
R3795 VDD.n2980 VDD.n26 19.3944
R3796 VDD.n2980 VDD.n2979 19.3944
R3797 VDD.n2979 VDD.n2978 19.3944
R3798 VDD.n2978 VDD.n2738 19.3944
R3799 VDD.n2842 VDD.n2738 19.3944
R3800 VDD.n2843 VDD.n2842 19.3944
R3801 VDD.n2843 VDD.n2839 19.3944
R3802 VDD.n2848 VDD.n2839 19.3944
R3803 VDD.n2849 VDD.n2848 19.3944
R3804 VDD.n2850 VDD.n2849 19.3944
R3805 VDD.n2850 VDD.n2837 19.3944
R3806 VDD.n2855 VDD.n2837 19.3944
R3807 VDD.n2856 VDD.n2855 19.3944
R3808 VDD.n2857 VDD.n2856 19.3944
R3809 VDD.n2891 VDD.n2821 19.3944
R3810 VDD.n2891 VDD.n2888 19.3944
R3811 VDD.n2888 VDD.n2885 19.3944
R3812 VDD.n2885 VDD.n2884 19.3944
R3813 VDD.n2884 VDD.n2881 19.3944
R3814 VDD.n2881 VDD.n2880 19.3944
R3815 VDD.n2880 VDD.n2877 19.3944
R3816 VDD.n2877 VDD.n2876 19.3944
R3817 VDD.n2876 VDD.n2873 19.3944
R3818 VDD.n2873 VDD.n2872 19.3944
R3819 VDD.n2872 VDD.n2869 19.3944
R3820 VDD.n2869 VDD.n2868 19.3944
R3821 VDD.n2868 VDD.n2865 19.3944
R3822 VDD.n2922 VDD.n2804 19.3944
R3823 VDD.n2922 VDD.n2919 19.3944
R3824 VDD.n2919 VDD.n2918 19.3944
R3825 VDD.n2918 VDD.n2915 19.3944
R3826 VDD.n2915 VDD.n2914 19.3944
R3827 VDD.n2914 VDD.n2911 19.3944
R3828 VDD.n2911 VDD.n2910 19.3944
R3829 VDD.n2910 VDD.n2907 19.3944
R3830 VDD.n2907 VDD.n2906 19.3944
R3831 VDD.n2906 VDD.n2903 19.3944
R3832 VDD.n2903 VDD.n2902 19.3944
R3833 VDD.n2902 VDD.n2899 19.3944
R3834 VDD.n2899 VDD.n2898 19.3944
R3835 VDD.n2950 VDD.n2949 19.3944
R3836 VDD.n2949 VDD.n2795 19.3944
R3837 VDD.n2945 VDD.n2795 19.3944
R3838 VDD.n2945 VDD.n2942 19.3944
R3839 VDD.n2942 VDD.n2939 19.3944
R3840 VDD.n2939 VDD.n2938 19.3944
R3841 VDD.n2938 VDD.n2935 19.3944
R3842 VDD.n2935 VDD.n2934 19.3944
R3843 VDD.n2934 VDD.n2931 19.3944
R3844 VDD.n2931 VDD.n2930 19.3944
R3845 VDD.n2930 VDD.n2927 19.3944
R3846 VDD.n2692 VDD.n58 19.3944
R3847 VDD.n2692 VDD.n56 19.3944
R3848 VDD.n2696 VDD.n56 19.3944
R3849 VDD.n2696 VDD.n46 19.3944
R3850 VDD.n2708 VDD.n46 19.3944
R3851 VDD.n2708 VDD.n44 19.3944
R3852 VDD.n2712 VDD.n44 19.3944
R3853 VDD.n2712 VDD.n34 19.3944
R3854 VDD.n2724 VDD.n34 19.3944
R3855 VDD.n2724 VDD.n32 19.3944
R3856 VDD.n2728 VDD.n32 19.3944
R3857 VDD.n2728 VDD.n18 19.3944
R3858 VDD.n2983 VDD.n18 19.3944
R3859 VDD.n2983 VDD.n19 19.3944
R3860 VDD.n2974 VDD.n19 19.3944
R3861 VDD.n2974 VDD.n2973 19.3944
R3862 VDD.n2973 VDD.n2972 19.3944
R3863 VDD.n2972 VDD.n2745 19.3944
R3864 VDD.n2966 VDD.n2745 19.3944
R3865 VDD.n2966 VDD.n2965 19.3944
R3866 VDD.n2965 VDD.n2964 19.3944
R3867 VDD.n2964 VDD.n2756 19.3944
R3868 VDD.n2958 VDD.n2756 19.3944
R3869 VDD.n2958 VDD.n2957 19.3944
R3870 VDD.n2957 VDD.n2956 19.3944
R3871 VDD.n2956 VDD.n2767 19.3944
R3872 VDD.n2651 VDD.n99 19.3944
R3873 VDD.n2651 VDD.n2648 19.3944
R3874 VDD.n2648 VDD.n2647 19.3944
R3875 VDD.n2647 VDD.n2644 19.3944
R3876 VDD.n2644 VDD.n2643 19.3944
R3877 VDD.n2643 VDD.n2640 19.3944
R3878 VDD.n2640 VDD.n2639 19.3944
R3879 VDD.n2639 VDD.n2636 19.3944
R3880 VDD.n2636 VDD.n2635 19.3944
R3881 VDD.n2635 VDD.n2632 19.3944
R3882 VDD.n2632 VDD.n2631 19.3944
R3883 VDD.n2631 VDD.n2628 19.3944
R3884 VDD.n2628 VDD.n2627 19.3944
R3885 VDD.n2678 VDD.n2677 19.3944
R3886 VDD.n2677 VDD.n2676 19.3944
R3887 VDD.n2676 VDD.n2675 19.3944
R3888 VDD.n2675 VDD.n2673 19.3944
R3889 VDD.n2673 VDD.n2670 19.3944
R3890 VDD.n2670 VDD.n2669 19.3944
R3891 VDD.n2666 VDD.n2665 19.3944
R3892 VDD.n2662 VDD.n2661 19.3944
R3893 VDD.n2661 VDD.n2658 19.3944
R3894 VDD.n2620 VDD.n114 19.3944
R3895 VDD.n2620 VDD.n2617 19.3944
R3896 VDD.n2617 VDD.n2614 19.3944
R3897 VDD.n2614 VDD.n2613 19.3944
R3898 VDD.n2613 VDD.n2610 19.3944
R3899 VDD.n2592 VDD.n120 19.3944
R3900 VDD.n2606 VDD.n2605 19.3944
R3901 VDD.n2605 VDD.n2603 19.3944
R3902 VDD.n2603 VDD.n2600 19.3944
R3903 VDD.n2600 VDD.n2599 19.3944
R3904 VDD.n2599 VDD.n2597 19.3944
R3905 VDD.n1164 VDD.n1066 19.0066
R3906 VDD.n1359 VDD.n778 19.0066
R3907 VDD.n2895 VDD.n2821 19.0066
R3908 VDD.n2624 VDD.n114 19.0066
R3909 VDD.n1044 VDD.t45 16.7974
R3910 VDD.t16 VDD.n978 16.7974
R3911 VDD.n2698 VDD.t8 16.7974
R3912 VDD.t12 VDD.n2960 16.7974
R3913 VDD.n1571 VDD.n718 13.2817
R3914 VDD.n1571 VDD.n712 13.2817
R3915 VDD.n1577 VDD.n712 13.2817
R3916 VDD.n1577 VDD.n706 13.2817
R3917 VDD.n1583 VDD.n706 13.2817
R3918 VDD.n1583 VDD.n700 13.2817
R3919 VDD.n1589 VDD.n700 13.2817
R3920 VDD.n1595 VDD.n694 13.2817
R3921 VDD.n1595 VDD.n688 13.2817
R3922 VDD.n1601 VDD.n688 13.2817
R3923 VDD.n1601 VDD.n682 13.2817
R3924 VDD.n1607 VDD.n682 13.2817
R3925 VDD.n1607 VDD.n676 13.2817
R3926 VDD.n1613 VDD.n676 13.2817
R3927 VDD.n1613 VDD.n670 13.2817
R3928 VDD.n1619 VDD.n670 13.2817
R3929 VDD.n1619 VDD.n664 13.2817
R3930 VDD.n1625 VDD.n664 13.2817
R3931 VDD.n1625 VDD.n658 13.2817
R3932 VDD.n1631 VDD.n658 13.2817
R3933 VDD.n1637 VDD.n651 13.2817
R3934 VDD.n1637 VDD.n654 13.2817
R3935 VDD.n1643 VDD.n640 13.2817
R3936 VDD.n1649 VDD.n640 13.2817
R3937 VDD.n1649 VDD.n634 13.2817
R3938 VDD.n1655 VDD.n634 13.2817
R3939 VDD.n1655 VDD.n628 13.2817
R3940 VDD.n1661 VDD.n628 13.2817
R3941 VDD.n1661 VDD.n622 13.2817
R3942 VDD.n1667 VDD.n622 13.2817
R3943 VDD.n1667 VDD.n616 13.2817
R3944 VDD.n1673 VDD.n616 13.2817
R3945 VDD.n1673 VDD.n609 13.2817
R3946 VDD.n1679 VDD.n609 13.2817
R3947 VDD.n1679 VDD.n612 13.2817
R3948 VDD.n1685 VDD.n597 13.2817
R3949 VDD.n1691 VDD.n597 13.2817
R3950 VDD.n1691 VDD.n600 13.2817
R3951 VDD.n1697 VDD.n586 13.2817
R3952 VDD.n1703 VDD.n586 13.2817
R3953 VDD.n1703 VDD.n580 13.2817
R3954 VDD.n1709 VDD.n580 13.2817
R3955 VDD.n1709 VDD.n574 13.2817
R3956 VDD.n1715 VDD.n574 13.2817
R3957 VDD.n1715 VDD.n568 13.2817
R3958 VDD.n1721 VDD.n568 13.2817
R3959 VDD.n1727 VDD.n562 13.2817
R3960 VDD.n1727 VDD.n556 13.2817
R3961 VDD.n1733 VDD.n556 13.2817
R3962 VDD.n1739 VDD.n550 13.2817
R3963 VDD.n1739 VDD.n544 13.2817
R3964 VDD.n1745 VDD.n544 13.2817
R3965 VDD.n1745 VDD.n538 13.2817
R3966 VDD.n1751 VDD.n538 13.2817
R3967 VDD.n1751 VDD.n532 13.2817
R3968 VDD.n1757 VDD.n532 13.2817
R3969 VDD.n1757 VDD.n526 13.2817
R3970 VDD.n1763 VDD.n526 13.2817
R3971 VDD.n1769 VDD.n520 13.2817
R3972 VDD.n1769 VDD.n514 13.2817
R3973 VDD.n1775 VDD.n514 13.2817
R3974 VDD.n1781 VDD.n508 13.2817
R3975 VDD.n1781 VDD.n502 13.2817
R3976 VDD.n1787 VDD.n502 13.2817
R3977 VDD.n1787 VDD.n496 13.2817
R3978 VDD.n1793 VDD.n496 13.2817
R3979 VDD.n1793 VDD.n490 13.2817
R3980 VDD.n1799 VDD.n490 13.2817
R3981 VDD.n1799 VDD.n484 13.2817
R3982 VDD.n1805 VDD.n484 13.2817
R3983 VDD.n1805 VDD.n477 13.2817
R3984 VDD.n1811 VDD.n477 13.2817
R3985 VDD.n1811 VDD.n480 13.2817
R3986 VDD.n1819 VDD.n465 13.2817
R3987 VDD.n1825 VDD.n465 13.2817
R3988 VDD.n1825 VDD.n455 13.2817
R3989 VDD.n1871 VDD.n455 13.2817
R3990 VDD.n1871 VDD.n449 13.2817
R3991 VDD.n1877 VDD.n449 13.2817
R3992 VDD.n1877 VDD.n424 13.2817
R3993 VDD.n2254 VDD.n418 13.2817
R3994 VDD.n2254 VDD.n412 13.2817
R3995 VDD.n2260 VDD.n412 13.2817
R3996 VDD.n2260 VDD.n406 13.2817
R3997 VDD.n2266 VDD.n406 13.2817
R3998 VDD.n2266 VDD.n400 13.2817
R3999 VDD.n2272 VDD.n400 13.2817
R4000 VDD.n2278 VDD.n394 13.2817
R4001 VDD.n2278 VDD.n388 13.2817
R4002 VDD.n2284 VDD.n388 13.2817
R4003 VDD.n2284 VDD.n382 13.2817
R4004 VDD.n2290 VDD.n382 13.2817
R4005 VDD.n2290 VDD.n376 13.2817
R4006 VDD.n2296 VDD.n376 13.2817
R4007 VDD.n2296 VDD.n370 13.2817
R4008 VDD.n2302 VDD.n370 13.2817
R4009 VDD.n2302 VDD.n363 13.2817
R4010 VDD.n2308 VDD.n363 13.2817
R4011 VDD.n2308 VDD.n366 13.2817
R4012 VDD.n2314 VDD.n351 13.2817
R4013 VDD.n2320 VDD.n351 13.2817
R4014 VDD.n2320 VDD.n354 13.2817
R4015 VDD.n2326 VDD.n340 13.2817
R4016 VDD.n2332 VDD.n340 13.2817
R4017 VDD.n2332 VDD.n334 13.2817
R4018 VDD.n2338 VDD.n334 13.2817
R4019 VDD.n2338 VDD.n328 13.2817
R4020 VDD.n2344 VDD.n328 13.2817
R4021 VDD.n2344 VDD.n321 13.2817
R4022 VDD.n2350 VDD.n321 13.2817
R4023 VDD.n2350 VDD.n324 13.2817
R4024 VDD.n2356 VDD.n309 13.2817
R4025 VDD.n2362 VDD.n309 13.2817
R4026 VDD.n2362 VDD.n312 13.2817
R4027 VDD.n2368 VDD.n298 13.2817
R4028 VDD.n2374 VDD.n298 13.2817
R4029 VDD.n2374 VDD.n292 13.2817
R4030 VDD.n2380 VDD.n292 13.2817
R4031 VDD.n2380 VDD.n286 13.2817
R4032 VDD.n2386 VDD.n286 13.2817
R4033 VDD.n2386 VDD.n280 13.2817
R4034 VDD.n2392 VDD.n280 13.2817
R4035 VDD.n2398 VDD.n274 13.2817
R4036 VDD.n2398 VDD.n268 13.2817
R4037 VDD.n2404 VDD.n268 13.2817
R4038 VDD.n2410 VDD.n262 13.2817
R4039 VDD.n2410 VDD.n256 13.2817
R4040 VDD.n2416 VDD.n256 13.2817
R4041 VDD.n2416 VDD.n250 13.2817
R4042 VDD.n2422 VDD.n250 13.2817
R4043 VDD.n2422 VDD.n244 13.2817
R4044 VDD.n2428 VDD.n244 13.2817
R4045 VDD.n2428 VDD.n238 13.2817
R4046 VDD.n2434 VDD.n238 13.2817
R4047 VDD.n2434 VDD.n232 13.2817
R4048 VDD.n2440 VDD.n232 13.2817
R4049 VDD.n2440 VDD.n226 13.2817
R4050 VDD.n2446 VDD.n226 13.2817
R4051 VDD.n2452 VDD.n219 13.2817
R4052 VDD.n2452 VDD.n222 13.2817
R4053 VDD.n2458 VDD.n208 13.2817
R4054 VDD.n2464 VDD.n208 13.2817
R4055 VDD.n2464 VDD.n202 13.2817
R4056 VDD.n2470 VDD.n202 13.2817
R4057 VDD.n2470 VDD.n196 13.2817
R4058 VDD.n2476 VDD.n196 13.2817
R4059 VDD.n2476 VDD.n190 13.2817
R4060 VDD.n2482 VDD.n190 13.2817
R4061 VDD.n2482 VDD.n184 13.2817
R4062 VDD.n2488 VDD.n184 13.2817
R4063 VDD.n2488 VDD.n177 13.2817
R4064 VDD.n2494 VDD.n177 13.2817
R4065 VDD.n2494 VDD.n180 13.2817
R4066 VDD.n2500 VDD.n165 13.2817
R4067 VDD.n2528 VDD.n165 13.2817
R4068 VDD.n2528 VDD.n159 13.2817
R4069 VDD.n2534 VDD.n159 13.2817
R4070 VDD.n2534 VDD.n136 13.2817
R4071 VDD.n2571 VDD.n136 13.2817
R4072 VDD.n2571 VDD.n138 13.2817
R4073 VDD.n1131 VDD.n1088 12.9944
R4074 VDD.n1127 VDD.n1088 12.9944
R4075 VDD.n1389 VDD.n749 12.9944
R4076 VDD.n1390 VDD.n1389 12.9944
R4077 VDD.n2926 VDD.n2804 12.9944
R4078 VDD.n2927 VDD.n2926 12.9944
R4079 VDD.n2657 VDD.n99 12.9944
R4080 VDD.n2658 VDD.n2657 12.9944
R4081 VDD.n1697 VDD.t85 12.8911
R4082 VDD.n2392 VDD.t88 12.8911
R4083 VDD.n1589 VDD.t20 11.9146
R4084 VDD.n2500 VDD.t4 11.9146
R4085 VDD.n7 VDD.t79 11.651
R4086 VDD.n7 VDD.t115 11.651
R4087 VDD.n8 VDD.t84 11.651
R4088 VDD.n8 VDD.t105 11.651
R4089 VDD.n10 VDD.t92 11.651
R4090 VDD.n10 VDD.t89 11.651
R4091 VDD.n12 VDD.t111 11.651
R4092 VDD.n12 VDD.t95 11.651
R4093 VDD.n5 VDD.t81 11.651
R4094 VDD.n5 VDD.t109 11.651
R4095 VDD.n3 VDD.t86 11.651
R4096 VDD.n3 VDD.t117 11.651
R4097 VDD.n1 VDD.t107 11.651
R4098 VDD.n1 VDD.t113 11.651
R4099 VDD.n0 VDD.t99 11.651
R4100 VDD.n0 VDD.t103 11.651
R4101 VDD.t80 VDD.n508 11.3286
R4102 VDD.n366 VDD.t94 11.3286
R4103 VDD.n1907 VDD.n1906 10.6151
R4104 VDD.n1906 VDD.n1905 10.6151
R4105 VDD.n1905 VDD.n1902 10.6151
R4106 VDD.n1902 VDD.n1901 10.6151
R4107 VDD.n1901 VDD.n1898 10.6151
R4108 VDD.n1898 VDD.n1897 10.6151
R4109 VDD.n1897 VDD.n1894 10.6151
R4110 VDD.n1894 VDD.n1893 10.6151
R4111 VDD.n1893 VDD.n1890 10.6151
R4112 VDD.n1890 VDD.n1889 10.6151
R4113 VDD.n1889 VDD.n1886 10.6151
R4114 VDD.n1886 VDD.n1885 10.6151
R4115 VDD.n1882 VDD.n1881 10.6151
R4116 VDD.n1537 VDD.n1536 10.6151
R4117 VDD.n1536 VDD.n1535 10.6151
R4118 VDD.n1535 VDD.n1533 10.6151
R4119 VDD.n1533 VDD.n1532 10.6151
R4120 VDD.n1532 VDD.n1530 10.6151
R4121 VDD.n1530 VDD.n1529 10.6151
R4122 VDD.n1529 VDD.n1527 10.6151
R4123 VDD.n1527 VDD.n1526 10.6151
R4124 VDD.n1526 VDD.n1524 10.6151
R4125 VDD.n1524 VDD.n1523 10.6151
R4126 VDD.n1523 VDD.n1521 10.6151
R4127 VDD.n1521 VDD.n1520 10.6151
R4128 VDD.n1520 VDD.n1518 10.6151
R4129 VDD.n1518 VDD.n1517 10.6151
R4130 VDD.n1517 VDD.n1515 10.6151
R4131 VDD.n1515 VDD.n1514 10.6151
R4132 VDD.n1514 VDD.n1512 10.6151
R4133 VDD.n1512 VDD.n1511 10.6151
R4134 VDD.n1511 VDD.n1509 10.6151
R4135 VDD.n1509 VDD.n1508 10.6151
R4136 VDD.n1508 VDD.n1506 10.6151
R4137 VDD.n1506 VDD.n1505 10.6151
R4138 VDD.n1505 VDD.n1503 10.6151
R4139 VDD.n1503 VDD.n1502 10.6151
R4140 VDD.n1502 VDD.n1500 10.6151
R4141 VDD.n1500 VDD.n1499 10.6151
R4142 VDD.n1499 VDD.n1497 10.6151
R4143 VDD.n1497 VDD.n1496 10.6151
R4144 VDD.n1496 VDD.n1494 10.6151
R4145 VDD.n1494 VDD.n1493 10.6151
R4146 VDD.n1493 VDD.n1491 10.6151
R4147 VDD.n1491 VDD.n1490 10.6151
R4148 VDD.n1490 VDD.n1488 10.6151
R4149 VDD.n1488 VDD.n1487 10.6151
R4150 VDD.n1487 VDD.n1485 10.6151
R4151 VDD.n1485 VDD.n1484 10.6151
R4152 VDD.n1484 VDD.n1482 10.6151
R4153 VDD.n1482 VDD.n1481 10.6151
R4154 VDD.n1481 VDD.n1479 10.6151
R4155 VDD.n1479 VDD.n1478 10.6151
R4156 VDD.n1478 VDD.n1476 10.6151
R4157 VDD.n1476 VDD.n1475 10.6151
R4158 VDD.n1475 VDD.n1473 10.6151
R4159 VDD.n1473 VDD.n1472 10.6151
R4160 VDD.n1472 VDD.n1470 10.6151
R4161 VDD.n1470 VDD.n1469 10.6151
R4162 VDD.n1469 VDD.n1467 10.6151
R4163 VDD.n1467 VDD.n1466 10.6151
R4164 VDD.n1466 VDD.n1464 10.6151
R4165 VDD.n1464 VDD.n1463 10.6151
R4166 VDD.n1463 VDD.n1461 10.6151
R4167 VDD.n1461 VDD.n1460 10.6151
R4168 VDD.n1460 VDD.n1458 10.6151
R4169 VDD.n1458 VDD.n1457 10.6151
R4170 VDD.n1457 VDD.n1455 10.6151
R4171 VDD.n1455 VDD.n1454 10.6151
R4172 VDD.n1454 VDD.n1452 10.6151
R4173 VDD.n1452 VDD.n1451 10.6151
R4174 VDD.n1451 VDD.n1449 10.6151
R4175 VDD.n1449 VDD.n1448 10.6151
R4176 VDD.n1448 VDD.n1446 10.6151
R4177 VDD.n1446 VDD.n1445 10.6151
R4178 VDD.n1445 VDD.n1443 10.6151
R4179 VDD.n1443 VDD.n1442 10.6151
R4180 VDD.n1442 VDD.n1440 10.6151
R4181 VDD.n1440 VDD.n1439 10.6151
R4182 VDD.n1439 VDD.n1437 10.6151
R4183 VDD.n1437 VDD.n1436 10.6151
R4184 VDD.n1436 VDD.n1434 10.6151
R4185 VDD.n1434 VDD.n1433 10.6151
R4186 VDD.n1433 VDD.n1431 10.6151
R4187 VDD.n1431 VDD.n1430 10.6151
R4188 VDD.n1430 VDD.n1428 10.6151
R4189 VDD.n1428 VDD.n1427 10.6151
R4190 VDD.n1427 VDD.n1425 10.6151
R4191 VDD.n1425 VDD.n1424 10.6151
R4192 VDD.n1424 VDD.n1422 10.6151
R4193 VDD.n1422 VDD.n1421 10.6151
R4194 VDD.n1421 VDD.n1419 10.6151
R4195 VDD.n1419 VDD.n1418 10.6151
R4196 VDD.n1418 VDD.n1416 10.6151
R4197 VDD.n1416 VDD.n1415 10.6151
R4198 VDD.n1415 VDD.n1413 10.6151
R4199 VDD.n1413 VDD.n1412 10.6151
R4200 VDD.n1412 VDD.n1410 10.6151
R4201 VDD.n1410 VDD.n1409 10.6151
R4202 VDD.n1409 VDD.n1407 10.6151
R4203 VDD.n1407 VDD.n1406 10.6151
R4204 VDD.n1406 VDD.n448 10.6151
R4205 VDD.n448 VDD.n446 10.6151
R4206 VDD.n1567 VDD.n722 10.6151
R4207 VDD.n1562 VDD.n722 10.6151
R4208 VDD.n1562 VDD.n1561 10.6151
R4209 VDD.n1561 VDD.n1560 10.6151
R4210 VDD.n1560 VDD.n1557 10.6151
R4211 VDD.n1557 VDD.n1556 10.6151
R4212 VDD.n1556 VDD.n1553 10.6151
R4213 VDD.n1553 VDD.n1552 10.6151
R4214 VDD.n1552 VDD.n1549 10.6151
R4215 VDD.n1549 VDD.n1548 10.6151
R4216 VDD.n1548 VDD.n1545 10.6151
R4217 VDD.n1545 VDD.n1544 10.6151
R4218 VDD.n1541 VDD.n1540 10.6151
R4219 VDD.n1569 VDD.n1568 10.6151
R4220 VDD.n1569 VDD.n710 10.6151
R4221 VDD.n1579 VDD.n710 10.6151
R4222 VDD.n1580 VDD.n1579 10.6151
R4223 VDD.n1581 VDD.n1580 10.6151
R4224 VDD.n1581 VDD.n698 10.6151
R4225 VDD.n1591 VDD.n698 10.6151
R4226 VDD.n1592 VDD.n1591 10.6151
R4227 VDD.n1593 VDD.n1592 10.6151
R4228 VDD.n1593 VDD.n686 10.6151
R4229 VDD.n1603 VDD.n686 10.6151
R4230 VDD.n1604 VDD.n1603 10.6151
R4231 VDD.n1605 VDD.n1604 10.6151
R4232 VDD.n1605 VDD.n674 10.6151
R4233 VDD.n1615 VDD.n674 10.6151
R4234 VDD.n1616 VDD.n1615 10.6151
R4235 VDD.n1617 VDD.n1616 10.6151
R4236 VDD.n1617 VDD.n662 10.6151
R4237 VDD.n1627 VDD.n662 10.6151
R4238 VDD.n1628 VDD.n1627 10.6151
R4239 VDD.n1629 VDD.n1628 10.6151
R4240 VDD.n1629 VDD.n649 10.6151
R4241 VDD.n1639 VDD.n649 10.6151
R4242 VDD.n1640 VDD.n1639 10.6151
R4243 VDD.n1641 VDD.n1640 10.6151
R4244 VDD.n1641 VDD.n638 10.6151
R4245 VDD.n1651 VDD.n638 10.6151
R4246 VDD.n1652 VDD.n1651 10.6151
R4247 VDD.n1653 VDD.n1652 10.6151
R4248 VDD.n1653 VDD.n626 10.6151
R4249 VDD.n1663 VDD.n626 10.6151
R4250 VDD.n1664 VDD.n1663 10.6151
R4251 VDD.n1665 VDD.n1664 10.6151
R4252 VDD.n1665 VDD.n614 10.6151
R4253 VDD.n1675 VDD.n614 10.6151
R4254 VDD.n1676 VDD.n1675 10.6151
R4255 VDD.n1677 VDD.n1676 10.6151
R4256 VDD.n1677 VDD.n602 10.6151
R4257 VDD.n1687 VDD.n602 10.6151
R4258 VDD.n1688 VDD.n1687 10.6151
R4259 VDD.n1689 VDD.n1688 10.6151
R4260 VDD.n1689 VDD.n590 10.6151
R4261 VDD.n1699 VDD.n590 10.6151
R4262 VDD.n1700 VDD.n1699 10.6151
R4263 VDD.n1701 VDD.n1700 10.6151
R4264 VDD.n1701 VDD.n578 10.6151
R4265 VDD.n1711 VDD.n578 10.6151
R4266 VDD.n1712 VDD.n1711 10.6151
R4267 VDD.n1713 VDD.n1712 10.6151
R4268 VDD.n1713 VDD.n566 10.6151
R4269 VDD.n1723 VDD.n566 10.6151
R4270 VDD.n1724 VDD.n1723 10.6151
R4271 VDD.n1725 VDD.n1724 10.6151
R4272 VDD.n1725 VDD.n554 10.6151
R4273 VDD.n1735 VDD.n554 10.6151
R4274 VDD.n1736 VDD.n1735 10.6151
R4275 VDD.n1737 VDD.n1736 10.6151
R4276 VDD.n1737 VDD.n542 10.6151
R4277 VDD.n1747 VDD.n542 10.6151
R4278 VDD.n1748 VDD.n1747 10.6151
R4279 VDD.n1749 VDD.n1748 10.6151
R4280 VDD.n1749 VDD.n530 10.6151
R4281 VDD.n1759 VDD.n530 10.6151
R4282 VDD.n1760 VDD.n1759 10.6151
R4283 VDD.n1761 VDD.n1760 10.6151
R4284 VDD.n1761 VDD.n518 10.6151
R4285 VDD.n1771 VDD.n518 10.6151
R4286 VDD.n1772 VDD.n1771 10.6151
R4287 VDD.n1773 VDD.n1772 10.6151
R4288 VDD.n1773 VDD.n506 10.6151
R4289 VDD.n1783 VDD.n506 10.6151
R4290 VDD.n1784 VDD.n1783 10.6151
R4291 VDD.n1785 VDD.n1784 10.6151
R4292 VDD.n1785 VDD.n494 10.6151
R4293 VDD.n1795 VDD.n494 10.6151
R4294 VDD.n1796 VDD.n1795 10.6151
R4295 VDD.n1797 VDD.n1796 10.6151
R4296 VDD.n1797 VDD.n482 10.6151
R4297 VDD.n1807 VDD.n482 10.6151
R4298 VDD.n1808 VDD.n1807 10.6151
R4299 VDD.n1809 VDD.n1808 10.6151
R4300 VDD.n1809 VDD.n469 10.6151
R4301 VDD.n1821 VDD.n469 10.6151
R4302 VDD.n1822 VDD.n1821 10.6151
R4303 VDD.n1823 VDD.n1822 10.6151
R4304 VDD.n1823 VDD.n453 10.6151
R4305 VDD.n1873 VDD.n453 10.6151
R4306 VDD.n1874 VDD.n1873 10.6151
R4307 VDD.n1875 VDD.n1874 10.6151
R4308 VDD.n1875 VDD.n442 10.6151
R4309 VDD.n2216 VDD.n2215 10.6151
R4310 VDD.n2215 VDD.n2214 10.6151
R4311 VDD.n2214 VDD.n2212 10.6151
R4312 VDD.n2212 VDD.n2211 10.6151
R4313 VDD.n2211 VDD.n2209 10.6151
R4314 VDD.n2209 VDD.n2208 10.6151
R4315 VDD.n2208 VDD.n2206 10.6151
R4316 VDD.n2206 VDD.n2205 10.6151
R4317 VDD.n2205 VDD.n2203 10.6151
R4318 VDD.n2203 VDD.n2202 10.6151
R4319 VDD.n2202 VDD.n2200 10.6151
R4320 VDD.n2200 VDD.n2199 10.6151
R4321 VDD.n2199 VDD.n2197 10.6151
R4322 VDD.n2197 VDD.n2196 10.6151
R4323 VDD.n2196 VDD.n2194 10.6151
R4324 VDD.n2194 VDD.n2193 10.6151
R4325 VDD.n2193 VDD.n2191 10.6151
R4326 VDD.n2191 VDD.n2190 10.6151
R4327 VDD.n2190 VDD.n2188 10.6151
R4328 VDD.n2188 VDD.n2187 10.6151
R4329 VDD.n2187 VDD.n2185 10.6151
R4330 VDD.n2185 VDD.n2184 10.6151
R4331 VDD.n2184 VDD.n2182 10.6151
R4332 VDD.n2182 VDD.n2181 10.6151
R4333 VDD.n2181 VDD.n2179 10.6151
R4334 VDD.n2179 VDD.n2178 10.6151
R4335 VDD.n2178 VDD.n2176 10.6151
R4336 VDD.n2176 VDD.n2175 10.6151
R4337 VDD.n2175 VDD.n2173 10.6151
R4338 VDD.n2173 VDD.n2172 10.6151
R4339 VDD.n2172 VDD.n2170 10.6151
R4340 VDD.n2170 VDD.n2169 10.6151
R4341 VDD.n2169 VDD.n2167 10.6151
R4342 VDD.n2167 VDD.n2166 10.6151
R4343 VDD.n2166 VDD.n2164 10.6151
R4344 VDD.n2164 VDD.n2163 10.6151
R4345 VDD.n2163 VDD.n2161 10.6151
R4346 VDD.n2161 VDD.n2160 10.6151
R4347 VDD.n2160 VDD.n2158 10.6151
R4348 VDD.n2158 VDD.n2157 10.6151
R4349 VDD.n2157 VDD.n2155 10.6151
R4350 VDD.n2155 VDD.n2154 10.6151
R4351 VDD.n2154 VDD.n2152 10.6151
R4352 VDD.n2152 VDD.n2151 10.6151
R4353 VDD.n2151 VDD.n2149 10.6151
R4354 VDD.n2149 VDD.n2148 10.6151
R4355 VDD.n2148 VDD.n2146 10.6151
R4356 VDD.n2146 VDD.n2145 10.6151
R4357 VDD.n2145 VDD.n2143 10.6151
R4358 VDD.n2143 VDD.n2142 10.6151
R4359 VDD.n2142 VDD.n2140 10.6151
R4360 VDD.n2140 VDD.n2139 10.6151
R4361 VDD.n2139 VDD.n2137 10.6151
R4362 VDD.n2137 VDD.n2136 10.6151
R4363 VDD.n2136 VDD.n2134 10.6151
R4364 VDD.n2134 VDD.n2133 10.6151
R4365 VDD.n2133 VDD.n2131 10.6151
R4366 VDD.n2131 VDD.n2130 10.6151
R4367 VDD.n2130 VDD.n2128 10.6151
R4368 VDD.n2128 VDD.n2127 10.6151
R4369 VDD.n2127 VDD.n2125 10.6151
R4370 VDD.n2125 VDD.n2124 10.6151
R4371 VDD.n2124 VDD.n2122 10.6151
R4372 VDD.n2122 VDD.n2121 10.6151
R4373 VDD.n2121 VDD.n2119 10.6151
R4374 VDD.n2119 VDD.n2118 10.6151
R4375 VDD.n2118 VDD.n2116 10.6151
R4376 VDD.n2116 VDD.n2115 10.6151
R4377 VDD.n2115 VDD.n2113 10.6151
R4378 VDD.n2113 VDD.n2112 10.6151
R4379 VDD.n2112 VDD.n2110 10.6151
R4380 VDD.n2110 VDD.n2109 10.6151
R4381 VDD.n2109 VDD.n2107 10.6151
R4382 VDD.n2107 VDD.n2106 10.6151
R4383 VDD.n2106 VDD.n2104 10.6151
R4384 VDD.n2104 VDD.n2103 10.6151
R4385 VDD.n2103 VDD.n2101 10.6151
R4386 VDD.n2101 VDD.n2100 10.6151
R4387 VDD.n2100 VDD.n2098 10.6151
R4388 VDD.n2098 VDD.n2097 10.6151
R4389 VDD.n2097 VDD.n2095 10.6151
R4390 VDD.n2095 VDD.n2094 10.6151
R4391 VDD.n2094 VDD.n2092 10.6151
R4392 VDD.n2092 VDD.n2091 10.6151
R4393 VDD.n2091 VDD.n2089 10.6151
R4394 VDD.n2089 VDD.n2088 10.6151
R4395 VDD.n2088 VDD.n157 10.6151
R4396 VDD.n2537 VDD.n157 10.6151
R4397 VDD.n2538 VDD.n2537 10.6151
R4398 VDD.n2539 VDD.n2538 10.6151
R4399 VDD.n2244 VDD.n2243 10.6151
R4400 VDD.n2243 VDD.n2242 10.6151
R4401 VDD.n2242 VDD.n2241 10.6151
R4402 VDD.n2241 VDD.n2239 10.6151
R4403 VDD.n2239 VDD.n2236 10.6151
R4404 VDD.n2236 VDD.n2235 10.6151
R4405 VDD.n2235 VDD.n2232 10.6151
R4406 VDD.n2232 VDD.n2231 10.6151
R4407 VDD.n2231 VDD.n2228 10.6151
R4408 VDD.n2228 VDD.n2227 10.6151
R4409 VDD.n2227 VDD.n2224 10.6151
R4410 VDD.n2224 VDD.n2223 10.6151
R4411 VDD.n2220 VDD.n2219 10.6151
R4412 VDD.n2256 VDD.n416 10.6151
R4413 VDD.n2257 VDD.n2256 10.6151
R4414 VDD.n2258 VDD.n2257 10.6151
R4415 VDD.n2258 VDD.n404 10.6151
R4416 VDD.n2268 VDD.n404 10.6151
R4417 VDD.n2269 VDD.n2268 10.6151
R4418 VDD.n2270 VDD.n2269 10.6151
R4419 VDD.n2270 VDD.n392 10.6151
R4420 VDD.n2280 VDD.n392 10.6151
R4421 VDD.n2281 VDD.n2280 10.6151
R4422 VDD.n2282 VDD.n2281 10.6151
R4423 VDD.n2282 VDD.n380 10.6151
R4424 VDD.n2292 VDD.n380 10.6151
R4425 VDD.n2293 VDD.n2292 10.6151
R4426 VDD.n2294 VDD.n2293 10.6151
R4427 VDD.n2294 VDD.n368 10.6151
R4428 VDD.n2304 VDD.n368 10.6151
R4429 VDD.n2305 VDD.n2304 10.6151
R4430 VDD.n2306 VDD.n2305 10.6151
R4431 VDD.n2306 VDD.n356 10.6151
R4432 VDD.n2316 VDD.n356 10.6151
R4433 VDD.n2317 VDD.n2316 10.6151
R4434 VDD.n2318 VDD.n2317 10.6151
R4435 VDD.n2318 VDD.n344 10.6151
R4436 VDD.n2328 VDD.n344 10.6151
R4437 VDD.n2329 VDD.n2328 10.6151
R4438 VDD.n2330 VDD.n2329 10.6151
R4439 VDD.n2330 VDD.n332 10.6151
R4440 VDD.n2340 VDD.n332 10.6151
R4441 VDD.n2341 VDD.n2340 10.6151
R4442 VDD.n2342 VDD.n2341 10.6151
R4443 VDD.n2342 VDD.n319 10.6151
R4444 VDD.n2352 VDD.n319 10.6151
R4445 VDD.n2353 VDD.n2352 10.6151
R4446 VDD.n2354 VDD.n2353 10.6151
R4447 VDD.n2354 VDD.n307 10.6151
R4448 VDD.n2364 VDD.n307 10.6151
R4449 VDD.n2365 VDD.n2364 10.6151
R4450 VDD.n2366 VDD.n2365 10.6151
R4451 VDD.n2366 VDD.n296 10.6151
R4452 VDD.n2376 VDD.n296 10.6151
R4453 VDD.n2377 VDD.n2376 10.6151
R4454 VDD.n2378 VDD.n2377 10.6151
R4455 VDD.n2378 VDD.n284 10.6151
R4456 VDD.n2388 VDD.n284 10.6151
R4457 VDD.n2389 VDD.n2388 10.6151
R4458 VDD.n2390 VDD.n2389 10.6151
R4459 VDD.n2390 VDD.n272 10.6151
R4460 VDD.n2400 VDD.n272 10.6151
R4461 VDD.n2401 VDD.n2400 10.6151
R4462 VDD.n2402 VDD.n2401 10.6151
R4463 VDD.n2402 VDD.n260 10.6151
R4464 VDD.n2412 VDD.n260 10.6151
R4465 VDD.n2413 VDD.n2412 10.6151
R4466 VDD.n2414 VDD.n2413 10.6151
R4467 VDD.n2414 VDD.n248 10.6151
R4468 VDD.n2424 VDD.n248 10.6151
R4469 VDD.n2425 VDD.n2424 10.6151
R4470 VDD.n2426 VDD.n2425 10.6151
R4471 VDD.n2426 VDD.n236 10.6151
R4472 VDD.n2436 VDD.n236 10.6151
R4473 VDD.n2437 VDD.n2436 10.6151
R4474 VDD.n2438 VDD.n2437 10.6151
R4475 VDD.n2438 VDD.n224 10.6151
R4476 VDD.n2448 VDD.n224 10.6151
R4477 VDD.n2449 VDD.n2448 10.6151
R4478 VDD.n2450 VDD.n2449 10.6151
R4479 VDD.n2450 VDD.n212 10.6151
R4480 VDD.n2460 VDD.n212 10.6151
R4481 VDD.n2461 VDD.n2460 10.6151
R4482 VDD.n2462 VDD.n2461 10.6151
R4483 VDD.n2462 VDD.n200 10.6151
R4484 VDD.n2472 VDD.n200 10.6151
R4485 VDD.n2473 VDD.n2472 10.6151
R4486 VDD.n2474 VDD.n2473 10.6151
R4487 VDD.n2474 VDD.n188 10.6151
R4488 VDD.n2484 VDD.n188 10.6151
R4489 VDD.n2485 VDD.n2484 10.6151
R4490 VDD.n2486 VDD.n2485 10.6151
R4491 VDD.n2486 VDD.n175 10.6151
R4492 VDD.n2496 VDD.n175 10.6151
R4493 VDD.n2497 VDD.n2496 10.6151
R4494 VDD.n2498 VDD.n2497 10.6151
R4495 VDD.n2498 VDD.n163 10.6151
R4496 VDD.n2530 VDD.n163 10.6151
R4497 VDD.n2531 VDD.n2530 10.6151
R4498 VDD.n2532 VDD.n2531 10.6151
R4499 VDD.n2532 VDD.n142 10.6151
R4500 VDD.n2569 VDD.n142 10.6151
R4501 VDD.n2569 VDD.n2568 10.6151
R4502 VDD.n2567 VDD.n143 10.6151
R4503 VDD.n2562 VDD.n143 10.6151
R4504 VDD.n2562 VDD.n2561 10.6151
R4505 VDD.n2561 VDD.n2560 10.6151
R4506 VDD.n2560 VDD.n145 10.6151
R4507 VDD.n2555 VDD.n145 10.6151
R4508 VDD.n2555 VDD.n2554 10.6151
R4509 VDD.n2554 VDD.n2552 10.6151
R4510 VDD.n2552 VDD.n148 10.6151
R4511 VDD.n2547 VDD.n148 10.6151
R4512 VDD.n2547 VDD.n2546 10.6151
R4513 VDD.n2546 VDD.n2545 10.6151
R4514 VDD.n2540 VDD.n155 10.6151
R4515 VDD.n2505 VDD.n2504 10.6151
R4516 VDD.n2514 VDD.n2505 10.6151
R4517 VDD.n2514 VDD.n2513 10.6151
R4518 VDD.n2513 VDD.n2512 10.6151
R4519 VDD.n2512 VDD.n2507 10.6151
R4520 VDD.n2507 VDD.n122 10.6151
R4521 VDD.n2589 VDD.n122 10.6151
R4522 VDD.n2589 VDD.n123 10.6151
R4523 VDD.n126 VDD.n123 10.6151
R4524 VDD.n2582 VDD.n126 10.6151
R4525 VDD.n2582 VDD.n2581 10.6151
R4526 VDD.n2581 VDD.n2580 10.6151
R4527 VDD.n2575 VDD.n132 10.6151
R4528 VDD.n2080 VDD.n2079 10.6151
R4529 VDD.n2079 VDD.n2078 10.6151
R4530 VDD.n2078 VDD.n2076 10.6151
R4531 VDD.n2076 VDD.n2075 10.6151
R4532 VDD.n2075 VDD.n2073 10.6151
R4533 VDD.n2073 VDD.n2072 10.6151
R4534 VDD.n2072 VDD.n2070 10.6151
R4535 VDD.n2070 VDD.n2069 10.6151
R4536 VDD.n2069 VDD.n2067 10.6151
R4537 VDD.n2067 VDD.n2066 10.6151
R4538 VDD.n2066 VDD.n2064 10.6151
R4539 VDD.n2064 VDD.n2063 10.6151
R4540 VDD.n2063 VDD.n2061 10.6151
R4541 VDD.n2061 VDD.n2060 10.6151
R4542 VDD.n2060 VDD.n2058 10.6151
R4543 VDD.n2058 VDD.n2057 10.6151
R4544 VDD.n2057 VDD.n2055 10.6151
R4545 VDD.n2055 VDD.n2054 10.6151
R4546 VDD.n2054 VDD.n2052 10.6151
R4547 VDD.n2052 VDD.n2051 10.6151
R4548 VDD.n2051 VDD.n2049 10.6151
R4549 VDD.n2049 VDD.n2048 10.6151
R4550 VDD.n2048 VDD.n2046 10.6151
R4551 VDD.n2046 VDD.n2045 10.6151
R4552 VDD.n2045 VDD.n2043 10.6151
R4553 VDD.n2043 VDD.n2042 10.6151
R4554 VDD.n2042 VDD.n2040 10.6151
R4555 VDD.n2040 VDD.n2039 10.6151
R4556 VDD.n2039 VDD.n2037 10.6151
R4557 VDD.n2037 VDD.n2036 10.6151
R4558 VDD.n2036 VDD.n2034 10.6151
R4559 VDD.n2034 VDD.n2033 10.6151
R4560 VDD.n2033 VDD.n2031 10.6151
R4561 VDD.n2031 VDD.n2030 10.6151
R4562 VDD.n2030 VDD.n2028 10.6151
R4563 VDD.n2028 VDD.n2027 10.6151
R4564 VDD.n2027 VDD.n2025 10.6151
R4565 VDD.n2025 VDD.n2024 10.6151
R4566 VDD.n2024 VDD.n2022 10.6151
R4567 VDD.n2022 VDD.n2021 10.6151
R4568 VDD.n2021 VDD.n2019 10.6151
R4569 VDD.n2019 VDD.n2018 10.6151
R4570 VDD.n2018 VDD.n2016 10.6151
R4571 VDD.n2016 VDD.n2015 10.6151
R4572 VDD.n2015 VDD.n2013 10.6151
R4573 VDD.n2013 VDD.n2012 10.6151
R4574 VDD.n2012 VDD.n2010 10.6151
R4575 VDD.n2010 VDD.n2009 10.6151
R4576 VDD.n2009 VDD.n2007 10.6151
R4577 VDD.n2007 VDD.n2006 10.6151
R4578 VDD.n2006 VDD.n2004 10.6151
R4579 VDD.n2004 VDD.n2003 10.6151
R4580 VDD.n2003 VDD.n2001 10.6151
R4581 VDD.n2001 VDD.n2000 10.6151
R4582 VDD.n2000 VDD.n1998 10.6151
R4583 VDD.n1998 VDD.n1997 10.6151
R4584 VDD.n1997 VDD.n1995 10.6151
R4585 VDD.n1995 VDD.n1994 10.6151
R4586 VDD.n1994 VDD.n1992 10.6151
R4587 VDD.n1992 VDD.n1991 10.6151
R4588 VDD.n1991 VDD.n1989 10.6151
R4589 VDD.n1989 VDD.n1988 10.6151
R4590 VDD.n1988 VDD.n1986 10.6151
R4591 VDD.n1986 VDD.n1985 10.6151
R4592 VDD.n1985 VDD.n1983 10.6151
R4593 VDD.n1983 VDD.n1982 10.6151
R4594 VDD.n1982 VDD.n1980 10.6151
R4595 VDD.n1980 VDD.n1979 10.6151
R4596 VDD.n1979 VDD.n1977 10.6151
R4597 VDD.n1977 VDD.n1976 10.6151
R4598 VDD.n1976 VDD.n1974 10.6151
R4599 VDD.n1974 VDD.n1973 10.6151
R4600 VDD.n1973 VDD.n1971 10.6151
R4601 VDD.n1971 VDD.n1970 10.6151
R4602 VDD.n1970 VDD.n1968 10.6151
R4603 VDD.n1968 VDD.n1967 10.6151
R4604 VDD.n1967 VDD.n1965 10.6151
R4605 VDD.n1965 VDD.n1964 10.6151
R4606 VDD.n1964 VDD.n1962 10.6151
R4607 VDD.n1962 VDD.n1961 10.6151
R4608 VDD.n1961 VDD.n1959 10.6151
R4609 VDD.n1959 VDD.n1958 10.6151
R4610 VDD.n1958 VDD.n1956 10.6151
R4611 VDD.n1956 VDD.n1955 10.6151
R4612 VDD.n1955 VDD.n1953 10.6151
R4613 VDD.n1953 VDD.n1952 10.6151
R4614 VDD.n1952 VDD.n1950 10.6151
R4615 VDD.n1950 VDD.n134 10.6151
R4616 VDD.n2573 VDD.n134 10.6151
R4617 VDD.n2574 VDD.n2573 10.6151
R4618 VDD.n2250 VDD.n422 10.6151
R4619 VDD.n1927 VDD.n422 10.6151
R4620 VDD.n1928 VDD.n1927 10.6151
R4621 VDD.n1931 VDD.n1928 10.6151
R4622 VDD.n1932 VDD.n1931 10.6151
R4623 VDD.n1935 VDD.n1932 10.6151
R4624 VDD.n1936 VDD.n1935 10.6151
R4625 VDD.n1939 VDD.n1936 10.6151
R4626 VDD.n1940 VDD.n1939 10.6151
R4627 VDD.n1943 VDD.n1940 10.6151
R4628 VDD.n1944 VDD.n1943 10.6151
R4629 VDD.n1947 VDD.n1944 10.6151
R4630 VDD.n2081 VDD.n1949 10.6151
R4631 VDD.n2252 VDD.n2251 10.6151
R4632 VDD.n2252 VDD.n410 10.6151
R4633 VDD.n2262 VDD.n410 10.6151
R4634 VDD.n2263 VDD.n2262 10.6151
R4635 VDD.n2264 VDD.n2263 10.6151
R4636 VDD.n2264 VDD.n398 10.6151
R4637 VDD.n2274 VDD.n398 10.6151
R4638 VDD.n2275 VDD.n2274 10.6151
R4639 VDD.n2276 VDD.n2275 10.6151
R4640 VDD.n2276 VDD.n386 10.6151
R4641 VDD.n2286 VDD.n386 10.6151
R4642 VDD.n2287 VDD.n2286 10.6151
R4643 VDD.n2288 VDD.n2287 10.6151
R4644 VDD.n2288 VDD.n374 10.6151
R4645 VDD.n2298 VDD.n374 10.6151
R4646 VDD.n2299 VDD.n2298 10.6151
R4647 VDD.n2300 VDD.n2299 10.6151
R4648 VDD.n2300 VDD.n361 10.6151
R4649 VDD.n2310 VDD.n361 10.6151
R4650 VDD.n2311 VDD.n2310 10.6151
R4651 VDD.n2312 VDD.n2311 10.6151
R4652 VDD.n2312 VDD.n349 10.6151
R4653 VDD.n2322 VDD.n349 10.6151
R4654 VDD.n2323 VDD.n2322 10.6151
R4655 VDD.n2324 VDD.n2323 10.6151
R4656 VDD.n2324 VDD.n338 10.6151
R4657 VDD.n2334 VDD.n338 10.6151
R4658 VDD.n2335 VDD.n2334 10.6151
R4659 VDD.n2336 VDD.n2335 10.6151
R4660 VDD.n2336 VDD.n326 10.6151
R4661 VDD.n2346 VDD.n326 10.6151
R4662 VDD.n2347 VDD.n2346 10.6151
R4663 VDD.n2348 VDD.n2347 10.6151
R4664 VDD.n2348 VDD.n314 10.6151
R4665 VDD.n2358 VDD.n314 10.6151
R4666 VDD.n2359 VDD.n2358 10.6151
R4667 VDD.n2360 VDD.n2359 10.6151
R4668 VDD.n2360 VDD.n302 10.6151
R4669 VDD.n2370 VDD.n302 10.6151
R4670 VDD.n2371 VDD.n2370 10.6151
R4671 VDD.n2372 VDD.n2371 10.6151
R4672 VDD.n2372 VDD.n290 10.6151
R4673 VDD.n2382 VDD.n290 10.6151
R4674 VDD.n2383 VDD.n2382 10.6151
R4675 VDD.n2384 VDD.n2383 10.6151
R4676 VDD.n2384 VDD.n278 10.6151
R4677 VDD.n2394 VDD.n278 10.6151
R4678 VDD.n2395 VDD.n2394 10.6151
R4679 VDD.n2396 VDD.n2395 10.6151
R4680 VDD.n2396 VDD.n266 10.6151
R4681 VDD.n2406 VDD.n266 10.6151
R4682 VDD.n2407 VDD.n2406 10.6151
R4683 VDD.n2408 VDD.n2407 10.6151
R4684 VDD.n2408 VDD.n254 10.6151
R4685 VDD.n2418 VDD.n254 10.6151
R4686 VDD.n2419 VDD.n2418 10.6151
R4687 VDD.n2420 VDD.n2419 10.6151
R4688 VDD.n2420 VDD.n242 10.6151
R4689 VDD.n2430 VDD.n242 10.6151
R4690 VDD.n2431 VDD.n2430 10.6151
R4691 VDD.n2432 VDD.n2431 10.6151
R4692 VDD.n2432 VDD.n230 10.6151
R4693 VDD.n2442 VDD.n230 10.6151
R4694 VDD.n2443 VDD.n2442 10.6151
R4695 VDD.n2444 VDD.n2443 10.6151
R4696 VDD.n2444 VDD.n217 10.6151
R4697 VDD.n2454 VDD.n217 10.6151
R4698 VDD.n2455 VDD.n2454 10.6151
R4699 VDD.n2456 VDD.n2455 10.6151
R4700 VDD.n2456 VDD.n206 10.6151
R4701 VDD.n2466 VDD.n206 10.6151
R4702 VDD.n2467 VDD.n2466 10.6151
R4703 VDD.n2468 VDD.n2467 10.6151
R4704 VDD.n2468 VDD.n194 10.6151
R4705 VDD.n2478 VDD.n194 10.6151
R4706 VDD.n2479 VDD.n2478 10.6151
R4707 VDD.n2480 VDD.n2479 10.6151
R4708 VDD.n2480 VDD.n182 10.6151
R4709 VDD.n2490 VDD.n182 10.6151
R4710 VDD.n2491 VDD.n2490 10.6151
R4711 VDD.n2492 VDD.n2491 10.6151
R4712 VDD.n2492 VDD.n170 10.6151
R4713 VDD.n2502 VDD.n170 10.6151
R4714 VDD.n2503 VDD.n2502 10.6151
R4715 VDD.n2526 VDD.n2503 10.6151
R4716 VDD.n2526 VDD.n2525 10.6151
R4717 VDD.n2525 VDD.n2524 10.6151
R4718 VDD.n2524 VDD.n2523 10.6151
R4719 VDD.n2523 VDD.n2521 10.6151
R4720 VDD.n2521 VDD.n2520 10.6151
R4721 VDD.n1573 VDD.n716 10.6151
R4722 VDD.n1574 VDD.n1573 10.6151
R4723 VDD.n1575 VDD.n1574 10.6151
R4724 VDD.n1575 VDD.n704 10.6151
R4725 VDD.n1585 VDD.n704 10.6151
R4726 VDD.n1586 VDD.n1585 10.6151
R4727 VDD.n1587 VDD.n1586 10.6151
R4728 VDD.n1587 VDD.n692 10.6151
R4729 VDD.n1597 VDD.n692 10.6151
R4730 VDD.n1598 VDD.n1597 10.6151
R4731 VDD.n1599 VDD.n1598 10.6151
R4732 VDD.n1599 VDD.n680 10.6151
R4733 VDD.n1609 VDD.n680 10.6151
R4734 VDD.n1610 VDD.n1609 10.6151
R4735 VDD.n1611 VDD.n1610 10.6151
R4736 VDD.n1611 VDD.n668 10.6151
R4737 VDD.n1621 VDD.n668 10.6151
R4738 VDD.n1622 VDD.n1621 10.6151
R4739 VDD.n1623 VDD.n1622 10.6151
R4740 VDD.n1623 VDD.n656 10.6151
R4741 VDD.n1633 VDD.n656 10.6151
R4742 VDD.n1634 VDD.n1633 10.6151
R4743 VDD.n1635 VDD.n1634 10.6151
R4744 VDD.n1635 VDD.n644 10.6151
R4745 VDD.n1645 VDD.n644 10.6151
R4746 VDD.n1646 VDD.n1645 10.6151
R4747 VDD.n1647 VDD.n1646 10.6151
R4748 VDD.n1647 VDD.n632 10.6151
R4749 VDD.n1657 VDD.n632 10.6151
R4750 VDD.n1658 VDD.n1657 10.6151
R4751 VDD.n1659 VDD.n1658 10.6151
R4752 VDD.n1659 VDD.n620 10.6151
R4753 VDD.n1669 VDD.n620 10.6151
R4754 VDD.n1670 VDD.n1669 10.6151
R4755 VDD.n1671 VDD.n1670 10.6151
R4756 VDD.n1671 VDD.n607 10.6151
R4757 VDD.n1681 VDD.n607 10.6151
R4758 VDD.n1682 VDD.n1681 10.6151
R4759 VDD.n1683 VDD.n1682 10.6151
R4760 VDD.n1683 VDD.n595 10.6151
R4761 VDD.n1693 VDD.n595 10.6151
R4762 VDD.n1694 VDD.n1693 10.6151
R4763 VDD.n1695 VDD.n1694 10.6151
R4764 VDD.n1695 VDD.n584 10.6151
R4765 VDD.n1705 VDD.n584 10.6151
R4766 VDD.n1706 VDD.n1705 10.6151
R4767 VDD.n1707 VDD.n1706 10.6151
R4768 VDD.n1707 VDD.n572 10.6151
R4769 VDD.n1717 VDD.n572 10.6151
R4770 VDD.n1718 VDD.n1717 10.6151
R4771 VDD.n1719 VDD.n1718 10.6151
R4772 VDD.n1719 VDD.n560 10.6151
R4773 VDD.n1729 VDD.n560 10.6151
R4774 VDD.n1730 VDD.n1729 10.6151
R4775 VDD.n1731 VDD.n1730 10.6151
R4776 VDD.n1731 VDD.n548 10.6151
R4777 VDD.n1741 VDD.n548 10.6151
R4778 VDD.n1742 VDD.n1741 10.6151
R4779 VDD.n1743 VDD.n1742 10.6151
R4780 VDD.n1743 VDD.n536 10.6151
R4781 VDD.n1753 VDD.n536 10.6151
R4782 VDD.n1754 VDD.n1753 10.6151
R4783 VDD.n1755 VDD.n1754 10.6151
R4784 VDD.n1755 VDD.n524 10.6151
R4785 VDD.n1765 VDD.n524 10.6151
R4786 VDD.n1766 VDD.n1765 10.6151
R4787 VDD.n1767 VDD.n1766 10.6151
R4788 VDD.n1767 VDD.n512 10.6151
R4789 VDD.n1777 VDD.n512 10.6151
R4790 VDD.n1778 VDD.n1777 10.6151
R4791 VDD.n1779 VDD.n1778 10.6151
R4792 VDD.n1779 VDD.n500 10.6151
R4793 VDD.n1789 VDD.n500 10.6151
R4794 VDD.n1790 VDD.n1789 10.6151
R4795 VDD.n1791 VDD.n1790 10.6151
R4796 VDD.n1791 VDD.n488 10.6151
R4797 VDD.n1801 VDD.n488 10.6151
R4798 VDD.n1802 VDD.n1801 10.6151
R4799 VDD.n1803 VDD.n1802 10.6151
R4800 VDD.n1803 VDD.n475 10.6151
R4801 VDD.n1813 VDD.n475 10.6151
R4802 VDD.n1814 VDD.n1813 10.6151
R4803 VDD.n1817 VDD.n1814 10.6151
R4804 VDD.n1817 VDD.n1816 10.6151
R4805 VDD.n1816 VDD.n1815 10.6151
R4806 VDD.n1815 VDD.n460 10.6151
R4807 VDD.n1869 VDD.n460 10.6151
R4808 VDD.n1869 VDD.n1868 10.6151
R4809 VDD.n1868 VDD.n1867 10.6151
R4810 VDD.n1867 VDD.n1866 10.6151
R4811 VDD.n1863 VDD.n1862 10.6151
R4812 VDD.n1862 VDD.n1859 10.6151
R4813 VDD.n1859 VDD.n1858 10.6151
R4814 VDD.n1858 VDD.n1855 10.6151
R4815 VDD.n1855 VDD.n1854 10.6151
R4816 VDD.n1854 VDD.n1851 10.6151
R4817 VDD.n1851 VDD.n1850 10.6151
R4818 VDD.n1850 VDD.n1847 10.6151
R4819 VDD.n1847 VDD.n1846 10.6151
R4820 VDD.n1846 VDD.n1843 10.6151
R4821 VDD.n1843 VDD.n1842 10.6151
R4822 VDD.n1842 VDD.n1839 10.6151
R4823 VDD.n1837 VDD.n1835 10.6151
R4824 VDD.n934 VDD.n932 10.6151
R4825 VDD.n932 VDD.n931 10.6151
R4826 VDD.n931 VDD.n929 10.6151
R4827 VDD.n929 VDD.n928 10.6151
R4828 VDD.n928 VDD.n926 10.6151
R4829 VDD.n926 VDD.n925 10.6151
R4830 VDD.n925 VDD.n923 10.6151
R4831 VDD.n923 VDD.n922 10.6151
R4832 VDD.n922 VDD.n920 10.6151
R4833 VDD.n920 VDD.n919 10.6151
R4834 VDD.n919 VDD.n917 10.6151
R4835 VDD.n917 VDD.n916 10.6151
R4836 VDD.n916 VDD.n914 10.6151
R4837 VDD.n914 VDD.n913 10.6151
R4838 VDD.n913 VDD.n911 10.6151
R4839 VDD.n911 VDD.n910 10.6151
R4840 VDD.n910 VDD.n908 10.6151
R4841 VDD.n908 VDD.n907 10.6151
R4842 VDD.n907 VDD.n905 10.6151
R4843 VDD.n905 VDD.n904 10.6151
R4844 VDD.n904 VDD.n902 10.6151
R4845 VDD.n902 VDD.n901 10.6151
R4846 VDD.n901 VDD.n899 10.6151
R4847 VDD.n899 VDD.n898 10.6151
R4848 VDD.n898 VDD.n896 10.6151
R4849 VDD.n896 VDD.n895 10.6151
R4850 VDD.n895 VDD.n893 10.6151
R4851 VDD.n893 VDD.n892 10.6151
R4852 VDD.n892 VDD.n890 10.6151
R4853 VDD.n890 VDD.n889 10.6151
R4854 VDD.n889 VDD.n887 10.6151
R4855 VDD.n887 VDD.n886 10.6151
R4856 VDD.n886 VDD.n884 10.6151
R4857 VDD.n884 VDD.n883 10.6151
R4858 VDD.n883 VDD.n881 10.6151
R4859 VDD.n881 VDD.n880 10.6151
R4860 VDD.n880 VDD.n878 10.6151
R4861 VDD.n878 VDD.n877 10.6151
R4862 VDD.n877 VDD.n875 10.6151
R4863 VDD.n875 VDD.n874 10.6151
R4864 VDD.n874 VDD.n872 10.6151
R4865 VDD.n872 VDD.n871 10.6151
R4866 VDD.n871 VDD.n869 10.6151
R4867 VDD.n869 VDD.n868 10.6151
R4868 VDD.n868 VDD.n866 10.6151
R4869 VDD.n866 VDD.n865 10.6151
R4870 VDD.n865 VDD.n863 10.6151
R4871 VDD.n863 VDD.n862 10.6151
R4872 VDD.n862 VDD.n860 10.6151
R4873 VDD.n860 VDD.n859 10.6151
R4874 VDD.n859 VDD.n857 10.6151
R4875 VDD.n857 VDD.n856 10.6151
R4876 VDD.n856 VDD.n854 10.6151
R4877 VDD.n854 VDD.n853 10.6151
R4878 VDD.n853 VDD.n851 10.6151
R4879 VDD.n851 VDD.n850 10.6151
R4880 VDD.n850 VDD.n848 10.6151
R4881 VDD.n848 VDD.n847 10.6151
R4882 VDD.n847 VDD.n845 10.6151
R4883 VDD.n845 VDD.n844 10.6151
R4884 VDD.n844 VDD.n842 10.6151
R4885 VDD.n842 VDD.n841 10.6151
R4886 VDD.n841 VDD.n839 10.6151
R4887 VDD.n839 VDD.n838 10.6151
R4888 VDD.n838 VDD.n836 10.6151
R4889 VDD.n836 VDD.n835 10.6151
R4890 VDD.n835 VDD.n833 10.6151
R4891 VDD.n833 VDD.n832 10.6151
R4892 VDD.n832 VDD.n830 10.6151
R4893 VDD.n830 VDD.n829 10.6151
R4894 VDD.n829 VDD.n827 10.6151
R4895 VDD.n827 VDD.n826 10.6151
R4896 VDD.n826 VDD.n824 10.6151
R4897 VDD.n824 VDD.n823 10.6151
R4898 VDD.n823 VDD.n821 10.6151
R4899 VDD.n821 VDD.n820 10.6151
R4900 VDD.n820 VDD.n818 10.6151
R4901 VDD.n818 VDD.n817 10.6151
R4902 VDD.n817 VDD.n815 10.6151
R4903 VDD.n815 VDD.n814 10.6151
R4904 VDD.n814 VDD.n812 10.6151
R4905 VDD.n812 VDD.n811 10.6151
R4906 VDD.n811 VDD.n809 10.6151
R4907 VDD.n809 VDD.n808 10.6151
R4908 VDD.n808 VDD.n463 10.6151
R4909 VDD.n1828 VDD.n463 10.6151
R4910 VDD.n1829 VDD.n1828 10.6151
R4911 VDD.n1831 VDD.n1829 10.6151
R4912 VDD.n1832 VDD.n1831 10.6151
R4913 VDD.n1834 VDD.n1832 10.6151
R4914 VDD.n793 VDD.n792 10.6151
R4915 VDD.n796 VDD.n793 10.6151
R4916 VDD.n797 VDD.n796 10.6151
R4917 VDD.n800 VDD.n797 10.6151
R4918 VDD.n801 VDD.n800 10.6151
R4919 VDD.n804 VDD.n801 10.6151
R4920 VDD.n949 VDD.n804 10.6151
R4921 VDD.n949 VDD.n948 10.6151
R4922 VDD.n948 VDD.n946 10.6151
R4923 VDD.n946 VDD.n943 10.6151
R4924 VDD.n943 VDD.n942 10.6151
R4925 VDD.n942 VDD.n939 10.6151
R4926 VDD.n937 VDD.n935 10.6151
R4927 VDD.n1553 VDD.n1402 10.4202
R4928 VDD.n2554 VDD.n2553 10.4202
R4929 VDD.n2608 VDD.n2589 10.4202
R4930 VDD.n1349 VDD.n949 10.4202
R4931 VDD.n1685 VDD.t101 10.3521
R4932 VDD.n1721 VDD.t100 10.3521
R4933 VDD.n2368 VDD.t93 10.3521
R4934 VDD.n2404 VDD.t90 10.3521
R4935 VDD.n1265 VDD.n1264 9.3005
R4936 VDD.n1001 VDD.n1000 9.3005
R4937 VDD.n1278 VDD.n1277 9.3005
R4938 VDD.n1279 VDD.n999 9.3005
R4939 VDD.n1281 VDD.n1280 9.3005
R4940 VDD.n989 VDD.n988 9.3005
R4941 VDD.n1294 VDD.n1293 9.3005
R4942 VDD.n1295 VDD.n987 9.3005
R4943 VDD.n1297 VDD.n1296 9.3005
R4944 VDD.n976 VDD.n975 9.3005
R4945 VDD.n1312 VDD.n1311 9.3005
R4946 VDD.n1313 VDD.n974 9.3005
R4947 VDD.n1332 VDD.n1331 9.3005
R4948 VDD.n1387 VDD.n749 9.3005
R4949 VDD.n1386 VDD.n1385 9.3005
R4950 VDD.n755 VDD.n754 9.3005
R4951 VDD.n1380 VDD.n759 9.3005
R4952 VDD.n1379 VDD.n760 9.3005
R4953 VDD.n1378 VDD.n761 9.3005
R4954 VDD.n765 VDD.n762 9.3005
R4955 VDD.n1373 VDD.n766 9.3005
R4956 VDD.n1372 VDD.n767 9.3005
R4957 VDD.n1371 VDD.n768 9.3005
R4958 VDD.n772 VDD.n769 9.3005
R4959 VDD.n1366 VDD.n773 9.3005
R4960 VDD.n1365 VDD.n774 9.3005
R4961 VDD.n1364 VDD.n775 9.3005
R4962 VDD.n781 VDD.n778 9.3005
R4963 VDD.n1359 VDD.n782 9.3005
R4964 VDD.n1358 VDD.n783 9.3005
R4965 VDD.n1357 VDD.n784 9.3005
R4966 VDD.n788 VDD.n785 9.3005
R4967 VDD.n1352 VDD.n789 9.3005
R4968 VDD.n1389 VDD.n1388 9.3005
R4969 VDD.n1328 VDD.n1314 9.3005
R4970 VDD.n1318 VDD.n1315 9.3005
R4971 VDD.n1319 VDD.n1316 9.3005
R4972 VDD.n1321 VDD.n1320 9.3005
R4973 VDD.n743 VDD.n739 9.3005
R4974 VDD.n1391 VDD.n740 9.3005
R4975 VDD.n1390 VDD.n748 9.3005
R4976 VDD.n1330 VDD.n1329 9.3005
R4977 VDD.n2624 VDD.n2623 9.3005
R4978 VDD.n2627 VDD.n113 9.3005
R4979 VDD.n2628 VDD.n112 9.3005
R4980 VDD.n2631 VDD.n111 9.3005
R4981 VDD.n2632 VDD.n110 9.3005
R4982 VDD.n2635 VDD.n109 9.3005
R4983 VDD.n2636 VDD.n108 9.3005
R4984 VDD.n2639 VDD.n107 9.3005
R4985 VDD.n2640 VDD.n106 9.3005
R4986 VDD.n2643 VDD.n105 9.3005
R4987 VDD.n2644 VDD.n104 9.3005
R4988 VDD.n2647 VDD.n103 9.3005
R4989 VDD.n2648 VDD.n102 9.3005
R4990 VDD.n2652 VDD.n2651 9.3005
R4991 VDD.n2653 VDD.n99 9.3005
R4992 VDD.n2657 VDD.n2654 9.3005
R4993 VDD.n2658 VDD.n98 9.3005
R4994 VDD.n2661 VDD.n97 9.3005
R4995 VDD.n2670 VDD.n94 9.3005
R4996 VDD.n2673 VDD.n93 9.3005
R4997 VDD.n2675 VDD.n92 9.3005
R4998 VDD.n2676 VDD.n91 9.3005
R4999 VDD.n2677 VDD.n90 9.3005
R5000 VDD.n2678 VDD.n89 9.3005
R5001 VDD.n58 VDD.n57 9.3005
R5002 VDD.n2693 VDD.n2692 9.3005
R5003 VDD.n2694 VDD.n56 9.3005
R5004 VDD.n2696 VDD.n2695 9.3005
R5005 VDD.n46 VDD.n45 9.3005
R5006 VDD.n2709 VDD.n2708 9.3005
R5007 VDD.n2710 VDD.n44 9.3005
R5008 VDD.n2712 VDD.n2711 9.3005
R5009 VDD.n34 VDD.n33 9.3005
R5010 VDD.n2725 VDD.n2724 9.3005
R5011 VDD.n2726 VDD.n32 9.3005
R5012 VDD.n2728 VDD.n2727 9.3005
R5013 VDD.n18 VDD.n16 9.3005
R5014 VDD.n2984 VDD.n2983 9.3005
R5015 VDD.n19 VDD.n17 9.3005
R5016 VDD.n2974 VDD.n2742 9.3005
R5017 VDD.n2973 VDD.n2743 9.3005
R5018 VDD.n2972 VDD.n2744 9.3005
R5019 VDD.n2752 VDD.n2745 9.3005
R5020 VDD.n2966 VDD.n2753 9.3005
R5021 VDD.n2965 VDD.n2754 9.3005
R5022 VDD.n2964 VDD.n2755 9.3005
R5023 VDD.n2763 VDD.n2756 9.3005
R5024 VDD.n2958 VDD.n2764 9.3005
R5025 VDD.n2957 VDD.n2765 9.3005
R5026 VDD.n2956 VDD.n2766 9.3005
R5027 VDD.n2793 VDD.n2767 9.3005
R5028 VDD.n2949 VDD.n2948 9.3005
R5029 VDD.n2947 VDD.n2795 9.3005
R5030 VDD.n2946 VDD.n2945 9.3005
R5031 VDD.n2942 VDD.n2796 9.3005
R5032 VDD.n2939 VDD.n2797 9.3005
R5033 VDD.n2938 VDD.n2798 9.3005
R5034 VDD.n2935 VDD.n2799 9.3005
R5035 VDD.n2934 VDD.n2800 9.3005
R5036 VDD.n2931 VDD.n2801 9.3005
R5037 VDD.n2930 VDD.n2802 9.3005
R5038 VDD.n2927 VDD.n2803 9.3005
R5039 VDD.n2926 VDD.n2925 9.3005
R5040 VDD.n2924 VDD.n2804 9.3005
R5041 VDD.n2923 VDD.n2922 9.3005
R5042 VDD.n2919 VDD.n2809 9.3005
R5043 VDD.n2918 VDD.n2810 9.3005
R5044 VDD.n2915 VDD.n2811 9.3005
R5045 VDD.n2914 VDD.n2812 9.3005
R5046 VDD.n2911 VDD.n2813 9.3005
R5047 VDD.n2910 VDD.n2814 9.3005
R5048 VDD.n2907 VDD.n2815 9.3005
R5049 VDD.n2906 VDD.n2816 9.3005
R5050 VDD.n2903 VDD.n2817 9.3005
R5051 VDD.n2902 VDD.n2818 9.3005
R5052 VDD.n2899 VDD.n2819 9.3005
R5053 VDD.n2898 VDD.n2820 9.3005
R5054 VDD.n2895 VDD.n2894 9.3005
R5055 VDD.n2893 VDD.n2821 9.3005
R5056 VDD.n2892 VDD.n2891 9.3005
R5057 VDD.n2888 VDD.n2824 9.3005
R5058 VDD.n2885 VDD.n2825 9.3005
R5059 VDD.n2884 VDD.n2826 9.3005
R5060 VDD.n2881 VDD.n2827 9.3005
R5061 VDD.n2880 VDD.n2828 9.3005
R5062 VDD.n2877 VDD.n2829 9.3005
R5063 VDD.n2876 VDD.n2830 9.3005
R5064 VDD.n2873 VDD.n2831 9.3005
R5065 VDD.n2872 VDD.n2832 9.3005
R5066 VDD.n2869 VDD.n2833 9.3005
R5067 VDD.n2868 VDD.n2834 9.3005
R5068 VDD.n2865 VDD.n2835 9.3005
R5069 VDD.n2861 VDD.n2859 9.3005
R5070 VDD.n2950 VDD.n2794 9.3005
R5071 VDD.n2688 VDD.n2687 9.3005
R5072 VDD.n52 VDD.n51 9.3005
R5073 VDD.n2701 VDD.n2700 9.3005
R5074 VDD.n2702 VDD.n50 9.3005
R5075 VDD.n2704 VDD.n2703 9.3005
R5076 VDD.n40 VDD.n39 9.3005
R5077 VDD.n2717 VDD.n2716 9.3005
R5078 VDD.n2718 VDD.n38 9.3005
R5079 VDD.n2720 VDD.n2719 9.3005
R5080 VDD.n28 VDD.n27 9.3005
R5081 VDD.n2733 VDD.n2732 9.3005
R5082 VDD.n2734 VDD.n26 9.3005
R5083 VDD.n2980 VDD.n2735 9.3005
R5084 VDD.n2979 VDD.n2736 9.3005
R5085 VDD.n2978 VDD.n2737 9.3005
R5086 VDD.n2840 VDD.n2738 9.3005
R5087 VDD.n2842 VDD.n2841 9.3005
R5088 VDD.n2844 VDD.n2843 9.3005
R5089 VDD.n2845 VDD.n2839 9.3005
R5090 VDD.n2848 VDD.n2846 9.3005
R5091 VDD.n2849 VDD.n2838 9.3005
R5092 VDD.n2851 VDD.n2850 9.3005
R5093 VDD.n2852 VDD.n2837 9.3005
R5094 VDD.n2855 VDD.n2853 9.3005
R5095 VDD.n2856 VDD.n2836 9.3005
R5096 VDD.n2858 VDD.n2857 9.3005
R5097 VDD.n2686 VDD.n62 9.3005
R5098 VDD.n2685 VDD.n2684 9.3005
R5099 VDD.n2597 VDD.n63 9.3005
R5100 VDD.n2599 VDD.n2596 9.3005
R5101 VDD.n2600 VDD.n2595 9.3005
R5102 VDD.n2603 VDD.n2594 9.3005
R5103 VDD.n2605 VDD.n121 9.3005
R5104 VDD.n2613 VDD.n119 9.3005
R5105 VDD.n2614 VDD.n118 9.3005
R5106 VDD.n2617 VDD.n117 9.3005
R5107 VDD.n2621 VDD.n2620 9.3005
R5108 VDD.n2622 VDD.n114 9.3005
R5109 VDD.n1348 VDD.n1347 9.3005
R5110 VDD.n1346 VDD.n951 9.3005
R5111 VDD.n1345 VDD.n1344 9.3005
R5112 VDD.n1343 VDD.n963 9.3005
R5113 VDD.n1342 VDD.n1341 9.3005
R5114 VDD.n1337 VDD.n964 9.3005
R5115 VDD.n1041 VDD.n1040 9.3005
R5116 VDD.n1219 VDD.n1218 9.3005
R5117 VDD.n1220 VDD.n1039 9.3005
R5118 VDD.n1222 VDD.n1221 9.3005
R5119 VDD.n1030 VDD.n1029 9.3005
R5120 VDD.n1235 VDD.n1234 9.3005
R5121 VDD.n1236 VDD.n1028 9.3005
R5122 VDD.n1238 VDD.n1237 9.3005
R5123 VDD.n1018 VDD.n1017 9.3005
R5124 VDD.n1251 VDD.n1250 9.3005
R5125 VDD.n1252 VDD.n1016 9.3005
R5126 VDD.n1254 VDD.n1253 9.3005
R5127 VDD.n1007 VDD.n1006 9.3005
R5128 VDD.n1270 VDD.n1269 9.3005
R5129 VDD.n1271 VDD.n1005 9.3005
R5130 VDD.n1273 VDD.n1272 9.3005
R5131 VDD.n995 VDD.n994 9.3005
R5132 VDD.n1286 VDD.n1285 9.3005
R5133 VDD.n1287 VDD.n993 9.3005
R5134 VDD.n1289 VDD.n1288 9.3005
R5135 VDD.n983 VDD.n982 9.3005
R5136 VDD.n1302 VDD.n1301 9.3005
R5137 VDD.n1303 VDD.n980 9.3005
R5138 VDD.n1307 VDD.n1306 9.3005
R5139 VDD.n1305 VDD.n981 9.3005
R5140 VDD.n1304 VDD.n970 9.3005
R5141 VDD.n1206 VDD.n1205 9.3005
R5142 VDD.n1201 VDD.n1051 9.3005
R5143 VDD.n1193 VDD.n1054 9.3005
R5144 VDD.n1195 VDD.n1194 9.3005
R5145 VDD.n1192 VDD.n1056 9.3005
R5146 VDD.n1191 VDD.n1190 9.3005
R5147 VDD.n1058 VDD.n1057 9.3005
R5148 VDD.n1184 VDD.n1183 9.3005
R5149 VDD.n1182 VDD.n1060 9.3005
R5150 VDD.n1181 VDD.n1180 9.3005
R5151 VDD.n1062 VDD.n1061 9.3005
R5152 VDD.n1174 VDD.n1173 9.3005
R5153 VDD.n1172 VDD.n1064 9.3005
R5154 VDD.n1171 VDD.n1170 9.3005
R5155 VDD.n1066 VDD.n1065 9.3005
R5156 VDD.n1164 VDD.n1068 9.3005
R5157 VDD.n1163 VDD.n1162 9.3005
R5158 VDD.n1161 VDD.n1071 9.3005
R5159 VDD.n1160 VDD.n1159 9.3005
R5160 VDD.n1073 VDD.n1072 9.3005
R5161 VDD.n1150 VDD.n1076 9.3005
R5162 VDD.n1152 VDD.n1151 9.3005
R5163 VDD.n1149 VDD.n1078 9.3005
R5164 VDD.n1148 VDD.n1147 9.3005
R5165 VDD.n1080 VDD.n1079 9.3005
R5166 VDD.n1141 VDD.n1140 9.3005
R5167 VDD.n1139 VDD.n1082 9.3005
R5168 VDD.n1138 VDD.n1137 9.3005
R5169 VDD.n1084 VDD.n1083 9.3005
R5170 VDD.n1131 VDD.n1130 9.3005
R5171 VDD.n1129 VDD.n1088 9.3005
R5172 VDD.n1128 VDD.n1127 9.3005
R5173 VDD.n1090 VDD.n1089 9.3005
R5174 VDD.n1121 VDD.n1120 9.3005
R5175 VDD.n1119 VDD.n1092 9.3005
R5176 VDD.n1118 VDD.n1117 9.3005
R5177 VDD.n1094 VDD.n1093 9.3005
R5178 VDD.n1111 VDD.n1110 9.3005
R5179 VDD.n1109 VDD.n1096 9.3005
R5180 VDD.n1108 VDD.n1107 9.3005
R5181 VDD.n1098 VDD.n1097 9.3005
R5182 VDD.n1101 VDD.n1100 9.3005
R5183 VDD.n1099 VDD.n1047 9.3005
R5184 VDD.n1204 VDD.n1203 9.3005
R5185 VDD.n1212 VDD.n1046 9.3005
R5186 VDD.n1214 VDD.n1213 9.3005
R5187 VDD.n1036 VDD.n1035 9.3005
R5188 VDD.n1227 VDD.n1226 9.3005
R5189 VDD.n1228 VDD.n1034 9.3005
R5190 VDD.n1230 VDD.n1229 9.3005
R5191 VDD.n1024 VDD.n1023 9.3005
R5192 VDD.n1243 VDD.n1242 9.3005
R5193 VDD.n1244 VDD.n1022 9.3005
R5194 VDD.n1246 VDD.n1245 9.3005
R5195 VDD.n1012 VDD.n1011 9.3005
R5196 VDD.n1259 VDD.n1258 9.3005
R5197 VDD.n1211 VDD.n1210 9.3005
R5198 VDD.n1263 VDD.n1010 9.3005
R5199 VDD.n654 VDD.t97 8.78956
R5200 VDD.t82 VDD.n520 8.78956
R5201 VDD.n354 VDD.t96 8.78956
R5202 VDD.t87 VDD.n219 8.78956
R5203 VDD.n15 VDD.n14 8.2489
R5204 VDD.t49 VDD.t108 8.00831
R5205 VDD.t110 VDD.t59 8.00831
R5206 VDD.n1733 VDD.t116 7.813
R5207 VDD.n2356 VDD.t91 7.813
R5208 VDD.n1882 VDD.n445 7.18099
R5209 VDD.n1541 VDD.n1405 7.18099
R5210 VDD.n2220 VDD.n2087 7.18099
R5211 VDD.n155 VDD.n153 7.18099
R5212 VDD.n132 VDD.n130 7.18099
R5213 VDD.n1949 VDD.n1948 7.18099
R5214 VDD.n1838 VDD.n1837 7.18099
R5215 VDD.n938 VDD.n937 7.18099
R5216 VDD.n1631 VDD.t112 7.03175
R5217 VDD.n2458 VDD.t83 7.03175
R5218 VDD.n1164 VDD.n1163 6.98232
R5219 VDD.n1364 VDD.n778 6.98232
R5220 VDD.n2898 VDD.n2895 6.98232
R5221 VDD.n2627 VDD.n2624 6.98232
R5222 VDD.t112 VDD.n651 6.2505
R5223 VDD.n222 VDD.t83 6.2505
R5224 VDD.n1203 VDD.n1202 5.62474
R5225 VDD.n1340 VDD.n1337 5.62474
R5226 VDD.n2864 VDD.n2861 5.62474
R5227 VDD.n2684 VDD.n66 5.62474
R5228 VDD.t116 VDD.n550 5.46925
R5229 VDD.n324 VDD.t91 5.46925
R5230 VDD.n11 VDD.n9 4.99188
R5231 VDD.n4 VDD.n2 4.99188
R5232 VDD.n1351 VDD.n1350 4.74817
R5233 VDD.n955 VDD.n950 4.74817
R5234 VDD.n1401 VDD.n1400 4.74817
R5235 VDD.n1395 VDD.n741 4.74817
R5236 VDD.n1401 VDD.n742 4.74817
R5237 VDD.n746 VDD.n741 4.74817
R5238 VDD.n2669 VDD.n95 4.74817
R5239 VDD.n2662 VDD.n96 4.74817
R5240 VDD.n2665 VDD.n96 4.74817
R5241 VDD.n2666 VDD.n95 4.74817
R5242 VDD.n2609 VDD.n120 4.74817
R5243 VDD.n2607 VDD.n2606 4.74817
R5244 VDD.n2607 VDD.n2592 4.74817
R5245 VDD.n2610 VDD.n2609 4.74817
R5246 VDD.n1350 VDD.n790 4.74817
R5247 VDD.n952 VDD.n950 4.74817
R5248 VDD.n1263 VDD.n1262 4.64712
R5249 VDD.n2987 VDD.n2984 4.64712
R5250 VDD.n1643 VDD.t97 4.49269
R5251 VDD.n1763 VDD.t82 4.49269
R5252 VDD.n2326 VDD.t96 4.49269
R5253 VDD.n2446 VDD.t87 4.49269
R5254 VDD.n13 VDD.n11 3.97464
R5255 VDD.n6 VDD.n4 3.97464
R5256 VDD.n1819 VDD.t108 3.90675
R5257 VDD.n2272 VDD.t110 3.90675
R5258 VDD.n1262 VDD.n15 3.50649
R5259 VDD VDD.n2987 3.49866
R5260 VDD.n1885 VDD.n445 3.43465
R5261 VDD.n1544 VDD.n1405 3.43465
R5262 VDD.n2223 VDD.n2087 3.43465
R5263 VDD.n2545 VDD.n153 3.43465
R5264 VDD.n2580 VDD.n130 3.43465
R5265 VDD.n1948 VDD.n1947 3.43465
R5266 VDD.n1839 VDD.n1838 3.43465
R5267 VDD.n939 VDD.n938 3.43465
R5268 VDD.n2986 VDD.n2985 3.1061
R5269 VDD.n1261 VDD.n1260 3.1061
R5270 VDD.n14 VDD.n13 3.06233
R5271 VDD.n14 VDD.n6 3.06233
R5272 VDD.n612 VDD.t101 2.93019
R5273 VDD.t100 VDD.n562 2.93019
R5274 VDD.n312 VDD.t93 2.93019
R5275 VDD.t90 VDD.n262 2.93019
R5276 VDD.n1224 VDD.t45 2.73488
R5277 VDD.n1299 VDD.t16 2.73488
R5278 VDD.t8 VDD.n48 2.73488
R5279 VDD.n2961 VDD.t12 2.73488
R5280 VDD.n1402 VDD.n1401 2.27742
R5281 VDD.n1402 VDD.n741 2.27742
R5282 VDD.n2553 VDD.n96 2.27742
R5283 VDD.n2553 VDD.n95 2.27742
R5284 VDD.n2608 VDD.n2607 2.27742
R5285 VDD.n2609 VDD.n2608 2.27742
R5286 VDD.n1350 VDD.n1349 2.27742
R5287 VDD.n1349 VDD.n950 2.27742
R5288 VDD.n1775 VDD.t80 1.95362
R5289 VDD.n2314 VDD.t94 1.95362
R5290 VDD.n1262 VDD.n1261 1.39158
R5291 VDD.n2987 VDD.n2986 1.39157
R5292 VDD.n480 VDD.t49 1.36769
R5293 VDD.t59 VDD.n394 1.36769
R5294 VDD.t20 VDD.t106 0.977062
R5295 VDD.t104 VDD.t4 0.977062
R5296 VDD.n1202 VDD.n1201 0.970197
R5297 VDD.n1341 VDD.n1340 0.970197
R5298 VDD.n2865 VDD.n2864 0.970197
R5299 VDD.n2597 VDD.n66 0.970197
R5300 VDD.n1331 VDD.n1330 0.466963
R5301 VDD.n89 VDD.n57 0.466963
R5302 VDD.n2794 VDD.n2793 0.466963
R5303 VDD.n2859 VDD.n2858 0.466963
R5304 VDD.n2686 VDD.n2685 0.466963
R5305 VDD.n1304 VDD.n964 0.466963
R5306 VDD.n1205 VDD.n1204 0.466963
R5307 VDD.n1211 VDD.n1047 0.466963
R5308 VDD.t106 VDD.n694 0.391125
R5309 VDD.n600 VDD.t85 0.391125
R5310 VDD.t88 VDD.n274 0.391125
R5311 VDD.n180 VDD.t104 0.391125
R5312 VDD.n1264 VDD.n1000 0.152939
R5313 VDD.n1278 VDD.n1000 0.152939
R5314 VDD.n1279 VDD.n1278 0.152939
R5315 VDD.n1280 VDD.n1279 0.152939
R5316 VDD.n1280 VDD.n988 0.152939
R5317 VDD.n1294 VDD.n988 0.152939
R5318 VDD.n1295 VDD.n1294 0.152939
R5319 VDD.n1296 VDD.n1295 0.152939
R5320 VDD.n1296 VDD.n975 0.152939
R5321 VDD.n1312 VDD.n975 0.152939
R5322 VDD.n1313 VDD.n1312 0.152939
R5323 VDD.n1331 VDD.n1313 0.152939
R5324 VDD.n1330 VDD.n1314 0.152939
R5325 VDD.n1318 VDD.n1314 0.152939
R5326 VDD.n1319 VDD.n1318 0.152939
R5327 VDD.n1320 VDD.n1319 0.152939
R5328 VDD.n1320 VDD.n739 0.152939
R5329 VDD.n748 VDD.n740 0.152939
R5330 VDD.n1388 VDD.n748 0.152939
R5331 VDD.n1388 VDD.n1387 0.152939
R5332 VDD.n1387 VDD.n1386 0.152939
R5333 VDD.n1386 VDD.n754 0.152939
R5334 VDD.n759 VDD.n754 0.152939
R5335 VDD.n760 VDD.n759 0.152939
R5336 VDD.n761 VDD.n760 0.152939
R5337 VDD.n765 VDD.n761 0.152939
R5338 VDD.n766 VDD.n765 0.152939
R5339 VDD.n767 VDD.n766 0.152939
R5340 VDD.n768 VDD.n767 0.152939
R5341 VDD.n772 VDD.n768 0.152939
R5342 VDD.n773 VDD.n772 0.152939
R5343 VDD.n774 VDD.n773 0.152939
R5344 VDD.n775 VDD.n774 0.152939
R5345 VDD.n781 VDD.n775 0.152939
R5346 VDD.n782 VDD.n781 0.152939
R5347 VDD.n783 VDD.n782 0.152939
R5348 VDD.n784 VDD.n783 0.152939
R5349 VDD.n788 VDD.n784 0.152939
R5350 VDD.n789 VDD.n788 0.152939
R5351 VDD.n98 VDD.n97 0.152939
R5352 VDD.n2654 VDD.n98 0.152939
R5353 VDD.n2654 VDD.n2653 0.152939
R5354 VDD.n2653 VDD.n2652 0.152939
R5355 VDD.n2652 VDD.n102 0.152939
R5356 VDD.n103 VDD.n102 0.152939
R5357 VDD.n104 VDD.n103 0.152939
R5358 VDD.n105 VDD.n104 0.152939
R5359 VDD.n106 VDD.n105 0.152939
R5360 VDD.n107 VDD.n106 0.152939
R5361 VDD.n108 VDD.n107 0.152939
R5362 VDD.n109 VDD.n108 0.152939
R5363 VDD.n110 VDD.n109 0.152939
R5364 VDD.n111 VDD.n110 0.152939
R5365 VDD.n112 VDD.n111 0.152939
R5366 VDD.n113 VDD.n112 0.152939
R5367 VDD.n2623 VDD.n113 0.152939
R5368 VDD.n2623 VDD.n2622 0.152939
R5369 VDD.n2622 VDD.n2621 0.152939
R5370 VDD.n2621 VDD.n117 0.152939
R5371 VDD.n118 VDD.n117 0.152939
R5372 VDD.n119 VDD.n118 0.152939
R5373 VDD.n90 VDD.n89 0.152939
R5374 VDD.n91 VDD.n90 0.152939
R5375 VDD.n92 VDD.n91 0.152939
R5376 VDD.n93 VDD.n92 0.152939
R5377 VDD.n94 VDD.n93 0.152939
R5378 VDD.n2693 VDD.n57 0.152939
R5379 VDD.n2694 VDD.n2693 0.152939
R5380 VDD.n2695 VDD.n2694 0.152939
R5381 VDD.n2695 VDD.n45 0.152939
R5382 VDD.n2709 VDD.n45 0.152939
R5383 VDD.n2710 VDD.n2709 0.152939
R5384 VDD.n2711 VDD.n2710 0.152939
R5385 VDD.n2711 VDD.n33 0.152939
R5386 VDD.n2725 VDD.n33 0.152939
R5387 VDD.n2726 VDD.n2725 0.152939
R5388 VDD.n2727 VDD.n2726 0.152939
R5389 VDD.n2727 VDD.n16 0.152939
R5390 VDD.n2742 VDD.n17 0.152939
R5391 VDD.n2743 VDD.n2742 0.152939
R5392 VDD.n2744 VDD.n2743 0.152939
R5393 VDD.n2752 VDD.n2744 0.152939
R5394 VDD.n2753 VDD.n2752 0.152939
R5395 VDD.n2754 VDD.n2753 0.152939
R5396 VDD.n2755 VDD.n2754 0.152939
R5397 VDD.n2763 VDD.n2755 0.152939
R5398 VDD.n2764 VDD.n2763 0.152939
R5399 VDD.n2765 VDD.n2764 0.152939
R5400 VDD.n2766 VDD.n2765 0.152939
R5401 VDD.n2793 VDD.n2766 0.152939
R5402 VDD.n2948 VDD.n2794 0.152939
R5403 VDD.n2948 VDD.n2947 0.152939
R5404 VDD.n2947 VDD.n2946 0.152939
R5405 VDD.n2946 VDD.n2796 0.152939
R5406 VDD.n2797 VDD.n2796 0.152939
R5407 VDD.n2798 VDD.n2797 0.152939
R5408 VDD.n2799 VDD.n2798 0.152939
R5409 VDD.n2800 VDD.n2799 0.152939
R5410 VDD.n2801 VDD.n2800 0.152939
R5411 VDD.n2802 VDD.n2801 0.152939
R5412 VDD.n2803 VDD.n2802 0.152939
R5413 VDD.n2925 VDD.n2803 0.152939
R5414 VDD.n2925 VDD.n2924 0.152939
R5415 VDD.n2924 VDD.n2923 0.152939
R5416 VDD.n2923 VDD.n2809 0.152939
R5417 VDD.n2810 VDD.n2809 0.152939
R5418 VDD.n2811 VDD.n2810 0.152939
R5419 VDD.n2812 VDD.n2811 0.152939
R5420 VDD.n2813 VDD.n2812 0.152939
R5421 VDD.n2814 VDD.n2813 0.152939
R5422 VDD.n2815 VDD.n2814 0.152939
R5423 VDD.n2816 VDD.n2815 0.152939
R5424 VDD.n2817 VDD.n2816 0.152939
R5425 VDD.n2818 VDD.n2817 0.152939
R5426 VDD.n2819 VDD.n2818 0.152939
R5427 VDD.n2820 VDD.n2819 0.152939
R5428 VDD.n2894 VDD.n2820 0.152939
R5429 VDD.n2894 VDD.n2893 0.152939
R5430 VDD.n2893 VDD.n2892 0.152939
R5431 VDD.n2892 VDD.n2824 0.152939
R5432 VDD.n2825 VDD.n2824 0.152939
R5433 VDD.n2826 VDD.n2825 0.152939
R5434 VDD.n2827 VDD.n2826 0.152939
R5435 VDD.n2828 VDD.n2827 0.152939
R5436 VDD.n2829 VDD.n2828 0.152939
R5437 VDD.n2830 VDD.n2829 0.152939
R5438 VDD.n2831 VDD.n2830 0.152939
R5439 VDD.n2832 VDD.n2831 0.152939
R5440 VDD.n2833 VDD.n2832 0.152939
R5441 VDD.n2834 VDD.n2833 0.152939
R5442 VDD.n2835 VDD.n2834 0.152939
R5443 VDD.n2859 VDD.n2835 0.152939
R5444 VDD.n2687 VDD.n2686 0.152939
R5445 VDD.n2687 VDD.n51 0.152939
R5446 VDD.n2701 VDD.n51 0.152939
R5447 VDD.n2702 VDD.n2701 0.152939
R5448 VDD.n2703 VDD.n2702 0.152939
R5449 VDD.n2703 VDD.n39 0.152939
R5450 VDD.n2717 VDD.n39 0.152939
R5451 VDD.n2718 VDD.n2717 0.152939
R5452 VDD.n2719 VDD.n2718 0.152939
R5453 VDD.n2719 VDD.n27 0.152939
R5454 VDD.n2733 VDD.n27 0.152939
R5455 VDD.n2734 VDD.n2733 0.152939
R5456 VDD.n2735 VDD.n2734 0.152939
R5457 VDD.n2736 VDD.n2735 0.152939
R5458 VDD.n2737 VDD.n2736 0.152939
R5459 VDD.n2840 VDD.n2737 0.152939
R5460 VDD.n2841 VDD.n2840 0.152939
R5461 VDD.n2844 VDD.n2841 0.152939
R5462 VDD.n2845 VDD.n2844 0.152939
R5463 VDD.n2846 VDD.n2845 0.152939
R5464 VDD.n2846 VDD.n2838 0.152939
R5465 VDD.n2851 VDD.n2838 0.152939
R5466 VDD.n2852 VDD.n2851 0.152939
R5467 VDD.n2853 VDD.n2852 0.152939
R5468 VDD.n2853 VDD.n2836 0.152939
R5469 VDD.n2858 VDD.n2836 0.152939
R5470 VDD.n2594 VDD.n121 0.152939
R5471 VDD.n2595 VDD.n2594 0.152939
R5472 VDD.n2596 VDD.n2595 0.152939
R5473 VDD.n2596 VDD.n63 0.152939
R5474 VDD.n2685 VDD.n63 0.152939
R5475 VDD.n1348 VDD.n951 0.152939
R5476 VDD.n1344 VDD.n951 0.152939
R5477 VDD.n1344 VDD.n1343 0.152939
R5478 VDD.n1343 VDD.n1342 0.152939
R5479 VDD.n1342 VDD.n964 0.152939
R5480 VDD.n1205 VDD.n1040 0.152939
R5481 VDD.n1219 VDD.n1040 0.152939
R5482 VDD.n1220 VDD.n1219 0.152939
R5483 VDD.n1221 VDD.n1220 0.152939
R5484 VDD.n1221 VDD.n1029 0.152939
R5485 VDD.n1235 VDD.n1029 0.152939
R5486 VDD.n1236 VDD.n1235 0.152939
R5487 VDD.n1237 VDD.n1236 0.152939
R5488 VDD.n1237 VDD.n1017 0.152939
R5489 VDD.n1251 VDD.n1017 0.152939
R5490 VDD.n1252 VDD.n1251 0.152939
R5491 VDD.n1253 VDD.n1252 0.152939
R5492 VDD.n1253 VDD.n1006 0.152939
R5493 VDD.n1270 VDD.n1006 0.152939
R5494 VDD.n1271 VDD.n1270 0.152939
R5495 VDD.n1272 VDD.n1271 0.152939
R5496 VDD.n1272 VDD.n994 0.152939
R5497 VDD.n1286 VDD.n994 0.152939
R5498 VDD.n1287 VDD.n1286 0.152939
R5499 VDD.n1288 VDD.n1287 0.152939
R5500 VDD.n1288 VDD.n982 0.152939
R5501 VDD.n1302 VDD.n982 0.152939
R5502 VDD.n1303 VDD.n1302 0.152939
R5503 VDD.n1306 VDD.n1303 0.152939
R5504 VDD.n1306 VDD.n1305 0.152939
R5505 VDD.n1305 VDD.n1304 0.152939
R5506 VDD.n1100 VDD.n1047 0.152939
R5507 VDD.n1100 VDD.n1097 0.152939
R5508 VDD.n1108 VDD.n1097 0.152939
R5509 VDD.n1109 VDD.n1108 0.152939
R5510 VDD.n1110 VDD.n1109 0.152939
R5511 VDD.n1110 VDD.n1093 0.152939
R5512 VDD.n1118 VDD.n1093 0.152939
R5513 VDD.n1119 VDD.n1118 0.152939
R5514 VDD.n1120 VDD.n1119 0.152939
R5515 VDD.n1120 VDD.n1089 0.152939
R5516 VDD.n1128 VDD.n1089 0.152939
R5517 VDD.n1129 VDD.n1128 0.152939
R5518 VDD.n1130 VDD.n1129 0.152939
R5519 VDD.n1130 VDD.n1083 0.152939
R5520 VDD.n1138 VDD.n1083 0.152939
R5521 VDD.n1139 VDD.n1138 0.152939
R5522 VDD.n1140 VDD.n1139 0.152939
R5523 VDD.n1140 VDD.n1079 0.152939
R5524 VDD.n1148 VDD.n1079 0.152939
R5525 VDD.n1149 VDD.n1148 0.152939
R5526 VDD.n1151 VDD.n1149 0.152939
R5527 VDD.n1151 VDD.n1150 0.152939
R5528 VDD.n1150 VDD.n1072 0.152939
R5529 VDD.n1160 VDD.n1072 0.152939
R5530 VDD.n1161 VDD.n1160 0.152939
R5531 VDD.n1162 VDD.n1161 0.152939
R5532 VDD.n1162 VDD.n1068 0.152939
R5533 VDD.n1068 VDD.n1065 0.152939
R5534 VDD.n1171 VDD.n1065 0.152939
R5535 VDD.n1172 VDD.n1171 0.152939
R5536 VDD.n1173 VDD.n1172 0.152939
R5537 VDD.n1173 VDD.n1061 0.152939
R5538 VDD.n1181 VDD.n1061 0.152939
R5539 VDD.n1182 VDD.n1181 0.152939
R5540 VDD.n1183 VDD.n1182 0.152939
R5541 VDD.n1183 VDD.n1057 0.152939
R5542 VDD.n1191 VDD.n1057 0.152939
R5543 VDD.n1192 VDD.n1191 0.152939
R5544 VDD.n1194 VDD.n1192 0.152939
R5545 VDD.n1194 VDD.n1193 0.152939
R5546 VDD.n1193 VDD.n1051 0.152939
R5547 VDD.n1204 VDD.n1051 0.152939
R5548 VDD.n1212 VDD.n1211 0.152939
R5549 VDD.n1213 VDD.n1212 0.152939
R5550 VDD.n1213 VDD.n1035 0.152939
R5551 VDD.n1227 VDD.n1035 0.152939
R5552 VDD.n1228 VDD.n1227 0.152939
R5553 VDD.n1229 VDD.n1228 0.152939
R5554 VDD.n1229 VDD.n1023 0.152939
R5555 VDD.n1243 VDD.n1023 0.152939
R5556 VDD.n1244 VDD.n1243 0.152939
R5557 VDD.n1245 VDD.n1244 0.152939
R5558 VDD.n1245 VDD.n1011 0.152939
R5559 VDD.n1259 VDD.n1011 0.152939
R5560 VDD.n1402 VDD.n739 0.146841
R5561 VDD.n2553 VDD.n94 0.146841
R5562 VDD.n2608 VDD.n121 0.146841
R5563 VDD.n1349 VDD.n1348 0.146841
R5564 VDD.n1264 VDD.n1263 0.145814
R5565 VDD.n2984 VDD.n16 0.145814
R5566 VDD.n2984 VDD.n17 0.145814
R5567 VDD.n1263 VDD.n1259 0.145814
R5568 VDD VDD.n15 0.00833333
R5569 VDD.n1402 VDD.n740 0.00659756
R5570 VDD.n1349 VDD.n789 0.00659756
R5571 VDD.n2553 VDD.n97 0.00659756
R5572 VDD.n2608 VDD.n119 0.00659756
R5573 GND.n6188 GND.n6187 2282.54
R5574 GND.n5421 GND.n1234 2075.9
R5575 GND.n522 GND.n441 833.646
R5576 GND.n6351 GND.n450 833.646
R5577 GND.n4865 GND.n2542 833.646
R5578 GND.n4955 GND.n2550 833.646
R5579 GND.n5293 GND.n1401 833.646
R5580 GND.n5295 GND.n1394 833.646
R5581 GND.n1935 GND.n1276 833.646
R5582 GND.n5378 GND.n1280 833.646
R5583 GND.n3474 GND.n1533 778.39
R5584 GND.n4981 GND.n2498 778.39
R5585 GND.n4983 GND.n2493 778.39
R5586 GND.n5158 GND.n1535 778.39
R5587 GND.n4687 GND.n446 775.989
R5588 GND.n4706 GND.n451 775.989
R5589 GND.n2613 GND.n2544 775.989
R5590 GND.n4959 GND.n2518 775.989
R5591 GND.n5174 GND.n1399 775.989
R5592 GND.n5193 GND.n1396 775.989
R5593 GND.n1962 GND.n1277 775.989
R5594 GND.n1943 GND.n1279 775.989
R5595 GND.n5516 GND.n1138 775.989
R5596 GND.n6186 GND.n736 775.989
R5597 GND.n6312 GND.n664 775.989
R5598 GND.n5420 GND.n1235 775.989
R5599 GND.n5516 GND.n5515 585
R5600 GND.n5517 GND.n5516 585
R5601 GND.n5514 GND.n1140 585
R5602 GND.n1140 GND.n1139 585
R5603 GND.n5513 GND.n5512 585
R5604 GND.n5512 GND.n5511 585
R5605 GND.n1145 GND.n1144 585
R5606 GND.n5510 GND.n1145 585
R5607 GND.n5508 GND.n5507 585
R5608 GND.n5509 GND.n5508 585
R5609 GND.n5506 GND.n1147 585
R5610 GND.n1147 GND.n1146 585
R5611 GND.n5505 GND.n5504 585
R5612 GND.n5504 GND.n5503 585
R5613 GND.n1153 GND.n1152 585
R5614 GND.n5502 GND.n1153 585
R5615 GND.n5500 GND.n5499 585
R5616 GND.n5501 GND.n5500 585
R5617 GND.n5498 GND.n1155 585
R5618 GND.n1155 GND.n1154 585
R5619 GND.n5497 GND.n5496 585
R5620 GND.n5496 GND.n5495 585
R5621 GND.n1161 GND.n1160 585
R5622 GND.n5494 GND.n1161 585
R5623 GND.n5492 GND.n5491 585
R5624 GND.n5493 GND.n5492 585
R5625 GND.n5490 GND.n1163 585
R5626 GND.n1163 GND.n1162 585
R5627 GND.n5489 GND.n5488 585
R5628 GND.n5488 GND.n5487 585
R5629 GND.n1169 GND.n1168 585
R5630 GND.n5486 GND.n1169 585
R5631 GND.n5484 GND.n5483 585
R5632 GND.n5485 GND.n5484 585
R5633 GND.n5482 GND.n1171 585
R5634 GND.n1171 GND.n1170 585
R5635 GND.n5481 GND.n5480 585
R5636 GND.n5480 GND.n5479 585
R5637 GND.n1177 GND.n1176 585
R5638 GND.n5478 GND.n1177 585
R5639 GND.n5476 GND.n5475 585
R5640 GND.n5477 GND.n5476 585
R5641 GND.n5474 GND.n1179 585
R5642 GND.n1179 GND.n1178 585
R5643 GND.n5473 GND.n5472 585
R5644 GND.n5472 GND.n5471 585
R5645 GND.n1185 GND.n1184 585
R5646 GND.n5470 GND.n1185 585
R5647 GND.n5468 GND.n5467 585
R5648 GND.n5469 GND.n5468 585
R5649 GND.n5466 GND.n1187 585
R5650 GND.n1187 GND.n1186 585
R5651 GND.n5465 GND.n5464 585
R5652 GND.n5464 GND.n5463 585
R5653 GND.n1193 GND.n1192 585
R5654 GND.n5462 GND.n1193 585
R5655 GND.n5460 GND.n5459 585
R5656 GND.n5461 GND.n5460 585
R5657 GND.n5458 GND.n1195 585
R5658 GND.n1195 GND.n1194 585
R5659 GND.n5457 GND.n5456 585
R5660 GND.n5456 GND.n5455 585
R5661 GND.n1201 GND.n1200 585
R5662 GND.n5454 GND.n1201 585
R5663 GND.n5452 GND.n5451 585
R5664 GND.n5453 GND.n5452 585
R5665 GND.n5450 GND.n1203 585
R5666 GND.n1203 GND.n1202 585
R5667 GND.n5449 GND.n5448 585
R5668 GND.n5448 GND.n5447 585
R5669 GND.n1209 GND.n1208 585
R5670 GND.n5446 GND.n1209 585
R5671 GND.n5444 GND.n5443 585
R5672 GND.n5445 GND.n5444 585
R5673 GND.n5442 GND.n1211 585
R5674 GND.n1211 GND.n1210 585
R5675 GND.n5441 GND.n5440 585
R5676 GND.n5440 GND.n5439 585
R5677 GND.n1217 GND.n1216 585
R5678 GND.n5438 GND.n1217 585
R5679 GND.n5436 GND.n5435 585
R5680 GND.n5437 GND.n5436 585
R5681 GND.n5434 GND.n1219 585
R5682 GND.n1219 GND.n1218 585
R5683 GND.n5433 GND.n5432 585
R5684 GND.n5432 GND.n5431 585
R5685 GND.n1225 GND.n1224 585
R5686 GND.n5430 GND.n1225 585
R5687 GND.n5428 GND.n5427 585
R5688 GND.n5429 GND.n5428 585
R5689 GND.n5426 GND.n1227 585
R5690 GND.n1227 GND.n1226 585
R5691 GND.n5425 GND.n5424 585
R5692 GND.n5424 GND.n5423 585
R5693 GND.n1233 GND.n1232 585
R5694 GND.n5422 GND.n1233 585
R5695 GND.n5420 GND.n5419 585
R5696 GND.n5421 GND.n5420 585
R5697 GND.n1138 GND.n1137 585
R5698 GND.n5518 GND.n1138 585
R5699 GND.n5521 GND.n5520 585
R5700 GND.n5520 GND.n5519 585
R5701 GND.n1135 GND.n1134 585
R5702 GND.n1134 GND.n1133 585
R5703 GND.n5526 GND.n5525 585
R5704 GND.n5527 GND.n5526 585
R5705 GND.n1132 GND.n1131 585
R5706 GND.n5528 GND.n1132 585
R5707 GND.n5531 GND.n5530 585
R5708 GND.n5530 GND.n5529 585
R5709 GND.n1129 GND.n1128 585
R5710 GND.n1128 GND.n1127 585
R5711 GND.n5536 GND.n5535 585
R5712 GND.n5537 GND.n5536 585
R5713 GND.n1126 GND.n1125 585
R5714 GND.n5538 GND.n1126 585
R5715 GND.n5541 GND.n5540 585
R5716 GND.n5540 GND.n5539 585
R5717 GND.n1123 GND.n1122 585
R5718 GND.n1122 GND.n1121 585
R5719 GND.n5546 GND.n5545 585
R5720 GND.n5547 GND.n5546 585
R5721 GND.n1120 GND.n1119 585
R5722 GND.n5548 GND.n1120 585
R5723 GND.n5551 GND.n5550 585
R5724 GND.n5550 GND.n5549 585
R5725 GND.n1117 GND.n1116 585
R5726 GND.n1116 GND.n1115 585
R5727 GND.n5556 GND.n5555 585
R5728 GND.n5557 GND.n5556 585
R5729 GND.n1114 GND.n1113 585
R5730 GND.n5558 GND.n1114 585
R5731 GND.n5561 GND.n5560 585
R5732 GND.n5560 GND.n5559 585
R5733 GND.n1111 GND.n1110 585
R5734 GND.n1110 GND.n1109 585
R5735 GND.n5566 GND.n5565 585
R5736 GND.n5567 GND.n5566 585
R5737 GND.n1108 GND.n1107 585
R5738 GND.n5568 GND.n1108 585
R5739 GND.n5571 GND.n5570 585
R5740 GND.n5570 GND.n5569 585
R5741 GND.n1105 GND.n1104 585
R5742 GND.n1104 GND.n1103 585
R5743 GND.n5576 GND.n5575 585
R5744 GND.n5577 GND.n5576 585
R5745 GND.n1102 GND.n1101 585
R5746 GND.n5578 GND.n1102 585
R5747 GND.n5581 GND.n5580 585
R5748 GND.n5580 GND.n5579 585
R5749 GND.n1099 GND.n1098 585
R5750 GND.n1098 GND.n1097 585
R5751 GND.n5586 GND.n5585 585
R5752 GND.n5587 GND.n5586 585
R5753 GND.n1096 GND.n1095 585
R5754 GND.n5588 GND.n1096 585
R5755 GND.n5591 GND.n5590 585
R5756 GND.n5590 GND.n5589 585
R5757 GND.n1093 GND.n1092 585
R5758 GND.n1092 GND.n1091 585
R5759 GND.n5596 GND.n5595 585
R5760 GND.n5597 GND.n5596 585
R5761 GND.n1090 GND.n1089 585
R5762 GND.n5598 GND.n1090 585
R5763 GND.n5601 GND.n5600 585
R5764 GND.n5600 GND.n5599 585
R5765 GND.n1087 GND.n1086 585
R5766 GND.n1086 GND.n1085 585
R5767 GND.n5606 GND.n5605 585
R5768 GND.n5607 GND.n5606 585
R5769 GND.n1084 GND.n1083 585
R5770 GND.n5608 GND.n1084 585
R5771 GND.n5611 GND.n5610 585
R5772 GND.n5610 GND.n5609 585
R5773 GND.n1081 GND.n1080 585
R5774 GND.n1080 GND.n1079 585
R5775 GND.n5616 GND.n5615 585
R5776 GND.n5617 GND.n5616 585
R5777 GND.n1078 GND.n1077 585
R5778 GND.n5618 GND.n1078 585
R5779 GND.n5621 GND.n5620 585
R5780 GND.n5620 GND.n5619 585
R5781 GND.n1075 GND.n1074 585
R5782 GND.n1074 GND.n1073 585
R5783 GND.n5626 GND.n5625 585
R5784 GND.n5627 GND.n5626 585
R5785 GND.n1072 GND.n1071 585
R5786 GND.n5628 GND.n1072 585
R5787 GND.n5631 GND.n5630 585
R5788 GND.n5630 GND.n5629 585
R5789 GND.n1069 GND.n1068 585
R5790 GND.n1068 GND.n1067 585
R5791 GND.n5636 GND.n5635 585
R5792 GND.n5637 GND.n5636 585
R5793 GND.n1066 GND.n1065 585
R5794 GND.n5638 GND.n1066 585
R5795 GND.n5641 GND.n5640 585
R5796 GND.n5640 GND.n5639 585
R5797 GND.n1063 GND.n1062 585
R5798 GND.n1062 GND.n1061 585
R5799 GND.n5646 GND.n5645 585
R5800 GND.n5647 GND.n5646 585
R5801 GND.n1060 GND.n1059 585
R5802 GND.n5648 GND.n1060 585
R5803 GND.n5651 GND.n5650 585
R5804 GND.n5650 GND.n5649 585
R5805 GND.n1057 GND.n1056 585
R5806 GND.n1056 GND.n1055 585
R5807 GND.n5656 GND.n5655 585
R5808 GND.n5657 GND.n5656 585
R5809 GND.n1054 GND.n1053 585
R5810 GND.n5658 GND.n1054 585
R5811 GND.n5661 GND.n5660 585
R5812 GND.n5660 GND.n5659 585
R5813 GND.n1051 GND.n1050 585
R5814 GND.n1050 GND.n1049 585
R5815 GND.n5666 GND.n5665 585
R5816 GND.n5667 GND.n5666 585
R5817 GND.n1048 GND.n1047 585
R5818 GND.n5668 GND.n1048 585
R5819 GND.n5671 GND.n5670 585
R5820 GND.n5670 GND.n5669 585
R5821 GND.n1045 GND.n1044 585
R5822 GND.n1044 GND.n1043 585
R5823 GND.n5676 GND.n5675 585
R5824 GND.n5677 GND.n5676 585
R5825 GND.n1042 GND.n1041 585
R5826 GND.n5678 GND.n1042 585
R5827 GND.n5681 GND.n5680 585
R5828 GND.n5680 GND.n5679 585
R5829 GND.n1039 GND.n1038 585
R5830 GND.n1038 GND.n1037 585
R5831 GND.n5686 GND.n5685 585
R5832 GND.n5687 GND.n5686 585
R5833 GND.n1036 GND.n1035 585
R5834 GND.n5688 GND.n1036 585
R5835 GND.n5691 GND.n5690 585
R5836 GND.n5690 GND.n5689 585
R5837 GND.n1033 GND.n1032 585
R5838 GND.n1032 GND.n1031 585
R5839 GND.n5696 GND.n5695 585
R5840 GND.n5697 GND.n5696 585
R5841 GND.n1030 GND.n1029 585
R5842 GND.n5698 GND.n1030 585
R5843 GND.n5701 GND.n5700 585
R5844 GND.n5700 GND.n5699 585
R5845 GND.n1027 GND.n1026 585
R5846 GND.n1026 GND.n1025 585
R5847 GND.n5706 GND.n5705 585
R5848 GND.n5707 GND.n5706 585
R5849 GND.n1024 GND.n1023 585
R5850 GND.n5708 GND.n1024 585
R5851 GND.n5711 GND.n5710 585
R5852 GND.n5710 GND.n5709 585
R5853 GND.n1021 GND.n1020 585
R5854 GND.n1020 GND.n1019 585
R5855 GND.n5716 GND.n5715 585
R5856 GND.n5717 GND.n5716 585
R5857 GND.n1018 GND.n1017 585
R5858 GND.n5718 GND.n1018 585
R5859 GND.n5721 GND.n5720 585
R5860 GND.n5720 GND.n5719 585
R5861 GND.n1015 GND.n1014 585
R5862 GND.n1014 GND.n1013 585
R5863 GND.n5726 GND.n5725 585
R5864 GND.n5727 GND.n5726 585
R5865 GND.n1012 GND.n1011 585
R5866 GND.n5728 GND.n1012 585
R5867 GND.n5731 GND.n5730 585
R5868 GND.n5730 GND.n5729 585
R5869 GND.n1009 GND.n1008 585
R5870 GND.n1008 GND.n1007 585
R5871 GND.n5736 GND.n5735 585
R5872 GND.n5737 GND.n5736 585
R5873 GND.n1006 GND.n1005 585
R5874 GND.n5738 GND.n1006 585
R5875 GND.n5741 GND.n5740 585
R5876 GND.n5740 GND.n5739 585
R5877 GND.n1003 GND.n1002 585
R5878 GND.n1002 GND.n1001 585
R5879 GND.n5746 GND.n5745 585
R5880 GND.n5747 GND.n5746 585
R5881 GND.n1000 GND.n999 585
R5882 GND.n5748 GND.n1000 585
R5883 GND.n5751 GND.n5750 585
R5884 GND.n5750 GND.n5749 585
R5885 GND.n997 GND.n996 585
R5886 GND.n996 GND.n995 585
R5887 GND.n5756 GND.n5755 585
R5888 GND.n5757 GND.n5756 585
R5889 GND.n994 GND.n993 585
R5890 GND.n5758 GND.n994 585
R5891 GND.n5761 GND.n5760 585
R5892 GND.n5760 GND.n5759 585
R5893 GND.n991 GND.n990 585
R5894 GND.n990 GND.n989 585
R5895 GND.n5766 GND.n5765 585
R5896 GND.n5767 GND.n5766 585
R5897 GND.n988 GND.n987 585
R5898 GND.n5768 GND.n988 585
R5899 GND.n5771 GND.n5770 585
R5900 GND.n5770 GND.n5769 585
R5901 GND.n985 GND.n984 585
R5902 GND.n984 GND.n983 585
R5903 GND.n5776 GND.n5775 585
R5904 GND.n5777 GND.n5776 585
R5905 GND.n982 GND.n981 585
R5906 GND.n5778 GND.n982 585
R5907 GND.n5781 GND.n5780 585
R5908 GND.n5780 GND.n5779 585
R5909 GND.n979 GND.n978 585
R5910 GND.n978 GND.n977 585
R5911 GND.n5786 GND.n5785 585
R5912 GND.n5787 GND.n5786 585
R5913 GND.n976 GND.n975 585
R5914 GND.n5788 GND.n976 585
R5915 GND.n5791 GND.n5790 585
R5916 GND.n5790 GND.n5789 585
R5917 GND.n973 GND.n972 585
R5918 GND.n972 GND.n971 585
R5919 GND.n5796 GND.n5795 585
R5920 GND.n5797 GND.n5796 585
R5921 GND.n970 GND.n969 585
R5922 GND.n5798 GND.n970 585
R5923 GND.n5801 GND.n5800 585
R5924 GND.n5800 GND.n5799 585
R5925 GND.n967 GND.n966 585
R5926 GND.n966 GND.n965 585
R5927 GND.n5806 GND.n5805 585
R5928 GND.n5807 GND.n5806 585
R5929 GND.n964 GND.n963 585
R5930 GND.n5808 GND.n964 585
R5931 GND.n5811 GND.n5810 585
R5932 GND.n5810 GND.n5809 585
R5933 GND.n961 GND.n960 585
R5934 GND.n960 GND.n959 585
R5935 GND.n5816 GND.n5815 585
R5936 GND.n5817 GND.n5816 585
R5937 GND.n958 GND.n957 585
R5938 GND.n5818 GND.n958 585
R5939 GND.n5821 GND.n5820 585
R5940 GND.n5820 GND.n5819 585
R5941 GND.n955 GND.n954 585
R5942 GND.n954 GND.n953 585
R5943 GND.n5826 GND.n5825 585
R5944 GND.n5827 GND.n5826 585
R5945 GND.n952 GND.n951 585
R5946 GND.n5828 GND.n952 585
R5947 GND.n5831 GND.n5830 585
R5948 GND.n5830 GND.n5829 585
R5949 GND.n949 GND.n948 585
R5950 GND.n948 GND.n947 585
R5951 GND.n5836 GND.n5835 585
R5952 GND.n5837 GND.n5836 585
R5953 GND.n946 GND.n945 585
R5954 GND.n5838 GND.n946 585
R5955 GND.n5841 GND.n5840 585
R5956 GND.n5840 GND.n5839 585
R5957 GND.n943 GND.n942 585
R5958 GND.n942 GND.n941 585
R5959 GND.n5846 GND.n5845 585
R5960 GND.n5847 GND.n5846 585
R5961 GND.n940 GND.n939 585
R5962 GND.n5848 GND.n940 585
R5963 GND.n5851 GND.n5850 585
R5964 GND.n5850 GND.n5849 585
R5965 GND.n937 GND.n936 585
R5966 GND.n936 GND.n935 585
R5967 GND.n5856 GND.n5855 585
R5968 GND.n5857 GND.n5856 585
R5969 GND.n934 GND.n933 585
R5970 GND.n5858 GND.n934 585
R5971 GND.n5861 GND.n5860 585
R5972 GND.n5860 GND.n5859 585
R5973 GND.n931 GND.n930 585
R5974 GND.n930 GND.n929 585
R5975 GND.n5866 GND.n5865 585
R5976 GND.n5867 GND.n5866 585
R5977 GND.n928 GND.n927 585
R5978 GND.n5868 GND.n928 585
R5979 GND.n5871 GND.n5870 585
R5980 GND.n5870 GND.n5869 585
R5981 GND.n925 GND.n924 585
R5982 GND.n924 GND.n923 585
R5983 GND.n5876 GND.n5875 585
R5984 GND.n5877 GND.n5876 585
R5985 GND.n922 GND.n921 585
R5986 GND.n5878 GND.n922 585
R5987 GND.n5881 GND.n5880 585
R5988 GND.n5880 GND.n5879 585
R5989 GND.n919 GND.n918 585
R5990 GND.n918 GND.n917 585
R5991 GND.n5886 GND.n5885 585
R5992 GND.n5887 GND.n5886 585
R5993 GND.n916 GND.n915 585
R5994 GND.n5888 GND.n916 585
R5995 GND.n5891 GND.n5890 585
R5996 GND.n5890 GND.n5889 585
R5997 GND.n913 GND.n912 585
R5998 GND.n912 GND.n911 585
R5999 GND.n5896 GND.n5895 585
R6000 GND.n5897 GND.n5896 585
R6001 GND.n910 GND.n909 585
R6002 GND.n5898 GND.n910 585
R6003 GND.n5901 GND.n5900 585
R6004 GND.n5900 GND.n5899 585
R6005 GND.n907 GND.n906 585
R6006 GND.n906 GND.n905 585
R6007 GND.n5906 GND.n5905 585
R6008 GND.n5907 GND.n5906 585
R6009 GND.n904 GND.n903 585
R6010 GND.n5908 GND.n904 585
R6011 GND.n5911 GND.n5910 585
R6012 GND.n5910 GND.n5909 585
R6013 GND.n901 GND.n900 585
R6014 GND.n900 GND.n899 585
R6015 GND.n5916 GND.n5915 585
R6016 GND.n5917 GND.n5916 585
R6017 GND.n898 GND.n897 585
R6018 GND.n5918 GND.n898 585
R6019 GND.n5921 GND.n5920 585
R6020 GND.n5920 GND.n5919 585
R6021 GND.n895 GND.n894 585
R6022 GND.n894 GND.n893 585
R6023 GND.n5926 GND.n5925 585
R6024 GND.n5927 GND.n5926 585
R6025 GND.n892 GND.n891 585
R6026 GND.n5928 GND.n892 585
R6027 GND.n5931 GND.n5930 585
R6028 GND.n5930 GND.n5929 585
R6029 GND.n889 GND.n888 585
R6030 GND.n888 GND.n887 585
R6031 GND.n5936 GND.n5935 585
R6032 GND.n5937 GND.n5936 585
R6033 GND.n886 GND.n885 585
R6034 GND.n5938 GND.n886 585
R6035 GND.n5941 GND.n5940 585
R6036 GND.n5940 GND.n5939 585
R6037 GND.n883 GND.n882 585
R6038 GND.n882 GND.n881 585
R6039 GND.n5946 GND.n5945 585
R6040 GND.n5947 GND.n5946 585
R6041 GND.n880 GND.n879 585
R6042 GND.n5948 GND.n880 585
R6043 GND.n5951 GND.n5950 585
R6044 GND.n5950 GND.n5949 585
R6045 GND.n877 GND.n876 585
R6046 GND.n876 GND.n875 585
R6047 GND.n5956 GND.n5955 585
R6048 GND.n5957 GND.n5956 585
R6049 GND.n874 GND.n873 585
R6050 GND.n5958 GND.n874 585
R6051 GND.n5961 GND.n5960 585
R6052 GND.n5960 GND.n5959 585
R6053 GND.n871 GND.n870 585
R6054 GND.n870 GND.n869 585
R6055 GND.n5966 GND.n5965 585
R6056 GND.n5967 GND.n5966 585
R6057 GND.n868 GND.n867 585
R6058 GND.n5968 GND.n868 585
R6059 GND.n5971 GND.n5970 585
R6060 GND.n5970 GND.n5969 585
R6061 GND.n865 GND.n864 585
R6062 GND.n864 GND.n863 585
R6063 GND.n5976 GND.n5975 585
R6064 GND.n5977 GND.n5976 585
R6065 GND.n862 GND.n861 585
R6066 GND.n5978 GND.n862 585
R6067 GND.n5981 GND.n5980 585
R6068 GND.n5980 GND.n5979 585
R6069 GND.n859 GND.n858 585
R6070 GND.n858 GND.n857 585
R6071 GND.n5986 GND.n5985 585
R6072 GND.n5987 GND.n5986 585
R6073 GND.n856 GND.n855 585
R6074 GND.n5988 GND.n856 585
R6075 GND.n5991 GND.n5990 585
R6076 GND.n5990 GND.n5989 585
R6077 GND.n853 GND.n852 585
R6078 GND.n852 GND.n851 585
R6079 GND.n5996 GND.n5995 585
R6080 GND.n5997 GND.n5996 585
R6081 GND.n850 GND.n849 585
R6082 GND.n5998 GND.n850 585
R6083 GND.n6001 GND.n6000 585
R6084 GND.n6000 GND.n5999 585
R6085 GND.n847 GND.n846 585
R6086 GND.n846 GND.n845 585
R6087 GND.n6006 GND.n6005 585
R6088 GND.n6007 GND.n6006 585
R6089 GND.n844 GND.n843 585
R6090 GND.n6008 GND.n844 585
R6091 GND.n6011 GND.n6010 585
R6092 GND.n6010 GND.n6009 585
R6093 GND.n841 GND.n840 585
R6094 GND.n840 GND.n839 585
R6095 GND.n6016 GND.n6015 585
R6096 GND.n6017 GND.n6016 585
R6097 GND.n838 GND.n837 585
R6098 GND.n6018 GND.n838 585
R6099 GND.n6021 GND.n6020 585
R6100 GND.n6020 GND.n6019 585
R6101 GND.n835 GND.n834 585
R6102 GND.n834 GND.n833 585
R6103 GND.n6026 GND.n6025 585
R6104 GND.n6027 GND.n6026 585
R6105 GND.n832 GND.n831 585
R6106 GND.n6028 GND.n832 585
R6107 GND.n6031 GND.n6030 585
R6108 GND.n6030 GND.n6029 585
R6109 GND.n829 GND.n828 585
R6110 GND.n828 GND.n827 585
R6111 GND.n6036 GND.n6035 585
R6112 GND.n6037 GND.n6036 585
R6113 GND.n826 GND.n825 585
R6114 GND.n6038 GND.n826 585
R6115 GND.n6041 GND.n6040 585
R6116 GND.n6040 GND.n6039 585
R6117 GND.n823 GND.n822 585
R6118 GND.n822 GND.n821 585
R6119 GND.n6046 GND.n6045 585
R6120 GND.n6047 GND.n6046 585
R6121 GND.n820 GND.n819 585
R6122 GND.n6048 GND.n820 585
R6123 GND.n6051 GND.n6050 585
R6124 GND.n6050 GND.n6049 585
R6125 GND.n817 GND.n816 585
R6126 GND.n816 GND.n815 585
R6127 GND.n6056 GND.n6055 585
R6128 GND.n6057 GND.n6056 585
R6129 GND.n814 GND.n813 585
R6130 GND.n6058 GND.n814 585
R6131 GND.n6061 GND.n6060 585
R6132 GND.n6060 GND.n6059 585
R6133 GND.n811 GND.n810 585
R6134 GND.n810 GND.n809 585
R6135 GND.n6066 GND.n6065 585
R6136 GND.n6067 GND.n6066 585
R6137 GND.n808 GND.n807 585
R6138 GND.n6068 GND.n808 585
R6139 GND.n6071 GND.n6070 585
R6140 GND.n6070 GND.n6069 585
R6141 GND.n805 GND.n804 585
R6142 GND.n804 GND.n803 585
R6143 GND.n6076 GND.n6075 585
R6144 GND.n6077 GND.n6076 585
R6145 GND.n802 GND.n801 585
R6146 GND.n6078 GND.n802 585
R6147 GND.n6081 GND.n6080 585
R6148 GND.n6080 GND.n6079 585
R6149 GND.n799 GND.n798 585
R6150 GND.n798 GND.n797 585
R6151 GND.n6086 GND.n6085 585
R6152 GND.n6087 GND.n6086 585
R6153 GND.n796 GND.n795 585
R6154 GND.n6088 GND.n796 585
R6155 GND.n6091 GND.n6090 585
R6156 GND.n6090 GND.n6089 585
R6157 GND.n793 GND.n792 585
R6158 GND.n792 GND.n791 585
R6159 GND.n6096 GND.n6095 585
R6160 GND.n6097 GND.n6096 585
R6161 GND.n790 GND.n789 585
R6162 GND.n6098 GND.n790 585
R6163 GND.n6101 GND.n6100 585
R6164 GND.n6100 GND.n6099 585
R6165 GND.n787 GND.n786 585
R6166 GND.n786 GND.n785 585
R6167 GND.n6106 GND.n6105 585
R6168 GND.n6107 GND.n6106 585
R6169 GND.n784 GND.n783 585
R6170 GND.n6108 GND.n784 585
R6171 GND.n6111 GND.n6110 585
R6172 GND.n6110 GND.n6109 585
R6173 GND.n781 GND.n780 585
R6174 GND.n780 GND.n779 585
R6175 GND.n6116 GND.n6115 585
R6176 GND.n6117 GND.n6116 585
R6177 GND.n778 GND.n777 585
R6178 GND.n6118 GND.n778 585
R6179 GND.n6121 GND.n6120 585
R6180 GND.n6120 GND.n6119 585
R6181 GND.n775 GND.n774 585
R6182 GND.n774 GND.n773 585
R6183 GND.n6126 GND.n6125 585
R6184 GND.n6127 GND.n6126 585
R6185 GND.n772 GND.n771 585
R6186 GND.n6128 GND.n772 585
R6187 GND.n6131 GND.n6130 585
R6188 GND.n6130 GND.n6129 585
R6189 GND.n769 GND.n768 585
R6190 GND.n768 GND.n767 585
R6191 GND.n6136 GND.n6135 585
R6192 GND.n6137 GND.n6136 585
R6193 GND.n766 GND.n765 585
R6194 GND.n6138 GND.n766 585
R6195 GND.n6141 GND.n6140 585
R6196 GND.n6140 GND.n6139 585
R6197 GND.n763 GND.n762 585
R6198 GND.n762 GND.n761 585
R6199 GND.n6146 GND.n6145 585
R6200 GND.n6147 GND.n6146 585
R6201 GND.n760 GND.n759 585
R6202 GND.n6148 GND.n760 585
R6203 GND.n6151 GND.n6150 585
R6204 GND.n6150 GND.n6149 585
R6205 GND.n757 GND.n756 585
R6206 GND.n756 GND.n755 585
R6207 GND.n6156 GND.n6155 585
R6208 GND.n6157 GND.n6156 585
R6209 GND.n754 GND.n753 585
R6210 GND.n6158 GND.n754 585
R6211 GND.n6161 GND.n6160 585
R6212 GND.n6160 GND.n6159 585
R6213 GND.n751 GND.n750 585
R6214 GND.n750 GND.n749 585
R6215 GND.n6166 GND.n6165 585
R6216 GND.n6167 GND.n6166 585
R6217 GND.n748 GND.n747 585
R6218 GND.n6168 GND.n748 585
R6219 GND.n6171 GND.n6170 585
R6220 GND.n6170 GND.n6169 585
R6221 GND.n745 GND.n744 585
R6222 GND.n744 GND.n743 585
R6223 GND.n6176 GND.n6175 585
R6224 GND.n6177 GND.n6176 585
R6225 GND.n742 GND.n741 585
R6226 GND.n6178 GND.n742 585
R6227 GND.n6181 GND.n6180 585
R6228 GND.n6180 GND.n6179 585
R6229 GND.n739 GND.n738 585
R6230 GND.n738 GND.n737 585
R6231 GND.n6186 GND.n6185 585
R6232 GND.n6187 GND.n6186 585
R6233 GND.n6306 GND.n664 585
R6234 GND.n6310 GND.n664 585
R6235 GND.n6308 GND.n6307 585
R6236 GND.n6309 GND.n6308 585
R6237 GND.n667 GND.n666 585
R6238 GND.n666 GND.n665 585
R6239 GND.n6301 GND.n6300 585
R6240 GND.n6300 GND.n6299 585
R6241 GND.n670 GND.n669 585
R6242 GND.n6298 GND.n670 585
R6243 GND.n6296 GND.n6295 585
R6244 GND.n6297 GND.n6296 585
R6245 GND.n673 GND.n672 585
R6246 GND.n672 GND.n671 585
R6247 GND.n6291 GND.n6290 585
R6248 GND.n6290 GND.n6289 585
R6249 GND.n676 GND.n675 585
R6250 GND.n6288 GND.n676 585
R6251 GND.n6286 GND.n6285 585
R6252 GND.n6287 GND.n6286 585
R6253 GND.n679 GND.n678 585
R6254 GND.n678 GND.n677 585
R6255 GND.n6281 GND.n6280 585
R6256 GND.n6280 GND.n6279 585
R6257 GND.n682 GND.n681 585
R6258 GND.n6278 GND.n682 585
R6259 GND.n6276 GND.n6275 585
R6260 GND.n6277 GND.n6276 585
R6261 GND.n685 GND.n684 585
R6262 GND.n684 GND.n683 585
R6263 GND.n6271 GND.n6270 585
R6264 GND.n6270 GND.n6269 585
R6265 GND.n688 GND.n687 585
R6266 GND.n6268 GND.n688 585
R6267 GND.n6266 GND.n6265 585
R6268 GND.n6267 GND.n6266 585
R6269 GND.n691 GND.n690 585
R6270 GND.n690 GND.n689 585
R6271 GND.n6261 GND.n6260 585
R6272 GND.n6260 GND.n6259 585
R6273 GND.n694 GND.n693 585
R6274 GND.n6258 GND.n694 585
R6275 GND.n6256 GND.n6255 585
R6276 GND.n6257 GND.n6256 585
R6277 GND.n697 GND.n696 585
R6278 GND.n696 GND.n695 585
R6279 GND.n6251 GND.n6250 585
R6280 GND.n6250 GND.n6249 585
R6281 GND.n700 GND.n699 585
R6282 GND.n6248 GND.n700 585
R6283 GND.n6246 GND.n6245 585
R6284 GND.n6247 GND.n6246 585
R6285 GND.n703 GND.n702 585
R6286 GND.n702 GND.n701 585
R6287 GND.n6241 GND.n6240 585
R6288 GND.n6240 GND.n6239 585
R6289 GND.n706 GND.n705 585
R6290 GND.n6238 GND.n706 585
R6291 GND.n6236 GND.n6235 585
R6292 GND.n6237 GND.n6236 585
R6293 GND.n709 GND.n708 585
R6294 GND.n708 GND.n707 585
R6295 GND.n6231 GND.n6230 585
R6296 GND.n6230 GND.n6229 585
R6297 GND.n712 GND.n711 585
R6298 GND.n6228 GND.n712 585
R6299 GND.n6226 GND.n6225 585
R6300 GND.n6227 GND.n6226 585
R6301 GND.n715 GND.n714 585
R6302 GND.n714 GND.n713 585
R6303 GND.n6221 GND.n6220 585
R6304 GND.n6220 GND.n6219 585
R6305 GND.n718 GND.n717 585
R6306 GND.n6218 GND.n718 585
R6307 GND.n6216 GND.n6215 585
R6308 GND.n6217 GND.n6216 585
R6309 GND.n721 GND.n720 585
R6310 GND.n720 GND.n719 585
R6311 GND.n6211 GND.n6210 585
R6312 GND.n6210 GND.n6209 585
R6313 GND.n724 GND.n723 585
R6314 GND.n6208 GND.n724 585
R6315 GND.n6206 GND.n6205 585
R6316 GND.n6207 GND.n6206 585
R6317 GND.n727 GND.n726 585
R6318 GND.n726 GND.n725 585
R6319 GND.n6201 GND.n6200 585
R6320 GND.n6200 GND.n6199 585
R6321 GND.n730 GND.n729 585
R6322 GND.n6198 GND.n730 585
R6323 GND.n6196 GND.n6195 585
R6324 GND.n6197 GND.n6196 585
R6325 GND.n733 GND.n732 585
R6326 GND.n732 GND.n731 585
R6327 GND.n6191 GND.n6190 585
R6328 GND.n6190 GND.n6189 585
R6329 GND.n736 GND.n735 585
R6330 GND.n6188 GND.n736 585
R6331 GND.n1399 GND.n1398 585
R6332 GND.n5294 GND.n1399 585
R6333 GND.n2344 GND.n1391 585
R6334 GND.n2345 GND.n2344 585
R6335 GND.n2343 GND.n1390 585
R6336 GND.n2343 GND.n2342 585
R6337 GND.n1542 GND.n1389 585
R6338 GND.n2278 GND.n1542 585
R6339 GND.n2333 GND.n2332 585
R6340 GND.n2334 GND.n2333 585
R6341 GND.n2331 GND.n1383 585
R6342 GND.n2331 GND.n2330 585
R6343 GND.n1552 GND.n1382 585
R6344 GND.n2305 GND.n1552 585
R6345 GND.n2294 GND.n1381 585
R6346 GND.n2294 GND.n1561 585
R6347 GND.n2296 GND.n2295 585
R6348 GND.n2297 GND.n2296 585
R6349 GND.n2293 GND.n1375 585
R6350 GND.n2293 GND.n2292 585
R6351 GND.n1572 GND.n1374 585
R6352 GND.n1585 GND.n1572 585
R6353 GND.n1582 GND.n1373 585
R6354 GND.n2269 GND.n1582 585
R6355 GND.n2257 GND.n2255 585
R6356 GND.n2257 GND.n2256 585
R6357 GND.n2258 GND.n1367 585
R6358 GND.n2259 GND.n2258 585
R6359 GND.n2254 GND.n1366 585
R6360 GND.n2254 GND.n2253 585
R6361 GND.n1594 GND.n1365 585
R6362 GND.n1608 GND.n1594 585
R6363 GND.n1606 GND.n1605 585
R6364 GND.n2244 GND.n1606 585
R6365 GND.n2232 GND.n1359 585
R6366 GND.n2232 GND.n2231 585
R6367 GND.n2233 GND.n1358 585
R6368 GND.n2234 GND.n2233 585
R6369 GND.n2230 GND.n1357 585
R6370 GND.n2230 GND.n2229 585
R6371 GND.n1619 GND.n1618 585
R6372 GND.n1631 GND.n1619 585
R6373 GND.n1629 GND.n1351 585
R6374 GND.n2220 GND.n1629 585
R6375 GND.n2139 GND.n1350 585
R6376 GND.n2140 GND.n2139 585
R6377 GND.n1671 GND.n1349 585
R6378 GND.n2136 GND.n1671 585
R6379 GND.n2192 GND.n1672 585
R6380 GND.n2192 GND.n2191 585
R6381 GND.n2193 GND.n1343 585
R6382 GND.n2194 GND.n2193 585
R6383 GND.n1664 GND.n1342 585
R6384 GND.n2199 GND.n1664 585
R6385 GND.n1663 GND.n1341 585
R6386 GND.n1663 GND.n1659 585
R6387 GND.n1650 GND.n1649 585
R6388 GND.n1652 GND.n1650 585
R6389 GND.n2209 GND.n1335 585
R6390 GND.n2209 GND.n2208 585
R6391 GND.n2210 GND.n1334 585
R6392 GND.n2211 GND.n2210 585
R6393 GND.n1648 GND.n1333 585
R6394 GND.n1684 GND.n1648 585
R6395 GND.n1687 GND.n1686 585
R6396 GND.n2112 GND.n1687 585
R6397 GND.n2102 GND.n1327 585
R6398 GND.n2102 GND.n2101 585
R6399 GND.n2103 GND.n1326 585
R6400 GND.n2104 GND.n2103 585
R6401 GND.n2100 GND.n1325 585
R6402 GND.n2100 GND.n2099 585
R6403 GND.n1698 GND.n1697 585
R6404 GND.n1709 GND.n1698 585
R6405 GND.n1707 GND.n1319 585
R6406 GND.n2090 GND.n1707 585
R6407 GND.n2078 GND.n1318 585
R6408 GND.n2078 GND.n2077 585
R6409 GND.n2079 GND.n1317 585
R6410 GND.n2080 GND.n2079 585
R6411 GND.n1719 GND.n1718 585
R6412 GND.n2046 GND.n1719 585
R6413 GND.n1737 GND.n1311 585
R6414 GND.n1737 GND.n1727 585
R6415 GND.n1738 GND.n1310 585
R6416 GND.n2037 GND.n1738 585
R6417 GND.n2024 GND.n1309 585
R6418 GND.n2024 GND.n2023 585
R6419 GND.n2026 GND.n2025 585
R6420 GND.n2027 GND.n2026 585
R6421 GND.n2022 GND.n1303 585
R6422 GND.n2022 GND.n2021 585
R6423 GND.n1748 GND.n1302 585
R6424 GND.n2004 GND.n1748 585
R6425 GND.n1974 GND.n1301 585
R6426 GND.n2012 GND.n1974 585
R6427 GND.n1294 GND.n1292 585
R6428 GND.n1972 GND.n1292 585
R6429 GND.n5372 GND.n5371 585
R6430 GND.n5373 GND.n5372 585
R6431 GND.n1293 GND.n1291 585
R6432 GND.n1755 GND.n1291 585
R6433 GND.n1938 GND.n1279 585
R6434 GND.n5379 GND.n1279 585
R6435 GND.n1944 GND.n1943 585
R6436 GND.n1767 GND.n1766 585
R6437 GND.n1949 GND.n1948 585
R6438 GND.n1951 GND.n1765 585
R6439 GND.n1954 GND.n1953 585
R6440 GND.n1763 GND.n1762 585
R6441 GND.n1959 GND.n1958 585
R6442 GND.n1961 GND.n1761 585
R6443 GND.n1963 GND.n1962 585
R6444 GND.n1962 GND.n1267 585
R6445 GND.n5194 GND.n5193 585
R6446 GND.n1504 GND.n1503 585
R6447 GND.n5169 GND.n1488 585
R6448 GND.n5207 GND.n1487 585
R6449 GND.n5208 GND.n1486 585
R6450 GND.n5171 GND.n1480 585
R6451 GND.n5215 GND.n1479 585
R6452 GND.n5216 GND.n1478 585
R6453 GND.n5174 GND.n1477 585
R6454 GND.n5191 GND.n5174 585
R6455 GND.n2348 GND.n1396 585
R6456 GND.n5294 GND.n1396 585
R6457 GND.n2347 GND.n2346 585
R6458 GND.n2346 GND.n2345 585
R6459 GND.n1540 GND.n1539 585
R6460 GND.n2342 GND.n1540 585
R6461 GND.n2280 GND.n2279 585
R6462 GND.n2279 GND.n2278 585
R6463 GND.n2276 GND.n1550 585
R6464 GND.n2334 GND.n1550 585
R6465 GND.n2284 GND.n1554 585
R6466 GND.n2330 GND.n1554 585
R6467 GND.n2285 GND.n1563 585
R6468 GND.n2305 GND.n1563 585
R6469 GND.n2286 GND.n2275 585
R6470 GND.n2275 GND.n1561 585
R6471 GND.n1576 GND.n1570 585
R6472 GND.n2297 GND.n1570 585
R6473 GND.n2291 GND.n2290 585
R6474 GND.n2292 GND.n2291 585
R6475 GND.n1575 GND.n1574 585
R6476 GND.n1585 GND.n1574 585
R6477 GND.n2271 GND.n2270 585
R6478 GND.n2270 GND.n2269 585
R6479 GND.n1579 GND.n1578 585
R6480 GND.n2256 GND.n1579 585
R6481 GND.n1599 GND.n1592 585
R6482 GND.n2259 GND.n1592 585
R6483 GND.n2252 GND.n2251 585
R6484 GND.n2253 GND.n2252 585
R6485 GND.n1598 GND.n1597 585
R6486 GND.n1608 GND.n1597 585
R6487 GND.n2246 GND.n2245 585
R6488 GND.n2245 GND.n2244 585
R6489 GND.n1602 GND.n1601 585
R6490 GND.n2231 GND.n1602 585
R6491 GND.n1623 GND.n1616 585
R6492 GND.n2234 GND.n1616 585
R6493 GND.n2228 GND.n2227 585
R6494 GND.n2229 GND.n2228 585
R6495 GND.n1622 GND.n1621 585
R6496 GND.n1631 GND.n1621 585
R6497 GND.n2222 GND.n2221 585
R6498 GND.n2221 GND.n2220 585
R6499 GND.n1626 GND.n1625 585
R6500 GND.n2140 GND.n1626 585
R6501 GND.n2132 GND.n2131 585
R6502 GND.n2136 GND.n2132 585
R6503 GND.n1674 GND.n1673 585
R6504 GND.n2191 GND.n1673 585
R6505 GND.n2127 GND.n1669 585
R6506 GND.n2194 GND.n1669 585
R6507 GND.n2126 GND.n1661 585
R6508 GND.n2199 GND.n1661 585
R6509 GND.n2120 GND.n1676 585
R6510 GND.n2120 GND.n1659 585
R6511 GND.n2122 GND.n2121 585
R6512 GND.n2121 GND.n1652 585
R6513 GND.n2119 GND.n1651 585
R6514 GND.n2208 GND.n1651 585
R6515 GND.n2118 GND.n1646 585
R6516 GND.n2211 GND.n1646 585
R6517 GND.n1682 GND.n1678 585
R6518 GND.n1684 GND.n1682 585
R6519 GND.n2114 GND.n2113 585
R6520 GND.n2113 GND.n2112 585
R6521 GND.n1681 GND.n1680 585
R6522 GND.n2101 GND.n1681 585
R6523 GND.n1702 GND.n1695 585
R6524 GND.n2104 GND.n1695 585
R6525 GND.n2098 GND.n2097 585
R6526 GND.n2099 GND.n2098 585
R6527 GND.n1701 GND.n1700 585
R6528 GND.n1709 GND.n1700 585
R6529 GND.n2092 GND.n2091 585
R6530 GND.n2091 GND.n2090 585
R6531 GND.n1705 GND.n1704 585
R6532 GND.n2077 GND.n1705 585
R6533 GND.n1730 GND.n1716 585
R6534 GND.n2080 GND.n1716 585
R6535 GND.n2045 GND.n2044 585
R6536 GND.n2046 GND.n2045 585
R6537 GND.n1729 GND.n1728 585
R6538 GND.n1728 GND.n1727 585
R6539 GND.n2039 GND.n2038 585
R6540 GND.n2038 GND.n2037 585
R6541 GND.n1733 GND.n1732 585
R6542 GND.n2023 GND.n1733 585
R6543 GND.n1752 GND.n1746 585
R6544 GND.n2027 GND.n1746 585
R6545 GND.n2020 GND.n2019 585
R6546 GND.n2021 GND.n2020 585
R6547 GND.n1751 GND.n1750 585
R6548 GND.n2004 GND.n1750 585
R6549 GND.n2014 GND.n2013 585
R6550 GND.n2013 GND.n2012 585
R6551 GND.n1971 GND.n1970 585
R6552 GND.n1972 GND.n1971 585
R6553 GND.n1969 GND.n1289 585
R6554 GND.n5373 GND.n1289 585
R6555 GND.n1757 GND.n1756 585
R6556 GND.n1756 GND.n1755 585
R6557 GND.n1965 GND.n1277 585
R6558 GND.n5379 GND.n1277 585
R6559 GND.n6354 GND.n446 585
R6560 GND.n6350 GND.n446 585
R6561 GND.n6356 GND.n6355 585
R6562 GND.n6357 GND.n6356 585
R6563 GND.n430 GND.n429 585
R6564 GND.n4714 GND.n430 585
R6565 GND.n6365 GND.n6364 585
R6566 GND.n6364 GND.n6363 585
R6567 GND.n6366 GND.n425 585
R6568 GND.n4720 GND.n425 585
R6569 GND.n6368 GND.n6367 585
R6570 GND.n6369 GND.n6368 585
R6571 GND.n409 GND.n408 585
R6572 GND.n4726 GND.n409 585
R6573 GND.n6377 GND.n6376 585
R6574 GND.n6376 GND.n6375 585
R6575 GND.n6378 GND.n404 585
R6576 GND.n4732 GND.n404 585
R6577 GND.n6380 GND.n6379 585
R6578 GND.n6381 GND.n6380 585
R6579 GND.n388 GND.n387 585
R6580 GND.n4738 GND.n388 585
R6581 GND.n6389 GND.n6388 585
R6582 GND.n6388 GND.n6387 585
R6583 GND.n6390 GND.n383 585
R6584 GND.n4744 GND.n383 585
R6585 GND.n6392 GND.n6391 585
R6586 GND.n6393 GND.n6392 585
R6587 GND.n367 GND.n366 585
R6588 GND.n4750 GND.n367 585
R6589 GND.n6401 GND.n6400 585
R6590 GND.n6400 GND.n6399 585
R6591 GND.n6402 GND.n362 585
R6592 GND.n4756 GND.n362 585
R6593 GND.n6404 GND.n6403 585
R6594 GND.n6405 GND.n6404 585
R6595 GND.n347 GND.n346 585
R6596 GND.n4762 GND.n347 585
R6597 GND.n6413 GND.n6412 585
R6598 GND.n6412 GND.n6411 585
R6599 GND.n6414 GND.n341 585
R6600 GND.n4768 GND.n341 585
R6601 GND.n6416 GND.n6415 585
R6602 GND.n6417 GND.n6416 585
R6603 GND.n342 GND.n340 585
R6604 GND.n4774 GND.n340 585
R6605 GND.n4780 GND.n4779 585
R6606 GND.n4783 GND.n4780 585
R6607 GND.n2877 GND.n2876 585
R6608 GND.n2876 GND.n2872 585
R6609 GND.n4632 GND.n320 585
R6610 GND.n6424 GND.n320 585
R6611 GND.n4631 GND.n4630 585
R6612 GND.n4630 GND.n2744 585
R6613 GND.n2736 GND.n2735 585
R6614 GND.n4793 GND.n2736 585
R6615 GND.n4798 GND.n4797 585
R6616 GND.n4797 GND.n4796 585
R6617 GND.n4799 GND.n2731 585
R6618 GND.n4623 GND.n2731 585
R6619 GND.n4801 GND.n4800 585
R6620 GND.n4802 GND.n4801 585
R6621 GND.n2717 GND.n2716 585
R6622 GND.n4611 GND.n2717 585
R6623 GND.n4810 GND.n4809 585
R6624 GND.n4809 GND.n4808 585
R6625 GND.n4811 GND.n2712 585
R6626 GND.n4604 GND.n2712 585
R6627 GND.n4813 GND.n4812 585
R6628 GND.n4814 GND.n4813 585
R6629 GND.n2696 GND.n2695 585
R6630 GND.n4596 GND.n2696 585
R6631 GND.n4822 GND.n4821 585
R6632 GND.n4821 GND.n4820 585
R6633 GND.n4823 GND.n2691 585
R6634 GND.n4589 GND.n2691 585
R6635 GND.n4825 GND.n4824 585
R6636 GND.n4826 GND.n4825 585
R6637 GND.n2675 GND.n2674 585
R6638 GND.n4581 GND.n2675 585
R6639 GND.n4834 GND.n4833 585
R6640 GND.n4833 GND.n4832 585
R6641 GND.n4835 GND.n2670 585
R6642 GND.n4574 GND.n2670 585
R6643 GND.n4837 GND.n4836 585
R6644 GND.n4838 GND.n4837 585
R6645 GND.n2654 GND.n2653 585
R6646 GND.n4566 GND.n2654 585
R6647 GND.n4846 GND.n4845 585
R6648 GND.n4845 GND.n4844 585
R6649 GND.n4847 GND.n2648 585
R6650 GND.n4559 GND.n2648 585
R6651 GND.n4849 GND.n4848 585
R6652 GND.n4850 GND.n4849 585
R6653 GND.n2649 GND.n2647 585
R6654 GND.n4551 GND.n2647 585
R6655 GND.n4546 GND.n2628 585
R6656 GND.n4856 GND.n2628 585
R6657 GND.n4545 GND.n4544 585
R6658 GND.n4544 GND.n2624 585
R6659 GND.n4543 GND.n4542 585
R6660 GND.n4543 GND.n2614 585
R6661 GND.n2608 GND.n2518 585
R6662 GND.n4864 GND.n2518 585
R6663 GND.n4960 GND.n4959 585
R6664 GND.n2519 GND.n2517 585
R6665 GND.n2939 GND.n2931 585
R6666 GND.n2941 GND.n2940 585
R6667 GND.n2943 GND.n2942 585
R6668 GND.n2911 GND.n2910 585
R6669 GND.n4522 GND.n2912 585
R6670 GND.n4523 GND.n2907 585
R6671 GND.n2906 GND.n2544 585
R6672 GND.n4957 GND.n2544 585
R6673 GND.n4707 GND.n4706 585
R6674 GND.n4704 GND.n4679 585
R6675 GND.n4703 GND.n4702 585
R6676 GND.n4696 GND.n4681 585
R6677 GND.n4698 GND.n4697 585
R6678 GND.n4694 GND.n4683 585
R6679 GND.n4693 GND.n4692 585
R6680 GND.n4686 GND.n4685 585
R6681 GND.n4688 GND.n4687 585
R6682 GND.n4687 GND.n633 585
R6683 GND.n4710 GND.n451 585
R6684 GND.n6350 GND.n451 585
R6685 GND.n4711 GND.n444 585
R6686 GND.n6357 GND.n444 585
R6687 GND.n4713 GND.n4712 585
R6688 GND.n4714 GND.n4713 585
R6689 GND.n4671 GND.n433 585
R6690 GND.n6363 GND.n433 585
R6691 GND.n4722 GND.n4721 585
R6692 GND.n4721 GND.n4720 585
R6693 GND.n4723 GND.n423 585
R6694 GND.n6369 GND.n423 585
R6695 GND.n4725 GND.n4724 585
R6696 GND.n4726 GND.n4725 585
R6697 GND.n4664 GND.n412 585
R6698 GND.n6375 GND.n412 585
R6699 GND.n4734 GND.n4733 585
R6700 GND.n4733 GND.n4732 585
R6701 GND.n4735 GND.n402 585
R6702 GND.n6381 GND.n402 585
R6703 GND.n4737 GND.n4736 585
R6704 GND.n4738 GND.n4737 585
R6705 GND.n4657 GND.n391 585
R6706 GND.n6387 GND.n391 585
R6707 GND.n4746 GND.n4745 585
R6708 GND.n4745 GND.n4744 585
R6709 GND.n4747 GND.n381 585
R6710 GND.n6393 GND.n381 585
R6711 GND.n4749 GND.n4748 585
R6712 GND.n4750 GND.n4749 585
R6713 GND.n4650 GND.n370 585
R6714 GND.n6399 GND.n370 585
R6715 GND.n4758 GND.n4757 585
R6716 GND.n4757 GND.n4756 585
R6717 GND.n4759 GND.n360 585
R6718 GND.n6405 GND.n360 585
R6719 GND.n4761 GND.n4760 585
R6720 GND.n4762 GND.n4761 585
R6721 GND.n4643 GND.n350 585
R6722 GND.n6411 GND.n350 585
R6723 GND.n4770 GND.n4769 585
R6724 GND.n4769 GND.n4768 585
R6725 GND.n4771 GND.n338 585
R6726 GND.n6417 GND.n338 585
R6727 GND.n4773 GND.n4772 585
R6728 GND.n4774 GND.n4773 585
R6729 GND.n4638 GND.n2874 585
R6730 GND.n4783 GND.n2874 585
R6731 GND.n316 GND.n314 585
R6732 GND.n2872 GND.n316 585
R6733 GND.n6426 GND.n6425 585
R6734 GND.n6425 GND.n6424 585
R6735 GND.n315 GND.n313 585
R6736 GND.n2744 GND.n315 585
R6737 GND.n4619 GND.n2743 585
R6738 GND.n4793 GND.n2743 585
R6739 GND.n4620 GND.n2739 585
R6740 GND.n4796 GND.n2739 585
R6741 GND.n4622 GND.n4621 585
R6742 GND.n4623 GND.n4622 585
R6743 GND.n2883 GND.n2729 585
R6744 GND.n4802 GND.n2729 585
R6745 GND.n4613 GND.n4612 585
R6746 GND.n4612 GND.n4611 585
R6747 GND.n2885 GND.n2720 585
R6748 GND.n4808 GND.n2720 585
R6749 GND.n4603 GND.n4602 585
R6750 GND.n4604 GND.n4603 585
R6751 GND.n2887 GND.n2710 585
R6752 GND.n4814 GND.n2710 585
R6753 GND.n4598 GND.n4597 585
R6754 GND.n4597 GND.n4596 585
R6755 GND.n2889 GND.n2699 585
R6756 GND.n4820 GND.n2699 585
R6757 GND.n4588 GND.n4587 585
R6758 GND.n4589 GND.n4588 585
R6759 GND.n2891 GND.n2689 585
R6760 GND.n4826 GND.n2689 585
R6761 GND.n4583 GND.n4582 585
R6762 GND.n4582 GND.n4581 585
R6763 GND.n2893 GND.n2678 585
R6764 GND.n4832 GND.n2678 585
R6765 GND.n4573 GND.n4572 585
R6766 GND.n4574 GND.n4573 585
R6767 GND.n2895 GND.n2668 585
R6768 GND.n4838 GND.n2668 585
R6769 GND.n4568 GND.n4567 585
R6770 GND.n4567 GND.n4566 585
R6771 GND.n2897 GND.n2657 585
R6772 GND.n4844 GND.n2657 585
R6773 GND.n4558 GND.n4557 585
R6774 GND.n4559 GND.n4558 585
R6775 GND.n2899 GND.n2645 585
R6776 GND.n4850 GND.n2645 585
R6777 GND.n4553 GND.n4552 585
R6778 GND.n4552 GND.n4551 585
R6779 GND.n4537 GND.n2626 585
R6780 GND.n4856 GND.n2626 585
R6781 GND.n4536 GND.n4535 585
R6782 GND.n4535 GND.n2624 585
R6783 GND.n4534 GND.n2901 585
R6784 GND.n4534 GND.n2614 585
R6785 GND.n4530 GND.n2613 585
R6786 GND.n4864 GND.n2613 585
R6787 GND.n4344 GND.n3053 585
R6788 GND.n3053 GND.n3029 585
R6789 GND.n4343 GND.n4342 585
R6790 GND.n4342 GND.n4341 585
R6791 GND.n3061 GND.n3060 585
R6792 GND.n3062 GND.n3061 585
R6793 GND.n4314 GND.n4313 585
R6794 GND.n4314 GND.n3071 585
R6795 GND.n4316 GND.n4315 585
R6796 GND.n4315 GND.n3070 585
R6797 GND.n4317 GND.n3085 585
R6798 GND.n4302 GND.n3085 585
R6799 GND.n4319 GND.n4318 585
R6800 GND.n4320 GND.n4319 585
R6801 GND.n4312 GND.n3084 585
R6802 GND.n3084 GND.n3079 585
R6803 GND.n4311 GND.n4310 585
R6804 GND.n4310 GND.n4309 585
R6805 GND.n3087 GND.n3086 585
R6806 GND.n3088 GND.n3087 585
R6807 GND.n4245 GND.n4244 585
R6808 GND.n4246 GND.n4245 585
R6809 GND.n4243 GND.n3097 585
R6810 GND.n4239 GND.n3097 585
R6811 GND.n4242 GND.n4241 585
R6812 GND.n4241 GND.n4240 585
R6813 GND.n3099 GND.n3098 585
R6814 GND.n3105 GND.n3099 585
R6815 GND.n4232 GND.n4231 585
R6816 GND.n4233 GND.n4232 585
R6817 GND.n4230 GND.n3107 585
R6818 GND.n3107 GND.n3104 585
R6819 GND.n4229 GND.n4228 585
R6820 GND.n4228 GND.n4227 585
R6821 GND.n3109 GND.n3108 585
R6822 GND.n3123 GND.n3109 585
R6823 GND.n4205 GND.n4204 585
R6824 GND.n4206 GND.n4205 585
R6825 GND.n4203 GND.n3124 585
R6826 GND.n3124 GND.n3120 585
R6827 GND.n4202 GND.n4201 585
R6828 GND.n4201 GND.n4200 585
R6829 GND.n3126 GND.n3125 585
R6830 GND.n3127 GND.n3126 585
R6831 GND.n4152 GND.n4151 585
R6832 GND.n4152 GND.n3136 585
R6833 GND.n4154 GND.n4153 585
R6834 GND.n4153 GND.n3135 585
R6835 GND.n4155 GND.n3150 585
R6836 GND.n4140 GND.n3150 585
R6837 GND.n4157 GND.n4156 585
R6838 GND.n4158 GND.n4157 585
R6839 GND.n4150 GND.n3149 585
R6840 GND.n3149 GND.n3145 585
R6841 GND.n4149 GND.n4148 585
R6842 GND.n4148 GND.n4147 585
R6843 GND.n3152 GND.n3151 585
R6844 GND.n3159 GND.n3152 585
R6845 GND.n4122 GND.n4121 585
R6846 GND.n4123 GND.n4122 585
R6847 GND.n4120 GND.n3162 585
R6848 GND.n3162 GND.n3158 585
R6849 GND.n4119 GND.n4118 585
R6850 GND.n4118 GND.n4117 585
R6851 GND.n3164 GND.n3163 585
R6852 GND.n3177 GND.n3164 585
R6853 GND.n4094 GND.n3175 585
R6854 GND.n4106 GND.n3175 585
R6855 GND.n4095 GND.n3184 585
R6856 GND.n3184 GND.n3174 585
R6857 GND.n4097 GND.n4096 585
R6858 GND.n4098 GND.n4097 585
R6859 GND.n4093 GND.n3183 585
R6860 GND.n4089 GND.n3183 585
R6861 GND.n4092 GND.n4091 585
R6862 GND.n4091 GND.n4090 585
R6863 GND.n3186 GND.n3185 585
R6864 GND.n3192 GND.n3186 585
R6865 GND.n4082 GND.n4081 585
R6866 GND.n4083 GND.n4082 585
R6867 GND.n4080 GND.n3194 585
R6868 GND.n3194 GND.n3191 585
R6869 GND.n4079 GND.n4078 585
R6870 GND.n4078 GND.n4077 585
R6871 GND.n3196 GND.n3195 585
R6872 GND.n3210 GND.n3196 585
R6873 GND.n4058 GND.n4057 585
R6874 GND.n4059 GND.n4058 585
R6875 GND.n4056 GND.n3211 585
R6876 GND.n3211 GND.n3207 585
R6877 GND.n4055 GND.n4054 585
R6878 GND.n4054 GND.n4053 585
R6879 GND.n3213 GND.n3212 585
R6880 GND.n3214 GND.n3213 585
R6881 GND.n3992 GND.n3991 585
R6882 GND.n3992 GND.n3223 585
R6883 GND.n3994 GND.n3993 585
R6884 GND.n3993 GND.n3222 585
R6885 GND.n3995 GND.n3237 585
R6886 GND.n3980 GND.n3237 585
R6887 GND.n3997 GND.n3996 585
R6888 GND.n3998 GND.n3997 585
R6889 GND.n3990 GND.n3236 585
R6890 GND.n3236 GND.n3232 585
R6891 GND.n3989 GND.n3988 585
R6892 GND.n3988 GND.n3987 585
R6893 GND.n3239 GND.n3238 585
R6894 GND.n3247 GND.n3239 585
R6895 GND.n3962 GND.n3961 585
R6896 GND.n3963 GND.n3962 585
R6897 GND.n3960 GND.n3249 585
R6898 GND.n3249 GND.n3246 585
R6899 GND.n3959 GND.n3958 585
R6900 GND.n3958 GND.n3957 585
R6901 GND.n3251 GND.n3250 585
R6902 GND.n3263 GND.n3251 585
R6903 GND.n3934 GND.n3261 585
R6904 GND.n3946 GND.n3261 585
R6905 GND.n3935 GND.n3272 585
R6906 GND.n3272 GND.n3260 585
R6907 GND.n3937 GND.n3936 585
R6908 GND.n3938 GND.n3937 585
R6909 GND.n3933 GND.n3271 585
R6910 GND.n3929 GND.n3271 585
R6911 GND.n3932 GND.n3931 585
R6912 GND.n3931 GND.n3930 585
R6913 GND.n3274 GND.n3273 585
R6914 GND.n3280 GND.n3274 585
R6915 GND.n3922 GND.n3921 585
R6916 GND.n3923 GND.n3922 585
R6917 GND.n3920 GND.n3283 585
R6918 GND.n3283 GND.n3279 585
R6919 GND.n3919 GND.n3918 585
R6920 GND.n3918 GND.n3917 585
R6921 GND.n3285 GND.n3284 585
R6922 GND.n3298 GND.n3285 585
R6923 GND.n3898 GND.n3897 585
R6924 GND.n3899 GND.n3898 585
R6925 GND.n3896 GND.n3299 585
R6926 GND.n3299 GND.n3295 585
R6927 GND.n3895 GND.n3894 585
R6928 GND.n3894 GND.n3893 585
R6929 GND.n3301 GND.n3300 585
R6930 GND.n3302 GND.n3301 585
R6931 GND.n3831 GND.n3830 585
R6932 GND.n3831 GND.n3311 585
R6933 GND.n3833 GND.n3832 585
R6934 GND.n3832 GND.n3310 585
R6935 GND.n3834 GND.n3324 585
R6936 GND.n3819 GND.n3324 585
R6937 GND.n3836 GND.n3835 585
R6938 GND.n3837 GND.n3836 585
R6939 GND.n3829 GND.n3323 585
R6940 GND.n3323 GND.n3319 585
R6941 GND.n3828 GND.n3827 585
R6942 GND.n3827 GND.n3826 585
R6943 GND.n3326 GND.n3325 585
R6944 GND.n3333 GND.n3326 585
R6945 GND.n3801 GND.n3800 585
R6946 GND.n3802 GND.n3801 585
R6947 GND.n3799 GND.n3335 585
R6948 GND.n3335 GND.n3332 585
R6949 GND.n3798 GND.n3797 585
R6950 GND.n3797 GND.n3796 585
R6951 GND.n3337 GND.n3336 585
R6952 GND.n3351 GND.n3337 585
R6953 GND.n3773 GND.n3349 585
R6954 GND.n3785 GND.n3349 585
R6955 GND.n3774 GND.n3359 585
R6956 GND.n3359 GND.n3348 585
R6957 GND.n3776 GND.n3775 585
R6958 GND.n3777 GND.n3776 585
R6959 GND.n3772 GND.n3358 585
R6960 GND.n3768 GND.n3358 585
R6961 GND.n3771 GND.n3770 585
R6962 GND.n3770 GND.n3769 585
R6963 GND.n3361 GND.n3360 585
R6964 GND.n3368 GND.n3361 585
R6965 GND.n3761 GND.n3760 585
R6966 GND.n3762 GND.n3761 585
R6967 GND.n3759 GND.n3370 585
R6968 GND.n3370 GND.n3367 585
R6969 GND.n3758 GND.n3757 585
R6970 GND.n3757 GND.n3756 585
R6971 GND.n3650 GND.n3377 585
R6972 GND.n3735 GND.n3734 585
R6973 GND.n3733 GND.n3649 585
R6974 GND.n3737 GND.n3649 585
R6975 GND.n3732 GND.n3731 585
R6976 GND.n3730 GND.n3729 585
R6977 GND.n3728 GND.n3727 585
R6978 GND.n3726 GND.n3725 585
R6979 GND.n3724 GND.n3723 585
R6980 GND.n3722 GND.n3721 585
R6981 GND.n3720 GND.n3719 585
R6982 GND.n3718 GND.n3717 585
R6983 GND.n3716 GND.n3715 585
R6984 GND.n3714 GND.n3713 585
R6985 GND.n3712 GND.n3711 585
R6986 GND.n3710 GND.n3709 585
R6987 GND.n3708 GND.n3707 585
R6988 GND.n3705 GND.n3704 585
R6989 GND.n3703 GND.n3702 585
R6990 GND.n3701 GND.n3700 585
R6991 GND.n3699 GND.n3698 585
R6992 GND.n3695 GND.n3694 585
R6993 GND.n3693 GND.n3692 585
R6994 GND.n3691 GND.n3690 585
R6995 GND.n3689 GND.n3688 585
R6996 GND.n3686 GND.n3685 585
R6997 GND.n3684 GND.n3683 585
R6998 GND.n3682 GND.n3681 585
R6999 GND.n3680 GND.n3679 585
R7000 GND.n3678 GND.n3677 585
R7001 GND.n3676 GND.n3675 585
R7002 GND.n3674 GND.n3673 585
R7003 GND.n3672 GND.n3671 585
R7004 GND.n3670 GND.n3669 585
R7005 GND.n3668 GND.n3667 585
R7006 GND.n3666 GND.n3665 585
R7007 GND.n3664 GND.n3663 585
R7008 GND.n3662 GND.n3661 585
R7009 GND.n3660 GND.n3659 585
R7010 GND.n3658 GND.n3657 585
R7011 GND.n3656 GND.n3407 585
R7012 GND.n3737 GND.n3407 585
R7013 GND.n4294 GND.n4293 585
R7014 GND.n4292 GND.n4291 585
R7015 GND.n4290 GND.n4289 585
R7016 GND.n4288 GND.n4287 585
R7017 GND.n4286 GND.n4285 585
R7018 GND.n4284 GND.n4283 585
R7019 GND.n4282 GND.n4281 585
R7020 GND.n4280 GND.n4279 585
R7021 GND.n4278 GND.n4277 585
R7022 GND.n4276 GND.n4275 585
R7023 GND.n4274 GND.n4273 585
R7024 GND.n4272 GND.n4271 585
R7025 GND.n4270 GND.n4269 585
R7026 GND.n4268 GND.n4267 585
R7027 GND.n4266 GND.n4265 585
R7028 GND.n4264 GND.n4263 585
R7029 GND.n4262 GND.n4261 585
R7030 GND.n4260 GND.n4259 585
R7031 GND.n4258 GND.n4257 585
R7032 GND.n4256 GND.n4255 585
R7033 GND.n4388 GND.n3031 585
R7034 GND.n4349 GND.n4348 585
R7035 GND.n4351 GND.n4350 585
R7036 GND.n4353 GND.n4352 585
R7037 GND.n4355 GND.n4354 585
R7038 GND.n4358 GND.n4357 585
R7039 GND.n4360 GND.n4359 585
R7040 GND.n4362 GND.n4361 585
R7041 GND.n4364 GND.n4363 585
R7042 GND.n4366 GND.n4365 585
R7043 GND.n4368 GND.n4367 585
R7044 GND.n4370 GND.n4369 585
R7045 GND.n4372 GND.n4371 585
R7046 GND.n4374 GND.n4373 585
R7047 GND.n4376 GND.n4375 585
R7048 GND.n4378 GND.n4377 585
R7049 GND.n4380 GND.n4379 585
R7050 GND.n4382 GND.n4381 585
R7051 GND.n4384 GND.n4383 585
R7052 GND.n4385 GND.n3054 585
R7053 GND.n4387 GND.n4386 585
R7054 GND.n4388 GND.n4387 585
R7055 GND.n4296 GND.n4295 585
R7056 GND.n4295 GND.n3029 585
R7057 GND.n4297 GND.n3063 585
R7058 GND.n4341 GND.n3063 585
R7059 GND.n4298 GND.n4251 585
R7060 GND.n4251 GND.n3062 585
R7061 GND.n4300 GND.n4299 585
R7062 GND.n4300 GND.n3071 585
R7063 GND.n4301 GND.n4250 585
R7064 GND.n4301 GND.n3070 585
R7065 GND.n4304 GND.n4303 585
R7066 GND.n4303 GND.n4302 585
R7067 GND.n4305 GND.n3081 585
R7068 GND.n4320 GND.n3081 585
R7069 GND.n4306 GND.n3091 585
R7070 GND.n3091 GND.n3079 585
R7071 GND.n4308 GND.n4307 585
R7072 GND.n4309 GND.n4308 585
R7073 GND.n4249 GND.n3090 585
R7074 GND.n3090 GND.n3088 585
R7075 GND.n4248 GND.n4247 585
R7076 GND.n4247 GND.n4246 585
R7077 GND.n3093 GND.n3092 585
R7078 GND.n4239 GND.n3093 585
R7079 GND.n4238 GND.n4237 585
R7080 GND.n4240 GND.n4238 585
R7081 GND.n4236 GND.n3101 585
R7082 GND.n3105 GND.n3101 585
R7083 GND.n4235 GND.n4234 585
R7084 GND.n4234 GND.n4233 585
R7085 GND.n3103 GND.n3102 585
R7086 GND.n3104 GND.n3103 585
R7087 GND.n4129 GND.n3112 585
R7088 GND.n4227 GND.n3112 585
R7089 GND.n4131 GND.n4130 585
R7090 GND.n4130 GND.n3123 585
R7091 GND.n4132 GND.n3122 585
R7092 GND.n4206 GND.n3122 585
R7093 GND.n4134 GND.n4133 585
R7094 GND.n4133 GND.n3120 585
R7095 GND.n4135 GND.n3128 585
R7096 GND.n4200 GND.n3128 585
R7097 GND.n4136 GND.n4128 585
R7098 GND.n4128 GND.n3127 585
R7099 GND.n4138 GND.n4137 585
R7100 GND.n4138 GND.n3136 585
R7101 GND.n4139 GND.n4127 585
R7102 GND.n4139 GND.n3135 585
R7103 GND.n4142 GND.n4141 585
R7104 GND.n4141 GND.n4140 585
R7105 GND.n4143 GND.n3147 585
R7106 GND.n4158 GND.n3147 585
R7107 GND.n4144 GND.n3155 585
R7108 GND.n3155 GND.n3145 585
R7109 GND.n4146 GND.n4145 585
R7110 GND.n4147 GND.n4146 585
R7111 GND.n4126 GND.n3154 585
R7112 GND.n3159 GND.n3154 585
R7113 GND.n4125 GND.n4124 585
R7114 GND.n4124 GND.n4123 585
R7115 GND.n3157 GND.n3156 585
R7116 GND.n3158 GND.n3157 585
R7117 GND.n4102 GND.n3166 585
R7118 GND.n4117 GND.n3166 585
R7119 GND.n4103 GND.n3179 585
R7120 GND.n3179 GND.n3177 585
R7121 GND.n4105 GND.n4104 585
R7122 GND.n4106 GND.n4105 585
R7123 GND.n4101 GND.n3178 585
R7124 GND.n3178 GND.n3174 585
R7125 GND.n4100 GND.n4099 585
R7126 GND.n4099 GND.n4098 585
R7127 GND.n3181 GND.n3180 585
R7128 GND.n4089 GND.n3181 585
R7129 GND.n4088 GND.n4087 585
R7130 GND.n4090 GND.n4088 585
R7131 GND.n4086 GND.n3188 585
R7132 GND.n3192 GND.n3188 585
R7133 GND.n4085 GND.n4084 585
R7134 GND.n4084 GND.n4083 585
R7135 GND.n3190 GND.n3189 585
R7136 GND.n3191 GND.n3190 585
R7137 GND.n3969 GND.n3198 585
R7138 GND.n4077 GND.n3198 585
R7139 GND.n3971 GND.n3970 585
R7140 GND.n3970 GND.n3210 585
R7141 GND.n3972 GND.n3209 585
R7142 GND.n4059 GND.n3209 585
R7143 GND.n3974 GND.n3973 585
R7144 GND.n3973 GND.n3207 585
R7145 GND.n3975 GND.n3215 585
R7146 GND.n4053 GND.n3215 585
R7147 GND.n3976 GND.n3968 585
R7148 GND.n3968 GND.n3214 585
R7149 GND.n3978 GND.n3977 585
R7150 GND.n3978 GND.n3223 585
R7151 GND.n3979 GND.n3967 585
R7152 GND.n3979 GND.n3222 585
R7153 GND.n3982 GND.n3981 585
R7154 GND.n3981 GND.n3980 585
R7155 GND.n3983 GND.n3234 585
R7156 GND.n3998 GND.n3234 585
R7157 GND.n3984 GND.n3243 585
R7158 GND.n3243 GND.n3232 585
R7159 GND.n3986 GND.n3985 585
R7160 GND.n3987 GND.n3986 585
R7161 GND.n3966 GND.n3242 585
R7162 GND.n3247 GND.n3242 585
R7163 GND.n3965 GND.n3964 585
R7164 GND.n3964 GND.n3963 585
R7165 GND.n3245 GND.n3244 585
R7166 GND.n3246 GND.n3245 585
R7167 GND.n3942 GND.n3252 585
R7168 GND.n3957 GND.n3252 585
R7169 GND.n3943 GND.n3266 585
R7170 GND.n3266 GND.n3263 585
R7171 GND.n3945 GND.n3944 585
R7172 GND.n3946 GND.n3945 585
R7173 GND.n3941 GND.n3265 585
R7174 GND.n3265 GND.n3260 585
R7175 GND.n3940 GND.n3939 585
R7176 GND.n3939 GND.n3938 585
R7177 GND.n3268 GND.n3267 585
R7178 GND.n3929 GND.n3268 585
R7179 GND.n3928 GND.n3927 585
R7180 GND.n3930 GND.n3928 585
R7181 GND.n3926 GND.n3276 585
R7182 GND.n3280 GND.n3276 585
R7183 GND.n3925 GND.n3924 585
R7184 GND.n3924 GND.n3923 585
R7185 GND.n3278 GND.n3277 585
R7186 GND.n3279 GND.n3278 585
R7187 GND.n3808 GND.n3287 585
R7188 GND.n3917 GND.n3287 585
R7189 GND.n3810 GND.n3809 585
R7190 GND.n3809 GND.n3298 585
R7191 GND.n3811 GND.n3297 585
R7192 GND.n3899 GND.n3297 585
R7193 GND.n3813 GND.n3812 585
R7194 GND.n3812 GND.n3295 585
R7195 GND.n3814 GND.n3303 585
R7196 GND.n3893 GND.n3303 585
R7197 GND.n3815 GND.n3807 585
R7198 GND.n3807 GND.n3302 585
R7199 GND.n3817 GND.n3816 585
R7200 GND.n3817 GND.n3311 585
R7201 GND.n3818 GND.n3806 585
R7202 GND.n3818 GND.n3310 585
R7203 GND.n3821 GND.n3820 585
R7204 GND.n3820 GND.n3819 585
R7205 GND.n3822 GND.n3321 585
R7206 GND.n3837 GND.n3321 585
R7207 GND.n3823 GND.n3329 585
R7208 GND.n3329 GND.n3319 585
R7209 GND.n3825 GND.n3824 585
R7210 GND.n3826 GND.n3825 585
R7211 GND.n3805 GND.n3328 585
R7212 GND.n3333 GND.n3328 585
R7213 GND.n3804 GND.n3803 585
R7214 GND.n3803 GND.n3802 585
R7215 GND.n3331 GND.n3330 585
R7216 GND.n3332 GND.n3331 585
R7217 GND.n3781 GND.n3340 585
R7218 GND.n3796 GND.n3340 585
R7219 GND.n3782 GND.n3353 585
R7220 GND.n3353 GND.n3351 585
R7221 GND.n3784 GND.n3783 585
R7222 GND.n3785 GND.n3784 585
R7223 GND.n3780 GND.n3352 585
R7224 GND.n3352 GND.n3348 585
R7225 GND.n3779 GND.n3778 585
R7226 GND.n3778 GND.n3777 585
R7227 GND.n3355 GND.n3354 585
R7228 GND.n3768 GND.n3355 585
R7229 GND.n3767 GND.n3766 585
R7230 GND.n3769 GND.n3767 585
R7231 GND.n3765 GND.n3364 585
R7232 GND.n3368 GND.n3364 585
R7233 GND.n3764 GND.n3763 585
R7234 GND.n3763 GND.n3762 585
R7235 GND.n3366 GND.n3365 585
R7236 GND.n3367 GND.n3366 585
R7237 GND.n3655 GND.n3378 585
R7238 GND.n3756 GND.n3378 585
R7239 GND.n5293 GND.n5292 585
R7240 GND.n5294 GND.n5293 585
R7241 GND.n1402 GND.n1400 585
R7242 GND.n2345 GND.n1400 585
R7243 GND.n2341 GND.n2340 585
R7244 GND.n2342 GND.n2341 585
R7245 GND.n1546 GND.n1545 585
R7246 GND.n2278 GND.n1545 585
R7247 GND.n2336 GND.n2335 585
R7248 GND.n2335 GND.n2334 585
R7249 GND.n1549 GND.n1548 585
R7250 GND.n2330 GND.n1549 585
R7251 GND.n2304 GND.n2303 585
R7252 GND.n2305 GND.n2304 585
R7253 GND.n1565 GND.n1564 585
R7254 GND.n1564 GND.n1561 585
R7255 GND.n2299 GND.n2298 585
R7256 GND.n2298 GND.n2297 585
R7257 GND.n1568 GND.n1567 585
R7258 GND.n2292 GND.n1568 585
R7259 GND.n2266 GND.n1586 585
R7260 GND.n1586 GND.n1585 585
R7261 GND.n2268 GND.n2267 585
R7262 GND.n2269 GND.n2268 585
R7263 GND.n1587 GND.n1583 585
R7264 GND.n2256 GND.n1583 585
R7265 GND.n2261 GND.n2260 585
R7266 GND.n2260 GND.n2259 585
R7267 GND.n1590 GND.n1589 585
R7268 GND.n2253 GND.n1590 585
R7269 GND.n2241 GND.n1609 585
R7270 GND.n1609 GND.n1608 585
R7271 GND.n2243 GND.n2242 585
R7272 GND.n2244 GND.n2243 585
R7273 GND.n1610 GND.n1607 585
R7274 GND.n2231 GND.n1607 585
R7275 GND.n2236 GND.n2235 585
R7276 GND.n2235 GND.n2234 585
R7277 GND.n1613 GND.n1612 585
R7278 GND.n2229 GND.n1613 585
R7279 GND.n2217 GND.n1632 585
R7280 GND.n1632 GND.n1631 585
R7281 GND.n2219 GND.n2218 585
R7282 GND.n2220 GND.n2219 585
R7283 GND.n1633 GND.n1630 585
R7284 GND.n2140 GND.n1630 585
R7285 GND.n2135 GND.n2134 585
R7286 GND.n2136 GND.n2135 585
R7287 GND.n2133 GND.n1668 585
R7288 GND.n2191 GND.n1668 585
R7289 GND.n2196 GND.n2195 585
R7290 GND.n2195 GND.n2194 585
R7291 GND.n2198 GND.n2197 585
R7292 GND.n2199 GND.n2198 585
R7293 GND.n1667 GND.n1666 585
R7294 GND.n1667 GND.n1659 585
R7295 GND.n1665 GND.n1639 585
R7296 GND.n1665 GND.n1652 585
R7297 GND.n1643 GND.n1640 585
R7298 GND.n2208 GND.n1643 585
R7299 GND.n2213 GND.n2212 585
R7300 GND.n2212 GND.n2211 585
R7301 GND.n1642 GND.n1641 585
R7302 GND.n1684 GND.n1642 585
R7303 GND.n2111 GND.n2110 585
R7304 GND.n2112 GND.n2111 585
R7305 GND.n1689 GND.n1688 585
R7306 GND.n2101 GND.n1688 585
R7307 GND.n2106 GND.n2105 585
R7308 GND.n2105 GND.n2104 585
R7309 GND.n1692 GND.n1691 585
R7310 GND.n2099 GND.n1692 585
R7311 GND.n2087 GND.n1710 585
R7312 GND.n1710 GND.n1709 585
R7313 GND.n2089 GND.n2088 585
R7314 GND.n2090 GND.n2089 585
R7315 GND.n1711 GND.n1708 585
R7316 GND.n2077 GND.n1708 585
R7317 GND.n2082 GND.n2081 585
R7318 GND.n2081 GND.n2080 585
R7319 GND.n1714 GND.n1713 585
R7320 GND.n2046 GND.n1714 585
R7321 GND.n2034 GND.n1740 585
R7322 GND.n1740 GND.n1727 585
R7323 GND.n2036 GND.n2035 585
R7324 GND.n2037 GND.n2036 585
R7325 GND.n1741 GND.n1739 585
R7326 GND.n2023 GND.n1739 585
R7327 GND.n2029 GND.n2028 585
R7328 GND.n2028 GND.n2027 585
R7329 GND.n1744 GND.n1743 585
R7330 GND.n2021 GND.n1744 585
R7331 GND.n2009 GND.n2005 585
R7332 GND.n2005 GND.n2004 585
R7333 GND.n2011 GND.n2010 585
R7334 GND.n2012 GND.n2011 585
R7335 GND.n1286 GND.n1285 585
R7336 GND.n1972 GND.n1286 585
R7337 GND.n5375 GND.n5374 585
R7338 GND.n5374 GND.n5373 585
R7339 GND.n5376 GND.n1281 585
R7340 GND.n1755 GND.n1281 585
R7341 GND.n5378 GND.n5377 585
R7342 GND.n5379 GND.n5378 585
R7343 GND.n1820 GND.n1280 585
R7344 GND.n1823 GND.n1822 585
R7345 GND.n1818 GND.n1817 585
R7346 GND.n1817 GND.n1267 585
R7347 GND.n1828 GND.n1827 585
R7348 GND.n1830 GND.n1816 585
R7349 GND.n1833 GND.n1832 585
R7350 GND.n1814 GND.n1813 585
R7351 GND.n1840 GND.n1839 585
R7352 GND.n1842 GND.n1812 585
R7353 GND.n1845 GND.n1844 585
R7354 GND.n1810 GND.n1809 585
R7355 GND.n1850 GND.n1849 585
R7356 GND.n1852 GND.n1808 585
R7357 GND.n1855 GND.n1854 585
R7358 GND.n1806 GND.n1805 585
R7359 GND.n1860 GND.n1859 585
R7360 GND.n1862 GND.n1804 585
R7361 GND.n1865 GND.n1864 585
R7362 GND.n1800 GND.n1799 585
R7363 GND.n1870 GND.n1869 585
R7364 GND.n1872 GND.n1798 585
R7365 GND.n1875 GND.n1874 585
R7366 GND.n1796 GND.n1795 585
R7367 GND.n1880 GND.n1879 585
R7368 GND.n1882 GND.n1791 585
R7369 GND.n1885 GND.n1884 585
R7370 GND.n1789 GND.n1788 585
R7371 GND.n1890 GND.n1889 585
R7372 GND.n1892 GND.n1787 585
R7373 GND.n1895 GND.n1894 585
R7374 GND.n1785 GND.n1784 585
R7375 GND.n1900 GND.n1899 585
R7376 GND.n1902 GND.n1783 585
R7377 GND.n1905 GND.n1904 585
R7378 GND.n1781 GND.n1780 585
R7379 GND.n1912 GND.n1911 585
R7380 GND.n1914 GND.n1779 585
R7381 GND.n1917 GND.n1916 585
R7382 GND.n1777 GND.n1776 585
R7383 GND.n1922 GND.n1921 585
R7384 GND.n1924 GND.n1775 585
R7385 GND.n1927 GND.n1926 585
R7386 GND.n1773 GND.n1772 585
R7387 GND.n1932 GND.n1931 585
R7388 GND.n1934 GND.n1771 585
R7389 GND.n1936 GND.n1935 585
R7390 GND.n1935 GND.n1267 585
R7391 GND.n5225 GND.n1394 585
R7392 GND.n5226 GND.n1469 585
R7393 GND.n5227 GND.n1465 585
R7394 GND.n5228 GND.n1464 585
R7395 GND.n1520 GND.n1462 585
R7396 GND.n5232 GND.n1461 585
R7397 GND.n5233 GND.n1460 585
R7398 GND.n5234 GND.n1459 585
R7399 GND.n1517 GND.n1457 585
R7400 GND.n5238 GND.n1456 585
R7401 GND.n5239 GND.n1455 585
R7402 GND.n5240 GND.n1452 585
R7403 GND.n1514 GND.n1450 585
R7404 GND.n5244 GND.n1449 585
R7405 GND.n5245 GND.n1448 585
R7406 GND.n5246 GND.n1447 585
R7407 GND.n1511 GND.n1445 585
R7408 GND.n5250 GND.n1444 585
R7409 GND.n5251 GND.n1443 585
R7410 GND.n5252 GND.n1442 585
R7411 GND.n1508 GND.n1437 585
R7412 GND.n5256 GND.n1436 585
R7413 GND.n5257 GND.n1435 585
R7414 GND.n5258 GND.n1434 585
R7415 GND.n5191 GND.n1506 585
R7416 GND.n5175 GND.n1431 585
R7417 GND.n5263 GND.n1430 585
R7418 GND.n5264 GND.n1429 585
R7419 GND.n5265 GND.n1428 585
R7420 GND.n5179 GND.n1424 585
R7421 GND.n5269 GND.n1423 585
R7422 GND.n5270 GND.n1422 585
R7423 GND.n5271 GND.n1421 585
R7424 GND.n5182 GND.n1419 585
R7425 GND.n5275 GND.n1418 585
R7426 GND.n5276 GND.n1417 585
R7427 GND.n5277 GND.n1416 585
R7428 GND.n5185 GND.n1414 585
R7429 GND.n5281 GND.n1411 585
R7430 GND.n5282 GND.n1410 585
R7431 GND.n5283 GND.n1409 585
R7432 GND.n5188 GND.n1407 585
R7433 GND.n5287 GND.n1406 585
R7434 GND.n5288 GND.n1405 585
R7435 GND.n5289 GND.n1401 585
R7436 GND.n5191 GND.n1401 585
R7437 GND.n5296 GND.n5295 585
R7438 GND.n5295 GND.n5294 585
R7439 GND.n5297 GND.n1393 585
R7440 GND.n2345 GND.n1393 585
R7441 GND.n1544 GND.n1388 585
R7442 GND.n2342 GND.n1544 585
R7443 GND.n5301 GND.n1387 585
R7444 GND.n2278 GND.n1387 585
R7445 GND.n5302 GND.n1386 585
R7446 GND.n2334 GND.n1386 585
R7447 GND.n5303 GND.n1385 585
R7448 GND.n2330 GND.n1385 585
R7449 GND.n1562 GND.n1380 585
R7450 GND.n2305 GND.n1562 585
R7451 GND.n5307 GND.n1379 585
R7452 GND.n1561 GND.n1379 585
R7453 GND.n5308 GND.n1378 585
R7454 GND.n2297 GND.n1378 585
R7455 GND.n5309 GND.n1377 585
R7456 GND.n2292 GND.n1377 585
R7457 GND.n1584 GND.n1372 585
R7458 GND.n1585 GND.n1584 585
R7459 GND.n5313 GND.n1371 585
R7460 GND.n2269 GND.n1371 585
R7461 GND.n5314 GND.n1370 585
R7462 GND.n2256 GND.n1370 585
R7463 GND.n5315 GND.n1369 585
R7464 GND.n2259 GND.n1369 585
R7465 GND.n1596 GND.n1364 585
R7466 GND.n2253 GND.n1596 585
R7467 GND.n5319 GND.n1363 585
R7468 GND.n1608 GND.n1363 585
R7469 GND.n5320 GND.n1362 585
R7470 GND.n2244 GND.n1362 585
R7471 GND.n5321 GND.n1361 585
R7472 GND.n2231 GND.n1361 585
R7473 GND.n1615 GND.n1356 585
R7474 GND.n2234 GND.n1615 585
R7475 GND.n5325 GND.n1355 585
R7476 GND.n2229 GND.n1355 585
R7477 GND.n5326 GND.n1354 585
R7478 GND.n1631 GND.n1354 585
R7479 GND.n5327 GND.n1353 585
R7480 GND.n2220 GND.n1353 585
R7481 GND.n2138 GND.n1348 585
R7482 GND.n2140 GND.n2138 585
R7483 GND.n5331 GND.n1347 585
R7484 GND.n2136 GND.n1347 585
R7485 GND.n5332 GND.n1346 585
R7486 GND.n2191 GND.n1346 585
R7487 GND.n5333 GND.n1345 585
R7488 GND.n2194 GND.n1345 585
R7489 GND.n1660 GND.n1340 585
R7490 GND.n2199 GND.n1660 585
R7491 GND.n5337 GND.n1339 585
R7492 GND.n1659 GND.n1339 585
R7493 GND.n5338 GND.n1338 585
R7494 GND.n1652 GND.n1338 585
R7495 GND.n5339 GND.n1337 585
R7496 GND.n2208 GND.n1337 585
R7497 GND.n1645 GND.n1332 585
R7498 GND.n2211 GND.n1645 585
R7499 GND.n5343 GND.n1331 585
R7500 GND.n1684 GND.n1331 585
R7501 GND.n5344 GND.n1330 585
R7502 GND.n2112 GND.n1330 585
R7503 GND.n5345 GND.n1329 585
R7504 GND.n2101 GND.n1329 585
R7505 GND.n1694 GND.n1324 585
R7506 GND.n2104 GND.n1694 585
R7507 GND.n5349 GND.n1323 585
R7508 GND.n2099 GND.n1323 585
R7509 GND.n5350 GND.n1322 585
R7510 GND.n1709 GND.n1322 585
R7511 GND.n5351 GND.n1321 585
R7512 GND.n2090 GND.n1321 585
R7513 GND.n1720 GND.n1316 585
R7514 GND.n2077 GND.n1720 585
R7515 GND.n5355 GND.n1315 585
R7516 GND.n2080 GND.n1315 585
R7517 GND.n5356 GND.n1314 585
R7518 GND.n2046 GND.n1314 585
R7519 GND.n5357 GND.n1313 585
R7520 GND.n1727 GND.n1313 585
R7521 GND.n1735 GND.n1308 585
R7522 GND.n2037 GND.n1735 585
R7523 GND.n5361 GND.n1307 585
R7524 GND.n2023 GND.n1307 585
R7525 GND.n5362 GND.n1306 585
R7526 GND.n2027 GND.n1306 585
R7527 GND.n5363 GND.n1305 585
R7528 GND.n2021 GND.n1305 585
R7529 GND.n2003 GND.n1300 585
R7530 GND.n2004 GND.n2003 585
R7531 GND.n5367 GND.n1299 585
R7532 GND.n2012 GND.n1299 585
R7533 GND.n5368 GND.n1298 585
R7534 GND.n1972 GND.n1298 585
R7535 GND.n5369 GND.n1288 585
R7536 GND.n5373 GND.n1288 585
R7537 GND.n1754 GND.n1297 585
R7538 GND.n1755 GND.n1754 585
R7539 GND.n1939 GND.n1276 585
R7540 GND.n5379 GND.n1276 585
R7541 GND.n441 GND.n440 585
R7542 GND.n6350 GND.n441 585
R7543 GND.n6359 GND.n6358 585
R7544 GND.n6358 GND.n6357 585
R7545 GND.n6360 GND.n435 585
R7546 GND.n4714 GND.n435 585
R7547 GND.n6362 GND.n6361 585
R7548 GND.n6363 GND.n6362 585
R7549 GND.n420 GND.n419 585
R7550 GND.n4720 GND.n420 585
R7551 GND.n6371 GND.n6370 585
R7552 GND.n6370 GND.n6369 585
R7553 GND.n6372 GND.n414 585
R7554 GND.n4726 GND.n414 585
R7555 GND.n6374 GND.n6373 585
R7556 GND.n6375 GND.n6374 585
R7557 GND.n399 GND.n398 585
R7558 GND.n4732 GND.n399 585
R7559 GND.n6383 GND.n6382 585
R7560 GND.n6382 GND.n6381 585
R7561 GND.n6384 GND.n393 585
R7562 GND.n4738 GND.n393 585
R7563 GND.n6386 GND.n6385 585
R7564 GND.n6387 GND.n6386 585
R7565 GND.n378 GND.n377 585
R7566 GND.n4744 GND.n378 585
R7567 GND.n6395 GND.n6394 585
R7568 GND.n6394 GND.n6393 585
R7569 GND.n6396 GND.n372 585
R7570 GND.n4750 GND.n372 585
R7571 GND.n6398 GND.n6397 585
R7572 GND.n6399 GND.n6398 585
R7573 GND.n357 GND.n356 585
R7574 GND.n4756 GND.n357 585
R7575 GND.n6407 GND.n6406 585
R7576 GND.n6406 GND.n6405 585
R7577 GND.n6408 GND.n352 585
R7578 GND.n4762 GND.n352 585
R7579 GND.n6410 GND.n6409 585
R7580 GND.n6411 GND.n6410 585
R7581 GND.n335 GND.n333 585
R7582 GND.n4768 GND.n335 585
R7583 GND.n6419 GND.n6418 585
R7584 GND.n6418 GND.n6417 585
R7585 GND.n334 GND.n332 585
R7586 GND.n4774 GND.n334 585
R7587 GND.n4782 GND.n4781 585
R7588 GND.n4783 GND.n4782 585
R7589 GND.n324 GND.n322 585
R7590 GND.n2872 GND.n322 585
R7591 GND.n6423 GND.n6422 585
R7592 GND.n6424 GND.n6423 585
R7593 GND.n323 GND.n321 585
R7594 GND.n2744 GND.n321 585
R7595 GND.n4794 GND.n2741 585
R7596 GND.n4794 GND.n4793 585
R7597 GND.n4795 GND.n330 585
R7598 GND.n4796 GND.n4795 585
R7599 GND.n2726 GND.n2725 585
R7600 GND.n4623 GND.n2726 585
R7601 GND.n4804 GND.n4803 585
R7602 GND.n4803 GND.n4802 585
R7603 GND.n4805 GND.n2722 585
R7604 GND.n4611 GND.n2722 585
R7605 GND.n4807 GND.n4806 585
R7606 GND.n4808 GND.n4807 585
R7607 GND.n2707 GND.n2706 585
R7608 GND.n4604 GND.n2707 585
R7609 GND.n4816 GND.n4815 585
R7610 GND.n4815 GND.n4814 585
R7611 GND.n4817 GND.n2701 585
R7612 GND.n4596 GND.n2701 585
R7613 GND.n4819 GND.n4818 585
R7614 GND.n4820 GND.n4819 585
R7615 GND.n2686 GND.n2685 585
R7616 GND.n4589 GND.n2686 585
R7617 GND.n4828 GND.n4827 585
R7618 GND.n4827 GND.n4826 585
R7619 GND.n4829 GND.n2680 585
R7620 GND.n4581 GND.n2680 585
R7621 GND.n4831 GND.n4830 585
R7622 GND.n4832 GND.n4831 585
R7623 GND.n2665 GND.n2664 585
R7624 GND.n4574 GND.n2665 585
R7625 GND.n4840 GND.n4839 585
R7626 GND.n4839 GND.n4838 585
R7627 GND.n4841 GND.n2659 585
R7628 GND.n4566 GND.n2659 585
R7629 GND.n4843 GND.n4842 585
R7630 GND.n4844 GND.n4843 585
R7631 GND.n2642 GND.n2641 585
R7632 GND.n4559 GND.n2642 585
R7633 GND.n4852 GND.n4851 585
R7634 GND.n4851 GND.n4850 585
R7635 GND.n4853 GND.n2630 585
R7636 GND.n4551 GND.n2630 585
R7637 GND.n4855 GND.n4854 585
R7638 GND.n4856 GND.n4855 585
R7639 GND.n2631 GND.n2629 585
R7640 GND.n2629 GND.n2624 585
R7641 GND.n2635 GND.n2634 585
R7642 GND.n2634 GND.n2614 585
R7643 GND.n2633 GND.n2550 585
R7644 GND.n4864 GND.n2550 585
R7645 GND.n4955 GND.n4954 585
R7646 GND.n4953 GND.n2549 585
R7647 GND.n4952 GND.n2548 585
R7648 GND.n4957 GND.n2548 585
R7649 GND.n4951 GND.n4950 585
R7650 GND.n4949 GND.n4948 585
R7651 GND.n4947 GND.n4946 585
R7652 GND.n4945 GND.n4944 585
R7653 GND.n4943 GND.n4942 585
R7654 GND.n4941 GND.n4940 585
R7655 GND.n4939 GND.n4938 585
R7656 GND.n4937 GND.n4936 585
R7657 GND.n4935 GND.n4934 585
R7658 GND.n4933 GND.n4932 585
R7659 GND.n4931 GND.n4930 585
R7660 GND.n4929 GND.n4928 585
R7661 GND.n4927 GND.n4926 585
R7662 GND.n4925 GND.n2569 585
R7663 GND.n4924 GND.n4923 585
R7664 GND.n4922 GND.n4921 585
R7665 GND.n4920 GND.n4919 585
R7666 GND.n4917 GND.n4916 585
R7667 GND.n4915 GND.n4914 585
R7668 GND.n4913 GND.n4912 585
R7669 GND.n4911 GND.n4910 585
R7670 GND.n4908 GND.n4907 585
R7671 GND.n4906 GND.n4905 585
R7672 GND.n4904 GND.n4903 585
R7673 GND.n4902 GND.n4901 585
R7674 GND.n4900 GND.n4899 585
R7675 GND.n4898 GND.n4897 585
R7676 GND.n4896 GND.n4895 585
R7677 GND.n4894 GND.n4893 585
R7678 GND.n4892 GND.n4891 585
R7679 GND.n4890 GND.n4889 585
R7680 GND.n4888 GND.n4887 585
R7681 GND.n4886 GND.n4885 585
R7682 GND.n4884 GND.n4883 585
R7683 GND.n4882 GND.n4881 585
R7684 GND.n4880 GND.n4879 585
R7685 GND.n4878 GND.n4877 585
R7686 GND.n4876 GND.n4875 585
R7687 GND.n4874 GND.n4873 585
R7688 GND.n2607 GND.n2604 585
R7689 GND.n4869 GND.n2542 585
R7690 GND.n4957 GND.n2542 585
R7691 GND.n484 GND.n450 585
R7692 GND.n631 GND.n630 585
R7693 GND.n629 GND.n483 585
R7694 GND.n623 GND.n489 585
R7695 GND.n625 GND.n624 585
R7696 GND.n622 GND.n621 585
R7697 GND.n620 GND.n619 585
R7698 GND.n613 GND.n491 585
R7699 GND.n615 GND.n614 585
R7700 GND.n612 GND.n611 585
R7701 GND.n610 GND.n609 585
R7702 GND.n608 GND.n607 585
R7703 GND.n606 GND.n496 585
R7704 GND.n602 GND.n601 585
R7705 GND.n600 GND.n599 585
R7706 GND.n598 GND.n597 585
R7707 GND.n596 GND.n498 585
R7708 GND.n592 GND.n591 585
R7709 GND.n590 GND.n589 585
R7710 GND.n588 GND.n587 585
R7711 GND.n586 GND.n585 585
R7712 GND.n579 GND.n504 585
R7713 GND.n581 GND.n580 585
R7714 GND.n578 GND.n577 585
R7715 GND.n576 GND.n575 585
R7716 GND.n569 GND.n506 585
R7717 GND.n571 GND.n570 585
R7718 GND.n568 GND.n567 585
R7719 GND.n566 GND.n565 585
R7720 GND.n559 GND.n510 585
R7721 GND.n561 GND.n560 585
R7722 GND.n558 GND.n557 585
R7723 GND.n556 GND.n555 585
R7724 GND.n549 GND.n512 585
R7725 GND.n551 GND.n550 585
R7726 GND.n548 GND.n547 585
R7727 GND.n546 GND.n545 585
R7728 GND.n518 GND.n514 585
R7729 GND.n541 GND.n519 585
R7730 GND.n540 GND.n539 585
R7731 GND.n538 GND.n537 585
R7732 GND.n531 GND.n520 585
R7733 GND.n533 GND.n532 585
R7734 GND.n530 GND.n529 585
R7735 GND.n528 GND.n527 585
R7736 GND.n523 GND.n522 585
R7737 GND.n6352 GND.n6351 585
R7738 GND.n6351 GND.n6350 585
R7739 GND.n449 GND.n443 585
R7740 GND.n6357 GND.n443 585
R7741 GND.n4716 GND.n4715 585
R7742 GND.n4715 GND.n4714 585
R7743 GND.n4717 GND.n432 585
R7744 GND.n6363 GND.n432 585
R7745 GND.n4719 GND.n4718 585
R7746 GND.n4720 GND.n4719 585
R7747 GND.n4666 GND.n422 585
R7748 GND.n6369 GND.n422 585
R7749 GND.n4728 GND.n4727 585
R7750 GND.n4727 GND.n4726 585
R7751 GND.n4729 GND.n411 585
R7752 GND.n6375 GND.n411 585
R7753 GND.n4731 GND.n4730 585
R7754 GND.n4732 GND.n4731 585
R7755 GND.n4659 GND.n401 585
R7756 GND.n6381 GND.n401 585
R7757 GND.n4740 GND.n4739 585
R7758 GND.n4739 GND.n4738 585
R7759 GND.n4741 GND.n390 585
R7760 GND.n6387 GND.n390 585
R7761 GND.n4743 GND.n4742 585
R7762 GND.n4744 GND.n4743 585
R7763 GND.n4652 GND.n380 585
R7764 GND.n6393 GND.n380 585
R7765 GND.n4752 GND.n4751 585
R7766 GND.n4751 GND.n4750 585
R7767 GND.n4753 GND.n369 585
R7768 GND.n6399 GND.n369 585
R7769 GND.n4755 GND.n4754 585
R7770 GND.n4756 GND.n4755 585
R7771 GND.n4645 GND.n359 585
R7772 GND.n6405 GND.n359 585
R7773 GND.n4764 GND.n4763 585
R7774 GND.n4763 GND.n4762 585
R7775 GND.n4765 GND.n349 585
R7776 GND.n6411 GND.n349 585
R7777 GND.n4767 GND.n4766 585
R7778 GND.n4768 GND.n4767 585
R7779 GND.n4637 GND.n337 585
R7780 GND.n6417 GND.n337 585
R7781 GND.n4776 GND.n4775 585
R7782 GND.n4775 GND.n4774 585
R7783 GND.n4777 GND.n2873 585
R7784 GND.n4783 GND.n2873 585
R7785 GND.n4636 GND.n4635 585
R7786 GND.n4635 GND.n2872 585
R7787 GND.n4634 GND.n318 585
R7788 GND.n6424 GND.n318 585
R7789 GND.n2881 GND.n2880 585
R7790 GND.n2880 GND.n2744 585
R7791 GND.n4627 GND.n2742 585
R7792 GND.n4793 GND.n2742 585
R7793 GND.n4626 GND.n2738 585
R7794 GND.n4796 GND.n2738 585
R7795 GND.n4625 GND.n4624 585
R7796 GND.n4624 GND.n4623 585
R7797 GND.n2882 GND.n2728 585
R7798 GND.n4802 GND.n2728 585
R7799 GND.n4610 GND.n4609 585
R7800 GND.n4611 GND.n4610 585
R7801 GND.n4607 GND.n2719 585
R7802 GND.n4808 GND.n2719 585
R7803 GND.n4606 GND.n4605 585
R7804 GND.n4605 GND.n4604 585
R7805 GND.n2886 GND.n2709 585
R7806 GND.n4814 GND.n2709 585
R7807 GND.n4595 GND.n4594 585
R7808 GND.n4596 GND.n4595 585
R7809 GND.n4592 GND.n2698 585
R7810 GND.n4820 GND.n2698 585
R7811 GND.n4591 GND.n4590 585
R7812 GND.n4590 GND.n4589 585
R7813 GND.n2890 GND.n2688 585
R7814 GND.n4826 GND.n2688 585
R7815 GND.n4580 GND.n4579 585
R7816 GND.n4581 GND.n4580 585
R7817 GND.n4577 GND.n2677 585
R7818 GND.n4832 GND.n2677 585
R7819 GND.n4576 GND.n4575 585
R7820 GND.n4575 GND.n4574 585
R7821 GND.n2894 GND.n2667 585
R7822 GND.n4838 GND.n2667 585
R7823 GND.n4565 GND.n4564 585
R7824 GND.n4566 GND.n4565 585
R7825 GND.n4562 GND.n2656 585
R7826 GND.n4844 GND.n2656 585
R7827 GND.n4561 GND.n4560 585
R7828 GND.n4560 GND.n4559 585
R7829 GND.n2898 GND.n2644 585
R7830 GND.n4850 GND.n2644 585
R7831 GND.n4550 GND.n4549 585
R7832 GND.n4551 GND.n4550 585
R7833 GND.n4538 GND.n2625 585
R7834 GND.n4856 GND.n2625 585
R7835 GND.n4540 GND.n4539 585
R7836 GND.n4539 GND.n2624 585
R7837 GND.n2611 GND.n2610 585
R7838 GND.n2614 GND.n2611 585
R7839 GND.n4866 GND.n4865 585
R7840 GND.n4865 GND.n4864 585
R7841 GND.n6313 GND.n6312 585
R7842 GND.n6312 GND.n6311 585
R7843 GND.n6314 GND.n659 585
R7844 GND.n659 GND.n658 585
R7845 GND.n6316 GND.n6315 585
R7846 GND.n6317 GND.n6316 585
R7847 GND.n657 GND.n656 585
R7848 GND.n6318 GND.n657 585
R7849 GND.n6321 GND.n6320 585
R7850 GND.n6320 GND.n6319 585
R7851 GND.n6322 GND.n651 585
R7852 GND.n651 GND.n650 585
R7853 GND.n6324 GND.n6323 585
R7854 GND.n6325 GND.n6324 585
R7855 GND.n649 GND.n648 585
R7856 GND.n6326 GND.n649 585
R7857 GND.n6329 GND.n6328 585
R7858 GND.n6328 GND.n6327 585
R7859 GND.n6330 GND.n643 585
R7860 GND.n643 GND.n642 585
R7861 GND.n6332 GND.n6331 585
R7862 GND.n6333 GND.n6332 585
R7863 GND.n641 GND.n640 585
R7864 GND.n6334 GND.n641 585
R7865 GND.n6337 GND.n6336 585
R7866 GND.n6336 GND.n6335 585
R7867 GND.n6338 GND.n635 585
R7868 GND.n635 GND.n634 585
R7869 GND.n6340 GND.n6339 585
R7870 GND.n6341 GND.n6340 585
R7871 GND.n460 GND.n459 585
R7872 GND.n6342 GND.n460 585
R7873 GND.n6345 GND.n6344 585
R7874 GND.n6344 GND.n6343 585
R7875 GND.n6346 GND.n454 585
R7876 GND.n454 GND.n452 585
R7877 GND.n6348 GND.n6347 585
R7878 GND.n6349 GND.n6348 585
R7879 GND.n455 GND.n453 585
R7880 GND.n453 GND.n445 585
R7881 GND.n2838 GND.n2833 585
R7882 GND.n2833 GND.n442 585
R7883 GND.n2840 GND.n2839 585
R7884 GND.n2840 GND.n434 585
R7885 GND.n2841 GND.n2832 585
R7886 GND.n2841 GND.n431 585
R7887 GND.n2843 GND.n2842 585
R7888 GND.n2842 GND.n424 585
R7889 GND.n2844 GND.n2827 585
R7890 GND.n2827 GND.n421 585
R7891 GND.n2846 GND.n2845 585
R7892 GND.n2846 GND.n413 585
R7893 GND.n2847 GND.n2826 585
R7894 GND.n2847 GND.n410 585
R7895 GND.n2849 GND.n2848 585
R7896 GND.n2848 GND.n403 585
R7897 GND.n2850 GND.n2821 585
R7898 GND.n2821 GND.n400 585
R7899 GND.n2852 GND.n2851 585
R7900 GND.n2852 GND.n392 585
R7901 GND.n2853 GND.n2820 585
R7902 GND.n2853 GND.n389 585
R7903 GND.n2855 GND.n2854 585
R7904 GND.n2854 GND.n382 585
R7905 GND.n2856 GND.n2815 585
R7906 GND.n2815 GND.n379 585
R7907 GND.n2858 GND.n2857 585
R7908 GND.n2858 GND.n371 585
R7909 GND.n2859 GND.n2814 585
R7910 GND.n2859 GND.n368 585
R7911 GND.n2861 GND.n2860 585
R7912 GND.n2860 GND.n361 585
R7913 GND.n2862 GND.n2809 585
R7914 GND.n2809 GND.n358 585
R7915 GND.n2864 GND.n2863 585
R7916 GND.n2864 GND.n351 585
R7917 GND.n2865 GND.n2808 585
R7918 GND.n2865 GND.n348 585
R7919 GND.n2867 GND.n2866 585
R7920 GND.n2866 GND.n339 585
R7921 GND.n2869 GND.n2806 585
R7922 GND.n2806 GND.n336 585
R7923 GND.n2871 GND.n2870 585
R7924 GND.n2875 GND.n2871 585
R7925 GND.n4785 GND.n2805 585
R7926 GND.n4785 GND.n4784 585
R7927 GND.n4787 GND.n4786 585
R7928 GND.n4786 GND.n319 585
R7929 GND.n4789 GND.n2746 585
R7930 GND.n2746 GND.n317 585
R7931 GND.n4791 GND.n4790 585
R7932 GND.n4792 GND.n4791 585
R7933 GND.n2803 GND.n2745 585
R7934 GND.n2745 GND.n2740 585
R7935 GND.n2802 GND.n2801 585
R7936 GND.n2801 GND.n2737 585
R7937 GND.n2800 GND.n2799 585
R7938 GND.n2800 GND.n2730 585
R7939 GND.n2798 GND.n2748 585
R7940 GND.n2748 GND.n2727 585
R7941 GND.n2797 GND.n2796 585
R7942 GND.n2796 GND.n2721 585
R7943 GND.n2795 GND.n2749 585
R7944 GND.n2795 GND.n2718 585
R7945 GND.n2794 GND.n2793 585
R7946 GND.n2794 GND.n2711 585
R7947 GND.n2752 GND.n2751 585
R7948 GND.n2751 GND.n2708 585
R7949 GND.n2788 GND.n2787 585
R7950 GND.n2787 GND.n2700 585
R7951 GND.n2786 GND.n2754 585
R7952 GND.n2786 GND.n2697 585
R7953 GND.n2785 GND.n2784 585
R7954 GND.n2785 GND.n2690 585
R7955 GND.n2756 GND.n2755 585
R7956 GND.n2755 GND.n2687 585
R7957 GND.n2780 GND.n2779 585
R7958 GND.n2779 GND.n2679 585
R7959 GND.n2778 GND.n2758 585
R7960 GND.n2778 GND.n2676 585
R7961 GND.n2777 GND.n2776 585
R7962 GND.n2777 GND.n2669 585
R7963 GND.n2760 GND.n2759 585
R7964 GND.n2759 GND.n2666 585
R7965 GND.n2772 GND.n2771 585
R7966 GND.n2771 GND.n2658 585
R7967 GND.n2770 GND.n2762 585
R7968 GND.n2770 GND.n2655 585
R7969 GND.n2769 GND.n2768 585
R7970 GND.n2769 GND.n2646 585
R7971 GND.n2764 GND.n2763 585
R7972 GND.n2763 GND.n2643 585
R7973 GND.n2622 GND.n2621 585
R7974 GND.n2627 GND.n2622 585
R7975 GND.n4859 GND.n4858 585
R7976 GND.n4858 GND.n4857 585
R7977 GND.n4860 GND.n2616 585
R7978 GND.n2623 GND.n2616 585
R7979 GND.n4862 GND.n4861 585
R7980 GND.n4863 GND.n4862 585
R7981 GND.n2617 GND.n2615 585
R7982 GND.n2615 GND.n2612 585
R7983 GND.n4508 GND.n4507 585
R7984 GND.n4508 GND.n2543 585
R7985 GND.n4510 GND.n4509 585
R7986 GND.n4509 GND.n2520 585
R7987 GND.n4511 GND.n2952 585
R7988 GND.n2952 GND.n2950 585
R7989 GND.n4513 GND.n4512 585
R7990 GND.n4514 GND.n4513 585
R7991 GND.n2953 GND.n2951 585
R7992 GND.n2951 GND.n2496 585
R7993 GND.n4499 GND.n2495 585
R7994 GND.n4982 GND.n2495 585
R7995 GND.n4498 GND.n4497 585
R7996 GND.n4497 GND.n2494 585
R7997 GND.n4496 GND.n2955 585
R7998 GND.n4496 GND.n4495 585
R7999 GND.n4483 GND.n2956 585
R8000 GND.n2957 GND.n2956 585
R8001 GND.n4485 GND.n4484 585
R8002 GND.n4486 GND.n4485 585
R8003 GND.n2965 GND.n2964 585
R8004 GND.n2964 GND.n2963 585
R8005 GND.n4477 GND.n4476 585
R8006 GND.n4476 GND.n4475 585
R8007 GND.n2968 GND.n2967 585
R8008 GND.n2975 GND.n2968 585
R8009 GND.n4465 GND.n4464 585
R8010 GND.n4466 GND.n4465 585
R8011 GND.n2977 GND.n2976 585
R8012 GND.n2976 GND.n2974 585
R8013 GND.n4460 GND.n4459 585
R8014 GND.n4459 GND.n4458 585
R8015 GND.n2980 GND.n2979 585
R8016 GND.n2981 GND.n2980 585
R8017 GND.n4448 GND.n4447 585
R8018 GND.n4449 GND.n4448 585
R8019 GND.n2989 GND.n2988 585
R8020 GND.n2988 GND.n2987 585
R8021 GND.n4443 GND.n4442 585
R8022 GND.n4442 GND.n4441 585
R8023 GND.n2992 GND.n2991 585
R8024 GND.n2993 GND.n2992 585
R8025 GND.n4431 GND.n4430 585
R8026 GND.n4432 GND.n4431 585
R8027 GND.n3001 GND.n3000 585
R8028 GND.n3000 GND.n2999 585
R8029 GND.n4426 GND.n4425 585
R8030 GND.n4425 GND.n4424 585
R8031 GND.n3004 GND.n3003 585
R8032 GND.n3005 GND.n3004 585
R8033 GND.n4414 GND.n4413 585
R8034 GND.n4415 GND.n4414 585
R8035 GND.n3013 GND.n3012 585
R8036 GND.n3012 GND.n3011 585
R8037 GND.n4409 GND.n4408 585
R8038 GND.n4408 GND.n4407 585
R8039 GND.n3016 GND.n3015 585
R8040 GND.n3017 GND.n3016 585
R8041 GND.n4397 GND.n4396 585
R8042 GND.n4398 GND.n4397 585
R8043 GND.n3025 GND.n3024 585
R8044 GND.n3024 GND.n3023 585
R8045 GND.n4392 GND.n4391 585
R8046 GND.n4391 GND.n4390 585
R8047 GND.n3028 GND.n3027 585
R8048 GND.n4340 GND.n3028 585
R8049 GND.n4328 GND.n3074 585
R8050 GND.n3074 GND.n3073 585
R8051 GND.n4330 GND.n4329 585
R8052 GND.n4331 GND.n4330 585
R8053 GND.n3075 GND.n3072 585
R8054 GND.n3083 GND.n3072 585
R8055 GND.n4323 GND.n4322 585
R8056 GND.n4322 GND.n4321 585
R8057 GND.n3078 GND.n3077 585
R8058 GND.n4309 GND.n3078 585
R8059 GND.n4219 GND.n4218 585
R8060 GND.n4219 GND.n3096 585
R8061 GND.n4220 GND.n4215 585
R8062 GND.n4220 GND.n3095 585
R8063 GND.n4222 GND.n4221 585
R8064 GND.n4221 GND.n3100 585
R8065 GND.n4223 GND.n3115 585
R8066 GND.n3115 GND.n3106 585
R8067 GND.n4225 GND.n4224 585
R8068 GND.n4226 GND.n4225 585
R8069 GND.n3116 GND.n3114 585
R8070 GND.n3114 GND.n3111 585
R8071 GND.n4209 GND.n4208 585
R8072 GND.n4208 GND.n4207 585
R8073 GND.n3119 GND.n3118 585
R8074 GND.n4199 GND.n3119 585
R8075 GND.n4166 GND.n3140 585
R8076 GND.n3140 GND.n3139 585
R8077 GND.n4168 GND.n4167 585
R8078 GND.n4169 GND.n4168 585
R8079 GND.n3141 GND.n3138 585
R8080 GND.n3148 GND.n3138 585
R8081 GND.n4161 GND.n4160 585
R8082 GND.n4160 GND.n4159 585
R8083 GND.n3144 GND.n3143 585
R8084 GND.n3153 GND.n3144 585
R8085 GND.n4113 GND.n3169 585
R8086 GND.n3169 GND.n3161 585
R8087 GND.n4115 GND.n4114 585
R8088 GND.n4116 GND.n4115 585
R8089 GND.n3170 GND.n3168 585
R8090 GND.n3168 GND.n3165 585
R8091 GND.n4108 GND.n4107 585
R8092 GND.n4107 GND.n4106 585
R8093 GND.n3173 GND.n3172 585
R8094 GND.n4022 GND.n3173 585
R8095 GND.n4070 GND.n4069 585
R8096 GND.n4070 GND.n3182 585
R8097 GND.n4072 GND.n4071 585
R8098 GND.n4071 GND.n3187 585
R8099 GND.n4073 GND.n3202 585
R8100 GND.n3202 GND.n3193 585
R8101 GND.n4075 GND.n4074 585
R8102 GND.n4076 GND.n4075 585
R8103 GND.n3203 GND.n3201 585
R8104 GND.n3201 GND.n3197 585
R8105 GND.n4062 GND.n4061 585
R8106 GND.n4061 GND.n4060 585
R8107 GND.n3206 GND.n3205 585
R8108 GND.n4052 GND.n3206 585
R8109 GND.n4006 GND.n3227 585
R8110 GND.n3227 GND.n3226 585
R8111 GND.n4008 GND.n4007 585
R8112 GND.n4009 GND.n4008 585
R8113 GND.n3228 GND.n3224 585
R8114 GND.n3235 GND.n3224 585
R8115 GND.n4001 GND.n4000 585
R8116 GND.n4000 GND.n3999 585
R8117 GND.n3231 GND.n3230 585
R8118 GND.n3241 GND.n3231 585
R8119 GND.n3953 GND.n3255 585
R8120 GND.n3255 GND.n3248 585
R8121 GND.n3955 GND.n3954 585
R8122 GND.n3956 GND.n3955 585
R8123 GND.n3256 GND.n3254 585
R8124 GND.n3862 GND.n3254 585
R8125 GND.n3948 GND.n3947 585
R8126 GND.n3947 GND.n3946 585
R8127 GND.n3259 GND.n3258 585
R8128 GND.n3270 GND.n3259 585
R8129 GND.n3910 GND.n3909 585
R8130 GND.n3910 GND.n3269 585
R8131 GND.n3912 GND.n3911 585
R8132 GND.n3911 GND.n3275 585
R8133 GND.n3913 GND.n3290 585
R8134 GND.n3290 GND.n3282 585
R8135 GND.n3915 GND.n3914 585
R8136 GND.n3916 GND.n3915 585
R8137 GND.n3291 GND.n3289 585
R8138 GND.n3289 GND.n3286 585
R8139 GND.n3902 GND.n3901 585
R8140 GND.n3901 GND.n3900 585
R8141 GND.n3294 GND.n3293 585
R8142 GND.n3892 GND.n3294 585
R8143 GND.n3846 GND.n3314 585
R8144 GND.n3314 GND.n3313 585
R8145 GND.n3848 GND.n3847 585
R8146 GND.n3849 GND.n3848 585
R8147 GND.n3315 GND.n3312 585
R8148 GND.n3322 GND.n3312 585
R8149 GND.n3841 GND.n3840 585
R8150 GND.n3840 GND.n3839 585
R8151 GND.n3318 GND.n3317 585
R8152 GND.n3327 GND.n3318 585
R8153 GND.n3792 GND.n3343 585
R8154 GND.n3343 GND.n3334 585
R8155 GND.n3794 GND.n3793 585
R8156 GND.n3795 GND.n3794 585
R8157 GND.n3344 GND.n3342 585
R8158 GND.n3342 GND.n3339 585
R8159 GND.n3787 GND.n3786 585
R8160 GND.n3786 GND.n3785 585
R8161 GND.n3347 GND.n3346 585
R8162 GND.n3357 GND.n3347 585
R8163 GND.n3749 GND.n3748 585
R8164 GND.n3749 GND.n3356 585
R8165 GND.n3751 GND.n3750 585
R8166 GND.n3750 GND.n3363 585
R8167 GND.n3752 GND.n3381 585
R8168 GND.n3381 GND.n3369 585
R8169 GND.n3754 GND.n3753 585
R8170 GND.n3755 GND.n3754 585
R8171 GND.n3382 GND.n3380 585
R8172 GND.n3648 GND.n3380 585
R8173 GND.n3741 GND.n3740 585
R8174 GND.n3740 GND.n3739 585
R8175 GND.n3385 GND.n3384 585
R8176 GND.n3386 GND.n3385 585
R8177 GND.n3610 GND.n3609 585
R8178 GND.n3611 GND.n3610 585
R8179 GND.n3415 GND.n3414 585
R8180 GND.n3414 GND.n3413 585
R8181 GND.n3605 GND.n3604 585
R8182 GND.n3604 GND.n3603 585
R8183 GND.n3418 GND.n3417 585
R8184 GND.n3419 GND.n3418 585
R8185 GND.n3592 GND.n3591 585
R8186 GND.n3593 GND.n3592 585
R8187 GND.n3428 GND.n3427 585
R8188 GND.n3427 GND.n3426 585
R8189 GND.n3587 GND.n3586 585
R8190 GND.n3586 GND.n3585 585
R8191 GND.n3431 GND.n3430 585
R8192 GND.n3432 GND.n3431 585
R8193 GND.n3575 GND.n3574 585
R8194 GND.n3576 GND.n3575 585
R8195 GND.n3440 GND.n3439 585
R8196 GND.n3439 GND.n3438 585
R8197 GND.n3570 GND.n3569 585
R8198 GND.n3569 GND.n3568 585
R8199 GND.n3443 GND.n3442 585
R8200 GND.n3444 GND.n3443 585
R8201 GND.n3558 GND.n3557 585
R8202 GND.n3559 GND.n3558 585
R8203 GND.n3452 GND.n3451 585
R8204 GND.n3451 GND.n3450 585
R8205 GND.n3553 GND.n3552 585
R8206 GND.n3552 GND.n3551 585
R8207 GND.n3455 GND.n3454 585
R8208 GND.n3456 GND.n3455 585
R8209 GND.n3541 GND.n3540 585
R8210 GND.n3542 GND.n3541 585
R8211 GND.n3463 GND.n3462 585
R8212 GND.n3532 GND.n3462 585
R8213 GND.n3536 GND.n3535 585
R8214 GND.n3535 GND.n3534 585
R8215 GND.n3466 GND.n3465 585
R8216 GND.n3467 GND.n3466 585
R8217 GND.n3523 GND.n3522 585
R8218 GND.n3524 GND.n3523 585
R8219 GND.n3513 GND.n3512 585
R8220 GND.n3512 GND.n3511 585
R8221 GND.n3518 GND.n3517 585
R8222 GND.n3517 GND.n1534 585
R8223 GND.n3516 GND.n1532 585
R8224 GND.n5159 GND.n1532 585
R8225 GND.n5161 GND.n1531 585
R8226 GND.n5161 GND.n5160 585
R8227 GND.n5164 GND.n5163 585
R8228 GND.n5163 GND.n5162 585
R8229 GND.n5165 GND.n1526 585
R8230 GND.n1526 GND.n1524 585
R8231 GND.n5167 GND.n5166 585
R8232 GND.n5168 GND.n5167 585
R8233 GND.n1527 GND.n1525 585
R8234 GND.n1525 GND.n1505 585
R8235 GND.n2320 GND.n2315 585
R8236 GND.n2315 GND.n1397 585
R8237 GND.n2322 GND.n2321 585
R8238 GND.n2322 GND.n1395 585
R8239 GND.n2323 GND.n2314 585
R8240 GND.n2323 GND.n1541 585
R8241 GND.n2325 GND.n2324 585
R8242 GND.n2324 GND.n1543 585
R8243 GND.n2326 GND.n1556 585
R8244 GND.n1556 GND.n1551 585
R8245 GND.n2328 GND.n2327 585
R8246 GND.n2329 GND.n2328 585
R8247 GND.n1557 GND.n1555 585
R8248 GND.n1555 GND.n1553 585
R8249 GND.n2308 GND.n2307 585
R8250 GND.n2307 GND.n2306 585
R8251 GND.n1560 GND.n1559 585
R8252 GND.n1571 GND.n1560 585
R8253 GND.n2165 GND.n2164 585
R8254 GND.n2165 GND.n1569 585
R8255 GND.n2166 GND.n2161 585
R8256 GND.n2166 GND.n1573 585
R8257 GND.n2168 GND.n2167 585
R8258 GND.n2167 GND.n1581 585
R8259 GND.n2169 GND.n2156 585
R8260 GND.n2156 GND.n1580 585
R8261 GND.n2171 GND.n2170 585
R8262 GND.n2171 GND.n1593 585
R8263 GND.n2172 GND.n2155 585
R8264 GND.n2172 GND.n1591 585
R8265 GND.n2174 GND.n2173 585
R8266 GND.n2173 GND.n1595 585
R8267 GND.n2175 GND.n2150 585
R8268 GND.n2150 GND.n1604 585
R8269 GND.n2177 GND.n2176 585
R8270 GND.n2177 GND.n1603 585
R8271 GND.n2178 GND.n2149 585
R8272 GND.n2178 GND.n1617 585
R8273 GND.n2180 GND.n2179 585
R8274 GND.n2179 GND.n1614 585
R8275 GND.n2181 GND.n2146 585
R8276 GND.n2146 GND.n1620 585
R8277 GND.n2183 GND.n2182 585
R8278 GND.n2183 GND.n1628 585
R8279 GND.n2185 GND.n2184 585
R8280 GND.n2184 GND.n1627 585
R8281 GND.n2186 GND.n2142 585
R8282 GND.n2142 GND.n2141 585
R8283 GND.n2189 GND.n2188 585
R8284 GND.n2190 GND.n2189 585
R8285 GND.n2144 GND.n2137 585
R8286 GND.n2137 GND.n1670 585
R8287 GND.n1657 GND.n1656 585
R8288 GND.n1662 GND.n1657 585
R8289 GND.n2202 GND.n2201 585
R8290 GND.n2201 GND.n2200 585
R8291 GND.n2204 GND.n1654 585
R8292 GND.n1658 GND.n1654 585
R8293 GND.n2206 GND.n2205 585
R8294 GND.n2207 GND.n2206 585
R8295 GND.n1655 GND.n1653 585
R8296 GND.n1653 GND.n1647 585
R8297 GND.n2064 GND.n2063 585
R8298 GND.n2064 GND.n1644 585
R8299 GND.n2066 GND.n2065 585
R8300 GND.n2065 GND.n1685 585
R8301 GND.n2067 GND.n2057 585
R8302 GND.n2057 GND.n1683 585
R8303 GND.n2069 GND.n2068 585
R8304 GND.n2069 GND.n1696 585
R8305 GND.n2070 GND.n2056 585
R8306 GND.n2070 GND.n1693 585
R8307 GND.n2072 GND.n2071 585
R8308 GND.n2071 GND.n1699 585
R8309 GND.n2073 GND.n1722 585
R8310 GND.n1722 GND.n1706 585
R8311 GND.n2075 GND.n2074 585
R8312 GND.n2076 GND.n2075 585
R8313 GND.n1723 GND.n1721 585
R8314 GND.n1721 GND.n1717 585
R8315 GND.n2050 GND.n2049 585
R8316 GND.n2049 GND.n1715 585
R8317 GND.n2048 GND.n1725 585
R8318 GND.n2048 GND.n2047 585
R8319 GND.n1993 GND.n1726 585
R8320 GND.n1736 GND.n1726 585
R8321 GND.n1995 GND.n1994 585
R8322 GND.n1995 GND.n1734 585
R8323 GND.n1996 GND.n1989 585
R8324 GND.n1996 GND.n1747 585
R8325 GND.n1998 GND.n1997 585
R8326 GND.n1997 GND.n1745 585
R8327 GND.n1999 GND.n1976 585
R8328 GND.n1976 GND.n1749 585
R8329 GND.n2001 GND.n2000 585
R8330 GND.n2002 GND.n2001 585
R8331 GND.n1977 GND.n1975 585
R8332 GND.n1975 GND.n1973 585
R8333 GND.n1983 GND.n1982 585
R8334 GND.n1982 GND.n1290 585
R8335 GND.n1981 GND.n1980 585
R8336 GND.n1981 GND.n1287 585
R8337 GND.n1274 GND.n1273 585
R8338 GND.n1278 GND.n1274 585
R8339 GND.n5382 GND.n5381 585
R8340 GND.n5381 GND.n5380 585
R8341 GND.n5383 GND.n1268 585
R8342 GND.n1275 GND.n1268 585
R8343 GND.n5385 GND.n5384 585
R8344 GND.n5386 GND.n5385 585
R8345 GND.n1266 GND.n1265 585
R8346 GND.n5387 GND.n1266 585
R8347 GND.n5390 GND.n5389 585
R8348 GND.n5389 GND.n5388 585
R8349 GND.n5391 GND.n1260 585
R8350 GND.n1260 GND.n1259 585
R8351 GND.n5393 GND.n5392 585
R8352 GND.n5394 GND.n5393 585
R8353 GND.n1258 GND.n1257 585
R8354 GND.n5395 GND.n1258 585
R8355 GND.n5398 GND.n5397 585
R8356 GND.n5397 GND.n5396 585
R8357 GND.n5399 GND.n1252 585
R8358 GND.n1252 GND.n1251 585
R8359 GND.n5401 GND.n5400 585
R8360 GND.n5402 GND.n5401 585
R8361 GND.n1250 GND.n1249 585
R8362 GND.n5403 GND.n1250 585
R8363 GND.n5406 GND.n5405 585
R8364 GND.n5405 GND.n5404 585
R8365 GND.n5407 GND.n1244 585
R8366 GND.n1244 GND.n1243 585
R8367 GND.n5409 GND.n5408 585
R8368 GND.n5410 GND.n5409 585
R8369 GND.n1241 GND.n1240 585
R8370 GND.n5411 GND.n1241 585
R8371 GND.n5414 GND.n5413 585
R8372 GND.n5413 GND.n5412 585
R8373 GND.n5415 GND.n1238 585
R8374 GND.n1242 GND.n1238 585
R8375 GND.n5416 GND.n1235 585
R8376 GND.n1235 GND.n1234 585
R8377 GND.n4981 GND.n4980 585
R8378 GND.n4982 GND.n4981 585
R8379 GND.n2499 GND.n2497 585
R8380 GND.n2497 GND.n2494 585
R8381 GND.n4493 GND.n4492 585
R8382 GND.n4495 GND.n4493 585
R8383 GND.n2959 GND.n2958 585
R8384 GND.n2958 GND.n2957 585
R8385 GND.n4488 GND.n4487 585
R8386 GND.n4487 GND.n4486 585
R8387 GND.n2962 GND.n2961 585
R8388 GND.n2963 GND.n2962 585
R8389 GND.n4473 GND.n4472 585
R8390 GND.n4475 GND.n4473 585
R8391 GND.n2970 GND.n2969 585
R8392 GND.n2975 GND.n2969 585
R8393 GND.n4468 GND.n4467 585
R8394 GND.n4467 GND.n4466 585
R8395 GND.n2973 GND.n2972 585
R8396 GND.n2974 GND.n2973 585
R8397 GND.n4456 GND.n4455 585
R8398 GND.n4458 GND.n4456 585
R8399 GND.n2983 GND.n2982 585
R8400 GND.n2982 GND.n2981 585
R8401 GND.n4451 GND.n4450 585
R8402 GND.n4450 GND.n4449 585
R8403 GND.n2986 GND.n2985 585
R8404 GND.n2987 GND.n2986 585
R8405 GND.n4439 GND.n4438 585
R8406 GND.n4441 GND.n4439 585
R8407 GND.n2995 GND.n2994 585
R8408 GND.n2994 GND.n2993 585
R8409 GND.n4434 GND.n4433 585
R8410 GND.n4433 GND.n4432 585
R8411 GND.n2998 GND.n2997 585
R8412 GND.n2999 GND.n2998 585
R8413 GND.n4422 GND.n4421 585
R8414 GND.n4424 GND.n4422 585
R8415 GND.n3007 GND.n3006 585
R8416 GND.n3006 GND.n3005 585
R8417 GND.n4417 GND.n4416 585
R8418 GND.n4416 GND.n4415 585
R8419 GND.n3010 GND.n3009 585
R8420 GND.n3011 GND.n3010 585
R8421 GND.n4405 GND.n4404 585
R8422 GND.n4407 GND.n4405 585
R8423 GND.n3019 GND.n3018 585
R8424 GND.n3018 GND.n3017 585
R8425 GND.n4400 GND.n4399 585
R8426 GND.n4399 GND.n4398 585
R8427 GND.n3022 GND.n3021 585
R8428 GND.n3023 GND.n3022 585
R8429 GND.n3066 GND.n3030 585
R8430 GND.n4390 GND.n3030 585
R8431 GND.n4339 GND.n4338 585
R8432 GND.n4340 GND.n4339 585
R8433 GND.n3065 GND.n3064 585
R8434 GND.n3073 GND.n3064 585
R8435 GND.n4333 GND.n4332 585
R8436 GND.n4332 GND.n4331 585
R8437 GND.n3069 GND.n3068 585
R8438 GND.n3083 GND.n3069 585
R8439 GND.n4182 GND.n3080 585
R8440 GND.n4321 GND.n3080 585
R8441 GND.n4185 GND.n3089 585
R8442 GND.n4309 GND.n3089 585
R8443 GND.n4186 GND.n4181 585
R8444 GND.n4181 GND.n3096 585
R8445 GND.n4187 GND.n4180 585
R8446 GND.n4180 GND.n3095 585
R8447 GND.n4179 GND.n4177 585
R8448 GND.n4179 GND.n3100 585
R8449 GND.n4191 GND.n4176 585
R8450 GND.n4176 GND.n3106 585
R8451 GND.n4192 GND.n3113 585
R8452 GND.n4226 GND.n3113 585
R8453 GND.n4193 GND.n4175 585
R8454 GND.n4175 GND.n3111 585
R8455 GND.n3131 GND.n3121 585
R8456 GND.n4207 GND.n3121 585
R8457 GND.n4198 GND.n4197 585
R8458 GND.n4199 GND.n4198 585
R8459 GND.n3130 GND.n3129 585
R8460 GND.n3139 GND.n3129 585
R8461 GND.n4171 GND.n4170 585
R8462 GND.n4170 GND.n4169 585
R8463 GND.n3134 GND.n3133 585
R8464 GND.n3148 GND.n3134 585
R8465 GND.n4029 GND.n3146 585
R8466 GND.n4159 GND.n3146 585
R8467 GND.n4032 GND.n4028 585
R8468 GND.n4028 GND.n3153 585
R8469 GND.n4033 GND.n4027 585
R8470 GND.n4027 GND.n3161 585
R8471 GND.n4034 GND.n3167 585
R8472 GND.n4116 GND.n3167 585
R8473 GND.n4025 GND.n4024 585
R8474 GND.n4024 GND.n3165 585
R8475 GND.n4038 GND.n3176 585
R8476 GND.n4106 GND.n3176 585
R8477 GND.n4039 GND.n4023 585
R8478 GND.n4023 GND.n4022 585
R8479 GND.n4040 GND.n4020 585
R8480 GND.n4020 GND.n3182 585
R8481 GND.n4019 GND.n4017 585
R8482 GND.n4019 GND.n3187 585
R8483 GND.n4044 GND.n4016 585
R8484 GND.n4016 GND.n3193 585
R8485 GND.n4045 GND.n3199 585
R8486 GND.n4076 GND.n3199 585
R8487 GND.n4046 GND.n4015 585
R8488 GND.n4015 GND.n3197 585
R8489 GND.n3218 GND.n3208 585
R8490 GND.n4060 GND.n3208 585
R8491 GND.n4051 GND.n4050 585
R8492 GND.n4052 GND.n4051 585
R8493 GND.n3217 GND.n3216 585
R8494 GND.n3226 GND.n3216 585
R8495 GND.n4011 GND.n4010 585
R8496 GND.n4010 GND.n4009 585
R8497 GND.n3221 GND.n3220 585
R8498 GND.n3235 GND.n3221 585
R8499 GND.n3868 GND.n3233 585
R8500 GND.n3999 GND.n3233 585
R8501 GND.n3871 GND.n3867 585
R8502 GND.n3867 GND.n3241 585
R8503 GND.n3872 GND.n3866 585
R8504 GND.n3866 GND.n3248 585
R8505 GND.n3873 GND.n3253 585
R8506 GND.n3956 GND.n3253 585
R8507 GND.n3864 GND.n3863 585
R8508 GND.n3863 GND.n3862 585
R8509 GND.n3877 GND.n3262 585
R8510 GND.n3946 GND.n3262 585
R8511 GND.n3878 GND.n3861 585
R8512 GND.n3861 GND.n3270 585
R8513 GND.n3879 GND.n3860 585
R8514 GND.n3860 GND.n3269 585
R8515 GND.n3859 GND.n3857 585
R8516 GND.n3859 GND.n3275 585
R8517 GND.n3883 GND.n3856 585
R8518 GND.n3856 GND.n3282 585
R8519 GND.n3884 GND.n3288 585
R8520 GND.n3916 GND.n3288 585
R8521 GND.n3885 GND.n3855 585
R8522 GND.n3855 GND.n3286 585
R8523 GND.n3306 GND.n3296 585
R8524 GND.n3900 GND.n3296 585
R8525 GND.n3890 GND.n3889 585
R8526 GND.n3892 GND.n3890 585
R8527 GND.n3305 GND.n3304 585
R8528 GND.n3313 GND.n3304 585
R8529 GND.n3851 GND.n3850 585
R8530 GND.n3850 GND.n3849 585
R8531 GND.n3309 GND.n3308 585
R8532 GND.n3322 GND.n3309 585
R8533 GND.n3629 GND.n3320 585
R8534 GND.n3839 GND.n3320 585
R8535 GND.n3630 GND.n3628 585
R8536 GND.n3628 GND.n3327 585
R8537 GND.n3627 GND.n3625 585
R8538 GND.n3627 GND.n3334 585
R8539 GND.n3634 GND.n3341 585
R8540 GND.n3795 GND.n3341 585
R8541 GND.n3635 GND.n3624 585
R8542 GND.n3624 GND.n3339 585
R8543 GND.n3636 GND.n3350 585
R8544 GND.n3785 GND.n3350 585
R8545 GND.n3622 GND.n3621 585
R8546 GND.n3621 GND.n3357 585
R8547 GND.n3640 GND.n3620 585
R8548 GND.n3620 GND.n3356 585
R8549 GND.n3641 GND.n3619 585
R8550 GND.n3619 GND.n3363 585
R8551 GND.n3642 GND.n3618 585
R8552 GND.n3618 GND.n3369 585
R8553 GND.n3409 GND.n3379 585
R8554 GND.n3755 GND.n3379 585
R8555 GND.n3647 GND.n3646 585
R8556 GND.n3648 GND.n3647 585
R8557 GND.n3408 GND.n3387 585
R8558 GND.n3739 GND.n3387 585
R8559 GND.n3614 GND.n3613 585
R8560 GND.n3613 GND.n3386 585
R8561 GND.n3612 GND.n3411 585
R8562 GND.n3612 GND.n3611 585
R8563 GND.n3422 GND.n3412 585
R8564 GND.n3413 GND.n3412 585
R8565 GND.n3601 GND.n3600 585
R8566 GND.n3603 GND.n3601 585
R8567 GND.n3421 GND.n3420 585
R8568 GND.n3420 GND.n3419 585
R8569 GND.n3595 GND.n3594 585
R8570 GND.n3594 GND.n3593 585
R8571 GND.n3425 GND.n3424 585
R8572 GND.n3426 GND.n3425 585
R8573 GND.n3583 GND.n3582 585
R8574 GND.n3585 GND.n3583 585
R8575 GND.n3434 GND.n3433 585
R8576 GND.n3433 GND.n3432 585
R8577 GND.n3578 GND.n3577 585
R8578 GND.n3577 GND.n3576 585
R8579 GND.n3437 GND.n3436 585
R8580 GND.n3438 GND.n3437 585
R8581 GND.n3566 GND.n3565 585
R8582 GND.n3568 GND.n3566 585
R8583 GND.n3446 GND.n3445 585
R8584 GND.n3445 GND.n3444 585
R8585 GND.n3561 GND.n3560 585
R8586 GND.n3560 GND.n3559 585
R8587 GND.n3449 GND.n3448 585
R8588 GND.n3450 GND.n3449 585
R8589 GND.n3549 GND.n3548 585
R8590 GND.n3551 GND.n3549 585
R8591 GND.n3458 GND.n3457 585
R8592 GND.n3457 GND.n3456 585
R8593 GND.n3544 GND.n3543 585
R8594 GND.n3543 GND.n3542 585
R8595 GND.n3461 GND.n3460 585
R8596 GND.n3532 GND.n3461 585
R8597 GND.n3531 GND.n3530 585
R8598 GND.n3534 GND.n3531 585
R8599 GND.n3469 GND.n3468 585
R8600 GND.n3468 GND.n3467 585
R8601 GND.n3526 GND.n3525 585
R8602 GND.n3525 GND.n3524 585
R8603 GND.n3510 GND.n3471 585
R8604 GND.n3511 GND.n3510 585
R8605 GND.n3509 GND.n3508 585
R8606 GND.n3509 GND.n1534 585
R8607 GND.n3472 GND.n1533 585
R8608 GND.n5159 GND.n1533 585
R8609 GND.n4527 GND.n2493 585
R8610 GND.n4526 GND.n2904 585
R8611 GND.n4516 GND.n2903 585
R8612 GND.n4519 GND.n4518 585
R8613 GND.n2917 GND.n2914 585
R8614 GND.n2947 GND.n2946 585
R8615 GND.n2928 GND.n2927 585
R8616 GND.n2935 GND.n2934 585
R8617 GND.n2933 GND.n2514 585
R8618 GND.n4963 GND.n2513 585
R8619 GND.n4964 GND.n2512 585
R8620 GND.n4965 GND.n2511 585
R8621 GND.n2922 GND.n2509 585
R8622 GND.n4969 GND.n2508 585
R8623 GND.n4970 GND.n2507 585
R8624 GND.n4971 GND.n2506 585
R8625 GND.n2919 GND.n2504 585
R8626 GND.n4975 GND.n2503 585
R8627 GND.n4976 GND.n2502 585
R8628 GND.n4977 GND.n2498 585
R8629 GND.n4984 GND.n4983 585
R8630 GND.n4983 GND.n4982 585
R8631 GND.n4985 GND.n2492 585
R8632 GND.n2494 GND.n2492 585
R8633 GND.n4494 GND.n2490 585
R8634 GND.n4495 GND.n4494 585
R8635 GND.n4989 GND.n2489 585
R8636 GND.n2957 GND.n2489 585
R8637 GND.n4990 GND.n2488 585
R8638 GND.n4486 GND.n2488 585
R8639 GND.n4991 GND.n2487 585
R8640 GND.n2963 GND.n2487 585
R8641 GND.n4474 GND.n2485 585
R8642 GND.n4475 GND.n4474 585
R8643 GND.n4995 GND.n2484 585
R8644 GND.n2975 GND.n2484 585
R8645 GND.n4996 GND.n2483 585
R8646 GND.n4466 GND.n2483 585
R8647 GND.n4997 GND.n2482 585
R8648 GND.n2974 GND.n2482 585
R8649 GND.n4457 GND.n2480 585
R8650 GND.n4458 GND.n4457 585
R8651 GND.n5001 GND.n2479 585
R8652 GND.n2981 GND.n2479 585
R8653 GND.n5002 GND.n2478 585
R8654 GND.n4449 GND.n2478 585
R8655 GND.n5003 GND.n2477 585
R8656 GND.n2987 GND.n2477 585
R8657 GND.n4440 GND.n2475 585
R8658 GND.n4441 GND.n4440 585
R8659 GND.n5007 GND.n2474 585
R8660 GND.n2993 GND.n2474 585
R8661 GND.n5008 GND.n2473 585
R8662 GND.n4432 GND.n2473 585
R8663 GND.n5009 GND.n2472 585
R8664 GND.n2999 GND.n2472 585
R8665 GND.n4423 GND.n2470 585
R8666 GND.n4424 GND.n4423 585
R8667 GND.n5013 GND.n2469 585
R8668 GND.n3005 GND.n2469 585
R8669 GND.n5014 GND.n2468 585
R8670 GND.n4415 GND.n2468 585
R8671 GND.n5015 GND.n2467 585
R8672 GND.n3011 GND.n2467 585
R8673 GND.n4406 GND.n2465 585
R8674 GND.n4407 GND.n4406 585
R8675 GND.n5019 GND.n2464 585
R8676 GND.n3017 GND.n2464 585
R8677 GND.n5020 GND.n2463 585
R8678 GND.n4398 GND.n2463 585
R8679 GND.n5021 GND.n2462 585
R8680 GND.n3023 GND.n2462 585
R8681 GND.n4389 GND.n2460 585
R8682 GND.n4390 GND.n4389 585
R8683 GND.n5025 GND.n2459 585
R8684 GND.n4340 GND.n2459 585
R8685 GND.n5026 GND.n2458 585
R8686 GND.n3073 GND.n2458 585
R8687 GND.n5027 GND.n2457 585
R8688 GND.n4331 GND.n2457 585
R8689 GND.n3082 GND.n2455 585
R8690 GND.n3083 GND.n3082 585
R8691 GND.n5031 GND.n2454 585
R8692 GND.n4321 GND.n2454 585
R8693 GND.n5032 GND.n2453 585
R8694 GND.n4309 GND.n2453 585
R8695 GND.n5033 GND.n2452 585
R8696 GND.n3096 GND.n2452 585
R8697 GND.n3094 GND.n2450 585
R8698 GND.n3095 GND.n3094 585
R8699 GND.n5037 GND.n2449 585
R8700 GND.n3100 GND.n2449 585
R8701 GND.n5038 GND.n2448 585
R8702 GND.n3106 GND.n2448 585
R8703 GND.n5039 GND.n2447 585
R8704 GND.n4226 GND.n2447 585
R8705 GND.n3110 GND.n2445 585
R8706 GND.n3111 GND.n3110 585
R8707 GND.n5043 GND.n2444 585
R8708 GND.n4207 GND.n2444 585
R8709 GND.n5044 GND.n2443 585
R8710 GND.n4199 GND.n2443 585
R8711 GND.n5045 GND.n2442 585
R8712 GND.n3139 GND.n2442 585
R8713 GND.n3137 GND.n2440 585
R8714 GND.n4169 GND.n3137 585
R8715 GND.n5049 GND.n2439 585
R8716 GND.n3148 GND.n2439 585
R8717 GND.n5050 GND.n2438 585
R8718 GND.n4159 GND.n2438 585
R8719 GND.n5051 GND.n2437 585
R8720 GND.n3153 GND.n2437 585
R8721 GND.n3160 GND.n2435 585
R8722 GND.n3161 GND.n3160 585
R8723 GND.n5055 GND.n2434 585
R8724 GND.n4116 GND.n2434 585
R8725 GND.n5056 GND.n2433 585
R8726 GND.n3165 GND.n2433 585
R8727 GND.n5057 GND.n2432 585
R8728 GND.n4106 GND.n2432 585
R8729 GND.n4021 GND.n2430 585
R8730 GND.n4022 GND.n4021 585
R8731 GND.n5061 GND.n2429 585
R8732 GND.n3182 GND.n2429 585
R8733 GND.n5062 GND.n2428 585
R8734 GND.n3187 GND.n2428 585
R8735 GND.n5063 GND.n2427 585
R8736 GND.n3193 GND.n2427 585
R8737 GND.n3200 GND.n2425 585
R8738 GND.n4076 GND.n3200 585
R8739 GND.n5067 GND.n2424 585
R8740 GND.n3197 GND.n2424 585
R8741 GND.n5068 GND.n2423 585
R8742 GND.n4060 GND.n2423 585
R8743 GND.n5069 GND.n2422 585
R8744 GND.n4052 GND.n2422 585
R8745 GND.n3225 GND.n2420 585
R8746 GND.n3226 GND.n3225 585
R8747 GND.n5073 GND.n2419 585
R8748 GND.n4009 GND.n2419 585
R8749 GND.n5074 GND.n2418 585
R8750 GND.n3235 GND.n2418 585
R8751 GND.n5075 GND.n2417 585
R8752 GND.n3999 GND.n2417 585
R8753 GND.n3240 GND.n2415 585
R8754 GND.n3241 GND.n3240 585
R8755 GND.n5079 GND.n2414 585
R8756 GND.n3248 GND.n2414 585
R8757 GND.n5080 GND.n2413 585
R8758 GND.n3956 GND.n2413 585
R8759 GND.n5081 GND.n2412 585
R8760 GND.n3862 GND.n2412 585
R8761 GND.n3264 GND.n2410 585
R8762 GND.n3946 GND.n3264 585
R8763 GND.n5085 GND.n2409 585
R8764 GND.n3270 GND.n2409 585
R8765 GND.n5086 GND.n2408 585
R8766 GND.n3269 GND.n2408 585
R8767 GND.n5087 GND.n2407 585
R8768 GND.n3275 GND.n2407 585
R8769 GND.n3281 GND.n2405 585
R8770 GND.n3282 GND.n3281 585
R8771 GND.n5091 GND.n2404 585
R8772 GND.n3916 GND.n2404 585
R8773 GND.n5092 GND.n2403 585
R8774 GND.n3286 GND.n2403 585
R8775 GND.n5093 GND.n2402 585
R8776 GND.n3900 GND.n2402 585
R8777 GND.n3891 GND.n2400 585
R8778 GND.n3892 GND.n3891 585
R8779 GND.n5097 GND.n2399 585
R8780 GND.n3313 GND.n2399 585
R8781 GND.n5098 GND.n2398 585
R8782 GND.n3849 GND.n2398 585
R8783 GND.n5099 GND.n2397 585
R8784 GND.n3322 GND.n2397 585
R8785 GND.n3838 GND.n2395 585
R8786 GND.n3839 GND.n3838 585
R8787 GND.n5103 GND.n2394 585
R8788 GND.n3327 GND.n2394 585
R8789 GND.n5104 GND.n2393 585
R8790 GND.n3334 GND.n2393 585
R8791 GND.n5105 GND.n2392 585
R8792 GND.n3795 GND.n2392 585
R8793 GND.n3338 GND.n2390 585
R8794 GND.n3339 GND.n3338 585
R8795 GND.n5109 GND.n2389 585
R8796 GND.n3785 GND.n2389 585
R8797 GND.n5110 GND.n2388 585
R8798 GND.n3357 GND.n2388 585
R8799 GND.n5111 GND.n2387 585
R8800 GND.n3356 GND.n2387 585
R8801 GND.n3362 GND.n2385 585
R8802 GND.n3363 GND.n3362 585
R8803 GND.n5115 GND.n2384 585
R8804 GND.n3369 GND.n2384 585
R8805 GND.n5116 GND.n2383 585
R8806 GND.n3755 GND.n2383 585
R8807 GND.n5117 GND.n2382 585
R8808 GND.n3648 GND.n2382 585
R8809 GND.n3738 GND.n2380 585
R8810 GND.n3739 GND.n3738 585
R8811 GND.n5121 GND.n2379 585
R8812 GND.n3386 GND.n2379 585
R8813 GND.n5122 GND.n2378 585
R8814 GND.n3611 GND.n2378 585
R8815 GND.n5123 GND.n2377 585
R8816 GND.n3413 GND.n2377 585
R8817 GND.n3602 GND.n2375 585
R8818 GND.n3603 GND.n3602 585
R8819 GND.n5127 GND.n2374 585
R8820 GND.n3419 GND.n2374 585
R8821 GND.n5128 GND.n2373 585
R8822 GND.n3593 GND.n2373 585
R8823 GND.n5129 GND.n2372 585
R8824 GND.n3426 GND.n2372 585
R8825 GND.n3584 GND.n2370 585
R8826 GND.n3585 GND.n3584 585
R8827 GND.n5133 GND.n2369 585
R8828 GND.n3432 GND.n2369 585
R8829 GND.n5134 GND.n2368 585
R8830 GND.n3576 GND.n2368 585
R8831 GND.n5135 GND.n2367 585
R8832 GND.n3438 GND.n2367 585
R8833 GND.n3567 GND.n2365 585
R8834 GND.n3568 GND.n3567 585
R8835 GND.n5139 GND.n2364 585
R8836 GND.n3444 GND.n2364 585
R8837 GND.n5140 GND.n2363 585
R8838 GND.n3559 GND.n2363 585
R8839 GND.n5141 GND.n2362 585
R8840 GND.n3450 GND.n2362 585
R8841 GND.n3550 GND.n2360 585
R8842 GND.n3551 GND.n3550 585
R8843 GND.n5145 GND.n2359 585
R8844 GND.n3456 GND.n2359 585
R8845 GND.n5146 GND.n2358 585
R8846 GND.n3542 GND.n2358 585
R8847 GND.n5147 GND.n2357 585
R8848 GND.n3532 GND.n2357 585
R8849 GND.n3533 GND.n2355 585
R8850 GND.n3534 GND.n3533 585
R8851 GND.n5151 GND.n2354 585
R8852 GND.n3467 GND.n2354 585
R8853 GND.n5152 GND.n2353 585
R8854 GND.n3524 GND.n2353 585
R8855 GND.n5153 GND.n2352 585
R8856 GND.n3511 GND.n2352 585
R8857 GND.n1537 GND.n1536 585
R8858 GND.n1536 GND.n1534 585
R8859 GND.n5158 GND.n5157 585
R8860 GND.n5159 GND.n5158 585
R8861 GND.n5199 GND.n1490 585
R8862 GND.n5198 GND.n5197 585
R8863 GND.n1535 GND.n1497 585
R8864 GND.n5204 GND.n5201 585
R8865 GND.n3504 GND.n3474 585
R8866 GND.n3503 GND.n3476 585
R8867 GND.n3502 GND.n3477 585
R8868 GND.n3477 GND.n1495 585
R8869 GND.n3480 GND.n3478 585
R8870 GND.n3498 GND.n3482 585
R8871 GND.n3497 GND.n3483 585
R8872 GND.n3496 GND.n3485 585
R8873 GND.n3489 GND.n3486 585
R8874 GND.n3492 GND.n3491 585
R8875 GND.n3488 GND.n1472 585
R8876 GND.n5220 GND.n1473 585
R8877 GND.n5219 GND.n1474 585
R8878 GND.n1492 GND.n1475 585
R8879 GND.n5212 GND.n1482 585
R8880 GND.n5211 GND.n1483 585
R8881 GND.n1491 GND.n1484 585
R8882 GND.n1495 GND.n1491 585
R8883 GND.n5518 GND.n5517 483.755
R8884 GND.n4387 GND.n3053 482.89
R8885 GND.n4295 GND.n4294 482.89
R8886 GND.n3407 GND.n3378 482.89
R8887 GND.n3757 GND.n3377 482.89
R8888 GND.n6311 GND.n6310 401.031
R8889 GND.n6189 GND.n6188 301.784
R8890 GND.n6189 GND.n731 301.784
R8891 GND.n6197 GND.n731 301.784
R8892 GND.n6198 GND.n6197 301.784
R8893 GND.n6199 GND.n6198 301.784
R8894 GND.n6199 GND.n725 301.784
R8895 GND.n6207 GND.n725 301.784
R8896 GND.n6208 GND.n6207 301.784
R8897 GND.n6209 GND.n6208 301.784
R8898 GND.n6209 GND.n719 301.784
R8899 GND.n6217 GND.n719 301.784
R8900 GND.n6218 GND.n6217 301.784
R8901 GND.n6219 GND.n6218 301.784
R8902 GND.n6219 GND.n713 301.784
R8903 GND.n6227 GND.n713 301.784
R8904 GND.n6228 GND.n6227 301.784
R8905 GND.n6229 GND.n6228 301.784
R8906 GND.n6229 GND.n707 301.784
R8907 GND.n6237 GND.n707 301.784
R8908 GND.n6238 GND.n6237 301.784
R8909 GND.n6239 GND.n6238 301.784
R8910 GND.n6239 GND.n701 301.784
R8911 GND.n6247 GND.n701 301.784
R8912 GND.n6248 GND.n6247 301.784
R8913 GND.n6249 GND.n6248 301.784
R8914 GND.n6249 GND.n695 301.784
R8915 GND.n6257 GND.n695 301.784
R8916 GND.n6258 GND.n6257 301.784
R8917 GND.n6259 GND.n6258 301.784
R8918 GND.n6259 GND.n689 301.784
R8919 GND.n6267 GND.n689 301.784
R8920 GND.n6268 GND.n6267 301.784
R8921 GND.n6269 GND.n6268 301.784
R8922 GND.n6269 GND.n683 301.784
R8923 GND.n6277 GND.n683 301.784
R8924 GND.n6278 GND.n6277 301.784
R8925 GND.n6279 GND.n6278 301.784
R8926 GND.n6279 GND.n677 301.784
R8927 GND.n6287 GND.n677 301.784
R8928 GND.n6288 GND.n6287 301.784
R8929 GND.n6289 GND.n6288 301.784
R8930 GND.n6289 GND.n671 301.784
R8931 GND.n6297 GND.n671 301.784
R8932 GND.n6298 GND.n6297 301.784
R8933 GND.n6299 GND.n6298 301.784
R8934 GND.n6299 GND.n665 301.784
R8935 GND.n6309 GND.n665 301.784
R8936 GND.n6310 GND.n6309 301.784
R8937 GND.n135 GND.n129 289.615
R8938 GND.n148 GND.n142 289.615
R8939 GND.n109 GND.n103 289.615
R8940 GND.n122 GND.n116 289.615
R8941 GND.n83 GND.n77 289.615
R8942 GND.n96 GND.n90 289.615
R8943 GND.n57 GND.n51 289.615
R8944 GND.n70 GND.n64 289.615
R8945 GND.n31 GND.n25 289.615
R8946 GND.n44 GND.n38 289.615
R8947 GND.n6 GND.n0 289.615
R8948 GND.n19 GND.n13 289.615
R8949 GND.n304 GND.n298 289.615
R8950 GND.n291 GND.n285 289.615
R8951 GND.n278 GND.n272 289.615
R8952 GND.n265 GND.n259 289.615
R8953 GND.n252 GND.n246 289.615
R8954 GND.n239 GND.n233 289.615
R8955 GND.n226 GND.n220 289.615
R8956 GND.n213 GND.n207 289.615
R8957 GND.n200 GND.n194 289.615
R8958 GND.n187 GND.n181 289.615
R8959 GND.n175 GND.n169 289.615
R8960 GND.n162 GND.n156 289.615
R8961 GND.n5519 GND.n5518 280.613
R8962 GND.n5519 GND.n1133 280.613
R8963 GND.n5527 GND.n1133 280.613
R8964 GND.n5528 GND.n5527 280.613
R8965 GND.n5529 GND.n5528 280.613
R8966 GND.n5529 GND.n1127 280.613
R8967 GND.n5537 GND.n1127 280.613
R8968 GND.n5538 GND.n5537 280.613
R8969 GND.n5539 GND.n5538 280.613
R8970 GND.n5539 GND.n1121 280.613
R8971 GND.n5547 GND.n1121 280.613
R8972 GND.n5548 GND.n5547 280.613
R8973 GND.n5549 GND.n5548 280.613
R8974 GND.n5549 GND.n1115 280.613
R8975 GND.n5557 GND.n1115 280.613
R8976 GND.n5558 GND.n5557 280.613
R8977 GND.n5559 GND.n5558 280.613
R8978 GND.n5559 GND.n1109 280.613
R8979 GND.n5567 GND.n1109 280.613
R8980 GND.n5568 GND.n5567 280.613
R8981 GND.n5569 GND.n5568 280.613
R8982 GND.n5569 GND.n1103 280.613
R8983 GND.n5577 GND.n1103 280.613
R8984 GND.n5578 GND.n5577 280.613
R8985 GND.n5579 GND.n5578 280.613
R8986 GND.n5579 GND.n1097 280.613
R8987 GND.n5587 GND.n1097 280.613
R8988 GND.n5588 GND.n5587 280.613
R8989 GND.n5589 GND.n5588 280.613
R8990 GND.n5589 GND.n1091 280.613
R8991 GND.n5597 GND.n1091 280.613
R8992 GND.n5598 GND.n5597 280.613
R8993 GND.n5599 GND.n5598 280.613
R8994 GND.n5599 GND.n1085 280.613
R8995 GND.n5607 GND.n1085 280.613
R8996 GND.n5608 GND.n5607 280.613
R8997 GND.n5609 GND.n5608 280.613
R8998 GND.n5609 GND.n1079 280.613
R8999 GND.n5617 GND.n1079 280.613
R9000 GND.n5618 GND.n5617 280.613
R9001 GND.n5619 GND.n5618 280.613
R9002 GND.n5619 GND.n1073 280.613
R9003 GND.n5627 GND.n1073 280.613
R9004 GND.n5628 GND.n5627 280.613
R9005 GND.n5629 GND.n5628 280.613
R9006 GND.n5629 GND.n1067 280.613
R9007 GND.n5637 GND.n1067 280.613
R9008 GND.n5638 GND.n5637 280.613
R9009 GND.n5639 GND.n5638 280.613
R9010 GND.n5639 GND.n1061 280.613
R9011 GND.n5647 GND.n1061 280.613
R9012 GND.n5648 GND.n5647 280.613
R9013 GND.n5649 GND.n5648 280.613
R9014 GND.n5649 GND.n1055 280.613
R9015 GND.n5657 GND.n1055 280.613
R9016 GND.n5658 GND.n5657 280.613
R9017 GND.n5659 GND.n5658 280.613
R9018 GND.n5659 GND.n1049 280.613
R9019 GND.n5667 GND.n1049 280.613
R9020 GND.n5668 GND.n5667 280.613
R9021 GND.n5669 GND.n5668 280.613
R9022 GND.n5669 GND.n1043 280.613
R9023 GND.n5677 GND.n1043 280.613
R9024 GND.n5678 GND.n5677 280.613
R9025 GND.n5679 GND.n5678 280.613
R9026 GND.n5679 GND.n1037 280.613
R9027 GND.n5687 GND.n1037 280.613
R9028 GND.n5688 GND.n5687 280.613
R9029 GND.n5689 GND.n5688 280.613
R9030 GND.n5689 GND.n1031 280.613
R9031 GND.n5697 GND.n1031 280.613
R9032 GND.n5698 GND.n5697 280.613
R9033 GND.n5699 GND.n5698 280.613
R9034 GND.n5699 GND.n1025 280.613
R9035 GND.n5707 GND.n1025 280.613
R9036 GND.n5708 GND.n5707 280.613
R9037 GND.n5709 GND.n5708 280.613
R9038 GND.n5709 GND.n1019 280.613
R9039 GND.n5717 GND.n1019 280.613
R9040 GND.n5718 GND.n5717 280.613
R9041 GND.n5719 GND.n5718 280.613
R9042 GND.n5719 GND.n1013 280.613
R9043 GND.n5727 GND.n1013 280.613
R9044 GND.n5728 GND.n5727 280.613
R9045 GND.n5729 GND.n5728 280.613
R9046 GND.n5729 GND.n1007 280.613
R9047 GND.n5737 GND.n1007 280.613
R9048 GND.n5738 GND.n5737 280.613
R9049 GND.n5739 GND.n5738 280.613
R9050 GND.n5739 GND.n1001 280.613
R9051 GND.n5747 GND.n1001 280.613
R9052 GND.n5748 GND.n5747 280.613
R9053 GND.n5749 GND.n5748 280.613
R9054 GND.n5749 GND.n995 280.613
R9055 GND.n5757 GND.n995 280.613
R9056 GND.n5758 GND.n5757 280.613
R9057 GND.n5759 GND.n5758 280.613
R9058 GND.n5759 GND.n989 280.613
R9059 GND.n5767 GND.n989 280.613
R9060 GND.n5768 GND.n5767 280.613
R9061 GND.n5769 GND.n5768 280.613
R9062 GND.n5769 GND.n983 280.613
R9063 GND.n5777 GND.n983 280.613
R9064 GND.n5778 GND.n5777 280.613
R9065 GND.n5779 GND.n5778 280.613
R9066 GND.n5779 GND.n977 280.613
R9067 GND.n5787 GND.n977 280.613
R9068 GND.n5788 GND.n5787 280.613
R9069 GND.n5789 GND.n5788 280.613
R9070 GND.n5789 GND.n971 280.613
R9071 GND.n5797 GND.n971 280.613
R9072 GND.n5798 GND.n5797 280.613
R9073 GND.n5799 GND.n5798 280.613
R9074 GND.n5799 GND.n965 280.613
R9075 GND.n5807 GND.n965 280.613
R9076 GND.n5808 GND.n5807 280.613
R9077 GND.n5809 GND.n5808 280.613
R9078 GND.n5809 GND.n959 280.613
R9079 GND.n5817 GND.n959 280.613
R9080 GND.n5818 GND.n5817 280.613
R9081 GND.n5819 GND.n5818 280.613
R9082 GND.n5819 GND.n953 280.613
R9083 GND.n5827 GND.n953 280.613
R9084 GND.n5828 GND.n5827 280.613
R9085 GND.n5829 GND.n5828 280.613
R9086 GND.n5829 GND.n947 280.613
R9087 GND.n5837 GND.n947 280.613
R9088 GND.n5838 GND.n5837 280.613
R9089 GND.n5839 GND.n5838 280.613
R9090 GND.n5839 GND.n941 280.613
R9091 GND.n5847 GND.n941 280.613
R9092 GND.n5848 GND.n5847 280.613
R9093 GND.n5849 GND.n5848 280.613
R9094 GND.n5849 GND.n935 280.613
R9095 GND.n5857 GND.n935 280.613
R9096 GND.n5858 GND.n5857 280.613
R9097 GND.n5859 GND.n5858 280.613
R9098 GND.n5859 GND.n929 280.613
R9099 GND.n5867 GND.n929 280.613
R9100 GND.n5868 GND.n5867 280.613
R9101 GND.n5869 GND.n5868 280.613
R9102 GND.n5869 GND.n923 280.613
R9103 GND.n5877 GND.n923 280.613
R9104 GND.n5878 GND.n5877 280.613
R9105 GND.n5879 GND.n5878 280.613
R9106 GND.n5879 GND.n917 280.613
R9107 GND.n5887 GND.n917 280.613
R9108 GND.n5888 GND.n5887 280.613
R9109 GND.n5889 GND.n5888 280.613
R9110 GND.n5889 GND.n911 280.613
R9111 GND.n5897 GND.n911 280.613
R9112 GND.n5898 GND.n5897 280.613
R9113 GND.n5899 GND.n5898 280.613
R9114 GND.n5899 GND.n905 280.613
R9115 GND.n5907 GND.n905 280.613
R9116 GND.n5908 GND.n5907 280.613
R9117 GND.n5909 GND.n5908 280.613
R9118 GND.n5909 GND.n899 280.613
R9119 GND.n5917 GND.n899 280.613
R9120 GND.n5918 GND.n5917 280.613
R9121 GND.n5919 GND.n5918 280.613
R9122 GND.n5919 GND.n893 280.613
R9123 GND.n5927 GND.n893 280.613
R9124 GND.n5928 GND.n5927 280.613
R9125 GND.n5929 GND.n5928 280.613
R9126 GND.n5929 GND.n887 280.613
R9127 GND.n5937 GND.n887 280.613
R9128 GND.n5938 GND.n5937 280.613
R9129 GND.n5939 GND.n5938 280.613
R9130 GND.n5939 GND.n881 280.613
R9131 GND.n5947 GND.n881 280.613
R9132 GND.n5948 GND.n5947 280.613
R9133 GND.n5949 GND.n5948 280.613
R9134 GND.n5949 GND.n875 280.613
R9135 GND.n5957 GND.n875 280.613
R9136 GND.n5958 GND.n5957 280.613
R9137 GND.n5959 GND.n5958 280.613
R9138 GND.n5959 GND.n869 280.613
R9139 GND.n5967 GND.n869 280.613
R9140 GND.n5968 GND.n5967 280.613
R9141 GND.n5969 GND.n5968 280.613
R9142 GND.n5969 GND.n863 280.613
R9143 GND.n5977 GND.n863 280.613
R9144 GND.n5978 GND.n5977 280.613
R9145 GND.n5979 GND.n5978 280.613
R9146 GND.n5979 GND.n857 280.613
R9147 GND.n5987 GND.n857 280.613
R9148 GND.n5988 GND.n5987 280.613
R9149 GND.n5989 GND.n5988 280.613
R9150 GND.n5989 GND.n851 280.613
R9151 GND.n5997 GND.n851 280.613
R9152 GND.n5998 GND.n5997 280.613
R9153 GND.n5999 GND.n5998 280.613
R9154 GND.n5999 GND.n845 280.613
R9155 GND.n6007 GND.n845 280.613
R9156 GND.n6008 GND.n6007 280.613
R9157 GND.n6009 GND.n6008 280.613
R9158 GND.n6009 GND.n839 280.613
R9159 GND.n6017 GND.n839 280.613
R9160 GND.n6018 GND.n6017 280.613
R9161 GND.n6019 GND.n6018 280.613
R9162 GND.n6019 GND.n833 280.613
R9163 GND.n6027 GND.n833 280.613
R9164 GND.n6028 GND.n6027 280.613
R9165 GND.n6029 GND.n6028 280.613
R9166 GND.n6029 GND.n827 280.613
R9167 GND.n6037 GND.n827 280.613
R9168 GND.n6038 GND.n6037 280.613
R9169 GND.n6039 GND.n6038 280.613
R9170 GND.n6039 GND.n821 280.613
R9171 GND.n6047 GND.n821 280.613
R9172 GND.n6048 GND.n6047 280.613
R9173 GND.n6049 GND.n6048 280.613
R9174 GND.n6049 GND.n815 280.613
R9175 GND.n6057 GND.n815 280.613
R9176 GND.n6058 GND.n6057 280.613
R9177 GND.n6059 GND.n6058 280.613
R9178 GND.n6059 GND.n809 280.613
R9179 GND.n6067 GND.n809 280.613
R9180 GND.n6068 GND.n6067 280.613
R9181 GND.n6069 GND.n6068 280.613
R9182 GND.n6069 GND.n803 280.613
R9183 GND.n6077 GND.n803 280.613
R9184 GND.n6078 GND.n6077 280.613
R9185 GND.n6079 GND.n6078 280.613
R9186 GND.n6079 GND.n797 280.613
R9187 GND.n6087 GND.n797 280.613
R9188 GND.n6088 GND.n6087 280.613
R9189 GND.n6089 GND.n6088 280.613
R9190 GND.n6089 GND.n791 280.613
R9191 GND.n6097 GND.n791 280.613
R9192 GND.n6098 GND.n6097 280.613
R9193 GND.n6099 GND.n6098 280.613
R9194 GND.n6099 GND.n785 280.613
R9195 GND.n6107 GND.n785 280.613
R9196 GND.n6108 GND.n6107 280.613
R9197 GND.n6109 GND.n6108 280.613
R9198 GND.n6109 GND.n779 280.613
R9199 GND.n6117 GND.n779 280.613
R9200 GND.n6118 GND.n6117 280.613
R9201 GND.n6119 GND.n6118 280.613
R9202 GND.n6119 GND.n773 280.613
R9203 GND.n6127 GND.n773 280.613
R9204 GND.n6128 GND.n6127 280.613
R9205 GND.n6129 GND.n6128 280.613
R9206 GND.n6129 GND.n767 280.613
R9207 GND.n6137 GND.n767 280.613
R9208 GND.n6138 GND.n6137 280.613
R9209 GND.n6139 GND.n6138 280.613
R9210 GND.n6139 GND.n761 280.613
R9211 GND.n6147 GND.n761 280.613
R9212 GND.n6148 GND.n6147 280.613
R9213 GND.n6149 GND.n6148 280.613
R9214 GND.n6149 GND.n755 280.613
R9215 GND.n6157 GND.n755 280.613
R9216 GND.n6158 GND.n6157 280.613
R9217 GND.n6159 GND.n6158 280.613
R9218 GND.n6159 GND.n749 280.613
R9219 GND.n6167 GND.n749 280.613
R9220 GND.n6168 GND.n6167 280.613
R9221 GND.n6169 GND.n6168 280.613
R9222 GND.n6169 GND.n743 280.613
R9223 GND.n6177 GND.n743 280.613
R9224 GND.n6178 GND.n6177 280.613
R9225 GND.n6179 GND.n6178 280.613
R9226 GND.n6179 GND.n737 280.613
R9227 GND.n6187 GND.n737 280.613
R9228 GND.n2915 GND.t82 275.661
R9229 GND.n5202 GND.t90 275.661
R9230 GND.n3653 GND.t75 258.24
R9231 GND.n4252 GND.t49 258.24
R9232 GND.n3651 GND.t156 258.24
R9233 GND.n4346 GND.t140 258.24
R9234 GND.n3737 GND.n3736 256.663
R9235 GND.n3737 GND.n3388 256.663
R9236 GND.n3737 GND.n3389 256.663
R9237 GND.n3737 GND.n3390 256.663
R9238 GND.n3737 GND.n3391 256.663
R9239 GND.n3737 GND.n3392 256.663
R9240 GND.n3737 GND.n3393 256.663
R9241 GND.n3737 GND.n3394 256.663
R9242 GND.n3737 GND.n3395 256.663
R9243 GND.n3737 GND.n3396 256.663
R9244 GND.n3697 GND.n3696 256.663
R9245 GND.n3737 GND.n3397 256.663
R9246 GND.n3737 GND.n3398 256.663
R9247 GND.n3737 GND.n3399 256.663
R9248 GND.n3737 GND.n3400 256.663
R9249 GND.n3737 GND.n3401 256.663
R9250 GND.n3737 GND.n3402 256.663
R9251 GND.n3737 GND.n3403 256.663
R9252 GND.n3737 GND.n3404 256.663
R9253 GND.n3737 GND.n3405 256.663
R9254 GND.n3737 GND.n3406 256.663
R9255 GND.n4388 GND.n3041 256.663
R9256 GND.n4388 GND.n3040 256.663
R9257 GND.n4388 GND.n3039 256.663
R9258 GND.n4388 GND.n3038 256.663
R9259 GND.n4388 GND.n3037 256.663
R9260 GND.n4388 GND.n3036 256.663
R9261 GND.n4388 GND.n3035 256.663
R9262 GND.n4388 GND.n3034 256.663
R9263 GND.n4388 GND.n3033 256.663
R9264 GND.n4388 GND.n3032 256.663
R9265 GND.n3042 GND.n2576 256.663
R9266 GND.n4388 GND.n3043 256.663
R9267 GND.n4388 GND.n3044 256.663
R9268 GND.n4388 GND.n3045 256.663
R9269 GND.n4388 GND.n3046 256.663
R9270 GND.n4388 GND.n3047 256.663
R9271 GND.n4388 GND.n3048 256.663
R9272 GND.n4388 GND.n3049 256.663
R9273 GND.n4388 GND.n3050 256.663
R9274 GND.n4388 GND.n3051 256.663
R9275 GND.n4388 GND.n3052 256.663
R9276 GND.n1942 GND.n1267 242.672
R9277 GND.n1950 GND.n1267 242.672
R9278 GND.n1952 GND.n1267 242.672
R9279 GND.n1960 GND.n1267 242.672
R9280 GND.n5192 GND.n5191 242.672
R9281 GND.n5191 GND.n5170 242.672
R9282 GND.n5191 GND.n5172 242.672
R9283 GND.n5191 GND.n5173 242.672
R9284 GND.n4958 GND.n4957 242.672
R9285 GND.n4957 GND.n2547 242.672
R9286 GND.n4957 GND.n2546 242.672
R9287 GND.n4957 GND.n2545 242.672
R9288 GND.n4705 GND.n633 242.672
R9289 GND.n4680 GND.n633 242.672
R9290 GND.n4695 GND.n633 242.672
R9291 GND.n4684 GND.n633 242.672
R9292 GND.n1821 GND.n1267 242.672
R9293 GND.n1829 GND.n1267 242.672
R9294 GND.n1831 GND.n1267 242.672
R9295 GND.n1841 GND.n1267 242.672
R9296 GND.n1843 GND.n1267 242.672
R9297 GND.n1851 GND.n1267 242.672
R9298 GND.n1853 GND.n1267 242.672
R9299 GND.n1861 GND.n1267 242.672
R9300 GND.n1863 GND.n1267 242.672
R9301 GND.n1871 GND.n1267 242.672
R9302 GND.n1873 GND.n1267 242.672
R9303 GND.n1881 GND.n1267 242.672
R9304 GND.n1883 GND.n1267 242.672
R9305 GND.n1891 GND.n1267 242.672
R9306 GND.n1893 GND.n1267 242.672
R9307 GND.n1901 GND.n1267 242.672
R9308 GND.n1903 GND.n1267 242.672
R9309 GND.n1913 GND.n1267 242.672
R9310 GND.n1915 GND.n1267 242.672
R9311 GND.n1923 GND.n1267 242.672
R9312 GND.n1925 GND.n1267 242.672
R9313 GND.n1933 GND.n1267 242.672
R9314 GND.n5191 GND.n1523 242.672
R9315 GND.n5191 GND.n1522 242.672
R9316 GND.n5191 GND.n1521 242.672
R9317 GND.n5191 GND.n1519 242.672
R9318 GND.n5191 GND.n1518 242.672
R9319 GND.n5191 GND.n1516 242.672
R9320 GND.n5191 GND.n1515 242.672
R9321 GND.n5191 GND.n1513 242.672
R9322 GND.n5191 GND.n1512 242.672
R9323 GND.n5191 GND.n1510 242.672
R9324 GND.n5191 GND.n1509 242.672
R9325 GND.n5191 GND.n1507 242.672
R9326 GND.n5176 GND.n1432 242.672
R9327 GND.n5191 GND.n5177 242.672
R9328 GND.n5191 GND.n5178 242.672
R9329 GND.n5191 GND.n5180 242.672
R9330 GND.n5191 GND.n5181 242.672
R9331 GND.n5191 GND.n5183 242.672
R9332 GND.n5191 GND.n5184 242.672
R9333 GND.n5191 GND.n5186 242.672
R9334 GND.n5191 GND.n5187 242.672
R9335 GND.n5191 GND.n5189 242.672
R9336 GND.n5191 GND.n5190 242.672
R9337 GND.n4957 GND.n4956 242.672
R9338 GND.n4957 GND.n2521 242.672
R9339 GND.n4957 GND.n2522 242.672
R9340 GND.n4957 GND.n2523 242.672
R9341 GND.n4957 GND.n2524 242.672
R9342 GND.n4957 GND.n2525 242.672
R9343 GND.n4957 GND.n2526 242.672
R9344 GND.n4957 GND.n2527 242.672
R9345 GND.n4957 GND.n2528 242.672
R9346 GND.n4957 GND.n2529 242.672
R9347 GND.n4918 GND.n2577 242.672
R9348 GND.n4957 GND.n2530 242.672
R9349 GND.n4957 GND.n2531 242.672
R9350 GND.n4957 GND.n2532 242.672
R9351 GND.n4957 GND.n2533 242.672
R9352 GND.n4957 GND.n2534 242.672
R9353 GND.n4957 GND.n2535 242.672
R9354 GND.n4957 GND.n2536 242.672
R9355 GND.n4957 GND.n2537 242.672
R9356 GND.n4957 GND.n2538 242.672
R9357 GND.n4957 GND.n2539 242.672
R9358 GND.n4957 GND.n2540 242.672
R9359 GND.n4957 GND.n2541 242.672
R9360 GND.n633 GND.n632 242.672
R9361 GND.n633 GND.n482 242.672
R9362 GND.n633 GND.n481 242.672
R9363 GND.n633 GND.n480 242.672
R9364 GND.n633 GND.n479 242.672
R9365 GND.n633 GND.n478 242.672
R9366 GND.n633 GND.n477 242.672
R9367 GND.n633 GND.n476 242.672
R9368 GND.n633 GND.n475 242.672
R9369 GND.n633 GND.n474 242.672
R9370 GND.n633 GND.n473 242.672
R9371 GND.n633 GND.n472 242.672
R9372 GND.n633 GND.n471 242.672
R9373 GND.n633 GND.n470 242.672
R9374 GND.n633 GND.n469 242.672
R9375 GND.n633 GND.n468 242.672
R9376 GND.n633 GND.n467 242.672
R9377 GND.n633 GND.n466 242.672
R9378 GND.n633 GND.n465 242.672
R9379 GND.n633 GND.n464 242.672
R9380 GND.n633 GND.n463 242.672
R9381 GND.n633 GND.n462 242.672
R9382 GND.n633 GND.n461 242.672
R9383 GND.n4515 GND.n2949 242.672
R9384 GND.n4517 GND.n4515 242.672
R9385 GND.n4515 GND.n2948 242.672
R9386 GND.n4515 GND.n2926 242.672
R9387 GND.n4515 GND.n2925 242.672
R9388 GND.n4515 GND.n2924 242.672
R9389 GND.n4515 GND.n2923 242.672
R9390 GND.n4515 GND.n2921 242.672
R9391 GND.n4515 GND.n2920 242.672
R9392 GND.n4515 GND.n2918 242.672
R9393 GND.n5200 GND.n1495 242.672
R9394 GND.n1496 GND.n1495 242.672
R9395 GND.n3475 GND.n1495 242.672
R9396 GND.n3481 GND.n1495 242.672
R9397 GND.n3484 GND.n1495 242.672
R9398 GND.n3490 GND.n1495 242.672
R9399 GND.n3487 GND.n1495 242.672
R9400 GND.n1495 GND.n1493 242.672
R9401 GND.n1495 GND.n1494 242.672
R9402 GND.n529 GND.n528 240.244
R9403 GND.n532 GND.n531 240.244
R9404 GND.n539 GND.n538 240.244
R9405 GND.n519 GND.n518 240.244
R9406 GND.n547 GND.n546 240.244
R9407 GND.n550 GND.n549 240.244
R9408 GND.n557 GND.n556 240.244
R9409 GND.n560 GND.n559 240.244
R9410 GND.n567 GND.n566 240.244
R9411 GND.n570 GND.n569 240.244
R9412 GND.n577 GND.n576 240.244
R9413 GND.n580 GND.n579 240.244
R9414 GND.n587 GND.n586 240.244
R9415 GND.n591 GND.n590 240.244
R9416 GND.n597 GND.n596 240.244
R9417 GND.n601 GND.n600 240.244
R9418 GND.n607 GND.n606 240.244
R9419 GND.n611 GND.n610 240.244
R9420 GND.n614 GND.n613 240.244
R9421 GND.n621 GND.n620 240.244
R9422 GND.n624 GND.n623 240.244
R9423 GND.n631 GND.n483 240.244
R9424 GND.n4865 GND.n2611 240.244
R9425 GND.n4539 GND.n2611 240.244
R9426 GND.n4539 GND.n2625 240.244
R9427 GND.n4550 GND.n2625 240.244
R9428 GND.n4550 GND.n2644 240.244
R9429 GND.n4560 GND.n2644 240.244
R9430 GND.n4560 GND.n2656 240.244
R9431 GND.n4565 GND.n2656 240.244
R9432 GND.n4565 GND.n2667 240.244
R9433 GND.n4575 GND.n2667 240.244
R9434 GND.n4575 GND.n2677 240.244
R9435 GND.n4580 GND.n2677 240.244
R9436 GND.n4580 GND.n2688 240.244
R9437 GND.n4590 GND.n2688 240.244
R9438 GND.n4590 GND.n2698 240.244
R9439 GND.n4595 GND.n2698 240.244
R9440 GND.n4595 GND.n2709 240.244
R9441 GND.n4605 GND.n2709 240.244
R9442 GND.n4605 GND.n2719 240.244
R9443 GND.n4610 GND.n2719 240.244
R9444 GND.n4610 GND.n2728 240.244
R9445 GND.n4624 GND.n2728 240.244
R9446 GND.n4624 GND.n2738 240.244
R9447 GND.n2742 GND.n2738 240.244
R9448 GND.n2880 GND.n2742 240.244
R9449 GND.n2880 GND.n318 240.244
R9450 GND.n4635 GND.n318 240.244
R9451 GND.n4635 GND.n2873 240.244
R9452 GND.n4775 GND.n2873 240.244
R9453 GND.n4775 GND.n337 240.244
R9454 GND.n4767 GND.n337 240.244
R9455 GND.n4767 GND.n349 240.244
R9456 GND.n4763 GND.n349 240.244
R9457 GND.n4763 GND.n359 240.244
R9458 GND.n4755 GND.n359 240.244
R9459 GND.n4755 GND.n369 240.244
R9460 GND.n4751 GND.n369 240.244
R9461 GND.n4751 GND.n380 240.244
R9462 GND.n4743 GND.n380 240.244
R9463 GND.n4743 GND.n390 240.244
R9464 GND.n4739 GND.n390 240.244
R9465 GND.n4739 GND.n401 240.244
R9466 GND.n4731 GND.n401 240.244
R9467 GND.n4731 GND.n411 240.244
R9468 GND.n4727 GND.n411 240.244
R9469 GND.n4727 GND.n422 240.244
R9470 GND.n4719 GND.n422 240.244
R9471 GND.n4719 GND.n432 240.244
R9472 GND.n4715 GND.n432 240.244
R9473 GND.n4715 GND.n443 240.244
R9474 GND.n6351 GND.n443 240.244
R9475 GND.n2549 GND.n2548 240.244
R9476 GND.n4950 GND.n2548 240.244
R9477 GND.n4948 GND.n4947 240.244
R9478 GND.n4944 GND.n4943 240.244
R9479 GND.n4940 GND.n4939 240.244
R9480 GND.n4936 GND.n4935 240.244
R9481 GND.n4932 GND.n4931 240.244
R9482 GND.n4928 GND.n4927 240.244
R9483 GND.n4923 GND.n2569 240.244
R9484 GND.n4921 GND.n4920 240.244
R9485 GND.n4916 GND.n4915 240.244
R9486 GND.n4912 GND.n4911 240.244
R9487 GND.n4907 GND.n4906 240.244
R9488 GND.n4903 GND.n4902 240.244
R9489 GND.n4899 GND.n4898 240.244
R9490 GND.n4895 GND.n4894 240.244
R9491 GND.n4891 GND.n4890 240.244
R9492 GND.n4887 GND.n4886 240.244
R9493 GND.n4883 GND.n4882 240.244
R9494 GND.n4879 GND.n4878 240.244
R9495 GND.n4875 GND.n4874 240.244
R9496 GND.n2604 GND.n2542 240.244
R9497 GND.n2634 GND.n2550 240.244
R9498 GND.n2634 GND.n2629 240.244
R9499 GND.n4855 GND.n2629 240.244
R9500 GND.n4855 GND.n2630 240.244
R9501 GND.n4851 GND.n2630 240.244
R9502 GND.n4851 GND.n2642 240.244
R9503 GND.n4843 GND.n2642 240.244
R9504 GND.n4843 GND.n2659 240.244
R9505 GND.n4839 GND.n2659 240.244
R9506 GND.n4839 GND.n2665 240.244
R9507 GND.n4831 GND.n2665 240.244
R9508 GND.n4831 GND.n2680 240.244
R9509 GND.n4827 GND.n2680 240.244
R9510 GND.n4827 GND.n2686 240.244
R9511 GND.n4819 GND.n2686 240.244
R9512 GND.n4819 GND.n2701 240.244
R9513 GND.n4815 GND.n2701 240.244
R9514 GND.n4815 GND.n2707 240.244
R9515 GND.n4807 GND.n2707 240.244
R9516 GND.n4807 GND.n2722 240.244
R9517 GND.n4803 GND.n2722 240.244
R9518 GND.n4803 GND.n2726 240.244
R9519 GND.n4795 GND.n2726 240.244
R9520 GND.n4795 GND.n4794 240.244
R9521 GND.n4794 GND.n321 240.244
R9522 GND.n6423 GND.n321 240.244
R9523 GND.n6423 GND.n322 240.244
R9524 GND.n4782 GND.n322 240.244
R9525 GND.n4782 GND.n334 240.244
R9526 GND.n6418 GND.n334 240.244
R9527 GND.n6418 GND.n335 240.244
R9528 GND.n6410 GND.n335 240.244
R9529 GND.n6410 GND.n352 240.244
R9530 GND.n6406 GND.n352 240.244
R9531 GND.n6406 GND.n357 240.244
R9532 GND.n6398 GND.n357 240.244
R9533 GND.n6398 GND.n372 240.244
R9534 GND.n6394 GND.n372 240.244
R9535 GND.n6394 GND.n378 240.244
R9536 GND.n6386 GND.n378 240.244
R9537 GND.n6386 GND.n393 240.244
R9538 GND.n6382 GND.n393 240.244
R9539 GND.n6382 GND.n399 240.244
R9540 GND.n6374 GND.n399 240.244
R9541 GND.n6374 GND.n414 240.244
R9542 GND.n6370 GND.n414 240.244
R9543 GND.n6370 GND.n420 240.244
R9544 GND.n6362 GND.n420 240.244
R9545 GND.n6362 GND.n435 240.244
R9546 GND.n6358 GND.n435 240.244
R9547 GND.n6358 GND.n441 240.244
R9548 GND.n1405 GND.n1401 240.244
R9549 GND.n5188 GND.n1406 240.244
R9550 GND.n1410 GND.n1409 240.244
R9551 GND.n5185 GND.n1411 240.244
R9552 GND.n1417 GND.n1416 240.244
R9553 GND.n5182 GND.n1418 240.244
R9554 GND.n1422 GND.n1421 240.244
R9555 GND.n5179 GND.n1423 240.244
R9556 GND.n1429 GND.n1428 240.244
R9557 GND.n5175 GND.n1430 240.244
R9558 GND.n1506 GND.n1434 240.244
R9559 GND.n1436 GND.n1435 240.244
R9560 GND.n1508 GND.n1442 240.244
R9561 GND.n1444 GND.n1443 240.244
R9562 GND.n1511 GND.n1447 240.244
R9563 GND.n1449 GND.n1448 240.244
R9564 GND.n1514 GND.n1452 240.244
R9565 GND.n1456 GND.n1455 240.244
R9566 GND.n1517 GND.n1459 240.244
R9567 GND.n1461 GND.n1460 240.244
R9568 GND.n1520 GND.n1464 240.244
R9569 GND.n1469 GND.n1465 240.244
R9570 GND.n1754 GND.n1276 240.244
R9571 GND.n1754 GND.n1288 240.244
R9572 GND.n1298 GND.n1288 240.244
R9573 GND.n1299 GND.n1298 240.244
R9574 GND.n2003 GND.n1299 240.244
R9575 GND.n2003 GND.n1305 240.244
R9576 GND.n1306 GND.n1305 240.244
R9577 GND.n1307 GND.n1306 240.244
R9578 GND.n1735 GND.n1307 240.244
R9579 GND.n1735 GND.n1313 240.244
R9580 GND.n1314 GND.n1313 240.244
R9581 GND.n1315 GND.n1314 240.244
R9582 GND.n1720 GND.n1315 240.244
R9583 GND.n1720 GND.n1321 240.244
R9584 GND.n1322 GND.n1321 240.244
R9585 GND.n1323 GND.n1322 240.244
R9586 GND.n1694 GND.n1323 240.244
R9587 GND.n1694 GND.n1329 240.244
R9588 GND.n1330 GND.n1329 240.244
R9589 GND.n1331 GND.n1330 240.244
R9590 GND.n1645 GND.n1331 240.244
R9591 GND.n1645 GND.n1337 240.244
R9592 GND.n1338 GND.n1337 240.244
R9593 GND.n1339 GND.n1338 240.244
R9594 GND.n1660 GND.n1339 240.244
R9595 GND.n1660 GND.n1345 240.244
R9596 GND.n1346 GND.n1345 240.244
R9597 GND.n1347 GND.n1346 240.244
R9598 GND.n2138 GND.n1347 240.244
R9599 GND.n2138 GND.n1353 240.244
R9600 GND.n1354 GND.n1353 240.244
R9601 GND.n1355 GND.n1354 240.244
R9602 GND.n1615 GND.n1355 240.244
R9603 GND.n1615 GND.n1361 240.244
R9604 GND.n1362 GND.n1361 240.244
R9605 GND.n1363 GND.n1362 240.244
R9606 GND.n1596 GND.n1363 240.244
R9607 GND.n1596 GND.n1369 240.244
R9608 GND.n1370 GND.n1369 240.244
R9609 GND.n1371 GND.n1370 240.244
R9610 GND.n1584 GND.n1371 240.244
R9611 GND.n1584 GND.n1377 240.244
R9612 GND.n1378 GND.n1377 240.244
R9613 GND.n1379 GND.n1378 240.244
R9614 GND.n1562 GND.n1379 240.244
R9615 GND.n1562 GND.n1385 240.244
R9616 GND.n1386 GND.n1385 240.244
R9617 GND.n1387 GND.n1386 240.244
R9618 GND.n1544 GND.n1387 240.244
R9619 GND.n1544 GND.n1393 240.244
R9620 GND.n5295 GND.n1393 240.244
R9621 GND.n1822 GND.n1817 240.244
R9622 GND.n1828 GND.n1817 240.244
R9623 GND.n1832 GND.n1830 240.244
R9624 GND.n1840 GND.n1813 240.244
R9625 GND.n1844 GND.n1842 240.244
R9626 GND.n1850 GND.n1809 240.244
R9627 GND.n1854 GND.n1852 240.244
R9628 GND.n1860 GND.n1805 240.244
R9629 GND.n1864 GND.n1862 240.244
R9630 GND.n1870 GND.n1799 240.244
R9631 GND.n1874 GND.n1872 240.244
R9632 GND.n1880 GND.n1795 240.244
R9633 GND.n1884 GND.n1882 240.244
R9634 GND.n1890 GND.n1788 240.244
R9635 GND.n1894 GND.n1892 240.244
R9636 GND.n1900 GND.n1784 240.244
R9637 GND.n1904 GND.n1902 240.244
R9638 GND.n1912 GND.n1780 240.244
R9639 GND.n1916 GND.n1914 240.244
R9640 GND.n1922 GND.n1776 240.244
R9641 GND.n1926 GND.n1924 240.244
R9642 GND.n1932 GND.n1772 240.244
R9643 GND.n1935 GND.n1934 240.244
R9644 GND.n5378 GND.n1281 240.244
R9645 GND.n5374 GND.n1281 240.244
R9646 GND.n5374 GND.n1286 240.244
R9647 GND.n2011 GND.n1286 240.244
R9648 GND.n2011 GND.n2005 240.244
R9649 GND.n2005 GND.n1744 240.244
R9650 GND.n2028 GND.n1744 240.244
R9651 GND.n2028 GND.n1739 240.244
R9652 GND.n2036 GND.n1739 240.244
R9653 GND.n2036 GND.n1740 240.244
R9654 GND.n1740 GND.n1714 240.244
R9655 GND.n2081 GND.n1714 240.244
R9656 GND.n2081 GND.n1708 240.244
R9657 GND.n2089 GND.n1708 240.244
R9658 GND.n2089 GND.n1710 240.244
R9659 GND.n1710 GND.n1692 240.244
R9660 GND.n2105 GND.n1692 240.244
R9661 GND.n2105 GND.n1688 240.244
R9662 GND.n2111 GND.n1688 240.244
R9663 GND.n2111 GND.n1642 240.244
R9664 GND.n2212 GND.n1642 240.244
R9665 GND.n2212 GND.n1643 240.244
R9666 GND.n1665 GND.n1643 240.244
R9667 GND.n1667 GND.n1665 240.244
R9668 GND.n2198 GND.n1667 240.244
R9669 GND.n2198 GND.n2195 240.244
R9670 GND.n2195 GND.n1668 240.244
R9671 GND.n2135 GND.n1668 240.244
R9672 GND.n2135 GND.n1630 240.244
R9673 GND.n2219 GND.n1630 240.244
R9674 GND.n2219 GND.n1632 240.244
R9675 GND.n1632 GND.n1613 240.244
R9676 GND.n2235 GND.n1613 240.244
R9677 GND.n2235 GND.n1607 240.244
R9678 GND.n2243 GND.n1607 240.244
R9679 GND.n2243 GND.n1609 240.244
R9680 GND.n1609 GND.n1590 240.244
R9681 GND.n2260 GND.n1590 240.244
R9682 GND.n2260 GND.n1583 240.244
R9683 GND.n2268 GND.n1583 240.244
R9684 GND.n2268 GND.n1586 240.244
R9685 GND.n1586 GND.n1568 240.244
R9686 GND.n2298 GND.n1568 240.244
R9687 GND.n2298 GND.n1564 240.244
R9688 GND.n2304 GND.n1564 240.244
R9689 GND.n2304 GND.n1549 240.244
R9690 GND.n2335 GND.n1549 240.244
R9691 GND.n2335 GND.n1545 240.244
R9692 GND.n2341 GND.n1545 240.244
R9693 GND.n2341 GND.n1400 240.244
R9694 GND.n5293 GND.n1400 240.244
R9695 GND.n4687 GND.n4686 240.244
R9696 GND.n4694 GND.n4693 240.244
R9697 GND.n4697 GND.n4696 240.244
R9698 GND.n4704 GND.n4703 240.244
R9699 GND.n4534 GND.n2613 240.244
R9700 GND.n4535 GND.n4534 240.244
R9701 GND.n4535 GND.n2626 240.244
R9702 GND.n4552 GND.n2626 240.244
R9703 GND.n4552 GND.n2645 240.244
R9704 GND.n4558 GND.n2645 240.244
R9705 GND.n4558 GND.n2657 240.244
R9706 GND.n4567 GND.n2657 240.244
R9707 GND.n4567 GND.n2668 240.244
R9708 GND.n4573 GND.n2668 240.244
R9709 GND.n4573 GND.n2678 240.244
R9710 GND.n4582 GND.n2678 240.244
R9711 GND.n4582 GND.n2689 240.244
R9712 GND.n4588 GND.n2689 240.244
R9713 GND.n4588 GND.n2699 240.244
R9714 GND.n4597 GND.n2699 240.244
R9715 GND.n4597 GND.n2710 240.244
R9716 GND.n4603 GND.n2710 240.244
R9717 GND.n4603 GND.n2720 240.244
R9718 GND.n4612 GND.n2720 240.244
R9719 GND.n4612 GND.n2729 240.244
R9720 GND.n4622 GND.n2729 240.244
R9721 GND.n4622 GND.n2739 240.244
R9722 GND.n2743 GND.n2739 240.244
R9723 GND.n2743 GND.n315 240.244
R9724 GND.n6425 GND.n315 240.244
R9725 GND.n6425 GND.n316 240.244
R9726 GND.n2874 GND.n316 240.244
R9727 GND.n4773 GND.n2874 240.244
R9728 GND.n4773 GND.n338 240.244
R9729 GND.n4769 GND.n338 240.244
R9730 GND.n4769 GND.n350 240.244
R9731 GND.n4761 GND.n350 240.244
R9732 GND.n4761 GND.n360 240.244
R9733 GND.n4757 GND.n360 240.244
R9734 GND.n4757 GND.n370 240.244
R9735 GND.n4749 GND.n370 240.244
R9736 GND.n4749 GND.n381 240.244
R9737 GND.n4745 GND.n381 240.244
R9738 GND.n4745 GND.n391 240.244
R9739 GND.n4737 GND.n391 240.244
R9740 GND.n4737 GND.n402 240.244
R9741 GND.n4733 GND.n402 240.244
R9742 GND.n4733 GND.n412 240.244
R9743 GND.n4725 GND.n412 240.244
R9744 GND.n4725 GND.n423 240.244
R9745 GND.n4721 GND.n423 240.244
R9746 GND.n4721 GND.n433 240.244
R9747 GND.n4713 GND.n433 240.244
R9748 GND.n4713 GND.n444 240.244
R9749 GND.n451 GND.n444 240.244
R9750 GND.n2931 GND.n2519 240.244
R9751 GND.n2942 GND.n2941 240.244
R9752 GND.n2912 GND.n2911 240.244
R9753 GND.n2907 GND.n2544 240.244
R9754 GND.n4543 GND.n2518 240.244
R9755 GND.n4544 GND.n4543 240.244
R9756 GND.n4544 GND.n2628 240.244
R9757 GND.n2647 GND.n2628 240.244
R9758 GND.n4849 GND.n2647 240.244
R9759 GND.n4849 GND.n2648 240.244
R9760 GND.n4845 GND.n2648 240.244
R9761 GND.n4845 GND.n2654 240.244
R9762 GND.n4837 GND.n2654 240.244
R9763 GND.n4837 GND.n2670 240.244
R9764 GND.n4833 GND.n2670 240.244
R9765 GND.n4833 GND.n2675 240.244
R9766 GND.n4825 GND.n2675 240.244
R9767 GND.n4825 GND.n2691 240.244
R9768 GND.n4821 GND.n2691 240.244
R9769 GND.n4821 GND.n2696 240.244
R9770 GND.n4813 GND.n2696 240.244
R9771 GND.n4813 GND.n2712 240.244
R9772 GND.n4809 GND.n2712 240.244
R9773 GND.n4809 GND.n2717 240.244
R9774 GND.n4801 GND.n2717 240.244
R9775 GND.n4801 GND.n2731 240.244
R9776 GND.n4797 GND.n2731 240.244
R9777 GND.n4797 GND.n2736 240.244
R9778 GND.n4630 GND.n2736 240.244
R9779 GND.n4630 GND.n320 240.244
R9780 GND.n2876 GND.n320 240.244
R9781 GND.n4780 GND.n2876 240.244
R9782 GND.n4780 GND.n340 240.244
R9783 GND.n6416 GND.n340 240.244
R9784 GND.n6416 GND.n341 240.244
R9785 GND.n6412 GND.n341 240.244
R9786 GND.n6412 GND.n347 240.244
R9787 GND.n6404 GND.n347 240.244
R9788 GND.n6404 GND.n362 240.244
R9789 GND.n6400 GND.n362 240.244
R9790 GND.n6400 GND.n367 240.244
R9791 GND.n6392 GND.n367 240.244
R9792 GND.n6392 GND.n383 240.244
R9793 GND.n6388 GND.n383 240.244
R9794 GND.n6388 GND.n388 240.244
R9795 GND.n6380 GND.n388 240.244
R9796 GND.n6380 GND.n404 240.244
R9797 GND.n6376 GND.n404 240.244
R9798 GND.n6376 GND.n409 240.244
R9799 GND.n6368 GND.n409 240.244
R9800 GND.n6368 GND.n425 240.244
R9801 GND.n6364 GND.n425 240.244
R9802 GND.n6364 GND.n430 240.244
R9803 GND.n6356 GND.n430 240.244
R9804 GND.n6356 GND.n446 240.244
R9805 GND.n5174 GND.n1478 240.244
R9806 GND.n5171 GND.n1479 240.244
R9807 GND.n1487 GND.n1486 240.244
R9808 GND.n5169 GND.n1504 240.244
R9809 GND.n1756 GND.n1277 240.244
R9810 GND.n1756 GND.n1289 240.244
R9811 GND.n1971 GND.n1289 240.244
R9812 GND.n2013 GND.n1971 240.244
R9813 GND.n2013 GND.n1750 240.244
R9814 GND.n2020 GND.n1750 240.244
R9815 GND.n2020 GND.n1746 240.244
R9816 GND.n1746 GND.n1733 240.244
R9817 GND.n2038 GND.n1733 240.244
R9818 GND.n2038 GND.n1728 240.244
R9819 GND.n2045 GND.n1728 240.244
R9820 GND.n2045 GND.n1716 240.244
R9821 GND.n1716 GND.n1705 240.244
R9822 GND.n2091 GND.n1705 240.244
R9823 GND.n2091 GND.n1700 240.244
R9824 GND.n2098 GND.n1700 240.244
R9825 GND.n2098 GND.n1695 240.244
R9826 GND.n1695 GND.n1681 240.244
R9827 GND.n2113 GND.n1681 240.244
R9828 GND.n2113 GND.n1682 240.244
R9829 GND.n1682 GND.n1646 240.244
R9830 GND.n1651 GND.n1646 240.244
R9831 GND.n2121 GND.n1651 240.244
R9832 GND.n2121 GND.n2120 240.244
R9833 GND.n2120 GND.n1661 240.244
R9834 GND.n1669 GND.n1661 240.244
R9835 GND.n1673 GND.n1669 240.244
R9836 GND.n2132 GND.n1673 240.244
R9837 GND.n2132 GND.n1626 240.244
R9838 GND.n2221 GND.n1626 240.244
R9839 GND.n2221 GND.n1621 240.244
R9840 GND.n2228 GND.n1621 240.244
R9841 GND.n2228 GND.n1616 240.244
R9842 GND.n1616 GND.n1602 240.244
R9843 GND.n2245 GND.n1602 240.244
R9844 GND.n2245 GND.n1597 240.244
R9845 GND.n2252 GND.n1597 240.244
R9846 GND.n2252 GND.n1592 240.244
R9847 GND.n1592 GND.n1579 240.244
R9848 GND.n2270 GND.n1579 240.244
R9849 GND.n2270 GND.n1574 240.244
R9850 GND.n2291 GND.n1574 240.244
R9851 GND.n2291 GND.n1570 240.244
R9852 GND.n2275 GND.n1570 240.244
R9853 GND.n2275 GND.n1563 240.244
R9854 GND.n1563 GND.n1554 240.244
R9855 GND.n1554 GND.n1550 240.244
R9856 GND.n2279 GND.n1550 240.244
R9857 GND.n2279 GND.n1540 240.244
R9858 GND.n2346 GND.n1540 240.244
R9859 GND.n2346 GND.n1396 240.244
R9860 GND.n1949 GND.n1766 240.244
R9861 GND.n1953 GND.n1951 240.244
R9862 GND.n1959 GND.n1762 240.244
R9863 GND.n1962 GND.n1961 240.244
R9864 GND.n1291 GND.n1279 240.244
R9865 GND.n5372 GND.n1291 240.244
R9866 GND.n5372 GND.n1292 240.244
R9867 GND.n1974 GND.n1292 240.244
R9868 GND.n1974 GND.n1748 240.244
R9869 GND.n2022 GND.n1748 240.244
R9870 GND.n2026 GND.n2022 240.244
R9871 GND.n2026 GND.n2024 240.244
R9872 GND.n2024 GND.n1738 240.244
R9873 GND.n1738 GND.n1737 240.244
R9874 GND.n1737 GND.n1719 240.244
R9875 GND.n2079 GND.n1719 240.244
R9876 GND.n2079 GND.n2078 240.244
R9877 GND.n2078 GND.n1707 240.244
R9878 GND.n1707 GND.n1698 240.244
R9879 GND.n2100 GND.n1698 240.244
R9880 GND.n2103 GND.n2100 240.244
R9881 GND.n2103 GND.n2102 240.244
R9882 GND.n2102 GND.n1687 240.244
R9883 GND.n1687 GND.n1648 240.244
R9884 GND.n2210 GND.n1648 240.244
R9885 GND.n2210 GND.n2209 240.244
R9886 GND.n2209 GND.n1650 240.244
R9887 GND.n1663 GND.n1650 240.244
R9888 GND.n1664 GND.n1663 240.244
R9889 GND.n2193 GND.n1664 240.244
R9890 GND.n2193 GND.n2192 240.244
R9891 GND.n2192 GND.n1671 240.244
R9892 GND.n2139 GND.n1671 240.244
R9893 GND.n2139 GND.n1629 240.244
R9894 GND.n1629 GND.n1619 240.244
R9895 GND.n2230 GND.n1619 240.244
R9896 GND.n2233 GND.n2230 240.244
R9897 GND.n2233 GND.n2232 240.244
R9898 GND.n2232 GND.n1606 240.244
R9899 GND.n1606 GND.n1594 240.244
R9900 GND.n2254 GND.n1594 240.244
R9901 GND.n2258 GND.n2254 240.244
R9902 GND.n2258 GND.n2257 240.244
R9903 GND.n2257 GND.n1582 240.244
R9904 GND.n1582 GND.n1572 240.244
R9905 GND.n2293 GND.n1572 240.244
R9906 GND.n2296 GND.n2293 240.244
R9907 GND.n2296 GND.n2294 240.244
R9908 GND.n2294 GND.n1552 240.244
R9909 GND.n2331 GND.n1552 240.244
R9910 GND.n2333 GND.n2331 240.244
R9911 GND.n2333 GND.n1542 240.244
R9912 GND.n2343 GND.n1542 240.244
R9913 GND.n2344 GND.n2343 240.244
R9914 GND.n2344 GND.n1399 240.244
R9915 GND.n5520 GND.n1138 240.244
R9916 GND.n5520 GND.n1134 240.244
R9917 GND.n5526 GND.n1134 240.244
R9918 GND.n5526 GND.n1132 240.244
R9919 GND.n5530 GND.n1132 240.244
R9920 GND.n5530 GND.n1128 240.244
R9921 GND.n5536 GND.n1128 240.244
R9922 GND.n5536 GND.n1126 240.244
R9923 GND.n5540 GND.n1126 240.244
R9924 GND.n5540 GND.n1122 240.244
R9925 GND.n5546 GND.n1122 240.244
R9926 GND.n5546 GND.n1120 240.244
R9927 GND.n5550 GND.n1120 240.244
R9928 GND.n5550 GND.n1116 240.244
R9929 GND.n5556 GND.n1116 240.244
R9930 GND.n5556 GND.n1114 240.244
R9931 GND.n5560 GND.n1114 240.244
R9932 GND.n5560 GND.n1110 240.244
R9933 GND.n5566 GND.n1110 240.244
R9934 GND.n5566 GND.n1108 240.244
R9935 GND.n5570 GND.n1108 240.244
R9936 GND.n5570 GND.n1104 240.244
R9937 GND.n5576 GND.n1104 240.244
R9938 GND.n5576 GND.n1102 240.244
R9939 GND.n5580 GND.n1102 240.244
R9940 GND.n5580 GND.n1098 240.244
R9941 GND.n5586 GND.n1098 240.244
R9942 GND.n5586 GND.n1096 240.244
R9943 GND.n5590 GND.n1096 240.244
R9944 GND.n5590 GND.n1092 240.244
R9945 GND.n5596 GND.n1092 240.244
R9946 GND.n5596 GND.n1090 240.244
R9947 GND.n5600 GND.n1090 240.244
R9948 GND.n5600 GND.n1086 240.244
R9949 GND.n5606 GND.n1086 240.244
R9950 GND.n5606 GND.n1084 240.244
R9951 GND.n5610 GND.n1084 240.244
R9952 GND.n5610 GND.n1080 240.244
R9953 GND.n5616 GND.n1080 240.244
R9954 GND.n5616 GND.n1078 240.244
R9955 GND.n5620 GND.n1078 240.244
R9956 GND.n5620 GND.n1074 240.244
R9957 GND.n5626 GND.n1074 240.244
R9958 GND.n5626 GND.n1072 240.244
R9959 GND.n5630 GND.n1072 240.244
R9960 GND.n5630 GND.n1068 240.244
R9961 GND.n5636 GND.n1068 240.244
R9962 GND.n5636 GND.n1066 240.244
R9963 GND.n5640 GND.n1066 240.244
R9964 GND.n5640 GND.n1062 240.244
R9965 GND.n5646 GND.n1062 240.244
R9966 GND.n5646 GND.n1060 240.244
R9967 GND.n5650 GND.n1060 240.244
R9968 GND.n5650 GND.n1056 240.244
R9969 GND.n5656 GND.n1056 240.244
R9970 GND.n5656 GND.n1054 240.244
R9971 GND.n5660 GND.n1054 240.244
R9972 GND.n5660 GND.n1050 240.244
R9973 GND.n5666 GND.n1050 240.244
R9974 GND.n5666 GND.n1048 240.244
R9975 GND.n5670 GND.n1048 240.244
R9976 GND.n5670 GND.n1044 240.244
R9977 GND.n5676 GND.n1044 240.244
R9978 GND.n5676 GND.n1042 240.244
R9979 GND.n5680 GND.n1042 240.244
R9980 GND.n5680 GND.n1038 240.244
R9981 GND.n5686 GND.n1038 240.244
R9982 GND.n5686 GND.n1036 240.244
R9983 GND.n5690 GND.n1036 240.244
R9984 GND.n5690 GND.n1032 240.244
R9985 GND.n5696 GND.n1032 240.244
R9986 GND.n5696 GND.n1030 240.244
R9987 GND.n5700 GND.n1030 240.244
R9988 GND.n5700 GND.n1026 240.244
R9989 GND.n5706 GND.n1026 240.244
R9990 GND.n5706 GND.n1024 240.244
R9991 GND.n5710 GND.n1024 240.244
R9992 GND.n5710 GND.n1020 240.244
R9993 GND.n5716 GND.n1020 240.244
R9994 GND.n5716 GND.n1018 240.244
R9995 GND.n5720 GND.n1018 240.244
R9996 GND.n5720 GND.n1014 240.244
R9997 GND.n5726 GND.n1014 240.244
R9998 GND.n5726 GND.n1012 240.244
R9999 GND.n5730 GND.n1012 240.244
R10000 GND.n5730 GND.n1008 240.244
R10001 GND.n5736 GND.n1008 240.244
R10002 GND.n5736 GND.n1006 240.244
R10003 GND.n5740 GND.n1006 240.244
R10004 GND.n5740 GND.n1002 240.244
R10005 GND.n5746 GND.n1002 240.244
R10006 GND.n5746 GND.n1000 240.244
R10007 GND.n5750 GND.n1000 240.244
R10008 GND.n5750 GND.n996 240.244
R10009 GND.n5756 GND.n996 240.244
R10010 GND.n5756 GND.n994 240.244
R10011 GND.n5760 GND.n994 240.244
R10012 GND.n5760 GND.n990 240.244
R10013 GND.n5766 GND.n990 240.244
R10014 GND.n5766 GND.n988 240.244
R10015 GND.n5770 GND.n988 240.244
R10016 GND.n5770 GND.n984 240.244
R10017 GND.n5776 GND.n984 240.244
R10018 GND.n5776 GND.n982 240.244
R10019 GND.n5780 GND.n982 240.244
R10020 GND.n5780 GND.n978 240.244
R10021 GND.n5786 GND.n978 240.244
R10022 GND.n5786 GND.n976 240.244
R10023 GND.n5790 GND.n976 240.244
R10024 GND.n5790 GND.n972 240.244
R10025 GND.n5796 GND.n972 240.244
R10026 GND.n5796 GND.n970 240.244
R10027 GND.n5800 GND.n970 240.244
R10028 GND.n5800 GND.n966 240.244
R10029 GND.n5806 GND.n966 240.244
R10030 GND.n5806 GND.n964 240.244
R10031 GND.n5810 GND.n964 240.244
R10032 GND.n5810 GND.n960 240.244
R10033 GND.n5816 GND.n960 240.244
R10034 GND.n5816 GND.n958 240.244
R10035 GND.n5820 GND.n958 240.244
R10036 GND.n5820 GND.n954 240.244
R10037 GND.n5826 GND.n954 240.244
R10038 GND.n5826 GND.n952 240.244
R10039 GND.n5830 GND.n952 240.244
R10040 GND.n5830 GND.n948 240.244
R10041 GND.n5836 GND.n948 240.244
R10042 GND.n5836 GND.n946 240.244
R10043 GND.n5840 GND.n946 240.244
R10044 GND.n5840 GND.n942 240.244
R10045 GND.n5846 GND.n942 240.244
R10046 GND.n5846 GND.n940 240.244
R10047 GND.n5850 GND.n940 240.244
R10048 GND.n5850 GND.n936 240.244
R10049 GND.n5856 GND.n936 240.244
R10050 GND.n5856 GND.n934 240.244
R10051 GND.n5860 GND.n934 240.244
R10052 GND.n5860 GND.n930 240.244
R10053 GND.n5866 GND.n930 240.244
R10054 GND.n5866 GND.n928 240.244
R10055 GND.n5870 GND.n928 240.244
R10056 GND.n5870 GND.n924 240.244
R10057 GND.n5876 GND.n924 240.244
R10058 GND.n5876 GND.n922 240.244
R10059 GND.n5880 GND.n922 240.244
R10060 GND.n5880 GND.n918 240.244
R10061 GND.n5886 GND.n918 240.244
R10062 GND.n5886 GND.n916 240.244
R10063 GND.n5890 GND.n916 240.244
R10064 GND.n5890 GND.n912 240.244
R10065 GND.n5896 GND.n912 240.244
R10066 GND.n5896 GND.n910 240.244
R10067 GND.n5900 GND.n910 240.244
R10068 GND.n5900 GND.n906 240.244
R10069 GND.n5906 GND.n906 240.244
R10070 GND.n5906 GND.n904 240.244
R10071 GND.n5910 GND.n904 240.244
R10072 GND.n5910 GND.n900 240.244
R10073 GND.n5916 GND.n900 240.244
R10074 GND.n5916 GND.n898 240.244
R10075 GND.n5920 GND.n898 240.244
R10076 GND.n5920 GND.n894 240.244
R10077 GND.n5926 GND.n894 240.244
R10078 GND.n5926 GND.n892 240.244
R10079 GND.n5930 GND.n892 240.244
R10080 GND.n5930 GND.n888 240.244
R10081 GND.n5936 GND.n888 240.244
R10082 GND.n5936 GND.n886 240.244
R10083 GND.n5940 GND.n886 240.244
R10084 GND.n5940 GND.n882 240.244
R10085 GND.n5946 GND.n882 240.244
R10086 GND.n5946 GND.n880 240.244
R10087 GND.n5950 GND.n880 240.244
R10088 GND.n5950 GND.n876 240.244
R10089 GND.n5956 GND.n876 240.244
R10090 GND.n5956 GND.n874 240.244
R10091 GND.n5960 GND.n874 240.244
R10092 GND.n5960 GND.n870 240.244
R10093 GND.n5966 GND.n870 240.244
R10094 GND.n5966 GND.n868 240.244
R10095 GND.n5970 GND.n868 240.244
R10096 GND.n5970 GND.n864 240.244
R10097 GND.n5976 GND.n864 240.244
R10098 GND.n5976 GND.n862 240.244
R10099 GND.n5980 GND.n862 240.244
R10100 GND.n5980 GND.n858 240.244
R10101 GND.n5986 GND.n858 240.244
R10102 GND.n5986 GND.n856 240.244
R10103 GND.n5990 GND.n856 240.244
R10104 GND.n5990 GND.n852 240.244
R10105 GND.n5996 GND.n852 240.244
R10106 GND.n5996 GND.n850 240.244
R10107 GND.n6000 GND.n850 240.244
R10108 GND.n6000 GND.n846 240.244
R10109 GND.n6006 GND.n846 240.244
R10110 GND.n6006 GND.n844 240.244
R10111 GND.n6010 GND.n844 240.244
R10112 GND.n6010 GND.n840 240.244
R10113 GND.n6016 GND.n840 240.244
R10114 GND.n6016 GND.n838 240.244
R10115 GND.n6020 GND.n838 240.244
R10116 GND.n6020 GND.n834 240.244
R10117 GND.n6026 GND.n834 240.244
R10118 GND.n6026 GND.n832 240.244
R10119 GND.n6030 GND.n832 240.244
R10120 GND.n6030 GND.n828 240.244
R10121 GND.n6036 GND.n828 240.244
R10122 GND.n6036 GND.n826 240.244
R10123 GND.n6040 GND.n826 240.244
R10124 GND.n6040 GND.n822 240.244
R10125 GND.n6046 GND.n822 240.244
R10126 GND.n6046 GND.n820 240.244
R10127 GND.n6050 GND.n820 240.244
R10128 GND.n6050 GND.n816 240.244
R10129 GND.n6056 GND.n816 240.244
R10130 GND.n6056 GND.n814 240.244
R10131 GND.n6060 GND.n814 240.244
R10132 GND.n6060 GND.n810 240.244
R10133 GND.n6066 GND.n810 240.244
R10134 GND.n6066 GND.n808 240.244
R10135 GND.n6070 GND.n808 240.244
R10136 GND.n6070 GND.n804 240.244
R10137 GND.n6076 GND.n804 240.244
R10138 GND.n6076 GND.n802 240.244
R10139 GND.n6080 GND.n802 240.244
R10140 GND.n6080 GND.n798 240.244
R10141 GND.n6086 GND.n798 240.244
R10142 GND.n6086 GND.n796 240.244
R10143 GND.n6090 GND.n796 240.244
R10144 GND.n6090 GND.n792 240.244
R10145 GND.n6096 GND.n792 240.244
R10146 GND.n6096 GND.n790 240.244
R10147 GND.n6100 GND.n790 240.244
R10148 GND.n6100 GND.n786 240.244
R10149 GND.n6106 GND.n786 240.244
R10150 GND.n6106 GND.n784 240.244
R10151 GND.n6110 GND.n784 240.244
R10152 GND.n6110 GND.n780 240.244
R10153 GND.n6116 GND.n780 240.244
R10154 GND.n6116 GND.n778 240.244
R10155 GND.n6120 GND.n778 240.244
R10156 GND.n6120 GND.n774 240.244
R10157 GND.n6126 GND.n774 240.244
R10158 GND.n6126 GND.n772 240.244
R10159 GND.n6130 GND.n772 240.244
R10160 GND.n6130 GND.n768 240.244
R10161 GND.n6136 GND.n768 240.244
R10162 GND.n6136 GND.n766 240.244
R10163 GND.n6140 GND.n766 240.244
R10164 GND.n6140 GND.n762 240.244
R10165 GND.n6146 GND.n762 240.244
R10166 GND.n6146 GND.n760 240.244
R10167 GND.n6150 GND.n760 240.244
R10168 GND.n6150 GND.n756 240.244
R10169 GND.n6156 GND.n756 240.244
R10170 GND.n6156 GND.n754 240.244
R10171 GND.n6160 GND.n754 240.244
R10172 GND.n6160 GND.n750 240.244
R10173 GND.n6166 GND.n750 240.244
R10174 GND.n6166 GND.n748 240.244
R10175 GND.n6170 GND.n748 240.244
R10176 GND.n6170 GND.n744 240.244
R10177 GND.n6176 GND.n744 240.244
R10178 GND.n6176 GND.n742 240.244
R10179 GND.n6180 GND.n742 240.244
R10180 GND.n6180 GND.n738 240.244
R10181 GND.n6186 GND.n738 240.244
R10182 GND.n6190 GND.n736 240.244
R10183 GND.n6190 GND.n732 240.244
R10184 GND.n6196 GND.n732 240.244
R10185 GND.n6196 GND.n730 240.244
R10186 GND.n6200 GND.n730 240.244
R10187 GND.n6200 GND.n726 240.244
R10188 GND.n6206 GND.n726 240.244
R10189 GND.n6206 GND.n724 240.244
R10190 GND.n6210 GND.n724 240.244
R10191 GND.n6210 GND.n720 240.244
R10192 GND.n6216 GND.n720 240.244
R10193 GND.n6216 GND.n718 240.244
R10194 GND.n6220 GND.n718 240.244
R10195 GND.n6220 GND.n714 240.244
R10196 GND.n6226 GND.n714 240.244
R10197 GND.n6226 GND.n712 240.244
R10198 GND.n6230 GND.n712 240.244
R10199 GND.n6230 GND.n708 240.244
R10200 GND.n6236 GND.n708 240.244
R10201 GND.n6236 GND.n706 240.244
R10202 GND.n6240 GND.n706 240.244
R10203 GND.n6240 GND.n702 240.244
R10204 GND.n6246 GND.n702 240.244
R10205 GND.n6246 GND.n700 240.244
R10206 GND.n6250 GND.n700 240.244
R10207 GND.n6250 GND.n696 240.244
R10208 GND.n6256 GND.n696 240.244
R10209 GND.n6256 GND.n694 240.244
R10210 GND.n6260 GND.n694 240.244
R10211 GND.n6260 GND.n690 240.244
R10212 GND.n6266 GND.n690 240.244
R10213 GND.n6266 GND.n688 240.244
R10214 GND.n6270 GND.n688 240.244
R10215 GND.n6270 GND.n684 240.244
R10216 GND.n6276 GND.n684 240.244
R10217 GND.n6276 GND.n682 240.244
R10218 GND.n6280 GND.n682 240.244
R10219 GND.n6280 GND.n678 240.244
R10220 GND.n6286 GND.n678 240.244
R10221 GND.n6286 GND.n676 240.244
R10222 GND.n6290 GND.n676 240.244
R10223 GND.n6290 GND.n672 240.244
R10224 GND.n6296 GND.n672 240.244
R10225 GND.n6296 GND.n670 240.244
R10226 GND.n6300 GND.n670 240.244
R10227 GND.n6300 GND.n666 240.244
R10228 GND.n6308 GND.n666 240.244
R10229 GND.n6308 GND.n664 240.244
R10230 GND.n1238 GND.n1235 240.244
R10231 GND.n5413 GND.n1238 240.244
R10232 GND.n5413 GND.n1241 240.244
R10233 GND.n5409 GND.n1241 240.244
R10234 GND.n5409 GND.n1244 240.244
R10235 GND.n5405 GND.n1244 240.244
R10236 GND.n5405 GND.n1250 240.244
R10237 GND.n5401 GND.n1250 240.244
R10238 GND.n5401 GND.n1252 240.244
R10239 GND.n5397 GND.n1252 240.244
R10240 GND.n5397 GND.n1258 240.244
R10241 GND.n5393 GND.n1258 240.244
R10242 GND.n5393 GND.n1260 240.244
R10243 GND.n5389 GND.n1260 240.244
R10244 GND.n5389 GND.n1266 240.244
R10245 GND.n5385 GND.n1266 240.244
R10246 GND.n5385 GND.n1268 240.244
R10247 GND.n5381 GND.n1268 240.244
R10248 GND.n5381 GND.n1274 240.244
R10249 GND.n1981 GND.n1274 240.244
R10250 GND.n1982 GND.n1981 240.244
R10251 GND.n1982 GND.n1975 240.244
R10252 GND.n2001 GND.n1975 240.244
R10253 GND.n2001 GND.n1976 240.244
R10254 GND.n1997 GND.n1976 240.244
R10255 GND.n1997 GND.n1996 240.244
R10256 GND.n1996 GND.n1995 240.244
R10257 GND.n1995 GND.n1726 240.244
R10258 GND.n2048 GND.n1726 240.244
R10259 GND.n2049 GND.n2048 240.244
R10260 GND.n2049 GND.n1721 240.244
R10261 GND.n2075 GND.n1721 240.244
R10262 GND.n2075 GND.n1722 240.244
R10263 GND.n2071 GND.n1722 240.244
R10264 GND.n2071 GND.n2070 240.244
R10265 GND.n2070 GND.n2069 240.244
R10266 GND.n2069 GND.n2057 240.244
R10267 GND.n2065 GND.n2057 240.244
R10268 GND.n2065 GND.n2064 240.244
R10269 GND.n2064 GND.n1653 240.244
R10270 GND.n2206 GND.n1653 240.244
R10271 GND.n2206 GND.n1654 240.244
R10272 GND.n2201 GND.n1654 240.244
R10273 GND.n2201 GND.n1657 240.244
R10274 GND.n2137 GND.n1657 240.244
R10275 GND.n2189 GND.n2137 240.244
R10276 GND.n2189 GND.n2142 240.244
R10277 GND.n2184 GND.n2142 240.244
R10278 GND.n2184 GND.n2183 240.244
R10279 GND.n2183 GND.n2146 240.244
R10280 GND.n2179 GND.n2146 240.244
R10281 GND.n2179 GND.n2178 240.244
R10282 GND.n2178 GND.n2177 240.244
R10283 GND.n2177 GND.n2150 240.244
R10284 GND.n2173 GND.n2150 240.244
R10285 GND.n2173 GND.n2172 240.244
R10286 GND.n2172 GND.n2171 240.244
R10287 GND.n2171 GND.n2156 240.244
R10288 GND.n2167 GND.n2156 240.244
R10289 GND.n2167 GND.n2166 240.244
R10290 GND.n2166 GND.n2165 240.244
R10291 GND.n2165 GND.n1560 240.244
R10292 GND.n2307 GND.n1560 240.244
R10293 GND.n2307 GND.n1555 240.244
R10294 GND.n2328 GND.n1555 240.244
R10295 GND.n2328 GND.n1556 240.244
R10296 GND.n2324 GND.n1556 240.244
R10297 GND.n2324 GND.n2323 240.244
R10298 GND.n2323 GND.n2322 240.244
R10299 GND.n2322 GND.n2315 240.244
R10300 GND.n2315 GND.n1525 240.244
R10301 GND.n5167 GND.n1525 240.244
R10302 GND.n5167 GND.n1526 240.244
R10303 GND.n5163 GND.n1526 240.244
R10304 GND.n5163 GND.n5161 240.244
R10305 GND.n5161 GND.n1532 240.244
R10306 GND.n3517 GND.n1532 240.244
R10307 GND.n3517 GND.n3512 240.244
R10308 GND.n3523 GND.n3512 240.244
R10309 GND.n3523 GND.n3466 240.244
R10310 GND.n3535 GND.n3466 240.244
R10311 GND.n3535 GND.n3462 240.244
R10312 GND.n3541 GND.n3462 240.244
R10313 GND.n3541 GND.n3455 240.244
R10314 GND.n3552 GND.n3455 240.244
R10315 GND.n3552 GND.n3451 240.244
R10316 GND.n3558 GND.n3451 240.244
R10317 GND.n3558 GND.n3443 240.244
R10318 GND.n3569 GND.n3443 240.244
R10319 GND.n3569 GND.n3439 240.244
R10320 GND.n3575 GND.n3439 240.244
R10321 GND.n3575 GND.n3431 240.244
R10322 GND.n3586 GND.n3431 240.244
R10323 GND.n3586 GND.n3427 240.244
R10324 GND.n3592 GND.n3427 240.244
R10325 GND.n3592 GND.n3418 240.244
R10326 GND.n3604 GND.n3418 240.244
R10327 GND.n3604 GND.n3414 240.244
R10328 GND.n3610 GND.n3414 240.244
R10329 GND.n3610 GND.n3385 240.244
R10330 GND.n3740 GND.n3385 240.244
R10331 GND.n3740 GND.n3380 240.244
R10332 GND.n3754 GND.n3380 240.244
R10333 GND.n3754 GND.n3381 240.244
R10334 GND.n3750 GND.n3381 240.244
R10335 GND.n3750 GND.n3749 240.244
R10336 GND.n3749 GND.n3347 240.244
R10337 GND.n3786 GND.n3347 240.244
R10338 GND.n3786 GND.n3342 240.244
R10339 GND.n3794 GND.n3342 240.244
R10340 GND.n3794 GND.n3343 240.244
R10341 GND.n3343 GND.n3318 240.244
R10342 GND.n3840 GND.n3318 240.244
R10343 GND.n3840 GND.n3312 240.244
R10344 GND.n3848 GND.n3312 240.244
R10345 GND.n3848 GND.n3314 240.244
R10346 GND.n3314 GND.n3294 240.244
R10347 GND.n3901 GND.n3294 240.244
R10348 GND.n3901 GND.n3289 240.244
R10349 GND.n3915 GND.n3289 240.244
R10350 GND.n3915 GND.n3290 240.244
R10351 GND.n3911 GND.n3290 240.244
R10352 GND.n3911 GND.n3910 240.244
R10353 GND.n3910 GND.n3259 240.244
R10354 GND.n3947 GND.n3259 240.244
R10355 GND.n3947 GND.n3254 240.244
R10356 GND.n3955 GND.n3254 240.244
R10357 GND.n3955 GND.n3255 240.244
R10358 GND.n3255 GND.n3231 240.244
R10359 GND.n4000 GND.n3231 240.244
R10360 GND.n4000 GND.n3224 240.244
R10361 GND.n4008 GND.n3224 240.244
R10362 GND.n4008 GND.n3227 240.244
R10363 GND.n3227 GND.n3206 240.244
R10364 GND.n4061 GND.n3206 240.244
R10365 GND.n4061 GND.n3201 240.244
R10366 GND.n4075 GND.n3201 240.244
R10367 GND.n4075 GND.n3202 240.244
R10368 GND.n4071 GND.n3202 240.244
R10369 GND.n4071 GND.n4070 240.244
R10370 GND.n4070 GND.n3173 240.244
R10371 GND.n4107 GND.n3173 240.244
R10372 GND.n4107 GND.n3168 240.244
R10373 GND.n4115 GND.n3168 240.244
R10374 GND.n4115 GND.n3169 240.244
R10375 GND.n3169 GND.n3144 240.244
R10376 GND.n4160 GND.n3144 240.244
R10377 GND.n4160 GND.n3138 240.244
R10378 GND.n4168 GND.n3138 240.244
R10379 GND.n4168 GND.n3140 240.244
R10380 GND.n3140 GND.n3119 240.244
R10381 GND.n4208 GND.n3119 240.244
R10382 GND.n4208 GND.n3114 240.244
R10383 GND.n4225 GND.n3114 240.244
R10384 GND.n4225 GND.n3115 240.244
R10385 GND.n4221 GND.n3115 240.244
R10386 GND.n4221 GND.n4220 240.244
R10387 GND.n4220 GND.n4219 240.244
R10388 GND.n4219 GND.n3078 240.244
R10389 GND.n4322 GND.n3078 240.244
R10390 GND.n4322 GND.n3072 240.244
R10391 GND.n4330 GND.n3072 240.244
R10392 GND.n4330 GND.n3074 240.244
R10393 GND.n3074 GND.n3028 240.244
R10394 GND.n4391 GND.n3028 240.244
R10395 GND.n4391 GND.n3024 240.244
R10396 GND.n4397 GND.n3024 240.244
R10397 GND.n4397 GND.n3016 240.244
R10398 GND.n4408 GND.n3016 240.244
R10399 GND.n4408 GND.n3012 240.244
R10400 GND.n4414 GND.n3012 240.244
R10401 GND.n4414 GND.n3004 240.244
R10402 GND.n4425 GND.n3004 240.244
R10403 GND.n4425 GND.n3000 240.244
R10404 GND.n4431 GND.n3000 240.244
R10405 GND.n4431 GND.n2992 240.244
R10406 GND.n4442 GND.n2992 240.244
R10407 GND.n4442 GND.n2988 240.244
R10408 GND.n4448 GND.n2988 240.244
R10409 GND.n4448 GND.n2980 240.244
R10410 GND.n4459 GND.n2980 240.244
R10411 GND.n4459 GND.n2976 240.244
R10412 GND.n4465 GND.n2976 240.244
R10413 GND.n4465 GND.n2968 240.244
R10414 GND.n4476 GND.n2968 240.244
R10415 GND.n4476 GND.n2964 240.244
R10416 GND.n4485 GND.n2964 240.244
R10417 GND.n4485 GND.n2956 240.244
R10418 GND.n4496 GND.n2956 240.244
R10419 GND.n4497 GND.n4496 240.244
R10420 GND.n4497 GND.n2495 240.244
R10421 GND.n2951 GND.n2495 240.244
R10422 GND.n4513 GND.n2951 240.244
R10423 GND.n4513 GND.n2952 240.244
R10424 GND.n4509 GND.n2952 240.244
R10425 GND.n4509 GND.n4508 240.244
R10426 GND.n4508 GND.n2615 240.244
R10427 GND.n4862 GND.n2615 240.244
R10428 GND.n4862 GND.n2616 240.244
R10429 GND.n4858 GND.n2616 240.244
R10430 GND.n4858 GND.n2622 240.244
R10431 GND.n2763 GND.n2622 240.244
R10432 GND.n2769 GND.n2763 240.244
R10433 GND.n2770 GND.n2769 240.244
R10434 GND.n2771 GND.n2770 240.244
R10435 GND.n2771 GND.n2759 240.244
R10436 GND.n2777 GND.n2759 240.244
R10437 GND.n2778 GND.n2777 240.244
R10438 GND.n2779 GND.n2778 240.244
R10439 GND.n2779 GND.n2755 240.244
R10440 GND.n2785 GND.n2755 240.244
R10441 GND.n2786 GND.n2785 240.244
R10442 GND.n2787 GND.n2786 240.244
R10443 GND.n2787 GND.n2751 240.244
R10444 GND.n2794 GND.n2751 240.244
R10445 GND.n2795 GND.n2794 240.244
R10446 GND.n2796 GND.n2795 240.244
R10447 GND.n2796 GND.n2748 240.244
R10448 GND.n2800 GND.n2748 240.244
R10449 GND.n2801 GND.n2800 240.244
R10450 GND.n2801 GND.n2745 240.244
R10451 GND.n4791 GND.n2745 240.244
R10452 GND.n4791 GND.n2746 240.244
R10453 GND.n4786 GND.n2746 240.244
R10454 GND.n4786 GND.n4785 240.244
R10455 GND.n4785 GND.n2871 240.244
R10456 GND.n2871 GND.n2806 240.244
R10457 GND.n2866 GND.n2806 240.244
R10458 GND.n2866 GND.n2865 240.244
R10459 GND.n2865 GND.n2864 240.244
R10460 GND.n2864 GND.n2809 240.244
R10461 GND.n2860 GND.n2809 240.244
R10462 GND.n2860 GND.n2859 240.244
R10463 GND.n2859 GND.n2858 240.244
R10464 GND.n2858 GND.n2815 240.244
R10465 GND.n2854 GND.n2815 240.244
R10466 GND.n2854 GND.n2853 240.244
R10467 GND.n2853 GND.n2852 240.244
R10468 GND.n2852 GND.n2821 240.244
R10469 GND.n2848 GND.n2821 240.244
R10470 GND.n2848 GND.n2847 240.244
R10471 GND.n2847 GND.n2846 240.244
R10472 GND.n2846 GND.n2827 240.244
R10473 GND.n2842 GND.n2827 240.244
R10474 GND.n2842 GND.n2841 240.244
R10475 GND.n2841 GND.n2840 240.244
R10476 GND.n2840 GND.n2833 240.244
R10477 GND.n2833 GND.n453 240.244
R10478 GND.n6348 GND.n453 240.244
R10479 GND.n6348 GND.n454 240.244
R10480 GND.n6344 GND.n454 240.244
R10481 GND.n6344 GND.n460 240.244
R10482 GND.n6340 GND.n460 240.244
R10483 GND.n6340 GND.n635 240.244
R10484 GND.n6336 GND.n635 240.244
R10485 GND.n6336 GND.n641 240.244
R10486 GND.n6332 GND.n641 240.244
R10487 GND.n6332 GND.n643 240.244
R10488 GND.n6328 GND.n643 240.244
R10489 GND.n6328 GND.n649 240.244
R10490 GND.n6324 GND.n649 240.244
R10491 GND.n6324 GND.n651 240.244
R10492 GND.n6320 GND.n651 240.244
R10493 GND.n6320 GND.n657 240.244
R10494 GND.n6316 GND.n657 240.244
R10495 GND.n6316 GND.n659 240.244
R10496 GND.n6312 GND.n659 240.244
R10497 GND.n5516 GND.n1140 240.244
R10498 GND.n5512 GND.n1140 240.244
R10499 GND.n5512 GND.n1145 240.244
R10500 GND.n5508 GND.n1145 240.244
R10501 GND.n5508 GND.n1147 240.244
R10502 GND.n5504 GND.n1147 240.244
R10503 GND.n5504 GND.n1153 240.244
R10504 GND.n5500 GND.n1153 240.244
R10505 GND.n5500 GND.n1155 240.244
R10506 GND.n5496 GND.n1155 240.244
R10507 GND.n5496 GND.n1161 240.244
R10508 GND.n5492 GND.n1161 240.244
R10509 GND.n5492 GND.n1163 240.244
R10510 GND.n5488 GND.n1163 240.244
R10511 GND.n5488 GND.n1169 240.244
R10512 GND.n5484 GND.n1169 240.244
R10513 GND.n5484 GND.n1171 240.244
R10514 GND.n5480 GND.n1171 240.244
R10515 GND.n5480 GND.n1177 240.244
R10516 GND.n5476 GND.n1177 240.244
R10517 GND.n5476 GND.n1179 240.244
R10518 GND.n5472 GND.n1179 240.244
R10519 GND.n5472 GND.n1185 240.244
R10520 GND.n5468 GND.n1185 240.244
R10521 GND.n5468 GND.n1187 240.244
R10522 GND.n5464 GND.n1187 240.244
R10523 GND.n5464 GND.n1193 240.244
R10524 GND.n5460 GND.n1193 240.244
R10525 GND.n5460 GND.n1195 240.244
R10526 GND.n5456 GND.n1195 240.244
R10527 GND.n5456 GND.n1201 240.244
R10528 GND.n5452 GND.n1201 240.244
R10529 GND.n5452 GND.n1203 240.244
R10530 GND.n5448 GND.n1203 240.244
R10531 GND.n5448 GND.n1209 240.244
R10532 GND.n5444 GND.n1209 240.244
R10533 GND.n5444 GND.n1211 240.244
R10534 GND.n5440 GND.n1211 240.244
R10535 GND.n5440 GND.n1217 240.244
R10536 GND.n5436 GND.n1217 240.244
R10537 GND.n5436 GND.n1219 240.244
R10538 GND.n5432 GND.n1219 240.244
R10539 GND.n5432 GND.n1225 240.244
R10540 GND.n5428 GND.n1225 240.244
R10541 GND.n5428 GND.n1227 240.244
R10542 GND.n5424 GND.n1227 240.244
R10543 GND.n5424 GND.n1233 240.244
R10544 GND.n5420 GND.n1233 240.244
R10545 GND.n3509 GND.n1533 240.244
R10546 GND.n3510 GND.n3509 240.244
R10547 GND.n3525 GND.n3510 240.244
R10548 GND.n3525 GND.n3468 240.244
R10549 GND.n3531 GND.n3468 240.244
R10550 GND.n3531 GND.n3461 240.244
R10551 GND.n3543 GND.n3461 240.244
R10552 GND.n3543 GND.n3457 240.244
R10553 GND.n3549 GND.n3457 240.244
R10554 GND.n3549 GND.n3449 240.244
R10555 GND.n3560 GND.n3449 240.244
R10556 GND.n3560 GND.n3445 240.244
R10557 GND.n3566 GND.n3445 240.244
R10558 GND.n3566 GND.n3437 240.244
R10559 GND.n3577 GND.n3437 240.244
R10560 GND.n3577 GND.n3433 240.244
R10561 GND.n3583 GND.n3433 240.244
R10562 GND.n3583 GND.n3425 240.244
R10563 GND.n3594 GND.n3425 240.244
R10564 GND.n3594 GND.n3420 240.244
R10565 GND.n3601 GND.n3420 240.244
R10566 GND.n3601 GND.n3412 240.244
R10567 GND.n3612 GND.n3412 240.244
R10568 GND.n3613 GND.n3612 240.244
R10569 GND.n3613 GND.n3387 240.244
R10570 GND.n3647 GND.n3387 240.244
R10571 GND.n3647 GND.n3379 240.244
R10572 GND.n3618 GND.n3379 240.244
R10573 GND.n3619 GND.n3618 240.244
R10574 GND.n3620 GND.n3619 240.244
R10575 GND.n3621 GND.n3620 240.244
R10576 GND.n3621 GND.n3350 240.244
R10577 GND.n3624 GND.n3350 240.244
R10578 GND.n3624 GND.n3341 240.244
R10579 GND.n3627 GND.n3341 240.244
R10580 GND.n3628 GND.n3627 240.244
R10581 GND.n3628 GND.n3320 240.244
R10582 GND.n3320 GND.n3309 240.244
R10583 GND.n3850 GND.n3309 240.244
R10584 GND.n3850 GND.n3304 240.244
R10585 GND.n3890 GND.n3304 240.244
R10586 GND.n3890 GND.n3296 240.244
R10587 GND.n3855 GND.n3296 240.244
R10588 GND.n3855 GND.n3288 240.244
R10589 GND.n3856 GND.n3288 240.244
R10590 GND.n3859 GND.n3856 240.244
R10591 GND.n3860 GND.n3859 240.244
R10592 GND.n3861 GND.n3860 240.244
R10593 GND.n3861 GND.n3262 240.244
R10594 GND.n3863 GND.n3262 240.244
R10595 GND.n3863 GND.n3253 240.244
R10596 GND.n3866 GND.n3253 240.244
R10597 GND.n3867 GND.n3866 240.244
R10598 GND.n3867 GND.n3233 240.244
R10599 GND.n3233 GND.n3221 240.244
R10600 GND.n4010 GND.n3221 240.244
R10601 GND.n4010 GND.n3216 240.244
R10602 GND.n4051 GND.n3216 240.244
R10603 GND.n4051 GND.n3208 240.244
R10604 GND.n4015 GND.n3208 240.244
R10605 GND.n4015 GND.n3199 240.244
R10606 GND.n4016 GND.n3199 240.244
R10607 GND.n4019 GND.n4016 240.244
R10608 GND.n4020 GND.n4019 240.244
R10609 GND.n4023 GND.n4020 240.244
R10610 GND.n4023 GND.n3176 240.244
R10611 GND.n4024 GND.n3176 240.244
R10612 GND.n4024 GND.n3167 240.244
R10613 GND.n4027 GND.n3167 240.244
R10614 GND.n4028 GND.n4027 240.244
R10615 GND.n4028 GND.n3146 240.244
R10616 GND.n3146 GND.n3134 240.244
R10617 GND.n4170 GND.n3134 240.244
R10618 GND.n4170 GND.n3129 240.244
R10619 GND.n4198 GND.n3129 240.244
R10620 GND.n4198 GND.n3121 240.244
R10621 GND.n4175 GND.n3121 240.244
R10622 GND.n4175 GND.n3113 240.244
R10623 GND.n4176 GND.n3113 240.244
R10624 GND.n4179 GND.n4176 240.244
R10625 GND.n4180 GND.n4179 240.244
R10626 GND.n4181 GND.n4180 240.244
R10627 GND.n4181 GND.n3089 240.244
R10628 GND.n3089 GND.n3080 240.244
R10629 GND.n3080 GND.n3069 240.244
R10630 GND.n4332 GND.n3069 240.244
R10631 GND.n4332 GND.n3064 240.244
R10632 GND.n4339 GND.n3064 240.244
R10633 GND.n4339 GND.n3030 240.244
R10634 GND.n3030 GND.n3022 240.244
R10635 GND.n4399 GND.n3022 240.244
R10636 GND.n4399 GND.n3018 240.244
R10637 GND.n4405 GND.n3018 240.244
R10638 GND.n4405 GND.n3010 240.244
R10639 GND.n4416 GND.n3010 240.244
R10640 GND.n4416 GND.n3006 240.244
R10641 GND.n4422 GND.n3006 240.244
R10642 GND.n4422 GND.n2998 240.244
R10643 GND.n4433 GND.n2998 240.244
R10644 GND.n4433 GND.n2994 240.244
R10645 GND.n4439 GND.n2994 240.244
R10646 GND.n4439 GND.n2986 240.244
R10647 GND.n4450 GND.n2986 240.244
R10648 GND.n4450 GND.n2982 240.244
R10649 GND.n4456 GND.n2982 240.244
R10650 GND.n4456 GND.n2973 240.244
R10651 GND.n4467 GND.n2973 240.244
R10652 GND.n4467 GND.n2969 240.244
R10653 GND.n4473 GND.n2969 240.244
R10654 GND.n4473 GND.n2962 240.244
R10655 GND.n4487 GND.n2962 240.244
R10656 GND.n4487 GND.n2958 240.244
R10657 GND.n4493 GND.n2958 240.244
R10658 GND.n4493 GND.n2497 240.244
R10659 GND.n4981 GND.n2497 240.244
R10660 GND.n2503 GND.n2502 240.244
R10661 GND.n2919 GND.n2506 240.244
R10662 GND.n2508 GND.n2507 240.244
R10663 GND.n2922 GND.n2511 240.244
R10664 GND.n2513 GND.n2512 240.244
R10665 GND.n2934 GND.n2933 240.244
R10666 GND.n2947 GND.n2927 240.244
R10667 GND.n4518 GND.n2917 240.244
R10668 GND.n4516 GND.n2904 240.244
R10669 GND.n5158 GND.n1536 240.244
R10670 GND.n2352 GND.n1536 240.244
R10671 GND.n2353 GND.n2352 240.244
R10672 GND.n2354 GND.n2353 240.244
R10673 GND.n3533 GND.n2354 240.244
R10674 GND.n3533 GND.n2357 240.244
R10675 GND.n2358 GND.n2357 240.244
R10676 GND.n2359 GND.n2358 240.244
R10677 GND.n3550 GND.n2359 240.244
R10678 GND.n3550 GND.n2362 240.244
R10679 GND.n2363 GND.n2362 240.244
R10680 GND.n2364 GND.n2363 240.244
R10681 GND.n3567 GND.n2364 240.244
R10682 GND.n3567 GND.n2367 240.244
R10683 GND.n2368 GND.n2367 240.244
R10684 GND.n2369 GND.n2368 240.244
R10685 GND.n3584 GND.n2369 240.244
R10686 GND.n3584 GND.n2372 240.244
R10687 GND.n2373 GND.n2372 240.244
R10688 GND.n2374 GND.n2373 240.244
R10689 GND.n3602 GND.n2374 240.244
R10690 GND.n3602 GND.n2377 240.244
R10691 GND.n2378 GND.n2377 240.244
R10692 GND.n2379 GND.n2378 240.244
R10693 GND.n3738 GND.n2379 240.244
R10694 GND.n3738 GND.n2382 240.244
R10695 GND.n2383 GND.n2382 240.244
R10696 GND.n2384 GND.n2383 240.244
R10697 GND.n3362 GND.n2384 240.244
R10698 GND.n3362 GND.n2387 240.244
R10699 GND.n2388 GND.n2387 240.244
R10700 GND.n2389 GND.n2388 240.244
R10701 GND.n3338 GND.n2389 240.244
R10702 GND.n3338 GND.n2392 240.244
R10703 GND.n2393 GND.n2392 240.244
R10704 GND.n2394 GND.n2393 240.244
R10705 GND.n3838 GND.n2394 240.244
R10706 GND.n3838 GND.n2397 240.244
R10707 GND.n2398 GND.n2397 240.244
R10708 GND.n2399 GND.n2398 240.244
R10709 GND.n3891 GND.n2399 240.244
R10710 GND.n3891 GND.n2402 240.244
R10711 GND.n2403 GND.n2402 240.244
R10712 GND.n2404 GND.n2403 240.244
R10713 GND.n3281 GND.n2404 240.244
R10714 GND.n3281 GND.n2407 240.244
R10715 GND.n2408 GND.n2407 240.244
R10716 GND.n2409 GND.n2408 240.244
R10717 GND.n3264 GND.n2409 240.244
R10718 GND.n3264 GND.n2412 240.244
R10719 GND.n2413 GND.n2412 240.244
R10720 GND.n2414 GND.n2413 240.244
R10721 GND.n3240 GND.n2414 240.244
R10722 GND.n3240 GND.n2417 240.244
R10723 GND.n2418 GND.n2417 240.244
R10724 GND.n2419 GND.n2418 240.244
R10725 GND.n3225 GND.n2419 240.244
R10726 GND.n3225 GND.n2422 240.244
R10727 GND.n2423 GND.n2422 240.244
R10728 GND.n2424 GND.n2423 240.244
R10729 GND.n3200 GND.n2424 240.244
R10730 GND.n3200 GND.n2427 240.244
R10731 GND.n2428 GND.n2427 240.244
R10732 GND.n2429 GND.n2428 240.244
R10733 GND.n4021 GND.n2429 240.244
R10734 GND.n4021 GND.n2432 240.244
R10735 GND.n2433 GND.n2432 240.244
R10736 GND.n2434 GND.n2433 240.244
R10737 GND.n3160 GND.n2434 240.244
R10738 GND.n3160 GND.n2437 240.244
R10739 GND.n2438 GND.n2437 240.244
R10740 GND.n2439 GND.n2438 240.244
R10741 GND.n3137 GND.n2439 240.244
R10742 GND.n3137 GND.n2442 240.244
R10743 GND.n2443 GND.n2442 240.244
R10744 GND.n2444 GND.n2443 240.244
R10745 GND.n3110 GND.n2444 240.244
R10746 GND.n3110 GND.n2447 240.244
R10747 GND.n2448 GND.n2447 240.244
R10748 GND.n2449 GND.n2448 240.244
R10749 GND.n3094 GND.n2449 240.244
R10750 GND.n3094 GND.n2452 240.244
R10751 GND.n2453 GND.n2452 240.244
R10752 GND.n2454 GND.n2453 240.244
R10753 GND.n3082 GND.n2454 240.244
R10754 GND.n3082 GND.n2457 240.244
R10755 GND.n2458 GND.n2457 240.244
R10756 GND.n2459 GND.n2458 240.244
R10757 GND.n4389 GND.n2459 240.244
R10758 GND.n4389 GND.n2462 240.244
R10759 GND.n2463 GND.n2462 240.244
R10760 GND.n2464 GND.n2463 240.244
R10761 GND.n4406 GND.n2464 240.244
R10762 GND.n4406 GND.n2467 240.244
R10763 GND.n2468 GND.n2467 240.244
R10764 GND.n2469 GND.n2468 240.244
R10765 GND.n4423 GND.n2469 240.244
R10766 GND.n4423 GND.n2472 240.244
R10767 GND.n2473 GND.n2472 240.244
R10768 GND.n2474 GND.n2473 240.244
R10769 GND.n4440 GND.n2474 240.244
R10770 GND.n4440 GND.n2477 240.244
R10771 GND.n2478 GND.n2477 240.244
R10772 GND.n2479 GND.n2478 240.244
R10773 GND.n4457 GND.n2479 240.244
R10774 GND.n4457 GND.n2482 240.244
R10775 GND.n2483 GND.n2482 240.244
R10776 GND.n2484 GND.n2483 240.244
R10777 GND.n4474 GND.n2484 240.244
R10778 GND.n4474 GND.n2487 240.244
R10779 GND.n2488 GND.n2487 240.244
R10780 GND.n2489 GND.n2488 240.244
R10781 GND.n4494 GND.n2489 240.244
R10782 GND.n4494 GND.n2492 240.244
R10783 GND.n4983 GND.n2492 240.244
R10784 GND.n3477 GND.n3476 240.244
R10785 GND.n3480 GND.n3477 240.244
R10786 GND.n3483 GND.n3482 240.244
R10787 GND.n3489 GND.n3485 240.244
R10788 GND.n3491 GND.n3488 240.244
R10789 GND.n1474 GND.n1473 240.244
R10790 GND.n1492 GND.n1482 240.244
R10791 GND.n1491 GND.n1483 240.244
R10792 GND.n5201 GND.n1491 240.244
R10793 GND.n5199 GND.n5198 240.244
R10794 GND.n2915 GND.t80 229.109
R10795 GND.n5202 GND.t87 229.109
R10796 GND.n3372 GND.n3371 228.118
R10797 GND.n3056 GND.n3055 228.118
R10798 GND.n1412 GND.t103 225.582
R10799 GND.n1426 GND.t124 225.582
R10800 GND.n1439 GND.t133 225.582
R10801 GND.n1453 GND.t76 225.582
R10802 GND.n1466 GND.t127 225.582
R10803 GND.n2908 GND.t94 225.582
R10804 GND.n1501 GND.t106 225.582
R10805 GND.n1759 GND.t130 225.582
R10806 GND.n2559 GND.t66 225.582
R10807 GND.n2571 GND.t84 225.582
R10808 GND.n2583 GND.t58 225.582
R10809 GND.n2595 GND.t136 225.582
R10810 GND.n2605 GND.t115 225.582
R10811 GND.n485 GND.t118 225.582
R10812 GND.n493 GND.t109 225.582
R10813 GND.n500 GND.t55 225.582
R10814 GND.n508 GND.t51 225.582
R10815 GND.n516 GND.t145 225.582
R10816 GND.n4677 GND.t100 225.582
R10817 GND.n1837 GND.t97 225.582
R10818 GND.n1802 GND.t112 225.582
R10819 GND.n1792 GND.t142 225.582
R10820 GND.n1909 GND.t62 225.582
R10821 GND.n1769 GND.t148 225.582
R10822 GND.n3651 GND.t154 223.94
R10823 GND.n3653 GND.t72 223.94
R10824 GND.n4252 GND.t47 223.94
R10825 GND.n4346 GND.t139 223.94
R10826 GND.n2577 GND.n2529 199.319
R10827 GND.n2577 GND.n2530 199.319
R10828 GND.n5177 GND.n5176 199.319
R10829 GND.n1412 GND.t104 195.232
R10830 GND.n1426 GND.t125 195.232
R10831 GND.n1439 GND.t134 195.232
R10832 GND.n1453 GND.t78 195.232
R10833 GND.n1466 GND.t128 195.232
R10834 GND.n2908 GND.t96 195.232
R10835 GND.n1501 GND.t107 195.232
R10836 GND.n1759 GND.t132 195.232
R10837 GND.n2559 GND.t68 195.232
R10838 GND.n2571 GND.t86 195.232
R10839 GND.n2583 GND.t61 195.232
R10840 GND.n2595 GND.t138 195.232
R10841 GND.n2605 GND.t117 195.232
R10842 GND.n485 GND.t119 195.232
R10843 GND.n493 GND.t110 195.232
R10844 GND.n500 GND.t56 195.232
R10845 GND.n508 GND.t53 195.232
R10846 GND.n516 GND.t146 195.232
R10847 GND.n4677 GND.t101 195.232
R10848 GND.n1837 GND.t99 195.232
R10849 GND.n1802 GND.t114 195.232
R10850 GND.n1792 GND.t144 195.232
R10851 GND.n1909 GND.t65 195.232
R10852 GND.n1769 GND.t150 195.232
R10853 GND.n3697 GND.n1432 191.936
R10854 GND.n4918 GND.n2576 191.936
R10855 GND.n136 GND.n135 185
R10856 GND.n134 GND.n133 185
R10857 GND.n149 GND.n148 185
R10858 GND.n147 GND.n146 185
R10859 GND.n110 GND.n109 185
R10860 GND.n108 GND.n107 185
R10861 GND.n123 GND.n122 185
R10862 GND.n121 GND.n120 185
R10863 GND.n84 GND.n83 185
R10864 GND.n82 GND.n81 185
R10865 GND.n97 GND.n96 185
R10866 GND.n95 GND.n94 185
R10867 GND.n58 GND.n57 185
R10868 GND.n56 GND.n55 185
R10869 GND.n71 GND.n70 185
R10870 GND.n69 GND.n68 185
R10871 GND.n32 GND.n31 185
R10872 GND.n30 GND.n29 185
R10873 GND.n45 GND.n44 185
R10874 GND.n43 GND.n42 185
R10875 GND.n7 GND.n6 185
R10876 GND.n5 GND.n4 185
R10877 GND.n20 GND.n19 185
R10878 GND.n18 GND.n17 185
R10879 GND.n305 GND.n304 185
R10880 GND.n303 GND.n302 185
R10881 GND.n292 GND.n291 185
R10882 GND.n290 GND.n289 185
R10883 GND.n279 GND.n278 185
R10884 GND.n277 GND.n276 185
R10885 GND.n266 GND.n265 185
R10886 GND.n264 GND.n263 185
R10887 GND.n253 GND.n252 185
R10888 GND.n251 GND.n250 185
R10889 GND.n240 GND.n239 185
R10890 GND.n238 GND.n237 185
R10891 GND.n227 GND.n226 185
R10892 GND.n225 GND.n224 185
R10893 GND.n214 GND.n213 185
R10894 GND.n212 GND.n211 185
R10895 GND.n201 GND.n200 185
R10896 GND.n199 GND.n198 185
R10897 GND.n188 GND.n187 185
R10898 GND.n186 GND.n185 185
R10899 GND.n176 GND.n175 185
R10900 GND.n174 GND.n173 185
R10901 GND.n163 GND.n162 185
R10902 GND.n161 GND.n160 185
R10903 GND.n4387 GND.n3054 163.367
R10904 GND.n4383 GND.n4382 163.367
R10905 GND.n4379 GND.n4378 163.367
R10906 GND.n4375 GND.n4374 163.367
R10907 GND.n4371 GND.n4370 163.367
R10908 GND.n4367 GND.n4366 163.367
R10909 GND.n4363 GND.n4362 163.367
R10910 GND.n4359 GND.n4358 163.367
R10911 GND.n4354 GND.n4353 163.367
R10912 GND.n4350 GND.n4349 163.367
R10913 GND.n4255 GND.n3031 163.367
R10914 GND.n4259 GND.n4258 163.367
R10915 GND.n4263 GND.n4262 163.367
R10916 GND.n4267 GND.n4266 163.367
R10917 GND.n4271 GND.n4270 163.367
R10918 GND.n4275 GND.n4274 163.367
R10919 GND.n4279 GND.n4278 163.367
R10920 GND.n4283 GND.n4282 163.367
R10921 GND.n4287 GND.n4286 163.367
R10922 GND.n4291 GND.n4290 163.367
R10923 GND.n3378 GND.n3366 163.367
R10924 GND.n3763 GND.n3366 163.367
R10925 GND.n3763 GND.n3364 163.367
R10926 GND.n3767 GND.n3364 163.367
R10927 GND.n3767 GND.n3355 163.367
R10928 GND.n3778 GND.n3355 163.367
R10929 GND.n3778 GND.n3352 163.367
R10930 GND.n3784 GND.n3352 163.367
R10931 GND.n3784 GND.n3353 163.367
R10932 GND.n3353 GND.n3340 163.367
R10933 GND.n3340 GND.n3331 163.367
R10934 GND.n3803 GND.n3331 163.367
R10935 GND.n3803 GND.n3328 163.367
R10936 GND.n3825 GND.n3328 163.367
R10937 GND.n3825 GND.n3329 163.367
R10938 GND.n3329 GND.n3321 163.367
R10939 GND.n3820 GND.n3321 163.367
R10940 GND.n3820 GND.n3818 163.367
R10941 GND.n3818 GND.n3817 163.367
R10942 GND.n3817 GND.n3807 163.367
R10943 GND.n3807 GND.n3303 163.367
R10944 GND.n3812 GND.n3303 163.367
R10945 GND.n3812 GND.n3297 163.367
R10946 GND.n3809 GND.n3297 163.367
R10947 GND.n3809 GND.n3287 163.367
R10948 GND.n3287 GND.n3278 163.367
R10949 GND.n3924 GND.n3278 163.367
R10950 GND.n3924 GND.n3276 163.367
R10951 GND.n3928 GND.n3276 163.367
R10952 GND.n3928 GND.n3268 163.367
R10953 GND.n3939 GND.n3268 163.367
R10954 GND.n3939 GND.n3265 163.367
R10955 GND.n3945 GND.n3265 163.367
R10956 GND.n3945 GND.n3266 163.367
R10957 GND.n3266 GND.n3252 163.367
R10958 GND.n3252 GND.n3245 163.367
R10959 GND.n3964 GND.n3245 163.367
R10960 GND.n3964 GND.n3242 163.367
R10961 GND.n3986 GND.n3242 163.367
R10962 GND.n3986 GND.n3243 163.367
R10963 GND.n3243 GND.n3234 163.367
R10964 GND.n3981 GND.n3234 163.367
R10965 GND.n3981 GND.n3979 163.367
R10966 GND.n3979 GND.n3978 163.367
R10967 GND.n3978 GND.n3968 163.367
R10968 GND.n3968 GND.n3215 163.367
R10969 GND.n3973 GND.n3215 163.367
R10970 GND.n3973 GND.n3209 163.367
R10971 GND.n3970 GND.n3209 163.367
R10972 GND.n3970 GND.n3198 163.367
R10973 GND.n3198 GND.n3190 163.367
R10974 GND.n4084 GND.n3190 163.367
R10975 GND.n4084 GND.n3188 163.367
R10976 GND.n4088 GND.n3188 163.367
R10977 GND.n4088 GND.n3181 163.367
R10978 GND.n4099 GND.n3181 163.367
R10979 GND.n4099 GND.n3178 163.367
R10980 GND.n4105 GND.n3178 163.367
R10981 GND.n4105 GND.n3179 163.367
R10982 GND.n3179 GND.n3166 163.367
R10983 GND.n3166 GND.n3157 163.367
R10984 GND.n4124 GND.n3157 163.367
R10985 GND.n4124 GND.n3154 163.367
R10986 GND.n4146 GND.n3154 163.367
R10987 GND.n4146 GND.n3155 163.367
R10988 GND.n3155 GND.n3147 163.367
R10989 GND.n4141 GND.n3147 163.367
R10990 GND.n4141 GND.n4139 163.367
R10991 GND.n4139 GND.n4138 163.367
R10992 GND.n4138 GND.n4128 163.367
R10993 GND.n4128 GND.n3128 163.367
R10994 GND.n4133 GND.n3128 163.367
R10995 GND.n4133 GND.n3122 163.367
R10996 GND.n4130 GND.n3122 163.367
R10997 GND.n4130 GND.n3112 163.367
R10998 GND.n3112 GND.n3103 163.367
R10999 GND.n4234 GND.n3103 163.367
R11000 GND.n4234 GND.n3101 163.367
R11001 GND.n4238 GND.n3101 163.367
R11002 GND.n4238 GND.n3093 163.367
R11003 GND.n4247 GND.n3093 163.367
R11004 GND.n4247 GND.n3090 163.367
R11005 GND.n4308 GND.n3090 163.367
R11006 GND.n4308 GND.n3091 163.367
R11007 GND.n3091 GND.n3081 163.367
R11008 GND.n4303 GND.n3081 163.367
R11009 GND.n4303 GND.n4301 163.367
R11010 GND.n4301 GND.n4300 163.367
R11011 GND.n4300 GND.n4251 163.367
R11012 GND.n4251 GND.n3063 163.367
R11013 GND.n4295 GND.n3063 163.367
R11014 GND.n3735 GND.n3649 163.367
R11015 GND.n3731 GND.n3649 163.367
R11016 GND.n3729 GND.n3728 163.367
R11017 GND.n3725 GND.n3724 163.367
R11018 GND.n3721 GND.n3720 163.367
R11019 GND.n3717 GND.n3716 163.367
R11020 GND.n3713 GND.n3712 163.367
R11021 GND.n3709 GND.n3708 163.367
R11022 GND.n3704 GND.n3703 163.367
R11023 GND.n3700 GND.n3699 163.367
R11024 GND.n3694 GND.n3693 163.367
R11025 GND.n3690 GND.n3689 163.367
R11026 GND.n3685 GND.n3684 163.367
R11027 GND.n3681 GND.n3680 163.367
R11028 GND.n3677 GND.n3676 163.367
R11029 GND.n3673 GND.n3672 163.367
R11030 GND.n3669 GND.n3668 163.367
R11031 GND.n3665 GND.n3664 163.367
R11032 GND.n3661 GND.n3660 163.367
R11033 GND.n3657 GND.n3407 163.367
R11034 GND.n3757 GND.n3370 163.367
R11035 GND.n3761 GND.n3370 163.367
R11036 GND.n3761 GND.n3361 163.367
R11037 GND.n3770 GND.n3361 163.367
R11038 GND.n3770 GND.n3358 163.367
R11039 GND.n3776 GND.n3358 163.367
R11040 GND.n3776 GND.n3359 163.367
R11041 GND.n3359 GND.n3349 163.367
R11042 GND.n3349 GND.n3337 163.367
R11043 GND.n3797 GND.n3337 163.367
R11044 GND.n3797 GND.n3335 163.367
R11045 GND.n3801 GND.n3335 163.367
R11046 GND.n3801 GND.n3326 163.367
R11047 GND.n3827 GND.n3326 163.367
R11048 GND.n3827 GND.n3323 163.367
R11049 GND.n3836 GND.n3323 163.367
R11050 GND.n3836 GND.n3324 163.367
R11051 GND.n3832 GND.n3324 163.367
R11052 GND.n3832 GND.n3831 163.367
R11053 GND.n3831 GND.n3301 163.367
R11054 GND.n3894 GND.n3301 163.367
R11055 GND.n3894 GND.n3299 163.367
R11056 GND.n3898 GND.n3299 163.367
R11057 GND.n3898 GND.n3285 163.367
R11058 GND.n3918 GND.n3285 163.367
R11059 GND.n3918 GND.n3283 163.367
R11060 GND.n3922 GND.n3283 163.367
R11061 GND.n3922 GND.n3274 163.367
R11062 GND.n3931 GND.n3274 163.367
R11063 GND.n3931 GND.n3271 163.367
R11064 GND.n3937 GND.n3271 163.367
R11065 GND.n3937 GND.n3272 163.367
R11066 GND.n3272 GND.n3261 163.367
R11067 GND.n3261 GND.n3251 163.367
R11068 GND.n3958 GND.n3251 163.367
R11069 GND.n3958 GND.n3249 163.367
R11070 GND.n3962 GND.n3249 163.367
R11071 GND.n3962 GND.n3239 163.367
R11072 GND.n3988 GND.n3239 163.367
R11073 GND.n3988 GND.n3236 163.367
R11074 GND.n3997 GND.n3236 163.367
R11075 GND.n3997 GND.n3237 163.367
R11076 GND.n3993 GND.n3237 163.367
R11077 GND.n3993 GND.n3992 163.367
R11078 GND.n3992 GND.n3213 163.367
R11079 GND.n4054 GND.n3213 163.367
R11080 GND.n4054 GND.n3211 163.367
R11081 GND.n4058 GND.n3211 163.367
R11082 GND.n4058 GND.n3196 163.367
R11083 GND.n4078 GND.n3196 163.367
R11084 GND.n4078 GND.n3194 163.367
R11085 GND.n4082 GND.n3194 163.367
R11086 GND.n4082 GND.n3186 163.367
R11087 GND.n4091 GND.n3186 163.367
R11088 GND.n4091 GND.n3183 163.367
R11089 GND.n4097 GND.n3183 163.367
R11090 GND.n4097 GND.n3184 163.367
R11091 GND.n3184 GND.n3175 163.367
R11092 GND.n3175 GND.n3164 163.367
R11093 GND.n4118 GND.n3164 163.367
R11094 GND.n4118 GND.n3162 163.367
R11095 GND.n4122 GND.n3162 163.367
R11096 GND.n4122 GND.n3152 163.367
R11097 GND.n4148 GND.n3152 163.367
R11098 GND.n4148 GND.n3149 163.367
R11099 GND.n4157 GND.n3149 163.367
R11100 GND.n4157 GND.n3150 163.367
R11101 GND.n4153 GND.n3150 163.367
R11102 GND.n4153 GND.n4152 163.367
R11103 GND.n4152 GND.n3126 163.367
R11104 GND.n4201 GND.n3126 163.367
R11105 GND.n4201 GND.n3124 163.367
R11106 GND.n4205 GND.n3124 163.367
R11107 GND.n4205 GND.n3109 163.367
R11108 GND.n4228 GND.n3109 163.367
R11109 GND.n4228 GND.n3107 163.367
R11110 GND.n4232 GND.n3107 163.367
R11111 GND.n4232 GND.n3099 163.367
R11112 GND.n4241 GND.n3099 163.367
R11113 GND.n4241 GND.n3097 163.367
R11114 GND.n4245 GND.n3097 163.367
R11115 GND.n4245 GND.n3087 163.367
R11116 GND.n4310 GND.n3087 163.367
R11117 GND.n4310 GND.n3084 163.367
R11118 GND.n4319 GND.n3084 163.367
R11119 GND.n4319 GND.n3085 163.367
R11120 GND.n4315 GND.n3085 163.367
R11121 GND.n4315 GND.n4314 163.367
R11122 GND.n4314 GND.n3061 163.367
R11123 GND.n4342 GND.n3061 163.367
R11124 GND.n4342 GND.n3053 163.367
R11125 GND.n2916 GND.t83 154.643
R11126 GND.n5203 GND.t89 154.643
R11127 GND.n3375 GND.n3374 152
R11128 GND.n3059 GND.n3058 152
R11129 GND.n132 GND.t38 151.613
R11130 GND.n145 GND.t6 151.613
R11131 GND.n106 GND.t45 151.613
R11132 GND.n119 GND.t7 151.613
R11133 GND.n80 GND.t8 151.613
R11134 GND.n93 GND.t14 151.613
R11135 GND.n54 GND.t18 151.613
R11136 GND.n67 GND.t27 151.613
R11137 GND.n28 GND.t11 151.613
R11138 GND.n41 GND.t35 151.613
R11139 GND.n3 GND.t3 151.613
R11140 GND.n16 GND.t26 151.613
R11141 GND.n301 GND.t44 151.613
R11142 GND.n288 GND.t17 151.613
R11143 GND.n275 GND.t31 151.613
R11144 GND.n262 GND.t32 151.613
R11145 GND.n249 GND.t22 151.613
R11146 GND.n236 GND.t46 151.613
R11147 GND.n223 GND.t173 151.613
R11148 GND.n210 GND.t29 151.613
R11149 GND.n197 GND.t172 151.613
R11150 GND.n184 GND.t13 151.613
R11151 GND.n172 GND.t40 151.613
R11152 GND.n159 GND.t171 151.613
R11153 GND.n3043 GND.n3042 143.351
R11154 GND.n3696 GND.n3396 143.351
R11155 GND.n3696 GND.n3397 143.351
R11156 GND.n3373 GND.t69 138.431
R11157 GND.n3057 GND.t121 138.431
R11158 GND.n3654 GND.t74 135.282
R11159 GND.n4253 GND.t50 135.282
R11160 GND.n3652 GND.t155 135.282
R11161 GND.n4347 GND.t141 135.282
R11162 GND.n3374 GND.t91 126.766
R11163 GND.n3058 GND.t151 126.766
R11164 GND.n3652 GND.n3651 122.959
R11165 GND.n3654 GND.n3653 122.959
R11166 GND.n4253 GND.n4252 122.959
R11167 GND.n4347 GND.n4346 122.959
R11168 GND.n2916 GND.n2915 121.019
R11169 GND.n5203 GND.n5202 121.019
R11170 GND.n1413 GND.t105 120.76
R11171 GND.n1427 GND.t126 120.76
R11172 GND.n1440 GND.t135 120.76
R11173 GND.n1454 GND.t79 120.76
R11174 GND.n1467 GND.t129 120.76
R11175 GND.n2909 GND.t95 120.76
R11176 GND.n1502 GND.t108 120.76
R11177 GND.n1760 GND.t131 120.76
R11178 GND.n2560 GND.t67 120.76
R11179 GND.n2572 GND.t85 120.76
R11180 GND.n2584 GND.t60 120.76
R11181 GND.n2596 GND.t137 120.76
R11182 GND.n2606 GND.t116 120.76
R11183 GND.n486 GND.t120 120.76
R11184 GND.n494 GND.t111 120.76
R11185 GND.n501 GND.t57 120.76
R11186 GND.n509 GND.t54 120.76
R11187 GND.n517 GND.t147 120.76
R11188 GND.n4678 GND.t102 120.76
R11189 GND.n1838 GND.t98 120.76
R11190 GND.n1803 GND.t113 120.76
R11191 GND.n1793 GND.t143 120.76
R11192 GND.n1910 GND.t64 120.76
R11193 GND.n1770 GND.t149 120.76
R11194 GND.n135 GND.n134 104.615
R11195 GND.n148 GND.n147 104.615
R11196 GND.n109 GND.n108 104.615
R11197 GND.n122 GND.n121 104.615
R11198 GND.n83 GND.n82 104.615
R11199 GND.n96 GND.n95 104.615
R11200 GND.n57 GND.n56 104.615
R11201 GND.n70 GND.n69 104.615
R11202 GND.n31 GND.n30 104.615
R11203 GND.n44 GND.n43 104.615
R11204 GND.n6 GND.n5 104.615
R11205 GND.n19 GND.n18 104.615
R11206 GND.n304 GND.n303 104.615
R11207 GND.n291 GND.n290 104.615
R11208 GND.n278 GND.n277 104.615
R11209 GND.n265 GND.n264 104.615
R11210 GND.n252 GND.n251 104.615
R11211 GND.n239 GND.n238 104.615
R11212 GND.n226 GND.n225 104.615
R11213 GND.n213 GND.n212 104.615
R11214 GND.n200 GND.n199 104.615
R11215 GND.n187 GND.n186 104.615
R11216 GND.n175 GND.n174 104.615
R11217 GND.n162 GND.n161 104.615
R11218 GND.n528 GND.n461 99.6594
R11219 GND.n532 GND.n462 99.6594
R11220 GND.n538 GND.n463 99.6594
R11221 GND.n519 GND.n464 99.6594
R11222 GND.n546 GND.n465 99.6594
R11223 GND.n550 GND.n466 99.6594
R11224 GND.n556 GND.n467 99.6594
R11225 GND.n560 GND.n468 99.6594
R11226 GND.n566 GND.n469 99.6594
R11227 GND.n570 GND.n470 99.6594
R11228 GND.n576 GND.n471 99.6594
R11229 GND.n580 GND.n472 99.6594
R11230 GND.n586 GND.n473 99.6594
R11231 GND.n590 GND.n474 99.6594
R11232 GND.n596 GND.n475 99.6594
R11233 GND.n600 GND.n476 99.6594
R11234 GND.n606 GND.n477 99.6594
R11235 GND.n610 GND.n478 99.6594
R11236 GND.n614 GND.n479 99.6594
R11237 GND.n620 GND.n480 99.6594
R11238 GND.n624 GND.n481 99.6594
R11239 GND.n483 GND.n482 99.6594
R11240 GND.n632 GND.n450 99.6594
R11241 GND.n4956 GND.n4955 99.6594
R11242 GND.n4950 GND.n2521 99.6594
R11243 GND.n4947 GND.n2522 99.6594
R11244 GND.n4943 GND.n2523 99.6594
R11245 GND.n4939 GND.n2524 99.6594
R11246 GND.n4935 GND.n2525 99.6594
R11247 GND.n4931 GND.n2526 99.6594
R11248 GND.n4927 GND.n2527 99.6594
R11249 GND.n4923 GND.n2528 99.6594
R11250 GND.n4920 GND.n2529 99.6594
R11251 GND.n4915 GND.n2531 99.6594
R11252 GND.n4911 GND.n2532 99.6594
R11253 GND.n4906 GND.n2533 99.6594
R11254 GND.n4902 GND.n2534 99.6594
R11255 GND.n4898 GND.n2535 99.6594
R11256 GND.n4894 GND.n2536 99.6594
R11257 GND.n4890 GND.n2537 99.6594
R11258 GND.n4886 GND.n2538 99.6594
R11259 GND.n4882 GND.n2539 99.6594
R11260 GND.n4878 GND.n2540 99.6594
R11261 GND.n4874 GND.n2541 99.6594
R11262 GND.n5190 GND.n1406 99.6594
R11263 GND.n5189 GND.n1409 99.6594
R11264 GND.n5187 GND.n1411 99.6594
R11265 GND.n5186 GND.n1416 99.6594
R11266 GND.n5184 GND.n1418 99.6594
R11267 GND.n5183 GND.n1421 99.6594
R11268 GND.n5181 GND.n1423 99.6594
R11269 GND.n5180 GND.n1428 99.6594
R11270 GND.n5178 GND.n1430 99.6594
R11271 GND.n5176 GND.n1506 99.6594
R11272 GND.n1507 GND.n1435 99.6594
R11273 GND.n1509 GND.n1508 99.6594
R11274 GND.n1510 GND.n1443 99.6594
R11275 GND.n1512 GND.n1511 99.6594
R11276 GND.n1513 GND.n1448 99.6594
R11277 GND.n1515 GND.n1514 99.6594
R11278 GND.n1516 GND.n1455 99.6594
R11279 GND.n1518 GND.n1517 99.6594
R11280 GND.n1519 GND.n1460 99.6594
R11281 GND.n1521 GND.n1520 99.6594
R11282 GND.n1522 GND.n1465 99.6594
R11283 GND.n1523 GND.n1394 99.6594
R11284 GND.n1821 GND.n1280 99.6594
R11285 GND.n1829 GND.n1828 99.6594
R11286 GND.n1832 GND.n1831 99.6594
R11287 GND.n1841 GND.n1840 99.6594
R11288 GND.n1844 GND.n1843 99.6594
R11289 GND.n1851 GND.n1850 99.6594
R11290 GND.n1854 GND.n1853 99.6594
R11291 GND.n1861 GND.n1860 99.6594
R11292 GND.n1864 GND.n1863 99.6594
R11293 GND.n1871 GND.n1870 99.6594
R11294 GND.n1874 GND.n1873 99.6594
R11295 GND.n1881 GND.n1880 99.6594
R11296 GND.n1884 GND.n1883 99.6594
R11297 GND.n1891 GND.n1890 99.6594
R11298 GND.n1894 GND.n1893 99.6594
R11299 GND.n1901 GND.n1900 99.6594
R11300 GND.n1904 GND.n1903 99.6594
R11301 GND.n1913 GND.n1912 99.6594
R11302 GND.n1916 GND.n1915 99.6594
R11303 GND.n1923 GND.n1922 99.6594
R11304 GND.n1926 GND.n1925 99.6594
R11305 GND.n1933 GND.n1932 99.6594
R11306 GND.n4693 GND.n4684 99.6594
R11307 GND.n4697 GND.n4695 99.6594
R11308 GND.n4703 GND.n4680 99.6594
R11309 GND.n4706 GND.n4705 99.6594
R11310 GND.n4959 GND.n4958 99.6594
R11311 GND.n2931 GND.n2547 99.6594
R11312 GND.n2942 GND.n2546 99.6594
R11313 GND.n2912 GND.n2545 99.6594
R11314 GND.n5173 GND.n1479 99.6594
R11315 GND.n5172 GND.n1486 99.6594
R11316 GND.n5170 GND.n5169 99.6594
R11317 GND.n5193 GND.n5192 99.6594
R11318 GND.n1943 GND.n1942 99.6594
R11319 GND.n1950 GND.n1949 99.6594
R11320 GND.n1953 GND.n1952 99.6594
R11321 GND.n1960 GND.n1959 99.6594
R11322 GND.n1942 GND.n1766 99.6594
R11323 GND.n1951 GND.n1950 99.6594
R11324 GND.n1952 GND.n1762 99.6594
R11325 GND.n1961 GND.n1960 99.6594
R11326 GND.n5192 GND.n1504 99.6594
R11327 GND.n5170 GND.n1487 99.6594
R11328 GND.n5172 GND.n5171 99.6594
R11329 GND.n5173 GND.n1478 99.6594
R11330 GND.n4958 GND.n2519 99.6594
R11331 GND.n2941 GND.n2547 99.6594
R11332 GND.n2911 GND.n2546 99.6594
R11333 GND.n2907 GND.n2545 99.6594
R11334 GND.n4705 GND.n4704 99.6594
R11335 GND.n4696 GND.n4680 99.6594
R11336 GND.n4695 GND.n4694 99.6594
R11337 GND.n4686 GND.n4684 99.6594
R11338 GND.n1822 GND.n1821 99.6594
R11339 GND.n1830 GND.n1829 99.6594
R11340 GND.n1831 GND.n1813 99.6594
R11341 GND.n1842 GND.n1841 99.6594
R11342 GND.n1843 GND.n1809 99.6594
R11343 GND.n1852 GND.n1851 99.6594
R11344 GND.n1853 GND.n1805 99.6594
R11345 GND.n1862 GND.n1861 99.6594
R11346 GND.n1863 GND.n1799 99.6594
R11347 GND.n1872 GND.n1871 99.6594
R11348 GND.n1873 GND.n1795 99.6594
R11349 GND.n1882 GND.n1881 99.6594
R11350 GND.n1883 GND.n1788 99.6594
R11351 GND.n1892 GND.n1891 99.6594
R11352 GND.n1893 GND.n1784 99.6594
R11353 GND.n1902 GND.n1901 99.6594
R11354 GND.n1903 GND.n1780 99.6594
R11355 GND.n1914 GND.n1913 99.6594
R11356 GND.n1915 GND.n1776 99.6594
R11357 GND.n1924 GND.n1923 99.6594
R11358 GND.n1925 GND.n1772 99.6594
R11359 GND.n1934 GND.n1933 99.6594
R11360 GND.n1523 GND.n1469 99.6594
R11361 GND.n1522 GND.n1464 99.6594
R11362 GND.n1521 GND.n1461 99.6594
R11363 GND.n1519 GND.n1459 99.6594
R11364 GND.n1518 GND.n1456 99.6594
R11365 GND.n1516 GND.n1452 99.6594
R11366 GND.n1515 GND.n1449 99.6594
R11367 GND.n1513 GND.n1447 99.6594
R11368 GND.n1512 GND.n1444 99.6594
R11369 GND.n1510 GND.n1442 99.6594
R11370 GND.n1509 GND.n1436 99.6594
R11371 GND.n1507 GND.n1434 99.6594
R11372 GND.n5177 GND.n5175 99.6594
R11373 GND.n5178 GND.n1429 99.6594
R11374 GND.n5180 GND.n5179 99.6594
R11375 GND.n5181 GND.n1422 99.6594
R11376 GND.n5183 GND.n5182 99.6594
R11377 GND.n5184 GND.n1417 99.6594
R11378 GND.n5186 GND.n5185 99.6594
R11379 GND.n5187 GND.n1410 99.6594
R11380 GND.n5189 GND.n5188 99.6594
R11381 GND.n5190 GND.n1405 99.6594
R11382 GND.n4956 GND.n2549 99.6594
R11383 GND.n4948 GND.n2521 99.6594
R11384 GND.n4944 GND.n2522 99.6594
R11385 GND.n4940 GND.n2523 99.6594
R11386 GND.n4936 GND.n2524 99.6594
R11387 GND.n4932 GND.n2525 99.6594
R11388 GND.n4928 GND.n2526 99.6594
R11389 GND.n2569 GND.n2527 99.6594
R11390 GND.n4921 GND.n2528 99.6594
R11391 GND.n4916 GND.n2530 99.6594
R11392 GND.n4912 GND.n2531 99.6594
R11393 GND.n4907 GND.n2532 99.6594
R11394 GND.n4903 GND.n2533 99.6594
R11395 GND.n4899 GND.n2534 99.6594
R11396 GND.n4895 GND.n2535 99.6594
R11397 GND.n4891 GND.n2536 99.6594
R11398 GND.n4887 GND.n2537 99.6594
R11399 GND.n4883 GND.n2538 99.6594
R11400 GND.n4879 GND.n2539 99.6594
R11401 GND.n4875 GND.n2540 99.6594
R11402 GND.n2604 GND.n2541 99.6594
R11403 GND.n632 GND.n631 99.6594
R11404 GND.n623 GND.n482 99.6594
R11405 GND.n621 GND.n481 99.6594
R11406 GND.n613 GND.n480 99.6594
R11407 GND.n611 GND.n479 99.6594
R11408 GND.n607 GND.n478 99.6594
R11409 GND.n601 GND.n477 99.6594
R11410 GND.n597 GND.n476 99.6594
R11411 GND.n591 GND.n475 99.6594
R11412 GND.n587 GND.n474 99.6594
R11413 GND.n579 GND.n473 99.6594
R11414 GND.n577 GND.n472 99.6594
R11415 GND.n569 GND.n471 99.6594
R11416 GND.n567 GND.n470 99.6594
R11417 GND.n559 GND.n469 99.6594
R11418 GND.n557 GND.n468 99.6594
R11419 GND.n549 GND.n467 99.6594
R11420 GND.n547 GND.n466 99.6594
R11421 GND.n518 GND.n465 99.6594
R11422 GND.n539 GND.n464 99.6594
R11423 GND.n531 GND.n463 99.6594
R11424 GND.n529 GND.n462 99.6594
R11425 GND.n522 GND.n461 99.6594
R11426 GND.n2918 GND.n2502 99.6594
R11427 GND.n2920 GND.n2919 99.6594
R11428 GND.n2921 GND.n2507 99.6594
R11429 GND.n2923 GND.n2922 99.6594
R11430 GND.n2924 GND.n2512 99.6594
R11431 GND.n2933 GND.n2925 99.6594
R11432 GND.n2927 GND.n2926 99.6594
R11433 GND.n2948 GND.n2917 99.6594
R11434 GND.n4517 GND.n4516 99.6594
R11435 GND.n2949 GND.n2493 99.6594
R11436 GND.n2949 GND.n2904 99.6594
R11437 GND.n4518 GND.n4517 99.6594
R11438 GND.n2948 GND.n2947 99.6594
R11439 GND.n2934 GND.n2926 99.6594
R11440 GND.n2925 GND.n2513 99.6594
R11441 GND.n2924 GND.n2511 99.6594
R11442 GND.n2923 GND.n2508 99.6594
R11443 GND.n2921 GND.n2506 99.6594
R11444 GND.n2920 GND.n2503 99.6594
R11445 GND.n2918 GND.n2498 99.6594
R11446 GND.n3475 GND.n3474 99.6594
R11447 GND.n3481 GND.n3480 99.6594
R11448 GND.n3484 GND.n3483 99.6594
R11449 GND.n3490 GND.n3489 99.6594
R11450 GND.n3488 GND.n3487 99.6594
R11451 GND.n1493 GND.n1474 99.6594
R11452 GND.n1494 GND.n1482 99.6594
R11453 GND.n5200 GND.n5199 99.6594
R11454 GND.n5198 GND.n1496 99.6594
R11455 GND.n1535 GND.n1496 99.6594
R11456 GND.n5201 GND.n5200 99.6594
R11457 GND.n3476 GND.n3475 99.6594
R11458 GND.n3482 GND.n3481 99.6594
R11459 GND.n3485 GND.n3484 99.6594
R11460 GND.n3491 GND.n3490 99.6594
R11461 GND.n3487 GND.n1473 99.6594
R11462 GND.n1493 GND.n1492 99.6594
R11463 GND.n1494 GND.n1483 99.6594
R11464 GND.n1413 GND.n1412 74.4732
R11465 GND.n1427 GND.n1426 74.4732
R11466 GND.n1440 GND.n1439 74.4732
R11467 GND.n1454 GND.n1453 74.4732
R11468 GND.n1467 GND.n1466 74.4732
R11469 GND.n2909 GND.n2908 74.4732
R11470 GND.n1502 GND.n1501 74.4732
R11471 GND.n1760 GND.n1759 74.4732
R11472 GND.n2560 GND.n2559 74.4732
R11473 GND.n2572 GND.n2571 74.4732
R11474 GND.n2584 GND.n2583 74.4732
R11475 GND.n2596 GND.n2595 74.4732
R11476 GND.n2606 GND.n2605 74.4732
R11477 GND.n486 GND.n485 74.4732
R11478 GND.n494 GND.n493 74.4732
R11479 GND.n501 GND.n500 74.4732
R11480 GND.n509 GND.n508 74.4732
R11481 GND.n517 GND.n516 74.4732
R11482 GND.n4678 GND.n4677 74.4732
R11483 GND.n1838 GND.n1837 74.4732
R11484 GND.n1803 GND.n1802 74.4732
R11485 GND.n1793 GND.n1792 74.4732
R11486 GND.n1910 GND.n1909 74.4732
R11487 GND.n1770 GND.n1769 74.4732
R11488 GND.n3373 GND.n3372 73.571
R11489 GND.n3057 GND.n3056 73.571
R11490 GND.n4383 GND.n3052 71.676
R11491 GND.n4379 GND.n3051 71.676
R11492 GND.n4375 GND.n3050 71.676
R11493 GND.n4371 GND.n3049 71.676
R11494 GND.n4367 GND.n3048 71.676
R11495 GND.n4363 GND.n3047 71.676
R11496 GND.n4359 GND.n3046 71.676
R11497 GND.n4354 GND.n3045 71.676
R11498 GND.n4350 GND.n3044 71.676
R11499 GND.n3042 GND.n3031 71.676
R11500 GND.n4258 GND.n3032 71.676
R11501 GND.n4262 GND.n3033 71.676
R11502 GND.n4266 GND.n3034 71.676
R11503 GND.n4270 GND.n3035 71.676
R11504 GND.n4274 GND.n3036 71.676
R11505 GND.n4278 GND.n3037 71.676
R11506 GND.n4282 GND.n3038 71.676
R11507 GND.n4286 GND.n3039 71.676
R11508 GND.n4290 GND.n3040 71.676
R11509 GND.n4294 GND.n3041 71.676
R11510 GND.n3736 GND.n3377 71.676
R11511 GND.n3731 GND.n3388 71.676
R11512 GND.n3728 GND.n3389 71.676
R11513 GND.n3724 GND.n3390 71.676
R11514 GND.n3720 GND.n3391 71.676
R11515 GND.n3716 GND.n3392 71.676
R11516 GND.n3712 GND.n3393 71.676
R11517 GND.n3708 GND.n3394 71.676
R11518 GND.n3703 GND.n3395 71.676
R11519 GND.n3699 GND.n3396 71.676
R11520 GND.n3693 GND.n3398 71.676
R11521 GND.n3689 GND.n3399 71.676
R11522 GND.n3684 GND.n3400 71.676
R11523 GND.n3680 GND.n3401 71.676
R11524 GND.n3676 GND.n3402 71.676
R11525 GND.n3672 GND.n3403 71.676
R11526 GND.n3668 GND.n3404 71.676
R11527 GND.n3664 GND.n3405 71.676
R11528 GND.n3660 GND.n3406 71.676
R11529 GND.n3736 GND.n3735 71.676
R11530 GND.n3729 GND.n3388 71.676
R11531 GND.n3725 GND.n3389 71.676
R11532 GND.n3721 GND.n3390 71.676
R11533 GND.n3717 GND.n3391 71.676
R11534 GND.n3713 GND.n3392 71.676
R11535 GND.n3709 GND.n3393 71.676
R11536 GND.n3704 GND.n3394 71.676
R11537 GND.n3700 GND.n3395 71.676
R11538 GND.n3694 GND.n3397 71.676
R11539 GND.n3690 GND.n3398 71.676
R11540 GND.n3685 GND.n3399 71.676
R11541 GND.n3681 GND.n3400 71.676
R11542 GND.n3677 GND.n3401 71.676
R11543 GND.n3673 GND.n3402 71.676
R11544 GND.n3669 GND.n3403 71.676
R11545 GND.n3665 GND.n3404 71.676
R11546 GND.n3661 GND.n3405 71.676
R11547 GND.n3657 GND.n3406 71.676
R11548 GND.n4291 GND.n3041 71.676
R11549 GND.n4287 GND.n3040 71.676
R11550 GND.n4283 GND.n3039 71.676
R11551 GND.n4279 GND.n3038 71.676
R11552 GND.n4275 GND.n3037 71.676
R11553 GND.n4271 GND.n3036 71.676
R11554 GND.n4267 GND.n3035 71.676
R11555 GND.n4263 GND.n3034 71.676
R11556 GND.n4259 GND.n3033 71.676
R11557 GND.n4255 GND.n3032 71.676
R11558 GND.n4349 GND.n3043 71.676
R11559 GND.n4353 GND.n3044 71.676
R11560 GND.n4358 GND.n3045 71.676
R11561 GND.n4362 GND.n3046 71.676
R11562 GND.n4366 GND.n3047 71.676
R11563 GND.n4370 GND.n3048 71.676
R11564 GND.n4374 GND.n3049 71.676
R11565 GND.n4378 GND.n3050 71.676
R11566 GND.n4382 GND.n3051 71.676
R11567 GND.n3054 GND.n3052 71.676
R11568 GND.n141 GND.n140 68.2805
R11569 GND.n115 GND.n114 68.2805
R11570 GND.n89 GND.n88 68.2805
R11571 GND.n63 GND.n62 68.2805
R11572 GND.n37 GND.n36 68.2805
R11573 GND.n12 GND.n11 68.2805
R11574 GND.n297 GND.n296 68.2805
R11575 GND.n271 GND.n270 68.2805
R11576 GND.n245 GND.n244 68.2805
R11577 GND.n219 GND.n218 68.2805
R11578 GND.n193 GND.n192 68.2805
R11579 GND.n168 GND.n167 68.2805
R11580 GND.n3376 GND.n3375 63.641
R11581 GND.n3706 GND.n3652 59.5399
R11582 GND.n3687 GND.n3654 59.5399
R11583 GND.n4254 GND.n4253 59.5399
R11584 GND.n4356 GND.n4347 59.5399
R11585 GND.n134 GND.t38 52.3082
R11586 GND.n147 GND.t6 52.3082
R11587 GND.n108 GND.t45 52.3082
R11588 GND.n121 GND.t7 52.3082
R11589 GND.n82 GND.t8 52.3082
R11590 GND.n95 GND.t14 52.3082
R11591 GND.n56 GND.t18 52.3082
R11592 GND.n69 GND.t27 52.3082
R11593 GND.n30 GND.t11 52.3082
R11594 GND.n43 GND.t35 52.3082
R11595 GND.n5 GND.t3 52.3082
R11596 GND.n18 GND.t26 52.3082
R11597 GND.n303 GND.t44 52.3082
R11598 GND.n290 GND.t17 52.3082
R11599 GND.n277 GND.t31 52.3082
R11600 GND.n264 GND.t32 52.3082
R11601 GND.n251 GND.t22 52.3082
R11602 GND.n238 GND.t46 52.3082
R11603 GND.n225 GND.t173 52.3082
R11604 GND.n212 GND.t29 52.3082
R11605 GND.n199 GND.t172 52.3082
R11606 GND.n186 GND.t13 52.3082
R11607 GND.n174 GND.t40 52.3082
R11608 GND.n161 GND.t171 52.3082
R11609 GND.n4345 GND.n3059 44.3322
R11610 GND.n4519 GND.n2916 42.2793
R11611 GND.n1414 GND.n1413 42.2793
R11612 GND.n5265 GND.n1427 42.2793
R11613 GND.n1441 GND.n1440 42.2793
R11614 GND.n5239 GND.n1454 42.2793
R11615 GND.n5226 GND.n1467 42.2793
R11616 GND.n4523 GND.n2909 42.2793
R11617 GND.n1503 GND.n1502 42.2793
R11618 GND.n1761 GND.n1760 42.2793
R11619 GND.n4942 GND.n2560 42.2793
R11620 GND.n4925 GND.n2572 42.2793
R11621 GND.n4909 GND.n2584 42.2793
R11622 GND.n4889 GND.n2596 42.2793
R11623 GND.n2607 GND.n2606 42.2793
R11624 GND.n630 GND.n486 42.2793
R11625 GND.n609 GND.n494 42.2793
R11626 GND.n502 GND.n501 42.2793
R11627 GND.n510 GND.n509 42.2793
R11628 GND.n541 GND.n517 42.2793
R11629 GND.n4679 GND.n4678 42.2793
R11630 GND.n1839 GND.n1838 42.2793
R11631 GND.n1804 GND.n1803 42.2793
R11632 GND.n1794 GND.n1793 42.2793
R11633 GND.n1911 GND.n1910 42.2793
R11634 GND.n1771 GND.n1770 42.2793
R11635 GND.n5204 GND.n5203 42.2793
R11636 GND.n5517 GND.n1139 42.0897
R11637 GND.n5511 GND.n1139 42.0897
R11638 GND.n5511 GND.n5510 42.0897
R11639 GND.n5510 GND.n5509 42.0897
R11640 GND.n5509 GND.n1146 42.0897
R11641 GND.n5503 GND.n1146 42.0897
R11642 GND.n5503 GND.n5502 42.0897
R11643 GND.n5502 GND.n5501 42.0897
R11644 GND.n5501 GND.n1154 42.0897
R11645 GND.n5495 GND.n1154 42.0897
R11646 GND.n5495 GND.n5494 42.0897
R11647 GND.n5494 GND.n5493 42.0897
R11648 GND.n5493 GND.n1162 42.0897
R11649 GND.n5487 GND.n1162 42.0897
R11650 GND.n5487 GND.n5486 42.0897
R11651 GND.n5486 GND.n5485 42.0897
R11652 GND.n5485 GND.n1170 42.0897
R11653 GND.n5479 GND.n1170 42.0897
R11654 GND.n5479 GND.n5478 42.0897
R11655 GND.n5478 GND.n5477 42.0897
R11656 GND.n5477 GND.n1178 42.0897
R11657 GND.n5471 GND.n1178 42.0897
R11658 GND.n5471 GND.n5470 42.0897
R11659 GND.n5470 GND.n5469 42.0897
R11660 GND.n5469 GND.n1186 42.0897
R11661 GND.n5463 GND.n1186 42.0897
R11662 GND.n5463 GND.n5462 42.0897
R11663 GND.n5462 GND.n5461 42.0897
R11664 GND.n5461 GND.n1194 42.0897
R11665 GND.n5455 GND.n1194 42.0897
R11666 GND.n5455 GND.n5454 42.0897
R11667 GND.n5454 GND.n5453 42.0897
R11668 GND.n5453 GND.n1202 42.0897
R11669 GND.n5447 GND.n1202 42.0897
R11670 GND.n5447 GND.n5446 42.0897
R11671 GND.n5446 GND.n5445 42.0897
R11672 GND.n5445 GND.n1210 42.0897
R11673 GND.n5439 GND.n1210 42.0897
R11674 GND.n5439 GND.n5438 42.0897
R11675 GND.n5438 GND.n5437 42.0897
R11676 GND.n5437 GND.n1218 42.0897
R11677 GND.n5431 GND.n1218 42.0897
R11678 GND.n5431 GND.n5430 42.0897
R11679 GND.n5430 GND.n5429 42.0897
R11680 GND.n5429 GND.n1226 42.0897
R11681 GND.n5423 GND.n1226 42.0897
R11682 GND.n5423 GND.n5422 42.0897
R11683 GND.n5422 GND.n5421 42.0897
R11684 GND.n1242 GND.n1234 39.0838
R11685 GND.n5412 GND.n1242 39.0838
R11686 GND.n5412 GND.n5411 39.0838
R11687 GND.n5411 GND.n5410 39.0838
R11688 GND.n5410 GND.n1243 39.0838
R11689 GND.n5404 GND.n1243 39.0838
R11690 GND.n5404 GND.n5403 39.0838
R11691 GND.n5403 GND.n5402 39.0838
R11692 GND.n5402 GND.n1251 39.0838
R11693 GND.n5396 GND.n1251 39.0838
R11694 GND.n5396 GND.n5395 39.0838
R11695 GND.n5395 GND.n5394 39.0838
R11696 GND.n5394 GND.n1259 39.0838
R11697 GND.n5388 GND.n1259 39.0838
R11698 GND.n5388 GND.n5387 39.0838
R11699 GND.n5387 GND.n5386 39.0838
R11700 GND.n5380 GND.n1275 39.0838
R11701 GND.n1505 GND.n1397 39.0838
R11702 GND.n5168 GND.n1524 39.0838
R11703 GND.n5162 GND.n1524 39.0838
R11704 GND.n5160 GND.n5159 39.0838
R11705 GND.n5159 GND.n1534 39.0838
R11706 GND.n3511 GND.n1534 39.0838
R11707 GND.n3524 GND.n3511 39.0838
R11708 GND.n3524 GND.n3467 39.0838
R11709 GND.n3534 GND.n3467 39.0838
R11710 GND.n3534 GND.n3532 39.0838
R11711 GND.n3542 GND.n3456 39.0838
R11712 GND.n3551 GND.n3456 39.0838
R11713 GND.n3551 GND.n3450 39.0838
R11714 GND.n3559 GND.n3450 39.0838
R11715 GND.n3559 GND.n3444 39.0838
R11716 GND.n3568 GND.n3444 39.0838
R11717 GND.n3568 GND.n3438 39.0838
R11718 GND.n3576 GND.n3438 39.0838
R11719 GND.n3576 GND.n3432 39.0838
R11720 GND.n3585 GND.n3432 39.0838
R11721 GND.n3585 GND.n3426 39.0838
R11722 GND.n3593 GND.n3426 39.0838
R11723 GND.n3593 GND.n3419 39.0838
R11724 GND.n3603 GND.n3419 39.0838
R11725 GND.n3611 GND.n3413 39.0838
R11726 GND.n3611 GND.n3386 39.0838
R11727 GND.n3739 GND.n3386 39.0838
R11728 GND.n4398 GND.n3023 39.0838
R11729 GND.n4398 GND.n3017 39.0838
R11730 GND.n4407 GND.n3017 39.0838
R11731 GND.n4415 GND.n3011 39.0838
R11732 GND.n4415 GND.n3005 39.0838
R11733 GND.n4424 GND.n3005 39.0838
R11734 GND.n4424 GND.n2999 39.0838
R11735 GND.n4432 GND.n2999 39.0838
R11736 GND.n4432 GND.n2993 39.0838
R11737 GND.n4441 GND.n2993 39.0838
R11738 GND.n4441 GND.n2987 39.0838
R11739 GND.n4449 GND.n2987 39.0838
R11740 GND.n4449 GND.n2981 39.0838
R11741 GND.n4458 GND.n2981 39.0838
R11742 GND.n4458 GND.n2974 39.0838
R11743 GND.n4466 GND.n2974 39.0838
R11744 GND.n4466 GND.n2975 39.0838
R11745 GND.n4475 GND.n2963 39.0838
R11746 GND.n4486 GND.n2963 39.0838
R11747 GND.n4486 GND.n2957 39.0838
R11748 GND.n4495 GND.n2957 39.0838
R11749 GND.n4495 GND.n2494 39.0838
R11750 GND.n4982 GND.n2494 39.0838
R11751 GND.n4982 GND.n2496 39.0838
R11752 GND.n4514 GND.n2950 39.0838
R11753 GND.n2950 GND.n2520 39.0838
R11754 GND.n2612 GND.n2543 39.0838
R11755 GND.n6349 GND.n452 39.0838
R11756 GND.n6343 GND.n6342 39.0838
R11757 GND.n6342 GND.n6341 39.0838
R11758 GND.n6341 GND.n634 39.0838
R11759 GND.n6335 GND.n634 39.0838
R11760 GND.n6335 GND.n6334 39.0838
R11761 GND.n6334 GND.n6333 39.0838
R11762 GND.n6333 GND.n642 39.0838
R11763 GND.n6327 GND.n642 39.0838
R11764 GND.n6327 GND.n6326 39.0838
R11765 GND.n6326 GND.n6325 39.0838
R11766 GND.n6325 GND.n650 39.0838
R11767 GND.n6319 GND.n650 39.0838
R11768 GND.n6319 GND.n6318 39.0838
R11769 GND.n6318 GND.n6317 39.0838
R11770 GND.n6317 GND.n658 39.0838
R11771 GND.n6311 GND.n658 39.0838
R11772 GND.n141 GND.n139 35.4957
R11773 GND.n115 GND.n113 35.4957
R11774 GND.n89 GND.n87 35.4957
R11775 GND.n63 GND.n61 35.4957
R11776 GND.n37 GND.n35 35.4957
R11777 GND.n12 GND.n10 35.4957
R11778 GND.n297 GND.n295 35.4957
R11779 GND.n271 GND.n269 35.4957
R11780 GND.n245 GND.n243 35.4957
R11781 GND.n219 GND.n217 35.4957
R11782 GND.n193 GND.n191 35.4957
R11783 GND.n168 GND.n166 35.4957
R11784 GND.n3374 GND.n3373 34.8345
R11785 GND.n3058 GND.n3057 34.8345
R11786 GND.n153 GND.n152 32.1853
R11787 GND.n127 GND.n126 32.1853
R11788 GND.n101 GND.n100 32.1853
R11789 GND.n75 GND.n74 32.1853
R11790 GND.n49 GND.n48 32.1853
R11791 GND.n24 GND.n23 32.1853
R11792 GND.n309 GND.n308 32.1853
R11793 GND.n283 GND.n282 32.1853
R11794 GND.n257 GND.n256 32.1853
R11795 GND.n231 GND.n230 32.1853
R11796 GND.n205 GND.n204 32.1853
R11797 GND.n180 GND.n179 32.1853
R11798 GND.n4296 GND.n4293 31.3761
R11799 GND.n3656 GND.n3655 31.3761
R11800 GND.n5160 GND.n1495 28.5313
R11801 GND.n4515 GND.n2496 28.5313
R11802 GND.n3532 GND.t88 26.968
R11803 GND.n4475 GND.t81 26.968
R11804 GND.n3762 GND.n3367 26.5772
R11805 GND.n3769 GND.n3768 26.5772
R11806 GND.n3785 GND.n3348 26.5772
R11807 GND.n3785 GND.n3351 26.5772
R11808 GND.n3802 GND.n3332 26.5772
R11809 GND.n3826 GND.n3319 26.5772
R11810 GND.n3819 GND.n3310 26.5772
R11811 GND.n3893 GND.n3302 26.5772
R11812 GND.n3899 GND.n3298 26.5772
R11813 GND.n3923 GND.n3279 26.5772
R11814 GND.n3930 GND.n3929 26.5772
R11815 GND.n3946 GND.n3260 26.5772
R11816 GND.n3946 GND.n3263 26.5772
R11817 GND.n3963 GND.n3246 26.5772
R11818 GND.n3987 GND.n3232 26.5772
R11819 GND.n3980 GND.n3222 26.5772
R11820 GND.n4053 GND.n3214 26.5772
R11821 GND.n4059 GND.n3210 26.5772
R11822 GND.n4083 GND.n3191 26.5772
R11823 GND.n4090 GND.n4089 26.5772
R11824 GND.n4106 GND.n3174 26.5772
R11825 GND.n4106 GND.n3177 26.5772
R11826 GND.n4123 GND.n3158 26.5772
R11827 GND.n4147 GND.n3145 26.5772
R11828 GND.n4140 GND.n3135 26.5772
R11829 GND.n4200 GND.n3127 26.5772
R11830 GND.n4206 GND.n3123 26.5772
R11831 GND.n4233 GND.n3104 26.5772
R11832 GND.n4240 GND.n4239 26.5772
R11833 GND.n4309 GND.n3088 26.5772
R11834 GND.n4309 GND.n3079 26.5772
R11835 GND.n4302 GND.n3070 26.5772
R11836 GND.n4341 GND.n3062 26.5772
R11837 GND.t159 GND.n3413 25.4047
R11838 GND.n4407 GND.t162 25.4047
R11839 GND.n3777 GND.n3356 25.0138
R11840 GND.n3796 GND.n3795 25.0138
R11841 GND.n3938 GND.n3269 25.0138
R11842 GND.n3957 GND.n3956 25.0138
R11843 GND.n4098 GND.n3182 25.0138
R11844 GND.n4117 GND.n4116 25.0138
R11845 GND.n4246 GND.n3095 25.0138
R11846 GND.n4320 GND.n3083 25.0138
R11847 GND.n3737 GND.n3648 23.8413
R11848 GND.n4390 GND.n4388 23.8413
R11849 GND.n5386 GND.n1267 23.4505
R11850 GND.n5191 GND.n5168 23.4505
R11851 GND.n3282 GND.n3280 23.4505
R11852 GND.n3247 GND.n3241 23.4505
R11853 GND.n3193 GND.n3192 23.4505
R11854 GND.n3159 GND.n3153 23.4505
R11855 GND.n3073 GND.n3071 23.4505
R11856 GND.n4957 GND.n2520 23.4505
R11857 GND.n6343 GND.n633 23.4505
R11858 GND.t70 GND.n3368 21.8872
R11859 GND.n3837 GND.n3322 21.8872
R11860 GND.n3917 GND.n3286 21.8872
R11861 GND.n3998 GND.n3235 21.8872
R11862 GND.n4077 GND.n3197 21.8872
R11863 GND.n4158 GND.n3148 21.8872
R11864 GND.n4227 GND.n3111 21.8872
R11865 GND.n4390 GND.n3029 21.8872
R11866 GND.n3313 GND.n3311 20.3238
R11867 GND.n3892 GND.n3295 20.3238
R11868 GND.n3226 GND.n3223 20.3238
R11869 GND.n4052 GND.n3207 20.3238
R11870 GND.n3139 GND.n3136 20.3238
R11871 GND.n4199 GND.n3120 20.3238
R11872 GND.n3371 GND.t93 19.8005
R11873 GND.n3371 GND.t71 19.8005
R11874 GND.n3055 GND.t123 19.8005
R11875 GND.n3055 GND.t153 19.8005
R11876 GND.n5380 GND.n5379 19.5422
R11877 GND.n5379 GND.n1278 19.5422
R11878 GND.n1755 GND.n1278 19.5422
R11879 GND.n1755 GND.n1287 19.5422
R11880 GND.n5373 GND.n1287 19.5422
R11881 GND.n5373 GND.n1290 19.5422
R11882 GND.n1972 GND.n1290 19.5422
R11883 GND.n1973 GND.n1972 19.5422
R11884 GND.n2012 GND.n1973 19.5422
R11885 GND.n2004 GND.n2002 19.5422
R11886 GND.n2004 GND.n1749 19.5422
R11887 GND.n2021 GND.n1749 19.5422
R11888 GND.n2021 GND.n1745 19.5422
R11889 GND.n2027 GND.n1745 19.5422
R11890 GND.n2027 GND.n1747 19.5422
R11891 GND.n2023 GND.n1747 19.5422
R11892 GND.n2023 GND.n1734 19.5422
R11893 GND.n2037 GND.n1734 19.5422
R11894 GND.n2037 GND.n1736 19.5422
R11895 GND.n1736 GND.n1727 19.5422
R11896 GND.n2047 GND.n1727 19.5422
R11897 GND.n2047 GND.n2046 19.5422
R11898 GND.n2046 GND.n1715 19.5422
R11899 GND.n2080 GND.n1715 19.5422
R11900 GND.n2080 GND.n1717 19.5422
R11901 GND.n2077 GND.n1717 19.5422
R11902 GND.n2077 GND.n2076 19.5422
R11903 GND.n2090 GND.n1706 19.5422
R11904 GND.n1709 GND.n1706 19.5422
R11905 GND.n1709 GND.n1699 19.5422
R11906 GND.n2099 GND.n1699 19.5422
R11907 GND.n2099 GND.n1693 19.5422
R11908 GND.n2104 GND.n1693 19.5422
R11909 GND.n2104 GND.n1696 19.5422
R11910 GND.n2101 GND.n1696 19.5422
R11911 GND.n2101 GND.n1683 19.5422
R11912 GND.n2112 GND.n1683 19.5422
R11913 GND.n2112 GND.n1685 19.5422
R11914 GND.n1685 GND.n1684 19.5422
R11915 GND.n1684 GND.n1644 19.5422
R11916 GND.n2211 GND.n1644 19.5422
R11917 GND.n2211 GND.n1647 19.5422
R11918 GND.n2208 GND.n2207 19.5422
R11919 GND.n2207 GND.n1652 19.5422
R11920 GND.n1658 GND.n1652 19.5422
R11921 GND.n1659 GND.n1658 19.5422
R11922 GND.n2200 GND.n1659 19.5422
R11923 GND.n2200 GND.n2199 19.5422
R11924 GND.n2199 GND.n1662 19.5422
R11925 GND.n2194 GND.n1662 19.5422
R11926 GND.n2194 GND.n1670 19.5422
R11927 GND.n2191 GND.n1670 19.5422
R11928 GND.n2191 GND.n2190 19.5422
R11929 GND.n2190 GND.n2136 19.5422
R11930 GND.n2141 GND.n2136 19.5422
R11931 GND.n2141 GND.n2140 19.5422
R11932 GND.n2220 GND.n1627 19.5422
R11933 GND.n2220 GND.n1628 19.5422
R11934 GND.n1631 GND.n1628 19.5422
R11935 GND.n1631 GND.n1620 19.5422
R11936 GND.n2229 GND.n1620 19.5422
R11937 GND.n2229 GND.n1614 19.5422
R11938 GND.n2234 GND.n1614 19.5422
R11939 GND.n2234 GND.n1617 19.5422
R11940 GND.n2231 GND.n1617 19.5422
R11941 GND.n2231 GND.n1603 19.5422
R11942 GND.n2244 GND.n1603 19.5422
R11943 GND.n2244 GND.n1604 19.5422
R11944 GND.n1608 GND.n1604 19.5422
R11945 GND.n1608 GND.n1595 19.5422
R11946 GND.n2253 GND.n1595 19.5422
R11947 GND.n2259 GND.n1591 19.5422
R11948 GND.n2259 GND.n1593 19.5422
R11949 GND.n2256 GND.n1593 19.5422
R11950 GND.n2256 GND.n1580 19.5422
R11951 GND.n2269 GND.n1580 19.5422
R11952 GND.n2269 GND.n1581 19.5422
R11953 GND.n1585 GND.n1581 19.5422
R11954 GND.n1585 GND.n1573 19.5422
R11955 GND.n2292 GND.n1573 19.5422
R11956 GND.n2292 GND.n1569 19.5422
R11957 GND.n2297 GND.n1569 19.5422
R11958 GND.n2297 GND.n1571 19.5422
R11959 GND.n1571 GND.n1561 19.5422
R11960 GND.n2306 GND.n1561 19.5422
R11961 GND.n2306 GND.n2305 19.5422
R11962 GND.n2305 GND.n1553 19.5422
R11963 GND.n2330 GND.n1553 19.5422
R11964 GND.n2330 GND.n2329 19.5422
R11965 GND.n2334 GND.n1551 19.5422
R11966 GND.n2278 GND.n1551 19.5422
R11967 GND.n2278 GND.n1543 19.5422
R11968 GND.n2342 GND.n1543 19.5422
R11969 GND.n2342 GND.n1541 19.5422
R11970 GND.n2345 GND.n1541 19.5422
R11971 GND.n2345 GND.n1395 19.5422
R11972 GND.n5294 GND.n1395 19.5422
R11973 GND.n5294 GND.n1397 19.5422
R11974 GND.n4864 GND.n2612 19.5422
R11975 GND.n4864 GND.n4863 19.5422
R11976 GND.n4863 GND.n2614 19.5422
R11977 GND.n2623 GND.n2614 19.5422
R11978 GND.n2624 GND.n2623 19.5422
R11979 GND.n4857 GND.n2624 19.5422
R11980 GND.n4857 GND.n4856 19.5422
R11981 GND.n4856 GND.n2627 19.5422
R11982 GND.n4551 GND.n2627 19.5422
R11983 GND.n4850 GND.n2643 19.5422
R11984 GND.n4850 GND.n2646 19.5422
R11985 GND.n4559 GND.n2646 19.5422
R11986 GND.n4559 GND.n2655 19.5422
R11987 GND.n4844 GND.n2655 19.5422
R11988 GND.n4844 GND.n2658 19.5422
R11989 GND.n4566 GND.n2658 19.5422
R11990 GND.n4566 GND.n2666 19.5422
R11991 GND.n4838 GND.n2666 19.5422
R11992 GND.n4838 GND.n2669 19.5422
R11993 GND.n4574 GND.n2669 19.5422
R11994 GND.n4574 GND.n2676 19.5422
R11995 GND.n4832 GND.n2676 19.5422
R11996 GND.n4832 GND.n2679 19.5422
R11997 GND.n4581 GND.n2679 19.5422
R11998 GND.n4581 GND.n2687 19.5422
R11999 GND.n4826 GND.n2687 19.5422
R12000 GND.n4826 GND.n2690 19.5422
R12001 GND.n4589 GND.n2697 19.5422
R12002 GND.n4820 GND.n2697 19.5422
R12003 GND.n4820 GND.n2700 19.5422
R12004 GND.n4596 GND.n2700 19.5422
R12005 GND.n4596 GND.n2708 19.5422
R12006 GND.n4814 GND.n2708 19.5422
R12007 GND.n4814 GND.n2711 19.5422
R12008 GND.n4604 GND.n2711 19.5422
R12009 GND.n4604 GND.n2718 19.5422
R12010 GND.n4808 GND.n2718 19.5422
R12011 GND.n4808 GND.n2721 19.5422
R12012 GND.n4611 GND.n2721 19.5422
R12013 GND.n4611 GND.n2727 19.5422
R12014 GND.n4802 GND.n2727 19.5422
R12015 GND.n4802 GND.n2730 19.5422
R12016 GND.n4623 GND.n2737 19.5422
R12017 GND.n4796 GND.n2737 19.5422
R12018 GND.n4796 GND.n2740 19.5422
R12019 GND.n4793 GND.n2740 19.5422
R12020 GND.n4793 GND.n4792 19.5422
R12021 GND.n4792 GND.n2744 19.5422
R12022 GND.n2744 GND.n317 19.5422
R12023 GND.n6424 GND.n317 19.5422
R12024 GND.n6424 GND.n319 19.5422
R12025 GND.n2872 GND.n319 19.5422
R12026 GND.n4784 GND.n2872 19.5422
R12027 GND.n4784 GND.n4783 19.5422
R12028 GND.n4783 GND.n2875 19.5422
R12029 GND.n4774 GND.n2875 19.5422
R12030 GND.n6417 GND.n336 19.5422
R12031 GND.n6417 GND.n339 19.5422
R12032 GND.n4768 GND.n339 19.5422
R12033 GND.n4768 GND.n348 19.5422
R12034 GND.n6411 GND.n348 19.5422
R12035 GND.n6411 GND.n351 19.5422
R12036 GND.n4762 GND.n351 19.5422
R12037 GND.n4762 GND.n358 19.5422
R12038 GND.n6405 GND.n358 19.5422
R12039 GND.n6405 GND.n361 19.5422
R12040 GND.n4756 GND.n361 19.5422
R12041 GND.n4756 GND.n368 19.5422
R12042 GND.n6399 GND.n368 19.5422
R12043 GND.n6399 GND.n371 19.5422
R12044 GND.n4750 GND.n371 19.5422
R12045 GND.n6393 GND.n379 19.5422
R12046 GND.n6393 GND.n382 19.5422
R12047 GND.n4744 GND.n382 19.5422
R12048 GND.n4744 GND.n389 19.5422
R12049 GND.n6387 GND.n389 19.5422
R12050 GND.n6387 GND.n392 19.5422
R12051 GND.n4738 GND.n392 19.5422
R12052 GND.n4738 GND.n400 19.5422
R12053 GND.n6381 GND.n400 19.5422
R12054 GND.n6381 GND.n403 19.5422
R12055 GND.n4732 GND.n403 19.5422
R12056 GND.n4732 GND.n410 19.5422
R12057 GND.n6375 GND.n410 19.5422
R12058 GND.n6375 GND.n413 19.5422
R12059 GND.n4726 GND.n413 19.5422
R12060 GND.n4726 GND.n421 19.5422
R12061 GND.n6369 GND.n421 19.5422
R12062 GND.n6369 GND.n424 19.5422
R12063 GND.n4720 GND.n431 19.5422
R12064 GND.n6363 GND.n431 19.5422
R12065 GND.n6363 GND.n434 19.5422
R12066 GND.n4714 GND.n434 19.5422
R12067 GND.n4714 GND.n442 19.5422
R12068 GND.n6357 GND.n442 19.5422
R12069 GND.n6357 GND.n445 19.5422
R12070 GND.n6350 GND.n445 19.5422
R12071 GND.n6350 GND.n6349 19.5422
R12072 GND.n5197 GND.n1490 19.3944
R12073 GND.n5197 GND.n1497 19.3944
R12074 GND.n5157 GND.n1537 19.3944
R12075 GND.n5153 GND.n1537 19.3944
R12076 GND.n5153 GND.n5152 19.3944
R12077 GND.n5152 GND.n5151 19.3944
R12078 GND.n5151 GND.n2355 19.3944
R12079 GND.n5147 GND.n2355 19.3944
R12080 GND.n5147 GND.n5146 19.3944
R12081 GND.n5146 GND.n5145 19.3944
R12082 GND.n5145 GND.n2360 19.3944
R12083 GND.n5141 GND.n2360 19.3944
R12084 GND.n5141 GND.n5140 19.3944
R12085 GND.n5140 GND.n5139 19.3944
R12086 GND.n5139 GND.n2365 19.3944
R12087 GND.n5135 GND.n2365 19.3944
R12088 GND.n5135 GND.n5134 19.3944
R12089 GND.n5134 GND.n5133 19.3944
R12090 GND.n5133 GND.n2370 19.3944
R12091 GND.n5129 GND.n2370 19.3944
R12092 GND.n5129 GND.n5128 19.3944
R12093 GND.n5128 GND.n5127 19.3944
R12094 GND.n5127 GND.n2375 19.3944
R12095 GND.n5123 GND.n2375 19.3944
R12096 GND.n5123 GND.n5122 19.3944
R12097 GND.n5122 GND.n5121 19.3944
R12098 GND.n5121 GND.n2380 19.3944
R12099 GND.n5117 GND.n2380 19.3944
R12100 GND.n5117 GND.n5116 19.3944
R12101 GND.n5116 GND.n5115 19.3944
R12102 GND.n5115 GND.n2385 19.3944
R12103 GND.n5111 GND.n2385 19.3944
R12104 GND.n5111 GND.n5110 19.3944
R12105 GND.n5110 GND.n5109 19.3944
R12106 GND.n5109 GND.n2390 19.3944
R12107 GND.n5105 GND.n2390 19.3944
R12108 GND.n5105 GND.n5104 19.3944
R12109 GND.n5104 GND.n5103 19.3944
R12110 GND.n5103 GND.n2395 19.3944
R12111 GND.n5099 GND.n2395 19.3944
R12112 GND.n5099 GND.n5098 19.3944
R12113 GND.n5098 GND.n5097 19.3944
R12114 GND.n5097 GND.n2400 19.3944
R12115 GND.n5093 GND.n2400 19.3944
R12116 GND.n5093 GND.n5092 19.3944
R12117 GND.n5092 GND.n5091 19.3944
R12118 GND.n5091 GND.n2405 19.3944
R12119 GND.n5087 GND.n2405 19.3944
R12120 GND.n5087 GND.n5086 19.3944
R12121 GND.n5086 GND.n5085 19.3944
R12122 GND.n5085 GND.n2410 19.3944
R12123 GND.n5081 GND.n2410 19.3944
R12124 GND.n5081 GND.n5080 19.3944
R12125 GND.n5080 GND.n5079 19.3944
R12126 GND.n5079 GND.n2415 19.3944
R12127 GND.n5075 GND.n2415 19.3944
R12128 GND.n5075 GND.n5074 19.3944
R12129 GND.n5074 GND.n5073 19.3944
R12130 GND.n5073 GND.n2420 19.3944
R12131 GND.n5069 GND.n2420 19.3944
R12132 GND.n5069 GND.n5068 19.3944
R12133 GND.n5068 GND.n5067 19.3944
R12134 GND.n5067 GND.n2425 19.3944
R12135 GND.n5063 GND.n2425 19.3944
R12136 GND.n5063 GND.n5062 19.3944
R12137 GND.n5062 GND.n5061 19.3944
R12138 GND.n5061 GND.n2430 19.3944
R12139 GND.n5057 GND.n2430 19.3944
R12140 GND.n5057 GND.n5056 19.3944
R12141 GND.n5056 GND.n5055 19.3944
R12142 GND.n5055 GND.n2435 19.3944
R12143 GND.n5051 GND.n2435 19.3944
R12144 GND.n5051 GND.n5050 19.3944
R12145 GND.n5050 GND.n5049 19.3944
R12146 GND.n5049 GND.n2440 19.3944
R12147 GND.n5045 GND.n2440 19.3944
R12148 GND.n5045 GND.n5044 19.3944
R12149 GND.n5044 GND.n5043 19.3944
R12150 GND.n5043 GND.n2445 19.3944
R12151 GND.n5039 GND.n2445 19.3944
R12152 GND.n5039 GND.n5038 19.3944
R12153 GND.n5038 GND.n5037 19.3944
R12154 GND.n5037 GND.n2450 19.3944
R12155 GND.n5033 GND.n2450 19.3944
R12156 GND.n5033 GND.n5032 19.3944
R12157 GND.n5032 GND.n5031 19.3944
R12158 GND.n5031 GND.n2455 19.3944
R12159 GND.n5027 GND.n2455 19.3944
R12160 GND.n5027 GND.n5026 19.3944
R12161 GND.n5026 GND.n5025 19.3944
R12162 GND.n5025 GND.n2460 19.3944
R12163 GND.n5021 GND.n2460 19.3944
R12164 GND.n5021 GND.n5020 19.3944
R12165 GND.n5020 GND.n5019 19.3944
R12166 GND.n5019 GND.n2465 19.3944
R12167 GND.n5015 GND.n2465 19.3944
R12168 GND.n5015 GND.n5014 19.3944
R12169 GND.n5014 GND.n5013 19.3944
R12170 GND.n5013 GND.n2470 19.3944
R12171 GND.n5009 GND.n2470 19.3944
R12172 GND.n5009 GND.n5008 19.3944
R12173 GND.n5008 GND.n5007 19.3944
R12174 GND.n5007 GND.n2475 19.3944
R12175 GND.n5003 GND.n2475 19.3944
R12176 GND.n5003 GND.n5002 19.3944
R12177 GND.n5002 GND.n5001 19.3944
R12178 GND.n5001 GND.n2480 19.3944
R12179 GND.n4997 GND.n2480 19.3944
R12180 GND.n4997 GND.n4996 19.3944
R12181 GND.n4996 GND.n4995 19.3944
R12182 GND.n4995 GND.n2485 19.3944
R12183 GND.n4991 GND.n2485 19.3944
R12184 GND.n4991 GND.n4990 19.3944
R12185 GND.n4990 GND.n4989 19.3944
R12186 GND.n4989 GND.n2490 19.3944
R12187 GND.n4985 GND.n2490 19.3944
R12188 GND.n4985 GND.n4984 19.3944
R12189 GND.n4977 GND.n4976 19.3944
R12190 GND.n4976 GND.n4975 19.3944
R12191 GND.n4975 GND.n2504 19.3944
R12192 GND.n4971 GND.n2504 19.3944
R12193 GND.n4971 GND.n4970 19.3944
R12194 GND.n4970 GND.n4969 19.3944
R12195 GND.n4969 GND.n2509 19.3944
R12196 GND.n4965 GND.n2509 19.3944
R12197 GND.n4965 GND.n4964 19.3944
R12198 GND.n4964 GND.n4963 19.3944
R12199 GND.n4963 GND.n2514 19.3944
R12200 GND.n2935 GND.n2514 19.3944
R12201 GND.n2935 GND.n2928 19.3944
R12202 GND.n2946 GND.n2928 19.3944
R12203 GND.n2946 GND.n2914 19.3944
R12204 GND.n4526 GND.n2903 19.3944
R12205 GND.n4527 GND.n4526 19.3944
R12206 GND.n1939 GND.n1297 19.3944
R12207 GND.n5369 GND.n1297 19.3944
R12208 GND.n5369 GND.n5368 19.3944
R12209 GND.n5368 GND.n5367 19.3944
R12210 GND.n5367 GND.n1300 19.3944
R12211 GND.n5363 GND.n1300 19.3944
R12212 GND.n5363 GND.n5362 19.3944
R12213 GND.n5362 GND.n5361 19.3944
R12214 GND.n5361 GND.n1308 19.3944
R12215 GND.n5357 GND.n1308 19.3944
R12216 GND.n5357 GND.n5356 19.3944
R12217 GND.n5356 GND.n5355 19.3944
R12218 GND.n5355 GND.n1316 19.3944
R12219 GND.n5351 GND.n1316 19.3944
R12220 GND.n5351 GND.n5350 19.3944
R12221 GND.n5350 GND.n5349 19.3944
R12222 GND.n5349 GND.n1324 19.3944
R12223 GND.n5345 GND.n1324 19.3944
R12224 GND.n5345 GND.n5344 19.3944
R12225 GND.n5344 GND.n5343 19.3944
R12226 GND.n5343 GND.n1332 19.3944
R12227 GND.n5339 GND.n1332 19.3944
R12228 GND.n5339 GND.n5338 19.3944
R12229 GND.n5338 GND.n5337 19.3944
R12230 GND.n5337 GND.n1340 19.3944
R12231 GND.n5333 GND.n1340 19.3944
R12232 GND.n5333 GND.n5332 19.3944
R12233 GND.n5332 GND.n5331 19.3944
R12234 GND.n5331 GND.n1348 19.3944
R12235 GND.n5327 GND.n1348 19.3944
R12236 GND.n5327 GND.n5326 19.3944
R12237 GND.n5326 GND.n5325 19.3944
R12238 GND.n5325 GND.n1356 19.3944
R12239 GND.n5321 GND.n1356 19.3944
R12240 GND.n5321 GND.n5320 19.3944
R12241 GND.n5320 GND.n5319 19.3944
R12242 GND.n5319 GND.n1364 19.3944
R12243 GND.n5315 GND.n1364 19.3944
R12244 GND.n5315 GND.n5314 19.3944
R12245 GND.n5314 GND.n5313 19.3944
R12246 GND.n5313 GND.n1372 19.3944
R12247 GND.n5309 GND.n1372 19.3944
R12248 GND.n5309 GND.n5308 19.3944
R12249 GND.n5308 GND.n5307 19.3944
R12250 GND.n5307 GND.n1380 19.3944
R12251 GND.n5303 GND.n1380 19.3944
R12252 GND.n5303 GND.n5302 19.3944
R12253 GND.n5302 GND.n5301 19.3944
R12254 GND.n5301 GND.n1388 19.3944
R12255 GND.n5297 GND.n1388 19.3944
R12256 GND.n5297 GND.n5296 19.3944
R12257 GND.n5289 GND.n5288 19.3944
R12258 GND.n5288 GND.n5287 19.3944
R12259 GND.n5287 GND.n1407 19.3944
R12260 GND.n5283 GND.n1407 19.3944
R12261 GND.n5283 GND.n5282 19.3944
R12262 GND.n5282 GND.n5281 19.3944
R12263 GND.n5277 GND.n5276 19.3944
R12264 GND.n5276 GND.n5275 19.3944
R12265 GND.n5275 GND.n1419 19.3944
R12266 GND.n5271 GND.n1419 19.3944
R12267 GND.n5271 GND.n5270 19.3944
R12268 GND.n5270 GND.n5269 19.3944
R12269 GND.n5269 GND.n1424 19.3944
R12270 GND.n5264 GND.n5263 19.3944
R12271 GND.n5263 GND.n1431 19.3944
R12272 GND.n5258 GND.n5257 19.3944
R12273 GND.n5257 GND.n5256 19.3944
R12274 GND.n5256 GND.n1437 19.3944
R12275 GND.n5252 GND.n5251 19.3944
R12276 GND.n5251 GND.n5250 19.3944
R12277 GND.n5250 GND.n1445 19.3944
R12278 GND.n5246 GND.n1445 19.3944
R12279 GND.n5246 GND.n5245 19.3944
R12280 GND.n5245 GND.n5244 19.3944
R12281 GND.n5244 GND.n1450 19.3944
R12282 GND.n5240 GND.n1450 19.3944
R12283 GND.n5238 GND.n1457 19.3944
R12284 GND.n5234 GND.n1457 19.3944
R12285 GND.n5234 GND.n5233 19.3944
R12286 GND.n5233 GND.n5232 19.3944
R12287 GND.n5232 GND.n1462 19.3944
R12288 GND.n5228 GND.n1462 19.3944
R12289 GND.n5228 GND.n5227 19.3944
R12290 GND.n4960 GND.n2517 19.3944
R12291 GND.n2939 GND.n2517 19.3944
R12292 GND.n2940 GND.n2939 19.3944
R12293 GND.n2943 GND.n2940 19.3944
R12294 GND.n2943 GND.n2910 19.3944
R12295 GND.n4522 GND.n2910 19.3944
R12296 GND.n1965 GND.n1757 19.3944
R12297 GND.n1969 GND.n1757 19.3944
R12298 GND.n1970 GND.n1969 19.3944
R12299 GND.n2014 GND.n1970 19.3944
R12300 GND.n2014 GND.n1751 19.3944
R12301 GND.n2019 GND.n1751 19.3944
R12302 GND.n2019 GND.n1752 19.3944
R12303 GND.n1752 GND.n1732 19.3944
R12304 GND.n2039 GND.n1732 19.3944
R12305 GND.n2039 GND.n1729 19.3944
R12306 GND.n2044 GND.n1729 19.3944
R12307 GND.n2044 GND.n1730 19.3944
R12308 GND.n1730 GND.n1704 19.3944
R12309 GND.n2092 GND.n1704 19.3944
R12310 GND.n2092 GND.n1701 19.3944
R12311 GND.n2097 GND.n1701 19.3944
R12312 GND.n2097 GND.n1702 19.3944
R12313 GND.n1702 GND.n1680 19.3944
R12314 GND.n2114 GND.n1680 19.3944
R12315 GND.n2114 GND.n1678 19.3944
R12316 GND.n2118 GND.n1678 19.3944
R12317 GND.n2119 GND.n2118 19.3944
R12318 GND.n2122 GND.n2119 19.3944
R12319 GND.n2122 GND.n1676 19.3944
R12320 GND.n2126 GND.n1676 19.3944
R12321 GND.n2127 GND.n2126 19.3944
R12322 GND.n2127 GND.n1674 19.3944
R12323 GND.n2131 GND.n1674 19.3944
R12324 GND.n2131 GND.n1625 19.3944
R12325 GND.n2222 GND.n1625 19.3944
R12326 GND.n2222 GND.n1622 19.3944
R12327 GND.n2227 GND.n1622 19.3944
R12328 GND.n2227 GND.n1623 19.3944
R12329 GND.n1623 GND.n1601 19.3944
R12330 GND.n2246 GND.n1601 19.3944
R12331 GND.n2246 GND.n1598 19.3944
R12332 GND.n2251 GND.n1598 19.3944
R12333 GND.n2251 GND.n1599 19.3944
R12334 GND.n1599 GND.n1578 19.3944
R12335 GND.n2271 GND.n1578 19.3944
R12336 GND.n2271 GND.n1575 19.3944
R12337 GND.n2290 GND.n1575 19.3944
R12338 GND.n2290 GND.n1576 19.3944
R12339 GND.n2286 GND.n1576 19.3944
R12340 GND.n2286 GND.n2285 19.3944
R12341 GND.n2285 GND.n2284 19.3944
R12342 GND.n2284 GND.n2276 19.3944
R12343 GND.n2280 GND.n2276 19.3944
R12344 GND.n2280 GND.n1539 19.3944
R12345 GND.n2347 GND.n1539 19.3944
R12346 GND.n2348 GND.n2347 19.3944
R12347 GND.n5216 GND.n1477 19.3944
R12348 GND.n5216 GND.n5215 19.3944
R12349 GND.n5215 GND.n1480 19.3944
R12350 GND.n5208 GND.n1480 19.3944
R12351 GND.n5208 GND.n5207 19.3944
R12352 GND.n5207 GND.n1488 19.3944
R12353 GND.n1944 GND.n1767 19.3944
R12354 GND.n1948 GND.n1767 19.3944
R12355 GND.n1948 GND.n1765 19.3944
R12356 GND.n1954 GND.n1765 19.3944
R12357 GND.n1954 GND.n1763 19.3944
R12358 GND.n1958 GND.n1763 19.3944
R12359 GND.n1938 GND.n1293 19.3944
R12360 GND.n5371 GND.n1293 19.3944
R12361 GND.n5371 GND.n1294 19.3944
R12362 GND.n1301 GND.n1294 19.3944
R12363 GND.n1302 GND.n1301 19.3944
R12364 GND.n1303 GND.n1302 19.3944
R12365 GND.n2025 GND.n1303 19.3944
R12366 GND.n2025 GND.n1309 19.3944
R12367 GND.n1310 GND.n1309 19.3944
R12368 GND.n1311 GND.n1310 19.3944
R12369 GND.n1718 GND.n1311 19.3944
R12370 GND.n1718 GND.n1317 19.3944
R12371 GND.n1318 GND.n1317 19.3944
R12372 GND.n1319 GND.n1318 19.3944
R12373 GND.n1697 GND.n1319 19.3944
R12374 GND.n1697 GND.n1325 19.3944
R12375 GND.n1326 GND.n1325 19.3944
R12376 GND.n1327 GND.n1326 19.3944
R12377 GND.n1686 GND.n1327 19.3944
R12378 GND.n1686 GND.n1333 19.3944
R12379 GND.n1334 GND.n1333 19.3944
R12380 GND.n1335 GND.n1334 19.3944
R12381 GND.n1649 GND.n1335 19.3944
R12382 GND.n1649 GND.n1341 19.3944
R12383 GND.n1342 GND.n1341 19.3944
R12384 GND.n1343 GND.n1342 19.3944
R12385 GND.n1672 GND.n1343 19.3944
R12386 GND.n1672 GND.n1349 19.3944
R12387 GND.n1350 GND.n1349 19.3944
R12388 GND.n1351 GND.n1350 19.3944
R12389 GND.n1618 GND.n1351 19.3944
R12390 GND.n1618 GND.n1357 19.3944
R12391 GND.n1358 GND.n1357 19.3944
R12392 GND.n1359 GND.n1358 19.3944
R12393 GND.n1605 GND.n1359 19.3944
R12394 GND.n1605 GND.n1365 19.3944
R12395 GND.n1366 GND.n1365 19.3944
R12396 GND.n1367 GND.n1366 19.3944
R12397 GND.n2255 GND.n1367 19.3944
R12398 GND.n2255 GND.n1373 19.3944
R12399 GND.n1374 GND.n1373 19.3944
R12400 GND.n1375 GND.n1374 19.3944
R12401 GND.n2295 GND.n1375 19.3944
R12402 GND.n2295 GND.n1381 19.3944
R12403 GND.n1382 GND.n1381 19.3944
R12404 GND.n1383 GND.n1382 19.3944
R12405 GND.n2332 GND.n1383 19.3944
R12406 GND.n2332 GND.n1389 19.3944
R12407 GND.n1390 GND.n1389 19.3944
R12408 GND.n1391 GND.n1390 19.3944
R12409 GND.n1398 GND.n1391 19.3944
R12410 GND.n6191 GND.n735 19.3944
R12411 GND.n6191 GND.n733 19.3944
R12412 GND.n6195 GND.n733 19.3944
R12413 GND.n6195 GND.n729 19.3944
R12414 GND.n6201 GND.n729 19.3944
R12415 GND.n6201 GND.n727 19.3944
R12416 GND.n6205 GND.n727 19.3944
R12417 GND.n6205 GND.n723 19.3944
R12418 GND.n6211 GND.n723 19.3944
R12419 GND.n6211 GND.n721 19.3944
R12420 GND.n6215 GND.n721 19.3944
R12421 GND.n6215 GND.n717 19.3944
R12422 GND.n6221 GND.n717 19.3944
R12423 GND.n6221 GND.n715 19.3944
R12424 GND.n6225 GND.n715 19.3944
R12425 GND.n6225 GND.n711 19.3944
R12426 GND.n6231 GND.n711 19.3944
R12427 GND.n6231 GND.n709 19.3944
R12428 GND.n6235 GND.n709 19.3944
R12429 GND.n6235 GND.n705 19.3944
R12430 GND.n6241 GND.n705 19.3944
R12431 GND.n6241 GND.n703 19.3944
R12432 GND.n6245 GND.n703 19.3944
R12433 GND.n6245 GND.n699 19.3944
R12434 GND.n6251 GND.n699 19.3944
R12435 GND.n6251 GND.n697 19.3944
R12436 GND.n6255 GND.n697 19.3944
R12437 GND.n6255 GND.n693 19.3944
R12438 GND.n6261 GND.n693 19.3944
R12439 GND.n6261 GND.n691 19.3944
R12440 GND.n6265 GND.n691 19.3944
R12441 GND.n6265 GND.n687 19.3944
R12442 GND.n6271 GND.n687 19.3944
R12443 GND.n6271 GND.n685 19.3944
R12444 GND.n6275 GND.n685 19.3944
R12445 GND.n6275 GND.n681 19.3944
R12446 GND.n6281 GND.n681 19.3944
R12447 GND.n6281 GND.n679 19.3944
R12448 GND.n6285 GND.n679 19.3944
R12449 GND.n6285 GND.n675 19.3944
R12450 GND.n6291 GND.n675 19.3944
R12451 GND.n6291 GND.n673 19.3944
R12452 GND.n6295 GND.n673 19.3944
R12453 GND.n6295 GND.n669 19.3944
R12454 GND.n6301 GND.n669 19.3944
R12455 GND.n6301 GND.n667 19.3944
R12456 GND.n6307 GND.n667 19.3944
R12457 GND.n6307 GND.n6306 19.3944
R12458 GND.n5521 GND.n1137 19.3944
R12459 GND.n5521 GND.n1135 19.3944
R12460 GND.n5525 GND.n1135 19.3944
R12461 GND.n5525 GND.n1131 19.3944
R12462 GND.n5531 GND.n1131 19.3944
R12463 GND.n5531 GND.n1129 19.3944
R12464 GND.n5535 GND.n1129 19.3944
R12465 GND.n5535 GND.n1125 19.3944
R12466 GND.n5541 GND.n1125 19.3944
R12467 GND.n5541 GND.n1123 19.3944
R12468 GND.n5545 GND.n1123 19.3944
R12469 GND.n5545 GND.n1119 19.3944
R12470 GND.n5551 GND.n1119 19.3944
R12471 GND.n5551 GND.n1117 19.3944
R12472 GND.n5555 GND.n1117 19.3944
R12473 GND.n5555 GND.n1113 19.3944
R12474 GND.n5561 GND.n1113 19.3944
R12475 GND.n5561 GND.n1111 19.3944
R12476 GND.n5565 GND.n1111 19.3944
R12477 GND.n5565 GND.n1107 19.3944
R12478 GND.n5571 GND.n1107 19.3944
R12479 GND.n5571 GND.n1105 19.3944
R12480 GND.n5575 GND.n1105 19.3944
R12481 GND.n5575 GND.n1101 19.3944
R12482 GND.n5581 GND.n1101 19.3944
R12483 GND.n5581 GND.n1099 19.3944
R12484 GND.n5585 GND.n1099 19.3944
R12485 GND.n5585 GND.n1095 19.3944
R12486 GND.n5591 GND.n1095 19.3944
R12487 GND.n5591 GND.n1093 19.3944
R12488 GND.n5595 GND.n1093 19.3944
R12489 GND.n5595 GND.n1089 19.3944
R12490 GND.n5601 GND.n1089 19.3944
R12491 GND.n5601 GND.n1087 19.3944
R12492 GND.n5605 GND.n1087 19.3944
R12493 GND.n5605 GND.n1083 19.3944
R12494 GND.n5611 GND.n1083 19.3944
R12495 GND.n5611 GND.n1081 19.3944
R12496 GND.n5615 GND.n1081 19.3944
R12497 GND.n5615 GND.n1077 19.3944
R12498 GND.n5621 GND.n1077 19.3944
R12499 GND.n5621 GND.n1075 19.3944
R12500 GND.n5625 GND.n1075 19.3944
R12501 GND.n5625 GND.n1071 19.3944
R12502 GND.n5631 GND.n1071 19.3944
R12503 GND.n5631 GND.n1069 19.3944
R12504 GND.n5635 GND.n1069 19.3944
R12505 GND.n5635 GND.n1065 19.3944
R12506 GND.n5641 GND.n1065 19.3944
R12507 GND.n5641 GND.n1063 19.3944
R12508 GND.n5645 GND.n1063 19.3944
R12509 GND.n5645 GND.n1059 19.3944
R12510 GND.n5651 GND.n1059 19.3944
R12511 GND.n5651 GND.n1057 19.3944
R12512 GND.n5655 GND.n1057 19.3944
R12513 GND.n5655 GND.n1053 19.3944
R12514 GND.n5661 GND.n1053 19.3944
R12515 GND.n5661 GND.n1051 19.3944
R12516 GND.n5665 GND.n1051 19.3944
R12517 GND.n5665 GND.n1047 19.3944
R12518 GND.n5671 GND.n1047 19.3944
R12519 GND.n5671 GND.n1045 19.3944
R12520 GND.n5675 GND.n1045 19.3944
R12521 GND.n5675 GND.n1041 19.3944
R12522 GND.n5681 GND.n1041 19.3944
R12523 GND.n5681 GND.n1039 19.3944
R12524 GND.n5685 GND.n1039 19.3944
R12525 GND.n5685 GND.n1035 19.3944
R12526 GND.n5691 GND.n1035 19.3944
R12527 GND.n5691 GND.n1033 19.3944
R12528 GND.n5695 GND.n1033 19.3944
R12529 GND.n5695 GND.n1029 19.3944
R12530 GND.n5701 GND.n1029 19.3944
R12531 GND.n5701 GND.n1027 19.3944
R12532 GND.n5705 GND.n1027 19.3944
R12533 GND.n5705 GND.n1023 19.3944
R12534 GND.n5711 GND.n1023 19.3944
R12535 GND.n5711 GND.n1021 19.3944
R12536 GND.n5715 GND.n1021 19.3944
R12537 GND.n5715 GND.n1017 19.3944
R12538 GND.n5721 GND.n1017 19.3944
R12539 GND.n5721 GND.n1015 19.3944
R12540 GND.n5725 GND.n1015 19.3944
R12541 GND.n5725 GND.n1011 19.3944
R12542 GND.n5731 GND.n1011 19.3944
R12543 GND.n5731 GND.n1009 19.3944
R12544 GND.n5735 GND.n1009 19.3944
R12545 GND.n5735 GND.n1005 19.3944
R12546 GND.n5741 GND.n1005 19.3944
R12547 GND.n5741 GND.n1003 19.3944
R12548 GND.n5745 GND.n1003 19.3944
R12549 GND.n5745 GND.n999 19.3944
R12550 GND.n5751 GND.n999 19.3944
R12551 GND.n5751 GND.n997 19.3944
R12552 GND.n5755 GND.n997 19.3944
R12553 GND.n5755 GND.n993 19.3944
R12554 GND.n5761 GND.n993 19.3944
R12555 GND.n5761 GND.n991 19.3944
R12556 GND.n5765 GND.n991 19.3944
R12557 GND.n5765 GND.n987 19.3944
R12558 GND.n5771 GND.n987 19.3944
R12559 GND.n5771 GND.n985 19.3944
R12560 GND.n5775 GND.n985 19.3944
R12561 GND.n5775 GND.n981 19.3944
R12562 GND.n5781 GND.n981 19.3944
R12563 GND.n5781 GND.n979 19.3944
R12564 GND.n5785 GND.n979 19.3944
R12565 GND.n5785 GND.n975 19.3944
R12566 GND.n5791 GND.n975 19.3944
R12567 GND.n5791 GND.n973 19.3944
R12568 GND.n5795 GND.n973 19.3944
R12569 GND.n5795 GND.n969 19.3944
R12570 GND.n5801 GND.n969 19.3944
R12571 GND.n5801 GND.n967 19.3944
R12572 GND.n5805 GND.n967 19.3944
R12573 GND.n5805 GND.n963 19.3944
R12574 GND.n5811 GND.n963 19.3944
R12575 GND.n5811 GND.n961 19.3944
R12576 GND.n5815 GND.n961 19.3944
R12577 GND.n5815 GND.n957 19.3944
R12578 GND.n5821 GND.n957 19.3944
R12579 GND.n5821 GND.n955 19.3944
R12580 GND.n5825 GND.n955 19.3944
R12581 GND.n5825 GND.n951 19.3944
R12582 GND.n5831 GND.n951 19.3944
R12583 GND.n5831 GND.n949 19.3944
R12584 GND.n5835 GND.n949 19.3944
R12585 GND.n5835 GND.n945 19.3944
R12586 GND.n5841 GND.n945 19.3944
R12587 GND.n5841 GND.n943 19.3944
R12588 GND.n5845 GND.n943 19.3944
R12589 GND.n5845 GND.n939 19.3944
R12590 GND.n5851 GND.n939 19.3944
R12591 GND.n5851 GND.n937 19.3944
R12592 GND.n5855 GND.n937 19.3944
R12593 GND.n5855 GND.n933 19.3944
R12594 GND.n5861 GND.n933 19.3944
R12595 GND.n5861 GND.n931 19.3944
R12596 GND.n5865 GND.n931 19.3944
R12597 GND.n5865 GND.n927 19.3944
R12598 GND.n5871 GND.n927 19.3944
R12599 GND.n5871 GND.n925 19.3944
R12600 GND.n5875 GND.n925 19.3944
R12601 GND.n5875 GND.n921 19.3944
R12602 GND.n5881 GND.n921 19.3944
R12603 GND.n5881 GND.n919 19.3944
R12604 GND.n5885 GND.n919 19.3944
R12605 GND.n5885 GND.n915 19.3944
R12606 GND.n5891 GND.n915 19.3944
R12607 GND.n5891 GND.n913 19.3944
R12608 GND.n5895 GND.n913 19.3944
R12609 GND.n5895 GND.n909 19.3944
R12610 GND.n5901 GND.n909 19.3944
R12611 GND.n5901 GND.n907 19.3944
R12612 GND.n5905 GND.n907 19.3944
R12613 GND.n5905 GND.n903 19.3944
R12614 GND.n5911 GND.n903 19.3944
R12615 GND.n5911 GND.n901 19.3944
R12616 GND.n5915 GND.n901 19.3944
R12617 GND.n5915 GND.n897 19.3944
R12618 GND.n5921 GND.n897 19.3944
R12619 GND.n5921 GND.n895 19.3944
R12620 GND.n5925 GND.n895 19.3944
R12621 GND.n5925 GND.n891 19.3944
R12622 GND.n5931 GND.n891 19.3944
R12623 GND.n5931 GND.n889 19.3944
R12624 GND.n5935 GND.n889 19.3944
R12625 GND.n5935 GND.n885 19.3944
R12626 GND.n5941 GND.n885 19.3944
R12627 GND.n5941 GND.n883 19.3944
R12628 GND.n5945 GND.n883 19.3944
R12629 GND.n5945 GND.n879 19.3944
R12630 GND.n5951 GND.n879 19.3944
R12631 GND.n5951 GND.n877 19.3944
R12632 GND.n5955 GND.n877 19.3944
R12633 GND.n5955 GND.n873 19.3944
R12634 GND.n5961 GND.n873 19.3944
R12635 GND.n5961 GND.n871 19.3944
R12636 GND.n5965 GND.n871 19.3944
R12637 GND.n5965 GND.n867 19.3944
R12638 GND.n5971 GND.n867 19.3944
R12639 GND.n5971 GND.n865 19.3944
R12640 GND.n5975 GND.n865 19.3944
R12641 GND.n5975 GND.n861 19.3944
R12642 GND.n5981 GND.n861 19.3944
R12643 GND.n5981 GND.n859 19.3944
R12644 GND.n5985 GND.n859 19.3944
R12645 GND.n5985 GND.n855 19.3944
R12646 GND.n5991 GND.n855 19.3944
R12647 GND.n5991 GND.n853 19.3944
R12648 GND.n5995 GND.n853 19.3944
R12649 GND.n5995 GND.n849 19.3944
R12650 GND.n6001 GND.n849 19.3944
R12651 GND.n6001 GND.n847 19.3944
R12652 GND.n6005 GND.n847 19.3944
R12653 GND.n6005 GND.n843 19.3944
R12654 GND.n6011 GND.n843 19.3944
R12655 GND.n6011 GND.n841 19.3944
R12656 GND.n6015 GND.n841 19.3944
R12657 GND.n6015 GND.n837 19.3944
R12658 GND.n6021 GND.n837 19.3944
R12659 GND.n6021 GND.n835 19.3944
R12660 GND.n6025 GND.n835 19.3944
R12661 GND.n6025 GND.n831 19.3944
R12662 GND.n6031 GND.n831 19.3944
R12663 GND.n6031 GND.n829 19.3944
R12664 GND.n6035 GND.n829 19.3944
R12665 GND.n6035 GND.n825 19.3944
R12666 GND.n6041 GND.n825 19.3944
R12667 GND.n6041 GND.n823 19.3944
R12668 GND.n6045 GND.n823 19.3944
R12669 GND.n6045 GND.n819 19.3944
R12670 GND.n6051 GND.n819 19.3944
R12671 GND.n6051 GND.n817 19.3944
R12672 GND.n6055 GND.n817 19.3944
R12673 GND.n6055 GND.n813 19.3944
R12674 GND.n6061 GND.n813 19.3944
R12675 GND.n6061 GND.n811 19.3944
R12676 GND.n6065 GND.n811 19.3944
R12677 GND.n6065 GND.n807 19.3944
R12678 GND.n6071 GND.n807 19.3944
R12679 GND.n6071 GND.n805 19.3944
R12680 GND.n6075 GND.n805 19.3944
R12681 GND.n6075 GND.n801 19.3944
R12682 GND.n6081 GND.n801 19.3944
R12683 GND.n6081 GND.n799 19.3944
R12684 GND.n6085 GND.n799 19.3944
R12685 GND.n6085 GND.n795 19.3944
R12686 GND.n6091 GND.n795 19.3944
R12687 GND.n6091 GND.n793 19.3944
R12688 GND.n6095 GND.n793 19.3944
R12689 GND.n6095 GND.n789 19.3944
R12690 GND.n6101 GND.n789 19.3944
R12691 GND.n6101 GND.n787 19.3944
R12692 GND.n6105 GND.n787 19.3944
R12693 GND.n6105 GND.n783 19.3944
R12694 GND.n6111 GND.n783 19.3944
R12695 GND.n6111 GND.n781 19.3944
R12696 GND.n6115 GND.n781 19.3944
R12697 GND.n6115 GND.n777 19.3944
R12698 GND.n6121 GND.n777 19.3944
R12699 GND.n6121 GND.n775 19.3944
R12700 GND.n6125 GND.n775 19.3944
R12701 GND.n6125 GND.n771 19.3944
R12702 GND.n6131 GND.n771 19.3944
R12703 GND.n6131 GND.n769 19.3944
R12704 GND.n6135 GND.n769 19.3944
R12705 GND.n6135 GND.n765 19.3944
R12706 GND.n6141 GND.n765 19.3944
R12707 GND.n6141 GND.n763 19.3944
R12708 GND.n6145 GND.n763 19.3944
R12709 GND.n6145 GND.n759 19.3944
R12710 GND.n6151 GND.n759 19.3944
R12711 GND.n6151 GND.n757 19.3944
R12712 GND.n6155 GND.n757 19.3944
R12713 GND.n6155 GND.n753 19.3944
R12714 GND.n6161 GND.n753 19.3944
R12715 GND.n6161 GND.n751 19.3944
R12716 GND.n6165 GND.n751 19.3944
R12717 GND.n6165 GND.n747 19.3944
R12718 GND.n6171 GND.n747 19.3944
R12719 GND.n6171 GND.n745 19.3944
R12720 GND.n6175 GND.n745 19.3944
R12721 GND.n6175 GND.n741 19.3944
R12722 GND.n6181 GND.n741 19.3944
R12723 GND.n6181 GND.n739 19.3944
R12724 GND.n6185 GND.n739 19.3944
R12725 GND.n4954 GND.n4953 19.3944
R12726 GND.n4953 GND.n4952 19.3944
R12727 GND.n4952 GND.n4951 19.3944
R12728 GND.n4951 GND.n4949 19.3944
R12729 GND.n4949 GND.n4946 19.3944
R12730 GND.n4946 GND.n4945 19.3944
R12731 GND.n4941 GND.n4938 19.3944
R12732 GND.n4938 GND.n4937 19.3944
R12733 GND.n4937 GND.n4934 19.3944
R12734 GND.n4934 GND.n4933 19.3944
R12735 GND.n4933 GND.n4930 19.3944
R12736 GND.n4930 GND.n4929 19.3944
R12737 GND.n4929 GND.n4926 19.3944
R12738 GND.n4924 GND.n4922 19.3944
R12739 GND.n4922 GND.n4919 19.3944
R12740 GND.n4917 GND.n4914 19.3944
R12741 GND.n4914 GND.n4913 19.3944
R12742 GND.n4913 GND.n4910 19.3944
R12743 GND.n4908 GND.n4905 19.3944
R12744 GND.n4905 GND.n4904 19.3944
R12745 GND.n4904 GND.n4901 19.3944
R12746 GND.n4901 GND.n4900 19.3944
R12747 GND.n4900 GND.n4897 19.3944
R12748 GND.n4897 GND.n4896 19.3944
R12749 GND.n4896 GND.n4893 19.3944
R12750 GND.n4893 GND.n4892 19.3944
R12751 GND.n4888 GND.n4885 19.3944
R12752 GND.n4885 GND.n4884 19.3944
R12753 GND.n4884 GND.n4881 19.3944
R12754 GND.n4881 GND.n4880 19.3944
R12755 GND.n4880 GND.n4877 19.3944
R12756 GND.n4877 GND.n4876 19.3944
R12757 GND.n4876 GND.n4873 19.3944
R12758 GND.n4866 GND.n2610 19.3944
R12759 GND.n4540 GND.n2610 19.3944
R12760 GND.n4540 GND.n4538 19.3944
R12761 GND.n4549 GND.n4538 19.3944
R12762 GND.n4549 GND.n2898 19.3944
R12763 GND.n4561 GND.n2898 19.3944
R12764 GND.n4562 GND.n4561 19.3944
R12765 GND.n4564 GND.n4562 19.3944
R12766 GND.n4564 GND.n2894 19.3944
R12767 GND.n4576 GND.n2894 19.3944
R12768 GND.n4577 GND.n4576 19.3944
R12769 GND.n4579 GND.n4577 19.3944
R12770 GND.n4579 GND.n2890 19.3944
R12771 GND.n4591 GND.n2890 19.3944
R12772 GND.n4592 GND.n4591 19.3944
R12773 GND.n4594 GND.n4592 19.3944
R12774 GND.n4594 GND.n2886 19.3944
R12775 GND.n4606 GND.n2886 19.3944
R12776 GND.n4607 GND.n4606 19.3944
R12777 GND.n4609 GND.n4607 19.3944
R12778 GND.n4609 GND.n2882 19.3944
R12779 GND.n4625 GND.n2882 19.3944
R12780 GND.n4626 GND.n4625 19.3944
R12781 GND.n4627 GND.n4626 19.3944
R12782 GND.n4627 GND.n2881 19.3944
R12783 GND.n4634 GND.n2881 19.3944
R12784 GND.n4636 GND.n4634 19.3944
R12785 GND.n4777 GND.n4636 19.3944
R12786 GND.n4777 GND.n4776 19.3944
R12787 GND.n4776 GND.n4637 19.3944
R12788 GND.n4766 GND.n4637 19.3944
R12789 GND.n4766 GND.n4765 19.3944
R12790 GND.n4765 GND.n4764 19.3944
R12791 GND.n4764 GND.n4645 19.3944
R12792 GND.n4754 GND.n4645 19.3944
R12793 GND.n4754 GND.n4753 19.3944
R12794 GND.n4753 GND.n4752 19.3944
R12795 GND.n4752 GND.n4652 19.3944
R12796 GND.n4742 GND.n4652 19.3944
R12797 GND.n4742 GND.n4741 19.3944
R12798 GND.n4741 GND.n4740 19.3944
R12799 GND.n4740 GND.n4659 19.3944
R12800 GND.n4730 GND.n4659 19.3944
R12801 GND.n4730 GND.n4729 19.3944
R12802 GND.n4729 GND.n4728 19.3944
R12803 GND.n4728 GND.n4666 19.3944
R12804 GND.n4718 GND.n4666 19.3944
R12805 GND.n4718 GND.n4717 19.3944
R12806 GND.n4717 GND.n4716 19.3944
R12807 GND.n4716 GND.n449 19.3944
R12808 GND.n6352 GND.n449 19.3944
R12809 GND.n4542 GND.n2608 19.3944
R12810 GND.n4545 GND.n4542 19.3944
R12811 GND.n4546 GND.n4545 19.3944
R12812 GND.n4546 GND.n2649 19.3944
R12813 GND.n4848 GND.n2649 19.3944
R12814 GND.n4848 GND.n4847 19.3944
R12815 GND.n4847 GND.n4846 19.3944
R12816 GND.n4846 GND.n2653 19.3944
R12817 GND.n4836 GND.n2653 19.3944
R12818 GND.n4836 GND.n4835 19.3944
R12819 GND.n4835 GND.n4834 19.3944
R12820 GND.n4834 GND.n2674 19.3944
R12821 GND.n4824 GND.n2674 19.3944
R12822 GND.n4824 GND.n4823 19.3944
R12823 GND.n4823 GND.n4822 19.3944
R12824 GND.n4822 GND.n2695 19.3944
R12825 GND.n4812 GND.n2695 19.3944
R12826 GND.n4812 GND.n4811 19.3944
R12827 GND.n4811 GND.n4810 19.3944
R12828 GND.n4810 GND.n2716 19.3944
R12829 GND.n4800 GND.n2716 19.3944
R12830 GND.n4800 GND.n4799 19.3944
R12831 GND.n4799 GND.n4798 19.3944
R12832 GND.n4798 GND.n2735 19.3944
R12833 GND.n4631 GND.n2735 19.3944
R12834 GND.n4632 GND.n4631 19.3944
R12835 GND.n4632 GND.n2877 19.3944
R12836 GND.n4779 GND.n2877 19.3944
R12837 GND.n4779 GND.n342 19.3944
R12838 GND.n6415 GND.n342 19.3944
R12839 GND.n6415 GND.n6414 19.3944
R12840 GND.n6414 GND.n6413 19.3944
R12841 GND.n6413 GND.n346 19.3944
R12842 GND.n6403 GND.n346 19.3944
R12843 GND.n6403 GND.n6402 19.3944
R12844 GND.n6402 GND.n6401 19.3944
R12845 GND.n6401 GND.n366 19.3944
R12846 GND.n6391 GND.n366 19.3944
R12847 GND.n6391 GND.n6390 19.3944
R12848 GND.n6390 GND.n6389 19.3944
R12849 GND.n6389 GND.n387 19.3944
R12850 GND.n6379 GND.n387 19.3944
R12851 GND.n6379 GND.n6378 19.3944
R12852 GND.n6378 GND.n6377 19.3944
R12853 GND.n6377 GND.n408 19.3944
R12854 GND.n6367 GND.n408 19.3944
R12855 GND.n6367 GND.n6366 19.3944
R12856 GND.n6366 GND.n6365 19.3944
R12857 GND.n6365 GND.n429 19.3944
R12858 GND.n6355 GND.n429 19.3944
R12859 GND.n6355 GND.n6354 19.3944
R12860 GND.n615 GND.n612 19.3944
R12861 GND.n615 GND.n491 19.3944
R12862 GND.n619 GND.n491 19.3944
R12863 GND.n622 GND.n619 19.3944
R12864 GND.n625 GND.n622 19.3944
R12865 GND.n625 GND.n489 19.3944
R12866 GND.n629 GND.n489 19.3944
R12867 GND.n589 GND.n588 19.3944
R12868 GND.n592 GND.n589 19.3944
R12869 GND.n592 GND.n498 19.3944
R12870 GND.n598 GND.n498 19.3944
R12871 GND.n599 GND.n598 19.3944
R12872 GND.n602 GND.n599 19.3944
R12873 GND.n602 GND.n496 19.3944
R12874 GND.n608 GND.n496 19.3944
R12875 GND.n568 GND.n565 19.3944
R12876 GND.n571 GND.n568 19.3944
R12877 GND.n571 GND.n506 19.3944
R12878 GND.n575 GND.n506 19.3944
R12879 GND.n578 GND.n575 19.3944
R12880 GND.n581 GND.n578 19.3944
R12881 GND.n581 GND.n504 19.3944
R12882 GND.n585 GND.n504 19.3944
R12883 GND.n545 GND.n514 19.3944
R12884 GND.n548 GND.n545 19.3944
R12885 GND.n551 GND.n548 19.3944
R12886 GND.n551 GND.n512 19.3944
R12887 GND.n555 GND.n512 19.3944
R12888 GND.n558 GND.n555 19.3944
R12889 GND.n561 GND.n558 19.3944
R12890 GND.n527 GND.n523 19.3944
R12891 GND.n530 GND.n527 19.3944
R12892 GND.n533 GND.n530 19.3944
R12893 GND.n533 GND.n520 19.3944
R12894 GND.n537 GND.n520 19.3944
R12895 GND.n540 GND.n537 19.3944
R12896 GND.n4688 GND.n4685 19.3944
R12897 GND.n4692 GND.n4685 19.3944
R12898 GND.n4692 GND.n4683 19.3944
R12899 GND.n4698 GND.n4683 19.3944
R12900 GND.n4698 GND.n4681 19.3944
R12901 GND.n4702 GND.n4681 19.3944
R12902 GND.n4530 GND.n2901 19.3944
R12903 GND.n4536 GND.n2901 19.3944
R12904 GND.n4537 GND.n4536 19.3944
R12905 GND.n4553 GND.n4537 19.3944
R12906 GND.n4553 GND.n2899 19.3944
R12907 GND.n4557 GND.n2899 19.3944
R12908 GND.n4557 GND.n2897 19.3944
R12909 GND.n4568 GND.n2897 19.3944
R12910 GND.n4568 GND.n2895 19.3944
R12911 GND.n4572 GND.n2895 19.3944
R12912 GND.n4572 GND.n2893 19.3944
R12913 GND.n4583 GND.n2893 19.3944
R12914 GND.n4583 GND.n2891 19.3944
R12915 GND.n4587 GND.n2891 19.3944
R12916 GND.n4587 GND.n2889 19.3944
R12917 GND.n4598 GND.n2889 19.3944
R12918 GND.n4598 GND.n2887 19.3944
R12919 GND.n4602 GND.n2887 19.3944
R12920 GND.n4602 GND.n2885 19.3944
R12921 GND.n4613 GND.n2885 19.3944
R12922 GND.n4613 GND.n2883 19.3944
R12923 GND.n4621 GND.n2883 19.3944
R12924 GND.n4621 GND.n4620 19.3944
R12925 GND.n4620 GND.n4619 19.3944
R12926 GND.n4619 GND.n313 19.3944
R12927 GND.n6426 GND.n313 19.3944
R12928 GND.n6426 GND.n314 19.3944
R12929 GND.n4638 GND.n314 19.3944
R12930 GND.n4772 GND.n4638 19.3944
R12931 GND.n4772 GND.n4771 19.3944
R12932 GND.n4771 GND.n4770 19.3944
R12933 GND.n4770 GND.n4643 19.3944
R12934 GND.n4760 GND.n4643 19.3944
R12935 GND.n4760 GND.n4759 19.3944
R12936 GND.n4759 GND.n4758 19.3944
R12937 GND.n4758 GND.n4650 19.3944
R12938 GND.n4748 GND.n4650 19.3944
R12939 GND.n4748 GND.n4747 19.3944
R12940 GND.n4747 GND.n4746 19.3944
R12941 GND.n4746 GND.n4657 19.3944
R12942 GND.n4736 GND.n4657 19.3944
R12943 GND.n4736 GND.n4735 19.3944
R12944 GND.n4735 GND.n4734 19.3944
R12945 GND.n4734 GND.n4664 19.3944
R12946 GND.n4724 GND.n4664 19.3944
R12947 GND.n4724 GND.n4723 19.3944
R12948 GND.n4723 GND.n4722 19.3944
R12949 GND.n4722 GND.n4671 19.3944
R12950 GND.n4712 GND.n4671 19.3944
R12951 GND.n4712 GND.n4711 19.3944
R12952 GND.n4711 GND.n4710 19.3944
R12953 GND.n2635 GND.n2633 19.3944
R12954 GND.n2635 GND.n2631 19.3944
R12955 GND.n4854 GND.n2631 19.3944
R12956 GND.n4854 GND.n4853 19.3944
R12957 GND.n4853 GND.n4852 19.3944
R12958 GND.n4852 GND.n2641 19.3944
R12959 GND.n4842 GND.n2641 19.3944
R12960 GND.n4842 GND.n4841 19.3944
R12961 GND.n4841 GND.n4840 19.3944
R12962 GND.n4840 GND.n2664 19.3944
R12963 GND.n4830 GND.n2664 19.3944
R12964 GND.n4830 GND.n4829 19.3944
R12965 GND.n4829 GND.n4828 19.3944
R12966 GND.n4828 GND.n2685 19.3944
R12967 GND.n4818 GND.n2685 19.3944
R12968 GND.n4818 GND.n4817 19.3944
R12969 GND.n4817 GND.n4816 19.3944
R12970 GND.n4816 GND.n2706 19.3944
R12971 GND.n4806 GND.n2706 19.3944
R12972 GND.n4806 GND.n4805 19.3944
R12973 GND.n4805 GND.n4804 19.3944
R12974 GND.n2725 GND.n330 19.3944
R12975 GND.n2741 GND.n330 19.3944
R12976 GND.n6422 GND.n323 19.3944
R12977 GND.n4781 GND.n324 19.3944
R12978 GND.n6419 GND.n332 19.3944
R12979 GND.n6419 GND.n333 19.3944
R12980 GND.n6409 GND.n333 19.3944
R12981 GND.n6409 GND.n6408 19.3944
R12982 GND.n6408 GND.n6407 19.3944
R12983 GND.n6407 GND.n356 19.3944
R12984 GND.n6397 GND.n356 19.3944
R12985 GND.n6397 GND.n6396 19.3944
R12986 GND.n6396 GND.n6395 19.3944
R12987 GND.n6395 GND.n377 19.3944
R12988 GND.n6385 GND.n377 19.3944
R12989 GND.n6385 GND.n6384 19.3944
R12990 GND.n6384 GND.n6383 19.3944
R12991 GND.n6383 GND.n398 19.3944
R12992 GND.n6373 GND.n398 19.3944
R12993 GND.n6373 GND.n6372 19.3944
R12994 GND.n6372 GND.n6371 19.3944
R12995 GND.n6371 GND.n419 19.3944
R12996 GND.n6361 GND.n419 19.3944
R12997 GND.n6361 GND.n6360 19.3944
R12998 GND.n6360 GND.n6359 19.3944
R12999 GND.n6359 GND.n440 19.3944
R13000 GND.n1823 GND.n1820 19.3944
R13001 GND.n1823 GND.n1818 19.3944
R13002 GND.n1827 GND.n1818 19.3944
R13003 GND.n1827 GND.n1816 19.3944
R13004 GND.n1833 GND.n1816 19.3944
R13005 GND.n1833 GND.n1814 19.3944
R13006 GND.n1845 GND.n1812 19.3944
R13007 GND.n1845 GND.n1810 19.3944
R13008 GND.n1849 GND.n1810 19.3944
R13009 GND.n1849 GND.n1808 19.3944
R13010 GND.n1855 GND.n1808 19.3944
R13011 GND.n1855 GND.n1806 19.3944
R13012 GND.n1859 GND.n1806 19.3944
R13013 GND.n1865 GND.n1800 19.3944
R13014 GND.n1869 GND.n1800 19.3944
R13015 GND.n1869 GND.n1798 19.3944
R13016 GND.n1875 GND.n1798 19.3944
R13017 GND.n1875 GND.n1796 19.3944
R13018 GND.n1879 GND.n1796 19.3944
R13019 GND.n1879 GND.n1791 19.3944
R13020 GND.n1885 GND.n1791 19.3944
R13021 GND.n1889 GND.n1789 19.3944
R13022 GND.n1889 GND.n1787 19.3944
R13023 GND.n1895 GND.n1787 19.3944
R13024 GND.n1895 GND.n1785 19.3944
R13025 GND.n1899 GND.n1785 19.3944
R13026 GND.n1899 GND.n1783 19.3944
R13027 GND.n1905 GND.n1783 19.3944
R13028 GND.n1905 GND.n1781 19.3944
R13029 GND.n1917 GND.n1779 19.3944
R13030 GND.n1917 GND.n1777 19.3944
R13031 GND.n1921 GND.n1777 19.3944
R13032 GND.n1921 GND.n1775 19.3944
R13033 GND.n1927 GND.n1775 19.3944
R13034 GND.n1927 GND.n1773 19.3944
R13035 GND.n1931 GND.n1773 19.3944
R13036 GND.n5377 GND.n5376 19.3944
R13037 GND.n5376 GND.n5375 19.3944
R13038 GND.n5375 GND.n1285 19.3944
R13039 GND.n2010 GND.n1285 19.3944
R13040 GND.n2010 GND.n2009 19.3944
R13041 GND.n2009 GND.n1743 19.3944
R13042 GND.n2029 GND.n1743 19.3944
R13043 GND.n2029 GND.n1741 19.3944
R13044 GND.n2035 GND.n1741 19.3944
R13045 GND.n2035 GND.n2034 19.3944
R13046 GND.n2034 GND.n1713 19.3944
R13047 GND.n2082 GND.n1713 19.3944
R13048 GND.n2082 GND.n1711 19.3944
R13049 GND.n2088 GND.n1711 19.3944
R13050 GND.n2088 GND.n2087 19.3944
R13051 GND.n2087 GND.n1691 19.3944
R13052 GND.n2106 GND.n1691 19.3944
R13053 GND.n2106 GND.n1689 19.3944
R13054 GND.n2110 GND.n1689 19.3944
R13055 GND.n2110 GND.n1641 19.3944
R13056 GND.n2213 GND.n1641 19.3944
R13057 GND.n1640 GND.n1639 19.3944
R13058 GND.n1666 GND.n1639 19.3944
R13059 GND.n2197 GND.n2196 19.3944
R13060 GND.n2134 GND.n2133 19.3944
R13061 GND.n2218 GND.n1633 19.3944
R13062 GND.n2218 GND.n2217 19.3944
R13063 GND.n2217 GND.n1612 19.3944
R13064 GND.n2236 GND.n1612 19.3944
R13065 GND.n2236 GND.n1610 19.3944
R13066 GND.n2242 GND.n1610 19.3944
R13067 GND.n2242 GND.n2241 19.3944
R13068 GND.n2241 GND.n1589 19.3944
R13069 GND.n2261 GND.n1589 19.3944
R13070 GND.n2261 GND.n1587 19.3944
R13071 GND.n2267 GND.n1587 19.3944
R13072 GND.n2267 GND.n2266 19.3944
R13073 GND.n2266 GND.n1567 19.3944
R13074 GND.n2299 GND.n1567 19.3944
R13075 GND.n2299 GND.n1565 19.3944
R13076 GND.n2303 GND.n1565 19.3944
R13077 GND.n2303 GND.n1548 19.3944
R13078 GND.n2336 GND.n1548 19.3944
R13079 GND.n2336 GND.n1546 19.3944
R13080 GND.n2340 GND.n1546 19.3944
R13081 GND.n2340 GND.n1402 19.3944
R13082 GND.n5292 GND.n1402 19.3944
R13083 GND.n5416 GND.n5415 19.3944
R13084 GND.n5415 GND.n5414 19.3944
R13085 GND.n5414 GND.n1240 19.3944
R13086 GND.n5408 GND.n1240 19.3944
R13087 GND.n5408 GND.n5407 19.3944
R13088 GND.n5407 GND.n5406 19.3944
R13089 GND.n5406 GND.n1249 19.3944
R13090 GND.n5400 GND.n1249 19.3944
R13091 GND.n5400 GND.n5399 19.3944
R13092 GND.n5399 GND.n5398 19.3944
R13093 GND.n5398 GND.n1257 19.3944
R13094 GND.n5392 GND.n1257 19.3944
R13095 GND.n5392 GND.n5391 19.3944
R13096 GND.n5391 GND.n5390 19.3944
R13097 GND.n5390 GND.n1265 19.3944
R13098 GND.n5384 GND.n1265 19.3944
R13099 GND.n5384 GND.n5383 19.3944
R13100 GND.n5383 GND.n5382 19.3944
R13101 GND.n5382 GND.n1273 19.3944
R13102 GND.n1980 GND.n1273 19.3944
R13103 GND.n1983 GND.n1980 19.3944
R13104 GND.n1983 GND.n1977 19.3944
R13105 GND.n2000 GND.n1977 19.3944
R13106 GND.n2000 GND.n1999 19.3944
R13107 GND.n1999 GND.n1998 19.3944
R13108 GND.n1998 GND.n1989 19.3944
R13109 GND.n1994 GND.n1989 19.3944
R13110 GND.n1994 GND.n1993 19.3944
R13111 GND.n1993 GND.n1725 19.3944
R13112 GND.n2050 GND.n1725 19.3944
R13113 GND.n2050 GND.n1723 19.3944
R13114 GND.n2074 GND.n1723 19.3944
R13115 GND.n2074 GND.n2073 19.3944
R13116 GND.n2073 GND.n2072 19.3944
R13117 GND.n2072 GND.n2056 19.3944
R13118 GND.n2068 GND.n2056 19.3944
R13119 GND.n2068 GND.n2067 19.3944
R13120 GND.n2067 GND.n2066 19.3944
R13121 GND.n2066 GND.n2063 19.3944
R13122 GND.n2205 GND.n1655 19.3944
R13123 GND.n2205 GND.n2204 19.3944
R13124 GND.n2202 GND.n1656 19.3944
R13125 GND.n2188 GND.n2144 19.3944
R13126 GND.n2186 GND.n2185 19.3944
R13127 GND.n2182 GND.n2181 19.3944
R13128 GND.n2181 GND.n2180 19.3944
R13129 GND.n2180 GND.n2149 19.3944
R13130 GND.n2176 GND.n2149 19.3944
R13131 GND.n2176 GND.n2175 19.3944
R13132 GND.n2175 GND.n2174 19.3944
R13133 GND.n2174 GND.n2155 19.3944
R13134 GND.n2170 GND.n2155 19.3944
R13135 GND.n2170 GND.n2169 19.3944
R13136 GND.n2169 GND.n2168 19.3944
R13137 GND.n2168 GND.n2161 19.3944
R13138 GND.n2164 GND.n2161 19.3944
R13139 GND.n2164 GND.n1559 19.3944
R13140 GND.n2308 GND.n1559 19.3944
R13141 GND.n2308 GND.n1557 19.3944
R13142 GND.n2327 GND.n1557 19.3944
R13143 GND.n2327 GND.n2326 19.3944
R13144 GND.n2326 GND.n2325 19.3944
R13145 GND.n2325 GND.n2314 19.3944
R13146 GND.n2321 GND.n2314 19.3944
R13147 GND.n2321 GND.n2320 19.3944
R13148 GND.n2320 GND.n1527 19.3944
R13149 GND.n5166 GND.n1527 19.3944
R13150 GND.n5166 GND.n5165 19.3944
R13151 GND.n5165 GND.n5164 19.3944
R13152 GND.n5164 GND.n1531 19.3944
R13153 GND.n3516 GND.n1531 19.3944
R13154 GND.n3518 GND.n3516 19.3944
R13155 GND.n3518 GND.n3513 19.3944
R13156 GND.n3522 GND.n3513 19.3944
R13157 GND.n3522 GND.n3465 19.3944
R13158 GND.n3536 GND.n3465 19.3944
R13159 GND.n3536 GND.n3463 19.3944
R13160 GND.n3540 GND.n3463 19.3944
R13161 GND.n3540 GND.n3454 19.3944
R13162 GND.n3553 GND.n3454 19.3944
R13163 GND.n3553 GND.n3452 19.3944
R13164 GND.n3557 GND.n3452 19.3944
R13165 GND.n3557 GND.n3442 19.3944
R13166 GND.n3570 GND.n3442 19.3944
R13167 GND.n3570 GND.n3440 19.3944
R13168 GND.n3574 GND.n3440 19.3944
R13169 GND.n3574 GND.n3430 19.3944
R13170 GND.n3587 GND.n3430 19.3944
R13171 GND.n3587 GND.n3428 19.3944
R13172 GND.n3591 GND.n3428 19.3944
R13173 GND.n3591 GND.n3417 19.3944
R13174 GND.n3605 GND.n3417 19.3944
R13175 GND.n3605 GND.n3415 19.3944
R13176 GND.n3609 GND.n3415 19.3944
R13177 GND.n3609 GND.n3384 19.3944
R13178 GND.n3741 GND.n3384 19.3944
R13179 GND.n3741 GND.n3382 19.3944
R13180 GND.n3753 GND.n3382 19.3944
R13181 GND.n3753 GND.n3752 19.3944
R13182 GND.n3752 GND.n3751 19.3944
R13183 GND.n3751 GND.n3748 19.3944
R13184 GND.n3748 GND.n3346 19.3944
R13185 GND.n3787 GND.n3346 19.3944
R13186 GND.n3787 GND.n3344 19.3944
R13187 GND.n3793 GND.n3344 19.3944
R13188 GND.n3793 GND.n3792 19.3944
R13189 GND.n3792 GND.n3317 19.3944
R13190 GND.n3841 GND.n3317 19.3944
R13191 GND.n3841 GND.n3315 19.3944
R13192 GND.n3847 GND.n3315 19.3944
R13193 GND.n3847 GND.n3846 19.3944
R13194 GND.n3846 GND.n3293 19.3944
R13195 GND.n3902 GND.n3293 19.3944
R13196 GND.n3902 GND.n3291 19.3944
R13197 GND.n3914 GND.n3291 19.3944
R13198 GND.n3914 GND.n3913 19.3944
R13199 GND.n3913 GND.n3912 19.3944
R13200 GND.n3912 GND.n3909 19.3944
R13201 GND.n3909 GND.n3258 19.3944
R13202 GND.n3948 GND.n3258 19.3944
R13203 GND.n3948 GND.n3256 19.3944
R13204 GND.n3954 GND.n3256 19.3944
R13205 GND.n3954 GND.n3953 19.3944
R13206 GND.n3953 GND.n3230 19.3944
R13207 GND.n4001 GND.n3230 19.3944
R13208 GND.n4001 GND.n3228 19.3944
R13209 GND.n4007 GND.n3228 19.3944
R13210 GND.n4007 GND.n4006 19.3944
R13211 GND.n4006 GND.n3205 19.3944
R13212 GND.n4062 GND.n3205 19.3944
R13213 GND.n4062 GND.n3203 19.3944
R13214 GND.n4074 GND.n3203 19.3944
R13215 GND.n4074 GND.n4073 19.3944
R13216 GND.n4073 GND.n4072 19.3944
R13217 GND.n4072 GND.n4069 19.3944
R13218 GND.n4069 GND.n3172 19.3944
R13219 GND.n4108 GND.n3172 19.3944
R13220 GND.n4108 GND.n3170 19.3944
R13221 GND.n4114 GND.n3170 19.3944
R13222 GND.n4114 GND.n4113 19.3944
R13223 GND.n4113 GND.n3143 19.3944
R13224 GND.n4161 GND.n3143 19.3944
R13225 GND.n4161 GND.n3141 19.3944
R13226 GND.n4167 GND.n3141 19.3944
R13227 GND.n4167 GND.n4166 19.3944
R13228 GND.n4166 GND.n3118 19.3944
R13229 GND.n4209 GND.n3118 19.3944
R13230 GND.n4209 GND.n3116 19.3944
R13231 GND.n4224 GND.n3116 19.3944
R13232 GND.n4224 GND.n4223 19.3944
R13233 GND.n4223 GND.n4222 19.3944
R13234 GND.n4222 GND.n4215 19.3944
R13235 GND.n4218 GND.n4215 19.3944
R13236 GND.n4218 GND.n3077 19.3944
R13237 GND.n4323 GND.n3077 19.3944
R13238 GND.n4323 GND.n3075 19.3944
R13239 GND.n4329 GND.n3075 19.3944
R13240 GND.n4329 GND.n4328 19.3944
R13241 GND.n4328 GND.n3027 19.3944
R13242 GND.n4392 GND.n3027 19.3944
R13243 GND.n4392 GND.n3025 19.3944
R13244 GND.n4396 GND.n3025 19.3944
R13245 GND.n4396 GND.n3015 19.3944
R13246 GND.n4409 GND.n3015 19.3944
R13247 GND.n4409 GND.n3013 19.3944
R13248 GND.n4413 GND.n3013 19.3944
R13249 GND.n4413 GND.n3003 19.3944
R13250 GND.n4426 GND.n3003 19.3944
R13251 GND.n4426 GND.n3001 19.3944
R13252 GND.n4430 GND.n3001 19.3944
R13253 GND.n4430 GND.n2991 19.3944
R13254 GND.n4443 GND.n2991 19.3944
R13255 GND.n4443 GND.n2989 19.3944
R13256 GND.n4447 GND.n2989 19.3944
R13257 GND.n4447 GND.n2979 19.3944
R13258 GND.n4460 GND.n2979 19.3944
R13259 GND.n4460 GND.n2977 19.3944
R13260 GND.n4464 GND.n2977 19.3944
R13261 GND.n4464 GND.n2967 19.3944
R13262 GND.n4477 GND.n2967 19.3944
R13263 GND.n4477 GND.n2965 19.3944
R13264 GND.n4484 GND.n2965 19.3944
R13265 GND.n4484 GND.n4483 19.3944
R13266 GND.n4483 GND.n2955 19.3944
R13267 GND.n4498 GND.n2955 19.3944
R13268 GND.n4499 GND.n4498 19.3944
R13269 GND.n4499 GND.n2953 19.3944
R13270 GND.n4512 GND.n2953 19.3944
R13271 GND.n4512 GND.n4511 19.3944
R13272 GND.n4511 GND.n4510 19.3944
R13273 GND.n4510 GND.n4507 19.3944
R13274 GND.n4507 GND.n2617 19.3944
R13275 GND.n4861 GND.n2617 19.3944
R13276 GND.n4861 GND.n4860 19.3944
R13277 GND.n4860 GND.n4859 19.3944
R13278 GND.n4859 GND.n2621 19.3944
R13279 GND.n2764 GND.n2621 19.3944
R13280 GND.n2768 GND.n2764 19.3944
R13281 GND.n2768 GND.n2762 19.3944
R13282 GND.n2772 GND.n2762 19.3944
R13283 GND.n2772 GND.n2760 19.3944
R13284 GND.n2776 GND.n2760 19.3944
R13285 GND.n2776 GND.n2758 19.3944
R13286 GND.n2780 GND.n2758 19.3944
R13287 GND.n2780 GND.n2756 19.3944
R13288 GND.n2784 GND.n2756 19.3944
R13289 GND.n2784 GND.n2754 19.3944
R13290 GND.n2788 GND.n2754 19.3944
R13291 GND.n2788 GND.n2752 19.3944
R13292 GND.n2793 GND.n2752 19.3944
R13293 GND.n2793 GND.n2749 19.3944
R13294 GND.n2797 GND.n2749 19.3944
R13295 GND.n2798 GND.n2797 19.3944
R13296 GND.n2799 GND.n2798 19.3944
R13297 GND.n2803 GND.n2802 19.3944
R13298 GND.n4790 GND.n4789 19.3944
R13299 GND.n4787 GND.n2805 19.3944
R13300 GND.n2870 GND.n2869 19.3944
R13301 GND.n2867 GND.n2808 19.3944
R13302 GND.n2863 GND.n2808 19.3944
R13303 GND.n2863 GND.n2862 19.3944
R13304 GND.n2862 GND.n2861 19.3944
R13305 GND.n2861 GND.n2814 19.3944
R13306 GND.n2857 GND.n2814 19.3944
R13307 GND.n2857 GND.n2856 19.3944
R13308 GND.n2856 GND.n2855 19.3944
R13309 GND.n2855 GND.n2820 19.3944
R13310 GND.n2851 GND.n2820 19.3944
R13311 GND.n2851 GND.n2850 19.3944
R13312 GND.n2850 GND.n2849 19.3944
R13313 GND.n2849 GND.n2826 19.3944
R13314 GND.n2845 GND.n2826 19.3944
R13315 GND.n2845 GND.n2844 19.3944
R13316 GND.n2844 GND.n2843 19.3944
R13317 GND.n2843 GND.n2832 19.3944
R13318 GND.n2839 GND.n2832 19.3944
R13319 GND.n2839 GND.n2838 19.3944
R13320 GND.n2838 GND.n455 19.3944
R13321 GND.n6347 GND.n455 19.3944
R13322 GND.n6347 GND.n6346 19.3944
R13323 GND.n6346 GND.n6345 19.3944
R13324 GND.n6345 GND.n459 19.3944
R13325 GND.n6339 GND.n459 19.3944
R13326 GND.n6339 GND.n6338 19.3944
R13327 GND.n6338 GND.n6337 19.3944
R13328 GND.n6337 GND.n640 19.3944
R13329 GND.n6331 GND.n640 19.3944
R13330 GND.n6331 GND.n6330 19.3944
R13331 GND.n6330 GND.n6329 19.3944
R13332 GND.n6329 GND.n648 19.3944
R13333 GND.n6323 GND.n648 19.3944
R13334 GND.n6323 GND.n6322 19.3944
R13335 GND.n6322 GND.n6321 19.3944
R13336 GND.n6321 GND.n656 19.3944
R13337 GND.n6315 GND.n656 19.3944
R13338 GND.n6315 GND.n6314 19.3944
R13339 GND.n6314 GND.n6313 19.3944
R13340 GND.n5515 GND.n5514 19.3944
R13341 GND.n5514 GND.n5513 19.3944
R13342 GND.n5513 GND.n1144 19.3944
R13343 GND.n5507 GND.n1144 19.3944
R13344 GND.n5507 GND.n5506 19.3944
R13345 GND.n5506 GND.n5505 19.3944
R13346 GND.n5505 GND.n1152 19.3944
R13347 GND.n5499 GND.n1152 19.3944
R13348 GND.n5499 GND.n5498 19.3944
R13349 GND.n5498 GND.n5497 19.3944
R13350 GND.n5497 GND.n1160 19.3944
R13351 GND.n5491 GND.n1160 19.3944
R13352 GND.n5491 GND.n5490 19.3944
R13353 GND.n5490 GND.n5489 19.3944
R13354 GND.n5489 GND.n1168 19.3944
R13355 GND.n5483 GND.n1168 19.3944
R13356 GND.n5483 GND.n5482 19.3944
R13357 GND.n5482 GND.n5481 19.3944
R13358 GND.n5481 GND.n1176 19.3944
R13359 GND.n5475 GND.n1176 19.3944
R13360 GND.n5475 GND.n5474 19.3944
R13361 GND.n5474 GND.n5473 19.3944
R13362 GND.n5473 GND.n1184 19.3944
R13363 GND.n5467 GND.n1184 19.3944
R13364 GND.n5467 GND.n5466 19.3944
R13365 GND.n5466 GND.n5465 19.3944
R13366 GND.n5465 GND.n1192 19.3944
R13367 GND.n5459 GND.n1192 19.3944
R13368 GND.n5459 GND.n5458 19.3944
R13369 GND.n5458 GND.n5457 19.3944
R13370 GND.n5457 GND.n1200 19.3944
R13371 GND.n5451 GND.n1200 19.3944
R13372 GND.n5451 GND.n5450 19.3944
R13373 GND.n5450 GND.n5449 19.3944
R13374 GND.n5449 GND.n1208 19.3944
R13375 GND.n5443 GND.n1208 19.3944
R13376 GND.n5443 GND.n5442 19.3944
R13377 GND.n5442 GND.n5441 19.3944
R13378 GND.n5441 GND.n1216 19.3944
R13379 GND.n5435 GND.n1216 19.3944
R13380 GND.n5435 GND.n5434 19.3944
R13381 GND.n5434 GND.n5433 19.3944
R13382 GND.n5433 GND.n1224 19.3944
R13383 GND.n5427 GND.n1224 19.3944
R13384 GND.n5427 GND.n5426 19.3944
R13385 GND.n5426 GND.n5425 19.3944
R13386 GND.n5425 GND.n1232 19.3944
R13387 GND.n5419 GND.n1232 19.3944
R13388 GND.n3508 GND.n3472 19.3944
R13389 GND.n3508 GND.n3471 19.3944
R13390 GND.n3526 GND.n3471 19.3944
R13391 GND.n3526 GND.n3469 19.3944
R13392 GND.n3530 GND.n3469 19.3944
R13393 GND.n3530 GND.n3460 19.3944
R13394 GND.n3544 GND.n3460 19.3944
R13395 GND.n3544 GND.n3458 19.3944
R13396 GND.n3548 GND.n3458 19.3944
R13397 GND.n3548 GND.n3448 19.3944
R13398 GND.n3561 GND.n3448 19.3944
R13399 GND.n3561 GND.n3446 19.3944
R13400 GND.n3565 GND.n3446 19.3944
R13401 GND.n3565 GND.n3436 19.3944
R13402 GND.n3578 GND.n3436 19.3944
R13403 GND.n3578 GND.n3434 19.3944
R13404 GND.n3582 GND.n3434 19.3944
R13405 GND.n3582 GND.n3424 19.3944
R13406 GND.n3595 GND.n3424 19.3944
R13407 GND.n3595 GND.n3421 19.3944
R13408 GND.n3600 GND.n3421 19.3944
R13409 GND.n3600 GND.n3422 19.3944
R13410 GND.n3422 GND.n3411 19.3944
R13411 GND.n3614 GND.n3411 19.3944
R13412 GND.n3614 GND.n3408 19.3944
R13413 GND.n3646 GND.n3408 19.3944
R13414 GND.n3646 GND.n3409 19.3944
R13415 GND.n3642 GND.n3409 19.3944
R13416 GND.n3642 GND.n3641 19.3944
R13417 GND.n3641 GND.n3640 19.3944
R13418 GND.n3640 GND.n3622 19.3944
R13419 GND.n3636 GND.n3622 19.3944
R13420 GND.n3636 GND.n3635 19.3944
R13421 GND.n3635 GND.n3634 19.3944
R13422 GND.n3634 GND.n3625 19.3944
R13423 GND.n3630 GND.n3625 19.3944
R13424 GND.n3630 GND.n3629 19.3944
R13425 GND.n3629 GND.n3308 19.3944
R13426 GND.n3851 GND.n3308 19.3944
R13427 GND.n3851 GND.n3305 19.3944
R13428 GND.n3889 GND.n3305 19.3944
R13429 GND.n3889 GND.n3306 19.3944
R13430 GND.n3885 GND.n3306 19.3944
R13431 GND.n3885 GND.n3884 19.3944
R13432 GND.n3884 GND.n3883 19.3944
R13433 GND.n3883 GND.n3857 19.3944
R13434 GND.n3879 GND.n3857 19.3944
R13435 GND.n3879 GND.n3878 19.3944
R13436 GND.n3878 GND.n3877 19.3944
R13437 GND.n3877 GND.n3864 19.3944
R13438 GND.n3873 GND.n3864 19.3944
R13439 GND.n3873 GND.n3872 19.3944
R13440 GND.n3872 GND.n3871 19.3944
R13441 GND.n3871 GND.n3868 19.3944
R13442 GND.n3868 GND.n3220 19.3944
R13443 GND.n4011 GND.n3220 19.3944
R13444 GND.n4011 GND.n3217 19.3944
R13445 GND.n4050 GND.n3217 19.3944
R13446 GND.n4050 GND.n3218 19.3944
R13447 GND.n4046 GND.n3218 19.3944
R13448 GND.n4046 GND.n4045 19.3944
R13449 GND.n4045 GND.n4044 19.3944
R13450 GND.n4044 GND.n4017 19.3944
R13451 GND.n4040 GND.n4017 19.3944
R13452 GND.n4040 GND.n4039 19.3944
R13453 GND.n4039 GND.n4038 19.3944
R13454 GND.n4038 GND.n4025 19.3944
R13455 GND.n4034 GND.n4025 19.3944
R13456 GND.n4034 GND.n4033 19.3944
R13457 GND.n4033 GND.n4032 19.3944
R13458 GND.n4032 GND.n4029 19.3944
R13459 GND.n4029 GND.n3133 19.3944
R13460 GND.n4171 GND.n3133 19.3944
R13461 GND.n4171 GND.n3130 19.3944
R13462 GND.n4197 GND.n3130 19.3944
R13463 GND.n4197 GND.n3131 19.3944
R13464 GND.n4193 GND.n3131 19.3944
R13465 GND.n4193 GND.n4192 19.3944
R13466 GND.n4192 GND.n4191 19.3944
R13467 GND.n4191 GND.n4177 19.3944
R13468 GND.n4187 GND.n4177 19.3944
R13469 GND.n4187 GND.n4186 19.3944
R13470 GND.n4186 GND.n4185 19.3944
R13471 GND.n4185 GND.n4182 19.3944
R13472 GND.n4182 GND.n3068 19.3944
R13473 GND.n4333 GND.n3068 19.3944
R13474 GND.n4333 GND.n3065 19.3944
R13475 GND.n4338 GND.n3065 19.3944
R13476 GND.n4338 GND.n3066 19.3944
R13477 GND.n3066 GND.n3021 19.3944
R13478 GND.n4400 GND.n3021 19.3944
R13479 GND.n4400 GND.n3019 19.3944
R13480 GND.n4404 GND.n3019 19.3944
R13481 GND.n4404 GND.n3009 19.3944
R13482 GND.n4417 GND.n3009 19.3944
R13483 GND.n4417 GND.n3007 19.3944
R13484 GND.n4421 GND.n3007 19.3944
R13485 GND.n4421 GND.n2997 19.3944
R13486 GND.n4434 GND.n2997 19.3944
R13487 GND.n4434 GND.n2995 19.3944
R13488 GND.n4438 GND.n2995 19.3944
R13489 GND.n4438 GND.n2985 19.3944
R13490 GND.n4451 GND.n2985 19.3944
R13491 GND.n4451 GND.n2983 19.3944
R13492 GND.n4455 GND.n2983 19.3944
R13493 GND.n4455 GND.n2972 19.3944
R13494 GND.n4468 GND.n2972 19.3944
R13495 GND.n4468 GND.n2970 19.3944
R13496 GND.n4472 GND.n2970 19.3944
R13497 GND.n4472 GND.n2961 19.3944
R13498 GND.n4488 GND.n2961 19.3944
R13499 GND.n4488 GND.n2959 19.3944
R13500 GND.n4492 GND.n2959 19.3944
R13501 GND.n4492 GND.n2499 19.3944
R13502 GND.n4980 GND.n2499 19.3944
R13503 GND.n3504 GND.n3503 19.3944
R13504 GND.n3503 GND.n3502 19.3944
R13505 GND.n3502 GND.n3478 19.3944
R13506 GND.n3498 GND.n3478 19.3944
R13507 GND.n3498 GND.n3497 19.3944
R13508 GND.n3497 GND.n3496 19.3944
R13509 GND.n3496 GND.n3486 19.3944
R13510 GND.n3492 GND.n3486 19.3944
R13511 GND.n3492 GND.n1472 19.3944
R13512 GND.n5220 GND.n1472 19.3944
R13513 GND.n5220 GND.n5219 19.3944
R13514 GND.n5219 GND.n1475 19.3944
R13515 GND.n5212 GND.n1475 19.3944
R13516 GND.n5212 GND.n5211 19.3944
R13517 GND.n5211 GND.n1484 19.3944
R13518 GND.n2076 GND.t5 18.7605
R13519 GND.t2 GND.n1591 18.7605
R13520 GND.n3849 GND.n3311 18.7605
R13521 GND.n3900 GND.n3295 18.7605
R13522 GND.n4009 GND.n3223 18.7605
R13523 GND.n4060 GND.n3207 18.7605
R13524 GND.n4169 GND.n3136 18.7605
R13525 GND.n4207 GND.n3120 18.7605
R13526 GND.t12 GND.n2690 18.7605
R13527 GND.t21 GND.n379 18.7605
R13528 GND.n3758 GND.n3376 18.2639
R13529 GND.n4345 GND.n4344 18.2639
R13530 GND.n5204 GND.n1490 17.455
R13531 GND.n4519 GND.n2903 17.455
R13532 GND.n3756 GND.n3755 17.1972
R13533 GND.n3839 GND.n3837 17.1972
R13534 GND.n3917 GND.n3916 17.1972
R13535 GND.n3999 GND.n3998 17.1972
R13536 GND.n4077 GND.n4076 17.1972
R13537 GND.n4159 GND.n4158 17.1972
R13538 GND.n4227 GND.n4226 17.1972
R13539 GND.n5265 GND.n1424 16.4853
R13540 GND.n4926 GND.n4925 16.4853
R13541 GND.n561 GND.n510 16.4853
R13542 GND.n1859 GND.n1804 16.4853
R13543 GND.n5227 GND.n5226 16.2914
R13544 GND.n4873 GND.n2607 16.2914
R13545 GND.n630 GND.n629 16.2914
R13546 GND.n1931 GND.n1771 16.2914
R13547 GND.n5239 GND.n5238 16.0975
R13548 GND.n4889 GND.n4888 16.0975
R13549 GND.n612 GND.n609 16.0975
R13550 GND.n1911 GND.n1779 16.0975
R13551 GND.n3333 GND.t161 16.0247
R13552 GND.t158 GND.n3105 16.0247
R13553 GND.n5277 GND.n1414 15.9035
R13554 GND.n4942 GND.n4941 15.9035
R13555 GND.n541 GND.n514 15.9035
R13556 GND.n1839 GND.n1812 15.9035
R13557 GND.n1275 GND.n1267 15.6338
R13558 GND.n5191 GND.n1505 15.6338
R13559 GND.n3368 GND.n3363 15.6338
R13560 GND.n3280 GND.n3275 15.6338
R13561 GND.n3248 GND.n3247 15.6338
R13562 GND.n3192 GND.n3187 15.6338
R13563 GND.n3161 GND.n3159 15.6338
R13564 GND.n4331 GND.n3071 15.6338
R13565 GND.n4957 GND.n2543 15.6338
R13566 GND.n633 GND.n452 15.6338
R13567 GND.n133 GND.n132 15.3979
R13568 GND.n146 GND.n145 15.3979
R13569 GND.n107 GND.n106 15.3979
R13570 GND.n120 GND.n119 15.3979
R13571 GND.n81 GND.n80 15.3979
R13572 GND.n94 GND.n93 15.3979
R13573 GND.n55 GND.n54 15.3979
R13574 GND.n68 GND.n67 15.3979
R13575 GND.n29 GND.n28 15.3979
R13576 GND.n42 GND.n41 15.3979
R13577 GND.n4 GND.n3 15.3979
R13578 GND.n17 GND.n16 15.3979
R13579 GND.n302 GND.n301 15.3979
R13580 GND.n289 GND.n288 15.3979
R13581 GND.n276 GND.n275 15.3979
R13582 GND.n263 GND.n262 15.3979
R13583 GND.n250 GND.n249 15.3979
R13584 GND.n237 GND.n236 15.3979
R13585 GND.n224 GND.n223 15.3979
R13586 GND.n211 GND.n210 15.3979
R13587 GND.n198 GND.n197 15.3979
R13588 GND.n185 GND.n184 15.3979
R13589 GND.n173 GND.n172 15.3979
R13590 GND.n160 GND.n159 15.3979
R13591 GND.n3739 GND.n3737 15.243
R13592 GND.n2002 GND.t63 14.8522
R13593 GND.n2329 GND.t77 14.8522
R13594 GND.n3648 GND.t92 14.8522
R13595 GND.t59 GND.n2643 14.8522
R13596 GND.t52 GND.n424 14.8522
R13597 GND.n4523 GND.n4522 14.7399
R13598 GND.n1503 GND.n1488 14.7399
R13599 GND.n1958 GND.n1761 14.7399
R13600 GND.n4702 GND.n4679 14.7399
R13601 GND.n3777 GND.n3357 14.0705
R13602 GND.n3796 GND.n3339 14.0705
R13603 GND.n3938 GND.n3270 14.0705
R13604 GND.n4117 GND.n3165 14.0705
R13605 GND.n4246 GND.n3096 14.0705
R13606 GND.n4321 GND.n4320 14.0705
R13607 GND.n3603 GND.t159 13.6797
R13608 GND.t162 GND.n3011 13.6797
R13609 GND.n2208 GND.t19 13.2888
R13610 GND.n2140 GND.t0 13.2888
R13611 GND.t122 GND.n3029 13.2888
R13612 GND.n4623 GND.t9 13.2888
R13613 GND.n4774 GND.t15 13.2888
R13614 GND.n3375 GND.n3372 13.1884
R13615 GND.n3059 GND.n3056 13.1884
R13616 GND.n3650 GND.n3376 13.1127
R13617 GND.n4386 GND.n4345 13.1127
R13618 GND.n136 GND.n131 12.8005
R13619 GND.n149 GND.n144 12.8005
R13620 GND.n110 GND.n105 12.8005
R13621 GND.n123 GND.n118 12.8005
R13622 GND.n84 GND.n79 12.8005
R13623 GND.n97 GND.n92 12.8005
R13624 GND.n58 GND.n53 12.8005
R13625 GND.n71 GND.n66 12.8005
R13626 GND.n32 GND.n27 12.8005
R13627 GND.n45 GND.n40 12.8005
R13628 GND.n7 GND.n2 12.8005
R13629 GND.n20 GND.n15 12.8005
R13630 GND.n305 GND.n300 12.8005
R13631 GND.n292 GND.n287 12.8005
R13632 GND.n279 GND.n274 12.8005
R13633 GND.n266 GND.n261 12.8005
R13634 GND.n253 GND.n248 12.8005
R13635 GND.n240 GND.n235 12.8005
R13636 GND.n227 GND.n222 12.8005
R13637 GND.n214 GND.n209 12.8005
R13638 GND.n201 GND.n196 12.8005
R13639 GND.n188 GND.n183 12.8005
R13640 GND.n176 GND.n171 12.8005
R13641 GND.n163 GND.n158 12.8005
R13642 GND.n3357 GND.n3348 12.5072
R13643 GND.n3351 GND.n3339 12.5072
R13644 GND.n3270 GND.n3260 12.5072
R13645 GND.n3862 GND.n3263 12.5072
R13646 GND.n4022 GND.n3174 12.5072
R13647 GND.n3177 GND.n3165 12.5072
R13648 GND.n3096 GND.n3088 12.5072
R13649 GND.n4321 GND.n3079 12.5072
R13650 GND.n3542 GND.t88 12.1163
R13651 GND.n2975 GND.t81 12.1163
R13652 GND.n137 GND.n129 12.0247
R13653 GND.n150 GND.n142 12.0247
R13654 GND.n111 GND.n103 12.0247
R13655 GND.n124 GND.n116 12.0247
R13656 GND.n85 GND.n77 12.0247
R13657 GND.n98 GND.n90 12.0247
R13658 GND.n59 GND.n51 12.0247
R13659 GND.n72 GND.n64 12.0247
R13660 GND.n33 GND.n25 12.0247
R13661 GND.n46 GND.n38 12.0247
R13662 GND.n8 GND.n0 12.0247
R13663 GND.n21 GND.n13 12.0247
R13664 GND.n306 GND.n298 12.0247
R13665 GND.n293 GND.n285 12.0247
R13666 GND.n280 GND.n272 12.0247
R13667 GND.n267 GND.n259 12.0247
R13668 GND.n254 GND.n246 12.0247
R13669 GND.n241 GND.n233 12.0247
R13670 GND.n228 GND.n220 12.0247
R13671 GND.n215 GND.n207 12.0247
R13672 GND.n202 GND.n194 12.0247
R13673 GND.n189 GND.n181 12.0247
R13674 GND.n177 GND.n169 12.0247
R13675 GND.n164 GND.n156 12.0247
R13676 GND.n4523 GND.n2906 11.249
R13677 GND.n5194 GND.n1503 11.249
R13678 GND.n1963 GND.n1761 11.249
R13679 GND.n4707 GND.n4679 11.249
R13680 GND.n3769 GND.n3363 10.9438
R13681 GND.n3802 GND.n3334 10.9438
R13682 GND.n3930 GND.n3275 10.9438
R13683 GND.n3963 GND.n3248 10.9438
R13684 GND.n4090 GND.n3187 10.9438
R13685 GND.n4123 GND.n3161 10.9438
R13686 GND.n4240 GND.n3100 10.9438
R13687 GND.n4331 GND.n3070 10.9438
R13688 GND.n5258 GND.n1432 10.6672
R13689 GND.n4918 GND.n4917 10.6672
R13690 GND.n4257 GND.n4256 10.6151
R13691 GND.n4260 GND.n4257 10.6151
R13692 GND.n4261 GND.n4260 10.6151
R13693 GND.n4265 GND.n4264 10.6151
R13694 GND.n4268 GND.n4265 10.6151
R13695 GND.n4269 GND.n4268 10.6151
R13696 GND.n4272 GND.n4269 10.6151
R13697 GND.n4273 GND.n4272 10.6151
R13698 GND.n4276 GND.n4273 10.6151
R13699 GND.n4277 GND.n4276 10.6151
R13700 GND.n4280 GND.n4277 10.6151
R13701 GND.n4281 GND.n4280 10.6151
R13702 GND.n4284 GND.n4281 10.6151
R13703 GND.n4285 GND.n4284 10.6151
R13704 GND.n4288 GND.n4285 10.6151
R13705 GND.n4289 GND.n4288 10.6151
R13706 GND.n4292 GND.n4289 10.6151
R13707 GND.n4293 GND.n4292 10.6151
R13708 GND.n3655 GND.n3365 10.6151
R13709 GND.n3764 GND.n3365 10.6151
R13710 GND.n3765 GND.n3764 10.6151
R13711 GND.n3766 GND.n3765 10.6151
R13712 GND.n3766 GND.n3354 10.6151
R13713 GND.n3779 GND.n3354 10.6151
R13714 GND.n3780 GND.n3779 10.6151
R13715 GND.n3783 GND.n3780 10.6151
R13716 GND.n3783 GND.n3782 10.6151
R13717 GND.n3782 GND.n3781 10.6151
R13718 GND.n3781 GND.n3330 10.6151
R13719 GND.n3804 GND.n3330 10.6151
R13720 GND.n3805 GND.n3804 10.6151
R13721 GND.n3824 GND.n3805 10.6151
R13722 GND.n3824 GND.n3823 10.6151
R13723 GND.n3823 GND.n3822 10.6151
R13724 GND.n3822 GND.n3821 10.6151
R13725 GND.n3821 GND.n3806 10.6151
R13726 GND.n3816 GND.n3806 10.6151
R13727 GND.n3816 GND.n3815 10.6151
R13728 GND.n3815 GND.n3814 10.6151
R13729 GND.n3814 GND.n3813 10.6151
R13730 GND.n3813 GND.n3811 10.6151
R13731 GND.n3811 GND.n3810 10.6151
R13732 GND.n3810 GND.n3808 10.6151
R13733 GND.n3808 GND.n3277 10.6151
R13734 GND.n3925 GND.n3277 10.6151
R13735 GND.n3926 GND.n3925 10.6151
R13736 GND.n3927 GND.n3926 10.6151
R13737 GND.n3927 GND.n3267 10.6151
R13738 GND.n3940 GND.n3267 10.6151
R13739 GND.n3941 GND.n3940 10.6151
R13740 GND.n3944 GND.n3941 10.6151
R13741 GND.n3944 GND.n3943 10.6151
R13742 GND.n3943 GND.n3942 10.6151
R13743 GND.n3942 GND.n3244 10.6151
R13744 GND.n3965 GND.n3244 10.6151
R13745 GND.n3966 GND.n3965 10.6151
R13746 GND.n3985 GND.n3966 10.6151
R13747 GND.n3985 GND.n3984 10.6151
R13748 GND.n3984 GND.n3983 10.6151
R13749 GND.n3983 GND.n3982 10.6151
R13750 GND.n3982 GND.n3967 10.6151
R13751 GND.n3977 GND.n3967 10.6151
R13752 GND.n3977 GND.n3976 10.6151
R13753 GND.n3976 GND.n3975 10.6151
R13754 GND.n3975 GND.n3974 10.6151
R13755 GND.n3974 GND.n3972 10.6151
R13756 GND.n3972 GND.n3971 10.6151
R13757 GND.n3971 GND.n3969 10.6151
R13758 GND.n3969 GND.n3189 10.6151
R13759 GND.n4085 GND.n3189 10.6151
R13760 GND.n4086 GND.n4085 10.6151
R13761 GND.n4087 GND.n4086 10.6151
R13762 GND.n4087 GND.n3180 10.6151
R13763 GND.n4100 GND.n3180 10.6151
R13764 GND.n4101 GND.n4100 10.6151
R13765 GND.n4104 GND.n4101 10.6151
R13766 GND.n4104 GND.n4103 10.6151
R13767 GND.n4103 GND.n4102 10.6151
R13768 GND.n4102 GND.n3156 10.6151
R13769 GND.n4125 GND.n3156 10.6151
R13770 GND.n4126 GND.n4125 10.6151
R13771 GND.n4145 GND.n4126 10.6151
R13772 GND.n4145 GND.n4144 10.6151
R13773 GND.n4144 GND.n4143 10.6151
R13774 GND.n4143 GND.n4142 10.6151
R13775 GND.n4142 GND.n4127 10.6151
R13776 GND.n4137 GND.n4127 10.6151
R13777 GND.n4137 GND.n4136 10.6151
R13778 GND.n4136 GND.n4135 10.6151
R13779 GND.n4135 GND.n4134 10.6151
R13780 GND.n4134 GND.n4132 10.6151
R13781 GND.n4132 GND.n4131 10.6151
R13782 GND.n4131 GND.n4129 10.6151
R13783 GND.n4129 GND.n3102 10.6151
R13784 GND.n4235 GND.n3102 10.6151
R13785 GND.n4236 GND.n4235 10.6151
R13786 GND.n4237 GND.n4236 10.6151
R13787 GND.n4237 GND.n3092 10.6151
R13788 GND.n4248 GND.n3092 10.6151
R13789 GND.n4249 GND.n4248 10.6151
R13790 GND.n4307 GND.n4249 10.6151
R13791 GND.n4307 GND.n4306 10.6151
R13792 GND.n4306 GND.n4305 10.6151
R13793 GND.n4305 GND.n4304 10.6151
R13794 GND.n4304 GND.n4250 10.6151
R13795 GND.n4299 GND.n4250 10.6151
R13796 GND.n4299 GND.n4298 10.6151
R13797 GND.n4298 GND.n4297 10.6151
R13798 GND.n4297 GND.n4296 10.6151
R13799 GND.n3695 GND.n3692 10.6151
R13800 GND.n3692 GND.n3691 10.6151
R13801 GND.n3691 GND.n3688 10.6151
R13802 GND.n3686 GND.n3683 10.6151
R13803 GND.n3683 GND.n3682 10.6151
R13804 GND.n3682 GND.n3679 10.6151
R13805 GND.n3679 GND.n3678 10.6151
R13806 GND.n3678 GND.n3675 10.6151
R13807 GND.n3675 GND.n3674 10.6151
R13808 GND.n3674 GND.n3671 10.6151
R13809 GND.n3671 GND.n3670 10.6151
R13810 GND.n3670 GND.n3667 10.6151
R13811 GND.n3667 GND.n3666 10.6151
R13812 GND.n3666 GND.n3663 10.6151
R13813 GND.n3663 GND.n3662 10.6151
R13814 GND.n3662 GND.n3659 10.6151
R13815 GND.n3659 GND.n3658 10.6151
R13816 GND.n3658 GND.n3656 10.6151
R13817 GND.n3734 GND.n3650 10.6151
R13818 GND.n3734 GND.n3733 10.6151
R13819 GND.n3733 GND.n3732 10.6151
R13820 GND.n3732 GND.n3730 10.6151
R13821 GND.n3730 GND.n3727 10.6151
R13822 GND.n3727 GND.n3726 10.6151
R13823 GND.n3726 GND.n3723 10.6151
R13824 GND.n3723 GND.n3722 10.6151
R13825 GND.n3722 GND.n3719 10.6151
R13826 GND.n3719 GND.n3718 10.6151
R13827 GND.n3718 GND.n3715 10.6151
R13828 GND.n3715 GND.n3714 10.6151
R13829 GND.n3714 GND.n3711 10.6151
R13830 GND.n3711 GND.n3710 10.6151
R13831 GND.n3710 GND.n3707 10.6151
R13832 GND.n3705 GND.n3702 10.6151
R13833 GND.n3702 GND.n3701 10.6151
R13834 GND.n3701 GND.n3698 10.6151
R13835 GND.n4386 GND.n4385 10.6151
R13836 GND.n4385 GND.n4384 10.6151
R13837 GND.n4384 GND.n4381 10.6151
R13838 GND.n4381 GND.n4380 10.6151
R13839 GND.n4380 GND.n4377 10.6151
R13840 GND.n4377 GND.n4376 10.6151
R13841 GND.n4376 GND.n4373 10.6151
R13842 GND.n4373 GND.n4372 10.6151
R13843 GND.n4372 GND.n4369 10.6151
R13844 GND.n4369 GND.n4368 10.6151
R13845 GND.n4368 GND.n4365 10.6151
R13846 GND.n4365 GND.n4364 10.6151
R13847 GND.n4364 GND.n4361 10.6151
R13848 GND.n4361 GND.n4360 10.6151
R13849 GND.n4360 GND.n4357 10.6151
R13850 GND.n4355 GND.n4352 10.6151
R13851 GND.n4352 GND.n4351 10.6151
R13852 GND.n4351 GND.n4348 10.6151
R13853 GND.n3759 GND.n3758 10.6151
R13854 GND.n3760 GND.n3759 10.6151
R13855 GND.n3760 GND.n3360 10.6151
R13856 GND.n3771 GND.n3360 10.6151
R13857 GND.n3772 GND.n3771 10.6151
R13858 GND.n3775 GND.n3772 10.6151
R13859 GND.n3775 GND.n3774 10.6151
R13860 GND.n3774 GND.n3773 10.6151
R13861 GND.n3773 GND.n3336 10.6151
R13862 GND.n3798 GND.n3336 10.6151
R13863 GND.n3799 GND.n3798 10.6151
R13864 GND.n3800 GND.n3799 10.6151
R13865 GND.n3800 GND.n3325 10.6151
R13866 GND.n3828 GND.n3325 10.6151
R13867 GND.n3829 GND.n3828 10.6151
R13868 GND.n3835 GND.n3829 10.6151
R13869 GND.n3835 GND.n3834 10.6151
R13870 GND.n3834 GND.n3833 10.6151
R13871 GND.n3833 GND.n3830 10.6151
R13872 GND.n3830 GND.n3300 10.6151
R13873 GND.n3895 GND.n3300 10.6151
R13874 GND.n3896 GND.n3895 10.6151
R13875 GND.n3897 GND.n3896 10.6151
R13876 GND.n3897 GND.n3284 10.6151
R13877 GND.n3919 GND.n3284 10.6151
R13878 GND.n3920 GND.n3919 10.6151
R13879 GND.n3921 GND.n3920 10.6151
R13880 GND.n3921 GND.n3273 10.6151
R13881 GND.n3932 GND.n3273 10.6151
R13882 GND.n3933 GND.n3932 10.6151
R13883 GND.n3936 GND.n3933 10.6151
R13884 GND.n3936 GND.n3935 10.6151
R13885 GND.n3935 GND.n3934 10.6151
R13886 GND.n3934 GND.n3250 10.6151
R13887 GND.n3959 GND.n3250 10.6151
R13888 GND.n3960 GND.n3959 10.6151
R13889 GND.n3961 GND.n3960 10.6151
R13890 GND.n3961 GND.n3238 10.6151
R13891 GND.n3989 GND.n3238 10.6151
R13892 GND.n3990 GND.n3989 10.6151
R13893 GND.n3996 GND.n3990 10.6151
R13894 GND.n3996 GND.n3995 10.6151
R13895 GND.n3995 GND.n3994 10.6151
R13896 GND.n3994 GND.n3991 10.6151
R13897 GND.n3991 GND.n3212 10.6151
R13898 GND.n4055 GND.n3212 10.6151
R13899 GND.n4056 GND.n4055 10.6151
R13900 GND.n4057 GND.n4056 10.6151
R13901 GND.n4057 GND.n3195 10.6151
R13902 GND.n4079 GND.n3195 10.6151
R13903 GND.n4080 GND.n4079 10.6151
R13904 GND.n4081 GND.n4080 10.6151
R13905 GND.n4081 GND.n3185 10.6151
R13906 GND.n4092 GND.n3185 10.6151
R13907 GND.n4093 GND.n4092 10.6151
R13908 GND.n4096 GND.n4093 10.6151
R13909 GND.n4096 GND.n4095 10.6151
R13910 GND.n4095 GND.n4094 10.6151
R13911 GND.n4094 GND.n3163 10.6151
R13912 GND.n4119 GND.n3163 10.6151
R13913 GND.n4120 GND.n4119 10.6151
R13914 GND.n4121 GND.n4120 10.6151
R13915 GND.n4121 GND.n3151 10.6151
R13916 GND.n4149 GND.n3151 10.6151
R13917 GND.n4150 GND.n4149 10.6151
R13918 GND.n4156 GND.n4150 10.6151
R13919 GND.n4156 GND.n4155 10.6151
R13920 GND.n4155 GND.n4154 10.6151
R13921 GND.n4154 GND.n4151 10.6151
R13922 GND.n4151 GND.n3125 10.6151
R13923 GND.n4202 GND.n3125 10.6151
R13924 GND.n4203 GND.n4202 10.6151
R13925 GND.n4204 GND.n4203 10.6151
R13926 GND.n4204 GND.n3108 10.6151
R13927 GND.n4229 GND.n3108 10.6151
R13928 GND.n4230 GND.n4229 10.6151
R13929 GND.n4231 GND.n4230 10.6151
R13930 GND.n4231 GND.n3098 10.6151
R13931 GND.n4242 GND.n3098 10.6151
R13932 GND.n4243 GND.n4242 10.6151
R13933 GND.n4244 GND.n4243 10.6151
R13934 GND.n4244 GND.n3086 10.6151
R13935 GND.n4311 GND.n3086 10.6151
R13936 GND.n4312 GND.n4311 10.6151
R13937 GND.n4318 GND.n4312 10.6151
R13938 GND.n4318 GND.n4317 10.6151
R13939 GND.n4317 GND.n4316 10.6151
R13940 GND.n4316 GND.n4313 10.6151
R13941 GND.n4313 GND.n3060 10.6151
R13942 GND.n4343 GND.n3060 10.6151
R13943 GND.n4344 GND.n4343 10.6151
R13944 GND.n5162 GND.n1495 10.553
R13945 GND.n4515 GND.n4514 10.553
R13946 GND.n5281 GND.n1414 10.0853
R13947 GND.n4945 GND.n4942 10.0853
R13948 GND.n541 GND.n540 10.0853
R13949 GND.n1839 GND.n1814 10.0853
R13950 GND.n5240 GND.n5239 9.89141
R13951 GND.n4892 GND.n4889 9.89141
R13952 GND.n609 GND.n608 9.89141
R13953 GND.n1911 GND.n1781 9.89141
R13954 GND.n5226 GND.n5225 9.69747
R13955 GND.n4869 GND.n2607 9.69747
R13956 GND.n630 GND.n484 9.69747
R13957 GND.n1936 GND.n1771 9.69747
R13958 GND.n5265 GND.n5264 9.50353
R13959 GND.n4925 GND.n4924 9.50353
R13960 GND.n565 GND.n510 9.50353
R13961 GND.n1865 GND.n1804 9.50353
R13962 GND.n139 GND.n138 9.45567
R13963 GND.n152 GND.n151 9.45567
R13964 GND.n113 GND.n112 9.45567
R13965 GND.n126 GND.n125 9.45567
R13966 GND.n87 GND.n86 9.45567
R13967 GND.n100 GND.n99 9.45567
R13968 GND.n61 GND.n60 9.45567
R13969 GND.n74 GND.n73 9.45567
R13970 GND.n35 GND.n34 9.45567
R13971 GND.n48 GND.n47 9.45567
R13972 GND.n10 GND.n9 9.45567
R13973 GND.n23 GND.n22 9.45567
R13974 GND.n308 GND.n307 9.45567
R13975 GND.n295 GND.n294 9.45567
R13976 GND.n282 GND.n281 9.45567
R13977 GND.n269 GND.n268 9.45567
R13978 GND.n256 GND.n255 9.45567
R13979 GND.n243 GND.n242 9.45567
R13980 GND.n230 GND.n229 9.45567
R13981 GND.n217 GND.n216 9.45567
R13982 GND.n204 GND.n203 9.45567
R13983 GND.n191 GND.n190 9.45567
R13984 GND.n179 GND.n178 9.45567
R13985 GND.n166 GND.n165 9.45567
R13986 GND.n3755 GND.n3367 9.3805
R13987 GND.n3839 GND.n3319 9.3805
R13988 GND.n3916 GND.n3279 9.3805
R13989 GND.n3999 GND.n3232 9.3805
R13990 GND.n4076 GND.n3191 9.3805
R13991 GND.n4159 GND.n3145 9.3805
R13992 GND.n4226 GND.n3104 9.3805
R13993 GND.n4341 GND.n4340 9.3805
R13994 GND.t152 GND.n3023 9.3805
R13995 GND.n4264 GND.n4254 9.36635
R13996 GND.n3687 GND.n3686 9.36635
R13997 GND.n3707 GND.n3706 9.36635
R13998 GND.n4357 GND.n4356 9.36635
R13999 GND.n138 GND.n137 9.3005
R14000 GND.n131 GND.n130 9.3005
R14001 GND.n151 GND.n150 9.3005
R14002 GND.n144 GND.n143 9.3005
R14003 GND.n112 GND.n111 9.3005
R14004 GND.n105 GND.n104 9.3005
R14005 GND.n125 GND.n124 9.3005
R14006 GND.n118 GND.n117 9.3005
R14007 GND.n86 GND.n85 9.3005
R14008 GND.n79 GND.n78 9.3005
R14009 GND.n99 GND.n98 9.3005
R14010 GND.n92 GND.n91 9.3005
R14011 GND.n60 GND.n59 9.3005
R14012 GND.n53 GND.n52 9.3005
R14013 GND.n73 GND.n72 9.3005
R14014 GND.n66 GND.n65 9.3005
R14015 GND.n34 GND.n33 9.3005
R14016 GND.n27 GND.n26 9.3005
R14017 GND.n47 GND.n46 9.3005
R14018 GND.n40 GND.n39 9.3005
R14019 GND.n9 GND.n8 9.3005
R14020 GND.n2 GND.n1 9.3005
R14021 GND.n22 GND.n21 9.3005
R14022 GND.n15 GND.n14 9.3005
R14023 GND.n1137 GND.n1136 9.3005
R14024 GND.n5522 GND.n5521 9.3005
R14025 GND.n5523 GND.n1135 9.3005
R14026 GND.n5525 GND.n5524 9.3005
R14027 GND.n1131 GND.n1130 9.3005
R14028 GND.n5532 GND.n5531 9.3005
R14029 GND.n5533 GND.n1129 9.3005
R14030 GND.n5535 GND.n5534 9.3005
R14031 GND.n1125 GND.n1124 9.3005
R14032 GND.n5542 GND.n5541 9.3005
R14033 GND.n5543 GND.n1123 9.3005
R14034 GND.n5545 GND.n5544 9.3005
R14035 GND.n1119 GND.n1118 9.3005
R14036 GND.n5552 GND.n5551 9.3005
R14037 GND.n5553 GND.n1117 9.3005
R14038 GND.n5555 GND.n5554 9.3005
R14039 GND.n1113 GND.n1112 9.3005
R14040 GND.n5562 GND.n5561 9.3005
R14041 GND.n5563 GND.n1111 9.3005
R14042 GND.n5565 GND.n5564 9.3005
R14043 GND.n1107 GND.n1106 9.3005
R14044 GND.n5572 GND.n5571 9.3005
R14045 GND.n5573 GND.n1105 9.3005
R14046 GND.n5575 GND.n5574 9.3005
R14047 GND.n1101 GND.n1100 9.3005
R14048 GND.n5582 GND.n5581 9.3005
R14049 GND.n5583 GND.n1099 9.3005
R14050 GND.n5585 GND.n5584 9.3005
R14051 GND.n1095 GND.n1094 9.3005
R14052 GND.n5592 GND.n5591 9.3005
R14053 GND.n5593 GND.n1093 9.3005
R14054 GND.n5595 GND.n5594 9.3005
R14055 GND.n1089 GND.n1088 9.3005
R14056 GND.n5602 GND.n5601 9.3005
R14057 GND.n5603 GND.n1087 9.3005
R14058 GND.n5605 GND.n5604 9.3005
R14059 GND.n1083 GND.n1082 9.3005
R14060 GND.n5612 GND.n5611 9.3005
R14061 GND.n5613 GND.n1081 9.3005
R14062 GND.n5615 GND.n5614 9.3005
R14063 GND.n1077 GND.n1076 9.3005
R14064 GND.n5622 GND.n5621 9.3005
R14065 GND.n5623 GND.n1075 9.3005
R14066 GND.n5625 GND.n5624 9.3005
R14067 GND.n1071 GND.n1070 9.3005
R14068 GND.n5632 GND.n5631 9.3005
R14069 GND.n5633 GND.n1069 9.3005
R14070 GND.n5635 GND.n5634 9.3005
R14071 GND.n1065 GND.n1064 9.3005
R14072 GND.n5642 GND.n5641 9.3005
R14073 GND.n5643 GND.n1063 9.3005
R14074 GND.n5645 GND.n5644 9.3005
R14075 GND.n1059 GND.n1058 9.3005
R14076 GND.n5652 GND.n5651 9.3005
R14077 GND.n5653 GND.n1057 9.3005
R14078 GND.n5655 GND.n5654 9.3005
R14079 GND.n1053 GND.n1052 9.3005
R14080 GND.n5662 GND.n5661 9.3005
R14081 GND.n5663 GND.n1051 9.3005
R14082 GND.n5665 GND.n5664 9.3005
R14083 GND.n1047 GND.n1046 9.3005
R14084 GND.n5672 GND.n5671 9.3005
R14085 GND.n5673 GND.n1045 9.3005
R14086 GND.n5675 GND.n5674 9.3005
R14087 GND.n1041 GND.n1040 9.3005
R14088 GND.n5682 GND.n5681 9.3005
R14089 GND.n5683 GND.n1039 9.3005
R14090 GND.n5685 GND.n5684 9.3005
R14091 GND.n1035 GND.n1034 9.3005
R14092 GND.n5692 GND.n5691 9.3005
R14093 GND.n5693 GND.n1033 9.3005
R14094 GND.n5695 GND.n5694 9.3005
R14095 GND.n1029 GND.n1028 9.3005
R14096 GND.n5702 GND.n5701 9.3005
R14097 GND.n5703 GND.n1027 9.3005
R14098 GND.n5705 GND.n5704 9.3005
R14099 GND.n1023 GND.n1022 9.3005
R14100 GND.n5712 GND.n5711 9.3005
R14101 GND.n5713 GND.n1021 9.3005
R14102 GND.n5715 GND.n5714 9.3005
R14103 GND.n1017 GND.n1016 9.3005
R14104 GND.n5722 GND.n5721 9.3005
R14105 GND.n5723 GND.n1015 9.3005
R14106 GND.n5725 GND.n5724 9.3005
R14107 GND.n1011 GND.n1010 9.3005
R14108 GND.n5732 GND.n5731 9.3005
R14109 GND.n5733 GND.n1009 9.3005
R14110 GND.n5735 GND.n5734 9.3005
R14111 GND.n1005 GND.n1004 9.3005
R14112 GND.n5742 GND.n5741 9.3005
R14113 GND.n5743 GND.n1003 9.3005
R14114 GND.n5745 GND.n5744 9.3005
R14115 GND.n999 GND.n998 9.3005
R14116 GND.n5752 GND.n5751 9.3005
R14117 GND.n5753 GND.n997 9.3005
R14118 GND.n5755 GND.n5754 9.3005
R14119 GND.n993 GND.n992 9.3005
R14120 GND.n5762 GND.n5761 9.3005
R14121 GND.n5763 GND.n991 9.3005
R14122 GND.n5765 GND.n5764 9.3005
R14123 GND.n987 GND.n986 9.3005
R14124 GND.n5772 GND.n5771 9.3005
R14125 GND.n5773 GND.n985 9.3005
R14126 GND.n5775 GND.n5774 9.3005
R14127 GND.n981 GND.n980 9.3005
R14128 GND.n5782 GND.n5781 9.3005
R14129 GND.n5783 GND.n979 9.3005
R14130 GND.n5785 GND.n5784 9.3005
R14131 GND.n975 GND.n974 9.3005
R14132 GND.n5792 GND.n5791 9.3005
R14133 GND.n5793 GND.n973 9.3005
R14134 GND.n5795 GND.n5794 9.3005
R14135 GND.n969 GND.n968 9.3005
R14136 GND.n5802 GND.n5801 9.3005
R14137 GND.n5803 GND.n967 9.3005
R14138 GND.n5805 GND.n5804 9.3005
R14139 GND.n963 GND.n962 9.3005
R14140 GND.n5812 GND.n5811 9.3005
R14141 GND.n5813 GND.n961 9.3005
R14142 GND.n5815 GND.n5814 9.3005
R14143 GND.n957 GND.n956 9.3005
R14144 GND.n5822 GND.n5821 9.3005
R14145 GND.n5823 GND.n955 9.3005
R14146 GND.n5825 GND.n5824 9.3005
R14147 GND.n951 GND.n950 9.3005
R14148 GND.n5832 GND.n5831 9.3005
R14149 GND.n5833 GND.n949 9.3005
R14150 GND.n5835 GND.n5834 9.3005
R14151 GND.n945 GND.n944 9.3005
R14152 GND.n5842 GND.n5841 9.3005
R14153 GND.n5843 GND.n943 9.3005
R14154 GND.n5845 GND.n5844 9.3005
R14155 GND.n939 GND.n938 9.3005
R14156 GND.n5852 GND.n5851 9.3005
R14157 GND.n5853 GND.n937 9.3005
R14158 GND.n5855 GND.n5854 9.3005
R14159 GND.n933 GND.n932 9.3005
R14160 GND.n5862 GND.n5861 9.3005
R14161 GND.n5863 GND.n931 9.3005
R14162 GND.n5865 GND.n5864 9.3005
R14163 GND.n927 GND.n926 9.3005
R14164 GND.n5872 GND.n5871 9.3005
R14165 GND.n5873 GND.n925 9.3005
R14166 GND.n5875 GND.n5874 9.3005
R14167 GND.n921 GND.n920 9.3005
R14168 GND.n5882 GND.n5881 9.3005
R14169 GND.n5883 GND.n919 9.3005
R14170 GND.n5885 GND.n5884 9.3005
R14171 GND.n915 GND.n914 9.3005
R14172 GND.n5892 GND.n5891 9.3005
R14173 GND.n5893 GND.n913 9.3005
R14174 GND.n5895 GND.n5894 9.3005
R14175 GND.n909 GND.n908 9.3005
R14176 GND.n5902 GND.n5901 9.3005
R14177 GND.n5903 GND.n907 9.3005
R14178 GND.n5905 GND.n5904 9.3005
R14179 GND.n903 GND.n902 9.3005
R14180 GND.n5912 GND.n5911 9.3005
R14181 GND.n5913 GND.n901 9.3005
R14182 GND.n5915 GND.n5914 9.3005
R14183 GND.n897 GND.n896 9.3005
R14184 GND.n5922 GND.n5921 9.3005
R14185 GND.n5923 GND.n895 9.3005
R14186 GND.n5925 GND.n5924 9.3005
R14187 GND.n891 GND.n890 9.3005
R14188 GND.n5932 GND.n5931 9.3005
R14189 GND.n5933 GND.n889 9.3005
R14190 GND.n5935 GND.n5934 9.3005
R14191 GND.n885 GND.n884 9.3005
R14192 GND.n5942 GND.n5941 9.3005
R14193 GND.n5943 GND.n883 9.3005
R14194 GND.n5945 GND.n5944 9.3005
R14195 GND.n879 GND.n878 9.3005
R14196 GND.n5952 GND.n5951 9.3005
R14197 GND.n5953 GND.n877 9.3005
R14198 GND.n5955 GND.n5954 9.3005
R14199 GND.n873 GND.n872 9.3005
R14200 GND.n5962 GND.n5961 9.3005
R14201 GND.n5963 GND.n871 9.3005
R14202 GND.n5965 GND.n5964 9.3005
R14203 GND.n867 GND.n866 9.3005
R14204 GND.n5972 GND.n5971 9.3005
R14205 GND.n5973 GND.n865 9.3005
R14206 GND.n5975 GND.n5974 9.3005
R14207 GND.n861 GND.n860 9.3005
R14208 GND.n5982 GND.n5981 9.3005
R14209 GND.n5983 GND.n859 9.3005
R14210 GND.n5985 GND.n5984 9.3005
R14211 GND.n855 GND.n854 9.3005
R14212 GND.n5992 GND.n5991 9.3005
R14213 GND.n5993 GND.n853 9.3005
R14214 GND.n5995 GND.n5994 9.3005
R14215 GND.n849 GND.n848 9.3005
R14216 GND.n6002 GND.n6001 9.3005
R14217 GND.n6003 GND.n847 9.3005
R14218 GND.n6005 GND.n6004 9.3005
R14219 GND.n843 GND.n842 9.3005
R14220 GND.n6012 GND.n6011 9.3005
R14221 GND.n6013 GND.n841 9.3005
R14222 GND.n6015 GND.n6014 9.3005
R14223 GND.n837 GND.n836 9.3005
R14224 GND.n6022 GND.n6021 9.3005
R14225 GND.n6023 GND.n835 9.3005
R14226 GND.n6025 GND.n6024 9.3005
R14227 GND.n831 GND.n830 9.3005
R14228 GND.n6032 GND.n6031 9.3005
R14229 GND.n6033 GND.n829 9.3005
R14230 GND.n6035 GND.n6034 9.3005
R14231 GND.n825 GND.n824 9.3005
R14232 GND.n6042 GND.n6041 9.3005
R14233 GND.n6043 GND.n823 9.3005
R14234 GND.n6045 GND.n6044 9.3005
R14235 GND.n819 GND.n818 9.3005
R14236 GND.n6052 GND.n6051 9.3005
R14237 GND.n6053 GND.n817 9.3005
R14238 GND.n6055 GND.n6054 9.3005
R14239 GND.n813 GND.n812 9.3005
R14240 GND.n6062 GND.n6061 9.3005
R14241 GND.n6063 GND.n811 9.3005
R14242 GND.n6065 GND.n6064 9.3005
R14243 GND.n807 GND.n806 9.3005
R14244 GND.n6072 GND.n6071 9.3005
R14245 GND.n6073 GND.n805 9.3005
R14246 GND.n6075 GND.n6074 9.3005
R14247 GND.n801 GND.n800 9.3005
R14248 GND.n6082 GND.n6081 9.3005
R14249 GND.n6083 GND.n799 9.3005
R14250 GND.n6085 GND.n6084 9.3005
R14251 GND.n795 GND.n794 9.3005
R14252 GND.n6092 GND.n6091 9.3005
R14253 GND.n6093 GND.n793 9.3005
R14254 GND.n6095 GND.n6094 9.3005
R14255 GND.n789 GND.n788 9.3005
R14256 GND.n6102 GND.n6101 9.3005
R14257 GND.n6103 GND.n787 9.3005
R14258 GND.n6105 GND.n6104 9.3005
R14259 GND.n783 GND.n782 9.3005
R14260 GND.n6112 GND.n6111 9.3005
R14261 GND.n6113 GND.n781 9.3005
R14262 GND.n6115 GND.n6114 9.3005
R14263 GND.n777 GND.n776 9.3005
R14264 GND.n6122 GND.n6121 9.3005
R14265 GND.n6123 GND.n775 9.3005
R14266 GND.n6125 GND.n6124 9.3005
R14267 GND.n771 GND.n770 9.3005
R14268 GND.n6132 GND.n6131 9.3005
R14269 GND.n6133 GND.n769 9.3005
R14270 GND.n6135 GND.n6134 9.3005
R14271 GND.n765 GND.n764 9.3005
R14272 GND.n6142 GND.n6141 9.3005
R14273 GND.n6143 GND.n763 9.3005
R14274 GND.n6145 GND.n6144 9.3005
R14275 GND.n759 GND.n758 9.3005
R14276 GND.n6152 GND.n6151 9.3005
R14277 GND.n6153 GND.n757 9.3005
R14278 GND.n6155 GND.n6154 9.3005
R14279 GND.n753 GND.n752 9.3005
R14280 GND.n6162 GND.n6161 9.3005
R14281 GND.n6163 GND.n751 9.3005
R14282 GND.n6165 GND.n6164 9.3005
R14283 GND.n747 GND.n746 9.3005
R14284 GND.n6172 GND.n6171 9.3005
R14285 GND.n6173 GND.n745 9.3005
R14286 GND.n6175 GND.n6174 9.3005
R14287 GND.n741 GND.n740 9.3005
R14288 GND.n6182 GND.n6181 9.3005
R14289 GND.n6183 GND.n739 9.3005
R14290 GND.n6185 GND.n6184 9.3005
R14291 GND.n6192 GND.n6191 9.3005
R14292 GND.n6193 GND.n733 9.3005
R14293 GND.n6195 GND.n6194 9.3005
R14294 GND.n729 GND.n728 9.3005
R14295 GND.n6202 GND.n6201 9.3005
R14296 GND.n6203 GND.n727 9.3005
R14297 GND.n6205 GND.n6204 9.3005
R14298 GND.n723 GND.n722 9.3005
R14299 GND.n6212 GND.n6211 9.3005
R14300 GND.n6213 GND.n721 9.3005
R14301 GND.n6215 GND.n6214 9.3005
R14302 GND.n717 GND.n716 9.3005
R14303 GND.n6222 GND.n6221 9.3005
R14304 GND.n6223 GND.n715 9.3005
R14305 GND.n6225 GND.n6224 9.3005
R14306 GND.n711 GND.n710 9.3005
R14307 GND.n6232 GND.n6231 9.3005
R14308 GND.n6233 GND.n709 9.3005
R14309 GND.n6235 GND.n6234 9.3005
R14310 GND.n705 GND.n704 9.3005
R14311 GND.n6242 GND.n6241 9.3005
R14312 GND.n6243 GND.n703 9.3005
R14313 GND.n6245 GND.n6244 9.3005
R14314 GND.n699 GND.n698 9.3005
R14315 GND.n6252 GND.n6251 9.3005
R14316 GND.n6253 GND.n697 9.3005
R14317 GND.n6255 GND.n6254 9.3005
R14318 GND.n693 GND.n692 9.3005
R14319 GND.n6262 GND.n6261 9.3005
R14320 GND.n6263 GND.n691 9.3005
R14321 GND.n6265 GND.n6264 9.3005
R14322 GND.n687 GND.n686 9.3005
R14323 GND.n6272 GND.n6271 9.3005
R14324 GND.n6273 GND.n685 9.3005
R14325 GND.n6275 GND.n6274 9.3005
R14326 GND.n681 GND.n680 9.3005
R14327 GND.n6282 GND.n6281 9.3005
R14328 GND.n6283 GND.n679 9.3005
R14329 GND.n6285 GND.n6284 9.3005
R14330 GND.n675 GND.n674 9.3005
R14331 GND.n6292 GND.n6291 9.3005
R14332 GND.n6293 GND.n673 9.3005
R14333 GND.n6295 GND.n6294 9.3005
R14334 GND.n669 GND.n668 9.3005
R14335 GND.n6302 GND.n6301 9.3005
R14336 GND.n6303 GND.n667 9.3005
R14337 GND.n6307 GND.n6304 9.3005
R14338 GND.n6306 GND.n6305 9.3005
R14339 GND.n735 GND.n734 9.3005
R14340 GND.n307 GND.n306 9.3005
R14341 GND.n300 GND.n299 9.3005
R14342 GND.n294 GND.n293 9.3005
R14343 GND.n287 GND.n286 9.3005
R14344 GND.n281 GND.n280 9.3005
R14345 GND.n274 GND.n273 9.3005
R14346 GND.n268 GND.n267 9.3005
R14347 GND.n261 GND.n260 9.3005
R14348 GND.n255 GND.n254 9.3005
R14349 GND.n248 GND.n247 9.3005
R14350 GND.n242 GND.n241 9.3005
R14351 GND.n235 GND.n234 9.3005
R14352 GND.n229 GND.n228 9.3005
R14353 GND.n222 GND.n221 9.3005
R14354 GND.n216 GND.n215 9.3005
R14355 GND.n209 GND.n208 9.3005
R14356 GND.n203 GND.n202 9.3005
R14357 GND.n196 GND.n195 9.3005
R14358 GND.n190 GND.n189 9.3005
R14359 GND.n183 GND.n182 9.3005
R14360 GND.n178 GND.n177 9.3005
R14361 GND.n171 GND.n170 9.3005
R14362 GND.n165 GND.n164 9.3005
R14363 GND.n158 GND.n157 9.3005
R14364 GND.n4532 GND.n2901 9.3005
R14365 GND.n4536 GND.n4533 9.3005
R14366 GND.n4537 GND.n2900 9.3005
R14367 GND.n4554 GND.n4553 9.3005
R14368 GND.n4555 GND.n2899 9.3005
R14369 GND.n4557 GND.n4556 9.3005
R14370 GND.n2897 GND.n2896 9.3005
R14371 GND.n4569 GND.n4568 9.3005
R14372 GND.n4570 GND.n2895 9.3005
R14373 GND.n4572 GND.n4571 9.3005
R14374 GND.n2893 GND.n2892 9.3005
R14375 GND.n4584 GND.n4583 9.3005
R14376 GND.n4585 GND.n2891 9.3005
R14377 GND.n4587 GND.n4586 9.3005
R14378 GND.n2889 GND.n2888 9.3005
R14379 GND.n4599 GND.n4598 9.3005
R14380 GND.n4600 GND.n2887 9.3005
R14381 GND.n4602 GND.n4601 9.3005
R14382 GND.n2885 GND.n2884 9.3005
R14383 GND.n4614 GND.n4613 9.3005
R14384 GND.n4615 GND.n2883 9.3005
R14385 GND.n4621 GND.n4616 9.3005
R14386 GND.n4620 GND.n4617 9.3005
R14387 GND.n4619 GND.n4618 9.3005
R14388 GND.n313 GND.n311 9.3005
R14389 GND.n4531 GND.n4530 9.3005
R14390 GND.n6427 GND.n6426 9.3005
R14391 GND.n314 GND.n312 9.3005
R14392 GND.n4639 GND.n4638 9.3005
R14393 GND.n4772 GND.n4640 9.3005
R14394 GND.n4771 GND.n4641 9.3005
R14395 GND.n4770 GND.n4642 9.3005
R14396 GND.n4646 GND.n4643 9.3005
R14397 GND.n4760 GND.n4647 9.3005
R14398 GND.n4759 GND.n4648 9.3005
R14399 GND.n4758 GND.n4649 9.3005
R14400 GND.n4653 GND.n4650 9.3005
R14401 GND.n4748 GND.n4654 9.3005
R14402 GND.n4747 GND.n4655 9.3005
R14403 GND.n4746 GND.n4656 9.3005
R14404 GND.n4660 GND.n4657 9.3005
R14405 GND.n4736 GND.n4661 9.3005
R14406 GND.n4735 GND.n4662 9.3005
R14407 GND.n4734 GND.n4663 9.3005
R14408 GND.n4667 GND.n4664 9.3005
R14409 GND.n4724 GND.n4668 9.3005
R14410 GND.n4723 GND.n4669 9.3005
R14411 GND.n4722 GND.n4670 9.3005
R14412 GND.n4673 GND.n4671 9.3005
R14413 GND.n4712 GND.n4674 9.3005
R14414 GND.n4711 GND.n4675 9.3005
R14415 GND.n4710 GND.n4709 9.3005
R14416 GND.n4690 GND.n4685 9.3005
R14417 GND.n4692 GND.n4691 9.3005
R14418 GND.n4683 GND.n4682 9.3005
R14419 GND.n4699 GND.n4698 9.3005
R14420 GND.n4700 GND.n4681 9.3005
R14421 GND.n4702 GND.n4701 9.3005
R14422 GND.n4679 GND.n4676 9.3005
R14423 GND.n4708 GND.n4707 9.3005
R14424 GND.n4689 GND.n4688 9.3005
R14425 GND.n527 GND.n526 9.3005
R14426 GND.n530 GND.n521 9.3005
R14427 GND.n534 GND.n533 9.3005
R14428 GND.n535 GND.n520 9.3005
R14429 GND.n537 GND.n536 9.3005
R14430 GND.n540 GND.n515 9.3005
R14431 GND.n542 GND.n541 9.3005
R14432 GND.n543 GND.n514 9.3005
R14433 GND.n545 GND.n544 9.3005
R14434 GND.n548 GND.n513 9.3005
R14435 GND.n552 GND.n551 9.3005
R14436 GND.n553 GND.n512 9.3005
R14437 GND.n555 GND.n554 9.3005
R14438 GND.n558 GND.n511 9.3005
R14439 GND.n562 GND.n561 9.3005
R14440 GND.n563 GND.n510 9.3005
R14441 GND.n565 GND.n564 9.3005
R14442 GND.n568 GND.n507 9.3005
R14443 GND.n572 GND.n571 9.3005
R14444 GND.n573 GND.n506 9.3005
R14445 GND.n575 GND.n574 9.3005
R14446 GND.n578 GND.n505 9.3005
R14447 GND.n582 GND.n581 9.3005
R14448 GND.n583 GND.n504 9.3005
R14449 GND.n585 GND.n584 9.3005
R14450 GND.n588 GND.n503 9.3005
R14451 GND.n589 GND.n499 9.3005
R14452 GND.n593 GND.n592 9.3005
R14453 GND.n594 GND.n498 9.3005
R14454 GND.n598 GND.n595 9.3005
R14455 GND.n599 GND.n497 9.3005
R14456 GND.n603 GND.n602 9.3005
R14457 GND.n604 GND.n496 9.3005
R14458 GND.n608 GND.n605 9.3005
R14459 GND.n609 GND.n495 9.3005
R14460 GND.n612 GND.n492 9.3005
R14461 GND.n616 GND.n615 9.3005
R14462 GND.n617 GND.n491 9.3005
R14463 GND.n619 GND.n618 9.3005
R14464 GND.n622 GND.n490 9.3005
R14465 GND.n626 GND.n625 9.3005
R14466 GND.n627 GND.n489 9.3005
R14467 GND.n629 GND.n628 9.3005
R14468 GND.n630 GND.n488 9.3005
R14469 GND.n487 GND.n484 9.3005
R14470 GND.n525 GND.n523 9.3005
R14471 GND.n4542 GND.n2609 9.3005
R14472 GND.n4545 GND.n4541 9.3005
R14473 GND.n4547 GND.n4546 9.3005
R14474 GND.n4548 GND.n2649 9.3005
R14475 GND.n4848 GND.n2650 9.3005
R14476 GND.n4847 GND.n2651 9.3005
R14477 GND.n4846 GND.n2652 9.3005
R14478 GND.n4563 GND.n2653 9.3005
R14479 GND.n4836 GND.n2671 9.3005
R14480 GND.n4835 GND.n2672 9.3005
R14481 GND.n4834 GND.n2673 9.3005
R14482 GND.n4578 GND.n2674 9.3005
R14483 GND.n4824 GND.n2692 9.3005
R14484 GND.n4823 GND.n2693 9.3005
R14485 GND.n4822 GND.n2694 9.3005
R14486 GND.n4593 GND.n2695 9.3005
R14487 GND.n4812 GND.n2713 9.3005
R14488 GND.n4811 GND.n2714 9.3005
R14489 GND.n4810 GND.n2715 9.3005
R14490 GND.n4608 GND.n2716 9.3005
R14491 GND.n4800 GND.n2732 9.3005
R14492 GND.n4799 GND.n2733 9.3005
R14493 GND.n4798 GND.n2734 9.3005
R14494 GND.n4628 GND.n2735 9.3005
R14495 GND.n4631 GND.n4629 9.3005
R14496 GND.n4633 GND.n4632 9.3005
R14497 GND.n2878 GND.n2877 9.3005
R14498 GND.n4779 GND.n4778 9.3005
R14499 GND.n2879 GND.n342 9.3005
R14500 GND.n6415 GND.n343 9.3005
R14501 GND.n6414 GND.n344 9.3005
R14502 GND.n6413 GND.n345 9.3005
R14503 GND.n4644 GND.n346 9.3005
R14504 GND.n6403 GND.n363 9.3005
R14505 GND.n6402 GND.n364 9.3005
R14506 GND.n6401 GND.n365 9.3005
R14507 GND.n4651 GND.n366 9.3005
R14508 GND.n6391 GND.n384 9.3005
R14509 GND.n6390 GND.n385 9.3005
R14510 GND.n6389 GND.n386 9.3005
R14511 GND.n4658 GND.n387 9.3005
R14512 GND.n6379 GND.n405 9.3005
R14513 GND.n6378 GND.n406 9.3005
R14514 GND.n6377 GND.n407 9.3005
R14515 GND.n4665 GND.n408 9.3005
R14516 GND.n6367 GND.n426 9.3005
R14517 GND.n6366 GND.n427 9.3005
R14518 GND.n6365 GND.n428 9.3005
R14519 GND.n4672 GND.n429 9.3005
R14520 GND.n6355 GND.n447 9.3005
R14521 GND.n6354 GND.n6353 9.3005
R14522 GND.n4867 GND.n2608 9.3005
R14523 GND.n2610 GND.n2609 9.3005
R14524 GND.n4541 GND.n4540 9.3005
R14525 GND.n4547 GND.n4538 9.3005
R14526 GND.n4549 GND.n4548 9.3005
R14527 GND.n2898 GND.n2650 9.3005
R14528 GND.n4561 GND.n2651 9.3005
R14529 GND.n4562 GND.n2652 9.3005
R14530 GND.n4564 GND.n4563 9.3005
R14531 GND.n2894 GND.n2671 9.3005
R14532 GND.n4576 GND.n2672 9.3005
R14533 GND.n4577 GND.n2673 9.3005
R14534 GND.n4579 GND.n4578 9.3005
R14535 GND.n2890 GND.n2692 9.3005
R14536 GND.n4591 GND.n2693 9.3005
R14537 GND.n4592 GND.n2694 9.3005
R14538 GND.n4594 GND.n4593 9.3005
R14539 GND.n2886 GND.n2713 9.3005
R14540 GND.n4606 GND.n2714 9.3005
R14541 GND.n4607 GND.n2715 9.3005
R14542 GND.n4609 GND.n4608 9.3005
R14543 GND.n2882 GND.n2732 9.3005
R14544 GND.n4625 GND.n2733 9.3005
R14545 GND.n4626 GND.n2734 9.3005
R14546 GND.n4628 GND.n4627 9.3005
R14547 GND.n4629 GND.n2881 9.3005
R14548 GND.n4634 GND.n4633 9.3005
R14549 GND.n4636 GND.n2878 9.3005
R14550 GND.n4778 GND.n4777 9.3005
R14551 GND.n4776 GND.n2879 9.3005
R14552 GND.n4637 GND.n343 9.3005
R14553 GND.n4766 GND.n344 9.3005
R14554 GND.n4765 GND.n345 9.3005
R14555 GND.n4764 GND.n4644 9.3005
R14556 GND.n4645 GND.n363 9.3005
R14557 GND.n4754 GND.n364 9.3005
R14558 GND.n4753 GND.n365 9.3005
R14559 GND.n4752 GND.n4651 9.3005
R14560 GND.n4652 GND.n384 9.3005
R14561 GND.n4742 GND.n385 9.3005
R14562 GND.n4741 GND.n386 9.3005
R14563 GND.n4740 GND.n4658 9.3005
R14564 GND.n4659 GND.n405 9.3005
R14565 GND.n4730 GND.n406 9.3005
R14566 GND.n4729 GND.n407 9.3005
R14567 GND.n4728 GND.n4665 9.3005
R14568 GND.n4666 GND.n426 9.3005
R14569 GND.n4718 GND.n427 9.3005
R14570 GND.n4717 GND.n428 9.3005
R14571 GND.n4716 GND.n4672 9.3005
R14572 GND.n449 GND.n447 9.3005
R14573 GND.n6353 GND.n6352 9.3005
R14574 GND.n4867 GND.n4866 9.3005
R14575 GND.n4873 GND.n4872 9.3005
R14576 GND.n4876 GND.n2603 9.3005
R14577 GND.n4877 GND.n2602 9.3005
R14578 GND.n4880 GND.n2601 9.3005
R14579 GND.n4881 GND.n2600 9.3005
R14580 GND.n4884 GND.n2599 9.3005
R14581 GND.n4885 GND.n2598 9.3005
R14582 GND.n4888 GND.n2597 9.3005
R14583 GND.n4889 GND.n2594 9.3005
R14584 GND.n4892 GND.n2593 9.3005
R14585 GND.n4893 GND.n2592 9.3005
R14586 GND.n4896 GND.n2591 9.3005
R14587 GND.n4897 GND.n2590 9.3005
R14588 GND.n4900 GND.n2589 9.3005
R14589 GND.n4901 GND.n2588 9.3005
R14590 GND.n4904 GND.n2587 9.3005
R14591 GND.n4905 GND.n2586 9.3005
R14592 GND.n4908 GND.n2585 9.3005
R14593 GND.n4910 GND.n2582 9.3005
R14594 GND.n4913 GND.n2581 9.3005
R14595 GND.n4914 GND.n2580 9.3005
R14596 GND.n4917 GND.n2579 9.3005
R14597 GND.n4919 GND.n2575 9.3005
R14598 GND.n4922 GND.n2574 9.3005
R14599 GND.n4924 GND.n2573 9.3005
R14600 GND.n4926 GND.n2568 9.3005
R14601 GND.n4929 GND.n2567 9.3005
R14602 GND.n4930 GND.n2566 9.3005
R14603 GND.n4933 GND.n2565 9.3005
R14604 GND.n4934 GND.n2564 9.3005
R14605 GND.n4937 GND.n2563 9.3005
R14606 GND.n4938 GND.n2562 9.3005
R14607 GND.n4941 GND.n2561 9.3005
R14608 GND.n4942 GND.n2558 9.3005
R14609 GND.n4945 GND.n2557 9.3005
R14610 GND.n4946 GND.n2556 9.3005
R14611 GND.n4949 GND.n2555 9.3005
R14612 GND.n4951 GND.n2554 9.3005
R14613 GND.n4952 GND.n2553 9.3005
R14614 GND.n4953 GND.n2552 9.3005
R14615 GND.n4954 GND.n2551 9.3005
R14616 GND.n4925 GND.n2570 9.3005
R14617 GND.n4871 GND.n2607 9.3005
R14618 GND.n4870 GND.n4869 9.3005
R14619 GND.n2636 GND.n2635 9.3005
R14620 GND.n2637 GND.n2631 9.3005
R14621 GND.n4854 GND.n2638 9.3005
R14622 GND.n4853 GND.n2639 9.3005
R14623 GND.n4852 GND.n2640 9.3005
R14624 GND.n2660 GND.n2641 9.3005
R14625 GND.n4842 GND.n2661 9.3005
R14626 GND.n4841 GND.n2662 9.3005
R14627 GND.n4840 GND.n2663 9.3005
R14628 GND.n2681 GND.n2664 9.3005
R14629 GND.n4830 GND.n2682 9.3005
R14630 GND.n4829 GND.n2683 9.3005
R14631 GND.n4828 GND.n2684 9.3005
R14632 GND.n2702 GND.n2685 9.3005
R14633 GND.n4818 GND.n2703 9.3005
R14634 GND.n4817 GND.n2704 9.3005
R14635 GND.n4816 GND.n2705 9.3005
R14636 GND.n2723 GND.n2706 9.3005
R14637 GND.n4806 GND.n2724 9.3005
R14638 GND.n4805 GND.n326 9.3005
R14639 GND.n333 GND.n325 9.3005
R14640 GND.n6409 GND.n353 9.3005
R14641 GND.n6408 GND.n354 9.3005
R14642 GND.n6407 GND.n355 9.3005
R14643 GND.n373 GND.n356 9.3005
R14644 GND.n6397 GND.n374 9.3005
R14645 GND.n6396 GND.n375 9.3005
R14646 GND.n6395 GND.n376 9.3005
R14647 GND.n394 GND.n377 9.3005
R14648 GND.n6385 GND.n395 9.3005
R14649 GND.n6384 GND.n396 9.3005
R14650 GND.n6383 GND.n397 9.3005
R14651 GND.n415 GND.n398 9.3005
R14652 GND.n6373 GND.n416 9.3005
R14653 GND.n6372 GND.n417 9.3005
R14654 GND.n6371 GND.n418 9.3005
R14655 GND.n436 GND.n419 9.3005
R14656 GND.n6361 GND.n437 9.3005
R14657 GND.n6360 GND.n438 9.3005
R14658 GND.n6359 GND.n439 9.3005
R14659 GND.n524 GND.n440 9.3005
R14660 GND.n2633 GND.n2632 9.3005
R14661 GND.n6420 GND.n330 9.3005
R14662 GND.n6420 GND.n6419 9.3005
R14663 GND.n1931 GND.n1930 9.3005
R14664 GND.n1929 GND.n1773 9.3005
R14665 GND.n1928 GND.n1927 9.3005
R14666 GND.n1775 GND.n1774 9.3005
R14667 GND.n1921 GND.n1920 9.3005
R14668 GND.n1919 GND.n1777 9.3005
R14669 GND.n1918 GND.n1917 9.3005
R14670 GND.n1779 GND.n1778 9.3005
R14671 GND.n1911 GND.n1908 9.3005
R14672 GND.n1907 GND.n1781 9.3005
R14673 GND.n1906 GND.n1905 9.3005
R14674 GND.n1783 GND.n1782 9.3005
R14675 GND.n1899 GND.n1898 9.3005
R14676 GND.n1897 GND.n1785 9.3005
R14677 GND.n1896 GND.n1895 9.3005
R14678 GND.n1787 GND.n1786 9.3005
R14679 GND.n1889 GND.n1888 9.3005
R14680 GND.n1887 GND.n1789 9.3005
R14681 GND.n1886 GND.n1885 9.3005
R14682 GND.n1791 GND.n1790 9.3005
R14683 GND.n1879 GND.n1878 9.3005
R14684 GND.n1877 GND.n1796 9.3005
R14685 GND.n1876 GND.n1875 9.3005
R14686 GND.n1798 GND.n1797 9.3005
R14687 GND.n1869 GND.n1868 9.3005
R14688 GND.n1867 GND.n1800 9.3005
R14689 GND.n1866 GND.n1865 9.3005
R14690 GND.n1859 GND.n1858 9.3005
R14691 GND.n1857 GND.n1806 9.3005
R14692 GND.n1856 GND.n1855 9.3005
R14693 GND.n1808 GND.n1807 9.3005
R14694 GND.n1849 GND.n1848 9.3005
R14695 GND.n1847 GND.n1810 9.3005
R14696 GND.n1846 GND.n1845 9.3005
R14697 GND.n1812 GND.n1811 9.3005
R14698 GND.n1839 GND.n1836 9.3005
R14699 GND.n1835 GND.n1814 9.3005
R14700 GND.n1834 GND.n1833 9.3005
R14701 GND.n1816 GND.n1815 9.3005
R14702 GND.n1827 GND.n1826 9.3005
R14703 GND.n1825 GND.n1818 9.3005
R14704 GND.n1824 GND.n1823 9.3005
R14705 GND.n1820 GND.n1819 9.3005
R14706 GND.n1804 GND.n1801 9.3005
R14707 GND.n1771 GND.n1768 9.3005
R14708 GND.n1937 GND.n1936 9.3005
R14709 GND.n5376 GND.n1283 9.3005
R14710 GND.n5375 GND.n1284 9.3005
R14711 GND.n2006 GND.n1285 9.3005
R14712 GND.n2010 GND.n2007 9.3005
R14713 GND.n2009 GND.n2008 9.3005
R14714 GND.n1743 GND.n1742 9.3005
R14715 GND.n2030 GND.n2029 9.3005
R14716 GND.n2031 GND.n1741 9.3005
R14717 GND.n2035 GND.n2032 9.3005
R14718 GND.n2034 GND.n2033 9.3005
R14719 GND.n1713 GND.n1712 9.3005
R14720 GND.n2083 GND.n2082 9.3005
R14721 GND.n2084 GND.n1711 9.3005
R14722 GND.n2088 GND.n2085 9.3005
R14723 GND.n2087 GND.n2086 9.3005
R14724 GND.n1691 GND.n1690 9.3005
R14725 GND.n2107 GND.n2106 9.3005
R14726 GND.n2108 GND.n1689 9.3005
R14727 GND.n2110 GND.n2109 9.3005
R14728 GND.n1641 GND.n1634 9.3005
R14729 GND.n2217 GND.n2216 9.3005
R14730 GND.n1612 GND.n1611 9.3005
R14731 GND.n2237 GND.n2236 9.3005
R14732 GND.n2238 GND.n1610 9.3005
R14733 GND.n2242 GND.n2239 9.3005
R14734 GND.n2241 GND.n2240 9.3005
R14735 GND.n1589 GND.n1588 9.3005
R14736 GND.n2262 GND.n2261 9.3005
R14737 GND.n2263 GND.n1587 9.3005
R14738 GND.n2267 GND.n2264 9.3005
R14739 GND.n2266 GND.n2265 9.3005
R14740 GND.n1567 GND.n1566 9.3005
R14741 GND.n2300 GND.n2299 9.3005
R14742 GND.n2301 GND.n1565 9.3005
R14743 GND.n2303 GND.n2302 9.3005
R14744 GND.n1548 GND.n1547 9.3005
R14745 GND.n2337 GND.n2336 9.3005
R14746 GND.n2338 GND.n1546 9.3005
R14747 GND.n2340 GND.n2339 9.3005
R14748 GND.n1403 GND.n1402 9.3005
R14749 GND.n5292 GND.n5291 9.3005
R14750 GND.n5377 GND.n1282 9.3005
R14751 GND.n2215 GND.n1639 9.3005
R14752 GND.n2218 GND.n2215 9.3005
R14753 GND.n2205 GND.n1635 9.3005
R14754 GND.n2181 GND.n2147 9.3005
R14755 GND.n2180 GND.n2148 9.3005
R14756 GND.n2151 GND.n2149 9.3005
R14757 GND.n2176 GND.n2152 9.3005
R14758 GND.n2175 GND.n2153 9.3005
R14759 GND.n2174 GND.n2154 9.3005
R14760 GND.n2157 GND.n2155 9.3005
R14761 GND.n2170 GND.n2158 9.3005
R14762 GND.n2169 GND.n2159 9.3005
R14763 GND.n2168 GND.n2160 9.3005
R14764 GND.n2162 GND.n2161 9.3005
R14765 GND.n2164 GND.n2163 9.3005
R14766 GND.n1559 GND.n1558 9.3005
R14767 GND.n2309 GND.n2308 9.3005
R14768 GND.n2310 GND.n1557 9.3005
R14769 GND.n2327 GND.n2311 9.3005
R14770 GND.n2326 GND.n2312 9.3005
R14771 GND.n2325 GND.n2313 9.3005
R14772 GND.n2316 GND.n2314 9.3005
R14773 GND.n2321 GND.n2317 9.3005
R14774 GND.n2320 GND.n2319 9.3005
R14775 GND.n2318 GND.n1527 9.3005
R14776 GND.n5166 GND.n1528 9.3005
R14777 GND.n5165 GND.n1529 9.3005
R14778 GND.n5164 GND.n1530 9.3005
R14779 GND.n3514 GND.n1531 9.3005
R14780 GND.n3516 GND.n3515 9.3005
R14781 GND.n3519 GND.n3518 9.3005
R14782 GND.n3520 GND.n3513 9.3005
R14783 GND.n3522 GND.n3521 9.3005
R14784 GND.n3465 GND.n3464 9.3005
R14785 GND.n3537 GND.n3536 9.3005
R14786 GND.n3538 GND.n3463 9.3005
R14787 GND.n3540 GND.n3539 9.3005
R14788 GND.n3454 GND.n3453 9.3005
R14789 GND.n3554 GND.n3553 9.3005
R14790 GND.n3555 GND.n3452 9.3005
R14791 GND.n3557 GND.n3556 9.3005
R14792 GND.n3442 GND.n3441 9.3005
R14793 GND.n3571 GND.n3570 9.3005
R14794 GND.n3572 GND.n3440 9.3005
R14795 GND.n3574 GND.n3573 9.3005
R14796 GND.n3430 GND.n3429 9.3005
R14797 GND.n3588 GND.n3587 9.3005
R14798 GND.n3589 GND.n3428 9.3005
R14799 GND.n3591 GND.n3590 9.3005
R14800 GND.n3417 GND.n3416 9.3005
R14801 GND.n3606 GND.n3605 9.3005
R14802 GND.n3607 GND.n3415 9.3005
R14803 GND.n3609 GND.n3608 9.3005
R14804 GND.n3384 GND.n3383 9.3005
R14805 GND.n3742 GND.n3741 9.3005
R14806 GND.n3743 GND.n3382 9.3005
R14807 GND.n3753 GND.n3744 9.3005
R14808 GND.n3752 GND.n3745 9.3005
R14809 GND.n3751 GND.n3746 9.3005
R14810 GND.n3748 GND.n3747 9.3005
R14811 GND.n3346 GND.n3345 9.3005
R14812 GND.n3788 GND.n3787 9.3005
R14813 GND.n3789 GND.n3344 9.3005
R14814 GND.n3793 GND.n3790 9.3005
R14815 GND.n3792 GND.n3791 9.3005
R14816 GND.n3317 GND.n3316 9.3005
R14817 GND.n3842 GND.n3841 9.3005
R14818 GND.n3843 GND.n3315 9.3005
R14819 GND.n3847 GND.n3844 9.3005
R14820 GND.n3846 GND.n3845 9.3005
R14821 GND.n3293 GND.n3292 9.3005
R14822 GND.n3903 GND.n3902 9.3005
R14823 GND.n3904 GND.n3291 9.3005
R14824 GND.n3914 GND.n3905 9.3005
R14825 GND.n3913 GND.n3906 9.3005
R14826 GND.n3912 GND.n3907 9.3005
R14827 GND.n3909 GND.n3908 9.3005
R14828 GND.n3258 GND.n3257 9.3005
R14829 GND.n3949 GND.n3948 9.3005
R14830 GND.n3950 GND.n3256 9.3005
R14831 GND.n3954 GND.n3951 9.3005
R14832 GND.n3953 GND.n3952 9.3005
R14833 GND.n3230 GND.n3229 9.3005
R14834 GND.n4002 GND.n4001 9.3005
R14835 GND.n4003 GND.n3228 9.3005
R14836 GND.n4007 GND.n4004 9.3005
R14837 GND.n4006 GND.n4005 9.3005
R14838 GND.n3205 GND.n3204 9.3005
R14839 GND.n4063 GND.n4062 9.3005
R14840 GND.n4064 GND.n3203 9.3005
R14841 GND.n4074 GND.n4065 9.3005
R14842 GND.n4073 GND.n4066 9.3005
R14843 GND.n4072 GND.n4067 9.3005
R14844 GND.n4069 GND.n4068 9.3005
R14845 GND.n3172 GND.n3171 9.3005
R14846 GND.n4109 GND.n4108 9.3005
R14847 GND.n4110 GND.n3170 9.3005
R14848 GND.n4114 GND.n4111 9.3005
R14849 GND.n4113 GND.n4112 9.3005
R14850 GND.n3143 GND.n3142 9.3005
R14851 GND.n4162 GND.n4161 9.3005
R14852 GND.n4163 GND.n3141 9.3005
R14853 GND.n4167 GND.n4164 9.3005
R14854 GND.n4166 GND.n4165 9.3005
R14855 GND.n3118 GND.n3117 9.3005
R14856 GND.n4210 GND.n4209 9.3005
R14857 GND.n4211 GND.n3116 9.3005
R14858 GND.n4224 GND.n4212 9.3005
R14859 GND.n4223 GND.n4213 9.3005
R14860 GND.n4222 GND.n4214 9.3005
R14861 GND.n4216 GND.n4215 9.3005
R14862 GND.n4218 GND.n4217 9.3005
R14863 GND.n3077 GND.n3076 9.3005
R14864 GND.n4324 GND.n4323 9.3005
R14865 GND.n4325 GND.n3075 9.3005
R14866 GND.n4329 GND.n4326 9.3005
R14867 GND.n4328 GND.n4327 9.3005
R14868 GND.n3027 GND.n3026 9.3005
R14869 GND.n4393 GND.n4392 9.3005
R14870 GND.n4394 GND.n3025 9.3005
R14871 GND.n4396 GND.n4395 9.3005
R14872 GND.n3015 GND.n3014 9.3005
R14873 GND.n4410 GND.n4409 9.3005
R14874 GND.n4411 GND.n3013 9.3005
R14875 GND.n4413 GND.n4412 9.3005
R14876 GND.n3003 GND.n3002 9.3005
R14877 GND.n4427 GND.n4426 9.3005
R14878 GND.n4428 GND.n3001 9.3005
R14879 GND.n4430 GND.n4429 9.3005
R14880 GND.n2991 GND.n2990 9.3005
R14881 GND.n4444 GND.n4443 9.3005
R14882 GND.n4445 GND.n2989 9.3005
R14883 GND.n4447 GND.n4446 9.3005
R14884 GND.n2979 GND.n2978 9.3005
R14885 GND.n4461 GND.n4460 9.3005
R14886 GND.n4462 GND.n2977 9.3005
R14887 GND.n4464 GND.n4463 9.3005
R14888 GND.n2967 GND.n2966 9.3005
R14889 GND.n4478 GND.n4477 9.3005
R14890 GND.n4479 GND.n2965 9.3005
R14891 GND.n4484 GND.n4480 9.3005
R14892 GND.n4483 GND.n4482 9.3005
R14893 GND.n4481 GND.n2955 9.3005
R14894 GND.n4498 GND.n2954 9.3005
R14895 GND.n4500 GND.n4499 9.3005
R14896 GND.n4501 GND.n2953 9.3005
R14897 GND.n4512 GND.n4502 9.3005
R14898 GND.n4511 GND.n4503 9.3005
R14899 GND.n4510 GND.n4504 9.3005
R14900 GND.n4507 GND.n4506 9.3005
R14901 GND.n4505 GND.n2617 9.3005
R14902 GND.n4861 GND.n2618 9.3005
R14903 GND.n4860 GND.n2619 9.3005
R14904 GND.n4859 GND.n2620 9.3005
R14905 GND.n2765 GND.n2621 9.3005
R14906 GND.n2766 GND.n2764 9.3005
R14907 GND.n2768 GND.n2767 9.3005
R14908 GND.n2762 GND.n2761 9.3005
R14909 GND.n2773 GND.n2772 9.3005
R14910 GND.n2774 GND.n2760 9.3005
R14911 GND.n2776 GND.n2775 9.3005
R14912 GND.n2758 GND.n2757 9.3005
R14913 GND.n2781 GND.n2780 9.3005
R14914 GND.n2782 GND.n2756 9.3005
R14915 GND.n2784 GND.n2783 9.3005
R14916 GND.n2754 GND.n2753 9.3005
R14917 GND.n2789 GND.n2788 9.3005
R14918 GND.n2790 GND.n2752 9.3005
R14919 GND.n2793 GND.n2792 9.3005
R14920 GND.n2791 GND.n2749 9.3005
R14921 GND.n2797 GND.n2750 9.3005
R14922 GND.n2798 GND.n327 9.3005
R14923 GND.n2810 GND.n2808 9.3005
R14924 GND.n2863 GND.n2811 9.3005
R14925 GND.n2862 GND.n2812 9.3005
R14926 GND.n2861 GND.n2813 9.3005
R14927 GND.n2816 GND.n2814 9.3005
R14928 GND.n2857 GND.n2817 9.3005
R14929 GND.n2856 GND.n2818 9.3005
R14930 GND.n2855 GND.n2819 9.3005
R14931 GND.n2822 GND.n2820 9.3005
R14932 GND.n2851 GND.n2823 9.3005
R14933 GND.n2850 GND.n2824 9.3005
R14934 GND.n2849 GND.n2825 9.3005
R14935 GND.n2828 GND.n2826 9.3005
R14936 GND.n2845 GND.n2829 9.3005
R14937 GND.n2844 GND.n2830 9.3005
R14938 GND.n2843 GND.n2831 9.3005
R14939 GND.n2834 GND.n2832 9.3005
R14940 GND.n2839 GND.n2835 9.3005
R14941 GND.n2838 GND.n2837 9.3005
R14942 GND.n2836 GND.n455 9.3005
R14943 GND.n6347 GND.n456 9.3005
R14944 GND.n6346 GND.n457 9.3005
R14945 GND.n6345 GND.n458 9.3005
R14946 GND.n636 GND.n459 9.3005
R14947 GND.n6339 GND.n637 9.3005
R14948 GND.n6338 GND.n638 9.3005
R14949 GND.n6337 GND.n639 9.3005
R14950 GND.n644 GND.n640 9.3005
R14951 GND.n6331 GND.n645 9.3005
R14952 GND.n6330 GND.n646 9.3005
R14953 GND.n6329 GND.n647 9.3005
R14954 GND.n652 GND.n648 9.3005
R14955 GND.n6323 GND.n653 9.3005
R14956 GND.n6322 GND.n654 9.3005
R14957 GND.n6321 GND.n655 9.3005
R14958 GND.n660 GND.n656 9.3005
R14959 GND.n6315 GND.n661 9.3005
R14960 GND.n6314 GND.n662 9.3005
R14961 GND.n6313 GND.n663 9.3005
R14962 GND.n5415 GND.n1237 9.3005
R14963 GND.n5414 GND.n1239 9.3005
R14964 GND.n1245 GND.n1240 9.3005
R14965 GND.n5408 GND.n1246 9.3005
R14966 GND.n5407 GND.n1247 9.3005
R14967 GND.n5406 GND.n1248 9.3005
R14968 GND.n1253 GND.n1249 9.3005
R14969 GND.n5400 GND.n1254 9.3005
R14970 GND.n5399 GND.n1255 9.3005
R14971 GND.n5398 GND.n1256 9.3005
R14972 GND.n1261 GND.n1257 9.3005
R14973 GND.n5392 GND.n1262 9.3005
R14974 GND.n5391 GND.n1263 9.3005
R14975 GND.n5390 GND.n1264 9.3005
R14976 GND.n1269 GND.n1265 9.3005
R14977 GND.n5384 GND.n1270 9.3005
R14978 GND.n5383 GND.n1271 9.3005
R14979 GND.n5382 GND.n1272 9.3005
R14980 GND.n1978 GND.n1273 9.3005
R14981 GND.n1980 GND.n1979 9.3005
R14982 GND.n1984 GND.n1983 9.3005
R14983 GND.n1985 GND.n1977 9.3005
R14984 GND.n2000 GND.n1986 9.3005
R14985 GND.n1999 GND.n1987 9.3005
R14986 GND.n1998 GND.n1988 9.3005
R14987 GND.n1990 GND.n1989 9.3005
R14988 GND.n1994 GND.n1991 9.3005
R14989 GND.n1993 GND.n1992 9.3005
R14990 GND.n1725 GND.n1724 9.3005
R14991 GND.n2051 GND.n2050 9.3005
R14992 GND.n2052 GND.n1723 9.3005
R14993 GND.n2074 GND.n2053 9.3005
R14994 GND.n2073 GND.n2054 9.3005
R14995 GND.n2072 GND.n2055 9.3005
R14996 GND.n2058 GND.n2056 9.3005
R14997 GND.n2068 GND.n2059 9.3005
R14998 GND.n2067 GND.n2060 9.3005
R14999 GND.n2066 GND.n2061 9.3005
R15000 GND.n5417 GND.n5416 9.3005
R15001 GND.n1236 GND.n1232 9.3005
R15002 GND.n5425 GND.n1231 9.3005
R15003 GND.n5426 GND.n1230 9.3005
R15004 GND.n5427 GND.n1229 9.3005
R15005 GND.n1228 GND.n1224 9.3005
R15006 GND.n5433 GND.n1223 9.3005
R15007 GND.n5434 GND.n1222 9.3005
R15008 GND.n5435 GND.n1221 9.3005
R15009 GND.n1220 GND.n1216 9.3005
R15010 GND.n5441 GND.n1215 9.3005
R15011 GND.n5442 GND.n1214 9.3005
R15012 GND.n5443 GND.n1213 9.3005
R15013 GND.n1212 GND.n1208 9.3005
R15014 GND.n5449 GND.n1207 9.3005
R15015 GND.n5450 GND.n1206 9.3005
R15016 GND.n5451 GND.n1205 9.3005
R15017 GND.n1204 GND.n1200 9.3005
R15018 GND.n5457 GND.n1199 9.3005
R15019 GND.n5458 GND.n1198 9.3005
R15020 GND.n5459 GND.n1197 9.3005
R15021 GND.n1196 GND.n1192 9.3005
R15022 GND.n5465 GND.n1191 9.3005
R15023 GND.n5466 GND.n1190 9.3005
R15024 GND.n5467 GND.n1189 9.3005
R15025 GND.n1188 GND.n1184 9.3005
R15026 GND.n5473 GND.n1183 9.3005
R15027 GND.n5474 GND.n1182 9.3005
R15028 GND.n5475 GND.n1181 9.3005
R15029 GND.n1180 GND.n1176 9.3005
R15030 GND.n5481 GND.n1175 9.3005
R15031 GND.n5482 GND.n1174 9.3005
R15032 GND.n5483 GND.n1173 9.3005
R15033 GND.n1172 GND.n1168 9.3005
R15034 GND.n5489 GND.n1167 9.3005
R15035 GND.n5490 GND.n1166 9.3005
R15036 GND.n5491 GND.n1165 9.3005
R15037 GND.n1164 GND.n1160 9.3005
R15038 GND.n5497 GND.n1159 9.3005
R15039 GND.n5498 GND.n1158 9.3005
R15040 GND.n5499 GND.n1157 9.3005
R15041 GND.n1156 GND.n1152 9.3005
R15042 GND.n5505 GND.n1151 9.3005
R15043 GND.n5506 GND.n1150 9.3005
R15044 GND.n5507 GND.n1149 9.3005
R15045 GND.n1148 GND.n1144 9.3005
R15046 GND.n5513 GND.n1143 9.3005
R15047 GND.n5514 GND.n1142 9.3005
R15048 GND.n5515 GND.n1141 9.3005
R15049 GND.n5419 GND.n5418 9.3005
R15050 GND.n1472 GND.n1470 9.3005
R15051 GND.n3493 GND.n3492 9.3005
R15052 GND.n3494 GND.n3486 9.3005
R15053 GND.n3496 GND.n3495 9.3005
R15054 GND.n3497 GND.n3479 9.3005
R15055 GND.n3499 GND.n3498 9.3005
R15056 GND.n3500 GND.n3478 9.3005
R15057 GND.n3502 GND.n3501 9.3005
R15058 GND.n3503 GND.n3473 9.3005
R15059 GND.n3505 GND.n3504 9.3005
R15060 GND.n3508 GND.n3507 9.3005
R15061 GND.n3471 GND.n3470 9.3005
R15062 GND.n3527 GND.n3526 9.3005
R15063 GND.n3528 GND.n3469 9.3005
R15064 GND.n3530 GND.n3529 9.3005
R15065 GND.n3460 GND.n3459 9.3005
R15066 GND.n3545 GND.n3544 9.3005
R15067 GND.n3546 GND.n3458 9.3005
R15068 GND.n3548 GND.n3547 9.3005
R15069 GND.n3448 GND.n3447 9.3005
R15070 GND.n3562 GND.n3561 9.3005
R15071 GND.n3563 GND.n3446 9.3005
R15072 GND.n3565 GND.n3564 9.3005
R15073 GND.n3436 GND.n3435 9.3005
R15074 GND.n3579 GND.n3578 9.3005
R15075 GND.n3580 GND.n3434 9.3005
R15076 GND.n3582 GND.n3581 9.3005
R15077 GND.n3424 GND.n3423 9.3005
R15078 GND.n3596 GND.n3595 9.3005
R15079 GND.n3597 GND.n3421 9.3005
R15080 GND.n3600 GND.n3599 9.3005
R15081 GND.n3598 GND.n3422 9.3005
R15082 GND.n3411 GND.n3410 9.3005
R15083 GND.n3615 GND.n3614 9.3005
R15084 GND.n3616 GND.n3408 9.3005
R15085 GND.n3646 GND.n3645 9.3005
R15086 GND.n3644 GND.n3409 9.3005
R15087 GND.n3643 GND.n3642 9.3005
R15088 GND.n3641 GND.n3617 9.3005
R15089 GND.n3640 GND.n3639 9.3005
R15090 GND.n3638 GND.n3622 9.3005
R15091 GND.n3637 GND.n3636 9.3005
R15092 GND.n3635 GND.n3623 9.3005
R15093 GND.n3634 GND.n3633 9.3005
R15094 GND.n3632 GND.n3625 9.3005
R15095 GND.n3631 GND.n3630 9.3005
R15096 GND.n3629 GND.n3626 9.3005
R15097 GND.n3308 GND.n3307 9.3005
R15098 GND.n3852 GND.n3851 9.3005
R15099 GND.n3853 GND.n3305 9.3005
R15100 GND.n3889 GND.n3888 9.3005
R15101 GND.n3887 GND.n3306 9.3005
R15102 GND.n3886 GND.n3885 9.3005
R15103 GND.n3884 GND.n3854 9.3005
R15104 GND.n3883 GND.n3882 9.3005
R15105 GND.n3881 GND.n3857 9.3005
R15106 GND.n3880 GND.n3879 9.3005
R15107 GND.n3878 GND.n3858 9.3005
R15108 GND.n3877 GND.n3876 9.3005
R15109 GND.n3875 GND.n3864 9.3005
R15110 GND.n3874 GND.n3873 9.3005
R15111 GND.n3872 GND.n3865 9.3005
R15112 GND.n3871 GND.n3870 9.3005
R15113 GND.n3869 GND.n3868 9.3005
R15114 GND.n3220 GND.n3219 9.3005
R15115 GND.n4012 GND.n4011 9.3005
R15116 GND.n4013 GND.n3217 9.3005
R15117 GND.n4050 GND.n4049 9.3005
R15118 GND.n4048 GND.n3218 9.3005
R15119 GND.n4047 GND.n4046 9.3005
R15120 GND.n4045 GND.n4014 9.3005
R15121 GND.n4044 GND.n4043 9.3005
R15122 GND.n4042 GND.n4017 9.3005
R15123 GND.n4041 GND.n4040 9.3005
R15124 GND.n4039 GND.n4018 9.3005
R15125 GND.n4038 GND.n4037 9.3005
R15126 GND.n4036 GND.n4025 9.3005
R15127 GND.n4035 GND.n4034 9.3005
R15128 GND.n4033 GND.n4026 9.3005
R15129 GND.n4032 GND.n4031 9.3005
R15130 GND.n4030 GND.n4029 9.3005
R15131 GND.n3133 GND.n3132 9.3005
R15132 GND.n4172 GND.n4171 9.3005
R15133 GND.n4173 GND.n3130 9.3005
R15134 GND.n4197 GND.n4196 9.3005
R15135 GND.n4195 GND.n3131 9.3005
R15136 GND.n4194 GND.n4193 9.3005
R15137 GND.n4192 GND.n4174 9.3005
R15138 GND.n4191 GND.n4190 9.3005
R15139 GND.n4189 GND.n4177 9.3005
R15140 GND.n4188 GND.n4187 9.3005
R15141 GND.n4186 GND.n4178 9.3005
R15142 GND.n4185 GND.n4184 9.3005
R15143 GND.n4183 GND.n4182 9.3005
R15144 GND.n3068 GND.n3067 9.3005
R15145 GND.n4334 GND.n4333 9.3005
R15146 GND.n4335 GND.n3065 9.3005
R15147 GND.n4338 GND.n4337 9.3005
R15148 GND.n4336 GND.n3066 9.3005
R15149 GND.n3021 GND.n3020 9.3005
R15150 GND.n4401 GND.n4400 9.3005
R15151 GND.n4402 GND.n3019 9.3005
R15152 GND.n4404 GND.n4403 9.3005
R15153 GND.n3009 GND.n3008 9.3005
R15154 GND.n4418 GND.n4417 9.3005
R15155 GND.n4419 GND.n3007 9.3005
R15156 GND.n4421 GND.n4420 9.3005
R15157 GND.n2997 GND.n2996 9.3005
R15158 GND.n4435 GND.n4434 9.3005
R15159 GND.n4436 GND.n2995 9.3005
R15160 GND.n4438 GND.n4437 9.3005
R15161 GND.n2985 GND.n2984 9.3005
R15162 GND.n4452 GND.n4451 9.3005
R15163 GND.n4453 GND.n2983 9.3005
R15164 GND.n4455 GND.n4454 9.3005
R15165 GND.n2972 GND.n2971 9.3005
R15166 GND.n4469 GND.n4468 9.3005
R15167 GND.n4470 GND.n2970 9.3005
R15168 GND.n4472 GND.n4471 9.3005
R15169 GND.n2961 GND.n2960 9.3005
R15170 GND.n4489 GND.n4488 9.3005
R15171 GND.n4490 GND.n2959 9.3005
R15172 GND.n4492 GND.n4491 9.3005
R15173 GND.n2500 GND.n2499 9.3005
R15174 GND.n4980 GND.n4979 9.3005
R15175 GND.n3506 GND.n3472 9.3005
R15176 GND.n4976 GND.n2501 9.3005
R15177 GND.n4975 GND.n4974 9.3005
R15178 GND.n4973 GND.n2504 9.3005
R15179 GND.n4972 GND.n4971 9.3005
R15180 GND.n4970 GND.n2505 9.3005
R15181 GND.n4969 GND.n4968 9.3005
R15182 GND.n4967 GND.n2509 9.3005
R15183 GND.n4966 GND.n4965 9.3005
R15184 GND.n4964 GND.n2510 9.3005
R15185 GND.n4978 GND.n4977 9.3005
R15186 GND.n4522 GND.n4521 9.3005
R15187 GND.n2913 GND.n2910 9.3005
R15188 GND.n2944 GND.n2943 9.3005
R15189 GND.n2940 GND.n2929 9.3005
R15190 GND.n2939 GND.n2938 9.3005
R15191 GND.n2932 GND.n2517 9.3005
R15192 GND.n4961 GND.n4960 9.3005
R15193 GND.n4524 GND.n4523 9.3005
R15194 GND.n2906 GND.n2902 9.3005
R15195 GND.n4963 GND.n4962 9.3005
R15196 GND.n2516 GND.n2514 9.3005
R15197 GND.n2936 GND.n2935 9.3005
R15198 GND.n2937 GND.n2928 9.3005
R15199 GND.n2946 GND.n2945 9.3005
R15200 GND.n2930 GND.n2914 9.3005
R15201 GND.n4520 GND.n4519 9.3005
R15202 GND.n2905 GND.n2903 9.3005
R15203 GND.n4526 GND.n4525 9.3005
R15204 GND.n4528 GND.n4527 9.3005
R15205 GND.n5155 GND.n1537 9.3005
R15206 GND.n5154 GND.n5153 9.3005
R15207 GND.n5152 GND.n2351 9.3005
R15208 GND.n5151 GND.n5150 9.3005
R15209 GND.n5149 GND.n2355 9.3005
R15210 GND.n5148 GND.n5147 9.3005
R15211 GND.n5146 GND.n2356 9.3005
R15212 GND.n5145 GND.n5144 9.3005
R15213 GND.n5143 GND.n2360 9.3005
R15214 GND.n5142 GND.n5141 9.3005
R15215 GND.n5140 GND.n2361 9.3005
R15216 GND.n5139 GND.n5138 9.3005
R15217 GND.n5137 GND.n2365 9.3005
R15218 GND.n5136 GND.n5135 9.3005
R15219 GND.n5134 GND.n2366 9.3005
R15220 GND.n5133 GND.n5132 9.3005
R15221 GND.n5131 GND.n2370 9.3005
R15222 GND.n5130 GND.n5129 9.3005
R15223 GND.n5128 GND.n2371 9.3005
R15224 GND.n5127 GND.n5126 9.3005
R15225 GND.n5125 GND.n2375 9.3005
R15226 GND.n5124 GND.n5123 9.3005
R15227 GND.n5122 GND.n2376 9.3005
R15228 GND.n5121 GND.n5120 9.3005
R15229 GND.n5119 GND.n2380 9.3005
R15230 GND.n5118 GND.n5117 9.3005
R15231 GND.n5116 GND.n2381 9.3005
R15232 GND.n5115 GND.n5114 9.3005
R15233 GND.n5113 GND.n2385 9.3005
R15234 GND.n5112 GND.n5111 9.3005
R15235 GND.n5110 GND.n2386 9.3005
R15236 GND.n5109 GND.n5108 9.3005
R15237 GND.n5107 GND.n2390 9.3005
R15238 GND.n5106 GND.n5105 9.3005
R15239 GND.n5104 GND.n2391 9.3005
R15240 GND.n5103 GND.n5102 9.3005
R15241 GND.n5101 GND.n2395 9.3005
R15242 GND.n5100 GND.n5099 9.3005
R15243 GND.n5098 GND.n2396 9.3005
R15244 GND.n5097 GND.n5096 9.3005
R15245 GND.n5095 GND.n2400 9.3005
R15246 GND.n5094 GND.n5093 9.3005
R15247 GND.n5092 GND.n2401 9.3005
R15248 GND.n5091 GND.n5090 9.3005
R15249 GND.n5089 GND.n2405 9.3005
R15250 GND.n5088 GND.n5087 9.3005
R15251 GND.n5086 GND.n2406 9.3005
R15252 GND.n5085 GND.n5084 9.3005
R15253 GND.n5083 GND.n2410 9.3005
R15254 GND.n5082 GND.n5081 9.3005
R15255 GND.n5080 GND.n2411 9.3005
R15256 GND.n5079 GND.n5078 9.3005
R15257 GND.n5077 GND.n2415 9.3005
R15258 GND.n5076 GND.n5075 9.3005
R15259 GND.n5074 GND.n2416 9.3005
R15260 GND.n5073 GND.n5072 9.3005
R15261 GND.n5071 GND.n2420 9.3005
R15262 GND.n5070 GND.n5069 9.3005
R15263 GND.n5068 GND.n2421 9.3005
R15264 GND.n5067 GND.n5066 9.3005
R15265 GND.n5065 GND.n2425 9.3005
R15266 GND.n5064 GND.n5063 9.3005
R15267 GND.n5062 GND.n2426 9.3005
R15268 GND.n5061 GND.n5060 9.3005
R15269 GND.n5059 GND.n2430 9.3005
R15270 GND.n5058 GND.n5057 9.3005
R15271 GND.n5056 GND.n2431 9.3005
R15272 GND.n5055 GND.n5054 9.3005
R15273 GND.n5053 GND.n2435 9.3005
R15274 GND.n5052 GND.n5051 9.3005
R15275 GND.n5050 GND.n2436 9.3005
R15276 GND.n5049 GND.n5048 9.3005
R15277 GND.n5047 GND.n2440 9.3005
R15278 GND.n5046 GND.n5045 9.3005
R15279 GND.n5044 GND.n2441 9.3005
R15280 GND.n5043 GND.n5042 9.3005
R15281 GND.n5041 GND.n2445 9.3005
R15282 GND.n5040 GND.n5039 9.3005
R15283 GND.n5038 GND.n2446 9.3005
R15284 GND.n5037 GND.n5036 9.3005
R15285 GND.n5035 GND.n2450 9.3005
R15286 GND.n5034 GND.n5033 9.3005
R15287 GND.n5032 GND.n2451 9.3005
R15288 GND.n5031 GND.n5030 9.3005
R15289 GND.n5029 GND.n2455 9.3005
R15290 GND.n5028 GND.n5027 9.3005
R15291 GND.n5026 GND.n2456 9.3005
R15292 GND.n5025 GND.n5024 9.3005
R15293 GND.n5023 GND.n2460 9.3005
R15294 GND.n5022 GND.n5021 9.3005
R15295 GND.n5020 GND.n2461 9.3005
R15296 GND.n5019 GND.n5018 9.3005
R15297 GND.n5017 GND.n2465 9.3005
R15298 GND.n5016 GND.n5015 9.3005
R15299 GND.n5014 GND.n2466 9.3005
R15300 GND.n5013 GND.n5012 9.3005
R15301 GND.n5011 GND.n2470 9.3005
R15302 GND.n5010 GND.n5009 9.3005
R15303 GND.n5008 GND.n2471 9.3005
R15304 GND.n5007 GND.n5006 9.3005
R15305 GND.n5005 GND.n2475 9.3005
R15306 GND.n5004 GND.n5003 9.3005
R15307 GND.n5002 GND.n2476 9.3005
R15308 GND.n5001 GND.n5000 9.3005
R15309 GND.n4999 GND.n2480 9.3005
R15310 GND.n4998 GND.n4997 9.3005
R15311 GND.n4996 GND.n2481 9.3005
R15312 GND.n4995 GND.n4994 9.3005
R15313 GND.n4993 GND.n2485 9.3005
R15314 GND.n4992 GND.n4991 9.3005
R15315 GND.n4990 GND.n2486 9.3005
R15316 GND.n4989 GND.n4988 9.3005
R15317 GND.n4987 GND.n2490 9.3005
R15318 GND.n4986 GND.n4985 9.3005
R15319 GND.n4984 GND.n2491 9.3005
R15320 GND.n5157 GND.n5156 9.3005
R15321 GND.n2128 GND.n2127 9.3005
R15322 GND.n2129 GND.n1674 9.3005
R15323 GND.n2131 GND.n2130 9.3005
R15324 GND.n1625 GND.n1624 9.3005
R15325 GND.n2223 GND.n2222 9.3005
R15326 GND.n2224 GND.n1622 9.3005
R15327 GND.n2227 GND.n2226 9.3005
R15328 GND.n2225 GND.n1623 9.3005
R15329 GND.n1601 GND.n1600 9.3005
R15330 GND.n2247 GND.n2246 9.3005
R15331 GND.n2248 GND.n1598 9.3005
R15332 GND.n2251 GND.n2250 9.3005
R15333 GND.n2249 GND.n1599 9.3005
R15334 GND.n1578 GND.n1577 9.3005
R15335 GND.n2272 GND.n2271 9.3005
R15336 GND.n2273 GND.n1575 9.3005
R15337 GND.n2290 GND.n2289 9.3005
R15338 GND.n2288 GND.n1576 9.3005
R15339 GND.n2287 GND.n2286 9.3005
R15340 GND.n2285 GND.n2274 9.3005
R15341 GND.n2284 GND.n2283 9.3005
R15342 GND.n2282 GND.n2276 9.3005
R15343 GND.n2281 GND.n2280 9.3005
R15344 GND.n2277 GND.n1539 9.3005
R15345 GND.n2347 GND.n1538 9.3005
R15346 GND.n2349 GND.n2348 9.3005
R15347 GND.n5217 GND.n5216 9.3005
R15348 GND.n5215 GND.n5214 9.3005
R15349 GND.n1481 GND.n1480 9.3005
R15350 GND.n5209 GND.n5208 9.3005
R15351 GND.n5207 GND.n5206 9.3005
R15352 GND.n1489 GND.n1488 9.3005
R15353 GND.n1503 GND.n1499 9.3005
R15354 GND.n5195 GND.n5194 9.3005
R15355 GND.n1477 GND.n1471 9.3005
R15356 GND.n5197 GND.n5196 9.3005
R15357 GND.n1498 GND.n1490 9.3005
R15358 GND.n5205 GND.n5204 9.3005
R15359 GND.n1485 GND.n1484 9.3005
R15360 GND.n5211 GND.n5210 9.3005
R15361 GND.n5213 GND.n5212 9.3005
R15362 GND.n1476 GND.n1475 9.3005
R15363 GND.n5219 GND.n5218 9.3005
R15364 GND.n5221 GND.n5220 9.3005
R15365 GND.n1500 GND.n1497 9.3005
R15366 GND.n5261 GND.n1431 9.3005
R15367 GND.n5263 GND.n5262 9.3005
R15368 GND.n5264 GND.n1425 9.3005
R15369 GND.n5266 GND.n5265 9.3005
R15370 GND.n5267 GND.n1424 9.3005
R15371 GND.n5269 GND.n5268 9.3005
R15372 GND.n5270 GND.n1420 9.3005
R15373 GND.n5272 GND.n5271 9.3005
R15374 GND.n5273 GND.n1419 9.3005
R15375 GND.n5275 GND.n5274 9.3005
R15376 GND.n5276 GND.n1415 9.3005
R15377 GND.n5278 GND.n5277 9.3005
R15378 GND.n5279 GND.n1414 9.3005
R15379 GND.n5281 GND.n5280 9.3005
R15380 GND.n5282 GND.n1408 9.3005
R15381 GND.n5284 GND.n5283 9.3005
R15382 GND.n5285 GND.n1407 9.3005
R15383 GND.n5287 GND.n5286 9.3005
R15384 GND.n5288 GND.n1404 9.3005
R15385 GND.n5290 GND.n5289 9.3005
R15386 GND.n5259 GND.n5258 9.3005
R15387 GND.n5257 GND.n1433 9.3005
R15388 GND.n5256 GND.n5255 9.3005
R15389 GND.n5254 GND.n1437 9.3005
R15390 GND.n5253 GND.n5252 9.3005
R15391 GND.n5251 GND.n1438 9.3005
R15392 GND.n5250 GND.n5249 9.3005
R15393 GND.n5248 GND.n1445 9.3005
R15394 GND.n5247 GND.n5246 9.3005
R15395 GND.n5245 GND.n1446 9.3005
R15396 GND.n5244 GND.n5243 9.3005
R15397 GND.n5242 GND.n1450 9.3005
R15398 GND.n5241 GND.n5240 9.3005
R15399 GND.n5239 GND.n1451 9.3005
R15400 GND.n5238 GND.n5237 9.3005
R15401 GND.n5236 GND.n1457 9.3005
R15402 GND.n5235 GND.n5234 9.3005
R15403 GND.n5233 GND.n1458 9.3005
R15404 GND.n5232 GND.n5231 9.3005
R15405 GND.n5230 GND.n1462 9.3005
R15406 GND.n5229 GND.n5228 9.3005
R15407 GND.n5227 GND.n1463 9.3005
R15408 GND.n5226 GND.n1468 9.3005
R15409 GND.n5225 GND.n5224 9.3005
R15410 GND.n1295 GND.n1293 9.3005
R15411 GND.n5371 GND.n5370 9.3005
R15412 GND.n1296 GND.n1294 9.3005
R15413 GND.n5366 GND.n1301 9.3005
R15414 GND.n5365 GND.n1302 9.3005
R15415 GND.n5364 GND.n1303 9.3005
R15416 GND.n2025 GND.n1304 9.3005
R15417 GND.n5360 GND.n1309 9.3005
R15418 GND.n5359 GND.n1310 9.3005
R15419 GND.n5358 GND.n1311 9.3005
R15420 GND.n1718 GND.n1312 9.3005
R15421 GND.n5354 GND.n1317 9.3005
R15422 GND.n5353 GND.n1318 9.3005
R15423 GND.n5352 GND.n1319 9.3005
R15424 GND.n1697 GND.n1320 9.3005
R15425 GND.n5348 GND.n1325 9.3005
R15426 GND.n5347 GND.n1326 9.3005
R15427 GND.n5346 GND.n1327 9.3005
R15428 GND.n1686 GND.n1328 9.3005
R15429 GND.n5342 GND.n1333 9.3005
R15430 GND.n5341 GND.n1334 9.3005
R15431 GND.n5340 GND.n1335 9.3005
R15432 GND.n1649 GND.n1336 9.3005
R15433 GND.n5336 GND.n1341 9.3005
R15434 GND.n5335 GND.n1342 9.3005
R15435 GND.n5334 GND.n1343 9.3005
R15436 GND.n1672 GND.n1344 9.3005
R15437 GND.n5330 GND.n1349 9.3005
R15438 GND.n5329 GND.n1350 9.3005
R15439 GND.n5328 GND.n1351 9.3005
R15440 GND.n1618 GND.n1352 9.3005
R15441 GND.n5324 GND.n1357 9.3005
R15442 GND.n5323 GND.n1358 9.3005
R15443 GND.n5322 GND.n1359 9.3005
R15444 GND.n1605 GND.n1360 9.3005
R15445 GND.n5318 GND.n1365 9.3005
R15446 GND.n5317 GND.n1366 9.3005
R15447 GND.n5316 GND.n1367 9.3005
R15448 GND.n2255 GND.n1368 9.3005
R15449 GND.n5312 GND.n1373 9.3005
R15450 GND.n5311 GND.n1374 9.3005
R15451 GND.n5310 GND.n1375 9.3005
R15452 GND.n2295 GND.n1376 9.3005
R15453 GND.n5306 GND.n1381 9.3005
R15454 GND.n5305 GND.n1382 9.3005
R15455 GND.n5304 GND.n1383 9.3005
R15456 GND.n2332 GND.n1384 9.3005
R15457 GND.n5300 GND.n1389 9.3005
R15458 GND.n5299 GND.n1390 9.3005
R15459 GND.n5298 GND.n1391 9.3005
R15460 GND.n1398 GND.n1392 9.3005
R15461 GND.n1940 GND.n1938 9.3005
R15462 GND.n1297 GND.n1295 9.3005
R15463 GND.n5370 GND.n5369 9.3005
R15464 GND.n5368 GND.n1296 9.3005
R15465 GND.n5367 GND.n5366 9.3005
R15466 GND.n5365 GND.n1300 9.3005
R15467 GND.n5364 GND.n5363 9.3005
R15468 GND.n5362 GND.n1304 9.3005
R15469 GND.n5361 GND.n5360 9.3005
R15470 GND.n5359 GND.n1308 9.3005
R15471 GND.n5358 GND.n5357 9.3005
R15472 GND.n5356 GND.n1312 9.3005
R15473 GND.n5355 GND.n5354 9.3005
R15474 GND.n5353 GND.n1316 9.3005
R15475 GND.n5352 GND.n5351 9.3005
R15476 GND.n5350 GND.n1320 9.3005
R15477 GND.n5349 GND.n5348 9.3005
R15478 GND.n5347 GND.n1324 9.3005
R15479 GND.n5346 GND.n5345 9.3005
R15480 GND.n5344 GND.n1328 9.3005
R15481 GND.n5343 GND.n5342 9.3005
R15482 GND.n5341 GND.n1332 9.3005
R15483 GND.n5340 GND.n5339 9.3005
R15484 GND.n5338 GND.n1336 9.3005
R15485 GND.n5337 GND.n5336 9.3005
R15486 GND.n5335 GND.n1340 9.3005
R15487 GND.n5334 GND.n5333 9.3005
R15488 GND.n5332 GND.n1344 9.3005
R15489 GND.n5331 GND.n5330 9.3005
R15490 GND.n5329 GND.n1348 9.3005
R15491 GND.n5328 GND.n5327 9.3005
R15492 GND.n5326 GND.n1352 9.3005
R15493 GND.n5325 GND.n5324 9.3005
R15494 GND.n5323 GND.n1356 9.3005
R15495 GND.n5322 GND.n5321 9.3005
R15496 GND.n5320 GND.n1360 9.3005
R15497 GND.n5319 GND.n5318 9.3005
R15498 GND.n5317 GND.n1364 9.3005
R15499 GND.n5316 GND.n5315 9.3005
R15500 GND.n5314 GND.n1368 9.3005
R15501 GND.n5313 GND.n5312 9.3005
R15502 GND.n5311 GND.n1372 9.3005
R15503 GND.n5310 GND.n5309 9.3005
R15504 GND.n5308 GND.n1376 9.3005
R15505 GND.n5307 GND.n5306 9.3005
R15506 GND.n5305 GND.n1380 9.3005
R15507 GND.n5304 GND.n5303 9.3005
R15508 GND.n5302 GND.n1384 9.3005
R15509 GND.n5301 GND.n5300 9.3005
R15510 GND.n5299 GND.n1388 9.3005
R15511 GND.n5298 GND.n5297 9.3005
R15512 GND.n5296 GND.n1392 9.3005
R15513 GND.n1940 GND.n1939 9.3005
R15514 GND.n1958 GND.n1957 9.3005
R15515 GND.n1956 GND.n1763 9.3005
R15516 GND.n1955 GND.n1954 9.3005
R15517 GND.n1765 GND.n1764 9.3005
R15518 GND.n1948 GND.n1947 9.3005
R15519 GND.n1946 GND.n1767 9.3005
R15520 GND.n1945 GND.n1944 9.3005
R15521 GND.n1761 GND.n1758 9.3005
R15522 GND.n1964 GND.n1963 9.3005
R15523 GND.n1967 GND.n1757 9.3005
R15524 GND.n1969 GND.n1968 9.3005
R15525 GND.n1970 GND.n1753 9.3005
R15526 GND.n2015 GND.n2014 9.3005
R15527 GND.n2016 GND.n1751 9.3005
R15528 GND.n2019 GND.n2018 9.3005
R15529 GND.n2017 GND.n1752 9.3005
R15530 GND.n1732 GND.n1731 9.3005
R15531 GND.n2040 GND.n2039 9.3005
R15532 GND.n2041 GND.n1729 9.3005
R15533 GND.n2044 GND.n2043 9.3005
R15534 GND.n2042 GND.n1730 9.3005
R15535 GND.n1704 GND.n1703 9.3005
R15536 GND.n2093 GND.n2092 9.3005
R15537 GND.n2094 GND.n1701 9.3005
R15538 GND.n2097 GND.n2096 9.3005
R15539 GND.n2095 GND.n1702 9.3005
R15540 GND.n1680 GND.n1679 9.3005
R15541 GND.n2115 GND.n2114 9.3005
R15542 GND.n2116 GND.n1678 9.3005
R15543 GND.n2118 GND.n2117 9.3005
R15544 GND.n2119 GND.n1677 9.3005
R15545 GND.n2123 GND.n2122 9.3005
R15546 GND.n2124 GND.n1676 9.3005
R15547 GND.n2126 GND.n2125 9.3005
R15548 GND.n1966 GND.n1965 9.3005
R15549 GND.n1432 GND.n1431 8.72777
R15550 GND.n4919 GND.n4918 8.72777
R15551 GND.n4519 GND.n2914 8.53383
R15552 GND.n5204 GND.n1484 8.53383
R15553 GND.n140 GND.t33 8.2505
R15554 GND.n140 GND.t1 8.2505
R15555 GND.n114 GND.t28 8.2505
R15556 GND.n114 GND.t166 8.2505
R15557 GND.n88 GND.t168 8.2505
R15558 GND.n88 GND.t163 8.2505
R15559 GND.n62 GND.t34 8.2505
R15560 GND.n62 GND.t167 8.2505
R15561 GND.n36 GND.t30 8.2505
R15562 GND.n36 GND.t42 8.2505
R15563 GND.n11 GND.t20 8.2505
R15564 GND.n11 GND.t39 8.2505
R15565 GND.n296 GND.t10 8.2505
R15566 GND.n296 GND.t37 8.2505
R15567 GND.n270 GND.t36 8.2505
R15568 GND.n270 GND.t43 8.2505
R15569 GND.n244 GND.t170 8.2505
R15570 GND.n244 GND.t16 8.2505
R15571 GND.n218 GND.t169 8.2505
R15572 GND.n218 GND.t23 8.2505
R15573 GND.n192 GND.t165 8.2505
R15574 GND.n192 GND.t41 8.2505
R15575 GND.n167 GND.t24 8.2505
R15576 GND.n167 GND.t25 8.2505
R15577 GND.n3334 GND.t73 8.208
R15578 GND.t48 GND.n3100 8.208
R15579 GND.n6429 GND.n6428 8.07081
R15580 GND.n1675 GND.n155 8.07081
R15581 GND.n3849 GND.n3310 7.81716
R15582 GND.n3900 GND.n3899 7.81716
R15583 GND.t4 GND.t157 7.81716
R15584 GND.n4009 GND.n3222 7.81716
R15585 GND.n4060 GND.n4059 7.81716
R15586 GND.t164 GND.t160 7.81716
R15587 GND.n4169 GND.n3135 7.81716
R15588 GND.n4207 GND.n4206 7.81716
R15589 GND.t73 GND.n3333 7.42633
R15590 GND.t161 GND.n3327 7.42633
R15591 GND.n3106 GND.t158 7.42633
R15592 GND.n3105 GND.t48 7.42633
R15593 GND.n3756 GND.t92 7.0355
R15594 GND.n50 GND.n24 6.83455
R15595 GND.n206 GND.n180 6.83455
R15596 GND.t19 GND.n1647 6.25383
R15597 GND.t0 GND.n1627 6.25383
R15598 GND.n3313 GND.n3302 6.25383
R15599 GND.n3893 GND.n3892 6.25383
R15600 GND.n3226 GND.n3214 6.25383
R15601 GND.n4053 GND.n4052 6.25383
R15602 GND.n3139 GND.n3127 6.25383
R15603 GND.n4200 GND.n4199 6.25383
R15604 GND.t9 GND.n2730 6.25383
R15605 GND.t15 GND.n336 6.25383
R15606 GND.n155 GND.n154 6.04028
R15607 GND.n6429 GND.n310 6.04028
R15608 GND.n4388 GND.t152 5.863
R15609 GND.n154 GND.n153 4.94662
R15610 GND.n310 GND.n309 4.94662
R15611 GND.n128 GND.n127 4.88412
R15612 GND.n102 GND.n101 4.88412
R15613 GND.n76 GND.n75 4.88412
R15614 GND.n50 GND.n49 4.88412
R15615 GND.n284 GND.n283 4.88412
R15616 GND.n258 GND.n257 4.88412
R15617 GND.n232 GND.n231 4.88412
R15618 GND.n206 GND.n205 4.88412
R15619 GND.n4804 GND.n331 4.74817
R15620 GND.n329 GND.n323 4.74817
R15621 GND.n6421 GND.n324 4.74817
R15622 GND.n332 GND.n328 4.74817
R15623 GND.n2725 GND.n331 4.74817
R15624 GND.n2741 GND.n329 4.74817
R15625 GND.n6422 GND.n6421 4.74817
R15626 GND.n4781 GND.n328 4.74817
R15627 GND.n2214 GND.n2213 4.74817
R15628 GND.n2197 GND.n1638 4.74817
R15629 GND.n2133 GND.n1637 4.74817
R15630 GND.n1636 GND.n1633 4.74817
R15631 GND.n2214 GND.n1640 4.74817
R15632 GND.n1666 GND.n1638 4.74817
R15633 GND.n2196 GND.n1637 4.74817
R15634 GND.n2134 GND.n1636 4.74817
R15635 GND.n2063 GND.n2062 4.74817
R15636 GND.n2203 GND.n2202 4.74817
R15637 GND.n2144 GND.n2143 4.74817
R15638 GND.n2187 GND.n2186 4.74817
R15639 GND.n2182 GND.n2145 4.74817
R15640 GND.n2802 GND.n2747 4.74817
R15641 GND.n4790 GND.n2804 4.74817
R15642 GND.n4788 GND.n4787 4.74817
R15643 GND.n2870 GND.n2807 4.74817
R15644 GND.n2868 GND.n2867 4.74817
R15645 GND.n2062 GND.n1655 4.74817
R15646 GND.n2204 GND.n2203 4.74817
R15647 GND.n2143 GND.n1656 4.74817
R15648 GND.n2188 GND.n2187 4.74817
R15649 GND.n2185 GND.n2145 4.74817
R15650 GND.n2799 GND.n2747 4.74817
R15651 GND.n2804 GND.n2803 4.74817
R15652 GND.n4789 GND.n4788 4.74817
R15653 GND.n2807 GND.n2805 4.74817
R15654 GND.n2869 GND.n2868 4.74817
R15655 GND.n132 GND.n130 4.69785
R15656 GND.n145 GND.n143 4.69785
R15657 GND.n106 GND.n104 4.69785
R15658 GND.n119 GND.n117 4.69785
R15659 GND.n80 GND.n78 4.69785
R15660 GND.n93 GND.n91 4.69785
R15661 GND.n54 GND.n52 4.69785
R15662 GND.n67 GND.n65 4.69785
R15663 GND.n28 GND.n26 4.69785
R15664 GND.n41 GND.n39 4.69785
R15665 GND.n3 GND.n1 4.69785
R15666 GND.n16 GND.n14 4.69785
R15667 GND.n301 GND.n299 4.69785
R15668 GND.n288 GND.n286 4.69785
R15669 GND.n275 GND.n273 4.69785
R15670 GND.n262 GND.n260 4.69785
R15671 GND.n249 GND.n247 4.69785
R15672 GND.n236 GND.n234 4.69785
R15673 GND.n223 GND.n221 4.69785
R15674 GND.n210 GND.n208 4.69785
R15675 GND.n197 GND.n195 4.69785
R15676 GND.n184 GND.n182 4.69785
R15677 GND.n172 GND.n170 4.69785
R15678 GND.n159 GND.n157 4.69785
R15679 GND.n2012 GND.t63 4.6905
R15680 GND.n2334 GND.t77 4.6905
R15681 GND.n3819 GND.n3322 4.6905
R15682 GND.n3298 GND.n3286 4.6905
R15683 GND.n3980 GND.n3235 4.6905
R15684 GND.n3210 GND.n3197 4.6905
R15685 GND.n4140 GND.n3148 4.6905
R15686 GND.n3123 GND.n3111 4.6905
R15687 GND.n4551 GND.t59 4.6905
R15688 GND.n4720 GND.t52 4.6905
R15689 GND.n4918 GND.n2578 4.6132
R15690 GND.n5260 GND.n1432 4.6132
R15691 GND.n4340 GND.t122 3.90883
R15692 GND.n3957 GND.t157 3.518
R15693 GND.n4098 GND.t160 3.518
R15694 GND.n1441 GND.n1437 3.49141
R15695 GND.n4910 GND.n4909 3.49141
R15696 GND.n585 GND.n502 3.49141
R15697 GND.n1885 GND.n1794 3.49141
R15698 GND.n153 GND.n141 3.31084
R15699 GND.n127 GND.n115 3.31084
R15700 GND.n101 GND.n89 3.31084
R15701 GND.n75 GND.n63 3.31084
R15702 GND.n49 GND.n37 3.31084
R15703 GND.n24 GND.n12 3.31084
R15704 GND.n309 GND.n297 3.31084
R15705 GND.n283 GND.n271 3.31084
R15706 GND.n257 GND.n245 3.31084
R15707 GND.n231 GND.n219 3.31084
R15708 GND.n205 GND.n193 3.31084
R15709 GND.n180 GND.n168 3.31084
R15710 GND.n3762 GND.n3369 3.12717
R15711 GND.n3826 GND.n3327 3.12717
R15712 GND.n3923 GND.n3282 3.12717
R15713 GND.n3987 GND.n3241 3.12717
R15714 GND.n4083 GND.n3193 3.12717
R15715 GND.n4147 GND.n3153 3.12717
R15716 GND.n4233 GND.n3106 3.12717
R15717 GND.n3073 GND.n3062 3.12717
R15718 GND.n5252 GND.n1441 3.10353
R15719 GND.n4909 GND.n4908 3.10353
R15720 GND.n588 GND.n502 3.10353
R15721 GND.n1794 GND.n1789 3.10353
R15722 GND.n154 GND.n128 3.03936
R15723 GND.n310 GND.n284 3.03936
R15724 GND.n3862 GND.t4 2.73633
R15725 GND.n4022 GND.t164 2.73633
R15726 GND.n6420 GND.n331 2.27742
R15727 GND.n6420 GND.n329 2.27742
R15728 GND.n6421 GND.n6420 2.27742
R15729 GND.n6420 GND.n328 2.27742
R15730 GND.n2215 GND.n2214 2.27742
R15731 GND.n2215 GND.n1638 2.27742
R15732 GND.n2215 GND.n1637 2.27742
R15733 GND.n2215 GND.n1636 2.27742
R15734 GND.n2203 GND.n1635 2.27742
R15735 GND.n2143 GND.n1635 2.27742
R15736 GND.n2187 GND.n1635 2.27742
R15737 GND.n2145 GND.n1635 2.27742
R15738 GND.n2747 GND.n327 2.27742
R15739 GND.n2804 GND.n327 2.27742
R15740 GND.n4788 GND.n327 2.27742
R15741 GND.n2807 GND.n327 2.27742
R15742 GND.n2868 GND.n327 2.27742
R15743 GND.n2062 GND.n1635 2.27742
R15744 GND.n76 GND.n50 1.95093
R15745 GND.n102 GND.n76 1.95093
R15746 GND.n128 GND.n102 1.95093
R15747 GND.n232 GND.n206 1.95093
R15748 GND.n258 GND.n232 1.95093
R15749 GND.n284 GND.n258 1.95093
R15750 GND.n139 GND.n129 1.93989
R15751 GND.n152 GND.n142 1.93989
R15752 GND.n113 GND.n103 1.93989
R15753 GND.n126 GND.n116 1.93989
R15754 GND.n87 GND.n77 1.93989
R15755 GND.n100 GND.n90 1.93989
R15756 GND.n61 GND.n51 1.93989
R15757 GND.n74 GND.n64 1.93989
R15758 GND.n35 GND.n25 1.93989
R15759 GND.n48 GND.n38 1.93989
R15760 GND.n10 GND.n0 1.93989
R15761 GND.n23 GND.n13 1.93989
R15762 GND.n308 GND.n298 1.93989
R15763 GND.n295 GND.n285 1.93989
R15764 GND.n282 GND.n272 1.93989
R15765 GND.n269 GND.n259 1.93989
R15766 GND.n256 GND.n246 1.93989
R15767 GND.n243 GND.n233 1.93989
R15768 GND.n230 GND.n220 1.93989
R15769 GND.n217 GND.n207 1.93989
R15770 GND.n204 GND.n194 1.93989
R15771 GND.n191 GND.n181 1.93989
R15772 GND.n179 GND.n169 1.93989
R15773 GND.n166 GND.n156 1.93989
R15774 GND.n3369 GND.t70 1.56383
R15775 GND.n3768 GND.n3356 1.56383
R15776 GND.n3795 GND.n3332 1.56383
R15777 GND.n3929 GND.n3269 1.56383
R15778 GND.n3956 GND.n3246 1.56383
R15779 GND.n4089 GND.n3182 1.56383
R15780 GND.n4116 GND.n3158 1.56383
R15781 GND.n4239 GND.n3095 1.56383
R15782 GND.n4302 GND.n3083 1.56383
R15783 GND GND.n155 1.37917
R15784 GND.n4261 GND.n4254 1.24928
R15785 GND.n3688 GND.n3687 1.24928
R15786 GND.n3706 GND.n3705 1.24928
R15787 GND.n4356 GND.n4355 1.24928
R15788 GND.n137 GND.n136 1.16414
R15789 GND.n150 GND.n149 1.16414
R15790 GND.n111 GND.n110 1.16414
R15791 GND.n124 GND.n123 1.16414
R15792 GND.n85 GND.n84 1.16414
R15793 GND.n98 GND.n97 1.16414
R15794 GND.n59 GND.n58 1.16414
R15795 GND.n72 GND.n71 1.16414
R15796 GND.n33 GND.n32 1.16414
R15797 GND.n46 GND.n45 1.16414
R15798 GND.n8 GND.n7 1.16414
R15799 GND.n21 GND.n20 1.16414
R15800 GND.n306 GND.n305 1.16414
R15801 GND.n293 GND.n292 1.16414
R15802 GND.n280 GND.n279 1.16414
R15803 GND.n267 GND.n266 1.16414
R15804 GND.n254 GND.n253 1.16414
R15805 GND.n241 GND.n240 1.16414
R15806 GND.n228 GND.n227 1.16414
R15807 GND.n215 GND.n214 1.16414
R15808 GND.n202 GND.n201 1.16414
R15809 GND.n189 GND.n188 1.16414
R15810 GND.n177 GND.n176 1.16414
R15811 GND.n164 GND.n163 1.16414
R15812 GND GND.n6429 1.03826
R15813 GND.n2090 GND.t5 0.782166
R15814 GND.n2253 GND.t2 0.782166
R15815 GND.n4589 GND.t12 0.782166
R15816 GND.n4750 GND.t21 0.782166
R15817 GND.n2632 GND.n2551 0.529463
R15818 GND.n1819 GND.n1282 0.529463
R15819 GND.n525 GND.n524 0.529463
R15820 GND.n5291 GND.n5290 0.529463
R15821 GND.n3506 GND.n3505 0.494402
R15822 GND.n4979 GND.n4978 0.494402
R15823 GND.n1141 GND.n1136 0.492878
R15824 GND.n6184 GND.n734 0.492878
R15825 GND.n6305 GND.n663 0.492878
R15826 GND.n4709 GND.n4708 0.492878
R15827 GND.n5418 GND.n5417 0.492878
R15828 GND.n1966 GND.n1964 0.492878
R15829 GND.n6420 GND.n327 0.413375
R15830 GND.n2215 GND.n1635 0.413375
R15831 GND.n133 GND.n131 0.388379
R15832 GND.n146 GND.n144 0.388379
R15833 GND.n107 GND.n105 0.388379
R15834 GND.n120 GND.n118 0.388379
R15835 GND.n81 GND.n79 0.388379
R15836 GND.n94 GND.n92 0.388379
R15837 GND.n55 GND.n53 0.388379
R15838 GND.n68 GND.n66 0.388379
R15839 GND.n29 GND.n27 0.388379
R15840 GND.n42 GND.n40 0.388379
R15841 GND.n4 GND.n2 0.388379
R15842 GND.n17 GND.n15 0.388379
R15843 GND.n302 GND.n300 0.388379
R15844 GND.n289 GND.n287 0.388379
R15845 GND.n276 GND.n274 0.388379
R15846 GND.n263 GND.n261 0.388379
R15847 GND.n250 GND.n248 0.388379
R15848 GND.n237 GND.n235 0.388379
R15849 GND.n224 GND.n222 0.388379
R15850 GND.n211 GND.n209 0.388379
R15851 GND.n198 GND.n196 0.388379
R15852 GND.n185 GND.n183 0.388379
R15853 GND.n173 GND.n171 0.388379
R15854 GND.n160 GND.n158 0.388379
R15855 GND.n4256 GND.n2576 0.312695
R15856 GND.n3697 GND.n3695 0.312695
R15857 GND.n3698 GND.n3697 0.312695
R15858 GND.n4348 GND.n2576 0.312695
R15859 GND.n487 GND.n448 0.302329
R15860 GND.n4870 GND.n4868 0.302329
R15861 GND.n1941 GND.n1937 0.302329
R15862 GND.n5224 GND.n5223 0.302329
R15863 GND.n4529 GND.n2491 0.294707
R15864 GND.n5156 GND.n2350 0.294707
R15865 GND.n4531 GND.n4529 0.290134
R15866 GND.n2350 GND.n2349 0.290134
R15867 GND.n4689 GND.n448 0.265744
R15868 GND.n1945 GND.n1941 0.265744
R15869 GND.n2578 GND.n2575 0.229039
R15870 GND.n2579 GND.n2578 0.229039
R15871 GND.n5261 GND.n5260 0.229039
R15872 GND.n5260 GND.n5259 0.229039
R15873 GND.n138 GND.n130 0.155672
R15874 GND.n151 GND.n143 0.155672
R15875 GND.n112 GND.n104 0.155672
R15876 GND.n125 GND.n117 0.155672
R15877 GND.n86 GND.n78 0.155672
R15878 GND.n99 GND.n91 0.155672
R15879 GND.n60 GND.n52 0.155672
R15880 GND.n73 GND.n65 0.155672
R15881 GND.n34 GND.n26 0.155672
R15882 GND.n47 GND.n39 0.155672
R15883 GND.n9 GND.n1 0.155672
R15884 GND.n22 GND.n14 0.155672
R15885 GND.n307 GND.n299 0.155672
R15886 GND.n294 GND.n286 0.155672
R15887 GND.n281 GND.n273 0.155672
R15888 GND.n268 GND.n260 0.155672
R15889 GND.n255 GND.n247 0.155672
R15890 GND.n242 GND.n234 0.155672
R15891 GND.n229 GND.n221 0.155672
R15892 GND.n216 GND.n208 0.155672
R15893 GND.n203 GND.n195 0.155672
R15894 GND.n190 GND.n182 0.155672
R15895 GND.n178 GND.n170 0.155672
R15896 GND.n165 GND.n157 0.155672
R15897 GND.n5522 GND.n1136 0.152939
R15898 GND.n5523 GND.n5522 0.152939
R15899 GND.n5524 GND.n5523 0.152939
R15900 GND.n5524 GND.n1130 0.152939
R15901 GND.n5532 GND.n1130 0.152939
R15902 GND.n5533 GND.n5532 0.152939
R15903 GND.n5534 GND.n5533 0.152939
R15904 GND.n5534 GND.n1124 0.152939
R15905 GND.n5542 GND.n1124 0.152939
R15906 GND.n5543 GND.n5542 0.152939
R15907 GND.n5544 GND.n5543 0.152939
R15908 GND.n5544 GND.n1118 0.152939
R15909 GND.n5552 GND.n1118 0.152939
R15910 GND.n5553 GND.n5552 0.152939
R15911 GND.n5554 GND.n5553 0.152939
R15912 GND.n5554 GND.n1112 0.152939
R15913 GND.n5562 GND.n1112 0.152939
R15914 GND.n5563 GND.n5562 0.152939
R15915 GND.n5564 GND.n5563 0.152939
R15916 GND.n5564 GND.n1106 0.152939
R15917 GND.n5572 GND.n1106 0.152939
R15918 GND.n5573 GND.n5572 0.152939
R15919 GND.n5574 GND.n5573 0.152939
R15920 GND.n5574 GND.n1100 0.152939
R15921 GND.n5582 GND.n1100 0.152939
R15922 GND.n5583 GND.n5582 0.152939
R15923 GND.n5584 GND.n5583 0.152939
R15924 GND.n5584 GND.n1094 0.152939
R15925 GND.n5592 GND.n1094 0.152939
R15926 GND.n5593 GND.n5592 0.152939
R15927 GND.n5594 GND.n5593 0.152939
R15928 GND.n5594 GND.n1088 0.152939
R15929 GND.n5602 GND.n1088 0.152939
R15930 GND.n5603 GND.n5602 0.152939
R15931 GND.n5604 GND.n5603 0.152939
R15932 GND.n5604 GND.n1082 0.152939
R15933 GND.n5612 GND.n1082 0.152939
R15934 GND.n5613 GND.n5612 0.152939
R15935 GND.n5614 GND.n5613 0.152939
R15936 GND.n5614 GND.n1076 0.152939
R15937 GND.n5622 GND.n1076 0.152939
R15938 GND.n5623 GND.n5622 0.152939
R15939 GND.n5624 GND.n5623 0.152939
R15940 GND.n5624 GND.n1070 0.152939
R15941 GND.n5632 GND.n1070 0.152939
R15942 GND.n5633 GND.n5632 0.152939
R15943 GND.n5634 GND.n5633 0.152939
R15944 GND.n5634 GND.n1064 0.152939
R15945 GND.n5642 GND.n1064 0.152939
R15946 GND.n5643 GND.n5642 0.152939
R15947 GND.n5644 GND.n5643 0.152939
R15948 GND.n5644 GND.n1058 0.152939
R15949 GND.n5652 GND.n1058 0.152939
R15950 GND.n5653 GND.n5652 0.152939
R15951 GND.n5654 GND.n5653 0.152939
R15952 GND.n5654 GND.n1052 0.152939
R15953 GND.n5662 GND.n1052 0.152939
R15954 GND.n5663 GND.n5662 0.152939
R15955 GND.n5664 GND.n5663 0.152939
R15956 GND.n5664 GND.n1046 0.152939
R15957 GND.n5672 GND.n1046 0.152939
R15958 GND.n5673 GND.n5672 0.152939
R15959 GND.n5674 GND.n5673 0.152939
R15960 GND.n5674 GND.n1040 0.152939
R15961 GND.n5682 GND.n1040 0.152939
R15962 GND.n5683 GND.n5682 0.152939
R15963 GND.n5684 GND.n5683 0.152939
R15964 GND.n5684 GND.n1034 0.152939
R15965 GND.n5692 GND.n1034 0.152939
R15966 GND.n5693 GND.n5692 0.152939
R15967 GND.n5694 GND.n5693 0.152939
R15968 GND.n5694 GND.n1028 0.152939
R15969 GND.n5702 GND.n1028 0.152939
R15970 GND.n5703 GND.n5702 0.152939
R15971 GND.n5704 GND.n5703 0.152939
R15972 GND.n5704 GND.n1022 0.152939
R15973 GND.n5712 GND.n1022 0.152939
R15974 GND.n5713 GND.n5712 0.152939
R15975 GND.n5714 GND.n5713 0.152939
R15976 GND.n5714 GND.n1016 0.152939
R15977 GND.n5722 GND.n1016 0.152939
R15978 GND.n5723 GND.n5722 0.152939
R15979 GND.n5724 GND.n5723 0.152939
R15980 GND.n5724 GND.n1010 0.152939
R15981 GND.n5732 GND.n1010 0.152939
R15982 GND.n5733 GND.n5732 0.152939
R15983 GND.n5734 GND.n5733 0.152939
R15984 GND.n5734 GND.n1004 0.152939
R15985 GND.n5742 GND.n1004 0.152939
R15986 GND.n5743 GND.n5742 0.152939
R15987 GND.n5744 GND.n5743 0.152939
R15988 GND.n5744 GND.n998 0.152939
R15989 GND.n5752 GND.n998 0.152939
R15990 GND.n5753 GND.n5752 0.152939
R15991 GND.n5754 GND.n5753 0.152939
R15992 GND.n5754 GND.n992 0.152939
R15993 GND.n5762 GND.n992 0.152939
R15994 GND.n5763 GND.n5762 0.152939
R15995 GND.n5764 GND.n5763 0.152939
R15996 GND.n5764 GND.n986 0.152939
R15997 GND.n5772 GND.n986 0.152939
R15998 GND.n5773 GND.n5772 0.152939
R15999 GND.n5774 GND.n5773 0.152939
R16000 GND.n5774 GND.n980 0.152939
R16001 GND.n5782 GND.n980 0.152939
R16002 GND.n5783 GND.n5782 0.152939
R16003 GND.n5784 GND.n5783 0.152939
R16004 GND.n5784 GND.n974 0.152939
R16005 GND.n5792 GND.n974 0.152939
R16006 GND.n5793 GND.n5792 0.152939
R16007 GND.n5794 GND.n5793 0.152939
R16008 GND.n5794 GND.n968 0.152939
R16009 GND.n5802 GND.n968 0.152939
R16010 GND.n5803 GND.n5802 0.152939
R16011 GND.n5804 GND.n5803 0.152939
R16012 GND.n5804 GND.n962 0.152939
R16013 GND.n5812 GND.n962 0.152939
R16014 GND.n5813 GND.n5812 0.152939
R16015 GND.n5814 GND.n5813 0.152939
R16016 GND.n5814 GND.n956 0.152939
R16017 GND.n5822 GND.n956 0.152939
R16018 GND.n5823 GND.n5822 0.152939
R16019 GND.n5824 GND.n5823 0.152939
R16020 GND.n5824 GND.n950 0.152939
R16021 GND.n5832 GND.n950 0.152939
R16022 GND.n5833 GND.n5832 0.152939
R16023 GND.n5834 GND.n5833 0.152939
R16024 GND.n5834 GND.n944 0.152939
R16025 GND.n5842 GND.n944 0.152939
R16026 GND.n5843 GND.n5842 0.152939
R16027 GND.n5844 GND.n5843 0.152939
R16028 GND.n5844 GND.n938 0.152939
R16029 GND.n5852 GND.n938 0.152939
R16030 GND.n5853 GND.n5852 0.152939
R16031 GND.n5854 GND.n5853 0.152939
R16032 GND.n5854 GND.n932 0.152939
R16033 GND.n5862 GND.n932 0.152939
R16034 GND.n5863 GND.n5862 0.152939
R16035 GND.n5864 GND.n5863 0.152939
R16036 GND.n5864 GND.n926 0.152939
R16037 GND.n5872 GND.n926 0.152939
R16038 GND.n5873 GND.n5872 0.152939
R16039 GND.n5874 GND.n5873 0.152939
R16040 GND.n5874 GND.n920 0.152939
R16041 GND.n5882 GND.n920 0.152939
R16042 GND.n5883 GND.n5882 0.152939
R16043 GND.n5884 GND.n5883 0.152939
R16044 GND.n5884 GND.n914 0.152939
R16045 GND.n5892 GND.n914 0.152939
R16046 GND.n5893 GND.n5892 0.152939
R16047 GND.n5894 GND.n5893 0.152939
R16048 GND.n5894 GND.n908 0.152939
R16049 GND.n5902 GND.n908 0.152939
R16050 GND.n5903 GND.n5902 0.152939
R16051 GND.n5904 GND.n5903 0.152939
R16052 GND.n5904 GND.n902 0.152939
R16053 GND.n5912 GND.n902 0.152939
R16054 GND.n5913 GND.n5912 0.152939
R16055 GND.n5914 GND.n5913 0.152939
R16056 GND.n5914 GND.n896 0.152939
R16057 GND.n5922 GND.n896 0.152939
R16058 GND.n5923 GND.n5922 0.152939
R16059 GND.n5924 GND.n5923 0.152939
R16060 GND.n5924 GND.n890 0.152939
R16061 GND.n5932 GND.n890 0.152939
R16062 GND.n5933 GND.n5932 0.152939
R16063 GND.n5934 GND.n5933 0.152939
R16064 GND.n5934 GND.n884 0.152939
R16065 GND.n5942 GND.n884 0.152939
R16066 GND.n5943 GND.n5942 0.152939
R16067 GND.n5944 GND.n5943 0.152939
R16068 GND.n5944 GND.n878 0.152939
R16069 GND.n5952 GND.n878 0.152939
R16070 GND.n5953 GND.n5952 0.152939
R16071 GND.n5954 GND.n5953 0.152939
R16072 GND.n5954 GND.n872 0.152939
R16073 GND.n5962 GND.n872 0.152939
R16074 GND.n5963 GND.n5962 0.152939
R16075 GND.n5964 GND.n5963 0.152939
R16076 GND.n5964 GND.n866 0.152939
R16077 GND.n5972 GND.n866 0.152939
R16078 GND.n5973 GND.n5972 0.152939
R16079 GND.n5974 GND.n5973 0.152939
R16080 GND.n5974 GND.n860 0.152939
R16081 GND.n5982 GND.n860 0.152939
R16082 GND.n5983 GND.n5982 0.152939
R16083 GND.n5984 GND.n5983 0.152939
R16084 GND.n5984 GND.n854 0.152939
R16085 GND.n5992 GND.n854 0.152939
R16086 GND.n5993 GND.n5992 0.152939
R16087 GND.n5994 GND.n5993 0.152939
R16088 GND.n5994 GND.n848 0.152939
R16089 GND.n6002 GND.n848 0.152939
R16090 GND.n6003 GND.n6002 0.152939
R16091 GND.n6004 GND.n6003 0.152939
R16092 GND.n6004 GND.n842 0.152939
R16093 GND.n6012 GND.n842 0.152939
R16094 GND.n6013 GND.n6012 0.152939
R16095 GND.n6014 GND.n6013 0.152939
R16096 GND.n6014 GND.n836 0.152939
R16097 GND.n6022 GND.n836 0.152939
R16098 GND.n6023 GND.n6022 0.152939
R16099 GND.n6024 GND.n6023 0.152939
R16100 GND.n6024 GND.n830 0.152939
R16101 GND.n6032 GND.n830 0.152939
R16102 GND.n6033 GND.n6032 0.152939
R16103 GND.n6034 GND.n6033 0.152939
R16104 GND.n6034 GND.n824 0.152939
R16105 GND.n6042 GND.n824 0.152939
R16106 GND.n6043 GND.n6042 0.152939
R16107 GND.n6044 GND.n6043 0.152939
R16108 GND.n6044 GND.n818 0.152939
R16109 GND.n6052 GND.n818 0.152939
R16110 GND.n6053 GND.n6052 0.152939
R16111 GND.n6054 GND.n6053 0.152939
R16112 GND.n6054 GND.n812 0.152939
R16113 GND.n6062 GND.n812 0.152939
R16114 GND.n6063 GND.n6062 0.152939
R16115 GND.n6064 GND.n6063 0.152939
R16116 GND.n6064 GND.n806 0.152939
R16117 GND.n6072 GND.n806 0.152939
R16118 GND.n6073 GND.n6072 0.152939
R16119 GND.n6074 GND.n6073 0.152939
R16120 GND.n6074 GND.n800 0.152939
R16121 GND.n6082 GND.n800 0.152939
R16122 GND.n6083 GND.n6082 0.152939
R16123 GND.n6084 GND.n6083 0.152939
R16124 GND.n6084 GND.n794 0.152939
R16125 GND.n6092 GND.n794 0.152939
R16126 GND.n6093 GND.n6092 0.152939
R16127 GND.n6094 GND.n6093 0.152939
R16128 GND.n6094 GND.n788 0.152939
R16129 GND.n6102 GND.n788 0.152939
R16130 GND.n6103 GND.n6102 0.152939
R16131 GND.n6104 GND.n6103 0.152939
R16132 GND.n6104 GND.n782 0.152939
R16133 GND.n6112 GND.n782 0.152939
R16134 GND.n6113 GND.n6112 0.152939
R16135 GND.n6114 GND.n6113 0.152939
R16136 GND.n6114 GND.n776 0.152939
R16137 GND.n6122 GND.n776 0.152939
R16138 GND.n6123 GND.n6122 0.152939
R16139 GND.n6124 GND.n6123 0.152939
R16140 GND.n6124 GND.n770 0.152939
R16141 GND.n6132 GND.n770 0.152939
R16142 GND.n6133 GND.n6132 0.152939
R16143 GND.n6134 GND.n6133 0.152939
R16144 GND.n6134 GND.n764 0.152939
R16145 GND.n6142 GND.n764 0.152939
R16146 GND.n6143 GND.n6142 0.152939
R16147 GND.n6144 GND.n6143 0.152939
R16148 GND.n6144 GND.n758 0.152939
R16149 GND.n6152 GND.n758 0.152939
R16150 GND.n6153 GND.n6152 0.152939
R16151 GND.n6154 GND.n6153 0.152939
R16152 GND.n6154 GND.n752 0.152939
R16153 GND.n6162 GND.n752 0.152939
R16154 GND.n6163 GND.n6162 0.152939
R16155 GND.n6164 GND.n6163 0.152939
R16156 GND.n6164 GND.n746 0.152939
R16157 GND.n6172 GND.n746 0.152939
R16158 GND.n6173 GND.n6172 0.152939
R16159 GND.n6174 GND.n6173 0.152939
R16160 GND.n6174 GND.n740 0.152939
R16161 GND.n6182 GND.n740 0.152939
R16162 GND.n6183 GND.n6182 0.152939
R16163 GND.n6184 GND.n6183 0.152939
R16164 GND.n6192 GND.n734 0.152939
R16165 GND.n6193 GND.n6192 0.152939
R16166 GND.n6194 GND.n6193 0.152939
R16167 GND.n6194 GND.n728 0.152939
R16168 GND.n6202 GND.n728 0.152939
R16169 GND.n6203 GND.n6202 0.152939
R16170 GND.n6204 GND.n6203 0.152939
R16171 GND.n6204 GND.n722 0.152939
R16172 GND.n6212 GND.n722 0.152939
R16173 GND.n6213 GND.n6212 0.152939
R16174 GND.n6214 GND.n6213 0.152939
R16175 GND.n6214 GND.n716 0.152939
R16176 GND.n6222 GND.n716 0.152939
R16177 GND.n6223 GND.n6222 0.152939
R16178 GND.n6224 GND.n6223 0.152939
R16179 GND.n6224 GND.n710 0.152939
R16180 GND.n6232 GND.n710 0.152939
R16181 GND.n6233 GND.n6232 0.152939
R16182 GND.n6234 GND.n6233 0.152939
R16183 GND.n6234 GND.n704 0.152939
R16184 GND.n6242 GND.n704 0.152939
R16185 GND.n6243 GND.n6242 0.152939
R16186 GND.n6244 GND.n6243 0.152939
R16187 GND.n6244 GND.n698 0.152939
R16188 GND.n6252 GND.n698 0.152939
R16189 GND.n6253 GND.n6252 0.152939
R16190 GND.n6254 GND.n6253 0.152939
R16191 GND.n6254 GND.n692 0.152939
R16192 GND.n6262 GND.n692 0.152939
R16193 GND.n6263 GND.n6262 0.152939
R16194 GND.n6264 GND.n6263 0.152939
R16195 GND.n6264 GND.n686 0.152939
R16196 GND.n6272 GND.n686 0.152939
R16197 GND.n6273 GND.n6272 0.152939
R16198 GND.n6274 GND.n6273 0.152939
R16199 GND.n6274 GND.n680 0.152939
R16200 GND.n6282 GND.n680 0.152939
R16201 GND.n6283 GND.n6282 0.152939
R16202 GND.n6284 GND.n6283 0.152939
R16203 GND.n6284 GND.n674 0.152939
R16204 GND.n6292 GND.n674 0.152939
R16205 GND.n6293 GND.n6292 0.152939
R16206 GND.n6294 GND.n6293 0.152939
R16207 GND.n6294 GND.n668 0.152939
R16208 GND.n6302 GND.n668 0.152939
R16209 GND.n6303 GND.n6302 0.152939
R16210 GND.n6304 GND.n6303 0.152939
R16211 GND.n6305 GND.n6304 0.152939
R16212 GND.n2810 GND.n327 0.152939
R16213 GND.n2811 GND.n2810 0.152939
R16214 GND.n2812 GND.n2811 0.152939
R16215 GND.n2813 GND.n2812 0.152939
R16216 GND.n2816 GND.n2813 0.152939
R16217 GND.n2817 GND.n2816 0.152939
R16218 GND.n2818 GND.n2817 0.152939
R16219 GND.n2819 GND.n2818 0.152939
R16220 GND.n2822 GND.n2819 0.152939
R16221 GND.n2823 GND.n2822 0.152939
R16222 GND.n2824 GND.n2823 0.152939
R16223 GND.n2825 GND.n2824 0.152939
R16224 GND.n2828 GND.n2825 0.152939
R16225 GND.n2829 GND.n2828 0.152939
R16226 GND.n2830 GND.n2829 0.152939
R16227 GND.n2831 GND.n2830 0.152939
R16228 GND.n2834 GND.n2831 0.152939
R16229 GND.n2835 GND.n2834 0.152939
R16230 GND.n2837 GND.n2835 0.152939
R16231 GND.n2837 GND.n2836 0.152939
R16232 GND.n2836 GND.n456 0.152939
R16233 GND.n457 GND.n456 0.152939
R16234 GND.n458 GND.n457 0.152939
R16235 GND.n636 GND.n458 0.152939
R16236 GND.n637 GND.n636 0.152939
R16237 GND.n638 GND.n637 0.152939
R16238 GND.n639 GND.n638 0.152939
R16239 GND.n644 GND.n639 0.152939
R16240 GND.n645 GND.n644 0.152939
R16241 GND.n646 GND.n645 0.152939
R16242 GND.n647 GND.n646 0.152939
R16243 GND.n652 GND.n647 0.152939
R16244 GND.n653 GND.n652 0.152939
R16245 GND.n654 GND.n653 0.152939
R16246 GND.n655 GND.n654 0.152939
R16247 GND.n660 GND.n655 0.152939
R16248 GND.n661 GND.n660 0.152939
R16249 GND.n662 GND.n661 0.152939
R16250 GND.n663 GND.n662 0.152939
R16251 GND.n353 GND.n325 0.152939
R16252 GND.n354 GND.n353 0.152939
R16253 GND.n355 GND.n354 0.152939
R16254 GND.n373 GND.n355 0.152939
R16255 GND.n374 GND.n373 0.152939
R16256 GND.n375 GND.n374 0.152939
R16257 GND.n376 GND.n375 0.152939
R16258 GND.n394 GND.n376 0.152939
R16259 GND.n395 GND.n394 0.152939
R16260 GND.n396 GND.n395 0.152939
R16261 GND.n397 GND.n396 0.152939
R16262 GND.n415 GND.n397 0.152939
R16263 GND.n416 GND.n415 0.152939
R16264 GND.n417 GND.n416 0.152939
R16265 GND.n418 GND.n417 0.152939
R16266 GND.n436 GND.n418 0.152939
R16267 GND.n437 GND.n436 0.152939
R16268 GND.n438 GND.n437 0.152939
R16269 GND.n439 GND.n438 0.152939
R16270 GND.n524 GND.n439 0.152939
R16271 GND.n4532 GND.n4531 0.152939
R16272 GND.n4533 GND.n4532 0.152939
R16273 GND.n4533 GND.n2900 0.152939
R16274 GND.n4554 GND.n2900 0.152939
R16275 GND.n4555 GND.n4554 0.152939
R16276 GND.n4556 GND.n4555 0.152939
R16277 GND.n4556 GND.n2896 0.152939
R16278 GND.n4569 GND.n2896 0.152939
R16279 GND.n4570 GND.n4569 0.152939
R16280 GND.n4571 GND.n4570 0.152939
R16281 GND.n4571 GND.n2892 0.152939
R16282 GND.n4584 GND.n2892 0.152939
R16283 GND.n4585 GND.n4584 0.152939
R16284 GND.n4586 GND.n4585 0.152939
R16285 GND.n4586 GND.n2888 0.152939
R16286 GND.n4599 GND.n2888 0.152939
R16287 GND.n4600 GND.n4599 0.152939
R16288 GND.n4601 GND.n4600 0.152939
R16289 GND.n4601 GND.n2884 0.152939
R16290 GND.n4614 GND.n2884 0.152939
R16291 GND.n4615 GND.n4614 0.152939
R16292 GND.n4616 GND.n4615 0.152939
R16293 GND.n4617 GND.n4616 0.152939
R16294 GND.n4618 GND.n4617 0.152939
R16295 GND.n4618 GND.n311 0.152939
R16296 GND.n6427 GND.n312 0.152939
R16297 GND.n4639 GND.n312 0.152939
R16298 GND.n4640 GND.n4639 0.152939
R16299 GND.n4641 GND.n4640 0.152939
R16300 GND.n4642 GND.n4641 0.152939
R16301 GND.n4646 GND.n4642 0.152939
R16302 GND.n4647 GND.n4646 0.152939
R16303 GND.n4648 GND.n4647 0.152939
R16304 GND.n4649 GND.n4648 0.152939
R16305 GND.n4653 GND.n4649 0.152939
R16306 GND.n4654 GND.n4653 0.152939
R16307 GND.n4655 GND.n4654 0.152939
R16308 GND.n4656 GND.n4655 0.152939
R16309 GND.n4660 GND.n4656 0.152939
R16310 GND.n4661 GND.n4660 0.152939
R16311 GND.n4662 GND.n4661 0.152939
R16312 GND.n4663 GND.n4662 0.152939
R16313 GND.n4667 GND.n4663 0.152939
R16314 GND.n4668 GND.n4667 0.152939
R16315 GND.n4669 GND.n4668 0.152939
R16316 GND.n4670 GND.n4669 0.152939
R16317 GND.n4673 GND.n4670 0.152939
R16318 GND.n4674 GND.n4673 0.152939
R16319 GND.n4675 GND.n4674 0.152939
R16320 GND.n4709 GND.n4675 0.152939
R16321 GND.n4690 GND.n4689 0.152939
R16322 GND.n4691 GND.n4690 0.152939
R16323 GND.n4691 GND.n4682 0.152939
R16324 GND.n4699 GND.n4682 0.152939
R16325 GND.n4700 GND.n4699 0.152939
R16326 GND.n4701 GND.n4700 0.152939
R16327 GND.n4701 GND.n4676 0.152939
R16328 GND.n4708 GND.n4676 0.152939
R16329 GND.n526 GND.n525 0.152939
R16330 GND.n526 GND.n521 0.152939
R16331 GND.n534 GND.n521 0.152939
R16332 GND.n535 GND.n534 0.152939
R16333 GND.n536 GND.n535 0.152939
R16334 GND.n536 GND.n515 0.152939
R16335 GND.n542 GND.n515 0.152939
R16336 GND.n543 GND.n542 0.152939
R16337 GND.n544 GND.n543 0.152939
R16338 GND.n544 GND.n513 0.152939
R16339 GND.n552 GND.n513 0.152939
R16340 GND.n553 GND.n552 0.152939
R16341 GND.n554 GND.n553 0.152939
R16342 GND.n554 GND.n511 0.152939
R16343 GND.n562 GND.n511 0.152939
R16344 GND.n563 GND.n562 0.152939
R16345 GND.n564 GND.n563 0.152939
R16346 GND.n564 GND.n507 0.152939
R16347 GND.n572 GND.n507 0.152939
R16348 GND.n573 GND.n572 0.152939
R16349 GND.n574 GND.n573 0.152939
R16350 GND.n574 GND.n505 0.152939
R16351 GND.n582 GND.n505 0.152939
R16352 GND.n583 GND.n582 0.152939
R16353 GND.n584 GND.n583 0.152939
R16354 GND.n584 GND.n503 0.152939
R16355 GND.n503 GND.n499 0.152939
R16356 GND.n593 GND.n499 0.152939
R16357 GND.n594 GND.n593 0.152939
R16358 GND.n595 GND.n594 0.152939
R16359 GND.n595 GND.n497 0.152939
R16360 GND.n603 GND.n497 0.152939
R16361 GND.n604 GND.n603 0.152939
R16362 GND.n605 GND.n604 0.152939
R16363 GND.n605 GND.n495 0.152939
R16364 GND.n495 GND.n492 0.152939
R16365 GND.n616 GND.n492 0.152939
R16366 GND.n617 GND.n616 0.152939
R16367 GND.n618 GND.n617 0.152939
R16368 GND.n618 GND.n490 0.152939
R16369 GND.n626 GND.n490 0.152939
R16370 GND.n627 GND.n626 0.152939
R16371 GND.n628 GND.n627 0.152939
R16372 GND.n628 GND.n488 0.152939
R16373 GND.n488 GND.n487 0.152939
R16374 GND.n2552 GND.n2551 0.152939
R16375 GND.n2553 GND.n2552 0.152939
R16376 GND.n2554 GND.n2553 0.152939
R16377 GND.n2555 GND.n2554 0.152939
R16378 GND.n2556 GND.n2555 0.152939
R16379 GND.n2557 GND.n2556 0.152939
R16380 GND.n2558 GND.n2557 0.152939
R16381 GND.n2561 GND.n2558 0.152939
R16382 GND.n2562 GND.n2561 0.152939
R16383 GND.n2563 GND.n2562 0.152939
R16384 GND.n2564 GND.n2563 0.152939
R16385 GND.n2565 GND.n2564 0.152939
R16386 GND.n2566 GND.n2565 0.152939
R16387 GND.n2567 GND.n2566 0.152939
R16388 GND.n2568 GND.n2567 0.152939
R16389 GND.n2570 GND.n2568 0.152939
R16390 GND.n2573 GND.n2570 0.152939
R16391 GND.n2574 GND.n2573 0.152939
R16392 GND.n2575 GND.n2574 0.152939
R16393 GND.n2580 GND.n2579 0.152939
R16394 GND.n2581 GND.n2580 0.152939
R16395 GND.n2582 GND.n2581 0.152939
R16396 GND.n2585 GND.n2582 0.152939
R16397 GND.n2586 GND.n2585 0.152939
R16398 GND.n2587 GND.n2586 0.152939
R16399 GND.n2588 GND.n2587 0.152939
R16400 GND.n2589 GND.n2588 0.152939
R16401 GND.n2590 GND.n2589 0.152939
R16402 GND.n2591 GND.n2590 0.152939
R16403 GND.n2592 GND.n2591 0.152939
R16404 GND.n2593 GND.n2592 0.152939
R16405 GND.n2594 GND.n2593 0.152939
R16406 GND.n2597 GND.n2594 0.152939
R16407 GND.n2598 GND.n2597 0.152939
R16408 GND.n2599 GND.n2598 0.152939
R16409 GND.n2600 GND.n2599 0.152939
R16410 GND.n2601 GND.n2600 0.152939
R16411 GND.n2602 GND.n2601 0.152939
R16412 GND.n2603 GND.n2602 0.152939
R16413 GND.n4872 GND.n2603 0.152939
R16414 GND.n4872 GND.n4871 0.152939
R16415 GND.n4871 GND.n4870 0.152939
R16416 GND.n2636 GND.n2632 0.152939
R16417 GND.n2637 GND.n2636 0.152939
R16418 GND.n2638 GND.n2637 0.152939
R16419 GND.n2639 GND.n2638 0.152939
R16420 GND.n2640 GND.n2639 0.152939
R16421 GND.n2660 GND.n2640 0.152939
R16422 GND.n2661 GND.n2660 0.152939
R16423 GND.n2662 GND.n2661 0.152939
R16424 GND.n2663 GND.n2662 0.152939
R16425 GND.n2681 GND.n2663 0.152939
R16426 GND.n2682 GND.n2681 0.152939
R16427 GND.n2683 GND.n2682 0.152939
R16428 GND.n2684 GND.n2683 0.152939
R16429 GND.n2702 GND.n2684 0.152939
R16430 GND.n2703 GND.n2702 0.152939
R16431 GND.n2704 GND.n2703 0.152939
R16432 GND.n2705 GND.n2704 0.152939
R16433 GND.n2723 GND.n2705 0.152939
R16434 GND.n2724 GND.n2723 0.152939
R16435 GND.n2724 GND.n326 0.152939
R16436 GND.n2147 GND.n1635 0.152939
R16437 GND.n2148 GND.n2147 0.152939
R16438 GND.n2151 GND.n2148 0.152939
R16439 GND.n2152 GND.n2151 0.152939
R16440 GND.n2153 GND.n2152 0.152939
R16441 GND.n2154 GND.n2153 0.152939
R16442 GND.n2157 GND.n2154 0.152939
R16443 GND.n2158 GND.n2157 0.152939
R16444 GND.n2159 GND.n2158 0.152939
R16445 GND.n2160 GND.n2159 0.152939
R16446 GND.n2162 GND.n2160 0.152939
R16447 GND.n2163 GND.n2162 0.152939
R16448 GND.n2163 GND.n1558 0.152939
R16449 GND.n2309 GND.n1558 0.152939
R16450 GND.n2310 GND.n2309 0.152939
R16451 GND.n2311 GND.n2310 0.152939
R16452 GND.n2312 GND.n2311 0.152939
R16453 GND.n2313 GND.n2312 0.152939
R16454 GND.n2316 GND.n2313 0.152939
R16455 GND.n2317 GND.n2316 0.152939
R16456 GND.n2319 GND.n2317 0.152939
R16457 GND.n2319 GND.n2318 0.152939
R16458 GND.n2318 GND.n1528 0.152939
R16459 GND.n1529 GND.n1528 0.152939
R16460 GND.n1530 GND.n1529 0.152939
R16461 GND.n3514 GND.n1530 0.152939
R16462 GND.n3515 GND.n3514 0.152939
R16463 GND.n3519 GND.n3515 0.152939
R16464 GND.n3520 GND.n3519 0.152939
R16465 GND.n3521 GND.n3520 0.152939
R16466 GND.n3521 GND.n3464 0.152939
R16467 GND.n3537 GND.n3464 0.152939
R16468 GND.n3538 GND.n3537 0.152939
R16469 GND.n3539 GND.n3538 0.152939
R16470 GND.n3539 GND.n3453 0.152939
R16471 GND.n3554 GND.n3453 0.152939
R16472 GND.n3555 GND.n3554 0.152939
R16473 GND.n3556 GND.n3555 0.152939
R16474 GND.n3556 GND.n3441 0.152939
R16475 GND.n3571 GND.n3441 0.152939
R16476 GND.n3572 GND.n3571 0.152939
R16477 GND.n3573 GND.n3572 0.152939
R16478 GND.n3573 GND.n3429 0.152939
R16479 GND.n3588 GND.n3429 0.152939
R16480 GND.n3589 GND.n3588 0.152939
R16481 GND.n3590 GND.n3589 0.152939
R16482 GND.n3590 GND.n3416 0.152939
R16483 GND.n3606 GND.n3416 0.152939
R16484 GND.n3607 GND.n3606 0.152939
R16485 GND.n3608 GND.n3607 0.152939
R16486 GND.n3608 GND.n3383 0.152939
R16487 GND.n3742 GND.n3383 0.152939
R16488 GND.n3743 GND.n3742 0.152939
R16489 GND.n3744 GND.n3743 0.152939
R16490 GND.n3745 GND.n3744 0.152939
R16491 GND.n3746 GND.n3745 0.152939
R16492 GND.n3747 GND.n3746 0.152939
R16493 GND.n3747 GND.n3345 0.152939
R16494 GND.n3788 GND.n3345 0.152939
R16495 GND.n3789 GND.n3788 0.152939
R16496 GND.n3790 GND.n3789 0.152939
R16497 GND.n3791 GND.n3790 0.152939
R16498 GND.n3791 GND.n3316 0.152939
R16499 GND.n3842 GND.n3316 0.152939
R16500 GND.n3843 GND.n3842 0.152939
R16501 GND.n3844 GND.n3843 0.152939
R16502 GND.n3845 GND.n3844 0.152939
R16503 GND.n3845 GND.n3292 0.152939
R16504 GND.n3903 GND.n3292 0.152939
R16505 GND.n3904 GND.n3903 0.152939
R16506 GND.n3905 GND.n3904 0.152939
R16507 GND.n3906 GND.n3905 0.152939
R16508 GND.n3907 GND.n3906 0.152939
R16509 GND.n3908 GND.n3907 0.152939
R16510 GND.n3908 GND.n3257 0.152939
R16511 GND.n3949 GND.n3257 0.152939
R16512 GND.n3950 GND.n3949 0.152939
R16513 GND.n3951 GND.n3950 0.152939
R16514 GND.n3952 GND.n3951 0.152939
R16515 GND.n3952 GND.n3229 0.152939
R16516 GND.n4002 GND.n3229 0.152939
R16517 GND.n4003 GND.n4002 0.152939
R16518 GND.n4004 GND.n4003 0.152939
R16519 GND.n4005 GND.n4004 0.152939
R16520 GND.n4005 GND.n3204 0.152939
R16521 GND.n4063 GND.n3204 0.152939
R16522 GND.n4064 GND.n4063 0.152939
R16523 GND.n4065 GND.n4064 0.152939
R16524 GND.n4066 GND.n4065 0.152939
R16525 GND.n4067 GND.n4066 0.152939
R16526 GND.n4068 GND.n4067 0.152939
R16527 GND.n4068 GND.n3171 0.152939
R16528 GND.n4109 GND.n3171 0.152939
R16529 GND.n4110 GND.n4109 0.152939
R16530 GND.n4111 GND.n4110 0.152939
R16531 GND.n4112 GND.n4111 0.152939
R16532 GND.n4112 GND.n3142 0.152939
R16533 GND.n4162 GND.n3142 0.152939
R16534 GND.n4163 GND.n4162 0.152939
R16535 GND.n4164 GND.n4163 0.152939
R16536 GND.n4165 GND.n4164 0.152939
R16537 GND.n4165 GND.n3117 0.152939
R16538 GND.n4210 GND.n3117 0.152939
R16539 GND.n4211 GND.n4210 0.152939
R16540 GND.n4212 GND.n4211 0.152939
R16541 GND.n4213 GND.n4212 0.152939
R16542 GND.n4214 GND.n4213 0.152939
R16543 GND.n4216 GND.n4214 0.152939
R16544 GND.n4217 GND.n4216 0.152939
R16545 GND.n4217 GND.n3076 0.152939
R16546 GND.n4324 GND.n3076 0.152939
R16547 GND.n4325 GND.n4324 0.152939
R16548 GND.n4326 GND.n4325 0.152939
R16549 GND.n4327 GND.n4326 0.152939
R16550 GND.n4327 GND.n3026 0.152939
R16551 GND.n4393 GND.n3026 0.152939
R16552 GND.n4394 GND.n4393 0.152939
R16553 GND.n4395 GND.n4394 0.152939
R16554 GND.n4395 GND.n3014 0.152939
R16555 GND.n4410 GND.n3014 0.152939
R16556 GND.n4411 GND.n4410 0.152939
R16557 GND.n4412 GND.n4411 0.152939
R16558 GND.n4412 GND.n3002 0.152939
R16559 GND.n4427 GND.n3002 0.152939
R16560 GND.n4428 GND.n4427 0.152939
R16561 GND.n4429 GND.n4428 0.152939
R16562 GND.n4429 GND.n2990 0.152939
R16563 GND.n4444 GND.n2990 0.152939
R16564 GND.n4445 GND.n4444 0.152939
R16565 GND.n4446 GND.n4445 0.152939
R16566 GND.n4446 GND.n2978 0.152939
R16567 GND.n4461 GND.n2978 0.152939
R16568 GND.n4462 GND.n4461 0.152939
R16569 GND.n4463 GND.n4462 0.152939
R16570 GND.n4463 GND.n2966 0.152939
R16571 GND.n4478 GND.n2966 0.152939
R16572 GND.n4479 GND.n4478 0.152939
R16573 GND.n4480 GND.n4479 0.152939
R16574 GND.n4482 GND.n4480 0.152939
R16575 GND.n4482 GND.n4481 0.152939
R16576 GND.n4481 GND.n2954 0.152939
R16577 GND.n4500 GND.n2954 0.152939
R16578 GND.n4501 GND.n4500 0.152939
R16579 GND.n4502 GND.n4501 0.152939
R16580 GND.n4503 GND.n4502 0.152939
R16581 GND.n4504 GND.n4503 0.152939
R16582 GND.n4506 GND.n4504 0.152939
R16583 GND.n4506 GND.n4505 0.152939
R16584 GND.n4505 GND.n2618 0.152939
R16585 GND.n2619 GND.n2618 0.152939
R16586 GND.n2620 GND.n2619 0.152939
R16587 GND.n2765 GND.n2620 0.152939
R16588 GND.n2766 GND.n2765 0.152939
R16589 GND.n2767 GND.n2766 0.152939
R16590 GND.n2767 GND.n2761 0.152939
R16591 GND.n2773 GND.n2761 0.152939
R16592 GND.n2774 GND.n2773 0.152939
R16593 GND.n2775 GND.n2774 0.152939
R16594 GND.n2775 GND.n2757 0.152939
R16595 GND.n2781 GND.n2757 0.152939
R16596 GND.n2782 GND.n2781 0.152939
R16597 GND.n2783 GND.n2782 0.152939
R16598 GND.n2783 GND.n2753 0.152939
R16599 GND.n2789 GND.n2753 0.152939
R16600 GND.n2790 GND.n2789 0.152939
R16601 GND.n2792 GND.n2790 0.152939
R16602 GND.n2792 GND.n2791 0.152939
R16603 GND.n2791 GND.n2750 0.152939
R16604 GND.n2750 GND.n327 0.152939
R16605 GND.n2216 GND.n1611 0.152939
R16606 GND.n2237 GND.n1611 0.152939
R16607 GND.n2238 GND.n2237 0.152939
R16608 GND.n2239 GND.n2238 0.152939
R16609 GND.n2240 GND.n2239 0.152939
R16610 GND.n2240 GND.n1588 0.152939
R16611 GND.n2262 GND.n1588 0.152939
R16612 GND.n2263 GND.n2262 0.152939
R16613 GND.n2264 GND.n2263 0.152939
R16614 GND.n2265 GND.n2264 0.152939
R16615 GND.n2265 GND.n1566 0.152939
R16616 GND.n2300 GND.n1566 0.152939
R16617 GND.n2301 GND.n2300 0.152939
R16618 GND.n2302 GND.n2301 0.152939
R16619 GND.n2302 GND.n1547 0.152939
R16620 GND.n2337 GND.n1547 0.152939
R16621 GND.n2338 GND.n2337 0.152939
R16622 GND.n2339 GND.n2338 0.152939
R16623 GND.n2339 GND.n1403 0.152939
R16624 GND.n5291 GND.n1403 0.152939
R16625 GND.n1824 GND.n1819 0.152939
R16626 GND.n1825 GND.n1824 0.152939
R16627 GND.n1826 GND.n1825 0.152939
R16628 GND.n1826 GND.n1815 0.152939
R16629 GND.n1834 GND.n1815 0.152939
R16630 GND.n1835 GND.n1834 0.152939
R16631 GND.n1836 GND.n1835 0.152939
R16632 GND.n1836 GND.n1811 0.152939
R16633 GND.n1846 GND.n1811 0.152939
R16634 GND.n1847 GND.n1846 0.152939
R16635 GND.n1848 GND.n1847 0.152939
R16636 GND.n1848 GND.n1807 0.152939
R16637 GND.n1856 GND.n1807 0.152939
R16638 GND.n1857 GND.n1856 0.152939
R16639 GND.n1858 GND.n1857 0.152939
R16640 GND.n1858 GND.n1801 0.152939
R16641 GND.n1866 GND.n1801 0.152939
R16642 GND.n1867 GND.n1866 0.152939
R16643 GND.n1868 GND.n1867 0.152939
R16644 GND.n1868 GND.n1797 0.152939
R16645 GND.n1876 GND.n1797 0.152939
R16646 GND.n1877 GND.n1876 0.152939
R16647 GND.n1878 GND.n1877 0.152939
R16648 GND.n1878 GND.n1790 0.152939
R16649 GND.n1886 GND.n1790 0.152939
R16650 GND.n1887 GND.n1886 0.152939
R16651 GND.n1888 GND.n1887 0.152939
R16652 GND.n1888 GND.n1786 0.152939
R16653 GND.n1896 GND.n1786 0.152939
R16654 GND.n1897 GND.n1896 0.152939
R16655 GND.n1898 GND.n1897 0.152939
R16656 GND.n1898 GND.n1782 0.152939
R16657 GND.n1906 GND.n1782 0.152939
R16658 GND.n1907 GND.n1906 0.152939
R16659 GND.n1908 GND.n1907 0.152939
R16660 GND.n1908 GND.n1778 0.152939
R16661 GND.n1918 GND.n1778 0.152939
R16662 GND.n1919 GND.n1918 0.152939
R16663 GND.n1920 GND.n1919 0.152939
R16664 GND.n1920 GND.n1774 0.152939
R16665 GND.n1928 GND.n1774 0.152939
R16666 GND.n1929 GND.n1928 0.152939
R16667 GND.n1930 GND.n1929 0.152939
R16668 GND.n1930 GND.n1768 0.152939
R16669 GND.n1937 GND.n1768 0.152939
R16670 GND.n1283 GND.n1282 0.152939
R16671 GND.n1284 GND.n1283 0.152939
R16672 GND.n2006 GND.n1284 0.152939
R16673 GND.n2007 GND.n2006 0.152939
R16674 GND.n2008 GND.n2007 0.152939
R16675 GND.n2008 GND.n1742 0.152939
R16676 GND.n2030 GND.n1742 0.152939
R16677 GND.n2031 GND.n2030 0.152939
R16678 GND.n2032 GND.n2031 0.152939
R16679 GND.n2033 GND.n2032 0.152939
R16680 GND.n2033 GND.n1712 0.152939
R16681 GND.n2083 GND.n1712 0.152939
R16682 GND.n2084 GND.n2083 0.152939
R16683 GND.n2085 GND.n2084 0.152939
R16684 GND.n2086 GND.n2085 0.152939
R16685 GND.n2086 GND.n1690 0.152939
R16686 GND.n2107 GND.n1690 0.152939
R16687 GND.n2108 GND.n2107 0.152939
R16688 GND.n2109 GND.n2108 0.152939
R16689 GND.n2109 GND.n1634 0.152939
R16690 GND.n5417 GND.n1237 0.152939
R16691 GND.n1239 GND.n1237 0.152939
R16692 GND.n1245 GND.n1239 0.152939
R16693 GND.n1246 GND.n1245 0.152939
R16694 GND.n1247 GND.n1246 0.152939
R16695 GND.n1248 GND.n1247 0.152939
R16696 GND.n1253 GND.n1248 0.152939
R16697 GND.n1254 GND.n1253 0.152939
R16698 GND.n1255 GND.n1254 0.152939
R16699 GND.n1256 GND.n1255 0.152939
R16700 GND.n1261 GND.n1256 0.152939
R16701 GND.n1262 GND.n1261 0.152939
R16702 GND.n1263 GND.n1262 0.152939
R16703 GND.n1264 GND.n1263 0.152939
R16704 GND.n1269 GND.n1264 0.152939
R16705 GND.n1270 GND.n1269 0.152939
R16706 GND.n1271 GND.n1270 0.152939
R16707 GND.n1272 GND.n1271 0.152939
R16708 GND.n1978 GND.n1272 0.152939
R16709 GND.n1979 GND.n1978 0.152939
R16710 GND.n1984 GND.n1979 0.152939
R16711 GND.n1985 GND.n1984 0.152939
R16712 GND.n1986 GND.n1985 0.152939
R16713 GND.n1987 GND.n1986 0.152939
R16714 GND.n1988 GND.n1987 0.152939
R16715 GND.n1990 GND.n1988 0.152939
R16716 GND.n1991 GND.n1990 0.152939
R16717 GND.n1992 GND.n1991 0.152939
R16718 GND.n1992 GND.n1724 0.152939
R16719 GND.n2051 GND.n1724 0.152939
R16720 GND.n2052 GND.n2051 0.152939
R16721 GND.n2053 GND.n2052 0.152939
R16722 GND.n2054 GND.n2053 0.152939
R16723 GND.n2055 GND.n2054 0.152939
R16724 GND.n2058 GND.n2055 0.152939
R16725 GND.n2059 GND.n2058 0.152939
R16726 GND.n2060 GND.n2059 0.152939
R16727 GND.n2061 GND.n2060 0.152939
R16728 GND.n2061 GND.n1635 0.152939
R16729 GND.n1142 GND.n1141 0.152939
R16730 GND.n1143 GND.n1142 0.152939
R16731 GND.n1148 GND.n1143 0.152939
R16732 GND.n1149 GND.n1148 0.152939
R16733 GND.n1150 GND.n1149 0.152939
R16734 GND.n1151 GND.n1150 0.152939
R16735 GND.n1156 GND.n1151 0.152939
R16736 GND.n1157 GND.n1156 0.152939
R16737 GND.n1158 GND.n1157 0.152939
R16738 GND.n1159 GND.n1158 0.152939
R16739 GND.n1164 GND.n1159 0.152939
R16740 GND.n1165 GND.n1164 0.152939
R16741 GND.n1166 GND.n1165 0.152939
R16742 GND.n1167 GND.n1166 0.152939
R16743 GND.n1172 GND.n1167 0.152939
R16744 GND.n1173 GND.n1172 0.152939
R16745 GND.n1174 GND.n1173 0.152939
R16746 GND.n1175 GND.n1174 0.152939
R16747 GND.n1180 GND.n1175 0.152939
R16748 GND.n1181 GND.n1180 0.152939
R16749 GND.n1182 GND.n1181 0.152939
R16750 GND.n1183 GND.n1182 0.152939
R16751 GND.n1188 GND.n1183 0.152939
R16752 GND.n1189 GND.n1188 0.152939
R16753 GND.n1190 GND.n1189 0.152939
R16754 GND.n1191 GND.n1190 0.152939
R16755 GND.n1196 GND.n1191 0.152939
R16756 GND.n1197 GND.n1196 0.152939
R16757 GND.n1198 GND.n1197 0.152939
R16758 GND.n1199 GND.n1198 0.152939
R16759 GND.n1204 GND.n1199 0.152939
R16760 GND.n1205 GND.n1204 0.152939
R16761 GND.n1206 GND.n1205 0.152939
R16762 GND.n1207 GND.n1206 0.152939
R16763 GND.n1212 GND.n1207 0.152939
R16764 GND.n1213 GND.n1212 0.152939
R16765 GND.n1214 GND.n1213 0.152939
R16766 GND.n1215 GND.n1214 0.152939
R16767 GND.n1220 GND.n1215 0.152939
R16768 GND.n1221 GND.n1220 0.152939
R16769 GND.n1222 GND.n1221 0.152939
R16770 GND.n1223 GND.n1222 0.152939
R16771 GND.n1228 GND.n1223 0.152939
R16772 GND.n1229 GND.n1228 0.152939
R16773 GND.n1230 GND.n1229 0.152939
R16774 GND.n1231 GND.n1230 0.152939
R16775 GND.n1236 GND.n1231 0.152939
R16776 GND.n5418 GND.n1236 0.152939
R16777 GND.n3505 GND.n3473 0.152939
R16778 GND.n3501 GND.n3473 0.152939
R16779 GND.n3501 GND.n3500 0.152939
R16780 GND.n3500 GND.n3499 0.152939
R16781 GND.n3499 GND.n3479 0.152939
R16782 GND.n3495 GND.n3479 0.152939
R16783 GND.n3495 GND.n3494 0.152939
R16784 GND.n3494 GND.n3493 0.152939
R16785 GND.n3493 GND.n1470 0.152939
R16786 GND.n3507 GND.n3506 0.152939
R16787 GND.n3507 GND.n3470 0.152939
R16788 GND.n3527 GND.n3470 0.152939
R16789 GND.n3528 GND.n3527 0.152939
R16790 GND.n3529 GND.n3528 0.152939
R16791 GND.n3529 GND.n3459 0.152939
R16792 GND.n3545 GND.n3459 0.152939
R16793 GND.n3546 GND.n3545 0.152939
R16794 GND.n3547 GND.n3546 0.152939
R16795 GND.n3547 GND.n3447 0.152939
R16796 GND.n3562 GND.n3447 0.152939
R16797 GND.n3563 GND.n3562 0.152939
R16798 GND.n3564 GND.n3563 0.152939
R16799 GND.n3564 GND.n3435 0.152939
R16800 GND.n3579 GND.n3435 0.152939
R16801 GND.n3580 GND.n3579 0.152939
R16802 GND.n3581 GND.n3580 0.152939
R16803 GND.n3581 GND.n3423 0.152939
R16804 GND.n3596 GND.n3423 0.152939
R16805 GND.n3597 GND.n3596 0.152939
R16806 GND.n3599 GND.n3597 0.152939
R16807 GND.n3599 GND.n3598 0.152939
R16808 GND.n3598 GND.n3410 0.152939
R16809 GND.n3615 GND.n3410 0.152939
R16810 GND.n3616 GND.n3615 0.152939
R16811 GND.n3645 GND.n3616 0.152939
R16812 GND.n3645 GND.n3644 0.152939
R16813 GND.n3644 GND.n3643 0.152939
R16814 GND.n3643 GND.n3617 0.152939
R16815 GND.n3639 GND.n3617 0.152939
R16816 GND.n3639 GND.n3638 0.152939
R16817 GND.n3638 GND.n3637 0.152939
R16818 GND.n3637 GND.n3623 0.152939
R16819 GND.n3633 GND.n3623 0.152939
R16820 GND.n3633 GND.n3632 0.152939
R16821 GND.n3632 GND.n3631 0.152939
R16822 GND.n3631 GND.n3626 0.152939
R16823 GND.n3626 GND.n3307 0.152939
R16824 GND.n3852 GND.n3307 0.152939
R16825 GND.n3853 GND.n3852 0.152939
R16826 GND.n3888 GND.n3853 0.152939
R16827 GND.n3888 GND.n3887 0.152939
R16828 GND.n3887 GND.n3886 0.152939
R16829 GND.n3886 GND.n3854 0.152939
R16830 GND.n3882 GND.n3854 0.152939
R16831 GND.n3882 GND.n3881 0.152939
R16832 GND.n3881 GND.n3880 0.152939
R16833 GND.n3880 GND.n3858 0.152939
R16834 GND.n3876 GND.n3858 0.152939
R16835 GND.n3876 GND.n3875 0.152939
R16836 GND.n3875 GND.n3874 0.152939
R16837 GND.n3874 GND.n3865 0.152939
R16838 GND.n3870 GND.n3865 0.152939
R16839 GND.n3870 GND.n3869 0.152939
R16840 GND.n3869 GND.n3219 0.152939
R16841 GND.n4012 GND.n3219 0.152939
R16842 GND.n4013 GND.n4012 0.152939
R16843 GND.n4049 GND.n4013 0.152939
R16844 GND.n4049 GND.n4048 0.152939
R16845 GND.n4048 GND.n4047 0.152939
R16846 GND.n4047 GND.n4014 0.152939
R16847 GND.n4043 GND.n4014 0.152939
R16848 GND.n4043 GND.n4042 0.152939
R16849 GND.n4042 GND.n4041 0.152939
R16850 GND.n4041 GND.n4018 0.152939
R16851 GND.n4037 GND.n4018 0.152939
R16852 GND.n4037 GND.n4036 0.152939
R16853 GND.n4036 GND.n4035 0.152939
R16854 GND.n4035 GND.n4026 0.152939
R16855 GND.n4031 GND.n4026 0.152939
R16856 GND.n4031 GND.n4030 0.152939
R16857 GND.n4030 GND.n3132 0.152939
R16858 GND.n4172 GND.n3132 0.152939
R16859 GND.n4173 GND.n4172 0.152939
R16860 GND.n4196 GND.n4173 0.152939
R16861 GND.n4196 GND.n4195 0.152939
R16862 GND.n4195 GND.n4194 0.152939
R16863 GND.n4194 GND.n4174 0.152939
R16864 GND.n4190 GND.n4174 0.152939
R16865 GND.n4190 GND.n4189 0.152939
R16866 GND.n4189 GND.n4188 0.152939
R16867 GND.n4188 GND.n4178 0.152939
R16868 GND.n4184 GND.n4178 0.152939
R16869 GND.n4184 GND.n4183 0.152939
R16870 GND.n4183 GND.n3067 0.152939
R16871 GND.n4334 GND.n3067 0.152939
R16872 GND.n4335 GND.n4334 0.152939
R16873 GND.n4337 GND.n4335 0.152939
R16874 GND.n4337 GND.n4336 0.152939
R16875 GND.n4336 GND.n3020 0.152939
R16876 GND.n4401 GND.n3020 0.152939
R16877 GND.n4402 GND.n4401 0.152939
R16878 GND.n4403 GND.n4402 0.152939
R16879 GND.n4403 GND.n3008 0.152939
R16880 GND.n4418 GND.n3008 0.152939
R16881 GND.n4419 GND.n4418 0.152939
R16882 GND.n4420 GND.n4419 0.152939
R16883 GND.n4420 GND.n2996 0.152939
R16884 GND.n4435 GND.n2996 0.152939
R16885 GND.n4436 GND.n4435 0.152939
R16886 GND.n4437 GND.n4436 0.152939
R16887 GND.n4437 GND.n2984 0.152939
R16888 GND.n4452 GND.n2984 0.152939
R16889 GND.n4453 GND.n4452 0.152939
R16890 GND.n4454 GND.n4453 0.152939
R16891 GND.n4454 GND.n2971 0.152939
R16892 GND.n4469 GND.n2971 0.152939
R16893 GND.n4470 GND.n4469 0.152939
R16894 GND.n4471 GND.n4470 0.152939
R16895 GND.n4471 GND.n2960 0.152939
R16896 GND.n4489 GND.n2960 0.152939
R16897 GND.n4490 GND.n4489 0.152939
R16898 GND.n4491 GND.n4490 0.152939
R16899 GND.n4491 GND.n2500 0.152939
R16900 GND.n4979 GND.n2500 0.152939
R16901 GND.n4978 GND.n2501 0.152939
R16902 GND.n4974 GND.n2501 0.152939
R16903 GND.n4974 GND.n4973 0.152939
R16904 GND.n4973 GND.n4972 0.152939
R16905 GND.n4972 GND.n2505 0.152939
R16906 GND.n4968 GND.n2505 0.152939
R16907 GND.n4968 GND.n4967 0.152939
R16908 GND.n4967 GND.n4966 0.152939
R16909 GND.n4966 GND.n2510 0.152939
R16910 GND.n5156 GND.n5155 0.152939
R16911 GND.n5155 GND.n5154 0.152939
R16912 GND.n5154 GND.n2351 0.152939
R16913 GND.n5150 GND.n2351 0.152939
R16914 GND.n5150 GND.n5149 0.152939
R16915 GND.n5149 GND.n5148 0.152939
R16916 GND.n5148 GND.n2356 0.152939
R16917 GND.n5144 GND.n2356 0.152939
R16918 GND.n5144 GND.n5143 0.152939
R16919 GND.n5143 GND.n5142 0.152939
R16920 GND.n5142 GND.n2361 0.152939
R16921 GND.n5138 GND.n2361 0.152939
R16922 GND.n5138 GND.n5137 0.152939
R16923 GND.n5137 GND.n5136 0.152939
R16924 GND.n5136 GND.n2366 0.152939
R16925 GND.n5132 GND.n2366 0.152939
R16926 GND.n5132 GND.n5131 0.152939
R16927 GND.n5131 GND.n5130 0.152939
R16928 GND.n5130 GND.n2371 0.152939
R16929 GND.n5126 GND.n2371 0.152939
R16930 GND.n5126 GND.n5125 0.152939
R16931 GND.n5125 GND.n5124 0.152939
R16932 GND.n5124 GND.n2376 0.152939
R16933 GND.n5120 GND.n2376 0.152939
R16934 GND.n5120 GND.n5119 0.152939
R16935 GND.n5119 GND.n5118 0.152939
R16936 GND.n5118 GND.n2381 0.152939
R16937 GND.n5114 GND.n2381 0.152939
R16938 GND.n5114 GND.n5113 0.152939
R16939 GND.n5113 GND.n5112 0.152939
R16940 GND.n5112 GND.n2386 0.152939
R16941 GND.n5108 GND.n2386 0.152939
R16942 GND.n5108 GND.n5107 0.152939
R16943 GND.n5107 GND.n5106 0.152939
R16944 GND.n5106 GND.n2391 0.152939
R16945 GND.n5102 GND.n2391 0.152939
R16946 GND.n5102 GND.n5101 0.152939
R16947 GND.n5101 GND.n5100 0.152939
R16948 GND.n5100 GND.n2396 0.152939
R16949 GND.n5096 GND.n2396 0.152939
R16950 GND.n5096 GND.n5095 0.152939
R16951 GND.n5095 GND.n5094 0.152939
R16952 GND.n5094 GND.n2401 0.152939
R16953 GND.n5090 GND.n2401 0.152939
R16954 GND.n5090 GND.n5089 0.152939
R16955 GND.n5089 GND.n5088 0.152939
R16956 GND.n5088 GND.n2406 0.152939
R16957 GND.n5084 GND.n2406 0.152939
R16958 GND.n5084 GND.n5083 0.152939
R16959 GND.n5083 GND.n5082 0.152939
R16960 GND.n5082 GND.n2411 0.152939
R16961 GND.n5078 GND.n2411 0.152939
R16962 GND.n5078 GND.n5077 0.152939
R16963 GND.n5077 GND.n5076 0.152939
R16964 GND.n5076 GND.n2416 0.152939
R16965 GND.n5072 GND.n2416 0.152939
R16966 GND.n5072 GND.n5071 0.152939
R16967 GND.n5071 GND.n5070 0.152939
R16968 GND.n5070 GND.n2421 0.152939
R16969 GND.n5066 GND.n2421 0.152939
R16970 GND.n5066 GND.n5065 0.152939
R16971 GND.n5065 GND.n5064 0.152939
R16972 GND.n5064 GND.n2426 0.152939
R16973 GND.n5060 GND.n2426 0.152939
R16974 GND.n5060 GND.n5059 0.152939
R16975 GND.n5059 GND.n5058 0.152939
R16976 GND.n5058 GND.n2431 0.152939
R16977 GND.n5054 GND.n2431 0.152939
R16978 GND.n5054 GND.n5053 0.152939
R16979 GND.n5053 GND.n5052 0.152939
R16980 GND.n5052 GND.n2436 0.152939
R16981 GND.n5048 GND.n2436 0.152939
R16982 GND.n5048 GND.n5047 0.152939
R16983 GND.n5047 GND.n5046 0.152939
R16984 GND.n5046 GND.n2441 0.152939
R16985 GND.n5042 GND.n2441 0.152939
R16986 GND.n5042 GND.n5041 0.152939
R16987 GND.n5041 GND.n5040 0.152939
R16988 GND.n5040 GND.n2446 0.152939
R16989 GND.n5036 GND.n2446 0.152939
R16990 GND.n5036 GND.n5035 0.152939
R16991 GND.n5035 GND.n5034 0.152939
R16992 GND.n5034 GND.n2451 0.152939
R16993 GND.n5030 GND.n2451 0.152939
R16994 GND.n5030 GND.n5029 0.152939
R16995 GND.n5029 GND.n5028 0.152939
R16996 GND.n5028 GND.n2456 0.152939
R16997 GND.n5024 GND.n2456 0.152939
R16998 GND.n5024 GND.n5023 0.152939
R16999 GND.n5023 GND.n5022 0.152939
R17000 GND.n5022 GND.n2461 0.152939
R17001 GND.n5018 GND.n2461 0.152939
R17002 GND.n5018 GND.n5017 0.152939
R17003 GND.n5017 GND.n5016 0.152939
R17004 GND.n5016 GND.n2466 0.152939
R17005 GND.n5012 GND.n2466 0.152939
R17006 GND.n5012 GND.n5011 0.152939
R17007 GND.n5011 GND.n5010 0.152939
R17008 GND.n5010 GND.n2471 0.152939
R17009 GND.n5006 GND.n2471 0.152939
R17010 GND.n5006 GND.n5005 0.152939
R17011 GND.n5005 GND.n5004 0.152939
R17012 GND.n5004 GND.n2476 0.152939
R17013 GND.n5000 GND.n2476 0.152939
R17014 GND.n5000 GND.n4999 0.152939
R17015 GND.n4999 GND.n4998 0.152939
R17016 GND.n4998 GND.n2481 0.152939
R17017 GND.n4994 GND.n2481 0.152939
R17018 GND.n4994 GND.n4993 0.152939
R17019 GND.n4993 GND.n4992 0.152939
R17020 GND.n4992 GND.n2486 0.152939
R17021 GND.n4988 GND.n2486 0.152939
R17022 GND.n4988 GND.n4987 0.152939
R17023 GND.n4987 GND.n4986 0.152939
R17024 GND.n4986 GND.n2491 0.152939
R17025 GND.n2129 GND.n2128 0.152939
R17026 GND.n2130 GND.n2129 0.152939
R17027 GND.n2130 GND.n1624 0.152939
R17028 GND.n2223 GND.n1624 0.152939
R17029 GND.n2224 GND.n2223 0.152939
R17030 GND.n2226 GND.n2224 0.152939
R17031 GND.n2226 GND.n2225 0.152939
R17032 GND.n2225 GND.n1600 0.152939
R17033 GND.n2247 GND.n1600 0.152939
R17034 GND.n2248 GND.n2247 0.152939
R17035 GND.n2250 GND.n2248 0.152939
R17036 GND.n2250 GND.n2249 0.152939
R17037 GND.n2249 GND.n1577 0.152939
R17038 GND.n2272 GND.n1577 0.152939
R17039 GND.n2273 GND.n2272 0.152939
R17040 GND.n2289 GND.n2273 0.152939
R17041 GND.n2289 GND.n2288 0.152939
R17042 GND.n2288 GND.n2287 0.152939
R17043 GND.n2287 GND.n2274 0.152939
R17044 GND.n2283 GND.n2274 0.152939
R17045 GND.n2283 GND.n2282 0.152939
R17046 GND.n2282 GND.n2281 0.152939
R17047 GND.n2281 GND.n2277 0.152939
R17048 GND.n2277 GND.n1538 0.152939
R17049 GND.n2349 GND.n1538 0.152939
R17050 GND.n5290 GND.n1404 0.152939
R17051 GND.n5286 GND.n1404 0.152939
R17052 GND.n5286 GND.n5285 0.152939
R17053 GND.n5285 GND.n5284 0.152939
R17054 GND.n5284 GND.n1408 0.152939
R17055 GND.n5280 GND.n1408 0.152939
R17056 GND.n5280 GND.n5279 0.152939
R17057 GND.n5279 GND.n5278 0.152939
R17058 GND.n5278 GND.n1415 0.152939
R17059 GND.n5274 GND.n1415 0.152939
R17060 GND.n5274 GND.n5273 0.152939
R17061 GND.n5273 GND.n5272 0.152939
R17062 GND.n5272 GND.n1420 0.152939
R17063 GND.n5268 GND.n1420 0.152939
R17064 GND.n5268 GND.n5267 0.152939
R17065 GND.n5267 GND.n5266 0.152939
R17066 GND.n5266 GND.n1425 0.152939
R17067 GND.n5262 GND.n1425 0.152939
R17068 GND.n5262 GND.n5261 0.152939
R17069 GND.n5259 GND.n1433 0.152939
R17070 GND.n5255 GND.n1433 0.152939
R17071 GND.n5255 GND.n5254 0.152939
R17072 GND.n5254 GND.n5253 0.152939
R17073 GND.n5253 GND.n1438 0.152939
R17074 GND.n5249 GND.n1438 0.152939
R17075 GND.n5249 GND.n5248 0.152939
R17076 GND.n5248 GND.n5247 0.152939
R17077 GND.n5247 GND.n1446 0.152939
R17078 GND.n5243 GND.n1446 0.152939
R17079 GND.n5243 GND.n5242 0.152939
R17080 GND.n5242 GND.n5241 0.152939
R17081 GND.n5241 GND.n1451 0.152939
R17082 GND.n5237 GND.n1451 0.152939
R17083 GND.n5237 GND.n5236 0.152939
R17084 GND.n5236 GND.n5235 0.152939
R17085 GND.n5235 GND.n1458 0.152939
R17086 GND.n5231 GND.n1458 0.152939
R17087 GND.n5231 GND.n5230 0.152939
R17088 GND.n5230 GND.n5229 0.152939
R17089 GND.n5229 GND.n1463 0.152939
R17090 GND.n1468 GND.n1463 0.152939
R17091 GND.n5224 GND.n1468 0.152939
R17092 GND.n1946 GND.n1945 0.152939
R17093 GND.n1947 GND.n1946 0.152939
R17094 GND.n1947 GND.n1764 0.152939
R17095 GND.n1955 GND.n1764 0.152939
R17096 GND.n1956 GND.n1955 0.152939
R17097 GND.n1957 GND.n1956 0.152939
R17098 GND.n1957 GND.n1758 0.152939
R17099 GND.n1964 GND.n1758 0.152939
R17100 GND.n1967 GND.n1966 0.152939
R17101 GND.n1968 GND.n1967 0.152939
R17102 GND.n1968 GND.n1753 0.152939
R17103 GND.n2015 GND.n1753 0.152939
R17104 GND.n2016 GND.n2015 0.152939
R17105 GND.n2018 GND.n2016 0.152939
R17106 GND.n2018 GND.n2017 0.152939
R17107 GND.n2017 GND.n1731 0.152939
R17108 GND.n2040 GND.n1731 0.152939
R17109 GND.n2041 GND.n2040 0.152939
R17110 GND.n2043 GND.n2041 0.152939
R17111 GND.n2043 GND.n2042 0.152939
R17112 GND.n2042 GND.n1703 0.152939
R17113 GND.n2093 GND.n1703 0.152939
R17114 GND.n2094 GND.n2093 0.152939
R17115 GND.n2096 GND.n2094 0.152939
R17116 GND.n2096 GND.n2095 0.152939
R17117 GND.n2095 GND.n1679 0.152939
R17118 GND.n2115 GND.n1679 0.152939
R17119 GND.n2116 GND.n2115 0.152939
R17120 GND.n2117 GND.n2116 0.152939
R17121 GND.n2117 GND.n1677 0.152939
R17122 GND.n2123 GND.n1677 0.152939
R17123 GND.n2124 GND.n2123 0.152939
R17124 GND.n2125 GND.n2124 0.152939
R17125 GND.n5222 GND.n1470 0.0995854
R17126 GND.n2515 GND.n2510 0.0995854
R17127 GND.n6420 GND.n325 0.0767195
R17128 GND.n6420 GND.n326 0.0767195
R17129 GND.n2216 GND.n2215 0.0767195
R17130 GND.n2215 GND.n1634 0.0767195
R17131 GND.n6428 GND.n311 0.0695946
R17132 GND.n6428 GND.n6427 0.0695946
R17133 GND.n2128 GND.n1675 0.0695946
R17134 GND.n2125 GND.n1675 0.0695946
R17135 GND.n4868 GND.n2515 0.063
R17136 GND.n5223 GND.n5222 0.063
R17137 GND.n4868 GND.n4867 0.0511114
R17138 GND.n6353 GND.n448 0.0511114
R17139 GND.n1941 GND.n1940 0.0511114
R17140 GND.n5223 GND.n1392 0.0511114
R17141 GND.n4529 GND.n4528 0.0448767
R17142 GND.n2350 GND.n1500 0.0448767
R17143 GND.n4867 GND.n2609 0.0344674
R17144 GND.n4541 GND.n2609 0.0344674
R17145 GND.n4547 GND.n4541 0.0344674
R17146 GND.n4548 GND.n4547 0.0344674
R17147 GND.n4548 GND.n2650 0.0344674
R17148 GND.n2651 GND.n2650 0.0344674
R17149 GND.n2652 GND.n2651 0.0344674
R17150 GND.n4563 GND.n2652 0.0344674
R17151 GND.n4563 GND.n2671 0.0344674
R17152 GND.n2672 GND.n2671 0.0344674
R17153 GND.n2673 GND.n2672 0.0344674
R17154 GND.n4578 GND.n2673 0.0344674
R17155 GND.n4578 GND.n2692 0.0344674
R17156 GND.n2693 GND.n2692 0.0344674
R17157 GND.n2694 GND.n2693 0.0344674
R17158 GND.n4593 GND.n2694 0.0344674
R17159 GND.n4593 GND.n2713 0.0344674
R17160 GND.n2714 GND.n2713 0.0344674
R17161 GND.n2715 GND.n2714 0.0344674
R17162 GND.n4608 GND.n2715 0.0344674
R17163 GND.n4608 GND.n2732 0.0344674
R17164 GND.n2733 GND.n2732 0.0344674
R17165 GND.n2734 GND.n2733 0.0344674
R17166 GND.n4628 GND.n2734 0.0344674
R17167 GND.n4629 GND.n4628 0.0344674
R17168 GND.n4633 GND.n4629 0.0344674
R17169 GND.n4633 GND.n2878 0.0344674
R17170 GND.n4778 GND.n2878 0.0344674
R17171 GND.n4778 GND.n2879 0.0344674
R17172 GND.n2879 GND.n343 0.0344674
R17173 GND.n344 GND.n343 0.0344674
R17174 GND.n345 GND.n344 0.0344674
R17175 GND.n4644 GND.n345 0.0344674
R17176 GND.n4644 GND.n363 0.0344674
R17177 GND.n364 GND.n363 0.0344674
R17178 GND.n365 GND.n364 0.0344674
R17179 GND.n4651 GND.n365 0.0344674
R17180 GND.n4651 GND.n384 0.0344674
R17181 GND.n385 GND.n384 0.0344674
R17182 GND.n386 GND.n385 0.0344674
R17183 GND.n4658 GND.n386 0.0344674
R17184 GND.n4658 GND.n405 0.0344674
R17185 GND.n406 GND.n405 0.0344674
R17186 GND.n407 GND.n406 0.0344674
R17187 GND.n4665 GND.n407 0.0344674
R17188 GND.n4665 GND.n426 0.0344674
R17189 GND.n427 GND.n426 0.0344674
R17190 GND.n428 GND.n427 0.0344674
R17191 GND.n4672 GND.n428 0.0344674
R17192 GND.n4672 GND.n447 0.0344674
R17193 GND.n6353 GND.n447 0.0344674
R17194 GND.n1940 GND.n1295 0.0344674
R17195 GND.n5370 GND.n1295 0.0344674
R17196 GND.n5370 GND.n1296 0.0344674
R17197 GND.n5366 GND.n1296 0.0344674
R17198 GND.n5366 GND.n5365 0.0344674
R17199 GND.n5365 GND.n5364 0.0344674
R17200 GND.n5364 GND.n1304 0.0344674
R17201 GND.n5360 GND.n1304 0.0344674
R17202 GND.n5360 GND.n5359 0.0344674
R17203 GND.n5359 GND.n5358 0.0344674
R17204 GND.n5358 GND.n1312 0.0344674
R17205 GND.n5354 GND.n1312 0.0344674
R17206 GND.n5354 GND.n5353 0.0344674
R17207 GND.n5353 GND.n5352 0.0344674
R17208 GND.n5352 GND.n1320 0.0344674
R17209 GND.n5348 GND.n1320 0.0344674
R17210 GND.n5348 GND.n5347 0.0344674
R17211 GND.n5347 GND.n5346 0.0344674
R17212 GND.n5346 GND.n1328 0.0344674
R17213 GND.n5342 GND.n1328 0.0344674
R17214 GND.n5342 GND.n5341 0.0344674
R17215 GND.n5341 GND.n5340 0.0344674
R17216 GND.n5340 GND.n1336 0.0344674
R17217 GND.n5336 GND.n1336 0.0344674
R17218 GND.n5336 GND.n5335 0.0344674
R17219 GND.n5335 GND.n5334 0.0344674
R17220 GND.n5334 GND.n1344 0.0344674
R17221 GND.n5330 GND.n1344 0.0344674
R17222 GND.n5330 GND.n5329 0.0344674
R17223 GND.n5329 GND.n5328 0.0344674
R17224 GND.n5328 GND.n1352 0.0344674
R17225 GND.n5324 GND.n1352 0.0344674
R17226 GND.n5324 GND.n5323 0.0344674
R17227 GND.n5323 GND.n5322 0.0344674
R17228 GND.n5322 GND.n1360 0.0344674
R17229 GND.n5318 GND.n1360 0.0344674
R17230 GND.n5318 GND.n5317 0.0344674
R17231 GND.n5317 GND.n5316 0.0344674
R17232 GND.n5316 GND.n1368 0.0344674
R17233 GND.n5312 GND.n1368 0.0344674
R17234 GND.n5312 GND.n5311 0.0344674
R17235 GND.n5311 GND.n5310 0.0344674
R17236 GND.n5310 GND.n1376 0.0344674
R17237 GND.n5306 GND.n1376 0.0344674
R17238 GND.n5306 GND.n5305 0.0344674
R17239 GND.n5305 GND.n5304 0.0344674
R17240 GND.n5304 GND.n1384 0.0344674
R17241 GND.n5300 GND.n1384 0.0344674
R17242 GND.n5300 GND.n5299 0.0344674
R17243 GND.n5299 GND.n5298 0.0344674
R17244 GND.n5298 GND.n1392 0.0344674
R17245 GND.n4962 GND.n4961 0.0336978
R17246 GND.n2932 GND.n2516 0.0336978
R17247 GND.n2938 GND.n2936 0.0336978
R17248 GND.n2937 GND.n2929 0.0336978
R17249 GND.n2945 GND.n2944 0.0336978
R17250 GND.n2930 GND.n2913 0.0336978
R17251 GND.n4521 GND.n4520 0.0336978
R17252 GND.n4524 GND.n2905 0.0336978
R17253 GND.n4525 GND.n2902 0.0336978
R17254 GND.n5221 GND.n1471 0.0336978
R17255 GND.n5218 GND.n5217 0.0336978
R17256 GND.n5214 GND.n1476 0.0336978
R17257 GND.n5213 GND.n1481 0.0336978
R17258 GND.n5210 GND.n5209 0.0336978
R17259 GND.n5206 GND.n1485 0.0336978
R17260 GND.n5205 GND.n1489 0.0336978
R17261 GND.n1499 GND.n1498 0.0336978
R17262 GND.n5196 GND.n5195 0.0336978
R17263 GND.n4962 GND.n2515 0.0123564
R17264 GND.n5222 GND.n5221 0.0123564
R17265 GND.n4961 GND.n2516 0.00117751
R17266 GND.n2936 GND.n2932 0.00117751
R17267 GND.n2938 GND.n2937 0.00117751
R17268 GND.n2945 GND.n2929 0.00117751
R17269 GND.n2944 GND.n2930 0.00117751
R17270 GND.n4520 GND.n2913 0.00117751
R17271 GND.n4521 GND.n2905 0.00117751
R17272 GND.n4525 GND.n4524 0.00117751
R17273 GND.n4528 GND.n2902 0.00117751
R17274 GND.n5218 GND.n1471 0.00117751
R17275 GND.n5217 GND.n1476 0.00117751
R17276 GND.n5214 GND.n5213 0.00117751
R17277 GND.n5210 GND.n1481 0.00117751
R17278 GND.n5209 GND.n1485 0.00117751
R17279 GND.n5206 GND.n5205 0.00117751
R17280 GND.n1498 GND.n1489 0.00117751
R17281 GND.n5196 GND.n1499 0.00117751
R17282 GND.n5195 GND.n1500 0.00117751
R17283 VP.n1 VP.t0 243.97
R17284 VP.n1 VP.t1 243.255
R17285 VP.n0 VP.t3 79.2009
R17286 VP.n0 VP.t2 58.4413
R17287 VP VP.n2 12.474
R17288 VP.n2 VP.n1 4.80222
R17289 VP.n2 VP.n0 0.972091
R17290 a_n5434_7417.n12 a_n5434_7417.t9 137.597
R17291 a_n5434_7417.n6 a_n5434_7417.t3 137.597
R17292 a_n5434_7417.n2 a_n5434_7417.t15 137.597
R17293 a_n5434_7417.n0 a_n5434_7417.t5 133.624
R17294 a_n5434_7417.n0 a_n5434_7417.t10 133.624
R17295 a_n5434_7417.n9 a_n5434_7417.t6 133.624
R17296 a_n5434_7417.n3 a_n5434_7417.t13 133.624
R17297 a_n5434_7417.n7 a_n5434_7417.t2 133.624
R17298 a_n5434_7417.n11 a_n5434_7417.n10 121.974
R17299 a_n5434_7417.n2 a_n5434_7417.n1 121.974
R17300 a_n5434_7417.n6 a_n5434_7417.n5 121.974
R17301 a_n5434_7417.n13 a_n5434_7417.n12 121.974
R17302 a_n5434_7417.n8 a_n5434_7417.n7 40.6178
R17303 a_n5434_7417.n4 a_n5434_7417.n3 13.8884
R17304 a_n5434_7417.n10 a_n5434_7417.t7 11.651
R17305 a_n5434_7417.n10 a_n5434_7417.t8 11.651
R17306 a_n5434_7417.n1 a_n5434_7417.t12 11.651
R17307 a_n5434_7417.n1 a_n5434_7417.t1 11.651
R17308 a_n5434_7417.n5 a_n5434_7417.t16 11.651
R17309 a_n5434_7417.n5 a_n5434_7417.t14 11.651
R17310 a_n5434_7417.t11 a_n5434_7417.n13 11.651
R17311 a_n5434_7417.n13 a_n5434_7417.t4 11.651
R17312 a_n5434_7417.n4 a_n5434_7417.t0 10.1951
R17313 a_n5434_7417.n9 a_n5434_7417.n8 7.46817
R17314 a_n5434_7417.n12 a_n5434_7417.n0 4.99188
R17315 a_n5434_7417.n3 a_n5434_7417.n2 3.97464
R17316 a_n5434_7417.n7 a_n5434_7417.n6 3.97464
R17317 a_n5434_7417.n11 a_n5434_7417.n9 3.97464
R17318 a_n5434_7417.n0 a_n5434_7417.n11 3.97464
R17319 a_n5434_7417.n8 a_n5434_7417.n4 2.44368
R17320 CS_BIAS.n215 CS_BIAS.n214 161.3
R17321 CS_BIAS.n213 CS_BIAS.n183 161.3
R17322 CS_BIAS.n212 CS_BIAS.n211 161.3
R17323 CS_BIAS.n210 CS_BIAS.n184 161.3
R17324 CS_BIAS.n209 CS_BIAS.n208 161.3
R17325 CS_BIAS.n207 CS_BIAS.n185 161.3
R17326 CS_BIAS.n206 CS_BIAS.n205 161.3
R17327 CS_BIAS.n204 CS_BIAS.n186 161.3
R17328 CS_BIAS.n203 CS_BIAS.n202 161.3
R17329 CS_BIAS.n201 CS_BIAS.n187 161.3
R17330 CS_BIAS.n200 CS_BIAS.n199 161.3
R17331 CS_BIAS.n198 CS_BIAS.n189 161.3
R17332 CS_BIAS.n197 CS_BIAS.n196 161.3
R17333 CS_BIAS.n195 CS_BIAS.n190 161.3
R17334 CS_BIAS.n194 CS_BIAS.n193 161.3
R17335 CS_BIAS.n158 CS_BIAS.n157 161.3
R17336 CS_BIAS.n159 CS_BIAS.n154 161.3
R17337 CS_BIAS.n161 CS_BIAS.n160 161.3
R17338 CS_BIAS.n162 CS_BIAS.n153 161.3
R17339 CS_BIAS.n164 CS_BIAS.n163 161.3
R17340 CS_BIAS.n165 CS_BIAS.n151 161.3
R17341 CS_BIAS.n167 CS_BIAS.n166 161.3
R17342 CS_BIAS.n168 CS_BIAS.n150 161.3
R17343 CS_BIAS.n170 CS_BIAS.n169 161.3
R17344 CS_BIAS.n171 CS_BIAS.n149 161.3
R17345 CS_BIAS.n173 CS_BIAS.n172 161.3
R17346 CS_BIAS.n174 CS_BIAS.n148 161.3
R17347 CS_BIAS.n176 CS_BIAS.n175 161.3
R17348 CS_BIAS.n177 CS_BIAS.n147 161.3
R17349 CS_BIAS.n179 CS_BIAS.n178 161.3
R17350 CS_BIAS.n122 CS_BIAS.n121 161.3
R17351 CS_BIAS.n123 CS_BIAS.n118 161.3
R17352 CS_BIAS.n125 CS_BIAS.n124 161.3
R17353 CS_BIAS.n126 CS_BIAS.n117 161.3
R17354 CS_BIAS.n128 CS_BIAS.n127 161.3
R17355 CS_BIAS.n129 CS_BIAS.n115 161.3
R17356 CS_BIAS.n131 CS_BIAS.n130 161.3
R17357 CS_BIAS.n132 CS_BIAS.n114 161.3
R17358 CS_BIAS.n134 CS_BIAS.n133 161.3
R17359 CS_BIAS.n135 CS_BIAS.n113 161.3
R17360 CS_BIAS.n137 CS_BIAS.n136 161.3
R17361 CS_BIAS.n138 CS_BIAS.n112 161.3
R17362 CS_BIAS.n140 CS_BIAS.n139 161.3
R17363 CS_BIAS.n141 CS_BIAS.n111 161.3
R17364 CS_BIAS.n143 CS_BIAS.n142 161.3
R17365 CS_BIAS.n86 CS_BIAS.n85 161.3
R17366 CS_BIAS.n87 CS_BIAS.n82 161.3
R17367 CS_BIAS.n89 CS_BIAS.n88 161.3
R17368 CS_BIAS.n90 CS_BIAS.n81 161.3
R17369 CS_BIAS.n92 CS_BIAS.n91 161.3
R17370 CS_BIAS.n93 CS_BIAS.n79 161.3
R17371 CS_BIAS.n95 CS_BIAS.n94 161.3
R17372 CS_BIAS.n96 CS_BIAS.n78 161.3
R17373 CS_BIAS.n98 CS_BIAS.n97 161.3
R17374 CS_BIAS.n99 CS_BIAS.n77 161.3
R17375 CS_BIAS.n101 CS_BIAS.n100 161.3
R17376 CS_BIAS.n102 CS_BIAS.n76 161.3
R17377 CS_BIAS.n104 CS_BIAS.n103 161.3
R17378 CS_BIAS.n105 CS_BIAS.n75 161.3
R17379 CS_BIAS.n107 CS_BIAS.n106 161.3
R17380 CS_BIAS.n20 CS_BIAS.n19 161.3
R17381 CS_BIAS.n21 CS_BIAS.n16 161.3
R17382 CS_BIAS.n23 CS_BIAS.n22 161.3
R17383 CS_BIAS.n24 CS_BIAS.n15 161.3
R17384 CS_BIAS.n26 CS_BIAS.n25 161.3
R17385 CS_BIAS.n27 CS_BIAS.n13 161.3
R17386 CS_BIAS.n29 CS_BIAS.n28 161.3
R17387 CS_BIAS.n30 CS_BIAS.n12 161.3
R17388 CS_BIAS.n32 CS_BIAS.n31 161.3
R17389 CS_BIAS.n33 CS_BIAS.n11 161.3
R17390 CS_BIAS.n35 CS_BIAS.n34 161.3
R17391 CS_BIAS.n36 CS_BIAS.n10 161.3
R17392 CS_BIAS.n38 CS_BIAS.n37 161.3
R17393 CS_BIAS.n39 CS_BIAS.n9 161.3
R17394 CS_BIAS.n41 CS_BIAS.n40 161.3
R17395 CS_BIAS.n51 CS_BIAS.n50 161.3
R17396 CS_BIAS.n52 CS_BIAS.n47 161.3
R17397 CS_BIAS.n54 CS_BIAS.n53 161.3
R17398 CS_BIAS.n55 CS_BIAS.n7 161.3
R17399 CS_BIAS.n57 CS_BIAS.n56 161.3
R17400 CS_BIAS.n58 CS_BIAS.n5 161.3
R17401 CS_BIAS.n60 CS_BIAS.n59 161.3
R17402 CS_BIAS.n61 CS_BIAS.n4 161.3
R17403 CS_BIAS.n63 CS_BIAS.n62 161.3
R17404 CS_BIAS.n64 CS_BIAS.n3 161.3
R17405 CS_BIAS.n66 CS_BIAS.n65 161.3
R17406 CS_BIAS.n67 CS_BIAS.n2 161.3
R17407 CS_BIAS.n69 CS_BIAS.n68 161.3
R17408 CS_BIAS.n70 CS_BIAS.n1 161.3
R17409 CS_BIAS.n72 CS_BIAS.n71 161.3
R17410 CS_BIAS.n433 CS_BIAS.n432 161.3
R17411 CS_BIAS.n431 CS_BIAS.n401 161.3
R17412 CS_BIAS.n430 CS_BIAS.n429 161.3
R17413 CS_BIAS.n428 CS_BIAS.n402 161.3
R17414 CS_BIAS.n427 CS_BIAS.n426 161.3
R17415 CS_BIAS.n425 CS_BIAS.n403 161.3
R17416 CS_BIAS.n424 CS_BIAS.n423 161.3
R17417 CS_BIAS.n422 CS_BIAS.n404 161.3
R17418 CS_BIAS.n421 CS_BIAS.n420 161.3
R17419 CS_BIAS.n418 CS_BIAS.n405 161.3
R17420 CS_BIAS.n417 CS_BIAS.n416 161.3
R17421 CS_BIAS.n415 CS_BIAS.n406 161.3
R17422 CS_BIAS.n414 CS_BIAS.n413 161.3
R17423 CS_BIAS.n412 CS_BIAS.n407 161.3
R17424 CS_BIAS.n411 CS_BIAS.n410 161.3
R17425 CS_BIAS.n397 CS_BIAS.n396 161.3
R17426 CS_BIAS.n395 CS_BIAS.n365 161.3
R17427 CS_BIAS.n394 CS_BIAS.n393 161.3
R17428 CS_BIAS.n392 CS_BIAS.n366 161.3
R17429 CS_BIAS.n391 CS_BIAS.n390 161.3
R17430 CS_BIAS.n389 CS_BIAS.n367 161.3
R17431 CS_BIAS.n388 CS_BIAS.n387 161.3
R17432 CS_BIAS.n386 CS_BIAS.n368 161.3
R17433 CS_BIAS.n385 CS_BIAS.n384 161.3
R17434 CS_BIAS.n382 CS_BIAS.n369 161.3
R17435 CS_BIAS.n381 CS_BIAS.n380 161.3
R17436 CS_BIAS.n379 CS_BIAS.n370 161.3
R17437 CS_BIAS.n378 CS_BIAS.n377 161.3
R17438 CS_BIAS.n376 CS_BIAS.n371 161.3
R17439 CS_BIAS.n375 CS_BIAS.n374 161.3
R17440 CS_BIAS.n361 CS_BIAS.n360 161.3
R17441 CS_BIAS.n359 CS_BIAS.n329 161.3
R17442 CS_BIAS.n358 CS_BIAS.n357 161.3
R17443 CS_BIAS.n356 CS_BIAS.n330 161.3
R17444 CS_BIAS.n355 CS_BIAS.n354 161.3
R17445 CS_BIAS.n353 CS_BIAS.n331 161.3
R17446 CS_BIAS.n352 CS_BIAS.n351 161.3
R17447 CS_BIAS.n350 CS_BIAS.n332 161.3
R17448 CS_BIAS.n349 CS_BIAS.n348 161.3
R17449 CS_BIAS.n346 CS_BIAS.n333 161.3
R17450 CS_BIAS.n345 CS_BIAS.n344 161.3
R17451 CS_BIAS.n343 CS_BIAS.n334 161.3
R17452 CS_BIAS.n342 CS_BIAS.n341 161.3
R17453 CS_BIAS.n340 CS_BIAS.n335 161.3
R17454 CS_BIAS.n339 CS_BIAS.n338 161.3
R17455 CS_BIAS.n325 CS_BIAS.n324 161.3
R17456 CS_BIAS.n323 CS_BIAS.n293 161.3
R17457 CS_BIAS.n322 CS_BIAS.n321 161.3
R17458 CS_BIAS.n320 CS_BIAS.n294 161.3
R17459 CS_BIAS.n319 CS_BIAS.n318 161.3
R17460 CS_BIAS.n317 CS_BIAS.n295 161.3
R17461 CS_BIAS.n316 CS_BIAS.n315 161.3
R17462 CS_BIAS.n314 CS_BIAS.n296 161.3
R17463 CS_BIAS.n313 CS_BIAS.n312 161.3
R17464 CS_BIAS.n310 CS_BIAS.n297 161.3
R17465 CS_BIAS.n309 CS_BIAS.n308 161.3
R17466 CS_BIAS.n307 CS_BIAS.n298 161.3
R17467 CS_BIAS.n306 CS_BIAS.n305 161.3
R17468 CS_BIAS.n304 CS_BIAS.n299 161.3
R17469 CS_BIAS.n303 CS_BIAS.n302 161.3
R17470 CS_BIAS.n267 CS_BIAS.n266 161.3
R17471 CS_BIAS.n265 CS_BIAS.n235 161.3
R17472 CS_BIAS.n264 CS_BIAS.n263 161.3
R17473 CS_BIAS.n262 CS_BIAS.n236 161.3
R17474 CS_BIAS.n261 CS_BIAS.n260 161.3
R17475 CS_BIAS.n259 CS_BIAS.n237 161.3
R17476 CS_BIAS.n258 CS_BIAS.n257 161.3
R17477 CS_BIAS.n256 CS_BIAS.n238 161.3
R17478 CS_BIAS.n255 CS_BIAS.n254 161.3
R17479 CS_BIAS.n252 CS_BIAS.n239 161.3
R17480 CS_BIAS.n251 CS_BIAS.n250 161.3
R17481 CS_BIAS.n249 CS_BIAS.n240 161.3
R17482 CS_BIAS.n248 CS_BIAS.n247 161.3
R17483 CS_BIAS.n246 CS_BIAS.n241 161.3
R17484 CS_BIAS.n245 CS_BIAS.n244 161.3
R17485 CS_BIAS.n232 CS_BIAS.n231 161.3
R17486 CS_BIAS.n230 CS_BIAS.n225 161.3
R17487 CS_BIAS.n229 CS_BIAS.n228 161.3
R17488 CS_BIAS.n272 CS_BIAS.n224 161.3
R17489 CS_BIAS.n290 CS_BIAS.n289 161.3
R17490 CS_BIAS.n288 CS_BIAS.n219 161.3
R17491 CS_BIAS.n287 CS_BIAS.n286 161.3
R17492 CS_BIAS.n285 CS_BIAS.n220 161.3
R17493 CS_BIAS.n284 CS_BIAS.n283 161.3
R17494 CS_BIAS.n282 CS_BIAS.n221 161.3
R17495 CS_BIAS.n281 CS_BIAS.n280 161.3
R17496 CS_BIAS.n279 CS_BIAS.n222 161.3
R17497 CS_BIAS.n278 CS_BIAS.n277 161.3
R17498 CS_BIAS.n275 CS_BIAS.n223 161.3
R17499 CS_BIAS.n274 CS_BIAS.n273 161.3
R17500 CS_BIAS.n46 CS_BIAS.n45 86.5843
R17501 CS_BIAS.n271 CS_BIAS.n233 86.5843
R17502 CS_BIAS.n44 CS_BIAS.n43 84.9593
R17503 CS_BIAS.n270 CS_BIAS.n269 84.9593
R17504 CS_BIAS.n216 CS_BIAS.n182 77.4578
R17505 CS_BIAS.n180 CS_BIAS.n146 77.4578
R17506 CS_BIAS.n144 CS_BIAS.n110 77.4578
R17507 CS_BIAS.n108 CS_BIAS.n74 77.4578
R17508 CS_BIAS.n42 CS_BIAS.n8 77.4578
R17509 CS_BIAS.n73 CS_BIAS.n0 77.4578
R17510 CS_BIAS.n434 CS_BIAS.n400 77.4578
R17511 CS_BIAS.n398 CS_BIAS.n364 77.4578
R17512 CS_BIAS.n362 CS_BIAS.n328 77.4578
R17513 CS_BIAS.n326 CS_BIAS.n292 77.4578
R17514 CS_BIAS.n268 CS_BIAS.n234 77.4578
R17515 CS_BIAS.n291 CS_BIAS.n218 77.4578
R17516 CS_BIAS.n208 CS_BIAS.n184 56.0773
R17517 CS_BIAS.n172 CS_BIAS.n148 56.0773
R17518 CS_BIAS.n136 CS_BIAS.n112 56.0773
R17519 CS_BIAS.n100 CS_BIAS.n76 56.0773
R17520 CS_BIAS.n34 CS_BIAS.n10 56.0773
R17521 CS_BIAS.n65 CS_BIAS.n2 56.0773
R17522 CS_BIAS.n426 CS_BIAS.n402 56.0773
R17523 CS_BIAS.n390 CS_BIAS.n366 56.0773
R17524 CS_BIAS.n354 CS_BIAS.n330 56.0773
R17525 CS_BIAS.n318 CS_BIAS.n294 56.0773
R17526 CS_BIAS.n260 CS_BIAS.n236 56.0773
R17527 CS_BIAS.n283 CS_BIAS.n220 56.0773
R17528 CS_BIAS.n156 CS_BIAS.n155 54.2621
R17529 CS_BIAS.n120 CS_BIAS.n119 54.2621
R17530 CS_BIAS.n84 CS_BIAS.n83 54.2621
R17531 CS_BIAS.n18 CS_BIAS.n17 54.2621
R17532 CS_BIAS.n49 CS_BIAS.n48 54.2621
R17533 CS_BIAS.n192 CS_BIAS.n191 54.2621
R17534 CS_BIAS.n409 CS_BIAS.n408 54.2621
R17535 CS_BIAS.n373 CS_BIAS.n372 54.2621
R17536 CS_BIAS.n337 CS_BIAS.n336 54.2621
R17537 CS_BIAS.n301 CS_BIAS.n300 54.2621
R17538 CS_BIAS.n243 CS_BIAS.n242 54.2621
R17539 CS_BIAS.n227 CS_BIAS.n226 54.2621
R17540 CS_BIAS.n192 CS_BIAS.t20 50.3417
R17541 CS_BIAS.n409 CS_BIAS.t46 50.3417
R17542 CS_BIAS.n373 CS_BIAS.t40 50.3417
R17543 CS_BIAS.n337 CS_BIAS.t50 50.3417
R17544 CS_BIAS.n301 CS_BIAS.t18 50.3417
R17545 CS_BIAS.n243 CS_BIAS.t10 50.3417
R17546 CS_BIAS.n227 CS_BIAS.t23 50.3417
R17547 CS_BIAS.n156 CS_BIAS.t55 50.3415
R17548 CS_BIAS.n120 CS_BIAS.t39 50.3415
R17549 CS_BIAS.n84 CS_BIAS.t35 50.3415
R17550 CS_BIAS.n18 CS_BIAS.t2 50.3415
R17551 CS_BIAS.n49 CS_BIAS.t44 50.3415
R17552 CS_BIAS.n196 CS_BIAS.n189 40.577
R17553 CS_BIAS.n200 CS_BIAS.n189 40.577
R17554 CS_BIAS.n164 CS_BIAS.n153 40.577
R17555 CS_BIAS.n160 CS_BIAS.n153 40.577
R17556 CS_BIAS.n128 CS_BIAS.n117 40.577
R17557 CS_BIAS.n124 CS_BIAS.n117 40.577
R17558 CS_BIAS.n92 CS_BIAS.n81 40.577
R17559 CS_BIAS.n88 CS_BIAS.n81 40.577
R17560 CS_BIAS.n26 CS_BIAS.n15 40.577
R17561 CS_BIAS.n22 CS_BIAS.n15 40.577
R17562 CS_BIAS.n57 CS_BIAS.n7 40.577
R17563 CS_BIAS.n53 CS_BIAS.n7 40.577
R17564 CS_BIAS.n413 CS_BIAS.n406 40.577
R17565 CS_BIAS.n417 CS_BIAS.n406 40.577
R17566 CS_BIAS.n377 CS_BIAS.n370 40.577
R17567 CS_BIAS.n381 CS_BIAS.n370 40.577
R17568 CS_BIAS.n341 CS_BIAS.n334 40.577
R17569 CS_BIAS.n345 CS_BIAS.n334 40.577
R17570 CS_BIAS.n305 CS_BIAS.n298 40.577
R17571 CS_BIAS.n309 CS_BIAS.n298 40.577
R17572 CS_BIAS.n247 CS_BIAS.n240 40.577
R17573 CS_BIAS.n251 CS_BIAS.n240 40.577
R17574 CS_BIAS.n274 CS_BIAS.n224 40.577
R17575 CS_BIAS.n231 CS_BIAS.n224 40.577
R17576 CS_BIAS.n212 CS_BIAS.n184 25.0767
R17577 CS_BIAS.n176 CS_BIAS.n148 25.0767
R17578 CS_BIAS.n140 CS_BIAS.n112 25.0767
R17579 CS_BIAS.n104 CS_BIAS.n76 25.0767
R17580 CS_BIAS.n38 CS_BIAS.n10 25.0767
R17581 CS_BIAS.n69 CS_BIAS.n2 25.0767
R17582 CS_BIAS.n430 CS_BIAS.n402 25.0767
R17583 CS_BIAS.n394 CS_BIAS.n366 25.0767
R17584 CS_BIAS.n358 CS_BIAS.n330 25.0767
R17585 CS_BIAS.n322 CS_BIAS.n294 25.0767
R17586 CS_BIAS.n264 CS_BIAS.n236 25.0767
R17587 CS_BIAS.n287 CS_BIAS.n220 25.0767
R17588 CS_BIAS.n196 CS_BIAS.n195 24.5923
R17589 CS_BIAS.n195 CS_BIAS.n194 24.5923
R17590 CS_BIAS.n208 CS_BIAS.n207 24.5923
R17591 CS_BIAS.n207 CS_BIAS.n206 24.5923
R17592 CS_BIAS.n206 CS_BIAS.n186 24.5923
R17593 CS_BIAS.n202 CS_BIAS.n201 24.5923
R17594 CS_BIAS.n201 CS_BIAS.n200 24.5923
R17595 CS_BIAS.n214 CS_BIAS.n213 24.5923
R17596 CS_BIAS.n213 CS_BIAS.n212 24.5923
R17597 CS_BIAS.n178 CS_BIAS.n177 24.5923
R17598 CS_BIAS.n177 CS_BIAS.n176 24.5923
R17599 CS_BIAS.n172 CS_BIAS.n171 24.5923
R17600 CS_BIAS.n171 CS_BIAS.n170 24.5923
R17601 CS_BIAS.n170 CS_BIAS.n150 24.5923
R17602 CS_BIAS.n166 CS_BIAS.n165 24.5923
R17603 CS_BIAS.n165 CS_BIAS.n164 24.5923
R17604 CS_BIAS.n160 CS_BIAS.n159 24.5923
R17605 CS_BIAS.n159 CS_BIAS.n158 24.5923
R17606 CS_BIAS.n142 CS_BIAS.n141 24.5923
R17607 CS_BIAS.n141 CS_BIAS.n140 24.5923
R17608 CS_BIAS.n136 CS_BIAS.n135 24.5923
R17609 CS_BIAS.n135 CS_BIAS.n134 24.5923
R17610 CS_BIAS.n134 CS_BIAS.n114 24.5923
R17611 CS_BIAS.n130 CS_BIAS.n129 24.5923
R17612 CS_BIAS.n129 CS_BIAS.n128 24.5923
R17613 CS_BIAS.n124 CS_BIAS.n123 24.5923
R17614 CS_BIAS.n123 CS_BIAS.n122 24.5923
R17615 CS_BIAS.n106 CS_BIAS.n105 24.5923
R17616 CS_BIAS.n105 CS_BIAS.n104 24.5923
R17617 CS_BIAS.n100 CS_BIAS.n99 24.5923
R17618 CS_BIAS.n99 CS_BIAS.n98 24.5923
R17619 CS_BIAS.n98 CS_BIAS.n78 24.5923
R17620 CS_BIAS.n94 CS_BIAS.n93 24.5923
R17621 CS_BIAS.n93 CS_BIAS.n92 24.5923
R17622 CS_BIAS.n88 CS_BIAS.n87 24.5923
R17623 CS_BIAS.n87 CS_BIAS.n86 24.5923
R17624 CS_BIAS.n40 CS_BIAS.n39 24.5923
R17625 CS_BIAS.n39 CS_BIAS.n38 24.5923
R17626 CS_BIAS.n34 CS_BIAS.n33 24.5923
R17627 CS_BIAS.n33 CS_BIAS.n32 24.5923
R17628 CS_BIAS.n32 CS_BIAS.n12 24.5923
R17629 CS_BIAS.n28 CS_BIAS.n27 24.5923
R17630 CS_BIAS.n27 CS_BIAS.n26 24.5923
R17631 CS_BIAS.n22 CS_BIAS.n21 24.5923
R17632 CS_BIAS.n21 CS_BIAS.n20 24.5923
R17633 CS_BIAS.n71 CS_BIAS.n70 24.5923
R17634 CS_BIAS.n70 CS_BIAS.n69 24.5923
R17635 CS_BIAS.n65 CS_BIAS.n64 24.5923
R17636 CS_BIAS.n64 CS_BIAS.n63 24.5923
R17637 CS_BIAS.n63 CS_BIAS.n4 24.5923
R17638 CS_BIAS.n59 CS_BIAS.n58 24.5923
R17639 CS_BIAS.n58 CS_BIAS.n57 24.5923
R17640 CS_BIAS.n53 CS_BIAS.n52 24.5923
R17641 CS_BIAS.n52 CS_BIAS.n51 24.5923
R17642 CS_BIAS.n412 CS_BIAS.n411 24.5923
R17643 CS_BIAS.n413 CS_BIAS.n412 24.5923
R17644 CS_BIAS.n418 CS_BIAS.n417 24.5923
R17645 CS_BIAS.n420 CS_BIAS.n418 24.5923
R17646 CS_BIAS.n424 CS_BIAS.n404 24.5923
R17647 CS_BIAS.n425 CS_BIAS.n424 24.5923
R17648 CS_BIAS.n426 CS_BIAS.n425 24.5923
R17649 CS_BIAS.n431 CS_BIAS.n430 24.5923
R17650 CS_BIAS.n432 CS_BIAS.n431 24.5923
R17651 CS_BIAS.n376 CS_BIAS.n375 24.5923
R17652 CS_BIAS.n377 CS_BIAS.n376 24.5923
R17653 CS_BIAS.n382 CS_BIAS.n381 24.5923
R17654 CS_BIAS.n384 CS_BIAS.n382 24.5923
R17655 CS_BIAS.n388 CS_BIAS.n368 24.5923
R17656 CS_BIAS.n389 CS_BIAS.n388 24.5923
R17657 CS_BIAS.n390 CS_BIAS.n389 24.5923
R17658 CS_BIAS.n395 CS_BIAS.n394 24.5923
R17659 CS_BIAS.n396 CS_BIAS.n395 24.5923
R17660 CS_BIAS.n340 CS_BIAS.n339 24.5923
R17661 CS_BIAS.n341 CS_BIAS.n340 24.5923
R17662 CS_BIAS.n346 CS_BIAS.n345 24.5923
R17663 CS_BIAS.n348 CS_BIAS.n346 24.5923
R17664 CS_BIAS.n352 CS_BIAS.n332 24.5923
R17665 CS_BIAS.n353 CS_BIAS.n352 24.5923
R17666 CS_BIAS.n354 CS_BIAS.n353 24.5923
R17667 CS_BIAS.n359 CS_BIAS.n358 24.5923
R17668 CS_BIAS.n360 CS_BIAS.n359 24.5923
R17669 CS_BIAS.n304 CS_BIAS.n303 24.5923
R17670 CS_BIAS.n305 CS_BIAS.n304 24.5923
R17671 CS_BIAS.n310 CS_BIAS.n309 24.5923
R17672 CS_BIAS.n312 CS_BIAS.n310 24.5923
R17673 CS_BIAS.n316 CS_BIAS.n296 24.5923
R17674 CS_BIAS.n317 CS_BIAS.n316 24.5923
R17675 CS_BIAS.n318 CS_BIAS.n317 24.5923
R17676 CS_BIAS.n323 CS_BIAS.n322 24.5923
R17677 CS_BIAS.n324 CS_BIAS.n323 24.5923
R17678 CS_BIAS.n246 CS_BIAS.n245 24.5923
R17679 CS_BIAS.n247 CS_BIAS.n246 24.5923
R17680 CS_BIAS.n252 CS_BIAS.n251 24.5923
R17681 CS_BIAS.n254 CS_BIAS.n252 24.5923
R17682 CS_BIAS.n258 CS_BIAS.n238 24.5923
R17683 CS_BIAS.n259 CS_BIAS.n258 24.5923
R17684 CS_BIAS.n260 CS_BIAS.n259 24.5923
R17685 CS_BIAS.n265 CS_BIAS.n264 24.5923
R17686 CS_BIAS.n266 CS_BIAS.n265 24.5923
R17687 CS_BIAS.n288 CS_BIAS.n287 24.5923
R17688 CS_BIAS.n289 CS_BIAS.n288 24.5923
R17689 CS_BIAS.n275 CS_BIAS.n274 24.5923
R17690 CS_BIAS.n277 CS_BIAS.n275 24.5923
R17691 CS_BIAS.n281 CS_BIAS.n222 24.5923
R17692 CS_BIAS.n282 CS_BIAS.n281 24.5923
R17693 CS_BIAS.n283 CS_BIAS.n282 24.5923
R17694 CS_BIAS.n230 CS_BIAS.n229 24.5923
R17695 CS_BIAS.n231 CS_BIAS.n230 24.5923
R17696 CS_BIAS.n194 CS_BIAS.n191 20.6576
R17697 CS_BIAS.n202 CS_BIAS.n188 20.6576
R17698 CS_BIAS.n166 CS_BIAS.n152 20.6576
R17699 CS_BIAS.n158 CS_BIAS.n155 20.6576
R17700 CS_BIAS.n130 CS_BIAS.n116 20.6576
R17701 CS_BIAS.n122 CS_BIAS.n119 20.6576
R17702 CS_BIAS.n94 CS_BIAS.n80 20.6576
R17703 CS_BIAS.n86 CS_BIAS.n83 20.6576
R17704 CS_BIAS.n28 CS_BIAS.n14 20.6576
R17705 CS_BIAS.n20 CS_BIAS.n17 20.6576
R17706 CS_BIAS.n59 CS_BIAS.n6 20.6576
R17707 CS_BIAS.n51 CS_BIAS.n48 20.6576
R17708 CS_BIAS.n411 CS_BIAS.n408 20.6576
R17709 CS_BIAS.n420 CS_BIAS.n419 20.6576
R17710 CS_BIAS.n375 CS_BIAS.n372 20.6576
R17711 CS_BIAS.n384 CS_BIAS.n383 20.6576
R17712 CS_BIAS.n339 CS_BIAS.n336 20.6576
R17713 CS_BIAS.n348 CS_BIAS.n347 20.6576
R17714 CS_BIAS.n303 CS_BIAS.n300 20.6576
R17715 CS_BIAS.n312 CS_BIAS.n311 20.6576
R17716 CS_BIAS.n245 CS_BIAS.n242 20.6576
R17717 CS_BIAS.n254 CS_BIAS.n253 20.6576
R17718 CS_BIAS.n277 CS_BIAS.n276 20.6576
R17719 CS_BIAS.n229 CS_BIAS.n226 20.6576
R17720 CS_BIAS.n191 CS_BIAS.t32 16.4791
R17721 CS_BIAS.n188 CS_BIAS.t28 16.4791
R17722 CS_BIAS.n182 CS_BIAS.t51 16.4791
R17723 CS_BIAS.n146 CS_BIAS.t45 16.4791
R17724 CS_BIAS.n152 CS_BIAS.t22 16.4791
R17725 CS_BIAS.n155 CS_BIAS.t24 16.4791
R17726 CS_BIAS.n110 CS_BIAS.t26 16.4791
R17727 CS_BIAS.n116 CS_BIAS.t27 16.4791
R17728 CS_BIAS.n119 CS_BIAS.t49 16.4791
R17729 CS_BIAS.n74 CS_BIAS.t21 16.4791
R17730 CS_BIAS.n80 CS_BIAS.t38 16.4791
R17731 CS_BIAS.n83 CS_BIAS.t42 16.4791
R17732 CS_BIAS.n8 CS_BIAS.t12 16.4791
R17733 CS_BIAS.n14 CS_BIAS.t6 16.4791
R17734 CS_BIAS.n17 CS_BIAS.t0 16.4791
R17735 CS_BIAS.n0 CS_BIAS.t16 16.4791
R17736 CS_BIAS.n6 CS_BIAS.t41 16.4791
R17737 CS_BIAS.n48 CS_BIAS.t48 16.4791
R17738 CS_BIAS.n408 CS_BIAS.t54 16.4791
R17739 CS_BIAS.n419 CS_BIAS.t25 16.4791
R17740 CS_BIAS.n400 CS_BIAS.t34 16.4791
R17741 CS_BIAS.n372 CS_BIAS.t52 16.4791
R17742 CS_BIAS.n383 CS_BIAS.t19 16.4791
R17743 CS_BIAS.n364 CS_BIAS.t31 16.4791
R17744 CS_BIAS.n336 CS_BIAS.t17 16.4791
R17745 CS_BIAS.n347 CS_BIAS.t29 16.4791
R17746 CS_BIAS.n328 CS_BIAS.t36 16.4791
R17747 CS_BIAS.n300 CS_BIAS.t30 16.4791
R17748 CS_BIAS.n311 CS_BIAS.t37 16.4791
R17749 CS_BIAS.n292 CS_BIAS.t47 16.4791
R17750 CS_BIAS.n242 CS_BIAS.t4 16.4791
R17751 CS_BIAS.n253 CS_BIAS.t8 16.4791
R17752 CS_BIAS.n234 CS_BIAS.t14 16.4791
R17753 CS_BIAS.n218 CS_BIAS.t53 16.4791
R17754 CS_BIAS.n276 CS_BIAS.t33 16.4791
R17755 CS_BIAS.n226 CS_BIAS.t43 16.4791
R17756 CS_BIAS.n44 CS_BIAS.n42 13.1696
R17757 CS_BIAS.n270 CS_BIAS.n268 13.1696
R17758 CS_BIAS.n214 CS_BIAS.n182 12.7883
R17759 CS_BIAS.n178 CS_BIAS.n146 12.7883
R17760 CS_BIAS.n142 CS_BIAS.n110 12.7883
R17761 CS_BIAS.n106 CS_BIAS.n74 12.7883
R17762 CS_BIAS.n40 CS_BIAS.n8 12.7883
R17763 CS_BIAS.n71 CS_BIAS.n0 12.7883
R17764 CS_BIAS.n432 CS_BIAS.n400 12.7883
R17765 CS_BIAS.n396 CS_BIAS.n364 12.7883
R17766 CS_BIAS.n360 CS_BIAS.n328 12.7883
R17767 CS_BIAS.n324 CS_BIAS.n292 12.7883
R17768 CS_BIAS.n266 CS_BIAS.n234 12.7883
R17769 CS_BIAS.n289 CS_BIAS.n218 12.7883
R17770 CS_BIAS.n55 CS_BIAS.n46 9.50363
R17771 CS_BIAS.n272 CS_BIAS.n271 9.50363
R17772 CS_BIAS.n436 CS_BIAS.n217 8.38478
R17773 CS_BIAS.n45 CS_BIAS.t1 8.2505
R17774 CS_BIAS.n45 CS_BIAS.t3 8.2505
R17775 CS_BIAS.n43 CS_BIAS.t13 8.2505
R17776 CS_BIAS.n43 CS_BIAS.t7 8.2505
R17777 CS_BIAS.n269 CS_BIAS.t9 8.2505
R17778 CS_BIAS.n269 CS_BIAS.t15 8.2505
R17779 CS_BIAS.n233 CS_BIAS.t11 8.2505
R17780 CS_BIAS.n233 CS_BIAS.t5 8.2505
R17781 CS_BIAS.n109 CS_BIAS.n73 6.92995
R17782 CS_BIAS.n327 CS_BIAS.n291 6.92995
R17783 CS_BIAS.n436 CS_BIAS.n435 6.0658
R17784 CS_BIAS.n217 CS_BIAS.n216 5.20078
R17785 CS_BIAS.n181 CS_BIAS.n180 5.20078
R17786 CS_BIAS.n145 CS_BIAS.n144 5.20078
R17787 CS_BIAS.n109 CS_BIAS.n108 5.20078
R17788 CS_BIAS.n435 CS_BIAS.n434 5.20078
R17789 CS_BIAS.n399 CS_BIAS.n398 5.20078
R17790 CS_BIAS.n363 CS_BIAS.n362 5.20078
R17791 CS_BIAS.n327 CS_BIAS.n326 5.20078
R17792 CS_BIAS.n188 CS_BIAS.n186 3.93519
R17793 CS_BIAS.n152 CS_BIAS.n150 3.93519
R17794 CS_BIAS.n116 CS_BIAS.n114 3.93519
R17795 CS_BIAS.n80 CS_BIAS.n78 3.93519
R17796 CS_BIAS.n14 CS_BIAS.n12 3.93519
R17797 CS_BIAS.n6 CS_BIAS.n4 3.93519
R17798 CS_BIAS.n419 CS_BIAS.n404 3.93519
R17799 CS_BIAS.n383 CS_BIAS.n368 3.93519
R17800 CS_BIAS.n347 CS_BIAS.n332 3.93519
R17801 CS_BIAS.n311 CS_BIAS.n296 3.93519
R17802 CS_BIAS.n253 CS_BIAS.n238 3.93519
R17803 CS_BIAS.n276 CS_BIAS.n222 3.93519
R17804 CS_BIAS CS_BIAS.n436 3.91321
R17805 CS_BIAS.n193 CS_BIAS.n192 3.05448
R17806 CS_BIAS.n410 CS_BIAS.n409 3.05448
R17807 CS_BIAS.n374 CS_BIAS.n373 3.05448
R17808 CS_BIAS.n338 CS_BIAS.n337 3.05448
R17809 CS_BIAS.n302 CS_BIAS.n301 3.05448
R17810 CS_BIAS.n244 CS_BIAS.n243 3.05448
R17811 CS_BIAS.n228 CS_BIAS.n227 3.05448
R17812 CS_BIAS.n157 CS_BIAS.n156 3.05446
R17813 CS_BIAS.n121 CS_BIAS.n120 3.05446
R17814 CS_BIAS.n85 CS_BIAS.n84 3.05446
R17815 CS_BIAS.n19 CS_BIAS.n18 3.05446
R17816 CS_BIAS.n50 CS_BIAS.n49 3.05446
R17817 CS_BIAS.n145 CS_BIAS.n109 1.72967
R17818 CS_BIAS.n181 CS_BIAS.n145 1.72967
R17819 CS_BIAS.n217 CS_BIAS.n181 1.72967
R17820 CS_BIAS.n363 CS_BIAS.n327 1.72967
R17821 CS_BIAS.n399 CS_BIAS.n363 1.72967
R17822 CS_BIAS.n435 CS_BIAS.n399 1.72967
R17823 CS_BIAS.n46 CS_BIAS.n44 1.6255
R17824 CS_BIAS.n271 CS_BIAS.n270 1.6255
R17825 CS_BIAS.n216 CS_BIAS.n215 0.354861
R17826 CS_BIAS.n180 CS_BIAS.n179 0.354861
R17827 CS_BIAS.n144 CS_BIAS.n143 0.354861
R17828 CS_BIAS.n108 CS_BIAS.n107 0.354861
R17829 CS_BIAS.n42 CS_BIAS.n41 0.354861
R17830 CS_BIAS.n73 CS_BIAS.n72 0.354861
R17831 CS_BIAS.n434 CS_BIAS.n433 0.354861
R17832 CS_BIAS.n398 CS_BIAS.n397 0.354861
R17833 CS_BIAS.n362 CS_BIAS.n361 0.354861
R17834 CS_BIAS.n326 CS_BIAS.n325 0.354861
R17835 CS_BIAS.n268 CS_BIAS.n267 0.354861
R17836 CS_BIAS.n291 CS_BIAS.n290 0.354861
R17837 CS_BIAS.n215 CS_BIAS.n183 0.189894
R17838 CS_BIAS.n211 CS_BIAS.n183 0.189894
R17839 CS_BIAS.n211 CS_BIAS.n210 0.189894
R17840 CS_BIAS.n210 CS_BIAS.n209 0.189894
R17841 CS_BIAS.n209 CS_BIAS.n185 0.189894
R17842 CS_BIAS.n205 CS_BIAS.n185 0.189894
R17843 CS_BIAS.n205 CS_BIAS.n204 0.189894
R17844 CS_BIAS.n204 CS_BIAS.n203 0.189894
R17845 CS_BIAS.n203 CS_BIAS.n187 0.189894
R17846 CS_BIAS.n199 CS_BIAS.n187 0.189894
R17847 CS_BIAS.n199 CS_BIAS.n198 0.189894
R17848 CS_BIAS.n198 CS_BIAS.n197 0.189894
R17849 CS_BIAS.n197 CS_BIAS.n190 0.189894
R17850 CS_BIAS.n193 CS_BIAS.n190 0.189894
R17851 CS_BIAS.n179 CS_BIAS.n147 0.189894
R17852 CS_BIAS.n175 CS_BIAS.n147 0.189894
R17853 CS_BIAS.n175 CS_BIAS.n174 0.189894
R17854 CS_BIAS.n174 CS_BIAS.n173 0.189894
R17855 CS_BIAS.n173 CS_BIAS.n149 0.189894
R17856 CS_BIAS.n169 CS_BIAS.n149 0.189894
R17857 CS_BIAS.n169 CS_BIAS.n168 0.189894
R17858 CS_BIAS.n168 CS_BIAS.n167 0.189894
R17859 CS_BIAS.n167 CS_BIAS.n151 0.189894
R17860 CS_BIAS.n163 CS_BIAS.n151 0.189894
R17861 CS_BIAS.n163 CS_BIAS.n162 0.189894
R17862 CS_BIAS.n162 CS_BIAS.n161 0.189894
R17863 CS_BIAS.n161 CS_BIAS.n154 0.189894
R17864 CS_BIAS.n157 CS_BIAS.n154 0.189894
R17865 CS_BIAS.n143 CS_BIAS.n111 0.189894
R17866 CS_BIAS.n139 CS_BIAS.n111 0.189894
R17867 CS_BIAS.n139 CS_BIAS.n138 0.189894
R17868 CS_BIAS.n138 CS_BIAS.n137 0.189894
R17869 CS_BIAS.n137 CS_BIAS.n113 0.189894
R17870 CS_BIAS.n133 CS_BIAS.n113 0.189894
R17871 CS_BIAS.n133 CS_BIAS.n132 0.189894
R17872 CS_BIAS.n132 CS_BIAS.n131 0.189894
R17873 CS_BIAS.n131 CS_BIAS.n115 0.189894
R17874 CS_BIAS.n127 CS_BIAS.n115 0.189894
R17875 CS_BIAS.n127 CS_BIAS.n126 0.189894
R17876 CS_BIAS.n126 CS_BIAS.n125 0.189894
R17877 CS_BIAS.n125 CS_BIAS.n118 0.189894
R17878 CS_BIAS.n121 CS_BIAS.n118 0.189894
R17879 CS_BIAS.n107 CS_BIAS.n75 0.189894
R17880 CS_BIAS.n103 CS_BIAS.n75 0.189894
R17881 CS_BIAS.n103 CS_BIAS.n102 0.189894
R17882 CS_BIAS.n102 CS_BIAS.n101 0.189894
R17883 CS_BIAS.n101 CS_BIAS.n77 0.189894
R17884 CS_BIAS.n97 CS_BIAS.n77 0.189894
R17885 CS_BIAS.n97 CS_BIAS.n96 0.189894
R17886 CS_BIAS.n96 CS_BIAS.n95 0.189894
R17887 CS_BIAS.n95 CS_BIAS.n79 0.189894
R17888 CS_BIAS.n91 CS_BIAS.n79 0.189894
R17889 CS_BIAS.n91 CS_BIAS.n90 0.189894
R17890 CS_BIAS.n90 CS_BIAS.n89 0.189894
R17891 CS_BIAS.n89 CS_BIAS.n82 0.189894
R17892 CS_BIAS.n85 CS_BIAS.n82 0.189894
R17893 CS_BIAS.n41 CS_BIAS.n9 0.189894
R17894 CS_BIAS.n37 CS_BIAS.n9 0.189894
R17895 CS_BIAS.n37 CS_BIAS.n36 0.189894
R17896 CS_BIAS.n36 CS_BIAS.n35 0.189894
R17897 CS_BIAS.n35 CS_BIAS.n11 0.189894
R17898 CS_BIAS.n31 CS_BIAS.n11 0.189894
R17899 CS_BIAS.n31 CS_BIAS.n30 0.189894
R17900 CS_BIAS.n30 CS_BIAS.n29 0.189894
R17901 CS_BIAS.n29 CS_BIAS.n13 0.189894
R17902 CS_BIAS.n25 CS_BIAS.n13 0.189894
R17903 CS_BIAS.n25 CS_BIAS.n24 0.189894
R17904 CS_BIAS.n24 CS_BIAS.n23 0.189894
R17905 CS_BIAS.n23 CS_BIAS.n16 0.189894
R17906 CS_BIAS.n19 CS_BIAS.n16 0.189894
R17907 CS_BIAS.n54 CS_BIAS.n47 0.189894
R17908 CS_BIAS.n50 CS_BIAS.n47 0.189894
R17909 CS_BIAS.n72 CS_BIAS.n1 0.189894
R17910 CS_BIAS.n68 CS_BIAS.n1 0.189894
R17911 CS_BIAS.n68 CS_BIAS.n67 0.189894
R17912 CS_BIAS.n67 CS_BIAS.n66 0.189894
R17913 CS_BIAS.n66 CS_BIAS.n3 0.189894
R17914 CS_BIAS.n62 CS_BIAS.n3 0.189894
R17915 CS_BIAS.n62 CS_BIAS.n61 0.189894
R17916 CS_BIAS.n61 CS_BIAS.n60 0.189894
R17917 CS_BIAS.n60 CS_BIAS.n5 0.189894
R17918 CS_BIAS.n56 CS_BIAS.n5 0.189894
R17919 CS_BIAS.n410 CS_BIAS.n407 0.189894
R17920 CS_BIAS.n414 CS_BIAS.n407 0.189894
R17921 CS_BIAS.n415 CS_BIAS.n414 0.189894
R17922 CS_BIAS.n416 CS_BIAS.n415 0.189894
R17923 CS_BIAS.n416 CS_BIAS.n405 0.189894
R17924 CS_BIAS.n421 CS_BIAS.n405 0.189894
R17925 CS_BIAS.n422 CS_BIAS.n421 0.189894
R17926 CS_BIAS.n423 CS_BIAS.n422 0.189894
R17927 CS_BIAS.n423 CS_BIAS.n403 0.189894
R17928 CS_BIAS.n427 CS_BIAS.n403 0.189894
R17929 CS_BIAS.n428 CS_BIAS.n427 0.189894
R17930 CS_BIAS.n429 CS_BIAS.n428 0.189894
R17931 CS_BIAS.n429 CS_BIAS.n401 0.189894
R17932 CS_BIAS.n433 CS_BIAS.n401 0.189894
R17933 CS_BIAS.n374 CS_BIAS.n371 0.189894
R17934 CS_BIAS.n378 CS_BIAS.n371 0.189894
R17935 CS_BIAS.n379 CS_BIAS.n378 0.189894
R17936 CS_BIAS.n380 CS_BIAS.n379 0.189894
R17937 CS_BIAS.n380 CS_BIAS.n369 0.189894
R17938 CS_BIAS.n385 CS_BIAS.n369 0.189894
R17939 CS_BIAS.n386 CS_BIAS.n385 0.189894
R17940 CS_BIAS.n387 CS_BIAS.n386 0.189894
R17941 CS_BIAS.n387 CS_BIAS.n367 0.189894
R17942 CS_BIAS.n391 CS_BIAS.n367 0.189894
R17943 CS_BIAS.n392 CS_BIAS.n391 0.189894
R17944 CS_BIAS.n393 CS_BIAS.n392 0.189894
R17945 CS_BIAS.n393 CS_BIAS.n365 0.189894
R17946 CS_BIAS.n397 CS_BIAS.n365 0.189894
R17947 CS_BIAS.n338 CS_BIAS.n335 0.189894
R17948 CS_BIAS.n342 CS_BIAS.n335 0.189894
R17949 CS_BIAS.n343 CS_BIAS.n342 0.189894
R17950 CS_BIAS.n344 CS_BIAS.n343 0.189894
R17951 CS_BIAS.n344 CS_BIAS.n333 0.189894
R17952 CS_BIAS.n349 CS_BIAS.n333 0.189894
R17953 CS_BIAS.n350 CS_BIAS.n349 0.189894
R17954 CS_BIAS.n351 CS_BIAS.n350 0.189894
R17955 CS_BIAS.n351 CS_BIAS.n331 0.189894
R17956 CS_BIAS.n355 CS_BIAS.n331 0.189894
R17957 CS_BIAS.n356 CS_BIAS.n355 0.189894
R17958 CS_BIAS.n357 CS_BIAS.n356 0.189894
R17959 CS_BIAS.n357 CS_BIAS.n329 0.189894
R17960 CS_BIAS.n361 CS_BIAS.n329 0.189894
R17961 CS_BIAS.n302 CS_BIAS.n299 0.189894
R17962 CS_BIAS.n306 CS_BIAS.n299 0.189894
R17963 CS_BIAS.n307 CS_BIAS.n306 0.189894
R17964 CS_BIAS.n308 CS_BIAS.n307 0.189894
R17965 CS_BIAS.n308 CS_BIAS.n297 0.189894
R17966 CS_BIAS.n313 CS_BIAS.n297 0.189894
R17967 CS_BIAS.n314 CS_BIAS.n313 0.189894
R17968 CS_BIAS.n315 CS_BIAS.n314 0.189894
R17969 CS_BIAS.n315 CS_BIAS.n295 0.189894
R17970 CS_BIAS.n319 CS_BIAS.n295 0.189894
R17971 CS_BIAS.n320 CS_BIAS.n319 0.189894
R17972 CS_BIAS.n321 CS_BIAS.n320 0.189894
R17973 CS_BIAS.n321 CS_BIAS.n293 0.189894
R17974 CS_BIAS.n325 CS_BIAS.n293 0.189894
R17975 CS_BIAS.n244 CS_BIAS.n241 0.189894
R17976 CS_BIAS.n248 CS_BIAS.n241 0.189894
R17977 CS_BIAS.n249 CS_BIAS.n248 0.189894
R17978 CS_BIAS.n250 CS_BIAS.n249 0.189894
R17979 CS_BIAS.n250 CS_BIAS.n239 0.189894
R17980 CS_BIAS.n255 CS_BIAS.n239 0.189894
R17981 CS_BIAS.n256 CS_BIAS.n255 0.189894
R17982 CS_BIAS.n257 CS_BIAS.n256 0.189894
R17983 CS_BIAS.n257 CS_BIAS.n237 0.189894
R17984 CS_BIAS.n261 CS_BIAS.n237 0.189894
R17985 CS_BIAS.n262 CS_BIAS.n261 0.189894
R17986 CS_BIAS.n263 CS_BIAS.n262 0.189894
R17987 CS_BIAS.n263 CS_BIAS.n235 0.189894
R17988 CS_BIAS.n267 CS_BIAS.n235 0.189894
R17989 CS_BIAS.n228 CS_BIAS.n225 0.189894
R17990 CS_BIAS.n232 CS_BIAS.n225 0.189894
R17991 CS_BIAS.n273 CS_BIAS.n223 0.189894
R17992 CS_BIAS.n278 CS_BIAS.n223 0.189894
R17993 CS_BIAS.n279 CS_BIAS.n278 0.189894
R17994 CS_BIAS.n280 CS_BIAS.n279 0.189894
R17995 CS_BIAS.n280 CS_BIAS.n221 0.189894
R17996 CS_BIAS.n284 CS_BIAS.n221 0.189894
R17997 CS_BIAS.n285 CS_BIAS.n284 0.189894
R17998 CS_BIAS.n286 CS_BIAS.n285 0.189894
R17999 CS_BIAS.n286 CS_BIAS.n219 0.189894
R18000 CS_BIAS.n290 CS_BIAS.n219 0.189894
R18001 CS_BIAS.n55 CS_BIAS.n54 0.170955
R18002 CS_BIAS.n56 CS_BIAS.n55 0.170955
R18003 CS_BIAS.n272 CS_BIAS.n232 0.170955
R18004 CS_BIAS.n273 CS_BIAS.n272 0.170955
R18005 VOUT.n9 VOUT.t41 119.948
R18006 VOUT.n0 VOUT.t44 118.448
R18007 VOUT.n9 VOUT.t43 116.844
R18008 VOUT.n10 VOUT.t40 116.844
R18009 VOUT.n1 VOUT.t42 115.344
R18010 VOUT.n0 VOUT.t45 115.344
R18011 VOUT.n29 VOUT.n27 88.2696
R18012 VOUT.n25 VOUT.n23 88.2696
R18013 VOUT.n21 VOUT.n19 88.2696
R18014 VOUT.n17 VOUT.n15 88.2696
R18015 VOUT.n14 VOUT.n12 88.2696
R18016 VOUT.n49 VOUT.n47 88.2696
R18017 VOUT.n45 VOUT.n43 88.2696
R18018 VOUT.n41 VOUT.n39 88.2696
R18019 VOUT.n37 VOUT.n35 88.2696
R18020 VOUT.n34 VOUT.n32 88.2696
R18021 VOUT.n29 VOUT.n28 84.9593
R18022 VOUT.n25 VOUT.n24 84.9593
R18023 VOUT.n21 VOUT.n20 84.9593
R18024 VOUT.n17 VOUT.n16 84.9593
R18025 VOUT.n14 VOUT.n13 84.9593
R18026 VOUT.n49 VOUT.n48 84.9593
R18027 VOUT.n45 VOUT.n44 84.9593
R18028 VOUT.n41 VOUT.n40 84.9593
R18029 VOUT.n37 VOUT.n36 84.9593
R18030 VOUT.n34 VOUT.n33 84.9593
R18031 VOUT.n18 VOUT.n14 9.00697
R18032 VOUT.n38 VOUT.n34 9.00697
R18033 VOUT.n31 VOUT.n11 8.54861
R18034 VOUT.n28 VOUT.t23 8.2505
R18035 VOUT.n28 VOUT.t35 8.2505
R18036 VOUT.n27 VOUT.t4 8.2505
R18037 VOUT.n27 VOUT.t27 8.2505
R18038 VOUT.n24 VOUT.t31 8.2505
R18039 VOUT.n24 VOUT.t0 8.2505
R18040 VOUT.n23 VOUT.t10 8.2505
R18041 VOUT.n23 VOUT.t33 8.2505
R18042 VOUT.n20 VOUT.t6 8.2505
R18043 VOUT.n20 VOUT.t16 8.2505
R18044 VOUT.n19 VOUT.t29 8.2505
R18045 VOUT.n19 VOUT.t28 8.2505
R18046 VOUT.n16 VOUT.t13 8.2505
R18047 VOUT.n16 VOUT.t20 8.2505
R18048 VOUT.n15 VOUT.t34 8.2505
R18049 VOUT.n15 VOUT.t17 8.2505
R18050 VOUT.n13 VOUT.t7 8.2505
R18051 VOUT.n13 VOUT.t11 8.2505
R18052 VOUT.n12 VOUT.t39 8.2505
R18053 VOUT.n12 VOUT.t14 8.2505
R18054 VOUT.n47 VOUT.t30 8.2505
R18055 VOUT.n47 VOUT.t21 8.2505
R18056 VOUT.n48 VOUT.t9 8.2505
R18057 VOUT.n48 VOUT.t1 8.2505
R18058 VOUT.n43 VOUT.t36 8.2505
R18059 VOUT.n43 VOUT.t24 8.2505
R18060 VOUT.n44 VOUT.t15 8.2505
R18061 VOUT.n44 VOUT.t3 8.2505
R18062 VOUT.n39 VOUT.t26 8.2505
R18063 VOUT.n39 VOUT.t19 8.2505
R18064 VOUT.n40 VOUT.t5 8.2505
R18065 VOUT.n40 VOUT.t38 8.2505
R18066 VOUT.n35 VOUT.t18 8.2505
R18067 VOUT.n35 VOUT.t8 8.2505
R18068 VOUT.n36 VOUT.t37 8.2505
R18069 VOUT.n36 VOUT.t25 8.2505
R18070 VOUT.n32 VOUT.t22 8.2505
R18071 VOUT.n32 VOUT.t2 8.2505
R18072 VOUT.n33 VOUT.t32 8.2505
R18073 VOUT.n33 VOUT.t12 8.2505
R18074 VOUT.n30 VOUT.n29 7.05653
R18075 VOUT.n26 VOUT.n25 7.05653
R18076 VOUT.n22 VOUT.n21 7.05653
R18077 VOUT.n18 VOUT.n17 7.05653
R18078 VOUT.n50 VOUT.n49 7.05653
R18079 VOUT.n46 VOUT.n45 7.05653
R18080 VOUT.n42 VOUT.n41 7.05653
R18081 VOUT.n38 VOUT.n37 7.05653
R18082 VOUT.n11 VOUT.n10 6.00964
R18083 VOUT.n2 VOUT.n1 6.00964
R18084 VOUT.n31 VOUT.n30 5.8049
R18085 VOUT.n51 VOUT.n50 5.8049
R18086 VOUT.n52 VOUT.n2 4.59255
R18087 VOUT.n8 VOUT 4.4044
R18088 VOUT.n11 VOUT.n2 3.98171
R18089 VOUT.n52 VOUT.n51 3.93706
R18090 VOUT.n51 VOUT.n31 3.38356
R18091 VOUT.n10 VOUT.n9 3.1061
R18092 VOUT.n1 VOUT.n0 3.1061
R18093 VOUT.n22 VOUT.n18 1.95093
R18094 VOUT.n26 VOUT.n22 1.95093
R18095 VOUT.n30 VOUT.n26 1.95093
R18096 VOUT.n42 VOUT.n38 1.95093
R18097 VOUT.n46 VOUT.n42 1.95093
R18098 VOUT.n50 VOUT.n46 1.95093
R18099 VOUT.n52 VOUT.n8 0.43149
R18100 VOUT.n8 VOUT.n7 0.400809
R18101 VOUT.n6 VOUT.n5 0.115454
R18102 VOUT.n4 VOUT.n3 0.112341
R18103 VOUT.n5 VOUT.n4 0.0612264
R18104 VOUT.n7 VOUT.n3 0.0544562
R18105 VOUT.n3 VOUT.t49 0.019303
R18106 VOUT.n4 VOUT.t47 0.0184469
R18107 VOUT.n5 VOUT.t48 0.0184262
R18108 VOUT.n6 VOUT.t46 0.0168887
R18109 VOUT.n7 VOUT.n6 0.0123828
R18110 VOUT VOUT.n52 0.0099
R18111 a_n1578_n2628.n73 a_n1578_n2628.n69 289.615
R18112 a_n1578_n2628.n61 a_n1578_n2628.n11 215.245
R18113 a_n1578_n2628.n57 a_n1578_n2628.n13 215.245
R18114 a_n1578_n2628.n53 a_n1578_n2628.n15 215.245
R18115 a_n1578_n2628.n1 a_n1578_n2628.n0 11.0009
R18116 a_n1578_n2628.n3 a_n1578_n2628.n2 11.0009
R18117 a_n1578_n2628.n5 a_n1578_n2628.n4 11.6603
R18118 a_n1578_n2628.n74 a_n1578_n2628.n73 185
R18119 a_n1578_n2628.n72 a_n1578_n2628.n71 185
R18120 a_n1578_n2628.n10 a_n1578_n2628.n11 7.50266
R18121 a_n1578_n2628.n61 a_n1578_n2628.n29 185
R18122 a_n1578_n2628.n35 a_n1578_n2628.n34 185
R18123 a_n1578_n2628.n43 a_n1578_n2628.n60 185
R18124 a_n1578_n2628.n59 a_n1578_n2628.n46 185
R18125 a_n1578_n2628.n12 a_n1578_n2628.n13 7.50266
R18126 a_n1578_n2628.n57 a_n1578_n2628.n31 185
R18127 a_n1578_n2628.n38 a_n1578_n2628.n37 185
R18128 a_n1578_n2628.n44 a_n1578_n2628.n56 185
R18129 a_n1578_n2628.n55 a_n1578_n2628.n47 185
R18130 a_n1578_n2628.n14 a_n1578_n2628.n15 7.50266
R18131 a_n1578_n2628.n53 a_n1578_n2628.n33 185
R18132 a_n1578_n2628.n41 a_n1578_n2628.n40 185
R18133 a_n1578_n2628.n45 a_n1578_n2628.n52 185
R18134 a_n1578_n2628.n51 a_n1578_n2628.n48 185
R18135 a_n1578_n2628.n68 a_n1578_n2628.n67 185
R18136 a_n1578_n2628.n65 a_n1578_n2628.n64 185
R18137 a_n1578_n2628.n78 a_n1578_n2628.n77 185
R18138 a_n1578_n2628.n22 a_n1578_n2628.t6 150.499
R18139 a_n1578_n2628.n25 a_n1578_n2628.t0 150.499
R18140 a_n1578_n2628.t5 a_n1578_n2628.n26 150.499
R18141 a_n1578_n2628.n19 a_n1578_n2628.t4 150.499
R18142 a_n1578_n2628.n28 a_n1578_n2628.t2 150.026
R18143 a_n1578_n2628.n30 a_n1578_n2628.t1 150.026
R18144 a_n1578_n2628.n32 a_n1578_n2628.t3 150.026
R18145 a_n1578_n2628.n6 a_n1578_n2628.n54 140.091
R18146 a_n1578_n2628.n9 a_n1578_n2628.n62 138.31
R18147 a_n1578_n2628.n6 a_n1578_n2628.n58 138.31
R18148 a_n1578_n2628.n73 a_n1578_n2628.n72 104.615
R18149 a_n1578_n2628.n72 a_n1578_n2628.n17 104.615
R18150 a_n1578_n2628.n61 a_n1578_n2628.n34 104.615
R18151 a_n1578_n2628.n60 a_n1578_n2628.n34 104.615
R18152 a_n1578_n2628.n60 a_n1578_n2628.n59 104.615
R18153 a_n1578_n2628.n57 a_n1578_n2628.n37 104.615
R18154 a_n1578_n2628.n56 a_n1578_n2628.n37 104.615
R18155 a_n1578_n2628.n56 a_n1578_n2628.n55 104.615
R18156 a_n1578_n2628.n53 a_n1578_n2628.n40 104.615
R18157 a_n1578_n2628.n52 a_n1578_n2628.n40 104.615
R18158 a_n1578_n2628.n52 a_n1578_n2628.n51 104.615
R18159 a_n1578_n2628.n68 a_n1578_n2628.n20 104.615
R18160 a_n1578_n2628.n1 a_n1578_n2628.n68 214.453
R18161 a_n1578_n2628.n65 a_n1578_n2628.n23 104.615
R18162 a_n1578_n2628.n3 a_n1578_n2628.n65 214.453
R18163 a_n1578_n2628.n77 a_n1578_n2628.n5 214.453
R18164 a_n1578_n2628.n77 a_n1578_n2628.n50 104.615
R18165 a_n1578_n2628.t4 a_n1578_n2628.n17 52.3082
R18166 a_n1578_n2628.n59 a_n1578_n2628.t2 52.3082
R18167 a_n1578_n2628.n55 a_n1578_n2628.t1 52.3082
R18168 a_n1578_n2628.n51 a_n1578_n2628.t3 52.3082
R18169 a_n1578_n2628.t6 a_n1578_n2628.n20 52.3082
R18170 a_n1578_n2628.t0 a_n1578_n2628.n23 52.3082
R18171 a_n1578_n2628.t5 a_n1578_n2628.n50 52.3082
R18172 a_n1578_n2628.n16 a_n1578_n2628.n76 29.8581
R18173 a_n1578_n2628.n8 a_n1578_n2628.n0 33.0811
R18174 a_n1578_n2628.n8 a_n1578_n2628.n2 33.0811
R18175 a_n1578_n2628.n4 a_n1578_n2628.n16 32.7555
R18176 a_n1578_n2628.n46 a_n1578_n2628.n28 5.10304
R18177 a_n1578_n2628.n47 a_n1578_n2628.n30 5.10304
R18178 a_n1578_n2628.n48 a_n1578_n2628.n32 5.10304
R18179 a_n1578_n2628.n7 a_n1578_n2628.n6 4.23592
R18180 a_n1578_n2628.n43 a_n1578_n2628.n46 12.8005
R18181 a_n1578_n2628.n44 a_n1578_n2628.n47 12.8005
R18182 a_n1578_n2628.n45 a_n1578_n2628.n48 12.8005
R18183 a_n1578_n2628.n4 a_n1578_n2628.n26 3.73448
R18184 a_n1578_n2628.n33 a_n1578_n2628.n14 3.56777
R18185 a_n1578_n2628.n31 a_n1578_n2628.n12 3.56777
R18186 a_n1578_n2628.n29 a_n1578_n2628.n10 3.56777
R18187 a_n1578_n2628.n36 a_n1578_n2628.n35 4.008
R18188 a_n1578_n2628.n39 a_n1578_n2628.n38 4.008
R18189 a_n1578_n2628.n42 a_n1578_n2628.n41 4.008
R18190 a_n1578_n2628.n29 a_n1578_n2628.n35 11.249
R18191 a_n1578_n2628.n31 a_n1578_n2628.n38 11.249
R18192 a_n1578_n2628.n33 a_n1578_n2628.n41 11.249
R18193 a_n1578_n2628.n8 a_n1578_n2628.n6 10.7289
R18194 a_n1578_n2628.n42 a_n1578_n2628.n45 3.73143
R18195 a_n1578_n2628.n39 a_n1578_n2628.n44 3.73143
R18196 a_n1578_n2628.n36 a_n1578_n2628.n43 3.73143
R18197 a_n1578_n2628.n19 a_n1578_n2628.n18 3.53826
R18198 a_n1578_n2628.n22 a_n1578_n2628.n21 3.53826
R18199 a_n1578_n2628.n25 a_n1578_n2628.n24 3.53826
R18200 a_n1578_n2628.n26 a_n1578_n2628.n27 3.53826
R18201 a_n1578_n2628.n76 a_n1578_n2628.n69 9.69747
R18202 a_n1578_n2628.n76 a_n1578_n2628.n19 9.45567
R18203 a_n1578_n2628.n62 a_n1578_n2628.n28 9.45567
R18204 a_n1578_n2628.n58 a_n1578_n2628.n30 9.45567
R18205 a_n1578_n2628.n54 a_n1578_n2628.n32 9.45567
R18206 a_n1578_n2628.n70 a_n1578_n2628.n19 9.3005
R18207 a_n1578_n2628.n22 a_n1578_n2628.n0 3.09156
R18208 a_n1578_n2628.n25 a_n1578_n2628.n2 3.09156
R18209 a_n1578_n2628.n26 a_n1578_n2628.n49 9.3005
R18210 a_n1578_n2628.n75 a_n1578_n2628.n74 8.92171
R18211 a_n1578_n2628.n71 a_n1578_n2628.n70 8.14595
R18212 a_n1578_n2628.n67 a_n1578_n2628.n66 8.14595
R18213 a_n1578_n2628.n64 a_n1578_n2628.n63 8.14595
R18214 a_n1578_n2628.n78 a_n1578_n2628.n49 8.14595
R18215 a_n1578_n2628.n18 a_n1578_n2628.n17 187.804
R18216 a_n1578_n2628.n21 a_n1578_n2628.n20 187.804
R18217 a_n1578_n2628.n24 a_n1578_n2628.n23 187.804
R18218 a_n1578_n2628.n50 a_n1578_n2628.n27 187.804
R18219 a_n1578_n2628.n49 a_n1578_n2628.n5 10.0449
R18220 a_n1578_n2628.n16 a_n1578_n2628.n7 5.43859
R18221 a_n1578_n2628.n28 a_n1578_n2628.n10 4.35729
R18222 a_n1578_n2628.n30 a_n1578_n2628.n12 4.35729
R18223 a_n1578_n2628.n32 a_n1578_n2628.n14 4.35729
R18224 a_n1578_n2628.n63 a_n1578_n2628.n25 12.4975
R18225 a_n1578_n2628.n66 a_n1578_n2628.n22 12.4975
R18226 a_n1578_n2628.n19 a_n1578_n2628.n75 12.4975
R18227 a_n1578_n2628.n9 a_n1578_n2628.n7 4.36906
R18228 a_n1578_n2628.n9 a_n1578_n2628.n8 11.1988
R18229 a_n1578_n2628.n71 a_n1578_n2628.n18 8.3669
R18230 a_n1578_n2628.n67 a_n1578_n2628.n21 8.3669
R18231 a_n1578_n2628.n64 a_n1578_n2628.n24 8.3669
R18232 a_n1578_n2628.n27 a_n1578_n2628.n78 8.3669
R18233 a_n1578_n2628.n36 a_n1578_n2628.n28 5.53918
R18234 a_n1578_n2628.n39 a_n1578_n2628.n30 5.53918
R18235 a_n1578_n2628.n42 a_n1578_n2628.n32 5.53918
R18236 a_n1578_n2628.n74 a_n1578_n2628.n70 5.04292
R18237 a_n1578_n2628.n1 a_n1578_n2628.n66 10.0449
R18238 a_n1578_n2628.n3 a_n1578_n2628.n63 10.0449
R18239 a_n1578_n2628.n75 a_n1578_n2628.n69 4.26717
R18240 a_n1578_n2628.n62 a_n1578_n2628.n11 10.0664
R18241 a_n1578_n2628.n58 a_n1578_n2628.n13 10.0664
R18242 a_n1578_n2628.n54 a_n1578_n2628.n15 10.0664
R18243 a_n12120_6849.n25 a_n12120_6849.n17 289.615
R18244 a_n12120_6849.n13 a_n12120_6849.n5 289.615
R18245 a_n12120_6849.n20 a_n12120_6849.n19 185
R18246 a_n12120_6849.n24 a_n12120_6849.n23 185
R18247 a_n12120_6849.n26 a_n12120_6849.n25 185
R18248 a_n12120_6849.n14 a_n12120_6849.n13 185
R18249 a_n12120_6849.n12 a_n12120_6849.n11 185
R18250 a_n12120_6849.n8 a_n12120_6849.n7 185
R18251 a_n12120_6849.n21 a_n12120_6849.t0 150.499
R18252 a_n12120_6849.n9 a_n12120_6849.t1 150.499
R18253 a_n12120_6849.n4 a_n12120_6849.n2 142.626
R18254 a_n12120_6849.n38 a_n12120_6849.n37 142.626
R18255 a_n12120_6849.n4 a_n12120_6849.n3 138.653
R18256 a_n12120_6849.n39 a_n12120_6849.n38 138.651
R18257 a_n12120_6849.n24 a_n12120_6849.n19 104.615
R18258 a_n12120_6849.n25 a_n12120_6849.n24 104.615
R18259 a_n12120_6849.n13 a_n12120_6849.n12 104.615
R18260 a_n12120_6849.n12 a_n12120_6849.n7 104.615
R18261 a_n12120_6849.n30 a_n12120_6849.t15 85.8441
R18262 a_n12120_6849.n32 a_n12120_6849.t14 85.8429
R18263 a_n12120_6849.n29 a_n12120_6849.n28 85.2565
R18264 a_n12120_6849.n31 a_n12120_6849.t13 83.0998
R18265 a_n12120_6849.n30 a_n12120_6849.t12 83.0998
R18266 a_n12120_6849.n33 a_n12120_6849.t10 83.0986
R18267 a_n12120_6849.n32 a_n12120_6849.t11 83.0986
R18268 a_n12120_6849.t0 a_n12120_6849.n19 52.3082
R18269 a_n12120_6849.t1 a_n12120_6849.n7 52.3082
R18270 a_n12120_6849.n38 a_n12120_6849.n36 50.7956
R18271 a_n12120_6849.n29 a_n12120_6849.n16 47.8638
R18272 a_n12120_6849.n36 a_n12120_6849.n4 42.6536
R18273 a_n12120_6849.n35 a_n12120_6849.n29 12.3668
R18274 a_n12120_6849.n37 a_n12120_6849.t8 11.651
R18275 a_n12120_6849.n37 a_n12120_6849.t7 11.651
R18276 a_n12120_6849.n3 a_n12120_6849.t3 11.651
R18277 a_n12120_6849.n3 a_n12120_6849.t2 11.651
R18278 a_n12120_6849.n2 a_n12120_6849.t5 11.651
R18279 a_n12120_6849.n2 a_n12120_6849.t4 11.651
R18280 a_n12120_6849.n39 a_n12120_6849.t6 11.651
R18281 a_n12120_6849.t9 a_n12120_6849.n39 11.651
R18282 a_n12120_6849.n36 a_n12120_6849.n35 11.5607
R18283 a_n12120_6849.n21 a_n12120_6849.n20 10.2326
R18284 a_n12120_6849.n9 a_n12120_6849.n8 10.2326
R18285 a_n12120_6849.n28 a_n12120_6849.n17 9.69747
R18286 a_n12120_6849.n16 a_n12120_6849.n5 9.69747
R18287 a_n12120_6849.n28 a_n12120_6849.n1 9.45567
R18288 a_n12120_6849.n16 a_n12120_6849.n0 9.45567
R18289 a_n12120_6849.n22 a_n12120_6849.n1 9.3005
R18290 a_n12120_6849.n18 a_n12120_6849.n1 9.3005
R18291 a_n12120_6849.n1 a_n12120_6849.n27 9.3005
R18292 a_n12120_6849.n6 a_n12120_6849.n0 9.3005
R18293 a_n12120_6849.n0 a_n12120_6849.n15 9.3005
R18294 a_n12120_6849.n10 a_n12120_6849.n0 9.3005
R18295 a_n12120_6849.n27 a_n12120_6849.n26 8.92171
R18296 a_n12120_6849.n15 a_n12120_6849.n14 8.92171
R18297 a_n12120_6849.n23 a_n12120_6849.n18 8.14595
R18298 a_n12120_6849.n11 a_n12120_6849.n6 8.14595
R18299 a_n12120_6849.n22 a_n12120_6849.n20 7.3702
R18300 a_n12120_6849.n10 a_n12120_6849.n8 7.3702
R18301 a_n12120_6849.n34 a_n12120_6849.n31 6.44791
R18302 a_n12120_6849.n34 a_n12120_6849.n33 6.2151
R18303 a_n12120_6849.n23 a_n12120_6849.n22 5.81868
R18304 a_n12120_6849.n11 a_n12120_6849.n10 5.81868
R18305 a_n12120_6849.n26 a_n12120_6849.n18 5.04292
R18306 a_n12120_6849.n14 a_n12120_6849.n6 5.04292
R18307 a_n12120_6849.n27 a_n12120_6849.n17 4.26717
R18308 a_n12120_6849.n15 a_n12120_6849.n5 4.26717
R18309 a_n12120_6849.n35 a_n12120_6849.n34 3.4105
R18310 a_n12120_6849.n1 a_n12120_6849.n21 3.19753
R18311 a_n12120_6849.n0 a_n12120_6849.n9 3.19753
R18312 a_n12120_6849.n33 a_n12120_6849.n32 2.74482
R18313 a_n12120_6849.n31 a_n12120_6849.n30 2.74482
R18314 VN.n1 VN.t0 243.97
R18315 VN.n1 VN.t1 243.255
R18316 VN.n0 VN.t2 78.9867
R18317 VN.n0 VN.t3 58.2236
R18318 VN VN.n2 15.5475
R18319 VN.n2 VN.n1 5.04791
R18320 VN.n2 VN.n0 1.188
R18321 DIFFPAIR_BIAS.n18 DIFFPAIR_BIAS.n0 289.615
R18322 DIFFPAIR_BIAS.n41 DIFFPAIR_BIAS.n23 289.615
R18323 DIFFPAIR_BIAS.n65 DIFFPAIR_BIAS.n47 289.615
R18324 DIFFPAIR_BIAS.n19 DIFFPAIR_BIAS.n18 185
R18325 DIFFPAIR_BIAS.n17 DIFFPAIR_BIAS.n16 185
R18326 DIFFPAIR_BIAS.n4 DIFFPAIR_BIAS.n3 185
R18327 DIFFPAIR_BIAS.n11 DIFFPAIR_BIAS.n10 185
R18328 DIFFPAIR_BIAS.n9 DIFFPAIR_BIAS.n8 185
R18329 DIFFPAIR_BIAS.n42 DIFFPAIR_BIAS.n41 185
R18330 DIFFPAIR_BIAS.n40 DIFFPAIR_BIAS.n39 185
R18331 DIFFPAIR_BIAS.n27 DIFFPAIR_BIAS.n26 185
R18332 DIFFPAIR_BIAS.n34 DIFFPAIR_BIAS.n33 185
R18333 DIFFPAIR_BIAS.n32 DIFFPAIR_BIAS.n31 185
R18334 DIFFPAIR_BIAS.n66 DIFFPAIR_BIAS.n65 185
R18335 DIFFPAIR_BIAS.n64 DIFFPAIR_BIAS.n63 185
R18336 DIFFPAIR_BIAS.n51 DIFFPAIR_BIAS.n50 185
R18337 DIFFPAIR_BIAS.n58 DIFFPAIR_BIAS.n57 185
R18338 DIFFPAIR_BIAS.n56 DIFFPAIR_BIAS.n55 185
R18339 DIFFPAIR_BIAS.n7 DIFFPAIR_BIAS.t1 147.714
R18340 DIFFPAIR_BIAS.n30 DIFFPAIR_BIAS.t5 147.714
R18341 DIFFPAIR_BIAS.n54 DIFFPAIR_BIAS.t3 147.714
R18342 DIFFPAIR_BIAS.n18 DIFFPAIR_BIAS.n17 104.615
R18343 DIFFPAIR_BIAS.n17 DIFFPAIR_BIAS.n3 104.615
R18344 DIFFPAIR_BIAS.n10 DIFFPAIR_BIAS.n3 104.615
R18345 DIFFPAIR_BIAS.n10 DIFFPAIR_BIAS.n9 104.615
R18346 DIFFPAIR_BIAS.n41 DIFFPAIR_BIAS.n40 104.615
R18347 DIFFPAIR_BIAS.n40 DIFFPAIR_BIAS.n26 104.615
R18348 DIFFPAIR_BIAS.n33 DIFFPAIR_BIAS.n26 104.615
R18349 DIFFPAIR_BIAS.n33 DIFFPAIR_BIAS.n32 104.615
R18350 DIFFPAIR_BIAS.n65 DIFFPAIR_BIAS.n64 104.615
R18351 DIFFPAIR_BIAS.n64 DIFFPAIR_BIAS.n50 104.615
R18352 DIFFPAIR_BIAS.n57 DIFFPAIR_BIAS.n50 104.615
R18353 DIFFPAIR_BIAS.n57 DIFFPAIR_BIAS.n56 104.615
R18354 DIFFPAIR_BIAS.n46 DIFFPAIR_BIAS.n22 74.2464
R18355 DIFFPAIR_BIAS.n46 DIFFPAIR_BIAS.n45 70.0429
R18356 DIFFPAIR_BIAS.n70 DIFFPAIR_BIAS.n69 70.0429
R18357 DIFFPAIR_BIAS.n9 DIFFPAIR_BIAS.t1 52.3082
R18358 DIFFPAIR_BIAS.n32 DIFFPAIR_BIAS.t5 52.3082
R18359 DIFFPAIR_BIAS.n56 DIFFPAIR_BIAS.t3 52.3082
R18360 DIFFPAIR_BIAS.n71 DIFFPAIR_BIAS.t0 50.1011
R18361 DIFFPAIR_BIAS.n76 DIFFPAIR_BIAS.t7 48.1263
R18362 DIFFPAIR_BIAS.n71 DIFFPAIR_BIAS.t4 45.8969
R18363 DIFFPAIR_BIAS.n72 DIFFPAIR_BIAS.t2 45.8969
R18364 DIFFPAIR_BIAS.n75 DIFFPAIR_BIAS.t8 45.1196
R18365 DIFFPAIR_BIAS.n74 DIFFPAIR_BIAS.t6 45.1196
R18366 DIFFPAIR_BIAS.n8 DIFFPAIR_BIAS.n7 15.6631
R18367 DIFFPAIR_BIAS.n31 DIFFPAIR_BIAS.n30 15.6631
R18368 DIFFPAIR_BIAS.n55 DIFFPAIR_BIAS.n54 15.6631
R18369 DIFFPAIR_BIAS.n11 DIFFPAIR_BIAS.n6 12.8005
R18370 DIFFPAIR_BIAS.n34 DIFFPAIR_BIAS.n29 12.8005
R18371 DIFFPAIR_BIAS.n58 DIFFPAIR_BIAS.n53 12.8005
R18372 DIFFPAIR_BIAS.n12 DIFFPAIR_BIAS.n4 12.0247
R18373 DIFFPAIR_BIAS.n35 DIFFPAIR_BIAS.n27 12.0247
R18374 DIFFPAIR_BIAS.n59 DIFFPAIR_BIAS.n51 12.0247
R18375 DIFFPAIR_BIAS.n16 DIFFPAIR_BIAS.n15 11.249
R18376 DIFFPAIR_BIAS.n39 DIFFPAIR_BIAS.n38 11.249
R18377 DIFFPAIR_BIAS.n63 DIFFPAIR_BIAS.n62 11.249
R18378 DIFFPAIR_BIAS.n19 DIFFPAIR_BIAS.n2 10.4732
R18379 DIFFPAIR_BIAS.n42 DIFFPAIR_BIAS.n25 10.4732
R18380 DIFFPAIR_BIAS.n66 DIFFPAIR_BIAS.n49 10.4732
R18381 DIFFPAIR_BIAS.n20 DIFFPAIR_BIAS.n0 9.69747
R18382 DIFFPAIR_BIAS.n43 DIFFPAIR_BIAS.n23 9.69747
R18383 DIFFPAIR_BIAS.n67 DIFFPAIR_BIAS.n47 9.69747
R18384 DIFFPAIR_BIAS.n22 DIFFPAIR_BIAS.n21 9.45567
R18385 DIFFPAIR_BIAS.n45 DIFFPAIR_BIAS.n44 9.45567
R18386 DIFFPAIR_BIAS.n69 DIFFPAIR_BIAS.n68 9.45567
R18387 DIFFPAIR_BIAS.n21 DIFFPAIR_BIAS.n20 9.3005
R18388 DIFFPAIR_BIAS.n2 DIFFPAIR_BIAS.n1 9.3005
R18389 DIFFPAIR_BIAS.n15 DIFFPAIR_BIAS.n14 9.3005
R18390 DIFFPAIR_BIAS.n13 DIFFPAIR_BIAS.n12 9.3005
R18391 DIFFPAIR_BIAS.n6 DIFFPAIR_BIAS.n5 9.3005
R18392 DIFFPAIR_BIAS.n44 DIFFPAIR_BIAS.n43 9.3005
R18393 DIFFPAIR_BIAS.n25 DIFFPAIR_BIAS.n24 9.3005
R18394 DIFFPAIR_BIAS.n38 DIFFPAIR_BIAS.n37 9.3005
R18395 DIFFPAIR_BIAS.n36 DIFFPAIR_BIAS.n35 9.3005
R18396 DIFFPAIR_BIAS.n29 DIFFPAIR_BIAS.n28 9.3005
R18397 DIFFPAIR_BIAS.n68 DIFFPAIR_BIAS.n67 9.3005
R18398 DIFFPAIR_BIAS.n49 DIFFPAIR_BIAS.n48 9.3005
R18399 DIFFPAIR_BIAS.n62 DIFFPAIR_BIAS.n61 9.3005
R18400 DIFFPAIR_BIAS.n60 DIFFPAIR_BIAS.n59 9.3005
R18401 DIFFPAIR_BIAS.n53 DIFFPAIR_BIAS.n52 9.3005
R18402 DIFFPAIR_BIAS.n73 DIFFPAIR_BIAS.n72 6.91702
R18403 DIFFPAIR_BIAS.n73 DIFFPAIR_BIAS.n70 6.21567
R18404 DIFFPAIR_BIAS.n74 DIFFPAIR_BIAS.n73 4.85213
R18405 DIFFPAIR_BIAS.n7 DIFFPAIR_BIAS.n5 4.39059
R18406 DIFFPAIR_BIAS.n30 DIFFPAIR_BIAS.n28 4.39059
R18407 DIFFPAIR_BIAS.n54 DIFFPAIR_BIAS.n52 4.39059
R18408 DIFFPAIR_BIAS.n22 DIFFPAIR_BIAS.n0 4.26717
R18409 DIFFPAIR_BIAS.n45 DIFFPAIR_BIAS.n23 4.26717
R18410 DIFFPAIR_BIAS.n69 DIFFPAIR_BIAS.n47 4.26717
R18411 DIFFPAIR_BIAS.n72 DIFFPAIR_BIAS.n71 4.20583
R18412 DIFFPAIR_BIAS.n75 DIFFPAIR_BIAS.n74 4.20559
R18413 DIFFPAIR_BIAS.n70 DIFFPAIR_BIAS.n46 4.20399
R18414 DIFFPAIR_BIAS.n20 DIFFPAIR_BIAS.n19 3.49141
R18415 DIFFPAIR_BIAS.n43 DIFFPAIR_BIAS.n42 3.49141
R18416 DIFFPAIR_BIAS.n67 DIFFPAIR_BIAS.n66 3.49141
R18417 DIFFPAIR_BIAS.n16 DIFFPAIR_BIAS.n2 2.71565
R18418 DIFFPAIR_BIAS.n39 DIFFPAIR_BIAS.n25 2.71565
R18419 DIFFPAIR_BIAS.n63 DIFFPAIR_BIAS.n49 2.71565
R18420 DIFFPAIR_BIAS.n15 DIFFPAIR_BIAS.n4 1.93989
R18421 DIFFPAIR_BIAS.n38 DIFFPAIR_BIAS.n27 1.93989
R18422 DIFFPAIR_BIAS.n62 DIFFPAIR_BIAS.n51 1.93989
R18423 DIFFPAIR_BIAS.n12 DIFFPAIR_BIAS.n11 1.16414
R18424 DIFFPAIR_BIAS.n35 DIFFPAIR_BIAS.n34 1.16414
R18425 DIFFPAIR_BIAS.n59 DIFFPAIR_BIAS.n58 1.16414
R18426 DIFFPAIR_BIAS.n76 DIFFPAIR_BIAS.n75 0.907034
R18427 DIFFPAIR_BIAS DIFFPAIR_BIAS.n76 0.683625
R18428 DIFFPAIR_BIAS.n8 DIFFPAIR_BIAS.n6 0.388379
R18429 DIFFPAIR_BIAS.n31 DIFFPAIR_BIAS.n29 0.388379
R18430 DIFFPAIR_BIAS.n55 DIFFPAIR_BIAS.n53 0.388379
R18431 DIFFPAIR_BIAS.n21 DIFFPAIR_BIAS.n1 0.155672
R18432 DIFFPAIR_BIAS.n14 DIFFPAIR_BIAS.n1 0.155672
R18433 DIFFPAIR_BIAS.n14 DIFFPAIR_BIAS.n13 0.155672
R18434 DIFFPAIR_BIAS.n13 DIFFPAIR_BIAS.n5 0.155672
R18435 DIFFPAIR_BIAS.n44 DIFFPAIR_BIAS.n24 0.155672
R18436 DIFFPAIR_BIAS.n37 DIFFPAIR_BIAS.n24 0.155672
R18437 DIFFPAIR_BIAS.n37 DIFFPAIR_BIAS.n36 0.155672
R18438 DIFFPAIR_BIAS.n36 DIFFPAIR_BIAS.n28 0.155672
R18439 DIFFPAIR_BIAS.n68 DIFFPAIR_BIAS.n48 0.155672
R18440 DIFFPAIR_BIAS.n61 DIFFPAIR_BIAS.n48 0.155672
R18441 DIFFPAIR_BIAS.n61 DIFFPAIR_BIAS.n60 0.155672
R18442 DIFFPAIR_BIAS.n60 DIFFPAIR_BIAS.n52 0.155672
R18443 a_n2838_n2628.n34 a_n2838_n2628.n1 215.245
R18444 a_n2838_n2628.n30 a_n2838_n2628.n3 215.245
R18445 a_n2838_n2628.n10 a_n2838_n2628.n5 215.245
R18446 a_n2838_n2628.n0 a_n2838_n2628.n1 7.50266
R18447 a_n2838_n2628.n34 a_n2838_n2628.n7 185
R18448 a_n2838_n2628.n14 a_n2838_n2628.n13 185
R18449 a_n2838_n2628.n21 a_n2838_n2628.n33 185
R18450 a_n2838_n2628.n32 a_n2838_n2628.n24 185
R18451 a_n2838_n2628.n2 a_n2838_n2628.n3 7.50266
R18452 a_n2838_n2628.n30 a_n2838_n2628.n9 185
R18453 a_n2838_n2628.n17 a_n2838_n2628.n16 185
R18454 a_n2838_n2628.n22 a_n2838_n2628.n29 185
R18455 a_n2838_n2628.n28 a_n2838_n2628.n25 185
R18456 a_n2838_n2628.n4 a_n2838_n2628.n5 7.50266
R18457 a_n2838_n2628.n11 a_n2838_n2628.n10 185
R18458 a_n2838_n2628.n38 a_n2838_n2628.n20 185
R18459 a_n2838_n2628.n23 a_n2838_n2628.n39 185
R18460 a_n2838_n2628.n27 a_n2838_n2628.n26 185
R18461 a_n2838_n2628.n6 a_n2838_n2628.t0 150.026
R18462 a_n2838_n2628.n8 a_n2838_n2628.t2 150.026
R18463 a_n2838_n2628.t1 a_n2838_n2628.n12 150.026
R18464 a_n2838_n2628.n36 a_n2838_n2628.n31 114.974
R18465 a_n2838_n2628.n37 a_n2838_n2628.n36 114.974
R18466 a_n2838_n2628.n36 a_n2838_n2628.n35 110.77
R18467 a_n2838_n2628.n34 a_n2838_n2628.n13 104.615
R18468 a_n2838_n2628.n33 a_n2838_n2628.n13 104.615
R18469 a_n2838_n2628.n33 a_n2838_n2628.n32 104.615
R18470 a_n2838_n2628.n30 a_n2838_n2628.n16 104.615
R18471 a_n2838_n2628.n29 a_n2838_n2628.n16 104.615
R18472 a_n2838_n2628.n29 a_n2838_n2628.n28 104.615
R18473 a_n2838_n2628.n38 a_n2838_n2628.n10 104.615
R18474 a_n2838_n2628.n39 a_n2838_n2628.n38 104.615
R18475 a_n2838_n2628.n39 a_n2838_n2628.n26 104.615
R18476 a_n2838_n2628.n32 a_n2838_n2628.t0 52.3082
R18477 a_n2838_n2628.n28 a_n2838_n2628.t2 52.3082
R18478 a_n2838_n2628.t1 a_n2838_n2628.n26 52.3082
R18479 a_n2838_n2628.n24 a_n2838_n2628.n6 5.10304
R18480 a_n2838_n2628.n25 a_n2838_n2628.n8 5.10304
R18481 a_n2838_n2628.n12 a_n2838_n2628.n27 5.10304
R18482 a_n2838_n2628.n21 a_n2838_n2628.n24 12.8005
R18483 a_n2838_n2628.n22 a_n2838_n2628.n25 12.8005
R18484 a_n2838_n2628.n27 a_n2838_n2628.n23 12.8005
R18485 a_n2838_n2628.n6 a_n2838_n2628.n0 4.35729
R18486 a_n2838_n2628.n8 a_n2838_n2628.n2 4.35729
R18487 a_n2838_n2628.n4 a_n2838_n2628.n12 4.35729
R18488 a_n2838_n2628.n4 a_n2838_n2628.n11 3.56777
R18489 a_n2838_n2628.n9 a_n2838_n2628.n2 3.56777
R18490 a_n2838_n2628.n7 a_n2838_n2628.n0 3.56777
R18491 a_n2838_n2628.n15 a_n2838_n2628.n14 4.008
R18492 a_n2838_n2628.n18 a_n2838_n2628.n17 4.008
R18493 a_n2838_n2628.n20 a_n2838_n2628.n19 4.008
R18494 a_n2838_n2628.n7 a_n2838_n2628.n14 11.249
R18495 a_n2838_n2628.n9 a_n2838_n2628.n17 11.249
R18496 a_n2838_n2628.n20 a_n2838_n2628.n11 11.249
R18497 a_n2838_n2628.n23 a_n2838_n2628.n19 3.73143
R18498 a_n2838_n2628.n18 a_n2838_n2628.n22 3.73143
R18499 a_n2838_n2628.n15 a_n2838_n2628.n21 3.73143
R18500 a_n2838_n2628.n35 a_n2838_n2628.n6 9.45567
R18501 a_n2838_n2628.n31 a_n2838_n2628.n8 9.45567
R18502 a_n2838_n2628.n37 a_n2838_n2628.n12 9.45567
R18503 a_n2838_n2628.n15 a_n2838_n2628.n6 5.53918
R18504 a_n2838_n2628.n18 a_n2838_n2628.n8 5.53918
R18505 a_n2838_n2628.n19 a_n2838_n2628.n12 5.53918
R18506 a_n2838_n2628.n35 a_n2838_n2628.n1 10.0664
R18507 a_n2838_n2628.n31 a_n2838_n2628.n3 10.0664
R18508 a_n2838_n2628.n5 a_n2838_n2628.n37 10.0664
R18509 a_n4284_n2628.n30 a_n4284_n2628.n1 215.245
R18510 a_n4284_n2628.n34 a_n4284_n2628.n3 215.245
R18511 a_n4284_n2628.n10 a_n4284_n2628.n5 215.245
R18512 a_n4284_n2628.n0 a_n4284_n2628.n1 7.50266
R18513 a_n4284_n2628.n30 a_n4284_n2628.n7 185
R18514 a_n4284_n2628.n14 a_n4284_n2628.n13 185
R18515 a_n4284_n2628.n21 a_n4284_n2628.n29 185
R18516 a_n4284_n2628.n28 a_n4284_n2628.n24 185
R18517 a_n4284_n2628.n2 a_n4284_n2628.n3 7.50266
R18518 a_n4284_n2628.n34 a_n4284_n2628.n9 185
R18519 a_n4284_n2628.n17 a_n4284_n2628.n16 185
R18520 a_n4284_n2628.n22 a_n4284_n2628.n33 185
R18521 a_n4284_n2628.n32 a_n4284_n2628.n25 185
R18522 a_n4284_n2628.n4 a_n4284_n2628.n5 7.50266
R18523 a_n4284_n2628.n11 a_n4284_n2628.n10 185
R18524 a_n4284_n2628.n38 a_n4284_n2628.n20 185
R18525 a_n4284_n2628.n23 a_n4284_n2628.n39 185
R18526 a_n4284_n2628.n27 a_n4284_n2628.n26 185
R18527 a_n4284_n2628.n6 a_n4284_n2628.t2 150.026
R18528 a_n4284_n2628.n8 a_n4284_n2628.t0 150.026
R18529 a_n4284_n2628.t1 a_n4284_n2628.n12 150.026
R18530 a_n4284_n2628.n30 a_n4284_n2628.n13 104.615
R18531 a_n4284_n2628.n29 a_n4284_n2628.n13 104.615
R18532 a_n4284_n2628.n29 a_n4284_n2628.n28 104.615
R18533 a_n4284_n2628.n34 a_n4284_n2628.n16 104.615
R18534 a_n4284_n2628.n33 a_n4284_n2628.n16 104.615
R18535 a_n4284_n2628.n33 a_n4284_n2628.n32 104.615
R18536 a_n4284_n2628.n38 a_n4284_n2628.n10 104.615
R18537 a_n4284_n2628.n39 a_n4284_n2628.n38 104.615
R18538 a_n4284_n2628.n39 a_n4284_n2628.n26 104.615
R18539 a_n4284_n2628.n28 a_n4284_n2628.t2 52.3082
R18540 a_n4284_n2628.n32 a_n4284_n2628.t0 52.3082
R18541 a_n4284_n2628.t1 a_n4284_n2628.n26 52.3082
R18542 a_n4284_n2628.n36 a_n4284_n2628.n31 46.707
R18543 a_n4284_n2628.n37 a_n4284_n2628.n36 46.707
R18544 a_n4284_n2628.n36 a_n4284_n2628.n35 42.5035
R18545 a_n4284_n2628.n24 a_n4284_n2628.n6 5.10304
R18546 a_n4284_n2628.n25 a_n4284_n2628.n8 5.10304
R18547 a_n4284_n2628.n12 a_n4284_n2628.n27 5.10304
R18548 a_n4284_n2628.n21 a_n4284_n2628.n24 12.8005
R18549 a_n4284_n2628.n22 a_n4284_n2628.n25 12.8005
R18550 a_n4284_n2628.n27 a_n4284_n2628.n23 12.8005
R18551 a_n4284_n2628.n6 a_n4284_n2628.n0 4.35729
R18552 a_n4284_n2628.n8 a_n4284_n2628.n2 4.35729
R18553 a_n4284_n2628.n4 a_n4284_n2628.n12 4.35729
R18554 a_n4284_n2628.n4 a_n4284_n2628.n11 3.56777
R18555 a_n4284_n2628.n9 a_n4284_n2628.n2 3.56777
R18556 a_n4284_n2628.n7 a_n4284_n2628.n0 3.56777
R18557 a_n4284_n2628.n15 a_n4284_n2628.n14 4.008
R18558 a_n4284_n2628.n18 a_n4284_n2628.n17 4.008
R18559 a_n4284_n2628.n20 a_n4284_n2628.n19 4.008
R18560 a_n4284_n2628.n7 a_n4284_n2628.n14 11.249
R18561 a_n4284_n2628.n9 a_n4284_n2628.n17 11.249
R18562 a_n4284_n2628.n20 a_n4284_n2628.n11 11.249
R18563 a_n4284_n2628.n23 a_n4284_n2628.n19 3.73143
R18564 a_n4284_n2628.n18 a_n4284_n2628.n22 3.73143
R18565 a_n4284_n2628.n15 a_n4284_n2628.n21 3.73143
R18566 a_n4284_n2628.n31 a_n4284_n2628.n6 9.45567
R18567 a_n4284_n2628.n35 a_n4284_n2628.n8 9.45567
R18568 a_n4284_n2628.n37 a_n4284_n2628.n12 9.45567
R18569 a_n4284_n2628.n15 a_n4284_n2628.n6 5.53918
R18570 a_n4284_n2628.n18 a_n4284_n2628.n8 5.53918
R18571 a_n4284_n2628.n19 a_n4284_n2628.n12 5.53918
R18572 a_n4284_n2628.n31 a_n4284_n2628.n1 10.0664
R18573 a_n4284_n2628.n35 a_n4284_n2628.n3 10.0664
R18574 a_n4284_n2628.n5 a_n4284_n2628.n37 10.0664
C0 VP VN 9.65165f
C1 VOUT CS_BIAS 25.108599f
C2 VP CS_BIAS 0.348579f
C3 VP DIFFPAIR_BIAS 0.01402f
C4 VN CS_BIAS 0.274753f
C5 VN DIFFPAIR_BIAS 0.01402f
C6 a_8541_8735# VDD 1.42517f
C7 VDD VOUT 18.403198f
C8 a_n9553_8735# VDD 1.42571f
C9 VOUT VP 3.53664f
C10 VDD VN 0.143758f
C11 VOUT VN 0.930007f
C12 DIFFPAIR_BIAS GND 32.17023f
C13 CS_BIAS GND 0.123317p
C14 VN GND 28.2066f
C15 VP GND 23.95313f
C16 VOUT GND 72.462234f
C17 VDD GND 0.408151p
C18 a_8541_8735# GND 0.544554f
C19 a_n9553_8735# GND 0.544554f
C20 a_n4284_n2628.n0 GND 0.010941f
C21 a_n4284_n2628.n1 GND 0.048872f
C22 a_n4284_n2628.n2 GND 0.010941f
C23 a_n4284_n2628.n3 GND 0.048872f
C24 a_n4284_n2628.n4 GND 0.010941f
C25 a_n4284_n2628.n5 GND 0.048872f
C26 a_n4284_n2628.n6 GND 0.530141f
C27 a_n4284_n2628.n7 GND 0.022157f
C28 a_n4284_n2628.n8 GND 0.530141f
C29 a_n4284_n2628.n9 GND 0.022157f
C30 a_n4284_n2628.n10 GND 0.053003f
C31 a_n4284_n2628.n11 GND 0.022157f
C32 a_n4284_n2628.n12 GND 0.530141f
C33 a_n4284_n2628.t0 GND 0.04293f
C34 a_n4284_n2628.t2 GND 0.04293f
C35 a_n4284_n2628.n13 GND 0.025437f
C36 a_n4284_n2628.n14 GND 0.022157f
C37 a_n4284_n2628.n16 GND 0.025437f
C38 a_n4284_n2628.n17 GND 0.022157f
C39 a_n4284_n2628.n20 GND 0.022157f
C40 a_n4284_n2628.n21 GND 0.022157f
C41 a_n4284_n2628.n22 GND 0.022157f
C42 a_n4284_n2628.n23 GND 0.022157f
C43 a_n4284_n2628.n24 GND 0.025774f
C44 a_n4284_n2628.n25 GND 0.025774f
C45 a_n4284_n2628.n26 GND 0.019078f
C46 a_n4284_n2628.n27 GND 0.025774f
C47 a_n4284_n2628.n28 GND 0.019078f
C48 a_n4284_n2628.n29 GND 0.025437f
C49 a_n4284_n2628.n30 GND 0.053003f
C50 a_n4284_n2628.n31 GND 0.188019f
C51 a_n4284_n2628.n32 GND 0.019078f
C52 a_n4284_n2628.n33 GND 0.025437f
C53 a_n4284_n2628.n34 GND 0.053003f
C54 a_n4284_n2628.n35 GND 0.105233f
C55 a_n4284_n2628.n36 GND 3.88858f
C56 a_n4284_n2628.n37 GND 0.273912f
C57 a_n4284_n2628.n38 GND 0.025437f
C58 a_n4284_n2628.n39 GND 0.025437f
C59 a_n4284_n2628.t1 GND 0.04293f
C60 a_n2838_n2628.n0 GND 0.014536f
C61 a_n2838_n2628.n1 GND 0.06493f
C62 a_n2838_n2628.n2 GND 0.014536f
C63 a_n2838_n2628.n3 GND 0.06493f
C64 a_n2838_n2628.n4 GND 0.014536f
C65 a_n2838_n2628.n5 GND 0.06493f
C66 a_n2838_n2628.n6 GND 0.704331f
C67 a_n2838_n2628.n7 GND 0.029437f
C68 a_n2838_n2628.n8 GND 0.704331f
C69 a_n2838_n2628.n9 GND 0.029437f
C70 a_n2838_n2628.n10 GND 0.070419f
C71 a_n2838_n2628.n11 GND 0.029437f
C72 a_n2838_n2628.n12 GND 0.704331f
C73 a_n2838_n2628.t2 GND 0.057035f
C74 a_n2838_n2628.t0 GND 0.057035f
C75 a_n2838_n2628.n13 GND 0.033795f
C76 a_n2838_n2628.n14 GND 0.029437f
C77 a_n2838_n2628.n16 GND 0.033795f
C78 a_n2838_n2628.n17 GND 0.029437f
C79 a_n2838_n2628.n20 GND 0.029437f
C80 a_n2838_n2628.n21 GND 0.029437f
C81 a_n2838_n2628.n22 GND 0.029437f
C82 a_n2838_n2628.n23 GND 0.029437f
C83 a_n2838_n2628.n24 GND 0.034242f
C84 a_n2838_n2628.n25 GND 0.034242f
C85 a_n2838_n2628.n26 GND 0.025346f
C86 a_n2838_n2628.n27 GND 0.034242f
C87 a_n2838_n2628.n28 GND 0.025346f
C88 a_n2838_n2628.n29 GND 0.033795f
C89 a_n2838_n2628.n30 GND 0.070419f
C90 a_n2838_n2628.n31 GND 0.215292f
C91 a_n2838_n2628.n32 GND 0.025346f
C92 a_n2838_n2628.n33 GND 0.033795f
C93 a_n2838_n2628.n34 GND 0.070419f
C94 a_n2838_n2628.n35 GND 0.153731f
C95 a_n2838_n2628.n36 GND 5.32388f
C96 a_n2838_n2628.n37 GND 0.226872f
C97 a_n2838_n2628.n38 GND 0.033795f
C98 a_n2838_n2628.n39 GND 0.033795f
C99 a_n2838_n2628.t1 GND 0.057035f
C100 DIFFPAIR_BIAS.t7 GND 1.01926f
C101 DIFFPAIR_BIAS.t8 GND 0.976948f
C102 DIFFPAIR_BIAS.t6 GND 0.976948f
C103 DIFFPAIR_BIAS.n0 GND 0.004953f
C104 DIFFPAIR_BIAS.n1 GND 0.003628f
C105 DIFFPAIR_BIAS.n2 GND 0.00195f
C106 DIFFPAIR_BIAS.n3 GND 0.004608f
C107 DIFFPAIR_BIAS.n4 GND 0.002064f
C108 DIFFPAIR_BIAS.n5 GND 0.06254f
C109 DIFFPAIR_BIAS.n6 GND 0.00195f
C110 DIFFPAIR_BIAS.t1 GND 0.007556f
C111 DIFFPAIR_BIAS.n7 GND 0.014349f
C112 DIFFPAIR_BIAS.n8 GND 0.002719f
C113 DIFFPAIR_BIAS.n9 GND 0.003456f
C114 DIFFPAIR_BIAS.n10 GND 0.004608f
C115 DIFFPAIR_BIAS.n11 GND 0.002064f
C116 DIFFPAIR_BIAS.n12 GND 0.00195f
C117 DIFFPAIR_BIAS.n13 GND 0.003628f
C118 DIFFPAIR_BIAS.n14 GND 0.003628f
C119 DIFFPAIR_BIAS.n15 GND 0.00195f
C120 DIFFPAIR_BIAS.n16 GND 0.002064f
C121 DIFFPAIR_BIAS.n17 GND 0.004608f
C122 DIFFPAIR_BIAS.n18 GND 0.009716f
C123 DIFFPAIR_BIAS.n19 GND 0.002064f
C124 DIFFPAIR_BIAS.n20 GND 0.00195f
C125 DIFFPAIR_BIAS.n21 GND 0.008485f
C126 DIFFPAIR_BIAS.n22 GND 0.028225f
C127 DIFFPAIR_BIAS.n23 GND 0.004953f
C128 DIFFPAIR_BIAS.n24 GND 0.003628f
C129 DIFFPAIR_BIAS.n25 GND 0.00195f
C130 DIFFPAIR_BIAS.n26 GND 0.004608f
C131 DIFFPAIR_BIAS.n27 GND 0.002064f
C132 DIFFPAIR_BIAS.n28 GND 0.06254f
C133 DIFFPAIR_BIAS.n29 GND 0.00195f
C134 DIFFPAIR_BIAS.t5 GND 0.007556f
C135 DIFFPAIR_BIAS.n30 GND 0.014349f
C136 DIFFPAIR_BIAS.n31 GND 0.002719f
C137 DIFFPAIR_BIAS.n32 GND 0.003456f
C138 DIFFPAIR_BIAS.n33 GND 0.004608f
C139 DIFFPAIR_BIAS.n34 GND 0.002064f
C140 DIFFPAIR_BIAS.n35 GND 0.00195f
C141 DIFFPAIR_BIAS.n36 GND 0.003628f
C142 DIFFPAIR_BIAS.n37 GND 0.003628f
C143 DIFFPAIR_BIAS.n38 GND 0.00195f
C144 DIFFPAIR_BIAS.n39 GND 0.002064f
C145 DIFFPAIR_BIAS.n40 GND 0.004608f
C146 DIFFPAIR_BIAS.n41 GND 0.009716f
C147 DIFFPAIR_BIAS.n42 GND 0.002064f
C148 DIFFPAIR_BIAS.n43 GND 0.00195f
C149 DIFFPAIR_BIAS.n44 GND 0.008485f
C150 DIFFPAIR_BIAS.n45 GND 0.015054f
C151 DIFFPAIR_BIAS.n46 GND 0.464448f
C152 DIFFPAIR_BIAS.n47 GND 0.004953f
C153 DIFFPAIR_BIAS.n48 GND 0.003628f
C154 DIFFPAIR_BIAS.n49 GND 0.00195f
C155 DIFFPAIR_BIAS.n50 GND 0.004608f
C156 DIFFPAIR_BIAS.n51 GND 0.002064f
C157 DIFFPAIR_BIAS.n52 GND 0.06254f
C158 DIFFPAIR_BIAS.n53 GND 0.00195f
C159 DIFFPAIR_BIAS.t3 GND 0.007556f
C160 DIFFPAIR_BIAS.n54 GND 0.014349f
C161 DIFFPAIR_BIAS.n55 GND 0.002719f
C162 DIFFPAIR_BIAS.n56 GND 0.003456f
C163 DIFFPAIR_BIAS.n57 GND 0.004608f
C164 DIFFPAIR_BIAS.n58 GND 0.002064f
C165 DIFFPAIR_BIAS.n59 GND 0.00195f
C166 DIFFPAIR_BIAS.n60 GND 0.003628f
C167 DIFFPAIR_BIAS.n61 GND 0.003628f
C168 DIFFPAIR_BIAS.n62 GND 0.00195f
C169 DIFFPAIR_BIAS.n63 GND 0.002064f
C170 DIFFPAIR_BIAS.n64 GND 0.004608f
C171 DIFFPAIR_BIAS.n65 GND 0.009716f
C172 DIFFPAIR_BIAS.n66 GND 0.002064f
C173 DIFFPAIR_BIAS.n67 GND 0.00195f
C174 DIFFPAIR_BIAS.n68 GND 0.008485f
C175 DIFFPAIR_BIAS.n69 GND 0.015054f
C176 DIFFPAIR_BIAS.n70 GND 0.250538f
C177 DIFFPAIR_BIAS.t2 GND 0.958021f
C178 DIFFPAIR_BIAS.t4 GND 0.958021f
C179 DIFFPAIR_BIAS.t0 GND 1.00798f
C180 DIFFPAIR_BIAS.n71 GND 1.20468f
C181 DIFFPAIR_BIAS.n72 GND 0.677808f
C182 DIFFPAIR_BIAS.n73 GND 0.582856f
C183 DIFFPAIR_BIAS.n74 GND 0.627104f
C184 DIFFPAIR_BIAS.n75 GND 0.531532f
C185 DIFFPAIR_BIAS.n76 GND 0.929837f
C186 VN.t3 GND 0.946763f
C187 VN.t2 GND 1.15252f
C188 VN.n0 GND 1.40068f
C189 VN.t0 GND 0.02016f
C190 VN.t1 GND 0.020037f
C191 VN.n1 GND 0.102363f
C192 VN.n2 GND 1.73607f
C193 a_n12120_6849.n0 GND 0.209893f
C194 a_n12120_6849.n1 GND 0.209894f
C195 a_n12120_6849.t6 GND 0.031001f
C196 a_n12120_6849.t5 GND 0.031001f
C197 a_n12120_6849.t4 GND 0.031001f
C198 a_n12120_6849.n2 GND 0.173914f
C199 a_n12120_6849.t3 GND 0.031001f
C200 a_n12120_6849.t2 GND 0.031001f
C201 a_n12120_6849.n3 GND 0.158934f
C202 a_n12120_6849.n4 GND 2.38935f
C203 a_n12120_6849.n5 GND 0.020523f
C204 a_n12120_6849.n6 GND 0.007556f
C205 a_n12120_6849.n7 GND 0.013394f
C206 a_n12120_6849.n8 GND 0.012504f
C207 a_n12120_6849.t1 GND 0.031195f
C208 a_n12120_6849.n9 GND 0.056531f
C209 a_n12120_6849.n10 GND 0.007556f
C210 a_n12120_6849.n11 GND 0.008f
C211 a_n12120_6849.n12 GND 0.017859f
C212 a_n12120_6849.n13 GND 0.040004f
C213 a_n12120_6849.n14 GND 0.008f
C214 a_n12120_6849.n15 GND 0.007556f
C215 a_n12120_6849.n16 GND 0.034564f
C216 a_n12120_6849.n17 GND 0.020523f
C217 a_n12120_6849.n18 GND 0.007556f
C218 a_n12120_6849.n19 GND 0.013394f
C219 a_n12120_6849.n20 GND 0.012504f
C220 a_n12120_6849.t0 GND 0.031195f
C221 a_n12120_6849.n21 GND 0.056531f
C222 a_n12120_6849.n22 GND 0.007556f
C223 a_n12120_6849.n23 GND 0.008f
C224 a_n12120_6849.n24 GND 0.017859f
C225 a_n12120_6849.n25 GND 0.040004f
C226 a_n12120_6849.n26 GND 0.008f
C227 a_n12120_6849.n27 GND 0.007556f
C228 a_n12120_6849.n28 GND 0.420855f
C229 a_n12120_6849.n29 GND 2.0809f
C230 a_n12120_6849.t15 GND 2.00804f
C231 a_n12120_6849.t12 GND 1.97782f
C232 a_n12120_6849.n30 GND 2.01396f
C233 a_n12120_6849.t13 GND 1.97782f
C234 a_n12120_6849.n31 GND 3.10266f
C235 a_n12120_6849.t14 GND 2.00803f
C236 a_n12120_6849.t11 GND 1.97781f
C237 a_n12120_6849.n32 GND 2.01398f
C238 a_n12120_6849.t10 GND 1.97781f
C239 a_n12120_6849.n33 GND 2.7377f
C240 a_n12120_6849.n34 GND 19.8504f
C241 a_n12120_6849.n35 GND 3.26759f
C242 a_n12120_6849.n36 GND 4.13936f
C243 a_n12120_6849.t8 GND 0.031001f
C244 a_n12120_6849.t7 GND 0.031001f
C245 a_n12120_6849.n37 GND 0.173913f
C246 a_n12120_6849.n38 GND 2.8265f
C247 a_n12120_6849.n39 GND 0.158934f
C248 a_n12120_6849.t9 GND 0.031001f
C249 a_n1578_n2628.n0 GND 0.048227f
C250 a_n1578_n2628.n1 GND 0.037892f
C251 a_n1578_n2628.n2 GND 0.048227f
C252 a_n1578_n2628.n3 GND 0.037892f
C253 a_n1578_n2628.n4 GND 0.047114f
C254 a_n1578_n2628.n5 GND 0.039246f
C255 a_n1578_n2628.n6 GND 2.83601f
C256 a_n1578_n2628.n8 GND 1.1779f
C257 a_n1578_n2628.n9 GND 2.43613f
C258 a_n1578_n2628.n10 GND 0.009204f
C259 a_n1578_n2628.n11 GND 0.041114f
C260 a_n1578_n2628.n12 GND 0.009204f
C261 a_n1578_n2628.n13 GND 0.041114f
C262 a_n1578_n2628.n14 GND 0.009204f
C263 a_n1578_n2628.n15 GND 0.041114f
C264 a_n1578_n2628.n16 GND 1.45774f
C265 a_n1578_n2628.n17 GND 0.016273f
C266 a_n1578_n2628.n18 GND 0.021056f
C267 a_n1578_n2628.n19 GND 0.319241f
C268 a_n1578_n2628.n20 GND 0.016273f
C269 a_n1578_n2628.n21 GND 0.021056f
C270 a_n1578_n2628.n22 GND 0.319241f
C271 a_n1578_n2628.n23 GND 0.016273f
C272 a_n1578_n2628.n24 GND 0.021056f
C273 a_n1578_n2628.n25 GND 0.319241f
C274 a_n1578_n2628.n26 GND 0.319241f
C275 a_n1578_n2628.n27 GND 0.021056f
C276 a_n1578_n2628.n28 GND 0.445989f
C277 a_n1578_n2628.n29 GND 0.01864f
C278 a_n1578_n2628.n30 GND 0.445989f
C279 a_n1578_n2628.n31 GND 0.01864f
C280 a_n1578_n2628.n32 GND 0.445989f
C281 a_n1578_n2628.n33 GND 0.01864f
C282 a_n1578_n2628.t3 GND 0.036115f
C283 a_n1578_n2628.t1 GND 0.036115f
C284 a_n1578_n2628.t2 GND 0.036115f
C285 a_n1578_n2628.n34 GND 0.021399f
C286 a_n1578_n2628.n35 GND 0.01864f
C287 a_n1578_n2628.n37 GND 0.021399f
C288 a_n1578_n2628.n38 GND 0.01864f
C289 a_n1578_n2628.n40 GND 0.021399f
C290 a_n1578_n2628.n41 GND 0.01864f
C291 a_n1578_n2628.n43 GND 0.01864f
C292 a_n1578_n2628.n44 GND 0.01864f
C293 a_n1578_n2628.n45 GND 0.01864f
C294 a_n1578_n2628.n46 GND 0.021683f
C295 a_n1578_n2628.n47 GND 0.021683f
C296 a_n1578_n2628.n48 GND 0.021683f
C297 a_n1578_n2628.n49 GND 0.013827f
C298 a_n1578_n2628.n50 GND 0.016273f
C299 a_n1578_n2628.n51 GND 0.01605f
C300 a_n1578_n2628.n52 GND 0.021399f
C301 a_n1578_n2628.n53 GND 0.04459f
C302 a_n1578_n2628.n54 GND 0.116234f
C303 a_n1578_n2628.n55 GND 0.01605f
C304 a_n1578_n2628.n56 GND 0.021399f
C305 a_n1578_n2628.n57 GND 0.04459f
C306 a_n1578_n2628.n58 GND 0.111985f
C307 a_n1578_n2628.n59 GND 0.01605f
C308 a_n1578_n2628.n60 GND 0.021399f
C309 a_n1578_n2628.n61 GND 0.04459f
C310 a_n1578_n2628.n62 GND 0.111985f
C311 a_n1578_n2628.n63 GND 0.013827f
C312 a_n1578_n2628.t0 GND 0.037379f
C313 a_n1578_n2628.n64 GND 0.012344f
C314 a_n1578_n2628.n65 GND 0.04595f
C315 a_n1578_n2628.n66 GND 0.013827f
C316 a_n1578_n2628.t6 GND 0.037379f
C317 a_n1578_n2628.n67 GND 0.012344f
C318 a_n1578_n2628.n68 GND 0.04595f
C319 a_n1578_n2628.n69 GND 0.024591f
C320 a_n1578_n2628.n70 GND 0.009054f
C321 a_n1578_n2628.t4 GND 0.037379f
C322 a_n1578_n2628.n71 GND 0.012344f
C323 a_n1578_n2628.n72 GND 0.021399f
C324 a_n1578_n2628.n73 GND 0.047935f
C325 a_n1578_n2628.n74 GND 0.009586f
C326 a_n1578_n2628.n75 GND 0.009054f
C327 a_n1578_n2628.n76 GND 0.026899f
C328 a_n1578_n2628.n77 GND 0.04595f
C329 a_n1578_n2628.n78 GND 0.012344f
C330 a_n1578_n2628.t5 GND 0.037379f
C331 VOUT.t44 GND 0.199457f
C332 VOUT.t45 GND 0.193241f
C333 VOUT.n0 GND 0.519384f
C334 VOUT.t42 GND 0.193241f
C335 VOUT.n1 GND 0.369833f
C336 VOUT.n2 GND 5.996f
C337 VOUT.t49 GND 10.2157f
C338 VOUT.n3 GND 6.8611f
C339 VOUT.t48 GND 10.3914f
C340 VOUT.t47 GND 10.442699f
C341 VOUT.n4 GND 7.79865f
C342 VOUT.n5 GND 7.856939f
C343 VOUT.t46 GND 10.2157f
C344 VOUT.n6 GND 3.34447f
C345 VOUT.n7 GND 7.91067f
C346 VOUT.n8 GND 1.76633f
C347 VOUT.t41 GND 0.200777f
C348 VOUT.t43 GND 0.194676f
C349 VOUT.n9 GND 0.516629f
C350 VOUT.t40 GND 0.194676f
C351 VOUT.n10 GND 0.368398f
C352 VOUT.n11 GND 7.829999f
C353 VOUT.t39 GND 0.010162f
C354 VOUT.t14 GND 0.010162f
C355 VOUT.n12 GND 0.077619f
C356 VOUT.t7 GND 0.010162f
C357 VOUT.t11 GND 0.010162f
C358 VOUT.n13 GND 0.071807f
C359 VOUT.n14 GND 0.334729f
C360 VOUT.t34 GND 0.010162f
C361 VOUT.t17 GND 0.010162f
C362 VOUT.n15 GND 0.077619f
C363 VOUT.t13 GND 0.010162f
C364 VOUT.t20 GND 0.010162f
C365 VOUT.n16 GND 0.071807f
C366 VOUT.n17 GND 0.321814f
C367 VOUT.n18 GND 0.137876f
C368 VOUT.t29 GND 0.010162f
C369 VOUT.t28 GND 0.010162f
C370 VOUT.n19 GND 0.077619f
C371 VOUT.t6 GND 0.010162f
C372 VOUT.t16 GND 0.010162f
C373 VOUT.n20 GND 0.071807f
C374 VOUT.n21 GND 0.321814f
C375 VOUT.n22 GND 0.091154f
C376 VOUT.t10 GND 0.010162f
C377 VOUT.t33 GND 0.010162f
C378 VOUT.n23 GND 0.077619f
C379 VOUT.t31 GND 0.010162f
C380 VOUT.t0 GND 0.010162f
C381 VOUT.n24 GND 0.071807f
C382 VOUT.n25 GND 0.321814f
C383 VOUT.n26 GND 0.091154f
C384 VOUT.t4 GND 0.010162f
C385 VOUT.t27 GND 0.010162f
C386 VOUT.n27 GND 0.077619f
C387 VOUT.t23 GND 0.010162f
C388 VOUT.t35 GND 0.010162f
C389 VOUT.n28 GND 0.071807f
C390 VOUT.n29 GND 0.321814f
C391 VOUT.n30 GND 0.189965f
C392 VOUT.n31 GND 7.606431f
C393 VOUT.t22 GND 0.010162f
C394 VOUT.t2 GND 0.010162f
C395 VOUT.n32 GND 0.077619f
C396 VOUT.t32 GND 0.010162f
C397 VOUT.t12 GND 0.010162f
C398 VOUT.n33 GND 0.071807f
C399 VOUT.n34 GND 0.334729f
C400 VOUT.t18 GND 0.010162f
C401 VOUT.t8 GND 0.010162f
C402 VOUT.n35 GND 0.077619f
C403 VOUT.t37 GND 0.010162f
C404 VOUT.t25 GND 0.010162f
C405 VOUT.n36 GND 0.071807f
C406 VOUT.n37 GND 0.321814f
C407 VOUT.n38 GND 0.137876f
C408 VOUT.t26 GND 0.010162f
C409 VOUT.t19 GND 0.010162f
C410 VOUT.n39 GND 0.077619f
C411 VOUT.t5 GND 0.010162f
C412 VOUT.t38 GND 0.010162f
C413 VOUT.n40 GND 0.071807f
C414 VOUT.n41 GND 0.321814f
C415 VOUT.n42 GND 0.091154f
C416 VOUT.t36 GND 0.010162f
C417 VOUT.t24 GND 0.010162f
C418 VOUT.n43 GND 0.077619f
C419 VOUT.t15 GND 0.010162f
C420 VOUT.t3 GND 0.010162f
C421 VOUT.n44 GND 0.071807f
C422 VOUT.n45 GND 0.321814f
C423 VOUT.n46 GND 0.091154f
C424 VOUT.t30 GND 0.010162f
C425 VOUT.t21 GND 0.010162f
C426 VOUT.n47 GND 0.077619f
C427 VOUT.t9 GND 0.010162f
C428 VOUT.t1 GND 0.010162f
C429 VOUT.n48 GND 0.071807f
C430 VOUT.n49 GND 0.321814f
C431 VOUT.n50 GND 0.189965f
C432 VOUT.n51 GND 5.47683f
C433 VOUT.n52 GND 4.10141f
C434 CS_BIAS.t16 GND 0.143123f
C435 CS_BIAS.n0 GND 0.090069f
C436 CS_BIAS.n1 GND 0.00704f
C437 CS_BIAS.n2 GND 0.008376f
C438 CS_BIAS.n3 GND 0.00704f
C439 CS_BIAS.n4 GND 0.007642f
C440 CS_BIAS.n5 GND 0.00704f
C441 CS_BIAS.t41 GND 0.143123f
C442 CS_BIAS.n6 GND 0.061848f
C443 CS_BIAS.n7 GND 0.005686f
C444 CS_BIAS.t12 GND 0.143123f
C445 CS_BIAS.n8 GND 0.090069f
C446 CS_BIAS.n9 GND 0.00704f
C447 CS_BIAS.n10 GND 0.008376f
C448 CS_BIAS.n11 GND 0.00704f
C449 CS_BIAS.n12 GND 0.007642f
C450 CS_BIAS.n13 GND 0.00704f
C451 CS_BIAS.t6 GND 0.143123f
C452 CS_BIAS.n14 GND 0.061848f
C453 CS_BIAS.n15 GND 0.005686f
C454 CS_BIAS.n16 GND 0.00704f
C455 CS_BIAS.t0 GND 0.143123f
C456 CS_BIAS.n17 GND 0.088437f
C457 CS_BIAS.t2 GND 0.220418f
C458 CS_BIAS.n18 GND 0.091063f
C459 CS_BIAS.n19 GND 0.086627f
C460 CS_BIAS.n20 GND 0.012024f
C461 CS_BIAS.n21 GND 0.013056f
C462 CS_BIAS.n22 GND 0.013919f
C463 CS_BIAS.n23 GND 0.00704f
C464 CS_BIAS.n24 GND 0.00704f
C465 CS_BIAS.n25 GND 0.00704f
C466 CS_BIAS.n26 GND 0.013919f
C467 CS_BIAS.n27 GND 0.013056f
C468 CS_BIAS.n28 GND 0.012024f
C469 CS_BIAS.n29 GND 0.00704f
C470 CS_BIAS.n30 GND 0.00704f
C471 CS_BIAS.n31 GND 0.00704f
C472 CS_BIAS.n32 GND 0.013056f
C473 CS_BIAS.n33 GND 0.013056f
C474 CS_BIAS.n34 GND 0.01197f
C475 CS_BIAS.n35 GND 0.00704f
C476 CS_BIAS.n36 GND 0.00704f
C477 CS_BIAS.n37 GND 0.00704f
C478 CS_BIAS.n38 GND 0.013178f
C479 CS_BIAS.n39 GND 0.013056f
C480 CS_BIAS.n40 GND 0.009962f
C481 CS_BIAS.n41 GND 0.011361f
C482 CS_BIAS.n42 GND 0.065582f
C483 CS_BIAS.t13 GND 0.005209f
C484 CS_BIAS.t7 GND 0.005209f
C485 CS_BIAS.n43 GND 0.036806f
C486 CS_BIAS.n44 GND 0.086504f
C487 CS_BIAS.t1 GND 0.005209f
C488 CS_BIAS.t3 GND 0.005209f
C489 CS_BIAS.n45 GND 0.038017f
C490 CS_BIAS.n46 GND 0.137358f
C491 CS_BIAS.n47 GND 0.00704f
C492 CS_BIAS.t48 GND 0.143123f
C493 CS_BIAS.n48 GND 0.088437f
C494 CS_BIAS.t44 GND 0.220418f
C495 CS_BIAS.n49 GND 0.091063f
C496 CS_BIAS.n50 GND 0.086627f
C497 CS_BIAS.n51 GND 0.012024f
C498 CS_BIAS.n52 GND 0.013056f
C499 CS_BIAS.n53 GND 0.013919f
C500 CS_BIAS.n54 GND 0.007007f
C501 CS_BIAS.n55 GND 0.050893f
C502 CS_BIAS.n56 GND 0.007007f
C503 CS_BIAS.n57 GND 0.013919f
C504 CS_BIAS.n58 GND 0.013056f
C505 CS_BIAS.n59 GND 0.012024f
C506 CS_BIAS.n60 GND 0.00704f
C507 CS_BIAS.n61 GND 0.00704f
C508 CS_BIAS.n62 GND 0.00704f
C509 CS_BIAS.n63 GND 0.013056f
C510 CS_BIAS.n64 GND 0.013056f
C511 CS_BIAS.n65 GND 0.01197f
C512 CS_BIAS.n66 GND 0.00704f
C513 CS_BIAS.n67 GND 0.00704f
C514 CS_BIAS.n68 GND 0.00704f
C515 CS_BIAS.n69 GND 0.013178f
C516 CS_BIAS.n70 GND 0.013056f
C517 CS_BIAS.n71 GND 0.009962f
C518 CS_BIAS.n72 GND 0.011361f
C519 CS_BIAS.n73 GND 0.047902f
C520 CS_BIAS.t21 GND 0.143123f
C521 CS_BIAS.n74 GND 0.090069f
C522 CS_BIAS.n75 GND 0.00704f
C523 CS_BIAS.n76 GND 0.008376f
C524 CS_BIAS.n77 GND 0.00704f
C525 CS_BIAS.n78 GND 0.007642f
C526 CS_BIAS.n79 GND 0.00704f
C527 CS_BIAS.t38 GND 0.143123f
C528 CS_BIAS.n80 GND 0.061848f
C529 CS_BIAS.n81 GND 0.005686f
C530 CS_BIAS.n82 GND 0.00704f
C531 CS_BIAS.t42 GND 0.143123f
C532 CS_BIAS.n83 GND 0.088437f
C533 CS_BIAS.t35 GND 0.220418f
C534 CS_BIAS.n84 GND 0.091063f
C535 CS_BIAS.n85 GND 0.086627f
C536 CS_BIAS.n86 GND 0.012024f
C537 CS_BIAS.n87 GND 0.013056f
C538 CS_BIAS.n88 GND 0.013919f
C539 CS_BIAS.n89 GND 0.00704f
C540 CS_BIAS.n90 GND 0.00704f
C541 CS_BIAS.n91 GND 0.00704f
C542 CS_BIAS.n92 GND 0.013919f
C543 CS_BIAS.n93 GND 0.013056f
C544 CS_BIAS.n94 GND 0.012024f
C545 CS_BIAS.n95 GND 0.00704f
C546 CS_BIAS.n96 GND 0.00704f
C547 CS_BIAS.n97 GND 0.00704f
C548 CS_BIAS.n98 GND 0.013056f
C549 CS_BIAS.n99 GND 0.013056f
C550 CS_BIAS.n100 GND 0.01197f
C551 CS_BIAS.n101 GND 0.00704f
C552 CS_BIAS.n102 GND 0.00704f
C553 CS_BIAS.n103 GND 0.00704f
C554 CS_BIAS.n104 GND 0.013178f
C555 CS_BIAS.n105 GND 0.013056f
C556 CS_BIAS.n106 GND 0.009962f
C557 CS_BIAS.n107 GND 0.011361f
C558 CS_BIAS.n108 GND 0.041603f
C559 CS_BIAS.n109 GND 0.062571f
C560 CS_BIAS.t26 GND 0.143123f
C561 CS_BIAS.n110 GND 0.090069f
C562 CS_BIAS.n111 GND 0.00704f
C563 CS_BIAS.n112 GND 0.008376f
C564 CS_BIAS.n113 GND 0.00704f
C565 CS_BIAS.n114 GND 0.007642f
C566 CS_BIAS.n115 GND 0.00704f
C567 CS_BIAS.t27 GND 0.143123f
C568 CS_BIAS.n116 GND 0.061848f
C569 CS_BIAS.n117 GND 0.005686f
C570 CS_BIAS.n118 GND 0.00704f
C571 CS_BIAS.t49 GND 0.143123f
C572 CS_BIAS.n119 GND 0.088437f
C573 CS_BIAS.t39 GND 0.220418f
C574 CS_BIAS.n120 GND 0.091063f
C575 CS_BIAS.n121 GND 0.086627f
C576 CS_BIAS.n122 GND 0.012024f
C577 CS_BIAS.n123 GND 0.013056f
C578 CS_BIAS.n124 GND 0.013919f
C579 CS_BIAS.n125 GND 0.00704f
C580 CS_BIAS.n126 GND 0.00704f
C581 CS_BIAS.n127 GND 0.00704f
C582 CS_BIAS.n128 GND 0.013919f
C583 CS_BIAS.n129 GND 0.013056f
C584 CS_BIAS.n130 GND 0.012024f
C585 CS_BIAS.n131 GND 0.00704f
C586 CS_BIAS.n132 GND 0.00704f
C587 CS_BIAS.n133 GND 0.00704f
C588 CS_BIAS.n134 GND 0.013056f
C589 CS_BIAS.n135 GND 0.013056f
C590 CS_BIAS.n136 GND 0.01197f
C591 CS_BIAS.n137 GND 0.00704f
C592 CS_BIAS.n138 GND 0.00704f
C593 CS_BIAS.n139 GND 0.00704f
C594 CS_BIAS.n140 GND 0.013178f
C595 CS_BIAS.n141 GND 0.013056f
C596 CS_BIAS.n142 GND 0.009962f
C597 CS_BIAS.n143 GND 0.011361f
C598 CS_BIAS.n144 GND 0.041603f
C599 CS_BIAS.n145 GND 0.043626f
C600 CS_BIAS.t45 GND 0.143123f
C601 CS_BIAS.n146 GND 0.090069f
C602 CS_BIAS.n147 GND 0.00704f
C603 CS_BIAS.n148 GND 0.008376f
C604 CS_BIAS.n149 GND 0.00704f
C605 CS_BIAS.n150 GND 0.007642f
C606 CS_BIAS.n151 GND 0.00704f
C607 CS_BIAS.t22 GND 0.143123f
C608 CS_BIAS.n152 GND 0.061848f
C609 CS_BIAS.n153 GND 0.005686f
C610 CS_BIAS.n154 GND 0.00704f
C611 CS_BIAS.t24 GND 0.143123f
C612 CS_BIAS.n155 GND 0.088437f
C613 CS_BIAS.t55 GND 0.220418f
C614 CS_BIAS.n156 GND 0.091063f
C615 CS_BIAS.n157 GND 0.086627f
C616 CS_BIAS.n158 GND 0.012024f
C617 CS_BIAS.n159 GND 0.013056f
C618 CS_BIAS.n160 GND 0.013919f
C619 CS_BIAS.n161 GND 0.00704f
C620 CS_BIAS.n162 GND 0.00704f
C621 CS_BIAS.n163 GND 0.00704f
C622 CS_BIAS.n164 GND 0.013919f
C623 CS_BIAS.n165 GND 0.013056f
C624 CS_BIAS.n166 GND 0.012024f
C625 CS_BIAS.n167 GND 0.00704f
C626 CS_BIAS.n168 GND 0.00704f
C627 CS_BIAS.n169 GND 0.00704f
C628 CS_BIAS.n170 GND 0.013056f
C629 CS_BIAS.n171 GND 0.013056f
C630 CS_BIAS.n172 GND 0.01197f
C631 CS_BIAS.n173 GND 0.00704f
C632 CS_BIAS.n174 GND 0.00704f
C633 CS_BIAS.n175 GND 0.00704f
C634 CS_BIAS.n176 GND 0.013178f
C635 CS_BIAS.n177 GND 0.013056f
C636 CS_BIAS.n178 GND 0.009962f
C637 CS_BIAS.n179 GND 0.011361f
C638 CS_BIAS.n180 GND 0.041603f
C639 CS_BIAS.n181 GND 0.043626f
C640 CS_BIAS.t51 GND 0.143123f
C641 CS_BIAS.n182 GND 0.090069f
C642 CS_BIAS.n183 GND 0.00704f
C643 CS_BIAS.n184 GND 0.008376f
C644 CS_BIAS.n185 GND 0.00704f
C645 CS_BIAS.n186 GND 0.007642f
C646 CS_BIAS.n187 GND 0.00704f
C647 CS_BIAS.t28 GND 0.143123f
C648 CS_BIAS.n188 GND 0.061848f
C649 CS_BIAS.n189 GND 0.005686f
C650 CS_BIAS.n190 GND 0.00704f
C651 CS_BIAS.t32 GND 0.143123f
C652 CS_BIAS.n191 GND 0.088437f
C653 CS_BIAS.t20 GND 0.220418f
C654 CS_BIAS.n192 GND 0.091063f
C655 CS_BIAS.n193 GND 0.086627f
C656 CS_BIAS.n194 GND 0.012024f
C657 CS_BIAS.n195 GND 0.013056f
C658 CS_BIAS.n196 GND 0.013919f
C659 CS_BIAS.n197 GND 0.00704f
C660 CS_BIAS.n198 GND 0.00704f
C661 CS_BIAS.n199 GND 0.00704f
C662 CS_BIAS.n200 GND 0.013919f
C663 CS_BIAS.n201 GND 0.013056f
C664 CS_BIAS.n202 GND 0.012024f
C665 CS_BIAS.n203 GND 0.00704f
C666 CS_BIAS.n204 GND 0.00704f
C667 CS_BIAS.n205 GND 0.00704f
C668 CS_BIAS.n206 GND 0.013056f
C669 CS_BIAS.n207 GND 0.013056f
C670 CS_BIAS.n208 GND 0.01197f
C671 CS_BIAS.n209 GND 0.00704f
C672 CS_BIAS.n210 GND 0.00704f
C673 CS_BIAS.n211 GND 0.00704f
C674 CS_BIAS.n212 GND 0.013178f
C675 CS_BIAS.n213 GND 0.013056f
C676 CS_BIAS.n214 GND 0.009962f
C677 CS_BIAS.n215 GND 0.011361f
C678 CS_BIAS.n216 GND 0.041603f
C679 CS_BIAS.n217 GND 0.526665f
C680 CS_BIAS.t53 GND 0.143123f
C681 CS_BIAS.n218 GND 0.090069f
C682 CS_BIAS.n219 GND 0.00704f
C683 CS_BIAS.n220 GND 0.008376f
C684 CS_BIAS.n221 GND 0.00704f
C685 CS_BIAS.n222 GND 0.007642f
C686 CS_BIAS.n223 GND 0.00704f
C687 CS_BIAS.n224 GND 0.005686f
C688 CS_BIAS.n225 GND 0.00704f
C689 CS_BIAS.t43 GND 0.143123f
C690 CS_BIAS.n226 GND 0.088437f
C691 CS_BIAS.t23 GND 0.220418f
C692 CS_BIAS.n227 GND 0.091063f
C693 CS_BIAS.n228 GND 0.086627f
C694 CS_BIAS.n229 GND 0.012024f
C695 CS_BIAS.n230 GND 0.013056f
C696 CS_BIAS.n231 GND 0.013919f
C697 CS_BIAS.n232 GND 0.007007f
C698 CS_BIAS.t11 GND 0.005209f
C699 CS_BIAS.t5 GND 0.005209f
C700 CS_BIAS.n233 GND 0.038017f
C701 CS_BIAS.t14 GND 0.143123f
C702 CS_BIAS.n234 GND 0.090069f
C703 CS_BIAS.n235 GND 0.00704f
C704 CS_BIAS.n236 GND 0.008376f
C705 CS_BIAS.n237 GND 0.00704f
C706 CS_BIAS.n238 GND 0.007642f
C707 CS_BIAS.n239 GND 0.00704f
C708 CS_BIAS.n240 GND 0.005686f
C709 CS_BIAS.n241 GND 0.00704f
C710 CS_BIAS.t4 GND 0.143123f
C711 CS_BIAS.n242 GND 0.088437f
C712 CS_BIAS.t10 GND 0.220418f
C713 CS_BIAS.n243 GND 0.091063f
C714 CS_BIAS.n244 GND 0.086627f
C715 CS_BIAS.n245 GND 0.012024f
C716 CS_BIAS.n246 GND 0.013056f
C717 CS_BIAS.n247 GND 0.013919f
C718 CS_BIAS.n248 GND 0.00704f
C719 CS_BIAS.n249 GND 0.00704f
C720 CS_BIAS.n250 GND 0.00704f
C721 CS_BIAS.n251 GND 0.013919f
C722 CS_BIAS.n252 GND 0.013056f
C723 CS_BIAS.t8 GND 0.143123f
C724 CS_BIAS.n253 GND 0.061848f
C725 CS_BIAS.n254 GND 0.012024f
C726 CS_BIAS.n255 GND 0.00704f
C727 CS_BIAS.n256 GND 0.00704f
C728 CS_BIAS.n257 GND 0.00704f
C729 CS_BIAS.n258 GND 0.013056f
C730 CS_BIAS.n259 GND 0.013056f
C731 CS_BIAS.n260 GND 0.01197f
C732 CS_BIAS.n261 GND 0.00704f
C733 CS_BIAS.n262 GND 0.00704f
C734 CS_BIAS.n263 GND 0.00704f
C735 CS_BIAS.n264 GND 0.013178f
C736 CS_BIAS.n265 GND 0.013056f
C737 CS_BIAS.n266 GND 0.009962f
C738 CS_BIAS.n267 GND 0.011361f
C739 CS_BIAS.n268 GND 0.065582f
C740 CS_BIAS.t9 GND 0.005209f
C741 CS_BIAS.t15 GND 0.005209f
C742 CS_BIAS.n269 GND 0.036806f
C743 CS_BIAS.n270 GND 0.086504f
C744 CS_BIAS.n271 GND 0.137358f
C745 CS_BIAS.n272 GND 0.050893f
C746 CS_BIAS.n273 GND 0.007007f
C747 CS_BIAS.n274 GND 0.013919f
C748 CS_BIAS.n275 GND 0.013056f
C749 CS_BIAS.t33 GND 0.143123f
C750 CS_BIAS.n276 GND 0.061848f
C751 CS_BIAS.n277 GND 0.012024f
C752 CS_BIAS.n278 GND 0.00704f
C753 CS_BIAS.n279 GND 0.00704f
C754 CS_BIAS.n280 GND 0.00704f
C755 CS_BIAS.n281 GND 0.013056f
C756 CS_BIAS.n282 GND 0.013056f
C757 CS_BIAS.n283 GND 0.01197f
C758 CS_BIAS.n284 GND 0.00704f
C759 CS_BIAS.n285 GND 0.00704f
C760 CS_BIAS.n286 GND 0.00704f
C761 CS_BIAS.n287 GND 0.013178f
C762 CS_BIAS.n288 GND 0.013056f
C763 CS_BIAS.n289 GND 0.009962f
C764 CS_BIAS.n290 GND 0.011361f
C765 CS_BIAS.n291 GND 0.047902f
C766 CS_BIAS.t47 GND 0.143123f
C767 CS_BIAS.n292 GND 0.090069f
C768 CS_BIAS.n293 GND 0.00704f
C769 CS_BIAS.n294 GND 0.008376f
C770 CS_BIAS.n295 GND 0.00704f
C771 CS_BIAS.n296 GND 0.007642f
C772 CS_BIAS.n297 GND 0.00704f
C773 CS_BIAS.n298 GND 0.005686f
C774 CS_BIAS.n299 GND 0.00704f
C775 CS_BIAS.t30 GND 0.143123f
C776 CS_BIAS.n300 GND 0.088437f
C777 CS_BIAS.t18 GND 0.220418f
C778 CS_BIAS.n301 GND 0.091063f
C779 CS_BIAS.n302 GND 0.086627f
C780 CS_BIAS.n303 GND 0.012024f
C781 CS_BIAS.n304 GND 0.013056f
C782 CS_BIAS.n305 GND 0.013919f
C783 CS_BIAS.n306 GND 0.00704f
C784 CS_BIAS.n307 GND 0.00704f
C785 CS_BIAS.n308 GND 0.00704f
C786 CS_BIAS.n309 GND 0.013919f
C787 CS_BIAS.n310 GND 0.013056f
C788 CS_BIAS.t37 GND 0.143123f
C789 CS_BIAS.n311 GND 0.061848f
C790 CS_BIAS.n312 GND 0.012024f
C791 CS_BIAS.n313 GND 0.00704f
C792 CS_BIAS.n314 GND 0.00704f
C793 CS_BIAS.n315 GND 0.00704f
C794 CS_BIAS.n316 GND 0.013056f
C795 CS_BIAS.n317 GND 0.013056f
C796 CS_BIAS.n318 GND 0.01197f
C797 CS_BIAS.n319 GND 0.00704f
C798 CS_BIAS.n320 GND 0.00704f
C799 CS_BIAS.n321 GND 0.00704f
C800 CS_BIAS.n322 GND 0.013178f
C801 CS_BIAS.n323 GND 0.013056f
C802 CS_BIAS.n324 GND 0.009962f
C803 CS_BIAS.n325 GND 0.011361f
C804 CS_BIAS.n326 GND 0.041603f
C805 CS_BIAS.n327 GND 0.062571f
C806 CS_BIAS.t36 GND 0.143123f
C807 CS_BIAS.n328 GND 0.090069f
C808 CS_BIAS.n329 GND 0.00704f
C809 CS_BIAS.n330 GND 0.008376f
C810 CS_BIAS.n331 GND 0.00704f
C811 CS_BIAS.n332 GND 0.007642f
C812 CS_BIAS.n333 GND 0.00704f
C813 CS_BIAS.n334 GND 0.005686f
C814 CS_BIAS.n335 GND 0.00704f
C815 CS_BIAS.t17 GND 0.143123f
C816 CS_BIAS.n336 GND 0.088437f
C817 CS_BIAS.t50 GND 0.220418f
C818 CS_BIAS.n337 GND 0.091063f
C819 CS_BIAS.n338 GND 0.086627f
C820 CS_BIAS.n339 GND 0.012024f
C821 CS_BIAS.n340 GND 0.013056f
C822 CS_BIAS.n341 GND 0.013919f
C823 CS_BIAS.n342 GND 0.00704f
C824 CS_BIAS.n343 GND 0.00704f
C825 CS_BIAS.n344 GND 0.00704f
C826 CS_BIAS.n345 GND 0.013919f
C827 CS_BIAS.n346 GND 0.013056f
C828 CS_BIAS.t29 GND 0.143123f
C829 CS_BIAS.n347 GND 0.061848f
C830 CS_BIAS.n348 GND 0.012024f
C831 CS_BIAS.n349 GND 0.00704f
C832 CS_BIAS.n350 GND 0.00704f
C833 CS_BIAS.n351 GND 0.00704f
C834 CS_BIAS.n352 GND 0.013056f
C835 CS_BIAS.n353 GND 0.013056f
C836 CS_BIAS.n354 GND 0.01197f
C837 CS_BIAS.n355 GND 0.00704f
C838 CS_BIAS.n356 GND 0.00704f
C839 CS_BIAS.n357 GND 0.00704f
C840 CS_BIAS.n358 GND 0.013178f
C841 CS_BIAS.n359 GND 0.013056f
C842 CS_BIAS.n360 GND 0.009962f
C843 CS_BIAS.n361 GND 0.011361f
C844 CS_BIAS.n362 GND 0.041603f
C845 CS_BIAS.n363 GND 0.043626f
C846 CS_BIAS.t31 GND 0.143123f
C847 CS_BIAS.n364 GND 0.090069f
C848 CS_BIAS.n365 GND 0.00704f
C849 CS_BIAS.n366 GND 0.008376f
C850 CS_BIAS.n367 GND 0.00704f
C851 CS_BIAS.n368 GND 0.007642f
C852 CS_BIAS.n369 GND 0.00704f
C853 CS_BIAS.n370 GND 0.005686f
C854 CS_BIAS.n371 GND 0.00704f
C855 CS_BIAS.t52 GND 0.143123f
C856 CS_BIAS.n372 GND 0.088437f
C857 CS_BIAS.t40 GND 0.220418f
C858 CS_BIAS.n373 GND 0.091063f
C859 CS_BIAS.n374 GND 0.086627f
C860 CS_BIAS.n375 GND 0.012024f
C861 CS_BIAS.n376 GND 0.013056f
C862 CS_BIAS.n377 GND 0.013919f
C863 CS_BIAS.n378 GND 0.00704f
C864 CS_BIAS.n379 GND 0.00704f
C865 CS_BIAS.n380 GND 0.00704f
C866 CS_BIAS.n381 GND 0.013919f
C867 CS_BIAS.n382 GND 0.013056f
C868 CS_BIAS.t19 GND 0.143123f
C869 CS_BIAS.n383 GND 0.061848f
C870 CS_BIAS.n384 GND 0.012024f
C871 CS_BIAS.n385 GND 0.00704f
C872 CS_BIAS.n386 GND 0.00704f
C873 CS_BIAS.n387 GND 0.00704f
C874 CS_BIAS.n388 GND 0.013056f
C875 CS_BIAS.n389 GND 0.013056f
C876 CS_BIAS.n390 GND 0.01197f
C877 CS_BIAS.n391 GND 0.00704f
C878 CS_BIAS.n392 GND 0.00704f
C879 CS_BIAS.n393 GND 0.00704f
C880 CS_BIAS.n394 GND 0.013178f
C881 CS_BIAS.n395 GND 0.013056f
C882 CS_BIAS.n396 GND 0.009962f
C883 CS_BIAS.n397 GND 0.011361f
C884 CS_BIAS.n398 GND 0.041603f
C885 CS_BIAS.n399 GND 0.043626f
C886 CS_BIAS.t34 GND 0.143123f
C887 CS_BIAS.n400 GND 0.090069f
C888 CS_BIAS.n401 GND 0.00704f
C889 CS_BIAS.n402 GND 0.008376f
C890 CS_BIAS.n403 GND 0.00704f
C891 CS_BIAS.n404 GND 0.007642f
C892 CS_BIAS.n405 GND 0.00704f
C893 CS_BIAS.n406 GND 0.005686f
C894 CS_BIAS.n407 GND 0.00704f
C895 CS_BIAS.t54 GND 0.143123f
C896 CS_BIAS.n408 GND 0.088437f
C897 CS_BIAS.t46 GND 0.220418f
C898 CS_BIAS.n409 GND 0.091063f
C899 CS_BIAS.n410 GND 0.086627f
C900 CS_BIAS.n411 GND 0.012024f
C901 CS_BIAS.n412 GND 0.013056f
C902 CS_BIAS.n413 GND 0.013919f
C903 CS_BIAS.n414 GND 0.00704f
C904 CS_BIAS.n415 GND 0.00704f
C905 CS_BIAS.n416 GND 0.00704f
C906 CS_BIAS.n417 GND 0.013919f
C907 CS_BIAS.n418 GND 0.013056f
C908 CS_BIAS.t25 GND 0.143123f
C909 CS_BIAS.n419 GND 0.061848f
C910 CS_BIAS.n420 GND 0.012024f
C911 CS_BIAS.n421 GND 0.00704f
C912 CS_BIAS.n422 GND 0.00704f
C913 CS_BIAS.n423 GND 0.00704f
C914 CS_BIAS.n424 GND 0.013056f
C915 CS_BIAS.n425 GND 0.013056f
C916 CS_BIAS.n426 GND 0.01197f
C917 CS_BIAS.n427 GND 0.00704f
C918 CS_BIAS.n428 GND 0.00704f
C919 CS_BIAS.n429 GND 0.00704f
C920 CS_BIAS.n430 GND 0.013178f
C921 CS_BIAS.n431 GND 0.013056f
C922 CS_BIAS.n432 GND 0.009962f
C923 CS_BIAS.n433 GND 0.011361f
C924 CS_BIAS.n434 GND 0.041603f
C925 CS_BIAS.n435 GND 0.103959f
C926 CS_BIAS.n436 GND 4.24078f
C927 a_n5434_7417.n0 GND 0.694499f
C928 a_n5434_7417.t0 GND 90.1449f
C929 a_n5434_7417.t4 GND 0.025723f
C930 a_n5434_7417.t15 GND 0.178199f
C931 a_n5434_7417.t12 GND 0.025723f
C932 a_n5434_7417.t1 GND 0.025723f
C933 a_n5434_7417.n1 GND 0.112684f
C934 a_n5434_7417.n2 GND 0.749359f
C935 a_n5434_7417.t13 GND 0.169139f
C936 a_n5434_7417.n3 GND 0.781481f
C937 a_n5434_7417.n4 GND 2.41553f
C938 a_n5434_7417.t3 GND 0.1782f
C939 a_n5434_7417.t16 GND 0.025723f
C940 a_n5434_7417.t14 GND 0.025723f
C941 a_n5434_7417.n5 GND 0.112684f
C942 a_n5434_7417.n6 GND 0.749358f
C943 a_n5434_7417.t2 GND 0.169139f
C944 a_n5434_7417.n7 GND 1.27297f
C945 a_n5434_7417.n8 GND 1.36362f
C946 a_n5434_7417.t6 GND 0.169139f
C947 a_n5434_7417.n9 GND 0.497448f
C948 a_n5434_7417.t7 GND 0.025723f
C949 a_n5434_7417.t8 GND 0.025723f
C950 a_n5434_7417.n10 GND 0.112684f
C951 a_n5434_7417.n11 GND 0.444713f
C952 a_n5434_7417.t10 GND 0.169139f
C953 a_n5434_7417.t5 GND 0.169139f
C954 a_n5434_7417.t9 GND 0.1782f
C955 a_n5434_7417.n12 GND 0.749358f
C956 a_n5434_7417.n13 GND 0.112684f
C957 a_n5434_7417.t11 GND 0.025723f
C958 VP.t2 GND 1.43239f
C959 VP.t3 GND 1.74455f
C960 VP.n0 GND 2.12514f
C961 VP.t0 GND 0.030433f
C962 VP.t1 GND 0.030248f
C963 VP.n1 GND 0.144962f
C964 VP.n2 GND 1.50704f
C965 VDD.t99 GND 0.007261f
C966 VDD.t103 GND 0.007261f
C967 VDD.n0 GND 0.040736f
C968 VDD.t107 GND 0.007261f
C969 VDD.t113 GND 0.007261f
C970 VDD.n1 GND 0.037227f
C971 VDD.n2 GND 0.257805f
C972 VDD.t86 GND 0.007261f
C973 VDD.t117 GND 0.007261f
C974 VDD.n3 GND 0.037227f
C975 VDD.n4 GND 0.135391f
C976 VDD.t81 GND 0.007261f
C977 VDD.t109 GND 0.007261f
C978 VDD.n5 GND 0.037227f
C979 VDD.n6 GND 0.114936f
C980 VDD.t79 GND 0.007261f
C981 VDD.t115 GND 0.007261f
C982 VDD.n7 GND 0.040736f
C983 VDD.t84 GND 0.007261f
C984 VDD.t105 GND 0.007261f
C985 VDD.n8 GND 0.037227f
C986 VDD.n9 GND 0.257805f
C987 VDD.t92 GND 0.007261f
C988 VDD.t89 GND 0.007261f
C989 VDD.n10 GND 0.037227f
C990 VDD.n11 GND 0.135391f
C991 VDD.t111 GND 0.007261f
C992 VDD.t95 GND 0.007261f
C993 VDD.n12 GND 0.037227f
C994 VDD.n13 GND 0.114936f
C995 VDD.n14 GND 0.087519f
C996 VDD.n15 GND 2.83343f
C997 VDD.n16 GND 0.006445f
C998 VDD.n17 GND 0.006445f
C999 VDD.n18 GND 0.005205f
C1000 VDD.n19 GND 0.005205f
C1001 VDD.n20 GND 0.006467f
C1002 VDD.n21 GND 0.006467f
C1003 VDD.n22 GND 0.38361f
C1004 VDD.n23 GND 0.38361f
C1005 VDD.n24 GND 0.006467f
C1006 VDD.n25 GND 0.006467f
C1007 VDD.n26 GND 0.005205f
C1008 VDD.n27 GND 0.006467f
C1009 VDD.n28 GND 0.005205f
C1010 VDD.n29 GND 0.006467f
C1011 VDD.n30 GND 0.38361f
C1012 VDD.n31 GND 0.006467f
C1013 VDD.n32 GND 0.005205f
C1014 VDD.n33 GND 0.006467f
C1015 VDD.n34 GND 0.005205f
C1016 VDD.n35 GND 0.006467f
C1017 VDD.n36 GND 0.38361f
C1018 VDD.n37 GND 0.006467f
C1019 VDD.n38 GND 0.005205f
C1020 VDD.n39 GND 0.006467f
C1021 VDD.n40 GND 0.005205f
C1022 VDD.n41 GND 0.006467f
C1023 VDD.n42 GND 0.38361f
C1024 VDD.n43 GND 0.006467f
C1025 VDD.n44 GND 0.005205f
C1026 VDD.n45 GND 0.006467f
C1027 VDD.n46 GND 0.005205f
C1028 VDD.n47 GND 0.006467f
C1029 VDD.n48 GND 0.218658f
C1030 VDD.n49 GND 0.006467f
C1031 VDD.n50 GND 0.005205f
C1032 VDD.n51 GND 0.006467f
C1033 VDD.n52 GND 0.005205f
C1034 VDD.n53 GND 0.006467f
C1035 VDD.n54 GND 0.38361f
C1036 VDD.t8 GND 0.191805f
C1037 VDD.n55 GND 0.006467f
C1038 VDD.n56 GND 0.005205f
C1039 VDD.n57 GND 0.014445f
C1040 VDD.n58 GND 0.00432f
C1041 VDD.n59 GND 0.014445f
C1042 VDD.n60 GND 0.487185f
C1043 VDD.n61 GND 0.014445f
C1044 VDD.n62 GND 0.00432f
C1045 VDD.n63 GND 0.006467f
C1046 VDD.t27 GND 0.089332f
C1047 VDD.t28 GND 0.10348f
C1048 VDD.t26 GND 0.482813f
C1049 VDD.n64 GND 0.068834f
C1050 VDD.n65 GND 0.04271f
C1051 VDD.n66 GND 0.008016f
C1052 VDD.n67 GND 0.006467f
C1053 VDD.t75 GND 4.68772f
C1054 VDD.n87 GND 0.006467f
C1055 VDD.n88 GND 0.006467f
C1056 VDD.n89 GND 0.014463f
C1057 VDD.n90 GND 0.006467f
C1058 VDD.n91 GND 0.006467f
C1059 VDD.n92 GND 0.006467f
C1060 VDD.n93 GND 0.006467f
C1061 VDD.n94 GND 0.006338f
C1062 VDD.n97 GND 0.003363f
C1063 VDD.n98 GND 0.006467f
C1064 VDD.n99 GND 0.004346f
C1065 VDD.n100 GND 0.006467f
C1066 VDD.n101 GND 0.006467f
C1067 VDD.n102 GND 0.006467f
C1068 VDD.n103 GND 0.006467f
C1069 VDD.n104 GND 0.006467f
C1070 VDD.n105 GND 0.006467f
C1071 VDD.n106 GND 0.006467f
C1072 VDD.n107 GND 0.006467f
C1073 VDD.n108 GND 0.006467f
C1074 VDD.n109 GND 0.006467f
C1075 VDD.n110 GND 0.006467f
C1076 VDD.n111 GND 0.006467f
C1077 VDD.n112 GND 0.006467f
C1078 VDD.n113 GND 0.006467f
C1079 VDD.n114 GND 0.005153f
C1080 VDD.t24 GND 0.089332f
C1081 VDD.t25 GND 0.10348f
C1082 VDD.t23 GND 0.482813f
C1083 VDD.n115 GND 0.068834f
C1084 VDD.n116 GND 0.04271f
C1085 VDD.n117 GND 0.006467f
C1086 VDD.n118 GND 0.006467f
C1087 VDD.n119 GND 0.003363f
C1088 VDD.n120 GND 0.005205f
C1089 VDD.n121 GND 0.006338f
C1090 VDD.n122 GND 0.004398f
C1091 VDD.n123 GND 0.004398f
C1092 VDD.n124 GND 0.004398f
C1093 VDD.t114 GND 3.95502f
C1094 VDD.t78 GND 2.2633f
C1095 VDD.n125 GND 0.72886f
C1096 VDD.n126 GND 0.004398f
C1097 VDD.n127 GND 0.004398f
C1098 VDD.t54 GND 0.041419f
C1099 VDD.t53 GND 0.056208f
C1100 VDD.t52 GND 0.369485f
C1101 VDD.n128 GND 0.058137f
C1102 VDD.n129 GND 0.040639f
C1103 VDD.n130 GND 0.006285f
C1104 VDD.n132 GND 0.003686f
C1105 VDD.n133 GND 0.009619f
C1106 VDD.n134 GND 0.004398f
C1107 VDD.n135 GND 0.004398f
C1108 VDD.n136 GND 0.260855f
C1109 VDD.n137 GND 0.004398f
C1110 VDD.n138 GND 0.36443f
C1111 VDD.n139 GND 0.004398f
C1112 VDD.n140 GND 0.004398f
C1113 VDD.n141 GND 0.009619f
C1114 VDD.n142 GND 0.004398f
C1115 VDD.n143 GND 0.004398f
C1116 VDD.n144 GND 0.004398f
C1117 VDD.n145 GND 0.004398f
C1118 VDD.n147 GND 0.004398f
C1119 VDD.n148 GND 0.004398f
C1120 VDD.n150 GND 0.004398f
C1121 VDD.t6 GND 0.041419f
C1122 VDD.t5 GND 0.056208f
C1123 VDD.t3 GND 0.369485f
C1124 VDD.n151 GND 0.058137f
C1125 VDD.n152 GND 0.040639f
C1126 VDD.n153 GND 0.006285f
C1127 VDD.n155 GND 0.003686f
C1128 VDD.n156 GND 0.009619f
C1129 VDD.n157 GND 0.004398f
C1130 VDD.n158 GND 0.004398f
C1131 VDD.n159 GND 0.260855f
C1132 VDD.n160 GND 0.004398f
C1133 VDD.n161 GND 0.004398f
C1134 VDD.n162 GND 0.004398f
C1135 VDD.n163 GND 0.004398f
C1136 VDD.n164 GND 0.004398f
C1137 VDD.n165 GND 0.260855f
C1138 VDD.n166 GND 0.004398f
C1139 VDD.n167 GND 0.004398f
C1140 VDD.n168 GND 0.004398f
C1141 VDD.n169 GND 0.004398f
C1142 VDD.n170 GND 0.004398f
C1143 VDD.n171 GND 0.004398f
C1144 VDD.t4 GND 0.126591f
C1145 VDD.n172 GND 0.004398f
C1146 VDD.n173 GND 0.004398f
C1147 VDD.n174 GND 0.004398f
C1148 VDD.n175 GND 0.004398f
C1149 VDD.n176 GND 0.004398f
C1150 VDD.n177 GND 0.260855f
C1151 VDD.n178 GND 0.004398f
C1152 VDD.n179 GND 0.004398f
C1153 VDD.t104 GND 0.013426f
C1154 VDD.n180 GND 0.134264f
C1155 VDD.n181 GND 0.004398f
C1156 VDD.n182 GND 0.004398f
C1157 VDD.n183 GND 0.004398f
C1158 VDD.n184 GND 0.260855f
C1159 VDD.n185 GND 0.004398f
C1160 VDD.n186 GND 0.004398f
C1161 VDD.n187 GND 0.004398f
C1162 VDD.n188 GND 0.004398f
C1163 VDD.n189 GND 0.004398f
C1164 VDD.n190 GND 0.260855f
C1165 VDD.n191 GND 0.004398f
C1166 VDD.n192 GND 0.004398f
C1167 VDD.n193 GND 0.004398f
C1168 VDD.n194 GND 0.004398f
C1169 VDD.n195 GND 0.004398f
C1170 VDD.n196 GND 0.260855f
C1171 VDD.n197 GND 0.004398f
C1172 VDD.n198 GND 0.004398f
C1173 VDD.n199 GND 0.004398f
C1174 VDD.n200 GND 0.004398f
C1175 VDD.n201 GND 0.004398f
C1176 VDD.n202 GND 0.260855f
C1177 VDD.n203 GND 0.004398f
C1178 VDD.n204 GND 0.004398f
C1179 VDD.n205 GND 0.004398f
C1180 VDD.n206 GND 0.004398f
C1181 VDD.n207 GND 0.004398f
C1182 VDD.n208 GND 0.260855f
C1183 VDD.n209 GND 0.004398f
C1184 VDD.n210 GND 0.004398f
C1185 VDD.n211 GND 0.004398f
C1186 VDD.n212 GND 0.004398f
C1187 VDD.n213 GND 0.004398f
C1188 VDD.t83 GND 0.130428f
C1189 VDD.n214 GND 0.004398f
C1190 VDD.n215 GND 0.004398f
C1191 VDD.n216 GND 0.004398f
C1192 VDD.n217 GND 0.004398f
C1193 VDD.n218 GND 0.004398f
C1194 VDD.n219 GND 0.21674f
C1195 VDD.n220 GND 0.004398f
C1196 VDD.n221 GND 0.004398f
C1197 VDD.n222 GND 0.191805f
C1198 VDD.n223 GND 0.004398f
C1199 VDD.n224 GND 0.004398f
C1200 VDD.n225 GND 0.004398f
C1201 VDD.n226 GND 0.260855f
C1202 VDD.n227 GND 0.004398f
C1203 VDD.n228 GND 0.004398f
C1204 VDD.t87 GND 0.130428f
C1205 VDD.n229 GND 0.004398f
C1206 VDD.n230 GND 0.004398f
C1207 VDD.n231 GND 0.004398f
C1208 VDD.n232 GND 0.260855f
C1209 VDD.n233 GND 0.004398f
C1210 VDD.n234 GND 0.004398f
C1211 VDD.n235 GND 0.004398f
C1212 VDD.n236 GND 0.004398f
C1213 VDD.n237 GND 0.004398f
C1214 VDD.n238 GND 0.260855f
C1215 VDD.n239 GND 0.004398f
C1216 VDD.n240 GND 0.004398f
C1217 VDD.n241 GND 0.004398f
C1218 VDD.n242 GND 0.004398f
C1219 VDD.n243 GND 0.004398f
C1220 VDD.n244 GND 0.260855f
C1221 VDD.n245 GND 0.004398f
C1222 VDD.n246 GND 0.004398f
C1223 VDD.n247 GND 0.004398f
C1224 VDD.n248 GND 0.004398f
C1225 VDD.n249 GND 0.004398f
C1226 VDD.n250 GND 0.260855f
C1227 VDD.n251 GND 0.004398f
C1228 VDD.n252 GND 0.004398f
C1229 VDD.n253 GND 0.004398f
C1230 VDD.n254 GND 0.004398f
C1231 VDD.n255 GND 0.004398f
C1232 VDD.n256 GND 0.260855f
C1233 VDD.n257 GND 0.004398f
C1234 VDD.n258 GND 0.004398f
C1235 VDD.n259 GND 0.004398f
C1236 VDD.n260 GND 0.004398f
C1237 VDD.n261 GND 0.004398f
C1238 VDD.n262 GND 0.159198f
C1239 VDD.n263 GND 0.004398f
C1240 VDD.n264 GND 0.004398f
C1241 VDD.n265 GND 0.004398f
C1242 VDD.n266 GND 0.004398f
C1243 VDD.n267 GND 0.004398f
C1244 VDD.n268 GND 0.260855f
C1245 VDD.n269 GND 0.004398f
C1246 VDD.n270 GND 0.004398f
C1247 VDD.t90 GND 0.130428f
C1248 VDD.n271 GND 0.004398f
C1249 VDD.n272 GND 0.004398f
C1250 VDD.n273 GND 0.004398f
C1251 VDD.n274 GND 0.134264f
C1252 VDD.n275 GND 0.004398f
C1253 VDD.n276 GND 0.004398f
C1254 VDD.n277 GND 0.004398f
C1255 VDD.n278 GND 0.004398f
C1256 VDD.n279 GND 0.004398f
C1257 VDD.n280 GND 0.260855f
C1258 VDD.n281 GND 0.004398f
C1259 VDD.n282 GND 0.004398f
C1260 VDD.t88 GND 0.130428f
C1261 VDD.n283 GND 0.004398f
C1262 VDD.n284 GND 0.004398f
C1263 VDD.n285 GND 0.004398f
C1264 VDD.n286 GND 0.260855f
C1265 VDD.n287 GND 0.004398f
C1266 VDD.n288 GND 0.004398f
C1267 VDD.n289 GND 0.004398f
C1268 VDD.n290 GND 0.004398f
C1269 VDD.n291 GND 0.004398f
C1270 VDD.n292 GND 0.260855f
C1271 VDD.n293 GND 0.004398f
C1272 VDD.n294 GND 0.004398f
C1273 VDD.n295 GND 0.004398f
C1274 VDD.n296 GND 0.004398f
C1275 VDD.n297 GND 0.004398f
C1276 VDD.n298 GND 0.260855f
C1277 VDD.n299 GND 0.004398f
C1278 VDD.n300 GND 0.004398f
C1279 VDD.n301 GND 0.004398f
C1280 VDD.n302 GND 0.004398f
C1281 VDD.n303 GND 0.004398f
C1282 VDD.t93 GND 0.130428f
C1283 VDD.n304 GND 0.004398f
C1284 VDD.n305 GND 0.004398f
C1285 VDD.n306 GND 0.004398f
C1286 VDD.n307 GND 0.004398f
C1287 VDD.n308 GND 0.004398f
C1288 VDD.n309 GND 0.260855f
C1289 VDD.n310 GND 0.004398f
C1290 VDD.n311 GND 0.004398f
C1291 VDD.n312 GND 0.159198f
C1292 VDD.n313 GND 0.004398f
C1293 VDD.n314 GND 0.004398f
C1294 VDD.n315 GND 0.004398f
C1295 VDD.t91 GND 0.130428f
C1296 VDD.n316 GND 0.004398f
C1297 VDD.n317 GND 0.004398f
C1298 VDD.n318 GND 0.004398f
C1299 VDD.n319 GND 0.004398f
C1300 VDD.n320 GND 0.004398f
C1301 VDD.n321 GND 0.260855f
C1302 VDD.n322 GND 0.004398f
C1303 VDD.n323 GND 0.004398f
C1304 VDD.n324 GND 0.184133f
C1305 VDD.n325 GND 0.004398f
C1306 VDD.n326 GND 0.004398f
C1307 VDD.n327 GND 0.004398f
C1308 VDD.n328 GND 0.260855f
C1309 VDD.n329 GND 0.004398f
C1310 VDD.n330 GND 0.004398f
C1311 VDD.n331 GND 0.004398f
C1312 VDD.n332 GND 0.004398f
C1313 VDD.n333 GND 0.004398f
C1314 VDD.n334 GND 0.260855f
C1315 VDD.n335 GND 0.004398f
C1316 VDD.n336 GND 0.004398f
C1317 VDD.n337 GND 0.004398f
C1318 VDD.n338 GND 0.004398f
C1319 VDD.n339 GND 0.004398f
C1320 VDD.n340 GND 0.260855f
C1321 VDD.n341 GND 0.004398f
C1322 VDD.n342 GND 0.004398f
C1323 VDD.n343 GND 0.004398f
C1324 VDD.n344 GND 0.004398f
C1325 VDD.n345 GND 0.004398f
C1326 VDD.t96 GND 0.130428f
C1327 VDD.n346 GND 0.004398f
C1328 VDD.n347 GND 0.004398f
C1329 VDD.n348 GND 0.004398f
C1330 VDD.n349 GND 0.004398f
C1331 VDD.n350 GND 0.004398f
C1332 VDD.n351 GND 0.260855f
C1333 VDD.n352 GND 0.004398f
C1334 VDD.n353 GND 0.004398f
C1335 VDD.n354 GND 0.21674f
C1336 VDD.n355 GND 0.004398f
C1337 VDD.n356 GND 0.004398f
C1338 VDD.n357 GND 0.004398f
C1339 VDD.t94 GND 0.130428f
C1340 VDD.n358 GND 0.004398f
C1341 VDD.n359 GND 0.004398f
C1342 VDD.n360 GND 0.004398f
C1343 VDD.n361 GND 0.004398f
C1344 VDD.n362 GND 0.004398f
C1345 VDD.n363 GND 0.260855f
C1346 VDD.n364 GND 0.004398f
C1347 VDD.n365 GND 0.004398f
C1348 VDD.n366 GND 0.241675f
C1349 VDD.n367 GND 0.004398f
C1350 VDD.n368 GND 0.004398f
C1351 VDD.n369 GND 0.004398f
C1352 VDD.n370 GND 0.260855f
C1353 VDD.n371 GND 0.004398f
C1354 VDD.n372 GND 0.004398f
C1355 VDD.n373 GND 0.004398f
C1356 VDD.n374 GND 0.004398f
C1357 VDD.n375 GND 0.004398f
C1358 VDD.n376 GND 0.260855f
C1359 VDD.n377 GND 0.004398f
C1360 VDD.n378 GND 0.004398f
C1361 VDD.n379 GND 0.004398f
C1362 VDD.n380 GND 0.004398f
C1363 VDD.n381 GND 0.004398f
C1364 VDD.n382 GND 0.260855f
C1365 VDD.n383 GND 0.004398f
C1366 VDD.n384 GND 0.004398f
C1367 VDD.n385 GND 0.004398f
C1368 VDD.n386 GND 0.004398f
C1369 VDD.n387 GND 0.004398f
C1370 VDD.n388 GND 0.260855f
C1371 VDD.n389 GND 0.004398f
C1372 VDD.n390 GND 0.004398f
C1373 VDD.n391 GND 0.004398f
C1374 VDD.n392 GND 0.004398f
C1375 VDD.n393 GND 0.004398f
C1376 VDD.n394 GND 0.143854f
C1377 VDD.n395 GND 0.004398f
C1378 VDD.n396 GND 0.004398f
C1379 VDD.n397 GND 0.004398f
C1380 VDD.n398 GND 0.004398f
C1381 VDD.n399 GND 0.004398f
C1382 VDD.n400 GND 0.260855f
C1383 VDD.n401 GND 0.004398f
C1384 VDD.n402 GND 0.004398f
C1385 VDD.t59 GND 0.092066f
C1386 VDD.t110 GND 0.117001f
C1387 VDD.n403 GND 0.004398f
C1388 VDD.n404 GND 0.004398f
C1389 VDD.n405 GND 0.004398f
C1390 VDD.n406 GND 0.260855f
C1391 VDD.n407 GND 0.004398f
C1392 VDD.n408 GND 0.004398f
C1393 VDD.n409 GND 0.004398f
C1394 VDD.n410 GND 0.004398f
C1395 VDD.n411 GND 0.004398f
C1396 VDD.n412 GND 0.260855f
C1397 VDD.n413 GND 0.004398f
C1398 VDD.n414 GND 0.004398f
C1399 VDD.n415 GND 0.004398f
C1400 VDD.n416 GND 0.009619f
C1401 VDD.n417 GND 0.009619f
C1402 VDD.n418 GND 0.36443f
C1403 VDD.n419 GND 0.004398f
C1404 VDD.n420 GND 0.004398f
C1405 VDD.n421 GND 0.009619f
C1406 VDD.n422 GND 0.004398f
C1407 VDD.n423 GND 0.004398f
C1408 VDD.n424 GND 0.36443f
C1409 VDD.n432 GND 0.010235f
C1410 VDD.n440 GND 0.009619f
C1411 VDD.n441 GND 0.004398f
C1412 VDD.n442 GND 0.009619f
C1413 VDD.t51 GND 0.041419f
C1414 VDD.t50 GND 0.056208f
C1415 VDD.t48 GND 0.369485f
C1416 VDD.n443 GND 0.058137f
C1417 VDD.n444 GND 0.040639f
C1418 VDD.n445 GND 0.006285f
C1419 VDD.n446 GND 0.010168f
C1420 VDD.n447 GND 0.004398f
C1421 VDD.n448 GND 0.004398f
C1422 VDD.n449 GND 0.260855f
C1423 VDD.n450 GND 0.004398f
C1424 VDD.n451 GND 0.004398f
C1425 VDD.n452 GND 0.004398f
C1426 VDD.n453 GND 0.004398f
C1427 VDD.n454 GND 0.004398f
C1428 VDD.n455 GND 0.260855f
C1429 VDD.n456 GND 0.004398f
C1430 VDD.n457 GND 0.004398f
C1431 VDD.n458 GND 0.004398f
C1432 VDD.n459 GND 0.004398f
C1433 VDD.n460 GND 0.004398f
C1434 VDD.t57 GND 0.041419f
C1435 VDD.t56 GND 0.056208f
C1436 VDD.t55 GND 0.369485f
C1437 VDD.n461 GND 0.058137f
C1438 VDD.n462 GND 0.040639f
C1439 VDD.n463 GND 0.004398f
C1440 VDD.n464 GND 0.004398f
C1441 VDD.n465 GND 0.260855f
C1442 VDD.n466 GND 0.004398f
C1443 VDD.n467 GND 0.004398f
C1444 VDD.n468 GND 0.004398f
C1445 VDD.n469 GND 0.004398f
C1446 VDD.n470 GND 0.004398f
C1447 VDD.t108 GND 0.117001f
C1448 VDD.n471 GND 0.004398f
C1449 VDD.n472 GND 0.004398f
C1450 VDD.n473 GND 0.004398f
C1451 VDD.n474 GND 0.004398f
C1452 VDD.n475 GND 0.004398f
C1453 VDD.n476 GND 0.004398f
C1454 VDD.n477 GND 0.260855f
C1455 VDD.n478 GND 0.004398f
C1456 VDD.n479 GND 0.004398f
C1457 VDD.t49 GND 0.092066f
C1458 VDD.n480 GND 0.143854f
C1459 VDD.n481 GND 0.004398f
C1460 VDD.n482 GND 0.004398f
C1461 VDD.n483 GND 0.004398f
C1462 VDD.n484 GND 0.260855f
C1463 VDD.n485 GND 0.004398f
C1464 VDD.n486 GND 0.004398f
C1465 VDD.n487 GND 0.004398f
C1466 VDD.n488 GND 0.004398f
C1467 VDD.n489 GND 0.004398f
C1468 VDD.n490 GND 0.260855f
C1469 VDD.n491 GND 0.004398f
C1470 VDD.n492 GND 0.004398f
C1471 VDD.n493 GND 0.004398f
C1472 VDD.n494 GND 0.004398f
C1473 VDD.n495 GND 0.004398f
C1474 VDD.n496 GND 0.260855f
C1475 VDD.n497 GND 0.004398f
C1476 VDD.n498 GND 0.004398f
C1477 VDD.n499 GND 0.004398f
C1478 VDD.n500 GND 0.004398f
C1479 VDD.n501 GND 0.004398f
C1480 VDD.n502 GND 0.260855f
C1481 VDD.n503 GND 0.004398f
C1482 VDD.n504 GND 0.004398f
C1483 VDD.n505 GND 0.004398f
C1484 VDD.n506 GND 0.004398f
C1485 VDD.n507 GND 0.004398f
C1486 VDD.n508 GND 0.241675f
C1487 VDD.n509 GND 0.004398f
C1488 VDD.n510 GND 0.004398f
C1489 VDD.n511 GND 0.004398f
C1490 VDD.n512 GND 0.004398f
C1491 VDD.n513 GND 0.004398f
C1492 VDD.n514 GND 0.260855f
C1493 VDD.n515 GND 0.004398f
C1494 VDD.n516 GND 0.004398f
C1495 VDD.t80 GND 0.130428f
C1496 VDD.n517 GND 0.004398f
C1497 VDD.n518 GND 0.004398f
C1498 VDD.n519 GND 0.004398f
C1499 VDD.n520 GND 0.21674f
C1500 VDD.n521 GND 0.004398f
C1501 VDD.n522 GND 0.004398f
C1502 VDD.n523 GND 0.004398f
C1503 VDD.n524 GND 0.004398f
C1504 VDD.n525 GND 0.004398f
C1505 VDD.n526 GND 0.260855f
C1506 VDD.n527 GND 0.004398f
C1507 VDD.n528 GND 0.004398f
C1508 VDD.t82 GND 0.130428f
C1509 VDD.n529 GND 0.004398f
C1510 VDD.n530 GND 0.004398f
C1511 VDD.n531 GND 0.004398f
C1512 VDD.n532 GND 0.260855f
C1513 VDD.n533 GND 0.004398f
C1514 VDD.n534 GND 0.004398f
C1515 VDD.n535 GND 0.004398f
C1516 VDD.n536 GND 0.004398f
C1517 VDD.n537 GND 0.004398f
C1518 VDD.n538 GND 0.260855f
C1519 VDD.n539 GND 0.004398f
C1520 VDD.n540 GND 0.004398f
C1521 VDD.n541 GND 0.004398f
C1522 VDD.n542 GND 0.004398f
C1523 VDD.n543 GND 0.004398f
C1524 VDD.n544 GND 0.260855f
C1525 VDD.n545 GND 0.004398f
C1526 VDD.n546 GND 0.004398f
C1527 VDD.n547 GND 0.004398f
C1528 VDD.n548 GND 0.004398f
C1529 VDD.n549 GND 0.004398f
C1530 VDD.n550 GND 0.184133f
C1531 VDD.n551 GND 0.004398f
C1532 VDD.n552 GND 0.004398f
C1533 VDD.n553 GND 0.004398f
C1534 VDD.n554 GND 0.004398f
C1535 VDD.n555 GND 0.004398f
C1536 VDD.n556 GND 0.260855f
C1537 VDD.n557 GND 0.004398f
C1538 VDD.n558 GND 0.004398f
C1539 VDD.t116 GND 0.130428f
C1540 VDD.n559 GND 0.004398f
C1541 VDD.n560 GND 0.004398f
C1542 VDD.n561 GND 0.004398f
C1543 VDD.n562 GND 0.159198f
C1544 VDD.n563 GND 0.004398f
C1545 VDD.n564 GND 0.004398f
C1546 VDD.n565 GND 0.004398f
C1547 VDD.n566 GND 0.004398f
C1548 VDD.n567 GND 0.004398f
C1549 VDD.n568 GND 0.260855f
C1550 VDD.n569 GND 0.004398f
C1551 VDD.n570 GND 0.004398f
C1552 VDD.t100 GND 0.130428f
C1553 VDD.n571 GND 0.004398f
C1554 VDD.n572 GND 0.004398f
C1555 VDD.n573 GND 0.004398f
C1556 VDD.n574 GND 0.260855f
C1557 VDD.n575 GND 0.004398f
C1558 VDD.n576 GND 0.004398f
C1559 VDD.n577 GND 0.004398f
C1560 VDD.n578 GND 0.004398f
C1561 VDD.n579 GND 0.004398f
C1562 VDD.n580 GND 0.260855f
C1563 VDD.n581 GND 0.004398f
C1564 VDD.n582 GND 0.004398f
C1565 VDD.n583 GND 0.004398f
C1566 VDD.n584 GND 0.004398f
C1567 VDD.n585 GND 0.004398f
C1568 VDD.n586 GND 0.260855f
C1569 VDD.n587 GND 0.004398f
C1570 VDD.n588 GND 0.004398f
C1571 VDD.n589 GND 0.004398f
C1572 VDD.n590 GND 0.004398f
C1573 VDD.n591 GND 0.004398f
C1574 VDD.t85 GND 0.130428f
C1575 VDD.n592 GND 0.004398f
C1576 VDD.n593 GND 0.004398f
C1577 VDD.n594 GND 0.004398f
C1578 VDD.n595 GND 0.004398f
C1579 VDD.n596 GND 0.004398f
C1580 VDD.n597 GND 0.260855f
C1581 VDD.n598 GND 0.004398f
C1582 VDD.n599 GND 0.004398f
C1583 VDD.n600 GND 0.134264f
C1584 VDD.n601 GND 0.004398f
C1585 VDD.n602 GND 0.004398f
C1586 VDD.n603 GND 0.004398f
C1587 VDD.t101 GND 0.130428f
C1588 VDD.n604 GND 0.004398f
C1589 VDD.n605 GND 0.004398f
C1590 VDD.n606 GND 0.004398f
C1591 VDD.n607 GND 0.004398f
C1592 VDD.n608 GND 0.004398f
C1593 VDD.n609 GND 0.260855f
C1594 VDD.n610 GND 0.004398f
C1595 VDD.n611 GND 0.004398f
C1596 VDD.n612 GND 0.159198f
C1597 VDD.n613 GND 0.004398f
C1598 VDD.n614 GND 0.004398f
C1599 VDD.n615 GND 0.004398f
C1600 VDD.n616 GND 0.260855f
C1601 VDD.n617 GND 0.004398f
C1602 VDD.n618 GND 0.004398f
C1603 VDD.n619 GND 0.004398f
C1604 VDD.n620 GND 0.004398f
C1605 VDD.n621 GND 0.004398f
C1606 VDD.n622 GND 0.260855f
C1607 VDD.n623 GND 0.004398f
C1608 VDD.n624 GND 0.004398f
C1609 VDD.n625 GND 0.004398f
C1610 VDD.n626 GND 0.004398f
C1611 VDD.n627 GND 0.004398f
C1612 VDD.n628 GND 0.260855f
C1613 VDD.n629 GND 0.004398f
C1614 VDD.n630 GND 0.004398f
C1615 VDD.n631 GND 0.004398f
C1616 VDD.n632 GND 0.004398f
C1617 VDD.n633 GND 0.004398f
C1618 VDD.n634 GND 0.260855f
C1619 VDD.n635 GND 0.004398f
C1620 VDD.n636 GND 0.004398f
C1621 VDD.n637 GND 0.004398f
C1622 VDD.n638 GND 0.004398f
C1623 VDD.n639 GND 0.004398f
C1624 VDD.n640 GND 0.260855f
C1625 VDD.n641 GND 0.004398f
C1626 VDD.n642 GND 0.004398f
C1627 VDD.n643 GND 0.004398f
C1628 VDD.n644 GND 0.004398f
C1629 VDD.n645 GND 0.004398f
C1630 VDD.t97 GND 0.130428f
C1631 VDD.n646 GND 0.004398f
C1632 VDD.n647 GND 0.004398f
C1633 VDD.n648 GND 0.004398f
C1634 VDD.n649 GND 0.004398f
C1635 VDD.n650 GND 0.004398f
C1636 VDD.n651 GND 0.191805f
C1637 VDD.n652 GND 0.004398f
C1638 VDD.n653 GND 0.004398f
C1639 VDD.n654 GND 0.21674f
C1640 VDD.n655 GND 0.004398f
C1641 VDD.n656 GND 0.004398f
C1642 VDD.n657 GND 0.004398f
C1643 VDD.n658 GND 0.260855f
C1644 VDD.n659 GND 0.004398f
C1645 VDD.n660 GND 0.004398f
C1646 VDD.t112 GND 0.130428f
C1647 VDD.n661 GND 0.004398f
C1648 VDD.n662 GND 0.004398f
C1649 VDD.n663 GND 0.004398f
C1650 VDD.n664 GND 0.260855f
C1651 VDD.n665 GND 0.004398f
C1652 VDD.n666 GND 0.004398f
C1653 VDD.n667 GND 0.004398f
C1654 VDD.n668 GND 0.004398f
C1655 VDD.n669 GND 0.004398f
C1656 VDD.n670 GND 0.260855f
C1657 VDD.n671 GND 0.004398f
C1658 VDD.n672 GND 0.004398f
C1659 VDD.n673 GND 0.004398f
C1660 VDD.n674 GND 0.004398f
C1661 VDD.n675 GND 0.004398f
C1662 VDD.n676 GND 0.260855f
C1663 VDD.n677 GND 0.004398f
C1664 VDD.n678 GND 0.004398f
C1665 VDD.n679 GND 0.004398f
C1666 VDD.n680 GND 0.004398f
C1667 VDD.n681 GND 0.004398f
C1668 VDD.n682 GND 0.260855f
C1669 VDD.n683 GND 0.004398f
C1670 VDD.n684 GND 0.004398f
C1671 VDD.n685 GND 0.004398f
C1672 VDD.n686 GND 0.004398f
C1673 VDD.n687 GND 0.004398f
C1674 VDD.n688 GND 0.260855f
C1675 VDD.n689 GND 0.004398f
C1676 VDD.n690 GND 0.004398f
C1677 VDD.n691 GND 0.004398f
C1678 VDD.n692 GND 0.004398f
C1679 VDD.n693 GND 0.004398f
C1680 VDD.n694 GND 0.134264f
C1681 VDD.n695 GND 0.004398f
C1682 VDD.n696 GND 0.004398f
C1683 VDD.n697 GND 0.004398f
C1684 VDD.n698 GND 0.004398f
C1685 VDD.n699 GND 0.004398f
C1686 VDD.n700 GND 0.260855f
C1687 VDD.n701 GND 0.004398f
C1688 VDD.n702 GND 0.004398f
C1689 VDD.t106 GND 0.013426f
C1690 VDD.t20 GND 0.126591f
C1691 VDD.n703 GND 0.004398f
C1692 VDD.n704 GND 0.004398f
C1693 VDD.n705 GND 0.004398f
C1694 VDD.n706 GND 0.260855f
C1695 VDD.n707 GND 0.004398f
C1696 VDD.n708 GND 0.004398f
C1697 VDD.n709 GND 0.004398f
C1698 VDD.n710 GND 0.004398f
C1699 VDD.n711 GND 0.004398f
C1700 VDD.n712 GND 0.260855f
C1701 VDD.n713 GND 0.004398f
C1702 VDD.n714 GND 0.004398f
C1703 VDD.n715 GND 0.004398f
C1704 VDD.n716 GND 0.009619f
C1705 VDD.n717 GND 0.009619f
C1706 VDD.n718 GND 0.36443f
C1707 VDD.n719 GND 0.004398f
C1708 VDD.n720 GND 0.004398f
C1709 VDD.n721 GND 0.009619f
C1710 VDD.n722 GND 0.004398f
C1711 VDD.n723 GND 0.004398f
C1712 VDD.t102 GND 2.2633f
C1713 VDD.n737 GND 0.010235f
C1714 VDD.n738 GND 0.004398f
C1715 VDD.n739 GND 0.006338f
C1716 VDD.n740 GND 0.003363f
C1717 VDD.n742 GND 0.005205f
C1718 VDD.n743 GND 0.005205f
C1719 VDD.t98 GND 3.95502f
C1720 VDD.t71 GND 4.68772f
C1721 VDD.n745 GND 2.79652f
C1722 VDD.n746 GND 0.005205f
C1723 VDD.n747 GND 0.006467f
C1724 VDD.n748 GND 0.006467f
C1725 VDD.n749 GND 0.004346f
C1726 VDD.t18 GND 0.089332f
C1727 VDD.t17 GND 0.10348f
C1728 VDD.t15 GND 0.482813f
C1729 VDD.n750 GND 0.068834f
C1730 VDD.n751 GND 0.04271f
C1731 VDD.n753 GND 0.006467f
C1732 VDD.n754 GND 0.006467f
C1733 VDD.n755 GND 0.005205f
C1734 VDD.n756 GND 0.006467f
C1735 VDD.n758 GND 0.006467f
C1736 VDD.n759 GND 0.006467f
C1737 VDD.n760 GND 0.006467f
C1738 VDD.n761 GND 0.006467f
C1739 VDD.n762 GND 0.005205f
C1740 VDD.n764 GND 0.006467f
C1741 VDD.n765 GND 0.006467f
C1742 VDD.n766 GND 0.006467f
C1743 VDD.n767 GND 0.006467f
C1744 VDD.n768 GND 0.006467f
C1745 VDD.n769 GND 0.005205f
C1746 VDD.n771 GND 0.006467f
C1747 VDD.n772 GND 0.006467f
C1748 VDD.n773 GND 0.006467f
C1749 VDD.n774 GND 0.006467f
C1750 VDD.n775 GND 0.006467f
C1751 VDD.t43 GND 0.089332f
C1752 VDD.t42 GND 0.10348f
C1753 VDD.t41 GND 0.482813f
C1754 VDD.n776 GND 0.068834f
C1755 VDD.n777 GND 0.04271f
C1756 VDD.n778 GND 0.010619f
C1757 VDD.n780 GND 0.006467f
C1758 VDD.n781 GND 0.006467f
C1759 VDD.n782 GND 0.006467f
C1760 VDD.n783 GND 0.006467f
C1761 VDD.n784 GND 0.006467f
C1762 VDD.n785 GND 0.005205f
C1763 VDD.n787 GND 0.006467f
C1764 VDD.n788 GND 0.006467f
C1765 VDD.n789 GND 0.003363f
C1766 VDD.n790 GND 0.005205f
C1767 VDD.n791 GND 0.010235f
C1768 VDD.n792 GND 0.010235f
C1769 VDD.n793 GND 0.004398f
C1770 VDD.n794 GND 0.004398f
C1771 VDD.n795 GND 0.004398f
C1772 VDD.n796 GND 0.004398f
C1773 VDD.n797 GND 0.004398f
C1774 VDD.n798 GND 0.004398f
C1775 VDD.n799 GND 0.004398f
C1776 VDD.n800 GND 0.004398f
C1777 VDD.n801 GND 0.004398f
C1778 VDD.n802 GND 0.004398f
C1779 VDD.n803 GND 0.004398f
C1780 VDD.n804 GND 0.004398f
C1781 VDD.n805 GND 0.004398f
C1782 VDD.t21 GND 0.041419f
C1783 VDD.t22 GND 0.056208f
C1784 VDD.t19 GND 0.369485f
C1785 VDD.n806 GND 0.058137f
C1786 VDD.n807 GND 0.040639f
C1787 VDD.n808 GND 0.004398f
C1788 VDD.n809 GND 0.004398f
C1789 VDD.n810 GND 0.004398f
C1790 VDD.n811 GND 0.004398f
C1791 VDD.n812 GND 0.004398f
C1792 VDD.n813 GND 0.004398f
C1793 VDD.n814 GND 0.004398f
C1794 VDD.n815 GND 0.004398f
C1795 VDD.n816 GND 0.004398f
C1796 VDD.n817 GND 0.004398f
C1797 VDD.n818 GND 0.004398f
C1798 VDD.n819 GND 0.004398f
C1799 VDD.n820 GND 0.004398f
C1800 VDD.n821 GND 0.004398f
C1801 VDD.n822 GND 0.004398f
C1802 VDD.n823 GND 0.004398f
C1803 VDD.n824 GND 0.004398f
C1804 VDD.n825 GND 0.004398f
C1805 VDD.n826 GND 0.004398f
C1806 VDD.n827 GND 0.004398f
C1807 VDD.n828 GND 0.004398f
C1808 VDD.n829 GND 0.004398f
C1809 VDD.n830 GND 0.004398f
C1810 VDD.n831 GND 0.004398f
C1811 VDD.n832 GND 0.004398f
C1812 VDD.n833 GND 0.004398f
C1813 VDD.n834 GND 0.004398f
C1814 VDD.n835 GND 0.004398f
C1815 VDD.n836 GND 0.004398f
C1816 VDD.n837 GND 0.004398f
C1817 VDD.n838 GND 0.004398f
C1818 VDD.n839 GND 0.004398f
C1819 VDD.n840 GND 0.004398f
C1820 VDD.n841 GND 0.004398f
C1821 VDD.n842 GND 0.004398f
C1822 VDD.n843 GND 0.004398f
C1823 VDD.n844 GND 0.004398f
C1824 VDD.n845 GND 0.004398f
C1825 VDD.n846 GND 0.004398f
C1826 VDD.n847 GND 0.004398f
C1827 VDD.n848 GND 0.004398f
C1828 VDD.n849 GND 0.004398f
C1829 VDD.n850 GND 0.004398f
C1830 VDD.n851 GND 0.004398f
C1831 VDD.n852 GND 0.004398f
C1832 VDD.n853 GND 0.004398f
C1833 VDD.n854 GND 0.004398f
C1834 VDD.n855 GND 0.004398f
C1835 VDD.n856 GND 0.004398f
C1836 VDD.n857 GND 0.004398f
C1837 VDD.n858 GND 0.004398f
C1838 VDD.n859 GND 0.004398f
C1839 VDD.n860 GND 0.004398f
C1840 VDD.n861 GND 0.004398f
C1841 VDD.n862 GND 0.004398f
C1842 VDD.n863 GND 0.004398f
C1843 VDD.n864 GND 0.004398f
C1844 VDD.n865 GND 0.004398f
C1845 VDD.n866 GND 0.004398f
C1846 VDD.n867 GND 0.004398f
C1847 VDD.n868 GND 0.004398f
C1848 VDD.n869 GND 0.004398f
C1849 VDD.n870 GND 0.004398f
C1850 VDD.n871 GND 0.004398f
C1851 VDD.n872 GND 0.004398f
C1852 VDD.n873 GND 0.004398f
C1853 VDD.n874 GND 0.004398f
C1854 VDD.n875 GND 0.004398f
C1855 VDD.n876 GND 0.004398f
C1856 VDD.n877 GND 0.004398f
C1857 VDD.n878 GND 0.004398f
C1858 VDD.n879 GND 0.004398f
C1859 VDD.n880 GND 0.004398f
C1860 VDD.n881 GND 0.004398f
C1861 VDD.n882 GND 0.004398f
C1862 VDD.n883 GND 0.004398f
C1863 VDD.n884 GND 0.004398f
C1864 VDD.n885 GND 0.004398f
C1865 VDD.n886 GND 0.004398f
C1866 VDD.n887 GND 0.004398f
C1867 VDD.n888 GND 0.004398f
C1868 VDD.n889 GND 0.004398f
C1869 VDD.n890 GND 0.004398f
C1870 VDD.n891 GND 0.004398f
C1871 VDD.n892 GND 0.004398f
C1872 VDD.n893 GND 0.004398f
C1873 VDD.n894 GND 0.004398f
C1874 VDD.n895 GND 0.004398f
C1875 VDD.n896 GND 0.004398f
C1876 VDD.n897 GND 0.004398f
C1877 VDD.n898 GND 0.004398f
C1878 VDD.n899 GND 0.004398f
C1879 VDD.n900 GND 0.004398f
C1880 VDD.n901 GND 0.004398f
C1881 VDD.n902 GND 0.004398f
C1882 VDD.n903 GND 0.004398f
C1883 VDD.n904 GND 0.004398f
C1884 VDD.n905 GND 0.004398f
C1885 VDD.n906 GND 0.004398f
C1886 VDD.n907 GND 0.004398f
C1887 VDD.n908 GND 0.004398f
C1888 VDD.n909 GND 0.004398f
C1889 VDD.n910 GND 0.004398f
C1890 VDD.n911 GND 0.004398f
C1891 VDD.n912 GND 0.004398f
C1892 VDD.n913 GND 0.004398f
C1893 VDD.n914 GND 0.004398f
C1894 VDD.n915 GND 0.004398f
C1895 VDD.n916 GND 0.004398f
C1896 VDD.n917 GND 0.004398f
C1897 VDD.n918 GND 0.004398f
C1898 VDD.n919 GND 0.004398f
C1899 VDD.n920 GND 0.004398f
C1900 VDD.n921 GND 0.004398f
C1901 VDD.n922 GND 0.004398f
C1902 VDD.n923 GND 0.004398f
C1903 VDD.n924 GND 0.004398f
C1904 VDD.n925 GND 0.004398f
C1905 VDD.n926 GND 0.004398f
C1906 VDD.n927 GND 0.004398f
C1907 VDD.n928 GND 0.004398f
C1908 VDD.n929 GND 0.004398f
C1909 VDD.n930 GND 0.004398f
C1910 VDD.n931 GND 0.004398f
C1911 VDD.n932 GND 0.004398f
C1912 VDD.n933 GND 0.009619f
C1913 VDD.n934 GND 0.009619f
C1914 VDD.n935 GND 0.010235f
C1915 VDD.n936 GND 0.004398f
C1916 VDD.n937 GND 0.003686f
C1917 VDD.n938 GND 0.006285f
C1918 VDD.n939 GND 0.00291f
C1919 VDD.n940 GND 0.004398f
C1920 VDD.n941 GND 0.004398f
C1921 VDD.n942 GND 0.004398f
C1922 VDD.n943 GND 0.004398f
C1923 VDD.n944 GND 0.004398f
C1924 VDD.n945 GND 0.004398f
C1925 VDD.n946 GND 0.004398f
C1926 VDD.n947 GND 0.004398f
C1927 VDD.n948 GND 0.004398f
C1928 VDD.n949 GND 0.066313f
C1929 VDD.n951 GND 0.006467f
C1930 VDD.n952 GND 0.005205f
C1931 VDD.n954 GND 0.006467f
C1932 VDD.n955 GND 0.005205f
C1933 VDD.n956 GND 0.006467f
C1934 VDD.n958 GND 0.006467f
C1935 VDD.n959 GND 0.006467f
C1936 VDD.n961 GND 0.006467f
C1937 VDD.n962 GND 0.006467f
C1938 VDD.n963 GND 0.005205f
C1939 VDD.n964 GND 0.014463f
C1940 VDD.n966 GND 0.006467f
C1941 VDD.n967 GND 0.006467f
C1942 VDD.n969 GND 0.006467f
C1943 VDD.n970 GND 0.00432f
C1944 VDD.n971 GND 0.38361f
C1945 VDD.n972 GND 0.006467f
C1946 VDD.n973 GND 0.014463f
C1947 VDD.n974 GND 0.005205f
C1948 VDD.n975 GND 0.006467f
C1949 VDD.n976 GND 0.005205f
C1950 VDD.n977 GND 0.006467f
C1951 VDD.n978 GND 0.356758f
C1952 VDD.n979 GND 0.006467f
C1953 VDD.n980 GND 0.005205f
C1954 VDD.n981 GND 0.005205f
C1955 VDD.n982 GND 0.006467f
C1956 VDD.n983 GND 0.005205f
C1957 VDD.n984 GND 0.006467f
C1958 VDD.n985 GND 0.38361f
C1959 VDD.t16 GND 0.191805f
C1960 VDD.n986 GND 0.006467f
C1961 VDD.n987 GND 0.005205f
C1962 VDD.n988 GND 0.006467f
C1963 VDD.n989 GND 0.005205f
C1964 VDD.n990 GND 0.006467f
C1965 VDD.n991 GND 0.38361f
C1966 VDD.n992 GND 0.006467f
C1967 VDD.n993 GND 0.005205f
C1968 VDD.n994 GND 0.006467f
C1969 VDD.n995 GND 0.005205f
C1970 VDD.n996 GND 0.006467f
C1971 VDD.n997 GND 0.38361f
C1972 VDD.n998 GND 0.006467f
C1973 VDD.n999 GND 0.005205f
C1974 VDD.n1000 GND 0.006467f
C1975 VDD.n1001 GND 0.005205f
C1976 VDD.n1002 GND 0.006467f
C1977 VDD.n1003 GND 0.38361f
C1978 VDD.n1004 GND 0.006467f
C1979 VDD.n1005 GND 0.005205f
C1980 VDD.n1006 GND 0.006467f
C1981 VDD.n1007 GND 0.005205f
C1982 VDD.n1008 GND 0.006467f
C1983 VDD.t72 GND 0.38361f
C1984 VDD.n1009 GND 0.006467f
C1985 VDD.n1010 GND 0.005205f
C1986 VDD.n1011 GND 0.006467f
C1987 VDD.n1012 GND 0.005205f
C1988 VDD.n1013 GND 0.006467f
C1989 VDD.n1014 GND 0.38361f
C1990 VDD.n1015 GND 0.006467f
C1991 VDD.n1016 GND 0.005205f
C1992 VDD.n1017 GND 0.006467f
C1993 VDD.n1018 GND 0.005205f
C1994 VDD.n1019 GND 0.006467f
C1995 VDD.n1020 GND 0.38361f
C1996 VDD.n1021 GND 0.006467f
C1997 VDD.n1022 GND 0.005205f
C1998 VDD.n1023 GND 0.006467f
C1999 VDD.n1024 GND 0.005205f
C2000 VDD.n1025 GND 0.006467f
C2001 VDD.n1026 GND 0.38361f
C2002 VDD.n1027 GND 0.006467f
C2003 VDD.n1028 GND 0.005205f
C2004 VDD.n1029 GND 0.006467f
C2005 VDD.n1030 GND 0.005205f
C2006 VDD.n1031 GND 0.006467f
C2007 VDD.n1032 GND 0.38361f
C2008 VDD.n1033 GND 0.006467f
C2009 VDD.n1034 GND 0.005205f
C2010 VDD.n1035 GND 0.006467f
C2011 VDD.n1036 GND 0.005205f
C2012 VDD.n1037 GND 0.006467f
C2013 VDD.t45 GND 0.191805f
C2014 VDD.n1038 GND 0.006467f
C2015 VDD.n1039 GND 0.005205f
C2016 VDD.n1040 GND 0.006467f
C2017 VDD.n1041 GND 0.005205f
C2018 VDD.n1042 GND 0.006467f
C2019 VDD.n1043 GND 0.38361f
C2020 VDD.n1044 GND 0.356758f
C2021 VDD.n1045 GND 0.006467f
C2022 VDD.n1046 GND 0.005205f
C2023 VDD.n1047 GND 0.014463f
C2024 VDD.n1048 GND 0.014463f
C2025 VDD.n1049 GND 0.836271f
C2026 VDD.n1050 GND 0.014463f
C2027 VDD.n1051 GND 0.006467f
C2028 VDD.t66 GND 0.089332f
C2029 VDD.t67 GND 0.10348f
C2030 VDD.t65 GND 0.482813f
C2031 VDD.n1052 GND 0.068834f
C2032 VDD.n1053 GND 0.04271f
C2033 VDD.n1054 GND 0.005205f
C2034 VDD.n1055 GND 0.006467f
C2035 VDD.n1056 GND 0.005205f
C2036 VDD.n1057 GND 0.006467f
C2037 VDD.n1058 GND 0.005205f
C2038 VDD.n1059 GND 0.006467f
C2039 VDD.n1060 GND 0.005205f
C2040 VDD.n1061 GND 0.006467f
C2041 VDD.n1062 GND 0.005205f
C2042 VDD.n1063 GND 0.006467f
C2043 VDD.n1064 GND 0.005205f
C2044 VDD.n1065 GND 0.006467f
C2045 VDD.n1066 GND 0.005153f
C2046 VDD.n1067 GND 0.006467f
C2047 VDD.n1068 GND 0.006467f
C2048 VDD.t69 GND 0.089332f
C2049 VDD.t70 GND 0.10348f
C2050 VDD.t68 GND 0.482813f
C2051 VDD.n1069 GND 0.068834f
C2052 VDD.n1070 GND 0.04271f
C2053 VDD.n1071 GND 0.005205f
C2054 VDD.n1072 GND 0.006467f
C2055 VDD.n1073 GND 0.005205f
C2056 VDD.n1075 GND 0.006467f
C2057 VDD.n1076 GND 0.005205f
C2058 VDD.n1077 GND 0.006467f
C2059 VDD.n1078 GND 0.005205f
C2060 VDD.n1079 GND 0.006467f
C2061 VDD.n1080 GND 0.005205f
C2062 VDD.n1081 GND 0.006467f
C2063 VDD.n1082 GND 0.005205f
C2064 VDD.n1083 GND 0.006467f
C2065 VDD.n1084 GND 0.005205f
C2066 VDD.n1085 GND 0.006467f
C2067 VDD.t46 GND 0.089332f
C2068 VDD.t47 GND 0.10348f
C2069 VDD.t44 GND 0.482813f
C2070 VDD.n1086 GND 0.068834f
C2071 VDD.n1087 GND 0.04271f
C2072 VDD.n1088 GND 0.010619f
C2073 VDD.n1089 GND 0.006467f
C2074 VDD.n1090 GND 0.005205f
C2075 VDD.n1091 GND 0.006467f
C2076 VDD.n1092 GND 0.005205f
C2077 VDD.n1093 GND 0.006467f
C2078 VDD.n1094 GND 0.005205f
C2079 VDD.n1095 GND 0.006467f
C2080 VDD.n1096 GND 0.005205f
C2081 VDD.n1097 GND 0.006467f
C2082 VDD.n1098 GND 0.005205f
C2083 VDD.n1099 GND 0.00432f
C2084 VDD.n1100 GND 0.006467f
C2085 VDD.n1101 GND 0.005205f
C2086 VDD.n1103 GND 0.006467f
C2087 VDD.n1104 GND 0.006467f
C2088 VDD.n1106 GND 0.006467f
C2089 VDD.n1107 GND 0.005205f
C2090 VDD.n1108 GND 0.006467f
C2091 VDD.n1109 GND 0.006467f
C2092 VDD.n1110 GND 0.006467f
C2093 VDD.n1111 GND 0.005205f
C2094 VDD.n1112 GND 0.006467f
C2095 VDD.n1114 GND 0.006467f
C2096 VDD.n1116 GND 0.006467f
C2097 VDD.n1117 GND 0.005205f
C2098 VDD.n1118 GND 0.006467f
C2099 VDD.n1119 GND 0.006467f
C2100 VDD.n1120 GND 0.006467f
C2101 VDD.n1121 GND 0.005205f
C2102 VDD.n1122 GND 0.006467f
C2103 VDD.n1124 GND 0.006467f
C2104 VDD.n1126 GND 0.006467f
C2105 VDD.n1127 GND 0.004346f
C2106 VDD.n1128 GND 0.006467f
C2107 VDD.n1129 GND 0.006467f
C2108 VDD.n1130 GND 0.006467f
C2109 VDD.n1131 GND 0.004346f
C2110 VDD.n1132 GND 0.006467f
C2111 VDD.n1134 GND 0.006467f
C2112 VDD.n1136 GND 0.006467f
C2113 VDD.n1137 GND 0.005205f
C2114 VDD.n1138 GND 0.006467f
C2115 VDD.n1139 GND 0.006467f
C2116 VDD.n1140 GND 0.006467f
C2117 VDD.n1141 GND 0.005205f
C2118 VDD.n1142 GND 0.006467f
C2119 VDD.n1144 GND 0.006467f
C2120 VDD.n1146 GND 0.006467f
C2121 VDD.n1147 GND 0.005205f
C2122 VDD.n1148 GND 0.006467f
C2123 VDD.n1149 GND 0.006467f
C2124 VDD.n1150 GND 0.006467f
C2125 VDD.n1151 GND 0.006467f
C2126 VDD.n1152 GND 0.005205f
C2127 VDD.n1153 GND 0.006467f
C2128 VDD.n1155 GND 0.006467f
C2129 VDD.n1156 GND 0.006467f
C2130 VDD.n1158 GND 0.006467f
C2131 VDD.n1159 GND 0.005205f
C2132 VDD.n1160 GND 0.006467f
C2133 VDD.n1161 GND 0.006467f
C2134 VDD.n1162 GND 0.006467f
C2135 VDD.n1163 GND 0.00354f
C2136 VDD.n1164 GND 0.010619f
C2137 VDD.n1165 GND 0.006467f
C2138 VDD.n1167 GND 0.006467f
C2139 VDD.n1169 GND 0.006467f
C2140 VDD.n1170 GND 0.005205f
C2141 VDD.n1171 GND 0.006467f
C2142 VDD.n1172 GND 0.006467f
C2143 VDD.n1173 GND 0.006467f
C2144 VDD.n1174 GND 0.005205f
C2145 VDD.n1175 GND 0.006467f
C2146 VDD.n1177 GND 0.006467f
C2147 VDD.n1179 GND 0.006467f
C2148 VDD.n1180 GND 0.005205f
C2149 VDD.n1181 GND 0.006467f
C2150 VDD.n1182 GND 0.006467f
C2151 VDD.n1183 GND 0.006467f
C2152 VDD.n1184 GND 0.005205f
C2153 VDD.n1185 GND 0.006467f
C2154 VDD.n1187 GND 0.006467f
C2155 VDD.n1189 GND 0.006467f
C2156 VDD.n1190 GND 0.005205f
C2157 VDD.n1191 GND 0.006467f
C2158 VDD.n1192 GND 0.006467f
C2159 VDD.n1193 GND 0.006467f
C2160 VDD.n1194 GND 0.006467f
C2161 VDD.n1195 GND 0.005205f
C2162 VDD.n1196 GND 0.006467f
C2163 VDD.n1198 GND 0.006467f
C2164 VDD.n1200 GND 0.006467f
C2165 VDD.n1201 GND 0.002733f
C2166 VDD.n1202 GND 0.008016f
C2167 VDD.n1203 GND 0.002472f
C2168 VDD.n1204 GND 0.014463f
C2169 VDD.n1205 GND 0.014445f
C2170 VDD.n1206 GND 0.00432f
C2171 VDD.n1207 GND 0.014445f
C2172 VDD.n1208 GND 0.487185f
C2173 VDD.n1209 GND 0.014445f
C2174 VDD.n1210 GND 0.00432f
C2175 VDD.n1211 GND 0.014445f
C2176 VDD.n1212 GND 0.006467f
C2177 VDD.n1213 GND 0.006467f
C2178 VDD.n1214 GND 0.005205f
C2179 VDD.n1215 GND 0.006467f
C2180 VDD.n1216 GND 0.38361f
C2181 VDD.n1217 GND 0.006467f
C2182 VDD.n1218 GND 0.005205f
C2183 VDD.n1219 GND 0.006467f
C2184 VDD.n1220 GND 0.006467f
C2185 VDD.n1221 GND 0.006467f
C2186 VDD.n1222 GND 0.005205f
C2187 VDD.n1223 GND 0.006467f
C2188 VDD.n1224 GND 0.218658f
C2189 VDD.n1225 GND 0.006467f
C2190 VDD.n1226 GND 0.005205f
C2191 VDD.n1227 GND 0.006467f
C2192 VDD.n1228 GND 0.006467f
C2193 VDD.n1229 GND 0.006467f
C2194 VDD.n1230 GND 0.005205f
C2195 VDD.n1231 GND 0.006467f
C2196 VDD.n1232 GND 0.38361f
C2197 VDD.n1233 GND 0.006467f
C2198 VDD.n1234 GND 0.005205f
C2199 VDD.n1235 GND 0.006467f
C2200 VDD.n1236 GND 0.006467f
C2201 VDD.n1237 GND 0.006467f
C2202 VDD.n1238 GND 0.005205f
C2203 VDD.n1239 GND 0.006467f
C2204 VDD.n1240 GND 0.38361f
C2205 VDD.n1241 GND 0.006467f
C2206 VDD.n1242 GND 0.005205f
C2207 VDD.n1243 GND 0.006467f
C2208 VDD.n1244 GND 0.006467f
C2209 VDD.n1245 GND 0.006467f
C2210 VDD.n1246 GND 0.005205f
C2211 VDD.n1247 GND 0.006467f
C2212 VDD.n1248 GND 0.38361f
C2213 VDD.n1249 GND 0.006467f
C2214 VDD.n1250 GND 0.005205f
C2215 VDD.n1251 GND 0.006467f
C2216 VDD.n1252 GND 0.006467f
C2217 VDD.n1253 GND 0.006467f
C2218 VDD.n1254 GND 0.005205f
C2219 VDD.n1255 GND 0.006467f
C2220 VDD.n1256 GND 0.38361f
C2221 VDD.n1257 GND 0.006467f
C2222 VDD.n1258 GND 0.005205f
C2223 VDD.n1259 GND 0.006445f
C2224 VDD.t76 GND 0.114213f
C2225 VDD.t77 GND 0.110011f
C2226 VDD.n1260 GND 0.30549f
C2227 VDD.t73 GND 0.110011f
C2228 VDD.n1261 GND 0.161408f
C2229 VDD.n1262 GND 1.16178f
C2230 VDD.n1263 GND 0.01174f
C2231 VDD.n1264 GND 0.006445f
C2232 VDD.n1265 GND 0.005205f
C2233 VDD.n1266 GND 0.006467f
C2234 VDD.n1267 GND 0.38361f
C2235 VDD.n1268 GND 0.006467f
C2236 VDD.n1269 GND 0.005205f
C2237 VDD.n1270 GND 0.006467f
C2238 VDD.n1271 GND 0.006467f
C2239 VDD.n1272 GND 0.006467f
C2240 VDD.n1273 GND 0.005205f
C2241 VDD.n1274 GND 0.006467f
C2242 VDD.n1275 GND 0.38361f
C2243 VDD.n1276 GND 0.006467f
C2244 VDD.n1277 GND 0.005205f
C2245 VDD.n1278 GND 0.006467f
C2246 VDD.n1279 GND 0.006467f
C2247 VDD.n1280 GND 0.006467f
C2248 VDD.n1281 GND 0.005205f
C2249 VDD.n1282 GND 0.006467f
C2250 VDD.n1283 GND 0.38361f
C2251 VDD.n1284 GND 0.006467f
C2252 VDD.n1285 GND 0.005205f
C2253 VDD.n1286 GND 0.006467f
C2254 VDD.n1287 GND 0.006467f
C2255 VDD.n1288 GND 0.006467f
C2256 VDD.n1289 GND 0.005205f
C2257 VDD.n1290 GND 0.006467f
C2258 VDD.n1291 GND 0.38361f
C2259 VDD.n1292 GND 0.006467f
C2260 VDD.n1293 GND 0.005205f
C2261 VDD.n1294 GND 0.006467f
C2262 VDD.n1295 GND 0.006467f
C2263 VDD.n1296 GND 0.006467f
C2264 VDD.n1297 GND 0.005205f
C2265 VDD.n1298 GND 0.006467f
C2266 VDD.n1299 GND 0.218658f
C2267 VDD.n1300 GND 0.006467f
C2268 VDD.n1301 GND 0.005205f
C2269 VDD.n1302 GND 0.006467f
C2270 VDD.n1303 GND 0.006467f
C2271 VDD.n1304 GND 0.014445f
C2272 VDD.n1305 GND 0.006467f
C2273 VDD.n1306 GND 0.006467f
C2274 VDD.n1307 GND 0.005205f
C2275 VDD.n1308 GND 0.006467f
C2276 VDD.n1309 GND 0.38361f
C2277 VDD.n1310 GND 0.006467f
C2278 VDD.n1311 GND 0.005205f
C2279 VDD.n1312 GND 0.006467f
C2280 VDD.n1313 GND 0.006467f
C2281 VDD.n1314 GND 0.006467f
C2282 VDD.n1315 GND 0.005205f
C2283 VDD.n1316 GND 0.005205f
C2284 VDD.n1317 GND 0.006467f
C2285 VDD.n1318 GND 0.006467f
C2286 VDD.n1319 GND 0.006467f
C2287 VDD.n1320 GND 0.006467f
C2288 VDD.n1321 GND 0.005205f
C2289 VDD.n1322 GND 0.006467f
C2290 VDD.n1324 GND 0.006467f
C2291 VDD.n1325 GND 0.006467f
C2292 VDD.n1327 GND 0.006467f
C2293 VDD.n1328 GND 0.005205f
C2294 VDD.n1329 GND 0.00432f
C2295 VDD.n1330 GND 0.014463f
C2296 VDD.n1331 GND 0.014445f
C2297 VDD.n1332 GND 0.00432f
C2298 VDD.n1333 GND 0.014445f
C2299 VDD.n1334 GND 0.487185f
C2300 VDD.n1335 GND 0.014445f
C2301 VDD.n1336 GND 0.014463f
C2302 VDD.n1337 GND 0.002472f
C2303 VDD.t40 GND 0.089332f
C2304 VDD.t39 GND 0.10348f
C2305 VDD.t38 GND 0.482813f
C2306 VDD.n1338 GND 0.068834f
C2307 VDD.n1339 GND 0.04271f
C2308 VDD.n1340 GND 0.008016f
C2309 VDD.n1341 GND 0.002733f
C2310 VDD.n1342 GND 0.006467f
C2311 VDD.n1343 GND 0.006467f
C2312 VDD.n1344 GND 0.006467f
C2313 VDD.n1345 GND 0.005205f
C2314 VDD.n1346 GND 0.005205f
C2315 VDD.n1347 GND 0.005205f
C2316 VDD.n1348 GND 0.006338f
C2317 VDD.n1349 GND 1.08458f
C2318 VDD.n1351 GND 0.005205f
C2319 VDD.n1352 GND 0.005205f
C2320 VDD.n1353 GND 0.006467f
C2321 VDD.n1355 GND 0.006467f
C2322 VDD.n1356 GND 0.006467f
C2323 VDD.n1357 GND 0.005205f
C2324 VDD.n1358 GND 0.005205f
C2325 VDD.n1359 GND 0.005153f
C2326 VDD.n1360 GND 0.006467f
C2327 VDD.n1362 GND 0.006467f
C2328 VDD.n1363 GND 0.006467f
C2329 VDD.n1364 GND 0.00354f
C2330 VDD.n1365 GND 0.005205f
C2331 VDD.n1366 GND 0.005205f
C2332 VDD.n1367 GND 0.006467f
C2333 VDD.n1369 GND 0.006467f
C2334 VDD.n1370 GND 0.006467f
C2335 VDD.n1371 GND 0.005205f
C2336 VDD.n1372 GND 0.005205f
C2337 VDD.n1373 GND 0.005205f
C2338 VDD.n1374 GND 0.006467f
C2339 VDD.n1376 GND 0.006467f
C2340 VDD.n1377 GND 0.006467f
C2341 VDD.n1378 GND 0.005205f
C2342 VDD.n1379 GND 0.005205f
C2343 VDD.n1380 GND 0.005205f
C2344 VDD.n1381 GND 0.006467f
C2345 VDD.n1383 GND 0.006467f
C2346 VDD.n1384 GND 0.006467f
C2347 VDD.n1385 GND 0.005205f
C2348 VDD.n1386 GND 0.006467f
C2349 VDD.n1387 GND 0.006467f
C2350 VDD.n1388 GND 0.006467f
C2351 VDD.n1389 GND 0.010619f
C2352 VDD.n1390 GND 0.004346f
C2353 VDD.n1391 GND 0.005205f
C2354 VDD.n1392 GND 0.006467f
C2355 VDD.n1394 GND 0.006467f
C2356 VDD.n1395 GND 0.005205f
C2357 VDD.n1396 GND 0.006467f
C2358 VDD.n1398 GND 0.006467f
C2359 VDD.n1399 GND 0.006467f
C2360 VDD.n1400 GND 0.005205f
C2361 VDD.n1402 GND 1.08458f
C2362 VDD.t36 GND 0.041419f
C2363 VDD.t37 GND 0.056208f
C2364 VDD.t35 GND 0.369485f
C2365 VDD.n1403 GND 0.058137f
C2366 VDD.n1404 GND 0.040639f
C2367 VDD.n1405 GND 0.006285f
C2368 VDD.n1406 GND 0.004398f
C2369 VDD.n1407 GND 0.004398f
C2370 VDD.n1408 GND 0.004398f
C2371 VDD.n1409 GND 0.004398f
C2372 VDD.n1410 GND 0.004398f
C2373 VDD.n1411 GND 0.004398f
C2374 VDD.n1412 GND 0.004398f
C2375 VDD.n1413 GND 0.004398f
C2376 VDD.n1414 GND 0.004398f
C2377 VDD.n1415 GND 0.004398f
C2378 VDD.n1416 GND 0.004398f
C2379 VDD.n1417 GND 0.004398f
C2380 VDD.n1418 GND 0.004398f
C2381 VDD.n1419 GND 0.004398f
C2382 VDD.n1420 GND 0.004398f
C2383 VDD.n1421 GND 0.004398f
C2384 VDD.n1422 GND 0.004398f
C2385 VDD.n1423 GND 0.004398f
C2386 VDD.n1424 GND 0.004398f
C2387 VDD.n1425 GND 0.004398f
C2388 VDD.n1426 GND 0.004398f
C2389 VDD.n1427 GND 0.004398f
C2390 VDD.n1428 GND 0.004398f
C2391 VDD.n1429 GND 0.004398f
C2392 VDD.n1430 GND 0.004398f
C2393 VDD.n1431 GND 0.004398f
C2394 VDD.n1432 GND 0.004398f
C2395 VDD.n1433 GND 0.004398f
C2396 VDD.n1434 GND 0.004398f
C2397 VDD.n1435 GND 0.004398f
C2398 VDD.n1436 GND 0.004398f
C2399 VDD.n1437 GND 0.004398f
C2400 VDD.n1438 GND 0.004398f
C2401 VDD.n1439 GND 0.004398f
C2402 VDD.n1440 GND 0.004398f
C2403 VDD.n1441 GND 0.004398f
C2404 VDD.n1442 GND 0.004398f
C2405 VDD.n1443 GND 0.004398f
C2406 VDD.n1444 GND 0.004398f
C2407 VDD.n1445 GND 0.004398f
C2408 VDD.n1446 GND 0.004398f
C2409 VDD.n1447 GND 0.004398f
C2410 VDD.n1448 GND 0.004398f
C2411 VDD.n1449 GND 0.004398f
C2412 VDD.n1450 GND 0.004398f
C2413 VDD.n1451 GND 0.004398f
C2414 VDD.n1452 GND 0.004398f
C2415 VDD.n1453 GND 0.004398f
C2416 VDD.n1454 GND 0.004398f
C2417 VDD.n1455 GND 0.004398f
C2418 VDD.n1456 GND 0.004398f
C2419 VDD.n1457 GND 0.004398f
C2420 VDD.n1458 GND 0.004398f
C2421 VDD.n1459 GND 0.004398f
C2422 VDD.n1460 GND 0.004398f
C2423 VDD.n1461 GND 0.004398f
C2424 VDD.n1462 GND 0.004398f
C2425 VDD.n1463 GND 0.004398f
C2426 VDD.n1464 GND 0.004398f
C2427 VDD.n1465 GND 0.004398f
C2428 VDD.n1466 GND 0.004398f
C2429 VDD.n1467 GND 0.004398f
C2430 VDD.n1468 GND 0.004398f
C2431 VDD.n1469 GND 0.004398f
C2432 VDD.n1470 GND 0.004398f
C2433 VDD.n1471 GND 0.004398f
C2434 VDD.n1472 GND 0.004398f
C2435 VDD.n1473 GND 0.004398f
C2436 VDD.n1474 GND 0.004398f
C2437 VDD.n1475 GND 0.004398f
C2438 VDD.n1476 GND 0.004398f
C2439 VDD.n1477 GND 0.004398f
C2440 VDD.n1478 GND 0.004398f
C2441 VDD.n1479 GND 0.004398f
C2442 VDD.n1480 GND 0.004398f
C2443 VDD.n1481 GND 0.004398f
C2444 VDD.n1482 GND 0.004398f
C2445 VDD.n1483 GND 0.004398f
C2446 VDD.n1484 GND 0.004398f
C2447 VDD.n1485 GND 0.004398f
C2448 VDD.n1486 GND 0.004398f
C2449 VDD.n1487 GND 0.004398f
C2450 VDD.n1488 GND 0.004398f
C2451 VDD.n1489 GND 0.004398f
C2452 VDD.n1490 GND 0.004398f
C2453 VDD.n1491 GND 0.004398f
C2454 VDD.n1492 GND 0.004398f
C2455 VDD.n1493 GND 0.004398f
C2456 VDD.n1494 GND 0.004398f
C2457 VDD.n1495 GND 0.004398f
C2458 VDD.n1496 GND 0.004398f
C2459 VDD.n1497 GND 0.004398f
C2460 VDD.n1498 GND 0.004398f
C2461 VDD.n1499 GND 0.004398f
C2462 VDD.n1500 GND 0.004398f
C2463 VDD.n1501 GND 0.004398f
C2464 VDD.n1502 GND 0.004398f
C2465 VDD.n1503 GND 0.004398f
C2466 VDD.n1504 GND 0.004398f
C2467 VDD.n1505 GND 0.004398f
C2468 VDD.n1506 GND 0.004398f
C2469 VDD.n1507 GND 0.004398f
C2470 VDD.n1508 GND 0.004398f
C2471 VDD.n1509 GND 0.004398f
C2472 VDD.n1510 GND 0.004398f
C2473 VDD.n1511 GND 0.004398f
C2474 VDD.n1512 GND 0.004398f
C2475 VDD.n1513 GND 0.004398f
C2476 VDD.n1514 GND 0.004398f
C2477 VDD.n1515 GND 0.004398f
C2478 VDD.n1516 GND 0.004398f
C2479 VDD.n1517 GND 0.004398f
C2480 VDD.n1518 GND 0.004398f
C2481 VDD.n1519 GND 0.004398f
C2482 VDD.n1520 GND 0.004398f
C2483 VDD.n1521 GND 0.004398f
C2484 VDD.n1522 GND 0.004398f
C2485 VDD.n1523 GND 0.004398f
C2486 VDD.n1524 GND 0.004398f
C2487 VDD.n1525 GND 0.004398f
C2488 VDD.n1526 GND 0.004398f
C2489 VDD.n1527 GND 0.004398f
C2490 VDD.n1528 GND 0.004398f
C2491 VDD.n1529 GND 0.004398f
C2492 VDD.n1530 GND 0.004398f
C2493 VDD.n1531 GND 0.004398f
C2494 VDD.n1532 GND 0.004398f
C2495 VDD.n1533 GND 0.004398f
C2496 VDD.n1534 GND 0.004398f
C2497 VDD.n1535 GND 0.004398f
C2498 VDD.n1536 GND 0.004398f
C2499 VDD.n1537 GND 0.009619f
C2500 VDD.n1538 GND 0.009619f
C2501 VDD.n1539 GND 0.010235f
C2502 VDD.n1540 GND 0.010235f
C2503 VDD.n1541 GND 0.003686f
C2504 VDD.n1542 GND 0.004398f
C2505 VDD.n1543 GND 0.004398f
C2506 VDD.n1544 GND 0.00291f
C2507 VDD.n1545 GND 0.004398f
C2508 VDD.n1546 GND 0.004398f
C2509 VDD.n1547 GND 0.004398f
C2510 VDD.n1548 GND 0.004398f
C2511 VDD.n1549 GND 0.004398f
C2512 VDD.n1550 GND 0.004398f
C2513 VDD.n1551 GND 0.004398f
C2514 VDD.n1552 GND 0.004398f
C2515 VDD.n1553 GND 0.066313f
C2516 VDD.n1554 GND 0.004398f
C2517 VDD.n1555 GND 0.004398f
C2518 VDD.n1556 GND 0.004398f
C2519 VDD.n1557 GND 0.004398f
C2520 VDD.n1558 GND 0.004398f
C2521 VDD.n1559 GND 0.004398f
C2522 VDD.n1560 GND 0.004398f
C2523 VDD.n1561 GND 0.004398f
C2524 VDD.n1562 GND 0.004398f
C2525 VDD.n1563 GND 0.004398f
C2526 VDD.n1564 GND 0.72886f
C2527 VDD.n1566 GND 0.010235f
C2528 VDD.n1567 GND 0.010235f
C2529 VDD.n1568 GND 0.009619f
C2530 VDD.n1569 GND 0.004398f
C2531 VDD.n1570 GND 0.004398f
C2532 VDD.n1571 GND 0.260855f
C2533 VDD.n1572 GND 0.004398f
C2534 VDD.n1573 GND 0.004398f
C2535 VDD.n1574 GND 0.004398f
C2536 VDD.n1575 GND 0.004398f
C2537 VDD.n1576 GND 0.004398f
C2538 VDD.n1577 GND 0.260855f
C2539 VDD.n1578 GND 0.004398f
C2540 VDD.n1579 GND 0.004398f
C2541 VDD.n1580 GND 0.004398f
C2542 VDD.n1581 GND 0.004398f
C2543 VDD.n1582 GND 0.004398f
C2544 VDD.n1583 GND 0.260855f
C2545 VDD.n1584 GND 0.004398f
C2546 VDD.n1585 GND 0.004398f
C2547 VDD.n1586 GND 0.004398f
C2548 VDD.n1587 GND 0.004398f
C2549 VDD.n1588 GND 0.004398f
C2550 VDD.n1589 GND 0.247429f
C2551 VDD.n1590 GND 0.004398f
C2552 VDD.n1591 GND 0.004398f
C2553 VDD.n1592 GND 0.004398f
C2554 VDD.n1593 GND 0.004398f
C2555 VDD.n1594 GND 0.004398f
C2556 VDD.n1595 GND 0.260855f
C2557 VDD.n1596 GND 0.004398f
C2558 VDD.n1597 GND 0.004398f
C2559 VDD.n1598 GND 0.004398f
C2560 VDD.n1599 GND 0.004398f
C2561 VDD.n1600 GND 0.004398f
C2562 VDD.n1601 GND 0.260855f
C2563 VDD.n1602 GND 0.004398f
C2564 VDD.n1603 GND 0.004398f
C2565 VDD.n1604 GND 0.004398f
C2566 VDD.n1605 GND 0.004398f
C2567 VDD.n1606 GND 0.004398f
C2568 VDD.n1607 GND 0.260855f
C2569 VDD.n1608 GND 0.004398f
C2570 VDD.n1609 GND 0.004398f
C2571 VDD.n1610 GND 0.004398f
C2572 VDD.n1611 GND 0.004398f
C2573 VDD.n1612 GND 0.004398f
C2574 VDD.n1613 GND 0.260855f
C2575 VDD.n1614 GND 0.004398f
C2576 VDD.n1615 GND 0.004398f
C2577 VDD.n1616 GND 0.004398f
C2578 VDD.n1617 GND 0.004398f
C2579 VDD.n1618 GND 0.004398f
C2580 VDD.n1619 GND 0.260855f
C2581 VDD.n1620 GND 0.004398f
C2582 VDD.n1621 GND 0.004398f
C2583 VDD.n1622 GND 0.004398f
C2584 VDD.n1623 GND 0.004398f
C2585 VDD.n1624 GND 0.004398f
C2586 VDD.n1625 GND 0.260855f
C2587 VDD.n1626 GND 0.004398f
C2588 VDD.n1627 GND 0.004398f
C2589 VDD.n1628 GND 0.004398f
C2590 VDD.n1629 GND 0.004398f
C2591 VDD.n1630 GND 0.004398f
C2592 VDD.n1631 GND 0.199477f
C2593 VDD.n1632 GND 0.004398f
C2594 VDD.n1633 GND 0.004398f
C2595 VDD.n1634 GND 0.004398f
C2596 VDD.n1635 GND 0.004398f
C2597 VDD.n1636 GND 0.004398f
C2598 VDD.n1637 GND 0.260855f
C2599 VDD.n1638 GND 0.004398f
C2600 VDD.n1639 GND 0.004398f
C2601 VDD.n1640 GND 0.004398f
C2602 VDD.n1641 GND 0.004398f
C2603 VDD.n1642 GND 0.004398f
C2604 VDD.n1643 GND 0.174543f
C2605 VDD.n1644 GND 0.004398f
C2606 VDD.n1645 GND 0.004398f
C2607 VDD.n1646 GND 0.004398f
C2608 VDD.n1647 GND 0.004398f
C2609 VDD.n1648 GND 0.004398f
C2610 VDD.n1649 GND 0.260855f
C2611 VDD.n1650 GND 0.004398f
C2612 VDD.n1651 GND 0.004398f
C2613 VDD.n1652 GND 0.004398f
C2614 VDD.n1653 GND 0.004398f
C2615 VDD.n1654 GND 0.004398f
C2616 VDD.n1655 GND 0.260855f
C2617 VDD.n1656 GND 0.004398f
C2618 VDD.n1657 GND 0.004398f
C2619 VDD.n1658 GND 0.004398f
C2620 VDD.n1659 GND 0.004398f
C2621 VDD.n1660 GND 0.004398f
C2622 VDD.n1661 GND 0.260855f
C2623 VDD.n1662 GND 0.004398f
C2624 VDD.n1663 GND 0.004398f
C2625 VDD.n1664 GND 0.004398f
C2626 VDD.n1665 GND 0.004398f
C2627 VDD.n1666 GND 0.004398f
C2628 VDD.n1667 GND 0.260855f
C2629 VDD.n1668 GND 0.004398f
C2630 VDD.n1669 GND 0.004398f
C2631 VDD.n1670 GND 0.004398f
C2632 VDD.n1671 GND 0.004398f
C2633 VDD.n1672 GND 0.004398f
C2634 VDD.n1673 GND 0.260855f
C2635 VDD.n1674 GND 0.004398f
C2636 VDD.n1675 GND 0.004398f
C2637 VDD.n1676 GND 0.004398f
C2638 VDD.n1677 GND 0.004398f
C2639 VDD.n1678 GND 0.004398f
C2640 VDD.n1679 GND 0.260855f
C2641 VDD.n1680 GND 0.004398f
C2642 VDD.n1681 GND 0.004398f
C2643 VDD.n1682 GND 0.004398f
C2644 VDD.n1683 GND 0.004398f
C2645 VDD.n1684 GND 0.004398f
C2646 VDD.n1685 GND 0.232084f
C2647 VDD.n1686 GND 0.004398f
C2648 VDD.n1687 GND 0.004398f
C2649 VDD.n1688 GND 0.004398f
C2650 VDD.n1689 GND 0.004398f
C2651 VDD.n1690 GND 0.004398f
C2652 VDD.n1691 GND 0.260855f
C2653 VDD.n1692 GND 0.004398f
C2654 VDD.n1693 GND 0.004398f
C2655 VDD.n1694 GND 0.004398f
C2656 VDD.n1695 GND 0.004398f
C2657 VDD.n1696 GND 0.004398f
C2658 VDD.n1697 GND 0.257019f
C2659 VDD.n1698 GND 0.004398f
C2660 VDD.n1699 GND 0.004398f
C2661 VDD.n1700 GND 0.004398f
C2662 VDD.n1701 GND 0.004398f
C2663 VDD.n1702 GND 0.004398f
C2664 VDD.n1703 GND 0.260855f
C2665 VDD.n1704 GND 0.004398f
C2666 VDD.n1705 GND 0.004398f
C2667 VDD.n1706 GND 0.004398f
C2668 VDD.n1707 GND 0.004398f
C2669 VDD.n1708 GND 0.004398f
C2670 VDD.n1709 GND 0.260855f
C2671 VDD.n1710 GND 0.004398f
C2672 VDD.n1711 GND 0.004398f
C2673 VDD.n1712 GND 0.004398f
C2674 VDD.n1713 GND 0.004398f
C2675 VDD.n1714 GND 0.004398f
C2676 VDD.n1715 GND 0.260855f
C2677 VDD.n1716 GND 0.004398f
C2678 VDD.n1717 GND 0.004398f
C2679 VDD.n1718 GND 0.004398f
C2680 VDD.n1719 GND 0.004398f
C2681 VDD.n1720 GND 0.004398f
C2682 VDD.n1721 GND 0.232084f
C2683 VDD.n1722 GND 0.004398f
C2684 VDD.n1723 GND 0.004398f
C2685 VDD.n1724 GND 0.004398f
C2686 VDD.n1725 GND 0.004398f
C2687 VDD.n1726 GND 0.004398f
C2688 VDD.n1727 GND 0.260855f
C2689 VDD.n1728 GND 0.004398f
C2690 VDD.n1729 GND 0.004398f
C2691 VDD.n1730 GND 0.004398f
C2692 VDD.n1731 GND 0.004398f
C2693 VDD.n1732 GND 0.004398f
C2694 VDD.n1733 GND 0.20715f
C2695 VDD.n1734 GND 0.004398f
C2696 VDD.n1735 GND 0.004398f
C2697 VDD.n1736 GND 0.004398f
C2698 VDD.n1737 GND 0.004398f
C2699 VDD.n1738 GND 0.004398f
C2700 VDD.n1739 GND 0.260855f
C2701 VDD.n1740 GND 0.004398f
C2702 VDD.n1741 GND 0.004398f
C2703 VDD.n1742 GND 0.004398f
C2704 VDD.n1743 GND 0.004398f
C2705 VDD.n1744 GND 0.004398f
C2706 VDD.n1745 GND 0.260855f
C2707 VDD.n1746 GND 0.004398f
C2708 VDD.n1747 GND 0.004398f
C2709 VDD.n1748 GND 0.004398f
C2710 VDD.n1749 GND 0.004398f
C2711 VDD.n1750 GND 0.004398f
C2712 VDD.n1751 GND 0.260855f
C2713 VDD.n1752 GND 0.004398f
C2714 VDD.n1753 GND 0.004398f
C2715 VDD.n1754 GND 0.004398f
C2716 VDD.n1755 GND 0.004398f
C2717 VDD.n1756 GND 0.004398f
C2718 VDD.n1757 GND 0.260855f
C2719 VDD.n1758 GND 0.004398f
C2720 VDD.n1759 GND 0.004398f
C2721 VDD.n1760 GND 0.004398f
C2722 VDD.n1761 GND 0.004398f
C2723 VDD.n1762 GND 0.004398f
C2724 VDD.n1763 GND 0.174543f
C2725 VDD.n1764 GND 0.004398f
C2726 VDD.n1765 GND 0.004398f
C2727 VDD.n1766 GND 0.004398f
C2728 VDD.n1767 GND 0.004398f
C2729 VDD.n1768 GND 0.004398f
C2730 VDD.n1769 GND 0.260855f
C2731 VDD.n1770 GND 0.004398f
C2732 VDD.n1771 GND 0.004398f
C2733 VDD.n1772 GND 0.004398f
C2734 VDD.n1773 GND 0.004398f
C2735 VDD.n1774 GND 0.004398f
C2736 VDD.n1775 GND 0.149608f
C2737 VDD.n1776 GND 0.004398f
C2738 VDD.n1777 GND 0.004398f
C2739 VDD.n1778 GND 0.004398f
C2740 VDD.n1779 GND 0.004398f
C2741 VDD.n1780 GND 0.004398f
C2742 VDD.n1781 GND 0.260855f
C2743 VDD.n1782 GND 0.004398f
C2744 VDD.n1783 GND 0.004398f
C2745 VDD.n1784 GND 0.004398f
C2746 VDD.n1785 GND 0.004398f
C2747 VDD.n1786 GND 0.004398f
C2748 VDD.n1787 GND 0.260855f
C2749 VDD.n1788 GND 0.004398f
C2750 VDD.n1789 GND 0.004398f
C2751 VDD.n1790 GND 0.004398f
C2752 VDD.n1791 GND 0.004398f
C2753 VDD.n1792 GND 0.004398f
C2754 VDD.n1793 GND 0.260855f
C2755 VDD.n1794 GND 0.004398f
C2756 VDD.n1795 GND 0.004398f
C2757 VDD.n1796 GND 0.004398f
C2758 VDD.n1797 GND 0.004398f
C2759 VDD.n1798 GND 0.004398f
C2760 VDD.n1799 GND 0.260855f
C2761 VDD.n1800 GND 0.004398f
C2762 VDD.n1801 GND 0.004398f
C2763 VDD.n1802 GND 0.004398f
C2764 VDD.n1803 GND 0.004398f
C2765 VDD.n1804 GND 0.004398f
C2766 VDD.n1805 GND 0.260855f
C2767 VDD.n1806 GND 0.004398f
C2768 VDD.n1807 GND 0.004398f
C2769 VDD.n1808 GND 0.004398f
C2770 VDD.n1809 GND 0.004398f
C2771 VDD.n1810 GND 0.004398f
C2772 VDD.n1811 GND 0.260855f
C2773 VDD.n1812 GND 0.004398f
C2774 VDD.n1813 GND 0.004398f
C2775 VDD.n1814 GND 0.004398f
C2776 VDD.n1815 GND 0.004398f
C2777 VDD.n1816 GND 0.004398f
C2778 VDD.n1817 GND 0.004398f
C2779 VDD.n1818 GND 0.004398f
C2780 VDD.n1819 GND 0.168789f
C2781 VDD.n1820 GND 0.004398f
C2782 VDD.n1821 GND 0.004398f
C2783 VDD.n1822 GND 0.004398f
C2784 VDD.n1823 GND 0.004398f
C2785 VDD.n1824 GND 0.004398f
C2786 VDD.n1825 GND 0.260855f
C2787 VDD.n1826 GND 0.004398f
C2788 VDD.n1827 GND 0.004398f
C2789 VDD.n1828 GND 0.004398f
C2790 VDD.n1829 GND 0.004398f
C2791 VDD.n1830 GND 0.004398f
C2792 VDD.n1831 GND 0.004398f
C2793 VDD.n1832 GND 0.004398f
C2794 VDD.n1833 GND 0.009619f
C2795 VDD.n1834 GND 0.010168f
C2796 VDD.n1835 GND 0.009686f
C2797 VDD.n1836 GND 0.004398f
C2798 VDD.n1837 GND 0.003686f
C2799 VDD.n1838 GND 0.006285f
C2800 VDD.n1839 GND 0.00291f
C2801 VDD.n1840 GND 0.004398f
C2802 VDD.n1841 GND 0.004398f
C2803 VDD.n1842 GND 0.004398f
C2804 VDD.n1843 GND 0.004398f
C2805 VDD.n1844 GND 0.004398f
C2806 VDD.n1845 GND 0.004398f
C2807 VDD.n1846 GND 0.004398f
C2808 VDD.n1847 GND 0.004398f
C2809 VDD.n1848 GND 0.004398f
C2810 VDD.n1849 GND 0.004398f
C2811 VDD.n1850 GND 0.004398f
C2812 VDD.n1851 GND 0.004398f
C2813 VDD.n1852 GND 0.004398f
C2814 VDD.n1853 GND 0.004398f
C2815 VDD.n1854 GND 0.004398f
C2816 VDD.n1855 GND 0.004398f
C2817 VDD.n1856 GND 0.004398f
C2818 VDD.n1857 GND 0.004398f
C2819 VDD.n1858 GND 0.004398f
C2820 VDD.n1859 GND 0.004398f
C2821 VDD.n1860 GND 0.004398f
C2822 VDD.n1861 GND 0.004398f
C2823 VDD.n1862 GND 0.004398f
C2824 VDD.n1863 GND 0.010235f
C2825 VDD.n1864 GND 0.010235f
C2826 VDD.n1865 GND 0.009619f
C2827 VDD.n1866 GND 0.009619f
C2828 VDD.n1867 GND 0.004398f
C2829 VDD.n1868 GND 0.004398f
C2830 VDD.n1869 GND 0.004398f
C2831 VDD.n1870 GND 0.004398f
C2832 VDD.n1871 GND 0.260855f
C2833 VDD.n1872 GND 0.004398f
C2834 VDD.n1873 GND 0.004398f
C2835 VDD.n1874 GND 0.004398f
C2836 VDD.n1875 GND 0.004398f
C2837 VDD.n1876 GND 0.004398f
C2838 VDD.n1877 GND 0.260855f
C2839 VDD.n1878 GND 0.004398f
C2840 VDD.n1879 GND 0.009619f
C2841 VDD.n1880 GND 0.010235f
C2842 VDD.n1881 GND 0.009686f
C2843 VDD.n1882 GND 0.003686f
C2844 VDD.n1883 GND 0.004398f
C2845 VDD.n1884 GND 0.004398f
C2846 VDD.n1885 GND 0.00291f
C2847 VDD.n1886 GND 0.004398f
C2848 VDD.n1887 GND 0.004398f
C2849 VDD.n1888 GND 0.004398f
C2850 VDD.n1889 GND 0.004398f
C2851 VDD.n1890 GND 0.004398f
C2852 VDD.n1891 GND 0.004398f
C2853 VDD.n1892 GND 0.004398f
C2854 VDD.n1893 GND 0.004398f
C2855 VDD.n1894 GND 0.004398f
C2856 VDD.n1895 GND 0.004398f
C2857 VDD.n1896 GND 0.004398f
C2858 VDD.n1897 GND 0.004398f
C2859 VDD.n1898 GND 0.004398f
C2860 VDD.n1899 GND 0.004398f
C2861 VDD.n1900 GND 0.004398f
C2862 VDD.n1901 GND 0.004398f
C2863 VDD.n1902 GND 0.004398f
C2864 VDD.n1903 GND 0.004398f
C2865 VDD.n1904 GND 0.004398f
C2866 VDD.n1905 GND 0.004398f
C2867 VDD.n1906 GND 0.004398f
C2868 VDD.n1907 GND 0.010235f
C2869 VDD.n1908 GND 0.010235f
C2870 VDD.n1909 GND 1.62651f
C2871 VDD.n1922 GND 0.004398f
C2872 VDD.n1923 GND 0.009619f
C2873 VDD.t63 GND 0.041419f
C2874 VDD.t64 GND 0.056208f
C2875 VDD.t62 GND 0.369485f
C2876 VDD.n1924 GND 0.058137f
C2877 VDD.n1925 GND 0.040639f
C2878 VDD.n1926 GND 0.004398f
C2879 VDD.n1927 GND 0.004398f
C2880 VDD.n1928 GND 0.004398f
C2881 VDD.n1929 GND 0.004398f
C2882 VDD.n1930 GND 0.004398f
C2883 VDD.n1931 GND 0.004398f
C2884 VDD.n1932 GND 0.004398f
C2885 VDD.n1933 GND 0.004398f
C2886 VDD.n1934 GND 0.004398f
C2887 VDD.n1935 GND 0.004398f
C2888 VDD.n1936 GND 0.004398f
C2889 VDD.n1937 GND 0.004398f
C2890 VDD.n1938 GND 0.004398f
C2891 VDD.n1939 GND 0.004398f
C2892 VDD.n1940 GND 0.004398f
C2893 VDD.n1941 GND 0.004398f
C2894 VDD.n1942 GND 0.004398f
C2895 VDD.n1943 GND 0.004398f
C2896 VDD.n1944 GND 0.004398f
C2897 VDD.n1945 GND 0.004398f
C2898 VDD.n1946 GND 0.004398f
C2899 VDD.n1947 GND 0.00291f
C2900 VDD.n1948 GND 0.006285f
C2901 VDD.n1949 GND 0.003686f
C2902 VDD.n1950 GND 0.004398f
C2903 VDD.n1951 GND 0.004398f
C2904 VDD.n1952 GND 0.004398f
C2905 VDD.n1953 GND 0.004398f
C2906 VDD.n1954 GND 0.004398f
C2907 VDD.n1955 GND 0.004398f
C2908 VDD.n1956 GND 0.004398f
C2909 VDD.n1957 GND 0.004398f
C2910 VDD.n1958 GND 0.004398f
C2911 VDD.n1959 GND 0.004398f
C2912 VDD.n1960 GND 0.004398f
C2913 VDD.n1961 GND 0.004398f
C2914 VDD.n1962 GND 0.004398f
C2915 VDD.n1963 GND 0.004398f
C2916 VDD.n1964 GND 0.004398f
C2917 VDD.n1965 GND 0.004398f
C2918 VDD.n1966 GND 0.004398f
C2919 VDD.n1967 GND 0.004398f
C2920 VDD.n1968 GND 0.004398f
C2921 VDD.n1969 GND 0.004398f
C2922 VDD.n1970 GND 0.004398f
C2923 VDD.n1971 GND 0.004398f
C2924 VDD.n1972 GND 0.004398f
C2925 VDD.n1973 GND 0.004398f
C2926 VDD.n1974 GND 0.004398f
C2927 VDD.n1975 GND 0.004398f
C2928 VDD.n1976 GND 0.004398f
C2929 VDD.n1977 GND 0.004398f
C2930 VDD.n1978 GND 0.004398f
C2931 VDD.n1979 GND 0.004398f
C2932 VDD.n1980 GND 0.004398f
C2933 VDD.n1981 GND 0.004398f
C2934 VDD.n1982 GND 0.004398f
C2935 VDD.n1983 GND 0.004398f
C2936 VDD.n1984 GND 0.004398f
C2937 VDD.n1985 GND 0.004398f
C2938 VDD.n1986 GND 0.004398f
C2939 VDD.n1987 GND 0.004398f
C2940 VDD.n1988 GND 0.004398f
C2941 VDD.n1989 GND 0.004398f
C2942 VDD.n1990 GND 0.004398f
C2943 VDD.n1991 GND 0.004398f
C2944 VDD.n1992 GND 0.004398f
C2945 VDD.n1993 GND 0.004398f
C2946 VDD.n1994 GND 0.004398f
C2947 VDD.n1995 GND 0.004398f
C2948 VDD.n1996 GND 0.004398f
C2949 VDD.n1997 GND 0.004398f
C2950 VDD.n1998 GND 0.004398f
C2951 VDD.n1999 GND 0.004398f
C2952 VDD.n2000 GND 0.004398f
C2953 VDD.n2001 GND 0.004398f
C2954 VDD.n2002 GND 0.004398f
C2955 VDD.n2003 GND 0.004398f
C2956 VDD.n2004 GND 0.004398f
C2957 VDD.n2005 GND 0.004398f
C2958 VDD.n2006 GND 0.004398f
C2959 VDD.n2007 GND 0.004398f
C2960 VDD.n2008 GND 0.004398f
C2961 VDD.n2009 GND 0.004398f
C2962 VDD.n2010 GND 0.004398f
C2963 VDD.n2011 GND 0.004398f
C2964 VDD.n2012 GND 0.004398f
C2965 VDD.n2013 GND 0.004398f
C2966 VDD.n2014 GND 0.004398f
C2967 VDD.n2015 GND 0.004398f
C2968 VDD.n2016 GND 0.004398f
C2969 VDD.n2017 GND 0.004398f
C2970 VDD.n2018 GND 0.004398f
C2971 VDD.n2019 GND 0.004398f
C2972 VDD.n2020 GND 0.004398f
C2973 VDD.n2021 GND 0.004398f
C2974 VDD.n2022 GND 0.004398f
C2975 VDD.n2023 GND 0.004398f
C2976 VDD.n2024 GND 0.004398f
C2977 VDD.n2025 GND 0.004398f
C2978 VDD.n2026 GND 0.004398f
C2979 VDD.n2027 GND 0.004398f
C2980 VDD.n2028 GND 0.004398f
C2981 VDD.n2029 GND 0.004398f
C2982 VDD.n2030 GND 0.004398f
C2983 VDD.n2031 GND 0.004398f
C2984 VDD.n2032 GND 0.004398f
C2985 VDD.n2033 GND 0.004398f
C2986 VDD.n2034 GND 0.004398f
C2987 VDD.n2035 GND 0.004398f
C2988 VDD.n2036 GND 0.004398f
C2989 VDD.n2037 GND 0.004398f
C2990 VDD.n2038 GND 0.004398f
C2991 VDD.n2039 GND 0.004398f
C2992 VDD.n2040 GND 0.004398f
C2993 VDD.n2041 GND 0.004398f
C2994 VDD.n2042 GND 0.004398f
C2995 VDD.n2043 GND 0.004398f
C2996 VDD.n2044 GND 0.004398f
C2997 VDD.n2045 GND 0.004398f
C2998 VDD.n2046 GND 0.004398f
C2999 VDD.n2047 GND 0.004398f
C3000 VDD.n2048 GND 0.004398f
C3001 VDD.n2049 GND 0.004398f
C3002 VDD.n2050 GND 0.004398f
C3003 VDD.n2051 GND 0.004398f
C3004 VDD.n2052 GND 0.004398f
C3005 VDD.n2053 GND 0.004398f
C3006 VDD.n2054 GND 0.004398f
C3007 VDD.n2055 GND 0.004398f
C3008 VDD.n2056 GND 0.004398f
C3009 VDD.n2057 GND 0.004398f
C3010 VDD.n2058 GND 0.004398f
C3011 VDD.n2059 GND 0.004398f
C3012 VDD.n2060 GND 0.004398f
C3013 VDD.n2061 GND 0.004398f
C3014 VDD.n2062 GND 0.004398f
C3015 VDD.n2063 GND 0.004398f
C3016 VDD.n2064 GND 0.004398f
C3017 VDD.n2065 GND 0.004398f
C3018 VDD.n2066 GND 0.004398f
C3019 VDD.n2067 GND 0.004398f
C3020 VDD.n2068 GND 0.004398f
C3021 VDD.n2069 GND 0.004398f
C3022 VDD.n2070 GND 0.004398f
C3023 VDD.n2071 GND 0.004398f
C3024 VDD.n2072 GND 0.004398f
C3025 VDD.n2073 GND 0.004398f
C3026 VDD.n2074 GND 0.004398f
C3027 VDD.n2075 GND 0.004398f
C3028 VDD.n2076 GND 0.004398f
C3029 VDD.n2077 GND 0.004398f
C3030 VDD.n2078 GND 0.004398f
C3031 VDD.n2079 GND 0.004398f
C3032 VDD.n2080 GND 0.009619f
C3033 VDD.n2081 GND 0.010235f
C3034 VDD.n2082 GND 0.010235f
C3035 VDD.n2083 GND 0.004398f
C3036 VDD.n2084 GND 0.004398f
C3037 VDD.t60 GND 0.041419f
C3038 VDD.t61 GND 0.056208f
C3039 VDD.t58 GND 0.369485f
C3040 VDD.n2085 GND 0.058137f
C3041 VDD.n2086 GND 0.040639f
C3042 VDD.n2087 GND 0.006285f
C3043 VDD.n2088 GND 0.004398f
C3044 VDD.n2089 GND 0.004398f
C3045 VDD.n2090 GND 0.004398f
C3046 VDD.n2091 GND 0.004398f
C3047 VDD.n2092 GND 0.004398f
C3048 VDD.n2093 GND 0.004398f
C3049 VDD.n2094 GND 0.004398f
C3050 VDD.n2095 GND 0.004398f
C3051 VDD.n2096 GND 0.004398f
C3052 VDD.n2097 GND 0.004398f
C3053 VDD.n2098 GND 0.004398f
C3054 VDD.n2099 GND 0.004398f
C3055 VDD.n2100 GND 0.004398f
C3056 VDD.n2101 GND 0.004398f
C3057 VDD.n2102 GND 0.004398f
C3058 VDD.n2103 GND 0.004398f
C3059 VDD.n2104 GND 0.004398f
C3060 VDD.n2105 GND 0.004398f
C3061 VDD.n2106 GND 0.004398f
C3062 VDD.n2107 GND 0.004398f
C3063 VDD.n2108 GND 0.004398f
C3064 VDD.n2109 GND 0.004398f
C3065 VDD.n2110 GND 0.004398f
C3066 VDD.n2111 GND 0.004398f
C3067 VDD.n2112 GND 0.004398f
C3068 VDD.n2113 GND 0.004398f
C3069 VDD.n2114 GND 0.004398f
C3070 VDD.n2115 GND 0.004398f
C3071 VDD.n2116 GND 0.004398f
C3072 VDD.n2117 GND 0.004398f
C3073 VDD.n2118 GND 0.004398f
C3074 VDD.n2119 GND 0.004398f
C3075 VDD.n2120 GND 0.004398f
C3076 VDD.n2121 GND 0.004398f
C3077 VDD.n2122 GND 0.004398f
C3078 VDD.n2123 GND 0.004398f
C3079 VDD.n2124 GND 0.004398f
C3080 VDD.n2125 GND 0.004398f
C3081 VDD.n2126 GND 0.004398f
C3082 VDD.n2127 GND 0.004398f
C3083 VDD.n2128 GND 0.004398f
C3084 VDD.n2129 GND 0.004398f
C3085 VDD.n2130 GND 0.004398f
C3086 VDD.n2131 GND 0.004398f
C3087 VDD.n2132 GND 0.004398f
C3088 VDD.n2133 GND 0.004398f
C3089 VDD.n2134 GND 0.004398f
C3090 VDD.n2135 GND 0.004398f
C3091 VDD.n2136 GND 0.004398f
C3092 VDD.n2137 GND 0.004398f
C3093 VDD.n2138 GND 0.004398f
C3094 VDD.n2139 GND 0.004398f
C3095 VDD.n2140 GND 0.004398f
C3096 VDD.n2141 GND 0.004398f
C3097 VDD.n2142 GND 0.004398f
C3098 VDD.n2143 GND 0.004398f
C3099 VDD.n2144 GND 0.004398f
C3100 VDD.n2145 GND 0.004398f
C3101 VDD.n2146 GND 0.004398f
C3102 VDD.n2147 GND 0.004398f
C3103 VDD.n2148 GND 0.004398f
C3104 VDD.n2149 GND 0.004398f
C3105 VDD.n2150 GND 0.004398f
C3106 VDD.n2151 GND 0.004398f
C3107 VDD.n2152 GND 0.004398f
C3108 VDD.n2153 GND 0.004398f
C3109 VDD.n2154 GND 0.004398f
C3110 VDD.n2155 GND 0.004398f
C3111 VDD.n2156 GND 0.004398f
C3112 VDD.n2157 GND 0.004398f
C3113 VDD.n2158 GND 0.004398f
C3114 VDD.n2159 GND 0.004398f
C3115 VDD.n2160 GND 0.004398f
C3116 VDD.n2161 GND 0.004398f
C3117 VDD.n2162 GND 0.004398f
C3118 VDD.n2163 GND 0.004398f
C3119 VDD.n2164 GND 0.004398f
C3120 VDD.n2165 GND 0.004398f
C3121 VDD.n2166 GND 0.004398f
C3122 VDD.n2167 GND 0.004398f
C3123 VDD.n2168 GND 0.004398f
C3124 VDD.n2169 GND 0.004398f
C3125 VDD.n2170 GND 0.004398f
C3126 VDD.n2171 GND 0.004398f
C3127 VDD.n2172 GND 0.004398f
C3128 VDD.n2173 GND 0.004398f
C3129 VDD.n2174 GND 0.004398f
C3130 VDD.n2175 GND 0.004398f
C3131 VDD.n2176 GND 0.004398f
C3132 VDD.n2177 GND 0.004398f
C3133 VDD.n2178 GND 0.004398f
C3134 VDD.n2179 GND 0.004398f
C3135 VDD.n2180 GND 0.004398f
C3136 VDD.n2181 GND 0.004398f
C3137 VDD.n2182 GND 0.004398f
C3138 VDD.n2183 GND 0.004398f
C3139 VDD.n2184 GND 0.004398f
C3140 VDD.n2185 GND 0.004398f
C3141 VDD.n2186 GND 0.004398f
C3142 VDD.n2187 GND 0.004398f
C3143 VDD.n2188 GND 0.004398f
C3144 VDD.n2189 GND 0.004398f
C3145 VDD.n2190 GND 0.004398f
C3146 VDD.n2191 GND 0.004398f
C3147 VDD.n2192 GND 0.004398f
C3148 VDD.n2193 GND 0.004398f
C3149 VDD.n2194 GND 0.004398f
C3150 VDD.n2195 GND 0.004398f
C3151 VDD.n2196 GND 0.004398f
C3152 VDD.n2197 GND 0.004398f
C3153 VDD.n2198 GND 0.004398f
C3154 VDD.n2199 GND 0.004398f
C3155 VDD.n2200 GND 0.004398f
C3156 VDD.n2201 GND 0.004398f
C3157 VDD.n2202 GND 0.004398f
C3158 VDD.n2203 GND 0.004398f
C3159 VDD.n2204 GND 0.004398f
C3160 VDD.n2205 GND 0.004398f
C3161 VDD.n2206 GND 0.004398f
C3162 VDD.n2207 GND 0.004398f
C3163 VDD.n2208 GND 0.004398f
C3164 VDD.n2209 GND 0.004398f
C3165 VDD.n2210 GND 0.004398f
C3166 VDD.n2211 GND 0.004398f
C3167 VDD.n2212 GND 0.004398f
C3168 VDD.n2213 GND 0.004398f
C3169 VDD.n2214 GND 0.004398f
C3170 VDD.n2215 GND 0.004398f
C3171 VDD.n2216 GND 0.009619f
C3172 VDD.n2217 GND 0.009619f
C3173 VDD.n2218 GND 0.010235f
C3174 VDD.n2219 GND 0.010235f
C3175 VDD.n2220 GND 0.003686f
C3176 VDD.n2221 GND 0.004398f
C3177 VDD.n2222 GND 0.004398f
C3178 VDD.n2223 GND 0.00291f
C3179 VDD.n2224 GND 0.004398f
C3180 VDD.n2225 GND 0.004398f
C3181 VDD.n2226 GND 0.004398f
C3182 VDD.n2227 GND 0.004398f
C3183 VDD.n2228 GND 0.004398f
C3184 VDD.n2229 GND 0.004398f
C3185 VDD.n2230 GND 0.004398f
C3186 VDD.n2231 GND 0.004398f
C3187 VDD.n2232 GND 0.004398f
C3188 VDD.n2233 GND 0.004398f
C3189 VDD.n2234 GND 0.004398f
C3190 VDD.n2235 GND 0.004398f
C3191 VDD.n2236 GND 0.004398f
C3192 VDD.n2237 GND 0.004398f
C3193 VDD.n2238 GND 0.004398f
C3194 VDD.n2239 GND 0.004398f
C3195 VDD.n2240 GND 0.004398f
C3196 VDD.n2241 GND 0.004398f
C3197 VDD.n2242 GND 0.004398f
C3198 VDD.n2243 GND 0.004398f
C3199 VDD.n2244 GND 0.010235f
C3200 VDD.n2245 GND 0.010235f
C3201 VDD.n2247 GND 1.62651f
C3202 VDD.n2249 GND 0.010235f
C3203 VDD.n2250 GND 0.010235f
C3204 VDD.n2251 GND 0.009619f
C3205 VDD.n2252 GND 0.004398f
C3206 VDD.n2253 GND 0.004398f
C3207 VDD.n2254 GND 0.260855f
C3208 VDD.n2255 GND 0.004398f
C3209 VDD.n2256 GND 0.004398f
C3210 VDD.n2257 GND 0.004398f
C3211 VDD.n2258 GND 0.004398f
C3212 VDD.n2259 GND 0.004398f
C3213 VDD.n2260 GND 0.260855f
C3214 VDD.n2261 GND 0.004398f
C3215 VDD.n2262 GND 0.004398f
C3216 VDD.n2263 GND 0.004398f
C3217 VDD.n2264 GND 0.004398f
C3218 VDD.n2265 GND 0.004398f
C3219 VDD.n2266 GND 0.260855f
C3220 VDD.n2267 GND 0.004398f
C3221 VDD.n2268 GND 0.004398f
C3222 VDD.n2269 GND 0.004398f
C3223 VDD.n2270 GND 0.004398f
C3224 VDD.n2271 GND 0.004398f
C3225 VDD.n2272 GND 0.168789f
C3226 VDD.n2273 GND 0.004398f
C3227 VDD.n2274 GND 0.004398f
C3228 VDD.n2275 GND 0.004398f
C3229 VDD.n2276 GND 0.004398f
C3230 VDD.n2277 GND 0.004398f
C3231 VDD.n2278 GND 0.260855f
C3232 VDD.n2279 GND 0.004398f
C3233 VDD.n2280 GND 0.004398f
C3234 VDD.n2281 GND 0.004398f
C3235 VDD.n2282 GND 0.004398f
C3236 VDD.n2283 GND 0.004398f
C3237 VDD.n2284 GND 0.260855f
C3238 VDD.n2285 GND 0.004398f
C3239 VDD.n2286 GND 0.004398f
C3240 VDD.n2287 GND 0.004398f
C3241 VDD.n2288 GND 0.004398f
C3242 VDD.n2289 GND 0.004398f
C3243 VDD.n2290 GND 0.260855f
C3244 VDD.n2291 GND 0.004398f
C3245 VDD.n2292 GND 0.004398f
C3246 VDD.n2293 GND 0.004398f
C3247 VDD.n2294 GND 0.004398f
C3248 VDD.n2295 GND 0.004398f
C3249 VDD.n2296 GND 0.260855f
C3250 VDD.n2297 GND 0.004398f
C3251 VDD.n2298 GND 0.004398f
C3252 VDD.n2299 GND 0.004398f
C3253 VDD.n2300 GND 0.004398f
C3254 VDD.n2301 GND 0.004398f
C3255 VDD.n2302 GND 0.260855f
C3256 VDD.n2303 GND 0.004398f
C3257 VDD.n2304 GND 0.004398f
C3258 VDD.n2305 GND 0.004398f
C3259 VDD.n2306 GND 0.004398f
C3260 VDD.n2307 GND 0.004398f
C3261 VDD.n2308 GND 0.260855f
C3262 VDD.n2309 GND 0.004398f
C3263 VDD.n2310 GND 0.004398f
C3264 VDD.n2311 GND 0.004398f
C3265 VDD.n2312 GND 0.004398f
C3266 VDD.n2313 GND 0.004398f
C3267 VDD.n2314 GND 0.149608f
C3268 VDD.n2315 GND 0.004398f
C3269 VDD.n2316 GND 0.004398f
C3270 VDD.n2317 GND 0.004398f
C3271 VDD.n2318 GND 0.004398f
C3272 VDD.n2319 GND 0.004398f
C3273 VDD.n2320 GND 0.260855f
C3274 VDD.n2321 GND 0.004398f
C3275 VDD.n2322 GND 0.004398f
C3276 VDD.n2323 GND 0.004398f
C3277 VDD.n2324 GND 0.004398f
C3278 VDD.n2325 GND 0.004398f
C3279 VDD.n2326 GND 0.174543f
C3280 VDD.n2327 GND 0.004398f
C3281 VDD.n2328 GND 0.004398f
C3282 VDD.n2329 GND 0.004398f
C3283 VDD.n2330 GND 0.004398f
C3284 VDD.n2331 GND 0.004398f
C3285 VDD.n2332 GND 0.260855f
C3286 VDD.n2333 GND 0.004398f
C3287 VDD.n2334 GND 0.004398f
C3288 VDD.n2335 GND 0.004398f
C3289 VDD.n2336 GND 0.004398f
C3290 VDD.n2337 GND 0.004398f
C3291 VDD.n2338 GND 0.260855f
C3292 VDD.n2339 GND 0.004398f
C3293 VDD.n2340 GND 0.004398f
C3294 VDD.n2341 GND 0.004398f
C3295 VDD.n2342 GND 0.004398f
C3296 VDD.n2343 GND 0.004398f
C3297 VDD.n2344 GND 0.260855f
C3298 VDD.n2345 GND 0.004398f
C3299 VDD.n2346 GND 0.004398f
C3300 VDD.n2347 GND 0.004398f
C3301 VDD.n2348 GND 0.004398f
C3302 VDD.n2349 GND 0.004398f
C3303 VDD.n2350 GND 0.260855f
C3304 VDD.n2351 GND 0.004398f
C3305 VDD.n2352 GND 0.004398f
C3306 VDD.n2353 GND 0.004398f
C3307 VDD.n2354 GND 0.004398f
C3308 VDD.n2355 GND 0.004398f
C3309 VDD.n2356 GND 0.20715f
C3310 VDD.n2357 GND 0.004398f
C3311 VDD.n2358 GND 0.004398f
C3312 VDD.n2359 GND 0.004398f
C3313 VDD.n2360 GND 0.004398f
C3314 VDD.n2361 GND 0.004398f
C3315 VDD.n2362 GND 0.260855f
C3316 VDD.n2363 GND 0.004398f
C3317 VDD.n2364 GND 0.004398f
C3318 VDD.n2365 GND 0.004398f
C3319 VDD.n2366 GND 0.004398f
C3320 VDD.n2367 GND 0.004398f
C3321 VDD.n2368 GND 0.232084f
C3322 VDD.n2369 GND 0.004398f
C3323 VDD.n2370 GND 0.004398f
C3324 VDD.n2371 GND 0.004398f
C3325 VDD.n2372 GND 0.004398f
C3326 VDD.n2373 GND 0.004398f
C3327 VDD.n2374 GND 0.260855f
C3328 VDD.n2375 GND 0.004398f
C3329 VDD.n2376 GND 0.004398f
C3330 VDD.n2377 GND 0.004398f
C3331 VDD.n2378 GND 0.004398f
C3332 VDD.n2379 GND 0.004398f
C3333 VDD.n2380 GND 0.260855f
C3334 VDD.n2381 GND 0.004398f
C3335 VDD.n2382 GND 0.004398f
C3336 VDD.n2383 GND 0.004398f
C3337 VDD.n2384 GND 0.004398f
C3338 VDD.n2385 GND 0.004398f
C3339 VDD.n2386 GND 0.260855f
C3340 VDD.n2387 GND 0.004398f
C3341 VDD.n2388 GND 0.004398f
C3342 VDD.n2389 GND 0.004398f
C3343 VDD.n2390 GND 0.004398f
C3344 VDD.n2391 GND 0.004398f
C3345 VDD.n2392 GND 0.257019f
C3346 VDD.n2393 GND 0.004398f
C3347 VDD.n2394 GND 0.004398f
C3348 VDD.n2395 GND 0.004398f
C3349 VDD.n2396 GND 0.004398f
C3350 VDD.n2397 GND 0.004398f
C3351 VDD.n2398 GND 0.260855f
C3352 VDD.n2399 GND 0.004398f
C3353 VDD.n2400 GND 0.004398f
C3354 VDD.n2401 GND 0.004398f
C3355 VDD.n2402 GND 0.004398f
C3356 VDD.n2403 GND 0.004398f
C3357 VDD.n2404 GND 0.232084f
C3358 VDD.n2405 GND 0.004398f
C3359 VDD.n2406 GND 0.004398f
C3360 VDD.n2407 GND 0.004398f
C3361 VDD.n2408 GND 0.004398f
C3362 VDD.n2409 GND 0.004398f
C3363 VDD.n2410 GND 0.260855f
C3364 VDD.n2411 GND 0.004398f
C3365 VDD.n2412 GND 0.004398f
C3366 VDD.n2413 GND 0.004398f
C3367 VDD.n2414 GND 0.004398f
C3368 VDD.n2415 GND 0.004398f
C3369 VDD.n2416 GND 0.260855f
C3370 VDD.n2417 GND 0.004398f
C3371 VDD.n2418 GND 0.004398f
C3372 VDD.n2419 GND 0.004398f
C3373 VDD.n2420 GND 0.004398f
C3374 VDD.n2421 GND 0.004398f
C3375 VDD.n2422 GND 0.260855f
C3376 VDD.n2423 GND 0.004398f
C3377 VDD.n2424 GND 0.004398f
C3378 VDD.n2425 GND 0.004398f
C3379 VDD.n2426 GND 0.004398f
C3380 VDD.n2427 GND 0.004398f
C3381 VDD.n2428 GND 0.260855f
C3382 VDD.n2429 GND 0.004398f
C3383 VDD.n2430 GND 0.004398f
C3384 VDD.n2431 GND 0.004398f
C3385 VDD.n2432 GND 0.004398f
C3386 VDD.n2433 GND 0.004398f
C3387 VDD.n2434 GND 0.260855f
C3388 VDD.n2435 GND 0.004398f
C3389 VDD.n2436 GND 0.004398f
C3390 VDD.n2437 GND 0.004398f
C3391 VDD.n2438 GND 0.004398f
C3392 VDD.n2439 GND 0.004398f
C3393 VDD.n2440 GND 0.260855f
C3394 VDD.n2441 GND 0.004398f
C3395 VDD.n2442 GND 0.004398f
C3396 VDD.n2443 GND 0.004398f
C3397 VDD.n2444 GND 0.004398f
C3398 VDD.n2445 GND 0.004398f
C3399 VDD.n2446 GND 0.174543f
C3400 VDD.n2447 GND 0.004398f
C3401 VDD.n2448 GND 0.004398f
C3402 VDD.n2449 GND 0.004398f
C3403 VDD.n2450 GND 0.004398f
C3404 VDD.n2451 GND 0.004398f
C3405 VDD.n2452 GND 0.260855f
C3406 VDD.n2453 GND 0.004398f
C3407 VDD.n2454 GND 0.004398f
C3408 VDD.n2455 GND 0.004398f
C3409 VDD.n2456 GND 0.004398f
C3410 VDD.n2457 GND 0.004398f
C3411 VDD.n2458 GND 0.199477f
C3412 VDD.n2459 GND 0.004398f
C3413 VDD.n2460 GND 0.004398f
C3414 VDD.n2461 GND 0.004398f
C3415 VDD.n2462 GND 0.004398f
C3416 VDD.n2463 GND 0.004398f
C3417 VDD.n2464 GND 0.260855f
C3418 VDD.n2465 GND 0.004398f
C3419 VDD.n2466 GND 0.004398f
C3420 VDD.n2467 GND 0.004398f
C3421 VDD.n2468 GND 0.004398f
C3422 VDD.n2469 GND 0.004398f
C3423 VDD.n2470 GND 0.260855f
C3424 VDD.n2471 GND 0.004398f
C3425 VDD.n2472 GND 0.004398f
C3426 VDD.n2473 GND 0.004398f
C3427 VDD.n2474 GND 0.004398f
C3428 VDD.n2475 GND 0.004398f
C3429 VDD.n2476 GND 0.260855f
C3430 VDD.n2477 GND 0.004398f
C3431 VDD.n2478 GND 0.004398f
C3432 VDD.n2479 GND 0.004398f
C3433 VDD.n2480 GND 0.004398f
C3434 VDD.n2481 GND 0.004398f
C3435 VDD.n2482 GND 0.260855f
C3436 VDD.n2483 GND 0.004398f
C3437 VDD.n2484 GND 0.004398f
C3438 VDD.n2485 GND 0.004398f
C3439 VDD.n2486 GND 0.004398f
C3440 VDD.n2487 GND 0.004398f
C3441 VDD.n2488 GND 0.260855f
C3442 VDD.n2489 GND 0.004398f
C3443 VDD.n2490 GND 0.004398f
C3444 VDD.n2491 GND 0.004398f
C3445 VDD.n2492 GND 0.004398f
C3446 VDD.n2493 GND 0.004398f
C3447 VDD.n2494 GND 0.260855f
C3448 VDD.n2495 GND 0.004398f
C3449 VDD.n2496 GND 0.004398f
C3450 VDD.n2497 GND 0.004398f
C3451 VDD.n2498 GND 0.004398f
C3452 VDD.n2499 GND 0.004398f
C3453 VDD.n2500 GND 0.247429f
C3454 VDD.n2501 GND 0.004398f
C3455 VDD.n2502 GND 0.004398f
C3456 VDD.n2503 GND 0.004398f
C3457 VDD.n2504 GND 0.010235f
C3458 VDD.n2505 GND 0.004398f
C3459 VDD.n2506 GND 0.004398f
C3460 VDD.n2507 GND 0.004398f
C3461 VDD.n2510 GND 0.004398f
C3462 VDD.n2511 GND 0.004398f
C3463 VDD.n2512 GND 0.004398f
C3464 VDD.n2513 GND 0.004398f
C3465 VDD.n2514 GND 0.004398f
C3466 VDD.n2515 GND 0.004398f
C3467 VDD.n2517 GND 0.004398f
C3468 VDD.n2518 GND 0.010235f
C3469 VDD.n2519 GND 0.009619f
C3470 VDD.n2520 GND 0.009619f
C3471 VDD.n2521 GND 0.004398f
C3472 VDD.n2522 GND 0.004398f
C3473 VDD.n2523 GND 0.004398f
C3474 VDD.n2524 GND 0.004398f
C3475 VDD.n2525 GND 0.004398f
C3476 VDD.n2526 GND 0.004398f
C3477 VDD.n2527 GND 0.004398f
C3478 VDD.n2528 GND 0.260855f
C3479 VDD.n2529 GND 0.004398f
C3480 VDD.n2530 GND 0.004398f
C3481 VDD.n2531 GND 0.004398f
C3482 VDD.n2532 GND 0.004398f
C3483 VDD.n2533 GND 0.004398f
C3484 VDD.n2534 GND 0.260855f
C3485 VDD.n2535 GND 0.004398f
C3486 VDD.n2536 GND 0.004398f
C3487 VDD.n2537 GND 0.004398f
C3488 VDD.n2538 GND 0.004398f
C3489 VDD.n2539 GND 0.010168f
C3490 VDD.n2540 GND 0.009686f
C3491 VDD.n2541 GND 0.010235f
C3492 VDD.n2543 GND 0.004398f
C3493 VDD.n2544 GND 0.004398f
C3494 VDD.n2545 GND 0.00291f
C3495 VDD.n2546 GND 0.004398f
C3496 VDD.n2547 GND 0.004398f
C3497 VDD.n2548 GND 0.004398f
C3498 VDD.n2550 GND 0.004398f
C3499 VDD.n2551 GND 0.004398f
C3500 VDD.n2552 GND 0.004398f
C3501 VDD.n2553 GND 1.08695f
C3502 VDD.n2554 GND 0.063945f
C3503 VDD.n2555 GND 0.004398f
C3504 VDD.n2556 GND 0.004398f
C3505 VDD.n2558 GND 0.004398f
C3506 VDD.n2559 GND 0.004398f
C3507 VDD.n2560 GND 0.004398f
C3508 VDD.n2561 GND 0.004398f
C3509 VDD.n2562 GND 0.004398f
C3510 VDD.n2563 GND 0.004398f
C3511 VDD.n2565 GND 0.004398f
C3512 VDD.n2566 GND 0.010235f
C3513 VDD.n2567 GND 0.010235f
C3514 VDD.n2568 GND 0.009619f
C3515 VDD.n2569 GND 0.004398f
C3516 VDD.n2570 GND 0.004398f
C3517 VDD.n2571 GND 0.260855f
C3518 VDD.n2572 GND 0.004398f
C3519 VDD.n2573 GND 0.004398f
C3520 VDD.n2574 GND 0.010168f
C3521 VDD.n2575 GND 0.009686f
C3522 VDD.n2576 GND 0.010235f
C3523 VDD.n2578 GND 0.004398f
C3524 VDD.n2579 GND 0.004398f
C3525 VDD.n2580 GND 0.00291f
C3526 VDD.n2581 GND 0.004398f
C3527 VDD.n2582 GND 0.004398f
C3528 VDD.n2583 GND 0.004398f
C3529 VDD.n2585 GND 0.004398f
C3530 VDD.n2586 GND 0.004398f
C3531 VDD.n2588 GND 0.004398f
C3532 VDD.n2589 GND 0.063945f
C3533 VDD.n2590 GND 0.006467f
C3534 VDD.n2591 GND 0.006467f
C3535 VDD.n2592 GND 0.005205f
C3536 VDD.n2593 GND 0.006467f
C3537 VDD.n2594 GND 0.006467f
C3538 VDD.n2595 GND 0.006467f
C3539 VDD.n2596 GND 0.006467f
C3540 VDD.n2597 GND 0.002733f
C3541 VDD.n2598 GND 0.006467f
C3542 VDD.n2599 GND 0.005205f
C3543 VDD.n2600 GND 0.005205f
C3544 VDD.n2601 GND 0.006467f
C3545 VDD.n2602 GND 0.006467f
C3546 VDD.n2603 GND 0.005205f
C3547 VDD.n2604 GND 0.006467f
C3548 VDD.n2605 GND 0.005205f
C3549 VDD.n2606 GND 0.005205f
C3550 VDD.n2608 GND 1.08695f
C3551 VDD.n2610 GND 0.005205f
C3552 VDD.n2611 GND 0.006467f
C3553 VDD.n2612 GND 0.006467f
C3554 VDD.n2613 GND 0.005205f
C3555 VDD.n2614 GND 0.005205f
C3556 VDD.n2615 GND 0.006467f
C3557 VDD.n2616 GND 0.006467f
C3558 VDD.n2617 GND 0.005205f
C3559 VDD.n2618 GND 0.006467f
C3560 VDD.n2619 GND 0.006467f
C3561 VDD.n2620 GND 0.005205f
C3562 VDD.n2621 GND 0.006467f
C3563 VDD.n2622 GND 0.006467f
C3564 VDD.n2623 GND 0.006467f
C3565 VDD.n2624 GND 0.010619f
C3566 VDD.n2625 GND 0.006467f
C3567 VDD.n2626 GND 0.006467f
C3568 VDD.n2627 GND 0.00354f
C3569 VDD.n2628 GND 0.005205f
C3570 VDD.n2629 GND 0.006467f
C3571 VDD.n2630 GND 0.006467f
C3572 VDD.n2631 GND 0.005205f
C3573 VDD.n2632 GND 0.005205f
C3574 VDD.n2633 GND 0.006467f
C3575 VDD.n2634 GND 0.006467f
C3576 VDD.n2635 GND 0.005205f
C3577 VDD.n2636 GND 0.005205f
C3578 VDD.n2637 GND 0.006467f
C3579 VDD.n2638 GND 0.006467f
C3580 VDD.n2639 GND 0.005205f
C3581 VDD.n2640 GND 0.005205f
C3582 VDD.n2641 GND 0.006467f
C3583 VDD.n2642 GND 0.006467f
C3584 VDD.n2643 GND 0.005205f
C3585 VDD.n2644 GND 0.005205f
C3586 VDD.n2645 GND 0.006467f
C3587 VDD.n2646 GND 0.006467f
C3588 VDD.n2647 GND 0.005205f
C3589 VDD.n2648 GND 0.005205f
C3590 VDD.n2649 GND 0.006467f
C3591 VDD.n2650 GND 0.006467f
C3592 VDD.n2651 GND 0.005205f
C3593 VDD.n2652 GND 0.006467f
C3594 VDD.n2653 GND 0.006467f
C3595 VDD.n2654 GND 0.006467f
C3596 VDD.t9 GND 0.089332f
C3597 VDD.t10 GND 0.10348f
C3598 VDD.t7 GND 0.482813f
C3599 VDD.n2655 GND 0.068834f
C3600 VDD.n2656 GND 0.04271f
C3601 VDD.n2657 GND 0.010619f
C3602 VDD.n2658 GND 0.004346f
C3603 VDD.n2659 GND 0.006467f
C3604 VDD.n2660 GND 0.006467f
C3605 VDD.n2661 GND 0.005205f
C3606 VDD.n2662 GND 0.005205f
C3607 VDD.n2663 GND 0.006467f
C3608 VDD.n2664 GND 0.006467f
C3609 VDD.n2665 GND 0.005205f
C3610 VDD.n2666 GND 0.005205f
C3611 VDD.n2667 GND 0.006467f
C3612 VDD.n2668 GND 0.006467f
C3613 VDD.n2669 GND 0.005205f
C3614 VDD.n2670 GND 0.005205f
C3615 VDD.n2671 GND 0.006467f
C3616 VDD.n2672 GND 0.006467f
C3617 VDD.n2673 GND 0.005205f
C3618 VDD.n2674 GND 0.006467f
C3619 VDD.n2675 GND 0.005205f
C3620 VDD.n2676 GND 0.005205f
C3621 VDD.n2677 GND 0.005205f
C3622 VDD.n2678 GND 0.00432f
C3623 VDD.n2679 GND 0.014463f
C3624 VDD.n2681 GND 2.79652f
C3625 VDD.n2683 GND 0.014463f
C3626 VDD.n2684 GND 0.002472f
C3627 VDD.n2685 GND 0.014463f
C3628 VDD.n2686 GND 0.014445f
C3629 VDD.n2687 GND 0.006467f
C3630 VDD.n2688 GND 0.005205f
C3631 VDD.n2689 GND 0.006467f
C3632 VDD.n2690 GND 0.38361f
C3633 VDD.n2691 GND 0.006467f
C3634 VDD.n2692 GND 0.005205f
C3635 VDD.n2693 GND 0.006467f
C3636 VDD.n2694 GND 0.006467f
C3637 VDD.n2695 GND 0.006467f
C3638 VDD.n2696 GND 0.005205f
C3639 VDD.n2697 GND 0.006467f
C3640 VDD.n2698 GND 0.356758f
C3641 VDD.n2699 GND 0.006467f
C3642 VDD.n2700 GND 0.005205f
C3643 VDD.n2701 GND 0.006467f
C3644 VDD.n2702 GND 0.006467f
C3645 VDD.n2703 GND 0.006467f
C3646 VDD.n2704 GND 0.005205f
C3647 VDD.n2705 GND 0.006467f
C3648 VDD.n2706 GND 0.38361f
C3649 VDD.n2707 GND 0.006467f
C3650 VDD.n2708 GND 0.005205f
C3651 VDD.n2709 GND 0.006467f
C3652 VDD.n2710 GND 0.006467f
C3653 VDD.n2711 GND 0.006467f
C3654 VDD.n2712 GND 0.005205f
C3655 VDD.n2713 GND 0.006467f
C3656 VDD.n2714 GND 0.38361f
C3657 VDD.n2715 GND 0.006467f
C3658 VDD.n2716 GND 0.005205f
C3659 VDD.n2717 GND 0.006467f
C3660 VDD.n2718 GND 0.006467f
C3661 VDD.n2719 GND 0.006467f
C3662 VDD.n2720 GND 0.005205f
C3663 VDD.n2721 GND 0.006467f
C3664 VDD.n2722 GND 0.38361f
C3665 VDD.n2723 GND 0.006467f
C3666 VDD.n2724 GND 0.005205f
C3667 VDD.n2725 GND 0.006467f
C3668 VDD.n2726 GND 0.006467f
C3669 VDD.n2727 GND 0.006467f
C3670 VDD.n2728 GND 0.005205f
C3671 VDD.n2729 GND 0.006467f
C3672 VDD.n2730 GND 0.38361f
C3673 VDD.n2731 GND 0.006467f
C3674 VDD.n2732 GND 0.005205f
C3675 VDD.n2733 GND 0.006467f
C3676 VDD.n2734 GND 0.006467f
C3677 VDD.n2735 GND 0.006467f
C3678 VDD.n2736 GND 0.006467f
C3679 VDD.n2737 GND 0.006467f
C3680 VDD.n2738 GND 0.005205f
C3681 VDD.n2739 GND 0.006467f
C3682 VDD.n2740 GND 0.38361f
C3683 VDD.n2741 GND 0.006467f
C3684 VDD.n2742 GND 0.006467f
C3685 VDD.n2743 GND 0.006467f
C3686 VDD.n2744 GND 0.006467f
C3687 VDD.n2745 GND 0.005205f
C3688 VDD.n2746 GND 0.006467f
C3689 VDD.n2747 GND 0.006467f
C3690 VDD.n2748 GND 0.006467f
C3691 VDD.n2749 GND 0.006467f
C3692 VDD.n2750 GND 0.38361f
C3693 VDD.n2751 GND 0.006467f
C3694 VDD.n2752 GND 0.006467f
C3695 VDD.n2753 GND 0.006467f
C3696 VDD.n2754 GND 0.006467f
C3697 VDD.n2755 GND 0.006467f
C3698 VDD.n2756 GND 0.005205f
C3699 VDD.n2757 GND 0.006467f
C3700 VDD.n2758 GND 0.006467f
C3701 VDD.n2759 GND 0.006467f
C3702 VDD.n2760 GND 0.006467f
C3703 VDD.n2761 GND 0.38361f
C3704 VDD.n2762 GND 0.006467f
C3705 VDD.n2763 GND 0.006467f
C3706 VDD.n2764 GND 0.006467f
C3707 VDD.n2765 GND 0.006467f
C3708 VDD.n2766 GND 0.006467f
C3709 VDD.n2767 GND 0.00432f
C3710 VDD.n2768 GND 0.014445f
C3711 VDD.n2769 GND 0.006467f
C3712 VDD.n2770 GND 0.014445f
C3713 VDD.n2792 GND 0.006467f
C3714 VDD.n2793 GND 0.014445f
C3715 VDD.n2794 GND 0.014463f
C3716 VDD.n2795 GND 0.005205f
C3717 VDD.n2796 GND 0.006467f
C3718 VDD.n2797 GND 0.006467f
C3719 VDD.n2798 GND 0.006467f
C3720 VDD.n2799 GND 0.006467f
C3721 VDD.n2800 GND 0.006467f
C3722 VDD.n2801 GND 0.006467f
C3723 VDD.n2802 GND 0.006467f
C3724 VDD.n2803 GND 0.006467f
C3725 VDD.n2804 GND 0.004346f
C3726 VDD.t14 GND 0.089332f
C3727 VDD.t13 GND 0.10348f
C3728 VDD.t11 GND 0.482813f
C3729 VDD.n2805 GND 0.068834f
C3730 VDD.n2806 GND 0.04271f
C3731 VDD.n2807 GND 0.006467f
C3732 VDD.n2808 GND 0.006467f
C3733 VDD.n2809 GND 0.006467f
C3734 VDD.n2810 GND 0.006467f
C3735 VDD.n2811 GND 0.006467f
C3736 VDD.n2812 GND 0.006467f
C3737 VDD.n2813 GND 0.006467f
C3738 VDD.n2814 GND 0.006467f
C3739 VDD.n2815 GND 0.006467f
C3740 VDD.n2816 GND 0.006467f
C3741 VDD.n2817 GND 0.006467f
C3742 VDD.n2818 GND 0.006467f
C3743 VDD.n2819 GND 0.006467f
C3744 VDD.n2820 GND 0.006467f
C3745 VDD.n2821 GND 0.005153f
C3746 VDD.t34 GND 0.089332f
C3747 VDD.t33 GND 0.10348f
C3748 VDD.t32 GND 0.482813f
C3749 VDD.n2822 GND 0.068834f
C3750 VDD.n2823 GND 0.04271f
C3751 VDD.n2824 GND 0.006467f
C3752 VDD.n2825 GND 0.006467f
C3753 VDD.n2826 GND 0.006467f
C3754 VDD.n2827 GND 0.006467f
C3755 VDD.n2828 GND 0.006467f
C3756 VDD.n2829 GND 0.006467f
C3757 VDD.n2830 GND 0.006467f
C3758 VDD.n2831 GND 0.006467f
C3759 VDD.n2832 GND 0.006467f
C3760 VDD.n2833 GND 0.006467f
C3761 VDD.n2834 GND 0.006467f
C3762 VDD.n2835 GND 0.006467f
C3763 VDD.n2836 GND 0.006467f
C3764 VDD.n2837 GND 0.005205f
C3765 VDD.n2838 GND 0.006467f
C3766 VDD.n2839 GND 0.005205f
C3767 VDD.n2840 GND 0.006467f
C3768 VDD.n2841 GND 0.006467f
C3769 VDD.n2842 GND 0.005205f
C3770 VDD.n2843 GND 0.005205f
C3771 VDD.n2844 GND 0.006467f
C3772 VDD.n2845 GND 0.006467f
C3773 VDD.n2846 GND 0.006467f
C3774 VDD.n2847 GND 0.006467f
C3775 VDD.n2848 GND 0.005205f
C3776 VDD.n2849 GND 0.005205f
C3777 VDD.n2850 GND 0.005205f
C3778 VDD.n2851 GND 0.006467f
C3779 VDD.n2852 GND 0.006467f
C3780 VDD.n2853 GND 0.006467f
C3781 VDD.n2854 GND 0.006467f
C3782 VDD.n2855 GND 0.005205f
C3783 VDD.n2856 GND 0.005205f
C3784 VDD.n2857 GND 0.00432f
C3785 VDD.n2858 GND 0.014445f
C3786 VDD.n2859 GND 0.014463f
C3787 VDD.n2860 GND 0.014463f
C3788 VDD.n2861 GND 0.002472f
C3789 VDD.t31 GND 0.089332f
C3790 VDD.t30 GND 0.10348f
C3791 VDD.t29 GND 0.482813f
C3792 VDD.n2862 GND 0.068834f
C3793 VDD.n2863 GND 0.04271f
C3794 VDD.n2864 GND 0.008016f
C3795 VDD.n2865 GND 0.002733f
C3796 VDD.n2866 GND 0.006467f
C3797 VDD.n2867 GND 0.006467f
C3798 VDD.n2868 GND 0.005205f
C3799 VDD.n2869 GND 0.005205f
C3800 VDD.n2870 GND 0.006467f
C3801 VDD.n2871 GND 0.006467f
C3802 VDD.n2872 GND 0.005205f
C3803 VDD.n2873 GND 0.005205f
C3804 VDD.n2874 GND 0.006467f
C3805 VDD.n2875 GND 0.006467f
C3806 VDD.n2876 GND 0.005205f
C3807 VDD.n2877 GND 0.005205f
C3808 VDD.n2878 GND 0.006467f
C3809 VDD.n2879 GND 0.006467f
C3810 VDD.n2880 GND 0.005205f
C3811 VDD.n2881 GND 0.005205f
C3812 VDD.n2882 GND 0.006467f
C3813 VDD.n2883 GND 0.006467f
C3814 VDD.n2884 GND 0.005205f
C3815 VDD.n2885 GND 0.005205f
C3816 VDD.n2886 GND 0.006467f
C3817 VDD.n2887 GND 0.006467f
C3818 VDD.n2888 GND 0.005205f
C3819 VDD.n2889 GND 0.006467f
C3820 VDD.n2890 GND 0.006467f
C3821 VDD.n2891 GND 0.005205f
C3822 VDD.n2892 GND 0.006467f
C3823 VDD.n2893 GND 0.006467f
C3824 VDD.n2894 GND 0.006467f
C3825 VDD.n2895 GND 0.010619f
C3826 VDD.n2896 GND 0.006467f
C3827 VDD.n2897 GND 0.006467f
C3828 VDD.n2898 GND 0.00354f
C3829 VDD.n2899 GND 0.005205f
C3830 VDD.n2900 GND 0.006467f
C3831 VDD.n2901 GND 0.006467f
C3832 VDD.n2902 GND 0.005205f
C3833 VDD.n2903 GND 0.005205f
C3834 VDD.n2904 GND 0.006467f
C3835 VDD.n2905 GND 0.006467f
C3836 VDD.n2906 GND 0.005205f
C3837 VDD.n2907 GND 0.005205f
C3838 VDD.n2908 GND 0.006467f
C3839 VDD.n2909 GND 0.006467f
C3840 VDD.n2910 GND 0.005205f
C3841 VDD.n2911 GND 0.005205f
C3842 VDD.n2912 GND 0.006467f
C3843 VDD.n2913 GND 0.006467f
C3844 VDD.n2914 GND 0.005205f
C3845 VDD.n2915 GND 0.005205f
C3846 VDD.n2916 GND 0.006467f
C3847 VDD.n2917 GND 0.006467f
C3848 VDD.n2918 GND 0.005205f
C3849 VDD.n2919 GND 0.005205f
C3850 VDD.n2920 GND 0.006467f
C3851 VDD.n2921 GND 0.006467f
C3852 VDD.n2922 GND 0.005205f
C3853 VDD.n2923 GND 0.006467f
C3854 VDD.n2924 GND 0.006467f
C3855 VDD.n2925 GND 0.006467f
C3856 VDD.n2926 GND 0.010619f
C3857 VDD.n2927 GND 0.004346f
C3858 VDD.n2928 GND 0.006467f
C3859 VDD.n2929 GND 0.006467f
C3860 VDD.n2930 GND 0.005205f
C3861 VDD.n2931 GND 0.005205f
C3862 VDD.n2932 GND 0.006467f
C3863 VDD.n2933 GND 0.006467f
C3864 VDD.n2934 GND 0.005205f
C3865 VDD.n2935 GND 0.005205f
C3866 VDD.n2936 GND 0.006467f
C3867 VDD.n2937 GND 0.006467f
C3868 VDD.n2938 GND 0.005205f
C3869 VDD.n2939 GND 0.005205f
C3870 VDD.n2940 GND 0.006467f
C3871 VDD.n2941 GND 0.006467f
C3872 VDD.n2942 GND 0.005205f
C3873 VDD.n2943 GND 0.006467f
C3874 VDD.n2944 GND 0.006467f
C3875 VDD.n2945 GND 0.005205f
C3876 VDD.n2946 GND 0.006467f
C3877 VDD.n2947 GND 0.006467f
C3878 VDD.n2948 GND 0.006467f
C3879 VDD.n2949 GND 0.005205f
C3880 VDD.n2950 GND 0.00432f
C3881 VDD.n2951 GND 0.014463f
C3882 VDD.n2952 GND 0.836271f
C3883 VDD.n2953 GND 0.487185f
C3884 VDD.n2954 GND 0.38361f
C3885 VDD.n2955 GND 0.006467f
C3886 VDD.n2956 GND 0.005205f
C3887 VDD.n2957 GND 0.005205f
C3888 VDD.n2958 GND 0.005205f
C3889 VDD.n2959 GND 0.006467f
C3890 VDD.n2960 GND 0.356758f
C3891 VDD.t12 GND 0.191805f
C3892 VDD.n2961 GND 0.218658f
C3893 VDD.n2962 GND 0.38361f
C3894 VDD.n2963 GND 0.006467f
C3895 VDD.n2964 GND 0.005205f
C3896 VDD.n2965 GND 0.005205f
C3897 VDD.n2966 GND 0.005205f
C3898 VDD.n2967 GND 0.006467f
C3899 VDD.n2968 GND 0.38361f
C3900 VDD.n2969 GND 0.38361f
C3901 VDD.n2970 GND 0.38361f
C3902 VDD.n2971 GND 0.006467f
C3903 VDD.n2972 GND 0.005205f
C3904 VDD.n2973 GND 0.005205f
C3905 VDD.n2974 GND 0.005205f
C3906 VDD.n2975 GND 0.006467f
C3907 VDD.n2976 GND 0.38361f
C3908 VDD.n2977 GND 0.006467f
C3909 VDD.n2978 GND 0.005205f
C3910 VDD.n2979 GND 0.005205f
C3911 VDD.n2980 GND 0.005205f
C3912 VDD.n2981 GND 0.006467f
C3913 VDD.t0 GND 0.38361f
C3914 VDD.n2982 GND 0.006467f
C3915 VDD.n2983 GND 0.005205f
C3916 VDD.n2984 GND 0.011738f
C3917 VDD.t2 GND 0.113194f
C3918 VDD.t74 GND 0.108896f
C3919 VDD.n2985 GND 0.307624f
C3920 VDD.t1 GND 0.108896f
C3921 VDD.n2986 GND 0.162532f
C3922 VDD.n2987 GND 1.15675f
C3923 a_n8413_8735.n0 GND 2.49088f
C3924 a_n8413_8735.t9 GND 0.092258f
C3925 a_n8413_8735.t10 GND 0.092258f
C3926 a_n8413_8735.t13 GND 0.092258f
C3927 a_n8413_8735.n1 GND 0.508889f
C3928 a_n8413_8735.t15 GND 0.092258f
C3929 a_n8413_8735.t8 GND 0.092258f
C3930 a_n8413_8735.n2 GND 0.472984f
C3931 a_n8413_8735.n3 GND 11.2455f
C3932 a_n8413_8735.t7 GND 0.639129f
C3933 a_n8413_8735.t5 GND 0.092258f
C3934 a_n8413_8735.t3 GND 0.092258f
C3935 a_n8413_8735.n4 GND 0.404151f
C3936 a_n8413_8735.n5 GND 2.68764f
C3937 a_n8413_8735.t2 GND 0.606632f
C3938 a_n8413_8735.t1 GND 0.606632f
C3939 a_n8413_8735.t0 GND 0.092258f
C3940 a_n8413_8735.t6 GND 0.092258f
C3941 a_n8413_8735.n6 GND 0.404151f
C3942 a_n8413_8735.n7 GND 1.595f
C3943 a_n8413_8735.t4 GND 0.606632f
C3944 a_n8413_8735.n8 GND 1.78414f
C3945 a_n8413_8735.n9 GND 5.540009f
C3946 a_n8413_8735.t11 GND 0.092258f
C3947 a_n8413_8735.t12 GND 0.092258f
C3948 a_n8413_8735.n10 GND 0.472982f
C3949 a_n8413_8735.n11 GND 4.81f
C3950 a_n8413_8735.n12 GND 0.517564f
C3951 a_n8413_8735.t14 GND 0.092258f
C3952 a_n8335_8538.n0 GND 12.5469f
C3953 a_n8335_8538.n1 GND 1.99566f
C3954 a_n8335_8538.n2 GND 16.563599f
C3955 a_n8335_8538.n3 GND 4.26795f
C3956 a_n8335_8538.n4 GND 0.853782f
C3957 a_n8335_8538.n5 GND 4.17681f
C3958 a_n8335_8538.n6 GND 0.853782f
C3959 a_n8335_8538.n7 GND 2.14042f
C3960 a_n8335_8538.n8 GND 2.18319f
C3961 a_n8335_8538.n9 GND 1.77969f
C3962 a_n8335_8538.t4 GND 0.195405f
C3963 a_n8335_8538.t16 GND 0.251585f
C3964 a_n8335_8538.t11 GND 1.82145f
C3965 a_n8335_8538.t3 GND 1.83952f
C3966 a_n8335_8538.t1 GND 1.78358f
C3967 a_n8335_8538.t29 GND 1.82145f
C3968 a_n8335_8538.t27 GND 1.83952f
C3969 a_n8335_8538.t26 GND 1.78358f
C3970 a_n8335_8538.t7 GND 1.81275f
C3971 a_n8335_8538.t13 GND 1.7913f
C3972 a_n8335_8538.t5 GND 1.83627f
C3973 a_n8335_8538.t31 GND 1.81275f
C3974 a_n8335_8538.t33 GND 1.78526f
C3975 a_n8335_8538.t35 GND 1.83329f
C3976 a_n8335_8538.t37 GND 1.82145f
C3977 a_n8335_8538.t17 GND 0.532239f
C3978 a_n8335_8538.t0 GND 0.260801f
C3979 a_n8335_8538.n10 GND 4.69113f
C3980 a_n8335_8538.t9 GND 1.82145f
C3981 a_n8335_8538.t10 GND 0.251585f
C3982 a_n8335_8538.t14 GND 0.195405f
C3983 a_n8335_8538.t6 GND 0.036316f
C3984 a_n8335_8538.t8 GND 0.238793f
C3985 a_n8335_8538.t28 GND 1.81275f
C3986 a_n8335_8538.t25 GND 1.79241f
C3987 a_n8335_8538.t24 GND 1.82358f
C3988 a_n8335_8538.t38 GND 1.81275f
C3989 a_n8335_8538.t18 GND 1.78445f
C3990 a_n8335_8538.t40 GND 1.78702f
C3991 a_n8335_8538.t22 GND 1.81275f
C3992 a_n8335_8538.t32 GND 1.78116f
C3993 a_n8335_8538.t34 GND 1.79221f
C3994 a_n8335_8538.t39 GND 1.81275f
C3995 a_n8335_8538.t20 GND 1.83276f
C3996 a_n8335_8538.t41 GND 1.78462f
C3997 a_n8335_8538.t19 GND 1.82145f
C3998 a_n8335_8538.t36 GND 1.85459f
C3999 a_n8335_8538.t23 GND 1.85485f
C4000 a_n8335_8538.t21 GND 1.82076f
C4001 a_n8335_8538.t30 GND 1.81275f
C4002 a_n8335_8538.t15 GND 1.81275f
C4003 a_n8335_8538.t12 GND 0.238792f
C4004 a_n8335_8538.t2 GND 0.036316f
.ends

