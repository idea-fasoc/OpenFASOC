* NGSPICE file created from diff_pair_sample_1649.ext - technology: sky130A

.subckt diff_pair_sample_1649 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VP.t0 VDD1.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=2.1294 pd=11.7 as=0.9009 ps=5.79 w=5.46 l=2.92
X1 VDD2.t3 VN.t0 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.9009 pd=5.79 as=2.1294 ps=11.7 w=5.46 l=2.92
X2 B.t17 B.t15 B.t16 B.t5 sky130_fd_pr__nfet_01v8 ad=2.1294 pd=11.7 as=0 ps=0 w=5.46 l=2.92
X3 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=2.1294 pd=11.7 as=0 ps=0 w=5.46 l=2.92
X4 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=2.1294 pd=11.7 as=0 ps=0 w=5.46 l=2.92
X5 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=2.1294 pd=11.7 as=0 ps=0 w=5.46 l=2.92
X6 VTAIL.t1 VN.t1 VDD2.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=2.1294 pd=11.7 as=0.9009 ps=5.79 w=5.46 l=2.92
X7 VDD2.t1 VN.t2 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.9009 pd=5.79 as=2.1294 ps=11.7 w=5.46 l=2.92
X8 VDD1.t0 VP.t1 VTAIL.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=0.9009 pd=5.79 as=2.1294 ps=11.7 w=5.46 l=2.92
X9 VDD1.t1 VP.t2 VTAIL.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=0.9009 pd=5.79 as=2.1294 ps=11.7 w=5.46 l=2.92
X10 VTAIL.t0 VN.t3 VDD2.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.1294 pd=11.7 as=0.9009 ps=5.79 w=5.46 l=2.92
X11 VTAIL.t4 VP.t3 VDD1.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=2.1294 pd=11.7 as=0.9009 ps=5.79 w=5.46 l=2.92
R0 VP.n15 VP.n14 161.3
R1 VP.n13 VP.n1 161.3
R2 VP.n12 VP.n11 161.3
R3 VP.n10 VP.n2 161.3
R4 VP.n9 VP.n8 161.3
R5 VP.n7 VP.n3 161.3
R6 VP.n4 VP.t3 79.4663
R7 VP.n4 VP.t1 78.4926
R8 VP.n6 VP.n5 71.8017
R9 VP.n16 VP.n0 71.8017
R10 VP.n12 VP.n2 56.5617
R11 VP.n5 VP.n4 45.4679
R12 VP.n6 VP.t0 45.0642
R13 VP.n0 VP.t2 45.0642
R14 VP.n8 VP.n7 24.5923
R15 VP.n8 VP.n2 24.5923
R16 VP.n13 VP.n12 24.5923
R17 VP.n14 VP.n13 24.5923
R18 VP.n7 VP.n6 18.4444
R19 VP.n14 VP.n0 18.4444
R20 VP.n5 VP.n3 0.354861
R21 VP.n16 VP.n15 0.354861
R22 VP VP.n16 0.267071
R23 VP.n9 VP.n3 0.189894
R24 VP.n10 VP.n9 0.189894
R25 VP.n11 VP.n10 0.189894
R26 VP.n11 VP.n1 0.189894
R27 VP.n15 VP.n1 0.189894
R28 VDD1 VDD1.n1 107.809
R29 VDD1 VDD1.n0 70.5149
R30 VDD1.n0 VDD1.t3 3.62687
R31 VDD1.n0 VDD1.t0 3.62687
R32 VDD1.n1 VDD1.t2 3.62687
R33 VDD1.n1 VDD1.t1 3.62687
R34 VTAIL.n5 VTAIL.t4 57.4053
R35 VTAIL.n4 VTAIL.t3 57.4053
R36 VTAIL.n3 VTAIL.t1 57.4053
R37 VTAIL.n6 VTAIL.t6 57.4043
R38 VTAIL.n7 VTAIL.t2 57.4043
R39 VTAIL.n0 VTAIL.t0 57.4043
R40 VTAIL.n1 VTAIL.t5 57.4043
R41 VTAIL.n2 VTAIL.t7 57.4043
R42 VTAIL.n7 VTAIL.n6 19.8755
R43 VTAIL.n3 VTAIL.n2 19.8755
R44 VTAIL.n4 VTAIL.n3 2.80222
R45 VTAIL.n6 VTAIL.n5 2.80222
R46 VTAIL.n2 VTAIL.n1 2.80222
R47 VTAIL VTAIL.n0 1.45955
R48 VTAIL VTAIL.n7 1.34317
R49 VTAIL.n5 VTAIL.n4 0.470328
R50 VTAIL.n1 VTAIL.n0 0.470328
R51 B.n579 B.n578 585
R52 B.n207 B.n96 585
R53 B.n206 B.n205 585
R54 B.n204 B.n203 585
R55 B.n202 B.n201 585
R56 B.n200 B.n199 585
R57 B.n198 B.n197 585
R58 B.n196 B.n195 585
R59 B.n194 B.n193 585
R60 B.n192 B.n191 585
R61 B.n190 B.n189 585
R62 B.n188 B.n187 585
R63 B.n186 B.n185 585
R64 B.n184 B.n183 585
R65 B.n182 B.n181 585
R66 B.n180 B.n179 585
R67 B.n178 B.n177 585
R68 B.n176 B.n175 585
R69 B.n174 B.n173 585
R70 B.n172 B.n171 585
R71 B.n170 B.n169 585
R72 B.n168 B.n167 585
R73 B.n166 B.n165 585
R74 B.n164 B.n163 585
R75 B.n162 B.n161 585
R76 B.n160 B.n159 585
R77 B.n158 B.n157 585
R78 B.n156 B.n155 585
R79 B.n154 B.n153 585
R80 B.n152 B.n151 585
R81 B.n150 B.n149 585
R82 B.n148 B.n147 585
R83 B.n146 B.n145 585
R84 B.n144 B.n143 585
R85 B.n142 B.n141 585
R86 B.n140 B.n139 585
R87 B.n138 B.n137 585
R88 B.n136 B.n135 585
R89 B.n134 B.n133 585
R90 B.n132 B.n131 585
R91 B.n130 B.n129 585
R92 B.n128 B.n127 585
R93 B.n126 B.n125 585
R94 B.n124 B.n123 585
R95 B.n122 B.n121 585
R96 B.n120 B.n119 585
R97 B.n118 B.n117 585
R98 B.n116 B.n115 585
R99 B.n114 B.n113 585
R100 B.n112 B.n111 585
R101 B.n110 B.n109 585
R102 B.n108 B.n107 585
R103 B.n106 B.n105 585
R104 B.n104 B.n103 585
R105 B.n577 B.n69 585
R106 B.n582 B.n69 585
R107 B.n576 B.n68 585
R108 B.n583 B.n68 585
R109 B.n575 B.n574 585
R110 B.n574 B.n64 585
R111 B.n573 B.n63 585
R112 B.n589 B.n63 585
R113 B.n572 B.n62 585
R114 B.n590 B.n62 585
R115 B.n571 B.n61 585
R116 B.n591 B.n61 585
R117 B.n570 B.n569 585
R118 B.n569 B.n57 585
R119 B.n568 B.n56 585
R120 B.n597 B.n56 585
R121 B.n567 B.n55 585
R122 B.n598 B.n55 585
R123 B.n566 B.n54 585
R124 B.n599 B.n54 585
R125 B.n565 B.n564 585
R126 B.n564 B.n50 585
R127 B.n563 B.n49 585
R128 B.n605 B.n49 585
R129 B.n562 B.n48 585
R130 B.n606 B.n48 585
R131 B.n561 B.n47 585
R132 B.n607 B.n47 585
R133 B.n560 B.n559 585
R134 B.n559 B.n43 585
R135 B.n558 B.n42 585
R136 B.n613 B.n42 585
R137 B.n557 B.n41 585
R138 B.n614 B.n41 585
R139 B.n556 B.n40 585
R140 B.n615 B.n40 585
R141 B.n555 B.n554 585
R142 B.n554 B.n36 585
R143 B.n553 B.n35 585
R144 B.n621 B.n35 585
R145 B.n552 B.n34 585
R146 B.n622 B.n34 585
R147 B.n551 B.n33 585
R148 B.n623 B.n33 585
R149 B.n550 B.n549 585
R150 B.n549 B.n29 585
R151 B.n548 B.n28 585
R152 B.n629 B.n28 585
R153 B.n547 B.n27 585
R154 B.n630 B.n27 585
R155 B.n546 B.n26 585
R156 B.n631 B.n26 585
R157 B.n545 B.n544 585
R158 B.n544 B.n22 585
R159 B.n543 B.n21 585
R160 B.n637 B.n21 585
R161 B.n542 B.n20 585
R162 B.n638 B.n20 585
R163 B.n541 B.n19 585
R164 B.n639 B.n19 585
R165 B.n540 B.n539 585
R166 B.n539 B.n18 585
R167 B.n538 B.n14 585
R168 B.n645 B.n14 585
R169 B.n537 B.n13 585
R170 B.n646 B.n13 585
R171 B.n536 B.n12 585
R172 B.n647 B.n12 585
R173 B.n535 B.n534 585
R174 B.n534 B.n8 585
R175 B.n533 B.n7 585
R176 B.n653 B.n7 585
R177 B.n532 B.n6 585
R178 B.n654 B.n6 585
R179 B.n531 B.n5 585
R180 B.n655 B.n5 585
R181 B.n530 B.n529 585
R182 B.n529 B.n4 585
R183 B.n528 B.n208 585
R184 B.n528 B.n527 585
R185 B.n518 B.n209 585
R186 B.n210 B.n209 585
R187 B.n520 B.n519 585
R188 B.n521 B.n520 585
R189 B.n517 B.n215 585
R190 B.n215 B.n214 585
R191 B.n516 B.n515 585
R192 B.n515 B.n514 585
R193 B.n217 B.n216 585
R194 B.n507 B.n217 585
R195 B.n506 B.n505 585
R196 B.n508 B.n506 585
R197 B.n504 B.n222 585
R198 B.n222 B.n221 585
R199 B.n503 B.n502 585
R200 B.n502 B.n501 585
R201 B.n224 B.n223 585
R202 B.n225 B.n224 585
R203 B.n494 B.n493 585
R204 B.n495 B.n494 585
R205 B.n492 B.n230 585
R206 B.n230 B.n229 585
R207 B.n491 B.n490 585
R208 B.n490 B.n489 585
R209 B.n232 B.n231 585
R210 B.n233 B.n232 585
R211 B.n482 B.n481 585
R212 B.n483 B.n482 585
R213 B.n480 B.n238 585
R214 B.n238 B.n237 585
R215 B.n479 B.n478 585
R216 B.n478 B.n477 585
R217 B.n240 B.n239 585
R218 B.n241 B.n240 585
R219 B.n470 B.n469 585
R220 B.n471 B.n470 585
R221 B.n468 B.n246 585
R222 B.n246 B.n245 585
R223 B.n467 B.n466 585
R224 B.n466 B.n465 585
R225 B.n248 B.n247 585
R226 B.n249 B.n248 585
R227 B.n458 B.n457 585
R228 B.n459 B.n458 585
R229 B.n456 B.n254 585
R230 B.n254 B.n253 585
R231 B.n455 B.n454 585
R232 B.n454 B.n453 585
R233 B.n256 B.n255 585
R234 B.n257 B.n256 585
R235 B.n446 B.n445 585
R236 B.n447 B.n446 585
R237 B.n444 B.n261 585
R238 B.n265 B.n261 585
R239 B.n443 B.n442 585
R240 B.n442 B.n441 585
R241 B.n263 B.n262 585
R242 B.n264 B.n263 585
R243 B.n434 B.n433 585
R244 B.n435 B.n434 585
R245 B.n432 B.n270 585
R246 B.n270 B.n269 585
R247 B.n431 B.n430 585
R248 B.n430 B.n429 585
R249 B.n272 B.n271 585
R250 B.n273 B.n272 585
R251 B.n422 B.n421 585
R252 B.n423 B.n422 585
R253 B.n420 B.n278 585
R254 B.n278 B.n277 585
R255 B.n415 B.n414 585
R256 B.n413 B.n307 585
R257 B.n412 B.n306 585
R258 B.n417 B.n306 585
R259 B.n411 B.n410 585
R260 B.n409 B.n408 585
R261 B.n407 B.n406 585
R262 B.n405 B.n404 585
R263 B.n403 B.n402 585
R264 B.n401 B.n400 585
R265 B.n399 B.n398 585
R266 B.n397 B.n396 585
R267 B.n395 B.n394 585
R268 B.n393 B.n392 585
R269 B.n391 B.n390 585
R270 B.n389 B.n388 585
R271 B.n387 B.n386 585
R272 B.n385 B.n384 585
R273 B.n383 B.n382 585
R274 B.n381 B.n380 585
R275 B.n379 B.n378 585
R276 B.n377 B.n376 585
R277 B.n375 B.n374 585
R278 B.n372 B.n371 585
R279 B.n370 B.n369 585
R280 B.n368 B.n367 585
R281 B.n366 B.n365 585
R282 B.n364 B.n363 585
R283 B.n362 B.n361 585
R284 B.n360 B.n359 585
R285 B.n358 B.n357 585
R286 B.n356 B.n355 585
R287 B.n354 B.n353 585
R288 B.n351 B.n350 585
R289 B.n349 B.n348 585
R290 B.n347 B.n346 585
R291 B.n345 B.n344 585
R292 B.n343 B.n342 585
R293 B.n341 B.n340 585
R294 B.n339 B.n338 585
R295 B.n337 B.n336 585
R296 B.n335 B.n334 585
R297 B.n333 B.n332 585
R298 B.n331 B.n330 585
R299 B.n329 B.n328 585
R300 B.n327 B.n326 585
R301 B.n325 B.n324 585
R302 B.n323 B.n322 585
R303 B.n321 B.n320 585
R304 B.n319 B.n318 585
R305 B.n317 B.n316 585
R306 B.n315 B.n314 585
R307 B.n313 B.n312 585
R308 B.n280 B.n279 585
R309 B.n419 B.n418 585
R310 B.n418 B.n417 585
R311 B.n276 B.n275 585
R312 B.n277 B.n276 585
R313 B.n425 B.n424 585
R314 B.n424 B.n423 585
R315 B.n426 B.n274 585
R316 B.n274 B.n273 585
R317 B.n428 B.n427 585
R318 B.n429 B.n428 585
R319 B.n268 B.n267 585
R320 B.n269 B.n268 585
R321 B.n437 B.n436 585
R322 B.n436 B.n435 585
R323 B.n438 B.n266 585
R324 B.n266 B.n264 585
R325 B.n440 B.n439 585
R326 B.n441 B.n440 585
R327 B.n260 B.n259 585
R328 B.n265 B.n260 585
R329 B.n449 B.n448 585
R330 B.n448 B.n447 585
R331 B.n450 B.n258 585
R332 B.n258 B.n257 585
R333 B.n452 B.n451 585
R334 B.n453 B.n452 585
R335 B.n252 B.n251 585
R336 B.n253 B.n252 585
R337 B.n461 B.n460 585
R338 B.n460 B.n459 585
R339 B.n462 B.n250 585
R340 B.n250 B.n249 585
R341 B.n464 B.n463 585
R342 B.n465 B.n464 585
R343 B.n244 B.n243 585
R344 B.n245 B.n244 585
R345 B.n473 B.n472 585
R346 B.n472 B.n471 585
R347 B.n474 B.n242 585
R348 B.n242 B.n241 585
R349 B.n476 B.n475 585
R350 B.n477 B.n476 585
R351 B.n236 B.n235 585
R352 B.n237 B.n236 585
R353 B.n485 B.n484 585
R354 B.n484 B.n483 585
R355 B.n486 B.n234 585
R356 B.n234 B.n233 585
R357 B.n488 B.n487 585
R358 B.n489 B.n488 585
R359 B.n228 B.n227 585
R360 B.n229 B.n228 585
R361 B.n497 B.n496 585
R362 B.n496 B.n495 585
R363 B.n498 B.n226 585
R364 B.n226 B.n225 585
R365 B.n500 B.n499 585
R366 B.n501 B.n500 585
R367 B.n220 B.n219 585
R368 B.n221 B.n220 585
R369 B.n510 B.n509 585
R370 B.n509 B.n508 585
R371 B.n511 B.n218 585
R372 B.n507 B.n218 585
R373 B.n513 B.n512 585
R374 B.n514 B.n513 585
R375 B.n213 B.n212 585
R376 B.n214 B.n213 585
R377 B.n523 B.n522 585
R378 B.n522 B.n521 585
R379 B.n524 B.n211 585
R380 B.n211 B.n210 585
R381 B.n526 B.n525 585
R382 B.n527 B.n526 585
R383 B.n2 B.n0 585
R384 B.n4 B.n2 585
R385 B.n3 B.n1 585
R386 B.n654 B.n3 585
R387 B.n652 B.n651 585
R388 B.n653 B.n652 585
R389 B.n650 B.n9 585
R390 B.n9 B.n8 585
R391 B.n649 B.n648 585
R392 B.n648 B.n647 585
R393 B.n11 B.n10 585
R394 B.n646 B.n11 585
R395 B.n644 B.n643 585
R396 B.n645 B.n644 585
R397 B.n642 B.n15 585
R398 B.n18 B.n15 585
R399 B.n641 B.n640 585
R400 B.n640 B.n639 585
R401 B.n17 B.n16 585
R402 B.n638 B.n17 585
R403 B.n636 B.n635 585
R404 B.n637 B.n636 585
R405 B.n634 B.n23 585
R406 B.n23 B.n22 585
R407 B.n633 B.n632 585
R408 B.n632 B.n631 585
R409 B.n25 B.n24 585
R410 B.n630 B.n25 585
R411 B.n628 B.n627 585
R412 B.n629 B.n628 585
R413 B.n626 B.n30 585
R414 B.n30 B.n29 585
R415 B.n625 B.n624 585
R416 B.n624 B.n623 585
R417 B.n32 B.n31 585
R418 B.n622 B.n32 585
R419 B.n620 B.n619 585
R420 B.n621 B.n620 585
R421 B.n618 B.n37 585
R422 B.n37 B.n36 585
R423 B.n617 B.n616 585
R424 B.n616 B.n615 585
R425 B.n39 B.n38 585
R426 B.n614 B.n39 585
R427 B.n612 B.n611 585
R428 B.n613 B.n612 585
R429 B.n610 B.n44 585
R430 B.n44 B.n43 585
R431 B.n609 B.n608 585
R432 B.n608 B.n607 585
R433 B.n46 B.n45 585
R434 B.n606 B.n46 585
R435 B.n604 B.n603 585
R436 B.n605 B.n604 585
R437 B.n602 B.n51 585
R438 B.n51 B.n50 585
R439 B.n601 B.n600 585
R440 B.n600 B.n599 585
R441 B.n53 B.n52 585
R442 B.n598 B.n53 585
R443 B.n596 B.n595 585
R444 B.n597 B.n596 585
R445 B.n594 B.n58 585
R446 B.n58 B.n57 585
R447 B.n593 B.n592 585
R448 B.n592 B.n591 585
R449 B.n60 B.n59 585
R450 B.n590 B.n60 585
R451 B.n588 B.n587 585
R452 B.n589 B.n588 585
R453 B.n586 B.n65 585
R454 B.n65 B.n64 585
R455 B.n585 B.n584 585
R456 B.n584 B.n583 585
R457 B.n67 B.n66 585
R458 B.n582 B.n67 585
R459 B.n657 B.n656 585
R460 B.n656 B.n655 585
R461 B.n415 B.n276 492.5
R462 B.n103 B.n67 492.5
R463 B.n418 B.n278 492.5
R464 B.n579 B.n69 492.5
R465 B.n581 B.n580 256.663
R466 B.n581 B.n95 256.663
R467 B.n581 B.n94 256.663
R468 B.n581 B.n93 256.663
R469 B.n581 B.n92 256.663
R470 B.n581 B.n91 256.663
R471 B.n581 B.n90 256.663
R472 B.n581 B.n89 256.663
R473 B.n581 B.n88 256.663
R474 B.n581 B.n87 256.663
R475 B.n581 B.n86 256.663
R476 B.n581 B.n85 256.663
R477 B.n581 B.n84 256.663
R478 B.n581 B.n83 256.663
R479 B.n581 B.n82 256.663
R480 B.n581 B.n81 256.663
R481 B.n581 B.n80 256.663
R482 B.n581 B.n79 256.663
R483 B.n581 B.n78 256.663
R484 B.n581 B.n77 256.663
R485 B.n581 B.n76 256.663
R486 B.n581 B.n75 256.663
R487 B.n581 B.n74 256.663
R488 B.n581 B.n73 256.663
R489 B.n581 B.n72 256.663
R490 B.n581 B.n71 256.663
R491 B.n581 B.n70 256.663
R492 B.n417 B.n416 256.663
R493 B.n417 B.n281 256.663
R494 B.n417 B.n282 256.663
R495 B.n417 B.n283 256.663
R496 B.n417 B.n284 256.663
R497 B.n417 B.n285 256.663
R498 B.n417 B.n286 256.663
R499 B.n417 B.n287 256.663
R500 B.n417 B.n288 256.663
R501 B.n417 B.n289 256.663
R502 B.n417 B.n290 256.663
R503 B.n417 B.n291 256.663
R504 B.n417 B.n292 256.663
R505 B.n417 B.n293 256.663
R506 B.n417 B.n294 256.663
R507 B.n417 B.n295 256.663
R508 B.n417 B.n296 256.663
R509 B.n417 B.n297 256.663
R510 B.n417 B.n298 256.663
R511 B.n417 B.n299 256.663
R512 B.n417 B.n300 256.663
R513 B.n417 B.n301 256.663
R514 B.n417 B.n302 256.663
R515 B.n417 B.n303 256.663
R516 B.n417 B.n304 256.663
R517 B.n417 B.n305 256.663
R518 B.n310 B.t8 253.548
R519 B.n308 B.t12 253.548
R520 B.n100 B.t15 253.548
R521 B.n97 B.t4 253.548
R522 B.n424 B.n276 163.367
R523 B.n424 B.n274 163.367
R524 B.n428 B.n274 163.367
R525 B.n428 B.n268 163.367
R526 B.n436 B.n268 163.367
R527 B.n436 B.n266 163.367
R528 B.n440 B.n266 163.367
R529 B.n440 B.n260 163.367
R530 B.n448 B.n260 163.367
R531 B.n448 B.n258 163.367
R532 B.n452 B.n258 163.367
R533 B.n452 B.n252 163.367
R534 B.n460 B.n252 163.367
R535 B.n460 B.n250 163.367
R536 B.n464 B.n250 163.367
R537 B.n464 B.n244 163.367
R538 B.n472 B.n244 163.367
R539 B.n472 B.n242 163.367
R540 B.n476 B.n242 163.367
R541 B.n476 B.n236 163.367
R542 B.n484 B.n236 163.367
R543 B.n484 B.n234 163.367
R544 B.n488 B.n234 163.367
R545 B.n488 B.n228 163.367
R546 B.n496 B.n228 163.367
R547 B.n496 B.n226 163.367
R548 B.n500 B.n226 163.367
R549 B.n500 B.n220 163.367
R550 B.n509 B.n220 163.367
R551 B.n509 B.n218 163.367
R552 B.n513 B.n218 163.367
R553 B.n513 B.n213 163.367
R554 B.n522 B.n213 163.367
R555 B.n522 B.n211 163.367
R556 B.n526 B.n211 163.367
R557 B.n526 B.n2 163.367
R558 B.n656 B.n2 163.367
R559 B.n656 B.n3 163.367
R560 B.n652 B.n3 163.367
R561 B.n652 B.n9 163.367
R562 B.n648 B.n9 163.367
R563 B.n648 B.n11 163.367
R564 B.n644 B.n11 163.367
R565 B.n644 B.n15 163.367
R566 B.n640 B.n15 163.367
R567 B.n640 B.n17 163.367
R568 B.n636 B.n17 163.367
R569 B.n636 B.n23 163.367
R570 B.n632 B.n23 163.367
R571 B.n632 B.n25 163.367
R572 B.n628 B.n25 163.367
R573 B.n628 B.n30 163.367
R574 B.n624 B.n30 163.367
R575 B.n624 B.n32 163.367
R576 B.n620 B.n32 163.367
R577 B.n620 B.n37 163.367
R578 B.n616 B.n37 163.367
R579 B.n616 B.n39 163.367
R580 B.n612 B.n39 163.367
R581 B.n612 B.n44 163.367
R582 B.n608 B.n44 163.367
R583 B.n608 B.n46 163.367
R584 B.n604 B.n46 163.367
R585 B.n604 B.n51 163.367
R586 B.n600 B.n51 163.367
R587 B.n600 B.n53 163.367
R588 B.n596 B.n53 163.367
R589 B.n596 B.n58 163.367
R590 B.n592 B.n58 163.367
R591 B.n592 B.n60 163.367
R592 B.n588 B.n60 163.367
R593 B.n588 B.n65 163.367
R594 B.n584 B.n65 163.367
R595 B.n584 B.n67 163.367
R596 B.n307 B.n306 163.367
R597 B.n410 B.n306 163.367
R598 B.n408 B.n407 163.367
R599 B.n404 B.n403 163.367
R600 B.n400 B.n399 163.367
R601 B.n396 B.n395 163.367
R602 B.n392 B.n391 163.367
R603 B.n388 B.n387 163.367
R604 B.n384 B.n383 163.367
R605 B.n380 B.n379 163.367
R606 B.n376 B.n375 163.367
R607 B.n371 B.n370 163.367
R608 B.n367 B.n366 163.367
R609 B.n363 B.n362 163.367
R610 B.n359 B.n358 163.367
R611 B.n355 B.n354 163.367
R612 B.n350 B.n349 163.367
R613 B.n346 B.n345 163.367
R614 B.n342 B.n341 163.367
R615 B.n338 B.n337 163.367
R616 B.n334 B.n333 163.367
R617 B.n330 B.n329 163.367
R618 B.n326 B.n325 163.367
R619 B.n322 B.n321 163.367
R620 B.n318 B.n317 163.367
R621 B.n314 B.n313 163.367
R622 B.n418 B.n280 163.367
R623 B.n422 B.n278 163.367
R624 B.n422 B.n272 163.367
R625 B.n430 B.n272 163.367
R626 B.n430 B.n270 163.367
R627 B.n434 B.n270 163.367
R628 B.n434 B.n263 163.367
R629 B.n442 B.n263 163.367
R630 B.n442 B.n261 163.367
R631 B.n446 B.n261 163.367
R632 B.n446 B.n256 163.367
R633 B.n454 B.n256 163.367
R634 B.n454 B.n254 163.367
R635 B.n458 B.n254 163.367
R636 B.n458 B.n248 163.367
R637 B.n466 B.n248 163.367
R638 B.n466 B.n246 163.367
R639 B.n470 B.n246 163.367
R640 B.n470 B.n240 163.367
R641 B.n478 B.n240 163.367
R642 B.n478 B.n238 163.367
R643 B.n482 B.n238 163.367
R644 B.n482 B.n232 163.367
R645 B.n490 B.n232 163.367
R646 B.n490 B.n230 163.367
R647 B.n494 B.n230 163.367
R648 B.n494 B.n224 163.367
R649 B.n502 B.n224 163.367
R650 B.n502 B.n222 163.367
R651 B.n506 B.n222 163.367
R652 B.n506 B.n217 163.367
R653 B.n515 B.n217 163.367
R654 B.n515 B.n215 163.367
R655 B.n520 B.n215 163.367
R656 B.n520 B.n209 163.367
R657 B.n528 B.n209 163.367
R658 B.n529 B.n528 163.367
R659 B.n529 B.n5 163.367
R660 B.n6 B.n5 163.367
R661 B.n7 B.n6 163.367
R662 B.n534 B.n7 163.367
R663 B.n534 B.n12 163.367
R664 B.n13 B.n12 163.367
R665 B.n14 B.n13 163.367
R666 B.n539 B.n14 163.367
R667 B.n539 B.n19 163.367
R668 B.n20 B.n19 163.367
R669 B.n21 B.n20 163.367
R670 B.n544 B.n21 163.367
R671 B.n544 B.n26 163.367
R672 B.n27 B.n26 163.367
R673 B.n28 B.n27 163.367
R674 B.n549 B.n28 163.367
R675 B.n549 B.n33 163.367
R676 B.n34 B.n33 163.367
R677 B.n35 B.n34 163.367
R678 B.n554 B.n35 163.367
R679 B.n554 B.n40 163.367
R680 B.n41 B.n40 163.367
R681 B.n42 B.n41 163.367
R682 B.n559 B.n42 163.367
R683 B.n559 B.n47 163.367
R684 B.n48 B.n47 163.367
R685 B.n49 B.n48 163.367
R686 B.n564 B.n49 163.367
R687 B.n564 B.n54 163.367
R688 B.n55 B.n54 163.367
R689 B.n56 B.n55 163.367
R690 B.n569 B.n56 163.367
R691 B.n569 B.n61 163.367
R692 B.n62 B.n61 163.367
R693 B.n63 B.n62 163.367
R694 B.n574 B.n63 163.367
R695 B.n574 B.n68 163.367
R696 B.n69 B.n68 163.367
R697 B.n107 B.n106 163.367
R698 B.n111 B.n110 163.367
R699 B.n115 B.n114 163.367
R700 B.n119 B.n118 163.367
R701 B.n123 B.n122 163.367
R702 B.n127 B.n126 163.367
R703 B.n131 B.n130 163.367
R704 B.n135 B.n134 163.367
R705 B.n139 B.n138 163.367
R706 B.n143 B.n142 163.367
R707 B.n147 B.n146 163.367
R708 B.n151 B.n150 163.367
R709 B.n155 B.n154 163.367
R710 B.n159 B.n158 163.367
R711 B.n163 B.n162 163.367
R712 B.n167 B.n166 163.367
R713 B.n171 B.n170 163.367
R714 B.n175 B.n174 163.367
R715 B.n179 B.n178 163.367
R716 B.n183 B.n182 163.367
R717 B.n187 B.n186 163.367
R718 B.n191 B.n190 163.367
R719 B.n195 B.n194 163.367
R720 B.n199 B.n198 163.367
R721 B.n203 B.n202 163.367
R722 B.n205 B.n96 163.367
R723 B.n310 B.t11 133.208
R724 B.n97 B.t6 133.208
R725 B.n308 B.t14 133.203
R726 B.n100 B.t16 133.203
R727 B.n417 B.n277 111.692
R728 B.n582 B.n581 111.692
R729 B.n416 B.n415 71.676
R730 B.n410 B.n281 71.676
R731 B.n407 B.n282 71.676
R732 B.n403 B.n283 71.676
R733 B.n399 B.n284 71.676
R734 B.n395 B.n285 71.676
R735 B.n391 B.n286 71.676
R736 B.n387 B.n287 71.676
R737 B.n383 B.n288 71.676
R738 B.n379 B.n289 71.676
R739 B.n375 B.n290 71.676
R740 B.n370 B.n291 71.676
R741 B.n366 B.n292 71.676
R742 B.n362 B.n293 71.676
R743 B.n358 B.n294 71.676
R744 B.n354 B.n295 71.676
R745 B.n349 B.n296 71.676
R746 B.n345 B.n297 71.676
R747 B.n341 B.n298 71.676
R748 B.n337 B.n299 71.676
R749 B.n333 B.n300 71.676
R750 B.n329 B.n301 71.676
R751 B.n325 B.n302 71.676
R752 B.n321 B.n303 71.676
R753 B.n317 B.n304 71.676
R754 B.n313 B.n305 71.676
R755 B.n103 B.n70 71.676
R756 B.n107 B.n71 71.676
R757 B.n111 B.n72 71.676
R758 B.n115 B.n73 71.676
R759 B.n119 B.n74 71.676
R760 B.n123 B.n75 71.676
R761 B.n127 B.n76 71.676
R762 B.n131 B.n77 71.676
R763 B.n135 B.n78 71.676
R764 B.n139 B.n79 71.676
R765 B.n143 B.n80 71.676
R766 B.n147 B.n81 71.676
R767 B.n151 B.n82 71.676
R768 B.n155 B.n83 71.676
R769 B.n159 B.n84 71.676
R770 B.n163 B.n85 71.676
R771 B.n167 B.n86 71.676
R772 B.n171 B.n87 71.676
R773 B.n175 B.n88 71.676
R774 B.n179 B.n89 71.676
R775 B.n183 B.n90 71.676
R776 B.n187 B.n91 71.676
R777 B.n191 B.n92 71.676
R778 B.n195 B.n93 71.676
R779 B.n199 B.n94 71.676
R780 B.n203 B.n95 71.676
R781 B.n580 B.n96 71.676
R782 B.n580 B.n579 71.676
R783 B.n205 B.n95 71.676
R784 B.n202 B.n94 71.676
R785 B.n198 B.n93 71.676
R786 B.n194 B.n92 71.676
R787 B.n190 B.n91 71.676
R788 B.n186 B.n90 71.676
R789 B.n182 B.n89 71.676
R790 B.n178 B.n88 71.676
R791 B.n174 B.n87 71.676
R792 B.n170 B.n86 71.676
R793 B.n166 B.n85 71.676
R794 B.n162 B.n84 71.676
R795 B.n158 B.n83 71.676
R796 B.n154 B.n82 71.676
R797 B.n150 B.n81 71.676
R798 B.n146 B.n80 71.676
R799 B.n142 B.n79 71.676
R800 B.n138 B.n78 71.676
R801 B.n134 B.n77 71.676
R802 B.n130 B.n76 71.676
R803 B.n126 B.n75 71.676
R804 B.n122 B.n74 71.676
R805 B.n118 B.n73 71.676
R806 B.n114 B.n72 71.676
R807 B.n110 B.n71 71.676
R808 B.n106 B.n70 71.676
R809 B.n416 B.n307 71.676
R810 B.n408 B.n281 71.676
R811 B.n404 B.n282 71.676
R812 B.n400 B.n283 71.676
R813 B.n396 B.n284 71.676
R814 B.n392 B.n285 71.676
R815 B.n388 B.n286 71.676
R816 B.n384 B.n287 71.676
R817 B.n380 B.n288 71.676
R818 B.n376 B.n289 71.676
R819 B.n371 B.n290 71.676
R820 B.n367 B.n291 71.676
R821 B.n363 B.n292 71.676
R822 B.n359 B.n293 71.676
R823 B.n355 B.n294 71.676
R824 B.n350 B.n295 71.676
R825 B.n346 B.n296 71.676
R826 B.n342 B.n297 71.676
R827 B.n338 B.n298 71.676
R828 B.n334 B.n299 71.676
R829 B.n330 B.n300 71.676
R830 B.n326 B.n301 71.676
R831 B.n322 B.n302 71.676
R832 B.n318 B.n303 71.676
R833 B.n314 B.n304 71.676
R834 B.n305 B.n280 71.676
R835 B.n311 B.t10 70.1786
R836 B.n98 B.t7 70.1786
R837 B.n309 B.t13 70.1728
R838 B.n101 B.t17 70.1728
R839 B.n423 B.n277 69.6791
R840 B.n423 B.n273 69.6791
R841 B.n429 B.n273 69.6791
R842 B.n429 B.n269 69.6791
R843 B.n435 B.n269 69.6791
R844 B.n435 B.n264 69.6791
R845 B.n441 B.n264 69.6791
R846 B.n441 B.n265 69.6791
R847 B.n447 B.n257 69.6791
R848 B.n453 B.n257 69.6791
R849 B.n453 B.n253 69.6791
R850 B.n459 B.n253 69.6791
R851 B.n459 B.n249 69.6791
R852 B.n465 B.n249 69.6791
R853 B.n465 B.n245 69.6791
R854 B.n471 B.n245 69.6791
R855 B.n471 B.n241 69.6791
R856 B.n477 B.n241 69.6791
R857 B.n477 B.n237 69.6791
R858 B.n483 B.n237 69.6791
R859 B.n489 B.n233 69.6791
R860 B.n489 B.n229 69.6791
R861 B.n495 B.n229 69.6791
R862 B.n495 B.n225 69.6791
R863 B.n501 B.n225 69.6791
R864 B.n501 B.n221 69.6791
R865 B.n508 B.n221 69.6791
R866 B.n508 B.n507 69.6791
R867 B.n514 B.n214 69.6791
R868 B.n521 B.n214 69.6791
R869 B.n521 B.n210 69.6791
R870 B.n527 B.n210 69.6791
R871 B.n527 B.n4 69.6791
R872 B.n655 B.n4 69.6791
R873 B.n655 B.n654 69.6791
R874 B.n654 B.n653 69.6791
R875 B.n653 B.n8 69.6791
R876 B.n647 B.n8 69.6791
R877 B.n647 B.n646 69.6791
R878 B.n646 B.n645 69.6791
R879 B.n639 B.n18 69.6791
R880 B.n639 B.n638 69.6791
R881 B.n638 B.n637 69.6791
R882 B.n637 B.n22 69.6791
R883 B.n631 B.n22 69.6791
R884 B.n631 B.n630 69.6791
R885 B.n630 B.n629 69.6791
R886 B.n629 B.n29 69.6791
R887 B.n623 B.n622 69.6791
R888 B.n622 B.n621 69.6791
R889 B.n621 B.n36 69.6791
R890 B.n615 B.n36 69.6791
R891 B.n615 B.n614 69.6791
R892 B.n614 B.n613 69.6791
R893 B.n613 B.n43 69.6791
R894 B.n607 B.n43 69.6791
R895 B.n607 B.n606 69.6791
R896 B.n606 B.n605 69.6791
R897 B.n605 B.n50 69.6791
R898 B.n599 B.n50 69.6791
R899 B.n598 B.n597 69.6791
R900 B.n597 B.n57 69.6791
R901 B.n591 B.n57 69.6791
R902 B.n591 B.n590 69.6791
R903 B.n590 B.n589 69.6791
R904 B.n589 B.n64 69.6791
R905 B.n583 B.n64 69.6791
R906 B.n583 B.n582 69.6791
R907 B.t1 B.n233 65.5804
R908 B.t2 B.n29 65.5804
R909 B.n311 B.n310 63.0308
R910 B.n309 B.n308 63.0308
R911 B.n101 B.n100 63.0308
R912 B.n98 B.n97 63.0308
R913 B.n352 B.n311 59.5399
R914 B.n373 B.n309 59.5399
R915 B.n102 B.n101 59.5399
R916 B.n99 B.n98 59.5399
R917 B.n447 B.t9 49.1854
R918 B.n599 B.t5 49.1854
R919 B.n507 B.t3 43.0373
R920 B.n18 B.t0 43.0373
R921 B.n104 B.n66 32.0005
R922 B.n578 B.n577 32.0005
R923 B.n420 B.n419 32.0005
R924 B.n414 B.n275 32.0005
R925 B.n514 B.t3 26.6423
R926 B.n645 B.t0 26.6423
R927 B.n265 B.t9 20.4942
R928 B.t5 B.n598 20.4942
R929 B B.n657 18.0485
R930 B.n105 B.n104 10.6151
R931 B.n108 B.n105 10.6151
R932 B.n109 B.n108 10.6151
R933 B.n112 B.n109 10.6151
R934 B.n113 B.n112 10.6151
R935 B.n116 B.n113 10.6151
R936 B.n117 B.n116 10.6151
R937 B.n120 B.n117 10.6151
R938 B.n121 B.n120 10.6151
R939 B.n124 B.n121 10.6151
R940 B.n125 B.n124 10.6151
R941 B.n128 B.n125 10.6151
R942 B.n129 B.n128 10.6151
R943 B.n132 B.n129 10.6151
R944 B.n133 B.n132 10.6151
R945 B.n136 B.n133 10.6151
R946 B.n137 B.n136 10.6151
R947 B.n140 B.n137 10.6151
R948 B.n141 B.n140 10.6151
R949 B.n144 B.n141 10.6151
R950 B.n145 B.n144 10.6151
R951 B.n149 B.n148 10.6151
R952 B.n152 B.n149 10.6151
R953 B.n153 B.n152 10.6151
R954 B.n156 B.n153 10.6151
R955 B.n157 B.n156 10.6151
R956 B.n160 B.n157 10.6151
R957 B.n161 B.n160 10.6151
R958 B.n164 B.n161 10.6151
R959 B.n165 B.n164 10.6151
R960 B.n169 B.n168 10.6151
R961 B.n172 B.n169 10.6151
R962 B.n173 B.n172 10.6151
R963 B.n176 B.n173 10.6151
R964 B.n177 B.n176 10.6151
R965 B.n180 B.n177 10.6151
R966 B.n181 B.n180 10.6151
R967 B.n184 B.n181 10.6151
R968 B.n185 B.n184 10.6151
R969 B.n188 B.n185 10.6151
R970 B.n189 B.n188 10.6151
R971 B.n192 B.n189 10.6151
R972 B.n193 B.n192 10.6151
R973 B.n196 B.n193 10.6151
R974 B.n197 B.n196 10.6151
R975 B.n200 B.n197 10.6151
R976 B.n201 B.n200 10.6151
R977 B.n204 B.n201 10.6151
R978 B.n206 B.n204 10.6151
R979 B.n207 B.n206 10.6151
R980 B.n578 B.n207 10.6151
R981 B.n421 B.n420 10.6151
R982 B.n421 B.n271 10.6151
R983 B.n431 B.n271 10.6151
R984 B.n432 B.n431 10.6151
R985 B.n433 B.n432 10.6151
R986 B.n433 B.n262 10.6151
R987 B.n443 B.n262 10.6151
R988 B.n444 B.n443 10.6151
R989 B.n445 B.n444 10.6151
R990 B.n445 B.n255 10.6151
R991 B.n455 B.n255 10.6151
R992 B.n456 B.n455 10.6151
R993 B.n457 B.n456 10.6151
R994 B.n457 B.n247 10.6151
R995 B.n467 B.n247 10.6151
R996 B.n468 B.n467 10.6151
R997 B.n469 B.n468 10.6151
R998 B.n469 B.n239 10.6151
R999 B.n479 B.n239 10.6151
R1000 B.n480 B.n479 10.6151
R1001 B.n481 B.n480 10.6151
R1002 B.n481 B.n231 10.6151
R1003 B.n491 B.n231 10.6151
R1004 B.n492 B.n491 10.6151
R1005 B.n493 B.n492 10.6151
R1006 B.n493 B.n223 10.6151
R1007 B.n503 B.n223 10.6151
R1008 B.n504 B.n503 10.6151
R1009 B.n505 B.n504 10.6151
R1010 B.n505 B.n216 10.6151
R1011 B.n516 B.n216 10.6151
R1012 B.n517 B.n516 10.6151
R1013 B.n519 B.n517 10.6151
R1014 B.n519 B.n518 10.6151
R1015 B.n518 B.n208 10.6151
R1016 B.n530 B.n208 10.6151
R1017 B.n531 B.n530 10.6151
R1018 B.n532 B.n531 10.6151
R1019 B.n533 B.n532 10.6151
R1020 B.n535 B.n533 10.6151
R1021 B.n536 B.n535 10.6151
R1022 B.n537 B.n536 10.6151
R1023 B.n538 B.n537 10.6151
R1024 B.n540 B.n538 10.6151
R1025 B.n541 B.n540 10.6151
R1026 B.n542 B.n541 10.6151
R1027 B.n543 B.n542 10.6151
R1028 B.n545 B.n543 10.6151
R1029 B.n546 B.n545 10.6151
R1030 B.n547 B.n546 10.6151
R1031 B.n548 B.n547 10.6151
R1032 B.n550 B.n548 10.6151
R1033 B.n551 B.n550 10.6151
R1034 B.n552 B.n551 10.6151
R1035 B.n553 B.n552 10.6151
R1036 B.n555 B.n553 10.6151
R1037 B.n556 B.n555 10.6151
R1038 B.n557 B.n556 10.6151
R1039 B.n558 B.n557 10.6151
R1040 B.n560 B.n558 10.6151
R1041 B.n561 B.n560 10.6151
R1042 B.n562 B.n561 10.6151
R1043 B.n563 B.n562 10.6151
R1044 B.n565 B.n563 10.6151
R1045 B.n566 B.n565 10.6151
R1046 B.n567 B.n566 10.6151
R1047 B.n568 B.n567 10.6151
R1048 B.n570 B.n568 10.6151
R1049 B.n571 B.n570 10.6151
R1050 B.n572 B.n571 10.6151
R1051 B.n573 B.n572 10.6151
R1052 B.n575 B.n573 10.6151
R1053 B.n576 B.n575 10.6151
R1054 B.n577 B.n576 10.6151
R1055 B.n414 B.n413 10.6151
R1056 B.n413 B.n412 10.6151
R1057 B.n412 B.n411 10.6151
R1058 B.n411 B.n409 10.6151
R1059 B.n409 B.n406 10.6151
R1060 B.n406 B.n405 10.6151
R1061 B.n405 B.n402 10.6151
R1062 B.n402 B.n401 10.6151
R1063 B.n401 B.n398 10.6151
R1064 B.n398 B.n397 10.6151
R1065 B.n397 B.n394 10.6151
R1066 B.n394 B.n393 10.6151
R1067 B.n393 B.n390 10.6151
R1068 B.n390 B.n389 10.6151
R1069 B.n389 B.n386 10.6151
R1070 B.n386 B.n385 10.6151
R1071 B.n385 B.n382 10.6151
R1072 B.n382 B.n381 10.6151
R1073 B.n381 B.n378 10.6151
R1074 B.n378 B.n377 10.6151
R1075 B.n377 B.n374 10.6151
R1076 B.n372 B.n369 10.6151
R1077 B.n369 B.n368 10.6151
R1078 B.n368 B.n365 10.6151
R1079 B.n365 B.n364 10.6151
R1080 B.n364 B.n361 10.6151
R1081 B.n361 B.n360 10.6151
R1082 B.n360 B.n357 10.6151
R1083 B.n357 B.n356 10.6151
R1084 B.n356 B.n353 10.6151
R1085 B.n351 B.n348 10.6151
R1086 B.n348 B.n347 10.6151
R1087 B.n347 B.n344 10.6151
R1088 B.n344 B.n343 10.6151
R1089 B.n343 B.n340 10.6151
R1090 B.n340 B.n339 10.6151
R1091 B.n339 B.n336 10.6151
R1092 B.n336 B.n335 10.6151
R1093 B.n335 B.n332 10.6151
R1094 B.n332 B.n331 10.6151
R1095 B.n331 B.n328 10.6151
R1096 B.n328 B.n327 10.6151
R1097 B.n327 B.n324 10.6151
R1098 B.n324 B.n323 10.6151
R1099 B.n323 B.n320 10.6151
R1100 B.n320 B.n319 10.6151
R1101 B.n319 B.n316 10.6151
R1102 B.n316 B.n315 10.6151
R1103 B.n315 B.n312 10.6151
R1104 B.n312 B.n279 10.6151
R1105 B.n419 B.n279 10.6151
R1106 B.n425 B.n275 10.6151
R1107 B.n426 B.n425 10.6151
R1108 B.n427 B.n426 10.6151
R1109 B.n427 B.n267 10.6151
R1110 B.n437 B.n267 10.6151
R1111 B.n438 B.n437 10.6151
R1112 B.n439 B.n438 10.6151
R1113 B.n439 B.n259 10.6151
R1114 B.n449 B.n259 10.6151
R1115 B.n450 B.n449 10.6151
R1116 B.n451 B.n450 10.6151
R1117 B.n451 B.n251 10.6151
R1118 B.n461 B.n251 10.6151
R1119 B.n462 B.n461 10.6151
R1120 B.n463 B.n462 10.6151
R1121 B.n463 B.n243 10.6151
R1122 B.n473 B.n243 10.6151
R1123 B.n474 B.n473 10.6151
R1124 B.n475 B.n474 10.6151
R1125 B.n475 B.n235 10.6151
R1126 B.n485 B.n235 10.6151
R1127 B.n486 B.n485 10.6151
R1128 B.n487 B.n486 10.6151
R1129 B.n487 B.n227 10.6151
R1130 B.n497 B.n227 10.6151
R1131 B.n498 B.n497 10.6151
R1132 B.n499 B.n498 10.6151
R1133 B.n499 B.n219 10.6151
R1134 B.n510 B.n219 10.6151
R1135 B.n511 B.n510 10.6151
R1136 B.n512 B.n511 10.6151
R1137 B.n512 B.n212 10.6151
R1138 B.n523 B.n212 10.6151
R1139 B.n524 B.n523 10.6151
R1140 B.n525 B.n524 10.6151
R1141 B.n525 B.n0 10.6151
R1142 B.n651 B.n1 10.6151
R1143 B.n651 B.n650 10.6151
R1144 B.n650 B.n649 10.6151
R1145 B.n649 B.n10 10.6151
R1146 B.n643 B.n10 10.6151
R1147 B.n643 B.n642 10.6151
R1148 B.n642 B.n641 10.6151
R1149 B.n641 B.n16 10.6151
R1150 B.n635 B.n16 10.6151
R1151 B.n635 B.n634 10.6151
R1152 B.n634 B.n633 10.6151
R1153 B.n633 B.n24 10.6151
R1154 B.n627 B.n24 10.6151
R1155 B.n627 B.n626 10.6151
R1156 B.n626 B.n625 10.6151
R1157 B.n625 B.n31 10.6151
R1158 B.n619 B.n31 10.6151
R1159 B.n619 B.n618 10.6151
R1160 B.n618 B.n617 10.6151
R1161 B.n617 B.n38 10.6151
R1162 B.n611 B.n38 10.6151
R1163 B.n611 B.n610 10.6151
R1164 B.n610 B.n609 10.6151
R1165 B.n609 B.n45 10.6151
R1166 B.n603 B.n45 10.6151
R1167 B.n603 B.n602 10.6151
R1168 B.n602 B.n601 10.6151
R1169 B.n601 B.n52 10.6151
R1170 B.n595 B.n52 10.6151
R1171 B.n595 B.n594 10.6151
R1172 B.n594 B.n593 10.6151
R1173 B.n593 B.n59 10.6151
R1174 B.n587 B.n59 10.6151
R1175 B.n587 B.n586 10.6151
R1176 B.n586 B.n585 10.6151
R1177 B.n585 B.n66 10.6151
R1178 B.n145 B.n102 9.36635
R1179 B.n168 B.n99 9.36635
R1180 B.n374 B.n373 9.36635
R1181 B.n352 B.n351 9.36635
R1182 B.n483 B.t1 4.09924
R1183 B.n623 B.t2 4.09924
R1184 B.n657 B.n0 2.81026
R1185 B.n657 B.n1 2.81026
R1186 B.n148 B.n102 1.24928
R1187 B.n165 B.n99 1.24928
R1188 B.n373 B.n372 1.24928
R1189 B.n353 B.n352 1.24928
R1190 VN.n1 VN.t2 79.4665
R1191 VN.n0 VN.t3 79.4665
R1192 VN.n0 VN.t0 78.4926
R1193 VN.n1 VN.t1 78.4926
R1194 VN VN.n1 45.6332
R1195 VN VN.n0 3.14452
R1196 VDD2.n2 VDD2.n0 107.284
R1197 VDD2.n2 VDD2.n1 70.4568
R1198 VDD2.n1 VDD2.t2 3.62687
R1199 VDD2.n1 VDD2.t1 3.62687
R1200 VDD2.n0 VDD2.t0 3.62687
R1201 VDD2.n0 VDD2.t3 3.62687
R1202 VDD2 VDD2.n2 0.0586897
C0 VTAIL VP 2.78359f
C1 VN VDD2 2.37919f
C2 VDD2 VP 0.418966f
C3 VDD2 VTAIL 4.03767f
C4 VN VDD1 0.149763f
C5 VDD1 VP 2.64373f
C6 VTAIL VDD1 3.98132f
C7 VN VP 5.21057f
C8 VN VTAIL 2.76948f
C9 VDD2 VDD1 1.10274f
C10 VDD2 B 3.444242f
C11 VDD1 B 7.08291f
C12 VTAIL B 6.03513f
C13 VN B 10.75654f
C14 VP B 9.048218f
C15 VDD2.t0 B 0.120276f
C16 VDD2.t3 B 0.120276f
C17 VDD2.n0 B 1.4473f
C18 VDD2.t2 B 0.120276f
C19 VDD2.t1 B 0.120276f
C20 VDD2.n1 B 1.00323f
C21 VDD2.n2 B 3.2107f
C22 VN.t0 B 1.41295f
C23 VN.t3 B 1.42049f
C24 VN.n0 B 0.870618f
C25 VN.t2 B 1.42049f
C26 VN.t1 B 1.41295f
C27 VN.n1 B 2.25265f
C28 VTAIL.t0 B 0.881158f
C29 VTAIL.n0 B 0.357073f
C30 VTAIL.t5 B 0.881158f
C31 VTAIL.n1 B 0.446028f
C32 VTAIL.t7 B 0.881158f
C33 VTAIL.n2 B 1.19166f
C34 VTAIL.t1 B 0.881158f
C35 VTAIL.n3 B 1.19166f
C36 VTAIL.t3 B 0.881158f
C37 VTAIL.n4 B 0.446027f
C38 VTAIL.t4 B 0.881158f
C39 VTAIL.n5 B 0.446027f
C40 VTAIL.t6 B 0.881154f
C41 VTAIL.n6 B 1.19166f
C42 VTAIL.t2 B 0.881158f
C43 VTAIL.n7 B 1.09499f
C44 VDD1.t3 B 0.122071f
C45 VDD1.t0 B 0.122071f
C46 VDD1.n0 B 1.0186f
C47 VDD1.t2 B 0.122071f
C48 VDD1.t1 B 0.122071f
C49 VDD1.n1 B 1.49278f
C50 VP.t2 B 1.17747f
C51 VP.n0 B 0.548246f
C52 VP.n1 B 0.028067f
C53 VP.n2 B 0.040799f
C54 VP.n3 B 0.045292f
C55 VP.t0 B 1.17747f
C56 VP.t3 B 1.4532f
C57 VP.t1 B 1.44548f
C58 VP.n4 B 2.29276f
C59 VP.n5 B 1.36635f
C60 VP.n6 B 0.548246f
C61 VP.n7 B 0.045624f
C62 VP.n8 B 0.052047f
C63 VP.n9 B 0.028067f
C64 VP.n10 B 0.028067f
C65 VP.n11 B 0.028067f
C66 VP.n12 B 0.040799f
C67 VP.n13 B 0.052047f
C68 VP.n14 B 0.045624f
C69 VP.n15 B 0.045292f
C70 VP.n16 B 0.059595f
.ends

