* NGSPICE file created from diff_pair_sample_0966.ext - technology: sky130A

.subckt diff_pair_sample_0966 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t1 w_n1422_n1224# sky130_fd_pr__pfet_01v8 ad=0.4914 pd=3.3 as=0.4914 ps=3.3 w=1.26 l=0.8
X1 B.t11 B.t9 B.t10 w_n1422_n1224# sky130_fd_pr__pfet_01v8 ad=0.4914 pd=3.3 as=0 ps=0 w=1.26 l=0.8
X2 B.t8 B.t6 B.t7 w_n1422_n1224# sky130_fd_pr__pfet_01v8 ad=0.4914 pd=3.3 as=0 ps=0 w=1.26 l=0.8
X3 B.t5 B.t3 B.t4 w_n1422_n1224# sky130_fd_pr__pfet_01v8 ad=0.4914 pd=3.3 as=0 ps=0 w=1.26 l=0.8
X4 B.t2 B.t0 B.t1 w_n1422_n1224# sky130_fd_pr__pfet_01v8 ad=0.4914 pd=3.3 as=0 ps=0 w=1.26 l=0.8
X5 VDD2.t1 VN.t0 VTAIL.t3 w_n1422_n1224# sky130_fd_pr__pfet_01v8 ad=0.4914 pd=3.3 as=0.4914 ps=3.3 w=1.26 l=0.8
X6 VDD2.t0 VN.t1 VTAIL.t0 w_n1422_n1224# sky130_fd_pr__pfet_01v8 ad=0.4914 pd=3.3 as=0.4914 ps=3.3 w=1.26 l=0.8
X7 VDD1.t0 VP.t1 VTAIL.t2 w_n1422_n1224# sky130_fd_pr__pfet_01v8 ad=0.4914 pd=3.3 as=0.4914 ps=3.3 w=1.26 l=0.8
R0 VP.n0 VP.t0 280.123
R1 VP.n0 VP.t1 248.362
R2 VP VP.n0 0.0516364
R3 VTAIL.n3 VTAIL.t3 372.312
R4 VTAIL.n0 VTAIL.t2 372.312
R5 VTAIL.n2 VTAIL.t1 372.312
R6 VTAIL.n1 VTAIL.t0 372.312
R7 VTAIL.n1 VTAIL.n0 15.4186
R8 VTAIL.n3 VTAIL.n2 14.4445
R9 VTAIL.n2 VTAIL.n1 0.957397
R10 VTAIL VTAIL.n0 0.772052
R11 VTAIL VTAIL.n3 0.185845
R12 VDD1 VDD1.t0 416.471
R13 VDD1 VDD1.t1 389.293
R14 B.n135 B.n134 585
R15 B.n133 B.n44 585
R16 B.n132 B.n131 585
R17 B.n130 B.n45 585
R18 B.n129 B.n128 585
R19 B.n127 B.n46 585
R20 B.n126 B.n125 585
R21 B.n124 B.n47 585
R22 B.n123 B.n122 585
R23 B.n121 B.n48 585
R24 B.n120 B.n119 585
R25 B.n115 B.n49 585
R26 B.n114 B.n113 585
R27 B.n112 B.n50 585
R28 B.n111 B.n110 585
R29 B.n109 B.n51 585
R30 B.n108 B.n107 585
R31 B.n106 B.n52 585
R32 B.n105 B.n104 585
R33 B.n103 B.n53 585
R34 B.n101 B.n100 585
R35 B.n99 B.n56 585
R36 B.n98 B.n97 585
R37 B.n96 B.n57 585
R38 B.n95 B.n94 585
R39 B.n93 B.n58 585
R40 B.n92 B.n91 585
R41 B.n90 B.n59 585
R42 B.n89 B.n88 585
R43 B.n87 B.n60 585
R44 B.n136 B.n43 585
R45 B.n138 B.n137 585
R46 B.n139 B.n42 585
R47 B.n141 B.n140 585
R48 B.n142 B.n41 585
R49 B.n144 B.n143 585
R50 B.n145 B.n40 585
R51 B.n147 B.n146 585
R52 B.n148 B.n39 585
R53 B.n150 B.n149 585
R54 B.n151 B.n38 585
R55 B.n153 B.n152 585
R56 B.n154 B.n37 585
R57 B.n156 B.n155 585
R58 B.n157 B.n36 585
R59 B.n159 B.n158 585
R60 B.n160 B.n35 585
R61 B.n162 B.n161 585
R62 B.n163 B.n34 585
R63 B.n165 B.n164 585
R64 B.n166 B.n33 585
R65 B.n168 B.n167 585
R66 B.n169 B.n32 585
R67 B.n171 B.n170 585
R68 B.n172 B.n31 585
R69 B.n174 B.n173 585
R70 B.n175 B.n30 585
R71 B.n177 B.n176 585
R72 B.n178 B.n29 585
R73 B.n180 B.n179 585
R74 B.n226 B.n9 585
R75 B.n225 B.n224 585
R76 B.n223 B.n10 585
R77 B.n222 B.n221 585
R78 B.n220 B.n11 585
R79 B.n219 B.n218 585
R80 B.n217 B.n12 585
R81 B.n216 B.n215 585
R82 B.n214 B.n13 585
R83 B.n213 B.n212 585
R84 B.n211 B.n210 585
R85 B.n209 B.n17 585
R86 B.n208 B.n207 585
R87 B.n206 B.n18 585
R88 B.n205 B.n204 585
R89 B.n203 B.n19 585
R90 B.n202 B.n201 585
R91 B.n200 B.n20 585
R92 B.n199 B.n198 585
R93 B.n197 B.n21 585
R94 B.n195 B.n194 585
R95 B.n193 B.n24 585
R96 B.n192 B.n191 585
R97 B.n190 B.n25 585
R98 B.n189 B.n188 585
R99 B.n187 B.n26 585
R100 B.n186 B.n185 585
R101 B.n184 B.n27 585
R102 B.n183 B.n182 585
R103 B.n181 B.n28 585
R104 B.n228 B.n227 585
R105 B.n229 B.n8 585
R106 B.n231 B.n230 585
R107 B.n232 B.n7 585
R108 B.n234 B.n233 585
R109 B.n235 B.n6 585
R110 B.n237 B.n236 585
R111 B.n238 B.n5 585
R112 B.n240 B.n239 585
R113 B.n241 B.n4 585
R114 B.n243 B.n242 585
R115 B.n244 B.n3 585
R116 B.n246 B.n245 585
R117 B.n247 B.n0 585
R118 B.n2 B.n1 585
R119 B.n68 B.n67 585
R120 B.n69 B.n66 585
R121 B.n71 B.n70 585
R122 B.n72 B.n65 585
R123 B.n74 B.n73 585
R124 B.n75 B.n64 585
R125 B.n77 B.n76 585
R126 B.n78 B.n63 585
R127 B.n80 B.n79 585
R128 B.n81 B.n62 585
R129 B.n83 B.n82 585
R130 B.n84 B.n61 585
R131 B.n86 B.n85 585
R132 B.n87 B.n86 521.33
R133 B.n134 B.n43 521.33
R134 B.n181 B.n180 521.33
R135 B.n228 B.n9 521.33
R136 B.n54 B.t4 388.156
R137 B.n116 B.t7 388.156
R138 B.n22 B.t2 388.156
R139 B.n14 B.t11 388.156
R140 B.n55 B.t5 366.241
R141 B.n117 B.t8 366.241
R142 B.n23 B.t1 366.241
R143 B.n15 B.t10 366.241
R144 B.n249 B.n248 256.663
R145 B.n54 B.t3 239.846
R146 B.n116 B.t6 239.846
R147 B.n22 B.t0 239.846
R148 B.n14 B.t9 239.846
R149 B.n248 B.n247 235.042
R150 B.n248 B.n2 235.042
R151 B.n88 B.n87 163.367
R152 B.n88 B.n59 163.367
R153 B.n92 B.n59 163.367
R154 B.n93 B.n92 163.367
R155 B.n94 B.n93 163.367
R156 B.n94 B.n57 163.367
R157 B.n98 B.n57 163.367
R158 B.n99 B.n98 163.367
R159 B.n100 B.n99 163.367
R160 B.n100 B.n53 163.367
R161 B.n105 B.n53 163.367
R162 B.n106 B.n105 163.367
R163 B.n107 B.n106 163.367
R164 B.n107 B.n51 163.367
R165 B.n111 B.n51 163.367
R166 B.n112 B.n111 163.367
R167 B.n113 B.n112 163.367
R168 B.n113 B.n49 163.367
R169 B.n120 B.n49 163.367
R170 B.n121 B.n120 163.367
R171 B.n122 B.n121 163.367
R172 B.n122 B.n47 163.367
R173 B.n126 B.n47 163.367
R174 B.n127 B.n126 163.367
R175 B.n128 B.n127 163.367
R176 B.n128 B.n45 163.367
R177 B.n132 B.n45 163.367
R178 B.n133 B.n132 163.367
R179 B.n134 B.n133 163.367
R180 B.n180 B.n29 163.367
R181 B.n176 B.n29 163.367
R182 B.n176 B.n175 163.367
R183 B.n175 B.n174 163.367
R184 B.n174 B.n31 163.367
R185 B.n170 B.n31 163.367
R186 B.n170 B.n169 163.367
R187 B.n169 B.n168 163.367
R188 B.n168 B.n33 163.367
R189 B.n164 B.n33 163.367
R190 B.n164 B.n163 163.367
R191 B.n163 B.n162 163.367
R192 B.n162 B.n35 163.367
R193 B.n158 B.n35 163.367
R194 B.n158 B.n157 163.367
R195 B.n157 B.n156 163.367
R196 B.n156 B.n37 163.367
R197 B.n152 B.n37 163.367
R198 B.n152 B.n151 163.367
R199 B.n151 B.n150 163.367
R200 B.n150 B.n39 163.367
R201 B.n146 B.n39 163.367
R202 B.n146 B.n145 163.367
R203 B.n145 B.n144 163.367
R204 B.n144 B.n41 163.367
R205 B.n140 B.n41 163.367
R206 B.n140 B.n139 163.367
R207 B.n139 B.n138 163.367
R208 B.n138 B.n43 163.367
R209 B.n224 B.n9 163.367
R210 B.n224 B.n223 163.367
R211 B.n223 B.n222 163.367
R212 B.n222 B.n11 163.367
R213 B.n218 B.n11 163.367
R214 B.n218 B.n217 163.367
R215 B.n217 B.n216 163.367
R216 B.n216 B.n13 163.367
R217 B.n212 B.n13 163.367
R218 B.n212 B.n211 163.367
R219 B.n211 B.n17 163.367
R220 B.n207 B.n17 163.367
R221 B.n207 B.n206 163.367
R222 B.n206 B.n205 163.367
R223 B.n205 B.n19 163.367
R224 B.n201 B.n19 163.367
R225 B.n201 B.n200 163.367
R226 B.n200 B.n199 163.367
R227 B.n199 B.n21 163.367
R228 B.n194 B.n21 163.367
R229 B.n194 B.n193 163.367
R230 B.n193 B.n192 163.367
R231 B.n192 B.n25 163.367
R232 B.n188 B.n25 163.367
R233 B.n188 B.n187 163.367
R234 B.n187 B.n186 163.367
R235 B.n186 B.n27 163.367
R236 B.n182 B.n27 163.367
R237 B.n182 B.n181 163.367
R238 B.n229 B.n228 163.367
R239 B.n230 B.n229 163.367
R240 B.n230 B.n7 163.367
R241 B.n234 B.n7 163.367
R242 B.n235 B.n234 163.367
R243 B.n236 B.n235 163.367
R244 B.n236 B.n5 163.367
R245 B.n240 B.n5 163.367
R246 B.n241 B.n240 163.367
R247 B.n242 B.n241 163.367
R248 B.n242 B.n3 163.367
R249 B.n246 B.n3 163.367
R250 B.n247 B.n246 163.367
R251 B.n68 B.n2 163.367
R252 B.n69 B.n68 163.367
R253 B.n70 B.n69 163.367
R254 B.n70 B.n65 163.367
R255 B.n74 B.n65 163.367
R256 B.n75 B.n74 163.367
R257 B.n76 B.n75 163.367
R258 B.n76 B.n63 163.367
R259 B.n80 B.n63 163.367
R260 B.n81 B.n80 163.367
R261 B.n82 B.n81 163.367
R262 B.n82 B.n61 163.367
R263 B.n86 B.n61 163.367
R264 B.n102 B.n55 59.5399
R265 B.n118 B.n117 59.5399
R266 B.n196 B.n23 59.5399
R267 B.n16 B.n15 59.5399
R268 B.n227 B.n226 33.8737
R269 B.n179 B.n28 33.8737
R270 B.n136 B.n135 33.8737
R271 B.n85 B.n60 33.8737
R272 B.n55 B.n54 21.9157
R273 B.n117 B.n116 21.9157
R274 B.n23 B.n22 21.9157
R275 B.n15 B.n14 21.9157
R276 B B.n249 18.0485
R277 B.n227 B.n8 10.6151
R278 B.n231 B.n8 10.6151
R279 B.n232 B.n231 10.6151
R280 B.n233 B.n232 10.6151
R281 B.n233 B.n6 10.6151
R282 B.n237 B.n6 10.6151
R283 B.n238 B.n237 10.6151
R284 B.n239 B.n238 10.6151
R285 B.n239 B.n4 10.6151
R286 B.n243 B.n4 10.6151
R287 B.n244 B.n243 10.6151
R288 B.n245 B.n244 10.6151
R289 B.n245 B.n0 10.6151
R290 B.n226 B.n225 10.6151
R291 B.n225 B.n10 10.6151
R292 B.n221 B.n10 10.6151
R293 B.n221 B.n220 10.6151
R294 B.n220 B.n219 10.6151
R295 B.n219 B.n12 10.6151
R296 B.n215 B.n12 10.6151
R297 B.n215 B.n214 10.6151
R298 B.n214 B.n213 10.6151
R299 B.n210 B.n209 10.6151
R300 B.n209 B.n208 10.6151
R301 B.n208 B.n18 10.6151
R302 B.n204 B.n18 10.6151
R303 B.n204 B.n203 10.6151
R304 B.n203 B.n202 10.6151
R305 B.n202 B.n20 10.6151
R306 B.n198 B.n20 10.6151
R307 B.n198 B.n197 10.6151
R308 B.n195 B.n24 10.6151
R309 B.n191 B.n24 10.6151
R310 B.n191 B.n190 10.6151
R311 B.n190 B.n189 10.6151
R312 B.n189 B.n26 10.6151
R313 B.n185 B.n26 10.6151
R314 B.n185 B.n184 10.6151
R315 B.n184 B.n183 10.6151
R316 B.n183 B.n28 10.6151
R317 B.n179 B.n178 10.6151
R318 B.n178 B.n177 10.6151
R319 B.n177 B.n30 10.6151
R320 B.n173 B.n30 10.6151
R321 B.n173 B.n172 10.6151
R322 B.n172 B.n171 10.6151
R323 B.n171 B.n32 10.6151
R324 B.n167 B.n32 10.6151
R325 B.n167 B.n166 10.6151
R326 B.n166 B.n165 10.6151
R327 B.n165 B.n34 10.6151
R328 B.n161 B.n34 10.6151
R329 B.n161 B.n160 10.6151
R330 B.n160 B.n159 10.6151
R331 B.n159 B.n36 10.6151
R332 B.n155 B.n36 10.6151
R333 B.n155 B.n154 10.6151
R334 B.n154 B.n153 10.6151
R335 B.n153 B.n38 10.6151
R336 B.n149 B.n38 10.6151
R337 B.n149 B.n148 10.6151
R338 B.n148 B.n147 10.6151
R339 B.n147 B.n40 10.6151
R340 B.n143 B.n40 10.6151
R341 B.n143 B.n142 10.6151
R342 B.n142 B.n141 10.6151
R343 B.n141 B.n42 10.6151
R344 B.n137 B.n42 10.6151
R345 B.n137 B.n136 10.6151
R346 B.n67 B.n1 10.6151
R347 B.n67 B.n66 10.6151
R348 B.n71 B.n66 10.6151
R349 B.n72 B.n71 10.6151
R350 B.n73 B.n72 10.6151
R351 B.n73 B.n64 10.6151
R352 B.n77 B.n64 10.6151
R353 B.n78 B.n77 10.6151
R354 B.n79 B.n78 10.6151
R355 B.n79 B.n62 10.6151
R356 B.n83 B.n62 10.6151
R357 B.n84 B.n83 10.6151
R358 B.n85 B.n84 10.6151
R359 B.n89 B.n60 10.6151
R360 B.n90 B.n89 10.6151
R361 B.n91 B.n90 10.6151
R362 B.n91 B.n58 10.6151
R363 B.n95 B.n58 10.6151
R364 B.n96 B.n95 10.6151
R365 B.n97 B.n96 10.6151
R366 B.n97 B.n56 10.6151
R367 B.n101 B.n56 10.6151
R368 B.n104 B.n103 10.6151
R369 B.n104 B.n52 10.6151
R370 B.n108 B.n52 10.6151
R371 B.n109 B.n108 10.6151
R372 B.n110 B.n109 10.6151
R373 B.n110 B.n50 10.6151
R374 B.n114 B.n50 10.6151
R375 B.n115 B.n114 10.6151
R376 B.n119 B.n115 10.6151
R377 B.n123 B.n48 10.6151
R378 B.n124 B.n123 10.6151
R379 B.n125 B.n124 10.6151
R380 B.n125 B.n46 10.6151
R381 B.n129 B.n46 10.6151
R382 B.n130 B.n129 10.6151
R383 B.n131 B.n130 10.6151
R384 B.n131 B.n44 10.6151
R385 B.n135 B.n44 10.6151
R386 B.n213 B.n16 8.74196
R387 B.n196 B.n195 8.74196
R388 B.n102 B.n101 8.74196
R389 B.n118 B.n48 8.74196
R390 B.n249 B.n0 8.11757
R391 B.n249 B.n1 8.11757
R392 B.n210 B.n16 1.87367
R393 B.n197 B.n196 1.87367
R394 B.n103 B.n102 1.87367
R395 B.n119 B.n118 1.87367
R396 VN VN.t1 280.503
R397 VN VN.t0 248.412
R398 VDD2.n0 VDD2.t1 415.702
R399 VDD2.n0 VDD2.t0 388.99
R400 VDD2 VDD2.n0 0.302224
C0 VP B 0.875633f
C1 VN B 0.592535f
C2 B VTAIL 0.742166f
C3 w_n1422_n1224# VDD2 0.789933f
C4 VDD1 B 0.64401f
C5 VP w_n1422_n1224# 1.72337f
C6 VN w_n1422_n1224# 1.55301f
C7 w_n1422_n1224# VTAIL 1.07091f
C8 w_n1422_n1224# VDD1 0.78522f
C9 VP VDD2 0.266192f
C10 VN VDD2 0.433701f
C11 VDD2 VTAIL 1.74805f
C12 VP VN 2.62435f
C13 VP VTAIL 0.553357f
C14 VDD1 VDD2 0.469029f
C15 VN VTAIL 0.539201f
C16 w_n1422_n1224# B 3.83889f
C17 VP VDD1 0.542026f
C18 VN VDD1 0.156341f
C19 VDD1 VTAIL 1.70749f
C20 B VDD2 0.659471f
C21 VDD2 VSUBS 0.334253f
C22 VDD1 VSUBS 0.489567f
C23 VTAIL VSUBS 0.201852f
C24 VN VSUBS 3.27698f
C25 VP VSUBS 0.655447f
C26 B VSUBS 1.583461f
C27 w_n1422_n1224# VSUBS 22.370901f
C28 VN.t0 VSUBS 0.205158f
C29 VN.t1 VSUBS 0.327764f
C30 B.n0 VSUBS 0.008828f
C31 B.n1 VSUBS 0.008828f
C32 B.n2 VSUBS 0.013057f
C33 B.n3 VSUBS 0.010006f
C34 B.n4 VSUBS 0.010006f
C35 B.n5 VSUBS 0.010006f
C36 B.n6 VSUBS 0.010006f
C37 B.n7 VSUBS 0.010006f
C38 B.n8 VSUBS 0.010006f
C39 B.n9 VSUBS 0.024887f
C40 B.n10 VSUBS 0.010006f
C41 B.n11 VSUBS 0.010006f
C42 B.n12 VSUBS 0.010006f
C43 B.n13 VSUBS 0.010006f
C44 B.t10 VSUBS 0.034017f
C45 B.t11 VSUBS 0.036705f
C46 B.t9 VSUBS 0.071912f
C47 B.n14 VSUBS 0.066564f
C48 B.n15 VSUBS 0.06189f
C49 B.n16 VSUBS 0.023182f
C50 B.n17 VSUBS 0.010006f
C51 B.n18 VSUBS 0.010006f
C52 B.n19 VSUBS 0.010006f
C53 B.n20 VSUBS 0.010006f
C54 B.n21 VSUBS 0.010006f
C55 B.t1 VSUBS 0.034017f
C56 B.t2 VSUBS 0.036705f
C57 B.t0 VSUBS 0.071912f
C58 B.n22 VSUBS 0.066564f
C59 B.n23 VSUBS 0.06189f
C60 B.n24 VSUBS 0.010006f
C61 B.n25 VSUBS 0.010006f
C62 B.n26 VSUBS 0.010006f
C63 B.n27 VSUBS 0.010006f
C64 B.n28 VSUBS 0.024887f
C65 B.n29 VSUBS 0.010006f
C66 B.n30 VSUBS 0.010006f
C67 B.n31 VSUBS 0.010006f
C68 B.n32 VSUBS 0.010006f
C69 B.n33 VSUBS 0.010006f
C70 B.n34 VSUBS 0.010006f
C71 B.n35 VSUBS 0.010006f
C72 B.n36 VSUBS 0.010006f
C73 B.n37 VSUBS 0.010006f
C74 B.n38 VSUBS 0.010006f
C75 B.n39 VSUBS 0.010006f
C76 B.n40 VSUBS 0.010006f
C77 B.n41 VSUBS 0.010006f
C78 B.n42 VSUBS 0.010006f
C79 B.n43 VSUBS 0.02308f
C80 B.n44 VSUBS 0.010006f
C81 B.n45 VSUBS 0.010006f
C82 B.n46 VSUBS 0.010006f
C83 B.n47 VSUBS 0.010006f
C84 B.n48 VSUBS 0.009123f
C85 B.n49 VSUBS 0.010006f
C86 B.n50 VSUBS 0.010006f
C87 B.n51 VSUBS 0.010006f
C88 B.n52 VSUBS 0.010006f
C89 B.n53 VSUBS 0.010006f
C90 B.t5 VSUBS 0.034017f
C91 B.t4 VSUBS 0.036705f
C92 B.t3 VSUBS 0.071912f
C93 B.n54 VSUBS 0.066564f
C94 B.n55 VSUBS 0.06189f
C95 B.n56 VSUBS 0.010006f
C96 B.n57 VSUBS 0.010006f
C97 B.n58 VSUBS 0.010006f
C98 B.n59 VSUBS 0.010006f
C99 B.n60 VSUBS 0.024887f
C100 B.n61 VSUBS 0.010006f
C101 B.n62 VSUBS 0.010006f
C102 B.n63 VSUBS 0.010006f
C103 B.n64 VSUBS 0.010006f
C104 B.n65 VSUBS 0.010006f
C105 B.n66 VSUBS 0.010006f
C106 B.n67 VSUBS 0.010006f
C107 B.n68 VSUBS 0.010006f
C108 B.n69 VSUBS 0.010006f
C109 B.n70 VSUBS 0.010006f
C110 B.n71 VSUBS 0.010006f
C111 B.n72 VSUBS 0.010006f
C112 B.n73 VSUBS 0.010006f
C113 B.n74 VSUBS 0.010006f
C114 B.n75 VSUBS 0.010006f
C115 B.n76 VSUBS 0.010006f
C116 B.n77 VSUBS 0.010006f
C117 B.n78 VSUBS 0.010006f
C118 B.n79 VSUBS 0.010006f
C119 B.n80 VSUBS 0.010006f
C120 B.n81 VSUBS 0.010006f
C121 B.n82 VSUBS 0.010006f
C122 B.n83 VSUBS 0.010006f
C123 B.n84 VSUBS 0.010006f
C124 B.n85 VSUBS 0.02308f
C125 B.n86 VSUBS 0.02308f
C126 B.n87 VSUBS 0.024887f
C127 B.n88 VSUBS 0.010006f
C128 B.n89 VSUBS 0.010006f
C129 B.n90 VSUBS 0.010006f
C130 B.n91 VSUBS 0.010006f
C131 B.n92 VSUBS 0.010006f
C132 B.n93 VSUBS 0.010006f
C133 B.n94 VSUBS 0.010006f
C134 B.n95 VSUBS 0.010006f
C135 B.n96 VSUBS 0.010006f
C136 B.n97 VSUBS 0.010006f
C137 B.n98 VSUBS 0.010006f
C138 B.n99 VSUBS 0.010006f
C139 B.n100 VSUBS 0.010006f
C140 B.n101 VSUBS 0.009123f
C141 B.n102 VSUBS 0.023182f
C142 B.n103 VSUBS 0.005886f
C143 B.n104 VSUBS 0.010006f
C144 B.n105 VSUBS 0.010006f
C145 B.n106 VSUBS 0.010006f
C146 B.n107 VSUBS 0.010006f
C147 B.n108 VSUBS 0.010006f
C148 B.n109 VSUBS 0.010006f
C149 B.n110 VSUBS 0.010006f
C150 B.n111 VSUBS 0.010006f
C151 B.n112 VSUBS 0.010006f
C152 B.n113 VSUBS 0.010006f
C153 B.n114 VSUBS 0.010006f
C154 B.n115 VSUBS 0.010006f
C155 B.t8 VSUBS 0.034017f
C156 B.t7 VSUBS 0.036705f
C157 B.t6 VSUBS 0.071912f
C158 B.n116 VSUBS 0.066564f
C159 B.n117 VSUBS 0.06189f
C160 B.n118 VSUBS 0.023182f
C161 B.n119 VSUBS 0.005886f
C162 B.n120 VSUBS 0.010006f
C163 B.n121 VSUBS 0.010006f
C164 B.n122 VSUBS 0.010006f
C165 B.n123 VSUBS 0.010006f
C166 B.n124 VSUBS 0.010006f
C167 B.n125 VSUBS 0.010006f
C168 B.n126 VSUBS 0.010006f
C169 B.n127 VSUBS 0.010006f
C170 B.n128 VSUBS 0.010006f
C171 B.n129 VSUBS 0.010006f
C172 B.n130 VSUBS 0.010006f
C173 B.n131 VSUBS 0.010006f
C174 B.n132 VSUBS 0.010006f
C175 B.n133 VSUBS 0.010006f
C176 B.n134 VSUBS 0.024887f
C177 B.n135 VSUBS 0.023748f
C178 B.n136 VSUBS 0.02422f
C179 B.n137 VSUBS 0.010006f
C180 B.n138 VSUBS 0.010006f
C181 B.n139 VSUBS 0.010006f
C182 B.n140 VSUBS 0.010006f
C183 B.n141 VSUBS 0.010006f
C184 B.n142 VSUBS 0.010006f
C185 B.n143 VSUBS 0.010006f
C186 B.n144 VSUBS 0.010006f
C187 B.n145 VSUBS 0.010006f
C188 B.n146 VSUBS 0.010006f
C189 B.n147 VSUBS 0.010006f
C190 B.n148 VSUBS 0.010006f
C191 B.n149 VSUBS 0.010006f
C192 B.n150 VSUBS 0.010006f
C193 B.n151 VSUBS 0.010006f
C194 B.n152 VSUBS 0.010006f
C195 B.n153 VSUBS 0.010006f
C196 B.n154 VSUBS 0.010006f
C197 B.n155 VSUBS 0.010006f
C198 B.n156 VSUBS 0.010006f
C199 B.n157 VSUBS 0.010006f
C200 B.n158 VSUBS 0.010006f
C201 B.n159 VSUBS 0.010006f
C202 B.n160 VSUBS 0.010006f
C203 B.n161 VSUBS 0.010006f
C204 B.n162 VSUBS 0.010006f
C205 B.n163 VSUBS 0.010006f
C206 B.n164 VSUBS 0.010006f
C207 B.n165 VSUBS 0.010006f
C208 B.n166 VSUBS 0.010006f
C209 B.n167 VSUBS 0.010006f
C210 B.n168 VSUBS 0.010006f
C211 B.n169 VSUBS 0.010006f
C212 B.n170 VSUBS 0.010006f
C213 B.n171 VSUBS 0.010006f
C214 B.n172 VSUBS 0.010006f
C215 B.n173 VSUBS 0.010006f
C216 B.n174 VSUBS 0.010006f
C217 B.n175 VSUBS 0.010006f
C218 B.n176 VSUBS 0.010006f
C219 B.n177 VSUBS 0.010006f
C220 B.n178 VSUBS 0.010006f
C221 B.n179 VSUBS 0.02308f
C222 B.n180 VSUBS 0.02308f
C223 B.n181 VSUBS 0.024887f
C224 B.n182 VSUBS 0.010006f
C225 B.n183 VSUBS 0.010006f
C226 B.n184 VSUBS 0.010006f
C227 B.n185 VSUBS 0.010006f
C228 B.n186 VSUBS 0.010006f
C229 B.n187 VSUBS 0.010006f
C230 B.n188 VSUBS 0.010006f
C231 B.n189 VSUBS 0.010006f
C232 B.n190 VSUBS 0.010006f
C233 B.n191 VSUBS 0.010006f
C234 B.n192 VSUBS 0.010006f
C235 B.n193 VSUBS 0.010006f
C236 B.n194 VSUBS 0.010006f
C237 B.n195 VSUBS 0.009123f
C238 B.n196 VSUBS 0.023182f
C239 B.n197 VSUBS 0.005886f
C240 B.n198 VSUBS 0.010006f
C241 B.n199 VSUBS 0.010006f
C242 B.n200 VSUBS 0.010006f
C243 B.n201 VSUBS 0.010006f
C244 B.n202 VSUBS 0.010006f
C245 B.n203 VSUBS 0.010006f
C246 B.n204 VSUBS 0.010006f
C247 B.n205 VSUBS 0.010006f
C248 B.n206 VSUBS 0.010006f
C249 B.n207 VSUBS 0.010006f
C250 B.n208 VSUBS 0.010006f
C251 B.n209 VSUBS 0.010006f
C252 B.n210 VSUBS 0.005886f
C253 B.n211 VSUBS 0.010006f
C254 B.n212 VSUBS 0.010006f
C255 B.n213 VSUBS 0.009123f
C256 B.n214 VSUBS 0.010006f
C257 B.n215 VSUBS 0.010006f
C258 B.n216 VSUBS 0.010006f
C259 B.n217 VSUBS 0.010006f
C260 B.n218 VSUBS 0.010006f
C261 B.n219 VSUBS 0.010006f
C262 B.n220 VSUBS 0.010006f
C263 B.n221 VSUBS 0.010006f
C264 B.n222 VSUBS 0.010006f
C265 B.n223 VSUBS 0.010006f
C266 B.n224 VSUBS 0.010006f
C267 B.n225 VSUBS 0.010006f
C268 B.n226 VSUBS 0.024887f
C269 B.n227 VSUBS 0.02308f
C270 B.n228 VSUBS 0.02308f
C271 B.n229 VSUBS 0.010006f
C272 B.n230 VSUBS 0.010006f
C273 B.n231 VSUBS 0.010006f
C274 B.n232 VSUBS 0.010006f
C275 B.n233 VSUBS 0.010006f
C276 B.n234 VSUBS 0.010006f
C277 B.n235 VSUBS 0.010006f
C278 B.n236 VSUBS 0.010006f
C279 B.n237 VSUBS 0.010006f
C280 B.n238 VSUBS 0.010006f
C281 B.n239 VSUBS 0.010006f
C282 B.n240 VSUBS 0.010006f
C283 B.n241 VSUBS 0.010006f
C284 B.n242 VSUBS 0.010006f
C285 B.n243 VSUBS 0.010006f
C286 B.n244 VSUBS 0.010006f
C287 B.n245 VSUBS 0.010006f
C288 B.n246 VSUBS 0.010006f
C289 B.n247 VSUBS 0.013057f
C290 B.n248 VSUBS 0.013909f
C291 B.n249 VSUBS 0.027659f
C292 VP.t0 VSUBS 0.330667f
C293 VP.t1 VSUBS 0.209764f
C294 VP.n0 VSUBS 2.04248f
.ends

