* NGSPICE file created from diff_pair_sample_0925.ext - technology: sky130A

.subckt diff_pair_sample_0925 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VP.t0 VDD1.t7 w_n2270_n1128# sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.97
X1 B.t11 B.t9 B.t10 w_n2270_n1128# sky130_fd_pr__pfet_01v8 ad=0.312 pd=2.38 as=0 ps=0 w=0.8 l=0.97
X2 B.t8 B.t6 B.t7 w_n2270_n1128# sky130_fd_pr__pfet_01v8 ad=0.312 pd=2.38 as=0 ps=0 w=0.8 l=0.97
X3 VDD2.t7 VN.t0 VTAIL.t3 w_n2270_n1128# sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.312 ps=2.38 w=0.8 l=0.97
X4 VDD2.t6 VN.t1 VTAIL.t7 w_n2270_n1128# sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.97
X5 VTAIL.t14 VP.t1 VDD1.t6 w_n2270_n1128# sky130_fd_pr__pfet_01v8 ad=0.312 pd=2.38 as=0.132 ps=1.13 w=0.8 l=0.97
X6 B.t5 B.t3 B.t4 w_n2270_n1128# sky130_fd_pr__pfet_01v8 ad=0.312 pd=2.38 as=0 ps=0 w=0.8 l=0.97
X7 B.t2 B.t0 B.t1 w_n2270_n1128# sky130_fd_pr__pfet_01v8 ad=0.312 pd=2.38 as=0 ps=0 w=0.8 l=0.97
X8 VDD2.t5 VN.t2 VTAIL.t4 w_n2270_n1128# sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.312 ps=2.38 w=0.8 l=0.97
X9 VDD2.t4 VN.t3 VTAIL.t5 w_n2270_n1128# sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.97
X10 VTAIL.t6 VN.t4 VDD2.t3 w_n2270_n1128# sky130_fd_pr__pfet_01v8 ad=0.312 pd=2.38 as=0.132 ps=1.13 w=0.8 l=0.97
X11 VDD1.t4 VP.t2 VTAIL.t13 w_n2270_n1128# sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.97
X12 VTAIL.t2 VN.t5 VDD2.t2 w_n2270_n1128# sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.97
X13 VTAIL.t0 VN.t6 VDD2.t1 w_n2270_n1128# sky130_fd_pr__pfet_01v8 ad=0.312 pd=2.38 as=0.132 ps=1.13 w=0.8 l=0.97
X14 VDD1.t5 VP.t3 VTAIL.t12 w_n2270_n1128# sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.312 ps=2.38 w=0.8 l=0.97
X15 VTAIL.t11 VP.t4 VDD1.t1 w_n2270_n1128# sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.97
X16 VTAIL.t10 VP.t5 VDD1.t3 w_n2270_n1128# sky130_fd_pr__pfet_01v8 ad=0.312 pd=2.38 as=0.132 ps=1.13 w=0.8 l=0.97
X17 VTAIL.t1 VN.t7 VDD2.t0 w_n2270_n1128# sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.97
X18 VDD1.t2 VP.t6 VTAIL.t9 w_n2270_n1128# sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.312 ps=2.38 w=0.8 l=0.97
X19 VDD1.t0 VP.t7 VTAIL.t8 w_n2270_n1128# sky130_fd_pr__pfet_01v8 ad=0.132 pd=1.13 as=0.132 ps=1.13 w=0.8 l=0.97
R0 VP.n8 VP.n7 161.3
R1 VP.n9 VP.n4 161.3
R2 VP.n11 VP.n10 161.3
R3 VP.n13 VP.n3 161.3
R4 VP.n26 VP.n0 161.3
R5 VP.n24 VP.n23 161.3
R6 VP.n22 VP.n1 161.3
R7 VP.n21 VP.n20 161.3
R8 VP.n18 VP.n2 161.3
R9 VP.n15 VP.n14 80.6037
R10 VP.n28 VP.n27 80.6037
R11 VP.n17 VP.n16 80.6037
R12 VP.n5 VP.t5 75.3094
R13 VP.n17 VP.t1 60.3747
R14 VP.n27 VP.t3 60.3747
R15 VP.n14 VP.t6 60.3747
R16 VP.n18 VP.n17 54.8403
R17 VP.n27 VP.n26 54.8403
R18 VP.n14 VP.n13 54.8403
R19 VP.n6 VP.n5 46.9959
R20 VP.n8 VP.n5 44.1162
R21 VP.n20 VP.n1 40.577
R22 VP.n24 VP.n1 40.577
R23 VP.n11 VP.n4 40.577
R24 VP.n7 VP.n4 40.577
R25 VP.n16 VP.n15 34.9559
R26 VP.n19 VP.t7 19.8768
R27 VP.n25 VP.t0 19.8768
R28 VP.n12 VP.t4 19.8768
R29 VP.n6 VP.t2 19.8768
R30 VP.n19 VP.n18 17.2148
R31 VP.n26 VP.n25 17.2148
R32 VP.n13 VP.n12 17.2148
R33 VP.n20 VP.n19 7.37805
R34 VP.n25 VP.n24 7.37805
R35 VP.n12 VP.n11 7.37805
R36 VP.n7 VP.n6 7.37805
R37 VP.n15 VP.n3 0.285035
R38 VP.n16 VP.n2 0.285035
R39 VP.n28 VP.n0 0.285035
R40 VP.n9 VP.n8 0.189894
R41 VP.n10 VP.n9 0.189894
R42 VP.n10 VP.n3 0.189894
R43 VP.n21 VP.n2 0.189894
R44 VP.n22 VP.n21 0.189894
R45 VP.n23 VP.n22 0.189894
R46 VP.n23 VP.n0 0.189894
R47 VP VP.n28 0.146778
R48 VDD1 VDD1.n0 638.361
R49 VDD1.n3 VDD1.n2 638.247
R50 VDD1.n3 VDD1.n1 638.247
R51 VDD1.n5 VDD1.n4 637.742
R52 VDD1.n4 VDD1.t1 40.6317
R53 VDD1.n4 VDD1.t2 40.6317
R54 VDD1.n0 VDD1.t3 40.6317
R55 VDD1.n0 VDD1.t4 40.6317
R56 VDD1.n2 VDD1.t7 40.6317
R57 VDD1.n2 VDD1.t5 40.6317
R58 VDD1.n1 VDD1.t6 40.6317
R59 VDD1.n1 VDD1.t0 40.6317
R60 VDD1.n5 VDD1.n3 30.0311
R61 VDD1 VDD1.n5 0.502655
R62 VTAIL.n15 VTAIL.t3 661.696
R63 VTAIL.n2 VTAIL.t6 661.696
R64 VTAIL.n3 VTAIL.t12 661.696
R65 VTAIL.n6 VTAIL.t14 661.696
R66 VTAIL.n14 VTAIL.t9 661.696
R67 VTAIL.n11 VTAIL.t10 661.696
R68 VTAIL.n10 VTAIL.t4 661.696
R69 VTAIL.n7 VTAIL.t0 661.696
R70 VTAIL.n1 VTAIL.n0 621.064
R71 VTAIL.n5 VTAIL.n4 621.064
R72 VTAIL.n13 VTAIL.n12 621.064
R73 VTAIL.n9 VTAIL.n8 621.064
R74 VTAIL.n0 VTAIL.t7 40.6317
R75 VTAIL.n0 VTAIL.t1 40.6317
R76 VTAIL.n4 VTAIL.t8 40.6317
R77 VTAIL.n4 VTAIL.t15 40.6317
R78 VTAIL.n12 VTAIL.t13 40.6317
R79 VTAIL.n12 VTAIL.t11 40.6317
R80 VTAIL.n8 VTAIL.t5 40.6317
R81 VTAIL.n8 VTAIL.t2 40.6317
R82 VTAIL.n15 VTAIL.n14 14.1772
R83 VTAIL.n7 VTAIL.n6 14.1772
R84 VTAIL.n9 VTAIL.n7 1.12119
R85 VTAIL.n10 VTAIL.n9 1.12119
R86 VTAIL.n13 VTAIL.n11 1.12119
R87 VTAIL.n14 VTAIL.n13 1.12119
R88 VTAIL.n6 VTAIL.n5 1.12119
R89 VTAIL.n5 VTAIL.n3 1.12119
R90 VTAIL.n2 VTAIL.n1 1.12119
R91 VTAIL VTAIL.n15 1.063
R92 VTAIL.n11 VTAIL.n10 0.470328
R93 VTAIL.n3 VTAIL.n2 0.470328
R94 VTAIL VTAIL.n1 0.0586897
R95 B.n66 B.t11 676.056
R96 B.n72 B.t5 676.056
R97 B.n20 B.t7 676.056
R98 B.n28 B.t1 676.056
R99 B.n67 B.t10 650.843
R100 B.n73 B.t4 650.843
R101 B.n21 B.t8 650.843
R102 B.n29 B.t2 650.843
R103 B.n256 B.n33 585
R104 B.n258 B.n257 585
R105 B.n259 B.n32 585
R106 B.n261 B.n260 585
R107 B.n262 B.n31 585
R108 B.n264 B.n263 585
R109 B.n265 B.n30 585
R110 B.n267 B.n266 585
R111 B.n268 B.n27 585
R112 B.n271 B.n270 585
R113 B.n272 B.n26 585
R114 B.n274 B.n273 585
R115 B.n275 B.n25 585
R116 B.n277 B.n276 585
R117 B.n278 B.n24 585
R118 B.n280 B.n279 585
R119 B.n281 B.n23 585
R120 B.n283 B.n282 585
R121 B.n285 B.n284 585
R122 B.n286 B.n19 585
R123 B.n288 B.n287 585
R124 B.n289 B.n18 585
R125 B.n291 B.n290 585
R126 B.n292 B.n17 585
R127 B.n294 B.n293 585
R128 B.n295 B.n16 585
R129 B.n297 B.n296 585
R130 B.n255 B.n254 585
R131 B.n253 B.n34 585
R132 B.n252 B.n251 585
R133 B.n250 B.n35 585
R134 B.n249 B.n248 585
R135 B.n247 B.n36 585
R136 B.n246 B.n245 585
R137 B.n244 B.n37 585
R138 B.n243 B.n242 585
R139 B.n241 B.n38 585
R140 B.n240 B.n239 585
R141 B.n238 B.n39 585
R142 B.n237 B.n236 585
R143 B.n235 B.n40 585
R144 B.n234 B.n233 585
R145 B.n232 B.n41 585
R146 B.n231 B.n230 585
R147 B.n229 B.n42 585
R148 B.n228 B.n227 585
R149 B.n226 B.n43 585
R150 B.n225 B.n224 585
R151 B.n223 B.n44 585
R152 B.n222 B.n221 585
R153 B.n220 B.n45 585
R154 B.n219 B.n218 585
R155 B.n217 B.n46 585
R156 B.n216 B.n215 585
R157 B.n214 B.n47 585
R158 B.n213 B.n212 585
R159 B.n211 B.n48 585
R160 B.n210 B.n209 585
R161 B.n208 B.n49 585
R162 B.n207 B.n206 585
R163 B.n205 B.n50 585
R164 B.n204 B.n203 585
R165 B.n202 B.n51 585
R166 B.n201 B.n200 585
R167 B.n199 B.n52 585
R168 B.n198 B.n197 585
R169 B.n196 B.n53 585
R170 B.n195 B.n194 585
R171 B.n193 B.n54 585
R172 B.n192 B.n191 585
R173 B.n190 B.n55 585
R174 B.n189 B.n188 585
R175 B.n187 B.n56 585
R176 B.n186 B.n185 585
R177 B.n184 B.n57 585
R178 B.n183 B.n182 585
R179 B.n181 B.n58 585
R180 B.n180 B.n179 585
R181 B.n178 B.n59 585
R182 B.n177 B.n176 585
R183 B.n175 B.n60 585
R184 B.n174 B.n173 585
R185 B.n132 B.n131 585
R186 B.n133 B.n78 585
R187 B.n135 B.n134 585
R188 B.n136 B.n77 585
R189 B.n138 B.n137 585
R190 B.n139 B.n76 585
R191 B.n141 B.n140 585
R192 B.n142 B.n75 585
R193 B.n144 B.n143 585
R194 B.n146 B.n145 585
R195 B.n147 B.n71 585
R196 B.n149 B.n148 585
R197 B.n150 B.n70 585
R198 B.n152 B.n151 585
R199 B.n153 B.n69 585
R200 B.n155 B.n154 585
R201 B.n156 B.n68 585
R202 B.n158 B.n157 585
R203 B.n160 B.n65 585
R204 B.n162 B.n161 585
R205 B.n163 B.n64 585
R206 B.n165 B.n164 585
R207 B.n166 B.n63 585
R208 B.n168 B.n167 585
R209 B.n169 B.n62 585
R210 B.n171 B.n170 585
R211 B.n172 B.n61 585
R212 B.n130 B.n79 585
R213 B.n129 B.n128 585
R214 B.n127 B.n80 585
R215 B.n126 B.n125 585
R216 B.n124 B.n81 585
R217 B.n123 B.n122 585
R218 B.n121 B.n82 585
R219 B.n120 B.n119 585
R220 B.n118 B.n83 585
R221 B.n117 B.n116 585
R222 B.n115 B.n84 585
R223 B.n114 B.n113 585
R224 B.n112 B.n85 585
R225 B.n111 B.n110 585
R226 B.n109 B.n86 585
R227 B.n108 B.n107 585
R228 B.n106 B.n87 585
R229 B.n105 B.n104 585
R230 B.n103 B.n88 585
R231 B.n102 B.n101 585
R232 B.n100 B.n89 585
R233 B.n99 B.n98 585
R234 B.n97 B.n90 585
R235 B.n96 B.n95 585
R236 B.n94 B.n91 585
R237 B.n93 B.n92 585
R238 B.n2 B.n0 585
R239 B.n337 B.n1 585
R240 B.n336 B.n335 585
R241 B.n334 B.n3 585
R242 B.n333 B.n332 585
R243 B.n331 B.n4 585
R244 B.n330 B.n329 585
R245 B.n328 B.n5 585
R246 B.n327 B.n326 585
R247 B.n325 B.n6 585
R248 B.n324 B.n323 585
R249 B.n322 B.n7 585
R250 B.n321 B.n320 585
R251 B.n319 B.n8 585
R252 B.n318 B.n317 585
R253 B.n316 B.n9 585
R254 B.n315 B.n314 585
R255 B.n313 B.n10 585
R256 B.n312 B.n311 585
R257 B.n310 B.n11 585
R258 B.n309 B.n308 585
R259 B.n307 B.n12 585
R260 B.n306 B.n305 585
R261 B.n304 B.n13 585
R262 B.n303 B.n302 585
R263 B.n301 B.n14 585
R264 B.n300 B.n299 585
R265 B.n298 B.n15 585
R266 B.n339 B.n338 585
R267 B.n132 B.n79 530.939
R268 B.n296 B.n15 530.939
R269 B.n174 B.n61 530.939
R270 B.n254 B.n33 530.939
R271 B.n66 B.t9 222.595
R272 B.n72 B.t3 222.595
R273 B.n20 B.t6 222.595
R274 B.n28 B.t0 222.595
R275 B.n128 B.n79 163.367
R276 B.n128 B.n127 163.367
R277 B.n127 B.n126 163.367
R278 B.n126 B.n81 163.367
R279 B.n122 B.n81 163.367
R280 B.n122 B.n121 163.367
R281 B.n121 B.n120 163.367
R282 B.n120 B.n83 163.367
R283 B.n116 B.n83 163.367
R284 B.n116 B.n115 163.367
R285 B.n115 B.n114 163.367
R286 B.n114 B.n85 163.367
R287 B.n110 B.n85 163.367
R288 B.n110 B.n109 163.367
R289 B.n109 B.n108 163.367
R290 B.n108 B.n87 163.367
R291 B.n104 B.n87 163.367
R292 B.n104 B.n103 163.367
R293 B.n103 B.n102 163.367
R294 B.n102 B.n89 163.367
R295 B.n98 B.n89 163.367
R296 B.n98 B.n97 163.367
R297 B.n97 B.n96 163.367
R298 B.n96 B.n91 163.367
R299 B.n92 B.n91 163.367
R300 B.n92 B.n2 163.367
R301 B.n338 B.n2 163.367
R302 B.n338 B.n337 163.367
R303 B.n337 B.n336 163.367
R304 B.n336 B.n3 163.367
R305 B.n332 B.n3 163.367
R306 B.n332 B.n331 163.367
R307 B.n331 B.n330 163.367
R308 B.n330 B.n5 163.367
R309 B.n326 B.n5 163.367
R310 B.n326 B.n325 163.367
R311 B.n325 B.n324 163.367
R312 B.n324 B.n7 163.367
R313 B.n320 B.n7 163.367
R314 B.n320 B.n319 163.367
R315 B.n319 B.n318 163.367
R316 B.n318 B.n9 163.367
R317 B.n314 B.n9 163.367
R318 B.n314 B.n313 163.367
R319 B.n313 B.n312 163.367
R320 B.n312 B.n11 163.367
R321 B.n308 B.n11 163.367
R322 B.n308 B.n307 163.367
R323 B.n307 B.n306 163.367
R324 B.n306 B.n13 163.367
R325 B.n302 B.n13 163.367
R326 B.n302 B.n301 163.367
R327 B.n301 B.n300 163.367
R328 B.n300 B.n15 163.367
R329 B.n133 B.n132 163.367
R330 B.n134 B.n133 163.367
R331 B.n134 B.n77 163.367
R332 B.n138 B.n77 163.367
R333 B.n139 B.n138 163.367
R334 B.n140 B.n139 163.367
R335 B.n140 B.n75 163.367
R336 B.n144 B.n75 163.367
R337 B.n145 B.n144 163.367
R338 B.n145 B.n71 163.367
R339 B.n149 B.n71 163.367
R340 B.n150 B.n149 163.367
R341 B.n151 B.n150 163.367
R342 B.n151 B.n69 163.367
R343 B.n155 B.n69 163.367
R344 B.n156 B.n155 163.367
R345 B.n157 B.n156 163.367
R346 B.n157 B.n65 163.367
R347 B.n162 B.n65 163.367
R348 B.n163 B.n162 163.367
R349 B.n164 B.n163 163.367
R350 B.n164 B.n63 163.367
R351 B.n168 B.n63 163.367
R352 B.n169 B.n168 163.367
R353 B.n170 B.n169 163.367
R354 B.n170 B.n61 163.367
R355 B.n175 B.n174 163.367
R356 B.n176 B.n175 163.367
R357 B.n176 B.n59 163.367
R358 B.n180 B.n59 163.367
R359 B.n181 B.n180 163.367
R360 B.n182 B.n181 163.367
R361 B.n182 B.n57 163.367
R362 B.n186 B.n57 163.367
R363 B.n187 B.n186 163.367
R364 B.n188 B.n187 163.367
R365 B.n188 B.n55 163.367
R366 B.n192 B.n55 163.367
R367 B.n193 B.n192 163.367
R368 B.n194 B.n193 163.367
R369 B.n194 B.n53 163.367
R370 B.n198 B.n53 163.367
R371 B.n199 B.n198 163.367
R372 B.n200 B.n199 163.367
R373 B.n200 B.n51 163.367
R374 B.n204 B.n51 163.367
R375 B.n205 B.n204 163.367
R376 B.n206 B.n205 163.367
R377 B.n206 B.n49 163.367
R378 B.n210 B.n49 163.367
R379 B.n211 B.n210 163.367
R380 B.n212 B.n211 163.367
R381 B.n212 B.n47 163.367
R382 B.n216 B.n47 163.367
R383 B.n217 B.n216 163.367
R384 B.n218 B.n217 163.367
R385 B.n218 B.n45 163.367
R386 B.n222 B.n45 163.367
R387 B.n223 B.n222 163.367
R388 B.n224 B.n223 163.367
R389 B.n224 B.n43 163.367
R390 B.n228 B.n43 163.367
R391 B.n229 B.n228 163.367
R392 B.n230 B.n229 163.367
R393 B.n230 B.n41 163.367
R394 B.n234 B.n41 163.367
R395 B.n235 B.n234 163.367
R396 B.n236 B.n235 163.367
R397 B.n236 B.n39 163.367
R398 B.n240 B.n39 163.367
R399 B.n241 B.n240 163.367
R400 B.n242 B.n241 163.367
R401 B.n242 B.n37 163.367
R402 B.n246 B.n37 163.367
R403 B.n247 B.n246 163.367
R404 B.n248 B.n247 163.367
R405 B.n248 B.n35 163.367
R406 B.n252 B.n35 163.367
R407 B.n253 B.n252 163.367
R408 B.n254 B.n253 163.367
R409 B.n296 B.n295 163.367
R410 B.n295 B.n294 163.367
R411 B.n294 B.n17 163.367
R412 B.n290 B.n17 163.367
R413 B.n290 B.n289 163.367
R414 B.n289 B.n288 163.367
R415 B.n288 B.n19 163.367
R416 B.n284 B.n19 163.367
R417 B.n284 B.n283 163.367
R418 B.n283 B.n23 163.367
R419 B.n279 B.n23 163.367
R420 B.n279 B.n278 163.367
R421 B.n278 B.n277 163.367
R422 B.n277 B.n25 163.367
R423 B.n273 B.n25 163.367
R424 B.n273 B.n272 163.367
R425 B.n272 B.n271 163.367
R426 B.n271 B.n27 163.367
R427 B.n266 B.n27 163.367
R428 B.n266 B.n265 163.367
R429 B.n265 B.n264 163.367
R430 B.n264 B.n31 163.367
R431 B.n260 B.n31 163.367
R432 B.n260 B.n259 163.367
R433 B.n259 B.n258 163.367
R434 B.n258 B.n33 163.367
R435 B.n159 B.n67 59.5399
R436 B.n74 B.n73 59.5399
R437 B.n22 B.n21 59.5399
R438 B.n269 B.n29 59.5399
R439 B.n298 B.n297 34.4981
R440 B.n256 B.n255 34.4981
R441 B.n173 B.n172 34.4981
R442 B.n131 B.n130 34.4981
R443 B.n67 B.n66 25.2126
R444 B.n73 B.n72 25.2126
R445 B.n21 B.n20 25.2126
R446 B.n29 B.n28 25.2126
R447 B B.n339 18.0485
R448 B.n297 B.n16 10.6151
R449 B.n293 B.n16 10.6151
R450 B.n293 B.n292 10.6151
R451 B.n292 B.n291 10.6151
R452 B.n291 B.n18 10.6151
R453 B.n287 B.n18 10.6151
R454 B.n287 B.n286 10.6151
R455 B.n286 B.n285 10.6151
R456 B.n282 B.n281 10.6151
R457 B.n281 B.n280 10.6151
R458 B.n280 B.n24 10.6151
R459 B.n276 B.n24 10.6151
R460 B.n276 B.n275 10.6151
R461 B.n275 B.n274 10.6151
R462 B.n274 B.n26 10.6151
R463 B.n270 B.n26 10.6151
R464 B.n268 B.n267 10.6151
R465 B.n267 B.n30 10.6151
R466 B.n263 B.n30 10.6151
R467 B.n263 B.n262 10.6151
R468 B.n262 B.n261 10.6151
R469 B.n261 B.n32 10.6151
R470 B.n257 B.n32 10.6151
R471 B.n257 B.n256 10.6151
R472 B.n173 B.n60 10.6151
R473 B.n177 B.n60 10.6151
R474 B.n178 B.n177 10.6151
R475 B.n179 B.n178 10.6151
R476 B.n179 B.n58 10.6151
R477 B.n183 B.n58 10.6151
R478 B.n184 B.n183 10.6151
R479 B.n185 B.n184 10.6151
R480 B.n185 B.n56 10.6151
R481 B.n189 B.n56 10.6151
R482 B.n190 B.n189 10.6151
R483 B.n191 B.n190 10.6151
R484 B.n191 B.n54 10.6151
R485 B.n195 B.n54 10.6151
R486 B.n196 B.n195 10.6151
R487 B.n197 B.n196 10.6151
R488 B.n197 B.n52 10.6151
R489 B.n201 B.n52 10.6151
R490 B.n202 B.n201 10.6151
R491 B.n203 B.n202 10.6151
R492 B.n203 B.n50 10.6151
R493 B.n207 B.n50 10.6151
R494 B.n208 B.n207 10.6151
R495 B.n209 B.n208 10.6151
R496 B.n209 B.n48 10.6151
R497 B.n213 B.n48 10.6151
R498 B.n214 B.n213 10.6151
R499 B.n215 B.n214 10.6151
R500 B.n215 B.n46 10.6151
R501 B.n219 B.n46 10.6151
R502 B.n220 B.n219 10.6151
R503 B.n221 B.n220 10.6151
R504 B.n221 B.n44 10.6151
R505 B.n225 B.n44 10.6151
R506 B.n226 B.n225 10.6151
R507 B.n227 B.n226 10.6151
R508 B.n227 B.n42 10.6151
R509 B.n231 B.n42 10.6151
R510 B.n232 B.n231 10.6151
R511 B.n233 B.n232 10.6151
R512 B.n233 B.n40 10.6151
R513 B.n237 B.n40 10.6151
R514 B.n238 B.n237 10.6151
R515 B.n239 B.n238 10.6151
R516 B.n239 B.n38 10.6151
R517 B.n243 B.n38 10.6151
R518 B.n244 B.n243 10.6151
R519 B.n245 B.n244 10.6151
R520 B.n245 B.n36 10.6151
R521 B.n249 B.n36 10.6151
R522 B.n250 B.n249 10.6151
R523 B.n251 B.n250 10.6151
R524 B.n251 B.n34 10.6151
R525 B.n255 B.n34 10.6151
R526 B.n131 B.n78 10.6151
R527 B.n135 B.n78 10.6151
R528 B.n136 B.n135 10.6151
R529 B.n137 B.n136 10.6151
R530 B.n137 B.n76 10.6151
R531 B.n141 B.n76 10.6151
R532 B.n142 B.n141 10.6151
R533 B.n143 B.n142 10.6151
R534 B.n147 B.n146 10.6151
R535 B.n148 B.n147 10.6151
R536 B.n148 B.n70 10.6151
R537 B.n152 B.n70 10.6151
R538 B.n153 B.n152 10.6151
R539 B.n154 B.n153 10.6151
R540 B.n154 B.n68 10.6151
R541 B.n158 B.n68 10.6151
R542 B.n161 B.n160 10.6151
R543 B.n161 B.n64 10.6151
R544 B.n165 B.n64 10.6151
R545 B.n166 B.n165 10.6151
R546 B.n167 B.n166 10.6151
R547 B.n167 B.n62 10.6151
R548 B.n171 B.n62 10.6151
R549 B.n172 B.n171 10.6151
R550 B.n130 B.n129 10.6151
R551 B.n129 B.n80 10.6151
R552 B.n125 B.n80 10.6151
R553 B.n125 B.n124 10.6151
R554 B.n124 B.n123 10.6151
R555 B.n123 B.n82 10.6151
R556 B.n119 B.n82 10.6151
R557 B.n119 B.n118 10.6151
R558 B.n118 B.n117 10.6151
R559 B.n117 B.n84 10.6151
R560 B.n113 B.n84 10.6151
R561 B.n113 B.n112 10.6151
R562 B.n112 B.n111 10.6151
R563 B.n111 B.n86 10.6151
R564 B.n107 B.n86 10.6151
R565 B.n107 B.n106 10.6151
R566 B.n106 B.n105 10.6151
R567 B.n105 B.n88 10.6151
R568 B.n101 B.n88 10.6151
R569 B.n101 B.n100 10.6151
R570 B.n100 B.n99 10.6151
R571 B.n99 B.n90 10.6151
R572 B.n95 B.n90 10.6151
R573 B.n95 B.n94 10.6151
R574 B.n94 B.n93 10.6151
R575 B.n93 B.n0 10.6151
R576 B.n335 B.n1 10.6151
R577 B.n335 B.n334 10.6151
R578 B.n334 B.n333 10.6151
R579 B.n333 B.n4 10.6151
R580 B.n329 B.n4 10.6151
R581 B.n329 B.n328 10.6151
R582 B.n328 B.n327 10.6151
R583 B.n327 B.n6 10.6151
R584 B.n323 B.n6 10.6151
R585 B.n323 B.n322 10.6151
R586 B.n322 B.n321 10.6151
R587 B.n321 B.n8 10.6151
R588 B.n317 B.n8 10.6151
R589 B.n317 B.n316 10.6151
R590 B.n316 B.n315 10.6151
R591 B.n315 B.n10 10.6151
R592 B.n311 B.n10 10.6151
R593 B.n311 B.n310 10.6151
R594 B.n310 B.n309 10.6151
R595 B.n309 B.n12 10.6151
R596 B.n305 B.n12 10.6151
R597 B.n305 B.n304 10.6151
R598 B.n304 B.n303 10.6151
R599 B.n303 B.n14 10.6151
R600 B.n299 B.n14 10.6151
R601 B.n299 B.n298 10.6151
R602 B.n282 B.n22 6.5566
R603 B.n270 B.n269 6.5566
R604 B.n146 B.n74 6.5566
R605 B.n159 B.n158 6.5566
R606 B.n285 B.n22 4.05904
R607 B.n269 B.n268 4.05904
R608 B.n143 B.n74 4.05904
R609 B.n160 B.n159 4.05904
R610 B.n339 B.n0 2.81026
R611 B.n339 B.n1 2.81026
R612 VN.n23 VN.n13 161.3
R613 VN.n21 VN.n20 161.3
R614 VN.n19 VN.n14 161.3
R615 VN.n18 VN.n17 161.3
R616 VN.n10 VN.n0 161.3
R617 VN.n8 VN.n7 161.3
R618 VN.n6 VN.n1 161.3
R619 VN.n5 VN.n4 161.3
R620 VN.n25 VN.n24 80.6037
R621 VN.n12 VN.n11 80.6037
R622 VN.n2 VN.t4 75.3094
R623 VN.n15 VN.t2 75.3094
R624 VN.n11 VN.t0 60.3747
R625 VN.n24 VN.t6 60.3747
R626 VN.n11 VN.n10 54.8403
R627 VN.n24 VN.n23 54.8403
R628 VN.n3 VN.n2 46.9959
R629 VN.n16 VN.n15 46.9959
R630 VN.n18 VN.n15 44.1163
R631 VN.n5 VN.n2 44.1163
R632 VN.n4 VN.n1 40.577
R633 VN.n8 VN.n1 40.577
R634 VN.n17 VN.n14 40.577
R635 VN.n21 VN.n14 40.577
R636 VN VN.n25 35.2415
R637 VN.n3 VN.t1 19.8768
R638 VN.n9 VN.t7 19.8768
R639 VN.n16 VN.t5 19.8768
R640 VN.n22 VN.t3 19.8768
R641 VN.n10 VN.n9 17.2148
R642 VN.n23 VN.n22 17.2148
R643 VN.n4 VN.n3 7.37805
R644 VN.n9 VN.n8 7.37805
R645 VN.n17 VN.n16 7.37805
R646 VN.n22 VN.n21 7.37805
R647 VN.n25 VN.n13 0.285035
R648 VN.n12 VN.n0 0.285035
R649 VN.n20 VN.n13 0.189894
R650 VN.n20 VN.n19 0.189894
R651 VN.n19 VN.n18 0.189894
R652 VN.n6 VN.n5 0.189894
R653 VN.n7 VN.n6 0.189894
R654 VN.n7 VN.n0 0.189894
R655 VN VN.n12 0.146778
R656 VDD2.n2 VDD2.n1 638.247
R657 VDD2.n2 VDD2.n0 638.247
R658 VDD2 VDD2.n5 638.245
R659 VDD2.n4 VDD2.n3 637.742
R660 VDD2.n5 VDD2.t2 40.6317
R661 VDD2.n5 VDD2.t5 40.6317
R662 VDD2.n3 VDD2.t1 40.6317
R663 VDD2.n3 VDD2.t4 40.6317
R664 VDD2.n1 VDD2.t0 40.6317
R665 VDD2.n1 VDD2.t7 40.6317
R666 VDD2.n0 VDD2.t3 40.6317
R667 VDD2.n0 VDD2.t6 40.6317
R668 VDD2.n4 VDD2.n2 29.4481
R669 VDD2 VDD2.n4 0.619035
C0 VP VDD2 0.355513f
C1 VN w_n2270_n1128# 3.91256f
C2 VN B 0.687206f
C3 w_n2270_n1128# VTAIL 1.33401f
C4 B VTAIL 0.805563f
C5 w_n2270_n1128# VDD2 1.13905f
C6 VP w_n2270_n1128# 4.19397f
C7 B VDD2 0.894518f
C8 VP B 1.16309f
C9 VN VDD1 0.156626f
C10 w_n2270_n1128# B 4.48033f
C11 VDD1 VTAIL 2.86668f
C12 VDD1 VDD2 0.961196f
C13 VP VDD1 0.999578f
C14 VN VTAIL 1.32955f
C15 w_n2270_n1128# VDD1 1.09417f
C16 VN VDD2 0.802868f
C17 VDD1 B 0.849113f
C18 VN VP 3.60111f
C19 VDD2 VTAIL 2.91017f
C20 VP VTAIL 1.34365f
C21 VDD2 VSUBS 0.645323f
C22 VDD1 VSUBS 0.98942f
C23 VTAIL VSUBS 0.324232f
C24 VN VSUBS 4.10874f
C25 VP VSUBS 1.404184f
C26 B VSUBS 2.120428f
C27 w_n2270_n1128# VSUBS 33.096603f
C28 VDD2.t3 VSUBS 0.013824f
C29 VDD2.t6 VSUBS 0.013824f
C30 VDD2.n0 VSUBS 0.029913f
C31 VDD2.t0 VSUBS 0.013824f
C32 VDD2.t7 VSUBS 0.013824f
C33 VDD2.n1 VSUBS 0.029913f
C34 VDD2.n2 VSUBS 1.22718f
C35 VDD2.t1 VSUBS 0.013824f
C36 VDD2.t4 VSUBS 0.013824f
C37 VDD2.n3 VSUBS 0.029767f
C38 VDD2.n4 VSUBS 1.18053f
C39 VDD2.t2 VSUBS 0.013824f
C40 VDD2.t5 VSUBS 0.013824f
C41 VDD2.n5 VSUBS 0.029911f
C42 VN.n0 VSUBS 0.080095f
C43 VN.t7 VSUBS 0.076146f
C44 VN.n1 VSUBS 0.04848f
C45 VN.t4 VSUBS 0.20184f
C46 VN.n2 VSUBS 0.179309f
C47 VN.t1 VSUBS 0.076146f
C48 VN.n3 VSUBS 0.148198f
C49 VN.n4 VSUBS 0.080204f
C50 VN.n5 VSUBS 0.25256f
C51 VN.n6 VSUBS 0.060024f
C52 VN.n7 VSUBS 0.060024f
C53 VN.n8 VSUBS 0.080204f
C54 VN.n9 VSUBS 0.098463f
C55 VN.n10 VSUBS 0.078484f
C56 VN.t0 VSUBS 0.164801f
C57 VN.n11 VSUBS 0.186369f
C58 VN.n12 VSUBS 0.056215f
C59 VN.n13 VSUBS 0.080095f
C60 VN.t3 VSUBS 0.076146f
C61 VN.n14 VSUBS 0.04848f
C62 VN.t2 VSUBS 0.20184f
C63 VN.n15 VSUBS 0.179309f
C64 VN.t5 VSUBS 0.076146f
C65 VN.n16 VSUBS 0.148198f
C66 VN.n17 VSUBS 0.080204f
C67 VN.n18 VSUBS 0.25256f
C68 VN.n19 VSUBS 0.060024f
C69 VN.n20 VSUBS 0.060024f
C70 VN.n21 VSUBS 0.080204f
C71 VN.n22 VSUBS 0.098463f
C72 VN.n23 VSUBS 0.078484f
C73 VN.t6 VSUBS 0.164801f
C74 VN.n24 VSUBS 0.186369f
C75 VN.n25 VSUBS 1.84039f
C76 B.n0 VSUBS 0.006406f
C77 B.n1 VSUBS 0.006406f
C78 B.n2 VSUBS 0.01013f
C79 B.n3 VSUBS 0.01013f
C80 B.n4 VSUBS 0.01013f
C81 B.n5 VSUBS 0.01013f
C82 B.n6 VSUBS 0.01013f
C83 B.n7 VSUBS 0.01013f
C84 B.n8 VSUBS 0.01013f
C85 B.n9 VSUBS 0.01013f
C86 B.n10 VSUBS 0.01013f
C87 B.n11 VSUBS 0.01013f
C88 B.n12 VSUBS 0.01013f
C89 B.n13 VSUBS 0.01013f
C90 B.n14 VSUBS 0.01013f
C91 B.n15 VSUBS 0.023794f
C92 B.n16 VSUBS 0.01013f
C93 B.n17 VSUBS 0.01013f
C94 B.n18 VSUBS 0.01013f
C95 B.n19 VSUBS 0.01013f
C96 B.t8 VSUBS 0.022231f
C97 B.t7 VSUBS 0.023625f
C98 B.t6 VSUBS 0.058778f
C99 B.n20 VSUBS 0.057098f
C100 B.n21 VSUBS 0.051823f
C101 B.n22 VSUBS 0.023471f
C102 B.n23 VSUBS 0.01013f
C103 B.n24 VSUBS 0.01013f
C104 B.n25 VSUBS 0.01013f
C105 B.n26 VSUBS 0.01013f
C106 B.n27 VSUBS 0.01013f
C107 B.t2 VSUBS 0.022231f
C108 B.t1 VSUBS 0.023625f
C109 B.t0 VSUBS 0.058778f
C110 B.n28 VSUBS 0.057098f
C111 B.n29 VSUBS 0.051823f
C112 B.n30 VSUBS 0.01013f
C113 B.n31 VSUBS 0.01013f
C114 B.n32 VSUBS 0.01013f
C115 B.n33 VSUBS 0.025369f
C116 B.n34 VSUBS 0.01013f
C117 B.n35 VSUBS 0.01013f
C118 B.n36 VSUBS 0.01013f
C119 B.n37 VSUBS 0.01013f
C120 B.n38 VSUBS 0.01013f
C121 B.n39 VSUBS 0.01013f
C122 B.n40 VSUBS 0.01013f
C123 B.n41 VSUBS 0.01013f
C124 B.n42 VSUBS 0.01013f
C125 B.n43 VSUBS 0.01013f
C126 B.n44 VSUBS 0.01013f
C127 B.n45 VSUBS 0.01013f
C128 B.n46 VSUBS 0.01013f
C129 B.n47 VSUBS 0.01013f
C130 B.n48 VSUBS 0.01013f
C131 B.n49 VSUBS 0.01013f
C132 B.n50 VSUBS 0.01013f
C133 B.n51 VSUBS 0.01013f
C134 B.n52 VSUBS 0.01013f
C135 B.n53 VSUBS 0.01013f
C136 B.n54 VSUBS 0.01013f
C137 B.n55 VSUBS 0.01013f
C138 B.n56 VSUBS 0.01013f
C139 B.n57 VSUBS 0.01013f
C140 B.n58 VSUBS 0.01013f
C141 B.n59 VSUBS 0.01013f
C142 B.n60 VSUBS 0.01013f
C143 B.n61 VSUBS 0.025369f
C144 B.n62 VSUBS 0.01013f
C145 B.n63 VSUBS 0.01013f
C146 B.n64 VSUBS 0.01013f
C147 B.n65 VSUBS 0.01013f
C148 B.t10 VSUBS 0.022231f
C149 B.t11 VSUBS 0.023625f
C150 B.t9 VSUBS 0.058778f
C151 B.n66 VSUBS 0.057098f
C152 B.n67 VSUBS 0.051823f
C153 B.n68 VSUBS 0.01013f
C154 B.n69 VSUBS 0.01013f
C155 B.n70 VSUBS 0.01013f
C156 B.n71 VSUBS 0.01013f
C157 B.t4 VSUBS 0.022231f
C158 B.t5 VSUBS 0.023625f
C159 B.t3 VSUBS 0.058778f
C160 B.n72 VSUBS 0.057098f
C161 B.n73 VSUBS 0.051823f
C162 B.n74 VSUBS 0.023471f
C163 B.n75 VSUBS 0.01013f
C164 B.n76 VSUBS 0.01013f
C165 B.n77 VSUBS 0.01013f
C166 B.n78 VSUBS 0.01013f
C167 B.n79 VSUBS 0.023794f
C168 B.n80 VSUBS 0.01013f
C169 B.n81 VSUBS 0.01013f
C170 B.n82 VSUBS 0.01013f
C171 B.n83 VSUBS 0.01013f
C172 B.n84 VSUBS 0.01013f
C173 B.n85 VSUBS 0.01013f
C174 B.n86 VSUBS 0.01013f
C175 B.n87 VSUBS 0.01013f
C176 B.n88 VSUBS 0.01013f
C177 B.n89 VSUBS 0.01013f
C178 B.n90 VSUBS 0.01013f
C179 B.n91 VSUBS 0.01013f
C180 B.n92 VSUBS 0.01013f
C181 B.n93 VSUBS 0.01013f
C182 B.n94 VSUBS 0.01013f
C183 B.n95 VSUBS 0.01013f
C184 B.n96 VSUBS 0.01013f
C185 B.n97 VSUBS 0.01013f
C186 B.n98 VSUBS 0.01013f
C187 B.n99 VSUBS 0.01013f
C188 B.n100 VSUBS 0.01013f
C189 B.n101 VSUBS 0.01013f
C190 B.n102 VSUBS 0.01013f
C191 B.n103 VSUBS 0.01013f
C192 B.n104 VSUBS 0.01013f
C193 B.n105 VSUBS 0.01013f
C194 B.n106 VSUBS 0.01013f
C195 B.n107 VSUBS 0.01013f
C196 B.n108 VSUBS 0.01013f
C197 B.n109 VSUBS 0.01013f
C198 B.n110 VSUBS 0.01013f
C199 B.n111 VSUBS 0.01013f
C200 B.n112 VSUBS 0.01013f
C201 B.n113 VSUBS 0.01013f
C202 B.n114 VSUBS 0.01013f
C203 B.n115 VSUBS 0.01013f
C204 B.n116 VSUBS 0.01013f
C205 B.n117 VSUBS 0.01013f
C206 B.n118 VSUBS 0.01013f
C207 B.n119 VSUBS 0.01013f
C208 B.n120 VSUBS 0.01013f
C209 B.n121 VSUBS 0.01013f
C210 B.n122 VSUBS 0.01013f
C211 B.n123 VSUBS 0.01013f
C212 B.n124 VSUBS 0.01013f
C213 B.n125 VSUBS 0.01013f
C214 B.n126 VSUBS 0.01013f
C215 B.n127 VSUBS 0.01013f
C216 B.n128 VSUBS 0.01013f
C217 B.n129 VSUBS 0.01013f
C218 B.n130 VSUBS 0.023794f
C219 B.n131 VSUBS 0.025369f
C220 B.n132 VSUBS 0.025369f
C221 B.n133 VSUBS 0.01013f
C222 B.n134 VSUBS 0.01013f
C223 B.n135 VSUBS 0.01013f
C224 B.n136 VSUBS 0.01013f
C225 B.n137 VSUBS 0.01013f
C226 B.n138 VSUBS 0.01013f
C227 B.n139 VSUBS 0.01013f
C228 B.n140 VSUBS 0.01013f
C229 B.n141 VSUBS 0.01013f
C230 B.n142 VSUBS 0.01013f
C231 B.n143 VSUBS 0.007002f
C232 B.n144 VSUBS 0.01013f
C233 B.n145 VSUBS 0.01013f
C234 B.n146 VSUBS 0.008194f
C235 B.n147 VSUBS 0.01013f
C236 B.n148 VSUBS 0.01013f
C237 B.n149 VSUBS 0.01013f
C238 B.n150 VSUBS 0.01013f
C239 B.n151 VSUBS 0.01013f
C240 B.n152 VSUBS 0.01013f
C241 B.n153 VSUBS 0.01013f
C242 B.n154 VSUBS 0.01013f
C243 B.n155 VSUBS 0.01013f
C244 B.n156 VSUBS 0.01013f
C245 B.n157 VSUBS 0.01013f
C246 B.n158 VSUBS 0.008194f
C247 B.n159 VSUBS 0.023471f
C248 B.n160 VSUBS 0.007002f
C249 B.n161 VSUBS 0.01013f
C250 B.n162 VSUBS 0.01013f
C251 B.n163 VSUBS 0.01013f
C252 B.n164 VSUBS 0.01013f
C253 B.n165 VSUBS 0.01013f
C254 B.n166 VSUBS 0.01013f
C255 B.n167 VSUBS 0.01013f
C256 B.n168 VSUBS 0.01013f
C257 B.n169 VSUBS 0.01013f
C258 B.n170 VSUBS 0.01013f
C259 B.n171 VSUBS 0.01013f
C260 B.n172 VSUBS 0.025369f
C261 B.n173 VSUBS 0.023794f
C262 B.n174 VSUBS 0.023794f
C263 B.n175 VSUBS 0.01013f
C264 B.n176 VSUBS 0.01013f
C265 B.n177 VSUBS 0.01013f
C266 B.n178 VSUBS 0.01013f
C267 B.n179 VSUBS 0.01013f
C268 B.n180 VSUBS 0.01013f
C269 B.n181 VSUBS 0.01013f
C270 B.n182 VSUBS 0.01013f
C271 B.n183 VSUBS 0.01013f
C272 B.n184 VSUBS 0.01013f
C273 B.n185 VSUBS 0.01013f
C274 B.n186 VSUBS 0.01013f
C275 B.n187 VSUBS 0.01013f
C276 B.n188 VSUBS 0.01013f
C277 B.n189 VSUBS 0.01013f
C278 B.n190 VSUBS 0.01013f
C279 B.n191 VSUBS 0.01013f
C280 B.n192 VSUBS 0.01013f
C281 B.n193 VSUBS 0.01013f
C282 B.n194 VSUBS 0.01013f
C283 B.n195 VSUBS 0.01013f
C284 B.n196 VSUBS 0.01013f
C285 B.n197 VSUBS 0.01013f
C286 B.n198 VSUBS 0.01013f
C287 B.n199 VSUBS 0.01013f
C288 B.n200 VSUBS 0.01013f
C289 B.n201 VSUBS 0.01013f
C290 B.n202 VSUBS 0.01013f
C291 B.n203 VSUBS 0.01013f
C292 B.n204 VSUBS 0.01013f
C293 B.n205 VSUBS 0.01013f
C294 B.n206 VSUBS 0.01013f
C295 B.n207 VSUBS 0.01013f
C296 B.n208 VSUBS 0.01013f
C297 B.n209 VSUBS 0.01013f
C298 B.n210 VSUBS 0.01013f
C299 B.n211 VSUBS 0.01013f
C300 B.n212 VSUBS 0.01013f
C301 B.n213 VSUBS 0.01013f
C302 B.n214 VSUBS 0.01013f
C303 B.n215 VSUBS 0.01013f
C304 B.n216 VSUBS 0.01013f
C305 B.n217 VSUBS 0.01013f
C306 B.n218 VSUBS 0.01013f
C307 B.n219 VSUBS 0.01013f
C308 B.n220 VSUBS 0.01013f
C309 B.n221 VSUBS 0.01013f
C310 B.n222 VSUBS 0.01013f
C311 B.n223 VSUBS 0.01013f
C312 B.n224 VSUBS 0.01013f
C313 B.n225 VSUBS 0.01013f
C314 B.n226 VSUBS 0.01013f
C315 B.n227 VSUBS 0.01013f
C316 B.n228 VSUBS 0.01013f
C317 B.n229 VSUBS 0.01013f
C318 B.n230 VSUBS 0.01013f
C319 B.n231 VSUBS 0.01013f
C320 B.n232 VSUBS 0.01013f
C321 B.n233 VSUBS 0.01013f
C322 B.n234 VSUBS 0.01013f
C323 B.n235 VSUBS 0.01013f
C324 B.n236 VSUBS 0.01013f
C325 B.n237 VSUBS 0.01013f
C326 B.n238 VSUBS 0.01013f
C327 B.n239 VSUBS 0.01013f
C328 B.n240 VSUBS 0.01013f
C329 B.n241 VSUBS 0.01013f
C330 B.n242 VSUBS 0.01013f
C331 B.n243 VSUBS 0.01013f
C332 B.n244 VSUBS 0.01013f
C333 B.n245 VSUBS 0.01013f
C334 B.n246 VSUBS 0.01013f
C335 B.n247 VSUBS 0.01013f
C336 B.n248 VSUBS 0.01013f
C337 B.n249 VSUBS 0.01013f
C338 B.n250 VSUBS 0.01013f
C339 B.n251 VSUBS 0.01013f
C340 B.n252 VSUBS 0.01013f
C341 B.n253 VSUBS 0.01013f
C342 B.n254 VSUBS 0.023794f
C343 B.n255 VSUBS 0.024927f
C344 B.n256 VSUBS 0.024236f
C345 B.n257 VSUBS 0.01013f
C346 B.n258 VSUBS 0.01013f
C347 B.n259 VSUBS 0.01013f
C348 B.n260 VSUBS 0.01013f
C349 B.n261 VSUBS 0.01013f
C350 B.n262 VSUBS 0.01013f
C351 B.n263 VSUBS 0.01013f
C352 B.n264 VSUBS 0.01013f
C353 B.n265 VSUBS 0.01013f
C354 B.n266 VSUBS 0.01013f
C355 B.n267 VSUBS 0.01013f
C356 B.n268 VSUBS 0.007002f
C357 B.n269 VSUBS 0.023471f
C358 B.n270 VSUBS 0.008194f
C359 B.n271 VSUBS 0.01013f
C360 B.n272 VSUBS 0.01013f
C361 B.n273 VSUBS 0.01013f
C362 B.n274 VSUBS 0.01013f
C363 B.n275 VSUBS 0.01013f
C364 B.n276 VSUBS 0.01013f
C365 B.n277 VSUBS 0.01013f
C366 B.n278 VSUBS 0.01013f
C367 B.n279 VSUBS 0.01013f
C368 B.n280 VSUBS 0.01013f
C369 B.n281 VSUBS 0.01013f
C370 B.n282 VSUBS 0.008194f
C371 B.n283 VSUBS 0.01013f
C372 B.n284 VSUBS 0.01013f
C373 B.n285 VSUBS 0.007002f
C374 B.n286 VSUBS 0.01013f
C375 B.n287 VSUBS 0.01013f
C376 B.n288 VSUBS 0.01013f
C377 B.n289 VSUBS 0.01013f
C378 B.n290 VSUBS 0.01013f
C379 B.n291 VSUBS 0.01013f
C380 B.n292 VSUBS 0.01013f
C381 B.n293 VSUBS 0.01013f
C382 B.n294 VSUBS 0.01013f
C383 B.n295 VSUBS 0.01013f
C384 B.n296 VSUBS 0.025369f
C385 B.n297 VSUBS 0.025369f
C386 B.n298 VSUBS 0.023794f
C387 B.n299 VSUBS 0.01013f
C388 B.n300 VSUBS 0.01013f
C389 B.n301 VSUBS 0.01013f
C390 B.n302 VSUBS 0.01013f
C391 B.n303 VSUBS 0.01013f
C392 B.n304 VSUBS 0.01013f
C393 B.n305 VSUBS 0.01013f
C394 B.n306 VSUBS 0.01013f
C395 B.n307 VSUBS 0.01013f
C396 B.n308 VSUBS 0.01013f
C397 B.n309 VSUBS 0.01013f
C398 B.n310 VSUBS 0.01013f
C399 B.n311 VSUBS 0.01013f
C400 B.n312 VSUBS 0.01013f
C401 B.n313 VSUBS 0.01013f
C402 B.n314 VSUBS 0.01013f
C403 B.n315 VSUBS 0.01013f
C404 B.n316 VSUBS 0.01013f
C405 B.n317 VSUBS 0.01013f
C406 B.n318 VSUBS 0.01013f
C407 B.n319 VSUBS 0.01013f
C408 B.n320 VSUBS 0.01013f
C409 B.n321 VSUBS 0.01013f
C410 B.n322 VSUBS 0.01013f
C411 B.n323 VSUBS 0.01013f
C412 B.n324 VSUBS 0.01013f
C413 B.n325 VSUBS 0.01013f
C414 B.n326 VSUBS 0.01013f
C415 B.n327 VSUBS 0.01013f
C416 B.n328 VSUBS 0.01013f
C417 B.n329 VSUBS 0.01013f
C418 B.n330 VSUBS 0.01013f
C419 B.n331 VSUBS 0.01013f
C420 B.n332 VSUBS 0.01013f
C421 B.n333 VSUBS 0.01013f
C422 B.n334 VSUBS 0.01013f
C423 B.n335 VSUBS 0.01013f
C424 B.n336 VSUBS 0.01013f
C425 B.n337 VSUBS 0.01013f
C426 B.n338 VSUBS 0.01013f
C427 B.n339 VSUBS 0.022939f
C428 VTAIL.t7 VSUBS 0.018956f
C429 VTAIL.t1 VSUBS 0.018956f
C430 VTAIL.n0 VSUBS 0.038754f
C431 VTAIL.n1 VSUBS 0.157796f
C432 VTAIL.t6 VSUBS 0.086063f
C433 VTAIL.n2 VSUBS 0.201958f
C434 VTAIL.t12 VSUBS 0.086063f
C435 VTAIL.n3 VSUBS 0.201958f
C436 VTAIL.t8 VSUBS 0.018956f
C437 VTAIL.t15 VSUBS 0.018956f
C438 VTAIL.n4 VSUBS 0.038754f
C439 VTAIL.n5 VSUBS 0.260454f
C440 VTAIL.t14 VSUBS 0.086063f
C441 VTAIL.n6 VSUBS 0.738795f
C442 VTAIL.t0 VSUBS 0.086063f
C443 VTAIL.n7 VSUBS 0.738795f
C444 VTAIL.t5 VSUBS 0.018956f
C445 VTAIL.t2 VSUBS 0.018956f
C446 VTAIL.n8 VSUBS 0.038754f
C447 VTAIL.n9 VSUBS 0.260454f
C448 VTAIL.t4 VSUBS 0.086063f
C449 VTAIL.n10 VSUBS 0.201958f
C450 VTAIL.t10 VSUBS 0.086063f
C451 VTAIL.n11 VSUBS 0.201958f
C452 VTAIL.t13 VSUBS 0.018956f
C453 VTAIL.t11 VSUBS 0.018956f
C454 VTAIL.n12 VSUBS 0.038754f
C455 VTAIL.n13 VSUBS 0.260454f
C456 VTAIL.t9 VSUBS 0.086063f
C457 VTAIL.n14 VSUBS 0.738795f
C458 VTAIL.t3 VSUBS 0.086063f
C459 VTAIL.n15 VSUBS 0.733173f
C460 VDD1.t3 VSUBS 0.013449f
C461 VDD1.t4 VSUBS 0.013449f
C462 VDD1.n0 VSUBS 0.029141f
C463 VDD1.t6 VSUBS 0.013449f
C464 VDD1.t0 VSUBS 0.013449f
C465 VDD1.n1 VSUBS 0.029102f
C466 VDD1.t7 VSUBS 0.013449f
C467 VDD1.t5 VSUBS 0.013449f
C468 VDD1.n2 VSUBS 0.029102f
C469 VDD1.n3 VSUBS 1.2393f
C470 VDD1.t1 VSUBS 0.013449f
C471 VDD1.t2 VSUBS 0.013449f
C472 VDD1.n4 VSUBS 0.02896f
C473 VDD1.n5 VSUBS 1.17377f
C474 VP.n0 VSUBS 0.084247f
C475 VP.t0 VSUBS 0.080093f
C476 VP.n1 VSUBS 0.050993f
C477 VP.n2 VSUBS 0.084247f
C478 VP.t7 VSUBS 0.080093f
C479 VP.n3 VSUBS 0.084247f
C480 VP.t6 VSUBS 0.173344f
C481 VP.t4 VSUBS 0.080093f
C482 VP.n4 VSUBS 0.050993f
C483 VP.t5 VSUBS 0.212302f
C484 VP.n5 VSUBS 0.188603f
C485 VP.t2 VSUBS 0.080093f
C486 VP.n6 VSUBS 0.15588f
C487 VP.n7 VSUBS 0.084361f
C488 VP.n8 VSUBS 0.265651f
C489 VP.n9 VSUBS 0.063136f
C490 VP.n10 VSUBS 0.063136f
C491 VP.n11 VSUBS 0.084361f
C492 VP.n12 VSUBS 0.103566f
C493 VP.n13 VSUBS 0.082553f
C494 VP.n14 VSUBS 0.196029f
C495 VP.n15 VSUBS 1.8991f
C496 VP.n16 VSUBS 1.96421f
C497 VP.t1 VSUBS 0.173344f
C498 VP.n17 VSUBS 0.196029f
C499 VP.n18 VSUBS 0.082553f
C500 VP.n19 VSUBS 0.103566f
C501 VP.n20 VSUBS 0.084361f
C502 VP.n21 VSUBS 0.063136f
C503 VP.n22 VSUBS 0.063136f
C504 VP.n23 VSUBS 0.063136f
C505 VP.n24 VSUBS 0.084361f
C506 VP.n25 VSUBS 0.103566f
C507 VP.n26 VSUBS 0.082553f
C508 VP.t3 VSUBS 0.173344f
C509 VP.n27 VSUBS 0.196029f
C510 VP.n28 VSUBS 0.059129f
.ends

