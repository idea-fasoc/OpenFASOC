* NGSPICE file created from diff_pair_sample_0607.ext - technology: sky130A

.subckt diff_pair_sample_0607 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t7 VN.t0 VTAIL.t3 B.t7 sky130_fd_pr__nfet_01v8 ad=2.83965 pd=17.54 as=6.7119 ps=35.2 w=17.21 l=0.56
X1 VDD1.t7 VP.t0 VTAIL.t15 B.t2 sky130_fd_pr__nfet_01v8 ad=2.83965 pd=17.54 as=6.7119 ps=35.2 w=17.21 l=0.56
X2 VTAIL.t9 VN.t1 VDD2.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=6.7119 pd=35.2 as=2.83965 ps=17.54 w=17.21 l=0.56
X3 VTAIL.t8 VN.t2 VDD2.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.83965 pd=17.54 as=2.83965 ps=17.54 w=17.21 l=0.56
X4 B.t21 B.t19 B.t20 B.t16 sky130_fd_pr__nfet_01v8 ad=6.7119 pd=35.2 as=0 ps=0 w=17.21 l=0.56
X5 VDD2.t4 VN.t3 VTAIL.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=2.83965 pd=17.54 as=2.83965 ps=17.54 w=17.21 l=0.56
X6 B.t18 B.t15 B.t17 B.t16 sky130_fd_pr__nfet_01v8 ad=6.7119 pd=35.2 as=0 ps=0 w=17.21 l=0.56
X7 VTAIL.t10 VP.t1 VDD1.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=6.7119 pd=35.2 as=2.83965 ps=17.54 w=17.21 l=0.56
X8 VTAIL.t4 VN.t4 VDD2.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=6.7119 pd=35.2 as=2.83965 ps=17.54 w=17.21 l=0.56
X9 VTAIL.t6 VN.t5 VDD2.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=2.83965 pd=17.54 as=2.83965 ps=17.54 w=17.21 l=0.56
X10 VTAIL.t1 VP.t2 VDD1.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=2.83965 pd=17.54 as=2.83965 ps=17.54 w=17.21 l=0.56
X11 VDD2.t1 VN.t6 VTAIL.t7 B.t0 sky130_fd_pr__nfet_01v8 ad=2.83965 pd=17.54 as=2.83965 ps=17.54 w=17.21 l=0.56
X12 VDD2.t0 VN.t7 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.83965 pd=17.54 as=6.7119 ps=35.2 w=17.21 l=0.56
X13 VTAIL.t14 VP.t3 VDD1.t4 B.t6 sky130_fd_pr__nfet_01v8 ad=6.7119 pd=35.2 as=2.83965 ps=17.54 w=17.21 l=0.56
X14 VDD1.t3 VP.t4 VTAIL.t13 B.t7 sky130_fd_pr__nfet_01v8 ad=2.83965 pd=17.54 as=6.7119 ps=35.2 w=17.21 l=0.56
X15 VDD1.t2 VP.t5 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.83965 pd=17.54 as=2.83965 ps=17.54 w=17.21 l=0.56
X16 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=6.7119 pd=35.2 as=0 ps=0 w=17.21 l=0.56
X17 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=6.7119 pd=35.2 as=0 ps=0 w=17.21 l=0.56
X18 VDD1.t1 VP.t6 VTAIL.t12 B.t4 sky130_fd_pr__nfet_01v8 ad=2.83965 pd=17.54 as=2.83965 ps=17.54 w=17.21 l=0.56
X19 VTAIL.t11 VP.t7 VDD1.t0 B.t5 sky130_fd_pr__nfet_01v8 ad=2.83965 pd=17.54 as=2.83965 ps=17.54 w=17.21 l=0.56
R0 VN.n2 VN.t4 837.266
R1 VN.n10 VN.t7 837.266
R2 VN.n1 VN.t3 811.223
R3 VN.n4 VN.t5 811.223
R4 VN.n6 VN.t0 811.223
R5 VN.n9 VN.t2 811.223
R6 VN.n12 VN.t6 811.223
R7 VN.n14 VN.t1 811.223
R8 VN.n7 VN.n6 161.3
R9 VN.n15 VN.n14 161.3
R10 VN.n13 VN.n8 161.3
R11 VN.n12 VN.n11 161.3
R12 VN.n5 VN.n0 161.3
R13 VN.n4 VN.n3 161.3
R14 VN.n4 VN.n1 48.2005
R15 VN.n12 VN.n9 48.2005
R16 VN VN.n15 45.6615
R17 VN.n11 VN.n10 45.057
R18 VN.n3 VN.n2 45.057
R19 VN.n6 VN.n5 44.549
R20 VN.n14 VN.n13 44.549
R21 VN.n2 VN.n1 14.6494
R22 VN.n10 VN.n9 14.6494
R23 VN.n5 VN.n4 3.65202
R24 VN.n13 VN.n12 3.65202
R25 VN.n15 VN.n8 0.189894
R26 VN.n11 VN.n8 0.189894
R27 VN.n3 VN.n0 0.189894
R28 VN.n7 VN.n0 0.189894
R29 VN VN.n7 0.0516364
R30 VTAIL.n11 VTAIL.t10 46.1434
R31 VTAIL.n10 VTAIL.t2 46.1434
R32 VTAIL.n7 VTAIL.t9 46.1434
R33 VTAIL.n15 VTAIL.t3 46.1433
R34 VTAIL.n2 VTAIL.t4 46.1433
R35 VTAIL.n3 VTAIL.t15 46.1433
R36 VTAIL.n6 VTAIL.t14 46.1433
R37 VTAIL.n14 VTAIL.t13 46.1433
R38 VTAIL.n13 VTAIL.n12 44.993
R39 VTAIL.n9 VTAIL.n8 44.993
R40 VTAIL.n1 VTAIL.n0 44.9927
R41 VTAIL.n5 VTAIL.n4 44.9927
R42 VTAIL.n15 VTAIL.n14 27.9703
R43 VTAIL.n7 VTAIL.n6 27.9703
R44 VTAIL.n0 VTAIL.t5 1.15099
R45 VTAIL.n0 VTAIL.t6 1.15099
R46 VTAIL.n4 VTAIL.t0 1.15099
R47 VTAIL.n4 VTAIL.t11 1.15099
R48 VTAIL.n12 VTAIL.t12 1.15099
R49 VTAIL.n12 VTAIL.t1 1.15099
R50 VTAIL.n8 VTAIL.t7 1.15099
R51 VTAIL.n8 VTAIL.t8 1.15099
R52 VTAIL.n9 VTAIL.n7 0.767741
R53 VTAIL.n10 VTAIL.n9 0.767741
R54 VTAIL.n13 VTAIL.n11 0.767741
R55 VTAIL.n14 VTAIL.n13 0.767741
R56 VTAIL.n6 VTAIL.n5 0.767741
R57 VTAIL.n5 VTAIL.n3 0.767741
R58 VTAIL.n2 VTAIL.n1 0.767741
R59 VTAIL VTAIL.n15 0.709552
R60 VTAIL.n11 VTAIL.n10 0.470328
R61 VTAIL.n3 VTAIL.n2 0.470328
R62 VTAIL VTAIL.n1 0.0586897
R63 VDD2.n2 VDD2.n1 61.9998
R64 VDD2.n2 VDD2.n0 61.9998
R65 VDD2 VDD2.n5 61.997
R66 VDD2.n4 VDD2.n3 61.6718
R67 VDD2.n4 VDD2.n2 42.0041
R68 VDD2.n5 VDD2.t5 1.15099
R69 VDD2.n5 VDD2.t0 1.15099
R70 VDD2.n3 VDD2.t6 1.15099
R71 VDD2.n3 VDD2.t1 1.15099
R72 VDD2.n1 VDD2.t2 1.15099
R73 VDD2.n1 VDD2.t7 1.15099
R74 VDD2.n0 VDD2.t3 1.15099
R75 VDD2.n0 VDD2.t4 1.15099
R76 VDD2 VDD2.n4 0.44231
R77 B.n457 B.t15 945.761
R78 B.n454 B.t19 945.761
R79 B.n107 B.t12 945.761
R80 B.n104 B.t8 945.761
R81 B.n797 B.n796 585
R82 B.n798 B.n797 585
R83 B.n352 B.n103 585
R84 B.n351 B.n350 585
R85 B.n349 B.n348 585
R86 B.n347 B.n346 585
R87 B.n345 B.n344 585
R88 B.n343 B.n342 585
R89 B.n341 B.n340 585
R90 B.n339 B.n338 585
R91 B.n337 B.n336 585
R92 B.n335 B.n334 585
R93 B.n333 B.n332 585
R94 B.n331 B.n330 585
R95 B.n329 B.n328 585
R96 B.n327 B.n326 585
R97 B.n325 B.n324 585
R98 B.n323 B.n322 585
R99 B.n321 B.n320 585
R100 B.n319 B.n318 585
R101 B.n317 B.n316 585
R102 B.n315 B.n314 585
R103 B.n313 B.n312 585
R104 B.n311 B.n310 585
R105 B.n309 B.n308 585
R106 B.n307 B.n306 585
R107 B.n305 B.n304 585
R108 B.n303 B.n302 585
R109 B.n301 B.n300 585
R110 B.n299 B.n298 585
R111 B.n297 B.n296 585
R112 B.n295 B.n294 585
R113 B.n293 B.n292 585
R114 B.n291 B.n290 585
R115 B.n289 B.n288 585
R116 B.n287 B.n286 585
R117 B.n285 B.n284 585
R118 B.n283 B.n282 585
R119 B.n281 B.n280 585
R120 B.n279 B.n278 585
R121 B.n277 B.n276 585
R122 B.n275 B.n274 585
R123 B.n273 B.n272 585
R124 B.n271 B.n270 585
R125 B.n269 B.n268 585
R126 B.n267 B.n266 585
R127 B.n265 B.n264 585
R128 B.n263 B.n262 585
R129 B.n261 B.n260 585
R130 B.n259 B.n258 585
R131 B.n257 B.n256 585
R132 B.n255 B.n254 585
R133 B.n253 B.n252 585
R134 B.n251 B.n250 585
R135 B.n249 B.n248 585
R136 B.n247 B.n246 585
R137 B.n245 B.n244 585
R138 B.n243 B.n242 585
R139 B.n241 B.n240 585
R140 B.n239 B.n238 585
R141 B.n237 B.n236 585
R142 B.n235 B.n234 585
R143 B.n233 B.n232 585
R144 B.n231 B.n230 585
R145 B.n229 B.n228 585
R146 B.n227 B.n226 585
R147 B.n225 B.n224 585
R148 B.n222 B.n221 585
R149 B.n220 B.n219 585
R150 B.n218 B.n217 585
R151 B.n216 B.n215 585
R152 B.n214 B.n213 585
R153 B.n212 B.n211 585
R154 B.n210 B.n209 585
R155 B.n208 B.n207 585
R156 B.n206 B.n205 585
R157 B.n204 B.n203 585
R158 B.n202 B.n201 585
R159 B.n200 B.n199 585
R160 B.n198 B.n197 585
R161 B.n196 B.n195 585
R162 B.n194 B.n193 585
R163 B.n192 B.n191 585
R164 B.n190 B.n189 585
R165 B.n188 B.n187 585
R166 B.n186 B.n185 585
R167 B.n184 B.n183 585
R168 B.n182 B.n181 585
R169 B.n180 B.n179 585
R170 B.n178 B.n177 585
R171 B.n176 B.n175 585
R172 B.n174 B.n173 585
R173 B.n172 B.n171 585
R174 B.n170 B.n169 585
R175 B.n168 B.n167 585
R176 B.n166 B.n165 585
R177 B.n164 B.n163 585
R178 B.n162 B.n161 585
R179 B.n160 B.n159 585
R180 B.n158 B.n157 585
R181 B.n156 B.n155 585
R182 B.n154 B.n153 585
R183 B.n152 B.n151 585
R184 B.n150 B.n149 585
R185 B.n148 B.n147 585
R186 B.n146 B.n145 585
R187 B.n144 B.n143 585
R188 B.n142 B.n141 585
R189 B.n140 B.n139 585
R190 B.n138 B.n137 585
R191 B.n136 B.n135 585
R192 B.n134 B.n133 585
R193 B.n132 B.n131 585
R194 B.n130 B.n129 585
R195 B.n128 B.n127 585
R196 B.n126 B.n125 585
R197 B.n124 B.n123 585
R198 B.n122 B.n121 585
R199 B.n120 B.n119 585
R200 B.n118 B.n117 585
R201 B.n116 B.n115 585
R202 B.n114 B.n113 585
R203 B.n112 B.n111 585
R204 B.n110 B.n109 585
R205 B.n795 B.n41 585
R206 B.n799 B.n41 585
R207 B.n794 B.n40 585
R208 B.n800 B.n40 585
R209 B.n793 B.n792 585
R210 B.n792 B.n36 585
R211 B.n791 B.n35 585
R212 B.n806 B.n35 585
R213 B.n790 B.n34 585
R214 B.n807 B.n34 585
R215 B.n789 B.n33 585
R216 B.n808 B.n33 585
R217 B.n788 B.n787 585
R218 B.n787 B.n29 585
R219 B.n786 B.n28 585
R220 B.n814 B.n28 585
R221 B.n785 B.n27 585
R222 B.n815 B.n27 585
R223 B.n784 B.n26 585
R224 B.n816 B.n26 585
R225 B.n783 B.n782 585
R226 B.n782 B.n25 585
R227 B.n781 B.n21 585
R228 B.n822 B.n21 585
R229 B.n780 B.n20 585
R230 B.n823 B.n20 585
R231 B.n779 B.n19 585
R232 B.n824 B.n19 585
R233 B.n778 B.n777 585
R234 B.n777 B.n15 585
R235 B.n776 B.n14 585
R236 B.n830 B.n14 585
R237 B.n775 B.n13 585
R238 B.n831 B.n13 585
R239 B.n774 B.n12 585
R240 B.n832 B.n12 585
R241 B.n773 B.n772 585
R242 B.n772 B.n11 585
R243 B.n771 B.n7 585
R244 B.n838 B.n7 585
R245 B.n770 B.n6 585
R246 B.n839 B.n6 585
R247 B.n769 B.n5 585
R248 B.n840 B.n5 585
R249 B.n768 B.n767 585
R250 B.n767 B.n4 585
R251 B.n766 B.n353 585
R252 B.n766 B.n765 585
R253 B.n755 B.n354 585
R254 B.n758 B.n354 585
R255 B.n757 B.n756 585
R256 B.n759 B.n757 585
R257 B.n754 B.n359 585
R258 B.n359 B.n358 585
R259 B.n753 B.n752 585
R260 B.n752 B.n751 585
R261 B.n361 B.n360 585
R262 B.n362 B.n361 585
R263 B.n744 B.n743 585
R264 B.n745 B.n744 585
R265 B.n742 B.n366 585
R266 B.n369 B.n366 585
R267 B.n741 B.n740 585
R268 B.n740 B.n739 585
R269 B.n368 B.n367 585
R270 B.n732 B.n368 585
R271 B.n731 B.n730 585
R272 B.n733 B.n731 585
R273 B.n729 B.n374 585
R274 B.n374 B.n373 585
R275 B.n728 B.n727 585
R276 B.n727 B.n726 585
R277 B.n376 B.n375 585
R278 B.n377 B.n376 585
R279 B.n719 B.n718 585
R280 B.n720 B.n719 585
R281 B.n717 B.n381 585
R282 B.n385 B.n381 585
R283 B.n716 B.n715 585
R284 B.n715 B.n714 585
R285 B.n383 B.n382 585
R286 B.n384 B.n383 585
R287 B.n707 B.n706 585
R288 B.n708 B.n707 585
R289 B.n705 B.n390 585
R290 B.n390 B.n389 585
R291 B.n699 B.n698 585
R292 B.n697 B.n453 585
R293 B.n696 B.n452 585
R294 B.n701 B.n452 585
R295 B.n695 B.n694 585
R296 B.n693 B.n692 585
R297 B.n691 B.n690 585
R298 B.n689 B.n688 585
R299 B.n687 B.n686 585
R300 B.n685 B.n684 585
R301 B.n683 B.n682 585
R302 B.n681 B.n680 585
R303 B.n679 B.n678 585
R304 B.n677 B.n676 585
R305 B.n675 B.n674 585
R306 B.n673 B.n672 585
R307 B.n671 B.n670 585
R308 B.n669 B.n668 585
R309 B.n667 B.n666 585
R310 B.n665 B.n664 585
R311 B.n663 B.n662 585
R312 B.n661 B.n660 585
R313 B.n659 B.n658 585
R314 B.n657 B.n656 585
R315 B.n655 B.n654 585
R316 B.n653 B.n652 585
R317 B.n651 B.n650 585
R318 B.n649 B.n648 585
R319 B.n647 B.n646 585
R320 B.n645 B.n644 585
R321 B.n643 B.n642 585
R322 B.n641 B.n640 585
R323 B.n639 B.n638 585
R324 B.n637 B.n636 585
R325 B.n635 B.n634 585
R326 B.n633 B.n632 585
R327 B.n631 B.n630 585
R328 B.n629 B.n628 585
R329 B.n627 B.n626 585
R330 B.n625 B.n624 585
R331 B.n623 B.n622 585
R332 B.n621 B.n620 585
R333 B.n619 B.n618 585
R334 B.n617 B.n616 585
R335 B.n615 B.n614 585
R336 B.n613 B.n612 585
R337 B.n611 B.n610 585
R338 B.n609 B.n608 585
R339 B.n607 B.n606 585
R340 B.n605 B.n604 585
R341 B.n603 B.n602 585
R342 B.n601 B.n600 585
R343 B.n599 B.n598 585
R344 B.n597 B.n596 585
R345 B.n595 B.n594 585
R346 B.n593 B.n592 585
R347 B.n591 B.n590 585
R348 B.n589 B.n588 585
R349 B.n587 B.n586 585
R350 B.n585 B.n584 585
R351 B.n583 B.n582 585
R352 B.n581 B.n580 585
R353 B.n579 B.n578 585
R354 B.n577 B.n576 585
R355 B.n575 B.n574 585
R356 B.n573 B.n572 585
R357 B.n571 B.n570 585
R358 B.n568 B.n567 585
R359 B.n566 B.n565 585
R360 B.n564 B.n563 585
R361 B.n562 B.n561 585
R362 B.n560 B.n559 585
R363 B.n558 B.n557 585
R364 B.n556 B.n555 585
R365 B.n554 B.n553 585
R366 B.n552 B.n551 585
R367 B.n550 B.n549 585
R368 B.n548 B.n547 585
R369 B.n546 B.n545 585
R370 B.n544 B.n543 585
R371 B.n542 B.n541 585
R372 B.n540 B.n539 585
R373 B.n538 B.n537 585
R374 B.n536 B.n535 585
R375 B.n534 B.n533 585
R376 B.n532 B.n531 585
R377 B.n530 B.n529 585
R378 B.n528 B.n527 585
R379 B.n526 B.n525 585
R380 B.n524 B.n523 585
R381 B.n522 B.n521 585
R382 B.n520 B.n519 585
R383 B.n518 B.n517 585
R384 B.n516 B.n515 585
R385 B.n514 B.n513 585
R386 B.n512 B.n511 585
R387 B.n510 B.n509 585
R388 B.n508 B.n507 585
R389 B.n506 B.n505 585
R390 B.n504 B.n503 585
R391 B.n502 B.n501 585
R392 B.n500 B.n499 585
R393 B.n498 B.n497 585
R394 B.n496 B.n495 585
R395 B.n494 B.n493 585
R396 B.n492 B.n491 585
R397 B.n490 B.n489 585
R398 B.n488 B.n487 585
R399 B.n486 B.n485 585
R400 B.n484 B.n483 585
R401 B.n482 B.n481 585
R402 B.n480 B.n479 585
R403 B.n478 B.n477 585
R404 B.n476 B.n475 585
R405 B.n474 B.n473 585
R406 B.n472 B.n471 585
R407 B.n470 B.n469 585
R408 B.n468 B.n467 585
R409 B.n466 B.n465 585
R410 B.n464 B.n463 585
R411 B.n462 B.n461 585
R412 B.n460 B.n459 585
R413 B.n392 B.n391 585
R414 B.n704 B.n703 585
R415 B.n388 B.n387 585
R416 B.n389 B.n388 585
R417 B.n710 B.n709 585
R418 B.n709 B.n708 585
R419 B.n711 B.n386 585
R420 B.n386 B.n384 585
R421 B.n713 B.n712 585
R422 B.n714 B.n713 585
R423 B.n380 B.n379 585
R424 B.n385 B.n380 585
R425 B.n722 B.n721 585
R426 B.n721 B.n720 585
R427 B.n723 B.n378 585
R428 B.n378 B.n377 585
R429 B.n725 B.n724 585
R430 B.n726 B.n725 585
R431 B.n372 B.n371 585
R432 B.n373 B.n372 585
R433 B.n735 B.n734 585
R434 B.n734 B.n733 585
R435 B.n736 B.n370 585
R436 B.n732 B.n370 585
R437 B.n738 B.n737 585
R438 B.n739 B.n738 585
R439 B.n365 B.n364 585
R440 B.n369 B.n365 585
R441 B.n747 B.n746 585
R442 B.n746 B.n745 585
R443 B.n748 B.n363 585
R444 B.n363 B.n362 585
R445 B.n750 B.n749 585
R446 B.n751 B.n750 585
R447 B.n357 B.n356 585
R448 B.n358 B.n357 585
R449 B.n761 B.n760 585
R450 B.n760 B.n759 585
R451 B.n762 B.n355 585
R452 B.n758 B.n355 585
R453 B.n764 B.n763 585
R454 B.n765 B.n764 585
R455 B.n2 B.n0 585
R456 B.n4 B.n2 585
R457 B.n3 B.n1 585
R458 B.n839 B.n3 585
R459 B.n837 B.n836 585
R460 B.n838 B.n837 585
R461 B.n835 B.n8 585
R462 B.n11 B.n8 585
R463 B.n834 B.n833 585
R464 B.n833 B.n832 585
R465 B.n10 B.n9 585
R466 B.n831 B.n10 585
R467 B.n829 B.n828 585
R468 B.n830 B.n829 585
R469 B.n827 B.n16 585
R470 B.n16 B.n15 585
R471 B.n826 B.n825 585
R472 B.n825 B.n824 585
R473 B.n18 B.n17 585
R474 B.n823 B.n18 585
R475 B.n821 B.n820 585
R476 B.n822 B.n821 585
R477 B.n819 B.n22 585
R478 B.n25 B.n22 585
R479 B.n818 B.n817 585
R480 B.n817 B.n816 585
R481 B.n24 B.n23 585
R482 B.n815 B.n24 585
R483 B.n813 B.n812 585
R484 B.n814 B.n813 585
R485 B.n811 B.n30 585
R486 B.n30 B.n29 585
R487 B.n810 B.n809 585
R488 B.n809 B.n808 585
R489 B.n32 B.n31 585
R490 B.n807 B.n32 585
R491 B.n805 B.n804 585
R492 B.n806 B.n805 585
R493 B.n803 B.n37 585
R494 B.n37 B.n36 585
R495 B.n802 B.n801 585
R496 B.n801 B.n800 585
R497 B.n39 B.n38 585
R498 B.n799 B.n39 585
R499 B.n842 B.n841 585
R500 B.n841 B.n840 585
R501 B.n699 B.n388 569.379
R502 B.n109 B.n39 569.379
R503 B.n703 B.n390 569.379
R504 B.n797 B.n41 569.379
R505 B.n798 B.n102 256.663
R506 B.n798 B.n101 256.663
R507 B.n798 B.n100 256.663
R508 B.n798 B.n99 256.663
R509 B.n798 B.n98 256.663
R510 B.n798 B.n97 256.663
R511 B.n798 B.n96 256.663
R512 B.n798 B.n95 256.663
R513 B.n798 B.n94 256.663
R514 B.n798 B.n93 256.663
R515 B.n798 B.n92 256.663
R516 B.n798 B.n91 256.663
R517 B.n798 B.n90 256.663
R518 B.n798 B.n89 256.663
R519 B.n798 B.n88 256.663
R520 B.n798 B.n87 256.663
R521 B.n798 B.n86 256.663
R522 B.n798 B.n85 256.663
R523 B.n798 B.n84 256.663
R524 B.n798 B.n83 256.663
R525 B.n798 B.n82 256.663
R526 B.n798 B.n81 256.663
R527 B.n798 B.n80 256.663
R528 B.n798 B.n79 256.663
R529 B.n798 B.n78 256.663
R530 B.n798 B.n77 256.663
R531 B.n798 B.n76 256.663
R532 B.n798 B.n75 256.663
R533 B.n798 B.n74 256.663
R534 B.n798 B.n73 256.663
R535 B.n798 B.n72 256.663
R536 B.n798 B.n71 256.663
R537 B.n798 B.n70 256.663
R538 B.n798 B.n69 256.663
R539 B.n798 B.n68 256.663
R540 B.n798 B.n67 256.663
R541 B.n798 B.n66 256.663
R542 B.n798 B.n65 256.663
R543 B.n798 B.n64 256.663
R544 B.n798 B.n63 256.663
R545 B.n798 B.n62 256.663
R546 B.n798 B.n61 256.663
R547 B.n798 B.n60 256.663
R548 B.n798 B.n59 256.663
R549 B.n798 B.n58 256.663
R550 B.n798 B.n57 256.663
R551 B.n798 B.n56 256.663
R552 B.n798 B.n55 256.663
R553 B.n798 B.n54 256.663
R554 B.n798 B.n53 256.663
R555 B.n798 B.n52 256.663
R556 B.n798 B.n51 256.663
R557 B.n798 B.n50 256.663
R558 B.n798 B.n49 256.663
R559 B.n798 B.n48 256.663
R560 B.n798 B.n47 256.663
R561 B.n798 B.n46 256.663
R562 B.n798 B.n45 256.663
R563 B.n798 B.n44 256.663
R564 B.n798 B.n43 256.663
R565 B.n798 B.n42 256.663
R566 B.n701 B.n700 256.663
R567 B.n701 B.n393 256.663
R568 B.n701 B.n394 256.663
R569 B.n701 B.n395 256.663
R570 B.n701 B.n396 256.663
R571 B.n701 B.n397 256.663
R572 B.n701 B.n398 256.663
R573 B.n701 B.n399 256.663
R574 B.n701 B.n400 256.663
R575 B.n701 B.n401 256.663
R576 B.n701 B.n402 256.663
R577 B.n701 B.n403 256.663
R578 B.n701 B.n404 256.663
R579 B.n701 B.n405 256.663
R580 B.n701 B.n406 256.663
R581 B.n701 B.n407 256.663
R582 B.n701 B.n408 256.663
R583 B.n701 B.n409 256.663
R584 B.n701 B.n410 256.663
R585 B.n701 B.n411 256.663
R586 B.n701 B.n412 256.663
R587 B.n701 B.n413 256.663
R588 B.n701 B.n414 256.663
R589 B.n701 B.n415 256.663
R590 B.n701 B.n416 256.663
R591 B.n701 B.n417 256.663
R592 B.n701 B.n418 256.663
R593 B.n701 B.n419 256.663
R594 B.n701 B.n420 256.663
R595 B.n701 B.n421 256.663
R596 B.n701 B.n422 256.663
R597 B.n701 B.n423 256.663
R598 B.n701 B.n424 256.663
R599 B.n701 B.n425 256.663
R600 B.n701 B.n426 256.663
R601 B.n701 B.n427 256.663
R602 B.n701 B.n428 256.663
R603 B.n701 B.n429 256.663
R604 B.n701 B.n430 256.663
R605 B.n701 B.n431 256.663
R606 B.n701 B.n432 256.663
R607 B.n701 B.n433 256.663
R608 B.n701 B.n434 256.663
R609 B.n701 B.n435 256.663
R610 B.n701 B.n436 256.663
R611 B.n701 B.n437 256.663
R612 B.n701 B.n438 256.663
R613 B.n701 B.n439 256.663
R614 B.n701 B.n440 256.663
R615 B.n701 B.n441 256.663
R616 B.n701 B.n442 256.663
R617 B.n701 B.n443 256.663
R618 B.n701 B.n444 256.663
R619 B.n701 B.n445 256.663
R620 B.n701 B.n446 256.663
R621 B.n701 B.n447 256.663
R622 B.n701 B.n448 256.663
R623 B.n701 B.n449 256.663
R624 B.n701 B.n450 256.663
R625 B.n701 B.n451 256.663
R626 B.n702 B.n701 256.663
R627 B.n709 B.n388 163.367
R628 B.n709 B.n386 163.367
R629 B.n713 B.n386 163.367
R630 B.n713 B.n380 163.367
R631 B.n721 B.n380 163.367
R632 B.n721 B.n378 163.367
R633 B.n725 B.n378 163.367
R634 B.n725 B.n372 163.367
R635 B.n734 B.n372 163.367
R636 B.n734 B.n370 163.367
R637 B.n738 B.n370 163.367
R638 B.n738 B.n365 163.367
R639 B.n746 B.n365 163.367
R640 B.n746 B.n363 163.367
R641 B.n750 B.n363 163.367
R642 B.n750 B.n357 163.367
R643 B.n760 B.n357 163.367
R644 B.n760 B.n355 163.367
R645 B.n764 B.n355 163.367
R646 B.n764 B.n2 163.367
R647 B.n841 B.n2 163.367
R648 B.n841 B.n3 163.367
R649 B.n837 B.n3 163.367
R650 B.n837 B.n8 163.367
R651 B.n833 B.n8 163.367
R652 B.n833 B.n10 163.367
R653 B.n829 B.n10 163.367
R654 B.n829 B.n16 163.367
R655 B.n825 B.n16 163.367
R656 B.n825 B.n18 163.367
R657 B.n821 B.n18 163.367
R658 B.n821 B.n22 163.367
R659 B.n817 B.n22 163.367
R660 B.n817 B.n24 163.367
R661 B.n813 B.n24 163.367
R662 B.n813 B.n30 163.367
R663 B.n809 B.n30 163.367
R664 B.n809 B.n32 163.367
R665 B.n805 B.n32 163.367
R666 B.n805 B.n37 163.367
R667 B.n801 B.n37 163.367
R668 B.n801 B.n39 163.367
R669 B.n453 B.n452 163.367
R670 B.n694 B.n452 163.367
R671 B.n692 B.n691 163.367
R672 B.n688 B.n687 163.367
R673 B.n684 B.n683 163.367
R674 B.n680 B.n679 163.367
R675 B.n676 B.n675 163.367
R676 B.n672 B.n671 163.367
R677 B.n668 B.n667 163.367
R678 B.n664 B.n663 163.367
R679 B.n660 B.n659 163.367
R680 B.n656 B.n655 163.367
R681 B.n652 B.n651 163.367
R682 B.n648 B.n647 163.367
R683 B.n644 B.n643 163.367
R684 B.n640 B.n639 163.367
R685 B.n636 B.n635 163.367
R686 B.n632 B.n631 163.367
R687 B.n628 B.n627 163.367
R688 B.n624 B.n623 163.367
R689 B.n620 B.n619 163.367
R690 B.n616 B.n615 163.367
R691 B.n612 B.n611 163.367
R692 B.n608 B.n607 163.367
R693 B.n604 B.n603 163.367
R694 B.n600 B.n599 163.367
R695 B.n596 B.n595 163.367
R696 B.n592 B.n591 163.367
R697 B.n588 B.n587 163.367
R698 B.n584 B.n583 163.367
R699 B.n580 B.n579 163.367
R700 B.n576 B.n575 163.367
R701 B.n572 B.n571 163.367
R702 B.n567 B.n566 163.367
R703 B.n563 B.n562 163.367
R704 B.n559 B.n558 163.367
R705 B.n555 B.n554 163.367
R706 B.n551 B.n550 163.367
R707 B.n547 B.n546 163.367
R708 B.n543 B.n542 163.367
R709 B.n539 B.n538 163.367
R710 B.n535 B.n534 163.367
R711 B.n531 B.n530 163.367
R712 B.n527 B.n526 163.367
R713 B.n523 B.n522 163.367
R714 B.n519 B.n518 163.367
R715 B.n515 B.n514 163.367
R716 B.n511 B.n510 163.367
R717 B.n507 B.n506 163.367
R718 B.n503 B.n502 163.367
R719 B.n499 B.n498 163.367
R720 B.n495 B.n494 163.367
R721 B.n491 B.n490 163.367
R722 B.n487 B.n486 163.367
R723 B.n483 B.n482 163.367
R724 B.n479 B.n478 163.367
R725 B.n475 B.n474 163.367
R726 B.n471 B.n470 163.367
R727 B.n467 B.n466 163.367
R728 B.n463 B.n462 163.367
R729 B.n459 B.n392 163.367
R730 B.n707 B.n390 163.367
R731 B.n707 B.n383 163.367
R732 B.n715 B.n383 163.367
R733 B.n715 B.n381 163.367
R734 B.n719 B.n381 163.367
R735 B.n719 B.n376 163.367
R736 B.n727 B.n376 163.367
R737 B.n727 B.n374 163.367
R738 B.n731 B.n374 163.367
R739 B.n731 B.n368 163.367
R740 B.n740 B.n368 163.367
R741 B.n740 B.n366 163.367
R742 B.n744 B.n366 163.367
R743 B.n744 B.n361 163.367
R744 B.n752 B.n361 163.367
R745 B.n752 B.n359 163.367
R746 B.n757 B.n359 163.367
R747 B.n757 B.n354 163.367
R748 B.n766 B.n354 163.367
R749 B.n767 B.n766 163.367
R750 B.n767 B.n5 163.367
R751 B.n6 B.n5 163.367
R752 B.n7 B.n6 163.367
R753 B.n772 B.n7 163.367
R754 B.n772 B.n12 163.367
R755 B.n13 B.n12 163.367
R756 B.n14 B.n13 163.367
R757 B.n777 B.n14 163.367
R758 B.n777 B.n19 163.367
R759 B.n20 B.n19 163.367
R760 B.n21 B.n20 163.367
R761 B.n782 B.n21 163.367
R762 B.n782 B.n26 163.367
R763 B.n27 B.n26 163.367
R764 B.n28 B.n27 163.367
R765 B.n787 B.n28 163.367
R766 B.n787 B.n33 163.367
R767 B.n34 B.n33 163.367
R768 B.n35 B.n34 163.367
R769 B.n792 B.n35 163.367
R770 B.n792 B.n40 163.367
R771 B.n41 B.n40 163.367
R772 B.n113 B.n112 163.367
R773 B.n117 B.n116 163.367
R774 B.n121 B.n120 163.367
R775 B.n125 B.n124 163.367
R776 B.n129 B.n128 163.367
R777 B.n133 B.n132 163.367
R778 B.n137 B.n136 163.367
R779 B.n141 B.n140 163.367
R780 B.n145 B.n144 163.367
R781 B.n149 B.n148 163.367
R782 B.n153 B.n152 163.367
R783 B.n157 B.n156 163.367
R784 B.n161 B.n160 163.367
R785 B.n165 B.n164 163.367
R786 B.n169 B.n168 163.367
R787 B.n173 B.n172 163.367
R788 B.n177 B.n176 163.367
R789 B.n181 B.n180 163.367
R790 B.n185 B.n184 163.367
R791 B.n189 B.n188 163.367
R792 B.n193 B.n192 163.367
R793 B.n197 B.n196 163.367
R794 B.n201 B.n200 163.367
R795 B.n205 B.n204 163.367
R796 B.n209 B.n208 163.367
R797 B.n213 B.n212 163.367
R798 B.n217 B.n216 163.367
R799 B.n221 B.n220 163.367
R800 B.n226 B.n225 163.367
R801 B.n230 B.n229 163.367
R802 B.n234 B.n233 163.367
R803 B.n238 B.n237 163.367
R804 B.n242 B.n241 163.367
R805 B.n246 B.n245 163.367
R806 B.n250 B.n249 163.367
R807 B.n254 B.n253 163.367
R808 B.n258 B.n257 163.367
R809 B.n262 B.n261 163.367
R810 B.n266 B.n265 163.367
R811 B.n270 B.n269 163.367
R812 B.n274 B.n273 163.367
R813 B.n278 B.n277 163.367
R814 B.n282 B.n281 163.367
R815 B.n286 B.n285 163.367
R816 B.n290 B.n289 163.367
R817 B.n294 B.n293 163.367
R818 B.n298 B.n297 163.367
R819 B.n302 B.n301 163.367
R820 B.n306 B.n305 163.367
R821 B.n310 B.n309 163.367
R822 B.n314 B.n313 163.367
R823 B.n318 B.n317 163.367
R824 B.n322 B.n321 163.367
R825 B.n326 B.n325 163.367
R826 B.n330 B.n329 163.367
R827 B.n334 B.n333 163.367
R828 B.n338 B.n337 163.367
R829 B.n342 B.n341 163.367
R830 B.n346 B.n345 163.367
R831 B.n350 B.n349 163.367
R832 B.n797 B.n103 163.367
R833 B.n457 B.t18 88.6312
R834 B.n104 B.t10 88.6312
R835 B.n454 B.t21 88.6085
R836 B.n107 B.t13 88.6085
R837 B.n700 B.n699 71.676
R838 B.n694 B.n393 71.676
R839 B.n691 B.n394 71.676
R840 B.n687 B.n395 71.676
R841 B.n683 B.n396 71.676
R842 B.n679 B.n397 71.676
R843 B.n675 B.n398 71.676
R844 B.n671 B.n399 71.676
R845 B.n667 B.n400 71.676
R846 B.n663 B.n401 71.676
R847 B.n659 B.n402 71.676
R848 B.n655 B.n403 71.676
R849 B.n651 B.n404 71.676
R850 B.n647 B.n405 71.676
R851 B.n643 B.n406 71.676
R852 B.n639 B.n407 71.676
R853 B.n635 B.n408 71.676
R854 B.n631 B.n409 71.676
R855 B.n627 B.n410 71.676
R856 B.n623 B.n411 71.676
R857 B.n619 B.n412 71.676
R858 B.n615 B.n413 71.676
R859 B.n611 B.n414 71.676
R860 B.n607 B.n415 71.676
R861 B.n603 B.n416 71.676
R862 B.n599 B.n417 71.676
R863 B.n595 B.n418 71.676
R864 B.n591 B.n419 71.676
R865 B.n587 B.n420 71.676
R866 B.n583 B.n421 71.676
R867 B.n579 B.n422 71.676
R868 B.n575 B.n423 71.676
R869 B.n571 B.n424 71.676
R870 B.n566 B.n425 71.676
R871 B.n562 B.n426 71.676
R872 B.n558 B.n427 71.676
R873 B.n554 B.n428 71.676
R874 B.n550 B.n429 71.676
R875 B.n546 B.n430 71.676
R876 B.n542 B.n431 71.676
R877 B.n538 B.n432 71.676
R878 B.n534 B.n433 71.676
R879 B.n530 B.n434 71.676
R880 B.n526 B.n435 71.676
R881 B.n522 B.n436 71.676
R882 B.n518 B.n437 71.676
R883 B.n514 B.n438 71.676
R884 B.n510 B.n439 71.676
R885 B.n506 B.n440 71.676
R886 B.n502 B.n441 71.676
R887 B.n498 B.n442 71.676
R888 B.n494 B.n443 71.676
R889 B.n490 B.n444 71.676
R890 B.n486 B.n445 71.676
R891 B.n482 B.n446 71.676
R892 B.n478 B.n447 71.676
R893 B.n474 B.n448 71.676
R894 B.n470 B.n449 71.676
R895 B.n466 B.n450 71.676
R896 B.n462 B.n451 71.676
R897 B.n702 B.n392 71.676
R898 B.n109 B.n42 71.676
R899 B.n113 B.n43 71.676
R900 B.n117 B.n44 71.676
R901 B.n121 B.n45 71.676
R902 B.n125 B.n46 71.676
R903 B.n129 B.n47 71.676
R904 B.n133 B.n48 71.676
R905 B.n137 B.n49 71.676
R906 B.n141 B.n50 71.676
R907 B.n145 B.n51 71.676
R908 B.n149 B.n52 71.676
R909 B.n153 B.n53 71.676
R910 B.n157 B.n54 71.676
R911 B.n161 B.n55 71.676
R912 B.n165 B.n56 71.676
R913 B.n169 B.n57 71.676
R914 B.n173 B.n58 71.676
R915 B.n177 B.n59 71.676
R916 B.n181 B.n60 71.676
R917 B.n185 B.n61 71.676
R918 B.n189 B.n62 71.676
R919 B.n193 B.n63 71.676
R920 B.n197 B.n64 71.676
R921 B.n201 B.n65 71.676
R922 B.n205 B.n66 71.676
R923 B.n209 B.n67 71.676
R924 B.n213 B.n68 71.676
R925 B.n217 B.n69 71.676
R926 B.n221 B.n70 71.676
R927 B.n226 B.n71 71.676
R928 B.n230 B.n72 71.676
R929 B.n234 B.n73 71.676
R930 B.n238 B.n74 71.676
R931 B.n242 B.n75 71.676
R932 B.n246 B.n76 71.676
R933 B.n250 B.n77 71.676
R934 B.n254 B.n78 71.676
R935 B.n258 B.n79 71.676
R936 B.n262 B.n80 71.676
R937 B.n266 B.n81 71.676
R938 B.n270 B.n82 71.676
R939 B.n274 B.n83 71.676
R940 B.n278 B.n84 71.676
R941 B.n282 B.n85 71.676
R942 B.n286 B.n86 71.676
R943 B.n290 B.n87 71.676
R944 B.n294 B.n88 71.676
R945 B.n298 B.n89 71.676
R946 B.n302 B.n90 71.676
R947 B.n306 B.n91 71.676
R948 B.n310 B.n92 71.676
R949 B.n314 B.n93 71.676
R950 B.n318 B.n94 71.676
R951 B.n322 B.n95 71.676
R952 B.n326 B.n96 71.676
R953 B.n330 B.n97 71.676
R954 B.n334 B.n98 71.676
R955 B.n338 B.n99 71.676
R956 B.n342 B.n100 71.676
R957 B.n346 B.n101 71.676
R958 B.n350 B.n102 71.676
R959 B.n103 B.n102 71.676
R960 B.n349 B.n101 71.676
R961 B.n345 B.n100 71.676
R962 B.n341 B.n99 71.676
R963 B.n337 B.n98 71.676
R964 B.n333 B.n97 71.676
R965 B.n329 B.n96 71.676
R966 B.n325 B.n95 71.676
R967 B.n321 B.n94 71.676
R968 B.n317 B.n93 71.676
R969 B.n313 B.n92 71.676
R970 B.n309 B.n91 71.676
R971 B.n305 B.n90 71.676
R972 B.n301 B.n89 71.676
R973 B.n297 B.n88 71.676
R974 B.n293 B.n87 71.676
R975 B.n289 B.n86 71.676
R976 B.n285 B.n85 71.676
R977 B.n281 B.n84 71.676
R978 B.n277 B.n83 71.676
R979 B.n273 B.n82 71.676
R980 B.n269 B.n81 71.676
R981 B.n265 B.n80 71.676
R982 B.n261 B.n79 71.676
R983 B.n257 B.n78 71.676
R984 B.n253 B.n77 71.676
R985 B.n249 B.n76 71.676
R986 B.n245 B.n75 71.676
R987 B.n241 B.n74 71.676
R988 B.n237 B.n73 71.676
R989 B.n233 B.n72 71.676
R990 B.n229 B.n71 71.676
R991 B.n225 B.n70 71.676
R992 B.n220 B.n69 71.676
R993 B.n216 B.n68 71.676
R994 B.n212 B.n67 71.676
R995 B.n208 B.n66 71.676
R996 B.n204 B.n65 71.676
R997 B.n200 B.n64 71.676
R998 B.n196 B.n63 71.676
R999 B.n192 B.n62 71.676
R1000 B.n188 B.n61 71.676
R1001 B.n184 B.n60 71.676
R1002 B.n180 B.n59 71.676
R1003 B.n176 B.n58 71.676
R1004 B.n172 B.n57 71.676
R1005 B.n168 B.n56 71.676
R1006 B.n164 B.n55 71.676
R1007 B.n160 B.n54 71.676
R1008 B.n156 B.n53 71.676
R1009 B.n152 B.n52 71.676
R1010 B.n148 B.n51 71.676
R1011 B.n144 B.n50 71.676
R1012 B.n140 B.n49 71.676
R1013 B.n136 B.n48 71.676
R1014 B.n132 B.n47 71.676
R1015 B.n128 B.n46 71.676
R1016 B.n124 B.n45 71.676
R1017 B.n120 B.n44 71.676
R1018 B.n116 B.n43 71.676
R1019 B.n112 B.n42 71.676
R1020 B.n700 B.n453 71.676
R1021 B.n692 B.n393 71.676
R1022 B.n688 B.n394 71.676
R1023 B.n684 B.n395 71.676
R1024 B.n680 B.n396 71.676
R1025 B.n676 B.n397 71.676
R1026 B.n672 B.n398 71.676
R1027 B.n668 B.n399 71.676
R1028 B.n664 B.n400 71.676
R1029 B.n660 B.n401 71.676
R1030 B.n656 B.n402 71.676
R1031 B.n652 B.n403 71.676
R1032 B.n648 B.n404 71.676
R1033 B.n644 B.n405 71.676
R1034 B.n640 B.n406 71.676
R1035 B.n636 B.n407 71.676
R1036 B.n632 B.n408 71.676
R1037 B.n628 B.n409 71.676
R1038 B.n624 B.n410 71.676
R1039 B.n620 B.n411 71.676
R1040 B.n616 B.n412 71.676
R1041 B.n612 B.n413 71.676
R1042 B.n608 B.n414 71.676
R1043 B.n604 B.n415 71.676
R1044 B.n600 B.n416 71.676
R1045 B.n596 B.n417 71.676
R1046 B.n592 B.n418 71.676
R1047 B.n588 B.n419 71.676
R1048 B.n584 B.n420 71.676
R1049 B.n580 B.n421 71.676
R1050 B.n576 B.n422 71.676
R1051 B.n572 B.n423 71.676
R1052 B.n567 B.n424 71.676
R1053 B.n563 B.n425 71.676
R1054 B.n559 B.n426 71.676
R1055 B.n555 B.n427 71.676
R1056 B.n551 B.n428 71.676
R1057 B.n547 B.n429 71.676
R1058 B.n543 B.n430 71.676
R1059 B.n539 B.n431 71.676
R1060 B.n535 B.n432 71.676
R1061 B.n531 B.n433 71.676
R1062 B.n527 B.n434 71.676
R1063 B.n523 B.n435 71.676
R1064 B.n519 B.n436 71.676
R1065 B.n515 B.n437 71.676
R1066 B.n511 B.n438 71.676
R1067 B.n507 B.n439 71.676
R1068 B.n503 B.n440 71.676
R1069 B.n499 B.n441 71.676
R1070 B.n495 B.n442 71.676
R1071 B.n491 B.n443 71.676
R1072 B.n487 B.n444 71.676
R1073 B.n483 B.n445 71.676
R1074 B.n479 B.n446 71.676
R1075 B.n475 B.n447 71.676
R1076 B.n471 B.n448 71.676
R1077 B.n467 B.n449 71.676
R1078 B.n463 B.n450 71.676
R1079 B.n459 B.n451 71.676
R1080 B.n703 B.n702 71.676
R1081 B.n458 B.t17 71.3706
R1082 B.n105 B.t11 71.3706
R1083 B.n455 B.t20 71.3479
R1084 B.n108 B.t14 71.3479
R1085 B.n701 B.n389 67.023
R1086 B.n799 B.n798 67.023
R1087 B.n569 B.n458 59.5399
R1088 B.n456 B.n455 59.5399
R1089 B.n223 B.n108 59.5399
R1090 B.n106 B.n105 59.5399
R1091 B.n110 B.n38 36.9956
R1092 B.n796 B.n795 36.9956
R1093 B.n705 B.n704 36.9956
R1094 B.n698 B.n387 36.9956
R1095 B.n708 B.n389 33.2671
R1096 B.n708 B.n384 33.2671
R1097 B.n714 B.n384 33.2671
R1098 B.n714 B.n385 33.2671
R1099 B.n720 B.n377 33.2671
R1100 B.n726 B.n377 33.2671
R1101 B.n726 B.n373 33.2671
R1102 B.n733 B.n373 33.2671
R1103 B.n733 B.n732 33.2671
R1104 B.n739 B.n369 33.2671
R1105 B.n745 B.n362 33.2671
R1106 B.n751 B.n362 33.2671
R1107 B.n759 B.n358 33.2671
R1108 B.n759 B.n758 33.2671
R1109 B.n765 B.n4 33.2671
R1110 B.n840 B.n4 33.2671
R1111 B.n840 B.n839 33.2671
R1112 B.n839 B.n838 33.2671
R1113 B.n832 B.n11 33.2671
R1114 B.n832 B.n831 33.2671
R1115 B.n830 B.n15 33.2671
R1116 B.n824 B.n15 33.2671
R1117 B.n823 B.n822 33.2671
R1118 B.n816 B.n25 33.2671
R1119 B.n816 B.n815 33.2671
R1120 B.n815 B.n814 33.2671
R1121 B.n814 B.n29 33.2671
R1122 B.n808 B.n29 33.2671
R1123 B.n807 B.n806 33.2671
R1124 B.n806 B.n36 33.2671
R1125 B.n800 B.n36 33.2671
R1126 B.n800 B.n799 33.2671
R1127 B.n765 B.t2 30.3318
R1128 B.n838 B.t3 30.3318
R1129 B.n369 B.t0 28.375
R1130 B.t1 B.n823 28.375
R1131 B.n739 B.t6 25.4397
R1132 B.n822 B.t7 25.4397
R1133 B.n720 B.t16 19.5691
R1134 B.n808 B.t9 19.5691
R1135 B B.n842 18.0485
R1136 B.t5 B.n358 17.6122
R1137 B.n831 B.t4 17.6122
R1138 B.n458 B.n457 17.2611
R1139 B.n455 B.n454 17.2611
R1140 B.n108 B.n107 17.2611
R1141 B.n105 B.n104 17.2611
R1142 B.n751 B.t5 15.6554
R1143 B.t4 B.n830 15.6554
R1144 B.n385 B.t16 13.6985
R1145 B.t9 B.n807 13.6985
R1146 B.n111 B.n110 10.6151
R1147 B.n114 B.n111 10.6151
R1148 B.n115 B.n114 10.6151
R1149 B.n118 B.n115 10.6151
R1150 B.n119 B.n118 10.6151
R1151 B.n122 B.n119 10.6151
R1152 B.n123 B.n122 10.6151
R1153 B.n126 B.n123 10.6151
R1154 B.n127 B.n126 10.6151
R1155 B.n130 B.n127 10.6151
R1156 B.n131 B.n130 10.6151
R1157 B.n134 B.n131 10.6151
R1158 B.n135 B.n134 10.6151
R1159 B.n138 B.n135 10.6151
R1160 B.n139 B.n138 10.6151
R1161 B.n142 B.n139 10.6151
R1162 B.n143 B.n142 10.6151
R1163 B.n146 B.n143 10.6151
R1164 B.n147 B.n146 10.6151
R1165 B.n150 B.n147 10.6151
R1166 B.n151 B.n150 10.6151
R1167 B.n154 B.n151 10.6151
R1168 B.n155 B.n154 10.6151
R1169 B.n158 B.n155 10.6151
R1170 B.n159 B.n158 10.6151
R1171 B.n162 B.n159 10.6151
R1172 B.n163 B.n162 10.6151
R1173 B.n166 B.n163 10.6151
R1174 B.n167 B.n166 10.6151
R1175 B.n170 B.n167 10.6151
R1176 B.n171 B.n170 10.6151
R1177 B.n174 B.n171 10.6151
R1178 B.n175 B.n174 10.6151
R1179 B.n178 B.n175 10.6151
R1180 B.n179 B.n178 10.6151
R1181 B.n182 B.n179 10.6151
R1182 B.n183 B.n182 10.6151
R1183 B.n186 B.n183 10.6151
R1184 B.n187 B.n186 10.6151
R1185 B.n190 B.n187 10.6151
R1186 B.n191 B.n190 10.6151
R1187 B.n194 B.n191 10.6151
R1188 B.n195 B.n194 10.6151
R1189 B.n198 B.n195 10.6151
R1190 B.n199 B.n198 10.6151
R1191 B.n202 B.n199 10.6151
R1192 B.n203 B.n202 10.6151
R1193 B.n206 B.n203 10.6151
R1194 B.n207 B.n206 10.6151
R1195 B.n210 B.n207 10.6151
R1196 B.n211 B.n210 10.6151
R1197 B.n214 B.n211 10.6151
R1198 B.n215 B.n214 10.6151
R1199 B.n218 B.n215 10.6151
R1200 B.n219 B.n218 10.6151
R1201 B.n222 B.n219 10.6151
R1202 B.n227 B.n224 10.6151
R1203 B.n228 B.n227 10.6151
R1204 B.n231 B.n228 10.6151
R1205 B.n232 B.n231 10.6151
R1206 B.n235 B.n232 10.6151
R1207 B.n236 B.n235 10.6151
R1208 B.n239 B.n236 10.6151
R1209 B.n240 B.n239 10.6151
R1210 B.n244 B.n243 10.6151
R1211 B.n247 B.n244 10.6151
R1212 B.n248 B.n247 10.6151
R1213 B.n251 B.n248 10.6151
R1214 B.n252 B.n251 10.6151
R1215 B.n255 B.n252 10.6151
R1216 B.n256 B.n255 10.6151
R1217 B.n259 B.n256 10.6151
R1218 B.n260 B.n259 10.6151
R1219 B.n263 B.n260 10.6151
R1220 B.n264 B.n263 10.6151
R1221 B.n267 B.n264 10.6151
R1222 B.n268 B.n267 10.6151
R1223 B.n271 B.n268 10.6151
R1224 B.n272 B.n271 10.6151
R1225 B.n275 B.n272 10.6151
R1226 B.n276 B.n275 10.6151
R1227 B.n279 B.n276 10.6151
R1228 B.n280 B.n279 10.6151
R1229 B.n283 B.n280 10.6151
R1230 B.n284 B.n283 10.6151
R1231 B.n287 B.n284 10.6151
R1232 B.n288 B.n287 10.6151
R1233 B.n291 B.n288 10.6151
R1234 B.n292 B.n291 10.6151
R1235 B.n295 B.n292 10.6151
R1236 B.n296 B.n295 10.6151
R1237 B.n299 B.n296 10.6151
R1238 B.n300 B.n299 10.6151
R1239 B.n303 B.n300 10.6151
R1240 B.n304 B.n303 10.6151
R1241 B.n307 B.n304 10.6151
R1242 B.n308 B.n307 10.6151
R1243 B.n311 B.n308 10.6151
R1244 B.n312 B.n311 10.6151
R1245 B.n315 B.n312 10.6151
R1246 B.n316 B.n315 10.6151
R1247 B.n319 B.n316 10.6151
R1248 B.n320 B.n319 10.6151
R1249 B.n323 B.n320 10.6151
R1250 B.n324 B.n323 10.6151
R1251 B.n327 B.n324 10.6151
R1252 B.n328 B.n327 10.6151
R1253 B.n331 B.n328 10.6151
R1254 B.n332 B.n331 10.6151
R1255 B.n335 B.n332 10.6151
R1256 B.n336 B.n335 10.6151
R1257 B.n339 B.n336 10.6151
R1258 B.n340 B.n339 10.6151
R1259 B.n343 B.n340 10.6151
R1260 B.n344 B.n343 10.6151
R1261 B.n347 B.n344 10.6151
R1262 B.n348 B.n347 10.6151
R1263 B.n351 B.n348 10.6151
R1264 B.n352 B.n351 10.6151
R1265 B.n796 B.n352 10.6151
R1266 B.n706 B.n705 10.6151
R1267 B.n706 B.n382 10.6151
R1268 B.n716 B.n382 10.6151
R1269 B.n717 B.n716 10.6151
R1270 B.n718 B.n717 10.6151
R1271 B.n718 B.n375 10.6151
R1272 B.n728 B.n375 10.6151
R1273 B.n729 B.n728 10.6151
R1274 B.n730 B.n729 10.6151
R1275 B.n730 B.n367 10.6151
R1276 B.n741 B.n367 10.6151
R1277 B.n742 B.n741 10.6151
R1278 B.n743 B.n742 10.6151
R1279 B.n743 B.n360 10.6151
R1280 B.n753 B.n360 10.6151
R1281 B.n754 B.n753 10.6151
R1282 B.n756 B.n754 10.6151
R1283 B.n756 B.n755 10.6151
R1284 B.n755 B.n353 10.6151
R1285 B.n768 B.n353 10.6151
R1286 B.n769 B.n768 10.6151
R1287 B.n770 B.n769 10.6151
R1288 B.n771 B.n770 10.6151
R1289 B.n773 B.n771 10.6151
R1290 B.n774 B.n773 10.6151
R1291 B.n775 B.n774 10.6151
R1292 B.n776 B.n775 10.6151
R1293 B.n778 B.n776 10.6151
R1294 B.n779 B.n778 10.6151
R1295 B.n780 B.n779 10.6151
R1296 B.n781 B.n780 10.6151
R1297 B.n783 B.n781 10.6151
R1298 B.n784 B.n783 10.6151
R1299 B.n785 B.n784 10.6151
R1300 B.n786 B.n785 10.6151
R1301 B.n788 B.n786 10.6151
R1302 B.n789 B.n788 10.6151
R1303 B.n790 B.n789 10.6151
R1304 B.n791 B.n790 10.6151
R1305 B.n793 B.n791 10.6151
R1306 B.n794 B.n793 10.6151
R1307 B.n795 B.n794 10.6151
R1308 B.n698 B.n697 10.6151
R1309 B.n697 B.n696 10.6151
R1310 B.n696 B.n695 10.6151
R1311 B.n695 B.n693 10.6151
R1312 B.n693 B.n690 10.6151
R1313 B.n690 B.n689 10.6151
R1314 B.n689 B.n686 10.6151
R1315 B.n686 B.n685 10.6151
R1316 B.n685 B.n682 10.6151
R1317 B.n682 B.n681 10.6151
R1318 B.n681 B.n678 10.6151
R1319 B.n678 B.n677 10.6151
R1320 B.n677 B.n674 10.6151
R1321 B.n674 B.n673 10.6151
R1322 B.n673 B.n670 10.6151
R1323 B.n670 B.n669 10.6151
R1324 B.n669 B.n666 10.6151
R1325 B.n666 B.n665 10.6151
R1326 B.n665 B.n662 10.6151
R1327 B.n662 B.n661 10.6151
R1328 B.n661 B.n658 10.6151
R1329 B.n658 B.n657 10.6151
R1330 B.n657 B.n654 10.6151
R1331 B.n654 B.n653 10.6151
R1332 B.n653 B.n650 10.6151
R1333 B.n650 B.n649 10.6151
R1334 B.n649 B.n646 10.6151
R1335 B.n646 B.n645 10.6151
R1336 B.n645 B.n642 10.6151
R1337 B.n642 B.n641 10.6151
R1338 B.n641 B.n638 10.6151
R1339 B.n638 B.n637 10.6151
R1340 B.n637 B.n634 10.6151
R1341 B.n634 B.n633 10.6151
R1342 B.n633 B.n630 10.6151
R1343 B.n630 B.n629 10.6151
R1344 B.n629 B.n626 10.6151
R1345 B.n626 B.n625 10.6151
R1346 B.n625 B.n622 10.6151
R1347 B.n622 B.n621 10.6151
R1348 B.n621 B.n618 10.6151
R1349 B.n618 B.n617 10.6151
R1350 B.n617 B.n614 10.6151
R1351 B.n614 B.n613 10.6151
R1352 B.n613 B.n610 10.6151
R1353 B.n610 B.n609 10.6151
R1354 B.n609 B.n606 10.6151
R1355 B.n606 B.n605 10.6151
R1356 B.n605 B.n602 10.6151
R1357 B.n602 B.n601 10.6151
R1358 B.n601 B.n598 10.6151
R1359 B.n598 B.n597 10.6151
R1360 B.n597 B.n594 10.6151
R1361 B.n594 B.n593 10.6151
R1362 B.n593 B.n590 10.6151
R1363 B.n590 B.n589 10.6151
R1364 B.n586 B.n585 10.6151
R1365 B.n585 B.n582 10.6151
R1366 B.n582 B.n581 10.6151
R1367 B.n581 B.n578 10.6151
R1368 B.n578 B.n577 10.6151
R1369 B.n577 B.n574 10.6151
R1370 B.n574 B.n573 10.6151
R1371 B.n573 B.n570 10.6151
R1372 B.n568 B.n565 10.6151
R1373 B.n565 B.n564 10.6151
R1374 B.n564 B.n561 10.6151
R1375 B.n561 B.n560 10.6151
R1376 B.n560 B.n557 10.6151
R1377 B.n557 B.n556 10.6151
R1378 B.n556 B.n553 10.6151
R1379 B.n553 B.n552 10.6151
R1380 B.n552 B.n549 10.6151
R1381 B.n549 B.n548 10.6151
R1382 B.n548 B.n545 10.6151
R1383 B.n545 B.n544 10.6151
R1384 B.n544 B.n541 10.6151
R1385 B.n541 B.n540 10.6151
R1386 B.n540 B.n537 10.6151
R1387 B.n537 B.n536 10.6151
R1388 B.n536 B.n533 10.6151
R1389 B.n533 B.n532 10.6151
R1390 B.n532 B.n529 10.6151
R1391 B.n529 B.n528 10.6151
R1392 B.n528 B.n525 10.6151
R1393 B.n525 B.n524 10.6151
R1394 B.n524 B.n521 10.6151
R1395 B.n521 B.n520 10.6151
R1396 B.n520 B.n517 10.6151
R1397 B.n517 B.n516 10.6151
R1398 B.n516 B.n513 10.6151
R1399 B.n513 B.n512 10.6151
R1400 B.n512 B.n509 10.6151
R1401 B.n509 B.n508 10.6151
R1402 B.n508 B.n505 10.6151
R1403 B.n505 B.n504 10.6151
R1404 B.n504 B.n501 10.6151
R1405 B.n501 B.n500 10.6151
R1406 B.n500 B.n497 10.6151
R1407 B.n497 B.n496 10.6151
R1408 B.n496 B.n493 10.6151
R1409 B.n493 B.n492 10.6151
R1410 B.n492 B.n489 10.6151
R1411 B.n489 B.n488 10.6151
R1412 B.n488 B.n485 10.6151
R1413 B.n485 B.n484 10.6151
R1414 B.n484 B.n481 10.6151
R1415 B.n481 B.n480 10.6151
R1416 B.n480 B.n477 10.6151
R1417 B.n477 B.n476 10.6151
R1418 B.n476 B.n473 10.6151
R1419 B.n473 B.n472 10.6151
R1420 B.n472 B.n469 10.6151
R1421 B.n469 B.n468 10.6151
R1422 B.n468 B.n465 10.6151
R1423 B.n465 B.n464 10.6151
R1424 B.n464 B.n461 10.6151
R1425 B.n461 B.n460 10.6151
R1426 B.n460 B.n391 10.6151
R1427 B.n704 B.n391 10.6151
R1428 B.n710 B.n387 10.6151
R1429 B.n711 B.n710 10.6151
R1430 B.n712 B.n711 10.6151
R1431 B.n712 B.n379 10.6151
R1432 B.n722 B.n379 10.6151
R1433 B.n723 B.n722 10.6151
R1434 B.n724 B.n723 10.6151
R1435 B.n724 B.n371 10.6151
R1436 B.n735 B.n371 10.6151
R1437 B.n736 B.n735 10.6151
R1438 B.n737 B.n736 10.6151
R1439 B.n737 B.n364 10.6151
R1440 B.n747 B.n364 10.6151
R1441 B.n748 B.n747 10.6151
R1442 B.n749 B.n748 10.6151
R1443 B.n749 B.n356 10.6151
R1444 B.n761 B.n356 10.6151
R1445 B.n762 B.n761 10.6151
R1446 B.n763 B.n762 10.6151
R1447 B.n763 B.n0 10.6151
R1448 B.n836 B.n1 10.6151
R1449 B.n836 B.n835 10.6151
R1450 B.n835 B.n834 10.6151
R1451 B.n834 B.n9 10.6151
R1452 B.n828 B.n9 10.6151
R1453 B.n828 B.n827 10.6151
R1454 B.n827 B.n826 10.6151
R1455 B.n826 B.n17 10.6151
R1456 B.n820 B.n17 10.6151
R1457 B.n820 B.n819 10.6151
R1458 B.n819 B.n818 10.6151
R1459 B.n818 B.n23 10.6151
R1460 B.n812 B.n23 10.6151
R1461 B.n812 B.n811 10.6151
R1462 B.n811 B.n810 10.6151
R1463 B.n810 B.n31 10.6151
R1464 B.n804 B.n31 10.6151
R1465 B.n804 B.n803 10.6151
R1466 B.n803 B.n802 10.6151
R1467 B.n802 B.n38 10.6151
R1468 B.n732 B.t6 7.82794
R1469 B.n25 B.t7 7.82794
R1470 B.n224 B.n223 6.5566
R1471 B.n240 B.n106 6.5566
R1472 B.n586 B.n456 6.5566
R1473 B.n570 B.n569 6.5566
R1474 B.n745 B.t0 4.89265
R1475 B.n824 B.t1 4.89265
R1476 B.n223 B.n222 4.05904
R1477 B.n243 B.n106 4.05904
R1478 B.n589 B.n456 4.05904
R1479 B.n569 B.n568 4.05904
R1480 B.n758 B.t2 2.93579
R1481 B.n11 B.t3 2.93579
R1482 B.n842 B.n0 2.81026
R1483 B.n842 B.n1 2.81026
R1484 VP.n4 VP.t1 837.266
R1485 VP.n11 VP.t3 811.223
R1486 VP.n1 VP.t5 811.223
R1487 VP.n16 VP.t7 811.223
R1488 VP.n18 VP.t0 811.223
R1489 VP.n8 VP.t4 811.223
R1490 VP.n6 VP.t2 811.223
R1491 VP.n5 VP.t6 811.223
R1492 VP.n19 VP.n18 161.3
R1493 VP.n6 VP.n3 161.3
R1494 VP.n7 VP.n2 161.3
R1495 VP.n9 VP.n8 161.3
R1496 VP.n17 VP.n0 161.3
R1497 VP.n16 VP.n15 161.3
R1498 VP.n14 VP.n1 161.3
R1499 VP.n13 VP.n12 161.3
R1500 VP.n11 VP.n10 161.3
R1501 VP.n16 VP.n1 48.2005
R1502 VP.n6 VP.n5 48.2005
R1503 VP.n10 VP.n9 45.2808
R1504 VP.n4 VP.n3 45.057
R1505 VP.n12 VP.n11 44.549
R1506 VP.n18 VP.n17 44.549
R1507 VP.n8 VP.n7 44.549
R1508 VP.n5 VP.n4 14.6494
R1509 VP.n12 VP.n1 3.65202
R1510 VP.n17 VP.n16 3.65202
R1511 VP.n7 VP.n6 3.65202
R1512 VP.n3 VP.n2 0.189894
R1513 VP.n9 VP.n2 0.189894
R1514 VP.n13 VP.n10 0.189894
R1515 VP.n14 VP.n13 0.189894
R1516 VP.n15 VP.n14 0.189894
R1517 VP.n15 VP.n0 0.189894
R1518 VP.n19 VP.n0 0.189894
R1519 VP VP.n19 0.0516364
R1520 VDD1 VDD1.n0 62.1136
R1521 VDD1.n3 VDD1.n2 61.9998
R1522 VDD1.n3 VDD1.n1 61.9998
R1523 VDD1.n5 VDD1.n4 61.6716
R1524 VDD1.n5 VDD1.n3 42.5871
R1525 VDD1.n4 VDD1.t5 1.15099
R1526 VDD1.n4 VDD1.t3 1.15099
R1527 VDD1.n0 VDD1.t6 1.15099
R1528 VDD1.n0 VDD1.t1 1.15099
R1529 VDD1.n2 VDD1.t0 1.15099
R1530 VDD1.n2 VDD1.t7 1.15099
R1531 VDD1.n1 VDD1.t4 1.15099
R1532 VDD1.n1 VDD1.t2 1.15099
R1533 VDD1 VDD1.n5 0.325931
C0 VN VP 6.13453f
C1 VTAIL VDD1 16.728498f
C2 VDD2 VDD1 0.756909f
C3 VTAIL VN 6.33615f
C4 VN VDD2 6.84135f
C5 VTAIL VP 6.35026f
C6 VDD2 VP 0.302526f
C7 VN VDD1 0.147972f
C8 VTAIL VDD2 16.7692f
C9 VP VDD1 6.99553f
C10 VDD2 B 3.768894f
C11 VDD1 B 3.988896f
C12 VTAIL B 11.688535f
C13 VN B 8.757951f
C14 VP B 6.436725f
C15 VDD1.t6 B 0.391002f
C16 VDD1.t1 B 0.391002f
C17 VDD1.n0 B 3.55927f
C18 VDD1.t4 B 0.391002f
C19 VDD1.t2 B 0.391002f
C20 VDD1.n1 B 3.55856f
C21 VDD1.t0 B 0.391002f
C22 VDD1.t7 B 0.391002f
C23 VDD1.n2 B 3.55856f
C24 VDD1.n3 B 2.83644f
C25 VDD1.t5 B 0.391002f
C26 VDD1.t3 B 0.391002f
C27 VDD1.n4 B 3.55669f
C28 VDD1.n5 B 3.07346f
C29 VP.n0 B 0.047853f
C30 VP.t5 B 1.30849f
C31 VP.n1 B 0.499995f
C32 VP.n2 B 0.047853f
C33 VP.t4 B 1.30849f
C34 VP.t2 B 1.30849f
C35 VP.n3 B 0.197231f
C36 VP.t6 B 1.30849f
C37 VP.t1 B 1.32401f
C38 VP.n4 B 0.485673f
C39 VP.n5 B 0.509146f
C40 VP.n6 B 0.499995f
C41 VP.n7 B 0.010859f
C42 VP.n8 B 0.49852f
C43 VP.n9 B 2.23225f
C44 VP.n10 B 2.27024f
C45 VP.t3 B 1.30849f
C46 VP.n11 B 0.49852f
C47 VP.n12 B 0.010859f
C48 VP.n13 B 0.047853f
C49 VP.n14 B 0.047853f
C50 VP.n15 B 0.047853f
C51 VP.t7 B 1.30849f
C52 VP.n16 B 0.499995f
C53 VP.n17 B 0.010859f
C54 VP.t0 B 1.30849f
C55 VP.n18 B 0.49852f
C56 VP.n19 B 0.037084f
C57 VDD2.t3 B 0.391104f
C58 VDD2.t4 B 0.391104f
C59 VDD2.n0 B 3.5595f
C60 VDD2.t2 B 0.391104f
C61 VDD2.t7 B 0.391104f
C62 VDD2.n1 B 3.5595f
C63 VDD2.n2 B 2.77606f
C64 VDD2.t6 B 0.391104f
C65 VDD2.t1 B 0.391104f
C66 VDD2.n3 B 3.55764f
C67 VDD2.n4 B 3.03995f
C68 VDD2.t5 B 0.391104f
C69 VDD2.t0 B 0.391104f
C70 VDD2.n5 B 3.55946f
C71 VTAIL.t5 B 0.276344f
C72 VTAIL.t6 B 0.276344f
C73 VTAIL.n0 B 2.4531f
C74 VTAIL.n1 B 0.25449f
C75 VTAIL.t4 B 3.13369f
C76 VTAIL.n2 B 0.354515f
C77 VTAIL.t15 B 3.13369f
C78 VTAIL.n3 B 0.354515f
C79 VTAIL.t0 B 0.276344f
C80 VTAIL.t11 B 0.276344f
C81 VTAIL.n4 B 2.4531f
C82 VTAIL.n5 B 0.300915f
C83 VTAIL.t14 B 3.13369f
C84 VTAIL.n6 B 1.6214f
C85 VTAIL.t9 B 3.13371f
C86 VTAIL.n7 B 1.62138f
C87 VTAIL.t7 B 0.276344f
C88 VTAIL.t8 B 0.276344f
C89 VTAIL.n8 B 2.4531f
C90 VTAIL.n9 B 0.300911f
C91 VTAIL.t2 B 3.13371f
C92 VTAIL.n10 B 0.354496f
C93 VTAIL.t10 B 3.13371f
C94 VTAIL.n11 B 0.354496f
C95 VTAIL.t12 B 0.276344f
C96 VTAIL.t1 B 0.276344f
C97 VTAIL.n12 B 2.4531f
C98 VTAIL.n13 B 0.300911f
C99 VTAIL.t13 B 3.13369f
C100 VTAIL.n14 B 1.6214f
C101 VTAIL.t3 B 3.13369f
C102 VTAIL.n15 B 1.61759f
C103 VN.n0 B 0.046955f
C104 VN.t3 B 1.28393f
C105 VN.n1 B 0.49959f
C106 VN.t4 B 1.29916f
C107 VN.n2 B 0.476557f
C108 VN.n3 B 0.193529f
C109 VN.t5 B 1.28393f
C110 VN.n4 B 0.490611f
C111 VN.n5 B 0.010655f
C112 VN.t0 B 1.28393f
C113 VN.n6 B 0.489163f
C114 VN.n7 B 0.036388f
C115 VN.n8 B 0.046955f
C116 VN.t2 B 1.28393f
C117 VN.n9 B 0.49959f
C118 VN.t6 B 1.28393f
C119 VN.t7 B 1.29916f
C120 VN.n10 B 0.476557f
C121 VN.n11 B 0.193529f
C122 VN.n12 B 0.490611f
C123 VN.n13 B 0.010655f
C124 VN.t1 B 1.28393f
C125 VN.n14 B 0.489163f
C126 VN.n15 B 2.22104f
.ends

