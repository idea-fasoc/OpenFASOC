* NGSPICE file created from diff_pair_sample_1079.ext - technology: sky130A

.subckt diff_pair_sample_1079 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t3 B.t5 sky130_fd_pr__nfet_01v8 ad=1.0395 pd=6.63 as=2.457 ps=13.38 w=6.3 l=1.51
X1 VTAIL.t7 VP.t1 VDD1.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=1.0395 pd=6.63 as=1.0395 ps=6.63 w=6.3 l=1.51
X2 VDD1.t3 VP.t2 VTAIL.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=2.457 pd=13.38 as=1.0395 ps=6.63 w=6.3 l=1.51
X3 VTAIL.t4 VP.t3 VDD1.t2 B.t4 sky130_fd_pr__nfet_01v8 ad=1.0395 pd=6.63 as=1.0395 ps=6.63 w=6.3 l=1.51
X4 VDD1.t1 VP.t4 VTAIL.t8 B.t0 sky130_fd_pr__nfet_01v8 ad=1.0395 pd=6.63 as=2.457 ps=13.38 w=6.3 l=1.51
X5 B.t19 B.t17 B.t18 B.t11 sky130_fd_pr__nfet_01v8 ad=2.457 pd=13.38 as=0 ps=0 w=6.3 l=1.51
X6 VDD2.t5 VN.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.0395 pd=6.63 as=2.457 ps=13.38 w=6.3 l=1.51
X7 B.t16 B.t14 B.t15 B.t7 sky130_fd_pr__nfet_01v8 ad=2.457 pd=13.38 as=0 ps=0 w=6.3 l=1.51
X8 VDD2.t4 VN.t1 VTAIL.t10 B.t5 sky130_fd_pr__nfet_01v8 ad=1.0395 pd=6.63 as=2.457 ps=13.38 w=6.3 l=1.51
X9 VDD2.t3 VN.t2 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.457 pd=13.38 as=1.0395 ps=6.63 w=6.3 l=1.51
X10 VTAIL.t2 VN.t3 VDD2.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.0395 pd=6.63 as=1.0395 ps=6.63 w=6.3 l=1.51
X11 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=2.457 pd=13.38 as=0 ps=0 w=6.3 l=1.51
X12 VTAIL.t9 VN.t4 VDD2.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=1.0395 pd=6.63 as=1.0395 ps=6.63 w=6.3 l=1.51
X13 VDD2.t0 VN.t5 VTAIL.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=2.457 pd=13.38 as=1.0395 ps=6.63 w=6.3 l=1.51
X14 VDD1.t0 VP.t5 VTAIL.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=2.457 pd=13.38 as=1.0395 ps=6.63 w=6.3 l=1.51
X15 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=2.457 pd=13.38 as=0 ps=0 w=6.3 l=1.51
R0 VP.n17 VP.n16 181.465
R1 VP.n32 VP.n31 181.465
R2 VP.n15 VP.n14 181.465
R3 VP.n9 VP.n8 161.3
R4 VP.n10 VP.n5 161.3
R5 VP.n12 VP.n11 161.3
R6 VP.n13 VP.n4 161.3
R7 VP.n30 VP.n0 161.3
R8 VP.n29 VP.n28 161.3
R9 VP.n27 VP.n1 161.3
R10 VP.n26 VP.n25 161.3
R11 VP.n23 VP.n2 161.3
R12 VP.n22 VP.n21 161.3
R13 VP.n20 VP.n3 161.3
R14 VP.n19 VP.n18 161.3
R15 VP.n6 VP.t5 131.316
R16 VP.n17 VP.t2 100.55
R17 VP.n24 VP.t3 100.55
R18 VP.n31 VP.t4 100.55
R19 VP.n14 VP.t0 100.55
R20 VP.n7 VP.t1 100.55
R21 VP.n22 VP.n3 56.5617
R22 VP.n29 VP.n1 56.5617
R23 VP.n12 VP.n5 56.5617
R24 VP.n7 VP.n6 53.734
R25 VP.n16 VP.n15 39.9247
R26 VP.n18 VP.n3 24.5923
R27 VP.n23 VP.n22 24.5923
R28 VP.n25 VP.n1 24.5923
R29 VP.n30 VP.n29 24.5923
R30 VP.n13 VP.n12 24.5923
R31 VP.n8 VP.n5 24.5923
R32 VP.n9 VP.n6 18.3138
R33 VP.n24 VP.n23 12.2964
R34 VP.n25 VP.n24 12.2964
R35 VP.n8 VP.n7 12.2964
R36 VP.n18 VP.n17 4.42703
R37 VP.n31 VP.n30 4.42703
R38 VP.n14 VP.n13 4.42703
R39 VP.n10 VP.n9 0.189894
R40 VP.n11 VP.n10 0.189894
R41 VP.n11 VP.n4 0.189894
R42 VP.n15 VP.n4 0.189894
R43 VP.n19 VP.n16 0.189894
R44 VP.n20 VP.n19 0.189894
R45 VP.n21 VP.n20 0.189894
R46 VP.n21 VP.n2 0.189894
R47 VP.n26 VP.n2 0.189894
R48 VP.n27 VP.n26 0.189894
R49 VP.n28 VP.n27 0.189894
R50 VP.n28 VP.n0 0.189894
R51 VP.n32 VP.n0 0.189894
R52 VP VP.n32 0.0516364
R53 VTAIL.n7 VTAIL.t0 51.8964
R54 VTAIL.n10 VTAIL.t3 51.8963
R55 VTAIL.n11 VTAIL.t10 51.8963
R56 VTAIL.n2 VTAIL.t8 51.8963
R57 VTAIL.n9 VTAIL.n8 48.7536
R58 VTAIL.n6 VTAIL.n5 48.7536
R59 VTAIL.n1 VTAIL.n0 48.7534
R60 VTAIL.n4 VTAIL.n3 48.7534
R61 VTAIL.n6 VTAIL.n4 20.9703
R62 VTAIL.n11 VTAIL.n10 19.3841
R63 VTAIL.n0 VTAIL.t11 3.14336
R64 VTAIL.n0 VTAIL.t2 3.14336
R65 VTAIL.n3 VTAIL.t5 3.14336
R66 VTAIL.n3 VTAIL.t4 3.14336
R67 VTAIL.n8 VTAIL.t6 3.14336
R68 VTAIL.n8 VTAIL.t7 3.14336
R69 VTAIL.n5 VTAIL.t1 3.14336
R70 VTAIL.n5 VTAIL.t9 3.14336
R71 VTAIL.n7 VTAIL.n6 1.58671
R72 VTAIL.n10 VTAIL.n9 1.58671
R73 VTAIL.n4 VTAIL.n2 1.58671
R74 VTAIL.n9 VTAIL.n7 1.26343
R75 VTAIL.n2 VTAIL.n1 1.26343
R76 VTAIL VTAIL.n11 1.13197
R77 VTAIL VTAIL.n1 0.455241
R78 VDD1 VDD1.t0 69.8231
R79 VDD1.n1 VDD1.t3 69.7094
R80 VDD1.n1 VDD1.n0 65.7734
R81 VDD1.n3 VDD1.n2 65.4322
R82 VDD1.n3 VDD1.n1 35.6776
R83 VDD1.n2 VDD1.t4 3.14336
R84 VDD1.n2 VDD1.t5 3.14336
R85 VDD1.n0 VDD1.t2 3.14336
R86 VDD1.n0 VDD1.t1 3.14336
R87 VDD1 VDD1.n3 0.338862
R88 B.n544 B.n543 585
R89 B.n545 B.n544 585
R90 B.n206 B.n85 585
R91 B.n205 B.n204 585
R92 B.n203 B.n202 585
R93 B.n201 B.n200 585
R94 B.n199 B.n198 585
R95 B.n197 B.n196 585
R96 B.n195 B.n194 585
R97 B.n193 B.n192 585
R98 B.n191 B.n190 585
R99 B.n189 B.n188 585
R100 B.n187 B.n186 585
R101 B.n185 B.n184 585
R102 B.n183 B.n182 585
R103 B.n181 B.n180 585
R104 B.n179 B.n178 585
R105 B.n177 B.n176 585
R106 B.n175 B.n174 585
R107 B.n173 B.n172 585
R108 B.n171 B.n170 585
R109 B.n169 B.n168 585
R110 B.n167 B.n166 585
R111 B.n165 B.n164 585
R112 B.n163 B.n162 585
R113 B.n161 B.n160 585
R114 B.n159 B.n158 585
R115 B.n157 B.n156 585
R116 B.n155 B.n154 585
R117 B.n153 B.n152 585
R118 B.n151 B.n150 585
R119 B.n149 B.n148 585
R120 B.n147 B.n146 585
R121 B.n145 B.n144 585
R122 B.n143 B.n142 585
R123 B.n140 B.n139 585
R124 B.n138 B.n137 585
R125 B.n136 B.n135 585
R126 B.n134 B.n133 585
R127 B.n132 B.n131 585
R128 B.n130 B.n129 585
R129 B.n128 B.n127 585
R130 B.n126 B.n125 585
R131 B.n124 B.n123 585
R132 B.n122 B.n121 585
R133 B.n120 B.n119 585
R134 B.n118 B.n117 585
R135 B.n116 B.n115 585
R136 B.n114 B.n113 585
R137 B.n112 B.n111 585
R138 B.n110 B.n109 585
R139 B.n108 B.n107 585
R140 B.n106 B.n105 585
R141 B.n104 B.n103 585
R142 B.n102 B.n101 585
R143 B.n100 B.n99 585
R144 B.n98 B.n97 585
R145 B.n96 B.n95 585
R146 B.n94 B.n93 585
R147 B.n92 B.n91 585
R148 B.n542 B.n55 585
R149 B.n546 B.n55 585
R150 B.n541 B.n54 585
R151 B.n547 B.n54 585
R152 B.n540 B.n539 585
R153 B.n539 B.n50 585
R154 B.n538 B.n49 585
R155 B.n553 B.n49 585
R156 B.n537 B.n48 585
R157 B.n554 B.n48 585
R158 B.n536 B.n47 585
R159 B.n555 B.n47 585
R160 B.n535 B.n534 585
R161 B.n534 B.n43 585
R162 B.n533 B.n42 585
R163 B.n561 B.n42 585
R164 B.n532 B.n41 585
R165 B.n562 B.n41 585
R166 B.n531 B.n40 585
R167 B.n563 B.n40 585
R168 B.n530 B.n529 585
R169 B.n529 B.n36 585
R170 B.n528 B.n35 585
R171 B.n569 B.n35 585
R172 B.n527 B.n34 585
R173 B.n570 B.n34 585
R174 B.n526 B.n33 585
R175 B.n571 B.n33 585
R176 B.n525 B.n524 585
R177 B.n524 B.n32 585
R178 B.n523 B.n28 585
R179 B.n577 B.n28 585
R180 B.n522 B.n27 585
R181 B.n578 B.n27 585
R182 B.n521 B.n26 585
R183 B.n579 B.n26 585
R184 B.n520 B.n519 585
R185 B.n519 B.n22 585
R186 B.n518 B.n21 585
R187 B.n585 B.n21 585
R188 B.n517 B.n20 585
R189 B.n586 B.n20 585
R190 B.n516 B.n19 585
R191 B.n587 B.n19 585
R192 B.n515 B.n514 585
R193 B.n514 B.n15 585
R194 B.n513 B.n14 585
R195 B.n593 B.n14 585
R196 B.n512 B.n13 585
R197 B.n594 B.n13 585
R198 B.n511 B.n12 585
R199 B.n595 B.n12 585
R200 B.n510 B.n509 585
R201 B.n509 B.n508 585
R202 B.n507 B.n506 585
R203 B.n507 B.n8 585
R204 B.n505 B.n7 585
R205 B.n602 B.n7 585
R206 B.n504 B.n6 585
R207 B.n603 B.n6 585
R208 B.n503 B.n5 585
R209 B.n604 B.n5 585
R210 B.n502 B.n501 585
R211 B.n501 B.n4 585
R212 B.n500 B.n207 585
R213 B.n500 B.n499 585
R214 B.n490 B.n208 585
R215 B.n209 B.n208 585
R216 B.n492 B.n491 585
R217 B.n493 B.n492 585
R218 B.n489 B.n214 585
R219 B.n214 B.n213 585
R220 B.n488 B.n487 585
R221 B.n487 B.n486 585
R222 B.n216 B.n215 585
R223 B.n217 B.n216 585
R224 B.n479 B.n478 585
R225 B.n480 B.n479 585
R226 B.n477 B.n222 585
R227 B.n222 B.n221 585
R228 B.n476 B.n475 585
R229 B.n475 B.n474 585
R230 B.n224 B.n223 585
R231 B.n225 B.n224 585
R232 B.n467 B.n466 585
R233 B.n468 B.n467 585
R234 B.n465 B.n230 585
R235 B.n230 B.n229 585
R236 B.n464 B.n463 585
R237 B.n463 B.n462 585
R238 B.n232 B.n231 585
R239 B.n455 B.n232 585
R240 B.n454 B.n453 585
R241 B.n456 B.n454 585
R242 B.n452 B.n237 585
R243 B.n237 B.n236 585
R244 B.n451 B.n450 585
R245 B.n450 B.n449 585
R246 B.n239 B.n238 585
R247 B.n240 B.n239 585
R248 B.n442 B.n441 585
R249 B.n443 B.n442 585
R250 B.n440 B.n245 585
R251 B.n245 B.n244 585
R252 B.n439 B.n438 585
R253 B.n438 B.n437 585
R254 B.n247 B.n246 585
R255 B.n248 B.n247 585
R256 B.n430 B.n429 585
R257 B.n431 B.n430 585
R258 B.n428 B.n253 585
R259 B.n253 B.n252 585
R260 B.n427 B.n426 585
R261 B.n426 B.n425 585
R262 B.n255 B.n254 585
R263 B.n256 B.n255 585
R264 B.n418 B.n417 585
R265 B.n419 B.n418 585
R266 B.n416 B.n261 585
R267 B.n261 B.n260 585
R268 B.n410 B.n409 585
R269 B.n408 B.n292 585
R270 B.n407 B.n291 585
R271 B.n412 B.n291 585
R272 B.n406 B.n405 585
R273 B.n404 B.n403 585
R274 B.n402 B.n401 585
R275 B.n400 B.n399 585
R276 B.n398 B.n397 585
R277 B.n396 B.n395 585
R278 B.n394 B.n393 585
R279 B.n392 B.n391 585
R280 B.n390 B.n389 585
R281 B.n388 B.n387 585
R282 B.n386 B.n385 585
R283 B.n384 B.n383 585
R284 B.n382 B.n381 585
R285 B.n380 B.n379 585
R286 B.n378 B.n377 585
R287 B.n376 B.n375 585
R288 B.n374 B.n373 585
R289 B.n372 B.n371 585
R290 B.n370 B.n369 585
R291 B.n368 B.n367 585
R292 B.n366 B.n365 585
R293 B.n364 B.n363 585
R294 B.n362 B.n361 585
R295 B.n360 B.n359 585
R296 B.n358 B.n357 585
R297 B.n356 B.n355 585
R298 B.n354 B.n353 585
R299 B.n352 B.n351 585
R300 B.n350 B.n349 585
R301 B.n348 B.n347 585
R302 B.n346 B.n345 585
R303 B.n343 B.n342 585
R304 B.n341 B.n340 585
R305 B.n339 B.n338 585
R306 B.n337 B.n336 585
R307 B.n335 B.n334 585
R308 B.n333 B.n332 585
R309 B.n331 B.n330 585
R310 B.n329 B.n328 585
R311 B.n327 B.n326 585
R312 B.n325 B.n324 585
R313 B.n323 B.n322 585
R314 B.n321 B.n320 585
R315 B.n319 B.n318 585
R316 B.n317 B.n316 585
R317 B.n315 B.n314 585
R318 B.n313 B.n312 585
R319 B.n311 B.n310 585
R320 B.n309 B.n308 585
R321 B.n307 B.n306 585
R322 B.n305 B.n304 585
R323 B.n303 B.n302 585
R324 B.n301 B.n300 585
R325 B.n299 B.n298 585
R326 B.n263 B.n262 585
R327 B.n415 B.n414 585
R328 B.n259 B.n258 585
R329 B.n260 B.n259 585
R330 B.n421 B.n420 585
R331 B.n420 B.n419 585
R332 B.n422 B.n257 585
R333 B.n257 B.n256 585
R334 B.n424 B.n423 585
R335 B.n425 B.n424 585
R336 B.n251 B.n250 585
R337 B.n252 B.n251 585
R338 B.n433 B.n432 585
R339 B.n432 B.n431 585
R340 B.n434 B.n249 585
R341 B.n249 B.n248 585
R342 B.n436 B.n435 585
R343 B.n437 B.n436 585
R344 B.n243 B.n242 585
R345 B.n244 B.n243 585
R346 B.n445 B.n444 585
R347 B.n444 B.n443 585
R348 B.n446 B.n241 585
R349 B.n241 B.n240 585
R350 B.n448 B.n447 585
R351 B.n449 B.n448 585
R352 B.n235 B.n234 585
R353 B.n236 B.n235 585
R354 B.n458 B.n457 585
R355 B.n457 B.n456 585
R356 B.n459 B.n233 585
R357 B.n455 B.n233 585
R358 B.n461 B.n460 585
R359 B.n462 B.n461 585
R360 B.n228 B.n227 585
R361 B.n229 B.n228 585
R362 B.n470 B.n469 585
R363 B.n469 B.n468 585
R364 B.n471 B.n226 585
R365 B.n226 B.n225 585
R366 B.n473 B.n472 585
R367 B.n474 B.n473 585
R368 B.n220 B.n219 585
R369 B.n221 B.n220 585
R370 B.n482 B.n481 585
R371 B.n481 B.n480 585
R372 B.n483 B.n218 585
R373 B.n218 B.n217 585
R374 B.n485 B.n484 585
R375 B.n486 B.n485 585
R376 B.n212 B.n211 585
R377 B.n213 B.n212 585
R378 B.n495 B.n494 585
R379 B.n494 B.n493 585
R380 B.n496 B.n210 585
R381 B.n210 B.n209 585
R382 B.n498 B.n497 585
R383 B.n499 B.n498 585
R384 B.n3 B.n0 585
R385 B.n4 B.n3 585
R386 B.n601 B.n1 585
R387 B.n602 B.n601 585
R388 B.n600 B.n599 585
R389 B.n600 B.n8 585
R390 B.n598 B.n9 585
R391 B.n508 B.n9 585
R392 B.n597 B.n596 585
R393 B.n596 B.n595 585
R394 B.n11 B.n10 585
R395 B.n594 B.n11 585
R396 B.n592 B.n591 585
R397 B.n593 B.n592 585
R398 B.n590 B.n16 585
R399 B.n16 B.n15 585
R400 B.n589 B.n588 585
R401 B.n588 B.n587 585
R402 B.n18 B.n17 585
R403 B.n586 B.n18 585
R404 B.n584 B.n583 585
R405 B.n585 B.n584 585
R406 B.n582 B.n23 585
R407 B.n23 B.n22 585
R408 B.n581 B.n580 585
R409 B.n580 B.n579 585
R410 B.n25 B.n24 585
R411 B.n578 B.n25 585
R412 B.n576 B.n575 585
R413 B.n577 B.n576 585
R414 B.n574 B.n29 585
R415 B.n32 B.n29 585
R416 B.n573 B.n572 585
R417 B.n572 B.n571 585
R418 B.n31 B.n30 585
R419 B.n570 B.n31 585
R420 B.n568 B.n567 585
R421 B.n569 B.n568 585
R422 B.n566 B.n37 585
R423 B.n37 B.n36 585
R424 B.n565 B.n564 585
R425 B.n564 B.n563 585
R426 B.n39 B.n38 585
R427 B.n562 B.n39 585
R428 B.n560 B.n559 585
R429 B.n561 B.n560 585
R430 B.n558 B.n44 585
R431 B.n44 B.n43 585
R432 B.n557 B.n556 585
R433 B.n556 B.n555 585
R434 B.n46 B.n45 585
R435 B.n554 B.n46 585
R436 B.n552 B.n551 585
R437 B.n553 B.n552 585
R438 B.n550 B.n51 585
R439 B.n51 B.n50 585
R440 B.n549 B.n548 585
R441 B.n548 B.n547 585
R442 B.n53 B.n52 585
R443 B.n546 B.n53 585
R444 B.n605 B.n604 585
R445 B.n603 B.n2 585
R446 B.n91 B.n53 564.573
R447 B.n544 B.n55 564.573
R448 B.n414 B.n261 564.573
R449 B.n410 B.n259 564.573
R450 B.n89 B.t10 306.026
R451 B.n86 B.t17 306.026
R452 B.n296 B.t6 306.026
R453 B.n293 B.t14 306.026
R454 B.n545 B.n84 256.663
R455 B.n545 B.n83 256.663
R456 B.n545 B.n82 256.663
R457 B.n545 B.n81 256.663
R458 B.n545 B.n80 256.663
R459 B.n545 B.n79 256.663
R460 B.n545 B.n78 256.663
R461 B.n545 B.n77 256.663
R462 B.n545 B.n76 256.663
R463 B.n545 B.n75 256.663
R464 B.n545 B.n74 256.663
R465 B.n545 B.n73 256.663
R466 B.n545 B.n72 256.663
R467 B.n545 B.n71 256.663
R468 B.n545 B.n70 256.663
R469 B.n545 B.n69 256.663
R470 B.n545 B.n68 256.663
R471 B.n545 B.n67 256.663
R472 B.n545 B.n66 256.663
R473 B.n545 B.n65 256.663
R474 B.n545 B.n64 256.663
R475 B.n545 B.n63 256.663
R476 B.n545 B.n62 256.663
R477 B.n545 B.n61 256.663
R478 B.n545 B.n60 256.663
R479 B.n545 B.n59 256.663
R480 B.n545 B.n58 256.663
R481 B.n545 B.n57 256.663
R482 B.n545 B.n56 256.663
R483 B.n412 B.n411 256.663
R484 B.n412 B.n264 256.663
R485 B.n412 B.n265 256.663
R486 B.n412 B.n266 256.663
R487 B.n412 B.n267 256.663
R488 B.n412 B.n268 256.663
R489 B.n412 B.n269 256.663
R490 B.n412 B.n270 256.663
R491 B.n412 B.n271 256.663
R492 B.n412 B.n272 256.663
R493 B.n412 B.n273 256.663
R494 B.n412 B.n274 256.663
R495 B.n412 B.n275 256.663
R496 B.n412 B.n276 256.663
R497 B.n412 B.n277 256.663
R498 B.n412 B.n278 256.663
R499 B.n412 B.n279 256.663
R500 B.n412 B.n280 256.663
R501 B.n412 B.n281 256.663
R502 B.n412 B.n282 256.663
R503 B.n412 B.n283 256.663
R504 B.n412 B.n284 256.663
R505 B.n412 B.n285 256.663
R506 B.n412 B.n286 256.663
R507 B.n412 B.n287 256.663
R508 B.n412 B.n288 256.663
R509 B.n412 B.n289 256.663
R510 B.n412 B.n290 256.663
R511 B.n413 B.n412 256.663
R512 B.n607 B.n606 256.663
R513 B.n95 B.n94 163.367
R514 B.n99 B.n98 163.367
R515 B.n103 B.n102 163.367
R516 B.n107 B.n106 163.367
R517 B.n111 B.n110 163.367
R518 B.n115 B.n114 163.367
R519 B.n119 B.n118 163.367
R520 B.n123 B.n122 163.367
R521 B.n127 B.n126 163.367
R522 B.n131 B.n130 163.367
R523 B.n135 B.n134 163.367
R524 B.n139 B.n138 163.367
R525 B.n144 B.n143 163.367
R526 B.n148 B.n147 163.367
R527 B.n152 B.n151 163.367
R528 B.n156 B.n155 163.367
R529 B.n160 B.n159 163.367
R530 B.n164 B.n163 163.367
R531 B.n168 B.n167 163.367
R532 B.n172 B.n171 163.367
R533 B.n176 B.n175 163.367
R534 B.n180 B.n179 163.367
R535 B.n184 B.n183 163.367
R536 B.n188 B.n187 163.367
R537 B.n192 B.n191 163.367
R538 B.n196 B.n195 163.367
R539 B.n200 B.n199 163.367
R540 B.n204 B.n203 163.367
R541 B.n544 B.n85 163.367
R542 B.n418 B.n261 163.367
R543 B.n418 B.n255 163.367
R544 B.n426 B.n255 163.367
R545 B.n426 B.n253 163.367
R546 B.n430 B.n253 163.367
R547 B.n430 B.n247 163.367
R548 B.n438 B.n247 163.367
R549 B.n438 B.n245 163.367
R550 B.n442 B.n245 163.367
R551 B.n442 B.n239 163.367
R552 B.n450 B.n239 163.367
R553 B.n450 B.n237 163.367
R554 B.n454 B.n237 163.367
R555 B.n454 B.n232 163.367
R556 B.n463 B.n232 163.367
R557 B.n463 B.n230 163.367
R558 B.n467 B.n230 163.367
R559 B.n467 B.n224 163.367
R560 B.n475 B.n224 163.367
R561 B.n475 B.n222 163.367
R562 B.n479 B.n222 163.367
R563 B.n479 B.n216 163.367
R564 B.n487 B.n216 163.367
R565 B.n487 B.n214 163.367
R566 B.n492 B.n214 163.367
R567 B.n492 B.n208 163.367
R568 B.n500 B.n208 163.367
R569 B.n501 B.n500 163.367
R570 B.n501 B.n5 163.367
R571 B.n6 B.n5 163.367
R572 B.n7 B.n6 163.367
R573 B.n507 B.n7 163.367
R574 B.n509 B.n507 163.367
R575 B.n509 B.n12 163.367
R576 B.n13 B.n12 163.367
R577 B.n14 B.n13 163.367
R578 B.n514 B.n14 163.367
R579 B.n514 B.n19 163.367
R580 B.n20 B.n19 163.367
R581 B.n21 B.n20 163.367
R582 B.n519 B.n21 163.367
R583 B.n519 B.n26 163.367
R584 B.n27 B.n26 163.367
R585 B.n28 B.n27 163.367
R586 B.n524 B.n28 163.367
R587 B.n524 B.n33 163.367
R588 B.n34 B.n33 163.367
R589 B.n35 B.n34 163.367
R590 B.n529 B.n35 163.367
R591 B.n529 B.n40 163.367
R592 B.n41 B.n40 163.367
R593 B.n42 B.n41 163.367
R594 B.n534 B.n42 163.367
R595 B.n534 B.n47 163.367
R596 B.n48 B.n47 163.367
R597 B.n49 B.n48 163.367
R598 B.n539 B.n49 163.367
R599 B.n539 B.n54 163.367
R600 B.n55 B.n54 163.367
R601 B.n292 B.n291 163.367
R602 B.n405 B.n291 163.367
R603 B.n403 B.n402 163.367
R604 B.n399 B.n398 163.367
R605 B.n395 B.n394 163.367
R606 B.n391 B.n390 163.367
R607 B.n387 B.n386 163.367
R608 B.n383 B.n382 163.367
R609 B.n379 B.n378 163.367
R610 B.n375 B.n374 163.367
R611 B.n371 B.n370 163.367
R612 B.n367 B.n366 163.367
R613 B.n363 B.n362 163.367
R614 B.n359 B.n358 163.367
R615 B.n355 B.n354 163.367
R616 B.n351 B.n350 163.367
R617 B.n347 B.n346 163.367
R618 B.n342 B.n341 163.367
R619 B.n338 B.n337 163.367
R620 B.n334 B.n333 163.367
R621 B.n330 B.n329 163.367
R622 B.n326 B.n325 163.367
R623 B.n322 B.n321 163.367
R624 B.n318 B.n317 163.367
R625 B.n314 B.n313 163.367
R626 B.n310 B.n309 163.367
R627 B.n306 B.n305 163.367
R628 B.n302 B.n301 163.367
R629 B.n298 B.n263 163.367
R630 B.n420 B.n259 163.367
R631 B.n420 B.n257 163.367
R632 B.n424 B.n257 163.367
R633 B.n424 B.n251 163.367
R634 B.n432 B.n251 163.367
R635 B.n432 B.n249 163.367
R636 B.n436 B.n249 163.367
R637 B.n436 B.n243 163.367
R638 B.n444 B.n243 163.367
R639 B.n444 B.n241 163.367
R640 B.n448 B.n241 163.367
R641 B.n448 B.n235 163.367
R642 B.n457 B.n235 163.367
R643 B.n457 B.n233 163.367
R644 B.n461 B.n233 163.367
R645 B.n461 B.n228 163.367
R646 B.n469 B.n228 163.367
R647 B.n469 B.n226 163.367
R648 B.n473 B.n226 163.367
R649 B.n473 B.n220 163.367
R650 B.n481 B.n220 163.367
R651 B.n481 B.n218 163.367
R652 B.n485 B.n218 163.367
R653 B.n485 B.n212 163.367
R654 B.n494 B.n212 163.367
R655 B.n494 B.n210 163.367
R656 B.n498 B.n210 163.367
R657 B.n498 B.n3 163.367
R658 B.n605 B.n3 163.367
R659 B.n601 B.n2 163.367
R660 B.n601 B.n600 163.367
R661 B.n600 B.n9 163.367
R662 B.n596 B.n9 163.367
R663 B.n596 B.n11 163.367
R664 B.n592 B.n11 163.367
R665 B.n592 B.n16 163.367
R666 B.n588 B.n16 163.367
R667 B.n588 B.n18 163.367
R668 B.n584 B.n18 163.367
R669 B.n584 B.n23 163.367
R670 B.n580 B.n23 163.367
R671 B.n580 B.n25 163.367
R672 B.n576 B.n25 163.367
R673 B.n576 B.n29 163.367
R674 B.n572 B.n29 163.367
R675 B.n572 B.n31 163.367
R676 B.n568 B.n31 163.367
R677 B.n568 B.n37 163.367
R678 B.n564 B.n37 163.367
R679 B.n564 B.n39 163.367
R680 B.n560 B.n39 163.367
R681 B.n560 B.n44 163.367
R682 B.n556 B.n44 163.367
R683 B.n556 B.n46 163.367
R684 B.n552 B.n46 163.367
R685 B.n552 B.n51 163.367
R686 B.n548 B.n51 163.367
R687 B.n548 B.n53 163.367
R688 B.n412 B.n260 133.996
R689 B.n546 B.n545 133.996
R690 B.n86 B.t18 108.462
R691 B.n296 B.t9 108.462
R692 B.n89 B.t12 108.454
R693 B.n293 B.t16 108.454
R694 B.n87 B.t19 72.7769
R695 B.n297 B.t8 72.7769
R696 B.n90 B.t13 72.7701
R697 B.n294 B.t15 72.7701
R698 B.n91 B.n56 71.676
R699 B.n95 B.n57 71.676
R700 B.n99 B.n58 71.676
R701 B.n103 B.n59 71.676
R702 B.n107 B.n60 71.676
R703 B.n111 B.n61 71.676
R704 B.n115 B.n62 71.676
R705 B.n119 B.n63 71.676
R706 B.n123 B.n64 71.676
R707 B.n127 B.n65 71.676
R708 B.n131 B.n66 71.676
R709 B.n135 B.n67 71.676
R710 B.n139 B.n68 71.676
R711 B.n144 B.n69 71.676
R712 B.n148 B.n70 71.676
R713 B.n152 B.n71 71.676
R714 B.n156 B.n72 71.676
R715 B.n160 B.n73 71.676
R716 B.n164 B.n74 71.676
R717 B.n168 B.n75 71.676
R718 B.n172 B.n76 71.676
R719 B.n176 B.n77 71.676
R720 B.n180 B.n78 71.676
R721 B.n184 B.n79 71.676
R722 B.n188 B.n80 71.676
R723 B.n192 B.n81 71.676
R724 B.n196 B.n82 71.676
R725 B.n200 B.n83 71.676
R726 B.n204 B.n84 71.676
R727 B.n85 B.n84 71.676
R728 B.n203 B.n83 71.676
R729 B.n199 B.n82 71.676
R730 B.n195 B.n81 71.676
R731 B.n191 B.n80 71.676
R732 B.n187 B.n79 71.676
R733 B.n183 B.n78 71.676
R734 B.n179 B.n77 71.676
R735 B.n175 B.n76 71.676
R736 B.n171 B.n75 71.676
R737 B.n167 B.n74 71.676
R738 B.n163 B.n73 71.676
R739 B.n159 B.n72 71.676
R740 B.n155 B.n71 71.676
R741 B.n151 B.n70 71.676
R742 B.n147 B.n69 71.676
R743 B.n143 B.n68 71.676
R744 B.n138 B.n67 71.676
R745 B.n134 B.n66 71.676
R746 B.n130 B.n65 71.676
R747 B.n126 B.n64 71.676
R748 B.n122 B.n63 71.676
R749 B.n118 B.n62 71.676
R750 B.n114 B.n61 71.676
R751 B.n110 B.n60 71.676
R752 B.n106 B.n59 71.676
R753 B.n102 B.n58 71.676
R754 B.n98 B.n57 71.676
R755 B.n94 B.n56 71.676
R756 B.n411 B.n410 71.676
R757 B.n405 B.n264 71.676
R758 B.n402 B.n265 71.676
R759 B.n398 B.n266 71.676
R760 B.n394 B.n267 71.676
R761 B.n390 B.n268 71.676
R762 B.n386 B.n269 71.676
R763 B.n382 B.n270 71.676
R764 B.n378 B.n271 71.676
R765 B.n374 B.n272 71.676
R766 B.n370 B.n273 71.676
R767 B.n366 B.n274 71.676
R768 B.n362 B.n275 71.676
R769 B.n358 B.n276 71.676
R770 B.n354 B.n277 71.676
R771 B.n350 B.n278 71.676
R772 B.n346 B.n279 71.676
R773 B.n341 B.n280 71.676
R774 B.n337 B.n281 71.676
R775 B.n333 B.n282 71.676
R776 B.n329 B.n283 71.676
R777 B.n325 B.n284 71.676
R778 B.n321 B.n285 71.676
R779 B.n317 B.n286 71.676
R780 B.n313 B.n287 71.676
R781 B.n309 B.n288 71.676
R782 B.n305 B.n289 71.676
R783 B.n301 B.n290 71.676
R784 B.n413 B.n263 71.676
R785 B.n411 B.n292 71.676
R786 B.n403 B.n264 71.676
R787 B.n399 B.n265 71.676
R788 B.n395 B.n266 71.676
R789 B.n391 B.n267 71.676
R790 B.n387 B.n268 71.676
R791 B.n383 B.n269 71.676
R792 B.n379 B.n270 71.676
R793 B.n375 B.n271 71.676
R794 B.n371 B.n272 71.676
R795 B.n367 B.n273 71.676
R796 B.n363 B.n274 71.676
R797 B.n359 B.n275 71.676
R798 B.n355 B.n276 71.676
R799 B.n351 B.n277 71.676
R800 B.n347 B.n278 71.676
R801 B.n342 B.n279 71.676
R802 B.n338 B.n280 71.676
R803 B.n334 B.n281 71.676
R804 B.n330 B.n282 71.676
R805 B.n326 B.n283 71.676
R806 B.n322 B.n284 71.676
R807 B.n318 B.n285 71.676
R808 B.n314 B.n286 71.676
R809 B.n310 B.n287 71.676
R810 B.n306 B.n288 71.676
R811 B.n302 B.n289 71.676
R812 B.n298 B.n290 71.676
R813 B.n414 B.n413 71.676
R814 B.n606 B.n605 71.676
R815 B.n606 B.n2 71.676
R816 B.n419 B.n260 64.6225
R817 B.n419 B.n256 64.6225
R818 B.n425 B.n256 64.6225
R819 B.n425 B.n252 64.6225
R820 B.n431 B.n252 64.6225
R821 B.n437 B.n248 64.6225
R822 B.n437 B.n244 64.6225
R823 B.n443 B.n244 64.6225
R824 B.n443 B.n240 64.6225
R825 B.n449 B.n240 64.6225
R826 B.n449 B.n236 64.6225
R827 B.n456 B.n236 64.6225
R828 B.n456 B.n455 64.6225
R829 B.n462 B.n229 64.6225
R830 B.n468 B.n229 64.6225
R831 B.n468 B.n225 64.6225
R832 B.n474 B.n225 64.6225
R833 B.n480 B.n221 64.6225
R834 B.n480 B.n217 64.6225
R835 B.n486 B.n217 64.6225
R836 B.n486 B.n213 64.6225
R837 B.n493 B.n213 64.6225
R838 B.n499 B.n209 64.6225
R839 B.n499 B.n4 64.6225
R840 B.n604 B.n4 64.6225
R841 B.n604 B.n603 64.6225
R842 B.n603 B.n602 64.6225
R843 B.n602 B.n8 64.6225
R844 B.n508 B.n8 64.6225
R845 B.n595 B.n594 64.6225
R846 B.n594 B.n593 64.6225
R847 B.n593 B.n15 64.6225
R848 B.n587 B.n15 64.6225
R849 B.n587 B.n586 64.6225
R850 B.n585 B.n22 64.6225
R851 B.n579 B.n22 64.6225
R852 B.n579 B.n578 64.6225
R853 B.n578 B.n577 64.6225
R854 B.n571 B.n32 64.6225
R855 B.n571 B.n570 64.6225
R856 B.n570 B.n569 64.6225
R857 B.n569 B.n36 64.6225
R858 B.n563 B.n36 64.6225
R859 B.n563 B.n562 64.6225
R860 B.n562 B.n561 64.6225
R861 B.n561 B.n43 64.6225
R862 B.n555 B.n554 64.6225
R863 B.n554 B.n553 64.6225
R864 B.n553 B.n50 64.6225
R865 B.n547 B.n50 64.6225
R866 B.n547 B.n546 64.6225
R867 B.n141 B.n90 59.5399
R868 B.n88 B.n87 59.5399
R869 B.n344 B.n297 59.5399
R870 B.n295 B.n294 59.5399
R871 B.t0 B.n209 52.2683
R872 B.n508 B.t3 52.2683
R873 B.n474 B.t4 50.3677
R874 B.t2 B.n585 50.3677
R875 B.n431 B.t7 48.467
R876 B.n555 B.t11 48.467
R877 B.n462 B.t1 40.8644
R878 B.n577 B.t5 40.8644
R879 B.n409 B.n258 36.6834
R880 B.n416 B.n415 36.6834
R881 B.n543 B.n542 36.6834
R882 B.n92 B.n52 36.6834
R883 B.n90 B.n89 35.6853
R884 B.n87 B.n86 35.6853
R885 B.n297 B.n296 35.6853
R886 B.n294 B.n293 35.6853
R887 B.n455 B.t1 23.7586
R888 B.n32 B.t5 23.7586
R889 B B.n607 18.0485
R890 B.t7 B.n248 16.156
R891 B.t11 B.n43 16.156
R892 B.t4 B.n221 14.2554
R893 B.n586 B.t2 14.2554
R894 B.n493 B.t0 12.3547
R895 B.n595 B.t3 12.3547
R896 B.n421 B.n258 10.6151
R897 B.n422 B.n421 10.6151
R898 B.n423 B.n422 10.6151
R899 B.n423 B.n250 10.6151
R900 B.n433 B.n250 10.6151
R901 B.n434 B.n433 10.6151
R902 B.n435 B.n434 10.6151
R903 B.n435 B.n242 10.6151
R904 B.n445 B.n242 10.6151
R905 B.n446 B.n445 10.6151
R906 B.n447 B.n446 10.6151
R907 B.n447 B.n234 10.6151
R908 B.n458 B.n234 10.6151
R909 B.n459 B.n458 10.6151
R910 B.n460 B.n459 10.6151
R911 B.n460 B.n227 10.6151
R912 B.n470 B.n227 10.6151
R913 B.n471 B.n470 10.6151
R914 B.n472 B.n471 10.6151
R915 B.n472 B.n219 10.6151
R916 B.n482 B.n219 10.6151
R917 B.n483 B.n482 10.6151
R918 B.n484 B.n483 10.6151
R919 B.n484 B.n211 10.6151
R920 B.n495 B.n211 10.6151
R921 B.n496 B.n495 10.6151
R922 B.n497 B.n496 10.6151
R923 B.n497 B.n0 10.6151
R924 B.n409 B.n408 10.6151
R925 B.n408 B.n407 10.6151
R926 B.n407 B.n406 10.6151
R927 B.n406 B.n404 10.6151
R928 B.n404 B.n401 10.6151
R929 B.n401 B.n400 10.6151
R930 B.n400 B.n397 10.6151
R931 B.n397 B.n396 10.6151
R932 B.n396 B.n393 10.6151
R933 B.n393 B.n392 10.6151
R934 B.n392 B.n389 10.6151
R935 B.n389 B.n388 10.6151
R936 B.n388 B.n385 10.6151
R937 B.n385 B.n384 10.6151
R938 B.n384 B.n381 10.6151
R939 B.n381 B.n380 10.6151
R940 B.n380 B.n377 10.6151
R941 B.n377 B.n376 10.6151
R942 B.n376 B.n373 10.6151
R943 B.n373 B.n372 10.6151
R944 B.n372 B.n369 10.6151
R945 B.n369 B.n368 10.6151
R946 B.n368 B.n365 10.6151
R947 B.n365 B.n364 10.6151
R948 B.n361 B.n360 10.6151
R949 B.n360 B.n357 10.6151
R950 B.n357 B.n356 10.6151
R951 B.n356 B.n353 10.6151
R952 B.n353 B.n352 10.6151
R953 B.n352 B.n349 10.6151
R954 B.n349 B.n348 10.6151
R955 B.n348 B.n345 10.6151
R956 B.n343 B.n340 10.6151
R957 B.n340 B.n339 10.6151
R958 B.n339 B.n336 10.6151
R959 B.n336 B.n335 10.6151
R960 B.n335 B.n332 10.6151
R961 B.n332 B.n331 10.6151
R962 B.n331 B.n328 10.6151
R963 B.n328 B.n327 10.6151
R964 B.n327 B.n324 10.6151
R965 B.n324 B.n323 10.6151
R966 B.n323 B.n320 10.6151
R967 B.n320 B.n319 10.6151
R968 B.n319 B.n316 10.6151
R969 B.n316 B.n315 10.6151
R970 B.n315 B.n312 10.6151
R971 B.n312 B.n311 10.6151
R972 B.n311 B.n308 10.6151
R973 B.n308 B.n307 10.6151
R974 B.n307 B.n304 10.6151
R975 B.n304 B.n303 10.6151
R976 B.n303 B.n300 10.6151
R977 B.n300 B.n299 10.6151
R978 B.n299 B.n262 10.6151
R979 B.n415 B.n262 10.6151
R980 B.n417 B.n416 10.6151
R981 B.n417 B.n254 10.6151
R982 B.n427 B.n254 10.6151
R983 B.n428 B.n427 10.6151
R984 B.n429 B.n428 10.6151
R985 B.n429 B.n246 10.6151
R986 B.n439 B.n246 10.6151
R987 B.n440 B.n439 10.6151
R988 B.n441 B.n440 10.6151
R989 B.n441 B.n238 10.6151
R990 B.n451 B.n238 10.6151
R991 B.n452 B.n451 10.6151
R992 B.n453 B.n452 10.6151
R993 B.n453 B.n231 10.6151
R994 B.n464 B.n231 10.6151
R995 B.n465 B.n464 10.6151
R996 B.n466 B.n465 10.6151
R997 B.n466 B.n223 10.6151
R998 B.n476 B.n223 10.6151
R999 B.n477 B.n476 10.6151
R1000 B.n478 B.n477 10.6151
R1001 B.n478 B.n215 10.6151
R1002 B.n488 B.n215 10.6151
R1003 B.n489 B.n488 10.6151
R1004 B.n491 B.n489 10.6151
R1005 B.n491 B.n490 10.6151
R1006 B.n490 B.n207 10.6151
R1007 B.n502 B.n207 10.6151
R1008 B.n503 B.n502 10.6151
R1009 B.n504 B.n503 10.6151
R1010 B.n505 B.n504 10.6151
R1011 B.n506 B.n505 10.6151
R1012 B.n510 B.n506 10.6151
R1013 B.n511 B.n510 10.6151
R1014 B.n512 B.n511 10.6151
R1015 B.n513 B.n512 10.6151
R1016 B.n515 B.n513 10.6151
R1017 B.n516 B.n515 10.6151
R1018 B.n517 B.n516 10.6151
R1019 B.n518 B.n517 10.6151
R1020 B.n520 B.n518 10.6151
R1021 B.n521 B.n520 10.6151
R1022 B.n522 B.n521 10.6151
R1023 B.n523 B.n522 10.6151
R1024 B.n525 B.n523 10.6151
R1025 B.n526 B.n525 10.6151
R1026 B.n527 B.n526 10.6151
R1027 B.n528 B.n527 10.6151
R1028 B.n530 B.n528 10.6151
R1029 B.n531 B.n530 10.6151
R1030 B.n532 B.n531 10.6151
R1031 B.n533 B.n532 10.6151
R1032 B.n535 B.n533 10.6151
R1033 B.n536 B.n535 10.6151
R1034 B.n537 B.n536 10.6151
R1035 B.n538 B.n537 10.6151
R1036 B.n540 B.n538 10.6151
R1037 B.n541 B.n540 10.6151
R1038 B.n542 B.n541 10.6151
R1039 B.n599 B.n1 10.6151
R1040 B.n599 B.n598 10.6151
R1041 B.n598 B.n597 10.6151
R1042 B.n597 B.n10 10.6151
R1043 B.n591 B.n10 10.6151
R1044 B.n591 B.n590 10.6151
R1045 B.n590 B.n589 10.6151
R1046 B.n589 B.n17 10.6151
R1047 B.n583 B.n17 10.6151
R1048 B.n583 B.n582 10.6151
R1049 B.n582 B.n581 10.6151
R1050 B.n581 B.n24 10.6151
R1051 B.n575 B.n24 10.6151
R1052 B.n575 B.n574 10.6151
R1053 B.n574 B.n573 10.6151
R1054 B.n573 B.n30 10.6151
R1055 B.n567 B.n30 10.6151
R1056 B.n567 B.n566 10.6151
R1057 B.n566 B.n565 10.6151
R1058 B.n565 B.n38 10.6151
R1059 B.n559 B.n38 10.6151
R1060 B.n559 B.n558 10.6151
R1061 B.n558 B.n557 10.6151
R1062 B.n557 B.n45 10.6151
R1063 B.n551 B.n45 10.6151
R1064 B.n551 B.n550 10.6151
R1065 B.n550 B.n549 10.6151
R1066 B.n549 B.n52 10.6151
R1067 B.n93 B.n92 10.6151
R1068 B.n96 B.n93 10.6151
R1069 B.n97 B.n96 10.6151
R1070 B.n100 B.n97 10.6151
R1071 B.n101 B.n100 10.6151
R1072 B.n104 B.n101 10.6151
R1073 B.n105 B.n104 10.6151
R1074 B.n108 B.n105 10.6151
R1075 B.n109 B.n108 10.6151
R1076 B.n112 B.n109 10.6151
R1077 B.n113 B.n112 10.6151
R1078 B.n116 B.n113 10.6151
R1079 B.n117 B.n116 10.6151
R1080 B.n120 B.n117 10.6151
R1081 B.n121 B.n120 10.6151
R1082 B.n124 B.n121 10.6151
R1083 B.n125 B.n124 10.6151
R1084 B.n128 B.n125 10.6151
R1085 B.n129 B.n128 10.6151
R1086 B.n132 B.n129 10.6151
R1087 B.n133 B.n132 10.6151
R1088 B.n136 B.n133 10.6151
R1089 B.n137 B.n136 10.6151
R1090 B.n140 B.n137 10.6151
R1091 B.n145 B.n142 10.6151
R1092 B.n146 B.n145 10.6151
R1093 B.n149 B.n146 10.6151
R1094 B.n150 B.n149 10.6151
R1095 B.n153 B.n150 10.6151
R1096 B.n154 B.n153 10.6151
R1097 B.n157 B.n154 10.6151
R1098 B.n158 B.n157 10.6151
R1099 B.n162 B.n161 10.6151
R1100 B.n165 B.n162 10.6151
R1101 B.n166 B.n165 10.6151
R1102 B.n169 B.n166 10.6151
R1103 B.n170 B.n169 10.6151
R1104 B.n173 B.n170 10.6151
R1105 B.n174 B.n173 10.6151
R1106 B.n177 B.n174 10.6151
R1107 B.n178 B.n177 10.6151
R1108 B.n181 B.n178 10.6151
R1109 B.n182 B.n181 10.6151
R1110 B.n185 B.n182 10.6151
R1111 B.n186 B.n185 10.6151
R1112 B.n189 B.n186 10.6151
R1113 B.n190 B.n189 10.6151
R1114 B.n193 B.n190 10.6151
R1115 B.n194 B.n193 10.6151
R1116 B.n197 B.n194 10.6151
R1117 B.n198 B.n197 10.6151
R1118 B.n201 B.n198 10.6151
R1119 B.n202 B.n201 10.6151
R1120 B.n205 B.n202 10.6151
R1121 B.n206 B.n205 10.6151
R1122 B.n543 B.n206 10.6151
R1123 B.n607 B.n0 8.11757
R1124 B.n607 B.n1 8.11757
R1125 B.n361 B.n295 6.5566
R1126 B.n345 B.n344 6.5566
R1127 B.n142 B.n141 6.5566
R1128 B.n158 B.n88 6.5566
R1129 B.n364 B.n295 4.05904
R1130 B.n344 B.n343 4.05904
R1131 B.n141 B.n140 4.05904
R1132 B.n161 B.n88 4.05904
R1133 VN.n11 VN.n10 181.465
R1134 VN.n23 VN.n22 181.465
R1135 VN.n21 VN.n12 161.3
R1136 VN.n20 VN.n19 161.3
R1137 VN.n18 VN.n13 161.3
R1138 VN.n17 VN.n16 161.3
R1139 VN.n9 VN.n0 161.3
R1140 VN.n8 VN.n7 161.3
R1141 VN.n6 VN.n1 161.3
R1142 VN.n5 VN.n4 161.3
R1143 VN.n2 VN.t5 131.316
R1144 VN.n14 VN.t0 131.316
R1145 VN.n3 VN.t3 100.55
R1146 VN.n10 VN.t1 100.55
R1147 VN.n15 VN.t4 100.55
R1148 VN.n22 VN.t2 100.55
R1149 VN.n8 VN.n1 56.5617
R1150 VN.n20 VN.n13 56.5617
R1151 VN.n3 VN.n2 53.734
R1152 VN.n15 VN.n14 53.734
R1153 VN VN.n23 40.3054
R1154 VN.n4 VN.n1 24.5923
R1155 VN.n9 VN.n8 24.5923
R1156 VN.n16 VN.n13 24.5923
R1157 VN.n21 VN.n20 24.5923
R1158 VN.n17 VN.n14 18.3138
R1159 VN.n5 VN.n2 18.3138
R1160 VN.n4 VN.n3 12.2964
R1161 VN.n16 VN.n15 12.2964
R1162 VN.n10 VN.n9 4.42703
R1163 VN.n22 VN.n21 4.42703
R1164 VN.n23 VN.n12 0.189894
R1165 VN.n19 VN.n12 0.189894
R1166 VN.n19 VN.n18 0.189894
R1167 VN.n18 VN.n17 0.189894
R1168 VN.n6 VN.n5 0.189894
R1169 VN.n7 VN.n6 0.189894
R1170 VN.n7 VN.n0 0.189894
R1171 VN.n11 VN.n0 0.189894
R1172 VN VN.n11 0.0516364
R1173 VDD2.n1 VDD2.t0 69.7094
R1174 VDD2.n2 VDD2.t3 68.5752
R1175 VDD2.n1 VDD2.n0 65.7734
R1176 VDD2 VDD2.n3 65.7706
R1177 VDD2.n2 VDD2.n1 34.3015
R1178 VDD2.n3 VDD2.t1 3.14336
R1179 VDD2.n3 VDD2.t5 3.14336
R1180 VDD2.n0 VDD2.t2 3.14336
R1181 VDD2.n0 VDD2.t4 3.14336
R1182 VDD2 VDD2.n2 1.24834
C0 VP VDD1 3.47741f
C1 VDD2 VDD1 1.01034f
C2 VN VTAIL 3.49191f
C3 VN VDD1 0.149649f
C4 VDD2 VP 0.365787f
C5 VDD1 VTAIL 5.38188f
C6 VP VN 4.81153f
C7 VP VTAIL 3.50618f
C8 VDD2 VN 3.26353f
C9 VDD2 VTAIL 5.42584f
C10 VDD2 B 4.103238f
C11 VDD1 B 4.370496f
C12 VTAIL B 4.643429f
C13 VN B 9.167411f
C14 VP B 7.712544f
C15 VDD2.t0 B 1.17429f
C16 VDD2.t2 B 0.109791f
C17 VDD2.t4 B 0.109791f
C18 VDD2.n0 B 0.922214f
C19 VDD2.n1 B 1.83795f
C20 VDD2.t3 B 1.16907f
C21 VDD2.n2 B 1.79815f
C22 VDD2.t1 B 0.109791f
C23 VDD2.t5 B 0.109791f
C24 VDD2.n3 B 0.92219f
C25 VN.n0 B 0.034485f
C26 VN.t1 B 0.870709f
C27 VN.n1 B 0.042496f
C28 VN.t5 B 0.980786f
C29 VN.n2 B 0.416381f
C30 VN.t3 B 0.870709f
C31 VN.n3 B 0.402053f
C32 VN.n4 B 0.048163f
C33 VN.n5 B 0.21522f
C34 VN.n6 B 0.034485f
C35 VN.n7 B 0.034485f
C36 VN.n8 B 0.057761f
C37 VN.n9 B 0.038061f
C38 VN.n10 B 0.400475f
C39 VN.n11 B 0.034532f
C40 VN.n12 B 0.034485f
C41 VN.t2 B 0.870709f
C42 VN.n13 B 0.042496f
C43 VN.t0 B 0.980786f
C44 VN.n14 B 0.416381f
C45 VN.t4 B 0.870709f
C46 VN.n15 B 0.402053f
C47 VN.n16 B 0.048163f
C48 VN.n17 B 0.21522f
C49 VN.n18 B 0.034485f
C50 VN.n19 B 0.034485f
C51 VN.n20 B 0.057761f
C52 VN.n21 B 0.038061f
C53 VN.n22 B 0.400475f
C54 VN.n23 B 1.33664f
C55 VDD1.t0 B 1.19081f
C56 VDD1.t3 B 1.19014f
C57 VDD1.t2 B 0.111274f
C58 VDD1.t1 B 0.111274f
C59 VDD1.n0 B 0.934663f
C60 VDD1.n1 B 1.9456f
C61 VDD1.t4 B 0.111274f
C62 VDD1.t5 B 0.111274f
C63 VDD1.n2 B 0.93294f
C64 VDD1.n3 B 1.81932f
C65 VTAIL.t11 B 0.127551f
C66 VTAIL.t2 B 0.127551f
C67 VTAIL.n0 B 0.999427f
C68 VTAIL.n1 B 0.386408f
C69 VTAIL.t8 B 1.27342f
C70 VTAIL.n2 B 0.553686f
C71 VTAIL.t5 B 0.127551f
C72 VTAIL.t4 B 0.127551f
C73 VTAIL.n3 B 0.999427f
C74 VTAIL.n4 B 1.43384f
C75 VTAIL.t1 B 0.127551f
C76 VTAIL.t9 B 0.127551f
C77 VTAIL.n5 B 0.999432f
C78 VTAIL.n6 B 1.43383f
C79 VTAIL.t0 B 1.27343f
C80 VTAIL.n7 B 0.553678f
C81 VTAIL.t6 B 0.127551f
C82 VTAIL.t7 B 0.127551f
C83 VTAIL.n8 B 0.999432f
C84 VTAIL.n9 B 0.479811f
C85 VTAIL.t3 B 1.27342f
C86 VTAIL.n10 B 1.37676f
C87 VTAIL.t10 B 1.27342f
C88 VTAIL.n11 B 1.33922f
C89 VP.n0 B 0.035226f
C90 VP.t4 B 0.889438f
C91 VP.n1 B 0.04341f
C92 VP.n2 B 0.035226f
C93 VP.t3 B 0.889438f
C94 VP.n3 B 0.059004f
C95 VP.n4 B 0.035226f
C96 VP.t0 B 0.889438f
C97 VP.n5 B 0.04341f
C98 VP.t5 B 1.00188f
C99 VP.n6 B 0.425338f
C100 VP.t1 B 0.889438f
C101 VP.n7 B 0.410701f
C102 VP.n8 B 0.0492f
C103 VP.n9 B 0.219849f
C104 VP.n10 B 0.035226f
C105 VP.n11 B 0.035226f
C106 VP.n12 B 0.059004f
C107 VP.n13 B 0.03888f
C108 VP.n14 B 0.409089f
C109 VP.n15 B 1.34219f
C110 VP.n16 B 1.374f
C111 VP.t2 B 0.889438f
C112 VP.n17 B 0.409089f
C113 VP.n18 B 0.03888f
C114 VP.n19 B 0.035226f
C115 VP.n20 B 0.035226f
C116 VP.n21 B 0.035226f
C117 VP.n22 B 0.04341f
C118 VP.n23 B 0.0492f
C119 VP.n24 B 0.345291f
C120 VP.n25 B 0.0492f
C121 VP.n26 B 0.035226f
C122 VP.n27 B 0.035226f
C123 VP.n28 B 0.035226f
C124 VP.n29 B 0.059004f
C125 VP.n30 B 0.03888f
C126 VP.n31 B 0.409089f
C127 VP.n32 B 0.035275f
.ends

