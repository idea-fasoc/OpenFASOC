* NGSPICE file created from diff_pair_sample_1684.ext - technology: sky130A

.subckt diff_pair_sample_1684 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n4306_n3544# sky130_fd_pr__pfet_01v8 ad=5.0232 pd=26.54 as=0 ps=0 w=12.88 l=3.84
X1 VDD1.t5 VP.t0 VTAIL.t7 w_n4306_n3544# sky130_fd_pr__pfet_01v8 ad=2.1252 pd=13.21 as=5.0232 ps=26.54 w=12.88 l=3.84
X2 B.t8 B.t6 B.t7 w_n4306_n3544# sky130_fd_pr__pfet_01v8 ad=5.0232 pd=26.54 as=0 ps=0 w=12.88 l=3.84
X3 B.t5 B.t3 B.t4 w_n4306_n3544# sky130_fd_pr__pfet_01v8 ad=5.0232 pd=26.54 as=0 ps=0 w=12.88 l=3.84
X4 VDD1.t4 VP.t1 VTAIL.t9 w_n4306_n3544# sky130_fd_pr__pfet_01v8 ad=2.1252 pd=13.21 as=5.0232 ps=26.54 w=12.88 l=3.84
X5 VDD1.t3 VP.t2 VTAIL.t10 w_n4306_n3544# sky130_fd_pr__pfet_01v8 ad=5.0232 pd=26.54 as=2.1252 ps=13.21 w=12.88 l=3.84
X6 VDD2.t5 VN.t0 VTAIL.t3 w_n4306_n3544# sky130_fd_pr__pfet_01v8 ad=2.1252 pd=13.21 as=5.0232 ps=26.54 w=12.88 l=3.84
X7 VDD2.t4 VN.t1 VTAIL.t1 w_n4306_n3544# sky130_fd_pr__pfet_01v8 ad=5.0232 pd=26.54 as=2.1252 ps=13.21 w=12.88 l=3.84
X8 VTAIL.t0 VN.t2 VDD2.t3 w_n4306_n3544# sky130_fd_pr__pfet_01v8 ad=2.1252 pd=13.21 as=2.1252 ps=13.21 w=12.88 l=3.84
X9 B.t2 B.t0 B.t1 w_n4306_n3544# sky130_fd_pr__pfet_01v8 ad=5.0232 pd=26.54 as=0 ps=0 w=12.88 l=3.84
X10 VTAIL.t8 VP.t3 VDD1.t2 w_n4306_n3544# sky130_fd_pr__pfet_01v8 ad=2.1252 pd=13.21 as=2.1252 ps=13.21 w=12.88 l=3.84
X11 VDD2.t2 VN.t3 VTAIL.t4 w_n4306_n3544# sky130_fd_pr__pfet_01v8 ad=2.1252 pd=13.21 as=5.0232 ps=26.54 w=12.88 l=3.84
X12 VTAIL.t6 VP.t4 VDD1.t1 w_n4306_n3544# sky130_fd_pr__pfet_01v8 ad=2.1252 pd=13.21 as=2.1252 ps=13.21 w=12.88 l=3.84
X13 VDD2.t1 VN.t4 VTAIL.t5 w_n4306_n3544# sky130_fd_pr__pfet_01v8 ad=5.0232 pd=26.54 as=2.1252 ps=13.21 w=12.88 l=3.84
X14 VDD1.t0 VP.t5 VTAIL.t11 w_n4306_n3544# sky130_fd_pr__pfet_01v8 ad=5.0232 pd=26.54 as=2.1252 ps=13.21 w=12.88 l=3.84
X15 VTAIL.t2 VN.t5 VDD2.t0 w_n4306_n3544# sky130_fd_pr__pfet_01v8 ad=2.1252 pd=13.21 as=2.1252 ps=13.21 w=12.88 l=3.84
R0 B.n629 B.n84 585
R1 B.n631 B.n630 585
R2 B.n632 B.n83 585
R3 B.n634 B.n633 585
R4 B.n635 B.n82 585
R5 B.n637 B.n636 585
R6 B.n638 B.n81 585
R7 B.n640 B.n639 585
R8 B.n641 B.n80 585
R9 B.n643 B.n642 585
R10 B.n644 B.n79 585
R11 B.n646 B.n645 585
R12 B.n647 B.n78 585
R13 B.n649 B.n648 585
R14 B.n650 B.n77 585
R15 B.n652 B.n651 585
R16 B.n653 B.n76 585
R17 B.n655 B.n654 585
R18 B.n656 B.n75 585
R19 B.n658 B.n657 585
R20 B.n659 B.n74 585
R21 B.n661 B.n660 585
R22 B.n662 B.n73 585
R23 B.n664 B.n663 585
R24 B.n665 B.n72 585
R25 B.n667 B.n666 585
R26 B.n668 B.n71 585
R27 B.n670 B.n669 585
R28 B.n671 B.n70 585
R29 B.n673 B.n672 585
R30 B.n674 B.n69 585
R31 B.n676 B.n675 585
R32 B.n677 B.n68 585
R33 B.n679 B.n678 585
R34 B.n680 B.n67 585
R35 B.n682 B.n681 585
R36 B.n683 B.n66 585
R37 B.n685 B.n684 585
R38 B.n686 B.n65 585
R39 B.n688 B.n687 585
R40 B.n689 B.n64 585
R41 B.n691 B.n690 585
R42 B.n692 B.n63 585
R43 B.n694 B.n693 585
R44 B.n696 B.n60 585
R45 B.n698 B.n697 585
R46 B.n699 B.n59 585
R47 B.n701 B.n700 585
R48 B.n702 B.n58 585
R49 B.n704 B.n703 585
R50 B.n705 B.n57 585
R51 B.n707 B.n706 585
R52 B.n708 B.n53 585
R53 B.n710 B.n709 585
R54 B.n711 B.n52 585
R55 B.n713 B.n712 585
R56 B.n714 B.n51 585
R57 B.n716 B.n715 585
R58 B.n717 B.n50 585
R59 B.n719 B.n718 585
R60 B.n720 B.n49 585
R61 B.n722 B.n721 585
R62 B.n723 B.n48 585
R63 B.n725 B.n724 585
R64 B.n726 B.n47 585
R65 B.n728 B.n727 585
R66 B.n729 B.n46 585
R67 B.n731 B.n730 585
R68 B.n732 B.n45 585
R69 B.n734 B.n733 585
R70 B.n735 B.n44 585
R71 B.n737 B.n736 585
R72 B.n738 B.n43 585
R73 B.n740 B.n739 585
R74 B.n741 B.n42 585
R75 B.n743 B.n742 585
R76 B.n744 B.n41 585
R77 B.n746 B.n745 585
R78 B.n747 B.n40 585
R79 B.n749 B.n748 585
R80 B.n750 B.n39 585
R81 B.n752 B.n751 585
R82 B.n753 B.n38 585
R83 B.n755 B.n754 585
R84 B.n756 B.n37 585
R85 B.n758 B.n757 585
R86 B.n759 B.n36 585
R87 B.n761 B.n760 585
R88 B.n762 B.n35 585
R89 B.n764 B.n763 585
R90 B.n765 B.n34 585
R91 B.n767 B.n766 585
R92 B.n768 B.n33 585
R93 B.n770 B.n769 585
R94 B.n771 B.n32 585
R95 B.n773 B.n772 585
R96 B.n774 B.n31 585
R97 B.n776 B.n775 585
R98 B.n628 B.n627 585
R99 B.n626 B.n85 585
R100 B.n625 B.n624 585
R101 B.n623 B.n86 585
R102 B.n622 B.n621 585
R103 B.n620 B.n87 585
R104 B.n619 B.n618 585
R105 B.n617 B.n88 585
R106 B.n616 B.n615 585
R107 B.n614 B.n89 585
R108 B.n613 B.n612 585
R109 B.n611 B.n90 585
R110 B.n610 B.n609 585
R111 B.n608 B.n91 585
R112 B.n607 B.n606 585
R113 B.n605 B.n92 585
R114 B.n604 B.n603 585
R115 B.n602 B.n93 585
R116 B.n601 B.n600 585
R117 B.n599 B.n94 585
R118 B.n598 B.n597 585
R119 B.n596 B.n95 585
R120 B.n595 B.n594 585
R121 B.n593 B.n96 585
R122 B.n592 B.n591 585
R123 B.n590 B.n97 585
R124 B.n589 B.n588 585
R125 B.n587 B.n98 585
R126 B.n586 B.n585 585
R127 B.n584 B.n99 585
R128 B.n583 B.n582 585
R129 B.n581 B.n100 585
R130 B.n580 B.n579 585
R131 B.n578 B.n101 585
R132 B.n577 B.n576 585
R133 B.n575 B.n102 585
R134 B.n574 B.n573 585
R135 B.n572 B.n103 585
R136 B.n571 B.n570 585
R137 B.n569 B.n104 585
R138 B.n568 B.n567 585
R139 B.n566 B.n105 585
R140 B.n565 B.n564 585
R141 B.n563 B.n106 585
R142 B.n562 B.n561 585
R143 B.n560 B.n107 585
R144 B.n559 B.n558 585
R145 B.n557 B.n108 585
R146 B.n556 B.n555 585
R147 B.n554 B.n109 585
R148 B.n553 B.n552 585
R149 B.n551 B.n110 585
R150 B.n550 B.n549 585
R151 B.n548 B.n111 585
R152 B.n547 B.n546 585
R153 B.n545 B.n112 585
R154 B.n544 B.n543 585
R155 B.n542 B.n113 585
R156 B.n541 B.n540 585
R157 B.n539 B.n114 585
R158 B.n538 B.n537 585
R159 B.n536 B.n115 585
R160 B.n535 B.n534 585
R161 B.n533 B.n116 585
R162 B.n532 B.n531 585
R163 B.n530 B.n117 585
R164 B.n529 B.n528 585
R165 B.n527 B.n118 585
R166 B.n526 B.n525 585
R167 B.n524 B.n119 585
R168 B.n523 B.n522 585
R169 B.n521 B.n120 585
R170 B.n520 B.n519 585
R171 B.n518 B.n121 585
R172 B.n517 B.n516 585
R173 B.n515 B.n122 585
R174 B.n514 B.n513 585
R175 B.n512 B.n123 585
R176 B.n511 B.n510 585
R177 B.n509 B.n124 585
R178 B.n508 B.n507 585
R179 B.n506 B.n125 585
R180 B.n505 B.n504 585
R181 B.n503 B.n126 585
R182 B.n502 B.n501 585
R183 B.n500 B.n127 585
R184 B.n499 B.n498 585
R185 B.n497 B.n128 585
R186 B.n496 B.n495 585
R187 B.n494 B.n129 585
R188 B.n493 B.n492 585
R189 B.n491 B.n130 585
R190 B.n490 B.n489 585
R191 B.n488 B.n131 585
R192 B.n487 B.n486 585
R193 B.n485 B.n132 585
R194 B.n484 B.n483 585
R195 B.n482 B.n133 585
R196 B.n481 B.n480 585
R197 B.n479 B.n134 585
R198 B.n478 B.n477 585
R199 B.n476 B.n135 585
R200 B.n475 B.n474 585
R201 B.n473 B.n136 585
R202 B.n472 B.n471 585
R203 B.n470 B.n137 585
R204 B.n469 B.n468 585
R205 B.n467 B.n138 585
R206 B.n466 B.n465 585
R207 B.n464 B.n139 585
R208 B.n463 B.n462 585
R209 B.n461 B.n140 585
R210 B.n460 B.n459 585
R211 B.n458 B.n141 585
R212 B.n457 B.n456 585
R213 B.n308 B.n195 585
R214 B.n310 B.n309 585
R215 B.n311 B.n194 585
R216 B.n313 B.n312 585
R217 B.n314 B.n193 585
R218 B.n316 B.n315 585
R219 B.n317 B.n192 585
R220 B.n319 B.n318 585
R221 B.n320 B.n191 585
R222 B.n322 B.n321 585
R223 B.n323 B.n190 585
R224 B.n325 B.n324 585
R225 B.n326 B.n189 585
R226 B.n328 B.n327 585
R227 B.n329 B.n188 585
R228 B.n331 B.n330 585
R229 B.n332 B.n187 585
R230 B.n334 B.n333 585
R231 B.n335 B.n186 585
R232 B.n337 B.n336 585
R233 B.n338 B.n185 585
R234 B.n340 B.n339 585
R235 B.n341 B.n184 585
R236 B.n343 B.n342 585
R237 B.n344 B.n183 585
R238 B.n346 B.n345 585
R239 B.n347 B.n182 585
R240 B.n349 B.n348 585
R241 B.n350 B.n181 585
R242 B.n352 B.n351 585
R243 B.n353 B.n180 585
R244 B.n355 B.n354 585
R245 B.n356 B.n179 585
R246 B.n358 B.n357 585
R247 B.n359 B.n178 585
R248 B.n361 B.n360 585
R249 B.n362 B.n177 585
R250 B.n364 B.n363 585
R251 B.n365 B.n176 585
R252 B.n367 B.n366 585
R253 B.n368 B.n175 585
R254 B.n370 B.n369 585
R255 B.n371 B.n174 585
R256 B.n373 B.n372 585
R257 B.n375 B.n374 585
R258 B.n376 B.n170 585
R259 B.n378 B.n377 585
R260 B.n379 B.n169 585
R261 B.n381 B.n380 585
R262 B.n382 B.n168 585
R263 B.n384 B.n383 585
R264 B.n385 B.n167 585
R265 B.n387 B.n386 585
R266 B.n388 B.n164 585
R267 B.n391 B.n390 585
R268 B.n392 B.n163 585
R269 B.n394 B.n393 585
R270 B.n395 B.n162 585
R271 B.n397 B.n396 585
R272 B.n398 B.n161 585
R273 B.n400 B.n399 585
R274 B.n401 B.n160 585
R275 B.n403 B.n402 585
R276 B.n404 B.n159 585
R277 B.n406 B.n405 585
R278 B.n407 B.n158 585
R279 B.n409 B.n408 585
R280 B.n410 B.n157 585
R281 B.n412 B.n411 585
R282 B.n413 B.n156 585
R283 B.n415 B.n414 585
R284 B.n416 B.n155 585
R285 B.n418 B.n417 585
R286 B.n419 B.n154 585
R287 B.n421 B.n420 585
R288 B.n422 B.n153 585
R289 B.n424 B.n423 585
R290 B.n425 B.n152 585
R291 B.n427 B.n426 585
R292 B.n428 B.n151 585
R293 B.n430 B.n429 585
R294 B.n431 B.n150 585
R295 B.n433 B.n432 585
R296 B.n434 B.n149 585
R297 B.n436 B.n435 585
R298 B.n437 B.n148 585
R299 B.n439 B.n438 585
R300 B.n440 B.n147 585
R301 B.n442 B.n441 585
R302 B.n443 B.n146 585
R303 B.n445 B.n444 585
R304 B.n446 B.n145 585
R305 B.n448 B.n447 585
R306 B.n449 B.n144 585
R307 B.n451 B.n450 585
R308 B.n452 B.n143 585
R309 B.n454 B.n453 585
R310 B.n455 B.n142 585
R311 B.n307 B.n306 585
R312 B.n305 B.n196 585
R313 B.n304 B.n303 585
R314 B.n302 B.n197 585
R315 B.n301 B.n300 585
R316 B.n299 B.n198 585
R317 B.n298 B.n297 585
R318 B.n296 B.n199 585
R319 B.n295 B.n294 585
R320 B.n293 B.n200 585
R321 B.n292 B.n291 585
R322 B.n290 B.n201 585
R323 B.n289 B.n288 585
R324 B.n287 B.n202 585
R325 B.n286 B.n285 585
R326 B.n284 B.n203 585
R327 B.n283 B.n282 585
R328 B.n281 B.n204 585
R329 B.n280 B.n279 585
R330 B.n278 B.n205 585
R331 B.n277 B.n276 585
R332 B.n275 B.n206 585
R333 B.n274 B.n273 585
R334 B.n272 B.n207 585
R335 B.n271 B.n270 585
R336 B.n269 B.n208 585
R337 B.n268 B.n267 585
R338 B.n266 B.n209 585
R339 B.n265 B.n264 585
R340 B.n263 B.n210 585
R341 B.n262 B.n261 585
R342 B.n260 B.n211 585
R343 B.n259 B.n258 585
R344 B.n257 B.n212 585
R345 B.n256 B.n255 585
R346 B.n254 B.n213 585
R347 B.n253 B.n252 585
R348 B.n251 B.n214 585
R349 B.n250 B.n249 585
R350 B.n248 B.n215 585
R351 B.n247 B.n246 585
R352 B.n245 B.n216 585
R353 B.n244 B.n243 585
R354 B.n242 B.n217 585
R355 B.n241 B.n240 585
R356 B.n239 B.n218 585
R357 B.n238 B.n237 585
R358 B.n236 B.n219 585
R359 B.n235 B.n234 585
R360 B.n233 B.n220 585
R361 B.n232 B.n231 585
R362 B.n230 B.n221 585
R363 B.n229 B.n228 585
R364 B.n227 B.n222 585
R365 B.n226 B.n225 585
R366 B.n224 B.n223 585
R367 B.n2 B.n0 585
R368 B.n861 B.n1 585
R369 B.n860 B.n859 585
R370 B.n858 B.n3 585
R371 B.n857 B.n856 585
R372 B.n855 B.n4 585
R373 B.n854 B.n853 585
R374 B.n852 B.n5 585
R375 B.n851 B.n850 585
R376 B.n849 B.n6 585
R377 B.n848 B.n847 585
R378 B.n846 B.n7 585
R379 B.n845 B.n844 585
R380 B.n843 B.n8 585
R381 B.n842 B.n841 585
R382 B.n840 B.n9 585
R383 B.n839 B.n838 585
R384 B.n837 B.n10 585
R385 B.n836 B.n835 585
R386 B.n834 B.n11 585
R387 B.n833 B.n832 585
R388 B.n831 B.n12 585
R389 B.n830 B.n829 585
R390 B.n828 B.n13 585
R391 B.n827 B.n826 585
R392 B.n825 B.n14 585
R393 B.n824 B.n823 585
R394 B.n822 B.n15 585
R395 B.n821 B.n820 585
R396 B.n819 B.n16 585
R397 B.n818 B.n817 585
R398 B.n816 B.n17 585
R399 B.n815 B.n814 585
R400 B.n813 B.n18 585
R401 B.n812 B.n811 585
R402 B.n810 B.n19 585
R403 B.n809 B.n808 585
R404 B.n807 B.n20 585
R405 B.n806 B.n805 585
R406 B.n804 B.n21 585
R407 B.n803 B.n802 585
R408 B.n801 B.n22 585
R409 B.n800 B.n799 585
R410 B.n798 B.n23 585
R411 B.n797 B.n796 585
R412 B.n795 B.n24 585
R413 B.n794 B.n793 585
R414 B.n792 B.n25 585
R415 B.n791 B.n790 585
R416 B.n789 B.n26 585
R417 B.n788 B.n787 585
R418 B.n786 B.n27 585
R419 B.n785 B.n784 585
R420 B.n783 B.n28 585
R421 B.n782 B.n781 585
R422 B.n780 B.n29 585
R423 B.n779 B.n778 585
R424 B.n777 B.n30 585
R425 B.n863 B.n862 585
R426 B.n308 B.n307 526.135
R427 B.n777 B.n776 526.135
R428 B.n457 B.n142 526.135
R429 B.n627 B.n84 526.135
R430 B.n165 B.t11 472.529
R431 B.n61 B.t4 472.529
R432 B.n171 B.t2 472.529
R433 B.n54 B.t7 472.529
R434 B.n166 B.t10 391.656
R435 B.n62 B.t5 391.656
R436 B.n172 B.t1 391.656
R437 B.n55 B.t8 391.656
R438 B.n165 B.t9 290.209
R439 B.n171 B.t0 290.209
R440 B.n54 B.t6 290.209
R441 B.n61 B.t3 290.209
R442 B.n307 B.n196 163.367
R443 B.n303 B.n196 163.367
R444 B.n303 B.n302 163.367
R445 B.n302 B.n301 163.367
R446 B.n301 B.n198 163.367
R447 B.n297 B.n198 163.367
R448 B.n297 B.n296 163.367
R449 B.n296 B.n295 163.367
R450 B.n295 B.n200 163.367
R451 B.n291 B.n200 163.367
R452 B.n291 B.n290 163.367
R453 B.n290 B.n289 163.367
R454 B.n289 B.n202 163.367
R455 B.n285 B.n202 163.367
R456 B.n285 B.n284 163.367
R457 B.n284 B.n283 163.367
R458 B.n283 B.n204 163.367
R459 B.n279 B.n204 163.367
R460 B.n279 B.n278 163.367
R461 B.n278 B.n277 163.367
R462 B.n277 B.n206 163.367
R463 B.n273 B.n206 163.367
R464 B.n273 B.n272 163.367
R465 B.n272 B.n271 163.367
R466 B.n271 B.n208 163.367
R467 B.n267 B.n208 163.367
R468 B.n267 B.n266 163.367
R469 B.n266 B.n265 163.367
R470 B.n265 B.n210 163.367
R471 B.n261 B.n210 163.367
R472 B.n261 B.n260 163.367
R473 B.n260 B.n259 163.367
R474 B.n259 B.n212 163.367
R475 B.n255 B.n212 163.367
R476 B.n255 B.n254 163.367
R477 B.n254 B.n253 163.367
R478 B.n253 B.n214 163.367
R479 B.n249 B.n214 163.367
R480 B.n249 B.n248 163.367
R481 B.n248 B.n247 163.367
R482 B.n247 B.n216 163.367
R483 B.n243 B.n216 163.367
R484 B.n243 B.n242 163.367
R485 B.n242 B.n241 163.367
R486 B.n241 B.n218 163.367
R487 B.n237 B.n218 163.367
R488 B.n237 B.n236 163.367
R489 B.n236 B.n235 163.367
R490 B.n235 B.n220 163.367
R491 B.n231 B.n220 163.367
R492 B.n231 B.n230 163.367
R493 B.n230 B.n229 163.367
R494 B.n229 B.n222 163.367
R495 B.n225 B.n222 163.367
R496 B.n225 B.n224 163.367
R497 B.n224 B.n2 163.367
R498 B.n862 B.n2 163.367
R499 B.n862 B.n861 163.367
R500 B.n861 B.n860 163.367
R501 B.n860 B.n3 163.367
R502 B.n856 B.n3 163.367
R503 B.n856 B.n855 163.367
R504 B.n855 B.n854 163.367
R505 B.n854 B.n5 163.367
R506 B.n850 B.n5 163.367
R507 B.n850 B.n849 163.367
R508 B.n849 B.n848 163.367
R509 B.n848 B.n7 163.367
R510 B.n844 B.n7 163.367
R511 B.n844 B.n843 163.367
R512 B.n843 B.n842 163.367
R513 B.n842 B.n9 163.367
R514 B.n838 B.n9 163.367
R515 B.n838 B.n837 163.367
R516 B.n837 B.n836 163.367
R517 B.n836 B.n11 163.367
R518 B.n832 B.n11 163.367
R519 B.n832 B.n831 163.367
R520 B.n831 B.n830 163.367
R521 B.n830 B.n13 163.367
R522 B.n826 B.n13 163.367
R523 B.n826 B.n825 163.367
R524 B.n825 B.n824 163.367
R525 B.n824 B.n15 163.367
R526 B.n820 B.n15 163.367
R527 B.n820 B.n819 163.367
R528 B.n819 B.n818 163.367
R529 B.n818 B.n17 163.367
R530 B.n814 B.n17 163.367
R531 B.n814 B.n813 163.367
R532 B.n813 B.n812 163.367
R533 B.n812 B.n19 163.367
R534 B.n808 B.n19 163.367
R535 B.n808 B.n807 163.367
R536 B.n807 B.n806 163.367
R537 B.n806 B.n21 163.367
R538 B.n802 B.n21 163.367
R539 B.n802 B.n801 163.367
R540 B.n801 B.n800 163.367
R541 B.n800 B.n23 163.367
R542 B.n796 B.n23 163.367
R543 B.n796 B.n795 163.367
R544 B.n795 B.n794 163.367
R545 B.n794 B.n25 163.367
R546 B.n790 B.n25 163.367
R547 B.n790 B.n789 163.367
R548 B.n789 B.n788 163.367
R549 B.n788 B.n27 163.367
R550 B.n784 B.n27 163.367
R551 B.n784 B.n783 163.367
R552 B.n783 B.n782 163.367
R553 B.n782 B.n29 163.367
R554 B.n778 B.n29 163.367
R555 B.n778 B.n777 163.367
R556 B.n309 B.n308 163.367
R557 B.n309 B.n194 163.367
R558 B.n313 B.n194 163.367
R559 B.n314 B.n313 163.367
R560 B.n315 B.n314 163.367
R561 B.n315 B.n192 163.367
R562 B.n319 B.n192 163.367
R563 B.n320 B.n319 163.367
R564 B.n321 B.n320 163.367
R565 B.n321 B.n190 163.367
R566 B.n325 B.n190 163.367
R567 B.n326 B.n325 163.367
R568 B.n327 B.n326 163.367
R569 B.n327 B.n188 163.367
R570 B.n331 B.n188 163.367
R571 B.n332 B.n331 163.367
R572 B.n333 B.n332 163.367
R573 B.n333 B.n186 163.367
R574 B.n337 B.n186 163.367
R575 B.n338 B.n337 163.367
R576 B.n339 B.n338 163.367
R577 B.n339 B.n184 163.367
R578 B.n343 B.n184 163.367
R579 B.n344 B.n343 163.367
R580 B.n345 B.n344 163.367
R581 B.n345 B.n182 163.367
R582 B.n349 B.n182 163.367
R583 B.n350 B.n349 163.367
R584 B.n351 B.n350 163.367
R585 B.n351 B.n180 163.367
R586 B.n355 B.n180 163.367
R587 B.n356 B.n355 163.367
R588 B.n357 B.n356 163.367
R589 B.n357 B.n178 163.367
R590 B.n361 B.n178 163.367
R591 B.n362 B.n361 163.367
R592 B.n363 B.n362 163.367
R593 B.n363 B.n176 163.367
R594 B.n367 B.n176 163.367
R595 B.n368 B.n367 163.367
R596 B.n369 B.n368 163.367
R597 B.n369 B.n174 163.367
R598 B.n373 B.n174 163.367
R599 B.n374 B.n373 163.367
R600 B.n374 B.n170 163.367
R601 B.n378 B.n170 163.367
R602 B.n379 B.n378 163.367
R603 B.n380 B.n379 163.367
R604 B.n380 B.n168 163.367
R605 B.n384 B.n168 163.367
R606 B.n385 B.n384 163.367
R607 B.n386 B.n385 163.367
R608 B.n386 B.n164 163.367
R609 B.n391 B.n164 163.367
R610 B.n392 B.n391 163.367
R611 B.n393 B.n392 163.367
R612 B.n393 B.n162 163.367
R613 B.n397 B.n162 163.367
R614 B.n398 B.n397 163.367
R615 B.n399 B.n398 163.367
R616 B.n399 B.n160 163.367
R617 B.n403 B.n160 163.367
R618 B.n404 B.n403 163.367
R619 B.n405 B.n404 163.367
R620 B.n405 B.n158 163.367
R621 B.n409 B.n158 163.367
R622 B.n410 B.n409 163.367
R623 B.n411 B.n410 163.367
R624 B.n411 B.n156 163.367
R625 B.n415 B.n156 163.367
R626 B.n416 B.n415 163.367
R627 B.n417 B.n416 163.367
R628 B.n417 B.n154 163.367
R629 B.n421 B.n154 163.367
R630 B.n422 B.n421 163.367
R631 B.n423 B.n422 163.367
R632 B.n423 B.n152 163.367
R633 B.n427 B.n152 163.367
R634 B.n428 B.n427 163.367
R635 B.n429 B.n428 163.367
R636 B.n429 B.n150 163.367
R637 B.n433 B.n150 163.367
R638 B.n434 B.n433 163.367
R639 B.n435 B.n434 163.367
R640 B.n435 B.n148 163.367
R641 B.n439 B.n148 163.367
R642 B.n440 B.n439 163.367
R643 B.n441 B.n440 163.367
R644 B.n441 B.n146 163.367
R645 B.n445 B.n146 163.367
R646 B.n446 B.n445 163.367
R647 B.n447 B.n446 163.367
R648 B.n447 B.n144 163.367
R649 B.n451 B.n144 163.367
R650 B.n452 B.n451 163.367
R651 B.n453 B.n452 163.367
R652 B.n453 B.n142 163.367
R653 B.n458 B.n457 163.367
R654 B.n459 B.n458 163.367
R655 B.n459 B.n140 163.367
R656 B.n463 B.n140 163.367
R657 B.n464 B.n463 163.367
R658 B.n465 B.n464 163.367
R659 B.n465 B.n138 163.367
R660 B.n469 B.n138 163.367
R661 B.n470 B.n469 163.367
R662 B.n471 B.n470 163.367
R663 B.n471 B.n136 163.367
R664 B.n475 B.n136 163.367
R665 B.n476 B.n475 163.367
R666 B.n477 B.n476 163.367
R667 B.n477 B.n134 163.367
R668 B.n481 B.n134 163.367
R669 B.n482 B.n481 163.367
R670 B.n483 B.n482 163.367
R671 B.n483 B.n132 163.367
R672 B.n487 B.n132 163.367
R673 B.n488 B.n487 163.367
R674 B.n489 B.n488 163.367
R675 B.n489 B.n130 163.367
R676 B.n493 B.n130 163.367
R677 B.n494 B.n493 163.367
R678 B.n495 B.n494 163.367
R679 B.n495 B.n128 163.367
R680 B.n499 B.n128 163.367
R681 B.n500 B.n499 163.367
R682 B.n501 B.n500 163.367
R683 B.n501 B.n126 163.367
R684 B.n505 B.n126 163.367
R685 B.n506 B.n505 163.367
R686 B.n507 B.n506 163.367
R687 B.n507 B.n124 163.367
R688 B.n511 B.n124 163.367
R689 B.n512 B.n511 163.367
R690 B.n513 B.n512 163.367
R691 B.n513 B.n122 163.367
R692 B.n517 B.n122 163.367
R693 B.n518 B.n517 163.367
R694 B.n519 B.n518 163.367
R695 B.n519 B.n120 163.367
R696 B.n523 B.n120 163.367
R697 B.n524 B.n523 163.367
R698 B.n525 B.n524 163.367
R699 B.n525 B.n118 163.367
R700 B.n529 B.n118 163.367
R701 B.n530 B.n529 163.367
R702 B.n531 B.n530 163.367
R703 B.n531 B.n116 163.367
R704 B.n535 B.n116 163.367
R705 B.n536 B.n535 163.367
R706 B.n537 B.n536 163.367
R707 B.n537 B.n114 163.367
R708 B.n541 B.n114 163.367
R709 B.n542 B.n541 163.367
R710 B.n543 B.n542 163.367
R711 B.n543 B.n112 163.367
R712 B.n547 B.n112 163.367
R713 B.n548 B.n547 163.367
R714 B.n549 B.n548 163.367
R715 B.n549 B.n110 163.367
R716 B.n553 B.n110 163.367
R717 B.n554 B.n553 163.367
R718 B.n555 B.n554 163.367
R719 B.n555 B.n108 163.367
R720 B.n559 B.n108 163.367
R721 B.n560 B.n559 163.367
R722 B.n561 B.n560 163.367
R723 B.n561 B.n106 163.367
R724 B.n565 B.n106 163.367
R725 B.n566 B.n565 163.367
R726 B.n567 B.n566 163.367
R727 B.n567 B.n104 163.367
R728 B.n571 B.n104 163.367
R729 B.n572 B.n571 163.367
R730 B.n573 B.n572 163.367
R731 B.n573 B.n102 163.367
R732 B.n577 B.n102 163.367
R733 B.n578 B.n577 163.367
R734 B.n579 B.n578 163.367
R735 B.n579 B.n100 163.367
R736 B.n583 B.n100 163.367
R737 B.n584 B.n583 163.367
R738 B.n585 B.n584 163.367
R739 B.n585 B.n98 163.367
R740 B.n589 B.n98 163.367
R741 B.n590 B.n589 163.367
R742 B.n591 B.n590 163.367
R743 B.n591 B.n96 163.367
R744 B.n595 B.n96 163.367
R745 B.n596 B.n595 163.367
R746 B.n597 B.n596 163.367
R747 B.n597 B.n94 163.367
R748 B.n601 B.n94 163.367
R749 B.n602 B.n601 163.367
R750 B.n603 B.n602 163.367
R751 B.n603 B.n92 163.367
R752 B.n607 B.n92 163.367
R753 B.n608 B.n607 163.367
R754 B.n609 B.n608 163.367
R755 B.n609 B.n90 163.367
R756 B.n613 B.n90 163.367
R757 B.n614 B.n613 163.367
R758 B.n615 B.n614 163.367
R759 B.n615 B.n88 163.367
R760 B.n619 B.n88 163.367
R761 B.n620 B.n619 163.367
R762 B.n621 B.n620 163.367
R763 B.n621 B.n86 163.367
R764 B.n625 B.n86 163.367
R765 B.n626 B.n625 163.367
R766 B.n627 B.n626 163.367
R767 B.n776 B.n31 163.367
R768 B.n772 B.n31 163.367
R769 B.n772 B.n771 163.367
R770 B.n771 B.n770 163.367
R771 B.n770 B.n33 163.367
R772 B.n766 B.n33 163.367
R773 B.n766 B.n765 163.367
R774 B.n765 B.n764 163.367
R775 B.n764 B.n35 163.367
R776 B.n760 B.n35 163.367
R777 B.n760 B.n759 163.367
R778 B.n759 B.n758 163.367
R779 B.n758 B.n37 163.367
R780 B.n754 B.n37 163.367
R781 B.n754 B.n753 163.367
R782 B.n753 B.n752 163.367
R783 B.n752 B.n39 163.367
R784 B.n748 B.n39 163.367
R785 B.n748 B.n747 163.367
R786 B.n747 B.n746 163.367
R787 B.n746 B.n41 163.367
R788 B.n742 B.n41 163.367
R789 B.n742 B.n741 163.367
R790 B.n741 B.n740 163.367
R791 B.n740 B.n43 163.367
R792 B.n736 B.n43 163.367
R793 B.n736 B.n735 163.367
R794 B.n735 B.n734 163.367
R795 B.n734 B.n45 163.367
R796 B.n730 B.n45 163.367
R797 B.n730 B.n729 163.367
R798 B.n729 B.n728 163.367
R799 B.n728 B.n47 163.367
R800 B.n724 B.n47 163.367
R801 B.n724 B.n723 163.367
R802 B.n723 B.n722 163.367
R803 B.n722 B.n49 163.367
R804 B.n718 B.n49 163.367
R805 B.n718 B.n717 163.367
R806 B.n717 B.n716 163.367
R807 B.n716 B.n51 163.367
R808 B.n712 B.n51 163.367
R809 B.n712 B.n711 163.367
R810 B.n711 B.n710 163.367
R811 B.n710 B.n53 163.367
R812 B.n706 B.n53 163.367
R813 B.n706 B.n705 163.367
R814 B.n705 B.n704 163.367
R815 B.n704 B.n58 163.367
R816 B.n700 B.n58 163.367
R817 B.n700 B.n699 163.367
R818 B.n699 B.n698 163.367
R819 B.n698 B.n60 163.367
R820 B.n693 B.n60 163.367
R821 B.n693 B.n692 163.367
R822 B.n692 B.n691 163.367
R823 B.n691 B.n64 163.367
R824 B.n687 B.n64 163.367
R825 B.n687 B.n686 163.367
R826 B.n686 B.n685 163.367
R827 B.n685 B.n66 163.367
R828 B.n681 B.n66 163.367
R829 B.n681 B.n680 163.367
R830 B.n680 B.n679 163.367
R831 B.n679 B.n68 163.367
R832 B.n675 B.n68 163.367
R833 B.n675 B.n674 163.367
R834 B.n674 B.n673 163.367
R835 B.n673 B.n70 163.367
R836 B.n669 B.n70 163.367
R837 B.n669 B.n668 163.367
R838 B.n668 B.n667 163.367
R839 B.n667 B.n72 163.367
R840 B.n663 B.n72 163.367
R841 B.n663 B.n662 163.367
R842 B.n662 B.n661 163.367
R843 B.n661 B.n74 163.367
R844 B.n657 B.n74 163.367
R845 B.n657 B.n656 163.367
R846 B.n656 B.n655 163.367
R847 B.n655 B.n76 163.367
R848 B.n651 B.n76 163.367
R849 B.n651 B.n650 163.367
R850 B.n650 B.n649 163.367
R851 B.n649 B.n78 163.367
R852 B.n645 B.n78 163.367
R853 B.n645 B.n644 163.367
R854 B.n644 B.n643 163.367
R855 B.n643 B.n80 163.367
R856 B.n639 B.n80 163.367
R857 B.n639 B.n638 163.367
R858 B.n638 B.n637 163.367
R859 B.n637 B.n82 163.367
R860 B.n633 B.n82 163.367
R861 B.n633 B.n632 163.367
R862 B.n632 B.n631 163.367
R863 B.n631 B.n84 163.367
R864 B.n166 B.n165 80.8732
R865 B.n172 B.n171 80.8732
R866 B.n55 B.n54 80.8732
R867 B.n62 B.n61 80.8732
R868 B.n389 B.n166 59.5399
R869 B.n173 B.n172 59.5399
R870 B.n56 B.n55 59.5399
R871 B.n695 B.n62 59.5399
R872 B.n775 B.n30 34.1859
R873 B.n629 B.n628 34.1859
R874 B.n456 B.n455 34.1859
R875 B.n306 B.n195 34.1859
R876 B B.n863 18.0485
R877 B.n775 B.n774 10.6151
R878 B.n774 B.n773 10.6151
R879 B.n773 B.n32 10.6151
R880 B.n769 B.n32 10.6151
R881 B.n769 B.n768 10.6151
R882 B.n768 B.n767 10.6151
R883 B.n767 B.n34 10.6151
R884 B.n763 B.n34 10.6151
R885 B.n763 B.n762 10.6151
R886 B.n762 B.n761 10.6151
R887 B.n761 B.n36 10.6151
R888 B.n757 B.n36 10.6151
R889 B.n757 B.n756 10.6151
R890 B.n756 B.n755 10.6151
R891 B.n755 B.n38 10.6151
R892 B.n751 B.n38 10.6151
R893 B.n751 B.n750 10.6151
R894 B.n750 B.n749 10.6151
R895 B.n749 B.n40 10.6151
R896 B.n745 B.n40 10.6151
R897 B.n745 B.n744 10.6151
R898 B.n744 B.n743 10.6151
R899 B.n743 B.n42 10.6151
R900 B.n739 B.n42 10.6151
R901 B.n739 B.n738 10.6151
R902 B.n738 B.n737 10.6151
R903 B.n737 B.n44 10.6151
R904 B.n733 B.n44 10.6151
R905 B.n733 B.n732 10.6151
R906 B.n732 B.n731 10.6151
R907 B.n731 B.n46 10.6151
R908 B.n727 B.n46 10.6151
R909 B.n727 B.n726 10.6151
R910 B.n726 B.n725 10.6151
R911 B.n725 B.n48 10.6151
R912 B.n721 B.n48 10.6151
R913 B.n721 B.n720 10.6151
R914 B.n720 B.n719 10.6151
R915 B.n719 B.n50 10.6151
R916 B.n715 B.n50 10.6151
R917 B.n715 B.n714 10.6151
R918 B.n714 B.n713 10.6151
R919 B.n713 B.n52 10.6151
R920 B.n709 B.n708 10.6151
R921 B.n708 B.n707 10.6151
R922 B.n707 B.n57 10.6151
R923 B.n703 B.n57 10.6151
R924 B.n703 B.n702 10.6151
R925 B.n702 B.n701 10.6151
R926 B.n701 B.n59 10.6151
R927 B.n697 B.n59 10.6151
R928 B.n697 B.n696 10.6151
R929 B.n694 B.n63 10.6151
R930 B.n690 B.n63 10.6151
R931 B.n690 B.n689 10.6151
R932 B.n689 B.n688 10.6151
R933 B.n688 B.n65 10.6151
R934 B.n684 B.n65 10.6151
R935 B.n684 B.n683 10.6151
R936 B.n683 B.n682 10.6151
R937 B.n682 B.n67 10.6151
R938 B.n678 B.n67 10.6151
R939 B.n678 B.n677 10.6151
R940 B.n677 B.n676 10.6151
R941 B.n676 B.n69 10.6151
R942 B.n672 B.n69 10.6151
R943 B.n672 B.n671 10.6151
R944 B.n671 B.n670 10.6151
R945 B.n670 B.n71 10.6151
R946 B.n666 B.n71 10.6151
R947 B.n666 B.n665 10.6151
R948 B.n665 B.n664 10.6151
R949 B.n664 B.n73 10.6151
R950 B.n660 B.n73 10.6151
R951 B.n660 B.n659 10.6151
R952 B.n659 B.n658 10.6151
R953 B.n658 B.n75 10.6151
R954 B.n654 B.n75 10.6151
R955 B.n654 B.n653 10.6151
R956 B.n653 B.n652 10.6151
R957 B.n652 B.n77 10.6151
R958 B.n648 B.n77 10.6151
R959 B.n648 B.n647 10.6151
R960 B.n647 B.n646 10.6151
R961 B.n646 B.n79 10.6151
R962 B.n642 B.n79 10.6151
R963 B.n642 B.n641 10.6151
R964 B.n641 B.n640 10.6151
R965 B.n640 B.n81 10.6151
R966 B.n636 B.n81 10.6151
R967 B.n636 B.n635 10.6151
R968 B.n635 B.n634 10.6151
R969 B.n634 B.n83 10.6151
R970 B.n630 B.n83 10.6151
R971 B.n630 B.n629 10.6151
R972 B.n456 B.n141 10.6151
R973 B.n460 B.n141 10.6151
R974 B.n461 B.n460 10.6151
R975 B.n462 B.n461 10.6151
R976 B.n462 B.n139 10.6151
R977 B.n466 B.n139 10.6151
R978 B.n467 B.n466 10.6151
R979 B.n468 B.n467 10.6151
R980 B.n468 B.n137 10.6151
R981 B.n472 B.n137 10.6151
R982 B.n473 B.n472 10.6151
R983 B.n474 B.n473 10.6151
R984 B.n474 B.n135 10.6151
R985 B.n478 B.n135 10.6151
R986 B.n479 B.n478 10.6151
R987 B.n480 B.n479 10.6151
R988 B.n480 B.n133 10.6151
R989 B.n484 B.n133 10.6151
R990 B.n485 B.n484 10.6151
R991 B.n486 B.n485 10.6151
R992 B.n486 B.n131 10.6151
R993 B.n490 B.n131 10.6151
R994 B.n491 B.n490 10.6151
R995 B.n492 B.n491 10.6151
R996 B.n492 B.n129 10.6151
R997 B.n496 B.n129 10.6151
R998 B.n497 B.n496 10.6151
R999 B.n498 B.n497 10.6151
R1000 B.n498 B.n127 10.6151
R1001 B.n502 B.n127 10.6151
R1002 B.n503 B.n502 10.6151
R1003 B.n504 B.n503 10.6151
R1004 B.n504 B.n125 10.6151
R1005 B.n508 B.n125 10.6151
R1006 B.n509 B.n508 10.6151
R1007 B.n510 B.n509 10.6151
R1008 B.n510 B.n123 10.6151
R1009 B.n514 B.n123 10.6151
R1010 B.n515 B.n514 10.6151
R1011 B.n516 B.n515 10.6151
R1012 B.n516 B.n121 10.6151
R1013 B.n520 B.n121 10.6151
R1014 B.n521 B.n520 10.6151
R1015 B.n522 B.n521 10.6151
R1016 B.n522 B.n119 10.6151
R1017 B.n526 B.n119 10.6151
R1018 B.n527 B.n526 10.6151
R1019 B.n528 B.n527 10.6151
R1020 B.n528 B.n117 10.6151
R1021 B.n532 B.n117 10.6151
R1022 B.n533 B.n532 10.6151
R1023 B.n534 B.n533 10.6151
R1024 B.n534 B.n115 10.6151
R1025 B.n538 B.n115 10.6151
R1026 B.n539 B.n538 10.6151
R1027 B.n540 B.n539 10.6151
R1028 B.n540 B.n113 10.6151
R1029 B.n544 B.n113 10.6151
R1030 B.n545 B.n544 10.6151
R1031 B.n546 B.n545 10.6151
R1032 B.n546 B.n111 10.6151
R1033 B.n550 B.n111 10.6151
R1034 B.n551 B.n550 10.6151
R1035 B.n552 B.n551 10.6151
R1036 B.n552 B.n109 10.6151
R1037 B.n556 B.n109 10.6151
R1038 B.n557 B.n556 10.6151
R1039 B.n558 B.n557 10.6151
R1040 B.n558 B.n107 10.6151
R1041 B.n562 B.n107 10.6151
R1042 B.n563 B.n562 10.6151
R1043 B.n564 B.n563 10.6151
R1044 B.n564 B.n105 10.6151
R1045 B.n568 B.n105 10.6151
R1046 B.n569 B.n568 10.6151
R1047 B.n570 B.n569 10.6151
R1048 B.n570 B.n103 10.6151
R1049 B.n574 B.n103 10.6151
R1050 B.n575 B.n574 10.6151
R1051 B.n576 B.n575 10.6151
R1052 B.n576 B.n101 10.6151
R1053 B.n580 B.n101 10.6151
R1054 B.n581 B.n580 10.6151
R1055 B.n582 B.n581 10.6151
R1056 B.n582 B.n99 10.6151
R1057 B.n586 B.n99 10.6151
R1058 B.n587 B.n586 10.6151
R1059 B.n588 B.n587 10.6151
R1060 B.n588 B.n97 10.6151
R1061 B.n592 B.n97 10.6151
R1062 B.n593 B.n592 10.6151
R1063 B.n594 B.n593 10.6151
R1064 B.n594 B.n95 10.6151
R1065 B.n598 B.n95 10.6151
R1066 B.n599 B.n598 10.6151
R1067 B.n600 B.n599 10.6151
R1068 B.n600 B.n93 10.6151
R1069 B.n604 B.n93 10.6151
R1070 B.n605 B.n604 10.6151
R1071 B.n606 B.n605 10.6151
R1072 B.n606 B.n91 10.6151
R1073 B.n610 B.n91 10.6151
R1074 B.n611 B.n610 10.6151
R1075 B.n612 B.n611 10.6151
R1076 B.n612 B.n89 10.6151
R1077 B.n616 B.n89 10.6151
R1078 B.n617 B.n616 10.6151
R1079 B.n618 B.n617 10.6151
R1080 B.n618 B.n87 10.6151
R1081 B.n622 B.n87 10.6151
R1082 B.n623 B.n622 10.6151
R1083 B.n624 B.n623 10.6151
R1084 B.n624 B.n85 10.6151
R1085 B.n628 B.n85 10.6151
R1086 B.n310 B.n195 10.6151
R1087 B.n311 B.n310 10.6151
R1088 B.n312 B.n311 10.6151
R1089 B.n312 B.n193 10.6151
R1090 B.n316 B.n193 10.6151
R1091 B.n317 B.n316 10.6151
R1092 B.n318 B.n317 10.6151
R1093 B.n318 B.n191 10.6151
R1094 B.n322 B.n191 10.6151
R1095 B.n323 B.n322 10.6151
R1096 B.n324 B.n323 10.6151
R1097 B.n324 B.n189 10.6151
R1098 B.n328 B.n189 10.6151
R1099 B.n329 B.n328 10.6151
R1100 B.n330 B.n329 10.6151
R1101 B.n330 B.n187 10.6151
R1102 B.n334 B.n187 10.6151
R1103 B.n335 B.n334 10.6151
R1104 B.n336 B.n335 10.6151
R1105 B.n336 B.n185 10.6151
R1106 B.n340 B.n185 10.6151
R1107 B.n341 B.n340 10.6151
R1108 B.n342 B.n341 10.6151
R1109 B.n342 B.n183 10.6151
R1110 B.n346 B.n183 10.6151
R1111 B.n347 B.n346 10.6151
R1112 B.n348 B.n347 10.6151
R1113 B.n348 B.n181 10.6151
R1114 B.n352 B.n181 10.6151
R1115 B.n353 B.n352 10.6151
R1116 B.n354 B.n353 10.6151
R1117 B.n354 B.n179 10.6151
R1118 B.n358 B.n179 10.6151
R1119 B.n359 B.n358 10.6151
R1120 B.n360 B.n359 10.6151
R1121 B.n360 B.n177 10.6151
R1122 B.n364 B.n177 10.6151
R1123 B.n365 B.n364 10.6151
R1124 B.n366 B.n365 10.6151
R1125 B.n366 B.n175 10.6151
R1126 B.n370 B.n175 10.6151
R1127 B.n371 B.n370 10.6151
R1128 B.n372 B.n371 10.6151
R1129 B.n376 B.n375 10.6151
R1130 B.n377 B.n376 10.6151
R1131 B.n377 B.n169 10.6151
R1132 B.n381 B.n169 10.6151
R1133 B.n382 B.n381 10.6151
R1134 B.n383 B.n382 10.6151
R1135 B.n383 B.n167 10.6151
R1136 B.n387 B.n167 10.6151
R1137 B.n388 B.n387 10.6151
R1138 B.n390 B.n163 10.6151
R1139 B.n394 B.n163 10.6151
R1140 B.n395 B.n394 10.6151
R1141 B.n396 B.n395 10.6151
R1142 B.n396 B.n161 10.6151
R1143 B.n400 B.n161 10.6151
R1144 B.n401 B.n400 10.6151
R1145 B.n402 B.n401 10.6151
R1146 B.n402 B.n159 10.6151
R1147 B.n406 B.n159 10.6151
R1148 B.n407 B.n406 10.6151
R1149 B.n408 B.n407 10.6151
R1150 B.n408 B.n157 10.6151
R1151 B.n412 B.n157 10.6151
R1152 B.n413 B.n412 10.6151
R1153 B.n414 B.n413 10.6151
R1154 B.n414 B.n155 10.6151
R1155 B.n418 B.n155 10.6151
R1156 B.n419 B.n418 10.6151
R1157 B.n420 B.n419 10.6151
R1158 B.n420 B.n153 10.6151
R1159 B.n424 B.n153 10.6151
R1160 B.n425 B.n424 10.6151
R1161 B.n426 B.n425 10.6151
R1162 B.n426 B.n151 10.6151
R1163 B.n430 B.n151 10.6151
R1164 B.n431 B.n430 10.6151
R1165 B.n432 B.n431 10.6151
R1166 B.n432 B.n149 10.6151
R1167 B.n436 B.n149 10.6151
R1168 B.n437 B.n436 10.6151
R1169 B.n438 B.n437 10.6151
R1170 B.n438 B.n147 10.6151
R1171 B.n442 B.n147 10.6151
R1172 B.n443 B.n442 10.6151
R1173 B.n444 B.n443 10.6151
R1174 B.n444 B.n145 10.6151
R1175 B.n448 B.n145 10.6151
R1176 B.n449 B.n448 10.6151
R1177 B.n450 B.n449 10.6151
R1178 B.n450 B.n143 10.6151
R1179 B.n454 B.n143 10.6151
R1180 B.n455 B.n454 10.6151
R1181 B.n306 B.n305 10.6151
R1182 B.n305 B.n304 10.6151
R1183 B.n304 B.n197 10.6151
R1184 B.n300 B.n197 10.6151
R1185 B.n300 B.n299 10.6151
R1186 B.n299 B.n298 10.6151
R1187 B.n298 B.n199 10.6151
R1188 B.n294 B.n199 10.6151
R1189 B.n294 B.n293 10.6151
R1190 B.n293 B.n292 10.6151
R1191 B.n292 B.n201 10.6151
R1192 B.n288 B.n201 10.6151
R1193 B.n288 B.n287 10.6151
R1194 B.n287 B.n286 10.6151
R1195 B.n286 B.n203 10.6151
R1196 B.n282 B.n203 10.6151
R1197 B.n282 B.n281 10.6151
R1198 B.n281 B.n280 10.6151
R1199 B.n280 B.n205 10.6151
R1200 B.n276 B.n205 10.6151
R1201 B.n276 B.n275 10.6151
R1202 B.n275 B.n274 10.6151
R1203 B.n274 B.n207 10.6151
R1204 B.n270 B.n207 10.6151
R1205 B.n270 B.n269 10.6151
R1206 B.n269 B.n268 10.6151
R1207 B.n268 B.n209 10.6151
R1208 B.n264 B.n209 10.6151
R1209 B.n264 B.n263 10.6151
R1210 B.n263 B.n262 10.6151
R1211 B.n262 B.n211 10.6151
R1212 B.n258 B.n211 10.6151
R1213 B.n258 B.n257 10.6151
R1214 B.n257 B.n256 10.6151
R1215 B.n256 B.n213 10.6151
R1216 B.n252 B.n213 10.6151
R1217 B.n252 B.n251 10.6151
R1218 B.n251 B.n250 10.6151
R1219 B.n250 B.n215 10.6151
R1220 B.n246 B.n215 10.6151
R1221 B.n246 B.n245 10.6151
R1222 B.n245 B.n244 10.6151
R1223 B.n244 B.n217 10.6151
R1224 B.n240 B.n217 10.6151
R1225 B.n240 B.n239 10.6151
R1226 B.n239 B.n238 10.6151
R1227 B.n238 B.n219 10.6151
R1228 B.n234 B.n219 10.6151
R1229 B.n234 B.n233 10.6151
R1230 B.n233 B.n232 10.6151
R1231 B.n232 B.n221 10.6151
R1232 B.n228 B.n221 10.6151
R1233 B.n228 B.n227 10.6151
R1234 B.n227 B.n226 10.6151
R1235 B.n226 B.n223 10.6151
R1236 B.n223 B.n0 10.6151
R1237 B.n859 B.n1 10.6151
R1238 B.n859 B.n858 10.6151
R1239 B.n858 B.n857 10.6151
R1240 B.n857 B.n4 10.6151
R1241 B.n853 B.n4 10.6151
R1242 B.n853 B.n852 10.6151
R1243 B.n852 B.n851 10.6151
R1244 B.n851 B.n6 10.6151
R1245 B.n847 B.n6 10.6151
R1246 B.n847 B.n846 10.6151
R1247 B.n846 B.n845 10.6151
R1248 B.n845 B.n8 10.6151
R1249 B.n841 B.n8 10.6151
R1250 B.n841 B.n840 10.6151
R1251 B.n840 B.n839 10.6151
R1252 B.n839 B.n10 10.6151
R1253 B.n835 B.n10 10.6151
R1254 B.n835 B.n834 10.6151
R1255 B.n834 B.n833 10.6151
R1256 B.n833 B.n12 10.6151
R1257 B.n829 B.n12 10.6151
R1258 B.n829 B.n828 10.6151
R1259 B.n828 B.n827 10.6151
R1260 B.n827 B.n14 10.6151
R1261 B.n823 B.n14 10.6151
R1262 B.n823 B.n822 10.6151
R1263 B.n822 B.n821 10.6151
R1264 B.n821 B.n16 10.6151
R1265 B.n817 B.n16 10.6151
R1266 B.n817 B.n816 10.6151
R1267 B.n816 B.n815 10.6151
R1268 B.n815 B.n18 10.6151
R1269 B.n811 B.n18 10.6151
R1270 B.n811 B.n810 10.6151
R1271 B.n810 B.n809 10.6151
R1272 B.n809 B.n20 10.6151
R1273 B.n805 B.n20 10.6151
R1274 B.n805 B.n804 10.6151
R1275 B.n804 B.n803 10.6151
R1276 B.n803 B.n22 10.6151
R1277 B.n799 B.n22 10.6151
R1278 B.n799 B.n798 10.6151
R1279 B.n798 B.n797 10.6151
R1280 B.n797 B.n24 10.6151
R1281 B.n793 B.n24 10.6151
R1282 B.n793 B.n792 10.6151
R1283 B.n792 B.n791 10.6151
R1284 B.n791 B.n26 10.6151
R1285 B.n787 B.n26 10.6151
R1286 B.n787 B.n786 10.6151
R1287 B.n786 B.n785 10.6151
R1288 B.n785 B.n28 10.6151
R1289 B.n781 B.n28 10.6151
R1290 B.n781 B.n780 10.6151
R1291 B.n780 B.n779 10.6151
R1292 B.n779 B.n30 10.6151
R1293 B.n56 B.n52 9.36635
R1294 B.n695 B.n694 9.36635
R1295 B.n372 B.n173 9.36635
R1296 B.n390 B.n389 9.36635
R1297 B.n863 B.n0 2.81026
R1298 B.n863 B.n1 2.81026
R1299 B.n709 B.n56 1.24928
R1300 B.n696 B.n695 1.24928
R1301 B.n375 B.n173 1.24928
R1302 B.n389 B.n388 1.24928
R1303 VP.n15 VP.n14 161.3
R1304 VP.n16 VP.n11 161.3
R1305 VP.n18 VP.n17 161.3
R1306 VP.n19 VP.n10 161.3
R1307 VP.n21 VP.n20 161.3
R1308 VP.n22 VP.n9 161.3
R1309 VP.n24 VP.n23 161.3
R1310 VP.n25 VP.n8 161.3
R1311 VP.n54 VP.n0 161.3
R1312 VP.n53 VP.n52 161.3
R1313 VP.n51 VP.n1 161.3
R1314 VP.n50 VP.n49 161.3
R1315 VP.n48 VP.n2 161.3
R1316 VP.n47 VP.n46 161.3
R1317 VP.n45 VP.n3 161.3
R1318 VP.n44 VP.n43 161.3
R1319 VP.n41 VP.n4 161.3
R1320 VP.n40 VP.n39 161.3
R1321 VP.n38 VP.n5 161.3
R1322 VP.n37 VP.n36 161.3
R1323 VP.n35 VP.n6 161.3
R1324 VP.n34 VP.n33 161.3
R1325 VP.n32 VP.n7 161.3
R1326 VP.n31 VP.n30 161.3
R1327 VP.n12 VP.t2 113.004
R1328 VP.n29 VP.t5 80.8359
R1329 VP.n42 VP.t3 80.8359
R1330 VP.n55 VP.t1 80.8359
R1331 VP.n26 VP.t0 80.8359
R1332 VP.n13 VP.t4 80.8359
R1333 VP.n13 VP.n12 62.6769
R1334 VP.n29 VP.n28 61.5371
R1335 VP.n56 VP.n55 61.5371
R1336 VP.n27 VP.n26 61.5371
R1337 VP.n36 VP.n35 56.4773
R1338 VP.n49 VP.n48 56.4773
R1339 VP.n20 VP.n19 56.4773
R1340 VP.n28 VP.n27 54.4164
R1341 VP.n30 VP.n7 24.3439
R1342 VP.n34 VP.n7 24.3439
R1343 VP.n35 VP.n34 24.3439
R1344 VP.n36 VP.n5 24.3439
R1345 VP.n40 VP.n5 24.3439
R1346 VP.n41 VP.n40 24.3439
R1347 VP.n43 VP.n3 24.3439
R1348 VP.n47 VP.n3 24.3439
R1349 VP.n48 VP.n47 24.3439
R1350 VP.n49 VP.n1 24.3439
R1351 VP.n53 VP.n1 24.3439
R1352 VP.n54 VP.n53 24.3439
R1353 VP.n20 VP.n9 24.3439
R1354 VP.n24 VP.n9 24.3439
R1355 VP.n25 VP.n24 24.3439
R1356 VP.n14 VP.n11 24.3439
R1357 VP.n18 VP.n11 24.3439
R1358 VP.n19 VP.n18 24.3439
R1359 VP.n30 VP.n29 20.449
R1360 VP.n55 VP.n54 20.449
R1361 VP.n26 VP.n25 20.449
R1362 VP.n42 VP.n41 12.1722
R1363 VP.n43 VP.n42 12.1722
R1364 VP.n14 VP.n13 12.1722
R1365 VP.n15 VP.n12 2.68622
R1366 VP.n27 VP.n8 0.417764
R1367 VP.n31 VP.n28 0.417764
R1368 VP.n56 VP.n0 0.417764
R1369 VP VP.n56 0.394061
R1370 VP.n16 VP.n15 0.189894
R1371 VP.n17 VP.n16 0.189894
R1372 VP.n17 VP.n10 0.189894
R1373 VP.n21 VP.n10 0.189894
R1374 VP.n22 VP.n21 0.189894
R1375 VP.n23 VP.n22 0.189894
R1376 VP.n23 VP.n8 0.189894
R1377 VP.n32 VP.n31 0.189894
R1378 VP.n33 VP.n32 0.189894
R1379 VP.n33 VP.n6 0.189894
R1380 VP.n37 VP.n6 0.189894
R1381 VP.n38 VP.n37 0.189894
R1382 VP.n39 VP.n38 0.189894
R1383 VP.n39 VP.n4 0.189894
R1384 VP.n44 VP.n4 0.189894
R1385 VP.n45 VP.n44 0.189894
R1386 VP.n46 VP.n45 0.189894
R1387 VP.n46 VP.n2 0.189894
R1388 VP.n50 VP.n2 0.189894
R1389 VP.n51 VP.n50 0.189894
R1390 VP.n52 VP.n51 0.189894
R1391 VP.n52 VP.n0 0.189894
R1392 VTAIL.n282 VTAIL.n218 756.745
R1393 VTAIL.n66 VTAIL.n2 756.745
R1394 VTAIL.n212 VTAIL.n148 756.745
R1395 VTAIL.n140 VTAIL.n76 756.745
R1396 VTAIL.n241 VTAIL.n240 585
R1397 VTAIL.n238 VTAIL.n237 585
R1398 VTAIL.n247 VTAIL.n246 585
R1399 VTAIL.n249 VTAIL.n248 585
R1400 VTAIL.n234 VTAIL.n233 585
R1401 VTAIL.n255 VTAIL.n254 585
R1402 VTAIL.n258 VTAIL.n257 585
R1403 VTAIL.n256 VTAIL.n230 585
R1404 VTAIL.n263 VTAIL.n229 585
R1405 VTAIL.n265 VTAIL.n264 585
R1406 VTAIL.n267 VTAIL.n266 585
R1407 VTAIL.n226 VTAIL.n225 585
R1408 VTAIL.n273 VTAIL.n272 585
R1409 VTAIL.n275 VTAIL.n274 585
R1410 VTAIL.n222 VTAIL.n221 585
R1411 VTAIL.n281 VTAIL.n280 585
R1412 VTAIL.n283 VTAIL.n282 585
R1413 VTAIL.n25 VTAIL.n24 585
R1414 VTAIL.n22 VTAIL.n21 585
R1415 VTAIL.n31 VTAIL.n30 585
R1416 VTAIL.n33 VTAIL.n32 585
R1417 VTAIL.n18 VTAIL.n17 585
R1418 VTAIL.n39 VTAIL.n38 585
R1419 VTAIL.n42 VTAIL.n41 585
R1420 VTAIL.n40 VTAIL.n14 585
R1421 VTAIL.n47 VTAIL.n13 585
R1422 VTAIL.n49 VTAIL.n48 585
R1423 VTAIL.n51 VTAIL.n50 585
R1424 VTAIL.n10 VTAIL.n9 585
R1425 VTAIL.n57 VTAIL.n56 585
R1426 VTAIL.n59 VTAIL.n58 585
R1427 VTAIL.n6 VTAIL.n5 585
R1428 VTAIL.n65 VTAIL.n64 585
R1429 VTAIL.n67 VTAIL.n66 585
R1430 VTAIL.n213 VTAIL.n212 585
R1431 VTAIL.n211 VTAIL.n210 585
R1432 VTAIL.n152 VTAIL.n151 585
R1433 VTAIL.n205 VTAIL.n204 585
R1434 VTAIL.n203 VTAIL.n202 585
R1435 VTAIL.n156 VTAIL.n155 585
R1436 VTAIL.n197 VTAIL.n196 585
R1437 VTAIL.n195 VTAIL.n194 585
R1438 VTAIL.n193 VTAIL.n159 585
R1439 VTAIL.n163 VTAIL.n160 585
R1440 VTAIL.n188 VTAIL.n187 585
R1441 VTAIL.n186 VTAIL.n185 585
R1442 VTAIL.n165 VTAIL.n164 585
R1443 VTAIL.n180 VTAIL.n179 585
R1444 VTAIL.n178 VTAIL.n177 585
R1445 VTAIL.n169 VTAIL.n168 585
R1446 VTAIL.n172 VTAIL.n171 585
R1447 VTAIL.n141 VTAIL.n140 585
R1448 VTAIL.n139 VTAIL.n138 585
R1449 VTAIL.n80 VTAIL.n79 585
R1450 VTAIL.n133 VTAIL.n132 585
R1451 VTAIL.n131 VTAIL.n130 585
R1452 VTAIL.n84 VTAIL.n83 585
R1453 VTAIL.n125 VTAIL.n124 585
R1454 VTAIL.n123 VTAIL.n122 585
R1455 VTAIL.n121 VTAIL.n87 585
R1456 VTAIL.n91 VTAIL.n88 585
R1457 VTAIL.n116 VTAIL.n115 585
R1458 VTAIL.n114 VTAIL.n113 585
R1459 VTAIL.n93 VTAIL.n92 585
R1460 VTAIL.n108 VTAIL.n107 585
R1461 VTAIL.n106 VTAIL.n105 585
R1462 VTAIL.n97 VTAIL.n96 585
R1463 VTAIL.n100 VTAIL.n99 585
R1464 VTAIL.t4 VTAIL.n239 329.036
R1465 VTAIL.t9 VTAIL.n23 329.036
R1466 VTAIL.t7 VTAIL.n170 329.036
R1467 VTAIL.t3 VTAIL.n98 329.036
R1468 VTAIL.n240 VTAIL.n237 171.744
R1469 VTAIL.n247 VTAIL.n237 171.744
R1470 VTAIL.n248 VTAIL.n247 171.744
R1471 VTAIL.n248 VTAIL.n233 171.744
R1472 VTAIL.n255 VTAIL.n233 171.744
R1473 VTAIL.n257 VTAIL.n255 171.744
R1474 VTAIL.n257 VTAIL.n256 171.744
R1475 VTAIL.n256 VTAIL.n229 171.744
R1476 VTAIL.n265 VTAIL.n229 171.744
R1477 VTAIL.n266 VTAIL.n265 171.744
R1478 VTAIL.n266 VTAIL.n225 171.744
R1479 VTAIL.n273 VTAIL.n225 171.744
R1480 VTAIL.n274 VTAIL.n273 171.744
R1481 VTAIL.n274 VTAIL.n221 171.744
R1482 VTAIL.n281 VTAIL.n221 171.744
R1483 VTAIL.n282 VTAIL.n281 171.744
R1484 VTAIL.n24 VTAIL.n21 171.744
R1485 VTAIL.n31 VTAIL.n21 171.744
R1486 VTAIL.n32 VTAIL.n31 171.744
R1487 VTAIL.n32 VTAIL.n17 171.744
R1488 VTAIL.n39 VTAIL.n17 171.744
R1489 VTAIL.n41 VTAIL.n39 171.744
R1490 VTAIL.n41 VTAIL.n40 171.744
R1491 VTAIL.n40 VTAIL.n13 171.744
R1492 VTAIL.n49 VTAIL.n13 171.744
R1493 VTAIL.n50 VTAIL.n49 171.744
R1494 VTAIL.n50 VTAIL.n9 171.744
R1495 VTAIL.n57 VTAIL.n9 171.744
R1496 VTAIL.n58 VTAIL.n57 171.744
R1497 VTAIL.n58 VTAIL.n5 171.744
R1498 VTAIL.n65 VTAIL.n5 171.744
R1499 VTAIL.n66 VTAIL.n65 171.744
R1500 VTAIL.n212 VTAIL.n211 171.744
R1501 VTAIL.n211 VTAIL.n151 171.744
R1502 VTAIL.n204 VTAIL.n151 171.744
R1503 VTAIL.n204 VTAIL.n203 171.744
R1504 VTAIL.n203 VTAIL.n155 171.744
R1505 VTAIL.n196 VTAIL.n155 171.744
R1506 VTAIL.n196 VTAIL.n195 171.744
R1507 VTAIL.n195 VTAIL.n159 171.744
R1508 VTAIL.n163 VTAIL.n159 171.744
R1509 VTAIL.n187 VTAIL.n163 171.744
R1510 VTAIL.n187 VTAIL.n186 171.744
R1511 VTAIL.n186 VTAIL.n164 171.744
R1512 VTAIL.n179 VTAIL.n164 171.744
R1513 VTAIL.n179 VTAIL.n178 171.744
R1514 VTAIL.n178 VTAIL.n168 171.744
R1515 VTAIL.n171 VTAIL.n168 171.744
R1516 VTAIL.n140 VTAIL.n139 171.744
R1517 VTAIL.n139 VTAIL.n79 171.744
R1518 VTAIL.n132 VTAIL.n79 171.744
R1519 VTAIL.n132 VTAIL.n131 171.744
R1520 VTAIL.n131 VTAIL.n83 171.744
R1521 VTAIL.n124 VTAIL.n83 171.744
R1522 VTAIL.n124 VTAIL.n123 171.744
R1523 VTAIL.n123 VTAIL.n87 171.744
R1524 VTAIL.n91 VTAIL.n87 171.744
R1525 VTAIL.n115 VTAIL.n91 171.744
R1526 VTAIL.n115 VTAIL.n114 171.744
R1527 VTAIL.n114 VTAIL.n92 171.744
R1528 VTAIL.n107 VTAIL.n92 171.744
R1529 VTAIL.n107 VTAIL.n106 171.744
R1530 VTAIL.n106 VTAIL.n96 171.744
R1531 VTAIL.n99 VTAIL.n96 171.744
R1532 VTAIL.n240 VTAIL.t4 85.8723
R1533 VTAIL.n24 VTAIL.t9 85.8723
R1534 VTAIL.n171 VTAIL.t7 85.8723
R1535 VTAIL.n99 VTAIL.t3 85.8723
R1536 VTAIL.n1 VTAIL.n0 57.1083
R1537 VTAIL.n73 VTAIL.n72 57.1083
R1538 VTAIL.n147 VTAIL.n146 57.1083
R1539 VTAIL.n75 VTAIL.n74 57.1083
R1540 VTAIL.n287 VTAIL.n286 32.9611
R1541 VTAIL.n71 VTAIL.n70 32.9611
R1542 VTAIL.n217 VTAIL.n216 32.9611
R1543 VTAIL.n145 VTAIL.n144 32.9611
R1544 VTAIL.n75 VTAIL.n73 30.66
R1545 VTAIL.n287 VTAIL.n217 27.0652
R1546 VTAIL.n264 VTAIL.n263 13.1884
R1547 VTAIL.n48 VTAIL.n47 13.1884
R1548 VTAIL.n194 VTAIL.n193 13.1884
R1549 VTAIL.n122 VTAIL.n121 13.1884
R1550 VTAIL.n262 VTAIL.n230 12.8005
R1551 VTAIL.n267 VTAIL.n228 12.8005
R1552 VTAIL.n46 VTAIL.n14 12.8005
R1553 VTAIL.n51 VTAIL.n12 12.8005
R1554 VTAIL.n197 VTAIL.n158 12.8005
R1555 VTAIL.n192 VTAIL.n160 12.8005
R1556 VTAIL.n125 VTAIL.n86 12.8005
R1557 VTAIL.n120 VTAIL.n88 12.8005
R1558 VTAIL.n259 VTAIL.n258 12.0247
R1559 VTAIL.n268 VTAIL.n226 12.0247
R1560 VTAIL.n43 VTAIL.n42 12.0247
R1561 VTAIL.n52 VTAIL.n10 12.0247
R1562 VTAIL.n198 VTAIL.n156 12.0247
R1563 VTAIL.n189 VTAIL.n188 12.0247
R1564 VTAIL.n126 VTAIL.n84 12.0247
R1565 VTAIL.n117 VTAIL.n116 12.0247
R1566 VTAIL.n254 VTAIL.n232 11.249
R1567 VTAIL.n272 VTAIL.n271 11.249
R1568 VTAIL.n38 VTAIL.n16 11.249
R1569 VTAIL.n56 VTAIL.n55 11.249
R1570 VTAIL.n202 VTAIL.n201 11.249
R1571 VTAIL.n185 VTAIL.n162 11.249
R1572 VTAIL.n130 VTAIL.n129 11.249
R1573 VTAIL.n113 VTAIL.n90 11.249
R1574 VTAIL.n241 VTAIL.n239 10.7239
R1575 VTAIL.n25 VTAIL.n23 10.7239
R1576 VTAIL.n172 VTAIL.n170 10.7239
R1577 VTAIL.n100 VTAIL.n98 10.7239
R1578 VTAIL.n253 VTAIL.n234 10.4732
R1579 VTAIL.n275 VTAIL.n224 10.4732
R1580 VTAIL.n37 VTAIL.n18 10.4732
R1581 VTAIL.n59 VTAIL.n8 10.4732
R1582 VTAIL.n205 VTAIL.n154 10.4732
R1583 VTAIL.n184 VTAIL.n165 10.4732
R1584 VTAIL.n133 VTAIL.n82 10.4732
R1585 VTAIL.n112 VTAIL.n93 10.4732
R1586 VTAIL.n250 VTAIL.n249 9.69747
R1587 VTAIL.n276 VTAIL.n222 9.69747
R1588 VTAIL.n34 VTAIL.n33 9.69747
R1589 VTAIL.n60 VTAIL.n6 9.69747
R1590 VTAIL.n206 VTAIL.n152 9.69747
R1591 VTAIL.n181 VTAIL.n180 9.69747
R1592 VTAIL.n134 VTAIL.n80 9.69747
R1593 VTAIL.n109 VTAIL.n108 9.69747
R1594 VTAIL.n286 VTAIL.n285 9.45567
R1595 VTAIL.n70 VTAIL.n69 9.45567
R1596 VTAIL.n216 VTAIL.n215 9.45567
R1597 VTAIL.n144 VTAIL.n143 9.45567
R1598 VTAIL.n220 VTAIL.n219 9.3005
R1599 VTAIL.n279 VTAIL.n278 9.3005
R1600 VTAIL.n277 VTAIL.n276 9.3005
R1601 VTAIL.n224 VTAIL.n223 9.3005
R1602 VTAIL.n271 VTAIL.n270 9.3005
R1603 VTAIL.n269 VTAIL.n268 9.3005
R1604 VTAIL.n228 VTAIL.n227 9.3005
R1605 VTAIL.n243 VTAIL.n242 9.3005
R1606 VTAIL.n245 VTAIL.n244 9.3005
R1607 VTAIL.n236 VTAIL.n235 9.3005
R1608 VTAIL.n251 VTAIL.n250 9.3005
R1609 VTAIL.n253 VTAIL.n252 9.3005
R1610 VTAIL.n232 VTAIL.n231 9.3005
R1611 VTAIL.n260 VTAIL.n259 9.3005
R1612 VTAIL.n262 VTAIL.n261 9.3005
R1613 VTAIL.n285 VTAIL.n284 9.3005
R1614 VTAIL.n4 VTAIL.n3 9.3005
R1615 VTAIL.n63 VTAIL.n62 9.3005
R1616 VTAIL.n61 VTAIL.n60 9.3005
R1617 VTAIL.n8 VTAIL.n7 9.3005
R1618 VTAIL.n55 VTAIL.n54 9.3005
R1619 VTAIL.n53 VTAIL.n52 9.3005
R1620 VTAIL.n12 VTAIL.n11 9.3005
R1621 VTAIL.n27 VTAIL.n26 9.3005
R1622 VTAIL.n29 VTAIL.n28 9.3005
R1623 VTAIL.n20 VTAIL.n19 9.3005
R1624 VTAIL.n35 VTAIL.n34 9.3005
R1625 VTAIL.n37 VTAIL.n36 9.3005
R1626 VTAIL.n16 VTAIL.n15 9.3005
R1627 VTAIL.n44 VTAIL.n43 9.3005
R1628 VTAIL.n46 VTAIL.n45 9.3005
R1629 VTAIL.n69 VTAIL.n68 9.3005
R1630 VTAIL.n174 VTAIL.n173 9.3005
R1631 VTAIL.n176 VTAIL.n175 9.3005
R1632 VTAIL.n167 VTAIL.n166 9.3005
R1633 VTAIL.n182 VTAIL.n181 9.3005
R1634 VTAIL.n184 VTAIL.n183 9.3005
R1635 VTAIL.n162 VTAIL.n161 9.3005
R1636 VTAIL.n190 VTAIL.n189 9.3005
R1637 VTAIL.n192 VTAIL.n191 9.3005
R1638 VTAIL.n215 VTAIL.n214 9.3005
R1639 VTAIL.n150 VTAIL.n149 9.3005
R1640 VTAIL.n209 VTAIL.n208 9.3005
R1641 VTAIL.n207 VTAIL.n206 9.3005
R1642 VTAIL.n154 VTAIL.n153 9.3005
R1643 VTAIL.n201 VTAIL.n200 9.3005
R1644 VTAIL.n199 VTAIL.n198 9.3005
R1645 VTAIL.n158 VTAIL.n157 9.3005
R1646 VTAIL.n102 VTAIL.n101 9.3005
R1647 VTAIL.n104 VTAIL.n103 9.3005
R1648 VTAIL.n95 VTAIL.n94 9.3005
R1649 VTAIL.n110 VTAIL.n109 9.3005
R1650 VTAIL.n112 VTAIL.n111 9.3005
R1651 VTAIL.n90 VTAIL.n89 9.3005
R1652 VTAIL.n118 VTAIL.n117 9.3005
R1653 VTAIL.n120 VTAIL.n119 9.3005
R1654 VTAIL.n143 VTAIL.n142 9.3005
R1655 VTAIL.n78 VTAIL.n77 9.3005
R1656 VTAIL.n137 VTAIL.n136 9.3005
R1657 VTAIL.n135 VTAIL.n134 9.3005
R1658 VTAIL.n82 VTAIL.n81 9.3005
R1659 VTAIL.n129 VTAIL.n128 9.3005
R1660 VTAIL.n127 VTAIL.n126 9.3005
R1661 VTAIL.n86 VTAIL.n85 9.3005
R1662 VTAIL.n246 VTAIL.n236 8.92171
R1663 VTAIL.n280 VTAIL.n279 8.92171
R1664 VTAIL.n30 VTAIL.n20 8.92171
R1665 VTAIL.n64 VTAIL.n63 8.92171
R1666 VTAIL.n210 VTAIL.n209 8.92171
R1667 VTAIL.n177 VTAIL.n167 8.92171
R1668 VTAIL.n138 VTAIL.n137 8.92171
R1669 VTAIL.n105 VTAIL.n95 8.92171
R1670 VTAIL.n245 VTAIL.n238 8.14595
R1671 VTAIL.n283 VTAIL.n220 8.14595
R1672 VTAIL.n29 VTAIL.n22 8.14595
R1673 VTAIL.n67 VTAIL.n4 8.14595
R1674 VTAIL.n213 VTAIL.n150 8.14595
R1675 VTAIL.n176 VTAIL.n169 8.14595
R1676 VTAIL.n141 VTAIL.n78 8.14595
R1677 VTAIL.n104 VTAIL.n97 8.14595
R1678 VTAIL.n242 VTAIL.n241 7.3702
R1679 VTAIL.n284 VTAIL.n218 7.3702
R1680 VTAIL.n26 VTAIL.n25 7.3702
R1681 VTAIL.n68 VTAIL.n2 7.3702
R1682 VTAIL.n214 VTAIL.n148 7.3702
R1683 VTAIL.n173 VTAIL.n172 7.3702
R1684 VTAIL.n142 VTAIL.n76 7.3702
R1685 VTAIL.n101 VTAIL.n100 7.3702
R1686 VTAIL.n286 VTAIL.n218 6.59444
R1687 VTAIL.n70 VTAIL.n2 6.59444
R1688 VTAIL.n216 VTAIL.n148 6.59444
R1689 VTAIL.n144 VTAIL.n76 6.59444
R1690 VTAIL.n242 VTAIL.n238 5.81868
R1691 VTAIL.n284 VTAIL.n283 5.81868
R1692 VTAIL.n26 VTAIL.n22 5.81868
R1693 VTAIL.n68 VTAIL.n67 5.81868
R1694 VTAIL.n214 VTAIL.n213 5.81868
R1695 VTAIL.n173 VTAIL.n169 5.81868
R1696 VTAIL.n142 VTAIL.n141 5.81868
R1697 VTAIL.n101 VTAIL.n97 5.81868
R1698 VTAIL.n246 VTAIL.n245 5.04292
R1699 VTAIL.n280 VTAIL.n220 5.04292
R1700 VTAIL.n30 VTAIL.n29 5.04292
R1701 VTAIL.n64 VTAIL.n4 5.04292
R1702 VTAIL.n210 VTAIL.n150 5.04292
R1703 VTAIL.n177 VTAIL.n176 5.04292
R1704 VTAIL.n138 VTAIL.n78 5.04292
R1705 VTAIL.n105 VTAIL.n104 5.04292
R1706 VTAIL.n249 VTAIL.n236 4.26717
R1707 VTAIL.n279 VTAIL.n222 4.26717
R1708 VTAIL.n33 VTAIL.n20 4.26717
R1709 VTAIL.n63 VTAIL.n6 4.26717
R1710 VTAIL.n209 VTAIL.n152 4.26717
R1711 VTAIL.n180 VTAIL.n167 4.26717
R1712 VTAIL.n137 VTAIL.n80 4.26717
R1713 VTAIL.n108 VTAIL.n95 4.26717
R1714 VTAIL.n145 VTAIL.n75 3.59533
R1715 VTAIL.n217 VTAIL.n147 3.59533
R1716 VTAIL.n73 VTAIL.n71 3.59533
R1717 VTAIL.n250 VTAIL.n234 3.49141
R1718 VTAIL.n276 VTAIL.n275 3.49141
R1719 VTAIL.n34 VTAIL.n18 3.49141
R1720 VTAIL.n60 VTAIL.n59 3.49141
R1721 VTAIL.n206 VTAIL.n205 3.49141
R1722 VTAIL.n181 VTAIL.n165 3.49141
R1723 VTAIL.n134 VTAIL.n133 3.49141
R1724 VTAIL.n109 VTAIL.n93 3.49141
R1725 VTAIL.n254 VTAIL.n253 2.71565
R1726 VTAIL.n272 VTAIL.n224 2.71565
R1727 VTAIL.n38 VTAIL.n37 2.71565
R1728 VTAIL.n56 VTAIL.n8 2.71565
R1729 VTAIL.n202 VTAIL.n154 2.71565
R1730 VTAIL.n185 VTAIL.n184 2.71565
R1731 VTAIL.n130 VTAIL.n82 2.71565
R1732 VTAIL.n113 VTAIL.n112 2.71565
R1733 VTAIL VTAIL.n287 2.63843
R1734 VTAIL.n0 VTAIL.t1 2.52418
R1735 VTAIL.n0 VTAIL.t0 2.52418
R1736 VTAIL.n72 VTAIL.t11 2.52418
R1737 VTAIL.n72 VTAIL.t8 2.52418
R1738 VTAIL.n146 VTAIL.t10 2.52418
R1739 VTAIL.n146 VTAIL.t6 2.52418
R1740 VTAIL.n74 VTAIL.t5 2.52418
R1741 VTAIL.n74 VTAIL.t2 2.52418
R1742 VTAIL.n243 VTAIL.n239 2.41282
R1743 VTAIL.n27 VTAIL.n23 2.41282
R1744 VTAIL.n174 VTAIL.n170 2.41282
R1745 VTAIL.n102 VTAIL.n98 2.41282
R1746 VTAIL.n147 VTAIL.n145 2.26774
R1747 VTAIL.n71 VTAIL.n1 2.26774
R1748 VTAIL.n258 VTAIL.n232 1.93989
R1749 VTAIL.n271 VTAIL.n226 1.93989
R1750 VTAIL.n42 VTAIL.n16 1.93989
R1751 VTAIL.n55 VTAIL.n10 1.93989
R1752 VTAIL.n201 VTAIL.n156 1.93989
R1753 VTAIL.n188 VTAIL.n162 1.93989
R1754 VTAIL.n129 VTAIL.n84 1.93989
R1755 VTAIL.n116 VTAIL.n90 1.93989
R1756 VTAIL.n259 VTAIL.n230 1.16414
R1757 VTAIL.n268 VTAIL.n267 1.16414
R1758 VTAIL.n43 VTAIL.n14 1.16414
R1759 VTAIL.n52 VTAIL.n51 1.16414
R1760 VTAIL.n198 VTAIL.n197 1.16414
R1761 VTAIL.n189 VTAIL.n160 1.16414
R1762 VTAIL.n126 VTAIL.n125 1.16414
R1763 VTAIL.n117 VTAIL.n88 1.16414
R1764 VTAIL VTAIL.n1 0.957397
R1765 VTAIL.n263 VTAIL.n262 0.388379
R1766 VTAIL.n264 VTAIL.n228 0.388379
R1767 VTAIL.n47 VTAIL.n46 0.388379
R1768 VTAIL.n48 VTAIL.n12 0.388379
R1769 VTAIL.n194 VTAIL.n158 0.388379
R1770 VTAIL.n193 VTAIL.n192 0.388379
R1771 VTAIL.n122 VTAIL.n86 0.388379
R1772 VTAIL.n121 VTAIL.n120 0.388379
R1773 VTAIL.n244 VTAIL.n243 0.155672
R1774 VTAIL.n244 VTAIL.n235 0.155672
R1775 VTAIL.n251 VTAIL.n235 0.155672
R1776 VTAIL.n252 VTAIL.n251 0.155672
R1777 VTAIL.n252 VTAIL.n231 0.155672
R1778 VTAIL.n260 VTAIL.n231 0.155672
R1779 VTAIL.n261 VTAIL.n260 0.155672
R1780 VTAIL.n261 VTAIL.n227 0.155672
R1781 VTAIL.n269 VTAIL.n227 0.155672
R1782 VTAIL.n270 VTAIL.n269 0.155672
R1783 VTAIL.n270 VTAIL.n223 0.155672
R1784 VTAIL.n277 VTAIL.n223 0.155672
R1785 VTAIL.n278 VTAIL.n277 0.155672
R1786 VTAIL.n278 VTAIL.n219 0.155672
R1787 VTAIL.n285 VTAIL.n219 0.155672
R1788 VTAIL.n28 VTAIL.n27 0.155672
R1789 VTAIL.n28 VTAIL.n19 0.155672
R1790 VTAIL.n35 VTAIL.n19 0.155672
R1791 VTAIL.n36 VTAIL.n35 0.155672
R1792 VTAIL.n36 VTAIL.n15 0.155672
R1793 VTAIL.n44 VTAIL.n15 0.155672
R1794 VTAIL.n45 VTAIL.n44 0.155672
R1795 VTAIL.n45 VTAIL.n11 0.155672
R1796 VTAIL.n53 VTAIL.n11 0.155672
R1797 VTAIL.n54 VTAIL.n53 0.155672
R1798 VTAIL.n54 VTAIL.n7 0.155672
R1799 VTAIL.n61 VTAIL.n7 0.155672
R1800 VTAIL.n62 VTAIL.n61 0.155672
R1801 VTAIL.n62 VTAIL.n3 0.155672
R1802 VTAIL.n69 VTAIL.n3 0.155672
R1803 VTAIL.n215 VTAIL.n149 0.155672
R1804 VTAIL.n208 VTAIL.n149 0.155672
R1805 VTAIL.n208 VTAIL.n207 0.155672
R1806 VTAIL.n207 VTAIL.n153 0.155672
R1807 VTAIL.n200 VTAIL.n153 0.155672
R1808 VTAIL.n200 VTAIL.n199 0.155672
R1809 VTAIL.n199 VTAIL.n157 0.155672
R1810 VTAIL.n191 VTAIL.n157 0.155672
R1811 VTAIL.n191 VTAIL.n190 0.155672
R1812 VTAIL.n190 VTAIL.n161 0.155672
R1813 VTAIL.n183 VTAIL.n161 0.155672
R1814 VTAIL.n183 VTAIL.n182 0.155672
R1815 VTAIL.n182 VTAIL.n166 0.155672
R1816 VTAIL.n175 VTAIL.n166 0.155672
R1817 VTAIL.n175 VTAIL.n174 0.155672
R1818 VTAIL.n143 VTAIL.n77 0.155672
R1819 VTAIL.n136 VTAIL.n77 0.155672
R1820 VTAIL.n136 VTAIL.n135 0.155672
R1821 VTAIL.n135 VTAIL.n81 0.155672
R1822 VTAIL.n128 VTAIL.n81 0.155672
R1823 VTAIL.n128 VTAIL.n127 0.155672
R1824 VTAIL.n127 VTAIL.n85 0.155672
R1825 VTAIL.n119 VTAIL.n85 0.155672
R1826 VTAIL.n119 VTAIL.n118 0.155672
R1827 VTAIL.n118 VTAIL.n89 0.155672
R1828 VTAIL.n111 VTAIL.n89 0.155672
R1829 VTAIL.n111 VTAIL.n110 0.155672
R1830 VTAIL.n110 VTAIL.n94 0.155672
R1831 VTAIL.n103 VTAIL.n94 0.155672
R1832 VTAIL.n103 VTAIL.n102 0.155672
R1833 VDD1.n64 VDD1.n0 756.745
R1834 VDD1.n133 VDD1.n69 756.745
R1835 VDD1.n65 VDD1.n64 585
R1836 VDD1.n63 VDD1.n62 585
R1837 VDD1.n4 VDD1.n3 585
R1838 VDD1.n57 VDD1.n56 585
R1839 VDD1.n55 VDD1.n54 585
R1840 VDD1.n8 VDD1.n7 585
R1841 VDD1.n49 VDD1.n48 585
R1842 VDD1.n47 VDD1.n46 585
R1843 VDD1.n45 VDD1.n11 585
R1844 VDD1.n15 VDD1.n12 585
R1845 VDD1.n40 VDD1.n39 585
R1846 VDD1.n38 VDD1.n37 585
R1847 VDD1.n17 VDD1.n16 585
R1848 VDD1.n32 VDD1.n31 585
R1849 VDD1.n30 VDD1.n29 585
R1850 VDD1.n21 VDD1.n20 585
R1851 VDD1.n24 VDD1.n23 585
R1852 VDD1.n92 VDD1.n91 585
R1853 VDD1.n89 VDD1.n88 585
R1854 VDD1.n98 VDD1.n97 585
R1855 VDD1.n100 VDD1.n99 585
R1856 VDD1.n85 VDD1.n84 585
R1857 VDD1.n106 VDD1.n105 585
R1858 VDD1.n109 VDD1.n108 585
R1859 VDD1.n107 VDD1.n81 585
R1860 VDD1.n114 VDD1.n80 585
R1861 VDD1.n116 VDD1.n115 585
R1862 VDD1.n118 VDD1.n117 585
R1863 VDD1.n77 VDD1.n76 585
R1864 VDD1.n124 VDD1.n123 585
R1865 VDD1.n126 VDD1.n125 585
R1866 VDD1.n73 VDD1.n72 585
R1867 VDD1.n132 VDD1.n131 585
R1868 VDD1.n134 VDD1.n133 585
R1869 VDD1.t0 VDD1.n90 329.036
R1870 VDD1.t3 VDD1.n22 329.036
R1871 VDD1.n64 VDD1.n63 171.744
R1872 VDD1.n63 VDD1.n3 171.744
R1873 VDD1.n56 VDD1.n3 171.744
R1874 VDD1.n56 VDD1.n55 171.744
R1875 VDD1.n55 VDD1.n7 171.744
R1876 VDD1.n48 VDD1.n7 171.744
R1877 VDD1.n48 VDD1.n47 171.744
R1878 VDD1.n47 VDD1.n11 171.744
R1879 VDD1.n15 VDD1.n11 171.744
R1880 VDD1.n39 VDD1.n15 171.744
R1881 VDD1.n39 VDD1.n38 171.744
R1882 VDD1.n38 VDD1.n16 171.744
R1883 VDD1.n31 VDD1.n16 171.744
R1884 VDD1.n31 VDD1.n30 171.744
R1885 VDD1.n30 VDD1.n20 171.744
R1886 VDD1.n23 VDD1.n20 171.744
R1887 VDD1.n91 VDD1.n88 171.744
R1888 VDD1.n98 VDD1.n88 171.744
R1889 VDD1.n99 VDD1.n98 171.744
R1890 VDD1.n99 VDD1.n84 171.744
R1891 VDD1.n106 VDD1.n84 171.744
R1892 VDD1.n108 VDD1.n106 171.744
R1893 VDD1.n108 VDD1.n107 171.744
R1894 VDD1.n107 VDD1.n80 171.744
R1895 VDD1.n116 VDD1.n80 171.744
R1896 VDD1.n117 VDD1.n116 171.744
R1897 VDD1.n117 VDD1.n76 171.744
R1898 VDD1.n124 VDD1.n76 171.744
R1899 VDD1.n125 VDD1.n124 171.744
R1900 VDD1.n125 VDD1.n72 171.744
R1901 VDD1.n132 VDD1.n72 171.744
R1902 VDD1.n133 VDD1.n132 171.744
R1903 VDD1.n23 VDD1.t3 85.8723
R1904 VDD1.n91 VDD1.t0 85.8723
R1905 VDD1.n139 VDD1.n138 74.6305
R1906 VDD1.n141 VDD1.n140 73.7869
R1907 VDD1 VDD1.n68 52.3942
R1908 VDD1.n139 VDD1.n137 52.2807
R1909 VDD1.n141 VDD1.n139 48.8824
R1910 VDD1.n46 VDD1.n45 13.1884
R1911 VDD1.n115 VDD1.n114 13.1884
R1912 VDD1.n49 VDD1.n10 12.8005
R1913 VDD1.n44 VDD1.n12 12.8005
R1914 VDD1.n113 VDD1.n81 12.8005
R1915 VDD1.n118 VDD1.n79 12.8005
R1916 VDD1.n50 VDD1.n8 12.0247
R1917 VDD1.n41 VDD1.n40 12.0247
R1918 VDD1.n110 VDD1.n109 12.0247
R1919 VDD1.n119 VDD1.n77 12.0247
R1920 VDD1.n54 VDD1.n53 11.249
R1921 VDD1.n37 VDD1.n14 11.249
R1922 VDD1.n105 VDD1.n83 11.249
R1923 VDD1.n123 VDD1.n122 11.249
R1924 VDD1.n24 VDD1.n22 10.7239
R1925 VDD1.n92 VDD1.n90 10.7239
R1926 VDD1.n57 VDD1.n6 10.4732
R1927 VDD1.n36 VDD1.n17 10.4732
R1928 VDD1.n104 VDD1.n85 10.4732
R1929 VDD1.n126 VDD1.n75 10.4732
R1930 VDD1.n58 VDD1.n4 9.69747
R1931 VDD1.n33 VDD1.n32 9.69747
R1932 VDD1.n101 VDD1.n100 9.69747
R1933 VDD1.n127 VDD1.n73 9.69747
R1934 VDD1.n68 VDD1.n67 9.45567
R1935 VDD1.n137 VDD1.n136 9.45567
R1936 VDD1.n26 VDD1.n25 9.3005
R1937 VDD1.n28 VDD1.n27 9.3005
R1938 VDD1.n19 VDD1.n18 9.3005
R1939 VDD1.n34 VDD1.n33 9.3005
R1940 VDD1.n36 VDD1.n35 9.3005
R1941 VDD1.n14 VDD1.n13 9.3005
R1942 VDD1.n42 VDD1.n41 9.3005
R1943 VDD1.n44 VDD1.n43 9.3005
R1944 VDD1.n67 VDD1.n66 9.3005
R1945 VDD1.n2 VDD1.n1 9.3005
R1946 VDD1.n61 VDD1.n60 9.3005
R1947 VDD1.n59 VDD1.n58 9.3005
R1948 VDD1.n6 VDD1.n5 9.3005
R1949 VDD1.n53 VDD1.n52 9.3005
R1950 VDD1.n51 VDD1.n50 9.3005
R1951 VDD1.n10 VDD1.n9 9.3005
R1952 VDD1.n71 VDD1.n70 9.3005
R1953 VDD1.n130 VDD1.n129 9.3005
R1954 VDD1.n128 VDD1.n127 9.3005
R1955 VDD1.n75 VDD1.n74 9.3005
R1956 VDD1.n122 VDD1.n121 9.3005
R1957 VDD1.n120 VDD1.n119 9.3005
R1958 VDD1.n79 VDD1.n78 9.3005
R1959 VDD1.n94 VDD1.n93 9.3005
R1960 VDD1.n96 VDD1.n95 9.3005
R1961 VDD1.n87 VDD1.n86 9.3005
R1962 VDD1.n102 VDD1.n101 9.3005
R1963 VDD1.n104 VDD1.n103 9.3005
R1964 VDD1.n83 VDD1.n82 9.3005
R1965 VDD1.n111 VDD1.n110 9.3005
R1966 VDD1.n113 VDD1.n112 9.3005
R1967 VDD1.n136 VDD1.n135 9.3005
R1968 VDD1.n62 VDD1.n61 8.92171
R1969 VDD1.n29 VDD1.n19 8.92171
R1970 VDD1.n97 VDD1.n87 8.92171
R1971 VDD1.n131 VDD1.n130 8.92171
R1972 VDD1.n65 VDD1.n2 8.14595
R1973 VDD1.n28 VDD1.n21 8.14595
R1974 VDD1.n96 VDD1.n89 8.14595
R1975 VDD1.n134 VDD1.n71 8.14595
R1976 VDD1.n66 VDD1.n0 7.3702
R1977 VDD1.n25 VDD1.n24 7.3702
R1978 VDD1.n93 VDD1.n92 7.3702
R1979 VDD1.n135 VDD1.n69 7.3702
R1980 VDD1.n68 VDD1.n0 6.59444
R1981 VDD1.n137 VDD1.n69 6.59444
R1982 VDD1.n66 VDD1.n65 5.81868
R1983 VDD1.n25 VDD1.n21 5.81868
R1984 VDD1.n93 VDD1.n89 5.81868
R1985 VDD1.n135 VDD1.n134 5.81868
R1986 VDD1.n62 VDD1.n2 5.04292
R1987 VDD1.n29 VDD1.n28 5.04292
R1988 VDD1.n97 VDD1.n96 5.04292
R1989 VDD1.n131 VDD1.n71 5.04292
R1990 VDD1.n61 VDD1.n4 4.26717
R1991 VDD1.n32 VDD1.n19 4.26717
R1992 VDD1.n100 VDD1.n87 4.26717
R1993 VDD1.n130 VDD1.n73 4.26717
R1994 VDD1.n58 VDD1.n57 3.49141
R1995 VDD1.n33 VDD1.n17 3.49141
R1996 VDD1.n101 VDD1.n85 3.49141
R1997 VDD1.n127 VDD1.n126 3.49141
R1998 VDD1.n54 VDD1.n6 2.71565
R1999 VDD1.n37 VDD1.n36 2.71565
R2000 VDD1.n105 VDD1.n104 2.71565
R2001 VDD1.n123 VDD1.n75 2.71565
R2002 VDD1.n140 VDD1.t1 2.52418
R2003 VDD1.n140 VDD1.t5 2.52418
R2004 VDD1.n138 VDD1.t2 2.52418
R2005 VDD1.n138 VDD1.t4 2.52418
R2006 VDD1.n26 VDD1.n22 2.41282
R2007 VDD1.n94 VDD1.n90 2.41282
R2008 VDD1.n53 VDD1.n8 1.93989
R2009 VDD1.n40 VDD1.n14 1.93989
R2010 VDD1.n109 VDD1.n83 1.93989
R2011 VDD1.n122 VDD1.n77 1.93989
R2012 VDD1.n50 VDD1.n49 1.16414
R2013 VDD1.n41 VDD1.n12 1.16414
R2014 VDD1.n110 VDD1.n81 1.16414
R2015 VDD1.n119 VDD1.n118 1.16414
R2016 VDD1 VDD1.n141 0.841017
R2017 VDD1.n46 VDD1.n10 0.388379
R2018 VDD1.n45 VDD1.n44 0.388379
R2019 VDD1.n114 VDD1.n113 0.388379
R2020 VDD1.n115 VDD1.n79 0.388379
R2021 VDD1.n67 VDD1.n1 0.155672
R2022 VDD1.n60 VDD1.n1 0.155672
R2023 VDD1.n60 VDD1.n59 0.155672
R2024 VDD1.n59 VDD1.n5 0.155672
R2025 VDD1.n52 VDD1.n5 0.155672
R2026 VDD1.n52 VDD1.n51 0.155672
R2027 VDD1.n51 VDD1.n9 0.155672
R2028 VDD1.n43 VDD1.n9 0.155672
R2029 VDD1.n43 VDD1.n42 0.155672
R2030 VDD1.n42 VDD1.n13 0.155672
R2031 VDD1.n35 VDD1.n13 0.155672
R2032 VDD1.n35 VDD1.n34 0.155672
R2033 VDD1.n34 VDD1.n18 0.155672
R2034 VDD1.n27 VDD1.n18 0.155672
R2035 VDD1.n27 VDD1.n26 0.155672
R2036 VDD1.n95 VDD1.n94 0.155672
R2037 VDD1.n95 VDD1.n86 0.155672
R2038 VDD1.n102 VDD1.n86 0.155672
R2039 VDD1.n103 VDD1.n102 0.155672
R2040 VDD1.n103 VDD1.n82 0.155672
R2041 VDD1.n111 VDD1.n82 0.155672
R2042 VDD1.n112 VDD1.n111 0.155672
R2043 VDD1.n112 VDD1.n78 0.155672
R2044 VDD1.n120 VDD1.n78 0.155672
R2045 VDD1.n121 VDD1.n120 0.155672
R2046 VDD1.n121 VDD1.n74 0.155672
R2047 VDD1.n128 VDD1.n74 0.155672
R2048 VDD1.n129 VDD1.n128 0.155672
R2049 VDD1.n129 VDD1.n70 0.155672
R2050 VDD1.n136 VDD1.n70 0.155672
R2051 VN.n37 VN.n20 161.3
R2052 VN.n36 VN.n35 161.3
R2053 VN.n34 VN.n21 161.3
R2054 VN.n33 VN.n32 161.3
R2055 VN.n31 VN.n22 161.3
R2056 VN.n30 VN.n29 161.3
R2057 VN.n28 VN.n23 161.3
R2058 VN.n27 VN.n26 161.3
R2059 VN.n17 VN.n0 161.3
R2060 VN.n16 VN.n15 161.3
R2061 VN.n14 VN.n1 161.3
R2062 VN.n13 VN.n12 161.3
R2063 VN.n11 VN.n2 161.3
R2064 VN.n10 VN.n9 161.3
R2065 VN.n8 VN.n3 161.3
R2066 VN.n7 VN.n6 161.3
R2067 VN.n4 VN.t1 113.004
R2068 VN.n24 VN.t0 113.004
R2069 VN.n5 VN.t2 80.8359
R2070 VN.n18 VN.t3 80.8359
R2071 VN.n25 VN.t5 80.8359
R2072 VN.n38 VN.t4 80.8359
R2073 VN.n5 VN.n4 62.6769
R2074 VN.n25 VN.n24 62.6769
R2075 VN.n19 VN.n18 61.5371
R2076 VN.n39 VN.n38 61.5371
R2077 VN.n12 VN.n11 56.4773
R2078 VN.n32 VN.n31 56.4773
R2079 VN VN.n39 54.4547
R2080 VN.n6 VN.n3 24.3439
R2081 VN.n10 VN.n3 24.3439
R2082 VN.n11 VN.n10 24.3439
R2083 VN.n12 VN.n1 24.3439
R2084 VN.n16 VN.n1 24.3439
R2085 VN.n17 VN.n16 24.3439
R2086 VN.n31 VN.n30 24.3439
R2087 VN.n30 VN.n23 24.3439
R2088 VN.n26 VN.n23 24.3439
R2089 VN.n37 VN.n36 24.3439
R2090 VN.n36 VN.n21 24.3439
R2091 VN.n32 VN.n21 24.3439
R2092 VN.n18 VN.n17 20.449
R2093 VN.n38 VN.n37 20.449
R2094 VN.n6 VN.n5 12.1722
R2095 VN.n26 VN.n25 12.1722
R2096 VN.n27 VN.n24 2.68625
R2097 VN.n7 VN.n4 2.68625
R2098 VN.n39 VN.n20 0.417764
R2099 VN.n19 VN.n0 0.417764
R2100 VN VN.n19 0.394061
R2101 VN.n35 VN.n20 0.189894
R2102 VN.n35 VN.n34 0.189894
R2103 VN.n34 VN.n33 0.189894
R2104 VN.n33 VN.n22 0.189894
R2105 VN.n29 VN.n22 0.189894
R2106 VN.n29 VN.n28 0.189894
R2107 VN.n28 VN.n27 0.189894
R2108 VN.n8 VN.n7 0.189894
R2109 VN.n9 VN.n8 0.189894
R2110 VN.n9 VN.n2 0.189894
R2111 VN.n13 VN.n2 0.189894
R2112 VN.n14 VN.n13 0.189894
R2113 VN.n15 VN.n14 0.189894
R2114 VN.n15 VN.n0 0.189894
R2115 VDD2.n135 VDD2.n71 756.745
R2116 VDD2.n64 VDD2.n0 756.745
R2117 VDD2.n136 VDD2.n135 585
R2118 VDD2.n134 VDD2.n133 585
R2119 VDD2.n75 VDD2.n74 585
R2120 VDD2.n128 VDD2.n127 585
R2121 VDD2.n126 VDD2.n125 585
R2122 VDD2.n79 VDD2.n78 585
R2123 VDD2.n120 VDD2.n119 585
R2124 VDD2.n118 VDD2.n117 585
R2125 VDD2.n116 VDD2.n82 585
R2126 VDD2.n86 VDD2.n83 585
R2127 VDD2.n111 VDD2.n110 585
R2128 VDD2.n109 VDD2.n108 585
R2129 VDD2.n88 VDD2.n87 585
R2130 VDD2.n103 VDD2.n102 585
R2131 VDD2.n101 VDD2.n100 585
R2132 VDD2.n92 VDD2.n91 585
R2133 VDD2.n95 VDD2.n94 585
R2134 VDD2.n23 VDD2.n22 585
R2135 VDD2.n20 VDD2.n19 585
R2136 VDD2.n29 VDD2.n28 585
R2137 VDD2.n31 VDD2.n30 585
R2138 VDD2.n16 VDD2.n15 585
R2139 VDD2.n37 VDD2.n36 585
R2140 VDD2.n40 VDD2.n39 585
R2141 VDD2.n38 VDD2.n12 585
R2142 VDD2.n45 VDD2.n11 585
R2143 VDD2.n47 VDD2.n46 585
R2144 VDD2.n49 VDD2.n48 585
R2145 VDD2.n8 VDD2.n7 585
R2146 VDD2.n55 VDD2.n54 585
R2147 VDD2.n57 VDD2.n56 585
R2148 VDD2.n4 VDD2.n3 585
R2149 VDD2.n63 VDD2.n62 585
R2150 VDD2.n65 VDD2.n64 585
R2151 VDD2.t4 VDD2.n21 329.036
R2152 VDD2.t1 VDD2.n93 329.036
R2153 VDD2.n135 VDD2.n134 171.744
R2154 VDD2.n134 VDD2.n74 171.744
R2155 VDD2.n127 VDD2.n74 171.744
R2156 VDD2.n127 VDD2.n126 171.744
R2157 VDD2.n126 VDD2.n78 171.744
R2158 VDD2.n119 VDD2.n78 171.744
R2159 VDD2.n119 VDD2.n118 171.744
R2160 VDD2.n118 VDD2.n82 171.744
R2161 VDD2.n86 VDD2.n82 171.744
R2162 VDD2.n110 VDD2.n86 171.744
R2163 VDD2.n110 VDD2.n109 171.744
R2164 VDD2.n109 VDD2.n87 171.744
R2165 VDD2.n102 VDD2.n87 171.744
R2166 VDD2.n102 VDD2.n101 171.744
R2167 VDD2.n101 VDD2.n91 171.744
R2168 VDD2.n94 VDD2.n91 171.744
R2169 VDD2.n22 VDD2.n19 171.744
R2170 VDD2.n29 VDD2.n19 171.744
R2171 VDD2.n30 VDD2.n29 171.744
R2172 VDD2.n30 VDD2.n15 171.744
R2173 VDD2.n37 VDD2.n15 171.744
R2174 VDD2.n39 VDD2.n37 171.744
R2175 VDD2.n39 VDD2.n38 171.744
R2176 VDD2.n38 VDD2.n11 171.744
R2177 VDD2.n47 VDD2.n11 171.744
R2178 VDD2.n48 VDD2.n47 171.744
R2179 VDD2.n48 VDD2.n7 171.744
R2180 VDD2.n55 VDD2.n7 171.744
R2181 VDD2.n56 VDD2.n55 171.744
R2182 VDD2.n56 VDD2.n3 171.744
R2183 VDD2.n63 VDD2.n3 171.744
R2184 VDD2.n64 VDD2.n63 171.744
R2185 VDD2.n94 VDD2.t1 85.8723
R2186 VDD2.n22 VDD2.t4 85.8723
R2187 VDD2.n70 VDD2.n69 74.6305
R2188 VDD2 VDD2.n141 74.6274
R2189 VDD2.n70 VDD2.n68 52.2807
R2190 VDD2.n140 VDD2.n139 49.6399
R2191 VDD2.n140 VDD2.n70 46.5019
R2192 VDD2.n117 VDD2.n116 13.1884
R2193 VDD2.n46 VDD2.n45 13.1884
R2194 VDD2.n120 VDD2.n81 12.8005
R2195 VDD2.n115 VDD2.n83 12.8005
R2196 VDD2.n44 VDD2.n12 12.8005
R2197 VDD2.n49 VDD2.n10 12.8005
R2198 VDD2.n121 VDD2.n79 12.0247
R2199 VDD2.n112 VDD2.n111 12.0247
R2200 VDD2.n41 VDD2.n40 12.0247
R2201 VDD2.n50 VDD2.n8 12.0247
R2202 VDD2.n125 VDD2.n124 11.249
R2203 VDD2.n108 VDD2.n85 11.249
R2204 VDD2.n36 VDD2.n14 11.249
R2205 VDD2.n54 VDD2.n53 11.249
R2206 VDD2.n95 VDD2.n93 10.7239
R2207 VDD2.n23 VDD2.n21 10.7239
R2208 VDD2.n128 VDD2.n77 10.4732
R2209 VDD2.n107 VDD2.n88 10.4732
R2210 VDD2.n35 VDD2.n16 10.4732
R2211 VDD2.n57 VDD2.n6 10.4732
R2212 VDD2.n129 VDD2.n75 9.69747
R2213 VDD2.n104 VDD2.n103 9.69747
R2214 VDD2.n32 VDD2.n31 9.69747
R2215 VDD2.n58 VDD2.n4 9.69747
R2216 VDD2.n139 VDD2.n138 9.45567
R2217 VDD2.n68 VDD2.n67 9.45567
R2218 VDD2.n97 VDD2.n96 9.3005
R2219 VDD2.n99 VDD2.n98 9.3005
R2220 VDD2.n90 VDD2.n89 9.3005
R2221 VDD2.n105 VDD2.n104 9.3005
R2222 VDD2.n107 VDD2.n106 9.3005
R2223 VDD2.n85 VDD2.n84 9.3005
R2224 VDD2.n113 VDD2.n112 9.3005
R2225 VDD2.n115 VDD2.n114 9.3005
R2226 VDD2.n138 VDD2.n137 9.3005
R2227 VDD2.n73 VDD2.n72 9.3005
R2228 VDD2.n132 VDD2.n131 9.3005
R2229 VDD2.n130 VDD2.n129 9.3005
R2230 VDD2.n77 VDD2.n76 9.3005
R2231 VDD2.n124 VDD2.n123 9.3005
R2232 VDD2.n122 VDD2.n121 9.3005
R2233 VDD2.n81 VDD2.n80 9.3005
R2234 VDD2.n2 VDD2.n1 9.3005
R2235 VDD2.n61 VDD2.n60 9.3005
R2236 VDD2.n59 VDD2.n58 9.3005
R2237 VDD2.n6 VDD2.n5 9.3005
R2238 VDD2.n53 VDD2.n52 9.3005
R2239 VDD2.n51 VDD2.n50 9.3005
R2240 VDD2.n10 VDD2.n9 9.3005
R2241 VDD2.n25 VDD2.n24 9.3005
R2242 VDD2.n27 VDD2.n26 9.3005
R2243 VDD2.n18 VDD2.n17 9.3005
R2244 VDD2.n33 VDD2.n32 9.3005
R2245 VDD2.n35 VDD2.n34 9.3005
R2246 VDD2.n14 VDD2.n13 9.3005
R2247 VDD2.n42 VDD2.n41 9.3005
R2248 VDD2.n44 VDD2.n43 9.3005
R2249 VDD2.n67 VDD2.n66 9.3005
R2250 VDD2.n133 VDD2.n132 8.92171
R2251 VDD2.n100 VDD2.n90 8.92171
R2252 VDD2.n28 VDD2.n18 8.92171
R2253 VDD2.n62 VDD2.n61 8.92171
R2254 VDD2.n136 VDD2.n73 8.14595
R2255 VDD2.n99 VDD2.n92 8.14595
R2256 VDD2.n27 VDD2.n20 8.14595
R2257 VDD2.n65 VDD2.n2 8.14595
R2258 VDD2.n137 VDD2.n71 7.3702
R2259 VDD2.n96 VDD2.n95 7.3702
R2260 VDD2.n24 VDD2.n23 7.3702
R2261 VDD2.n66 VDD2.n0 7.3702
R2262 VDD2.n139 VDD2.n71 6.59444
R2263 VDD2.n68 VDD2.n0 6.59444
R2264 VDD2.n137 VDD2.n136 5.81868
R2265 VDD2.n96 VDD2.n92 5.81868
R2266 VDD2.n24 VDD2.n20 5.81868
R2267 VDD2.n66 VDD2.n65 5.81868
R2268 VDD2.n133 VDD2.n73 5.04292
R2269 VDD2.n100 VDD2.n99 5.04292
R2270 VDD2.n28 VDD2.n27 5.04292
R2271 VDD2.n62 VDD2.n2 5.04292
R2272 VDD2.n132 VDD2.n75 4.26717
R2273 VDD2.n103 VDD2.n90 4.26717
R2274 VDD2.n31 VDD2.n18 4.26717
R2275 VDD2.n61 VDD2.n4 4.26717
R2276 VDD2.n129 VDD2.n128 3.49141
R2277 VDD2.n104 VDD2.n88 3.49141
R2278 VDD2.n32 VDD2.n16 3.49141
R2279 VDD2.n58 VDD2.n57 3.49141
R2280 VDD2 VDD2.n140 2.75481
R2281 VDD2.n125 VDD2.n77 2.71565
R2282 VDD2.n108 VDD2.n107 2.71565
R2283 VDD2.n36 VDD2.n35 2.71565
R2284 VDD2.n54 VDD2.n6 2.71565
R2285 VDD2.n141 VDD2.t0 2.52418
R2286 VDD2.n141 VDD2.t5 2.52418
R2287 VDD2.n69 VDD2.t3 2.52418
R2288 VDD2.n69 VDD2.t2 2.52418
R2289 VDD2.n97 VDD2.n93 2.41282
R2290 VDD2.n25 VDD2.n21 2.41282
R2291 VDD2.n124 VDD2.n79 1.93989
R2292 VDD2.n111 VDD2.n85 1.93989
R2293 VDD2.n40 VDD2.n14 1.93989
R2294 VDD2.n53 VDD2.n8 1.93989
R2295 VDD2.n121 VDD2.n120 1.16414
R2296 VDD2.n112 VDD2.n83 1.16414
R2297 VDD2.n41 VDD2.n12 1.16414
R2298 VDD2.n50 VDD2.n49 1.16414
R2299 VDD2.n117 VDD2.n81 0.388379
R2300 VDD2.n116 VDD2.n115 0.388379
R2301 VDD2.n45 VDD2.n44 0.388379
R2302 VDD2.n46 VDD2.n10 0.388379
R2303 VDD2.n138 VDD2.n72 0.155672
R2304 VDD2.n131 VDD2.n72 0.155672
R2305 VDD2.n131 VDD2.n130 0.155672
R2306 VDD2.n130 VDD2.n76 0.155672
R2307 VDD2.n123 VDD2.n76 0.155672
R2308 VDD2.n123 VDD2.n122 0.155672
R2309 VDD2.n122 VDD2.n80 0.155672
R2310 VDD2.n114 VDD2.n80 0.155672
R2311 VDD2.n114 VDD2.n113 0.155672
R2312 VDD2.n113 VDD2.n84 0.155672
R2313 VDD2.n106 VDD2.n84 0.155672
R2314 VDD2.n106 VDD2.n105 0.155672
R2315 VDD2.n105 VDD2.n89 0.155672
R2316 VDD2.n98 VDD2.n89 0.155672
R2317 VDD2.n98 VDD2.n97 0.155672
R2318 VDD2.n26 VDD2.n25 0.155672
R2319 VDD2.n26 VDD2.n17 0.155672
R2320 VDD2.n33 VDD2.n17 0.155672
R2321 VDD2.n34 VDD2.n33 0.155672
R2322 VDD2.n34 VDD2.n13 0.155672
R2323 VDD2.n42 VDD2.n13 0.155672
R2324 VDD2.n43 VDD2.n42 0.155672
R2325 VDD2.n43 VDD2.n9 0.155672
R2326 VDD2.n51 VDD2.n9 0.155672
R2327 VDD2.n52 VDD2.n51 0.155672
R2328 VDD2.n52 VDD2.n5 0.155672
R2329 VDD2.n59 VDD2.n5 0.155672
R2330 VDD2.n60 VDD2.n59 0.155672
R2331 VDD2.n60 VDD2.n1 0.155672
R2332 VDD2.n67 VDD2.n1 0.155672
C0 VDD1 VTAIL 8.46143f
C1 w_n4306_n3544# B 11.6354f
C2 B VP 2.37584f
C3 VDD2 VTAIL 8.521429f
C4 VDD1 VN 0.152192f
C5 w_n4306_n3544# VP 9.05284f
C6 VDD2 VN 7.64988f
C7 B VTAIL 4.36068f
C8 w_n4306_n3544# VTAIL 3.20392f
C9 VP VTAIL 8.0802f
C10 VDD1 VDD2 1.89161f
C11 B VN 1.43435f
C12 w_n4306_n3544# VN 8.49268f
C13 VP VN 8.30611f
C14 VDD1 B 2.48588f
C15 VDD1 w_n4306_n3544# 2.65132f
C16 VDD1 VP 8.057831f
C17 VDD2 B 2.58971f
C18 VN VTAIL 8.065351f
C19 VDD2 w_n4306_n3544# 2.77604f
C20 VDD2 VP 0.562677f
C21 VDD2 VSUBS 2.268074f
C22 VDD1 VSUBS 2.295718f
C23 VTAIL VSUBS 1.460607f
C24 VN VSUBS 7.11114f
C25 VP VSUBS 3.948563f
C26 B VSUBS 5.936007f
C27 w_n4306_n3544# VSUBS 0.187621p
C28 VDD2.n0 VSUBS 0.031966f
C29 VDD2.n1 VSUBS 0.028326f
C30 VDD2.n2 VSUBS 0.015221f
C31 VDD2.n3 VSUBS 0.035977f
C32 VDD2.n4 VSUBS 0.016117f
C33 VDD2.n5 VSUBS 0.028326f
C34 VDD2.n6 VSUBS 0.015221f
C35 VDD2.n7 VSUBS 0.035977f
C36 VDD2.n8 VSUBS 0.016117f
C37 VDD2.n9 VSUBS 0.028326f
C38 VDD2.n10 VSUBS 0.015221f
C39 VDD2.n11 VSUBS 0.035977f
C40 VDD2.n12 VSUBS 0.016117f
C41 VDD2.n13 VSUBS 0.028326f
C42 VDD2.n14 VSUBS 0.015221f
C43 VDD2.n15 VSUBS 0.035977f
C44 VDD2.n16 VSUBS 0.016117f
C45 VDD2.n17 VSUBS 0.028326f
C46 VDD2.n18 VSUBS 0.015221f
C47 VDD2.n19 VSUBS 0.035977f
C48 VDD2.n20 VSUBS 0.016117f
C49 VDD2.n21 VSUBS 0.234353f
C50 VDD2.t4 VSUBS 0.07761f
C51 VDD2.n22 VSUBS 0.026983f
C52 VDD2.n23 VSUBS 0.027064f
C53 VDD2.n24 VSUBS 0.015221f
C54 VDD2.n25 VSUBS 1.50097f
C55 VDD2.n26 VSUBS 0.028326f
C56 VDD2.n27 VSUBS 0.015221f
C57 VDD2.n28 VSUBS 0.016117f
C58 VDD2.n29 VSUBS 0.035977f
C59 VDD2.n30 VSUBS 0.035977f
C60 VDD2.n31 VSUBS 0.016117f
C61 VDD2.n32 VSUBS 0.015221f
C62 VDD2.n33 VSUBS 0.028326f
C63 VDD2.n34 VSUBS 0.028326f
C64 VDD2.n35 VSUBS 0.015221f
C65 VDD2.n36 VSUBS 0.016117f
C66 VDD2.n37 VSUBS 0.035977f
C67 VDD2.n38 VSUBS 0.035977f
C68 VDD2.n39 VSUBS 0.035977f
C69 VDD2.n40 VSUBS 0.016117f
C70 VDD2.n41 VSUBS 0.015221f
C71 VDD2.n42 VSUBS 0.028326f
C72 VDD2.n43 VSUBS 0.028326f
C73 VDD2.n44 VSUBS 0.015221f
C74 VDD2.n45 VSUBS 0.015669f
C75 VDD2.n46 VSUBS 0.015669f
C76 VDD2.n47 VSUBS 0.035977f
C77 VDD2.n48 VSUBS 0.035977f
C78 VDD2.n49 VSUBS 0.016117f
C79 VDD2.n50 VSUBS 0.015221f
C80 VDD2.n51 VSUBS 0.028326f
C81 VDD2.n52 VSUBS 0.028326f
C82 VDD2.n53 VSUBS 0.015221f
C83 VDD2.n54 VSUBS 0.016117f
C84 VDD2.n55 VSUBS 0.035977f
C85 VDD2.n56 VSUBS 0.035977f
C86 VDD2.n57 VSUBS 0.016117f
C87 VDD2.n58 VSUBS 0.015221f
C88 VDD2.n59 VSUBS 0.028326f
C89 VDD2.n60 VSUBS 0.028326f
C90 VDD2.n61 VSUBS 0.015221f
C91 VDD2.n62 VSUBS 0.016117f
C92 VDD2.n63 VSUBS 0.035977f
C93 VDD2.n64 VSUBS 0.089965f
C94 VDD2.n65 VSUBS 0.016117f
C95 VDD2.n66 VSUBS 0.015221f
C96 VDD2.n67 VSUBS 0.067022f
C97 VDD2.n68 VSUBS 0.079951f
C98 VDD2.t3 VSUBS 0.288306f
C99 VDD2.t2 VSUBS 0.288306f
C100 VDD2.n69 VSUBS 2.28967f
C101 VDD2.n70 VSUBS 4.00368f
C102 VDD2.n71 VSUBS 0.031966f
C103 VDD2.n72 VSUBS 0.028326f
C104 VDD2.n73 VSUBS 0.015221f
C105 VDD2.n74 VSUBS 0.035977f
C106 VDD2.n75 VSUBS 0.016117f
C107 VDD2.n76 VSUBS 0.028326f
C108 VDD2.n77 VSUBS 0.015221f
C109 VDD2.n78 VSUBS 0.035977f
C110 VDD2.n79 VSUBS 0.016117f
C111 VDD2.n80 VSUBS 0.028326f
C112 VDD2.n81 VSUBS 0.015221f
C113 VDD2.n82 VSUBS 0.035977f
C114 VDD2.n83 VSUBS 0.016117f
C115 VDD2.n84 VSUBS 0.028326f
C116 VDD2.n85 VSUBS 0.015221f
C117 VDD2.n86 VSUBS 0.035977f
C118 VDD2.n87 VSUBS 0.035977f
C119 VDD2.n88 VSUBS 0.016117f
C120 VDD2.n89 VSUBS 0.028326f
C121 VDD2.n90 VSUBS 0.015221f
C122 VDD2.n91 VSUBS 0.035977f
C123 VDD2.n92 VSUBS 0.016117f
C124 VDD2.n93 VSUBS 0.234353f
C125 VDD2.t1 VSUBS 0.07761f
C126 VDD2.n94 VSUBS 0.026983f
C127 VDD2.n95 VSUBS 0.027064f
C128 VDD2.n96 VSUBS 0.015221f
C129 VDD2.n97 VSUBS 1.50097f
C130 VDD2.n98 VSUBS 0.028326f
C131 VDD2.n99 VSUBS 0.015221f
C132 VDD2.n100 VSUBS 0.016117f
C133 VDD2.n101 VSUBS 0.035977f
C134 VDD2.n102 VSUBS 0.035977f
C135 VDD2.n103 VSUBS 0.016117f
C136 VDD2.n104 VSUBS 0.015221f
C137 VDD2.n105 VSUBS 0.028326f
C138 VDD2.n106 VSUBS 0.028326f
C139 VDD2.n107 VSUBS 0.015221f
C140 VDD2.n108 VSUBS 0.016117f
C141 VDD2.n109 VSUBS 0.035977f
C142 VDD2.n110 VSUBS 0.035977f
C143 VDD2.n111 VSUBS 0.016117f
C144 VDD2.n112 VSUBS 0.015221f
C145 VDD2.n113 VSUBS 0.028326f
C146 VDD2.n114 VSUBS 0.028326f
C147 VDD2.n115 VSUBS 0.015221f
C148 VDD2.n116 VSUBS 0.015669f
C149 VDD2.n117 VSUBS 0.015669f
C150 VDD2.n118 VSUBS 0.035977f
C151 VDD2.n119 VSUBS 0.035977f
C152 VDD2.n120 VSUBS 0.016117f
C153 VDD2.n121 VSUBS 0.015221f
C154 VDD2.n122 VSUBS 0.028326f
C155 VDD2.n123 VSUBS 0.028326f
C156 VDD2.n124 VSUBS 0.015221f
C157 VDD2.n125 VSUBS 0.016117f
C158 VDD2.n126 VSUBS 0.035977f
C159 VDD2.n127 VSUBS 0.035977f
C160 VDD2.n128 VSUBS 0.016117f
C161 VDD2.n129 VSUBS 0.015221f
C162 VDD2.n130 VSUBS 0.028326f
C163 VDD2.n131 VSUBS 0.028326f
C164 VDD2.n132 VSUBS 0.015221f
C165 VDD2.n133 VSUBS 0.016117f
C166 VDD2.n134 VSUBS 0.035977f
C167 VDD2.n135 VSUBS 0.089965f
C168 VDD2.n136 VSUBS 0.016117f
C169 VDD2.n137 VSUBS 0.015221f
C170 VDD2.n138 VSUBS 0.067022f
C171 VDD2.n139 VSUBS 0.064964f
C172 VDD2.n140 VSUBS 3.36351f
C173 VDD2.t0 VSUBS 0.288306f
C174 VDD2.t5 VSUBS 0.288306f
C175 VDD2.n141 VSUBS 2.28962f
C176 VN.n0 VSUBS 0.04548f
C177 VN.t3 VSUBS 3.26367f
C178 VN.n1 VSUBS 0.045276f
C179 VN.n2 VSUBS 0.024172f
C180 VN.n3 VSUBS 0.045276f
C181 VN.t1 VSUBS 3.64173f
C182 VN.n4 VSUBS 1.17015f
C183 VN.t2 VSUBS 3.26367f
C184 VN.n5 VSUBS 1.2268f
C185 VN.n6 VSUBS 0.034098f
C186 VN.n7 VSUBS 0.318352f
C187 VN.n8 VSUBS 0.024172f
C188 VN.n9 VSUBS 0.024172f
C189 VN.n10 VSUBS 0.045276f
C190 VN.n11 VSUBS 0.041206f
C191 VN.n12 VSUBS 0.029674f
C192 VN.n13 VSUBS 0.024172f
C193 VN.n14 VSUBS 0.024172f
C194 VN.n15 VSUBS 0.024172f
C195 VN.n16 VSUBS 0.045276f
C196 VN.n17 VSUBS 0.041699f
C197 VN.n18 VSUBS 1.24369f
C198 VN.n19 VSUBS 0.075265f
C199 VN.n20 VSUBS 0.04548f
C200 VN.t4 VSUBS 3.26367f
C201 VN.n21 VSUBS 0.045276f
C202 VN.n22 VSUBS 0.024172f
C203 VN.n23 VSUBS 0.045276f
C204 VN.t0 VSUBS 3.64173f
C205 VN.n24 VSUBS 1.17015f
C206 VN.t5 VSUBS 3.26367f
C207 VN.n25 VSUBS 1.2268f
C208 VN.n26 VSUBS 0.034098f
C209 VN.n27 VSUBS 0.318352f
C210 VN.n28 VSUBS 0.024172f
C211 VN.n29 VSUBS 0.024172f
C212 VN.n30 VSUBS 0.045276f
C213 VN.n31 VSUBS 0.041206f
C214 VN.n32 VSUBS 0.029674f
C215 VN.n33 VSUBS 0.024172f
C216 VN.n34 VSUBS 0.024172f
C217 VN.n35 VSUBS 0.024172f
C218 VN.n36 VSUBS 0.045276f
C219 VN.n37 VSUBS 0.041699f
C220 VN.n38 VSUBS 1.24369f
C221 VN.n39 VSUBS 1.58466f
C222 VDD1.n0 VSUBS 0.032255f
C223 VDD1.n1 VSUBS 0.028582f
C224 VDD1.n2 VSUBS 0.015359f
C225 VDD1.n3 VSUBS 0.036303f
C226 VDD1.n4 VSUBS 0.016262f
C227 VDD1.n5 VSUBS 0.028582f
C228 VDD1.n6 VSUBS 0.015359f
C229 VDD1.n7 VSUBS 0.036303f
C230 VDD1.n8 VSUBS 0.016262f
C231 VDD1.n9 VSUBS 0.028582f
C232 VDD1.n10 VSUBS 0.015359f
C233 VDD1.n11 VSUBS 0.036303f
C234 VDD1.n12 VSUBS 0.016262f
C235 VDD1.n13 VSUBS 0.028582f
C236 VDD1.n14 VSUBS 0.015359f
C237 VDD1.n15 VSUBS 0.036303f
C238 VDD1.n16 VSUBS 0.036303f
C239 VDD1.n17 VSUBS 0.016262f
C240 VDD1.n18 VSUBS 0.028582f
C241 VDD1.n19 VSUBS 0.015359f
C242 VDD1.n20 VSUBS 0.036303f
C243 VDD1.n21 VSUBS 0.016262f
C244 VDD1.n22 VSUBS 0.236472f
C245 VDD1.t3 VSUBS 0.078312f
C246 VDD1.n23 VSUBS 0.027227f
C247 VDD1.n24 VSUBS 0.027309f
C248 VDD1.n25 VSUBS 0.015359f
C249 VDD1.n26 VSUBS 1.51454f
C250 VDD1.n27 VSUBS 0.028582f
C251 VDD1.n28 VSUBS 0.015359f
C252 VDD1.n29 VSUBS 0.016262f
C253 VDD1.n30 VSUBS 0.036303f
C254 VDD1.n31 VSUBS 0.036303f
C255 VDD1.n32 VSUBS 0.016262f
C256 VDD1.n33 VSUBS 0.015359f
C257 VDD1.n34 VSUBS 0.028582f
C258 VDD1.n35 VSUBS 0.028582f
C259 VDD1.n36 VSUBS 0.015359f
C260 VDD1.n37 VSUBS 0.016262f
C261 VDD1.n38 VSUBS 0.036303f
C262 VDD1.n39 VSUBS 0.036303f
C263 VDD1.n40 VSUBS 0.016262f
C264 VDD1.n41 VSUBS 0.015359f
C265 VDD1.n42 VSUBS 0.028582f
C266 VDD1.n43 VSUBS 0.028582f
C267 VDD1.n44 VSUBS 0.015359f
C268 VDD1.n45 VSUBS 0.015811f
C269 VDD1.n46 VSUBS 0.015811f
C270 VDD1.n47 VSUBS 0.036303f
C271 VDD1.n48 VSUBS 0.036303f
C272 VDD1.n49 VSUBS 0.016262f
C273 VDD1.n50 VSUBS 0.015359f
C274 VDD1.n51 VSUBS 0.028582f
C275 VDD1.n52 VSUBS 0.028582f
C276 VDD1.n53 VSUBS 0.015359f
C277 VDD1.n54 VSUBS 0.016262f
C278 VDD1.n55 VSUBS 0.036303f
C279 VDD1.n56 VSUBS 0.036303f
C280 VDD1.n57 VSUBS 0.016262f
C281 VDD1.n58 VSUBS 0.015359f
C282 VDD1.n59 VSUBS 0.028582f
C283 VDD1.n60 VSUBS 0.028582f
C284 VDD1.n61 VSUBS 0.015359f
C285 VDD1.n62 VSUBS 0.016262f
C286 VDD1.n63 VSUBS 0.036303f
C287 VDD1.n64 VSUBS 0.090779f
C288 VDD1.n65 VSUBS 0.016262f
C289 VDD1.n66 VSUBS 0.015359f
C290 VDD1.n67 VSUBS 0.067628f
C291 VDD1.n68 VSUBS 0.081827f
C292 VDD1.n69 VSUBS 0.032255f
C293 VDD1.n70 VSUBS 0.028582f
C294 VDD1.n71 VSUBS 0.015359f
C295 VDD1.n72 VSUBS 0.036303f
C296 VDD1.n73 VSUBS 0.016262f
C297 VDD1.n74 VSUBS 0.028582f
C298 VDD1.n75 VSUBS 0.015359f
C299 VDD1.n76 VSUBS 0.036303f
C300 VDD1.n77 VSUBS 0.016262f
C301 VDD1.n78 VSUBS 0.028582f
C302 VDD1.n79 VSUBS 0.015359f
C303 VDD1.n80 VSUBS 0.036303f
C304 VDD1.n81 VSUBS 0.016262f
C305 VDD1.n82 VSUBS 0.028582f
C306 VDD1.n83 VSUBS 0.015359f
C307 VDD1.n84 VSUBS 0.036303f
C308 VDD1.n85 VSUBS 0.016262f
C309 VDD1.n86 VSUBS 0.028582f
C310 VDD1.n87 VSUBS 0.015359f
C311 VDD1.n88 VSUBS 0.036303f
C312 VDD1.n89 VSUBS 0.016262f
C313 VDD1.n90 VSUBS 0.236472f
C314 VDD1.t0 VSUBS 0.078312f
C315 VDD1.n91 VSUBS 0.027227f
C316 VDD1.n92 VSUBS 0.027309f
C317 VDD1.n93 VSUBS 0.015359f
C318 VDD1.n94 VSUBS 1.51454f
C319 VDD1.n95 VSUBS 0.028582f
C320 VDD1.n96 VSUBS 0.015359f
C321 VDD1.n97 VSUBS 0.016262f
C322 VDD1.n98 VSUBS 0.036303f
C323 VDD1.n99 VSUBS 0.036303f
C324 VDD1.n100 VSUBS 0.016262f
C325 VDD1.n101 VSUBS 0.015359f
C326 VDD1.n102 VSUBS 0.028582f
C327 VDD1.n103 VSUBS 0.028582f
C328 VDD1.n104 VSUBS 0.015359f
C329 VDD1.n105 VSUBS 0.016262f
C330 VDD1.n106 VSUBS 0.036303f
C331 VDD1.n107 VSUBS 0.036303f
C332 VDD1.n108 VSUBS 0.036303f
C333 VDD1.n109 VSUBS 0.016262f
C334 VDD1.n110 VSUBS 0.015359f
C335 VDD1.n111 VSUBS 0.028582f
C336 VDD1.n112 VSUBS 0.028582f
C337 VDD1.n113 VSUBS 0.015359f
C338 VDD1.n114 VSUBS 0.015811f
C339 VDD1.n115 VSUBS 0.015811f
C340 VDD1.n116 VSUBS 0.036303f
C341 VDD1.n117 VSUBS 0.036303f
C342 VDD1.n118 VSUBS 0.016262f
C343 VDD1.n119 VSUBS 0.015359f
C344 VDD1.n120 VSUBS 0.028582f
C345 VDD1.n121 VSUBS 0.028582f
C346 VDD1.n122 VSUBS 0.015359f
C347 VDD1.n123 VSUBS 0.016262f
C348 VDD1.n124 VSUBS 0.036303f
C349 VDD1.n125 VSUBS 0.036303f
C350 VDD1.n126 VSUBS 0.016262f
C351 VDD1.n127 VSUBS 0.015359f
C352 VDD1.n128 VSUBS 0.028582f
C353 VDD1.n129 VSUBS 0.028582f
C354 VDD1.n130 VSUBS 0.015359f
C355 VDD1.n131 VSUBS 0.016262f
C356 VDD1.n132 VSUBS 0.036303f
C357 VDD1.n133 VSUBS 0.090779f
C358 VDD1.n134 VSUBS 0.016262f
C359 VDD1.n135 VSUBS 0.015359f
C360 VDD1.n136 VSUBS 0.067628f
C361 VDD1.n137 VSUBS 0.080674f
C362 VDD1.t2 VSUBS 0.290913f
C363 VDD1.t4 VSUBS 0.290913f
C364 VDD1.n138 VSUBS 2.31037f
C365 VDD1.n139 VSUBS 4.22064f
C366 VDD1.t1 VSUBS 0.290913f
C367 VDD1.t5 VSUBS 0.290913f
C368 VDD1.n140 VSUBS 2.2995f
C369 VDD1.n141 VSUBS 3.97046f
C370 VTAIL.t1 VSUBS 0.304103f
C371 VTAIL.t0 VSUBS 0.304103f
C372 VTAIL.n0 VSUBS 2.24016f
C373 VTAIL.n1 VSUBS 0.999248f
C374 VTAIL.n2 VSUBS 0.033718f
C375 VTAIL.n3 VSUBS 0.029878f
C376 VTAIL.n4 VSUBS 0.016055f
C377 VTAIL.n5 VSUBS 0.037949f
C378 VTAIL.n6 VSUBS 0.017f
C379 VTAIL.n7 VSUBS 0.029878f
C380 VTAIL.n8 VSUBS 0.016055f
C381 VTAIL.n9 VSUBS 0.037949f
C382 VTAIL.n10 VSUBS 0.017f
C383 VTAIL.n11 VSUBS 0.029878f
C384 VTAIL.n12 VSUBS 0.016055f
C385 VTAIL.n13 VSUBS 0.037949f
C386 VTAIL.n14 VSUBS 0.017f
C387 VTAIL.n15 VSUBS 0.029878f
C388 VTAIL.n16 VSUBS 0.016055f
C389 VTAIL.n17 VSUBS 0.037949f
C390 VTAIL.n18 VSUBS 0.017f
C391 VTAIL.n19 VSUBS 0.029878f
C392 VTAIL.n20 VSUBS 0.016055f
C393 VTAIL.n21 VSUBS 0.037949f
C394 VTAIL.n22 VSUBS 0.017f
C395 VTAIL.n23 VSUBS 0.247194f
C396 VTAIL.t9 VSUBS 0.081862f
C397 VTAIL.n24 VSUBS 0.028461f
C398 VTAIL.n25 VSUBS 0.028547f
C399 VTAIL.n26 VSUBS 0.016055f
C400 VTAIL.n27 VSUBS 1.58321f
C401 VTAIL.n28 VSUBS 0.029878f
C402 VTAIL.n29 VSUBS 0.016055f
C403 VTAIL.n30 VSUBS 0.017f
C404 VTAIL.n31 VSUBS 0.037949f
C405 VTAIL.n32 VSUBS 0.037949f
C406 VTAIL.n33 VSUBS 0.017f
C407 VTAIL.n34 VSUBS 0.016055f
C408 VTAIL.n35 VSUBS 0.029878f
C409 VTAIL.n36 VSUBS 0.029878f
C410 VTAIL.n37 VSUBS 0.016055f
C411 VTAIL.n38 VSUBS 0.017f
C412 VTAIL.n39 VSUBS 0.037949f
C413 VTAIL.n40 VSUBS 0.037949f
C414 VTAIL.n41 VSUBS 0.037949f
C415 VTAIL.n42 VSUBS 0.017f
C416 VTAIL.n43 VSUBS 0.016055f
C417 VTAIL.n44 VSUBS 0.029878f
C418 VTAIL.n45 VSUBS 0.029878f
C419 VTAIL.n46 VSUBS 0.016055f
C420 VTAIL.n47 VSUBS 0.016527f
C421 VTAIL.n48 VSUBS 0.016527f
C422 VTAIL.n49 VSUBS 0.037949f
C423 VTAIL.n50 VSUBS 0.037949f
C424 VTAIL.n51 VSUBS 0.017f
C425 VTAIL.n52 VSUBS 0.016055f
C426 VTAIL.n53 VSUBS 0.029878f
C427 VTAIL.n54 VSUBS 0.029878f
C428 VTAIL.n55 VSUBS 0.016055f
C429 VTAIL.n56 VSUBS 0.017f
C430 VTAIL.n57 VSUBS 0.037949f
C431 VTAIL.n58 VSUBS 0.037949f
C432 VTAIL.n59 VSUBS 0.017f
C433 VTAIL.n60 VSUBS 0.016055f
C434 VTAIL.n61 VSUBS 0.029878f
C435 VTAIL.n62 VSUBS 0.029878f
C436 VTAIL.n63 VSUBS 0.016055f
C437 VTAIL.n64 VSUBS 0.017f
C438 VTAIL.n65 VSUBS 0.037949f
C439 VTAIL.n66 VSUBS 0.094895f
C440 VTAIL.n67 VSUBS 0.017f
C441 VTAIL.n68 VSUBS 0.016055f
C442 VTAIL.n69 VSUBS 0.070694f
C443 VTAIL.n70 VSUBS 0.047906f
C444 VTAIL.n71 VSUBS 0.590803f
C445 VTAIL.t11 VSUBS 0.304103f
C446 VTAIL.t8 VSUBS 0.304103f
C447 VTAIL.n72 VSUBS 2.24016f
C448 VTAIL.n73 VSUBS 3.20194f
C449 VTAIL.t5 VSUBS 0.304103f
C450 VTAIL.t2 VSUBS 0.304103f
C451 VTAIL.n74 VSUBS 2.24017f
C452 VTAIL.n75 VSUBS 3.20193f
C453 VTAIL.n76 VSUBS 0.033718f
C454 VTAIL.n77 VSUBS 0.029878f
C455 VTAIL.n78 VSUBS 0.016055f
C456 VTAIL.n79 VSUBS 0.037949f
C457 VTAIL.n80 VSUBS 0.017f
C458 VTAIL.n81 VSUBS 0.029878f
C459 VTAIL.n82 VSUBS 0.016055f
C460 VTAIL.n83 VSUBS 0.037949f
C461 VTAIL.n84 VSUBS 0.017f
C462 VTAIL.n85 VSUBS 0.029878f
C463 VTAIL.n86 VSUBS 0.016055f
C464 VTAIL.n87 VSUBS 0.037949f
C465 VTAIL.n88 VSUBS 0.017f
C466 VTAIL.n89 VSUBS 0.029878f
C467 VTAIL.n90 VSUBS 0.016055f
C468 VTAIL.n91 VSUBS 0.037949f
C469 VTAIL.n92 VSUBS 0.037949f
C470 VTAIL.n93 VSUBS 0.017f
C471 VTAIL.n94 VSUBS 0.029878f
C472 VTAIL.n95 VSUBS 0.016055f
C473 VTAIL.n96 VSUBS 0.037949f
C474 VTAIL.n97 VSUBS 0.017f
C475 VTAIL.n98 VSUBS 0.247194f
C476 VTAIL.t3 VSUBS 0.081862f
C477 VTAIL.n99 VSUBS 0.028461f
C478 VTAIL.n100 VSUBS 0.028547f
C479 VTAIL.n101 VSUBS 0.016055f
C480 VTAIL.n102 VSUBS 1.58321f
C481 VTAIL.n103 VSUBS 0.029878f
C482 VTAIL.n104 VSUBS 0.016055f
C483 VTAIL.n105 VSUBS 0.017f
C484 VTAIL.n106 VSUBS 0.037949f
C485 VTAIL.n107 VSUBS 0.037949f
C486 VTAIL.n108 VSUBS 0.017f
C487 VTAIL.n109 VSUBS 0.016055f
C488 VTAIL.n110 VSUBS 0.029878f
C489 VTAIL.n111 VSUBS 0.029878f
C490 VTAIL.n112 VSUBS 0.016055f
C491 VTAIL.n113 VSUBS 0.017f
C492 VTAIL.n114 VSUBS 0.037949f
C493 VTAIL.n115 VSUBS 0.037949f
C494 VTAIL.n116 VSUBS 0.017f
C495 VTAIL.n117 VSUBS 0.016055f
C496 VTAIL.n118 VSUBS 0.029878f
C497 VTAIL.n119 VSUBS 0.029878f
C498 VTAIL.n120 VSUBS 0.016055f
C499 VTAIL.n121 VSUBS 0.016527f
C500 VTAIL.n122 VSUBS 0.016527f
C501 VTAIL.n123 VSUBS 0.037949f
C502 VTAIL.n124 VSUBS 0.037949f
C503 VTAIL.n125 VSUBS 0.017f
C504 VTAIL.n126 VSUBS 0.016055f
C505 VTAIL.n127 VSUBS 0.029878f
C506 VTAIL.n128 VSUBS 0.029878f
C507 VTAIL.n129 VSUBS 0.016055f
C508 VTAIL.n130 VSUBS 0.017f
C509 VTAIL.n131 VSUBS 0.037949f
C510 VTAIL.n132 VSUBS 0.037949f
C511 VTAIL.n133 VSUBS 0.017f
C512 VTAIL.n134 VSUBS 0.016055f
C513 VTAIL.n135 VSUBS 0.029878f
C514 VTAIL.n136 VSUBS 0.029878f
C515 VTAIL.n137 VSUBS 0.016055f
C516 VTAIL.n138 VSUBS 0.017f
C517 VTAIL.n139 VSUBS 0.037949f
C518 VTAIL.n140 VSUBS 0.094895f
C519 VTAIL.n141 VSUBS 0.017f
C520 VTAIL.n142 VSUBS 0.016055f
C521 VTAIL.n143 VSUBS 0.070694f
C522 VTAIL.n144 VSUBS 0.047906f
C523 VTAIL.n145 VSUBS 0.590803f
C524 VTAIL.t10 VSUBS 0.304103f
C525 VTAIL.t6 VSUBS 0.304103f
C526 VTAIL.n146 VSUBS 2.24017f
C527 VTAIL.n147 VSUBS 1.2532f
C528 VTAIL.n148 VSUBS 0.033718f
C529 VTAIL.n149 VSUBS 0.029878f
C530 VTAIL.n150 VSUBS 0.016055f
C531 VTAIL.n151 VSUBS 0.037949f
C532 VTAIL.n152 VSUBS 0.017f
C533 VTAIL.n153 VSUBS 0.029878f
C534 VTAIL.n154 VSUBS 0.016055f
C535 VTAIL.n155 VSUBS 0.037949f
C536 VTAIL.n156 VSUBS 0.017f
C537 VTAIL.n157 VSUBS 0.029878f
C538 VTAIL.n158 VSUBS 0.016055f
C539 VTAIL.n159 VSUBS 0.037949f
C540 VTAIL.n160 VSUBS 0.017f
C541 VTAIL.n161 VSUBS 0.029878f
C542 VTAIL.n162 VSUBS 0.016055f
C543 VTAIL.n163 VSUBS 0.037949f
C544 VTAIL.n164 VSUBS 0.037949f
C545 VTAIL.n165 VSUBS 0.017f
C546 VTAIL.n166 VSUBS 0.029878f
C547 VTAIL.n167 VSUBS 0.016055f
C548 VTAIL.n168 VSUBS 0.037949f
C549 VTAIL.n169 VSUBS 0.017f
C550 VTAIL.n170 VSUBS 0.247194f
C551 VTAIL.t7 VSUBS 0.081862f
C552 VTAIL.n171 VSUBS 0.028461f
C553 VTAIL.n172 VSUBS 0.028547f
C554 VTAIL.n173 VSUBS 0.016055f
C555 VTAIL.n174 VSUBS 1.58321f
C556 VTAIL.n175 VSUBS 0.029878f
C557 VTAIL.n176 VSUBS 0.016055f
C558 VTAIL.n177 VSUBS 0.017f
C559 VTAIL.n178 VSUBS 0.037949f
C560 VTAIL.n179 VSUBS 0.037949f
C561 VTAIL.n180 VSUBS 0.017f
C562 VTAIL.n181 VSUBS 0.016055f
C563 VTAIL.n182 VSUBS 0.029878f
C564 VTAIL.n183 VSUBS 0.029878f
C565 VTAIL.n184 VSUBS 0.016055f
C566 VTAIL.n185 VSUBS 0.017f
C567 VTAIL.n186 VSUBS 0.037949f
C568 VTAIL.n187 VSUBS 0.037949f
C569 VTAIL.n188 VSUBS 0.017f
C570 VTAIL.n189 VSUBS 0.016055f
C571 VTAIL.n190 VSUBS 0.029878f
C572 VTAIL.n191 VSUBS 0.029878f
C573 VTAIL.n192 VSUBS 0.016055f
C574 VTAIL.n193 VSUBS 0.016527f
C575 VTAIL.n194 VSUBS 0.016527f
C576 VTAIL.n195 VSUBS 0.037949f
C577 VTAIL.n196 VSUBS 0.037949f
C578 VTAIL.n197 VSUBS 0.017f
C579 VTAIL.n198 VSUBS 0.016055f
C580 VTAIL.n199 VSUBS 0.029878f
C581 VTAIL.n200 VSUBS 0.029878f
C582 VTAIL.n201 VSUBS 0.016055f
C583 VTAIL.n202 VSUBS 0.017f
C584 VTAIL.n203 VSUBS 0.037949f
C585 VTAIL.n204 VSUBS 0.037949f
C586 VTAIL.n205 VSUBS 0.017f
C587 VTAIL.n206 VSUBS 0.016055f
C588 VTAIL.n207 VSUBS 0.029878f
C589 VTAIL.n208 VSUBS 0.029878f
C590 VTAIL.n209 VSUBS 0.016055f
C591 VTAIL.n210 VSUBS 0.017f
C592 VTAIL.n211 VSUBS 0.037949f
C593 VTAIL.n212 VSUBS 0.094895f
C594 VTAIL.n213 VSUBS 0.017f
C595 VTAIL.n214 VSUBS 0.016055f
C596 VTAIL.n215 VSUBS 0.070694f
C597 VTAIL.n216 VSUBS 0.047906f
C598 VTAIL.n217 VSUBS 2.19344f
C599 VTAIL.n218 VSUBS 0.033718f
C600 VTAIL.n219 VSUBS 0.029878f
C601 VTAIL.n220 VSUBS 0.016055f
C602 VTAIL.n221 VSUBS 0.037949f
C603 VTAIL.n222 VSUBS 0.017f
C604 VTAIL.n223 VSUBS 0.029878f
C605 VTAIL.n224 VSUBS 0.016055f
C606 VTAIL.n225 VSUBS 0.037949f
C607 VTAIL.n226 VSUBS 0.017f
C608 VTAIL.n227 VSUBS 0.029878f
C609 VTAIL.n228 VSUBS 0.016055f
C610 VTAIL.n229 VSUBS 0.037949f
C611 VTAIL.n230 VSUBS 0.017f
C612 VTAIL.n231 VSUBS 0.029878f
C613 VTAIL.n232 VSUBS 0.016055f
C614 VTAIL.n233 VSUBS 0.037949f
C615 VTAIL.n234 VSUBS 0.017f
C616 VTAIL.n235 VSUBS 0.029878f
C617 VTAIL.n236 VSUBS 0.016055f
C618 VTAIL.n237 VSUBS 0.037949f
C619 VTAIL.n238 VSUBS 0.017f
C620 VTAIL.n239 VSUBS 0.247194f
C621 VTAIL.t4 VSUBS 0.081862f
C622 VTAIL.n240 VSUBS 0.028461f
C623 VTAIL.n241 VSUBS 0.028547f
C624 VTAIL.n242 VSUBS 0.016055f
C625 VTAIL.n243 VSUBS 1.58321f
C626 VTAIL.n244 VSUBS 0.029878f
C627 VTAIL.n245 VSUBS 0.016055f
C628 VTAIL.n246 VSUBS 0.017f
C629 VTAIL.n247 VSUBS 0.037949f
C630 VTAIL.n248 VSUBS 0.037949f
C631 VTAIL.n249 VSUBS 0.017f
C632 VTAIL.n250 VSUBS 0.016055f
C633 VTAIL.n251 VSUBS 0.029878f
C634 VTAIL.n252 VSUBS 0.029878f
C635 VTAIL.n253 VSUBS 0.016055f
C636 VTAIL.n254 VSUBS 0.017f
C637 VTAIL.n255 VSUBS 0.037949f
C638 VTAIL.n256 VSUBS 0.037949f
C639 VTAIL.n257 VSUBS 0.037949f
C640 VTAIL.n258 VSUBS 0.017f
C641 VTAIL.n259 VSUBS 0.016055f
C642 VTAIL.n260 VSUBS 0.029878f
C643 VTAIL.n261 VSUBS 0.029878f
C644 VTAIL.n262 VSUBS 0.016055f
C645 VTAIL.n263 VSUBS 0.016527f
C646 VTAIL.n264 VSUBS 0.016527f
C647 VTAIL.n265 VSUBS 0.037949f
C648 VTAIL.n266 VSUBS 0.037949f
C649 VTAIL.n267 VSUBS 0.017f
C650 VTAIL.n268 VSUBS 0.016055f
C651 VTAIL.n269 VSUBS 0.029878f
C652 VTAIL.n270 VSUBS 0.029878f
C653 VTAIL.n271 VSUBS 0.016055f
C654 VTAIL.n272 VSUBS 0.017f
C655 VTAIL.n273 VSUBS 0.037949f
C656 VTAIL.n274 VSUBS 0.037949f
C657 VTAIL.n275 VSUBS 0.017f
C658 VTAIL.n276 VSUBS 0.016055f
C659 VTAIL.n277 VSUBS 0.029878f
C660 VTAIL.n278 VSUBS 0.029878f
C661 VTAIL.n279 VSUBS 0.016055f
C662 VTAIL.n280 VSUBS 0.017f
C663 VTAIL.n281 VSUBS 0.037949f
C664 VTAIL.n282 VSUBS 0.094895f
C665 VTAIL.n283 VSUBS 0.017f
C666 VTAIL.n284 VSUBS 0.016055f
C667 VTAIL.n285 VSUBS 0.070694f
C668 VTAIL.n286 VSUBS 0.047906f
C669 VTAIL.n287 VSUBS 2.10132f
C670 VP.n0 VSUBS 0.05043f
C671 VP.t1 VSUBS 3.61892f
C672 VP.n1 VSUBS 0.050204f
C673 VP.n2 VSUBS 0.026803f
C674 VP.n3 VSUBS 0.050204f
C675 VP.n4 VSUBS 0.026803f
C676 VP.t3 VSUBS 3.61892f
C677 VP.n5 VSUBS 0.050204f
C678 VP.n6 VSUBS 0.026803f
C679 VP.n7 VSUBS 0.050204f
C680 VP.n8 VSUBS 0.05043f
C681 VP.t0 VSUBS 3.61892f
C682 VP.n9 VSUBS 0.050204f
C683 VP.n10 VSUBS 0.026803f
C684 VP.n11 VSUBS 0.050204f
C685 VP.t2 VSUBS 4.03813f
C686 VP.n12 VSUBS 1.29752f
C687 VP.t4 VSUBS 3.61892f
C688 VP.n13 VSUBS 1.36034f
C689 VP.n14 VSUBS 0.03781f
C690 VP.n15 VSUBS 0.353007f
C691 VP.n16 VSUBS 0.026803f
C692 VP.n17 VSUBS 0.026803f
C693 VP.n18 VSUBS 0.050204f
C694 VP.n19 VSUBS 0.045691f
C695 VP.n20 VSUBS 0.032904f
C696 VP.n21 VSUBS 0.026803f
C697 VP.n22 VSUBS 0.026803f
C698 VP.n23 VSUBS 0.026803f
C699 VP.n24 VSUBS 0.050204f
C700 VP.n25 VSUBS 0.046238f
C701 VP.n26 VSUBS 1.37907f
C702 VP.n27 VSUBS 1.75055f
C703 VP.n28 VSUBS 1.76821f
C704 VP.t5 VSUBS 3.61892f
C705 VP.n29 VSUBS 1.37907f
C706 VP.n30 VSUBS 0.046238f
C707 VP.n31 VSUBS 0.05043f
C708 VP.n32 VSUBS 0.026803f
C709 VP.n33 VSUBS 0.026803f
C710 VP.n34 VSUBS 0.050204f
C711 VP.n35 VSUBS 0.032904f
C712 VP.n36 VSUBS 0.045691f
C713 VP.n37 VSUBS 0.026803f
C714 VP.n38 VSUBS 0.026803f
C715 VP.n39 VSUBS 0.026803f
C716 VP.n40 VSUBS 0.050204f
C717 VP.n41 VSUBS 0.03781f
C718 VP.n42 VSUBS 1.26314f
C719 VP.n43 VSUBS 0.03781f
C720 VP.n44 VSUBS 0.026803f
C721 VP.n45 VSUBS 0.026803f
C722 VP.n46 VSUBS 0.026803f
C723 VP.n47 VSUBS 0.050204f
C724 VP.n48 VSUBS 0.045691f
C725 VP.n49 VSUBS 0.032904f
C726 VP.n50 VSUBS 0.026803f
C727 VP.n51 VSUBS 0.026803f
C728 VP.n52 VSUBS 0.026803f
C729 VP.n53 VSUBS 0.050204f
C730 VP.n54 VSUBS 0.046238f
C731 VP.n55 VSUBS 1.37907f
C732 VP.n56 VSUBS 0.083457f
C733 B.n0 VSUBS 0.00514f
C734 B.n1 VSUBS 0.00514f
C735 B.n2 VSUBS 0.008128f
C736 B.n3 VSUBS 0.008128f
C737 B.n4 VSUBS 0.008128f
C738 B.n5 VSUBS 0.008128f
C739 B.n6 VSUBS 0.008128f
C740 B.n7 VSUBS 0.008128f
C741 B.n8 VSUBS 0.008128f
C742 B.n9 VSUBS 0.008128f
C743 B.n10 VSUBS 0.008128f
C744 B.n11 VSUBS 0.008128f
C745 B.n12 VSUBS 0.008128f
C746 B.n13 VSUBS 0.008128f
C747 B.n14 VSUBS 0.008128f
C748 B.n15 VSUBS 0.008128f
C749 B.n16 VSUBS 0.008128f
C750 B.n17 VSUBS 0.008128f
C751 B.n18 VSUBS 0.008128f
C752 B.n19 VSUBS 0.008128f
C753 B.n20 VSUBS 0.008128f
C754 B.n21 VSUBS 0.008128f
C755 B.n22 VSUBS 0.008128f
C756 B.n23 VSUBS 0.008128f
C757 B.n24 VSUBS 0.008128f
C758 B.n25 VSUBS 0.008128f
C759 B.n26 VSUBS 0.008128f
C760 B.n27 VSUBS 0.008128f
C761 B.n28 VSUBS 0.008128f
C762 B.n29 VSUBS 0.008128f
C763 B.n30 VSUBS 0.019032f
C764 B.n31 VSUBS 0.008128f
C765 B.n32 VSUBS 0.008128f
C766 B.n33 VSUBS 0.008128f
C767 B.n34 VSUBS 0.008128f
C768 B.n35 VSUBS 0.008128f
C769 B.n36 VSUBS 0.008128f
C770 B.n37 VSUBS 0.008128f
C771 B.n38 VSUBS 0.008128f
C772 B.n39 VSUBS 0.008128f
C773 B.n40 VSUBS 0.008128f
C774 B.n41 VSUBS 0.008128f
C775 B.n42 VSUBS 0.008128f
C776 B.n43 VSUBS 0.008128f
C777 B.n44 VSUBS 0.008128f
C778 B.n45 VSUBS 0.008128f
C779 B.n46 VSUBS 0.008128f
C780 B.n47 VSUBS 0.008128f
C781 B.n48 VSUBS 0.008128f
C782 B.n49 VSUBS 0.008128f
C783 B.n50 VSUBS 0.008128f
C784 B.n51 VSUBS 0.008128f
C785 B.n52 VSUBS 0.00765f
C786 B.n53 VSUBS 0.008128f
C787 B.t8 VSUBS 0.268205f
C788 B.t7 VSUBS 0.319645f
C789 B.t6 VSUBS 2.66996f
C790 B.n54 VSUBS 0.509461f
C791 B.n55 VSUBS 0.312151f
C792 B.n56 VSUBS 0.018832f
C793 B.n57 VSUBS 0.008128f
C794 B.n58 VSUBS 0.008128f
C795 B.n59 VSUBS 0.008128f
C796 B.n60 VSUBS 0.008128f
C797 B.t5 VSUBS 0.268208f
C798 B.t4 VSUBS 0.319648f
C799 B.t3 VSUBS 2.66996f
C800 B.n61 VSUBS 0.509458f
C801 B.n62 VSUBS 0.312147f
C802 B.n63 VSUBS 0.008128f
C803 B.n64 VSUBS 0.008128f
C804 B.n65 VSUBS 0.008128f
C805 B.n66 VSUBS 0.008128f
C806 B.n67 VSUBS 0.008128f
C807 B.n68 VSUBS 0.008128f
C808 B.n69 VSUBS 0.008128f
C809 B.n70 VSUBS 0.008128f
C810 B.n71 VSUBS 0.008128f
C811 B.n72 VSUBS 0.008128f
C812 B.n73 VSUBS 0.008128f
C813 B.n74 VSUBS 0.008128f
C814 B.n75 VSUBS 0.008128f
C815 B.n76 VSUBS 0.008128f
C816 B.n77 VSUBS 0.008128f
C817 B.n78 VSUBS 0.008128f
C818 B.n79 VSUBS 0.008128f
C819 B.n80 VSUBS 0.008128f
C820 B.n81 VSUBS 0.008128f
C821 B.n82 VSUBS 0.008128f
C822 B.n83 VSUBS 0.008128f
C823 B.n84 VSUBS 0.020174f
C824 B.n85 VSUBS 0.008128f
C825 B.n86 VSUBS 0.008128f
C826 B.n87 VSUBS 0.008128f
C827 B.n88 VSUBS 0.008128f
C828 B.n89 VSUBS 0.008128f
C829 B.n90 VSUBS 0.008128f
C830 B.n91 VSUBS 0.008128f
C831 B.n92 VSUBS 0.008128f
C832 B.n93 VSUBS 0.008128f
C833 B.n94 VSUBS 0.008128f
C834 B.n95 VSUBS 0.008128f
C835 B.n96 VSUBS 0.008128f
C836 B.n97 VSUBS 0.008128f
C837 B.n98 VSUBS 0.008128f
C838 B.n99 VSUBS 0.008128f
C839 B.n100 VSUBS 0.008128f
C840 B.n101 VSUBS 0.008128f
C841 B.n102 VSUBS 0.008128f
C842 B.n103 VSUBS 0.008128f
C843 B.n104 VSUBS 0.008128f
C844 B.n105 VSUBS 0.008128f
C845 B.n106 VSUBS 0.008128f
C846 B.n107 VSUBS 0.008128f
C847 B.n108 VSUBS 0.008128f
C848 B.n109 VSUBS 0.008128f
C849 B.n110 VSUBS 0.008128f
C850 B.n111 VSUBS 0.008128f
C851 B.n112 VSUBS 0.008128f
C852 B.n113 VSUBS 0.008128f
C853 B.n114 VSUBS 0.008128f
C854 B.n115 VSUBS 0.008128f
C855 B.n116 VSUBS 0.008128f
C856 B.n117 VSUBS 0.008128f
C857 B.n118 VSUBS 0.008128f
C858 B.n119 VSUBS 0.008128f
C859 B.n120 VSUBS 0.008128f
C860 B.n121 VSUBS 0.008128f
C861 B.n122 VSUBS 0.008128f
C862 B.n123 VSUBS 0.008128f
C863 B.n124 VSUBS 0.008128f
C864 B.n125 VSUBS 0.008128f
C865 B.n126 VSUBS 0.008128f
C866 B.n127 VSUBS 0.008128f
C867 B.n128 VSUBS 0.008128f
C868 B.n129 VSUBS 0.008128f
C869 B.n130 VSUBS 0.008128f
C870 B.n131 VSUBS 0.008128f
C871 B.n132 VSUBS 0.008128f
C872 B.n133 VSUBS 0.008128f
C873 B.n134 VSUBS 0.008128f
C874 B.n135 VSUBS 0.008128f
C875 B.n136 VSUBS 0.008128f
C876 B.n137 VSUBS 0.008128f
C877 B.n138 VSUBS 0.008128f
C878 B.n139 VSUBS 0.008128f
C879 B.n140 VSUBS 0.008128f
C880 B.n141 VSUBS 0.008128f
C881 B.n142 VSUBS 0.020174f
C882 B.n143 VSUBS 0.008128f
C883 B.n144 VSUBS 0.008128f
C884 B.n145 VSUBS 0.008128f
C885 B.n146 VSUBS 0.008128f
C886 B.n147 VSUBS 0.008128f
C887 B.n148 VSUBS 0.008128f
C888 B.n149 VSUBS 0.008128f
C889 B.n150 VSUBS 0.008128f
C890 B.n151 VSUBS 0.008128f
C891 B.n152 VSUBS 0.008128f
C892 B.n153 VSUBS 0.008128f
C893 B.n154 VSUBS 0.008128f
C894 B.n155 VSUBS 0.008128f
C895 B.n156 VSUBS 0.008128f
C896 B.n157 VSUBS 0.008128f
C897 B.n158 VSUBS 0.008128f
C898 B.n159 VSUBS 0.008128f
C899 B.n160 VSUBS 0.008128f
C900 B.n161 VSUBS 0.008128f
C901 B.n162 VSUBS 0.008128f
C902 B.n163 VSUBS 0.008128f
C903 B.n164 VSUBS 0.008128f
C904 B.t10 VSUBS 0.268208f
C905 B.t11 VSUBS 0.319648f
C906 B.t9 VSUBS 2.66996f
C907 B.n165 VSUBS 0.509458f
C908 B.n166 VSUBS 0.312147f
C909 B.n167 VSUBS 0.008128f
C910 B.n168 VSUBS 0.008128f
C911 B.n169 VSUBS 0.008128f
C912 B.n170 VSUBS 0.008128f
C913 B.t1 VSUBS 0.268205f
C914 B.t2 VSUBS 0.319645f
C915 B.t0 VSUBS 2.66996f
C916 B.n171 VSUBS 0.509461f
C917 B.n172 VSUBS 0.312151f
C918 B.n173 VSUBS 0.018832f
C919 B.n174 VSUBS 0.008128f
C920 B.n175 VSUBS 0.008128f
C921 B.n176 VSUBS 0.008128f
C922 B.n177 VSUBS 0.008128f
C923 B.n178 VSUBS 0.008128f
C924 B.n179 VSUBS 0.008128f
C925 B.n180 VSUBS 0.008128f
C926 B.n181 VSUBS 0.008128f
C927 B.n182 VSUBS 0.008128f
C928 B.n183 VSUBS 0.008128f
C929 B.n184 VSUBS 0.008128f
C930 B.n185 VSUBS 0.008128f
C931 B.n186 VSUBS 0.008128f
C932 B.n187 VSUBS 0.008128f
C933 B.n188 VSUBS 0.008128f
C934 B.n189 VSUBS 0.008128f
C935 B.n190 VSUBS 0.008128f
C936 B.n191 VSUBS 0.008128f
C937 B.n192 VSUBS 0.008128f
C938 B.n193 VSUBS 0.008128f
C939 B.n194 VSUBS 0.008128f
C940 B.n195 VSUBS 0.020174f
C941 B.n196 VSUBS 0.008128f
C942 B.n197 VSUBS 0.008128f
C943 B.n198 VSUBS 0.008128f
C944 B.n199 VSUBS 0.008128f
C945 B.n200 VSUBS 0.008128f
C946 B.n201 VSUBS 0.008128f
C947 B.n202 VSUBS 0.008128f
C948 B.n203 VSUBS 0.008128f
C949 B.n204 VSUBS 0.008128f
C950 B.n205 VSUBS 0.008128f
C951 B.n206 VSUBS 0.008128f
C952 B.n207 VSUBS 0.008128f
C953 B.n208 VSUBS 0.008128f
C954 B.n209 VSUBS 0.008128f
C955 B.n210 VSUBS 0.008128f
C956 B.n211 VSUBS 0.008128f
C957 B.n212 VSUBS 0.008128f
C958 B.n213 VSUBS 0.008128f
C959 B.n214 VSUBS 0.008128f
C960 B.n215 VSUBS 0.008128f
C961 B.n216 VSUBS 0.008128f
C962 B.n217 VSUBS 0.008128f
C963 B.n218 VSUBS 0.008128f
C964 B.n219 VSUBS 0.008128f
C965 B.n220 VSUBS 0.008128f
C966 B.n221 VSUBS 0.008128f
C967 B.n222 VSUBS 0.008128f
C968 B.n223 VSUBS 0.008128f
C969 B.n224 VSUBS 0.008128f
C970 B.n225 VSUBS 0.008128f
C971 B.n226 VSUBS 0.008128f
C972 B.n227 VSUBS 0.008128f
C973 B.n228 VSUBS 0.008128f
C974 B.n229 VSUBS 0.008128f
C975 B.n230 VSUBS 0.008128f
C976 B.n231 VSUBS 0.008128f
C977 B.n232 VSUBS 0.008128f
C978 B.n233 VSUBS 0.008128f
C979 B.n234 VSUBS 0.008128f
C980 B.n235 VSUBS 0.008128f
C981 B.n236 VSUBS 0.008128f
C982 B.n237 VSUBS 0.008128f
C983 B.n238 VSUBS 0.008128f
C984 B.n239 VSUBS 0.008128f
C985 B.n240 VSUBS 0.008128f
C986 B.n241 VSUBS 0.008128f
C987 B.n242 VSUBS 0.008128f
C988 B.n243 VSUBS 0.008128f
C989 B.n244 VSUBS 0.008128f
C990 B.n245 VSUBS 0.008128f
C991 B.n246 VSUBS 0.008128f
C992 B.n247 VSUBS 0.008128f
C993 B.n248 VSUBS 0.008128f
C994 B.n249 VSUBS 0.008128f
C995 B.n250 VSUBS 0.008128f
C996 B.n251 VSUBS 0.008128f
C997 B.n252 VSUBS 0.008128f
C998 B.n253 VSUBS 0.008128f
C999 B.n254 VSUBS 0.008128f
C1000 B.n255 VSUBS 0.008128f
C1001 B.n256 VSUBS 0.008128f
C1002 B.n257 VSUBS 0.008128f
C1003 B.n258 VSUBS 0.008128f
C1004 B.n259 VSUBS 0.008128f
C1005 B.n260 VSUBS 0.008128f
C1006 B.n261 VSUBS 0.008128f
C1007 B.n262 VSUBS 0.008128f
C1008 B.n263 VSUBS 0.008128f
C1009 B.n264 VSUBS 0.008128f
C1010 B.n265 VSUBS 0.008128f
C1011 B.n266 VSUBS 0.008128f
C1012 B.n267 VSUBS 0.008128f
C1013 B.n268 VSUBS 0.008128f
C1014 B.n269 VSUBS 0.008128f
C1015 B.n270 VSUBS 0.008128f
C1016 B.n271 VSUBS 0.008128f
C1017 B.n272 VSUBS 0.008128f
C1018 B.n273 VSUBS 0.008128f
C1019 B.n274 VSUBS 0.008128f
C1020 B.n275 VSUBS 0.008128f
C1021 B.n276 VSUBS 0.008128f
C1022 B.n277 VSUBS 0.008128f
C1023 B.n278 VSUBS 0.008128f
C1024 B.n279 VSUBS 0.008128f
C1025 B.n280 VSUBS 0.008128f
C1026 B.n281 VSUBS 0.008128f
C1027 B.n282 VSUBS 0.008128f
C1028 B.n283 VSUBS 0.008128f
C1029 B.n284 VSUBS 0.008128f
C1030 B.n285 VSUBS 0.008128f
C1031 B.n286 VSUBS 0.008128f
C1032 B.n287 VSUBS 0.008128f
C1033 B.n288 VSUBS 0.008128f
C1034 B.n289 VSUBS 0.008128f
C1035 B.n290 VSUBS 0.008128f
C1036 B.n291 VSUBS 0.008128f
C1037 B.n292 VSUBS 0.008128f
C1038 B.n293 VSUBS 0.008128f
C1039 B.n294 VSUBS 0.008128f
C1040 B.n295 VSUBS 0.008128f
C1041 B.n296 VSUBS 0.008128f
C1042 B.n297 VSUBS 0.008128f
C1043 B.n298 VSUBS 0.008128f
C1044 B.n299 VSUBS 0.008128f
C1045 B.n300 VSUBS 0.008128f
C1046 B.n301 VSUBS 0.008128f
C1047 B.n302 VSUBS 0.008128f
C1048 B.n303 VSUBS 0.008128f
C1049 B.n304 VSUBS 0.008128f
C1050 B.n305 VSUBS 0.008128f
C1051 B.n306 VSUBS 0.019032f
C1052 B.n307 VSUBS 0.019032f
C1053 B.n308 VSUBS 0.020174f
C1054 B.n309 VSUBS 0.008128f
C1055 B.n310 VSUBS 0.008128f
C1056 B.n311 VSUBS 0.008128f
C1057 B.n312 VSUBS 0.008128f
C1058 B.n313 VSUBS 0.008128f
C1059 B.n314 VSUBS 0.008128f
C1060 B.n315 VSUBS 0.008128f
C1061 B.n316 VSUBS 0.008128f
C1062 B.n317 VSUBS 0.008128f
C1063 B.n318 VSUBS 0.008128f
C1064 B.n319 VSUBS 0.008128f
C1065 B.n320 VSUBS 0.008128f
C1066 B.n321 VSUBS 0.008128f
C1067 B.n322 VSUBS 0.008128f
C1068 B.n323 VSUBS 0.008128f
C1069 B.n324 VSUBS 0.008128f
C1070 B.n325 VSUBS 0.008128f
C1071 B.n326 VSUBS 0.008128f
C1072 B.n327 VSUBS 0.008128f
C1073 B.n328 VSUBS 0.008128f
C1074 B.n329 VSUBS 0.008128f
C1075 B.n330 VSUBS 0.008128f
C1076 B.n331 VSUBS 0.008128f
C1077 B.n332 VSUBS 0.008128f
C1078 B.n333 VSUBS 0.008128f
C1079 B.n334 VSUBS 0.008128f
C1080 B.n335 VSUBS 0.008128f
C1081 B.n336 VSUBS 0.008128f
C1082 B.n337 VSUBS 0.008128f
C1083 B.n338 VSUBS 0.008128f
C1084 B.n339 VSUBS 0.008128f
C1085 B.n340 VSUBS 0.008128f
C1086 B.n341 VSUBS 0.008128f
C1087 B.n342 VSUBS 0.008128f
C1088 B.n343 VSUBS 0.008128f
C1089 B.n344 VSUBS 0.008128f
C1090 B.n345 VSUBS 0.008128f
C1091 B.n346 VSUBS 0.008128f
C1092 B.n347 VSUBS 0.008128f
C1093 B.n348 VSUBS 0.008128f
C1094 B.n349 VSUBS 0.008128f
C1095 B.n350 VSUBS 0.008128f
C1096 B.n351 VSUBS 0.008128f
C1097 B.n352 VSUBS 0.008128f
C1098 B.n353 VSUBS 0.008128f
C1099 B.n354 VSUBS 0.008128f
C1100 B.n355 VSUBS 0.008128f
C1101 B.n356 VSUBS 0.008128f
C1102 B.n357 VSUBS 0.008128f
C1103 B.n358 VSUBS 0.008128f
C1104 B.n359 VSUBS 0.008128f
C1105 B.n360 VSUBS 0.008128f
C1106 B.n361 VSUBS 0.008128f
C1107 B.n362 VSUBS 0.008128f
C1108 B.n363 VSUBS 0.008128f
C1109 B.n364 VSUBS 0.008128f
C1110 B.n365 VSUBS 0.008128f
C1111 B.n366 VSUBS 0.008128f
C1112 B.n367 VSUBS 0.008128f
C1113 B.n368 VSUBS 0.008128f
C1114 B.n369 VSUBS 0.008128f
C1115 B.n370 VSUBS 0.008128f
C1116 B.n371 VSUBS 0.008128f
C1117 B.n372 VSUBS 0.00765f
C1118 B.n373 VSUBS 0.008128f
C1119 B.n374 VSUBS 0.008128f
C1120 B.n375 VSUBS 0.004542f
C1121 B.n376 VSUBS 0.008128f
C1122 B.n377 VSUBS 0.008128f
C1123 B.n378 VSUBS 0.008128f
C1124 B.n379 VSUBS 0.008128f
C1125 B.n380 VSUBS 0.008128f
C1126 B.n381 VSUBS 0.008128f
C1127 B.n382 VSUBS 0.008128f
C1128 B.n383 VSUBS 0.008128f
C1129 B.n384 VSUBS 0.008128f
C1130 B.n385 VSUBS 0.008128f
C1131 B.n386 VSUBS 0.008128f
C1132 B.n387 VSUBS 0.008128f
C1133 B.n388 VSUBS 0.004542f
C1134 B.n389 VSUBS 0.018832f
C1135 B.n390 VSUBS 0.00765f
C1136 B.n391 VSUBS 0.008128f
C1137 B.n392 VSUBS 0.008128f
C1138 B.n393 VSUBS 0.008128f
C1139 B.n394 VSUBS 0.008128f
C1140 B.n395 VSUBS 0.008128f
C1141 B.n396 VSUBS 0.008128f
C1142 B.n397 VSUBS 0.008128f
C1143 B.n398 VSUBS 0.008128f
C1144 B.n399 VSUBS 0.008128f
C1145 B.n400 VSUBS 0.008128f
C1146 B.n401 VSUBS 0.008128f
C1147 B.n402 VSUBS 0.008128f
C1148 B.n403 VSUBS 0.008128f
C1149 B.n404 VSUBS 0.008128f
C1150 B.n405 VSUBS 0.008128f
C1151 B.n406 VSUBS 0.008128f
C1152 B.n407 VSUBS 0.008128f
C1153 B.n408 VSUBS 0.008128f
C1154 B.n409 VSUBS 0.008128f
C1155 B.n410 VSUBS 0.008128f
C1156 B.n411 VSUBS 0.008128f
C1157 B.n412 VSUBS 0.008128f
C1158 B.n413 VSUBS 0.008128f
C1159 B.n414 VSUBS 0.008128f
C1160 B.n415 VSUBS 0.008128f
C1161 B.n416 VSUBS 0.008128f
C1162 B.n417 VSUBS 0.008128f
C1163 B.n418 VSUBS 0.008128f
C1164 B.n419 VSUBS 0.008128f
C1165 B.n420 VSUBS 0.008128f
C1166 B.n421 VSUBS 0.008128f
C1167 B.n422 VSUBS 0.008128f
C1168 B.n423 VSUBS 0.008128f
C1169 B.n424 VSUBS 0.008128f
C1170 B.n425 VSUBS 0.008128f
C1171 B.n426 VSUBS 0.008128f
C1172 B.n427 VSUBS 0.008128f
C1173 B.n428 VSUBS 0.008128f
C1174 B.n429 VSUBS 0.008128f
C1175 B.n430 VSUBS 0.008128f
C1176 B.n431 VSUBS 0.008128f
C1177 B.n432 VSUBS 0.008128f
C1178 B.n433 VSUBS 0.008128f
C1179 B.n434 VSUBS 0.008128f
C1180 B.n435 VSUBS 0.008128f
C1181 B.n436 VSUBS 0.008128f
C1182 B.n437 VSUBS 0.008128f
C1183 B.n438 VSUBS 0.008128f
C1184 B.n439 VSUBS 0.008128f
C1185 B.n440 VSUBS 0.008128f
C1186 B.n441 VSUBS 0.008128f
C1187 B.n442 VSUBS 0.008128f
C1188 B.n443 VSUBS 0.008128f
C1189 B.n444 VSUBS 0.008128f
C1190 B.n445 VSUBS 0.008128f
C1191 B.n446 VSUBS 0.008128f
C1192 B.n447 VSUBS 0.008128f
C1193 B.n448 VSUBS 0.008128f
C1194 B.n449 VSUBS 0.008128f
C1195 B.n450 VSUBS 0.008128f
C1196 B.n451 VSUBS 0.008128f
C1197 B.n452 VSUBS 0.008128f
C1198 B.n453 VSUBS 0.008128f
C1199 B.n454 VSUBS 0.008128f
C1200 B.n455 VSUBS 0.020174f
C1201 B.n456 VSUBS 0.019032f
C1202 B.n457 VSUBS 0.019032f
C1203 B.n458 VSUBS 0.008128f
C1204 B.n459 VSUBS 0.008128f
C1205 B.n460 VSUBS 0.008128f
C1206 B.n461 VSUBS 0.008128f
C1207 B.n462 VSUBS 0.008128f
C1208 B.n463 VSUBS 0.008128f
C1209 B.n464 VSUBS 0.008128f
C1210 B.n465 VSUBS 0.008128f
C1211 B.n466 VSUBS 0.008128f
C1212 B.n467 VSUBS 0.008128f
C1213 B.n468 VSUBS 0.008128f
C1214 B.n469 VSUBS 0.008128f
C1215 B.n470 VSUBS 0.008128f
C1216 B.n471 VSUBS 0.008128f
C1217 B.n472 VSUBS 0.008128f
C1218 B.n473 VSUBS 0.008128f
C1219 B.n474 VSUBS 0.008128f
C1220 B.n475 VSUBS 0.008128f
C1221 B.n476 VSUBS 0.008128f
C1222 B.n477 VSUBS 0.008128f
C1223 B.n478 VSUBS 0.008128f
C1224 B.n479 VSUBS 0.008128f
C1225 B.n480 VSUBS 0.008128f
C1226 B.n481 VSUBS 0.008128f
C1227 B.n482 VSUBS 0.008128f
C1228 B.n483 VSUBS 0.008128f
C1229 B.n484 VSUBS 0.008128f
C1230 B.n485 VSUBS 0.008128f
C1231 B.n486 VSUBS 0.008128f
C1232 B.n487 VSUBS 0.008128f
C1233 B.n488 VSUBS 0.008128f
C1234 B.n489 VSUBS 0.008128f
C1235 B.n490 VSUBS 0.008128f
C1236 B.n491 VSUBS 0.008128f
C1237 B.n492 VSUBS 0.008128f
C1238 B.n493 VSUBS 0.008128f
C1239 B.n494 VSUBS 0.008128f
C1240 B.n495 VSUBS 0.008128f
C1241 B.n496 VSUBS 0.008128f
C1242 B.n497 VSUBS 0.008128f
C1243 B.n498 VSUBS 0.008128f
C1244 B.n499 VSUBS 0.008128f
C1245 B.n500 VSUBS 0.008128f
C1246 B.n501 VSUBS 0.008128f
C1247 B.n502 VSUBS 0.008128f
C1248 B.n503 VSUBS 0.008128f
C1249 B.n504 VSUBS 0.008128f
C1250 B.n505 VSUBS 0.008128f
C1251 B.n506 VSUBS 0.008128f
C1252 B.n507 VSUBS 0.008128f
C1253 B.n508 VSUBS 0.008128f
C1254 B.n509 VSUBS 0.008128f
C1255 B.n510 VSUBS 0.008128f
C1256 B.n511 VSUBS 0.008128f
C1257 B.n512 VSUBS 0.008128f
C1258 B.n513 VSUBS 0.008128f
C1259 B.n514 VSUBS 0.008128f
C1260 B.n515 VSUBS 0.008128f
C1261 B.n516 VSUBS 0.008128f
C1262 B.n517 VSUBS 0.008128f
C1263 B.n518 VSUBS 0.008128f
C1264 B.n519 VSUBS 0.008128f
C1265 B.n520 VSUBS 0.008128f
C1266 B.n521 VSUBS 0.008128f
C1267 B.n522 VSUBS 0.008128f
C1268 B.n523 VSUBS 0.008128f
C1269 B.n524 VSUBS 0.008128f
C1270 B.n525 VSUBS 0.008128f
C1271 B.n526 VSUBS 0.008128f
C1272 B.n527 VSUBS 0.008128f
C1273 B.n528 VSUBS 0.008128f
C1274 B.n529 VSUBS 0.008128f
C1275 B.n530 VSUBS 0.008128f
C1276 B.n531 VSUBS 0.008128f
C1277 B.n532 VSUBS 0.008128f
C1278 B.n533 VSUBS 0.008128f
C1279 B.n534 VSUBS 0.008128f
C1280 B.n535 VSUBS 0.008128f
C1281 B.n536 VSUBS 0.008128f
C1282 B.n537 VSUBS 0.008128f
C1283 B.n538 VSUBS 0.008128f
C1284 B.n539 VSUBS 0.008128f
C1285 B.n540 VSUBS 0.008128f
C1286 B.n541 VSUBS 0.008128f
C1287 B.n542 VSUBS 0.008128f
C1288 B.n543 VSUBS 0.008128f
C1289 B.n544 VSUBS 0.008128f
C1290 B.n545 VSUBS 0.008128f
C1291 B.n546 VSUBS 0.008128f
C1292 B.n547 VSUBS 0.008128f
C1293 B.n548 VSUBS 0.008128f
C1294 B.n549 VSUBS 0.008128f
C1295 B.n550 VSUBS 0.008128f
C1296 B.n551 VSUBS 0.008128f
C1297 B.n552 VSUBS 0.008128f
C1298 B.n553 VSUBS 0.008128f
C1299 B.n554 VSUBS 0.008128f
C1300 B.n555 VSUBS 0.008128f
C1301 B.n556 VSUBS 0.008128f
C1302 B.n557 VSUBS 0.008128f
C1303 B.n558 VSUBS 0.008128f
C1304 B.n559 VSUBS 0.008128f
C1305 B.n560 VSUBS 0.008128f
C1306 B.n561 VSUBS 0.008128f
C1307 B.n562 VSUBS 0.008128f
C1308 B.n563 VSUBS 0.008128f
C1309 B.n564 VSUBS 0.008128f
C1310 B.n565 VSUBS 0.008128f
C1311 B.n566 VSUBS 0.008128f
C1312 B.n567 VSUBS 0.008128f
C1313 B.n568 VSUBS 0.008128f
C1314 B.n569 VSUBS 0.008128f
C1315 B.n570 VSUBS 0.008128f
C1316 B.n571 VSUBS 0.008128f
C1317 B.n572 VSUBS 0.008128f
C1318 B.n573 VSUBS 0.008128f
C1319 B.n574 VSUBS 0.008128f
C1320 B.n575 VSUBS 0.008128f
C1321 B.n576 VSUBS 0.008128f
C1322 B.n577 VSUBS 0.008128f
C1323 B.n578 VSUBS 0.008128f
C1324 B.n579 VSUBS 0.008128f
C1325 B.n580 VSUBS 0.008128f
C1326 B.n581 VSUBS 0.008128f
C1327 B.n582 VSUBS 0.008128f
C1328 B.n583 VSUBS 0.008128f
C1329 B.n584 VSUBS 0.008128f
C1330 B.n585 VSUBS 0.008128f
C1331 B.n586 VSUBS 0.008128f
C1332 B.n587 VSUBS 0.008128f
C1333 B.n588 VSUBS 0.008128f
C1334 B.n589 VSUBS 0.008128f
C1335 B.n590 VSUBS 0.008128f
C1336 B.n591 VSUBS 0.008128f
C1337 B.n592 VSUBS 0.008128f
C1338 B.n593 VSUBS 0.008128f
C1339 B.n594 VSUBS 0.008128f
C1340 B.n595 VSUBS 0.008128f
C1341 B.n596 VSUBS 0.008128f
C1342 B.n597 VSUBS 0.008128f
C1343 B.n598 VSUBS 0.008128f
C1344 B.n599 VSUBS 0.008128f
C1345 B.n600 VSUBS 0.008128f
C1346 B.n601 VSUBS 0.008128f
C1347 B.n602 VSUBS 0.008128f
C1348 B.n603 VSUBS 0.008128f
C1349 B.n604 VSUBS 0.008128f
C1350 B.n605 VSUBS 0.008128f
C1351 B.n606 VSUBS 0.008128f
C1352 B.n607 VSUBS 0.008128f
C1353 B.n608 VSUBS 0.008128f
C1354 B.n609 VSUBS 0.008128f
C1355 B.n610 VSUBS 0.008128f
C1356 B.n611 VSUBS 0.008128f
C1357 B.n612 VSUBS 0.008128f
C1358 B.n613 VSUBS 0.008128f
C1359 B.n614 VSUBS 0.008128f
C1360 B.n615 VSUBS 0.008128f
C1361 B.n616 VSUBS 0.008128f
C1362 B.n617 VSUBS 0.008128f
C1363 B.n618 VSUBS 0.008128f
C1364 B.n619 VSUBS 0.008128f
C1365 B.n620 VSUBS 0.008128f
C1366 B.n621 VSUBS 0.008128f
C1367 B.n622 VSUBS 0.008128f
C1368 B.n623 VSUBS 0.008128f
C1369 B.n624 VSUBS 0.008128f
C1370 B.n625 VSUBS 0.008128f
C1371 B.n626 VSUBS 0.008128f
C1372 B.n627 VSUBS 0.019032f
C1373 B.n628 VSUBS 0.01995f
C1374 B.n629 VSUBS 0.019256f
C1375 B.n630 VSUBS 0.008128f
C1376 B.n631 VSUBS 0.008128f
C1377 B.n632 VSUBS 0.008128f
C1378 B.n633 VSUBS 0.008128f
C1379 B.n634 VSUBS 0.008128f
C1380 B.n635 VSUBS 0.008128f
C1381 B.n636 VSUBS 0.008128f
C1382 B.n637 VSUBS 0.008128f
C1383 B.n638 VSUBS 0.008128f
C1384 B.n639 VSUBS 0.008128f
C1385 B.n640 VSUBS 0.008128f
C1386 B.n641 VSUBS 0.008128f
C1387 B.n642 VSUBS 0.008128f
C1388 B.n643 VSUBS 0.008128f
C1389 B.n644 VSUBS 0.008128f
C1390 B.n645 VSUBS 0.008128f
C1391 B.n646 VSUBS 0.008128f
C1392 B.n647 VSUBS 0.008128f
C1393 B.n648 VSUBS 0.008128f
C1394 B.n649 VSUBS 0.008128f
C1395 B.n650 VSUBS 0.008128f
C1396 B.n651 VSUBS 0.008128f
C1397 B.n652 VSUBS 0.008128f
C1398 B.n653 VSUBS 0.008128f
C1399 B.n654 VSUBS 0.008128f
C1400 B.n655 VSUBS 0.008128f
C1401 B.n656 VSUBS 0.008128f
C1402 B.n657 VSUBS 0.008128f
C1403 B.n658 VSUBS 0.008128f
C1404 B.n659 VSUBS 0.008128f
C1405 B.n660 VSUBS 0.008128f
C1406 B.n661 VSUBS 0.008128f
C1407 B.n662 VSUBS 0.008128f
C1408 B.n663 VSUBS 0.008128f
C1409 B.n664 VSUBS 0.008128f
C1410 B.n665 VSUBS 0.008128f
C1411 B.n666 VSUBS 0.008128f
C1412 B.n667 VSUBS 0.008128f
C1413 B.n668 VSUBS 0.008128f
C1414 B.n669 VSUBS 0.008128f
C1415 B.n670 VSUBS 0.008128f
C1416 B.n671 VSUBS 0.008128f
C1417 B.n672 VSUBS 0.008128f
C1418 B.n673 VSUBS 0.008128f
C1419 B.n674 VSUBS 0.008128f
C1420 B.n675 VSUBS 0.008128f
C1421 B.n676 VSUBS 0.008128f
C1422 B.n677 VSUBS 0.008128f
C1423 B.n678 VSUBS 0.008128f
C1424 B.n679 VSUBS 0.008128f
C1425 B.n680 VSUBS 0.008128f
C1426 B.n681 VSUBS 0.008128f
C1427 B.n682 VSUBS 0.008128f
C1428 B.n683 VSUBS 0.008128f
C1429 B.n684 VSUBS 0.008128f
C1430 B.n685 VSUBS 0.008128f
C1431 B.n686 VSUBS 0.008128f
C1432 B.n687 VSUBS 0.008128f
C1433 B.n688 VSUBS 0.008128f
C1434 B.n689 VSUBS 0.008128f
C1435 B.n690 VSUBS 0.008128f
C1436 B.n691 VSUBS 0.008128f
C1437 B.n692 VSUBS 0.008128f
C1438 B.n693 VSUBS 0.008128f
C1439 B.n694 VSUBS 0.00765f
C1440 B.n695 VSUBS 0.018832f
C1441 B.n696 VSUBS 0.004542f
C1442 B.n697 VSUBS 0.008128f
C1443 B.n698 VSUBS 0.008128f
C1444 B.n699 VSUBS 0.008128f
C1445 B.n700 VSUBS 0.008128f
C1446 B.n701 VSUBS 0.008128f
C1447 B.n702 VSUBS 0.008128f
C1448 B.n703 VSUBS 0.008128f
C1449 B.n704 VSUBS 0.008128f
C1450 B.n705 VSUBS 0.008128f
C1451 B.n706 VSUBS 0.008128f
C1452 B.n707 VSUBS 0.008128f
C1453 B.n708 VSUBS 0.008128f
C1454 B.n709 VSUBS 0.004542f
C1455 B.n710 VSUBS 0.008128f
C1456 B.n711 VSUBS 0.008128f
C1457 B.n712 VSUBS 0.008128f
C1458 B.n713 VSUBS 0.008128f
C1459 B.n714 VSUBS 0.008128f
C1460 B.n715 VSUBS 0.008128f
C1461 B.n716 VSUBS 0.008128f
C1462 B.n717 VSUBS 0.008128f
C1463 B.n718 VSUBS 0.008128f
C1464 B.n719 VSUBS 0.008128f
C1465 B.n720 VSUBS 0.008128f
C1466 B.n721 VSUBS 0.008128f
C1467 B.n722 VSUBS 0.008128f
C1468 B.n723 VSUBS 0.008128f
C1469 B.n724 VSUBS 0.008128f
C1470 B.n725 VSUBS 0.008128f
C1471 B.n726 VSUBS 0.008128f
C1472 B.n727 VSUBS 0.008128f
C1473 B.n728 VSUBS 0.008128f
C1474 B.n729 VSUBS 0.008128f
C1475 B.n730 VSUBS 0.008128f
C1476 B.n731 VSUBS 0.008128f
C1477 B.n732 VSUBS 0.008128f
C1478 B.n733 VSUBS 0.008128f
C1479 B.n734 VSUBS 0.008128f
C1480 B.n735 VSUBS 0.008128f
C1481 B.n736 VSUBS 0.008128f
C1482 B.n737 VSUBS 0.008128f
C1483 B.n738 VSUBS 0.008128f
C1484 B.n739 VSUBS 0.008128f
C1485 B.n740 VSUBS 0.008128f
C1486 B.n741 VSUBS 0.008128f
C1487 B.n742 VSUBS 0.008128f
C1488 B.n743 VSUBS 0.008128f
C1489 B.n744 VSUBS 0.008128f
C1490 B.n745 VSUBS 0.008128f
C1491 B.n746 VSUBS 0.008128f
C1492 B.n747 VSUBS 0.008128f
C1493 B.n748 VSUBS 0.008128f
C1494 B.n749 VSUBS 0.008128f
C1495 B.n750 VSUBS 0.008128f
C1496 B.n751 VSUBS 0.008128f
C1497 B.n752 VSUBS 0.008128f
C1498 B.n753 VSUBS 0.008128f
C1499 B.n754 VSUBS 0.008128f
C1500 B.n755 VSUBS 0.008128f
C1501 B.n756 VSUBS 0.008128f
C1502 B.n757 VSUBS 0.008128f
C1503 B.n758 VSUBS 0.008128f
C1504 B.n759 VSUBS 0.008128f
C1505 B.n760 VSUBS 0.008128f
C1506 B.n761 VSUBS 0.008128f
C1507 B.n762 VSUBS 0.008128f
C1508 B.n763 VSUBS 0.008128f
C1509 B.n764 VSUBS 0.008128f
C1510 B.n765 VSUBS 0.008128f
C1511 B.n766 VSUBS 0.008128f
C1512 B.n767 VSUBS 0.008128f
C1513 B.n768 VSUBS 0.008128f
C1514 B.n769 VSUBS 0.008128f
C1515 B.n770 VSUBS 0.008128f
C1516 B.n771 VSUBS 0.008128f
C1517 B.n772 VSUBS 0.008128f
C1518 B.n773 VSUBS 0.008128f
C1519 B.n774 VSUBS 0.008128f
C1520 B.n775 VSUBS 0.020174f
C1521 B.n776 VSUBS 0.020174f
C1522 B.n777 VSUBS 0.019032f
C1523 B.n778 VSUBS 0.008128f
C1524 B.n779 VSUBS 0.008128f
C1525 B.n780 VSUBS 0.008128f
C1526 B.n781 VSUBS 0.008128f
C1527 B.n782 VSUBS 0.008128f
C1528 B.n783 VSUBS 0.008128f
C1529 B.n784 VSUBS 0.008128f
C1530 B.n785 VSUBS 0.008128f
C1531 B.n786 VSUBS 0.008128f
C1532 B.n787 VSUBS 0.008128f
C1533 B.n788 VSUBS 0.008128f
C1534 B.n789 VSUBS 0.008128f
C1535 B.n790 VSUBS 0.008128f
C1536 B.n791 VSUBS 0.008128f
C1537 B.n792 VSUBS 0.008128f
C1538 B.n793 VSUBS 0.008128f
C1539 B.n794 VSUBS 0.008128f
C1540 B.n795 VSUBS 0.008128f
C1541 B.n796 VSUBS 0.008128f
C1542 B.n797 VSUBS 0.008128f
C1543 B.n798 VSUBS 0.008128f
C1544 B.n799 VSUBS 0.008128f
C1545 B.n800 VSUBS 0.008128f
C1546 B.n801 VSUBS 0.008128f
C1547 B.n802 VSUBS 0.008128f
C1548 B.n803 VSUBS 0.008128f
C1549 B.n804 VSUBS 0.008128f
C1550 B.n805 VSUBS 0.008128f
C1551 B.n806 VSUBS 0.008128f
C1552 B.n807 VSUBS 0.008128f
C1553 B.n808 VSUBS 0.008128f
C1554 B.n809 VSUBS 0.008128f
C1555 B.n810 VSUBS 0.008128f
C1556 B.n811 VSUBS 0.008128f
C1557 B.n812 VSUBS 0.008128f
C1558 B.n813 VSUBS 0.008128f
C1559 B.n814 VSUBS 0.008128f
C1560 B.n815 VSUBS 0.008128f
C1561 B.n816 VSUBS 0.008128f
C1562 B.n817 VSUBS 0.008128f
C1563 B.n818 VSUBS 0.008128f
C1564 B.n819 VSUBS 0.008128f
C1565 B.n820 VSUBS 0.008128f
C1566 B.n821 VSUBS 0.008128f
C1567 B.n822 VSUBS 0.008128f
C1568 B.n823 VSUBS 0.008128f
C1569 B.n824 VSUBS 0.008128f
C1570 B.n825 VSUBS 0.008128f
C1571 B.n826 VSUBS 0.008128f
C1572 B.n827 VSUBS 0.008128f
C1573 B.n828 VSUBS 0.008128f
C1574 B.n829 VSUBS 0.008128f
C1575 B.n830 VSUBS 0.008128f
C1576 B.n831 VSUBS 0.008128f
C1577 B.n832 VSUBS 0.008128f
C1578 B.n833 VSUBS 0.008128f
C1579 B.n834 VSUBS 0.008128f
C1580 B.n835 VSUBS 0.008128f
C1581 B.n836 VSUBS 0.008128f
C1582 B.n837 VSUBS 0.008128f
C1583 B.n838 VSUBS 0.008128f
C1584 B.n839 VSUBS 0.008128f
C1585 B.n840 VSUBS 0.008128f
C1586 B.n841 VSUBS 0.008128f
C1587 B.n842 VSUBS 0.008128f
C1588 B.n843 VSUBS 0.008128f
C1589 B.n844 VSUBS 0.008128f
C1590 B.n845 VSUBS 0.008128f
C1591 B.n846 VSUBS 0.008128f
C1592 B.n847 VSUBS 0.008128f
C1593 B.n848 VSUBS 0.008128f
C1594 B.n849 VSUBS 0.008128f
C1595 B.n850 VSUBS 0.008128f
C1596 B.n851 VSUBS 0.008128f
C1597 B.n852 VSUBS 0.008128f
C1598 B.n853 VSUBS 0.008128f
C1599 B.n854 VSUBS 0.008128f
C1600 B.n855 VSUBS 0.008128f
C1601 B.n856 VSUBS 0.008128f
C1602 B.n857 VSUBS 0.008128f
C1603 B.n858 VSUBS 0.008128f
C1604 B.n859 VSUBS 0.008128f
C1605 B.n860 VSUBS 0.008128f
C1606 B.n861 VSUBS 0.008128f
C1607 B.n862 VSUBS 0.008128f
C1608 B.n863 VSUBS 0.018405f
.ends

