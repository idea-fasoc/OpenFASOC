* NGSPICE file created from diff_pair_sample_0645.ext - technology: sky130A

.subckt diff_pair_sample_0645 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t8 w_n3906_n4216# sky130_fd_pr__pfet_01v8 ad=2.6796 pd=16.57 as=6.3336 ps=33.26 w=16.24 l=3.34
X1 VDD2.t5 VN.t0 VTAIL.t11 w_n3906_n4216# sky130_fd_pr__pfet_01v8 ad=6.3336 pd=33.26 as=2.6796 ps=16.57 w=16.24 l=3.34
X2 B.t11 B.t9 B.t10 w_n3906_n4216# sky130_fd_pr__pfet_01v8 ad=6.3336 pd=33.26 as=0 ps=0 w=16.24 l=3.34
X3 VTAIL.t0 VN.t1 VDD2.t4 w_n3906_n4216# sky130_fd_pr__pfet_01v8 ad=2.6796 pd=16.57 as=2.6796 ps=16.57 w=16.24 l=3.34
X4 VTAIL.t5 VP.t1 VDD1.t4 w_n3906_n4216# sky130_fd_pr__pfet_01v8 ad=2.6796 pd=16.57 as=2.6796 ps=16.57 w=16.24 l=3.34
X5 VTAIL.t3 VN.t2 VDD2.t3 w_n3906_n4216# sky130_fd_pr__pfet_01v8 ad=2.6796 pd=16.57 as=2.6796 ps=16.57 w=16.24 l=3.34
X6 B.t8 B.t6 B.t7 w_n3906_n4216# sky130_fd_pr__pfet_01v8 ad=6.3336 pd=33.26 as=0 ps=0 w=16.24 l=3.34
X7 VTAIL.t9 VP.t2 VDD1.t3 w_n3906_n4216# sky130_fd_pr__pfet_01v8 ad=2.6796 pd=16.57 as=2.6796 ps=16.57 w=16.24 l=3.34
X8 VDD2.t2 VN.t3 VTAIL.t1 w_n3906_n4216# sky130_fd_pr__pfet_01v8 ad=2.6796 pd=16.57 as=6.3336 ps=33.26 w=16.24 l=3.34
X9 VDD2.t1 VN.t4 VTAIL.t4 w_n3906_n4216# sky130_fd_pr__pfet_01v8 ad=6.3336 pd=33.26 as=2.6796 ps=16.57 w=16.24 l=3.34
X10 VDD2.t0 VN.t5 VTAIL.t2 w_n3906_n4216# sky130_fd_pr__pfet_01v8 ad=2.6796 pd=16.57 as=6.3336 ps=33.26 w=16.24 l=3.34
X11 B.t5 B.t3 B.t4 w_n3906_n4216# sky130_fd_pr__pfet_01v8 ad=6.3336 pd=33.26 as=0 ps=0 w=16.24 l=3.34
X12 VDD1.t2 VP.t3 VTAIL.t6 w_n3906_n4216# sky130_fd_pr__pfet_01v8 ad=6.3336 pd=33.26 as=2.6796 ps=16.57 w=16.24 l=3.34
X13 VDD1.t1 VP.t4 VTAIL.t10 w_n3906_n4216# sky130_fd_pr__pfet_01v8 ad=6.3336 pd=33.26 as=2.6796 ps=16.57 w=16.24 l=3.34
X14 VDD1.t0 VP.t5 VTAIL.t7 w_n3906_n4216# sky130_fd_pr__pfet_01v8 ad=2.6796 pd=16.57 as=6.3336 ps=33.26 w=16.24 l=3.34
X15 B.t2 B.t0 B.t1 w_n3906_n4216# sky130_fd_pr__pfet_01v8 ad=6.3336 pd=33.26 as=0 ps=0 w=16.24 l=3.34
R0 VP.n16 VP.n15 161.3
R1 VP.n17 VP.n12 161.3
R2 VP.n19 VP.n18 161.3
R3 VP.n20 VP.n11 161.3
R4 VP.n22 VP.n21 161.3
R5 VP.n23 VP.n10 161.3
R6 VP.n25 VP.n24 161.3
R7 VP.n50 VP.n49 161.3
R8 VP.n48 VP.n1 161.3
R9 VP.n47 VP.n46 161.3
R10 VP.n45 VP.n2 161.3
R11 VP.n44 VP.n43 161.3
R12 VP.n42 VP.n3 161.3
R13 VP.n41 VP.n40 161.3
R14 VP.n39 VP.n4 161.3
R15 VP.n38 VP.n37 161.3
R16 VP.n36 VP.n5 161.3
R17 VP.n35 VP.n34 161.3
R18 VP.n33 VP.n6 161.3
R19 VP.n32 VP.n31 161.3
R20 VP.n30 VP.n7 161.3
R21 VP.n29 VP.n28 161.3
R22 VP.n14 VP.t4 150.376
R23 VP.n4 VP.t1 117.181
R24 VP.n8 VP.t3 117.181
R25 VP.n0 VP.t5 117.181
R26 VP.n13 VP.t2 117.181
R27 VP.n9 VP.t0 117.181
R28 VP.n27 VP.n8 81.8843
R29 VP.n51 VP.n0 81.8843
R30 VP.n26 VP.n9 81.8843
R31 VP.n35 VP.n6 56.5617
R32 VP.n43 VP.n2 56.5617
R33 VP.n18 VP.n11 56.5617
R34 VP.n27 VP.n26 54.8139
R35 VP.n14 VP.n13 50.1906
R36 VP.n30 VP.n29 24.5923
R37 VP.n31 VP.n30 24.5923
R38 VP.n31 VP.n6 24.5923
R39 VP.n36 VP.n35 24.5923
R40 VP.n37 VP.n36 24.5923
R41 VP.n37 VP.n4 24.5923
R42 VP.n41 VP.n4 24.5923
R43 VP.n42 VP.n41 24.5923
R44 VP.n43 VP.n42 24.5923
R45 VP.n47 VP.n2 24.5923
R46 VP.n48 VP.n47 24.5923
R47 VP.n49 VP.n48 24.5923
R48 VP.n22 VP.n11 24.5923
R49 VP.n23 VP.n22 24.5923
R50 VP.n24 VP.n23 24.5923
R51 VP.n16 VP.n13 24.5923
R52 VP.n17 VP.n16 24.5923
R53 VP.n18 VP.n17 24.5923
R54 VP.n29 VP.n8 8.36172
R55 VP.n49 VP.n0 8.36172
R56 VP.n24 VP.n9 8.36172
R57 VP.n15 VP.n14 3.19892
R58 VP.n26 VP.n25 0.354861
R59 VP.n28 VP.n27 0.354861
R60 VP.n51 VP.n50 0.354861
R61 VP VP.n51 0.267071
R62 VP.n15 VP.n12 0.189894
R63 VP.n19 VP.n12 0.189894
R64 VP.n20 VP.n19 0.189894
R65 VP.n21 VP.n20 0.189894
R66 VP.n21 VP.n10 0.189894
R67 VP.n25 VP.n10 0.189894
R68 VP.n28 VP.n7 0.189894
R69 VP.n32 VP.n7 0.189894
R70 VP.n33 VP.n32 0.189894
R71 VP.n34 VP.n33 0.189894
R72 VP.n34 VP.n5 0.189894
R73 VP.n38 VP.n5 0.189894
R74 VP.n39 VP.n38 0.189894
R75 VP.n40 VP.n39 0.189894
R76 VP.n40 VP.n3 0.189894
R77 VP.n44 VP.n3 0.189894
R78 VP.n45 VP.n44 0.189894
R79 VP.n46 VP.n45 0.189894
R80 VP.n46 VP.n1 0.189894
R81 VP.n50 VP.n1 0.189894
R82 VTAIL.n362 VTAIL.n278 756.745
R83 VTAIL.n86 VTAIL.n2 756.745
R84 VTAIL.n272 VTAIL.n188 756.745
R85 VTAIL.n180 VTAIL.n96 756.745
R86 VTAIL.n306 VTAIL.n305 585
R87 VTAIL.n311 VTAIL.n310 585
R88 VTAIL.n313 VTAIL.n312 585
R89 VTAIL.n302 VTAIL.n301 585
R90 VTAIL.n319 VTAIL.n318 585
R91 VTAIL.n321 VTAIL.n320 585
R92 VTAIL.n298 VTAIL.n297 585
R93 VTAIL.n327 VTAIL.n326 585
R94 VTAIL.n329 VTAIL.n328 585
R95 VTAIL.n294 VTAIL.n293 585
R96 VTAIL.n335 VTAIL.n334 585
R97 VTAIL.n337 VTAIL.n336 585
R98 VTAIL.n290 VTAIL.n289 585
R99 VTAIL.n343 VTAIL.n342 585
R100 VTAIL.n345 VTAIL.n344 585
R101 VTAIL.n286 VTAIL.n285 585
R102 VTAIL.n352 VTAIL.n351 585
R103 VTAIL.n353 VTAIL.n284 585
R104 VTAIL.n355 VTAIL.n354 585
R105 VTAIL.n282 VTAIL.n281 585
R106 VTAIL.n361 VTAIL.n360 585
R107 VTAIL.n363 VTAIL.n362 585
R108 VTAIL.n30 VTAIL.n29 585
R109 VTAIL.n35 VTAIL.n34 585
R110 VTAIL.n37 VTAIL.n36 585
R111 VTAIL.n26 VTAIL.n25 585
R112 VTAIL.n43 VTAIL.n42 585
R113 VTAIL.n45 VTAIL.n44 585
R114 VTAIL.n22 VTAIL.n21 585
R115 VTAIL.n51 VTAIL.n50 585
R116 VTAIL.n53 VTAIL.n52 585
R117 VTAIL.n18 VTAIL.n17 585
R118 VTAIL.n59 VTAIL.n58 585
R119 VTAIL.n61 VTAIL.n60 585
R120 VTAIL.n14 VTAIL.n13 585
R121 VTAIL.n67 VTAIL.n66 585
R122 VTAIL.n69 VTAIL.n68 585
R123 VTAIL.n10 VTAIL.n9 585
R124 VTAIL.n76 VTAIL.n75 585
R125 VTAIL.n77 VTAIL.n8 585
R126 VTAIL.n79 VTAIL.n78 585
R127 VTAIL.n6 VTAIL.n5 585
R128 VTAIL.n85 VTAIL.n84 585
R129 VTAIL.n87 VTAIL.n86 585
R130 VTAIL.n273 VTAIL.n272 585
R131 VTAIL.n271 VTAIL.n270 585
R132 VTAIL.n192 VTAIL.n191 585
R133 VTAIL.n265 VTAIL.n264 585
R134 VTAIL.n263 VTAIL.n194 585
R135 VTAIL.n262 VTAIL.n261 585
R136 VTAIL.n197 VTAIL.n195 585
R137 VTAIL.n256 VTAIL.n255 585
R138 VTAIL.n254 VTAIL.n253 585
R139 VTAIL.n201 VTAIL.n200 585
R140 VTAIL.n248 VTAIL.n247 585
R141 VTAIL.n246 VTAIL.n245 585
R142 VTAIL.n205 VTAIL.n204 585
R143 VTAIL.n240 VTAIL.n239 585
R144 VTAIL.n238 VTAIL.n237 585
R145 VTAIL.n209 VTAIL.n208 585
R146 VTAIL.n232 VTAIL.n231 585
R147 VTAIL.n230 VTAIL.n229 585
R148 VTAIL.n213 VTAIL.n212 585
R149 VTAIL.n224 VTAIL.n223 585
R150 VTAIL.n222 VTAIL.n221 585
R151 VTAIL.n217 VTAIL.n216 585
R152 VTAIL.n181 VTAIL.n180 585
R153 VTAIL.n179 VTAIL.n178 585
R154 VTAIL.n100 VTAIL.n99 585
R155 VTAIL.n173 VTAIL.n172 585
R156 VTAIL.n171 VTAIL.n102 585
R157 VTAIL.n170 VTAIL.n169 585
R158 VTAIL.n105 VTAIL.n103 585
R159 VTAIL.n164 VTAIL.n163 585
R160 VTAIL.n162 VTAIL.n161 585
R161 VTAIL.n109 VTAIL.n108 585
R162 VTAIL.n156 VTAIL.n155 585
R163 VTAIL.n154 VTAIL.n153 585
R164 VTAIL.n113 VTAIL.n112 585
R165 VTAIL.n148 VTAIL.n147 585
R166 VTAIL.n146 VTAIL.n145 585
R167 VTAIL.n117 VTAIL.n116 585
R168 VTAIL.n140 VTAIL.n139 585
R169 VTAIL.n138 VTAIL.n137 585
R170 VTAIL.n121 VTAIL.n120 585
R171 VTAIL.n132 VTAIL.n131 585
R172 VTAIL.n130 VTAIL.n129 585
R173 VTAIL.n125 VTAIL.n124 585
R174 VTAIL.n307 VTAIL.t2 327.466
R175 VTAIL.n31 VTAIL.t7 327.466
R176 VTAIL.n218 VTAIL.t8 327.466
R177 VTAIL.n126 VTAIL.t1 327.466
R178 VTAIL.n311 VTAIL.n305 171.744
R179 VTAIL.n312 VTAIL.n311 171.744
R180 VTAIL.n312 VTAIL.n301 171.744
R181 VTAIL.n319 VTAIL.n301 171.744
R182 VTAIL.n320 VTAIL.n319 171.744
R183 VTAIL.n320 VTAIL.n297 171.744
R184 VTAIL.n327 VTAIL.n297 171.744
R185 VTAIL.n328 VTAIL.n327 171.744
R186 VTAIL.n328 VTAIL.n293 171.744
R187 VTAIL.n335 VTAIL.n293 171.744
R188 VTAIL.n336 VTAIL.n335 171.744
R189 VTAIL.n336 VTAIL.n289 171.744
R190 VTAIL.n343 VTAIL.n289 171.744
R191 VTAIL.n344 VTAIL.n343 171.744
R192 VTAIL.n344 VTAIL.n285 171.744
R193 VTAIL.n352 VTAIL.n285 171.744
R194 VTAIL.n353 VTAIL.n352 171.744
R195 VTAIL.n354 VTAIL.n353 171.744
R196 VTAIL.n354 VTAIL.n281 171.744
R197 VTAIL.n361 VTAIL.n281 171.744
R198 VTAIL.n362 VTAIL.n361 171.744
R199 VTAIL.n35 VTAIL.n29 171.744
R200 VTAIL.n36 VTAIL.n35 171.744
R201 VTAIL.n36 VTAIL.n25 171.744
R202 VTAIL.n43 VTAIL.n25 171.744
R203 VTAIL.n44 VTAIL.n43 171.744
R204 VTAIL.n44 VTAIL.n21 171.744
R205 VTAIL.n51 VTAIL.n21 171.744
R206 VTAIL.n52 VTAIL.n51 171.744
R207 VTAIL.n52 VTAIL.n17 171.744
R208 VTAIL.n59 VTAIL.n17 171.744
R209 VTAIL.n60 VTAIL.n59 171.744
R210 VTAIL.n60 VTAIL.n13 171.744
R211 VTAIL.n67 VTAIL.n13 171.744
R212 VTAIL.n68 VTAIL.n67 171.744
R213 VTAIL.n68 VTAIL.n9 171.744
R214 VTAIL.n76 VTAIL.n9 171.744
R215 VTAIL.n77 VTAIL.n76 171.744
R216 VTAIL.n78 VTAIL.n77 171.744
R217 VTAIL.n78 VTAIL.n5 171.744
R218 VTAIL.n85 VTAIL.n5 171.744
R219 VTAIL.n86 VTAIL.n85 171.744
R220 VTAIL.n272 VTAIL.n271 171.744
R221 VTAIL.n271 VTAIL.n191 171.744
R222 VTAIL.n264 VTAIL.n191 171.744
R223 VTAIL.n264 VTAIL.n263 171.744
R224 VTAIL.n263 VTAIL.n262 171.744
R225 VTAIL.n262 VTAIL.n195 171.744
R226 VTAIL.n255 VTAIL.n195 171.744
R227 VTAIL.n255 VTAIL.n254 171.744
R228 VTAIL.n254 VTAIL.n200 171.744
R229 VTAIL.n247 VTAIL.n200 171.744
R230 VTAIL.n247 VTAIL.n246 171.744
R231 VTAIL.n246 VTAIL.n204 171.744
R232 VTAIL.n239 VTAIL.n204 171.744
R233 VTAIL.n239 VTAIL.n238 171.744
R234 VTAIL.n238 VTAIL.n208 171.744
R235 VTAIL.n231 VTAIL.n208 171.744
R236 VTAIL.n231 VTAIL.n230 171.744
R237 VTAIL.n230 VTAIL.n212 171.744
R238 VTAIL.n223 VTAIL.n212 171.744
R239 VTAIL.n223 VTAIL.n222 171.744
R240 VTAIL.n222 VTAIL.n216 171.744
R241 VTAIL.n180 VTAIL.n179 171.744
R242 VTAIL.n179 VTAIL.n99 171.744
R243 VTAIL.n172 VTAIL.n99 171.744
R244 VTAIL.n172 VTAIL.n171 171.744
R245 VTAIL.n171 VTAIL.n170 171.744
R246 VTAIL.n170 VTAIL.n103 171.744
R247 VTAIL.n163 VTAIL.n103 171.744
R248 VTAIL.n163 VTAIL.n162 171.744
R249 VTAIL.n162 VTAIL.n108 171.744
R250 VTAIL.n155 VTAIL.n108 171.744
R251 VTAIL.n155 VTAIL.n154 171.744
R252 VTAIL.n154 VTAIL.n112 171.744
R253 VTAIL.n147 VTAIL.n112 171.744
R254 VTAIL.n147 VTAIL.n146 171.744
R255 VTAIL.n146 VTAIL.n116 171.744
R256 VTAIL.n139 VTAIL.n116 171.744
R257 VTAIL.n139 VTAIL.n138 171.744
R258 VTAIL.n138 VTAIL.n120 171.744
R259 VTAIL.n131 VTAIL.n120 171.744
R260 VTAIL.n131 VTAIL.n130 171.744
R261 VTAIL.n130 VTAIL.n124 171.744
R262 VTAIL.t2 VTAIL.n305 85.8723
R263 VTAIL.t7 VTAIL.n29 85.8723
R264 VTAIL.t8 VTAIL.n216 85.8723
R265 VTAIL.t1 VTAIL.n124 85.8723
R266 VTAIL.n187 VTAIL.n186 56.2264
R267 VTAIL.n95 VTAIL.n94 56.2264
R268 VTAIL.n1 VTAIL.n0 56.2262
R269 VTAIL.n93 VTAIL.n92 56.2262
R270 VTAIL.n367 VTAIL.n366 35.2884
R271 VTAIL.n91 VTAIL.n90 35.2884
R272 VTAIL.n277 VTAIL.n276 35.2884
R273 VTAIL.n185 VTAIL.n184 35.2884
R274 VTAIL.n95 VTAIL.n93 32.6945
R275 VTAIL.n367 VTAIL.n277 29.5307
R276 VTAIL.n307 VTAIL.n306 16.3895
R277 VTAIL.n31 VTAIL.n30 16.3895
R278 VTAIL.n218 VTAIL.n217 16.3895
R279 VTAIL.n126 VTAIL.n125 16.3895
R280 VTAIL.n355 VTAIL.n284 13.1884
R281 VTAIL.n79 VTAIL.n8 13.1884
R282 VTAIL.n265 VTAIL.n194 13.1884
R283 VTAIL.n173 VTAIL.n102 13.1884
R284 VTAIL.n310 VTAIL.n309 12.8005
R285 VTAIL.n351 VTAIL.n350 12.8005
R286 VTAIL.n356 VTAIL.n282 12.8005
R287 VTAIL.n34 VTAIL.n33 12.8005
R288 VTAIL.n75 VTAIL.n74 12.8005
R289 VTAIL.n80 VTAIL.n6 12.8005
R290 VTAIL.n266 VTAIL.n192 12.8005
R291 VTAIL.n261 VTAIL.n196 12.8005
R292 VTAIL.n221 VTAIL.n220 12.8005
R293 VTAIL.n174 VTAIL.n100 12.8005
R294 VTAIL.n169 VTAIL.n104 12.8005
R295 VTAIL.n129 VTAIL.n128 12.8005
R296 VTAIL.n313 VTAIL.n304 12.0247
R297 VTAIL.n349 VTAIL.n286 12.0247
R298 VTAIL.n360 VTAIL.n359 12.0247
R299 VTAIL.n37 VTAIL.n28 12.0247
R300 VTAIL.n73 VTAIL.n10 12.0247
R301 VTAIL.n84 VTAIL.n83 12.0247
R302 VTAIL.n270 VTAIL.n269 12.0247
R303 VTAIL.n260 VTAIL.n197 12.0247
R304 VTAIL.n224 VTAIL.n215 12.0247
R305 VTAIL.n178 VTAIL.n177 12.0247
R306 VTAIL.n168 VTAIL.n105 12.0247
R307 VTAIL.n132 VTAIL.n123 12.0247
R308 VTAIL.n314 VTAIL.n302 11.249
R309 VTAIL.n346 VTAIL.n345 11.249
R310 VTAIL.n363 VTAIL.n280 11.249
R311 VTAIL.n38 VTAIL.n26 11.249
R312 VTAIL.n70 VTAIL.n69 11.249
R313 VTAIL.n87 VTAIL.n4 11.249
R314 VTAIL.n273 VTAIL.n190 11.249
R315 VTAIL.n257 VTAIL.n256 11.249
R316 VTAIL.n225 VTAIL.n213 11.249
R317 VTAIL.n181 VTAIL.n98 11.249
R318 VTAIL.n165 VTAIL.n164 11.249
R319 VTAIL.n133 VTAIL.n121 11.249
R320 VTAIL.n318 VTAIL.n317 10.4732
R321 VTAIL.n342 VTAIL.n288 10.4732
R322 VTAIL.n364 VTAIL.n278 10.4732
R323 VTAIL.n42 VTAIL.n41 10.4732
R324 VTAIL.n66 VTAIL.n12 10.4732
R325 VTAIL.n88 VTAIL.n2 10.4732
R326 VTAIL.n274 VTAIL.n188 10.4732
R327 VTAIL.n253 VTAIL.n199 10.4732
R328 VTAIL.n229 VTAIL.n228 10.4732
R329 VTAIL.n182 VTAIL.n96 10.4732
R330 VTAIL.n161 VTAIL.n107 10.4732
R331 VTAIL.n137 VTAIL.n136 10.4732
R332 VTAIL.n321 VTAIL.n300 9.69747
R333 VTAIL.n341 VTAIL.n290 9.69747
R334 VTAIL.n45 VTAIL.n24 9.69747
R335 VTAIL.n65 VTAIL.n14 9.69747
R336 VTAIL.n252 VTAIL.n201 9.69747
R337 VTAIL.n232 VTAIL.n211 9.69747
R338 VTAIL.n160 VTAIL.n109 9.69747
R339 VTAIL.n140 VTAIL.n119 9.69747
R340 VTAIL.n366 VTAIL.n365 9.45567
R341 VTAIL.n90 VTAIL.n89 9.45567
R342 VTAIL.n276 VTAIL.n275 9.45567
R343 VTAIL.n184 VTAIL.n183 9.45567
R344 VTAIL.n365 VTAIL.n364 9.3005
R345 VTAIL.n280 VTAIL.n279 9.3005
R346 VTAIL.n359 VTAIL.n358 9.3005
R347 VTAIL.n357 VTAIL.n356 9.3005
R348 VTAIL.n296 VTAIL.n295 9.3005
R349 VTAIL.n325 VTAIL.n324 9.3005
R350 VTAIL.n323 VTAIL.n322 9.3005
R351 VTAIL.n300 VTAIL.n299 9.3005
R352 VTAIL.n317 VTAIL.n316 9.3005
R353 VTAIL.n315 VTAIL.n314 9.3005
R354 VTAIL.n304 VTAIL.n303 9.3005
R355 VTAIL.n309 VTAIL.n308 9.3005
R356 VTAIL.n331 VTAIL.n330 9.3005
R357 VTAIL.n333 VTAIL.n332 9.3005
R358 VTAIL.n292 VTAIL.n291 9.3005
R359 VTAIL.n339 VTAIL.n338 9.3005
R360 VTAIL.n341 VTAIL.n340 9.3005
R361 VTAIL.n288 VTAIL.n287 9.3005
R362 VTAIL.n347 VTAIL.n346 9.3005
R363 VTAIL.n349 VTAIL.n348 9.3005
R364 VTAIL.n350 VTAIL.n283 9.3005
R365 VTAIL.n89 VTAIL.n88 9.3005
R366 VTAIL.n4 VTAIL.n3 9.3005
R367 VTAIL.n83 VTAIL.n82 9.3005
R368 VTAIL.n81 VTAIL.n80 9.3005
R369 VTAIL.n20 VTAIL.n19 9.3005
R370 VTAIL.n49 VTAIL.n48 9.3005
R371 VTAIL.n47 VTAIL.n46 9.3005
R372 VTAIL.n24 VTAIL.n23 9.3005
R373 VTAIL.n41 VTAIL.n40 9.3005
R374 VTAIL.n39 VTAIL.n38 9.3005
R375 VTAIL.n28 VTAIL.n27 9.3005
R376 VTAIL.n33 VTAIL.n32 9.3005
R377 VTAIL.n55 VTAIL.n54 9.3005
R378 VTAIL.n57 VTAIL.n56 9.3005
R379 VTAIL.n16 VTAIL.n15 9.3005
R380 VTAIL.n63 VTAIL.n62 9.3005
R381 VTAIL.n65 VTAIL.n64 9.3005
R382 VTAIL.n12 VTAIL.n11 9.3005
R383 VTAIL.n71 VTAIL.n70 9.3005
R384 VTAIL.n73 VTAIL.n72 9.3005
R385 VTAIL.n74 VTAIL.n7 9.3005
R386 VTAIL.n244 VTAIL.n243 9.3005
R387 VTAIL.n203 VTAIL.n202 9.3005
R388 VTAIL.n250 VTAIL.n249 9.3005
R389 VTAIL.n252 VTAIL.n251 9.3005
R390 VTAIL.n199 VTAIL.n198 9.3005
R391 VTAIL.n258 VTAIL.n257 9.3005
R392 VTAIL.n260 VTAIL.n259 9.3005
R393 VTAIL.n196 VTAIL.n193 9.3005
R394 VTAIL.n275 VTAIL.n274 9.3005
R395 VTAIL.n190 VTAIL.n189 9.3005
R396 VTAIL.n269 VTAIL.n268 9.3005
R397 VTAIL.n267 VTAIL.n266 9.3005
R398 VTAIL.n242 VTAIL.n241 9.3005
R399 VTAIL.n207 VTAIL.n206 9.3005
R400 VTAIL.n236 VTAIL.n235 9.3005
R401 VTAIL.n234 VTAIL.n233 9.3005
R402 VTAIL.n211 VTAIL.n210 9.3005
R403 VTAIL.n228 VTAIL.n227 9.3005
R404 VTAIL.n226 VTAIL.n225 9.3005
R405 VTAIL.n215 VTAIL.n214 9.3005
R406 VTAIL.n220 VTAIL.n219 9.3005
R407 VTAIL.n152 VTAIL.n151 9.3005
R408 VTAIL.n111 VTAIL.n110 9.3005
R409 VTAIL.n158 VTAIL.n157 9.3005
R410 VTAIL.n160 VTAIL.n159 9.3005
R411 VTAIL.n107 VTAIL.n106 9.3005
R412 VTAIL.n166 VTAIL.n165 9.3005
R413 VTAIL.n168 VTAIL.n167 9.3005
R414 VTAIL.n104 VTAIL.n101 9.3005
R415 VTAIL.n183 VTAIL.n182 9.3005
R416 VTAIL.n98 VTAIL.n97 9.3005
R417 VTAIL.n177 VTAIL.n176 9.3005
R418 VTAIL.n175 VTAIL.n174 9.3005
R419 VTAIL.n150 VTAIL.n149 9.3005
R420 VTAIL.n115 VTAIL.n114 9.3005
R421 VTAIL.n144 VTAIL.n143 9.3005
R422 VTAIL.n142 VTAIL.n141 9.3005
R423 VTAIL.n119 VTAIL.n118 9.3005
R424 VTAIL.n136 VTAIL.n135 9.3005
R425 VTAIL.n134 VTAIL.n133 9.3005
R426 VTAIL.n123 VTAIL.n122 9.3005
R427 VTAIL.n128 VTAIL.n127 9.3005
R428 VTAIL.n322 VTAIL.n298 8.92171
R429 VTAIL.n338 VTAIL.n337 8.92171
R430 VTAIL.n46 VTAIL.n22 8.92171
R431 VTAIL.n62 VTAIL.n61 8.92171
R432 VTAIL.n249 VTAIL.n248 8.92171
R433 VTAIL.n233 VTAIL.n209 8.92171
R434 VTAIL.n157 VTAIL.n156 8.92171
R435 VTAIL.n141 VTAIL.n117 8.92171
R436 VTAIL.n326 VTAIL.n325 8.14595
R437 VTAIL.n334 VTAIL.n292 8.14595
R438 VTAIL.n50 VTAIL.n49 8.14595
R439 VTAIL.n58 VTAIL.n16 8.14595
R440 VTAIL.n245 VTAIL.n203 8.14595
R441 VTAIL.n237 VTAIL.n236 8.14595
R442 VTAIL.n153 VTAIL.n111 8.14595
R443 VTAIL.n145 VTAIL.n144 8.14595
R444 VTAIL.n329 VTAIL.n296 7.3702
R445 VTAIL.n333 VTAIL.n294 7.3702
R446 VTAIL.n53 VTAIL.n20 7.3702
R447 VTAIL.n57 VTAIL.n18 7.3702
R448 VTAIL.n244 VTAIL.n205 7.3702
R449 VTAIL.n240 VTAIL.n207 7.3702
R450 VTAIL.n152 VTAIL.n113 7.3702
R451 VTAIL.n148 VTAIL.n115 7.3702
R452 VTAIL.n330 VTAIL.n329 6.59444
R453 VTAIL.n330 VTAIL.n294 6.59444
R454 VTAIL.n54 VTAIL.n53 6.59444
R455 VTAIL.n54 VTAIL.n18 6.59444
R456 VTAIL.n241 VTAIL.n205 6.59444
R457 VTAIL.n241 VTAIL.n240 6.59444
R458 VTAIL.n149 VTAIL.n113 6.59444
R459 VTAIL.n149 VTAIL.n148 6.59444
R460 VTAIL.n326 VTAIL.n296 5.81868
R461 VTAIL.n334 VTAIL.n333 5.81868
R462 VTAIL.n50 VTAIL.n20 5.81868
R463 VTAIL.n58 VTAIL.n57 5.81868
R464 VTAIL.n245 VTAIL.n244 5.81868
R465 VTAIL.n237 VTAIL.n207 5.81868
R466 VTAIL.n153 VTAIL.n152 5.81868
R467 VTAIL.n145 VTAIL.n115 5.81868
R468 VTAIL.n325 VTAIL.n298 5.04292
R469 VTAIL.n337 VTAIL.n292 5.04292
R470 VTAIL.n49 VTAIL.n22 5.04292
R471 VTAIL.n61 VTAIL.n16 5.04292
R472 VTAIL.n248 VTAIL.n203 5.04292
R473 VTAIL.n236 VTAIL.n209 5.04292
R474 VTAIL.n156 VTAIL.n111 5.04292
R475 VTAIL.n144 VTAIL.n117 5.04292
R476 VTAIL.n322 VTAIL.n321 4.26717
R477 VTAIL.n338 VTAIL.n290 4.26717
R478 VTAIL.n46 VTAIL.n45 4.26717
R479 VTAIL.n62 VTAIL.n14 4.26717
R480 VTAIL.n249 VTAIL.n201 4.26717
R481 VTAIL.n233 VTAIL.n232 4.26717
R482 VTAIL.n157 VTAIL.n109 4.26717
R483 VTAIL.n141 VTAIL.n140 4.26717
R484 VTAIL.n308 VTAIL.n307 3.70982
R485 VTAIL.n32 VTAIL.n31 3.70982
R486 VTAIL.n219 VTAIL.n218 3.70982
R487 VTAIL.n127 VTAIL.n126 3.70982
R488 VTAIL.n318 VTAIL.n300 3.49141
R489 VTAIL.n342 VTAIL.n341 3.49141
R490 VTAIL.n366 VTAIL.n278 3.49141
R491 VTAIL.n42 VTAIL.n24 3.49141
R492 VTAIL.n66 VTAIL.n65 3.49141
R493 VTAIL.n90 VTAIL.n2 3.49141
R494 VTAIL.n276 VTAIL.n188 3.49141
R495 VTAIL.n253 VTAIL.n252 3.49141
R496 VTAIL.n229 VTAIL.n211 3.49141
R497 VTAIL.n184 VTAIL.n96 3.49141
R498 VTAIL.n161 VTAIL.n160 3.49141
R499 VTAIL.n137 VTAIL.n119 3.49141
R500 VTAIL.n185 VTAIL.n95 3.16429
R501 VTAIL.n277 VTAIL.n187 3.16429
R502 VTAIL.n93 VTAIL.n91 3.16429
R503 VTAIL.n317 VTAIL.n302 2.71565
R504 VTAIL.n345 VTAIL.n288 2.71565
R505 VTAIL.n364 VTAIL.n363 2.71565
R506 VTAIL.n41 VTAIL.n26 2.71565
R507 VTAIL.n69 VTAIL.n12 2.71565
R508 VTAIL.n88 VTAIL.n87 2.71565
R509 VTAIL.n274 VTAIL.n273 2.71565
R510 VTAIL.n256 VTAIL.n199 2.71565
R511 VTAIL.n228 VTAIL.n213 2.71565
R512 VTAIL.n182 VTAIL.n181 2.71565
R513 VTAIL.n164 VTAIL.n107 2.71565
R514 VTAIL.n136 VTAIL.n121 2.71565
R515 VTAIL VTAIL.n367 2.31516
R516 VTAIL.n187 VTAIL.n185 2.05222
R517 VTAIL.n91 VTAIL.n1 2.05222
R518 VTAIL.n0 VTAIL.t11 2.00204
R519 VTAIL.n0 VTAIL.t0 2.00204
R520 VTAIL.n92 VTAIL.t6 2.00204
R521 VTAIL.n92 VTAIL.t5 2.00204
R522 VTAIL.n186 VTAIL.t10 2.00204
R523 VTAIL.n186 VTAIL.t9 2.00204
R524 VTAIL.n94 VTAIL.t4 2.00204
R525 VTAIL.n94 VTAIL.t3 2.00204
R526 VTAIL.n314 VTAIL.n313 1.93989
R527 VTAIL.n346 VTAIL.n286 1.93989
R528 VTAIL.n360 VTAIL.n280 1.93989
R529 VTAIL.n38 VTAIL.n37 1.93989
R530 VTAIL.n70 VTAIL.n10 1.93989
R531 VTAIL.n84 VTAIL.n4 1.93989
R532 VTAIL.n270 VTAIL.n190 1.93989
R533 VTAIL.n257 VTAIL.n197 1.93989
R534 VTAIL.n225 VTAIL.n224 1.93989
R535 VTAIL.n178 VTAIL.n98 1.93989
R536 VTAIL.n165 VTAIL.n105 1.93989
R537 VTAIL.n133 VTAIL.n132 1.93989
R538 VTAIL.n310 VTAIL.n304 1.16414
R539 VTAIL.n351 VTAIL.n349 1.16414
R540 VTAIL.n359 VTAIL.n282 1.16414
R541 VTAIL.n34 VTAIL.n28 1.16414
R542 VTAIL.n75 VTAIL.n73 1.16414
R543 VTAIL.n83 VTAIL.n6 1.16414
R544 VTAIL.n269 VTAIL.n192 1.16414
R545 VTAIL.n261 VTAIL.n260 1.16414
R546 VTAIL.n221 VTAIL.n215 1.16414
R547 VTAIL.n177 VTAIL.n100 1.16414
R548 VTAIL.n169 VTAIL.n168 1.16414
R549 VTAIL.n129 VTAIL.n123 1.16414
R550 VTAIL VTAIL.n1 0.849638
R551 VTAIL.n309 VTAIL.n306 0.388379
R552 VTAIL.n350 VTAIL.n284 0.388379
R553 VTAIL.n356 VTAIL.n355 0.388379
R554 VTAIL.n33 VTAIL.n30 0.388379
R555 VTAIL.n74 VTAIL.n8 0.388379
R556 VTAIL.n80 VTAIL.n79 0.388379
R557 VTAIL.n266 VTAIL.n265 0.388379
R558 VTAIL.n196 VTAIL.n194 0.388379
R559 VTAIL.n220 VTAIL.n217 0.388379
R560 VTAIL.n174 VTAIL.n173 0.388379
R561 VTAIL.n104 VTAIL.n102 0.388379
R562 VTAIL.n128 VTAIL.n125 0.388379
R563 VTAIL.n308 VTAIL.n303 0.155672
R564 VTAIL.n315 VTAIL.n303 0.155672
R565 VTAIL.n316 VTAIL.n315 0.155672
R566 VTAIL.n316 VTAIL.n299 0.155672
R567 VTAIL.n323 VTAIL.n299 0.155672
R568 VTAIL.n324 VTAIL.n323 0.155672
R569 VTAIL.n324 VTAIL.n295 0.155672
R570 VTAIL.n331 VTAIL.n295 0.155672
R571 VTAIL.n332 VTAIL.n331 0.155672
R572 VTAIL.n332 VTAIL.n291 0.155672
R573 VTAIL.n339 VTAIL.n291 0.155672
R574 VTAIL.n340 VTAIL.n339 0.155672
R575 VTAIL.n340 VTAIL.n287 0.155672
R576 VTAIL.n347 VTAIL.n287 0.155672
R577 VTAIL.n348 VTAIL.n347 0.155672
R578 VTAIL.n348 VTAIL.n283 0.155672
R579 VTAIL.n357 VTAIL.n283 0.155672
R580 VTAIL.n358 VTAIL.n357 0.155672
R581 VTAIL.n358 VTAIL.n279 0.155672
R582 VTAIL.n365 VTAIL.n279 0.155672
R583 VTAIL.n32 VTAIL.n27 0.155672
R584 VTAIL.n39 VTAIL.n27 0.155672
R585 VTAIL.n40 VTAIL.n39 0.155672
R586 VTAIL.n40 VTAIL.n23 0.155672
R587 VTAIL.n47 VTAIL.n23 0.155672
R588 VTAIL.n48 VTAIL.n47 0.155672
R589 VTAIL.n48 VTAIL.n19 0.155672
R590 VTAIL.n55 VTAIL.n19 0.155672
R591 VTAIL.n56 VTAIL.n55 0.155672
R592 VTAIL.n56 VTAIL.n15 0.155672
R593 VTAIL.n63 VTAIL.n15 0.155672
R594 VTAIL.n64 VTAIL.n63 0.155672
R595 VTAIL.n64 VTAIL.n11 0.155672
R596 VTAIL.n71 VTAIL.n11 0.155672
R597 VTAIL.n72 VTAIL.n71 0.155672
R598 VTAIL.n72 VTAIL.n7 0.155672
R599 VTAIL.n81 VTAIL.n7 0.155672
R600 VTAIL.n82 VTAIL.n81 0.155672
R601 VTAIL.n82 VTAIL.n3 0.155672
R602 VTAIL.n89 VTAIL.n3 0.155672
R603 VTAIL.n275 VTAIL.n189 0.155672
R604 VTAIL.n268 VTAIL.n189 0.155672
R605 VTAIL.n268 VTAIL.n267 0.155672
R606 VTAIL.n267 VTAIL.n193 0.155672
R607 VTAIL.n259 VTAIL.n193 0.155672
R608 VTAIL.n259 VTAIL.n258 0.155672
R609 VTAIL.n258 VTAIL.n198 0.155672
R610 VTAIL.n251 VTAIL.n198 0.155672
R611 VTAIL.n251 VTAIL.n250 0.155672
R612 VTAIL.n250 VTAIL.n202 0.155672
R613 VTAIL.n243 VTAIL.n202 0.155672
R614 VTAIL.n243 VTAIL.n242 0.155672
R615 VTAIL.n242 VTAIL.n206 0.155672
R616 VTAIL.n235 VTAIL.n206 0.155672
R617 VTAIL.n235 VTAIL.n234 0.155672
R618 VTAIL.n234 VTAIL.n210 0.155672
R619 VTAIL.n227 VTAIL.n210 0.155672
R620 VTAIL.n227 VTAIL.n226 0.155672
R621 VTAIL.n226 VTAIL.n214 0.155672
R622 VTAIL.n219 VTAIL.n214 0.155672
R623 VTAIL.n183 VTAIL.n97 0.155672
R624 VTAIL.n176 VTAIL.n97 0.155672
R625 VTAIL.n176 VTAIL.n175 0.155672
R626 VTAIL.n175 VTAIL.n101 0.155672
R627 VTAIL.n167 VTAIL.n101 0.155672
R628 VTAIL.n167 VTAIL.n166 0.155672
R629 VTAIL.n166 VTAIL.n106 0.155672
R630 VTAIL.n159 VTAIL.n106 0.155672
R631 VTAIL.n159 VTAIL.n158 0.155672
R632 VTAIL.n158 VTAIL.n110 0.155672
R633 VTAIL.n151 VTAIL.n110 0.155672
R634 VTAIL.n151 VTAIL.n150 0.155672
R635 VTAIL.n150 VTAIL.n114 0.155672
R636 VTAIL.n143 VTAIL.n114 0.155672
R637 VTAIL.n143 VTAIL.n142 0.155672
R638 VTAIL.n142 VTAIL.n118 0.155672
R639 VTAIL.n135 VTAIL.n118 0.155672
R640 VTAIL.n135 VTAIL.n134 0.155672
R641 VTAIL.n134 VTAIL.n122 0.155672
R642 VTAIL.n127 VTAIL.n122 0.155672
R643 VDD1.n84 VDD1.n0 756.745
R644 VDD1.n173 VDD1.n89 756.745
R645 VDD1.n85 VDD1.n84 585
R646 VDD1.n83 VDD1.n82 585
R647 VDD1.n4 VDD1.n3 585
R648 VDD1.n77 VDD1.n76 585
R649 VDD1.n75 VDD1.n6 585
R650 VDD1.n74 VDD1.n73 585
R651 VDD1.n9 VDD1.n7 585
R652 VDD1.n68 VDD1.n67 585
R653 VDD1.n66 VDD1.n65 585
R654 VDD1.n13 VDD1.n12 585
R655 VDD1.n60 VDD1.n59 585
R656 VDD1.n58 VDD1.n57 585
R657 VDD1.n17 VDD1.n16 585
R658 VDD1.n52 VDD1.n51 585
R659 VDD1.n50 VDD1.n49 585
R660 VDD1.n21 VDD1.n20 585
R661 VDD1.n44 VDD1.n43 585
R662 VDD1.n42 VDD1.n41 585
R663 VDD1.n25 VDD1.n24 585
R664 VDD1.n36 VDD1.n35 585
R665 VDD1.n34 VDD1.n33 585
R666 VDD1.n29 VDD1.n28 585
R667 VDD1.n117 VDD1.n116 585
R668 VDD1.n122 VDD1.n121 585
R669 VDD1.n124 VDD1.n123 585
R670 VDD1.n113 VDD1.n112 585
R671 VDD1.n130 VDD1.n129 585
R672 VDD1.n132 VDD1.n131 585
R673 VDD1.n109 VDD1.n108 585
R674 VDD1.n138 VDD1.n137 585
R675 VDD1.n140 VDD1.n139 585
R676 VDD1.n105 VDD1.n104 585
R677 VDD1.n146 VDD1.n145 585
R678 VDD1.n148 VDD1.n147 585
R679 VDD1.n101 VDD1.n100 585
R680 VDD1.n154 VDD1.n153 585
R681 VDD1.n156 VDD1.n155 585
R682 VDD1.n97 VDD1.n96 585
R683 VDD1.n163 VDD1.n162 585
R684 VDD1.n164 VDD1.n95 585
R685 VDD1.n166 VDD1.n165 585
R686 VDD1.n93 VDD1.n92 585
R687 VDD1.n172 VDD1.n171 585
R688 VDD1.n174 VDD1.n173 585
R689 VDD1.n30 VDD1.t1 327.466
R690 VDD1.n118 VDD1.t2 327.466
R691 VDD1.n84 VDD1.n83 171.744
R692 VDD1.n83 VDD1.n3 171.744
R693 VDD1.n76 VDD1.n3 171.744
R694 VDD1.n76 VDD1.n75 171.744
R695 VDD1.n75 VDD1.n74 171.744
R696 VDD1.n74 VDD1.n7 171.744
R697 VDD1.n67 VDD1.n7 171.744
R698 VDD1.n67 VDD1.n66 171.744
R699 VDD1.n66 VDD1.n12 171.744
R700 VDD1.n59 VDD1.n12 171.744
R701 VDD1.n59 VDD1.n58 171.744
R702 VDD1.n58 VDD1.n16 171.744
R703 VDD1.n51 VDD1.n16 171.744
R704 VDD1.n51 VDD1.n50 171.744
R705 VDD1.n50 VDD1.n20 171.744
R706 VDD1.n43 VDD1.n20 171.744
R707 VDD1.n43 VDD1.n42 171.744
R708 VDD1.n42 VDD1.n24 171.744
R709 VDD1.n35 VDD1.n24 171.744
R710 VDD1.n35 VDD1.n34 171.744
R711 VDD1.n34 VDD1.n28 171.744
R712 VDD1.n122 VDD1.n116 171.744
R713 VDD1.n123 VDD1.n122 171.744
R714 VDD1.n123 VDD1.n112 171.744
R715 VDD1.n130 VDD1.n112 171.744
R716 VDD1.n131 VDD1.n130 171.744
R717 VDD1.n131 VDD1.n108 171.744
R718 VDD1.n138 VDD1.n108 171.744
R719 VDD1.n139 VDD1.n138 171.744
R720 VDD1.n139 VDD1.n104 171.744
R721 VDD1.n146 VDD1.n104 171.744
R722 VDD1.n147 VDD1.n146 171.744
R723 VDD1.n147 VDD1.n100 171.744
R724 VDD1.n154 VDD1.n100 171.744
R725 VDD1.n155 VDD1.n154 171.744
R726 VDD1.n155 VDD1.n96 171.744
R727 VDD1.n163 VDD1.n96 171.744
R728 VDD1.n164 VDD1.n163 171.744
R729 VDD1.n165 VDD1.n164 171.744
R730 VDD1.n165 VDD1.n92 171.744
R731 VDD1.n172 VDD1.n92 171.744
R732 VDD1.n173 VDD1.n172 171.744
R733 VDD1.t1 VDD1.n28 85.8723
R734 VDD1.t2 VDD1.n116 85.8723
R735 VDD1.n179 VDD1.n178 73.6406
R736 VDD1.n181 VDD1.n180 72.905
R737 VDD1 VDD1.n88 54.3982
R738 VDD1.n179 VDD1.n177 54.2847
R739 VDD1.n181 VDD1.n179 50.1625
R740 VDD1.n30 VDD1.n29 16.3895
R741 VDD1.n118 VDD1.n117 16.3895
R742 VDD1.n77 VDD1.n6 13.1884
R743 VDD1.n166 VDD1.n95 13.1884
R744 VDD1.n78 VDD1.n4 12.8005
R745 VDD1.n73 VDD1.n8 12.8005
R746 VDD1.n33 VDD1.n32 12.8005
R747 VDD1.n121 VDD1.n120 12.8005
R748 VDD1.n162 VDD1.n161 12.8005
R749 VDD1.n167 VDD1.n93 12.8005
R750 VDD1.n82 VDD1.n81 12.0247
R751 VDD1.n72 VDD1.n9 12.0247
R752 VDD1.n36 VDD1.n27 12.0247
R753 VDD1.n124 VDD1.n115 12.0247
R754 VDD1.n160 VDD1.n97 12.0247
R755 VDD1.n171 VDD1.n170 12.0247
R756 VDD1.n85 VDD1.n2 11.249
R757 VDD1.n69 VDD1.n68 11.249
R758 VDD1.n37 VDD1.n25 11.249
R759 VDD1.n125 VDD1.n113 11.249
R760 VDD1.n157 VDD1.n156 11.249
R761 VDD1.n174 VDD1.n91 11.249
R762 VDD1.n86 VDD1.n0 10.4732
R763 VDD1.n65 VDD1.n11 10.4732
R764 VDD1.n41 VDD1.n40 10.4732
R765 VDD1.n129 VDD1.n128 10.4732
R766 VDD1.n153 VDD1.n99 10.4732
R767 VDD1.n175 VDD1.n89 10.4732
R768 VDD1.n64 VDD1.n13 9.69747
R769 VDD1.n44 VDD1.n23 9.69747
R770 VDD1.n132 VDD1.n111 9.69747
R771 VDD1.n152 VDD1.n101 9.69747
R772 VDD1.n88 VDD1.n87 9.45567
R773 VDD1.n177 VDD1.n176 9.45567
R774 VDD1.n56 VDD1.n55 9.3005
R775 VDD1.n15 VDD1.n14 9.3005
R776 VDD1.n62 VDD1.n61 9.3005
R777 VDD1.n64 VDD1.n63 9.3005
R778 VDD1.n11 VDD1.n10 9.3005
R779 VDD1.n70 VDD1.n69 9.3005
R780 VDD1.n72 VDD1.n71 9.3005
R781 VDD1.n8 VDD1.n5 9.3005
R782 VDD1.n87 VDD1.n86 9.3005
R783 VDD1.n2 VDD1.n1 9.3005
R784 VDD1.n81 VDD1.n80 9.3005
R785 VDD1.n79 VDD1.n78 9.3005
R786 VDD1.n54 VDD1.n53 9.3005
R787 VDD1.n19 VDD1.n18 9.3005
R788 VDD1.n48 VDD1.n47 9.3005
R789 VDD1.n46 VDD1.n45 9.3005
R790 VDD1.n23 VDD1.n22 9.3005
R791 VDD1.n40 VDD1.n39 9.3005
R792 VDD1.n38 VDD1.n37 9.3005
R793 VDD1.n27 VDD1.n26 9.3005
R794 VDD1.n32 VDD1.n31 9.3005
R795 VDD1.n176 VDD1.n175 9.3005
R796 VDD1.n91 VDD1.n90 9.3005
R797 VDD1.n170 VDD1.n169 9.3005
R798 VDD1.n168 VDD1.n167 9.3005
R799 VDD1.n107 VDD1.n106 9.3005
R800 VDD1.n136 VDD1.n135 9.3005
R801 VDD1.n134 VDD1.n133 9.3005
R802 VDD1.n111 VDD1.n110 9.3005
R803 VDD1.n128 VDD1.n127 9.3005
R804 VDD1.n126 VDD1.n125 9.3005
R805 VDD1.n115 VDD1.n114 9.3005
R806 VDD1.n120 VDD1.n119 9.3005
R807 VDD1.n142 VDD1.n141 9.3005
R808 VDD1.n144 VDD1.n143 9.3005
R809 VDD1.n103 VDD1.n102 9.3005
R810 VDD1.n150 VDD1.n149 9.3005
R811 VDD1.n152 VDD1.n151 9.3005
R812 VDD1.n99 VDD1.n98 9.3005
R813 VDD1.n158 VDD1.n157 9.3005
R814 VDD1.n160 VDD1.n159 9.3005
R815 VDD1.n161 VDD1.n94 9.3005
R816 VDD1.n61 VDD1.n60 8.92171
R817 VDD1.n45 VDD1.n21 8.92171
R818 VDD1.n133 VDD1.n109 8.92171
R819 VDD1.n149 VDD1.n148 8.92171
R820 VDD1.n57 VDD1.n15 8.14595
R821 VDD1.n49 VDD1.n48 8.14595
R822 VDD1.n137 VDD1.n136 8.14595
R823 VDD1.n145 VDD1.n103 8.14595
R824 VDD1.n56 VDD1.n17 7.3702
R825 VDD1.n52 VDD1.n19 7.3702
R826 VDD1.n140 VDD1.n107 7.3702
R827 VDD1.n144 VDD1.n105 7.3702
R828 VDD1.n53 VDD1.n17 6.59444
R829 VDD1.n53 VDD1.n52 6.59444
R830 VDD1.n141 VDD1.n140 6.59444
R831 VDD1.n141 VDD1.n105 6.59444
R832 VDD1.n57 VDD1.n56 5.81868
R833 VDD1.n49 VDD1.n19 5.81868
R834 VDD1.n137 VDD1.n107 5.81868
R835 VDD1.n145 VDD1.n144 5.81868
R836 VDD1.n60 VDD1.n15 5.04292
R837 VDD1.n48 VDD1.n21 5.04292
R838 VDD1.n136 VDD1.n109 5.04292
R839 VDD1.n148 VDD1.n103 5.04292
R840 VDD1.n61 VDD1.n13 4.26717
R841 VDD1.n45 VDD1.n44 4.26717
R842 VDD1.n133 VDD1.n132 4.26717
R843 VDD1.n149 VDD1.n101 4.26717
R844 VDD1.n31 VDD1.n30 3.70982
R845 VDD1.n119 VDD1.n118 3.70982
R846 VDD1.n88 VDD1.n0 3.49141
R847 VDD1.n65 VDD1.n64 3.49141
R848 VDD1.n41 VDD1.n23 3.49141
R849 VDD1.n129 VDD1.n111 3.49141
R850 VDD1.n153 VDD1.n152 3.49141
R851 VDD1.n177 VDD1.n89 3.49141
R852 VDD1.n86 VDD1.n85 2.71565
R853 VDD1.n68 VDD1.n11 2.71565
R854 VDD1.n40 VDD1.n25 2.71565
R855 VDD1.n128 VDD1.n113 2.71565
R856 VDD1.n156 VDD1.n99 2.71565
R857 VDD1.n175 VDD1.n174 2.71565
R858 VDD1.n180 VDD1.t3 2.00204
R859 VDD1.n180 VDD1.t5 2.00204
R860 VDD1.n178 VDD1.t4 2.00204
R861 VDD1.n178 VDD1.t0 2.00204
R862 VDD1.n82 VDD1.n2 1.93989
R863 VDD1.n69 VDD1.n9 1.93989
R864 VDD1.n37 VDD1.n36 1.93989
R865 VDD1.n125 VDD1.n124 1.93989
R866 VDD1.n157 VDD1.n97 1.93989
R867 VDD1.n171 VDD1.n91 1.93989
R868 VDD1.n81 VDD1.n4 1.16414
R869 VDD1.n73 VDD1.n72 1.16414
R870 VDD1.n33 VDD1.n27 1.16414
R871 VDD1.n121 VDD1.n115 1.16414
R872 VDD1.n162 VDD1.n160 1.16414
R873 VDD1.n170 VDD1.n93 1.16414
R874 VDD1 VDD1.n181 0.733259
R875 VDD1.n78 VDD1.n77 0.388379
R876 VDD1.n8 VDD1.n6 0.388379
R877 VDD1.n32 VDD1.n29 0.388379
R878 VDD1.n120 VDD1.n117 0.388379
R879 VDD1.n161 VDD1.n95 0.388379
R880 VDD1.n167 VDD1.n166 0.388379
R881 VDD1.n87 VDD1.n1 0.155672
R882 VDD1.n80 VDD1.n1 0.155672
R883 VDD1.n80 VDD1.n79 0.155672
R884 VDD1.n79 VDD1.n5 0.155672
R885 VDD1.n71 VDD1.n5 0.155672
R886 VDD1.n71 VDD1.n70 0.155672
R887 VDD1.n70 VDD1.n10 0.155672
R888 VDD1.n63 VDD1.n10 0.155672
R889 VDD1.n63 VDD1.n62 0.155672
R890 VDD1.n62 VDD1.n14 0.155672
R891 VDD1.n55 VDD1.n14 0.155672
R892 VDD1.n55 VDD1.n54 0.155672
R893 VDD1.n54 VDD1.n18 0.155672
R894 VDD1.n47 VDD1.n18 0.155672
R895 VDD1.n47 VDD1.n46 0.155672
R896 VDD1.n46 VDD1.n22 0.155672
R897 VDD1.n39 VDD1.n22 0.155672
R898 VDD1.n39 VDD1.n38 0.155672
R899 VDD1.n38 VDD1.n26 0.155672
R900 VDD1.n31 VDD1.n26 0.155672
R901 VDD1.n119 VDD1.n114 0.155672
R902 VDD1.n126 VDD1.n114 0.155672
R903 VDD1.n127 VDD1.n126 0.155672
R904 VDD1.n127 VDD1.n110 0.155672
R905 VDD1.n134 VDD1.n110 0.155672
R906 VDD1.n135 VDD1.n134 0.155672
R907 VDD1.n135 VDD1.n106 0.155672
R908 VDD1.n142 VDD1.n106 0.155672
R909 VDD1.n143 VDD1.n142 0.155672
R910 VDD1.n143 VDD1.n102 0.155672
R911 VDD1.n150 VDD1.n102 0.155672
R912 VDD1.n151 VDD1.n150 0.155672
R913 VDD1.n151 VDD1.n98 0.155672
R914 VDD1.n158 VDD1.n98 0.155672
R915 VDD1.n159 VDD1.n158 0.155672
R916 VDD1.n159 VDD1.n94 0.155672
R917 VDD1.n168 VDD1.n94 0.155672
R918 VDD1.n169 VDD1.n168 0.155672
R919 VDD1.n169 VDD1.n90 0.155672
R920 VDD1.n176 VDD1.n90 0.155672
R921 VN.n34 VN.n33 161.3
R922 VN.n32 VN.n19 161.3
R923 VN.n31 VN.n30 161.3
R924 VN.n29 VN.n20 161.3
R925 VN.n28 VN.n27 161.3
R926 VN.n26 VN.n21 161.3
R927 VN.n25 VN.n24 161.3
R928 VN.n16 VN.n15 161.3
R929 VN.n14 VN.n1 161.3
R930 VN.n13 VN.n12 161.3
R931 VN.n11 VN.n2 161.3
R932 VN.n10 VN.n9 161.3
R933 VN.n8 VN.n3 161.3
R934 VN.n7 VN.n6 161.3
R935 VN.n23 VN.t3 150.376
R936 VN.n5 VN.t0 150.376
R937 VN.n4 VN.t1 117.181
R938 VN.n0 VN.t5 117.181
R939 VN.n22 VN.t2 117.181
R940 VN.n18 VN.t4 117.181
R941 VN.n17 VN.n0 81.8843
R942 VN.n35 VN.n18 81.8843
R943 VN.n9 VN.n2 56.5617
R944 VN.n27 VN.n20 56.5617
R945 VN VN.n35 54.9792
R946 VN.n5 VN.n4 50.1906
R947 VN.n23 VN.n22 50.1906
R948 VN.n7 VN.n4 24.5923
R949 VN.n8 VN.n7 24.5923
R950 VN.n9 VN.n8 24.5923
R951 VN.n13 VN.n2 24.5923
R952 VN.n14 VN.n13 24.5923
R953 VN.n15 VN.n14 24.5923
R954 VN.n27 VN.n26 24.5923
R955 VN.n26 VN.n25 24.5923
R956 VN.n25 VN.n22 24.5923
R957 VN.n33 VN.n32 24.5923
R958 VN.n32 VN.n31 24.5923
R959 VN.n31 VN.n20 24.5923
R960 VN.n15 VN.n0 8.36172
R961 VN.n33 VN.n18 8.36172
R962 VN.n6 VN.n5 3.19893
R963 VN.n24 VN.n23 3.19893
R964 VN.n35 VN.n34 0.354861
R965 VN.n17 VN.n16 0.354861
R966 VN VN.n17 0.267071
R967 VN.n34 VN.n19 0.189894
R968 VN.n30 VN.n19 0.189894
R969 VN.n30 VN.n29 0.189894
R970 VN.n29 VN.n28 0.189894
R971 VN.n28 VN.n21 0.189894
R972 VN.n24 VN.n21 0.189894
R973 VN.n6 VN.n3 0.189894
R974 VN.n10 VN.n3 0.189894
R975 VN.n11 VN.n10 0.189894
R976 VN.n12 VN.n11 0.189894
R977 VN.n12 VN.n1 0.189894
R978 VN.n16 VN.n1 0.189894
R979 VDD2.n175 VDD2.n91 756.745
R980 VDD2.n84 VDD2.n0 756.745
R981 VDD2.n176 VDD2.n175 585
R982 VDD2.n174 VDD2.n173 585
R983 VDD2.n95 VDD2.n94 585
R984 VDD2.n168 VDD2.n167 585
R985 VDD2.n166 VDD2.n97 585
R986 VDD2.n165 VDD2.n164 585
R987 VDD2.n100 VDD2.n98 585
R988 VDD2.n159 VDD2.n158 585
R989 VDD2.n157 VDD2.n156 585
R990 VDD2.n104 VDD2.n103 585
R991 VDD2.n151 VDD2.n150 585
R992 VDD2.n149 VDD2.n148 585
R993 VDD2.n108 VDD2.n107 585
R994 VDD2.n143 VDD2.n142 585
R995 VDD2.n141 VDD2.n140 585
R996 VDD2.n112 VDD2.n111 585
R997 VDD2.n135 VDD2.n134 585
R998 VDD2.n133 VDD2.n132 585
R999 VDD2.n116 VDD2.n115 585
R1000 VDD2.n127 VDD2.n126 585
R1001 VDD2.n125 VDD2.n124 585
R1002 VDD2.n120 VDD2.n119 585
R1003 VDD2.n28 VDD2.n27 585
R1004 VDD2.n33 VDD2.n32 585
R1005 VDD2.n35 VDD2.n34 585
R1006 VDD2.n24 VDD2.n23 585
R1007 VDD2.n41 VDD2.n40 585
R1008 VDD2.n43 VDD2.n42 585
R1009 VDD2.n20 VDD2.n19 585
R1010 VDD2.n49 VDD2.n48 585
R1011 VDD2.n51 VDD2.n50 585
R1012 VDD2.n16 VDD2.n15 585
R1013 VDD2.n57 VDD2.n56 585
R1014 VDD2.n59 VDD2.n58 585
R1015 VDD2.n12 VDD2.n11 585
R1016 VDD2.n65 VDD2.n64 585
R1017 VDD2.n67 VDD2.n66 585
R1018 VDD2.n8 VDD2.n7 585
R1019 VDD2.n74 VDD2.n73 585
R1020 VDD2.n75 VDD2.n6 585
R1021 VDD2.n77 VDD2.n76 585
R1022 VDD2.n4 VDD2.n3 585
R1023 VDD2.n83 VDD2.n82 585
R1024 VDD2.n85 VDD2.n84 585
R1025 VDD2.n121 VDD2.t1 327.466
R1026 VDD2.n29 VDD2.t5 327.466
R1027 VDD2.n175 VDD2.n174 171.744
R1028 VDD2.n174 VDD2.n94 171.744
R1029 VDD2.n167 VDD2.n94 171.744
R1030 VDD2.n167 VDD2.n166 171.744
R1031 VDD2.n166 VDD2.n165 171.744
R1032 VDD2.n165 VDD2.n98 171.744
R1033 VDD2.n158 VDD2.n98 171.744
R1034 VDD2.n158 VDD2.n157 171.744
R1035 VDD2.n157 VDD2.n103 171.744
R1036 VDD2.n150 VDD2.n103 171.744
R1037 VDD2.n150 VDD2.n149 171.744
R1038 VDD2.n149 VDD2.n107 171.744
R1039 VDD2.n142 VDD2.n107 171.744
R1040 VDD2.n142 VDD2.n141 171.744
R1041 VDD2.n141 VDD2.n111 171.744
R1042 VDD2.n134 VDD2.n111 171.744
R1043 VDD2.n134 VDD2.n133 171.744
R1044 VDD2.n133 VDD2.n115 171.744
R1045 VDD2.n126 VDD2.n115 171.744
R1046 VDD2.n126 VDD2.n125 171.744
R1047 VDD2.n125 VDD2.n119 171.744
R1048 VDD2.n33 VDD2.n27 171.744
R1049 VDD2.n34 VDD2.n33 171.744
R1050 VDD2.n34 VDD2.n23 171.744
R1051 VDD2.n41 VDD2.n23 171.744
R1052 VDD2.n42 VDD2.n41 171.744
R1053 VDD2.n42 VDD2.n19 171.744
R1054 VDD2.n49 VDD2.n19 171.744
R1055 VDD2.n50 VDD2.n49 171.744
R1056 VDD2.n50 VDD2.n15 171.744
R1057 VDD2.n57 VDD2.n15 171.744
R1058 VDD2.n58 VDD2.n57 171.744
R1059 VDD2.n58 VDD2.n11 171.744
R1060 VDD2.n65 VDD2.n11 171.744
R1061 VDD2.n66 VDD2.n65 171.744
R1062 VDD2.n66 VDD2.n7 171.744
R1063 VDD2.n74 VDD2.n7 171.744
R1064 VDD2.n75 VDD2.n74 171.744
R1065 VDD2.n76 VDD2.n75 171.744
R1066 VDD2.n76 VDD2.n3 171.744
R1067 VDD2.n83 VDD2.n3 171.744
R1068 VDD2.n84 VDD2.n83 171.744
R1069 VDD2.t1 VDD2.n119 85.8723
R1070 VDD2.t5 VDD2.n27 85.8723
R1071 VDD2.n90 VDD2.n89 73.6406
R1072 VDD2 VDD2.n181 73.6377
R1073 VDD2.n90 VDD2.n88 54.2847
R1074 VDD2.n180 VDD2.n179 51.9672
R1075 VDD2.n180 VDD2.n90 47.9976
R1076 VDD2.n121 VDD2.n120 16.3895
R1077 VDD2.n29 VDD2.n28 16.3895
R1078 VDD2.n168 VDD2.n97 13.1884
R1079 VDD2.n77 VDD2.n6 13.1884
R1080 VDD2.n169 VDD2.n95 12.8005
R1081 VDD2.n164 VDD2.n99 12.8005
R1082 VDD2.n124 VDD2.n123 12.8005
R1083 VDD2.n32 VDD2.n31 12.8005
R1084 VDD2.n73 VDD2.n72 12.8005
R1085 VDD2.n78 VDD2.n4 12.8005
R1086 VDD2.n173 VDD2.n172 12.0247
R1087 VDD2.n163 VDD2.n100 12.0247
R1088 VDD2.n127 VDD2.n118 12.0247
R1089 VDD2.n35 VDD2.n26 12.0247
R1090 VDD2.n71 VDD2.n8 12.0247
R1091 VDD2.n82 VDD2.n81 12.0247
R1092 VDD2.n176 VDD2.n93 11.249
R1093 VDD2.n160 VDD2.n159 11.249
R1094 VDD2.n128 VDD2.n116 11.249
R1095 VDD2.n36 VDD2.n24 11.249
R1096 VDD2.n68 VDD2.n67 11.249
R1097 VDD2.n85 VDD2.n2 11.249
R1098 VDD2.n177 VDD2.n91 10.4732
R1099 VDD2.n156 VDD2.n102 10.4732
R1100 VDD2.n132 VDD2.n131 10.4732
R1101 VDD2.n40 VDD2.n39 10.4732
R1102 VDD2.n64 VDD2.n10 10.4732
R1103 VDD2.n86 VDD2.n0 10.4732
R1104 VDD2.n155 VDD2.n104 9.69747
R1105 VDD2.n135 VDD2.n114 9.69747
R1106 VDD2.n43 VDD2.n22 9.69747
R1107 VDD2.n63 VDD2.n12 9.69747
R1108 VDD2.n179 VDD2.n178 9.45567
R1109 VDD2.n88 VDD2.n87 9.45567
R1110 VDD2.n147 VDD2.n146 9.3005
R1111 VDD2.n106 VDD2.n105 9.3005
R1112 VDD2.n153 VDD2.n152 9.3005
R1113 VDD2.n155 VDD2.n154 9.3005
R1114 VDD2.n102 VDD2.n101 9.3005
R1115 VDD2.n161 VDD2.n160 9.3005
R1116 VDD2.n163 VDD2.n162 9.3005
R1117 VDD2.n99 VDD2.n96 9.3005
R1118 VDD2.n178 VDD2.n177 9.3005
R1119 VDD2.n93 VDD2.n92 9.3005
R1120 VDD2.n172 VDD2.n171 9.3005
R1121 VDD2.n170 VDD2.n169 9.3005
R1122 VDD2.n145 VDD2.n144 9.3005
R1123 VDD2.n110 VDD2.n109 9.3005
R1124 VDD2.n139 VDD2.n138 9.3005
R1125 VDD2.n137 VDD2.n136 9.3005
R1126 VDD2.n114 VDD2.n113 9.3005
R1127 VDD2.n131 VDD2.n130 9.3005
R1128 VDD2.n129 VDD2.n128 9.3005
R1129 VDD2.n118 VDD2.n117 9.3005
R1130 VDD2.n123 VDD2.n122 9.3005
R1131 VDD2.n87 VDD2.n86 9.3005
R1132 VDD2.n2 VDD2.n1 9.3005
R1133 VDD2.n81 VDD2.n80 9.3005
R1134 VDD2.n79 VDD2.n78 9.3005
R1135 VDD2.n18 VDD2.n17 9.3005
R1136 VDD2.n47 VDD2.n46 9.3005
R1137 VDD2.n45 VDD2.n44 9.3005
R1138 VDD2.n22 VDD2.n21 9.3005
R1139 VDD2.n39 VDD2.n38 9.3005
R1140 VDD2.n37 VDD2.n36 9.3005
R1141 VDD2.n26 VDD2.n25 9.3005
R1142 VDD2.n31 VDD2.n30 9.3005
R1143 VDD2.n53 VDD2.n52 9.3005
R1144 VDD2.n55 VDD2.n54 9.3005
R1145 VDD2.n14 VDD2.n13 9.3005
R1146 VDD2.n61 VDD2.n60 9.3005
R1147 VDD2.n63 VDD2.n62 9.3005
R1148 VDD2.n10 VDD2.n9 9.3005
R1149 VDD2.n69 VDD2.n68 9.3005
R1150 VDD2.n71 VDD2.n70 9.3005
R1151 VDD2.n72 VDD2.n5 9.3005
R1152 VDD2.n152 VDD2.n151 8.92171
R1153 VDD2.n136 VDD2.n112 8.92171
R1154 VDD2.n44 VDD2.n20 8.92171
R1155 VDD2.n60 VDD2.n59 8.92171
R1156 VDD2.n148 VDD2.n106 8.14595
R1157 VDD2.n140 VDD2.n139 8.14595
R1158 VDD2.n48 VDD2.n47 8.14595
R1159 VDD2.n56 VDD2.n14 8.14595
R1160 VDD2.n147 VDD2.n108 7.3702
R1161 VDD2.n143 VDD2.n110 7.3702
R1162 VDD2.n51 VDD2.n18 7.3702
R1163 VDD2.n55 VDD2.n16 7.3702
R1164 VDD2.n144 VDD2.n108 6.59444
R1165 VDD2.n144 VDD2.n143 6.59444
R1166 VDD2.n52 VDD2.n51 6.59444
R1167 VDD2.n52 VDD2.n16 6.59444
R1168 VDD2.n148 VDD2.n147 5.81868
R1169 VDD2.n140 VDD2.n110 5.81868
R1170 VDD2.n48 VDD2.n18 5.81868
R1171 VDD2.n56 VDD2.n55 5.81868
R1172 VDD2.n151 VDD2.n106 5.04292
R1173 VDD2.n139 VDD2.n112 5.04292
R1174 VDD2.n47 VDD2.n20 5.04292
R1175 VDD2.n59 VDD2.n14 5.04292
R1176 VDD2.n152 VDD2.n104 4.26717
R1177 VDD2.n136 VDD2.n135 4.26717
R1178 VDD2.n44 VDD2.n43 4.26717
R1179 VDD2.n60 VDD2.n12 4.26717
R1180 VDD2.n122 VDD2.n121 3.70982
R1181 VDD2.n30 VDD2.n29 3.70982
R1182 VDD2.n179 VDD2.n91 3.49141
R1183 VDD2.n156 VDD2.n155 3.49141
R1184 VDD2.n132 VDD2.n114 3.49141
R1185 VDD2.n40 VDD2.n22 3.49141
R1186 VDD2.n64 VDD2.n63 3.49141
R1187 VDD2.n88 VDD2.n0 3.49141
R1188 VDD2.n177 VDD2.n176 2.71565
R1189 VDD2.n159 VDD2.n102 2.71565
R1190 VDD2.n131 VDD2.n116 2.71565
R1191 VDD2.n39 VDD2.n24 2.71565
R1192 VDD2.n67 VDD2.n10 2.71565
R1193 VDD2.n86 VDD2.n85 2.71565
R1194 VDD2 VDD2.n180 2.43153
R1195 VDD2.n181 VDD2.t3 2.00204
R1196 VDD2.n181 VDD2.t2 2.00204
R1197 VDD2.n89 VDD2.t4 2.00204
R1198 VDD2.n89 VDD2.t0 2.00204
R1199 VDD2.n173 VDD2.n93 1.93989
R1200 VDD2.n160 VDD2.n100 1.93989
R1201 VDD2.n128 VDD2.n127 1.93989
R1202 VDD2.n36 VDD2.n35 1.93989
R1203 VDD2.n68 VDD2.n8 1.93989
R1204 VDD2.n82 VDD2.n2 1.93989
R1205 VDD2.n172 VDD2.n95 1.16414
R1206 VDD2.n164 VDD2.n163 1.16414
R1207 VDD2.n124 VDD2.n118 1.16414
R1208 VDD2.n32 VDD2.n26 1.16414
R1209 VDD2.n73 VDD2.n71 1.16414
R1210 VDD2.n81 VDD2.n4 1.16414
R1211 VDD2.n169 VDD2.n168 0.388379
R1212 VDD2.n99 VDD2.n97 0.388379
R1213 VDD2.n123 VDD2.n120 0.388379
R1214 VDD2.n31 VDD2.n28 0.388379
R1215 VDD2.n72 VDD2.n6 0.388379
R1216 VDD2.n78 VDD2.n77 0.388379
R1217 VDD2.n178 VDD2.n92 0.155672
R1218 VDD2.n171 VDD2.n92 0.155672
R1219 VDD2.n171 VDD2.n170 0.155672
R1220 VDD2.n170 VDD2.n96 0.155672
R1221 VDD2.n162 VDD2.n96 0.155672
R1222 VDD2.n162 VDD2.n161 0.155672
R1223 VDD2.n161 VDD2.n101 0.155672
R1224 VDD2.n154 VDD2.n101 0.155672
R1225 VDD2.n154 VDD2.n153 0.155672
R1226 VDD2.n153 VDD2.n105 0.155672
R1227 VDD2.n146 VDD2.n105 0.155672
R1228 VDD2.n146 VDD2.n145 0.155672
R1229 VDD2.n145 VDD2.n109 0.155672
R1230 VDD2.n138 VDD2.n109 0.155672
R1231 VDD2.n138 VDD2.n137 0.155672
R1232 VDD2.n137 VDD2.n113 0.155672
R1233 VDD2.n130 VDD2.n113 0.155672
R1234 VDD2.n130 VDD2.n129 0.155672
R1235 VDD2.n129 VDD2.n117 0.155672
R1236 VDD2.n122 VDD2.n117 0.155672
R1237 VDD2.n30 VDD2.n25 0.155672
R1238 VDD2.n37 VDD2.n25 0.155672
R1239 VDD2.n38 VDD2.n37 0.155672
R1240 VDD2.n38 VDD2.n21 0.155672
R1241 VDD2.n45 VDD2.n21 0.155672
R1242 VDD2.n46 VDD2.n45 0.155672
R1243 VDD2.n46 VDD2.n17 0.155672
R1244 VDD2.n53 VDD2.n17 0.155672
R1245 VDD2.n54 VDD2.n53 0.155672
R1246 VDD2.n54 VDD2.n13 0.155672
R1247 VDD2.n61 VDD2.n13 0.155672
R1248 VDD2.n62 VDD2.n61 0.155672
R1249 VDD2.n62 VDD2.n9 0.155672
R1250 VDD2.n69 VDD2.n9 0.155672
R1251 VDD2.n70 VDD2.n69 0.155672
R1252 VDD2.n70 VDD2.n5 0.155672
R1253 VDD2.n79 VDD2.n5 0.155672
R1254 VDD2.n80 VDD2.n79 0.155672
R1255 VDD2.n80 VDD2.n1 0.155672
R1256 VDD2.n87 VDD2.n1 0.155672
R1257 B.n485 B.n484 585
R1258 B.n483 B.n144 585
R1259 B.n482 B.n481 585
R1260 B.n480 B.n145 585
R1261 B.n479 B.n478 585
R1262 B.n477 B.n146 585
R1263 B.n476 B.n475 585
R1264 B.n474 B.n147 585
R1265 B.n473 B.n472 585
R1266 B.n471 B.n148 585
R1267 B.n470 B.n469 585
R1268 B.n468 B.n149 585
R1269 B.n467 B.n466 585
R1270 B.n465 B.n150 585
R1271 B.n464 B.n463 585
R1272 B.n462 B.n151 585
R1273 B.n461 B.n460 585
R1274 B.n459 B.n152 585
R1275 B.n458 B.n457 585
R1276 B.n456 B.n153 585
R1277 B.n455 B.n454 585
R1278 B.n453 B.n154 585
R1279 B.n452 B.n451 585
R1280 B.n450 B.n155 585
R1281 B.n449 B.n448 585
R1282 B.n447 B.n156 585
R1283 B.n446 B.n445 585
R1284 B.n444 B.n157 585
R1285 B.n443 B.n442 585
R1286 B.n441 B.n158 585
R1287 B.n440 B.n439 585
R1288 B.n438 B.n159 585
R1289 B.n437 B.n436 585
R1290 B.n435 B.n160 585
R1291 B.n434 B.n433 585
R1292 B.n432 B.n161 585
R1293 B.n431 B.n430 585
R1294 B.n429 B.n162 585
R1295 B.n428 B.n427 585
R1296 B.n426 B.n163 585
R1297 B.n425 B.n424 585
R1298 B.n423 B.n164 585
R1299 B.n422 B.n421 585
R1300 B.n420 B.n165 585
R1301 B.n419 B.n418 585
R1302 B.n417 B.n166 585
R1303 B.n416 B.n415 585
R1304 B.n414 B.n167 585
R1305 B.n413 B.n412 585
R1306 B.n411 B.n168 585
R1307 B.n410 B.n409 585
R1308 B.n408 B.n169 585
R1309 B.n407 B.n406 585
R1310 B.n405 B.n170 585
R1311 B.n403 B.n402 585
R1312 B.n401 B.n173 585
R1313 B.n400 B.n399 585
R1314 B.n398 B.n174 585
R1315 B.n397 B.n396 585
R1316 B.n395 B.n175 585
R1317 B.n394 B.n393 585
R1318 B.n392 B.n176 585
R1319 B.n391 B.n390 585
R1320 B.n389 B.n177 585
R1321 B.n388 B.n387 585
R1322 B.n383 B.n178 585
R1323 B.n382 B.n381 585
R1324 B.n380 B.n179 585
R1325 B.n379 B.n378 585
R1326 B.n377 B.n180 585
R1327 B.n376 B.n375 585
R1328 B.n374 B.n181 585
R1329 B.n373 B.n372 585
R1330 B.n371 B.n182 585
R1331 B.n370 B.n369 585
R1332 B.n368 B.n183 585
R1333 B.n367 B.n366 585
R1334 B.n365 B.n184 585
R1335 B.n364 B.n363 585
R1336 B.n362 B.n185 585
R1337 B.n361 B.n360 585
R1338 B.n359 B.n186 585
R1339 B.n358 B.n357 585
R1340 B.n356 B.n187 585
R1341 B.n355 B.n354 585
R1342 B.n353 B.n188 585
R1343 B.n352 B.n351 585
R1344 B.n350 B.n189 585
R1345 B.n349 B.n348 585
R1346 B.n347 B.n190 585
R1347 B.n346 B.n345 585
R1348 B.n344 B.n191 585
R1349 B.n343 B.n342 585
R1350 B.n341 B.n192 585
R1351 B.n340 B.n339 585
R1352 B.n338 B.n193 585
R1353 B.n337 B.n336 585
R1354 B.n335 B.n194 585
R1355 B.n334 B.n333 585
R1356 B.n332 B.n195 585
R1357 B.n331 B.n330 585
R1358 B.n329 B.n196 585
R1359 B.n328 B.n327 585
R1360 B.n326 B.n197 585
R1361 B.n325 B.n324 585
R1362 B.n323 B.n198 585
R1363 B.n322 B.n321 585
R1364 B.n320 B.n199 585
R1365 B.n319 B.n318 585
R1366 B.n317 B.n200 585
R1367 B.n316 B.n315 585
R1368 B.n314 B.n201 585
R1369 B.n313 B.n312 585
R1370 B.n311 B.n202 585
R1371 B.n310 B.n309 585
R1372 B.n308 B.n203 585
R1373 B.n307 B.n306 585
R1374 B.n305 B.n204 585
R1375 B.n486 B.n143 585
R1376 B.n488 B.n487 585
R1377 B.n489 B.n142 585
R1378 B.n491 B.n490 585
R1379 B.n492 B.n141 585
R1380 B.n494 B.n493 585
R1381 B.n495 B.n140 585
R1382 B.n497 B.n496 585
R1383 B.n498 B.n139 585
R1384 B.n500 B.n499 585
R1385 B.n501 B.n138 585
R1386 B.n503 B.n502 585
R1387 B.n504 B.n137 585
R1388 B.n506 B.n505 585
R1389 B.n507 B.n136 585
R1390 B.n509 B.n508 585
R1391 B.n510 B.n135 585
R1392 B.n512 B.n511 585
R1393 B.n513 B.n134 585
R1394 B.n515 B.n514 585
R1395 B.n516 B.n133 585
R1396 B.n518 B.n517 585
R1397 B.n519 B.n132 585
R1398 B.n521 B.n520 585
R1399 B.n522 B.n131 585
R1400 B.n524 B.n523 585
R1401 B.n525 B.n130 585
R1402 B.n527 B.n526 585
R1403 B.n528 B.n129 585
R1404 B.n530 B.n529 585
R1405 B.n531 B.n128 585
R1406 B.n533 B.n532 585
R1407 B.n534 B.n127 585
R1408 B.n536 B.n535 585
R1409 B.n537 B.n126 585
R1410 B.n539 B.n538 585
R1411 B.n540 B.n125 585
R1412 B.n542 B.n541 585
R1413 B.n543 B.n124 585
R1414 B.n545 B.n544 585
R1415 B.n546 B.n123 585
R1416 B.n548 B.n547 585
R1417 B.n549 B.n122 585
R1418 B.n551 B.n550 585
R1419 B.n552 B.n121 585
R1420 B.n554 B.n553 585
R1421 B.n555 B.n120 585
R1422 B.n557 B.n556 585
R1423 B.n558 B.n119 585
R1424 B.n560 B.n559 585
R1425 B.n561 B.n118 585
R1426 B.n563 B.n562 585
R1427 B.n564 B.n117 585
R1428 B.n566 B.n565 585
R1429 B.n567 B.n116 585
R1430 B.n569 B.n568 585
R1431 B.n570 B.n115 585
R1432 B.n572 B.n571 585
R1433 B.n573 B.n114 585
R1434 B.n575 B.n574 585
R1435 B.n576 B.n113 585
R1436 B.n578 B.n577 585
R1437 B.n579 B.n112 585
R1438 B.n581 B.n580 585
R1439 B.n582 B.n111 585
R1440 B.n584 B.n583 585
R1441 B.n585 B.n110 585
R1442 B.n587 B.n586 585
R1443 B.n588 B.n109 585
R1444 B.n590 B.n589 585
R1445 B.n591 B.n108 585
R1446 B.n593 B.n592 585
R1447 B.n594 B.n107 585
R1448 B.n596 B.n595 585
R1449 B.n597 B.n106 585
R1450 B.n599 B.n598 585
R1451 B.n600 B.n105 585
R1452 B.n602 B.n601 585
R1453 B.n603 B.n104 585
R1454 B.n605 B.n604 585
R1455 B.n606 B.n103 585
R1456 B.n608 B.n607 585
R1457 B.n609 B.n102 585
R1458 B.n611 B.n610 585
R1459 B.n612 B.n101 585
R1460 B.n614 B.n613 585
R1461 B.n615 B.n100 585
R1462 B.n617 B.n616 585
R1463 B.n618 B.n99 585
R1464 B.n620 B.n619 585
R1465 B.n621 B.n98 585
R1466 B.n623 B.n622 585
R1467 B.n624 B.n97 585
R1468 B.n626 B.n625 585
R1469 B.n627 B.n96 585
R1470 B.n629 B.n628 585
R1471 B.n630 B.n95 585
R1472 B.n632 B.n631 585
R1473 B.n633 B.n94 585
R1474 B.n635 B.n634 585
R1475 B.n636 B.n93 585
R1476 B.n638 B.n637 585
R1477 B.n639 B.n92 585
R1478 B.n641 B.n640 585
R1479 B.n819 B.n818 585
R1480 B.n817 B.n28 585
R1481 B.n816 B.n815 585
R1482 B.n814 B.n29 585
R1483 B.n813 B.n812 585
R1484 B.n811 B.n30 585
R1485 B.n810 B.n809 585
R1486 B.n808 B.n31 585
R1487 B.n807 B.n806 585
R1488 B.n805 B.n32 585
R1489 B.n804 B.n803 585
R1490 B.n802 B.n33 585
R1491 B.n801 B.n800 585
R1492 B.n799 B.n34 585
R1493 B.n798 B.n797 585
R1494 B.n796 B.n35 585
R1495 B.n795 B.n794 585
R1496 B.n793 B.n36 585
R1497 B.n792 B.n791 585
R1498 B.n790 B.n37 585
R1499 B.n789 B.n788 585
R1500 B.n787 B.n38 585
R1501 B.n786 B.n785 585
R1502 B.n784 B.n39 585
R1503 B.n783 B.n782 585
R1504 B.n781 B.n40 585
R1505 B.n780 B.n779 585
R1506 B.n778 B.n41 585
R1507 B.n777 B.n776 585
R1508 B.n775 B.n42 585
R1509 B.n774 B.n773 585
R1510 B.n772 B.n43 585
R1511 B.n771 B.n770 585
R1512 B.n769 B.n44 585
R1513 B.n768 B.n767 585
R1514 B.n766 B.n45 585
R1515 B.n765 B.n764 585
R1516 B.n763 B.n46 585
R1517 B.n762 B.n761 585
R1518 B.n760 B.n47 585
R1519 B.n759 B.n758 585
R1520 B.n757 B.n48 585
R1521 B.n756 B.n755 585
R1522 B.n754 B.n49 585
R1523 B.n753 B.n752 585
R1524 B.n751 B.n50 585
R1525 B.n750 B.n749 585
R1526 B.n748 B.n51 585
R1527 B.n747 B.n746 585
R1528 B.n745 B.n52 585
R1529 B.n744 B.n743 585
R1530 B.n742 B.n53 585
R1531 B.n741 B.n740 585
R1532 B.n739 B.n54 585
R1533 B.n738 B.n737 585
R1534 B.n736 B.n55 585
R1535 B.n735 B.n734 585
R1536 B.n733 B.n59 585
R1537 B.n732 B.n731 585
R1538 B.n730 B.n60 585
R1539 B.n729 B.n728 585
R1540 B.n727 B.n61 585
R1541 B.n726 B.n725 585
R1542 B.n724 B.n62 585
R1543 B.n722 B.n721 585
R1544 B.n720 B.n65 585
R1545 B.n719 B.n718 585
R1546 B.n717 B.n66 585
R1547 B.n716 B.n715 585
R1548 B.n714 B.n67 585
R1549 B.n713 B.n712 585
R1550 B.n711 B.n68 585
R1551 B.n710 B.n709 585
R1552 B.n708 B.n69 585
R1553 B.n707 B.n706 585
R1554 B.n705 B.n70 585
R1555 B.n704 B.n703 585
R1556 B.n702 B.n71 585
R1557 B.n701 B.n700 585
R1558 B.n699 B.n72 585
R1559 B.n698 B.n697 585
R1560 B.n696 B.n73 585
R1561 B.n695 B.n694 585
R1562 B.n693 B.n74 585
R1563 B.n692 B.n691 585
R1564 B.n690 B.n75 585
R1565 B.n689 B.n688 585
R1566 B.n687 B.n76 585
R1567 B.n686 B.n685 585
R1568 B.n684 B.n77 585
R1569 B.n683 B.n682 585
R1570 B.n681 B.n78 585
R1571 B.n680 B.n679 585
R1572 B.n678 B.n79 585
R1573 B.n677 B.n676 585
R1574 B.n675 B.n80 585
R1575 B.n674 B.n673 585
R1576 B.n672 B.n81 585
R1577 B.n671 B.n670 585
R1578 B.n669 B.n82 585
R1579 B.n668 B.n667 585
R1580 B.n666 B.n83 585
R1581 B.n665 B.n664 585
R1582 B.n663 B.n84 585
R1583 B.n662 B.n661 585
R1584 B.n660 B.n85 585
R1585 B.n659 B.n658 585
R1586 B.n657 B.n86 585
R1587 B.n656 B.n655 585
R1588 B.n654 B.n87 585
R1589 B.n653 B.n652 585
R1590 B.n651 B.n88 585
R1591 B.n650 B.n649 585
R1592 B.n648 B.n89 585
R1593 B.n647 B.n646 585
R1594 B.n645 B.n90 585
R1595 B.n644 B.n643 585
R1596 B.n642 B.n91 585
R1597 B.n820 B.n27 585
R1598 B.n822 B.n821 585
R1599 B.n823 B.n26 585
R1600 B.n825 B.n824 585
R1601 B.n826 B.n25 585
R1602 B.n828 B.n827 585
R1603 B.n829 B.n24 585
R1604 B.n831 B.n830 585
R1605 B.n832 B.n23 585
R1606 B.n834 B.n833 585
R1607 B.n835 B.n22 585
R1608 B.n837 B.n836 585
R1609 B.n838 B.n21 585
R1610 B.n840 B.n839 585
R1611 B.n841 B.n20 585
R1612 B.n843 B.n842 585
R1613 B.n844 B.n19 585
R1614 B.n846 B.n845 585
R1615 B.n847 B.n18 585
R1616 B.n849 B.n848 585
R1617 B.n850 B.n17 585
R1618 B.n852 B.n851 585
R1619 B.n853 B.n16 585
R1620 B.n855 B.n854 585
R1621 B.n856 B.n15 585
R1622 B.n858 B.n857 585
R1623 B.n859 B.n14 585
R1624 B.n861 B.n860 585
R1625 B.n862 B.n13 585
R1626 B.n864 B.n863 585
R1627 B.n865 B.n12 585
R1628 B.n867 B.n866 585
R1629 B.n868 B.n11 585
R1630 B.n870 B.n869 585
R1631 B.n871 B.n10 585
R1632 B.n873 B.n872 585
R1633 B.n874 B.n9 585
R1634 B.n876 B.n875 585
R1635 B.n877 B.n8 585
R1636 B.n879 B.n878 585
R1637 B.n880 B.n7 585
R1638 B.n882 B.n881 585
R1639 B.n883 B.n6 585
R1640 B.n885 B.n884 585
R1641 B.n886 B.n5 585
R1642 B.n888 B.n887 585
R1643 B.n889 B.n4 585
R1644 B.n891 B.n890 585
R1645 B.n892 B.n3 585
R1646 B.n894 B.n893 585
R1647 B.n895 B.n0 585
R1648 B.n2 B.n1 585
R1649 B.n230 B.n229 585
R1650 B.n232 B.n231 585
R1651 B.n233 B.n228 585
R1652 B.n235 B.n234 585
R1653 B.n236 B.n227 585
R1654 B.n238 B.n237 585
R1655 B.n239 B.n226 585
R1656 B.n241 B.n240 585
R1657 B.n242 B.n225 585
R1658 B.n244 B.n243 585
R1659 B.n245 B.n224 585
R1660 B.n247 B.n246 585
R1661 B.n248 B.n223 585
R1662 B.n250 B.n249 585
R1663 B.n251 B.n222 585
R1664 B.n253 B.n252 585
R1665 B.n254 B.n221 585
R1666 B.n256 B.n255 585
R1667 B.n257 B.n220 585
R1668 B.n259 B.n258 585
R1669 B.n260 B.n219 585
R1670 B.n262 B.n261 585
R1671 B.n263 B.n218 585
R1672 B.n265 B.n264 585
R1673 B.n266 B.n217 585
R1674 B.n268 B.n267 585
R1675 B.n269 B.n216 585
R1676 B.n271 B.n270 585
R1677 B.n272 B.n215 585
R1678 B.n274 B.n273 585
R1679 B.n275 B.n214 585
R1680 B.n277 B.n276 585
R1681 B.n278 B.n213 585
R1682 B.n280 B.n279 585
R1683 B.n281 B.n212 585
R1684 B.n283 B.n282 585
R1685 B.n284 B.n211 585
R1686 B.n286 B.n285 585
R1687 B.n287 B.n210 585
R1688 B.n289 B.n288 585
R1689 B.n290 B.n209 585
R1690 B.n292 B.n291 585
R1691 B.n293 B.n208 585
R1692 B.n295 B.n294 585
R1693 B.n296 B.n207 585
R1694 B.n298 B.n297 585
R1695 B.n299 B.n206 585
R1696 B.n301 B.n300 585
R1697 B.n302 B.n205 585
R1698 B.n304 B.n303 585
R1699 B.n171 B.t10 523.295
R1700 B.n63 B.t2 523.295
R1701 B.n384 B.t7 523.295
R1702 B.n56 B.t5 523.295
R1703 B.n172 B.t11 452.12
R1704 B.n64 B.t1 452.12
R1705 B.n385 B.t8 452.12
R1706 B.n57 B.t4 452.12
R1707 B.n303 B.n204 444.452
R1708 B.n486 B.n485 444.452
R1709 B.n642 B.n641 444.452
R1710 B.n818 B.n27 444.452
R1711 B.n384 B.t6 326.125
R1712 B.n171 B.t9 326.125
R1713 B.n63 B.t0 326.125
R1714 B.n56 B.t3 326.125
R1715 B.n897 B.n896 256.663
R1716 B.n896 B.n895 235.042
R1717 B.n896 B.n2 235.042
R1718 B.n307 B.n204 163.367
R1719 B.n308 B.n307 163.367
R1720 B.n309 B.n308 163.367
R1721 B.n309 B.n202 163.367
R1722 B.n313 B.n202 163.367
R1723 B.n314 B.n313 163.367
R1724 B.n315 B.n314 163.367
R1725 B.n315 B.n200 163.367
R1726 B.n319 B.n200 163.367
R1727 B.n320 B.n319 163.367
R1728 B.n321 B.n320 163.367
R1729 B.n321 B.n198 163.367
R1730 B.n325 B.n198 163.367
R1731 B.n326 B.n325 163.367
R1732 B.n327 B.n326 163.367
R1733 B.n327 B.n196 163.367
R1734 B.n331 B.n196 163.367
R1735 B.n332 B.n331 163.367
R1736 B.n333 B.n332 163.367
R1737 B.n333 B.n194 163.367
R1738 B.n337 B.n194 163.367
R1739 B.n338 B.n337 163.367
R1740 B.n339 B.n338 163.367
R1741 B.n339 B.n192 163.367
R1742 B.n343 B.n192 163.367
R1743 B.n344 B.n343 163.367
R1744 B.n345 B.n344 163.367
R1745 B.n345 B.n190 163.367
R1746 B.n349 B.n190 163.367
R1747 B.n350 B.n349 163.367
R1748 B.n351 B.n350 163.367
R1749 B.n351 B.n188 163.367
R1750 B.n355 B.n188 163.367
R1751 B.n356 B.n355 163.367
R1752 B.n357 B.n356 163.367
R1753 B.n357 B.n186 163.367
R1754 B.n361 B.n186 163.367
R1755 B.n362 B.n361 163.367
R1756 B.n363 B.n362 163.367
R1757 B.n363 B.n184 163.367
R1758 B.n367 B.n184 163.367
R1759 B.n368 B.n367 163.367
R1760 B.n369 B.n368 163.367
R1761 B.n369 B.n182 163.367
R1762 B.n373 B.n182 163.367
R1763 B.n374 B.n373 163.367
R1764 B.n375 B.n374 163.367
R1765 B.n375 B.n180 163.367
R1766 B.n379 B.n180 163.367
R1767 B.n380 B.n379 163.367
R1768 B.n381 B.n380 163.367
R1769 B.n381 B.n178 163.367
R1770 B.n388 B.n178 163.367
R1771 B.n389 B.n388 163.367
R1772 B.n390 B.n389 163.367
R1773 B.n390 B.n176 163.367
R1774 B.n394 B.n176 163.367
R1775 B.n395 B.n394 163.367
R1776 B.n396 B.n395 163.367
R1777 B.n396 B.n174 163.367
R1778 B.n400 B.n174 163.367
R1779 B.n401 B.n400 163.367
R1780 B.n402 B.n401 163.367
R1781 B.n402 B.n170 163.367
R1782 B.n407 B.n170 163.367
R1783 B.n408 B.n407 163.367
R1784 B.n409 B.n408 163.367
R1785 B.n409 B.n168 163.367
R1786 B.n413 B.n168 163.367
R1787 B.n414 B.n413 163.367
R1788 B.n415 B.n414 163.367
R1789 B.n415 B.n166 163.367
R1790 B.n419 B.n166 163.367
R1791 B.n420 B.n419 163.367
R1792 B.n421 B.n420 163.367
R1793 B.n421 B.n164 163.367
R1794 B.n425 B.n164 163.367
R1795 B.n426 B.n425 163.367
R1796 B.n427 B.n426 163.367
R1797 B.n427 B.n162 163.367
R1798 B.n431 B.n162 163.367
R1799 B.n432 B.n431 163.367
R1800 B.n433 B.n432 163.367
R1801 B.n433 B.n160 163.367
R1802 B.n437 B.n160 163.367
R1803 B.n438 B.n437 163.367
R1804 B.n439 B.n438 163.367
R1805 B.n439 B.n158 163.367
R1806 B.n443 B.n158 163.367
R1807 B.n444 B.n443 163.367
R1808 B.n445 B.n444 163.367
R1809 B.n445 B.n156 163.367
R1810 B.n449 B.n156 163.367
R1811 B.n450 B.n449 163.367
R1812 B.n451 B.n450 163.367
R1813 B.n451 B.n154 163.367
R1814 B.n455 B.n154 163.367
R1815 B.n456 B.n455 163.367
R1816 B.n457 B.n456 163.367
R1817 B.n457 B.n152 163.367
R1818 B.n461 B.n152 163.367
R1819 B.n462 B.n461 163.367
R1820 B.n463 B.n462 163.367
R1821 B.n463 B.n150 163.367
R1822 B.n467 B.n150 163.367
R1823 B.n468 B.n467 163.367
R1824 B.n469 B.n468 163.367
R1825 B.n469 B.n148 163.367
R1826 B.n473 B.n148 163.367
R1827 B.n474 B.n473 163.367
R1828 B.n475 B.n474 163.367
R1829 B.n475 B.n146 163.367
R1830 B.n479 B.n146 163.367
R1831 B.n480 B.n479 163.367
R1832 B.n481 B.n480 163.367
R1833 B.n481 B.n144 163.367
R1834 B.n485 B.n144 163.367
R1835 B.n641 B.n92 163.367
R1836 B.n637 B.n92 163.367
R1837 B.n637 B.n636 163.367
R1838 B.n636 B.n635 163.367
R1839 B.n635 B.n94 163.367
R1840 B.n631 B.n94 163.367
R1841 B.n631 B.n630 163.367
R1842 B.n630 B.n629 163.367
R1843 B.n629 B.n96 163.367
R1844 B.n625 B.n96 163.367
R1845 B.n625 B.n624 163.367
R1846 B.n624 B.n623 163.367
R1847 B.n623 B.n98 163.367
R1848 B.n619 B.n98 163.367
R1849 B.n619 B.n618 163.367
R1850 B.n618 B.n617 163.367
R1851 B.n617 B.n100 163.367
R1852 B.n613 B.n100 163.367
R1853 B.n613 B.n612 163.367
R1854 B.n612 B.n611 163.367
R1855 B.n611 B.n102 163.367
R1856 B.n607 B.n102 163.367
R1857 B.n607 B.n606 163.367
R1858 B.n606 B.n605 163.367
R1859 B.n605 B.n104 163.367
R1860 B.n601 B.n104 163.367
R1861 B.n601 B.n600 163.367
R1862 B.n600 B.n599 163.367
R1863 B.n599 B.n106 163.367
R1864 B.n595 B.n106 163.367
R1865 B.n595 B.n594 163.367
R1866 B.n594 B.n593 163.367
R1867 B.n593 B.n108 163.367
R1868 B.n589 B.n108 163.367
R1869 B.n589 B.n588 163.367
R1870 B.n588 B.n587 163.367
R1871 B.n587 B.n110 163.367
R1872 B.n583 B.n110 163.367
R1873 B.n583 B.n582 163.367
R1874 B.n582 B.n581 163.367
R1875 B.n581 B.n112 163.367
R1876 B.n577 B.n112 163.367
R1877 B.n577 B.n576 163.367
R1878 B.n576 B.n575 163.367
R1879 B.n575 B.n114 163.367
R1880 B.n571 B.n114 163.367
R1881 B.n571 B.n570 163.367
R1882 B.n570 B.n569 163.367
R1883 B.n569 B.n116 163.367
R1884 B.n565 B.n116 163.367
R1885 B.n565 B.n564 163.367
R1886 B.n564 B.n563 163.367
R1887 B.n563 B.n118 163.367
R1888 B.n559 B.n118 163.367
R1889 B.n559 B.n558 163.367
R1890 B.n558 B.n557 163.367
R1891 B.n557 B.n120 163.367
R1892 B.n553 B.n120 163.367
R1893 B.n553 B.n552 163.367
R1894 B.n552 B.n551 163.367
R1895 B.n551 B.n122 163.367
R1896 B.n547 B.n122 163.367
R1897 B.n547 B.n546 163.367
R1898 B.n546 B.n545 163.367
R1899 B.n545 B.n124 163.367
R1900 B.n541 B.n124 163.367
R1901 B.n541 B.n540 163.367
R1902 B.n540 B.n539 163.367
R1903 B.n539 B.n126 163.367
R1904 B.n535 B.n126 163.367
R1905 B.n535 B.n534 163.367
R1906 B.n534 B.n533 163.367
R1907 B.n533 B.n128 163.367
R1908 B.n529 B.n128 163.367
R1909 B.n529 B.n528 163.367
R1910 B.n528 B.n527 163.367
R1911 B.n527 B.n130 163.367
R1912 B.n523 B.n130 163.367
R1913 B.n523 B.n522 163.367
R1914 B.n522 B.n521 163.367
R1915 B.n521 B.n132 163.367
R1916 B.n517 B.n132 163.367
R1917 B.n517 B.n516 163.367
R1918 B.n516 B.n515 163.367
R1919 B.n515 B.n134 163.367
R1920 B.n511 B.n134 163.367
R1921 B.n511 B.n510 163.367
R1922 B.n510 B.n509 163.367
R1923 B.n509 B.n136 163.367
R1924 B.n505 B.n136 163.367
R1925 B.n505 B.n504 163.367
R1926 B.n504 B.n503 163.367
R1927 B.n503 B.n138 163.367
R1928 B.n499 B.n138 163.367
R1929 B.n499 B.n498 163.367
R1930 B.n498 B.n497 163.367
R1931 B.n497 B.n140 163.367
R1932 B.n493 B.n140 163.367
R1933 B.n493 B.n492 163.367
R1934 B.n492 B.n491 163.367
R1935 B.n491 B.n142 163.367
R1936 B.n487 B.n142 163.367
R1937 B.n487 B.n486 163.367
R1938 B.n818 B.n817 163.367
R1939 B.n817 B.n816 163.367
R1940 B.n816 B.n29 163.367
R1941 B.n812 B.n29 163.367
R1942 B.n812 B.n811 163.367
R1943 B.n811 B.n810 163.367
R1944 B.n810 B.n31 163.367
R1945 B.n806 B.n31 163.367
R1946 B.n806 B.n805 163.367
R1947 B.n805 B.n804 163.367
R1948 B.n804 B.n33 163.367
R1949 B.n800 B.n33 163.367
R1950 B.n800 B.n799 163.367
R1951 B.n799 B.n798 163.367
R1952 B.n798 B.n35 163.367
R1953 B.n794 B.n35 163.367
R1954 B.n794 B.n793 163.367
R1955 B.n793 B.n792 163.367
R1956 B.n792 B.n37 163.367
R1957 B.n788 B.n37 163.367
R1958 B.n788 B.n787 163.367
R1959 B.n787 B.n786 163.367
R1960 B.n786 B.n39 163.367
R1961 B.n782 B.n39 163.367
R1962 B.n782 B.n781 163.367
R1963 B.n781 B.n780 163.367
R1964 B.n780 B.n41 163.367
R1965 B.n776 B.n41 163.367
R1966 B.n776 B.n775 163.367
R1967 B.n775 B.n774 163.367
R1968 B.n774 B.n43 163.367
R1969 B.n770 B.n43 163.367
R1970 B.n770 B.n769 163.367
R1971 B.n769 B.n768 163.367
R1972 B.n768 B.n45 163.367
R1973 B.n764 B.n45 163.367
R1974 B.n764 B.n763 163.367
R1975 B.n763 B.n762 163.367
R1976 B.n762 B.n47 163.367
R1977 B.n758 B.n47 163.367
R1978 B.n758 B.n757 163.367
R1979 B.n757 B.n756 163.367
R1980 B.n756 B.n49 163.367
R1981 B.n752 B.n49 163.367
R1982 B.n752 B.n751 163.367
R1983 B.n751 B.n750 163.367
R1984 B.n750 B.n51 163.367
R1985 B.n746 B.n51 163.367
R1986 B.n746 B.n745 163.367
R1987 B.n745 B.n744 163.367
R1988 B.n744 B.n53 163.367
R1989 B.n740 B.n53 163.367
R1990 B.n740 B.n739 163.367
R1991 B.n739 B.n738 163.367
R1992 B.n738 B.n55 163.367
R1993 B.n734 B.n55 163.367
R1994 B.n734 B.n733 163.367
R1995 B.n733 B.n732 163.367
R1996 B.n732 B.n60 163.367
R1997 B.n728 B.n60 163.367
R1998 B.n728 B.n727 163.367
R1999 B.n727 B.n726 163.367
R2000 B.n726 B.n62 163.367
R2001 B.n721 B.n62 163.367
R2002 B.n721 B.n720 163.367
R2003 B.n720 B.n719 163.367
R2004 B.n719 B.n66 163.367
R2005 B.n715 B.n66 163.367
R2006 B.n715 B.n714 163.367
R2007 B.n714 B.n713 163.367
R2008 B.n713 B.n68 163.367
R2009 B.n709 B.n68 163.367
R2010 B.n709 B.n708 163.367
R2011 B.n708 B.n707 163.367
R2012 B.n707 B.n70 163.367
R2013 B.n703 B.n70 163.367
R2014 B.n703 B.n702 163.367
R2015 B.n702 B.n701 163.367
R2016 B.n701 B.n72 163.367
R2017 B.n697 B.n72 163.367
R2018 B.n697 B.n696 163.367
R2019 B.n696 B.n695 163.367
R2020 B.n695 B.n74 163.367
R2021 B.n691 B.n74 163.367
R2022 B.n691 B.n690 163.367
R2023 B.n690 B.n689 163.367
R2024 B.n689 B.n76 163.367
R2025 B.n685 B.n76 163.367
R2026 B.n685 B.n684 163.367
R2027 B.n684 B.n683 163.367
R2028 B.n683 B.n78 163.367
R2029 B.n679 B.n78 163.367
R2030 B.n679 B.n678 163.367
R2031 B.n678 B.n677 163.367
R2032 B.n677 B.n80 163.367
R2033 B.n673 B.n80 163.367
R2034 B.n673 B.n672 163.367
R2035 B.n672 B.n671 163.367
R2036 B.n671 B.n82 163.367
R2037 B.n667 B.n82 163.367
R2038 B.n667 B.n666 163.367
R2039 B.n666 B.n665 163.367
R2040 B.n665 B.n84 163.367
R2041 B.n661 B.n84 163.367
R2042 B.n661 B.n660 163.367
R2043 B.n660 B.n659 163.367
R2044 B.n659 B.n86 163.367
R2045 B.n655 B.n86 163.367
R2046 B.n655 B.n654 163.367
R2047 B.n654 B.n653 163.367
R2048 B.n653 B.n88 163.367
R2049 B.n649 B.n88 163.367
R2050 B.n649 B.n648 163.367
R2051 B.n648 B.n647 163.367
R2052 B.n647 B.n90 163.367
R2053 B.n643 B.n90 163.367
R2054 B.n643 B.n642 163.367
R2055 B.n822 B.n27 163.367
R2056 B.n823 B.n822 163.367
R2057 B.n824 B.n823 163.367
R2058 B.n824 B.n25 163.367
R2059 B.n828 B.n25 163.367
R2060 B.n829 B.n828 163.367
R2061 B.n830 B.n829 163.367
R2062 B.n830 B.n23 163.367
R2063 B.n834 B.n23 163.367
R2064 B.n835 B.n834 163.367
R2065 B.n836 B.n835 163.367
R2066 B.n836 B.n21 163.367
R2067 B.n840 B.n21 163.367
R2068 B.n841 B.n840 163.367
R2069 B.n842 B.n841 163.367
R2070 B.n842 B.n19 163.367
R2071 B.n846 B.n19 163.367
R2072 B.n847 B.n846 163.367
R2073 B.n848 B.n847 163.367
R2074 B.n848 B.n17 163.367
R2075 B.n852 B.n17 163.367
R2076 B.n853 B.n852 163.367
R2077 B.n854 B.n853 163.367
R2078 B.n854 B.n15 163.367
R2079 B.n858 B.n15 163.367
R2080 B.n859 B.n858 163.367
R2081 B.n860 B.n859 163.367
R2082 B.n860 B.n13 163.367
R2083 B.n864 B.n13 163.367
R2084 B.n865 B.n864 163.367
R2085 B.n866 B.n865 163.367
R2086 B.n866 B.n11 163.367
R2087 B.n870 B.n11 163.367
R2088 B.n871 B.n870 163.367
R2089 B.n872 B.n871 163.367
R2090 B.n872 B.n9 163.367
R2091 B.n876 B.n9 163.367
R2092 B.n877 B.n876 163.367
R2093 B.n878 B.n877 163.367
R2094 B.n878 B.n7 163.367
R2095 B.n882 B.n7 163.367
R2096 B.n883 B.n882 163.367
R2097 B.n884 B.n883 163.367
R2098 B.n884 B.n5 163.367
R2099 B.n888 B.n5 163.367
R2100 B.n889 B.n888 163.367
R2101 B.n890 B.n889 163.367
R2102 B.n890 B.n3 163.367
R2103 B.n894 B.n3 163.367
R2104 B.n895 B.n894 163.367
R2105 B.n230 B.n2 163.367
R2106 B.n231 B.n230 163.367
R2107 B.n231 B.n228 163.367
R2108 B.n235 B.n228 163.367
R2109 B.n236 B.n235 163.367
R2110 B.n237 B.n236 163.367
R2111 B.n237 B.n226 163.367
R2112 B.n241 B.n226 163.367
R2113 B.n242 B.n241 163.367
R2114 B.n243 B.n242 163.367
R2115 B.n243 B.n224 163.367
R2116 B.n247 B.n224 163.367
R2117 B.n248 B.n247 163.367
R2118 B.n249 B.n248 163.367
R2119 B.n249 B.n222 163.367
R2120 B.n253 B.n222 163.367
R2121 B.n254 B.n253 163.367
R2122 B.n255 B.n254 163.367
R2123 B.n255 B.n220 163.367
R2124 B.n259 B.n220 163.367
R2125 B.n260 B.n259 163.367
R2126 B.n261 B.n260 163.367
R2127 B.n261 B.n218 163.367
R2128 B.n265 B.n218 163.367
R2129 B.n266 B.n265 163.367
R2130 B.n267 B.n266 163.367
R2131 B.n267 B.n216 163.367
R2132 B.n271 B.n216 163.367
R2133 B.n272 B.n271 163.367
R2134 B.n273 B.n272 163.367
R2135 B.n273 B.n214 163.367
R2136 B.n277 B.n214 163.367
R2137 B.n278 B.n277 163.367
R2138 B.n279 B.n278 163.367
R2139 B.n279 B.n212 163.367
R2140 B.n283 B.n212 163.367
R2141 B.n284 B.n283 163.367
R2142 B.n285 B.n284 163.367
R2143 B.n285 B.n210 163.367
R2144 B.n289 B.n210 163.367
R2145 B.n290 B.n289 163.367
R2146 B.n291 B.n290 163.367
R2147 B.n291 B.n208 163.367
R2148 B.n295 B.n208 163.367
R2149 B.n296 B.n295 163.367
R2150 B.n297 B.n296 163.367
R2151 B.n297 B.n206 163.367
R2152 B.n301 B.n206 163.367
R2153 B.n302 B.n301 163.367
R2154 B.n303 B.n302 163.367
R2155 B.n385 B.n384 71.1763
R2156 B.n172 B.n171 71.1763
R2157 B.n64 B.n63 71.1763
R2158 B.n57 B.n56 71.1763
R2159 B.n386 B.n385 59.5399
R2160 B.n404 B.n172 59.5399
R2161 B.n723 B.n64 59.5399
R2162 B.n58 B.n57 59.5399
R2163 B.n820 B.n819 28.8785
R2164 B.n640 B.n91 28.8785
R2165 B.n305 B.n304 28.8785
R2166 B.n484 B.n143 28.8785
R2167 B B.n897 18.0485
R2168 B.n821 B.n820 10.6151
R2169 B.n821 B.n26 10.6151
R2170 B.n825 B.n26 10.6151
R2171 B.n826 B.n825 10.6151
R2172 B.n827 B.n826 10.6151
R2173 B.n827 B.n24 10.6151
R2174 B.n831 B.n24 10.6151
R2175 B.n832 B.n831 10.6151
R2176 B.n833 B.n832 10.6151
R2177 B.n833 B.n22 10.6151
R2178 B.n837 B.n22 10.6151
R2179 B.n838 B.n837 10.6151
R2180 B.n839 B.n838 10.6151
R2181 B.n839 B.n20 10.6151
R2182 B.n843 B.n20 10.6151
R2183 B.n844 B.n843 10.6151
R2184 B.n845 B.n844 10.6151
R2185 B.n845 B.n18 10.6151
R2186 B.n849 B.n18 10.6151
R2187 B.n850 B.n849 10.6151
R2188 B.n851 B.n850 10.6151
R2189 B.n851 B.n16 10.6151
R2190 B.n855 B.n16 10.6151
R2191 B.n856 B.n855 10.6151
R2192 B.n857 B.n856 10.6151
R2193 B.n857 B.n14 10.6151
R2194 B.n861 B.n14 10.6151
R2195 B.n862 B.n861 10.6151
R2196 B.n863 B.n862 10.6151
R2197 B.n863 B.n12 10.6151
R2198 B.n867 B.n12 10.6151
R2199 B.n868 B.n867 10.6151
R2200 B.n869 B.n868 10.6151
R2201 B.n869 B.n10 10.6151
R2202 B.n873 B.n10 10.6151
R2203 B.n874 B.n873 10.6151
R2204 B.n875 B.n874 10.6151
R2205 B.n875 B.n8 10.6151
R2206 B.n879 B.n8 10.6151
R2207 B.n880 B.n879 10.6151
R2208 B.n881 B.n880 10.6151
R2209 B.n881 B.n6 10.6151
R2210 B.n885 B.n6 10.6151
R2211 B.n886 B.n885 10.6151
R2212 B.n887 B.n886 10.6151
R2213 B.n887 B.n4 10.6151
R2214 B.n891 B.n4 10.6151
R2215 B.n892 B.n891 10.6151
R2216 B.n893 B.n892 10.6151
R2217 B.n893 B.n0 10.6151
R2218 B.n819 B.n28 10.6151
R2219 B.n815 B.n28 10.6151
R2220 B.n815 B.n814 10.6151
R2221 B.n814 B.n813 10.6151
R2222 B.n813 B.n30 10.6151
R2223 B.n809 B.n30 10.6151
R2224 B.n809 B.n808 10.6151
R2225 B.n808 B.n807 10.6151
R2226 B.n807 B.n32 10.6151
R2227 B.n803 B.n32 10.6151
R2228 B.n803 B.n802 10.6151
R2229 B.n802 B.n801 10.6151
R2230 B.n801 B.n34 10.6151
R2231 B.n797 B.n34 10.6151
R2232 B.n797 B.n796 10.6151
R2233 B.n796 B.n795 10.6151
R2234 B.n795 B.n36 10.6151
R2235 B.n791 B.n36 10.6151
R2236 B.n791 B.n790 10.6151
R2237 B.n790 B.n789 10.6151
R2238 B.n789 B.n38 10.6151
R2239 B.n785 B.n38 10.6151
R2240 B.n785 B.n784 10.6151
R2241 B.n784 B.n783 10.6151
R2242 B.n783 B.n40 10.6151
R2243 B.n779 B.n40 10.6151
R2244 B.n779 B.n778 10.6151
R2245 B.n778 B.n777 10.6151
R2246 B.n777 B.n42 10.6151
R2247 B.n773 B.n42 10.6151
R2248 B.n773 B.n772 10.6151
R2249 B.n772 B.n771 10.6151
R2250 B.n771 B.n44 10.6151
R2251 B.n767 B.n44 10.6151
R2252 B.n767 B.n766 10.6151
R2253 B.n766 B.n765 10.6151
R2254 B.n765 B.n46 10.6151
R2255 B.n761 B.n46 10.6151
R2256 B.n761 B.n760 10.6151
R2257 B.n760 B.n759 10.6151
R2258 B.n759 B.n48 10.6151
R2259 B.n755 B.n48 10.6151
R2260 B.n755 B.n754 10.6151
R2261 B.n754 B.n753 10.6151
R2262 B.n753 B.n50 10.6151
R2263 B.n749 B.n50 10.6151
R2264 B.n749 B.n748 10.6151
R2265 B.n748 B.n747 10.6151
R2266 B.n747 B.n52 10.6151
R2267 B.n743 B.n52 10.6151
R2268 B.n743 B.n742 10.6151
R2269 B.n742 B.n741 10.6151
R2270 B.n741 B.n54 10.6151
R2271 B.n737 B.n736 10.6151
R2272 B.n736 B.n735 10.6151
R2273 B.n735 B.n59 10.6151
R2274 B.n731 B.n59 10.6151
R2275 B.n731 B.n730 10.6151
R2276 B.n730 B.n729 10.6151
R2277 B.n729 B.n61 10.6151
R2278 B.n725 B.n61 10.6151
R2279 B.n725 B.n724 10.6151
R2280 B.n722 B.n65 10.6151
R2281 B.n718 B.n65 10.6151
R2282 B.n718 B.n717 10.6151
R2283 B.n717 B.n716 10.6151
R2284 B.n716 B.n67 10.6151
R2285 B.n712 B.n67 10.6151
R2286 B.n712 B.n711 10.6151
R2287 B.n711 B.n710 10.6151
R2288 B.n710 B.n69 10.6151
R2289 B.n706 B.n69 10.6151
R2290 B.n706 B.n705 10.6151
R2291 B.n705 B.n704 10.6151
R2292 B.n704 B.n71 10.6151
R2293 B.n700 B.n71 10.6151
R2294 B.n700 B.n699 10.6151
R2295 B.n699 B.n698 10.6151
R2296 B.n698 B.n73 10.6151
R2297 B.n694 B.n73 10.6151
R2298 B.n694 B.n693 10.6151
R2299 B.n693 B.n692 10.6151
R2300 B.n692 B.n75 10.6151
R2301 B.n688 B.n75 10.6151
R2302 B.n688 B.n687 10.6151
R2303 B.n687 B.n686 10.6151
R2304 B.n686 B.n77 10.6151
R2305 B.n682 B.n77 10.6151
R2306 B.n682 B.n681 10.6151
R2307 B.n681 B.n680 10.6151
R2308 B.n680 B.n79 10.6151
R2309 B.n676 B.n79 10.6151
R2310 B.n676 B.n675 10.6151
R2311 B.n675 B.n674 10.6151
R2312 B.n674 B.n81 10.6151
R2313 B.n670 B.n81 10.6151
R2314 B.n670 B.n669 10.6151
R2315 B.n669 B.n668 10.6151
R2316 B.n668 B.n83 10.6151
R2317 B.n664 B.n83 10.6151
R2318 B.n664 B.n663 10.6151
R2319 B.n663 B.n662 10.6151
R2320 B.n662 B.n85 10.6151
R2321 B.n658 B.n85 10.6151
R2322 B.n658 B.n657 10.6151
R2323 B.n657 B.n656 10.6151
R2324 B.n656 B.n87 10.6151
R2325 B.n652 B.n87 10.6151
R2326 B.n652 B.n651 10.6151
R2327 B.n651 B.n650 10.6151
R2328 B.n650 B.n89 10.6151
R2329 B.n646 B.n89 10.6151
R2330 B.n646 B.n645 10.6151
R2331 B.n645 B.n644 10.6151
R2332 B.n644 B.n91 10.6151
R2333 B.n640 B.n639 10.6151
R2334 B.n639 B.n638 10.6151
R2335 B.n638 B.n93 10.6151
R2336 B.n634 B.n93 10.6151
R2337 B.n634 B.n633 10.6151
R2338 B.n633 B.n632 10.6151
R2339 B.n632 B.n95 10.6151
R2340 B.n628 B.n95 10.6151
R2341 B.n628 B.n627 10.6151
R2342 B.n627 B.n626 10.6151
R2343 B.n626 B.n97 10.6151
R2344 B.n622 B.n97 10.6151
R2345 B.n622 B.n621 10.6151
R2346 B.n621 B.n620 10.6151
R2347 B.n620 B.n99 10.6151
R2348 B.n616 B.n99 10.6151
R2349 B.n616 B.n615 10.6151
R2350 B.n615 B.n614 10.6151
R2351 B.n614 B.n101 10.6151
R2352 B.n610 B.n101 10.6151
R2353 B.n610 B.n609 10.6151
R2354 B.n609 B.n608 10.6151
R2355 B.n608 B.n103 10.6151
R2356 B.n604 B.n103 10.6151
R2357 B.n604 B.n603 10.6151
R2358 B.n603 B.n602 10.6151
R2359 B.n602 B.n105 10.6151
R2360 B.n598 B.n105 10.6151
R2361 B.n598 B.n597 10.6151
R2362 B.n597 B.n596 10.6151
R2363 B.n596 B.n107 10.6151
R2364 B.n592 B.n107 10.6151
R2365 B.n592 B.n591 10.6151
R2366 B.n591 B.n590 10.6151
R2367 B.n590 B.n109 10.6151
R2368 B.n586 B.n109 10.6151
R2369 B.n586 B.n585 10.6151
R2370 B.n585 B.n584 10.6151
R2371 B.n584 B.n111 10.6151
R2372 B.n580 B.n111 10.6151
R2373 B.n580 B.n579 10.6151
R2374 B.n579 B.n578 10.6151
R2375 B.n578 B.n113 10.6151
R2376 B.n574 B.n113 10.6151
R2377 B.n574 B.n573 10.6151
R2378 B.n573 B.n572 10.6151
R2379 B.n572 B.n115 10.6151
R2380 B.n568 B.n115 10.6151
R2381 B.n568 B.n567 10.6151
R2382 B.n567 B.n566 10.6151
R2383 B.n566 B.n117 10.6151
R2384 B.n562 B.n117 10.6151
R2385 B.n562 B.n561 10.6151
R2386 B.n561 B.n560 10.6151
R2387 B.n560 B.n119 10.6151
R2388 B.n556 B.n119 10.6151
R2389 B.n556 B.n555 10.6151
R2390 B.n555 B.n554 10.6151
R2391 B.n554 B.n121 10.6151
R2392 B.n550 B.n121 10.6151
R2393 B.n550 B.n549 10.6151
R2394 B.n549 B.n548 10.6151
R2395 B.n548 B.n123 10.6151
R2396 B.n544 B.n123 10.6151
R2397 B.n544 B.n543 10.6151
R2398 B.n543 B.n542 10.6151
R2399 B.n542 B.n125 10.6151
R2400 B.n538 B.n125 10.6151
R2401 B.n538 B.n537 10.6151
R2402 B.n537 B.n536 10.6151
R2403 B.n536 B.n127 10.6151
R2404 B.n532 B.n127 10.6151
R2405 B.n532 B.n531 10.6151
R2406 B.n531 B.n530 10.6151
R2407 B.n530 B.n129 10.6151
R2408 B.n526 B.n129 10.6151
R2409 B.n526 B.n525 10.6151
R2410 B.n525 B.n524 10.6151
R2411 B.n524 B.n131 10.6151
R2412 B.n520 B.n131 10.6151
R2413 B.n520 B.n519 10.6151
R2414 B.n519 B.n518 10.6151
R2415 B.n518 B.n133 10.6151
R2416 B.n514 B.n133 10.6151
R2417 B.n514 B.n513 10.6151
R2418 B.n513 B.n512 10.6151
R2419 B.n512 B.n135 10.6151
R2420 B.n508 B.n135 10.6151
R2421 B.n508 B.n507 10.6151
R2422 B.n507 B.n506 10.6151
R2423 B.n506 B.n137 10.6151
R2424 B.n502 B.n137 10.6151
R2425 B.n502 B.n501 10.6151
R2426 B.n501 B.n500 10.6151
R2427 B.n500 B.n139 10.6151
R2428 B.n496 B.n139 10.6151
R2429 B.n496 B.n495 10.6151
R2430 B.n495 B.n494 10.6151
R2431 B.n494 B.n141 10.6151
R2432 B.n490 B.n141 10.6151
R2433 B.n490 B.n489 10.6151
R2434 B.n489 B.n488 10.6151
R2435 B.n488 B.n143 10.6151
R2436 B.n229 B.n1 10.6151
R2437 B.n232 B.n229 10.6151
R2438 B.n233 B.n232 10.6151
R2439 B.n234 B.n233 10.6151
R2440 B.n234 B.n227 10.6151
R2441 B.n238 B.n227 10.6151
R2442 B.n239 B.n238 10.6151
R2443 B.n240 B.n239 10.6151
R2444 B.n240 B.n225 10.6151
R2445 B.n244 B.n225 10.6151
R2446 B.n245 B.n244 10.6151
R2447 B.n246 B.n245 10.6151
R2448 B.n246 B.n223 10.6151
R2449 B.n250 B.n223 10.6151
R2450 B.n251 B.n250 10.6151
R2451 B.n252 B.n251 10.6151
R2452 B.n252 B.n221 10.6151
R2453 B.n256 B.n221 10.6151
R2454 B.n257 B.n256 10.6151
R2455 B.n258 B.n257 10.6151
R2456 B.n258 B.n219 10.6151
R2457 B.n262 B.n219 10.6151
R2458 B.n263 B.n262 10.6151
R2459 B.n264 B.n263 10.6151
R2460 B.n264 B.n217 10.6151
R2461 B.n268 B.n217 10.6151
R2462 B.n269 B.n268 10.6151
R2463 B.n270 B.n269 10.6151
R2464 B.n270 B.n215 10.6151
R2465 B.n274 B.n215 10.6151
R2466 B.n275 B.n274 10.6151
R2467 B.n276 B.n275 10.6151
R2468 B.n276 B.n213 10.6151
R2469 B.n280 B.n213 10.6151
R2470 B.n281 B.n280 10.6151
R2471 B.n282 B.n281 10.6151
R2472 B.n282 B.n211 10.6151
R2473 B.n286 B.n211 10.6151
R2474 B.n287 B.n286 10.6151
R2475 B.n288 B.n287 10.6151
R2476 B.n288 B.n209 10.6151
R2477 B.n292 B.n209 10.6151
R2478 B.n293 B.n292 10.6151
R2479 B.n294 B.n293 10.6151
R2480 B.n294 B.n207 10.6151
R2481 B.n298 B.n207 10.6151
R2482 B.n299 B.n298 10.6151
R2483 B.n300 B.n299 10.6151
R2484 B.n300 B.n205 10.6151
R2485 B.n304 B.n205 10.6151
R2486 B.n306 B.n305 10.6151
R2487 B.n306 B.n203 10.6151
R2488 B.n310 B.n203 10.6151
R2489 B.n311 B.n310 10.6151
R2490 B.n312 B.n311 10.6151
R2491 B.n312 B.n201 10.6151
R2492 B.n316 B.n201 10.6151
R2493 B.n317 B.n316 10.6151
R2494 B.n318 B.n317 10.6151
R2495 B.n318 B.n199 10.6151
R2496 B.n322 B.n199 10.6151
R2497 B.n323 B.n322 10.6151
R2498 B.n324 B.n323 10.6151
R2499 B.n324 B.n197 10.6151
R2500 B.n328 B.n197 10.6151
R2501 B.n329 B.n328 10.6151
R2502 B.n330 B.n329 10.6151
R2503 B.n330 B.n195 10.6151
R2504 B.n334 B.n195 10.6151
R2505 B.n335 B.n334 10.6151
R2506 B.n336 B.n335 10.6151
R2507 B.n336 B.n193 10.6151
R2508 B.n340 B.n193 10.6151
R2509 B.n341 B.n340 10.6151
R2510 B.n342 B.n341 10.6151
R2511 B.n342 B.n191 10.6151
R2512 B.n346 B.n191 10.6151
R2513 B.n347 B.n346 10.6151
R2514 B.n348 B.n347 10.6151
R2515 B.n348 B.n189 10.6151
R2516 B.n352 B.n189 10.6151
R2517 B.n353 B.n352 10.6151
R2518 B.n354 B.n353 10.6151
R2519 B.n354 B.n187 10.6151
R2520 B.n358 B.n187 10.6151
R2521 B.n359 B.n358 10.6151
R2522 B.n360 B.n359 10.6151
R2523 B.n360 B.n185 10.6151
R2524 B.n364 B.n185 10.6151
R2525 B.n365 B.n364 10.6151
R2526 B.n366 B.n365 10.6151
R2527 B.n366 B.n183 10.6151
R2528 B.n370 B.n183 10.6151
R2529 B.n371 B.n370 10.6151
R2530 B.n372 B.n371 10.6151
R2531 B.n372 B.n181 10.6151
R2532 B.n376 B.n181 10.6151
R2533 B.n377 B.n376 10.6151
R2534 B.n378 B.n377 10.6151
R2535 B.n378 B.n179 10.6151
R2536 B.n382 B.n179 10.6151
R2537 B.n383 B.n382 10.6151
R2538 B.n387 B.n383 10.6151
R2539 B.n391 B.n177 10.6151
R2540 B.n392 B.n391 10.6151
R2541 B.n393 B.n392 10.6151
R2542 B.n393 B.n175 10.6151
R2543 B.n397 B.n175 10.6151
R2544 B.n398 B.n397 10.6151
R2545 B.n399 B.n398 10.6151
R2546 B.n399 B.n173 10.6151
R2547 B.n403 B.n173 10.6151
R2548 B.n406 B.n405 10.6151
R2549 B.n406 B.n169 10.6151
R2550 B.n410 B.n169 10.6151
R2551 B.n411 B.n410 10.6151
R2552 B.n412 B.n411 10.6151
R2553 B.n412 B.n167 10.6151
R2554 B.n416 B.n167 10.6151
R2555 B.n417 B.n416 10.6151
R2556 B.n418 B.n417 10.6151
R2557 B.n418 B.n165 10.6151
R2558 B.n422 B.n165 10.6151
R2559 B.n423 B.n422 10.6151
R2560 B.n424 B.n423 10.6151
R2561 B.n424 B.n163 10.6151
R2562 B.n428 B.n163 10.6151
R2563 B.n429 B.n428 10.6151
R2564 B.n430 B.n429 10.6151
R2565 B.n430 B.n161 10.6151
R2566 B.n434 B.n161 10.6151
R2567 B.n435 B.n434 10.6151
R2568 B.n436 B.n435 10.6151
R2569 B.n436 B.n159 10.6151
R2570 B.n440 B.n159 10.6151
R2571 B.n441 B.n440 10.6151
R2572 B.n442 B.n441 10.6151
R2573 B.n442 B.n157 10.6151
R2574 B.n446 B.n157 10.6151
R2575 B.n447 B.n446 10.6151
R2576 B.n448 B.n447 10.6151
R2577 B.n448 B.n155 10.6151
R2578 B.n452 B.n155 10.6151
R2579 B.n453 B.n452 10.6151
R2580 B.n454 B.n453 10.6151
R2581 B.n454 B.n153 10.6151
R2582 B.n458 B.n153 10.6151
R2583 B.n459 B.n458 10.6151
R2584 B.n460 B.n459 10.6151
R2585 B.n460 B.n151 10.6151
R2586 B.n464 B.n151 10.6151
R2587 B.n465 B.n464 10.6151
R2588 B.n466 B.n465 10.6151
R2589 B.n466 B.n149 10.6151
R2590 B.n470 B.n149 10.6151
R2591 B.n471 B.n470 10.6151
R2592 B.n472 B.n471 10.6151
R2593 B.n472 B.n147 10.6151
R2594 B.n476 B.n147 10.6151
R2595 B.n477 B.n476 10.6151
R2596 B.n478 B.n477 10.6151
R2597 B.n478 B.n145 10.6151
R2598 B.n482 B.n145 10.6151
R2599 B.n483 B.n482 10.6151
R2600 B.n484 B.n483 10.6151
R2601 B.n58 B.n54 9.36635
R2602 B.n723 B.n722 9.36635
R2603 B.n387 B.n386 9.36635
R2604 B.n405 B.n404 9.36635
R2605 B.n897 B.n0 8.11757
R2606 B.n897 B.n1 8.11757
R2607 B.n737 B.n58 1.24928
R2608 B.n724 B.n723 1.24928
R2609 B.n386 B.n177 1.24928
R2610 B.n404 B.n403 1.24928
C0 VTAIL VDD1 9.3593f
C1 B VP 2.22785f
C2 B VDD1 2.62629f
C3 VDD1 VP 9.72042f
C4 w_n3906_n4216# VN 7.656971f
C5 w_n3906_n4216# VDD2 2.87197f
C6 w_n3906_n4216# VTAIL 3.61939f
C7 w_n3906_n4216# B 11.8868f
C8 w_n3906_n4216# VP 8.164021f
C9 w_n3906_n4216# VDD1 2.76325f
C10 VDD2 VN 9.3545f
C11 VTAIL VN 9.494269f
C12 VTAIL VDD2 9.41499f
C13 B VN 1.37755f
C14 B VDD2 2.71813f
C15 VP VN 8.42986f
C16 VDD2 VP 0.521761f
C17 B VTAIL 4.96906f
C18 VDD1 VN 0.152167f
C19 VDD1 VDD2 1.69661f
C20 VTAIL VP 9.50855f
C21 VDD2 VSUBS 2.20151f
C22 VDD1 VSUBS 2.198644f
C23 VTAIL VSUBS 1.485307f
C24 VN VSUBS 6.70643f
C25 VP VSUBS 3.66557f
C26 B VSUBS 5.726858f
C27 w_n3906_n4216# VSUBS 0.20169p
C28 B.n0 VSUBS 0.006739f
C29 B.n1 VSUBS 0.006739f
C30 B.n2 VSUBS 0.009967f
C31 B.n3 VSUBS 0.007638f
C32 B.n4 VSUBS 0.007638f
C33 B.n5 VSUBS 0.007638f
C34 B.n6 VSUBS 0.007638f
C35 B.n7 VSUBS 0.007638f
C36 B.n8 VSUBS 0.007638f
C37 B.n9 VSUBS 0.007638f
C38 B.n10 VSUBS 0.007638f
C39 B.n11 VSUBS 0.007638f
C40 B.n12 VSUBS 0.007638f
C41 B.n13 VSUBS 0.007638f
C42 B.n14 VSUBS 0.007638f
C43 B.n15 VSUBS 0.007638f
C44 B.n16 VSUBS 0.007638f
C45 B.n17 VSUBS 0.007638f
C46 B.n18 VSUBS 0.007638f
C47 B.n19 VSUBS 0.007638f
C48 B.n20 VSUBS 0.007638f
C49 B.n21 VSUBS 0.007638f
C50 B.n22 VSUBS 0.007638f
C51 B.n23 VSUBS 0.007638f
C52 B.n24 VSUBS 0.007638f
C53 B.n25 VSUBS 0.007638f
C54 B.n26 VSUBS 0.007638f
C55 B.n27 VSUBS 0.016101f
C56 B.n28 VSUBS 0.007638f
C57 B.n29 VSUBS 0.007638f
C58 B.n30 VSUBS 0.007638f
C59 B.n31 VSUBS 0.007638f
C60 B.n32 VSUBS 0.007638f
C61 B.n33 VSUBS 0.007638f
C62 B.n34 VSUBS 0.007638f
C63 B.n35 VSUBS 0.007638f
C64 B.n36 VSUBS 0.007638f
C65 B.n37 VSUBS 0.007638f
C66 B.n38 VSUBS 0.007638f
C67 B.n39 VSUBS 0.007638f
C68 B.n40 VSUBS 0.007638f
C69 B.n41 VSUBS 0.007638f
C70 B.n42 VSUBS 0.007638f
C71 B.n43 VSUBS 0.007638f
C72 B.n44 VSUBS 0.007638f
C73 B.n45 VSUBS 0.007638f
C74 B.n46 VSUBS 0.007638f
C75 B.n47 VSUBS 0.007638f
C76 B.n48 VSUBS 0.007638f
C77 B.n49 VSUBS 0.007638f
C78 B.n50 VSUBS 0.007638f
C79 B.n51 VSUBS 0.007638f
C80 B.n52 VSUBS 0.007638f
C81 B.n53 VSUBS 0.007638f
C82 B.n54 VSUBS 0.007189f
C83 B.n55 VSUBS 0.007638f
C84 B.t4 VSUBS 0.337164f
C85 B.t5 VSUBS 0.381722f
C86 B.t3 VSUBS 2.69081f
C87 B.n56 VSUBS 0.603381f
C88 B.n57 VSUBS 0.338495f
C89 B.n58 VSUBS 0.017696f
C90 B.n59 VSUBS 0.007638f
C91 B.n60 VSUBS 0.007638f
C92 B.n61 VSUBS 0.007638f
C93 B.n62 VSUBS 0.007638f
C94 B.t1 VSUBS 0.337168f
C95 B.t2 VSUBS 0.381725f
C96 B.t0 VSUBS 2.69081f
C97 B.n63 VSUBS 0.603378f
C98 B.n64 VSUBS 0.338491f
C99 B.n65 VSUBS 0.007638f
C100 B.n66 VSUBS 0.007638f
C101 B.n67 VSUBS 0.007638f
C102 B.n68 VSUBS 0.007638f
C103 B.n69 VSUBS 0.007638f
C104 B.n70 VSUBS 0.007638f
C105 B.n71 VSUBS 0.007638f
C106 B.n72 VSUBS 0.007638f
C107 B.n73 VSUBS 0.007638f
C108 B.n74 VSUBS 0.007638f
C109 B.n75 VSUBS 0.007638f
C110 B.n76 VSUBS 0.007638f
C111 B.n77 VSUBS 0.007638f
C112 B.n78 VSUBS 0.007638f
C113 B.n79 VSUBS 0.007638f
C114 B.n80 VSUBS 0.007638f
C115 B.n81 VSUBS 0.007638f
C116 B.n82 VSUBS 0.007638f
C117 B.n83 VSUBS 0.007638f
C118 B.n84 VSUBS 0.007638f
C119 B.n85 VSUBS 0.007638f
C120 B.n86 VSUBS 0.007638f
C121 B.n87 VSUBS 0.007638f
C122 B.n88 VSUBS 0.007638f
C123 B.n89 VSUBS 0.007638f
C124 B.n90 VSUBS 0.007638f
C125 B.n91 VSUBS 0.016922f
C126 B.n92 VSUBS 0.007638f
C127 B.n93 VSUBS 0.007638f
C128 B.n94 VSUBS 0.007638f
C129 B.n95 VSUBS 0.007638f
C130 B.n96 VSUBS 0.007638f
C131 B.n97 VSUBS 0.007638f
C132 B.n98 VSUBS 0.007638f
C133 B.n99 VSUBS 0.007638f
C134 B.n100 VSUBS 0.007638f
C135 B.n101 VSUBS 0.007638f
C136 B.n102 VSUBS 0.007638f
C137 B.n103 VSUBS 0.007638f
C138 B.n104 VSUBS 0.007638f
C139 B.n105 VSUBS 0.007638f
C140 B.n106 VSUBS 0.007638f
C141 B.n107 VSUBS 0.007638f
C142 B.n108 VSUBS 0.007638f
C143 B.n109 VSUBS 0.007638f
C144 B.n110 VSUBS 0.007638f
C145 B.n111 VSUBS 0.007638f
C146 B.n112 VSUBS 0.007638f
C147 B.n113 VSUBS 0.007638f
C148 B.n114 VSUBS 0.007638f
C149 B.n115 VSUBS 0.007638f
C150 B.n116 VSUBS 0.007638f
C151 B.n117 VSUBS 0.007638f
C152 B.n118 VSUBS 0.007638f
C153 B.n119 VSUBS 0.007638f
C154 B.n120 VSUBS 0.007638f
C155 B.n121 VSUBS 0.007638f
C156 B.n122 VSUBS 0.007638f
C157 B.n123 VSUBS 0.007638f
C158 B.n124 VSUBS 0.007638f
C159 B.n125 VSUBS 0.007638f
C160 B.n126 VSUBS 0.007638f
C161 B.n127 VSUBS 0.007638f
C162 B.n128 VSUBS 0.007638f
C163 B.n129 VSUBS 0.007638f
C164 B.n130 VSUBS 0.007638f
C165 B.n131 VSUBS 0.007638f
C166 B.n132 VSUBS 0.007638f
C167 B.n133 VSUBS 0.007638f
C168 B.n134 VSUBS 0.007638f
C169 B.n135 VSUBS 0.007638f
C170 B.n136 VSUBS 0.007638f
C171 B.n137 VSUBS 0.007638f
C172 B.n138 VSUBS 0.007638f
C173 B.n139 VSUBS 0.007638f
C174 B.n140 VSUBS 0.007638f
C175 B.n141 VSUBS 0.007638f
C176 B.n142 VSUBS 0.007638f
C177 B.n143 VSUBS 0.017121f
C178 B.n144 VSUBS 0.007638f
C179 B.n145 VSUBS 0.007638f
C180 B.n146 VSUBS 0.007638f
C181 B.n147 VSUBS 0.007638f
C182 B.n148 VSUBS 0.007638f
C183 B.n149 VSUBS 0.007638f
C184 B.n150 VSUBS 0.007638f
C185 B.n151 VSUBS 0.007638f
C186 B.n152 VSUBS 0.007638f
C187 B.n153 VSUBS 0.007638f
C188 B.n154 VSUBS 0.007638f
C189 B.n155 VSUBS 0.007638f
C190 B.n156 VSUBS 0.007638f
C191 B.n157 VSUBS 0.007638f
C192 B.n158 VSUBS 0.007638f
C193 B.n159 VSUBS 0.007638f
C194 B.n160 VSUBS 0.007638f
C195 B.n161 VSUBS 0.007638f
C196 B.n162 VSUBS 0.007638f
C197 B.n163 VSUBS 0.007638f
C198 B.n164 VSUBS 0.007638f
C199 B.n165 VSUBS 0.007638f
C200 B.n166 VSUBS 0.007638f
C201 B.n167 VSUBS 0.007638f
C202 B.n168 VSUBS 0.007638f
C203 B.n169 VSUBS 0.007638f
C204 B.n170 VSUBS 0.007638f
C205 B.t11 VSUBS 0.337168f
C206 B.t10 VSUBS 0.381725f
C207 B.t9 VSUBS 2.69081f
C208 B.n171 VSUBS 0.603378f
C209 B.n172 VSUBS 0.338491f
C210 B.n173 VSUBS 0.007638f
C211 B.n174 VSUBS 0.007638f
C212 B.n175 VSUBS 0.007638f
C213 B.n176 VSUBS 0.007638f
C214 B.n177 VSUBS 0.004268f
C215 B.n178 VSUBS 0.007638f
C216 B.n179 VSUBS 0.007638f
C217 B.n180 VSUBS 0.007638f
C218 B.n181 VSUBS 0.007638f
C219 B.n182 VSUBS 0.007638f
C220 B.n183 VSUBS 0.007638f
C221 B.n184 VSUBS 0.007638f
C222 B.n185 VSUBS 0.007638f
C223 B.n186 VSUBS 0.007638f
C224 B.n187 VSUBS 0.007638f
C225 B.n188 VSUBS 0.007638f
C226 B.n189 VSUBS 0.007638f
C227 B.n190 VSUBS 0.007638f
C228 B.n191 VSUBS 0.007638f
C229 B.n192 VSUBS 0.007638f
C230 B.n193 VSUBS 0.007638f
C231 B.n194 VSUBS 0.007638f
C232 B.n195 VSUBS 0.007638f
C233 B.n196 VSUBS 0.007638f
C234 B.n197 VSUBS 0.007638f
C235 B.n198 VSUBS 0.007638f
C236 B.n199 VSUBS 0.007638f
C237 B.n200 VSUBS 0.007638f
C238 B.n201 VSUBS 0.007638f
C239 B.n202 VSUBS 0.007638f
C240 B.n203 VSUBS 0.007638f
C241 B.n204 VSUBS 0.016922f
C242 B.n205 VSUBS 0.007638f
C243 B.n206 VSUBS 0.007638f
C244 B.n207 VSUBS 0.007638f
C245 B.n208 VSUBS 0.007638f
C246 B.n209 VSUBS 0.007638f
C247 B.n210 VSUBS 0.007638f
C248 B.n211 VSUBS 0.007638f
C249 B.n212 VSUBS 0.007638f
C250 B.n213 VSUBS 0.007638f
C251 B.n214 VSUBS 0.007638f
C252 B.n215 VSUBS 0.007638f
C253 B.n216 VSUBS 0.007638f
C254 B.n217 VSUBS 0.007638f
C255 B.n218 VSUBS 0.007638f
C256 B.n219 VSUBS 0.007638f
C257 B.n220 VSUBS 0.007638f
C258 B.n221 VSUBS 0.007638f
C259 B.n222 VSUBS 0.007638f
C260 B.n223 VSUBS 0.007638f
C261 B.n224 VSUBS 0.007638f
C262 B.n225 VSUBS 0.007638f
C263 B.n226 VSUBS 0.007638f
C264 B.n227 VSUBS 0.007638f
C265 B.n228 VSUBS 0.007638f
C266 B.n229 VSUBS 0.007638f
C267 B.n230 VSUBS 0.007638f
C268 B.n231 VSUBS 0.007638f
C269 B.n232 VSUBS 0.007638f
C270 B.n233 VSUBS 0.007638f
C271 B.n234 VSUBS 0.007638f
C272 B.n235 VSUBS 0.007638f
C273 B.n236 VSUBS 0.007638f
C274 B.n237 VSUBS 0.007638f
C275 B.n238 VSUBS 0.007638f
C276 B.n239 VSUBS 0.007638f
C277 B.n240 VSUBS 0.007638f
C278 B.n241 VSUBS 0.007638f
C279 B.n242 VSUBS 0.007638f
C280 B.n243 VSUBS 0.007638f
C281 B.n244 VSUBS 0.007638f
C282 B.n245 VSUBS 0.007638f
C283 B.n246 VSUBS 0.007638f
C284 B.n247 VSUBS 0.007638f
C285 B.n248 VSUBS 0.007638f
C286 B.n249 VSUBS 0.007638f
C287 B.n250 VSUBS 0.007638f
C288 B.n251 VSUBS 0.007638f
C289 B.n252 VSUBS 0.007638f
C290 B.n253 VSUBS 0.007638f
C291 B.n254 VSUBS 0.007638f
C292 B.n255 VSUBS 0.007638f
C293 B.n256 VSUBS 0.007638f
C294 B.n257 VSUBS 0.007638f
C295 B.n258 VSUBS 0.007638f
C296 B.n259 VSUBS 0.007638f
C297 B.n260 VSUBS 0.007638f
C298 B.n261 VSUBS 0.007638f
C299 B.n262 VSUBS 0.007638f
C300 B.n263 VSUBS 0.007638f
C301 B.n264 VSUBS 0.007638f
C302 B.n265 VSUBS 0.007638f
C303 B.n266 VSUBS 0.007638f
C304 B.n267 VSUBS 0.007638f
C305 B.n268 VSUBS 0.007638f
C306 B.n269 VSUBS 0.007638f
C307 B.n270 VSUBS 0.007638f
C308 B.n271 VSUBS 0.007638f
C309 B.n272 VSUBS 0.007638f
C310 B.n273 VSUBS 0.007638f
C311 B.n274 VSUBS 0.007638f
C312 B.n275 VSUBS 0.007638f
C313 B.n276 VSUBS 0.007638f
C314 B.n277 VSUBS 0.007638f
C315 B.n278 VSUBS 0.007638f
C316 B.n279 VSUBS 0.007638f
C317 B.n280 VSUBS 0.007638f
C318 B.n281 VSUBS 0.007638f
C319 B.n282 VSUBS 0.007638f
C320 B.n283 VSUBS 0.007638f
C321 B.n284 VSUBS 0.007638f
C322 B.n285 VSUBS 0.007638f
C323 B.n286 VSUBS 0.007638f
C324 B.n287 VSUBS 0.007638f
C325 B.n288 VSUBS 0.007638f
C326 B.n289 VSUBS 0.007638f
C327 B.n290 VSUBS 0.007638f
C328 B.n291 VSUBS 0.007638f
C329 B.n292 VSUBS 0.007638f
C330 B.n293 VSUBS 0.007638f
C331 B.n294 VSUBS 0.007638f
C332 B.n295 VSUBS 0.007638f
C333 B.n296 VSUBS 0.007638f
C334 B.n297 VSUBS 0.007638f
C335 B.n298 VSUBS 0.007638f
C336 B.n299 VSUBS 0.007638f
C337 B.n300 VSUBS 0.007638f
C338 B.n301 VSUBS 0.007638f
C339 B.n302 VSUBS 0.007638f
C340 B.n303 VSUBS 0.016101f
C341 B.n304 VSUBS 0.016101f
C342 B.n305 VSUBS 0.016922f
C343 B.n306 VSUBS 0.007638f
C344 B.n307 VSUBS 0.007638f
C345 B.n308 VSUBS 0.007638f
C346 B.n309 VSUBS 0.007638f
C347 B.n310 VSUBS 0.007638f
C348 B.n311 VSUBS 0.007638f
C349 B.n312 VSUBS 0.007638f
C350 B.n313 VSUBS 0.007638f
C351 B.n314 VSUBS 0.007638f
C352 B.n315 VSUBS 0.007638f
C353 B.n316 VSUBS 0.007638f
C354 B.n317 VSUBS 0.007638f
C355 B.n318 VSUBS 0.007638f
C356 B.n319 VSUBS 0.007638f
C357 B.n320 VSUBS 0.007638f
C358 B.n321 VSUBS 0.007638f
C359 B.n322 VSUBS 0.007638f
C360 B.n323 VSUBS 0.007638f
C361 B.n324 VSUBS 0.007638f
C362 B.n325 VSUBS 0.007638f
C363 B.n326 VSUBS 0.007638f
C364 B.n327 VSUBS 0.007638f
C365 B.n328 VSUBS 0.007638f
C366 B.n329 VSUBS 0.007638f
C367 B.n330 VSUBS 0.007638f
C368 B.n331 VSUBS 0.007638f
C369 B.n332 VSUBS 0.007638f
C370 B.n333 VSUBS 0.007638f
C371 B.n334 VSUBS 0.007638f
C372 B.n335 VSUBS 0.007638f
C373 B.n336 VSUBS 0.007638f
C374 B.n337 VSUBS 0.007638f
C375 B.n338 VSUBS 0.007638f
C376 B.n339 VSUBS 0.007638f
C377 B.n340 VSUBS 0.007638f
C378 B.n341 VSUBS 0.007638f
C379 B.n342 VSUBS 0.007638f
C380 B.n343 VSUBS 0.007638f
C381 B.n344 VSUBS 0.007638f
C382 B.n345 VSUBS 0.007638f
C383 B.n346 VSUBS 0.007638f
C384 B.n347 VSUBS 0.007638f
C385 B.n348 VSUBS 0.007638f
C386 B.n349 VSUBS 0.007638f
C387 B.n350 VSUBS 0.007638f
C388 B.n351 VSUBS 0.007638f
C389 B.n352 VSUBS 0.007638f
C390 B.n353 VSUBS 0.007638f
C391 B.n354 VSUBS 0.007638f
C392 B.n355 VSUBS 0.007638f
C393 B.n356 VSUBS 0.007638f
C394 B.n357 VSUBS 0.007638f
C395 B.n358 VSUBS 0.007638f
C396 B.n359 VSUBS 0.007638f
C397 B.n360 VSUBS 0.007638f
C398 B.n361 VSUBS 0.007638f
C399 B.n362 VSUBS 0.007638f
C400 B.n363 VSUBS 0.007638f
C401 B.n364 VSUBS 0.007638f
C402 B.n365 VSUBS 0.007638f
C403 B.n366 VSUBS 0.007638f
C404 B.n367 VSUBS 0.007638f
C405 B.n368 VSUBS 0.007638f
C406 B.n369 VSUBS 0.007638f
C407 B.n370 VSUBS 0.007638f
C408 B.n371 VSUBS 0.007638f
C409 B.n372 VSUBS 0.007638f
C410 B.n373 VSUBS 0.007638f
C411 B.n374 VSUBS 0.007638f
C412 B.n375 VSUBS 0.007638f
C413 B.n376 VSUBS 0.007638f
C414 B.n377 VSUBS 0.007638f
C415 B.n378 VSUBS 0.007638f
C416 B.n379 VSUBS 0.007638f
C417 B.n380 VSUBS 0.007638f
C418 B.n381 VSUBS 0.007638f
C419 B.n382 VSUBS 0.007638f
C420 B.n383 VSUBS 0.007638f
C421 B.t8 VSUBS 0.337164f
C422 B.t7 VSUBS 0.381722f
C423 B.t6 VSUBS 2.69081f
C424 B.n384 VSUBS 0.603381f
C425 B.n385 VSUBS 0.338495f
C426 B.n386 VSUBS 0.017696f
C427 B.n387 VSUBS 0.007189f
C428 B.n388 VSUBS 0.007638f
C429 B.n389 VSUBS 0.007638f
C430 B.n390 VSUBS 0.007638f
C431 B.n391 VSUBS 0.007638f
C432 B.n392 VSUBS 0.007638f
C433 B.n393 VSUBS 0.007638f
C434 B.n394 VSUBS 0.007638f
C435 B.n395 VSUBS 0.007638f
C436 B.n396 VSUBS 0.007638f
C437 B.n397 VSUBS 0.007638f
C438 B.n398 VSUBS 0.007638f
C439 B.n399 VSUBS 0.007638f
C440 B.n400 VSUBS 0.007638f
C441 B.n401 VSUBS 0.007638f
C442 B.n402 VSUBS 0.007638f
C443 B.n403 VSUBS 0.004268f
C444 B.n404 VSUBS 0.017696f
C445 B.n405 VSUBS 0.007189f
C446 B.n406 VSUBS 0.007638f
C447 B.n407 VSUBS 0.007638f
C448 B.n408 VSUBS 0.007638f
C449 B.n409 VSUBS 0.007638f
C450 B.n410 VSUBS 0.007638f
C451 B.n411 VSUBS 0.007638f
C452 B.n412 VSUBS 0.007638f
C453 B.n413 VSUBS 0.007638f
C454 B.n414 VSUBS 0.007638f
C455 B.n415 VSUBS 0.007638f
C456 B.n416 VSUBS 0.007638f
C457 B.n417 VSUBS 0.007638f
C458 B.n418 VSUBS 0.007638f
C459 B.n419 VSUBS 0.007638f
C460 B.n420 VSUBS 0.007638f
C461 B.n421 VSUBS 0.007638f
C462 B.n422 VSUBS 0.007638f
C463 B.n423 VSUBS 0.007638f
C464 B.n424 VSUBS 0.007638f
C465 B.n425 VSUBS 0.007638f
C466 B.n426 VSUBS 0.007638f
C467 B.n427 VSUBS 0.007638f
C468 B.n428 VSUBS 0.007638f
C469 B.n429 VSUBS 0.007638f
C470 B.n430 VSUBS 0.007638f
C471 B.n431 VSUBS 0.007638f
C472 B.n432 VSUBS 0.007638f
C473 B.n433 VSUBS 0.007638f
C474 B.n434 VSUBS 0.007638f
C475 B.n435 VSUBS 0.007638f
C476 B.n436 VSUBS 0.007638f
C477 B.n437 VSUBS 0.007638f
C478 B.n438 VSUBS 0.007638f
C479 B.n439 VSUBS 0.007638f
C480 B.n440 VSUBS 0.007638f
C481 B.n441 VSUBS 0.007638f
C482 B.n442 VSUBS 0.007638f
C483 B.n443 VSUBS 0.007638f
C484 B.n444 VSUBS 0.007638f
C485 B.n445 VSUBS 0.007638f
C486 B.n446 VSUBS 0.007638f
C487 B.n447 VSUBS 0.007638f
C488 B.n448 VSUBS 0.007638f
C489 B.n449 VSUBS 0.007638f
C490 B.n450 VSUBS 0.007638f
C491 B.n451 VSUBS 0.007638f
C492 B.n452 VSUBS 0.007638f
C493 B.n453 VSUBS 0.007638f
C494 B.n454 VSUBS 0.007638f
C495 B.n455 VSUBS 0.007638f
C496 B.n456 VSUBS 0.007638f
C497 B.n457 VSUBS 0.007638f
C498 B.n458 VSUBS 0.007638f
C499 B.n459 VSUBS 0.007638f
C500 B.n460 VSUBS 0.007638f
C501 B.n461 VSUBS 0.007638f
C502 B.n462 VSUBS 0.007638f
C503 B.n463 VSUBS 0.007638f
C504 B.n464 VSUBS 0.007638f
C505 B.n465 VSUBS 0.007638f
C506 B.n466 VSUBS 0.007638f
C507 B.n467 VSUBS 0.007638f
C508 B.n468 VSUBS 0.007638f
C509 B.n469 VSUBS 0.007638f
C510 B.n470 VSUBS 0.007638f
C511 B.n471 VSUBS 0.007638f
C512 B.n472 VSUBS 0.007638f
C513 B.n473 VSUBS 0.007638f
C514 B.n474 VSUBS 0.007638f
C515 B.n475 VSUBS 0.007638f
C516 B.n476 VSUBS 0.007638f
C517 B.n477 VSUBS 0.007638f
C518 B.n478 VSUBS 0.007638f
C519 B.n479 VSUBS 0.007638f
C520 B.n480 VSUBS 0.007638f
C521 B.n481 VSUBS 0.007638f
C522 B.n482 VSUBS 0.007638f
C523 B.n483 VSUBS 0.007638f
C524 B.n484 VSUBS 0.015902f
C525 B.n485 VSUBS 0.016922f
C526 B.n486 VSUBS 0.016101f
C527 B.n487 VSUBS 0.007638f
C528 B.n488 VSUBS 0.007638f
C529 B.n489 VSUBS 0.007638f
C530 B.n490 VSUBS 0.007638f
C531 B.n491 VSUBS 0.007638f
C532 B.n492 VSUBS 0.007638f
C533 B.n493 VSUBS 0.007638f
C534 B.n494 VSUBS 0.007638f
C535 B.n495 VSUBS 0.007638f
C536 B.n496 VSUBS 0.007638f
C537 B.n497 VSUBS 0.007638f
C538 B.n498 VSUBS 0.007638f
C539 B.n499 VSUBS 0.007638f
C540 B.n500 VSUBS 0.007638f
C541 B.n501 VSUBS 0.007638f
C542 B.n502 VSUBS 0.007638f
C543 B.n503 VSUBS 0.007638f
C544 B.n504 VSUBS 0.007638f
C545 B.n505 VSUBS 0.007638f
C546 B.n506 VSUBS 0.007638f
C547 B.n507 VSUBS 0.007638f
C548 B.n508 VSUBS 0.007638f
C549 B.n509 VSUBS 0.007638f
C550 B.n510 VSUBS 0.007638f
C551 B.n511 VSUBS 0.007638f
C552 B.n512 VSUBS 0.007638f
C553 B.n513 VSUBS 0.007638f
C554 B.n514 VSUBS 0.007638f
C555 B.n515 VSUBS 0.007638f
C556 B.n516 VSUBS 0.007638f
C557 B.n517 VSUBS 0.007638f
C558 B.n518 VSUBS 0.007638f
C559 B.n519 VSUBS 0.007638f
C560 B.n520 VSUBS 0.007638f
C561 B.n521 VSUBS 0.007638f
C562 B.n522 VSUBS 0.007638f
C563 B.n523 VSUBS 0.007638f
C564 B.n524 VSUBS 0.007638f
C565 B.n525 VSUBS 0.007638f
C566 B.n526 VSUBS 0.007638f
C567 B.n527 VSUBS 0.007638f
C568 B.n528 VSUBS 0.007638f
C569 B.n529 VSUBS 0.007638f
C570 B.n530 VSUBS 0.007638f
C571 B.n531 VSUBS 0.007638f
C572 B.n532 VSUBS 0.007638f
C573 B.n533 VSUBS 0.007638f
C574 B.n534 VSUBS 0.007638f
C575 B.n535 VSUBS 0.007638f
C576 B.n536 VSUBS 0.007638f
C577 B.n537 VSUBS 0.007638f
C578 B.n538 VSUBS 0.007638f
C579 B.n539 VSUBS 0.007638f
C580 B.n540 VSUBS 0.007638f
C581 B.n541 VSUBS 0.007638f
C582 B.n542 VSUBS 0.007638f
C583 B.n543 VSUBS 0.007638f
C584 B.n544 VSUBS 0.007638f
C585 B.n545 VSUBS 0.007638f
C586 B.n546 VSUBS 0.007638f
C587 B.n547 VSUBS 0.007638f
C588 B.n548 VSUBS 0.007638f
C589 B.n549 VSUBS 0.007638f
C590 B.n550 VSUBS 0.007638f
C591 B.n551 VSUBS 0.007638f
C592 B.n552 VSUBS 0.007638f
C593 B.n553 VSUBS 0.007638f
C594 B.n554 VSUBS 0.007638f
C595 B.n555 VSUBS 0.007638f
C596 B.n556 VSUBS 0.007638f
C597 B.n557 VSUBS 0.007638f
C598 B.n558 VSUBS 0.007638f
C599 B.n559 VSUBS 0.007638f
C600 B.n560 VSUBS 0.007638f
C601 B.n561 VSUBS 0.007638f
C602 B.n562 VSUBS 0.007638f
C603 B.n563 VSUBS 0.007638f
C604 B.n564 VSUBS 0.007638f
C605 B.n565 VSUBS 0.007638f
C606 B.n566 VSUBS 0.007638f
C607 B.n567 VSUBS 0.007638f
C608 B.n568 VSUBS 0.007638f
C609 B.n569 VSUBS 0.007638f
C610 B.n570 VSUBS 0.007638f
C611 B.n571 VSUBS 0.007638f
C612 B.n572 VSUBS 0.007638f
C613 B.n573 VSUBS 0.007638f
C614 B.n574 VSUBS 0.007638f
C615 B.n575 VSUBS 0.007638f
C616 B.n576 VSUBS 0.007638f
C617 B.n577 VSUBS 0.007638f
C618 B.n578 VSUBS 0.007638f
C619 B.n579 VSUBS 0.007638f
C620 B.n580 VSUBS 0.007638f
C621 B.n581 VSUBS 0.007638f
C622 B.n582 VSUBS 0.007638f
C623 B.n583 VSUBS 0.007638f
C624 B.n584 VSUBS 0.007638f
C625 B.n585 VSUBS 0.007638f
C626 B.n586 VSUBS 0.007638f
C627 B.n587 VSUBS 0.007638f
C628 B.n588 VSUBS 0.007638f
C629 B.n589 VSUBS 0.007638f
C630 B.n590 VSUBS 0.007638f
C631 B.n591 VSUBS 0.007638f
C632 B.n592 VSUBS 0.007638f
C633 B.n593 VSUBS 0.007638f
C634 B.n594 VSUBS 0.007638f
C635 B.n595 VSUBS 0.007638f
C636 B.n596 VSUBS 0.007638f
C637 B.n597 VSUBS 0.007638f
C638 B.n598 VSUBS 0.007638f
C639 B.n599 VSUBS 0.007638f
C640 B.n600 VSUBS 0.007638f
C641 B.n601 VSUBS 0.007638f
C642 B.n602 VSUBS 0.007638f
C643 B.n603 VSUBS 0.007638f
C644 B.n604 VSUBS 0.007638f
C645 B.n605 VSUBS 0.007638f
C646 B.n606 VSUBS 0.007638f
C647 B.n607 VSUBS 0.007638f
C648 B.n608 VSUBS 0.007638f
C649 B.n609 VSUBS 0.007638f
C650 B.n610 VSUBS 0.007638f
C651 B.n611 VSUBS 0.007638f
C652 B.n612 VSUBS 0.007638f
C653 B.n613 VSUBS 0.007638f
C654 B.n614 VSUBS 0.007638f
C655 B.n615 VSUBS 0.007638f
C656 B.n616 VSUBS 0.007638f
C657 B.n617 VSUBS 0.007638f
C658 B.n618 VSUBS 0.007638f
C659 B.n619 VSUBS 0.007638f
C660 B.n620 VSUBS 0.007638f
C661 B.n621 VSUBS 0.007638f
C662 B.n622 VSUBS 0.007638f
C663 B.n623 VSUBS 0.007638f
C664 B.n624 VSUBS 0.007638f
C665 B.n625 VSUBS 0.007638f
C666 B.n626 VSUBS 0.007638f
C667 B.n627 VSUBS 0.007638f
C668 B.n628 VSUBS 0.007638f
C669 B.n629 VSUBS 0.007638f
C670 B.n630 VSUBS 0.007638f
C671 B.n631 VSUBS 0.007638f
C672 B.n632 VSUBS 0.007638f
C673 B.n633 VSUBS 0.007638f
C674 B.n634 VSUBS 0.007638f
C675 B.n635 VSUBS 0.007638f
C676 B.n636 VSUBS 0.007638f
C677 B.n637 VSUBS 0.007638f
C678 B.n638 VSUBS 0.007638f
C679 B.n639 VSUBS 0.007638f
C680 B.n640 VSUBS 0.016101f
C681 B.n641 VSUBS 0.016101f
C682 B.n642 VSUBS 0.016922f
C683 B.n643 VSUBS 0.007638f
C684 B.n644 VSUBS 0.007638f
C685 B.n645 VSUBS 0.007638f
C686 B.n646 VSUBS 0.007638f
C687 B.n647 VSUBS 0.007638f
C688 B.n648 VSUBS 0.007638f
C689 B.n649 VSUBS 0.007638f
C690 B.n650 VSUBS 0.007638f
C691 B.n651 VSUBS 0.007638f
C692 B.n652 VSUBS 0.007638f
C693 B.n653 VSUBS 0.007638f
C694 B.n654 VSUBS 0.007638f
C695 B.n655 VSUBS 0.007638f
C696 B.n656 VSUBS 0.007638f
C697 B.n657 VSUBS 0.007638f
C698 B.n658 VSUBS 0.007638f
C699 B.n659 VSUBS 0.007638f
C700 B.n660 VSUBS 0.007638f
C701 B.n661 VSUBS 0.007638f
C702 B.n662 VSUBS 0.007638f
C703 B.n663 VSUBS 0.007638f
C704 B.n664 VSUBS 0.007638f
C705 B.n665 VSUBS 0.007638f
C706 B.n666 VSUBS 0.007638f
C707 B.n667 VSUBS 0.007638f
C708 B.n668 VSUBS 0.007638f
C709 B.n669 VSUBS 0.007638f
C710 B.n670 VSUBS 0.007638f
C711 B.n671 VSUBS 0.007638f
C712 B.n672 VSUBS 0.007638f
C713 B.n673 VSUBS 0.007638f
C714 B.n674 VSUBS 0.007638f
C715 B.n675 VSUBS 0.007638f
C716 B.n676 VSUBS 0.007638f
C717 B.n677 VSUBS 0.007638f
C718 B.n678 VSUBS 0.007638f
C719 B.n679 VSUBS 0.007638f
C720 B.n680 VSUBS 0.007638f
C721 B.n681 VSUBS 0.007638f
C722 B.n682 VSUBS 0.007638f
C723 B.n683 VSUBS 0.007638f
C724 B.n684 VSUBS 0.007638f
C725 B.n685 VSUBS 0.007638f
C726 B.n686 VSUBS 0.007638f
C727 B.n687 VSUBS 0.007638f
C728 B.n688 VSUBS 0.007638f
C729 B.n689 VSUBS 0.007638f
C730 B.n690 VSUBS 0.007638f
C731 B.n691 VSUBS 0.007638f
C732 B.n692 VSUBS 0.007638f
C733 B.n693 VSUBS 0.007638f
C734 B.n694 VSUBS 0.007638f
C735 B.n695 VSUBS 0.007638f
C736 B.n696 VSUBS 0.007638f
C737 B.n697 VSUBS 0.007638f
C738 B.n698 VSUBS 0.007638f
C739 B.n699 VSUBS 0.007638f
C740 B.n700 VSUBS 0.007638f
C741 B.n701 VSUBS 0.007638f
C742 B.n702 VSUBS 0.007638f
C743 B.n703 VSUBS 0.007638f
C744 B.n704 VSUBS 0.007638f
C745 B.n705 VSUBS 0.007638f
C746 B.n706 VSUBS 0.007638f
C747 B.n707 VSUBS 0.007638f
C748 B.n708 VSUBS 0.007638f
C749 B.n709 VSUBS 0.007638f
C750 B.n710 VSUBS 0.007638f
C751 B.n711 VSUBS 0.007638f
C752 B.n712 VSUBS 0.007638f
C753 B.n713 VSUBS 0.007638f
C754 B.n714 VSUBS 0.007638f
C755 B.n715 VSUBS 0.007638f
C756 B.n716 VSUBS 0.007638f
C757 B.n717 VSUBS 0.007638f
C758 B.n718 VSUBS 0.007638f
C759 B.n719 VSUBS 0.007638f
C760 B.n720 VSUBS 0.007638f
C761 B.n721 VSUBS 0.007638f
C762 B.n722 VSUBS 0.007189f
C763 B.n723 VSUBS 0.017696f
C764 B.n724 VSUBS 0.004268f
C765 B.n725 VSUBS 0.007638f
C766 B.n726 VSUBS 0.007638f
C767 B.n727 VSUBS 0.007638f
C768 B.n728 VSUBS 0.007638f
C769 B.n729 VSUBS 0.007638f
C770 B.n730 VSUBS 0.007638f
C771 B.n731 VSUBS 0.007638f
C772 B.n732 VSUBS 0.007638f
C773 B.n733 VSUBS 0.007638f
C774 B.n734 VSUBS 0.007638f
C775 B.n735 VSUBS 0.007638f
C776 B.n736 VSUBS 0.007638f
C777 B.n737 VSUBS 0.004268f
C778 B.n738 VSUBS 0.007638f
C779 B.n739 VSUBS 0.007638f
C780 B.n740 VSUBS 0.007638f
C781 B.n741 VSUBS 0.007638f
C782 B.n742 VSUBS 0.007638f
C783 B.n743 VSUBS 0.007638f
C784 B.n744 VSUBS 0.007638f
C785 B.n745 VSUBS 0.007638f
C786 B.n746 VSUBS 0.007638f
C787 B.n747 VSUBS 0.007638f
C788 B.n748 VSUBS 0.007638f
C789 B.n749 VSUBS 0.007638f
C790 B.n750 VSUBS 0.007638f
C791 B.n751 VSUBS 0.007638f
C792 B.n752 VSUBS 0.007638f
C793 B.n753 VSUBS 0.007638f
C794 B.n754 VSUBS 0.007638f
C795 B.n755 VSUBS 0.007638f
C796 B.n756 VSUBS 0.007638f
C797 B.n757 VSUBS 0.007638f
C798 B.n758 VSUBS 0.007638f
C799 B.n759 VSUBS 0.007638f
C800 B.n760 VSUBS 0.007638f
C801 B.n761 VSUBS 0.007638f
C802 B.n762 VSUBS 0.007638f
C803 B.n763 VSUBS 0.007638f
C804 B.n764 VSUBS 0.007638f
C805 B.n765 VSUBS 0.007638f
C806 B.n766 VSUBS 0.007638f
C807 B.n767 VSUBS 0.007638f
C808 B.n768 VSUBS 0.007638f
C809 B.n769 VSUBS 0.007638f
C810 B.n770 VSUBS 0.007638f
C811 B.n771 VSUBS 0.007638f
C812 B.n772 VSUBS 0.007638f
C813 B.n773 VSUBS 0.007638f
C814 B.n774 VSUBS 0.007638f
C815 B.n775 VSUBS 0.007638f
C816 B.n776 VSUBS 0.007638f
C817 B.n777 VSUBS 0.007638f
C818 B.n778 VSUBS 0.007638f
C819 B.n779 VSUBS 0.007638f
C820 B.n780 VSUBS 0.007638f
C821 B.n781 VSUBS 0.007638f
C822 B.n782 VSUBS 0.007638f
C823 B.n783 VSUBS 0.007638f
C824 B.n784 VSUBS 0.007638f
C825 B.n785 VSUBS 0.007638f
C826 B.n786 VSUBS 0.007638f
C827 B.n787 VSUBS 0.007638f
C828 B.n788 VSUBS 0.007638f
C829 B.n789 VSUBS 0.007638f
C830 B.n790 VSUBS 0.007638f
C831 B.n791 VSUBS 0.007638f
C832 B.n792 VSUBS 0.007638f
C833 B.n793 VSUBS 0.007638f
C834 B.n794 VSUBS 0.007638f
C835 B.n795 VSUBS 0.007638f
C836 B.n796 VSUBS 0.007638f
C837 B.n797 VSUBS 0.007638f
C838 B.n798 VSUBS 0.007638f
C839 B.n799 VSUBS 0.007638f
C840 B.n800 VSUBS 0.007638f
C841 B.n801 VSUBS 0.007638f
C842 B.n802 VSUBS 0.007638f
C843 B.n803 VSUBS 0.007638f
C844 B.n804 VSUBS 0.007638f
C845 B.n805 VSUBS 0.007638f
C846 B.n806 VSUBS 0.007638f
C847 B.n807 VSUBS 0.007638f
C848 B.n808 VSUBS 0.007638f
C849 B.n809 VSUBS 0.007638f
C850 B.n810 VSUBS 0.007638f
C851 B.n811 VSUBS 0.007638f
C852 B.n812 VSUBS 0.007638f
C853 B.n813 VSUBS 0.007638f
C854 B.n814 VSUBS 0.007638f
C855 B.n815 VSUBS 0.007638f
C856 B.n816 VSUBS 0.007638f
C857 B.n817 VSUBS 0.007638f
C858 B.n818 VSUBS 0.016922f
C859 B.n819 VSUBS 0.016922f
C860 B.n820 VSUBS 0.016101f
C861 B.n821 VSUBS 0.007638f
C862 B.n822 VSUBS 0.007638f
C863 B.n823 VSUBS 0.007638f
C864 B.n824 VSUBS 0.007638f
C865 B.n825 VSUBS 0.007638f
C866 B.n826 VSUBS 0.007638f
C867 B.n827 VSUBS 0.007638f
C868 B.n828 VSUBS 0.007638f
C869 B.n829 VSUBS 0.007638f
C870 B.n830 VSUBS 0.007638f
C871 B.n831 VSUBS 0.007638f
C872 B.n832 VSUBS 0.007638f
C873 B.n833 VSUBS 0.007638f
C874 B.n834 VSUBS 0.007638f
C875 B.n835 VSUBS 0.007638f
C876 B.n836 VSUBS 0.007638f
C877 B.n837 VSUBS 0.007638f
C878 B.n838 VSUBS 0.007638f
C879 B.n839 VSUBS 0.007638f
C880 B.n840 VSUBS 0.007638f
C881 B.n841 VSUBS 0.007638f
C882 B.n842 VSUBS 0.007638f
C883 B.n843 VSUBS 0.007638f
C884 B.n844 VSUBS 0.007638f
C885 B.n845 VSUBS 0.007638f
C886 B.n846 VSUBS 0.007638f
C887 B.n847 VSUBS 0.007638f
C888 B.n848 VSUBS 0.007638f
C889 B.n849 VSUBS 0.007638f
C890 B.n850 VSUBS 0.007638f
C891 B.n851 VSUBS 0.007638f
C892 B.n852 VSUBS 0.007638f
C893 B.n853 VSUBS 0.007638f
C894 B.n854 VSUBS 0.007638f
C895 B.n855 VSUBS 0.007638f
C896 B.n856 VSUBS 0.007638f
C897 B.n857 VSUBS 0.007638f
C898 B.n858 VSUBS 0.007638f
C899 B.n859 VSUBS 0.007638f
C900 B.n860 VSUBS 0.007638f
C901 B.n861 VSUBS 0.007638f
C902 B.n862 VSUBS 0.007638f
C903 B.n863 VSUBS 0.007638f
C904 B.n864 VSUBS 0.007638f
C905 B.n865 VSUBS 0.007638f
C906 B.n866 VSUBS 0.007638f
C907 B.n867 VSUBS 0.007638f
C908 B.n868 VSUBS 0.007638f
C909 B.n869 VSUBS 0.007638f
C910 B.n870 VSUBS 0.007638f
C911 B.n871 VSUBS 0.007638f
C912 B.n872 VSUBS 0.007638f
C913 B.n873 VSUBS 0.007638f
C914 B.n874 VSUBS 0.007638f
C915 B.n875 VSUBS 0.007638f
C916 B.n876 VSUBS 0.007638f
C917 B.n877 VSUBS 0.007638f
C918 B.n878 VSUBS 0.007638f
C919 B.n879 VSUBS 0.007638f
C920 B.n880 VSUBS 0.007638f
C921 B.n881 VSUBS 0.007638f
C922 B.n882 VSUBS 0.007638f
C923 B.n883 VSUBS 0.007638f
C924 B.n884 VSUBS 0.007638f
C925 B.n885 VSUBS 0.007638f
C926 B.n886 VSUBS 0.007638f
C927 B.n887 VSUBS 0.007638f
C928 B.n888 VSUBS 0.007638f
C929 B.n889 VSUBS 0.007638f
C930 B.n890 VSUBS 0.007638f
C931 B.n891 VSUBS 0.007638f
C932 B.n892 VSUBS 0.007638f
C933 B.n893 VSUBS 0.007638f
C934 B.n894 VSUBS 0.007638f
C935 B.n895 VSUBS 0.009967f
C936 B.n896 VSUBS 0.010618f
C937 B.n897 VSUBS 0.021114f
C938 VDD2.n0 VSUBS 0.030595f
C939 VDD2.n1 VSUBS 0.027524f
C940 VDD2.n2 VSUBS 0.01479f
C941 VDD2.n3 VSUBS 0.034959f
C942 VDD2.n4 VSUBS 0.01566f
C943 VDD2.n5 VSUBS 0.027524f
C944 VDD2.n6 VSUBS 0.015225f
C945 VDD2.n7 VSUBS 0.034959f
C946 VDD2.n8 VSUBS 0.01566f
C947 VDD2.n9 VSUBS 0.027524f
C948 VDD2.n10 VSUBS 0.01479f
C949 VDD2.n11 VSUBS 0.034959f
C950 VDD2.n12 VSUBS 0.01566f
C951 VDD2.n13 VSUBS 0.027524f
C952 VDD2.n14 VSUBS 0.01479f
C953 VDD2.n15 VSUBS 0.034959f
C954 VDD2.n16 VSUBS 0.01566f
C955 VDD2.n17 VSUBS 0.027524f
C956 VDD2.n18 VSUBS 0.01479f
C957 VDD2.n19 VSUBS 0.034959f
C958 VDD2.n20 VSUBS 0.01566f
C959 VDD2.n21 VSUBS 0.027524f
C960 VDD2.n22 VSUBS 0.01479f
C961 VDD2.n23 VSUBS 0.034959f
C962 VDD2.n24 VSUBS 0.01566f
C963 VDD2.n25 VSUBS 0.027524f
C964 VDD2.n26 VSUBS 0.01479f
C965 VDD2.n27 VSUBS 0.026219f
C966 VDD2.n28 VSUBS 0.022239f
C967 VDD2.t5 VSUBS 0.074925f
C968 VDD2.n29 VSUBS 0.20409f
C969 VDD2.n30 VSUBS 1.91243f
C970 VDD2.n31 VSUBS 0.01479f
C971 VDD2.n32 VSUBS 0.01566f
C972 VDD2.n33 VSUBS 0.034959f
C973 VDD2.n34 VSUBS 0.034959f
C974 VDD2.n35 VSUBS 0.01566f
C975 VDD2.n36 VSUBS 0.01479f
C976 VDD2.n37 VSUBS 0.027524f
C977 VDD2.n38 VSUBS 0.027524f
C978 VDD2.n39 VSUBS 0.01479f
C979 VDD2.n40 VSUBS 0.01566f
C980 VDD2.n41 VSUBS 0.034959f
C981 VDD2.n42 VSUBS 0.034959f
C982 VDD2.n43 VSUBS 0.01566f
C983 VDD2.n44 VSUBS 0.01479f
C984 VDD2.n45 VSUBS 0.027524f
C985 VDD2.n46 VSUBS 0.027524f
C986 VDD2.n47 VSUBS 0.01479f
C987 VDD2.n48 VSUBS 0.01566f
C988 VDD2.n49 VSUBS 0.034959f
C989 VDD2.n50 VSUBS 0.034959f
C990 VDD2.n51 VSUBS 0.01566f
C991 VDD2.n52 VSUBS 0.01479f
C992 VDD2.n53 VSUBS 0.027524f
C993 VDD2.n54 VSUBS 0.027524f
C994 VDD2.n55 VSUBS 0.01479f
C995 VDD2.n56 VSUBS 0.01566f
C996 VDD2.n57 VSUBS 0.034959f
C997 VDD2.n58 VSUBS 0.034959f
C998 VDD2.n59 VSUBS 0.01566f
C999 VDD2.n60 VSUBS 0.01479f
C1000 VDD2.n61 VSUBS 0.027524f
C1001 VDD2.n62 VSUBS 0.027524f
C1002 VDD2.n63 VSUBS 0.01479f
C1003 VDD2.n64 VSUBS 0.01566f
C1004 VDD2.n65 VSUBS 0.034959f
C1005 VDD2.n66 VSUBS 0.034959f
C1006 VDD2.n67 VSUBS 0.01566f
C1007 VDD2.n68 VSUBS 0.01479f
C1008 VDD2.n69 VSUBS 0.027524f
C1009 VDD2.n70 VSUBS 0.027524f
C1010 VDD2.n71 VSUBS 0.01479f
C1011 VDD2.n72 VSUBS 0.01479f
C1012 VDD2.n73 VSUBS 0.01566f
C1013 VDD2.n74 VSUBS 0.034959f
C1014 VDD2.n75 VSUBS 0.034959f
C1015 VDD2.n76 VSUBS 0.034959f
C1016 VDD2.n77 VSUBS 0.015225f
C1017 VDD2.n78 VSUBS 0.01479f
C1018 VDD2.n79 VSUBS 0.027524f
C1019 VDD2.n80 VSUBS 0.027524f
C1020 VDD2.n81 VSUBS 0.01479f
C1021 VDD2.n82 VSUBS 0.01566f
C1022 VDD2.n83 VSUBS 0.034959f
C1023 VDD2.n84 VSUBS 0.08583f
C1024 VDD2.n85 VSUBS 0.01566f
C1025 VDD2.n86 VSUBS 0.01479f
C1026 VDD2.n87 VSUBS 0.069637f
C1027 VDD2.n88 VSUBS 0.073552f
C1028 VDD2.t4 VSUBS 0.353229f
C1029 VDD2.t0 VSUBS 0.353229f
C1030 VDD2.n89 VSUBS 2.91878f
C1031 VDD2.n90 VSUBS 3.88808f
C1032 VDD2.n91 VSUBS 0.030595f
C1033 VDD2.n92 VSUBS 0.027524f
C1034 VDD2.n93 VSUBS 0.01479f
C1035 VDD2.n94 VSUBS 0.034959f
C1036 VDD2.n95 VSUBS 0.01566f
C1037 VDD2.n96 VSUBS 0.027524f
C1038 VDD2.n97 VSUBS 0.015225f
C1039 VDD2.n98 VSUBS 0.034959f
C1040 VDD2.n99 VSUBS 0.01479f
C1041 VDD2.n100 VSUBS 0.01566f
C1042 VDD2.n101 VSUBS 0.027524f
C1043 VDD2.n102 VSUBS 0.01479f
C1044 VDD2.n103 VSUBS 0.034959f
C1045 VDD2.n104 VSUBS 0.01566f
C1046 VDD2.n105 VSUBS 0.027524f
C1047 VDD2.n106 VSUBS 0.01479f
C1048 VDD2.n107 VSUBS 0.034959f
C1049 VDD2.n108 VSUBS 0.01566f
C1050 VDD2.n109 VSUBS 0.027524f
C1051 VDD2.n110 VSUBS 0.01479f
C1052 VDD2.n111 VSUBS 0.034959f
C1053 VDD2.n112 VSUBS 0.01566f
C1054 VDD2.n113 VSUBS 0.027524f
C1055 VDD2.n114 VSUBS 0.01479f
C1056 VDD2.n115 VSUBS 0.034959f
C1057 VDD2.n116 VSUBS 0.01566f
C1058 VDD2.n117 VSUBS 0.027524f
C1059 VDD2.n118 VSUBS 0.01479f
C1060 VDD2.n119 VSUBS 0.026219f
C1061 VDD2.n120 VSUBS 0.022239f
C1062 VDD2.t1 VSUBS 0.074925f
C1063 VDD2.n121 VSUBS 0.20409f
C1064 VDD2.n122 VSUBS 1.91243f
C1065 VDD2.n123 VSUBS 0.01479f
C1066 VDD2.n124 VSUBS 0.01566f
C1067 VDD2.n125 VSUBS 0.034959f
C1068 VDD2.n126 VSUBS 0.034959f
C1069 VDD2.n127 VSUBS 0.01566f
C1070 VDD2.n128 VSUBS 0.01479f
C1071 VDD2.n129 VSUBS 0.027524f
C1072 VDD2.n130 VSUBS 0.027524f
C1073 VDD2.n131 VSUBS 0.01479f
C1074 VDD2.n132 VSUBS 0.01566f
C1075 VDD2.n133 VSUBS 0.034959f
C1076 VDD2.n134 VSUBS 0.034959f
C1077 VDD2.n135 VSUBS 0.01566f
C1078 VDD2.n136 VSUBS 0.01479f
C1079 VDD2.n137 VSUBS 0.027524f
C1080 VDD2.n138 VSUBS 0.027524f
C1081 VDD2.n139 VSUBS 0.01479f
C1082 VDD2.n140 VSUBS 0.01566f
C1083 VDD2.n141 VSUBS 0.034959f
C1084 VDD2.n142 VSUBS 0.034959f
C1085 VDD2.n143 VSUBS 0.01566f
C1086 VDD2.n144 VSUBS 0.01479f
C1087 VDD2.n145 VSUBS 0.027524f
C1088 VDD2.n146 VSUBS 0.027524f
C1089 VDD2.n147 VSUBS 0.01479f
C1090 VDD2.n148 VSUBS 0.01566f
C1091 VDD2.n149 VSUBS 0.034959f
C1092 VDD2.n150 VSUBS 0.034959f
C1093 VDD2.n151 VSUBS 0.01566f
C1094 VDD2.n152 VSUBS 0.01479f
C1095 VDD2.n153 VSUBS 0.027524f
C1096 VDD2.n154 VSUBS 0.027524f
C1097 VDD2.n155 VSUBS 0.01479f
C1098 VDD2.n156 VSUBS 0.01566f
C1099 VDD2.n157 VSUBS 0.034959f
C1100 VDD2.n158 VSUBS 0.034959f
C1101 VDD2.n159 VSUBS 0.01566f
C1102 VDD2.n160 VSUBS 0.01479f
C1103 VDD2.n161 VSUBS 0.027524f
C1104 VDD2.n162 VSUBS 0.027524f
C1105 VDD2.n163 VSUBS 0.01479f
C1106 VDD2.n164 VSUBS 0.01566f
C1107 VDD2.n165 VSUBS 0.034959f
C1108 VDD2.n166 VSUBS 0.034959f
C1109 VDD2.n167 VSUBS 0.034959f
C1110 VDD2.n168 VSUBS 0.015225f
C1111 VDD2.n169 VSUBS 0.01479f
C1112 VDD2.n170 VSUBS 0.027524f
C1113 VDD2.n171 VSUBS 0.027524f
C1114 VDD2.n172 VSUBS 0.01479f
C1115 VDD2.n173 VSUBS 0.01566f
C1116 VDD2.n174 VSUBS 0.034959f
C1117 VDD2.n175 VSUBS 0.08583f
C1118 VDD2.n176 VSUBS 0.01566f
C1119 VDD2.n177 VSUBS 0.01479f
C1120 VDD2.n178 VSUBS 0.069637f
C1121 VDD2.n179 VSUBS 0.062356f
C1122 VDD2.n180 VSUBS 3.40259f
C1123 VDD2.t3 VSUBS 0.353229f
C1124 VDD2.t2 VSUBS 0.353229f
C1125 VDD2.n181 VSUBS 2.91873f
C1126 VN.t5 VSUBS 3.62211f
C1127 VN.n0 VSUBS 1.34196f
C1128 VN.n1 VSUBS 0.024327f
C1129 VN.n2 VSUBS 0.029642f
C1130 VN.n3 VSUBS 0.024327f
C1131 VN.t1 VSUBS 3.62211f
C1132 VN.n4 VSUBS 1.34977f
C1133 VN.t0 VSUBS 3.93783f
C1134 VN.n5 VSUBS 1.28288f
C1135 VN.n6 VSUBS 0.296362f
C1136 VN.n7 VSUBS 0.045113f
C1137 VN.n8 VSUBS 0.045113f
C1138 VN.n9 VSUBS 0.041085f
C1139 VN.n10 VSUBS 0.024327f
C1140 VN.n11 VSUBS 0.024327f
C1141 VN.n12 VSUBS 0.024327f
C1142 VN.n13 VSUBS 0.045113f
C1143 VN.n14 VSUBS 0.045113f
C1144 VN.n15 VSUBS 0.030414f
C1145 VN.n16 VSUBS 0.039258f
C1146 VN.n17 VSUBS 0.064743f
C1147 VN.t4 VSUBS 3.62211f
C1148 VN.n18 VSUBS 1.34196f
C1149 VN.n19 VSUBS 0.024327f
C1150 VN.n20 VSUBS 0.029642f
C1151 VN.n21 VSUBS 0.024327f
C1152 VN.t2 VSUBS 3.62211f
C1153 VN.n22 VSUBS 1.34977f
C1154 VN.t3 VSUBS 3.93783f
C1155 VN.n23 VSUBS 1.28288f
C1156 VN.n24 VSUBS 0.296362f
C1157 VN.n25 VSUBS 0.045113f
C1158 VN.n26 VSUBS 0.045113f
C1159 VN.n27 VSUBS 0.041085f
C1160 VN.n28 VSUBS 0.024327f
C1161 VN.n29 VSUBS 0.024327f
C1162 VN.n30 VSUBS 0.024327f
C1163 VN.n31 VSUBS 0.045113f
C1164 VN.n32 VSUBS 0.045113f
C1165 VN.n33 VSUBS 0.030414f
C1166 VN.n34 VSUBS 0.039258f
C1167 VN.n35 VSUBS 1.58905f
C1168 VDD1.n0 VSUBS 0.030593f
C1169 VDD1.n1 VSUBS 0.027522f
C1170 VDD1.n2 VSUBS 0.014789f
C1171 VDD1.n3 VSUBS 0.034957f
C1172 VDD1.n4 VSUBS 0.015659f
C1173 VDD1.n5 VSUBS 0.027522f
C1174 VDD1.n6 VSUBS 0.015224f
C1175 VDD1.n7 VSUBS 0.034957f
C1176 VDD1.n8 VSUBS 0.014789f
C1177 VDD1.n9 VSUBS 0.015659f
C1178 VDD1.n10 VSUBS 0.027522f
C1179 VDD1.n11 VSUBS 0.014789f
C1180 VDD1.n12 VSUBS 0.034957f
C1181 VDD1.n13 VSUBS 0.015659f
C1182 VDD1.n14 VSUBS 0.027522f
C1183 VDD1.n15 VSUBS 0.014789f
C1184 VDD1.n16 VSUBS 0.034957f
C1185 VDD1.n17 VSUBS 0.015659f
C1186 VDD1.n18 VSUBS 0.027522f
C1187 VDD1.n19 VSUBS 0.014789f
C1188 VDD1.n20 VSUBS 0.034957f
C1189 VDD1.n21 VSUBS 0.015659f
C1190 VDD1.n22 VSUBS 0.027522f
C1191 VDD1.n23 VSUBS 0.014789f
C1192 VDD1.n24 VSUBS 0.034957f
C1193 VDD1.n25 VSUBS 0.015659f
C1194 VDD1.n26 VSUBS 0.027522f
C1195 VDD1.n27 VSUBS 0.014789f
C1196 VDD1.n28 VSUBS 0.026218f
C1197 VDD1.n29 VSUBS 0.022238f
C1198 VDD1.t1 VSUBS 0.07492f
C1199 VDD1.n30 VSUBS 0.204076f
C1200 VDD1.n31 VSUBS 1.9123f
C1201 VDD1.n32 VSUBS 0.014789f
C1202 VDD1.n33 VSUBS 0.015659f
C1203 VDD1.n34 VSUBS 0.034957f
C1204 VDD1.n35 VSUBS 0.034957f
C1205 VDD1.n36 VSUBS 0.015659f
C1206 VDD1.n37 VSUBS 0.014789f
C1207 VDD1.n38 VSUBS 0.027522f
C1208 VDD1.n39 VSUBS 0.027522f
C1209 VDD1.n40 VSUBS 0.014789f
C1210 VDD1.n41 VSUBS 0.015659f
C1211 VDD1.n42 VSUBS 0.034957f
C1212 VDD1.n43 VSUBS 0.034957f
C1213 VDD1.n44 VSUBS 0.015659f
C1214 VDD1.n45 VSUBS 0.014789f
C1215 VDD1.n46 VSUBS 0.027522f
C1216 VDD1.n47 VSUBS 0.027522f
C1217 VDD1.n48 VSUBS 0.014789f
C1218 VDD1.n49 VSUBS 0.015659f
C1219 VDD1.n50 VSUBS 0.034957f
C1220 VDD1.n51 VSUBS 0.034957f
C1221 VDD1.n52 VSUBS 0.015659f
C1222 VDD1.n53 VSUBS 0.014789f
C1223 VDD1.n54 VSUBS 0.027522f
C1224 VDD1.n55 VSUBS 0.027522f
C1225 VDD1.n56 VSUBS 0.014789f
C1226 VDD1.n57 VSUBS 0.015659f
C1227 VDD1.n58 VSUBS 0.034957f
C1228 VDD1.n59 VSUBS 0.034957f
C1229 VDD1.n60 VSUBS 0.015659f
C1230 VDD1.n61 VSUBS 0.014789f
C1231 VDD1.n62 VSUBS 0.027522f
C1232 VDD1.n63 VSUBS 0.027522f
C1233 VDD1.n64 VSUBS 0.014789f
C1234 VDD1.n65 VSUBS 0.015659f
C1235 VDD1.n66 VSUBS 0.034957f
C1236 VDD1.n67 VSUBS 0.034957f
C1237 VDD1.n68 VSUBS 0.015659f
C1238 VDD1.n69 VSUBS 0.014789f
C1239 VDD1.n70 VSUBS 0.027522f
C1240 VDD1.n71 VSUBS 0.027522f
C1241 VDD1.n72 VSUBS 0.014789f
C1242 VDD1.n73 VSUBS 0.015659f
C1243 VDD1.n74 VSUBS 0.034957f
C1244 VDD1.n75 VSUBS 0.034957f
C1245 VDD1.n76 VSUBS 0.034957f
C1246 VDD1.n77 VSUBS 0.015224f
C1247 VDD1.n78 VSUBS 0.014789f
C1248 VDD1.n79 VSUBS 0.027522f
C1249 VDD1.n80 VSUBS 0.027522f
C1250 VDD1.n81 VSUBS 0.014789f
C1251 VDD1.n82 VSUBS 0.015659f
C1252 VDD1.n83 VSUBS 0.034957f
C1253 VDD1.n84 VSUBS 0.085824f
C1254 VDD1.n85 VSUBS 0.015659f
C1255 VDD1.n86 VSUBS 0.014789f
C1256 VDD1.n87 VSUBS 0.069633f
C1257 VDD1.n88 VSUBS 0.074509f
C1258 VDD1.n89 VSUBS 0.030593f
C1259 VDD1.n90 VSUBS 0.027522f
C1260 VDD1.n91 VSUBS 0.014789f
C1261 VDD1.n92 VSUBS 0.034957f
C1262 VDD1.n93 VSUBS 0.015659f
C1263 VDD1.n94 VSUBS 0.027522f
C1264 VDD1.n95 VSUBS 0.015224f
C1265 VDD1.n96 VSUBS 0.034957f
C1266 VDD1.n97 VSUBS 0.015659f
C1267 VDD1.n98 VSUBS 0.027522f
C1268 VDD1.n99 VSUBS 0.014789f
C1269 VDD1.n100 VSUBS 0.034957f
C1270 VDD1.n101 VSUBS 0.015659f
C1271 VDD1.n102 VSUBS 0.027522f
C1272 VDD1.n103 VSUBS 0.014789f
C1273 VDD1.n104 VSUBS 0.034957f
C1274 VDD1.n105 VSUBS 0.015659f
C1275 VDD1.n106 VSUBS 0.027522f
C1276 VDD1.n107 VSUBS 0.014789f
C1277 VDD1.n108 VSUBS 0.034957f
C1278 VDD1.n109 VSUBS 0.015659f
C1279 VDD1.n110 VSUBS 0.027522f
C1280 VDD1.n111 VSUBS 0.014789f
C1281 VDD1.n112 VSUBS 0.034957f
C1282 VDD1.n113 VSUBS 0.015659f
C1283 VDD1.n114 VSUBS 0.027522f
C1284 VDD1.n115 VSUBS 0.014789f
C1285 VDD1.n116 VSUBS 0.026218f
C1286 VDD1.n117 VSUBS 0.022238f
C1287 VDD1.t2 VSUBS 0.07492f
C1288 VDD1.n118 VSUBS 0.204076f
C1289 VDD1.n119 VSUBS 1.9123f
C1290 VDD1.n120 VSUBS 0.014789f
C1291 VDD1.n121 VSUBS 0.015659f
C1292 VDD1.n122 VSUBS 0.034957f
C1293 VDD1.n123 VSUBS 0.034957f
C1294 VDD1.n124 VSUBS 0.015659f
C1295 VDD1.n125 VSUBS 0.014789f
C1296 VDD1.n126 VSUBS 0.027522f
C1297 VDD1.n127 VSUBS 0.027522f
C1298 VDD1.n128 VSUBS 0.014789f
C1299 VDD1.n129 VSUBS 0.015659f
C1300 VDD1.n130 VSUBS 0.034957f
C1301 VDD1.n131 VSUBS 0.034957f
C1302 VDD1.n132 VSUBS 0.015659f
C1303 VDD1.n133 VSUBS 0.014789f
C1304 VDD1.n134 VSUBS 0.027522f
C1305 VDD1.n135 VSUBS 0.027522f
C1306 VDD1.n136 VSUBS 0.014789f
C1307 VDD1.n137 VSUBS 0.015659f
C1308 VDD1.n138 VSUBS 0.034957f
C1309 VDD1.n139 VSUBS 0.034957f
C1310 VDD1.n140 VSUBS 0.015659f
C1311 VDD1.n141 VSUBS 0.014789f
C1312 VDD1.n142 VSUBS 0.027522f
C1313 VDD1.n143 VSUBS 0.027522f
C1314 VDD1.n144 VSUBS 0.014789f
C1315 VDD1.n145 VSUBS 0.015659f
C1316 VDD1.n146 VSUBS 0.034957f
C1317 VDD1.n147 VSUBS 0.034957f
C1318 VDD1.n148 VSUBS 0.015659f
C1319 VDD1.n149 VSUBS 0.014789f
C1320 VDD1.n150 VSUBS 0.027522f
C1321 VDD1.n151 VSUBS 0.027522f
C1322 VDD1.n152 VSUBS 0.014789f
C1323 VDD1.n153 VSUBS 0.015659f
C1324 VDD1.n154 VSUBS 0.034957f
C1325 VDD1.n155 VSUBS 0.034957f
C1326 VDD1.n156 VSUBS 0.015659f
C1327 VDD1.n157 VSUBS 0.014789f
C1328 VDD1.n158 VSUBS 0.027522f
C1329 VDD1.n159 VSUBS 0.027522f
C1330 VDD1.n160 VSUBS 0.014789f
C1331 VDD1.n161 VSUBS 0.014789f
C1332 VDD1.n162 VSUBS 0.015659f
C1333 VDD1.n163 VSUBS 0.034957f
C1334 VDD1.n164 VSUBS 0.034957f
C1335 VDD1.n165 VSUBS 0.034957f
C1336 VDD1.n166 VSUBS 0.015224f
C1337 VDD1.n167 VSUBS 0.014789f
C1338 VDD1.n168 VSUBS 0.027522f
C1339 VDD1.n169 VSUBS 0.027522f
C1340 VDD1.n170 VSUBS 0.014789f
C1341 VDD1.n171 VSUBS 0.015659f
C1342 VDD1.n172 VSUBS 0.034957f
C1343 VDD1.n173 VSUBS 0.085824f
C1344 VDD1.n174 VSUBS 0.015659f
C1345 VDD1.n175 VSUBS 0.014789f
C1346 VDD1.n176 VSUBS 0.069633f
C1347 VDD1.n177 VSUBS 0.073547f
C1348 VDD1.t4 VSUBS 0.353205f
C1349 VDD1.t0 VSUBS 0.353205f
C1350 VDD1.n178 VSUBS 2.91858f
C1351 VDD1.n179 VSUBS 4.04976f
C1352 VDD1.t3 VSUBS 0.353205f
C1353 VDD1.t5 VSUBS 0.353205f
C1354 VDD1.n180 VSUBS 2.9098f
C1355 VDD1.n181 VSUBS 3.94771f
C1356 VTAIL.t11 VSUBS 0.364649f
C1357 VTAIL.t0 VSUBS 0.364649f
C1358 VTAIL.n0 VSUBS 2.84612f
C1359 VTAIL.n1 VSUBS 0.922848f
C1360 VTAIL.n2 VSUBS 0.031584f
C1361 VTAIL.n3 VSUBS 0.028414f
C1362 VTAIL.n4 VSUBS 0.015269f
C1363 VTAIL.n5 VSUBS 0.036089f
C1364 VTAIL.n6 VSUBS 0.016167f
C1365 VTAIL.n7 VSUBS 0.028414f
C1366 VTAIL.n8 VSUBS 0.015718f
C1367 VTAIL.n9 VSUBS 0.036089f
C1368 VTAIL.n10 VSUBS 0.016167f
C1369 VTAIL.n11 VSUBS 0.028414f
C1370 VTAIL.n12 VSUBS 0.015269f
C1371 VTAIL.n13 VSUBS 0.036089f
C1372 VTAIL.n14 VSUBS 0.016167f
C1373 VTAIL.n15 VSUBS 0.028414f
C1374 VTAIL.n16 VSUBS 0.015269f
C1375 VTAIL.n17 VSUBS 0.036089f
C1376 VTAIL.n18 VSUBS 0.016167f
C1377 VTAIL.n19 VSUBS 0.028414f
C1378 VTAIL.n20 VSUBS 0.015269f
C1379 VTAIL.n21 VSUBS 0.036089f
C1380 VTAIL.n22 VSUBS 0.016167f
C1381 VTAIL.n23 VSUBS 0.028414f
C1382 VTAIL.n24 VSUBS 0.015269f
C1383 VTAIL.n25 VSUBS 0.036089f
C1384 VTAIL.n26 VSUBS 0.016167f
C1385 VTAIL.n27 VSUBS 0.028414f
C1386 VTAIL.n28 VSUBS 0.015269f
C1387 VTAIL.n29 VSUBS 0.027067f
C1388 VTAIL.n30 VSUBS 0.022958f
C1389 VTAIL.t7 VSUBS 0.077348f
C1390 VTAIL.n31 VSUBS 0.210688f
C1391 VTAIL.n32 VSUBS 1.97426f
C1392 VTAIL.n33 VSUBS 0.015269f
C1393 VTAIL.n34 VSUBS 0.016167f
C1394 VTAIL.n35 VSUBS 0.036089f
C1395 VTAIL.n36 VSUBS 0.036089f
C1396 VTAIL.n37 VSUBS 0.016167f
C1397 VTAIL.n38 VSUBS 0.015269f
C1398 VTAIL.n39 VSUBS 0.028414f
C1399 VTAIL.n40 VSUBS 0.028414f
C1400 VTAIL.n41 VSUBS 0.015269f
C1401 VTAIL.n42 VSUBS 0.016167f
C1402 VTAIL.n43 VSUBS 0.036089f
C1403 VTAIL.n44 VSUBS 0.036089f
C1404 VTAIL.n45 VSUBS 0.016167f
C1405 VTAIL.n46 VSUBS 0.015269f
C1406 VTAIL.n47 VSUBS 0.028414f
C1407 VTAIL.n48 VSUBS 0.028414f
C1408 VTAIL.n49 VSUBS 0.015269f
C1409 VTAIL.n50 VSUBS 0.016167f
C1410 VTAIL.n51 VSUBS 0.036089f
C1411 VTAIL.n52 VSUBS 0.036089f
C1412 VTAIL.n53 VSUBS 0.016167f
C1413 VTAIL.n54 VSUBS 0.015269f
C1414 VTAIL.n55 VSUBS 0.028414f
C1415 VTAIL.n56 VSUBS 0.028414f
C1416 VTAIL.n57 VSUBS 0.015269f
C1417 VTAIL.n58 VSUBS 0.016167f
C1418 VTAIL.n59 VSUBS 0.036089f
C1419 VTAIL.n60 VSUBS 0.036089f
C1420 VTAIL.n61 VSUBS 0.016167f
C1421 VTAIL.n62 VSUBS 0.015269f
C1422 VTAIL.n63 VSUBS 0.028414f
C1423 VTAIL.n64 VSUBS 0.028414f
C1424 VTAIL.n65 VSUBS 0.015269f
C1425 VTAIL.n66 VSUBS 0.016167f
C1426 VTAIL.n67 VSUBS 0.036089f
C1427 VTAIL.n68 VSUBS 0.036089f
C1428 VTAIL.n69 VSUBS 0.016167f
C1429 VTAIL.n70 VSUBS 0.015269f
C1430 VTAIL.n71 VSUBS 0.028414f
C1431 VTAIL.n72 VSUBS 0.028414f
C1432 VTAIL.n73 VSUBS 0.015269f
C1433 VTAIL.n74 VSUBS 0.015269f
C1434 VTAIL.n75 VSUBS 0.016167f
C1435 VTAIL.n76 VSUBS 0.036089f
C1436 VTAIL.n77 VSUBS 0.036089f
C1437 VTAIL.n78 VSUBS 0.036089f
C1438 VTAIL.n79 VSUBS 0.015718f
C1439 VTAIL.n80 VSUBS 0.015269f
C1440 VTAIL.n81 VSUBS 0.028414f
C1441 VTAIL.n82 VSUBS 0.028414f
C1442 VTAIL.n83 VSUBS 0.015269f
C1443 VTAIL.n84 VSUBS 0.016167f
C1444 VTAIL.n85 VSUBS 0.036089f
C1445 VTAIL.n86 VSUBS 0.088605f
C1446 VTAIL.n87 VSUBS 0.016167f
C1447 VTAIL.n88 VSUBS 0.015269f
C1448 VTAIL.n89 VSUBS 0.071889f
C1449 VTAIL.n90 VSUBS 0.044797f
C1450 VTAIL.n91 VSUBS 0.505298f
C1451 VTAIL.t6 VSUBS 0.364649f
C1452 VTAIL.t5 VSUBS 0.364649f
C1453 VTAIL.n92 VSUBS 2.84612f
C1454 VTAIL.n93 VSUBS 3.19403f
C1455 VTAIL.t4 VSUBS 0.364649f
C1456 VTAIL.t3 VSUBS 0.364649f
C1457 VTAIL.n94 VSUBS 2.84614f
C1458 VTAIL.n95 VSUBS 3.19401f
C1459 VTAIL.n96 VSUBS 0.031584f
C1460 VTAIL.n97 VSUBS 0.028414f
C1461 VTAIL.n98 VSUBS 0.015269f
C1462 VTAIL.n99 VSUBS 0.036089f
C1463 VTAIL.n100 VSUBS 0.016167f
C1464 VTAIL.n101 VSUBS 0.028414f
C1465 VTAIL.n102 VSUBS 0.015718f
C1466 VTAIL.n103 VSUBS 0.036089f
C1467 VTAIL.n104 VSUBS 0.015269f
C1468 VTAIL.n105 VSUBS 0.016167f
C1469 VTAIL.n106 VSUBS 0.028414f
C1470 VTAIL.n107 VSUBS 0.015269f
C1471 VTAIL.n108 VSUBS 0.036089f
C1472 VTAIL.n109 VSUBS 0.016167f
C1473 VTAIL.n110 VSUBS 0.028414f
C1474 VTAIL.n111 VSUBS 0.015269f
C1475 VTAIL.n112 VSUBS 0.036089f
C1476 VTAIL.n113 VSUBS 0.016167f
C1477 VTAIL.n114 VSUBS 0.028414f
C1478 VTAIL.n115 VSUBS 0.015269f
C1479 VTAIL.n116 VSUBS 0.036089f
C1480 VTAIL.n117 VSUBS 0.016167f
C1481 VTAIL.n118 VSUBS 0.028414f
C1482 VTAIL.n119 VSUBS 0.015269f
C1483 VTAIL.n120 VSUBS 0.036089f
C1484 VTAIL.n121 VSUBS 0.016167f
C1485 VTAIL.n122 VSUBS 0.028414f
C1486 VTAIL.n123 VSUBS 0.015269f
C1487 VTAIL.n124 VSUBS 0.027067f
C1488 VTAIL.n125 VSUBS 0.022958f
C1489 VTAIL.t1 VSUBS 0.077348f
C1490 VTAIL.n126 VSUBS 0.210688f
C1491 VTAIL.n127 VSUBS 1.97426f
C1492 VTAIL.n128 VSUBS 0.015269f
C1493 VTAIL.n129 VSUBS 0.016167f
C1494 VTAIL.n130 VSUBS 0.036089f
C1495 VTAIL.n131 VSUBS 0.036089f
C1496 VTAIL.n132 VSUBS 0.016167f
C1497 VTAIL.n133 VSUBS 0.015269f
C1498 VTAIL.n134 VSUBS 0.028414f
C1499 VTAIL.n135 VSUBS 0.028414f
C1500 VTAIL.n136 VSUBS 0.015269f
C1501 VTAIL.n137 VSUBS 0.016167f
C1502 VTAIL.n138 VSUBS 0.036089f
C1503 VTAIL.n139 VSUBS 0.036089f
C1504 VTAIL.n140 VSUBS 0.016167f
C1505 VTAIL.n141 VSUBS 0.015269f
C1506 VTAIL.n142 VSUBS 0.028414f
C1507 VTAIL.n143 VSUBS 0.028414f
C1508 VTAIL.n144 VSUBS 0.015269f
C1509 VTAIL.n145 VSUBS 0.016167f
C1510 VTAIL.n146 VSUBS 0.036089f
C1511 VTAIL.n147 VSUBS 0.036089f
C1512 VTAIL.n148 VSUBS 0.016167f
C1513 VTAIL.n149 VSUBS 0.015269f
C1514 VTAIL.n150 VSUBS 0.028414f
C1515 VTAIL.n151 VSUBS 0.028414f
C1516 VTAIL.n152 VSUBS 0.015269f
C1517 VTAIL.n153 VSUBS 0.016167f
C1518 VTAIL.n154 VSUBS 0.036089f
C1519 VTAIL.n155 VSUBS 0.036089f
C1520 VTAIL.n156 VSUBS 0.016167f
C1521 VTAIL.n157 VSUBS 0.015269f
C1522 VTAIL.n158 VSUBS 0.028414f
C1523 VTAIL.n159 VSUBS 0.028414f
C1524 VTAIL.n160 VSUBS 0.015269f
C1525 VTAIL.n161 VSUBS 0.016167f
C1526 VTAIL.n162 VSUBS 0.036089f
C1527 VTAIL.n163 VSUBS 0.036089f
C1528 VTAIL.n164 VSUBS 0.016167f
C1529 VTAIL.n165 VSUBS 0.015269f
C1530 VTAIL.n166 VSUBS 0.028414f
C1531 VTAIL.n167 VSUBS 0.028414f
C1532 VTAIL.n168 VSUBS 0.015269f
C1533 VTAIL.n169 VSUBS 0.016167f
C1534 VTAIL.n170 VSUBS 0.036089f
C1535 VTAIL.n171 VSUBS 0.036089f
C1536 VTAIL.n172 VSUBS 0.036089f
C1537 VTAIL.n173 VSUBS 0.015718f
C1538 VTAIL.n174 VSUBS 0.015269f
C1539 VTAIL.n175 VSUBS 0.028414f
C1540 VTAIL.n176 VSUBS 0.028414f
C1541 VTAIL.n177 VSUBS 0.015269f
C1542 VTAIL.n178 VSUBS 0.016167f
C1543 VTAIL.n179 VSUBS 0.036089f
C1544 VTAIL.n180 VSUBS 0.088605f
C1545 VTAIL.n181 VSUBS 0.016167f
C1546 VTAIL.n182 VSUBS 0.015269f
C1547 VTAIL.n183 VSUBS 0.071889f
C1548 VTAIL.n184 VSUBS 0.044797f
C1549 VTAIL.n185 VSUBS 0.505298f
C1550 VTAIL.t10 VSUBS 0.364649f
C1551 VTAIL.t9 VSUBS 0.364649f
C1552 VTAIL.n186 VSUBS 2.84614f
C1553 VTAIL.n187 VSUBS 1.13475f
C1554 VTAIL.n188 VSUBS 0.031584f
C1555 VTAIL.n189 VSUBS 0.028414f
C1556 VTAIL.n190 VSUBS 0.015269f
C1557 VTAIL.n191 VSUBS 0.036089f
C1558 VTAIL.n192 VSUBS 0.016167f
C1559 VTAIL.n193 VSUBS 0.028414f
C1560 VTAIL.n194 VSUBS 0.015718f
C1561 VTAIL.n195 VSUBS 0.036089f
C1562 VTAIL.n196 VSUBS 0.015269f
C1563 VTAIL.n197 VSUBS 0.016167f
C1564 VTAIL.n198 VSUBS 0.028414f
C1565 VTAIL.n199 VSUBS 0.015269f
C1566 VTAIL.n200 VSUBS 0.036089f
C1567 VTAIL.n201 VSUBS 0.016167f
C1568 VTAIL.n202 VSUBS 0.028414f
C1569 VTAIL.n203 VSUBS 0.015269f
C1570 VTAIL.n204 VSUBS 0.036089f
C1571 VTAIL.n205 VSUBS 0.016167f
C1572 VTAIL.n206 VSUBS 0.028414f
C1573 VTAIL.n207 VSUBS 0.015269f
C1574 VTAIL.n208 VSUBS 0.036089f
C1575 VTAIL.n209 VSUBS 0.016167f
C1576 VTAIL.n210 VSUBS 0.028414f
C1577 VTAIL.n211 VSUBS 0.015269f
C1578 VTAIL.n212 VSUBS 0.036089f
C1579 VTAIL.n213 VSUBS 0.016167f
C1580 VTAIL.n214 VSUBS 0.028414f
C1581 VTAIL.n215 VSUBS 0.015269f
C1582 VTAIL.n216 VSUBS 0.027067f
C1583 VTAIL.n217 VSUBS 0.022958f
C1584 VTAIL.t8 VSUBS 0.077348f
C1585 VTAIL.n218 VSUBS 0.210688f
C1586 VTAIL.n219 VSUBS 1.97426f
C1587 VTAIL.n220 VSUBS 0.015269f
C1588 VTAIL.n221 VSUBS 0.016167f
C1589 VTAIL.n222 VSUBS 0.036089f
C1590 VTAIL.n223 VSUBS 0.036089f
C1591 VTAIL.n224 VSUBS 0.016167f
C1592 VTAIL.n225 VSUBS 0.015269f
C1593 VTAIL.n226 VSUBS 0.028414f
C1594 VTAIL.n227 VSUBS 0.028414f
C1595 VTAIL.n228 VSUBS 0.015269f
C1596 VTAIL.n229 VSUBS 0.016167f
C1597 VTAIL.n230 VSUBS 0.036089f
C1598 VTAIL.n231 VSUBS 0.036089f
C1599 VTAIL.n232 VSUBS 0.016167f
C1600 VTAIL.n233 VSUBS 0.015269f
C1601 VTAIL.n234 VSUBS 0.028414f
C1602 VTAIL.n235 VSUBS 0.028414f
C1603 VTAIL.n236 VSUBS 0.015269f
C1604 VTAIL.n237 VSUBS 0.016167f
C1605 VTAIL.n238 VSUBS 0.036089f
C1606 VTAIL.n239 VSUBS 0.036089f
C1607 VTAIL.n240 VSUBS 0.016167f
C1608 VTAIL.n241 VSUBS 0.015269f
C1609 VTAIL.n242 VSUBS 0.028414f
C1610 VTAIL.n243 VSUBS 0.028414f
C1611 VTAIL.n244 VSUBS 0.015269f
C1612 VTAIL.n245 VSUBS 0.016167f
C1613 VTAIL.n246 VSUBS 0.036089f
C1614 VTAIL.n247 VSUBS 0.036089f
C1615 VTAIL.n248 VSUBS 0.016167f
C1616 VTAIL.n249 VSUBS 0.015269f
C1617 VTAIL.n250 VSUBS 0.028414f
C1618 VTAIL.n251 VSUBS 0.028414f
C1619 VTAIL.n252 VSUBS 0.015269f
C1620 VTAIL.n253 VSUBS 0.016167f
C1621 VTAIL.n254 VSUBS 0.036089f
C1622 VTAIL.n255 VSUBS 0.036089f
C1623 VTAIL.n256 VSUBS 0.016167f
C1624 VTAIL.n257 VSUBS 0.015269f
C1625 VTAIL.n258 VSUBS 0.028414f
C1626 VTAIL.n259 VSUBS 0.028414f
C1627 VTAIL.n260 VSUBS 0.015269f
C1628 VTAIL.n261 VSUBS 0.016167f
C1629 VTAIL.n262 VSUBS 0.036089f
C1630 VTAIL.n263 VSUBS 0.036089f
C1631 VTAIL.n264 VSUBS 0.036089f
C1632 VTAIL.n265 VSUBS 0.015718f
C1633 VTAIL.n266 VSUBS 0.015269f
C1634 VTAIL.n267 VSUBS 0.028414f
C1635 VTAIL.n268 VSUBS 0.028414f
C1636 VTAIL.n269 VSUBS 0.015269f
C1637 VTAIL.n270 VSUBS 0.016167f
C1638 VTAIL.n271 VSUBS 0.036089f
C1639 VTAIL.n272 VSUBS 0.088605f
C1640 VTAIL.n273 VSUBS 0.016167f
C1641 VTAIL.n274 VSUBS 0.015269f
C1642 VTAIL.n275 VSUBS 0.071889f
C1643 VTAIL.n276 VSUBS 0.044797f
C1644 VTAIL.n277 VSUBS 2.27489f
C1645 VTAIL.n278 VSUBS 0.031584f
C1646 VTAIL.n279 VSUBS 0.028414f
C1647 VTAIL.n280 VSUBS 0.015269f
C1648 VTAIL.n281 VSUBS 0.036089f
C1649 VTAIL.n282 VSUBS 0.016167f
C1650 VTAIL.n283 VSUBS 0.028414f
C1651 VTAIL.n284 VSUBS 0.015718f
C1652 VTAIL.n285 VSUBS 0.036089f
C1653 VTAIL.n286 VSUBS 0.016167f
C1654 VTAIL.n287 VSUBS 0.028414f
C1655 VTAIL.n288 VSUBS 0.015269f
C1656 VTAIL.n289 VSUBS 0.036089f
C1657 VTAIL.n290 VSUBS 0.016167f
C1658 VTAIL.n291 VSUBS 0.028414f
C1659 VTAIL.n292 VSUBS 0.015269f
C1660 VTAIL.n293 VSUBS 0.036089f
C1661 VTAIL.n294 VSUBS 0.016167f
C1662 VTAIL.n295 VSUBS 0.028414f
C1663 VTAIL.n296 VSUBS 0.015269f
C1664 VTAIL.n297 VSUBS 0.036089f
C1665 VTAIL.n298 VSUBS 0.016167f
C1666 VTAIL.n299 VSUBS 0.028414f
C1667 VTAIL.n300 VSUBS 0.015269f
C1668 VTAIL.n301 VSUBS 0.036089f
C1669 VTAIL.n302 VSUBS 0.016167f
C1670 VTAIL.n303 VSUBS 0.028414f
C1671 VTAIL.n304 VSUBS 0.015269f
C1672 VTAIL.n305 VSUBS 0.027067f
C1673 VTAIL.n306 VSUBS 0.022958f
C1674 VTAIL.t2 VSUBS 0.077348f
C1675 VTAIL.n307 VSUBS 0.210688f
C1676 VTAIL.n308 VSUBS 1.97426f
C1677 VTAIL.n309 VSUBS 0.015269f
C1678 VTAIL.n310 VSUBS 0.016167f
C1679 VTAIL.n311 VSUBS 0.036089f
C1680 VTAIL.n312 VSUBS 0.036089f
C1681 VTAIL.n313 VSUBS 0.016167f
C1682 VTAIL.n314 VSUBS 0.015269f
C1683 VTAIL.n315 VSUBS 0.028414f
C1684 VTAIL.n316 VSUBS 0.028414f
C1685 VTAIL.n317 VSUBS 0.015269f
C1686 VTAIL.n318 VSUBS 0.016167f
C1687 VTAIL.n319 VSUBS 0.036089f
C1688 VTAIL.n320 VSUBS 0.036089f
C1689 VTAIL.n321 VSUBS 0.016167f
C1690 VTAIL.n322 VSUBS 0.015269f
C1691 VTAIL.n323 VSUBS 0.028414f
C1692 VTAIL.n324 VSUBS 0.028414f
C1693 VTAIL.n325 VSUBS 0.015269f
C1694 VTAIL.n326 VSUBS 0.016167f
C1695 VTAIL.n327 VSUBS 0.036089f
C1696 VTAIL.n328 VSUBS 0.036089f
C1697 VTAIL.n329 VSUBS 0.016167f
C1698 VTAIL.n330 VSUBS 0.015269f
C1699 VTAIL.n331 VSUBS 0.028414f
C1700 VTAIL.n332 VSUBS 0.028414f
C1701 VTAIL.n333 VSUBS 0.015269f
C1702 VTAIL.n334 VSUBS 0.016167f
C1703 VTAIL.n335 VSUBS 0.036089f
C1704 VTAIL.n336 VSUBS 0.036089f
C1705 VTAIL.n337 VSUBS 0.016167f
C1706 VTAIL.n338 VSUBS 0.015269f
C1707 VTAIL.n339 VSUBS 0.028414f
C1708 VTAIL.n340 VSUBS 0.028414f
C1709 VTAIL.n341 VSUBS 0.015269f
C1710 VTAIL.n342 VSUBS 0.016167f
C1711 VTAIL.n343 VSUBS 0.036089f
C1712 VTAIL.n344 VSUBS 0.036089f
C1713 VTAIL.n345 VSUBS 0.016167f
C1714 VTAIL.n346 VSUBS 0.015269f
C1715 VTAIL.n347 VSUBS 0.028414f
C1716 VTAIL.n348 VSUBS 0.028414f
C1717 VTAIL.n349 VSUBS 0.015269f
C1718 VTAIL.n350 VSUBS 0.015269f
C1719 VTAIL.n351 VSUBS 0.016167f
C1720 VTAIL.n352 VSUBS 0.036089f
C1721 VTAIL.n353 VSUBS 0.036089f
C1722 VTAIL.n354 VSUBS 0.036089f
C1723 VTAIL.n355 VSUBS 0.015718f
C1724 VTAIL.n356 VSUBS 0.015269f
C1725 VTAIL.n357 VSUBS 0.028414f
C1726 VTAIL.n358 VSUBS 0.028414f
C1727 VTAIL.n359 VSUBS 0.015269f
C1728 VTAIL.n360 VSUBS 0.016167f
C1729 VTAIL.n361 VSUBS 0.036089f
C1730 VTAIL.n362 VSUBS 0.088605f
C1731 VTAIL.n363 VSUBS 0.016167f
C1732 VTAIL.n364 VSUBS 0.015269f
C1733 VTAIL.n365 VSUBS 0.071889f
C1734 VTAIL.n366 VSUBS 0.044797f
C1735 VTAIL.n367 VSUBS 2.19714f
C1736 VP.t5 VSUBS 3.93642f
C1737 VP.n0 VSUBS 1.45841f
C1738 VP.n1 VSUBS 0.026438f
C1739 VP.n2 VSUBS 0.032215f
C1740 VP.n3 VSUBS 0.026438f
C1741 VP.t1 VSUBS 3.93642f
C1742 VP.n4 VSUBS 1.38866f
C1743 VP.n5 VSUBS 0.026438f
C1744 VP.n6 VSUBS 0.032215f
C1745 VP.n7 VSUBS 0.026438f
C1746 VP.t3 VSUBS 3.93642f
C1747 VP.n8 VSUBS 1.45841f
C1748 VP.t0 VSUBS 3.93642f
C1749 VP.n9 VSUBS 1.45841f
C1750 VP.n10 VSUBS 0.026438f
C1751 VP.n11 VSUBS 0.032215f
C1752 VP.n12 VSUBS 0.026438f
C1753 VP.t2 VSUBS 3.93642f
C1754 VP.n13 VSUBS 1.4669f
C1755 VP.t4 VSUBS 4.27954f
C1756 VP.n14 VSUBS 1.3942f
C1757 VP.n15 VSUBS 0.322079f
C1758 VP.n16 VSUBS 0.049028f
C1759 VP.n17 VSUBS 0.049028f
C1760 VP.n18 VSUBS 0.04465f
C1761 VP.n19 VSUBS 0.026438f
C1762 VP.n20 VSUBS 0.026438f
C1763 VP.n21 VSUBS 0.026438f
C1764 VP.n22 VSUBS 0.049028f
C1765 VP.n23 VSUBS 0.049028f
C1766 VP.n24 VSUBS 0.033053f
C1767 VP.n25 VSUBS 0.042664f
C1768 VP.n26 VSUBS 1.71645f
C1769 VP.n27 VSUBS 1.73384f
C1770 VP.n28 VSUBS 0.042664f
C1771 VP.n29 VSUBS 0.033053f
C1772 VP.n30 VSUBS 0.049028f
C1773 VP.n31 VSUBS 0.049028f
C1774 VP.n32 VSUBS 0.026438f
C1775 VP.n33 VSUBS 0.026438f
C1776 VP.n34 VSUBS 0.026438f
C1777 VP.n35 VSUBS 0.04465f
C1778 VP.n36 VSUBS 0.049028f
C1779 VP.n37 VSUBS 0.049028f
C1780 VP.n38 VSUBS 0.026438f
C1781 VP.n39 VSUBS 0.026438f
C1782 VP.n40 VSUBS 0.026438f
C1783 VP.n41 VSUBS 0.049028f
C1784 VP.n42 VSUBS 0.049028f
C1785 VP.n43 VSUBS 0.04465f
C1786 VP.n44 VSUBS 0.026438f
C1787 VP.n45 VSUBS 0.026438f
C1788 VP.n46 VSUBS 0.026438f
C1789 VP.n47 VSUBS 0.049028f
C1790 VP.n48 VSUBS 0.049028f
C1791 VP.n49 VSUBS 0.033053f
C1792 VP.n50 VSUBS 0.042664f
C1793 VP.n51 VSUBS 0.070361f
.ends

