* NGSPICE file created from diff_pair_sample_1431.ext - technology: sky130A

.subckt diff_pair_sample_1431 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t3 w_n1522_n3816# sky130_fd_pr__pfet_01v8 ad=2.3496 pd=14.57 as=5.5536 ps=29.26 w=14.24 l=0.36
X1 VDD1.t4 VP.t1 VTAIL.t8 w_n1522_n3816# sky130_fd_pr__pfet_01v8 ad=5.5536 pd=29.26 as=2.3496 ps=14.57 w=14.24 l=0.36
X2 B.t11 B.t9 B.t10 w_n1522_n3816# sky130_fd_pr__pfet_01v8 ad=5.5536 pd=29.26 as=0 ps=0 w=14.24 l=0.36
X3 B.t8 B.t6 B.t7 w_n1522_n3816# sky130_fd_pr__pfet_01v8 ad=5.5536 pd=29.26 as=0 ps=0 w=14.24 l=0.36
X4 VDD2.t5 VN.t0 VTAIL.t0 w_n1522_n3816# sky130_fd_pr__pfet_01v8 ad=5.5536 pd=29.26 as=2.3496 ps=14.57 w=14.24 l=0.36
X5 VDD2.t4 VN.t1 VTAIL.t11 w_n1522_n3816# sky130_fd_pr__pfet_01v8 ad=5.5536 pd=29.26 as=2.3496 ps=14.57 w=14.24 l=0.36
X6 VDD2.t3 VN.t2 VTAIL.t10 w_n1522_n3816# sky130_fd_pr__pfet_01v8 ad=2.3496 pd=14.57 as=5.5536 ps=29.26 w=14.24 l=0.36
X7 VTAIL.t7 VP.t2 VDD1.t3 w_n1522_n3816# sky130_fd_pr__pfet_01v8 ad=2.3496 pd=14.57 as=2.3496 ps=14.57 w=14.24 l=0.36
X8 B.t5 B.t3 B.t4 w_n1522_n3816# sky130_fd_pr__pfet_01v8 ad=5.5536 pd=29.26 as=0 ps=0 w=14.24 l=0.36
X9 VTAIL.t6 VP.t3 VDD1.t2 w_n1522_n3816# sky130_fd_pr__pfet_01v8 ad=2.3496 pd=14.57 as=2.3496 ps=14.57 w=14.24 l=0.36
X10 VDD2.t2 VN.t3 VTAIL.t1 w_n1522_n3816# sky130_fd_pr__pfet_01v8 ad=2.3496 pd=14.57 as=5.5536 ps=29.26 w=14.24 l=0.36
X11 VDD1.t1 VP.t4 VTAIL.t5 w_n1522_n3816# sky130_fd_pr__pfet_01v8 ad=5.5536 pd=29.26 as=2.3496 ps=14.57 w=14.24 l=0.36
X12 VTAIL.t9 VN.t4 VDD2.t1 w_n1522_n3816# sky130_fd_pr__pfet_01v8 ad=2.3496 pd=14.57 as=2.3496 ps=14.57 w=14.24 l=0.36
X13 VDD1.t0 VP.t5 VTAIL.t4 w_n1522_n3816# sky130_fd_pr__pfet_01v8 ad=2.3496 pd=14.57 as=5.5536 ps=29.26 w=14.24 l=0.36
X14 VTAIL.t2 VN.t5 VDD2.t0 w_n1522_n3816# sky130_fd_pr__pfet_01v8 ad=2.3496 pd=14.57 as=2.3496 ps=14.57 w=14.24 l=0.36
X15 B.t2 B.t0 B.t1 w_n1522_n3816# sky130_fd_pr__pfet_01v8 ad=5.5536 pd=29.26 as=0 ps=0 w=14.24 l=0.36
R0 VP.n1 VP.t1 1085.63
R1 VP.n8 VP.t0 1065.21
R2 VP.n6 VP.t4 1065.21
R3 VP.n3 VP.t5 1065.21
R4 VP.n7 VP.t3 1063.75
R5 VP.n2 VP.t2 1063.75
R6 VP.n9 VP.n8 161.3
R7 VP.n4 VP.n3 161.3
R8 VP.n7 VP.n0 161.3
R9 VP.n6 VP.n5 161.3
R10 VP.n4 VP.n1 70.6808
R11 VP.n7 VP.n6 46.7399
R12 VP.n8 VP.n7 46.7399
R13 VP.n3 VP.n2 46.7399
R14 VP.n5 VP.n4 41.6028
R15 VP.n2 VP.n1 20.4028
R16 VP.n5 VP.n0 0.189894
R17 VP.n9 VP.n0 0.189894
R18 VP VP.n9 0.0516364
R19 VTAIL.n314 VTAIL.n242 756.745
R20 VTAIL.n74 VTAIL.n2 756.745
R21 VTAIL.n236 VTAIL.n164 756.745
R22 VTAIL.n156 VTAIL.n84 756.745
R23 VTAIL.n266 VTAIL.n265 585
R24 VTAIL.n271 VTAIL.n270 585
R25 VTAIL.n273 VTAIL.n272 585
R26 VTAIL.n262 VTAIL.n261 585
R27 VTAIL.n279 VTAIL.n278 585
R28 VTAIL.n281 VTAIL.n280 585
R29 VTAIL.n258 VTAIL.n257 585
R30 VTAIL.n288 VTAIL.n287 585
R31 VTAIL.n289 VTAIL.n256 585
R32 VTAIL.n291 VTAIL.n290 585
R33 VTAIL.n254 VTAIL.n253 585
R34 VTAIL.n297 VTAIL.n296 585
R35 VTAIL.n299 VTAIL.n298 585
R36 VTAIL.n250 VTAIL.n249 585
R37 VTAIL.n305 VTAIL.n304 585
R38 VTAIL.n307 VTAIL.n306 585
R39 VTAIL.n246 VTAIL.n245 585
R40 VTAIL.n313 VTAIL.n312 585
R41 VTAIL.n315 VTAIL.n314 585
R42 VTAIL.n26 VTAIL.n25 585
R43 VTAIL.n31 VTAIL.n30 585
R44 VTAIL.n33 VTAIL.n32 585
R45 VTAIL.n22 VTAIL.n21 585
R46 VTAIL.n39 VTAIL.n38 585
R47 VTAIL.n41 VTAIL.n40 585
R48 VTAIL.n18 VTAIL.n17 585
R49 VTAIL.n48 VTAIL.n47 585
R50 VTAIL.n49 VTAIL.n16 585
R51 VTAIL.n51 VTAIL.n50 585
R52 VTAIL.n14 VTAIL.n13 585
R53 VTAIL.n57 VTAIL.n56 585
R54 VTAIL.n59 VTAIL.n58 585
R55 VTAIL.n10 VTAIL.n9 585
R56 VTAIL.n65 VTAIL.n64 585
R57 VTAIL.n67 VTAIL.n66 585
R58 VTAIL.n6 VTAIL.n5 585
R59 VTAIL.n73 VTAIL.n72 585
R60 VTAIL.n75 VTAIL.n74 585
R61 VTAIL.n237 VTAIL.n236 585
R62 VTAIL.n235 VTAIL.n234 585
R63 VTAIL.n168 VTAIL.n167 585
R64 VTAIL.n229 VTAIL.n228 585
R65 VTAIL.n227 VTAIL.n226 585
R66 VTAIL.n172 VTAIL.n171 585
R67 VTAIL.n221 VTAIL.n220 585
R68 VTAIL.n219 VTAIL.n218 585
R69 VTAIL.n176 VTAIL.n175 585
R70 VTAIL.n213 VTAIL.n212 585
R71 VTAIL.n211 VTAIL.n178 585
R72 VTAIL.n210 VTAIL.n209 585
R73 VTAIL.n181 VTAIL.n179 585
R74 VTAIL.n204 VTAIL.n203 585
R75 VTAIL.n202 VTAIL.n201 585
R76 VTAIL.n185 VTAIL.n184 585
R77 VTAIL.n196 VTAIL.n195 585
R78 VTAIL.n194 VTAIL.n193 585
R79 VTAIL.n189 VTAIL.n188 585
R80 VTAIL.n157 VTAIL.n156 585
R81 VTAIL.n155 VTAIL.n154 585
R82 VTAIL.n88 VTAIL.n87 585
R83 VTAIL.n149 VTAIL.n148 585
R84 VTAIL.n147 VTAIL.n146 585
R85 VTAIL.n92 VTAIL.n91 585
R86 VTAIL.n141 VTAIL.n140 585
R87 VTAIL.n139 VTAIL.n138 585
R88 VTAIL.n96 VTAIL.n95 585
R89 VTAIL.n133 VTAIL.n132 585
R90 VTAIL.n131 VTAIL.n98 585
R91 VTAIL.n130 VTAIL.n129 585
R92 VTAIL.n101 VTAIL.n99 585
R93 VTAIL.n124 VTAIL.n123 585
R94 VTAIL.n122 VTAIL.n121 585
R95 VTAIL.n105 VTAIL.n104 585
R96 VTAIL.n116 VTAIL.n115 585
R97 VTAIL.n114 VTAIL.n113 585
R98 VTAIL.n109 VTAIL.n108 585
R99 VTAIL.n267 VTAIL.t1 329.036
R100 VTAIL.n27 VTAIL.t3 329.036
R101 VTAIL.n110 VTAIL.t10 329.036
R102 VTAIL.n190 VTAIL.t4 329.036
R103 VTAIL.n271 VTAIL.n265 171.744
R104 VTAIL.n272 VTAIL.n271 171.744
R105 VTAIL.n272 VTAIL.n261 171.744
R106 VTAIL.n279 VTAIL.n261 171.744
R107 VTAIL.n280 VTAIL.n279 171.744
R108 VTAIL.n280 VTAIL.n257 171.744
R109 VTAIL.n288 VTAIL.n257 171.744
R110 VTAIL.n289 VTAIL.n288 171.744
R111 VTAIL.n290 VTAIL.n289 171.744
R112 VTAIL.n290 VTAIL.n253 171.744
R113 VTAIL.n297 VTAIL.n253 171.744
R114 VTAIL.n298 VTAIL.n297 171.744
R115 VTAIL.n298 VTAIL.n249 171.744
R116 VTAIL.n305 VTAIL.n249 171.744
R117 VTAIL.n306 VTAIL.n305 171.744
R118 VTAIL.n306 VTAIL.n245 171.744
R119 VTAIL.n313 VTAIL.n245 171.744
R120 VTAIL.n314 VTAIL.n313 171.744
R121 VTAIL.n31 VTAIL.n25 171.744
R122 VTAIL.n32 VTAIL.n31 171.744
R123 VTAIL.n32 VTAIL.n21 171.744
R124 VTAIL.n39 VTAIL.n21 171.744
R125 VTAIL.n40 VTAIL.n39 171.744
R126 VTAIL.n40 VTAIL.n17 171.744
R127 VTAIL.n48 VTAIL.n17 171.744
R128 VTAIL.n49 VTAIL.n48 171.744
R129 VTAIL.n50 VTAIL.n49 171.744
R130 VTAIL.n50 VTAIL.n13 171.744
R131 VTAIL.n57 VTAIL.n13 171.744
R132 VTAIL.n58 VTAIL.n57 171.744
R133 VTAIL.n58 VTAIL.n9 171.744
R134 VTAIL.n65 VTAIL.n9 171.744
R135 VTAIL.n66 VTAIL.n65 171.744
R136 VTAIL.n66 VTAIL.n5 171.744
R137 VTAIL.n73 VTAIL.n5 171.744
R138 VTAIL.n74 VTAIL.n73 171.744
R139 VTAIL.n236 VTAIL.n235 171.744
R140 VTAIL.n235 VTAIL.n167 171.744
R141 VTAIL.n228 VTAIL.n167 171.744
R142 VTAIL.n228 VTAIL.n227 171.744
R143 VTAIL.n227 VTAIL.n171 171.744
R144 VTAIL.n220 VTAIL.n171 171.744
R145 VTAIL.n220 VTAIL.n219 171.744
R146 VTAIL.n219 VTAIL.n175 171.744
R147 VTAIL.n212 VTAIL.n175 171.744
R148 VTAIL.n212 VTAIL.n211 171.744
R149 VTAIL.n211 VTAIL.n210 171.744
R150 VTAIL.n210 VTAIL.n179 171.744
R151 VTAIL.n203 VTAIL.n179 171.744
R152 VTAIL.n203 VTAIL.n202 171.744
R153 VTAIL.n202 VTAIL.n184 171.744
R154 VTAIL.n195 VTAIL.n184 171.744
R155 VTAIL.n195 VTAIL.n194 171.744
R156 VTAIL.n194 VTAIL.n188 171.744
R157 VTAIL.n156 VTAIL.n155 171.744
R158 VTAIL.n155 VTAIL.n87 171.744
R159 VTAIL.n148 VTAIL.n87 171.744
R160 VTAIL.n148 VTAIL.n147 171.744
R161 VTAIL.n147 VTAIL.n91 171.744
R162 VTAIL.n140 VTAIL.n91 171.744
R163 VTAIL.n140 VTAIL.n139 171.744
R164 VTAIL.n139 VTAIL.n95 171.744
R165 VTAIL.n132 VTAIL.n95 171.744
R166 VTAIL.n132 VTAIL.n131 171.744
R167 VTAIL.n131 VTAIL.n130 171.744
R168 VTAIL.n130 VTAIL.n99 171.744
R169 VTAIL.n123 VTAIL.n99 171.744
R170 VTAIL.n123 VTAIL.n122 171.744
R171 VTAIL.n122 VTAIL.n104 171.744
R172 VTAIL.n115 VTAIL.n104 171.744
R173 VTAIL.n115 VTAIL.n114 171.744
R174 VTAIL.n114 VTAIL.n108 171.744
R175 VTAIL.t1 VTAIL.n265 85.8723
R176 VTAIL.t3 VTAIL.n25 85.8723
R177 VTAIL.t4 VTAIL.n188 85.8723
R178 VTAIL.t10 VTAIL.n108 85.8723
R179 VTAIL.n1 VTAIL.n0 54.1784
R180 VTAIL.n81 VTAIL.n80 54.1784
R181 VTAIL.n163 VTAIL.n162 54.1784
R182 VTAIL.n83 VTAIL.n82 54.1784
R183 VTAIL.n319 VTAIL.n318 31.4096
R184 VTAIL.n79 VTAIL.n78 31.4096
R185 VTAIL.n241 VTAIL.n240 31.4096
R186 VTAIL.n161 VTAIL.n160 31.4096
R187 VTAIL.n83 VTAIL.n81 25.8324
R188 VTAIL.n319 VTAIL.n241 25.2376
R189 VTAIL.n291 VTAIL.n256 13.1884
R190 VTAIL.n51 VTAIL.n16 13.1884
R191 VTAIL.n213 VTAIL.n178 13.1884
R192 VTAIL.n133 VTAIL.n98 13.1884
R193 VTAIL.n287 VTAIL.n286 12.8005
R194 VTAIL.n292 VTAIL.n254 12.8005
R195 VTAIL.n47 VTAIL.n46 12.8005
R196 VTAIL.n52 VTAIL.n14 12.8005
R197 VTAIL.n214 VTAIL.n176 12.8005
R198 VTAIL.n209 VTAIL.n180 12.8005
R199 VTAIL.n134 VTAIL.n96 12.8005
R200 VTAIL.n129 VTAIL.n100 12.8005
R201 VTAIL.n285 VTAIL.n258 12.0247
R202 VTAIL.n296 VTAIL.n295 12.0247
R203 VTAIL.n45 VTAIL.n18 12.0247
R204 VTAIL.n56 VTAIL.n55 12.0247
R205 VTAIL.n218 VTAIL.n217 12.0247
R206 VTAIL.n208 VTAIL.n181 12.0247
R207 VTAIL.n138 VTAIL.n137 12.0247
R208 VTAIL.n128 VTAIL.n101 12.0247
R209 VTAIL.n282 VTAIL.n281 11.249
R210 VTAIL.n299 VTAIL.n252 11.249
R211 VTAIL.n42 VTAIL.n41 11.249
R212 VTAIL.n59 VTAIL.n12 11.249
R213 VTAIL.n221 VTAIL.n174 11.249
R214 VTAIL.n205 VTAIL.n204 11.249
R215 VTAIL.n141 VTAIL.n94 11.249
R216 VTAIL.n125 VTAIL.n124 11.249
R217 VTAIL.n267 VTAIL.n266 10.7239
R218 VTAIL.n27 VTAIL.n26 10.7239
R219 VTAIL.n190 VTAIL.n189 10.7239
R220 VTAIL.n110 VTAIL.n109 10.7239
R221 VTAIL.n278 VTAIL.n260 10.4732
R222 VTAIL.n300 VTAIL.n250 10.4732
R223 VTAIL.n38 VTAIL.n20 10.4732
R224 VTAIL.n60 VTAIL.n10 10.4732
R225 VTAIL.n222 VTAIL.n172 10.4732
R226 VTAIL.n201 VTAIL.n183 10.4732
R227 VTAIL.n142 VTAIL.n92 10.4732
R228 VTAIL.n121 VTAIL.n103 10.4732
R229 VTAIL.n277 VTAIL.n262 9.69747
R230 VTAIL.n304 VTAIL.n303 9.69747
R231 VTAIL.n37 VTAIL.n22 9.69747
R232 VTAIL.n64 VTAIL.n63 9.69747
R233 VTAIL.n226 VTAIL.n225 9.69747
R234 VTAIL.n200 VTAIL.n185 9.69747
R235 VTAIL.n146 VTAIL.n145 9.69747
R236 VTAIL.n120 VTAIL.n105 9.69747
R237 VTAIL.n318 VTAIL.n317 9.45567
R238 VTAIL.n78 VTAIL.n77 9.45567
R239 VTAIL.n240 VTAIL.n239 9.45567
R240 VTAIL.n160 VTAIL.n159 9.45567
R241 VTAIL.n244 VTAIL.n243 9.3005
R242 VTAIL.n317 VTAIL.n316 9.3005
R243 VTAIL.n309 VTAIL.n308 9.3005
R244 VTAIL.n248 VTAIL.n247 9.3005
R245 VTAIL.n303 VTAIL.n302 9.3005
R246 VTAIL.n301 VTAIL.n300 9.3005
R247 VTAIL.n252 VTAIL.n251 9.3005
R248 VTAIL.n295 VTAIL.n294 9.3005
R249 VTAIL.n293 VTAIL.n292 9.3005
R250 VTAIL.n269 VTAIL.n268 9.3005
R251 VTAIL.n264 VTAIL.n263 9.3005
R252 VTAIL.n275 VTAIL.n274 9.3005
R253 VTAIL.n277 VTAIL.n276 9.3005
R254 VTAIL.n260 VTAIL.n259 9.3005
R255 VTAIL.n283 VTAIL.n282 9.3005
R256 VTAIL.n285 VTAIL.n284 9.3005
R257 VTAIL.n286 VTAIL.n255 9.3005
R258 VTAIL.n311 VTAIL.n310 9.3005
R259 VTAIL.n4 VTAIL.n3 9.3005
R260 VTAIL.n77 VTAIL.n76 9.3005
R261 VTAIL.n69 VTAIL.n68 9.3005
R262 VTAIL.n8 VTAIL.n7 9.3005
R263 VTAIL.n63 VTAIL.n62 9.3005
R264 VTAIL.n61 VTAIL.n60 9.3005
R265 VTAIL.n12 VTAIL.n11 9.3005
R266 VTAIL.n55 VTAIL.n54 9.3005
R267 VTAIL.n53 VTAIL.n52 9.3005
R268 VTAIL.n29 VTAIL.n28 9.3005
R269 VTAIL.n24 VTAIL.n23 9.3005
R270 VTAIL.n35 VTAIL.n34 9.3005
R271 VTAIL.n37 VTAIL.n36 9.3005
R272 VTAIL.n20 VTAIL.n19 9.3005
R273 VTAIL.n43 VTAIL.n42 9.3005
R274 VTAIL.n45 VTAIL.n44 9.3005
R275 VTAIL.n46 VTAIL.n15 9.3005
R276 VTAIL.n71 VTAIL.n70 9.3005
R277 VTAIL.n166 VTAIL.n165 9.3005
R278 VTAIL.n233 VTAIL.n232 9.3005
R279 VTAIL.n231 VTAIL.n230 9.3005
R280 VTAIL.n170 VTAIL.n169 9.3005
R281 VTAIL.n225 VTAIL.n224 9.3005
R282 VTAIL.n223 VTAIL.n222 9.3005
R283 VTAIL.n174 VTAIL.n173 9.3005
R284 VTAIL.n217 VTAIL.n216 9.3005
R285 VTAIL.n215 VTAIL.n214 9.3005
R286 VTAIL.n180 VTAIL.n177 9.3005
R287 VTAIL.n208 VTAIL.n207 9.3005
R288 VTAIL.n206 VTAIL.n205 9.3005
R289 VTAIL.n183 VTAIL.n182 9.3005
R290 VTAIL.n200 VTAIL.n199 9.3005
R291 VTAIL.n198 VTAIL.n197 9.3005
R292 VTAIL.n187 VTAIL.n186 9.3005
R293 VTAIL.n192 VTAIL.n191 9.3005
R294 VTAIL.n239 VTAIL.n238 9.3005
R295 VTAIL.n112 VTAIL.n111 9.3005
R296 VTAIL.n107 VTAIL.n106 9.3005
R297 VTAIL.n118 VTAIL.n117 9.3005
R298 VTAIL.n120 VTAIL.n119 9.3005
R299 VTAIL.n103 VTAIL.n102 9.3005
R300 VTAIL.n126 VTAIL.n125 9.3005
R301 VTAIL.n128 VTAIL.n127 9.3005
R302 VTAIL.n100 VTAIL.n97 9.3005
R303 VTAIL.n159 VTAIL.n158 9.3005
R304 VTAIL.n86 VTAIL.n85 9.3005
R305 VTAIL.n153 VTAIL.n152 9.3005
R306 VTAIL.n151 VTAIL.n150 9.3005
R307 VTAIL.n90 VTAIL.n89 9.3005
R308 VTAIL.n145 VTAIL.n144 9.3005
R309 VTAIL.n143 VTAIL.n142 9.3005
R310 VTAIL.n94 VTAIL.n93 9.3005
R311 VTAIL.n137 VTAIL.n136 9.3005
R312 VTAIL.n135 VTAIL.n134 9.3005
R313 VTAIL.n274 VTAIL.n273 8.92171
R314 VTAIL.n307 VTAIL.n248 8.92171
R315 VTAIL.n34 VTAIL.n33 8.92171
R316 VTAIL.n67 VTAIL.n8 8.92171
R317 VTAIL.n229 VTAIL.n170 8.92171
R318 VTAIL.n197 VTAIL.n196 8.92171
R319 VTAIL.n149 VTAIL.n90 8.92171
R320 VTAIL.n117 VTAIL.n116 8.92171
R321 VTAIL.n270 VTAIL.n264 8.14595
R322 VTAIL.n308 VTAIL.n246 8.14595
R323 VTAIL.n318 VTAIL.n242 8.14595
R324 VTAIL.n30 VTAIL.n24 8.14595
R325 VTAIL.n68 VTAIL.n6 8.14595
R326 VTAIL.n78 VTAIL.n2 8.14595
R327 VTAIL.n240 VTAIL.n164 8.14595
R328 VTAIL.n230 VTAIL.n168 8.14595
R329 VTAIL.n193 VTAIL.n187 8.14595
R330 VTAIL.n160 VTAIL.n84 8.14595
R331 VTAIL.n150 VTAIL.n88 8.14595
R332 VTAIL.n113 VTAIL.n107 8.14595
R333 VTAIL.n269 VTAIL.n266 7.3702
R334 VTAIL.n312 VTAIL.n311 7.3702
R335 VTAIL.n316 VTAIL.n315 7.3702
R336 VTAIL.n29 VTAIL.n26 7.3702
R337 VTAIL.n72 VTAIL.n71 7.3702
R338 VTAIL.n76 VTAIL.n75 7.3702
R339 VTAIL.n238 VTAIL.n237 7.3702
R340 VTAIL.n234 VTAIL.n233 7.3702
R341 VTAIL.n192 VTAIL.n189 7.3702
R342 VTAIL.n158 VTAIL.n157 7.3702
R343 VTAIL.n154 VTAIL.n153 7.3702
R344 VTAIL.n112 VTAIL.n109 7.3702
R345 VTAIL.n312 VTAIL.n244 6.59444
R346 VTAIL.n315 VTAIL.n244 6.59444
R347 VTAIL.n72 VTAIL.n4 6.59444
R348 VTAIL.n75 VTAIL.n4 6.59444
R349 VTAIL.n237 VTAIL.n166 6.59444
R350 VTAIL.n234 VTAIL.n166 6.59444
R351 VTAIL.n157 VTAIL.n86 6.59444
R352 VTAIL.n154 VTAIL.n86 6.59444
R353 VTAIL.n270 VTAIL.n269 5.81868
R354 VTAIL.n311 VTAIL.n246 5.81868
R355 VTAIL.n316 VTAIL.n242 5.81868
R356 VTAIL.n30 VTAIL.n29 5.81868
R357 VTAIL.n71 VTAIL.n6 5.81868
R358 VTAIL.n76 VTAIL.n2 5.81868
R359 VTAIL.n238 VTAIL.n164 5.81868
R360 VTAIL.n233 VTAIL.n168 5.81868
R361 VTAIL.n193 VTAIL.n192 5.81868
R362 VTAIL.n158 VTAIL.n84 5.81868
R363 VTAIL.n153 VTAIL.n88 5.81868
R364 VTAIL.n113 VTAIL.n112 5.81868
R365 VTAIL.n273 VTAIL.n264 5.04292
R366 VTAIL.n308 VTAIL.n307 5.04292
R367 VTAIL.n33 VTAIL.n24 5.04292
R368 VTAIL.n68 VTAIL.n67 5.04292
R369 VTAIL.n230 VTAIL.n229 5.04292
R370 VTAIL.n196 VTAIL.n187 5.04292
R371 VTAIL.n150 VTAIL.n149 5.04292
R372 VTAIL.n116 VTAIL.n107 5.04292
R373 VTAIL.n274 VTAIL.n262 4.26717
R374 VTAIL.n304 VTAIL.n248 4.26717
R375 VTAIL.n34 VTAIL.n22 4.26717
R376 VTAIL.n64 VTAIL.n8 4.26717
R377 VTAIL.n226 VTAIL.n170 4.26717
R378 VTAIL.n197 VTAIL.n185 4.26717
R379 VTAIL.n146 VTAIL.n90 4.26717
R380 VTAIL.n117 VTAIL.n105 4.26717
R381 VTAIL.n278 VTAIL.n277 3.49141
R382 VTAIL.n303 VTAIL.n250 3.49141
R383 VTAIL.n38 VTAIL.n37 3.49141
R384 VTAIL.n63 VTAIL.n10 3.49141
R385 VTAIL.n225 VTAIL.n172 3.49141
R386 VTAIL.n201 VTAIL.n200 3.49141
R387 VTAIL.n145 VTAIL.n92 3.49141
R388 VTAIL.n121 VTAIL.n120 3.49141
R389 VTAIL.n281 VTAIL.n260 2.71565
R390 VTAIL.n300 VTAIL.n299 2.71565
R391 VTAIL.n41 VTAIL.n20 2.71565
R392 VTAIL.n60 VTAIL.n59 2.71565
R393 VTAIL.n222 VTAIL.n221 2.71565
R394 VTAIL.n204 VTAIL.n183 2.71565
R395 VTAIL.n142 VTAIL.n141 2.71565
R396 VTAIL.n124 VTAIL.n103 2.71565
R397 VTAIL.n191 VTAIL.n190 2.41282
R398 VTAIL.n111 VTAIL.n110 2.41282
R399 VTAIL.n268 VTAIL.n267 2.41282
R400 VTAIL.n28 VTAIL.n27 2.41282
R401 VTAIL.n0 VTAIL.t0 2.28315
R402 VTAIL.n0 VTAIL.t2 2.28315
R403 VTAIL.n80 VTAIL.t5 2.28315
R404 VTAIL.n80 VTAIL.t6 2.28315
R405 VTAIL.n162 VTAIL.t8 2.28315
R406 VTAIL.n162 VTAIL.t7 2.28315
R407 VTAIL.n82 VTAIL.t11 2.28315
R408 VTAIL.n82 VTAIL.t9 2.28315
R409 VTAIL.n282 VTAIL.n258 1.93989
R410 VTAIL.n296 VTAIL.n252 1.93989
R411 VTAIL.n42 VTAIL.n18 1.93989
R412 VTAIL.n56 VTAIL.n12 1.93989
R413 VTAIL.n218 VTAIL.n174 1.93989
R414 VTAIL.n205 VTAIL.n181 1.93989
R415 VTAIL.n138 VTAIL.n94 1.93989
R416 VTAIL.n125 VTAIL.n101 1.93989
R417 VTAIL.n287 VTAIL.n285 1.16414
R418 VTAIL.n295 VTAIL.n254 1.16414
R419 VTAIL.n47 VTAIL.n45 1.16414
R420 VTAIL.n55 VTAIL.n14 1.16414
R421 VTAIL.n217 VTAIL.n176 1.16414
R422 VTAIL.n209 VTAIL.n208 1.16414
R423 VTAIL.n137 VTAIL.n96 1.16414
R424 VTAIL.n129 VTAIL.n128 1.16414
R425 VTAIL.n163 VTAIL.n161 0.767741
R426 VTAIL.n79 VTAIL.n1 0.767741
R427 VTAIL.n161 VTAIL.n83 0.595328
R428 VTAIL.n241 VTAIL.n163 0.595328
R429 VTAIL.n81 VTAIL.n79 0.595328
R430 VTAIL VTAIL.n319 0.388431
R431 VTAIL.n286 VTAIL.n256 0.388379
R432 VTAIL.n292 VTAIL.n291 0.388379
R433 VTAIL.n46 VTAIL.n16 0.388379
R434 VTAIL.n52 VTAIL.n51 0.388379
R435 VTAIL.n214 VTAIL.n213 0.388379
R436 VTAIL.n180 VTAIL.n178 0.388379
R437 VTAIL.n134 VTAIL.n133 0.388379
R438 VTAIL.n100 VTAIL.n98 0.388379
R439 VTAIL VTAIL.n1 0.207397
R440 VTAIL.n268 VTAIL.n263 0.155672
R441 VTAIL.n275 VTAIL.n263 0.155672
R442 VTAIL.n276 VTAIL.n275 0.155672
R443 VTAIL.n276 VTAIL.n259 0.155672
R444 VTAIL.n283 VTAIL.n259 0.155672
R445 VTAIL.n284 VTAIL.n283 0.155672
R446 VTAIL.n284 VTAIL.n255 0.155672
R447 VTAIL.n293 VTAIL.n255 0.155672
R448 VTAIL.n294 VTAIL.n293 0.155672
R449 VTAIL.n294 VTAIL.n251 0.155672
R450 VTAIL.n301 VTAIL.n251 0.155672
R451 VTAIL.n302 VTAIL.n301 0.155672
R452 VTAIL.n302 VTAIL.n247 0.155672
R453 VTAIL.n309 VTAIL.n247 0.155672
R454 VTAIL.n310 VTAIL.n309 0.155672
R455 VTAIL.n310 VTAIL.n243 0.155672
R456 VTAIL.n317 VTAIL.n243 0.155672
R457 VTAIL.n28 VTAIL.n23 0.155672
R458 VTAIL.n35 VTAIL.n23 0.155672
R459 VTAIL.n36 VTAIL.n35 0.155672
R460 VTAIL.n36 VTAIL.n19 0.155672
R461 VTAIL.n43 VTAIL.n19 0.155672
R462 VTAIL.n44 VTAIL.n43 0.155672
R463 VTAIL.n44 VTAIL.n15 0.155672
R464 VTAIL.n53 VTAIL.n15 0.155672
R465 VTAIL.n54 VTAIL.n53 0.155672
R466 VTAIL.n54 VTAIL.n11 0.155672
R467 VTAIL.n61 VTAIL.n11 0.155672
R468 VTAIL.n62 VTAIL.n61 0.155672
R469 VTAIL.n62 VTAIL.n7 0.155672
R470 VTAIL.n69 VTAIL.n7 0.155672
R471 VTAIL.n70 VTAIL.n69 0.155672
R472 VTAIL.n70 VTAIL.n3 0.155672
R473 VTAIL.n77 VTAIL.n3 0.155672
R474 VTAIL.n239 VTAIL.n165 0.155672
R475 VTAIL.n232 VTAIL.n165 0.155672
R476 VTAIL.n232 VTAIL.n231 0.155672
R477 VTAIL.n231 VTAIL.n169 0.155672
R478 VTAIL.n224 VTAIL.n169 0.155672
R479 VTAIL.n224 VTAIL.n223 0.155672
R480 VTAIL.n223 VTAIL.n173 0.155672
R481 VTAIL.n216 VTAIL.n173 0.155672
R482 VTAIL.n216 VTAIL.n215 0.155672
R483 VTAIL.n215 VTAIL.n177 0.155672
R484 VTAIL.n207 VTAIL.n177 0.155672
R485 VTAIL.n207 VTAIL.n206 0.155672
R486 VTAIL.n206 VTAIL.n182 0.155672
R487 VTAIL.n199 VTAIL.n182 0.155672
R488 VTAIL.n199 VTAIL.n198 0.155672
R489 VTAIL.n198 VTAIL.n186 0.155672
R490 VTAIL.n191 VTAIL.n186 0.155672
R491 VTAIL.n159 VTAIL.n85 0.155672
R492 VTAIL.n152 VTAIL.n85 0.155672
R493 VTAIL.n152 VTAIL.n151 0.155672
R494 VTAIL.n151 VTAIL.n89 0.155672
R495 VTAIL.n144 VTAIL.n89 0.155672
R496 VTAIL.n144 VTAIL.n143 0.155672
R497 VTAIL.n143 VTAIL.n93 0.155672
R498 VTAIL.n136 VTAIL.n93 0.155672
R499 VTAIL.n136 VTAIL.n135 0.155672
R500 VTAIL.n135 VTAIL.n97 0.155672
R501 VTAIL.n127 VTAIL.n97 0.155672
R502 VTAIL.n127 VTAIL.n126 0.155672
R503 VTAIL.n126 VTAIL.n102 0.155672
R504 VTAIL.n119 VTAIL.n102 0.155672
R505 VTAIL.n119 VTAIL.n118 0.155672
R506 VTAIL.n118 VTAIL.n106 0.155672
R507 VTAIL.n111 VTAIL.n106 0.155672
R508 VDD1.n72 VDD1.n0 756.745
R509 VDD1.n149 VDD1.n77 756.745
R510 VDD1.n73 VDD1.n72 585
R511 VDD1.n71 VDD1.n70 585
R512 VDD1.n4 VDD1.n3 585
R513 VDD1.n65 VDD1.n64 585
R514 VDD1.n63 VDD1.n62 585
R515 VDD1.n8 VDD1.n7 585
R516 VDD1.n57 VDD1.n56 585
R517 VDD1.n55 VDD1.n54 585
R518 VDD1.n12 VDD1.n11 585
R519 VDD1.n49 VDD1.n48 585
R520 VDD1.n47 VDD1.n14 585
R521 VDD1.n46 VDD1.n45 585
R522 VDD1.n17 VDD1.n15 585
R523 VDD1.n40 VDD1.n39 585
R524 VDD1.n38 VDD1.n37 585
R525 VDD1.n21 VDD1.n20 585
R526 VDD1.n32 VDD1.n31 585
R527 VDD1.n30 VDD1.n29 585
R528 VDD1.n25 VDD1.n24 585
R529 VDD1.n101 VDD1.n100 585
R530 VDD1.n106 VDD1.n105 585
R531 VDD1.n108 VDD1.n107 585
R532 VDD1.n97 VDD1.n96 585
R533 VDD1.n114 VDD1.n113 585
R534 VDD1.n116 VDD1.n115 585
R535 VDD1.n93 VDD1.n92 585
R536 VDD1.n123 VDD1.n122 585
R537 VDD1.n124 VDD1.n91 585
R538 VDD1.n126 VDD1.n125 585
R539 VDD1.n89 VDD1.n88 585
R540 VDD1.n132 VDD1.n131 585
R541 VDD1.n134 VDD1.n133 585
R542 VDD1.n85 VDD1.n84 585
R543 VDD1.n140 VDD1.n139 585
R544 VDD1.n142 VDD1.n141 585
R545 VDD1.n81 VDD1.n80 585
R546 VDD1.n148 VDD1.n147 585
R547 VDD1.n150 VDD1.n149 585
R548 VDD1.n26 VDD1.t4 329.036
R549 VDD1.n102 VDD1.t1 329.036
R550 VDD1.n72 VDD1.n71 171.744
R551 VDD1.n71 VDD1.n3 171.744
R552 VDD1.n64 VDD1.n3 171.744
R553 VDD1.n64 VDD1.n63 171.744
R554 VDD1.n63 VDD1.n7 171.744
R555 VDD1.n56 VDD1.n7 171.744
R556 VDD1.n56 VDD1.n55 171.744
R557 VDD1.n55 VDD1.n11 171.744
R558 VDD1.n48 VDD1.n11 171.744
R559 VDD1.n48 VDD1.n47 171.744
R560 VDD1.n47 VDD1.n46 171.744
R561 VDD1.n46 VDD1.n15 171.744
R562 VDD1.n39 VDD1.n15 171.744
R563 VDD1.n39 VDD1.n38 171.744
R564 VDD1.n38 VDD1.n20 171.744
R565 VDD1.n31 VDD1.n20 171.744
R566 VDD1.n31 VDD1.n30 171.744
R567 VDD1.n30 VDD1.n24 171.744
R568 VDD1.n106 VDD1.n100 171.744
R569 VDD1.n107 VDD1.n106 171.744
R570 VDD1.n107 VDD1.n96 171.744
R571 VDD1.n114 VDD1.n96 171.744
R572 VDD1.n115 VDD1.n114 171.744
R573 VDD1.n115 VDD1.n92 171.744
R574 VDD1.n123 VDD1.n92 171.744
R575 VDD1.n124 VDD1.n123 171.744
R576 VDD1.n125 VDD1.n124 171.744
R577 VDD1.n125 VDD1.n88 171.744
R578 VDD1.n132 VDD1.n88 171.744
R579 VDD1.n133 VDD1.n132 171.744
R580 VDD1.n133 VDD1.n84 171.744
R581 VDD1.n140 VDD1.n84 171.744
R582 VDD1.n141 VDD1.n140 171.744
R583 VDD1.n141 VDD1.n80 171.744
R584 VDD1.n148 VDD1.n80 171.744
R585 VDD1.n149 VDD1.n148 171.744
R586 VDD1.t4 VDD1.n24 85.8723
R587 VDD1.t1 VDD1.n100 85.8723
R588 VDD1.n155 VDD1.n154 70.9506
R589 VDD1.n157 VDD1.n156 70.8572
R590 VDD1 VDD1.n76 48.5927
R591 VDD1.n155 VDD1.n153 48.4792
R592 VDD1.n157 VDD1.n155 38.8048
R593 VDD1.n49 VDD1.n14 13.1884
R594 VDD1.n126 VDD1.n91 13.1884
R595 VDD1.n50 VDD1.n12 12.8005
R596 VDD1.n45 VDD1.n16 12.8005
R597 VDD1.n122 VDD1.n121 12.8005
R598 VDD1.n127 VDD1.n89 12.8005
R599 VDD1.n54 VDD1.n53 12.0247
R600 VDD1.n44 VDD1.n17 12.0247
R601 VDD1.n120 VDD1.n93 12.0247
R602 VDD1.n131 VDD1.n130 12.0247
R603 VDD1.n57 VDD1.n10 11.249
R604 VDD1.n41 VDD1.n40 11.249
R605 VDD1.n117 VDD1.n116 11.249
R606 VDD1.n134 VDD1.n87 11.249
R607 VDD1.n26 VDD1.n25 10.7239
R608 VDD1.n102 VDD1.n101 10.7239
R609 VDD1.n58 VDD1.n8 10.4732
R610 VDD1.n37 VDD1.n19 10.4732
R611 VDD1.n113 VDD1.n95 10.4732
R612 VDD1.n135 VDD1.n85 10.4732
R613 VDD1.n62 VDD1.n61 9.69747
R614 VDD1.n36 VDD1.n21 9.69747
R615 VDD1.n112 VDD1.n97 9.69747
R616 VDD1.n139 VDD1.n138 9.69747
R617 VDD1.n76 VDD1.n75 9.45567
R618 VDD1.n153 VDD1.n152 9.45567
R619 VDD1.n28 VDD1.n27 9.3005
R620 VDD1.n23 VDD1.n22 9.3005
R621 VDD1.n34 VDD1.n33 9.3005
R622 VDD1.n36 VDD1.n35 9.3005
R623 VDD1.n19 VDD1.n18 9.3005
R624 VDD1.n42 VDD1.n41 9.3005
R625 VDD1.n44 VDD1.n43 9.3005
R626 VDD1.n16 VDD1.n13 9.3005
R627 VDD1.n75 VDD1.n74 9.3005
R628 VDD1.n2 VDD1.n1 9.3005
R629 VDD1.n69 VDD1.n68 9.3005
R630 VDD1.n67 VDD1.n66 9.3005
R631 VDD1.n6 VDD1.n5 9.3005
R632 VDD1.n61 VDD1.n60 9.3005
R633 VDD1.n59 VDD1.n58 9.3005
R634 VDD1.n10 VDD1.n9 9.3005
R635 VDD1.n53 VDD1.n52 9.3005
R636 VDD1.n51 VDD1.n50 9.3005
R637 VDD1.n79 VDD1.n78 9.3005
R638 VDD1.n152 VDD1.n151 9.3005
R639 VDD1.n144 VDD1.n143 9.3005
R640 VDD1.n83 VDD1.n82 9.3005
R641 VDD1.n138 VDD1.n137 9.3005
R642 VDD1.n136 VDD1.n135 9.3005
R643 VDD1.n87 VDD1.n86 9.3005
R644 VDD1.n130 VDD1.n129 9.3005
R645 VDD1.n128 VDD1.n127 9.3005
R646 VDD1.n104 VDD1.n103 9.3005
R647 VDD1.n99 VDD1.n98 9.3005
R648 VDD1.n110 VDD1.n109 9.3005
R649 VDD1.n112 VDD1.n111 9.3005
R650 VDD1.n95 VDD1.n94 9.3005
R651 VDD1.n118 VDD1.n117 9.3005
R652 VDD1.n120 VDD1.n119 9.3005
R653 VDD1.n121 VDD1.n90 9.3005
R654 VDD1.n146 VDD1.n145 9.3005
R655 VDD1.n65 VDD1.n6 8.92171
R656 VDD1.n33 VDD1.n32 8.92171
R657 VDD1.n109 VDD1.n108 8.92171
R658 VDD1.n142 VDD1.n83 8.92171
R659 VDD1.n76 VDD1.n0 8.14595
R660 VDD1.n66 VDD1.n4 8.14595
R661 VDD1.n29 VDD1.n23 8.14595
R662 VDD1.n105 VDD1.n99 8.14595
R663 VDD1.n143 VDD1.n81 8.14595
R664 VDD1.n153 VDD1.n77 8.14595
R665 VDD1.n74 VDD1.n73 7.3702
R666 VDD1.n70 VDD1.n69 7.3702
R667 VDD1.n28 VDD1.n25 7.3702
R668 VDD1.n104 VDD1.n101 7.3702
R669 VDD1.n147 VDD1.n146 7.3702
R670 VDD1.n151 VDD1.n150 7.3702
R671 VDD1.n73 VDD1.n2 6.59444
R672 VDD1.n70 VDD1.n2 6.59444
R673 VDD1.n147 VDD1.n79 6.59444
R674 VDD1.n150 VDD1.n79 6.59444
R675 VDD1.n74 VDD1.n0 5.81868
R676 VDD1.n69 VDD1.n4 5.81868
R677 VDD1.n29 VDD1.n28 5.81868
R678 VDD1.n105 VDD1.n104 5.81868
R679 VDD1.n146 VDD1.n81 5.81868
R680 VDD1.n151 VDD1.n77 5.81868
R681 VDD1.n66 VDD1.n65 5.04292
R682 VDD1.n32 VDD1.n23 5.04292
R683 VDD1.n108 VDD1.n99 5.04292
R684 VDD1.n143 VDD1.n142 5.04292
R685 VDD1.n62 VDD1.n6 4.26717
R686 VDD1.n33 VDD1.n21 4.26717
R687 VDD1.n109 VDD1.n97 4.26717
R688 VDD1.n139 VDD1.n83 4.26717
R689 VDD1.n61 VDD1.n8 3.49141
R690 VDD1.n37 VDD1.n36 3.49141
R691 VDD1.n113 VDD1.n112 3.49141
R692 VDD1.n138 VDD1.n85 3.49141
R693 VDD1.n58 VDD1.n57 2.71565
R694 VDD1.n40 VDD1.n19 2.71565
R695 VDD1.n116 VDD1.n95 2.71565
R696 VDD1.n135 VDD1.n134 2.71565
R697 VDD1.n27 VDD1.n26 2.41282
R698 VDD1.n103 VDD1.n102 2.41282
R699 VDD1.n156 VDD1.t3 2.28315
R700 VDD1.n156 VDD1.t0 2.28315
R701 VDD1.n154 VDD1.t2 2.28315
R702 VDD1.n154 VDD1.t5 2.28315
R703 VDD1.n54 VDD1.n10 1.93989
R704 VDD1.n41 VDD1.n17 1.93989
R705 VDD1.n117 VDD1.n93 1.93989
R706 VDD1.n131 VDD1.n87 1.93989
R707 VDD1.n53 VDD1.n12 1.16414
R708 VDD1.n45 VDD1.n44 1.16414
R709 VDD1.n122 VDD1.n120 1.16414
R710 VDD1.n130 VDD1.n89 1.16414
R711 VDD1.n50 VDD1.n49 0.388379
R712 VDD1.n16 VDD1.n14 0.388379
R713 VDD1.n121 VDD1.n91 0.388379
R714 VDD1.n127 VDD1.n126 0.388379
R715 VDD1.n75 VDD1.n1 0.155672
R716 VDD1.n68 VDD1.n1 0.155672
R717 VDD1.n68 VDD1.n67 0.155672
R718 VDD1.n67 VDD1.n5 0.155672
R719 VDD1.n60 VDD1.n5 0.155672
R720 VDD1.n60 VDD1.n59 0.155672
R721 VDD1.n59 VDD1.n9 0.155672
R722 VDD1.n52 VDD1.n9 0.155672
R723 VDD1.n52 VDD1.n51 0.155672
R724 VDD1.n51 VDD1.n13 0.155672
R725 VDD1.n43 VDD1.n13 0.155672
R726 VDD1.n43 VDD1.n42 0.155672
R727 VDD1.n42 VDD1.n18 0.155672
R728 VDD1.n35 VDD1.n18 0.155672
R729 VDD1.n35 VDD1.n34 0.155672
R730 VDD1.n34 VDD1.n22 0.155672
R731 VDD1.n27 VDD1.n22 0.155672
R732 VDD1.n103 VDD1.n98 0.155672
R733 VDD1.n110 VDD1.n98 0.155672
R734 VDD1.n111 VDD1.n110 0.155672
R735 VDD1.n111 VDD1.n94 0.155672
R736 VDD1.n118 VDD1.n94 0.155672
R737 VDD1.n119 VDD1.n118 0.155672
R738 VDD1.n119 VDD1.n90 0.155672
R739 VDD1.n128 VDD1.n90 0.155672
R740 VDD1.n129 VDD1.n128 0.155672
R741 VDD1.n129 VDD1.n86 0.155672
R742 VDD1.n136 VDD1.n86 0.155672
R743 VDD1.n137 VDD1.n136 0.155672
R744 VDD1.n137 VDD1.n82 0.155672
R745 VDD1.n144 VDD1.n82 0.155672
R746 VDD1.n145 VDD1.n144 0.155672
R747 VDD1.n145 VDD1.n78 0.155672
R748 VDD1.n152 VDD1.n78 0.155672
R749 VDD1 VDD1.n157 0.0910172
R750 B.n108 B.t9 1164.38
R751 B.n116 B.t6 1164.38
R752 B.n34 B.t0 1164.38
R753 B.n42 B.t3 1164.38
R754 B.n382 B.n67 585
R755 B.n384 B.n383 585
R756 B.n385 B.n66 585
R757 B.n387 B.n386 585
R758 B.n388 B.n65 585
R759 B.n390 B.n389 585
R760 B.n391 B.n64 585
R761 B.n393 B.n392 585
R762 B.n394 B.n63 585
R763 B.n396 B.n395 585
R764 B.n397 B.n62 585
R765 B.n399 B.n398 585
R766 B.n400 B.n61 585
R767 B.n402 B.n401 585
R768 B.n403 B.n60 585
R769 B.n405 B.n404 585
R770 B.n406 B.n59 585
R771 B.n408 B.n407 585
R772 B.n409 B.n58 585
R773 B.n411 B.n410 585
R774 B.n412 B.n57 585
R775 B.n414 B.n413 585
R776 B.n415 B.n56 585
R777 B.n417 B.n416 585
R778 B.n418 B.n55 585
R779 B.n420 B.n419 585
R780 B.n421 B.n54 585
R781 B.n423 B.n422 585
R782 B.n424 B.n53 585
R783 B.n426 B.n425 585
R784 B.n427 B.n52 585
R785 B.n429 B.n428 585
R786 B.n430 B.n51 585
R787 B.n432 B.n431 585
R788 B.n433 B.n50 585
R789 B.n435 B.n434 585
R790 B.n436 B.n49 585
R791 B.n438 B.n437 585
R792 B.n439 B.n48 585
R793 B.n441 B.n440 585
R794 B.n442 B.n47 585
R795 B.n444 B.n443 585
R796 B.n445 B.n46 585
R797 B.n447 B.n446 585
R798 B.n448 B.n45 585
R799 B.n450 B.n449 585
R800 B.n451 B.n44 585
R801 B.n453 B.n452 585
R802 B.n455 B.n41 585
R803 B.n457 B.n456 585
R804 B.n458 B.n40 585
R805 B.n460 B.n459 585
R806 B.n461 B.n39 585
R807 B.n463 B.n462 585
R808 B.n464 B.n38 585
R809 B.n466 B.n465 585
R810 B.n467 B.n37 585
R811 B.n469 B.n468 585
R812 B.n471 B.n470 585
R813 B.n472 B.n33 585
R814 B.n474 B.n473 585
R815 B.n475 B.n32 585
R816 B.n477 B.n476 585
R817 B.n478 B.n31 585
R818 B.n480 B.n479 585
R819 B.n481 B.n30 585
R820 B.n483 B.n482 585
R821 B.n484 B.n29 585
R822 B.n486 B.n485 585
R823 B.n487 B.n28 585
R824 B.n489 B.n488 585
R825 B.n490 B.n27 585
R826 B.n492 B.n491 585
R827 B.n493 B.n26 585
R828 B.n495 B.n494 585
R829 B.n496 B.n25 585
R830 B.n498 B.n497 585
R831 B.n499 B.n24 585
R832 B.n501 B.n500 585
R833 B.n502 B.n23 585
R834 B.n504 B.n503 585
R835 B.n505 B.n22 585
R836 B.n507 B.n506 585
R837 B.n508 B.n21 585
R838 B.n510 B.n509 585
R839 B.n511 B.n20 585
R840 B.n513 B.n512 585
R841 B.n514 B.n19 585
R842 B.n516 B.n515 585
R843 B.n517 B.n18 585
R844 B.n519 B.n518 585
R845 B.n520 B.n17 585
R846 B.n522 B.n521 585
R847 B.n523 B.n16 585
R848 B.n525 B.n524 585
R849 B.n526 B.n15 585
R850 B.n528 B.n527 585
R851 B.n529 B.n14 585
R852 B.n531 B.n530 585
R853 B.n532 B.n13 585
R854 B.n534 B.n533 585
R855 B.n535 B.n12 585
R856 B.n537 B.n536 585
R857 B.n538 B.n11 585
R858 B.n540 B.n539 585
R859 B.n541 B.n10 585
R860 B.n381 B.n380 585
R861 B.n379 B.n68 585
R862 B.n378 B.n377 585
R863 B.n376 B.n69 585
R864 B.n375 B.n374 585
R865 B.n373 B.n70 585
R866 B.n372 B.n371 585
R867 B.n370 B.n71 585
R868 B.n369 B.n368 585
R869 B.n367 B.n72 585
R870 B.n366 B.n365 585
R871 B.n364 B.n73 585
R872 B.n363 B.n362 585
R873 B.n361 B.n74 585
R874 B.n360 B.n359 585
R875 B.n358 B.n75 585
R876 B.n357 B.n356 585
R877 B.n355 B.n76 585
R878 B.n354 B.n353 585
R879 B.n352 B.n77 585
R880 B.n351 B.n350 585
R881 B.n349 B.n78 585
R882 B.n348 B.n347 585
R883 B.n346 B.n79 585
R884 B.n345 B.n344 585
R885 B.n343 B.n80 585
R886 B.n342 B.n341 585
R887 B.n340 B.n81 585
R888 B.n339 B.n338 585
R889 B.n337 B.n82 585
R890 B.n336 B.n335 585
R891 B.n334 B.n83 585
R892 B.n333 B.n332 585
R893 B.n172 B.n141 585
R894 B.n174 B.n173 585
R895 B.n175 B.n140 585
R896 B.n177 B.n176 585
R897 B.n178 B.n139 585
R898 B.n180 B.n179 585
R899 B.n181 B.n138 585
R900 B.n183 B.n182 585
R901 B.n184 B.n137 585
R902 B.n186 B.n185 585
R903 B.n187 B.n136 585
R904 B.n189 B.n188 585
R905 B.n190 B.n135 585
R906 B.n192 B.n191 585
R907 B.n193 B.n134 585
R908 B.n195 B.n194 585
R909 B.n196 B.n133 585
R910 B.n198 B.n197 585
R911 B.n199 B.n132 585
R912 B.n201 B.n200 585
R913 B.n202 B.n131 585
R914 B.n204 B.n203 585
R915 B.n205 B.n130 585
R916 B.n207 B.n206 585
R917 B.n208 B.n129 585
R918 B.n210 B.n209 585
R919 B.n211 B.n128 585
R920 B.n213 B.n212 585
R921 B.n214 B.n127 585
R922 B.n216 B.n215 585
R923 B.n217 B.n126 585
R924 B.n219 B.n218 585
R925 B.n220 B.n125 585
R926 B.n222 B.n221 585
R927 B.n223 B.n124 585
R928 B.n225 B.n224 585
R929 B.n226 B.n123 585
R930 B.n228 B.n227 585
R931 B.n229 B.n122 585
R932 B.n231 B.n230 585
R933 B.n232 B.n121 585
R934 B.n234 B.n233 585
R935 B.n235 B.n120 585
R936 B.n237 B.n236 585
R937 B.n238 B.n119 585
R938 B.n240 B.n239 585
R939 B.n241 B.n118 585
R940 B.n243 B.n242 585
R941 B.n245 B.n115 585
R942 B.n247 B.n246 585
R943 B.n248 B.n114 585
R944 B.n250 B.n249 585
R945 B.n251 B.n113 585
R946 B.n253 B.n252 585
R947 B.n254 B.n112 585
R948 B.n256 B.n255 585
R949 B.n257 B.n111 585
R950 B.n259 B.n258 585
R951 B.n261 B.n260 585
R952 B.n262 B.n107 585
R953 B.n264 B.n263 585
R954 B.n265 B.n106 585
R955 B.n267 B.n266 585
R956 B.n268 B.n105 585
R957 B.n270 B.n269 585
R958 B.n271 B.n104 585
R959 B.n273 B.n272 585
R960 B.n274 B.n103 585
R961 B.n276 B.n275 585
R962 B.n277 B.n102 585
R963 B.n279 B.n278 585
R964 B.n280 B.n101 585
R965 B.n282 B.n281 585
R966 B.n283 B.n100 585
R967 B.n285 B.n284 585
R968 B.n286 B.n99 585
R969 B.n288 B.n287 585
R970 B.n289 B.n98 585
R971 B.n291 B.n290 585
R972 B.n292 B.n97 585
R973 B.n294 B.n293 585
R974 B.n295 B.n96 585
R975 B.n297 B.n296 585
R976 B.n298 B.n95 585
R977 B.n300 B.n299 585
R978 B.n301 B.n94 585
R979 B.n303 B.n302 585
R980 B.n304 B.n93 585
R981 B.n306 B.n305 585
R982 B.n307 B.n92 585
R983 B.n309 B.n308 585
R984 B.n310 B.n91 585
R985 B.n312 B.n311 585
R986 B.n313 B.n90 585
R987 B.n315 B.n314 585
R988 B.n316 B.n89 585
R989 B.n318 B.n317 585
R990 B.n319 B.n88 585
R991 B.n321 B.n320 585
R992 B.n322 B.n87 585
R993 B.n324 B.n323 585
R994 B.n325 B.n86 585
R995 B.n327 B.n326 585
R996 B.n328 B.n85 585
R997 B.n330 B.n329 585
R998 B.n331 B.n84 585
R999 B.n171 B.n170 585
R1000 B.n169 B.n142 585
R1001 B.n168 B.n167 585
R1002 B.n166 B.n143 585
R1003 B.n165 B.n164 585
R1004 B.n163 B.n144 585
R1005 B.n162 B.n161 585
R1006 B.n160 B.n145 585
R1007 B.n159 B.n158 585
R1008 B.n157 B.n146 585
R1009 B.n156 B.n155 585
R1010 B.n154 B.n147 585
R1011 B.n153 B.n152 585
R1012 B.n151 B.n148 585
R1013 B.n150 B.n149 585
R1014 B.n2 B.n0 585
R1015 B.n565 B.n1 585
R1016 B.n564 B.n563 585
R1017 B.n562 B.n3 585
R1018 B.n561 B.n560 585
R1019 B.n559 B.n4 585
R1020 B.n558 B.n557 585
R1021 B.n556 B.n5 585
R1022 B.n555 B.n554 585
R1023 B.n553 B.n6 585
R1024 B.n552 B.n551 585
R1025 B.n550 B.n7 585
R1026 B.n549 B.n548 585
R1027 B.n547 B.n8 585
R1028 B.n546 B.n545 585
R1029 B.n544 B.n9 585
R1030 B.n543 B.n542 585
R1031 B.n567 B.n566 585
R1032 B.n170 B.n141 535.745
R1033 B.n542 B.n541 535.745
R1034 B.n332 B.n331 535.745
R1035 B.n380 B.n67 535.745
R1036 B.n108 B.t11 429.533
R1037 B.n42 B.t4 429.533
R1038 B.n116 B.t8 429.533
R1039 B.n34 B.t1 429.533
R1040 B.n109 B.t10 416.151
R1041 B.n43 B.t5 416.151
R1042 B.n117 B.t7 416.151
R1043 B.n35 B.t2 416.151
R1044 B.n170 B.n169 163.367
R1045 B.n169 B.n168 163.367
R1046 B.n168 B.n143 163.367
R1047 B.n164 B.n143 163.367
R1048 B.n164 B.n163 163.367
R1049 B.n163 B.n162 163.367
R1050 B.n162 B.n145 163.367
R1051 B.n158 B.n145 163.367
R1052 B.n158 B.n157 163.367
R1053 B.n157 B.n156 163.367
R1054 B.n156 B.n147 163.367
R1055 B.n152 B.n147 163.367
R1056 B.n152 B.n151 163.367
R1057 B.n151 B.n150 163.367
R1058 B.n150 B.n2 163.367
R1059 B.n566 B.n2 163.367
R1060 B.n566 B.n565 163.367
R1061 B.n565 B.n564 163.367
R1062 B.n564 B.n3 163.367
R1063 B.n560 B.n3 163.367
R1064 B.n560 B.n559 163.367
R1065 B.n559 B.n558 163.367
R1066 B.n558 B.n5 163.367
R1067 B.n554 B.n5 163.367
R1068 B.n554 B.n553 163.367
R1069 B.n553 B.n552 163.367
R1070 B.n552 B.n7 163.367
R1071 B.n548 B.n7 163.367
R1072 B.n548 B.n547 163.367
R1073 B.n547 B.n546 163.367
R1074 B.n546 B.n9 163.367
R1075 B.n542 B.n9 163.367
R1076 B.n174 B.n141 163.367
R1077 B.n175 B.n174 163.367
R1078 B.n176 B.n175 163.367
R1079 B.n176 B.n139 163.367
R1080 B.n180 B.n139 163.367
R1081 B.n181 B.n180 163.367
R1082 B.n182 B.n181 163.367
R1083 B.n182 B.n137 163.367
R1084 B.n186 B.n137 163.367
R1085 B.n187 B.n186 163.367
R1086 B.n188 B.n187 163.367
R1087 B.n188 B.n135 163.367
R1088 B.n192 B.n135 163.367
R1089 B.n193 B.n192 163.367
R1090 B.n194 B.n193 163.367
R1091 B.n194 B.n133 163.367
R1092 B.n198 B.n133 163.367
R1093 B.n199 B.n198 163.367
R1094 B.n200 B.n199 163.367
R1095 B.n200 B.n131 163.367
R1096 B.n204 B.n131 163.367
R1097 B.n205 B.n204 163.367
R1098 B.n206 B.n205 163.367
R1099 B.n206 B.n129 163.367
R1100 B.n210 B.n129 163.367
R1101 B.n211 B.n210 163.367
R1102 B.n212 B.n211 163.367
R1103 B.n212 B.n127 163.367
R1104 B.n216 B.n127 163.367
R1105 B.n217 B.n216 163.367
R1106 B.n218 B.n217 163.367
R1107 B.n218 B.n125 163.367
R1108 B.n222 B.n125 163.367
R1109 B.n223 B.n222 163.367
R1110 B.n224 B.n223 163.367
R1111 B.n224 B.n123 163.367
R1112 B.n228 B.n123 163.367
R1113 B.n229 B.n228 163.367
R1114 B.n230 B.n229 163.367
R1115 B.n230 B.n121 163.367
R1116 B.n234 B.n121 163.367
R1117 B.n235 B.n234 163.367
R1118 B.n236 B.n235 163.367
R1119 B.n236 B.n119 163.367
R1120 B.n240 B.n119 163.367
R1121 B.n241 B.n240 163.367
R1122 B.n242 B.n241 163.367
R1123 B.n242 B.n115 163.367
R1124 B.n247 B.n115 163.367
R1125 B.n248 B.n247 163.367
R1126 B.n249 B.n248 163.367
R1127 B.n249 B.n113 163.367
R1128 B.n253 B.n113 163.367
R1129 B.n254 B.n253 163.367
R1130 B.n255 B.n254 163.367
R1131 B.n255 B.n111 163.367
R1132 B.n259 B.n111 163.367
R1133 B.n260 B.n259 163.367
R1134 B.n260 B.n107 163.367
R1135 B.n264 B.n107 163.367
R1136 B.n265 B.n264 163.367
R1137 B.n266 B.n265 163.367
R1138 B.n266 B.n105 163.367
R1139 B.n270 B.n105 163.367
R1140 B.n271 B.n270 163.367
R1141 B.n272 B.n271 163.367
R1142 B.n272 B.n103 163.367
R1143 B.n276 B.n103 163.367
R1144 B.n277 B.n276 163.367
R1145 B.n278 B.n277 163.367
R1146 B.n278 B.n101 163.367
R1147 B.n282 B.n101 163.367
R1148 B.n283 B.n282 163.367
R1149 B.n284 B.n283 163.367
R1150 B.n284 B.n99 163.367
R1151 B.n288 B.n99 163.367
R1152 B.n289 B.n288 163.367
R1153 B.n290 B.n289 163.367
R1154 B.n290 B.n97 163.367
R1155 B.n294 B.n97 163.367
R1156 B.n295 B.n294 163.367
R1157 B.n296 B.n295 163.367
R1158 B.n296 B.n95 163.367
R1159 B.n300 B.n95 163.367
R1160 B.n301 B.n300 163.367
R1161 B.n302 B.n301 163.367
R1162 B.n302 B.n93 163.367
R1163 B.n306 B.n93 163.367
R1164 B.n307 B.n306 163.367
R1165 B.n308 B.n307 163.367
R1166 B.n308 B.n91 163.367
R1167 B.n312 B.n91 163.367
R1168 B.n313 B.n312 163.367
R1169 B.n314 B.n313 163.367
R1170 B.n314 B.n89 163.367
R1171 B.n318 B.n89 163.367
R1172 B.n319 B.n318 163.367
R1173 B.n320 B.n319 163.367
R1174 B.n320 B.n87 163.367
R1175 B.n324 B.n87 163.367
R1176 B.n325 B.n324 163.367
R1177 B.n326 B.n325 163.367
R1178 B.n326 B.n85 163.367
R1179 B.n330 B.n85 163.367
R1180 B.n331 B.n330 163.367
R1181 B.n332 B.n83 163.367
R1182 B.n336 B.n83 163.367
R1183 B.n337 B.n336 163.367
R1184 B.n338 B.n337 163.367
R1185 B.n338 B.n81 163.367
R1186 B.n342 B.n81 163.367
R1187 B.n343 B.n342 163.367
R1188 B.n344 B.n343 163.367
R1189 B.n344 B.n79 163.367
R1190 B.n348 B.n79 163.367
R1191 B.n349 B.n348 163.367
R1192 B.n350 B.n349 163.367
R1193 B.n350 B.n77 163.367
R1194 B.n354 B.n77 163.367
R1195 B.n355 B.n354 163.367
R1196 B.n356 B.n355 163.367
R1197 B.n356 B.n75 163.367
R1198 B.n360 B.n75 163.367
R1199 B.n361 B.n360 163.367
R1200 B.n362 B.n361 163.367
R1201 B.n362 B.n73 163.367
R1202 B.n366 B.n73 163.367
R1203 B.n367 B.n366 163.367
R1204 B.n368 B.n367 163.367
R1205 B.n368 B.n71 163.367
R1206 B.n372 B.n71 163.367
R1207 B.n373 B.n372 163.367
R1208 B.n374 B.n373 163.367
R1209 B.n374 B.n69 163.367
R1210 B.n378 B.n69 163.367
R1211 B.n379 B.n378 163.367
R1212 B.n380 B.n379 163.367
R1213 B.n541 B.n540 163.367
R1214 B.n540 B.n11 163.367
R1215 B.n536 B.n11 163.367
R1216 B.n536 B.n535 163.367
R1217 B.n535 B.n534 163.367
R1218 B.n534 B.n13 163.367
R1219 B.n530 B.n13 163.367
R1220 B.n530 B.n529 163.367
R1221 B.n529 B.n528 163.367
R1222 B.n528 B.n15 163.367
R1223 B.n524 B.n15 163.367
R1224 B.n524 B.n523 163.367
R1225 B.n523 B.n522 163.367
R1226 B.n522 B.n17 163.367
R1227 B.n518 B.n17 163.367
R1228 B.n518 B.n517 163.367
R1229 B.n517 B.n516 163.367
R1230 B.n516 B.n19 163.367
R1231 B.n512 B.n19 163.367
R1232 B.n512 B.n511 163.367
R1233 B.n511 B.n510 163.367
R1234 B.n510 B.n21 163.367
R1235 B.n506 B.n21 163.367
R1236 B.n506 B.n505 163.367
R1237 B.n505 B.n504 163.367
R1238 B.n504 B.n23 163.367
R1239 B.n500 B.n23 163.367
R1240 B.n500 B.n499 163.367
R1241 B.n499 B.n498 163.367
R1242 B.n498 B.n25 163.367
R1243 B.n494 B.n25 163.367
R1244 B.n494 B.n493 163.367
R1245 B.n493 B.n492 163.367
R1246 B.n492 B.n27 163.367
R1247 B.n488 B.n27 163.367
R1248 B.n488 B.n487 163.367
R1249 B.n487 B.n486 163.367
R1250 B.n486 B.n29 163.367
R1251 B.n482 B.n29 163.367
R1252 B.n482 B.n481 163.367
R1253 B.n481 B.n480 163.367
R1254 B.n480 B.n31 163.367
R1255 B.n476 B.n31 163.367
R1256 B.n476 B.n475 163.367
R1257 B.n475 B.n474 163.367
R1258 B.n474 B.n33 163.367
R1259 B.n470 B.n33 163.367
R1260 B.n470 B.n469 163.367
R1261 B.n469 B.n37 163.367
R1262 B.n465 B.n37 163.367
R1263 B.n465 B.n464 163.367
R1264 B.n464 B.n463 163.367
R1265 B.n463 B.n39 163.367
R1266 B.n459 B.n39 163.367
R1267 B.n459 B.n458 163.367
R1268 B.n458 B.n457 163.367
R1269 B.n457 B.n41 163.367
R1270 B.n452 B.n41 163.367
R1271 B.n452 B.n451 163.367
R1272 B.n451 B.n450 163.367
R1273 B.n450 B.n45 163.367
R1274 B.n446 B.n45 163.367
R1275 B.n446 B.n445 163.367
R1276 B.n445 B.n444 163.367
R1277 B.n444 B.n47 163.367
R1278 B.n440 B.n47 163.367
R1279 B.n440 B.n439 163.367
R1280 B.n439 B.n438 163.367
R1281 B.n438 B.n49 163.367
R1282 B.n434 B.n49 163.367
R1283 B.n434 B.n433 163.367
R1284 B.n433 B.n432 163.367
R1285 B.n432 B.n51 163.367
R1286 B.n428 B.n51 163.367
R1287 B.n428 B.n427 163.367
R1288 B.n427 B.n426 163.367
R1289 B.n426 B.n53 163.367
R1290 B.n422 B.n53 163.367
R1291 B.n422 B.n421 163.367
R1292 B.n421 B.n420 163.367
R1293 B.n420 B.n55 163.367
R1294 B.n416 B.n55 163.367
R1295 B.n416 B.n415 163.367
R1296 B.n415 B.n414 163.367
R1297 B.n414 B.n57 163.367
R1298 B.n410 B.n57 163.367
R1299 B.n410 B.n409 163.367
R1300 B.n409 B.n408 163.367
R1301 B.n408 B.n59 163.367
R1302 B.n404 B.n59 163.367
R1303 B.n404 B.n403 163.367
R1304 B.n403 B.n402 163.367
R1305 B.n402 B.n61 163.367
R1306 B.n398 B.n61 163.367
R1307 B.n398 B.n397 163.367
R1308 B.n397 B.n396 163.367
R1309 B.n396 B.n63 163.367
R1310 B.n392 B.n63 163.367
R1311 B.n392 B.n391 163.367
R1312 B.n391 B.n390 163.367
R1313 B.n390 B.n65 163.367
R1314 B.n386 B.n65 163.367
R1315 B.n386 B.n385 163.367
R1316 B.n385 B.n384 163.367
R1317 B.n384 B.n67 163.367
R1318 B.n110 B.n109 59.5399
R1319 B.n244 B.n117 59.5399
R1320 B.n36 B.n35 59.5399
R1321 B.n454 B.n43 59.5399
R1322 B.n543 B.n10 34.8103
R1323 B.n382 B.n381 34.8103
R1324 B.n333 B.n84 34.8103
R1325 B.n172 B.n171 34.8103
R1326 B B.n567 18.0485
R1327 B.n109 B.n108 13.3823
R1328 B.n117 B.n116 13.3823
R1329 B.n35 B.n34 13.3823
R1330 B.n43 B.n42 13.3823
R1331 B.n539 B.n10 10.6151
R1332 B.n539 B.n538 10.6151
R1333 B.n538 B.n537 10.6151
R1334 B.n537 B.n12 10.6151
R1335 B.n533 B.n12 10.6151
R1336 B.n533 B.n532 10.6151
R1337 B.n532 B.n531 10.6151
R1338 B.n531 B.n14 10.6151
R1339 B.n527 B.n14 10.6151
R1340 B.n527 B.n526 10.6151
R1341 B.n526 B.n525 10.6151
R1342 B.n525 B.n16 10.6151
R1343 B.n521 B.n16 10.6151
R1344 B.n521 B.n520 10.6151
R1345 B.n520 B.n519 10.6151
R1346 B.n519 B.n18 10.6151
R1347 B.n515 B.n18 10.6151
R1348 B.n515 B.n514 10.6151
R1349 B.n514 B.n513 10.6151
R1350 B.n513 B.n20 10.6151
R1351 B.n509 B.n20 10.6151
R1352 B.n509 B.n508 10.6151
R1353 B.n508 B.n507 10.6151
R1354 B.n507 B.n22 10.6151
R1355 B.n503 B.n22 10.6151
R1356 B.n503 B.n502 10.6151
R1357 B.n502 B.n501 10.6151
R1358 B.n501 B.n24 10.6151
R1359 B.n497 B.n24 10.6151
R1360 B.n497 B.n496 10.6151
R1361 B.n496 B.n495 10.6151
R1362 B.n495 B.n26 10.6151
R1363 B.n491 B.n26 10.6151
R1364 B.n491 B.n490 10.6151
R1365 B.n490 B.n489 10.6151
R1366 B.n489 B.n28 10.6151
R1367 B.n485 B.n28 10.6151
R1368 B.n485 B.n484 10.6151
R1369 B.n484 B.n483 10.6151
R1370 B.n483 B.n30 10.6151
R1371 B.n479 B.n30 10.6151
R1372 B.n479 B.n478 10.6151
R1373 B.n478 B.n477 10.6151
R1374 B.n477 B.n32 10.6151
R1375 B.n473 B.n32 10.6151
R1376 B.n473 B.n472 10.6151
R1377 B.n472 B.n471 10.6151
R1378 B.n468 B.n467 10.6151
R1379 B.n467 B.n466 10.6151
R1380 B.n466 B.n38 10.6151
R1381 B.n462 B.n38 10.6151
R1382 B.n462 B.n461 10.6151
R1383 B.n461 B.n460 10.6151
R1384 B.n460 B.n40 10.6151
R1385 B.n456 B.n40 10.6151
R1386 B.n456 B.n455 10.6151
R1387 B.n453 B.n44 10.6151
R1388 B.n449 B.n44 10.6151
R1389 B.n449 B.n448 10.6151
R1390 B.n448 B.n447 10.6151
R1391 B.n447 B.n46 10.6151
R1392 B.n443 B.n46 10.6151
R1393 B.n443 B.n442 10.6151
R1394 B.n442 B.n441 10.6151
R1395 B.n441 B.n48 10.6151
R1396 B.n437 B.n48 10.6151
R1397 B.n437 B.n436 10.6151
R1398 B.n436 B.n435 10.6151
R1399 B.n435 B.n50 10.6151
R1400 B.n431 B.n50 10.6151
R1401 B.n431 B.n430 10.6151
R1402 B.n430 B.n429 10.6151
R1403 B.n429 B.n52 10.6151
R1404 B.n425 B.n52 10.6151
R1405 B.n425 B.n424 10.6151
R1406 B.n424 B.n423 10.6151
R1407 B.n423 B.n54 10.6151
R1408 B.n419 B.n54 10.6151
R1409 B.n419 B.n418 10.6151
R1410 B.n418 B.n417 10.6151
R1411 B.n417 B.n56 10.6151
R1412 B.n413 B.n56 10.6151
R1413 B.n413 B.n412 10.6151
R1414 B.n412 B.n411 10.6151
R1415 B.n411 B.n58 10.6151
R1416 B.n407 B.n58 10.6151
R1417 B.n407 B.n406 10.6151
R1418 B.n406 B.n405 10.6151
R1419 B.n405 B.n60 10.6151
R1420 B.n401 B.n60 10.6151
R1421 B.n401 B.n400 10.6151
R1422 B.n400 B.n399 10.6151
R1423 B.n399 B.n62 10.6151
R1424 B.n395 B.n62 10.6151
R1425 B.n395 B.n394 10.6151
R1426 B.n394 B.n393 10.6151
R1427 B.n393 B.n64 10.6151
R1428 B.n389 B.n64 10.6151
R1429 B.n389 B.n388 10.6151
R1430 B.n388 B.n387 10.6151
R1431 B.n387 B.n66 10.6151
R1432 B.n383 B.n66 10.6151
R1433 B.n383 B.n382 10.6151
R1434 B.n334 B.n333 10.6151
R1435 B.n335 B.n334 10.6151
R1436 B.n335 B.n82 10.6151
R1437 B.n339 B.n82 10.6151
R1438 B.n340 B.n339 10.6151
R1439 B.n341 B.n340 10.6151
R1440 B.n341 B.n80 10.6151
R1441 B.n345 B.n80 10.6151
R1442 B.n346 B.n345 10.6151
R1443 B.n347 B.n346 10.6151
R1444 B.n347 B.n78 10.6151
R1445 B.n351 B.n78 10.6151
R1446 B.n352 B.n351 10.6151
R1447 B.n353 B.n352 10.6151
R1448 B.n353 B.n76 10.6151
R1449 B.n357 B.n76 10.6151
R1450 B.n358 B.n357 10.6151
R1451 B.n359 B.n358 10.6151
R1452 B.n359 B.n74 10.6151
R1453 B.n363 B.n74 10.6151
R1454 B.n364 B.n363 10.6151
R1455 B.n365 B.n364 10.6151
R1456 B.n365 B.n72 10.6151
R1457 B.n369 B.n72 10.6151
R1458 B.n370 B.n369 10.6151
R1459 B.n371 B.n370 10.6151
R1460 B.n371 B.n70 10.6151
R1461 B.n375 B.n70 10.6151
R1462 B.n376 B.n375 10.6151
R1463 B.n377 B.n376 10.6151
R1464 B.n377 B.n68 10.6151
R1465 B.n381 B.n68 10.6151
R1466 B.n173 B.n172 10.6151
R1467 B.n173 B.n140 10.6151
R1468 B.n177 B.n140 10.6151
R1469 B.n178 B.n177 10.6151
R1470 B.n179 B.n178 10.6151
R1471 B.n179 B.n138 10.6151
R1472 B.n183 B.n138 10.6151
R1473 B.n184 B.n183 10.6151
R1474 B.n185 B.n184 10.6151
R1475 B.n185 B.n136 10.6151
R1476 B.n189 B.n136 10.6151
R1477 B.n190 B.n189 10.6151
R1478 B.n191 B.n190 10.6151
R1479 B.n191 B.n134 10.6151
R1480 B.n195 B.n134 10.6151
R1481 B.n196 B.n195 10.6151
R1482 B.n197 B.n196 10.6151
R1483 B.n197 B.n132 10.6151
R1484 B.n201 B.n132 10.6151
R1485 B.n202 B.n201 10.6151
R1486 B.n203 B.n202 10.6151
R1487 B.n203 B.n130 10.6151
R1488 B.n207 B.n130 10.6151
R1489 B.n208 B.n207 10.6151
R1490 B.n209 B.n208 10.6151
R1491 B.n209 B.n128 10.6151
R1492 B.n213 B.n128 10.6151
R1493 B.n214 B.n213 10.6151
R1494 B.n215 B.n214 10.6151
R1495 B.n215 B.n126 10.6151
R1496 B.n219 B.n126 10.6151
R1497 B.n220 B.n219 10.6151
R1498 B.n221 B.n220 10.6151
R1499 B.n221 B.n124 10.6151
R1500 B.n225 B.n124 10.6151
R1501 B.n226 B.n225 10.6151
R1502 B.n227 B.n226 10.6151
R1503 B.n227 B.n122 10.6151
R1504 B.n231 B.n122 10.6151
R1505 B.n232 B.n231 10.6151
R1506 B.n233 B.n232 10.6151
R1507 B.n233 B.n120 10.6151
R1508 B.n237 B.n120 10.6151
R1509 B.n238 B.n237 10.6151
R1510 B.n239 B.n238 10.6151
R1511 B.n239 B.n118 10.6151
R1512 B.n243 B.n118 10.6151
R1513 B.n246 B.n245 10.6151
R1514 B.n246 B.n114 10.6151
R1515 B.n250 B.n114 10.6151
R1516 B.n251 B.n250 10.6151
R1517 B.n252 B.n251 10.6151
R1518 B.n252 B.n112 10.6151
R1519 B.n256 B.n112 10.6151
R1520 B.n257 B.n256 10.6151
R1521 B.n258 B.n257 10.6151
R1522 B.n262 B.n261 10.6151
R1523 B.n263 B.n262 10.6151
R1524 B.n263 B.n106 10.6151
R1525 B.n267 B.n106 10.6151
R1526 B.n268 B.n267 10.6151
R1527 B.n269 B.n268 10.6151
R1528 B.n269 B.n104 10.6151
R1529 B.n273 B.n104 10.6151
R1530 B.n274 B.n273 10.6151
R1531 B.n275 B.n274 10.6151
R1532 B.n275 B.n102 10.6151
R1533 B.n279 B.n102 10.6151
R1534 B.n280 B.n279 10.6151
R1535 B.n281 B.n280 10.6151
R1536 B.n281 B.n100 10.6151
R1537 B.n285 B.n100 10.6151
R1538 B.n286 B.n285 10.6151
R1539 B.n287 B.n286 10.6151
R1540 B.n287 B.n98 10.6151
R1541 B.n291 B.n98 10.6151
R1542 B.n292 B.n291 10.6151
R1543 B.n293 B.n292 10.6151
R1544 B.n293 B.n96 10.6151
R1545 B.n297 B.n96 10.6151
R1546 B.n298 B.n297 10.6151
R1547 B.n299 B.n298 10.6151
R1548 B.n299 B.n94 10.6151
R1549 B.n303 B.n94 10.6151
R1550 B.n304 B.n303 10.6151
R1551 B.n305 B.n304 10.6151
R1552 B.n305 B.n92 10.6151
R1553 B.n309 B.n92 10.6151
R1554 B.n310 B.n309 10.6151
R1555 B.n311 B.n310 10.6151
R1556 B.n311 B.n90 10.6151
R1557 B.n315 B.n90 10.6151
R1558 B.n316 B.n315 10.6151
R1559 B.n317 B.n316 10.6151
R1560 B.n317 B.n88 10.6151
R1561 B.n321 B.n88 10.6151
R1562 B.n322 B.n321 10.6151
R1563 B.n323 B.n322 10.6151
R1564 B.n323 B.n86 10.6151
R1565 B.n327 B.n86 10.6151
R1566 B.n328 B.n327 10.6151
R1567 B.n329 B.n328 10.6151
R1568 B.n329 B.n84 10.6151
R1569 B.n171 B.n142 10.6151
R1570 B.n167 B.n142 10.6151
R1571 B.n167 B.n166 10.6151
R1572 B.n166 B.n165 10.6151
R1573 B.n165 B.n144 10.6151
R1574 B.n161 B.n144 10.6151
R1575 B.n161 B.n160 10.6151
R1576 B.n160 B.n159 10.6151
R1577 B.n159 B.n146 10.6151
R1578 B.n155 B.n146 10.6151
R1579 B.n155 B.n154 10.6151
R1580 B.n154 B.n153 10.6151
R1581 B.n153 B.n148 10.6151
R1582 B.n149 B.n148 10.6151
R1583 B.n149 B.n0 10.6151
R1584 B.n563 B.n1 10.6151
R1585 B.n563 B.n562 10.6151
R1586 B.n562 B.n561 10.6151
R1587 B.n561 B.n4 10.6151
R1588 B.n557 B.n4 10.6151
R1589 B.n557 B.n556 10.6151
R1590 B.n556 B.n555 10.6151
R1591 B.n555 B.n6 10.6151
R1592 B.n551 B.n6 10.6151
R1593 B.n551 B.n550 10.6151
R1594 B.n550 B.n549 10.6151
R1595 B.n549 B.n8 10.6151
R1596 B.n545 B.n8 10.6151
R1597 B.n545 B.n544 10.6151
R1598 B.n544 B.n543 10.6151
R1599 B.n471 B.n36 9.36635
R1600 B.n454 B.n453 9.36635
R1601 B.n244 B.n243 9.36635
R1602 B.n261 B.n110 9.36635
R1603 B.n567 B.n0 2.81026
R1604 B.n567 B.n1 2.81026
R1605 B.n468 B.n36 1.24928
R1606 B.n455 B.n454 1.24928
R1607 B.n245 B.n244 1.24928
R1608 B.n258 B.n110 1.24928
R1609 VN.n0 VN.t0 1085.63
R1610 VN.n4 VN.t2 1085.63
R1611 VN.n2 VN.t3 1065.21
R1612 VN.n6 VN.t1 1065.21
R1613 VN.n1 VN.t5 1063.75
R1614 VN.n5 VN.t4 1063.75
R1615 VN.n3 VN.n2 161.3
R1616 VN.n7 VN.n6 161.3
R1617 VN.n7 VN.n4 70.6808
R1618 VN.n3 VN.n0 70.6808
R1619 VN.n2 VN.n1 46.7399
R1620 VN.n6 VN.n5 46.7399
R1621 VN VN.n7 41.9835
R1622 VN.n5 VN.n4 20.4028
R1623 VN.n1 VN.n0 20.4028
R1624 VN VN.n3 0.0516364
R1625 VDD2.n151 VDD2.n79 756.745
R1626 VDD2.n72 VDD2.n0 756.745
R1627 VDD2.n152 VDD2.n151 585
R1628 VDD2.n150 VDD2.n149 585
R1629 VDD2.n83 VDD2.n82 585
R1630 VDD2.n144 VDD2.n143 585
R1631 VDD2.n142 VDD2.n141 585
R1632 VDD2.n87 VDD2.n86 585
R1633 VDD2.n136 VDD2.n135 585
R1634 VDD2.n134 VDD2.n133 585
R1635 VDD2.n91 VDD2.n90 585
R1636 VDD2.n128 VDD2.n127 585
R1637 VDD2.n126 VDD2.n93 585
R1638 VDD2.n125 VDD2.n124 585
R1639 VDD2.n96 VDD2.n94 585
R1640 VDD2.n119 VDD2.n118 585
R1641 VDD2.n117 VDD2.n116 585
R1642 VDD2.n100 VDD2.n99 585
R1643 VDD2.n111 VDD2.n110 585
R1644 VDD2.n109 VDD2.n108 585
R1645 VDD2.n104 VDD2.n103 585
R1646 VDD2.n24 VDD2.n23 585
R1647 VDD2.n29 VDD2.n28 585
R1648 VDD2.n31 VDD2.n30 585
R1649 VDD2.n20 VDD2.n19 585
R1650 VDD2.n37 VDD2.n36 585
R1651 VDD2.n39 VDD2.n38 585
R1652 VDD2.n16 VDD2.n15 585
R1653 VDD2.n46 VDD2.n45 585
R1654 VDD2.n47 VDD2.n14 585
R1655 VDD2.n49 VDD2.n48 585
R1656 VDD2.n12 VDD2.n11 585
R1657 VDD2.n55 VDD2.n54 585
R1658 VDD2.n57 VDD2.n56 585
R1659 VDD2.n8 VDD2.n7 585
R1660 VDD2.n63 VDD2.n62 585
R1661 VDD2.n65 VDD2.n64 585
R1662 VDD2.n4 VDD2.n3 585
R1663 VDD2.n71 VDD2.n70 585
R1664 VDD2.n73 VDD2.n72 585
R1665 VDD2.n105 VDD2.t4 329.036
R1666 VDD2.n25 VDD2.t5 329.036
R1667 VDD2.n151 VDD2.n150 171.744
R1668 VDD2.n150 VDD2.n82 171.744
R1669 VDD2.n143 VDD2.n82 171.744
R1670 VDD2.n143 VDD2.n142 171.744
R1671 VDD2.n142 VDD2.n86 171.744
R1672 VDD2.n135 VDD2.n86 171.744
R1673 VDD2.n135 VDD2.n134 171.744
R1674 VDD2.n134 VDD2.n90 171.744
R1675 VDD2.n127 VDD2.n90 171.744
R1676 VDD2.n127 VDD2.n126 171.744
R1677 VDD2.n126 VDD2.n125 171.744
R1678 VDD2.n125 VDD2.n94 171.744
R1679 VDD2.n118 VDD2.n94 171.744
R1680 VDD2.n118 VDD2.n117 171.744
R1681 VDD2.n117 VDD2.n99 171.744
R1682 VDD2.n110 VDD2.n99 171.744
R1683 VDD2.n110 VDD2.n109 171.744
R1684 VDD2.n109 VDD2.n103 171.744
R1685 VDD2.n29 VDD2.n23 171.744
R1686 VDD2.n30 VDD2.n29 171.744
R1687 VDD2.n30 VDD2.n19 171.744
R1688 VDD2.n37 VDD2.n19 171.744
R1689 VDD2.n38 VDD2.n37 171.744
R1690 VDD2.n38 VDD2.n15 171.744
R1691 VDD2.n46 VDD2.n15 171.744
R1692 VDD2.n47 VDD2.n46 171.744
R1693 VDD2.n48 VDD2.n47 171.744
R1694 VDD2.n48 VDD2.n11 171.744
R1695 VDD2.n55 VDD2.n11 171.744
R1696 VDD2.n56 VDD2.n55 171.744
R1697 VDD2.n56 VDD2.n7 171.744
R1698 VDD2.n63 VDD2.n7 171.744
R1699 VDD2.n64 VDD2.n63 171.744
R1700 VDD2.n64 VDD2.n3 171.744
R1701 VDD2.n71 VDD2.n3 171.744
R1702 VDD2.n72 VDD2.n71 171.744
R1703 VDD2.t4 VDD2.n103 85.8723
R1704 VDD2.t5 VDD2.n23 85.8723
R1705 VDD2.n78 VDD2.n77 70.9506
R1706 VDD2 VDD2.n157 70.9477
R1707 VDD2.n78 VDD2.n76 48.4792
R1708 VDD2.n156 VDD2.n155 48.0884
R1709 VDD2.n156 VDD2.n78 37.9243
R1710 VDD2.n128 VDD2.n93 13.1884
R1711 VDD2.n49 VDD2.n14 13.1884
R1712 VDD2.n129 VDD2.n91 12.8005
R1713 VDD2.n124 VDD2.n95 12.8005
R1714 VDD2.n45 VDD2.n44 12.8005
R1715 VDD2.n50 VDD2.n12 12.8005
R1716 VDD2.n133 VDD2.n132 12.0247
R1717 VDD2.n123 VDD2.n96 12.0247
R1718 VDD2.n43 VDD2.n16 12.0247
R1719 VDD2.n54 VDD2.n53 12.0247
R1720 VDD2.n136 VDD2.n89 11.249
R1721 VDD2.n120 VDD2.n119 11.249
R1722 VDD2.n40 VDD2.n39 11.249
R1723 VDD2.n57 VDD2.n10 11.249
R1724 VDD2.n105 VDD2.n104 10.7239
R1725 VDD2.n25 VDD2.n24 10.7239
R1726 VDD2.n137 VDD2.n87 10.4732
R1727 VDD2.n116 VDD2.n98 10.4732
R1728 VDD2.n36 VDD2.n18 10.4732
R1729 VDD2.n58 VDD2.n8 10.4732
R1730 VDD2.n141 VDD2.n140 9.69747
R1731 VDD2.n115 VDD2.n100 9.69747
R1732 VDD2.n35 VDD2.n20 9.69747
R1733 VDD2.n62 VDD2.n61 9.69747
R1734 VDD2.n155 VDD2.n154 9.45567
R1735 VDD2.n76 VDD2.n75 9.45567
R1736 VDD2.n107 VDD2.n106 9.3005
R1737 VDD2.n102 VDD2.n101 9.3005
R1738 VDD2.n113 VDD2.n112 9.3005
R1739 VDD2.n115 VDD2.n114 9.3005
R1740 VDD2.n98 VDD2.n97 9.3005
R1741 VDD2.n121 VDD2.n120 9.3005
R1742 VDD2.n123 VDD2.n122 9.3005
R1743 VDD2.n95 VDD2.n92 9.3005
R1744 VDD2.n154 VDD2.n153 9.3005
R1745 VDD2.n81 VDD2.n80 9.3005
R1746 VDD2.n148 VDD2.n147 9.3005
R1747 VDD2.n146 VDD2.n145 9.3005
R1748 VDD2.n85 VDD2.n84 9.3005
R1749 VDD2.n140 VDD2.n139 9.3005
R1750 VDD2.n138 VDD2.n137 9.3005
R1751 VDD2.n89 VDD2.n88 9.3005
R1752 VDD2.n132 VDD2.n131 9.3005
R1753 VDD2.n130 VDD2.n129 9.3005
R1754 VDD2.n2 VDD2.n1 9.3005
R1755 VDD2.n75 VDD2.n74 9.3005
R1756 VDD2.n67 VDD2.n66 9.3005
R1757 VDD2.n6 VDD2.n5 9.3005
R1758 VDD2.n61 VDD2.n60 9.3005
R1759 VDD2.n59 VDD2.n58 9.3005
R1760 VDD2.n10 VDD2.n9 9.3005
R1761 VDD2.n53 VDD2.n52 9.3005
R1762 VDD2.n51 VDD2.n50 9.3005
R1763 VDD2.n27 VDD2.n26 9.3005
R1764 VDD2.n22 VDD2.n21 9.3005
R1765 VDD2.n33 VDD2.n32 9.3005
R1766 VDD2.n35 VDD2.n34 9.3005
R1767 VDD2.n18 VDD2.n17 9.3005
R1768 VDD2.n41 VDD2.n40 9.3005
R1769 VDD2.n43 VDD2.n42 9.3005
R1770 VDD2.n44 VDD2.n13 9.3005
R1771 VDD2.n69 VDD2.n68 9.3005
R1772 VDD2.n144 VDD2.n85 8.92171
R1773 VDD2.n112 VDD2.n111 8.92171
R1774 VDD2.n32 VDD2.n31 8.92171
R1775 VDD2.n65 VDD2.n6 8.92171
R1776 VDD2.n155 VDD2.n79 8.14595
R1777 VDD2.n145 VDD2.n83 8.14595
R1778 VDD2.n108 VDD2.n102 8.14595
R1779 VDD2.n28 VDD2.n22 8.14595
R1780 VDD2.n66 VDD2.n4 8.14595
R1781 VDD2.n76 VDD2.n0 8.14595
R1782 VDD2.n153 VDD2.n152 7.3702
R1783 VDD2.n149 VDD2.n148 7.3702
R1784 VDD2.n107 VDD2.n104 7.3702
R1785 VDD2.n27 VDD2.n24 7.3702
R1786 VDD2.n70 VDD2.n69 7.3702
R1787 VDD2.n74 VDD2.n73 7.3702
R1788 VDD2.n152 VDD2.n81 6.59444
R1789 VDD2.n149 VDD2.n81 6.59444
R1790 VDD2.n70 VDD2.n2 6.59444
R1791 VDD2.n73 VDD2.n2 6.59444
R1792 VDD2.n153 VDD2.n79 5.81868
R1793 VDD2.n148 VDD2.n83 5.81868
R1794 VDD2.n108 VDD2.n107 5.81868
R1795 VDD2.n28 VDD2.n27 5.81868
R1796 VDD2.n69 VDD2.n4 5.81868
R1797 VDD2.n74 VDD2.n0 5.81868
R1798 VDD2.n145 VDD2.n144 5.04292
R1799 VDD2.n111 VDD2.n102 5.04292
R1800 VDD2.n31 VDD2.n22 5.04292
R1801 VDD2.n66 VDD2.n65 5.04292
R1802 VDD2.n141 VDD2.n85 4.26717
R1803 VDD2.n112 VDD2.n100 4.26717
R1804 VDD2.n32 VDD2.n20 4.26717
R1805 VDD2.n62 VDD2.n6 4.26717
R1806 VDD2.n140 VDD2.n87 3.49141
R1807 VDD2.n116 VDD2.n115 3.49141
R1808 VDD2.n36 VDD2.n35 3.49141
R1809 VDD2.n61 VDD2.n8 3.49141
R1810 VDD2.n137 VDD2.n136 2.71565
R1811 VDD2.n119 VDD2.n98 2.71565
R1812 VDD2.n39 VDD2.n18 2.71565
R1813 VDD2.n58 VDD2.n57 2.71565
R1814 VDD2.n106 VDD2.n105 2.41282
R1815 VDD2.n26 VDD2.n25 2.41282
R1816 VDD2.n157 VDD2.t1 2.28315
R1817 VDD2.n157 VDD2.t3 2.28315
R1818 VDD2.n77 VDD2.t0 2.28315
R1819 VDD2.n77 VDD2.t2 2.28315
R1820 VDD2.n133 VDD2.n89 1.93989
R1821 VDD2.n120 VDD2.n96 1.93989
R1822 VDD2.n40 VDD2.n16 1.93989
R1823 VDD2.n54 VDD2.n10 1.93989
R1824 VDD2.n132 VDD2.n91 1.16414
R1825 VDD2.n124 VDD2.n123 1.16414
R1826 VDD2.n45 VDD2.n43 1.16414
R1827 VDD2.n53 VDD2.n12 1.16414
R1828 VDD2 VDD2.n156 0.50481
R1829 VDD2.n129 VDD2.n128 0.388379
R1830 VDD2.n95 VDD2.n93 0.388379
R1831 VDD2.n44 VDD2.n14 0.388379
R1832 VDD2.n50 VDD2.n49 0.388379
R1833 VDD2.n154 VDD2.n80 0.155672
R1834 VDD2.n147 VDD2.n80 0.155672
R1835 VDD2.n147 VDD2.n146 0.155672
R1836 VDD2.n146 VDD2.n84 0.155672
R1837 VDD2.n139 VDD2.n84 0.155672
R1838 VDD2.n139 VDD2.n138 0.155672
R1839 VDD2.n138 VDD2.n88 0.155672
R1840 VDD2.n131 VDD2.n88 0.155672
R1841 VDD2.n131 VDD2.n130 0.155672
R1842 VDD2.n130 VDD2.n92 0.155672
R1843 VDD2.n122 VDD2.n92 0.155672
R1844 VDD2.n122 VDD2.n121 0.155672
R1845 VDD2.n121 VDD2.n97 0.155672
R1846 VDD2.n114 VDD2.n97 0.155672
R1847 VDD2.n114 VDD2.n113 0.155672
R1848 VDD2.n113 VDD2.n101 0.155672
R1849 VDD2.n106 VDD2.n101 0.155672
R1850 VDD2.n26 VDD2.n21 0.155672
R1851 VDD2.n33 VDD2.n21 0.155672
R1852 VDD2.n34 VDD2.n33 0.155672
R1853 VDD2.n34 VDD2.n17 0.155672
R1854 VDD2.n41 VDD2.n17 0.155672
R1855 VDD2.n42 VDD2.n41 0.155672
R1856 VDD2.n42 VDD2.n13 0.155672
R1857 VDD2.n51 VDD2.n13 0.155672
R1858 VDD2.n52 VDD2.n51 0.155672
R1859 VDD2.n52 VDD2.n9 0.155672
R1860 VDD2.n59 VDD2.n9 0.155672
R1861 VDD2.n60 VDD2.n59 0.155672
R1862 VDD2.n60 VDD2.n5 0.155672
R1863 VDD2.n67 VDD2.n5 0.155672
R1864 VDD2.n68 VDD2.n67 0.155672
R1865 VDD2.n68 VDD2.n1 0.155672
R1866 VDD2.n75 VDD2.n1 0.155672
C0 VDD2 w_n1522_n3816# 1.89656f
C1 VN B 0.714378f
C2 VDD1 B 1.61f
C3 VTAIL w_n1522_n3816# 3.34929f
C4 VN VDD1 0.147371f
C5 VP VDD2 0.269079f
C6 w_n1522_n3816# B 7.21447f
C7 VN w_n1522_n3816# 2.38726f
C8 VTAIL VP 3.00414f
C9 VDD1 w_n1522_n3816# 1.88278f
C10 VTAIL VDD2 15.086301f
C11 VP B 1.02121f
C12 VDD2 B 1.63142f
C13 VN VP 5.16897f
C14 VN VDD2 3.52008f
C15 VDD1 VP 3.63587f
C16 VDD1 VDD2 0.591931f
C17 VTAIL B 2.83806f
C18 VN VTAIL 2.98929f
C19 VDD1 VTAIL 15.0575f
C20 VP w_n1522_n3816# 2.57779f
C21 VDD2 VSUBS 1.419973f
C22 VDD1 VSUBS 1.114718f
C23 VTAIL VSUBS 0.66604f
C24 VN VSUBS 4.64579f
C25 VP VSUBS 1.295179f
C26 B VSUBS 2.597827f
C27 w_n1522_n3816# VSUBS 71.28439f
C28 VDD2.n0 VSUBS 0.030124f
C29 VDD2.n1 VSUBS 0.026693f
C30 VDD2.n2 VSUBS 0.014344f
C31 VDD2.n3 VSUBS 0.033903f
C32 VDD2.n4 VSUBS 0.015187f
C33 VDD2.n5 VSUBS 0.026693f
C34 VDD2.n6 VSUBS 0.014344f
C35 VDD2.n7 VSUBS 0.033903f
C36 VDD2.n8 VSUBS 0.015187f
C37 VDD2.n9 VSUBS 0.026693f
C38 VDD2.n10 VSUBS 0.014344f
C39 VDD2.n11 VSUBS 0.033903f
C40 VDD2.n12 VSUBS 0.015187f
C41 VDD2.n13 VSUBS 0.026693f
C42 VDD2.n14 VSUBS 0.014766f
C43 VDD2.n15 VSUBS 0.033903f
C44 VDD2.n16 VSUBS 0.015187f
C45 VDD2.n17 VSUBS 0.026693f
C46 VDD2.n18 VSUBS 0.014344f
C47 VDD2.n19 VSUBS 0.033903f
C48 VDD2.n20 VSUBS 0.015187f
C49 VDD2.n21 VSUBS 0.026693f
C50 VDD2.n22 VSUBS 0.014344f
C51 VDD2.n23 VSUBS 0.025427f
C52 VDD2.n24 VSUBS 0.025504f
C53 VDD2.t5 VSUBS 0.073257f
C54 VDD2.n25 VSUBS 0.237257f
C55 VDD2.n26 VSUBS 1.57351f
C56 VDD2.n27 VSUBS 0.014344f
C57 VDD2.n28 VSUBS 0.015187f
C58 VDD2.n29 VSUBS 0.033903f
C59 VDD2.n30 VSUBS 0.033903f
C60 VDD2.n31 VSUBS 0.015187f
C61 VDD2.n32 VSUBS 0.014344f
C62 VDD2.n33 VSUBS 0.026693f
C63 VDD2.n34 VSUBS 0.026693f
C64 VDD2.n35 VSUBS 0.014344f
C65 VDD2.n36 VSUBS 0.015187f
C66 VDD2.n37 VSUBS 0.033903f
C67 VDD2.n38 VSUBS 0.033903f
C68 VDD2.n39 VSUBS 0.015187f
C69 VDD2.n40 VSUBS 0.014344f
C70 VDD2.n41 VSUBS 0.026693f
C71 VDD2.n42 VSUBS 0.026693f
C72 VDD2.n43 VSUBS 0.014344f
C73 VDD2.n44 VSUBS 0.014344f
C74 VDD2.n45 VSUBS 0.015187f
C75 VDD2.n46 VSUBS 0.033903f
C76 VDD2.n47 VSUBS 0.033903f
C77 VDD2.n48 VSUBS 0.033903f
C78 VDD2.n49 VSUBS 0.014766f
C79 VDD2.n50 VSUBS 0.014344f
C80 VDD2.n51 VSUBS 0.026693f
C81 VDD2.n52 VSUBS 0.026693f
C82 VDD2.n53 VSUBS 0.014344f
C83 VDD2.n54 VSUBS 0.015187f
C84 VDD2.n55 VSUBS 0.033903f
C85 VDD2.n56 VSUBS 0.033903f
C86 VDD2.n57 VSUBS 0.015187f
C87 VDD2.n58 VSUBS 0.014344f
C88 VDD2.n59 VSUBS 0.026693f
C89 VDD2.n60 VSUBS 0.026693f
C90 VDD2.n61 VSUBS 0.014344f
C91 VDD2.n62 VSUBS 0.015187f
C92 VDD2.n63 VSUBS 0.033903f
C93 VDD2.n64 VSUBS 0.033903f
C94 VDD2.n65 VSUBS 0.015187f
C95 VDD2.n66 VSUBS 0.014344f
C96 VDD2.n67 VSUBS 0.026693f
C97 VDD2.n68 VSUBS 0.026693f
C98 VDD2.n69 VSUBS 0.014344f
C99 VDD2.n70 VSUBS 0.015187f
C100 VDD2.n71 VSUBS 0.033903f
C101 VDD2.n72 VSUBS 0.08478f
C102 VDD2.n73 VSUBS 0.015187f
C103 VDD2.n74 VSUBS 0.014344f
C104 VDD2.n75 VSUBS 0.060241f
C105 VDD2.n76 VSUBS 0.061844f
C106 VDD2.t0 VSUBS 0.300374f
C107 VDD2.t2 VSUBS 0.300374f
C108 VDD2.n77 VSUBS 2.40554f
C109 VDD2.n78 VSUBS 2.26524f
C110 VDD2.n79 VSUBS 0.030124f
C111 VDD2.n80 VSUBS 0.026693f
C112 VDD2.n81 VSUBS 0.014344f
C113 VDD2.n82 VSUBS 0.033903f
C114 VDD2.n83 VSUBS 0.015187f
C115 VDD2.n84 VSUBS 0.026693f
C116 VDD2.n85 VSUBS 0.014344f
C117 VDD2.n86 VSUBS 0.033903f
C118 VDD2.n87 VSUBS 0.015187f
C119 VDD2.n88 VSUBS 0.026693f
C120 VDD2.n89 VSUBS 0.014344f
C121 VDD2.n90 VSUBS 0.033903f
C122 VDD2.n91 VSUBS 0.015187f
C123 VDD2.n92 VSUBS 0.026693f
C124 VDD2.n93 VSUBS 0.014766f
C125 VDD2.n94 VSUBS 0.033903f
C126 VDD2.n95 VSUBS 0.014344f
C127 VDD2.n96 VSUBS 0.015187f
C128 VDD2.n97 VSUBS 0.026693f
C129 VDD2.n98 VSUBS 0.014344f
C130 VDD2.n99 VSUBS 0.033903f
C131 VDD2.n100 VSUBS 0.015187f
C132 VDD2.n101 VSUBS 0.026693f
C133 VDD2.n102 VSUBS 0.014344f
C134 VDD2.n103 VSUBS 0.025427f
C135 VDD2.n104 VSUBS 0.025504f
C136 VDD2.t4 VSUBS 0.073257f
C137 VDD2.n105 VSUBS 0.237257f
C138 VDD2.n106 VSUBS 1.57351f
C139 VDD2.n107 VSUBS 0.014344f
C140 VDD2.n108 VSUBS 0.015187f
C141 VDD2.n109 VSUBS 0.033903f
C142 VDD2.n110 VSUBS 0.033903f
C143 VDD2.n111 VSUBS 0.015187f
C144 VDD2.n112 VSUBS 0.014344f
C145 VDD2.n113 VSUBS 0.026693f
C146 VDD2.n114 VSUBS 0.026693f
C147 VDD2.n115 VSUBS 0.014344f
C148 VDD2.n116 VSUBS 0.015187f
C149 VDD2.n117 VSUBS 0.033903f
C150 VDD2.n118 VSUBS 0.033903f
C151 VDD2.n119 VSUBS 0.015187f
C152 VDD2.n120 VSUBS 0.014344f
C153 VDD2.n121 VSUBS 0.026693f
C154 VDD2.n122 VSUBS 0.026693f
C155 VDD2.n123 VSUBS 0.014344f
C156 VDD2.n124 VSUBS 0.015187f
C157 VDD2.n125 VSUBS 0.033903f
C158 VDD2.n126 VSUBS 0.033903f
C159 VDD2.n127 VSUBS 0.033903f
C160 VDD2.n128 VSUBS 0.014766f
C161 VDD2.n129 VSUBS 0.014344f
C162 VDD2.n130 VSUBS 0.026693f
C163 VDD2.n131 VSUBS 0.026693f
C164 VDD2.n132 VSUBS 0.014344f
C165 VDD2.n133 VSUBS 0.015187f
C166 VDD2.n134 VSUBS 0.033903f
C167 VDD2.n135 VSUBS 0.033903f
C168 VDD2.n136 VSUBS 0.015187f
C169 VDD2.n137 VSUBS 0.014344f
C170 VDD2.n138 VSUBS 0.026693f
C171 VDD2.n139 VSUBS 0.026693f
C172 VDD2.n140 VSUBS 0.014344f
C173 VDD2.n141 VSUBS 0.015187f
C174 VDD2.n142 VSUBS 0.033903f
C175 VDD2.n143 VSUBS 0.033903f
C176 VDD2.n144 VSUBS 0.015187f
C177 VDD2.n145 VSUBS 0.014344f
C178 VDD2.n146 VSUBS 0.026693f
C179 VDD2.n147 VSUBS 0.026693f
C180 VDD2.n148 VSUBS 0.014344f
C181 VDD2.n149 VSUBS 0.015187f
C182 VDD2.n150 VSUBS 0.033903f
C183 VDD2.n151 VSUBS 0.08478f
C184 VDD2.n152 VSUBS 0.015187f
C185 VDD2.n153 VSUBS 0.014344f
C186 VDD2.n154 VSUBS 0.060241f
C187 VDD2.n155 VSUBS 0.061152f
C188 VDD2.n156 VSUBS 2.2693f
C189 VDD2.t1 VSUBS 0.300374f
C190 VDD2.t3 VSUBS 0.300374f
C191 VDD2.n157 VSUBS 2.40552f
C192 VN.t0 VSUBS 0.984814f
C193 VN.n0 VSUBS 0.381101f
C194 VN.t5 VSUBS 0.977001f
C195 VN.n1 VSUBS 0.400827f
C196 VN.t3 VSUBS 0.977513f
C197 VN.n2 VSUBS 0.387926f
C198 VN.n3 VSUBS 0.19532f
C199 VN.t2 VSUBS 0.984814f
C200 VN.n4 VSUBS 0.381101f
C201 VN.t1 VSUBS 0.977513f
C202 VN.t4 VSUBS 0.977001f
C203 VN.n5 VSUBS 0.400827f
C204 VN.n6 VSUBS 0.387926f
C205 VN.n7 VSUBS 2.90888f
C206 B.n0 VSUBS 0.004695f
C207 B.n1 VSUBS 0.004695f
C208 B.n2 VSUBS 0.007425f
C209 B.n3 VSUBS 0.007425f
C210 B.n4 VSUBS 0.007425f
C211 B.n5 VSUBS 0.007425f
C212 B.n6 VSUBS 0.007425f
C213 B.n7 VSUBS 0.007425f
C214 B.n8 VSUBS 0.007425f
C215 B.n9 VSUBS 0.007425f
C216 B.n10 VSUBS 0.018677f
C217 B.n11 VSUBS 0.007425f
C218 B.n12 VSUBS 0.007425f
C219 B.n13 VSUBS 0.007425f
C220 B.n14 VSUBS 0.007425f
C221 B.n15 VSUBS 0.007425f
C222 B.n16 VSUBS 0.007425f
C223 B.n17 VSUBS 0.007425f
C224 B.n18 VSUBS 0.007425f
C225 B.n19 VSUBS 0.007425f
C226 B.n20 VSUBS 0.007425f
C227 B.n21 VSUBS 0.007425f
C228 B.n22 VSUBS 0.007425f
C229 B.n23 VSUBS 0.007425f
C230 B.n24 VSUBS 0.007425f
C231 B.n25 VSUBS 0.007425f
C232 B.n26 VSUBS 0.007425f
C233 B.n27 VSUBS 0.007425f
C234 B.n28 VSUBS 0.007425f
C235 B.n29 VSUBS 0.007425f
C236 B.n30 VSUBS 0.007425f
C237 B.n31 VSUBS 0.007425f
C238 B.n32 VSUBS 0.007425f
C239 B.n33 VSUBS 0.007425f
C240 B.t2 VSUBS 0.278037f
C241 B.t1 VSUBS 0.28671f
C242 B.t0 VSUBS 0.213953f
C243 B.n34 VSUBS 0.340662f
C244 B.n35 VSUBS 0.28897f
C245 B.n36 VSUBS 0.017203f
C246 B.n37 VSUBS 0.007425f
C247 B.n38 VSUBS 0.007425f
C248 B.n39 VSUBS 0.007425f
C249 B.n40 VSUBS 0.007425f
C250 B.n41 VSUBS 0.007425f
C251 B.t5 VSUBS 0.278041f
C252 B.t4 VSUBS 0.286713f
C253 B.t3 VSUBS 0.213953f
C254 B.n42 VSUBS 0.340658f
C255 B.n43 VSUBS 0.288966f
C256 B.n44 VSUBS 0.007425f
C257 B.n45 VSUBS 0.007425f
C258 B.n46 VSUBS 0.007425f
C259 B.n47 VSUBS 0.007425f
C260 B.n48 VSUBS 0.007425f
C261 B.n49 VSUBS 0.007425f
C262 B.n50 VSUBS 0.007425f
C263 B.n51 VSUBS 0.007425f
C264 B.n52 VSUBS 0.007425f
C265 B.n53 VSUBS 0.007425f
C266 B.n54 VSUBS 0.007425f
C267 B.n55 VSUBS 0.007425f
C268 B.n56 VSUBS 0.007425f
C269 B.n57 VSUBS 0.007425f
C270 B.n58 VSUBS 0.007425f
C271 B.n59 VSUBS 0.007425f
C272 B.n60 VSUBS 0.007425f
C273 B.n61 VSUBS 0.007425f
C274 B.n62 VSUBS 0.007425f
C275 B.n63 VSUBS 0.007425f
C276 B.n64 VSUBS 0.007425f
C277 B.n65 VSUBS 0.007425f
C278 B.n66 VSUBS 0.007425f
C279 B.n67 VSUBS 0.018677f
C280 B.n68 VSUBS 0.007425f
C281 B.n69 VSUBS 0.007425f
C282 B.n70 VSUBS 0.007425f
C283 B.n71 VSUBS 0.007425f
C284 B.n72 VSUBS 0.007425f
C285 B.n73 VSUBS 0.007425f
C286 B.n74 VSUBS 0.007425f
C287 B.n75 VSUBS 0.007425f
C288 B.n76 VSUBS 0.007425f
C289 B.n77 VSUBS 0.007425f
C290 B.n78 VSUBS 0.007425f
C291 B.n79 VSUBS 0.007425f
C292 B.n80 VSUBS 0.007425f
C293 B.n81 VSUBS 0.007425f
C294 B.n82 VSUBS 0.007425f
C295 B.n83 VSUBS 0.007425f
C296 B.n84 VSUBS 0.018677f
C297 B.n85 VSUBS 0.007425f
C298 B.n86 VSUBS 0.007425f
C299 B.n87 VSUBS 0.007425f
C300 B.n88 VSUBS 0.007425f
C301 B.n89 VSUBS 0.007425f
C302 B.n90 VSUBS 0.007425f
C303 B.n91 VSUBS 0.007425f
C304 B.n92 VSUBS 0.007425f
C305 B.n93 VSUBS 0.007425f
C306 B.n94 VSUBS 0.007425f
C307 B.n95 VSUBS 0.007425f
C308 B.n96 VSUBS 0.007425f
C309 B.n97 VSUBS 0.007425f
C310 B.n98 VSUBS 0.007425f
C311 B.n99 VSUBS 0.007425f
C312 B.n100 VSUBS 0.007425f
C313 B.n101 VSUBS 0.007425f
C314 B.n102 VSUBS 0.007425f
C315 B.n103 VSUBS 0.007425f
C316 B.n104 VSUBS 0.007425f
C317 B.n105 VSUBS 0.007425f
C318 B.n106 VSUBS 0.007425f
C319 B.n107 VSUBS 0.007425f
C320 B.t10 VSUBS 0.278041f
C321 B.t11 VSUBS 0.286713f
C322 B.t9 VSUBS 0.213953f
C323 B.n108 VSUBS 0.340658f
C324 B.n109 VSUBS 0.288966f
C325 B.n110 VSUBS 0.017203f
C326 B.n111 VSUBS 0.007425f
C327 B.n112 VSUBS 0.007425f
C328 B.n113 VSUBS 0.007425f
C329 B.n114 VSUBS 0.007425f
C330 B.n115 VSUBS 0.007425f
C331 B.t7 VSUBS 0.278037f
C332 B.t8 VSUBS 0.28671f
C333 B.t6 VSUBS 0.213953f
C334 B.n116 VSUBS 0.340662f
C335 B.n117 VSUBS 0.28897f
C336 B.n118 VSUBS 0.007425f
C337 B.n119 VSUBS 0.007425f
C338 B.n120 VSUBS 0.007425f
C339 B.n121 VSUBS 0.007425f
C340 B.n122 VSUBS 0.007425f
C341 B.n123 VSUBS 0.007425f
C342 B.n124 VSUBS 0.007425f
C343 B.n125 VSUBS 0.007425f
C344 B.n126 VSUBS 0.007425f
C345 B.n127 VSUBS 0.007425f
C346 B.n128 VSUBS 0.007425f
C347 B.n129 VSUBS 0.007425f
C348 B.n130 VSUBS 0.007425f
C349 B.n131 VSUBS 0.007425f
C350 B.n132 VSUBS 0.007425f
C351 B.n133 VSUBS 0.007425f
C352 B.n134 VSUBS 0.007425f
C353 B.n135 VSUBS 0.007425f
C354 B.n136 VSUBS 0.007425f
C355 B.n137 VSUBS 0.007425f
C356 B.n138 VSUBS 0.007425f
C357 B.n139 VSUBS 0.007425f
C358 B.n140 VSUBS 0.007425f
C359 B.n141 VSUBS 0.018677f
C360 B.n142 VSUBS 0.007425f
C361 B.n143 VSUBS 0.007425f
C362 B.n144 VSUBS 0.007425f
C363 B.n145 VSUBS 0.007425f
C364 B.n146 VSUBS 0.007425f
C365 B.n147 VSUBS 0.007425f
C366 B.n148 VSUBS 0.007425f
C367 B.n149 VSUBS 0.007425f
C368 B.n150 VSUBS 0.007425f
C369 B.n151 VSUBS 0.007425f
C370 B.n152 VSUBS 0.007425f
C371 B.n153 VSUBS 0.007425f
C372 B.n154 VSUBS 0.007425f
C373 B.n155 VSUBS 0.007425f
C374 B.n156 VSUBS 0.007425f
C375 B.n157 VSUBS 0.007425f
C376 B.n158 VSUBS 0.007425f
C377 B.n159 VSUBS 0.007425f
C378 B.n160 VSUBS 0.007425f
C379 B.n161 VSUBS 0.007425f
C380 B.n162 VSUBS 0.007425f
C381 B.n163 VSUBS 0.007425f
C382 B.n164 VSUBS 0.007425f
C383 B.n165 VSUBS 0.007425f
C384 B.n166 VSUBS 0.007425f
C385 B.n167 VSUBS 0.007425f
C386 B.n168 VSUBS 0.007425f
C387 B.n169 VSUBS 0.007425f
C388 B.n170 VSUBS 0.017573f
C389 B.n171 VSUBS 0.017573f
C390 B.n172 VSUBS 0.018677f
C391 B.n173 VSUBS 0.007425f
C392 B.n174 VSUBS 0.007425f
C393 B.n175 VSUBS 0.007425f
C394 B.n176 VSUBS 0.007425f
C395 B.n177 VSUBS 0.007425f
C396 B.n178 VSUBS 0.007425f
C397 B.n179 VSUBS 0.007425f
C398 B.n180 VSUBS 0.007425f
C399 B.n181 VSUBS 0.007425f
C400 B.n182 VSUBS 0.007425f
C401 B.n183 VSUBS 0.007425f
C402 B.n184 VSUBS 0.007425f
C403 B.n185 VSUBS 0.007425f
C404 B.n186 VSUBS 0.007425f
C405 B.n187 VSUBS 0.007425f
C406 B.n188 VSUBS 0.007425f
C407 B.n189 VSUBS 0.007425f
C408 B.n190 VSUBS 0.007425f
C409 B.n191 VSUBS 0.007425f
C410 B.n192 VSUBS 0.007425f
C411 B.n193 VSUBS 0.007425f
C412 B.n194 VSUBS 0.007425f
C413 B.n195 VSUBS 0.007425f
C414 B.n196 VSUBS 0.007425f
C415 B.n197 VSUBS 0.007425f
C416 B.n198 VSUBS 0.007425f
C417 B.n199 VSUBS 0.007425f
C418 B.n200 VSUBS 0.007425f
C419 B.n201 VSUBS 0.007425f
C420 B.n202 VSUBS 0.007425f
C421 B.n203 VSUBS 0.007425f
C422 B.n204 VSUBS 0.007425f
C423 B.n205 VSUBS 0.007425f
C424 B.n206 VSUBS 0.007425f
C425 B.n207 VSUBS 0.007425f
C426 B.n208 VSUBS 0.007425f
C427 B.n209 VSUBS 0.007425f
C428 B.n210 VSUBS 0.007425f
C429 B.n211 VSUBS 0.007425f
C430 B.n212 VSUBS 0.007425f
C431 B.n213 VSUBS 0.007425f
C432 B.n214 VSUBS 0.007425f
C433 B.n215 VSUBS 0.007425f
C434 B.n216 VSUBS 0.007425f
C435 B.n217 VSUBS 0.007425f
C436 B.n218 VSUBS 0.007425f
C437 B.n219 VSUBS 0.007425f
C438 B.n220 VSUBS 0.007425f
C439 B.n221 VSUBS 0.007425f
C440 B.n222 VSUBS 0.007425f
C441 B.n223 VSUBS 0.007425f
C442 B.n224 VSUBS 0.007425f
C443 B.n225 VSUBS 0.007425f
C444 B.n226 VSUBS 0.007425f
C445 B.n227 VSUBS 0.007425f
C446 B.n228 VSUBS 0.007425f
C447 B.n229 VSUBS 0.007425f
C448 B.n230 VSUBS 0.007425f
C449 B.n231 VSUBS 0.007425f
C450 B.n232 VSUBS 0.007425f
C451 B.n233 VSUBS 0.007425f
C452 B.n234 VSUBS 0.007425f
C453 B.n235 VSUBS 0.007425f
C454 B.n236 VSUBS 0.007425f
C455 B.n237 VSUBS 0.007425f
C456 B.n238 VSUBS 0.007425f
C457 B.n239 VSUBS 0.007425f
C458 B.n240 VSUBS 0.007425f
C459 B.n241 VSUBS 0.007425f
C460 B.n242 VSUBS 0.007425f
C461 B.n243 VSUBS 0.006988f
C462 B.n244 VSUBS 0.017203f
C463 B.n245 VSUBS 0.004149f
C464 B.n246 VSUBS 0.007425f
C465 B.n247 VSUBS 0.007425f
C466 B.n248 VSUBS 0.007425f
C467 B.n249 VSUBS 0.007425f
C468 B.n250 VSUBS 0.007425f
C469 B.n251 VSUBS 0.007425f
C470 B.n252 VSUBS 0.007425f
C471 B.n253 VSUBS 0.007425f
C472 B.n254 VSUBS 0.007425f
C473 B.n255 VSUBS 0.007425f
C474 B.n256 VSUBS 0.007425f
C475 B.n257 VSUBS 0.007425f
C476 B.n258 VSUBS 0.004149f
C477 B.n259 VSUBS 0.007425f
C478 B.n260 VSUBS 0.007425f
C479 B.n261 VSUBS 0.006988f
C480 B.n262 VSUBS 0.007425f
C481 B.n263 VSUBS 0.007425f
C482 B.n264 VSUBS 0.007425f
C483 B.n265 VSUBS 0.007425f
C484 B.n266 VSUBS 0.007425f
C485 B.n267 VSUBS 0.007425f
C486 B.n268 VSUBS 0.007425f
C487 B.n269 VSUBS 0.007425f
C488 B.n270 VSUBS 0.007425f
C489 B.n271 VSUBS 0.007425f
C490 B.n272 VSUBS 0.007425f
C491 B.n273 VSUBS 0.007425f
C492 B.n274 VSUBS 0.007425f
C493 B.n275 VSUBS 0.007425f
C494 B.n276 VSUBS 0.007425f
C495 B.n277 VSUBS 0.007425f
C496 B.n278 VSUBS 0.007425f
C497 B.n279 VSUBS 0.007425f
C498 B.n280 VSUBS 0.007425f
C499 B.n281 VSUBS 0.007425f
C500 B.n282 VSUBS 0.007425f
C501 B.n283 VSUBS 0.007425f
C502 B.n284 VSUBS 0.007425f
C503 B.n285 VSUBS 0.007425f
C504 B.n286 VSUBS 0.007425f
C505 B.n287 VSUBS 0.007425f
C506 B.n288 VSUBS 0.007425f
C507 B.n289 VSUBS 0.007425f
C508 B.n290 VSUBS 0.007425f
C509 B.n291 VSUBS 0.007425f
C510 B.n292 VSUBS 0.007425f
C511 B.n293 VSUBS 0.007425f
C512 B.n294 VSUBS 0.007425f
C513 B.n295 VSUBS 0.007425f
C514 B.n296 VSUBS 0.007425f
C515 B.n297 VSUBS 0.007425f
C516 B.n298 VSUBS 0.007425f
C517 B.n299 VSUBS 0.007425f
C518 B.n300 VSUBS 0.007425f
C519 B.n301 VSUBS 0.007425f
C520 B.n302 VSUBS 0.007425f
C521 B.n303 VSUBS 0.007425f
C522 B.n304 VSUBS 0.007425f
C523 B.n305 VSUBS 0.007425f
C524 B.n306 VSUBS 0.007425f
C525 B.n307 VSUBS 0.007425f
C526 B.n308 VSUBS 0.007425f
C527 B.n309 VSUBS 0.007425f
C528 B.n310 VSUBS 0.007425f
C529 B.n311 VSUBS 0.007425f
C530 B.n312 VSUBS 0.007425f
C531 B.n313 VSUBS 0.007425f
C532 B.n314 VSUBS 0.007425f
C533 B.n315 VSUBS 0.007425f
C534 B.n316 VSUBS 0.007425f
C535 B.n317 VSUBS 0.007425f
C536 B.n318 VSUBS 0.007425f
C537 B.n319 VSUBS 0.007425f
C538 B.n320 VSUBS 0.007425f
C539 B.n321 VSUBS 0.007425f
C540 B.n322 VSUBS 0.007425f
C541 B.n323 VSUBS 0.007425f
C542 B.n324 VSUBS 0.007425f
C543 B.n325 VSUBS 0.007425f
C544 B.n326 VSUBS 0.007425f
C545 B.n327 VSUBS 0.007425f
C546 B.n328 VSUBS 0.007425f
C547 B.n329 VSUBS 0.007425f
C548 B.n330 VSUBS 0.007425f
C549 B.n331 VSUBS 0.018677f
C550 B.n332 VSUBS 0.017573f
C551 B.n333 VSUBS 0.017573f
C552 B.n334 VSUBS 0.007425f
C553 B.n335 VSUBS 0.007425f
C554 B.n336 VSUBS 0.007425f
C555 B.n337 VSUBS 0.007425f
C556 B.n338 VSUBS 0.007425f
C557 B.n339 VSUBS 0.007425f
C558 B.n340 VSUBS 0.007425f
C559 B.n341 VSUBS 0.007425f
C560 B.n342 VSUBS 0.007425f
C561 B.n343 VSUBS 0.007425f
C562 B.n344 VSUBS 0.007425f
C563 B.n345 VSUBS 0.007425f
C564 B.n346 VSUBS 0.007425f
C565 B.n347 VSUBS 0.007425f
C566 B.n348 VSUBS 0.007425f
C567 B.n349 VSUBS 0.007425f
C568 B.n350 VSUBS 0.007425f
C569 B.n351 VSUBS 0.007425f
C570 B.n352 VSUBS 0.007425f
C571 B.n353 VSUBS 0.007425f
C572 B.n354 VSUBS 0.007425f
C573 B.n355 VSUBS 0.007425f
C574 B.n356 VSUBS 0.007425f
C575 B.n357 VSUBS 0.007425f
C576 B.n358 VSUBS 0.007425f
C577 B.n359 VSUBS 0.007425f
C578 B.n360 VSUBS 0.007425f
C579 B.n361 VSUBS 0.007425f
C580 B.n362 VSUBS 0.007425f
C581 B.n363 VSUBS 0.007425f
C582 B.n364 VSUBS 0.007425f
C583 B.n365 VSUBS 0.007425f
C584 B.n366 VSUBS 0.007425f
C585 B.n367 VSUBS 0.007425f
C586 B.n368 VSUBS 0.007425f
C587 B.n369 VSUBS 0.007425f
C588 B.n370 VSUBS 0.007425f
C589 B.n371 VSUBS 0.007425f
C590 B.n372 VSUBS 0.007425f
C591 B.n373 VSUBS 0.007425f
C592 B.n374 VSUBS 0.007425f
C593 B.n375 VSUBS 0.007425f
C594 B.n376 VSUBS 0.007425f
C595 B.n377 VSUBS 0.007425f
C596 B.n378 VSUBS 0.007425f
C597 B.n379 VSUBS 0.007425f
C598 B.n380 VSUBS 0.017573f
C599 B.n381 VSUBS 0.018396f
C600 B.n382 VSUBS 0.017854f
C601 B.n383 VSUBS 0.007425f
C602 B.n384 VSUBS 0.007425f
C603 B.n385 VSUBS 0.007425f
C604 B.n386 VSUBS 0.007425f
C605 B.n387 VSUBS 0.007425f
C606 B.n388 VSUBS 0.007425f
C607 B.n389 VSUBS 0.007425f
C608 B.n390 VSUBS 0.007425f
C609 B.n391 VSUBS 0.007425f
C610 B.n392 VSUBS 0.007425f
C611 B.n393 VSUBS 0.007425f
C612 B.n394 VSUBS 0.007425f
C613 B.n395 VSUBS 0.007425f
C614 B.n396 VSUBS 0.007425f
C615 B.n397 VSUBS 0.007425f
C616 B.n398 VSUBS 0.007425f
C617 B.n399 VSUBS 0.007425f
C618 B.n400 VSUBS 0.007425f
C619 B.n401 VSUBS 0.007425f
C620 B.n402 VSUBS 0.007425f
C621 B.n403 VSUBS 0.007425f
C622 B.n404 VSUBS 0.007425f
C623 B.n405 VSUBS 0.007425f
C624 B.n406 VSUBS 0.007425f
C625 B.n407 VSUBS 0.007425f
C626 B.n408 VSUBS 0.007425f
C627 B.n409 VSUBS 0.007425f
C628 B.n410 VSUBS 0.007425f
C629 B.n411 VSUBS 0.007425f
C630 B.n412 VSUBS 0.007425f
C631 B.n413 VSUBS 0.007425f
C632 B.n414 VSUBS 0.007425f
C633 B.n415 VSUBS 0.007425f
C634 B.n416 VSUBS 0.007425f
C635 B.n417 VSUBS 0.007425f
C636 B.n418 VSUBS 0.007425f
C637 B.n419 VSUBS 0.007425f
C638 B.n420 VSUBS 0.007425f
C639 B.n421 VSUBS 0.007425f
C640 B.n422 VSUBS 0.007425f
C641 B.n423 VSUBS 0.007425f
C642 B.n424 VSUBS 0.007425f
C643 B.n425 VSUBS 0.007425f
C644 B.n426 VSUBS 0.007425f
C645 B.n427 VSUBS 0.007425f
C646 B.n428 VSUBS 0.007425f
C647 B.n429 VSUBS 0.007425f
C648 B.n430 VSUBS 0.007425f
C649 B.n431 VSUBS 0.007425f
C650 B.n432 VSUBS 0.007425f
C651 B.n433 VSUBS 0.007425f
C652 B.n434 VSUBS 0.007425f
C653 B.n435 VSUBS 0.007425f
C654 B.n436 VSUBS 0.007425f
C655 B.n437 VSUBS 0.007425f
C656 B.n438 VSUBS 0.007425f
C657 B.n439 VSUBS 0.007425f
C658 B.n440 VSUBS 0.007425f
C659 B.n441 VSUBS 0.007425f
C660 B.n442 VSUBS 0.007425f
C661 B.n443 VSUBS 0.007425f
C662 B.n444 VSUBS 0.007425f
C663 B.n445 VSUBS 0.007425f
C664 B.n446 VSUBS 0.007425f
C665 B.n447 VSUBS 0.007425f
C666 B.n448 VSUBS 0.007425f
C667 B.n449 VSUBS 0.007425f
C668 B.n450 VSUBS 0.007425f
C669 B.n451 VSUBS 0.007425f
C670 B.n452 VSUBS 0.007425f
C671 B.n453 VSUBS 0.006988f
C672 B.n454 VSUBS 0.017203f
C673 B.n455 VSUBS 0.004149f
C674 B.n456 VSUBS 0.007425f
C675 B.n457 VSUBS 0.007425f
C676 B.n458 VSUBS 0.007425f
C677 B.n459 VSUBS 0.007425f
C678 B.n460 VSUBS 0.007425f
C679 B.n461 VSUBS 0.007425f
C680 B.n462 VSUBS 0.007425f
C681 B.n463 VSUBS 0.007425f
C682 B.n464 VSUBS 0.007425f
C683 B.n465 VSUBS 0.007425f
C684 B.n466 VSUBS 0.007425f
C685 B.n467 VSUBS 0.007425f
C686 B.n468 VSUBS 0.004149f
C687 B.n469 VSUBS 0.007425f
C688 B.n470 VSUBS 0.007425f
C689 B.n471 VSUBS 0.006988f
C690 B.n472 VSUBS 0.007425f
C691 B.n473 VSUBS 0.007425f
C692 B.n474 VSUBS 0.007425f
C693 B.n475 VSUBS 0.007425f
C694 B.n476 VSUBS 0.007425f
C695 B.n477 VSUBS 0.007425f
C696 B.n478 VSUBS 0.007425f
C697 B.n479 VSUBS 0.007425f
C698 B.n480 VSUBS 0.007425f
C699 B.n481 VSUBS 0.007425f
C700 B.n482 VSUBS 0.007425f
C701 B.n483 VSUBS 0.007425f
C702 B.n484 VSUBS 0.007425f
C703 B.n485 VSUBS 0.007425f
C704 B.n486 VSUBS 0.007425f
C705 B.n487 VSUBS 0.007425f
C706 B.n488 VSUBS 0.007425f
C707 B.n489 VSUBS 0.007425f
C708 B.n490 VSUBS 0.007425f
C709 B.n491 VSUBS 0.007425f
C710 B.n492 VSUBS 0.007425f
C711 B.n493 VSUBS 0.007425f
C712 B.n494 VSUBS 0.007425f
C713 B.n495 VSUBS 0.007425f
C714 B.n496 VSUBS 0.007425f
C715 B.n497 VSUBS 0.007425f
C716 B.n498 VSUBS 0.007425f
C717 B.n499 VSUBS 0.007425f
C718 B.n500 VSUBS 0.007425f
C719 B.n501 VSUBS 0.007425f
C720 B.n502 VSUBS 0.007425f
C721 B.n503 VSUBS 0.007425f
C722 B.n504 VSUBS 0.007425f
C723 B.n505 VSUBS 0.007425f
C724 B.n506 VSUBS 0.007425f
C725 B.n507 VSUBS 0.007425f
C726 B.n508 VSUBS 0.007425f
C727 B.n509 VSUBS 0.007425f
C728 B.n510 VSUBS 0.007425f
C729 B.n511 VSUBS 0.007425f
C730 B.n512 VSUBS 0.007425f
C731 B.n513 VSUBS 0.007425f
C732 B.n514 VSUBS 0.007425f
C733 B.n515 VSUBS 0.007425f
C734 B.n516 VSUBS 0.007425f
C735 B.n517 VSUBS 0.007425f
C736 B.n518 VSUBS 0.007425f
C737 B.n519 VSUBS 0.007425f
C738 B.n520 VSUBS 0.007425f
C739 B.n521 VSUBS 0.007425f
C740 B.n522 VSUBS 0.007425f
C741 B.n523 VSUBS 0.007425f
C742 B.n524 VSUBS 0.007425f
C743 B.n525 VSUBS 0.007425f
C744 B.n526 VSUBS 0.007425f
C745 B.n527 VSUBS 0.007425f
C746 B.n528 VSUBS 0.007425f
C747 B.n529 VSUBS 0.007425f
C748 B.n530 VSUBS 0.007425f
C749 B.n531 VSUBS 0.007425f
C750 B.n532 VSUBS 0.007425f
C751 B.n533 VSUBS 0.007425f
C752 B.n534 VSUBS 0.007425f
C753 B.n535 VSUBS 0.007425f
C754 B.n536 VSUBS 0.007425f
C755 B.n537 VSUBS 0.007425f
C756 B.n538 VSUBS 0.007425f
C757 B.n539 VSUBS 0.007425f
C758 B.n540 VSUBS 0.007425f
C759 B.n541 VSUBS 0.018677f
C760 B.n542 VSUBS 0.017573f
C761 B.n543 VSUBS 0.017573f
C762 B.n544 VSUBS 0.007425f
C763 B.n545 VSUBS 0.007425f
C764 B.n546 VSUBS 0.007425f
C765 B.n547 VSUBS 0.007425f
C766 B.n548 VSUBS 0.007425f
C767 B.n549 VSUBS 0.007425f
C768 B.n550 VSUBS 0.007425f
C769 B.n551 VSUBS 0.007425f
C770 B.n552 VSUBS 0.007425f
C771 B.n553 VSUBS 0.007425f
C772 B.n554 VSUBS 0.007425f
C773 B.n555 VSUBS 0.007425f
C774 B.n556 VSUBS 0.007425f
C775 B.n557 VSUBS 0.007425f
C776 B.n558 VSUBS 0.007425f
C777 B.n559 VSUBS 0.007425f
C778 B.n560 VSUBS 0.007425f
C779 B.n561 VSUBS 0.007425f
C780 B.n562 VSUBS 0.007425f
C781 B.n563 VSUBS 0.007425f
C782 B.n564 VSUBS 0.007425f
C783 B.n565 VSUBS 0.007425f
C784 B.n566 VSUBS 0.007425f
C785 B.n567 VSUBS 0.016812f
C786 VDD1.n0 VSUBS 0.030126f
C787 VDD1.n1 VSUBS 0.026695f
C788 VDD1.n2 VSUBS 0.014345f
C789 VDD1.n3 VSUBS 0.033906f
C790 VDD1.n4 VSUBS 0.015189f
C791 VDD1.n5 VSUBS 0.026695f
C792 VDD1.n6 VSUBS 0.014345f
C793 VDD1.n7 VSUBS 0.033906f
C794 VDD1.n8 VSUBS 0.015189f
C795 VDD1.n9 VSUBS 0.026695f
C796 VDD1.n10 VSUBS 0.014345f
C797 VDD1.n11 VSUBS 0.033906f
C798 VDD1.n12 VSUBS 0.015189f
C799 VDD1.n13 VSUBS 0.026695f
C800 VDD1.n14 VSUBS 0.014767f
C801 VDD1.n15 VSUBS 0.033906f
C802 VDD1.n16 VSUBS 0.014345f
C803 VDD1.n17 VSUBS 0.015189f
C804 VDD1.n18 VSUBS 0.026695f
C805 VDD1.n19 VSUBS 0.014345f
C806 VDD1.n20 VSUBS 0.033906f
C807 VDD1.n21 VSUBS 0.015189f
C808 VDD1.n22 VSUBS 0.026695f
C809 VDD1.n23 VSUBS 0.014345f
C810 VDD1.n24 VSUBS 0.025429f
C811 VDD1.n25 VSUBS 0.025506f
C812 VDD1.t4 VSUBS 0.073262f
C813 VDD1.n26 VSUBS 0.237275f
C814 VDD1.n27 VSUBS 1.57363f
C815 VDD1.n28 VSUBS 0.014345f
C816 VDD1.n29 VSUBS 0.015189f
C817 VDD1.n30 VSUBS 0.033906f
C818 VDD1.n31 VSUBS 0.033906f
C819 VDD1.n32 VSUBS 0.015189f
C820 VDD1.n33 VSUBS 0.014345f
C821 VDD1.n34 VSUBS 0.026695f
C822 VDD1.n35 VSUBS 0.026695f
C823 VDD1.n36 VSUBS 0.014345f
C824 VDD1.n37 VSUBS 0.015189f
C825 VDD1.n38 VSUBS 0.033906f
C826 VDD1.n39 VSUBS 0.033906f
C827 VDD1.n40 VSUBS 0.015189f
C828 VDD1.n41 VSUBS 0.014345f
C829 VDD1.n42 VSUBS 0.026695f
C830 VDD1.n43 VSUBS 0.026695f
C831 VDD1.n44 VSUBS 0.014345f
C832 VDD1.n45 VSUBS 0.015189f
C833 VDD1.n46 VSUBS 0.033906f
C834 VDD1.n47 VSUBS 0.033906f
C835 VDD1.n48 VSUBS 0.033906f
C836 VDD1.n49 VSUBS 0.014767f
C837 VDD1.n50 VSUBS 0.014345f
C838 VDD1.n51 VSUBS 0.026695f
C839 VDD1.n52 VSUBS 0.026695f
C840 VDD1.n53 VSUBS 0.014345f
C841 VDD1.n54 VSUBS 0.015189f
C842 VDD1.n55 VSUBS 0.033906f
C843 VDD1.n56 VSUBS 0.033906f
C844 VDD1.n57 VSUBS 0.015189f
C845 VDD1.n58 VSUBS 0.014345f
C846 VDD1.n59 VSUBS 0.026695f
C847 VDD1.n60 VSUBS 0.026695f
C848 VDD1.n61 VSUBS 0.014345f
C849 VDD1.n62 VSUBS 0.015189f
C850 VDD1.n63 VSUBS 0.033906f
C851 VDD1.n64 VSUBS 0.033906f
C852 VDD1.n65 VSUBS 0.015189f
C853 VDD1.n66 VSUBS 0.014345f
C854 VDD1.n67 VSUBS 0.026695f
C855 VDD1.n68 VSUBS 0.026695f
C856 VDD1.n69 VSUBS 0.014345f
C857 VDD1.n70 VSUBS 0.015189f
C858 VDD1.n71 VSUBS 0.033906f
C859 VDD1.n72 VSUBS 0.084786f
C860 VDD1.n73 VSUBS 0.015189f
C861 VDD1.n74 VSUBS 0.014345f
C862 VDD1.n75 VSUBS 0.060246f
C863 VDD1.n76 VSUBS 0.062132f
C864 VDD1.n77 VSUBS 0.030126f
C865 VDD1.n78 VSUBS 0.026695f
C866 VDD1.n79 VSUBS 0.014345f
C867 VDD1.n80 VSUBS 0.033906f
C868 VDD1.n81 VSUBS 0.015189f
C869 VDD1.n82 VSUBS 0.026695f
C870 VDD1.n83 VSUBS 0.014345f
C871 VDD1.n84 VSUBS 0.033906f
C872 VDD1.n85 VSUBS 0.015189f
C873 VDD1.n86 VSUBS 0.026695f
C874 VDD1.n87 VSUBS 0.014345f
C875 VDD1.n88 VSUBS 0.033906f
C876 VDD1.n89 VSUBS 0.015189f
C877 VDD1.n90 VSUBS 0.026695f
C878 VDD1.n91 VSUBS 0.014767f
C879 VDD1.n92 VSUBS 0.033906f
C880 VDD1.n93 VSUBS 0.015189f
C881 VDD1.n94 VSUBS 0.026695f
C882 VDD1.n95 VSUBS 0.014345f
C883 VDD1.n96 VSUBS 0.033906f
C884 VDD1.n97 VSUBS 0.015189f
C885 VDD1.n98 VSUBS 0.026695f
C886 VDD1.n99 VSUBS 0.014345f
C887 VDD1.n100 VSUBS 0.025429f
C888 VDD1.n101 VSUBS 0.025506f
C889 VDD1.t1 VSUBS 0.073262f
C890 VDD1.n102 VSUBS 0.237275f
C891 VDD1.n103 VSUBS 1.57363f
C892 VDD1.n104 VSUBS 0.014345f
C893 VDD1.n105 VSUBS 0.015189f
C894 VDD1.n106 VSUBS 0.033906f
C895 VDD1.n107 VSUBS 0.033906f
C896 VDD1.n108 VSUBS 0.015189f
C897 VDD1.n109 VSUBS 0.014345f
C898 VDD1.n110 VSUBS 0.026695f
C899 VDD1.n111 VSUBS 0.026695f
C900 VDD1.n112 VSUBS 0.014345f
C901 VDD1.n113 VSUBS 0.015189f
C902 VDD1.n114 VSUBS 0.033906f
C903 VDD1.n115 VSUBS 0.033906f
C904 VDD1.n116 VSUBS 0.015189f
C905 VDD1.n117 VSUBS 0.014345f
C906 VDD1.n118 VSUBS 0.026695f
C907 VDD1.n119 VSUBS 0.026695f
C908 VDD1.n120 VSUBS 0.014345f
C909 VDD1.n121 VSUBS 0.014345f
C910 VDD1.n122 VSUBS 0.015189f
C911 VDD1.n123 VSUBS 0.033906f
C912 VDD1.n124 VSUBS 0.033906f
C913 VDD1.n125 VSUBS 0.033906f
C914 VDD1.n126 VSUBS 0.014767f
C915 VDD1.n127 VSUBS 0.014345f
C916 VDD1.n128 VSUBS 0.026695f
C917 VDD1.n129 VSUBS 0.026695f
C918 VDD1.n130 VSUBS 0.014345f
C919 VDD1.n131 VSUBS 0.015189f
C920 VDD1.n132 VSUBS 0.033906f
C921 VDD1.n133 VSUBS 0.033906f
C922 VDD1.n134 VSUBS 0.015189f
C923 VDD1.n135 VSUBS 0.014345f
C924 VDD1.n136 VSUBS 0.026695f
C925 VDD1.n137 VSUBS 0.026695f
C926 VDD1.n138 VSUBS 0.014345f
C927 VDD1.n139 VSUBS 0.015189f
C928 VDD1.n140 VSUBS 0.033906f
C929 VDD1.n141 VSUBS 0.033906f
C930 VDD1.n142 VSUBS 0.015189f
C931 VDD1.n143 VSUBS 0.014345f
C932 VDD1.n144 VSUBS 0.026695f
C933 VDD1.n145 VSUBS 0.026695f
C934 VDD1.n146 VSUBS 0.014345f
C935 VDD1.n147 VSUBS 0.015189f
C936 VDD1.n148 VSUBS 0.033906f
C937 VDD1.n149 VSUBS 0.084786f
C938 VDD1.n150 VSUBS 0.015189f
C939 VDD1.n151 VSUBS 0.014345f
C940 VDD1.n152 VSUBS 0.060246f
C941 VDD1.n153 VSUBS 0.061848f
C942 VDD1.t2 VSUBS 0.300397f
C943 VDD1.t5 VSUBS 0.300397f
C944 VDD1.n154 VSUBS 2.40573f
C945 VDD1.n155 VSUBS 2.3399f
C946 VDD1.t3 VSUBS 0.300397f
C947 VDD1.t0 VSUBS 0.300397f
C948 VDD1.n156 VSUBS 2.40495f
C949 VDD1.n157 VSUBS 2.79064f
C950 VTAIL.t0 VSUBS 0.358397f
C951 VTAIL.t2 VSUBS 0.358397f
C952 VTAIL.n0 VSUBS 2.67968f
C953 VTAIL.n1 VSUBS 0.86825f
C954 VTAIL.n2 VSUBS 0.035943f
C955 VTAIL.n3 VSUBS 0.031849f
C956 VTAIL.n4 VSUBS 0.017114f
C957 VTAIL.n5 VSUBS 0.040452f
C958 VTAIL.n6 VSUBS 0.018121f
C959 VTAIL.n7 VSUBS 0.031849f
C960 VTAIL.n8 VSUBS 0.017114f
C961 VTAIL.n9 VSUBS 0.040452f
C962 VTAIL.n10 VSUBS 0.018121f
C963 VTAIL.n11 VSUBS 0.031849f
C964 VTAIL.n12 VSUBS 0.017114f
C965 VTAIL.n13 VSUBS 0.040452f
C966 VTAIL.n14 VSUBS 0.018121f
C967 VTAIL.n15 VSUBS 0.031849f
C968 VTAIL.n16 VSUBS 0.017618f
C969 VTAIL.n17 VSUBS 0.040452f
C970 VTAIL.n18 VSUBS 0.018121f
C971 VTAIL.n19 VSUBS 0.031849f
C972 VTAIL.n20 VSUBS 0.017114f
C973 VTAIL.n21 VSUBS 0.040452f
C974 VTAIL.n22 VSUBS 0.018121f
C975 VTAIL.n23 VSUBS 0.031849f
C976 VTAIL.n24 VSUBS 0.017114f
C977 VTAIL.n25 VSUBS 0.030339f
C978 VTAIL.n26 VSUBS 0.03043f
C979 VTAIL.t3 VSUBS 0.087408f
C980 VTAIL.n27 VSUBS 0.283087f
C981 VTAIL.n28 VSUBS 1.87746f
C982 VTAIL.n29 VSUBS 0.017114f
C983 VTAIL.n30 VSUBS 0.018121f
C984 VTAIL.n31 VSUBS 0.040452f
C985 VTAIL.n32 VSUBS 0.040452f
C986 VTAIL.n33 VSUBS 0.018121f
C987 VTAIL.n34 VSUBS 0.017114f
C988 VTAIL.n35 VSUBS 0.031849f
C989 VTAIL.n36 VSUBS 0.031849f
C990 VTAIL.n37 VSUBS 0.017114f
C991 VTAIL.n38 VSUBS 0.018121f
C992 VTAIL.n39 VSUBS 0.040452f
C993 VTAIL.n40 VSUBS 0.040452f
C994 VTAIL.n41 VSUBS 0.018121f
C995 VTAIL.n42 VSUBS 0.017114f
C996 VTAIL.n43 VSUBS 0.031849f
C997 VTAIL.n44 VSUBS 0.031849f
C998 VTAIL.n45 VSUBS 0.017114f
C999 VTAIL.n46 VSUBS 0.017114f
C1000 VTAIL.n47 VSUBS 0.018121f
C1001 VTAIL.n48 VSUBS 0.040452f
C1002 VTAIL.n49 VSUBS 0.040452f
C1003 VTAIL.n50 VSUBS 0.040452f
C1004 VTAIL.n51 VSUBS 0.017618f
C1005 VTAIL.n52 VSUBS 0.017114f
C1006 VTAIL.n53 VSUBS 0.031849f
C1007 VTAIL.n54 VSUBS 0.031849f
C1008 VTAIL.n55 VSUBS 0.017114f
C1009 VTAIL.n56 VSUBS 0.018121f
C1010 VTAIL.n57 VSUBS 0.040452f
C1011 VTAIL.n58 VSUBS 0.040452f
C1012 VTAIL.n59 VSUBS 0.018121f
C1013 VTAIL.n60 VSUBS 0.017114f
C1014 VTAIL.n61 VSUBS 0.031849f
C1015 VTAIL.n62 VSUBS 0.031849f
C1016 VTAIL.n63 VSUBS 0.017114f
C1017 VTAIL.n64 VSUBS 0.018121f
C1018 VTAIL.n65 VSUBS 0.040452f
C1019 VTAIL.n66 VSUBS 0.040452f
C1020 VTAIL.n67 VSUBS 0.018121f
C1021 VTAIL.n68 VSUBS 0.017114f
C1022 VTAIL.n69 VSUBS 0.031849f
C1023 VTAIL.n70 VSUBS 0.031849f
C1024 VTAIL.n71 VSUBS 0.017114f
C1025 VTAIL.n72 VSUBS 0.018121f
C1026 VTAIL.n73 VSUBS 0.040452f
C1027 VTAIL.n74 VSUBS 0.101156f
C1028 VTAIL.n75 VSUBS 0.018121f
C1029 VTAIL.n76 VSUBS 0.017114f
C1030 VTAIL.n77 VSUBS 0.071878f
C1031 VTAIL.n78 VSUBS 0.05096f
C1032 VTAIL.n79 VSUBS 0.166003f
C1033 VTAIL.t5 VSUBS 0.358397f
C1034 VTAIL.t6 VSUBS 0.358397f
C1035 VTAIL.n80 VSUBS 2.67968f
C1036 VTAIL.n81 VSUBS 2.64387f
C1037 VTAIL.t11 VSUBS 0.358397f
C1038 VTAIL.t9 VSUBS 0.358397f
C1039 VTAIL.n82 VSUBS 2.67969f
C1040 VTAIL.n83 VSUBS 2.64386f
C1041 VTAIL.n84 VSUBS 0.035943f
C1042 VTAIL.n85 VSUBS 0.031849f
C1043 VTAIL.n86 VSUBS 0.017114f
C1044 VTAIL.n87 VSUBS 0.040452f
C1045 VTAIL.n88 VSUBS 0.018121f
C1046 VTAIL.n89 VSUBS 0.031849f
C1047 VTAIL.n90 VSUBS 0.017114f
C1048 VTAIL.n91 VSUBS 0.040452f
C1049 VTAIL.n92 VSUBS 0.018121f
C1050 VTAIL.n93 VSUBS 0.031849f
C1051 VTAIL.n94 VSUBS 0.017114f
C1052 VTAIL.n95 VSUBS 0.040452f
C1053 VTAIL.n96 VSUBS 0.018121f
C1054 VTAIL.n97 VSUBS 0.031849f
C1055 VTAIL.n98 VSUBS 0.017618f
C1056 VTAIL.n99 VSUBS 0.040452f
C1057 VTAIL.n100 VSUBS 0.017114f
C1058 VTAIL.n101 VSUBS 0.018121f
C1059 VTAIL.n102 VSUBS 0.031849f
C1060 VTAIL.n103 VSUBS 0.017114f
C1061 VTAIL.n104 VSUBS 0.040452f
C1062 VTAIL.n105 VSUBS 0.018121f
C1063 VTAIL.n106 VSUBS 0.031849f
C1064 VTAIL.n107 VSUBS 0.017114f
C1065 VTAIL.n108 VSUBS 0.030339f
C1066 VTAIL.n109 VSUBS 0.03043f
C1067 VTAIL.t10 VSUBS 0.087408f
C1068 VTAIL.n110 VSUBS 0.283087f
C1069 VTAIL.n111 VSUBS 1.87746f
C1070 VTAIL.n112 VSUBS 0.017114f
C1071 VTAIL.n113 VSUBS 0.018121f
C1072 VTAIL.n114 VSUBS 0.040452f
C1073 VTAIL.n115 VSUBS 0.040452f
C1074 VTAIL.n116 VSUBS 0.018121f
C1075 VTAIL.n117 VSUBS 0.017114f
C1076 VTAIL.n118 VSUBS 0.031849f
C1077 VTAIL.n119 VSUBS 0.031849f
C1078 VTAIL.n120 VSUBS 0.017114f
C1079 VTAIL.n121 VSUBS 0.018121f
C1080 VTAIL.n122 VSUBS 0.040452f
C1081 VTAIL.n123 VSUBS 0.040452f
C1082 VTAIL.n124 VSUBS 0.018121f
C1083 VTAIL.n125 VSUBS 0.017114f
C1084 VTAIL.n126 VSUBS 0.031849f
C1085 VTAIL.n127 VSUBS 0.031849f
C1086 VTAIL.n128 VSUBS 0.017114f
C1087 VTAIL.n129 VSUBS 0.018121f
C1088 VTAIL.n130 VSUBS 0.040452f
C1089 VTAIL.n131 VSUBS 0.040452f
C1090 VTAIL.n132 VSUBS 0.040452f
C1091 VTAIL.n133 VSUBS 0.017618f
C1092 VTAIL.n134 VSUBS 0.017114f
C1093 VTAIL.n135 VSUBS 0.031849f
C1094 VTAIL.n136 VSUBS 0.031849f
C1095 VTAIL.n137 VSUBS 0.017114f
C1096 VTAIL.n138 VSUBS 0.018121f
C1097 VTAIL.n139 VSUBS 0.040452f
C1098 VTAIL.n140 VSUBS 0.040452f
C1099 VTAIL.n141 VSUBS 0.018121f
C1100 VTAIL.n142 VSUBS 0.017114f
C1101 VTAIL.n143 VSUBS 0.031849f
C1102 VTAIL.n144 VSUBS 0.031849f
C1103 VTAIL.n145 VSUBS 0.017114f
C1104 VTAIL.n146 VSUBS 0.018121f
C1105 VTAIL.n147 VSUBS 0.040452f
C1106 VTAIL.n148 VSUBS 0.040452f
C1107 VTAIL.n149 VSUBS 0.018121f
C1108 VTAIL.n150 VSUBS 0.017114f
C1109 VTAIL.n151 VSUBS 0.031849f
C1110 VTAIL.n152 VSUBS 0.031849f
C1111 VTAIL.n153 VSUBS 0.017114f
C1112 VTAIL.n154 VSUBS 0.018121f
C1113 VTAIL.n155 VSUBS 0.040452f
C1114 VTAIL.n156 VSUBS 0.101156f
C1115 VTAIL.n157 VSUBS 0.018121f
C1116 VTAIL.n158 VSUBS 0.017114f
C1117 VTAIL.n159 VSUBS 0.071878f
C1118 VTAIL.n160 VSUBS 0.05096f
C1119 VTAIL.n161 VSUBS 0.166003f
C1120 VTAIL.t8 VSUBS 0.358397f
C1121 VTAIL.t7 VSUBS 0.358397f
C1122 VTAIL.n162 VSUBS 2.67969f
C1123 VTAIL.n163 VSUBS 0.908049f
C1124 VTAIL.n164 VSUBS 0.035943f
C1125 VTAIL.n165 VSUBS 0.031849f
C1126 VTAIL.n166 VSUBS 0.017114f
C1127 VTAIL.n167 VSUBS 0.040452f
C1128 VTAIL.n168 VSUBS 0.018121f
C1129 VTAIL.n169 VSUBS 0.031849f
C1130 VTAIL.n170 VSUBS 0.017114f
C1131 VTAIL.n171 VSUBS 0.040452f
C1132 VTAIL.n172 VSUBS 0.018121f
C1133 VTAIL.n173 VSUBS 0.031849f
C1134 VTAIL.n174 VSUBS 0.017114f
C1135 VTAIL.n175 VSUBS 0.040452f
C1136 VTAIL.n176 VSUBS 0.018121f
C1137 VTAIL.n177 VSUBS 0.031849f
C1138 VTAIL.n178 VSUBS 0.017618f
C1139 VTAIL.n179 VSUBS 0.040452f
C1140 VTAIL.n180 VSUBS 0.017114f
C1141 VTAIL.n181 VSUBS 0.018121f
C1142 VTAIL.n182 VSUBS 0.031849f
C1143 VTAIL.n183 VSUBS 0.017114f
C1144 VTAIL.n184 VSUBS 0.040452f
C1145 VTAIL.n185 VSUBS 0.018121f
C1146 VTAIL.n186 VSUBS 0.031849f
C1147 VTAIL.n187 VSUBS 0.017114f
C1148 VTAIL.n188 VSUBS 0.030339f
C1149 VTAIL.n189 VSUBS 0.03043f
C1150 VTAIL.t4 VSUBS 0.087408f
C1151 VTAIL.n190 VSUBS 0.283087f
C1152 VTAIL.n191 VSUBS 1.87746f
C1153 VTAIL.n192 VSUBS 0.017114f
C1154 VTAIL.n193 VSUBS 0.018121f
C1155 VTAIL.n194 VSUBS 0.040452f
C1156 VTAIL.n195 VSUBS 0.040452f
C1157 VTAIL.n196 VSUBS 0.018121f
C1158 VTAIL.n197 VSUBS 0.017114f
C1159 VTAIL.n198 VSUBS 0.031849f
C1160 VTAIL.n199 VSUBS 0.031849f
C1161 VTAIL.n200 VSUBS 0.017114f
C1162 VTAIL.n201 VSUBS 0.018121f
C1163 VTAIL.n202 VSUBS 0.040452f
C1164 VTAIL.n203 VSUBS 0.040452f
C1165 VTAIL.n204 VSUBS 0.018121f
C1166 VTAIL.n205 VSUBS 0.017114f
C1167 VTAIL.n206 VSUBS 0.031849f
C1168 VTAIL.n207 VSUBS 0.031849f
C1169 VTAIL.n208 VSUBS 0.017114f
C1170 VTAIL.n209 VSUBS 0.018121f
C1171 VTAIL.n210 VSUBS 0.040452f
C1172 VTAIL.n211 VSUBS 0.040452f
C1173 VTAIL.n212 VSUBS 0.040452f
C1174 VTAIL.n213 VSUBS 0.017618f
C1175 VTAIL.n214 VSUBS 0.017114f
C1176 VTAIL.n215 VSUBS 0.031849f
C1177 VTAIL.n216 VSUBS 0.031849f
C1178 VTAIL.n217 VSUBS 0.017114f
C1179 VTAIL.n218 VSUBS 0.018121f
C1180 VTAIL.n219 VSUBS 0.040452f
C1181 VTAIL.n220 VSUBS 0.040452f
C1182 VTAIL.n221 VSUBS 0.018121f
C1183 VTAIL.n222 VSUBS 0.017114f
C1184 VTAIL.n223 VSUBS 0.031849f
C1185 VTAIL.n224 VSUBS 0.031849f
C1186 VTAIL.n225 VSUBS 0.017114f
C1187 VTAIL.n226 VSUBS 0.018121f
C1188 VTAIL.n227 VSUBS 0.040452f
C1189 VTAIL.n228 VSUBS 0.040452f
C1190 VTAIL.n229 VSUBS 0.018121f
C1191 VTAIL.n230 VSUBS 0.017114f
C1192 VTAIL.n231 VSUBS 0.031849f
C1193 VTAIL.n232 VSUBS 0.031849f
C1194 VTAIL.n233 VSUBS 0.017114f
C1195 VTAIL.n234 VSUBS 0.018121f
C1196 VTAIL.n235 VSUBS 0.040452f
C1197 VTAIL.n236 VSUBS 0.101156f
C1198 VTAIL.n237 VSUBS 0.018121f
C1199 VTAIL.n238 VSUBS 0.017114f
C1200 VTAIL.n239 VSUBS 0.071878f
C1201 VTAIL.n240 VSUBS 0.05096f
C1202 VTAIL.n241 VSUBS 1.84077f
C1203 VTAIL.n242 VSUBS 0.035943f
C1204 VTAIL.n243 VSUBS 0.031849f
C1205 VTAIL.n244 VSUBS 0.017114f
C1206 VTAIL.n245 VSUBS 0.040452f
C1207 VTAIL.n246 VSUBS 0.018121f
C1208 VTAIL.n247 VSUBS 0.031849f
C1209 VTAIL.n248 VSUBS 0.017114f
C1210 VTAIL.n249 VSUBS 0.040452f
C1211 VTAIL.n250 VSUBS 0.018121f
C1212 VTAIL.n251 VSUBS 0.031849f
C1213 VTAIL.n252 VSUBS 0.017114f
C1214 VTAIL.n253 VSUBS 0.040452f
C1215 VTAIL.n254 VSUBS 0.018121f
C1216 VTAIL.n255 VSUBS 0.031849f
C1217 VTAIL.n256 VSUBS 0.017618f
C1218 VTAIL.n257 VSUBS 0.040452f
C1219 VTAIL.n258 VSUBS 0.018121f
C1220 VTAIL.n259 VSUBS 0.031849f
C1221 VTAIL.n260 VSUBS 0.017114f
C1222 VTAIL.n261 VSUBS 0.040452f
C1223 VTAIL.n262 VSUBS 0.018121f
C1224 VTAIL.n263 VSUBS 0.031849f
C1225 VTAIL.n264 VSUBS 0.017114f
C1226 VTAIL.n265 VSUBS 0.030339f
C1227 VTAIL.n266 VSUBS 0.03043f
C1228 VTAIL.t1 VSUBS 0.087408f
C1229 VTAIL.n267 VSUBS 0.283087f
C1230 VTAIL.n268 VSUBS 1.87746f
C1231 VTAIL.n269 VSUBS 0.017114f
C1232 VTAIL.n270 VSUBS 0.018121f
C1233 VTAIL.n271 VSUBS 0.040452f
C1234 VTAIL.n272 VSUBS 0.040452f
C1235 VTAIL.n273 VSUBS 0.018121f
C1236 VTAIL.n274 VSUBS 0.017114f
C1237 VTAIL.n275 VSUBS 0.031849f
C1238 VTAIL.n276 VSUBS 0.031849f
C1239 VTAIL.n277 VSUBS 0.017114f
C1240 VTAIL.n278 VSUBS 0.018121f
C1241 VTAIL.n279 VSUBS 0.040452f
C1242 VTAIL.n280 VSUBS 0.040452f
C1243 VTAIL.n281 VSUBS 0.018121f
C1244 VTAIL.n282 VSUBS 0.017114f
C1245 VTAIL.n283 VSUBS 0.031849f
C1246 VTAIL.n284 VSUBS 0.031849f
C1247 VTAIL.n285 VSUBS 0.017114f
C1248 VTAIL.n286 VSUBS 0.017114f
C1249 VTAIL.n287 VSUBS 0.018121f
C1250 VTAIL.n288 VSUBS 0.040452f
C1251 VTAIL.n289 VSUBS 0.040452f
C1252 VTAIL.n290 VSUBS 0.040452f
C1253 VTAIL.n291 VSUBS 0.017618f
C1254 VTAIL.n292 VSUBS 0.017114f
C1255 VTAIL.n293 VSUBS 0.031849f
C1256 VTAIL.n294 VSUBS 0.031849f
C1257 VTAIL.n295 VSUBS 0.017114f
C1258 VTAIL.n296 VSUBS 0.018121f
C1259 VTAIL.n297 VSUBS 0.040452f
C1260 VTAIL.n298 VSUBS 0.040452f
C1261 VTAIL.n299 VSUBS 0.018121f
C1262 VTAIL.n300 VSUBS 0.017114f
C1263 VTAIL.n301 VSUBS 0.031849f
C1264 VTAIL.n302 VSUBS 0.031849f
C1265 VTAIL.n303 VSUBS 0.017114f
C1266 VTAIL.n304 VSUBS 0.018121f
C1267 VTAIL.n305 VSUBS 0.040452f
C1268 VTAIL.n306 VSUBS 0.040452f
C1269 VTAIL.n307 VSUBS 0.018121f
C1270 VTAIL.n308 VSUBS 0.017114f
C1271 VTAIL.n309 VSUBS 0.031849f
C1272 VTAIL.n310 VSUBS 0.031849f
C1273 VTAIL.n311 VSUBS 0.017114f
C1274 VTAIL.n312 VSUBS 0.018121f
C1275 VTAIL.n313 VSUBS 0.040452f
C1276 VTAIL.n314 VSUBS 0.101156f
C1277 VTAIL.n315 VSUBS 0.018121f
C1278 VTAIL.n316 VSUBS 0.017114f
C1279 VTAIL.n317 VSUBS 0.071878f
C1280 VTAIL.n318 VSUBS 0.05096f
C1281 VTAIL.n319 VSUBS 1.81953f
C1282 VP.n0 VSUBS 0.068871f
C1283 VP.t4 VSUBS 1.00502f
C1284 VP.t1 VSUBS 1.01253f
C1285 VP.n1 VSUBS 0.391826f
C1286 VP.t2 VSUBS 1.0045f
C1287 VP.n2 VSUBS 0.412108f
C1288 VP.t5 VSUBS 1.00502f
C1289 VP.n3 VSUBS 0.398843f
C1290 VP.n4 VSUBS 2.94551f
C1291 VP.n5 VSUBS 2.8574f
C1292 VP.n6 VSUBS 0.398843f
C1293 VP.t3 VSUBS 1.0045f
C1294 VP.n7 VSUBS 0.412108f
C1295 VP.t0 VSUBS 1.00502f
C1296 VP.n8 VSUBS 0.398843f
C1297 VP.n9 VSUBS 0.053373f
.ends

