* NGSPICE file created from diff_pair_sample_0033.ext - technology: sky130A

.subckt diff_pair_sample_0033 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t9 VN.t0 VTAIL.t11 B.t1 sky130_fd_pr__nfet_01v8 ad=0.3993 pd=2.75 as=0.3993 ps=2.75 w=2.42 l=1.33
X1 VTAIL.t18 VN.t1 VDD2.t8 B.t0 sky130_fd_pr__nfet_01v8 ad=0.3993 pd=2.75 as=0.3993 ps=2.75 w=2.42 l=1.33
X2 B.t23 B.t21 B.t22 B.t18 sky130_fd_pr__nfet_01v8 ad=0.9438 pd=5.62 as=0 ps=0 w=2.42 l=1.33
X3 VTAIL.t0 VP.t0 VDD1.t9 B.t0 sky130_fd_pr__nfet_01v8 ad=0.3993 pd=2.75 as=0.3993 ps=2.75 w=2.42 l=1.33
X4 VDD2.t7 VN.t2 VTAIL.t10 B.t4 sky130_fd_pr__nfet_01v8 ad=0.3993 pd=2.75 as=0.3993 ps=2.75 w=2.42 l=1.33
X5 VDD1.t8 VP.t1 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=0.9438 pd=5.62 as=0.3993 ps=2.75 w=2.42 l=1.33
X6 VTAIL.t19 VN.t3 VDD2.t6 B.t8 sky130_fd_pr__nfet_01v8 ad=0.3993 pd=2.75 as=0.3993 ps=2.75 w=2.42 l=1.33
X7 VDD1.t7 VP.t2 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.3993 pd=2.75 as=0.3993 ps=2.75 w=2.42 l=1.33
X8 VTAIL.t9 VP.t3 VDD1.t6 B.t9 sky130_fd_pr__nfet_01v8 ad=0.3993 pd=2.75 as=0.3993 ps=2.75 w=2.42 l=1.33
X9 VDD2.t5 VN.t4 VTAIL.t16 B.t7 sky130_fd_pr__nfet_01v8 ad=0.3993 pd=2.75 as=0.9438 ps=5.62 w=2.42 l=1.33
X10 B.t20 B.t17 B.t19 B.t18 sky130_fd_pr__nfet_01v8 ad=0.9438 pd=5.62 as=0 ps=0 w=2.42 l=1.33
X11 VDD1.t5 VP.t4 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=0.3993 pd=2.75 as=0.9438 ps=5.62 w=2.42 l=1.33
X12 VDD2.t4 VN.t5 VTAIL.t12 B.t3 sky130_fd_pr__nfet_01v8 ad=0.3993 pd=2.75 as=0.9438 ps=5.62 w=2.42 l=1.33
X13 VTAIL.t15 VN.t6 VDD2.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=0.3993 pd=2.75 as=0.3993 ps=2.75 w=2.42 l=1.33
X14 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=0.9438 pd=5.62 as=0 ps=0 w=2.42 l=1.33
X15 VDD1.t4 VP.t5 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=0.9438 pd=5.62 as=0.3993 ps=2.75 w=2.42 l=1.33
X16 VDD2.t2 VN.t7 VTAIL.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=0.9438 pd=5.62 as=0.3993 ps=2.75 w=2.42 l=1.33
X17 VTAIL.t8 VP.t6 VDD1.t3 B.t8 sky130_fd_pr__nfet_01v8 ad=0.3993 pd=2.75 as=0.3993 ps=2.75 w=2.42 l=1.33
X18 VTAIL.t14 VN.t8 VDD2.t1 B.t9 sky130_fd_pr__nfet_01v8 ad=0.3993 pd=2.75 as=0.3993 ps=2.75 w=2.42 l=1.33
X19 VDD1.t2 VP.t7 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.3993 pd=2.75 as=0.9438 ps=5.62 w=2.42 l=1.33
X20 VTAIL.t2 VP.t8 VDD1.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=0.3993 pd=2.75 as=0.3993 ps=2.75 w=2.42 l=1.33
X21 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=0.9438 pd=5.62 as=0 ps=0 w=2.42 l=1.33
X22 VDD1.t0 VP.t9 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.3993 pd=2.75 as=0.3993 ps=2.75 w=2.42 l=1.33
X23 VDD2.t0 VN.t9 VTAIL.t17 B.t6 sky130_fd_pr__nfet_01v8 ad=0.9438 pd=5.62 as=0.3993 ps=2.75 w=2.42 l=1.33
R0 VN.n24 VN.n23 170.154
R1 VN.n49 VN.n48 170.154
R2 VN.n47 VN.n25 161.3
R3 VN.n46 VN.n45 161.3
R4 VN.n44 VN.n26 161.3
R5 VN.n43 VN.n42 161.3
R6 VN.n41 VN.n27 161.3
R7 VN.n40 VN.n39 161.3
R8 VN.n38 VN.n29 161.3
R9 VN.n37 VN.n36 161.3
R10 VN.n35 VN.n30 161.3
R11 VN.n34 VN.n33 161.3
R12 VN.n22 VN.n0 161.3
R13 VN.n21 VN.n20 161.3
R14 VN.n19 VN.n1 161.3
R15 VN.n18 VN.n17 161.3
R16 VN.n15 VN.n2 161.3
R17 VN.n14 VN.n13 161.3
R18 VN.n12 VN.n3 161.3
R19 VN.n11 VN.n10 161.3
R20 VN.n9 VN.n4 161.3
R21 VN.n8 VN.n7 161.3
R22 VN.n6 VN.t9 75.5805
R23 VN.n32 VN.t5 75.5805
R24 VN.n6 VN.n5 56.6996
R25 VN.n32 VN.n31 56.6996
R26 VN.n10 VN.n9 56.5617
R27 VN.n15 VN.n14 56.5617
R28 VN.n36 VN.n35 56.5617
R29 VN.n41 VN.n40 56.5617
R30 VN.n3 VN.t0 43.8516
R31 VN.n5 VN.t8 43.8516
R32 VN.n16 VN.t6 43.8516
R33 VN.n23 VN.t4 43.8516
R34 VN.n29 VN.t2 43.8516
R35 VN.n31 VN.t3 43.8516
R36 VN.n28 VN.t1 43.8516
R37 VN.n48 VN.t7 43.8516
R38 VN.n21 VN.n1 41.5458
R39 VN.n46 VN.n26 41.5458
R40 VN.n22 VN.n21 39.6083
R41 VN.n47 VN.n46 39.6083
R42 VN VN.n49 39.3054
R43 VN.n33 VN.n32 26.5036
R44 VN.n7 VN.n6 26.5036
R45 VN.n9 VN.n8 24.5923
R46 VN.n10 VN.n3 24.5923
R47 VN.n14 VN.n3 24.5923
R48 VN.n17 VN.n15 24.5923
R49 VN.n35 VN.n34 24.5923
R50 VN.n40 VN.n29 24.5923
R51 VN.n36 VN.n29 24.5923
R52 VN.n42 VN.n41 24.5923
R53 VN.n16 VN.n1 16.7229
R54 VN.n28 VN.n26 16.7229
R55 VN.n23 VN.n22 15.7393
R56 VN.n48 VN.n47 15.7393
R57 VN.n8 VN.n5 7.86989
R58 VN.n17 VN.n16 7.86989
R59 VN.n34 VN.n31 7.86989
R60 VN.n42 VN.n28 7.86989
R61 VN.n49 VN.n25 0.189894
R62 VN.n45 VN.n25 0.189894
R63 VN.n45 VN.n44 0.189894
R64 VN.n44 VN.n43 0.189894
R65 VN.n43 VN.n27 0.189894
R66 VN.n39 VN.n27 0.189894
R67 VN.n39 VN.n38 0.189894
R68 VN.n38 VN.n37 0.189894
R69 VN.n37 VN.n30 0.189894
R70 VN.n33 VN.n30 0.189894
R71 VN.n7 VN.n4 0.189894
R72 VN.n11 VN.n4 0.189894
R73 VN.n12 VN.n11 0.189894
R74 VN.n13 VN.n12 0.189894
R75 VN.n13 VN.n2 0.189894
R76 VN.n18 VN.n2 0.189894
R77 VN.n19 VN.n18 0.189894
R78 VN.n20 VN.n19 0.189894
R79 VN.n20 VN.n0 0.189894
R80 VN.n24 VN.n0 0.189894
R81 VN VN.n24 0.0516364
R82 VTAIL.n56 VTAIL.n50 289.615
R83 VTAIL.n8 VTAIL.n2 289.615
R84 VTAIL.n44 VTAIL.n38 289.615
R85 VTAIL.n28 VTAIL.n22 289.615
R86 VTAIL.n55 VTAIL.n54 185
R87 VTAIL.n57 VTAIL.n56 185
R88 VTAIL.n7 VTAIL.n6 185
R89 VTAIL.n9 VTAIL.n8 185
R90 VTAIL.n45 VTAIL.n44 185
R91 VTAIL.n43 VTAIL.n42 185
R92 VTAIL.n29 VTAIL.n28 185
R93 VTAIL.n27 VTAIL.n26 185
R94 VTAIL.n53 VTAIL.t16 151.613
R95 VTAIL.n5 VTAIL.t3 151.613
R96 VTAIL.n41 VTAIL.t7 151.613
R97 VTAIL.n25 VTAIL.t12 151.613
R98 VTAIL.n56 VTAIL.n55 104.615
R99 VTAIL.n8 VTAIL.n7 104.615
R100 VTAIL.n44 VTAIL.n43 104.615
R101 VTAIL.n28 VTAIL.n27 104.615
R102 VTAIL.n37 VTAIL.n36 68.6684
R103 VTAIL.n35 VTAIL.n34 68.6684
R104 VTAIL.n21 VTAIL.n20 68.6684
R105 VTAIL.n19 VTAIL.n18 68.6684
R106 VTAIL.n63 VTAIL.n62 68.6683
R107 VTAIL.n1 VTAIL.n0 68.6683
R108 VTAIL.n15 VTAIL.n14 68.6683
R109 VTAIL.n17 VTAIL.n16 68.6683
R110 VTAIL.n55 VTAIL.t16 52.3082
R111 VTAIL.n7 VTAIL.t3 52.3082
R112 VTAIL.n43 VTAIL.t7 52.3082
R113 VTAIL.n27 VTAIL.t12 52.3082
R114 VTAIL.n61 VTAIL.n60 32.5732
R115 VTAIL.n13 VTAIL.n12 32.5732
R116 VTAIL.n49 VTAIL.n48 32.5732
R117 VTAIL.n33 VTAIL.n32 32.5732
R118 VTAIL.n19 VTAIL.n17 17.3152
R119 VTAIL.n61 VTAIL.n49 15.8841
R120 VTAIL.n54 VTAIL.n53 15.3979
R121 VTAIL.n6 VTAIL.n5 15.3979
R122 VTAIL.n42 VTAIL.n41 15.3979
R123 VTAIL.n26 VTAIL.n25 15.3979
R124 VTAIL.n57 VTAIL.n52 12.8005
R125 VTAIL.n9 VTAIL.n4 12.8005
R126 VTAIL.n45 VTAIL.n40 12.8005
R127 VTAIL.n29 VTAIL.n24 12.8005
R128 VTAIL.n58 VTAIL.n50 12.0247
R129 VTAIL.n10 VTAIL.n2 12.0247
R130 VTAIL.n46 VTAIL.n38 12.0247
R131 VTAIL.n30 VTAIL.n22 12.0247
R132 VTAIL.n60 VTAIL.n59 9.45567
R133 VTAIL.n12 VTAIL.n11 9.45567
R134 VTAIL.n48 VTAIL.n47 9.45567
R135 VTAIL.n32 VTAIL.n31 9.45567
R136 VTAIL.n59 VTAIL.n58 9.3005
R137 VTAIL.n52 VTAIL.n51 9.3005
R138 VTAIL.n11 VTAIL.n10 9.3005
R139 VTAIL.n4 VTAIL.n3 9.3005
R140 VTAIL.n47 VTAIL.n46 9.3005
R141 VTAIL.n40 VTAIL.n39 9.3005
R142 VTAIL.n31 VTAIL.n30 9.3005
R143 VTAIL.n24 VTAIL.n23 9.3005
R144 VTAIL.n62 VTAIL.t11 8.18232
R145 VTAIL.n62 VTAIL.t15 8.18232
R146 VTAIL.n0 VTAIL.t17 8.18232
R147 VTAIL.n0 VTAIL.t14 8.18232
R148 VTAIL.n14 VTAIL.t4 8.18232
R149 VTAIL.n14 VTAIL.t8 8.18232
R150 VTAIL.n16 VTAIL.t5 8.18232
R151 VTAIL.n16 VTAIL.t0 8.18232
R152 VTAIL.n36 VTAIL.t1 8.18232
R153 VTAIL.n36 VTAIL.t2 8.18232
R154 VTAIL.n34 VTAIL.t6 8.18232
R155 VTAIL.n34 VTAIL.t9 8.18232
R156 VTAIL.n20 VTAIL.t10 8.18232
R157 VTAIL.n20 VTAIL.t19 8.18232
R158 VTAIL.n18 VTAIL.t13 8.18232
R159 VTAIL.n18 VTAIL.t18 8.18232
R160 VTAIL.n53 VTAIL.n51 4.69785
R161 VTAIL.n5 VTAIL.n3 4.69785
R162 VTAIL.n41 VTAIL.n39 4.69785
R163 VTAIL.n25 VTAIL.n23 4.69785
R164 VTAIL.n60 VTAIL.n50 1.93989
R165 VTAIL.n12 VTAIL.n2 1.93989
R166 VTAIL.n48 VTAIL.n38 1.93989
R167 VTAIL.n32 VTAIL.n22 1.93989
R168 VTAIL.n21 VTAIL.n19 1.43153
R169 VTAIL.n33 VTAIL.n21 1.43153
R170 VTAIL.n37 VTAIL.n35 1.43153
R171 VTAIL.n49 VTAIL.n37 1.43153
R172 VTAIL.n17 VTAIL.n15 1.43153
R173 VTAIL.n15 VTAIL.n13 1.43153
R174 VTAIL.n63 VTAIL.n61 1.43153
R175 VTAIL.n35 VTAIL.n33 1.18584
R176 VTAIL.n13 VTAIL.n1 1.18584
R177 VTAIL.n58 VTAIL.n57 1.16414
R178 VTAIL.n10 VTAIL.n9 1.16414
R179 VTAIL.n46 VTAIL.n45 1.16414
R180 VTAIL.n30 VTAIL.n29 1.16414
R181 VTAIL VTAIL.n1 1.13197
R182 VTAIL.n54 VTAIL.n52 0.388379
R183 VTAIL.n6 VTAIL.n4 0.388379
R184 VTAIL.n42 VTAIL.n40 0.388379
R185 VTAIL.n26 VTAIL.n24 0.388379
R186 VTAIL VTAIL.n63 0.300069
R187 VTAIL.n59 VTAIL.n51 0.155672
R188 VTAIL.n11 VTAIL.n3 0.155672
R189 VTAIL.n47 VTAIL.n39 0.155672
R190 VTAIL.n31 VTAIL.n23 0.155672
R191 VDD2.n21 VDD2.n15 289.615
R192 VDD2.n6 VDD2.n0 289.615
R193 VDD2.n22 VDD2.n21 185
R194 VDD2.n20 VDD2.n19 185
R195 VDD2.n5 VDD2.n4 185
R196 VDD2.n7 VDD2.n6 185
R197 VDD2.n18 VDD2.t2 151.613
R198 VDD2.n3 VDD2.t0 151.613
R199 VDD2.n21 VDD2.n20 104.615
R200 VDD2.n6 VDD2.n5 104.615
R201 VDD2.n14 VDD2.n13 86.365
R202 VDD2 VDD2.n29 86.3621
R203 VDD2.n28 VDD2.n27 85.3472
R204 VDD2.n12 VDD2.n11 85.3471
R205 VDD2.n20 VDD2.t2 52.3082
R206 VDD2.n5 VDD2.t0 52.3082
R207 VDD2.n12 VDD2.n10 50.6831
R208 VDD2.n26 VDD2.n25 49.252
R209 VDD2.n26 VDD2.n14 32.5989
R210 VDD2.n19 VDD2.n18 15.3979
R211 VDD2.n4 VDD2.n3 15.3979
R212 VDD2.n22 VDD2.n17 12.8005
R213 VDD2.n7 VDD2.n2 12.8005
R214 VDD2.n23 VDD2.n15 12.0247
R215 VDD2.n8 VDD2.n0 12.0247
R216 VDD2.n25 VDD2.n24 9.45567
R217 VDD2.n10 VDD2.n9 9.45567
R218 VDD2.n24 VDD2.n23 9.3005
R219 VDD2.n17 VDD2.n16 9.3005
R220 VDD2.n9 VDD2.n8 9.3005
R221 VDD2.n2 VDD2.n1 9.3005
R222 VDD2.n29 VDD2.t6 8.18232
R223 VDD2.n29 VDD2.t4 8.18232
R224 VDD2.n27 VDD2.t8 8.18232
R225 VDD2.n27 VDD2.t7 8.18232
R226 VDD2.n13 VDD2.t3 8.18232
R227 VDD2.n13 VDD2.t5 8.18232
R228 VDD2.n11 VDD2.t1 8.18232
R229 VDD2.n11 VDD2.t9 8.18232
R230 VDD2.n18 VDD2.n16 4.69785
R231 VDD2.n3 VDD2.n1 4.69785
R232 VDD2.n25 VDD2.n15 1.93989
R233 VDD2.n10 VDD2.n0 1.93989
R234 VDD2.n28 VDD2.n26 1.43153
R235 VDD2.n23 VDD2.n22 1.16414
R236 VDD2.n8 VDD2.n7 1.16414
R237 VDD2 VDD2.n28 0.416448
R238 VDD2.n19 VDD2.n17 0.388379
R239 VDD2.n4 VDD2.n2 0.388379
R240 VDD2.n14 VDD2.n12 0.302913
R241 VDD2.n24 VDD2.n16 0.155672
R242 VDD2.n9 VDD2.n1 0.155672
R243 B.n492 B.n491 585
R244 B.n162 B.n87 585
R245 B.n161 B.n160 585
R246 B.n159 B.n158 585
R247 B.n157 B.n156 585
R248 B.n155 B.n154 585
R249 B.n153 B.n152 585
R250 B.n151 B.n150 585
R251 B.n149 B.n148 585
R252 B.n147 B.n146 585
R253 B.n145 B.n144 585
R254 B.n143 B.n142 585
R255 B.n141 B.n140 585
R256 B.n138 B.n137 585
R257 B.n136 B.n135 585
R258 B.n134 B.n133 585
R259 B.n132 B.n131 585
R260 B.n130 B.n129 585
R261 B.n128 B.n127 585
R262 B.n126 B.n125 585
R263 B.n124 B.n123 585
R264 B.n122 B.n121 585
R265 B.n120 B.n119 585
R266 B.n117 B.n116 585
R267 B.n115 B.n114 585
R268 B.n113 B.n112 585
R269 B.n111 B.n110 585
R270 B.n109 B.n108 585
R271 B.n107 B.n106 585
R272 B.n105 B.n104 585
R273 B.n103 B.n102 585
R274 B.n101 B.n100 585
R275 B.n99 B.n98 585
R276 B.n97 B.n96 585
R277 B.n95 B.n94 585
R278 B.n93 B.n92 585
R279 B.n490 B.n69 585
R280 B.n495 B.n69 585
R281 B.n489 B.n68 585
R282 B.n496 B.n68 585
R283 B.n488 B.n487 585
R284 B.n487 B.n64 585
R285 B.n486 B.n63 585
R286 B.n502 B.n63 585
R287 B.n485 B.n62 585
R288 B.n503 B.n62 585
R289 B.n484 B.n61 585
R290 B.n504 B.n61 585
R291 B.n483 B.n482 585
R292 B.n482 B.n57 585
R293 B.n481 B.n56 585
R294 B.n510 B.n56 585
R295 B.n480 B.n55 585
R296 B.n511 B.n55 585
R297 B.n479 B.n54 585
R298 B.n512 B.n54 585
R299 B.n478 B.n477 585
R300 B.n477 B.n50 585
R301 B.n476 B.n49 585
R302 B.n518 B.n49 585
R303 B.n475 B.n48 585
R304 B.n519 B.n48 585
R305 B.n474 B.n47 585
R306 B.n520 B.n47 585
R307 B.n473 B.n472 585
R308 B.n472 B.n43 585
R309 B.n471 B.n42 585
R310 B.n526 B.n42 585
R311 B.n470 B.n41 585
R312 B.n527 B.n41 585
R313 B.n469 B.n40 585
R314 B.n528 B.n40 585
R315 B.n468 B.n467 585
R316 B.n467 B.n39 585
R317 B.n466 B.n35 585
R318 B.n534 B.n35 585
R319 B.n465 B.n34 585
R320 B.n535 B.n34 585
R321 B.n464 B.n33 585
R322 B.n536 B.n33 585
R323 B.n463 B.n462 585
R324 B.n462 B.n29 585
R325 B.n461 B.n28 585
R326 B.n542 B.n28 585
R327 B.n460 B.n27 585
R328 B.n543 B.n27 585
R329 B.n459 B.n26 585
R330 B.n544 B.n26 585
R331 B.n458 B.n457 585
R332 B.n457 B.n22 585
R333 B.n456 B.n21 585
R334 B.n550 B.n21 585
R335 B.n455 B.n20 585
R336 B.n551 B.n20 585
R337 B.n454 B.n19 585
R338 B.n552 B.n19 585
R339 B.n453 B.n452 585
R340 B.n452 B.n15 585
R341 B.n451 B.n14 585
R342 B.n558 B.n14 585
R343 B.n450 B.n13 585
R344 B.n559 B.n13 585
R345 B.n449 B.n12 585
R346 B.n560 B.n12 585
R347 B.n448 B.n447 585
R348 B.n447 B.n446 585
R349 B.n445 B.n444 585
R350 B.n445 B.n8 585
R351 B.n443 B.n7 585
R352 B.n567 B.n7 585
R353 B.n442 B.n6 585
R354 B.n568 B.n6 585
R355 B.n441 B.n5 585
R356 B.n569 B.n5 585
R357 B.n440 B.n439 585
R358 B.n439 B.n4 585
R359 B.n438 B.n163 585
R360 B.n438 B.n437 585
R361 B.n428 B.n164 585
R362 B.n165 B.n164 585
R363 B.n430 B.n429 585
R364 B.n431 B.n430 585
R365 B.n427 B.n170 585
R366 B.n170 B.n169 585
R367 B.n426 B.n425 585
R368 B.n425 B.n424 585
R369 B.n172 B.n171 585
R370 B.n173 B.n172 585
R371 B.n417 B.n416 585
R372 B.n418 B.n417 585
R373 B.n415 B.n177 585
R374 B.n181 B.n177 585
R375 B.n414 B.n413 585
R376 B.n413 B.n412 585
R377 B.n179 B.n178 585
R378 B.n180 B.n179 585
R379 B.n405 B.n404 585
R380 B.n406 B.n405 585
R381 B.n403 B.n186 585
R382 B.n186 B.n185 585
R383 B.n402 B.n401 585
R384 B.n401 B.n400 585
R385 B.n188 B.n187 585
R386 B.n189 B.n188 585
R387 B.n393 B.n392 585
R388 B.n394 B.n393 585
R389 B.n391 B.n194 585
R390 B.n194 B.n193 585
R391 B.n390 B.n389 585
R392 B.n389 B.n388 585
R393 B.n196 B.n195 585
R394 B.n381 B.n196 585
R395 B.n380 B.n379 585
R396 B.n382 B.n380 585
R397 B.n378 B.n201 585
R398 B.n201 B.n200 585
R399 B.n377 B.n376 585
R400 B.n376 B.n375 585
R401 B.n203 B.n202 585
R402 B.n204 B.n203 585
R403 B.n368 B.n367 585
R404 B.n369 B.n368 585
R405 B.n366 B.n209 585
R406 B.n209 B.n208 585
R407 B.n365 B.n364 585
R408 B.n364 B.n363 585
R409 B.n211 B.n210 585
R410 B.n212 B.n211 585
R411 B.n356 B.n355 585
R412 B.n357 B.n356 585
R413 B.n354 B.n217 585
R414 B.n217 B.n216 585
R415 B.n353 B.n352 585
R416 B.n352 B.n351 585
R417 B.n219 B.n218 585
R418 B.n220 B.n219 585
R419 B.n344 B.n343 585
R420 B.n345 B.n344 585
R421 B.n342 B.n225 585
R422 B.n225 B.n224 585
R423 B.n341 B.n340 585
R424 B.n340 B.n339 585
R425 B.n227 B.n226 585
R426 B.n228 B.n227 585
R427 B.n332 B.n331 585
R428 B.n333 B.n332 585
R429 B.n330 B.n233 585
R430 B.n233 B.n232 585
R431 B.n325 B.n324 585
R432 B.n323 B.n253 585
R433 B.n322 B.n252 585
R434 B.n327 B.n252 585
R435 B.n321 B.n320 585
R436 B.n319 B.n318 585
R437 B.n317 B.n316 585
R438 B.n315 B.n314 585
R439 B.n313 B.n312 585
R440 B.n311 B.n310 585
R441 B.n309 B.n308 585
R442 B.n307 B.n306 585
R443 B.n305 B.n304 585
R444 B.n303 B.n302 585
R445 B.n301 B.n300 585
R446 B.n299 B.n298 585
R447 B.n297 B.n296 585
R448 B.n295 B.n294 585
R449 B.n293 B.n292 585
R450 B.n291 B.n290 585
R451 B.n289 B.n288 585
R452 B.n287 B.n286 585
R453 B.n285 B.n284 585
R454 B.n283 B.n282 585
R455 B.n281 B.n280 585
R456 B.n279 B.n278 585
R457 B.n277 B.n276 585
R458 B.n275 B.n274 585
R459 B.n273 B.n272 585
R460 B.n271 B.n270 585
R461 B.n269 B.n268 585
R462 B.n267 B.n266 585
R463 B.n265 B.n264 585
R464 B.n263 B.n262 585
R465 B.n261 B.n260 585
R466 B.n235 B.n234 585
R467 B.n329 B.n328 585
R468 B.n328 B.n327 585
R469 B.n231 B.n230 585
R470 B.n232 B.n231 585
R471 B.n335 B.n334 585
R472 B.n334 B.n333 585
R473 B.n336 B.n229 585
R474 B.n229 B.n228 585
R475 B.n338 B.n337 585
R476 B.n339 B.n338 585
R477 B.n223 B.n222 585
R478 B.n224 B.n223 585
R479 B.n347 B.n346 585
R480 B.n346 B.n345 585
R481 B.n348 B.n221 585
R482 B.n221 B.n220 585
R483 B.n350 B.n349 585
R484 B.n351 B.n350 585
R485 B.n215 B.n214 585
R486 B.n216 B.n215 585
R487 B.n359 B.n358 585
R488 B.n358 B.n357 585
R489 B.n360 B.n213 585
R490 B.n213 B.n212 585
R491 B.n362 B.n361 585
R492 B.n363 B.n362 585
R493 B.n207 B.n206 585
R494 B.n208 B.n207 585
R495 B.n371 B.n370 585
R496 B.n370 B.n369 585
R497 B.n372 B.n205 585
R498 B.n205 B.n204 585
R499 B.n374 B.n373 585
R500 B.n375 B.n374 585
R501 B.n199 B.n198 585
R502 B.n200 B.n199 585
R503 B.n384 B.n383 585
R504 B.n383 B.n382 585
R505 B.n385 B.n197 585
R506 B.n381 B.n197 585
R507 B.n387 B.n386 585
R508 B.n388 B.n387 585
R509 B.n192 B.n191 585
R510 B.n193 B.n192 585
R511 B.n396 B.n395 585
R512 B.n395 B.n394 585
R513 B.n397 B.n190 585
R514 B.n190 B.n189 585
R515 B.n399 B.n398 585
R516 B.n400 B.n399 585
R517 B.n184 B.n183 585
R518 B.n185 B.n184 585
R519 B.n408 B.n407 585
R520 B.n407 B.n406 585
R521 B.n409 B.n182 585
R522 B.n182 B.n180 585
R523 B.n411 B.n410 585
R524 B.n412 B.n411 585
R525 B.n176 B.n175 585
R526 B.n181 B.n176 585
R527 B.n420 B.n419 585
R528 B.n419 B.n418 585
R529 B.n421 B.n174 585
R530 B.n174 B.n173 585
R531 B.n423 B.n422 585
R532 B.n424 B.n423 585
R533 B.n168 B.n167 585
R534 B.n169 B.n168 585
R535 B.n433 B.n432 585
R536 B.n432 B.n431 585
R537 B.n434 B.n166 585
R538 B.n166 B.n165 585
R539 B.n436 B.n435 585
R540 B.n437 B.n436 585
R541 B.n3 B.n0 585
R542 B.n4 B.n3 585
R543 B.n566 B.n1 585
R544 B.n567 B.n566 585
R545 B.n565 B.n564 585
R546 B.n565 B.n8 585
R547 B.n563 B.n9 585
R548 B.n446 B.n9 585
R549 B.n562 B.n561 585
R550 B.n561 B.n560 585
R551 B.n11 B.n10 585
R552 B.n559 B.n11 585
R553 B.n557 B.n556 585
R554 B.n558 B.n557 585
R555 B.n555 B.n16 585
R556 B.n16 B.n15 585
R557 B.n554 B.n553 585
R558 B.n553 B.n552 585
R559 B.n18 B.n17 585
R560 B.n551 B.n18 585
R561 B.n549 B.n548 585
R562 B.n550 B.n549 585
R563 B.n547 B.n23 585
R564 B.n23 B.n22 585
R565 B.n546 B.n545 585
R566 B.n545 B.n544 585
R567 B.n25 B.n24 585
R568 B.n543 B.n25 585
R569 B.n541 B.n540 585
R570 B.n542 B.n541 585
R571 B.n539 B.n30 585
R572 B.n30 B.n29 585
R573 B.n538 B.n537 585
R574 B.n537 B.n536 585
R575 B.n32 B.n31 585
R576 B.n535 B.n32 585
R577 B.n533 B.n532 585
R578 B.n534 B.n533 585
R579 B.n531 B.n36 585
R580 B.n39 B.n36 585
R581 B.n530 B.n529 585
R582 B.n529 B.n528 585
R583 B.n38 B.n37 585
R584 B.n527 B.n38 585
R585 B.n525 B.n524 585
R586 B.n526 B.n525 585
R587 B.n523 B.n44 585
R588 B.n44 B.n43 585
R589 B.n522 B.n521 585
R590 B.n521 B.n520 585
R591 B.n46 B.n45 585
R592 B.n519 B.n46 585
R593 B.n517 B.n516 585
R594 B.n518 B.n517 585
R595 B.n515 B.n51 585
R596 B.n51 B.n50 585
R597 B.n514 B.n513 585
R598 B.n513 B.n512 585
R599 B.n53 B.n52 585
R600 B.n511 B.n53 585
R601 B.n509 B.n508 585
R602 B.n510 B.n509 585
R603 B.n507 B.n58 585
R604 B.n58 B.n57 585
R605 B.n506 B.n505 585
R606 B.n505 B.n504 585
R607 B.n60 B.n59 585
R608 B.n503 B.n60 585
R609 B.n501 B.n500 585
R610 B.n502 B.n501 585
R611 B.n499 B.n65 585
R612 B.n65 B.n64 585
R613 B.n498 B.n497 585
R614 B.n497 B.n496 585
R615 B.n67 B.n66 585
R616 B.n495 B.n67 585
R617 B.n570 B.n569 585
R618 B.n568 B.n2 585
R619 B.n92 B.n67 521.33
R620 B.n492 B.n69 521.33
R621 B.n328 B.n233 521.33
R622 B.n325 B.n231 521.33
R623 B.n494 B.n493 256.663
R624 B.n494 B.n86 256.663
R625 B.n494 B.n85 256.663
R626 B.n494 B.n84 256.663
R627 B.n494 B.n83 256.663
R628 B.n494 B.n82 256.663
R629 B.n494 B.n81 256.663
R630 B.n494 B.n80 256.663
R631 B.n494 B.n79 256.663
R632 B.n494 B.n78 256.663
R633 B.n494 B.n77 256.663
R634 B.n494 B.n76 256.663
R635 B.n494 B.n75 256.663
R636 B.n494 B.n74 256.663
R637 B.n494 B.n73 256.663
R638 B.n494 B.n72 256.663
R639 B.n494 B.n71 256.663
R640 B.n494 B.n70 256.663
R641 B.n327 B.n326 256.663
R642 B.n327 B.n236 256.663
R643 B.n327 B.n237 256.663
R644 B.n327 B.n238 256.663
R645 B.n327 B.n239 256.663
R646 B.n327 B.n240 256.663
R647 B.n327 B.n241 256.663
R648 B.n327 B.n242 256.663
R649 B.n327 B.n243 256.663
R650 B.n327 B.n244 256.663
R651 B.n327 B.n245 256.663
R652 B.n327 B.n246 256.663
R653 B.n327 B.n247 256.663
R654 B.n327 B.n248 256.663
R655 B.n327 B.n249 256.663
R656 B.n327 B.n250 256.663
R657 B.n327 B.n251 256.663
R658 B.n572 B.n571 256.663
R659 B.n90 B.t17 248.597
R660 B.n88 B.t21 248.597
R661 B.n257 B.t14 248.597
R662 B.n254 B.t10 248.597
R663 B.n327 B.n232 167.251
R664 B.n495 B.n494 167.251
R665 B.n96 B.n95 163.367
R666 B.n100 B.n99 163.367
R667 B.n104 B.n103 163.367
R668 B.n108 B.n107 163.367
R669 B.n112 B.n111 163.367
R670 B.n116 B.n115 163.367
R671 B.n121 B.n120 163.367
R672 B.n125 B.n124 163.367
R673 B.n129 B.n128 163.367
R674 B.n133 B.n132 163.367
R675 B.n137 B.n136 163.367
R676 B.n142 B.n141 163.367
R677 B.n146 B.n145 163.367
R678 B.n150 B.n149 163.367
R679 B.n154 B.n153 163.367
R680 B.n158 B.n157 163.367
R681 B.n160 B.n87 163.367
R682 B.n332 B.n233 163.367
R683 B.n332 B.n227 163.367
R684 B.n340 B.n227 163.367
R685 B.n340 B.n225 163.367
R686 B.n344 B.n225 163.367
R687 B.n344 B.n219 163.367
R688 B.n352 B.n219 163.367
R689 B.n352 B.n217 163.367
R690 B.n356 B.n217 163.367
R691 B.n356 B.n211 163.367
R692 B.n364 B.n211 163.367
R693 B.n364 B.n209 163.367
R694 B.n368 B.n209 163.367
R695 B.n368 B.n203 163.367
R696 B.n376 B.n203 163.367
R697 B.n376 B.n201 163.367
R698 B.n380 B.n201 163.367
R699 B.n380 B.n196 163.367
R700 B.n389 B.n196 163.367
R701 B.n389 B.n194 163.367
R702 B.n393 B.n194 163.367
R703 B.n393 B.n188 163.367
R704 B.n401 B.n188 163.367
R705 B.n401 B.n186 163.367
R706 B.n405 B.n186 163.367
R707 B.n405 B.n179 163.367
R708 B.n413 B.n179 163.367
R709 B.n413 B.n177 163.367
R710 B.n417 B.n177 163.367
R711 B.n417 B.n172 163.367
R712 B.n425 B.n172 163.367
R713 B.n425 B.n170 163.367
R714 B.n430 B.n170 163.367
R715 B.n430 B.n164 163.367
R716 B.n438 B.n164 163.367
R717 B.n439 B.n438 163.367
R718 B.n439 B.n5 163.367
R719 B.n6 B.n5 163.367
R720 B.n7 B.n6 163.367
R721 B.n445 B.n7 163.367
R722 B.n447 B.n445 163.367
R723 B.n447 B.n12 163.367
R724 B.n13 B.n12 163.367
R725 B.n14 B.n13 163.367
R726 B.n452 B.n14 163.367
R727 B.n452 B.n19 163.367
R728 B.n20 B.n19 163.367
R729 B.n21 B.n20 163.367
R730 B.n457 B.n21 163.367
R731 B.n457 B.n26 163.367
R732 B.n27 B.n26 163.367
R733 B.n28 B.n27 163.367
R734 B.n462 B.n28 163.367
R735 B.n462 B.n33 163.367
R736 B.n34 B.n33 163.367
R737 B.n35 B.n34 163.367
R738 B.n467 B.n35 163.367
R739 B.n467 B.n40 163.367
R740 B.n41 B.n40 163.367
R741 B.n42 B.n41 163.367
R742 B.n472 B.n42 163.367
R743 B.n472 B.n47 163.367
R744 B.n48 B.n47 163.367
R745 B.n49 B.n48 163.367
R746 B.n477 B.n49 163.367
R747 B.n477 B.n54 163.367
R748 B.n55 B.n54 163.367
R749 B.n56 B.n55 163.367
R750 B.n482 B.n56 163.367
R751 B.n482 B.n61 163.367
R752 B.n62 B.n61 163.367
R753 B.n63 B.n62 163.367
R754 B.n487 B.n63 163.367
R755 B.n487 B.n68 163.367
R756 B.n69 B.n68 163.367
R757 B.n253 B.n252 163.367
R758 B.n320 B.n252 163.367
R759 B.n318 B.n317 163.367
R760 B.n314 B.n313 163.367
R761 B.n310 B.n309 163.367
R762 B.n306 B.n305 163.367
R763 B.n302 B.n301 163.367
R764 B.n298 B.n297 163.367
R765 B.n294 B.n293 163.367
R766 B.n290 B.n289 163.367
R767 B.n286 B.n285 163.367
R768 B.n282 B.n281 163.367
R769 B.n278 B.n277 163.367
R770 B.n274 B.n273 163.367
R771 B.n270 B.n269 163.367
R772 B.n266 B.n265 163.367
R773 B.n262 B.n261 163.367
R774 B.n328 B.n235 163.367
R775 B.n334 B.n231 163.367
R776 B.n334 B.n229 163.367
R777 B.n338 B.n229 163.367
R778 B.n338 B.n223 163.367
R779 B.n346 B.n223 163.367
R780 B.n346 B.n221 163.367
R781 B.n350 B.n221 163.367
R782 B.n350 B.n215 163.367
R783 B.n358 B.n215 163.367
R784 B.n358 B.n213 163.367
R785 B.n362 B.n213 163.367
R786 B.n362 B.n207 163.367
R787 B.n370 B.n207 163.367
R788 B.n370 B.n205 163.367
R789 B.n374 B.n205 163.367
R790 B.n374 B.n199 163.367
R791 B.n383 B.n199 163.367
R792 B.n383 B.n197 163.367
R793 B.n387 B.n197 163.367
R794 B.n387 B.n192 163.367
R795 B.n395 B.n192 163.367
R796 B.n395 B.n190 163.367
R797 B.n399 B.n190 163.367
R798 B.n399 B.n184 163.367
R799 B.n407 B.n184 163.367
R800 B.n407 B.n182 163.367
R801 B.n411 B.n182 163.367
R802 B.n411 B.n176 163.367
R803 B.n419 B.n176 163.367
R804 B.n419 B.n174 163.367
R805 B.n423 B.n174 163.367
R806 B.n423 B.n168 163.367
R807 B.n432 B.n168 163.367
R808 B.n432 B.n166 163.367
R809 B.n436 B.n166 163.367
R810 B.n436 B.n3 163.367
R811 B.n570 B.n3 163.367
R812 B.n566 B.n2 163.367
R813 B.n566 B.n565 163.367
R814 B.n565 B.n9 163.367
R815 B.n561 B.n9 163.367
R816 B.n561 B.n11 163.367
R817 B.n557 B.n11 163.367
R818 B.n557 B.n16 163.367
R819 B.n553 B.n16 163.367
R820 B.n553 B.n18 163.367
R821 B.n549 B.n18 163.367
R822 B.n549 B.n23 163.367
R823 B.n545 B.n23 163.367
R824 B.n545 B.n25 163.367
R825 B.n541 B.n25 163.367
R826 B.n541 B.n30 163.367
R827 B.n537 B.n30 163.367
R828 B.n537 B.n32 163.367
R829 B.n533 B.n32 163.367
R830 B.n533 B.n36 163.367
R831 B.n529 B.n36 163.367
R832 B.n529 B.n38 163.367
R833 B.n525 B.n38 163.367
R834 B.n525 B.n44 163.367
R835 B.n521 B.n44 163.367
R836 B.n521 B.n46 163.367
R837 B.n517 B.n46 163.367
R838 B.n517 B.n51 163.367
R839 B.n513 B.n51 163.367
R840 B.n513 B.n53 163.367
R841 B.n509 B.n53 163.367
R842 B.n509 B.n58 163.367
R843 B.n505 B.n58 163.367
R844 B.n505 B.n60 163.367
R845 B.n501 B.n60 163.367
R846 B.n501 B.n65 163.367
R847 B.n497 B.n65 163.367
R848 B.n497 B.n67 163.367
R849 B.n88 B.t22 153.341
R850 B.n257 B.t16 153.341
R851 B.n90 B.t19 153.341
R852 B.n254 B.t13 153.341
R853 B.n89 B.t23 121.147
R854 B.n258 B.t15 121.147
R855 B.n91 B.t20 121.147
R856 B.n255 B.t12 121.147
R857 B.n333 B.n232 97.2065
R858 B.n333 B.n228 97.2065
R859 B.n339 B.n228 97.2065
R860 B.n339 B.n224 97.2065
R861 B.n345 B.n224 97.2065
R862 B.n351 B.n220 97.2065
R863 B.n351 B.n216 97.2065
R864 B.n357 B.n216 97.2065
R865 B.n357 B.n212 97.2065
R866 B.n363 B.n212 97.2065
R867 B.n363 B.n208 97.2065
R868 B.n369 B.n208 97.2065
R869 B.n375 B.n204 97.2065
R870 B.n375 B.n200 97.2065
R871 B.n382 B.n200 97.2065
R872 B.n382 B.n381 97.2065
R873 B.n388 B.n193 97.2065
R874 B.n394 B.n193 97.2065
R875 B.n394 B.n189 97.2065
R876 B.n400 B.n189 97.2065
R877 B.n406 B.n185 97.2065
R878 B.n406 B.n180 97.2065
R879 B.n412 B.n180 97.2065
R880 B.n412 B.n181 97.2065
R881 B.n418 B.n173 97.2065
R882 B.n424 B.n173 97.2065
R883 B.n424 B.n169 97.2065
R884 B.n431 B.n169 97.2065
R885 B.n437 B.n165 97.2065
R886 B.n437 B.n4 97.2065
R887 B.n569 B.n4 97.2065
R888 B.n569 B.n568 97.2065
R889 B.n568 B.n567 97.2065
R890 B.n567 B.n8 97.2065
R891 B.n446 B.n8 97.2065
R892 B.n560 B.n559 97.2065
R893 B.n559 B.n558 97.2065
R894 B.n558 B.n15 97.2065
R895 B.n552 B.n15 97.2065
R896 B.n551 B.n550 97.2065
R897 B.n550 B.n22 97.2065
R898 B.n544 B.n22 97.2065
R899 B.n544 B.n543 97.2065
R900 B.n542 B.n29 97.2065
R901 B.n536 B.n29 97.2065
R902 B.n536 B.n535 97.2065
R903 B.n535 B.n534 97.2065
R904 B.n528 B.n39 97.2065
R905 B.n528 B.n527 97.2065
R906 B.n527 B.n526 97.2065
R907 B.n526 B.n43 97.2065
R908 B.n520 B.n519 97.2065
R909 B.n519 B.n518 97.2065
R910 B.n518 B.n50 97.2065
R911 B.n512 B.n50 97.2065
R912 B.n512 B.n511 97.2065
R913 B.n511 B.n510 97.2065
R914 B.n510 B.n57 97.2065
R915 B.n504 B.n503 97.2065
R916 B.n503 B.n502 97.2065
R917 B.n502 B.n64 97.2065
R918 B.n496 B.n64 97.2065
R919 B.n496 B.n495 97.2065
R920 B.n369 B.t5 90.059
R921 B.n520 B.t7 90.059
R922 B.n345 B.t11 81.482
R923 B.n504 B.t18 81.482
R924 B.n381 B.t0 78.623
R925 B.n39 B.t2 78.623
R926 B.n92 B.n70 71.676
R927 B.n96 B.n71 71.676
R928 B.n100 B.n72 71.676
R929 B.n104 B.n73 71.676
R930 B.n108 B.n74 71.676
R931 B.n112 B.n75 71.676
R932 B.n116 B.n76 71.676
R933 B.n121 B.n77 71.676
R934 B.n125 B.n78 71.676
R935 B.n129 B.n79 71.676
R936 B.n133 B.n80 71.676
R937 B.n137 B.n81 71.676
R938 B.n142 B.n82 71.676
R939 B.n146 B.n83 71.676
R940 B.n150 B.n84 71.676
R941 B.n154 B.n85 71.676
R942 B.n158 B.n86 71.676
R943 B.n493 B.n87 71.676
R944 B.n493 B.n492 71.676
R945 B.n160 B.n86 71.676
R946 B.n157 B.n85 71.676
R947 B.n153 B.n84 71.676
R948 B.n149 B.n83 71.676
R949 B.n145 B.n82 71.676
R950 B.n141 B.n81 71.676
R951 B.n136 B.n80 71.676
R952 B.n132 B.n79 71.676
R953 B.n128 B.n78 71.676
R954 B.n124 B.n77 71.676
R955 B.n120 B.n76 71.676
R956 B.n115 B.n75 71.676
R957 B.n111 B.n74 71.676
R958 B.n107 B.n73 71.676
R959 B.n103 B.n72 71.676
R960 B.n99 B.n71 71.676
R961 B.n95 B.n70 71.676
R962 B.n326 B.n325 71.676
R963 B.n320 B.n236 71.676
R964 B.n317 B.n237 71.676
R965 B.n313 B.n238 71.676
R966 B.n309 B.n239 71.676
R967 B.n305 B.n240 71.676
R968 B.n301 B.n241 71.676
R969 B.n297 B.n242 71.676
R970 B.n293 B.n243 71.676
R971 B.n289 B.n244 71.676
R972 B.n285 B.n245 71.676
R973 B.n281 B.n246 71.676
R974 B.n277 B.n247 71.676
R975 B.n273 B.n248 71.676
R976 B.n269 B.n249 71.676
R977 B.n265 B.n250 71.676
R978 B.n261 B.n251 71.676
R979 B.n326 B.n253 71.676
R980 B.n318 B.n236 71.676
R981 B.n314 B.n237 71.676
R982 B.n310 B.n238 71.676
R983 B.n306 B.n239 71.676
R984 B.n302 B.n240 71.676
R985 B.n298 B.n241 71.676
R986 B.n294 B.n242 71.676
R987 B.n290 B.n243 71.676
R988 B.n286 B.n244 71.676
R989 B.n282 B.n245 71.676
R990 B.n278 B.n246 71.676
R991 B.n274 B.n247 71.676
R992 B.n270 B.n248 71.676
R993 B.n266 B.n249 71.676
R994 B.n262 B.n250 71.676
R995 B.n251 B.n235 71.676
R996 B.n571 B.n570 71.676
R997 B.n571 B.n2 71.676
R998 B.n400 B.t4 67.187
R999 B.t1 B.n542 67.187
R1000 B.n118 B.n91 59.5399
R1001 B.n139 B.n89 59.5399
R1002 B.n259 B.n258 59.5399
R1003 B.n256 B.n255 59.5399
R1004 B.n181 B.t8 55.751
R1005 B.t9 B.n551 55.751
R1006 B.t3 B.n165 52.892
R1007 B.n446 B.t6 52.892
R1008 B.n431 B.t3 44.315
R1009 B.n560 B.t6 44.315
R1010 B.n418 B.t8 41.456
R1011 B.n552 B.t9 41.456
R1012 B.n324 B.n230 33.8737
R1013 B.n330 B.n329 33.8737
R1014 B.n491 B.n490 33.8737
R1015 B.n93 B.n66 33.8737
R1016 B.n91 B.n90 32.1944
R1017 B.n89 B.n88 32.1944
R1018 B.n258 B.n257 32.1944
R1019 B.n255 B.n254 32.1944
R1020 B.t4 B.n185 30.02
R1021 B.n543 B.t1 30.02
R1022 B.n388 B.t0 18.584
R1023 B.n534 B.t2 18.584
R1024 B B.n572 18.0485
R1025 B.t11 B.n220 15.725
R1026 B.t18 B.n57 15.725
R1027 B.n335 B.n230 10.6151
R1028 B.n336 B.n335 10.6151
R1029 B.n337 B.n336 10.6151
R1030 B.n337 B.n222 10.6151
R1031 B.n347 B.n222 10.6151
R1032 B.n348 B.n347 10.6151
R1033 B.n349 B.n348 10.6151
R1034 B.n349 B.n214 10.6151
R1035 B.n359 B.n214 10.6151
R1036 B.n360 B.n359 10.6151
R1037 B.n361 B.n360 10.6151
R1038 B.n361 B.n206 10.6151
R1039 B.n371 B.n206 10.6151
R1040 B.n372 B.n371 10.6151
R1041 B.n373 B.n372 10.6151
R1042 B.n373 B.n198 10.6151
R1043 B.n384 B.n198 10.6151
R1044 B.n385 B.n384 10.6151
R1045 B.n386 B.n385 10.6151
R1046 B.n386 B.n191 10.6151
R1047 B.n396 B.n191 10.6151
R1048 B.n397 B.n396 10.6151
R1049 B.n398 B.n397 10.6151
R1050 B.n398 B.n183 10.6151
R1051 B.n408 B.n183 10.6151
R1052 B.n409 B.n408 10.6151
R1053 B.n410 B.n409 10.6151
R1054 B.n410 B.n175 10.6151
R1055 B.n420 B.n175 10.6151
R1056 B.n421 B.n420 10.6151
R1057 B.n422 B.n421 10.6151
R1058 B.n422 B.n167 10.6151
R1059 B.n433 B.n167 10.6151
R1060 B.n434 B.n433 10.6151
R1061 B.n435 B.n434 10.6151
R1062 B.n435 B.n0 10.6151
R1063 B.n324 B.n323 10.6151
R1064 B.n323 B.n322 10.6151
R1065 B.n322 B.n321 10.6151
R1066 B.n321 B.n319 10.6151
R1067 B.n319 B.n316 10.6151
R1068 B.n316 B.n315 10.6151
R1069 B.n315 B.n312 10.6151
R1070 B.n312 B.n311 10.6151
R1071 B.n311 B.n308 10.6151
R1072 B.n308 B.n307 10.6151
R1073 B.n307 B.n304 10.6151
R1074 B.n304 B.n303 10.6151
R1075 B.n300 B.n299 10.6151
R1076 B.n299 B.n296 10.6151
R1077 B.n296 B.n295 10.6151
R1078 B.n295 B.n292 10.6151
R1079 B.n292 B.n291 10.6151
R1080 B.n291 B.n288 10.6151
R1081 B.n288 B.n287 10.6151
R1082 B.n287 B.n284 10.6151
R1083 B.n284 B.n283 10.6151
R1084 B.n280 B.n279 10.6151
R1085 B.n279 B.n276 10.6151
R1086 B.n276 B.n275 10.6151
R1087 B.n275 B.n272 10.6151
R1088 B.n272 B.n271 10.6151
R1089 B.n271 B.n268 10.6151
R1090 B.n268 B.n267 10.6151
R1091 B.n267 B.n264 10.6151
R1092 B.n264 B.n263 10.6151
R1093 B.n263 B.n260 10.6151
R1094 B.n260 B.n234 10.6151
R1095 B.n329 B.n234 10.6151
R1096 B.n331 B.n330 10.6151
R1097 B.n331 B.n226 10.6151
R1098 B.n341 B.n226 10.6151
R1099 B.n342 B.n341 10.6151
R1100 B.n343 B.n342 10.6151
R1101 B.n343 B.n218 10.6151
R1102 B.n353 B.n218 10.6151
R1103 B.n354 B.n353 10.6151
R1104 B.n355 B.n354 10.6151
R1105 B.n355 B.n210 10.6151
R1106 B.n365 B.n210 10.6151
R1107 B.n366 B.n365 10.6151
R1108 B.n367 B.n366 10.6151
R1109 B.n367 B.n202 10.6151
R1110 B.n377 B.n202 10.6151
R1111 B.n378 B.n377 10.6151
R1112 B.n379 B.n378 10.6151
R1113 B.n379 B.n195 10.6151
R1114 B.n390 B.n195 10.6151
R1115 B.n391 B.n390 10.6151
R1116 B.n392 B.n391 10.6151
R1117 B.n392 B.n187 10.6151
R1118 B.n402 B.n187 10.6151
R1119 B.n403 B.n402 10.6151
R1120 B.n404 B.n403 10.6151
R1121 B.n404 B.n178 10.6151
R1122 B.n414 B.n178 10.6151
R1123 B.n415 B.n414 10.6151
R1124 B.n416 B.n415 10.6151
R1125 B.n416 B.n171 10.6151
R1126 B.n426 B.n171 10.6151
R1127 B.n427 B.n426 10.6151
R1128 B.n429 B.n427 10.6151
R1129 B.n429 B.n428 10.6151
R1130 B.n428 B.n163 10.6151
R1131 B.n440 B.n163 10.6151
R1132 B.n441 B.n440 10.6151
R1133 B.n442 B.n441 10.6151
R1134 B.n443 B.n442 10.6151
R1135 B.n444 B.n443 10.6151
R1136 B.n448 B.n444 10.6151
R1137 B.n449 B.n448 10.6151
R1138 B.n450 B.n449 10.6151
R1139 B.n451 B.n450 10.6151
R1140 B.n453 B.n451 10.6151
R1141 B.n454 B.n453 10.6151
R1142 B.n455 B.n454 10.6151
R1143 B.n456 B.n455 10.6151
R1144 B.n458 B.n456 10.6151
R1145 B.n459 B.n458 10.6151
R1146 B.n460 B.n459 10.6151
R1147 B.n461 B.n460 10.6151
R1148 B.n463 B.n461 10.6151
R1149 B.n464 B.n463 10.6151
R1150 B.n465 B.n464 10.6151
R1151 B.n466 B.n465 10.6151
R1152 B.n468 B.n466 10.6151
R1153 B.n469 B.n468 10.6151
R1154 B.n470 B.n469 10.6151
R1155 B.n471 B.n470 10.6151
R1156 B.n473 B.n471 10.6151
R1157 B.n474 B.n473 10.6151
R1158 B.n475 B.n474 10.6151
R1159 B.n476 B.n475 10.6151
R1160 B.n478 B.n476 10.6151
R1161 B.n479 B.n478 10.6151
R1162 B.n480 B.n479 10.6151
R1163 B.n481 B.n480 10.6151
R1164 B.n483 B.n481 10.6151
R1165 B.n484 B.n483 10.6151
R1166 B.n485 B.n484 10.6151
R1167 B.n486 B.n485 10.6151
R1168 B.n488 B.n486 10.6151
R1169 B.n489 B.n488 10.6151
R1170 B.n490 B.n489 10.6151
R1171 B.n564 B.n1 10.6151
R1172 B.n564 B.n563 10.6151
R1173 B.n563 B.n562 10.6151
R1174 B.n562 B.n10 10.6151
R1175 B.n556 B.n10 10.6151
R1176 B.n556 B.n555 10.6151
R1177 B.n555 B.n554 10.6151
R1178 B.n554 B.n17 10.6151
R1179 B.n548 B.n17 10.6151
R1180 B.n548 B.n547 10.6151
R1181 B.n547 B.n546 10.6151
R1182 B.n546 B.n24 10.6151
R1183 B.n540 B.n24 10.6151
R1184 B.n540 B.n539 10.6151
R1185 B.n539 B.n538 10.6151
R1186 B.n538 B.n31 10.6151
R1187 B.n532 B.n31 10.6151
R1188 B.n532 B.n531 10.6151
R1189 B.n531 B.n530 10.6151
R1190 B.n530 B.n37 10.6151
R1191 B.n524 B.n37 10.6151
R1192 B.n524 B.n523 10.6151
R1193 B.n523 B.n522 10.6151
R1194 B.n522 B.n45 10.6151
R1195 B.n516 B.n45 10.6151
R1196 B.n516 B.n515 10.6151
R1197 B.n515 B.n514 10.6151
R1198 B.n514 B.n52 10.6151
R1199 B.n508 B.n52 10.6151
R1200 B.n508 B.n507 10.6151
R1201 B.n507 B.n506 10.6151
R1202 B.n506 B.n59 10.6151
R1203 B.n500 B.n59 10.6151
R1204 B.n500 B.n499 10.6151
R1205 B.n499 B.n498 10.6151
R1206 B.n498 B.n66 10.6151
R1207 B.n94 B.n93 10.6151
R1208 B.n97 B.n94 10.6151
R1209 B.n98 B.n97 10.6151
R1210 B.n101 B.n98 10.6151
R1211 B.n102 B.n101 10.6151
R1212 B.n105 B.n102 10.6151
R1213 B.n106 B.n105 10.6151
R1214 B.n109 B.n106 10.6151
R1215 B.n110 B.n109 10.6151
R1216 B.n113 B.n110 10.6151
R1217 B.n114 B.n113 10.6151
R1218 B.n117 B.n114 10.6151
R1219 B.n122 B.n119 10.6151
R1220 B.n123 B.n122 10.6151
R1221 B.n126 B.n123 10.6151
R1222 B.n127 B.n126 10.6151
R1223 B.n130 B.n127 10.6151
R1224 B.n131 B.n130 10.6151
R1225 B.n134 B.n131 10.6151
R1226 B.n135 B.n134 10.6151
R1227 B.n138 B.n135 10.6151
R1228 B.n143 B.n140 10.6151
R1229 B.n144 B.n143 10.6151
R1230 B.n147 B.n144 10.6151
R1231 B.n148 B.n147 10.6151
R1232 B.n151 B.n148 10.6151
R1233 B.n152 B.n151 10.6151
R1234 B.n155 B.n152 10.6151
R1235 B.n156 B.n155 10.6151
R1236 B.n159 B.n156 10.6151
R1237 B.n161 B.n159 10.6151
R1238 B.n162 B.n161 10.6151
R1239 B.n491 B.n162 10.6151
R1240 B.n303 B.n256 9.36635
R1241 B.n280 B.n259 9.36635
R1242 B.n118 B.n117 9.36635
R1243 B.n140 B.n139 9.36635
R1244 B.n572 B.n0 8.11757
R1245 B.n572 B.n1 8.11757
R1246 B.t5 B.n204 7.148
R1247 B.t7 B.n43 7.148
R1248 B.n300 B.n256 1.24928
R1249 B.n283 B.n259 1.24928
R1250 B.n119 B.n118 1.24928
R1251 B.n139 B.n138 1.24928
R1252 VP.n33 VP.n7 170.154
R1253 VP.n56 VP.n55 170.154
R1254 VP.n32 VP.n31 170.154
R1255 VP.n16 VP.n15 161.3
R1256 VP.n17 VP.n12 161.3
R1257 VP.n19 VP.n18 161.3
R1258 VP.n20 VP.n11 161.3
R1259 VP.n22 VP.n21 161.3
R1260 VP.n23 VP.n10 161.3
R1261 VP.n26 VP.n25 161.3
R1262 VP.n27 VP.n9 161.3
R1263 VP.n29 VP.n28 161.3
R1264 VP.n30 VP.n8 161.3
R1265 VP.n54 VP.n0 161.3
R1266 VP.n53 VP.n52 161.3
R1267 VP.n51 VP.n1 161.3
R1268 VP.n50 VP.n49 161.3
R1269 VP.n47 VP.n2 161.3
R1270 VP.n46 VP.n45 161.3
R1271 VP.n44 VP.n3 161.3
R1272 VP.n43 VP.n42 161.3
R1273 VP.n41 VP.n4 161.3
R1274 VP.n40 VP.n39 161.3
R1275 VP.n38 VP.n37 161.3
R1276 VP.n36 VP.n6 161.3
R1277 VP.n35 VP.n34 161.3
R1278 VP.n14 VP.t5 75.5805
R1279 VP.n14 VP.n13 56.6996
R1280 VP.n42 VP.n41 56.5617
R1281 VP.n47 VP.n46 56.5617
R1282 VP.n23 VP.n22 56.5617
R1283 VP.n18 VP.n17 56.5617
R1284 VP.n3 VP.t2 43.8516
R1285 VP.n7 VP.t1 43.8516
R1286 VP.n5 VP.t0 43.8516
R1287 VP.n48 VP.t6 43.8516
R1288 VP.n55 VP.t7 43.8516
R1289 VP.n11 VP.t9 43.8516
R1290 VP.n31 VP.t4 43.8516
R1291 VP.n24 VP.t8 43.8516
R1292 VP.n13 VP.t3 43.8516
R1293 VP.n37 VP.n36 41.5458
R1294 VP.n53 VP.n1 41.5458
R1295 VP.n29 VP.n9 41.5458
R1296 VP.n36 VP.n35 39.6083
R1297 VP.n54 VP.n53 39.6083
R1298 VP.n30 VP.n29 39.6083
R1299 VP.n33 VP.n32 38.9247
R1300 VP.n15 VP.n14 26.5036
R1301 VP.n41 VP.n40 24.5923
R1302 VP.n42 VP.n3 24.5923
R1303 VP.n46 VP.n3 24.5923
R1304 VP.n49 VP.n47 24.5923
R1305 VP.n25 VP.n23 24.5923
R1306 VP.n18 VP.n11 24.5923
R1307 VP.n22 VP.n11 24.5923
R1308 VP.n17 VP.n16 24.5923
R1309 VP.n37 VP.n5 16.7229
R1310 VP.n48 VP.n1 16.7229
R1311 VP.n24 VP.n9 16.7229
R1312 VP.n35 VP.n7 15.7393
R1313 VP.n55 VP.n54 15.7393
R1314 VP.n31 VP.n30 15.7393
R1315 VP.n40 VP.n5 7.86989
R1316 VP.n49 VP.n48 7.86989
R1317 VP.n25 VP.n24 7.86989
R1318 VP.n16 VP.n13 7.86989
R1319 VP.n15 VP.n12 0.189894
R1320 VP.n19 VP.n12 0.189894
R1321 VP.n20 VP.n19 0.189894
R1322 VP.n21 VP.n20 0.189894
R1323 VP.n21 VP.n10 0.189894
R1324 VP.n26 VP.n10 0.189894
R1325 VP.n27 VP.n26 0.189894
R1326 VP.n28 VP.n27 0.189894
R1327 VP.n28 VP.n8 0.189894
R1328 VP.n32 VP.n8 0.189894
R1329 VP.n34 VP.n33 0.189894
R1330 VP.n34 VP.n6 0.189894
R1331 VP.n38 VP.n6 0.189894
R1332 VP.n39 VP.n38 0.189894
R1333 VP.n39 VP.n4 0.189894
R1334 VP.n43 VP.n4 0.189894
R1335 VP.n44 VP.n43 0.189894
R1336 VP.n45 VP.n44 0.189894
R1337 VP.n45 VP.n2 0.189894
R1338 VP.n50 VP.n2 0.189894
R1339 VP.n51 VP.n50 0.189894
R1340 VP.n52 VP.n51 0.189894
R1341 VP.n52 VP.n0 0.189894
R1342 VP.n56 VP.n0 0.189894
R1343 VP VP.n56 0.0516364
R1344 VDD1.n6 VDD1.n0 289.615
R1345 VDD1.n19 VDD1.n13 289.615
R1346 VDD1.n7 VDD1.n6 185
R1347 VDD1.n5 VDD1.n4 185
R1348 VDD1.n18 VDD1.n17 185
R1349 VDD1.n20 VDD1.n19 185
R1350 VDD1.n3 VDD1.t4 151.613
R1351 VDD1.n16 VDD1.t8 151.613
R1352 VDD1.n6 VDD1.n5 104.615
R1353 VDD1.n19 VDD1.n18 104.615
R1354 VDD1.n27 VDD1.n26 86.365
R1355 VDD1.n12 VDD1.n11 85.3472
R1356 VDD1.n29 VDD1.n28 85.3471
R1357 VDD1.n25 VDD1.n24 85.3471
R1358 VDD1.n5 VDD1.t4 52.3082
R1359 VDD1.n18 VDD1.t8 52.3082
R1360 VDD1.n12 VDD1.n10 50.6831
R1361 VDD1.n25 VDD1.n23 50.6831
R1362 VDD1.n29 VDD1.n27 33.8974
R1363 VDD1.n4 VDD1.n3 15.3979
R1364 VDD1.n17 VDD1.n16 15.3979
R1365 VDD1.n7 VDD1.n2 12.8005
R1366 VDD1.n20 VDD1.n15 12.8005
R1367 VDD1.n8 VDD1.n0 12.0247
R1368 VDD1.n21 VDD1.n13 12.0247
R1369 VDD1.n10 VDD1.n9 9.45567
R1370 VDD1.n23 VDD1.n22 9.45567
R1371 VDD1.n9 VDD1.n8 9.3005
R1372 VDD1.n2 VDD1.n1 9.3005
R1373 VDD1.n22 VDD1.n21 9.3005
R1374 VDD1.n15 VDD1.n14 9.3005
R1375 VDD1.n28 VDD1.t1 8.18232
R1376 VDD1.n28 VDD1.t5 8.18232
R1377 VDD1.n11 VDD1.t6 8.18232
R1378 VDD1.n11 VDD1.t0 8.18232
R1379 VDD1.n26 VDD1.t3 8.18232
R1380 VDD1.n26 VDD1.t2 8.18232
R1381 VDD1.n24 VDD1.t9 8.18232
R1382 VDD1.n24 VDD1.t7 8.18232
R1383 VDD1.n3 VDD1.n1 4.69785
R1384 VDD1.n16 VDD1.n14 4.69785
R1385 VDD1.n10 VDD1.n0 1.93989
R1386 VDD1.n23 VDD1.n13 1.93989
R1387 VDD1.n8 VDD1.n7 1.16414
R1388 VDD1.n21 VDD1.n20 1.16414
R1389 VDD1 VDD1.n29 1.01559
R1390 VDD1 VDD1.n12 0.416448
R1391 VDD1.n4 VDD1.n2 0.388379
R1392 VDD1.n17 VDD1.n15 0.388379
R1393 VDD1.n27 VDD1.n25 0.302913
R1394 VDD1.n9 VDD1.n1 0.155672
R1395 VDD1.n22 VDD1.n14 0.155672
C0 VDD2 VTAIL 4.9293f
C1 VDD2 VP 0.427443f
C2 VDD2 VN 2.17275f
C3 VTAIL VDD1 4.88512f
C4 VDD1 VP 2.44114f
C5 VTAIL VP 2.86079f
C6 VDD1 VN 0.156513f
C7 VTAIL VN 2.84662f
C8 VDD2 VDD1 1.34863f
C9 VN VP 4.75327f
C10 VDD2 B 3.99639f
C11 VDD1 B 3.970054f
C12 VTAIL B 3.195377f
C13 VN B 11.211711f
C14 VP B 9.68928f
C15 VDD1.n0 B 0.030624f
C16 VDD1.n1 B 0.172947f
C17 VDD1.n2 B 0.012815f
C18 VDD1.t4 B 0.051512f
C19 VDD1.n3 B 0.082166f
C20 VDD1.n4 B 0.017146f
C21 VDD1.n5 B 0.022717f
C22 VDD1.n6 B 0.06045f
C23 VDD1.n7 B 0.013568f
C24 VDD1.n8 B 0.012815f
C25 VDD1.n9 B 0.055774f
C26 VDD1.n10 B 0.054191f
C27 VDD1.t6 B 0.045605f
C28 VDD1.t0 B 0.045605f
C29 VDD1.n11 B 0.322509f
C30 VDD1.n12 B 0.465887f
C31 VDD1.n13 B 0.030624f
C32 VDD1.n14 B 0.172947f
C33 VDD1.n15 B 0.012815f
C34 VDD1.t8 B 0.051512f
C35 VDD1.n16 B 0.082166f
C36 VDD1.n17 B 0.017146f
C37 VDD1.n18 B 0.022717f
C38 VDD1.n19 B 0.06045f
C39 VDD1.n20 B 0.013568f
C40 VDD1.n21 B 0.012815f
C41 VDD1.n22 B 0.055774f
C42 VDD1.n23 B 0.054191f
C43 VDD1.t9 B 0.045605f
C44 VDD1.t7 B 0.045605f
C45 VDD1.n24 B 0.322507f
C46 VDD1.n25 B 0.458992f
C47 VDD1.t3 B 0.045605f
C48 VDD1.t2 B 0.045605f
C49 VDD1.n26 B 0.326874f
C50 VDD1.n27 B 1.65434f
C51 VDD1.t1 B 0.045605f
C52 VDD1.t5 B 0.045605f
C53 VDD1.n28 B 0.322507f
C54 VDD1.n29 B 1.77812f
C55 VP.n0 B 0.038479f
C56 VP.t7 B 0.299271f
C57 VP.n1 B 0.064395f
C58 VP.n2 B 0.038479f
C59 VP.t2 B 0.299271f
C60 VP.n3 B 0.187048f
C61 VP.n4 B 0.038479f
C62 VP.t0 B 0.299271f
C63 VP.n5 B 0.150919f
C64 VP.n6 B 0.038479f
C65 VP.t1 B 0.299271f
C66 VP.n7 B 0.228579f
C67 VP.n8 B 0.038479f
C68 VP.t4 B 0.299271f
C69 VP.n9 B 0.064395f
C70 VP.n10 B 0.038479f
C71 VP.t9 B 0.299271f
C72 VP.n11 B 0.187048f
C73 VP.n12 B 0.038479f
C74 VP.t3 B 0.299271f
C75 VP.n13 B 0.207549f
C76 VP.t5 B 0.416185f
C77 VP.n14 B 0.216343f
C78 VP.n15 B 0.205768f
C79 VP.n16 B 0.047401f
C80 VP.n17 B 0.047418f
C81 VP.n18 B 0.064451f
C82 VP.n19 B 0.038479f
C83 VP.n20 B 0.038479f
C84 VP.n21 B 0.038479f
C85 VP.n22 B 0.064451f
C86 VP.n23 B 0.047418f
C87 VP.t8 B 0.299271f
C88 VP.n24 B 0.150919f
C89 VP.n25 B 0.047401f
C90 VP.n26 B 0.038479f
C91 VP.n27 B 0.038479f
C92 VP.n28 B 0.038479f
C93 VP.n29 B 0.031127f
C94 VP.n30 B 0.063749f
C95 VP.n31 B 0.228579f
C96 VP.n32 B 1.39858f
C97 VP.n33 B 1.43422f
C98 VP.n34 B 0.038479f
C99 VP.n35 B 0.063749f
C100 VP.n36 B 0.031127f
C101 VP.n37 B 0.064395f
C102 VP.n38 B 0.038479f
C103 VP.n39 B 0.038479f
C104 VP.n40 B 0.047401f
C105 VP.n41 B 0.047418f
C106 VP.n42 B 0.064451f
C107 VP.n43 B 0.038479f
C108 VP.n44 B 0.038479f
C109 VP.n45 B 0.038479f
C110 VP.n46 B 0.064451f
C111 VP.n47 B 0.047418f
C112 VP.t6 B 0.299271f
C113 VP.n48 B 0.150919f
C114 VP.n49 B 0.047401f
C115 VP.n50 B 0.038479f
C116 VP.n51 B 0.038479f
C117 VP.n52 B 0.038479f
C118 VP.n53 B 0.031127f
C119 VP.n54 B 0.063749f
C120 VP.n55 B 0.228579f
C121 VP.n56 B 0.034082f
C122 VDD2.n0 B 0.030149f
C123 VDD2.n1 B 0.170263f
C124 VDD2.n2 B 0.012616f
C125 VDD2.t0 B 0.050712f
C126 VDD2.n3 B 0.080891f
C127 VDD2.n4 B 0.01688f
C128 VDD2.n5 B 0.022365f
C129 VDD2.n6 B 0.059512f
C130 VDD2.n7 B 0.013358f
C131 VDD2.n8 B 0.012616f
C132 VDD2.n9 B 0.054909f
C133 VDD2.n10 B 0.05335f
C134 VDD2.t1 B 0.044898f
C135 VDD2.t9 B 0.044898f
C136 VDD2.n11 B 0.317503f
C137 VDD2.n12 B 0.451869f
C138 VDD2.t3 B 0.044898f
C139 VDD2.t5 B 0.044898f
C140 VDD2.n13 B 0.321801f
C141 VDD2.n14 B 1.54812f
C142 VDD2.n15 B 0.030149f
C143 VDD2.n16 B 0.170263f
C144 VDD2.n17 B 0.012616f
C145 VDD2.t2 B 0.050712f
C146 VDD2.n18 B 0.080891f
C147 VDD2.n19 B 0.01688f
C148 VDD2.n20 B 0.022365f
C149 VDD2.n21 B 0.059512f
C150 VDD2.n22 B 0.013358f
C151 VDD2.n23 B 0.012616f
C152 VDD2.n24 B 0.054909f
C153 VDD2.n25 B 0.049006f
C154 VDD2.n26 B 1.53425f
C155 VDD2.t8 B 0.044898f
C156 VDD2.t7 B 0.044898f
C157 VDD2.n27 B 0.317504f
C158 VDD2.n28 B 0.309167f
C159 VDD2.t6 B 0.044898f
C160 VDD2.t4 B 0.044898f
C161 VDD2.n29 B 0.32178f
C162 VTAIL.t17 B 0.061499f
C163 VTAIL.t14 B 0.061499f
C164 VTAIL.n0 B 0.380013f
C165 VTAIL.n1 B 0.483347f
C166 VTAIL.n2 B 0.041296f
C167 VTAIL.n3 B 0.233219f
C168 VTAIL.n4 B 0.017281f
C169 VTAIL.t3 B 0.069463f
C170 VTAIL.n5 B 0.110801f
C171 VTAIL.n6 B 0.023122f
C172 VTAIL.n7 B 0.030634f
C173 VTAIL.n8 B 0.081516f
C174 VTAIL.n9 B 0.018297f
C175 VTAIL.n10 B 0.017281f
C176 VTAIL.n11 B 0.075212f
C177 VTAIL.n12 B 0.044929f
C178 VTAIL.n13 B 0.299076f
C179 VTAIL.t4 B 0.061499f
C180 VTAIL.t8 B 0.061499f
C181 VTAIL.n14 B 0.380013f
C182 VTAIL.n15 B 0.539848f
C183 VTAIL.t5 B 0.061499f
C184 VTAIL.t0 B 0.061499f
C185 VTAIL.n16 B 0.380013f
C186 VTAIL.n17 B 1.34115f
C187 VTAIL.t13 B 0.061499f
C188 VTAIL.t18 B 0.061499f
C189 VTAIL.n18 B 0.380016f
C190 VTAIL.n19 B 1.34115f
C191 VTAIL.t10 B 0.061499f
C192 VTAIL.t19 B 0.061499f
C193 VTAIL.n20 B 0.380016f
C194 VTAIL.n21 B 0.539845f
C195 VTAIL.n22 B 0.041296f
C196 VTAIL.n23 B 0.233219f
C197 VTAIL.n24 B 0.017281f
C198 VTAIL.t12 B 0.069463f
C199 VTAIL.n25 B 0.110801f
C200 VTAIL.n26 B 0.023122f
C201 VTAIL.n27 B 0.030634f
C202 VTAIL.n28 B 0.081516f
C203 VTAIL.n29 B 0.018297f
C204 VTAIL.n30 B 0.017281f
C205 VTAIL.n31 B 0.075212f
C206 VTAIL.n32 B 0.044929f
C207 VTAIL.n33 B 0.299076f
C208 VTAIL.t6 B 0.061499f
C209 VTAIL.t9 B 0.061499f
C210 VTAIL.n34 B 0.380016f
C211 VTAIL.n35 B 0.514386f
C212 VTAIL.t1 B 0.061499f
C213 VTAIL.t2 B 0.061499f
C214 VTAIL.n36 B 0.380016f
C215 VTAIL.n37 B 0.539845f
C216 VTAIL.n38 B 0.041296f
C217 VTAIL.n39 B 0.233219f
C218 VTAIL.n40 B 0.017281f
C219 VTAIL.t7 B 0.069463f
C220 VTAIL.n41 B 0.110801f
C221 VTAIL.n42 B 0.023122f
C222 VTAIL.n43 B 0.030634f
C223 VTAIL.n44 B 0.081516f
C224 VTAIL.n45 B 0.018297f
C225 VTAIL.n46 B 0.017281f
C226 VTAIL.n47 B 0.075212f
C227 VTAIL.n48 B 0.044929f
C228 VTAIL.n49 B 0.977548f
C229 VTAIL.n50 B 0.041296f
C230 VTAIL.n51 B 0.233219f
C231 VTAIL.n52 B 0.017281f
C232 VTAIL.t16 B 0.069463f
C233 VTAIL.n53 B 0.110801f
C234 VTAIL.n54 B 0.023122f
C235 VTAIL.n55 B 0.030634f
C236 VTAIL.n56 B 0.081516f
C237 VTAIL.n57 B 0.018297f
C238 VTAIL.n58 B 0.017281f
C239 VTAIL.n59 B 0.075212f
C240 VTAIL.n60 B 0.044929f
C241 VTAIL.n61 B 0.977548f
C242 VTAIL.t11 B 0.061499f
C243 VTAIL.t15 B 0.061499f
C244 VTAIL.n62 B 0.380013f
C245 VTAIL.n63 B 0.422603f
C246 VN.n0 B 0.037137f
C247 VN.t4 B 0.288835f
C248 VN.n1 B 0.06215f
C249 VN.n2 B 0.037137f
C250 VN.t0 B 0.288835f
C251 VN.n3 B 0.180525f
C252 VN.n4 B 0.037137f
C253 VN.t8 B 0.288835f
C254 VN.n5 B 0.200312f
C255 VN.t9 B 0.401672f
C256 VN.n6 B 0.208799f
C257 VN.n7 B 0.198592f
C258 VN.n8 B 0.045748f
C259 VN.n9 B 0.045764f
C260 VN.n10 B 0.062204f
C261 VN.n11 B 0.037137f
C262 VN.n12 B 0.037137f
C263 VN.n13 B 0.037137f
C264 VN.n14 B 0.062204f
C265 VN.n15 B 0.045764f
C266 VN.t6 B 0.288835f
C267 VN.n16 B 0.145656f
C268 VN.n17 B 0.045748f
C269 VN.n18 B 0.037137f
C270 VN.n19 B 0.037137f
C271 VN.n20 B 0.037137f
C272 VN.n21 B 0.030041f
C273 VN.n22 B 0.061526f
C274 VN.n23 B 0.220608f
C275 VN.n24 B 0.032893f
C276 VN.n25 B 0.037137f
C277 VN.t7 B 0.288835f
C278 VN.n26 B 0.06215f
C279 VN.n27 B 0.037137f
C280 VN.t1 B 0.288835f
C281 VN.n28 B 0.145656f
C282 VN.t2 B 0.288835f
C283 VN.n29 B 0.180525f
C284 VN.n30 B 0.037137f
C285 VN.t3 B 0.288835f
C286 VN.n31 B 0.200312f
C287 VN.t5 B 0.401672f
C288 VN.n32 B 0.208799f
C289 VN.n33 B 0.198592f
C290 VN.n34 B 0.045748f
C291 VN.n35 B 0.045764f
C292 VN.n36 B 0.062204f
C293 VN.n37 B 0.037137f
C294 VN.n38 B 0.037137f
C295 VN.n39 B 0.037137f
C296 VN.n40 B 0.062204f
C297 VN.n41 B 0.045764f
C298 VN.n42 B 0.045748f
C299 VN.n43 B 0.037137f
C300 VN.n44 B 0.037137f
C301 VN.n45 B 0.037137f
C302 VN.n46 B 0.030041f
C303 VN.n47 B 0.061526f
C304 VN.n48 B 0.220608f
C305 VN.n49 B 1.37431f
.ends

