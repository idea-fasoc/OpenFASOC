* NGSPICE file created from diff_pair_sample_0164.ext - technology: sky130A

.subckt diff_pair_sample_0164 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t3 sky130_fd_pr__nfet_01v8 ad=2.6403 pd=14.32 as=0 ps=0 w=6.77 l=2.74
X1 VDD1.t1 VP.t0 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=2.6403 pd=14.32 as=2.6403 ps=14.32 w=6.77 l=2.74
X2 VDD1.t0 VP.t1 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=2.6403 pd=14.32 as=2.6403 ps=14.32 w=6.77 l=2.74
X3 VDD2.t1 VN.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.6403 pd=14.32 as=2.6403 ps=14.32 w=6.77 l=2.74
X4 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=2.6403 pd=14.32 as=0 ps=0 w=6.77 l=2.74
X5 VDD2.t0 VN.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.6403 pd=14.32 as=2.6403 ps=14.32 w=6.77 l=2.74
X6 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=2.6403 pd=14.32 as=0 ps=0 w=6.77 l=2.74
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=2.6403 pd=14.32 as=0 ps=0 w=6.77 l=2.74
R0 B.n411 B.n410 585
R1 B.n412 B.n87 585
R2 B.n414 B.n413 585
R3 B.n416 B.n86 585
R4 B.n419 B.n418 585
R5 B.n420 B.n85 585
R6 B.n422 B.n421 585
R7 B.n424 B.n84 585
R8 B.n427 B.n426 585
R9 B.n428 B.n83 585
R10 B.n430 B.n429 585
R11 B.n432 B.n82 585
R12 B.n435 B.n434 585
R13 B.n436 B.n81 585
R14 B.n438 B.n437 585
R15 B.n440 B.n80 585
R16 B.n443 B.n442 585
R17 B.n444 B.n79 585
R18 B.n446 B.n445 585
R19 B.n448 B.n78 585
R20 B.n451 B.n450 585
R21 B.n452 B.n77 585
R22 B.n454 B.n453 585
R23 B.n456 B.n76 585
R24 B.n458 B.n457 585
R25 B.n460 B.n459 585
R26 B.n463 B.n462 585
R27 B.n464 B.n71 585
R28 B.n466 B.n465 585
R29 B.n468 B.n70 585
R30 B.n471 B.n470 585
R31 B.n472 B.n69 585
R32 B.n474 B.n473 585
R33 B.n476 B.n68 585
R34 B.n478 B.n477 585
R35 B.n480 B.n479 585
R36 B.n483 B.n482 585
R37 B.n484 B.n63 585
R38 B.n486 B.n485 585
R39 B.n488 B.n62 585
R40 B.n491 B.n490 585
R41 B.n492 B.n61 585
R42 B.n494 B.n493 585
R43 B.n496 B.n60 585
R44 B.n499 B.n498 585
R45 B.n500 B.n59 585
R46 B.n502 B.n501 585
R47 B.n504 B.n58 585
R48 B.n507 B.n506 585
R49 B.n508 B.n57 585
R50 B.n510 B.n509 585
R51 B.n512 B.n56 585
R52 B.n515 B.n514 585
R53 B.n516 B.n55 585
R54 B.n518 B.n517 585
R55 B.n520 B.n54 585
R56 B.n523 B.n522 585
R57 B.n524 B.n53 585
R58 B.n526 B.n525 585
R59 B.n528 B.n52 585
R60 B.n531 B.n530 585
R61 B.n532 B.n51 585
R62 B.n408 B.n49 585
R63 B.n535 B.n49 585
R64 B.n407 B.n48 585
R65 B.n536 B.n48 585
R66 B.n406 B.n47 585
R67 B.n537 B.n47 585
R68 B.n405 B.n404 585
R69 B.n404 B.n43 585
R70 B.n403 B.n42 585
R71 B.n543 B.n42 585
R72 B.n402 B.n41 585
R73 B.n544 B.n41 585
R74 B.n401 B.n40 585
R75 B.n545 B.n40 585
R76 B.n400 B.n399 585
R77 B.n399 B.n39 585
R78 B.n398 B.n35 585
R79 B.n551 B.n35 585
R80 B.n397 B.n34 585
R81 B.n552 B.n34 585
R82 B.n396 B.n33 585
R83 B.n553 B.n33 585
R84 B.n395 B.n394 585
R85 B.n394 B.n29 585
R86 B.n393 B.n28 585
R87 B.n559 B.n28 585
R88 B.n392 B.n27 585
R89 B.n560 B.n27 585
R90 B.n391 B.n26 585
R91 B.n561 B.n26 585
R92 B.n390 B.n389 585
R93 B.n389 B.n22 585
R94 B.n388 B.n21 585
R95 B.n567 B.n21 585
R96 B.n387 B.n20 585
R97 B.n568 B.n20 585
R98 B.n386 B.n19 585
R99 B.n569 B.n19 585
R100 B.n385 B.n384 585
R101 B.n384 B.n18 585
R102 B.n383 B.n14 585
R103 B.n575 B.n14 585
R104 B.n382 B.n13 585
R105 B.n576 B.n13 585
R106 B.n381 B.n12 585
R107 B.n577 B.n12 585
R108 B.n380 B.n379 585
R109 B.n379 B.n8 585
R110 B.n378 B.n7 585
R111 B.n583 B.n7 585
R112 B.n377 B.n6 585
R113 B.n584 B.n6 585
R114 B.n376 B.n5 585
R115 B.n585 B.n5 585
R116 B.n375 B.n374 585
R117 B.n374 B.n4 585
R118 B.n373 B.n88 585
R119 B.n373 B.n372 585
R120 B.n363 B.n89 585
R121 B.n90 B.n89 585
R122 B.n365 B.n364 585
R123 B.n366 B.n365 585
R124 B.n362 B.n95 585
R125 B.n95 B.n94 585
R126 B.n361 B.n360 585
R127 B.n360 B.n359 585
R128 B.n97 B.n96 585
R129 B.n352 B.n97 585
R130 B.n351 B.n350 585
R131 B.n353 B.n351 585
R132 B.n349 B.n102 585
R133 B.n102 B.n101 585
R134 B.n348 B.n347 585
R135 B.n347 B.n346 585
R136 B.n104 B.n103 585
R137 B.n105 B.n104 585
R138 B.n339 B.n338 585
R139 B.n340 B.n339 585
R140 B.n337 B.n110 585
R141 B.n110 B.n109 585
R142 B.n336 B.n335 585
R143 B.n335 B.n334 585
R144 B.n112 B.n111 585
R145 B.n113 B.n112 585
R146 B.n327 B.n326 585
R147 B.n328 B.n327 585
R148 B.n325 B.n118 585
R149 B.n118 B.n117 585
R150 B.n324 B.n323 585
R151 B.n323 B.n322 585
R152 B.n120 B.n119 585
R153 B.n315 B.n120 585
R154 B.n314 B.n313 585
R155 B.n316 B.n314 585
R156 B.n312 B.n125 585
R157 B.n125 B.n124 585
R158 B.n311 B.n310 585
R159 B.n310 B.n309 585
R160 B.n127 B.n126 585
R161 B.n128 B.n127 585
R162 B.n302 B.n301 585
R163 B.n303 B.n302 585
R164 B.n300 B.n133 585
R165 B.n133 B.n132 585
R166 B.n299 B.n298 585
R167 B.n298 B.n297 585
R168 B.n294 B.n137 585
R169 B.n293 B.n292 585
R170 B.n290 B.n138 585
R171 B.n290 B.n136 585
R172 B.n289 B.n288 585
R173 B.n287 B.n286 585
R174 B.n285 B.n140 585
R175 B.n283 B.n282 585
R176 B.n281 B.n141 585
R177 B.n280 B.n279 585
R178 B.n277 B.n142 585
R179 B.n275 B.n274 585
R180 B.n273 B.n143 585
R181 B.n272 B.n271 585
R182 B.n269 B.n144 585
R183 B.n267 B.n266 585
R184 B.n265 B.n145 585
R185 B.n264 B.n263 585
R186 B.n261 B.n146 585
R187 B.n259 B.n258 585
R188 B.n257 B.n147 585
R189 B.n256 B.n255 585
R190 B.n253 B.n148 585
R191 B.n251 B.n250 585
R192 B.n249 B.n149 585
R193 B.n248 B.n247 585
R194 B.n245 B.n150 585
R195 B.n243 B.n242 585
R196 B.n241 B.n151 585
R197 B.n240 B.n239 585
R198 B.n237 B.n155 585
R199 B.n235 B.n234 585
R200 B.n233 B.n156 585
R201 B.n232 B.n231 585
R202 B.n229 B.n157 585
R203 B.n227 B.n226 585
R204 B.n225 B.n158 585
R205 B.n223 B.n222 585
R206 B.n220 B.n161 585
R207 B.n218 B.n217 585
R208 B.n216 B.n162 585
R209 B.n215 B.n214 585
R210 B.n212 B.n163 585
R211 B.n210 B.n209 585
R212 B.n208 B.n164 585
R213 B.n207 B.n206 585
R214 B.n204 B.n165 585
R215 B.n202 B.n201 585
R216 B.n200 B.n166 585
R217 B.n199 B.n198 585
R218 B.n196 B.n167 585
R219 B.n194 B.n193 585
R220 B.n192 B.n168 585
R221 B.n191 B.n190 585
R222 B.n188 B.n169 585
R223 B.n186 B.n185 585
R224 B.n184 B.n170 585
R225 B.n183 B.n182 585
R226 B.n180 B.n171 585
R227 B.n178 B.n177 585
R228 B.n176 B.n172 585
R229 B.n175 B.n174 585
R230 B.n135 B.n134 585
R231 B.n136 B.n135 585
R232 B.n296 B.n295 585
R233 B.n297 B.n296 585
R234 B.n131 B.n130 585
R235 B.n132 B.n131 585
R236 B.n305 B.n304 585
R237 B.n304 B.n303 585
R238 B.n306 B.n129 585
R239 B.n129 B.n128 585
R240 B.n308 B.n307 585
R241 B.n309 B.n308 585
R242 B.n123 B.n122 585
R243 B.n124 B.n123 585
R244 B.n318 B.n317 585
R245 B.n317 B.n316 585
R246 B.n319 B.n121 585
R247 B.n315 B.n121 585
R248 B.n321 B.n320 585
R249 B.n322 B.n321 585
R250 B.n116 B.n115 585
R251 B.n117 B.n116 585
R252 B.n330 B.n329 585
R253 B.n329 B.n328 585
R254 B.n331 B.n114 585
R255 B.n114 B.n113 585
R256 B.n333 B.n332 585
R257 B.n334 B.n333 585
R258 B.n108 B.n107 585
R259 B.n109 B.n108 585
R260 B.n342 B.n341 585
R261 B.n341 B.n340 585
R262 B.n343 B.n106 585
R263 B.n106 B.n105 585
R264 B.n345 B.n344 585
R265 B.n346 B.n345 585
R266 B.n100 B.n99 585
R267 B.n101 B.n100 585
R268 B.n355 B.n354 585
R269 B.n354 B.n353 585
R270 B.n356 B.n98 585
R271 B.n352 B.n98 585
R272 B.n358 B.n357 585
R273 B.n359 B.n358 585
R274 B.n93 B.n92 585
R275 B.n94 B.n93 585
R276 B.n368 B.n367 585
R277 B.n367 B.n366 585
R278 B.n369 B.n91 585
R279 B.n91 B.n90 585
R280 B.n371 B.n370 585
R281 B.n372 B.n371 585
R282 B.n2 B.n0 585
R283 B.n4 B.n2 585
R284 B.n3 B.n1 585
R285 B.n584 B.n3 585
R286 B.n582 B.n581 585
R287 B.n583 B.n582 585
R288 B.n580 B.n9 585
R289 B.n9 B.n8 585
R290 B.n579 B.n578 585
R291 B.n578 B.n577 585
R292 B.n11 B.n10 585
R293 B.n576 B.n11 585
R294 B.n574 B.n573 585
R295 B.n575 B.n574 585
R296 B.n572 B.n15 585
R297 B.n18 B.n15 585
R298 B.n571 B.n570 585
R299 B.n570 B.n569 585
R300 B.n17 B.n16 585
R301 B.n568 B.n17 585
R302 B.n566 B.n565 585
R303 B.n567 B.n566 585
R304 B.n564 B.n23 585
R305 B.n23 B.n22 585
R306 B.n563 B.n562 585
R307 B.n562 B.n561 585
R308 B.n25 B.n24 585
R309 B.n560 B.n25 585
R310 B.n558 B.n557 585
R311 B.n559 B.n558 585
R312 B.n556 B.n30 585
R313 B.n30 B.n29 585
R314 B.n555 B.n554 585
R315 B.n554 B.n553 585
R316 B.n32 B.n31 585
R317 B.n552 B.n32 585
R318 B.n550 B.n549 585
R319 B.n551 B.n550 585
R320 B.n548 B.n36 585
R321 B.n39 B.n36 585
R322 B.n547 B.n546 585
R323 B.n546 B.n545 585
R324 B.n38 B.n37 585
R325 B.n544 B.n38 585
R326 B.n542 B.n541 585
R327 B.n543 B.n542 585
R328 B.n540 B.n44 585
R329 B.n44 B.n43 585
R330 B.n539 B.n538 585
R331 B.n538 B.n537 585
R332 B.n46 B.n45 585
R333 B.n536 B.n46 585
R334 B.n534 B.n533 585
R335 B.n535 B.n534 585
R336 B.n587 B.n586 585
R337 B.n586 B.n585 585
R338 B.n296 B.n137 530.939
R339 B.n534 B.n51 530.939
R340 B.n298 B.n135 530.939
R341 B.n410 B.n49 530.939
R342 B.n159 B.t13 267.796
R343 B.n152 B.t2 267.796
R344 B.n64 B.t6 267.796
R345 B.n72 B.t10 267.796
R346 B.n409 B.n50 256.663
R347 B.n415 B.n50 256.663
R348 B.n417 B.n50 256.663
R349 B.n423 B.n50 256.663
R350 B.n425 B.n50 256.663
R351 B.n431 B.n50 256.663
R352 B.n433 B.n50 256.663
R353 B.n439 B.n50 256.663
R354 B.n441 B.n50 256.663
R355 B.n447 B.n50 256.663
R356 B.n449 B.n50 256.663
R357 B.n455 B.n50 256.663
R358 B.n75 B.n50 256.663
R359 B.n461 B.n50 256.663
R360 B.n467 B.n50 256.663
R361 B.n469 B.n50 256.663
R362 B.n475 B.n50 256.663
R363 B.n67 B.n50 256.663
R364 B.n481 B.n50 256.663
R365 B.n487 B.n50 256.663
R366 B.n489 B.n50 256.663
R367 B.n495 B.n50 256.663
R368 B.n497 B.n50 256.663
R369 B.n503 B.n50 256.663
R370 B.n505 B.n50 256.663
R371 B.n511 B.n50 256.663
R372 B.n513 B.n50 256.663
R373 B.n519 B.n50 256.663
R374 B.n521 B.n50 256.663
R375 B.n527 B.n50 256.663
R376 B.n529 B.n50 256.663
R377 B.n291 B.n136 256.663
R378 B.n139 B.n136 256.663
R379 B.n284 B.n136 256.663
R380 B.n278 B.n136 256.663
R381 B.n276 B.n136 256.663
R382 B.n270 B.n136 256.663
R383 B.n268 B.n136 256.663
R384 B.n262 B.n136 256.663
R385 B.n260 B.n136 256.663
R386 B.n254 B.n136 256.663
R387 B.n252 B.n136 256.663
R388 B.n246 B.n136 256.663
R389 B.n244 B.n136 256.663
R390 B.n238 B.n136 256.663
R391 B.n236 B.n136 256.663
R392 B.n230 B.n136 256.663
R393 B.n228 B.n136 256.663
R394 B.n221 B.n136 256.663
R395 B.n219 B.n136 256.663
R396 B.n213 B.n136 256.663
R397 B.n211 B.n136 256.663
R398 B.n205 B.n136 256.663
R399 B.n203 B.n136 256.663
R400 B.n197 B.n136 256.663
R401 B.n195 B.n136 256.663
R402 B.n189 B.n136 256.663
R403 B.n187 B.n136 256.663
R404 B.n181 B.n136 256.663
R405 B.n179 B.n136 256.663
R406 B.n173 B.n136 256.663
R407 B.n159 B.t15 251.95
R408 B.n72 B.t11 251.95
R409 B.n152 B.t5 251.95
R410 B.n64 B.t8 251.95
R411 B.n160 B.t14 192.411
R412 B.n73 B.t12 192.411
R413 B.n153 B.t4 192.411
R414 B.n65 B.t9 192.411
R415 B.n296 B.n131 163.367
R416 B.n304 B.n131 163.367
R417 B.n304 B.n129 163.367
R418 B.n308 B.n129 163.367
R419 B.n308 B.n123 163.367
R420 B.n317 B.n123 163.367
R421 B.n317 B.n121 163.367
R422 B.n321 B.n121 163.367
R423 B.n321 B.n116 163.367
R424 B.n329 B.n116 163.367
R425 B.n329 B.n114 163.367
R426 B.n333 B.n114 163.367
R427 B.n333 B.n108 163.367
R428 B.n341 B.n108 163.367
R429 B.n341 B.n106 163.367
R430 B.n345 B.n106 163.367
R431 B.n345 B.n100 163.367
R432 B.n354 B.n100 163.367
R433 B.n354 B.n98 163.367
R434 B.n358 B.n98 163.367
R435 B.n358 B.n93 163.367
R436 B.n367 B.n93 163.367
R437 B.n367 B.n91 163.367
R438 B.n371 B.n91 163.367
R439 B.n371 B.n2 163.367
R440 B.n586 B.n2 163.367
R441 B.n586 B.n3 163.367
R442 B.n582 B.n3 163.367
R443 B.n582 B.n9 163.367
R444 B.n578 B.n9 163.367
R445 B.n578 B.n11 163.367
R446 B.n574 B.n11 163.367
R447 B.n574 B.n15 163.367
R448 B.n570 B.n15 163.367
R449 B.n570 B.n17 163.367
R450 B.n566 B.n17 163.367
R451 B.n566 B.n23 163.367
R452 B.n562 B.n23 163.367
R453 B.n562 B.n25 163.367
R454 B.n558 B.n25 163.367
R455 B.n558 B.n30 163.367
R456 B.n554 B.n30 163.367
R457 B.n554 B.n32 163.367
R458 B.n550 B.n32 163.367
R459 B.n550 B.n36 163.367
R460 B.n546 B.n36 163.367
R461 B.n546 B.n38 163.367
R462 B.n542 B.n38 163.367
R463 B.n542 B.n44 163.367
R464 B.n538 B.n44 163.367
R465 B.n538 B.n46 163.367
R466 B.n534 B.n46 163.367
R467 B.n292 B.n290 163.367
R468 B.n290 B.n289 163.367
R469 B.n286 B.n285 163.367
R470 B.n283 B.n141 163.367
R471 B.n279 B.n277 163.367
R472 B.n275 B.n143 163.367
R473 B.n271 B.n269 163.367
R474 B.n267 B.n145 163.367
R475 B.n263 B.n261 163.367
R476 B.n259 B.n147 163.367
R477 B.n255 B.n253 163.367
R478 B.n251 B.n149 163.367
R479 B.n247 B.n245 163.367
R480 B.n243 B.n151 163.367
R481 B.n239 B.n237 163.367
R482 B.n235 B.n156 163.367
R483 B.n231 B.n229 163.367
R484 B.n227 B.n158 163.367
R485 B.n222 B.n220 163.367
R486 B.n218 B.n162 163.367
R487 B.n214 B.n212 163.367
R488 B.n210 B.n164 163.367
R489 B.n206 B.n204 163.367
R490 B.n202 B.n166 163.367
R491 B.n198 B.n196 163.367
R492 B.n194 B.n168 163.367
R493 B.n190 B.n188 163.367
R494 B.n186 B.n170 163.367
R495 B.n182 B.n180 163.367
R496 B.n178 B.n172 163.367
R497 B.n174 B.n135 163.367
R498 B.n298 B.n133 163.367
R499 B.n302 B.n133 163.367
R500 B.n302 B.n127 163.367
R501 B.n310 B.n127 163.367
R502 B.n310 B.n125 163.367
R503 B.n314 B.n125 163.367
R504 B.n314 B.n120 163.367
R505 B.n323 B.n120 163.367
R506 B.n323 B.n118 163.367
R507 B.n327 B.n118 163.367
R508 B.n327 B.n112 163.367
R509 B.n335 B.n112 163.367
R510 B.n335 B.n110 163.367
R511 B.n339 B.n110 163.367
R512 B.n339 B.n104 163.367
R513 B.n347 B.n104 163.367
R514 B.n347 B.n102 163.367
R515 B.n351 B.n102 163.367
R516 B.n351 B.n97 163.367
R517 B.n360 B.n97 163.367
R518 B.n360 B.n95 163.367
R519 B.n365 B.n95 163.367
R520 B.n365 B.n89 163.367
R521 B.n373 B.n89 163.367
R522 B.n374 B.n373 163.367
R523 B.n374 B.n5 163.367
R524 B.n6 B.n5 163.367
R525 B.n7 B.n6 163.367
R526 B.n379 B.n7 163.367
R527 B.n379 B.n12 163.367
R528 B.n13 B.n12 163.367
R529 B.n14 B.n13 163.367
R530 B.n384 B.n14 163.367
R531 B.n384 B.n19 163.367
R532 B.n20 B.n19 163.367
R533 B.n21 B.n20 163.367
R534 B.n389 B.n21 163.367
R535 B.n389 B.n26 163.367
R536 B.n27 B.n26 163.367
R537 B.n28 B.n27 163.367
R538 B.n394 B.n28 163.367
R539 B.n394 B.n33 163.367
R540 B.n34 B.n33 163.367
R541 B.n35 B.n34 163.367
R542 B.n399 B.n35 163.367
R543 B.n399 B.n40 163.367
R544 B.n41 B.n40 163.367
R545 B.n42 B.n41 163.367
R546 B.n404 B.n42 163.367
R547 B.n404 B.n47 163.367
R548 B.n48 B.n47 163.367
R549 B.n49 B.n48 163.367
R550 B.n530 B.n528 163.367
R551 B.n526 B.n53 163.367
R552 B.n522 B.n520 163.367
R553 B.n518 B.n55 163.367
R554 B.n514 B.n512 163.367
R555 B.n510 B.n57 163.367
R556 B.n506 B.n504 163.367
R557 B.n502 B.n59 163.367
R558 B.n498 B.n496 163.367
R559 B.n494 B.n61 163.367
R560 B.n490 B.n488 163.367
R561 B.n486 B.n63 163.367
R562 B.n482 B.n480 163.367
R563 B.n477 B.n476 163.367
R564 B.n474 B.n69 163.367
R565 B.n470 B.n468 163.367
R566 B.n466 B.n71 163.367
R567 B.n462 B.n460 163.367
R568 B.n457 B.n456 163.367
R569 B.n454 B.n77 163.367
R570 B.n450 B.n448 163.367
R571 B.n446 B.n79 163.367
R572 B.n442 B.n440 163.367
R573 B.n438 B.n81 163.367
R574 B.n434 B.n432 163.367
R575 B.n430 B.n83 163.367
R576 B.n426 B.n424 163.367
R577 B.n422 B.n85 163.367
R578 B.n418 B.n416 163.367
R579 B.n414 B.n87 163.367
R580 B.n297 B.n136 123.288
R581 B.n535 B.n50 123.288
R582 B.n291 B.n137 71.676
R583 B.n289 B.n139 71.676
R584 B.n285 B.n284 71.676
R585 B.n278 B.n141 71.676
R586 B.n277 B.n276 71.676
R587 B.n270 B.n143 71.676
R588 B.n269 B.n268 71.676
R589 B.n262 B.n145 71.676
R590 B.n261 B.n260 71.676
R591 B.n254 B.n147 71.676
R592 B.n253 B.n252 71.676
R593 B.n246 B.n149 71.676
R594 B.n245 B.n244 71.676
R595 B.n238 B.n151 71.676
R596 B.n237 B.n236 71.676
R597 B.n230 B.n156 71.676
R598 B.n229 B.n228 71.676
R599 B.n221 B.n158 71.676
R600 B.n220 B.n219 71.676
R601 B.n213 B.n162 71.676
R602 B.n212 B.n211 71.676
R603 B.n205 B.n164 71.676
R604 B.n204 B.n203 71.676
R605 B.n197 B.n166 71.676
R606 B.n196 B.n195 71.676
R607 B.n189 B.n168 71.676
R608 B.n188 B.n187 71.676
R609 B.n181 B.n170 71.676
R610 B.n180 B.n179 71.676
R611 B.n173 B.n172 71.676
R612 B.n529 B.n51 71.676
R613 B.n528 B.n527 71.676
R614 B.n521 B.n53 71.676
R615 B.n520 B.n519 71.676
R616 B.n513 B.n55 71.676
R617 B.n512 B.n511 71.676
R618 B.n505 B.n57 71.676
R619 B.n504 B.n503 71.676
R620 B.n497 B.n59 71.676
R621 B.n496 B.n495 71.676
R622 B.n489 B.n61 71.676
R623 B.n488 B.n487 71.676
R624 B.n481 B.n63 71.676
R625 B.n480 B.n67 71.676
R626 B.n476 B.n475 71.676
R627 B.n469 B.n69 71.676
R628 B.n468 B.n467 71.676
R629 B.n461 B.n71 71.676
R630 B.n460 B.n75 71.676
R631 B.n456 B.n455 71.676
R632 B.n449 B.n77 71.676
R633 B.n448 B.n447 71.676
R634 B.n441 B.n79 71.676
R635 B.n440 B.n439 71.676
R636 B.n433 B.n81 71.676
R637 B.n432 B.n431 71.676
R638 B.n425 B.n83 71.676
R639 B.n424 B.n423 71.676
R640 B.n417 B.n85 71.676
R641 B.n416 B.n415 71.676
R642 B.n409 B.n87 71.676
R643 B.n410 B.n409 71.676
R644 B.n415 B.n414 71.676
R645 B.n418 B.n417 71.676
R646 B.n423 B.n422 71.676
R647 B.n426 B.n425 71.676
R648 B.n431 B.n430 71.676
R649 B.n434 B.n433 71.676
R650 B.n439 B.n438 71.676
R651 B.n442 B.n441 71.676
R652 B.n447 B.n446 71.676
R653 B.n450 B.n449 71.676
R654 B.n455 B.n454 71.676
R655 B.n457 B.n75 71.676
R656 B.n462 B.n461 71.676
R657 B.n467 B.n466 71.676
R658 B.n470 B.n469 71.676
R659 B.n475 B.n474 71.676
R660 B.n477 B.n67 71.676
R661 B.n482 B.n481 71.676
R662 B.n487 B.n486 71.676
R663 B.n490 B.n489 71.676
R664 B.n495 B.n494 71.676
R665 B.n498 B.n497 71.676
R666 B.n503 B.n502 71.676
R667 B.n506 B.n505 71.676
R668 B.n511 B.n510 71.676
R669 B.n514 B.n513 71.676
R670 B.n519 B.n518 71.676
R671 B.n522 B.n521 71.676
R672 B.n527 B.n526 71.676
R673 B.n530 B.n529 71.676
R674 B.n292 B.n291 71.676
R675 B.n286 B.n139 71.676
R676 B.n284 B.n283 71.676
R677 B.n279 B.n278 71.676
R678 B.n276 B.n275 71.676
R679 B.n271 B.n270 71.676
R680 B.n268 B.n267 71.676
R681 B.n263 B.n262 71.676
R682 B.n260 B.n259 71.676
R683 B.n255 B.n254 71.676
R684 B.n252 B.n251 71.676
R685 B.n247 B.n246 71.676
R686 B.n244 B.n243 71.676
R687 B.n239 B.n238 71.676
R688 B.n236 B.n235 71.676
R689 B.n231 B.n230 71.676
R690 B.n228 B.n227 71.676
R691 B.n222 B.n221 71.676
R692 B.n219 B.n218 71.676
R693 B.n214 B.n213 71.676
R694 B.n211 B.n210 71.676
R695 B.n206 B.n205 71.676
R696 B.n203 B.n202 71.676
R697 B.n198 B.n197 71.676
R698 B.n195 B.n194 71.676
R699 B.n190 B.n189 71.676
R700 B.n187 B.n186 71.676
R701 B.n182 B.n181 71.676
R702 B.n179 B.n178 71.676
R703 B.n174 B.n173 71.676
R704 B.n297 B.n132 62.101
R705 B.n303 B.n132 62.101
R706 B.n303 B.n128 62.101
R707 B.n309 B.n128 62.101
R708 B.n309 B.n124 62.101
R709 B.n316 B.n124 62.101
R710 B.n316 B.n315 62.101
R711 B.n322 B.n117 62.101
R712 B.n328 B.n117 62.101
R713 B.n328 B.n113 62.101
R714 B.n334 B.n113 62.101
R715 B.n334 B.n109 62.101
R716 B.n340 B.n109 62.101
R717 B.n340 B.n105 62.101
R718 B.n346 B.n105 62.101
R719 B.n346 B.n101 62.101
R720 B.n353 B.n101 62.101
R721 B.n353 B.n352 62.101
R722 B.n359 B.n94 62.101
R723 B.n366 B.n94 62.101
R724 B.n366 B.n90 62.101
R725 B.n372 B.n90 62.101
R726 B.n372 B.n4 62.101
R727 B.n585 B.n4 62.101
R728 B.n585 B.n584 62.101
R729 B.n584 B.n583 62.101
R730 B.n583 B.n8 62.101
R731 B.n577 B.n8 62.101
R732 B.n577 B.n576 62.101
R733 B.n576 B.n575 62.101
R734 B.n569 B.n18 62.101
R735 B.n569 B.n568 62.101
R736 B.n568 B.n567 62.101
R737 B.n567 B.n22 62.101
R738 B.n561 B.n22 62.101
R739 B.n561 B.n560 62.101
R740 B.n560 B.n559 62.101
R741 B.n559 B.n29 62.101
R742 B.n553 B.n29 62.101
R743 B.n553 B.n552 62.101
R744 B.n552 B.n551 62.101
R745 B.n545 B.n39 62.101
R746 B.n545 B.n544 62.101
R747 B.n544 B.n543 62.101
R748 B.n543 B.n43 62.101
R749 B.n537 B.n43 62.101
R750 B.n537 B.n536 62.101
R751 B.n536 B.n535 62.101
R752 B.n224 B.n160 59.5399
R753 B.n160 B.n159 59.5399
R754 B.n154 B.n153 59.5399
R755 B.n153 B.n152 59.5399
R756 B.n65 B.n64 59.5399
R757 B.n66 B.n65 59.5399
R758 B.n73 B.n72 59.5399
R759 B.n74 B.n73 59.5399
R760 B.n352 B.t0 54.795
R761 B.n18 B.t1 54.795
R762 B.n315 B.t3 40.1831
R763 B.n39 B.t7 40.1831
R764 B.n533 B.n532 34.4981
R765 B.n411 B.n408 34.4981
R766 B.n299 B.n134 34.4981
R767 B.n295 B.n294 34.4981
R768 B.n322 B.t3 21.9183
R769 B.n551 B.t7 21.9183
R770 B B.n587 18.0485
R771 B.n532 B.n531 10.6151
R772 B.n531 B.n52 10.6151
R773 B.n525 B.n52 10.6151
R774 B.n525 B.n524 10.6151
R775 B.n524 B.n523 10.6151
R776 B.n523 B.n54 10.6151
R777 B.n517 B.n54 10.6151
R778 B.n517 B.n516 10.6151
R779 B.n516 B.n515 10.6151
R780 B.n515 B.n56 10.6151
R781 B.n509 B.n56 10.6151
R782 B.n509 B.n508 10.6151
R783 B.n508 B.n507 10.6151
R784 B.n507 B.n58 10.6151
R785 B.n501 B.n58 10.6151
R786 B.n501 B.n500 10.6151
R787 B.n500 B.n499 10.6151
R788 B.n499 B.n60 10.6151
R789 B.n493 B.n60 10.6151
R790 B.n493 B.n492 10.6151
R791 B.n492 B.n491 10.6151
R792 B.n491 B.n62 10.6151
R793 B.n485 B.n62 10.6151
R794 B.n485 B.n484 10.6151
R795 B.n484 B.n483 10.6151
R796 B.n479 B.n478 10.6151
R797 B.n478 B.n68 10.6151
R798 B.n473 B.n68 10.6151
R799 B.n473 B.n472 10.6151
R800 B.n472 B.n471 10.6151
R801 B.n471 B.n70 10.6151
R802 B.n465 B.n70 10.6151
R803 B.n465 B.n464 10.6151
R804 B.n464 B.n463 10.6151
R805 B.n459 B.n458 10.6151
R806 B.n458 B.n76 10.6151
R807 B.n453 B.n76 10.6151
R808 B.n453 B.n452 10.6151
R809 B.n452 B.n451 10.6151
R810 B.n451 B.n78 10.6151
R811 B.n445 B.n78 10.6151
R812 B.n445 B.n444 10.6151
R813 B.n444 B.n443 10.6151
R814 B.n443 B.n80 10.6151
R815 B.n437 B.n80 10.6151
R816 B.n437 B.n436 10.6151
R817 B.n436 B.n435 10.6151
R818 B.n435 B.n82 10.6151
R819 B.n429 B.n82 10.6151
R820 B.n429 B.n428 10.6151
R821 B.n428 B.n427 10.6151
R822 B.n427 B.n84 10.6151
R823 B.n421 B.n84 10.6151
R824 B.n421 B.n420 10.6151
R825 B.n420 B.n419 10.6151
R826 B.n419 B.n86 10.6151
R827 B.n413 B.n86 10.6151
R828 B.n413 B.n412 10.6151
R829 B.n412 B.n411 10.6151
R830 B.n300 B.n299 10.6151
R831 B.n301 B.n300 10.6151
R832 B.n301 B.n126 10.6151
R833 B.n311 B.n126 10.6151
R834 B.n312 B.n311 10.6151
R835 B.n313 B.n312 10.6151
R836 B.n313 B.n119 10.6151
R837 B.n324 B.n119 10.6151
R838 B.n325 B.n324 10.6151
R839 B.n326 B.n325 10.6151
R840 B.n326 B.n111 10.6151
R841 B.n336 B.n111 10.6151
R842 B.n337 B.n336 10.6151
R843 B.n338 B.n337 10.6151
R844 B.n338 B.n103 10.6151
R845 B.n348 B.n103 10.6151
R846 B.n349 B.n348 10.6151
R847 B.n350 B.n349 10.6151
R848 B.n350 B.n96 10.6151
R849 B.n361 B.n96 10.6151
R850 B.n362 B.n361 10.6151
R851 B.n364 B.n362 10.6151
R852 B.n364 B.n363 10.6151
R853 B.n363 B.n88 10.6151
R854 B.n375 B.n88 10.6151
R855 B.n376 B.n375 10.6151
R856 B.n377 B.n376 10.6151
R857 B.n378 B.n377 10.6151
R858 B.n380 B.n378 10.6151
R859 B.n381 B.n380 10.6151
R860 B.n382 B.n381 10.6151
R861 B.n383 B.n382 10.6151
R862 B.n385 B.n383 10.6151
R863 B.n386 B.n385 10.6151
R864 B.n387 B.n386 10.6151
R865 B.n388 B.n387 10.6151
R866 B.n390 B.n388 10.6151
R867 B.n391 B.n390 10.6151
R868 B.n392 B.n391 10.6151
R869 B.n393 B.n392 10.6151
R870 B.n395 B.n393 10.6151
R871 B.n396 B.n395 10.6151
R872 B.n397 B.n396 10.6151
R873 B.n398 B.n397 10.6151
R874 B.n400 B.n398 10.6151
R875 B.n401 B.n400 10.6151
R876 B.n402 B.n401 10.6151
R877 B.n403 B.n402 10.6151
R878 B.n405 B.n403 10.6151
R879 B.n406 B.n405 10.6151
R880 B.n407 B.n406 10.6151
R881 B.n408 B.n407 10.6151
R882 B.n294 B.n293 10.6151
R883 B.n293 B.n138 10.6151
R884 B.n288 B.n138 10.6151
R885 B.n288 B.n287 10.6151
R886 B.n287 B.n140 10.6151
R887 B.n282 B.n140 10.6151
R888 B.n282 B.n281 10.6151
R889 B.n281 B.n280 10.6151
R890 B.n280 B.n142 10.6151
R891 B.n274 B.n142 10.6151
R892 B.n274 B.n273 10.6151
R893 B.n273 B.n272 10.6151
R894 B.n272 B.n144 10.6151
R895 B.n266 B.n144 10.6151
R896 B.n266 B.n265 10.6151
R897 B.n265 B.n264 10.6151
R898 B.n264 B.n146 10.6151
R899 B.n258 B.n146 10.6151
R900 B.n258 B.n257 10.6151
R901 B.n257 B.n256 10.6151
R902 B.n256 B.n148 10.6151
R903 B.n250 B.n148 10.6151
R904 B.n250 B.n249 10.6151
R905 B.n249 B.n248 10.6151
R906 B.n248 B.n150 10.6151
R907 B.n242 B.n241 10.6151
R908 B.n241 B.n240 10.6151
R909 B.n240 B.n155 10.6151
R910 B.n234 B.n155 10.6151
R911 B.n234 B.n233 10.6151
R912 B.n233 B.n232 10.6151
R913 B.n232 B.n157 10.6151
R914 B.n226 B.n157 10.6151
R915 B.n226 B.n225 10.6151
R916 B.n223 B.n161 10.6151
R917 B.n217 B.n161 10.6151
R918 B.n217 B.n216 10.6151
R919 B.n216 B.n215 10.6151
R920 B.n215 B.n163 10.6151
R921 B.n209 B.n163 10.6151
R922 B.n209 B.n208 10.6151
R923 B.n208 B.n207 10.6151
R924 B.n207 B.n165 10.6151
R925 B.n201 B.n165 10.6151
R926 B.n201 B.n200 10.6151
R927 B.n200 B.n199 10.6151
R928 B.n199 B.n167 10.6151
R929 B.n193 B.n167 10.6151
R930 B.n193 B.n192 10.6151
R931 B.n192 B.n191 10.6151
R932 B.n191 B.n169 10.6151
R933 B.n185 B.n169 10.6151
R934 B.n185 B.n184 10.6151
R935 B.n184 B.n183 10.6151
R936 B.n183 B.n171 10.6151
R937 B.n177 B.n171 10.6151
R938 B.n177 B.n176 10.6151
R939 B.n176 B.n175 10.6151
R940 B.n175 B.n134 10.6151
R941 B.n295 B.n130 10.6151
R942 B.n305 B.n130 10.6151
R943 B.n306 B.n305 10.6151
R944 B.n307 B.n306 10.6151
R945 B.n307 B.n122 10.6151
R946 B.n318 B.n122 10.6151
R947 B.n319 B.n318 10.6151
R948 B.n320 B.n319 10.6151
R949 B.n320 B.n115 10.6151
R950 B.n330 B.n115 10.6151
R951 B.n331 B.n330 10.6151
R952 B.n332 B.n331 10.6151
R953 B.n332 B.n107 10.6151
R954 B.n342 B.n107 10.6151
R955 B.n343 B.n342 10.6151
R956 B.n344 B.n343 10.6151
R957 B.n344 B.n99 10.6151
R958 B.n355 B.n99 10.6151
R959 B.n356 B.n355 10.6151
R960 B.n357 B.n356 10.6151
R961 B.n357 B.n92 10.6151
R962 B.n368 B.n92 10.6151
R963 B.n369 B.n368 10.6151
R964 B.n370 B.n369 10.6151
R965 B.n370 B.n0 10.6151
R966 B.n581 B.n1 10.6151
R967 B.n581 B.n580 10.6151
R968 B.n580 B.n579 10.6151
R969 B.n579 B.n10 10.6151
R970 B.n573 B.n10 10.6151
R971 B.n573 B.n572 10.6151
R972 B.n572 B.n571 10.6151
R973 B.n571 B.n16 10.6151
R974 B.n565 B.n16 10.6151
R975 B.n565 B.n564 10.6151
R976 B.n564 B.n563 10.6151
R977 B.n563 B.n24 10.6151
R978 B.n557 B.n24 10.6151
R979 B.n557 B.n556 10.6151
R980 B.n556 B.n555 10.6151
R981 B.n555 B.n31 10.6151
R982 B.n549 B.n31 10.6151
R983 B.n549 B.n548 10.6151
R984 B.n548 B.n547 10.6151
R985 B.n547 B.n37 10.6151
R986 B.n541 B.n37 10.6151
R987 B.n541 B.n540 10.6151
R988 B.n540 B.n539 10.6151
R989 B.n539 B.n45 10.6151
R990 B.n533 B.n45 10.6151
R991 B.n483 B.n66 9.36635
R992 B.n459 B.n74 9.36635
R993 B.n154 B.n150 9.36635
R994 B.n224 B.n223 9.36635
R995 B.n359 B.t0 7.30644
R996 B.n575 B.t1 7.30644
R997 B.n587 B.n0 2.81026
R998 B.n587 B.n1 2.81026
R999 B.n479 B.n66 1.24928
R1000 B.n463 B.n74 1.24928
R1001 B.n242 B.n154 1.24928
R1002 B.n225 B.n224 1.24928
R1003 VP.n0 VP.t1 141.708
R1004 VP.n0 VP.t0 100.642
R1005 VP VP.n0 0.431811
R1006 VTAIL.n138 VTAIL.n108 289.615
R1007 VTAIL.n30 VTAIL.n0 289.615
R1008 VTAIL.n102 VTAIL.n72 289.615
R1009 VTAIL.n66 VTAIL.n36 289.615
R1010 VTAIL.n121 VTAIL.n120 185
R1011 VTAIL.n123 VTAIL.n122 185
R1012 VTAIL.n116 VTAIL.n115 185
R1013 VTAIL.n129 VTAIL.n128 185
R1014 VTAIL.n131 VTAIL.n130 185
R1015 VTAIL.n112 VTAIL.n111 185
R1016 VTAIL.n137 VTAIL.n136 185
R1017 VTAIL.n139 VTAIL.n138 185
R1018 VTAIL.n13 VTAIL.n12 185
R1019 VTAIL.n15 VTAIL.n14 185
R1020 VTAIL.n8 VTAIL.n7 185
R1021 VTAIL.n21 VTAIL.n20 185
R1022 VTAIL.n23 VTAIL.n22 185
R1023 VTAIL.n4 VTAIL.n3 185
R1024 VTAIL.n29 VTAIL.n28 185
R1025 VTAIL.n31 VTAIL.n30 185
R1026 VTAIL.n103 VTAIL.n102 185
R1027 VTAIL.n101 VTAIL.n100 185
R1028 VTAIL.n76 VTAIL.n75 185
R1029 VTAIL.n95 VTAIL.n94 185
R1030 VTAIL.n93 VTAIL.n92 185
R1031 VTAIL.n80 VTAIL.n79 185
R1032 VTAIL.n87 VTAIL.n86 185
R1033 VTAIL.n85 VTAIL.n84 185
R1034 VTAIL.n67 VTAIL.n66 185
R1035 VTAIL.n65 VTAIL.n64 185
R1036 VTAIL.n40 VTAIL.n39 185
R1037 VTAIL.n59 VTAIL.n58 185
R1038 VTAIL.n57 VTAIL.n56 185
R1039 VTAIL.n44 VTAIL.n43 185
R1040 VTAIL.n51 VTAIL.n50 185
R1041 VTAIL.n49 VTAIL.n48 185
R1042 VTAIL.n119 VTAIL.t1 147.659
R1043 VTAIL.n11 VTAIL.t2 147.659
R1044 VTAIL.n83 VTAIL.t3 147.659
R1045 VTAIL.n47 VTAIL.t0 147.659
R1046 VTAIL.n122 VTAIL.n121 104.615
R1047 VTAIL.n122 VTAIL.n115 104.615
R1048 VTAIL.n129 VTAIL.n115 104.615
R1049 VTAIL.n130 VTAIL.n129 104.615
R1050 VTAIL.n130 VTAIL.n111 104.615
R1051 VTAIL.n137 VTAIL.n111 104.615
R1052 VTAIL.n138 VTAIL.n137 104.615
R1053 VTAIL.n14 VTAIL.n13 104.615
R1054 VTAIL.n14 VTAIL.n7 104.615
R1055 VTAIL.n21 VTAIL.n7 104.615
R1056 VTAIL.n22 VTAIL.n21 104.615
R1057 VTAIL.n22 VTAIL.n3 104.615
R1058 VTAIL.n29 VTAIL.n3 104.615
R1059 VTAIL.n30 VTAIL.n29 104.615
R1060 VTAIL.n102 VTAIL.n101 104.615
R1061 VTAIL.n101 VTAIL.n75 104.615
R1062 VTAIL.n94 VTAIL.n75 104.615
R1063 VTAIL.n94 VTAIL.n93 104.615
R1064 VTAIL.n93 VTAIL.n79 104.615
R1065 VTAIL.n86 VTAIL.n79 104.615
R1066 VTAIL.n86 VTAIL.n85 104.615
R1067 VTAIL.n66 VTAIL.n65 104.615
R1068 VTAIL.n65 VTAIL.n39 104.615
R1069 VTAIL.n58 VTAIL.n39 104.615
R1070 VTAIL.n58 VTAIL.n57 104.615
R1071 VTAIL.n57 VTAIL.n43 104.615
R1072 VTAIL.n50 VTAIL.n43 104.615
R1073 VTAIL.n50 VTAIL.n49 104.615
R1074 VTAIL.n121 VTAIL.t1 52.3082
R1075 VTAIL.n13 VTAIL.t2 52.3082
R1076 VTAIL.n85 VTAIL.t3 52.3082
R1077 VTAIL.n49 VTAIL.t0 52.3082
R1078 VTAIL.n143 VTAIL.n142 33.155
R1079 VTAIL.n35 VTAIL.n34 33.155
R1080 VTAIL.n107 VTAIL.n106 33.155
R1081 VTAIL.n71 VTAIL.n70 33.155
R1082 VTAIL.n71 VTAIL.n35 23.4962
R1083 VTAIL.n143 VTAIL.n107 20.8496
R1084 VTAIL.n120 VTAIL.n119 15.6676
R1085 VTAIL.n12 VTAIL.n11 15.6676
R1086 VTAIL.n84 VTAIL.n83 15.6676
R1087 VTAIL.n48 VTAIL.n47 15.6676
R1088 VTAIL.n123 VTAIL.n118 12.8005
R1089 VTAIL.n15 VTAIL.n10 12.8005
R1090 VTAIL.n87 VTAIL.n82 12.8005
R1091 VTAIL.n51 VTAIL.n46 12.8005
R1092 VTAIL.n124 VTAIL.n116 12.0247
R1093 VTAIL.n16 VTAIL.n8 12.0247
R1094 VTAIL.n88 VTAIL.n80 12.0247
R1095 VTAIL.n52 VTAIL.n44 12.0247
R1096 VTAIL.n128 VTAIL.n127 11.249
R1097 VTAIL.n20 VTAIL.n19 11.249
R1098 VTAIL.n92 VTAIL.n91 11.249
R1099 VTAIL.n56 VTAIL.n55 11.249
R1100 VTAIL.n131 VTAIL.n114 10.4732
R1101 VTAIL.n23 VTAIL.n6 10.4732
R1102 VTAIL.n95 VTAIL.n78 10.4732
R1103 VTAIL.n59 VTAIL.n42 10.4732
R1104 VTAIL.n132 VTAIL.n112 9.69747
R1105 VTAIL.n24 VTAIL.n4 9.69747
R1106 VTAIL.n96 VTAIL.n76 9.69747
R1107 VTAIL.n60 VTAIL.n40 9.69747
R1108 VTAIL.n142 VTAIL.n141 9.45567
R1109 VTAIL.n34 VTAIL.n33 9.45567
R1110 VTAIL.n106 VTAIL.n105 9.45567
R1111 VTAIL.n70 VTAIL.n69 9.45567
R1112 VTAIL.n110 VTAIL.n109 9.3005
R1113 VTAIL.n135 VTAIL.n134 9.3005
R1114 VTAIL.n133 VTAIL.n132 9.3005
R1115 VTAIL.n114 VTAIL.n113 9.3005
R1116 VTAIL.n127 VTAIL.n126 9.3005
R1117 VTAIL.n125 VTAIL.n124 9.3005
R1118 VTAIL.n118 VTAIL.n117 9.3005
R1119 VTAIL.n141 VTAIL.n140 9.3005
R1120 VTAIL.n2 VTAIL.n1 9.3005
R1121 VTAIL.n27 VTAIL.n26 9.3005
R1122 VTAIL.n25 VTAIL.n24 9.3005
R1123 VTAIL.n6 VTAIL.n5 9.3005
R1124 VTAIL.n19 VTAIL.n18 9.3005
R1125 VTAIL.n17 VTAIL.n16 9.3005
R1126 VTAIL.n10 VTAIL.n9 9.3005
R1127 VTAIL.n33 VTAIL.n32 9.3005
R1128 VTAIL.n105 VTAIL.n104 9.3005
R1129 VTAIL.n74 VTAIL.n73 9.3005
R1130 VTAIL.n99 VTAIL.n98 9.3005
R1131 VTAIL.n97 VTAIL.n96 9.3005
R1132 VTAIL.n78 VTAIL.n77 9.3005
R1133 VTAIL.n91 VTAIL.n90 9.3005
R1134 VTAIL.n89 VTAIL.n88 9.3005
R1135 VTAIL.n82 VTAIL.n81 9.3005
R1136 VTAIL.n69 VTAIL.n68 9.3005
R1137 VTAIL.n38 VTAIL.n37 9.3005
R1138 VTAIL.n63 VTAIL.n62 9.3005
R1139 VTAIL.n61 VTAIL.n60 9.3005
R1140 VTAIL.n42 VTAIL.n41 9.3005
R1141 VTAIL.n55 VTAIL.n54 9.3005
R1142 VTAIL.n53 VTAIL.n52 9.3005
R1143 VTAIL.n46 VTAIL.n45 9.3005
R1144 VTAIL.n136 VTAIL.n135 8.92171
R1145 VTAIL.n28 VTAIL.n27 8.92171
R1146 VTAIL.n100 VTAIL.n99 8.92171
R1147 VTAIL.n64 VTAIL.n63 8.92171
R1148 VTAIL.n139 VTAIL.n110 8.14595
R1149 VTAIL.n31 VTAIL.n2 8.14595
R1150 VTAIL.n103 VTAIL.n74 8.14595
R1151 VTAIL.n67 VTAIL.n38 8.14595
R1152 VTAIL.n140 VTAIL.n108 7.3702
R1153 VTAIL.n32 VTAIL.n0 7.3702
R1154 VTAIL.n104 VTAIL.n72 7.3702
R1155 VTAIL.n68 VTAIL.n36 7.3702
R1156 VTAIL.n142 VTAIL.n108 6.59444
R1157 VTAIL.n34 VTAIL.n0 6.59444
R1158 VTAIL.n106 VTAIL.n72 6.59444
R1159 VTAIL.n70 VTAIL.n36 6.59444
R1160 VTAIL.n140 VTAIL.n139 5.81868
R1161 VTAIL.n32 VTAIL.n31 5.81868
R1162 VTAIL.n104 VTAIL.n103 5.81868
R1163 VTAIL.n68 VTAIL.n67 5.81868
R1164 VTAIL.n136 VTAIL.n110 5.04292
R1165 VTAIL.n28 VTAIL.n2 5.04292
R1166 VTAIL.n100 VTAIL.n74 5.04292
R1167 VTAIL.n64 VTAIL.n38 5.04292
R1168 VTAIL.n119 VTAIL.n117 4.38571
R1169 VTAIL.n11 VTAIL.n9 4.38571
R1170 VTAIL.n83 VTAIL.n81 4.38571
R1171 VTAIL.n47 VTAIL.n45 4.38571
R1172 VTAIL.n135 VTAIL.n112 4.26717
R1173 VTAIL.n27 VTAIL.n4 4.26717
R1174 VTAIL.n99 VTAIL.n76 4.26717
R1175 VTAIL.n63 VTAIL.n40 4.26717
R1176 VTAIL.n132 VTAIL.n131 3.49141
R1177 VTAIL.n24 VTAIL.n23 3.49141
R1178 VTAIL.n96 VTAIL.n95 3.49141
R1179 VTAIL.n60 VTAIL.n59 3.49141
R1180 VTAIL.n128 VTAIL.n114 2.71565
R1181 VTAIL.n20 VTAIL.n6 2.71565
R1182 VTAIL.n92 VTAIL.n78 2.71565
R1183 VTAIL.n56 VTAIL.n42 2.71565
R1184 VTAIL.n127 VTAIL.n116 1.93989
R1185 VTAIL.n19 VTAIL.n8 1.93989
R1186 VTAIL.n91 VTAIL.n80 1.93989
R1187 VTAIL.n55 VTAIL.n44 1.93989
R1188 VTAIL.n107 VTAIL.n71 1.7936
R1189 VTAIL VTAIL.n35 1.19016
R1190 VTAIL.n124 VTAIL.n123 1.16414
R1191 VTAIL.n16 VTAIL.n15 1.16414
R1192 VTAIL.n88 VTAIL.n87 1.16414
R1193 VTAIL.n52 VTAIL.n51 1.16414
R1194 VTAIL VTAIL.n143 0.603948
R1195 VTAIL.n120 VTAIL.n118 0.388379
R1196 VTAIL.n12 VTAIL.n10 0.388379
R1197 VTAIL.n84 VTAIL.n82 0.388379
R1198 VTAIL.n48 VTAIL.n46 0.388379
R1199 VTAIL.n125 VTAIL.n117 0.155672
R1200 VTAIL.n126 VTAIL.n125 0.155672
R1201 VTAIL.n126 VTAIL.n113 0.155672
R1202 VTAIL.n133 VTAIL.n113 0.155672
R1203 VTAIL.n134 VTAIL.n133 0.155672
R1204 VTAIL.n134 VTAIL.n109 0.155672
R1205 VTAIL.n141 VTAIL.n109 0.155672
R1206 VTAIL.n17 VTAIL.n9 0.155672
R1207 VTAIL.n18 VTAIL.n17 0.155672
R1208 VTAIL.n18 VTAIL.n5 0.155672
R1209 VTAIL.n25 VTAIL.n5 0.155672
R1210 VTAIL.n26 VTAIL.n25 0.155672
R1211 VTAIL.n26 VTAIL.n1 0.155672
R1212 VTAIL.n33 VTAIL.n1 0.155672
R1213 VTAIL.n105 VTAIL.n73 0.155672
R1214 VTAIL.n98 VTAIL.n73 0.155672
R1215 VTAIL.n98 VTAIL.n97 0.155672
R1216 VTAIL.n97 VTAIL.n77 0.155672
R1217 VTAIL.n90 VTAIL.n77 0.155672
R1218 VTAIL.n90 VTAIL.n89 0.155672
R1219 VTAIL.n89 VTAIL.n81 0.155672
R1220 VTAIL.n69 VTAIL.n37 0.155672
R1221 VTAIL.n62 VTAIL.n37 0.155672
R1222 VTAIL.n62 VTAIL.n61 0.155672
R1223 VTAIL.n61 VTAIL.n41 0.155672
R1224 VTAIL.n54 VTAIL.n41 0.155672
R1225 VTAIL.n54 VTAIL.n53 0.155672
R1226 VTAIL.n53 VTAIL.n45 0.155672
R1227 VDD1.n30 VDD1.n0 289.615
R1228 VDD1.n65 VDD1.n35 289.615
R1229 VDD1.n31 VDD1.n30 185
R1230 VDD1.n29 VDD1.n28 185
R1231 VDD1.n4 VDD1.n3 185
R1232 VDD1.n23 VDD1.n22 185
R1233 VDD1.n21 VDD1.n20 185
R1234 VDD1.n8 VDD1.n7 185
R1235 VDD1.n15 VDD1.n14 185
R1236 VDD1.n13 VDD1.n12 185
R1237 VDD1.n48 VDD1.n47 185
R1238 VDD1.n50 VDD1.n49 185
R1239 VDD1.n43 VDD1.n42 185
R1240 VDD1.n56 VDD1.n55 185
R1241 VDD1.n58 VDD1.n57 185
R1242 VDD1.n39 VDD1.n38 185
R1243 VDD1.n64 VDD1.n63 185
R1244 VDD1.n66 VDD1.n65 185
R1245 VDD1.n11 VDD1.t0 147.659
R1246 VDD1.n46 VDD1.t1 147.659
R1247 VDD1.n30 VDD1.n29 104.615
R1248 VDD1.n29 VDD1.n3 104.615
R1249 VDD1.n22 VDD1.n3 104.615
R1250 VDD1.n22 VDD1.n21 104.615
R1251 VDD1.n21 VDD1.n7 104.615
R1252 VDD1.n14 VDD1.n7 104.615
R1253 VDD1.n14 VDD1.n13 104.615
R1254 VDD1.n49 VDD1.n48 104.615
R1255 VDD1.n49 VDD1.n42 104.615
R1256 VDD1.n56 VDD1.n42 104.615
R1257 VDD1.n57 VDD1.n56 104.615
R1258 VDD1.n57 VDD1.n38 104.615
R1259 VDD1.n64 VDD1.n38 104.615
R1260 VDD1.n65 VDD1.n64 104.615
R1261 VDD1 VDD1.n69 85.809
R1262 VDD1.n13 VDD1.t0 52.3082
R1263 VDD1.n48 VDD1.t1 52.3082
R1264 VDD1 VDD1.n34 50.5537
R1265 VDD1.n12 VDD1.n11 15.6676
R1266 VDD1.n47 VDD1.n46 15.6676
R1267 VDD1.n15 VDD1.n10 12.8005
R1268 VDD1.n50 VDD1.n45 12.8005
R1269 VDD1.n16 VDD1.n8 12.0247
R1270 VDD1.n51 VDD1.n43 12.0247
R1271 VDD1.n20 VDD1.n19 11.249
R1272 VDD1.n55 VDD1.n54 11.249
R1273 VDD1.n23 VDD1.n6 10.4732
R1274 VDD1.n58 VDD1.n41 10.4732
R1275 VDD1.n24 VDD1.n4 9.69747
R1276 VDD1.n59 VDD1.n39 9.69747
R1277 VDD1.n34 VDD1.n33 9.45567
R1278 VDD1.n69 VDD1.n68 9.45567
R1279 VDD1.n33 VDD1.n32 9.3005
R1280 VDD1.n2 VDD1.n1 9.3005
R1281 VDD1.n27 VDD1.n26 9.3005
R1282 VDD1.n25 VDD1.n24 9.3005
R1283 VDD1.n6 VDD1.n5 9.3005
R1284 VDD1.n19 VDD1.n18 9.3005
R1285 VDD1.n17 VDD1.n16 9.3005
R1286 VDD1.n10 VDD1.n9 9.3005
R1287 VDD1.n37 VDD1.n36 9.3005
R1288 VDD1.n62 VDD1.n61 9.3005
R1289 VDD1.n60 VDD1.n59 9.3005
R1290 VDD1.n41 VDD1.n40 9.3005
R1291 VDD1.n54 VDD1.n53 9.3005
R1292 VDD1.n52 VDD1.n51 9.3005
R1293 VDD1.n45 VDD1.n44 9.3005
R1294 VDD1.n68 VDD1.n67 9.3005
R1295 VDD1.n28 VDD1.n27 8.92171
R1296 VDD1.n63 VDD1.n62 8.92171
R1297 VDD1.n31 VDD1.n2 8.14595
R1298 VDD1.n66 VDD1.n37 8.14595
R1299 VDD1.n32 VDD1.n0 7.3702
R1300 VDD1.n67 VDD1.n35 7.3702
R1301 VDD1.n34 VDD1.n0 6.59444
R1302 VDD1.n69 VDD1.n35 6.59444
R1303 VDD1.n32 VDD1.n31 5.81868
R1304 VDD1.n67 VDD1.n66 5.81868
R1305 VDD1.n28 VDD1.n2 5.04292
R1306 VDD1.n63 VDD1.n37 5.04292
R1307 VDD1.n11 VDD1.n9 4.38571
R1308 VDD1.n46 VDD1.n44 4.38571
R1309 VDD1.n27 VDD1.n4 4.26717
R1310 VDD1.n62 VDD1.n39 4.26717
R1311 VDD1.n24 VDD1.n23 3.49141
R1312 VDD1.n59 VDD1.n58 3.49141
R1313 VDD1.n20 VDD1.n6 2.71565
R1314 VDD1.n55 VDD1.n41 2.71565
R1315 VDD1.n19 VDD1.n8 1.93989
R1316 VDD1.n54 VDD1.n43 1.93989
R1317 VDD1.n16 VDD1.n15 1.16414
R1318 VDD1.n51 VDD1.n50 1.16414
R1319 VDD1.n12 VDD1.n10 0.388379
R1320 VDD1.n47 VDD1.n45 0.388379
R1321 VDD1.n33 VDD1.n1 0.155672
R1322 VDD1.n26 VDD1.n1 0.155672
R1323 VDD1.n26 VDD1.n25 0.155672
R1324 VDD1.n25 VDD1.n5 0.155672
R1325 VDD1.n18 VDD1.n5 0.155672
R1326 VDD1.n18 VDD1.n17 0.155672
R1327 VDD1.n17 VDD1.n9 0.155672
R1328 VDD1.n52 VDD1.n44 0.155672
R1329 VDD1.n53 VDD1.n52 0.155672
R1330 VDD1.n53 VDD1.n40 0.155672
R1331 VDD1.n60 VDD1.n40 0.155672
R1332 VDD1.n61 VDD1.n60 0.155672
R1333 VDD1.n61 VDD1.n36 0.155672
R1334 VDD1.n68 VDD1.n36 0.155672
R1335 VN VN.t1 141.71
R1336 VN VN.t0 101.073
R1337 VDD2.n65 VDD2.n35 289.615
R1338 VDD2.n30 VDD2.n0 289.615
R1339 VDD2.n66 VDD2.n65 185
R1340 VDD2.n64 VDD2.n63 185
R1341 VDD2.n39 VDD2.n38 185
R1342 VDD2.n58 VDD2.n57 185
R1343 VDD2.n56 VDD2.n55 185
R1344 VDD2.n43 VDD2.n42 185
R1345 VDD2.n50 VDD2.n49 185
R1346 VDD2.n48 VDD2.n47 185
R1347 VDD2.n13 VDD2.n12 185
R1348 VDD2.n15 VDD2.n14 185
R1349 VDD2.n8 VDD2.n7 185
R1350 VDD2.n21 VDD2.n20 185
R1351 VDD2.n23 VDD2.n22 185
R1352 VDD2.n4 VDD2.n3 185
R1353 VDD2.n29 VDD2.n28 185
R1354 VDD2.n31 VDD2.n30 185
R1355 VDD2.n46 VDD2.t0 147.659
R1356 VDD2.n11 VDD2.t1 147.659
R1357 VDD2.n65 VDD2.n64 104.615
R1358 VDD2.n64 VDD2.n38 104.615
R1359 VDD2.n57 VDD2.n38 104.615
R1360 VDD2.n57 VDD2.n56 104.615
R1361 VDD2.n56 VDD2.n42 104.615
R1362 VDD2.n49 VDD2.n42 104.615
R1363 VDD2.n49 VDD2.n48 104.615
R1364 VDD2.n14 VDD2.n13 104.615
R1365 VDD2.n14 VDD2.n7 104.615
R1366 VDD2.n21 VDD2.n7 104.615
R1367 VDD2.n22 VDD2.n21 104.615
R1368 VDD2.n22 VDD2.n3 104.615
R1369 VDD2.n29 VDD2.n3 104.615
R1370 VDD2.n30 VDD2.n29 104.615
R1371 VDD2.n70 VDD2.n34 84.6226
R1372 VDD2.n48 VDD2.t0 52.3082
R1373 VDD2.n13 VDD2.t1 52.3082
R1374 VDD2.n70 VDD2.n69 49.8338
R1375 VDD2.n47 VDD2.n46 15.6676
R1376 VDD2.n12 VDD2.n11 15.6676
R1377 VDD2.n50 VDD2.n45 12.8005
R1378 VDD2.n15 VDD2.n10 12.8005
R1379 VDD2.n51 VDD2.n43 12.0247
R1380 VDD2.n16 VDD2.n8 12.0247
R1381 VDD2.n55 VDD2.n54 11.249
R1382 VDD2.n20 VDD2.n19 11.249
R1383 VDD2.n58 VDD2.n41 10.4732
R1384 VDD2.n23 VDD2.n6 10.4732
R1385 VDD2.n59 VDD2.n39 9.69747
R1386 VDD2.n24 VDD2.n4 9.69747
R1387 VDD2.n69 VDD2.n68 9.45567
R1388 VDD2.n34 VDD2.n33 9.45567
R1389 VDD2.n68 VDD2.n67 9.3005
R1390 VDD2.n37 VDD2.n36 9.3005
R1391 VDD2.n62 VDD2.n61 9.3005
R1392 VDD2.n60 VDD2.n59 9.3005
R1393 VDD2.n41 VDD2.n40 9.3005
R1394 VDD2.n54 VDD2.n53 9.3005
R1395 VDD2.n52 VDD2.n51 9.3005
R1396 VDD2.n45 VDD2.n44 9.3005
R1397 VDD2.n2 VDD2.n1 9.3005
R1398 VDD2.n27 VDD2.n26 9.3005
R1399 VDD2.n25 VDD2.n24 9.3005
R1400 VDD2.n6 VDD2.n5 9.3005
R1401 VDD2.n19 VDD2.n18 9.3005
R1402 VDD2.n17 VDD2.n16 9.3005
R1403 VDD2.n10 VDD2.n9 9.3005
R1404 VDD2.n33 VDD2.n32 9.3005
R1405 VDD2.n63 VDD2.n62 8.92171
R1406 VDD2.n28 VDD2.n27 8.92171
R1407 VDD2.n66 VDD2.n37 8.14595
R1408 VDD2.n31 VDD2.n2 8.14595
R1409 VDD2.n67 VDD2.n35 7.3702
R1410 VDD2.n32 VDD2.n0 7.3702
R1411 VDD2.n69 VDD2.n35 6.59444
R1412 VDD2.n34 VDD2.n0 6.59444
R1413 VDD2.n67 VDD2.n66 5.81868
R1414 VDD2.n32 VDD2.n31 5.81868
R1415 VDD2.n63 VDD2.n37 5.04292
R1416 VDD2.n28 VDD2.n2 5.04292
R1417 VDD2.n46 VDD2.n44 4.38571
R1418 VDD2.n11 VDD2.n9 4.38571
R1419 VDD2.n62 VDD2.n39 4.26717
R1420 VDD2.n27 VDD2.n4 4.26717
R1421 VDD2.n59 VDD2.n58 3.49141
R1422 VDD2.n24 VDD2.n23 3.49141
R1423 VDD2.n55 VDD2.n41 2.71565
R1424 VDD2.n20 VDD2.n6 2.71565
R1425 VDD2.n54 VDD2.n43 1.93989
R1426 VDD2.n19 VDD2.n8 1.93989
R1427 VDD2.n51 VDD2.n50 1.16414
R1428 VDD2.n16 VDD2.n15 1.16414
R1429 VDD2 VDD2.n70 0.720328
R1430 VDD2.n47 VDD2.n45 0.388379
R1431 VDD2.n12 VDD2.n10 0.388379
R1432 VDD2.n68 VDD2.n36 0.155672
R1433 VDD2.n61 VDD2.n36 0.155672
R1434 VDD2.n61 VDD2.n60 0.155672
R1435 VDD2.n60 VDD2.n40 0.155672
R1436 VDD2.n53 VDD2.n40 0.155672
R1437 VDD2.n53 VDD2.n52 0.155672
R1438 VDD2.n52 VDD2.n44 0.155672
R1439 VDD2.n17 VDD2.n9 0.155672
R1440 VDD2.n18 VDD2.n17 0.155672
R1441 VDD2.n18 VDD2.n5 0.155672
R1442 VDD2.n25 VDD2.n5 0.155672
R1443 VDD2.n26 VDD2.n25 0.155672
R1444 VDD2.n26 VDD2.n1 0.155672
R1445 VDD2.n33 VDD2.n1 0.155672
C0 VDD2 VN 1.68911f
C1 VDD2 VDD1 0.690937f
C2 VP VN 4.55544f
C3 VP VDD1 1.87788f
C4 VTAIL VN 1.68953f
C5 VTAIL VDD1 3.71849f
C6 VDD2 VP 0.338542f
C7 VDD2 VTAIL 3.77134f
C8 VN VDD1 0.148186f
C9 VTAIL VP 1.70373f
C10 VDD2 B 3.502231f
C11 VDD1 B 5.14827f
C12 VTAIL B 5.0769f
C13 VN B 8.1622f
C14 VP B 6.100295f
C15 VDD2.n0 B 0.021321f
C16 VDD2.n1 B 0.014541f
C17 VDD2.n2 B 0.007814f
C18 VDD2.n3 B 0.018468f
C19 VDD2.n4 B 0.008273f
C20 VDD2.n5 B 0.014541f
C21 VDD2.n6 B 0.007814f
C22 VDD2.n7 B 0.018468f
C23 VDD2.n8 B 0.008273f
C24 VDD2.n9 B 0.397418f
C25 VDD2.n10 B 0.007814f
C26 VDD2.t1 B 0.030098f
C27 VDD2.n11 B 0.064951f
C28 VDD2.n12 B 0.01091f
C29 VDD2.n13 B 0.013851f
C30 VDD2.n14 B 0.018468f
C31 VDD2.n15 B 0.008273f
C32 VDD2.n16 B 0.007814f
C33 VDD2.n17 B 0.014541f
C34 VDD2.n18 B 0.014541f
C35 VDD2.n19 B 0.007814f
C36 VDD2.n20 B 0.008273f
C37 VDD2.n21 B 0.018468f
C38 VDD2.n22 B 0.018468f
C39 VDD2.n23 B 0.008273f
C40 VDD2.n24 B 0.007814f
C41 VDD2.n25 B 0.014541f
C42 VDD2.n26 B 0.014541f
C43 VDD2.n27 B 0.007814f
C44 VDD2.n28 B 0.008273f
C45 VDD2.n29 B 0.018468f
C46 VDD2.n30 B 0.041543f
C47 VDD2.n31 B 0.008273f
C48 VDD2.n32 B 0.007814f
C49 VDD2.n33 B 0.034603f
C50 VDD2.n34 B 0.328011f
C51 VDD2.n35 B 0.021321f
C52 VDD2.n36 B 0.014541f
C53 VDD2.n37 B 0.007814f
C54 VDD2.n38 B 0.018468f
C55 VDD2.n39 B 0.008273f
C56 VDD2.n40 B 0.014541f
C57 VDD2.n41 B 0.007814f
C58 VDD2.n42 B 0.018468f
C59 VDD2.n43 B 0.008273f
C60 VDD2.n44 B 0.397418f
C61 VDD2.n45 B 0.007814f
C62 VDD2.t0 B 0.030098f
C63 VDD2.n46 B 0.064951f
C64 VDD2.n47 B 0.01091f
C65 VDD2.n48 B 0.013851f
C66 VDD2.n49 B 0.018468f
C67 VDD2.n50 B 0.008273f
C68 VDD2.n51 B 0.007814f
C69 VDD2.n52 B 0.014541f
C70 VDD2.n53 B 0.014541f
C71 VDD2.n54 B 0.007814f
C72 VDD2.n55 B 0.008273f
C73 VDD2.n56 B 0.018468f
C74 VDD2.n57 B 0.018468f
C75 VDD2.n58 B 0.008273f
C76 VDD2.n59 B 0.007814f
C77 VDD2.n60 B 0.014541f
C78 VDD2.n61 B 0.014541f
C79 VDD2.n62 B 0.007814f
C80 VDD2.n63 B 0.008273f
C81 VDD2.n64 B 0.018468f
C82 VDD2.n65 B 0.041543f
C83 VDD2.n66 B 0.008273f
C84 VDD2.n67 B 0.007814f
C85 VDD2.n68 B 0.034603f
C86 VDD2.n69 B 0.033468f
C87 VDD2.n70 B 1.47605f
C88 VN.t0 B 1.13911f
C89 VN.t1 B 1.46959f
C90 VDD1.n0 B 0.020471f
C91 VDD1.n1 B 0.013961f
C92 VDD1.n2 B 0.007502f
C93 VDD1.n3 B 0.017732f
C94 VDD1.n4 B 0.007943f
C95 VDD1.n5 B 0.013961f
C96 VDD1.n6 B 0.007502f
C97 VDD1.n7 B 0.017732f
C98 VDD1.n8 B 0.007943f
C99 VDD1.n9 B 0.381567f
C100 VDD1.n10 B 0.007502f
C101 VDD1.t0 B 0.028898f
C102 VDD1.n11 B 0.06236f
C103 VDD1.n12 B 0.010475f
C104 VDD1.n13 B 0.013299f
C105 VDD1.n14 B 0.017732f
C106 VDD1.n15 B 0.007943f
C107 VDD1.n16 B 0.007502f
C108 VDD1.n17 B 0.013961f
C109 VDD1.n18 B 0.013961f
C110 VDD1.n19 B 0.007502f
C111 VDD1.n20 B 0.007943f
C112 VDD1.n21 B 0.017732f
C113 VDD1.n22 B 0.017732f
C114 VDD1.n23 B 0.007943f
C115 VDD1.n24 B 0.007502f
C116 VDD1.n25 B 0.013961f
C117 VDD1.n26 B 0.013961f
C118 VDD1.n27 B 0.007502f
C119 VDD1.n28 B 0.007943f
C120 VDD1.n29 B 0.017732f
C121 VDD1.n30 B 0.039886f
C122 VDD1.n31 B 0.007943f
C123 VDD1.n32 B 0.007502f
C124 VDD1.n33 B 0.033223f
C125 VDD1.n34 B 0.032985f
C126 VDD1.n35 B 0.020471f
C127 VDD1.n36 B 0.013961f
C128 VDD1.n37 B 0.007502f
C129 VDD1.n38 B 0.017732f
C130 VDD1.n39 B 0.007943f
C131 VDD1.n40 B 0.013961f
C132 VDD1.n41 B 0.007502f
C133 VDD1.n42 B 0.017732f
C134 VDD1.n43 B 0.007943f
C135 VDD1.n44 B 0.381567f
C136 VDD1.n45 B 0.007502f
C137 VDD1.t1 B 0.028898f
C138 VDD1.n46 B 0.06236f
C139 VDD1.n47 B 0.010475f
C140 VDD1.n48 B 0.013299f
C141 VDD1.n49 B 0.017732f
C142 VDD1.n50 B 0.007943f
C143 VDD1.n51 B 0.007502f
C144 VDD1.n52 B 0.013961f
C145 VDD1.n53 B 0.013961f
C146 VDD1.n54 B 0.007502f
C147 VDD1.n55 B 0.007943f
C148 VDD1.n56 B 0.017732f
C149 VDD1.n57 B 0.017732f
C150 VDD1.n58 B 0.007943f
C151 VDD1.n59 B 0.007502f
C152 VDD1.n60 B 0.013961f
C153 VDD1.n61 B 0.013961f
C154 VDD1.n62 B 0.007502f
C155 VDD1.n63 B 0.007943f
C156 VDD1.n64 B 0.017732f
C157 VDD1.n65 B 0.039886f
C158 VDD1.n66 B 0.007943f
C159 VDD1.n67 B 0.007502f
C160 VDD1.n68 B 0.033223f
C161 VDD1.n69 B 0.340027f
C162 VTAIL.n0 B 0.023371f
C163 VTAIL.n1 B 0.015938f
C164 VTAIL.n2 B 0.008565f
C165 VTAIL.n3 B 0.020244f
C166 VTAIL.n4 B 0.009068f
C167 VTAIL.n5 B 0.015938f
C168 VTAIL.n6 B 0.008565f
C169 VTAIL.n7 B 0.020244f
C170 VTAIL.n8 B 0.009068f
C171 VTAIL.n9 B 0.435621f
C172 VTAIL.n10 B 0.008565f
C173 VTAIL.t2 B 0.032992f
C174 VTAIL.n11 B 0.071194f
C175 VTAIL.n12 B 0.011958f
C176 VTAIL.n13 B 0.015183f
C177 VTAIL.n14 B 0.020244f
C178 VTAIL.n15 B 0.009068f
C179 VTAIL.n16 B 0.008565f
C180 VTAIL.n17 B 0.015938f
C181 VTAIL.n18 B 0.015938f
C182 VTAIL.n19 B 0.008565f
C183 VTAIL.n20 B 0.009068f
C184 VTAIL.n21 B 0.020244f
C185 VTAIL.n22 B 0.020244f
C186 VTAIL.n23 B 0.009068f
C187 VTAIL.n24 B 0.008565f
C188 VTAIL.n25 B 0.015938f
C189 VTAIL.n26 B 0.015938f
C190 VTAIL.n27 B 0.008565f
C191 VTAIL.n28 B 0.009068f
C192 VTAIL.n29 B 0.020244f
C193 VTAIL.n30 B 0.045536f
C194 VTAIL.n31 B 0.009068f
C195 VTAIL.n32 B 0.008565f
C196 VTAIL.n33 B 0.03793f
C197 VTAIL.n34 B 0.025688f
C198 VTAIL.n35 B 0.863405f
C199 VTAIL.n36 B 0.023371f
C200 VTAIL.n37 B 0.015938f
C201 VTAIL.n38 B 0.008565f
C202 VTAIL.n39 B 0.020244f
C203 VTAIL.n40 B 0.009068f
C204 VTAIL.n41 B 0.015938f
C205 VTAIL.n42 B 0.008565f
C206 VTAIL.n43 B 0.020244f
C207 VTAIL.n44 B 0.009068f
C208 VTAIL.n45 B 0.435621f
C209 VTAIL.n46 B 0.008565f
C210 VTAIL.t0 B 0.032992f
C211 VTAIL.n47 B 0.071194f
C212 VTAIL.n48 B 0.011958f
C213 VTAIL.n49 B 0.015183f
C214 VTAIL.n50 B 0.020244f
C215 VTAIL.n51 B 0.009068f
C216 VTAIL.n52 B 0.008565f
C217 VTAIL.n53 B 0.015938f
C218 VTAIL.n54 B 0.015938f
C219 VTAIL.n55 B 0.008565f
C220 VTAIL.n56 B 0.009068f
C221 VTAIL.n57 B 0.020244f
C222 VTAIL.n58 B 0.020244f
C223 VTAIL.n59 B 0.009068f
C224 VTAIL.n60 B 0.008565f
C225 VTAIL.n61 B 0.015938f
C226 VTAIL.n62 B 0.015938f
C227 VTAIL.n63 B 0.008565f
C228 VTAIL.n64 B 0.009068f
C229 VTAIL.n65 B 0.020244f
C230 VTAIL.n66 B 0.045536f
C231 VTAIL.n67 B 0.009068f
C232 VTAIL.n68 B 0.008565f
C233 VTAIL.n69 B 0.03793f
C234 VTAIL.n70 B 0.025688f
C235 VTAIL.n71 B 0.894397f
C236 VTAIL.n72 B 0.023371f
C237 VTAIL.n73 B 0.015938f
C238 VTAIL.n74 B 0.008565f
C239 VTAIL.n75 B 0.020244f
C240 VTAIL.n76 B 0.009068f
C241 VTAIL.n77 B 0.015938f
C242 VTAIL.n78 B 0.008565f
C243 VTAIL.n79 B 0.020244f
C244 VTAIL.n80 B 0.009068f
C245 VTAIL.n81 B 0.435621f
C246 VTAIL.n82 B 0.008565f
C247 VTAIL.t3 B 0.032992f
C248 VTAIL.n83 B 0.071194f
C249 VTAIL.n84 B 0.011958f
C250 VTAIL.n85 B 0.015183f
C251 VTAIL.n86 B 0.020244f
C252 VTAIL.n87 B 0.009068f
C253 VTAIL.n88 B 0.008565f
C254 VTAIL.n89 B 0.015938f
C255 VTAIL.n90 B 0.015938f
C256 VTAIL.n91 B 0.008565f
C257 VTAIL.n92 B 0.009068f
C258 VTAIL.n93 B 0.020244f
C259 VTAIL.n94 B 0.020244f
C260 VTAIL.n95 B 0.009068f
C261 VTAIL.n96 B 0.008565f
C262 VTAIL.n97 B 0.015938f
C263 VTAIL.n98 B 0.015938f
C264 VTAIL.n99 B 0.008565f
C265 VTAIL.n100 B 0.009068f
C266 VTAIL.n101 B 0.020244f
C267 VTAIL.n102 B 0.045536f
C268 VTAIL.n103 B 0.009068f
C269 VTAIL.n104 B 0.008565f
C270 VTAIL.n105 B 0.03793f
C271 VTAIL.n106 B 0.025688f
C272 VTAIL.n107 B 0.758477f
C273 VTAIL.n108 B 0.023371f
C274 VTAIL.n109 B 0.015938f
C275 VTAIL.n110 B 0.008565f
C276 VTAIL.n111 B 0.020244f
C277 VTAIL.n112 B 0.009068f
C278 VTAIL.n113 B 0.015938f
C279 VTAIL.n114 B 0.008565f
C280 VTAIL.n115 B 0.020244f
C281 VTAIL.n116 B 0.009068f
C282 VTAIL.n117 B 0.435621f
C283 VTAIL.n118 B 0.008565f
C284 VTAIL.t1 B 0.032992f
C285 VTAIL.n119 B 0.071194f
C286 VTAIL.n120 B 0.011958f
C287 VTAIL.n121 B 0.015183f
C288 VTAIL.n122 B 0.020244f
C289 VTAIL.n123 B 0.009068f
C290 VTAIL.n124 B 0.008565f
C291 VTAIL.n125 B 0.015938f
C292 VTAIL.n126 B 0.015938f
C293 VTAIL.n127 B 0.008565f
C294 VTAIL.n128 B 0.009068f
C295 VTAIL.n129 B 0.020244f
C296 VTAIL.n130 B 0.020244f
C297 VTAIL.n131 B 0.009068f
C298 VTAIL.n132 B 0.008565f
C299 VTAIL.n133 B 0.015938f
C300 VTAIL.n134 B 0.015938f
C301 VTAIL.n135 B 0.008565f
C302 VTAIL.n136 B 0.009068f
C303 VTAIL.n137 B 0.020244f
C304 VTAIL.n138 B 0.045536f
C305 VTAIL.n139 B 0.009068f
C306 VTAIL.n140 B 0.008565f
C307 VTAIL.n141 B 0.03793f
C308 VTAIL.n142 B 0.025688f
C309 VTAIL.n143 B 0.697379f
C310 VP.t0 B 1.14416f
C311 VP.t1 B 1.47669f
C312 VP.n0 B 1.92729f
.ends

